* NGSPICE file created from diff_pair_sample_1691.ext - technology: sky130A

.subckt diff_pair_sample_1691 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=7.722 pd=40.38 as=7.722 ps=40.38 w=19.8 l=0.84
X1 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=7.722 pd=40.38 as=0 ps=0 w=19.8 l=0.84
X2 VDD2.t0 VN.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=7.722 pd=40.38 as=7.722 ps=40.38 w=19.8 l=0.84
X3 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=7.722 pd=40.38 as=0 ps=0 w=19.8 l=0.84
X4 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=7.722 pd=40.38 as=0 ps=0 w=19.8 l=0.84
X5 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=7.722 pd=40.38 as=7.722 ps=40.38 w=19.8 l=0.84
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=7.722 pd=40.38 as=0 ps=0 w=19.8 l=0.84
X7 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.722 pd=40.38 as=7.722 ps=40.38 w=19.8 l=0.84
R0 VN VN.t0 822.431
R1 VN VN.t1 776.188
R2 VTAIL.n1 VTAIL.t2 46.8533
R3 VTAIL.n2 VTAIL.t0 46.8531
R4 VTAIL.n3 VTAIL.t3 46.8531
R5 VTAIL.n0 VTAIL.t1 46.8531
R6 VTAIL.n1 VTAIL.n0 31.4703
R7 VTAIL.n3 VTAIL.n2 30.4617
R8 VTAIL.n2 VTAIL.n1 0.974638
R9 VTAIL VTAIL.n0 0.780672
R10 VTAIL VTAIL.n3 0.194466
R11 VDD2.n0 VDD2.t0 106.294
R12 VDD2.n0 VDD2.t1 63.5319
R13 VDD2 VDD2.n0 0.310845
R14 B.n482 B.t6 769.774
R15 B.n479 B.t2 769.774
R16 B.n106 B.t9 769.774
R17 B.n103 B.t13 769.774
R18 B.n826 B.n825 585
R19 B.n827 B.n826 585
R20 B.n379 B.n101 585
R21 B.n378 B.n377 585
R22 B.n376 B.n375 585
R23 B.n374 B.n373 585
R24 B.n372 B.n371 585
R25 B.n370 B.n369 585
R26 B.n368 B.n367 585
R27 B.n366 B.n365 585
R28 B.n364 B.n363 585
R29 B.n362 B.n361 585
R30 B.n360 B.n359 585
R31 B.n358 B.n357 585
R32 B.n356 B.n355 585
R33 B.n354 B.n353 585
R34 B.n352 B.n351 585
R35 B.n350 B.n349 585
R36 B.n348 B.n347 585
R37 B.n346 B.n345 585
R38 B.n344 B.n343 585
R39 B.n342 B.n341 585
R40 B.n340 B.n339 585
R41 B.n338 B.n337 585
R42 B.n336 B.n335 585
R43 B.n334 B.n333 585
R44 B.n332 B.n331 585
R45 B.n330 B.n329 585
R46 B.n328 B.n327 585
R47 B.n326 B.n325 585
R48 B.n324 B.n323 585
R49 B.n322 B.n321 585
R50 B.n320 B.n319 585
R51 B.n318 B.n317 585
R52 B.n316 B.n315 585
R53 B.n314 B.n313 585
R54 B.n312 B.n311 585
R55 B.n310 B.n309 585
R56 B.n308 B.n307 585
R57 B.n306 B.n305 585
R58 B.n304 B.n303 585
R59 B.n302 B.n301 585
R60 B.n300 B.n299 585
R61 B.n298 B.n297 585
R62 B.n296 B.n295 585
R63 B.n294 B.n293 585
R64 B.n292 B.n291 585
R65 B.n290 B.n289 585
R66 B.n288 B.n287 585
R67 B.n286 B.n285 585
R68 B.n284 B.n283 585
R69 B.n282 B.n281 585
R70 B.n280 B.n279 585
R71 B.n278 B.n277 585
R72 B.n276 B.n275 585
R73 B.n274 B.n273 585
R74 B.n272 B.n271 585
R75 B.n270 B.n269 585
R76 B.n268 B.n267 585
R77 B.n266 B.n265 585
R78 B.n264 B.n263 585
R79 B.n262 B.n261 585
R80 B.n260 B.n259 585
R81 B.n258 B.n257 585
R82 B.n256 B.n255 585
R83 B.n254 B.n253 585
R84 B.n252 B.n251 585
R85 B.n250 B.n249 585
R86 B.n248 B.n247 585
R87 B.n246 B.n245 585
R88 B.n244 B.n243 585
R89 B.n242 B.n241 585
R90 B.n240 B.n239 585
R91 B.n238 B.n237 585
R92 B.n236 B.n235 585
R93 B.n233 B.n232 585
R94 B.n231 B.n230 585
R95 B.n229 B.n228 585
R96 B.n227 B.n226 585
R97 B.n225 B.n224 585
R98 B.n223 B.n222 585
R99 B.n221 B.n220 585
R100 B.n219 B.n218 585
R101 B.n217 B.n216 585
R102 B.n215 B.n214 585
R103 B.n213 B.n212 585
R104 B.n211 B.n210 585
R105 B.n209 B.n208 585
R106 B.n207 B.n206 585
R107 B.n205 B.n204 585
R108 B.n203 B.n202 585
R109 B.n201 B.n200 585
R110 B.n199 B.n198 585
R111 B.n197 B.n196 585
R112 B.n195 B.n194 585
R113 B.n193 B.n192 585
R114 B.n191 B.n190 585
R115 B.n189 B.n188 585
R116 B.n187 B.n186 585
R117 B.n185 B.n184 585
R118 B.n183 B.n182 585
R119 B.n181 B.n180 585
R120 B.n179 B.n178 585
R121 B.n177 B.n176 585
R122 B.n175 B.n174 585
R123 B.n173 B.n172 585
R124 B.n171 B.n170 585
R125 B.n169 B.n168 585
R126 B.n167 B.n166 585
R127 B.n165 B.n164 585
R128 B.n163 B.n162 585
R129 B.n161 B.n160 585
R130 B.n159 B.n158 585
R131 B.n157 B.n156 585
R132 B.n155 B.n154 585
R133 B.n153 B.n152 585
R134 B.n151 B.n150 585
R135 B.n149 B.n148 585
R136 B.n147 B.n146 585
R137 B.n145 B.n144 585
R138 B.n143 B.n142 585
R139 B.n141 B.n140 585
R140 B.n139 B.n138 585
R141 B.n137 B.n136 585
R142 B.n135 B.n134 585
R143 B.n133 B.n132 585
R144 B.n131 B.n130 585
R145 B.n129 B.n128 585
R146 B.n127 B.n126 585
R147 B.n125 B.n124 585
R148 B.n123 B.n122 585
R149 B.n121 B.n120 585
R150 B.n119 B.n118 585
R151 B.n117 B.n116 585
R152 B.n115 B.n114 585
R153 B.n113 B.n112 585
R154 B.n111 B.n110 585
R155 B.n109 B.n108 585
R156 B.n32 B.n31 585
R157 B.n830 B.n829 585
R158 B.n824 B.n102 585
R159 B.n102 B.n29 585
R160 B.n823 B.n28 585
R161 B.n834 B.n28 585
R162 B.n822 B.n27 585
R163 B.n835 B.n27 585
R164 B.n821 B.n26 585
R165 B.n836 B.n26 585
R166 B.n820 B.n819 585
R167 B.n819 B.n22 585
R168 B.n818 B.n21 585
R169 B.n842 B.n21 585
R170 B.n817 B.n20 585
R171 B.n843 B.n20 585
R172 B.n816 B.n19 585
R173 B.n844 B.n19 585
R174 B.n815 B.n814 585
R175 B.n814 B.n15 585
R176 B.n813 B.n14 585
R177 B.n850 B.n14 585
R178 B.n812 B.n13 585
R179 B.n851 B.n13 585
R180 B.n811 B.n12 585
R181 B.n852 B.n12 585
R182 B.n810 B.n809 585
R183 B.n809 B.n8 585
R184 B.n808 B.n7 585
R185 B.n858 B.n7 585
R186 B.n807 B.n6 585
R187 B.n859 B.n6 585
R188 B.n806 B.n5 585
R189 B.n860 B.n5 585
R190 B.n805 B.n804 585
R191 B.n804 B.n4 585
R192 B.n803 B.n380 585
R193 B.n803 B.n802 585
R194 B.n793 B.n381 585
R195 B.n382 B.n381 585
R196 B.n795 B.n794 585
R197 B.n796 B.n795 585
R198 B.n792 B.n387 585
R199 B.n387 B.n386 585
R200 B.n791 B.n790 585
R201 B.n790 B.n789 585
R202 B.n389 B.n388 585
R203 B.n390 B.n389 585
R204 B.n782 B.n781 585
R205 B.n783 B.n782 585
R206 B.n780 B.n395 585
R207 B.n395 B.n394 585
R208 B.n779 B.n778 585
R209 B.n778 B.n777 585
R210 B.n397 B.n396 585
R211 B.n398 B.n397 585
R212 B.n770 B.n769 585
R213 B.n771 B.n770 585
R214 B.n768 B.n403 585
R215 B.n403 B.n402 585
R216 B.n767 B.n766 585
R217 B.n766 B.n765 585
R218 B.n405 B.n404 585
R219 B.n406 B.n405 585
R220 B.n761 B.n760 585
R221 B.n409 B.n408 585
R222 B.n757 B.n756 585
R223 B.n758 B.n757 585
R224 B.n755 B.n478 585
R225 B.n754 B.n753 585
R226 B.n752 B.n751 585
R227 B.n750 B.n749 585
R228 B.n748 B.n747 585
R229 B.n746 B.n745 585
R230 B.n744 B.n743 585
R231 B.n742 B.n741 585
R232 B.n740 B.n739 585
R233 B.n738 B.n737 585
R234 B.n736 B.n735 585
R235 B.n734 B.n733 585
R236 B.n732 B.n731 585
R237 B.n730 B.n729 585
R238 B.n728 B.n727 585
R239 B.n726 B.n725 585
R240 B.n724 B.n723 585
R241 B.n722 B.n721 585
R242 B.n720 B.n719 585
R243 B.n718 B.n717 585
R244 B.n716 B.n715 585
R245 B.n714 B.n713 585
R246 B.n712 B.n711 585
R247 B.n710 B.n709 585
R248 B.n708 B.n707 585
R249 B.n706 B.n705 585
R250 B.n704 B.n703 585
R251 B.n702 B.n701 585
R252 B.n700 B.n699 585
R253 B.n698 B.n697 585
R254 B.n696 B.n695 585
R255 B.n694 B.n693 585
R256 B.n692 B.n691 585
R257 B.n690 B.n689 585
R258 B.n688 B.n687 585
R259 B.n686 B.n685 585
R260 B.n684 B.n683 585
R261 B.n682 B.n681 585
R262 B.n680 B.n679 585
R263 B.n678 B.n677 585
R264 B.n676 B.n675 585
R265 B.n674 B.n673 585
R266 B.n672 B.n671 585
R267 B.n670 B.n669 585
R268 B.n668 B.n667 585
R269 B.n666 B.n665 585
R270 B.n664 B.n663 585
R271 B.n662 B.n661 585
R272 B.n660 B.n659 585
R273 B.n658 B.n657 585
R274 B.n656 B.n655 585
R275 B.n654 B.n653 585
R276 B.n652 B.n651 585
R277 B.n650 B.n649 585
R278 B.n648 B.n647 585
R279 B.n646 B.n645 585
R280 B.n644 B.n643 585
R281 B.n642 B.n641 585
R282 B.n640 B.n639 585
R283 B.n638 B.n637 585
R284 B.n636 B.n635 585
R285 B.n634 B.n633 585
R286 B.n632 B.n631 585
R287 B.n630 B.n629 585
R288 B.n628 B.n627 585
R289 B.n626 B.n625 585
R290 B.n624 B.n623 585
R291 B.n622 B.n621 585
R292 B.n620 B.n619 585
R293 B.n618 B.n617 585
R294 B.n616 B.n615 585
R295 B.n613 B.n612 585
R296 B.n611 B.n610 585
R297 B.n609 B.n608 585
R298 B.n607 B.n606 585
R299 B.n605 B.n604 585
R300 B.n603 B.n602 585
R301 B.n601 B.n600 585
R302 B.n599 B.n598 585
R303 B.n597 B.n596 585
R304 B.n595 B.n594 585
R305 B.n593 B.n592 585
R306 B.n591 B.n590 585
R307 B.n589 B.n588 585
R308 B.n587 B.n586 585
R309 B.n585 B.n584 585
R310 B.n583 B.n582 585
R311 B.n581 B.n580 585
R312 B.n579 B.n578 585
R313 B.n577 B.n576 585
R314 B.n575 B.n574 585
R315 B.n573 B.n572 585
R316 B.n571 B.n570 585
R317 B.n569 B.n568 585
R318 B.n567 B.n566 585
R319 B.n565 B.n564 585
R320 B.n563 B.n562 585
R321 B.n561 B.n560 585
R322 B.n559 B.n558 585
R323 B.n557 B.n556 585
R324 B.n555 B.n554 585
R325 B.n553 B.n552 585
R326 B.n551 B.n550 585
R327 B.n549 B.n548 585
R328 B.n547 B.n546 585
R329 B.n545 B.n544 585
R330 B.n543 B.n542 585
R331 B.n541 B.n540 585
R332 B.n539 B.n538 585
R333 B.n537 B.n536 585
R334 B.n535 B.n534 585
R335 B.n533 B.n532 585
R336 B.n531 B.n530 585
R337 B.n529 B.n528 585
R338 B.n527 B.n526 585
R339 B.n525 B.n524 585
R340 B.n523 B.n522 585
R341 B.n521 B.n520 585
R342 B.n519 B.n518 585
R343 B.n517 B.n516 585
R344 B.n515 B.n514 585
R345 B.n513 B.n512 585
R346 B.n511 B.n510 585
R347 B.n509 B.n508 585
R348 B.n507 B.n506 585
R349 B.n505 B.n504 585
R350 B.n503 B.n502 585
R351 B.n501 B.n500 585
R352 B.n499 B.n498 585
R353 B.n497 B.n496 585
R354 B.n495 B.n494 585
R355 B.n493 B.n492 585
R356 B.n491 B.n490 585
R357 B.n489 B.n488 585
R358 B.n487 B.n486 585
R359 B.n485 B.n484 585
R360 B.n762 B.n407 585
R361 B.n407 B.n406 585
R362 B.n764 B.n763 585
R363 B.n765 B.n764 585
R364 B.n401 B.n400 585
R365 B.n402 B.n401 585
R366 B.n773 B.n772 585
R367 B.n772 B.n771 585
R368 B.n774 B.n399 585
R369 B.n399 B.n398 585
R370 B.n776 B.n775 585
R371 B.n777 B.n776 585
R372 B.n393 B.n392 585
R373 B.n394 B.n393 585
R374 B.n785 B.n784 585
R375 B.n784 B.n783 585
R376 B.n786 B.n391 585
R377 B.n391 B.n390 585
R378 B.n788 B.n787 585
R379 B.n789 B.n788 585
R380 B.n385 B.n384 585
R381 B.n386 B.n385 585
R382 B.n798 B.n797 585
R383 B.n797 B.n796 585
R384 B.n799 B.n383 585
R385 B.n383 B.n382 585
R386 B.n801 B.n800 585
R387 B.n802 B.n801 585
R388 B.n2 B.n0 585
R389 B.n4 B.n2 585
R390 B.n3 B.n1 585
R391 B.n859 B.n3 585
R392 B.n857 B.n856 585
R393 B.n858 B.n857 585
R394 B.n855 B.n9 585
R395 B.n9 B.n8 585
R396 B.n854 B.n853 585
R397 B.n853 B.n852 585
R398 B.n11 B.n10 585
R399 B.n851 B.n11 585
R400 B.n849 B.n848 585
R401 B.n850 B.n849 585
R402 B.n847 B.n16 585
R403 B.n16 B.n15 585
R404 B.n846 B.n845 585
R405 B.n845 B.n844 585
R406 B.n18 B.n17 585
R407 B.n843 B.n18 585
R408 B.n841 B.n840 585
R409 B.n842 B.n841 585
R410 B.n839 B.n23 585
R411 B.n23 B.n22 585
R412 B.n838 B.n837 585
R413 B.n837 B.n836 585
R414 B.n25 B.n24 585
R415 B.n835 B.n25 585
R416 B.n833 B.n832 585
R417 B.n834 B.n833 585
R418 B.n831 B.n30 585
R419 B.n30 B.n29 585
R420 B.n862 B.n861 585
R421 B.n861 B.n860 585
R422 B.n760 B.n407 482.89
R423 B.n829 B.n30 482.89
R424 B.n484 B.n405 482.89
R425 B.n826 B.n102 482.89
R426 B.n827 B.n100 256.663
R427 B.n827 B.n99 256.663
R428 B.n827 B.n98 256.663
R429 B.n827 B.n97 256.663
R430 B.n827 B.n96 256.663
R431 B.n827 B.n95 256.663
R432 B.n827 B.n94 256.663
R433 B.n827 B.n93 256.663
R434 B.n827 B.n92 256.663
R435 B.n827 B.n91 256.663
R436 B.n827 B.n90 256.663
R437 B.n827 B.n89 256.663
R438 B.n827 B.n88 256.663
R439 B.n827 B.n87 256.663
R440 B.n827 B.n86 256.663
R441 B.n827 B.n85 256.663
R442 B.n827 B.n84 256.663
R443 B.n827 B.n83 256.663
R444 B.n827 B.n82 256.663
R445 B.n827 B.n81 256.663
R446 B.n827 B.n80 256.663
R447 B.n827 B.n79 256.663
R448 B.n827 B.n78 256.663
R449 B.n827 B.n77 256.663
R450 B.n827 B.n76 256.663
R451 B.n827 B.n75 256.663
R452 B.n827 B.n74 256.663
R453 B.n827 B.n73 256.663
R454 B.n827 B.n72 256.663
R455 B.n827 B.n71 256.663
R456 B.n827 B.n70 256.663
R457 B.n827 B.n69 256.663
R458 B.n827 B.n68 256.663
R459 B.n827 B.n67 256.663
R460 B.n827 B.n66 256.663
R461 B.n827 B.n65 256.663
R462 B.n827 B.n64 256.663
R463 B.n827 B.n63 256.663
R464 B.n827 B.n62 256.663
R465 B.n827 B.n61 256.663
R466 B.n827 B.n60 256.663
R467 B.n827 B.n59 256.663
R468 B.n827 B.n58 256.663
R469 B.n827 B.n57 256.663
R470 B.n827 B.n56 256.663
R471 B.n827 B.n55 256.663
R472 B.n827 B.n54 256.663
R473 B.n827 B.n53 256.663
R474 B.n827 B.n52 256.663
R475 B.n827 B.n51 256.663
R476 B.n827 B.n50 256.663
R477 B.n827 B.n49 256.663
R478 B.n827 B.n48 256.663
R479 B.n827 B.n47 256.663
R480 B.n827 B.n46 256.663
R481 B.n827 B.n45 256.663
R482 B.n827 B.n44 256.663
R483 B.n827 B.n43 256.663
R484 B.n827 B.n42 256.663
R485 B.n827 B.n41 256.663
R486 B.n827 B.n40 256.663
R487 B.n827 B.n39 256.663
R488 B.n827 B.n38 256.663
R489 B.n827 B.n37 256.663
R490 B.n827 B.n36 256.663
R491 B.n827 B.n35 256.663
R492 B.n827 B.n34 256.663
R493 B.n827 B.n33 256.663
R494 B.n828 B.n827 256.663
R495 B.n759 B.n758 256.663
R496 B.n758 B.n410 256.663
R497 B.n758 B.n411 256.663
R498 B.n758 B.n412 256.663
R499 B.n758 B.n413 256.663
R500 B.n758 B.n414 256.663
R501 B.n758 B.n415 256.663
R502 B.n758 B.n416 256.663
R503 B.n758 B.n417 256.663
R504 B.n758 B.n418 256.663
R505 B.n758 B.n419 256.663
R506 B.n758 B.n420 256.663
R507 B.n758 B.n421 256.663
R508 B.n758 B.n422 256.663
R509 B.n758 B.n423 256.663
R510 B.n758 B.n424 256.663
R511 B.n758 B.n425 256.663
R512 B.n758 B.n426 256.663
R513 B.n758 B.n427 256.663
R514 B.n758 B.n428 256.663
R515 B.n758 B.n429 256.663
R516 B.n758 B.n430 256.663
R517 B.n758 B.n431 256.663
R518 B.n758 B.n432 256.663
R519 B.n758 B.n433 256.663
R520 B.n758 B.n434 256.663
R521 B.n758 B.n435 256.663
R522 B.n758 B.n436 256.663
R523 B.n758 B.n437 256.663
R524 B.n758 B.n438 256.663
R525 B.n758 B.n439 256.663
R526 B.n758 B.n440 256.663
R527 B.n758 B.n441 256.663
R528 B.n758 B.n442 256.663
R529 B.n758 B.n443 256.663
R530 B.n758 B.n444 256.663
R531 B.n758 B.n445 256.663
R532 B.n758 B.n446 256.663
R533 B.n758 B.n447 256.663
R534 B.n758 B.n448 256.663
R535 B.n758 B.n449 256.663
R536 B.n758 B.n450 256.663
R537 B.n758 B.n451 256.663
R538 B.n758 B.n452 256.663
R539 B.n758 B.n453 256.663
R540 B.n758 B.n454 256.663
R541 B.n758 B.n455 256.663
R542 B.n758 B.n456 256.663
R543 B.n758 B.n457 256.663
R544 B.n758 B.n458 256.663
R545 B.n758 B.n459 256.663
R546 B.n758 B.n460 256.663
R547 B.n758 B.n461 256.663
R548 B.n758 B.n462 256.663
R549 B.n758 B.n463 256.663
R550 B.n758 B.n464 256.663
R551 B.n758 B.n465 256.663
R552 B.n758 B.n466 256.663
R553 B.n758 B.n467 256.663
R554 B.n758 B.n468 256.663
R555 B.n758 B.n469 256.663
R556 B.n758 B.n470 256.663
R557 B.n758 B.n471 256.663
R558 B.n758 B.n472 256.663
R559 B.n758 B.n473 256.663
R560 B.n758 B.n474 256.663
R561 B.n758 B.n475 256.663
R562 B.n758 B.n476 256.663
R563 B.n758 B.n477 256.663
R564 B.n764 B.n407 163.367
R565 B.n764 B.n401 163.367
R566 B.n772 B.n401 163.367
R567 B.n772 B.n399 163.367
R568 B.n776 B.n399 163.367
R569 B.n776 B.n393 163.367
R570 B.n784 B.n393 163.367
R571 B.n784 B.n391 163.367
R572 B.n788 B.n391 163.367
R573 B.n788 B.n385 163.367
R574 B.n797 B.n385 163.367
R575 B.n797 B.n383 163.367
R576 B.n801 B.n383 163.367
R577 B.n801 B.n2 163.367
R578 B.n861 B.n2 163.367
R579 B.n861 B.n3 163.367
R580 B.n857 B.n3 163.367
R581 B.n857 B.n9 163.367
R582 B.n853 B.n9 163.367
R583 B.n853 B.n11 163.367
R584 B.n849 B.n11 163.367
R585 B.n849 B.n16 163.367
R586 B.n845 B.n16 163.367
R587 B.n845 B.n18 163.367
R588 B.n841 B.n18 163.367
R589 B.n841 B.n23 163.367
R590 B.n837 B.n23 163.367
R591 B.n837 B.n25 163.367
R592 B.n833 B.n25 163.367
R593 B.n833 B.n30 163.367
R594 B.n757 B.n409 163.367
R595 B.n757 B.n478 163.367
R596 B.n753 B.n752 163.367
R597 B.n749 B.n748 163.367
R598 B.n745 B.n744 163.367
R599 B.n741 B.n740 163.367
R600 B.n737 B.n736 163.367
R601 B.n733 B.n732 163.367
R602 B.n729 B.n728 163.367
R603 B.n725 B.n724 163.367
R604 B.n721 B.n720 163.367
R605 B.n717 B.n716 163.367
R606 B.n713 B.n712 163.367
R607 B.n709 B.n708 163.367
R608 B.n705 B.n704 163.367
R609 B.n701 B.n700 163.367
R610 B.n697 B.n696 163.367
R611 B.n693 B.n692 163.367
R612 B.n689 B.n688 163.367
R613 B.n685 B.n684 163.367
R614 B.n681 B.n680 163.367
R615 B.n677 B.n676 163.367
R616 B.n673 B.n672 163.367
R617 B.n669 B.n668 163.367
R618 B.n665 B.n664 163.367
R619 B.n661 B.n660 163.367
R620 B.n657 B.n656 163.367
R621 B.n653 B.n652 163.367
R622 B.n649 B.n648 163.367
R623 B.n645 B.n644 163.367
R624 B.n641 B.n640 163.367
R625 B.n637 B.n636 163.367
R626 B.n633 B.n632 163.367
R627 B.n629 B.n628 163.367
R628 B.n625 B.n624 163.367
R629 B.n621 B.n620 163.367
R630 B.n617 B.n616 163.367
R631 B.n612 B.n611 163.367
R632 B.n608 B.n607 163.367
R633 B.n604 B.n603 163.367
R634 B.n600 B.n599 163.367
R635 B.n596 B.n595 163.367
R636 B.n592 B.n591 163.367
R637 B.n588 B.n587 163.367
R638 B.n584 B.n583 163.367
R639 B.n580 B.n579 163.367
R640 B.n576 B.n575 163.367
R641 B.n572 B.n571 163.367
R642 B.n568 B.n567 163.367
R643 B.n564 B.n563 163.367
R644 B.n560 B.n559 163.367
R645 B.n556 B.n555 163.367
R646 B.n552 B.n551 163.367
R647 B.n548 B.n547 163.367
R648 B.n544 B.n543 163.367
R649 B.n540 B.n539 163.367
R650 B.n536 B.n535 163.367
R651 B.n532 B.n531 163.367
R652 B.n528 B.n527 163.367
R653 B.n524 B.n523 163.367
R654 B.n520 B.n519 163.367
R655 B.n516 B.n515 163.367
R656 B.n512 B.n511 163.367
R657 B.n508 B.n507 163.367
R658 B.n504 B.n503 163.367
R659 B.n500 B.n499 163.367
R660 B.n496 B.n495 163.367
R661 B.n492 B.n491 163.367
R662 B.n488 B.n487 163.367
R663 B.n766 B.n405 163.367
R664 B.n766 B.n403 163.367
R665 B.n770 B.n403 163.367
R666 B.n770 B.n397 163.367
R667 B.n778 B.n397 163.367
R668 B.n778 B.n395 163.367
R669 B.n782 B.n395 163.367
R670 B.n782 B.n389 163.367
R671 B.n790 B.n389 163.367
R672 B.n790 B.n387 163.367
R673 B.n795 B.n387 163.367
R674 B.n795 B.n381 163.367
R675 B.n803 B.n381 163.367
R676 B.n804 B.n803 163.367
R677 B.n804 B.n5 163.367
R678 B.n6 B.n5 163.367
R679 B.n7 B.n6 163.367
R680 B.n809 B.n7 163.367
R681 B.n809 B.n12 163.367
R682 B.n13 B.n12 163.367
R683 B.n14 B.n13 163.367
R684 B.n814 B.n14 163.367
R685 B.n814 B.n19 163.367
R686 B.n20 B.n19 163.367
R687 B.n21 B.n20 163.367
R688 B.n819 B.n21 163.367
R689 B.n819 B.n26 163.367
R690 B.n27 B.n26 163.367
R691 B.n28 B.n27 163.367
R692 B.n102 B.n28 163.367
R693 B.n108 B.n32 163.367
R694 B.n112 B.n111 163.367
R695 B.n116 B.n115 163.367
R696 B.n120 B.n119 163.367
R697 B.n124 B.n123 163.367
R698 B.n128 B.n127 163.367
R699 B.n132 B.n131 163.367
R700 B.n136 B.n135 163.367
R701 B.n140 B.n139 163.367
R702 B.n144 B.n143 163.367
R703 B.n148 B.n147 163.367
R704 B.n152 B.n151 163.367
R705 B.n156 B.n155 163.367
R706 B.n160 B.n159 163.367
R707 B.n164 B.n163 163.367
R708 B.n168 B.n167 163.367
R709 B.n172 B.n171 163.367
R710 B.n176 B.n175 163.367
R711 B.n180 B.n179 163.367
R712 B.n184 B.n183 163.367
R713 B.n188 B.n187 163.367
R714 B.n192 B.n191 163.367
R715 B.n196 B.n195 163.367
R716 B.n200 B.n199 163.367
R717 B.n204 B.n203 163.367
R718 B.n208 B.n207 163.367
R719 B.n212 B.n211 163.367
R720 B.n216 B.n215 163.367
R721 B.n220 B.n219 163.367
R722 B.n224 B.n223 163.367
R723 B.n228 B.n227 163.367
R724 B.n232 B.n231 163.367
R725 B.n237 B.n236 163.367
R726 B.n241 B.n240 163.367
R727 B.n245 B.n244 163.367
R728 B.n249 B.n248 163.367
R729 B.n253 B.n252 163.367
R730 B.n257 B.n256 163.367
R731 B.n261 B.n260 163.367
R732 B.n265 B.n264 163.367
R733 B.n269 B.n268 163.367
R734 B.n273 B.n272 163.367
R735 B.n277 B.n276 163.367
R736 B.n281 B.n280 163.367
R737 B.n285 B.n284 163.367
R738 B.n289 B.n288 163.367
R739 B.n293 B.n292 163.367
R740 B.n297 B.n296 163.367
R741 B.n301 B.n300 163.367
R742 B.n305 B.n304 163.367
R743 B.n309 B.n308 163.367
R744 B.n313 B.n312 163.367
R745 B.n317 B.n316 163.367
R746 B.n321 B.n320 163.367
R747 B.n325 B.n324 163.367
R748 B.n329 B.n328 163.367
R749 B.n333 B.n332 163.367
R750 B.n337 B.n336 163.367
R751 B.n341 B.n340 163.367
R752 B.n345 B.n344 163.367
R753 B.n349 B.n348 163.367
R754 B.n353 B.n352 163.367
R755 B.n357 B.n356 163.367
R756 B.n361 B.n360 163.367
R757 B.n365 B.n364 163.367
R758 B.n369 B.n368 163.367
R759 B.n373 B.n372 163.367
R760 B.n377 B.n376 163.367
R761 B.n826 B.n101 163.367
R762 B.n482 B.t8 91.3938
R763 B.n103 B.t14 91.3938
R764 B.n479 B.t5 91.3671
R765 B.n106 B.t11 91.3671
R766 B.n760 B.n759 71.676
R767 B.n478 B.n410 71.676
R768 B.n752 B.n411 71.676
R769 B.n748 B.n412 71.676
R770 B.n744 B.n413 71.676
R771 B.n740 B.n414 71.676
R772 B.n736 B.n415 71.676
R773 B.n732 B.n416 71.676
R774 B.n728 B.n417 71.676
R775 B.n724 B.n418 71.676
R776 B.n720 B.n419 71.676
R777 B.n716 B.n420 71.676
R778 B.n712 B.n421 71.676
R779 B.n708 B.n422 71.676
R780 B.n704 B.n423 71.676
R781 B.n700 B.n424 71.676
R782 B.n696 B.n425 71.676
R783 B.n692 B.n426 71.676
R784 B.n688 B.n427 71.676
R785 B.n684 B.n428 71.676
R786 B.n680 B.n429 71.676
R787 B.n676 B.n430 71.676
R788 B.n672 B.n431 71.676
R789 B.n668 B.n432 71.676
R790 B.n664 B.n433 71.676
R791 B.n660 B.n434 71.676
R792 B.n656 B.n435 71.676
R793 B.n652 B.n436 71.676
R794 B.n648 B.n437 71.676
R795 B.n644 B.n438 71.676
R796 B.n640 B.n439 71.676
R797 B.n636 B.n440 71.676
R798 B.n632 B.n441 71.676
R799 B.n628 B.n442 71.676
R800 B.n624 B.n443 71.676
R801 B.n620 B.n444 71.676
R802 B.n616 B.n445 71.676
R803 B.n611 B.n446 71.676
R804 B.n607 B.n447 71.676
R805 B.n603 B.n448 71.676
R806 B.n599 B.n449 71.676
R807 B.n595 B.n450 71.676
R808 B.n591 B.n451 71.676
R809 B.n587 B.n452 71.676
R810 B.n583 B.n453 71.676
R811 B.n579 B.n454 71.676
R812 B.n575 B.n455 71.676
R813 B.n571 B.n456 71.676
R814 B.n567 B.n457 71.676
R815 B.n563 B.n458 71.676
R816 B.n559 B.n459 71.676
R817 B.n555 B.n460 71.676
R818 B.n551 B.n461 71.676
R819 B.n547 B.n462 71.676
R820 B.n543 B.n463 71.676
R821 B.n539 B.n464 71.676
R822 B.n535 B.n465 71.676
R823 B.n531 B.n466 71.676
R824 B.n527 B.n467 71.676
R825 B.n523 B.n468 71.676
R826 B.n519 B.n469 71.676
R827 B.n515 B.n470 71.676
R828 B.n511 B.n471 71.676
R829 B.n507 B.n472 71.676
R830 B.n503 B.n473 71.676
R831 B.n499 B.n474 71.676
R832 B.n495 B.n475 71.676
R833 B.n491 B.n476 71.676
R834 B.n487 B.n477 71.676
R835 B.n829 B.n828 71.676
R836 B.n108 B.n33 71.676
R837 B.n112 B.n34 71.676
R838 B.n116 B.n35 71.676
R839 B.n120 B.n36 71.676
R840 B.n124 B.n37 71.676
R841 B.n128 B.n38 71.676
R842 B.n132 B.n39 71.676
R843 B.n136 B.n40 71.676
R844 B.n140 B.n41 71.676
R845 B.n144 B.n42 71.676
R846 B.n148 B.n43 71.676
R847 B.n152 B.n44 71.676
R848 B.n156 B.n45 71.676
R849 B.n160 B.n46 71.676
R850 B.n164 B.n47 71.676
R851 B.n168 B.n48 71.676
R852 B.n172 B.n49 71.676
R853 B.n176 B.n50 71.676
R854 B.n180 B.n51 71.676
R855 B.n184 B.n52 71.676
R856 B.n188 B.n53 71.676
R857 B.n192 B.n54 71.676
R858 B.n196 B.n55 71.676
R859 B.n200 B.n56 71.676
R860 B.n204 B.n57 71.676
R861 B.n208 B.n58 71.676
R862 B.n212 B.n59 71.676
R863 B.n216 B.n60 71.676
R864 B.n220 B.n61 71.676
R865 B.n224 B.n62 71.676
R866 B.n228 B.n63 71.676
R867 B.n232 B.n64 71.676
R868 B.n237 B.n65 71.676
R869 B.n241 B.n66 71.676
R870 B.n245 B.n67 71.676
R871 B.n249 B.n68 71.676
R872 B.n253 B.n69 71.676
R873 B.n257 B.n70 71.676
R874 B.n261 B.n71 71.676
R875 B.n265 B.n72 71.676
R876 B.n269 B.n73 71.676
R877 B.n273 B.n74 71.676
R878 B.n277 B.n75 71.676
R879 B.n281 B.n76 71.676
R880 B.n285 B.n77 71.676
R881 B.n289 B.n78 71.676
R882 B.n293 B.n79 71.676
R883 B.n297 B.n80 71.676
R884 B.n301 B.n81 71.676
R885 B.n305 B.n82 71.676
R886 B.n309 B.n83 71.676
R887 B.n313 B.n84 71.676
R888 B.n317 B.n85 71.676
R889 B.n321 B.n86 71.676
R890 B.n325 B.n87 71.676
R891 B.n329 B.n88 71.676
R892 B.n333 B.n89 71.676
R893 B.n337 B.n90 71.676
R894 B.n341 B.n91 71.676
R895 B.n345 B.n92 71.676
R896 B.n349 B.n93 71.676
R897 B.n353 B.n94 71.676
R898 B.n357 B.n95 71.676
R899 B.n361 B.n96 71.676
R900 B.n365 B.n97 71.676
R901 B.n369 B.n98 71.676
R902 B.n373 B.n99 71.676
R903 B.n377 B.n100 71.676
R904 B.n101 B.n100 71.676
R905 B.n376 B.n99 71.676
R906 B.n372 B.n98 71.676
R907 B.n368 B.n97 71.676
R908 B.n364 B.n96 71.676
R909 B.n360 B.n95 71.676
R910 B.n356 B.n94 71.676
R911 B.n352 B.n93 71.676
R912 B.n348 B.n92 71.676
R913 B.n344 B.n91 71.676
R914 B.n340 B.n90 71.676
R915 B.n336 B.n89 71.676
R916 B.n332 B.n88 71.676
R917 B.n328 B.n87 71.676
R918 B.n324 B.n86 71.676
R919 B.n320 B.n85 71.676
R920 B.n316 B.n84 71.676
R921 B.n312 B.n83 71.676
R922 B.n308 B.n82 71.676
R923 B.n304 B.n81 71.676
R924 B.n300 B.n80 71.676
R925 B.n296 B.n79 71.676
R926 B.n292 B.n78 71.676
R927 B.n288 B.n77 71.676
R928 B.n284 B.n76 71.676
R929 B.n280 B.n75 71.676
R930 B.n276 B.n74 71.676
R931 B.n272 B.n73 71.676
R932 B.n268 B.n72 71.676
R933 B.n264 B.n71 71.676
R934 B.n260 B.n70 71.676
R935 B.n256 B.n69 71.676
R936 B.n252 B.n68 71.676
R937 B.n248 B.n67 71.676
R938 B.n244 B.n66 71.676
R939 B.n240 B.n65 71.676
R940 B.n236 B.n64 71.676
R941 B.n231 B.n63 71.676
R942 B.n227 B.n62 71.676
R943 B.n223 B.n61 71.676
R944 B.n219 B.n60 71.676
R945 B.n215 B.n59 71.676
R946 B.n211 B.n58 71.676
R947 B.n207 B.n57 71.676
R948 B.n203 B.n56 71.676
R949 B.n199 B.n55 71.676
R950 B.n195 B.n54 71.676
R951 B.n191 B.n53 71.676
R952 B.n187 B.n52 71.676
R953 B.n183 B.n51 71.676
R954 B.n179 B.n50 71.676
R955 B.n175 B.n49 71.676
R956 B.n171 B.n48 71.676
R957 B.n167 B.n47 71.676
R958 B.n163 B.n46 71.676
R959 B.n159 B.n45 71.676
R960 B.n155 B.n44 71.676
R961 B.n151 B.n43 71.676
R962 B.n147 B.n42 71.676
R963 B.n143 B.n41 71.676
R964 B.n139 B.n40 71.676
R965 B.n135 B.n39 71.676
R966 B.n131 B.n38 71.676
R967 B.n127 B.n37 71.676
R968 B.n123 B.n36 71.676
R969 B.n119 B.n35 71.676
R970 B.n115 B.n34 71.676
R971 B.n111 B.n33 71.676
R972 B.n828 B.n32 71.676
R973 B.n759 B.n409 71.676
R974 B.n753 B.n410 71.676
R975 B.n749 B.n411 71.676
R976 B.n745 B.n412 71.676
R977 B.n741 B.n413 71.676
R978 B.n737 B.n414 71.676
R979 B.n733 B.n415 71.676
R980 B.n729 B.n416 71.676
R981 B.n725 B.n417 71.676
R982 B.n721 B.n418 71.676
R983 B.n717 B.n419 71.676
R984 B.n713 B.n420 71.676
R985 B.n709 B.n421 71.676
R986 B.n705 B.n422 71.676
R987 B.n701 B.n423 71.676
R988 B.n697 B.n424 71.676
R989 B.n693 B.n425 71.676
R990 B.n689 B.n426 71.676
R991 B.n685 B.n427 71.676
R992 B.n681 B.n428 71.676
R993 B.n677 B.n429 71.676
R994 B.n673 B.n430 71.676
R995 B.n669 B.n431 71.676
R996 B.n665 B.n432 71.676
R997 B.n661 B.n433 71.676
R998 B.n657 B.n434 71.676
R999 B.n653 B.n435 71.676
R1000 B.n649 B.n436 71.676
R1001 B.n645 B.n437 71.676
R1002 B.n641 B.n438 71.676
R1003 B.n637 B.n439 71.676
R1004 B.n633 B.n440 71.676
R1005 B.n629 B.n441 71.676
R1006 B.n625 B.n442 71.676
R1007 B.n621 B.n443 71.676
R1008 B.n617 B.n444 71.676
R1009 B.n612 B.n445 71.676
R1010 B.n608 B.n446 71.676
R1011 B.n604 B.n447 71.676
R1012 B.n600 B.n448 71.676
R1013 B.n596 B.n449 71.676
R1014 B.n592 B.n450 71.676
R1015 B.n588 B.n451 71.676
R1016 B.n584 B.n452 71.676
R1017 B.n580 B.n453 71.676
R1018 B.n576 B.n454 71.676
R1019 B.n572 B.n455 71.676
R1020 B.n568 B.n456 71.676
R1021 B.n564 B.n457 71.676
R1022 B.n560 B.n458 71.676
R1023 B.n556 B.n459 71.676
R1024 B.n552 B.n460 71.676
R1025 B.n548 B.n461 71.676
R1026 B.n544 B.n462 71.676
R1027 B.n540 B.n463 71.676
R1028 B.n536 B.n464 71.676
R1029 B.n532 B.n465 71.676
R1030 B.n528 B.n466 71.676
R1031 B.n524 B.n467 71.676
R1032 B.n520 B.n468 71.676
R1033 B.n516 B.n469 71.676
R1034 B.n512 B.n470 71.676
R1035 B.n508 B.n471 71.676
R1036 B.n504 B.n472 71.676
R1037 B.n500 B.n473 71.676
R1038 B.n496 B.n474 71.676
R1039 B.n492 B.n475 71.676
R1040 B.n488 B.n476 71.676
R1041 B.n484 B.n477 71.676
R1042 B.n483 B.t7 68.7029
R1043 B.n104 B.t15 68.7029
R1044 B.n480 B.t4 68.6762
R1045 B.n107 B.t12 68.6762
R1046 B.n614 B.n483 59.5399
R1047 B.n481 B.n480 59.5399
R1048 B.n234 B.n107 59.5399
R1049 B.n105 B.n104 59.5399
R1050 B.n758 B.n406 53.9156
R1051 B.n827 B.n29 53.9156
R1052 B.n831 B.n830 31.3761
R1053 B.n825 B.n824 31.3761
R1054 B.n485 B.n404 31.3761
R1055 B.n762 B.n761 31.3761
R1056 B.n765 B.n406 29.8072
R1057 B.n765 B.n402 29.8072
R1058 B.n771 B.n402 29.8072
R1059 B.n771 B.n398 29.8072
R1060 B.n777 B.n398 29.8072
R1061 B.n783 B.n394 29.8072
R1062 B.n783 B.n390 29.8072
R1063 B.n789 B.n390 29.8072
R1064 B.n789 B.n386 29.8072
R1065 B.n796 B.n386 29.8072
R1066 B.n802 B.n382 29.8072
R1067 B.n802 B.n4 29.8072
R1068 B.n860 B.n4 29.8072
R1069 B.n860 B.n859 29.8072
R1070 B.n859 B.n858 29.8072
R1071 B.n858 B.n8 29.8072
R1072 B.n852 B.n851 29.8072
R1073 B.n851 B.n850 29.8072
R1074 B.n850 B.n15 29.8072
R1075 B.n844 B.n15 29.8072
R1076 B.n844 B.n843 29.8072
R1077 B.n842 B.n22 29.8072
R1078 B.n836 B.n22 29.8072
R1079 B.n836 B.n835 29.8072
R1080 B.n835 B.n834 29.8072
R1081 B.n834 B.n29 29.8072
R1082 B.t3 B.n394 28.9306
R1083 B.n843 B.t10 28.9306
R1084 B.n483 B.n482 22.6914
R1085 B.n480 B.n479 22.6914
R1086 B.n107 B.n106 22.6914
R1087 B.n104 B.n103 22.6914
R1088 B.n796 B.t1 20.1639
R1089 B.n852 B.t0 20.1639
R1090 B B.n862 18.0485
R1091 B.n830 B.n31 10.6151
R1092 B.n109 B.n31 10.6151
R1093 B.n110 B.n109 10.6151
R1094 B.n113 B.n110 10.6151
R1095 B.n114 B.n113 10.6151
R1096 B.n117 B.n114 10.6151
R1097 B.n118 B.n117 10.6151
R1098 B.n121 B.n118 10.6151
R1099 B.n122 B.n121 10.6151
R1100 B.n125 B.n122 10.6151
R1101 B.n126 B.n125 10.6151
R1102 B.n129 B.n126 10.6151
R1103 B.n130 B.n129 10.6151
R1104 B.n133 B.n130 10.6151
R1105 B.n134 B.n133 10.6151
R1106 B.n137 B.n134 10.6151
R1107 B.n138 B.n137 10.6151
R1108 B.n141 B.n138 10.6151
R1109 B.n142 B.n141 10.6151
R1110 B.n145 B.n142 10.6151
R1111 B.n146 B.n145 10.6151
R1112 B.n149 B.n146 10.6151
R1113 B.n150 B.n149 10.6151
R1114 B.n153 B.n150 10.6151
R1115 B.n154 B.n153 10.6151
R1116 B.n157 B.n154 10.6151
R1117 B.n158 B.n157 10.6151
R1118 B.n161 B.n158 10.6151
R1119 B.n162 B.n161 10.6151
R1120 B.n165 B.n162 10.6151
R1121 B.n166 B.n165 10.6151
R1122 B.n169 B.n166 10.6151
R1123 B.n170 B.n169 10.6151
R1124 B.n173 B.n170 10.6151
R1125 B.n174 B.n173 10.6151
R1126 B.n177 B.n174 10.6151
R1127 B.n178 B.n177 10.6151
R1128 B.n181 B.n178 10.6151
R1129 B.n182 B.n181 10.6151
R1130 B.n185 B.n182 10.6151
R1131 B.n186 B.n185 10.6151
R1132 B.n189 B.n186 10.6151
R1133 B.n190 B.n189 10.6151
R1134 B.n193 B.n190 10.6151
R1135 B.n194 B.n193 10.6151
R1136 B.n197 B.n194 10.6151
R1137 B.n198 B.n197 10.6151
R1138 B.n201 B.n198 10.6151
R1139 B.n202 B.n201 10.6151
R1140 B.n205 B.n202 10.6151
R1141 B.n206 B.n205 10.6151
R1142 B.n209 B.n206 10.6151
R1143 B.n210 B.n209 10.6151
R1144 B.n213 B.n210 10.6151
R1145 B.n214 B.n213 10.6151
R1146 B.n217 B.n214 10.6151
R1147 B.n218 B.n217 10.6151
R1148 B.n221 B.n218 10.6151
R1149 B.n222 B.n221 10.6151
R1150 B.n225 B.n222 10.6151
R1151 B.n226 B.n225 10.6151
R1152 B.n229 B.n226 10.6151
R1153 B.n230 B.n229 10.6151
R1154 B.n233 B.n230 10.6151
R1155 B.n238 B.n235 10.6151
R1156 B.n239 B.n238 10.6151
R1157 B.n242 B.n239 10.6151
R1158 B.n243 B.n242 10.6151
R1159 B.n246 B.n243 10.6151
R1160 B.n247 B.n246 10.6151
R1161 B.n250 B.n247 10.6151
R1162 B.n251 B.n250 10.6151
R1163 B.n255 B.n254 10.6151
R1164 B.n258 B.n255 10.6151
R1165 B.n259 B.n258 10.6151
R1166 B.n262 B.n259 10.6151
R1167 B.n263 B.n262 10.6151
R1168 B.n266 B.n263 10.6151
R1169 B.n267 B.n266 10.6151
R1170 B.n270 B.n267 10.6151
R1171 B.n271 B.n270 10.6151
R1172 B.n274 B.n271 10.6151
R1173 B.n275 B.n274 10.6151
R1174 B.n278 B.n275 10.6151
R1175 B.n279 B.n278 10.6151
R1176 B.n282 B.n279 10.6151
R1177 B.n283 B.n282 10.6151
R1178 B.n286 B.n283 10.6151
R1179 B.n287 B.n286 10.6151
R1180 B.n290 B.n287 10.6151
R1181 B.n291 B.n290 10.6151
R1182 B.n294 B.n291 10.6151
R1183 B.n295 B.n294 10.6151
R1184 B.n298 B.n295 10.6151
R1185 B.n299 B.n298 10.6151
R1186 B.n302 B.n299 10.6151
R1187 B.n303 B.n302 10.6151
R1188 B.n306 B.n303 10.6151
R1189 B.n307 B.n306 10.6151
R1190 B.n310 B.n307 10.6151
R1191 B.n311 B.n310 10.6151
R1192 B.n314 B.n311 10.6151
R1193 B.n315 B.n314 10.6151
R1194 B.n318 B.n315 10.6151
R1195 B.n319 B.n318 10.6151
R1196 B.n322 B.n319 10.6151
R1197 B.n323 B.n322 10.6151
R1198 B.n326 B.n323 10.6151
R1199 B.n327 B.n326 10.6151
R1200 B.n330 B.n327 10.6151
R1201 B.n331 B.n330 10.6151
R1202 B.n334 B.n331 10.6151
R1203 B.n335 B.n334 10.6151
R1204 B.n338 B.n335 10.6151
R1205 B.n339 B.n338 10.6151
R1206 B.n342 B.n339 10.6151
R1207 B.n343 B.n342 10.6151
R1208 B.n346 B.n343 10.6151
R1209 B.n347 B.n346 10.6151
R1210 B.n350 B.n347 10.6151
R1211 B.n351 B.n350 10.6151
R1212 B.n354 B.n351 10.6151
R1213 B.n355 B.n354 10.6151
R1214 B.n358 B.n355 10.6151
R1215 B.n359 B.n358 10.6151
R1216 B.n362 B.n359 10.6151
R1217 B.n363 B.n362 10.6151
R1218 B.n366 B.n363 10.6151
R1219 B.n367 B.n366 10.6151
R1220 B.n370 B.n367 10.6151
R1221 B.n371 B.n370 10.6151
R1222 B.n374 B.n371 10.6151
R1223 B.n375 B.n374 10.6151
R1224 B.n378 B.n375 10.6151
R1225 B.n379 B.n378 10.6151
R1226 B.n825 B.n379 10.6151
R1227 B.n767 B.n404 10.6151
R1228 B.n768 B.n767 10.6151
R1229 B.n769 B.n768 10.6151
R1230 B.n769 B.n396 10.6151
R1231 B.n779 B.n396 10.6151
R1232 B.n780 B.n779 10.6151
R1233 B.n781 B.n780 10.6151
R1234 B.n781 B.n388 10.6151
R1235 B.n791 B.n388 10.6151
R1236 B.n792 B.n791 10.6151
R1237 B.n794 B.n792 10.6151
R1238 B.n794 B.n793 10.6151
R1239 B.n793 B.n380 10.6151
R1240 B.n805 B.n380 10.6151
R1241 B.n806 B.n805 10.6151
R1242 B.n807 B.n806 10.6151
R1243 B.n808 B.n807 10.6151
R1244 B.n810 B.n808 10.6151
R1245 B.n811 B.n810 10.6151
R1246 B.n812 B.n811 10.6151
R1247 B.n813 B.n812 10.6151
R1248 B.n815 B.n813 10.6151
R1249 B.n816 B.n815 10.6151
R1250 B.n817 B.n816 10.6151
R1251 B.n818 B.n817 10.6151
R1252 B.n820 B.n818 10.6151
R1253 B.n821 B.n820 10.6151
R1254 B.n822 B.n821 10.6151
R1255 B.n823 B.n822 10.6151
R1256 B.n824 B.n823 10.6151
R1257 B.n761 B.n408 10.6151
R1258 B.n756 B.n408 10.6151
R1259 B.n756 B.n755 10.6151
R1260 B.n755 B.n754 10.6151
R1261 B.n754 B.n751 10.6151
R1262 B.n751 B.n750 10.6151
R1263 B.n750 B.n747 10.6151
R1264 B.n747 B.n746 10.6151
R1265 B.n746 B.n743 10.6151
R1266 B.n743 B.n742 10.6151
R1267 B.n742 B.n739 10.6151
R1268 B.n739 B.n738 10.6151
R1269 B.n738 B.n735 10.6151
R1270 B.n735 B.n734 10.6151
R1271 B.n734 B.n731 10.6151
R1272 B.n731 B.n730 10.6151
R1273 B.n730 B.n727 10.6151
R1274 B.n727 B.n726 10.6151
R1275 B.n726 B.n723 10.6151
R1276 B.n723 B.n722 10.6151
R1277 B.n722 B.n719 10.6151
R1278 B.n719 B.n718 10.6151
R1279 B.n718 B.n715 10.6151
R1280 B.n715 B.n714 10.6151
R1281 B.n714 B.n711 10.6151
R1282 B.n711 B.n710 10.6151
R1283 B.n710 B.n707 10.6151
R1284 B.n707 B.n706 10.6151
R1285 B.n706 B.n703 10.6151
R1286 B.n703 B.n702 10.6151
R1287 B.n702 B.n699 10.6151
R1288 B.n699 B.n698 10.6151
R1289 B.n698 B.n695 10.6151
R1290 B.n695 B.n694 10.6151
R1291 B.n694 B.n691 10.6151
R1292 B.n691 B.n690 10.6151
R1293 B.n690 B.n687 10.6151
R1294 B.n687 B.n686 10.6151
R1295 B.n686 B.n683 10.6151
R1296 B.n683 B.n682 10.6151
R1297 B.n682 B.n679 10.6151
R1298 B.n679 B.n678 10.6151
R1299 B.n678 B.n675 10.6151
R1300 B.n675 B.n674 10.6151
R1301 B.n674 B.n671 10.6151
R1302 B.n671 B.n670 10.6151
R1303 B.n670 B.n667 10.6151
R1304 B.n667 B.n666 10.6151
R1305 B.n666 B.n663 10.6151
R1306 B.n663 B.n662 10.6151
R1307 B.n662 B.n659 10.6151
R1308 B.n659 B.n658 10.6151
R1309 B.n658 B.n655 10.6151
R1310 B.n655 B.n654 10.6151
R1311 B.n654 B.n651 10.6151
R1312 B.n651 B.n650 10.6151
R1313 B.n650 B.n647 10.6151
R1314 B.n647 B.n646 10.6151
R1315 B.n646 B.n643 10.6151
R1316 B.n643 B.n642 10.6151
R1317 B.n642 B.n639 10.6151
R1318 B.n639 B.n638 10.6151
R1319 B.n638 B.n635 10.6151
R1320 B.n635 B.n634 10.6151
R1321 B.n631 B.n630 10.6151
R1322 B.n630 B.n627 10.6151
R1323 B.n627 B.n626 10.6151
R1324 B.n626 B.n623 10.6151
R1325 B.n623 B.n622 10.6151
R1326 B.n622 B.n619 10.6151
R1327 B.n619 B.n618 10.6151
R1328 B.n618 B.n615 10.6151
R1329 B.n613 B.n610 10.6151
R1330 B.n610 B.n609 10.6151
R1331 B.n609 B.n606 10.6151
R1332 B.n606 B.n605 10.6151
R1333 B.n605 B.n602 10.6151
R1334 B.n602 B.n601 10.6151
R1335 B.n601 B.n598 10.6151
R1336 B.n598 B.n597 10.6151
R1337 B.n597 B.n594 10.6151
R1338 B.n594 B.n593 10.6151
R1339 B.n593 B.n590 10.6151
R1340 B.n590 B.n589 10.6151
R1341 B.n589 B.n586 10.6151
R1342 B.n586 B.n585 10.6151
R1343 B.n585 B.n582 10.6151
R1344 B.n582 B.n581 10.6151
R1345 B.n581 B.n578 10.6151
R1346 B.n578 B.n577 10.6151
R1347 B.n577 B.n574 10.6151
R1348 B.n574 B.n573 10.6151
R1349 B.n573 B.n570 10.6151
R1350 B.n570 B.n569 10.6151
R1351 B.n569 B.n566 10.6151
R1352 B.n566 B.n565 10.6151
R1353 B.n565 B.n562 10.6151
R1354 B.n562 B.n561 10.6151
R1355 B.n561 B.n558 10.6151
R1356 B.n558 B.n557 10.6151
R1357 B.n557 B.n554 10.6151
R1358 B.n554 B.n553 10.6151
R1359 B.n553 B.n550 10.6151
R1360 B.n550 B.n549 10.6151
R1361 B.n549 B.n546 10.6151
R1362 B.n546 B.n545 10.6151
R1363 B.n545 B.n542 10.6151
R1364 B.n542 B.n541 10.6151
R1365 B.n541 B.n538 10.6151
R1366 B.n538 B.n537 10.6151
R1367 B.n537 B.n534 10.6151
R1368 B.n534 B.n533 10.6151
R1369 B.n533 B.n530 10.6151
R1370 B.n530 B.n529 10.6151
R1371 B.n529 B.n526 10.6151
R1372 B.n526 B.n525 10.6151
R1373 B.n525 B.n522 10.6151
R1374 B.n522 B.n521 10.6151
R1375 B.n521 B.n518 10.6151
R1376 B.n518 B.n517 10.6151
R1377 B.n517 B.n514 10.6151
R1378 B.n514 B.n513 10.6151
R1379 B.n513 B.n510 10.6151
R1380 B.n510 B.n509 10.6151
R1381 B.n509 B.n506 10.6151
R1382 B.n506 B.n505 10.6151
R1383 B.n505 B.n502 10.6151
R1384 B.n502 B.n501 10.6151
R1385 B.n501 B.n498 10.6151
R1386 B.n498 B.n497 10.6151
R1387 B.n497 B.n494 10.6151
R1388 B.n494 B.n493 10.6151
R1389 B.n493 B.n490 10.6151
R1390 B.n490 B.n489 10.6151
R1391 B.n489 B.n486 10.6151
R1392 B.n486 B.n485 10.6151
R1393 B.n763 B.n762 10.6151
R1394 B.n763 B.n400 10.6151
R1395 B.n773 B.n400 10.6151
R1396 B.n774 B.n773 10.6151
R1397 B.n775 B.n774 10.6151
R1398 B.n775 B.n392 10.6151
R1399 B.n785 B.n392 10.6151
R1400 B.n786 B.n785 10.6151
R1401 B.n787 B.n786 10.6151
R1402 B.n787 B.n384 10.6151
R1403 B.n798 B.n384 10.6151
R1404 B.n799 B.n798 10.6151
R1405 B.n800 B.n799 10.6151
R1406 B.n800 B.n0 10.6151
R1407 B.n856 B.n1 10.6151
R1408 B.n856 B.n855 10.6151
R1409 B.n855 B.n854 10.6151
R1410 B.n854 B.n10 10.6151
R1411 B.n848 B.n10 10.6151
R1412 B.n848 B.n847 10.6151
R1413 B.n847 B.n846 10.6151
R1414 B.n846 B.n17 10.6151
R1415 B.n840 B.n17 10.6151
R1416 B.n840 B.n839 10.6151
R1417 B.n839 B.n838 10.6151
R1418 B.n838 B.n24 10.6151
R1419 B.n832 B.n24 10.6151
R1420 B.n832 B.n831 10.6151
R1421 B.t1 B.n382 9.64386
R1422 B.t0 B.n8 9.64386
R1423 B.n235 B.n234 7.18099
R1424 B.n251 B.n105 7.18099
R1425 B.n631 B.n481 7.18099
R1426 B.n615 B.n614 7.18099
R1427 B.n234 B.n233 3.43465
R1428 B.n254 B.n105 3.43465
R1429 B.n634 B.n481 3.43465
R1430 B.n614 B.n613 3.43465
R1431 B.n862 B.n0 2.81026
R1432 B.n862 B.n1 2.81026
R1433 B.n777 B.t3 0.877169
R1434 B.t10 B.n842 0.877169
R1435 VP.n0 VP.t0 822.051
R1436 VP.n0 VP.t1 776.138
R1437 VP VP.n0 0.0516364
R1438 VDD1 VDD1.t0 107.072
R1439 VDD1 VDD1.t1 63.8423
C0 VP VTAIL 2.52356f
C1 VDD2 VN 3.3366f
C2 VDD2 VTAIL 8.206f
C3 VN VTAIL 2.5087f
C4 VDD1 VP 3.44322f
C5 VDD1 VDD2 0.477838f
C6 VDD1 VN 0.148986f
C7 VDD1 VTAIL 8.174701f
C8 VDD2 VP 0.262271f
C9 VN VP 6.06731f
C10 VDD2 B 5.211534f
C11 VDD1 B 8.66966f
C12 VTAIL B 9.453226f
C13 VN B 11.204141f
C14 VP B 4.731881f
C15 VDD1.t1 B 3.75963f
C16 VDD1.t0 B 4.46368f
C17 VP.t0 B 2.88194f
C18 VP.t1 B 2.69874f
C19 VP.n0 B 6.39618f
C20 VDD2.t0 B 4.42554f
C21 VDD2.t1 B 3.7505f
C22 VDD2.n0 B 3.2697f
C23 VTAIL.t1 B 3.56663f
C24 VTAIL.n0 B 1.80323f
C25 VTAIL.t2 B 3.56663f
C26 VTAIL.n1 B 1.81564f
C27 VTAIL.t0 B 3.56663f
C28 VTAIL.n2 B 1.7511f
C29 VTAIL.t3 B 3.56663f
C30 VTAIL.n3 B 1.70117f
C31 VN.t1 B 2.65972f
C32 VN.t0 B 2.84356f
.ends

