* NGSPICE file created from diff_pair_sample_0503.ext - technology: sky130A

.subckt diff_pair_sample_0503 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1650_n2202# sky130_fd_pr__pfet_01v8 ad=2.4063 pd=13.12 as=0 ps=0 w=6.17 l=1.37
X1 B.t8 B.t6 B.t7 w_n1650_n2202# sky130_fd_pr__pfet_01v8 ad=2.4063 pd=13.12 as=0 ps=0 w=6.17 l=1.37
X2 VDD2.t1 VN.t0 VTAIL.t3 w_n1650_n2202# sky130_fd_pr__pfet_01v8 ad=2.4063 pd=13.12 as=2.4063 ps=13.12 w=6.17 l=1.37
X3 VDD2.t0 VN.t1 VTAIL.t2 w_n1650_n2202# sky130_fd_pr__pfet_01v8 ad=2.4063 pd=13.12 as=2.4063 ps=13.12 w=6.17 l=1.37
X4 B.t5 B.t3 B.t4 w_n1650_n2202# sky130_fd_pr__pfet_01v8 ad=2.4063 pd=13.12 as=0 ps=0 w=6.17 l=1.37
X5 VDD1.t1 VP.t0 VTAIL.t1 w_n1650_n2202# sky130_fd_pr__pfet_01v8 ad=2.4063 pd=13.12 as=2.4063 ps=13.12 w=6.17 l=1.37
X6 B.t2 B.t0 B.t1 w_n1650_n2202# sky130_fd_pr__pfet_01v8 ad=2.4063 pd=13.12 as=0 ps=0 w=6.17 l=1.37
X7 VDD1.t0 VP.t1 VTAIL.t0 w_n1650_n2202# sky130_fd_pr__pfet_01v8 ad=2.4063 pd=13.12 as=2.4063 ps=13.12 w=6.17 l=1.37
R0 B.n275 B.n44 585
R1 B.n277 B.n276 585
R2 B.n278 B.n43 585
R3 B.n280 B.n279 585
R4 B.n281 B.n42 585
R5 B.n283 B.n282 585
R6 B.n284 B.n41 585
R7 B.n286 B.n285 585
R8 B.n287 B.n40 585
R9 B.n289 B.n288 585
R10 B.n290 B.n39 585
R11 B.n292 B.n291 585
R12 B.n293 B.n38 585
R13 B.n295 B.n294 585
R14 B.n296 B.n37 585
R15 B.n298 B.n297 585
R16 B.n299 B.n36 585
R17 B.n301 B.n300 585
R18 B.n302 B.n35 585
R19 B.n304 B.n303 585
R20 B.n305 B.n34 585
R21 B.n307 B.n306 585
R22 B.n308 B.n33 585
R23 B.n310 B.n309 585
R24 B.n312 B.n311 585
R25 B.n313 B.n29 585
R26 B.n315 B.n314 585
R27 B.n316 B.n28 585
R28 B.n318 B.n317 585
R29 B.n319 B.n27 585
R30 B.n321 B.n320 585
R31 B.n322 B.n26 585
R32 B.n324 B.n323 585
R33 B.n325 B.n23 585
R34 B.n328 B.n327 585
R35 B.n329 B.n22 585
R36 B.n331 B.n330 585
R37 B.n332 B.n21 585
R38 B.n334 B.n333 585
R39 B.n335 B.n20 585
R40 B.n337 B.n336 585
R41 B.n338 B.n19 585
R42 B.n340 B.n339 585
R43 B.n341 B.n18 585
R44 B.n343 B.n342 585
R45 B.n344 B.n17 585
R46 B.n346 B.n345 585
R47 B.n347 B.n16 585
R48 B.n349 B.n348 585
R49 B.n350 B.n15 585
R50 B.n352 B.n351 585
R51 B.n353 B.n14 585
R52 B.n355 B.n354 585
R53 B.n356 B.n13 585
R54 B.n358 B.n357 585
R55 B.n359 B.n12 585
R56 B.n361 B.n360 585
R57 B.n362 B.n11 585
R58 B.n274 B.n273 585
R59 B.n272 B.n45 585
R60 B.n271 B.n270 585
R61 B.n269 B.n46 585
R62 B.n268 B.n267 585
R63 B.n266 B.n47 585
R64 B.n265 B.n264 585
R65 B.n263 B.n48 585
R66 B.n262 B.n261 585
R67 B.n260 B.n49 585
R68 B.n259 B.n258 585
R69 B.n257 B.n50 585
R70 B.n256 B.n255 585
R71 B.n254 B.n51 585
R72 B.n253 B.n252 585
R73 B.n251 B.n52 585
R74 B.n250 B.n249 585
R75 B.n248 B.n53 585
R76 B.n247 B.n246 585
R77 B.n245 B.n54 585
R78 B.n244 B.n243 585
R79 B.n242 B.n55 585
R80 B.n241 B.n240 585
R81 B.n239 B.n56 585
R82 B.n238 B.n237 585
R83 B.n236 B.n57 585
R84 B.n235 B.n234 585
R85 B.n233 B.n58 585
R86 B.n232 B.n231 585
R87 B.n230 B.n59 585
R88 B.n229 B.n228 585
R89 B.n227 B.n60 585
R90 B.n226 B.n225 585
R91 B.n224 B.n61 585
R92 B.n223 B.n222 585
R93 B.n221 B.n62 585
R94 B.n220 B.n219 585
R95 B.n131 B.n96 585
R96 B.n133 B.n132 585
R97 B.n134 B.n95 585
R98 B.n136 B.n135 585
R99 B.n137 B.n94 585
R100 B.n139 B.n138 585
R101 B.n140 B.n93 585
R102 B.n142 B.n141 585
R103 B.n143 B.n92 585
R104 B.n145 B.n144 585
R105 B.n146 B.n91 585
R106 B.n148 B.n147 585
R107 B.n149 B.n90 585
R108 B.n151 B.n150 585
R109 B.n152 B.n89 585
R110 B.n154 B.n153 585
R111 B.n155 B.n88 585
R112 B.n157 B.n156 585
R113 B.n158 B.n87 585
R114 B.n160 B.n159 585
R115 B.n161 B.n86 585
R116 B.n163 B.n162 585
R117 B.n164 B.n85 585
R118 B.n166 B.n165 585
R119 B.n168 B.n167 585
R120 B.n169 B.n81 585
R121 B.n171 B.n170 585
R122 B.n172 B.n80 585
R123 B.n174 B.n173 585
R124 B.n175 B.n79 585
R125 B.n177 B.n176 585
R126 B.n178 B.n78 585
R127 B.n180 B.n179 585
R128 B.n181 B.n75 585
R129 B.n184 B.n183 585
R130 B.n185 B.n74 585
R131 B.n187 B.n186 585
R132 B.n188 B.n73 585
R133 B.n190 B.n189 585
R134 B.n191 B.n72 585
R135 B.n193 B.n192 585
R136 B.n194 B.n71 585
R137 B.n196 B.n195 585
R138 B.n197 B.n70 585
R139 B.n199 B.n198 585
R140 B.n200 B.n69 585
R141 B.n202 B.n201 585
R142 B.n203 B.n68 585
R143 B.n205 B.n204 585
R144 B.n206 B.n67 585
R145 B.n208 B.n207 585
R146 B.n209 B.n66 585
R147 B.n211 B.n210 585
R148 B.n212 B.n65 585
R149 B.n214 B.n213 585
R150 B.n215 B.n64 585
R151 B.n217 B.n216 585
R152 B.n218 B.n63 585
R153 B.n130 B.n129 585
R154 B.n128 B.n97 585
R155 B.n127 B.n126 585
R156 B.n125 B.n98 585
R157 B.n124 B.n123 585
R158 B.n122 B.n99 585
R159 B.n121 B.n120 585
R160 B.n119 B.n100 585
R161 B.n118 B.n117 585
R162 B.n116 B.n101 585
R163 B.n115 B.n114 585
R164 B.n113 B.n102 585
R165 B.n112 B.n111 585
R166 B.n110 B.n103 585
R167 B.n109 B.n108 585
R168 B.n107 B.n104 585
R169 B.n106 B.n105 585
R170 B.n2 B.n0 585
R171 B.n389 B.n1 585
R172 B.n388 B.n387 585
R173 B.n386 B.n3 585
R174 B.n385 B.n384 585
R175 B.n383 B.n4 585
R176 B.n382 B.n381 585
R177 B.n380 B.n5 585
R178 B.n379 B.n378 585
R179 B.n377 B.n6 585
R180 B.n376 B.n375 585
R181 B.n374 B.n7 585
R182 B.n373 B.n372 585
R183 B.n371 B.n8 585
R184 B.n370 B.n369 585
R185 B.n368 B.n9 585
R186 B.n367 B.n366 585
R187 B.n365 B.n10 585
R188 B.n364 B.n363 585
R189 B.n391 B.n390 585
R190 B.n131 B.n130 559.769
R191 B.n364 B.n11 559.769
R192 B.n220 B.n63 559.769
R193 B.n275 B.n274 559.769
R194 B.n76 B.t0 313.459
R195 B.n82 B.t6 313.459
R196 B.n24 B.t3 313.459
R197 B.n30 B.t9 313.459
R198 B.n130 B.n97 163.367
R199 B.n126 B.n97 163.367
R200 B.n126 B.n125 163.367
R201 B.n125 B.n124 163.367
R202 B.n124 B.n99 163.367
R203 B.n120 B.n99 163.367
R204 B.n120 B.n119 163.367
R205 B.n119 B.n118 163.367
R206 B.n118 B.n101 163.367
R207 B.n114 B.n101 163.367
R208 B.n114 B.n113 163.367
R209 B.n113 B.n112 163.367
R210 B.n112 B.n103 163.367
R211 B.n108 B.n103 163.367
R212 B.n108 B.n107 163.367
R213 B.n107 B.n106 163.367
R214 B.n106 B.n2 163.367
R215 B.n390 B.n2 163.367
R216 B.n390 B.n389 163.367
R217 B.n389 B.n388 163.367
R218 B.n388 B.n3 163.367
R219 B.n384 B.n3 163.367
R220 B.n384 B.n383 163.367
R221 B.n383 B.n382 163.367
R222 B.n382 B.n5 163.367
R223 B.n378 B.n5 163.367
R224 B.n378 B.n377 163.367
R225 B.n377 B.n376 163.367
R226 B.n376 B.n7 163.367
R227 B.n372 B.n7 163.367
R228 B.n372 B.n371 163.367
R229 B.n371 B.n370 163.367
R230 B.n370 B.n9 163.367
R231 B.n366 B.n9 163.367
R232 B.n366 B.n365 163.367
R233 B.n365 B.n364 163.367
R234 B.n132 B.n131 163.367
R235 B.n132 B.n95 163.367
R236 B.n136 B.n95 163.367
R237 B.n137 B.n136 163.367
R238 B.n138 B.n137 163.367
R239 B.n138 B.n93 163.367
R240 B.n142 B.n93 163.367
R241 B.n143 B.n142 163.367
R242 B.n144 B.n143 163.367
R243 B.n144 B.n91 163.367
R244 B.n148 B.n91 163.367
R245 B.n149 B.n148 163.367
R246 B.n150 B.n149 163.367
R247 B.n150 B.n89 163.367
R248 B.n154 B.n89 163.367
R249 B.n155 B.n154 163.367
R250 B.n156 B.n155 163.367
R251 B.n156 B.n87 163.367
R252 B.n160 B.n87 163.367
R253 B.n161 B.n160 163.367
R254 B.n162 B.n161 163.367
R255 B.n162 B.n85 163.367
R256 B.n166 B.n85 163.367
R257 B.n167 B.n166 163.367
R258 B.n167 B.n81 163.367
R259 B.n171 B.n81 163.367
R260 B.n172 B.n171 163.367
R261 B.n173 B.n172 163.367
R262 B.n173 B.n79 163.367
R263 B.n177 B.n79 163.367
R264 B.n178 B.n177 163.367
R265 B.n179 B.n178 163.367
R266 B.n179 B.n75 163.367
R267 B.n184 B.n75 163.367
R268 B.n185 B.n184 163.367
R269 B.n186 B.n185 163.367
R270 B.n186 B.n73 163.367
R271 B.n190 B.n73 163.367
R272 B.n191 B.n190 163.367
R273 B.n192 B.n191 163.367
R274 B.n192 B.n71 163.367
R275 B.n196 B.n71 163.367
R276 B.n197 B.n196 163.367
R277 B.n198 B.n197 163.367
R278 B.n198 B.n69 163.367
R279 B.n202 B.n69 163.367
R280 B.n203 B.n202 163.367
R281 B.n204 B.n203 163.367
R282 B.n204 B.n67 163.367
R283 B.n208 B.n67 163.367
R284 B.n209 B.n208 163.367
R285 B.n210 B.n209 163.367
R286 B.n210 B.n65 163.367
R287 B.n214 B.n65 163.367
R288 B.n215 B.n214 163.367
R289 B.n216 B.n215 163.367
R290 B.n216 B.n63 163.367
R291 B.n221 B.n220 163.367
R292 B.n222 B.n221 163.367
R293 B.n222 B.n61 163.367
R294 B.n226 B.n61 163.367
R295 B.n227 B.n226 163.367
R296 B.n228 B.n227 163.367
R297 B.n228 B.n59 163.367
R298 B.n232 B.n59 163.367
R299 B.n233 B.n232 163.367
R300 B.n234 B.n233 163.367
R301 B.n234 B.n57 163.367
R302 B.n238 B.n57 163.367
R303 B.n239 B.n238 163.367
R304 B.n240 B.n239 163.367
R305 B.n240 B.n55 163.367
R306 B.n244 B.n55 163.367
R307 B.n245 B.n244 163.367
R308 B.n246 B.n245 163.367
R309 B.n246 B.n53 163.367
R310 B.n250 B.n53 163.367
R311 B.n251 B.n250 163.367
R312 B.n252 B.n251 163.367
R313 B.n252 B.n51 163.367
R314 B.n256 B.n51 163.367
R315 B.n257 B.n256 163.367
R316 B.n258 B.n257 163.367
R317 B.n258 B.n49 163.367
R318 B.n262 B.n49 163.367
R319 B.n263 B.n262 163.367
R320 B.n264 B.n263 163.367
R321 B.n264 B.n47 163.367
R322 B.n268 B.n47 163.367
R323 B.n269 B.n268 163.367
R324 B.n270 B.n269 163.367
R325 B.n270 B.n45 163.367
R326 B.n274 B.n45 163.367
R327 B.n360 B.n11 163.367
R328 B.n360 B.n359 163.367
R329 B.n359 B.n358 163.367
R330 B.n358 B.n13 163.367
R331 B.n354 B.n13 163.367
R332 B.n354 B.n353 163.367
R333 B.n353 B.n352 163.367
R334 B.n352 B.n15 163.367
R335 B.n348 B.n15 163.367
R336 B.n348 B.n347 163.367
R337 B.n347 B.n346 163.367
R338 B.n346 B.n17 163.367
R339 B.n342 B.n17 163.367
R340 B.n342 B.n341 163.367
R341 B.n341 B.n340 163.367
R342 B.n340 B.n19 163.367
R343 B.n336 B.n19 163.367
R344 B.n336 B.n335 163.367
R345 B.n335 B.n334 163.367
R346 B.n334 B.n21 163.367
R347 B.n330 B.n21 163.367
R348 B.n330 B.n329 163.367
R349 B.n329 B.n328 163.367
R350 B.n328 B.n23 163.367
R351 B.n323 B.n23 163.367
R352 B.n323 B.n322 163.367
R353 B.n322 B.n321 163.367
R354 B.n321 B.n27 163.367
R355 B.n317 B.n27 163.367
R356 B.n317 B.n316 163.367
R357 B.n316 B.n315 163.367
R358 B.n315 B.n29 163.367
R359 B.n311 B.n29 163.367
R360 B.n311 B.n310 163.367
R361 B.n310 B.n33 163.367
R362 B.n306 B.n33 163.367
R363 B.n306 B.n305 163.367
R364 B.n305 B.n304 163.367
R365 B.n304 B.n35 163.367
R366 B.n300 B.n35 163.367
R367 B.n300 B.n299 163.367
R368 B.n299 B.n298 163.367
R369 B.n298 B.n37 163.367
R370 B.n294 B.n37 163.367
R371 B.n294 B.n293 163.367
R372 B.n293 B.n292 163.367
R373 B.n292 B.n39 163.367
R374 B.n288 B.n39 163.367
R375 B.n288 B.n287 163.367
R376 B.n287 B.n286 163.367
R377 B.n286 B.n41 163.367
R378 B.n282 B.n41 163.367
R379 B.n282 B.n281 163.367
R380 B.n281 B.n280 163.367
R381 B.n280 B.n43 163.367
R382 B.n276 B.n43 163.367
R383 B.n276 B.n275 163.367
R384 B.n76 B.t2 144.669
R385 B.n30 B.t10 144.669
R386 B.n82 B.t8 144.662
R387 B.n24 B.t4 144.662
R388 B.n77 B.t1 111.7
R389 B.n31 B.t11 111.7
R390 B.n83 B.t7 111.694
R391 B.n25 B.t5 111.694
R392 B.n182 B.n77 59.5399
R393 B.n84 B.n83 59.5399
R394 B.n326 B.n25 59.5399
R395 B.n32 B.n31 59.5399
R396 B.n363 B.n362 36.3712
R397 B.n219 B.n218 36.3712
R398 B.n129 B.n96 36.3712
R399 B.n273 B.n44 36.3712
R400 B.n77 B.n76 32.9702
R401 B.n83 B.n82 32.9702
R402 B.n25 B.n24 32.9702
R403 B.n31 B.n30 32.9702
R404 B B.n391 18.0485
R405 B.n362 B.n361 10.6151
R406 B.n361 B.n12 10.6151
R407 B.n357 B.n12 10.6151
R408 B.n357 B.n356 10.6151
R409 B.n356 B.n355 10.6151
R410 B.n355 B.n14 10.6151
R411 B.n351 B.n14 10.6151
R412 B.n351 B.n350 10.6151
R413 B.n350 B.n349 10.6151
R414 B.n349 B.n16 10.6151
R415 B.n345 B.n16 10.6151
R416 B.n345 B.n344 10.6151
R417 B.n344 B.n343 10.6151
R418 B.n343 B.n18 10.6151
R419 B.n339 B.n18 10.6151
R420 B.n339 B.n338 10.6151
R421 B.n338 B.n337 10.6151
R422 B.n337 B.n20 10.6151
R423 B.n333 B.n20 10.6151
R424 B.n333 B.n332 10.6151
R425 B.n332 B.n331 10.6151
R426 B.n331 B.n22 10.6151
R427 B.n327 B.n22 10.6151
R428 B.n325 B.n324 10.6151
R429 B.n324 B.n26 10.6151
R430 B.n320 B.n26 10.6151
R431 B.n320 B.n319 10.6151
R432 B.n319 B.n318 10.6151
R433 B.n318 B.n28 10.6151
R434 B.n314 B.n28 10.6151
R435 B.n314 B.n313 10.6151
R436 B.n313 B.n312 10.6151
R437 B.n309 B.n308 10.6151
R438 B.n308 B.n307 10.6151
R439 B.n307 B.n34 10.6151
R440 B.n303 B.n34 10.6151
R441 B.n303 B.n302 10.6151
R442 B.n302 B.n301 10.6151
R443 B.n301 B.n36 10.6151
R444 B.n297 B.n36 10.6151
R445 B.n297 B.n296 10.6151
R446 B.n296 B.n295 10.6151
R447 B.n295 B.n38 10.6151
R448 B.n291 B.n38 10.6151
R449 B.n291 B.n290 10.6151
R450 B.n290 B.n289 10.6151
R451 B.n289 B.n40 10.6151
R452 B.n285 B.n40 10.6151
R453 B.n285 B.n284 10.6151
R454 B.n284 B.n283 10.6151
R455 B.n283 B.n42 10.6151
R456 B.n279 B.n42 10.6151
R457 B.n279 B.n278 10.6151
R458 B.n278 B.n277 10.6151
R459 B.n277 B.n44 10.6151
R460 B.n219 B.n62 10.6151
R461 B.n223 B.n62 10.6151
R462 B.n224 B.n223 10.6151
R463 B.n225 B.n224 10.6151
R464 B.n225 B.n60 10.6151
R465 B.n229 B.n60 10.6151
R466 B.n230 B.n229 10.6151
R467 B.n231 B.n230 10.6151
R468 B.n231 B.n58 10.6151
R469 B.n235 B.n58 10.6151
R470 B.n236 B.n235 10.6151
R471 B.n237 B.n236 10.6151
R472 B.n237 B.n56 10.6151
R473 B.n241 B.n56 10.6151
R474 B.n242 B.n241 10.6151
R475 B.n243 B.n242 10.6151
R476 B.n243 B.n54 10.6151
R477 B.n247 B.n54 10.6151
R478 B.n248 B.n247 10.6151
R479 B.n249 B.n248 10.6151
R480 B.n249 B.n52 10.6151
R481 B.n253 B.n52 10.6151
R482 B.n254 B.n253 10.6151
R483 B.n255 B.n254 10.6151
R484 B.n255 B.n50 10.6151
R485 B.n259 B.n50 10.6151
R486 B.n260 B.n259 10.6151
R487 B.n261 B.n260 10.6151
R488 B.n261 B.n48 10.6151
R489 B.n265 B.n48 10.6151
R490 B.n266 B.n265 10.6151
R491 B.n267 B.n266 10.6151
R492 B.n267 B.n46 10.6151
R493 B.n271 B.n46 10.6151
R494 B.n272 B.n271 10.6151
R495 B.n273 B.n272 10.6151
R496 B.n133 B.n96 10.6151
R497 B.n134 B.n133 10.6151
R498 B.n135 B.n134 10.6151
R499 B.n135 B.n94 10.6151
R500 B.n139 B.n94 10.6151
R501 B.n140 B.n139 10.6151
R502 B.n141 B.n140 10.6151
R503 B.n141 B.n92 10.6151
R504 B.n145 B.n92 10.6151
R505 B.n146 B.n145 10.6151
R506 B.n147 B.n146 10.6151
R507 B.n147 B.n90 10.6151
R508 B.n151 B.n90 10.6151
R509 B.n152 B.n151 10.6151
R510 B.n153 B.n152 10.6151
R511 B.n153 B.n88 10.6151
R512 B.n157 B.n88 10.6151
R513 B.n158 B.n157 10.6151
R514 B.n159 B.n158 10.6151
R515 B.n159 B.n86 10.6151
R516 B.n163 B.n86 10.6151
R517 B.n164 B.n163 10.6151
R518 B.n165 B.n164 10.6151
R519 B.n169 B.n168 10.6151
R520 B.n170 B.n169 10.6151
R521 B.n170 B.n80 10.6151
R522 B.n174 B.n80 10.6151
R523 B.n175 B.n174 10.6151
R524 B.n176 B.n175 10.6151
R525 B.n176 B.n78 10.6151
R526 B.n180 B.n78 10.6151
R527 B.n181 B.n180 10.6151
R528 B.n183 B.n74 10.6151
R529 B.n187 B.n74 10.6151
R530 B.n188 B.n187 10.6151
R531 B.n189 B.n188 10.6151
R532 B.n189 B.n72 10.6151
R533 B.n193 B.n72 10.6151
R534 B.n194 B.n193 10.6151
R535 B.n195 B.n194 10.6151
R536 B.n195 B.n70 10.6151
R537 B.n199 B.n70 10.6151
R538 B.n200 B.n199 10.6151
R539 B.n201 B.n200 10.6151
R540 B.n201 B.n68 10.6151
R541 B.n205 B.n68 10.6151
R542 B.n206 B.n205 10.6151
R543 B.n207 B.n206 10.6151
R544 B.n207 B.n66 10.6151
R545 B.n211 B.n66 10.6151
R546 B.n212 B.n211 10.6151
R547 B.n213 B.n212 10.6151
R548 B.n213 B.n64 10.6151
R549 B.n217 B.n64 10.6151
R550 B.n218 B.n217 10.6151
R551 B.n129 B.n128 10.6151
R552 B.n128 B.n127 10.6151
R553 B.n127 B.n98 10.6151
R554 B.n123 B.n98 10.6151
R555 B.n123 B.n122 10.6151
R556 B.n122 B.n121 10.6151
R557 B.n121 B.n100 10.6151
R558 B.n117 B.n100 10.6151
R559 B.n117 B.n116 10.6151
R560 B.n116 B.n115 10.6151
R561 B.n115 B.n102 10.6151
R562 B.n111 B.n102 10.6151
R563 B.n111 B.n110 10.6151
R564 B.n110 B.n109 10.6151
R565 B.n109 B.n104 10.6151
R566 B.n105 B.n104 10.6151
R567 B.n105 B.n0 10.6151
R568 B.n387 B.n1 10.6151
R569 B.n387 B.n386 10.6151
R570 B.n386 B.n385 10.6151
R571 B.n385 B.n4 10.6151
R572 B.n381 B.n4 10.6151
R573 B.n381 B.n380 10.6151
R574 B.n380 B.n379 10.6151
R575 B.n379 B.n6 10.6151
R576 B.n375 B.n6 10.6151
R577 B.n375 B.n374 10.6151
R578 B.n374 B.n373 10.6151
R579 B.n373 B.n8 10.6151
R580 B.n369 B.n8 10.6151
R581 B.n369 B.n368 10.6151
R582 B.n368 B.n367 10.6151
R583 B.n367 B.n10 10.6151
R584 B.n363 B.n10 10.6151
R585 B.n327 B.n326 9.36635
R586 B.n309 B.n32 9.36635
R587 B.n165 B.n84 9.36635
R588 B.n183 B.n182 9.36635
R589 B.n391 B.n0 2.81026
R590 B.n391 B.n1 2.81026
R591 B.n326 B.n325 1.24928
R592 B.n312 B.n32 1.24928
R593 B.n168 B.n84 1.24928
R594 B.n182 B.n181 1.24928
R595 VN VN.t1 255.255
R596 VN VN.t0 218.137
R597 VTAIL.n1 VTAIL.t2 81.5112
R598 VTAIL.n3 VTAIL.t3 81.5103
R599 VTAIL.n0 VTAIL.t1 81.5103
R600 VTAIL.n2 VTAIL.t0 81.5102
R601 VTAIL.n1 VTAIL.n0 20.6169
R602 VTAIL.n3 VTAIL.n2 19.1514
R603 VTAIL.n2 VTAIL.n1 1.20309
R604 VTAIL VTAIL.n0 0.894897
R605 VTAIL VTAIL.n3 0.30869
R606 VDD2.n0 VDD2.t1 130.099
R607 VDD2.n0 VDD2.t0 98.189
R608 VDD2 VDD2.n0 0.425069
R609 VP.n0 VP.t1 254.97
R610 VP.n0 VP.t0 217.992
R611 VP VP.n0 0.146778
R612 VDD1 VDD1.t1 130.989
R613 VDD1 VDD1.t0 98.6136
C0 VN w_n1650_n2202# 2.05891f
C1 VTAIL w_n1650_n2202# 1.90899f
C2 VDD1 VP 1.50764f
C3 VN B 0.77105f
C4 VN VDD2 1.37624f
C5 VTAIL B 1.92161f
C6 VTAIL VDD2 3.37516f
C7 VP w_n1650_n2202# 2.26644f
C8 VP B 1.1073f
C9 VDD2 VP 0.280872f
C10 VDD1 w_n1650_n2202# 1.22551f
C11 VTAIL VN 1.2628f
C12 VDD1 B 1.08646f
C13 VDD1 VDD2 0.53062f
C14 VN VP 3.79839f
C15 VTAIL VP 1.27707f
C16 B w_n1650_n2202# 5.84926f
C17 VDD2 w_n1650_n2202# 1.23693f
C18 VDD1 VN 0.147558f
C19 VDD2 B 1.10588f
C20 VDD1 VTAIL 3.33248f
C21 VDD2 VSUBS 0.579327f
C22 VDD1 VSUBS 2.533275f
C23 VTAIL VSUBS 0.464514f
C24 VN VSUBS 4.89168f
C25 VP VSUBS 1.023637f
C26 B VSUBS 2.491012f
C27 w_n1650_n2202# VSUBS 45.322197f
C28 VDD1.t0 VSUBS 0.629086f
C29 VDD1.t1 VSUBS 0.844339f
C30 VP.t1 VSUBS 1.50456f
C31 VP.t0 VSUBS 1.246f
C32 VP.n0 VSUBS 3.30764f
C33 VDD2.t1 VSUBS 0.869371f
C34 VDD2.t0 VSUBS 0.657335f
C35 VDD2.n0 VSUBS 1.81758f
C36 VTAIL.t1 VSUBS 0.664714f
C37 VTAIL.n0 VSUBS 1.03263f
C38 VTAIL.t2 VSUBS 0.664716f
C39 VTAIL.n1 VSUBS 1.04885f
C40 VTAIL.t0 VSUBS 0.664712f
C41 VTAIL.n2 VSUBS 0.971726f
C42 VTAIL.t3 VSUBS 0.664714f
C43 VTAIL.n3 VSUBS 0.924654f
C44 VN.t0 VSUBS 1.19338f
C45 VN.t1 VSUBS 1.44587f
C46 B.n0 VSUBS 0.003887f
C47 B.n1 VSUBS 0.003887f
C48 B.n2 VSUBS 0.006147f
C49 B.n3 VSUBS 0.006147f
C50 B.n4 VSUBS 0.006147f
C51 B.n5 VSUBS 0.006147f
C52 B.n6 VSUBS 0.006147f
C53 B.n7 VSUBS 0.006147f
C54 B.n8 VSUBS 0.006147f
C55 B.n9 VSUBS 0.006147f
C56 B.n10 VSUBS 0.006147f
C57 B.n11 VSUBS 0.015688f
C58 B.n12 VSUBS 0.006147f
C59 B.n13 VSUBS 0.006147f
C60 B.n14 VSUBS 0.006147f
C61 B.n15 VSUBS 0.006147f
C62 B.n16 VSUBS 0.006147f
C63 B.n17 VSUBS 0.006147f
C64 B.n18 VSUBS 0.006147f
C65 B.n19 VSUBS 0.006147f
C66 B.n20 VSUBS 0.006147f
C67 B.n21 VSUBS 0.006147f
C68 B.n22 VSUBS 0.006147f
C69 B.n23 VSUBS 0.006147f
C70 B.t5 VSUBS 0.159165f
C71 B.t4 VSUBS 0.17032f
C72 B.t3 VSUBS 0.337414f
C73 B.n24 VSUBS 0.090275f
C74 B.n25 VSUBS 0.057711f
C75 B.n26 VSUBS 0.006147f
C76 B.n27 VSUBS 0.006147f
C77 B.n28 VSUBS 0.006147f
C78 B.n29 VSUBS 0.006147f
C79 B.t11 VSUBS 0.159165f
C80 B.t10 VSUBS 0.170319f
C81 B.t9 VSUBS 0.337414f
C82 B.n30 VSUBS 0.090276f
C83 B.n31 VSUBS 0.057712f
C84 B.n32 VSUBS 0.014241f
C85 B.n33 VSUBS 0.006147f
C86 B.n34 VSUBS 0.006147f
C87 B.n35 VSUBS 0.006147f
C88 B.n36 VSUBS 0.006147f
C89 B.n37 VSUBS 0.006147f
C90 B.n38 VSUBS 0.006147f
C91 B.n39 VSUBS 0.006147f
C92 B.n40 VSUBS 0.006147f
C93 B.n41 VSUBS 0.006147f
C94 B.n42 VSUBS 0.006147f
C95 B.n43 VSUBS 0.006147f
C96 B.n44 VSUBS 0.015036f
C97 B.n45 VSUBS 0.006147f
C98 B.n46 VSUBS 0.006147f
C99 B.n47 VSUBS 0.006147f
C100 B.n48 VSUBS 0.006147f
C101 B.n49 VSUBS 0.006147f
C102 B.n50 VSUBS 0.006147f
C103 B.n51 VSUBS 0.006147f
C104 B.n52 VSUBS 0.006147f
C105 B.n53 VSUBS 0.006147f
C106 B.n54 VSUBS 0.006147f
C107 B.n55 VSUBS 0.006147f
C108 B.n56 VSUBS 0.006147f
C109 B.n57 VSUBS 0.006147f
C110 B.n58 VSUBS 0.006147f
C111 B.n59 VSUBS 0.006147f
C112 B.n60 VSUBS 0.006147f
C113 B.n61 VSUBS 0.006147f
C114 B.n62 VSUBS 0.006147f
C115 B.n63 VSUBS 0.015688f
C116 B.n64 VSUBS 0.006147f
C117 B.n65 VSUBS 0.006147f
C118 B.n66 VSUBS 0.006147f
C119 B.n67 VSUBS 0.006147f
C120 B.n68 VSUBS 0.006147f
C121 B.n69 VSUBS 0.006147f
C122 B.n70 VSUBS 0.006147f
C123 B.n71 VSUBS 0.006147f
C124 B.n72 VSUBS 0.006147f
C125 B.n73 VSUBS 0.006147f
C126 B.n74 VSUBS 0.006147f
C127 B.n75 VSUBS 0.006147f
C128 B.t1 VSUBS 0.159165f
C129 B.t2 VSUBS 0.170319f
C130 B.t0 VSUBS 0.337414f
C131 B.n76 VSUBS 0.090276f
C132 B.n77 VSUBS 0.057712f
C133 B.n78 VSUBS 0.006147f
C134 B.n79 VSUBS 0.006147f
C135 B.n80 VSUBS 0.006147f
C136 B.n81 VSUBS 0.006147f
C137 B.t7 VSUBS 0.159165f
C138 B.t8 VSUBS 0.17032f
C139 B.t6 VSUBS 0.337414f
C140 B.n82 VSUBS 0.090275f
C141 B.n83 VSUBS 0.057711f
C142 B.n84 VSUBS 0.014241f
C143 B.n85 VSUBS 0.006147f
C144 B.n86 VSUBS 0.006147f
C145 B.n87 VSUBS 0.006147f
C146 B.n88 VSUBS 0.006147f
C147 B.n89 VSUBS 0.006147f
C148 B.n90 VSUBS 0.006147f
C149 B.n91 VSUBS 0.006147f
C150 B.n92 VSUBS 0.006147f
C151 B.n93 VSUBS 0.006147f
C152 B.n94 VSUBS 0.006147f
C153 B.n95 VSUBS 0.006147f
C154 B.n96 VSUBS 0.015688f
C155 B.n97 VSUBS 0.006147f
C156 B.n98 VSUBS 0.006147f
C157 B.n99 VSUBS 0.006147f
C158 B.n100 VSUBS 0.006147f
C159 B.n101 VSUBS 0.006147f
C160 B.n102 VSUBS 0.006147f
C161 B.n103 VSUBS 0.006147f
C162 B.n104 VSUBS 0.006147f
C163 B.n105 VSUBS 0.006147f
C164 B.n106 VSUBS 0.006147f
C165 B.n107 VSUBS 0.006147f
C166 B.n108 VSUBS 0.006147f
C167 B.n109 VSUBS 0.006147f
C168 B.n110 VSUBS 0.006147f
C169 B.n111 VSUBS 0.006147f
C170 B.n112 VSUBS 0.006147f
C171 B.n113 VSUBS 0.006147f
C172 B.n114 VSUBS 0.006147f
C173 B.n115 VSUBS 0.006147f
C174 B.n116 VSUBS 0.006147f
C175 B.n117 VSUBS 0.006147f
C176 B.n118 VSUBS 0.006147f
C177 B.n119 VSUBS 0.006147f
C178 B.n120 VSUBS 0.006147f
C179 B.n121 VSUBS 0.006147f
C180 B.n122 VSUBS 0.006147f
C181 B.n123 VSUBS 0.006147f
C182 B.n124 VSUBS 0.006147f
C183 B.n125 VSUBS 0.006147f
C184 B.n126 VSUBS 0.006147f
C185 B.n127 VSUBS 0.006147f
C186 B.n128 VSUBS 0.006147f
C187 B.n129 VSUBS 0.015227f
C188 B.n130 VSUBS 0.015227f
C189 B.n131 VSUBS 0.015688f
C190 B.n132 VSUBS 0.006147f
C191 B.n133 VSUBS 0.006147f
C192 B.n134 VSUBS 0.006147f
C193 B.n135 VSUBS 0.006147f
C194 B.n136 VSUBS 0.006147f
C195 B.n137 VSUBS 0.006147f
C196 B.n138 VSUBS 0.006147f
C197 B.n139 VSUBS 0.006147f
C198 B.n140 VSUBS 0.006147f
C199 B.n141 VSUBS 0.006147f
C200 B.n142 VSUBS 0.006147f
C201 B.n143 VSUBS 0.006147f
C202 B.n144 VSUBS 0.006147f
C203 B.n145 VSUBS 0.006147f
C204 B.n146 VSUBS 0.006147f
C205 B.n147 VSUBS 0.006147f
C206 B.n148 VSUBS 0.006147f
C207 B.n149 VSUBS 0.006147f
C208 B.n150 VSUBS 0.006147f
C209 B.n151 VSUBS 0.006147f
C210 B.n152 VSUBS 0.006147f
C211 B.n153 VSUBS 0.006147f
C212 B.n154 VSUBS 0.006147f
C213 B.n155 VSUBS 0.006147f
C214 B.n156 VSUBS 0.006147f
C215 B.n157 VSUBS 0.006147f
C216 B.n158 VSUBS 0.006147f
C217 B.n159 VSUBS 0.006147f
C218 B.n160 VSUBS 0.006147f
C219 B.n161 VSUBS 0.006147f
C220 B.n162 VSUBS 0.006147f
C221 B.n163 VSUBS 0.006147f
C222 B.n164 VSUBS 0.006147f
C223 B.n165 VSUBS 0.005785f
C224 B.n166 VSUBS 0.006147f
C225 B.n167 VSUBS 0.006147f
C226 B.n168 VSUBS 0.003435f
C227 B.n169 VSUBS 0.006147f
C228 B.n170 VSUBS 0.006147f
C229 B.n171 VSUBS 0.006147f
C230 B.n172 VSUBS 0.006147f
C231 B.n173 VSUBS 0.006147f
C232 B.n174 VSUBS 0.006147f
C233 B.n175 VSUBS 0.006147f
C234 B.n176 VSUBS 0.006147f
C235 B.n177 VSUBS 0.006147f
C236 B.n178 VSUBS 0.006147f
C237 B.n179 VSUBS 0.006147f
C238 B.n180 VSUBS 0.006147f
C239 B.n181 VSUBS 0.003435f
C240 B.n182 VSUBS 0.014241f
C241 B.n183 VSUBS 0.005785f
C242 B.n184 VSUBS 0.006147f
C243 B.n185 VSUBS 0.006147f
C244 B.n186 VSUBS 0.006147f
C245 B.n187 VSUBS 0.006147f
C246 B.n188 VSUBS 0.006147f
C247 B.n189 VSUBS 0.006147f
C248 B.n190 VSUBS 0.006147f
C249 B.n191 VSUBS 0.006147f
C250 B.n192 VSUBS 0.006147f
C251 B.n193 VSUBS 0.006147f
C252 B.n194 VSUBS 0.006147f
C253 B.n195 VSUBS 0.006147f
C254 B.n196 VSUBS 0.006147f
C255 B.n197 VSUBS 0.006147f
C256 B.n198 VSUBS 0.006147f
C257 B.n199 VSUBS 0.006147f
C258 B.n200 VSUBS 0.006147f
C259 B.n201 VSUBS 0.006147f
C260 B.n202 VSUBS 0.006147f
C261 B.n203 VSUBS 0.006147f
C262 B.n204 VSUBS 0.006147f
C263 B.n205 VSUBS 0.006147f
C264 B.n206 VSUBS 0.006147f
C265 B.n207 VSUBS 0.006147f
C266 B.n208 VSUBS 0.006147f
C267 B.n209 VSUBS 0.006147f
C268 B.n210 VSUBS 0.006147f
C269 B.n211 VSUBS 0.006147f
C270 B.n212 VSUBS 0.006147f
C271 B.n213 VSUBS 0.006147f
C272 B.n214 VSUBS 0.006147f
C273 B.n215 VSUBS 0.006147f
C274 B.n216 VSUBS 0.006147f
C275 B.n217 VSUBS 0.006147f
C276 B.n218 VSUBS 0.015688f
C277 B.n219 VSUBS 0.015227f
C278 B.n220 VSUBS 0.015227f
C279 B.n221 VSUBS 0.006147f
C280 B.n222 VSUBS 0.006147f
C281 B.n223 VSUBS 0.006147f
C282 B.n224 VSUBS 0.006147f
C283 B.n225 VSUBS 0.006147f
C284 B.n226 VSUBS 0.006147f
C285 B.n227 VSUBS 0.006147f
C286 B.n228 VSUBS 0.006147f
C287 B.n229 VSUBS 0.006147f
C288 B.n230 VSUBS 0.006147f
C289 B.n231 VSUBS 0.006147f
C290 B.n232 VSUBS 0.006147f
C291 B.n233 VSUBS 0.006147f
C292 B.n234 VSUBS 0.006147f
C293 B.n235 VSUBS 0.006147f
C294 B.n236 VSUBS 0.006147f
C295 B.n237 VSUBS 0.006147f
C296 B.n238 VSUBS 0.006147f
C297 B.n239 VSUBS 0.006147f
C298 B.n240 VSUBS 0.006147f
C299 B.n241 VSUBS 0.006147f
C300 B.n242 VSUBS 0.006147f
C301 B.n243 VSUBS 0.006147f
C302 B.n244 VSUBS 0.006147f
C303 B.n245 VSUBS 0.006147f
C304 B.n246 VSUBS 0.006147f
C305 B.n247 VSUBS 0.006147f
C306 B.n248 VSUBS 0.006147f
C307 B.n249 VSUBS 0.006147f
C308 B.n250 VSUBS 0.006147f
C309 B.n251 VSUBS 0.006147f
C310 B.n252 VSUBS 0.006147f
C311 B.n253 VSUBS 0.006147f
C312 B.n254 VSUBS 0.006147f
C313 B.n255 VSUBS 0.006147f
C314 B.n256 VSUBS 0.006147f
C315 B.n257 VSUBS 0.006147f
C316 B.n258 VSUBS 0.006147f
C317 B.n259 VSUBS 0.006147f
C318 B.n260 VSUBS 0.006147f
C319 B.n261 VSUBS 0.006147f
C320 B.n262 VSUBS 0.006147f
C321 B.n263 VSUBS 0.006147f
C322 B.n264 VSUBS 0.006147f
C323 B.n265 VSUBS 0.006147f
C324 B.n266 VSUBS 0.006147f
C325 B.n267 VSUBS 0.006147f
C326 B.n268 VSUBS 0.006147f
C327 B.n269 VSUBS 0.006147f
C328 B.n270 VSUBS 0.006147f
C329 B.n271 VSUBS 0.006147f
C330 B.n272 VSUBS 0.006147f
C331 B.n273 VSUBS 0.015879f
C332 B.n274 VSUBS 0.015227f
C333 B.n275 VSUBS 0.015688f
C334 B.n276 VSUBS 0.006147f
C335 B.n277 VSUBS 0.006147f
C336 B.n278 VSUBS 0.006147f
C337 B.n279 VSUBS 0.006147f
C338 B.n280 VSUBS 0.006147f
C339 B.n281 VSUBS 0.006147f
C340 B.n282 VSUBS 0.006147f
C341 B.n283 VSUBS 0.006147f
C342 B.n284 VSUBS 0.006147f
C343 B.n285 VSUBS 0.006147f
C344 B.n286 VSUBS 0.006147f
C345 B.n287 VSUBS 0.006147f
C346 B.n288 VSUBS 0.006147f
C347 B.n289 VSUBS 0.006147f
C348 B.n290 VSUBS 0.006147f
C349 B.n291 VSUBS 0.006147f
C350 B.n292 VSUBS 0.006147f
C351 B.n293 VSUBS 0.006147f
C352 B.n294 VSUBS 0.006147f
C353 B.n295 VSUBS 0.006147f
C354 B.n296 VSUBS 0.006147f
C355 B.n297 VSUBS 0.006147f
C356 B.n298 VSUBS 0.006147f
C357 B.n299 VSUBS 0.006147f
C358 B.n300 VSUBS 0.006147f
C359 B.n301 VSUBS 0.006147f
C360 B.n302 VSUBS 0.006147f
C361 B.n303 VSUBS 0.006147f
C362 B.n304 VSUBS 0.006147f
C363 B.n305 VSUBS 0.006147f
C364 B.n306 VSUBS 0.006147f
C365 B.n307 VSUBS 0.006147f
C366 B.n308 VSUBS 0.006147f
C367 B.n309 VSUBS 0.005785f
C368 B.n310 VSUBS 0.006147f
C369 B.n311 VSUBS 0.006147f
C370 B.n312 VSUBS 0.003435f
C371 B.n313 VSUBS 0.006147f
C372 B.n314 VSUBS 0.006147f
C373 B.n315 VSUBS 0.006147f
C374 B.n316 VSUBS 0.006147f
C375 B.n317 VSUBS 0.006147f
C376 B.n318 VSUBS 0.006147f
C377 B.n319 VSUBS 0.006147f
C378 B.n320 VSUBS 0.006147f
C379 B.n321 VSUBS 0.006147f
C380 B.n322 VSUBS 0.006147f
C381 B.n323 VSUBS 0.006147f
C382 B.n324 VSUBS 0.006147f
C383 B.n325 VSUBS 0.003435f
C384 B.n326 VSUBS 0.014241f
C385 B.n327 VSUBS 0.005785f
C386 B.n328 VSUBS 0.006147f
C387 B.n329 VSUBS 0.006147f
C388 B.n330 VSUBS 0.006147f
C389 B.n331 VSUBS 0.006147f
C390 B.n332 VSUBS 0.006147f
C391 B.n333 VSUBS 0.006147f
C392 B.n334 VSUBS 0.006147f
C393 B.n335 VSUBS 0.006147f
C394 B.n336 VSUBS 0.006147f
C395 B.n337 VSUBS 0.006147f
C396 B.n338 VSUBS 0.006147f
C397 B.n339 VSUBS 0.006147f
C398 B.n340 VSUBS 0.006147f
C399 B.n341 VSUBS 0.006147f
C400 B.n342 VSUBS 0.006147f
C401 B.n343 VSUBS 0.006147f
C402 B.n344 VSUBS 0.006147f
C403 B.n345 VSUBS 0.006147f
C404 B.n346 VSUBS 0.006147f
C405 B.n347 VSUBS 0.006147f
C406 B.n348 VSUBS 0.006147f
C407 B.n349 VSUBS 0.006147f
C408 B.n350 VSUBS 0.006147f
C409 B.n351 VSUBS 0.006147f
C410 B.n352 VSUBS 0.006147f
C411 B.n353 VSUBS 0.006147f
C412 B.n354 VSUBS 0.006147f
C413 B.n355 VSUBS 0.006147f
C414 B.n356 VSUBS 0.006147f
C415 B.n357 VSUBS 0.006147f
C416 B.n358 VSUBS 0.006147f
C417 B.n359 VSUBS 0.006147f
C418 B.n360 VSUBS 0.006147f
C419 B.n361 VSUBS 0.006147f
C420 B.n362 VSUBS 0.015688f
C421 B.n363 VSUBS 0.015227f
C422 B.n364 VSUBS 0.015227f
C423 B.n365 VSUBS 0.006147f
C424 B.n366 VSUBS 0.006147f
C425 B.n367 VSUBS 0.006147f
C426 B.n368 VSUBS 0.006147f
C427 B.n369 VSUBS 0.006147f
C428 B.n370 VSUBS 0.006147f
C429 B.n371 VSUBS 0.006147f
C430 B.n372 VSUBS 0.006147f
C431 B.n373 VSUBS 0.006147f
C432 B.n374 VSUBS 0.006147f
C433 B.n375 VSUBS 0.006147f
C434 B.n376 VSUBS 0.006147f
C435 B.n377 VSUBS 0.006147f
C436 B.n378 VSUBS 0.006147f
C437 B.n379 VSUBS 0.006147f
C438 B.n380 VSUBS 0.006147f
C439 B.n381 VSUBS 0.006147f
C440 B.n382 VSUBS 0.006147f
C441 B.n383 VSUBS 0.006147f
C442 B.n384 VSUBS 0.006147f
C443 B.n385 VSUBS 0.006147f
C444 B.n386 VSUBS 0.006147f
C445 B.n387 VSUBS 0.006147f
C446 B.n388 VSUBS 0.006147f
C447 B.n389 VSUBS 0.006147f
C448 B.n390 VSUBS 0.006147f
C449 B.n391 VSUBS 0.013919f
.ends

