* NGSPICE file created from diff_pair_sample_1504.ext - technology: sky130A

.subckt diff_pair_sample_1504 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t7 w_n2922_n3092# sky130_fd_pr__pfet_01v8 ad=1.7523 pd=10.95 as=4.1418 ps=22.02 w=10.62 l=2.11
X1 VDD2.t4 VN.t1 VTAIL.t6 w_n2922_n3092# sky130_fd_pr__pfet_01v8 ad=4.1418 pd=22.02 as=1.7523 ps=10.95 w=10.62 l=2.11
X2 VDD1.t5 VP.t0 VTAIL.t5 w_n2922_n3092# sky130_fd_pr__pfet_01v8 ad=4.1418 pd=22.02 as=1.7523 ps=10.95 w=10.62 l=2.11
X3 VTAIL.t0 VP.t1 VDD1.t4 w_n2922_n3092# sky130_fd_pr__pfet_01v8 ad=1.7523 pd=10.95 as=1.7523 ps=10.95 w=10.62 l=2.11
X4 B.t11 B.t9 B.t10 w_n2922_n3092# sky130_fd_pr__pfet_01v8 ad=4.1418 pd=22.02 as=0 ps=0 w=10.62 l=2.11
X5 VDD2.t3 VN.t2 VTAIL.t11 w_n2922_n3092# sky130_fd_pr__pfet_01v8 ad=4.1418 pd=22.02 as=1.7523 ps=10.95 w=10.62 l=2.11
X6 VDD1.t3 VP.t2 VTAIL.t3 w_n2922_n3092# sky130_fd_pr__pfet_01v8 ad=1.7523 pd=10.95 as=4.1418 ps=22.02 w=10.62 l=2.11
X7 B.t8 B.t6 B.t7 w_n2922_n3092# sky130_fd_pr__pfet_01v8 ad=4.1418 pd=22.02 as=0 ps=0 w=10.62 l=2.11
X8 VDD2.t2 VN.t3 VTAIL.t8 w_n2922_n3092# sky130_fd_pr__pfet_01v8 ad=1.7523 pd=10.95 as=4.1418 ps=22.02 w=10.62 l=2.11
X9 B.t5 B.t3 B.t4 w_n2922_n3092# sky130_fd_pr__pfet_01v8 ad=4.1418 pd=22.02 as=0 ps=0 w=10.62 l=2.11
X10 B.t2 B.t0 B.t1 w_n2922_n3092# sky130_fd_pr__pfet_01v8 ad=4.1418 pd=22.02 as=0 ps=0 w=10.62 l=2.11
X11 VTAIL.t10 VN.t4 VDD2.t1 w_n2922_n3092# sky130_fd_pr__pfet_01v8 ad=1.7523 pd=10.95 as=1.7523 ps=10.95 w=10.62 l=2.11
X12 VDD1.t2 VP.t3 VTAIL.t1 w_n2922_n3092# sky130_fd_pr__pfet_01v8 ad=1.7523 pd=10.95 as=4.1418 ps=22.02 w=10.62 l=2.11
X13 VTAIL.t2 VP.t4 VDD1.t1 w_n2922_n3092# sky130_fd_pr__pfet_01v8 ad=1.7523 pd=10.95 as=1.7523 ps=10.95 w=10.62 l=2.11
X14 VTAIL.t9 VN.t5 VDD2.t0 w_n2922_n3092# sky130_fd_pr__pfet_01v8 ad=1.7523 pd=10.95 as=1.7523 ps=10.95 w=10.62 l=2.11
X15 VDD1.t0 VP.t5 VTAIL.t4 w_n2922_n3092# sky130_fd_pr__pfet_01v8 ad=4.1418 pd=22.02 as=1.7523 ps=10.95 w=10.62 l=2.11
R0 VN.n21 VN.n12 161.3
R1 VN.n20 VN.n19 161.3
R2 VN.n18 VN.n13 161.3
R3 VN.n17 VN.n16 161.3
R4 VN.n9 VN.n0 161.3
R5 VN.n8 VN.n7 161.3
R6 VN.n6 VN.n1 161.3
R7 VN.n5 VN.n4 161.3
R8 VN.n2 VN.t1 155.772
R9 VN.n14 VN.t3 155.772
R10 VN.n3 VN.t4 121.3
R11 VN.n10 VN.t0 121.3
R12 VN.n15 VN.t5 121.3
R13 VN.n22 VN.t2 121.3
R14 VN.n11 VN.n10 89.2674
R15 VN.n23 VN.n22 89.2674
R16 VN.n8 VN.n1 56.5617
R17 VN.n20 VN.n13 56.5617
R18 VN.n15 VN.n14 46.3186
R19 VN.n3 VN.n2 46.3186
R20 VN VN.n23 46.0664
R21 VN.n4 VN.n3 24.5923
R22 VN.n4 VN.n1 24.5923
R23 VN.n9 VN.n8 24.5923
R24 VN.n16 VN.n13 24.5923
R25 VN.n16 VN.n15 24.5923
R26 VN.n21 VN.n20 24.5923
R27 VN.n10 VN.n9 21.6413
R28 VN.n22 VN.n21 21.6413
R29 VN.n17 VN.n14 8.80512
R30 VN.n5 VN.n2 8.80512
R31 VN.n23 VN.n12 0.278335
R32 VN.n11 VN.n0 0.278335
R33 VN.n19 VN.n12 0.189894
R34 VN.n19 VN.n18 0.189894
R35 VN.n18 VN.n17 0.189894
R36 VN.n6 VN.n5 0.189894
R37 VN.n7 VN.n6 0.189894
R38 VN.n7 VN.n0 0.189894
R39 VN VN.n11 0.153485
R40 VTAIL.n234 VTAIL.n182 756.745
R41 VTAIL.n54 VTAIL.n2 756.745
R42 VTAIL.n176 VTAIL.n124 756.745
R43 VTAIL.n116 VTAIL.n64 756.745
R44 VTAIL.n201 VTAIL.n200 585
R45 VTAIL.n198 VTAIL.n197 585
R46 VTAIL.n207 VTAIL.n206 585
R47 VTAIL.n209 VTAIL.n208 585
R48 VTAIL.n194 VTAIL.n193 585
R49 VTAIL.n215 VTAIL.n214 585
R50 VTAIL.n218 VTAIL.n217 585
R51 VTAIL.n216 VTAIL.n190 585
R52 VTAIL.n223 VTAIL.n189 585
R53 VTAIL.n225 VTAIL.n224 585
R54 VTAIL.n227 VTAIL.n226 585
R55 VTAIL.n186 VTAIL.n185 585
R56 VTAIL.n233 VTAIL.n232 585
R57 VTAIL.n235 VTAIL.n234 585
R58 VTAIL.n21 VTAIL.n20 585
R59 VTAIL.n18 VTAIL.n17 585
R60 VTAIL.n27 VTAIL.n26 585
R61 VTAIL.n29 VTAIL.n28 585
R62 VTAIL.n14 VTAIL.n13 585
R63 VTAIL.n35 VTAIL.n34 585
R64 VTAIL.n38 VTAIL.n37 585
R65 VTAIL.n36 VTAIL.n10 585
R66 VTAIL.n43 VTAIL.n9 585
R67 VTAIL.n45 VTAIL.n44 585
R68 VTAIL.n47 VTAIL.n46 585
R69 VTAIL.n6 VTAIL.n5 585
R70 VTAIL.n53 VTAIL.n52 585
R71 VTAIL.n55 VTAIL.n54 585
R72 VTAIL.n177 VTAIL.n176 585
R73 VTAIL.n175 VTAIL.n174 585
R74 VTAIL.n128 VTAIL.n127 585
R75 VTAIL.n169 VTAIL.n168 585
R76 VTAIL.n167 VTAIL.n166 585
R77 VTAIL.n165 VTAIL.n131 585
R78 VTAIL.n135 VTAIL.n132 585
R79 VTAIL.n160 VTAIL.n159 585
R80 VTAIL.n158 VTAIL.n157 585
R81 VTAIL.n137 VTAIL.n136 585
R82 VTAIL.n152 VTAIL.n151 585
R83 VTAIL.n150 VTAIL.n149 585
R84 VTAIL.n141 VTAIL.n140 585
R85 VTAIL.n144 VTAIL.n143 585
R86 VTAIL.n117 VTAIL.n116 585
R87 VTAIL.n115 VTAIL.n114 585
R88 VTAIL.n68 VTAIL.n67 585
R89 VTAIL.n109 VTAIL.n108 585
R90 VTAIL.n107 VTAIL.n106 585
R91 VTAIL.n105 VTAIL.n71 585
R92 VTAIL.n75 VTAIL.n72 585
R93 VTAIL.n100 VTAIL.n99 585
R94 VTAIL.n98 VTAIL.n97 585
R95 VTAIL.n77 VTAIL.n76 585
R96 VTAIL.n92 VTAIL.n91 585
R97 VTAIL.n90 VTAIL.n89 585
R98 VTAIL.n81 VTAIL.n80 585
R99 VTAIL.n84 VTAIL.n83 585
R100 VTAIL.t1 VTAIL.n142 329.038
R101 VTAIL.t8 VTAIL.n82 329.038
R102 VTAIL.t7 VTAIL.n199 329.038
R103 VTAIL.t3 VTAIL.n19 329.038
R104 VTAIL.n200 VTAIL.n197 171.744
R105 VTAIL.n207 VTAIL.n197 171.744
R106 VTAIL.n208 VTAIL.n207 171.744
R107 VTAIL.n208 VTAIL.n193 171.744
R108 VTAIL.n215 VTAIL.n193 171.744
R109 VTAIL.n217 VTAIL.n215 171.744
R110 VTAIL.n217 VTAIL.n216 171.744
R111 VTAIL.n216 VTAIL.n189 171.744
R112 VTAIL.n225 VTAIL.n189 171.744
R113 VTAIL.n226 VTAIL.n225 171.744
R114 VTAIL.n226 VTAIL.n185 171.744
R115 VTAIL.n233 VTAIL.n185 171.744
R116 VTAIL.n234 VTAIL.n233 171.744
R117 VTAIL.n20 VTAIL.n17 171.744
R118 VTAIL.n27 VTAIL.n17 171.744
R119 VTAIL.n28 VTAIL.n27 171.744
R120 VTAIL.n28 VTAIL.n13 171.744
R121 VTAIL.n35 VTAIL.n13 171.744
R122 VTAIL.n37 VTAIL.n35 171.744
R123 VTAIL.n37 VTAIL.n36 171.744
R124 VTAIL.n36 VTAIL.n9 171.744
R125 VTAIL.n45 VTAIL.n9 171.744
R126 VTAIL.n46 VTAIL.n45 171.744
R127 VTAIL.n46 VTAIL.n5 171.744
R128 VTAIL.n53 VTAIL.n5 171.744
R129 VTAIL.n54 VTAIL.n53 171.744
R130 VTAIL.n176 VTAIL.n175 171.744
R131 VTAIL.n175 VTAIL.n127 171.744
R132 VTAIL.n168 VTAIL.n127 171.744
R133 VTAIL.n168 VTAIL.n167 171.744
R134 VTAIL.n167 VTAIL.n131 171.744
R135 VTAIL.n135 VTAIL.n131 171.744
R136 VTAIL.n159 VTAIL.n135 171.744
R137 VTAIL.n159 VTAIL.n158 171.744
R138 VTAIL.n158 VTAIL.n136 171.744
R139 VTAIL.n151 VTAIL.n136 171.744
R140 VTAIL.n151 VTAIL.n150 171.744
R141 VTAIL.n150 VTAIL.n140 171.744
R142 VTAIL.n143 VTAIL.n140 171.744
R143 VTAIL.n116 VTAIL.n115 171.744
R144 VTAIL.n115 VTAIL.n67 171.744
R145 VTAIL.n108 VTAIL.n67 171.744
R146 VTAIL.n108 VTAIL.n107 171.744
R147 VTAIL.n107 VTAIL.n71 171.744
R148 VTAIL.n75 VTAIL.n71 171.744
R149 VTAIL.n99 VTAIL.n75 171.744
R150 VTAIL.n99 VTAIL.n98 171.744
R151 VTAIL.n98 VTAIL.n76 171.744
R152 VTAIL.n91 VTAIL.n76 171.744
R153 VTAIL.n91 VTAIL.n90 171.744
R154 VTAIL.n90 VTAIL.n80 171.744
R155 VTAIL.n83 VTAIL.n80 171.744
R156 VTAIL.n200 VTAIL.t7 85.8723
R157 VTAIL.n20 VTAIL.t3 85.8723
R158 VTAIL.n143 VTAIL.t1 85.8723
R159 VTAIL.n83 VTAIL.t8 85.8723
R160 VTAIL.n123 VTAIL.n122 58.0237
R161 VTAIL.n63 VTAIL.n62 58.0237
R162 VTAIL.n1 VTAIL.n0 58.0236
R163 VTAIL.n61 VTAIL.n60 58.0236
R164 VTAIL.n239 VTAIL.n238 31.0217
R165 VTAIL.n59 VTAIL.n58 31.0217
R166 VTAIL.n181 VTAIL.n180 31.0217
R167 VTAIL.n121 VTAIL.n120 31.0217
R168 VTAIL.n63 VTAIL.n61 25.7289
R169 VTAIL.n239 VTAIL.n181 23.6255
R170 VTAIL.n224 VTAIL.n223 13.1884
R171 VTAIL.n44 VTAIL.n43 13.1884
R172 VTAIL.n166 VTAIL.n165 13.1884
R173 VTAIL.n106 VTAIL.n105 13.1884
R174 VTAIL.n222 VTAIL.n190 12.8005
R175 VTAIL.n227 VTAIL.n188 12.8005
R176 VTAIL.n42 VTAIL.n10 12.8005
R177 VTAIL.n47 VTAIL.n8 12.8005
R178 VTAIL.n169 VTAIL.n130 12.8005
R179 VTAIL.n164 VTAIL.n132 12.8005
R180 VTAIL.n109 VTAIL.n70 12.8005
R181 VTAIL.n104 VTAIL.n72 12.8005
R182 VTAIL.n219 VTAIL.n218 12.0247
R183 VTAIL.n228 VTAIL.n186 12.0247
R184 VTAIL.n39 VTAIL.n38 12.0247
R185 VTAIL.n48 VTAIL.n6 12.0247
R186 VTAIL.n170 VTAIL.n128 12.0247
R187 VTAIL.n161 VTAIL.n160 12.0247
R188 VTAIL.n110 VTAIL.n68 12.0247
R189 VTAIL.n101 VTAIL.n100 12.0247
R190 VTAIL.n214 VTAIL.n192 11.249
R191 VTAIL.n232 VTAIL.n231 11.249
R192 VTAIL.n34 VTAIL.n12 11.249
R193 VTAIL.n52 VTAIL.n51 11.249
R194 VTAIL.n174 VTAIL.n173 11.249
R195 VTAIL.n157 VTAIL.n134 11.249
R196 VTAIL.n114 VTAIL.n113 11.249
R197 VTAIL.n97 VTAIL.n74 11.249
R198 VTAIL.n201 VTAIL.n199 10.7239
R199 VTAIL.n21 VTAIL.n19 10.7239
R200 VTAIL.n144 VTAIL.n142 10.7239
R201 VTAIL.n84 VTAIL.n82 10.7239
R202 VTAIL.n213 VTAIL.n194 10.4732
R203 VTAIL.n235 VTAIL.n184 10.4732
R204 VTAIL.n33 VTAIL.n14 10.4732
R205 VTAIL.n55 VTAIL.n4 10.4732
R206 VTAIL.n177 VTAIL.n126 10.4732
R207 VTAIL.n156 VTAIL.n137 10.4732
R208 VTAIL.n117 VTAIL.n66 10.4732
R209 VTAIL.n96 VTAIL.n77 10.4732
R210 VTAIL.n210 VTAIL.n209 9.69747
R211 VTAIL.n236 VTAIL.n182 9.69747
R212 VTAIL.n30 VTAIL.n29 9.69747
R213 VTAIL.n56 VTAIL.n2 9.69747
R214 VTAIL.n178 VTAIL.n124 9.69747
R215 VTAIL.n153 VTAIL.n152 9.69747
R216 VTAIL.n118 VTAIL.n64 9.69747
R217 VTAIL.n93 VTAIL.n92 9.69747
R218 VTAIL.n238 VTAIL.n237 9.45567
R219 VTAIL.n58 VTAIL.n57 9.45567
R220 VTAIL.n180 VTAIL.n179 9.45567
R221 VTAIL.n120 VTAIL.n119 9.45567
R222 VTAIL.n237 VTAIL.n236 9.3005
R223 VTAIL.n184 VTAIL.n183 9.3005
R224 VTAIL.n231 VTAIL.n230 9.3005
R225 VTAIL.n229 VTAIL.n228 9.3005
R226 VTAIL.n188 VTAIL.n187 9.3005
R227 VTAIL.n203 VTAIL.n202 9.3005
R228 VTAIL.n205 VTAIL.n204 9.3005
R229 VTAIL.n196 VTAIL.n195 9.3005
R230 VTAIL.n211 VTAIL.n210 9.3005
R231 VTAIL.n213 VTAIL.n212 9.3005
R232 VTAIL.n192 VTAIL.n191 9.3005
R233 VTAIL.n220 VTAIL.n219 9.3005
R234 VTAIL.n222 VTAIL.n221 9.3005
R235 VTAIL.n57 VTAIL.n56 9.3005
R236 VTAIL.n4 VTAIL.n3 9.3005
R237 VTAIL.n51 VTAIL.n50 9.3005
R238 VTAIL.n49 VTAIL.n48 9.3005
R239 VTAIL.n8 VTAIL.n7 9.3005
R240 VTAIL.n23 VTAIL.n22 9.3005
R241 VTAIL.n25 VTAIL.n24 9.3005
R242 VTAIL.n16 VTAIL.n15 9.3005
R243 VTAIL.n31 VTAIL.n30 9.3005
R244 VTAIL.n33 VTAIL.n32 9.3005
R245 VTAIL.n12 VTAIL.n11 9.3005
R246 VTAIL.n40 VTAIL.n39 9.3005
R247 VTAIL.n42 VTAIL.n41 9.3005
R248 VTAIL.n146 VTAIL.n145 9.3005
R249 VTAIL.n148 VTAIL.n147 9.3005
R250 VTAIL.n139 VTAIL.n138 9.3005
R251 VTAIL.n154 VTAIL.n153 9.3005
R252 VTAIL.n156 VTAIL.n155 9.3005
R253 VTAIL.n134 VTAIL.n133 9.3005
R254 VTAIL.n162 VTAIL.n161 9.3005
R255 VTAIL.n164 VTAIL.n163 9.3005
R256 VTAIL.n179 VTAIL.n178 9.3005
R257 VTAIL.n126 VTAIL.n125 9.3005
R258 VTAIL.n173 VTAIL.n172 9.3005
R259 VTAIL.n171 VTAIL.n170 9.3005
R260 VTAIL.n130 VTAIL.n129 9.3005
R261 VTAIL.n86 VTAIL.n85 9.3005
R262 VTAIL.n88 VTAIL.n87 9.3005
R263 VTAIL.n79 VTAIL.n78 9.3005
R264 VTAIL.n94 VTAIL.n93 9.3005
R265 VTAIL.n96 VTAIL.n95 9.3005
R266 VTAIL.n74 VTAIL.n73 9.3005
R267 VTAIL.n102 VTAIL.n101 9.3005
R268 VTAIL.n104 VTAIL.n103 9.3005
R269 VTAIL.n119 VTAIL.n118 9.3005
R270 VTAIL.n66 VTAIL.n65 9.3005
R271 VTAIL.n113 VTAIL.n112 9.3005
R272 VTAIL.n111 VTAIL.n110 9.3005
R273 VTAIL.n70 VTAIL.n69 9.3005
R274 VTAIL.n206 VTAIL.n196 8.92171
R275 VTAIL.n26 VTAIL.n16 8.92171
R276 VTAIL.n149 VTAIL.n139 8.92171
R277 VTAIL.n89 VTAIL.n79 8.92171
R278 VTAIL.n205 VTAIL.n198 8.14595
R279 VTAIL.n25 VTAIL.n18 8.14595
R280 VTAIL.n148 VTAIL.n141 8.14595
R281 VTAIL.n88 VTAIL.n81 8.14595
R282 VTAIL.n202 VTAIL.n201 7.3702
R283 VTAIL.n22 VTAIL.n21 7.3702
R284 VTAIL.n145 VTAIL.n144 7.3702
R285 VTAIL.n85 VTAIL.n84 7.3702
R286 VTAIL.n202 VTAIL.n198 5.81868
R287 VTAIL.n22 VTAIL.n18 5.81868
R288 VTAIL.n145 VTAIL.n141 5.81868
R289 VTAIL.n85 VTAIL.n81 5.81868
R290 VTAIL.n206 VTAIL.n205 5.04292
R291 VTAIL.n26 VTAIL.n25 5.04292
R292 VTAIL.n149 VTAIL.n148 5.04292
R293 VTAIL.n89 VTAIL.n88 5.04292
R294 VTAIL.n209 VTAIL.n196 4.26717
R295 VTAIL.n238 VTAIL.n182 4.26717
R296 VTAIL.n29 VTAIL.n16 4.26717
R297 VTAIL.n58 VTAIL.n2 4.26717
R298 VTAIL.n180 VTAIL.n124 4.26717
R299 VTAIL.n152 VTAIL.n139 4.26717
R300 VTAIL.n120 VTAIL.n64 4.26717
R301 VTAIL.n92 VTAIL.n79 4.26717
R302 VTAIL.n210 VTAIL.n194 3.49141
R303 VTAIL.n236 VTAIL.n235 3.49141
R304 VTAIL.n30 VTAIL.n14 3.49141
R305 VTAIL.n56 VTAIL.n55 3.49141
R306 VTAIL.n178 VTAIL.n177 3.49141
R307 VTAIL.n153 VTAIL.n137 3.49141
R308 VTAIL.n118 VTAIL.n117 3.49141
R309 VTAIL.n93 VTAIL.n77 3.49141
R310 VTAIL.n0 VTAIL.t6 3.06123
R311 VTAIL.n0 VTAIL.t10 3.06123
R312 VTAIL.n60 VTAIL.t5 3.06123
R313 VTAIL.n60 VTAIL.t2 3.06123
R314 VTAIL.n122 VTAIL.t4 3.06123
R315 VTAIL.n122 VTAIL.t0 3.06123
R316 VTAIL.n62 VTAIL.t11 3.06123
R317 VTAIL.n62 VTAIL.t9 3.06123
R318 VTAIL.n214 VTAIL.n213 2.71565
R319 VTAIL.n232 VTAIL.n184 2.71565
R320 VTAIL.n34 VTAIL.n33 2.71565
R321 VTAIL.n52 VTAIL.n4 2.71565
R322 VTAIL.n174 VTAIL.n126 2.71565
R323 VTAIL.n157 VTAIL.n156 2.71565
R324 VTAIL.n114 VTAIL.n66 2.71565
R325 VTAIL.n97 VTAIL.n96 2.71565
R326 VTAIL.n203 VTAIL.n199 2.41282
R327 VTAIL.n23 VTAIL.n19 2.41282
R328 VTAIL.n146 VTAIL.n142 2.41282
R329 VTAIL.n86 VTAIL.n82 2.41282
R330 VTAIL.n121 VTAIL.n63 2.10395
R331 VTAIL.n181 VTAIL.n123 2.10395
R332 VTAIL.n61 VTAIL.n59 2.10395
R333 VTAIL.n218 VTAIL.n192 1.93989
R334 VTAIL.n231 VTAIL.n186 1.93989
R335 VTAIL.n38 VTAIL.n12 1.93989
R336 VTAIL.n51 VTAIL.n6 1.93989
R337 VTAIL.n173 VTAIL.n128 1.93989
R338 VTAIL.n160 VTAIL.n134 1.93989
R339 VTAIL.n113 VTAIL.n68 1.93989
R340 VTAIL.n100 VTAIL.n74 1.93989
R341 VTAIL.n123 VTAIL.n121 1.52205
R342 VTAIL.n59 VTAIL.n1 1.52205
R343 VTAIL VTAIL.n239 1.5199
R344 VTAIL.n219 VTAIL.n190 1.16414
R345 VTAIL.n228 VTAIL.n227 1.16414
R346 VTAIL.n39 VTAIL.n10 1.16414
R347 VTAIL.n48 VTAIL.n47 1.16414
R348 VTAIL.n170 VTAIL.n169 1.16414
R349 VTAIL.n161 VTAIL.n132 1.16414
R350 VTAIL.n110 VTAIL.n109 1.16414
R351 VTAIL.n101 VTAIL.n72 1.16414
R352 VTAIL VTAIL.n1 0.584552
R353 VTAIL.n223 VTAIL.n222 0.388379
R354 VTAIL.n224 VTAIL.n188 0.388379
R355 VTAIL.n43 VTAIL.n42 0.388379
R356 VTAIL.n44 VTAIL.n8 0.388379
R357 VTAIL.n166 VTAIL.n130 0.388379
R358 VTAIL.n165 VTAIL.n164 0.388379
R359 VTAIL.n106 VTAIL.n70 0.388379
R360 VTAIL.n105 VTAIL.n104 0.388379
R361 VTAIL.n204 VTAIL.n203 0.155672
R362 VTAIL.n204 VTAIL.n195 0.155672
R363 VTAIL.n211 VTAIL.n195 0.155672
R364 VTAIL.n212 VTAIL.n211 0.155672
R365 VTAIL.n212 VTAIL.n191 0.155672
R366 VTAIL.n220 VTAIL.n191 0.155672
R367 VTAIL.n221 VTAIL.n220 0.155672
R368 VTAIL.n221 VTAIL.n187 0.155672
R369 VTAIL.n229 VTAIL.n187 0.155672
R370 VTAIL.n230 VTAIL.n229 0.155672
R371 VTAIL.n230 VTAIL.n183 0.155672
R372 VTAIL.n237 VTAIL.n183 0.155672
R373 VTAIL.n24 VTAIL.n23 0.155672
R374 VTAIL.n24 VTAIL.n15 0.155672
R375 VTAIL.n31 VTAIL.n15 0.155672
R376 VTAIL.n32 VTAIL.n31 0.155672
R377 VTAIL.n32 VTAIL.n11 0.155672
R378 VTAIL.n40 VTAIL.n11 0.155672
R379 VTAIL.n41 VTAIL.n40 0.155672
R380 VTAIL.n41 VTAIL.n7 0.155672
R381 VTAIL.n49 VTAIL.n7 0.155672
R382 VTAIL.n50 VTAIL.n49 0.155672
R383 VTAIL.n50 VTAIL.n3 0.155672
R384 VTAIL.n57 VTAIL.n3 0.155672
R385 VTAIL.n179 VTAIL.n125 0.155672
R386 VTAIL.n172 VTAIL.n125 0.155672
R387 VTAIL.n172 VTAIL.n171 0.155672
R388 VTAIL.n171 VTAIL.n129 0.155672
R389 VTAIL.n163 VTAIL.n129 0.155672
R390 VTAIL.n163 VTAIL.n162 0.155672
R391 VTAIL.n162 VTAIL.n133 0.155672
R392 VTAIL.n155 VTAIL.n133 0.155672
R393 VTAIL.n155 VTAIL.n154 0.155672
R394 VTAIL.n154 VTAIL.n138 0.155672
R395 VTAIL.n147 VTAIL.n138 0.155672
R396 VTAIL.n147 VTAIL.n146 0.155672
R397 VTAIL.n119 VTAIL.n65 0.155672
R398 VTAIL.n112 VTAIL.n65 0.155672
R399 VTAIL.n112 VTAIL.n111 0.155672
R400 VTAIL.n111 VTAIL.n69 0.155672
R401 VTAIL.n103 VTAIL.n69 0.155672
R402 VTAIL.n103 VTAIL.n102 0.155672
R403 VTAIL.n102 VTAIL.n73 0.155672
R404 VTAIL.n95 VTAIL.n73 0.155672
R405 VTAIL.n95 VTAIL.n94 0.155672
R406 VTAIL.n94 VTAIL.n78 0.155672
R407 VTAIL.n87 VTAIL.n78 0.155672
R408 VTAIL.n87 VTAIL.n86 0.155672
R409 VDD2.n111 VDD2.n59 756.745
R410 VDD2.n52 VDD2.n0 756.745
R411 VDD2.n112 VDD2.n111 585
R412 VDD2.n110 VDD2.n109 585
R413 VDD2.n63 VDD2.n62 585
R414 VDD2.n104 VDD2.n103 585
R415 VDD2.n102 VDD2.n101 585
R416 VDD2.n100 VDD2.n66 585
R417 VDD2.n70 VDD2.n67 585
R418 VDD2.n95 VDD2.n94 585
R419 VDD2.n93 VDD2.n92 585
R420 VDD2.n72 VDD2.n71 585
R421 VDD2.n87 VDD2.n86 585
R422 VDD2.n85 VDD2.n84 585
R423 VDD2.n76 VDD2.n75 585
R424 VDD2.n79 VDD2.n78 585
R425 VDD2.n19 VDD2.n18 585
R426 VDD2.n16 VDD2.n15 585
R427 VDD2.n25 VDD2.n24 585
R428 VDD2.n27 VDD2.n26 585
R429 VDD2.n12 VDD2.n11 585
R430 VDD2.n33 VDD2.n32 585
R431 VDD2.n36 VDD2.n35 585
R432 VDD2.n34 VDD2.n8 585
R433 VDD2.n41 VDD2.n7 585
R434 VDD2.n43 VDD2.n42 585
R435 VDD2.n45 VDD2.n44 585
R436 VDD2.n4 VDD2.n3 585
R437 VDD2.n51 VDD2.n50 585
R438 VDD2.n53 VDD2.n52 585
R439 VDD2.t3 VDD2.n77 329.038
R440 VDD2.t4 VDD2.n17 329.038
R441 VDD2.n111 VDD2.n110 171.744
R442 VDD2.n110 VDD2.n62 171.744
R443 VDD2.n103 VDD2.n62 171.744
R444 VDD2.n103 VDD2.n102 171.744
R445 VDD2.n102 VDD2.n66 171.744
R446 VDD2.n70 VDD2.n66 171.744
R447 VDD2.n94 VDD2.n70 171.744
R448 VDD2.n94 VDD2.n93 171.744
R449 VDD2.n93 VDD2.n71 171.744
R450 VDD2.n86 VDD2.n71 171.744
R451 VDD2.n86 VDD2.n85 171.744
R452 VDD2.n85 VDD2.n75 171.744
R453 VDD2.n78 VDD2.n75 171.744
R454 VDD2.n18 VDD2.n15 171.744
R455 VDD2.n25 VDD2.n15 171.744
R456 VDD2.n26 VDD2.n25 171.744
R457 VDD2.n26 VDD2.n11 171.744
R458 VDD2.n33 VDD2.n11 171.744
R459 VDD2.n35 VDD2.n33 171.744
R460 VDD2.n35 VDD2.n34 171.744
R461 VDD2.n34 VDD2.n7 171.744
R462 VDD2.n43 VDD2.n7 171.744
R463 VDD2.n44 VDD2.n43 171.744
R464 VDD2.n44 VDD2.n3 171.744
R465 VDD2.n51 VDD2.n3 171.744
R466 VDD2.n52 VDD2.n51 171.744
R467 VDD2.n78 VDD2.t3 85.8723
R468 VDD2.n18 VDD2.t4 85.8723
R469 VDD2.n58 VDD2.n57 75.1729
R470 VDD2 VDD2.n117 75.17
R471 VDD2.n58 VDD2.n56 49.2227
R472 VDD2.n116 VDD2.n115 47.7005
R473 VDD2.n116 VDD2.n58 39.7067
R474 VDD2.n101 VDD2.n100 13.1884
R475 VDD2.n42 VDD2.n41 13.1884
R476 VDD2.n104 VDD2.n65 12.8005
R477 VDD2.n99 VDD2.n67 12.8005
R478 VDD2.n40 VDD2.n8 12.8005
R479 VDD2.n45 VDD2.n6 12.8005
R480 VDD2.n105 VDD2.n63 12.0247
R481 VDD2.n96 VDD2.n95 12.0247
R482 VDD2.n37 VDD2.n36 12.0247
R483 VDD2.n46 VDD2.n4 12.0247
R484 VDD2.n109 VDD2.n108 11.249
R485 VDD2.n92 VDD2.n69 11.249
R486 VDD2.n32 VDD2.n10 11.249
R487 VDD2.n50 VDD2.n49 11.249
R488 VDD2.n79 VDD2.n77 10.7239
R489 VDD2.n19 VDD2.n17 10.7239
R490 VDD2.n112 VDD2.n61 10.4732
R491 VDD2.n91 VDD2.n72 10.4732
R492 VDD2.n31 VDD2.n12 10.4732
R493 VDD2.n53 VDD2.n2 10.4732
R494 VDD2.n113 VDD2.n59 9.69747
R495 VDD2.n88 VDD2.n87 9.69747
R496 VDD2.n28 VDD2.n27 9.69747
R497 VDD2.n54 VDD2.n0 9.69747
R498 VDD2.n115 VDD2.n114 9.45567
R499 VDD2.n56 VDD2.n55 9.45567
R500 VDD2.n81 VDD2.n80 9.3005
R501 VDD2.n83 VDD2.n82 9.3005
R502 VDD2.n74 VDD2.n73 9.3005
R503 VDD2.n89 VDD2.n88 9.3005
R504 VDD2.n91 VDD2.n90 9.3005
R505 VDD2.n69 VDD2.n68 9.3005
R506 VDD2.n97 VDD2.n96 9.3005
R507 VDD2.n99 VDD2.n98 9.3005
R508 VDD2.n114 VDD2.n113 9.3005
R509 VDD2.n61 VDD2.n60 9.3005
R510 VDD2.n108 VDD2.n107 9.3005
R511 VDD2.n106 VDD2.n105 9.3005
R512 VDD2.n65 VDD2.n64 9.3005
R513 VDD2.n55 VDD2.n54 9.3005
R514 VDD2.n2 VDD2.n1 9.3005
R515 VDD2.n49 VDD2.n48 9.3005
R516 VDD2.n47 VDD2.n46 9.3005
R517 VDD2.n6 VDD2.n5 9.3005
R518 VDD2.n21 VDD2.n20 9.3005
R519 VDD2.n23 VDD2.n22 9.3005
R520 VDD2.n14 VDD2.n13 9.3005
R521 VDD2.n29 VDD2.n28 9.3005
R522 VDD2.n31 VDD2.n30 9.3005
R523 VDD2.n10 VDD2.n9 9.3005
R524 VDD2.n38 VDD2.n37 9.3005
R525 VDD2.n40 VDD2.n39 9.3005
R526 VDD2.n84 VDD2.n74 8.92171
R527 VDD2.n24 VDD2.n14 8.92171
R528 VDD2.n83 VDD2.n76 8.14595
R529 VDD2.n23 VDD2.n16 8.14595
R530 VDD2.n80 VDD2.n79 7.3702
R531 VDD2.n20 VDD2.n19 7.3702
R532 VDD2.n80 VDD2.n76 5.81868
R533 VDD2.n20 VDD2.n16 5.81868
R534 VDD2.n84 VDD2.n83 5.04292
R535 VDD2.n24 VDD2.n23 5.04292
R536 VDD2.n115 VDD2.n59 4.26717
R537 VDD2.n87 VDD2.n74 4.26717
R538 VDD2.n27 VDD2.n14 4.26717
R539 VDD2.n56 VDD2.n0 4.26717
R540 VDD2.n113 VDD2.n112 3.49141
R541 VDD2.n88 VDD2.n72 3.49141
R542 VDD2.n28 VDD2.n12 3.49141
R543 VDD2.n54 VDD2.n53 3.49141
R544 VDD2.n117 VDD2.t0 3.06123
R545 VDD2.n117 VDD2.t2 3.06123
R546 VDD2.n57 VDD2.t1 3.06123
R547 VDD2.n57 VDD2.t5 3.06123
R548 VDD2.n109 VDD2.n61 2.71565
R549 VDD2.n92 VDD2.n91 2.71565
R550 VDD2.n32 VDD2.n31 2.71565
R551 VDD2.n50 VDD2.n2 2.71565
R552 VDD2.n81 VDD2.n77 2.41282
R553 VDD2.n21 VDD2.n17 2.41282
R554 VDD2.n108 VDD2.n63 1.93989
R555 VDD2.n95 VDD2.n69 1.93989
R556 VDD2.n36 VDD2.n10 1.93989
R557 VDD2.n49 VDD2.n4 1.93989
R558 VDD2 VDD2.n116 1.63628
R559 VDD2.n105 VDD2.n104 1.16414
R560 VDD2.n96 VDD2.n67 1.16414
R561 VDD2.n37 VDD2.n8 1.16414
R562 VDD2.n46 VDD2.n45 1.16414
R563 VDD2.n101 VDD2.n65 0.388379
R564 VDD2.n100 VDD2.n99 0.388379
R565 VDD2.n41 VDD2.n40 0.388379
R566 VDD2.n42 VDD2.n6 0.388379
R567 VDD2.n114 VDD2.n60 0.155672
R568 VDD2.n107 VDD2.n60 0.155672
R569 VDD2.n107 VDD2.n106 0.155672
R570 VDD2.n106 VDD2.n64 0.155672
R571 VDD2.n98 VDD2.n64 0.155672
R572 VDD2.n98 VDD2.n97 0.155672
R573 VDD2.n97 VDD2.n68 0.155672
R574 VDD2.n90 VDD2.n68 0.155672
R575 VDD2.n90 VDD2.n89 0.155672
R576 VDD2.n89 VDD2.n73 0.155672
R577 VDD2.n82 VDD2.n73 0.155672
R578 VDD2.n82 VDD2.n81 0.155672
R579 VDD2.n22 VDD2.n21 0.155672
R580 VDD2.n22 VDD2.n13 0.155672
R581 VDD2.n29 VDD2.n13 0.155672
R582 VDD2.n30 VDD2.n29 0.155672
R583 VDD2.n30 VDD2.n9 0.155672
R584 VDD2.n38 VDD2.n9 0.155672
R585 VDD2.n39 VDD2.n38 0.155672
R586 VDD2.n39 VDD2.n5 0.155672
R587 VDD2.n47 VDD2.n5 0.155672
R588 VDD2.n48 VDD2.n47 0.155672
R589 VDD2.n48 VDD2.n1 0.155672
R590 VDD2.n55 VDD2.n1 0.155672
R591 VP.n10 VP.n9 161.3
R592 VP.n11 VP.n6 161.3
R593 VP.n13 VP.n12 161.3
R594 VP.n14 VP.n5 161.3
R595 VP.n31 VP.n0 161.3
R596 VP.n30 VP.n29 161.3
R597 VP.n28 VP.n1 161.3
R598 VP.n27 VP.n26 161.3
R599 VP.n25 VP.n2 161.3
R600 VP.n24 VP.n23 161.3
R601 VP.n22 VP.n3 161.3
R602 VP.n21 VP.n20 161.3
R603 VP.n19 VP.n4 161.3
R604 VP.n7 VP.t5 155.772
R605 VP.n25 VP.t4 121.3
R606 VP.n18 VP.t0 121.3
R607 VP.n32 VP.t2 121.3
R608 VP.n8 VP.t1 121.3
R609 VP.n15 VP.t3 121.3
R610 VP.n18 VP.n17 89.2674
R611 VP.n33 VP.n32 89.2674
R612 VP.n16 VP.n15 89.2674
R613 VP.n20 VP.n3 56.5617
R614 VP.n30 VP.n1 56.5617
R615 VP.n13 VP.n6 56.5617
R616 VP.n8 VP.n7 46.3186
R617 VP.n17 VP.n16 45.7875
R618 VP.n20 VP.n19 24.5923
R619 VP.n24 VP.n3 24.5923
R620 VP.n25 VP.n24 24.5923
R621 VP.n26 VP.n25 24.5923
R622 VP.n26 VP.n1 24.5923
R623 VP.n31 VP.n30 24.5923
R624 VP.n14 VP.n13 24.5923
R625 VP.n9 VP.n8 24.5923
R626 VP.n9 VP.n6 24.5923
R627 VP.n19 VP.n18 21.6413
R628 VP.n32 VP.n31 21.6413
R629 VP.n15 VP.n14 21.6413
R630 VP.n10 VP.n7 8.80512
R631 VP.n16 VP.n5 0.278335
R632 VP.n17 VP.n4 0.278335
R633 VP.n33 VP.n0 0.278335
R634 VP.n11 VP.n10 0.189894
R635 VP.n12 VP.n11 0.189894
R636 VP.n12 VP.n5 0.189894
R637 VP.n21 VP.n4 0.189894
R638 VP.n22 VP.n21 0.189894
R639 VP.n23 VP.n22 0.189894
R640 VP.n23 VP.n2 0.189894
R641 VP.n27 VP.n2 0.189894
R642 VP.n28 VP.n27 0.189894
R643 VP.n29 VP.n28 0.189894
R644 VP.n29 VP.n0 0.189894
R645 VP VP.n33 0.153485
R646 VDD1.n52 VDD1.n0 756.745
R647 VDD1.n109 VDD1.n57 756.745
R648 VDD1.n53 VDD1.n52 585
R649 VDD1.n51 VDD1.n50 585
R650 VDD1.n4 VDD1.n3 585
R651 VDD1.n45 VDD1.n44 585
R652 VDD1.n43 VDD1.n42 585
R653 VDD1.n41 VDD1.n7 585
R654 VDD1.n11 VDD1.n8 585
R655 VDD1.n36 VDD1.n35 585
R656 VDD1.n34 VDD1.n33 585
R657 VDD1.n13 VDD1.n12 585
R658 VDD1.n28 VDD1.n27 585
R659 VDD1.n26 VDD1.n25 585
R660 VDD1.n17 VDD1.n16 585
R661 VDD1.n20 VDD1.n19 585
R662 VDD1.n76 VDD1.n75 585
R663 VDD1.n73 VDD1.n72 585
R664 VDD1.n82 VDD1.n81 585
R665 VDD1.n84 VDD1.n83 585
R666 VDD1.n69 VDD1.n68 585
R667 VDD1.n90 VDD1.n89 585
R668 VDD1.n93 VDD1.n92 585
R669 VDD1.n91 VDD1.n65 585
R670 VDD1.n98 VDD1.n64 585
R671 VDD1.n100 VDD1.n99 585
R672 VDD1.n102 VDD1.n101 585
R673 VDD1.n61 VDD1.n60 585
R674 VDD1.n108 VDD1.n107 585
R675 VDD1.n110 VDD1.n109 585
R676 VDD1.t0 VDD1.n18 329.038
R677 VDD1.t5 VDD1.n74 329.038
R678 VDD1.n52 VDD1.n51 171.744
R679 VDD1.n51 VDD1.n3 171.744
R680 VDD1.n44 VDD1.n3 171.744
R681 VDD1.n44 VDD1.n43 171.744
R682 VDD1.n43 VDD1.n7 171.744
R683 VDD1.n11 VDD1.n7 171.744
R684 VDD1.n35 VDD1.n11 171.744
R685 VDD1.n35 VDD1.n34 171.744
R686 VDD1.n34 VDD1.n12 171.744
R687 VDD1.n27 VDD1.n12 171.744
R688 VDD1.n27 VDD1.n26 171.744
R689 VDD1.n26 VDD1.n16 171.744
R690 VDD1.n19 VDD1.n16 171.744
R691 VDD1.n75 VDD1.n72 171.744
R692 VDD1.n82 VDD1.n72 171.744
R693 VDD1.n83 VDD1.n82 171.744
R694 VDD1.n83 VDD1.n68 171.744
R695 VDD1.n90 VDD1.n68 171.744
R696 VDD1.n92 VDD1.n90 171.744
R697 VDD1.n92 VDD1.n91 171.744
R698 VDD1.n91 VDD1.n64 171.744
R699 VDD1.n100 VDD1.n64 171.744
R700 VDD1.n101 VDD1.n100 171.744
R701 VDD1.n101 VDD1.n60 171.744
R702 VDD1.n108 VDD1.n60 171.744
R703 VDD1.n109 VDD1.n108 171.744
R704 VDD1.n19 VDD1.t0 85.8723
R705 VDD1.n75 VDD1.t5 85.8723
R706 VDD1.n115 VDD1.n114 75.1729
R707 VDD1.n117 VDD1.n116 74.7023
R708 VDD1 VDD1.n56 49.3363
R709 VDD1.n115 VDD1.n113 49.2227
R710 VDD1.n117 VDD1.n115 41.3414
R711 VDD1.n42 VDD1.n41 13.1884
R712 VDD1.n99 VDD1.n98 13.1884
R713 VDD1.n45 VDD1.n6 12.8005
R714 VDD1.n40 VDD1.n8 12.8005
R715 VDD1.n97 VDD1.n65 12.8005
R716 VDD1.n102 VDD1.n63 12.8005
R717 VDD1.n46 VDD1.n4 12.0247
R718 VDD1.n37 VDD1.n36 12.0247
R719 VDD1.n94 VDD1.n93 12.0247
R720 VDD1.n103 VDD1.n61 12.0247
R721 VDD1.n50 VDD1.n49 11.249
R722 VDD1.n33 VDD1.n10 11.249
R723 VDD1.n89 VDD1.n67 11.249
R724 VDD1.n107 VDD1.n106 11.249
R725 VDD1.n20 VDD1.n18 10.7239
R726 VDD1.n76 VDD1.n74 10.7239
R727 VDD1.n53 VDD1.n2 10.4732
R728 VDD1.n32 VDD1.n13 10.4732
R729 VDD1.n88 VDD1.n69 10.4732
R730 VDD1.n110 VDD1.n59 10.4732
R731 VDD1.n54 VDD1.n0 9.69747
R732 VDD1.n29 VDD1.n28 9.69747
R733 VDD1.n85 VDD1.n84 9.69747
R734 VDD1.n111 VDD1.n57 9.69747
R735 VDD1.n56 VDD1.n55 9.45567
R736 VDD1.n113 VDD1.n112 9.45567
R737 VDD1.n22 VDD1.n21 9.3005
R738 VDD1.n24 VDD1.n23 9.3005
R739 VDD1.n15 VDD1.n14 9.3005
R740 VDD1.n30 VDD1.n29 9.3005
R741 VDD1.n32 VDD1.n31 9.3005
R742 VDD1.n10 VDD1.n9 9.3005
R743 VDD1.n38 VDD1.n37 9.3005
R744 VDD1.n40 VDD1.n39 9.3005
R745 VDD1.n55 VDD1.n54 9.3005
R746 VDD1.n2 VDD1.n1 9.3005
R747 VDD1.n49 VDD1.n48 9.3005
R748 VDD1.n47 VDD1.n46 9.3005
R749 VDD1.n6 VDD1.n5 9.3005
R750 VDD1.n112 VDD1.n111 9.3005
R751 VDD1.n59 VDD1.n58 9.3005
R752 VDD1.n106 VDD1.n105 9.3005
R753 VDD1.n104 VDD1.n103 9.3005
R754 VDD1.n63 VDD1.n62 9.3005
R755 VDD1.n78 VDD1.n77 9.3005
R756 VDD1.n80 VDD1.n79 9.3005
R757 VDD1.n71 VDD1.n70 9.3005
R758 VDD1.n86 VDD1.n85 9.3005
R759 VDD1.n88 VDD1.n87 9.3005
R760 VDD1.n67 VDD1.n66 9.3005
R761 VDD1.n95 VDD1.n94 9.3005
R762 VDD1.n97 VDD1.n96 9.3005
R763 VDD1.n25 VDD1.n15 8.92171
R764 VDD1.n81 VDD1.n71 8.92171
R765 VDD1.n24 VDD1.n17 8.14595
R766 VDD1.n80 VDD1.n73 8.14595
R767 VDD1.n21 VDD1.n20 7.3702
R768 VDD1.n77 VDD1.n76 7.3702
R769 VDD1.n21 VDD1.n17 5.81868
R770 VDD1.n77 VDD1.n73 5.81868
R771 VDD1.n25 VDD1.n24 5.04292
R772 VDD1.n81 VDD1.n80 5.04292
R773 VDD1.n56 VDD1.n0 4.26717
R774 VDD1.n28 VDD1.n15 4.26717
R775 VDD1.n84 VDD1.n71 4.26717
R776 VDD1.n113 VDD1.n57 4.26717
R777 VDD1.n54 VDD1.n53 3.49141
R778 VDD1.n29 VDD1.n13 3.49141
R779 VDD1.n85 VDD1.n69 3.49141
R780 VDD1.n111 VDD1.n110 3.49141
R781 VDD1.n116 VDD1.t4 3.06123
R782 VDD1.n116 VDD1.t2 3.06123
R783 VDD1.n114 VDD1.t1 3.06123
R784 VDD1.n114 VDD1.t3 3.06123
R785 VDD1.n50 VDD1.n2 2.71565
R786 VDD1.n33 VDD1.n32 2.71565
R787 VDD1.n89 VDD1.n88 2.71565
R788 VDD1.n107 VDD1.n59 2.71565
R789 VDD1.n22 VDD1.n18 2.41282
R790 VDD1.n78 VDD1.n74 2.41282
R791 VDD1.n49 VDD1.n4 1.93989
R792 VDD1.n36 VDD1.n10 1.93989
R793 VDD1.n93 VDD1.n67 1.93989
R794 VDD1.n106 VDD1.n61 1.93989
R795 VDD1.n46 VDD1.n45 1.16414
R796 VDD1.n37 VDD1.n8 1.16414
R797 VDD1.n94 VDD1.n65 1.16414
R798 VDD1.n103 VDD1.n102 1.16414
R799 VDD1 VDD1.n117 0.468172
R800 VDD1.n42 VDD1.n6 0.388379
R801 VDD1.n41 VDD1.n40 0.388379
R802 VDD1.n98 VDD1.n97 0.388379
R803 VDD1.n99 VDD1.n63 0.388379
R804 VDD1.n55 VDD1.n1 0.155672
R805 VDD1.n48 VDD1.n1 0.155672
R806 VDD1.n48 VDD1.n47 0.155672
R807 VDD1.n47 VDD1.n5 0.155672
R808 VDD1.n39 VDD1.n5 0.155672
R809 VDD1.n39 VDD1.n38 0.155672
R810 VDD1.n38 VDD1.n9 0.155672
R811 VDD1.n31 VDD1.n9 0.155672
R812 VDD1.n31 VDD1.n30 0.155672
R813 VDD1.n30 VDD1.n14 0.155672
R814 VDD1.n23 VDD1.n14 0.155672
R815 VDD1.n23 VDD1.n22 0.155672
R816 VDD1.n79 VDD1.n78 0.155672
R817 VDD1.n79 VDD1.n70 0.155672
R818 VDD1.n86 VDD1.n70 0.155672
R819 VDD1.n87 VDD1.n86 0.155672
R820 VDD1.n87 VDD1.n66 0.155672
R821 VDD1.n95 VDD1.n66 0.155672
R822 VDD1.n96 VDD1.n95 0.155672
R823 VDD1.n96 VDD1.n62 0.155672
R824 VDD1.n104 VDD1.n62 0.155672
R825 VDD1.n105 VDD1.n104 0.155672
R826 VDD1.n105 VDD1.n58 0.155672
R827 VDD1.n112 VDD1.n58 0.155672
R828 B.n466 B.n67 585
R829 B.n468 B.n467 585
R830 B.n469 B.n66 585
R831 B.n471 B.n470 585
R832 B.n472 B.n65 585
R833 B.n474 B.n473 585
R834 B.n475 B.n64 585
R835 B.n477 B.n476 585
R836 B.n478 B.n63 585
R837 B.n480 B.n479 585
R838 B.n481 B.n62 585
R839 B.n483 B.n482 585
R840 B.n484 B.n61 585
R841 B.n486 B.n485 585
R842 B.n487 B.n60 585
R843 B.n489 B.n488 585
R844 B.n490 B.n59 585
R845 B.n492 B.n491 585
R846 B.n493 B.n58 585
R847 B.n495 B.n494 585
R848 B.n496 B.n57 585
R849 B.n498 B.n497 585
R850 B.n499 B.n56 585
R851 B.n501 B.n500 585
R852 B.n502 B.n55 585
R853 B.n504 B.n503 585
R854 B.n505 B.n54 585
R855 B.n507 B.n506 585
R856 B.n508 B.n53 585
R857 B.n510 B.n509 585
R858 B.n511 B.n52 585
R859 B.n513 B.n512 585
R860 B.n514 B.n51 585
R861 B.n516 B.n515 585
R862 B.n517 B.n50 585
R863 B.n519 B.n518 585
R864 B.n520 B.n49 585
R865 B.n522 B.n521 585
R866 B.n524 B.n523 585
R867 B.n525 B.n45 585
R868 B.n527 B.n526 585
R869 B.n528 B.n44 585
R870 B.n530 B.n529 585
R871 B.n531 B.n43 585
R872 B.n533 B.n532 585
R873 B.n534 B.n42 585
R874 B.n536 B.n535 585
R875 B.n538 B.n39 585
R876 B.n540 B.n539 585
R877 B.n541 B.n38 585
R878 B.n543 B.n542 585
R879 B.n544 B.n37 585
R880 B.n546 B.n545 585
R881 B.n547 B.n36 585
R882 B.n549 B.n548 585
R883 B.n550 B.n35 585
R884 B.n552 B.n551 585
R885 B.n553 B.n34 585
R886 B.n555 B.n554 585
R887 B.n556 B.n33 585
R888 B.n558 B.n557 585
R889 B.n559 B.n32 585
R890 B.n561 B.n560 585
R891 B.n562 B.n31 585
R892 B.n564 B.n563 585
R893 B.n565 B.n30 585
R894 B.n567 B.n566 585
R895 B.n568 B.n29 585
R896 B.n570 B.n569 585
R897 B.n571 B.n28 585
R898 B.n573 B.n572 585
R899 B.n574 B.n27 585
R900 B.n576 B.n575 585
R901 B.n577 B.n26 585
R902 B.n579 B.n578 585
R903 B.n580 B.n25 585
R904 B.n582 B.n581 585
R905 B.n583 B.n24 585
R906 B.n585 B.n584 585
R907 B.n586 B.n23 585
R908 B.n588 B.n587 585
R909 B.n589 B.n22 585
R910 B.n591 B.n590 585
R911 B.n592 B.n21 585
R912 B.n594 B.n593 585
R913 B.n465 B.n464 585
R914 B.n463 B.n68 585
R915 B.n462 B.n461 585
R916 B.n460 B.n69 585
R917 B.n459 B.n458 585
R918 B.n457 B.n70 585
R919 B.n456 B.n455 585
R920 B.n454 B.n71 585
R921 B.n453 B.n452 585
R922 B.n451 B.n72 585
R923 B.n450 B.n449 585
R924 B.n448 B.n73 585
R925 B.n447 B.n446 585
R926 B.n445 B.n74 585
R927 B.n444 B.n443 585
R928 B.n442 B.n75 585
R929 B.n441 B.n440 585
R930 B.n439 B.n76 585
R931 B.n438 B.n437 585
R932 B.n436 B.n77 585
R933 B.n435 B.n434 585
R934 B.n433 B.n78 585
R935 B.n432 B.n431 585
R936 B.n430 B.n79 585
R937 B.n429 B.n428 585
R938 B.n427 B.n80 585
R939 B.n426 B.n425 585
R940 B.n424 B.n81 585
R941 B.n423 B.n422 585
R942 B.n421 B.n82 585
R943 B.n420 B.n419 585
R944 B.n418 B.n83 585
R945 B.n417 B.n416 585
R946 B.n415 B.n84 585
R947 B.n414 B.n413 585
R948 B.n412 B.n85 585
R949 B.n411 B.n410 585
R950 B.n409 B.n86 585
R951 B.n408 B.n407 585
R952 B.n406 B.n87 585
R953 B.n405 B.n404 585
R954 B.n403 B.n88 585
R955 B.n402 B.n401 585
R956 B.n400 B.n89 585
R957 B.n399 B.n398 585
R958 B.n397 B.n90 585
R959 B.n396 B.n395 585
R960 B.n394 B.n91 585
R961 B.n393 B.n392 585
R962 B.n391 B.n92 585
R963 B.n390 B.n389 585
R964 B.n388 B.n93 585
R965 B.n387 B.n386 585
R966 B.n385 B.n94 585
R967 B.n384 B.n383 585
R968 B.n382 B.n95 585
R969 B.n381 B.n380 585
R970 B.n379 B.n96 585
R971 B.n378 B.n377 585
R972 B.n376 B.n97 585
R973 B.n375 B.n374 585
R974 B.n373 B.n98 585
R975 B.n372 B.n371 585
R976 B.n370 B.n99 585
R977 B.n369 B.n368 585
R978 B.n367 B.n100 585
R979 B.n366 B.n365 585
R980 B.n364 B.n101 585
R981 B.n363 B.n362 585
R982 B.n361 B.n102 585
R983 B.n360 B.n359 585
R984 B.n358 B.n103 585
R985 B.n357 B.n356 585
R986 B.n355 B.n104 585
R987 B.n354 B.n353 585
R988 B.n225 B.n224 585
R989 B.n226 B.n151 585
R990 B.n228 B.n227 585
R991 B.n229 B.n150 585
R992 B.n231 B.n230 585
R993 B.n232 B.n149 585
R994 B.n234 B.n233 585
R995 B.n235 B.n148 585
R996 B.n237 B.n236 585
R997 B.n238 B.n147 585
R998 B.n240 B.n239 585
R999 B.n241 B.n146 585
R1000 B.n243 B.n242 585
R1001 B.n244 B.n145 585
R1002 B.n246 B.n245 585
R1003 B.n247 B.n144 585
R1004 B.n249 B.n248 585
R1005 B.n250 B.n143 585
R1006 B.n252 B.n251 585
R1007 B.n253 B.n142 585
R1008 B.n255 B.n254 585
R1009 B.n256 B.n141 585
R1010 B.n258 B.n257 585
R1011 B.n259 B.n140 585
R1012 B.n261 B.n260 585
R1013 B.n262 B.n139 585
R1014 B.n264 B.n263 585
R1015 B.n265 B.n138 585
R1016 B.n267 B.n266 585
R1017 B.n268 B.n137 585
R1018 B.n270 B.n269 585
R1019 B.n271 B.n136 585
R1020 B.n273 B.n272 585
R1021 B.n274 B.n135 585
R1022 B.n276 B.n275 585
R1023 B.n277 B.n134 585
R1024 B.n279 B.n278 585
R1025 B.n280 B.n131 585
R1026 B.n283 B.n282 585
R1027 B.n284 B.n130 585
R1028 B.n286 B.n285 585
R1029 B.n287 B.n129 585
R1030 B.n289 B.n288 585
R1031 B.n290 B.n128 585
R1032 B.n292 B.n291 585
R1033 B.n293 B.n127 585
R1034 B.n295 B.n294 585
R1035 B.n297 B.n296 585
R1036 B.n298 B.n123 585
R1037 B.n300 B.n299 585
R1038 B.n301 B.n122 585
R1039 B.n303 B.n302 585
R1040 B.n304 B.n121 585
R1041 B.n306 B.n305 585
R1042 B.n307 B.n120 585
R1043 B.n309 B.n308 585
R1044 B.n310 B.n119 585
R1045 B.n312 B.n311 585
R1046 B.n313 B.n118 585
R1047 B.n315 B.n314 585
R1048 B.n316 B.n117 585
R1049 B.n318 B.n317 585
R1050 B.n319 B.n116 585
R1051 B.n321 B.n320 585
R1052 B.n322 B.n115 585
R1053 B.n324 B.n323 585
R1054 B.n325 B.n114 585
R1055 B.n327 B.n326 585
R1056 B.n328 B.n113 585
R1057 B.n330 B.n329 585
R1058 B.n331 B.n112 585
R1059 B.n333 B.n332 585
R1060 B.n334 B.n111 585
R1061 B.n336 B.n335 585
R1062 B.n337 B.n110 585
R1063 B.n339 B.n338 585
R1064 B.n340 B.n109 585
R1065 B.n342 B.n341 585
R1066 B.n343 B.n108 585
R1067 B.n345 B.n344 585
R1068 B.n346 B.n107 585
R1069 B.n348 B.n347 585
R1070 B.n349 B.n106 585
R1071 B.n351 B.n350 585
R1072 B.n352 B.n105 585
R1073 B.n223 B.n152 585
R1074 B.n222 B.n221 585
R1075 B.n220 B.n153 585
R1076 B.n219 B.n218 585
R1077 B.n217 B.n154 585
R1078 B.n216 B.n215 585
R1079 B.n214 B.n155 585
R1080 B.n213 B.n212 585
R1081 B.n211 B.n156 585
R1082 B.n210 B.n209 585
R1083 B.n208 B.n157 585
R1084 B.n207 B.n206 585
R1085 B.n205 B.n158 585
R1086 B.n204 B.n203 585
R1087 B.n202 B.n159 585
R1088 B.n201 B.n200 585
R1089 B.n199 B.n160 585
R1090 B.n198 B.n197 585
R1091 B.n196 B.n161 585
R1092 B.n195 B.n194 585
R1093 B.n193 B.n162 585
R1094 B.n192 B.n191 585
R1095 B.n190 B.n163 585
R1096 B.n189 B.n188 585
R1097 B.n187 B.n164 585
R1098 B.n186 B.n185 585
R1099 B.n184 B.n165 585
R1100 B.n183 B.n182 585
R1101 B.n181 B.n166 585
R1102 B.n180 B.n179 585
R1103 B.n178 B.n167 585
R1104 B.n177 B.n176 585
R1105 B.n175 B.n168 585
R1106 B.n174 B.n173 585
R1107 B.n172 B.n169 585
R1108 B.n171 B.n170 585
R1109 B.n2 B.n0 585
R1110 B.n649 B.n1 585
R1111 B.n648 B.n647 585
R1112 B.n646 B.n3 585
R1113 B.n645 B.n644 585
R1114 B.n643 B.n4 585
R1115 B.n642 B.n641 585
R1116 B.n640 B.n5 585
R1117 B.n639 B.n638 585
R1118 B.n637 B.n6 585
R1119 B.n636 B.n635 585
R1120 B.n634 B.n7 585
R1121 B.n633 B.n632 585
R1122 B.n631 B.n8 585
R1123 B.n630 B.n629 585
R1124 B.n628 B.n9 585
R1125 B.n627 B.n626 585
R1126 B.n625 B.n10 585
R1127 B.n624 B.n623 585
R1128 B.n622 B.n11 585
R1129 B.n621 B.n620 585
R1130 B.n619 B.n12 585
R1131 B.n618 B.n617 585
R1132 B.n616 B.n13 585
R1133 B.n615 B.n614 585
R1134 B.n613 B.n14 585
R1135 B.n612 B.n611 585
R1136 B.n610 B.n15 585
R1137 B.n609 B.n608 585
R1138 B.n607 B.n16 585
R1139 B.n606 B.n605 585
R1140 B.n604 B.n17 585
R1141 B.n603 B.n602 585
R1142 B.n601 B.n18 585
R1143 B.n600 B.n599 585
R1144 B.n598 B.n19 585
R1145 B.n597 B.n596 585
R1146 B.n595 B.n20 585
R1147 B.n651 B.n650 585
R1148 B.n224 B.n223 444.452
R1149 B.n595 B.n594 444.452
R1150 B.n354 B.n105 444.452
R1151 B.n464 B.n67 444.452
R1152 B.n124 B.t2 397.974
R1153 B.n46 B.t4 397.974
R1154 B.n132 B.t11 397.974
R1155 B.n40 B.t7 397.974
R1156 B.n125 B.t1 350.652
R1157 B.n47 B.t5 350.652
R1158 B.n133 B.t10 350.652
R1159 B.n41 B.t8 350.652
R1160 B.n124 B.t0 328.464
R1161 B.n132 B.t9 328.464
R1162 B.n40 B.t6 328.464
R1163 B.n46 B.t3 328.464
R1164 B.n223 B.n222 163.367
R1165 B.n222 B.n153 163.367
R1166 B.n218 B.n153 163.367
R1167 B.n218 B.n217 163.367
R1168 B.n217 B.n216 163.367
R1169 B.n216 B.n155 163.367
R1170 B.n212 B.n155 163.367
R1171 B.n212 B.n211 163.367
R1172 B.n211 B.n210 163.367
R1173 B.n210 B.n157 163.367
R1174 B.n206 B.n157 163.367
R1175 B.n206 B.n205 163.367
R1176 B.n205 B.n204 163.367
R1177 B.n204 B.n159 163.367
R1178 B.n200 B.n159 163.367
R1179 B.n200 B.n199 163.367
R1180 B.n199 B.n198 163.367
R1181 B.n198 B.n161 163.367
R1182 B.n194 B.n161 163.367
R1183 B.n194 B.n193 163.367
R1184 B.n193 B.n192 163.367
R1185 B.n192 B.n163 163.367
R1186 B.n188 B.n163 163.367
R1187 B.n188 B.n187 163.367
R1188 B.n187 B.n186 163.367
R1189 B.n186 B.n165 163.367
R1190 B.n182 B.n165 163.367
R1191 B.n182 B.n181 163.367
R1192 B.n181 B.n180 163.367
R1193 B.n180 B.n167 163.367
R1194 B.n176 B.n167 163.367
R1195 B.n176 B.n175 163.367
R1196 B.n175 B.n174 163.367
R1197 B.n174 B.n169 163.367
R1198 B.n170 B.n169 163.367
R1199 B.n170 B.n2 163.367
R1200 B.n650 B.n2 163.367
R1201 B.n650 B.n649 163.367
R1202 B.n649 B.n648 163.367
R1203 B.n648 B.n3 163.367
R1204 B.n644 B.n3 163.367
R1205 B.n644 B.n643 163.367
R1206 B.n643 B.n642 163.367
R1207 B.n642 B.n5 163.367
R1208 B.n638 B.n5 163.367
R1209 B.n638 B.n637 163.367
R1210 B.n637 B.n636 163.367
R1211 B.n636 B.n7 163.367
R1212 B.n632 B.n7 163.367
R1213 B.n632 B.n631 163.367
R1214 B.n631 B.n630 163.367
R1215 B.n630 B.n9 163.367
R1216 B.n626 B.n9 163.367
R1217 B.n626 B.n625 163.367
R1218 B.n625 B.n624 163.367
R1219 B.n624 B.n11 163.367
R1220 B.n620 B.n11 163.367
R1221 B.n620 B.n619 163.367
R1222 B.n619 B.n618 163.367
R1223 B.n618 B.n13 163.367
R1224 B.n614 B.n13 163.367
R1225 B.n614 B.n613 163.367
R1226 B.n613 B.n612 163.367
R1227 B.n612 B.n15 163.367
R1228 B.n608 B.n15 163.367
R1229 B.n608 B.n607 163.367
R1230 B.n607 B.n606 163.367
R1231 B.n606 B.n17 163.367
R1232 B.n602 B.n17 163.367
R1233 B.n602 B.n601 163.367
R1234 B.n601 B.n600 163.367
R1235 B.n600 B.n19 163.367
R1236 B.n596 B.n19 163.367
R1237 B.n596 B.n595 163.367
R1238 B.n224 B.n151 163.367
R1239 B.n228 B.n151 163.367
R1240 B.n229 B.n228 163.367
R1241 B.n230 B.n229 163.367
R1242 B.n230 B.n149 163.367
R1243 B.n234 B.n149 163.367
R1244 B.n235 B.n234 163.367
R1245 B.n236 B.n235 163.367
R1246 B.n236 B.n147 163.367
R1247 B.n240 B.n147 163.367
R1248 B.n241 B.n240 163.367
R1249 B.n242 B.n241 163.367
R1250 B.n242 B.n145 163.367
R1251 B.n246 B.n145 163.367
R1252 B.n247 B.n246 163.367
R1253 B.n248 B.n247 163.367
R1254 B.n248 B.n143 163.367
R1255 B.n252 B.n143 163.367
R1256 B.n253 B.n252 163.367
R1257 B.n254 B.n253 163.367
R1258 B.n254 B.n141 163.367
R1259 B.n258 B.n141 163.367
R1260 B.n259 B.n258 163.367
R1261 B.n260 B.n259 163.367
R1262 B.n260 B.n139 163.367
R1263 B.n264 B.n139 163.367
R1264 B.n265 B.n264 163.367
R1265 B.n266 B.n265 163.367
R1266 B.n266 B.n137 163.367
R1267 B.n270 B.n137 163.367
R1268 B.n271 B.n270 163.367
R1269 B.n272 B.n271 163.367
R1270 B.n272 B.n135 163.367
R1271 B.n276 B.n135 163.367
R1272 B.n277 B.n276 163.367
R1273 B.n278 B.n277 163.367
R1274 B.n278 B.n131 163.367
R1275 B.n283 B.n131 163.367
R1276 B.n284 B.n283 163.367
R1277 B.n285 B.n284 163.367
R1278 B.n285 B.n129 163.367
R1279 B.n289 B.n129 163.367
R1280 B.n290 B.n289 163.367
R1281 B.n291 B.n290 163.367
R1282 B.n291 B.n127 163.367
R1283 B.n295 B.n127 163.367
R1284 B.n296 B.n295 163.367
R1285 B.n296 B.n123 163.367
R1286 B.n300 B.n123 163.367
R1287 B.n301 B.n300 163.367
R1288 B.n302 B.n301 163.367
R1289 B.n302 B.n121 163.367
R1290 B.n306 B.n121 163.367
R1291 B.n307 B.n306 163.367
R1292 B.n308 B.n307 163.367
R1293 B.n308 B.n119 163.367
R1294 B.n312 B.n119 163.367
R1295 B.n313 B.n312 163.367
R1296 B.n314 B.n313 163.367
R1297 B.n314 B.n117 163.367
R1298 B.n318 B.n117 163.367
R1299 B.n319 B.n318 163.367
R1300 B.n320 B.n319 163.367
R1301 B.n320 B.n115 163.367
R1302 B.n324 B.n115 163.367
R1303 B.n325 B.n324 163.367
R1304 B.n326 B.n325 163.367
R1305 B.n326 B.n113 163.367
R1306 B.n330 B.n113 163.367
R1307 B.n331 B.n330 163.367
R1308 B.n332 B.n331 163.367
R1309 B.n332 B.n111 163.367
R1310 B.n336 B.n111 163.367
R1311 B.n337 B.n336 163.367
R1312 B.n338 B.n337 163.367
R1313 B.n338 B.n109 163.367
R1314 B.n342 B.n109 163.367
R1315 B.n343 B.n342 163.367
R1316 B.n344 B.n343 163.367
R1317 B.n344 B.n107 163.367
R1318 B.n348 B.n107 163.367
R1319 B.n349 B.n348 163.367
R1320 B.n350 B.n349 163.367
R1321 B.n350 B.n105 163.367
R1322 B.n355 B.n354 163.367
R1323 B.n356 B.n355 163.367
R1324 B.n356 B.n103 163.367
R1325 B.n360 B.n103 163.367
R1326 B.n361 B.n360 163.367
R1327 B.n362 B.n361 163.367
R1328 B.n362 B.n101 163.367
R1329 B.n366 B.n101 163.367
R1330 B.n367 B.n366 163.367
R1331 B.n368 B.n367 163.367
R1332 B.n368 B.n99 163.367
R1333 B.n372 B.n99 163.367
R1334 B.n373 B.n372 163.367
R1335 B.n374 B.n373 163.367
R1336 B.n374 B.n97 163.367
R1337 B.n378 B.n97 163.367
R1338 B.n379 B.n378 163.367
R1339 B.n380 B.n379 163.367
R1340 B.n380 B.n95 163.367
R1341 B.n384 B.n95 163.367
R1342 B.n385 B.n384 163.367
R1343 B.n386 B.n385 163.367
R1344 B.n386 B.n93 163.367
R1345 B.n390 B.n93 163.367
R1346 B.n391 B.n390 163.367
R1347 B.n392 B.n391 163.367
R1348 B.n392 B.n91 163.367
R1349 B.n396 B.n91 163.367
R1350 B.n397 B.n396 163.367
R1351 B.n398 B.n397 163.367
R1352 B.n398 B.n89 163.367
R1353 B.n402 B.n89 163.367
R1354 B.n403 B.n402 163.367
R1355 B.n404 B.n403 163.367
R1356 B.n404 B.n87 163.367
R1357 B.n408 B.n87 163.367
R1358 B.n409 B.n408 163.367
R1359 B.n410 B.n409 163.367
R1360 B.n410 B.n85 163.367
R1361 B.n414 B.n85 163.367
R1362 B.n415 B.n414 163.367
R1363 B.n416 B.n415 163.367
R1364 B.n416 B.n83 163.367
R1365 B.n420 B.n83 163.367
R1366 B.n421 B.n420 163.367
R1367 B.n422 B.n421 163.367
R1368 B.n422 B.n81 163.367
R1369 B.n426 B.n81 163.367
R1370 B.n427 B.n426 163.367
R1371 B.n428 B.n427 163.367
R1372 B.n428 B.n79 163.367
R1373 B.n432 B.n79 163.367
R1374 B.n433 B.n432 163.367
R1375 B.n434 B.n433 163.367
R1376 B.n434 B.n77 163.367
R1377 B.n438 B.n77 163.367
R1378 B.n439 B.n438 163.367
R1379 B.n440 B.n439 163.367
R1380 B.n440 B.n75 163.367
R1381 B.n444 B.n75 163.367
R1382 B.n445 B.n444 163.367
R1383 B.n446 B.n445 163.367
R1384 B.n446 B.n73 163.367
R1385 B.n450 B.n73 163.367
R1386 B.n451 B.n450 163.367
R1387 B.n452 B.n451 163.367
R1388 B.n452 B.n71 163.367
R1389 B.n456 B.n71 163.367
R1390 B.n457 B.n456 163.367
R1391 B.n458 B.n457 163.367
R1392 B.n458 B.n69 163.367
R1393 B.n462 B.n69 163.367
R1394 B.n463 B.n462 163.367
R1395 B.n464 B.n463 163.367
R1396 B.n594 B.n21 163.367
R1397 B.n590 B.n21 163.367
R1398 B.n590 B.n589 163.367
R1399 B.n589 B.n588 163.367
R1400 B.n588 B.n23 163.367
R1401 B.n584 B.n23 163.367
R1402 B.n584 B.n583 163.367
R1403 B.n583 B.n582 163.367
R1404 B.n582 B.n25 163.367
R1405 B.n578 B.n25 163.367
R1406 B.n578 B.n577 163.367
R1407 B.n577 B.n576 163.367
R1408 B.n576 B.n27 163.367
R1409 B.n572 B.n27 163.367
R1410 B.n572 B.n571 163.367
R1411 B.n571 B.n570 163.367
R1412 B.n570 B.n29 163.367
R1413 B.n566 B.n29 163.367
R1414 B.n566 B.n565 163.367
R1415 B.n565 B.n564 163.367
R1416 B.n564 B.n31 163.367
R1417 B.n560 B.n31 163.367
R1418 B.n560 B.n559 163.367
R1419 B.n559 B.n558 163.367
R1420 B.n558 B.n33 163.367
R1421 B.n554 B.n33 163.367
R1422 B.n554 B.n553 163.367
R1423 B.n553 B.n552 163.367
R1424 B.n552 B.n35 163.367
R1425 B.n548 B.n35 163.367
R1426 B.n548 B.n547 163.367
R1427 B.n547 B.n546 163.367
R1428 B.n546 B.n37 163.367
R1429 B.n542 B.n37 163.367
R1430 B.n542 B.n541 163.367
R1431 B.n541 B.n540 163.367
R1432 B.n540 B.n39 163.367
R1433 B.n535 B.n39 163.367
R1434 B.n535 B.n534 163.367
R1435 B.n534 B.n533 163.367
R1436 B.n533 B.n43 163.367
R1437 B.n529 B.n43 163.367
R1438 B.n529 B.n528 163.367
R1439 B.n528 B.n527 163.367
R1440 B.n527 B.n45 163.367
R1441 B.n523 B.n45 163.367
R1442 B.n523 B.n522 163.367
R1443 B.n522 B.n49 163.367
R1444 B.n518 B.n49 163.367
R1445 B.n518 B.n517 163.367
R1446 B.n517 B.n516 163.367
R1447 B.n516 B.n51 163.367
R1448 B.n512 B.n51 163.367
R1449 B.n512 B.n511 163.367
R1450 B.n511 B.n510 163.367
R1451 B.n510 B.n53 163.367
R1452 B.n506 B.n53 163.367
R1453 B.n506 B.n505 163.367
R1454 B.n505 B.n504 163.367
R1455 B.n504 B.n55 163.367
R1456 B.n500 B.n55 163.367
R1457 B.n500 B.n499 163.367
R1458 B.n499 B.n498 163.367
R1459 B.n498 B.n57 163.367
R1460 B.n494 B.n57 163.367
R1461 B.n494 B.n493 163.367
R1462 B.n493 B.n492 163.367
R1463 B.n492 B.n59 163.367
R1464 B.n488 B.n59 163.367
R1465 B.n488 B.n487 163.367
R1466 B.n487 B.n486 163.367
R1467 B.n486 B.n61 163.367
R1468 B.n482 B.n61 163.367
R1469 B.n482 B.n481 163.367
R1470 B.n481 B.n480 163.367
R1471 B.n480 B.n63 163.367
R1472 B.n476 B.n63 163.367
R1473 B.n476 B.n475 163.367
R1474 B.n475 B.n474 163.367
R1475 B.n474 B.n65 163.367
R1476 B.n470 B.n65 163.367
R1477 B.n470 B.n469 163.367
R1478 B.n469 B.n468 163.367
R1479 B.n468 B.n67 163.367
R1480 B.n126 B.n125 59.5399
R1481 B.n281 B.n133 59.5399
R1482 B.n537 B.n41 59.5399
R1483 B.n48 B.n47 59.5399
R1484 B.n125 B.n124 47.3217
R1485 B.n133 B.n132 47.3217
R1486 B.n41 B.n40 47.3217
R1487 B.n47 B.n46 47.3217
R1488 B.n593 B.n20 28.8785
R1489 B.n353 B.n352 28.8785
R1490 B.n225 B.n152 28.8785
R1491 B.n466 B.n465 28.8785
R1492 B B.n651 18.0485
R1493 B.n593 B.n592 10.6151
R1494 B.n592 B.n591 10.6151
R1495 B.n591 B.n22 10.6151
R1496 B.n587 B.n22 10.6151
R1497 B.n587 B.n586 10.6151
R1498 B.n586 B.n585 10.6151
R1499 B.n585 B.n24 10.6151
R1500 B.n581 B.n24 10.6151
R1501 B.n581 B.n580 10.6151
R1502 B.n580 B.n579 10.6151
R1503 B.n579 B.n26 10.6151
R1504 B.n575 B.n26 10.6151
R1505 B.n575 B.n574 10.6151
R1506 B.n574 B.n573 10.6151
R1507 B.n573 B.n28 10.6151
R1508 B.n569 B.n28 10.6151
R1509 B.n569 B.n568 10.6151
R1510 B.n568 B.n567 10.6151
R1511 B.n567 B.n30 10.6151
R1512 B.n563 B.n30 10.6151
R1513 B.n563 B.n562 10.6151
R1514 B.n562 B.n561 10.6151
R1515 B.n561 B.n32 10.6151
R1516 B.n557 B.n32 10.6151
R1517 B.n557 B.n556 10.6151
R1518 B.n556 B.n555 10.6151
R1519 B.n555 B.n34 10.6151
R1520 B.n551 B.n34 10.6151
R1521 B.n551 B.n550 10.6151
R1522 B.n550 B.n549 10.6151
R1523 B.n549 B.n36 10.6151
R1524 B.n545 B.n36 10.6151
R1525 B.n545 B.n544 10.6151
R1526 B.n544 B.n543 10.6151
R1527 B.n543 B.n38 10.6151
R1528 B.n539 B.n38 10.6151
R1529 B.n539 B.n538 10.6151
R1530 B.n536 B.n42 10.6151
R1531 B.n532 B.n42 10.6151
R1532 B.n532 B.n531 10.6151
R1533 B.n531 B.n530 10.6151
R1534 B.n530 B.n44 10.6151
R1535 B.n526 B.n44 10.6151
R1536 B.n526 B.n525 10.6151
R1537 B.n525 B.n524 10.6151
R1538 B.n521 B.n520 10.6151
R1539 B.n520 B.n519 10.6151
R1540 B.n519 B.n50 10.6151
R1541 B.n515 B.n50 10.6151
R1542 B.n515 B.n514 10.6151
R1543 B.n514 B.n513 10.6151
R1544 B.n513 B.n52 10.6151
R1545 B.n509 B.n52 10.6151
R1546 B.n509 B.n508 10.6151
R1547 B.n508 B.n507 10.6151
R1548 B.n507 B.n54 10.6151
R1549 B.n503 B.n54 10.6151
R1550 B.n503 B.n502 10.6151
R1551 B.n502 B.n501 10.6151
R1552 B.n501 B.n56 10.6151
R1553 B.n497 B.n56 10.6151
R1554 B.n497 B.n496 10.6151
R1555 B.n496 B.n495 10.6151
R1556 B.n495 B.n58 10.6151
R1557 B.n491 B.n58 10.6151
R1558 B.n491 B.n490 10.6151
R1559 B.n490 B.n489 10.6151
R1560 B.n489 B.n60 10.6151
R1561 B.n485 B.n60 10.6151
R1562 B.n485 B.n484 10.6151
R1563 B.n484 B.n483 10.6151
R1564 B.n483 B.n62 10.6151
R1565 B.n479 B.n62 10.6151
R1566 B.n479 B.n478 10.6151
R1567 B.n478 B.n477 10.6151
R1568 B.n477 B.n64 10.6151
R1569 B.n473 B.n64 10.6151
R1570 B.n473 B.n472 10.6151
R1571 B.n472 B.n471 10.6151
R1572 B.n471 B.n66 10.6151
R1573 B.n467 B.n66 10.6151
R1574 B.n467 B.n466 10.6151
R1575 B.n353 B.n104 10.6151
R1576 B.n357 B.n104 10.6151
R1577 B.n358 B.n357 10.6151
R1578 B.n359 B.n358 10.6151
R1579 B.n359 B.n102 10.6151
R1580 B.n363 B.n102 10.6151
R1581 B.n364 B.n363 10.6151
R1582 B.n365 B.n364 10.6151
R1583 B.n365 B.n100 10.6151
R1584 B.n369 B.n100 10.6151
R1585 B.n370 B.n369 10.6151
R1586 B.n371 B.n370 10.6151
R1587 B.n371 B.n98 10.6151
R1588 B.n375 B.n98 10.6151
R1589 B.n376 B.n375 10.6151
R1590 B.n377 B.n376 10.6151
R1591 B.n377 B.n96 10.6151
R1592 B.n381 B.n96 10.6151
R1593 B.n382 B.n381 10.6151
R1594 B.n383 B.n382 10.6151
R1595 B.n383 B.n94 10.6151
R1596 B.n387 B.n94 10.6151
R1597 B.n388 B.n387 10.6151
R1598 B.n389 B.n388 10.6151
R1599 B.n389 B.n92 10.6151
R1600 B.n393 B.n92 10.6151
R1601 B.n394 B.n393 10.6151
R1602 B.n395 B.n394 10.6151
R1603 B.n395 B.n90 10.6151
R1604 B.n399 B.n90 10.6151
R1605 B.n400 B.n399 10.6151
R1606 B.n401 B.n400 10.6151
R1607 B.n401 B.n88 10.6151
R1608 B.n405 B.n88 10.6151
R1609 B.n406 B.n405 10.6151
R1610 B.n407 B.n406 10.6151
R1611 B.n407 B.n86 10.6151
R1612 B.n411 B.n86 10.6151
R1613 B.n412 B.n411 10.6151
R1614 B.n413 B.n412 10.6151
R1615 B.n413 B.n84 10.6151
R1616 B.n417 B.n84 10.6151
R1617 B.n418 B.n417 10.6151
R1618 B.n419 B.n418 10.6151
R1619 B.n419 B.n82 10.6151
R1620 B.n423 B.n82 10.6151
R1621 B.n424 B.n423 10.6151
R1622 B.n425 B.n424 10.6151
R1623 B.n425 B.n80 10.6151
R1624 B.n429 B.n80 10.6151
R1625 B.n430 B.n429 10.6151
R1626 B.n431 B.n430 10.6151
R1627 B.n431 B.n78 10.6151
R1628 B.n435 B.n78 10.6151
R1629 B.n436 B.n435 10.6151
R1630 B.n437 B.n436 10.6151
R1631 B.n437 B.n76 10.6151
R1632 B.n441 B.n76 10.6151
R1633 B.n442 B.n441 10.6151
R1634 B.n443 B.n442 10.6151
R1635 B.n443 B.n74 10.6151
R1636 B.n447 B.n74 10.6151
R1637 B.n448 B.n447 10.6151
R1638 B.n449 B.n448 10.6151
R1639 B.n449 B.n72 10.6151
R1640 B.n453 B.n72 10.6151
R1641 B.n454 B.n453 10.6151
R1642 B.n455 B.n454 10.6151
R1643 B.n455 B.n70 10.6151
R1644 B.n459 B.n70 10.6151
R1645 B.n460 B.n459 10.6151
R1646 B.n461 B.n460 10.6151
R1647 B.n461 B.n68 10.6151
R1648 B.n465 B.n68 10.6151
R1649 B.n226 B.n225 10.6151
R1650 B.n227 B.n226 10.6151
R1651 B.n227 B.n150 10.6151
R1652 B.n231 B.n150 10.6151
R1653 B.n232 B.n231 10.6151
R1654 B.n233 B.n232 10.6151
R1655 B.n233 B.n148 10.6151
R1656 B.n237 B.n148 10.6151
R1657 B.n238 B.n237 10.6151
R1658 B.n239 B.n238 10.6151
R1659 B.n239 B.n146 10.6151
R1660 B.n243 B.n146 10.6151
R1661 B.n244 B.n243 10.6151
R1662 B.n245 B.n244 10.6151
R1663 B.n245 B.n144 10.6151
R1664 B.n249 B.n144 10.6151
R1665 B.n250 B.n249 10.6151
R1666 B.n251 B.n250 10.6151
R1667 B.n251 B.n142 10.6151
R1668 B.n255 B.n142 10.6151
R1669 B.n256 B.n255 10.6151
R1670 B.n257 B.n256 10.6151
R1671 B.n257 B.n140 10.6151
R1672 B.n261 B.n140 10.6151
R1673 B.n262 B.n261 10.6151
R1674 B.n263 B.n262 10.6151
R1675 B.n263 B.n138 10.6151
R1676 B.n267 B.n138 10.6151
R1677 B.n268 B.n267 10.6151
R1678 B.n269 B.n268 10.6151
R1679 B.n269 B.n136 10.6151
R1680 B.n273 B.n136 10.6151
R1681 B.n274 B.n273 10.6151
R1682 B.n275 B.n274 10.6151
R1683 B.n275 B.n134 10.6151
R1684 B.n279 B.n134 10.6151
R1685 B.n280 B.n279 10.6151
R1686 B.n282 B.n130 10.6151
R1687 B.n286 B.n130 10.6151
R1688 B.n287 B.n286 10.6151
R1689 B.n288 B.n287 10.6151
R1690 B.n288 B.n128 10.6151
R1691 B.n292 B.n128 10.6151
R1692 B.n293 B.n292 10.6151
R1693 B.n294 B.n293 10.6151
R1694 B.n298 B.n297 10.6151
R1695 B.n299 B.n298 10.6151
R1696 B.n299 B.n122 10.6151
R1697 B.n303 B.n122 10.6151
R1698 B.n304 B.n303 10.6151
R1699 B.n305 B.n304 10.6151
R1700 B.n305 B.n120 10.6151
R1701 B.n309 B.n120 10.6151
R1702 B.n310 B.n309 10.6151
R1703 B.n311 B.n310 10.6151
R1704 B.n311 B.n118 10.6151
R1705 B.n315 B.n118 10.6151
R1706 B.n316 B.n315 10.6151
R1707 B.n317 B.n316 10.6151
R1708 B.n317 B.n116 10.6151
R1709 B.n321 B.n116 10.6151
R1710 B.n322 B.n321 10.6151
R1711 B.n323 B.n322 10.6151
R1712 B.n323 B.n114 10.6151
R1713 B.n327 B.n114 10.6151
R1714 B.n328 B.n327 10.6151
R1715 B.n329 B.n328 10.6151
R1716 B.n329 B.n112 10.6151
R1717 B.n333 B.n112 10.6151
R1718 B.n334 B.n333 10.6151
R1719 B.n335 B.n334 10.6151
R1720 B.n335 B.n110 10.6151
R1721 B.n339 B.n110 10.6151
R1722 B.n340 B.n339 10.6151
R1723 B.n341 B.n340 10.6151
R1724 B.n341 B.n108 10.6151
R1725 B.n345 B.n108 10.6151
R1726 B.n346 B.n345 10.6151
R1727 B.n347 B.n346 10.6151
R1728 B.n347 B.n106 10.6151
R1729 B.n351 B.n106 10.6151
R1730 B.n352 B.n351 10.6151
R1731 B.n221 B.n152 10.6151
R1732 B.n221 B.n220 10.6151
R1733 B.n220 B.n219 10.6151
R1734 B.n219 B.n154 10.6151
R1735 B.n215 B.n154 10.6151
R1736 B.n215 B.n214 10.6151
R1737 B.n214 B.n213 10.6151
R1738 B.n213 B.n156 10.6151
R1739 B.n209 B.n156 10.6151
R1740 B.n209 B.n208 10.6151
R1741 B.n208 B.n207 10.6151
R1742 B.n207 B.n158 10.6151
R1743 B.n203 B.n158 10.6151
R1744 B.n203 B.n202 10.6151
R1745 B.n202 B.n201 10.6151
R1746 B.n201 B.n160 10.6151
R1747 B.n197 B.n160 10.6151
R1748 B.n197 B.n196 10.6151
R1749 B.n196 B.n195 10.6151
R1750 B.n195 B.n162 10.6151
R1751 B.n191 B.n162 10.6151
R1752 B.n191 B.n190 10.6151
R1753 B.n190 B.n189 10.6151
R1754 B.n189 B.n164 10.6151
R1755 B.n185 B.n164 10.6151
R1756 B.n185 B.n184 10.6151
R1757 B.n184 B.n183 10.6151
R1758 B.n183 B.n166 10.6151
R1759 B.n179 B.n166 10.6151
R1760 B.n179 B.n178 10.6151
R1761 B.n178 B.n177 10.6151
R1762 B.n177 B.n168 10.6151
R1763 B.n173 B.n168 10.6151
R1764 B.n173 B.n172 10.6151
R1765 B.n172 B.n171 10.6151
R1766 B.n171 B.n0 10.6151
R1767 B.n647 B.n1 10.6151
R1768 B.n647 B.n646 10.6151
R1769 B.n646 B.n645 10.6151
R1770 B.n645 B.n4 10.6151
R1771 B.n641 B.n4 10.6151
R1772 B.n641 B.n640 10.6151
R1773 B.n640 B.n639 10.6151
R1774 B.n639 B.n6 10.6151
R1775 B.n635 B.n6 10.6151
R1776 B.n635 B.n634 10.6151
R1777 B.n634 B.n633 10.6151
R1778 B.n633 B.n8 10.6151
R1779 B.n629 B.n8 10.6151
R1780 B.n629 B.n628 10.6151
R1781 B.n628 B.n627 10.6151
R1782 B.n627 B.n10 10.6151
R1783 B.n623 B.n10 10.6151
R1784 B.n623 B.n622 10.6151
R1785 B.n622 B.n621 10.6151
R1786 B.n621 B.n12 10.6151
R1787 B.n617 B.n12 10.6151
R1788 B.n617 B.n616 10.6151
R1789 B.n616 B.n615 10.6151
R1790 B.n615 B.n14 10.6151
R1791 B.n611 B.n14 10.6151
R1792 B.n611 B.n610 10.6151
R1793 B.n610 B.n609 10.6151
R1794 B.n609 B.n16 10.6151
R1795 B.n605 B.n16 10.6151
R1796 B.n605 B.n604 10.6151
R1797 B.n604 B.n603 10.6151
R1798 B.n603 B.n18 10.6151
R1799 B.n599 B.n18 10.6151
R1800 B.n599 B.n598 10.6151
R1801 B.n598 B.n597 10.6151
R1802 B.n597 B.n20 10.6151
R1803 B.n537 B.n536 6.5566
R1804 B.n524 B.n48 6.5566
R1805 B.n282 B.n281 6.5566
R1806 B.n294 B.n126 6.5566
R1807 B.n538 B.n537 4.05904
R1808 B.n521 B.n48 4.05904
R1809 B.n281 B.n280 4.05904
R1810 B.n297 B.n126 4.05904
R1811 B.n651 B.n0 2.81026
R1812 B.n651 B.n1 2.81026
C0 w_n2922_n3092# VTAIL 2.74602f
C1 VDD2 VN 5.73638f
C2 VDD2 VTAIL 7.21566f
C3 w_n2922_n3092# B 8.611879f
C4 VP VN 6.18937f
C5 w_n2922_n3092# VDD1 2.07739f
C6 VDD2 B 1.91779f
C7 VTAIL VP 5.85443f
C8 VTAIL VN 5.84012f
C9 VDD2 VDD1 1.21885f
C10 B VP 1.6769f
C11 B VN 1.05092f
C12 VP VDD1 5.99991f
C13 B VTAIL 3.18611f
C14 VDD1 VN 0.150477f
C15 VDD2 w_n2922_n3092# 2.14684f
C16 VTAIL VDD1 7.16834f
C17 B VDD1 1.85545f
C18 w_n2922_n3092# VP 5.75523f
C19 w_n2922_n3092# VN 5.37883f
C20 VDD2 VP 0.417087f
C21 VDD2 VSUBS 1.638532f
C22 VDD1 VSUBS 1.583763f
C23 VTAIL VSUBS 1.048337f
C24 VN VSUBS 5.32226f
C25 VP VSUBS 2.514159f
C26 B VSUBS 4.033748f
C27 w_n2922_n3092# VSUBS 0.111468p
C28 B.n0 VSUBS 0.00417f
C29 B.n1 VSUBS 0.00417f
C30 B.n2 VSUBS 0.006595f
C31 B.n3 VSUBS 0.006595f
C32 B.n4 VSUBS 0.006595f
C33 B.n5 VSUBS 0.006595f
C34 B.n6 VSUBS 0.006595f
C35 B.n7 VSUBS 0.006595f
C36 B.n8 VSUBS 0.006595f
C37 B.n9 VSUBS 0.006595f
C38 B.n10 VSUBS 0.006595f
C39 B.n11 VSUBS 0.006595f
C40 B.n12 VSUBS 0.006595f
C41 B.n13 VSUBS 0.006595f
C42 B.n14 VSUBS 0.006595f
C43 B.n15 VSUBS 0.006595f
C44 B.n16 VSUBS 0.006595f
C45 B.n17 VSUBS 0.006595f
C46 B.n18 VSUBS 0.006595f
C47 B.n19 VSUBS 0.006595f
C48 B.n20 VSUBS 0.013859f
C49 B.n21 VSUBS 0.006595f
C50 B.n22 VSUBS 0.006595f
C51 B.n23 VSUBS 0.006595f
C52 B.n24 VSUBS 0.006595f
C53 B.n25 VSUBS 0.006595f
C54 B.n26 VSUBS 0.006595f
C55 B.n27 VSUBS 0.006595f
C56 B.n28 VSUBS 0.006595f
C57 B.n29 VSUBS 0.006595f
C58 B.n30 VSUBS 0.006595f
C59 B.n31 VSUBS 0.006595f
C60 B.n32 VSUBS 0.006595f
C61 B.n33 VSUBS 0.006595f
C62 B.n34 VSUBS 0.006595f
C63 B.n35 VSUBS 0.006595f
C64 B.n36 VSUBS 0.006595f
C65 B.n37 VSUBS 0.006595f
C66 B.n38 VSUBS 0.006595f
C67 B.n39 VSUBS 0.006595f
C68 B.t8 VSUBS 0.17018f
C69 B.t7 VSUBS 0.194861f
C70 B.t6 VSUBS 0.955135f
C71 B.n40 VSUBS 0.312071f
C72 B.n41 VSUBS 0.216975f
C73 B.n42 VSUBS 0.006595f
C74 B.n43 VSUBS 0.006595f
C75 B.n44 VSUBS 0.006595f
C76 B.n45 VSUBS 0.006595f
C77 B.t5 VSUBS 0.170183f
C78 B.t4 VSUBS 0.194864f
C79 B.t3 VSUBS 0.955135f
C80 B.n46 VSUBS 0.312069f
C81 B.n47 VSUBS 0.216973f
C82 B.n48 VSUBS 0.01528f
C83 B.n49 VSUBS 0.006595f
C84 B.n50 VSUBS 0.006595f
C85 B.n51 VSUBS 0.006595f
C86 B.n52 VSUBS 0.006595f
C87 B.n53 VSUBS 0.006595f
C88 B.n54 VSUBS 0.006595f
C89 B.n55 VSUBS 0.006595f
C90 B.n56 VSUBS 0.006595f
C91 B.n57 VSUBS 0.006595f
C92 B.n58 VSUBS 0.006595f
C93 B.n59 VSUBS 0.006595f
C94 B.n60 VSUBS 0.006595f
C95 B.n61 VSUBS 0.006595f
C96 B.n62 VSUBS 0.006595f
C97 B.n63 VSUBS 0.006595f
C98 B.n64 VSUBS 0.006595f
C99 B.n65 VSUBS 0.006595f
C100 B.n66 VSUBS 0.006595f
C101 B.n67 VSUBS 0.014654f
C102 B.n68 VSUBS 0.006595f
C103 B.n69 VSUBS 0.006595f
C104 B.n70 VSUBS 0.006595f
C105 B.n71 VSUBS 0.006595f
C106 B.n72 VSUBS 0.006595f
C107 B.n73 VSUBS 0.006595f
C108 B.n74 VSUBS 0.006595f
C109 B.n75 VSUBS 0.006595f
C110 B.n76 VSUBS 0.006595f
C111 B.n77 VSUBS 0.006595f
C112 B.n78 VSUBS 0.006595f
C113 B.n79 VSUBS 0.006595f
C114 B.n80 VSUBS 0.006595f
C115 B.n81 VSUBS 0.006595f
C116 B.n82 VSUBS 0.006595f
C117 B.n83 VSUBS 0.006595f
C118 B.n84 VSUBS 0.006595f
C119 B.n85 VSUBS 0.006595f
C120 B.n86 VSUBS 0.006595f
C121 B.n87 VSUBS 0.006595f
C122 B.n88 VSUBS 0.006595f
C123 B.n89 VSUBS 0.006595f
C124 B.n90 VSUBS 0.006595f
C125 B.n91 VSUBS 0.006595f
C126 B.n92 VSUBS 0.006595f
C127 B.n93 VSUBS 0.006595f
C128 B.n94 VSUBS 0.006595f
C129 B.n95 VSUBS 0.006595f
C130 B.n96 VSUBS 0.006595f
C131 B.n97 VSUBS 0.006595f
C132 B.n98 VSUBS 0.006595f
C133 B.n99 VSUBS 0.006595f
C134 B.n100 VSUBS 0.006595f
C135 B.n101 VSUBS 0.006595f
C136 B.n102 VSUBS 0.006595f
C137 B.n103 VSUBS 0.006595f
C138 B.n104 VSUBS 0.006595f
C139 B.n105 VSUBS 0.014654f
C140 B.n106 VSUBS 0.006595f
C141 B.n107 VSUBS 0.006595f
C142 B.n108 VSUBS 0.006595f
C143 B.n109 VSUBS 0.006595f
C144 B.n110 VSUBS 0.006595f
C145 B.n111 VSUBS 0.006595f
C146 B.n112 VSUBS 0.006595f
C147 B.n113 VSUBS 0.006595f
C148 B.n114 VSUBS 0.006595f
C149 B.n115 VSUBS 0.006595f
C150 B.n116 VSUBS 0.006595f
C151 B.n117 VSUBS 0.006595f
C152 B.n118 VSUBS 0.006595f
C153 B.n119 VSUBS 0.006595f
C154 B.n120 VSUBS 0.006595f
C155 B.n121 VSUBS 0.006595f
C156 B.n122 VSUBS 0.006595f
C157 B.n123 VSUBS 0.006595f
C158 B.t1 VSUBS 0.170183f
C159 B.t2 VSUBS 0.194864f
C160 B.t0 VSUBS 0.955135f
C161 B.n124 VSUBS 0.312069f
C162 B.n125 VSUBS 0.216973f
C163 B.n126 VSUBS 0.01528f
C164 B.n127 VSUBS 0.006595f
C165 B.n128 VSUBS 0.006595f
C166 B.n129 VSUBS 0.006595f
C167 B.n130 VSUBS 0.006595f
C168 B.n131 VSUBS 0.006595f
C169 B.t10 VSUBS 0.17018f
C170 B.t11 VSUBS 0.194861f
C171 B.t9 VSUBS 0.955135f
C172 B.n132 VSUBS 0.312071f
C173 B.n133 VSUBS 0.216975f
C174 B.n134 VSUBS 0.006595f
C175 B.n135 VSUBS 0.006595f
C176 B.n136 VSUBS 0.006595f
C177 B.n137 VSUBS 0.006595f
C178 B.n138 VSUBS 0.006595f
C179 B.n139 VSUBS 0.006595f
C180 B.n140 VSUBS 0.006595f
C181 B.n141 VSUBS 0.006595f
C182 B.n142 VSUBS 0.006595f
C183 B.n143 VSUBS 0.006595f
C184 B.n144 VSUBS 0.006595f
C185 B.n145 VSUBS 0.006595f
C186 B.n146 VSUBS 0.006595f
C187 B.n147 VSUBS 0.006595f
C188 B.n148 VSUBS 0.006595f
C189 B.n149 VSUBS 0.006595f
C190 B.n150 VSUBS 0.006595f
C191 B.n151 VSUBS 0.006595f
C192 B.n152 VSUBS 0.013859f
C193 B.n153 VSUBS 0.006595f
C194 B.n154 VSUBS 0.006595f
C195 B.n155 VSUBS 0.006595f
C196 B.n156 VSUBS 0.006595f
C197 B.n157 VSUBS 0.006595f
C198 B.n158 VSUBS 0.006595f
C199 B.n159 VSUBS 0.006595f
C200 B.n160 VSUBS 0.006595f
C201 B.n161 VSUBS 0.006595f
C202 B.n162 VSUBS 0.006595f
C203 B.n163 VSUBS 0.006595f
C204 B.n164 VSUBS 0.006595f
C205 B.n165 VSUBS 0.006595f
C206 B.n166 VSUBS 0.006595f
C207 B.n167 VSUBS 0.006595f
C208 B.n168 VSUBS 0.006595f
C209 B.n169 VSUBS 0.006595f
C210 B.n170 VSUBS 0.006595f
C211 B.n171 VSUBS 0.006595f
C212 B.n172 VSUBS 0.006595f
C213 B.n173 VSUBS 0.006595f
C214 B.n174 VSUBS 0.006595f
C215 B.n175 VSUBS 0.006595f
C216 B.n176 VSUBS 0.006595f
C217 B.n177 VSUBS 0.006595f
C218 B.n178 VSUBS 0.006595f
C219 B.n179 VSUBS 0.006595f
C220 B.n180 VSUBS 0.006595f
C221 B.n181 VSUBS 0.006595f
C222 B.n182 VSUBS 0.006595f
C223 B.n183 VSUBS 0.006595f
C224 B.n184 VSUBS 0.006595f
C225 B.n185 VSUBS 0.006595f
C226 B.n186 VSUBS 0.006595f
C227 B.n187 VSUBS 0.006595f
C228 B.n188 VSUBS 0.006595f
C229 B.n189 VSUBS 0.006595f
C230 B.n190 VSUBS 0.006595f
C231 B.n191 VSUBS 0.006595f
C232 B.n192 VSUBS 0.006595f
C233 B.n193 VSUBS 0.006595f
C234 B.n194 VSUBS 0.006595f
C235 B.n195 VSUBS 0.006595f
C236 B.n196 VSUBS 0.006595f
C237 B.n197 VSUBS 0.006595f
C238 B.n198 VSUBS 0.006595f
C239 B.n199 VSUBS 0.006595f
C240 B.n200 VSUBS 0.006595f
C241 B.n201 VSUBS 0.006595f
C242 B.n202 VSUBS 0.006595f
C243 B.n203 VSUBS 0.006595f
C244 B.n204 VSUBS 0.006595f
C245 B.n205 VSUBS 0.006595f
C246 B.n206 VSUBS 0.006595f
C247 B.n207 VSUBS 0.006595f
C248 B.n208 VSUBS 0.006595f
C249 B.n209 VSUBS 0.006595f
C250 B.n210 VSUBS 0.006595f
C251 B.n211 VSUBS 0.006595f
C252 B.n212 VSUBS 0.006595f
C253 B.n213 VSUBS 0.006595f
C254 B.n214 VSUBS 0.006595f
C255 B.n215 VSUBS 0.006595f
C256 B.n216 VSUBS 0.006595f
C257 B.n217 VSUBS 0.006595f
C258 B.n218 VSUBS 0.006595f
C259 B.n219 VSUBS 0.006595f
C260 B.n220 VSUBS 0.006595f
C261 B.n221 VSUBS 0.006595f
C262 B.n222 VSUBS 0.006595f
C263 B.n223 VSUBS 0.013859f
C264 B.n224 VSUBS 0.014654f
C265 B.n225 VSUBS 0.014654f
C266 B.n226 VSUBS 0.006595f
C267 B.n227 VSUBS 0.006595f
C268 B.n228 VSUBS 0.006595f
C269 B.n229 VSUBS 0.006595f
C270 B.n230 VSUBS 0.006595f
C271 B.n231 VSUBS 0.006595f
C272 B.n232 VSUBS 0.006595f
C273 B.n233 VSUBS 0.006595f
C274 B.n234 VSUBS 0.006595f
C275 B.n235 VSUBS 0.006595f
C276 B.n236 VSUBS 0.006595f
C277 B.n237 VSUBS 0.006595f
C278 B.n238 VSUBS 0.006595f
C279 B.n239 VSUBS 0.006595f
C280 B.n240 VSUBS 0.006595f
C281 B.n241 VSUBS 0.006595f
C282 B.n242 VSUBS 0.006595f
C283 B.n243 VSUBS 0.006595f
C284 B.n244 VSUBS 0.006595f
C285 B.n245 VSUBS 0.006595f
C286 B.n246 VSUBS 0.006595f
C287 B.n247 VSUBS 0.006595f
C288 B.n248 VSUBS 0.006595f
C289 B.n249 VSUBS 0.006595f
C290 B.n250 VSUBS 0.006595f
C291 B.n251 VSUBS 0.006595f
C292 B.n252 VSUBS 0.006595f
C293 B.n253 VSUBS 0.006595f
C294 B.n254 VSUBS 0.006595f
C295 B.n255 VSUBS 0.006595f
C296 B.n256 VSUBS 0.006595f
C297 B.n257 VSUBS 0.006595f
C298 B.n258 VSUBS 0.006595f
C299 B.n259 VSUBS 0.006595f
C300 B.n260 VSUBS 0.006595f
C301 B.n261 VSUBS 0.006595f
C302 B.n262 VSUBS 0.006595f
C303 B.n263 VSUBS 0.006595f
C304 B.n264 VSUBS 0.006595f
C305 B.n265 VSUBS 0.006595f
C306 B.n266 VSUBS 0.006595f
C307 B.n267 VSUBS 0.006595f
C308 B.n268 VSUBS 0.006595f
C309 B.n269 VSUBS 0.006595f
C310 B.n270 VSUBS 0.006595f
C311 B.n271 VSUBS 0.006595f
C312 B.n272 VSUBS 0.006595f
C313 B.n273 VSUBS 0.006595f
C314 B.n274 VSUBS 0.006595f
C315 B.n275 VSUBS 0.006595f
C316 B.n276 VSUBS 0.006595f
C317 B.n277 VSUBS 0.006595f
C318 B.n278 VSUBS 0.006595f
C319 B.n279 VSUBS 0.006595f
C320 B.n280 VSUBS 0.004558f
C321 B.n281 VSUBS 0.01528f
C322 B.n282 VSUBS 0.005334f
C323 B.n283 VSUBS 0.006595f
C324 B.n284 VSUBS 0.006595f
C325 B.n285 VSUBS 0.006595f
C326 B.n286 VSUBS 0.006595f
C327 B.n287 VSUBS 0.006595f
C328 B.n288 VSUBS 0.006595f
C329 B.n289 VSUBS 0.006595f
C330 B.n290 VSUBS 0.006595f
C331 B.n291 VSUBS 0.006595f
C332 B.n292 VSUBS 0.006595f
C333 B.n293 VSUBS 0.006595f
C334 B.n294 VSUBS 0.005334f
C335 B.n295 VSUBS 0.006595f
C336 B.n296 VSUBS 0.006595f
C337 B.n297 VSUBS 0.004558f
C338 B.n298 VSUBS 0.006595f
C339 B.n299 VSUBS 0.006595f
C340 B.n300 VSUBS 0.006595f
C341 B.n301 VSUBS 0.006595f
C342 B.n302 VSUBS 0.006595f
C343 B.n303 VSUBS 0.006595f
C344 B.n304 VSUBS 0.006595f
C345 B.n305 VSUBS 0.006595f
C346 B.n306 VSUBS 0.006595f
C347 B.n307 VSUBS 0.006595f
C348 B.n308 VSUBS 0.006595f
C349 B.n309 VSUBS 0.006595f
C350 B.n310 VSUBS 0.006595f
C351 B.n311 VSUBS 0.006595f
C352 B.n312 VSUBS 0.006595f
C353 B.n313 VSUBS 0.006595f
C354 B.n314 VSUBS 0.006595f
C355 B.n315 VSUBS 0.006595f
C356 B.n316 VSUBS 0.006595f
C357 B.n317 VSUBS 0.006595f
C358 B.n318 VSUBS 0.006595f
C359 B.n319 VSUBS 0.006595f
C360 B.n320 VSUBS 0.006595f
C361 B.n321 VSUBS 0.006595f
C362 B.n322 VSUBS 0.006595f
C363 B.n323 VSUBS 0.006595f
C364 B.n324 VSUBS 0.006595f
C365 B.n325 VSUBS 0.006595f
C366 B.n326 VSUBS 0.006595f
C367 B.n327 VSUBS 0.006595f
C368 B.n328 VSUBS 0.006595f
C369 B.n329 VSUBS 0.006595f
C370 B.n330 VSUBS 0.006595f
C371 B.n331 VSUBS 0.006595f
C372 B.n332 VSUBS 0.006595f
C373 B.n333 VSUBS 0.006595f
C374 B.n334 VSUBS 0.006595f
C375 B.n335 VSUBS 0.006595f
C376 B.n336 VSUBS 0.006595f
C377 B.n337 VSUBS 0.006595f
C378 B.n338 VSUBS 0.006595f
C379 B.n339 VSUBS 0.006595f
C380 B.n340 VSUBS 0.006595f
C381 B.n341 VSUBS 0.006595f
C382 B.n342 VSUBS 0.006595f
C383 B.n343 VSUBS 0.006595f
C384 B.n344 VSUBS 0.006595f
C385 B.n345 VSUBS 0.006595f
C386 B.n346 VSUBS 0.006595f
C387 B.n347 VSUBS 0.006595f
C388 B.n348 VSUBS 0.006595f
C389 B.n349 VSUBS 0.006595f
C390 B.n350 VSUBS 0.006595f
C391 B.n351 VSUBS 0.006595f
C392 B.n352 VSUBS 0.014654f
C393 B.n353 VSUBS 0.013859f
C394 B.n354 VSUBS 0.013859f
C395 B.n355 VSUBS 0.006595f
C396 B.n356 VSUBS 0.006595f
C397 B.n357 VSUBS 0.006595f
C398 B.n358 VSUBS 0.006595f
C399 B.n359 VSUBS 0.006595f
C400 B.n360 VSUBS 0.006595f
C401 B.n361 VSUBS 0.006595f
C402 B.n362 VSUBS 0.006595f
C403 B.n363 VSUBS 0.006595f
C404 B.n364 VSUBS 0.006595f
C405 B.n365 VSUBS 0.006595f
C406 B.n366 VSUBS 0.006595f
C407 B.n367 VSUBS 0.006595f
C408 B.n368 VSUBS 0.006595f
C409 B.n369 VSUBS 0.006595f
C410 B.n370 VSUBS 0.006595f
C411 B.n371 VSUBS 0.006595f
C412 B.n372 VSUBS 0.006595f
C413 B.n373 VSUBS 0.006595f
C414 B.n374 VSUBS 0.006595f
C415 B.n375 VSUBS 0.006595f
C416 B.n376 VSUBS 0.006595f
C417 B.n377 VSUBS 0.006595f
C418 B.n378 VSUBS 0.006595f
C419 B.n379 VSUBS 0.006595f
C420 B.n380 VSUBS 0.006595f
C421 B.n381 VSUBS 0.006595f
C422 B.n382 VSUBS 0.006595f
C423 B.n383 VSUBS 0.006595f
C424 B.n384 VSUBS 0.006595f
C425 B.n385 VSUBS 0.006595f
C426 B.n386 VSUBS 0.006595f
C427 B.n387 VSUBS 0.006595f
C428 B.n388 VSUBS 0.006595f
C429 B.n389 VSUBS 0.006595f
C430 B.n390 VSUBS 0.006595f
C431 B.n391 VSUBS 0.006595f
C432 B.n392 VSUBS 0.006595f
C433 B.n393 VSUBS 0.006595f
C434 B.n394 VSUBS 0.006595f
C435 B.n395 VSUBS 0.006595f
C436 B.n396 VSUBS 0.006595f
C437 B.n397 VSUBS 0.006595f
C438 B.n398 VSUBS 0.006595f
C439 B.n399 VSUBS 0.006595f
C440 B.n400 VSUBS 0.006595f
C441 B.n401 VSUBS 0.006595f
C442 B.n402 VSUBS 0.006595f
C443 B.n403 VSUBS 0.006595f
C444 B.n404 VSUBS 0.006595f
C445 B.n405 VSUBS 0.006595f
C446 B.n406 VSUBS 0.006595f
C447 B.n407 VSUBS 0.006595f
C448 B.n408 VSUBS 0.006595f
C449 B.n409 VSUBS 0.006595f
C450 B.n410 VSUBS 0.006595f
C451 B.n411 VSUBS 0.006595f
C452 B.n412 VSUBS 0.006595f
C453 B.n413 VSUBS 0.006595f
C454 B.n414 VSUBS 0.006595f
C455 B.n415 VSUBS 0.006595f
C456 B.n416 VSUBS 0.006595f
C457 B.n417 VSUBS 0.006595f
C458 B.n418 VSUBS 0.006595f
C459 B.n419 VSUBS 0.006595f
C460 B.n420 VSUBS 0.006595f
C461 B.n421 VSUBS 0.006595f
C462 B.n422 VSUBS 0.006595f
C463 B.n423 VSUBS 0.006595f
C464 B.n424 VSUBS 0.006595f
C465 B.n425 VSUBS 0.006595f
C466 B.n426 VSUBS 0.006595f
C467 B.n427 VSUBS 0.006595f
C468 B.n428 VSUBS 0.006595f
C469 B.n429 VSUBS 0.006595f
C470 B.n430 VSUBS 0.006595f
C471 B.n431 VSUBS 0.006595f
C472 B.n432 VSUBS 0.006595f
C473 B.n433 VSUBS 0.006595f
C474 B.n434 VSUBS 0.006595f
C475 B.n435 VSUBS 0.006595f
C476 B.n436 VSUBS 0.006595f
C477 B.n437 VSUBS 0.006595f
C478 B.n438 VSUBS 0.006595f
C479 B.n439 VSUBS 0.006595f
C480 B.n440 VSUBS 0.006595f
C481 B.n441 VSUBS 0.006595f
C482 B.n442 VSUBS 0.006595f
C483 B.n443 VSUBS 0.006595f
C484 B.n444 VSUBS 0.006595f
C485 B.n445 VSUBS 0.006595f
C486 B.n446 VSUBS 0.006595f
C487 B.n447 VSUBS 0.006595f
C488 B.n448 VSUBS 0.006595f
C489 B.n449 VSUBS 0.006595f
C490 B.n450 VSUBS 0.006595f
C491 B.n451 VSUBS 0.006595f
C492 B.n452 VSUBS 0.006595f
C493 B.n453 VSUBS 0.006595f
C494 B.n454 VSUBS 0.006595f
C495 B.n455 VSUBS 0.006595f
C496 B.n456 VSUBS 0.006595f
C497 B.n457 VSUBS 0.006595f
C498 B.n458 VSUBS 0.006595f
C499 B.n459 VSUBS 0.006595f
C500 B.n460 VSUBS 0.006595f
C501 B.n461 VSUBS 0.006595f
C502 B.n462 VSUBS 0.006595f
C503 B.n463 VSUBS 0.006595f
C504 B.n464 VSUBS 0.013859f
C505 B.n465 VSUBS 0.01474f
C506 B.n466 VSUBS 0.013773f
C507 B.n467 VSUBS 0.006595f
C508 B.n468 VSUBS 0.006595f
C509 B.n469 VSUBS 0.006595f
C510 B.n470 VSUBS 0.006595f
C511 B.n471 VSUBS 0.006595f
C512 B.n472 VSUBS 0.006595f
C513 B.n473 VSUBS 0.006595f
C514 B.n474 VSUBS 0.006595f
C515 B.n475 VSUBS 0.006595f
C516 B.n476 VSUBS 0.006595f
C517 B.n477 VSUBS 0.006595f
C518 B.n478 VSUBS 0.006595f
C519 B.n479 VSUBS 0.006595f
C520 B.n480 VSUBS 0.006595f
C521 B.n481 VSUBS 0.006595f
C522 B.n482 VSUBS 0.006595f
C523 B.n483 VSUBS 0.006595f
C524 B.n484 VSUBS 0.006595f
C525 B.n485 VSUBS 0.006595f
C526 B.n486 VSUBS 0.006595f
C527 B.n487 VSUBS 0.006595f
C528 B.n488 VSUBS 0.006595f
C529 B.n489 VSUBS 0.006595f
C530 B.n490 VSUBS 0.006595f
C531 B.n491 VSUBS 0.006595f
C532 B.n492 VSUBS 0.006595f
C533 B.n493 VSUBS 0.006595f
C534 B.n494 VSUBS 0.006595f
C535 B.n495 VSUBS 0.006595f
C536 B.n496 VSUBS 0.006595f
C537 B.n497 VSUBS 0.006595f
C538 B.n498 VSUBS 0.006595f
C539 B.n499 VSUBS 0.006595f
C540 B.n500 VSUBS 0.006595f
C541 B.n501 VSUBS 0.006595f
C542 B.n502 VSUBS 0.006595f
C543 B.n503 VSUBS 0.006595f
C544 B.n504 VSUBS 0.006595f
C545 B.n505 VSUBS 0.006595f
C546 B.n506 VSUBS 0.006595f
C547 B.n507 VSUBS 0.006595f
C548 B.n508 VSUBS 0.006595f
C549 B.n509 VSUBS 0.006595f
C550 B.n510 VSUBS 0.006595f
C551 B.n511 VSUBS 0.006595f
C552 B.n512 VSUBS 0.006595f
C553 B.n513 VSUBS 0.006595f
C554 B.n514 VSUBS 0.006595f
C555 B.n515 VSUBS 0.006595f
C556 B.n516 VSUBS 0.006595f
C557 B.n517 VSUBS 0.006595f
C558 B.n518 VSUBS 0.006595f
C559 B.n519 VSUBS 0.006595f
C560 B.n520 VSUBS 0.006595f
C561 B.n521 VSUBS 0.004558f
C562 B.n522 VSUBS 0.006595f
C563 B.n523 VSUBS 0.006595f
C564 B.n524 VSUBS 0.005334f
C565 B.n525 VSUBS 0.006595f
C566 B.n526 VSUBS 0.006595f
C567 B.n527 VSUBS 0.006595f
C568 B.n528 VSUBS 0.006595f
C569 B.n529 VSUBS 0.006595f
C570 B.n530 VSUBS 0.006595f
C571 B.n531 VSUBS 0.006595f
C572 B.n532 VSUBS 0.006595f
C573 B.n533 VSUBS 0.006595f
C574 B.n534 VSUBS 0.006595f
C575 B.n535 VSUBS 0.006595f
C576 B.n536 VSUBS 0.005334f
C577 B.n537 VSUBS 0.01528f
C578 B.n538 VSUBS 0.004558f
C579 B.n539 VSUBS 0.006595f
C580 B.n540 VSUBS 0.006595f
C581 B.n541 VSUBS 0.006595f
C582 B.n542 VSUBS 0.006595f
C583 B.n543 VSUBS 0.006595f
C584 B.n544 VSUBS 0.006595f
C585 B.n545 VSUBS 0.006595f
C586 B.n546 VSUBS 0.006595f
C587 B.n547 VSUBS 0.006595f
C588 B.n548 VSUBS 0.006595f
C589 B.n549 VSUBS 0.006595f
C590 B.n550 VSUBS 0.006595f
C591 B.n551 VSUBS 0.006595f
C592 B.n552 VSUBS 0.006595f
C593 B.n553 VSUBS 0.006595f
C594 B.n554 VSUBS 0.006595f
C595 B.n555 VSUBS 0.006595f
C596 B.n556 VSUBS 0.006595f
C597 B.n557 VSUBS 0.006595f
C598 B.n558 VSUBS 0.006595f
C599 B.n559 VSUBS 0.006595f
C600 B.n560 VSUBS 0.006595f
C601 B.n561 VSUBS 0.006595f
C602 B.n562 VSUBS 0.006595f
C603 B.n563 VSUBS 0.006595f
C604 B.n564 VSUBS 0.006595f
C605 B.n565 VSUBS 0.006595f
C606 B.n566 VSUBS 0.006595f
C607 B.n567 VSUBS 0.006595f
C608 B.n568 VSUBS 0.006595f
C609 B.n569 VSUBS 0.006595f
C610 B.n570 VSUBS 0.006595f
C611 B.n571 VSUBS 0.006595f
C612 B.n572 VSUBS 0.006595f
C613 B.n573 VSUBS 0.006595f
C614 B.n574 VSUBS 0.006595f
C615 B.n575 VSUBS 0.006595f
C616 B.n576 VSUBS 0.006595f
C617 B.n577 VSUBS 0.006595f
C618 B.n578 VSUBS 0.006595f
C619 B.n579 VSUBS 0.006595f
C620 B.n580 VSUBS 0.006595f
C621 B.n581 VSUBS 0.006595f
C622 B.n582 VSUBS 0.006595f
C623 B.n583 VSUBS 0.006595f
C624 B.n584 VSUBS 0.006595f
C625 B.n585 VSUBS 0.006595f
C626 B.n586 VSUBS 0.006595f
C627 B.n587 VSUBS 0.006595f
C628 B.n588 VSUBS 0.006595f
C629 B.n589 VSUBS 0.006595f
C630 B.n590 VSUBS 0.006595f
C631 B.n591 VSUBS 0.006595f
C632 B.n592 VSUBS 0.006595f
C633 B.n593 VSUBS 0.014654f
C634 B.n594 VSUBS 0.014654f
C635 B.n595 VSUBS 0.013859f
C636 B.n596 VSUBS 0.006595f
C637 B.n597 VSUBS 0.006595f
C638 B.n598 VSUBS 0.006595f
C639 B.n599 VSUBS 0.006595f
C640 B.n600 VSUBS 0.006595f
C641 B.n601 VSUBS 0.006595f
C642 B.n602 VSUBS 0.006595f
C643 B.n603 VSUBS 0.006595f
C644 B.n604 VSUBS 0.006595f
C645 B.n605 VSUBS 0.006595f
C646 B.n606 VSUBS 0.006595f
C647 B.n607 VSUBS 0.006595f
C648 B.n608 VSUBS 0.006595f
C649 B.n609 VSUBS 0.006595f
C650 B.n610 VSUBS 0.006595f
C651 B.n611 VSUBS 0.006595f
C652 B.n612 VSUBS 0.006595f
C653 B.n613 VSUBS 0.006595f
C654 B.n614 VSUBS 0.006595f
C655 B.n615 VSUBS 0.006595f
C656 B.n616 VSUBS 0.006595f
C657 B.n617 VSUBS 0.006595f
C658 B.n618 VSUBS 0.006595f
C659 B.n619 VSUBS 0.006595f
C660 B.n620 VSUBS 0.006595f
C661 B.n621 VSUBS 0.006595f
C662 B.n622 VSUBS 0.006595f
C663 B.n623 VSUBS 0.006595f
C664 B.n624 VSUBS 0.006595f
C665 B.n625 VSUBS 0.006595f
C666 B.n626 VSUBS 0.006595f
C667 B.n627 VSUBS 0.006595f
C668 B.n628 VSUBS 0.006595f
C669 B.n629 VSUBS 0.006595f
C670 B.n630 VSUBS 0.006595f
C671 B.n631 VSUBS 0.006595f
C672 B.n632 VSUBS 0.006595f
C673 B.n633 VSUBS 0.006595f
C674 B.n634 VSUBS 0.006595f
C675 B.n635 VSUBS 0.006595f
C676 B.n636 VSUBS 0.006595f
C677 B.n637 VSUBS 0.006595f
C678 B.n638 VSUBS 0.006595f
C679 B.n639 VSUBS 0.006595f
C680 B.n640 VSUBS 0.006595f
C681 B.n641 VSUBS 0.006595f
C682 B.n642 VSUBS 0.006595f
C683 B.n643 VSUBS 0.006595f
C684 B.n644 VSUBS 0.006595f
C685 B.n645 VSUBS 0.006595f
C686 B.n646 VSUBS 0.006595f
C687 B.n647 VSUBS 0.006595f
C688 B.n648 VSUBS 0.006595f
C689 B.n649 VSUBS 0.006595f
C690 B.n650 VSUBS 0.006595f
C691 B.n651 VSUBS 0.014933f
C692 VDD1.n0 VSUBS 0.026171f
C693 VDD1.n1 VSUBS 0.02528f
C694 VDD1.n2 VSUBS 0.013584f
C695 VDD1.n3 VSUBS 0.032108f
C696 VDD1.n4 VSUBS 0.014383f
C697 VDD1.n5 VSUBS 0.02528f
C698 VDD1.n6 VSUBS 0.013584f
C699 VDD1.n7 VSUBS 0.032108f
C700 VDD1.n8 VSUBS 0.014383f
C701 VDD1.n9 VSUBS 0.02528f
C702 VDD1.n10 VSUBS 0.013584f
C703 VDD1.n11 VSUBS 0.032108f
C704 VDD1.n12 VSUBS 0.032108f
C705 VDD1.n13 VSUBS 0.014383f
C706 VDD1.n14 VSUBS 0.02528f
C707 VDD1.n15 VSUBS 0.013584f
C708 VDD1.n16 VSUBS 0.032108f
C709 VDD1.n17 VSUBS 0.014383f
C710 VDD1.n18 VSUBS 0.183323f
C711 VDD1.t0 VSUBS 0.069078f
C712 VDD1.n19 VSUBS 0.024081f
C713 VDD1.n20 VSUBS 0.024153f
C714 VDD1.n21 VSUBS 0.013584f
C715 VDD1.n22 VSUBS 1.0892f
C716 VDD1.n23 VSUBS 0.02528f
C717 VDD1.n24 VSUBS 0.013584f
C718 VDD1.n25 VSUBS 0.014383f
C719 VDD1.n26 VSUBS 0.032108f
C720 VDD1.n27 VSUBS 0.032108f
C721 VDD1.n28 VSUBS 0.014383f
C722 VDD1.n29 VSUBS 0.013584f
C723 VDD1.n30 VSUBS 0.02528f
C724 VDD1.n31 VSUBS 0.02528f
C725 VDD1.n32 VSUBS 0.013584f
C726 VDD1.n33 VSUBS 0.014383f
C727 VDD1.n34 VSUBS 0.032108f
C728 VDD1.n35 VSUBS 0.032108f
C729 VDD1.n36 VSUBS 0.014383f
C730 VDD1.n37 VSUBS 0.013584f
C731 VDD1.n38 VSUBS 0.02528f
C732 VDD1.n39 VSUBS 0.02528f
C733 VDD1.n40 VSUBS 0.013584f
C734 VDD1.n41 VSUBS 0.013984f
C735 VDD1.n42 VSUBS 0.013984f
C736 VDD1.n43 VSUBS 0.032108f
C737 VDD1.n44 VSUBS 0.032108f
C738 VDD1.n45 VSUBS 0.014383f
C739 VDD1.n46 VSUBS 0.013584f
C740 VDD1.n47 VSUBS 0.02528f
C741 VDD1.n48 VSUBS 0.02528f
C742 VDD1.n49 VSUBS 0.013584f
C743 VDD1.n50 VSUBS 0.014383f
C744 VDD1.n51 VSUBS 0.032108f
C745 VDD1.n52 VSUBS 0.07226f
C746 VDD1.n53 VSUBS 0.014383f
C747 VDD1.n54 VSUBS 0.013584f
C748 VDD1.n55 VSUBS 0.05636f
C749 VDD1.n56 VSUBS 0.059496f
C750 VDD1.n57 VSUBS 0.026171f
C751 VDD1.n58 VSUBS 0.02528f
C752 VDD1.n59 VSUBS 0.013584f
C753 VDD1.n60 VSUBS 0.032108f
C754 VDD1.n61 VSUBS 0.014383f
C755 VDD1.n62 VSUBS 0.02528f
C756 VDD1.n63 VSUBS 0.013584f
C757 VDD1.n64 VSUBS 0.032108f
C758 VDD1.n65 VSUBS 0.014383f
C759 VDD1.n66 VSUBS 0.02528f
C760 VDD1.n67 VSUBS 0.013584f
C761 VDD1.n68 VSUBS 0.032108f
C762 VDD1.n69 VSUBS 0.014383f
C763 VDD1.n70 VSUBS 0.02528f
C764 VDD1.n71 VSUBS 0.013584f
C765 VDD1.n72 VSUBS 0.032108f
C766 VDD1.n73 VSUBS 0.014383f
C767 VDD1.n74 VSUBS 0.183323f
C768 VDD1.t5 VSUBS 0.069078f
C769 VDD1.n75 VSUBS 0.024081f
C770 VDD1.n76 VSUBS 0.024153f
C771 VDD1.n77 VSUBS 0.013584f
C772 VDD1.n78 VSUBS 1.0892f
C773 VDD1.n79 VSUBS 0.02528f
C774 VDD1.n80 VSUBS 0.013584f
C775 VDD1.n81 VSUBS 0.014383f
C776 VDD1.n82 VSUBS 0.032108f
C777 VDD1.n83 VSUBS 0.032108f
C778 VDD1.n84 VSUBS 0.014383f
C779 VDD1.n85 VSUBS 0.013584f
C780 VDD1.n86 VSUBS 0.02528f
C781 VDD1.n87 VSUBS 0.02528f
C782 VDD1.n88 VSUBS 0.013584f
C783 VDD1.n89 VSUBS 0.014383f
C784 VDD1.n90 VSUBS 0.032108f
C785 VDD1.n91 VSUBS 0.032108f
C786 VDD1.n92 VSUBS 0.032108f
C787 VDD1.n93 VSUBS 0.014383f
C788 VDD1.n94 VSUBS 0.013584f
C789 VDD1.n95 VSUBS 0.02528f
C790 VDD1.n96 VSUBS 0.02528f
C791 VDD1.n97 VSUBS 0.013584f
C792 VDD1.n98 VSUBS 0.013984f
C793 VDD1.n99 VSUBS 0.013984f
C794 VDD1.n100 VSUBS 0.032108f
C795 VDD1.n101 VSUBS 0.032108f
C796 VDD1.n102 VSUBS 0.014383f
C797 VDD1.n103 VSUBS 0.013584f
C798 VDD1.n104 VSUBS 0.02528f
C799 VDD1.n105 VSUBS 0.02528f
C800 VDD1.n106 VSUBS 0.013584f
C801 VDD1.n107 VSUBS 0.014383f
C802 VDD1.n108 VSUBS 0.032108f
C803 VDD1.n109 VSUBS 0.07226f
C804 VDD1.n110 VSUBS 0.014383f
C805 VDD1.n111 VSUBS 0.013584f
C806 VDD1.n112 VSUBS 0.05636f
C807 VDD1.n113 VSUBS 0.058819f
C808 VDD1.t1 VSUBS 0.212152f
C809 VDD1.t3 VSUBS 0.212152f
C810 VDD1.n114 VSUBS 1.62027f
C811 VDD1.n115 VSUBS 2.77645f
C812 VDD1.t4 VSUBS 0.212152f
C813 VDD1.t2 VSUBS 0.212152f
C814 VDD1.n116 VSUBS 1.61596f
C815 VDD1.n117 VSUBS 2.83278f
C816 VP.n0 VSUBS 0.047823f
C817 VP.t2 VSUBS 2.20657f
C818 VP.n1 VSUBS 0.049722f
C819 VP.n2 VSUBS 0.036276f
C820 VP.t4 VSUBS 2.20657f
C821 VP.n3 VSUBS 0.049722f
C822 VP.n4 VSUBS 0.047823f
C823 VP.t0 VSUBS 2.20657f
C824 VP.n5 VSUBS 0.047823f
C825 VP.t3 VSUBS 2.20657f
C826 VP.n6 VSUBS 0.049722f
C827 VP.t5 VSUBS 2.42569f
C828 VP.n7 VSUBS 0.868329f
C829 VP.t1 VSUBS 2.20657f
C830 VP.n8 VSUBS 0.901394f
C831 VP.n9 VSUBS 0.067271f
C832 VP.n10 VSUBS 0.305397f
C833 VP.n11 VSUBS 0.036276f
C834 VP.n12 VSUBS 0.036276f
C835 VP.n13 VSUBS 0.055744f
C836 VP.n14 VSUBS 0.063285f
C837 VP.n15 VSUBS 0.913103f
C838 VP.n16 VSUBS 1.75227f
C839 VP.n17 VSUBS 1.78083f
C840 VP.n18 VSUBS 0.913103f
C841 VP.n19 VSUBS 0.063285f
C842 VP.n20 VSUBS 0.055744f
C843 VP.n21 VSUBS 0.036276f
C844 VP.n22 VSUBS 0.036276f
C845 VP.n23 VSUBS 0.036276f
C846 VP.n24 VSUBS 0.067271f
C847 VP.n25 VSUBS 0.826628f
C848 VP.n26 VSUBS 0.067271f
C849 VP.n27 VSUBS 0.036276f
C850 VP.n28 VSUBS 0.036276f
C851 VP.n29 VSUBS 0.036276f
C852 VP.n30 VSUBS 0.055744f
C853 VP.n31 VSUBS 0.063285f
C854 VP.n32 VSUBS 0.913103f
C855 VP.n33 VSUBS 0.04266f
C856 VDD2.n0 VSUBS 0.025815f
C857 VDD2.n1 VSUBS 0.024936f
C858 VDD2.n2 VSUBS 0.0134f
C859 VDD2.n3 VSUBS 0.031672f
C860 VDD2.n4 VSUBS 0.014188f
C861 VDD2.n5 VSUBS 0.024936f
C862 VDD2.n6 VSUBS 0.0134f
C863 VDD2.n7 VSUBS 0.031672f
C864 VDD2.n8 VSUBS 0.014188f
C865 VDD2.n9 VSUBS 0.024936f
C866 VDD2.n10 VSUBS 0.0134f
C867 VDD2.n11 VSUBS 0.031672f
C868 VDD2.n12 VSUBS 0.014188f
C869 VDD2.n13 VSUBS 0.024936f
C870 VDD2.n14 VSUBS 0.0134f
C871 VDD2.n15 VSUBS 0.031672f
C872 VDD2.n16 VSUBS 0.014188f
C873 VDD2.n17 VSUBS 0.180832f
C874 VDD2.t4 VSUBS 0.068139f
C875 VDD2.n18 VSUBS 0.023754f
C876 VDD2.n19 VSUBS 0.023825f
C877 VDD2.n20 VSUBS 0.0134f
C878 VDD2.n21 VSUBS 1.0744f
C879 VDD2.n22 VSUBS 0.024936f
C880 VDD2.n23 VSUBS 0.0134f
C881 VDD2.n24 VSUBS 0.014188f
C882 VDD2.n25 VSUBS 0.031672f
C883 VDD2.n26 VSUBS 0.031672f
C884 VDD2.n27 VSUBS 0.014188f
C885 VDD2.n28 VSUBS 0.0134f
C886 VDD2.n29 VSUBS 0.024936f
C887 VDD2.n30 VSUBS 0.024936f
C888 VDD2.n31 VSUBS 0.0134f
C889 VDD2.n32 VSUBS 0.014188f
C890 VDD2.n33 VSUBS 0.031672f
C891 VDD2.n34 VSUBS 0.031672f
C892 VDD2.n35 VSUBS 0.031672f
C893 VDD2.n36 VSUBS 0.014188f
C894 VDD2.n37 VSUBS 0.0134f
C895 VDD2.n38 VSUBS 0.024936f
C896 VDD2.n39 VSUBS 0.024936f
C897 VDD2.n40 VSUBS 0.0134f
C898 VDD2.n41 VSUBS 0.013794f
C899 VDD2.n42 VSUBS 0.013794f
C900 VDD2.n43 VSUBS 0.031672f
C901 VDD2.n44 VSUBS 0.031672f
C902 VDD2.n45 VSUBS 0.014188f
C903 VDD2.n46 VSUBS 0.0134f
C904 VDD2.n47 VSUBS 0.024936f
C905 VDD2.n48 VSUBS 0.024936f
C906 VDD2.n49 VSUBS 0.0134f
C907 VDD2.n50 VSUBS 0.014188f
C908 VDD2.n51 VSUBS 0.031672f
C909 VDD2.n52 VSUBS 0.071278f
C910 VDD2.n53 VSUBS 0.014188f
C911 VDD2.n54 VSUBS 0.0134f
C912 VDD2.n55 VSUBS 0.055595f
C913 VDD2.n56 VSUBS 0.058019f
C914 VDD2.t1 VSUBS 0.209269f
C915 VDD2.t5 VSUBS 0.209269f
C916 VDD2.n57 VSUBS 1.59825f
C917 VDD2.n58 VSUBS 2.62849f
C918 VDD2.n59 VSUBS 0.025815f
C919 VDD2.n60 VSUBS 0.024936f
C920 VDD2.n61 VSUBS 0.0134f
C921 VDD2.n62 VSUBS 0.031672f
C922 VDD2.n63 VSUBS 0.014188f
C923 VDD2.n64 VSUBS 0.024936f
C924 VDD2.n65 VSUBS 0.0134f
C925 VDD2.n66 VSUBS 0.031672f
C926 VDD2.n67 VSUBS 0.014188f
C927 VDD2.n68 VSUBS 0.024936f
C928 VDD2.n69 VSUBS 0.0134f
C929 VDD2.n70 VSUBS 0.031672f
C930 VDD2.n71 VSUBS 0.031672f
C931 VDD2.n72 VSUBS 0.014188f
C932 VDD2.n73 VSUBS 0.024936f
C933 VDD2.n74 VSUBS 0.0134f
C934 VDD2.n75 VSUBS 0.031672f
C935 VDD2.n76 VSUBS 0.014188f
C936 VDD2.n77 VSUBS 0.180832f
C937 VDD2.t3 VSUBS 0.068139f
C938 VDD2.n78 VSUBS 0.023754f
C939 VDD2.n79 VSUBS 0.023825f
C940 VDD2.n80 VSUBS 0.0134f
C941 VDD2.n81 VSUBS 1.0744f
C942 VDD2.n82 VSUBS 0.024936f
C943 VDD2.n83 VSUBS 0.0134f
C944 VDD2.n84 VSUBS 0.014188f
C945 VDD2.n85 VSUBS 0.031672f
C946 VDD2.n86 VSUBS 0.031672f
C947 VDD2.n87 VSUBS 0.014188f
C948 VDD2.n88 VSUBS 0.0134f
C949 VDD2.n89 VSUBS 0.024936f
C950 VDD2.n90 VSUBS 0.024936f
C951 VDD2.n91 VSUBS 0.0134f
C952 VDD2.n92 VSUBS 0.014188f
C953 VDD2.n93 VSUBS 0.031672f
C954 VDD2.n94 VSUBS 0.031672f
C955 VDD2.n95 VSUBS 0.014188f
C956 VDD2.n96 VSUBS 0.0134f
C957 VDD2.n97 VSUBS 0.024936f
C958 VDD2.n98 VSUBS 0.024936f
C959 VDD2.n99 VSUBS 0.0134f
C960 VDD2.n100 VSUBS 0.013794f
C961 VDD2.n101 VSUBS 0.013794f
C962 VDD2.n102 VSUBS 0.031672f
C963 VDD2.n103 VSUBS 0.031672f
C964 VDD2.n104 VSUBS 0.014188f
C965 VDD2.n105 VSUBS 0.0134f
C966 VDD2.n106 VSUBS 0.024936f
C967 VDD2.n107 VSUBS 0.024936f
C968 VDD2.n108 VSUBS 0.0134f
C969 VDD2.n109 VSUBS 0.014188f
C970 VDD2.n110 VSUBS 0.031672f
C971 VDD2.n111 VSUBS 0.071278f
C972 VDD2.n112 VSUBS 0.014188f
C973 VDD2.n113 VSUBS 0.0134f
C974 VDD2.n114 VSUBS 0.055595f
C975 VDD2.n115 VSUBS 0.052776f
C976 VDD2.n116 VSUBS 2.31339f
C977 VDD2.t0 VSUBS 0.209269f
C978 VDD2.t2 VSUBS 0.209269f
C979 VDD2.n117 VSUBS 1.59822f
C980 VTAIL.t6 VSUBS 0.245514f
C981 VTAIL.t10 VSUBS 0.245514f
C982 VTAIL.n0 VSUBS 1.71632f
C983 VTAIL.n1 VSUBS 0.852946f
C984 VTAIL.n2 VSUBS 0.030286f
C985 VTAIL.n3 VSUBS 0.029255f
C986 VTAIL.n4 VSUBS 0.01572f
C987 VTAIL.n5 VSUBS 0.037157f
C988 VTAIL.n6 VSUBS 0.016645f
C989 VTAIL.n7 VSUBS 0.029255f
C990 VTAIL.n8 VSUBS 0.01572f
C991 VTAIL.n9 VSUBS 0.037157f
C992 VTAIL.n10 VSUBS 0.016645f
C993 VTAIL.n11 VSUBS 0.029255f
C994 VTAIL.n12 VSUBS 0.01572f
C995 VTAIL.n13 VSUBS 0.037157f
C996 VTAIL.n14 VSUBS 0.016645f
C997 VTAIL.n15 VSUBS 0.029255f
C998 VTAIL.n16 VSUBS 0.01572f
C999 VTAIL.n17 VSUBS 0.037157f
C1000 VTAIL.n18 VSUBS 0.016645f
C1001 VTAIL.n19 VSUBS 0.212151f
C1002 VTAIL.t3 VSUBS 0.07994f
C1003 VTAIL.n20 VSUBS 0.027868f
C1004 VTAIL.n21 VSUBS 0.027951f
C1005 VTAIL.n22 VSUBS 0.01572f
C1006 VTAIL.n23 VSUBS 1.26048f
C1007 VTAIL.n24 VSUBS 0.029255f
C1008 VTAIL.n25 VSUBS 0.01572f
C1009 VTAIL.n26 VSUBS 0.016645f
C1010 VTAIL.n27 VSUBS 0.037157f
C1011 VTAIL.n28 VSUBS 0.037157f
C1012 VTAIL.n29 VSUBS 0.016645f
C1013 VTAIL.n30 VSUBS 0.01572f
C1014 VTAIL.n31 VSUBS 0.029255f
C1015 VTAIL.n32 VSUBS 0.029255f
C1016 VTAIL.n33 VSUBS 0.01572f
C1017 VTAIL.n34 VSUBS 0.016645f
C1018 VTAIL.n35 VSUBS 0.037157f
C1019 VTAIL.n36 VSUBS 0.037157f
C1020 VTAIL.n37 VSUBS 0.037157f
C1021 VTAIL.n38 VSUBS 0.016645f
C1022 VTAIL.n39 VSUBS 0.01572f
C1023 VTAIL.n40 VSUBS 0.029255f
C1024 VTAIL.n41 VSUBS 0.029255f
C1025 VTAIL.n42 VSUBS 0.01572f
C1026 VTAIL.n43 VSUBS 0.016183f
C1027 VTAIL.n44 VSUBS 0.016183f
C1028 VTAIL.n45 VSUBS 0.037157f
C1029 VTAIL.n46 VSUBS 0.037157f
C1030 VTAIL.n47 VSUBS 0.016645f
C1031 VTAIL.n48 VSUBS 0.01572f
C1032 VTAIL.n49 VSUBS 0.029255f
C1033 VTAIL.n50 VSUBS 0.029255f
C1034 VTAIL.n51 VSUBS 0.01572f
C1035 VTAIL.n52 VSUBS 0.016645f
C1036 VTAIL.n53 VSUBS 0.037157f
C1037 VTAIL.n54 VSUBS 0.083623f
C1038 VTAIL.n55 VSUBS 0.016645f
C1039 VTAIL.n56 VSUBS 0.01572f
C1040 VTAIL.n57 VSUBS 0.065223f
C1041 VTAIL.n58 VSUBS 0.041697f
C1042 VTAIL.n59 VSUBS 0.365347f
C1043 VTAIL.t5 VSUBS 0.245514f
C1044 VTAIL.t2 VSUBS 0.245514f
C1045 VTAIL.n60 VSUBS 1.71632f
C1046 VTAIL.n61 VSUBS 2.50972f
C1047 VTAIL.t11 VSUBS 0.245514f
C1048 VTAIL.t9 VSUBS 0.245514f
C1049 VTAIL.n62 VSUBS 1.71633f
C1050 VTAIL.n63 VSUBS 2.50971f
C1051 VTAIL.n64 VSUBS 0.030286f
C1052 VTAIL.n65 VSUBS 0.029255f
C1053 VTAIL.n66 VSUBS 0.01572f
C1054 VTAIL.n67 VSUBS 0.037157f
C1055 VTAIL.n68 VSUBS 0.016645f
C1056 VTAIL.n69 VSUBS 0.029255f
C1057 VTAIL.n70 VSUBS 0.01572f
C1058 VTAIL.n71 VSUBS 0.037157f
C1059 VTAIL.n72 VSUBS 0.016645f
C1060 VTAIL.n73 VSUBS 0.029255f
C1061 VTAIL.n74 VSUBS 0.01572f
C1062 VTAIL.n75 VSUBS 0.037157f
C1063 VTAIL.n76 VSUBS 0.037157f
C1064 VTAIL.n77 VSUBS 0.016645f
C1065 VTAIL.n78 VSUBS 0.029255f
C1066 VTAIL.n79 VSUBS 0.01572f
C1067 VTAIL.n80 VSUBS 0.037157f
C1068 VTAIL.n81 VSUBS 0.016645f
C1069 VTAIL.n82 VSUBS 0.212151f
C1070 VTAIL.t8 VSUBS 0.07994f
C1071 VTAIL.n83 VSUBS 0.027868f
C1072 VTAIL.n84 VSUBS 0.027951f
C1073 VTAIL.n85 VSUBS 0.01572f
C1074 VTAIL.n86 VSUBS 1.26048f
C1075 VTAIL.n87 VSUBS 0.029255f
C1076 VTAIL.n88 VSUBS 0.01572f
C1077 VTAIL.n89 VSUBS 0.016645f
C1078 VTAIL.n90 VSUBS 0.037157f
C1079 VTAIL.n91 VSUBS 0.037157f
C1080 VTAIL.n92 VSUBS 0.016645f
C1081 VTAIL.n93 VSUBS 0.01572f
C1082 VTAIL.n94 VSUBS 0.029255f
C1083 VTAIL.n95 VSUBS 0.029255f
C1084 VTAIL.n96 VSUBS 0.01572f
C1085 VTAIL.n97 VSUBS 0.016645f
C1086 VTAIL.n98 VSUBS 0.037157f
C1087 VTAIL.n99 VSUBS 0.037157f
C1088 VTAIL.n100 VSUBS 0.016645f
C1089 VTAIL.n101 VSUBS 0.01572f
C1090 VTAIL.n102 VSUBS 0.029255f
C1091 VTAIL.n103 VSUBS 0.029255f
C1092 VTAIL.n104 VSUBS 0.01572f
C1093 VTAIL.n105 VSUBS 0.016183f
C1094 VTAIL.n106 VSUBS 0.016183f
C1095 VTAIL.n107 VSUBS 0.037157f
C1096 VTAIL.n108 VSUBS 0.037157f
C1097 VTAIL.n109 VSUBS 0.016645f
C1098 VTAIL.n110 VSUBS 0.01572f
C1099 VTAIL.n111 VSUBS 0.029255f
C1100 VTAIL.n112 VSUBS 0.029255f
C1101 VTAIL.n113 VSUBS 0.01572f
C1102 VTAIL.n114 VSUBS 0.016645f
C1103 VTAIL.n115 VSUBS 0.037157f
C1104 VTAIL.n116 VSUBS 0.083623f
C1105 VTAIL.n117 VSUBS 0.016645f
C1106 VTAIL.n118 VSUBS 0.01572f
C1107 VTAIL.n119 VSUBS 0.065223f
C1108 VTAIL.n120 VSUBS 0.041697f
C1109 VTAIL.n121 VSUBS 0.365347f
C1110 VTAIL.t4 VSUBS 0.245514f
C1111 VTAIL.t0 VSUBS 0.245514f
C1112 VTAIL.n122 VSUBS 1.71633f
C1113 VTAIL.n123 VSUBS 0.99616f
C1114 VTAIL.n124 VSUBS 0.030286f
C1115 VTAIL.n125 VSUBS 0.029255f
C1116 VTAIL.n126 VSUBS 0.01572f
C1117 VTAIL.n127 VSUBS 0.037157f
C1118 VTAIL.n128 VSUBS 0.016645f
C1119 VTAIL.n129 VSUBS 0.029255f
C1120 VTAIL.n130 VSUBS 0.01572f
C1121 VTAIL.n131 VSUBS 0.037157f
C1122 VTAIL.n132 VSUBS 0.016645f
C1123 VTAIL.n133 VSUBS 0.029255f
C1124 VTAIL.n134 VSUBS 0.01572f
C1125 VTAIL.n135 VSUBS 0.037157f
C1126 VTAIL.n136 VSUBS 0.037157f
C1127 VTAIL.n137 VSUBS 0.016645f
C1128 VTAIL.n138 VSUBS 0.029255f
C1129 VTAIL.n139 VSUBS 0.01572f
C1130 VTAIL.n140 VSUBS 0.037157f
C1131 VTAIL.n141 VSUBS 0.016645f
C1132 VTAIL.n142 VSUBS 0.212151f
C1133 VTAIL.t1 VSUBS 0.07994f
C1134 VTAIL.n143 VSUBS 0.027868f
C1135 VTAIL.n144 VSUBS 0.027951f
C1136 VTAIL.n145 VSUBS 0.01572f
C1137 VTAIL.n146 VSUBS 1.26048f
C1138 VTAIL.n147 VSUBS 0.029255f
C1139 VTAIL.n148 VSUBS 0.01572f
C1140 VTAIL.n149 VSUBS 0.016645f
C1141 VTAIL.n150 VSUBS 0.037157f
C1142 VTAIL.n151 VSUBS 0.037157f
C1143 VTAIL.n152 VSUBS 0.016645f
C1144 VTAIL.n153 VSUBS 0.01572f
C1145 VTAIL.n154 VSUBS 0.029255f
C1146 VTAIL.n155 VSUBS 0.029255f
C1147 VTAIL.n156 VSUBS 0.01572f
C1148 VTAIL.n157 VSUBS 0.016645f
C1149 VTAIL.n158 VSUBS 0.037157f
C1150 VTAIL.n159 VSUBS 0.037157f
C1151 VTAIL.n160 VSUBS 0.016645f
C1152 VTAIL.n161 VSUBS 0.01572f
C1153 VTAIL.n162 VSUBS 0.029255f
C1154 VTAIL.n163 VSUBS 0.029255f
C1155 VTAIL.n164 VSUBS 0.01572f
C1156 VTAIL.n165 VSUBS 0.016183f
C1157 VTAIL.n166 VSUBS 0.016183f
C1158 VTAIL.n167 VSUBS 0.037157f
C1159 VTAIL.n168 VSUBS 0.037157f
C1160 VTAIL.n169 VSUBS 0.016645f
C1161 VTAIL.n170 VSUBS 0.01572f
C1162 VTAIL.n171 VSUBS 0.029255f
C1163 VTAIL.n172 VSUBS 0.029255f
C1164 VTAIL.n173 VSUBS 0.01572f
C1165 VTAIL.n174 VSUBS 0.016645f
C1166 VTAIL.n175 VSUBS 0.037157f
C1167 VTAIL.n176 VSUBS 0.083623f
C1168 VTAIL.n177 VSUBS 0.016645f
C1169 VTAIL.n178 VSUBS 0.01572f
C1170 VTAIL.n179 VSUBS 0.065223f
C1171 VTAIL.n180 VSUBS 0.041697f
C1172 VTAIL.n181 VSUBS 1.68061f
C1173 VTAIL.n182 VSUBS 0.030286f
C1174 VTAIL.n183 VSUBS 0.029255f
C1175 VTAIL.n184 VSUBS 0.01572f
C1176 VTAIL.n185 VSUBS 0.037157f
C1177 VTAIL.n186 VSUBS 0.016645f
C1178 VTAIL.n187 VSUBS 0.029255f
C1179 VTAIL.n188 VSUBS 0.01572f
C1180 VTAIL.n189 VSUBS 0.037157f
C1181 VTAIL.n190 VSUBS 0.016645f
C1182 VTAIL.n191 VSUBS 0.029255f
C1183 VTAIL.n192 VSUBS 0.01572f
C1184 VTAIL.n193 VSUBS 0.037157f
C1185 VTAIL.n194 VSUBS 0.016645f
C1186 VTAIL.n195 VSUBS 0.029255f
C1187 VTAIL.n196 VSUBS 0.01572f
C1188 VTAIL.n197 VSUBS 0.037157f
C1189 VTAIL.n198 VSUBS 0.016645f
C1190 VTAIL.n199 VSUBS 0.212151f
C1191 VTAIL.t7 VSUBS 0.07994f
C1192 VTAIL.n200 VSUBS 0.027868f
C1193 VTAIL.n201 VSUBS 0.027951f
C1194 VTAIL.n202 VSUBS 0.01572f
C1195 VTAIL.n203 VSUBS 1.26048f
C1196 VTAIL.n204 VSUBS 0.029255f
C1197 VTAIL.n205 VSUBS 0.01572f
C1198 VTAIL.n206 VSUBS 0.016645f
C1199 VTAIL.n207 VSUBS 0.037157f
C1200 VTAIL.n208 VSUBS 0.037157f
C1201 VTAIL.n209 VSUBS 0.016645f
C1202 VTAIL.n210 VSUBS 0.01572f
C1203 VTAIL.n211 VSUBS 0.029255f
C1204 VTAIL.n212 VSUBS 0.029255f
C1205 VTAIL.n213 VSUBS 0.01572f
C1206 VTAIL.n214 VSUBS 0.016645f
C1207 VTAIL.n215 VSUBS 0.037157f
C1208 VTAIL.n216 VSUBS 0.037157f
C1209 VTAIL.n217 VSUBS 0.037157f
C1210 VTAIL.n218 VSUBS 0.016645f
C1211 VTAIL.n219 VSUBS 0.01572f
C1212 VTAIL.n220 VSUBS 0.029255f
C1213 VTAIL.n221 VSUBS 0.029255f
C1214 VTAIL.n222 VSUBS 0.01572f
C1215 VTAIL.n223 VSUBS 0.016183f
C1216 VTAIL.n224 VSUBS 0.016183f
C1217 VTAIL.n225 VSUBS 0.037157f
C1218 VTAIL.n226 VSUBS 0.037157f
C1219 VTAIL.n227 VSUBS 0.016645f
C1220 VTAIL.n228 VSUBS 0.01572f
C1221 VTAIL.n229 VSUBS 0.029255f
C1222 VTAIL.n230 VSUBS 0.029255f
C1223 VTAIL.n231 VSUBS 0.01572f
C1224 VTAIL.n232 VSUBS 0.016645f
C1225 VTAIL.n233 VSUBS 0.037157f
C1226 VTAIL.n234 VSUBS 0.083623f
C1227 VTAIL.n235 VSUBS 0.016645f
C1228 VTAIL.n236 VSUBS 0.01572f
C1229 VTAIL.n237 VSUBS 0.065223f
C1230 VTAIL.n238 VSUBS 0.041697f
C1231 VTAIL.n239 VSUBS 1.62555f
C1232 VN.n0 VSUBS 0.046124f
C1233 VN.t0 VSUBS 2.12817f
C1234 VN.n1 VSUBS 0.047955f
C1235 VN.t1 VSUBS 2.33951f
C1236 VN.n2 VSUBS 0.837477f
C1237 VN.t4 VSUBS 2.12817f
C1238 VN.n3 VSUBS 0.869367f
C1239 VN.n4 VSUBS 0.06488f
C1240 VN.n5 VSUBS 0.294546f
C1241 VN.n6 VSUBS 0.034987f
C1242 VN.n7 VSUBS 0.034987f
C1243 VN.n8 VSUBS 0.053763f
C1244 VN.n9 VSUBS 0.061037f
C1245 VN.n10 VSUBS 0.88066f
C1246 VN.n11 VSUBS 0.041144f
C1247 VN.n12 VSUBS 0.046124f
C1248 VN.t2 VSUBS 2.12817f
C1249 VN.n13 VSUBS 0.047955f
C1250 VN.t3 VSUBS 2.33951f
C1251 VN.n14 VSUBS 0.837477f
C1252 VN.t5 VSUBS 2.12817f
C1253 VN.n15 VSUBS 0.869367f
C1254 VN.n16 VSUBS 0.06488f
C1255 VN.n17 VSUBS 0.294546f
C1256 VN.n18 VSUBS 0.034987f
C1257 VN.n19 VSUBS 0.034987f
C1258 VN.n20 VSUBS 0.053763f
C1259 VN.n21 VSUBS 0.061037f
C1260 VN.n22 VSUBS 0.88066f
C1261 VN.n23 VSUBS 1.70908f
.ends

