* NGSPICE file created from opamp_sample_0002.ext - technology: sky130A

.subckt opamp_sample_0002 GND VOUT VDD VN VP CS_BIAS DIFFPAIR_BIAS
X0 a_n11986_8880.t13 a_n5004_9136.t22 a_n3584_7550.t1 VDD.t112 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=1.6536 ps=9.26 w=4.24 l=2.43
X1 a_n1672_n179.t10 DIFFPAIR_BIAS.t6 GND.t171 GND.t170 sky130_fd_pr__nfet_01v8 ad=1.5678 pd=8.82 as=1.5678 ps=8.82 w=4.02 l=3.07
X2 GND.t153 GND.t151 GND.t152 GND.t34 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=4.65
X3 VOUT.t35 CS_BIAS.t12 GND.t22 GND.t20 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=1.3572 ps=7.74 w=3.48 l=4.65
X4 a_n3584_7550.t14 a_n5004_9136.t23 VDD.t114 VDD.t113 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=0.6996 ps=4.57 w=4.24 l=2.43
X5 VDD.t55 VDD.t53 VDD.t54 VDD.t50 sky130_fd_pr__pfet_01v8 ad=1.6536 pd=9.26 as=0 ps=0 w=4.24 l=2.43
X6 a_n5004_9136.t3 VP.t7 a_n1672_n179.t6 GND.t8 sky130_fd_pr__nfet_01v8 ad=1.6107 pd=9.04 as=0.68145 ps=4.46 w=4.13 l=2.2
X7 GND.t150 GND.t148 GND.t149 GND.t84 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=4.65
X8 GND.t147 GND.t145 VN.t6 GND.t146 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X9 a_n11986_8880.t2 VN.t7 a_n1672_n179.t5 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.68145 pd=4.46 as=1.6107 ps=9.04 w=4.13 l=2.2
X10 a_n3584_7550.t2 a_n5004_9136.t24 a_n11986_8880.t12 VDD.t93 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=0.6996 ps=4.57 w=4.24 l=2.43
X11 a_n5082_9332.t15 a_n5004_9136.t14 a_n5004_9136.t15 VDD.t77 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=1.6536 ps=9.26 w=4.24 l=2.43
X12 GND.t15 CS_BIAS.t13 VOUT.t34 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=0.5742 ps=3.81 w=3.48 l=4.65
X13 GND.t23 CS_BIAS.t14 VOUT.t33 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=0.5742 ps=3.81 w=3.48 l=4.65
X14 VDD.t52 VDD.t49 VDD.t51 VDD.t50 sky130_fd_pr__pfet_01v8 ad=1.6536 pd=9.26 as=0 ps=0 w=4.24 l=2.43
X15 VOUT.t11 a_n11986_8880.t14 VDD.t74 VDD.t62 sky130_fd_pr__pfet_01v8 ad=0.33165 pd=2.34 as=0.7839 ps=4.8 w=2.01 l=5.87
X16 CS_BIAS.t11 CS_BIAS.t10 GND.t159 GND.t20 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=1.3572 ps=7.74 w=3.48 l=4.65
X17 GND.t144 GND.t142 GND.t143 GND.t74 sky130_fd_pr__nfet_01v8 ad=1.6107 pd=9.04 as=0 ps=0 w=4.13 l=2.2
X18 GND.t126 GND.t124 VN.t5 GND.t125 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X19 a_n3584_7550.t11 a_n5004_9136.t25 a_n11986_8880.t11 VDD.t111 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=0.6996 ps=4.57 w=4.24 l=2.43
X20 a_n5082_9332.t14 a_n5004_9136.t8 a_n5004_9136.t9 VDD.t112 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=1.6536 ps=9.26 w=4.24 l=2.43
X21 GND.t141 GND.t139 GND.t140 GND.t61 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=4.65
X22 VP.t6 GND.t136 GND.t138 GND.t137 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X23 VOUT.t10 a_n11986_8880.t15 VDD.t73 VDD.t59 sky130_fd_pr__pfet_01v8 ad=0.33165 pd=2.34 as=0.7839 ps=4.8 w=2.01 l=5.87
X24 a_n5004_9136.t11 a_n5004_9136.t10 a_n5082_9332.t13 VDD.t111 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=0.6996 ps=4.57 w=4.24 l=2.43
X25 VDD.t48 VDD.t46 VDD.t47 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0.7839 pd=4.8 as=0 ps=0 w=2.01 l=5.87
X26 VOUT.t32 CS_BIAS.t15 GND.t12 GND.t11 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0.5742 ps=3.81 w=3.48 l=4.65
X27 VDD.t110 a_n5004_9136.t26 a_n3584_7550.t5 VDD.t109 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=1.6536 ps=9.26 w=4.24 l=2.43
X28 VOUT.t9 a_n11986_8880.t16 VDD.t72 VDD.t70 sky130_fd_pr__pfet_01v8 ad=0.7839 pd=4.8 as=0.33165 ps=2.34 w=2.01 l=5.87
X29 GND.t135 GND.t133 GND.t134 GND.t34 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=4.65
X30 VOUT.t8 a_n11986_8880.t17 VDD.t71 VDD.t70 sky130_fd_pr__pfet_01v8 ad=0.7839 pd=4.8 as=0.33165 ps=2.34 w=2.01 l=5.87
X31 DIFFPAIR_BIAS.t5 DIFFPAIR_BIAS.t4 GND.t169 GND.t168 sky130_fd_pr__nfet_01v8 ad=1.5678 pd=8.82 as=1.5678 ps=8.82 w=4.02 l=3.07
X32 VDD.t108 a_n5004_9136.t27 a_n3584_7550.t4 VDD.t107 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=1.6536 ps=9.26 w=4.24 l=2.43
X33 VOUT.t31 CS_BIAS.t16 GND.t180 GND.t11 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0.5742 ps=3.81 w=3.48 l=4.65
X34 GND.t132 GND.t130 VN.t4 GND.t131 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X35 VP.t5 GND.t127 GND.t129 GND.t128 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X36 VDD.t45 VDD.t43 VDD.t44 VDD.t40 sky130_fd_pr__pfet_01v8 ad=1.6536 pd=9.26 as=0 ps=0 w=4.24 l=2.43
X37 VDD.t42 VDD.t39 VDD.t41 VDD.t40 sky130_fd_pr__pfet_01v8 ad=1.6536 pd=9.26 as=0 ps=0 w=4.24 l=2.43
X38 GND.t123 GND.t121 GND.t122 GND.t44 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=4.65
X39 a_5210_9332# a_5210_9332# a_5210_9332# VDD.t115 sky130_fd_pr__pfet_01v8 ad=1.6536 pd=9.26 as=3.3072 ps=18.52 w=4.24 l=2.43
X40 a_n3584_7550.t8 a_n5004_9136.t28 a_n11986_8880.t10 VDD.t88 sky130_fd_pr__pfet_01v8 ad=1.6536 pd=9.26 as=0.6996 ps=4.57 w=4.24 l=2.43
X41 GND.t175 CS_BIAS.t17 VOUT.t30 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=0.5742 ps=3.81 w=3.48 l=4.65
X42 GND.t120 GND.t118 VN.t3 GND.t119 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X43 VDD.t38 VDD.t36 VDD.t37 VDD.t16 sky130_fd_pr__pfet_01v8 ad=1.6536 pd=9.26 as=0 ps=0 w=4.24 l=2.43
X44 GND.t117 GND.t115 GND.t116 GND.t44 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=4.65
X45 a_n5004_9136.t1 VP.t8 a_n1672_n179.t1 GND.t1 sky130_fd_pr__nfet_01v8 ad=1.6107 pd=9.04 as=0.68145 ps=4.46 w=4.13 l=2.2
X46 VOUT.t29 CS_BIAS.t18 GND.t158 GND.t20 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=1.3572 ps=7.74 w=3.48 l=4.65
X47 VDD.t35 VDD.t33 VDD.t34 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.7839 pd=4.8 as=0 ps=0 w=2.01 l=5.87
X48 VOUT.t28 CS_BIAS.t19 GND.t155 GND.t11 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0.5742 ps=3.81 w=3.48 l=4.65
X49 VOUT.t36 a_n3584_7550.t0 sky130_fd_pr__cap_mim_m3_1 l=10.17 w=15.34
X50 VOUT.t27 CS_BIAS.t20 GND.t7 GND.t3 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=1.3572 ps=7.74 w=3.48 l=4.65
X51 a_n1672_n179.t11 VN.t8 a_n11986_8880.t4 GND.t176 sky130_fd_pr__nfet_01v8 ad=0.68145 pd=4.46 as=0.68145 ps=4.46 w=4.13 l=2.2
X52 VP.t4 GND.t112 GND.t114 GND.t113 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X53 GND.t111 GND.t109 GND.t110 GND.t44 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=4.65
X54 a_n11986_8880.t9 a_n5004_9136.t29 a_n3584_7550.t15 VDD.t102 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=0.6996 ps=4.57 w=4.24 l=2.43
X55 a_n11986_8880.t1 VN.t9 a_n1672_n179.t4 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.68145 pd=4.46 as=1.6107 ps=9.04 w=4.13 l=2.2
X56 VDD.t69 a_n11986_8880.t18 VOUT.t7 VDD.t64 sky130_fd_pr__pfet_01v8 ad=0.33165 pd=2.34 as=0.33165 ps=2.34 w=2.01 l=5.87
X57 GND.t17 CS_BIAS.t21 VOUT.t26 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=0.5742 ps=3.81 w=3.48 l=4.65
X58 a_n1672_n179.t2 VP.t9 a_n5004_9136.t2 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.68145 pd=4.46 as=0.68145 ps=4.46 w=4.13 l=2.2
X59 VDD.t106 a_n5004_9136.t30 a_n5082_9332.t7 VDD.t105 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=1.6536 ps=9.26 w=4.24 l=2.43
X60 VDD.t104 a_n5004_9136.t31 a_n5082_9332.t6 VDD.t103 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=0.6996 ps=4.57 w=4.24 l=2.43
X61 GND.t108 GND.t105 GND.t107 GND.t106 sky130_fd_pr__nfet_01v8 ad=1.5678 pd=8.82 as=0 ps=0 w=4.02 l=3.07
X62 VDD.t32 VDD.t30 VDD.t31 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.7839 pd=4.8 as=0 ps=0 w=2.01 l=5.87
X63 VOUT.t37 a_n3584_7550.t0 sky130_fd_pr__cap_mim_m3_1 l=10.17 w=15.34
X64 a_n5082_9332.t12 a_n5004_9136.t6 a_n5004_9136.t7 VDD.t102 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=0.6996 ps=4.57 w=4.24 l=2.43
X65 a_n3584_7550.t10 a_n5004_9136.t32 a_n11986_8880.t8 VDD.t80 sky130_fd_pr__pfet_01v8 ad=1.6536 pd=9.26 as=0.6996 ps=4.57 w=4.24 l=2.43
X66 GND.t104 GND.t102 GND.t103 GND.t84 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=4.65
X67 a_n5082_9332.t5 a_n5004_9136.t33 VDD.t101 VDD.t100 sky130_fd_pr__pfet_01v8 ad=1.6536 pd=9.26 as=0.6996 ps=4.57 w=4.24 l=2.43
X68 VOUT.t25 CS_BIAS.t22 GND.t156 GND.t5 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0.5742 ps=3.81 w=3.48 l=4.65
X69 VOUT.t24 CS_BIAS.t23 GND.t21 GND.t20 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=1.3572 ps=7.74 w=3.48 l=4.65
X70 GND.t101 GND.t99 GND.t100 GND.t44 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=4.65
X71 VOUT.t23 CS_BIAS.t24 GND.t25 GND.t3 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=1.3572 ps=7.74 w=3.48 l=4.65
X72 a_n1672_n179.t9 DIFFPAIR_BIAS.t7 GND.t167 GND.t166 sky130_fd_pr__nfet_01v8 ad=1.5678 pd=8.82 as=1.5678 ps=8.82 w=4.02 l=3.07
X73 GND.t98 GND.t96 GND.t97 GND.t84 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=4.65
X74 GND.t95 GND.t93 GND.t94 GND.t61 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=4.65
X75 GND.t39 GND.t37 GND.t38 GND.t27 sky130_fd_pr__nfet_01v8 ad=1.6107 pd=9.04 as=0 ps=0 w=4.13 l=2.2
X76 GND.t18 CS_BIAS.t25 VOUT.t22 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=0.5742 ps=3.81 w=3.48 l=4.65
X77 a_n5082_9332.t4 a_n5004_9136.t34 VDD.t99 VDD.t98 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=0.6996 ps=4.57 w=4.24 l=2.43
X78 CS_BIAS.t9 CS_BIAS.t8 GND.t24 GND.t5 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0.5742 ps=3.81 w=3.48 l=4.65
X79 GND.t92 GND.t90 GND.t91 GND.t61 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=4.65
X80 VDD.t29 VDD.t27 VDD.t28 VDD.t24 sky130_fd_pr__pfet_01v8 ad=1.6536 pd=9.26 as=0 ps=0 w=4.24 l=2.43
X81 DIFFPAIR_BIAS.t3 DIFFPAIR_BIAS.t2 GND.t165 GND.t164 sky130_fd_pr__nfet_01v8 ad=1.5678 pd=8.82 as=1.5678 ps=8.82 w=4.02 l=3.07
X82 a_n11986_8880.t0 VN.t10 a_n1672_n179.t3 GND.t8 sky130_fd_pr__nfet_01v8 ad=1.6107 pd=9.04 as=0.68145 ps=4.46 w=4.13 l=2.2
X83 a_n3584_7550.t9 a_n5004_9136.t35 VDD.t97 VDD.t96 sky130_fd_pr__pfet_01v8 ad=1.6536 pd=9.26 as=0.6996 ps=4.57 w=4.24 l=2.43
X84 a_n5004_9136.t0 VP.t10 a_n1672_n179.t0 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.68145 pd=4.46 as=1.6107 ps=9.04 w=4.13 l=2.2
X85 VOUT.t21 CS_BIAS.t26 GND.t177 GND.t20 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=1.3572 ps=7.74 w=3.48 l=4.65
X86 GND.t89 GND.t87 GND.t88 GND.t84 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=4.65
X87 a_n5852_9332# a_n5852_9332# a_n5852_9332# VDD.t56 sky130_fd_pr__pfet_01v8 ad=1.6536 pd=9.26 as=3.3072 ps=18.52 w=4.24 l=2.43
X88 GND.t86 GND.t83 GND.t85 GND.t84 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=4.65
X89 a_n5082_9332.t3 a_n5004_9136.t36 VDD.t95 VDD.t94 sky130_fd_pr__pfet_01v8 ad=1.6536 pd=9.26 as=0.6996 ps=4.57 w=4.24 l=2.43
X90 GND.t19 CS_BIAS.t27 VOUT.t20 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=0.5742 ps=3.81 w=3.48 l=4.65
X91 GND.t66 GND.t64 GND.t65 GND.t34 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=4.65
X92 GND.t82 GND.t80 VP.t3 GND.t81 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X93 GND.t79 GND.t77 GND.t78 GND.t61 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=4.65
X94 GND.t76 GND.t73 GND.t75 GND.t74 sky130_fd_pr__nfet_01v8 ad=1.6107 pd=9.04 as=0 ps=0 w=4.13 l=2.2
X95 VDD.t26 VDD.t23 VDD.t25 VDD.t24 sky130_fd_pr__pfet_01v8 ad=1.6536 pd=9.26 as=0 ps=0 w=4.24 l=2.43
X96 GND.t63 GND.t60 GND.t62 GND.t61 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=4.65
X97 a_n5004_9136.t13 a_n5004_9136.t12 a_n5082_9332.t11 VDD.t93 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=0.6996 ps=4.57 w=4.24 l=2.43
X98 VDD.t22 VDD.t19 VDD.t21 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.7839 pd=4.8 as=0 ps=0 w=2.01 l=5.87
X99 GND.t72 GND.t70 GND.t71 GND.t34 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=4.65
X100 VOUT.t6 a_n11986_8880.t19 VDD.t68 VDD.t66 sky130_fd_pr__pfet_01v8 ad=0.7839 pd=4.8 as=0.33165 ps=2.34 w=2.01 l=5.87
X101 VDD.t92 a_n5004_9136.t37 a_n3584_7550.t12 VDD.t91 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=0.6996 ps=4.57 w=4.24 l=2.43
X102 a_n3584_7550.t13 a_n5004_9136.t38 VDD.t90 VDD.t89 sky130_fd_pr__pfet_01v8 ad=1.6536 pd=9.26 as=0.6996 ps=4.57 w=4.24 l=2.43
X103 VOUT.t19 CS_BIAS.t28 GND.t179 GND.t5 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0.5742 ps=3.81 w=3.48 l=4.65
X104 VN.t2 GND.t67 GND.t69 GND.t68 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X105 VDD.t18 VDD.t15 VDD.t17 VDD.t16 sky130_fd_pr__pfet_01v8 ad=1.6536 pd=9.26 as=0 ps=0 w=4.24 l=2.43
X106 a_n11986_8880.t7 a_n5004_9136.t39 a_n3584_7550.t16 VDD.t85 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=0.6996 ps=4.57 w=4.24 l=2.43
X107 GND.t59 GND.t57 VP.t2 GND.t58 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X108 a_n5004_9136.t17 a_n5004_9136.t16 a_n5082_9332.t10 VDD.t88 sky130_fd_pr__pfet_01v8 ad=1.6536 pd=9.26 as=0.6996 ps=4.57 w=4.24 l=2.43
X109 CS_BIAS.t7 CS_BIAS.t6 GND.t10 GND.t3 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=1.3572 ps=7.74 w=3.48 l=4.65
X110 a_n1672_n179.t8 DIFFPAIR_BIAS.t8 GND.t163 GND.t162 sky130_fd_pr__nfet_01v8 ad=1.5678 pd=8.82 as=1.5678 ps=8.82 w=4.02 l=3.07
X111 GND.t56 GND.t53 GND.t55 GND.t54 sky130_fd_pr__nfet_01v8 ad=1.5678 pd=8.82 as=0 ps=0 w=4.02 l=3.07
X112 VN.t1 GND.t50 GND.t52 GND.t51 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X113 VOUT.t5 a_n11986_8880.t20 VDD.t67 VDD.t66 sky130_fd_pr__pfet_01v8 ad=0.7839 pd=4.8 as=0.33165 ps=2.34 w=2.01 l=5.87
X114 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.t0 GND.t161 GND.t160 sky130_fd_pr__nfet_01v8 ad=1.5678 pd=8.82 as=1.5678 ps=8.82 w=4.02 l=3.07
X115 GND.t49 GND.t47 VP.t1 GND.t48 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X116 a_n5082_9332.t2 a_n5004_9136.t40 VDD.t87 VDD.t86 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=0.6996 ps=4.57 w=4.24 l=2.43
X117 VOUT.t18 CS_BIAS.t29 GND.t13 GND.t11 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0.5742 ps=3.81 w=3.48 l=4.65
X118 a_n5082_9332.t9 a_n5004_9136.t18 a_n5004_9136.t19 VDD.t85 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=0.6996 ps=4.57 w=4.24 l=2.43
X119 a_n1672_n179.t13 VP.t11 a_n5004_9136.t5 GND.t176 sky130_fd_pr__nfet_01v8 ad=0.68145 pd=4.46 as=0.68145 ps=4.46 w=4.13 l=2.2
X120 VDD.t14 VDD.t12 VDD.t13 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.7839 pd=4.8 as=0 ps=0 w=2.01 l=5.87
X121 VDD.t65 a_n11986_8880.t21 VOUT.t4 VDD.t64 sky130_fd_pr__pfet_01v8 ad=0.33165 pd=2.34 as=0.33165 ps=2.34 w=2.01 l=5.87
X122 VDD.t11 VDD.t8 VDD.t10 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0.7839 pd=4.8 as=0 ps=0 w=2.01 l=5.87
X123 GND.t157 CS_BIAS.t4 CS_BIAS.t5 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=0.5742 ps=3.81 w=3.48 l=4.65
X124 a_n11986_8880.t5 VN.t11 a_n1672_n179.t14 GND.t1 sky130_fd_pr__nfet_01v8 ad=1.6107 pd=9.04 as=0.68145 ps=4.46 w=4.13 l=2.2
X125 VDD.t84 a_n5004_9136.t41 a_n3584_7550.t7 VDD.t83 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=0.6996 ps=4.57 w=4.24 l=2.43
X126 GND.t46 GND.t43 GND.t45 GND.t44 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=4.65
X127 VOUT.t3 a_n11986_8880.t22 VDD.t63 VDD.t62 sky130_fd_pr__pfet_01v8 ad=0.33165 pd=2.34 as=0.7839 ps=4.8 w=2.01 l=5.87
X128 VOUT.t17 CS_BIAS.t30 GND.t173 GND.t5 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0.5742 ps=3.81 w=3.48 l=4.65
X129 GND.t36 GND.t33 GND.t35 GND.t34 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0 ps=0 w=3.48 l=4.65
X130 GND.t172 CS_BIAS.t31 VOUT.t16 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=0.5742 ps=3.81 w=3.48 l=4.65
X131 a_n1672_n179.t7 VN.t12 a_n11986_8880.t3 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.68145 pd=4.46 as=0.68145 ps=4.46 w=4.13 l=2.2
X132 VDD.t7 VDD.t4 VDD.t6 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.7839 pd=4.8 as=0 ps=0 w=2.01 l=5.87
X133 VDD.t61 a_n11986_8880.t23 VOUT.t2 VDD.t57 sky130_fd_pr__pfet_01v8 ad=0.33165 pd=2.34 as=0.33165 ps=2.34 w=2.01 l=5.87
X134 VOUT.t15 CS_BIAS.t32 GND.t4 GND.t3 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=1.3572 ps=7.74 w=3.48 l=4.65
X135 a_n5004_9136.t4 VP.t12 a_n1672_n179.t12 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.68145 pd=4.46 as=1.6107 ps=9.04 w=4.13 l=2.2
X136 VN.t0 GND.t40 GND.t42 GND.t41 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X137 GND.t32 GND.t30 VP.t0 GND.t31 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X138 VDD.t82 a_n5004_9136.t42 a_n5082_9332.t1 VDD.t81 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=1.6536 ps=9.26 w=4.24 l=2.43
X139 VOUT.t38 a_n3584_7550.t0 sky130_fd_pr__cap_mim_m3_1 l=10.17 w=15.34
X140 a_n5004_9136.t21 a_n5004_9136.t20 a_n5082_9332.t8 VDD.t80 sky130_fd_pr__pfet_01v8 ad=1.6536 pd=9.26 as=0.6996 ps=4.57 w=4.24 l=2.43
X141 VOUT.t14 CS_BIAS.t33 GND.t178 GND.t3 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=1.3572 ps=7.74 w=3.48 l=4.65
X142 a_n3584_7550.t6 a_n5004_9136.t43 VDD.t79 VDD.t78 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=0.6996 ps=4.57 w=4.24 l=2.43
X143 GND.t181 CS_BIAS.t2 CS_BIAS.t3 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=0.5742 ps=3.81 w=3.48 l=4.65
X144 VOUT.t13 CS_BIAS.t34 GND.t6 GND.t5 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0.5742 ps=3.81 w=3.48 l=4.65
X145 GND.t29 GND.t26 GND.t28 GND.t27 sky130_fd_pr__nfet_01v8 ad=1.6107 pd=9.04 as=0 ps=0 w=4.13 l=2.2
X146 GND.t174 CS_BIAS.t35 VOUT.t12 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.5742 pd=3.81 as=0.5742 ps=3.81 w=3.48 l=4.65
X147 VOUT.t1 a_n11986_8880.t24 VDD.t60 VDD.t59 sky130_fd_pr__pfet_01v8 ad=0.33165 pd=2.34 as=0.7839 ps=4.8 w=2.01 l=5.87
X148 CS_BIAS.t1 CS_BIAS.t0 GND.t154 GND.t11 sky130_fd_pr__nfet_01v8 ad=1.3572 pd=7.74 as=0.5742 ps=3.81 w=3.48 l=4.65
X149 VOUT.t39 a_n3584_7550.t0 sky130_fd_pr__cap_mim_m3_1 l=10.17 w=15.34
X150 a_n11986_8880.t6 a_n5004_9136.t44 a_n3584_7550.t3 VDD.t77 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=1.6536 ps=9.26 w=4.24 l=2.43
X151 VDD.t58 a_n11986_8880.t25 VOUT.t0 VDD.t57 sky130_fd_pr__pfet_01v8 ad=0.33165 pd=2.34 as=0.33165 ps=2.34 w=2.01 l=5.87
X152 VDD.t76 a_n5004_9136.t45 a_n5082_9332.t0 VDD.t75 sky130_fd_pr__pfet_01v8 ad=0.6996 pd=4.57 as=0.6996 ps=4.57 w=4.24 l=2.43
X153 VDD.t3 VDD.t0 VDD.t2 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.7839 pd=4.8 as=0 ps=0 w=2.01 l=5.87
R0 a_n5004_9136.n11 a_n5004_9136.n27 15.8745
R1 a_n5004_9136.n9 a_n5004_9136.n28 15.8745
R2 a_n5004_9136.n0 a_n5004_9136.n29 15.8745
R3 a_n5004_9136.n8 a_n5004_9136.n0 6.564
R4 a_n5004_9136.n4 a_n5004_9136.n3 6.56383
R5 a_n5004_9136.n3 a_n5004_9136.n30 15.8745
R6 a_n5004_9136.n21 a_n5004_9136.n3 6.56383
R7 a_n5004_9136.n3 a_n5004_9136.n31 15.8745
R8 a_n5004_9136.n36 a_n5004_9136.n5 74.9385
R9 a_n5004_9136.n5 a_n5004_9136.n32 15.8745
R10 a_n5004_9136.n6 a_n5004_9136.n33 15.8745
R11 a_n5004_9136.n7 a_n5004_9136.n6 6.564
R12 a_n5004_9136.n1 a_n5004_9136.n34 15.8745
R13 a_n5004_9136.n24 a_n5004_9136.t17 106.963
R14 a_n5004_9136.n25 a_n5004_9136.t9 106.963
R15 a_n5004_9136.n25 a_n5004_9136.t21 105.775
R16 a_n5004_9136.n24 a_n5004_9136.t15 105.773
R17 a_n5004_9136.n2 a_n5004_9136.n1 6.56383
R18 a_n5004_9136.n6 a_n5004_9136.n22 6.56383
R19 a_n5004_9136.n5 a_n5004_9136.n15 6.564
R20 a_n5004_9136.n6 a_n5004_9136.n35 15.4804
R21 a_n5004_9136.n3 a_n5004_9136.n16 6.564
R22 a_n5004_9136.n3 a_n5004_9136.n17 6.564
R23 a_n5004_9136.n9 a_n5004_9136.n10 6.564
R24 a_n5004_9136.n11 a_n5004_9136.n12 6.564
R25 a_n5004_9136.n11 a_n5004_9136.n18 6.56383
R26 a_n5004_9136.n0 a_n5004_9136.n20 6.56383
R27 a_n5004_9136.n24 a_n5004_9136.n38 98.1078
R28 a_n5004_9136.n25 a_n5004_9136.n49 98.1078
R29 a_n5004_9136.n56 a_n5004_9136.t3 93.0454
R30 a_n5004_9136.n26 a_n5004_9136.t1 92.2278
R31 a_n5004_9136.n57 a_n5004_9136.n26 87.7061
R32 a_n5004_9136.n56 a_n5004_9136.n55 87.706
R33 a_n5004_9136.n14 a_n5004_9136.t20 74.392
R34 a_n5004_9136.n47 a_n5004_9136.t18 42.0515
R35 a_n5004_9136.n48 a_n5004_9136.t12 42.0515
R36 a_n5004_9136.n2 a_n5004_9136.t8 74.3922
R37 a_n5004_9136.n7 a_n5004_9136.t36 74.392
R38 a_n5004_9136.n53 a_n5004_9136.t31 42.0515
R39 a_n5004_9136.n39 a_n5004_9136.t34 42.0515
R40 a_n5004_9136.n22 a_n5004_9136.t30 74.3922
R41 a_n5004_9136.n15 a_n5004_9136.t33 74.392
R42 a_n5004_9136.n52 a_n5004_9136.t45 42.0515
R43 a_n5004_9136.n40 a_n5004_9136.t40 42.0515
R44 a_n5004_9136.n35 a_n5004_9136.t42 66.8303
R45 a_n5004_9136.n16 a_n5004_9136.t35 74.392
R46 a_n5004_9136.n51 a_n5004_9136.t37 42.0515
R47 a_n5004_9136.n41 a_n5004_9136.t43 42.0515
R48 a_n5004_9136.n21 a_n5004_9136.t26 74.3922
R49 a_n5004_9136.n17 a_n5004_9136.t38 74.392
R50 a_n5004_9136.n50 a_n5004_9136.t41 42.0515
R51 a_n5004_9136.n42 a_n5004_9136.t23 42.0515
R52 a_n5004_9136.n4 a_n5004_9136.t27 74.3922
R53 a_n5004_9136.n10 a_n5004_9136.t16 74.392
R54 a_n5004_9136.n44 a_n5004_9136.t6 42.0515
R55 a_n5004_9136.n45 a_n5004_9136.t10 42.0515
R56 a_n5004_9136.n19 a_n5004_9136.t14 74.3922
R57 a_n5004_9136.n12 a_n5004_9136.t32 74.392
R58 a_n5004_9136.n43 a_n5004_9136.t39 42.0515
R59 a_n5004_9136.n46 a_n5004_9136.t24 42.0515
R60 a_n5004_9136.n18 a_n5004_9136.t22 74.3922
R61 a_n5004_9136.n8 a_n5004_9136.t28 74.392
R62 a_n5004_9136.n37 a_n5004_9136.t29 42.0515
R63 a_n5004_9136.n54 a_n5004_9136.t25 42.0515
R64 a_n5004_9136.n20 a_n5004_9136.t44 74.3922
R65 a_n5004_9136.n26 a_n5004_9136.n56 29.3882
R66 a_n5004_9136.n48 a_n5004_9136.n34 60.8154
R67 a_n5004_9136.n53 a_n5004_9136.n7 53.9331
R68 a_n5004_9136.n39 a_n5004_9136.n33 60.8154
R69 a_n5004_9136.n40 a_n5004_9136.n32 60.8154
R70 a_n5004_9136.n35 a_n5004_9136.n36 86.3406
R71 a_n5004_9136.n41 a_n5004_9136.n31 60.8154
R72 a_n5004_9136.n21 a_n5004_9136.n41 53.9331
R73 a_n5004_9136.n42 a_n5004_9136.n30 60.8154
R74 a_n5004_9136.n4 a_n5004_9136.n42 53.9331
R75 a_n5004_9136.n45 a_n5004_9136.n28 60.8154
R76 a_n5004_9136.n46 a_n5004_9136.n27 60.8154
R77 a_n5004_9136.n8 a_n5004_9136.n37 53.9331
R78 a_n5004_9136.n54 a_n5004_9136.n29 60.8154
R79 a_n5004_9136.n34 a_n5004_9136.n47 60.8156
R80 a_n5004_9136.n33 a_n5004_9136.n53 60.8156
R81 a_n5004_9136.n32 a_n5004_9136.n52 60.8156
R82 a_n5004_9136.n31 a_n5004_9136.n51 60.8156
R83 a_n5004_9136.n30 a_n5004_9136.n50 60.8156
R84 a_n5004_9136.n28 a_n5004_9136.n44 60.8156
R85 a_n5004_9136.n27 a_n5004_9136.n43 60.8156
R86 a_n5004_9136.n29 a_n5004_9136.n37 60.8156
R87 a_n5004_9136.n26 a_n5004_9136.n1 24.7357
R88 a_n5004_9136.n23 a_n5004_9136.n11 12.7766
R89 a_n5004_9136.n0 a_n5004_9136.n13 12.572
R90 a_n5004_9136.n23 a_n5004_9136.n1 11.2671
R91 a_n5004_9136.n9 a_n5004_9136.n13 9.23493
R92 a_n5004_9136.n38 a_n5004_9136.t7 7.66677
R93 a_n5004_9136.n38 a_n5004_9136.t11 7.66677
R94 a_n5004_9136.n49 a_n5004_9136.t19 7.66677
R95 a_n5004_9136.n49 a_n5004_9136.t13 7.66677
R96 a_n5004_9136.n14 a_n5004_9136.n47 53.9331
R97 a_n5004_9136.n48 a_n5004_9136.n2 53.9331
R98 a_n5004_9136.n22 a_n5004_9136.n39 53.9331
R99 a_n5004_9136.n52 a_n5004_9136.n15 53.9331
R100 a_n5004_9136.n36 a_n5004_9136.n40 17.328
R101 a_n5004_9136.n51 a_n5004_9136.n16 53.9331
R102 a_n5004_9136.n50 a_n5004_9136.n17 53.9331
R103 a_n5004_9136.n10 a_n5004_9136.n44 53.9331
R104 a_n5004_9136.n45 a_n5004_9136.n19 53.9331
R105 a_n5004_9136.n12 a_n5004_9136.n43 53.9331
R106 a_n5004_9136.n46 a_n5004_9136.n18 53.9331
R107 a_n5004_9136.n54 a_n5004_9136.n20 53.9331
R108 a_n5004_9136.n1 a_n5004_9136.n14 11.3067
R109 a_n5004_9136.n13 a_n5004_9136.n24 10.265
R110 a_n5004_9136.n5 a_n5004_9136.n3 10.1802
R111 a_n5004_9136.n9 a_n5004_9136.n19 10.1498
R112 a_n5004_9136.n13 a_n5004_9136.n6 9.93947
R113 a_n5004_9136.n11 a_n5004_9136.n9 9.22578
R114 a_n5004_9136.n6 a_n5004_9136.n5 8.30986
R115 a_n5004_9136.n23 a_n5004_9136.n25 8.22464
R116 a_n5004_9136.n1 a_n5004_9136.n0 8.03113
R117 a_n5004_9136.n3 a_n5004_9136.n23 7.70273
R118 a_n5004_9136.n55 a_n5004_9136.t2 4.79469
R119 a_n5004_9136.n55 a_n5004_9136.t4 4.79469
R120 a_n5004_9136.n57 a_n5004_9136.t5 4.79469
R121 a_n5004_9136.t0 a_n5004_9136.n57 4.79469
R122 a_n3584_7550.n0 a_n3584_7550.t5 106.963
R123 a_n3584_7550.n2 a_n3584_7550.t3 106.963
R124 a_n3584_7550.t1 a_n3584_7550.n3 106.963
R125 a_n3584_7550.n3 a_n3584_7550.t10 105.775
R126 a_n3584_7550.n0 a_n3584_7550.t9 105.775
R127 a_n3584_7550.n0 a_n3584_7550.t4 105.775
R128 a_n3584_7550.n0 a_n3584_7550.t13 105.775
R129 a_n3584_7550.n2 a_n3584_7550.t8 105.775
R130 a_n3584_7550.n3 a_n3584_7550.n7 98.1078
R131 a_n3584_7550.n0 a_n3584_7550.n5 98.1078
R132 a_n3584_7550.n0 a_n3584_7550.n6 98.1078
R133 a_n3584_7550.n2 a_n3584_7550.n4 98.1078
R134 a_n3584_7550.n1 a_n3584_7550.n2 25.6573
R135 a_n3584_7550.n1 a_n3584_7550.n0 13.0174
R136 a_n3584_7550.n1 a_n3584_7550.t0 10.5469
R137 a_n3584_7550.n3 a_n3584_7550.n1 8.40352
R138 a_n3584_7550.n7 a_n3584_7550.t16 7.66677
R139 a_n3584_7550.n7 a_n3584_7550.t2 7.66677
R140 a_n3584_7550.n5 a_n3584_7550.t12 7.66677
R141 a_n3584_7550.n5 a_n3584_7550.t6 7.66677
R142 a_n3584_7550.n6 a_n3584_7550.t7 7.66677
R143 a_n3584_7550.n6 a_n3584_7550.t14 7.66677
R144 a_n3584_7550.n4 a_n3584_7550.t15 7.66677
R145 a_n3584_7550.n4 a_n3584_7550.t11 7.66677
R146 a_n11986_8880.n22 a_n11986_8880.n27 74.9655
R147 a_n11986_8880.n23 a_n11986_8880.n24 28.5074
R148 a_n11986_8880.n4 a_n11986_8880.n25 28.3431
R149 a_n11986_8880.n18 a_n11986_8880.n28 74.9655
R150 a_n11986_8880.n19 a_n11986_8880.n20 28.5074
R151 a_n11986_8880.n7 a_n11986_8880.n21 28.3431
R152 a_n11986_8880.n17 a_n11986_8880.n10 28.3431
R153 a_n11986_8880.n2 a_n11986_8880.n3 12.6734
R154 a_n11986_8880.n16 a_n11986_8880.n13 28.3431
R155 a_n11986_8880.n0 a_n11986_8880.n1 12.6734
R156 a_n11986_8880.n31 a_n11986_8880.n29 127.225
R157 a_n11986_8880.n50 a_n11986_8880.n49 127.225
R158 a_n11986_8880.n49 a_n11986_8880.n48 126.035
R159 a_n11986_8880.n31 a_n11986_8880.n30 126.035
R160 a_n11986_8880.n26 a_n11986_8880.t0 93.0457
R161 a_n11986_8880.n33 a_n11986_8880.t5 93.0454
R162 a_n11986_8880.n33 a_n11986_8880.n32 87.706
R163 a_n11986_8880.n26 a_n11986_8880.n34 87.4336
R164 a_n11986_8880.n43 a_n11986_8880.n42 63.6066
R165 a_n11986_8880.n41 a_n11986_8880.n40 63.6066
R166 a_n11986_8880.n38 a_n11986_8880.n37 63.6066
R167 a_n11986_8880.n36 a_n11986_8880.n35 63.6066
R168 a_n11986_8880.n5 a_n11986_8880.n6 25.329
R169 a_n11986_8880.n8 a_n11986_8880.n9 25.329
R170 a_n11986_8880.n11 a_n11986_8880.n12 25.329
R171 a_n11986_8880.n14 a_n11986_8880.n15 25.329
R172 a_n11986_8880.n37 a_n11986_8880.t16 41.0691
R173 a_n11986_8880.n35 a_n11986_8880.t17 41.0691
R174 a_n11986_8880.n42 a_n11986_8880.t14 41.0687
R175 a_n11986_8880.n40 a_n11986_8880.t22 41.0687
R176 a_n11986_8880.n26 a_n11986_8880.n33 30.6721
R177 a_n11986_8880.n49 a_n11986_8880.n47 29.9047
R178 a_n11986_8880.n17 a_n11986_8880.n3 125.487
R179 a_n11986_8880.n16 a_n11986_8880.n1 125.487
R180 a_n11986_8880.n25 a_n11986_8880.n6 80.6698
R181 a_n11986_8880.n24 a_n11986_8880.n25 114.472
R182 a_n11986_8880.n24 a_n11986_8880.n27 65.1634
R183 a_n11986_8880.n43 a_n11986_8880.n27 23.6056
R184 a_n11986_8880.n21 a_n11986_8880.n9 80.6698
R185 a_n11986_8880.n20 a_n11986_8880.n21 114.472
R186 a_n11986_8880.n20 a_n11986_8880.n28 65.1634
R187 a_n11986_8880.n41 a_n11986_8880.n28 23.6056
R188 a_n11986_8880.n17 a_n11986_8880.n12 80.6698
R189 a_n11986_8880.n16 a_n11986_8880.n15 80.6698
R190 a_n11986_8880.n47 a_n11986_8880.n31 21.1173
R191 a_n11986_8880.n3 a_n11986_8880.n38 52.5736
R192 a_n11986_8880.n1 a_n11986_8880.n36 52.5736
R193 a_n11986_8880.n46 a_n11986_8880.n26 12.6334
R194 a_n11986_8880.n47 a_n11986_8880.n46 11.4887
R195 a_n11986_8880.n45 a_n11986_8880.n39 9.04282
R196 a_n11986_8880.n45 a_n11986_8880.n44 8.77084
R197 a_n11986_8880.n6 a_n11986_8880.t19 19.5352
R198 a_n11986_8880.n43 a_n11986_8880.t23 8.2528
R199 a_n11986_8880.n9 a_n11986_8880.t20 19.5352
R200 a_n11986_8880.n41 a_n11986_8880.t25 8.2528
R201 a_n11986_8880.n38 a_n11986_8880.t18 8.2528
R202 a_n11986_8880.n12 a_n11986_8880.t15 19.5352
R203 a_n11986_8880.n36 a_n11986_8880.t21 8.2528
R204 a_n11986_8880.n15 a_n11986_8880.t24 19.5352
R205 a_n11986_8880.n48 a_n11986_8880.t8 7.66677
R206 a_n11986_8880.n48 a_n11986_8880.t7 7.66677
R207 a_n11986_8880.n30 a_n11986_8880.t11 7.66677
R208 a_n11986_8880.n30 a_n11986_8880.t6 7.66677
R209 a_n11986_8880.n29 a_n11986_8880.t10 7.66677
R210 a_n11986_8880.n29 a_n11986_8880.t9 7.66677
R211 a_n11986_8880.n50 a_n11986_8880.t12 7.66677
R212 a_n11986_8880.t13 a_n11986_8880.n50 7.66677
R213 a_n11986_8880.n44 a_n11986_8880.n8 7.37588
R214 a_n11986_8880.n39 a_n11986_8880.n14 7.37588
R215 a_n11986_8880.n44 a_n11986_8880.n5 5.57285
R216 a_n11986_8880.n39 a_n11986_8880.n11 5.57285
R217 a_n11986_8880.n34 a_n11986_8880.t3 4.79469
R218 a_n11986_8880.n34 a_n11986_8880.t1 4.79469
R219 a_n11986_8880.n32 a_n11986_8880.t4 4.79469
R220 a_n11986_8880.n32 a_n11986_8880.t2 4.79469
R221 a_n11986_8880.n46 a_n11986_8880.n45 3.4105
R222 a_n11986_8880.n10 a_n11986_8880.n2 1.32626
R223 a_n11986_8880.n13 a_n11986_8880.n0 1.32626
R224 a_n11986_8880.n14 a_n11986_8880.n13 1.2602
R225 a_n11986_8880.n11 a_n11986_8880.n10 1.2602
R226 a_n11986_8880.n8 a_n11986_8880.n7 1.0708
R227 a_n11986_8880.n5 a_n11986_8880.n4 1.0708
R228 a_n11986_8880.n2 a_n11986_8880.n37 0.986657
R229 a_n11986_8880.n0 a_n11986_8880.n35 0.986657
R230 a_n11986_8880.n22 a_n11986_8880.n42 0.986652
R231 a_n11986_8880.n18 a_n11986_8880.n40 0.986652
R232 a_n11986_8880.n4 a_n11986_8880.n23 0.758076
R233 a_n11986_8880.n23 a_n11986_8880.n22 0.758076
R234 a_n11986_8880.n7 a_n11986_8880.n19 0.758076
R235 a_n11986_8880.n19 a_n11986_8880.n18 0.758076
R236 VDD.n28 VDD.n26 756.745
R237 VDD.n19 VDD.n17 756.745
R238 VDD.n1112 VDD.n1110 756.745
R239 VDD.n1103 VDD.n1101 756.745
R240 VDD.n29 VDD.n28 585
R241 VDD.n20 VDD.n19 585
R242 VDD.n1113 VDD.n1112 585
R243 VDD.n1104 VDD.n1103 585
R244 VDD.t63 VDD.n27 417.779
R245 VDD.t74 VDD.n18 417.779
R246 VDD.t60 VDD.n1111 417.779
R247 VDD.t73 VDD.n1102 417.779
R248 VDD.n2709 VDD.n127 411.221
R249 VDD.n156 VDD.n129 411.221
R250 VDD.n2475 VDD.n275 411.221
R251 VDD.n2473 VDD.n2402 411.221
R252 VDD.n1253 VDD.n699 411.221
R253 VDD.n1317 VDD.n689 411.221
R254 VDD.n965 VDD.n894 411.221
R255 VDD.n967 VDD.n892 411.221
R256 VDD.n898 VDD.t48 368.774
R257 VDD.n913 VDD.t11 368.774
R258 VDD.n2414 VDD.t22 368.774
R259 VDD.n2433 VDD.t35 368.774
R260 VDD.n158 VDD.t6 368.774
R261 VDD.n2690 VDD.t13 368.774
R262 VDD.n1264 VDD.t2 368.774
R263 VDD.n690 VDD.t31 368.774
R264 VDD.n2133 VDD.n1863 305.854
R265 VDD.n2399 VDD.n298 305.854
R266 VDD.n2358 VDD.n2357 305.854
R267 VDD.n2092 VDD.n1860 305.854
R268 VDD.n1857 VDD.n498 305.854
R269 VDD.n1816 VDD.n1815 305.854
R270 VDD.n1550 VDD.n1320 305.854
R271 VDD.n1591 VDD.n1452 305.854
R272 VDD.n2343 VDD.n277 305.854
R273 VDD.n2301 VDD.n2300 305.854
R274 VDD.n1984 VDD.n1861 305.854
R275 VDD.n2135 VDD.n475 305.854
R276 VDD.n1801 VDD.n477 305.854
R277 VDD.n1759 VDD.n1758 305.854
R278 VDD.n1451 VDD.n1321 305.854
R279 VDD.n1593 VDD.n677 305.854
R280 VDD.n1874 VDD.t15 249.827
R281 VDD.n301 VDD.t23 249.827
R282 VDD.n1463 VDD.t53 249.827
R283 VDD.n501 VDD.t43 249.827
R284 VDD.n1935 VDD.t36 249.827
R285 VDD.n318 VDD.t27 249.827
R286 VDD.n1324 VDD.t49 249.827
R287 VDD.n518 VDD.t39 249.827
R288 VDD.n899 VDD.t47 248.531
R289 VDD.n914 VDD.t10 248.531
R290 VDD.n2415 VDD.t21 248.531
R291 VDD.n2434 VDD.t34 248.531
R292 VDD.n159 VDD.t7 248.531
R293 VDD.n2691 VDD.t14 248.531
R294 VDD.n1265 VDD.t3 248.531
R295 VDD.n691 VDD.t32 248.531
R296 VDD.n898 VDD.t46 210.659
R297 VDD.n913 VDD.t8 210.659
R298 VDD.n2414 VDD.t19 210.659
R299 VDD.n2433 VDD.t33 210.659
R300 VDD.n158 VDD.t4 210.659
R301 VDD.n2690 VDD.t12 210.659
R302 VDD.n1264 VDD.t0 210.659
R303 VDD.n690 VDD.t30 210.659
R304 VDD.n33 VDD.n25 192.643
R305 VDD.n24 VDD.n16 192.643
R306 VDD.t115 VDD.n1318 192.27
R307 VDD.n2401 VDD.t56 192.27
R308 VDD.n1118 VDD.n1117 189.97
R309 VDD.n1109 VDD.n1108 189.97
R310 VDD.n1802 VDD.n1801 185
R311 VDD.n1801 VDD.n476 185
R312 VDD.n1803 VDD.n507 185
R313 VDD.n1813 VDD.n507 185
R314 VDD.n1804 VDD.n516 185
R315 VDD.n516 VDD.n514 185
R316 VDD.n1806 VDD.n1805 185
R317 VDD.n1807 VDD.n1806 185
R318 VDD.n517 VDD.n515 185
R319 VDD.n515 VDD.n511 185
R320 VDD.n1740 VDD.n523 185
R321 VDD.t40 VDD.n523 185
R322 VDD.n1741 VDD.n532 185
R323 VDD.n532 VDD.n522 185
R324 VDD.n1743 VDD.n1742 185
R325 VDD.n1744 VDD.n1743 185
R326 VDD.n1739 VDD.n531 185
R327 VDD.n531 VDD.n528 185
R328 VDD.n1738 VDD.n1737 185
R329 VDD.n1737 VDD.n1736 185
R330 VDD.n534 VDD.n533 185
R331 VDD.n543 VDD.n534 185
R332 VDD.n1729 VDD.n1728 185
R333 VDD.n1730 VDD.n1729 185
R334 VDD.n1727 VDD.n544 185
R335 VDD.n544 VDD.n540 185
R336 VDD.n1726 VDD.n1725 185
R337 VDD.n1725 VDD.n1724 185
R338 VDD.n546 VDD.n545 185
R339 VDD.n547 VDD.n546 185
R340 VDD.n1717 VDD.n1716 185
R341 VDD.n1718 VDD.n1717 185
R342 VDD.n1715 VDD.n556 185
R343 VDD.n556 VDD.n553 185
R344 VDD.n1714 VDD.n1713 185
R345 VDD.n1713 VDD.n1712 185
R346 VDD.n558 VDD.n557 185
R347 VDD.n567 VDD.n558 185
R348 VDD.n1705 VDD.n1704 185
R349 VDD.n1706 VDD.n1705 185
R350 VDD.n1703 VDD.n568 185
R351 VDD.n568 VDD.n564 185
R352 VDD.n1702 VDD.n1701 185
R353 VDD.n1701 VDD.n1700 185
R354 VDD.n570 VDD.n569 185
R355 VDD.n571 VDD.n570 185
R356 VDD.n1693 VDD.n1692 185
R357 VDD.n1694 VDD.n1693 185
R358 VDD.n1691 VDD.n580 185
R359 VDD.n580 VDD.n577 185
R360 VDD.n1690 VDD.n1689 185
R361 VDD.n1689 VDD.n1688 185
R362 VDD.n582 VDD.n581 185
R363 VDD.n583 VDD.n582 185
R364 VDD.n1681 VDD.n1680 185
R365 VDD.n1682 VDD.n1681 185
R366 VDD.n1679 VDD.n592 185
R367 VDD.n592 VDD.n589 185
R368 VDD.n1678 VDD.n1677 185
R369 VDD.n1677 VDD.n1676 185
R370 VDD.n594 VDD.n593 185
R371 VDD.n595 VDD.n594 185
R372 VDD.n1669 VDD.n1668 185
R373 VDD.n1670 VDD.n1669 185
R374 VDD.n1667 VDD.n604 185
R375 VDD.n604 VDD.n601 185
R376 VDD.n1666 VDD.n1665 185
R377 VDD.n1665 VDD.n1664 185
R378 VDD.n606 VDD.n605 185
R379 VDD.n607 VDD.n606 185
R380 VDD.n1657 VDD.n1656 185
R381 VDD.n1658 VDD.n1657 185
R382 VDD.n1655 VDD.n616 185
R383 VDD.n616 VDD.n613 185
R384 VDD.n1654 VDD.n1653 185
R385 VDD.n1653 VDD.n1652 185
R386 VDD.n618 VDD.n617 185
R387 VDD.n619 VDD.n618 185
R388 VDD.n1645 VDD.n1644 185
R389 VDD.n1646 VDD.n1645 185
R390 VDD.n1643 VDD.n628 185
R391 VDD.n628 VDD.n625 185
R392 VDD.n1642 VDD.n1641 185
R393 VDD.n1641 VDD.n1640 185
R394 VDD.n630 VDD.n629 185
R395 VDD.n631 VDD.n630 185
R396 VDD.n1633 VDD.n1632 185
R397 VDD.n1634 VDD.n1633 185
R398 VDD.n1631 VDD.n640 185
R399 VDD.n640 VDD.n637 185
R400 VDD.n1630 VDD.n1629 185
R401 VDD.n1629 VDD.n1628 185
R402 VDD.n642 VDD.n641 185
R403 VDD.n643 VDD.n642 185
R404 VDD.n1621 VDD.n1620 185
R405 VDD.n1622 VDD.n1621 185
R406 VDD.n1619 VDD.n652 185
R407 VDD.n652 VDD.n649 185
R408 VDD.n1618 VDD.n1617 185
R409 VDD.n1617 VDD.n1616 185
R410 VDD.n654 VDD.n653 185
R411 VDD.n655 VDD.n654 185
R412 VDD.n1609 VDD.n1608 185
R413 VDD.n1610 VDD.n1609 185
R414 VDD.n1607 VDD.n663 185
R415 VDD.n663 VDD.t50 185
R416 VDD.n1606 VDD.n1605 185
R417 VDD.n1605 VDD.n1604 185
R418 VDD.n665 VDD.n664 185
R419 VDD.n666 VDD.n665 185
R420 VDD.n1597 VDD.n1596 185
R421 VDD.n1598 VDD.n1597 185
R422 VDD.n1595 VDD.n675 185
R423 VDD.n675 VDD.n672 185
R424 VDD.n1594 VDD.n1593 185
R425 VDD.n1593 VDD.n1592 185
R426 VDD.n677 VDD.n676 185
R427 VDD.n1337 VDD.n1335 185
R428 VDD.n1340 VDD.n1339 185
R429 VDD.n1341 VDD.n1334 185
R430 VDD.n1343 VDD.n1342 185
R431 VDD.n1345 VDD.n1333 185
R432 VDD.n1348 VDD.n1347 185
R433 VDD.n1349 VDD.n1332 185
R434 VDD.n1351 VDD.n1350 185
R435 VDD.n1353 VDD.n1331 185
R436 VDD.n1356 VDD.n1355 185
R437 VDD.n1357 VDD.n1330 185
R438 VDD.n1359 VDD.n1358 185
R439 VDD.n1361 VDD.n1329 185
R440 VDD.n1364 VDD.n1363 185
R441 VDD.n1365 VDD.n1328 185
R442 VDD.n1367 VDD.n1366 185
R443 VDD.n1369 VDD.n1327 185
R444 VDD.n1370 VDD.n1323 185
R445 VDD.n1373 VDD.n1372 185
R446 VDD.n1374 VDD.n1321 185
R447 VDD.n1321 VDD.n1319 185
R448 VDD.n1760 VDD.n1759 185
R449 VDD.n1762 VDD.n1761 185
R450 VDD.n1764 VDD.n1763 185
R451 VDD.n1767 VDD.n1766 185
R452 VDD.n1769 VDD.n1768 185
R453 VDD.n1771 VDD.n1770 185
R454 VDD.n1773 VDD.n1772 185
R455 VDD.n1775 VDD.n1774 185
R456 VDD.n1777 VDD.n1776 185
R457 VDD.n1779 VDD.n1778 185
R458 VDD.n1781 VDD.n1780 185
R459 VDD.n1783 VDD.n1782 185
R460 VDD.n1785 VDD.n1784 185
R461 VDD.n1787 VDD.n1786 185
R462 VDD.n1789 VDD.n1788 185
R463 VDD.n1791 VDD.n1790 185
R464 VDD.n1793 VDD.n1792 185
R465 VDD.n1795 VDD.n1794 185
R466 VDD.n1797 VDD.n1796 185
R467 VDD.n1799 VDD.n1798 185
R468 VDD.n1800 VDD.n477 185
R469 VDD.n1858 VDD.n477 185
R470 VDD.n1758 VDD.n1757 185
R471 VDD.n1758 VDD.n476 185
R472 VDD.n1756 VDD.n506 185
R473 VDD.n1813 VDD.n506 185
R474 VDD.n1755 VDD.n1754 185
R475 VDD.n1754 VDD.n514 185
R476 VDD.n1753 VDD.n513 185
R477 VDD.n1807 VDD.n513 185
R478 VDD.n1752 VDD.n1751 185
R479 VDD.n1751 VDD.n511 185
R480 VDD.n1750 VDD.n520 185
R481 VDD.n1750 VDD.t40 185
R482 VDD.n1375 VDD.n521 185
R483 VDD.n522 VDD.n521 185
R484 VDD.n1376 VDD.n530 185
R485 VDD.n1744 VDD.n530 185
R486 VDD.n1378 VDD.n1377 185
R487 VDD.n1377 VDD.n528 185
R488 VDD.n1379 VDD.n536 185
R489 VDD.n1736 VDD.n536 185
R490 VDD.n1381 VDD.n1380 185
R491 VDD.n1380 VDD.n543 185
R492 VDD.n1382 VDD.n542 185
R493 VDD.n1730 VDD.n542 185
R494 VDD.n1384 VDD.n1383 185
R495 VDD.n1383 VDD.n540 185
R496 VDD.n1385 VDD.n549 185
R497 VDD.n1724 VDD.n549 185
R498 VDD.n1387 VDD.n1386 185
R499 VDD.n1386 VDD.n547 185
R500 VDD.n1388 VDD.n555 185
R501 VDD.n1718 VDD.n555 185
R502 VDD.n1390 VDD.n1389 185
R503 VDD.n1389 VDD.n553 185
R504 VDD.n1391 VDD.n560 185
R505 VDD.n1712 VDD.n560 185
R506 VDD.n1393 VDD.n1392 185
R507 VDD.n1392 VDD.n567 185
R508 VDD.n1394 VDD.n566 185
R509 VDD.n1706 VDD.n566 185
R510 VDD.n1396 VDD.n1395 185
R511 VDD.n1395 VDD.n564 185
R512 VDD.n1397 VDD.n573 185
R513 VDD.n1700 VDD.n573 185
R514 VDD.n1399 VDD.n1398 185
R515 VDD.n1398 VDD.n571 185
R516 VDD.n1400 VDD.n579 185
R517 VDD.n1694 VDD.n579 185
R518 VDD.n1402 VDD.n1401 185
R519 VDD.n1401 VDD.n577 185
R520 VDD.n1403 VDD.n585 185
R521 VDD.n1688 VDD.n585 185
R522 VDD.n1405 VDD.n1404 185
R523 VDD.n1404 VDD.n583 185
R524 VDD.n1406 VDD.n591 185
R525 VDD.n1682 VDD.n591 185
R526 VDD.n1408 VDD.n1407 185
R527 VDD.n1407 VDD.n589 185
R528 VDD.n1409 VDD.n597 185
R529 VDD.n1676 VDD.n597 185
R530 VDD.n1411 VDD.n1410 185
R531 VDD.n1410 VDD.n595 185
R532 VDD.n1412 VDD.n603 185
R533 VDD.n1670 VDD.n603 185
R534 VDD.n1414 VDD.n1413 185
R535 VDD.n1413 VDD.n601 185
R536 VDD.n1415 VDD.n609 185
R537 VDD.n1664 VDD.n609 185
R538 VDD.n1417 VDD.n1416 185
R539 VDD.n1416 VDD.n607 185
R540 VDD.n1418 VDD.n615 185
R541 VDD.n1658 VDD.n615 185
R542 VDD.n1420 VDD.n1419 185
R543 VDD.n1419 VDD.n613 185
R544 VDD.n1421 VDD.n621 185
R545 VDD.n1652 VDD.n621 185
R546 VDD.n1423 VDD.n1422 185
R547 VDD.n1422 VDD.n619 185
R548 VDD.n1424 VDD.n627 185
R549 VDD.n1646 VDD.n627 185
R550 VDD.n1426 VDD.n1425 185
R551 VDD.n1425 VDD.n625 185
R552 VDD.n1427 VDD.n633 185
R553 VDD.n1640 VDD.n633 185
R554 VDD.n1429 VDD.n1428 185
R555 VDD.n1428 VDD.n631 185
R556 VDD.n1430 VDD.n639 185
R557 VDD.n1634 VDD.n639 185
R558 VDD.n1432 VDD.n1431 185
R559 VDD.n1431 VDD.n637 185
R560 VDD.n1433 VDD.n645 185
R561 VDD.n1628 VDD.n645 185
R562 VDD.n1435 VDD.n1434 185
R563 VDD.n1434 VDD.n643 185
R564 VDD.n1436 VDD.n651 185
R565 VDD.n1622 VDD.n651 185
R566 VDD.n1438 VDD.n1437 185
R567 VDD.n1437 VDD.n649 185
R568 VDD.n1439 VDD.n657 185
R569 VDD.n1616 VDD.n657 185
R570 VDD.n1441 VDD.n1440 185
R571 VDD.n1440 VDD.n655 185
R572 VDD.n1442 VDD.n662 185
R573 VDD.n1610 VDD.n662 185
R574 VDD.n1444 VDD.n1443 185
R575 VDD.n1443 VDD.t50 185
R576 VDD.n1445 VDD.n668 185
R577 VDD.n1604 VDD.n668 185
R578 VDD.n1447 VDD.n1446 185
R579 VDD.n1446 VDD.n666 185
R580 VDD.n1448 VDD.n674 185
R581 VDD.n1598 VDD.n674 185
R582 VDD.n1449 VDD.n1322 185
R583 VDD.n1322 VDD.n672 185
R584 VDD.n1451 VDD.n1450 185
R585 VDD.n1592 VDD.n1451 185
R586 VDD.n2344 VDD.n2343 185
R587 VDD.n2343 VDD.n276 185
R588 VDD.n2345 VDD.n308 185
R589 VDD.n2355 VDD.n308 185
R590 VDD.n2346 VDD.n316 185
R591 VDD.n316 VDD.n306 185
R592 VDD.n2348 VDD.n2347 185
R593 VDD.n2349 VDD.n2348 185
R594 VDD.n317 VDD.n315 185
R595 VDD.n315 VDD.n312 185
R596 VDD.n2282 VDD.n323 185
R597 VDD.t24 VDD.n323 185
R598 VDD.n2283 VDD.n332 185
R599 VDD.n332 VDD.n322 185
R600 VDD.n2285 VDD.n2284 185
R601 VDD.n2286 VDD.n2285 185
R602 VDD.n2281 VDD.n331 185
R603 VDD.n331 VDD.n328 185
R604 VDD.n2280 VDD.n2279 185
R605 VDD.n2279 VDD.n2278 185
R606 VDD.n334 VDD.n333 185
R607 VDD.n335 VDD.n334 185
R608 VDD.n2271 VDD.n2270 185
R609 VDD.n2272 VDD.n2271 185
R610 VDD.n2269 VDD.n344 185
R611 VDD.n344 VDD.n341 185
R612 VDD.n2268 VDD.n2267 185
R613 VDD.n2267 VDD.n2266 185
R614 VDD.n346 VDD.n345 185
R615 VDD.n347 VDD.n346 185
R616 VDD.n2259 VDD.n2258 185
R617 VDD.n2260 VDD.n2259 185
R618 VDD.n2257 VDD.n356 185
R619 VDD.n356 VDD.n353 185
R620 VDD.n2256 VDD.n2255 185
R621 VDD.n2255 VDD.n2254 185
R622 VDD.n358 VDD.n357 185
R623 VDD.n359 VDD.n358 185
R624 VDD.n2247 VDD.n2246 185
R625 VDD.n2248 VDD.n2247 185
R626 VDD.n2245 VDD.n368 185
R627 VDD.n368 VDD.n365 185
R628 VDD.n2244 VDD.n2243 185
R629 VDD.n2243 VDD.n2242 185
R630 VDD.n370 VDD.n369 185
R631 VDD.n371 VDD.n370 185
R632 VDD.n2235 VDD.n2234 185
R633 VDD.n2236 VDD.n2235 185
R634 VDD.n2233 VDD.n380 185
R635 VDD.n380 VDD.n377 185
R636 VDD.n2232 VDD.n2231 185
R637 VDD.n2231 VDD.n2230 185
R638 VDD.n382 VDD.n381 185
R639 VDD.n383 VDD.n382 185
R640 VDD.n2223 VDD.n2222 185
R641 VDD.n2224 VDD.n2223 185
R642 VDD.n2221 VDD.n392 185
R643 VDD.n392 VDD.n389 185
R644 VDD.n2220 VDD.n2219 185
R645 VDD.n2219 VDD.n2218 185
R646 VDD.n394 VDD.n393 185
R647 VDD.n395 VDD.n394 185
R648 VDD.n2211 VDD.n2210 185
R649 VDD.n2212 VDD.n2211 185
R650 VDD.n2209 VDD.n404 185
R651 VDD.n404 VDD.n401 185
R652 VDD.n2208 VDD.n2207 185
R653 VDD.n2207 VDD.n2206 185
R654 VDD.n406 VDD.n405 185
R655 VDD.n407 VDD.n406 185
R656 VDD.n2199 VDD.n2198 185
R657 VDD.n2200 VDD.n2199 185
R658 VDD.n2197 VDD.n416 185
R659 VDD.n416 VDD.n413 185
R660 VDD.n2196 VDD.n2195 185
R661 VDD.n2195 VDD.n2194 185
R662 VDD.n418 VDD.n417 185
R663 VDD.n419 VDD.n418 185
R664 VDD.n2187 VDD.n2186 185
R665 VDD.n2188 VDD.n2187 185
R666 VDD.n2185 VDD.n427 185
R667 VDD.n2063 VDD.n427 185
R668 VDD.n2184 VDD.n2183 185
R669 VDD.n2183 VDD.n2182 185
R670 VDD.n429 VDD.n428 185
R671 VDD.n430 VDD.n429 185
R672 VDD.n2175 VDD.n2174 185
R673 VDD.n2176 VDD.n2175 185
R674 VDD.n2173 VDD.n439 185
R675 VDD.n439 VDD.n436 185
R676 VDD.n2172 VDD.n2171 185
R677 VDD.n2171 VDD.n2170 185
R678 VDD.n441 VDD.n440 185
R679 VDD.n442 VDD.n441 185
R680 VDD.n2163 VDD.n2162 185
R681 VDD.n2164 VDD.n2163 185
R682 VDD.n2161 VDD.n450 185
R683 VDD.n456 VDD.n450 185
R684 VDD.n2160 VDD.n2159 185
R685 VDD.n2159 VDD.n2158 185
R686 VDD.n452 VDD.n451 185
R687 VDD.n453 VDD.n452 185
R688 VDD.n2151 VDD.n2150 185
R689 VDD.n2152 VDD.n2151 185
R690 VDD.n2149 VDD.n462 185
R691 VDD.n462 VDD.t16 185
R692 VDD.n2148 VDD.n2147 185
R693 VDD.n2147 VDD.n2146 185
R694 VDD.n464 VDD.n463 185
R695 VDD.n465 VDD.n464 185
R696 VDD.n2139 VDD.n2138 185
R697 VDD.n2140 VDD.n2139 185
R698 VDD.n2137 VDD.n473 185
R699 VDD.n1862 VDD.n473 185
R700 VDD.n2136 VDD.n2135 185
R701 VDD.n2135 VDD.n2134 185
R702 VDD.n475 VDD.n474 185
R703 VDD.n1946 VDD.n1945 185
R704 VDD.n1948 VDD.n1947 185
R705 VDD.n1950 VDD.n1943 185
R706 VDD.n1953 VDD.n1952 185
R707 VDD.n1954 VDD.n1942 185
R708 VDD.n1956 VDD.n1955 185
R709 VDD.n1958 VDD.n1941 185
R710 VDD.n1961 VDD.n1960 185
R711 VDD.n1962 VDD.n1940 185
R712 VDD.n1964 VDD.n1963 185
R713 VDD.n1966 VDD.n1939 185
R714 VDD.n1969 VDD.n1968 185
R715 VDD.n1970 VDD.n1938 185
R716 VDD.n1972 VDD.n1971 185
R717 VDD.n1974 VDD.n1937 185
R718 VDD.n1977 VDD.n1976 185
R719 VDD.n1978 VDD.n1934 185
R720 VDD.n1981 VDD.n1980 185
R721 VDD.n1983 VDD.n1933 185
R722 VDD.n1985 VDD.n1984 185
R723 VDD.n1984 VDD.n1859 185
R724 VDD.n2302 VDD.n2301 185
R725 VDD.n2304 VDD.n2303 185
R726 VDD.n2306 VDD.n2305 185
R727 VDD.n2309 VDD.n2308 185
R728 VDD.n2311 VDD.n2310 185
R729 VDD.n2313 VDD.n2312 185
R730 VDD.n2315 VDD.n2314 185
R731 VDD.n2317 VDD.n2316 185
R732 VDD.n2319 VDD.n2318 185
R733 VDD.n2321 VDD.n2320 185
R734 VDD.n2323 VDD.n2322 185
R735 VDD.n2325 VDD.n2324 185
R736 VDD.n2327 VDD.n2326 185
R737 VDD.n2329 VDD.n2328 185
R738 VDD.n2331 VDD.n2330 185
R739 VDD.n2333 VDD.n2332 185
R740 VDD.n2335 VDD.n2334 185
R741 VDD.n2337 VDD.n2336 185
R742 VDD.n2339 VDD.n2338 185
R743 VDD.n2341 VDD.n2340 185
R744 VDD.n2342 VDD.n277 185
R745 VDD.n2400 VDD.n277 185
R746 VDD.n2300 VDD.n2299 185
R747 VDD.n2300 VDD.n276 185
R748 VDD.n2298 VDD.n307 185
R749 VDD.n2355 VDD.n307 185
R750 VDD.n2297 VDD.n2296 185
R751 VDD.n2296 VDD.n306 185
R752 VDD.n2295 VDD.n314 185
R753 VDD.n2349 VDD.n314 185
R754 VDD.n2294 VDD.n2293 185
R755 VDD.n2293 VDD.n312 185
R756 VDD.n2292 VDD.n320 185
R757 VDD.n2292 VDD.t24 185
R758 VDD.n2011 VDD.n321 185
R759 VDD.n322 VDD.n321 185
R760 VDD.n2012 VDD.n330 185
R761 VDD.n2286 VDD.n330 185
R762 VDD.n2014 VDD.n2013 185
R763 VDD.n2013 VDD.n328 185
R764 VDD.n2015 VDD.n337 185
R765 VDD.n2278 VDD.n337 185
R766 VDD.n2017 VDD.n2016 185
R767 VDD.n2016 VDD.n335 185
R768 VDD.n2018 VDD.n343 185
R769 VDD.n2272 VDD.n343 185
R770 VDD.n2020 VDD.n2019 185
R771 VDD.n2019 VDD.n341 185
R772 VDD.n2021 VDD.n349 185
R773 VDD.n2266 VDD.n349 185
R774 VDD.n2023 VDD.n2022 185
R775 VDD.n2022 VDD.n347 185
R776 VDD.n2024 VDD.n355 185
R777 VDD.n2260 VDD.n355 185
R778 VDD.n2026 VDD.n2025 185
R779 VDD.n2025 VDD.n353 185
R780 VDD.n2027 VDD.n361 185
R781 VDD.n2254 VDD.n361 185
R782 VDD.n2029 VDD.n2028 185
R783 VDD.n2028 VDD.n359 185
R784 VDD.n2030 VDD.n367 185
R785 VDD.n2248 VDD.n367 185
R786 VDD.n2032 VDD.n2031 185
R787 VDD.n2031 VDD.n365 185
R788 VDD.n2033 VDD.n373 185
R789 VDD.n2242 VDD.n373 185
R790 VDD.n2035 VDD.n2034 185
R791 VDD.n2034 VDD.n371 185
R792 VDD.n2036 VDD.n379 185
R793 VDD.n2236 VDD.n379 185
R794 VDD.n2038 VDD.n2037 185
R795 VDD.n2037 VDD.n377 185
R796 VDD.n2039 VDD.n385 185
R797 VDD.n2230 VDD.n385 185
R798 VDD.n2041 VDD.n2040 185
R799 VDD.n2040 VDD.n383 185
R800 VDD.n2042 VDD.n391 185
R801 VDD.n2224 VDD.n391 185
R802 VDD.n2044 VDD.n2043 185
R803 VDD.n2043 VDD.n389 185
R804 VDD.n2045 VDD.n397 185
R805 VDD.n2218 VDD.n397 185
R806 VDD.n2047 VDD.n2046 185
R807 VDD.n2046 VDD.n395 185
R808 VDD.n2048 VDD.n403 185
R809 VDD.n2212 VDD.n403 185
R810 VDD.n2050 VDD.n2049 185
R811 VDD.n2049 VDD.n401 185
R812 VDD.n2051 VDD.n409 185
R813 VDD.n2206 VDD.n409 185
R814 VDD.n2053 VDD.n2052 185
R815 VDD.n2052 VDD.n407 185
R816 VDD.n2054 VDD.n415 185
R817 VDD.n2200 VDD.n415 185
R818 VDD.n2056 VDD.n2055 185
R819 VDD.n2055 VDD.n413 185
R820 VDD.n2057 VDD.n421 185
R821 VDD.n2194 VDD.n421 185
R822 VDD.n2059 VDD.n2058 185
R823 VDD.n2058 VDD.n419 185
R824 VDD.n2060 VDD.n426 185
R825 VDD.n2188 VDD.n426 185
R826 VDD.n2062 VDD.n2061 185
R827 VDD.n2063 VDD.n2062 185
R828 VDD.n2010 VDD.n432 185
R829 VDD.n2182 VDD.n432 185
R830 VDD.n2009 VDD.n2008 185
R831 VDD.n2008 VDD.n430 185
R832 VDD.n2007 VDD.n438 185
R833 VDD.n2176 VDD.n438 185
R834 VDD.n2006 VDD.n2005 185
R835 VDD.n2005 VDD.n436 185
R836 VDD.n2004 VDD.n444 185
R837 VDD.n2170 VDD.n444 185
R838 VDD.n2003 VDD.n2002 185
R839 VDD.n2002 VDD.n442 185
R840 VDD.n2001 VDD.n449 185
R841 VDD.n2164 VDD.n449 185
R842 VDD.n2000 VDD.n1999 185
R843 VDD.n1999 VDD.n456 185
R844 VDD.n1998 VDD.n455 185
R845 VDD.n2158 VDD.n455 185
R846 VDD.n1997 VDD.n1996 185
R847 VDD.n1996 VDD.n453 185
R848 VDD.n1995 VDD.n461 185
R849 VDD.n2152 VDD.n461 185
R850 VDD.n1994 VDD.n1993 185
R851 VDD.n1993 VDD.t16 185
R852 VDD.n1992 VDD.n467 185
R853 VDD.n2146 VDD.n467 185
R854 VDD.n1991 VDD.n1990 185
R855 VDD.n1990 VDD.n465 185
R856 VDD.n1989 VDD.n472 185
R857 VDD.n2140 VDD.n472 185
R858 VDD.n1988 VDD.n1987 185
R859 VDD.n1987 VDD.n1862 185
R860 VDD.n1986 VDD.n1861 185
R861 VDD.n2134 VDD.n1861 185
R862 VDD.n500 VDD.n498 185
R863 VDD.n498 VDD.n476 185
R864 VDD.n1812 VDD.n1811 185
R865 VDD.n1813 VDD.n1812 185
R866 VDD.n1810 VDD.n508 185
R867 VDD.n514 VDD.n508 185
R868 VDD.n1809 VDD.n1808 185
R869 VDD.n1808 VDD.n1807 185
R870 VDD.n510 VDD.n509 185
R871 VDD.n511 VDD.n510 185
R872 VDD.n1749 VDD.n1748 185
R873 VDD.t40 VDD.n1749 185
R874 VDD.n1747 VDD.n525 185
R875 VDD.n525 VDD.n522 185
R876 VDD.n1746 VDD.n1745 185
R877 VDD.n1745 VDD.n1744 185
R878 VDD.n527 VDD.n526 185
R879 VDD.n528 VDD.n527 185
R880 VDD.n1735 VDD.n1734 185
R881 VDD.n1736 VDD.n1735 185
R882 VDD.n1733 VDD.n537 185
R883 VDD.n543 VDD.n537 185
R884 VDD.n1732 VDD.n1731 185
R885 VDD.n1731 VDD.n1730 185
R886 VDD.n539 VDD.n538 185
R887 VDD.n540 VDD.n539 185
R888 VDD.n1723 VDD.n1722 185
R889 VDD.n1724 VDD.n1723 185
R890 VDD.n1721 VDD.n550 185
R891 VDD.n550 VDD.n547 185
R892 VDD.n1720 VDD.n1719 185
R893 VDD.n1719 VDD.n1718 185
R894 VDD.n552 VDD.n551 185
R895 VDD.n553 VDD.n552 185
R896 VDD.n1711 VDD.n1710 185
R897 VDD.n1712 VDD.n1711 185
R898 VDD.n1709 VDD.n561 185
R899 VDD.n567 VDD.n561 185
R900 VDD.n1708 VDD.n1707 185
R901 VDD.n1707 VDD.n1706 185
R902 VDD.n563 VDD.n562 185
R903 VDD.n564 VDD.n563 185
R904 VDD.n1699 VDD.n1698 185
R905 VDD.n1700 VDD.n1699 185
R906 VDD.n1697 VDD.n574 185
R907 VDD.n574 VDD.n571 185
R908 VDD.n1696 VDD.n1695 185
R909 VDD.n1695 VDD.n1694 185
R910 VDD.n576 VDD.n575 185
R911 VDD.n577 VDD.n576 185
R912 VDD.n1687 VDD.n1686 185
R913 VDD.n1688 VDD.n1687 185
R914 VDD.n1685 VDD.n586 185
R915 VDD.n586 VDD.n583 185
R916 VDD.n1684 VDD.n1683 185
R917 VDD.n1683 VDD.n1682 185
R918 VDD.n588 VDD.n587 185
R919 VDD.n589 VDD.n588 185
R920 VDD.n1675 VDD.n1674 185
R921 VDD.n1676 VDD.n1675 185
R922 VDD.n1673 VDD.n598 185
R923 VDD.n598 VDD.n595 185
R924 VDD.n1672 VDD.n1671 185
R925 VDD.n1671 VDD.n1670 185
R926 VDD.n600 VDD.n599 185
R927 VDD.n601 VDD.n600 185
R928 VDD.n1663 VDD.n1662 185
R929 VDD.n1664 VDD.n1663 185
R930 VDD.n1661 VDD.n610 185
R931 VDD.n610 VDD.n607 185
R932 VDD.n1660 VDD.n1659 185
R933 VDD.n1659 VDD.n1658 185
R934 VDD.n612 VDD.n611 185
R935 VDD.n613 VDD.n612 185
R936 VDD.n1651 VDD.n1650 185
R937 VDD.n1652 VDD.n1651 185
R938 VDD.n1649 VDD.n622 185
R939 VDD.n622 VDD.n619 185
R940 VDD.n1648 VDD.n1647 185
R941 VDD.n1647 VDD.n1646 185
R942 VDD.n624 VDD.n623 185
R943 VDD.n625 VDD.n624 185
R944 VDD.n1639 VDD.n1638 185
R945 VDD.n1640 VDD.n1639 185
R946 VDD.n1637 VDD.n634 185
R947 VDD.n634 VDD.n631 185
R948 VDD.n1636 VDD.n1635 185
R949 VDD.n1635 VDD.n1634 185
R950 VDD.n636 VDD.n635 185
R951 VDD.n637 VDD.n636 185
R952 VDD.n1627 VDD.n1626 185
R953 VDD.n1628 VDD.n1627 185
R954 VDD.n1625 VDD.n646 185
R955 VDD.n646 VDD.n643 185
R956 VDD.n1624 VDD.n1623 185
R957 VDD.n1623 VDD.n1622 185
R958 VDD.n648 VDD.n647 185
R959 VDD.n649 VDD.n648 185
R960 VDD.n1615 VDD.n1614 185
R961 VDD.n1616 VDD.n1615 185
R962 VDD.n1613 VDD.n658 185
R963 VDD.n658 VDD.n655 185
R964 VDD.n1612 VDD.n1611 185
R965 VDD.n1611 VDD.n1610 185
R966 VDD.n660 VDD.n659 185
R967 VDD.t50 VDD.n660 185
R968 VDD.n1603 VDD.n1602 185
R969 VDD.n1604 VDD.n1603 185
R970 VDD.n1601 VDD.n669 185
R971 VDD.n669 VDD.n666 185
R972 VDD.n1600 VDD.n1599 185
R973 VDD.n1599 VDD.n1598 185
R974 VDD.n671 VDD.n670 185
R975 VDD.n672 VDD.n671 185
R976 VDD.n1591 VDD.n1590 185
R977 VDD.n1592 VDD.n1591 185
R978 VDD.n1589 VDD.n1452 185
R979 VDD.n1588 VDD.n1587 185
R980 VDD.n1585 VDD.n1453 185
R981 VDD.n1585 VDD.n1319 185
R982 VDD.n1584 VDD.n1583 185
R983 VDD.n1582 VDD.n1581 185
R984 VDD.n1580 VDD.n1455 185
R985 VDD.n1578 VDD.n1577 185
R986 VDD.n1576 VDD.n1456 185
R987 VDD.n1575 VDD.n1574 185
R988 VDD.n1572 VDD.n1457 185
R989 VDD.n1570 VDD.n1569 185
R990 VDD.n1568 VDD.n1458 185
R991 VDD.n1567 VDD.n1566 185
R992 VDD.n1564 VDD.n1459 185
R993 VDD.n1562 VDD.n1561 185
R994 VDD.n1560 VDD.n1460 185
R995 VDD.n1559 VDD.n1558 185
R996 VDD.n1556 VDD.n1461 185
R997 VDD.n1554 VDD.n1553 185
R998 VDD.n1552 VDD.n1462 185
R999 VDD.n1551 VDD.n1550 185
R1000 VDD.n1817 VDD.n1816 185
R1001 VDD.n1819 VDD.n1818 185
R1002 VDD.n1821 VDD.n1820 185
R1003 VDD.n1824 VDD.n1823 185
R1004 VDD.n1826 VDD.n1825 185
R1005 VDD.n1828 VDD.n1827 185
R1006 VDD.n1830 VDD.n1829 185
R1007 VDD.n1832 VDD.n1831 185
R1008 VDD.n1834 VDD.n1833 185
R1009 VDD.n1836 VDD.n1835 185
R1010 VDD.n1838 VDD.n1837 185
R1011 VDD.n1840 VDD.n1839 185
R1012 VDD.n1842 VDD.n1841 185
R1013 VDD.n1844 VDD.n1843 185
R1014 VDD.n1846 VDD.n1845 185
R1015 VDD.n1848 VDD.n1847 185
R1016 VDD.n1850 VDD.n1849 185
R1017 VDD.n1852 VDD.n1851 185
R1018 VDD.n1854 VDD.n1853 185
R1019 VDD.n1855 VDD.n499 185
R1020 VDD.n1857 VDD.n1856 185
R1021 VDD.n1858 VDD.n1857 185
R1022 VDD.n1815 VDD.n503 185
R1023 VDD.n1815 VDD.n476 185
R1024 VDD.n1814 VDD.n505 185
R1025 VDD.n1814 VDD.n1813 185
R1026 VDD.n1466 VDD.n504 185
R1027 VDD.n514 VDD.n504 185
R1028 VDD.n1467 VDD.n512 185
R1029 VDD.n1807 VDD.n512 185
R1030 VDD.n1469 VDD.n1468 185
R1031 VDD.n1468 VDD.n511 185
R1032 VDD.n1470 VDD.n524 185
R1033 VDD.t40 VDD.n524 185
R1034 VDD.n1472 VDD.n1471 185
R1035 VDD.n1471 VDD.n522 185
R1036 VDD.n1473 VDD.n529 185
R1037 VDD.n1744 VDD.n529 185
R1038 VDD.n1475 VDD.n1474 185
R1039 VDD.n1474 VDD.n528 185
R1040 VDD.n1476 VDD.n535 185
R1041 VDD.n1736 VDD.n535 185
R1042 VDD.n1478 VDD.n1477 185
R1043 VDD.n1477 VDD.n543 185
R1044 VDD.n1479 VDD.n541 185
R1045 VDD.n1730 VDD.n541 185
R1046 VDD.n1481 VDD.n1480 185
R1047 VDD.n1480 VDD.n540 185
R1048 VDD.n1482 VDD.n548 185
R1049 VDD.n1724 VDD.n548 185
R1050 VDD.n1484 VDD.n1483 185
R1051 VDD.n1483 VDD.n547 185
R1052 VDD.n1485 VDD.n554 185
R1053 VDD.n1718 VDD.n554 185
R1054 VDD.n1487 VDD.n1486 185
R1055 VDD.n1486 VDD.n553 185
R1056 VDD.n1488 VDD.n559 185
R1057 VDD.n1712 VDD.n559 185
R1058 VDD.n1490 VDD.n1489 185
R1059 VDD.n1489 VDD.n567 185
R1060 VDD.n1491 VDD.n565 185
R1061 VDD.n1706 VDD.n565 185
R1062 VDD.n1493 VDD.n1492 185
R1063 VDD.n1492 VDD.n564 185
R1064 VDD.n1494 VDD.n572 185
R1065 VDD.n1700 VDD.n572 185
R1066 VDD.n1496 VDD.n1495 185
R1067 VDD.n1495 VDD.n571 185
R1068 VDD.n1497 VDD.n578 185
R1069 VDD.n1694 VDD.n578 185
R1070 VDD.n1499 VDD.n1498 185
R1071 VDD.n1498 VDD.n577 185
R1072 VDD.n1500 VDD.n584 185
R1073 VDD.n1688 VDD.n584 185
R1074 VDD.n1502 VDD.n1501 185
R1075 VDD.n1501 VDD.n583 185
R1076 VDD.n1503 VDD.n590 185
R1077 VDD.n1682 VDD.n590 185
R1078 VDD.n1505 VDD.n1504 185
R1079 VDD.n1504 VDD.n589 185
R1080 VDD.n1506 VDD.n596 185
R1081 VDD.n1676 VDD.n596 185
R1082 VDD.n1508 VDD.n1507 185
R1083 VDD.n1507 VDD.n595 185
R1084 VDD.n1509 VDD.n602 185
R1085 VDD.n1670 VDD.n602 185
R1086 VDD.n1511 VDD.n1510 185
R1087 VDD.n1510 VDD.n601 185
R1088 VDD.n1512 VDD.n608 185
R1089 VDD.n1664 VDD.n608 185
R1090 VDD.n1514 VDD.n1513 185
R1091 VDD.n1513 VDD.n607 185
R1092 VDD.n1515 VDD.n614 185
R1093 VDD.n1658 VDD.n614 185
R1094 VDD.n1517 VDD.n1516 185
R1095 VDD.n1516 VDD.n613 185
R1096 VDD.n1518 VDD.n620 185
R1097 VDD.n1652 VDD.n620 185
R1098 VDD.n1520 VDD.n1519 185
R1099 VDD.n1519 VDD.n619 185
R1100 VDD.n1521 VDD.n626 185
R1101 VDD.n1646 VDD.n626 185
R1102 VDD.n1523 VDD.n1522 185
R1103 VDD.n1522 VDD.n625 185
R1104 VDD.n1524 VDD.n632 185
R1105 VDD.n1640 VDD.n632 185
R1106 VDD.n1526 VDD.n1525 185
R1107 VDD.n1525 VDD.n631 185
R1108 VDD.n1527 VDD.n638 185
R1109 VDD.n1634 VDD.n638 185
R1110 VDD.n1529 VDD.n1528 185
R1111 VDD.n1528 VDD.n637 185
R1112 VDD.n1530 VDD.n644 185
R1113 VDD.n1628 VDD.n644 185
R1114 VDD.n1532 VDD.n1531 185
R1115 VDD.n1531 VDD.n643 185
R1116 VDD.n1533 VDD.n650 185
R1117 VDD.n1622 VDD.n650 185
R1118 VDD.n1535 VDD.n1534 185
R1119 VDD.n1534 VDD.n649 185
R1120 VDD.n1536 VDD.n656 185
R1121 VDD.n1616 VDD.n656 185
R1122 VDD.n1538 VDD.n1537 185
R1123 VDD.n1537 VDD.n655 185
R1124 VDD.n1539 VDD.n661 185
R1125 VDD.n1610 VDD.n661 185
R1126 VDD.n1541 VDD.n1540 185
R1127 VDD.n1540 VDD.t50 185
R1128 VDD.n1542 VDD.n667 185
R1129 VDD.n1604 VDD.n667 185
R1130 VDD.n1544 VDD.n1543 185
R1131 VDD.n1543 VDD.n666 185
R1132 VDD.n1545 VDD.n673 185
R1133 VDD.n1598 VDD.n673 185
R1134 VDD.n1547 VDD.n1546 185
R1135 VDD.n1546 VDD.n672 185
R1136 VDD.n1548 VDD.n1320 185
R1137 VDD.n1592 VDD.n1320 185
R1138 VDD.n127 VDD.n126 185
R1139 VDD.n2711 VDD.n127 185
R1140 VDD.n2714 VDD.n2713 185
R1141 VDD.n2713 VDD.n2712 185
R1142 VDD.n2715 VDD.n121 185
R1143 VDD.n121 VDD.n120 185
R1144 VDD.n2717 VDD.n2716 185
R1145 VDD.n2718 VDD.n2717 185
R1146 VDD.n115 VDD.n114 185
R1147 VDD.n2719 VDD.n115 185
R1148 VDD.n2722 VDD.n2721 185
R1149 VDD.n2721 VDD.n2720 185
R1150 VDD.n2723 VDD.n109 185
R1151 VDD.n116 VDD.n109 185
R1152 VDD.n2725 VDD.n2724 185
R1153 VDD.n2726 VDD.n2725 185
R1154 VDD.n105 VDD.n104 185
R1155 VDD.n2727 VDD.n105 185
R1156 VDD.n2730 VDD.n2729 185
R1157 VDD.n2729 VDD.n2728 185
R1158 VDD.n2731 VDD.n99 185
R1159 VDD.n99 VDD.n98 185
R1160 VDD.n2733 VDD.n2732 185
R1161 VDD.n2734 VDD.n2733 185
R1162 VDD.n94 VDD.n93 185
R1163 VDD.n2735 VDD.n94 185
R1164 VDD.n2738 VDD.n2737 185
R1165 VDD.n2737 VDD.n2736 185
R1166 VDD.n2739 VDD.n88 185
R1167 VDD.n88 VDD.n87 185
R1168 VDD.n2741 VDD.n2740 185
R1169 VDD.n2742 VDD.n2741 185
R1170 VDD.n83 VDD.n82 185
R1171 VDD.n2743 VDD.n83 185
R1172 VDD.n2746 VDD.n2745 185
R1173 VDD.n2745 VDD.n2744 185
R1174 VDD.n2747 VDD.n77 185
R1175 VDD.n77 VDD.n76 185
R1176 VDD.n2749 VDD.n2748 185
R1177 VDD.n2750 VDD.n2749 185
R1178 VDD.n72 VDD.n71 185
R1179 VDD.n2751 VDD.n72 185
R1180 VDD.n2754 VDD.n2753 185
R1181 VDD.n2753 VDD.n2752 185
R1182 VDD.n2755 VDD.n66 185
R1183 VDD.n66 VDD.n65 185
R1184 VDD.n2757 VDD.n2756 185
R1185 VDD.n2758 VDD.n2757 185
R1186 VDD.n61 VDD.n60 185
R1187 VDD.n2759 VDD.n61 185
R1188 VDD.n2762 VDD.n2761 185
R1189 VDD.n2761 VDD.n2760 185
R1190 VDD.n2763 VDD.n55 185
R1191 VDD.n55 VDD.n54 185
R1192 VDD.n2765 VDD.n2764 185
R1193 VDD.n2766 VDD.n2765 185
R1194 VDD.n50 VDD.n49 185
R1195 VDD.n2767 VDD.n50 185
R1196 VDD.n2770 VDD.n2769 185
R1197 VDD.n2769 VDD.n2768 185
R1198 VDD.n2771 VDD.n45 185
R1199 VDD.n45 VDD.n44 185
R1200 VDD.n2773 VDD.n2772 185
R1201 VDD.n2774 VDD.n2773 185
R1202 VDD.n40 VDD.n38 185
R1203 VDD.n2775 VDD.n40 185
R1204 VDD.n2778 VDD.n2777 185
R1205 VDD.n2777 VDD.n2776 185
R1206 VDD.n39 VDD.n37 185
R1207 VDD.n2606 VDD.n39 185
R1208 VDD.n2604 VDD.n2603 185
R1209 VDD.n2605 VDD.n2604 185
R1210 VDD.n182 VDD.n181 185
R1211 VDD.n181 VDD.n180 185
R1212 VDD.n2599 VDD.n2598 185
R1213 VDD.n2598 VDD.n2597 185
R1214 VDD.n185 VDD.n184 185
R1215 VDD.n186 VDD.n185 185
R1216 VDD.n2585 VDD.n2584 185
R1217 VDD.n2586 VDD.n2585 185
R1218 VDD.n195 VDD.n194 185
R1219 VDD.n194 VDD.n193 185
R1220 VDD.n2580 VDD.n2579 185
R1221 VDD.n2579 VDD.n2578 185
R1222 VDD.n198 VDD.n197 185
R1223 VDD.n199 VDD.n198 185
R1224 VDD.n2569 VDD.n2568 185
R1225 VDD.n2570 VDD.n2569 185
R1226 VDD.n207 VDD.n206 185
R1227 VDD.n206 VDD.n205 185
R1228 VDD.n2564 VDD.n2563 185
R1229 VDD.n2563 VDD.n2562 185
R1230 VDD.n210 VDD.n209 185
R1231 VDD.n217 VDD.n210 185
R1232 VDD.n2553 VDD.n2552 185
R1233 VDD.n2554 VDD.n2553 185
R1234 VDD.n219 VDD.n218 185
R1235 VDD.n218 VDD.n216 185
R1236 VDD.n2548 VDD.n2547 185
R1237 VDD.n2547 VDD.n2546 185
R1238 VDD.n222 VDD.n221 185
R1239 VDD.n223 VDD.n222 185
R1240 VDD.n2537 VDD.n2536 185
R1241 VDD.n2538 VDD.n2537 185
R1242 VDD.n231 VDD.n230 185
R1243 VDD.n230 VDD.n229 185
R1244 VDD.n2532 VDD.n2531 185
R1245 VDD.n2531 VDD.n2530 185
R1246 VDD.n234 VDD.n233 185
R1247 VDD.n235 VDD.n234 185
R1248 VDD.n2521 VDD.n2520 185
R1249 VDD.n2522 VDD.n2521 185
R1250 VDD.n243 VDD.n242 185
R1251 VDD.n242 VDD.n241 185
R1252 VDD.n2516 VDD.n2515 185
R1253 VDD.n2515 VDD.n2514 185
R1254 VDD.n246 VDD.n245 185
R1255 VDD.n247 VDD.n246 185
R1256 VDD.n2505 VDD.n2504 185
R1257 VDD.n2506 VDD.n2505 185
R1258 VDD.n255 VDD.n254 185
R1259 VDD.n254 VDD.n253 185
R1260 VDD.n2500 VDD.n2499 185
R1261 VDD.n2499 VDD.n2498 185
R1262 VDD.n258 VDD.n257 185
R1263 VDD.n259 VDD.n258 185
R1264 VDD.n2489 VDD.n2488 185
R1265 VDD.n2490 VDD.n2489 185
R1266 VDD.n267 VDD.n266 185
R1267 VDD.n266 VDD.n265 185
R1268 VDD.n2484 VDD.n2483 185
R1269 VDD.n2483 VDD.n2482 185
R1270 VDD.n270 VDD.n269 185
R1271 VDD.n271 VDD.n270 185
R1272 VDD.n2473 VDD.n2472 185
R1273 VDD.n2474 VDD.n2473 185
R1274 VDD.n2469 VDD.n2402 185
R1275 VDD.n2468 VDD.n2467 185
R1276 VDD.n2465 VDD.n2404 185
R1277 VDD.n2465 VDD.n2401 185
R1278 VDD.n2464 VDD.n2463 185
R1279 VDD.n2462 VDD.n2461 185
R1280 VDD.n2460 VDD.n2409 185
R1281 VDD.n2458 VDD.n2457 185
R1282 VDD.n2456 VDD.n2410 185
R1283 VDD.n2454 VDD.n2453 185
R1284 VDD.n2451 VDD.n2417 185
R1285 VDD.n2449 VDD.n2448 185
R1286 VDD.n2447 VDD.n2418 185
R1287 VDD.n2446 VDD.n2445 185
R1288 VDD.n2443 VDD.n2423 185
R1289 VDD.n2441 VDD.n2440 185
R1290 VDD.n2439 VDD.n2424 185
R1291 VDD.n2438 VDD.n2429 185
R1292 VDD.n2435 VDD.n2432 185
R1293 VDD.n2430 VDD.n275 185
R1294 VDD.n157 VDD.n156 185
R1295 VDD.n2671 VDD.n2670 185
R1296 VDD.n2673 VDD.n2672 185
R1297 VDD.n2675 VDD.n2674 185
R1298 VDD.n2677 VDD.n2676 185
R1299 VDD.n2679 VDD.n2678 185
R1300 VDD.n2681 VDD.n2680 185
R1301 VDD.n2683 VDD.n2682 185
R1302 VDD.n2685 VDD.n2684 185
R1303 VDD.n2687 VDD.n2686 185
R1304 VDD.n2689 VDD.n2688 185
R1305 VDD.n2694 VDD.n2693 185
R1306 VDD.n2696 VDD.n2695 185
R1307 VDD.n2698 VDD.n2697 185
R1308 VDD.n2700 VDD.n2699 185
R1309 VDD.n2703 VDD.n2702 185
R1310 VDD.n2701 VDD.n142 185
R1311 VDD.n2707 VDD.n139 185
R1312 VDD.n2709 VDD.n2708 185
R1313 VDD.n2710 VDD.n2709 185
R1314 VDD.n2666 VDD.n129 185
R1315 VDD.n2711 VDD.n129 185
R1316 VDD.n2665 VDD.n128 185
R1317 VDD.n2712 VDD.n128 185
R1318 VDD.n2664 VDD.n2663 185
R1319 VDD.n2663 VDD.n120 185
R1320 VDD.n161 VDD.n119 185
R1321 VDD.n2718 VDD.n119 185
R1322 VDD.n2659 VDD.n118 185
R1323 VDD.n2719 VDD.n118 185
R1324 VDD.n2658 VDD.n117 185
R1325 VDD.n2720 VDD.n117 185
R1326 VDD.n2657 VDD.n2656 185
R1327 VDD.n2656 VDD.n116 185
R1328 VDD.n163 VDD.n108 185
R1329 VDD.n2726 VDD.n108 185
R1330 VDD.n2652 VDD.n107 185
R1331 VDD.n2727 VDD.n107 185
R1332 VDD.n2651 VDD.n106 185
R1333 VDD.n2728 VDD.n106 185
R1334 VDD.n2650 VDD.n2649 185
R1335 VDD.n2649 VDD.n98 185
R1336 VDD.n165 VDD.n97 185
R1337 VDD.n2734 VDD.n97 185
R1338 VDD.n2645 VDD.n96 185
R1339 VDD.n2735 VDD.n96 185
R1340 VDD.n2644 VDD.n95 185
R1341 VDD.n2736 VDD.n95 185
R1342 VDD.n2643 VDD.n2642 185
R1343 VDD.n2642 VDD.n87 185
R1344 VDD.n167 VDD.n86 185
R1345 VDD.n2742 VDD.n86 185
R1346 VDD.n2638 VDD.n85 185
R1347 VDD.n2743 VDD.n85 185
R1348 VDD.n2637 VDD.n84 185
R1349 VDD.n2744 VDD.n84 185
R1350 VDD.n2636 VDD.n2635 185
R1351 VDD.n2635 VDD.n76 185
R1352 VDD.n169 VDD.n75 185
R1353 VDD.n2750 VDD.n75 185
R1354 VDD.n2631 VDD.n74 185
R1355 VDD.n2751 VDD.n74 185
R1356 VDD.n2630 VDD.n73 185
R1357 VDD.n2752 VDD.n73 185
R1358 VDD.n2629 VDD.n2628 185
R1359 VDD.n2628 VDD.n65 185
R1360 VDD.n171 VDD.n64 185
R1361 VDD.n2758 VDD.n64 185
R1362 VDD.n2624 VDD.n63 185
R1363 VDD.n2759 VDD.n63 185
R1364 VDD.n2623 VDD.n62 185
R1365 VDD.n2760 VDD.n62 185
R1366 VDD.n2622 VDD.n2621 185
R1367 VDD.n2621 VDD.n54 185
R1368 VDD.n173 VDD.n53 185
R1369 VDD.n2766 VDD.n53 185
R1370 VDD.n2617 VDD.n52 185
R1371 VDD.n2767 VDD.n52 185
R1372 VDD.n2616 VDD.n51 185
R1373 VDD.n2768 VDD.n51 185
R1374 VDD.n2615 VDD.n2614 185
R1375 VDD.n2614 VDD.n44 185
R1376 VDD.n175 VDD.n43 185
R1377 VDD.n2774 VDD.n43 185
R1378 VDD.n2610 VDD.n42 185
R1379 VDD.n2775 VDD.n42 185
R1380 VDD.n2609 VDD.n41 185
R1381 VDD.n2776 VDD.n41 185
R1382 VDD.n2608 VDD.n2607 185
R1383 VDD.n2607 VDD.n2606 185
R1384 VDD.n179 VDD.n177 185
R1385 VDD.n2605 VDD.n179 185
R1386 VDD.n2594 VDD.n188 185
R1387 VDD.n188 VDD.n180 185
R1388 VDD.n2596 VDD.n2595 185
R1389 VDD.n2597 VDD.n2596 185
R1390 VDD.n189 VDD.n187 185
R1391 VDD.n187 VDD.n186 185
R1392 VDD.n2588 VDD.n2587 185
R1393 VDD.n2587 VDD.n2586 185
R1394 VDD.n192 VDD.n191 185
R1395 VDD.n193 VDD.n192 185
R1396 VDD.n2577 VDD.n2576 185
R1397 VDD.n2578 VDD.n2577 185
R1398 VDD.n201 VDD.n200 185
R1399 VDD.n200 VDD.n199 185
R1400 VDD.n2572 VDD.n2571 185
R1401 VDD.n2571 VDD.n2570 185
R1402 VDD.n204 VDD.n203 185
R1403 VDD.n205 VDD.n204 185
R1404 VDD.n2561 VDD.n2560 185
R1405 VDD.n2562 VDD.n2561 185
R1406 VDD.n212 VDD.n211 185
R1407 VDD.n217 VDD.n211 185
R1408 VDD.n2556 VDD.n2555 185
R1409 VDD.n2555 VDD.n2554 185
R1410 VDD.n215 VDD.n214 185
R1411 VDD.n216 VDD.n215 185
R1412 VDD.n2545 VDD.n2544 185
R1413 VDD.n2546 VDD.n2545 185
R1414 VDD.n225 VDD.n224 185
R1415 VDD.n224 VDD.n223 185
R1416 VDD.n2540 VDD.n2539 185
R1417 VDD.n2539 VDD.n2538 185
R1418 VDD.n228 VDD.n227 185
R1419 VDD.n229 VDD.n228 185
R1420 VDD.n2529 VDD.n2528 185
R1421 VDD.n2530 VDD.n2529 185
R1422 VDD.n237 VDD.n236 185
R1423 VDD.n236 VDD.n235 185
R1424 VDD.n2524 VDD.n2523 185
R1425 VDD.n2523 VDD.n2522 185
R1426 VDD.n240 VDD.n239 185
R1427 VDD.n241 VDD.n240 185
R1428 VDD.n2513 VDD.n2512 185
R1429 VDD.n2514 VDD.n2513 185
R1430 VDD.n249 VDD.n248 185
R1431 VDD.n248 VDD.n247 185
R1432 VDD.n2508 VDD.n2507 185
R1433 VDD.n2507 VDD.n2506 185
R1434 VDD.n252 VDD.n251 185
R1435 VDD.n253 VDD.n252 185
R1436 VDD.n2497 VDD.n2496 185
R1437 VDD.n2498 VDD.n2497 185
R1438 VDD.n261 VDD.n260 185
R1439 VDD.n260 VDD.n259 185
R1440 VDD.n2492 VDD.n2491 185
R1441 VDD.n2491 VDD.n2490 185
R1442 VDD.n264 VDD.n263 185
R1443 VDD.n265 VDD.n264 185
R1444 VDD.n2481 VDD.n2480 185
R1445 VDD.n2482 VDD.n2481 185
R1446 VDD.n273 VDD.n272 185
R1447 VDD.n272 VDD.n271 185
R1448 VDD.n2476 VDD.n2475 185
R1449 VDD.n2475 VDD.n2474 185
R1450 VDD.n2131 VDD.n1863 185
R1451 VDD.n2130 VDD.n2129 185
R1452 VDD.n2127 VDD.n1864 185
R1453 VDD.n2127 VDD.n1859 185
R1454 VDD.n2126 VDD.n2125 185
R1455 VDD.n2124 VDD.n2123 185
R1456 VDD.n2122 VDD.n1866 185
R1457 VDD.n2120 VDD.n2119 185
R1458 VDD.n2118 VDD.n1867 185
R1459 VDD.n2117 VDD.n2116 185
R1460 VDD.n2114 VDD.n1868 185
R1461 VDD.n2112 VDD.n2111 185
R1462 VDD.n2110 VDD.n1869 185
R1463 VDD.n2109 VDD.n2108 185
R1464 VDD.n2106 VDD.n1870 185
R1465 VDD.n2104 VDD.n2103 185
R1466 VDD.n2102 VDD.n1871 185
R1467 VDD.n2101 VDD.n2100 185
R1468 VDD.n2098 VDD.n1872 185
R1469 VDD.n2096 VDD.n2095 185
R1470 VDD.n2094 VDD.n1873 185
R1471 VDD.n2093 VDD.n2092 185
R1472 VDD.n2359 VDD.n2358 185
R1473 VDD.n2361 VDD.n2360 185
R1474 VDD.n2363 VDD.n2362 185
R1475 VDD.n2366 VDD.n2365 185
R1476 VDD.n2368 VDD.n2367 185
R1477 VDD.n2370 VDD.n2369 185
R1478 VDD.n2372 VDD.n2371 185
R1479 VDD.n2374 VDD.n2373 185
R1480 VDD.n2376 VDD.n2375 185
R1481 VDD.n2378 VDD.n2377 185
R1482 VDD.n2380 VDD.n2379 185
R1483 VDD.n2382 VDD.n2381 185
R1484 VDD.n2384 VDD.n2383 185
R1485 VDD.n2386 VDD.n2385 185
R1486 VDD.n2388 VDD.n2387 185
R1487 VDD.n2390 VDD.n2389 185
R1488 VDD.n2392 VDD.n2391 185
R1489 VDD.n2394 VDD.n2393 185
R1490 VDD.n2396 VDD.n2395 185
R1491 VDD.n2397 VDD.n299 185
R1492 VDD.n2399 VDD.n2398 185
R1493 VDD.n2400 VDD.n2399 185
R1494 VDD.n2357 VDD.n303 185
R1495 VDD.n2357 VDD.n276 185
R1496 VDD.n2356 VDD.n305 185
R1497 VDD.n2356 VDD.n2355 185
R1498 VDD.n1877 VDD.n304 185
R1499 VDD.n306 VDD.n304 185
R1500 VDD.n1878 VDD.n313 185
R1501 VDD.n2349 VDD.n313 185
R1502 VDD.n1880 VDD.n1879 185
R1503 VDD.n1879 VDD.n312 185
R1504 VDD.n1881 VDD.n324 185
R1505 VDD.t24 VDD.n324 185
R1506 VDD.n1883 VDD.n1882 185
R1507 VDD.n1882 VDD.n322 185
R1508 VDD.n1884 VDD.n329 185
R1509 VDD.n2286 VDD.n329 185
R1510 VDD.n1886 VDD.n1885 185
R1511 VDD.n1885 VDD.n328 185
R1512 VDD.n1887 VDD.n336 185
R1513 VDD.n2278 VDD.n336 185
R1514 VDD.n1889 VDD.n1888 185
R1515 VDD.n1888 VDD.n335 185
R1516 VDD.n1890 VDD.n342 185
R1517 VDD.n2272 VDD.n342 185
R1518 VDD.n1892 VDD.n1891 185
R1519 VDD.n1891 VDD.n341 185
R1520 VDD.n1893 VDD.n348 185
R1521 VDD.n2266 VDD.n348 185
R1522 VDD.n1895 VDD.n1894 185
R1523 VDD.n1894 VDD.n347 185
R1524 VDD.n1896 VDD.n354 185
R1525 VDD.n2260 VDD.n354 185
R1526 VDD.n1898 VDD.n1897 185
R1527 VDD.n1897 VDD.n353 185
R1528 VDD.n1899 VDD.n360 185
R1529 VDD.n2254 VDD.n360 185
R1530 VDD.n1901 VDD.n1900 185
R1531 VDD.n1900 VDD.n359 185
R1532 VDD.n1902 VDD.n366 185
R1533 VDD.n2248 VDD.n366 185
R1534 VDD.n1904 VDD.n1903 185
R1535 VDD.n1903 VDD.n365 185
R1536 VDD.n1905 VDD.n372 185
R1537 VDD.n2242 VDD.n372 185
R1538 VDD.n1907 VDD.n1906 185
R1539 VDD.n1906 VDD.n371 185
R1540 VDD.n1908 VDD.n378 185
R1541 VDD.n2236 VDD.n378 185
R1542 VDD.n1910 VDD.n1909 185
R1543 VDD.n1909 VDD.n377 185
R1544 VDD.n1911 VDD.n384 185
R1545 VDD.n2230 VDD.n384 185
R1546 VDD.n1913 VDD.n1912 185
R1547 VDD.n1912 VDD.n383 185
R1548 VDD.n1914 VDD.n390 185
R1549 VDD.n2224 VDD.n390 185
R1550 VDD.n1916 VDD.n1915 185
R1551 VDD.n1915 VDD.n389 185
R1552 VDD.n1917 VDD.n396 185
R1553 VDD.n2218 VDD.n396 185
R1554 VDD.n1919 VDD.n1918 185
R1555 VDD.n1918 VDD.n395 185
R1556 VDD.n1920 VDD.n402 185
R1557 VDD.n2212 VDD.n402 185
R1558 VDD.n1922 VDD.n1921 185
R1559 VDD.n1921 VDD.n401 185
R1560 VDD.n1923 VDD.n408 185
R1561 VDD.n2206 VDD.n408 185
R1562 VDD.n1925 VDD.n1924 185
R1563 VDD.n1924 VDD.n407 185
R1564 VDD.n1926 VDD.n414 185
R1565 VDD.n2200 VDD.n414 185
R1566 VDD.n1928 VDD.n1927 185
R1567 VDD.n1927 VDD.n413 185
R1568 VDD.n1929 VDD.n420 185
R1569 VDD.n2194 VDD.n420 185
R1570 VDD.n1931 VDD.n1930 185
R1571 VDD.n1930 VDD.n419 185
R1572 VDD.n1932 VDD.n425 185
R1573 VDD.n2188 VDD.n425 185
R1574 VDD.n2065 VDD.n2064 185
R1575 VDD.n2064 VDD.n2063 185
R1576 VDD.n2066 VDD.n431 185
R1577 VDD.n2182 VDD.n431 185
R1578 VDD.n2068 VDD.n2067 185
R1579 VDD.n2067 VDD.n430 185
R1580 VDD.n2069 VDD.n437 185
R1581 VDD.n2176 VDD.n437 185
R1582 VDD.n2071 VDD.n2070 185
R1583 VDD.n2070 VDD.n436 185
R1584 VDD.n2072 VDD.n443 185
R1585 VDD.n2170 VDD.n443 185
R1586 VDD.n2074 VDD.n2073 185
R1587 VDD.n2073 VDD.n442 185
R1588 VDD.n2075 VDD.n448 185
R1589 VDD.n2164 VDD.n448 185
R1590 VDD.n2077 VDD.n2076 185
R1591 VDD.n2076 VDD.n456 185
R1592 VDD.n2078 VDD.n454 185
R1593 VDD.n2158 VDD.n454 185
R1594 VDD.n2080 VDD.n2079 185
R1595 VDD.n2079 VDD.n453 185
R1596 VDD.n2081 VDD.n460 185
R1597 VDD.n2152 VDD.n460 185
R1598 VDD.n2083 VDD.n2082 185
R1599 VDD.n2082 VDD.t16 185
R1600 VDD.n2084 VDD.n466 185
R1601 VDD.n2146 VDD.n466 185
R1602 VDD.n2086 VDD.n2085 185
R1603 VDD.n2085 VDD.n465 185
R1604 VDD.n2087 VDD.n471 185
R1605 VDD.n2140 VDD.n471 185
R1606 VDD.n2089 VDD.n2088 185
R1607 VDD.n2088 VDD.n1862 185
R1608 VDD.n2090 VDD.n1860 185
R1609 VDD.n2134 VDD.n1860 185
R1610 VDD.n2133 VDD.n2132 185
R1611 VDD.n2134 VDD.n2133 185
R1612 VDD.n470 VDD.n469 185
R1613 VDD.n1862 VDD.n470 185
R1614 VDD.n2142 VDD.n2141 185
R1615 VDD.n2141 VDD.n2140 185
R1616 VDD.n2143 VDD.n468 185
R1617 VDD.n468 VDD.n465 185
R1618 VDD.n2145 VDD.n2144 185
R1619 VDD.n2146 VDD.n2145 185
R1620 VDD.n459 VDD.n458 185
R1621 VDD.t16 VDD.n459 185
R1622 VDD.n2154 VDD.n2153 185
R1623 VDD.n2153 VDD.n2152 185
R1624 VDD.n2155 VDD.n457 185
R1625 VDD.n457 VDD.n453 185
R1626 VDD.n2157 VDD.n2156 185
R1627 VDD.n2158 VDD.n2157 185
R1628 VDD.n447 VDD.n446 185
R1629 VDD.n456 VDD.n447 185
R1630 VDD.n2166 VDD.n2165 185
R1631 VDD.n2165 VDD.n2164 185
R1632 VDD.n2167 VDD.n445 185
R1633 VDD.n445 VDD.n442 185
R1634 VDD.n2169 VDD.n2168 185
R1635 VDD.n2170 VDD.n2169 185
R1636 VDD.n435 VDD.n434 185
R1637 VDD.n436 VDD.n435 185
R1638 VDD.n2178 VDD.n2177 185
R1639 VDD.n2177 VDD.n2176 185
R1640 VDD.n2179 VDD.n433 185
R1641 VDD.n433 VDD.n430 185
R1642 VDD.n2181 VDD.n2180 185
R1643 VDD.n2182 VDD.n2181 185
R1644 VDD.n424 VDD.n423 185
R1645 VDD.n2063 VDD.n424 185
R1646 VDD.n2190 VDD.n2189 185
R1647 VDD.n2189 VDD.n2188 185
R1648 VDD.n2191 VDD.n422 185
R1649 VDD.n422 VDD.n419 185
R1650 VDD.n2193 VDD.n2192 185
R1651 VDD.n2194 VDD.n2193 185
R1652 VDD.n412 VDD.n411 185
R1653 VDD.n413 VDD.n412 185
R1654 VDD.n2202 VDD.n2201 185
R1655 VDD.n2201 VDD.n2200 185
R1656 VDD.n2203 VDD.n410 185
R1657 VDD.n410 VDD.n407 185
R1658 VDD.n2205 VDD.n2204 185
R1659 VDD.n2206 VDD.n2205 185
R1660 VDD.n400 VDD.n399 185
R1661 VDD.n401 VDD.n400 185
R1662 VDD.n2214 VDD.n2213 185
R1663 VDD.n2213 VDD.n2212 185
R1664 VDD.n2215 VDD.n398 185
R1665 VDD.n398 VDD.n395 185
R1666 VDD.n2217 VDD.n2216 185
R1667 VDD.n2218 VDD.n2217 185
R1668 VDD.n388 VDD.n387 185
R1669 VDD.n389 VDD.n388 185
R1670 VDD.n2226 VDD.n2225 185
R1671 VDD.n2225 VDD.n2224 185
R1672 VDD.n2227 VDD.n386 185
R1673 VDD.n386 VDD.n383 185
R1674 VDD.n2229 VDD.n2228 185
R1675 VDD.n2230 VDD.n2229 185
R1676 VDD.n376 VDD.n375 185
R1677 VDD.n377 VDD.n376 185
R1678 VDD.n2238 VDD.n2237 185
R1679 VDD.n2237 VDD.n2236 185
R1680 VDD.n2239 VDD.n374 185
R1681 VDD.n374 VDD.n371 185
R1682 VDD.n2241 VDD.n2240 185
R1683 VDD.n2242 VDD.n2241 185
R1684 VDD.n364 VDD.n363 185
R1685 VDD.n365 VDD.n364 185
R1686 VDD.n2250 VDD.n2249 185
R1687 VDD.n2249 VDD.n2248 185
R1688 VDD.n2251 VDD.n362 185
R1689 VDD.n362 VDD.n359 185
R1690 VDD.n2253 VDD.n2252 185
R1691 VDD.n2254 VDD.n2253 185
R1692 VDD.n352 VDD.n351 185
R1693 VDD.n353 VDD.n352 185
R1694 VDD.n2262 VDD.n2261 185
R1695 VDD.n2261 VDD.n2260 185
R1696 VDD.n2263 VDD.n350 185
R1697 VDD.n350 VDD.n347 185
R1698 VDD.n2265 VDD.n2264 185
R1699 VDD.n2266 VDD.n2265 185
R1700 VDD.n340 VDD.n339 185
R1701 VDD.n341 VDD.n340 185
R1702 VDD.n2274 VDD.n2273 185
R1703 VDD.n2273 VDD.n2272 185
R1704 VDD.n2275 VDD.n338 185
R1705 VDD.n338 VDD.n335 185
R1706 VDD.n2277 VDD.n2276 185
R1707 VDD.n2278 VDD.n2277 185
R1708 VDD.n327 VDD.n326 185
R1709 VDD.n328 VDD.n327 185
R1710 VDD.n2288 VDD.n2287 185
R1711 VDD.n2287 VDD.n2286 185
R1712 VDD.n2289 VDD.n325 185
R1713 VDD.n325 VDD.n322 185
R1714 VDD.n2291 VDD.n2290 185
R1715 VDD.t24 VDD.n2291 185
R1716 VDD.n311 VDD.n310 185
R1717 VDD.n312 VDD.n311 185
R1718 VDD.n2351 VDD.n2350 185
R1719 VDD.n2350 VDD.n2349 185
R1720 VDD.n2352 VDD.n309 185
R1721 VDD.n309 VDD.n306 185
R1722 VDD.n2354 VDD.n2353 185
R1723 VDD.n2355 VDD.n2354 185
R1724 VDD.n300 VDD.n298 185
R1725 VDD.n298 VDD.n276 185
R1726 VDD.n1317 VDD.n1316 185
R1727 VDD.n1318 VDD.n1317 185
R1728 VDD.n692 VDD.n688 185
R1729 VDD.n1280 VDD.n1279 185
R1730 VDD.n1278 VDD.n1277 185
R1731 VDD.n1284 VDD.n1276 185
R1732 VDD.n1285 VDD.n1275 185
R1733 VDD.n1286 VDD.n1274 185
R1734 VDD.n1273 VDD.n1271 185
R1735 VDD.n1290 VDD.n1270 185
R1736 VDD.n1291 VDD.n1269 185
R1737 VDD.n1292 VDD.n1268 185
R1738 VDD.n1267 VDD.n1262 185
R1739 VDD.n1296 VDD.n1261 185
R1740 VDD.n1297 VDD.n1260 185
R1741 VDD.n1298 VDD.n1259 185
R1742 VDD.n1258 VDD.n1256 185
R1743 VDD.n1302 VDD.n1255 185
R1744 VDD.n1303 VDD.n1254 185
R1745 VDD.n1304 VDD.n1253 185
R1746 VDD.n1313 VDD.n689 185
R1747 VDD.n689 VDD.n678 185
R1748 VDD.n1312 VDD.n1311 185
R1749 VDD.n1311 VDD.n1310 185
R1750 VDD.n696 VDD.n695 185
R1751 VDD.n697 VDD.n696 185
R1752 VDD.n1246 VDD.n1245 185
R1753 VDD.n1247 VDD.n1246 185
R1754 VDD.n707 VDD.n706 185
R1755 VDD.n706 VDD.n705 185
R1756 VDD.n1240 VDD.n1239 185
R1757 VDD.n1239 VDD.n1238 185
R1758 VDD.n710 VDD.n709 185
R1759 VDD.n711 VDD.n710 185
R1760 VDD.n1229 VDD.n1228 185
R1761 VDD.n1230 VDD.n1229 185
R1762 VDD.n719 VDD.n718 185
R1763 VDD.n718 VDD.n717 185
R1764 VDD.n1224 VDD.n1223 185
R1765 VDD.n1223 VDD.n1222 185
R1766 VDD.n722 VDD.n721 185
R1767 VDD.n723 VDD.n722 185
R1768 VDD.n1213 VDD.n1212 185
R1769 VDD.n1214 VDD.n1213 185
R1770 VDD.n731 VDD.n730 185
R1771 VDD.n730 VDD.n729 185
R1772 VDD.n1208 VDD.n1207 185
R1773 VDD.n1207 VDD.n1206 185
R1774 VDD.n734 VDD.n733 185
R1775 VDD.n735 VDD.n734 185
R1776 VDD.n1197 VDD.n1196 185
R1777 VDD.n1198 VDD.n1197 185
R1778 VDD.n743 VDD.n742 185
R1779 VDD.n742 VDD.n741 185
R1780 VDD.n1192 VDD.n1191 185
R1781 VDD.n1191 VDD.n1190 185
R1782 VDD.n746 VDD.n745 185
R1783 VDD.n747 VDD.n746 185
R1784 VDD.n1181 VDD.n1180 185
R1785 VDD.n1182 VDD.n1181 185
R1786 VDD.n755 VDD.n754 185
R1787 VDD.n754 VDD.n753 185
R1788 VDD.n1176 VDD.n1175 185
R1789 VDD.n1175 VDD.n1174 185
R1790 VDD.n758 VDD.n757 185
R1791 VDD.n1165 VDD.n758 185
R1792 VDD.n1164 VDD.n1163 185
R1793 VDD.n1166 VDD.n1164 185
R1794 VDD.n766 VDD.n765 185
R1795 VDD.n765 VDD.n764 185
R1796 VDD.n1159 VDD.n1158 185
R1797 VDD.n1158 VDD.n1157 185
R1798 VDD.n769 VDD.n768 185
R1799 VDD.n770 VDD.n769 185
R1800 VDD.n1148 VDD.n1147 185
R1801 VDD.n1149 VDD.n1148 185
R1802 VDD.n778 VDD.n777 185
R1803 VDD.n777 VDD.n776 185
R1804 VDD.n1143 VDD.n1142 185
R1805 VDD.n1142 VDD.n1141 185
R1806 VDD.n781 VDD.n780 185
R1807 VDD.n782 VDD.n781 185
R1808 VDD.n1132 VDD.n1131 185
R1809 VDD.n1133 VDD.n1132 185
R1810 VDD.n790 VDD.n789 185
R1811 VDD.n789 VDD.n788 185
R1812 VDD.n1127 VDD.n1126 185
R1813 VDD.n1126 VDD.n1125 185
R1814 VDD.n793 VDD.n792 185
R1815 VDD.n1095 VDD.n793 185
R1816 VDD.n1094 VDD.n1093 185
R1817 VDD.n1096 VDD.n1094 185
R1818 VDD.n801 VDD.n800 185
R1819 VDD.n800 VDD.n799 185
R1820 VDD.n1089 VDD.n1088 185
R1821 VDD.n1088 VDD.n1087 185
R1822 VDD.n804 VDD.n803 185
R1823 VDD.n805 VDD.n804 185
R1824 VDD.n1078 VDD.n1077 185
R1825 VDD.n1079 VDD.n1078 185
R1826 VDD.n813 VDD.n812 185
R1827 VDD.n812 VDD.n811 185
R1828 VDD.n1073 VDD.n1072 185
R1829 VDD.n1072 VDD.n1071 185
R1830 VDD.n816 VDD.n815 185
R1831 VDD.n817 VDD.n816 185
R1832 VDD.n1062 VDD.n1061 185
R1833 VDD.n1063 VDD.n1062 185
R1834 VDD.n825 VDD.n824 185
R1835 VDD.n824 VDD.n823 185
R1836 VDD.n1057 VDD.n1056 185
R1837 VDD.n1056 VDD.n1055 185
R1838 VDD.n828 VDD.n827 185
R1839 VDD.n1046 VDD.n828 185
R1840 VDD.n1045 VDD.n1044 185
R1841 VDD.n1047 VDD.n1045 185
R1842 VDD.n836 VDD.n835 185
R1843 VDD.n835 VDD.n834 185
R1844 VDD.n1040 VDD.n1039 185
R1845 VDD.n1039 VDD.n1038 185
R1846 VDD.n839 VDD.n838 185
R1847 VDD.n840 VDD.n839 185
R1848 VDD.n1029 VDD.n1028 185
R1849 VDD.n1030 VDD.n1029 185
R1850 VDD.n848 VDD.n847 185
R1851 VDD.n847 VDD.n846 185
R1852 VDD.n1024 VDD.n1023 185
R1853 VDD.n1023 VDD.n1022 185
R1854 VDD.n851 VDD.n850 185
R1855 VDD.n852 VDD.n851 185
R1856 VDD.n1013 VDD.n1012 185
R1857 VDD.n1014 VDD.n1013 185
R1858 VDD.n860 VDD.n859 185
R1859 VDD.n859 VDD.n858 185
R1860 VDD.n1008 VDD.n1007 185
R1861 VDD.n1007 VDD.n1006 185
R1862 VDD.n863 VDD.n862 185
R1863 VDD.n864 VDD.n863 185
R1864 VDD.n997 VDD.n996 185
R1865 VDD.n998 VDD.n997 185
R1866 VDD.n872 VDD.n871 185
R1867 VDD.n871 VDD.n870 185
R1868 VDD.n992 VDD.n991 185
R1869 VDD.n991 VDD.n990 185
R1870 VDD.n875 VDD.n874 185
R1871 VDD.n876 VDD.n875 185
R1872 VDD.n981 VDD.n980 185
R1873 VDD.n982 VDD.n981 185
R1874 VDD.n884 VDD.n883 185
R1875 VDD.n883 VDD.n882 185
R1876 VDD.n976 VDD.n975 185
R1877 VDD.n975 VDD.n974 185
R1878 VDD.n887 VDD.n886 185
R1879 VDD.n888 VDD.n887 185
R1880 VDD.n965 VDD.n964 185
R1881 VDD.n966 VDD.n965 185
R1882 VDD.n920 VDD.n892 185
R1883 VDD.n923 VDD.n922 185
R1884 VDD.n919 VDD.n918 185
R1885 VDD.n918 VDD.n893 185
R1886 VDD.n928 VDD.n927 185
R1887 VDD.n930 VDD.n917 185
R1888 VDD.n933 VDD.n932 185
R1889 VDD.n912 VDD.n911 185
R1890 VDD.n938 VDD.n937 185
R1891 VDD.n940 VDD.n910 185
R1892 VDD.n943 VDD.n942 185
R1893 VDD.n908 VDD.n907 185
R1894 VDD.n949 VDD.n948 185
R1895 VDD.n951 VDD.n906 185
R1896 VDD.n952 VDD.n903 185
R1897 VDD.n955 VDD.n954 185
R1898 VDD.n905 VDD.n900 185
R1899 VDD.n959 VDD.n901 185
R1900 VDD.n960 VDD.n897 185
R1901 VDD.n961 VDD.n894 185
R1902 VDD.n701 VDD.n699 185
R1903 VDD.n699 VDD.n678 185
R1904 VDD.n1309 VDD.n1308 185
R1905 VDD.n1310 VDD.n1309 185
R1906 VDD.n700 VDD.n698 185
R1907 VDD.n698 VDD.n697 185
R1908 VDD.n1249 VDD.n1248 185
R1909 VDD.n1248 VDD.n1247 185
R1910 VDD.n704 VDD.n703 185
R1911 VDD.n705 VDD.n704 185
R1912 VDD.n1237 VDD.n1236 185
R1913 VDD.n1238 VDD.n1237 185
R1914 VDD.n713 VDD.n712 185
R1915 VDD.n712 VDD.n711 185
R1916 VDD.n1232 VDD.n1231 185
R1917 VDD.n1231 VDD.n1230 185
R1918 VDD.n716 VDD.n715 185
R1919 VDD.n717 VDD.n716 185
R1920 VDD.n1221 VDD.n1220 185
R1921 VDD.n1222 VDD.n1221 185
R1922 VDD.n725 VDD.n724 185
R1923 VDD.n724 VDD.n723 185
R1924 VDD.n1216 VDD.n1215 185
R1925 VDD.n1215 VDD.n1214 185
R1926 VDD.n728 VDD.n727 185
R1927 VDD.n729 VDD.n728 185
R1928 VDD.n1205 VDD.n1204 185
R1929 VDD.n1206 VDD.n1205 185
R1930 VDD.n737 VDD.n736 185
R1931 VDD.n736 VDD.n735 185
R1932 VDD.n1200 VDD.n1199 185
R1933 VDD.n1199 VDD.n1198 185
R1934 VDD.n740 VDD.n739 185
R1935 VDD.n741 VDD.n740 185
R1936 VDD.n1189 VDD.n1188 185
R1937 VDD.n1190 VDD.n1189 185
R1938 VDD.n749 VDD.n748 185
R1939 VDD.n748 VDD.n747 185
R1940 VDD.n1184 VDD.n1183 185
R1941 VDD.n1183 VDD.n1182 185
R1942 VDD.n752 VDD.n751 185
R1943 VDD.n753 VDD.n752 185
R1944 VDD.n1173 VDD.n1172 185
R1945 VDD.n1174 VDD.n1173 185
R1946 VDD.n760 VDD.n759 185
R1947 VDD.n1165 VDD.n759 185
R1948 VDD.n1168 VDD.n1167 185
R1949 VDD.n1167 VDD.n1166 185
R1950 VDD.n763 VDD.n762 185
R1951 VDD.n764 VDD.n763 185
R1952 VDD.n1156 VDD.n1155 185
R1953 VDD.n1157 VDD.n1156 185
R1954 VDD.n772 VDD.n771 185
R1955 VDD.n771 VDD.n770 185
R1956 VDD.n1151 VDD.n1150 185
R1957 VDD.n1150 VDD.n1149 185
R1958 VDD.n775 VDD.n774 185
R1959 VDD.n776 VDD.n775 185
R1960 VDD.n1140 VDD.n1139 185
R1961 VDD.n1141 VDD.n1140 185
R1962 VDD.n784 VDD.n783 185
R1963 VDD.n783 VDD.n782 185
R1964 VDD.n1135 VDD.n1134 185
R1965 VDD.n1134 VDD.n1133 185
R1966 VDD.n787 VDD.n786 185
R1967 VDD.n788 VDD.n787 185
R1968 VDD.n1124 VDD.n1123 185
R1969 VDD.n1125 VDD.n1124 185
R1970 VDD.n795 VDD.n794 185
R1971 VDD.n1095 VDD.n794 185
R1972 VDD.n1098 VDD.n1097 185
R1973 VDD.n1097 VDD.n1096 185
R1974 VDD.n798 VDD.n797 185
R1975 VDD.n799 VDD.n798 185
R1976 VDD.n1086 VDD.n1085 185
R1977 VDD.n1087 VDD.n1086 185
R1978 VDD.n807 VDD.n806 185
R1979 VDD.n806 VDD.n805 185
R1980 VDD.n1081 VDD.n1080 185
R1981 VDD.n1080 VDD.n1079 185
R1982 VDD.n810 VDD.n809 185
R1983 VDD.n811 VDD.n810 185
R1984 VDD.n1070 VDD.n1069 185
R1985 VDD.n1071 VDD.n1070 185
R1986 VDD.n819 VDD.n818 185
R1987 VDD.n818 VDD.n817 185
R1988 VDD.n1065 VDD.n1064 185
R1989 VDD.n1064 VDD.n1063 185
R1990 VDD.n822 VDD.n821 185
R1991 VDD.n823 VDD.n822 185
R1992 VDD.n1054 VDD.n1053 185
R1993 VDD.n1055 VDD.n1054 185
R1994 VDD.n830 VDD.n829 185
R1995 VDD.n1046 VDD.n829 185
R1996 VDD.n1049 VDD.n1048 185
R1997 VDD.n1048 VDD.n1047 185
R1998 VDD.n833 VDD.n832 185
R1999 VDD.n834 VDD.n833 185
R2000 VDD.n1037 VDD.n1036 185
R2001 VDD.n1038 VDD.n1037 185
R2002 VDD.n842 VDD.n841 185
R2003 VDD.n841 VDD.n840 185
R2004 VDD.n1032 VDD.n1031 185
R2005 VDD.n1031 VDD.n1030 185
R2006 VDD.n845 VDD.n844 185
R2007 VDD.n846 VDD.n845 185
R2008 VDD.n1021 VDD.n1020 185
R2009 VDD.n1022 VDD.n1021 185
R2010 VDD.n854 VDD.n853 185
R2011 VDD.n853 VDD.n852 185
R2012 VDD.n1016 VDD.n1015 185
R2013 VDD.n1015 VDD.n1014 185
R2014 VDD.n857 VDD.n856 185
R2015 VDD.n858 VDD.n857 185
R2016 VDD.n1005 VDD.n1004 185
R2017 VDD.n1006 VDD.n1005 185
R2018 VDD.n866 VDD.n865 185
R2019 VDD.n865 VDD.n864 185
R2020 VDD.n1000 VDD.n999 185
R2021 VDD.n999 VDD.n998 185
R2022 VDD.n869 VDD.n868 185
R2023 VDD.n870 VDD.n869 185
R2024 VDD.n989 VDD.n988 185
R2025 VDD.n990 VDD.n989 185
R2026 VDD.n878 VDD.n877 185
R2027 VDD.n877 VDD.n876 185
R2028 VDD.n984 VDD.n983 185
R2029 VDD.n983 VDD.n982 185
R2030 VDD.n881 VDD.n880 185
R2031 VDD.n882 VDD.n881 185
R2032 VDD.n973 VDD.n972 185
R2033 VDD.n974 VDD.n973 185
R2034 VDD.n890 VDD.n889 185
R2035 VDD.n889 VDD.n888 185
R2036 VDD.n968 VDD.n967 185
R2037 VDD.n967 VDD.n966 185
R2038 VDD.n1874 VDD.t18 175.417
R2039 VDD.n301 VDD.t25 175.417
R2040 VDD.n1463 VDD.t55 175.417
R2041 VDD.n501 VDD.t44 175.417
R2042 VDD.n1935 VDD.t38 175.417
R2043 VDD.n318 VDD.t28 175.417
R2044 VDD.n1324 VDD.t52 175.417
R2045 VDD.n518 VDD.t41 175.417
R2046 VDD.n2709 VDD.n139 146.341
R2047 VDD.n2702 VDD.n2701 146.341
R2048 VDD.n2699 VDD.n2698 146.341
R2049 VDD.n2695 VDD.n2694 146.341
R2050 VDD.n2688 VDD.n2687 146.341
R2051 VDD.n2684 VDD.n2683 146.341
R2052 VDD.n2680 VDD.n2679 146.341
R2053 VDD.n2676 VDD.n2675 146.341
R2054 VDD.n2672 VDD.n2671 146.341
R2055 VDD.n2475 VDD.n272 146.341
R2056 VDD.n2481 VDD.n272 146.341
R2057 VDD.n2481 VDD.n264 146.341
R2058 VDD.n2491 VDD.n264 146.341
R2059 VDD.n2491 VDD.n260 146.341
R2060 VDD.n2497 VDD.n260 146.341
R2061 VDD.n2497 VDD.n252 146.341
R2062 VDD.n2507 VDD.n252 146.341
R2063 VDD.n2507 VDD.n248 146.341
R2064 VDD.n2513 VDD.n248 146.341
R2065 VDD.n2513 VDD.n240 146.341
R2066 VDD.n2523 VDD.n240 146.341
R2067 VDD.n2523 VDD.n236 146.341
R2068 VDD.n2529 VDD.n236 146.341
R2069 VDD.n2529 VDD.n228 146.341
R2070 VDD.n2539 VDD.n228 146.341
R2071 VDD.n2539 VDD.n224 146.341
R2072 VDD.n2545 VDD.n224 146.341
R2073 VDD.n2545 VDD.n215 146.341
R2074 VDD.n2555 VDD.n215 146.341
R2075 VDD.n2555 VDD.n211 146.341
R2076 VDD.n2561 VDD.n211 146.341
R2077 VDD.n2561 VDD.n204 146.341
R2078 VDD.n2571 VDD.n204 146.341
R2079 VDD.n2571 VDD.n200 146.341
R2080 VDD.n2577 VDD.n200 146.341
R2081 VDD.n2577 VDD.n192 146.341
R2082 VDD.n2587 VDD.n192 146.341
R2083 VDD.n2587 VDD.n187 146.341
R2084 VDD.n2596 VDD.n187 146.341
R2085 VDD.n2596 VDD.n188 146.341
R2086 VDD.n188 VDD.n179 146.341
R2087 VDD.n2607 VDD.n179 146.341
R2088 VDD.n2607 VDD.n41 146.341
R2089 VDD.n42 VDD.n41 146.341
R2090 VDD.n43 VDD.n42 146.341
R2091 VDD.n2614 VDD.n43 146.341
R2092 VDD.n2614 VDD.n51 146.341
R2093 VDD.n52 VDD.n51 146.341
R2094 VDD.n53 VDD.n52 146.341
R2095 VDD.n2621 VDD.n53 146.341
R2096 VDD.n2621 VDD.n62 146.341
R2097 VDD.n63 VDD.n62 146.341
R2098 VDD.n64 VDD.n63 146.341
R2099 VDD.n2628 VDD.n64 146.341
R2100 VDD.n2628 VDD.n73 146.341
R2101 VDD.n74 VDD.n73 146.341
R2102 VDD.n75 VDD.n74 146.341
R2103 VDD.n2635 VDD.n75 146.341
R2104 VDD.n2635 VDD.n84 146.341
R2105 VDD.n85 VDD.n84 146.341
R2106 VDD.n86 VDD.n85 146.341
R2107 VDD.n2642 VDD.n86 146.341
R2108 VDD.n2642 VDD.n95 146.341
R2109 VDD.n96 VDD.n95 146.341
R2110 VDD.n97 VDD.n96 146.341
R2111 VDD.n2649 VDD.n97 146.341
R2112 VDD.n2649 VDD.n106 146.341
R2113 VDD.n107 VDD.n106 146.341
R2114 VDD.n108 VDD.n107 146.341
R2115 VDD.n2656 VDD.n108 146.341
R2116 VDD.n2656 VDD.n117 146.341
R2117 VDD.n118 VDD.n117 146.341
R2118 VDD.n119 VDD.n118 146.341
R2119 VDD.n2663 VDD.n119 146.341
R2120 VDD.n2663 VDD.n128 146.341
R2121 VDD.n129 VDD.n128 146.341
R2122 VDD.n2467 VDD.n2465 146.341
R2123 VDD.n2465 VDD.n2464 146.341
R2124 VDD.n2461 VDD.n2460 146.341
R2125 VDD.n2458 VDD.n2410 146.341
R2126 VDD.n2453 VDD.n2451 146.341
R2127 VDD.n2449 VDD.n2418 146.341
R2128 VDD.n2445 VDD.n2443 146.341
R2129 VDD.n2441 VDD.n2424 146.341
R2130 VDD.n2432 VDD.n2429 146.341
R2131 VDD.n2473 VDD.n270 146.341
R2132 VDD.n2483 VDD.n270 146.341
R2133 VDD.n2483 VDD.n266 146.341
R2134 VDD.n2489 VDD.n266 146.341
R2135 VDD.n2489 VDD.n258 146.341
R2136 VDD.n2499 VDD.n258 146.341
R2137 VDD.n2499 VDD.n254 146.341
R2138 VDD.n2505 VDD.n254 146.341
R2139 VDD.n2505 VDD.n246 146.341
R2140 VDD.n2515 VDD.n246 146.341
R2141 VDD.n2515 VDD.n242 146.341
R2142 VDD.n2521 VDD.n242 146.341
R2143 VDD.n2521 VDD.n234 146.341
R2144 VDD.n2531 VDD.n234 146.341
R2145 VDD.n2531 VDD.n230 146.341
R2146 VDD.n2537 VDD.n230 146.341
R2147 VDD.n2537 VDD.n222 146.341
R2148 VDD.n2547 VDD.n222 146.341
R2149 VDD.n2547 VDD.n218 146.341
R2150 VDD.n2553 VDD.n218 146.341
R2151 VDD.n2553 VDD.n210 146.341
R2152 VDD.n2563 VDD.n210 146.341
R2153 VDD.n2563 VDD.n206 146.341
R2154 VDD.n2569 VDD.n206 146.341
R2155 VDD.n2569 VDD.n198 146.341
R2156 VDD.n2579 VDD.n198 146.341
R2157 VDD.n2579 VDD.n194 146.341
R2158 VDD.n2585 VDD.n194 146.341
R2159 VDD.n2585 VDD.n185 146.341
R2160 VDD.n2598 VDD.n185 146.341
R2161 VDD.n2598 VDD.n181 146.341
R2162 VDD.n2604 VDD.n181 146.341
R2163 VDD.n2604 VDD.n39 146.341
R2164 VDD.n2777 VDD.n39 146.341
R2165 VDD.n2777 VDD.n40 146.341
R2166 VDD.n2773 VDD.n40 146.341
R2167 VDD.n2773 VDD.n45 146.341
R2168 VDD.n2769 VDD.n45 146.341
R2169 VDD.n2769 VDD.n50 146.341
R2170 VDD.n2765 VDD.n50 146.341
R2171 VDD.n2765 VDD.n55 146.341
R2172 VDD.n2761 VDD.n55 146.341
R2173 VDD.n2761 VDD.n61 146.341
R2174 VDD.n2757 VDD.n61 146.341
R2175 VDD.n2757 VDD.n66 146.341
R2176 VDD.n2753 VDD.n66 146.341
R2177 VDD.n2753 VDD.n72 146.341
R2178 VDD.n2749 VDD.n72 146.341
R2179 VDD.n2749 VDD.n77 146.341
R2180 VDD.n2745 VDD.n77 146.341
R2181 VDD.n2745 VDD.n83 146.341
R2182 VDD.n2741 VDD.n83 146.341
R2183 VDD.n2741 VDD.n88 146.341
R2184 VDD.n2737 VDD.n88 146.341
R2185 VDD.n2737 VDD.n94 146.341
R2186 VDD.n2733 VDD.n94 146.341
R2187 VDD.n2733 VDD.n99 146.341
R2188 VDD.n2729 VDD.n99 146.341
R2189 VDD.n2729 VDD.n105 146.341
R2190 VDD.n2725 VDD.n105 146.341
R2191 VDD.n2725 VDD.n109 146.341
R2192 VDD.n2721 VDD.n109 146.341
R2193 VDD.n2721 VDD.n115 146.341
R2194 VDD.n2717 VDD.n115 146.341
R2195 VDD.n2717 VDD.n121 146.341
R2196 VDD.n2713 VDD.n121 146.341
R2197 VDD.n2713 VDD.n127 146.341
R2198 VDD.n1255 VDD.n1254 146.341
R2199 VDD.n1259 VDD.n1258 146.341
R2200 VDD.n1261 VDD.n1260 146.341
R2201 VDD.n1268 VDD.n1267 146.341
R2202 VDD.n1270 VDD.n1269 146.341
R2203 VDD.n1274 VDD.n1273 146.341
R2204 VDD.n1276 VDD.n1275 146.341
R2205 VDD.n1279 VDD.n1278 146.341
R2206 VDD.n1317 VDD.n688 146.341
R2207 VDD.n965 VDD.n887 146.341
R2208 VDD.n975 VDD.n887 146.341
R2209 VDD.n975 VDD.n883 146.341
R2210 VDD.n981 VDD.n883 146.341
R2211 VDD.n981 VDD.n875 146.341
R2212 VDD.n991 VDD.n875 146.341
R2213 VDD.n991 VDD.n871 146.341
R2214 VDD.n997 VDD.n871 146.341
R2215 VDD.n997 VDD.n863 146.341
R2216 VDD.n1007 VDD.n863 146.341
R2217 VDD.n1007 VDD.n859 146.341
R2218 VDD.n1013 VDD.n859 146.341
R2219 VDD.n1013 VDD.n851 146.341
R2220 VDD.n1023 VDD.n851 146.341
R2221 VDD.n1023 VDD.n847 146.341
R2222 VDD.n1029 VDD.n847 146.341
R2223 VDD.n1029 VDD.n839 146.341
R2224 VDD.n1039 VDD.n839 146.341
R2225 VDD.n1039 VDD.n835 146.341
R2226 VDD.n1045 VDD.n835 146.341
R2227 VDD.n1045 VDD.n828 146.341
R2228 VDD.n1056 VDD.n828 146.341
R2229 VDD.n1056 VDD.n824 146.341
R2230 VDD.n1062 VDD.n824 146.341
R2231 VDD.n1062 VDD.n816 146.341
R2232 VDD.n1072 VDD.n816 146.341
R2233 VDD.n1072 VDD.n812 146.341
R2234 VDD.n1078 VDD.n812 146.341
R2235 VDD.n1078 VDD.n804 146.341
R2236 VDD.n1088 VDD.n804 146.341
R2237 VDD.n1088 VDD.n800 146.341
R2238 VDD.n1094 VDD.n800 146.341
R2239 VDD.n1094 VDD.n793 146.341
R2240 VDD.n1126 VDD.n793 146.341
R2241 VDD.n1126 VDD.n789 146.341
R2242 VDD.n1132 VDD.n789 146.341
R2243 VDD.n1132 VDD.n781 146.341
R2244 VDD.n1142 VDD.n781 146.341
R2245 VDD.n1142 VDD.n777 146.341
R2246 VDD.n1148 VDD.n777 146.341
R2247 VDD.n1148 VDD.n769 146.341
R2248 VDD.n1158 VDD.n769 146.341
R2249 VDD.n1158 VDD.n765 146.341
R2250 VDD.n1164 VDD.n765 146.341
R2251 VDD.n1164 VDD.n758 146.341
R2252 VDD.n1175 VDD.n758 146.341
R2253 VDD.n1175 VDD.n754 146.341
R2254 VDD.n1181 VDD.n754 146.341
R2255 VDD.n1181 VDD.n746 146.341
R2256 VDD.n1191 VDD.n746 146.341
R2257 VDD.n1191 VDD.n742 146.341
R2258 VDD.n1197 VDD.n742 146.341
R2259 VDD.n1197 VDD.n734 146.341
R2260 VDD.n1207 VDD.n734 146.341
R2261 VDD.n1207 VDD.n730 146.341
R2262 VDD.n1213 VDD.n730 146.341
R2263 VDD.n1213 VDD.n722 146.341
R2264 VDD.n1223 VDD.n722 146.341
R2265 VDD.n1223 VDD.n718 146.341
R2266 VDD.n1229 VDD.n718 146.341
R2267 VDD.n1229 VDD.n710 146.341
R2268 VDD.n1239 VDD.n710 146.341
R2269 VDD.n1239 VDD.n706 146.341
R2270 VDD.n1246 VDD.n706 146.341
R2271 VDD.n1246 VDD.n696 146.341
R2272 VDD.n1311 VDD.n696 146.341
R2273 VDD.n1311 VDD.n689 146.341
R2274 VDD.n922 VDD.n918 146.341
R2275 VDD.n928 VDD.n918 146.341
R2276 VDD.n932 VDD.n930 146.341
R2277 VDD.n938 VDD.n911 146.341
R2278 VDD.n942 VDD.n940 146.341
R2279 VDD.n949 VDD.n907 146.341
R2280 VDD.n952 VDD.n951 146.341
R2281 VDD.n954 VDD.n905 146.341
R2282 VDD.n901 VDD.n897 146.341
R2283 VDD.n967 VDD.n889 146.341
R2284 VDD.n973 VDD.n889 146.341
R2285 VDD.n973 VDD.n881 146.341
R2286 VDD.n983 VDD.n881 146.341
R2287 VDD.n983 VDD.n877 146.341
R2288 VDD.n989 VDD.n877 146.341
R2289 VDD.n989 VDD.n869 146.341
R2290 VDD.n999 VDD.n869 146.341
R2291 VDD.n999 VDD.n865 146.341
R2292 VDD.n1005 VDD.n865 146.341
R2293 VDD.n1005 VDD.n857 146.341
R2294 VDD.n1015 VDD.n857 146.341
R2295 VDD.n1015 VDD.n853 146.341
R2296 VDD.n1021 VDD.n853 146.341
R2297 VDD.n1021 VDD.n845 146.341
R2298 VDD.n1031 VDD.n845 146.341
R2299 VDD.n1031 VDD.n841 146.341
R2300 VDD.n1037 VDD.n841 146.341
R2301 VDD.n1037 VDD.n833 146.341
R2302 VDD.n1048 VDD.n833 146.341
R2303 VDD.n1048 VDD.n829 146.341
R2304 VDD.n1054 VDD.n829 146.341
R2305 VDD.n1054 VDD.n822 146.341
R2306 VDD.n1064 VDD.n822 146.341
R2307 VDD.n1064 VDD.n818 146.341
R2308 VDD.n1070 VDD.n818 146.341
R2309 VDD.n1070 VDD.n810 146.341
R2310 VDD.n1080 VDD.n810 146.341
R2311 VDD.n1080 VDD.n806 146.341
R2312 VDD.n1086 VDD.n806 146.341
R2313 VDD.n1086 VDD.n798 146.341
R2314 VDD.n1097 VDD.n798 146.341
R2315 VDD.n1097 VDD.n794 146.341
R2316 VDD.n1124 VDD.n794 146.341
R2317 VDD.n1124 VDD.n787 146.341
R2318 VDD.n1134 VDD.n787 146.341
R2319 VDD.n1134 VDD.n783 146.341
R2320 VDD.n1140 VDD.n783 146.341
R2321 VDD.n1140 VDD.n775 146.341
R2322 VDD.n1150 VDD.n775 146.341
R2323 VDD.n1150 VDD.n771 146.341
R2324 VDD.n1156 VDD.n771 146.341
R2325 VDD.n1156 VDD.n763 146.341
R2326 VDD.n1167 VDD.n763 146.341
R2327 VDD.n1167 VDD.n759 146.341
R2328 VDD.n1173 VDD.n759 146.341
R2329 VDD.n1173 VDD.n752 146.341
R2330 VDD.n1183 VDD.n752 146.341
R2331 VDD.n1183 VDD.n748 146.341
R2332 VDD.n1189 VDD.n748 146.341
R2333 VDD.n1189 VDD.n740 146.341
R2334 VDD.n1199 VDD.n740 146.341
R2335 VDD.n1199 VDD.n736 146.341
R2336 VDD.n1205 VDD.n736 146.341
R2337 VDD.n1205 VDD.n728 146.341
R2338 VDD.n1215 VDD.n728 146.341
R2339 VDD.n1215 VDD.n724 146.341
R2340 VDD.n1221 VDD.n724 146.341
R2341 VDD.n1221 VDD.n716 146.341
R2342 VDD.n1231 VDD.n716 146.341
R2343 VDD.n1231 VDD.n712 146.341
R2344 VDD.n1237 VDD.n712 146.341
R2345 VDD.n1237 VDD.n704 146.341
R2346 VDD.n1248 VDD.n704 146.341
R2347 VDD.n1248 VDD.n698 146.341
R2348 VDD.n1309 VDD.n698 146.341
R2349 VDD.n1309 VDD.n699 146.341
R2350 VDD.t89 VDD.t115 132.423
R2351 VDD.t56 VDD.t105 132.423
R2352 VDD.n9 VDD.n7 127.225
R2353 VDD.n2 VDD.n0 127.225
R2354 VDD.n9 VDD.n8 126.035
R2355 VDD.n11 VDD.n10 126.035
R2356 VDD.n13 VDD.n12 126.035
R2357 VDD.n6 VDD.n5 126.035
R2358 VDD.n4 VDD.n3 126.035
R2359 VDD.n2 VDD.n1 126.035
R2360 VDD.n1859 VDD.n1858 124.856
R2361 VDD.n1875 VDD.t17 121.889
R2362 VDD.n302 VDD.t26 121.889
R2363 VDD.n1464 VDD.t54 121.889
R2364 VDD.n502 VDD.t45 121.889
R2365 VDD.n1936 VDD.t37 121.889
R2366 VDD.n319 VDD.t29 121.889
R2367 VDD.n1325 VDD.t51 121.889
R2368 VDD.n519 VDD.t42 121.889
R2369 VDD.n899 VDD.n898 120.243
R2370 VDD.n914 VDD.n913 120.243
R2371 VDD.n2415 VDD.n2414 120.243
R2372 VDD.n2434 VDD.n2433 120.243
R2373 VDD.n159 VDD.n158 120.243
R2374 VDD.n2691 VDD.n2690 120.243
R2375 VDD.n1265 VDD.n1264 120.243
R2376 VDD.n691 VDD.n690 120.243
R2377 VDD.n2133 VDD.n470 99.5127
R2378 VDD.n2141 VDD.n470 99.5127
R2379 VDD.n2141 VDD.n468 99.5127
R2380 VDD.n2145 VDD.n468 99.5127
R2381 VDD.n2145 VDD.n459 99.5127
R2382 VDD.n2153 VDD.n459 99.5127
R2383 VDD.n2153 VDD.n457 99.5127
R2384 VDD.n2157 VDD.n457 99.5127
R2385 VDD.n2157 VDD.n447 99.5127
R2386 VDD.n2165 VDD.n447 99.5127
R2387 VDD.n2165 VDD.n445 99.5127
R2388 VDD.n2169 VDD.n445 99.5127
R2389 VDD.n2169 VDD.n435 99.5127
R2390 VDD.n2177 VDD.n435 99.5127
R2391 VDD.n2177 VDD.n433 99.5127
R2392 VDD.n2181 VDD.n433 99.5127
R2393 VDD.n2181 VDD.n424 99.5127
R2394 VDD.n2189 VDD.n424 99.5127
R2395 VDD.n2189 VDD.n422 99.5127
R2396 VDD.n2193 VDD.n422 99.5127
R2397 VDD.n2193 VDD.n412 99.5127
R2398 VDD.n2201 VDD.n412 99.5127
R2399 VDD.n2201 VDD.n410 99.5127
R2400 VDD.n2205 VDD.n410 99.5127
R2401 VDD.n2205 VDD.n400 99.5127
R2402 VDD.n2213 VDD.n400 99.5127
R2403 VDD.n2213 VDD.n398 99.5127
R2404 VDD.n2217 VDD.n398 99.5127
R2405 VDD.n2217 VDD.n388 99.5127
R2406 VDD.n2225 VDD.n388 99.5127
R2407 VDD.n2225 VDD.n386 99.5127
R2408 VDD.n2229 VDD.n386 99.5127
R2409 VDD.n2229 VDD.n376 99.5127
R2410 VDD.n2237 VDD.n376 99.5127
R2411 VDD.n2237 VDD.n374 99.5127
R2412 VDD.n2241 VDD.n374 99.5127
R2413 VDD.n2241 VDD.n364 99.5127
R2414 VDD.n2249 VDD.n364 99.5127
R2415 VDD.n2249 VDD.n362 99.5127
R2416 VDD.n2253 VDD.n362 99.5127
R2417 VDD.n2253 VDD.n352 99.5127
R2418 VDD.n2261 VDD.n352 99.5127
R2419 VDD.n2261 VDD.n350 99.5127
R2420 VDD.n2265 VDD.n350 99.5127
R2421 VDD.n2265 VDD.n340 99.5127
R2422 VDD.n2273 VDD.n340 99.5127
R2423 VDD.n2273 VDD.n338 99.5127
R2424 VDD.n2277 VDD.n338 99.5127
R2425 VDD.n2277 VDD.n327 99.5127
R2426 VDD.n2287 VDD.n327 99.5127
R2427 VDD.n2287 VDD.n325 99.5127
R2428 VDD.n2291 VDD.n325 99.5127
R2429 VDD.n2291 VDD.n311 99.5127
R2430 VDD.n2350 VDD.n311 99.5127
R2431 VDD.n2350 VDD.n309 99.5127
R2432 VDD.n2354 VDD.n309 99.5127
R2433 VDD.n2354 VDD.n298 99.5127
R2434 VDD.n2399 VDD.n299 99.5127
R2435 VDD.n2395 VDD.n2394 99.5127
R2436 VDD.n2391 VDD.n2390 99.5127
R2437 VDD.n2387 VDD.n2386 99.5127
R2438 VDD.n2383 VDD.n2382 99.5127
R2439 VDD.n2379 VDD.n2378 99.5127
R2440 VDD.n2375 VDD.n2374 99.5127
R2441 VDD.n2371 VDD.n2370 99.5127
R2442 VDD.n2367 VDD.n2366 99.5127
R2443 VDD.n2362 VDD.n2361 99.5127
R2444 VDD.n2088 VDD.n1860 99.5127
R2445 VDD.n2088 VDD.n471 99.5127
R2446 VDD.n2085 VDD.n471 99.5127
R2447 VDD.n2085 VDD.n466 99.5127
R2448 VDD.n2082 VDD.n466 99.5127
R2449 VDD.n2082 VDD.n460 99.5127
R2450 VDD.n2079 VDD.n460 99.5127
R2451 VDD.n2079 VDD.n454 99.5127
R2452 VDD.n2076 VDD.n454 99.5127
R2453 VDD.n2076 VDD.n448 99.5127
R2454 VDD.n2073 VDD.n448 99.5127
R2455 VDD.n2073 VDD.n443 99.5127
R2456 VDD.n2070 VDD.n443 99.5127
R2457 VDD.n2070 VDD.n437 99.5127
R2458 VDD.n2067 VDD.n437 99.5127
R2459 VDD.n2067 VDD.n431 99.5127
R2460 VDD.n2064 VDD.n431 99.5127
R2461 VDD.n2064 VDD.n425 99.5127
R2462 VDD.n1930 VDD.n425 99.5127
R2463 VDD.n1930 VDD.n420 99.5127
R2464 VDD.n1927 VDD.n420 99.5127
R2465 VDD.n1927 VDD.n414 99.5127
R2466 VDD.n1924 VDD.n414 99.5127
R2467 VDD.n1924 VDD.n408 99.5127
R2468 VDD.n1921 VDD.n408 99.5127
R2469 VDD.n1921 VDD.n402 99.5127
R2470 VDD.n1918 VDD.n402 99.5127
R2471 VDD.n1918 VDD.n396 99.5127
R2472 VDD.n1915 VDD.n396 99.5127
R2473 VDD.n1915 VDD.n390 99.5127
R2474 VDD.n1912 VDD.n390 99.5127
R2475 VDD.n1912 VDD.n384 99.5127
R2476 VDD.n1909 VDD.n384 99.5127
R2477 VDD.n1909 VDD.n378 99.5127
R2478 VDD.n1906 VDD.n378 99.5127
R2479 VDD.n1906 VDD.n372 99.5127
R2480 VDD.n1903 VDD.n372 99.5127
R2481 VDD.n1903 VDD.n366 99.5127
R2482 VDD.n1900 VDD.n366 99.5127
R2483 VDD.n1900 VDD.n360 99.5127
R2484 VDD.n1897 VDD.n360 99.5127
R2485 VDD.n1897 VDD.n354 99.5127
R2486 VDD.n1894 VDD.n354 99.5127
R2487 VDD.n1894 VDD.n348 99.5127
R2488 VDD.n1891 VDD.n348 99.5127
R2489 VDD.n1891 VDD.n342 99.5127
R2490 VDD.n1888 VDD.n342 99.5127
R2491 VDD.n1888 VDD.n336 99.5127
R2492 VDD.n1885 VDD.n336 99.5127
R2493 VDD.n1885 VDD.n329 99.5127
R2494 VDD.n1882 VDD.n329 99.5127
R2495 VDD.n1882 VDD.n324 99.5127
R2496 VDD.n1879 VDD.n324 99.5127
R2497 VDD.n1879 VDD.n313 99.5127
R2498 VDD.n313 VDD.n304 99.5127
R2499 VDD.n2356 VDD.n304 99.5127
R2500 VDD.n2357 VDD.n2356 99.5127
R2501 VDD.n2129 VDD.n2127 99.5127
R2502 VDD.n2127 VDD.n2126 99.5127
R2503 VDD.n2123 VDD.n2122 99.5127
R2504 VDD.n2120 VDD.n1867 99.5127
R2505 VDD.n2116 VDD.n2114 99.5127
R2506 VDD.n2112 VDD.n1869 99.5127
R2507 VDD.n2108 VDD.n2106 99.5127
R2508 VDD.n2104 VDD.n1871 99.5127
R2509 VDD.n2100 VDD.n2098 99.5127
R2510 VDD.n2096 VDD.n1873 99.5127
R2511 VDD.n1857 VDD.n499 99.5127
R2512 VDD.n1853 VDD.n1852 99.5127
R2513 VDD.n1849 VDD.n1848 99.5127
R2514 VDD.n1845 VDD.n1844 99.5127
R2515 VDD.n1841 VDD.n1840 99.5127
R2516 VDD.n1837 VDD.n1836 99.5127
R2517 VDD.n1833 VDD.n1832 99.5127
R2518 VDD.n1829 VDD.n1828 99.5127
R2519 VDD.n1825 VDD.n1824 99.5127
R2520 VDD.n1820 VDD.n1819 99.5127
R2521 VDD.n1546 VDD.n1320 99.5127
R2522 VDD.n1546 VDD.n673 99.5127
R2523 VDD.n1543 VDD.n673 99.5127
R2524 VDD.n1543 VDD.n667 99.5127
R2525 VDD.n1540 VDD.n667 99.5127
R2526 VDD.n1540 VDD.n661 99.5127
R2527 VDD.n1537 VDD.n661 99.5127
R2528 VDD.n1537 VDD.n656 99.5127
R2529 VDD.n1534 VDD.n656 99.5127
R2530 VDD.n1534 VDD.n650 99.5127
R2531 VDD.n1531 VDD.n650 99.5127
R2532 VDD.n1531 VDD.n644 99.5127
R2533 VDD.n1528 VDD.n644 99.5127
R2534 VDD.n1528 VDD.n638 99.5127
R2535 VDD.n1525 VDD.n638 99.5127
R2536 VDD.n1525 VDD.n632 99.5127
R2537 VDD.n1522 VDD.n632 99.5127
R2538 VDD.n1522 VDD.n626 99.5127
R2539 VDD.n1519 VDD.n626 99.5127
R2540 VDD.n1519 VDD.n620 99.5127
R2541 VDD.n1516 VDD.n620 99.5127
R2542 VDD.n1516 VDD.n614 99.5127
R2543 VDD.n1513 VDD.n614 99.5127
R2544 VDD.n1513 VDD.n608 99.5127
R2545 VDD.n1510 VDD.n608 99.5127
R2546 VDD.n1510 VDD.n602 99.5127
R2547 VDD.n1507 VDD.n602 99.5127
R2548 VDD.n1507 VDD.n596 99.5127
R2549 VDD.n1504 VDD.n596 99.5127
R2550 VDD.n1504 VDD.n590 99.5127
R2551 VDD.n1501 VDD.n590 99.5127
R2552 VDD.n1501 VDD.n584 99.5127
R2553 VDD.n1498 VDD.n584 99.5127
R2554 VDD.n1498 VDD.n578 99.5127
R2555 VDD.n1495 VDD.n578 99.5127
R2556 VDD.n1495 VDD.n572 99.5127
R2557 VDD.n1492 VDD.n572 99.5127
R2558 VDD.n1492 VDD.n565 99.5127
R2559 VDD.n1489 VDD.n565 99.5127
R2560 VDD.n1489 VDD.n559 99.5127
R2561 VDD.n1486 VDD.n559 99.5127
R2562 VDD.n1486 VDD.n554 99.5127
R2563 VDD.n1483 VDD.n554 99.5127
R2564 VDD.n1483 VDD.n548 99.5127
R2565 VDD.n1480 VDD.n548 99.5127
R2566 VDD.n1480 VDD.n541 99.5127
R2567 VDD.n1477 VDD.n541 99.5127
R2568 VDD.n1477 VDD.n535 99.5127
R2569 VDD.n1474 VDD.n535 99.5127
R2570 VDD.n1474 VDD.n529 99.5127
R2571 VDD.n1471 VDD.n529 99.5127
R2572 VDD.n1471 VDD.n524 99.5127
R2573 VDD.n1468 VDD.n524 99.5127
R2574 VDD.n1468 VDD.n512 99.5127
R2575 VDD.n512 VDD.n504 99.5127
R2576 VDD.n1814 VDD.n504 99.5127
R2577 VDD.n1815 VDD.n1814 99.5127
R2578 VDD.n1587 VDD.n1585 99.5127
R2579 VDD.n1585 VDD.n1584 99.5127
R2580 VDD.n1581 VDD.n1580 99.5127
R2581 VDD.n1578 VDD.n1456 99.5127
R2582 VDD.n1574 VDD.n1572 99.5127
R2583 VDD.n1570 VDD.n1458 99.5127
R2584 VDD.n1566 VDD.n1564 99.5127
R2585 VDD.n1562 VDD.n1460 99.5127
R2586 VDD.n1558 VDD.n1556 99.5127
R2587 VDD.n1554 VDD.n1462 99.5127
R2588 VDD.n1591 VDD.n671 99.5127
R2589 VDD.n1599 VDD.n671 99.5127
R2590 VDD.n1599 VDD.n669 99.5127
R2591 VDD.n1603 VDD.n669 99.5127
R2592 VDD.n1603 VDD.n660 99.5127
R2593 VDD.n1611 VDD.n660 99.5127
R2594 VDD.n1611 VDD.n658 99.5127
R2595 VDD.n1615 VDD.n658 99.5127
R2596 VDD.n1615 VDD.n648 99.5127
R2597 VDD.n1623 VDD.n648 99.5127
R2598 VDD.n1623 VDD.n646 99.5127
R2599 VDD.n1627 VDD.n646 99.5127
R2600 VDD.n1627 VDD.n636 99.5127
R2601 VDD.n1635 VDD.n636 99.5127
R2602 VDD.n1635 VDD.n634 99.5127
R2603 VDD.n1639 VDD.n634 99.5127
R2604 VDD.n1639 VDD.n624 99.5127
R2605 VDD.n1647 VDD.n624 99.5127
R2606 VDD.n1647 VDD.n622 99.5127
R2607 VDD.n1651 VDD.n622 99.5127
R2608 VDD.n1651 VDD.n612 99.5127
R2609 VDD.n1659 VDD.n612 99.5127
R2610 VDD.n1659 VDD.n610 99.5127
R2611 VDD.n1663 VDD.n610 99.5127
R2612 VDD.n1663 VDD.n600 99.5127
R2613 VDD.n1671 VDD.n600 99.5127
R2614 VDD.n1671 VDD.n598 99.5127
R2615 VDD.n1675 VDD.n598 99.5127
R2616 VDD.n1675 VDD.n588 99.5127
R2617 VDD.n1683 VDD.n588 99.5127
R2618 VDD.n1683 VDD.n586 99.5127
R2619 VDD.n1687 VDD.n586 99.5127
R2620 VDD.n1687 VDD.n576 99.5127
R2621 VDD.n1695 VDD.n576 99.5127
R2622 VDD.n1695 VDD.n574 99.5127
R2623 VDD.n1699 VDD.n574 99.5127
R2624 VDD.n1699 VDD.n563 99.5127
R2625 VDD.n1707 VDD.n563 99.5127
R2626 VDD.n1707 VDD.n561 99.5127
R2627 VDD.n1711 VDD.n561 99.5127
R2628 VDD.n1711 VDD.n552 99.5127
R2629 VDD.n1719 VDD.n552 99.5127
R2630 VDD.n1719 VDD.n550 99.5127
R2631 VDD.n1723 VDD.n550 99.5127
R2632 VDD.n1723 VDD.n539 99.5127
R2633 VDD.n1731 VDD.n539 99.5127
R2634 VDD.n1731 VDD.n537 99.5127
R2635 VDD.n1735 VDD.n537 99.5127
R2636 VDD.n1735 VDD.n527 99.5127
R2637 VDD.n1745 VDD.n527 99.5127
R2638 VDD.n1745 VDD.n525 99.5127
R2639 VDD.n1749 VDD.n525 99.5127
R2640 VDD.n1749 VDD.n510 99.5127
R2641 VDD.n1808 VDD.n510 99.5127
R2642 VDD.n1808 VDD.n508 99.5127
R2643 VDD.n1812 VDD.n508 99.5127
R2644 VDD.n1812 VDD.n498 99.5127
R2645 VDD.n2340 VDD.n277 99.5127
R2646 VDD.n2338 VDD.n2337 99.5127
R2647 VDD.n2334 VDD.n2333 99.5127
R2648 VDD.n2330 VDD.n2329 99.5127
R2649 VDD.n2326 VDD.n2325 99.5127
R2650 VDD.n2322 VDD.n2321 99.5127
R2651 VDD.n2318 VDD.n2317 99.5127
R2652 VDD.n2314 VDD.n2313 99.5127
R2653 VDD.n2310 VDD.n2309 99.5127
R2654 VDD.n2305 VDD.n2304 99.5127
R2655 VDD.n1987 VDD.n1861 99.5127
R2656 VDD.n1987 VDD.n472 99.5127
R2657 VDD.n1990 VDD.n472 99.5127
R2658 VDD.n1990 VDD.n467 99.5127
R2659 VDD.n1993 VDD.n467 99.5127
R2660 VDD.n1993 VDD.n461 99.5127
R2661 VDD.n1996 VDD.n461 99.5127
R2662 VDD.n1996 VDD.n455 99.5127
R2663 VDD.n1999 VDD.n455 99.5127
R2664 VDD.n1999 VDD.n449 99.5127
R2665 VDD.n2002 VDD.n449 99.5127
R2666 VDD.n2002 VDD.n444 99.5127
R2667 VDD.n2005 VDD.n444 99.5127
R2668 VDD.n2005 VDD.n438 99.5127
R2669 VDD.n2008 VDD.n438 99.5127
R2670 VDD.n2008 VDD.n432 99.5127
R2671 VDD.n2062 VDD.n432 99.5127
R2672 VDD.n2062 VDD.n426 99.5127
R2673 VDD.n2058 VDD.n426 99.5127
R2674 VDD.n2058 VDD.n421 99.5127
R2675 VDD.n2055 VDD.n421 99.5127
R2676 VDD.n2055 VDD.n415 99.5127
R2677 VDD.n2052 VDD.n415 99.5127
R2678 VDD.n2052 VDD.n409 99.5127
R2679 VDD.n2049 VDD.n409 99.5127
R2680 VDD.n2049 VDD.n403 99.5127
R2681 VDD.n2046 VDD.n403 99.5127
R2682 VDD.n2046 VDD.n397 99.5127
R2683 VDD.n2043 VDD.n397 99.5127
R2684 VDD.n2043 VDD.n391 99.5127
R2685 VDD.n2040 VDD.n391 99.5127
R2686 VDD.n2040 VDD.n385 99.5127
R2687 VDD.n2037 VDD.n385 99.5127
R2688 VDD.n2037 VDD.n379 99.5127
R2689 VDD.n2034 VDD.n379 99.5127
R2690 VDD.n2034 VDD.n373 99.5127
R2691 VDD.n2031 VDD.n373 99.5127
R2692 VDD.n2031 VDD.n367 99.5127
R2693 VDD.n2028 VDD.n367 99.5127
R2694 VDD.n2028 VDD.n361 99.5127
R2695 VDD.n2025 VDD.n361 99.5127
R2696 VDD.n2025 VDD.n355 99.5127
R2697 VDD.n2022 VDD.n355 99.5127
R2698 VDD.n2022 VDD.n349 99.5127
R2699 VDD.n2019 VDD.n349 99.5127
R2700 VDD.n2019 VDD.n343 99.5127
R2701 VDD.n2016 VDD.n343 99.5127
R2702 VDD.n2016 VDD.n337 99.5127
R2703 VDD.n2013 VDD.n337 99.5127
R2704 VDD.n2013 VDD.n330 99.5127
R2705 VDD.n330 VDD.n321 99.5127
R2706 VDD.n2292 VDD.n321 99.5127
R2707 VDD.n2293 VDD.n2292 99.5127
R2708 VDD.n2293 VDD.n314 99.5127
R2709 VDD.n2296 VDD.n314 99.5127
R2710 VDD.n2296 VDD.n307 99.5127
R2711 VDD.n2300 VDD.n307 99.5127
R2712 VDD.n1948 VDD.n1945 99.5127
R2713 VDD.n1952 VDD.n1950 99.5127
R2714 VDD.n1956 VDD.n1942 99.5127
R2715 VDD.n1960 VDD.n1958 99.5127
R2716 VDD.n1964 VDD.n1940 99.5127
R2717 VDD.n1968 VDD.n1966 99.5127
R2718 VDD.n1972 VDD.n1938 99.5127
R2719 VDD.n1976 VDD.n1974 99.5127
R2720 VDD.n1981 VDD.n1934 99.5127
R2721 VDD.n1984 VDD.n1983 99.5127
R2722 VDD.n2135 VDD.n473 99.5127
R2723 VDD.n2139 VDD.n473 99.5127
R2724 VDD.n2139 VDD.n464 99.5127
R2725 VDD.n2147 VDD.n464 99.5127
R2726 VDD.n2147 VDD.n462 99.5127
R2727 VDD.n2151 VDD.n462 99.5127
R2728 VDD.n2151 VDD.n452 99.5127
R2729 VDD.n2159 VDD.n452 99.5127
R2730 VDD.n2159 VDD.n450 99.5127
R2731 VDD.n2163 VDD.n450 99.5127
R2732 VDD.n2163 VDD.n441 99.5127
R2733 VDD.n2171 VDD.n441 99.5127
R2734 VDD.n2171 VDD.n439 99.5127
R2735 VDD.n2175 VDD.n439 99.5127
R2736 VDD.n2175 VDD.n429 99.5127
R2737 VDD.n2183 VDD.n429 99.5127
R2738 VDD.n2183 VDD.n427 99.5127
R2739 VDD.n2187 VDD.n427 99.5127
R2740 VDD.n2187 VDD.n418 99.5127
R2741 VDD.n2195 VDD.n418 99.5127
R2742 VDD.n2195 VDD.n416 99.5127
R2743 VDD.n2199 VDD.n416 99.5127
R2744 VDD.n2199 VDD.n406 99.5127
R2745 VDD.n2207 VDD.n406 99.5127
R2746 VDD.n2207 VDD.n404 99.5127
R2747 VDD.n2211 VDD.n404 99.5127
R2748 VDD.n2211 VDD.n394 99.5127
R2749 VDD.n2219 VDD.n394 99.5127
R2750 VDD.n2219 VDD.n392 99.5127
R2751 VDD.n2223 VDD.n392 99.5127
R2752 VDD.n2223 VDD.n382 99.5127
R2753 VDD.n2231 VDD.n382 99.5127
R2754 VDD.n2231 VDD.n380 99.5127
R2755 VDD.n2235 VDD.n380 99.5127
R2756 VDD.n2235 VDD.n370 99.5127
R2757 VDD.n2243 VDD.n370 99.5127
R2758 VDD.n2243 VDD.n368 99.5127
R2759 VDD.n2247 VDD.n368 99.5127
R2760 VDD.n2247 VDD.n358 99.5127
R2761 VDD.n2255 VDD.n358 99.5127
R2762 VDD.n2255 VDD.n356 99.5127
R2763 VDD.n2259 VDD.n356 99.5127
R2764 VDD.n2259 VDD.n346 99.5127
R2765 VDD.n2267 VDD.n346 99.5127
R2766 VDD.n2267 VDD.n344 99.5127
R2767 VDD.n2271 VDD.n344 99.5127
R2768 VDD.n2271 VDD.n334 99.5127
R2769 VDD.n2279 VDD.n334 99.5127
R2770 VDD.n2279 VDD.n331 99.5127
R2771 VDD.n2285 VDD.n331 99.5127
R2772 VDD.n2285 VDD.n332 99.5127
R2773 VDD.n332 VDD.n323 99.5127
R2774 VDD.n323 VDD.n315 99.5127
R2775 VDD.n2348 VDD.n315 99.5127
R2776 VDD.n2348 VDD.n316 99.5127
R2777 VDD.n316 VDD.n308 99.5127
R2778 VDD.n2343 VDD.n308 99.5127
R2779 VDD.n1798 VDD.n477 99.5127
R2780 VDD.n1796 VDD.n1795 99.5127
R2781 VDD.n1792 VDD.n1791 99.5127
R2782 VDD.n1788 VDD.n1787 99.5127
R2783 VDD.n1784 VDD.n1783 99.5127
R2784 VDD.n1780 VDD.n1779 99.5127
R2785 VDD.n1776 VDD.n1775 99.5127
R2786 VDD.n1772 VDD.n1771 99.5127
R2787 VDD.n1768 VDD.n1767 99.5127
R2788 VDD.n1763 VDD.n1762 99.5127
R2789 VDD.n1451 VDD.n1322 99.5127
R2790 VDD.n1322 VDD.n674 99.5127
R2791 VDD.n1446 VDD.n674 99.5127
R2792 VDD.n1446 VDD.n668 99.5127
R2793 VDD.n1443 VDD.n668 99.5127
R2794 VDD.n1443 VDD.n662 99.5127
R2795 VDD.n1440 VDD.n662 99.5127
R2796 VDD.n1440 VDD.n657 99.5127
R2797 VDD.n1437 VDD.n657 99.5127
R2798 VDD.n1437 VDD.n651 99.5127
R2799 VDD.n1434 VDD.n651 99.5127
R2800 VDD.n1434 VDD.n645 99.5127
R2801 VDD.n1431 VDD.n645 99.5127
R2802 VDD.n1431 VDD.n639 99.5127
R2803 VDD.n1428 VDD.n639 99.5127
R2804 VDD.n1428 VDD.n633 99.5127
R2805 VDD.n1425 VDD.n633 99.5127
R2806 VDD.n1425 VDD.n627 99.5127
R2807 VDD.n1422 VDD.n627 99.5127
R2808 VDD.n1422 VDD.n621 99.5127
R2809 VDD.n1419 VDD.n621 99.5127
R2810 VDD.n1419 VDD.n615 99.5127
R2811 VDD.n1416 VDD.n615 99.5127
R2812 VDD.n1416 VDD.n609 99.5127
R2813 VDD.n1413 VDD.n609 99.5127
R2814 VDD.n1413 VDD.n603 99.5127
R2815 VDD.n1410 VDD.n603 99.5127
R2816 VDD.n1410 VDD.n597 99.5127
R2817 VDD.n1407 VDD.n597 99.5127
R2818 VDD.n1407 VDD.n591 99.5127
R2819 VDD.n1404 VDD.n591 99.5127
R2820 VDD.n1404 VDD.n585 99.5127
R2821 VDD.n1401 VDD.n585 99.5127
R2822 VDD.n1401 VDD.n579 99.5127
R2823 VDD.n1398 VDD.n579 99.5127
R2824 VDD.n1398 VDD.n573 99.5127
R2825 VDD.n1395 VDD.n573 99.5127
R2826 VDD.n1395 VDD.n566 99.5127
R2827 VDD.n1392 VDD.n566 99.5127
R2828 VDD.n1392 VDD.n560 99.5127
R2829 VDD.n1389 VDD.n560 99.5127
R2830 VDD.n1389 VDD.n555 99.5127
R2831 VDD.n1386 VDD.n555 99.5127
R2832 VDD.n1386 VDD.n549 99.5127
R2833 VDD.n1383 VDD.n549 99.5127
R2834 VDD.n1383 VDD.n542 99.5127
R2835 VDD.n1380 VDD.n542 99.5127
R2836 VDD.n1380 VDD.n536 99.5127
R2837 VDD.n1377 VDD.n536 99.5127
R2838 VDD.n1377 VDD.n530 99.5127
R2839 VDD.n530 VDD.n521 99.5127
R2840 VDD.n1750 VDD.n521 99.5127
R2841 VDD.n1751 VDD.n1750 99.5127
R2842 VDD.n1751 VDD.n513 99.5127
R2843 VDD.n1754 VDD.n513 99.5127
R2844 VDD.n1754 VDD.n506 99.5127
R2845 VDD.n1758 VDD.n506 99.5127
R2846 VDD.n1339 VDD.n1337 99.5127
R2847 VDD.n1343 VDD.n1334 99.5127
R2848 VDD.n1347 VDD.n1345 99.5127
R2849 VDD.n1351 VDD.n1332 99.5127
R2850 VDD.n1355 VDD.n1353 99.5127
R2851 VDD.n1359 VDD.n1330 99.5127
R2852 VDD.n1363 VDD.n1361 99.5127
R2853 VDD.n1367 VDD.n1328 99.5127
R2854 VDD.n1370 VDD.n1369 99.5127
R2855 VDD.n1372 VDD.n1321 99.5127
R2856 VDD.n1593 VDD.n675 99.5127
R2857 VDD.n1597 VDD.n675 99.5127
R2858 VDD.n1597 VDD.n665 99.5127
R2859 VDD.n1605 VDD.n665 99.5127
R2860 VDD.n1605 VDD.n663 99.5127
R2861 VDD.n1609 VDD.n663 99.5127
R2862 VDD.n1609 VDD.n654 99.5127
R2863 VDD.n1617 VDD.n654 99.5127
R2864 VDD.n1617 VDD.n652 99.5127
R2865 VDD.n1621 VDD.n652 99.5127
R2866 VDD.n1621 VDD.n642 99.5127
R2867 VDD.n1629 VDD.n642 99.5127
R2868 VDD.n1629 VDD.n640 99.5127
R2869 VDD.n1633 VDD.n640 99.5127
R2870 VDD.n1633 VDD.n630 99.5127
R2871 VDD.n1641 VDD.n630 99.5127
R2872 VDD.n1641 VDD.n628 99.5127
R2873 VDD.n1645 VDD.n628 99.5127
R2874 VDD.n1645 VDD.n618 99.5127
R2875 VDD.n1653 VDD.n618 99.5127
R2876 VDD.n1653 VDD.n616 99.5127
R2877 VDD.n1657 VDD.n616 99.5127
R2878 VDD.n1657 VDD.n606 99.5127
R2879 VDD.n1665 VDD.n606 99.5127
R2880 VDD.n1665 VDD.n604 99.5127
R2881 VDD.n1669 VDD.n604 99.5127
R2882 VDD.n1669 VDD.n594 99.5127
R2883 VDD.n1677 VDD.n594 99.5127
R2884 VDD.n1677 VDD.n592 99.5127
R2885 VDD.n1681 VDD.n592 99.5127
R2886 VDD.n1681 VDD.n582 99.5127
R2887 VDD.n1689 VDD.n582 99.5127
R2888 VDD.n1689 VDD.n580 99.5127
R2889 VDD.n1693 VDD.n580 99.5127
R2890 VDD.n1693 VDD.n570 99.5127
R2891 VDD.n1701 VDD.n570 99.5127
R2892 VDD.n1701 VDD.n568 99.5127
R2893 VDD.n1705 VDD.n568 99.5127
R2894 VDD.n1705 VDD.n558 99.5127
R2895 VDD.n1713 VDD.n558 99.5127
R2896 VDD.n1713 VDD.n556 99.5127
R2897 VDD.n1717 VDD.n556 99.5127
R2898 VDD.n1717 VDD.n546 99.5127
R2899 VDD.n1725 VDD.n546 99.5127
R2900 VDD.n1725 VDD.n544 99.5127
R2901 VDD.n1729 VDD.n544 99.5127
R2902 VDD.n1729 VDD.n534 99.5127
R2903 VDD.n1737 VDD.n534 99.5127
R2904 VDD.n1737 VDD.n531 99.5127
R2905 VDD.n1743 VDD.n531 99.5127
R2906 VDD.n1743 VDD.n532 99.5127
R2907 VDD.n532 VDD.n523 99.5127
R2908 VDD.n523 VDD.n515 99.5127
R2909 VDD.n1806 VDD.n515 99.5127
R2910 VDD.n1806 VDD.n516 99.5127
R2911 VDD.n516 VDD.n507 99.5127
R2912 VDD.n1801 VDD.n507 99.5127
R2913 VDD.n28 VDD.t63 85.8723
R2914 VDD.n19 VDD.t74 85.8723
R2915 VDD.n1112 VDD.t60 85.8723
R2916 VDD.n1103 VDD.t73 85.8723
R2917 VDD.n1336 VDD.n1319 72.8958
R2918 VDD.n1338 VDD.n1319 72.8958
R2919 VDD.n1344 VDD.n1319 72.8958
R2920 VDD.n1346 VDD.n1319 72.8958
R2921 VDD.n1352 VDD.n1319 72.8958
R2922 VDD.n1354 VDD.n1319 72.8958
R2923 VDD.n1360 VDD.n1319 72.8958
R2924 VDD.n1362 VDD.n1319 72.8958
R2925 VDD.n1368 VDD.n1319 72.8958
R2926 VDD.n1371 VDD.n1319 72.8958
R2927 VDD.n1858 VDD.n487 72.8958
R2928 VDD.n1858 VDD.n486 72.8958
R2929 VDD.n1858 VDD.n485 72.8958
R2930 VDD.n1858 VDD.n484 72.8958
R2931 VDD.n1858 VDD.n483 72.8958
R2932 VDD.n1858 VDD.n482 72.8958
R2933 VDD.n1858 VDD.n481 72.8958
R2934 VDD.n1858 VDD.n480 72.8958
R2935 VDD.n1858 VDD.n479 72.8958
R2936 VDD.n1858 VDD.n478 72.8958
R2937 VDD.n1944 VDD.n1859 72.8958
R2938 VDD.n1949 VDD.n1859 72.8958
R2939 VDD.n1951 VDD.n1859 72.8958
R2940 VDD.n1957 VDD.n1859 72.8958
R2941 VDD.n1959 VDD.n1859 72.8958
R2942 VDD.n1965 VDD.n1859 72.8958
R2943 VDD.n1967 VDD.n1859 72.8958
R2944 VDD.n1973 VDD.n1859 72.8958
R2945 VDD.n1975 VDD.n1859 72.8958
R2946 VDD.n1982 VDD.n1859 72.8958
R2947 VDD.n2400 VDD.n287 72.8958
R2948 VDD.n2400 VDD.n286 72.8958
R2949 VDD.n2400 VDD.n285 72.8958
R2950 VDD.n2400 VDD.n284 72.8958
R2951 VDD.n2400 VDD.n283 72.8958
R2952 VDD.n2400 VDD.n282 72.8958
R2953 VDD.n2400 VDD.n281 72.8958
R2954 VDD.n2400 VDD.n280 72.8958
R2955 VDD.n2400 VDD.n279 72.8958
R2956 VDD.n2400 VDD.n278 72.8958
R2957 VDD.n1586 VDD.n1319 72.8958
R2958 VDD.n1454 VDD.n1319 72.8958
R2959 VDD.n1579 VDD.n1319 72.8958
R2960 VDD.n1573 VDD.n1319 72.8958
R2961 VDD.n1571 VDD.n1319 72.8958
R2962 VDD.n1565 VDD.n1319 72.8958
R2963 VDD.n1563 VDD.n1319 72.8958
R2964 VDD.n1557 VDD.n1319 72.8958
R2965 VDD.n1555 VDD.n1319 72.8958
R2966 VDD.n1549 VDD.n1319 72.8958
R2967 VDD.n1858 VDD.n488 72.8958
R2968 VDD.n1858 VDD.n489 72.8958
R2969 VDD.n1858 VDD.n490 72.8958
R2970 VDD.n1858 VDD.n491 72.8958
R2971 VDD.n1858 VDD.n492 72.8958
R2972 VDD.n1858 VDD.n493 72.8958
R2973 VDD.n1858 VDD.n494 72.8958
R2974 VDD.n1858 VDD.n495 72.8958
R2975 VDD.n1858 VDD.n496 72.8958
R2976 VDD.n1858 VDD.n497 72.8958
R2977 VDD.n2128 VDD.n1859 72.8958
R2978 VDD.n1865 VDD.n1859 72.8958
R2979 VDD.n2121 VDD.n1859 72.8958
R2980 VDD.n2115 VDD.n1859 72.8958
R2981 VDD.n2113 VDD.n1859 72.8958
R2982 VDD.n2107 VDD.n1859 72.8958
R2983 VDD.n2105 VDD.n1859 72.8958
R2984 VDD.n2099 VDD.n1859 72.8958
R2985 VDD.n2097 VDD.n1859 72.8958
R2986 VDD.n2091 VDD.n1859 72.8958
R2987 VDD.n2400 VDD.n288 72.8958
R2988 VDD.n2400 VDD.n289 72.8958
R2989 VDD.n2400 VDD.n290 72.8958
R2990 VDD.n2400 VDD.n291 72.8958
R2991 VDD.n2400 VDD.n292 72.8958
R2992 VDD.n2400 VDD.n293 72.8958
R2993 VDD.n2400 VDD.n294 72.8958
R2994 VDD.n2400 VDD.n295 72.8958
R2995 VDD.n2400 VDD.n296 72.8958
R2996 VDD.n2400 VDD.n297 72.8958
R2997 VDD.n2466 VDD.n2401 66.2847
R2998 VDD.n2405 VDD.n2401 66.2847
R2999 VDD.n2459 VDD.n2401 66.2847
R3000 VDD.n2452 VDD.n2401 66.2847
R3001 VDD.n2450 VDD.n2401 66.2847
R3002 VDD.n2444 VDD.n2401 66.2847
R3003 VDD.n2442 VDD.n2401 66.2847
R3004 VDD.n2428 VDD.n2401 66.2847
R3005 VDD.n2431 VDD.n2401 66.2847
R3006 VDD.n2710 VDD.n130 66.2847
R3007 VDD.n2710 VDD.n131 66.2847
R3008 VDD.n2710 VDD.n132 66.2847
R3009 VDD.n2710 VDD.n133 66.2847
R3010 VDD.n2710 VDD.n134 66.2847
R3011 VDD.n2710 VDD.n135 66.2847
R3012 VDD.n2710 VDD.n136 66.2847
R3013 VDD.n2710 VDD.n137 66.2847
R3014 VDD.n2710 VDD.n138 66.2847
R3015 VDD.n1318 VDD.n687 66.2847
R3016 VDD.n1318 VDD.n686 66.2847
R3017 VDD.n1318 VDD.n685 66.2847
R3018 VDD.n1318 VDD.n684 66.2847
R3019 VDD.n1318 VDD.n683 66.2847
R3020 VDD.n1318 VDD.n682 66.2847
R3021 VDD.n1318 VDD.n681 66.2847
R3022 VDD.n1318 VDD.n680 66.2847
R3023 VDD.n1318 VDD.n679 66.2847
R3024 VDD.n921 VDD.n893 66.2847
R3025 VDD.n929 VDD.n893 66.2847
R3026 VDD.n931 VDD.n893 66.2847
R3027 VDD.n939 VDD.n893 66.2847
R3028 VDD.n941 VDD.n893 66.2847
R3029 VDD.n950 VDD.n893 66.2847
R3030 VDD.n953 VDD.n893 66.2847
R3031 VDD.n904 VDD.n893 66.2847
R3032 VDD.n896 VDD.n893 66.2847
R3033 VDD.n1875 VDD.n1874 53.5278
R3034 VDD.n302 VDD.n301 53.5278
R3035 VDD.n1464 VDD.n1463 53.5278
R3036 VDD.n502 VDD.n501 53.5278
R3037 VDD.n1936 VDD.n1935 53.5278
R3038 VDD.n319 VDD.n318 53.5278
R3039 VDD.n1325 VDD.n1324 53.5278
R3040 VDD.n519 VDD.n518 53.5278
R3041 VDD.n2701 VDD.n138 52.4337
R3042 VDD.n2699 VDD.n137 52.4337
R3043 VDD.n2695 VDD.n136 52.4337
R3044 VDD.n2688 VDD.n135 52.4337
R3045 VDD.n2684 VDD.n134 52.4337
R3046 VDD.n2680 VDD.n133 52.4337
R3047 VDD.n2676 VDD.n132 52.4337
R3048 VDD.n2672 VDD.n131 52.4337
R3049 VDD.n156 VDD.n130 52.4337
R3050 VDD.n2466 VDD.n2402 52.4337
R3051 VDD.n2464 VDD.n2405 52.4337
R3052 VDD.n2460 VDD.n2459 52.4337
R3053 VDD.n2452 VDD.n2410 52.4337
R3054 VDD.n2451 VDD.n2450 52.4337
R3055 VDD.n2444 VDD.n2418 52.4337
R3056 VDD.n2443 VDD.n2442 52.4337
R3057 VDD.n2428 VDD.n2424 52.4337
R3058 VDD.n2432 VDD.n2431 52.4337
R3059 VDD.n2467 VDD.n2466 52.4337
R3060 VDD.n2461 VDD.n2405 52.4337
R3061 VDD.n2459 VDD.n2458 52.4337
R3062 VDD.n2453 VDD.n2452 52.4337
R3063 VDD.n2450 VDD.n2449 52.4337
R3064 VDD.n2445 VDD.n2444 52.4337
R3065 VDD.n2442 VDD.n2441 52.4337
R3066 VDD.n2429 VDD.n2428 52.4337
R3067 VDD.n2431 VDD.n275 52.4337
R3068 VDD.n2671 VDD.n130 52.4337
R3069 VDD.n2675 VDD.n131 52.4337
R3070 VDD.n2679 VDD.n132 52.4337
R3071 VDD.n2683 VDD.n133 52.4337
R3072 VDD.n2687 VDD.n134 52.4337
R3073 VDD.n2694 VDD.n135 52.4337
R3074 VDD.n2698 VDD.n136 52.4337
R3075 VDD.n2702 VDD.n137 52.4337
R3076 VDD.n139 VDD.n138 52.4337
R3077 VDD.n1253 VDD.n679 52.4337
R3078 VDD.n1255 VDD.n680 52.4337
R3079 VDD.n1259 VDD.n681 52.4337
R3080 VDD.n1261 VDD.n682 52.4337
R3081 VDD.n1268 VDD.n683 52.4337
R3082 VDD.n1270 VDD.n684 52.4337
R3083 VDD.n1274 VDD.n685 52.4337
R3084 VDD.n1276 VDD.n686 52.4337
R3085 VDD.n1279 VDD.n687 52.4337
R3086 VDD.n688 VDD.n687 52.4337
R3087 VDD.n1278 VDD.n686 52.4337
R3088 VDD.n1275 VDD.n685 52.4337
R3089 VDD.n1273 VDD.n684 52.4337
R3090 VDD.n1269 VDD.n683 52.4337
R3091 VDD.n1267 VDD.n682 52.4337
R3092 VDD.n1260 VDD.n681 52.4337
R3093 VDD.n1258 VDD.n680 52.4337
R3094 VDD.n1254 VDD.n679 52.4337
R3095 VDD.n921 VDD.n892 52.4337
R3096 VDD.n929 VDD.n928 52.4337
R3097 VDD.n932 VDD.n931 52.4337
R3098 VDD.n939 VDD.n938 52.4337
R3099 VDD.n942 VDD.n941 52.4337
R3100 VDD.n950 VDD.n949 52.4337
R3101 VDD.n953 VDD.n952 52.4337
R3102 VDD.n905 VDD.n904 52.4337
R3103 VDD.n897 VDD.n896 52.4337
R3104 VDD.n922 VDD.n921 52.4337
R3105 VDD.n930 VDD.n929 52.4337
R3106 VDD.n931 VDD.n911 52.4337
R3107 VDD.n940 VDD.n939 52.4337
R3108 VDD.n941 VDD.n907 52.4337
R3109 VDD.n951 VDD.n950 52.4337
R3110 VDD.n954 VDD.n953 52.4337
R3111 VDD.n904 VDD.n901 52.4337
R3112 VDD.n896 VDD.n894 52.4337
R3113 VDD.n1319 VDD.t89 43.6826
R3114 VDD.t105 VDD.n2400 43.6826
R3115 VDD.n1118 VDD.n1116 39.9002
R3116 VDD.n1109 VDD.n1107 39.9002
R3117 VDD.n2395 VDD.n297 39.2114
R3118 VDD.n2391 VDD.n296 39.2114
R3119 VDD.n2387 VDD.n295 39.2114
R3120 VDD.n2383 VDD.n294 39.2114
R3121 VDD.n2379 VDD.n293 39.2114
R3122 VDD.n2375 VDD.n292 39.2114
R3123 VDD.n2371 VDD.n291 39.2114
R3124 VDD.n2367 VDD.n290 39.2114
R3125 VDD.n2362 VDD.n289 39.2114
R3126 VDD.n2358 VDD.n288 39.2114
R3127 VDD.n2128 VDD.n1863 39.2114
R3128 VDD.n2126 VDD.n1865 39.2114
R3129 VDD.n2122 VDD.n2121 39.2114
R3130 VDD.n2115 VDD.n1867 39.2114
R3131 VDD.n2114 VDD.n2113 39.2114
R3132 VDD.n2107 VDD.n1869 39.2114
R3133 VDD.n2106 VDD.n2105 39.2114
R3134 VDD.n2099 VDD.n1871 39.2114
R3135 VDD.n2098 VDD.n2097 39.2114
R3136 VDD.n2091 VDD.n1873 39.2114
R3137 VDD.n1853 VDD.n497 39.2114
R3138 VDD.n1849 VDD.n496 39.2114
R3139 VDD.n1845 VDD.n495 39.2114
R3140 VDD.n1841 VDD.n494 39.2114
R3141 VDD.n1837 VDD.n493 39.2114
R3142 VDD.n1833 VDD.n492 39.2114
R3143 VDD.n1829 VDD.n491 39.2114
R3144 VDD.n1825 VDD.n490 39.2114
R3145 VDD.n1820 VDD.n489 39.2114
R3146 VDD.n1816 VDD.n488 39.2114
R3147 VDD.n1586 VDD.n1452 39.2114
R3148 VDD.n1584 VDD.n1454 39.2114
R3149 VDD.n1580 VDD.n1579 39.2114
R3150 VDD.n1573 VDD.n1456 39.2114
R3151 VDD.n1572 VDD.n1571 39.2114
R3152 VDD.n1565 VDD.n1458 39.2114
R3153 VDD.n1564 VDD.n1563 39.2114
R3154 VDD.n1557 VDD.n1460 39.2114
R3155 VDD.n1556 VDD.n1555 39.2114
R3156 VDD.n1549 VDD.n1462 39.2114
R3157 VDD.n2338 VDD.n278 39.2114
R3158 VDD.n2334 VDD.n279 39.2114
R3159 VDD.n2330 VDD.n280 39.2114
R3160 VDD.n2326 VDD.n281 39.2114
R3161 VDD.n2322 VDD.n282 39.2114
R3162 VDD.n2318 VDD.n283 39.2114
R3163 VDD.n2314 VDD.n284 39.2114
R3164 VDD.n2310 VDD.n285 39.2114
R3165 VDD.n2305 VDD.n286 39.2114
R3166 VDD.n2301 VDD.n287 39.2114
R3167 VDD.n1944 VDD.n475 39.2114
R3168 VDD.n1949 VDD.n1948 39.2114
R3169 VDD.n1952 VDD.n1951 39.2114
R3170 VDD.n1957 VDD.n1956 39.2114
R3171 VDD.n1960 VDD.n1959 39.2114
R3172 VDD.n1965 VDD.n1964 39.2114
R3173 VDD.n1968 VDD.n1967 39.2114
R3174 VDD.n1973 VDD.n1972 39.2114
R3175 VDD.n1976 VDD.n1975 39.2114
R3176 VDD.n1982 VDD.n1981 39.2114
R3177 VDD.n1796 VDD.n478 39.2114
R3178 VDD.n1792 VDD.n479 39.2114
R3179 VDD.n1788 VDD.n480 39.2114
R3180 VDD.n1784 VDD.n481 39.2114
R3181 VDD.n1780 VDD.n482 39.2114
R3182 VDD.n1776 VDD.n483 39.2114
R3183 VDD.n1772 VDD.n484 39.2114
R3184 VDD.n1768 VDD.n485 39.2114
R3185 VDD.n1763 VDD.n486 39.2114
R3186 VDD.n1759 VDD.n487 39.2114
R3187 VDD.n1336 VDD.n677 39.2114
R3188 VDD.n1339 VDD.n1338 39.2114
R3189 VDD.n1344 VDD.n1343 39.2114
R3190 VDD.n1347 VDD.n1346 39.2114
R3191 VDD.n1352 VDD.n1351 39.2114
R3192 VDD.n1355 VDD.n1354 39.2114
R3193 VDD.n1360 VDD.n1359 39.2114
R3194 VDD.n1363 VDD.n1362 39.2114
R3195 VDD.n1368 VDD.n1367 39.2114
R3196 VDD.n1371 VDD.n1370 39.2114
R3197 VDD.n1337 VDD.n1336 39.2114
R3198 VDD.n1338 VDD.n1334 39.2114
R3199 VDD.n1345 VDD.n1344 39.2114
R3200 VDD.n1346 VDD.n1332 39.2114
R3201 VDD.n1353 VDD.n1352 39.2114
R3202 VDD.n1354 VDD.n1330 39.2114
R3203 VDD.n1361 VDD.n1360 39.2114
R3204 VDD.n1362 VDD.n1328 39.2114
R3205 VDD.n1369 VDD.n1368 39.2114
R3206 VDD.n1372 VDD.n1371 39.2114
R3207 VDD.n1762 VDD.n487 39.2114
R3208 VDD.n1767 VDD.n486 39.2114
R3209 VDD.n1771 VDD.n485 39.2114
R3210 VDD.n1775 VDD.n484 39.2114
R3211 VDD.n1779 VDD.n483 39.2114
R3212 VDD.n1783 VDD.n482 39.2114
R3213 VDD.n1787 VDD.n481 39.2114
R3214 VDD.n1791 VDD.n480 39.2114
R3215 VDD.n1795 VDD.n479 39.2114
R3216 VDD.n1798 VDD.n478 39.2114
R3217 VDD.n1945 VDD.n1944 39.2114
R3218 VDD.n1950 VDD.n1949 39.2114
R3219 VDD.n1951 VDD.n1942 39.2114
R3220 VDD.n1958 VDD.n1957 39.2114
R3221 VDD.n1959 VDD.n1940 39.2114
R3222 VDD.n1966 VDD.n1965 39.2114
R3223 VDD.n1967 VDD.n1938 39.2114
R3224 VDD.n1974 VDD.n1973 39.2114
R3225 VDD.n1975 VDD.n1934 39.2114
R3226 VDD.n1983 VDD.n1982 39.2114
R3227 VDD.n2304 VDD.n287 39.2114
R3228 VDD.n2309 VDD.n286 39.2114
R3229 VDD.n2313 VDD.n285 39.2114
R3230 VDD.n2317 VDD.n284 39.2114
R3231 VDD.n2321 VDD.n283 39.2114
R3232 VDD.n2325 VDD.n282 39.2114
R3233 VDD.n2329 VDD.n281 39.2114
R3234 VDD.n2333 VDD.n280 39.2114
R3235 VDD.n2337 VDD.n279 39.2114
R3236 VDD.n2340 VDD.n278 39.2114
R3237 VDD.n1587 VDD.n1586 39.2114
R3238 VDD.n1581 VDD.n1454 39.2114
R3239 VDD.n1579 VDD.n1578 39.2114
R3240 VDD.n1574 VDD.n1573 39.2114
R3241 VDD.n1571 VDD.n1570 39.2114
R3242 VDD.n1566 VDD.n1565 39.2114
R3243 VDD.n1563 VDD.n1562 39.2114
R3244 VDD.n1558 VDD.n1557 39.2114
R3245 VDD.n1555 VDD.n1554 39.2114
R3246 VDD.n1550 VDD.n1549 39.2114
R3247 VDD.n1819 VDD.n488 39.2114
R3248 VDD.n1824 VDD.n489 39.2114
R3249 VDD.n1828 VDD.n490 39.2114
R3250 VDD.n1832 VDD.n491 39.2114
R3251 VDD.n1836 VDD.n492 39.2114
R3252 VDD.n1840 VDD.n493 39.2114
R3253 VDD.n1844 VDD.n494 39.2114
R3254 VDD.n1848 VDD.n495 39.2114
R3255 VDD.n1852 VDD.n496 39.2114
R3256 VDD.n499 VDD.n497 39.2114
R3257 VDD.n2129 VDD.n2128 39.2114
R3258 VDD.n2123 VDD.n1865 39.2114
R3259 VDD.n2121 VDD.n2120 39.2114
R3260 VDD.n2116 VDD.n2115 39.2114
R3261 VDD.n2113 VDD.n2112 39.2114
R3262 VDD.n2108 VDD.n2107 39.2114
R3263 VDD.n2105 VDD.n2104 39.2114
R3264 VDD.n2100 VDD.n2099 39.2114
R3265 VDD.n2097 VDD.n2096 39.2114
R3266 VDD.n2092 VDD.n2091 39.2114
R3267 VDD.n2361 VDD.n288 39.2114
R3268 VDD.n2366 VDD.n289 39.2114
R3269 VDD.n2370 VDD.n290 39.2114
R3270 VDD.n2374 VDD.n291 39.2114
R3271 VDD.n2378 VDD.n292 39.2114
R3272 VDD.n2382 VDD.n293 39.2114
R3273 VDD.n2386 VDD.n294 39.2114
R3274 VDD.n2390 VDD.n295 39.2114
R3275 VDD.n2394 VDD.n296 39.2114
R3276 VDD.n299 VDD.n297 39.2114
R3277 VDD.n960 VDD.n899 37.2369
R3278 VDD.n915 VDD.n914 37.2369
R3279 VDD.n2455 VDD.n2415 37.2369
R3280 VDD.n2435 VDD.n2434 37.2369
R3281 VDD.n2670 VDD.n159 37.2369
R3282 VDD.n2692 VDD.n2691 37.2369
R3283 VDD.n1266 VDD.n1265 37.2369
R3284 VDD.n692 VDD.n691 37.2369
R3285 VDD.n33 VDD.n32 37.2278
R3286 VDD.n24 VDD.n23 37.2278
R3287 VDD.n2132 VDD.n2131 32.6249
R3288 VDD.n2398 VDD.n300 32.6249
R3289 VDD.n2359 VDD.n303 32.6249
R3290 VDD.n2093 VDD.n2090 32.6249
R3291 VDD.n1856 VDD.n500 32.6249
R3292 VDD.n1817 VDD.n503 32.6249
R3293 VDD.n1551 VDD.n1548 32.6249
R3294 VDD.n1590 VDD.n1589 32.6249
R3295 VDD.n2344 VDD.n2342 32.6249
R3296 VDD.n2302 VDD.n2299 32.6249
R3297 VDD.n1986 VDD.n1985 32.6249
R3298 VDD.n2136 VDD.n474 32.6249
R3299 VDD.n1802 VDD.n1800 32.6249
R3300 VDD.n1760 VDD.n1757 32.6249
R3301 VDD.n1450 VDD.n1374 32.6249
R3302 VDD.n1594 VDD.n676 32.6249
R3303 VDD.n1876 VDD.n1875 30.449
R3304 VDD.n2364 VDD.n302 30.449
R3305 VDD.n1465 VDD.n1464 30.449
R3306 VDD.n1822 VDD.n502 30.449
R3307 VDD.n1979 VDD.n1936 30.449
R3308 VDD.n2307 VDD.n319 30.449
R3309 VDD.n1326 VDD.n1325 30.449
R3310 VDD.n1765 VDD.n519 30.449
R3311 VDD.n966 VDD.n893 27.5168
R3312 VDD.n1318 VDD.n678 27.5168
R3313 VDD.n2474 VDD.n2401 27.5168
R3314 VDD.n2711 VDD.n2710 27.5168
R3315 VDD.n1592 VDD.n1319 23.0454
R3316 VDD.n1858 VDD.n476 23.0454
R3317 VDD.n2134 VDD.n1859 23.0454
R3318 VDD.n2400 VDD.n276 23.0454
R3319 VDD.n943 VDD.n910 19.3944
R3320 VDD.n943 VDD.n908 19.3944
R3321 VDD.n948 VDD.n908 19.3944
R3322 VDD.n948 VDD.n906 19.3944
R3323 VDD.n906 VDD.n903 19.3944
R3324 VDD.n955 VDD.n903 19.3944
R3325 VDD.n955 VDD.n900 19.3944
R3326 VDD.n959 VDD.n900 19.3944
R3327 VDD.n923 VDD.n920 19.3944
R3328 VDD.n923 VDD.n919 19.3944
R3329 VDD.n927 VDD.n919 19.3944
R3330 VDD.n927 VDD.n917 19.3944
R3331 VDD.n933 VDD.n917 19.3944
R3332 VDD.n933 VDD.n912 19.3944
R3333 VDD.n937 VDD.n912 19.3944
R3334 VDD.n964 VDD.n886 19.3944
R3335 VDD.n976 VDD.n886 19.3944
R3336 VDD.n976 VDD.n884 19.3944
R3337 VDD.n980 VDD.n884 19.3944
R3338 VDD.n980 VDD.n874 19.3944
R3339 VDD.n992 VDD.n874 19.3944
R3340 VDD.n992 VDD.n872 19.3944
R3341 VDD.n996 VDD.n872 19.3944
R3342 VDD.n996 VDD.n862 19.3944
R3343 VDD.n1008 VDD.n862 19.3944
R3344 VDD.n1008 VDD.n860 19.3944
R3345 VDD.n1012 VDD.n860 19.3944
R3346 VDD.n1012 VDD.n850 19.3944
R3347 VDD.n1024 VDD.n850 19.3944
R3348 VDD.n1024 VDD.n848 19.3944
R3349 VDD.n1028 VDD.n848 19.3944
R3350 VDD.n1028 VDD.n838 19.3944
R3351 VDD.n1040 VDD.n838 19.3944
R3352 VDD.n1040 VDD.n836 19.3944
R3353 VDD.n1044 VDD.n836 19.3944
R3354 VDD.n1044 VDD.n827 19.3944
R3355 VDD.n1057 VDD.n827 19.3944
R3356 VDD.n1057 VDD.n825 19.3944
R3357 VDD.n1061 VDD.n825 19.3944
R3358 VDD.n1061 VDD.n815 19.3944
R3359 VDD.n1073 VDD.n815 19.3944
R3360 VDD.n1073 VDD.n813 19.3944
R3361 VDD.n1077 VDD.n813 19.3944
R3362 VDD.n1077 VDD.n803 19.3944
R3363 VDD.n1089 VDD.n803 19.3944
R3364 VDD.n1089 VDD.n801 19.3944
R3365 VDD.n1093 VDD.n801 19.3944
R3366 VDD.n1093 VDD.n792 19.3944
R3367 VDD.n1127 VDD.n792 19.3944
R3368 VDD.n1127 VDD.n790 19.3944
R3369 VDD.n1131 VDD.n790 19.3944
R3370 VDD.n1131 VDD.n780 19.3944
R3371 VDD.n1143 VDD.n780 19.3944
R3372 VDD.n1143 VDD.n778 19.3944
R3373 VDD.n1147 VDD.n778 19.3944
R3374 VDD.n1147 VDD.n768 19.3944
R3375 VDD.n1159 VDD.n768 19.3944
R3376 VDD.n1159 VDD.n766 19.3944
R3377 VDD.n1163 VDD.n766 19.3944
R3378 VDD.n1163 VDD.n757 19.3944
R3379 VDD.n1176 VDD.n757 19.3944
R3380 VDD.n1176 VDD.n755 19.3944
R3381 VDD.n1180 VDD.n755 19.3944
R3382 VDD.n1180 VDD.n745 19.3944
R3383 VDD.n1192 VDD.n745 19.3944
R3384 VDD.n1192 VDD.n743 19.3944
R3385 VDD.n1196 VDD.n743 19.3944
R3386 VDD.n1196 VDD.n733 19.3944
R3387 VDD.n1208 VDD.n733 19.3944
R3388 VDD.n1208 VDD.n731 19.3944
R3389 VDD.n1212 VDD.n731 19.3944
R3390 VDD.n1212 VDD.n721 19.3944
R3391 VDD.n1224 VDD.n721 19.3944
R3392 VDD.n1224 VDD.n719 19.3944
R3393 VDD.n1228 VDD.n719 19.3944
R3394 VDD.n1228 VDD.n709 19.3944
R3395 VDD.n1240 VDD.n709 19.3944
R3396 VDD.n1240 VDD.n707 19.3944
R3397 VDD.n1245 VDD.n707 19.3944
R3398 VDD.n1245 VDD.n695 19.3944
R3399 VDD.n1312 VDD.n695 19.3944
R3400 VDD.n1313 VDD.n1312 19.3944
R3401 VDD.n2469 VDD.n2468 19.3944
R3402 VDD.n2468 VDD.n2404 19.3944
R3403 VDD.n2463 VDD.n2404 19.3944
R3404 VDD.n2463 VDD.n2462 19.3944
R3405 VDD.n2462 VDD.n2409 19.3944
R3406 VDD.n2457 VDD.n2409 19.3944
R3407 VDD.n2457 VDD.n2456 19.3944
R3408 VDD.n2454 VDD.n2417 19.3944
R3409 VDD.n2448 VDD.n2417 19.3944
R3410 VDD.n2448 VDD.n2447 19.3944
R3411 VDD.n2447 VDD.n2446 19.3944
R3412 VDD.n2446 VDD.n2423 19.3944
R3413 VDD.n2440 VDD.n2423 19.3944
R3414 VDD.n2440 VDD.n2439 19.3944
R3415 VDD.n2439 VDD.n2438 19.3944
R3416 VDD.n2476 VDD.n273 19.3944
R3417 VDD.n2480 VDD.n273 19.3944
R3418 VDD.n2480 VDD.n263 19.3944
R3419 VDD.n2492 VDD.n263 19.3944
R3420 VDD.n2492 VDD.n261 19.3944
R3421 VDD.n2496 VDD.n261 19.3944
R3422 VDD.n2496 VDD.n251 19.3944
R3423 VDD.n2508 VDD.n251 19.3944
R3424 VDD.n2508 VDD.n249 19.3944
R3425 VDD.n2512 VDD.n249 19.3944
R3426 VDD.n2512 VDD.n239 19.3944
R3427 VDD.n2524 VDD.n239 19.3944
R3428 VDD.n2524 VDD.n237 19.3944
R3429 VDD.n2528 VDD.n237 19.3944
R3430 VDD.n2528 VDD.n227 19.3944
R3431 VDD.n2540 VDD.n227 19.3944
R3432 VDD.n2540 VDD.n225 19.3944
R3433 VDD.n2544 VDD.n225 19.3944
R3434 VDD.n2544 VDD.n214 19.3944
R3435 VDD.n2556 VDD.n214 19.3944
R3436 VDD.n2556 VDD.n212 19.3944
R3437 VDD.n2560 VDD.n212 19.3944
R3438 VDD.n2560 VDD.n203 19.3944
R3439 VDD.n2572 VDD.n203 19.3944
R3440 VDD.n2572 VDD.n201 19.3944
R3441 VDD.n2576 VDD.n201 19.3944
R3442 VDD.n2576 VDD.n191 19.3944
R3443 VDD.n2588 VDD.n191 19.3944
R3444 VDD.n2588 VDD.n189 19.3944
R3445 VDD.n2595 VDD.n189 19.3944
R3446 VDD.n2595 VDD.n2594 19.3944
R3447 VDD.n2594 VDD.n177 19.3944
R3448 VDD.n2608 VDD.n177 19.3944
R3449 VDD.n2609 VDD.n2608 19.3944
R3450 VDD.n2610 VDD.n2609 19.3944
R3451 VDD.n2610 VDD.n175 19.3944
R3452 VDD.n2615 VDD.n175 19.3944
R3453 VDD.n2616 VDD.n2615 19.3944
R3454 VDD.n2617 VDD.n2616 19.3944
R3455 VDD.n2617 VDD.n173 19.3944
R3456 VDD.n2622 VDD.n173 19.3944
R3457 VDD.n2623 VDD.n2622 19.3944
R3458 VDD.n2624 VDD.n2623 19.3944
R3459 VDD.n2624 VDD.n171 19.3944
R3460 VDD.n2629 VDD.n171 19.3944
R3461 VDD.n2630 VDD.n2629 19.3944
R3462 VDD.n2631 VDD.n2630 19.3944
R3463 VDD.n2631 VDD.n169 19.3944
R3464 VDD.n2636 VDD.n169 19.3944
R3465 VDD.n2637 VDD.n2636 19.3944
R3466 VDD.n2638 VDD.n2637 19.3944
R3467 VDD.n2638 VDD.n167 19.3944
R3468 VDD.n2643 VDD.n167 19.3944
R3469 VDD.n2644 VDD.n2643 19.3944
R3470 VDD.n2645 VDD.n2644 19.3944
R3471 VDD.n2645 VDD.n165 19.3944
R3472 VDD.n2650 VDD.n165 19.3944
R3473 VDD.n2651 VDD.n2650 19.3944
R3474 VDD.n2652 VDD.n2651 19.3944
R3475 VDD.n2652 VDD.n163 19.3944
R3476 VDD.n2657 VDD.n163 19.3944
R3477 VDD.n2658 VDD.n2657 19.3944
R3478 VDD.n2659 VDD.n2658 19.3944
R3479 VDD.n2659 VDD.n161 19.3944
R3480 VDD.n2664 VDD.n161 19.3944
R3481 VDD.n2665 VDD.n2664 19.3944
R3482 VDD.n2666 VDD.n2665 19.3944
R3483 VDD.n2689 VDD.n2686 19.3944
R3484 VDD.n2686 VDD.n2685 19.3944
R3485 VDD.n2685 VDD.n2682 19.3944
R3486 VDD.n2682 VDD.n2681 19.3944
R3487 VDD.n2681 VDD.n2678 19.3944
R3488 VDD.n2678 VDD.n2677 19.3944
R3489 VDD.n2677 VDD.n2674 19.3944
R3490 VDD.n2674 VDD.n2673 19.3944
R3491 VDD.n2708 VDD.n2707 19.3944
R3492 VDD.n2707 VDD.n142 19.3944
R3493 VDD.n2703 VDD.n142 19.3944
R3494 VDD.n2703 VDD.n2700 19.3944
R3495 VDD.n2700 VDD.n2697 19.3944
R3496 VDD.n2697 VDD.n2696 19.3944
R3497 VDD.n2696 VDD.n2693 19.3944
R3498 VDD.n2472 VDD.n269 19.3944
R3499 VDD.n2484 VDD.n269 19.3944
R3500 VDD.n2484 VDD.n267 19.3944
R3501 VDD.n2488 VDD.n267 19.3944
R3502 VDD.n2488 VDD.n257 19.3944
R3503 VDD.n2500 VDD.n257 19.3944
R3504 VDD.n2500 VDD.n255 19.3944
R3505 VDD.n2504 VDD.n255 19.3944
R3506 VDD.n2504 VDD.n245 19.3944
R3507 VDD.n2516 VDD.n245 19.3944
R3508 VDD.n2516 VDD.n243 19.3944
R3509 VDD.n2520 VDD.n243 19.3944
R3510 VDD.n2520 VDD.n233 19.3944
R3511 VDD.n2532 VDD.n233 19.3944
R3512 VDD.n2532 VDD.n231 19.3944
R3513 VDD.n2536 VDD.n231 19.3944
R3514 VDD.n2536 VDD.n221 19.3944
R3515 VDD.n2548 VDD.n221 19.3944
R3516 VDD.n2548 VDD.n219 19.3944
R3517 VDD.n2552 VDD.n219 19.3944
R3518 VDD.n2552 VDD.n209 19.3944
R3519 VDD.n2564 VDD.n209 19.3944
R3520 VDD.n2564 VDD.n207 19.3944
R3521 VDD.n2568 VDD.n207 19.3944
R3522 VDD.n2568 VDD.n197 19.3944
R3523 VDD.n2580 VDD.n197 19.3944
R3524 VDD.n2580 VDD.n195 19.3944
R3525 VDD.n2584 VDD.n195 19.3944
R3526 VDD.n2584 VDD.n184 19.3944
R3527 VDD.n2599 VDD.n184 19.3944
R3528 VDD.n2599 VDD.n182 19.3944
R3529 VDD.n2603 VDD.n182 19.3944
R3530 VDD.n2603 VDD.n37 19.3944
R3531 VDD.n2778 VDD.n37 19.3944
R3532 VDD.n2778 VDD.n38 19.3944
R3533 VDD.n2772 VDD.n38 19.3944
R3534 VDD.n2772 VDD.n2771 19.3944
R3535 VDD.n2771 VDD.n2770 19.3944
R3536 VDD.n2770 VDD.n49 19.3944
R3537 VDD.n2764 VDD.n49 19.3944
R3538 VDD.n2764 VDD.n2763 19.3944
R3539 VDD.n2763 VDD.n2762 19.3944
R3540 VDD.n2762 VDD.n60 19.3944
R3541 VDD.n2756 VDD.n60 19.3944
R3542 VDD.n2756 VDD.n2755 19.3944
R3543 VDD.n2755 VDD.n2754 19.3944
R3544 VDD.n2754 VDD.n71 19.3944
R3545 VDD.n2748 VDD.n71 19.3944
R3546 VDD.n2748 VDD.n2747 19.3944
R3547 VDD.n2747 VDD.n2746 19.3944
R3548 VDD.n2746 VDD.n82 19.3944
R3549 VDD.n2740 VDD.n82 19.3944
R3550 VDD.n2740 VDD.n2739 19.3944
R3551 VDD.n2739 VDD.n2738 19.3944
R3552 VDD.n2738 VDD.n93 19.3944
R3553 VDD.n2732 VDD.n93 19.3944
R3554 VDD.n2732 VDD.n2731 19.3944
R3555 VDD.n2731 VDD.n2730 19.3944
R3556 VDD.n2730 VDD.n104 19.3944
R3557 VDD.n2724 VDD.n104 19.3944
R3558 VDD.n2724 VDD.n2723 19.3944
R3559 VDD.n2723 VDD.n2722 19.3944
R3560 VDD.n2722 VDD.n114 19.3944
R3561 VDD.n2716 VDD.n114 19.3944
R3562 VDD.n2716 VDD.n2715 19.3944
R3563 VDD.n2715 VDD.n2714 19.3944
R3564 VDD.n2714 VDD.n126 19.3944
R3565 VDD.n1304 VDD.n1303 19.3944
R3566 VDD.n1303 VDD.n1302 19.3944
R3567 VDD.n1302 VDD.n1256 19.3944
R3568 VDD.n1298 VDD.n1256 19.3944
R3569 VDD.n1298 VDD.n1297 19.3944
R3570 VDD.n1297 VDD.n1296 19.3944
R3571 VDD.n1296 VDD.n1262 19.3944
R3572 VDD.n1292 VDD.n1291 19.3944
R3573 VDD.n1291 VDD.n1290 19.3944
R3574 VDD.n1290 VDD.n1271 19.3944
R3575 VDD.n1286 VDD.n1271 19.3944
R3576 VDD.n1286 VDD.n1285 19.3944
R3577 VDD.n1285 VDD.n1284 19.3944
R3578 VDD.n1284 VDD.n1277 19.3944
R3579 VDD.n1280 VDD.n1277 19.3944
R3580 VDD.n968 VDD.n890 19.3944
R3581 VDD.n972 VDD.n890 19.3944
R3582 VDD.n972 VDD.n880 19.3944
R3583 VDD.n984 VDD.n880 19.3944
R3584 VDD.n984 VDD.n878 19.3944
R3585 VDD.n988 VDD.n878 19.3944
R3586 VDD.n988 VDD.n868 19.3944
R3587 VDD.n1000 VDD.n868 19.3944
R3588 VDD.n1000 VDD.n866 19.3944
R3589 VDD.n1004 VDD.n866 19.3944
R3590 VDD.n1004 VDD.n856 19.3944
R3591 VDD.n1016 VDD.n856 19.3944
R3592 VDD.n1016 VDD.n854 19.3944
R3593 VDD.n1020 VDD.n854 19.3944
R3594 VDD.n1020 VDD.n844 19.3944
R3595 VDD.n1032 VDD.n844 19.3944
R3596 VDD.n1032 VDD.n842 19.3944
R3597 VDD.n1036 VDD.n842 19.3944
R3598 VDD.n1036 VDD.n832 19.3944
R3599 VDD.n1049 VDD.n832 19.3944
R3600 VDD.n1049 VDD.n830 19.3944
R3601 VDD.n1053 VDD.n830 19.3944
R3602 VDD.n1053 VDD.n821 19.3944
R3603 VDD.n1065 VDD.n821 19.3944
R3604 VDD.n1065 VDD.n819 19.3944
R3605 VDD.n1069 VDD.n819 19.3944
R3606 VDD.n1069 VDD.n809 19.3944
R3607 VDD.n1081 VDD.n809 19.3944
R3608 VDD.n1081 VDD.n807 19.3944
R3609 VDD.n1085 VDD.n807 19.3944
R3610 VDD.n1085 VDD.n797 19.3944
R3611 VDD.n1098 VDD.n797 19.3944
R3612 VDD.n1098 VDD.n795 19.3944
R3613 VDD.n1123 VDD.n795 19.3944
R3614 VDD.n1123 VDD.n786 19.3944
R3615 VDD.n1135 VDD.n786 19.3944
R3616 VDD.n1135 VDD.n784 19.3944
R3617 VDD.n1139 VDD.n784 19.3944
R3618 VDD.n1139 VDD.n774 19.3944
R3619 VDD.n1151 VDD.n774 19.3944
R3620 VDD.n1151 VDD.n772 19.3944
R3621 VDD.n1155 VDD.n772 19.3944
R3622 VDD.n1155 VDD.n762 19.3944
R3623 VDD.n1168 VDD.n762 19.3944
R3624 VDD.n1168 VDD.n760 19.3944
R3625 VDD.n1172 VDD.n760 19.3944
R3626 VDD.n1172 VDD.n751 19.3944
R3627 VDD.n1184 VDD.n751 19.3944
R3628 VDD.n1184 VDD.n749 19.3944
R3629 VDD.n1188 VDD.n749 19.3944
R3630 VDD.n1188 VDD.n739 19.3944
R3631 VDD.n1200 VDD.n739 19.3944
R3632 VDD.n1200 VDD.n737 19.3944
R3633 VDD.n1204 VDD.n737 19.3944
R3634 VDD.n1204 VDD.n727 19.3944
R3635 VDD.n1216 VDD.n727 19.3944
R3636 VDD.n1216 VDD.n725 19.3944
R3637 VDD.n1220 VDD.n725 19.3944
R3638 VDD.n1220 VDD.n715 19.3944
R3639 VDD.n1232 VDD.n715 19.3944
R3640 VDD.n1232 VDD.n713 19.3944
R3641 VDD.n1236 VDD.n713 19.3944
R3642 VDD.n1236 VDD.n703 19.3944
R3643 VDD.n1249 VDD.n703 19.3944
R3644 VDD.n1249 VDD.n700 19.3944
R3645 VDD.n1308 VDD.n700 19.3944
R3646 VDD.n1308 VDD.n701 19.3944
R3647 VDD.n966 VDD.n888 17.1982
R3648 VDD.n974 VDD.n888 17.1982
R3649 VDD.n974 VDD.n882 17.1982
R3650 VDD.n982 VDD.n882 17.1982
R3651 VDD.n982 VDD.n876 17.1982
R3652 VDD.n990 VDD.n876 17.1982
R3653 VDD.n998 VDD.n870 17.1982
R3654 VDD.n998 VDD.n864 17.1982
R3655 VDD.n1006 VDD.n864 17.1982
R3656 VDD.n1006 VDD.n858 17.1982
R3657 VDD.n1014 VDD.n858 17.1982
R3658 VDD.n1014 VDD.n852 17.1982
R3659 VDD.n1022 VDD.n852 17.1982
R3660 VDD.n1022 VDD.n846 17.1982
R3661 VDD.n1030 VDD.n846 17.1982
R3662 VDD.n1030 VDD.n840 17.1982
R3663 VDD.n1038 VDD.n840 17.1982
R3664 VDD.n1038 VDD.n834 17.1982
R3665 VDD.n1047 VDD.n834 17.1982
R3666 VDD.n1047 VDD.n1046 17.1982
R3667 VDD.n1055 VDD.n823 17.1982
R3668 VDD.n1063 VDD.n823 17.1982
R3669 VDD.n1063 VDD.n817 17.1982
R3670 VDD.n1071 VDD.n817 17.1982
R3671 VDD.n1071 VDD.n811 17.1982
R3672 VDD.n1079 VDD.n811 17.1982
R3673 VDD.n1079 VDD.n805 17.1982
R3674 VDD.n1087 VDD.n805 17.1982
R3675 VDD.n1087 VDD.n799 17.1982
R3676 VDD.n1096 VDD.n799 17.1982
R3677 VDD.n1096 VDD.n1095 17.1982
R3678 VDD.n1125 VDD.n788 17.1982
R3679 VDD.n1133 VDD.n788 17.1982
R3680 VDD.n1133 VDD.n782 17.1982
R3681 VDD.n1141 VDD.n782 17.1982
R3682 VDD.n1141 VDD.n776 17.1982
R3683 VDD.n1149 VDD.n776 17.1982
R3684 VDD.n1149 VDD.n770 17.1982
R3685 VDD.n1157 VDD.n770 17.1982
R3686 VDD.n1157 VDD.n764 17.1982
R3687 VDD.n1166 VDD.n764 17.1982
R3688 VDD.n1166 VDD.n1165 17.1982
R3689 VDD.n1174 VDD.n753 17.1982
R3690 VDD.n1182 VDD.n753 17.1982
R3691 VDD.n1182 VDD.n747 17.1982
R3692 VDD.n1190 VDD.n747 17.1982
R3693 VDD.n1190 VDD.n741 17.1982
R3694 VDD.n1198 VDD.n741 17.1982
R3695 VDD.n1198 VDD.n735 17.1982
R3696 VDD.n1206 VDD.n735 17.1982
R3697 VDD.n1206 VDD.n729 17.1982
R3698 VDD.n1214 VDD.n729 17.1982
R3699 VDD.n1214 VDD.n723 17.1982
R3700 VDD.n1222 VDD.n723 17.1982
R3701 VDD.n1222 VDD.n717 17.1982
R3702 VDD.n1230 VDD.n717 17.1982
R3703 VDD.n1238 VDD.n711 17.1982
R3704 VDD.n1238 VDD.n705 17.1982
R3705 VDD.n1247 VDD.n705 17.1982
R3706 VDD.n1247 VDD.n697 17.1982
R3707 VDD.n1310 VDD.n697 17.1982
R3708 VDD.n1310 VDD.n678 17.1982
R3709 VDD.n2474 VDD.n271 17.1982
R3710 VDD.n2482 VDD.n271 17.1982
R3711 VDD.n2482 VDD.n265 17.1982
R3712 VDD.n2490 VDD.n265 17.1982
R3713 VDD.n2490 VDD.n259 17.1982
R3714 VDD.n2498 VDD.n259 17.1982
R3715 VDD.n2506 VDD.n253 17.1982
R3716 VDD.n2506 VDD.n247 17.1982
R3717 VDD.n2514 VDD.n247 17.1982
R3718 VDD.n2514 VDD.n241 17.1982
R3719 VDD.n2522 VDD.n241 17.1982
R3720 VDD.n2522 VDD.n235 17.1982
R3721 VDD.n2530 VDD.n235 17.1982
R3722 VDD.n2530 VDD.n229 17.1982
R3723 VDD.n2538 VDD.n229 17.1982
R3724 VDD.n2538 VDD.n223 17.1982
R3725 VDD.n2546 VDD.n223 17.1982
R3726 VDD.n2546 VDD.n216 17.1982
R3727 VDD.n2554 VDD.n216 17.1982
R3728 VDD.n2554 VDD.n217 17.1982
R3729 VDD.n2562 VDD.n205 17.1982
R3730 VDD.n2570 VDD.n205 17.1982
R3731 VDD.n2570 VDD.n199 17.1982
R3732 VDD.n2578 VDD.n199 17.1982
R3733 VDD.n2578 VDD.n193 17.1982
R3734 VDD.n2586 VDD.n193 17.1982
R3735 VDD.n2586 VDD.n186 17.1982
R3736 VDD.n2597 VDD.n186 17.1982
R3737 VDD.n2597 VDD.n180 17.1982
R3738 VDD.n2605 VDD.n180 17.1982
R3739 VDD.n2606 VDD.n2605 17.1982
R3740 VDD.n2776 VDD.n2775 17.1982
R3741 VDD.n2775 VDD.n2774 17.1982
R3742 VDD.n2774 VDD.n44 17.1982
R3743 VDD.n2768 VDD.n44 17.1982
R3744 VDD.n2768 VDD.n2767 17.1982
R3745 VDD.n2767 VDD.n2766 17.1982
R3746 VDD.n2766 VDD.n54 17.1982
R3747 VDD.n2760 VDD.n54 17.1982
R3748 VDD.n2760 VDD.n2759 17.1982
R3749 VDD.n2759 VDD.n2758 17.1982
R3750 VDD.n2758 VDD.n65 17.1982
R3751 VDD.n2752 VDD.n2751 17.1982
R3752 VDD.n2751 VDD.n2750 17.1982
R3753 VDD.n2750 VDD.n76 17.1982
R3754 VDD.n2744 VDD.n76 17.1982
R3755 VDD.n2744 VDD.n2743 17.1982
R3756 VDD.n2743 VDD.n2742 17.1982
R3757 VDD.n2742 VDD.n87 17.1982
R3758 VDD.n2736 VDD.n87 17.1982
R3759 VDD.n2736 VDD.n2735 17.1982
R3760 VDD.n2735 VDD.n2734 17.1982
R3761 VDD.n2734 VDD.n98 17.1982
R3762 VDD.n2728 VDD.n98 17.1982
R3763 VDD.n2728 VDD.n2727 17.1982
R3764 VDD.n2727 VDD.n2726 17.1982
R3765 VDD.n2720 VDD.n116 17.1982
R3766 VDD.n2720 VDD.n2719 17.1982
R3767 VDD.n2719 VDD.n2718 17.1982
R3768 VDD.n2718 VDD.n120 17.1982
R3769 VDD.n2712 VDD.n120 17.1982
R3770 VDD.n2712 VDD.n2711 17.1982
R3771 VDD.n25 VDD.t67 16.1721
R3772 VDD.n25 VDD.t58 16.1721
R3773 VDD.n16 VDD.t68 16.1721
R3774 VDD.n16 VDD.t61 16.1721
R3775 VDD.n1117 VDD.t71 16.1721
R3776 VDD.n1117 VDD.t65 16.1721
R3777 VDD.n1108 VDD.t72 16.1721
R3778 VDD.n1108 VDD.t69 16.1721
R3779 VDD.n1055 VDD.t70 15.4784
R3780 VDD.n1165 VDD.t59 15.4784
R3781 VDD.n2562 VDD.t66 15.4784
R3782 VDD.t62 VDD.n65 15.4784
R3783 VDD.n960 VDD.n959 14.1581
R3784 VDD.n2438 VDD.n2435 14.1581
R3785 VDD.n2673 VDD.n2670 14.1581
R3786 VDD.n1280 VDD.n692 14.1581
R3787 VDD.n961 VDD.n960 11.8308
R3788 VDD.n2435 VDD.n2430 11.8308
R3789 VDD.n2670 VDD.n157 11.8308
R3790 VDD.n1316 VDD.n692 11.8308
R3791 VDD.n1592 VDD.n672 11.6949
R3792 VDD.n1598 VDD.n672 11.6949
R3793 VDD.n1604 VDD.n666 11.6949
R3794 VDD.n1604 VDD.t50 11.6949
R3795 VDD.n1610 VDD.t50 11.6949
R3796 VDD.n1610 VDD.n655 11.6949
R3797 VDD.n1616 VDD.n655 11.6949
R3798 VDD.n1616 VDD.n649 11.6949
R3799 VDD.n1622 VDD.n649 11.6949
R3800 VDD.n1628 VDD.n643 11.6949
R3801 VDD.n1628 VDD.n637 11.6949
R3802 VDD.n1634 VDD.n637 11.6949
R3803 VDD.n1634 VDD.n631 11.6949
R3804 VDD.n1640 VDD.n631 11.6949
R3805 VDD.n1646 VDD.n625 11.6949
R3806 VDD.n1652 VDD.n619 11.6949
R3807 VDD.n1652 VDD.n613 11.6949
R3808 VDD.n1658 VDD.n613 11.6949
R3809 VDD.n1658 VDD.n607 11.6949
R3810 VDD.n1664 VDD.n607 11.6949
R3811 VDD.n1670 VDD.n601 11.6949
R3812 VDD.n1670 VDD.n595 11.6949
R3813 VDD.n1676 VDD.n595 11.6949
R3814 VDD.n1676 VDD.n589 11.6949
R3815 VDD.n1682 VDD.n589 11.6949
R3816 VDD.n1688 VDD.n583 11.6949
R3817 VDD.n1694 VDD.n577 11.6949
R3818 VDD.n1694 VDD.n571 11.6949
R3819 VDD.n1700 VDD.n571 11.6949
R3820 VDD.n1700 VDD.n564 11.6949
R3821 VDD.n1706 VDD.n564 11.6949
R3822 VDD.n1706 VDD.n567 11.6949
R3823 VDD.n1718 VDD.n553 11.6949
R3824 VDD.n1718 VDD.n547 11.6949
R3825 VDD.n1724 VDD.n547 11.6949
R3826 VDD.n1724 VDD.n540 11.6949
R3827 VDD.n1730 VDD.n540 11.6949
R3828 VDD.n1730 VDD.n543 11.6949
R3829 VDD.n1736 VDD.n528 11.6949
R3830 VDD.n1744 VDD.n528 11.6949
R3831 VDD.n1744 VDD.n522 11.6949
R3832 VDD.t40 VDD.n522 11.6949
R3833 VDD.t40 VDD.n511 11.6949
R3834 VDD.n1807 VDD.n511 11.6949
R3835 VDD.n1807 VDD.n514 11.6949
R3836 VDD.n1813 VDD.n476 11.6949
R3837 VDD.n2134 VDD.n1862 11.6949
R3838 VDD.n2140 VDD.n465 11.6949
R3839 VDD.n2146 VDD.n465 11.6949
R3840 VDD.n2146 VDD.t16 11.6949
R3841 VDD.n2152 VDD.t16 11.6949
R3842 VDD.n2152 VDD.n453 11.6949
R3843 VDD.n2158 VDD.n453 11.6949
R3844 VDD.n2158 VDD.n456 11.6949
R3845 VDD.n2164 VDD.n442 11.6949
R3846 VDD.n2170 VDD.n442 11.6949
R3847 VDD.n2170 VDD.n436 11.6949
R3848 VDD.n2176 VDD.n436 11.6949
R3849 VDD.n2176 VDD.n430 11.6949
R3850 VDD.n2182 VDD.n430 11.6949
R3851 VDD.n2188 VDD.n419 11.6949
R3852 VDD.n2194 VDD.n419 11.6949
R3853 VDD.n2194 VDD.n413 11.6949
R3854 VDD.n2200 VDD.n413 11.6949
R3855 VDD.n2200 VDD.n407 11.6949
R3856 VDD.n2206 VDD.n407 11.6949
R3857 VDD.n2212 VDD.n401 11.6949
R3858 VDD.n2218 VDD.n395 11.6949
R3859 VDD.n2218 VDD.n389 11.6949
R3860 VDD.n2224 VDD.n389 11.6949
R3861 VDD.n2224 VDD.n383 11.6949
R3862 VDD.n2230 VDD.n383 11.6949
R3863 VDD.n2236 VDD.n377 11.6949
R3864 VDD.n2236 VDD.n371 11.6949
R3865 VDD.n2242 VDD.n371 11.6949
R3866 VDD.n2242 VDD.n365 11.6949
R3867 VDD.n2248 VDD.n365 11.6949
R3868 VDD.n2254 VDD.n359 11.6949
R3869 VDD.n2260 VDD.n353 11.6949
R3870 VDD.n2260 VDD.n347 11.6949
R3871 VDD.n2266 VDD.n347 11.6949
R3872 VDD.n2266 VDD.n341 11.6949
R3873 VDD.n2272 VDD.n341 11.6949
R3874 VDD.n2278 VDD.n335 11.6949
R3875 VDD.n2278 VDD.n328 11.6949
R3876 VDD.n2286 VDD.n328 11.6949
R3877 VDD.n2286 VDD.n322 11.6949
R3878 VDD.t24 VDD.n322 11.6949
R3879 VDD.t24 VDD.n312 11.6949
R3880 VDD.n2349 VDD.n312 11.6949
R3881 VDD.n2355 VDD.n306 11.6949
R3882 VDD.n2355 VDD.n276 11.6949
R3883 VDD.n1682 VDD.t96 11.179
R3884 VDD.t81 VDD.n395 11.179
R3885 VDD.n1712 VDD.t91 10.835
R3886 VDD.n2063 VDD.t86 10.835
R3887 VDD.n2132 VDD.n469 10.6151
R3888 VDD.n2142 VDD.n469 10.6151
R3889 VDD.n2143 VDD.n2142 10.6151
R3890 VDD.n2144 VDD.n2143 10.6151
R3891 VDD.n2144 VDD.n458 10.6151
R3892 VDD.n2154 VDD.n458 10.6151
R3893 VDD.n2155 VDD.n2154 10.6151
R3894 VDD.n2156 VDD.n2155 10.6151
R3895 VDD.n2156 VDD.n446 10.6151
R3896 VDD.n2166 VDD.n446 10.6151
R3897 VDD.n2167 VDD.n2166 10.6151
R3898 VDD.n2168 VDD.n2167 10.6151
R3899 VDD.n2168 VDD.n434 10.6151
R3900 VDD.n2178 VDD.n434 10.6151
R3901 VDD.n2179 VDD.n2178 10.6151
R3902 VDD.n2180 VDD.n2179 10.6151
R3903 VDD.n2180 VDD.n423 10.6151
R3904 VDD.n2190 VDD.n423 10.6151
R3905 VDD.n2191 VDD.n2190 10.6151
R3906 VDD.n2192 VDD.n2191 10.6151
R3907 VDD.n2192 VDD.n411 10.6151
R3908 VDD.n2202 VDD.n411 10.6151
R3909 VDD.n2203 VDD.n2202 10.6151
R3910 VDD.n2204 VDD.n2203 10.6151
R3911 VDD.n2204 VDD.n399 10.6151
R3912 VDD.n2214 VDD.n399 10.6151
R3913 VDD.n2215 VDD.n2214 10.6151
R3914 VDD.n2216 VDD.n2215 10.6151
R3915 VDD.n2216 VDD.n387 10.6151
R3916 VDD.n2226 VDD.n387 10.6151
R3917 VDD.n2227 VDD.n2226 10.6151
R3918 VDD.n2228 VDD.n2227 10.6151
R3919 VDD.n2228 VDD.n375 10.6151
R3920 VDD.n2238 VDD.n375 10.6151
R3921 VDD.n2239 VDD.n2238 10.6151
R3922 VDD.n2240 VDD.n2239 10.6151
R3923 VDD.n2240 VDD.n363 10.6151
R3924 VDD.n2250 VDD.n363 10.6151
R3925 VDD.n2251 VDD.n2250 10.6151
R3926 VDD.n2252 VDD.n2251 10.6151
R3927 VDD.n2252 VDD.n351 10.6151
R3928 VDD.n2262 VDD.n351 10.6151
R3929 VDD.n2263 VDD.n2262 10.6151
R3930 VDD.n2264 VDD.n2263 10.6151
R3931 VDD.n2264 VDD.n339 10.6151
R3932 VDD.n2274 VDD.n339 10.6151
R3933 VDD.n2275 VDD.n2274 10.6151
R3934 VDD.n2276 VDD.n2275 10.6151
R3935 VDD.n2276 VDD.n326 10.6151
R3936 VDD.n2288 VDD.n326 10.6151
R3937 VDD.n2289 VDD.n2288 10.6151
R3938 VDD.n2290 VDD.n2289 10.6151
R3939 VDD.n2290 VDD.n310 10.6151
R3940 VDD.n2351 VDD.n310 10.6151
R3941 VDD.n2352 VDD.n2351 10.6151
R3942 VDD.n2353 VDD.n2352 10.6151
R3943 VDD.n2353 VDD.n300 10.6151
R3944 VDD.n2398 VDD.n2397 10.6151
R3945 VDD.n2397 VDD.n2396 10.6151
R3946 VDD.n2396 VDD.n2393 10.6151
R3947 VDD.n2393 VDD.n2392 10.6151
R3948 VDD.n2392 VDD.n2389 10.6151
R3949 VDD.n2389 VDD.n2388 10.6151
R3950 VDD.n2388 VDD.n2385 10.6151
R3951 VDD.n2385 VDD.n2384 10.6151
R3952 VDD.n2384 VDD.n2381 10.6151
R3953 VDD.n2381 VDD.n2380 10.6151
R3954 VDD.n2380 VDD.n2377 10.6151
R3955 VDD.n2377 VDD.n2376 10.6151
R3956 VDD.n2376 VDD.n2373 10.6151
R3957 VDD.n2373 VDD.n2372 10.6151
R3958 VDD.n2372 VDD.n2369 10.6151
R3959 VDD.n2369 VDD.n2368 10.6151
R3960 VDD.n2368 VDD.n2365 10.6151
R3961 VDD.n2363 VDD.n2360 10.6151
R3962 VDD.n2360 VDD.n2359 10.6151
R3963 VDD.n2090 VDD.n2089 10.6151
R3964 VDD.n2089 VDD.n2087 10.6151
R3965 VDD.n2087 VDD.n2086 10.6151
R3966 VDD.n2086 VDD.n2084 10.6151
R3967 VDD.n2084 VDD.n2083 10.6151
R3968 VDD.n2083 VDD.n2081 10.6151
R3969 VDD.n2081 VDD.n2080 10.6151
R3970 VDD.n2080 VDD.n2078 10.6151
R3971 VDD.n2078 VDD.n2077 10.6151
R3972 VDD.n2077 VDD.n2075 10.6151
R3973 VDD.n2075 VDD.n2074 10.6151
R3974 VDD.n2074 VDD.n2072 10.6151
R3975 VDD.n2072 VDD.n2071 10.6151
R3976 VDD.n2071 VDD.n2069 10.6151
R3977 VDD.n2069 VDD.n2068 10.6151
R3978 VDD.n2068 VDD.n2066 10.6151
R3979 VDD.n2066 VDD.n2065 10.6151
R3980 VDD.n2065 VDD.n1932 10.6151
R3981 VDD.n1932 VDD.n1931 10.6151
R3982 VDD.n1931 VDD.n1929 10.6151
R3983 VDD.n1929 VDD.n1928 10.6151
R3984 VDD.n1928 VDD.n1926 10.6151
R3985 VDD.n1926 VDD.n1925 10.6151
R3986 VDD.n1925 VDD.n1923 10.6151
R3987 VDD.n1923 VDD.n1922 10.6151
R3988 VDD.n1922 VDD.n1920 10.6151
R3989 VDD.n1920 VDD.n1919 10.6151
R3990 VDD.n1919 VDD.n1917 10.6151
R3991 VDD.n1917 VDD.n1916 10.6151
R3992 VDD.n1916 VDD.n1914 10.6151
R3993 VDD.n1914 VDD.n1913 10.6151
R3994 VDD.n1913 VDD.n1911 10.6151
R3995 VDD.n1911 VDD.n1910 10.6151
R3996 VDD.n1910 VDD.n1908 10.6151
R3997 VDD.n1908 VDD.n1907 10.6151
R3998 VDD.n1907 VDD.n1905 10.6151
R3999 VDD.n1905 VDD.n1904 10.6151
R4000 VDD.n1904 VDD.n1902 10.6151
R4001 VDD.n1902 VDD.n1901 10.6151
R4002 VDD.n1901 VDD.n1899 10.6151
R4003 VDD.n1899 VDD.n1898 10.6151
R4004 VDD.n1898 VDD.n1896 10.6151
R4005 VDD.n1896 VDD.n1895 10.6151
R4006 VDD.n1895 VDD.n1893 10.6151
R4007 VDD.n1893 VDD.n1892 10.6151
R4008 VDD.n1892 VDD.n1890 10.6151
R4009 VDD.n1890 VDD.n1889 10.6151
R4010 VDD.n1889 VDD.n1887 10.6151
R4011 VDD.n1887 VDD.n1886 10.6151
R4012 VDD.n1886 VDD.n1884 10.6151
R4013 VDD.n1884 VDD.n1883 10.6151
R4014 VDD.n1883 VDD.n1881 10.6151
R4015 VDD.n1881 VDD.n1880 10.6151
R4016 VDD.n1880 VDD.n1878 10.6151
R4017 VDD.n1878 VDD.n1877 10.6151
R4018 VDD.n1877 VDD.n305 10.6151
R4019 VDD.n305 VDD.n303 10.6151
R4020 VDD.n2131 VDD.n2130 10.6151
R4021 VDD.n2130 VDD.n1864 10.6151
R4022 VDD.n2125 VDD.n1864 10.6151
R4023 VDD.n2125 VDD.n2124 10.6151
R4024 VDD.n2124 VDD.n1866 10.6151
R4025 VDD.n2119 VDD.n1866 10.6151
R4026 VDD.n2119 VDD.n2118 10.6151
R4027 VDD.n2118 VDD.n2117 10.6151
R4028 VDD.n2117 VDD.n1868 10.6151
R4029 VDD.n2111 VDD.n1868 10.6151
R4030 VDD.n2111 VDD.n2110 10.6151
R4031 VDD.n2110 VDD.n2109 10.6151
R4032 VDD.n2109 VDD.n1870 10.6151
R4033 VDD.n2103 VDD.n1870 10.6151
R4034 VDD.n2103 VDD.n2102 10.6151
R4035 VDD.n2102 VDD.n2101 10.6151
R4036 VDD.n2101 VDD.n1872 10.6151
R4037 VDD.n2095 VDD.n2094 10.6151
R4038 VDD.n2094 VDD.n2093 10.6151
R4039 VDD.n1856 VDD.n1855 10.6151
R4040 VDD.n1855 VDD.n1854 10.6151
R4041 VDD.n1854 VDD.n1851 10.6151
R4042 VDD.n1851 VDD.n1850 10.6151
R4043 VDD.n1850 VDD.n1847 10.6151
R4044 VDD.n1847 VDD.n1846 10.6151
R4045 VDD.n1846 VDD.n1843 10.6151
R4046 VDD.n1843 VDD.n1842 10.6151
R4047 VDD.n1842 VDD.n1839 10.6151
R4048 VDD.n1839 VDD.n1838 10.6151
R4049 VDD.n1838 VDD.n1835 10.6151
R4050 VDD.n1835 VDD.n1834 10.6151
R4051 VDD.n1834 VDD.n1831 10.6151
R4052 VDD.n1831 VDD.n1830 10.6151
R4053 VDD.n1830 VDD.n1827 10.6151
R4054 VDD.n1827 VDD.n1826 10.6151
R4055 VDD.n1826 VDD.n1823 10.6151
R4056 VDD.n1821 VDD.n1818 10.6151
R4057 VDD.n1818 VDD.n1817 10.6151
R4058 VDD.n1548 VDD.n1547 10.6151
R4059 VDD.n1547 VDD.n1545 10.6151
R4060 VDD.n1545 VDD.n1544 10.6151
R4061 VDD.n1544 VDD.n1542 10.6151
R4062 VDD.n1542 VDD.n1541 10.6151
R4063 VDD.n1541 VDD.n1539 10.6151
R4064 VDD.n1539 VDD.n1538 10.6151
R4065 VDD.n1538 VDD.n1536 10.6151
R4066 VDD.n1536 VDD.n1535 10.6151
R4067 VDD.n1535 VDD.n1533 10.6151
R4068 VDD.n1533 VDD.n1532 10.6151
R4069 VDD.n1532 VDD.n1530 10.6151
R4070 VDD.n1530 VDD.n1529 10.6151
R4071 VDD.n1529 VDD.n1527 10.6151
R4072 VDD.n1527 VDD.n1526 10.6151
R4073 VDD.n1526 VDD.n1524 10.6151
R4074 VDD.n1524 VDD.n1523 10.6151
R4075 VDD.n1523 VDD.n1521 10.6151
R4076 VDD.n1521 VDD.n1520 10.6151
R4077 VDD.n1520 VDD.n1518 10.6151
R4078 VDD.n1518 VDD.n1517 10.6151
R4079 VDD.n1517 VDD.n1515 10.6151
R4080 VDD.n1515 VDD.n1514 10.6151
R4081 VDD.n1514 VDD.n1512 10.6151
R4082 VDD.n1512 VDD.n1511 10.6151
R4083 VDD.n1511 VDD.n1509 10.6151
R4084 VDD.n1509 VDD.n1508 10.6151
R4085 VDD.n1508 VDD.n1506 10.6151
R4086 VDD.n1506 VDD.n1505 10.6151
R4087 VDD.n1505 VDD.n1503 10.6151
R4088 VDD.n1503 VDD.n1502 10.6151
R4089 VDD.n1502 VDD.n1500 10.6151
R4090 VDD.n1500 VDD.n1499 10.6151
R4091 VDD.n1499 VDD.n1497 10.6151
R4092 VDD.n1497 VDD.n1496 10.6151
R4093 VDD.n1496 VDD.n1494 10.6151
R4094 VDD.n1494 VDD.n1493 10.6151
R4095 VDD.n1493 VDD.n1491 10.6151
R4096 VDD.n1491 VDD.n1490 10.6151
R4097 VDD.n1490 VDD.n1488 10.6151
R4098 VDD.n1488 VDD.n1487 10.6151
R4099 VDD.n1487 VDD.n1485 10.6151
R4100 VDD.n1485 VDD.n1484 10.6151
R4101 VDD.n1484 VDD.n1482 10.6151
R4102 VDD.n1482 VDD.n1481 10.6151
R4103 VDD.n1481 VDD.n1479 10.6151
R4104 VDD.n1479 VDD.n1478 10.6151
R4105 VDD.n1478 VDD.n1476 10.6151
R4106 VDD.n1476 VDD.n1475 10.6151
R4107 VDD.n1475 VDD.n1473 10.6151
R4108 VDD.n1473 VDD.n1472 10.6151
R4109 VDD.n1472 VDD.n1470 10.6151
R4110 VDD.n1470 VDD.n1469 10.6151
R4111 VDD.n1469 VDD.n1467 10.6151
R4112 VDD.n1467 VDD.n1466 10.6151
R4113 VDD.n1466 VDD.n505 10.6151
R4114 VDD.n505 VDD.n503 10.6151
R4115 VDD.n1589 VDD.n1588 10.6151
R4116 VDD.n1588 VDD.n1453 10.6151
R4117 VDD.n1583 VDD.n1453 10.6151
R4118 VDD.n1583 VDD.n1582 10.6151
R4119 VDD.n1582 VDD.n1455 10.6151
R4120 VDD.n1577 VDD.n1455 10.6151
R4121 VDD.n1577 VDD.n1576 10.6151
R4122 VDD.n1576 VDD.n1575 10.6151
R4123 VDD.n1575 VDD.n1457 10.6151
R4124 VDD.n1569 VDD.n1457 10.6151
R4125 VDD.n1569 VDD.n1568 10.6151
R4126 VDD.n1568 VDD.n1567 10.6151
R4127 VDD.n1567 VDD.n1459 10.6151
R4128 VDD.n1561 VDD.n1459 10.6151
R4129 VDD.n1561 VDD.n1560 10.6151
R4130 VDD.n1560 VDD.n1559 10.6151
R4131 VDD.n1559 VDD.n1461 10.6151
R4132 VDD.n1553 VDD.n1552 10.6151
R4133 VDD.n1552 VDD.n1551 10.6151
R4134 VDD.n1590 VDD.n670 10.6151
R4135 VDD.n1600 VDD.n670 10.6151
R4136 VDD.n1601 VDD.n1600 10.6151
R4137 VDD.n1602 VDD.n1601 10.6151
R4138 VDD.n1602 VDD.n659 10.6151
R4139 VDD.n1612 VDD.n659 10.6151
R4140 VDD.n1613 VDD.n1612 10.6151
R4141 VDD.n1614 VDD.n1613 10.6151
R4142 VDD.n1614 VDD.n647 10.6151
R4143 VDD.n1624 VDD.n647 10.6151
R4144 VDD.n1625 VDD.n1624 10.6151
R4145 VDD.n1626 VDD.n1625 10.6151
R4146 VDD.n1626 VDD.n635 10.6151
R4147 VDD.n1636 VDD.n635 10.6151
R4148 VDD.n1637 VDD.n1636 10.6151
R4149 VDD.n1638 VDD.n1637 10.6151
R4150 VDD.n1638 VDD.n623 10.6151
R4151 VDD.n1648 VDD.n623 10.6151
R4152 VDD.n1649 VDD.n1648 10.6151
R4153 VDD.n1650 VDD.n1649 10.6151
R4154 VDD.n1650 VDD.n611 10.6151
R4155 VDD.n1660 VDD.n611 10.6151
R4156 VDD.n1661 VDD.n1660 10.6151
R4157 VDD.n1662 VDD.n1661 10.6151
R4158 VDD.n1662 VDD.n599 10.6151
R4159 VDD.n1672 VDD.n599 10.6151
R4160 VDD.n1673 VDD.n1672 10.6151
R4161 VDD.n1674 VDD.n1673 10.6151
R4162 VDD.n1674 VDD.n587 10.6151
R4163 VDD.n1684 VDD.n587 10.6151
R4164 VDD.n1685 VDD.n1684 10.6151
R4165 VDD.n1686 VDD.n1685 10.6151
R4166 VDD.n1686 VDD.n575 10.6151
R4167 VDD.n1696 VDD.n575 10.6151
R4168 VDD.n1697 VDD.n1696 10.6151
R4169 VDD.n1698 VDD.n1697 10.6151
R4170 VDD.n1698 VDD.n562 10.6151
R4171 VDD.n1708 VDD.n562 10.6151
R4172 VDD.n1709 VDD.n1708 10.6151
R4173 VDD.n1710 VDD.n1709 10.6151
R4174 VDD.n1710 VDD.n551 10.6151
R4175 VDD.n1720 VDD.n551 10.6151
R4176 VDD.n1721 VDD.n1720 10.6151
R4177 VDD.n1722 VDD.n1721 10.6151
R4178 VDD.n1722 VDD.n538 10.6151
R4179 VDD.n1732 VDD.n538 10.6151
R4180 VDD.n1733 VDD.n1732 10.6151
R4181 VDD.n1734 VDD.n1733 10.6151
R4182 VDD.n1734 VDD.n526 10.6151
R4183 VDD.n1746 VDD.n526 10.6151
R4184 VDD.n1747 VDD.n1746 10.6151
R4185 VDD.n1748 VDD.n1747 10.6151
R4186 VDD.n1748 VDD.n509 10.6151
R4187 VDD.n1809 VDD.n509 10.6151
R4188 VDD.n1810 VDD.n1809 10.6151
R4189 VDD.n1811 VDD.n1810 10.6151
R4190 VDD.n1811 VDD.n500 10.6151
R4191 VDD.n2342 VDD.n2341 10.6151
R4192 VDD.n2341 VDD.n2339 10.6151
R4193 VDD.n2339 VDD.n2336 10.6151
R4194 VDD.n2336 VDD.n2335 10.6151
R4195 VDD.n2335 VDD.n2332 10.6151
R4196 VDD.n2332 VDD.n2331 10.6151
R4197 VDD.n2331 VDD.n2328 10.6151
R4198 VDD.n2328 VDD.n2327 10.6151
R4199 VDD.n2327 VDD.n2324 10.6151
R4200 VDD.n2324 VDD.n2323 10.6151
R4201 VDD.n2323 VDD.n2320 10.6151
R4202 VDD.n2320 VDD.n2319 10.6151
R4203 VDD.n2319 VDD.n2316 10.6151
R4204 VDD.n2316 VDD.n2315 10.6151
R4205 VDD.n2315 VDD.n2312 10.6151
R4206 VDD.n2312 VDD.n2311 10.6151
R4207 VDD.n2311 VDD.n2308 10.6151
R4208 VDD.n2306 VDD.n2303 10.6151
R4209 VDD.n2303 VDD.n2302 10.6151
R4210 VDD.n1988 VDD.n1986 10.6151
R4211 VDD.n1989 VDD.n1988 10.6151
R4212 VDD.n1991 VDD.n1989 10.6151
R4213 VDD.n1992 VDD.n1991 10.6151
R4214 VDD.n1994 VDD.n1992 10.6151
R4215 VDD.n1995 VDD.n1994 10.6151
R4216 VDD.n1997 VDD.n1995 10.6151
R4217 VDD.n1998 VDD.n1997 10.6151
R4218 VDD.n2000 VDD.n1998 10.6151
R4219 VDD.n2001 VDD.n2000 10.6151
R4220 VDD.n2003 VDD.n2001 10.6151
R4221 VDD.n2004 VDD.n2003 10.6151
R4222 VDD.n2006 VDD.n2004 10.6151
R4223 VDD.n2007 VDD.n2006 10.6151
R4224 VDD.n2009 VDD.n2007 10.6151
R4225 VDD.n2010 VDD.n2009 10.6151
R4226 VDD.n2061 VDD.n2010 10.6151
R4227 VDD.n2061 VDD.n2060 10.6151
R4228 VDD.n2060 VDD.n2059 10.6151
R4229 VDD.n2059 VDD.n2057 10.6151
R4230 VDD.n2057 VDD.n2056 10.6151
R4231 VDD.n2056 VDD.n2054 10.6151
R4232 VDD.n2054 VDD.n2053 10.6151
R4233 VDD.n2053 VDD.n2051 10.6151
R4234 VDD.n2051 VDD.n2050 10.6151
R4235 VDD.n2050 VDD.n2048 10.6151
R4236 VDD.n2048 VDD.n2047 10.6151
R4237 VDD.n2047 VDD.n2045 10.6151
R4238 VDD.n2045 VDD.n2044 10.6151
R4239 VDD.n2044 VDD.n2042 10.6151
R4240 VDD.n2042 VDD.n2041 10.6151
R4241 VDD.n2041 VDD.n2039 10.6151
R4242 VDD.n2039 VDD.n2038 10.6151
R4243 VDD.n2038 VDD.n2036 10.6151
R4244 VDD.n2036 VDD.n2035 10.6151
R4245 VDD.n2035 VDD.n2033 10.6151
R4246 VDD.n2033 VDD.n2032 10.6151
R4247 VDD.n2032 VDD.n2030 10.6151
R4248 VDD.n2030 VDD.n2029 10.6151
R4249 VDD.n2029 VDD.n2027 10.6151
R4250 VDD.n2027 VDD.n2026 10.6151
R4251 VDD.n2026 VDD.n2024 10.6151
R4252 VDD.n2024 VDD.n2023 10.6151
R4253 VDD.n2023 VDD.n2021 10.6151
R4254 VDD.n2021 VDD.n2020 10.6151
R4255 VDD.n2020 VDD.n2018 10.6151
R4256 VDD.n2018 VDD.n2017 10.6151
R4257 VDD.n2017 VDD.n2015 10.6151
R4258 VDD.n2015 VDD.n2014 10.6151
R4259 VDD.n2014 VDD.n2012 10.6151
R4260 VDD.n2012 VDD.n2011 10.6151
R4261 VDD.n2011 VDD.n320 10.6151
R4262 VDD.n2294 VDD.n320 10.6151
R4263 VDD.n2295 VDD.n2294 10.6151
R4264 VDD.n2297 VDD.n2295 10.6151
R4265 VDD.n2298 VDD.n2297 10.6151
R4266 VDD.n2299 VDD.n2298 10.6151
R4267 VDD.n1946 VDD.n474 10.6151
R4268 VDD.n1947 VDD.n1946 10.6151
R4269 VDD.n1947 VDD.n1943 10.6151
R4270 VDD.n1953 VDD.n1943 10.6151
R4271 VDD.n1954 VDD.n1953 10.6151
R4272 VDD.n1955 VDD.n1954 10.6151
R4273 VDD.n1955 VDD.n1941 10.6151
R4274 VDD.n1961 VDD.n1941 10.6151
R4275 VDD.n1962 VDD.n1961 10.6151
R4276 VDD.n1963 VDD.n1962 10.6151
R4277 VDD.n1963 VDD.n1939 10.6151
R4278 VDD.n1969 VDD.n1939 10.6151
R4279 VDD.n1970 VDD.n1969 10.6151
R4280 VDD.n1971 VDD.n1970 10.6151
R4281 VDD.n1971 VDD.n1937 10.6151
R4282 VDD.n1977 VDD.n1937 10.6151
R4283 VDD.n1978 VDD.n1977 10.6151
R4284 VDD.n1980 VDD.n1933 10.6151
R4285 VDD.n1985 VDD.n1933 10.6151
R4286 VDD.n2137 VDD.n2136 10.6151
R4287 VDD.n2138 VDD.n2137 10.6151
R4288 VDD.n2138 VDD.n463 10.6151
R4289 VDD.n2148 VDD.n463 10.6151
R4290 VDD.n2149 VDD.n2148 10.6151
R4291 VDD.n2150 VDD.n2149 10.6151
R4292 VDD.n2150 VDD.n451 10.6151
R4293 VDD.n2160 VDD.n451 10.6151
R4294 VDD.n2161 VDD.n2160 10.6151
R4295 VDD.n2162 VDD.n2161 10.6151
R4296 VDD.n2162 VDD.n440 10.6151
R4297 VDD.n2172 VDD.n440 10.6151
R4298 VDD.n2173 VDD.n2172 10.6151
R4299 VDD.n2174 VDD.n2173 10.6151
R4300 VDD.n2174 VDD.n428 10.6151
R4301 VDD.n2184 VDD.n428 10.6151
R4302 VDD.n2185 VDD.n2184 10.6151
R4303 VDD.n2186 VDD.n2185 10.6151
R4304 VDD.n2186 VDD.n417 10.6151
R4305 VDD.n2196 VDD.n417 10.6151
R4306 VDD.n2197 VDD.n2196 10.6151
R4307 VDD.n2198 VDD.n2197 10.6151
R4308 VDD.n2198 VDD.n405 10.6151
R4309 VDD.n2208 VDD.n405 10.6151
R4310 VDD.n2209 VDD.n2208 10.6151
R4311 VDD.n2210 VDD.n2209 10.6151
R4312 VDD.n2210 VDD.n393 10.6151
R4313 VDD.n2220 VDD.n393 10.6151
R4314 VDD.n2221 VDD.n2220 10.6151
R4315 VDD.n2222 VDD.n2221 10.6151
R4316 VDD.n2222 VDD.n381 10.6151
R4317 VDD.n2232 VDD.n381 10.6151
R4318 VDD.n2233 VDD.n2232 10.6151
R4319 VDD.n2234 VDD.n2233 10.6151
R4320 VDD.n2234 VDD.n369 10.6151
R4321 VDD.n2244 VDD.n369 10.6151
R4322 VDD.n2245 VDD.n2244 10.6151
R4323 VDD.n2246 VDD.n2245 10.6151
R4324 VDD.n2246 VDD.n357 10.6151
R4325 VDD.n2256 VDD.n357 10.6151
R4326 VDD.n2257 VDD.n2256 10.6151
R4327 VDD.n2258 VDD.n2257 10.6151
R4328 VDD.n2258 VDD.n345 10.6151
R4329 VDD.n2268 VDD.n345 10.6151
R4330 VDD.n2269 VDD.n2268 10.6151
R4331 VDD.n2270 VDD.n2269 10.6151
R4332 VDD.n2270 VDD.n333 10.6151
R4333 VDD.n2280 VDD.n333 10.6151
R4334 VDD.n2281 VDD.n2280 10.6151
R4335 VDD.n2284 VDD.n2281 10.6151
R4336 VDD.n2284 VDD.n2283 10.6151
R4337 VDD.n2283 VDD.n2282 10.6151
R4338 VDD.n2282 VDD.n317 10.6151
R4339 VDD.n2347 VDD.n317 10.6151
R4340 VDD.n2347 VDD.n2346 10.6151
R4341 VDD.n2346 VDD.n2345 10.6151
R4342 VDD.n2345 VDD.n2344 10.6151
R4343 VDD.n1800 VDD.n1799 10.6151
R4344 VDD.n1799 VDD.n1797 10.6151
R4345 VDD.n1797 VDD.n1794 10.6151
R4346 VDD.n1794 VDD.n1793 10.6151
R4347 VDD.n1793 VDD.n1790 10.6151
R4348 VDD.n1790 VDD.n1789 10.6151
R4349 VDD.n1789 VDD.n1786 10.6151
R4350 VDD.n1786 VDD.n1785 10.6151
R4351 VDD.n1785 VDD.n1782 10.6151
R4352 VDD.n1782 VDD.n1781 10.6151
R4353 VDD.n1781 VDD.n1778 10.6151
R4354 VDD.n1778 VDD.n1777 10.6151
R4355 VDD.n1777 VDD.n1774 10.6151
R4356 VDD.n1774 VDD.n1773 10.6151
R4357 VDD.n1773 VDD.n1770 10.6151
R4358 VDD.n1770 VDD.n1769 10.6151
R4359 VDD.n1769 VDD.n1766 10.6151
R4360 VDD.n1764 VDD.n1761 10.6151
R4361 VDD.n1761 VDD.n1760 10.6151
R4362 VDD.n1450 VDD.n1449 10.6151
R4363 VDD.n1449 VDD.n1448 10.6151
R4364 VDD.n1448 VDD.n1447 10.6151
R4365 VDD.n1447 VDD.n1445 10.6151
R4366 VDD.n1445 VDD.n1444 10.6151
R4367 VDD.n1444 VDD.n1442 10.6151
R4368 VDD.n1442 VDD.n1441 10.6151
R4369 VDD.n1441 VDD.n1439 10.6151
R4370 VDD.n1439 VDD.n1438 10.6151
R4371 VDD.n1438 VDD.n1436 10.6151
R4372 VDD.n1436 VDD.n1435 10.6151
R4373 VDD.n1435 VDD.n1433 10.6151
R4374 VDD.n1433 VDD.n1432 10.6151
R4375 VDD.n1432 VDD.n1430 10.6151
R4376 VDD.n1430 VDD.n1429 10.6151
R4377 VDD.n1429 VDD.n1427 10.6151
R4378 VDD.n1427 VDD.n1426 10.6151
R4379 VDD.n1426 VDD.n1424 10.6151
R4380 VDD.n1424 VDD.n1423 10.6151
R4381 VDD.n1423 VDD.n1421 10.6151
R4382 VDD.n1421 VDD.n1420 10.6151
R4383 VDD.n1420 VDD.n1418 10.6151
R4384 VDD.n1418 VDD.n1417 10.6151
R4385 VDD.n1417 VDD.n1415 10.6151
R4386 VDD.n1415 VDD.n1414 10.6151
R4387 VDD.n1414 VDD.n1412 10.6151
R4388 VDD.n1412 VDD.n1411 10.6151
R4389 VDD.n1411 VDD.n1409 10.6151
R4390 VDD.n1409 VDD.n1408 10.6151
R4391 VDD.n1408 VDD.n1406 10.6151
R4392 VDD.n1406 VDD.n1405 10.6151
R4393 VDD.n1405 VDD.n1403 10.6151
R4394 VDD.n1403 VDD.n1402 10.6151
R4395 VDD.n1402 VDD.n1400 10.6151
R4396 VDD.n1400 VDD.n1399 10.6151
R4397 VDD.n1399 VDD.n1397 10.6151
R4398 VDD.n1397 VDD.n1396 10.6151
R4399 VDD.n1396 VDD.n1394 10.6151
R4400 VDD.n1394 VDD.n1393 10.6151
R4401 VDD.n1393 VDD.n1391 10.6151
R4402 VDD.n1391 VDD.n1390 10.6151
R4403 VDD.n1390 VDD.n1388 10.6151
R4404 VDD.n1388 VDD.n1387 10.6151
R4405 VDD.n1387 VDD.n1385 10.6151
R4406 VDD.n1385 VDD.n1384 10.6151
R4407 VDD.n1384 VDD.n1382 10.6151
R4408 VDD.n1382 VDD.n1381 10.6151
R4409 VDD.n1381 VDD.n1379 10.6151
R4410 VDD.n1379 VDD.n1378 10.6151
R4411 VDD.n1378 VDD.n1376 10.6151
R4412 VDD.n1376 VDD.n1375 10.6151
R4413 VDD.n1375 VDD.n520 10.6151
R4414 VDD.n1752 VDD.n520 10.6151
R4415 VDD.n1753 VDD.n1752 10.6151
R4416 VDD.n1755 VDD.n1753 10.6151
R4417 VDD.n1756 VDD.n1755 10.6151
R4418 VDD.n1757 VDD.n1756 10.6151
R4419 VDD.n1335 VDD.n676 10.6151
R4420 VDD.n1340 VDD.n1335 10.6151
R4421 VDD.n1341 VDD.n1340 10.6151
R4422 VDD.n1342 VDD.n1341 10.6151
R4423 VDD.n1342 VDD.n1333 10.6151
R4424 VDD.n1348 VDD.n1333 10.6151
R4425 VDD.n1349 VDD.n1348 10.6151
R4426 VDD.n1350 VDD.n1349 10.6151
R4427 VDD.n1350 VDD.n1331 10.6151
R4428 VDD.n1356 VDD.n1331 10.6151
R4429 VDD.n1357 VDD.n1356 10.6151
R4430 VDD.n1358 VDD.n1357 10.6151
R4431 VDD.n1358 VDD.n1329 10.6151
R4432 VDD.n1364 VDD.n1329 10.6151
R4433 VDD.n1365 VDD.n1364 10.6151
R4434 VDD.n1366 VDD.n1365 10.6151
R4435 VDD.n1366 VDD.n1327 10.6151
R4436 VDD.n1373 VDD.n1323 10.6151
R4437 VDD.n1374 VDD.n1373 10.6151
R4438 VDD.n1595 VDD.n1594 10.6151
R4439 VDD.n1596 VDD.n1595 10.6151
R4440 VDD.n1596 VDD.n664 10.6151
R4441 VDD.n1606 VDD.n664 10.6151
R4442 VDD.n1607 VDD.n1606 10.6151
R4443 VDD.n1608 VDD.n1607 10.6151
R4444 VDD.n1608 VDD.n653 10.6151
R4445 VDD.n1618 VDD.n653 10.6151
R4446 VDD.n1619 VDD.n1618 10.6151
R4447 VDD.n1620 VDD.n1619 10.6151
R4448 VDD.n1620 VDD.n641 10.6151
R4449 VDD.n1630 VDD.n641 10.6151
R4450 VDD.n1631 VDD.n1630 10.6151
R4451 VDD.n1632 VDD.n1631 10.6151
R4452 VDD.n1632 VDD.n629 10.6151
R4453 VDD.n1642 VDD.n629 10.6151
R4454 VDD.n1643 VDD.n1642 10.6151
R4455 VDD.n1644 VDD.n1643 10.6151
R4456 VDD.n1644 VDD.n617 10.6151
R4457 VDD.n1654 VDD.n617 10.6151
R4458 VDD.n1655 VDD.n1654 10.6151
R4459 VDD.n1656 VDD.n1655 10.6151
R4460 VDD.n1656 VDD.n605 10.6151
R4461 VDD.n1666 VDD.n605 10.6151
R4462 VDD.n1667 VDD.n1666 10.6151
R4463 VDD.n1668 VDD.n1667 10.6151
R4464 VDD.n1668 VDD.n593 10.6151
R4465 VDD.n1678 VDD.n593 10.6151
R4466 VDD.n1679 VDD.n1678 10.6151
R4467 VDD.n1680 VDD.n1679 10.6151
R4468 VDD.n1680 VDD.n581 10.6151
R4469 VDD.n1690 VDD.n581 10.6151
R4470 VDD.n1691 VDD.n1690 10.6151
R4471 VDD.n1692 VDD.n1691 10.6151
R4472 VDD.n1692 VDD.n569 10.6151
R4473 VDD.n1702 VDD.n569 10.6151
R4474 VDD.n1703 VDD.n1702 10.6151
R4475 VDD.n1704 VDD.n1703 10.6151
R4476 VDD.n1704 VDD.n557 10.6151
R4477 VDD.n1714 VDD.n557 10.6151
R4478 VDD.n1715 VDD.n1714 10.6151
R4479 VDD.n1716 VDD.n1715 10.6151
R4480 VDD.n1716 VDD.n545 10.6151
R4481 VDD.n1726 VDD.n545 10.6151
R4482 VDD.n1727 VDD.n1726 10.6151
R4483 VDD.n1728 VDD.n1727 10.6151
R4484 VDD.n1728 VDD.n533 10.6151
R4485 VDD.n1738 VDD.n533 10.6151
R4486 VDD.n1739 VDD.n1738 10.6151
R4487 VDD.n1742 VDD.n1739 10.6151
R4488 VDD.n1742 VDD.n1741 10.6151
R4489 VDD.n1741 VDD.n1740 10.6151
R4490 VDD.n1740 VDD.n517 10.6151
R4491 VDD.n1805 VDD.n517 10.6151
R4492 VDD.n1805 VDD.n1804 10.6151
R4493 VDD.n1804 VDD.n1803 10.6151
R4494 VDD.n1803 VDD.n1802 10.6151
R4495 VDD.n29 VDD.n27 9.84608
R4496 VDD.n20 VDD.n18 9.84608
R4497 VDD.n1113 VDD.n1111 9.84608
R4498 VDD.n1104 VDD.n1102 9.84608
R4499 VDD.n1736 VDD.t78 9.45923
R4500 VDD.n456 VDD.t75 9.45923
R4501 VDD.n32 VDD.n31 9.45567
R4502 VDD.n23 VDD.n22 9.45567
R4503 VDD.n1116 VDD.n1115 9.45567
R4504 VDD.n1107 VDD.n1106 9.45567
R4505 VDD.n31 VDD.n30 9.3005
R4506 VDD.n22 VDD.n21 9.3005
R4507 VDD.n2707 VDD.n2706 9.3005
R4508 VDD.n2705 VDD.n142 9.3005
R4509 VDD.n2704 VDD.n2703 9.3005
R4510 VDD.n2700 VDD.n143 9.3005
R4511 VDD.n2697 VDD.n144 9.3005
R4512 VDD.n2696 VDD.n145 9.3005
R4513 VDD.n2693 VDD.n146 9.3005
R4514 VDD.n2689 VDD.n147 9.3005
R4515 VDD.n2686 VDD.n148 9.3005
R4516 VDD.n2685 VDD.n149 9.3005
R4517 VDD.n2682 VDD.n150 9.3005
R4518 VDD.n2681 VDD.n151 9.3005
R4519 VDD.n2678 VDD.n152 9.3005
R4520 VDD.n2677 VDD.n153 9.3005
R4521 VDD.n2674 VDD.n154 9.3005
R4522 VDD.n2673 VDD.n155 9.3005
R4523 VDD.n2670 VDD.n2669 9.3005
R4524 VDD.n2668 VDD.n157 9.3005
R4525 VDD.n2708 VDD.n141 9.3005
R4526 VDD.n2478 VDD.n273 9.3005
R4527 VDD.n2480 VDD.n2479 9.3005
R4528 VDD.n263 VDD.n262 9.3005
R4529 VDD.n2493 VDD.n2492 9.3005
R4530 VDD.n2494 VDD.n261 9.3005
R4531 VDD.n2496 VDD.n2495 9.3005
R4532 VDD.n251 VDD.n250 9.3005
R4533 VDD.n2509 VDD.n2508 9.3005
R4534 VDD.n2510 VDD.n249 9.3005
R4535 VDD.n2512 VDD.n2511 9.3005
R4536 VDD.n239 VDD.n238 9.3005
R4537 VDD.n2525 VDD.n2524 9.3005
R4538 VDD.n2526 VDD.n237 9.3005
R4539 VDD.n2528 VDD.n2527 9.3005
R4540 VDD.n227 VDD.n226 9.3005
R4541 VDD.n2541 VDD.n2540 9.3005
R4542 VDD.n2542 VDD.n225 9.3005
R4543 VDD.n2544 VDD.n2543 9.3005
R4544 VDD.n214 VDD.n213 9.3005
R4545 VDD.n2557 VDD.n2556 9.3005
R4546 VDD.n2558 VDD.n212 9.3005
R4547 VDD.n2560 VDD.n2559 9.3005
R4548 VDD.n203 VDD.n202 9.3005
R4549 VDD.n2573 VDD.n2572 9.3005
R4550 VDD.n2574 VDD.n201 9.3005
R4551 VDD.n2576 VDD.n2575 9.3005
R4552 VDD.n191 VDD.n190 9.3005
R4553 VDD.n2589 VDD.n2588 9.3005
R4554 VDD.n2590 VDD.n189 9.3005
R4555 VDD.n2595 VDD.n2591 9.3005
R4556 VDD.n2594 VDD.n2593 9.3005
R4557 VDD.n2592 VDD.n177 9.3005
R4558 VDD.n2608 VDD.n178 9.3005
R4559 VDD.n2609 VDD.n176 9.3005
R4560 VDD.n2611 VDD.n2610 9.3005
R4561 VDD.n2612 VDD.n175 9.3005
R4562 VDD.n2615 VDD.n2613 9.3005
R4563 VDD.n2616 VDD.n174 9.3005
R4564 VDD.n2618 VDD.n2617 9.3005
R4565 VDD.n2619 VDD.n173 9.3005
R4566 VDD.n2622 VDD.n2620 9.3005
R4567 VDD.n2623 VDD.n172 9.3005
R4568 VDD.n2625 VDD.n2624 9.3005
R4569 VDD.n2626 VDD.n171 9.3005
R4570 VDD.n2629 VDD.n2627 9.3005
R4571 VDD.n2630 VDD.n170 9.3005
R4572 VDD.n2632 VDD.n2631 9.3005
R4573 VDD.n2633 VDD.n169 9.3005
R4574 VDD.n2636 VDD.n2634 9.3005
R4575 VDD.n2637 VDD.n168 9.3005
R4576 VDD.n2639 VDD.n2638 9.3005
R4577 VDD.n2640 VDD.n167 9.3005
R4578 VDD.n2643 VDD.n2641 9.3005
R4579 VDD.n2644 VDD.n166 9.3005
R4580 VDD.n2646 VDD.n2645 9.3005
R4581 VDD.n2647 VDD.n165 9.3005
R4582 VDD.n2650 VDD.n2648 9.3005
R4583 VDD.n2651 VDD.n164 9.3005
R4584 VDD.n2653 VDD.n2652 9.3005
R4585 VDD.n2654 VDD.n163 9.3005
R4586 VDD.n2657 VDD.n2655 9.3005
R4587 VDD.n2658 VDD.n162 9.3005
R4588 VDD.n2660 VDD.n2659 9.3005
R4589 VDD.n2661 VDD.n161 9.3005
R4590 VDD.n2664 VDD.n2662 9.3005
R4591 VDD.n2665 VDD.n160 9.3005
R4592 VDD.n2667 VDD.n2666 9.3005
R4593 VDD.n2477 VDD.n2476 9.3005
R4594 VDD.n2438 VDD.n2437 9.3005
R4595 VDD.n2439 VDD.n2427 9.3005
R4596 VDD.n2440 VDD.n2426 9.3005
R4597 VDD.n2425 VDD.n2423 9.3005
R4598 VDD.n2446 VDD.n2422 9.3005
R4599 VDD.n2447 VDD.n2421 9.3005
R4600 VDD.n2448 VDD.n2420 9.3005
R4601 VDD.n2419 VDD.n2417 9.3005
R4602 VDD.n2454 VDD.n2416 9.3005
R4603 VDD.n2457 VDD.n2412 9.3005
R4604 VDD.n2411 VDD.n2409 9.3005
R4605 VDD.n2462 VDD.n2408 9.3005
R4606 VDD.n2463 VDD.n2407 9.3005
R4607 VDD.n2406 VDD.n2404 9.3005
R4608 VDD.n2468 VDD.n2403 9.3005
R4609 VDD.n2470 VDD.n2469 9.3005
R4610 VDD.n2456 VDD.n2413 9.3005
R4611 VDD.n2436 VDD.n2435 9.3005
R4612 VDD.n2430 VDD.n274 9.3005
R4613 VDD.n269 VDD.n268 9.3005
R4614 VDD.n2485 VDD.n2484 9.3005
R4615 VDD.n2486 VDD.n267 9.3005
R4616 VDD.n2488 VDD.n2487 9.3005
R4617 VDD.n257 VDD.n256 9.3005
R4618 VDD.n2501 VDD.n2500 9.3005
R4619 VDD.n2502 VDD.n255 9.3005
R4620 VDD.n2504 VDD.n2503 9.3005
R4621 VDD.n245 VDD.n244 9.3005
R4622 VDD.n2517 VDD.n2516 9.3005
R4623 VDD.n2518 VDD.n243 9.3005
R4624 VDD.n2520 VDD.n2519 9.3005
R4625 VDD.n233 VDD.n232 9.3005
R4626 VDD.n2533 VDD.n2532 9.3005
R4627 VDD.n2534 VDD.n231 9.3005
R4628 VDD.n2536 VDD.n2535 9.3005
R4629 VDD.n221 VDD.n220 9.3005
R4630 VDD.n2549 VDD.n2548 9.3005
R4631 VDD.n2550 VDD.n219 9.3005
R4632 VDD.n2552 VDD.n2551 9.3005
R4633 VDD.n209 VDD.n208 9.3005
R4634 VDD.n2565 VDD.n2564 9.3005
R4635 VDD.n2566 VDD.n207 9.3005
R4636 VDD.n2568 VDD.n2567 9.3005
R4637 VDD.n197 VDD.n196 9.3005
R4638 VDD.n2581 VDD.n2580 9.3005
R4639 VDD.n2582 VDD.n195 9.3005
R4640 VDD.n2584 VDD.n2583 9.3005
R4641 VDD.n184 VDD.n183 9.3005
R4642 VDD.n2600 VDD.n2599 9.3005
R4643 VDD.n2601 VDD.n182 9.3005
R4644 VDD.n2603 VDD.n2602 9.3005
R4645 VDD.n37 VDD.n35 9.3005
R4646 VDD.n2779 VDD.n2778 9.3005
R4647 VDD.n38 VDD.n36 9.3005
R4648 VDD.n2772 VDD.n46 9.3005
R4649 VDD.n2771 VDD.n47 9.3005
R4650 VDD.n2770 VDD.n48 9.3005
R4651 VDD.n56 VDD.n49 9.3005
R4652 VDD.n2764 VDD.n57 9.3005
R4653 VDD.n2763 VDD.n58 9.3005
R4654 VDD.n2762 VDD.n59 9.3005
R4655 VDD.n67 VDD.n60 9.3005
R4656 VDD.n2756 VDD.n68 9.3005
R4657 VDD.n2755 VDD.n69 9.3005
R4658 VDD.n2754 VDD.n70 9.3005
R4659 VDD.n78 VDD.n71 9.3005
R4660 VDD.n2748 VDD.n79 9.3005
R4661 VDD.n2747 VDD.n80 9.3005
R4662 VDD.n2746 VDD.n81 9.3005
R4663 VDD.n89 VDD.n82 9.3005
R4664 VDD.n2740 VDD.n90 9.3005
R4665 VDD.n2739 VDD.n91 9.3005
R4666 VDD.n2738 VDD.n92 9.3005
R4667 VDD.n100 VDD.n93 9.3005
R4668 VDD.n2732 VDD.n101 9.3005
R4669 VDD.n2731 VDD.n102 9.3005
R4670 VDD.n2730 VDD.n103 9.3005
R4671 VDD.n110 VDD.n104 9.3005
R4672 VDD.n2724 VDD.n111 9.3005
R4673 VDD.n2723 VDD.n112 9.3005
R4674 VDD.n2722 VDD.n113 9.3005
R4675 VDD.n122 VDD.n114 9.3005
R4676 VDD.n2716 VDD.n123 9.3005
R4677 VDD.n2715 VDD.n124 9.3005
R4678 VDD.n2714 VDD.n125 9.3005
R4679 VDD.n140 VDD.n126 9.3005
R4680 VDD.n2472 VDD.n2471 9.3005
R4681 VDD.n1123 VDD.n1122 9.3005
R4682 VDD.n786 VDD.n785 9.3005
R4683 VDD.n1136 VDD.n1135 9.3005
R4684 VDD.n1137 VDD.n784 9.3005
R4685 VDD.n1139 VDD.n1138 9.3005
R4686 VDD.n774 VDD.n773 9.3005
R4687 VDD.n1152 VDD.n1151 9.3005
R4688 VDD.n1153 VDD.n772 9.3005
R4689 VDD.n1155 VDD.n1154 9.3005
R4690 VDD.n762 VDD.n761 9.3005
R4691 VDD.n1169 VDD.n1168 9.3005
R4692 VDD.n1170 VDD.n760 9.3005
R4693 VDD.n1172 VDD.n1171 9.3005
R4694 VDD.n751 VDD.n750 9.3005
R4695 VDD.n1185 VDD.n1184 9.3005
R4696 VDD.n1186 VDD.n749 9.3005
R4697 VDD.n1188 VDD.n1187 9.3005
R4698 VDD.n739 VDD.n738 9.3005
R4699 VDD.n1201 VDD.n1200 9.3005
R4700 VDD.n1202 VDD.n737 9.3005
R4701 VDD.n1204 VDD.n1203 9.3005
R4702 VDD.n727 VDD.n726 9.3005
R4703 VDD.n1217 VDD.n1216 9.3005
R4704 VDD.n1218 VDD.n725 9.3005
R4705 VDD.n1220 VDD.n1219 9.3005
R4706 VDD.n715 VDD.n714 9.3005
R4707 VDD.n1233 VDD.n1232 9.3005
R4708 VDD.n1234 VDD.n713 9.3005
R4709 VDD.n1236 VDD.n1235 9.3005
R4710 VDD.n703 VDD.n702 9.3005
R4711 VDD.n1250 VDD.n1249 9.3005
R4712 VDD.n1251 VDD.n700 9.3005
R4713 VDD.n1308 VDD.n1307 9.3005
R4714 VDD.n1306 VDD.n701 9.3005
R4715 VDD.n1303 VDD.n1252 9.3005
R4716 VDD.n1302 VDD.n1301 9.3005
R4717 VDD.n1300 VDD.n1256 9.3005
R4718 VDD.n1299 VDD.n1298 9.3005
R4719 VDD.n1297 VDD.n1257 9.3005
R4720 VDD.n1296 VDD.n1295 9.3005
R4721 VDD.n1294 VDD.n1262 9.3005
R4722 VDD.n1293 VDD.n1292 9.3005
R4723 VDD.n1291 VDD.n1263 9.3005
R4724 VDD.n1290 VDD.n1289 9.3005
R4725 VDD.n1288 VDD.n1271 9.3005
R4726 VDD.n1287 VDD.n1286 9.3005
R4727 VDD.n1285 VDD.n1272 9.3005
R4728 VDD.n1284 VDD.n1283 9.3005
R4729 VDD.n1282 VDD.n1277 9.3005
R4730 VDD.n1281 VDD.n1280 9.3005
R4731 VDD.n693 VDD.n692 9.3005
R4732 VDD.n1316 VDD.n1315 9.3005
R4733 VDD.n1305 VDD.n1304 9.3005
R4734 VDD.n886 VDD.n885 9.3005
R4735 VDD.n977 VDD.n976 9.3005
R4736 VDD.n978 VDD.n884 9.3005
R4737 VDD.n980 VDD.n979 9.3005
R4738 VDD.n874 VDD.n873 9.3005
R4739 VDD.n993 VDD.n992 9.3005
R4740 VDD.n994 VDD.n872 9.3005
R4741 VDD.n996 VDD.n995 9.3005
R4742 VDD.n862 VDD.n861 9.3005
R4743 VDD.n1009 VDD.n1008 9.3005
R4744 VDD.n1010 VDD.n860 9.3005
R4745 VDD.n1012 VDD.n1011 9.3005
R4746 VDD.n850 VDD.n849 9.3005
R4747 VDD.n1025 VDD.n1024 9.3005
R4748 VDD.n1026 VDD.n848 9.3005
R4749 VDD.n1028 VDD.n1027 9.3005
R4750 VDD.n838 VDD.n837 9.3005
R4751 VDD.n1041 VDD.n1040 9.3005
R4752 VDD.n1042 VDD.n836 9.3005
R4753 VDD.n1044 VDD.n1043 9.3005
R4754 VDD.n827 VDD.n826 9.3005
R4755 VDD.n1058 VDD.n1057 9.3005
R4756 VDD.n1059 VDD.n825 9.3005
R4757 VDD.n1061 VDD.n1060 9.3005
R4758 VDD.n815 VDD.n814 9.3005
R4759 VDD.n1074 VDD.n1073 9.3005
R4760 VDD.n1075 VDD.n813 9.3005
R4761 VDD.n1077 VDD.n1076 9.3005
R4762 VDD.n803 VDD.n802 9.3005
R4763 VDD.n1090 VDD.n1089 9.3005
R4764 VDD.n1091 VDD.n801 9.3005
R4765 VDD.n1093 VDD.n1092 9.3005
R4766 VDD.n792 VDD.n791 9.3005
R4767 VDD.n1128 VDD.n1127 9.3005
R4768 VDD.n1129 VDD.n790 9.3005
R4769 VDD.n1131 VDD.n1130 9.3005
R4770 VDD.n780 VDD.n779 9.3005
R4771 VDD.n1144 VDD.n1143 9.3005
R4772 VDD.n1145 VDD.n778 9.3005
R4773 VDD.n1147 VDD.n1146 9.3005
R4774 VDD.n768 VDD.n767 9.3005
R4775 VDD.n1160 VDD.n1159 9.3005
R4776 VDD.n1161 VDD.n766 9.3005
R4777 VDD.n1163 VDD.n1162 9.3005
R4778 VDD.n757 VDD.n756 9.3005
R4779 VDD.n1177 VDD.n1176 9.3005
R4780 VDD.n1178 VDD.n755 9.3005
R4781 VDD.n1180 VDD.n1179 9.3005
R4782 VDD.n745 VDD.n744 9.3005
R4783 VDD.n1193 VDD.n1192 9.3005
R4784 VDD.n1194 VDD.n743 9.3005
R4785 VDD.n1196 VDD.n1195 9.3005
R4786 VDD.n733 VDD.n732 9.3005
R4787 VDD.n1209 VDD.n1208 9.3005
R4788 VDD.n1210 VDD.n731 9.3005
R4789 VDD.n1212 VDD.n1211 9.3005
R4790 VDD.n721 VDD.n720 9.3005
R4791 VDD.n1225 VDD.n1224 9.3005
R4792 VDD.n1226 VDD.n719 9.3005
R4793 VDD.n1228 VDD.n1227 9.3005
R4794 VDD.n709 VDD.n708 9.3005
R4795 VDD.n1241 VDD.n1240 9.3005
R4796 VDD.n1242 VDD.n707 9.3005
R4797 VDD.n1245 VDD.n1244 9.3005
R4798 VDD.n1243 VDD.n695 9.3005
R4799 VDD.n1312 VDD.n694 9.3005
R4800 VDD.n1314 VDD.n1313 9.3005
R4801 VDD.n964 VDD.n963 9.3005
R4802 VDD.n959 VDD.n958 9.3005
R4803 VDD.n957 VDD.n900 9.3005
R4804 VDD.n956 VDD.n955 9.3005
R4805 VDD.n903 VDD.n902 9.3005
R4806 VDD.n946 VDD.n906 9.3005
R4807 VDD.n948 VDD.n947 9.3005
R4808 VDD.n945 VDD.n908 9.3005
R4809 VDD.n944 VDD.n943 9.3005
R4810 VDD.n910 VDD.n909 9.3005
R4811 VDD.n935 VDD.n912 9.3005
R4812 VDD.n934 VDD.n933 9.3005
R4813 VDD.n917 VDD.n916 9.3005
R4814 VDD.n927 VDD.n926 9.3005
R4815 VDD.n925 VDD.n919 9.3005
R4816 VDD.n924 VDD.n923 9.3005
R4817 VDD.n920 VDD.n891 9.3005
R4818 VDD.n937 VDD.n936 9.3005
R4819 VDD.n960 VDD.n895 9.3005
R4820 VDD.n962 VDD.n961 9.3005
R4821 VDD.n970 VDD.n890 9.3005
R4822 VDD.n972 VDD.n971 9.3005
R4823 VDD.n880 VDD.n879 9.3005
R4824 VDD.n985 VDD.n984 9.3005
R4825 VDD.n986 VDD.n878 9.3005
R4826 VDD.n988 VDD.n987 9.3005
R4827 VDD.n868 VDD.n867 9.3005
R4828 VDD.n1001 VDD.n1000 9.3005
R4829 VDD.n1002 VDD.n866 9.3005
R4830 VDD.n1004 VDD.n1003 9.3005
R4831 VDD.n856 VDD.n855 9.3005
R4832 VDD.n1017 VDD.n1016 9.3005
R4833 VDD.n1018 VDD.n854 9.3005
R4834 VDD.n1020 VDD.n1019 9.3005
R4835 VDD.n844 VDD.n843 9.3005
R4836 VDD.n1033 VDD.n1032 9.3005
R4837 VDD.n1034 VDD.n842 9.3005
R4838 VDD.n1036 VDD.n1035 9.3005
R4839 VDD.n832 VDD.n831 9.3005
R4840 VDD.n1050 VDD.n1049 9.3005
R4841 VDD.n1051 VDD.n830 9.3005
R4842 VDD.n1053 VDD.n1052 9.3005
R4843 VDD.n821 VDD.n820 9.3005
R4844 VDD.n1066 VDD.n1065 9.3005
R4845 VDD.n1067 VDD.n819 9.3005
R4846 VDD.n1069 VDD.n1068 9.3005
R4847 VDD.n809 VDD.n808 9.3005
R4848 VDD.n1082 VDD.n1081 9.3005
R4849 VDD.n1083 VDD.n807 9.3005
R4850 VDD.n1085 VDD.n1084 9.3005
R4851 VDD.n797 VDD.n796 9.3005
R4852 VDD.n1099 VDD.n1098 9.3005
R4853 VDD.n1100 VDD.n795 9.3005
R4854 VDD.n969 VDD.n968 9.3005
R4855 VDD.n1115 VDD.n1114 9.3005
R4856 VDD.n1106 VDD.n1105 9.3005
R4857 VDD.n990 VDD.t9 8.94329
R4858 VDD.t1 VDD.n711 8.94329
R4859 VDD.n2498 VDD.t20 8.94329
R4860 VDD.n116 VDD.t5 8.94329
R4861 VDD.n1095 VDD.t64 8.59934
R4862 VDD.n1125 VDD.t64 8.59934
R4863 VDD.n2606 VDD.t57 8.59934
R4864 VDD.n2776 VDD.t57 8.59934
R4865 VDD.n15 VDD.n14 8.27334
R4866 VDD.n2781 VDD.n2780 8.26888
R4867 VDD.n1121 VDD.n1120 8.26888
R4868 VDD.t9 VDD.n870 8.25539
R4869 VDD.n1230 VDD.t1 8.25539
R4870 VDD.t20 VDD.n253 8.25539
R4871 VDD.n2726 VDD.t5 8.25539
R4872 VDD.n32 VDD.n26 8.14595
R4873 VDD.n23 VDD.n17 8.14595
R4874 VDD.n1116 VDD.n1110 8.14595
R4875 VDD.n1107 VDD.n1101 8.14595
R4876 VDD.n1813 VDD.t109 8.08341
R4877 VDD.n1862 VDD.t100 8.08341
R4878 VDD.t80 VDD.n625 7.91143
R4879 VDD.n1712 VDD.t112 7.91143
R4880 VDD.n2063 VDD.t88 7.91143
R4881 VDD.n2254 VDD.t77 7.91143
R4882 VDD.n7 VDD.t99 7.66677
R4883 VDD.n7 VDD.t106 7.66677
R4884 VDD.n8 VDD.t95 7.66677
R4885 VDD.n8 VDD.t104 7.66677
R4886 VDD.n10 VDD.t87 7.66677
R4887 VDD.n10 VDD.t82 7.66677
R4888 VDD.n12 VDD.t101 7.66677
R4889 VDD.n12 VDD.t76 7.66677
R4890 VDD.n5 VDD.t79 7.66677
R4891 VDD.n5 VDD.t110 7.66677
R4892 VDD.n3 VDD.t97 7.66677
R4893 VDD.n3 VDD.t92 7.66677
R4894 VDD.n1 VDD.t114 7.66677
R4895 VDD.n1 VDD.t108 7.66677
R4896 VDD.n0 VDD.t90 7.66677
R4897 VDD.n0 VDD.t84 7.66677
R4898 VDD.n1646 VDD.t107 7.56748
R4899 VDD.t94 VDD.n359 7.56748
R4900 VDD.n30 VDD.n29 7.3702
R4901 VDD.n21 VDD.n20 7.3702
R4902 VDD.n1114 VDD.n1113 7.3702
R4903 VDD.n1105 VDD.n1104 7.3702
R4904 VDD.n1119 VDD.n1109 7.09102
R4905 VDD.t83 VDD.n666 6.87957
R4906 VDD.n2349 VDD.t98 6.87957
R4907 VDD.t85 VDD.n601 6.53562
R4908 VDD.n1688 VDD.t93 6.53562
R4909 VDD.t102 VDD.n401 6.53562
R4910 VDD.n2230 VDD.t111 6.53562
R4911 VDD.n915 VDD.n910 6.4005
R4912 VDD.n2455 VDD.n2454 6.4005
R4913 VDD.n2692 VDD.n2689 6.4005
R4914 VDD.n1292 VDD.n1266 6.4005
R4915 VDD.n2781 VDD.n34 6.2014
R4916 VDD.n1120 VDD.n1119 6.2014
R4917 VDD.n1622 VDD.t113 6.19167
R4918 VDD.t103 VDD.n335 6.19167
R4919 VDD.n1119 VDD.n1118 6.0436
R4920 VDD.n30 VDD.n26 5.81868
R4921 VDD.n21 VDD.n17 5.81868
R4922 VDD.n1114 VDD.n1110 5.81868
R4923 VDD.n1105 VDD.n1101 5.81868
R4924 VDD.n2364 VDD.n2363 5.77611
R4925 VDD.n2095 VDD.n1876 5.77611
R4926 VDD.n1822 VDD.n1821 5.77611
R4927 VDD.n1553 VDD.n1465 5.77611
R4928 VDD.n2307 VDD.n2306 5.77611
R4929 VDD.n1980 VDD.n1979 5.77611
R4930 VDD.n1765 VDD.n1764 5.77611
R4931 VDD.n1326 VDD.n1323 5.77611
R4932 VDD.n34 VDD.n24 5.75481
R4933 VDD.t113 VDD.n643 5.50376
R4934 VDD.n2272 VDD.t103 5.50376
R4935 VDD.n1664 VDD.t85 5.1598
R4936 VDD.t93 VDD.n577 5.1598
R4937 VDD.n2206 VDD.t102 5.1598
R4938 VDD.t111 VDD.n377 5.1598
R4939 VDD.n2365 VDD.n2364 4.83952
R4940 VDD.n1876 VDD.n1872 4.83952
R4941 VDD.n1823 VDD.n1822 4.83952
R4942 VDD.n1465 VDD.n1461 4.83952
R4943 VDD.n2308 VDD.n2307 4.83952
R4944 VDD.n1979 VDD.n1978 4.83952
R4945 VDD.n1766 VDD.n1765 4.83952
R4946 VDD.n1327 VDD.n1326 4.83952
R4947 VDD.n1598 VDD.t83 4.81585
R4948 VDD.t98 VDD.n306 4.81585
R4949 VDD.n34 VDD.n33 4.7074
R4950 VDD.t107 VDD.n619 4.12794
R4951 VDD.n2248 VDD.t94 4.12794
R4952 VDD.n1640 VDD.t80 3.78399
R4953 VDD.t112 VDD.n553 3.78399
R4954 VDD.n2182 VDD.t88 3.78399
R4955 VDD.t77 VDD.n353 3.78399
R4956 VDD.n514 VDD.t109 3.61201
R4957 VDD.n2140 VDD.t100 3.61201
R4958 VDD.n31 VDD.n27 3.32369
R4959 VDD.n22 VDD.n18 3.32369
R4960 VDD.n1115 VDD.n1111 3.32369
R4961 VDD.n1106 VDD.n1102 3.32369
R4962 VDD.n543 VDD.t78 2.2362
R4963 VDD.n2164 VDD.t75 2.2362
R4964 VDD.n1046 VDD.t70 1.72027
R4965 VDD.n1174 VDD.t59 1.72027
R4966 VDD.n217 VDD.t66 1.72027
R4967 VDD.n2752 VDD.t62 1.72027
R4968 VDD.n1120 VDD.n15 1.55291
R4969 VDD VDD.n2781 1.54508
R4970 VDD.n4 VDD.n2 1.49727
R4971 VDD.n11 VDD.n9 1.49727
R4972 VDD.n6 VDD.n4 1.19016
R4973 VDD.n13 VDD.n11 1.19016
R4974 VDD.n14 VDD.n6 0.957397
R4975 VDD.n14 VDD.n13 0.957397
R4976 VDD.n567 VDD.t91 0.860384
R4977 VDD.n2188 VDD.t86 0.860384
R4978 VDD.t96 VDD.n583 0.51643
R4979 VDD.n2212 VDD.t81 0.51643
R4980 VDD.n141 VDD.n140 0.428854
R4981 VDD.n2668 VDD.n2667 0.428854
R4982 VDD.n2477 VDD.n274 0.428854
R4983 VDD.n2471 VDD.n2470 0.428854
R4984 VDD.n1306 VDD.n1305 0.428854
R4985 VDD.n1315 VDD.n1314 0.428854
R4986 VDD.n963 VDD.n962 0.428854
R4987 VDD.n969 VDD.n891 0.428854
R4988 VDD.n937 VDD.n915 0.194439
R4989 VDD.n2456 VDD.n2455 0.194439
R4990 VDD.n2693 VDD.n2692 0.194439
R4991 VDD.n1266 VDD.n1262 0.194439
R4992 VDD.n2779 VDD.n36 0.152939
R4993 VDD.n46 VDD.n36 0.152939
R4994 VDD.n47 VDD.n46 0.152939
R4995 VDD.n48 VDD.n47 0.152939
R4996 VDD.n56 VDD.n48 0.152939
R4997 VDD.n57 VDD.n56 0.152939
R4998 VDD.n58 VDD.n57 0.152939
R4999 VDD.n59 VDD.n58 0.152939
R5000 VDD.n67 VDD.n59 0.152939
R5001 VDD.n68 VDD.n67 0.152939
R5002 VDD.n69 VDD.n68 0.152939
R5003 VDD.n70 VDD.n69 0.152939
R5004 VDD.n78 VDD.n70 0.152939
R5005 VDD.n79 VDD.n78 0.152939
R5006 VDD.n80 VDD.n79 0.152939
R5007 VDD.n81 VDD.n80 0.152939
R5008 VDD.n89 VDD.n81 0.152939
R5009 VDD.n90 VDD.n89 0.152939
R5010 VDD.n91 VDD.n90 0.152939
R5011 VDD.n92 VDD.n91 0.152939
R5012 VDD.n100 VDD.n92 0.152939
R5013 VDD.n101 VDD.n100 0.152939
R5014 VDD.n102 VDD.n101 0.152939
R5015 VDD.n103 VDD.n102 0.152939
R5016 VDD.n110 VDD.n103 0.152939
R5017 VDD.n111 VDD.n110 0.152939
R5018 VDD.n112 VDD.n111 0.152939
R5019 VDD.n113 VDD.n112 0.152939
R5020 VDD.n122 VDD.n113 0.152939
R5021 VDD.n123 VDD.n122 0.152939
R5022 VDD.n124 VDD.n123 0.152939
R5023 VDD.n125 VDD.n124 0.152939
R5024 VDD.n140 VDD.n125 0.152939
R5025 VDD.n2706 VDD.n141 0.152939
R5026 VDD.n2706 VDD.n2705 0.152939
R5027 VDD.n2705 VDD.n2704 0.152939
R5028 VDD.n2704 VDD.n143 0.152939
R5029 VDD.n144 VDD.n143 0.152939
R5030 VDD.n145 VDD.n144 0.152939
R5031 VDD.n146 VDD.n145 0.152939
R5032 VDD.n147 VDD.n146 0.152939
R5033 VDD.n148 VDD.n147 0.152939
R5034 VDD.n149 VDD.n148 0.152939
R5035 VDD.n150 VDD.n149 0.152939
R5036 VDD.n151 VDD.n150 0.152939
R5037 VDD.n152 VDD.n151 0.152939
R5038 VDD.n153 VDD.n152 0.152939
R5039 VDD.n154 VDD.n153 0.152939
R5040 VDD.n155 VDD.n154 0.152939
R5041 VDD.n2669 VDD.n155 0.152939
R5042 VDD.n2669 VDD.n2668 0.152939
R5043 VDD.n2478 VDD.n2477 0.152939
R5044 VDD.n2479 VDD.n2478 0.152939
R5045 VDD.n2479 VDD.n262 0.152939
R5046 VDD.n2493 VDD.n262 0.152939
R5047 VDD.n2494 VDD.n2493 0.152939
R5048 VDD.n2495 VDD.n2494 0.152939
R5049 VDD.n2495 VDD.n250 0.152939
R5050 VDD.n2509 VDD.n250 0.152939
R5051 VDD.n2510 VDD.n2509 0.152939
R5052 VDD.n2511 VDD.n2510 0.152939
R5053 VDD.n2511 VDD.n238 0.152939
R5054 VDD.n2525 VDD.n238 0.152939
R5055 VDD.n2526 VDD.n2525 0.152939
R5056 VDD.n2527 VDD.n2526 0.152939
R5057 VDD.n2527 VDD.n226 0.152939
R5058 VDD.n2541 VDD.n226 0.152939
R5059 VDD.n2542 VDD.n2541 0.152939
R5060 VDD.n2543 VDD.n2542 0.152939
R5061 VDD.n2543 VDD.n213 0.152939
R5062 VDD.n2557 VDD.n213 0.152939
R5063 VDD.n2558 VDD.n2557 0.152939
R5064 VDD.n2559 VDD.n2558 0.152939
R5065 VDD.n2559 VDD.n202 0.152939
R5066 VDD.n2573 VDD.n202 0.152939
R5067 VDD.n2574 VDD.n2573 0.152939
R5068 VDD.n2575 VDD.n2574 0.152939
R5069 VDD.n2575 VDD.n190 0.152939
R5070 VDD.n2589 VDD.n190 0.152939
R5071 VDD.n2590 VDD.n2589 0.152939
R5072 VDD.n2591 VDD.n2590 0.152939
R5073 VDD.n2593 VDD.n2591 0.152939
R5074 VDD.n2593 VDD.n2592 0.152939
R5075 VDD.n2592 VDD.n178 0.152939
R5076 VDD.n178 VDD.n176 0.152939
R5077 VDD.n2611 VDD.n176 0.152939
R5078 VDD.n2612 VDD.n2611 0.152939
R5079 VDD.n2613 VDD.n2612 0.152939
R5080 VDD.n2613 VDD.n174 0.152939
R5081 VDD.n2618 VDD.n174 0.152939
R5082 VDD.n2619 VDD.n2618 0.152939
R5083 VDD.n2620 VDD.n2619 0.152939
R5084 VDD.n2620 VDD.n172 0.152939
R5085 VDD.n2625 VDD.n172 0.152939
R5086 VDD.n2626 VDD.n2625 0.152939
R5087 VDD.n2627 VDD.n2626 0.152939
R5088 VDD.n2627 VDD.n170 0.152939
R5089 VDD.n2632 VDD.n170 0.152939
R5090 VDD.n2633 VDD.n2632 0.152939
R5091 VDD.n2634 VDD.n2633 0.152939
R5092 VDD.n2634 VDD.n168 0.152939
R5093 VDD.n2639 VDD.n168 0.152939
R5094 VDD.n2640 VDD.n2639 0.152939
R5095 VDD.n2641 VDD.n2640 0.152939
R5096 VDD.n2641 VDD.n166 0.152939
R5097 VDD.n2646 VDD.n166 0.152939
R5098 VDD.n2647 VDD.n2646 0.152939
R5099 VDD.n2648 VDD.n2647 0.152939
R5100 VDD.n2648 VDD.n164 0.152939
R5101 VDD.n2653 VDD.n164 0.152939
R5102 VDD.n2654 VDD.n2653 0.152939
R5103 VDD.n2655 VDD.n2654 0.152939
R5104 VDD.n2655 VDD.n162 0.152939
R5105 VDD.n2660 VDD.n162 0.152939
R5106 VDD.n2661 VDD.n2660 0.152939
R5107 VDD.n2662 VDD.n2661 0.152939
R5108 VDD.n2662 VDD.n160 0.152939
R5109 VDD.n2667 VDD.n160 0.152939
R5110 VDD.n2470 VDD.n2403 0.152939
R5111 VDD.n2406 VDD.n2403 0.152939
R5112 VDD.n2407 VDD.n2406 0.152939
R5113 VDD.n2408 VDD.n2407 0.152939
R5114 VDD.n2411 VDD.n2408 0.152939
R5115 VDD.n2412 VDD.n2411 0.152939
R5116 VDD.n2413 VDD.n2412 0.152939
R5117 VDD.n2416 VDD.n2413 0.152939
R5118 VDD.n2419 VDD.n2416 0.152939
R5119 VDD.n2420 VDD.n2419 0.152939
R5120 VDD.n2421 VDD.n2420 0.152939
R5121 VDD.n2422 VDD.n2421 0.152939
R5122 VDD.n2425 VDD.n2422 0.152939
R5123 VDD.n2426 VDD.n2425 0.152939
R5124 VDD.n2427 VDD.n2426 0.152939
R5125 VDD.n2437 VDD.n2427 0.152939
R5126 VDD.n2437 VDD.n2436 0.152939
R5127 VDD.n2436 VDD.n274 0.152939
R5128 VDD.n2471 VDD.n268 0.152939
R5129 VDD.n2485 VDD.n268 0.152939
R5130 VDD.n2486 VDD.n2485 0.152939
R5131 VDD.n2487 VDD.n2486 0.152939
R5132 VDD.n2487 VDD.n256 0.152939
R5133 VDD.n2501 VDD.n256 0.152939
R5134 VDD.n2502 VDD.n2501 0.152939
R5135 VDD.n2503 VDD.n2502 0.152939
R5136 VDD.n2503 VDD.n244 0.152939
R5137 VDD.n2517 VDD.n244 0.152939
R5138 VDD.n2518 VDD.n2517 0.152939
R5139 VDD.n2519 VDD.n2518 0.152939
R5140 VDD.n2519 VDD.n232 0.152939
R5141 VDD.n2533 VDD.n232 0.152939
R5142 VDD.n2534 VDD.n2533 0.152939
R5143 VDD.n2535 VDD.n2534 0.152939
R5144 VDD.n2535 VDD.n220 0.152939
R5145 VDD.n2549 VDD.n220 0.152939
R5146 VDD.n2550 VDD.n2549 0.152939
R5147 VDD.n2551 VDD.n2550 0.152939
R5148 VDD.n2551 VDD.n208 0.152939
R5149 VDD.n2565 VDD.n208 0.152939
R5150 VDD.n2566 VDD.n2565 0.152939
R5151 VDD.n2567 VDD.n2566 0.152939
R5152 VDD.n2567 VDD.n196 0.152939
R5153 VDD.n2581 VDD.n196 0.152939
R5154 VDD.n2582 VDD.n2581 0.152939
R5155 VDD.n2583 VDD.n2582 0.152939
R5156 VDD.n2583 VDD.n183 0.152939
R5157 VDD.n2600 VDD.n183 0.152939
R5158 VDD.n2601 VDD.n2600 0.152939
R5159 VDD.n2602 VDD.n2601 0.152939
R5160 VDD.n2602 VDD.n35 0.152939
R5161 VDD.n1122 VDD.n785 0.152939
R5162 VDD.n1136 VDD.n785 0.152939
R5163 VDD.n1137 VDD.n1136 0.152939
R5164 VDD.n1138 VDD.n1137 0.152939
R5165 VDD.n1138 VDD.n773 0.152939
R5166 VDD.n1152 VDD.n773 0.152939
R5167 VDD.n1153 VDD.n1152 0.152939
R5168 VDD.n1154 VDD.n1153 0.152939
R5169 VDD.n1154 VDD.n761 0.152939
R5170 VDD.n1169 VDD.n761 0.152939
R5171 VDD.n1170 VDD.n1169 0.152939
R5172 VDD.n1171 VDD.n1170 0.152939
R5173 VDD.n1171 VDD.n750 0.152939
R5174 VDD.n1185 VDD.n750 0.152939
R5175 VDD.n1186 VDD.n1185 0.152939
R5176 VDD.n1187 VDD.n1186 0.152939
R5177 VDD.n1187 VDD.n738 0.152939
R5178 VDD.n1201 VDD.n738 0.152939
R5179 VDD.n1202 VDD.n1201 0.152939
R5180 VDD.n1203 VDD.n1202 0.152939
R5181 VDD.n1203 VDD.n726 0.152939
R5182 VDD.n1217 VDD.n726 0.152939
R5183 VDD.n1218 VDD.n1217 0.152939
R5184 VDD.n1219 VDD.n1218 0.152939
R5185 VDD.n1219 VDD.n714 0.152939
R5186 VDD.n1233 VDD.n714 0.152939
R5187 VDD.n1234 VDD.n1233 0.152939
R5188 VDD.n1235 VDD.n1234 0.152939
R5189 VDD.n1235 VDD.n702 0.152939
R5190 VDD.n1250 VDD.n702 0.152939
R5191 VDD.n1251 VDD.n1250 0.152939
R5192 VDD.n1307 VDD.n1251 0.152939
R5193 VDD.n1307 VDD.n1306 0.152939
R5194 VDD.n1305 VDD.n1252 0.152939
R5195 VDD.n1301 VDD.n1252 0.152939
R5196 VDD.n1301 VDD.n1300 0.152939
R5197 VDD.n1300 VDD.n1299 0.152939
R5198 VDD.n1299 VDD.n1257 0.152939
R5199 VDD.n1295 VDD.n1257 0.152939
R5200 VDD.n1295 VDD.n1294 0.152939
R5201 VDD.n1294 VDD.n1293 0.152939
R5202 VDD.n1293 VDD.n1263 0.152939
R5203 VDD.n1289 VDD.n1263 0.152939
R5204 VDD.n1289 VDD.n1288 0.152939
R5205 VDD.n1288 VDD.n1287 0.152939
R5206 VDD.n1287 VDD.n1272 0.152939
R5207 VDD.n1283 VDD.n1272 0.152939
R5208 VDD.n1283 VDD.n1282 0.152939
R5209 VDD.n1282 VDD.n1281 0.152939
R5210 VDD.n1281 VDD.n693 0.152939
R5211 VDD.n1315 VDD.n693 0.152939
R5212 VDD.n963 VDD.n885 0.152939
R5213 VDD.n977 VDD.n885 0.152939
R5214 VDD.n978 VDD.n977 0.152939
R5215 VDD.n979 VDD.n978 0.152939
R5216 VDD.n979 VDD.n873 0.152939
R5217 VDD.n993 VDD.n873 0.152939
R5218 VDD.n994 VDD.n993 0.152939
R5219 VDD.n995 VDD.n994 0.152939
R5220 VDD.n995 VDD.n861 0.152939
R5221 VDD.n1009 VDD.n861 0.152939
R5222 VDD.n1010 VDD.n1009 0.152939
R5223 VDD.n1011 VDD.n1010 0.152939
R5224 VDD.n1011 VDD.n849 0.152939
R5225 VDD.n1025 VDD.n849 0.152939
R5226 VDD.n1026 VDD.n1025 0.152939
R5227 VDD.n1027 VDD.n1026 0.152939
R5228 VDD.n1027 VDD.n837 0.152939
R5229 VDD.n1041 VDD.n837 0.152939
R5230 VDD.n1042 VDD.n1041 0.152939
R5231 VDD.n1043 VDD.n1042 0.152939
R5232 VDD.n1043 VDD.n826 0.152939
R5233 VDD.n1058 VDD.n826 0.152939
R5234 VDD.n1059 VDD.n1058 0.152939
R5235 VDD.n1060 VDD.n1059 0.152939
R5236 VDD.n1060 VDD.n814 0.152939
R5237 VDD.n1074 VDD.n814 0.152939
R5238 VDD.n1075 VDD.n1074 0.152939
R5239 VDD.n1076 VDD.n1075 0.152939
R5240 VDD.n1076 VDD.n802 0.152939
R5241 VDD.n1090 VDD.n802 0.152939
R5242 VDD.n1091 VDD.n1090 0.152939
R5243 VDD.n1092 VDD.n1091 0.152939
R5244 VDD.n1092 VDD.n791 0.152939
R5245 VDD.n1128 VDD.n791 0.152939
R5246 VDD.n1129 VDD.n1128 0.152939
R5247 VDD.n1130 VDD.n1129 0.152939
R5248 VDD.n1130 VDD.n779 0.152939
R5249 VDD.n1144 VDD.n779 0.152939
R5250 VDD.n1145 VDD.n1144 0.152939
R5251 VDD.n1146 VDD.n1145 0.152939
R5252 VDD.n1146 VDD.n767 0.152939
R5253 VDD.n1160 VDD.n767 0.152939
R5254 VDD.n1161 VDD.n1160 0.152939
R5255 VDD.n1162 VDD.n1161 0.152939
R5256 VDD.n1162 VDD.n756 0.152939
R5257 VDD.n1177 VDD.n756 0.152939
R5258 VDD.n1178 VDD.n1177 0.152939
R5259 VDD.n1179 VDD.n1178 0.152939
R5260 VDD.n1179 VDD.n744 0.152939
R5261 VDD.n1193 VDD.n744 0.152939
R5262 VDD.n1194 VDD.n1193 0.152939
R5263 VDD.n1195 VDD.n1194 0.152939
R5264 VDD.n1195 VDD.n732 0.152939
R5265 VDD.n1209 VDD.n732 0.152939
R5266 VDD.n1210 VDD.n1209 0.152939
R5267 VDD.n1211 VDD.n1210 0.152939
R5268 VDD.n1211 VDD.n720 0.152939
R5269 VDD.n1225 VDD.n720 0.152939
R5270 VDD.n1226 VDD.n1225 0.152939
R5271 VDD.n1227 VDD.n1226 0.152939
R5272 VDD.n1227 VDD.n708 0.152939
R5273 VDD.n1241 VDD.n708 0.152939
R5274 VDD.n1242 VDD.n1241 0.152939
R5275 VDD.n1244 VDD.n1242 0.152939
R5276 VDD.n1244 VDD.n1243 0.152939
R5277 VDD.n1243 VDD.n694 0.152939
R5278 VDD.n1314 VDD.n694 0.152939
R5279 VDD.n924 VDD.n891 0.152939
R5280 VDD.n925 VDD.n924 0.152939
R5281 VDD.n926 VDD.n925 0.152939
R5282 VDD.n926 VDD.n916 0.152939
R5283 VDD.n934 VDD.n916 0.152939
R5284 VDD.n935 VDD.n934 0.152939
R5285 VDD.n936 VDD.n935 0.152939
R5286 VDD.n936 VDD.n909 0.152939
R5287 VDD.n944 VDD.n909 0.152939
R5288 VDD.n945 VDD.n944 0.152939
R5289 VDD.n947 VDD.n945 0.152939
R5290 VDD.n947 VDD.n946 0.152939
R5291 VDD.n946 VDD.n902 0.152939
R5292 VDD.n956 VDD.n902 0.152939
R5293 VDD.n957 VDD.n956 0.152939
R5294 VDD.n958 VDD.n957 0.152939
R5295 VDD.n958 VDD.n895 0.152939
R5296 VDD.n962 VDD.n895 0.152939
R5297 VDD.n970 VDD.n969 0.152939
R5298 VDD.n971 VDD.n970 0.152939
R5299 VDD.n971 VDD.n879 0.152939
R5300 VDD.n985 VDD.n879 0.152939
R5301 VDD.n986 VDD.n985 0.152939
R5302 VDD.n987 VDD.n986 0.152939
R5303 VDD.n987 VDD.n867 0.152939
R5304 VDD.n1001 VDD.n867 0.152939
R5305 VDD.n1002 VDD.n1001 0.152939
R5306 VDD.n1003 VDD.n1002 0.152939
R5307 VDD.n1003 VDD.n855 0.152939
R5308 VDD.n1017 VDD.n855 0.152939
R5309 VDD.n1018 VDD.n1017 0.152939
R5310 VDD.n1019 VDD.n1018 0.152939
R5311 VDD.n1019 VDD.n843 0.152939
R5312 VDD.n1033 VDD.n843 0.152939
R5313 VDD.n1034 VDD.n1033 0.152939
R5314 VDD.n1035 VDD.n1034 0.152939
R5315 VDD.n1035 VDD.n831 0.152939
R5316 VDD.n1050 VDD.n831 0.152939
R5317 VDD.n1051 VDD.n1050 0.152939
R5318 VDD.n1052 VDD.n1051 0.152939
R5319 VDD.n1052 VDD.n820 0.152939
R5320 VDD.n1066 VDD.n820 0.152939
R5321 VDD.n1067 VDD.n1066 0.152939
R5322 VDD.n1068 VDD.n1067 0.152939
R5323 VDD.n1068 VDD.n808 0.152939
R5324 VDD.n1082 VDD.n808 0.152939
R5325 VDD.n1083 VDD.n1082 0.152939
R5326 VDD.n1084 VDD.n1083 0.152939
R5327 VDD.n1084 VDD.n796 0.152939
R5328 VDD.n1099 VDD.n796 0.152939
R5329 VDD.n1100 VDD.n1099 0.152939
R5330 VDD.n2780 VDD.n35 0.0695946
R5331 VDD.n2780 VDD.n2779 0.0695946
R5332 VDD.n1122 VDD.n1121 0.0695946
R5333 VDD.n1121 VDD.n1100 0.0695946
R5334 VDD VDD.n15 0.00833333
R5335 DIFFPAIR_BIAS.n14 DIFFPAIR_BIAS.n0 289.615
R5336 DIFFPAIR_BIAS.n33 DIFFPAIR_BIAS.n19 289.615
R5337 DIFFPAIR_BIAS.n53 DIFFPAIR_BIAS.n39 289.615
R5338 DIFFPAIR_BIAS.n15 DIFFPAIR_BIAS.n14 185
R5339 DIFFPAIR_BIAS.n13 DIFFPAIR_BIAS.n12 185
R5340 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.n3 185
R5341 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.n6 185
R5342 DIFFPAIR_BIAS.n34 DIFFPAIR_BIAS.n33 185
R5343 DIFFPAIR_BIAS.n32 DIFFPAIR_BIAS.n31 185
R5344 DIFFPAIR_BIAS.n23 DIFFPAIR_BIAS.n22 185
R5345 DIFFPAIR_BIAS.n26 DIFFPAIR_BIAS.n25 185
R5346 DIFFPAIR_BIAS.n54 DIFFPAIR_BIAS.n53 185
R5347 DIFFPAIR_BIAS.n52 DIFFPAIR_BIAS.n51 185
R5348 DIFFPAIR_BIAS.n43 DIFFPAIR_BIAS.n42 185
R5349 DIFFPAIR_BIAS.n46 DIFFPAIR_BIAS.n45 185
R5350 DIFFPAIR_BIAS.t5 DIFFPAIR_BIAS.n5 147.888
R5351 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.n24 147.888
R5352 DIFFPAIR_BIAS.t3 DIFFPAIR_BIAS.n44 147.888
R5353 DIFFPAIR_BIAS.n64 DIFFPAIR_BIAS.t6 106.936
R5354 DIFFPAIR_BIAS.n63 DIFFPAIR_BIAS.t7 105.168
R5355 DIFFPAIR_BIAS.n62 DIFFPAIR_BIAS.t8 105.168
R5356 DIFFPAIR_BIAS.n14 DIFFPAIR_BIAS.n13 104.615
R5357 DIFFPAIR_BIAS.n13 DIFFPAIR_BIAS.n3 104.615
R5358 DIFFPAIR_BIAS.n6 DIFFPAIR_BIAS.n3 104.615
R5359 DIFFPAIR_BIAS.n33 DIFFPAIR_BIAS.n32 104.615
R5360 DIFFPAIR_BIAS.n32 DIFFPAIR_BIAS.n22 104.615
R5361 DIFFPAIR_BIAS.n25 DIFFPAIR_BIAS.n22 104.615
R5362 DIFFPAIR_BIAS.n53 DIFFPAIR_BIAS.n52 104.615
R5363 DIFFPAIR_BIAS.n52 DIFFPAIR_BIAS.n42 104.615
R5364 DIFFPAIR_BIAS.n45 DIFFPAIR_BIAS.n42 104.615
R5365 DIFFPAIR_BIAS.n38 DIFFPAIR_BIAS.n18 99.4403
R5366 DIFFPAIR_BIAS.n38 DIFFPAIR_BIAS.n37 98.1641
R5367 DIFFPAIR_BIAS.n58 DIFFPAIR_BIAS.n57 98.1641
R5368 DIFFPAIR_BIAS.n59 DIFFPAIR_BIAS.t4 80.4932
R5369 DIFFPAIR_BIAS.n59 DIFFPAIR_BIAS.t0 77.9396
R5370 DIFFPAIR_BIAS.n60 DIFFPAIR_BIAS.t2 77.9396
R5371 DIFFPAIR_BIAS.n6 DIFFPAIR_BIAS.t5 52.3082
R5372 DIFFPAIR_BIAS.n25 DIFFPAIR_BIAS.t1 52.3082
R5373 DIFFPAIR_BIAS.n45 DIFFPAIR_BIAS.t3 52.3082
R5374 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.n5 15.6496
R5375 DIFFPAIR_BIAS.n26 DIFFPAIR_BIAS.n24 15.6496
R5376 DIFFPAIR_BIAS.n46 DIFFPAIR_BIAS.n44 15.6496
R5377 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.n4 12.8005
R5378 DIFFPAIR_BIAS.n27 DIFFPAIR_BIAS.n23 12.8005
R5379 DIFFPAIR_BIAS.n47 DIFFPAIR_BIAS.n43 12.8005
R5380 DIFFPAIR_BIAS.n12 DIFFPAIR_BIAS.n11 12.0247
R5381 DIFFPAIR_BIAS.n31 DIFFPAIR_BIAS.n30 12.0247
R5382 DIFFPAIR_BIAS.n51 DIFFPAIR_BIAS.n50 12.0247
R5383 DIFFPAIR_BIAS.n15 DIFFPAIR_BIAS.n2 11.249
R5384 DIFFPAIR_BIAS.n34 DIFFPAIR_BIAS.n21 11.249
R5385 DIFFPAIR_BIAS.n54 DIFFPAIR_BIAS.n41 11.249
R5386 DIFFPAIR_BIAS.n16 DIFFPAIR_BIAS.n0 10.4732
R5387 DIFFPAIR_BIAS.n35 DIFFPAIR_BIAS.n19 10.4732
R5388 DIFFPAIR_BIAS.n55 DIFFPAIR_BIAS.n39 10.4732
R5389 DIFFPAIR_BIAS.n18 DIFFPAIR_BIAS.n17 9.45567
R5390 DIFFPAIR_BIAS.n37 DIFFPAIR_BIAS.n36 9.45567
R5391 DIFFPAIR_BIAS.n57 DIFFPAIR_BIAS.n56 9.45567
R5392 DIFFPAIR_BIAS.n17 DIFFPAIR_BIAS.n16 9.3005
R5393 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.n1 9.3005
R5394 DIFFPAIR_BIAS.n11 DIFFPAIR_BIAS.n10 9.3005
R5395 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.n8 9.3005
R5396 DIFFPAIR_BIAS.n36 DIFFPAIR_BIAS.n35 9.3005
R5397 DIFFPAIR_BIAS.n21 DIFFPAIR_BIAS.n20 9.3005
R5398 DIFFPAIR_BIAS.n30 DIFFPAIR_BIAS.n29 9.3005
R5399 DIFFPAIR_BIAS.n28 DIFFPAIR_BIAS.n27 9.3005
R5400 DIFFPAIR_BIAS.n56 DIFFPAIR_BIAS.n55 9.3005
R5401 DIFFPAIR_BIAS.n41 DIFFPAIR_BIAS.n40 9.3005
R5402 DIFFPAIR_BIAS.n50 DIFFPAIR_BIAS.n49 9.3005
R5403 DIFFPAIR_BIAS.n48 DIFFPAIR_BIAS.n47 9.3005
R5404 DIFFPAIR_BIAS.n61 DIFFPAIR_BIAS.n60 5.67907
R5405 DIFFPAIR_BIAS.n61 DIFFPAIR_BIAS.n58 4.51702
R5406 DIFFPAIR_BIAS.n62 DIFFPAIR_BIAS.n61 4.44014
R5407 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.n5 4.40546
R5408 DIFFPAIR_BIAS.n28 DIFFPAIR_BIAS.n24 4.40546
R5409 DIFFPAIR_BIAS.n48 DIFFPAIR_BIAS.n44 4.40546
R5410 DIFFPAIR_BIAS.n18 DIFFPAIR_BIAS.n0 3.49141
R5411 DIFFPAIR_BIAS.n37 DIFFPAIR_BIAS.n19 3.49141
R5412 DIFFPAIR_BIAS.n57 DIFFPAIR_BIAS.n39 3.49141
R5413 DIFFPAIR_BIAS.n16 DIFFPAIR_BIAS.n15 2.71565
R5414 DIFFPAIR_BIAS.n35 DIFFPAIR_BIAS.n34 2.71565
R5415 DIFFPAIR_BIAS.n55 DIFFPAIR_BIAS.n54 2.71565
R5416 DIFFPAIR_BIAS.n60 DIFFPAIR_BIAS.n59 2.55507
R5417 DIFFPAIR_BIAS.n63 DIFFPAIR_BIAS.n62 2.55497
R5418 DIFFPAIR_BIAS.n12 DIFFPAIR_BIAS.n2 1.93989
R5419 DIFFPAIR_BIAS.n31 DIFFPAIR_BIAS.n21 1.93989
R5420 DIFFPAIR_BIAS.n51 DIFFPAIR_BIAS.n41 1.93989
R5421 DIFFPAIR_BIAS.n58 DIFFPAIR_BIAS.n38 1.27666
R5422 DIFFPAIR_BIAS.n11 DIFFPAIR_BIAS.n4 1.16414
R5423 DIFFPAIR_BIAS.n30 DIFFPAIR_BIAS.n23 1.16414
R5424 DIFFPAIR_BIAS.n50 DIFFPAIR_BIAS.n43 1.16414
R5425 DIFFPAIR_BIAS DIFFPAIR_BIAS.n64 0.6855
R5426 DIFFPAIR_BIAS.n64 DIFFPAIR_BIAS.n63 0.494303
R5427 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.n7 0.388379
R5428 DIFFPAIR_BIAS.n27 DIFFPAIR_BIAS.n26 0.388379
R5429 DIFFPAIR_BIAS.n47 DIFFPAIR_BIAS.n46 0.388379
R5430 DIFFPAIR_BIAS.n17 DIFFPAIR_BIAS.n1 0.155672
R5431 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.n1 0.155672
R5432 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.n9 0.155672
R5433 DIFFPAIR_BIAS.n36 DIFFPAIR_BIAS.n20 0.155672
R5434 DIFFPAIR_BIAS.n29 DIFFPAIR_BIAS.n20 0.155672
R5435 DIFFPAIR_BIAS.n29 DIFFPAIR_BIAS.n28 0.155672
R5436 DIFFPAIR_BIAS.n56 DIFFPAIR_BIAS.n40 0.155672
R5437 DIFFPAIR_BIAS.n49 DIFFPAIR_BIAS.n40 0.155672
R5438 DIFFPAIR_BIAS.n49 DIFFPAIR_BIAS.n48 0.155672
R5439 GND.n5930 GND.n553 2335.17
R5440 GND.n5134 GND.n1076 1694.82
R5441 GND.n5241 GND.n968 819.232
R5442 GND.n5931 GND.n554 819.232
R5443 GND.n6071 GND.n469 819.232
R5444 GND.n5127 GND.n1077 819.232
R5445 GND.n6255 GND.n290 795.207
R5446 GND.n6160 GND.n385 795.207
R5447 GND.n4588 GND.n1589 795.207
R5448 GND.n4686 GND.n1599 795.207
R5449 GND.n4952 GND.n1296 795.207
R5450 GND.n4954 GND.n1289 795.207
R5451 GND.n3487 GND.n1163 795.207
R5452 GND.n5043 GND.n1167 795.207
R5453 GND.n4403 GND.n285 780.793
R5454 GND.n4430 GND.n386 780.793
R5455 GND.n2031 GND.n1665 780.793
R5456 GND.n4586 GND.n1667 780.793
R5457 GND.n1408 GND.n1294 780.793
R5458 GND.n4834 GND.n1291 780.793
R5459 GND.n3522 GND.n1164 780.793
R5460 GND.n3496 GND.n1166 780.793
R5461 GND.n4824 GND.n1465 771.183
R5462 GND.n4698 GND.n1553 771.183
R5463 GND.n2039 GND.n1556 771.183
R5464 GND.n4828 GND.n1446 771.183
R5465 GND.n5242 GND.n5241 585
R5466 GND.n5241 GND.n5240 585
R5467 GND.n972 GND.n971 585
R5468 GND.n5239 GND.n972 585
R5469 GND.n5237 GND.n5236 585
R5470 GND.n5238 GND.n5237 585
R5471 GND.n5235 GND.n974 585
R5472 GND.n974 GND.n973 585
R5473 GND.n5234 GND.n5233 585
R5474 GND.n5233 GND.n5232 585
R5475 GND.n979 GND.n978 585
R5476 GND.n5231 GND.n979 585
R5477 GND.n5229 GND.n5228 585
R5478 GND.n5230 GND.n5229 585
R5479 GND.n5227 GND.n981 585
R5480 GND.n981 GND.n980 585
R5481 GND.n5226 GND.n5225 585
R5482 GND.n5225 GND.n5224 585
R5483 GND.n987 GND.n986 585
R5484 GND.n5223 GND.n987 585
R5485 GND.n5221 GND.n5220 585
R5486 GND.n5222 GND.n5221 585
R5487 GND.n5219 GND.n989 585
R5488 GND.n989 GND.n988 585
R5489 GND.n5218 GND.n5217 585
R5490 GND.n5217 GND.n5216 585
R5491 GND.n995 GND.n994 585
R5492 GND.n5215 GND.n995 585
R5493 GND.n5213 GND.n5212 585
R5494 GND.n5214 GND.n5213 585
R5495 GND.n5211 GND.n997 585
R5496 GND.n997 GND.n996 585
R5497 GND.n5210 GND.n5209 585
R5498 GND.n5209 GND.n5208 585
R5499 GND.n1003 GND.n1002 585
R5500 GND.n5207 GND.n1003 585
R5501 GND.n5205 GND.n5204 585
R5502 GND.n5206 GND.n5205 585
R5503 GND.n5203 GND.n1005 585
R5504 GND.n1005 GND.n1004 585
R5505 GND.n5202 GND.n5201 585
R5506 GND.n5201 GND.n5200 585
R5507 GND.n1011 GND.n1010 585
R5508 GND.n5199 GND.n1011 585
R5509 GND.n5197 GND.n5196 585
R5510 GND.n5198 GND.n5197 585
R5511 GND.n5195 GND.n1013 585
R5512 GND.n1013 GND.n1012 585
R5513 GND.n5194 GND.n5193 585
R5514 GND.n5193 GND.n5192 585
R5515 GND.n1019 GND.n1018 585
R5516 GND.n5191 GND.n1019 585
R5517 GND.n5189 GND.n5188 585
R5518 GND.n5190 GND.n5189 585
R5519 GND.n5187 GND.n1021 585
R5520 GND.n1021 GND.n1020 585
R5521 GND.n5186 GND.n5185 585
R5522 GND.n5185 GND.n5184 585
R5523 GND.n1027 GND.n1026 585
R5524 GND.n5183 GND.n1027 585
R5525 GND.n5181 GND.n5180 585
R5526 GND.n5182 GND.n5181 585
R5527 GND.n5179 GND.n1029 585
R5528 GND.n1029 GND.n1028 585
R5529 GND.n5178 GND.n5177 585
R5530 GND.n5177 GND.n5176 585
R5531 GND.n1035 GND.n1034 585
R5532 GND.n5175 GND.n1035 585
R5533 GND.n5173 GND.n5172 585
R5534 GND.n5174 GND.n5173 585
R5535 GND.n5171 GND.n1037 585
R5536 GND.n1037 GND.n1036 585
R5537 GND.n5170 GND.n5169 585
R5538 GND.n5169 GND.n5168 585
R5539 GND.n1043 GND.n1042 585
R5540 GND.n5167 GND.n1043 585
R5541 GND.n5165 GND.n5164 585
R5542 GND.n5166 GND.n5165 585
R5543 GND.n5163 GND.n1045 585
R5544 GND.n1045 GND.n1044 585
R5545 GND.n5162 GND.n5161 585
R5546 GND.n5161 GND.n5160 585
R5547 GND.n1051 GND.n1050 585
R5548 GND.n5159 GND.n1051 585
R5549 GND.n5157 GND.n5156 585
R5550 GND.n5158 GND.n5157 585
R5551 GND.n5155 GND.n1053 585
R5552 GND.n1053 GND.n1052 585
R5553 GND.n5154 GND.n5153 585
R5554 GND.n5153 GND.n5152 585
R5555 GND.n1059 GND.n1058 585
R5556 GND.n5151 GND.n1059 585
R5557 GND.n5149 GND.n5148 585
R5558 GND.n5150 GND.n5149 585
R5559 GND.n5147 GND.n1061 585
R5560 GND.n1061 GND.n1060 585
R5561 GND.n5146 GND.n5145 585
R5562 GND.n5145 GND.n5144 585
R5563 GND.n1067 GND.n1066 585
R5564 GND.n5143 GND.n1067 585
R5565 GND.n5141 GND.n5140 585
R5566 GND.n5142 GND.n5141 585
R5567 GND.n5139 GND.n1069 585
R5568 GND.n1069 GND.n1068 585
R5569 GND.n5138 GND.n5137 585
R5570 GND.n5137 GND.n5136 585
R5571 GND.n1075 GND.n1074 585
R5572 GND.n5135 GND.n1075 585
R5573 GND.n5133 GND.n5132 585
R5574 GND.n5134 GND.n5133 585
R5575 GND.n969 GND.n968 585
R5576 GND.n968 GND.n967 585
R5577 GND.n5247 GND.n5246 585
R5578 GND.n5248 GND.n5247 585
R5579 GND.n966 GND.n965 585
R5580 GND.n5249 GND.n966 585
R5581 GND.n5252 GND.n5251 585
R5582 GND.n5251 GND.n5250 585
R5583 GND.n963 GND.n962 585
R5584 GND.n962 GND.n961 585
R5585 GND.n5257 GND.n5256 585
R5586 GND.n5258 GND.n5257 585
R5587 GND.n960 GND.n959 585
R5588 GND.n5259 GND.n960 585
R5589 GND.n5262 GND.n5261 585
R5590 GND.n5261 GND.n5260 585
R5591 GND.n957 GND.n956 585
R5592 GND.n956 GND.n955 585
R5593 GND.n5267 GND.n5266 585
R5594 GND.n5268 GND.n5267 585
R5595 GND.n954 GND.n953 585
R5596 GND.n5269 GND.n954 585
R5597 GND.n5272 GND.n5271 585
R5598 GND.n5271 GND.n5270 585
R5599 GND.n951 GND.n950 585
R5600 GND.n950 GND.n949 585
R5601 GND.n5277 GND.n5276 585
R5602 GND.n5278 GND.n5277 585
R5603 GND.n948 GND.n947 585
R5604 GND.n5279 GND.n948 585
R5605 GND.n5282 GND.n5281 585
R5606 GND.n5281 GND.n5280 585
R5607 GND.n945 GND.n944 585
R5608 GND.n944 GND.n943 585
R5609 GND.n5287 GND.n5286 585
R5610 GND.n5288 GND.n5287 585
R5611 GND.n942 GND.n941 585
R5612 GND.n5289 GND.n942 585
R5613 GND.n5292 GND.n5291 585
R5614 GND.n5291 GND.n5290 585
R5615 GND.n939 GND.n938 585
R5616 GND.n938 GND.n937 585
R5617 GND.n5297 GND.n5296 585
R5618 GND.n5298 GND.n5297 585
R5619 GND.n936 GND.n935 585
R5620 GND.n5299 GND.n936 585
R5621 GND.n5302 GND.n5301 585
R5622 GND.n5301 GND.n5300 585
R5623 GND.n933 GND.n932 585
R5624 GND.n932 GND.n931 585
R5625 GND.n5307 GND.n5306 585
R5626 GND.n5308 GND.n5307 585
R5627 GND.n930 GND.n929 585
R5628 GND.n5309 GND.n930 585
R5629 GND.n5312 GND.n5311 585
R5630 GND.n5311 GND.n5310 585
R5631 GND.n927 GND.n926 585
R5632 GND.n926 GND.n925 585
R5633 GND.n5317 GND.n5316 585
R5634 GND.n5318 GND.n5317 585
R5635 GND.n924 GND.n923 585
R5636 GND.n5319 GND.n924 585
R5637 GND.n5322 GND.n5321 585
R5638 GND.n5321 GND.n5320 585
R5639 GND.n921 GND.n920 585
R5640 GND.n920 GND.n919 585
R5641 GND.n5327 GND.n5326 585
R5642 GND.n5328 GND.n5327 585
R5643 GND.n918 GND.n917 585
R5644 GND.n5329 GND.n918 585
R5645 GND.n5332 GND.n5331 585
R5646 GND.n5331 GND.n5330 585
R5647 GND.n915 GND.n914 585
R5648 GND.n914 GND.n913 585
R5649 GND.n5337 GND.n5336 585
R5650 GND.n5338 GND.n5337 585
R5651 GND.n912 GND.n911 585
R5652 GND.n5339 GND.n912 585
R5653 GND.n5342 GND.n5341 585
R5654 GND.n5341 GND.n5340 585
R5655 GND.n909 GND.n908 585
R5656 GND.n908 GND.n907 585
R5657 GND.n5347 GND.n5346 585
R5658 GND.n5348 GND.n5347 585
R5659 GND.n906 GND.n905 585
R5660 GND.n5349 GND.n906 585
R5661 GND.n5352 GND.n5351 585
R5662 GND.n5351 GND.n5350 585
R5663 GND.n903 GND.n902 585
R5664 GND.n902 GND.n901 585
R5665 GND.n5357 GND.n5356 585
R5666 GND.n5358 GND.n5357 585
R5667 GND.n900 GND.n899 585
R5668 GND.n5359 GND.n900 585
R5669 GND.n5362 GND.n5361 585
R5670 GND.n5361 GND.n5360 585
R5671 GND.n897 GND.n896 585
R5672 GND.n896 GND.n895 585
R5673 GND.n5367 GND.n5366 585
R5674 GND.n5368 GND.n5367 585
R5675 GND.n894 GND.n893 585
R5676 GND.n5369 GND.n894 585
R5677 GND.n5372 GND.n5371 585
R5678 GND.n5371 GND.n5370 585
R5679 GND.n891 GND.n890 585
R5680 GND.n890 GND.n889 585
R5681 GND.n5377 GND.n5376 585
R5682 GND.n5378 GND.n5377 585
R5683 GND.n888 GND.n887 585
R5684 GND.n5379 GND.n888 585
R5685 GND.n5382 GND.n5381 585
R5686 GND.n5381 GND.n5380 585
R5687 GND.n885 GND.n884 585
R5688 GND.n884 GND.n883 585
R5689 GND.n5387 GND.n5386 585
R5690 GND.n5388 GND.n5387 585
R5691 GND.n882 GND.n881 585
R5692 GND.n5389 GND.n882 585
R5693 GND.n5392 GND.n5391 585
R5694 GND.n5391 GND.n5390 585
R5695 GND.n879 GND.n878 585
R5696 GND.n878 GND.n877 585
R5697 GND.n5397 GND.n5396 585
R5698 GND.n5398 GND.n5397 585
R5699 GND.n876 GND.n875 585
R5700 GND.n5399 GND.n876 585
R5701 GND.n5402 GND.n5401 585
R5702 GND.n5401 GND.n5400 585
R5703 GND.n873 GND.n872 585
R5704 GND.n872 GND.n871 585
R5705 GND.n5407 GND.n5406 585
R5706 GND.n5408 GND.n5407 585
R5707 GND.n870 GND.n869 585
R5708 GND.n5409 GND.n870 585
R5709 GND.n5412 GND.n5411 585
R5710 GND.n5411 GND.n5410 585
R5711 GND.n867 GND.n866 585
R5712 GND.n866 GND.n865 585
R5713 GND.n5417 GND.n5416 585
R5714 GND.n5418 GND.n5417 585
R5715 GND.n864 GND.n863 585
R5716 GND.n5419 GND.n864 585
R5717 GND.n5422 GND.n5421 585
R5718 GND.n5421 GND.n5420 585
R5719 GND.n861 GND.n860 585
R5720 GND.n860 GND.n859 585
R5721 GND.n5427 GND.n5426 585
R5722 GND.n5428 GND.n5427 585
R5723 GND.n858 GND.n857 585
R5724 GND.n5429 GND.n858 585
R5725 GND.n5432 GND.n5431 585
R5726 GND.n5431 GND.n5430 585
R5727 GND.n855 GND.n854 585
R5728 GND.n854 GND.n853 585
R5729 GND.n5437 GND.n5436 585
R5730 GND.n5438 GND.n5437 585
R5731 GND.n852 GND.n851 585
R5732 GND.n5439 GND.n852 585
R5733 GND.n5442 GND.n5441 585
R5734 GND.n5441 GND.n5440 585
R5735 GND.n849 GND.n848 585
R5736 GND.n848 GND.n847 585
R5737 GND.n5447 GND.n5446 585
R5738 GND.n5448 GND.n5447 585
R5739 GND.n846 GND.n845 585
R5740 GND.n5449 GND.n846 585
R5741 GND.n5452 GND.n5451 585
R5742 GND.n5451 GND.n5450 585
R5743 GND.n843 GND.n842 585
R5744 GND.n842 GND.n841 585
R5745 GND.n5457 GND.n5456 585
R5746 GND.n5458 GND.n5457 585
R5747 GND.n840 GND.n839 585
R5748 GND.n5459 GND.n840 585
R5749 GND.n5462 GND.n5461 585
R5750 GND.n5461 GND.n5460 585
R5751 GND.n837 GND.n836 585
R5752 GND.n836 GND.n835 585
R5753 GND.n5467 GND.n5466 585
R5754 GND.n5468 GND.n5467 585
R5755 GND.n834 GND.n833 585
R5756 GND.n5469 GND.n834 585
R5757 GND.n5472 GND.n5471 585
R5758 GND.n5471 GND.n5470 585
R5759 GND.n831 GND.n830 585
R5760 GND.n830 GND.n829 585
R5761 GND.n5477 GND.n5476 585
R5762 GND.n5478 GND.n5477 585
R5763 GND.n828 GND.n827 585
R5764 GND.n5479 GND.n828 585
R5765 GND.n5482 GND.n5481 585
R5766 GND.n5481 GND.n5480 585
R5767 GND.n825 GND.n824 585
R5768 GND.n824 GND.n823 585
R5769 GND.n5487 GND.n5486 585
R5770 GND.n5488 GND.n5487 585
R5771 GND.n822 GND.n821 585
R5772 GND.n5489 GND.n822 585
R5773 GND.n5492 GND.n5491 585
R5774 GND.n5491 GND.n5490 585
R5775 GND.n819 GND.n818 585
R5776 GND.n818 GND.n817 585
R5777 GND.n5497 GND.n5496 585
R5778 GND.n5498 GND.n5497 585
R5779 GND.n816 GND.n815 585
R5780 GND.n5499 GND.n816 585
R5781 GND.n5502 GND.n5501 585
R5782 GND.n5501 GND.n5500 585
R5783 GND.n813 GND.n812 585
R5784 GND.n812 GND.n811 585
R5785 GND.n5507 GND.n5506 585
R5786 GND.n5508 GND.n5507 585
R5787 GND.n810 GND.n809 585
R5788 GND.n5509 GND.n810 585
R5789 GND.n5512 GND.n5511 585
R5790 GND.n5511 GND.n5510 585
R5791 GND.n807 GND.n806 585
R5792 GND.n806 GND.n805 585
R5793 GND.n5517 GND.n5516 585
R5794 GND.n5518 GND.n5517 585
R5795 GND.n804 GND.n803 585
R5796 GND.n5519 GND.n804 585
R5797 GND.n5522 GND.n5521 585
R5798 GND.n5521 GND.n5520 585
R5799 GND.n801 GND.n800 585
R5800 GND.n800 GND.n799 585
R5801 GND.n5527 GND.n5526 585
R5802 GND.n5528 GND.n5527 585
R5803 GND.n798 GND.n797 585
R5804 GND.n5529 GND.n798 585
R5805 GND.n5532 GND.n5531 585
R5806 GND.n5531 GND.n5530 585
R5807 GND.n795 GND.n794 585
R5808 GND.n794 GND.n793 585
R5809 GND.n5537 GND.n5536 585
R5810 GND.n5538 GND.n5537 585
R5811 GND.n792 GND.n791 585
R5812 GND.n5539 GND.n792 585
R5813 GND.n5542 GND.n5541 585
R5814 GND.n5541 GND.n5540 585
R5815 GND.n789 GND.n788 585
R5816 GND.n788 GND.n787 585
R5817 GND.n5547 GND.n5546 585
R5818 GND.n5548 GND.n5547 585
R5819 GND.n786 GND.n785 585
R5820 GND.n5549 GND.n786 585
R5821 GND.n5552 GND.n5551 585
R5822 GND.n5551 GND.n5550 585
R5823 GND.n783 GND.n782 585
R5824 GND.n782 GND.n781 585
R5825 GND.n5557 GND.n5556 585
R5826 GND.n5558 GND.n5557 585
R5827 GND.n780 GND.n779 585
R5828 GND.n5559 GND.n780 585
R5829 GND.n5562 GND.n5561 585
R5830 GND.n5561 GND.n5560 585
R5831 GND.n777 GND.n776 585
R5832 GND.n776 GND.n775 585
R5833 GND.n5567 GND.n5566 585
R5834 GND.n5568 GND.n5567 585
R5835 GND.n774 GND.n773 585
R5836 GND.n5569 GND.n774 585
R5837 GND.n5572 GND.n5571 585
R5838 GND.n5571 GND.n5570 585
R5839 GND.n771 GND.n770 585
R5840 GND.n770 GND.n769 585
R5841 GND.n5577 GND.n5576 585
R5842 GND.n5578 GND.n5577 585
R5843 GND.n768 GND.n767 585
R5844 GND.n5579 GND.n768 585
R5845 GND.n5582 GND.n5581 585
R5846 GND.n5581 GND.n5580 585
R5847 GND.n765 GND.n764 585
R5848 GND.n764 GND.n763 585
R5849 GND.n5587 GND.n5586 585
R5850 GND.n5588 GND.n5587 585
R5851 GND.n762 GND.n761 585
R5852 GND.n5589 GND.n762 585
R5853 GND.n5592 GND.n5591 585
R5854 GND.n5591 GND.n5590 585
R5855 GND.n759 GND.n758 585
R5856 GND.n758 GND.n757 585
R5857 GND.n5597 GND.n5596 585
R5858 GND.n5598 GND.n5597 585
R5859 GND.n756 GND.n755 585
R5860 GND.n5599 GND.n756 585
R5861 GND.n5602 GND.n5601 585
R5862 GND.n5601 GND.n5600 585
R5863 GND.n753 GND.n752 585
R5864 GND.n752 GND.n751 585
R5865 GND.n5607 GND.n5606 585
R5866 GND.n5608 GND.n5607 585
R5867 GND.n750 GND.n749 585
R5868 GND.n5609 GND.n750 585
R5869 GND.n5612 GND.n5611 585
R5870 GND.n5611 GND.n5610 585
R5871 GND.n747 GND.n746 585
R5872 GND.n746 GND.n745 585
R5873 GND.n5617 GND.n5616 585
R5874 GND.n5618 GND.n5617 585
R5875 GND.n744 GND.n743 585
R5876 GND.n5619 GND.n744 585
R5877 GND.n5622 GND.n5621 585
R5878 GND.n5621 GND.n5620 585
R5879 GND.n741 GND.n740 585
R5880 GND.n740 GND.n739 585
R5881 GND.n5627 GND.n5626 585
R5882 GND.n5628 GND.n5627 585
R5883 GND.n738 GND.n737 585
R5884 GND.n5629 GND.n738 585
R5885 GND.n5632 GND.n5631 585
R5886 GND.n5631 GND.n5630 585
R5887 GND.n735 GND.n734 585
R5888 GND.n734 GND.n733 585
R5889 GND.n5637 GND.n5636 585
R5890 GND.n5638 GND.n5637 585
R5891 GND.n732 GND.n731 585
R5892 GND.n5639 GND.n732 585
R5893 GND.n5642 GND.n5641 585
R5894 GND.n5641 GND.n5640 585
R5895 GND.n729 GND.n728 585
R5896 GND.n728 GND.n727 585
R5897 GND.n5647 GND.n5646 585
R5898 GND.n5648 GND.n5647 585
R5899 GND.n726 GND.n725 585
R5900 GND.n5649 GND.n726 585
R5901 GND.n5652 GND.n5651 585
R5902 GND.n5651 GND.n5650 585
R5903 GND.n723 GND.n722 585
R5904 GND.n722 GND.n721 585
R5905 GND.n5657 GND.n5656 585
R5906 GND.n5658 GND.n5657 585
R5907 GND.n720 GND.n719 585
R5908 GND.n5659 GND.n720 585
R5909 GND.n5662 GND.n5661 585
R5910 GND.n5661 GND.n5660 585
R5911 GND.n717 GND.n716 585
R5912 GND.n716 GND.n715 585
R5913 GND.n5667 GND.n5666 585
R5914 GND.n5668 GND.n5667 585
R5915 GND.n714 GND.n713 585
R5916 GND.n5669 GND.n714 585
R5917 GND.n5672 GND.n5671 585
R5918 GND.n5671 GND.n5670 585
R5919 GND.n711 GND.n710 585
R5920 GND.n710 GND.n709 585
R5921 GND.n5677 GND.n5676 585
R5922 GND.n5678 GND.n5677 585
R5923 GND.n708 GND.n707 585
R5924 GND.n5679 GND.n708 585
R5925 GND.n5682 GND.n5681 585
R5926 GND.n5681 GND.n5680 585
R5927 GND.n705 GND.n704 585
R5928 GND.n704 GND.n703 585
R5929 GND.n5687 GND.n5686 585
R5930 GND.n5688 GND.n5687 585
R5931 GND.n702 GND.n701 585
R5932 GND.n5689 GND.n702 585
R5933 GND.n5692 GND.n5691 585
R5934 GND.n5691 GND.n5690 585
R5935 GND.n699 GND.n698 585
R5936 GND.n698 GND.n697 585
R5937 GND.n5697 GND.n5696 585
R5938 GND.n5698 GND.n5697 585
R5939 GND.n696 GND.n695 585
R5940 GND.n5699 GND.n696 585
R5941 GND.n5702 GND.n5701 585
R5942 GND.n5701 GND.n5700 585
R5943 GND.n693 GND.n692 585
R5944 GND.n692 GND.n691 585
R5945 GND.n5707 GND.n5706 585
R5946 GND.n5708 GND.n5707 585
R5947 GND.n690 GND.n689 585
R5948 GND.n5709 GND.n690 585
R5949 GND.n5712 GND.n5711 585
R5950 GND.n5711 GND.n5710 585
R5951 GND.n687 GND.n686 585
R5952 GND.n686 GND.n685 585
R5953 GND.n5717 GND.n5716 585
R5954 GND.n5718 GND.n5717 585
R5955 GND.n684 GND.n683 585
R5956 GND.n5719 GND.n684 585
R5957 GND.n5722 GND.n5721 585
R5958 GND.n5721 GND.n5720 585
R5959 GND.n681 GND.n680 585
R5960 GND.n680 GND.n679 585
R5961 GND.n5727 GND.n5726 585
R5962 GND.n5728 GND.n5727 585
R5963 GND.n678 GND.n677 585
R5964 GND.n5729 GND.n678 585
R5965 GND.n5732 GND.n5731 585
R5966 GND.n5731 GND.n5730 585
R5967 GND.n675 GND.n674 585
R5968 GND.n674 GND.n673 585
R5969 GND.n5737 GND.n5736 585
R5970 GND.n5738 GND.n5737 585
R5971 GND.n672 GND.n671 585
R5972 GND.n5739 GND.n672 585
R5973 GND.n5742 GND.n5741 585
R5974 GND.n5741 GND.n5740 585
R5975 GND.n669 GND.n668 585
R5976 GND.n668 GND.n667 585
R5977 GND.n5747 GND.n5746 585
R5978 GND.n5748 GND.n5747 585
R5979 GND.n666 GND.n665 585
R5980 GND.n5749 GND.n666 585
R5981 GND.n5752 GND.n5751 585
R5982 GND.n5751 GND.n5750 585
R5983 GND.n663 GND.n662 585
R5984 GND.n662 GND.n661 585
R5985 GND.n5757 GND.n5756 585
R5986 GND.n5758 GND.n5757 585
R5987 GND.n660 GND.n659 585
R5988 GND.n5759 GND.n660 585
R5989 GND.n5762 GND.n5761 585
R5990 GND.n5761 GND.n5760 585
R5991 GND.n657 GND.n656 585
R5992 GND.n656 GND.n655 585
R5993 GND.n5767 GND.n5766 585
R5994 GND.n5768 GND.n5767 585
R5995 GND.n654 GND.n653 585
R5996 GND.n5769 GND.n654 585
R5997 GND.n5772 GND.n5771 585
R5998 GND.n5771 GND.n5770 585
R5999 GND.n651 GND.n650 585
R6000 GND.n650 GND.n649 585
R6001 GND.n5777 GND.n5776 585
R6002 GND.n5778 GND.n5777 585
R6003 GND.n648 GND.n647 585
R6004 GND.n5779 GND.n648 585
R6005 GND.n5782 GND.n5781 585
R6006 GND.n5781 GND.n5780 585
R6007 GND.n645 GND.n644 585
R6008 GND.n644 GND.n643 585
R6009 GND.n5787 GND.n5786 585
R6010 GND.n5788 GND.n5787 585
R6011 GND.n642 GND.n641 585
R6012 GND.n5789 GND.n642 585
R6013 GND.n5792 GND.n5791 585
R6014 GND.n5791 GND.n5790 585
R6015 GND.n639 GND.n638 585
R6016 GND.n638 GND.n637 585
R6017 GND.n5797 GND.n5796 585
R6018 GND.n5798 GND.n5797 585
R6019 GND.n636 GND.n635 585
R6020 GND.n5799 GND.n636 585
R6021 GND.n5802 GND.n5801 585
R6022 GND.n5801 GND.n5800 585
R6023 GND.n633 GND.n632 585
R6024 GND.n632 GND.n631 585
R6025 GND.n5807 GND.n5806 585
R6026 GND.n5808 GND.n5807 585
R6027 GND.n630 GND.n629 585
R6028 GND.n5809 GND.n630 585
R6029 GND.n5812 GND.n5811 585
R6030 GND.n5811 GND.n5810 585
R6031 GND.n627 GND.n626 585
R6032 GND.n626 GND.n625 585
R6033 GND.n5817 GND.n5816 585
R6034 GND.n5818 GND.n5817 585
R6035 GND.n624 GND.n623 585
R6036 GND.n5819 GND.n624 585
R6037 GND.n5822 GND.n5821 585
R6038 GND.n5821 GND.n5820 585
R6039 GND.n621 GND.n620 585
R6040 GND.n620 GND.n619 585
R6041 GND.n5827 GND.n5826 585
R6042 GND.n5828 GND.n5827 585
R6043 GND.n618 GND.n617 585
R6044 GND.n5829 GND.n618 585
R6045 GND.n5832 GND.n5831 585
R6046 GND.n5831 GND.n5830 585
R6047 GND.n615 GND.n614 585
R6048 GND.n614 GND.n613 585
R6049 GND.n5837 GND.n5836 585
R6050 GND.n5838 GND.n5837 585
R6051 GND.n612 GND.n611 585
R6052 GND.n5839 GND.n612 585
R6053 GND.n5842 GND.n5841 585
R6054 GND.n5841 GND.n5840 585
R6055 GND.n609 GND.n608 585
R6056 GND.n608 GND.n607 585
R6057 GND.n5847 GND.n5846 585
R6058 GND.n5848 GND.n5847 585
R6059 GND.n606 GND.n605 585
R6060 GND.n5849 GND.n606 585
R6061 GND.n5852 GND.n5851 585
R6062 GND.n5851 GND.n5850 585
R6063 GND.n603 GND.n602 585
R6064 GND.n602 GND.n601 585
R6065 GND.n5857 GND.n5856 585
R6066 GND.n5858 GND.n5857 585
R6067 GND.n600 GND.n599 585
R6068 GND.n5859 GND.n600 585
R6069 GND.n5862 GND.n5861 585
R6070 GND.n5861 GND.n5860 585
R6071 GND.n597 GND.n596 585
R6072 GND.n596 GND.n595 585
R6073 GND.n5867 GND.n5866 585
R6074 GND.n5868 GND.n5867 585
R6075 GND.n594 GND.n593 585
R6076 GND.n5869 GND.n594 585
R6077 GND.n5872 GND.n5871 585
R6078 GND.n5871 GND.n5870 585
R6079 GND.n591 GND.n590 585
R6080 GND.n590 GND.n589 585
R6081 GND.n5877 GND.n5876 585
R6082 GND.n5878 GND.n5877 585
R6083 GND.n588 GND.n587 585
R6084 GND.n5879 GND.n588 585
R6085 GND.n5882 GND.n5881 585
R6086 GND.n5881 GND.n5880 585
R6087 GND.n585 GND.n584 585
R6088 GND.n584 GND.n583 585
R6089 GND.n5887 GND.n5886 585
R6090 GND.n5888 GND.n5887 585
R6091 GND.n582 GND.n581 585
R6092 GND.n5889 GND.n582 585
R6093 GND.n5892 GND.n5891 585
R6094 GND.n5891 GND.n5890 585
R6095 GND.n579 GND.n578 585
R6096 GND.n578 GND.n577 585
R6097 GND.n5897 GND.n5896 585
R6098 GND.n5898 GND.n5897 585
R6099 GND.n576 GND.n575 585
R6100 GND.n5899 GND.n576 585
R6101 GND.n5902 GND.n5901 585
R6102 GND.n5901 GND.n5900 585
R6103 GND.n573 GND.n572 585
R6104 GND.n572 GND.n571 585
R6105 GND.n5907 GND.n5906 585
R6106 GND.n5908 GND.n5907 585
R6107 GND.n570 GND.n569 585
R6108 GND.n5909 GND.n570 585
R6109 GND.n5912 GND.n5911 585
R6110 GND.n5911 GND.n5910 585
R6111 GND.n567 GND.n566 585
R6112 GND.n566 GND.n565 585
R6113 GND.n5917 GND.n5916 585
R6114 GND.n5918 GND.n5917 585
R6115 GND.n564 GND.n563 585
R6116 GND.n5919 GND.n564 585
R6117 GND.n5922 GND.n5921 585
R6118 GND.n5921 GND.n5920 585
R6119 GND.n561 GND.n560 585
R6120 GND.n560 GND.n559 585
R6121 GND.n5927 GND.n5926 585
R6122 GND.n5928 GND.n5927 585
R6123 GND.n558 GND.n557 585
R6124 GND.n5929 GND.n558 585
R6125 GND.n5932 GND.n5931 585
R6126 GND.n5931 GND.n5930 585
R6127 GND.n474 GND.n473 585
R6128 GND.n6069 GND.n474 585
R6129 GND.n6067 GND.n6066 585
R6130 GND.n6068 GND.n6067 585
R6131 GND.n477 GND.n476 585
R6132 GND.n476 GND.n475 585
R6133 GND.n6062 GND.n6061 585
R6134 GND.n6061 GND.n6060 585
R6135 GND.n480 GND.n479 585
R6136 GND.n6059 GND.n480 585
R6137 GND.n6057 GND.n6056 585
R6138 GND.n6058 GND.n6057 585
R6139 GND.n483 GND.n482 585
R6140 GND.n482 GND.n481 585
R6141 GND.n6052 GND.n6051 585
R6142 GND.n6051 GND.n6050 585
R6143 GND.n486 GND.n485 585
R6144 GND.n6049 GND.n486 585
R6145 GND.n6047 GND.n6046 585
R6146 GND.n6048 GND.n6047 585
R6147 GND.n489 GND.n488 585
R6148 GND.n488 GND.n487 585
R6149 GND.n6042 GND.n6041 585
R6150 GND.n6041 GND.n6040 585
R6151 GND.n492 GND.n491 585
R6152 GND.n6039 GND.n492 585
R6153 GND.n6037 GND.n6036 585
R6154 GND.n6038 GND.n6037 585
R6155 GND.n495 GND.n494 585
R6156 GND.n494 GND.n493 585
R6157 GND.n6032 GND.n6031 585
R6158 GND.n6031 GND.n6030 585
R6159 GND.n498 GND.n497 585
R6160 GND.n6029 GND.n498 585
R6161 GND.n6027 GND.n6026 585
R6162 GND.n6028 GND.n6027 585
R6163 GND.n501 GND.n500 585
R6164 GND.n500 GND.n499 585
R6165 GND.n6022 GND.n6021 585
R6166 GND.n6021 GND.n6020 585
R6167 GND.n504 GND.n503 585
R6168 GND.n6019 GND.n504 585
R6169 GND.n6017 GND.n6016 585
R6170 GND.n6018 GND.n6017 585
R6171 GND.n507 GND.n506 585
R6172 GND.n506 GND.n505 585
R6173 GND.n6012 GND.n6011 585
R6174 GND.n6011 GND.n6010 585
R6175 GND.n510 GND.n509 585
R6176 GND.n6009 GND.n510 585
R6177 GND.n6007 GND.n6006 585
R6178 GND.n6008 GND.n6007 585
R6179 GND.n513 GND.n512 585
R6180 GND.n512 GND.n511 585
R6181 GND.n6002 GND.n6001 585
R6182 GND.n6001 GND.n6000 585
R6183 GND.n516 GND.n515 585
R6184 GND.n5999 GND.n516 585
R6185 GND.n5997 GND.n5996 585
R6186 GND.n5998 GND.n5997 585
R6187 GND.n519 GND.n518 585
R6188 GND.n518 GND.n517 585
R6189 GND.n5992 GND.n5991 585
R6190 GND.n5991 GND.n5990 585
R6191 GND.n522 GND.n521 585
R6192 GND.n5989 GND.n522 585
R6193 GND.n5987 GND.n5986 585
R6194 GND.n5988 GND.n5987 585
R6195 GND.n525 GND.n524 585
R6196 GND.n524 GND.n523 585
R6197 GND.n5982 GND.n5981 585
R6198 GND.n5981 GND.n5980 585
R6199 GND.n528 GND.n527 585
R6200 GND.n5979 GND.n528 585
R6201 GND.n5977 GND.n5976 585
R6202 GND.n5978 GND.n5977 585
R6203 GND.n531 GND.n530 585
R6204 GND.n530 GND.n529 585
R6205 GND.n5972 GND.n5971 585
R6206 GND.n5971 GND.n5970 585
R6207 GND.n534 GND.n533 585
R6208 GND.n5969 GND.n534 585
R6209 GND.n5967 GND.n5966 585
R6210 GND.n5968 GND.n5967 585
R6211 GND.n537 GND.n536 585
R6212 GND.n536 GND.n535 585
R6213 GND.n5962 GND.n5961 585
R6214 GND.n5961 GND.n5960 585
R6215 GND.n540 GND.n539 585
R6216 GND.n5959 GND.n540 585
R6217 GND.n5957 GND.n5956 585
R6218 GND.n5958 GND.n5957 585
R6219 GND.n543 GND.n542 585
R6220 GND.n542 GND.n541 585
R6221 GND.n5952 GND.n5951 585
R6222 GND.n5951 GND.n5950 585
R6223 GND.n546 GND.n545 585
R6224 GND.n5949 GND.n546 585
R6225 GND.n5947 GND.n5946 585
R6226 GND.n5948 GND.n5947 585
R6227 GND.n549 GND.n548 585
R6228 GND.n548 GND.n547 585
R6229 GND.n5942 GND.n5941 585
R6230 GND.n5941 GND.n5940 585
R6231 GND.n552 GND.n551 585
R6232 GND.n5939 GND.n552 585
R6233 GND.n5937 GND.n5936 585
R6234 GND.n5938 GND.n5937 585
R6235 GND.n555 GND.n554 585
R6236 GND.n554 GND.n553 585
R6237 GND.n1294 GND.n1293 585
R6238 GND.n4953 GND.n1294 585
R6239 GND.n3868 GND.n1286 585
R6240 GND.n3869 GND.n3868 585
R6241 GND.n3867 GND.n1285 585
R6242 GND.n3867 GND.n3866 585
R6243 GND.n2972 GND.n1284 585
R6244 GND.n3846 GND.n2972 585
R6245 GND.n3857 GND.n3856 585
R6246 GND.n3858 GND.n3857 585
R6247 GND.n3855 GND.n1278 585
R6248 GND.n3855 GND.n3854 585
R6249 GND.n2983 GND.n1277 585
R6250 GND.n2996 GND.n2983 585
R6251 GND.n2993 GND.n1276 585
R6252 GND.n3840 GND.n2993 585
R6253 GND.n3828 GND.n3826 585
R6254 GND.n3828 GND.n3827 585
R6255 GND.n3829 GND.n1270 585
R6256 GND.n3830 GND.n3829 585
R6257 GND.n3825 GND.n1269 585
R6258 GND.n3825 GND.n3824 585
R6259 GND.n3005 GND.n1268 585
R6260 GND.n3019 GND.n3005 585
R6261 GND.n3017 GND.n3016 585
R6262 GND.n3815 GND.n3017 585
R6263 GND.n3803 GND.n1262 585
R6264 GND.n3803 GND.n3802 585
R6265 GND.n3804 GND.n1261 585
R6266 GND.n3805 GND.n3804 585
R6267 GND.n3801 GND.n1260 585
R6268 GND.n3801 GND.n3800 585
R6269 GND.n3030 GND.n3029 585
R6270 GND.n3042 GND.n3030 585
R6271 GND.n3040 GND.n1254 585
R6272 GND.n3791 GND.n3040 585
R6273 GND.n3779 GND.n1253 585
R6274 GND.n3779 GND.n3778 585
R6275 GND.n3780 GND.n1252 585
R6276 GND.n3781 GND.n3780 585
R6277 GND.n3776 GND.n3052 585
R6278 GND.n3776 GND.n3775 585
R6279 GND.n3051 GND.n1246 585
R6280 GND.n3065 GND.n3051 585
R6281 GND.n3063 GND.n1245 585
R6282 GND.n3766 GND.n3063 585
R6283 GND.n3725 GND.n1244 585
R6284 GND.n3726 GND.n3725 585
R6285 GND.n3724 GND.n3723 585
R6286 GND.n3724 GND.n3722 585
R6287 GND.n3104 GND.n1238 585
R6288 GND.n3107 GND.n3104 585
R6289 GND.n3736 GND.n1237 585
R6290 GND.n3736 GND.n3735 585
R6291 GND.n3737 GND.n1236 585
R6292 GND.n3738 GND.n3737 585
R6293 GND.n3096 GND.n3095 585
R6294 GND.n3743 GND.n3096 585
R6295 GND.n3094 GND.n1230 585
R6296 GND.n3094 GND.n3092 585
R6297 GND.n3082 GND.n1229 585
R6298 GND.n3085 GND.n3082 585
R6299 GND.n3753 GND.n1228 585
R6300 GND.n3753 GND.n3752 585
R6301 GND.n3755 GND.n3754 585
R6302 GND.n3756 GND.n3755 585
R6303 GND.n3081 GND.n1222 585
R6304 GND.n3216 GND.n3081 585
R6305 GND.n3218 GND.n1221 585
R6306 GND.n3694 GND.n3218 585
R6307 GND.n3683 GND.n1220 585
R6308 GND.n3683 GND.n3682 585
R6309 GND.n3685 GND.n3684 585
R6310 GND.n3686 GND.n3685 585
R6311 GND.n3681 GND.n1214 585
R6312 GND.n3681 GND.n3680 585
R6313 GND.n3227 GND.n1213 585
R6314 GND.n3240 GND.n3227 585
R6315 GND.n3237 GND.n1212 585
R6316 GND.n3671 GND.n3237 585
R6317 GND.n3659 GND.n3657 585
R6318 GND.n3659 GND.n3658 585
R6319 GND.n3660 GND.n1206 585
R6320 GND.n3661 GND.n3660 585
R6321 GND.n3656 GND.n1205 585
R6322 GND.n3656 GND.n3655 585
R6323 GND.n3249 GND.n1204 585
R6324 GND.n3263 GND.n3249 585
R6325 GND.n3261 GND.n3260 585
R6326 GND.n3646 GND.n3261 585
R6327 GND.n3634 GND.n1198 585
R6328 GND.n3634 GND.n3633 585
R6329 GND.n3635 GND.n1197 585
R6330 GND.n3636 GND.n3635 585
R6331 GND.n3632 GND.n1196 585
R6332 GND.n3632 GND.n3631 585
R6333 GND.n3274 GND.n3273 585
R6334 GND.n3286 GND.n3274 585
R6335 GND.n3284 GND.n1190 585
R6336 GND.n3622 GND.n3284 585
R6337 GND.n3610 GND.n1189 585
R6338 GND.n3610 GND.n3609 585
R6339 GND.n3611 GND.n1188 585
R6340 GND.n3612 GND.n3611 585
R6341 GND.n1181 GND.n1179 585
R6342 GND.n3291 GND.n1179 585
R6343 GND.n5037 GND.n5036 585
R6344 GND.n5038 GND.n5037 585
R6345 GND.n1180 GND.n1178 585
R6346 GND.n3528 GND.n1178 585
R6347 GND.n3490 GND.n1166 585
R6348 GND.n5044 GND.n1166 585
R6349 GND.n3496 GND.n3495 585
R6350 GND.n3498 GND.n3307 585
R6351 GND.n3501 GND.n3500 585
R6352 GND.n3305 GND.n3304 585
R6353 GND.n3506 GND.n3505 585
R6354 GND.n3508 GND.n3303 585
R6355 GND.n3511 GND.n3510 585
R6356 GND.n3301 GND.n3300 585
R6357 GND.n3517 GND.n3516 585
R6358 GND.n3519 GND.n3299 585
R6359 GND.n3520 GND.n3298 585
R6360 GND.n3523 GND.n3522 585
R6361 GND.n4835 GND.n4834 585
R6362 GND.n4836 GND.n1443 585
R6363 GND.n1442 GND.n1433 585
R6364 GND.n4846 GND.n1432 585
R6365 GND.n4847 GND.n1431 585
R6366 GND.n1429 GND.n1423 585
R6367 GND.n4854 GND.n1422 585
R6368 GND.n4855 GND.n1420 585
R6369 GND.n1419 GND.n1412 585
R6370 GND.n4862 GND.n1411 585
R6371 GND.n4863 GND.n1410 585
R6372 GND.n1408 GND.n1407 585
R6373 GND.n3872 GND.n1291 585
R6374 GND.n4953 GND.n1291 585
R6375 GND.n3871 GND.n3870 585
R6376 GND.n3870 GND.n3869 585
R6377 GND.n2970 GND.n2969 585
R6378 GND.n3866 GND.n2970 585
R6379 GND.n3848 GND.n3847 585
R6380 GND.n3847 GND.n3846 585
R6381 GND.n2987 GND.n2981 585
R6382 GND.n3858 GND.n2981 585
R6383 GND.n3853 GND.n3852 585
R6384 GND.n3854 GND.n3853 585
R6385 GND.n2986 GND.n2985 585
R6386 GND.n2996 GND.n2985 585
R6387 GND.n3842 GND.n3841 585
R6388 GND.n3841 GND.n3840 585
R6389 GND.n2990 GND.n2989 585
R6390 GND.n3827 GND.n2990 585
R6391 GND.n3010 GND.n3003 585
R6392 GND.n3830 GND.n3003 585
R6393 GND.n3823 GND.n3822 585
R6394 GND.n3824 GND.n3823 585
R6395 GND.n3009 GND.n3008 585
R6396 GND.n3019 GND.n3008 585
R6397 GND.n3817 GND.n3816 585
R6398 GND.n3816 GND.n3815 585
R6399 GND.n3013 GND.n3012 585
R6400 GND.n3802 GND.n3013 585
R6401 GND.n3034 GND.n3027 585
R6402 GND.n3805 GND.n3027 585
R6403 GND.n3799 GND.n3798 585
R6404 GND.n3800 GND.n3799 585
R6405 GND.n3033 GND.n3032 585
R6406 GND.n3042 GND.n3032 585
R6407 GND.n3793 GND.n3792 585
R6408 GND.n3792 GND.n3791 585
R6409 GND.n3037 GND.n3036 585
R6410 GND.n3778 GND.n3037 585
R6411 GND.n3056 GND.n3049 585
R6412 GND.n3781 GND.n3049 585
R6413 GND.n3774 GND.n3773 585
R6414 GND.n3775 GND.n3774 585
R6415 GND.n3055 GND.n3054 585
R6416 GND.n3065 GND.n3054 585
R6417 GND.n3768 GND.n3767 585
R6418 GND.n3767 GND.n3766 585
R6419 GND.n3059 GND.n3058 585
R6420 GND.n3726 GND.n3059 585
R6421 GND.n3716 GND.n3715 585
R6422 GND.n3722 GND.n3716 585
R6423 GND.n3205 GND.n3204 585
R6424 GND.n3204 GND.n3107 585
R6425 GND.n3711 GND.n3106 585
R6426 GND.n3735 GND.n3106 585
R6427 GND.n3710 GND.n3102 585
R6428 GND.n3738 GND.n3102 585
R6429 GND.n3709 GND.n3093 585
R6430 GND.n3743 GND.n3093 585
R6431 GND.n3702 GND.n3207 585
R6432 GND.n3702 GND.n3092 585
R6433 GND.n3704 GND.n3703 585
R6434 GND.n3703 GND.n3085 585
R6435 GND.n3701 GND.n3083 585
R6436 GND.n3752 GND.n3083 585
R6437 GND.n3700 GND.n3079 585
R6438 GND.n3756 GND.n3079 585
R6439 GND.n3213 GND.n3209 585
R6440 GND.n3216 GND.n3213 585
R6441 GND.n3696 GND.n3695 585
R6442 GND.n3695 GND.n3694 585
R6443 GND.n3212 GND.n3211 585
R6444 GND.n3682 GND.n3212 585
R6445 GND.n3231 GND.n3225 585
R6446 GND.n3686 GND.n3225 585
R6447 GND.n3679 GND.n3678 585
R6448 GND.n3680 GND.n3679 585
R6449 GND.n3230 GND.n3229 585
R6450 GND.n3240 GND.n3229 585
R6451 GND.n3673 GND.n3672 585
R6452 GND.n3672 GND.n3671 585
R6453 GND.n3234 GND.n3233 585
R6454 GND.n3658 GND.n3234 585
R6455 GND.n3254 GND.n3247 585
R6456 GND.n3661 GND.n3247 585
R6457 GND.n3654 GND.n3653 585
R6458 GND.n3655 GND.n3654 585
R6459 GND.n3253 GND.n3252 585
R6460 GND.n3263 GND.n3252 585
R6461 GND.n3648 GND.n3647 585
R6462 GND.n3647 GND.n3646 585
R6463 GND.n3257 GND.n3256 585
R6464 GND.n3633 GND.n3257 585
R6465 GND.n3278 GND.n3271 585
R6466 GND.n3636 GND.n3271 585
R6467 GND.n3630 GND.n3629 585
R6468 GND.n3631 GND.n3630 585
R6469 GND.n3277 GND.n3276 585
R6470 GND.n3286 GND.n3276 585
R6471 GND.n3624 GND.n3623 585
R6472 GND.n3623 GND.n3622 585
R6473 GND.n3281 GND.n3280 585
R6474 GND.n3609 GND.n3281 585
R6475 GND.n3536 GND.n3535 585
R6476 GND.n3612 GND.n3536 585
R6477 GND.n3293 GND.n3292 585
R6478 GND.n3292 GND.n3291 585
R6479 GND.n3531 GND.n1176 585
R6480 GND.n5038 GND.n1176 585
R6481 GND.n3530 GND.n3529 585
R6482 GND.n3529 GND.n3528 585
R6483 GND.n3526 GND.n1164 585
R6484 GND.n5044 GND.n1164 585
R6485 GND.n285 GND.n284 585
R6486 GND.n6159 GND.n285 585
R6487 GND.n6264 GND.n6263 585
R6488 GND.n6263 GND.n6262 585
R6489 GND.n6265 GND.n280 585
R6490 GND.n4438 GND.n280 585
R6491 GND.n6267 GND.n6266 585
R6492 GND.n6268 GND.n6267 585
R6493 GND.n265 GND.n264 585
R6494 GND.n4444 GND.n265 585
R6495 GND.n6276 GND.n6275 585
R6496 GND.n6275 GND.n6274 585
R6497 GND.n6277 GND.n260 585
R6498 GND.n4450 GND.n260 585
R6499 GND.n6279 GND.n6278 585
R6500 GND.n6280 GND.n6279 585
R6501 GND.n244 GND.n243 585
R6502 GND.n4380 GND.n244 585
R6503 GND.n6288 GND.n6287 585
R6504 GND.n6287 GND.n6286 585
R6505 GND.n6289 GND.n239 585
R6506 GND.n4371 GND.n239 585
R6507 GND.n6291 GND.n6290 585
R6508 GND.n6292 GND.n6291 585
R6509 GND.n223 GND.n222 585
R6510 GND.n4365 GND.n223 585
R6511 GND.n6300 GND.n6299 585
R6512 GND.n6299 GND.n6298 585
R6513 GND.n6301 GND.n218 585
R6514 GND.n4357 GND.n218 585
R6515 GND.n6303 GND.n6302 585
R6516 GND.n6304 GND.n6303 585
R6517 GND.n203 GND.n202 585
R6518 GND.n4351 GND.n203 585
R6519 GND.n6312 GND.n6311 585
R6520 GND.n6311 GND.n6310 585
R6521 GND.n6313 GND.n198 585
R6522 GND.n4472 GND.n198 585
R6523 GND.n6315 GND.n6314 585
R6524 GND.n6316 GND.n6315 585
R6525 GND.n183 GND.n182 585
R6526 GND.n4478 GND.n183 585
R6527 GND.n6324 GND.n6323 585
R6528 GND.n6323 GND.n6322 585
R6529 GND.n6325 GND.n177 585
R6530 GND.n4484 GND.n177 585
R6531 GND.n6327 GND.n6326 585
R6532 GND.n6328 GND.n6327 585
R6533 GND.n178 GND.n176 585
R6534 GND.n4490 GND.n176 585
R6535 GND.n4496 GND.n4495 585
R6536 GND.n4499 GND.n4496 585
R6537 GND.n1895 GND.n1894 585
R6538 GND.n1894 GND.n1890 585
R6539 GND.n4256 GND.n156 585
R6540 GND.n6335 GND.n156 585
R6541 GND.n4255 GND.n4254 585
R6542 GND.n4254 GND.n1801 585
R6543 GND.n1793 GND.n1792 585
R6544 GND.n4509 GND.n1793 585
R6545 GND.n4514 GND.n4513 585
R6546 GND.n4513 GND.n4512 585
R6547 GND.n4515 GND.n1788 585
R6548 GND.n4247 GND.n1788 585
R6549 GND.n4517 GND.n4516 585
R6550 GND.n4518 GND.n4517 585
R6551 GND.n1774 GND.n1773 585
R6552 GND.n4235 GND.n1774 585
R6553 GND.n4526 GND.n4525 585
R6554 GND.n4525 GND.n4524 585
R6555 GND.n4527 GND.n1769 585
R6556 GND.n4228 GND.n1769 585
R6557 GND.n4529 GND.n4528 585
R6558 GND.n4530 GND.n4529 585
R6559 GND.n1753 GND.n1752 585
R6560 GND.n4220 GND.n1753 585
R6561 GND.n4538 GND.n4537 585
R6562 GND.n4537 GND.n4536 585
R6563 GND.n4539 GND.n1748 585
R6564 GND.n4213 GND.n1748 585
R6565 GND.n4541 GND.n4540 585
R6566 GND.n4542 GND.n4541 585
R6567 GND.n1732 GND.n1731 585
R6568 GND.n4205 GND.n1732 585
R6569 GND.n4550 GND.n4549 585
R6570 GND.n4549 GND.n4548 585
R6571 GND.n4551 GND.n1727 585
R6572 GND.n4198 GND.n1727 585
R6573 GND.n4553 GND.n4552 585
R6574 GND.n4554 GND.n4553 585
R6575 GND.n1711 GND.n1710 585
R6576 GND.n4190 GND.n1711 585
R6577 GND.n4562 GND.n4561 585
R6578 GND.n4561 GND.n4560 585
R6579 GND.n4563 GND.n1706 585
R6580 GND.n4183 GND.n1706 585
R6581 GND.n4565 GND.n4564 585
R6582 GND.n4566 GND.n4565 585
R6583 GND.n1690 GND.n1689 585
R6584 GND.n4175 GND.n1690 585
R6585 GND.n4574 GND.n4573 585
R6586 GND.n4573 GND.n4572 585
R6587 GND.n4575 GND.n1684 585
R6588 GND.n4168 GND.n1684 585
R6589 GND.n4577 GND.n4576 585
R6590 GND.n4578 GND.n4577 585
R6591 GND.n1685 GND.n1668 585
R6592 GND.n4160 GND.n1668 585
R6593 GND.n4585 GND.n1669 585
R6594 GND.n4585 GND.n4584 585
R6595 GND.n4586 GND.n1660 585
R6596 GND.n4587 GND.n4586 585
R6597 GND.n1946 GND.n1667 585
R6598 GND.n1989 GND.n1988 585
R6599 GND.n1991 GND.n1990 585
R6600 GND.n1994 GND.n1993 585
R6601 GND.n1992 GND.n1939 585
R6602 GND.n2008 GND.n2007 585
R6603 GND.n2010 GND.n2009 585
R6604 GND.n2013 GND.n2012 585
R6605 GND.n2011 GND.n1931 585
R6606 GND.n2029 GND.n1932 585
R6607 GND.n2030 GND.n1928 585
R6608 GND.n2032 GND.n2031 585
R6609 GND.n4431 GND.n4430 585
R6610 GND.n4428 GND.n4393 585
R6611 GND.n4427 GND.n4426 585
R6612 GND.n4420 GND.n4395 585
R6613 GND.n4422 GND.n4421 585
R6614 GND.n4418 GND.n4397 585
R6615 GND.n4417 GND.n4416 585
R6616 GND.n4410 GND.n4399 585
R6617 GND.n4412 GND.n4411 585
R6618 GND.n4408 GND.n4401 585
R6619 GND.n4407 GND.n4406 585
R6620 GND.n4404 GND.n4403 585
R6621 GND.n4434 GND.n386 585
R6622 GND.n6159 GND.n386 585
R6623 GND.n4435 GND.n288 585
R6624 GND.n6262 GND.n288 585
R6625 GND.n4437 GND.n4436 585
R6626 GND.n4438 GND.n4437 585
R6627 GND.n4333 GND.n278 585
R6628 GND.n6268 GND.n278 585
R6629 GND.n4446 GND.n4445 585
R6630 GND.n4445 GND.n4444 585
R6631 GND.n4447 GND.n267 585
R6632 GND.n6274 GND.n267 585
R6633 GND.n4449 GND.n4448 585
R6634 GND.n4450 GND.n4449 585
R6635 GND.n4329 GND.n258 585
R6636 GND.n6280 GND.n258 585
R6637 GND.n4379 GND.n4378 585
R6638 GND.n4380 GND.n4379 585
R6639 GND.n4336 GND.n247 585
R6640 GND.n6286 GND.n247 585
R6641 GND.n4373 GND.n4372 585
R6642 GND.n4372 GND.n4371 585
R6643 GND.n4338 GND.n237 585
R6644 GND.n6292 GND.n237 585
R6645 GND.n4364 GND.n4363 585
R6646 GND.n4365 GND.n4364 585
R6647 GND.n4341 GND.n226 585
R6648 GND.n6298 GND.n226 585
R6649 GND.n4359 GND.n4358 585
R6650 GND.n4358 GND.n4357 585
R6651 GND.n4343 GND.n216 585
R6652 GND.n6304 GND.n216 585
R6653 GND.n4350 GND.n4349 585
R6654 GND.n4351 GND.n4350 585
R6655 GND.n4274 GND.n205 585
R6656 GND.n6310 GND.n205 585
R6657 GND.n4474 GND.n4473 585
R6658 GND.n4473 GND.n4472 585
R6659 GND.n4475 GND.n196 585
R6660 GND.n6316 GND.n196 585
R6661 GND.n4477 GND.n4476 585
R6662 GND.n4478 GND.n4477 585
R6663 GND.n4267 GND.n186 585
R6664 GND.n6322 GND.n186 585
R6665 GND.n4486 GND.n4485 585
R6666 GND.n4485 GND.n4484 585
R6667 GND.n4487 GND.n174 585
R6668 GND.n6328 GND.n174 585
R6669 GND.n4489 GND.n4488 585
R6670 GND.n4490 GND.n4489 585
R6671 GND.n4262 GND.n1892 585
R6672 GND.n4499 GND.n1892 585
R6673 GND.n153 GND.n151 585
R6674 GND.n1890 GND.n153 585
R6675 GND.n6337 GND.n6336 585
R6676 GND.n6336 GND.n6335 585
R6677 GND.n152 GND.n150 585
R6678 GND.n1801 GND.n152 585
R6679 GND.n4243 GND.n1800 585
R6680 GND.n4509 GND.n1800 585
R6681 GND.n4244 GND.n1796 585
R6682 GND.n4512 GND.n1796 585
R6683 GND.n4246 GND.n4245 585
R6684 GND.n4247 GND.n4246 585
R6685 GND.n1901 GND.n1786 585
R6686 GND.n4518 GND.n1786 585
R6687 GND.n4237 GND.n4236 585
R6688 GND.n4236 GND.n4235 585
R6689 GND.n1903 GND.n1777 585
R6690 GND.n4524 GND.n1777 585
R6691 GND.n4227 GND.n4226 585
R6692 GND.n4228 GND.n4227 585
R6693 GND.n1905 GND.n1767 585
R6694 GND.n4530 GND.n1767 585
R6695 GND.n4222 GND.n4221 585
R6696 GND.n4221 GND.n4220 585
R6697 GND.n1907 GND.n1756 585
R6698 GND.n4536 GND.n1756 585
R6699 GND.n4212 GND.n4211 585
R6700 GND.n4213 GND.n4212 585
R6701 GND.n1909 GND.n1746 585
R6702 GND.n4542 GND.n1746 585
R6703 GND.n4207 GND.n4206 585
R6704 GND.n4206 GND.n4205 585
R6705 GND.n1911 GND.n1735 585
R6706 GND.n4548 GND.n1735 585
R6707 GND.n4197 GND.n4196 585
R6708 GND.n4198 GND.n4197 585
R6709 GND.n1913 GND.n1725 585
R6710 GND.n4554 GND.n1725 585
R6711 GND.n4192 GND.n4191 585
R6712 GND.n4191 GND.n4190 585
R6713 GND.n1915 GND.n1714 585
R6714 GND.n4560 GND.n1714 585
R6715 GND.n4182 GND.n4181 585
R6716 GND.n4183 GND.n4182 585
R6717 GND.n1917 GND.n1704 585
R6718 GND.n4566 GND.n1704 585
R6719 GND.n4177 GND.n4176 585
R6720 GND.n4176 GND.n4175 585
R6721 GND.n1919 GND.n1693 585
R6722 GND.n4572 GND.n1693 585
R6723 GND.n4167 GND.n4166 585
R6724 GND.n4168 GND.n4167 585
R6725 GND.n1921 GND.n1682 585
R6726 GND.n4578 GND.n1682 585
R6727 GND.n4162 GND.n4161 585
R6728 GND.n4161 GND.n4160 585
R6729 GND.n4156 GND.n1670 585
R6730 GND.n4584 GND.n1670 585
R6731 GND.n4155 GND.n1665 585
R6732 GND.n4587 GND.n1665 585
R6733 GND.n2671 GND.n2507 585
R6734 GND.n2671 GND.n2067 585
R6735 GND.n2673 GND.n2672 585
R6736 GND.n2672 GND.n2077 585
R6737 GND.n2674 GND.n2502 585
R6738 GND.n2502 GND.n2074 585
R6739 GND.n2676 GND.n2675 585
R6740 GND.n2677 GND.n2676 585
R6741 GND.n2506 GND.n2501 585
R6742 GND.n2501 GND.n2084 585
R6743 GND.n2505 GND.n2504 585
R6744 GND.n2504 GND.n2083 585
R6745 GND.n2503 GND.n2492 585
R6746 GND.n2684 GND.n2492 585
R6747 GND.n2687 GND.n2491 585
R6748 GND.n2687 GND.n2686 585
R6749 GND.n2689 GND.n2688 585
R6750 GND.n2688 GND.n2090 585
R6751 GND.n2690 GND.n2489 585
R6752 GND.n2489 GND.n2488 585
R6753 GND.n2692 GND.n2691 585
R6754 GND.n2693 GND.n2692 585
R6755 GND.n2490 GND.n2479 585
R6756 GND.n2479 GND.n2097 585
R6757 GND.n2700 GND.n2478 585
R6758 GND.n2700 GND.n2699 585
R6759 GND.n2702 GND.n2701 585
R6760 GND.n2701 GND.n2105 585
R6761 GND.n2703 GND.n2475 585
R6762 GND.n2475 GND.n2103 585
R6763 GND.n2705 GND.n2704 585
R6764 GND.n2706 GND.n2705 585
R6765 GND.n2477 GND.n2474 585
R6766 GND.n2474 GND.n2112 585
R6767 GND.n2476 GND.n2465 585
R6768 GND.n2465 GND.n2111 585
R6769 GND.n2714 GND.n2464 585
R6770 GND.n2714 GND.n2713 585
R6771 GND.n2716 GND.n2715 585
R6772 GND.n2715 GND.n2120 585
R6773 GND.n2717 GND.n2460 585
R6774 GND.n2460 GND.n2118 585
R6775 GND.n2719 GND.n2718 585
R6776 GND.n2720 GND.n2719 585
R6777 GND.n2463 GND.n2459 585
R6778 GND.n2459 GND.n2127 585
R6779 GND.n2462 GND.n2461 585
R6780 GND.n2461 GND.n2126 585
R6781 GND.n2451 GND.n2450 585
R6782 GND.n2727 GND.n2451 585
R6783 GND.n2731 GND.n2730 585
R6784 GND.n2730 GND.n2729 585
R6785 GND.n2732 GND.n2447 585
R6786 GND.n2447 GND.n2133 585
R6787 GND.n2734 GND.n2733 585
R6788 GND.n2735 GND.n2734 585
R6789 GND.n2449 GND.n2446 585
R6790 GND.n2446 GND.n2141 585
R6791 GND.n2448 GND.n2438 585
R6792 GND.n2438 GND.n2140 585
R6793 GND.n2744 GND.n2437 585
R6794 GND.n2744 GND.n2743 585
R6795 GND.n2746 GND.n2745 585
R6796 GND.n2745 GND.n2148 585
R6797 GND.n2747 GND.n2434 585
R6798 GND.n2434 GND.n2433 585
R6799 GND.n2749 GND.n2748 585
R6800 GND.n2750 GND.n2749 585
R6801 GND.n2436 GND.n2432 585
R6802 GND.n2432 GND.n2155 585
R6803 GND.n2435 GND.n2424 585
R6804 GND.n2424 GND.n2154 585
R6805 GND.n2759 GND.n2423 585
R6806 GND.n2759 GND.n2758 585
R6807 GND.n2761 GND.n2760 585
R6808 GND.n2760 GND.n2163 585
R6809 GND.n2762 GND.n2420 585
R6810 GND.n2420 GND.n2161 585
R6811 GND.n2764 GND.n2763 585
R6812 GND.n2765 GND.n2764 585
R6813 GND.n2422 GND.n2419 585
R6814 GND.n2419 GND.n2170 585
R6815 GND.n2421 GND.n2411 585
R6816 GND.n2411 GND.n2169 585
R6817 GND.n2774 GND.n2410 585
R6818 GND.n2774 GND.n2773 585
R6819 GND.n2776 GND.n2775 585
R6820 GND.n2775 GND.n2177 585
R6821 GND.n2777 GND.n2395 585
R6822 GND.n2395 GND.n2394 585
R6823 GND.n2779 GND.n2778 585
R6824 GND.n2780 GND.n2779 585
R6825 GND.n2409 GND.n2393 585
R6826 GND.n2393 GND.n2184 585
R6827 GND.n2408 GND.n2407 585
R6828 GND.n2407 GND.n2183 585
R6829 GND.n2406 GND.n2396 585
R6830 GND.n2406 GND.n2405 585
R6831 GND.n2403 GND.n2402 585
R6832 GND.n2403 GND.n2192 585
R6833 GND.n2401 GND.n2397 585
R6834 GND.n2397 GND.n2190 585
R6835 GND.n2400 GND.n2399 585
R6836 GND.n2399 GND.n2200 585
R6837 GND.n2398 GND.n2379 585
R6838 GND.n2379 GND.n2198 585
R6839 GND.n2795 GND.n2380 585
R6840 GND.n2795 GND.n2794 585
R6841 GND.n2796 GND.n2378 585
R6842 GND.n2796 GND.n2208 585
R6843 GND.n2798 GND.n2797 585
R6844 GND.n2797 GND.n2206 585
R6845 GND.n2799 GND.n2376 585
R6846 GND.n2376 GND.n2375 585
R6847 GND.n2801 GND.n2800 585
R6848 GND.n2802 GND.n2801 585
R6849 GND.n2377 GND.n2366 585
R6850 GND.n2366 GND.n2214 585
R6851 GND.n2809 GND.n2365 585
R6852 GND.n2809 GND.n2808 585
R6853 GND.n2811 GND.n2810 585
R6854 GND.n2810 GND.n2222 585
R6855 GND.n2812 GND.n2361 585
R6856 GND.n2361 GND.n2220 585
R6857 GND.n2814 GND.n2813 585
R6858 GND.n2815 GND.n2814 585
R6859 GND.n2364 GND.n2360 585
R6860 GND.n2360 GND.n2229 585
R6861 GND.n2363 GND.n2362 585
R6862 GND.n2362 GND.n2228 585
R6863 GND.n2352 GND.n2351 585
R6864 GND.n2822 GND.n2352 585
R6865 GND.n2826 GND.n2825 585
R6866 GND.n2825 GND.n2824 585
R6867 GND.n2827 GND.n2348 585
R6868 GND.n2348 GND.n2235 585
R6869 GND.n2829 GND.n2828 585
R6870 GND.n2830 GND.n2829 585
R6871 GND.n2350 GND.n2347 585
R6872 GND.n2347 GND.n2243 585
R6873 GND.n2349 GND.n2338 585
R6874 GND.n2338 GND.n2242 585
R6875 GND.n2838 GND.n2337 585
R6876 GND.n2838 GND.n2837 585
R6877 GND.n2840 GND.n2839 585
R6878 GND.n2839 GND.n2251 585
R6879 GND.n2841 GND.n2334 585
R6880 GND.n2334 GND.n2249 585
R6881 GND.n2843 GND.n2842 585
R6882 GND.n2844 GND.n2843 585
R6883 GND.n2336 GND.n2333 585
R6884 GND.n2333 GND.n2258 585
R6885 GND.n2335 GND.n2293 585
R6886 GND.n2293 GND.n2257 585
R6887 GND.n2945 GND.n2944 585
R6888 GND.n2943 GND.n2292 585
R6889 GND.n2942 GND.n2291 585
R6890 GND.n2947 GND.n2291 585
R6891 GND.n2941 GND.n2940 585
R6892 GND.n2939 GND.n2938 585
R6893 GND.n2937 GND.n2936 585
R6894 GND.n2935 GND.n2934 585
R6895 GND.n2933 GND.n2932 585
R6896 GND.n2931 GND.n2930 585
R6897 GND.n2929 GND.n2928 585
R6898 GND.n2927 GND.n2926 585
R6899 GND.n2925 GND.n2924 585
R6900 GND.n2923 GND.n2922 585
R6901 GND.n2921 GND.n2920 585
R6902 GND.n2919 GND.n2918 585
R6903 GND.n2917 GND.n2916 585
R6904 GND.n2915 GND.n2914 585
R6905 GND.n2913 GND.n2912 585
R6906 GND.n2911 GND.n2910 585
R6907 GND.n2909 GND.n2908 585
R6908 GND.n2906 GND.n2905 585
R6909 GND.n2904 GND.n2903 585
R6910 GND.n2902 GND.n2901 585
R6911 GND.n2900 GND.n2899 585
R6912 GND.n2896 GND.n2895 585
R6913 GND.n2894 GND.n2893 585
R6914 GND.n2892 GND.n2891 585
R6915 GND.n2890 GND.n2889 585
R6916 GND.n2887 GND.n2886 585
R6917 GND.n2885 GND.n2884 585
R6918 GND.n2883 GND.n2882 585
R6919 GND.n2881 GND.n2880 585
R6920 GND.n2879 GND.n2878 585
R6921 GND.n2877 GND.n2876 585
R6922 GND.n2875 GND.n2874 585
R6923 GND.n2873 GND.n2872 585
R6924 GND.n2871 GND.n2870 585
R6925 GND.n2869 GND.n2868 585
R6926 GND.n2867 GND.n2866 585
R6927 GND.n2865 GND.n2864 585
R6928 GND.n2863 GND.n2862 585
R6929 GND.n2861 GND.n2860 585
R6930 GND.n2859 GND.n2858 585
R6931 GND.n2857 GND.n2856 585
R6932 GND.n2855 GND.n2854 585
R6933 GND.n2853 GND.n2852 585
R6934 GND.n2851 GND.n2850 585
R6935 GND.n2849 GND.n2289 585
R6936 GND.n2947 GND.n2289 585
R6937 GND.n2586 GND.n2585 585
R6938 GND.n2587 GND.n2578 585
R6939 GND.n2589 GND.n2588 585
R6940 GND.n2591 GND.n2576 585
R6941 GND.n2593 GND.n2592 585
R6942 GND.n2594 GND.n2575 585
R6943 GND.n2596 GND.n2595 585
R6944 GND.n2598 GND.n2573 585
R6945 GND.n2600 GND.n2599 585
R6946 GND.n2601 GND.n2572 585
R6947 GND.n2603 GND.n2602 585
R6948 GND.n2605 GND.n2570 585
R6949 GND.n2607 GND.n2606 585
R6950 GND.n2608 GND.n2569 585
R6951 GND.n2610 GND.n2609 585
R6952 GND.n2612 GND.n2567 585
R6953 GND.n2614 GND.n2613 585
R6954 GND.n2615 GND.n2566 585
R6955 GND.n2617 GND.n2616 585
R6956 GND.n2619 GND.n2565 585
R6957 GND.n2621 GND.n2620 585
R6958 GND.n2622 GND.n2560 585
R6959 GND.n2624 GND.n2623 585
R6960 GND.n2626 GND.n2559 585
R6961 GND.n2627 GND.n2068 585
R6962 GND.n2630 GND.n2557 585
R6963 GND.n2632 GND.n2631 585
R6964 GND.n2633 GND.n2553 585
R6965 GND.n2635 GND.n2634 585
R6966 GND.n2637 GND.n2551 585
R6967 GND.n2639 GND.n2638 585
R6968 GND.n2640 GND.n2550 585
R6969 GND.n2642 GND.n2641 585
R6970 GND.n2644 GND.n2548 585
R6971 GND.n2646 GND.n2645 585
R6972 GND.n2647 GND.n2547 585
R6973 GND.n2649 GND.n2648 585
R6974 GND.n2651 GND.n2545 585
R6975 GND.n2653 GND.n2652 585
R6976 GND.n2654 GND.n2544 585
R6977 GND.n2656 GND.n2655 585
R6978 GND.n2658 GND.n2542 585
R6979 GND.n2660 GND.n2659 585
R6980 GND.n2661 GND.n2541 585
R6981 GND.n2663 GND.n2662 585
R6982 GND.n2665 GND.n2539 585
R6983 GND.n2667 GND.n2666 585
R6984 GND.n2668 GND.n2508 585
R6985 GND.n2670 GND.n2669 585
R6986 GND.n2670 GND.n2068 585
R6987 GND.n2584 GND.n2579 585
R6988 GND.n2584 GND.n2067 585
R6989 GND.n2583 GND.n2582 585
R6990 GND.n2583 GND.n2077 585
R6991 GND.n2581 GND.n2499 585
R6992 GND.n2499 GND.n2074 585
R6993 GND.n2678 GND.n2498 585
R6994 GND.n2678 GND.n2677 585
R6995 GND.n2680 GND.n2679 585
R6996 GND.n2679 GND.n2084 585
R6997 GND.n2681 GND.n2494 585
R6998 GND.n2494 GND.n2083 585
R6999 GND.n2683 GND.n2682 585
R7000 GND.n2684 GND.n2683 585
R7001 GND.n2497 GND.n2493 585
R7002 GND.n2686 GND.n2493 585
R7003 GND.n2496 GND.n2495 585
R7004 GND.n2495 GND.n2090 585
R7005 GND.n2486 GND.n2485 585
R7006 GND.n2488 GND.n2486 585
R7007 GND.n2695 GND.n2694 585
R7008 GND.n2694 GND.n2693 585
R7009 GND.n2696 GND.n2482 585
R7010 GND.n2482 GND.n2097 585
R7011 GND.n2698 GND.n2697 585
R7012 GND.n2699 GND.n2698 585
R7013 GND.n2484 GND.n2481 585
R7014 GND.n2481 GND.n2105 585
R7015 GND.n2483 GND.n2472 585
R7016 GND.n2472 GND.n2103 585
R7017 GND.n2707 GND.n2471 585
R7018 GND.n2707 GND.n2706 585
R7019 GND.n2709 GND.n2708 585
R7020 GND.n2708 GND.n2112 585
R7021 GND.n2710 GND.n2468 585
R7022 GND.n2468 GND.n2111 585
R7023 GND.n2712 GND.n2711 585
R7024 GND.n2713 GND.n2712 585
R7025 GND.n2470 GND.n2467 585
R7026 GND.n2467 GND.n2120 585
R7027 GND.n2469 GND.n2457 585
R7028 GND.n2457 GND.n2118 585
R7029 GND.n2721 GND.n2456 585
R7030 GND.n2721 GND.n2720 585
R7031 GND.n2723 GND.n2722 585
R7032 GND.n2722 GND.n2127 585
R7033 GND.n2724 GND.n2453 585
R7034 GND.n2453 GND.n2126 585
R7035 GND.n2726 GND.n2725 585
R7036 GND.n2727 GND.n2726 585
R7037 GND.n2455 GND.n2452 585
R7038 GND.n2729 GND.n2452 585
R7039 GND.n2454 GND.n2444 585
R7040 GND.n2444 GND.n2133 585
R7041 GND.n2736 GND.n2443 585
R7042 GND.n2736 GND.n2735 585
R7043 GND.n2738 GND.n2737 585
R7044 GND.n2737 GND.n2141 585
R7045 GND.n2739 GND.n2440 585
R7046 GND.n2440 GND.n2140 585
R7047 GND.n2741 GND.n2740 585
R7048 GND.n2743 GND.n2741 585
R7049 GND.n2442 GND.n2439 585
R7050 GND.n2439 GND.n2148 585
R7051 GND.n2441 GND.n2430 585
R7052 GND.n2433 GND.n2430 585
R7053 GND.n2751 GND.n2429 585
R7054 GND.n2751 GND.n2750 585
R7055 GND.n2753 GND.n2752 585
R7056 GND.n2752 GND.n2155 585
R7057 GND.n2754 GND.n2426 585
R7058 GND.n2426 GND.n2154 585
R7059 GND.n2756 GND.n2755 585
R7060 GND.n2758 GND.n2756 585
R7061 GND.n2428 GND.n2425 585
R7062 GND.n2425 GND.n2163 585
R7063 GND.n2427 GND.n2417 585
R7064 GND.n2417 GND.n2161 585
R7065 GND.n2766 GND.n2416 585
R7066 GND.n2766 GND.n2765 585
R7067 GND.n2768 GND.n2767 585
R7068 GND.n2767 GND.n2170 585
R7069 GND.n2769 GND.n2413 585
R7070 GND.n2413 GND.n2169 585
R7071 GND.n2771 GND.n2770 585
R7072 GND.n2773 GND.n2771 585
R7073 GND.n2415 GND.n2412 585
R7074 GND.n2412 GND.n2177 585
R7075 GND.n2414 GND.n2390 585
R7076 GND.n2394 GND.n2390 585
R7077 GND.n2781 GND.n2391 585
R7078 GND.n2781 GND.n2780 585
R7079 GND.n2782 GND.n2389 585
R7080 GND.n2782 GND.n2184 585
R7081 GND.n2784 GND.n2783 585
R7082 GND.n2783 GND.n2183 585
R7083 GND.n2785 GND.n2388 585
R7084 GND.n2405 GND.n2388 585
R7085 GND.n2787 GND.n2786 585
R7086 GND.n2787 GND.n2192 585
R7087 GND.n2788 GND.n2387 585
R7088 GND.n2788 GND.n2190 585
R7089 GND.n2790 GND.n2789 585
R7090 GND.n2789 GND.n2200 585
R7091 GND.n2791 GND.n2383 585
R7092 GND.n2383 GND.n2198 585
R7093 GND.n2793 GND.n2792 585
R7094 GND.n2794 GND.n2793 585
R7095 GND.n2386 GND.n2382 585
R7096 GND.n2382 GND.n2208 585
R7097 GND.n2385 GND.n2384 585
R7098 GND.n2384 GND.n2206 585
R7099 GND.n2373 GND.n2372 585
R7100 GND.n2375 GND.n2373 585
R7101 GND.n2804 GND.n2803 585
R7102 GND.n2803 GND.n2802 585
R7103 GND.n2805 GND.n2369 585
R7104 GND.n2369 GND.n2214 585
R7105 GND.n2807 GND.n2806 585
R7106 GND.n2808 GND.n2807 585
R7107 GND.n2371 GND.n2368 585
R7108 GND.n2368 GND.n2222 585
R7109 GND.n2370 GND.n2358 585
R7110 GND.n2358 GND.n2220 585
R7111 GND.n2816 GND.n2357 585
R7112 GND.n2816 GND.n2815 585
R7113 GND.n2818 GND.n2817 585
R7114 GND.n2817 GND.n2229 585
R7115 GND.n2819 GND.n2354 585
R7116 GND.n2354 GND.n2228 585
R7117 GND.n2821 GND.n2820 585
R7118 GND.n2822 GND.n2821 585
R7119 GND.n2356 GND.n2353 585
R7120 GND.n2824 GND.n2353 585
R7121 GND.n2355 GND.n2345 585
R7122 GND.n2345 GND.n2235 585
R7123 GND.n2831 GND.n2344 585
R7124 GND.n2831 GND.n2830 585
R7125 GND.n2833 GND.n2832 585
R7126 GND.n2832 GND.n2243 585
R7127 GND.n2834 GND.n2341 585
R7128 GND.n2341 GND.n2242 585
R7129 GND.n2836 GND.n2835 585
R7130 GND.n2837 GND.n2836 585
R7131 GND.n2343 GND.n2340 585
R7132 GND.n2340 GND.n2251 585
R7133 GND.n2342 GND.n2330 585
R7134 GND.n2330 GND.n2249 585
R7135 GND.n2845 GND.n2331 585
R7136 GND.n2845 GND.n2844 585
R7137 GND.n2846 GND.n2329 585
R7138 GND.n2846 GND.n2258 585
R7139 GND.n2848 GND.n2847 585
R7140 GND.n2847 GND.n2257 585
R7141 GND.n4952 GND.n4951 585
R7142 GND.n4953 GND.n4952 585
R7143 GND.n1297 GND.n1295 585
R7144 GND.n3869 GND.n1295 585
R7145 GND.n3865 GND.n3864 585
R7146 GND.n3866 GND.n3865 585
R7147 GND.n2976 GND.n2975 585
R7148 GND.n3846 GND.n2975 585
R7149 GND.n3860 GND.n3859 585
R7150 GND.n3859 GND.n3858 585
R7151 GND.n2979 GND.n2978 585
R7152 GND.n3854 GND.n2979 585
R7153 GND.n3837 GND.n2997 585
R7154 GND.n2997 GND.n2996 585
R7155 GND.n3839 GND.n3838 585
R7156 GND.n3840 GND.n3839 585
R7157 GND.n2998 GND.n2994 585
R7158 GND.n3827 GND.n2994 585
R7159 GND.n3832 GND.n3831 585
R7160 GND.n3831 GND.n3830 585
R7161 GND.n3001 GND.n3000 585
R7162 GND.n3824 GND.n3001 585
R7163 GND.n3812 GND.n3020 585
R7164 GND.n3020 GND.n3019 585
R7165 GND.n3814 GND.n3813 585
R7166 GND.n3815 GND.n3814 585
R7167 GND.n3021 GND.n3018 585
R7168 GND.n3802 GND.n3018 585
R7169 GND.n3807 GND.n3806 585
R7170 GND.n3806 GND.n3805 585
R7171 GND.n3024 GND.n3023 585
R7172 GND.n3800 GND.n3024 585
R7173 GND.n3788 GND.n3043 585
R7174 GND.n3043 GND.n3042 585
R7175 GND.n3790 GND.n3789 585
R7176 GND.n3791 GND.n3790 585
R7177 GND.n3044 GND.n3041 585
R7178 GND.n3778 GND.n3041 585
R7179 GND.n3783 GND.n3782 585
R7180 GND.n3782 GND.n3781 585
R7181 GND.n3047 GND.n3046 585
R7182 GND.n3775 GND.n3047 585
R7183 GND.n3763 GND.n3066 585
R7184 GND.n3066 GND.n3065 585
R7185 GND.n3765 GND.n3764 585
R7186 GND.n3766 GND.n3765 585
R7187 GND.n3067 GND.n3064 585
R7188 GND.n3726 GND.n3064 585
R7189 GND.n3721 GND.n3720 585
R7190 GND.n3722 GND.n3721 585
R7191 GND.n3719 GND.n3718 585
R7192 GND.n3719 GND.n3107 585
R7193 GND.n3717 GND.n3100 585
R7194 GND.n3735 GND.n3100 585
R7195 GND.n3740 GND.n3739 585
R7196 GND.n3739 GND.n3738 585
R7197 GND.n3742 GND.n3741 585
R7198 GND.n3743 GND.n3742 585
R7199 GND.n3099 GND.n3098 585
R7200 GND.n3099 GND.n3092 585
R7201 GND.n3097 GND.n3073 585
R7202 GND.n3097 GND.n3085 585
R7203 GND.n3077 GND.n3074 585
R7204 GND.n3752 GND.n3077 585
R7205 GND.n3758 GND.n3757 585
R7206 GND.n3757 GND.n3756 585
R7207 GND.n3076 GND.n3075 585
R7208 GND.n3216 GND.n3076 585
R7209 GND.n3693 GND.n3692 585
R7210 GND.n3694 GND.n3693 585
R7211 GND.n3220 GND.n3219 585
R7212 GND.n3682 GND.n3219 585
R7213 GND.n3688 GND.n3687 585
R7214 GND.n3687 GND.n3686 585
R7215 GND.n3223 GND.n3222 585
R7216 GND.n3680 GND.n3223 585
R7217 GND.n3668 GND.n3241 585
R7218 GND.n3241 GND.n3240 585
R7219 GND.n3670 GND.n3669 585
R7220 GND.n3671 GND.n3670 585
R7221 GND.n3242 GND.n3238 585
R7222 GND.n3658 GND.n3238 585
R7223 GND.n3663 GND.n3662 585
R7224 GND.n3662 GND.n3661 585
R7225 GND.n3245 GND.n3244 585
R7226 GND.n3655 GND.n3245 585
R7227 GND.n3643 GND.n3264 585
R7228 GND.n3264 GND.n3263 585
R7229 GND.n3645 GND.n3644 585
R7230 GND.n3646 GND.n3645 585
R7231 GND.n3265 GND.n3262 585
R7232 GND.n3633 GND.n3262 585
R7233 GND.n3638 GND.n3637 585
R7234 GND.n3637 GND.n3636 585
R7235 GND.n3268 GND.n3267 585
R7236 GND.n3631 GND.n3268 585
R7237 GND.n3619 GND.n3287 585
R7238 GND.n3287 GND.n3286 585
R7239 GND.n3621 GND.n3620 585
R7240 GND.n3622 GND.n3621 585
R7241 GND.n3288 GND.n3285 585
R7242 GND.n3609 GND.n3285 585
R7243 GND.n3614 GND.n3613 585
R7244 GND.n3613 GND.n3612 585
R7245 GND.n1173 GND.n1172 585
R7246 GND.n3291 GND.n1173 585
R7247 GND.n5040 GND.n5039 585
R7248 GND.n5039 GND.n5038 585
R7249 GND.n5041 GND.n1168 585
R7250 GND.n3528 GND.n1168 585
R7251 GND.n5043 GND.n5042 585
R7252 GND.n5044 GND.n5043 585
R7253 GND.n3361 GND.n1167 585
R7254 GND.n3364 GND.n3363 585
R7255 GND.n3359 GND.n3358 585
R7256 GND.n3358 GND.n1162 585
R7257 GND.n3369 GND.n3368 585
R7258 GND.n3371 GND.n3357 585
R7259 GND.n3374 GND.n3373 585
R7260 GND.n3355 GND.n3354 585
R7261 GND.n3379 GND.n3378 585
R7262 GND.n3381 GND.n3353 585
R7263 GND.n3384 GND.n3383 585
R7264 GND.n3351 GND.n3348 585
R7265 GND.n3389 GND.n3388 585
R7266 GND.n3391 GND.n3347 585
R7267 GND.n3394 GND.n3393 585
R7268 GND.n3345 GND.n3344 585
R7269 GND.n3399 GND.n3398 585
R7270 GND.n3401 GND.n3343 585
R7271 GND.n3404 GND.n3403 585
R7272 GND.n3341 GND.n3340 585
R7273 GND.n3409 GND.n3408 585
R7274 GND.n3411 GND.n3339 585
R7275 GND.n3414 GND.n3413 585
R7276 GND.n3337 GND.n3336 585
R7277 GND.n3421 GND.n3420 585
R7278 GND.n3423 GND.n3335 585
R7279 GND.n3426 GND.n3425 585
R7280 GND.n3333 GND.n3332 585
R7281 GND.n3431 GND.n3430 585
R7282 GND.n3433 GND.n3331 585
R7283 GND.n3436 GND.n3435 585
R7284 GND.n3329 GND.n3328 585
R7285 GND.n3441 GND.n3440 585
R7286 GND.n3443 GND.n3327 585
R7287 GND.n3446 GND.n3445 585
R7288 GND.n3325 GND.n3324 585
R7289 GND.n3454 GND.n3453 585
R7290 GND.n3456 GND.n3323 585
R7291 GND.n3459 GND.n3458 585
R7292 GND.n3321 GND.n3320 585
R7293 GND.n3464 GND.n3463 585
R7294 GND.n3466 GND.n3319 585
R7295 GND.n3469 GND.n3468 585
R7296 GND.n3317 GND.n3316 585
R7297 GND.n3474 GND.n3473 585
R7298 GND.n3476 GND.n3315 585
R7299 GND.n3479 GND.n3478 585
R7300 GND.n3313 GND.n3312 585
R7301 GND.n3484 GND.n3483 585
R7302 GND.n3486 GND.n3311 585
R7303 GND.n3488 GND.n3487 585
R7304 GND.n3487 GND.n1162 585
R7305 GND.n4872 GND.n1289 585
R7306 GND.n4873 GND.n1399 585
R7307 GND.n4874 GND.n1395 585
R7308 GND.n1393 GND.n1391 585
R7309 GND.n4878 GND.n1390 585
R7310 GND.n4879 GND.n1388 585
R7311 GND.n4880 GND.n1387 585
R7312 GND.n1385 GND.n1383 585
R7313 GND.n4884 GND.n1382 585
R7314 GND.n4885 GND.n1380 585
R7315 GND.n4886 GND.n1379 585
R7316 GND.n1377 GND.n1375 585
R7317 GND.n4890 GND.n1374 585
R7318 GND.n4891 GND.n1372 585
R7319 GND.n4893 GND.n1369 585
R7320 GND.n1367 GND.n1365 585
R7321 GND.n4897 GND.n1364 585
R7322 GND.n4898 GND.n1362 585
R7323 GND.n4899 GND.n1361 585
R7324 GND.n1359 GND.n1357 585
R7325 GND.n4903 GND.n1356 585
R7326 GND.n4904 GND.n1354 585
R7327 GND.n4905 GND.n1353 585
R7328 GND.n1349 GND.n1348 585
R7329 GND.n4910 GND.n4909 585
R7330 GND.n4912 GND.n1347 585
R7331 GND.n4913 GND.n1346 585
R7332 GND.n4917 GND.n4916 585
R7333 GND.n1331 GND.n1326 585
R7334 GND.n4921 GND.n1325 585
R7335 GND.n4922 GND.n1324 585
R7336 GND.n4923 GND.n1323 585
R7337 GND.n1334 GND.n1321 585
R7338 GND.n4927 GND.n1320 585
R7339 GND.n4928 GND.n1319 585
R7340 GND.n4929 GND.n1318 585
R7341 GND.n1337 GND.n1316 585
R7342 GND.n4933 GND.n1315 585
R7343 GND.n4934 GND.n1314 585
R7344 GND.n4935 GND.n1310 585
R7345 GND.n4936 GND.n1309 585
R7346 GND.n1340 GND.n1307 585
R7347 GND.n4940 GND.n1306 585
R7348 GND.n4941 GND.n1305 585
R7349 GND.n4942 GND.n1304 585
R7350 GND.n1343 GND.n1302 585
R7351 GND.n4946 GND.n1301 585
R7352 GND.n4947 GND.n1300 585
R7353 GND.n4948 GND.n1296 585
R7354 GND.n1346 GND.n1296 585
R7355 GND.n4955 GND.n4954 585
R7356 GND.n4954 GND.n4953 585
R7357 GND.n4956 GND.n1288 585
R7358 GND.n3869 GND.n1288 585
R7359 GND.n2974 GND.n1283 585
R7360 GND.n3866 GND.n2974 585
R7361 GND.n4960 GND.n1282 585
R7362 GND.n3846 GND.n1282 585
R7363 GND.n4961 GND.n1281 585
R7364 GND.n3858 GND.n1281 585
R7365 GND.n4962 GND.n1280 585
R7366 GND.n3854 GND.n1280 585
R7367 GND.n2995 GND.n1275 585
R7368 GND.n2996 GND.n2995 585
R7369 GND.n4966 GND.n1274 585
R7370 GND.n3840 GND.n1274 585
R7371 GND.n4967 GND.n1273 585
R7372 GND.n3827 GND.n1273 585
R7373 GND.n4968 GND.n1272 585
R7374 GND.n3830 GND.n1272 585
R7375 GND.n3007 GND.n1267 585
R7376 GND.n3824 GND.n3007 585
R7377 GND.n4972 GND.n1266 585
R7378 GND.n3019 GND.n1266 585
R7379 GND.n4973 GND.n1265 585
R7380 GND.n3815 GND.n1265 585
R7381 GND.n4974 GND.n1264 585
R7382 GND.n3802 GND.n1264 585
R7383 GND.n3026 GND.n1259 585
R7384 GND.n3805 GND.n3026 585
R7385 GND.n4978 GND.n1258 585
R7386 GND.n3800 GND.n1258 585
R7387 GND.n4979 GND.n1257 585
R7388 GND.n3042 GND.n1257 585
R7389 GND.n4980 GND.n1256 585
R7390 GND.n3791 GND.n1256 585
R7391 GND.n3777 GND.n1251 585
R7392 GND.n3778 GND.n3777 585
R7393 GND.n4984 GND.n1250 585
R7394 GND.n3781 GND.n1250 585
R7395 GND.n4985 GND.n1249 585
R7396 GND.n3775 GND.n1249 585
R7397 GND.n4986 GND.n1248 585
R7398 GND.n3065 GND.n1248 585
R7399 GND.n3061 GND.n1243 585
R7400 GND.n3766 GND.n3061 585
R7401 GND.n4990 GND.n1242 585
R7402 GND.n3726 GND.n1242 585
R7403 GND.n4991 GND.n1241 585
R7404 GND.n3722 GND.n1241 585
R7405 GND.n4992 GND.n1240 585
R7406 GND.n3107 GND.n1240 585
R7407 GND.n3105 GND.n1235 585
R7408 GND.n3735 GND.n3105 585
R7409 GND.n4996 GND.n1234 585
R7410 GND.n3738 GND.n1234 585
R7411 GND.n4997 GND.n1233 585
R7412 GND.n3743 GND.n1233 585
R7413 GND.n4998 GND.n1232 585
R7414 GND.n3092 GND.n1232 585
R7415 GND.n3084 GND.n1227 585
R7416 GND.n3085 GND.n3084 585
R7417 GND.n5002 GND.n1226 585
R7418 GND.n3752 GND.n1226 585
R7419 GND.n5003 GND.n1225 585
R7420 GND.n3756 GND.n1225 585
R7421 GND.n5004 GND.n1224 585
R7422 GND.n3216 GND.n1224 585
R7423 GND.n3215 GND.n1219 585
R7424 GND.n3694 GND.n3215 585
R7425 GND.n5008 GND.n1218 585
R7426 GND.n3682 GND.n1218 585
R7427 GND.n5009 GND.n1217 585
R7428 GND.n3686 GND.n1217 585
R7429 GND.n5010 GND.n1216 585
R7430 GND.n3680 GND.n1216 585
R7431 GND.n3239 GND.n1211 585
R7432 GND.n3240 GND.n3239 585
R7433 GND.n5014 GND.n1210 585
R7434 GND.n3671 GND.n1210 585
R7435 GND.n5015 GND.n1209 585
R7436 GND.n3658 GND.n1209 585
R7437 GND.n5016 GND.n1208 585
R7438 GND.n3661 GND.n1208 585
R7439 GND.n3251 GND.n1203 585
R7440 GND.n3655 GND.n3251 585
R7441 GND.n5020 GND.n1202 585
R7442 GND.n3263 GND.n1202 585
R7443 GND.n5021 GND.n1201 585
R7444 GND.n3646 GND.n1201 585
R7445 GND.n5022 GND.n1200 585
R7446 GND.n3633 GND.n1200 585
R7447 GND.n3270 GND.n1195 585
R7448 GND.n3636 GND.n3270 585
R7449 GND.n5026 GND.n1194 585
R7450 GND.n3631 GND.n1194 585
R7451 GND.n5027 GND.n1193 585
R7452 GND.n3286 GND.n1193 585
R7453 GND.n5028 GND.n1192 585
R7454 GND.n3622 GND.n1192 585
R7455 GND.n3608 GND.n1187 585
R7456 GND.n3609 GND.n3608 585
R7457 GND.n5032 GND.n1186 585
R7458 GND.n3612 GND.n1186 585
R7459 GND.n5033 GND.n1185 585
R7460 GND.n3291 GND.n1185 585
R7461 GND.n5034 GND.n1175 585
R7462 GND.n5038 GND.n1175 585
R7463 GND.n3527 GND.n1184 585
R7464 GND.n3528 GND.n3527 585
R7465 GND.n3491 GND.n1163 585
R7466 GND.n5044 GND.n1163 585
R7467 GND.n6259 GND.n290 585
R7468 GND.n6159 GND.n290 585
R7469 GND.n6261 GND.n6260 585
R7470 GND.n6262 GND.n6261 585
R7471 GND.n275 GND.n274 585
R7472 GND.n4438 GND.n275 585
R7473 GND.n6270 GND.n6269 585
R7474 GND.n6269 GND.n6268 585
R7475 GND.n6271 GND.n269 585
R7476 GND.n4444 GND.n269 585
R7477 GND.n6273 GND.n6272 585
R7478 GND.n6274 GND.n6273 585
R7479 GND.n255 GND.n254 585
R7480 GND.n4450 GND.n255 585
R7481 GND.n6282 GND.n6281 585
R7482 GND.n6281 GND.n6280 585
R7483 GND.n6283 GND.n249 585
R7484 GND.n4380 GND.n249 585
R7485 GND.n6285 GND.n6284 585
R7486 GND.n6286 GND.n6285 585
R7487 GND.n234 GND.n233 585
R7488 GND.n4371 GND.n234 585
R7489 GND.n6294 GND.n6293 585
R7490 GND.n6293 GND.n6292 585
R7491 GND.n6295 GND.n228 585
R7492 GND.n4365 GND.n228 585
R7493 GND.n6297 GND.n6296 585
R7494 GND.n6298 GND.n6297 585
R7495 GND.n213 GND.n212 585
R7496 GND.n4357 GND.n213 585
R7497 GND.n6306 GND.n6305 585
R7498 GND.n6305 GND.n6304 585
R7499 GND.n6307 GND.n207 585
R7500 GND.n4351 GND.n207 585
R7501 GND.n6309 GND.n6308 585
R7502 GND.n6310 GND.n6309 585
R7503 GND.n193 GND.n192 585
R7504 GND.n4472 GND.n193 585
R7505 GND.n6318 GND.n6317 585
R7506 GND.n6317 GND.n6316 585
R7507 GND.n6319 GND.n188 585
R7508 GND.n4478 GND.n188 585
R7509 GND.n6321 GND.n6320 585
R7510 GND.n6322 GND.n6321 585
R7511 GND.n171 GND.n169 585
R7512 GND.n4484 GND.n171 585
R7513 GND.n6330 GND.n6329 585
R7514 GND.n6329 GND.n6328 585
R7515 GND.n170 GND.n168 585
R7516 GND.n4490 GND.n170 585
R7517 GND.n4498 GND.n4497 585
R7518 GND.n4499 GND.n4498 585
R7519 GND.n160 GND.n158 585
R7520 GND.n1890 GND.n158 585
R7521 GND.n6334 GND.n6333 585
R7522 GND.n6335 GND.n6334 585
R7523 GND.n159 GND.n157 585
R7524 GND.n1801 GND.n157 585
R7525 GND.n4510 GND.n1798 585
R7526 GND.n4510 GND.n4509 585
R7527 GND.n4511 GND.n166 585
R7528 GND.n4512 GND.n4511 585
R7529 GND.n1783 GND.n1782 585
R7530 GND.n4247 GND.n1783 585
R7531 GND.n4520 GND.n4519 585
R7532 GND.n4519 GND.n4518 585
R7533 GND.n4521 GND.n1779 585
R7534 GND.n4235 GND.n1779 585
R7535 GND.n4523 GND.n4522 585
R7536 GND.n4524 GND.n4523 585
R7537 GND.n1764 GND.n1763 585
R7538 GND.n4228 GND.n1764 585
R7539 GND.n4532 GND.n4531 585
R7540 GND.n4531 GND.n4530 585
R7541 GND.n4533 GND.n1758 585
R7542 GND.n4220 GND.n1758 585
R7543 GND.n4535 GND.n4534 585
R7544 GND.n4536 GND.n4535 585
R7545 GND.n1743 GND.n1742 585
R7546 GND.n4213 GND.n1743 585
R7547 GND.n4544 GND.n4543 585
R7548 GND.n4543 GND.n4542 585
R7549 GND.n4545 GND.n1737 585
R7550 GND.n4205 GND.n1737 585
R7551 GND.n4547 GND.n4546 585
R7552 GND.n4548 GND.n4547 585
R7553 GND.n1722 GND.n1721 585
R7554 GND.n4198 GND.n1722 585
R7555 GND.n4556 GND.n4555 585
R7556 GND.n4555 GND.n4554 585
R7557 GND.n4557 GND.n1716 585
R7558 GND.n4190 GND.n1716 585
R7559 GND.n4559 GND.n4558 585
R7560 GND.n4560 GND.n4559 585
R7561 GND.n1701 GND.n1700 585
R7562 GND.n4183 GND.n1701 585
R7563 GND.n4568 GND.n4567 585
R7564 GND.n4567 GND.n4566 585
R7565 GND.n4569 GND.n1695 585
R7566 GND.n4175 GND.n1695 585
R7567 GND.n4571 GND.n4570 585
R7568 GND.n4572 GND.n4571 585
R7569 GND.n1679 GND.n1678 585
R7570 GND.n4168 GND.n1679 585
R7571 GND.n4580 GND.n4579 585
R7572 GND.n4579 GND.n4578 585
R7573 GND.n4581 GND.n1672 585
R7574 GND.n4160 GND.n1672 585
R7575 GND.n4583 GND.n4582 585
R7576 GND.n4584 GND.n4583 585
R7577 GND.n1673 GND.n1599 585
R7578 GND.n4587 GND.n1599 585
R7579 GND.n4686 GND.n4685 585
R7580 GND.n4684 GND.n1598 585
R7581 GND.n4683 GND.n1597 585
R7582 GND.n4688 GND.n1597 585
R7583 GND.n4682 GND.n4681 585
R7584 GND.n4680 GND.n4679 585
R7585 GND.n4678 GND.n4677 585
R7586 GND.n4676 GND.n4675 585
R7587 GND.n4674 GND.n4673 585
R7588 GND.n4672 GND.n4671 585
R7589 GND.n4670 GND.n4669 585
R7590 GND.n4668 GND.n1610 585
R7591 GND.n4667 GND.n4666 585
R7592 GND.n4665 GND.n4664 585
R7593 GND.n4663 GND.n4662 585
R7594 GND.n4661 GND.n4660 585
R7595 GND.n4659 GND.n4658 585
R7596 GND.n4657 GND.n4656 585
R7597 GND.n4655 GND.n4654 585
R7598 GND.n4653 GND.n4652 585
R7599 GND.n4651 GND.n4650 585
R7600 GND.n4649 GND.n4648 585
R7601 GND.n4647 GND.n4646 585
R7602 GND.n4644 GND.n4643 585
R7603 GND.n4642 GND.n4641 585
R7604 GND.n4640 GND.n4639 585
R7605 GND.n4638 GND.n4637 585
R7606 GND.n4636 GND.n4635 585
R7607 GND.n4634 GND.n4633 585
R7608 GND.n4632 GND.n4631 585
R7609 GND.n4630 GND.n4629 585
R7610 GND.n4628 GND.n4627 585
R7611 GND.n4626 GND.n4625 585
R7612 GND.n4624 GND.n4623 585
R7613 GND.n4622 GND.n4621 585
R7614 GND.n4619 GND.n4618 585
R7615 GND.n4617 GND.n4616 585
R7616 GND.n4615 GND.n4614 585
R7617 GND.n4613 GND.n4612 585
R7618 GND.n4611 GND.n4610 585
R7619 GND.n4609 GND.n4608 585
R7620 GND.n4607 GND.n4606 585
R7621 GND.n4605 GND.n4604 585
R7622 GND.n4603 GND.n4602 585
R7623 GND.n4601 GND.n4600 585
R7624 GND.n4599 GND.n4598 585
R7625 GND.n4597 GND.n4596 585
R7626 GND.n1658 GND.n1655 585
R7627 GND.n4592 GND.n1589 585
R7628 GND.n4688 GND.n1589 585
R7629 GND.n385 GND.n379 585
R7630 GND.n6166 GND.n376 585
R7631 GND.n6168 GND.n6167 585
R7632 GND.n6170 GND.n374 585
R7633 GND.n6172 GND.n6171 585
R7634 GND.n6173 GND.n369 585
R7635 GND.n6175 GND.n6174 585
R7636 GND.n6177 GND.n367 585
R7637 GND.n6179 GND.n6178 585
R7638 GND.n6180 GND.n362 585
R7639 GND.n6182 GND.n6181 585
R7640 GND.n6184 GND.n360 585
R7641 GND.n6186 GND.n6185 585
R7642 GND.n6187 GND.n355 585
R7643 GND.n6192 GND.n6191 585
R7644 GND.n6194 GND.n353 585
R7645 GND.n6196 GND.n6195 585
R7646 GND.n6197 GND.n348 585
R7647 GND.n6199 GND.n6198 585
R7648 GND.n6201 GND.n346 585
R7649 GND.n6203 GND.n6202 585
R7650 GND.n6204 GND.n342 585
R7651 GND.n6206 GND.n6205 585
R7652 GND.n6208 GND.n340 585
R7653 GND.n6210 GND.n6209 585
R7654 GND.n335 GND.n334 585
R7655 GND.n6215 GND.n6214 585
R7656 GND.n6217 GND.n332 585
R7657 GND.n6219 GND.n6218 585
R7658 GND.n6220 GND.n327 585
R7659 GND.n6222 GND.n6221 585
R7660 GND.n6224 GND.n325 585
R7661 GND.n6226 GND.n6225 585
R7662 GND.n6227 GND.n320 585
R7663 GND.n6229 GND.n6228 585
R7664 GND.n6231 GND.n318 585
R7665 GND.n6233 GND.n6232 585
R7666 GND.n6234 GND.n313 585
R7667 GND.n6236 GND.n6235 585
R7668 GND.n6238 GND.n311 585
R7669 GND.n6240 GND.n6239 585
R7670 GND.n6241 GND.n304 585
R7671 GND.n6243 GND.n6242 585
R7672 GND.n6245 GND.n302 585
R7673 GND.n6247 GND.n6246 585
R7674 GND.n6248 GND.n297 585
R7675 GND.n6250 GND.n6249 585
R7676 GND.n6252 GND.n296 585
R7677 GND.n6253 GND.n294 585
R7678 GND.n6256 GND.n6255 585
R7679 GND.n6161 GND.n6160 585
R7680 GND.n6160 GND.n6159 585
R7681 GND.n383 GND.n287 585
R7682 GND.n6262 GND.n287 585
R7683 GND.n4440 GND.n4439 585
R7684 GND.n4439 GND.n4438 585
R7685 GND.n4441 GND.n277 585
R7686 GND.n6268 GND.n277 585
R7687 GND.n4443 GND.n4442 585
R7688 GND.n4444 GND.n4443 585
R7689 GND.n4385 GND.n266 585
R7690 GND.n6274 GND.n266 585
R7691 GND.n4384 GND.n4328 585
R7692 GND.n4450 GND.n4328 585
R7693 GND.n4383 GND.n257 585
R7694 GND.n6280 GND.n257 585
R7695 GND.n4382 GND.n4381 585
R7696 GND.n4381 GND.n4380 585
R7697 GND.n4334 GND.n246 585
R7698 GND.n6286 GND.n246 585
R7699 GND.n4370 GND.n4369 585
R7700 GND.n4371 GND.n4370 585
R7701 GND.n4368 GND.n236 585
R7702 GND.n6292 GND.n236 585
R7703 GND.n4367 GND.n4366 585
R7704 GND.n4366 GND.n4365 585
R7705 GND.n4339 GND.n225 585
R7706 GND.n6298 GND.n225 585
R7707 GND.n4356 GND.n4355 585
R7708 GND.n4357 GND.n4356 585
R7709 GND.n4354 GND.n215 585
R7710 GND.n6304 GND.n215 585
R7711 GND.n4353 GND.n4352 585
R7712 GND.n4352 GND.n4351 585
R7713 GND.n4345 GND.n204 585
R7714 GND.n6310 GND.n204 585
R7715 GND.n4344 GND.n4275 585
R7716 GND.n4472 GND.n4275 585
R7717 GND.n4269 GND.n195 585
R7718 GND.n6316 GND.n195 585
R7719 GND.n4480 GND.n4479 585
R7720 GND.n4479 GND.n4478 585
R7721 GND.n4481 GND.n185 585
R7722 GND.n6322 GND.n185 585
R7723 GND.n4483 GND.n4482 585
R7724 GND.n4484 GND.n4483 585
R7725 GND.n4261 GND.n173 585
R7726 GND.n6328 GND.n173 585
R7727 GND.n4492 GND.n4491 585
R7728 GND.n4491 GND.n4490 585
R7729 GND.n4493 GND.n1891 585
R7730 GND.n4499 GND.n1891 585
R7731 GND.n4260 GND.n4259 585
R7732 GND.n4259 GND.n1890 585
R7733 GND.n4258 GND.n154 585
R7734 GND.n6335 GND.n154 585
R7735 GND.n1899 GND.n1898 585
R7736 GND.n1898 GND.n1801 585
R7737 GND.n4251 GND.n1799 585
R7738 GND.n4509 GND.n1799 585
R7739 GND.n4250 GND.n1795 585
R7740 GND.n4512 GND.n1795 585
R7741 GND.n4249 GND.n4248 585
R7742 GND.n4248 GND.n4247 585
R7743 GND.n1900 GND.n1785 585
R7744 GND.n4518 GND.n1785 585
R7745 GND.n4234 GND.n4233 585
R7746 GND.n4235 GND.n4234 585
R7747 GND.n4231 GND.n1776 585
R7748 GND.n4524 GND.n1776 585
R7749 GND.n4230 GND.n4229 585
R7750 GND.n4229 GND.n4228 585
R7751 GND.n1904 GND.n1766 585
R7752 GND.n4530 GND.n1766 585
R7753 GND.n4219 GND.n4218 585
R7754 GND.n4220 GND.n4219 585
R7755 GND.n4216 GND.n1755 585
R7756 GND.n4536 GND.n1755 585
R7757 GND.n4215 GND.n4214 585
R7758 GND.n4214 GND.n4213 585
R7759 GND.n1908 GND.n1745 585
R7760 GND.n4542 GND.n1745 585
R7761 GND.n4204 GND.n4203 585
R7762 GND.n4205 GND.n4204 585
R7763 GND.n4201 GND.n1734 585
R7764 GND.n4548 GND.n1734 585
R7765 GND.n4200 GND.n4199 585
R7766 GND.n4199 GND.n4198 585
R7767 GND.n1912 GND.n1724 585
R7768 GND.n4554 GND.n1724 585
R7769 GND.n4189 GND.n4188 585
R7770 GND.n4190 GND.n4189 585
R7771 GND.n4186 GND.n1713 585
R7772 GND.n4560 GND.n1713 585
R7773 GND.n4185 GND.n4184 585
R7774 GND.n4184 GND.n4183 585
R7775 GND.n1916 GND.n1703 585
R7776 GND.n4566 GND.n1703 585
R7777 GND.n4174 GND.n4173 585
R7778 GND.n4175 GND.n4174 585
R7779 GND.n4171 GND.n1692 585
R7780 GND.n4572 GND.n1692 585
R7781 GND.n4170 GND.n4169 585
R7782 GND.n4169 GND.n4168 585
R7783 GND.n1920 GND.n1681 585
R7784 GND.n4578 GND.n1681 585
R7785 GND.n4159 GND.n4158 585
R7786 GND.n4160 GND.n4159 585
R7787 GND.n1663 GND.n1662 585
R7788 GND.n4584 GND.n1663 585
R7789 GND.n4589 GND.n4588 585
R7790 GND.n4588 GND.n4587 585
R7791 GND.n5131 GND.n1077 585
R7792 GND.n1077 GND.n1076 585
R7793 GND.n6072 GND.n6071 585
R7794 GND.n6071 GND.n6070 585
R7795 GND.n6075 GND.n469 585
R7796 GND.n469 GND.n468 585
R7797 GND.n6077 GND.n6076 585
R7798 GND.n6078 GND.n6077 585
R7799 GND.n467 GND.n466 585
R7800 GND.n6079 GND.n467 585
R7801 GND.n6082 GND.n6081 585
R7802 GND.n6081 GND.n6080 585
R7803 GND.n6083 GND.n461 585
R7804 GND.n461 GND.n460 585
R7805 GND.n6085 GND.n6084 585
R7806 GND.n6086 GND.n6085 585
R7807 GND.n459 GND.n458 585
R7808 GND.n6087 GND.n459 585
R7809 GND.n6090 GND.n6089 585
R7810 GND.n6089 GND.n6088 585
R7811 GND.n6091 GND.n453 585
R7812 GND.n453 GND.n452 585
R7813 GND.n6093 GND.n6092 585
R7814 GND.n6094 GND.n6093 585
R7815 GND.n451 GND.n450 585
R7816 GND.n6095 GND.n451 585
R7817 GND.n6098 GND.n6097 585
R7818 GND.n6097 GND.n6096 585
R7819 GND.n6099 GND.n445 585
R7820 GND.n445 GND.n444 585
R7821 GND.n6101 GND.n6100 585
R7822 GND.n6102 GND.n6101 585
R7823 GND.n443 GND.n442 585
R7824 GND.n6103 GND.n443 585
R7825 GND.n6106 GND.n6105 585
R7826 GND.n6105 GND.n6104 585
R7827 GND.n6107 GND.n437 585
R7828 GND.n437 GND.n436 585
R7829 GND.n6109 GND.n6108 585
R7830 GND.n6110 GND.n6109 585
R7831 GND.n435 GND.n434 585
R7832 GND.n6111 GND.n435 585
R7833 GND.n6114 GND.n6113 585
R7834 GND.n6113 GND.n6112 585
R7835 GND.n6115 GND.n429 585
R7836 GND.n429 GND.n428 585
R7837 GND.n6117 GND.n6116 585
R7838 GND.n6118 GND.n6117 585
R7839 GND.n427 GND.n426 585
R7840 GND.n6119 GND.n427 585
R7841 GND.n6122 GND.n6121 585
R7842 GND.n6121 GND.n6120 585
R7843 GND.n6123 GND.n421 585
R7844 GND.n421 GND.n420 585
R7845 GND.n6125 GND.n6124 585
R7846 GND.n6126 GND.n6125 585
R7847 GND.n419 GND.n418 585
R7848 GND.n6127 GND.n419 585
R7849 GND.n6130 GND.n6129 585
R7850 GND.n6129 GND.n6128 585
R7851 GND.n6131 GND.n413 585
R7852 GND.n413 GND.n412 585
R7853 GND.n6133 GND.n6132 585
R7854 GND.n6134 GND.n6133 585
R7855 GND.n411 GND.n410 585
R7856 GND.n6135 GND.n411 585
R7857 GND.n6138 GND.n6137 585
R7858 GND.n6137 GND.n6136 585
R7859 GND.n6139 GND.n405 585
R7860 GND.n405 GND.n404 585
R7861 GND.n6141 GND.n6140 585
R7862 GND.n6142 GND.n6141 585
R7863 GND.n403 GND.n402 585
R7864 GND.n6143 GND.n403 585
R7865 GND.n6146 GND.n6145 585
R7866 GND.n6145 GND.n6144 585
R7867 GND.n6147 GND.n397 585
R7868 GND.n397 GND.n396 585
R7869 GND.n6149 GND.n6148 585
R7870 GND.n6150 GND.n6149 585
R7871 GND.n395 GND.n394 585
R7872 GND.n6151 GND.n395 585
R7873 GND.n6154 GND.n6153 585
R7874 GND.n6153 GND.n6152 585
R7875 GND.n6155 GND.n389 585
R7876 GND.n389 GND.n387 585
R7877 GND.n6157 GND.n6156 585
R7878 GND.n6158 GND.n6157 585
R7879 GND.n390 GND.n388 585
R7880 GND.n388 GND.n289 585
R7881 GND.n4322 GND.n4321 585
R7882 GND.n4322 GND.n286 585
R7883 GND.n4323 GND.n4317 585
R7884 GND.n4323 GND.n279 585
R7885 GND.n4325 GND.n4324 585
R7886 GND.n4324 GND.n276 585
R7887 GND.n4326 GND.n4312 585
R7888 GND.n4312 GND.n268 585
R7889 GND.n4452 GND.n4327 585
R7890 GND.n4452 GND.n4451 585
R7891 GND.n4453 GND.n4311 585
R7892 GND.n4453 GND.n259 585
R7893 GND.n4455 GND.n4454 585
R7894 GND.n4454 GND.n256 585
R7895 GND.n4456 GND.n4306 585
R7896 GND.n4306 GND.n248 585
R7897 GND.n4458 GND.n4457 585
R7898 GND.n4458 GND.n245 585
R7899 GND.n4459 GND.n4305 585
R7900 GND.n4459 GND.n238 585
R7901 GND.n4461 GND.n4460 585
R7902 GND.n4460 GND.n235 585
R7903 GND.n4462 GND.n4300 585
R7904 GND.n4300 GND.n227 585
R7905 GND.n4464 GND.n4463 585
R7906 GND.n4464 GND.n224 585
R7907 GND.n4465 GND.n4299 585
R7908 GND.n4465 GND.n217 585
R7909 GND.n4467 GND.n4466 585
R7910 GND.n4466 GND.n214 585
R7911 GND.n4468 GND.n4277 585
R7912 GND.n4277 GND.n206 585
R7913 GND.n4470 GND.n4469 585
R7914 GND.n4471 GND.n4470 585
R7915 GND.n4278 GND.n4276 585
R7916 GND.n4276 GND.n197 585
R7917 GND.n4293 GND.n4292 585
R7918 GND.n4292 GND.n194 585
R7919 GND.n4291 GND.n4280 585
R7920 GND.n4291 GND.n187 585
R7921 GND.n4290 GND.n4289 585
R7922 GND.n4290 GND.n184 585
R7923 GND.n4287 GND.n4281 585
R7924 GND.n4281 GND.n175 585
R7925 GND.n4285 GND.n4284 585
R7926 GND.n4284 GND.n172 585
R7927 GND.n4283 GND.n1889 585
R7928 GND.n1893 GND.n1889 585
R7929 GND.n4501 GND.n1888 585
R7930 GND.n4501 GND.n4500 585
R7931 GND.n4503 GND.n4502 585
R7932 GND.n4502 GND.n155 585
R7933 GND.n4505 GND.n1804 585
R7934 GND.n1804 GND.n1803 585
R7935 GND.n4507 GND.n4506 585
R7936 GND.n4508 GND.n4507 585
R7937 GND.n1886 GND.n1802 585
R7938 GND.n1802 GND.n1797 585
R7939 GND.n1885 GND.n1884 585
R7940 GND.n1884 GND.n1794 585
R7941 GND.n1883 GND.n1882 585
R7942 GND.n1883 GND.n1787 585
R7943 GND.n1881 GND.n1806 585
R7944 GND.n1806 GND.n1784 585
R7945 GND.n1875 GND.n1807 585
R7946 GND.n1875 GND.n1778 585
R7947 GND.n1877 GND.n1876 585
R7948 GND.n1876 GND.n1775 585
R7949 GND.n1874 GND.n1809 585
R7950 GND.n1874 GND.n1768 585
R7951 GND.n1873 GND.n1872 585
R7952 GND.n1873 GND.n1765 585
R7953 GND.n1811 GND.n1810 585
R7954 GND.n1810 GND.n1757 585
R7955 GND.n1868 GND.n1867 585
R7956 GND.n1867 GND.n1754 585
R7957 GND.n1866 GND.n1813 585
R7958 GND.n1866 GND.n1747 585
R7959 GND.n1865 GND.n1864 585
R7960 GND.n1865 GND.n1744 585
R7961 GND.n1815 GND.n1814 585
R7962 GND.n1814 GND.n1736 585
R7963 GND.n1860 GND.n1859 585
R7964 GND.n1859 GND.n1733 585
R7965 GND.n1858 GND.n1817 585
R7966 GND.n1858 GND.n1726 585
R7967 GND.n1857 GND.n1856 585
R7968 GND.n1857 GND.n1723 585
R7969 GND.n1819 GND.n1818 585
R7970 GND.n1818 GND.n1715 585
R7971 GND.n1852 GND.n1851 585
R7972 GND.n1851 GND.n1712 585
R7973 GND.n1850 GND.n1821 585
R7974 GND.n1850 GND.n1705 585
R7975 GND.n1849 GND.n1848 585
R7976 GND.n1849 GND.n1702 585
R7977 GND.n1823 GND.n1822 585
R7978 GND.n1822 GND.n1694 585
R7979 GND.n1844 GND.n1843 585
R7980 GND.n1843 GND.n1691 585
R7981 GND.n1842 GND.n1825 585
R7982 GND.n1842 GND.n1683 585
R7983 GND.n1841 GND.n1840 585
R7984 GND.n1841 GND.n1680 585
R7985 GND.n1827 GND.n1826 585
R7986 GND.n1826 GND.n1671 585
R7987 GND.n1836 GND.n1835 585
R7988 GND.n1835 GND.n1666 585
R7989 GND.n1834 GND.n1829 585
R7990 GND.n1834 GND.n1664 585
R7991 GND.n1833 GND.n1832 585
R7992 GND.n1833 GND.n1590 585
R7993 GND.n1564 GND.n1563 585
R7994 GND.n4689 GND.n1564 585
R7995 GND.n4692 GND.n4691 585
R7996 GND.n4691 GND.n4690 585
R7997 GND.n4693 GND.n1558 585
R7998 GND.n1558 GND.n1557 585
R7999 GND.n4695 GND.n4694 585
R8000 GND.n4696 GND.n4695 585
R8001 GND.n1559 GND.n1555 585
R8002 GND.n4697 GND.n1555 585
R8003 GND.n4144 GND.n2048 585
R8004 GND.n2048 GND.n1554 585
R8005 GND.n4146 GND.n4145 585
R8006 GND.n4147 GND.n4146 585
R8007 GND.n2049 GND.n2047 585
R8008 GND.n2047 GND.n2045 585
R8009 GND.n4138 GND.n4137 585
R8010 GND.n4137 GND.n4136 585
R8011 GND.n2052 GND.n2051 585
R8012 GND.n2053 GND.n2052 585
R8013 GND.n4125 GND.n4124 585
R8014 GND.n4126 GND.n4125 585
R8015 GND.n2063 GND.n2062 585
R8016 GND.n2062 GND.n2060 585
R8017 GND.n4120 GND.n4119 585
R8018 GND.n4119 GND.n4118 585
R8019 GND.n2066 GND.n2065 585
R8020 GND.n2076 GND.n2066 585
R8021 GND.n4109 GND.n4108 585
R8022 GND.n4110 GND.n4109 585
R8023 GND.n2079 GND.n2078 585
R8024 GND.n2500 GND.n2078 585
R8025 GND.n4104 GND.n4103 585
R8026 GND.n4103 GND.n4102 585
R8027 GND.n2082 GND.n2081 585
R8028 GND.n2685 GND.n2082 585
R8029 GND.n4094 GND.n4093 585
R8030 GND.t31 GND.n4094 585
R8031 GND.n2093 GND.n2092 585
R8032 GND.n2487 GND.n2092 585
R8033 GND.n4089 GND.n4088 585
R8034 GND.n4088 GND.n4087 585
R8035 GND.n2096 GND.n2095 585
R8036 GND.n2480 GND.n2096 585
R8037 GND.n4078 GND.n4077 585
R8038 GND.n4079 GND.n4078 585
R8039 GND.n2107 GND.n2106 585
R8040 GND.n2473 GND.n2106 585
R8041 GND.n4073 GND.n4072 585
R8042 GND.n4072 GND.n4071 585
R8043 GND.n2110 GND.n2109 585
R8044 GND.n2466 GND.n2110 585
R8045 GND.n4062 GND.n4061 585
R8046 GND.n4063 GND.n4062 585
R8047 GND.n2122 GND.n2121 585
R8048 GND.n2458 GND.n2121 585
R8049 GND.n4057 GND.n4056 585
R8050 GND.n4056 GND.n4055 585
R8051 GND.n2125 GND.n2124 585
R8052 GND.n2728 GND.n2125 585
R8053 GND.n4046 GND.n4045 585
R8054 GND.n4047 GND.n4046 585
R8055 GND.n2136 GND.n2135 585
R8056 GND.n2445 GND.n2135 585
R8057 GND.n4041 GND.n4040 585
R8058 GND.n4040 GND.n4039 585
R8059 GND.n2139 GND.n2138 585
R8060 GND.n2742 GND.n2139 585
R8061 GND.n4030 GND.n4029 585
R8062 GND.n4031 GND.n4030 585
R8063 GND.n2150 GND.n2149 585
R8064 GND.n2431 GND.n2149 585
R8065 GND.n4025 GND.n4024 585
R8066 GND.n4024 GND.n4023 585
R8067 GND.n2153 GND.n2152 585
R8068 GND.n2757 GND.n2153 585
R8069 GND.n4014 GND.n4013 585
R8070 GND.n4015 GND.n4014 585
R8071 GND.n2165 GND.n2164 585
R8072 GND.n2418 GND.n2164 585
R8073 GND.n4009 GND.n4008 585
R8074 GND.n4008 GND.n4007 585
R8075 GND.n2168 GND.n2167 585
R8076 GND.n2772 GND.n2168 585
R8077 GND.n3998 GND.n3997 585
R8078 GND.n3999 GND.n3998 585
R8079 GND.n2179 GND.n2178 585
R8080 GND.n2392 GND.n2178 585
R8081 GND.n3993 GND.n3992 585
R8082 GND.n3992 GND.n3991 585
R8083 GND.n2182 GND.n2181 585
R8084 GND.n2404 GND.n2182 585
R8085 GND.n3982 GND.n3981 585
R8086 GND.n3983 GND.n3982 585
R8087 GND.n2194 GND.n2193 585
R8088 GND.n2199 GND.n2193 585
R8089 GND.n3977 GND.n3976 585
R8090 GND.n3976 GND.n3975 585
R8091 GND.n2197 GND.n2196 585
R8092 GND.n2381 GND.n2197 585
R8093 GND.n3966 GND.n3965 585
R8094 GND.n3967 GND.n3966 585
R8095 GND.n2210 GND.n2209 585
R8096 GND.n2374 GND.n2209 585
R8097 GND.n3961 GND.n3960 585
R8098 GND.n3960 GND.n3959 585
R8099 GND.n2213 GND.n2212 585
R8100 GND.n2367 GND.n2213 585
R8101 GND.n3950 GND.n3949 585
R8102 GND.n3951 GND.n3950 585
R8103 GND.n2224 GND.n2223 585
R8104 GND.n2359 GND.n2223 585
R8105 GND.n3945 GND.n3944 585
R8106 GND.n3944 GND.n3943 585
R8107 GND.n2227 GND.n2226 585
R8108 GND.n2823 GND.n2227 585
R8109 GND.n3934 GND.n3933 585
R8110 GND.n3935 GND.n3934 585
R8111 GND.n2238 GND.n2237 585
R8112 GND.n2346 GND.n2237 585
R8113 GND.n3929 GND.n3928 585
R8114 GND.n3928 GND.n3927 585
R8115 GND.n2241 GND.n2240 585
R8116 GND.n2339 GND.n2241 585
R8117 GND.n3918 GND.n3917 585
R8118 GND.n3919 GND.n3918 585
R8119 GND.n2253 GND.n2252 585
R8120 GND.n2332 GND.n2252 585
R8121 GND.n3913 GND.n3912 585
R8122 GND.n3912 GND.n3911 585
R8123 GND.n2256 GND.n2255 585
R8124 GND.n2290 GND.n2256 585
R8125 GND.n3902 GND.n3901 585
R8126 GND.n3903 GND.n3902 585
R8127 GND.n2949 GND.n2948 585
R8128 GND.n2948 GND.n2264 585
R8129 GND.n3897 GND.n3896 585
R8130 GND.n3896 GND.n3895 585
R8131 GND.n2952 GND.n2951 585
R8132 GND.n2953 GND.n2952 585
R8133 GND.n3886 GND.n3885 585
R8134 GND.n3887 GND.n3886 585
R8135 GND.n2962 GND.n2961 585
R8136 GND.n2961 GND.n2959 585
R8137 GND.n3881 GND.n3880 585
R8138 GND.n3880 GND.n3879 585
R8139 GND.n2965 GND.n2964 585
R8140 GND.n2966 GND.n2965 585
R8141 GND.n3158 GND.n3156 585
R8142 GND.n3158 GND.n3157 585
R8143 GND.n3160 GND.n3159 585
R8144 GND.n3159 GND.n1460 585
R8145 GND.n3161 GND.n3150 585
R8146 GND.n3150 GND.n1447 585
R8147 GND.n3164 GND.n3162 585
R8148 GND.n3164 GND.n3163 585
R8149 GND.n3166 GND.n3149 585
R8150 GND.n3166 GND.n3165 585
R8151 GND.n3168 GND.n3167 585
R8152 GND.n3167 GND.n1292 585
R8153 GND.n3169 GND.n3144 585
R8154 GND.n3144 GND.n1290 585
R8155 GND.n3171 GND.n3170 585
R8156 GND.n3171 GND.n2971 585
R8157 GND.n3172 GND.n3143 585
R8158 GND.n3172 GND.n2973 585
R8159 GND.n3174 GND.n3173 585
R8160 GND.n3173 GND.n2982 585
R8161 GND.n3175 GND.n3138 585
R8162 GND.n3138 GND.n2980 585
R8163 GND.n3177 GND.n3176 585
R8164 GND.n3177 GND.n2984 585
R8165 GND.n3178 GND.n3137 585
R8166 GND.n3178 GND.n2992 585
R8167 GND.n3180 GND.n3179 585
R8168 GND.n3179 GND.n2991 585
R8169 GND.n3181 GND.n3132 585
R8170 GND.n3132 GND.n3004 585
R8171 GND.n3183 GND.n3182 585
R8172 GND.n3183 GND.n3002 585
R8173 GND.n3184 GND.n3131 585
R8174 GND.n3184 GND.n3006 585
R8175 GND.n3186 GND.n3185 585
R8176 GND.n3185 GND.n3015 585
R8177 GND.n3187 GND.n3126 585
R8178 GND.n3126 GND.n3014 585
R8179 GND.n3189 GND.n3188 585
R8180 GND.n3189 GND.n3028 585
R8181 GND.n3190 GND.n3125 585
R8182 GND.n3190 GND.n3025 585
R8183 GND.n3192 GND.n3191 585
R8184 GND.n3191 GND.n3031 585
R8185 GND.n3193 GND.n3120 585
R8186 GND.n3120 GND.n3039 585
R8187 GND.n3195 GND.n3194 585
R8188 GND.n3195 GND.n3038 585
R8189 GND.n3196 GND.n3119 585
R8190 GND.n3196 GND.n3050 585
R8191 GND.n3198 GND.n3197 585
R8192 GND.n3197 GND.n3048 585
R8193 GND.n3199 GND.n3114 585
R8194 GND.n3114 GND.n3053 585
R8195 GND.n3201 GND.n3200 585
R8196 GND.n3201 GND.n3062 585
R8197 GND.n3202 GND.n3113 585
R8198 GND.n3202 GND.n3060 585
R8199 GND.n3729 GND.n3728 585
R8200 GND.n3728 GND.n3727 585
R8201 GND.n3731 GND.n3109 585
R8202 GND.n3203 GND.n3109 585
R8203 GND.n3733 GND.n3732 585
R8204 GND.n3734 GND.n3733 585
R8205 GND.n3111 GND.n3108 585
R8206 GND.n3108 GND.n3103 585
R8207 GND.n3110 GND.n3090 585
R8208 GND.n3101 GND.n3090 585
R8209 GND.n3746 GND.n3745 585
R8210 GND.n3745 GND.n3744 585
R8211 GND.n3747 GND.n3087 585
R8212 GND.n3091 GND.n3087 585
R8213 GND.n3750 GND.n3749 585
R8214 GND.n3751 GND.n3750 585
R8215 GND.n3088 GND.n3086 585
R8216 GND.n3086 GND.n3080 585
R8217 GND.n3579 GND.n3577 585
R8218 GND.n3577 GND.n3078 585
R8219 GND.n3580 GND.n3573 585
R8220 GND.n3573 GND.n3217 585
R8221 GND.n3582 GND.n3581 585
R8222 GND.n3582 GND.n3214 585
R8223 GND.n3583 GND.n3572 585
R8224 GND.n3583 GND.n3226 585
R8225 GND.n3585 GND.n3584 585
R8226 GND.n3584 GND.n3224 585
R8227 GND.n3586 GND.n3567 585
R8228 GND.n3567 GND.n3228 585
R8229 GND.n3588 GND.n3587 585
R8230 GND.n3588 GND.n3236 585
R8231 GND.n3589 GND.n3566 585
R8232 GND.n3589 GND.n3235 585
R8233 GND.n3591 GND.n3590 585
R8234 GND.n3590 GND.n3248 585
R8235 GND.n3592 GND.n3561 585
R8236 GND.n3561 GND.n3246 585
R8237 GND.n3594 GND.n3593 585
R8238 GND.n3594 GND.n3250 585
R8239 GND.n3595 GND.n3560 585
R8240 GND.n3595 GND.n3259 585
R8241 GND.n3597 GND.n3596 585
R8242 GND.n3596 GND.n3258 585
R8243 GND.n3598 GND.n3555 585
R8244 GND.n3555 GND.n3272 585
R8245 GND.n3600 GND.n3599 585
R8246 GND.n3600 GND.n3269 585
R8247 GND.n3601 GND.n3554 585
R8248 GND.n3601 GND.n3275 585
R8249 GND.n3603 GND.n3602 585
R8250 GND.n3602 GND.n3283 585
R8251 GND.n3604 GND.n3538 585
R8252 GND.n3538 GND.n3282 585
R8253 GND.n3606 GND.n3605 585
R8254 GND.n3607 GND.n3606 585
R8255 GND.n3539 GND.n3537 585
R8256 GND.n3537 GND.n3290 585
R8257 GND.n3548 GND.n3547 585
R8258 GND.n3547 GND.n1177 585
R8259 GND.n3546 GND.n3541 585
R8260 GND.n3546 GND.n1174 585
R8261 GND.n3545 GND.n3544 585
R8262 GND.n3545 GND.n1165 585
R8263 GND.n1161 GND.n1160 585
R8264 GND.n5045 GND.n1161 585
R8265 GND.n5048 GND.n5047 585
R8266 GND.n5047 GND.n5046 585
R8267 GND.n5049 GND.n1155 585
R8268 GND.n1155 GND.n1154 585
R8269 GND.n5051 GND.n5050 585
R8270 GND.n5052 GND.n5051 585
R8271 GND.n1153 GND.n1152 585
R8272 GND.n5053 GND.n1153 585
R8273 GND.n5056 GND.n5055 585
R8274 GND.n5055 GND.n5054 585
R8275 GND.n5057 GND.n1147 585
R8276 GND.n1147 GND.n1146 585
R8277 GND.n5059 GND.n5058 585
R8278 GND.n5060 GND.n5059 585
R8279 GND.n1145 GND.n1144 585
R8280 GND.n5061 GND.n1145 585
R8281 GND.n5064 GND.n5063 585
R8282 GND.n5063 GND.n5062 585
R8283 GND.n5065 GND.n1139 585
R8284 GND.n1139 GND.n1138 585
R8285 GND.n5067 GND.n5066 585
R8286 GND.n5068 GND.n5067 585
R8287 GND.n1137 GND.n1136 585
R8288 GND.n5069 GND.n1137 585
R8289 GND.n5072 GND.n5071 585
R8290 GND.n5071 GND.n5070 585
R8291 GND.n5073 GND.n1131 585
R8292 GND.n1131 GND.n1130 585
R8293 GND.n5075 GND.n5074 585
R8294 GND.n5076 GND.n5075 585
R8295 GND.n1129 GND.n1128 585
R8296 GND.n5077 GND.n1129 585
R8297 GND.n5080 GND.n5079 585
R8298 GND.n5079 GND.n5078 585
R8299 GND.n5081 GND.n1123 585
R8300 GND.n1123 GND.n1122 585
R8301 GND.n5083 GND.n5082 585
R8302 GND.n5084 GND.n5083 585
R8303 GND.n1121 GND.n1120 585
R8304 GND.n5085 GND.n1121 585
R8305 GND.n5088 GND.n5087 585
R8306 GND.n5087 GND.n5086 585
R8307 GND.n5089 GND.n1115 585
R8308 GND.n1115 GND.n1114 585
R8309 GND.n5091 GND.n5090 585
R8310 GND.n5092 GND.n5091 585
R8311 GND.n1113 GND.n1112 585
R8312 GND.n5093 GND.n1113 585
R8313 GND.n5096 GND.n5095 585
R8314 GND.n5095 GND.n5094 585
R8315 GND.n5097 GND.n1107 585
R8316 GND.n1107 GND.n1106 585
R8317 GND.n5099 GND.n5098 585
R8318 GND.n5100 GND.n5099 585
R8319 GND.n1105 GND.n1104 585
R8320 GND.n5101 GND.n1105 585
R8321 GND.n5104 GND.n5103 585
R8322 GND.n5103 GND.n5102 585
R8323 GND.n5105 GND.n1099 585
R8324 GND.n1099 GND.n1098 585
R8325 GND.n5107 GND.n5106 585
R8326 GND.n5108 GND.n5107 585
R8327 GND.n1097 GND.n1096 585
R8328 GND.n5109 GND.n1097 585
R8329 GND.n5112 GND.n5111 585
R8330 GND.n5111 GND.n5110 585
R8331 GND.n5113 GND.n1091 585
R8332 GND.n1091 GND.n1090 585
R8333 GND.n5115 GND.n5114 585
R8334 GND.n5116 GND.n5115 585
R8335 GND.n1089 GND.n1088 585
R8336 GND.n5117 GND.n1089 585
R8337 GND.n5120 GND.n5119 585
R8338 GND.n5119 GND.n5118 585
R8339 GND.n5121 GND.n1084 585
R8340 GND.n1084 GND.n1083 585
R8341 GND.n5123 GND.n5122 585
R8342 GND.n5124 GND.n5123 585
R8343 GND.n1082 GND.n1081 585
R8344 GND.n5125 GND.n1082 585
R8345 GND.n5128 GND.n5127 585
R8346 GND.n5127 GND.n5126 585
R8347 GND.n4699 GND.n4698 585
R8348 GND.n4698 GND.n4697 585
R8349 GND.n4700 GND.n1552 585
R8350 GND.n1554 GND.n1552 585
R8351 GND.n2046 GND.n1550 585
R8352 GND.n4147 GND.n2046 585
R8353 GND.n4704 GND.n1549 585
R8354 GND.n2045 GND.n1549 585
R8355 GND.n4705 GND.n1548 585
R8356 GND.n4136 GND.n1548 585
R8357 GND.n4706 GND.n1547 585
R8358 GND.n2053 GND.n1547 585
R8359 GND.n2061 GND.n1545 585
R8360 GND.n4126 GND.n2061 585
R8361 GND.n4710 GND.n1544 585
R8362 GND.n2060 GND.n1544 585
R8363 GND.n4711 GND.n1543 585
R8364 GND.n4118 GND.n1543 585
R8365 GND.n4712 GND.n1542 585
R8366 GND.n2076 GND.n1542 585
R8367 GND.n2075 GND.n1540 585
R8368 GND.n4110 GND.n2075 585
R8369 GND.n4716 GND.n1539 585
R8370 GND.n2500 GND.n1539 585
R8371 GND.n4717 GND.n1538 585
R8372 GND.n4102 GND.n1538 585
R8373 GND.n4718 GND.n1537 585
R8374 GND.n2685 GND.n1537 585
R8375 GND.n2091 GND.n1535 585
R8376 GND.t31 GND.n2091 585
R8377 GND.n4722 GND.n1534 585
R8378 GND.n2487 GND.n1534 585
R8379 GND.n4723 GND.n1533 585
R8380 GND.n4087 GND.n1533 585
R8381 GND.n4724 GND.n1532 585
R8382 GND.n2480 GND.n1532 585
R8383 GND.n2104 GND.n1530 585
R8384 GND.n4079 GND.n2104 585
R8385 GND.n4728 GND.n1529 585
R8386 GND.n2473 GND.n1529 585
R8387 GND.n4729 GND.n1528 585
R8388 GND.n4071 GND.n1528 585
R8389 GND.n4730 GND.n1527 585
R8390 GND.n2466 GND.n1527 585
R8391 GND.n2119 GND.n1525 585
R8392 GND.n4063 GND.n2119 585
R8393 GND.n4734 GND.n1524 585
R8394 GND.n2458 GND.n1524 585
R8395 GND.n4735 GND.n1523 585
R8396 GND.n4055 GND.n1523 585
R8397 GND.n4736 GND.n1522 585
R8398 GND.n2728 GND.n1522 585
R8399 GND.n2134 GND.n1520 585
R8400 GND.n4047 GND.n2134 585
R8401 GND.n4740 GND.n1519 585
R8402 GND.n2445 GND.n1519 585
R8403 GND.n4741 GND.n1518 585
R8404 GND.n4039 GND.n1518 585
R8405 GND.n4742 GND.n1517 585
R8406 GND.n2742 GND.n1517 585
R8407 GND.n2147 GND.n1515 585
R8408 GND.n4031 GND.n2147 585
R8409 GND.n4746 GND.n1514 585
R8410 GND.n2431 GND.n1514 585
R8411 GND.n4747 GND.n1513 585
R8412 GND.n4023 GND.n1513 585
R8413 GND.n4748 GND.n1512 585
R8414 GND.n2757 GND.n1512 585
R8415 GND.n2162 GND.n1510 585
R8416 GND.n4015 GND.n2162 585
R8417 GND.n4752 GND.n1509 585
R8418 GND.n2418 GND.n1509 585
R8419 GND.n4753 GND.n1508 585
R8420 GND.n4007 GND.n1508 585
R8421 GND.n4754 GND.n1507 585
R8422 GND.n2772 GND.n1507 585
R8423 GND.n2176 GND.n1505 585
R8424 GND.n3999 GND.n2176 585
R8425 GND.n4758 GND.n1504 585
R8426 GND.n2392 GND.n1504 585
R8427 GND.n4759 GND.n1503 585
R8428 GND.n3991 GND.n1503 585
R8429 GND.n4760 GND.n1502 585
R8430 GND.n2404 GND.n1502 585
R8431 GND.n2191 GND.n1500 585
R8432 GND.n3983 GND.n2191 585
R8433 GND.n4764 GND.n1499 585
R8434 GND.n2199 GND.n1499 585
R8435 GND.n4765 GND.n1498 585
R8436 GND.n3975 GND.n1498 585
R8437 GND.n4766 GND.n1497 585
R8438 GND.n2381 GND.n1497 585
R8439 GND.n2207 GND.n1495 585
R8440 GND.n3967 GND.n2207 585
R8441 GND.n4770 GND.n1494 585
R8442 GND.n2374 GND.n1494 585
R8443 GND.n4771 GND.n1493 585
R8444 GND.n3959 GND.n1493 585
R8445 GND.n4772 GND.n1492 585
R8446 GND.n2367 GND.n1492 585
R8447 GND.n2221 GND.n1490 585
R8448 GND.n3951 GND.n2221 585
R8449 GND.n4776 GND.n1489 585
R8450 GND.n2359 GND.n1489 585
R8451 GND.n4777 GND.n1488 585
R8452 GND.n3943 GND.n1488 585
R8453 GND.n4778 GND.n1487 585
R8454 GND.n2823 GND.n1487 585
R8455 GND.n2236 GND.n1485 585
R8456 GND.n3935 GND.n2236 585
R8457 GND.n4782 GND.n1484 585
R8458 GND.n2346 GND.n1484 585
R8459 GND.n4783 GND.n1483 585
R8460 GND.n3927 GND.n1483 585
R8461 GND.n4784 GND.n1482 585
R8462 GND.n2339 GND.n1482 585
R8463 GND.n2250 GND.n1480 585
R8464 GND.n3919 GND.n2250 585
R8465 GND.n4788 GND.n1479 585
R8466 GND.n2332 GND.n1479 585
R8467 GND.n4789 GND.n1478 585
R8468 GND.n3911 GND.n1478 585
R8469 GND.n4790 GND.n1477 585
R8470 GND.n2290 GND.n1477 585
R8471 GND.n2265 GND.n1475 585
R8472 GND.n3903 GND.n2265 585
R8473 GND.n4794 GND.n1474 585
R8474 GND.n2264 GND.n1474 585
R8475 GND.n4795 GND.n1473 585
R8476 GND.n3895 GND.n1473 585
R8477 GND.n4796 GND.n1472 585
R8478 GND.n2953 GND.n1472 585
R8479 GND.n2960 GND.n1470 585
R8480 GND.n3887 GND.n2960 585
R8481 GND.n4800 GND.n1469 585
R8482 GND.n2959 GND.n1469 585
R8483 GND.n4801 GND.n1468 585
R8484 GND.n3879 GND.n1468 585
R8485 GND.n4802 GND.n1465 585
R8486 GND.n2966 GND.n1465 585
R8487 GND.n2040 GND.n2039 585
R8488 GND.n2037 GND.n1924 585
R8489 GND.n2036 GND.n2035 585
R8490 GND.n2020 GND.n1926 585
R8491 GND.n2025 GND.n2021 585
R8492 GND.n2018 GND.n1934 585
R8493 GND.n2017 GND.n2016 585
R8494 GND.n2001 GND.n1936 585
R8495 GND.n2003 GND.n2002 585
R8496 GND.n1999 GND.n1941 585
R8497 GND.n1998 GND.n1997 585
R8498 GND.n1982 GND.n1943 585
R8499 GND.n1984 GND.n1983 585
R8500 GND.n1980 GND.n1949 585
R8501 GND.n1979 GND.n1978 585
R8502 GND.n1972 GND.n1951 585
R8503 GND.n1974 GND.n1973 585
R8504 GND.n1970 GND.n1953 585
R8505 GND.n1969 GND.n1968 585
R8506 GND.n1962 GND.n1955 585
R8507 GND.n1964 GND.n1963 585
R8508 GND.n1960 GND.n1959 585
R8509 GND.n1958 GND.n1553 585
R8510 GND.n1565 GND.n1553 585
R8511 GND.n4151 GND.n1556 585
R8512 GND.n4697 GND.n1556 585
R8513 GND.n4150 GND.n4149 585
R8514 GND.n4149 GND.n1554 585
R8515 GND.n4148 GND.n2043 585
R8516 GND.n4148 GND.n4147 585
R8517 GND.n2056 GND.n2044 585
R8518 GND.n2045 GND.n2044 585
R8519 GND.n4135 GND.n4134 585
R8520 GND.n4136 GND.n4135 585
R8521 GND.n2055 GND.n2054 585
R8522 GND.n2054 GND.n2053 585
R8523 GND.n4128 GND.n4127 585
R8524 GND.n4127 GND.n4126 585
R8525 GND.n2059 GND.n2058 585
R8526 GND.n2060 GND.n2059 585
R8527 GND.n4117 GND.n4116 585
R8528 GND.n4118 GND.n4117 585
R8529 GND.n2070 GND.n2069 585
R8530 GND.n2076 GND.n2069 585
R8531 GND.n4112 GND.n4111 585
R8532 GND.n4111 GND.n4110 585
R8533 GND.n2073 GND.n2072 585
R8534 GND.n2500 GND.n2073 585
R8535 GND.n4101 GND.n4100 585
R8536 GND.n4102 GND.n4101 585
R8537 GND.n2086 GND.n2085 585
R8538 GND.n2685 GND.n2085 585
R8539 GND.n4096 GND.n4095 585
R8540 GND.n4095 GND.t31 585
R8541 GND.n2089 GND.n2088 585
R8542 GND.n2487 GND.n2089 585
R8543 GND.n4086 GND.n4085 585
R8544 GND.n4087 GND.n4086 585
R8545 GND.n2099 GND.n2098 585
R8546 GND.n2480 GND.n2098 585
R8547 GND.n4081 GND.n4080 585
R8548 GND.n4080 GND.n4079 585
R8549 GND.n2102 GND.n2101 585
R8550 GND.n2473 GND.n2102 585
R8551 GND.n4070 GND.n4069 585
R8552 GND.n4071 GND.n4070 585
R8553 GND.n2114 GND.n2113 585
R8554 GND.n2466 GND.n2113 585
R8555 GND.n4065 GND.n4064 585
R8556 GND.n4064 GND.n4063 585
R8557 GND.n2117 GND.n2116 585
R8558 GND.n2458 GND.n2117 585
R8559 GND.n4054 GND.n4053 585
R8560 GND.n4055 GND.n4054 585
R8561 GND.n2129 GND.n2128 585
R8562 GND.n2728 GND.n2128 585
R8563 GND.n4049 GND.n4048 585
R8564 GND.n4048 GND.n4047 585
R8565 GND.n2132 GND.n2131 585
R8566 GND.n2445 GND.n2132 585
R8567 GND.n4038 GND.n4037 585
R8568 GND.n4039 GND.n4038 585
R8569 GND.n2143 GND.n2142 585
R8570 GND.n2742 GND.n2142 585
R8571 GND.n4033 GND.n4032 585
R8572 GND.n4032 GND.n4031 585
R8573 GND.n2146 GND.n2145 585
R8574 GND.n2431 GND.n2146 585
R8575 GND.n4022 GND.n4021 585
R8576 GND.n4023 GND.n4022 585
R8577 GND.n2157 GND.n2156 585
R8578 GND.n2757 GND.n2156 585
R8579 GND.n4017 GND.n4016 585
R8580 GND.n4016 GND.n4015 585
R8581 GND.n2160 GND.n2159 585
R8582 GND.n2418 GND.n2160 585
R8583 GND.n4006 GND.n4005 585
R8584 GND.n4007 GND.n4006 585
R8585 GND.n2172 GND.n2171 585
R8586 GND.n2772 GND.n2171 585
R8587 GND.n4001 GND.n4000 585
R8588 GND.n4000 GND.n3999 585
R8589 GND.n2175 GND.n2174 585
R8590 GND.n2392 GND.n2175 585
R8591 GND.n3990 GND.n3989 585
R8592 GND.n3991 GND.n3990 585
R8593 GND.n2186 GND.n2185 585
R8594 GND.n2404 GND.n2185 585
R8595 GND.n3985 GND.n3984 585
R8596 GND.n3984 GND.n3983 585
R8597 GND.n2189 GND.n2188 585
R8598 GND.n2199 GND.n2189 585
R8599 GND.n3974 GND.n3973 585
R8600 GND.n3975 GND.n3974 585
R8601 GND.n2202 GND.n2201 585
R8602 GND.n2381 GND.n2201 585
R8603 GND.n3969 GND.n3968 585
R8604 GND.n3968 GND.n3967 585
R8605 GND.n2205 GND.n2204 585
R8606 GND.n2374 GND.n2205 585
R8607 GND.n3958 GND.n3957 585
R8608 GND.n3959 GND.n3958 585
R8609 GND.n2216 GND.n2215 585
R8610 GND.n2367 GND.n2215 585
R8611 GND.n3953 GND.n3952 585
R8612 GND.n3952 GND.n3951 585
R8613 GND.n2219 GND.n2218 585
R8614 GND.n2359 GND.n2219 585
R8615 GND.n3942 GND.n3941 585
R8616 GND.n3943 GND.n3942 585
R8617 GND.n2231 GND.n2230 585
R8618 GND.n2823 GND.n2230 585
R8619 GND.n3937 GND.n3936 585
R8620 GND.n3936 GND.n3935 585
R8621 GND.n2234 GND.n2233 585
R8622 GND.n2346 GND.n2234 585
R8623 GND.n3926 GND.n3925 585
R8624 GND.n3927 GND.n3926 585
R8625 GND.n2245 GND.n2244 585
R8626 GND.n2339 GND.n2244 585
R8627 GND.n3921 GND.n3920 585
R8628 GND.n3920 GND.n3919 585
R8629 GND.n2248 GND.n2247 585
R8630 GND.n2332 GND.n2248 585
R8631 GND.n3910 GND.n3909 585
R8632 GND.n3911 GND.n3910 585
R8633 GND.n2260 GND.n2259 585
R8634 GND.n2290 GND.n2259 585
R8635 GND.n3905 GND.n3904 585
R8636 GND.n3904 GND.n3903 585
R8637 GND.n2263 GND.n2262 585
R8638 GND.n2264 GND.n2263 585
R8639 GND.n3894 GND.n3893 585
R8640 GND.n3895 GND.n3894 585
R8641 GND.n2955 GND.n2954 585
R8642 GND.n2954 GND.n2953 585
R8643 GND.n3889 GND.n3888 585
R8644 GND.n3888 GND.n3887 585
R8645 GND.n2958 GND.n2957 585
R8646 GND.n2959 GND.n2958 585
R8647 GND.n3878 GND.n3877 585
R8648 GND.n3879 GND.n3878 585
R8649 GND.n2967 GND.n1446 585
R8650 GND.n2966 GND.n1446 585
R8651 GND.n4839 GND.n1436 585
R8652 GND.n1461 GND.n1437 585
R8653 GND.n4830 GND.n1445 585
R8654 GND.n4829 GND.n4828 585
R8655 GND.n4824 GND.n4823 585
R8656 GND.n1466 GND.n1464 585
R8657 GND.n4819 GND.n1463 585
R8658 GND.n4826 GND.n1463 585
R8659 GND.n4818 GND.n4805 585
R8660 GND.n4817 GND.n4806 585
R8661 GND.n4808 GND.n4807 585
R8662 GND.n4813 GND.n4810 585
R8663 GND.n4812 GND.n4811 585
R8664 GND.n1450 GND.n1402 585
R8665 GND.n4867 GND.n1403 585
R8666 GND.n4866 GND.n1404 585
R8667 GND.n1453 GND.n1405 585
R8668 GND.n4859 GND.n1414 585
R8669 GND.n4858 GND.n1415 585
R8670 GND.n1455 GND.n1416 585
R8671 GND.n4851 GND.n1425 585
R8672 GND.n4850 GND.n1426 585
R8673 GND.n1458 GND.n1427 585
R8674 GND.n4843 GND.n1435 585
R8675 GND.n5240 GND.n967 547.755
R8676 GND.n2671 GND.n2670 473.281
R8677 GND.n2585 GND.n2584 473.281
R8678 GND.n2847 GND.n2289 473.281
R8679 GND.n2945 GND.n2293 473.281
R8680 GND.n6070 GND.n6069 460.19
R8681 GND.n5938 GND.n553 301.784
R8682 GND.n5939 GND.n5938 301.784
R8683 GND.n5940 GND.n5939 301.784
R8684 GND.n5940 GND.n547 301.784
R8685 GND.n5948 GND.n547 301.784
R8686 GND.n5949 GND.n5948 301.784
R8687 GND.n5950 GND.n5949 301.784
R8688 GND.n5950 GND.n541 301.784
R8689 GND.n5958 GND.n541 301.784
R8690 GND.n5959 GND.n5958 301.784
R8691 GND.n5960 GND.n5959 301.784
R8692 GND.n5960 GND.n535 301.784
R8693 GND.n5968 GND.n535 301.784
R8694 GND.n5969 GND.n5968 301.784
R8695 GND.n5970 GND.n5969 301.784
R8696 GND.n5970 GND.n529 301.784
R8697 GND.n5978 GND.n529 301.784
R8698 GND.n5979 GND.n5978 301.784
R8699 GND.n5980 GND.n5979 301.784
R8700 GND.n5980 GND.n523 301.784
R8701 GND.n5988 GND.n523 301.784
R8702 GND.n5989 GND.n5988 301.784
R8703 GND.n5990 GND.n5989 301.784
R8704 GND.n5990 GND.n517 301.784
R8705 GND.n5998 GND.n517 301.784
R8706 GND.n5999 GND.n5998 301.784
R8707 GND.n6000 GND.n5999 301.784
R8708 GND.n6000 GND.n511 301.784
R8709 GND.n6008 GND.n511 301.784
R8710 GND.n6009 GND.n6008 301.784
R8711 GND.n6010 GND.n6009 301.784
R8712 GND.n6010 GND.n505 301.784
R8713 GND.n6018 GND.n505 301.784
R8714 GND.n6019 GND.n6018 301.784
R8715 GND.n6020 GND.n6019 301.784
R8716 GND.n6020 GND.n499 301.784
R8717 GND.n6028 GND.n499 301.784
R8718 GND.n6029 GND.n6028 301.784
R8719 GND.n6030 GND.n6029 301.784
R8720 GND.n6030 GND.n493 301.784
R8721 GND.n6038 GND.n493 301.784
R8722 GND.n6039 GND.n6038 301.784
R8723 GND.n6040 GND.n6039 301.784
R8724 GND.n6040 GND.n487 301.784
R8725 GND.n6048 GND.n487 301.784
R8726 GND.n6049 GND.n6048 301.784
R8727 GND.n6050 GND.n6049 301.784
R8728 GND.n6050 GND.n481 301.784
R8729 GND.n6058 GND.n481 301.784
R8730 GND.n6059 GND.n6058 301.784
R8731 GND.n6060 GND.n6059 301.784
R8732 GND.n6060 GND.n475 301.784
R8733 GND.n6068 GND.n475 301.784
R8734 GND.n6069 GND.n6068 301.784
R8735 GND.n68 GND.n54 289.615
R8736 GND.n48 GND.n34 289.615
R8737 GND.n29 GND.n15 289.615
R8738 GND.n127 GND.n113 289.615
R8739 GND.n107 GND.n93 289.615
R8740 GND.n88 GND.n74 289.615
R8741 GND.n5248 GND.n967 280.613
R8742 GND.n5249 GND.n5248 280.613
R8743 GND.n5250 GND.n5249 280.613
R8744 GND.n5250 GND.n961 280.613
R8745 GND.n5258 GND.n961 280.613
R8746 GND.n5259 GND.n5258 280.613
R8747 GND.n5260 GND.n5259 280.613
R8748 GND.n5260 GND.n955 280.613
R8749 GND.n5268 GND.n955 280.613
R8750 GND.n5269 GND.n5268 280.613
R8751 GND.n5270 GND.n5269 280.613
R8752 GND.n5270 GND.n949 280.613
R8753 GND.n5278 GND.n949 280.613
R8754 GND.n5279 GND.n5278 280.613
R8755 GND.n5280 GND.n5279 280.613
R8756 GND.n5280 GND.n943 280.613
R8757 GND.n5288 GND.n943 280.613
R8758 GND.n5289 GND.n5288 280.613
R8759 GND.n5290 GND.n5289 280.613
R8760 GND.n5290 GND.n937 280.613
R8761 GND.n5298 GND.n937 280.613
R8762 GND.n5299 GND.n5298 280.613
R8763 GND.n5300 GND.n5299 280.613
R8764 GND.n5300 GND.n931 280.613
R8765 GND.n5308 GND.n931 280.613
R8766 GND.n5309 GND.n5308 280.613
R8767 GND.n5310 GND.n5309 280.613
R8768 GND.n5310 GND.n925 280.613
R8769 GND.n5318 GND.n925 280.613
R8770 GND.n5319 GND.n5318 280.613
R8771 GND.n5320 GND.n5319 280.613
R8772 GND.n5320 GND.n919 280.613
R8773 GND.n5328 GND.n919 280.613
R8774 GND.n5329 GND.n5328 280.613
R8775 GND.n5330 GND.n5329 280.613
R8776 GND.n5330 GND.n913 280.613
R8777 GND.n5338 GND.n913 280.613
R8778 GND.n5339 GND.n5338 280.613
R8779 GND.n5340 GND.n5339 280.613
R8780 GND.n5340 GND.n907 280.613
R8781 GND.n5348 GND.n907 280.613
R8782 GND.n5349 GND.n5348 280.613
R8783 GND.n5350 GND.n5349 280.613
R8784 GND.n5350 GND.n901 280.613
R8785 GND.n5358 GND.n901 280.613
R8786 GND.n5359 GND.n5358 280.613
R8787 GND.n5360 GND.n5359 280.613
R8788 GND.n5360 GND.n895 280.613
R8789 GND.n5368 GND.n895 280.613
R8790 GND.n5369 GND.n5368 280.613
R8791 GND.n5370 GND.n5369 280.613
R8792 GND.n5370 GND.n889 280.613
R8793 GND.n5378 GND.n889 280.613
R8794 GND.n5379 GND.n5378 280.613
R8795 GND.n5380 GND.n5379 280.613
R8796 GND.n5380 GND.n883 280.613
R8797 GND.n5388 GND.n883 280.613
R8798 GND.n5389 GND.n5388 280.613
R8799 GND.n5390 GND.n5389 280.613
R8800 GND.n5390 GND.n877 280.613
R8801 GND.n5398 GND.n877 280.613
R8802 GND.n5399 GND.n5398 280.613
R8803 GND.n5400 GND.n5399 280.613
R8804 GND.n5400 GND.n871 280.613
R8805 GND.n5408 GND.n871 280.613
R8806 GND.n5409 GND.n5408 280.613
R8807 GND.n5410 GND.n5409 280.613
R8808 GND.n5410 GND.n865 280.613
R8809 GND.n5418 GND.n865 280.613
R8810 GND.n5419 GND.n5418 280.613
R8811 GND.n5420 GND.n5419 280.613
R8812 GND.n5420 GND.n859 280.613
R8813 GND.n5428 GND.n859 280.613
R8814 GND.n5429 GND.n5428 280.613
R8815 GND.n5430 GND.n5429 280.613
R8816 GND.n5430 GND.n853 280.613
R8817 GND.n5438 GND.n853 280.613
R8818 GND.n5439 GND.n5438 280.613
R8819 GND.n5440 GND.n5439 280.613
R8820 GND.n5440 GND.n847 280.613
R8821 GND.n5448 GND.n847 280.613
R8822 GND.n5449 GND.n5448 280.613
R8823 GND.n5450 GND.n5449 280.613
R8824 GND.n5450 GND.n841 280.613
R8825 GND.n5458 GND.n841 280.613
R8826 GND.n5459 GND.n5458 280.613
R8827 GND.n5460 GND.n5459 280.613
R8828 GND.n5460 GND.n835 280.613
R8829 GND.n5468 GND.n835 280.613
R8830 GND.n5469 GND.n5468 280.613
R8831 GND.n5470 GND.n5469 280.613
R8832 GND.n5470 GND.n829 280.613
R8833 GND.n5478 GND.n829 280.613
R8834 GND.n5479 GND.n5478 280.613
R8835 GND.n5480 GND.n5479 280.613
R8836 GND.n5480 GND.n823 280.613
R8837 GND.n5488 GND.n823 280.613
R8838 GND.n5489 GND.n5488 280.613
R8839 GND.n5490 GND.n5489 280.613
R8840 GND.n5490 GND.n817 280.613
R8841 GND.n5498 GND.n817 280.613
R8842 GND.n5499 GND.n5498 280.613
R8843 GND.n5500 GND.n5499 280.613
R8844 GND.n5500 GND.n811 280.613
R8845 GND.n5508 GND.n811 280.613
R8846 GND.n5509 GND.n5508 280.613
R8847 GND.n5510 GND.n5509 280.613
R8848 GND.n5510 GND.n805 280.613
R8849 GND.n5518 GND.n805 280.613
R8850 GND.n5519 GND.n5518 280.613
R8851 GND.n5520 GND.n5519 280.613
R8852 GND.n5520 GND.n799 280.613
R8853 GND.n5528 GND.n799 280.613
R8854 GND.n5529 GND.n5528 280.613
R8855 GND.n5530 GND.n5529 280.613
R8856 GND.n5530 GND.n793 280.613
R8857 GND.n5538 GND.n793 280.613
R8858 GND.n5539 GND.n5538 280.613
R8859 GND.n5540 GND.n5539 280.613
R8860 GND.n5540 GND.n787 280.613
R8861 GND.n5548 GND.n787 280.613
R8862 GND.n5549 GND.n5548 280.613
R8863 GND.n5550 GND.n5549 280.613
R8864 GND.n5550 GND.n781 280.613
R8865 GND.n5558 GND.n781 280.613
R8866 GND.n5559 GND.n5558 280.613
R8867 GND.n5560 GND.n5559 280.613
R8868 GND.n5560 GND.n775 280.613
R8869 GND.n5568 GND.n775 280.613
R8870 GND.n5569 GND.n5568 280.613
R8871 GND.n5570 GND.n5569 280.613
R8872 GND.n5570 GND.n769 280.613
R8873 GND.n5578 GND.n769 280.613
R8874 GND.n5579 GND.n5578 280.613
R8875 GND.n5580 GND.n5579 280.613
R8876 GND.n5580 GND.n763 280.613
R8877 GND.n5588 GND.n763 280.613
R8878 GND.n5589 GND.n5588 280.613
R8879 GND.n5590 GND.n5589 280.613
R8880 GND.n5590 GND.n757 280.613
R8881 GND.n5598 GND.n757 280.613
R8882 GND.n5599 GND.n5598 280.613
R8883 GND.n5600 GND.n5599 280.613
R8884 GND.n5600 GND.n751 280.613
R8885 GND.n5608 GND.n751 280.613
R8886 GND.n5609 GND.n5608 280.613
R8887 GND.n5610 GND.n5609 280.613
R8888 GND.n5610 GND.n745 280.613
R8889 GND.n5618 GND.n745 280.613
R8890 GND.n5619 GND.n5618 280.613
R8891 GND.n5620 GND.n5619 280.613
R8892 GND.n5620 GND.n739 280.613
R8893 GND.n5628 GND.n739 280.613
R8894 GND.n5629 GND.n5628 280.613
R8895 GND.n5630 GND.n5629 280.613
R8896 GND.n5630 GND.n733 280.613
R8897 GND.n5638 GND.n733 280.613
R8898 GND.n5639 GND.n5638 280.613
R8899 GND.n5640 GND.n5639 280.613
R8900 GND.n5640 GND.n727 280.613
R8901 GND.n5648 GND.n727 280.613
R8902 GND.n5649 GND.n5648 280.613
R8903 GND.n5650 GND.n5649 280.613
R8904 GND.n5650 GND.n721 280.613
R8905 GND.n5658 GND.n721 280.613
R8906 GND.n5659 GND.n5658 280.613
R8907 GND.n5660 GND.n5659 280.613
R8908 GND.n5660 GND.n715 280.613
R8909 GND.n5668 GND.n715 280.613
R8910 GND.n5669 GND.n5668 280.613
R8911 GND.n5670 GND.n5669 280.613
R8912 GND.n5670 GND.n709 280.613
R8913 GND.n5678 GND.n709 280.613
R8914 GND.n5679 GND.n5678 280.613
R8915 GND.n5680 GND.n5679 280.613
R8916 GND.n5680 GND.n703 280.613
R8917 GND.n5688 GND.n703 280.613
R8918 GND.n5689 GND.n5688 280.613
R8919 GND.n5690 GND.n5689 280.613
R8920 GND.n5690 GND.n697 280.613
R8921 GND.n5698 GND.n697 280.613
R8922 GND.n5699 GND.n5698 280.613
R8923 GND.n5700 GND.n5699 280.613
R8924 GND.n5700 GND.n691 280.613
R8925 GND.n5708 GND.n691 280.613
R8926 GND.n5709 GND.n5708 280.613
R8927 GND.n5710 GND.n5709 280.613
R8928 GND.n5710 GND.n685 280.613
R8929 GND.n5718 GND.n685 280.613
R8930 GND.n5719 GND.n5718 280.613
R8931 GND.n5720 GND.n5719 280.613
R8932 GND.n5720 GND.n679 280.613
R8933 GND.n5728 GND.n679 280.613
R8934 GND.n5729 GND.n5728 280.613
R8935 GND.n5730 GND.n5729 280.613
R8936 GND.n5730 GND.n673 280.613
R8937 GND.n5738 GND.n673 280.613
R8938 GND.n5739 GND.n5738 280.613
R8939 GND.n5740 GND.n5739 280.613
R8940 GND.n5740 GND.n667 280.613
R8941 GND.n5748 GND.n667 280.613
R8942 GND.n5749 GND.n5748 280.613
R8943 GND.n5750 GND.n5749 280.613
R8944 GND.n5750 GND.n661 280.613
R8945 GND.n5758 GND.n661 280.613
R8946 GND.n5759 GND.n5758 280.613
R8947 GND.n5760 GND.n5759 280.613
R8948 GND.n5760 GND.n655 280.613
R8949 GND.n5768 GND.n655 280.613
R8950 GND.n5769 GND.n5768 280.613
R8951 GND.n5770 GND.n5769 280.613
R8952 GND.n5770 GND.n649 280.613
R8953 GND.n5778 GND.n649 280.613
R8954 GND.n5779 GND.n5778 280.613
R8955 GND.n5780 GND.n5779 280.613
R8956 GND.n5780 GND.n643 280.613
R8957 GND.n5788 GND.n643 280.613
R8958 GND.n5789 GND.n5788 280.613
R8959 GND.n5790 GND.n5789 280.613
R8960 GND.n5790 GND.n637 280.613
R8961 GND.n5798 GND.n637 280.613
R8962 GND.n5799 GND.n5798 280.613
R8963 GND.n5800 GND.n5799 280.613
R8964 GND.n5800 GND.n631 280.613
R8965 GND.n5808 GND.n631 280.613
R8966 GND.n5809 GND.n5808 280.613
R8967 GND.n5810 GND.n5809 280.613
R8968 GND.n5810 GND.n625 280.613
R8969 GND.n5818 GND.n625 280.613
R8970 GND.n5819 GND.n5818 280.613
R8971 GND.n5820 GND.n5819 280.613
R8972 GND.n5820 GND.n619 280.613
R8973 GND.n5828 GND.n619 280.613
R8974 GND.n5829 GND.n5828 280.613
R8975 GND.n5830 GND.n5829 280.613
R8976 GND.n5830 GND.n613 280.613
R8977 GND.n5838 GND.n613 280.613
R8978 GND.n5839 GND.n5838 280.613
R8979 GND.n5840 GND.n5839 280.613
R8980 GND.n5840 GND.n607 280.613
R8981 GND.n5848 GND.n607 280.613
R8982 GND.n5849 GND.n5848 280.613
R8983 GND.n5850 GND.n5849 280.613
R8984 GND.n5850 GND.n601 280.613
R8985 GND.n5858 GND.n601 280.613
R8986 GND.n5859 GND.n5858 280.613
R8987 GND.n5860 GND.n5859 280.613
R8988 GND.n5860 GND.n595 280.613
R8989 GND.n5868 GND.n595 280.613
R8990 GND.n5869 GND.n5868 280.613
R8991 GND.n5870 GND.n5869 280.613
R8992 GND.n5870 GND.n589 280.613
R8993 GND.n5878 GND.n589 280.613
R8994 GND.n5879 GND.n5878 280.613
R8995 GND.n5880 GND.n5879 280.613
R8996 GND.n5880 GND.n583 280.613
R8997 GND.n5888 GND.n583 280.613
R8998 GND.n5889 GND.n5888 280.613
R8999 GND.n5890 GND.n5889 280.613
R9000 GND.n5890 GND.n577 280.613
R9001 GND.n5898 GND.n577 280.613
R9002 GND.n5899 GND.n5898 280.613
R9003 GND.n5900 GND.n5899 280.613
R9004 GND.n5900 GND.n571 280.613
R9005 GND.n5908 GND.n571 280.613
R9006 GND.n5909 GND.n5908 280.613
R9007 GND.n5910 GND.n5909 280.613
R9008 GND.n5910 GND.n565 280.613
R9009 GND.n5918 GND.n565 280.613
R9010 GND.n5919 GND.n5918 280.613
R9011 GND.n5920 GND.n5919 280.613
R9012 GND.n5920 GND.n559 280.613
R9013 GND.n5928 GND.n559 280.613
R9014 GND.n5929 GND.n5928 280.613
R9015 GND.n5930 GND.n5929 280.613
R9016 GND.n2302 GND.t132 260.649
R9017 GND.n2528 GND.t59 260.649
R9018 GND.n2947 GND.n2946 256.663
R9019 GND.n2947 GND.n2266 256.663
R9020 GND.n2947 GND.n2267 256.663
R9021 GND.n2947 GND.n2268 256.663
R9022 GND.n2947 GND.n2269 256.663
R9023 GND.n2947 GND.n2270 256.663
R9024 GND.n2947 GND.n2271 256.663
R9025 GND.n2947 GND.n2272 256.663
R9026 GND.n2947 GND.n2273 256.663
R9027 GND.n2947 GND.n2274 256.663
R9028 GND.n2947 GND.n2275 256.663
R9029 GND.n2947 GND.n2276 256.663
R9030 GND.n2898 GND.n2897 256.663
R9031 GND.n2947 GND.n2277 256.663
R9032 GND.n2947 GND.n2278 256.663
R9033 GND.n2947 GND.n2279 256.663
R9034 GND.n2947 GND.n2280 256.663
R9035 GND.n2947 GND.n2281 256.663
R9036 GND.n2947 GND.n2282 256.663
R9037 GND.n2947 GND.n2283 256.663
R9038 GND.n2947 GND.n2284 256.663
R9039 GND.n2947 GND.n2285 256.663
R9040 GND.n2947 GND.n2286 256.663
R9041 GND.n2947 GND.n2287 256.663
R9042 GND.n2947 GND.n2288 256.663
R9043 GND.n2580 GND.n2068 256.663
R9044 GND.n2590 GND.n2068 256.663
R9045 GND.n2577 GND.n2068 256.663
R9046 GND.n2597 GND.n2068 256.663
R9047 GND.n2574 GND.n2068 256.663
R9048 GND.n2604 GND.n2068 256.663
R9049 GND.n2571 GND.n2068 256.663
R9050 GND.n2611 GND.n2068 256.663
R9051 GND.n2568 GND.n2068 256.663
R9052 GND.n2618 GND.n2068 256.663
R9053 GND.n2564 GND.n2068 256.663
R9054 GND.n2625 GND.n2068 256.663
R9055 GND.n2628 GND.n1625 256.663
R9056 GND.n2629 GND.n2068 256.663
R9057 GND.n2558 GND.n2068 256.663
R9058 GND.n2636 GND.n2068 256.663
R9059 GND.n2552 GND.n2068 256.663
R9060 GND.n2643 GND.n2068 256.663
R9061 GND.n2549 GND.n2068 256.663
R9062 GND.n2650 GND.n2068 256.663
R9063 GND.n2546 GND.n2068 256.663
R9064 GND.n2657 GND.n2068 256.663
R9065 GND.n2543 GND.n2068 256.663
R9066 GND.n2664 GND.n2068 256.663
R9067 GND.n2540 GND.n2068 256.663
R9068 GND.n2325 GND.t26 252.594
R9069 GND.n2327 GND.t37 252.594
R9070 GND.n2561 GND.t73 252.594
R9071 GND.n2554 GND.t142 252.594
R9072 GND.n3497 GND.n1162 242.672
R9073 GND.n3499 GND.n1162 242.672
R9074 GND.n3507 GND.n1162 242.672
R9075 GND.n3509 GND.n1162 242.672
R9076 GND.n3518 GND.n1162 242.672
R9077 GND.n3521 GND.n1162 242.672
R9078 GND.n4833 GND.n1346 242.672
R9079 GND.n1441 GND.n1346 242.672
R9080 GND.n1430 GND.n1346 242.672
R9081 GND.n1421 GND.n1346 242.672
R9082 GND.n1418 GND.n1346 242.672
R9083 GND.n1409 GND.n1346 242.672
R9084 GND.n4688 GND.n1596 242.672
R9085 GND.n4688 GND.n1595 242.672
R9086 GND.n4688 GND.n1594 242.672
R9087 GND.n4688 GND.n1593 242.672
R9088 GND.n4688 GND.n1592 242.672
R9089 GND.n4688 GND.n1591 242.672
R9090 GND.n4429 GND.n295 242.672
R9091 GND.n4394 GND.n295 242.672
R9092 GND.n4419 GND.n295 242.672
R9093 GND.n4398 GND.n295 242.672
R9094 GND.n4409 GND.n295 242.672
R9095 GND.n4402 GND.n295 242.672
R9096 GND.n3362 GND.n1162 242.672
R9097 GND.n3370 GND.n1162 242.672
R9098 GND.n3372 GND.n1162 242.672
R9099 GND.n3380 GND.n1162 242.672
R9100 GND.n3382 GND.n1162 242.672
R9101 GND.n3390 GND.n1162 242.672
R9102 GND.n3392 GND.n1162 242.672
R9103 GND.n3400 GND.n1162 242.672
R9104 GND.n3402 GND.n1162 242.672
R9105 GND.n3410 GND.n1162 242.672
R9106 GND.n3412 GND.n1162 242.672
R9107 GND.n3422 GND.n1162 242.672
R9108 GND.n3424 GND.n1162 242.672
R9109 GND.n3432 GND.n1162 242.672
R9110 GND.n3434 GND.n1162 242.672
R9111 GND.n3442 GND.n1162 242.672
R9112 GND.n3444 GND.n1162 242.672
R9113 GND.n3455 GND.n1162 242.672
R9114 GND.n3457 GND.n1162 242.672
R9115 GND.n3465 GND.n1162 242.672
R9116 GND.n3467 GND.n1162 242.672
R9117 GND.n3475 GND.n1162 242.672
R9118 GND.n3477 GND.n1162 242.672
R9119 GND.n3485 GND.n1162 242.672
R9120 GND.n1398 GND.n1346 242.672
R9121 GND.n1394 GND.n1346 242.672
R9122 GND.n1389 GND.n1346 242.672
R9123 GND.n1386 GND.n1346 242.672
R9124 GND.n1381 GND.n1346 242.672
R9125 GND.n1378 GND.n1346 242.672
R9126 GND.n1373 GND.n1346 242.672
R9127 GND.n1368 GND.n1346 242.672
R9128 GND.n1363 GND.n1346 242.672
R9129 GND.n1360 GND.n1346 242.672
R9130 GND.n1355 GND.n1346 242.672
R9131 GND.n1352 GND.n1346 242.672
R9132 GND.n4911 GND.n1346 242.672
R9133 GND.n4914 GND.n1330 242.672
R9134 GND.n4915 GND.n1346 242.672
R9135 GND.n1346 GND.n1332 242.672
R9136 GND.n1346 GND.n1333 242.672
R9137 GND.n1346 GND.n1335 242.672
R9138 GND.n1346 GND.n1336 242.672
R9139 GND.n1346 GND.n1338 242.672
R9140 GND.n1346 GND.n1339 242.672
R9141 GND.n1346 GND.n1341 242.672
R9142 GND.n1346 GND.n1342 242.672
R9143 GND.n1346 GND.n1344 242.672
R9144 GND.n1346 GND.n1345 242.672
R9145 GND.n4688 GND.n4687 242.672
R9146 GND.n4688 GND.n1566 242.672
R9147 GND.n4688 GND.n1567 242.672
R9148 GND.n4688 GND.n1568 242.672
R9149 GND.n4688 GND.n1569 242.672
R9150 GND.n4688 GND.n1570 242.672
R9151 GND.n4688 GND.n1571 242.672
R9152 GND.n4688 GND.n1572 242.672
R9153 GND.n4688 GND.n1573 242.672
R9154 GND.n4688 GND.n1574 242.672
R9155 GND.n4688 GND.n1575 242.672
R9156 GND.n4645 GND.n1626 242.672
R9157 GND.n4688 GND.n1576 242.672
R9158 GND.n4688 GND.n1577 242.672
R9159 GND.n4688 GND.n1578 242.672
R9160 GND.n4688 GND.n1579 242.672
R9161 GND.n4688 GND.n1580 242.672
R9162 GND.n4688 GND.n1581 242.672
R9163 GND.n4688 GND.n1582 242.672
R9164 GND.n4688 GND.n1583 242.672
R9165 GND.n4688 GND.n1584 242.672
R9166 GND.n4688 GND.n1585 242.672
R9167 GND.n4688 GND.n1586 242.672
R9168 GND.n4688 GND.n1587 242.672
R9169 GND.n4688 GND.n1588 242.672
R9170 GND.n384 GND.n295 242.672
R9171 GND.n6169 GND.n295 242.672
R9172 GND.n375 GND.n295 242.672
R9173 GND.n6176 GND.n295 242.672
R9174 GND.n368 GND.n295 242.672
R9175 GND.n6183 GND.n295 242.672
R9176 GND.n361 GND.n295 242.672
R9177 GND.n6193 GND.n295 242.672
R9178 GND.n354 GND.n295 242.672
R9179 GND.n6200 GND.n295 242.672
R9180 GND.n347 GND.n295 242.672
R9181 GND.n6207 GND.n295 242.672
R9182 GND.n341 GND.n295 242.672
R9183 GND.n6216 GND.n295 242.672
R9184 GND.n333 GND.n295 242.672
R9185 GND.n6223 GND.n295 242.672
R9186 GND.n326 GND.n295 242.672
R9187 GND.n6230 GND.n295 242.672
R9188 GND.n319 GND.n295 242.672
R9189 GND.n6237 GND.n295 242.672
R9190 GND.n312 GND.n295 242.672
R9191 GND.n6244 GND.n295 242.672
R9192 GND.n303 GND.n295 242.672
R9193 GND.n6251 GND.n295 242.672
R9194 GND.n6254 GND.n295 242.672
R9195 GND.n2038 GND.n1565 242.672
R9196 GND.n1925 GND.n1565 242.672
R9197 GND.n2019 GND.n1565 242.672
R9198 GND.n1935 GND.n1565 242.672
R9199 GND.n2000 GND.n1565 242.672
R9200 GND.n1942 GND.n1565 242.672
R9201 GND.n1981 GND.n1565 242.672
R9202 GND.n1950 GND.n1565 242.672
R9203 GND.n1971 GND.n1565 242.672
R9204 GND.n1954 GND.n1565 242.672
R9205 GND.n1961 GND.n1565 242.672
R9206 GND.n4826 GND.n1462 242.672
R9207 GND.n4827 GND.n4826 242.672
R9208 GND.n4826 GND.n4825 242.672
R9209 GND.n4826 GND.n1448 242.672
R9210 GND.n4826 GND.n1449 242.672
R9211 GND.n4826 GND.n1451 242.672
R9212 GND.n4826 GND.n1452 242.672
R9213 GND.n4826 GND.n1454 242.672
R9214 GND.n4826 GND.n1456 242.672
R9215 GND.n4826 GND.n1457 242.672
R9216 GND.n4826 GND.n1459 242.672
R9217 GND.n6253 GND.n6252 240.244
R9218 GND.n6250 GND.n297 240.244
R9219 GND.n6246 GND.n6245 240.244
R9220 GND.n6243 GND.n304 240.244
R9221 GND.n6239 GND.n6238 240.244
R9222 GND.n6236 GND.n313 240.244
R9223 GND.n6232 GND.n6231 240.244
R9224 GND.n6229 GND.n320 240.244
R9225 GND.n6225 GND.n6224 240.244
R9226 GND.n6222 GND.n327 240.244
R9227 GND.n6218 GND.n6217 240.244
R9228 GND.n6215 GND.n334 240.244
R9229 GND.n6209 GND.n6208 240.244
R9230 GND.n6206 GND.n342 240.244
R9231 GND.n6202 GND.n6201 240.244
R9232 GND.n6199 GND.n348 240.244
R9233 GND.n6195 GND.n6194 240.244
R9234 GND.n6192 GND.n355 240.244
R9235 GND.n6185 GND.n6184 240.244
R9236 GND.n6182 GND.n362 240.244
R9237 GND.n6178 GND.n6177 240.244
R9238 GND.n6175 GND.n369 240.244
R9239 GND.n6171 GND.n6170 240.244
R9240 GND.n6168 GND.n376 240.244
R9241 GND.n4588 GND.n1663 240.244
R9242 GND.n4159 GND.n1663 240.244
R9243 GND.n4159 GND.n1681 240.244
R9244 GND.n4169 GND.n1681 240.244
R9245 GND.n4169 GND.n1692 240.244
R9246 GND.n4174 GND.n1692 240.244
R9247 GND.n4174 GND.n1703 240.244
R9248 GND.n4184 GND.n1703 240.244
R9249 GND.n4184 GND.n1713 240.244
R9250 GND.n4189 GND.n1713 240.244
R9251 GND.n4189 GND.n1724 240.244
R9252 GND.n4199 GND.n1724 240.244
R9253 GND.n4199 GND.n1734 240.244
R9254 GND.n4204 GND.n1734 240.244
R9255 GND.n4204 GND.n1745 240.244
R9256 GND.n4214 GND.n1745 240.244
R9257 GND.n4214 GND.n1755 240.244
R9258 GND.n4219 GND.n1755 240.244
R9259 GND.n4219 GND.n1766 240.244
R9260 GND.n4229 GND.n1766 240.244
R9261 GND.n4229 GND.n1776 240.244
R9262 GND.n4234 GND.n1776 240.244
R9263 GND.n4234 GND.n1785 240.244
R9264 GND.n4248 GND.n1785 240.244
R9265 GND.n4248 GND.n1795 240.244
R9266 GND.n1799 GND.n1795 240.244
R9267 GND.n1898 GND.n1799 240.244
R9268 GND.n1898 GND.n154 240.244
R9269 GND.n4259 GND.n154 240.244
R9270 GND.n4259 GND.n1891 240.244
R9271 GND.n4491 GND.n1891 240.244
R9272 GND.n4491 GND.n173 240.244
R9273 GND.n4483 GND.n173 240.244
R9274 GND.n4483 GND.n185 240.244
R9275 GND.n4479 GND.n185 240.244
R9276 GND.n4479 GND.n195 240.244
R9277 GND.n4275 GND.n195 240.244
R9278 GND.n4275 GND.n204 240.244
R9279 GND.n4352 GND.n204 240.244
R9280 GND.n4352 GND.n215 240.244
R9281 GND.n4356 GND.n215 240.244
R9282 GND.n4356 GND.n225 240.244
R9283 GND.n4366 GND.n225 240.244
R9284 GND.n4366 GND.n236 240.244
R9285 GND.n4370 GND.n236 240.244
R9286 GND.n4370 GND.n246 240.244
R9287 GND.n4381 GND.n246 240.244
R9288 GND.n4381 GND.n257 240.244
R9289 GND.n4328 GND.n257 240.244
R9290 GND.n4328 GND.n266 240.244
R9291 GND.n4443 GND.n266 240.244
R9292 GND.n4443 GND.n277 240.244
R9293 GND.n4439 GND.n277 240.244
R9294 GND.n4439 GND.n287 240.244
R9295 GND.n6160 GND.n287 240.244
R9296 GND.n1598 GND.n1597 240.244
R9297 GND.n4681 GND.n1597 240.244
R9298 GND.n4679 GND.n4678 240.244
R9299 GND.n4675 GND.n4674 240.244
R9300 GND.n4671 GND.n4670 240.244
R9301 GND.n4666 GND.n1610 240.244
R9302 GND.n4664 GND.n4663 240.244
R9303 GND.n4660 GND.n4659 240.244
R9304 GND.n4656 GND.n4655 240.244
R9305 GND.n4652 GND.n4651 240.244
R9306 GND.n4648 GND.n4647 240.244
R9307 GND.n4643 GND.n4642 240.244
R9308 GND.n4639 GND.n4638 240.244
R9309 GND.n4635 GND.n4634 240.244
R9310 GND.n4631 GND.n4630 240.244
R9311 GND.n4627 GND.n4626 240.244
R9312 GND.n4623 GND.n4622 240.244
R9313 GND.n4618 GND.n4617 240.244
R9314 GND.n4614 GND.n4613 240.244
R9315 GND.n4610 GND.n4609 240.244
R9316 GND.n4606 GND.n4605 240.244
R9317 GND.n4602 GND.n4601 240.244
R9318 GND.n4598 GND.n4597 240.244
R9319 GND.n1655 GND.n1589 240.244
R9320 GND.n4583 GND.n1599 240.244
R9321 GND.n4583 GND.n1672 240.244
R9322 GND.n4579 GND.n1672 240.244
R9323 GND.n4579 GND.n1679 240.244
R9324 GND.n4571 GND.n1679 240.244
R9325 GND.n4571 GND.n1695 240.244
R9326 GND.n4567 GND.n1695 240.244
R9327 GND.n4567 GND.n1701 240.244
R9328 GND.n4559 GND.n1701 240.244
R9329 GND.n4559 GND.n1716 240.244
R9330 GND.n4555 GND.n1716 240.244
R9331 GND.n4555 GND.n1722 240.244
R9332 GND.n4547 GND.n1722 240.244
R9333 GND.n4547 GND.n1737 240.244
R9334 GND.n4543 GND.n1737 240.244
R9335 GND.n4543 GND.n1743 240.244
R9336 GND.n4535 GND.n1743 240.244
R9337 GND.n4535 GND.n1758 240.244
R9338 GND.n4531 GND.n1758 240.244
R9339 GND.n4531 GND.n1764 240.244
R9340 GND.n4523 GND.n1764 240.244
R9341 GND.n4523 GND.n1779 240.244
R9342 GND.n4519 GND.n1779 240.244
R9343 GND.n4519 GND.n1783 240.244
R9344 GND.n4511 GND.n1783 240.244
R9345 GND.n4511 GND.n4510 240.244
R9346 GND.n4510 GND.n157 240.244
R9347 GND.n6334 GND.n157 240.244
R9348 GND.n6334 GND.n158 240.244
R9349 GND.n4498 GND.n158 240.244
R9350 GND.n4498 GND.n170 240.244
R9351 GND.n6329 GND.n170 240.244
R9352 GND.n6329 GND.n171 240.244
R9353 GND.n6321 GND.n171 240.244
R9354 GND.n6321 GND.n188 240.244
R9355 GND.n6317 GND.n188 240.244
R9356 GND.n6317 GND.n193 240.244
R9357 GND.n6309 GND.n193 240.244
R9358 GND.n6309 GND.n207 240.244
R9359 GND.n6305 GND.n207 240.244
R9360 GND.n6305 GND.n213 240.244
R9361 GND.n6297 GND.n213 240.244
R9362 GND.n6297 GND.n228 240.244
R9363 GND.n6293 GND.n228 240.244
R9364 GND.n6293 GND.n234 240.244
R9365 GND.n6285 GND.n234 240.244
R9366 GND.n6285 GND.n249 240.244
R9367 GND.n6281 GND.n249 240.244
R9368 GND.n6281 GND.n255 240.244
R9369 GND.n6273 GND.n255 240.244
R9370 GND.n6273 GND.n269 240.244
R9371 GND.n6269 GND.n269 240.244
R9372 GND.n6269 GND.n275 240.244
R9373 GND.n6261 GND.n275 240.244
R9374 GND.n6261 GND.n290 240.244
R9375 GND.n1300 GND.n1296 240.244
R9376 GND.n1343 GND.n1301 240.244
R9377 GND.n1305 GND.n1304 240.244
R9378 GND.n1340 GND.n1306 240.244
R9379 GND.n1310 GND.n1309 240.244
R9380 GND.n1315 GND.n1314 240.244
R9381 GND.n1337 GND.n1318 240.244
R9382 GND.n1320 GND.n1319 240.244
R9383 GND.n1334 GND.n1323 240.244
R9384 GND.n1325 GND.n1324 240.244
R9385 GND.n4916 GND.n1331 240.244
R9386 GND.n4913 GND.n4912 240.244
R9387 GND.n4910 GND.n1348 240.244
R9388 GND.n1354 GND.n1353 240.244
R9389 GND.n1359 GND.n1356 240.244
R9390 GND.n1362 GND.n1361 240.244
R9391 GND.n1367 GND.n1364 240.244
R9392 GND.n1372 GND.n1369 240.244
R9393 GND.n1377 GND.n1374 240.244
R9394 GND.n1380 GND.n1379 240.244
R9395 GND.n1385 GND.n1382 240.244
R9396 GND.n1388 GND.n1387 240.244
R9397 GND.n1393 GND.n1390 240.244
R9398 GND.n1399 GND.n1395 240.244
R9399 GND.n3527 GND.n1163 240.244
R9400 GND.n3527 GND.n1175 240.244
R9401 GND.n1185 GND.n1175 240.244
R9402 GND.n1186 GND.n1185 240.244
R9403 GND.n3608 GND.n1186 240.244
R9404 GND.n3608 GND.n1192 240.244
R9405 GND.n1193 GND.n1192 240.244
R9406 GND.n1194 GND.n1193 240.244
R9407 GND.n3270 GND.n1194 240.244
R9408 GND.n3270 GND.n1200 240.244
R9409 GND.n1201 GND.n1200 240.244
R9410 GND.n1202 GND.n1201 240.244
R9411 GND.n3251 GND.n1202 240.244
R9412 GND.n3251 GND.n1208 240.244
R9413 GND.n1209 GND.n1208 240.244
R9414 GND.n1210 GND.n1209 240.244
R9415 GND.n3239 GND.n1210 240.244
R9416 GND.n3239 GND.n1216 240.244
R9417 GND.n1217 GND.n1216 240.244
R9418 GND.n1218 GND.n1217 240.244
R9419 GND.n3215 GND.n1218 240.244
R9420 GND.n3215 GND.n1224 240.244
R9421 GND.n1225 GND.n1224 240.244
R9422 GND.n1226 GND.n1225 240.244
R9423 GND.n3084 GND.n1226 240.244
R9424 GND.n3084 GND.n1232 240.244
R9425 GND.n1233 GND.n1232 240.244
R9426 GND.n1234 GND.n1233 240.244
R9427 GND.n3105 GND.n1234 240.244
R9428 GND.n3105 GND.n1240 240.244
R9429 GND.n1241 GND.n1240 240.244
R9430 GND.n1242 GND.n1241 240.244
R9431 GND.n3061 GND.n1242 240.244
R9432 GND.n3061 GND.n1248 240.244
R9433 GND.n1249 GND.n1248 240.244
R9434 GND.n1250 GND.n1249 240.244
R9435 GND.n3777 GND.n1250 240.244
R9436 GND.n3777 GND.n1256 240.244
R9437 GND.n1257 GND.n1256 240.244
R9438 GND.n1258 GND.n1257 240.244
R9439 GND.n3026 GND.n1258 240.244
R9440 GND.n3026 GND.n1264 240.244
R9441 GND.n1265 GND.n1264 240.244
R9442 GND.n1266 GND.n1265 240.244
R9443 GND.n3007 GND.n1266 240.244
R9444 GND.n3007 GND.n1272 240.244
R9445 GND.n1273 GND.n1272 240.244
R9446 GND.n1274 GND.n1273 240.244
R9447 GND.n2995 GND.n1274 240.244
R9448 GND.n2995 GND.n1280 240.244
R9449 GND.n1281 GND.n1280 240.244
R9450 GND.n1282 GND.n1281 240.244
R9451 GND.n2974 GND.n1282 240.244
R9452 GND.n2974 GND.n1288 240.244
R9453 GND.n4954 GND.n1288 240.244
R9454 GND.n3363 GND.n3358 240.244
R9455 GND.n3369 GND.n3358 240.244
R9456 GND.n3373 GND.n3371 240.244
R9457 GND.n3379 GND.n3354 240.244
R9458 GND.n3383 GND.n3381 240.244
R9459 GND.n3389 GND.n3348 240.244
R9460 GND.n3393 GND.n3391 240.244
R9461 GND.n3399 GND.n3344 240.244
R9462 GND.n3403 GND.n3401 240.244
R9463 GND.n3409 GND.n3340 240.244
R9464 GND.n3413 GND.n3411 240.244
R9465 GND.n3421 GND.n3336 240.244
R9466 GND.n3425 GND.n3423 240.244
R9467 GND.n3431 GND.n3332 240.244
R9468 GND.n3435 GND.n3433 240.244
R9469 GND.n3441 GND.n3328 240.244
R9470 GND.n3445 GND.n3443 240.244
R9471 GND.n3454 GND.n3324 240.244
R9472 GND.n3458 GND.n3456 240.244
R9473 GND.n3464 GND.n3320 240.244
R9474 GND.n3468 GND.n3466 240.244
R9475 GND.n3474 GND.n3316 240.244
R9476 GND.n3478 GND.n3476 240.244
R9477 GND.n3484 GND.n3312 240.244
R9478 GND.n3487 GND.n3486 240.244
R9479 GND.n5043 GND.n1168 240.244
R9480 GND.n5039 GND.n1168 240.244
R9481 GND.n5039 GND.n1173 240.244
R9482 GND.n3613 GND.n1173 240.244
R9483 GND.n3613 GND.n3285 240.244
R9484 GND.n3621 GND.n3285 240.244
R9485 GND.n3621 GND.n3287 240.244
R9486 GND.n3287 GND.n3268 240.244
R9487 GND.n3637 GND.n3268 240.244
R9488 GND.n3637 GND.n3262 240.244
R9489 GND.n3645 GND.n3262 240.244
R9490 GND.n3645 GND.n3264 240.244
R9491 GND.n3264 GND.n3245 240.244
R9492 GND.n3662 GND.n3245 240.244
R9493 GND.n3662 GND.n3238 240.244
R9494 GND.n3670 GND.n3238 240.244
R9495 GND.n3670 GND.n3241 240.244
R9496 GND.n3241 GND.n3223 240.244
R9497 GND.n3687 GND.n3223 240.244
R9498 GND.n3687 GND.n3219 240.244
R9499 GND.n3693 GND.n3219 240.244
R9500 GND.n3693 GND.n3076 240.244
R9501 GND.n3757 GND.n3076 240.244
R9502 GND.n3757 GND.n3077 240.244
R9503 GND.n3097 GND.n3077 240.244
R9504 GND.n3099 GND.n3097 240.244
R9505 GND.n3742 GND.n3099 240.244
R9506 GND.n3742 GND.n3739 240.244
R9507 GND.n3739 GND.n3100 240.244
R9508 GND.n3719 GND.n3100 240.244
R9509 GND.n3721 GND.n3719 240.244
R9510 GND.n3721 GND.n3064 240.244
R9511 GND.n3765 GND.n3064 240.244
R9512 GND.n3765 GND.n3066 240.244
R9513 GND.n3066 GND.n3047 240.244
R9514 GND.n3782 GND.n3047 240.244
R9515 GND.n3782 GND.n3041 240.244
R9516 GND.n3790 GND.n3041 240.244
R9517 GND.n3790 GND.n3043 240.244
R9518 GND.n3043 GND.n3024 240.244
R9519 GND.n3806 GND.n3024 240.244
R9520 GND.n3806 GND.n3018 240.244
R9521 GND.n3814 GND.n3018 240.244
R9522 GND.n3814 GND.n3020 240.244
R9523 GND.n3020 GND.n3001 240.244
R9524 GND.n3831 GND.n3001 240.244
R9525 GND.n3831 GND.n2994 240.244
R9526 GND.n3839 GND.n2994 240.244
R9527 GND.n3839 GND.n2997 240.244
R9528 GND.n2997 GND.n2979 240.244
R9529 GND.n3859 GND.n2979 240.244
R9530 GND.n3859 GND.n2975 240.244
R9531 GND.n3865 GND.n2975 240.244
R9532 GND.n3865 GND.n1295 240.244
R9533 GND.n4952 GND.n1295 240.244
R9534 GND.n4408 GND.n4407 240.244
R9535 GND.n4411 GND.n4410 240.244
R9536 GND.n4418 GND.n4417 240.244
R9537 GND.n4421 GND.n4420 240.244
R9538 GND.n4428 GND.n4427 240.244
R9539 GND.n1670 GND.n1665 240.244
R9540 GND.n4161 GND.n1670 240.244
R9541 GND.n4161 GND.n1682 240.244
R9542 GND.n4167 GND.n1682 240.244
R9543 GND.n4167 GND.n1693 240.244
R9544 GND.n4176 GND.n1693 240.244
R9545 GND.n4176 GND.n1704 240.244
R9546 GND.n4182 GND.n1704 240.244
R9547 GND.n4182 GND.n1714 240.244
R9548 GND.n4191 GND.n1714 240.244
R9549 GND.n4191 GND.n1725 240.244
R9550 GND.n4197 GND.n1725 240.244
R9551 GND.n4197 GND.n1735 240.244
R9552 GND.n4206 GND.n1735 240.244
R9553 GND.n4206 GND.n1746 240.244
R9554 GND.n4212 GND.n1746 240.244
R9555 GND.n4212 GND.n1756 240.244
R9556 GND.n4221 GND.n1756 240.244
R9557 GND.n4221 GND.n1767 240.244
R9558 GND.n4227 GND.n1767 240.244
R9559 GND.n4227 GND.n1777 240.244
R9560 GND.n4236 GND.n1777 240.244
R9561 GND.n4236 GND.n1786 240.244
R9562 GND.n4246 GND.n1786 240.244
R9563 GND.n4246 GND.n1796 240.244
R9564 GND.n1800 GND.n1796 240.244
R9565 GND.n1800 GND.n152 240.244
R9566 GND.n6336 GND.n152 240.244
R9567 GND.n6336 GND.n153 240.244
R9568 GND.n1892 GND.n153 240.244
R9569 GND.n4489 GND.n1892 240.244
R9570 GND.n4489 GND.n174 240.244
R9571 GND.n4485 GND.n174 240.244
R9572 GND.n4485 GND.n186 240.244
R9573 GND.n4477 GND.n186 240.244
R9574 GND.n4477 GND.n196 240.244
R9575 GND.n4473 GND.n196 240.244
R9576 GND.n4473 GND.n205 240.244
R9577 GND.n4350 GND.n205 240.244
R9578 GND.n4350 GND.n216 240.244
R9579 GND.n4358 GND.n216 240.244
R9580 GND.n4358 GND.n226 240.244
R9581 GND.n4364 GND.n226 240.244
R9582 GND.n4364 GND.n237 240.244
R9583 GND.n4372 GND.n237 240.244
R9584 GND.n4372 GND.n247 240.244
R9585 GND.n4379 GND.n247 240.244
R9586 GND.n4379 GND.n258 240.244
R9587 GND.n4449 GND.n258 240.244
R9588 GND.n4449 GND.n267 240.244
R9589 GND.n4445 GND.n267 240.244
R9590 GND.n4445 GND.n278 240.244
R9591 GND.n4437 GND.n278 240.244
R9592 GND.n4437 GND.n288 240.244
R9593 GND.n386 GND.n288 240.244
R9594 GND.n1990 GND.n1989 240.244
R9595 GND.n1993 GND.n1992 240.244
R9596 GND.n2009 GND.n2008 240.244
R9597 GND.n2012 GND.n2011 240.244
R9598 GND.n1932 GND.n1928 240.244
R9599 GND.n4586 GND.n4585 240.244
R9600 GND.n4585 GND.n1668 240.244
R9601 GND.n4577 GND.n1668 240.244
R9602 GND.n4577 GND.n1684 240.244
R9603 GND.n4573 GND.n1684 240.244
R9604 GND.n4573 GND.n1690 240.244
R9605 GND.n4565 GND.n1690 240.244
R9606 GND.n4565 GND.n1706 240.244
R9607 GND.n4561 GND.n1706 240.244
R9608 GND.n4561 GND.n1711 240.244
R9609 GND.n4553 GND.n1711 240.244
R9610 GND.n4553 GND.n1727 240.244
R9611 GND.n4549 GND.n1727 240.244
R9612 GND.n4549 GND.n1732 240.244
R9613 GND.n4541 GND.n1732 240.244
R9614 GND.n4541 GND.n1748 240.244
R9615 GND.n4537 GND.n1748 240.244
R9616 GND.n4537 GND.n1753 240.244
R9617 GND.n4529 GND.n1753 240.244
R9618 GND.n4529 GND.n1769 240.244
R9619 GND.n4525 GND.n1769 240.244
R9620 GND.n4525 GND.n1774 240.244
R9621 GND.n4517 GND.n1774 240.244
R9622 GND.n4517 GND.n1788 240.244
R9623 GND.n4513 GND.n1788 240.244
R9624 GND.n4513 GND.n1793 240.244
R9625 GND.n4254 GND.n1793 240.244
R9626 GND.n4254 GND.n156 240.244
R9627 GND.n1894 GND.n156 240.244
R9628 GND.n4496 GND.n1894 240.244
R9629 GND.n4496 GND.n176 240.244
R9630 GND.n6327 GND.n176 240.244
R9631 GND.n6327 GND.n177 240.244
R9632 GND.n6323 GND.n177 240.244
R9633 GND.n6323 GND.n183 240.244
R9634 GND.n6315 GND.n183 240.244
R9635 GND.n6315 GND.n198 240.244
R9636 GND.n6311 GND.n198 240.244
R9637 GND.n6311 GND.n203 240.244
R9638 GND.n6303 GND.n203 240.244
R9639 GND.n6303 GND.n218 240.244
R9640 GND.n6299 GND.n218 240.244
R9641 GND.n6299 GND.n223 240.244
R9642 GND.n6291 GND.n223 240.244
R9643 GND.n6291 GND.n239 240.244
R9644 GND.n6287 GND.n239 240.244
R9645 GND.n6287 GND.n244 240.244
R9646 GND.n6279 GND.n244 240.244
R9647 GND.n6279 GND.n260 240.244
R9648 GND.n6275 GND.n260 240.244
R9649 GND.n6275 GND.n265 240.244
R9650 GND.n6267 GND.n265 240.244
R9651 GND.n6267 GND.n280 240.244
R9652 GND.n6263 GND.n280 240.244
R9653 GND.n6263 GND.n285 240.244
R9654 GND.n1411 GND.n1410 240.244
R9655 GND.n1420 GND.n1419 240.244
R9656 GND.n1429 GND.n1422 240.244
R9657 GND.n1432 GND.n1431 240.244
R9658 GND.n1443 GND.n1442 240.244
R9659 GND.n3529 GND.n1164 240.244
R9660 GND.n3529 GND.n1176 240.244
R9661 GND.n3292 GND.n1176 240.244
R9662 GND.n3536 GND.n3292 240.244
R9663 GND.n3536 GND.n3281 240.244
R9664 GND.n3623 GND.n3281 240.244
R9665 GND.n3623 GND.n3276 240.244
R9666 GND.n3630 GND.n3276 240.244
R9667 GND.n3630 GND.n3271 240.244
R9668 GND.n3271 GND.n3257 240.244
R9669 GND.n3647 GND.n3257 240.244
R9670 GND.n3647 GND.n3252 240.244
R9671 GND.n3654 GND.n3252 240.244
R9672 GND.n3654 GND.n3247 240.244
R9673 GND.n3247 GND.n3234 240.244
R9674 GND.n3672 GND.n3234 240.244
R9675 GND.n3672 GND.n3229 240.244
R9676 GND.n3679 GND.n3229 240.244
R9677 GND.n3679 GND.n3225 240.244
R9678 GND.n3225 GND.n3212 240.244
R9679 GND.n3695 GND.n3212 240.244
R9680 GND.n3695 GND.n3213 240.244
R9681 GND.n3213 GND.n3079 240.244
R9682 GND.n3083 GND.n3079 240.244
R9683 GND.n3703 GND.n3083 240.244
R9684 GND.n3703 GND.n3702 240.244
R9685 GND.n3702 GND.n3093 240.244
R9686 GND.n3102 GND.n3093 240.244
R9687 GND.n3106 GND.n3102 240.244
R9688 GND.n3204 GND.n3106 240.244
R9689 GND.n3716 GND.n3204 240.244
R9690 GND.n3716 GND.n3059 240.244
R9691 GND.n3767 GND.n3059 240.244
R9692 GND.n3767 GND.n3054 240.244
R9693 GND.n3774 GND.n3054 240.244
R9694 GND.n3774 GND.n3049 240.244
R9695 GND.n3049 GND.n3037 240.244
R9696 GND.n3792 GND.n3037 240.244
R9697 GND.n3792 GND.n3032 240.244
R9698 GND.n3799 GND.n3032 240.244
R9699 GND.n3799 GND.n3027 240.244
R9700 GND.n3027 GND.n3013 240.244
R9701 GND.n3816 GND.n3013 240.244
R9702 GND.n3816 GND.n3008 240.244
R9703 GND.n3823 GND.n3008 240.244
R9704 GND.n3823 GND.n3003 240.244
R9705 GND.n3003 GND.n2990 240.244
R9706 GND.n3841 GND.n2990 240.244
R9707 GND.n3841 GND.n2985 240.244
R9708 GND.n3853 GND.n2985 240.244
R9709 GND.n3853 GND.n2981 240.244
R9710 GND.n3847 GND.n2981 240.244
R9711 GND.n3847 GND.n2970 240.244
R9712 GND.n3870 GND.n2970 240.244
R9713 GND.n3870 GND.n1291 240.244
R9714 GND.n3500 GND.n3498 240.244
R9715 GND.n3506 GND.n3304 240.244
R9716 GND.n3510 GND.n3508 240.244
R9717 GND.n3517 GND.n3300 240.244
R9718 GND.n3520 GND.n3519 240.244
R9719 GND.n1178 GND.n1166 240.244
R9720 GND.n5037 GND.n1178 240.244
R9721 GND.n5037 GND.n1179 240.244
R9722 GND.n3611 GND.n1179 240.244
R9723 GND.n3611 GND.n3610 240.244
R9724 GND.n3610 GND.n3284 240.244
R9725 GND.n3284 GND.n3274 240.244
R9726 GND.n3632 GND.n3274 240.244
R9727 GND.n3635 GND.n3632 240.244
R9728 GND.n3635 GND.n3634 240.244
R9729 GND.n3634 GND.n3261 240.244
R9730 GND.n3261 GND.n3249 240.244
R9731 GND.n3656 GND.n3249 240.244
R9732 GND.n3660 GND.n3656 240.244
R9733 GND.n3660 GND.n3659 240.244
R9734 GND.n3659 GND.n3237 240.244
R9735 GND.n3237 GND.n3227 240.244
R9736 GND.n3681 GND.n3227 240.244
R9737 GND.n3685 GND.n3681 240.244
R9738 GND.n3685 GND.n3683 240.244
R9739 GND.n3683 GND.n3218 240.244
R9740 GND.n3218 GND.n3081 240.244
R9741 GND.n3755 GND.n3081 240.244
R9742 GND.n3755 GND.n3753 240.244
R9743 GND.n3753 GND.n3082 240.244
R9744 GND.n3094 GND.n3082 240.244
R9745 GND.n3096 GND.n3094 240.244
R9746 GND.n3737 GND.n3096 240.244
R9747 GND.n3737 GND.n3736 240.244
R9748 GND.n3736 GND.n3104 240.244
R9749 GND.n3724 GND.n3104 240.244
R9750 GND.n3725 GND.n3724 240.244
R9751 GND.n3725 GND.n3063 240.244
R9752 GND.n3063 GND.n3051 240.244
R9753 GND.n3776 GND.n3051 240.244
R9754 GND.n3780 GND.n3776 240.244
R9755 GND.n3780 GND.n3779 240.244
R9756 GND.n3779 GND.n3040 240.244
R9757 GND.n3040 GND.n3030 240.244
R9758 GND.n3801 GND.n3030 240.244
R9759 GND.n3804 GND.n3801 240.244
R9760 GND.n3804 GND.n3803 240.244
R9761 GND.n3803 GND.n3017 240.244
R9762 GND.n3017 GND.n3005 240.244
R9763 GND.n3825 GND.n3005 240.244
R9764 GND.n3829 GND.n3825 240.244
R9765 GND.n3829 GND.n3828 240.244
R9766 GND.n3828 GND.n2993 240.244
R9767 GND.n2993 GND.n2983 240.244
R9768 GND.n3855 GND.n2983 240.244
R9769 GND.n3857 GND.n3855 240.244
R9770 GND.n3857 GND.n2972 240.244
R9771 GND.n3867 GND.n2972 240.244
R9772 GND.n3868 GND.n3867 240.244
R9773 GND.n3868 GND.n1294 240.244
R9774 GND.n5247 GND.n968 240.244
R9775 GND.n5247 GND.n966 240.244
R9776 GND.n5251 GND.n966 240.244
R9777 GND.n5251 GND.n962 240.244
R9778 GND.n5257 GND.n962 240.244
R9779 GND.n5257 GND.n960 240.244
R9780 GND.n5261 GND.n960 240.244
R9781 GND.n5261 GND.n956 240.244
R9782 GND.n5267 GND.n956 240.244
R9783 GND.n5267 GND.n954 240.244
R9784 GND.n5271 GND.n954 240.244
R9785 GND.n5271 GND.n950 240.244
R9786 GND.n5277 GND.n950 240.244
R9787 GND.n5277 GND.n948 240.244
R9788 GND.n5281 GND.n948 240.244
R9789 GND.n5281 GND.n944 240.244
R9790 GND.n5287 GND.n944 240.244
R9791 GND.n5287 GND.n942 240.244
R9792 GND.n5291 GND.n942 240.244
R9793 GND.n5291 GND.n938 240.244
R9794 GND.n5297 GND.n938 240.244
R9795 GND.n5297 GND.n936 240.244
R9796 GND.n5301 GND.n936 240.244
R9797 GND.n5301 GND.n932 240.244
R9798 GND.n5307 GND.n932 240.244
R9799 GND.n5307 GND.n930 240.244
R9800 GND.n5311 GND.n930 240.244
R9801 GND.n5311 GND.n926 240.244
R9802 GND.n5317 GND.n926 240.244
R9803 GND.n5317 GND.n924 240.244
R9804 GND.n5321 GND.n924 240.244
R9805 GND.n5321 GND.n920 240.244
R9806 GND.n5327 GND.n920 240.244
R9807 GND.n5327 GND.n918 240.244
R9808 GND.n5331 GND.n918 240.244
R9809 GND.n5331 GND.n914 240.244
R9810 GND.n5337 GND.n914 240.244
R9811 GND.n5337 GND.n912 240.244
R9812 GND.n5341 GND.n912 240.244
R9813 GND.n5341 GND.n908 240.244
R9814 GND.n5347 GND.n908 240.244
R9815 GND.n5347 GND.n906 240.244
R9816 GND.n5351 GND.n906 240.244
R9817 GND.n5351 GND.n902 240.244
R9818 GND.n5357 GND.n902 240.244
R9819 GND.n5357 GND.n900 240.244
R9820 GND.n5361 GND.n900 240.244
R9821 GND.n5361 GND.n896 240.244
R9822 GND.n5367 GND.n896 240.244
R9823 GND.n5367 GND.n894 240.244
R9824 GND.n5371 GND.n894 240.244
R9825 GND.n5371 GND.n890 240.244
R9826 GND.n5377 GND.n890 240.244
R9827 GND.n5377 GND.n888 240.244
R9828 GND.n5381 GND.n888 240.244
R9829 GND.n5381 GND.n884 240.244
R9830 GND.n5387 GND.n884 240.244
R9831 GND.n5387 GND.n882 240.244
R9832 GND.n5391 GND.n882 240.244
R9833 GND.n5391 GND.n878 240.244
R9834 GND.n5397 GND.n878 240.244
R9835 GND.n5397 GND.n876 240.244
R9836 GND.n5401 GND.n876 240.244
R9837 GND.n5401 GND.n872 240.244
R9838 GND.n5407 GND.n872 240.244
R9839 GND.n5407 GND.n870 240.244
R9840 GND.n5411 GND.n870 240.244
R9841 GND.n5411 GND.n866 240.244
R9842 GND.n5417 GND.n866 240.244
R9843 GND.n5417 GND.n864 240.244
R9844 GND.n5421 GND.n864 240.244
R9845 GND.n5421 GND.n860 240.244
R9846 GND.n5427 GND.n860 240.244
R9847 GND.n5427 GND.n858 240.244
R9848 GND.n5431 GND.n858 240.244
R9849 GND.n5431 GND.n854 240.244
R9850 GND.n5437 GND.n854 240.244
R9851 GND.n5437 GND.n852 240.244
R9852 GND.n5441 GND.n852 240.244
R9853 GND.n5441 GND.n848 240.244
R9854 GND.n5447 GND.n848 240.244
R9855 GND.n5447 GND.n846 240.244
R9856 GND.n5451 GND.n846 240.244
R9857 GND.n5451 GND.n842 240.244
R9858 GND.n5457 GND.n842 240.244
R9859 GND.n5457 GND.n840 240.244
R9860 GND.n5461 GND.n840 240.244
R9861 GND.n5461 GND.n836 240.244
R9862 GND.n5467 GND.n836 240.244
R9863 GND.n5467 GND.n834 240.244
R9864 GND.n5471 GND.n834 240.244
R9865 GND.n5471 GND.n830 240.244
R9866 GND.n5477 GND.n830 240.244
R9867 GND.n5477 GND.n828 240.244
R9868 GND.n5481 GND.n828 240.244
R9869 GND.n5481 GND.n824 240.244
R9870 GND.n5487 GND.n824 240.244
R9871 GND.n5487 GND.n822 240.244
R9872 GND.n5491 GND.n822 240.244
R9873 GND.n5491 GND.n818 240.244
R9874 GND.n5497 GND.n818 240.244
R9875 GND.n5497 GND.n816 240.244
R9876 GND.n5501 GND.n816 240.244
R9877 GND.n5501 GND.n812 240.244
R9878 GND.n5507 GND.n812 240.244
R9879 GND.n5507 GND.n810 240.244
R9880 GND.n5511 GND.n810 240.244
R9881 GND.n5511 GND.n806 240.244
R9882 GND.n5517 GND.n806 240.244
R9883 GND.n5517 GND.n804 240.244
R9884 GND.n5521 GND.n804 240.244
R9885 GND.n5521 GND.n800 240.244
R9886 GND.n5527 GND.n800 240.244
R9887 GND.n5527 GND.n798 240.244
R9888 GND.n5531 GND.n798 240.244
R9889 GND.n5531 GND.n794 240.244
R9890 GND.n5537 GND.n794 240.244
R9891 GND.n5537 GND.n792 240.244
R9892 GND.n5541 GND.n792 240.244
R9893 GND.n5541 GND.n788 240.244
R9894 GND.n5547 GND.n788 240.244
R9895 GND.n5547 GND.n786 240.244
R9896 GND.n5551 GND.n786 240.244
R9897 GND.n5551 GND.n782 240.244
R9898 GND.n5557 GND.n782 240.244
R9899 GND.n5557 GND.n780 240.244
R9900 GND.n5561 GND.n780 240.244
R9901 GND.n5561 GND.n776 240.244
R9902 GND.n5567 GND.n776 240.244
R9903 GND.n5567 GND.n774 240.244
R9904 GND.n5571 GND.n774 240.244
R9905 GND.n5571 GND.n770 240.244
R9906 GND.n5577 GND.n770 240.244
R9907 GND.n5577 GND.n768 240.244
R9908 GND.n5581 GND.n768 240.244
R9909 GND.n5581 GND.n764 240.244
R9910 GND.n5587 GND.n764 240.244
R9911 GND.n5587 GND.n762 240.244
R9912 GND.n5591 GND.n762 240.244
R9913 GND.n5591 GND.n758 240.244
R9914 GND.n5597 GND.n758 240.244
R9915 GND.n5597 GND.n756 240.244
R9916 GND.n5601 GND.n756 240.244
R9917 GND.n5601 GND.n752 240.244
R9918 GND.n5607 GND.n752 240.244
R9919 GND.n5607 GND.n750 240.244
R9920 GND.n5611 GND.n750 240.244
R9921 GND.n5611 GND.n746 240.244
R9922 GND.n5617 GND.n746 240.244
R9923 GND.n5617 GND.n744 240.244
R9924 GND.n5621 GND.n744 240.244
R9925 GND.n5621 GND.n740 240.244
R9926 GND.n5627 GND.n740 240.244
R9927 GND.n5627 GND.n738 240.244
R9928 GND.n5631 GND.n738 240.244
R9929 GND.n5631 GND.n734 240.244
R9930 GND.n5637 GND.n734 240.244
R9931 GND.n5637 GND.n732 240.244
R9932 GND.n5641 GND.n732 240.244
R9933 GND.n5641 GND.n728 240.244
R9934 GND.n5647 GND.n728 240.244
R9935 GND.n5647 GND.n726 240.244
R9936 GND.n5651 GND.n726 240.244
R9937 GND.n5651 GND.n722 240.244
R9938 GND.n5657 GND.n722 240.244
R9939 GND.n5657 GND.n720 240.244
R9940 GND.n5661 GND.n720 240.244
R9941 GND.n5661 GND.n716 240.244
R9942 GND.n5667 GND.n716 240.244
R9943 GND.n5667 GND.n714 240.244
R9944 GND.n5671 GND.n714 240.244
R9945 GND.n5671 GND.n710 240.244
R9946 GND.n5677 GND.n710 240.244
R9947 GND.n5677 GND.n708 240.244
R9948 GND.n5681 GND.n708 240.244
R9949 GND.n5681 GND.n704 240.244
R9950 GND.n5687 GND.n704 240.244
R9951 GND.n5687 GND.n702 240.244
R9952 GND.n5691 GND.n702 240.244
R9953 GND.n5691 GND.n698 240.244
R9954 GND.n5697 GND.n698 240.244
R9955 GND.n5697 GND.n696 240.244
R9956 GND.n5701 GND.n696 240.244
R9957 GND.n5701 GND.n692 240.244
R9958 GND.n5707 GND.n692 240.244
R9959 GND.n5707 GND.n690 240.244
R9960 GND.n5711 GND.n690 240.244
R9961 GND.n5711 GND.n686 240.244
R9962 GND.n5717 GND.n686 240.244
R9963 GND.n5717 GND.n684 240.244
R9964 GND.n5721 GND.n684 240.244
R9965 GND.n5721 GND.n680 240.244
R9966 GND.n5727 GND.n680 240.244
R9967 GND.n5727 GND.n678 240.244
R9968 GND.n5731 GND.n678 240.244
R9969 GND.n5731 GND.n674 240.244
R9970 GND.n5737 GND.n674 240.244
R9971 GND.n5737 GND.n672 240.244
R9972 GND.n5741 GND.n672 240.244
R9973 GND.n5741 GND.n668 240.244
R9974 GND.n5747 GND.n668 240.244
R9975 GND.n5747 GND.n666 240.244
R9976 GND.n5751 GND.n666 240.244
R9977 GND.n5751 GND.n662 240.244
R9978 GND.n5757 GND.n662 240.244
R9979 GND.n5757 GND.n660 240.244
R9980 GND.n5761 GND.n660 240.244
R9981 GND.n5761 GND.n656 240.244
R9982 GND.n5767 GND.n656 240.244
R9983 GND.n5767 GND.n654 240.244
R9984 GND.n5771 GND.n654 240.244
R9985 GND.n5771 GND.n650 240.244
R9986 GND.n5777 GND.n650 240.244
R9987 GND.n5777 GND.n648 240.244
R9988 GND.n5781 GND.n648 240.244
R9989 GND.n5781 GND.n644 240.244
R9990 GND.n5787 GND.n644 240.244
R9991 GND.n5787 GND.n642 240.244
R9992 GND.n5791 GND.n642 240.244
R9993 GND.n5791 GND.n638 240.244
R9994 GND.n5797 GND.n638 240.244
R9995 GND.n5797 GND.n636 240.244
R9996 GND.n5801 GND.n636 240.244
R9997 GND.n5801 GND.n632 240.244
R9998 GND.n5807 GND.n632 240.244
R9999 GND.n5807 GND.n630 240.244
R10000 GND.n5811 GND.n630 240.244
R10001 GND.n5811 GND.n626 240.244
R10002 GND.n5817 GND.n626 240.244
R10003 GND.n5817 GND.n624 240.244
R10004 GND.n5821 GND.n624 240.244
R10005 GND.n5821 GND.n620 240.244
R10006 GND.n5827 GND.n620 240.244
R10007 GND.n5827 GND.n618 240.244
R10008 GND.n5831 GND.n618 240.244
R10009 GND.n5831 GND.n614 240.244
R10010 GND.n5837 GND.n614 240.244
R10011 GND.n5837 GND.n612 240.244
R10012 GND.n5841 GND.n612 240.244
R10013 GND.n5841 GND.n608 240.244
R10014 GND.n5847 GND.n608 240.244
R10015 GND.n5847 GND.n606 240.244
R10016 GND.n5851 GND.n606 240.244
R10017 GND.n5851 GND.n602 240.244
R10018 GND.n5857 GND.n602 240.244
R10019 GND.n5857 GND.n600 240.244
R10020 GND.n5861 GND.n600 240.244
R10021 GND.n5861 GND.n596 240.244
R10022 GND.n5867 GND.n596 240.244
R10023 GND.n5867 GND.n594 240.244
R10024 GND.n5871 GND.n594 240.244
R10025 GND.n5871 GND.n590 240.244
R10026 GND.n5877 GND.n590 240.244
R10027 GND.n5877 GND.n588 240.244
R10028 GND.n5881 GND.n588 240.244
R10029 GND.n5881 GND.n584 240.244
R10030 GND.n5887 GND.n584 240.244
R10031 GND.n5887 GND.n582 240.244
R10032 GND.n5891 GND.n582 240.244
R10033 GND.n5891 GND.n578 240.244
R10034 GND.n5897 GND.n578 240.244
R10035 GND.n5897 GND.n576 240.244
R10036 GND.n5901 GND.n576 240.244
R10037 GND.n5901 GND.n572 240.244
R10038 GND.n5907 GND.n572 240.244
R10039 GND.n5907 GND.n570 240.244
R10040 GND.n5911 GND.n570 240.244
R10041 GND.n5911 GND.n566 240.244
R10042 GND.n5917 GND.n566 240.244
R10043 GND.n5917 GND.n564 240.244
R10044 GND.n5921 GND.n564 240.244
R10045 GND.n5921 GND.n560 240.244
R10046 GND.n5927 GND.n560 240.244
R10047 GND.n5927 GND.n558 240.244
R10048 GND.n5931 GND.n558 240.244
R10049 GND.n5937 GND.n554 240.244
R10050 GND.n5937 GND.n552 240.244
R10051 GND.n5941 GND.n552 240.244
R10052 GND.n5941 GND.n548 240.244
R10053 GND.n5947 GND.n548 240.244
R10054 GND.n5947 GND.n546 240.244
R10055 GND.n5951 GND.n546 240.244
R10056 GND.n5951 GND.n542 240.244
R10057 GND.n5957 GND.n542 240.244
R10058 GND.n5957 GND.n540 240.244
R10059 GND.n5961 GND.n540 240.244
R10060 GND.n5961 GND.n536 240.244
R10061 GND.n5967 GND.n536 240.244
R10062 GND.n5967 GND.n534 240.244
R10063 GND.n5971 GND.n534 240.244
R10064 GND.n5971 GND.n530 240.244
R10065 GND.n5977 GND.n530 240.244
R10066 GND.n5977 GND.n528 240.244
R10067 GND.n5981 GND.n528 240.244
R10068 GND.n5981 GND.n524 240.244
R10069 GND.n5987 GND.n524 240.244
R10070 GND.n5987 GND.n522 240.244
R10071 GND.n5991 GND.n522 240.244
R10072 GND.n5991 GND.n518 240.244
R10073 GND.n5997 GND.n518 240.244
R10074 GND.n5997 GND.n516 240.244
R10075 GND.n6001 GND.n516 240.244
R10076 GND.n6001 GND.n512 240.244
R10077 GND.n6007 GND.n512 240.244
R10078 GND.n6007 GND.n510 240.244
R10079 GND.n6011 GND.n510 240.244
R10080 GND.n6011 GND.n506 240.244
R10081 GND.n6017 GND.n506 240.244
R10082 GND.n6017 GND.n504 240.244
R10083 GND.n6021 GND.n504 240.244
R10084 GND.n6021 GND.n500 240.244
R10085 GND.n6027 GND.n500 240.244
R10086 GND.n6027 GND.n498 240.244
R10087 GND.n6031 GND.n498 240.244
R10088 GND.n6031 GND.n494 240.244
R10089 GND.n6037 GND.n494 240.244
R10090 GND.n6037 GND.n492 240.244
R10091 GND.n6041 GND.n492 240.244
R10092 GND.n6041 GND.n488 240.244
R10093 GND.n6047 GND.n488 240.244
R10094 GND.n6047 GND.n486 240.244
R10095 GND.n6051 GND.n486 240.244
R10096 GND.n6051 GND.n482 240.244
R10097 GND.n6057 GND.n482 240.244
R10098 GND.n6057 GND.n480 240.244
R10099 GND.n6061 GND.n480 240.244
R10100 GND.n6061 GND.n476 240.244
R10101 GND.n6067 GND.n476 240.244
R10102 GND.n6067 GND.n474 240.244
R10103 GND.n6071 GND.n474 240.244
R10104 GND.n5127 GND.n1082 240.244
R10105 GND.n5123 GND.n1082 240.244
R10106 GND.n5123 GND.n1084 240.244
R10107 GND.n5119 GND.n1084 240.244
R10108 GND.n5119 GND.n1089 240.244
R10109 GND.n5115 GND.n1089 240.244
R10110 GND.n5115 GND.n1091 240.244
R10111 GND.n5111 GND.n1091 240.244
R10112 GND.n5111 GND.n1097 240.244
R10113 GND.n5107 GND.n1097 240.244
R10114 GND.n5107 GND.n1099 240.244
R10115 GND.n5103 GND.n1099 240.244
R10116 GND.n5103 GND.n1105 240.244
R10117 GND.n5099 GND.n1105 240.244
R10118 GND.n5099 GND.n1107 240.244
R10119 GND.n5095 GND.n1107 240.244
R10120 GND.n5095 GND.n1113 240.244
R10121 GND.n5091 GND.n1113 240.244
R10122 GND.n5091 GND.n1115 240.244
R10123 GND.n5087 GND.n1115 240.244
R10124 GND.n5087 GND.n1121 240.244
R10125 GND.n5083 GND.n1121 240.244
R10126 GND.n5083 GND.n1123 240.244
R10127 GND.n5079 GND.n1123 240.244
R10128 GND.n5079 GND.n1129 240.244
R10129 GND.n5075 GND.n1129 240.244
R10130 GND.n5075 GND.n1131 240.244
R10131 GND.n5071 GND.n1131 240.244
R10132 GND.n5071 GND.n1137 240.244
R10133 GND.n5067 GND.n1137 240.244
R10134 GND.n5067 GND.n1139 240.244
R10135 GND.n5063 GND.n1139 240.244
R10136 GND.n5063 GND.n1145 240.244
R10137 GND.n5059 GND.n1145 240.244
R10138 GND.n5059 GND.n1147 240.244
R10139 GND.n5055 GND.n1147 240.244
R10140 GND.n5055 GND.n1153 240.244
R10141 GND.n5051 GND.n1153 240.244
R10142 GND.n5051 GND.n1155 240.244
R10143 GND.n5047 GND.n1155 240.244
R10144 GND.n5047 GND.n1161 240.244
R10145 GND.n3545 GND.n1161 240.244
R10146 GND.n3546 GND.n3545 240.244
R10147 GND.n3547 GND.n3546 240.244
R10148 GND.n3547 GND.n3537 240.244
R10149 GND.n3606 GND.n3537 240.244
R10150 GND.n3606 GND.n3538 240.244
R10151 GND.n3602 GND.n3538 240.244
R10152 GND.n3602 GND.n3601 240.244
R10153 GND.n3601 GND.n3600 240.244
R10154 GND.n3600 GND.n3555 240.244
R10155 GND.n3596 GND.n3555 240.244
R10156 GND.n3596 GND.n3595 240.244
R10157 GND.n3595 GND.n3594 240.244
R10158 GND.n3594 GND.n3561 240.244
R10159 GND.n3590 GND.n3561 240.244
R10160 GND.n3590 GND.n3589 240.244
R10161 GND.n3589 GND.n3588 240.244
R10162 GND.n3588 GND.n3567 240.244
R10163 GND.n3584 GND.n3567 240.244
R10164 GND.n3584 GND.n3583 240.244
R10165 GND.n3583 GND.n3582 240.244
R10166 GND.n3582 GND.n3573 240.244
R10167 GND.n3577 GND.n3573 240.244
R10168 GND.n3577 GND.n3086 240.244
R10169 GND.n3750 GND.n3086 240.244
R10170 GND.n3750 GND.n3087 240.244
R10171 GND.n3745 GND.n3087 240.244
R10172 GND.n3745 GND.n3090 240.244
R10173 GND.n3108 GND.n3090 240.244
R10174 GND.n3733 GND.n3108 240.244
R10175 GND.n3733 GND.n3109 240.244
R10176 GND.n3728 GND.n3109 240.244
R10177 GND.n3728 GND.n3202 240.244
R10178 GND.n3202 GND.n3201 240.244
R10179 GND.n3201 GND.n3114 240.244
R10180 GND.n3197 GND.n3114 240.244
R10181 GND.n3197 GND.n3196 240.244
R10182 GND.n3196 GND.n3195 240.244
R10183 GND.n3195 GND.n3120 240.244
R10184 GND.n3191 GND.n3120 240.244
R10185 GND.n3191 GND.n3190 240.244
R10186 GND.n3190 GND.n3189 240.244
R10187 GND.n3189 GND.n3126 240.244
R10188 GND.n3185 GND.n3126 240.244
R10189 GND.n3185 GND.n3184 240.244
R10190 GND.n3184 GND.n3183 240.244
R10191 GND.n3183 GND.n3132 240.244
R10192 GND.n3179 GND.n3132 240.244
R10193 GND.n3179 GND.n3178 240.244
R10194 GND.n3178 GND.n3177 240.244
R10195 GND.n3177 GND.n3138 240.244
R10196 GND.n3173 GND.n3138 240.244
R10197 GND.n3173 GND.n3172 240.244
R10198 GND.n3172 GND.n3171 240.244
R10199 GND.n3171 GND.n3144 240.244
R10200 GND.n3167 GND.n3144 240.244
R10201 GND.n3167 GND.n3166 240.244
R10202 GND.n3166 GND.n3164 240.244
R10203 GND.n3164 GND.n3150 240.244
R10204 GND.n3159 GND.n3150 240.244
R10205 GND.n3159 GND.n3158 240.244
R10206 GND.n3158 GND.n2965 240.244
R10207 GND.n3880 GND.n2965 240.244
R10208 GND.n3880 GND.n2961 240.244
R10209 GND.n3886 GND.n2961 240.244
R10210 GND.n3886 GND.n2952 240.244
R10211 GND.n3896 GND.n2952 240.244
R10212 GND.n3896 GND.n2948 240.244
R10213 GND.n3902 GND.n2948 240.244
R10214 GND.n3902 GND.n2256 240.244
R10215 GND.n3912 GND.n2256 240.244
R10216 GND.n3912 GND.n2252 240.244
R10217 GND.n3918 GND.n2252 240.244
R10218 GND.n3918 GND.n2241 240.244
R10219 GND.n3928 GND.n2241 240.244
R10220 GND.n3928 GND.n2237 240.244
R10221 GND.n3934 GND.n2237 240.244
R10222 GND.n3934 GND.n2227 240.244
R10223 GND.n3944 GND.n2227 240.244
R10224 GND.n3944 GND.n2223 240.244
R10225 GND.n3950 GND.n2223 240.244
R10226 GND.n3950 GND.n2213 240.244
R10227 GND.n3960 GND.n2213 240.244
R10228 GND.n3960 GND.n2209 240.244
R10229 GND.n3966 GND.n2209 240.244
R10230 GND.n3966 GND.n2197 240.244
R10231 GND.n3976 GND.n2197 240.244
R10232 GND.n3976 GND.n2193 240.244
R10233 GND.n3982 GND.n2193 240.244
R10234 GND.n3982 GND.n2182 240.244
R10235 GND.n3992 GND.n2182 240.244
R10236 GND.n3992 GND.n2178 240.244
R10237 GND.n3998 GND.n2178 240.244
R10238 GND.n3998 GND.n2168 240.244
R10239 GND.n4008 GND.n2168 240.244
R10240 GND.n4008 GND.n2164 240.244
R10241 GND.n4014 GND.n2164 240.244
R10242 GND.n4014 GND.n2153 240.244
R10243 GND.n4024 GND.n2153 240.244
R10244 GND.n4024 GND.n2149 240.244
R10245 GND.n4030 GND.n2149 240.244
R10246 GND.n4030 GND.n2139 240.244
R10247 GND.n4040 GND.n2139 240.244
R10248 GND.n4040 GND.n2135 240.244
R10249 GND.n4046 GND.n2135 240.244
R10250 GND.n4046 GND.n2125 240.244
R10251 GND.n4056 GND.n2125 240.244
R10252 GND.n4056 GND.n2121 240.244
R10253 GND.n4062 GND.n2121 240.244
R10254 GND.n4062 GND.n2110 240.244
R10255 GND.n4072 GND.n2110 240.244
R10256 GND.n4072 GND.n2106 240.244
R10257 GND.n4078 GND.n2106 240.244
R10258 GND.n4078 GND.n2096 240.244
R10259 GND.n4088 GND.n2096 240.244
R10260 GND.n4088 GND.n2092 240.244
R10261 GND.n4094 GND.n2092 240.244
R10262 GND.n4094 GND.n2082 240.244
R10263 GND.n4103 GND.n2082 240.244
R10264 GND.n4103 GND.n2078 240.244
R10265 GND.n4109 GND.n2078 240.244
R10266 GND.n4109 GND.n2066 240.244
R10267 GND.n4119 GND.n2066 240.244
R10268 GND.n4119 GND.n2062 240.244
R10269 GND.n4125 GND.n2062 240.244
R10270 GND.n4125 GND.n2052 240.244
R10271 GND.n4137 GND.n2052 240.244
R10272 GND.n4137 GND.n2047 240.244
R10273 GND.n4146 GND.n2047 240.244
R10274 GND.n4146 GND.n2048 240.244
R10275 GND.n2048 GND.n1555 240.244
R10276 GND.n4695 GND.n1555 240.244
R10277 GND.n4695 GND.n1558 240.244
R10278 GND.n4691 GND.n1558 240.244
R10279 GND.n4691 GND.n1564 240.244
R10280 GND.n1833 GND.n1564 240.244
R10281 GND.n1834 GND.n1833 240.244
R10282 GND.n1835 GND.n1834 240.244
R10283 GND.n1835 GND.n1826 240.244
R10284 GND.n1841 GND.n1826 240.244
R10285 GND.n1842 GND.n1841 240.244
R10286 GND.n1843 GND.n1842 240.244
R10287 GND.n1843 GND.n1822 240.244
R10288 GND.n1849 GND.n1822 240.244
R10289 GND.n1850 GND.n1849 240.244
R10290 GND.n1851 GND.n1850 240.244
R10291 GND.n1851 GND.n1818 240.244
R10292 GND.n1857 GND.n1818 240.244
R10293 GND.n1858 GND.n1857 240.244
R10294 GND.n1859 GND.n1858 240.244
R10295 GND.n1859 GND.n1814 240.244
R10296 GND.n1865 GND.n1814 240.244
R10297 GND.n1866 GND.n1865 240.244
R10298 GND.n1867 GND.n1866 240.244
R10299 GND.n1867 GND.n1810 240.244
R10300 GND.n1873 GND.n1810 240.244
R10301 GND.n1874 GND.n1873 240.244
R10302 GND.n1876 GND.n1874 240.244
R10303 GND.n1876 GND.n1875 240.244
R10304 GND.n1875 GND.n1806 240.244
R10305 GND.n1883 GND.n1806 240.244
R10306 GND.n1884 GND.n1883 240.244
R10307 GND.n1884 GND.n1802 240.244
R10308 GND.n4507 GND.n1802 240.244
R10309 GND.n4507 GND.n1804 240.244
R10310 GND.n4502 GND.n1804 240.244
R10311 GND.n4502 GND.n4501 240.244
R10312 GND.n4501 GND.n1889 240.244
R10313 GND.n4284 GND.n1889 240.244
R10314 GND.n4284 GND.n4281 240.244
R10315 GND.n4290 GND.n4281 240.244
R10316 GND.n4291 GND.n4290 240.244
R10317 GND.n4292 GND.n4291 240.244
R10318 GND.n4292 GND.n4276 240.244
R10319 GND.n4470 GND.n4276 240.244
R10320 GND.n4470 GND.n4277 240.244
R10321 GND.n4466 GND.n4277 240.244
R10322 GND.n4466 GND.n4465 240.244
R10323 GND.n4465 GND.n4464 240.244
R10324 GND.n4464 GND.n4300 240.244
R10325 GND.n4460 GND.n4300 240.244
R10326 GND.n4460 GND.n4459 240.244
R10327 GND.n4459 GND.n4458 240.244
R10328 GND.n4458 GND.n4306 240.244
R10329 GND.n4454 GND.n4306 240.244
R10330 GND.n4454 GND.n4453 240.244
R10331 GND.n4453 GND.n4452 240.244
R10332 GND.n4452 GND.n4312 240.244
R10333 GND.n4324 GND.n4312 240.244
R10334 GND.n4324 GND.n4323 240.244
R10335 GND.n4323 GND.n4322 240.244
R10336 GND.n4322 GND.n388 240.244
R10337 GND.n6157 GND.n388 240.244
R10338 GND.n6157 GND.n389 240.244
R10339 GND.n6153 GND.n389 240.244
R10340 GND.n6153 GND.n395 240.244
R10341 GND.n6149 GND.n395 240.244
R10342 GND.n6149 GND.n397 240.244
R10343 GND.n6145 GND.n397 240.244
R10344 GND.n6145 GND.n403 240.244
R10345 GND.n6141 GND.n403 240.244
R10346 GND.n6141 GND.n405 240.244
R10347 GND.n6137 GND.n405 240.244
R10348 GND.n6137 GND.n411 240.244
R10349 GND.n6133 GND.n411 240.244
R10350 GND.n6133 GND.n413 240.244
R10351 GND.n6129 GND.n413 240.244
R10352 GND.n6129 GND.n419 240.244
R10353 GND.n6125 GND.n419 240.244
R10354 GND.n6125 GND.n421 240.244
R10355 GND.n6121 GND.n421 240.244
R10356 GND.n6121 GND.n427 240.244
R10357 GND.n6117 GND.n427 240.244
R10358 GND.n6117 GND.n429 240.244
R10359 GND.n6113 GND.n429 240.244
R10360 GND.n6113 GND.n435 240.244
R10361 GND.n6109 GND.n435 240.244
R10362 GND.n6109 GND.n437 240.244
R10363 GND.n6105 GND.n437 240.244
R10364 GND.n6105 GND.n443 240.244
R10365 GND.n6101 GND.n443 240.244
R10366 GND.n6101 GND.n445 240.244
R10367 GND.n6097 GND.n445 240.244
R10368 GND.n6097 GND.n451 240.244
R10369 GND.n6093 GND.n451 240.244
R10370 GND.n6093 GND.n453 240.244
R10371 GND.n6089 GND.n453 240.244
R10372 GND.n6089 GND.n459 240.244
R10373 GND.n6085 GND.n459 240.244
R10374 GND.n6085 GND.n461 240.244
R10375 GND.n6081 GND.n461 240.244
R10376 GND.n6081 GND.n467 240.244
R10377 GND.n6077 GND.n467 240.244
R10378 GND.n6077 GND.n469 240.244
R10379 GND.n5241 GND.n972 240.244
R10380 GND.n5237 GND.n972 240.244
R10381 GND.n5237 GND.n974 240.244
R10382 GND.n5233 GND.n974 240.244
R10383 GND.n5233 GND.n979 240.244
R10384 GND.n5229 GND.n979 240.244
R10385 GND.n5229 GND.n981 240.244
R10386 GND.n5225 GND.n981 240.244
R10387 GND.n5225 GND.n987 240.244
R10388 GND.n5221 GND.n987 240.244
R10389 GND.n5221 GND.n989 240.244
R10390 GND.n5217 GND.n989 240.244
R10391 GND.n5217 GND.n995 240.244
R10392 GND.n5213 GND.n995 240.244
R10393 GND.n5213 GND.n997 240.244
R10394 GND.n5209 GND.n997 240.244
R10395 GND.n5209 GND.n1003 240.244
R10396 GND.n5205 GND.n1003 240.244
R10397 GND.n5205 GND.n1005 240.244
R10398 GND.n5201 GND.n1005 240.244
R10399 GND.n5201 GND.n1011 240.244
R10400 GND.n5197 GND.n1011 240.244
R10401 GND.n5197 GND.n1013 240.244
R10402 GND.n5193 GND.n1013 240.244
R10403 GND.n5193 GND.n1019 240.244
R10404 GND.n5189 GND.n1019 240.244
R10405 GND.n5189 GND.n1021 240.244
R10406 GND.n5185 GND.n1021 240.244
R10407 GND.n5185 GND.n1027 240.244
R10408 GND.n5181 GND.n1027 240.244
R10409 GND.n5181 GND.n1029 240.244
R10410 GND.n5177 GND.n1029 240.244
R10411 GND.n5177 GND.n1035 240.244
R10412 GND.n5173 GND.n1035 240.244
R10413 GND.n5173 GND.n1037 240.244
R10414 GND.n5169 GND.n1037 240.244
R10415 GND.n5169 GND.n1043 240.244
R10416 GND.n5165 GND.n1043 240.244
R10417 GND.n5165 GND.n1045 240.244
R10418 GND.n5161 GND.n1045 240.244
R10419 GND.n5161 GND.n1051 240.244
R10420 GND.n5157 GND.n1051 240.244
R10421 GND.n5157 GND.n1053 240.244
R10422 GND.n5153 GND.n1053 240.244
R10423 GND.n5153 GND.n1059 240.244
R10424 GND.n5149 GND.n1059 240.244
R10425 GND.n5149 GND.n1061 240.244
R10426 GND.n5145 GND.n1061 240.244
R10427 GND.n5145 GND.n1067 240.244
R10428 GND.n5141 GND.n1067 240.244
R10429 GND.n5141 GND.n1069 240.244
R10430 GND.n5137 GND.n1069 240.244
R10431 GND.n5137 GND.n1075 240.244
R10432 GND.n5133 GND.n1075 240.244
R10433 GND.n5133 GND.n1077 240.244
R10434 GND.n1468 GND.n1465 240.244
R10435 GND.n1469 GND.n1468 240.244
R10436 GND.n2960 GND.n1469 240.244
R10437 GND.n2960 GND.n1472 240.244
R10438 GND.n1473 GND.n1472 240.244
R10439 GND.n1474 GND.n1473 240.244
R10440 GND.n2265 GND.n1474 240.244
R10441 GND.n2265 GND.n1477 240.244
R10442 GND.n1478 GND.n1477 240.244
R10443 GND.n1479 GND.n1478 240.244
R10444 GND.n2250 GND.n1479 240.244
R10445 GND.n2250 GND.n1482 240.244
R10446 GND.n1483 GND.n1482 240.244
R10447 GND.n1484 GND.n1483 240.244
R10448 GND.n2236 GND.n1484 240.244
R10449 GND.n2236 GND.n1487 240.244
R10450 GND.n1488 GND.n1487 240.244
R10451 GND.n1489 GND.n1488 240.244
R10452 GND.n2221 GND.n1489 240.244
R10453 GND.n2221 GND.n1492 240.244
R10454 GND.n1493 GND.n1492 240.244
R10455 GND.n1494 GND.n1493 240.244
R10456 GND.n2207 GND.n1494 240.244
R10457 GND.n2207 GND.n1497 240.244
R10458 GND.n1498 GND.n1497 240.244
R10459 GND.n1499 GND.n1498 240.244
R10460 GND.n2191 GND.n1499 240.244
R10461 GND.n2191 GND.n1502 240.244
R10462 GND.n1503 GND.n1502 240.244
R10463 GND.n1504 GND.n1503 240.244
R10464 GND.n2176 GND.n1504 240.244
R10465 GND.n2176 GND.n1507 240.244
R10466 GND.n1508 GND.n1507 240.244
R10467 GND.n1509 GND.n1508 240.244
R10468 GND.n2162 GND.n1509 240.244
R10469 GND.n2162 GND.n1512 240.244
R10470 GND.n1513 GND.n1512 240.244
R10471 GND.n1514 GND.n1513 240.244
R10472 GND.n2147 GND.n1514 240.244
R10473 GND.n2147 GND.n1517 240.244
R10474 GND.n1518 GND.n1517 240.244
R10475 GND.n1519 GND.n1518 240.244
R10476 GND.n2134 GND.n1519 240.244
R10477 GND.n2134 GND.n1522 240.244
R10478 GND.n1523 GND.n1522 240.244
R10479 GND.n1524 GND.n1523 240.244
R10480 GND.n2119 GND.n1524 240.244
R10481 GND.n2119 GND.n1527 240.244
R10482 GND.n1528 GND.n1527 240.244
R10483 GND.n1529 GND.n1528 240.244
R10484 GND.n2104 GND.n1529 240.244
R10485 GND.n2104 GND.n1532 240.244
R10486 GND.n1533 GND.n1532 240.244
R10487 GND.n1534 GND.n1533 240.244
R10488 GND.n2091 GND.n1534 240.244
R10489 GND.n2091 GND.n1537 240.244
R10490 GND.n1538 GND.n1537 240.244
R10491 GND.n1539 GND.n1538 240.244
R10492 GND.n2075 GND.n1539 240.244
R10493 GND.n2075 GND.n1542 240.244
R10494 GND.n1543 GND.n1542 240.244
R10495 GND.n1544 GND.n1543 240.244
R10496 GND.n2061 GND.n1544 240.244
R10497 GND.n2061 GND.n1547 240.244
R10498 GND.n1548 GND.n1547 240.244
R10499 GND.n1549 GND.n1548 240.244
R10500 GND.n2046 GND.n1549 240.244
R10501 GND.n2046 GND.n1552 240.244
R10502 GND.n4698 GND.n1552 240.244
R10503 GND.n1960 GND.n1553 240.244
R10504 GND.n1963 GND.n1962 240.244
R10505 GND.n1970 GND.n1969 240.244
R10506 GND.n1973 GND.n1972 240.244
R10507 GND.n1980 GND.n1979 240.244
R10508 GND.n1983 GND.n1982 240.244
R10509 GND.n1999 GND.n1998 240.244
R10510 GND.n2002 GND.n2001 240.244
R10511 GND.n2018 GND.n2017 240.244
R10512 GND.n2021 GND.n2020 240.244
R10513 GND.n2037 GND.n2036 240.244
R10514 GND.n3878 GND.n1446 240.244
R10515 GND.n3878 GND.n2958 240.244
R10516 GND.n3888 GND.n2958 240.244
R10517 GND.n3888 GND.n2954 240.244
R10518 GND.n3894 GND.n2954 240.244
R10519 GND.n3894 GND.n2263 240.244
R10520 GND.n3904 GND.n2263 240.244
R10521 GND.n3904 GND.n2259 240.244
R10522 GND.n3910 GND.n2259 240.244
R10523 GND.n3910 GND.n2248 240.244
R10524 GND.n3920 GND.n2248 240.244
R10525 GND.n3920 GND.n2244 240.244
R10526 GND.n3926 GND.n2244 240.244
R10527 GND.n3926 GND.n2234 240.244
R10528 GND.n3936 GND.n2234 240.244
R10529 GND.n3936 GND.n2230 240.244
R10530 GND.n3942 GND.n2230 240.244
R10531 GND.n3942 GND.n2219 240.244
R10532 GND.n3952 GND.n2219 240.244
R10533 GND.n3952 GND.n2215 240.244
R10534 GND.n3958 GND.n2215 240.244
R10535 GND.n3958 GND.n2205 240.244
R10536 GND.n3968 GND.n2205 240.244
R10537 GND.n3968 GND.n2201 240.244
R10538 GND.n3974 GND.n2201 240.244
R10539 GND.n3974 GND.n2189 240.244
R10540 GND.n3984 GND.n2189 240.244
R10541 GND.n3984 GND.n2185 240.244
R10542 GND.n3990 GND.n2185 240.244
R10543 GND.n3990 GND.n2175 240.244
R10544 GND.n4000 GND.n2175 240.244
R10545 GND.n4000 GND.n2171 240.244
R10546 GND.n4006 GND.n2171 240.244
R10547 GND.n4006 GND.n2160 240.244
R10548 GND.n4016 GND.n2160 240.244
R10549 GND.n4016 GND.n2156 240.244
R10550 GND.n4022 GND.n2156 240.244
R10551 GND.n4022 GND.n2146 240.244
R10552 GND.n4032 GND.n2146 240.244
R10553 GND.n4032 GND.n2142 240.244
R10554 GND.n4038 GND.n2142 240.244
R10555 GND.n4038 GND.n2132 240.244
R10556 GND.n4048 GND.n2132 240.244
R10557 GND.n4048 GND.n2128 240.244
R10558 GND.n4054 GND.n2128 240.244
R10559 GND.n4054 GND.n2117 240.244
R10560 GND.n4064 GND.n2117 240.244
R10561 GND.n4064 GND.n2113 240.244
R10562 GND.n4070 GND.n2113 240.244
R10563 GND.n4070 GND.n2102 240.244
R10564 GND.n4080 GND.n2102 240.244
R10565 GND.n4080 GND.n2098 240.244
R10566 GND.n4086 GND.n2098 240.244
R10567 GND.n4086 GND.n2089 240.244
R10568 GND.n4095 GND.n2089 240.244
R10569 GND.n4095 GND.n2085 240.244
R10570 GND.n4101 GND.n2085 240.244
R10571 GND.n4101 GND.n2073 240.244
R10572 GND.n4111 GND.n2073 240.244
R10573 GND.n4111 GND.n2069 240.244
R10574 GND.n4117 GND.n2069 240.244
R10575 GND.n4117 GND.n2059 240.244
R10576 GND.n4127 GND.n2059 240.244
R10577 GND.n4127 GND.n2054 240.244
R10578 GND.n4135 GND.n2054 240.244
R10579 GND.n4135 GND.n2044 240.244
R10580 GND.n4148 GND.n2044 240.244
R10581 GND.n4149 GND.n4148 240.244
R10582 GND.n4149 GND.n1556 240.244
R10583 GND.n1464 GND.n1463 240.244
R10584 GND.n4805 GND.n1463 240.244
R10585 GND.n4807 GND.n4806 240.244
R10586 GND.n4811 GND.n4810 240.244
R10587 GND.n1450 GND.n1403 240.244
R10588 GND.n1453 GND.n1404 240.244
R10589 GND.n1415 GND.n1414 240.244
R10590 GND.n1455 GND.n1425 240.244
R10591 GND.n1458 GND.n1426 240.244
R10592 GND.n1436 GND.n1435 240.244
R10593 GND.n1461 GND.n1445 240.244
R10594 GND.n2022 GND.t53 240.219
R10595 GND.n4840 GND.t105 240.219
R10596 GND.n2304 GND.n2303 240.132
R10597 GND.n2302 GND.n2301 240.132
R10598 GND.n2530 GND.n2529 240.132
R10599 GND.n2528 GND.n2527 240.132
R10600 GND.n1311 GND.t43 227.928
R10601 GND.n1370 GND.t109 227.928
R10602 GND.n1396 GND.t99 227.928
R10603 GND.n1328 GND.t121 227.928
R10604 GND.n1929 GND.t102 227.928
R10605 GND.n1439 GND.t115 227.928
R10606 GND.n3296 GND.t70 227.928
R10607 GND.n1612 GND.t148 227.928
R10608 GND.n1628 GND.t96 227.928
R10609 GND.n1642 GND.t83 227.928
R10610 GND.n1656 GND.t87 227.928
R10611 GND.n380 GND.t77 227.928
R10612 GND.n6188 GND.t60 227.928
R10613 GND.n336 GND.t90 227.928
R10614 GND.n309 GND.t139 227.928
R10615 GND.n4391 GND.t93 227.928
R10616 GND.n3349 GND.t64 227.928
R10617 GND.n3418 GND.t151 227.928
R10618 GND.n3450 GND.t133 227.928
R10619 GND.n3309 GND.t33 227.928
R10620 GND.n2022 GND.t55 211.588
R10621 GND.n4840 GND.t108 211.588
R10622 GND.n1626 GND.n1575 199.319
R10623 GND.n1626 GND.n1576 199.319
R10624 GND.n4915 GND.n4914 199.319
R10625 GND.n2305 GND.n2300 186.49
R10626 GND.n2531 GND.n2526 186.49
R10627 GND.n69 GND.n68 185
R10628 GND.n67 GND.n66 185
R10629 GND.n58 GND.n57 185
R10630 GND.n61 GND.n60 185
R10631 GND.n49 GND.n48 185
R10632 GND.n47 GND.n46 185
R10633 GND.n38 GND.n37 185
R10634 GND.n41 GND.n40 185
R10635 GND.n30 GND.n29 185
R10636 GND.n28 GND.n27 185
R10637 GND.n19 GND.n18 185
R10638 GND.n22 GND.n21 185
R10639 GND.n128 GND.n127 185
R10640 GND.n126 GND.n125 185
R10641 GND.n117 GND.n116 185
R10642 GND.n120 GND.n119 185
R10643 GND.n108 GND.n107 185
R10644 GND.n106 GND.n105 185
R10645 GND.n97 GND.n96 185
R10646 GND.n100 GND.n99 185
R10647 GND.n89 GND.n88 185
R10648 GND.n87 GND.n86 185
R10649 GND.n78 GND.n77 185
R10650 GND.n81 GND.n80 185
R10651 GND.n1311 GND.t45 170.781
R10652 GND.n1370 GND.t110 170.781
R10653 GND.n1396 GND.t100 170.781
R10654 GND.n1328 GND.t122 170.781
R10655 GND.n1929 GND.t104 170.781
R10656 GND.n1439 GND.t116 170.781
R10657 GND.n3296 GND.t72 170.781
R10658 GND.n1612 GND.t150 170.781
R10659 GND.n1628 GND.t98 170.781
R10660 GND.n1642 GND.t86 170.781
R10661 GND.n1656 GND.t89 170.781
R10662 GND.n380 GND.t78 170.781
R10663 GND.n6188 GND.t62 170.781
R10664 GND.n336 GND.t91 170.781
R10665 GND.n309 GND.t140 170.781
R10666 GND.n4391 GND.t94 170.781
R10667 GND.n3349 GND.t66 170.781
R10668 GND.n3418 GND.t153 170.781
R10669 GND.n3450 GND.t135 170.781
R10670 GND.n3309 GND.t36 170.781
R10671 GND.n2670 GND.n2508 163.367
R10672 GND.n2666 GND.n2665 163.367
R10673 GND.n2663 GND.n2541 163.367
R10674 GND.n2659 GND.n2658 163.367
R10675 GND.n2656 GND.n2544 163.367
R10676 GND.n2652 GND.n2651 163.367
R10677 GND.n2649 GND.n2547 163.367
R10678 GND.n2645 GND.n2644 163.367
R10679 GND.n2642 GND.n2550 163.367
R10680 GND.n2638 GND.n2637 163.367
R10681 GND.n2635 GND.n2553 163.367
R10682 GND.n2631 GND.n2630 163.367
R10683 GND.n2627 GND.n2626 163.367
R10684 GND.n2624 GND.n2560 163.367
R10685 GND.n2620 GND.n2619 163.367
R10686 GND.n2617 GND.n2566 163.367
R10687 GND.n2613 GND.n2612 163.367
R10688 GND.n2610 GND.n2569 163.367
R10689 GND.n2606 GND.n2605 163.367
R10690 GND.n2603 GND.n2572 163.367
R10691 GND.n2599 GND.n2598 163.367
R10692 GND.n2596 GND.n2575 163.367
R10693 GND.n2592 GND.n2591 163.367
R10694 GND.n2589 GND.n2578 163.367
R10695 GND.n2847 GND.n2846 163.367
R10696 GND.n2846 GND.n2845 163.367
R10697 GND.n2845 GND.n2330 163.367
R10698 GND.n2340 GND.n2330 163.367
R10699 GND.n2836 GND.n2340 163.367
R10700 GND.n2836 GND.n2341 163.367
R10701 GND.n2832 GND.n2341 163.367
R10702 GND.n2832 GND.n2831 163.367
R10703 GND.n2831 GND.n2345 163.367
R10704 GND.n2353 GND.n2345 163.367
R10705 GND.n2821 GND.n2353 163.367
R10706 GND.n2821 GND.n2354 163.367
R10707 GND.n2817 GND.n2354 163.367
R10708 GND.n2817 GND.n2816 163.367
R10709 GND.n2816 GND.n2358 163.367
R10710 GND.n2368 GND.n2358 163.367
R10711 GND.n2807 GND.n2368 163.367
R10712 GND.n2807 GND.n2369 163.367
R10713 GND.n2803 GND.n2369 163.367
R10714 GND.n2803 GND.n2373 163.367
R10715 GND.n2384 GND.n2373 163.367
R10716 GND.n2384 GND.n2382 163.367
R10717 GND.n2793 GND.n2382 163.367
R10718 GND.n2793 GND.n2383 163.367
R10719 GND.n2789 GND.n2383 163.367
R10720 GND.n2789 GND.n2788 163.367
R10721 GND.n2788 GND.n2787 163.367
R10722 GND.n2787 GND.n2388 163.367
R10723 GND.n2783 GND.n2388 163.367
R10724 GND.n2783 GND.n2782 163.367
R10725 GND.n2782 GND.n2781 163.367
R10726 GND.n2781 GND.n2390 163.367
R10727 GND.n2412 GND.n2390 163.367
R10728 GND.n2771 GND.n2412 163.367
R10729 GND.n2771 GND.n2413 163.367
R10730 GND.n2767 GND.n2413 163.367
R10731 GND.n2767 GND.n2766 163.367
R10732 GND.n2766 GND.n2417 163.367
R10733 GND.n2425 GND.n2417 163.367
R10734 GND.n2756 GND.n2425 163.367
R10735 GND.n2756 GND.n2426 163.367
R10736 GND.n2752 GND.n2426 163.367
R10737 GND.n2752 GND.n2751 163.367
R10738 GND.n2751 GND.n2430 163.367
R10739 GND.n2439 GND.n2430 163.367
R10740 GND.n2741 GND.n2439 163.367
R10741 GND.n2741 GND.n2440 163.367
R10742 GND.n2737 GND.n2440 163.367
R10743 GND.n2737 GND.n2736 163.367
R10744 GND.n2736 GND.n2444 163.367
R10745 GND.n2452 GND.n2444 163.367
R10746 GND.n2726 GND.n2452 163.367
R10747 GND.n2726 GND.n2453 163.367
R10748 GND.n2722 GND.n2453 163.367
R10749 GND.n2722 GND.n2721 163.367
R10750 GND.n2721 GND.n2457 163.367
R10751 GND.n2467 GND.n2457 163.367
R10752 GND.n2712 GND.n2467 163.367
R10753 GND.n2712 GND.n2468 163.367
R10754 GND.n2708 GND.n2468 163.367
R10755 GND.n2708 GND.n2707 163.367
R10756 GND.n2707 GND.n2472 163.367
R10757 GND.n2481 GND.n2472 163.367
R10758 GND.n2698 GND.n2481 163.367
R10759 GND.n2698 GND.n2482 163.367
R10760 GND.n2694 GND.n2482 163.367
R10761 GND.n2694 GND.n2486 163.367
R10762 GND.n2495 GND.n2486 163.367
R10763 GND.n2495 GND.n2493 163.367
R10764 GND.n2683 GND.n2493 163.367
R10765 GND.n2683 GND.n2494 163.367
R10766 GND.n2679 GND.n2494 163.367
R10767 GND.n2679 GND.n2678 163.367
R10768 GND.n2678 GND.n2499 163.367
R10769 GND.n2583 GND.n2499 163.367
R10770 GND.n2584 GND.n2583 163.367
R10771 GND.n2292 GND.n2291 163.367
R10772 GND.n2940 GND.n2291 163.367
R10773 GND.n2938 GND.n2937 163.367
R10774 GND.n2934 GND.n2933 163.367
R10775 GND.n2930 GND.n2929 163.367
R10776 GND.n2926 GND.n2925 163.367
R10777 GND.n2922 GND.n2921 163.367
R10778 GND.n2918 GND.n2917 163.367
R10779 GND.n2914 GND.n2913 163.367
R10780 GND.n2910 GND.n2909 163.367
R10781 GND.n2905 GND.n2904 163.367
R10782 GND.n2901 GND.n2900 163.367
R10783 GND.n2895 GND.n2894 163.367
R10784 GND.n2891 GND.n2890 163.367
R10785 GND.n2886 GND.n2885 163.367
R10786 GND.n2882 GND.n2881 163.367
R10787 GND.n2878 GND.n2877 163.367
R10788 GND.n2874 GND.n2873 163.367
R10789 GND.n2870 GND.n2869 163.367
R10790 GND.n2866 GND.n2865 163.367
R10791 GND.n2862 GND.n2861 163.367
R10792 GND.n2858 GND.n2857 163.367
R10793 GND.n2854 GND.n2853 163.367
R10794 GND.n2850 GND.n2289 163.367
R10795 GND.n2333 GND.n2293 163.367
R10796 GND.n2843 GND.n2333 163.367
R10797 GND.n2843 GND.n2334 163.367
R10798 GND.n2839 GND.n2334 163.367
R10799 GND.n2839 GND.n2838 163.367
R10800 GND.n2838 GND.n2338 163.367
R10801 GND.n2347 GND.n2338 163.367
R10802 GND.n2829 GND.n2347 163.367
R10803 GND.n2829 GND.n2348 163.367
R10804 GND.n2825 GND.n2348 163.367
R10805 GND.n2825 GND.n2352 163.367
R10806 GND.n2362 GND.n2352 163.367
R10807 GND.n2362 GND.n2360 163.367
R10808 GND.n2814 GND.n2360 163.367
R10809 GND.n2814 GND.n2361 163.367
R10810 GND.n2810 GND.n2361 163.367
R10811 GND.n2810 GND.n2809 163.367
R10812 GND.n2809 GND.n2366 163.367
R10813 GND.n2801 GND.n2366 163.367
R10814 GND.n2801 GND.n2376 163.367
R10815 GND.n2797 GND.n2376 163.367
R10816 GND.n2797 GND.n2796 163.367
R10817 GND.n2796 GND.n2795 163.367
R10818 GND.n2795 GND.n2379 163.367
R10819 GND.n2399 GND.n2379 163.367
R10820 GND.n2399 GND.n2397 163.367
R10821 GND.n2403 GND.n2397 163.367
R10822 GND.n2406 GND.n2403 163.367
R10823 GND.n2407 GND.n2406 163.367
R10824 GND.n2407 GND.n2393 163.367
R10825 GND.n2779 GND.n2393 163.367
R10826 GND.n2779 GND.n2395 163.367
R10827 GND.n2775 GND.n2395 163.367
R10828 GND.n2775 GND.n2774 163.367
R10829 GND.n2774 GND.n2411 163.367
R10830 GND.n2419 GND.n2411 163.367
R10831 GND.n2764 GND.n2419 163.367
R10832 GND.n2764 GND.n2420 163.367
R10833 GND.n2760 GND.n2420 163.367
R10834 GND.n2760 GND.n2759 163.367
R10835 GND.n2759 GND.n2424 163.367
R10836 GND.n2432 GND.n2424 163.367
R10837 GND.n2749 GND.n2432 163.367
R10838 GND.n2749 GND.n2434 163.367
R10839 GND.n2745 GND.n2434 163.367
R10840 GND.n2745 GND.n2744 163.367
R10841 GND.n2744 GND.n2438 163.367
R10842 GND.n2446 GND.n2438 163.367
R10843 GND.n2734 GND.n2446 163.367
R10844 GND.n2734 GND.n2447 163.367
R10845 GND.n2730 GND.n2447 163.367
R10846 GND.n2730 GND.n2451 163.367
R10847 GND.n2461 GND.n2451 163.367
R10848 GND.n2461 GND.n2459 163.367
R10849 GND.n2719 GND.n2459 163.367
R10850 GND.n2719 GND.n2460 163.367
R10851 GND.n2715 GND.n2460 163.367
R10852 GND.n2715 GND.n2714 163.367
R10853 GND.n2714 GND.n2465 163.367
R10854 GND.n2474 GND.n2465 163.367
R10855 GND.n2705 GND.n2474 163.367
R10856 GND.n2705 GND.n2475 163.367
R10857 GND.n2701 GND.n2475 163.367
R10858 GND.n2701 GND.n2700 163.367
R10859 GND.n2700 GND.n2479 163.367
R10860 GND.n2692 GND.n2479 163.367
R10861 GND.n2692 GND.n2489 163.367
R10862 GND.n2688 GND.n2489 163.367
R10863 GND.n2688 GND.n2687 163.367
R10864 GND.n2687 GND.n2492 163.367
R10865 GND.n2504 GND.n2492 163.367
R10866 GND.n2504 GND.n2501 163.367
R10867 GND.n2676 GND.n2501 163.367
R10868 GND.n2676 GND.n2502 163.367
R10869 GND.n2672 GND.n2502 163.367
R10870 GND.n2672 GND.n2671 163.367
R10871 GND.n2537 GND.n2536 157.237
R10872 GND.n53 GND.n33 156.846
R10873 GND.n73 GND.n72 155.571
R10874 GND.n53 GND.n52 155.571
R10875 GND.n2310 GND.n2309 152
R10876 GND.n2311 GND.n2298 152
R10877 GND.n2313 GND.n2312 152
R10878 GND.n2316 GND.n2315 152
R10879 GND.n2317 GND.n2296 152
R10880 GND.n2319 GND.n2318 152
R10881 GND.n2321 GND.n2294 152
R10882 GND.n2323 GND.n2322 152
R10883 GND.n2535 GND.n2509 152
R10884 GND.n2525 GND.n2510 152
R10885 GND.n2524 GND.n2523 152
R10886 GND.n2522 GND.n2511 152
R10887 GND.n2519 GND.n2512 152
R10888 GND.n2518 GND.n2517 152
R10889 GND.n2516 GND.n2513 152
R10890 GND.n2514 GND.t57 149.72
R10891 GND.t171 GND.n59 147.888
R10892 GND.t167 GND.n39 147.888
R10893 GND.t163 GND.n20 147.888
R10894 GND.t169 GND.n118 147.888
R10895 GND.t161 GND.n98 147.888
R10896 GND.t165 GND.n79 147.888
R10897 GND.n2023 GND.t56 145.649
R10898 GND.n4841 GND.t107 145.649
R10899 GND.n2629 GND.n2628 143.351
R10900 GND.n2897 GND.n2276 143.351
R10901 GND.n2897 GND.n2277 143.351
R10902 GND.n2307 GND.t118 129.018
R10903 GND.n2322 GND.t130 126.766
R10904 GND.n2320 GND.t50 126.766
R10905 GND.n2296 GND.t145 126.766
R10906 GND.n2314 GND.t40 126.766
R10907 GND.n2298 GND.t124 126.766
R10908 GND.n2308 GND.t67 126.766
R10909 GND.n2515 GND.t136 126.766
R10910 GND.n2517 GND.t30 126.766
R10911 GND.n2521 GND.t112 126.766
R10912 GND.n2523 GND.t47 126.766
R10913 GND.n2534 GND.t127 126.766
R10914 GND.n2536 GND.t80 126.766
R10915 GND.n2327 GND.t39 121.246
R10916 GND.n2561 GND.t75 121.246
R10917 GND.n2325 GND.t29 121.242
R10918 GND.n2554 GND.t143 121.242
R10919 GND.n68 GND.n67 104.615
R10920 GND.n67 GND.n57 104.615
R10921 GND.n60 GND.n57 104.615
R10922 GND.n48 GND.n47 104.615
R10923 GND.n47 GND.n37 104.615
R10924 GND.n40 GND.n37 104.615
R10925 GND.n29 GND.n28 104.615
R10926 GND.n28 GND.n18 104.615
R10927 GND.n21 GND.n18 104.615
R10928 GND.n127 GND.n126 104.615
R10929 GND.n126 GND.n116 104.615
R10930 GND.n119 GND.n116 104.615
R10931 GND.n107 GND.n106 104.615
R10932 GND.n106 GND.n96 104.615
R10933 GND.n99 GND.n96 104.615
R10934 GND.n88 GND.n87 104.615
R10935 GND.n87 GND.n77 104.615
R10936 GND.n80 GND.n77 104.615
R10937 GND.n6254 GND.n6253 99.6594
R10938 GND.n6251 GND.n6250 99.6594
R10939 GND.n6246 GND.n303 99.6594
R10940 GND.n6244 GND.n6243 99.6594
R10941 GND.n6239 GND.n312 99.6594
R10942 GND.n6237 GND.n6236 99.6594
R10943 GND.n6232 GND.n319 99.6594
R10944 GND.n6230 GND.n6229 99.6594
R10945 GND.n6225 GND.n326 99.6594
R10946 GND.n6223 GND.n6222 99.6594
R10947 GND.n6218 GND.n333 99.6594
R10948 GND.n6216 GND.n6215 99.6594
R10949 GND.n6209 GND.n341 99.6594
R10950 GND.n6207 GND.n6206 99.6594
R10951 GND.n6202 GND.n347 99.6594
R10952 GND.n6200 GND.n6199 99.6594
R10953 GND.n6195 GND.n354 99.6594
R10954 GND.n6193 GND.n6192 99.6594
R10955 GND.n6185 GND.n361 99.6594
R10956 GND.n6183 GND.n6182 99.6594
R10957 GND.n6178 GND.n368 99.6594
R10958 GND.n6176 GND.n6175 99.6594
R10959 GND.n6171 GND.n375 99.6594
R10960 GND.n6169 GND.n6168 99.6594
R10961 GND.n385 GND.n384 99.6594
R10962 GND.n4687 GND.n4686 99.6594
R10963 GND.n4681 GND.n1566 99.6594
R10964 GND.n4678 GND.n1567 99.6594
R10965 GND.n4674 GND.n1568 99.6594
R10966 GND.n4670 GND.n1569 99.6594
R10967 GND.n4666 GND.n1570 99.6594
R10968 GND.n4663 GND.n1571 99.6594
R10969 GND.n4659 GND.n1572 99.6594
R10970 GND.n4655 GND.n1573 99.6594
R10971 GND.n4651 GND.n1574 99.6594
R10972 GND.n4647 GND.n1575 99.6594
R10973 GND.n4642 GND.n1577 99.6594
R10974 GND.n4638 GND.n1578 99.6594
R10975 GND.n4634 GND.n1579 99.6594
R10976 GND.n4630 GND.n1580 99.6594
R10977 GND.n4626 GND.n1581 99.6594
R10978 GND.n4622 GND.n1582 99.6594
R10979 GND.n4617 GND.n1583 99.6594
R10980 GND.n4613 GND.n1584 99.6594
R10981 GND.n4609 GND.n1585 99.6594
R10982 GND.n4605 GND.n1586 99.6594
R10983 GND.n4601 GND.n1587 99.6594
R10984 GND.n4597 GND.n1588 99.6594
R10985 GND.n1345 GND.n1301 99.6594
R10986 GND.n1344 GND.n1304 99.6594
R10987 GND.n1342 GND.n1306 99.6594
R10988 GND.n1341 GND.n1309 99.6594
R10989 GND.n1339 GND.n1314 99.6594
R10990 GND.n1338 GND.n1337 99.6594
R10991 GND.n1336 GND.n1319 99.6594
R10992 GND.n1335 GND.n1334 99.6594
R10993 GND.n1333 GND.n1324 99.6594
R10994 GND.n1332 GND.n1331 99.6594
R10995 GND.n4914 GND.n4913 99.6594
R10996 GND.n4911 GND.n4910 99.6594
R10997 GND.n1353 GND.n1352 99.6594
R10998 GND.n1356 GND.n1355 99.6594
R10999 GND.n1361 GND.n1360 99.6594
R11000 GND.n1364 GND.n1363 99.6594
R11001 GND.n1369 GND.n1368 99.6594
R11002 GND.n1374 GND.n1373 99.6594
R11003 GND.n1379 GND.n1378 99.6594
R11004 GND.n1382 GND.n1381 99.6594
R11005 GND.n1387 GND.n1386 99.6594
R11006 GND.n1390 GND.n1389 99.6594
R11007 GND.n1395 GND.n1394 99.6594
R11008 GND.n1398 GND.n1289 99.6594
R11009 GND.n3362 GND.n1167 99.6594
R11010 GND.n3370 GND.n3369 99.6594
R11011 GND.n3373 GND.n3372 99.6594
R11012 GND.n3380 GND.n3379 99.6594
R11013 GND.n3383 GND.n3382 99.6594
R11014 GND.n3390 GND.n3389 99.6594
R11015 GND.n3393 GND.n3392 99.6594
R11016 GND.n3400 GND.n3399 99.6594
R11017 GND.n3403 GND.n3402 99.6594
R11018 GND.n3410 GND.n3409 99.6594
R11019 GND.n3413 GND.n3412 99.6594
R11020 GND.n3422 GND.n3421 99.6594
R11021 GND.n3425 GND.n3424 99.6594
R11022 GND.n3432 GND.n3431 99.6594
R11023 GND.n3435 GND.n3434 99.6594
R11024 GND.n3442 GND.n3441 99.6594
R11025 GND.n3445 GND.n3444 99.6594
R11026 GND.n3455 GND.n3454 99.6594
R11027 GND.n3458 GND.n3457 99.6594
R11028 GND.n3465 GND.n3464 99.6594
R11029 GND.n3468 GND.n3467 99.6594
R11030 GND.n3475 GND.n3474 99.6594
R11031 GND.n3478 GND.n3477 99.6594
R11032 GND.n3485 GND.n3484 99.6594
R11033 GND.n4407 GND.n4402 99.6594
R11034 GND.n4411 GND.n4409 99.6594
R11035 GND.n4417 GND.n4398 99.6594
R11036 GND.n4421 GND.n4419 99.6594
R11037 GND.n4427 GND.n4394 99.6594
R11038 GND.n4430 GND.n4429 99.6594
R11039 GND.n1667 GND.n1596 99.6594
R11040 GND.n1990 GND.n1595 99.6594
R11041 GND.n1992 GND.n1594 99.6594
R11042 GND.n2009 GND.n1593 99.6594
R11043 GND.n2011 GND.n1592 99.6594
R11044 GND.n1928 GND.n1591 99.6594
R11045 GND.n1410 GND.n1409 99.6594
R11046 GND.n1419 GND.n1418 99.6594
R11047 GND.n1422 GND.n1421 99.6594
R11048 GND.n1431 GND.n1430 99.6594
R11049 GND.n1442 GND.n1441 99.6594
R11050 GND.n4834 GND.n4833 99.6594
R11051 GND.n3497 GND.n3496 99.6594
R11052 GND.n3500 GND.n3499 99.6594
R11053 GND.n3507 GND.n3506 99.6594
R11054 GND.n3510 GND.n3509 99.6594
R11055 GND.n3518 GND.n3517 99.6594
R11056 GND.n3521 GND.n3520 99.6594
R11057 GND.n3498 GND.n3497 99.6594
R11058 GND.n3499 GND.n3304 99.6594
R11059 GND.n3508 GND.n3507 99.6594
R11060 GND.n3509 GND.n3300 99.6594
R11061 GND.n3519 GND.n3518 99.6594
R11062 GND.n3522 GND.n3521 99.6594
R11063 GND.n4833 GND.n1443 99.6594
R11064 GND.n1441 GND.n1432 99.6594
R11065 GND.n1430 GND.n1429 99.6594
R11066 GND.n1421 GND.n1420 99.6594
R11067 GND.n1418 GND.n1411 99.6594
R11068 GND.n1409 GND.n1408 99.6594
R11069 GND.n1989 GND.n1596 99.6594
R11070 GND.n1993 GND.n1595 99.6594
R11071 GND.n2008 GND.n1594 99.6594
R11072 GND.n2012 GND.n1593 99.6594
R11073 GND.n1932 GND.n1592 99.6594
R11074 GND.n2031 GND.n1591 99.6594
R11075 GND.n4429 GND.n4428 99.6594
R11076 GND.n4420 GND.n4394 99.6594
R11077 GND.n4419 GND.n4418 99.6594
R11078 GND.n4410 GND.n4398 99.6594
R11079 GND.n4409 GND.n4408 99.6594
R11080 GND.n4403 GND.n4402 99.6594
R11081 GND.n3363 GND.n3362 99.6594
R11082 GND.n3371 GND.n3370 99.6594
R11083 GND.n3372 GND.n3354 99.6594
R11084 GND.n3381 GND.n3380 99.6594
R11085 GND.n3382 GND.n3348 99.6594
R11086 GND.n3391 GND.n3390 99.6594
R11087 GND.n3392 GND.n3344 99.6594
R11088 GND.n3401 GND.n3400 99.6594
R11089 GND.n3402 GND.n3340 99.6594
R11090 GND.n3411 GND.n3410 99.6594
R11091 GND.n3412 GND.n3336 99.6594
R11092 GND.n3423 GND.n3422 99.6594
R11093 GND.n3424 GND.n3332 99.6594
R11094 GND.n3433 GND.n3432 99.6594
R11095 GND.n3434 GND.n3328 99.6594
R11096 GND.n3443 GND.n3442 99.6594
R11097 GND.n3444 GND.n3324 99.6594
R11098 GND.n3456 GND.n3455 99.6594
R11099 GND.n3457 GND.n3320 99.6594
R11100 GND.n3466 GND.n3465 99.6594
R11101 GND.n3467 GND.n3316 99.6594
R11102 GND.n3476 GND.n3475 99.6594
R11103 GND.n3477 GND.n3312 99.6594
R11104 GND.n3486 GND.n3485 99.6594
R11105 GND.n1399 GND.n1398 99.6594
R11106 GND.n1394 GND.n1393 99.6594
R11107 GND.n1389 GND.n1388 99.6594
R11108 GND.n1386 GND.n1385 99.6594
R11109 GND.n1381 GND.n1380 99.6594
R11110 GND.n1378 GND.n1377 99.6594
R11111 GND.n1373 GND.n1372 99.6594
R11112 GND.n1368 GND.n1367 99.6594
R11113 GND.n1363 GND.n1362 99.6594
R11114 GND.n1360 GND.n1359 99.6594
R11115 GND.n1355 GND.n1354 99.6594
R11116 GND.n1352 GND.n1348 99.6594
R11117 GND.n4912 GND.n4911 99.6594
R11118 GND.n4916 GND.n4915 99.6594
R11119 GND.n1332 GND.n1325 99.6594
R11120 GND.n1333 GND.n1323 99.6594
R11121 GND.n1335 GND.n1320 99.6594
R11122 GND.n1336 GND.n1318 99.6594
R11123 GND.n1338 GND.n1315 99.6594
R11124 GND.n1339 GND.n1310 99.6594
R11125 GND.n1341 GND.n1340 99.6594
R11126 GND.n1342 GND.n1305 99.6594
R11127 GND.n1344 GND.n1343 99.6594
R11128 GND.n1345 GND.n1300 99.6594
R11129 GND.n4687 GND.n1598 99.6594
R11130 GND.n4679 GND.n1566 99.6594
R11131 GND.n4675 GND.n1567 99.6594
R11132 GND.n4671 GND.n1568 99.6594
R11133 GND.n1610 GND.n1569 99.6594
R11134 GND.n4664 GND.n1570 99.6594
R11135 GND.n4660 GND.n1571 99.6594
R11136 GND.n4656 GND.n1572 99.6594
R11137 GND.n4652 GND.n1573 99.6594
R11138 GND.n4648 GND.n1574 99.6594
R11139 GND.n4643 GND.n1576 99.6594
R11140 GND.n4639 GND.n1577 99.6594
R11141 GND.n4635 GND.n1578 99.6594
R11142 GND.n4631 GND.n1579 99.6594
R11143 GND.n4627 GND.n1580 99.6594
R11144 GND.n4623 GND.n1581 99.6594
R11145 GND.n4618 GND.n1582 99.6594
R11146 GND.n4614 GND.n1583 99.6594
R11147 GND.n4610 GND.n1584 99.6594
R11148 GND.n4606 GND.n1585 99.6594
R11149 GND.n4602 GND.n1586 99.6594
R11150 GND.n4598 GND.n1587 99.6594
R11151 GND.n1655 GND.n1588 99.6594
R11152 GND.n384 GND.n376 99.6594
R11153 GND.n6170 GND.n6169 99.6594
R11154 GND.n375 GND.n369 99.6594
R11155 GND.n6177 GND.n6176 99.6594
R11156 GND.n368 GND.n362 99.6594
R11157 GND.n6184 GND.n6183 99.6594
R11158 GND.n361 GND.n355 99.6594
R11159 GND.n6194 GND.n6193 99.6594
R11160 GND.n354 GND.n348 99.6594
R11161 GND.n6201 GND.n6200 99.6594
R11162 GND.n347 GND.n342 99.6594
R11163 GND.n6208 GND.n6207 99.6594
R11164 GND.n341 GND.n334 99.6594
R11165 GND.n6217 GND.n6216 99.6594
R11166 GND.n333 GND.n327 99.6594
R11167 GND.n6224 GND.n6223 99.6594
R11168 GND.n326 GND.n320 99.6594
R11169 GND.n6231 GND.n6230 99.6594
R11170 GND.n319 GND.n313 99.6594
R11171 GND.n6238 GND.n6237 99.6594
R11172 GND.n312 GND.n304 99.6594
R11173 GND.n6245 GND.n6244 99.6594
R11174 GND.n303 GND.n297 99.6594
R11175 GND.n6252 GND.n6251 99.6594
R11176 GND.n6255 GND.n6254 99.6594
R11177 GND.n1963 GND.n1961 99.6594
R11178 GND.n1969 GND.n1954 99.6594
R11179 GND.n1973 GND.n1971 99.6594
R11180 GND.n1979 GND.n1950 99.6594
R11181 GND.n1983 GND.n1981 99.6594
R11182 GND.n1998 GND.n1942 99.6594
R11183 GND.n2002 GND.n2000 99.6594
R11184 GND.n2017 GND.n1935 99.6594
R11185 GND.n2021 GND.n2019 99.6594
R11186 GND.n2036 GND.n1925 99.6594
R11187 GND.n2039 GND.n2038 99.6594
R11188 GND.n2038 GND.n2037 99.6594
R11189 GND.n2020 GND.n1925 99.6594
R11190 GND.n2019 GND.n2018 99.6594
R11191 GND.n2001 GND.n1935 99.6594
R11192 GND.n2000 GND.n1999 99.6594
R11193 GND.n1982 GND.n1942 99.6594
R11194 GND.n1981 GND.n1980 99.6594
R11195 GND.n1972 GND.n1950 99.6594
R11196 GND.n1971 GND.n1970 99.6594
R11197 GND.n1962 GND.n1954 99.6594
R11198 GND.n1961 GND.n1960 99.6594
R11199 GND.n4825 GND.n4824 99.6594
R11200 GND.n4805 GND.n1448 99.6594
R11201 GND.n4807 GND.n1449 99.6594
R11202 GND.n4811 GND.n1451 99.6594
R11203 GND.n1452 GND.n1403 99.6594
R11204 GND.n1454 GND.n1453 99.6594
R11205 GND.n1456 GND.n1415 99.6594
R11206 GND.n1457 GND.n1425 99.6594
R11207 GND.n1459 GND.n1458 99.6594
R11208 GND.n1462 GND.n1461 99.6594
R11209 GND.n4827 GND.n1445 99.6594
R11210 GND.n1462 GND.n1436 99.6594
R11211 GND.n4828 GND.n4827 99.6594
R11212 GND.n4825 GND.n1464 99.6594
R11213 GND.n4806 GND.n1448 99.6594
R11214 GND.n4810 GND.n1449 99.6594
R11215 GND.n1451 GND.n1450 99.6594
R11216 GND.n1452 GND.n1404 99.6594
R11217 GND.n1454 GND.n1414 99.6594
R11218 GND.n1456 GND.n1455 99.6594
R11219 GND.n1457 GND.n1426 99.6594
R11220 GND.n1459 GND.n1435 99.6594
R11221 GND.n1312 GND.n1311 96.5823
R11222 GND.n1371 GND.n1370 96.5823
R11223 GND.n1397 GND.n1396 96.5823
R11224 GND.n1329 GND.n1328 96.5823
R11225 GND.n1930 GND.n1929 96.5823
R11226 GND.n1440 GND.n1439 96.5823
R11227 GND.n3297 GND.n3296 96.5823
R11228 GND.n1613 GND.n1612 96.5823
R11229 GND.n1629 GND.n1628 96.5823
R11230 GND.n1643 GND.n1642 96.5823
R11231 GND.n1657 GND.n1656 96.5823
R11232 GND.n381 GND.n380 96.5823
R11233 GND.n6189 GND.n6188 96.5823
R11234 GND.n337 GND.n336 96.5823
R11235 GND.n310 GND.n309 96.5823
R11236 GND.n4392 GND.n4391 96.5823
R11237 GND.n3350 GND.n3349 96.5823
R11238 GND.n3419 GND.n3418 96.5823
R11239 GND.n3451 GND.n3450 96.5823
R11240 GND.n3310 GND.n3309 96.5823
R11241 GND.n2307 GND.n2306 83.3186
R11242 GND.n2898 GND.n1330 79.2965
R11243 GND.n4645 GND.n1625 79.2965
R11244 GND.n1312 GND.t46 74.1998
R11245 GND.n1371 GND.t111 74.1998
R11246 GND.n1397 GND.t101 74.1998
R11247 GND.n1329 GND.t123 74.1998
R11248 GND.n1930 GND.t103 74.1998
R11249 GND.n1440 GND.t117 74.1998
R11250 GND.n3297 GND.t71 74.1998
R11251 GND.n1613 GND.t149 74.1998
R11252 GND.n1629 GND.t97 74.1998
R11253 GND.n1643 GND.t85 74.1998
R11254 GND.n1657 GND.t88 74.1998
R11255 GND.n381 GND.t79 74.1998
R11256 GND.n6189 GND.t63 74.1998
R11257 GND.n337 GND.t92 74.1998
R11258 GND.n310 GND.t141 74.1998
R11259 GND.n4392 GND.t95 74.1998
R11260 GND.n3350 GND.t65 74.1998
R11261 GND.n3419 GND.t152 74.1998
R11262 GND.n3451 GND.t134 74.1998
R11263 GND.n3310 GND.t35 74.1998
R11264 GND.n2308 GND.n2299 72.8411
R11265 GND.n2314 GND.n2297 72.8411
R11266 GND.n2320 GND.n2295 72.8411
R11267 GND.n2534 GND.n2533 72.8411
R11268 GND.n2521 GND.n2520 72.8411
R11269 GND.n2328 GND.t38 72.1784
R11270 GND.n2562 GND.t76 72.1784
R11271 GND.n2326 GND.t28 72.1745
R11272 GND.n2555 GND.t144 72.1745
R11273 GND.n3 GND.t178 72.1422
R11274 GND.n5 GND.t7 72.1422
R11275 GND.n8 GND.t25 72.1422
R11276 GND.n11 GND.t4 72.1422
R11277 GND.n1 GND.t10 72.1422
R11278 GND.n5126 GND.n1076 71.9952
R11279 GND.n6070 GND.n468 71.9952
R11280 GND.n2666 GND.n2540 71.676
R11281 GND.n2664 GND.n2663 71.676
R11282 GND.n2659 GND.n2543 71.676
R11283 GND.n2657 GND.n2656 71.676
R11284 GND.n2652 GND.n2546 71.676
R11285 GND.n2650 GND.n2649 71.676
R11286 GND.n2645 GND.n2549 71.676
R11287 GND.n2643 GND.n2642 71.676
R11288 GND.n2638 GND.n2552 71.676
R11289 GND.n2636 GND.n2635 71.676
R11290 GND.n2631 GND.n2558 71.676
R11291 GND.n2628 GND.n2627 71.676
R11292 GND.n2625 GND.n2624 71.676
R11293 GND.n2620 GND.n2564 71.676
R11294 GND.n2618 GND.n2617 71.676
R11295 GND.n2613 GND.n2568 71.676
R11296 GND.n2611 GND.n2610 71.676
R11297 GND.n2606 GND.n2571 71.676
R11298 GND.n2604 GND.n2603 71.676
R11299 GND.n2599 GND.n2574 71.676
R11300 GND.n2597 GND.n2596 71.676
R11301 GND.n2592 GND.n2577 71.676
R11302 GND.n2590 GND.n2589 71.676
R11303 GND.n2585 GND.n2580 71.676
R11304 GND.n2946 GND.n2945 71.676
R11305 GND.n2940 GND.n2266 71.676
R11306 GND.n2937 GND.n2267 71.676
R11307 GND.n2933 GND.n2268 71.676
R11308 GND.n2929 GND.n2269 71.676
R11309 GND.n2925 GND.n2270 71.676
R11310 GND.n2921 GND.n2271 71.676
R11311 GND.n2917 GND.n2272 71.676
R11312 GND.n2913 GND.n2273 71.676
R11313 GND.n2909 GND.n2274 71.676
R11314 GND.n2904 GND.n2275 71.676
R11315 GND.n2900 GND.n2276 71.676
R11316 GND.n2894 GND.n2278 71.676
R11317 GND.n2890 GND.n2279 71.676
R11318 GND.n2885 GND.n2280 71.676
R11319 GND.n2881 GND.n2281 71.676
R11320 GND.n2877 GND.n2282 71.676
R11321 GND.n2873 GND.n2283 71.676
R11322 GND.n2869 GND.n2284 71.676
R11323 GND.n2865 GND.n2285 71.676
R11324 GND.n2861 GND.n2286 71.676
R11325 GND.n2857 GND.n2287 71.676
R11326 GND.n2853 GND.n2288 71.676
R11327 GND.n2946 GND.n2292 71.676
R11328 GND.n2938 GND.n2266 71.676
R11329 GND.n2934 GND.n2267 71.676
R11330 GND.n2930 GND.n2268 71.676
R11331 GND.n2926 GND.n2269 71.676
R11332 GND.n2922 GND.n2270 71.676
R11333 GND.n2918 GND.n2271 71.676
R11334 GND.n2914 GND.n2272 71.676
R11335 GND.n2910 GND.n2273 71.676
R11336 GND.n2905 GND.n2274 71.676
R11337 GND.n2901 GND.n2275 71.676
R11338 GND.n2895 GND.n2277 71.676
R11339 GND.n2891 GND.n2278 71.676
R11340 GND.n2886 GND.n2279 71.676
R11341 GND.n2882 GND.n2280 71.676
R11342 GND.n2878 GND.n2281 71.676
R11343 GND.n2874 GND.n2282 71.676
R11344 GND.n2870 GND.n2283 71.676
R11345 GND.n2866 GND.n2284 71.676
R11346 GND.n2862 GND.n2285 71.676
R11347 GND.n2858 GND.n2286 71.676
R11348 GND.n2854 GND.n2287 71.676
R11349 GND.n2850 GND.n2288 71.676
R11350 GND.n2580 GND.n2578 71.676
R11351 GND.n2591 GND.n2590 71.676
R11352 GND.n2577 GND.n2575 71.676
R11353 GND.n2598 GND.n2597 71.676
R11354 GND.n2574 GND.n2572 71.676
R11355 GND.n2605 GND.n2604 71.676
R11356 GND.n2571 GND.n2569 71.676
R11357 GND.n2612 GND.n2611 71.676
R11358 GND.n2568 GND.n2566 71.676
R11359 GND.n2619 GND.n2618 71.676
R11360 GND.n2564 GND.n2560 71.676
R11361 GND.n2626 GND.n2625 71.676
R11362 GND.n2630 GND.n2629 71.676
R11363 GND.n2558 GND.n2553 71.676
R11364 GND.n2637 GND.n2636 71.676
R11365 GND.n2552 GND.n2550 71.676
R11366 GND.n2644 GND.n2643 71.676
R11367 GND.n2549 GND.n2547 71.676
R11368 GND.n2651 GND.n2650 71.676
R11369 GND.n2546 GND.n2544 71.676
R11370 GND.n2658 GND.n2657 71.676
R11371 GND.n2543 GND.n2541 71.676
R11372 GND.n2665 GND.n2664 71.676
R11373 GND.n2540 GND.n2508 71.676
R11374 GND.n135 GND.t22 69.9957
R11375 GND.n137 GND.t21 69.9957
R11376 GND.n140 GND.t177 69.9957
R11377 GND.n143 GND.t158 69.9957
R11378 GND.n146 GND.t159 69.9957
R11379 GND.n135 GND.n134 66.4527
R11380 GND.n137 GND.n136 66.4527
R11381 GND.n140 GND.n139 66.4527
R11382 GND.n143 GND.n142 66.4527
R11383 GND.n146 GND.n145 66.4527
R11384 GND.n2023 GND.n2022 65.9399
R11385 GND.n4841 GND.n4840 65.9399
R11386 GND.n3 GND.n2 64.3061
R11387 GND.n5 GND.n4 64.3061
R11388 GND.n8 GND.n7 64.3061
R11389 GND.n11 GND.n10 64.3061
R11390 GND.n1 GND.n0 64.3061
R11391 GND.n2907 GND.n2326 59.5399
R11392 GND.n2888 GND.n2328 59.5399
R11393 GND.n2563 GND.n2562 59.5399
R11394 GND.n2556 GND.n2555 59.5399
R11395 GND.n2324 GND.n2323 58.4046
R11396 GND.n112 GND.n92 55.2221
R11397 GND.n2305 GND.n2304 54.358
R11398 GND.n2531 GND.n2530 54.358
R11399 GND.n132 GND.n131 53.946
R11400 GND.n112 GND.n111 53.946
R11401 GND.n2514 GND.n2513 52.3702
R11402 GND.n60 GND.t171 52.3082
R11403 GND.n40 GND.t167 52.3082
R11404 GND.n21 GND.t163 52.3082
R11405 GND.n119 GND.t169 52.3082
R11406 GND.n99 GND.t161 52.3082
R11407 GND.n80 GND.t165 52.3082
R11408 GND.n2326 GND.n2325 49.0672
R11409 GND.n2328 GND.n2327 49.0672
R11410 GND.n2562 GND.n2561 49.0672
R11411 GND.n2555 GND.n2554 49.0672
R11412 GND.n5240 GND.n5239 46.6107
R11413 GND.n5239 GND.n5238 46.6107
R11414 GND.n5238 GND.n973 46.6107
R11415 GND.n5232 GND.n973 46.6107
R11416 GND.n5232 GND.n5231 46.6107
R11417 GND.n5231 GND.n5230 46.6107
R11418 GND.n5230 GND.n980 46.6107
R11419 GND.n5224 GND.n980 46.6107
R11420 GND.n5224 GND.n5223 46.6107
R11421 GND.n5223 GND.n5222 46.6107
R11422 GND.n5222 GND.n988 46.6107
R11423 GND.n5216 GND.n988 46.6107
R11424 GND.n5216 GND.n5215 46.6107
R11425 GND.n5215 GND.n5214 46.6107
R11426 GND.n5214 GND.n996 46.6107
R11427 GND.n5208 GND.n996 46.6107
R11428 GND.n5208 GND.n5207 46.6107
R11429 GND.n5207 GND.n5206 46.6107
R11430 GND.n5206 GND.n1004 46.6107
R11431 GND.n5200 GND.n1004 46.6107
R11432 GND.n5200 GND.n5199 46.6107
R11433 GND.n5199 GND.n5198 46.6107
R11434 GND.n5198 GND.n1012 46.6107
R11435 GND.n5192 GND.n1012 46.6107
R11436 GND.n5192 GND.n5191 46.6107
R11437 GND.n5191 GND.n5190 46.6107
R11438 GND.n5190 GND.n1020 46.6107
R11439 GND.n5184 GND.n1020 46.6107
R11440 GND.n5184 GND.n5183 46.6107
R11441 GND.n5183 GND.n5182 46.6107
R11442 GND.n5182 GND.n1028 46.6107
R11443 GND.n5176 GND.n1028 46.6107
R11444 GND.n5176 GND.n5175 46.6107
R11445 GND.n5175 GND.n5174 46.6107
R11446 GND.n5174 GND.n1036 46.6107
R11447 GND.n5168 GND.n1036 46.6107
R11448 GND.n5168 GND.n5167 46.6107
R11449 GND.n5167 GND.n5166 46.6107
R11450 GND.n5166 GND.n1044 46.6107
R11451 GND.n5160 GND.n1044 46.6107
R11452 GND.n5160 GND.n5159 46.6107
R11453 GND.n5159 GND.n5158 46.6107
R11454 GND.n5158 GND.n1052 46.6107
R11455 GND.n5152 GND.n1052 46.6107
R11456 GND.n5152 GND.n5151 46.6107
R11457 GND.n5151 GND.n5150 46.6107
R11458 GND.n5150 GND.n1060 46.6107
R11459 GND.n5144 GND.n1060 46.6107
R11460 GND.n5144 GND.n5143 46.6107
R11461 GND.n5143 GND.n5142 46.6107
R11462 GND.n5142 GND.n1068 46.6107
R11463 GND.n5136 GND.n1068 46.6107
R11464 GND.n5136 GND.n5135 46.6107
R11465 GND.n5135 GND.n5134 46.6107
R11466 GND.n2308 GND.n2307 45.8904
R11467 GND.n2538 GND.n2537 44.3322
R11468 GND.n2321 GND.n2320 43.8187
R11469 GND.n2535 GND.n2534 43.8187
R11470 GND.n2024 GND.n2023 42.2793
R11471 GND.n4934 GND.n1312 42.2793
R11472 GND.n4892 GND.n1371 42.2793
R11473 GND.n4873 GND.n1397 42.2793
R11474 GND.n2030 GND.n1930 42.2793
R11475 GND.n4836 GND.n1440 42.2793
R11476 GND.n3298 GND.n3297 42.2793
R11477 GND.n4668 GND.n1613 42.2793
R11478 GND.n4620 GND.n1643 42.2793
R11479 GND.n1658 GND.n1657 42.2793
R11480 GND.n6166 GND.n381 42.2793
R11481 GND.n6190 GND.n6189 42.2793
R11482 GND.n6214 GND.n337 42.2793
R11483 GND.n311 GND.n310 42.2793
R11484 GND.n4393 GND.n4392 42.2793
R11485 GND.n3351 GND.n3350 42.2793
R11486 GND.n3420 GND.n3419 42.2793
R11487 GND.n3452 GND.n3451 42.2793
R11488 GND.n3311 GND.n3310 42.2793
R11489 GND.n4842 GND.n4841 42.2793
R11490 GND.n2306 GND.n2305 41.6274
R11491 GND.n2532 GND.n2531 41.6274
R11492 GND.n2315 GND.n2314 37.9763
R11493 GND.n2314 GND.n2313 37.9763
R11494 GND.n2521 GND.n2512 37.9763
R11495 GND.n2522 GND.n2521 37.9763
R11496 GND.n1330 GND.n1329 36.9518
R11497 GND.n4645 GND.n1629 36.9518
R11498 GND.n5126 GND.n5125 36.1788
R11499 GND.n5125 GND.n5124 36.1788
R11500 GND.n5124 GND.n1083 36.1788
R11501 GND.n5118 GND.n1083 36.1788
R11502 GND.n5118 GND.n5117 36.1788
R11503 GND.n5117 GND.n5116 36.1788
R11504 GND.n5116 GND.n1090 36.1788
R11505 GND.n5110 GND.n1090 36.1788
R11506 GND.n5110 GND.n5109 36.1788
R11507 GND.n5109 GND.n5108 36.1788
R11508 GND.n5108 GND.n1098 36.1788
R11509 GND.n5102 GND.n1098 36.1788
R11510 GND.n5102 GND.n5101 36.1788
R11511 GND.n5101 GND.n5100 36.1788
R11512 GND.n5100 GND.n1106 36.1788
R11513 GND.n5094 GND.n1106 36.1788
R11514 GND.n5094 GND.n5093 36.1788
R11515 GND.n5093 GND.n5092 36.1788
R11516 GND.n5092 GND.n1114 36.1788
R11517 GND.n5086 GND.n1114 36.1788
R11518 GND.n5086 GND.n5085 36.1788
R11519 GND.n5085 GND.n5084 36.1788
R11520 GND.n5084 GND.n1122 36.1788
R11521 GND.n5078 GND.n1122 36.1788
R11522 GND.n5078 GND.n5077 36.1788
R11523 GND.n5077 GND.n5076 36.1788
R11524 GND.n5076 GND.n1130 36.1788
R11525 GND.n5070 GND.n1130 36.1788
R11526 GND.n5070 GND.n5069 36.1788
R11527 GND.n5069 GND.n5068 36.1788
R11528 GND.n5068 GND.n1138 36.1788
R11529 GND.n5062 GND.n1138 36.1788
R11530 GND.n5062 GND.n5061 36.1788
R11531 GND.n5061 GND.n5060 36.1788
R11532 GND.n5060 GND.n1146 36.1788
R11533 GND.n5054 GND.n1146 36.1788
R11534 GND.n5054 GND.n5053 36.1788
R11535 GND.n5053 GND.n5052 36.1788
R11536 GND.n5052 GND.n1154 36.1788
R11537 GND.n5046 GND.n5045 36.1788
R11538 GND.n3165 GND.n1292 36.1788
R11539 GND.n3163 GND.n1447 36.1788
R11540 GND.n3157 GND.n1460 36.1788
R11541 GND.n3157 GND.n2966 36.1788
R11542 GND.n3879 GND.n2966 36.1788
R11543 GND.n3879 GND.n2959 36.1788
R11544 GND.n3887 GND.n2959 36.1788
R11545 GND.n3895 GND.n2953 36.1788
R11546 GND.n3895 GND.n2264 36.1788
R11547 GND.n3903 GND.n2264 36.1788
R11548 GND.n4126 GND.n2060 36.1788
R11549 GND.n4126 GND.n2053 36.1788
R11550 GND.n4136 GND.n2053 36.1788
R11551 GND.n4147 GND.n2045 36.1788
R11552 GND.n4147 GND.n1554 36.1788
R11553 GND.n4697 GND.n1554 36.1788
R11554 GND.n4697 GND.n4696 36.1788
R11555 GND.n4696 GND.n1557 36.1788
R11556 GND.n4690 GND.n4689 36.1788
R11557 GND.n1664 GND.n1590 36.1788
R11558 GND.n6158 GND.n387 36.1788
R11559 GND.n6152 GND.n6151 36.1788
R11560 GND.n6151 GND.n6150 36.1788
R11561 GND.n6150 GND.n396 36.1788
R11562 GND.n6144 GND.n396 36.1788
R11563 GND.n6144 GND.n6143 36.1788
R11564 GND.n6143 GND.n6142 36.1788
R11565 GND.n6142 GND.n404 36.1788
R11566 GND.n6136 GND.n404 36.1788
R11567 GND.n6136 GND.n6135 36.1788
R11568 GND.n6135 GND.n6134 36.1788
R11569 GND.n6134 GND.n412 36.1788
R11570 GND.n6128 GND.n412 36.1788
R11571 GND.n6128 GND.n6127 36.1788
R11572 GND.n6127 GND.n6126 36.1788
R11573 GND.n6126 GND.n420 36.1788
R11574 GND.n6120 GND.n420 36.1788
R11575 GND.n6120 GND.n6119 36.1788
R11576 GND.n6119 GND.n6118 36.1788
R11577 GND.n6118 GND.n428 36.1788
R11578 GND.n6112 GND.n428 36.1788
R11579 GND.n6112 GND.n6111 36.1788
R11580 GND.n6111 GND.n6110 36.1788
R11581 GND.n6110 GND.n436 36.1788
R11582 GND.n6104 GND.n436 36.1788
R11583 GND.n6104 GND.n6103 36.1788
R11584 GND.n6103 GND.n6102 36.1788
R11585 GND.n6102 GND.n444 36.1788
R11586 GND.n6096 GND.n444 36.1788
R11587 GND.n6096 GND.n6095 36.1788
R11588 GND.n6095 GND.n6094 36.1788
R11589 GND.n6094 GND.n452 36.1788
R11590 GND.n6088 GND.n452 36.1788
R11591 GND.n6088 GND.n6087 36.1788
R11592 GND.n6087 GND.n6086 36.1788
R11593 GND.n6086 GND.n460 36.1788
R11594 GND.n6080 GND.n460 36.1788
R11595 GND.n6080 GND.n6079 36.1788
R11596 GND.n6079 GND.n6078 36.1788
R11597 GND.n6078 GND.n468 36.1788
R11598 GND.n4826 GND.n1447 35.817
R11599 GND.n4690 GND.n1565 35.817
R11600 GND.n2320 GND.n2319 32.1338
R11601 GND.n2309 GND.n2308 32.1338
R11602 GND.n2516 GND.n2515 32.1338
R11603 GND.n2534 GND.n2510 32.1338
R11604 GND.n3163 GND.n1346 31.8374
R11605 GND.n4689 GND.n4688 31.8374
R11606 GND.n2586 GND.n2579 30.7517
R11607 GND.n2849 GND.n2848 30.7517
R11608 GND.n2830 GND.n2235 24.6017
R11609 GND.n2375 GND.n2206 24.6017
R11610 GND.n2794 GND.n2198 24.6017
R11611 GND.n2405 GND.n2192 24.6017
R11612 GND.n2780 GND.n2184 24.6017
R11613 GND.n2773 GND.n2177 24.6017
R11614 GND.n2765 GND.n2170 24.6017
R11615 GND.n2758 GND.n2163 24.6017
R11616 GND.n2750 GND.n2155 24.6017
R11617 GND.n2743 GND.n2148 24.6017
R11618 GND.n2735 GND.n2141 24.6017
R11619 GND.n2727 GND.n2126 24.6017
R11620 GND.n2720 GND.n2118 24.6017
R11621 GND.n2706 GND.n2103 24.6017
R11622 GND.n2699 GND.n2097 24.6017
R11623 GND.n2488 GND.n2090 24.6017
R11624 GND.n2332 GND.n2258 23.8782
R11625 GND.n2822 GND.t68 23.8782
R11626 GND.n3975 GND.n2200 23.8782
R11627 GND.n3983 GND.n2190 23.8782
R11628 GND.n2445 GND.n2133 23.8782
R11629 GND.n2729 GND.n2728 23.8782
R11630 GND.t48 GND.n2074 23.8782
R11631 GND.n4110 GND.n2077 23.8782
R11632 GND.n4118 GND.n2067 23.8782
R11633 GND.n5044 GND.n1165 23.1546
R11634 GND.n3528 GND.n1174 23.1546
R11635 GND.n5038 GND.n1177 23.1546
R11636 GND.n3291 GND.n3290 23.1546
R11637 GND.n3612 GND.n3607 23.1546
R11638 GND.n3622 GND.n3283 23.1546
R11639 GND.n3286 GND.n3275 23.1546
R11640 GND.n3631 GND.n3269 23.1546
R11641 GND.n3636 GND.n3272 23.1546
R11642 GND.n3633 GND.n3258 23.1546
R11643 GND.n3646 GND.n3259 23.1546
R11644 GND.n3263 GND.n3250 23.1546
R11645 GND.n3655 GND.n3246 23.1546
R11646 GND.n3661 GND.n3248 23.1546
R11647 GND.n3658 GND.n3235 23.1546
R11648 GND.n3671 GND.n3236 23.1546
R11649 GND.n3680 GND.n3224 23.1546
R11650 GND.n3686 GND.n3226 23.1546
R11651 GND.n3682 GND.n3214 23.1546
R11652 GND.n3694 GND.n3217 23.1546
R11653 GND.n3216 GND.n3078 23.1546
R11654 GND.n3756 GND.n3080 23.1546
R11655 GND.n3752 GND.n3751 23.1546
R11656 GND.n3091 GND.n3085 23.1546
R11657 GND.n3744 GND.n3092 23.1546
R11658 GND.n3738 GND.n3103 23.1546
R11659 GND.n3735 GND.n3734 23.1546
R11660 GND.n3203 GND.n3107 23.1546
R11661 GND.n3727 GND.n3722 23.1546
R11662 GND.n3726 GND.n3060 23.1546
R11663 GND.n3766 GND.n3062 23.1546
R11664 GND.n3065 GND.n3053 23.1546
R11665 GND.n3775 GND.n3048 23.1546
R11666 GND.n3781 GND.n3050 23.1546
R11667 GND.n3791 GND.n3039 23.1546
R11668 GND.n3042 GND.n3031 23.1546
R11669 GND.n3800 GND.n3025 23.1546
R11670 GND.n3805 GND.n3028 23.1546
R11671 GND.n3802 GND.n3014 23.1546
R11672 GND.n3815 GND.n3015 23.1546
R11673 GND.n3019 GND.n3006 23.1546
R11674 GND.n3824 GND.n3002 23.1546
R11675 GND.n3830 GND.n3004 23.1546
R11676 GND.n3827 GND.n2991 23.1546
R11677 GND.n3840 GND.n2992 23.1546
R11678 GND.n3854 GND.n2980 23.1546
R11679 GND.n3858 GND.n2982 23.1546
R11680 GND.n3846 GND.n2973 23.1546
R11681 GND.n3866 GND.n2971 23.1546
R11682 GND.n3869 GND.n1290 23.1546
R11683 GND.n4953 GND.n1292 23.1546
R11684 GND.n4587 GND.n1664 23.1546
R11685 GND.n4584 GND.n1666 23.1546
R11686 GND.n4160 GND.n1671 23.1546
R11687 GND.n4578 GND.n1680 23.1546
R11688 GND.n4168 GND.n1683 23.1546
R11689 GND.n4572 GND.n1691 23.1546
R11690 GND.n4566 GND.n1702 23.1546
R11691 GND.n4183 GND.n1705 23.1546
R11692 GND.n4560 GND.n1712 23.1546
R11693 GND.n4190 GND.n1715 23.1546
R11694 GND.n4554 GND.n1723 23.1546
R11695 GND.n4198 GND.n1726 23.1546
R11696 GND.n4548 GND.n1733 23.1546
R11697 GND.n4205 GND.n1736 23.1546
R11698 GND.n4542 GND.n1744 23.1546
R11699 GND.n4213 GND.n1747 23.1546
R11700 GND.n4536 GND.n1754 23.1546
R11701 GND.n4530 GND.n1765 23.1546
R11702 GND.n4228 GND.n1768 23.1546
R11703 GND.n4524 GND.n1775 23.1546
R11704 GND.n4235 GND.n1778 23.1546
R11705 GND.n4518 GND.n1784 23.1546
R11706 GND.n4247 GND.n1787 23.1546
R11707 GND.n4512 GND.n1794 23.1546
R11708 GND.n4509 GND.n1797 23.1546
R11709 GND.n4508 GND.n1801 23.1546
R11710 GND.n1890 GND.n155 23.1546
R11711 GND.n4500 GND.n4499 23.1546
R11712 GND.n4490 GND.n1893 23.1546
R11713 GND.n6328 GND.n172 23.1546
R11714 GND.n4484 GND.n175 23.1546
R11715 GND.n6322 GND.n184 23.1546
R11716 GND.n4478 GND.n187 23.1546
R11717 GND.n6316 GND.n194 23.1546
R11718 GND.n4472 GND.n197 23.1546
R11719 GND.n4351 GND.n206 23.1546
R11720 GND.n6304 GND.n214 23.1546
R11721 GND.n4357 GND.n217 23.1546
R11722 GND.n6298 GND.n224 23.1546
R11723 GND.n4365 GND.n227 23.1546
R11724 GND.n6292 GND.n235 23.1546
R11725 GND.n4371 GND.n238 23.1546
R11726 GND.n6286 GND.n245 23.1546
R11727 GND.n4380 GND.n248 23.1546
R11728 GND.n6280 GND.n256 23.1546
R11729 GND.n4450 GND.n259 23.1546
R11730 GND.n4444 GND.n268 23.1546
R11731 GND.n6268 GND.n276 23.1546
R11732 GND.n4438 GND.n279 23.1546
R11733 GND.n6262 GND.n286 23.1546
R11734 GND.n6159 GND.n289 23.1546
R11735 GND.n3967 GND.n2208 22.431
R11736 GND.n3991 GND.n2183 22.431
R11737 GND.n2742 GND.n2140 22.431
R11738 GND.n2458 GND.n2127 22.431
R11739 GND.n4102 GND.n2084 22.431
R11740 GND.n1162 GND.n1154 21.7075
R11741 GND.n2996 GND.t44 21.7075
R11742 GND.n4175 GND.t84 21.7075
R11743 GND.n6152 GND.n295 21.7075
R11744 GND.n3887 GND.t106 20.6221
R11745 GND.t54 GND.n2045 20.6221
R11746 GND.n2303 GND.t42 19.8005
R11747 GND.n2303 GND.t126 19.8005
R11748 GND.n2301 GND.t52 19.8005
R11749 GND.n2301 GND.t147 19.8005
R11750 GND.n2300 GND.t69 19.8005
R11751 GND.n2300 GND.t120 19.8005
R11752 GND.n2529 GND.t114 19.8005
R11753 GND.n2529 GND.t49 19.8005
R11754 GND.n2527 GND.t138 19.8005
R11755 GND.n2527 GND.t32 19.8005
R11756 GND.n2526 GND.t129 19.8005
R11757 GND.n2526 GND.t82 19.8005
R11758 GND.n3240 GND.t11 19.5368
R11759 GND.t51 GND.n2249 19.5368
R11760 GND.n2824 GND.n2823 19.5368
R11761 GND.n3951 GND.n2222 19.5368
R11762 GND.n2808 GND.t1 19.5368
R11763 GND.n4007 GND.n2169 19.5368
R11764 GND.n2757 GND.n2154 19.5368
R11765 GND.t9 GND.n2111 19.5368
R11766 GND.n2473 GND.n2112 19.5368
R11767 GND.n6310 GND.t20 19.5368
R11768 GND.n2295 GND.n2294 19.5087
R11769 GND.n2318 GND.n2295 19.5087
R11770 GND.n2316 GND.n2297 19.5087
R11771 GND.n2312 GND.n2297 19.5087
R11772 GND.n2310 GND.n2299 19.5087
R11773 GND.n2520 GND.n2519 19.5087
R11774 GND.n2520 GND.n2511 19.5087
R11775 GND.n2533 GND.n2525 19.5087
R11776 GND.n3877 GND.n2967 19.3944
R11777 GND.n3877 GND.n2957 19.3944
R11778 GND.n3889 GND.n2957 19.3944
R11779 GND.n3889 GND.n2955 19.3944
R11780 GND.n3893 GND.n2955 19.3944
R11781 GND.n3893 GND.n2262 19.3944
R11782 GND.n3905 GND.n2262 19.3944
R11783 GND.n3905 GND.n2260 19.3944
R11784 GND.n3909 GND.n2260 19.3944
R11785 GND.n3909 GND.n2247 19.3944
R11786 GND.n3921 GND.n2247 19.3944
R11787 GND.n3921 GND.n2245 19.3944
R11788 GND.n3925 GND.n2245 19.3944
R11789 GND.n3925 GND.n2233 19.3944
R11790 GND.n3937 GND.n2233 19.3944
R11791 GND.n3937 GND.n2231 19.3944
R11792 GND.n3941 GND.n2231 19.3944
R11793 GND.n3941 GND.n2218 19.3944
R11794 GND.n3953 GND.n2218 19.3944
R11795 GND.n3953 GND.n2216 19.3944
R11796 GND.n3957 GND.n2216 19.3944
R11797 GND.n3957 GND.n2204 19.3944
R11798 GND.n3969 GND.n2204 19.3944
R11799 GND.n3969 GND.n2202 19.3944
R11800 GND.n3973 GND.n2202 19.3944
R11801 GND.n3973 GND.n2188 19.3944
R11802 GND.n3985 GND.n2188 19.3944
R11803 GND.n3985 GND.n2186 19.3944
R11804 GND.n3989 GND.n2186 19.3944
R11805 GND.n3989 GND.n2174 19.3944
R11806 GND.n4001 GND.n2174 19.3944
R11807 GND.n4001 GND.n2172 19.3944
R11808 GND.n4005 GND.n2172 19.3944
R11809 GND.n4005 GND.n2159 19.3944
R11810 GND.n4017 GND.n2159 19.3944
R11811 GND.n4017 GND.n2157 19.3944
R11812 GND.n4021 GND.n2157 19.3944
R11813 GND.n4021 GND.n2145 19.3944
R11814 GND.n4033 GND.n2145 19.3944
R11815 GND.n4033 GND.n2143 19.3944
R11816 GND.n4037 GND.n2143 19.3944
R11817 GND.n4037 GND.n2131 19.3944
R11818 GND.n4049 GND.n2131 19.3944
R11819 GND.n4049 GND.n2129 19.3944
R11820 GND.n4053 GND.n2129 19.3944
R11821 GND.n4053 GND.n2116 19.3944
R11822 GND.n4065 GND.n2116 19.3944
R11823 GND.n4065 GND.n2114 19.3944
R11824 GND.n4069 GND.n2114 19.3944
R11825 GND.n4069 GND.n2101 19.3944
R11826 GND.n4081 GND.n2101 19.3944
R11827 GND.n4081 GND.n2099 19.3944
R11828 GND.n4085 GND.n2099 19.3944
R11829 GND.n4085 GND.n2088 19.3944
R11830 GND.n4096 GND.n2088 19.3944
R11831 GND.n4096 GND.n2086 19.3944
R11832 GND.n4100 GND.n2086 19.3944
R11833 GND.n4100 GND.n2072 19.3944
R11834 GND.n4112 GND.n2072 19.3944
R11835 GND.n4112 GND.n2070 19.3944
R11836 GND.n4116 GND.n2070 19.3944
R11837 GND.n4116 GND.n2058 19.3944
R11838 GND.n4128 GND.n2058 19.3944
R11839 GND.n4128 GND.n2055 19.3944
R11840 GND.n4134 GND.n2055 19.3944
R11841 GND.n4134 GND.n2056 19.3944
R11842 GND.n2056 GND.n2043 19.3944
R11843 GND.n4150 GND.n2043 19.3944
R11844 GND.n4151 GND.n4150 19.3944
R11845 GND.n1959 GND.n1958 19.3944
R11846 GND.n1964 GND.n1959 19.3944
R11847 GND.n1964 GND.n1955 19.3944
R11848 GND.n1968 GND.n1955 19.3944
R11849 GND.n1968 GND.n1953 19.3944
R11850 GND.n1974 GND.n1953 19.3944
R11851 GND.n1974 GND.n1951 19.3944
R11852 GND.n1978 GND.n1951 19.3944
R11853 GND.n1978 GND.n1949 19.3944
R11854 GND.n1984 GND.n1949 19.3944
R11855 GND.n1984 GND.n1943 19.3944
R11856 GND.n1997 GND.n1943 19.3944
R11857 GND.n1997 GND.n1941 19.3944
R11858 GND.n2003 GND.n1941 19.3944
R11859 GND.n2003 GND.n1936 19.3944
R11860 GND.n2016 GND.n1936 19.3944
R11861 GND.n2016 GND.n1934 19.3944
R11862 GND.n2025 GND.n1934 19.3944
R11863 GND.n2035 GND.n1926 19.3944
R11864 GND.n2035 GND.n1924 19.3944
R11865 GND.n2040 GND.n1924 19.3944
R11866 GND.n3491 GND.n1184 19.3944
R11867 GND.n5034 GND.n1184 19.3944
R11868 GND.n5034 GND.n5033 19.3944
R11869 GND.n5033 GND.n5032 19.3944
R11870 GND.n5032 GND.n1187 19.3944
R11871 GND.n5028 GND.n1187 19.3944
R11872 GND.n5028 GND.n5027 19.3944
R11873 GND.n5027 GND.n5026 19.3944
R11874 GND.n5026 GND.n1195 19.3944
R11875 GND.n5022 GND.n1195 19.3944
R11876 GND.n5022 GND.n5021 19.3944
R11877 GND.n5021 GND.n5020 19.3944
R11878 GND.n5020 GND.n1203 19.3944
R11879 GND.n5016 GND.n1203 19.3944
R11880 GND.n5016 GND.n5015 19.3944
R11881 GND.n5015 GND.n5014 19.3944
R11882 GND.n5014 GND.n1211 19.3944
R11883 GND.n5010 GND.n1211 19.3944
R11884 GND.n5010 GND.n5009 19.3944
R11885 GND.n5009 GND.n5008 19.3944
R11886 GND.n5008 GND.n1219 19.3944
R11887 GND.n5004 GND.n1219 19.3944
R11888 GND.n5004 GND.n5003 19.3944
R11889 GND.n5003 GND.n5002 19.3944
R11890 GND.n5002 GND.n1227 19.3944
R11891 GND.n4998 GND.n1227 19.3944
R11892 GND.n4998 GND.n4997 19.3944
R11893 GND.n4997 GND.n4996 19.3944
R11894 GND.n4996 GND.n1235 19.3944
R11895 GND.n4992 GND.n1235 19.3944
R11896 GND.n4992 GND.n4991 19.3944
R11897 GND.n4991 GND.n4990 19.3944
R11898 GND.n4990 GND.n1243 19.3944
R11899 GND.n4986 GND.n1243 19.3944
R11900 GND.n4986 GND.n4985 19.3944
R11901 GND.n4985 GND.n4984 19.3944
R11902 GND.n4984 GND.n1251 19.3944
R11903 GND.n4980 GND.n1251 19.3944
R11904 GND.n4980 GND.n4979 19.3944
R11905 GND.n4979 GND.n4978 19.3944
R11906 GND.n4978 GND.n1259 19.3944
R11907 GND.n4974 GND.n1259 19.3944
R11908 GND.n4974 GND.n4973 19.3944
R11909 GND.n4973 GND.n4972 19.3944
R11910 GND.n4972 GND.n1267 19.3944
R11911 GND.n4968 GND.n1267 19.3944
R11912 GND.n4968 GND.n4967 19.3944
R11913 GND.n4967 GND.n4966 19.3944
R11914 GND.n4966 GND.n1275 19.3944
R11915 GND.n4962 GND.n1275 19.3944
R11916 GND.n4962 GND.n4961 19.3944
R11917 GND.n4961 GND.n4960 19.3944
R11918 GND.n4960 GND.n1283 19.3944
R11919 GND.n4956 GND.n1283 19.3944
R11920 GND.n4956 GND.n4955 19.3944
R11921 GND.n4948 GND.n4947 19.3944
R11922 GND.n4947 GND.n4946 19.3944
R11923 GND.n4946 GND.n1302 19.3944
R11924 GND.n4942 GND.n1302 19.3944
R11925 GND.n4942 GND.n4941 19.3944
R11926 GND.n4941 GND.n4940 19.3944
R11927 GND.n4940 GND.n1307 19.3944
R11928 GND.n4936 GND.n1307 19.3944
R11929 GND.n4936 GND.n4935 19.3944
R11930 GND.n4933 GND.n1316 19.3944
R11931 GND.n4929 GND.n1316 19.3944
R11932 GND.n4929 GND.n4928 19.3944
R11933 GND.n4928 GND.n4927 19.3944
R11934 GND.n4927 GND.n1321 19.3944
R11935 GND.n4923 GND.n1321 19.3944
R11936 GND.n4923 GND.n4922 19.3944
R11937 GND.n4922 GND.n4921 19.3944
R11938 GND.n4921 GND.n1326 19.3944
R11939 GND.n4917 GND.n1326 19.3944
R11940 GND.n4909 GND.n1347 19.3944
R11941 GND.n4909 GND.n1349 19.3944
R11942 GND.n4905 GND.n1349 19.3944
R11943 GND.n4905 GND.n4904 19.3944
R11944 GND.n4904 GND.n4903 19.3944
R11945 GND.n4903 GND.n1357 19.3944
R11946 GND.n4899 GND.n1357 19.3944
R11947 GND.n4899 GND.n4898 19.3944
R11948 GND.n4898 GND.n4897 19.3944
R11949 GND.n4897 GND.n1365 19.3944
R11950 GND.n4893 GND.n1365 19.3944
R11951 GND.n4891 GND.n4890 19.3944
R11952 GND.n4890 GND.n1375 19.3944
R11953 GND.n4886 GND.n1375 19.3944
R11954 GND.n4886 GND.n4885 19.3944
R11955 GND.n4885 GND.n4884 19.3944
R11956 GND.n4884 GND.n1383 19.3944
R11957 GND.n4880 GND.n1383 19.3944
R11958 GND.n4880 GND.n4879 19.3944
R11959 GND.n4879 GND.n4878 19.3944
R11960 GND.n4878 GND.n1391 19.3944
R11961 GND.n4874 GND.n1391 19.3944
R11962 GND.n1988 GND.n1946 19.3944
R11963 GND.n1991 GND.n1988 19.3944
R11964 GND.n1994 GND.n1991 19.3944
R11965 GND.n1994 GND.n1939 19.3944
R11966 GND.n2007 GND.n1939 19.3944
R11967 GND.n2010 GND.n2007 19.3944
R11968 GND.n2013 GND.n2010 19.3944
R11969 GND.n2013 GND.n1931 19.3944
R11970 GND.n2029 GND.n1931 19.3944
R11971 GND.n3530 GND.n3526 19.3944
R11972 GND.n3531 GND.n3530 19.3944
R11973 GND.n3531 GND.n3293 19.3944
R11974 GND.n3535 GND.n3293 19.3944
R11975 GND.n3535 GND.n3280 19.3944
R11976 GND.n3624 GND.n3280 19.3944
R11977 GND.n3624 GND.n3277 19.3944
R11978 GND.n3629 GND.n3277 19.3944
R11979 GND.n3629 GND.n3278 19.3944
R11980 GND.n3278 GND.n3256 19.3944
R11981 GND.n3648 GND.n3256 19.3944
R11982 GND.n3648 GND.n3253 19.3944
R11983 GND.n3653 GND.n3253 19.3944
R11984 GND.n3653 GND.n3254 19.3944
R11985 GND.n3254 GND.n3233 19.3944
R11986 GND.n3673 GND.n3233 19.3944
R11987 GND.n3673 GND.n3230 19.3944
R11988 GND.n3678 GND.n3230 19.3944
R11989 GND.n3678 GND.n3231 19.3944
R11990 GND.n3231 GND.n3211 19.3944
R11991 GND.n3696 GND.n3211 19.3944
R11992 GND.n3696 GND.n3209 19.3944
R11993 GND.n3700 GND.n3209 19.3944
R11994 GND.n3701 GND.n3700 19.3944
R11995 GND.n3704 GND.n3701 19.3944
R11996 GND.n3704 GND.n3207 19.3944
R11997 GND.n3709 GND.n3207 19.3944
R11998 GND.n3710 GND.n3709 19.3944
R11999 GND.n3711 GND.n3710 19.3944
R12000 GND.n3711 GND.n3205 19.3944
R12001 GND.n3715 GND.n3205 19.3944
R12002 GND.n3715 GND.n3058 19.3944
R12003 GND.n3768 GND.n3058 19.3944
R12004 GND.n3768 GND.n3055 19.3944
R12005 GND.n3773 GND.n3055 19.3944
R12006 GND.n3773 GND.n3056 19.3944
R12007 GND.n3056 GND.n3036 19.3944
R12008 GND.n3793 GND.n3036 19.3944
R12009 GND.n3793 GND.n3033 19.3944
R12010 GND.n3798 GND.n3033 19.3944
R12011 GND.n3798 GND.n3034 19.3944
R12012 GND.n3034 GND.n3012 19.3944
R12013 GND.n3817 GND.n3012 19.3944
R12014 GND.n3817 GND.n3009 19.3944
R12015 GND.n3822 GND.n3009 19.3944
R12016 GND.n3822 GND.n3010 19.3944
R12017 GND.n3010 GND.n2989 19.3944
R12018 GND.n3842 GND.n2989 19.3944
R12019 GND.n3842 GND.n2986 19.3944
R12020 GND.n3852 GND.n2986 19.3944
R12021 GND.n3852 GND.n2987 19.3944
R12022 GND.n3848 GND.n2987 19.3944
R12023 GND.n3848 GND.n2969 19.3944
R12024 GND.n3871 GND.n2969 19.3944
R12025 GND.n3872 GND.n3871 19.3944
R12026 GND.n4863 GND.n1407 19.3944
R12027 GND.n4863 GND.n4862 19.3944
R12028 GND.n4862 GND.n1412 19.3944
R12029 GND.n4855 GND.n1412 19.3944
R12030 GND.n4855 GND.n4854 19.3944
R12031 GND.n4854 GND.n1423 19.3944
R12032 GND.n4847 GND.n1423 19.3944
R12033 GND.n4847 GND.n4846 19.3944
R12034 GND.n4846 GND.n1433 19.3944
R12035 GND.n3495 GND.n3307 19.3944
R12036 GND.n3501 GND.n3307 19.3944
R12037 GND.n3501 GND.n3305 19.3944
R12038 GND.n3505 GND.n3305 19.3944
R12039 GND.n3505 GND.n3303 19.3944
R12040 GND.n3511 GND.n3303 19.3944
R12041 GND.n3511 GND.n3301 19.3944
R12042 GND.n3516 GND.n3301 19.3944
R12043 GND.n3516 GND.n3299 19.3944
R12044 GND.n3490 GND.n1180 19.3944
R12045 GND.n5036 GND.n1180 19.3944
R12046 GND.n5036 GND.n1181 19.3944
R12047 GND.n1188 GND.n1181 19.3944
R12048 GND.n1189 GND.n1188 19.3944
R12049 GND.n1190 GND.n1189 19.3944
R12050 GND.n3273 GND.n1190 19.3944
R12051 GND.n3273 GND.n1196 19.3944
R12052 GND.n1197 GND.n1196 19.3944
R12053 GND.n1198 GND.n1197 19.3944
R12054 GND.n3260 GND.n1198 19.3944
R12055 GND.n3260 GND.n1204 19.3944
R12056 GND.n1205 GND.n1204 19.3944
R12057 GND.n1206 GND.n1205 19.3944
R12058 GND.n3657 GND.n1206 19.3944
R12059 GND.n3657 GND.n1212 19.3944
R12060 GND.n1213 GND.n1212 19.3944
R12061 GND.n1214 GND.n1213 19.3944
R12062 GND.n3684 GND.n1214 19.3944
R12063 GND.n3684 GND.n1220 19.3944
R12064 GND.n1221 GND.n1220 19.3944
R12065 GND.n1222 GND.n1221 19.3944
R12066 GND.n3754 GND.n1222 19.3944
R12067 GND.n3754 GND.n1228 19.3944
R12068 GND.n1229 GND.n1228 19.3944
R12069 GND.n1230 GND.n1229 19.3944
R12070 GND.n3095 GND.n1230 19.3944
R12071 GND.n3095 GND.n1236 19.3944
R12072 GND.n1237 GND.n1236 19.3944
R12073 GND.n1238 GND.n1237 19.3944
R12074 GND.n3723 GND.n1238 19.3944
R12075 GND.n3723 GND.n1244 19.3944
R12076 GND.n1245 GND.n1244 19.3944
R12077 GND.n1246 GND.n1245 19.3944
R12078 GND.n3052 GND.n1246 19.3944
R12079 GND.n3052 GND.n1252 19.3944
R12080 GND.n1253 GND.n1252 19.3944
R12081 GND.n1254 GND.n1253 19.3944
R12082 GND.n3029 GND.n1254 19.3944
R12083 GND.n3029 GND.n1260 19.3944
R12084 GND.n1261 GND.n1260 19.3944
R12085 GND.n1262 GND.n1261 19.3944
R12086 GND.n3016 GND.n1262 19.3944
R12087 GND.n3016 GND.n1268 19.3944
R12088 GND.n1269 GND.n1268 19.3944
R12089 GND.n1270 GND.n1269 19.3944
R12090 GND.n3826 GND.n1270 19.3944
R12091 GND.n3826 GND.n1276 19.3944
R12092 GND.n1277 GND.n1276 19.3944
R12093 GND.n1278 GND.n1277 19.3944
R12094 GND.n3856 GND.n1278 19.3944
R12095 GND.n3856 GND.n1284 19.3944
R12096 GND.n1285 GND.n1284 19.3944
R12097 GND.n1286 GND.n1285 19.3944
R12098 GND.n1293 GND.n1286 19.3944
R12099 GND.n5936 GND.n555 19.3944
R12100 GND.n5936 GND.n551 19.3944
R12101 GND.n5942 GND.n551 19.3944
R12102 GND.n5942 GND.n549 19.3944
R12103 GND.n5946 GND.n549 19.3944
R12104 GND.n5946 GND.n545 19.3944
R12105 GND.n5952 GND.n545 19.3944
R12106 GND.n5952 GND.n543 19.3944
R12107 GND.n5956 GND.n543 19.3944
R12108 GND.n5956 GND.n539 19.3944
R12109 GND.n5962 GND.n539 19.3944
R12110 GND.n5962 GND.n537 19.3944
R12111 GND.n5966 GND.n537 19.3944
R12112 GND.n5966 GND.n533 19.3944
R12113 GND.n5972 GND.n533 19.3944
R12114 GND.n5972 GND.n531 19.3944
R12115 GND.n5976 GND.n531 19.3944
R12116 GND.n5976 GND.n527 19.3944
R12117 GND.n5982 GND.n527 19.3944
R12118 GND.n5982 GND.n525 19.3944
R12119 GND.n5986 GND.n525 19.3944
R12120 GND.n5986 GND.n521 19.3944
R12121 GND.n5992 GND.n521 19.3944
R12122 GND.n5992 GND.n519 19.3944
R12123 GND.n5996 GND.n519 19.3944
R12124 GND.n5996 GND.n515 19.3944
R12125 GND.n6002 GND.n515 19.3944
R12126 GND.n6002 GND.n513 19.3944
R12127 GND.n6006 GND.n513 19.3944
R12128 GND.n6006 GND.n509 19.3944
R12129 GND.n6012 GND.n509 19.3944
R12130 GND.n6012 GND.n507 19.3944
R12131 GND.n6016 GND.n507 19.3944
R12132 GND.n6016 GND.n503 19.3944
R12133 GND.n6022 GND.n503 19.3944
R12134 GND.n6022 GND.n501 19.3944
R12135 GND.n6026 GND.n501 19.3944
R12136 GND.n6026 GND.n497 19.3944
R12137 GND.n6032 GND.n497 19.3944
R12138 GND.n6032 GND.n495 19.3944
R12139 GND.n6036 GND.n495 19.3944
R12140 GND.n6036 GND.n491 19.3944
R12141 GND.n6042 GND.n491 19.3944
R12142 GND.n6042 GND.n489 19.3944
R12143 GND.n6046 GND.n489 19.3944
R12144 GND.n6046 GND.n485 19.3944
R12145 GND.n6052 GND.n485 19.3944
R12146 GND.n6052 GND.n483 19.3944
R12147 GND.n6056 GND.n483 19.3944
R12148 GND.n6056 GND.n479 19.3944
R12149 GND.n6062 GND.n479 19.3944
R12150 GND.n6062 GND.n477 19.3944
R12151 GND.n6066 GND.n477 19.3944
R12152 GND.n6066 GND.n473 19.3944
R12153 GND.n6072 GND.n473 19.3944
R12154 GND.n5246 GND.n969 19.3944
R12155 GND.n5246 GND.n965 19.3944
R12156 GND.n5252 GND.n965 19.3944
R12157 GND.n5252 GND.n963 19.3944
R12158 GND.n5256 GND.n963 19.3944
R12159 GND.n5256 GND.n959 19.3944
R12160 GND.n5262 GND.n959 19.3944
R12161 GND.n5262 GND.n957 19.3944
R12162 GND.n5266 GND.n957 19.3944
R12163 GND.n5266 GND.n953 19.3944
R12164 GND.n5272 GND.n953 19.3944
R12165 GND.n5272 GND.n951 19.3944
R12166 GND.n5276 GND.n951 19.3944
R12167 GND.n5276 GND.n947 19.3944
R12168 GND.n5282 GND.n947 19.3944
R12169 GND.n5282 GND.n945 19.3944
R12170 GND.n5286 GND.n945 19.3944
R12171 GND.n5286 GND.n941 19.3944
R12172 GND.n5292 GND.n941 19.3944
R12173 GND.n5292 GND.n939 19.3944
R12174 GND.n5296 GND.n939 19.3944
R12175 GND.n5296 GND.n935 19.3944
R12176 GND.n5302 GND.n935 19.3944
R12177 GND.n5302 GND.n933 19.3944
R12178 GND.n5306 GND.n933 19.3944
R12179 GND.n5306 GND.n929 19.3944
R12180 GND.n5312 GND.n929 19.3944
R12181 GND.n5312 GND.n927 19.3944
R12182 GND.n5316 GND.n927 19.3944
R12183 GND.n5316 GND.n923 19.3944
R12184 GND.n5322 GND.n923 19.3944
R12185 GND.n5322 GND.n921 19.3944
R12186 GND.n5326 GND.n921 19.3944
R12187 GND.n5326 GND.n917 19.3944
R12188 GND.n5332 GND.n917 19.3944
R12189 GND.n5332 GND.n915 19.3944
R12190 GND.n5336 GND.n915 19.3944
R12191 GND.n5336 GND.n911 19.3944
R12192 GND.n5342 GND.n911 19.3944
R12193 GND.n5342 GND.n909 19.3944
R12194 GND.n5346 GND.n909 19.3944
R12195 GND.n5346 GND.n905 19.3944
R12196 GND.n5352 GND.n905 19.3944
R12197 GND.n5352 GND.n903 19.3944
R12198 GND.n5356 GND.n903 19.3944
R12199 GND.n5356 GND.n899 19.3944
R12200 GND.n5362 GND.n899 19.3944
R12201 GND.n5362 GND.n897 19.3944
R12202 GND.n5366 GND.n897 19.3944
R12203 GND.n5366 GND.n893 19.3944
R12204 GND.n5372 GND.n893 19.3944
R12205 GND.n5372 GND.n891 19.3944
R12206 GND.n5376 GND.n891 19.3944
R12207 GND.n5376 GND.n887 19.3944
R12208 GND.n5382 GND.n887 19.3944
R12209 GND.n5382 GND.n885 19.3944
R12210 GND.n5386 GND.n885 19.3944
R12211 GND.n5386 GND.n881 19.3944
R12212 GND.n5392 GND.n881 19.3944
R12213 GND.n5392 GND.n879 19.3944
R12214 GND.n5396 GND.n879 19.3944
R12215 GND.n5396 GND.n875 19.3944
R12216 GND.n5402 GND.n875 19.3944
R12217 GND.n5402 GND.n873 19.3944
R12218 GND.n5406 GND.n873 19.3944
R12219 GND.n5406 GND.n869 19.3944
R12220 GND.n5412 GND.n869 19.3944
R12221 GND.n5412 GND.n867 19.3944
R12222 GND.n5416 GND.n867 19.3944
R12223 GND.n5416 GND.n863 19.3944
R12224 GND.n5422 GND.n863 19.3944
R12225 GND.n5422 GND.n861 19.3944
R12226 GND.n5426 GND.n861 19.3944
R12227 GND.n5426 GND.n857 19.3944
R12228 GND.n5432 GND.n857 19.3944
R12229 GND.n5432 GND.n855 19.3944
R12230 GND.n5436 GND.n855 19.3944
R12231 GND.n5436 GND.n851 19.3944
R12232 GND.n5442 GND.n851 19.3944
R12233 GND.n5442 GND.n849 19.3944
R12234 GND.n5446 GND.n849 19.3944
R12235 GND.n5446 GND.n845 19.3944
R12236 GND.n5452 GND.n845 19.3944
R12237 GND.n5452 GND.n843 19.3944
R12238 GND.n5456 GND.n843 19.3944
R12239 GND.n5456 GND.n839 19.3944
R12240 GND.n5462 GND.n839 19.3944
R12241 GND.n5462 GND.n837 19.3944
R12242 GND.n5466 GND.n837 19.3944
R12243 GND.n5466 GND.n833 19.3944
R12244 GND.n5472 GND.n833 19.3944
R12245 GND.n5472 GND.n831 19.3944
R12246 GND.n5476 GND.n831 19.3944
R12247 GND.n5476 GND.n827 19.3944
R12248 GND.n5482 GND.n827 19.3944
R12249 GND.n5482 GND.n825 19.3944
R12250 GND.n5486 GND.n825 19.3944
R12251 GND.n5486 GND.n821 19.3944
R12252 GND.n5492 GND.n821 19.3944
R12253 GND.n5492 GND.n819 19.3944
R12254 GND.n5496 GND.n819 19.3944
R12255 GND.n5496 GND.n815 19.3944
R12256 GND.n5502 GND.n815 19.3944
R12257 GND.n5502 GND.n813 19.3944
R12258 GND.n5506 GND.n813 19.3944
R12259 GND.n5506 GND.n809 19.3944
R12260 GND.n5512 GND.n809 19.3944
R12261 GND.n5512 GND.n807 19.3944
R12262 GND.n5516 GND.n807 19.3944
R12263 GND.n5516 GND.n803 19.3944
R12264 GND.n5522 GND.n803 19.3944
R12265 GND.n5522 GND.n801 19.3944
R12266 GND.n5526 GND.n801 19.3944
R12267 GND.n5526 GND.n797 19.3944
R12268 GND.n5532 GND.n797 19.3944
R12269 GND.n5532 GND.n795 19.3944
R12270 GND.n5536 GND.n795 19.3944
R12271 GND.n5536 GND.n791 19.3944
R12272 GND.n5542 GND.n791 19.3944
R12273 GND.n5542 GND.n789 19.3944
R12274 GND.n5546 GND.n789 19.3944
R12275 GND.n5546 GND.n785 19.3944
R12276 GND.n5552 GND.n785 19.3944
R12277 GND.n5552 GND.n783 19.3944
R12278 GND.n5556 GND.n783 19.3944
R12279 GND.n5556 GND.n779 19.3944
R12280 GND.n5562 GND.n779 19.3944
R12281 GND.n5562 GND.n777 19.3944
R12282 GND.n5566 GND.n777 19.3944
R12283 GND.n5566 GND.n773 19.3944
R12284 GND.n5572 GND.n773 19.3944
R12285 GND.n5572 GND.n771 19.3944
R12286 GND.n5576 GND.n771 19.3944
R12287 GND.n5576 GND.n767 19.3944
R12288 GND.n5582 GND.n767 19.3944
R12289 GND.n5582 GND.n765 19.3944
R12290 GND.n5586 GND.n765 19.3944
R12291 GND.n5586 GND.n761 19.3944
R12292 GND.n5592 GND.n761 19.3944
R12293 GND.n5592 GND.n759 19.3944
R12294 GND.n5596 GND.n759 19.3944
R12295 GND.n5596 GND.n755 19.3944
R12296 GND.n5602 GND.n755 19.3944
R12297 GND.n5602 GND.n753 19.3944
R12298 GND.n5606 GND.n753 19.3944
R12299 GND.n5606 GND.n749 19.3944
R12300 GND.n5612 GND.n749 19.3944
R12301 GND.n5612 GND.n747 19.3944
R12302 GND.n5616 GND.n747 19.3944
R12303 GND.n5616 GND.n743 19.3944
R12304 GND.n5622 GND.n743 19.3944
R12305 GND.n5622 GND.n741 19.3944
R12306 GND.n5626 GND.n741 19.3944
R12307 GND.n5626 GND.n737 19.3944
R12308 GND.n5632 GND.n737 19.3944
R12309 GND.n5632 GND.n735 19.3944
R12310 GND.n5636 GND.n735 19.3944
R12311 GND.n5636 GND.n731 19.3944
R12312 GND.n5642 GND.n731 19.3944
R12313 GND.n5642 GND.n729 19.3944
R12314 GND.n5646 GND.n729 19.3944
R12315 GND.n5646 GND.n725 19.3944
R12316 GND.n5652 GND.n725 19.3944
R12317 GND.n5652 GND.n723 19.3944
R12318 GND.n5656 GND.n723 19.3944
R12319 GND.n5656 GND.n719 19.3944
R12320 GND.n5662 GND.n719 19.3944
R12321 GND.n5662 GND.n717 19.3944
R12322 GND.n5666 GND.n717 19.3944
R12323 GND.n5666 GND.n713 19.3944
R12324 GND.n5672 GND.n713 19.3944
R12325 GND.n5672 GND.n711 19.3944
R12326 GND.n5676 GND.n711 19.3944
R12327 GND.n5676 GND.n707 19.3944
R12328 GND.n5682 GND.n707 19.3944
R12329 GND.n5682 GND.n705 19.3944
R12330 GND.n5686 GND.n705 19.3944
R12331 GND.n5686 GND.n701 19.3944
R12332 GND.n5692 GND.n701 19.3944
R12333 GND.n5692 GND.n699 19.3944
R12334 GND.n5696 GND.n699 19.3944
R12335 GND.n5696 GND.n695 19.3944
R12336 GND.n5702 GND.n695 19.3944
R12337 GND.n5702 GND.n693 19.3944
R12338 GND.n5706 GND.n693 19.3944
R12339 GND.n5706 GND.n689 19.3944
R12340 GND.n5712 GND.n689 19.3944
R12341 GND.n5712 GND.n687 19.3944
R12342 GND.n5716 GND.n687 19.3944
R12343 GND.n5716 GND.n683 19.3944
R12344 GND.n5722 GND.n683 19.3944
R12345 GND.n5722 GND.n681 19.3944
R12346 GND.n5726 GND.n681 19.3944
R12347 GND.n5726 GND.n677 19.3944
R12348 GND.n5732 GND.n677 19.3944
R12349 GND.n5732 GND.n675 19.3944
R12350 GND.n5736 GND.n675 19.3944
R12351 GND.n5736 GND.n671 19.3944
R12352 GND.n5742 GND.n671 19.3944
R12353 GND.n5742 GND.n669 19.3944
R12354 GND.n5746 GND.n669 19.3944
R12355 GND.n5746 GND.n665 19.3944
R12356 GND.n5752 GND.n665 19.3944
R12357 GND.n5752 GND.n663 19.3944
R12358 GND.n5756 GND.n663 19.3944
R12359 GND.n5756 GND.n659 19.3944
R12360 GND.n5762 GND.n659 19.3944
R12361 GND.n5762 GND.n657 19.3944
R12362 GND.n5766 GND.n657 19.3944
R12363 GND.n5766 GND.n653 19.3944
R12364 GND.n5772 GND.n653 19.3944
R12365 GND.n5772 GND.n651 19.3944
R12366 GND.n5776 GND.n651 19.3944
R12367 GND.n5776 GND.n647 19.3944
R12368 GND.n5782 GND.n647 19.3944
R12369 GND.n5782 GND.n645 19.3944
R12370 GND.n5786 GND.n645 19.3944
R12371 GND.n5786 GND.n641 19.3944
R12372 GND.n5792 GND.n641 19.3944
R12373 GND.n5792 GND.n639 19.3944
R12374 GND.n5796 GND.n639 19.3944
R12375 GND.n5796 GND.n635 19.3944
R12376 GND.n5802 GND.n635 19.3944
R12377 GND.n5802 GND.n633 19.3944
R12378 GND.n5806 GND.n633 19.3944
R12379 GND.n5806 GND.n629 19.3944
R12380 GND.n5812 GND.n629 19.3944
R12381 GND.n5812 GND.n627 19.3944
R12382 GND.n5816 GND.n627 19.3944
R12383 GND.n5816 GND.n623 19.3944
R12384 GND.n5822 GND.n623 19.3944
R12385 GND.n5822 GND.n621 19.3944
R12386 GND.n5826 GND.n621 19.3944
R12387 GND.n5826 GND.n617 19.3944
R12388 GND.n5832 GND.n617 19.3944
R12389 GND.n5832 GND.n615 19.3944
R12390 GND.n5836 GND.n615 19.3944
R12391 GND.n5836 GND.n611 19.3944
R12392 GND.n5842 GND.n611 19.3944
R12393 GND.n5842 GND.n609 19.3944
R12394 GND.n5846 GND.n609 19.3944
R12395 GND.n5846 GND.n605 19.3944
R12396 GND.n5852 GND.n605 19.3944
R12397 GND.n5852 GND.n603 19.3944
R12398 GND.n5856 GND.n603 19.3944
R12399 GND.n5856 GND.n599 19.3944
R12400 GND.n5862 GND.n599 19.3944
R12401 GND.n5862 GND.n597 19.3944
R12402 GND.n5866 GND.n597 19.3944
R12403 GND.n5866 GND.n593 19.3944
R12404 GND.n5872 GND.n593 19.3944
R12405 GND.n5872 GND.n591 19.3944
R12406 GND.n5876 GND.n591 19.3944
R12407 GND.n5876 GND.n587 19.3944
R12408 GND.n5882 GND.n587 19.3944
R12409 GND.n5882 GND.n585 19.3944
R12410 GND.n5886 GND.n585 19.3944
R12411 GND.n5886 GND.n581 19.3944
R12412 GND.n5892 GND.n581 19.3944
R12413 GND.n5892 GND.n579 19.3944
R12414 GND.n5896 GND.n579 19.3944
R12415 GND.n5896 GND.n575 19.3944
R12416 GND.n5902 GND.n575 19.3944
R12417 GND.n5902 GND.n573 19.3944
R12418 GND.n5906 GND.n573 19.3944
R12419 GND.n5906 GND.n569 19.3944
R12420 GND.n5912 GND.n569 19.3944
R12421 GND.n5912 GND.n567 19.3944
R12422 GND.n5916 GND.n567 19.3944
R12423 GND.n5916 GND.n563 19.3944
R12424 GND.n5922 GND.n563 19.3944
R12425 GND.n5922 GND.n561 19.3944
R12426 GND.n5926 GND.n561 19.3944
R12427 GND.n5926 GND.n557 19.3944
R12428 GND.n5932 GND.n557 19.3944
R12429 GND.n4685 GND.n4684 19.3944
R12430 GND.n4684 GND.n4683 19.3944
R12431 GND.n4683 GND.n4682 19.3944
R12432 GND.n4682 GND.n4680 19.3944
R12433 GND.n4680 GND.n4677 19.3944
R12434 GND.n4677 GND.n4676 19.3944
R12435 GND.n4676 GND.n4673 19.3944
R12436 GND.n4673 GND.n4672 19.3944
R12437 GND.n4672 GND.n4669 19.3944
R12438 GND.n4667 GND.n4665 19.3944
R12439 GND.n4665 GND.n4662 19.3944
R12440 GND.n4662 GND.n4661 19.3944
R12441 GND.n4661 GND.n4658 19.3944
R12442 GND.n4658 GND.n4657 19.3944
R12443 GND.n4657 GND.n4654 19.3944
R12444 GND.n4654 GND.n4653 19.3944
R12445 GND.n4653 GND.n4650 19.3944
R12446 GND.n4650 GND.n4649 19.3944
R12447 GND.n4649 GND.n4646 19.3944
R12448 GND.n4644 GND.n4641 19.3944
R12449 GND.n4641 GND.n4640 19.3944
R12450 GND.n4640 GND.n4637 19.3944
R12451 GND.n4637 GND.n4636 19.3944
R12452 GND.n4636 GND.n4633 19.3944
R12453 GND.n4633 GND.n4632 19.3944
R12454 GND.n4632 GND.n4629 19.3944
R12455 GND.n4629 GND.n4628 19.3944
R12456 GND.n4628 GND.n4625 19.3944
R12457 GND.n4625 GND.n4624 19.3944
R12458 GND.n4624 GND.n4621 19.3944
R12459 GND.n4619 GND.n4616 19.3944
R12460 GND.n4616 GND.n4615 19.3944
R12461 GND.n4615 GND.n4612 19.3944
R12462 GND.n4612 GND.n4611 19.3944
R12463 GND.n4611 GND.n4608 19.3944
R12464 GND.n4608 GND.n4607 19.3944
R12465 GND.n4607 GND.n4604 19.3944
R12466 GND.n4604 GND.n4603 19.3944
R12467 GND.n4603 GND.n4600 19.3944
R12468 GND.n4600 GND.n4599 19.3944
R12469 GND.n4599 GND.n4596 19.3944
R12470 GND.n4589 GND.n1662 19.3944
R12471 GND.n4158 GND.n1662 19.3944
R12472 GND.n4158 GND.n1920 19.3944
R12473 GND.n4170 GND.n1920 19.3944
R12474 GND.n4171 GND.n4170 19.3944
R12475 GND.n4173 GND.n4171 19.3944
R12476 GND.n4173 GND.n1916 19.3944
R12477 GND.n4185 GND.n1916 19.3944
R12478 GND.n4186 GND.n4185 19.3944
R12479 GND.n4188 GND.n4186 19.3944
R12480 GND.n4188 GND.n1912 19.3944
R12481 GND.n4200 GND.n1912 19.3944
R12482 GND.n4201 GND.n4200 19.3944
R12483 GND.n4203 GND.n4201 19.3944
R12484 GND.n4203 GND.n1908 19.3944
R12485 GND.n4215 GND.n1908 19.3944
R12486 GND.n4216 GND.n4215 19.3944
R12487 GND.n4218 GND.n4216 19.3944
R12488 GND.n4218 GND.n1904 19.3944
R12489 GND.n4230 GND.n1904 19.3944
R12490 GND.n4231 GND.n4230 19.3944
R12491 GND.n4233 GND.n4231 19.3944
R12492 GND.n4233 GND.n1900 19.3944
R12493 GND.n4249 GND.n1900 19.3944
R12494 GND.n4250 GND.n4249 19.3944
R12495 GND.n4251 GND.n4250 19.3944
R12496 GND.n4251 GND.n1899 19.3944
R12497 GND.n4258 GND.n1899 19.3944
R12498 GND.n4260 GND.n4258 19.3944
R12499 GND.n4493 GND.n4260 19.3944
R12500 GND.n4493 GND.n4492 19.3944
R12501 GND.n4492 GND.n4261 19.3944
R12502 GND.n4482 GND.n4261 19.3944
R12503 GND.n4482 GND.n4481 19.3944
R12504 GND.n4481 GND.n4480 19.3944
R12505 GND.n4480 GND.n4269 19.3944
R12506 GND.n4344 GND.n4269 19.3944
R12507 GND.n4345 GND.n4344 19.3944
R12508 GND.n4353 GND.n4345 19.3944
R12509 GND.n4354 GND.n4353 19.3944
R12510 GND.n4355 GND.n4354 19.3944
R12511 GND.n4355 GND.n4339 19.3944
R12512 GND.n4367 GND.n4339 19.3944
R12513 GND.n4368 GND.n4367 19.3944
R12514 GND.n4369 GND.n4368 19.3944
R12515 GND.n4369 GND.n4334 19.3944
R12516 GND.n4382 GND.n4334 19.3944
R12517 GND.n4383 GND.n4382 19.3944
R12518 GND.n4384 GND.n4383 19.3944
R12519 GND.n4385 GND.n4384 19.3944
R12520 GND.n4442 GND.n4385 19.3944
R12521 GND.n4442 GND.n4441 19.3944
R12522 GND.n4441 GND.n4440 19.3944
R12523 GND.n4440 GND.n383 19.3944
R12524 GND.n6161 GND.n383 19.3944
R12525 GND.n1669 GND.n1660 19.3944
R12526 GND.n1685 GND.n1669 19.3944
R12527 GND.n4576 GND.n1685 19.3944
R12528 GND.n4576 GND.n4575 19.3944
R12529 GND.n4575 GND.n4574 19.3944
R12530 GND.n4574 GND.n1689 19.3944
R12531 GND.n4564 GND.n1689 19.3944
R12532 GND.n4564 GND.n4563 19.3944
R12533 GND.n4563 GND.n4562 19.3944
R12534 GND.n4562 GND.n1710 19.3944
R12535 GND.n4552 GND.n1710 19.3944
R12536 GND.n4552 GND.n4551 19.3944
R12537 GND.n4551 GND.n4550 19.3944
R12538 GND.n4550 GND.n1731 19.3944
R12539 GND.n4540 GND.n1731 19.3944
R12540 GND.n4540 GND.n4539 19.3944
R12541 GND.n4539 GND.n4538 19.3944
R12542 GND.n4538 GND.n1752 19.3944
R12543 GND.n4528 GND.n1752 19.3944
R12544 GND.n4528 GND.n4527 19.3944
R12545 GND.n4527 GND.n4526 19.3944
R12546 GND.n4526 GND.n1773 19.3944
R12547 GND.n4516 GND.n1773 19.3944
R12548 GND.n4516 GND.n4515 19.3944
R12549 GND.n4515 GND.n4514 19.3944
R12550 GND.n4514 GND.n1792 19.3944
R12551 GND.n4255 GND.n1792 19.3944
R12552 GND.n4256 GND.n4255 19.3944
R12553 GND.n4256 GND.n1895 19.3944
R12554 GND.n4495 GND.n1895 19.3944
R12555 GND.n4495 GND.n178 19.3944
R12556 GND.n6326 GND.n178 19.3944
R12557 GND.n6326 GND.n6325 19.3944
R12558 GND.n6325 GND.n6324 19.3944
R12559 GND.n6324 GND.n182 19.3944
R12560 GND.n6314 GND.n182 19.3944
R12561 GND.n6314 GND.n6313 19.3944
R12562 GND.n6313 GND.n6312 19.3944
R12563 GND.n6312 GND.n202 19.3944
R12564 GND.n6302 GND.n202 19.3944
R12565 GND.n6302 GND.n6301 19.3944
R12566 GND.n6301 GND.n6300 19.3944
R12567 GND.n6300 GND.n222 19.3944
R12568 GND.n6290 GND.n222 19.3944
R12569 GND.n6290 GND.n6289 19.3944
R12570 GND.n6289 GND.n6288 19.3944
R12571 GND.n6288 GND.n243 19.3944
R12572 GND.n6278 GND.n243 19.3944
R12573 GND.n6278 GND.n6277 19.3944
R12574 GND.n6277 GND.n6276 19.3944
R12575 GND.n6276 GND.n264 19.3944
R12576 GND.n6266 GND.n264 19.3944
R12577 GND.n6266 GND.n6265 19.3944
R12578 GND.n6265 GND.n6264 19.3944
R12579 GND.n6264 GND.n284 19.3944
R12580 GND.n6187 GND.n6186 19.3944
R12581 GND.n6186 GND.n360 19.3944
R12582 GND.n6181 GND.n360 19.3944
R12583 GND.n6181 GND.n6180 19.3944
R12584 GND.n6180 GND.n6179 19.3944
R12585 GND.n6179 GND.n367 19.3944
R12586 GND.n6174 GND.n367 19.3944
R12587 GND.n6174 GND.n6173 19.3944
R12588 GND.n6173 GND.n6172 19.3944
R12589 GND.n6172 GND.n374 19.3944
R12590 GND.n6167 GND.n374 19.3944
R12591 GND.n6210 GND.n335 19.3944
R12592 GND.n6210 GND.n340 19.3944
R12593 GND.n6205 GND.n340 19.3944
R12594 GND.n6205 GND.n6204 19.3944
R12595 GND.n6204 GND.n6203 19.3944
R12596 GND.n6203 GND.n346 19.3944
R12597 GND.n6198 GND.n346 19.3944
R12598 GND.n6198 GND.n6197 19.3944
R12599 GND.n6197 GND.n6196 19.3944
R12600 GND.n6196 GND.n353 19.3944
R12601 GND.n6191 GND.n353 19.3944
R12602 GND.n6235 GND.n6234 19.3944
R12603 GND.n6234 GND.n6233 19.3944
R12604 GND.n6233 GND.n318 19.3944
R12605 GND.n6228 GND.n318 19.3944
R12606 GND.n6228 GND.n6227 19.3944
R12607 GND.n6227 GND.n6226 19.3944
R12608 GND.n6226 GND.n325 19.3944
R12609 GND.n6221 GND.n325 19.3944
R12610 GND.n6221 GND.n6220 19.3944
R12611 GND.n6220 GND.n6219 19.3944
R12612 GND.n6219 GND.n332 19.3944
R12613 GND.n6256 GND.n294 19.3944
R12614 GND.n296 GND.n294 19.3944
R12615 GND.n6249 GND.n296 19.3944
R12616 GND.n6249 GND.n6248 19.3944
R12617 GND.n6248 GND.n6247 19.3944
R12618 GND.n6247 GND.n302 19.3944
R12619 GND.n6242 GND.n302 19.3944
R12620 GND.n6242 GND.n6241 19.3944
R12621 GND.n6241 GND.n6240 19.3944
R12622 GND.n4406 GND.n4404 19.3944
R12623 GND.n4406 GND.n4401 19.3944
R12624 GND.n4412 GND.n4401 19.3944
R12625 GND.n4412 GND.n4399 19.3944
R12626 GND.n4416 GND.n4399 19.3944
R12627 GND.n4416 GND.n4397 19.3944
R12628 GND.n4422 GND.n4397 19.3944
R12629 GND.n4422 GND.n4395 19.3944
R12630 GND.n4426 GND.n4395 19.3944
R12631 GND.n4156 GND.n4155 19.3944
R12632 GND.n4162 GND.n4156 19.3944
R12633 GND.n4162 GND.n1921 19.3944
R12634 GND.n4166 GND.n1921 19.3944
R12635 GND.n4166 GND.n1919 19.3944
R12636 GND.n4177 GND.n1919 19.3944
R12637 GND.n4177 GND.n1917 19.3944
R12638 GND.n4181 GND.n1917 19.3944
R12639 GND.n4181 GND.n1915 19.3944
R12640 GND.n4192 GND.n1915 19.3944
R12641 GND.n4192 GND.n1913 19.3944
R12642 GND.n4196 GND.n1913 19.3944
R12643 GND.n4196 GND.n1911 19.3944
R12644 GND.n4207 GND.n1911 19.3944
R12645 GND.n4207 GND.n1909 19.3944
R12646 GND.n4211 GND.n1909 19.3944
R12647 GND.n4211 GND.n1907 19.3944
R12648 GND.n4222 GND.n1907 19.3944
R12649 GND.n4222 GND.n1905 19.3944
R12650 GND.n4226 GND.n1905 19.3944
R12651 GND.n4226 GND.n1903 19.3944
R12652 GND.n4237 GND.n1903 19.3944
R12653 GND.n4237 GND.n1901 19.3944
R12654 GND.n4245 GND.n1901 19.3944
R12655 GND.n4245 GND.n4244 19.3944
R12656 GND.n4244 GND.n4243 19.3944
R12657 GND.n4243 GND.n150 19.3944
R12658 GND.n6337 GND.n150 19.3944
R12659 GND.n6337 GND.n151 19.3944
R12660 GND.n4262 GND.n151 19.3944
R12661 GND.n4488 GND.n4262 19.3944
R12662 GND.n4488 GND.n4487 19.3944
R12663 GND.n4487 GND.n4486 19.3944
R12664 GND.n4486 GND.n4267 19.3944
R12665 GND.n4476 GND.n4267 19.3944
R12666 GND.n4476 GND.n4475 19.3944
R12667 GND.n4475 GND.n4474 19.3944
R12668 GND.n4474 GND.n4274 19.3944
R12669 GND.n4349 GND.n4274 19.3944
R12670 GND.n4349 GND.n4343 19.3944
R12671 GND.n4359 GND.n4343 19.3944
R12672 GND.n4359 GND.n4341 19.3944
R12673 GND.n4363 GND.n4341 19.3944
R12674 GND.n4363 GND.n4338 19.3944
R12675 GND.n4373 GND.n4338 19.3944
R12676 GND.n4373 GND.n4336 19.3944
R12677 GND.n4378 GND.n4336 19.3944
R12678 GND.n4378 GND.n4329 19.3944
R12679 GND.n4448 GND.n4329 19.3944
R12680 GND.n4448 GND.n4447 19.3944
R12681 GND.n4447 GND.n4446 19.3944
R12682 GND.n4446 GND.n4333 19.3944
R12683 GND.n4436 GND.n4333 19.3944
R12684 GND.n4436 GND.n4435 19.3944
R12685 GND.n4435 GND.n4434 19.3944
R12686 GND.n4582 GND.n1673 19.3944
R12687 GND.n4582 GND.n4581 19.3944
R12688 GND.n4581 GND.n4580 19.3944
R12689 GND.n4580 GND.n1678 19.3944
R12690 GND.n4570 GND.n1678 19.3944
R12691 GND.n4570 GND.n4569 19.3944
R12692 GND.n4569 GND.n4568 19.3944
R12693 GND.n4568 GND.n1700 19.3944
R12694 GND.n4558 GND.n1700 19.3944
R12695 GND.n4558 GND.n4557 19.3944
R12696 GND.n4557 GND.n4556 19.3944
R12697 GND.n4556 GND.n1721 19.3944
R12698 GND.n4546 GND.n1721 19.3944
R12699 GND.n4546 GND.n4545 19.3944
R12700 GND.n4545 GND.n4544 19.3944
R12701 GND.n4544 GND.n1742 19.3944
R12702 GND.n4534 GND.n1742 19.3944
R12703 GND.n4534 GND.n4533 19.3944
R12704 GND.n4533 GND.n4532 19.3944
R12705 GND.n4532 GND.n1763 19.3944
R12706 GND.n4522 GND.n1763 19.3944
R12707 GND.n4522 GND.n4521 19.3944
R12708 GND.n4521 GND.n4520 19.3944
R12709 GND.n1782 GND.n166 19.3944
R12710 GND.n1798 GND.n166 19.3944
R12711 GND.n6333 GND.n159 19.3944
R12712 GND.n4497 GND.n160 19.3944
R12713 GND.n6330 GND.n168 19.3944
R12714 GND.n6330 GND.n169 19.3944
R12715 GND.n6320 GND.n169 19.3944
R12716 GND.n6320 GND.n6319 19.3944
R12717 GND.n6319 GND.n6318 19.3944
R12718 GND.n6318 GND.n192 19.3944
R12719 GND.n6308 GND.n192 19.3944
R12720 GND.n6308 GND.n6307 19.3944
R12721 GND.n6307 GND.n6306 19.3944
R12722 GND.n6306 GND.n212 19.3944
R12723 GND.n6296 GND.n212 19.3944
R12724 GND.n6296 GND.n6295 19.3944
R12725 GND.n6295 GND.n6294 19.3944
R12726 GND.n6294 GND.n233 19.3944
R12727 GND.n6284 GND.n233 19.3944
R12728 GND.n6284 GND.n6283 19.3944
R12729 GND.n6283 GND.n6282 19.3944
R12730 GND.n6282 GND.n254 19.3944
R12731 GND.n6272 GND.n254 19.3944
R12732 GND.n6272 GND.n6271 19.3944
R12733 GND.n6271 GND.n6270 19.3944
R12734 GND.n6270 GND.n274 19.3944
R12735 GND.n6260 GND.n274 19.3944
R12736 GND.n6260 GND.n6259 19.3944
R12737 GND.n5128 GND.n1081 19.3944
R12738 GND.n5122 GND.n1081 19.3944
R12739 GND.n5122 GND.n5121 19.3944
R12740 GND.n5121 GND.n5120 19.3944
R12741 GND.n5120 GND.n1088 19.3944
R12742 GND.n5114 GND.n1088 19.3944
R12743 GND.n5114 GND.n5113 19.3944
R12744 GND.n5113 GND.n5112 19.3944
R12745 GND.n5112 GND.n1096 19.3944
R12746 GND.n5106 GND.n1096 19.3944
R12747 GND.n5106 GND.n5105 19.3944
R12748 GND.n5105 GND.n5104 19.3944
R12749 GND.n5104 GND.n1104 19.3944
R12750 GND.n5098 GND.n1104 19.3944
R12751 GND.n5098 GND.n5097 19.3944
R12752 GND.n5097 GND.n5096 19.3944
R12753 GND.n5096 GND.n1112 19.3944
R12754 GND.n5090 GND.n1112 19.3944
R12755 GND.n5090 GND.n5089 19.3944
R12756 GND.n5089 GND.n5088 19.3944
R12757 GND.n5088 GND.n1120 19.3944
R12758 GND.n5082 GND.n1120 19.3944
R12759 GND.n5082 GND.n5081 19.3944
R12760 GND.n5081 GND.n5080 19.3944
R12761 GND.n5080 GND.n1128 19.3944
R12762 GND.n5074 GND.n1128 19.3944
R12763 GND.n5074 GND.n5073 19.3944
R12764 GND.n5073 GND.n5072 19.3944
R12765 GND.n5072 GND.n1136 19.3944
R12766 GND.n5066 GND.n1136 19.3944
R12767 GND.n5066 GND.n5065 19.3944
R12768 GND.n5065 GND.n5064 19.3944
R12769 GND.n5064 GND.n1144 19.3944
R12770 GND.n5058 GND.n1144 19.3944
R12771 GND.n5058 GND.n5057 19.3944
R12772 GND.n5057 GND.n5056 19.3944
R12773 GND.n5056 GND.n1152 19.3944
R12774 GND.n5050 GND.n1152 19.3944
R12775 GND.n5050 GND.n5049 19.3944
R12776 GND.n5049 GND.n5048 19.3944
R12777 GND.n5048 GND.n1160 19.3944
R12778 GND.n3544 GND.n1160 19.3944
R12779 GND.n3544 GND.n3541 19.3944
R12780 GND.n3548 GND.n3541 19.3944
R12781 GND.n3548 GND.n3539 19.3944
R12782 GND.n3605 GND.n3539 19.3944
R12783 GND.n3605 GND.n3604 19.3944
R12784 GND.n3604 GND.n3603 19.3944
R12785 GND.n3603 GND.n3554 19.3944
R12786 GND.n3599 GND.n3554 19.3944
R12787 GND.n3599 GND.n3598 19.3944
R12788 GND.n3598 GND.n3597 19.3944
R12789 GND.n3597 GND.n3560 19.3944
R12790 GND.n3593 GND.n3560 19.3944
R12791 GND.n3593 GND.n3592 19.3944
R12792 GND.n3592 GND.n3591 19.3944
R12793 GND.n3591 GND.n3566 19.3944
R12794 GND.n3587 GND.n3566 19.3944
R12795 GND.n3587 GND.n3586 19.3944
R12796 GND.n3586 GND.n3585 19.3944
R12797 GND.n3585 GND.n3572 19.3944
R12798 GND.n3581 GND.n3572 19.3944
R12799 GND.n3581 GND.n3580 19.3944
R12800 GND.n3580 GND.n3579 19.3944
R12801 GND.n3749 GND.n3088 19.3944
R12802 GND.n3747 GND.n3746 19.3944
R12803 GND.n3111 GND.n3110 19.3944
R12804 GND.n3732 GND.n3731 19.3944
R12805 GND.n3729 GND.n3113 19.3944
R12806 GND.n3200 GND.n3113 19.3944
R12807 GND.n3200 GND.n3199 19.3944
R12808 GND.n3199 GND.n3198 19.3944
R12809 GND.n3198 GND.n3119 19.3944
R12810 GND.n3194 GND.n3119 19.3944
R12811 GND.n3194 GND.n3193 19.3944
R12812 GND.n3193 GND.n3192 19.3944
R12813 GND.n3192 GND.n3125 19.3944
R12814 GND.n3188 GND.n3125 19.3944
R12815 GND.n3188 GND.n3187 19.3944
R12816 GND.n3187 GND.n3186 19.3944
R12817 GND.n3186 GND.n3131 19.3944
R12818 GND.n3182 GND.n3131 19.3944
R12819 GND.n3182 GND.n3181 19.3944
R12820 GND.n3181 GND.n3180 19.3944
R12821 GND.n3180 GND.n3137 19.3944
R12822 GND.n3176 GND.n3137 19.3944
R12823 GND.n3176 GND.n3175 19.3944
R12824 GND.n3175 GND.n3174 19.3944
R12825 GND.n3174 GND.n3143 19.3944
R12826 GND.n3170 GND.n3143 19.3944
R12827 GND.n3170 GND.n3169 19.3944
R12828 GND.n3169 GND.n3168 19.3944
R12829 GND.n3168 GND.n3149 19.3944
R12830 GND.n3162 GND.n3149 19.3944
R12831 GND.n3162 GND.n3161 19.3944
R12832 GND.n3161 GND.n3160 19.3944
R12833 GND.n3160 GND.n3156 19.3944
R12834 GND.n3156 GND.n2964 19.3944
R12835 GND.n3881 GND.n2964 19.3944
R12836 GND.n3881 GND.n2962 19.3944
R12837 GND.n3885 GND.n2962 19.3944
R12838 GND.n3885 GND.n2951 19.3944
R12839 GND.n3897 GND.n2951 19.3944
R12840 GND.n3897 GND.n2949 19.3944
R12841 GND.n3901 GND.n2949 19.3944
R12842 GND.n3901 GND.n2255 19.3944
R12843 GND.n3913 GND.n2255 19.3944
R12844 GND.n3913 GND.n2253 19.3944
R12845 GND.n3917 GND.n2253 19.3944
R12846 GND.n3917 GND.n2240 19.3944
R12847 GND.n3929 GND.n2240 19.3944
R12848 GND.n3929 GND.n2238 19.3944
R12849 GND.n3933 GND.n2238 19.3944
R12850 GND.n3933 GND.n2226 19.3944
R12851 GND.n3945 GND.n2226 19.3944
R12852 GND.n3945 GND.n2224 19.3944
R12853 GND.n3949 GND.n2224 19.3944
R12854 GND.n3949 GND.n2212 19.3944
R12855 GND.n3961 GND.n2212 19.3944
R12856 GND.n3961 GND.n2210 19.3944
R12857 GND.n3965 GND.n2210 19.3944
R12858 GND.n3965 GND.n2196 19.3944
R12859 GND.n3977 GND.n2196 19.3944
R12860 GND.n3977 GND.n2194 19.3944
R12861 GND.n3981 GND.n2194 19.3944
R12862 GND.n3981 GND.n2181 19.3944
R12863 GND.n3993 GND.n2181 19.3944
R12864 GND.n3993 GND.n2179 19.3944
R12865 GND.n3997 GND.n2179 19.3944
R12866 GND.n3997 GND.n2167 19.3944
R12867 GND.n4009 GND.n2167 19.3944
R12868 GND.n4009 GND.n2165 19.3944
R12869 GND.n4013 GND.n2165 19.3944
R12870 GND.n4013 GND.n2152 19.3944
R12871 GND.n4025 GND.n2152 19.3944
R12872 GND.n4025 GND.n2150 19.3944
R12873 GND.n4029 GND.n2150 19.3944
R12874 GND.n4029 GND.n2138 19.3944
R12875 GND.n4041 GND.n2138 19.3944
R12876 GND.n4041 GND.n2136 19.3944
R12877 GND.n4045 GND.n2136 19.3944
R12878 GND.n4045 GND.n2124 19.3944
R12879 GND.n4057 GND.n2124 19.3944
R12880 GND.n4057 GND.n2122 19.3944
R12881 GND.n4061 GND.n2122 19.3944
R12882 GND.n4061 GND.n2109 19.3944
R12883 GND.n4073 GND.n2109 19.3944
R12884 GND.n4073 GND.n2107 19.3944
R12885 GND.n4077 GND.n2107 19.3944
R12886 GND.n4077 GND.n2095 19.3944
R12887 GND.n4089 GND.n2095 19.3944
R12888 GND.n4089 GND.n2093 19.3944
R12889 GND.n4093 GND.n2093 19.3944
R12890 GND.n4093 GND.n2081 19.3944
R12891 GND.n4104 GND.n2081 19.3944
R12892 GND.n4104 GND.n2079 19.3944
R12893 GND.n4108 GND.n2079 19.3944
R12894 GND.n4108 GND.n2065 19.3944
R12895 GND.n4120 GND.n2065 19.3944
R12896 GND.n4120 GND.n2063 19.3944
R12897 GND.n4124 GND.n2063 19.3944
R12898 GND.n4124 GND.n2051 19.3944
R12899 GND.n4138 GND.n2051 19.3944
R12900 GND.n4138 GND.n2049 19.3944
R12901 GND.n4145 GND.n2049 19.3944
R12902 GND.n4145 GND.n4144 19.3944
R12903 GND.n4144 GND.n1559 19.3944
R12904 GND.n4694 GND.n1559 19.3944
R12905 GND.n4694 GND.n4693 19.3944
R12906 GND.n4693 GND.n4692 19.3944
R12907 GND.n4692 GND.n1563 19.3944
R12908 GND.n1832 GND.n1563 19.3944
R12909 GND.n1832 GND.n1829 19.3944
R12910 GND.n1836 GND.n1829 19.3944
R12911 GND.n1836 GND.n1827 19.3944
R12912 GND.n1840 GND.n1827 19.3944
R12913 GND.n1840 GND.n1825 19.3944
R12914 GND.n1844 GND.n1825 19.3944
R12915 GND.n1844 GND.n1823 19.3944
R12916 GND.n1848 GND.n1823 19.3944
R12917 GND.n1848 GND.n1821 19.3944
R12918 GND.n1852 GND.n1821 19.3944
R12919 GND.n1852 GND.n1819 19.3944
R12920 GND.n1856 GND.n1819 19.3944
R12921 GND.n1856 GND.n1817 19.3944
R12922 GND.n1860 GND.n1817 19.3944
R12923 GND.n1860 GND.n1815 19.3944
R12924 GND.n1864 GND.n1815 19.3944
R12925 GND.n1864 GND.n1813 19.3944
R12926 GND.n1868 GND.n1813 19.3944
R12927 GND.n1868 GND.n1811 19.3944
R12928 GND.n1872 GND.n1811 19.3944
R12929 GND.n1872 GND.n1809 19.3944
R12930 GND.n1877 GND.n1809 19.3944
R12931 GND.n1877 GND.n1807 19.3944
R12932 GND.n1881 GND.n1807 19.3944
R12933 GND.n1882 GND.n1881 19.3944
R12934 GND.n1886 GND.n1885 19.3944
R12935 GND.n4506 GND.n4505 19.3944
R12936 GND.n4503 GND.n1888 19.3944
R12937 GND.n4285 GND.n4283 19.3944
R12938 GND.n4289 GND.n4287 19.3944
R12939 GND.n4289 GND.n4280 19.3944
R12940 GND.n4293 GND.n4280 19.3944
R12941 GND.n4293 GND.n4278 19.3944
R12942 GND.n4469 GND.n4278 19.3944
R12943 GND.n4469 GND.n4468 19.3944
R12944 GND.n4468 GND.n4467 19.3944
R12945 GND.n4467 GND.n4299 19.3944
R12946 GND.n4463 GND.n4299 19.3944
R12947 GND.n4463 GND.n4462 19.3944
R12948 GND.n4462 GND.n4461 19.3944
R12949 GND.n4461 GND.n4305 19.3944
R12950 GND.n4457 GND.n4305 19.3944
R12951 GND.n4457 GND.n4456 19.3944
R12952 GND.n4456 GND.n4455 19.3944
R12953 GND.n4455 GND.n4311 19.3944
R12954 GND.n4327 GND.n4311 19.3944
R12955 GND.n4327 GND.n4326 19.3944
R12956 GND.n4326 GND.n4325 19.3944
R12957 GND.n4325 GND.n4317 19.3944
R12958 GND.n4321 GND.n4317 19.3944
R12959 GND.n4321 GND.n390 19.3944
R12960 GND.n6156 GND.n390 19.3944
R12961 GND.n6156 GND.n6155 19.3944
R12962 GND.n6155 GND.n6154 19.3944
R12963 GND.n6154 GND.n394 19.3944
R12964 GND.n6148 GND.n394 19.3944
R12965 GND.n6148 GND.n6147 19.3944
R12966 GND.n6147 GND.n6146 19.3944
R12967 GND.n6146 GND.n402 19.3944
R12968 GND.n6140 GND.n402 19.3944
R12969 GND.n6140 GND.n6139 19.3944
R12970 GND.n6139 GND.n6138 19.3944
R12971 GND.n6138 GND.n410 19.3944
R12972 GND.n6132 GND.n410 19.3944
R12973 GND.n6132 GND.n6131 19.3944
R12974 GND.n6131 GND.n6130 19.3944
R12975 GND.n6130 GND.n418 19.3944
R12976 GND.n6124 GND.n418 19.3944
R12977 GND.n6124 GND.n6123 19.3944
R12978 GND.n6123 GND.n6122 19.3944
R12979 GND.n6122 GND.n426 19.3944
R12980 GND.n6116 GND.n426 19.3944
R12981 GND.n6116 GND.n6115 19.3944
R12982 GND.n6115 GND.n6114 19.3944
R12983 GND.n6114 GND.n434 19.3944
R12984 GND.n6108 GND.n434 19.3944
R12985 GND.n6108 GND.n6107 19.3944
R12986 GND.n6107 GND.n6106 19.3944
R12987 GND.n6106 GND.n442 19.3944
R12988 GND.n6100 GND.n442 19.3944
R12989 GND.n6100 GND.n6099 19.3944
R12990 GND.n6099 GND.n6098 19.3944
R12991 GND.n6098 GND.n450 19.3944
R12992 GND.n6092 GND.n450 19.3944
R12993 GND.n6092 GND.n6091 19.3944
R12994 GND.n6091 GND.n6090 19.3944
R12995 GND.n6090 GND.n458 19.3944
R12996 GND.n6084 GND.n458 19.3944
R12997 GND.n6084 GND.n6083 19.3944
R12998 GND.n6083 GND.n6082 19.3944
R12999 GND.n6082 GND.n466 19.3944
R13000 GND.n6076 GND.n466 19.3944
R13001 GND.n6076 GND.n6075 19.3944
R13002 GND.n3364 GND.n3361 19.3944
R13003 GND.n3364 GND.n3359 19.3944
R13004 GND.n3368 GND.n3359 19.3944
R13005 GND.n3368 GND.n3357 19.3944
R13006 GND.n3374 GND.n3357 19.3944
R13007 GND.n3374 GND.n3355 19.3944
R13008 GND.n3378 GND.n3355 19.3944
R13009 GND.n3378 GND.n3353 19.3944
R13010 GND.n3384 GND.n3353 19.3944
R13011 GND.n3388 GND.n3347 19.3944
R13012 GND.n3394 GND.n3347 19.3944
R13013 GND.n3394 GND.n3345 19.3944
R13014 GND.n3398 GND.n3345 19.3944
R13015 GND.n3398 GND.n3343 19.3944
R13016 GND.n3404 GND.n3343 19.3944
R13017 GND.n3404 GND.n3341 19.3944
R13018 GND.n3408 GND.n3341 19.3944
R13019 GND.n3408 GND.n3339 19.3944
R13020 GND.n3414 GND.n3339 19.3944
R13021 GND.n3414 GND.n3337 19.3944
R13022 GND.n3426 GND.n3335 19.3944
R13023 GND.n3426 GND.n3333 19.3944
R13024 GND.n3430 GND.n3333 19.3944
R13025 GND.n3430 GND.n3331 19.3944
R13026 GND.n3436 GND.n3331 19.3944
R13027 GND.n3436 GND.n3329 19.3944
R13028 GND.n3440 GND.n3329 19.3944
R13029 GND.n3440 GND.n3327 19.3944
R13030 GND.n3446 GND.n3327 19.3944
R13031 GND.n3446 GND.n3325 19.3944
R13032 GND.n3453 GND.n3325 19.3944
R13033 GND.n3459 GND.n3323 19.3944
R13034 GND.n3459 GND.n3321 19.3944
R13035 GND.n3463 GND.n3321 19.3944
R13036 GND.n3463 GND.n3319 19.3944
R13037 GND.n3469 GND.n3319 19.3944
R13038 GND.n3469 GND.n3317 19.3944
R13039 GND.n3473 GND.n3317 19.3944
R13040 GND.n3473 GND.n3315 19.3944
R13041 GND.n3479 GND.n3315 19.3944
R13042 GND.n3479 GND.n3313 19.3944
R13043 GND.n3483 GND.n3313 19.3944
R13044 GND.n5042 GND.n5041 19.3944
R13045 GND.n5041 GND.n5040 19.3944
R13046 GND.n5040 GND.n1172 19.3944
R13047 GND.n3614 GND.n1172 19.3944
R13048 GND.n3614 GND.n3288 19.3944
R13049 GND.n3620 GND.n3288 19.3944
R13050 GND.n3620 GND.n3619 19.3944
R13051 GND.n3619 GND.n3267 19.3944
R13052 GND.n3638 GND.n3267 19.3944
R13053 GND.n3638 GND.n3265 19.3944
R13054 GND.n3644 GND.n3265 19.3944
R13055 GND.n3644 GND.n3643 19.3944
R13056 GND.n3643 GND.n3244 19.3944
R13057 GND.n3663 GND.n3244 19.3944
R13058 GND.n3663 GND.n3242 19.3944
R13059 GND.n3669 GND.n3242 19.3944
R13060 GND.n3669 GND.n3668 19.3944
R13061 GND.n3668 GND.n3222 19.3944
R13062 GND.n3688 GND.n3222 19.3944
R13063 GND.n3688 GND.n3220 19.3944
R13064 GND.n3692 GND.n3220 19.3944
R13065 GND.n3692 GND.n3075 19.3944
R13066 GND.n3758 GND.n3075 19.3944
R13067 GND.n3074 GND.n3073 19.3944
R13068 GND.n3098 GND.n3073 19.3944
R13069 GND.n3741 GND.n3740 19.3944
R13070 GND.n3718 GND.n3717 19.3944
R13071 GND.n3720 GND.n3067 19.3944
R13072 GND.n3764 GND.n3067 19.3944
R13073 GND.n3764 GND.n3763 19.3944
R13074 GND.n3763 GND.n3046 19.3944
R13075 GND.n3783 GND.n3046 19.3944
R13076 GND.n3783 GND.n3044 19.3944
R13077 GND.n3789 GND.n3044 19.3944
R13078 GND.n3789 GND.n3788 19.3944
R13079 GND.n3788 GND.n3023 19.3944
R13080 GND.n3807 GND.n3023 19.3944
R13081 GND.n3807 GND.n3021 19.3944
R13082 GND.n3813 GND.n3021 19.3944
R13083 GND.n3813 GND.n3812 19.3944
R13084 GND.n3812 GND.n3000 19.3944
R13085 GND.n3832 GND.n3000 19.3944
R13086 GND.n3832 GND.n2998 19.3944
R13087 GND.n3838 GND.n2998 19.3944
R13088 GND.n3838 GND.n3837 19.3944
R13089 GND.n3837 GND.n2978 19.3944
R13090 GND.n3860 GND.n2978 19.3944
R13091 GND.n3860 GND.n2976 19.3944
R13092 GND.n3864 GND.n2976 19.3944
R13093 GND.n3864 GND.n1297 19.3944
R13094 GND.n4951 GND.n1297 19.3944
R13095 GND.n5242 GND.n971 19.3944
R13096 GND.n5236 GND.n971 19.3944
R13097 GND.n5236 GND.n5235 19.3944
R13098 GND.n5235 GND.n5234 19.3944
R13099 GND.n5234 GND.n978 19.3944
R13100 GND.n5228 GND.n978 19.3944
R13101 GND.n5228 GND.n5227 19.3944
R13102 GND.n5227 GND.n5226 19.3944
R13103 GND.n5226 GND.n986 19.3944
R13104 GND.n5220 GND.n986 19.3944
R13105 GND.n5220 GND.n5219 19.3944
R13106 GND.n5219 GND.n5218 19.3944
R13107 GND.n5218 GND.n994 19.3944
R13108 GND.n5212 GND.n994 19.3944
R13109 GND.n5212 GND.n5211 19.3944
R13110 GND.n5211 GND.n5210 19.3944
R13111 GND.n5210 GND.n1002 19.3944
R13112 GND.n5204 GND.n1002 19.3944
R13113 GND.n5204 GND.n5203 19.3944
R13114 GND.n5203 GND.n5202 19.3944
R13115 GND.n5202 GND.n1010 19.3944
R13116 GND.n5196 GND.n1010 19.3944
R13117 GND.n5196 GND.n5195 19.3944
R13118 GND.n5195 GND.n5194 19.3944
R13119 GND.n5194 GND.n1018 19.3944
R13120 GND.n5188 GND.n1018 19.3944
R13121 GND.n5188 GND.n5187 19.3944
R13122 GND.n5187 GND.n5186 19.3944
R13123 GND.n5186 GND.n1026 19.3944
R13124 GND.n5180 GND.n1026 19.3944
R13125 GND.n5180 GND.n5179 19.3944
R13126 GND.n5179 GND.n5178 19.3944
R13127 GND.n5178 GND.n1034 19.3944
R13128 GND.n5172 GND.n1034 19.3944
R13129 GND.n5172 GND.n5171 19.3944
R13130 GND.n5171 GND.n5170 19.3944
R13131 GND.n5170 GND.n1042 19.3944
R13132 GND.n5164 GND.n1042 19.3944
R13133 GND.n5164 GND.n5163 19.3944
R13134 GND.n5163 GND.n5162 19.3944
R13135 GND.n5162 GND.n1050 19.3944
R13136 GND.n5156 GND.n1050 19.3944
R13137 GND.n5156 GND.n5155 19.3944
R13138 GND.n5155 GND.n5154 19.3944
R13139 GND.n5154 GND.n1058 19.3944
R13140 GND.n5148 GND.n1058 19.3944
R13141 GND.n5148 GND.n5147 19.3944
R13142 GND.n5147 GND.n5146 19.3944
R13143 GND.n5146 GND.n1066 19.3944
R13144 GND.n5140 GND.n1066 19.3944
R13145 GND.n5140 GND.n5139 19.3944
R13146 GND.n5139 GND.n5138 19.3944
R13147 GND.n5138 GND.n1074 19.3944
R13148 GND.n5132 GND.n1074 19.3944
R13149 GND.n5132 GND.n5131 19.3944
R13150 GND.n4802 GND.n4801 19.3944
R13151 GND.n4801 GND.n4800 19.3944
R13152 GND.n4800 GND.n1470 19.3944
R13153 GND.n4796 GND.n1470 19.3944
R13154 GND.n4796 GND.n4795 19.3944
R13155 GND.n4795 GND.n4794 19.3944
R13156 GND.n4794 GND.n1475 19.3944
R13157 GND.n4790 GND.n1475 19.3944
R13158 GND.n4790 GND.n4789 19.3944
R13159 GND.n4789 GND.n4788 19.3944
R13160 GND.n4788 GND.n1480 19.3944
R13161 GND.n4784 GND.n1480 19.3944
R13162 GND.n4784 GND.n4783 19.3944
R13163 GND.n4783 GND.n4782 19.3944
R13164 GND.n4782 GND.n1485 19.3944
R13165 GND.n4778 GND.n1485 19.3944
R13166 GND.n4778 GND.n4777 19.3944
R13167 GND.n4777 GND.n4776 19.3944
R13168 GND.n4776 GND.n1490 19.3944
R13169 GND.n4772 GND.n1490 19.3944
R13170 GND.n4772 GND.n4771 19.3944
R13171 GND.n4771 GND.n4770 19.3944
R13172 GND.n4770 GND.n1495 19.3944
R13173 GND.n4766 GND.n1495 19.3944
R13174 GND.n4766 GND.n4765 19.3944
R13175 GND.n4765 GND.n4764 19.3944
R13176 GND.n4764 GND.n1500 19.3944
R13177 GND.n4760 GND.n1500 19.3944
R13178 GND.n4760 GND.n4759 19.3944
R13179 GND.n4759 GND.n4758 19.3944
R13180 GND.n4758 GND.n1505 19.3944
R13181 GND.n4754 GND.n1505 19.3944
R13182 GND.n4754 GND.n4753 19.3944
R13183 GND.n4753 GND.n4752 19.3944
R13184 GND.n4752 GND.n1510 19.3944
R13185 GND.n4748 GND.n1510 19.3944
R13186 GND.n4748 GND.n4747 19.3944
R13187 GND.n4747 GND.n4746 19.3944
R13188 GND.n4746 GND.n1515 19.3944
R13189 GND.n4742 GND.n1515 19.3944
R13190 GND.n4742 GND.n4741 19.3944
R13191 GND.n4741 GND.n4740 19.3944
R13192 GND.n4740 GND.n1520 19.3944
R13193 GND.n4736 GND.n1520 19.3944
R13194 GND.n4736 GND.n4735 19.3944
R13195 GND.n4735 GND.n4734 19.3944
R13196 GND.n4734 GND.n1525 19.3944
R13197 GND.n4730 GND.n1525 19.3944
R13198 GND.n4730 GND.n4729 19.3944
R13199 GND.n4729 GND.n4728 19.3944
R13200 GND.n4728 GND.n1530 19.3944
R13201 GND.n4724 GND.n1530 19.3944
R13202 GND.n4724 GND.n4723 19.3944
R13203 GND.n4723 GND.n4722 19.3944
R13204 GND.n4722 GND.n1535 19.3944
R13205 GND.n4718 GND.n1535 19.3944
R13206 GND.n4718 GND.n4717 19.3944
R13207 GND.n4717 GND.n4716 19.3944
R13208 GND.n4716 GND.n1540 19.3944
R13209 GND.n4712 GND.n1540 19.3944
R13210 GND.n4712 GND.n4711 19.3944
R13211 GND.n4711 GND.n4710 19.3944
R13212 GND.n4710 GND.n1545 19.3944
R13213 GND.n4706 GND.n1545 19.3944
R13214 GND.n4706 GND.n4705 19.3944
R13215 GND.n4705 GND.n4704 19.3944
R13216 GND.n4704 GND.n1550 19.3944
R13217 GND.n4700 GND.n1550 19.3944
R13218 GND.n4700 GND.n4699 19.3944
R13219 GND.n4839 GND.n1437 19.3944
R13220 GND.n4830 GND.n1437 19.3944
R13221 GND.n4830 GND.n4829 19.3944
R13222 GND.n4823 GND.n1466 19.3944
R13223 GND.n4819 GND.n1466 19.3944
R13224 GND.n4819 GND.n4818 19.3944
R13225 GND.n4818 GND.n4817 19.3944
R13226 GND.n4817 GND.n4808 19.3944
R13227 GND.n4813 GND.n4808 19.3944
R13228 GND.n4813 GND.n4812 19.3944
R13229 GND.n4812 GND.n1402 19.3944
R13230 GND.n4867 GND.n1402 19.3944
R13231 GND.n4867 GND.n4866 19.3944
R13232 GND.n4866 GND.n1405 19.3944
R13233 GND.n4859 GND.n1405 19.3944
R13234 GND.n4859 GND.n4858 19.3944
R13235 GND.n4858 GND.n1416 19.3944
R13236 GND.n4851 GND.n1416 19.3944
R13237 GND.n4851 GND.n4850 19.3944
R13238 GND.n4850 GND.n1427 19.3944
R13239 GND.n4843 GND.n1427 19.3944
R13240 GND.n3903 GND.n2947 18.4514
R13241 GND.n3743 GND.t16 18.0896
R13242 GND.n2290 GND.t131 18.0896
R13243 GND.n3943 GND.n2229 18.0896
R13244 GND.n2359 GND.n2229 18.0896
R13245 GND.n2418 GND.n2161 18.0896
R13246 GND.n4015 GND.n2161 18.0896
R13247 GND.n4079 GND.n2105 18.0896
R13248 GND.n6335 GND.t14 18.0896
R13249 GND.n2335 GND.n2324 17.9517
R13250 GND.n2538 GND.n2507 17.9517
R13251 GND.n2030 GND.n2029 17.8429
R13252 GND.n4836 GND.n1433 17.8429
R13253 GND.n3299 GND.n3298 17.8429
R13254 GND.n4426 GND.n4393 17.8429
R13255 GND.n2947 GND.n2290 17.7278
R13256 GND.n2837 GND.t162 17.7278
R13257 GND.n4118 GND.n2068 17.7278
R13258 GND.n2346 GND.t27 17.3661
R13259 GND.t31 GND.t74 17.3661
R13260 GND.n4935 GND.n4934 16.6793
R13261 GND.n4669 GND.n4668 16.6793
R13262 GND.n6240 GND.n311 16.6793
R13263 GND.n3384 GND.n3351 16.6793
R13264 GND.n3778 GND.t3 16.6425
R13265 GND.n2367 GND.n2222 16.6425
R13266 GND.n2394 GND.t0 16.6425
R13267 GND.n2772 GND.n2169 16.6425
R13268 GND.n4023 GND.n2154 16.6425
R13269 GND.n2433 GND.t8 16.6425
R13270 GND.n4071 GND.n2112 16.6425
R13271 GND.n2693 GND.n2487 16.6425
R13272 GND.n4220 GND.t5 16.6425
R13273 GND.n2319 GND.n2296 16.0672
R13274 GND.n2309 GND.n2298 16.0672
R13275 GND.n2517 GND.n2516 16.0672
R13276 GND.n2523 GND.n2510 16.0672
R13277 GND.t146 GND.n2251 15.9189
R13278 GND.n4874 GND.n4873 15.9035
R13279 GND.n4596 GND.n1658 15.9035
R13280 GND.n6167 GND.n6166 15.9035
R13281 GND.n6214 GND.n335 15.9035
R13282 GND.n3420 GND.n3335 15.9035
R13283 GND.n3483 GND.n3311 15.9035
R13284 GND.n61 GND.n59 15.6496
R13285 GND.n41 GND.n39 15.6496
R13286 GND.n22 GND.n20 15.6496
R13287 GND.n120 GND.n118 15.6496
R13288 GND.n100 GND.n98 15.6496
R13289 GND.n81 GND.n79 15.6496
R13290 GND.t106 GND.n2953 15.5572
R13291 GND.n4136 GND.t54 15.5572
R13292 GND.n2515 GND.n2514 15.4533
R13293 GND.n3927 GND.n2243 15.1954
R13294 GND.n2802 GND.n2374 15.1954
R13295 GND.n4063 GND.n2120 15.1954
R13296 GND.n2686 GND.n2685 15.1954
R13297 GND.n5046 GND.n1162 14.4718
R13298 GND.n3609 GND.t34 14.4718
R13299 GND.t119 GND.n2220 14.4718
R13300 GND.n6274 GND.t61 14.4718
R13301 GND.n387 GND.n295 14.4718
R13302 GND.n2306 GND.n2299 14.2723
R13303 GND.n2533 GND.n2532 14.2723
R13304 GND.n3919 GND.n2251 13.7482
R13305 GND.n2381 GND.n2208 13.7482
R13306 GND.n2404 GND.n2183 13.7482
R13307 GND.n4039 GND.n2140 13.7482
R13308 GND.n4055 GND.n2127 13.7482
R13309 GND.n2500 GND.n2084 13.7482
R13310 GND.n2323 GND.n2294 13.1884
R13311 GND.n2318 GND.n2317 13.1884
R13312 GND.n2317 GND.n2316 13.1884
R13313 GND.n2312 GND.n2311 13.1884
R13314 GND.n2311 GND.n2310 13.1884
R13315 GND.n2518 GND.n2513 13.1884
R13316 GND.n2519 GND.n2518 13.1884
R13317 GND.n2524 GND.n2511 13.1884
R13318 GND.n2525 GND.n2524 13.1884
R13319 GND.n5045 GND.n5044 13.0247
R13320 GND.n3528 GND.n1165 13.0247
R13321 GND.n5038 GND.n1174 13.0247
R13322 GND.n3291 GND.n1177 13.0247
R13323 GND.n3612 GND.n3290 13.0247
R13324 GND.n3609 GND.n3607 13.0247
R13325 GND.n3622 GND.n3282 13.0247
R13326 GND.n3286 GND.n3283 13.0247
R13327 GND.n3631 GND.n3275 13.0247
R13328 GND.n3636 GND.n3269 13.0247
R13329 GND.n3633 GND.n3272 13.0247
R13330 GND.n3646 GND.n3258 13.0247
R13331 GND.n3263 GND.n3259 13.0247
R13332 GND.n3655 GND.n3250 13.0247
R13333 GND.n3661 GND.n3246 13.0247
R13334 GND.n3658 GND.n3248 13.0247
R13335 GND.n3671 GND.n3235 13.0247
R13336 GND.n3240 GND.n3236 13.0247
R13337 GND.n3680 GND.n3228 13.0247
R13338 GND.n3686 GND.n3224 13.0247
R13339 GND.n3682 GND.n3226 13.0247
R13340 GND.n3694 GND.n3214 13.0247
R13341 GND.n3217 GND.n3216 13.0247
R13342 GND.n3756 GND.n3078 13.0247
R13343 GND.n3752 GND.n3080 13.0247
R13344 GND.n3751 GND.n3085 13.0247
R13345 GND.n3092 GND.n3091 13.0247
R13346 GND.n3744 GND.n3743 13.0247
R13347 GND.n3738 GND.n3101 13.0247
R13348 GND.n3735 GND.n3103 13.0247
R13349 GND.n3734 GND.n3107 13.0247
R13350 GND.n3722 GND.n3203 13.0247
R13351 GND.n3727 GND.n3726 13.0247
R13352 GND.n3766 GND.n3060 13.0247
R13353 GND.n3065 GND.n3062 13.0247
R13354 GND.n3775 GND.n3053 13.0247
R13355 GND.n3781 GND.n3048 13.0247
R13356 GND.n3778 GND.n3050 13.0247
R13357 GND.n3791 GND.n3038 13.0247
R13358 GND.n3042 GND.n3039 13.0247
R13359 GND.n3800 GND.n3031 13.0247
R13360 GND.n3805 GND.n3025 13.0247
R13361 GND.n3802 GND.n3028 13.0247
R13362 GND.n3815 GND.n3014 13.0247
R13363 GND.n3019 GND.n3015 13.0247
R13364 GND.n3824 GND.n3006 13.0247
R13365 GND.n3830 GND.n3002 13.0247
R13366 GND.n3827 GND.n3004 13.0247
R13367 GND.n3840 GND.n2991 13.0247
R13368 GND.n2996 GND.n2992 13.0247
R13369 GND.n3854 GND.n2984 13.0247
R13370 GND.n3858 GND.n2980 13.0247
R13371 GND.n3846 GND.n2982 13.0247
R13372 GND.n3866 GND.n2973 13.0247
R13373 GND.n3869 GND.n2971 13.0247
R13374 GND.n4953 GND.n1290 13.0247
R13375 GND.t81 GND.n2060 13.0247
R13376 GND.n4587 GND.n1666 13.0247
R13377 GND.n4584 GND.n1671 13.0247
R13378 GND.n4160 GND.n1680 13.0247
R13379 GND.n4578 GND.n1683 13.0247
R13380 GND.n4168 GND.n1691 13.0247
R13381 GND.n4572 GND.n1694 13.0247
R13382 GND.n4175 GND.n1702 13.0247
R13383 GND.n4566 GND.n1705 13.0247
R13384 GND.n4183 GND.n1712 13.0247
R13385 GND.n4560 GND.n1715 13.0247
R13386 GND.n4190 GND.n1723 13.0247
R13387 GND.n4554 GND.n1726 13.0247
R13388 GND.n4198 GND.n1733 13.0247
R13389 GND.n4548 GND.n1736 13.0247
R13390 GND.n4205 GND.n1744 13.0247
R13391 GND.n4542 GND.n1747 13.0247
R13392 GND.n4213 GND.n1754 13.0247
R13393 GND.n4536 GND.n1757 13.0247
R13394 GND.n4220 GND.n1765 13.0247
R13395 GND.n4530 GND.n1768 13.0247
R13396 GND.n4228 GND.n1775 13.0247
R13397 GND.n4524 GND.n1778 13.0247
R13398 GND.n4235 GND.n1784 13.0247
R13399 GND.n4518 GND.n1787 13.0247
R13400 GND.n4247 GND.n1794 13.0247
R13401 GND.n4512 GND.n1797 13.0247
R13402 GND.n4509 GND.n4508 13.0247
R13403 GND.n1803 GND.n1801 13.0247
R13404 GND.n6335 GND.n155 13.0247
R13405 GND.n4500 GND.n1890 13.0247
R13406 GND.n4499 GND.n1893 13.0247
R13407 GND.n4490 GND.n172 13.0247
R13408 GND.n6328 GND.n175 13.0247
R13409 GND.n4484 GND.n184 13.0247
R13410 GND.n6322 GND.n187 13.0247
R13411 GND.n4478 GND.n194 13.0247
R13412 GND.n6316 GND.n197 13.0247
R13413 GND.n4472 GND.n4471 13.0247
R13414 GND.n6310 GND.n206 13.0247
R13415 GND.n4351 GND.n214 13.0247
R13416 GND.n6304 GND.n217 13.0247
R13417 GND.n4357 GND.n224 13.0247
R13418 GND.n6298 GND.n227 13.0247
R13419 GND.n4365 GND.n235 13.0247
R13420 GND.n6292 GND.n238 13.0247
R13421 GND.n4371 GND.n245 13.0247
R13422 GND.n6286 GND.n248 13.0247
R13423 GND.n4380 GND.n256 13.0247
R13424 GND.n6280 GND.n259 13.0247
R13425 GND.n4451 GND.n4450 13.0247
R13426 GND.n6274 GND.n268 13.0247
R13427 GND.n4444 GND.n276 13.0247
R13428 GND.n6268 GND.n279 13.0247
R13429 GND.n4438 GND.n286 13.0247
R13430 GND.n6262 GND.n289 13.0247
R13431 GND.n6159 GND.n6158 13.0247
R13432 GND.n2944 GND.n2324 12.8005
R13433 GND.n2669 GND.n2538 12.8005
R13434 GND.n62 GND.n58 12.8005
R13435 GND.n42 GND.n38 12.8005
R13436 GND.n23 GND.n19 12.8005
R13437 GND.n121 GND.n117 12.8005
R13438 GND.n101 GND.n97 12.8005
R13439 GND.n82 GND.n78 12.8005
R13440 GND.n3911 GND.n2257 12.3011
R13441 GND.n3911 GND.n2258 12.3011
R13442 GND.n2199 GND.n2190 12.3011
R13443 GND.n4047 GND.n2133 12.3011
R13444 GND.n4087 GND.t137 12.3011
R13445 GND.n2076 GND.n2067 12.3011
R13446 GND.n66 GND.n65 12.0247
R13447 GND.n46 GND.n45 12.0247
R13448 GND.n27 GND.n26 12.0247
R13449 GND.n125 GND.n124 12.0247
R13450 GND.n105 GND.n104 12.0247
R13451 GND.n86 GND.n85 12.0247
R13452 GND.n3959 GND.t164 11.9393
R13453 GND.n2466 GND.t170 11.9393
R13454 GND.n2824 GND.t125 11.5775
R13455 GND.n2480 GND.t58 11.5775
R13456 GND.n2077 GND.t128 11.5775
R13457 GND.n69 GND.n56 11.249
R13458 GND.n49 GND.n36 11.249
R13459 GND.n30 GND.n17 11.249
R13460 GND.n128 GND.n115 11.249
R13461 GND.n108 GND.n95 11.249
R13462 GND.n89 GND.n76 11.249
R13463 GND.n2394 GND.t166 11.2158
R13464 GND.n2433 GND.t160 11.2158
R13465 GND.n3919 GND.n2249 10.854
R13466 GND.n2794 GND.n2381 10.854
R13467 GND.n2405 GND.n2404 10.854
R13468 GND.n4039 GND.n2141 10.854
R13469 GND.n4055 GND.n2126 10.854
R13470 GND.n2677 GND.n2500 10.854
R13471 GND.n2623 GND.n2559 10.6151
R13472 GND.n2623 GND.n2622 10.6151
R13473 GND.n2622 GND.n2621 10.6151
R13474 GND.n2616 GND.n2565 10.6151
R13475 GND.n2616 GND.n2615 10.6151
R13476 GND.n2615 GND.n2614 10.6151
R13477 GND.n2614 GND.n2567 10.6151
R13478 GND.n2609 GND.n2567 10.6151
R13479 GND.n2609 GND.n2608 10.6151
R13480 GND.n2608 GND.n2607 10.6151
R13481 GND.n2607 GND.n2570 10.6151
R13482 GND.n2602 GND.n2570 10.6151
R13483 GND.n2602 GND.n2601 10.6151
R13484 GND.n2601 GND.n2600 10.6151
R13485 GND.n2600 GND.n2573 10.6151
R13486 GND.n2595 GND.n2573 10.6151
R13487 GND.n2595 GND.n2594 10.6151
R13488 GND.n2594 GND.n2593 10.6151
R13489 GND.n2593 GND.n2576 10.6151
R13490 GND.n2588 GND.n2576 10.6151
R13491 GND.n2588 GND.n2587 10.6151
R13492 GND.n2587 GND.n2586 10.6151
R13493 GND.n2848 GND.n2329 10.6151
R13494 GND.n2331 GND.n2329 10.6151
R13495 GND.n2342 GND.n2331 10.6151
R13496 GND.n2343 GND.n2342 10.6151
R13497 GND.n2835 GND.n2343 10.6151
R13498 GND.n2835 GND.n2834 10.6151
R13499 GND.n2834 GND.n2833 10.6151
R13500 GND.n2833 GND.n2344 10.6151
R13501 GND.n2355 GND.n2344 10.6151
R13502 GND.n2356 GND.n2355 10.6151
R13503 GND.n2820 GND.n2356 10.6151
R13504 GND.n2820 GND.n2819 10.6151
R13505 GND.n2819 GND.n2818 10.6151
R13506 GND.n2818 GND.n2357 10.6151
R13507 GND.n2370 GND.n2357 10.6151
R13508 GND.n2371 GND.n2370 10.6151
R13509 GND.n2806 GND.n2371 10.6151
R13510 GND.n2806 GND.n2805 10.6151
R13511 GND.n2805 GND.n2804 10.6151
R13512 GND.n2804 GND.n2372 10.6151
R13513 GND.n2385 GND.n2372 10.6151
R13514 GND.n2386 GND.n2385 10.6151
R13515 GND.n2792 GND.n2386 10.6151
R13516 GND.n2792 GND.n2791 10.6151
R13517 GND.n2791 GND.n2790 10.6151
R13518 GND.n2790 GND.n2387 10.6151
R13519 GND.n2786 GND.n2387 10.6151
R13520 GND.n2786 GND.n2785 10.6151
R13521 GND.n2785 GND.n2784 10.6151
R13522 GND.n2784 GND.n2389 10.6151
R13523 GND.n2391 GND.n2389 10.6151
R13524 GND.n2414 GND.n2391 10.6151
R13525 GND.n2415 GND.n2414 10.6151
R13526 GND.n2770 GND.n2415 10.6151
R13527 GND.n2770 GND.n2769 10.6151
R13528 GND.n2769 GND.n2768 10.6151
R13529 GND.n2768 GND.n2416 10.6151
R13530 GND.n2427 GND.n2416 10.6151
R13531 GND.n2428 GND.n2427 10.6151
R13532 GND.n2755 GND.n2428 10.6151
R13533 GND.n2755 GND.n2754 10.6151
R13534 GND.n2754 GND.n2753 10.6151
R13535 GND.n2753 GND.n2429 10.6151
R13536 GND.n2441 GND.n2429 10.6151
R13537 GND.n2442 GND.n2441 10.6151
R13538 GND.n2740 GND.n2442 10.6151
R13539 GND.n2740 GND.n2739 10.6151
R13540 GND.n2739 GND.n2738 10.6151
R13541 GND.n2738 GND.n2443 10.6151
R13542 GND.n2454 GND.n2443 10.6151
R13543 GND.n2455 GND.n2454 10.6151
R13544 GND.n2725 GND.n2455 10.6151
R13545 GND.n2725 GND.n2724 10.6151
R13546 GND.n2724 GND.n2723 10.6151
R13547 GND.n2723 GND.n2456 10.6151
R13548 GND.n2469 GND.n2456 10.6151
R13549 GND.n2470 GND.n2469 10.6151
R13550 GND.n2711 GND.n2470 10.6151
R13551 GND.n2711 GND.n2710 10.6151
R13552 GND.n2710 GND.n2709 10.6151
R13553 GND.n2709 GND.n2471 10.6151
R13554 GND.n2483 GND.n2471 10.6151
R13555 GND.n2484 GND.n2483 10.6151
R13556 GND.n2697 GND.n2484 10.6151
R13557 GND.n2697 GND.n2696 10.6151
R13558 GND.n2696 GND.n2695 10.6151
R13559 GND.n2695 GND.n2485 10.6151
R13560 GND.n2496 GND.n2485 10.6151
R13561 GND.n2497 GND.n2496 10.6151
R13562 GND.n2682 GND.n2497 10.6151
R13563 GND.n2682 GND.n2681 10.6151
R13564 GND.n2681 GND.n2680 10.6151
R13565 GND.n2680 GND.n2498 10.6151
R13566 GND.n2581 GND.n2498 10.6151
R13567 GND.n2582 GND.n2581 10.6151
R13568 GND.n2582 GND.n2579 10.6151
R13569 GND.n2896 GND.n2893 10.6151
R13570 GND.n2893 GND.n2892 10.6151
R13571 GND.n2892 GND.n2889 10.6151
R13572 GND.n2887 GND.n2884 10.6151
R13573 GND.n2884 GND.n2883 10.6151
R13574 GND.n2883 GND.n2880 10.6151
R13575 GND.n2880 GND.n2879 10.6151
R13576 GND.n2879 GND.n2876 10.6151
R13577 GND.n2876 GND.n2875 10.6151
R13578 GND.n2875 GND.n2872 10.6151
R13579 GND.n2872 GND.n2871 10.6151
R13580 GND.n2871 GND.n2868 10.6151
R13581 GND.n2868 GND.n2867 10.6151
R13582 GND.n2867 GND.n2864 10.6151
R13583 GND.n2864 GND.n2863 10.6151
R13584 GND.n2863 GND.n2860 10.6151
R13585 GND.n2860 GND.n2859 10.6151
R13586 GND.n2859 GND.n2856 10.6151
R13587 GND.n2856 GND.n2855 10.6151
R13588 GND.n2855 GND.n2852 10.6151
R13589 GND.n2852 GND.n2851 10.6151
R13590 GND.n2851 GND.n2849 10.6151
R13591 GND.n2944 GND.n2943 10.6151
R13592 GND.n2943 GND.n2942 10.6151
R13593 GND.n2942 GND.n2941 10.6151
R13594 GND.n2941 GND.n2939 10.6151
R13595 GND.n2939 GND.n2936 10.6151
R13596 GND.n2936 GND.n2935 10.6151
R13597 GND.n2935 GND.n2932 10.6151
R13598 GND.n2932 GND.n2931 10.6151
R13599 GND.n2931 GND.n2928 10.6151
R13600 GND.n2928 GND.n2927 10.6151
R13601 GND.n2927 GND.n2924 10.6151
R13602 GND.n2924 GND.n2923 10.6151
R13603 GND.n2923 GND.n2920 10.6151
R13604 GND.n2920 GND.n2919 10.6151
R13605 GND.n2919 GND.n2916 10.6151
R13606 GND.n2916 GND.n2915 10.6151
R13607 GND.n2915 GND.n2912 10.6151
R13608 GND.n2912 GND.n2911 10.6151
R13609 GND.n2911 GND.n2908 10.6151
R13610 GND.n2906 GND.n2903 10.6151
R13611 GND.n2903 GND.n2902 10.6151
R13612 GND.n2902 GND.n2899 10.6151
R13613 GND.n2669 GND.n2668 10.6151
R13614 GND.n2668 GND.n2667 10.6151
R13615 GND.n2667 GND.n2539 10.6151
R13616 GND.n2662 GND.n2539 10.6151
R13617 GND.n2662 GND.n2661 10.6151
R13618 GND.n2661 GND.n2660 10.6151
R13619 GND.n2660 GND.n2542 10.6151
R13620 GND.n2655 GND.n2542 10.6151
R13621 GND.n2655 GND.n2654 10.6151
R13622 GND.n2654 GND.n2653 10.6151
R13623 GND.n2653 GND.n2545 10.6151
R13624 GND.n2648 GND.n2545 10.6151
R13625 GND.n2648 GND.n2647 10.6151
R13626 GND.n2647 GND.n2646 10.6151
R13627 GND.n2646 GND.n2548 10.6151
R13628 GND.n2641 GND.n2548 10.6151
R13629 GND.n2641 GND.n2640 10.6151
R13630 GND.n2640 GND.n2639 10.6151
R13631 GND.n2639 GND.n2551 10.6151
R13632 GND.n2634 GND.n2633 10.6151
R13633 GND.n2633 GND.n2632 10.6151
R13634 GND.n2632 GND.n2557 10.6151
R13635 GND.n2336 GND.n2335 10.6151
R13636 GND.n2842 GND.n2336 10.6151
R13637 GND.n2842 GND.n2841 10.6151
R13638 GND.n2841 GND.n2840 10.6151
R13639 GND.n2840 GND.n2337 10.6151
R13640 GND.n2349 GND.n2337 10.6151
R13641 GND.n2350 GND.n2349 10.6151
R13642 GND.n2828 GND.n2350 10.6151
R13643 GND.n2828 GND.n2827 10.6151
R13644 GND.n2827 GND.n2826 10.6151
R13645 GND.n2826 GND.n2351 10.6151
R13646 GND.n2363 GND.n2351 10.6151
R13647 GND.n2364 GND.n2363 10.6151
R13648 GND.n2813 GND.n2364 10.6151
R13649 GND.n2813 GND.n2812 10.6151
R13650 GND.n2812 GND.n2811 10.6151
R13651 GND.n2811 GND.n2365 10.6151
R13652 GND.n2377 GND.n2365 10.6151
R13653 GND.n2800 GND.n2377 10.6151
R13654 GND.n2800 GND.n2799 10.6151
R13655 GND.n2799 GND.n2798 10.6151
R13656 GND.n2798 GND.n2378 10.6151
R13657 GND.n2380 GND.n2378 10.6151
R13658 GND.n2398 GND.n2380 10.6151
R13659 GND.n2400 GND.n2398 10.6151
R13660 GND.n2401 GND.n2400 10.6151
R13661 GND.n2402 GND.n2401 10.6151
R13662 GND.n2402 GND.n2396 10.6151
R13663 GND.n2408 GND.n2396 10.6151
R13664 GND.n2409 GND.n2408 10.6151
R13665 GND.n2778 GND.n2409 10.6151
R13666 GND.n2778 GND.n2777 10.6151
R13667 GND.n2777 GND.n2776 10.6151
R13668 GND.n2776 GND.n2410 10.6151
R13669 GND.n2421 GND.n2410 10.6151
R13670 GND.n2422 GND.n2421 10.6151
R13671 GND.n2763 GND.n2422 10.6151
R13672 GND.n2763 GND.n2762 10.6151
R13673 GND.n2762 GND.n2761 10.6151
R13674 GND.n2761 GND.n2423 10.6151
R13675 GND.n2435 GND.n2423 10.6151
R13676 GND.n2436 GND.n2435 10.6151
R13677 GND.n2748 GND.n2436 10.6151
R13678 GND.n2748 GND.n2747 10.6151
R13679 GND.n2747 GND.n2746 10.6151
R13680 GND.n2746 GND.n2437 10.6151
R13681 GND.n2448 GND.n2437 10.6151
R13682 GND.n2449 GND.n2448 10.6151
R13683 GND.n2733 GND.n2449 10.6151
R13684 GND.n2733 GND.n2732 10.6151
R13685 GND.n2732 GND.n2731 10.6151
R13686 GND.n2731 GND.n2450 10.6151
R13687 GND.n2462 GND.n2450 10.6151
R13688 GND.n2463 GND.n2462 10.6151
R13689 GND.n2718 GND.n2463 10.6151
R13690 GND.n2718 GND.n2717 10.6151
R13691 GND.n2717 GND.n2716 10.6151
R13692 GND.n2716 GND.n2464 10.6151
R13693 GND.n2476 GND.n2464 10.6151
R13694 GND.n2477 GND.n2476 10.6151
R13695 GND.n2704 GND.n2477 10.6151
R13696 GND.n2704 GND.n2703 10.6151
R13697 GND.n2703 GND.n2702 10.6151
R13698 GND.n2702 GND.n2478 10.6151
R13699 GND.n2490 GND.n2478 10.6151
R13700 GND.n2691 GND.n2490 10.6151
R13701 GND.n2691 GND.n2690 10.6151
R13702 GND.n2690 GND.n2689 10.6151
R13703 GND.n2689 GND.n2491 10.6151
R13704 GND.n2503 GND.n2491 10.6151
R13705 GND.n2505 GND.n2503 10.6151
R13706 GND.n2506 GND.n2505 10.6151
R13707 GND.n2675 GND.n2506 10.6151
R13708 GND.n2675 GND.n2674 10.6151
R13709 GND.n2674 GND.n2673 10.6151
R13710 GND.n2673 GND.n2507 10.6151
R13711 GND.n1347 GND.n1330 10.4732
R13712 GND.n4645 GND.n4644 10.4732
R13713 GND.n70 GND.n54 10.4732
R13714 GND.n50 GND.n34 10.4732
R13715 GND.n31 GND.n15 10.4732
R13716 GND.n129 GND.n113 10.4732
R13717 GND.n109 GND.n93 10.4732
R13718 GND.n90 GND.n74 10.4732
R13719 GND.n2315 GND.n2296 10.2247
R13720 GND.n2313 GND.n2298 10.2247
R13721 GND.n2517 GND.n2512 10.2247
R13722 GND.n2523 GND.n2522 10.2247
R13723 GND.n2815 GND.t119 10.1304
R13724 GND.t113 GND.n2083 10.1304
R13725 GND.n4873 GND.n4872 10.0853
R13726 GND.n4592 GND.n1658 10.0853
R13727 GND.n6166 GND.n379 10.0853
R13728 GND.n6214 GND.n332 10.0853
R13729 GND.n3420 GND.n3337 10.0853
R13730 GND.n3488 GND.n3311 10.0853
R13731 GND.n72 GND.n71 9.45567
R13732 GND.n52 GND.n51 9.45567
R13733 GND.n33 GND.n32 9.45567
R13734 GND.n131 GND.n130 9.45567
R13735 GND.n111 GND.n110 9.45567
R13736 GND.n92 GND.n91 9.45567
R13737 GND.n3927 GND.n2242 9.40685
R13738 GND.n2375 GND.n2374 9.40685
R13739 GND.n2780 GND.n2392 9.40685
R13740 GND.n4031 GND.n2148 9.40685
R13741 GND.n4063 GND.n2118 9.40685
R13742 GND.n2685 GND.n2684 9.40685
R13743 GND.n2565 GND.n2563 9.36635
R13744 GND.n2888 GND.n2887 9.36635
R13745 GND.n2908 GND.n2907 9.36635
R13746 GND.n2556 GND.n2551 9.36635
R13747 GND.n4934 GND.n4933 9.30959
R13748 GND.n4668 GND.n4667 9.30959
R13749 GND.n6235 GND.n311 9.30959
R13750 GND.n3388 GND.n3351 9.30959
R13751 GND.n5244 GND.n969 9.3005
R13752 GND.n5246 GND.n5245 9.3005
R13753 GND.n965 GND.n964 9.3005
R13754 GND.n5253 GND.n5252 9.3005
R13755 GND.n5254 GND.n963 9.3005
R13756 GND.n5256 GND.n5255 9.3005
R13757 GND.n959 GND.n958 9.3005
R13758 GND.n5263 GND.n5262 9.3005
R13759 GND.n5264 GND.n957 9.3005
R13760 GND.n5266 GND.n5265 9.3005
R13761 GND.n953 GND.n952 9.3005
R13762 GND.n5273 GND.n5272 9.3005
R13763 GND.n5274 GND.n951 9.3005
R13764 GND.n5276 GND.n5275 9.3005
R13765 GND.n947 GND.n946 9.3005
R13766 GND.n5283 GND.n5282 9.3005
R13767 GND.n5284 GND.n945 9.3005
R13768 GND.n5286 GND.n5285 9.3005
R13769 GND.n941 GND.n940 9.3005
R13770 GND.n5293 GND.n5292 9.3005
R13771 GND.n5294 GND.n939 9.3005
R13772 GND.n5296 GND.n5295 9.3005
R13773 GND.n935 GND.n934 9.3005
R13774 GND.n5303 GND.n5302 9.3005
R13775 GND.n5304 GND.n933 9.3005
R13776 GND.n5306 GND.n5305 9.3005
R13777 GND.n929 GND.n928 9.3005
R13778 GND.n5313 GND.n5312 9.3005
R13779 GND.n5314 GND.n927 9.3005
R13780 GND.n5316 GND.n5315 9.3005
R13781 GND.n923 GND.n922 9.3005
R13782 GND.n5323 GND.n5322 9.3005
R13783 GND.n5324 GND.n921 9.3005
R13784 GND.n5326 GND.n5325 9.3005
R13785 GND.n917 GND.n916 9.3005
R13786 GND.n5333 GND.n5332 9.3005
R13787 GND.n5334 GND.n915 9.3005
R13788 GND.n5336 GND.n5335 9.3005
R13789 GND.n911 GND.n910 9.3005
R13790 GND.n5343 GND.n5342 9.3005
R13791 GND.n5344 GND.n909 9.3005
R13792 GND.n5346 GND.n5345 9.3005
R13793 GND.n905 GND.n904 9.3005
R13794 GND.n5353 GND.n5352 9.3005
R13795 GND.n5354 GND.n903 9.3005
R13796 GND.n5356 GND.n5355 9.3005
R13797 GND.n899 GND.n898 9.3005
R13798 GND.n5363 GND.n5362 9.3005
R13799 GND.n5364 GND.n897 9.3005
R13800 GND.n5366 GND.n5365 9.3005
R13801 GND.n893 GND.n892 9.3005
R13802 GND.n5373 GND.n5372 9.3005
R13803 GND.n5374 GND.n891 9.3005
R13804 GND.n5376 GND.n5375 9.3005
R13805 GND.n887 GND.n886 9.3005
R13806 GND.n5383 GND.n5382 9.3005
R13807 GND.n5384 GND.n885 9.3005
R13808 GND.n5386 GND.n5385 9.3005
R13809 GND.n881 GND.n880 9.3005
R13810 GND.n5393 GND.n5392 9.3005
R13811 GND.n5394 GND.n879 9.3005
R13812 GND.n5396 GND.n5395 9.3005
R13813 GND.n875 GND.n874 9.3005
R13814 GND.n5403 GND.n5402 9.3005
R13815 GND.n5404 GND.n873 9.3005
R13816 GND.n5406 GND.n5405 9.3005
R13817 GND.n869 GND.n868 9.3005
R13818 GND.n5413 GND.n5412 9.3005
R13819 GND.n5414 GND.n867 9.3005
R13820 GND.n5416 GND.n5415 9.3005
R13821 GND.n863 GND.n862 9.3005
R13822 GND.n5423 GND.n5422 9.3005
R13823 GND.n5424 GND.n861 9.3005
R13824 GND.n5426 GND.n5425 9.3005
R13825 GND.n857 GND.n856 9.3005
R13826 GND.n5433 GND.n5432 9.3005
R13827 GND.n5434 GND.n855 9.3005
R13828 GND.n5436 GND.n5435 9.3005
R13829 GND.n851 GND.n850 9.3005
R13830 GND.n5443 GND.n5442 9.3005
R13831 GND.n5444 GND.n849 9.3005
R13832 GND.n5446 GND.n5445 9.3005
R13833 GND.n845 GND.n844 9.3005
R13834 GND.n5453 GND.n5452 9.3005
R13835 GND.n5454 GND.n843 9.3005
R13836 GND.n5456 GND.n5455 9.3005
R13837 GND.n839 GND.n838 9.3005
R13838 GND.n5463 GND.n5462 9.3005
R13839 GND.n5464 GND.n837 9.3005
R13840 GND.n5466 GND.n5465 9.3005
R13841 GND.n833 GND.n832 9.3005
R13842 GND.n5473 GND.n5472 9.3005
R13843 GND.n5474 GND.n831 9.3005
R13844 GND.n5476 GND.n5475 9.3005
R13845 GND.n827 GND.n826 9.3005
R13846 GND.n5483 GND.n5482 9.3005
R13847 GND.n5484 GND.n825 9.3005
R13848 GND.n5486 GND.n5485 9.3005
R13849 GND.n821 GND.n820 9.3005
R13850 GND.n5493 GND.n5492 9.3005
R13851 GND.n5494 GND.n819 9.3005
R13852 GND.n5496 GND.n5495 9.3005
R13853 GND.n815 GND.n814 9.3005
R13854 GND.n5503 GND.n5502 9.3005
R13855 GND.n5504 GND.n813 9.3005
R13856 GND.n5506 GND.n5505 9.3005
R13857 GND.n809 GND.n808 9.3005
R13858 GND.n5513 GND.n5512 9.3005
R13859 GND.n5514 GND.n807 9.3005
R13860 GND.n5516 GND.n5515 9.3005
R13861 GND.n803 GND.n802 9.3005
R13862 GND.n5523 GND.n5522 9.3005
R13863 GND.n5524 GND.n801 9.3005
R13864 GND.n5526 GND.n5525 9.3005
R13865 GND.n797 GND.n796 9.3005
R13866 GND.n5533 GND.n5532 9.3005
R13867 GND.n5534 GND.n795 9.3005
R13868 GND.n5536 GND.n5535 9.3005
R13869 GND.n791 GND.n790 9.3005
R13870 GND.n5543 GND.n5542 9.3005
R13871 GND.n5544 GND.n789 9.3005
R13872 GND.n5546 GND.n5545 9.3005
R13873 GND.n785 GND.n784 9.3005
R13874 GND.n5553 GND.n5552 9.3005
R13875 GND.n5554 GND.n783 9.3005
R13876 GND.n5556 GND.n5555 9.3005
R13877 GND.n779 GND.n778 9.3005
R13878 GND.n5563 GND.n5562 9.3005
R13879 GND.n5564 GND.n777 9.3005
R13880 GND.n5566 GND.n5565 9.3005
R13881 GND.n773 GND.n772 9.3005
R13882 GND.n5573 GND.n5572 9.3005
R13883 GND.n5574 GND.n771 9.3005
R13884 GND.n5576 GND.n5575 9.3005
R13885 GND.n767 GND.n766 9.3005
R13886 GND.n5583 GND.n5582 9.3005
R13887 GND.n5584 GND.n765 9.3005
R13888 GND.n5586 GND.n5585 9.3005
R13889 GND.n761 GND.n760 9.3005
R13890 GND.n5593 GND.n5592 9.3005
R13891 GND.n5594 GND.n759 9.3005
R13892 GND.n5596 GND.n5595 9.3005
R13893 GND.n755 GND.n754 9.3005
R13894 GND.n5603 GND.n5602 9.3005
R13895 GND.n5604 GND.n753 9.3005
R13896 GND.n5606 GND.n5605 9.3005
R13897 GND.n749 GND.n748 9.3005
R13898 GND.n5613 GND.n5612 9.3005
R13899 GND.n5614 GND.n747 9.3005
R13900 GND.n5616 GND.n5615 9.3005
R13901 GND.n743 GND.n742 9.3005
R13902 GND.n5623 GND.n5622 9.3005
R13903 GND.n5624 GND.n741 9.3005
R13904 GND.n5626 GND.n5625 9.3005
R13905 GND.n737 GND.n736 9.3005
R13906 GND.n5633 GND.n5632 9.3005
R13907 GND.n5634 GND.n735 9.3005
R13908 GND.n5636 GND.n5635 9.3005
R13909 GND.n731 GND.n730 9.3005
R13910 GND.n5643 GND.n5642 9.3005
R13911 GND.n5644 GND.n729 9.3005
R13912 GND.n5646 GND.n5645 9.3005
R13913 GND.n725 GND.n724 9.3005
R13914 GND.n5653 GND.n5652 9.3005
R13915 GND.n5654 GND.n723 9.3005
R13916 GND.n5656 GND.n5655 9.3005
R13917 GND.n719 GND.n718 9.3005
R13918 GND.n5663 GND.n5662 9.3005
R13919 GND.n5664 GND.n717 9.3005
R13920 GND.n5666 GND.n5665 9.3005
R13921 GND.n713 GND.n712 9.3005
R13922 GND.n5673 GND.n5672 9.3005
R13923 GND.n5674 GND.n711 9.3005
R13924 GND.n5676 GND.n5675 9.3005
R13925 GND.n707 GND.n706 9.3005
R13926 GND.n5683 GND.n5682 9.3005
R13927 GND.n5684 GND.n705 9.3005
R13928 GND.n5686 GND.n5685 9.3005
R13929 GND.n701 GND.n700 9.3005
R13930 GND.n5693 GND.n5692 9.3005
R13931 GND.n5694 GND.n699 9.3005
R13932 GND.n5696 GND.n5695 9.3005
R13933 GND.n695 GND.n694 9.3005
R13934 GND.n5703 GND.n5702 9.3005
R13935 GND.n5704 GND.n693 9.3005
R13936 GND.n5706 GND.n5705 9.3005
R13937 GND.n689 GND.n688 9.3005
R13938 GND.n5713 GND.n5712 9.3005
R13939 GND.n5714 GND.n687 9.3005
R13940 GND.n5716 GND.n5715 9.3005
R13941 GND.n683 GND.n682 9.3005
R13942 GND.n5723 GND.n5722 9.3005
R13943 GND.n5724 GND.n681 9.3005
R13944 GND.n5726 GND.n5725 9.3005
R13945 GND.n677 GND.n676 9.3005
R13946 GND.n5733 GND.n5732 9.3005
R13947 GND.n5734 GND.n675 9.3005
R13948 GND.n5736 GND.n5735 9.3005
R13949 GND.n671 GND.n670 9.3005
R13950 GND.n5743 GND.n5742 9.3005
R13951 GND.n5744 GND.n669 9.3005
R13952 GND.n5746 GND.n5745 9.3005
R13953 GND.n665 GND.n664 9.3005
R13954 GND.n5753 GND.n5752 9.3005
R13955 GND.n5754 GND.n663 9.3005
R13956 GND.n5756 GND.n5755 9.3005
R13957 GND.n659 GND.n658 9.3005
R13958 GND.n5763 GND.n5762 9.3005
R13959 GND.n5764 GND.n657 9.3005
R13960 GND.n5766 GND.n5765 9.3005
R13961 GND.n653 GND.n652 9.3005
R13962 GND.n5773 GND.n5772 9.3005
R13963 GND.n5774 GND.n651 9.3005
R13964 GND.n5776 GND.n5775 9.3005
R13965 GND.n647 GND.n646 9.3005
R13966 GND.n5783 GND.n5782 9.3005
R13967 GND.n5784 GND.n645 9.3005
R13968 GND.n5786 GND.n5785 9.3005
R13969 GND.n641 GND.n640 9.3005
R13970 GND.n5793 GND.n5792 9.3005
R13971 GND.n5794 GND.n639 9.3005
R13972 GND.n5796 GND.n5795 9.3005
R13973 GND.n635 GND.n634 9.3005
R13974 GND.n5803 GND.n5802 9.3005
R13975 GND.n5804 GND.n633 9.3005
R13976 GND.n5806 GND.n5805 9.3005
R13977 GND.n629 GND.n628 9.3005
R13978 GND.n5813 GND.n5812 9.3005
R13979 GND.n5814 GND.n627 9.3005
R13980 GND.n5816 GND.n5815 9.3005
R13981 GND.n623 GND.n622 9.3005
R13982 GND.n5823 GND.n5822 9.3005
R13983 GND.n5824 GND.n621 9.3005
R13984 GND.n5826 GND.n5825 9.3005
R13985 GND.n617 GND.n616 9.3005
R13986 GND.n5833 GND.n5832 9.3005
R13987 GND.n5834 GND.n615 9.3005
R13988 GND.n5836 GND.n5835 9.3005
R13989 GND.n611 GND.n610 9.3005
R13990 GND.n5843 GND.n5842 9.3005
R13991 GND.n5844 GND.n609 9.3005
R13992 GND.n5846 GND.n5845 9.3005
R13993 GND.n605 GND.n604 9.3005
R13994 GND.n5853 GND.n5852 9.3005
R13995 GND.n5854 GND.n603 9.3005
R13996 GND.n5856 GND.n5855 9.3005
R13997 GND.n599 GND.n598 9.3005
R13998 GND.n5863 GND.n5862 9.3005
R13999 GND.n5864 GND.n597 9.3005
R14000 GND.n5866 GND.n5865 9.3005
R14001 GND.n593 GND.n592 9.3005
R14002 GND.n5873 GND.n5872 9.3005
R14003 GND.n5874 GND.n591 9.3005
R14004 GND.n5876 GND.n5875 9.3005
R14005 GND.n587 GND.n586 9.3005
R14006 GND.n5883 GND.n5882 9.3005
R14007 GND.n5884 GND.n585 9.3005
R14008 GND.n5886 GND.n5885 9.3005
R14009 GND.n581 GND.n580 9.3005
R14010 GND.n5893 GND.n5892 9.3005
R14011 GND.n5894 GND.n579 9.3005
R14012 GND.n5896 GND.n5895 9.3005
R14013 GND.n575 GND.n574 9.3005
R14014 GND.n5903 GND.n5902 9.3005
R14015 GND.n5904 GND.n573 9.3005
R14016 GND.n5906 GND.n5905 9.3005
R14017 GND.n569 GND.n568 9.3005
R14018 GND.n5913 GND.n5912 9.3005
R14019 GND.n5914 GND.n567 9.3005
R14020 GND.n5916 GND.n5915 9.3005
R14021 GND.n563 GND.n562 9.3005
R14022 GND.n5923 GND.n5922 9.3005
R14023 GND.n5924 GND.n561 9.3005
R14024 GND.n5926 GND.n5925 9.3005
R14025 GND.n557 GND.n556 9.3005
R14026 GND.n5933 GND.n5932 9.3005
R14027 GND.n5936 GND.n5935 9.3005
R14028 GND.n551 GND.n550 9.3005
R14029 GND.n5943 GND.n5942 9.3005
R14030 GND.n5944 GND.n549 9.3005
R14031 GND.n5946 GND.n5945 9.3005
R14032 GND.n545 GND.n544 9.3005
R14033 GND.n5953 GND.n5952 9.3005
R14034 GND.n5954 GND.n543 9.3005
R14035 GND.n5956 GND.n5955 9.3005
R14036 GND.n539 GND.n538 9.3005
R14037 GND.n5963 GND.n5962 9.3005
R14038 GND.n5964 GND.n537 9.3005
R14039 GND.n5966 GND.n5965 9.3005
R14040 GND.n533 GND.n532 9.3005
R14041 GND.n5973 GND.n5972 9.3005
R14042 GND.n5974 GND.n531 9.3005
R14043 GND.n5976 GND.n5975 9.3005
R14044 GND.n527 GND.n526 9.3005
R14045 GND.n5983 GND.n5982 9.3005
R14046 GND.n5984 GND.n525 9.3005
R14047 GND.n5986 GND.n5985 9.3005
R14048 GND.n521 GND.n520 9.3005
R14049 GND.n5993 GND.n5992 9.3005
R14050 GND.n5994 GND.n519 9.3005
R14051 GND.n5996 GND.n5995 9.3005
R14052 GND.n515 GND.n514 9.3005
R14053 GND.n6003 GND.n6002 9.3005
R14054 GND.n6004 GND.n513 9.3005
R14055 GND.n6006 GND.n6005 9.3005
R14056 GND.n509 GND.n508 9.3005
R14057 GND.n6013 GND.n6012 9.3005
R14058 GND.n6014 GND.n507 9.3005
R14059 GND.n6016 GND.n6015 9.3005
R14060 GND.n503 GND.n502 9.3005
R14061 GND.n6023 GND.n6022 9.3005
R14062 GND.n6024 GND.n501 9.3005
R14063 GND.n6026 GND.n6025 9.3005
R14064 GND.n497 GND.n496 9.3005
R14065 GND.n6033 GND.n6032 9.3005
R14066 GND.n6034 GND.n495 9.3005
R14067 GND.n6036 GND.n6035 9.3005
R14068 GND.n491 GND.n490 9.3005
R14069 GND.n6043 GND.n6042 9.3005
R14070 GND.n6044 GND.n489 9.3005
R14071 GND.n6046 GND.n6045 9.3005
R14072 GND.n485 GND.n484 9.3005
R14073 GND.n6053 GND.n6052 9.3005
R14074 GND.n6054 GND.n483 9.3005
R14075 GND.n6056 GND.n6055 9.3005
R14076 GND.n479 GND.n478 9.3005
R14077 GND.n6063 GND.n6062 9.3005
R14078 GND.n6064 GND.n477 9.3005
R14079 GND.n6066 GND.n6065 9.3005
R14080 GND.n473 GND.n472 9.3005
R14081 GND.n6073 GND.n6072 9.3005
R14082 GND.n5934 GND.n555 9.3005
R14083 GND.n4156 GND.n1922 9.3005
R14084 GND.n4163 GND.n4162 9.3005
R14085 GND.n4164 GND.n1921 9.3005
R14086 GND.n4166 GND.n4165 9.3005
R14087 GND.n1919 GND.n1918 9.3005
R14088 GND.n4178 GND.n4177 9.3005
R14089 GND.n4179 GND.n1917 9.3005
R14090 GND.n4181 GND.n4180 9.3005
R14091 GND.n1915 GND.n1914 9.3005
R14092 GND.n4193 GND.n4192 9.3005
R14093 GND.n4194 GND.n1913 9.3005
R14094 GND.n4196 GND.n4195 9.3005
R14095 GND.n1911 GND.n1910 9.3005
R14096 GND.n4208 GND.n4207 9.3005
R14097 GND.n4209 GND.n1909 9.3005
R14098 GND.n4211 GND.n4210 9.3005
R14099 GND.n1907 GND.n1906 9.3005
R14100 GND.n4223 GND.n4222 9.3005
R14101 GND.n4224 GND.n1905 9.3005
R14102 GND.n4226 GND.n4225 9.3005
R14103 GND.n1903 GND.n1902 9.3005
R14104 GND.n4238 GND.n4237 9.3005
R14105 GND.n4239 GND.n1901 9.3005
R14106 GND.n4245 GND.n4240 9.3005
R14107 GND.n4244 GND.n4241 9.3005
R14108 GND.n4243 GND.n4242 9.3005
R14109 GND.n150 GND.n148 9.3005
R14110 GND.n4155 GND.n4154 9.3005
R14111 GND.n6338 GND.n6337 9.3005
R14112 GND.n151 GND.n149 9.3005
R14113 GND.n4263 GND.n4262 9.3005
R14114 GND.n4488 GND.n4264 9.3005
R14115 GND.n4487 GND.n4265 9.3005
R14116 GND.n4486 GND.n4266 9.3005
R14117 GND.n4270 GND.n4267 9.3005
R14118 GND.n4476 GND.n4271 9.3005
R14119 GND.n4475 GND.n4272 9.3005
R14120 GND.n4474 GND.n4273 9.3005
R14121 GND.n4347 GND.n4274 9.3005
R14122 GND.n4349 GND.n4348 9.3005
R14123 GND.n4343 GND.n4342 9.3005
R14124 GND.n4360 GND.n4359 9.3005
R14125 GND.n4361 GND.n4341 9.3005
R14126 GND.n4363 GND.n4362 9.3005
R14127 GND.n4338 GND.n4337 9.3005
R14128 GND.n4374 GND.n4373 9.3005
R14129 GND.n4375 GND.n4336 9.3005
R14130 GND.n4378 GND.n4377 9.3005
R14131 GND.n4376 GND.n4329 9.3005
R14132 GND.n4448 GND.n4330 9.3005
R14133 GND.n4447 GND.n4331 9.3005
R14134 GND.n4446 GND.n4332 9.3005
R14135 GND.n4387 GND.n4333 9.3005
R14136 GND.n4436 GND.n4388 9.3005
R14137 GND.n4435 GND.n4389 9.3005
R14138 GND.n4434 GND.n4433 9.3005
R14139 GND.n4406 GND.n4405 9.3005
R14140 GND.n4401 GND.n4400 9.3005
R14141 GND.n4413 GND.n4412 9.3005
R14142 GND.n4414 GND.n4399 9.3005
R14143 GND.n4416 GND.n4415 9.3005
R14144 GND.n4397 GND.n4396 9.3005
R14145 GND.n4423 GND.n4422 9.3005
R14146 GND.n4424 GND.n4395 9.3005
R14147 GND.n4426 GND.n4425 9.3005
R14148 GND.n4393 GND.n4390 9.3005
R14149 GND.n4432 GND.n4431 9.3005
R14150 GND.n4404 GND.n382 9.3005
R14151 GND.n294 GND.n293 9.3005
R14152 GND.n298 GND.n296 9.3005
R14153 GND.n6249 GND.n299 9.3005
R14154 GND.n6248 GND.n300 9.3005
R14155 GND.n6247 GND.n301 9.3005
R14156 GND.n305 GND.n302 9.3005
R14157 GND.n6242 GND.n306 9.3005
R14158 GND.n6241 GND.n307 9.3005
R14159 GND.n6240 GND.n308 9.3005
R14160 GND.n314 GND.n311 9.3005
R14161 GND.n6235 GND.n315 9.3005
R14162 GND.n6234 GND.n316 9.3005
R14163 GND.n6233 GND.n317 9.3005
R14164 GND.n321 GND.n318 9.3005
R14165 GND.n6228 GND.n322 9.3005
R14166 GND.n6227 GND.n323 9.3005
R14167 GND.n6226 GND.n324 9.3005
R14168 GND.n328 GND.n325 9.3005
R14169 GND.n6221 GND.n329 9.3005
R14170 GND.n6220 GND.n330 9.3005
R14171 GND.n6219 GND.n331 9.3005
R14172 GND.n338 GND.n332 9.3005
R14173 GND.n6214 GND.n6213 9.3005
R14174 GND.n6212 GND.n335 9.3005
R14175 GND.n6211 GND.n6210 9.3005
R14176 GND.n340 GND.n339 9.3005
R14177 GND.n6205 GND.n343 9.3005
R14178 GND.n6204 GND.n344 9.3005
R14179 GND.n6203 GND.n345 9.3005
R14180 GND.n349 GND.n346 9.3005
R14181 GND.n6198 GND.n350 9.3005
R14182 GND.n6197 GND.n351 9.3005
R14183 GND.n6196 GND.n352 9.3005
R14184 GND.n356 GND.n353 9.3005
R14185 GND.n6191 GND.n357 9.3005
R14186 GND.n6187 GND.n358 9.3005
R14187 GND.n6186 GND.n359 9.3005
R14188 GND.n363 GND.n360 9.3005
R14189 GND.n6181 GND.n364 9.3005
R14190 GND.n6180 GND.n365 9.3005
R14191 GND.n6179 GND.n366 9.3005
R14192 GND.n370 GND.n367 9.3005
R14193 GND.n6174 GND.n371 9.3005
R14194 GND.n6173 GND.n372 9.3005
R14195 GND.n6172 GND.n373 9.3005
R14196 GND.n377 GND.n374 9.3005
R14197 GND.n6167 GND.n378 9.3005
R14198 GND.n6166 GND.n6165 9.3005
R14199 GND.n6164 GND.n379 9.3005
R14200 GND.n6257 GND.n6256 9.3005
R14201 GND.n1669 GND.n1661 9.3005
R14202 GND.n4157 GND.n1685 9.3005
R14203 GND.n4576 GND.n1686 9.3005
R14204 GND.n4575 GND.n1687 9.3005
R14205 GND.n4574 GND.n1688 9.3005
R14206 GND.n4172 GND.n1689 9.3005
R14207 GND.n4564 GND.n1707 9.3005
R14208 GND.n4563 GND.n1708 9.3005
R14209 GND.n4562 GND.n1709 9.3005
R14210 GND.n4187 GND.n1710 9.3005
R14211 GND.n4552 GND.n1728 9.3005
R14212 GND.n4551 GND.n1729 9.3005
R14213 GND.n4550 GND.n1730 9.3005
R14214 GND.n4202 GND.n1731 9.3005
R14215 GND.n4540 GND.n1749 9.3005
R14216 GND.n4539 GND.n1750 9.3005
R14217 GND.n4538 GND.n1751 9.3005
R14218 GND.n4217 GND.n1752 9.3005
R14219 GND.n4528 GND.n1770 9.3005
R14220 GND.n4527 GND.n1771 9.3005
R14221 GND.n4526 GND.n1772 9.3005
R14222 GND.n4232 GND.n1773 9.3005
R14223 GND.n4516 GND.n1789 9.3005
R14224 GND.n4515 GND.n1790 9.3005
R14225 GND.n4514 GND.n1791 9.3005
R14226 GND.n4252 GND.n1792 9.3005
R14227 GND.n4255 GND.n4253 9.3005
R14228 GND.n4257 GND.n4256 9.3005
R14229 GND.n1896 GND.n1895 9.3005
R14230 GND.n4495 GND.n4494 9.3005
R14231 GND.n1897 GND.n178 9.3005
R14232 GND.n6326 GND.n179 9.3005
R14233 GND.n6325 GND.n180 9.3005
R14234 GND.n6324 GND.n181 9.3005
R14235 GND.n4268 GND.n182 9.3005
R14236 GND.n6314 GND.n199 9.3005
R14237 GND.n6313 GND.n200 9.3005
R14238 GND.n6312 GND.n201 9.3005
R14239 GND.n4346 GND.n202 9.3005
R14240 GND.n6302 GND.n219 9.3005
R14241 GND.n6301 GND.n220 9.3005
R14242 GND.n6300 GND.n221 9.3005
R14243 GND.n4340 GND.n222 9.3005
R14244 GND.n6290 GND.n240 9.3005
R14245 GND.n6289 GND.n241 9.3005
R14246 GND.n6288 GND.n242 9.3005
R14247 GND.n4335 GND.n243 9.3005
R14248 GND.n6278 GND.n261 9.3005
R14249 GND.n6277 GND.n262 9.3005
R14250 GND.n6276 GND.n263 9.3005
R14251 GND.n4386 GND.n264 9.3005
R14252 GND.n6266 GND.n281 9.3005
R14253 GND.n6265 GND.n282 9.3005
R14254 GND.n6264 GND.n283 9.3005
R14255 GND.n6162 GND.n284 9.3005
R14256 GND.n4590 GND.n1660 9.3005
R14257 GND.n1662 GND.n1661 9.3005
R14258 GND.n4158 GND.n4157 9.3005
R14259 GND.n1920 GND.n1686 9.3005
R14260 GND.n4170 GND.n1687 9.3005
R14261 GND.n4171 GND.n1688 9.3005
R14262 GND.n4173 GND.n4172 9.3005
R14263 GND.n1916 GND.n1707 9.3005
R14264 GND.n4185 GND.n1708 9.3005
R14265 GND.n4186 GND.n1709 9.3005
R14266 GND.n4188 GND.n4187 9.3005
R14267 GND.n1912 GND.n1728 9.3005
R14268 GND.n4200 GND.n1729 9.3005
R14269 GND.n4201 GND.n1730 9.3005
R14270 GND.n4203 GND.n4202 9.3005
R14271 GND.n1908 GND.n1749 9.3005
R14272 GND.n4215 GND.n1750 9.3005
R14273 GND.n4216 GND.n1751 9.3005
R14274 GND.n4218 GND.n4217 9.3005
R14275 GND.n1904 GND.n1770 9.3005
R14276 GND.n4230 GND.n1771 9.3005
R14277 GND.n4231 GND.n1772 9.3005
R14278 GND.n4233 GND.n4232 9.3005
R14279 GND.n1900 GND.n1789 9.3005
R14280 GND.n4249 GND.n1790 9.3005
R14281 GND.n4250 GND.n1791 9.3005
R14282 GND.n4252 GND.n4251 9.3005
R14283 GND.n4253 GND.n1899 9.3005
R14284 GND.n4258 GND.n4257 9.3005
R14285 GND.n4260 GND.n1896 9.3005
R14286 GND.n4494 GND.n4493 9.3005
R14287 GND.n4492 GND.n1897 9.3005
R14288 GND.n4261 GND.n179 9.3005
R14289 GND.n4482 GND.n180 9.3005
R14290 GND.n4481 GND.n181 9.3005
R14291 GND.n4480 GND.n4268 9.3005
R14292 GND.n4269 GND.n199 9.3005
R14293 GND.n4344 GND.n200 9.3005
R14294 GND.n4345 GND.n201 9.3005
R14295 GND.n4353 GND.n4346 9.3005
R14296 GND.n4354 GND.n219 9.3005
R14297 GND.n4355 GND.n220 9.3005
R14298 GND.n4339 GND.n221 9.3005
R14299 GND.n4367 GND.n4340 9.3005
R14300 GND.n4368 GND.n240 9.3005
R14301 GND.n4369 GND.n241 9.3005
R14302 GND.n4334 GND.n242 9.3005
R14303 GND.n4382 GND.n4335 9.3005
R14304 GND.n4383 GND.n261 9.3005
R14305 GND.n4384 GND.n262 9.3005
R14306 GND.n4385 GND.n263 9.3005
R14307 GND.n4442 GND.n4386 9.3005
R14308 GND.n4441 GND.n281 9.3005
R14309 GND.n4440 GND.n282 9.3005
R14310 GND.n383 GND.n283 9.3005
R14311 GND.n6162 GND.n6161 9.3005
R14312 GND.n4590 GND.n4589 9.3005
R14313 GND.n4596 GND.n4595 9.3005
R14314 GND.n4599 GND.n1654 9.3005
R14315 GND.n4600 GND.n1653 9.3005
R14316 GND.n4603 GND.n1652 9.3005
R14317 GND.n4604 GND.n1651 9.3005
R14318 GND.n4607 GND.n1650 9.3005
R14319 GND.n4608 GND.n1649 9.3005
R14320 GND.n4611 GND.n1648 9.3005
R14321 GND.n4612 GND.n1647 9.3005
R14322 GND.n4615 GND.n1646 9.3005
R14323 GND.n4616 GND.n1645 9.3005
R14324 GND.n4619 GND.n1644 9.3005
R14325 GND.n4621 GND.n1641 9.3005
R14326 GND.n4624 GND.n1640 9.3005
R14327 GND.n4625 GND.n1639 9.3005
R14328 GND.n4628 GND.n1638 9.3005
R14329 GND.n4629 GND.n1637 9.3005
R14330 GND.n4632 GND.n1636 9.3005
R14331 GND.n4633 GND.n1635 9.3005
R14332 GND.n4636 GND.n1634 9.3005
R14333 GND.n4637 GND.n1633 9.3005
R14334 GND.n4640 GND.n1632 9.3005
R14335 GND.n4641 GND.n1631 9.3005
R14336 GND.n4644 GND.n1630 9.3005
R14337 GND.n4646 GND.n1624 9.3005
R14338 GND.n4649 GND.n1623 9.3005
R14339 GND.n4650 GND.n1622 9.3005
R14340 GND.n4653 GND.n1621 9.3005
R14341 GND.n4654 GND.n1620 9.3005
R14342 GND.n4657 GND.n1619 9.3005
R14343 GND.n4658 GND.n1618 9.3005
R14344 GND.n4661 GND.n1617 9.3005
R14345 GND.n4662 GND.n1616 9.3005
R14346 GND.n4665 GND.n1615 9.3005
R14347 GND.n4667 GND.n1614 9.3005
R14348 GND.n4669 GND.n1609 9.3005
R14349 GND.n4672 GND.n1608 9.3005
R14350 GND.n4673 GND.n1607 9.3005
R14351 GND.n4676 GND.n1606 9.3005
R14352 GND.n4677 GND.n1605 9.3005
R14353 GND.n4680 GND.n1604 9.3005
R14354 GND.n4682 GND.n1603 9.3005
R14355 GND.n4683 GND.n1602 9.3005
R14356 GND.n4684 GND.n1601 9.3005
R14357 GND.n4685 GND.n1600 9.3005
R14358 GND.n4668 GND.n1611 9.3005
R14359 GND.n4594 GND.n1658 9.3005
R14360 GND.n4593 GND.n4592 9.3005
R14361 GND.n4582 GND.n1675 9.3005
R14362 GND.n4581 GND.n1676 9.3005
R14363 GND.n4580 GND.n1677 9.3005
R14364 GND.n1696 GND.n1678 9.3005
R14365 GND.n4570 GND.n1697 9.3005
R14366 GND.n4569 GND.n1698 9.3005
R14367 GND.n4568 GND.n1699 9.3005
R14368 GND.n1717 GND.n1700 9.3005
R14369 GND.n4558 GND.n1718 9.3005
R14370 GND.n4557 GND.n1719 9.3005
R14371 GND.n4556 GND.n1720 9.3005
R14372 GND.n1738 GND.n1721 9.3005
R14373 GND.n4546 GND.n1739 9.3005
R14374 GND.n4545 GND.n1740 9.3005
R14375 GND.n4544 GND.n1741 9.3005
R14376 GND.n1759 GND.n1742 9.3005
R14377 GND.n4534 GND.n1760 9.3005
R14378 GND.n4533 GND.n1761 9.3005
R14379 GND.n4532 GND.n1762 9.3005
R14380 GND.n1780 GND.n1763 9.3005
R14381 GND.n4522 GND.n1781 9.3005
R14382 GND.n4521 GND.n162 9.3005
R14383 GND.n169 GND.n161 9.3005
R14384 GND.n6320 GND.n189 9.3005
R14385 GND.n6319 GND.n190 9.3005
R14386 GND.n6318 GND.n191 9.3005
R14387 GND.n208 GND.n192 9.3005
R14388 GND.n6308 GND.n209 9.3005
R14389 GND.n6307 GND.n210 9.3005
R14390 GND.n6306 GND.n211 9.3005
R14391 GND.n229 GND.n212 9.3005
R14392 GND.n6296 GND.n230 9.3005
R14393 GND.n6295 GND.n231 9.3005
R14394 GND.n6294 GND.n232 9.3005
R14395 GND.n250 GND.n233 9.3005
R14396 GND.n6284 GND.n251 9.3005
R14397 GND.n6283 GND.n252 9.3005
R14398 GND.n6282 GND.n253 9.3005
R14399 GND.n270 GND.n254 9.3005
R14400 GND.n6272 GND.n271 9.3005
R14401 GND.n6271 GND.n272 9.3005
R14402 GND.n6270 GND.n273 9.3005
R14403 GND.n291 GND.n274 9.3005
R14404 GND.n6260 GND.n292 9.3005
R14405 GND.n6259 GND.n6258 9.3005
R14406 GND.n1674 GND.n1673 9.3005
R14407 GND.n6331 GND.n166 9.3005
R14408 GND.n6331 GND.n6330 9.3005
R14409 GND.n3115 GND.n3113 9.3005
R14410 GND.n3200 GND.n3116 9.3005
R14411 GND.n3199 GND.n3117 9.3005
R14412 GND.n3198 GND.n3118 9.3005
R14413 GND.n3121 GND.n3119 9.3005
R14414 GND.n3194 GND.n3122 9.3005
R14415 GND.n3193 GND.n3123 9.3005
R14416 GND.n3192 GND.n3124 9.3005
R14417 GND.n3127 GND.n3125 9.3005
R14418 GND.n3188 GND.n3128 9.3005
R14419 GND.n3187 GND.n3129 9.3005
R14420 GND.n3186 GND.n3130 9.3005
R14421 GND.n3133 GND.n3131 9.3005
R14422 GND.n3182 GND.n3134 9.3005
R14423 GND.n3181 GND.n3135 9.3005
R14424 GND.n3180 GND.n3136 9.3005
R14425 GND.n3139 GND.n3137 9.3005
R14426 GND.n3176 GND.n3140 9.3005
R14427 GND.n3175 GND.n3141 9.3005
R14428 GND.n3174 GND.n3142 9.3005
R14429 GND.n3145 GND.n3143 9.3005
R14430 GND.n3170 GND.n3146 9.3005
R14431 GND.n3169 GND.n3147 9.3005
R14432 GND.n3168 GND.n3148 9.3005
R14433 GND.n3151 GND.n3149 9.3005
R14434 GND.n3162 GND.n3152 9.3005
R14435 GND.n3161 GND.n3153 9.3005
R14436 GND.n3160 GND.n3154 9.3005
R14437 GND.n3156 GND.n3155 9.3005
R14438 GND.n2964 GND.n2963 9.3005
R14439 GND.n3882 GND.n3881 9.3005
R14440 GND.n3883 GND.n2962 9.3005
R14441 GND.n3885 GND.n3884 9.3005
R14442 GND.n2951 GND.n2950 9.3005
R14443 GND.n3898 GND.n3897 9.3005
R14444 GND.n3899 GND.n2949 9.3005
R14445 GND.n3901 GND.n3900 9.3005
R14446 GND.n2255 GND.n2254 9.3005
R14447 GND.n3914 GND.n3913 9.3005
R14448 GND.n3915 GND.n2253 9.3005
R14449 GND.n3917 GND.n3916 9.3005
R14450 GND.n2240 GND.n2239 9.3005
R14451 GND.n3930 GND.n3929 9.3005
R14452 GND.n3931 GND.n2238 9.3005
R14453 GND.n3933 GND.n3932 9.3005
R14454 GND.n2226 GND.n2225 9.3005
R14455 GND.n3946 GND.n3945 9.3005
R14456 GND.n3947 GND.n2224 9.3005
R14457 GND.n3949 GND.n3948 9.3005
R14458 GND.n2212 GND.n2211 9.3005
R14459 GND.n3962 GND.n3961 9.3005
R14460 GND.n3963 GND.n2210 9.3005
R14461 GND.n3965 GND.n3964 9.3005
R14462 GND.n2196 GND.n2195 9.3005
R14463 GND.n3978 GND.n3977 9.3005
R14464 GND.n3979 GND.n2194 9.3005
R14465 GND.n3981 GND.n3980 9.3005
R14466 GND.n2181 GND.n2180 9.3005
R14467 GND.n3994 GND.n3993 9.3005
R14468 GND.n3995 GND.n2179 9.3005
R14469 GND.n3997 GND.n3996 9.3005
R14470 GND.n2167 GND.n2166 9.3005
R14471 GND.n4010 GND.n4009 9.3005
R14472 GND.n4011 GND.n2165 9.3005
R14473 GND.n4013 GND.n4012 9.3005
R14474 GND.n2152 GND.n2151 9.3005
R14475 GND.n4026 GND.n4025 9.3005
R14476 GND.n4027 GND.n2150 9.3005
R14477 GND.n4029 GND.n4028 9.3005
R14478 GND.n2138 GND.n2137 9.3005
R14479 GND.n4042 GND.n4041 9.3005
R14480 GND.n4043 GND.n2136 9.3005
R14481 GND.n4045 GND.n4044 9.3005
R14482 GND.n2124 GND.n2123 9.3005
R14483 GND.n4058 GND.n4057 9.3005
R14484 GND.n4059 GND.n2122 9.3005
R14485 GND.n4061 GND.n4060 9.3005
R14486 GND.n2109 GND.n2108 9.3005
R14487 GND.n4074 GND.n4073 9.3005
R14488 GND.n4075 GND.n2107 9.3005
R14489 GND.n4077 GND.n4076 9.3005
R14490 GND.n2095 GND.n2094 9.3005
R14491 GND.n4090 GND.n4089 9.3005
R14492 GND.n4091 GND.n2093 9.3005
R14493 GND.n4093 GND.n4092 9.3005
R14494 GND.n2081 GND.n2080 9.3005
R14495 GND.n4105 GND.n4104 9.3005
R14496 GND.n4106 GND.n2079 9.3005
R14497 GND.n4108 GND.n4107 9.3005
R14498 GND.n2065 GND.n2064 9.3005
R14499 GND.n4121 GND.n4120 9.3005
R14500 GND.n4122 GND.n2063 9.3005
R14501 GND.n4124 GND.n4123 9.3005
R14502 GND.n2051 GND.n2050 9.3005
R14503 GND.n4139 GND.n4138 9.3005
R14504 GND.n4140 GND.n2049 9.3005
R14505 GND.n4145 GND.n4141 9.3005
R14506 GND.n4144 GND.n4143 9.3005
R14507 GND.n4142 GND.n1559 9.3005
R14508 GND.n4694 GND.n1560 9.3005
R14509 GND.n4693 GND.n1561 9.3005
R14510 GND.n4692 GND.n1562 9.3005
R14511 GND.n1830 GND.n1563 9.3005
R14512 GND.n1832 GND.n1831 9.3005
R14513 GND.n1829 GND.n1828 9.3005
R14514 GND.n1837 GND.n1836 9.3005
R14515 GND.n1838 GND.n1827 9.3005
R14516 GND.n1840 GND.n1839 9.3005
R14517 GND.n1825 GND.n1824 9.3005
R14518 GND.n1845 GND.n1844 9.3005
R14519 GND.n1846 GND.n1823 9.3005
R14520 GND.n1848 GND.n1847 9.3005
R14521 GND.n1821 GND.n1820 9.3005
R14522 GND.n1853 GND.n1852 9.3005
R14523 GND.n1854 GND.n1819 9.3005
R14524 GND.n1856 GND.n1855 9.3005
R14525 GND.n1817 GND.n1816 9.3005
R14526 GND.n1861 GND.n1860 9.3005
R14527 GND.n1862 GND.n1815 9.3005
R14528 GND.n1864 GND.n1863 9.3005
R14529 GND.n1813 GND.n1812 9.3005
R14530 GND.n1869 GND.n1868 9.3005
R14531 GND.n1870 GND.n1811 9.3005
R14532 GND.n1872 GND.n1871 9.3005
R14533 GND.n1809 GND.n1808 9.3005
R14534 GND.n1878 GND.n1877 9.3005
R14535 GND.n1879 GND.n1807 9.3005
R14536 GND.n1881 GND.n1880 9.3005
R14537 GND.n4289 GND.n4288 9.3005
R14538 GND.n4280 GND.n4279 9.3005
R14539 GND.n4294 GND.n4293 9.3005
R14540 GND.n4295 GND.n4278 9.3005
R14541 GND.n4469 GND.n4296 9.3005
R14542 GND.n4468 GND.n4297 9.3005
R14543 GND.n4467 GND.n4298 9.3005
R14544 GND.n4301 GND.n4299 9.3005
R14545 GND.n4463 GND.n4302 9.3005
R14546 GND.n4462 GND.n4303 9.3005
R14547 GND.n4461 GND.n4304 9.3005
R14548 GND.n4307 GND.n4305 9.3005
R14549 GND.n4457 GND.n4308 9.3005
R14550 GND.n4456 GND.n4309 9.3005
R14551 GND.n4455 GND.n4310 9.3005
R14552 GND.n4313 GND.n4311 9.3005
R14553 GND.n4327 GND.n4314 9.3005
R14554 GND.n4326 GND.n4315 9.3005
R14555 GND.n4325 GND.n4316 9.3005
R14556 GND.n4318 GND.n4317 9.3005
R14557 GND.n4321 GND.n4320 9.3005
R14558 GND.n4319 GND.n390 9.3005
R14559 GND.n6156 GND.n391 9.3005
R14560 GND.n6155 GND.n392 9.3005
R14561 GND.n6154 GND.n393 9.3005
R14562 GND.n398 GND.n394 9.3005
R14563 GND.n6148 GND.n399 9.3005
R14564 GND.n6147 GND.n400 9.3005
R14565 GND.n6146 GND.n401 9.3005
R14566 GND.n406 GND.n402 9.3005
R14567 GND.n6140 GND.n407 9.3005
R14568 GND.n6139 GND.n408 9.3005
R14569 GND.n6138 GND.n409 9.3005
R14570 GND.n414 GND.n410 9.3005
R14571 GND.n6132 GND.n415 9.3005
R14572 GND.n6131 GND.n416 9.3005
R14573 GND.n6130 GND.n417 9.3005
R14574 GND.n422 GND.n418 9.3005
R14575 GND.n6124 GND.n423 9.3005
R14576 GND.n6123 GND.n424 9.3005
R14577 GND.n6122 GND.n425 9.3005
R14578 GND.n430 GND.n426 9.3005
R14579 GND.n6116 GND.n431 9.3005
R14580 GND.n6115 GND.n432 9.3005
R14581 GND.n6114 GND.n433 9.3005
R14582 GND.n438 GND.n434 9.3005
R14583 GND.n6108 GND.n439 9.3005
R14584 GND.n6107 GND.n440 9.3005
R14585 GND.n6106 GND.n441 9.3005
R14586 GND.n446 GND.n442 9.3005
R14587 GND.n6100 GND.n447 9.3005
R14588 GND.n6099 GND.n448 9.3005
R14589 GND.n6098 GND.n449 9.3005
R14590 GND.n454 GND.n450 9.3005
R14591 GND.n6092 GND.n455 9.3005
R14592 GND.n6091 GND.n456 9.3005
R14593 GND.n6090 GND.n457 9.3005
R14594 GND.n462 GND.n458 9.3005
R14595 GND.n6084 GND.n463 9.3005
R14596 GND.n6083 GND.n464 9.3005
R14597 GND.n6082 GND.n465 9.3005
R14598 GND.n470 GND.n466 9.3005
R14599 GND.n6076 GND.n471 9.3005
R14600 GND.n6075 GND.n6074 9.3005
R14601 GND.n3483 GND.n3482 9.3005
R14602 GND.n3481 GND.n3313 9.3005
R14603 GND.n3480 GND.n3479 9.3005
R14604 GND.n3315 GND.n3314 9.3005
R14605 GND.n3473 GND.n3472 9.3005
R14606 GND.n3471 GND.n3317 9.3005
R14607 GND.n3470 GND.n3469 9.3005
R14608 GND.n3319 GND.n3318 9.3005
R14609 GND.n3463 GND.n3462 9.3005
R14610 GND.n3461 GND.n3321 9.3005
R14611 GND.n3460 GND.n3459 9.3005
R14612 GND.n3323 GND.n3322 9.3005
R14613 GND.n3453 GND.n3449 9.3005
R14614 GND.n3448 GND.n3325 9.3005
R14615 GND.n3447 GND.n3446 9.3005
R14616 GND.n3327 GND.n3326 9.3005
R14617 GND.n3440 GND.n3439 9.3005
R14618 GND.n3438 GND.n3329 9.3005
R14619 GND.n3437 GND.n3436 9.3005
R14620 GND.n3331 GND.n3330 9.3005
R14621 GND.n3430 GND.n3429 9.3005
R14622 GND.n3428 GND.n3333 9.3005
R14623 GND.n3427 GND.n3426 9.3005
R14624 GND.n3335 GND.n3334 9.3005
R14625 GND.n3420 GND.n3417 9.3005
R14626 GND.n3416 GND.n3337 9.3005
R14627 GND.n3415 GND.n3414 9.3005
R14628 GND.n3339 GND.n3338 9.3005
R14629 GND.n3408 GND.n3407 9.3005
R14630 GND.n3406 GND.n3341 9.3005
R14631 GND.n3405 GND.n3404 9.3005
R14632 GND.n3343 GND.n3342 9.3005
R14633 GND.n3398 GND.n3397 9.3005
R14634 GND.n3396 GND.n3345 9.3005
R14635 GND.n3395 GND.n3394 9.3005
R14636 GND.n3347 GND.n3346 9.3005
R14637 GND.n3388 GND.n3387 9.3005
R14638 GND.n3385 GND.n3384 9.3005
R14639 GND.n3353 GND.n3352 9.3005
R14640 GND.n3378 GND.n3377 9.3005
R14641 GND.n3376 GND.n3355 9.3005
R14642 GND.n3375 GND.n3374 9.3005
R14643 GND.n3357 GND.n3356 9.3005
R14644 GND.n3368 GND.n3367 9.3005
R14645 GND.n3366 GND.n3359 9.3005
R14646 GND.n3365 GND.n3364 9.3005
R14647 GND.n3361 GND.n3360 9.3005
R14648 GND.n3386 GND.n3351 9.3005
R14649 GND.n3311 GND.n3308 9.3005
R14650 GND.n3489 GND.n3488 9.3005
R14651 GND.n5041 GND.n1170 9.3005
R14652 GND.n5040 GND.n1171 9.3005
R14653 GND.n3289 GND.n1172 9.3005
R14654 GND.n3615 GND.n3614 9.3005
R14655 GND.n3616 GND.n3288 9.3005
R14656 GND.n3620 GND.n3617 9.3005
R14657 GND.n3619 GND.n3618 9.3005
R14658 GND.n3267 GND.n3266 9.3005
R14659 GND.n3639 GND.n3638 9.3005
R14660 GND.n3640 GND.n3265 9.3005
R14661 GND.n3644 GND.n3641 9.3005
R14662 GND.n3643 GND.n3642 9.3005
R14663 GND.n3244 GND.n3243 9.3005
R14664 GND.n3664 GND.n3663 9.3005
R14665 GND.n3665 GND.n3242 9.3005
R14666 GND.n3669 GND.n3666 9.3005
R14667 GND.n3668 GND.n3667 9.3005
R14668 GND.n3222 GND.n3221 9.3005
R14669 GND.n3689 GND.n3688 9.3005
R14670 GND.n3690 GND.n3220 9.3005
R14671 GND.n3692 GND.n3691 9.3005
R14672 GND.n3075 GND.n3068 9.3005
R14673 GND.n3764 GND.n3761 9.3005
R14674 GND.n3763 GND.n3762 9.3005
R14675 GND.n3046 GND.n3045 9.3005
R14676 GND.n3784 GND.n3783 9.3005
R14677 GND.n3785 GND.n3044 9.3005
R14678 GND.n3789 GND.n3786 9.3005
R14679 GND.n3788 GND.n3787 9.3005
R14680 GND.n3023 GND.n3022 9.3005
R14681 GND.n3808 GND.n3807 9.3005
R14682 GND.n3809 GND.n3021 9.3005
R14683 GND.n3813 GND.n3810 9.3005
R14684 GND.n3812 GND.n3811 9.3005
R14685 GND.n3000 GND.n2999 9.3005
R14686 GND.n3833 GND.n3832 9.3005
R14687 GND.n3834 GND.n2998 9.3005
R14688 GND.n3838 GND.n3835 9.3005
R14689 GND.n3837 GND.n3836 9.3005
R14690 GND.n2978 GND.n2977 9.3005
R14691 GND.n3861 GND.n3860 9.3005
R14692 GND.n3862 GND.n2976 9.3005
R14693 GND.n3864 GND.n3863 9.3005
R14694 GND.n1298 GND.n1297 9.3005
R14695 GND.n4951 GND.n4950 9.3005
R14696 GND.n5042 GND.n1169 9.3005
R14697 GND.n3760 GND.n3073 9.3005
R14698 GND.n3760 GND.n3067 9.3005
R14699 GND.n1081 GND.n1080 9.3005
R14700 GND.n5122 GND.n1085 9.3005
R14701 GND.n5121 GND.n1086 9.3005
R14702 GND.n5120 GND.n1087 9.3005
R14703 GND.n1092 GND.n1088 9.3005
R14704 GND.n5114 GND.n1093 9.3005
R14705 GND.n5113 GND.n1094 9.3005
R14706 GND.n5112 GND.n1095 9.3005
R14707 GND.n1100 GND.n1096 9.3005
R14708 GND.n5106 GND.n1101 9.3005
R14709 GND.n5105 GND.n1102 9.3005
R14710 GND.n5104 GND.n1103 9.3005
R14711 GND.n1108 GND.n1104 9.3005
R14712 GND.n5098 GND.n1109 9.3005
R14713 GND.n5097 GND.n1110 9.3005
R14714 GND.n5096 GND.n1111 9.3005
R14715 GND.n1116 GND.n1112 9.3005
R14716 GND.n5090 GND.n1117 9.3005
R14717 GND.n5089 GND.n1118 9.3005
R14718 GND.n5088 GND.n1119 9.3005
R14719 GND.n1124 GND.n1120 9.3005
R14720 GND.n5082 GND.n1125 9.3005
R14721 GND.n5081 GND.n1126 9.3005
R14722 GND.n5080 GND.n1127 9.3005
R14723 GND.n1132 GND.n1128 9.3005
R14724 GND.n5074 GND.n1133 9.3005
R14725 GND.n5073 GND.n1134 9.3005
R14726 GND.n5072 GND.n1135 9.3005
R14727 GND.n1140 GND.n1136 9.3005
R14728 GND.n5066 GND.n1141 9.3005
R14729 GND.n5065 GND.n1142 9.3005
R14730 GND.n5064 GND.n1143 9.3005
R14731 GND.n1148 GND.n1144 9.3005
R14732 GND.n5058 GND.n1149 9.3005
R14733 GND.n5057 GND.n1150 9.3005
R14734 GND.n5056 GND.n1151 9.3005
R14735 GND.n1156 GND.n1152 9.3005
R14736 GND.n5050 GND.n1157 9.3005
R14737 GND.n5049 GND.n1158 9.3005
R14738 GND.n5048 GND.n1159 9.3005
R14739 GND.n3542 GND.n1160 9.3005
R14740 GND.n3544 GND.n3543 9.3005
R14741 GND.n3541 GND.n3540 9.3005
R14742 GND.n3549 GND.n3548 9.3005
R14743 GND.n3550 GND.n3539 9.3005
R14744 GND.n3605 GND.n3551 9.3005
R14745 GND.n3604 GND.n3552 9.3005
R14746 GND.n3603 GND.n3553 9.3005
R14747 GND.n3556 GND.n3554 9.3005
R14748 GND.n3599 GND.n3557 9.3005
R14749 GND.n3598 GND.n3558 9.3005
R14750 GND.n3597 GND.n3559 9.3005
R14751 GND.n3562 GND.n3560 9.3005
R14752 GND.n3593 GND.n3563 9.3005
R14753 GND.n3592 GND.n3564 9.3005
R14754 GND.n3591 GND.n3565 9.3005
R14755 GND.n3568 GND.n3566 9.3005
R14756 GND.n3587 GND.n3569 9.3005
R14757 GND.n3586 GND.n3570 9.3005
R14758 GND.n3585 GND.n3571 9.3005
R14759 GND.n3574 GND.n3572 9.3005
R14760 GND.n3581 GND.n3575 9.3005
R14761 GND.n3580 GND.n3576 9.3005
R14762 GND.n5129 GND.n5128 9.3005
R14763 GND.n5132 GND.n1079 9.3005
R14764 GND.n1078 GND.n1074 9.3005
R14765 GND.n5138 GND.n1073 9.3005
R14766 GND.n5139 GND.n1072 9.3005
R14767 GND.n5140 GND.n1071 9.3005
R14768 GND.n1070 GND.n1066 9.3005
R14769 GND.n5146 GND.n1065 9.3005
R14770 GND.n5147 GND.n1064 9.3005
R14771 GND.n5148 GND.n1063 9.3005
R14772 GND.n1062 GND.n1058 9.3005
R14773 GND.n5154 GND.n1057 9.3005
R14774 GND.n5155 GND.n1056 9.3005
R14775 GND.n5156 GND.n1055 9.3005
R14776 GND.n1054 GND.n1050 9.3005
R14777 GND.n5162 GND.n1049 9.3005
R14778 GND.n5163 GND.n1048 9.3005
R14779 GND.n5164 GND.n1047 9.3005
R14780 GND.n1046 GND.n1042 9.3005
R14781 GND.n5170 GND.n1041 9.3005
R14782 GND.n5171 GND.n1040 9.3005
R14783 GND.n5172 GND.n1039 9.3005
R14784 GND.n1038 GND.n1034 9.3005
R14785 GND.n5178 GND.n1033 9.3005
R14786 GND.n5179 GND.n1032 9.3005
R14787 GND.n5180 GND.n1031 9.3005
R14788 GND.n1030 GND.n1026 9.3005
R14789 GND.n5186 GND.n1025 9.3005
R14790 GND.n5187 GND.n1024 9.3005
R14791 GND.n5188 GND.n1023 9.3005
R14792 GND.n1022 GND.n1018 9.3005
R14793 GND.n5194 GND.n1017 9.3005
R14794 GND.n5195 GND.n1016 9.3005
R14795 GND.n5196 GND.n1015 9.3005
R14796 GND.n1014 GND.n1010 9.3005
R14797 GND.n5202 GND.n1009 9.3005
R14798 GND.n5203 GND.n1008 9.3005
R14799 GND.n5204 GND.n1007 9.3005
R14800 GND.n1006 GND.n1002 9.3005
R14801 GND.n5210 GND.n1001 9.3005
R14802 GND.n5211 GND.n1000 9.3005
R14803 GND.n5212 GND.n999 9.3005
R14804 GND.n998 GND.n994 9.3005
R14805 GND.n5218 GND.n993 9.3005
R14806 GND.n5219 GND.n992 9.3005
R14807 GND.n5220 GND.n991 9.3005
R14808 GND.n990 GND.n986 9.3005
R14809 GND.n5226 GND.n985 9.3005
R14810 GND.n5227 GND.n984 9.3005
R14811 GND.n5228 GND.n983 9.3005
R14812 GND.n982 GND.n978 9.3005
R14813 GND.n5234 GND.n977 9.3005
R14814 GND.n5235 GND.n976 9.3005
R14815 GND.n5236 GND.n975 9.3005
R14816 GND.n971 GND.n970 9.3005
R14817 GND.n5243 GND.n5242 9.3005
R14818 GND.n5131 GND.n5130 9.3005
R14819 GND.n1402 GND.n1400 9.3005
R14820 GND.n4812 GND.n4809 9.3005
R14821 GND.n4814 GND.n4813 9.3005
R14822 GND.n4815 GND.n4808 9.3005
R14823 GND.n4817 GND.n4816 9.3005
R14824 GND.n4818 GND.n4804 9.3005
R14825 GND.n4820 GND.n4819 9.3005
R14826 GND.n4821 GND.n1466 9.3005
R14827 GND.n4823 GND.n4822 9.3005
R14828 GND.n4801 GND.n1467 9.3005
R14829 GND.n4800 GND.n4799 9.3005
R14830 GND.n4798 GND.n1470 9.3005
R14831 GND.n4797 GND.n4796 9.3005
R14832 GND.n4795 GND.n1471 9.3005
R14833 GND.n4794 GND.n4793 9.3005
R14834 GND.n4792 GND.n1475 9.3005
R14835 GND.n4791 GND.n4790 9.3005
R14836 GND.n4789 GND.n1476 9.3005
R14837 GND.n4788 GND.n4787 9.3005
R14838 GND.n4786 GND.n1480 9.3005
R14839 GND.n4785 GND.n4784 9.3005
R14840 GND.n4783 GND.n1481 9.3005
R14841 GND.n4782 GND.n4781 9.3005
R14842 GND.n4780 GND.n1485 9.3005
R14843 GND.n4779 GND.n4778 9.3005
R14844 GND.n4777 GND.n1486 9.3005
R14845 GND.n4776 GND.n4775 9.3005
R14846 GND.n4774 GND.n1490 9.3005
R14847 GND.n4773 GND.n4772 9.3005
R14848 GND.n4771 GND.n1491 9.3005
R14849 GND.n4770 GND.n4769 9.3005
R14850 GND.n4768 GND.n1495 9.3005
R14851 GND.n4767 GND.n4766 9.3005
R14852 GND.n4765 GND.n1496 9.3005
R14853 GND.n4764 GND.n4763 9.3005
R14854 GND.n4762 GND.n1500 9.3005
R14855 GND.n4761 GND.n4760 9.3005
R14856 GND.n4759 GND.n1501 9.3005
R14857 GND.n4758 GND.n4757 9.3005
R14858 GND.n4756 GND.n1505 9.3005
R14859 GND.n4755 GND.n4754 9.3005
R14860 GND.n4753 GND.n1506 9.3005
R14861 GND.n4752 GND.n4751 9.3005
R14862 GND.n4750 GND.n1510 9.3005
R14863 GND.n4749 GND.n4748 9.3005
R14864 GND.n4747 GND.n1511 9.3005
R14865 GND.n4746 GND.n4745 9.3005
R14866 GND.n4744 GND.n1515 9.3005
R14867 GND.n4743 GND.n4742 9.3005
R14868 GND.n4741 GND.n1516 9.3005
R14869 GND.n4740 GND.n4739 9.3005
R14870 GND.n4738 GND.n1520 9.3005
R14871 GND.n4737 GND.n4736 9.3005
R14872 GND.n4735 GND.n1521 9.3005
R14873 GND.n4734 GND.n4733 9.3005
R14874 GND.n4732 GND.n1525 9.3005
R14875 GND.n4731 GND.n4730 9.3005
R14876 GND.n4729 GND.n1526 9.3005
R14877 GND.n4728 GND.n4727 9.3005
R14878 GND.n4726 GND.n1530 9.3005
R14879 GND.n4725 GND.n4724 9.3005
R14880 GND.n4723 GND.n1531 9.3005
R14881 GND.n4722 GND.n4721 9.3005
R14882 GND.n4720 GND.n1535 9.3005
R14883 GND.n4719 GND.n4718 9.3005
R14884 GND.n4717 GND.n1536 9.3005
R14885 GND.n4716 GND.n4715 9.3005
R14886 GND.n4714 GND.n1540 9.3005
R14887 GND.n4713 GND.n4712 9.3005
R14888 GND.n4711 GND.n1541 9.3005
R14889 GND.n4710 GND.n4709 9.3005
R14890 GND.n4708 GND.n1545 9.3005
R14891 GND.n4707 GND.n4706 9.3005
R14892 GND.n4705 GND.n1546 9.3005
R14893 GND.n4704 GND.n4703 9.3005
R14894 GND.n4702 GND.n1550 9.3005
R14895 GND.n4701 GND.n4700 9.3005
R14896 GND.n4699 GND.n1551 9.3005
R14897 GND.n4803 GND.n4802 9.3005
R14898 GND.n1959 GND.n1956 9.3005
R14899 GND.n1965 GND.n1964 9.3005
R14900 GND.n1966 GND.n1955 9.3005
R14901 GND.n1968 GND.n1967 9.3005
R14902 GND.n1953 GND.n1952 9.3005
R14903 GND.n1975 GND.n1974 9.3005
R14904 GND.n1976 GND.n1951 9.3005
R14905 GND.n1978 GND.n1977 9.3005
R14906 GND.n1958 GND.n1957 9.3005
R14907 GND.n2029 GND.n2028 9.3005
R14908 GND.n1933 GND.n1931 9.3005
R14909 GND.n2014 GND.n2013 9.3005
R14910 GND.n2010 GND.n1937 9.3005
R14911 GND.n2007 GND.n2006 9.3005
R14912 GND.n1940 GND.n1939 9.3005
R14913 GND.n1995 GND.n1994 9.3005
R14914 GND.n1991 GND.n1944 9.3005
R14915 GND.n1988 GND.n1987 9.3005
R14916 GND.n1947 GND.n1946 9.3005
R14917 GND.n2030 GND.n1927 9.3005
R14918 GND.n2033 GND.n2032 9.3005
R14919 GND.n1949 GND.n1948 9.3005
R14920 GND.n1985 GND.n1984 9.3005
R14921 GND.n1986 GND.n1943 9.3005
R14922 GND.n1997 GND.n1996 9.3005
R14923 GND.n1945 GND.n1941 9.3005
R14924 GND.n2004 GND.n2003 9.3005
R14925 GND.n2005 GND.n1936 9.3005
R14926 GND.n2016 GND.n2015 9.3005
R14927 GND.n1938 GND.n1934 9.3005
R14928 GND.n2026 GND.n2025 9.3005
R14929 GND.n2027 GND.n1926 9.3005
R14930 GND.n2035 GND.n2034 9.3005
R14931 GND.n1924 GND.n1923 9.3005
R14932 GND.n2041 GND.n2040 9.3005
R14933 GND.n3877 GND.n3876 9.3005
R14934 GND.n2957 GND.n2956 9.3005
R14935 GND.n3890 GND.n3889 9.3005
R14936 GND.n3891 GND.n2955 9.3005
R14937 GND.n3893 GND.n3892 9.3005
R14938 GND.n2262 GND.n2261 9.3005
R14939 GND.n3906 GND.n3905 9.3005
R14940 GND.n3907 GND.n2260 9.3005
R14941 GND.n3909 GND.n3908 9.3005
R14942 GND.n2247 GND.n2246 9.3005
R14943 GND.n3922 GND.n3921 9.3005
R14944 GND.n3923 GND.n2245 9.3005
R14945 GND.n3925 GND.n3924 9.3005
R14946 GND.n2233 GND.n2232 9.3005
R14947 GND.n3938 GND.n3937 9.3005
R14948 GND.n3939 GND.n2231 9.3005
R14949 GND.n3941 GND.n3940 9.3005
R14950 GND.n2218 GND.n2217 9.3005
R14951 GND.n3954 GND.n3953 9.3005
R14952 GND.n3955 GND.n2216 9.3005
R14953 GND.n3957 GND.n3956 9.3005
R14954 GND.n2204 GND.n2203 9.3005
R14955 GND.n3970 GND.n3969 9.3005
R14956 GND.n3971 GND.n2202 9.3005
R14957 GND.n3973 GND.n3972 9.3005
R14958 GND.n2188 GND.n2187 9.3005
R14959 GND.n3986 GND.n3985 9.3005
R14960 GND.n3987 GND.n2186 9.3005
R14961 GND.n3989 GND.n3988 9.3005
R14962 GND.n2174 GND.n2173 9.3005
R14963 GND.n4002 GND.n4001 9.3005
R14964 GND.n4003 GND.n2172 9.3005
R14965 GND.n4005 GND.n4004 9.3005
R14966 GND.n2159 GND.n2158 9.3005
R14967 GND.n4018 GND.n4017 9.3005
R14968 GND.n4019 GND.n2157 9.3005
R14969 GND.n4021 GND.n4020 9.3005
R14970 GND.n2145 GND.n2144 9.3005
R14971 GND.n4034 GND.n4033 9.3005
R14972 GND.n4035 GND.n2143 9.3005
R14973 GND.n4037 GND.n4036 9.3005
R14974 GND.n2131 GND.n2130 9.3005
R14975 GND.n4050 GND.n4049 9.3005
R14976 GND.n4051 GND.n2129 9.3005
R14977 GND.n4053 GND.n4052 9.3005
R14978 GND.n2116 GND.n2115 9.3005
R14979 GND.n4066 GND.n4065 9.3005
R14980 GND.n4067 GND.n2114 9.3005
R14981 GND.n4069 GND.n4068 9.3005
R14982 GND.n2101 GND.n2100 9.3005
R14983 GND.n4082 GND.n4081 9.3005
R14984 GND.n4083 GND.n2099 9.3005
R14985 GND.n4085 GND.n4084 9.3005
R14986 GND.n2088 GND.n2087 9.3005
R14987 GND.n4097 GND.n4096 9.3005
R14988 GND.n4098 GND.n2086 9.3005
R14989 GND.n4100 GND.n4099 9.3005
R14990 GND.n2072 GND.n2071 9.3005
R14991 GND.n4113 GND.n4112 9.3005
R14992 GND.n4114 GND.n2070 9.3005
R14993 GND.n4116 GND.n4115 9.3005
R14994 GND.n2058 GND.n2057 9.3005
R14995 GND.n4129 GND.n4128 9.3005
R14996 GND.n4130 GND.n2055 9.3005
R14997 GND.n4134 GND.n4133 9.3005
R14998 GND.n4132 GND.n2056 9.3005
R14999 GND.n4131 GND.n2043 9.3005
R15000 GND.n4150 GND.n2042 9.3005
R15001 GND.n4152 GND.n4151 9.3005
R15002 GND.n3875 GND.n2967 9.3005
R15003 GND.n3710 GND.n3206 9.3005
R15004 GND.n3712 GND.n3711 9.3005
R15005 GND.n3713 GND.n3205 9.3005
R15006 GND.n3715 GND.n3714 9.3005
R15007 GND.n3058 GND.n3057 9.3005
R15008 GND.n3769 GND.n3768 9.3005
R15009 GND.n3770 GND.n3055 9.3005
R15010 GND.n3773 GND.n3772 9.3005
R15011 GND.n3771 GND.n3056 9.3005
R15012 GND.n3036 GND.n3035 9.3005
R15013 GND.n3794 GND.n3793 9.3005
R15014 GND.n3795 GND.n3033 9.3005
R15015 GND.n3798 GND.n3797 9.3005
R15016 GND.n3796 GND.n3034 9.3005
R15017 GND.n3012 GND.n3011 9.3005
R15018 GND.n3818 GND.n3817 9.3005
R15019 GND.n3819 GND.n3009 9.3005
R15020 GND.n3822 GND.n3821 9.3005
R15021 GND.n3820 GND.n3010 9.3005
R15022 GND.n2989 GND.n2988 9.3005
R15023 GND.n3843 GND.n3842 9.3005
R15024 GND.n3844 GND.n2986 9.3005
R15025 GND.n3852 GND.n3851 9.3005
R15026 GND.n3850 GND.n2987 9.3005
R15027 GND.n3849 GND.n3848 9.3005
R15028 GND.n3845 GND.n2969 9.3005
R15029 GND.n3871 GND.n2968 9.3005
R15030 GND.n3873 GND.n3872 9.3005
R15031 GND.n4864 GND.n4863 9.3005
R15032 GND.n4862 GND.n4861 9.3005
R15033 GND.n1413 GND.n1412 9.3005
R15034 GND.n4856 GND.n4855 9.3005
R15035 GND.n4854 GND.n4853 9.3005
R15036 GND.n1424 GND.n1423 9.3005
R15037 GND.n4848 GND.n4847 9.3005
R15038 GND.n4846 GND.n4845 9.3005
R15039 GND.n1434 GND.n1433 9.3005
R15040 GND.n4837 GND.n4836 9.3005
R15041 GND.n4835 GND.n4832 9.3005
R15042 GND.n1407 GND.n1401 9.3005
R15043 GND.n4831 GND.n4830 9.3005
R15044 GND.n1438 GND.n1437 9.3005
R15045 GND.n4839 GND.n4838 9.3005
R15046 GND.n4844 GND.n4843 9.3005
R15047 GND.n1428 GND.n1427 9.3005
R15048 GND.n4850 GND.n4849 9.3005
R15049 GND.n4852 GND.n4851 9.3005
R15050 GND.n1417 GND.n1416 9.3005
R15051 GND.n4858 GND.n4857 9.3005
R15052 GND.n4860 GND.n4859 9.3005
R15053 GND.n1406 GND.n1405 9.3005
R15054 GND.n4866 GND.n4865 9.3005
R15055 GND.n4868 GND.n4867 9.3005
R15056 GND.n4829 GND.n1444 9.3005
R15057 GND.n4918 GND.n4917 9.3005
R15058 GND.n4919 GND.n1326 9.3005
R15059 GND.n4921 GND.n4920 9.3005
R15060 GND.n4922 GND.n1322 9.3005
R15061 GND.n4924 GND.n4923 9.3005
R15062 GND.n4925 GND.n1321 9.3005
R15063 GND.n4927 GND.n4926 9.3005
R15064 GND.n4928 GND.n1317 9.3005
R15065 GND.n4930 GND.n4929 9.3005
R15066 GND.n4931 GND.n1316 9.3005
R15067 GND.n4933 GND.n4932 9.3005
R15068 GND.n4934 GND.n1313 9.3005
R15069 GND.n4935 GND.n1308 9.3005
R15070 GND.n4937 GND.n4936 9.3005
R15071 GND.n4938 GND.n1307 9.3005
R15072 GND.n4940 GND.n4939 9.3005
R15073 GND.n4941 GND.n1303 9.3005
R15074 GND.n4943 GND.n4942 9.3005
R15075 GND.n4944 GND.n1302 9.3005
R15076 GND.n4946 GND.n4945 9.3005
R15077 GND.n4947 GND.n1299 9.3005
R15078 GND.n4949 GND.n4948 9.3005
R15079 GND.n1350 GND.n1347 9.3005
R15080 GND.n4909 GND.n4908 9.3005
R15081 GND.n4907 GND.n1349 9.3005
R15082 GND.n4906 GND.n4905 9.3005
R15083 GND.n4904 GND.n1351 9.3005
R15084 GND.n4903 GND.n4902 9.3005
R15085 GND.n4901 GND.n1357 9.3005
R15086 GND.n4900 GND.n4899 9.3005
R15087 GND.n4898 GND.n1358 9.3005
R15088 GND.n4897 GND.n4896 9.3005
R15089 GND.n4895 GND.n1365 9.3005
R15090 GND.n4894 GND.n4893 9.3005
R15091 GND.n4891 GND.n1366 9.3005
R15092 GND.n4890 GND.n4889 9.3005
R15093 GND.n4888 GND.n1375 9.3005
R15094 GND.n4887 GND.n4886 9.3005
R15095 GND.n4885 GND.n1376 9.3005
R15096 GND.n4884 GND.n4883 9.3005
R15097 GND.n4882 GND.n1383 9.3005
R15098 GND.n4881 GND.n4880 9.3005
R15099 GND.n4879 GND.n1384 9.3005
R15100 GND.n4878 GND.n4877 9.3005
R15101 GND.n4876 GND.n1391 9.3005
R15102 GND.n4875 GND.n4874 9.3005
R15103 GND.n4873 GND.n1392 9.3005
R15104 GND.n4872 GND.n4871 9.3005
R15105 GND.n1182 GND.n1180 9.3005
R15106 GND.n5036 GND.n5035 9.3005
R15107 GND.n1183 GND.n1181 9.3005
R15108 GND.n5031 GND.n1188 9.3005
R15109 GND.n5030 GND.n1189 9.3005
R15110 GND.n5029 GND.n1190 9.3005
R15111 GND.n3273 GND.n1191 9.3005
R15112 GND.n5025 GND.n1196 9.3005
R15113 GND.n5024 GND.n1197 9.3005
R15114 GND.n5023 GND.n1198 9.3005
R15115 GND.n3260 GND.n1199 9.3005
R15116 GND.n5019 GND.n1204 9.3005
R15117 GND.n5018 GND.n1205 9.3005
R15118 GND.n5017 GND.n1206 9.3005
R15119 GND.n3657 GND.n1207 9.3005
R15120 GND.n5013 GND.n1212 9.3005
R15121 GND.n5012 GND.n1213 9.3005
R15122 GND.n5011 GND.n1214 9.3005
R15123 GND.n3684 GND.n1215 9.3005
R15124 GND.n5007 GND.n1220 9.3005
R15125 GND.n5006 GND.n1221 9.3005
R15126 GND.n5005 GND.n1222 9.3005
R15127 GND.n3754 GND.n1223 9.3005
R15128 GND.n5001 GND.n1228 9.3005
R15129 GND.n5000 GND.n1229 9.3005
R15130 GND.n4999 GND.n1230 9.3005
R15131 GND.n3095 GND.n1231 9.3005
R15132 GND.n4995 GND.n1236 9.3005
R15133 GND.n4994 GND.n1237 9.3005
R15134 GND.n4993 GND.n1238 9.3005
R15135 GND.n3723 GND.n1239 9.3005
R15136 GND.n4989 GND.n1244 9.3005
R15137 GND.n4988 GND.n1245 9.3005
R15138 GND.n4987 GND.n1246 9.3005
R15139 GND.n3052 GND.n1247 9.3005
R15140 GND.n4983 GND.n1252 9.3005
R15141 GND.n4982 GND.n1253 9.3005
R15142 GND.n4981 GND.n1254 9.3005
R15143 GND.n3029 GND.n1255 9.3005
R15144 GND.n4977 GND.n1260 9.3005
R15145 GND.n4976 GND.n1261 9.3005
R15146 GND.n4975 GND.n1262 9.3005
R15147 GND.n3016 GND.n1263 9.3005
R15148 GND.n4971 GND.n1268 9.3005
R15149 GND.n4970 GND.n1269 9.3005
R15150 GND.n4969 GND.n1270 9.3005
R15151 GND.n3826 GND.n1271 9.3005
R15152 GND.n4965 GND.n1276 9.3005
R15153 GND.n4964 GND.n1277 9.3005
R15154 GND.n4963 GND.n1278 9.3005
R15155 GND.n3856 GND.n1279 9.3005
R15156 GND.n4959 GND.n1284 9.3005
R15157 GND.n4958 GND.n1285 9.3005
R15158 GND.n4957 GND.n1286 9.3005
R15159 GND.n1293 GND.n1287 9.3005
R15160 GND.n3492 GND.n3490 9.3005
R15161 GND.n1184 GND.n1182 9.3005
R15162 GND.n5035 GND.n5034 9.3005
R15163 GND.n5033 GND.n1183 9.3005
R15164 GND.n5032 GND.n5031 9.3005
R15165 GND.n5030 GND.n1187 9.3005
R15166 GND.n5029 GND.n5028 9.3005
R15167 GND.n5027 GND.n1191 9.3005
R15168 GND.n5026 GND.n5025 9.3005
R15169 GND.n5024 GND.n1195 9.3005
R15170 GND.n5023 GND.n5022 9.3005
R15171 GND.n5021 GND.n1199 9.3005
R15172 GND.n5020 GND.n5019 9.3005
R15173 GND.n5018 GND.n1203 9.3005
R15174 GND.n5017 GND.n5016 9.3005
R15175 GND.n5015 GND.n1207 9.3005
R15176 GND.n5014 GND.n5013 9.3005
R15177 GND.n5012 GND.n1211 9.3005
R15178 GND.n5011 GND.n5010 9.3005
R15179 GND.n5009 GND.n1215 9.3005
R15180 GND.n5008 GND.n5007 9.3005
R15181 GND.n5006 GND.n1219 9.3005
R15182 GND.n5005 GND.n5004 9.3005
R15183 GND.n5003 GND.n1223 9.3005
R15184 GND.n5002 GND.n5001 9.3005
R15185 GND.n5000 GND.n1227 9.3005
R15186 GND.n4999 GND.n4998 9.3005
R15187 GND.n4997 GND.n1231 9.3005
R15188 GND.n4996 GND.n4995 9.3005
R15189 GND.n4994 GND.n1235 9.3005
R15190 GND.n4993 GND.n4992 9.3005
R15191 GND.n4991 GND.n1239 9.3005
R15192 GND.n4990 GND.n4989 9.3005
R15193 GND.n4988 GND.n1243 9.3005
R15194 GND.n4987 GND.n4986 9.3005
R15195 GND.n4985 GND.n1247 9.3005
R15196 GND.n4984 GND.n4983 9.3005
R15197 GND.n4982 GND.n1251 9.3005
R15198 GND.n4981 GND.n4980 9.3005
R15199 GND.n4979 GND.n1255 9.3005
R15200 GND.n4978 GND.n4977 9.3005
R15201 GND.n4976 GND.n1259 9.3005
R15202 GND.n4975 GND.n4974 9.3005
R15203 GND.n4973 GND.n1263 9.3005
R15204 GND.n4972 GND.n4971 9.3005
R15205 GND.n4970 GND.n1267 9.3005
R15206 GND.n4969 GND.n4968 9.3005
R15207 GND.n4967 GND.n1271 9.3005
R15208 GND.n4966 GND.n4965 9.3005
R15209 GND.n4964 GND.n1275 9.3005
R15210 GND.n4963 GND.n4962 9.3005
R15211 GND.n4961 GND.n1279 9.3005
R15212 GND.n4960 GND.n4959 9.3005
R15213 GND.n4958 GND.n1283 9.3005
R15214 GND.n4957 GND.n4956 9.3005
R15215 GND.n4955 GND.n1287 9.3005
R15216 GND.n3492 GND.n3491 9.3005
R15217 GND.n3514 GND.n3299 9.3005
R15218 GND.n3516 GND.n3515 9.3005
R15219 GND.n3513 GND.n3301 9.3005
R15220 GND.n3512 GND.n3511 9.3005
R15221 GND.n3303 GND.n3302 9.3005
R15222 GND.n3505 GND.n3504 9.3005
R15223 GND.n3503 GND.n3305 9.3005
R15224 GND.n3502 GND.n3501 9.3005
R15225 GND.n3307 GND.n3306 9.3005
R15226 GND.n3495 GND.n3494 9.3005
R15227 GND.n3298 GND.n3295 9.3005
R15228 GND.n3524 GND.n3523 9.3005
R15229 GND.n3530 GND.n3294 9.3005
R15230 GND.n3532 GND.n3531 9.3005
R15231 GND.n3533 GND.n3293 9.3005
R15232 GND.n3535 GND.n3534 9.3005
R15233 GND.n3280 GND.n3279 9.3005
R15234 GND.n3625 GND.n3624 9.3005
R15235 GND.n3626 GND.n3277 9.3005
R15236 GND.n3629 GND.n3628 9.3005
R15237 GND.n3627 GND.n3278 9.3005
R15238 GND.n3256 GND.n3255 9.3005
R15239 GND.n3649 GND.n3648 9.3005
R15240 GND.n3650 GND.n3253 9.3005
R15241 GND.n3653 GND.n3652 9.3005
R15242 GND.n3651 GND.n3254 9.3005
R15243 GND.n3233 GND.n3232 9.3005
R15244 GND.n3674 GND.n3673 9.3005
R15245 GND.n3675 GND.n3230 9.3005
R15246 GND.n3678 GND.n3677 9.3005
R15247 GND.n3676 GND.n3231 9.3005
R15248 GND.n3211 GND.n3210 9.3005
R15249 GND.n3697 GND.n3696 9.3005
R15250 GND.n3698 GND.n3209 9.3005
R15251 GND.n3700 GND.n3699 9.3005
R15252 GND.n3701 GND.n3208 9.3005
R15253 GND.n3705 GND.n3704 9.3005
R15254 GND.n3706 GND.n3207 9.3005
R15255 GND.n3709 GND.n3708 9.3005
R15256 GND.n3526 GND.n3525 9.3005
R15257 GND.n71 GND.n70 9.3005
R15258 GND.n56 GND.n55 9.3005
R15259 GND.n65 GND.n64 9.3005
R15260 GND.n63 GND.n62 9.3005
R15261 GND.n51 GND.n50 9.3005
R15262 GND.n36 GND.n35 9.3005
R15263 GND.n45 GND.n44 9.3005
R15264 GND.n43 GND.n42 9.3005
R15265 GND.n32 GND.n31 9.3005
R15266 GND.n17 GND.n16 9.3005
R15267 GND.n26 GND.n25 9.3005
R15268 GND.n24 GND.n23 9.3005
R15269 GND.n130 GND.n129 9.3005
R15270 GND.n115 GND.n114 9.3005
R15271 GND.n124 GND.n123 9.3005
R15272 GND.n122 GND.n121 9.3005
R15273 GND.n110 GND.n109 9.3005
R15274 GND.n95 GND.n94 9.3005
R15275 GND.n104 GND.n103 9.3005
R15276 GND.n102 GND.n101 9.3005
R15277 GND.n91 GND.n90 9.3005
R15278 GND.n76 GND.n75 9.3005
R15279 GND.n85 GND.n84 9.3005
R15280 GND.n83 GND.n82 9.3005
R15281 GND.n2802 GND.t164 9.04507
R15282 GND.t170 GND.n2120 9.04507
R15283 GND.n4917 GND.n1330 8.92171
R15284 GND.n4646 GND.n4645 8.92171
R15285 GND.t34 GND.n3282 8.68328
R15286 GND.n4451 GND.t61 8.68328
R15287 GND.n2032 GND.n2030 8.14595
R15288 GND.n4836 GND.n4835 8.14595
R15289 GND.n3523 GND.n3298 8.14595
R15290 GND.n4431 GND.n4393 8.14595
R15291 GND.n6340 GND.n6339 8.09206
R15292 GND.n3707 GND.n14 8.09206
R15293 GND.n3935 GND.n2235 7.95972
R15294 GND.n2808 GND.n2367 7.95972
R15295 GND.n2773 GND.n2772 7.95972
R15296 GND.n4023 GND.n2155 7.95972
R15297 GND.n4071 GND.n2111 7.95972
R15298 GND.n2488 GND.n2487 7.95972
R15299 GND.n2537 GND.n2509 7.95202
R15300 GND.t168 GND.t113 7.59793
R15301 GND.n2693 GND.t137 7.23615
R15302 GND.n6 GND.n3 7.1449
R15303 GND.t162 GND.n2242 6.87437
R15304 GND.n2684 GND.t168 6.87437
R15305 GND.t3 GND.n3038 6.51259
R15306 GND.n2339 GND.t146 6.51259
R15307 GND.n3943 GND.n2228 6.51259
R15308 GND.n2815 GND.n2359 6.51259
R15309 GND.t176 GND.n2199 6.51259
R15310 GND.n2765 GND.n2418 6.51259
R15311 GND.n4015 GND.n2163 6.51259
R15312 GND.n4047 GND.t2 6.51259
R15313 GND.n4079 GND.n2103 6.51259
R15314 GND.t58 GND.n2105 6.51259
R15315 GND.n2699 GND.n2480 6.51259
R15316 GND.t5 GND.n1757 6.51259
R15317 GND.n138 GND.n135 6.07162
R15318 GND.n13 GND.n1 5.84317
R15319 GND.t131 GND.n2257 5.78902
R15320 GND.n2200 GND.t176 5.78902
R15321 GND.n2729 GND.t2 5.78902
R15322 GND.n6 GND.n5 5.78067
R15323 GND.n9 GND.n8 5.78067
R15324 GND.n12 GND.n11 5.78067
R15325 GND.n2 GND.t13 5.69016
R15326 GND.n2 GND.t172 5.69016
R15327 GND.n4 GND.t180 5.69016
R15328 GND.n4 GND.t175 5.69016
R15329 GND.n7 GND.t155 5.69016
R15330 GND.n7 GND.t17 5.69016
R15331 GND.n10 GND.t12 5.69016
R15332 GND.n10 GND.t174 5.69016
R15333 GND.n0 GND.t154 5.69016
R15334 GND.n0 GND.t157 5.69016
R15335 GND.n134 GND.t156 5.69016
R15336 GND.n134 GND.t15 5.69016
R15337 GND.n136 GND.t173 5.69016
R15338 GND.n136 GND.t18 5.69016
R15339 GND.n139 GND.t6 5.69016
R15340 GND.n139 GND.t19 5.69016
R15341 GND.n142 GND.t179 5.69016
R15342 GND.n142 GND.t23 5.69016
R15343 GND.n145 GND.t24 5.69016
R15344 GND.n145 GND.t181 5.69016
R15345 GND.n2068 GND.t81 5.42724
R15346 GND.n2532 GND.n2509 5.23686
R15347 GND.n14 GND.n13 5.22675
R15348 GND.n6340 GND.n147 5.22675
R15349 GND.n3101 GND.t16 5.06546
R15350 GND.n2844 GND.t51 5.06546
R15351 GND.n3935 GND.t125 5.06546
R15352 GND.n2823 GND.n2822 5.06546
R15353 GND.n3951 GND.n2220 5.06546
R15354 GND.t1 GND.n2214 5.06546
R15355 GND.n4007 GND.n2170 5.06546
R15356 GND.n2758 GND.n2757 5.06546
R15357 GND.n2713 GND.t9 5.06546
R15358 GND.n2706 GND.n2473 5.06546
R15359 GND.n4087 GND.n2097 5.06546
R15360 GND.n1803 GND.t14 5.06546
R15361 GND.n2024 GND.n1926 5.04292
R15362 GND.n4842 GND.n4839 5.04292
R15363 GND.n147 GND.n146 4.7699
R15364 GND.n4520 GND.n167 4.74817
R15365 GND.n165 GND.n159 4.74817
R15366 GND.n6332 GND.n160 4.74817
R15367 GND.n168 GND.n164 4.74817
R15368 GND.n1782 GND.n167 4.74817
R15369 GND.n1798 GND.n165 4.74817
R15370 GND.n6333 GND.n6332 4.74817
R15371 GND.n4497 GND.n164 4.74817
R15372 GND.n3579 GND.n3578 4.74817
R15373 GND.n3748 GND.n3747 4.74817
R15374 GND.n3110 GND.n3089 4.74817
R15375 GND.n3732 GND.n3112 4.74817
R15376 GND.n3730 GND.n3729 4.74817
R15377 GND.n1885 GND.n1805 4.74817
R15378 GND.n4506 GND.n1887 4.74817
R15379 GND.n4504 GND.n4503 4.74817
R15380 GND.n4283 GND.n4282 4.74817
R15381 GND.n4287 GND.n4286 4.74817
R15382 GND.n1882 GND.n1805 4.74817
R15383 GND.n1887 GND.n1886 4.74817
R15384 GND.n4505 GND.n4504 4.74817
R15385 GND.n4282 GND.n1888 4.74817
R15386 GND.n4286 GND.n4285 4.74817
R15387 GND.n3759 GND.n3758 4.74817
R15388 GND.n3741 GND.n3072 4.74817
R15389 GND.n3717 GND.n3071 4.74817
R15390 GND.n3720 GND.n3070 4.74817
R15391 GND.n3759 GND.n3074 4.74817
R15392 GND.n3098 GND.n3072 4.74817
R15393 GND.n3740 GND.n3071 4.74817
R15394 GND.n3718 GND.n3070 4.74817
R15395 GND.n3578 GND.n3088 4.74817
R15396 GND.n3749 GND.n3748 4.74817
R15397 GND.n3746 GND.n3089 4.74817
R15398 GND.n3112 GND.n3111 4.74817
R15399 GND.n3731 GND.n3730 4.74817
R15400 GND.n138 GND.n137 4.7074
R15401 GND.n141 GND.n140 4.7074
R15402 GND.n144 GND.n143 4.7074
R15403 GND.n4645 GND.n1627 4.6132
R15404 GND.n1330 GND.n1327 4.6132
R15405 GND.n63 GND.n59 4.40546
R15406 GND.n43 GND.n39 4.40546
R15407 GND.n24 GND.n20 4.40546
R15408 GND.n122 GND.n118 4.40546
R15409 GND.n102 GND.n98 4.40546
R15410 GND.n83 GND.n79 4.40546
R15411 GND.n2322 GND.n2321 4.38232
R15412 GND.n2536 GND.n2535 4.38232
R15413 GND.n3165 GND.n1346 4.34189
R15414 GND.n3999 GND.t0 4.34189
R15415 GND.t8 GND.n2431 4.34189
R15416 GND.n4688 GND.n1590 4.34189
R15417 GND.n133 GND.n73 4.30175
R15418 GND.t166 GND.n2392 3.98011
R15419 GND.n4031 GND.t160 3.98011
R15420 GND.t11 GND.n3228 3.61833
R15421 GND.n2830 GND.n2346 3.61833
R15422 GND.n3959 GND.n2214 3.61833
R15423 GND.n3999 GND.n2177 3.61833
R15424 GND.n2750 GND.n2431 3.61833
R15425 GND.n2713 GND.n2466 3.61833
R15426 GND.t31 GND.n2090 3.61833
R15427 GND.n2686 GND.t74 3.61833
R15428 GND.n4471 GND.t20 3.61833
R15429 GND.n133 GND.n132 3.60163
R15430 GND.n4892 GND.n4891 3.49141
R15431 GND.n4620 GND.n4619 3.49141
R15432 GND.n6190 GND.n6187 3.49141
R15433 GND.n3452 GND.n3323 3.49141
R15434 GND.n72 GND.n54 3.49141
R15435 GND.n52 GND.n34 3.49141
R15436 GND.n33 GND.n15 3.49141
R15437 GND.n131 GND.n113 3.49141
R15438 GND.n111 GND.n93 3.49141
R15439 GND.n92 GND.n74 3.49141
R15440 GND.n4893 GND.n4892 3.10353
R15441 GND.n4621 GND.n4620 3.10353
R15442 GND.n6191 GND.n6190 3.10353
R15443 GND.n3453 GND.n3452 3.10353
R15444 GND.n70 GND.n69 2.71565
R15445 GND.n50 GND.n49 2.71565
R15446 GND.n31 GND.n30 2.71565
R15447 GND.n129 GND.n128 2.71565
R15448 GND.n109 GND.n108 2.71565
R15449 GND.n90 GND.n89 2.71565
R15450 GND.n6331 GND.n167 2.27742
R15451 GND.n6331 GND.n165 2.27742
R15452 GND.n6332 GND.n6331 2.27742
R15453 GND.n6331 GND.n164 2.27742
R15454 GND.n1805 GND.n163 2.27742
R15455 GND.n1887 GND.n163 2.27742
R15456 GND.n4504 GND.n163 2.27742
R15457 GND.n4282 GND.n163 2.27742
R15458 GND.n4286 GND.n163 2.27742
R15459 GND.n3760 GND.n3759 2.27742
R15460 GND.n3760 GND.n3072 2.27742
R15461 GND.n3760 GND.n3071 2.27742
R15462 GND.n3760 GND.n3070 2.27742
R15463 GND.n3578 GND.n3069 2.27742
R15464 GND.n3748 GND.n3069 2.27742
R15465 GND.n3089 GND.n3069 2.27742
R15466 GND.n3112 GND.n3069 2.27742
R15467 GND.n3730 GND.n3069 2.27742
R15468 GND.n2837 GND.n2339 2.1712
R15469 GND.t41 GND.n2243 2.1712
R15470 GND.n3967 GND.n2206 2.1712
R15471 GND.n3991 GND.n2184 2.1712
R15472 GND.n2743 GND.n2742 2.1712
R15473 GND.n2720 GND.n2458 2.1712
R15474 GND.n4102 GND.n2083 2.1712
R15475 GND.n66 GND.n56 1.93989
R15476 GND.n46 GND.n36 1.93989
R15477 GND.n27 GND.n17 1.93989
R15478 GND.n125 GND.n115 1.93989
R15479 GND.n105 GND.n95 1.93989
R15480 GND.n86 GND.n76 1.93989
R15481 GND.n13 GND.n12 1.90459
R15482 GND.n147 GND.n144 1.90459
R15483 GND.n2025 GND.n2024 1.55202
R15484 GND.n4843 GND.n4842 1.55202
R15485 GND.t44 GND.n2984 1.44763
R15486 GND.t27 GND.t41 1.44763
R15487 GND.t84 GND.n1694 1.44763
R15488 GND.n12 GND.n9 1.36472
R15489 GND.n144 GND.n141 1.36472
R15490 GND.n9 GND.n6 1.36257
R15491 GND.n141 GND.n138 1.36257
R15492 GND.n73 GND.n53 1.27666
R15493 GND.n132 GND.n112 1.27666
R15494 GND.n2621 GND.n2563 1.24928
R15495 GND.n2889 GND.n2888 1.24928
R15496 GND.n2907 GND.n2906 1.24928
R15497 GND.n2634 GND.n2556 1.24928
R15498 GND.n65 GND.n58 1.16414
R15499 GND.n45 GND.n38 1.16414
R15500 GND.n26 GND.n19 1.16414
R15501 GND.n124 GND.n117 1.16414
R15502 GND.n104 GND.n97 1.16414
R15503 GND.n85 GND.n78 1.16414
R15504 GND GND.n14 1.05236
R15505 GND.n2844 GND.n2332 0.724065
R15506 GND.t68 GND.n2228 0.724065
R15507 GND.n3975 GND.n2198 0.724065
R15508 GND.n3983 GND.n2192 0.724065
R15509 GND.n2735 GND.n2445 0.724065
R15510 GND.n2728 GND.n2727 0.724065
R15511 GND.n2677 GND.t48 0.724065
R15512 GND.n4110 GND.n2074 0.724065
R15513 GND.t128 GND.n2076 0.724065
R15514 GND.n2304 GND.n2302 0.716017
R15515 GND.n2530 GND.n2528 0.716017
R15516 GND.n6341 GND.n6340 0.63359
R15517 GND.n5244 GND.n5243 0.520317
R15518 GND.n5934 GND.n5933 0.520317
R15519 GND.n6074 GND.n6073 0.520317
R15520 GND.n5130 GND.n5129 0.520317
R15521 GND.n6258 GND.n6257 0.505073
R15522 GND.n1674 GND.n1600 0.505073
R15523 GND.n4950 GND.n4949 0.505073
R15524 GND.n3360 GND.n1169 0.505073
R15525 GND.n4433 GND.n4432 0.495927
R15526 GND.n3525 GND.n3524 0.495927
R15527 GND.n4822 GND.n4803 0.489829
R15528 GND.n1957 GND.n1551 0.489829
R15529 GND.n4153 GND.n4152 0.441049
R15530 GND.n3875 GND.n3874 0.441049
R15531 GND.n6331 GND.n163 0.419375
R15532 GND.n3760 GND.n3069 0.419375
R15533 GND.n62 GND.n61 0.388379
R15534 GND.n42 GND.n41 0.388379
R15535 GND.n23 GND.n22 0.388379
R15536 GND.n121 GND.n120 0.388379
R15537 GND.n101 GND.n100 0.388379
R15538 GND.n82 GND.n81 0.388379
R15539 GND.n4826 GND.n1460 0.362283
R15540 GND.n1565 GND.n1557 0.362283
R15541 GND.n2559 GND.n1625 0.312695
R15542 GND.n2898 GND.n2896 0.312695
R15543 GND.n2899 GND.n2898 0.312695
R15544 GND.n2557 GND.n1625 0.312695
R15545 GND.n6164 GND.n6163 0.299281
R15546 GND.n4593 GND.n4591 0.299281
R15547 GND.n3493 GND.n3489 0.299281
R15548 GND.n4871 GND.n4870 0.299281
R15549 GND.n6163 GND.n382 0.290134
R15550 GND.n3494 GND.n3493 0.290134
R15551 GND.n6341 GND.n133 0.279993
R15552 GND.n4154 GND.n4153 0.268793
R15553 GND.n3874 GND.n3873 0.268793
R15554 GND.n1627 GND.n1624 0.229039
R15555 GND.n1630 GND.n1627 0.229039
R15556 GND.n4918 GND.n1327 0.229039
R15557 GND.n1350 GND.n1327 0.229039
R15558 GND GND.n6341 0.211843
R15559 GND.n71 GND.n55 0.155672
R15560 GND.n64 GND.n55 0.155672
R15561 GND.n64 GND.n63 0.155672
R15562 GND.n51 GND.n35 0.155672
R15563 GND.n44 GND.n35 0.155672
R15564 GND.n44 GND.n43 0.155672
R15565 GND.n32 GND.n16 0.155672
R15566 GND.n25 GND.n16 0.155672
R15567 GND.n25 GND.n24 0.155672
R15568 GND.n130 GND.n114 0.155672
R15569 GND.n123 GND.n114 0.155672
R15570 GND.n123 GND.n122 0.155672
R15571 GND.n110 GND.n94 0.155672
R15572 GND.n103 GND.n94 0.155672
R15573 GND.n103 GND.n102 0.155672
R15574 GND.n91 GND.n75 0.155672
R15575 GND.n84 GND.n75 0.155672
R15576 GND.n84 GND.n83 0.155672
R15577 GND.n5245 GND.n5244 0.152939
R15578 GND.n5245 GND.n964 0.152939
R15579 GND.n5253 GND.n964 0.152939
R15580 GND.n5254 GND.n5253 0.152939
R15581 GND.n5255 GND.n5254 0.152939
R15582 GND.n5255 GND.n958 0.152939
R15583 GND.n5263 GND.n958 0.152939
R15584 GND.n5264 GND.n5263 0.152939
R15585 GND.n5265 GND.n5264 0.152939
R15586 GND.n5265 GND.n952 0.152939
R15587 GND.n5273 GND.n952 0.152939
R15588 GND.n5274 GND.n5273 0.152939
R15589 GND.n5275 GND.n5274 0.152939
R15590 GND.n5275 GND.n946 0.152939
R15591 GND.n5283 GND.n946 0.152939
R15592 GND.n5284 GND.n5283 0.152939
R15593 GND.n5285 GND.n5284 0.152939
R15594 GND.n5285 GND.n940 0.152939
R15595 GND.n5293 GND.n940 0.152939
R15596 GND.n5294 GND.n5293 0.152939
R15597 GND.n5295 GND.n5294 0.152939
R15598 GND.n5295 GND.n934 0.152939
R15599 GND.n5303 GND.n934 0.152939
R15600 GND.n5304 GND.n5303 0.152939
R15601 GND.n5305 GND.n5304 0.152939
R15602 GND.n5305 GND.n928 0.152939
R15603 GND.n5313 GND.n928 0.152939
R15604 GND.n5314 GND.n5313 0.152939
R15605 GND.n5315 GND.n5314 0.152939
R15606 GND.n5315 GND.n922 0.152939
R15607 GND.n5323 GND.n922 0.152939
R15608 GND.n5324 GND.n5323 0.152939
R15609 GND.n5325 GND.n5324 0.152939
R15610 GND.n5325 GND.n916 0.152939
R15611 GND.n5333 GND.n916 0.152939
R15612 GND.n5334 GND.n5333 0.152939
R15613 GND.n5335 GND.n5334 0.152939
R15614 GND.n5335 GND.n910 0.152939
R15615 GND.n5343 GND.n910 0.152939
R15616 GND.n5344 GND.n5343 0.152939
R15617 GND.n5345 GND.n5344 0.152939
R15618 GND.n5345 GND.n904 0.152939
R15619 GND.n5353 GND.n904 0.152939
R15620 GND.n5354 GND.n5353 0.152939
R15621 GND.n5355 GND.n5354 0.152939
R15622 GND.n5355 GND.n898 0.152939
R15623 GND.n5363 GND.n898 0.152939
R15624 GND.n5364 GND.n5363 0.152939
R15625 GND.n5365 GND.n5364 0.152939
R15626 GND.n5365 GND.n892 0.152939
R15627 GND.n5373 GND.n892 0.152939
R15628 GND.n5374 GND.n5373 0.152939
R15629 GND.n5375 GND.n5374 0.152939
R15630 GND.n5375 GND.n886 0.152939
R15631 GND.n5383 GND.n886 0.152939
R15632 GND.n5384 GND.n5383 0.152939
R15633 GND.n5385 GND.n5384 0.152939
R15634 GND.n5385 GND.n880 0.152939
R15635 GND.n5393 GND.n880 0.152939
R15636 GND.n5394 GND.n5393 0.152939
R15637 GND.n5395 GND.n5394 0.152939
R15638 GND.n5395 GND.n874 0.152939
R15639 GND.n5403 GND.n874 0.152939
R15640 GND.n5404 GND.n5403 0.152939
R15641 GND.n5405 GND.n5404 0.152939
R15642 GND.n5405 GND.n868 0.152939
R15643 GND.n5413 GND.n868 0.152939
R15644 GND.n5414 GND.n5413 0.152939
R15645 GND.n5415 GND.n5414 0.152939
R15646 GND.n5415 GND.n862 0.152939
R15647 GND.n5423 GND.n862 0.152939
R15648 GND.n5424 GND.n5423 0.152939
R15649 GND.n5425 GND.n5424 0.152939
R15650 GND.n5425 GND.n856 0.152939
R15651 GND.n5433 GND.n856 0.152939
R15652 GND.n5434 GND.n5433 0.152939
R15653 GND.n5435 GND.n5434 0.152939
R15654 GND.n5435 GND.n850 0.152939
R15655 GND.n5443 GND.n850 0.152939
R15656 GND.n5444 GND.n5443 0.152939
R15657 GND.n5445 GND.n5444 0.152939
R15658 GND.n5445 GND.n844 0.152939
R15659 GND.n5453 GND.n844 0.152939
R15660 GND.n5454 GND.n5453 0.152939
R15661 GND.n5455 GND.n5454 0.152939
R15662 GND.n5455 GND.n838 0.152939
R15663 GND.n5463 GND.n838 0.152939
R15664 GND.n5464 GND.n5463 0.152939
R15665 GND.n5465 GND.n5464 0.152939
R15666 GND.n5465 GND.n832 0.152939
R15667 GND.n5473 GND.n832 0.152939
R15668 GND.n5474 GND.n5473 0.152939
R15669 GND.n5475 GND.n5474 0.152939
R15670 GND.n5475 GND.n826 0.152939
R15671 GND.n5483 GND.n826 0.152939
R15672 GND.n5484 GND.n5483 0.152939
R15673 GND.n5485 GND.n5484 0.152939
R15674 GND.n5485 GND.n820 0.152939
R15675 GND.n5493 GND.n820 0.152939
R15676 GND.n5494 GND.n5493 0.152939
R15677 GND.n5495 GND.n5494 0.152939
R15678 GND.n5495 GND.n814 0.152939
R15679 GND.n5503 GND.n814 0.152939
R15680 GND.n5504 GND.n5503 0.152939
R15681 GND.n5505 GND.n5504 0.152939
R15682 GND.n5505 GND.n808 0.152939
R15683 GND.n5513 GND.n808 0.152939
R15684 GND.n5514 GND.n5513 0.152939
R15685 GND.n5515 GND.n5514 0.152939
R15686 GND.n5515 GND.n802 0.152939
R15687 GND.n5523 GND.n802 0.152939
R15688 GND.n5524 GND.n5523 0.152939
R15689 GND.n5525 GND.n5524 0.152939
R15690 GND.n5525 GND.n796 0.152939
R15691 GND.n5533 GND.n796 0.152939
R15692 GND.n5534 GND.n5533 0.152939
R15693 GND.n5535 GND.n5534 0.152939
R15694 GND.n5535 GND.n790 0.152939
R15695 GND.n5543 GND.n790 0.152939
R15696 GND.n5544 GND.n5543 0.152939
R15697 GND.n5545 GND.n5544 0.152939
R15698 GND.n5545 GND.n784 0.152939
R15699 GND.n5553 GND.n784 0.152939
R15700 GND.n5554 GND.n5553 0.152939
R15701 GND.n5555 GND.n5554 0.152939
R15702 GND.n5555 GND.n778 0.152939
R15703 GND.n5563 GND.n778 0.152939
R15704 GND.n5564 GND.n5563 0.152939
R15705 GND.n5565 GND.n5564 0.152939
R15706 GND.n5565 GND.n772 0.152939
R15707 GND.n5573 GND.n772 0.152939
R15708 GND.n5574 GND.n5573 0.152939
R15709 GND.n5575 GND.n5574 0.152939
R15710 GND.n5575 GND.n766 0.152939
R15711 GND.n5583 GND.n766 0.152939
R15712 GND.n5584 GND.n5583 0.152939
R15713 GND.n5585 GND.n5584 0.152939
R15714 GND.n5585 GND.n760 0.152939
R15715 GND.n5593 GND.n760 0.152939
R15716 GND.n5594 GND.n5593 0.152939
R15717 GND.n5595 GND.n5594 0.152939
R15718 GND.n5595 GND.n754 0.152939
R15719 GND.n5603 GND.n754 0.152939
R15720 GND.n5604 GND.n5603 0.152939
R15721 GND.n5605 GND.n5604 0.152939
R15722 GND.n5605 GND.n748 0.152939
R15723 GND.n5613 GND.n748 0.152939
R15724 GND.n5614 GND.n5613 0.152939
R15725 GND.n5615 GND.n5614 0.152939
R15726 GND.n5615 GND.n742 0.152939
R15727 GND.n5623 GND.n742 0.152939
R15728 GND.n5624 GND.n5623 0.152939
R15729 GND.n5625 GND.n5624 0.152939
R15730 GND.n5625 GND.n736 0.152939
R15731 GND.n5633 GND.n736 0.152939
R15732 GND.n5634 GND.n5633 0.152939
R15733 GND.n5635 GND.n5634 0.152939
R15734 GND.n5635 GND.n730 0.152939
R15735 GND.n5643 GND.n730 0.152939
R15736 GND.n5644 GND.n5643 0.152939
R15737 GND.n5645 GND.n5644 0.152939
R15738 GND.n5645 GND.n724 0.152939
R15739 GND.n5653 GND.n724 0.152939
R15740 GND.n5654 GND.n5653 0.152939
R15741 GND.n5655 GND.n5654 0.152939
R15742 GND.n5655 GND.n718 0.152939
R15743 GND.n5663 GND.n718 0.152939
R15744 GND.n5664 GND.n5663 0.152939
R15745 GND.n5665 GND.n5664 0.152939
R15746 GND.n5665 GND.n712 0.152939
R15747 GND.n5673 GND.n712 0.152939
R15748 GND.n5674 GND.n5673 0.152939
R15749 GND.n5675 GND.n5674 0.152939
R15750 GND.n5675 GND.n706 0.152939
R15751 GND.n5683 GND.n706 0.152939
R15752 GND.n5684 GND.n5683 0.152939
R15753 GND.n5685 GND.n5684 0.152939
R15754 GND.n5685 GND.n700 0.152939
R15755 GND.n5693 GND.n700 0.152939
R15756 GND.n5694 GND.n5693 0.152939
R15757 GND.n5695 GND.n5694 0.152939
R15758 GND.n5695 GND.n694 0.152939
R15759 GND.n5703 GND.n694 0.152939
R15760 GND.n5704 GND.n5703 0.152939
R15761 GND.n5705 GND.n5704 0.152939
R15762 GND.n5705 GND.n688 0.152939
R15763 GND.n5713 GND.n688 0.152939
R15764 GND.n5714 GND.n5713 0.152939
R15765 GND.n5715 GND.n5714 0.152939
R15766 GND.n5715 GND.n682 0.152939
R15767 GND.n5723 GND.n682 0.152939
R15768 GND.n5724 GND.n5723 0.152939
R15769 GND.n5725 GND.n5724 0.152939
R15770 GND.n5725 GND.n676 0.152939
R15771 GND.n5733 GND.n676 0.152939
R15772 GND.n5734 GND.n5733 0.152939
R15773 GND.n5735 GND.n5734 0.152939
R15774 GND.n5735 GND.n670 0.152939
R15775 GND.n5743 GND.n670 0.152939
R15776 GND.n5744 GND.n5743 0.152939
R15777 GND.n5745 GND.n5744 0.152939
R15778 GND.n5745 GND.n664 0.152939
R15779 GND.n5753 GND.n664 0.152939
R15780 GND.n5754 GND.n5753 0.152939
R15781 GND.n5755 GND.n5754 0.152939
R15782 GND.n5755 GND.n658 0.152939
R15783 GND.n5763 GND.n658 0.152939
R15784 GND.n5764 GND.n5763 0.152939
R15785 GND.n5765 GND.n5764 0.152939
R15786 GND.n5765 GND.n652 0.152939
R15787 GND.n5773 GND.n652 0.152939
R15788 GND.n5774 GND.n5773 0.152939
R15789 GND.n5775 GND.n5774 0.152939
R15790 GND.n5775 GND.n646 0.152939
R15791 GND.n5783 GND.n646 0.152939
R15792 GND.n5784 GND.n5783 0.152939
R15793 GND.n5785 GND.n5784 0.152939
R15794 GND.n5785 GND.n640 0.152939
R15795 GND.n5793 GND.n640 0.152939
R15796 GND.n5794 GND.n5793 0.152939
R15797 GND.n5795 GND.n5794 0.152939
R15798 GND.n5795 GND.n634 0.152939
R15799 GND.n5803 GND.n634 0.152939
R15800 GND.n5804 GND.n5803 0.152939
R15801 GND.n5805 GND.n5804 0.152939
R15802 GND.n5805 GND.n628 0.152939
R15803 GND.n5813 GND.n628 0.152939
R15804 GND.n5814 GND.n5813 0.152939
R15805 GND.n5815 GND.n5814 0.152939
R15806 GND.n5815 GND.n622 0.152939
R15807 GND.n5823 GND.n622 0.152939
R15808 GND.n5824 GND.n5823 0.152939
R15809 GND.n5825 GND.n5824 0.152939
R15810 GND.n5825 GND.n616 0.152939
R15811 GND.n5833 GND.n616 0.152939
R15812 GND.n5834 GND.n5833 0.152939
R15813 GND.n5835 GND.n5834 0.152939
R15814 GND.n5835 GND.n610 0.152939
R15815 GND.n5843 GND.n610 0.152939
R15816 GND.n5844 GND.n5843 0.152939
R15817 GND.n5845 GND.n5844 0.152939
R15818 GND.n5845 GND.n604 0.152939
R15819 GND.n5853 GND.n604 0.152939
R15820 GND.n5854 GND.n5853 0.152939
R15821 GND.n5855 GND.n5854 0.152939
R15822 GND.n5855 GND.n598 0.152939
R15823 GND.n5863 GND.n598 0.152939
R15824 GND.n5864 GND.n5863 0.152939
R15825 GND.n5865 GND.n5864 0.152939
R15826 GND.n5865 GND.n592 0.152939
R15827 GND.n5873 GND.n592 0.152939
R15828 GND.n5874 GND.n5873 0.152939
R15829 GND.n5875 GND.n5874 0.152939
R15830 GND.n5875 GND.n586 0.152939
R15831 GND.n5883 GND.n586 0.152939
R15832 GND.n5884 GND.n5883 0.152939
R15833 GND.n5885 GND.n5884 0.152939
R15834 GND.n5885 GND.n580 0.152939
R15835 GND.n5893 GND.n580 0.152939
R15836 GND.n5894 GND.n5893 0.152939
R15837 GND.n5895 GND.n5894 0.152939
R15838 GND.n5895 GND.n574 0.152939
R15839 GND.n5903 GND.n574 0.152939
R15840 GND.n5904 GND.n5903 0.152939
R15841 GND.n5905 GND.n5904 0.152939
R15842 GND.n5905 GND.n568 0.152939
R15843 GND.n5913 GND.n568 0.152939
R15844 GND.n5914 GND.n5913 0.152939
R15845 GND.n5915 GND.n5914 0.152939
R15846 GND.n5915 GND.n562 0.152939
R15847 GND.n5923 GND.n562 0.152939
R15848 GND.n5924 GND.n5923 0.152939
R15849 GND.n5925 GND.n5924 0.152939
R15850 GND.n5925 GND.n556 0.152939
R15851 GND.n5933 GND.n556 0.152939
R15852 GND.n5935 GND.n5934 0.152939
R15853 GND.n5935 GND.n550 0.152939
R15854 GND.n5943 GND.n550 0.152939
R15855 GND.n5944 GND.n5943 0.152939
R15856 GND.n5945 GND.n5944 0.152939
R15857 GND.n5945 GND.n544 0.152939
R15858 GND.n5953 GND.n544 0.152939
R15859 GND.n5954 GND.n5953 0.152939
R15860 GND.n5955 GND.n5954 0.152939
R15861 GND.n5955 GND.n538 0.152939
R15862 GND.n5963 GND.n538 0.152939
R15863 GND.n5964 GND.n5963 0.152939
R15864 GND.n5965 GND.n5964 0.152939
R15865 GND.n5965 GND.n532 0.152939
R15866 GND.n5973 GND.n532 0.152939
R15867 GND.n5974 GND.n5973 0.152939
R15868 GND.n5975 GND.n5974 0.152939
R15869 GND.n5975 GND.n526 0.152939
R15870 GND.n5983 GND.n526 0.152939
R15871 GND.n5984 GND.n5983 0.152939
R15872 GND.n5985 GND.n5984 0.152939
R15873 GND.n5985 GND.n520 0.152939
R15874 GND.n5993 GND.n520 0.152939
R15875 GND.n5994 GND.n5993 0.152939
R15876 GND.n5995 GND.n5994 0.152939
R15877 GND.n5995 GND.n514 0.152939
R15878 GND.n6003 GND.n514 0.152939
R15879 GND.n6004 GND.n6003 0.152939
R15880 GND.n6005 GND.n6004 0.152939
R15881 GND.n6005 GND.n508 0.152939
R15882 GND.n6013 GND.n508 0.152939
R15883 GND.n6014 GND.n6013 0.152939
R15884 GND.n6015 GND.n6014 0.152939
R15885 GND.n6015 GND.n502 0.152939
R15886 GND.n6023 GND.n502 0.152939
R15887 GND.n6024 GND.n6023 0.152939
R15888 GND.n6025 GND.n6024 0.152939
R15889 GND.n6025 GND.n496 0.152939
R15890 GND.n6033 GND.n496 0.152939
R15891 GND.n6034 GND.n6033 0.152939
R15892 GND.n6035 GND.n6034 0.152939
R15893 GND.n6035 GND.n490 0.152939
R15894 GND.n6043 GND.n490 0.152939
R15895 GND.n6044 GND.n6043 0.152939
R15896 GND.n6045 GND.n6044 0.152939
R15897 GND.n6045 GND.n484 0.152939
R15898 GND.n6053 GND.n484 0.152939
R15899 GND.n6054 GND.n6053 0.152939
R15900 GND.n6055 GND.n6054 0.152939
R15901 GND.n6055 GND.n478 0.152939
R15902 GND.n6063 GND.n478 0.152939
R15903 GND.n6064 GND.n6063 0.152939
R15904 GND.n6065 GND.n6064 0.152939
R15905 GND.n6065 GND.n472 0.152939
R15906 GND.n6073 GND.n472 0.152939
R15907 GND.n4288 GND.n4279 0.152939
R15908 GND.n4294 GND.n4279 0.152939
R15909 GND.n4295 GND.n4294 0.152939
R15910 GND.n4296 GND.n4295 0.152939
R15911 GND.n4297 GND.n4296 0.152939
R15912 GND.n4298 GND.n4297 0.152939
R15913 GND.n4301 GND.n4298 0.152939
R15914 GND.n4302 GND.n4301 0.152939
R15915 GND.n4303 GND.n4302 0.152939
R15916 GND.n4304 GND.n4303 0.152939
R15917 GND.n4307 GND.n4304 0.152939
R15918 GND.n4308 GND.n4307 0.152939
R15919 GND.n4309 GND.n4308 0.152939
R15920 GND.n4310 GND.n4309 0.152939
R15921 GND.n4313 GND.n4310 0.152939
R15922 GND.n4314 GND.n4313 0.152939
R15923 GND.n4315 GND.n4314 0.152939
R15924 GND.n4316 GND.n4315 0.152939
R15925 GND.n4318 GND.n4316 0.152939
R15926 GND.n4320 GND.n4318 0.152939
R15927 GND.n4320 GND.n4319 0.152939
R15928 GND.n4319 GND.n391 0.152939
R15929 GND.n392 GND.n391 0.152939
R15930 GND.n393 GND.n392 0.152939
R15931 GND.n398 GND.n393 0.152939
R15932 GND.n399 GND.n398 0.152939
R15933 GND.n400 GND.n399 0.152939
R15934 GND.n401 GND.n400 0.152939
R15935 GND.n406 GND.n401 0.152939
R15936 GND.n407 GND.n406 0.152939
R15937 GND.n408 GND.n407 0.152939
R15938 GND.n409 GND.n408 0.152939
R15939 GND.n414 GND.n409 0.152939
R15940 GND.n415 GND.n414 0.152939
R15941 GND.n416 GND.n415 0.152939
R15942 GND.n417 GND.n416 0.152939
R15943 GND.n422 GND.n417 0.152939
R15944 GND.n423 GND.n422 0.152939
R15945 GND.n424 GND.n423 0.152939
R15946 GND.n425 GND.n424 0.152939
R15947 GND.n430 GND.n425 0.152939
R15948 GND.n431 GND.n430 0.152939
R15949 GND.n432 GND.n431 0.152939
R15950 GND.n433 GND.n432 0.152939
R15951 GND.n438 GND.n433 0.152939
R15952 GND.n439 GND.n438 0.152939
R15953 GND.n440 GND.n439 0.152939
R15954 GND.n441 GND.n440 0.152939
R15955 GND.n446 GND.n441 0.152939
R15956 GND.n447 GND.n446 0.152939
R15957 GND.n448 GND.n447 0.152939
R15958 GND.n449 GND.n448 0.152939
R15959 GND.n454 GND.n449 0.152939
R15960 GND.n455 GND.n454 0.152939
R15961 GND.n456 GND.n455 0.152939
R15962 GND.n457 GND.n456 0.152939
R15963 GND.n462 GND.n457 0.152939
R15964 GND.n463 GND.n462 0.152939
R15965 GND.n464 GND.n463 0.152939
R15966 GND.n465 GND.n464 0.152939
R15967 GND.n470 GND.n465 0.152939
R15968 GND.n471 GND.n470 0.152939
R15969 GND.n6074 GND.n471 0.152939
R15970 GND.n189 GND.n161 0.152939
R15971 GND.n190 GND.n189 0.152939
R15972 GND.n191 GND.n190 0.152939
R15973 GND.n208 GND.n191 0.152939
R15974 GND.n209 GND.n208 0.152939
R15975 GND.n210 GND.n209 0.152939
R15976 GND.n211 GND.n210 0.152939
R15977 GND.n229 GND.n211 0.152939
R15978 GND.n230 GND.n229 0.152939
R15979 GND.n231 GND.n230 0.152939
R15980 GND.n232 GND.n231 0.152939
R15981 GND.n250 GND.n232 0.152939
R15982 GND.n251 GND.n250 0.152939
R15983 GND.n252 GND.n251 0.152939
R15984 GND.n253 GND.n252 0.152939
R15985 GND.n270 GND.n253 0.152939
R15986 GND.n271 GND.n270 0.152939
R15987 GND.n272 GND.n271 0.152939
R15988 GND.n273 GND.n272 0.152939
R15989 GND.n291 GND.n273 0.152939
R15990 GND.n292 GND.n291 0.152939
R15991 GND.n6258 GND.n292 0.152939
R15992 GND.n4154 GND.n1922 0.152939
R15993 GND.n4163 GND.n1922 0.152939
R15994 GND.n4164 GND.n4163 0.152939
R15995 GND.n4165 GND.n4164 0.152939
R15996 GND.n4165 GND.n1918 0.152939
R15997 GND.n4178 GND.n1918 0.152939
R15998 GND.n4179 GND.n4178 0.152939
R15999 GND.n4180 GND.n4179 0.152939
R16000 GND.n4180 GND.n1914 0.152939
R16001 GND.n4193 GND.n1914 0.152939
R16002 GND.n4194 GND.n4193 0.152939
R16003 GND.n4195 GND.n4194 0.152939
R16004 GND.n4195 GND.n1910 0.152939
R16005 GND.n4208 GND.n1910 0.152939
R16006 GND.n4209 GND.n4208 0.152939
R16007 GND.n4210 GND.n4209 0.152939
R16008 GND.n4210 GND.n1906 0.152939
R16009 GND.n4223 GND.n1906 0.152939
R16010 GND.n4224 GND.n4223 0.152939
R16011 GND.n4225 GND.n4224 0.152939
R16012 GND.n4225 GND.n1902 0.152939
R16013 GND.n4238 GND.n1902 0.152939
R16014 GND.n4239 GND.n4238 0.152939
R16015 GND.n4240 GND.n4239 0.152939
R16016 GND.n4241 GND.n4240 0.152939
R16017 GND.n4242 GND.n4241 0.152939
R16018 GND.n4242 GND.n148 0.152939
R16019 GND.n6338 GND.n149 0.152939
R16020 GND.n4263 GND.n149 0.152939
R16021 GND.n4264 GND.n4263 0.152939
R16022 GND.n4265 GND.n4264 0.152939
R16023 GND.n4266 GND.n4265 0.152939
R16024 GND.n4270 GND.n4266 0.152939
R16025 GND.n4271 GND.n4270 0.152939
R16026 GND.n4272 GND.n4271 0.152939
R16027 GND.n4273 GND.n4272 0.152939
R16028 GND.n4347 GND.n4273 0.152939
R16029 GND.n4348 GND.n4347 0.152939
R16030 GND.n4348 GND.n4342 0.152939
R16031 GND.n4360 GND.n4342 0.152939
R16032 GND.n4361 GND.n4360 0.152939
R16033 GND.n4362 GND.n4361 0.152939
R16034 GND.n4362 GND.n4337 0.152939
R16035 GND.n4374 GND.n4337 0.152939
R16036 GND.n4375 GND.n4374 0.152939
R16037 GND.n4377 GND.n4375 0.152939
R16038 GND.n4377 GND.n4376 0.152939
R16039 GND.n4376 GND.n4330 0.152939
R16040 GND.n4331 GND.n4330 0.152939
R16041 GND.n4332 GND.n4331 0.152939
R16042 GND.n4387 GND.n4332 0.152939
R16043 GND.n4388 GND.n4387 0.152939
R16044 GND.n4389 GND.n4388 0.152939
R16045 GND.n4433 GND.n4389 0.152939
R16046 GND.n4405 GND.n382 0.152939
R16047 GND.n4405 GND.n4400 0.152939
R16048 GND.n4413 GND.n4400 0.152939
R16049 GND.n4414 GND.n4413 0.152939
R16050 GND.n4415 GND.n4414 0.152939
R16051 GND.n4415 GND.n4396 0.152939
R16052 GND.n4423 GND.n4396 0.152939
R16053 GND.n4424 GND.n4423 0.152939
R16054 GND.n4425 GND.n4424 0.152939
R16055 GND.n4425 GND.n4390 0.152939
R16056 GND.n4432 GND.n4390 0.152939
R16057 GND.n6257 GND.n293 0.152939
R16058 GND.n298 GND.n293 0.152939
R16059 GND.n299 GND.n298 0.152939
R16060 GND.n300 GND.n299 0.152939
R16061 GND.n301 GND.n300 0.152939
R16062 GND.n305 GND.n301 0.152939
R16063 GND.n306 GND.n305 0.152939
R16064 GND.n307 GND.n306 0.152939
R16065 GND.n308 GND.n307 0.152939
R16066 GND.n314 GND.n308 0.152939
R16067 GND.n315 GND.n314 0.152939
R16068 GND.n316 GND.n315 0.152939
R16069 GND.n317 GND.n316 0.152939
R16070 GND.n321 GND.n317 0.152939
R16071 GND.n322 GND.n321 0.152939
R16072 GND.n323 GND.n322 0.152939
R16073 GND.n324 GND.n323 0.152939
R16074 GND.n328 GND.n324 0.152939
R16075 GND.n329 GND.n328 0.152939
R16076 GND.n330 GND.n329 0.152939
R16077 GND.n331 GND.n330 0.152939
R16078 GND.n338 GND.n331 0.152939
R16079 GND.n6213 GND.n338 0.152939
R16080 GND.n6213 GND.n6212 0.152939
R16081 GND.n6212 GND.n6211 0.152939
R16082 GND.n6211 GND.n339 0.152939
R16083 GND.n343 GND.n339 0.152939
R16084 GND.n344 GND.n343 0.152939
R16085 GND.n345 GND.n344 0.152939
R16086 GND.n349 GND.n345 0.152939
R16087 GND.n350 GND.n349 0.152939
R16088 GND.n351 GND.n350 0.152939
R16089 GND.n352 GND.n351 0.152939
R16090 GND.n356 GND.n352 0.152939
R16091 GND.n357 GND.n356 0.152939
R16092 GND.n358 GND.n357 0.152939
R16093 GND.n359 GND.n358 0.152939
R16094 GND.n363 GND.n359 0.152939
R16095 GND.n364 GND.n363 0.152939
R16096 GND.n365 GND.n364 0.152939
R16097 GND.n366 GND.n365 0.152939
R16098 GND.n370 GND.n366 0.152939
R16099 GND.n371 GND.n370 0.152939
R16100 GND.n372 GND.n371 0.152939
R16101 GND.n373 GND.n372 0.152939
R16102 GND.n377 GND.n373 0.152939
R16103 GND.n378 GND.n377 0.152939
R16104 GND.n6165 GND.n378 0.152939
R16105 GND.n6165 GND.n6164 0.152939
R16106 GND.n1601 GND.n1600 0.152939
R16107 GND.n1602 GND.n1601 0.152939
R16108 GND.n1603 GND.n1602 0.152939
R16109 GND.n1604 GND.n1603 0.152939
R16110 GND.n1605 GND.n1604 0.152939
R16111 GND.n1606 GND.n1605 0.152939
R16112 GND.n1607 GND.n1606 0.152939
R16113 GND.n1608 GND.n1607 0.152939
R16114 GND.n1609 GND.n1608 0.152939
R16115 GND.n1611 GND.n1609 0.152939
R16116 GND.n1614 GND.n1611 0.152939
R16117 GND.n1615 GND.n1614 0.152939
R16118 GND.n1616 GND.n1615 0.152939
R16119 GND.n1617 GND.n1616 0.152939
R16120 GND.n1618 GND.n1617 0.152939
R16121 GND.n1619 GND.n1618 0.152939
R16122 GND.n1620 GND.n1619 0.152939
R16123 GND.n1621 GND.n1620 0.152939
R16124 GND.n1622 GND.n1621 0.152939
R16125 GND.n1623 GND.n1622 0.152939
R16126 GND.n1624 GND.n1623 0.152939
R16127 GND.n1631 GND.n1630 0.152939
R16128 GND.n1632 GND.n1631 0.152939
R16129 GND.n1633 GND.n1632 0.152939
R16130 GND.n1634 GND.n1633 0.152939
R16131 GND.n1635 GND.n1634 0.152939
R16132 GND.n1636 GND.n1635 0.152939
R16133 GND.n1637 GND.n1636 0.152939
R16134 GND.n1638 GND.n1637 0.152939
R16135 GND.n1639 GND.n1638 0.152939
R16136 GND.n1640 GND.n1639 0.152939
R16137 GND.n1641 GND.n1640 0.152939
R16138 GND.n1644 GND.n1641 0.152939
R16139 GND.n1645 GND.n1644 0.152939
R16140 GND.n1646 GND.n1645 0.152939
R16141 GND.n1647 GND.n1646 0.152939
R16142 GND.n1648 GND.n1647 0.152939
R16143 GND.n1649 GND.n1648 0.152939
R16144 GND.n1650 GND.n1649 0.152939
R16145 GND.n1651 GND.n1650 0.152939
R16146 GND.n1652 GND.n1651 0.152939
R16147 GND.n1653 GND.n1652 0.152939
R16148 GND.n1654 GND.n1653 0.152939
R16149 GND.n4595 GND.n1654 0.152939
R16150 GND.n4595 GND.n4594 0.152939
R16151 GND.n4594 GND.n4593 0.152939
R16152 GND.n1675 GND.n1674 0.152939
R16153 GND.n1676 GND.n1675 0.152939
R16154 GND.n1677 GND.n1676 0.152939
R16155 GND.n1696 GND.n1677 0.152939
R16156 GND.n1697 GND.n1696 0.152939
R16157 GND.n1698 GND.n1697 0.152939
R16158 GND.n1699 GND.n1698 0.152939
R16159 GND.n1717 GND.n1699 0.152939
R16160 GND.n1718 GND.n1717 0.152939
R16161 GND.n1719 GND.n1718 0.152939
R16162 GND.n1720 GND.n1719 0.152939
R16163 GND.n1738 GND.n1720 0.152939
R16164 GND.n1739 GND.n1738 0.152939
R16165 GND.n1740 GND.n1739 0.152939
R16166 GND.n1741 GND.n1740 0.152939
R16167 GND.n1759 GND.n1741 0.152939
R16168 GND.n1760 GND.n1759 0.152939
R16169 GND.n1761 GND.n1760 0.152939
R16170 GND.n1762 GND.n1761 0.152939
R16171 GND.n1780 GND.n1762 0.152939
R16172 GND.n1781 GND.n1780 0.152939
R16173 GND.n1781 GND.n162 0.152939
R16174 GND.n3116 GND.n3115 0.152939
R16175 GND.n3117 GND.n3116 0.152939
R16176 GND.n3118 GND.n3117 0.152939
R16177 GND.n3121 GND.n3118 0.152939
R16178 GND.n3122 GND.n3121 0.152939
R16179 GND.n3123 GND.n3122 0.152939
R16180 GND.n3124 GND.n3123 0.152939
R16181 GND.n3127 GND.n3124 0.152939
R16182 GND.n3128 GND.n3127 0.152939
R16183 GND.n3129 GND.n3128 0.152939
R16184 GND.n3130 GND.n3129 0.152939
R16185 GND.n3133 GND.n3130 0.152939
R16186 GND.n3134 GND.n3133 0.152939
R16187 GND.n3135 GND.n3134 0.152939
R16188 GND.n3136 GND.n3135 0.152939
R16189 GND.n3139 GND.n3136 0.152939
R16190 GND.n3140 GND.n3139 0.152939
R16191 GND.n3141 GND.n3140 0.152939
R16192 GND.n3142 GND.n3141 0.152939
R16193 GND.n3145 GND.n3142 0.152939
R16194 GND.n3146 GND.n3145 0.152939
R16195 GND.n3147 GND.n3146 0.152939
R16196 GND.n3148 GND.n3147 0.152939
R16197 GND.n3151 GND.n3148 0.152939
R16198 GND.n3152 GND.n3151 0.152939
R16199 GND.n3153 GND.n3152 0.152939
R16200 GND.n3154 GND.n3153 0.152939
R16201 GND.n3155 GND.n3154 0.152939
R16202 GND.n3155 GND.n2963 0.152939
R16203 GND.n3882 GND.n2963 0.152939
R16204 GND.n3883 GND.n3882 0.152939
R16205 GND.n3884 GND.n3883 0.152939
R16206 GND.n3884 GND.n2950 0.152939
R16207 GND.n3898 GND.n2950 0.152939
R16208 GND.n3899 GND.n3898 0.152939
R16209 GND.n3900 GND.n3899 0.152939
R16210 GND.n3900 GND.n2254 0.152939
R16211 GND.n3914 GND.n2254 0.152939
R16212 GND.n3915 GND.n3914 0.152939
R16213 GND.n3916 GND.n3915 0.152939
R16214 GND.n3916 GND.n2239 0.152939
R16215 GND.n3930 GND.n2239 0.152939
R16216 GND.n3931 GND.n3930 0.152939
R16217 GND.n3932 GND.n3931 0.152939
R16218 GND.n3932 GND.n2225 0.152939
R16219 GND.n3946 GND.n2225 0.152939
R16220 GND.n3947 GND.n3946 0.152939
R16221 GND.n3948 GND.n3947 0.152939
R16222 GND.n3948 GND.n2211 0.152939
R16223 GND.n3962 GND.n2211 0.152939
R16224 GND.n3963 GND.n3962 0.152939
R16225 GND.n3964 GND.n3963 0.152939
R16226 GND.n3964 GND.n2195 0.152939
R16227 GND.n3978 GND.n2195 0.152939
R16228 GND.n3979 GND.n3978 0.152939
R16229 GND.n3980 GND.n3979 0.152939
R16230 GND.n3980 GND.n2180 0.152939
R16231 GND.n3994 GND.n2180 0.152939
R16232 GND.n3995 GND.n3994 0.152939
R16233 GND.n3996 GND.n3995 0.152939
R16234 GND.n3996 GND.n2166 0.152939
R16235 GND.n4010 GND.n2166 0.152939
R16236 GND.n4011 GND.n4010 0.152939
R16237 GND.n4012 GND.n4011 0.152939
R16238 GND.n4012 GND.n2151 0.152939
R16239 GND.n4026 GND.n2151 0.152939
R16240 GND.n4027 GND.n4026 0.152939
R16241 GND.n4028 GND.n4027 0.152939
R16242 GND.n4028 GND.n2137 0.152939
R16243 GND.n4042 GND.n2137 0.152939
R16244 GND.n4043 GND.n4042 0.152939
R16245 GND.n4044 GND.n4043 0.152939
R16246 GND.n4044 GND.n2123 0.152939
R16247 GND.n4058 GND.n2123 0.152939
R16248 GND.n4059 GND.n4058 0.152939
R16249 GND.n4060 GND.n4059 0.152939
R16250 GND.n4060 GND.n2108 0.152939
R16251 GND.n4074 GND.n2108 0.152939
R16252 GND.n4075 GND.n4074 0.152939
R16253 GND.n4076 GND.n4075 0.152939
R16254 GND.n4076 GND.n2094 0.152939
R16255 GND.n4090 GND.n2094 0.152939
R16256 GND.n4091 GND.n4090 0.152939
R16257 GND.n4092 GND.n4091 0.152939
R16258 GND.n4092 GND.n2080 0.152939
R16259 GND.n4105 GND.n2080 0.152939
R16260 GND.n4106 GND.n4105 0.152939
R16261 GND.n4107 GND.n4106 0.152939
R16262 GND.n4107 GND.n2064 0.152939
R16263 GND.n4121 GND.n2064 0.152939
R16264 GND.n4122 GND.n4121 0.152939
R16265 GND.n4123 GND.n4122 0.152939
R16266 GND.n4123 GND.n2050 0.152939
R16267 GND.n4139 GND.n2050 0.152939
R16268 GND.n4140 GND.n4139 0.152939
R16269 GND.n4141 GND.n4140 0.152939
R16270 GND.n4143 GND.n4141 0.152939
R16271 GND.n4143 GND.n4142 0.152939
R16272 GND.n4142 GND.n1560 0.152939
R16273 GND.n1561 GND.n1560 0.152939
R16274 GND.n1562 GND.n1561 0.152939
R16275 GND.n1830 GND.n1562 0.152939
R16276 GND.n1831 GND.n1830 0.152939
R16277 GND.n1831 GND.n1828 0.152939
R16278 GND.n1837 GND.n1828 0.152939
R16279 GND.n1838 GND.n1837 0.152939
R16280 GND.n1839 GND.n1838 0.152939
R16281 GND.n1839 GND.n1824 0.152939
R16282 GND.n1845 GND.n1824 0.152939
R16283 GND.n1846 GND.n1845 0.152939
R16284 GND.n1847 GND.n1846 0.152939
R16285 GND.n1847 GND.n1820 0.152939
R16286 GND.n1853 GND.n1820 0.152939
R16287 GND.n1854 GND.n1853 0.152939
R16288 GND.n1855 GND.n1854 0.152939
R16289 GND.n1855 GND.n1816 0.152939
R16290 GND.n1861 GND.n1816 0.152939
R16291 GND.n1862 GND.n1861 0.152939
R16292 GND.n1863 GND.n1862 0.152939
R16293 GND.n1863 GND.n1812 0.152939
R16294 GND.n1869 GND.n1812 0.152939
R16295 GND.n1870 GND.n1869 0.152939
R16296 GND.n1871 GND.n1870 0.152939
R16297 GND.n1871 GND.n1808 0.152939
R16298 GND.n1878 GND.n1808 0.152939
R16299 GND.n1879 GND.n1878 0.152939
R16300 GND.n1880 GND.n1879 0.152939
R16301 GND.n3762 GND.n3761 0.152939
R16302 GND.n3762 GND.n3045 0.152939
R16303 GND.n3784 GND.n3045 0.152939
R16304 GND.n3785 GND.n3784 0.152939
R16305 GND.n3786 GND.n3785 0.152939
R16306 GND.n3787 GND.n3786 0.152939
R16307 GND.n3787 GND.n3022 0.152939
R16308 GND.n3808 GND.n3022 0.152939
R16309 GND.n3809 GND.n3808 0.152939
R16310 GND.n3810 GND.n3809 0.152939
R16311 GND.n3811 GND.n3810 0.152939
R16312 GND.n3811 GND.n2999 0.152939
R16313 GND.n3833 GND.n2999 0.152939
R16314 GND.n3834 GND.n3833 0.152939
R16315 GND.n3835 GND.n3834 0.152939
R16316 GND.n3836 GND.n3835 0.152939
R16317 GND.n3836 GND.n2977 0.152939
R16318 GND.n3861 GND.n2977 0.152939
R16319 GND.n3862 GND.n3861 0.152939
R16320 GND.n3863 GND.n3862 0.152939
R16321 GND.n3863 GND.n1298 0.152939
R16322 GND.n4950 GND.n1298 0.152939
R16323 GND.n3365 GND.n3360 0.152939
R16324 GND.n3366 GND.n3365 0.152939
R16325 GND.n3367 GND.n3366 0.152939
R16326 GND.n3367 GND.n3356 0.152939
R16327 GND.n3375 GND.n3356 0.152939
R16328 GND.n3376 GND.n3375 0.152939
R16329 GND.n3377 GND.n3376 0.152939
R16330 GND.n3377 GND.n3352 0.152939
R16331 GND.n3385 GND.n3352 0.152939
R16332 GND.n3386 GND.n3385 0.152939
R16333 GND.n3387 GND.n3386 0.152939
R16334 GND.n3387 GND.n3346 0.152939
R16335 GND.n3395 GND.n3346 0.152939
R16336 GND.n3396 GND.n3395 0.152939
R16337 GND.n3397 GND.n3396 0.152939
R16338 GND.n3397 GND.n3342 0.152939
R16339 GND.n3405 GND.n3342 0.152939
R16340 GND.n3406 GND.n3405 0.152939
R16341 GND.n3407 GND.n3406 0.152939
R16342 GND.n3407 GND.n3338 0.152939
R16343 GND.n3415 GND.n3338 0.152939
R16344 GND.n3416 GND.n3415 0.152939
R16345 GND.n3417 GND.n3416 0.152939
R16346 GND.n3417 GND.n3334 0.152939
R16347 GND.n3427 GND.n3334 0.152939
R16348 GND.n3428 GND.n3427 0.152939
R16349 GND.n3429 GND.n3428 0.152939
R16350 GND.n3429 GND.n3330 0.152939
R16351 GND.n3437 GND.n3330 0.152939
R16352 GND.n3438 GND.n3437 0.152939
R16353 GND.n3439 GND.n3438 0.152939
R16354 GND.n3439 GND.n3326 0.152939
R16355 GND.n3447 GND.n3326 0.152939
R16356 GND.n3448 GND.n3447 0.152939
R16357 GND.n3449 GND.n3448 0.152939
R16358 GND.n3449 GND.n3322 0.152939
R16359 GND.n3460 GND.n3322 0.152939
R16360 GND.n3461 GND.n3460 0.152939
R16361 GND.n3462 GND.n3461 0.152939
R16362 GND.n3462 GND.n3318 0.152939
R16363 GND.n3470 GND.n3318 0.152939
R16364 GND.n3471 GND.n3470 0.152939
R16365 GND.n3472 GND.n3471 0.152939
R16366 GND.n3472 GND.n3314 0.152939
R16367 GND.n3480 GND.n3314 0.152939
R16368 GND.n3481 GND.n3480 0.152939
R16369 GND.n3482 GND.n3481 0.152939
R16370 GND.n3482 GND.n3308 0.152939
R16371 GND.n3489 GND.n3308 0.152939
R16372 GND.n1170 GND.n1169 0.152939
R16373 GND.n1171 GND.n1170 0.152939
R16374 GND.n3289 GND.n1171 0.152939
R16375 GND.n3615 GND.n3289 0.152939
R16376 GND.n3616 GND.n3615 0.152939
R16377 GND.n3617 GND.n3616 0.152939
R16378 GND.n3618 GND.n3617 0.152939
R16379 GND.n3618 GND.n3266 0.152939
R16380 GND.n3639 GND.n3266 0.152939
R16381 GND.n3640 GND.n3639 0.152939
R16382 GND.n3641 GND.n3640 0.152939
R16383 GND.n3642 GND.n3641 0.152939
R16384 GND.n3642 GND.n3243 0.152939
R16385 GND.n3664 GND.n3243 0.152939
R16386 GND.n3665 GND.n3664 0.152939
R16387 GND.n3666 GND.n3665 0.152939
R16388 GND.n3667 GND.n3666 0.152939
R16389 GND.n3667 GND.n3221 0.152939
R16390 GND.n3689 GND.n3221 0.152939
R16391 GND.n3690 GND.n3689 0.152939
R16392 GND.n3691 GND.n3690 0.152939
R16393 GND.n3691 GND.n3068 0.152939
R16394 GND.n5129 GND.n1080 0.152939
R16395 GND.n1085 GND.n1080 0.152939
R16396 GND.n1086 GND.n1085 0.152939
R16397 GND.n1087 GND.n1086 0.152939
R16398 GND.n1092 GND.n1087 0.152939
R16399 GND.n1093 GND.n1092 0.152939
R16400 GND.n1094 GND.n1093 0.152939
R16401 GND.n1095 GND.n1094 0.152939
R16402 GND.n1100 GND.n1095 0.152939
R16403 GND.n1101 GND.n1100 0.152939
R16404 GND.n1102 GND.n1101 0.152939
R16405 GND.n1103 GND.n1102 0.152939
R16406 GND.n1108 GND.n1103 0.152939
R16407 GND.n1109 GND.n1108 0.152939
R16408 GND.n1110 GND.n1109 0.152939
R16409 GND.n1111 GND.n1110 0.152939
R16410 GND.n1116 GND.n1111 0.152939
R16411 GND.n1117 GND.n1116 0.152939
R16412 GND.n1118 GND.n1117 0.152939
R16413 GND.n1119 GND.n1118 0.152939
R16414 GND.n1124 GND.n1119 0.152939
R16415 GND.n1125 GND.n1124 0.152939
R16416 GND.n1126 GND.n1125 0.152939
R16417 GND.n1127 GND.n1126 0.152939
R16418 GND.n1132 GND.n1127 0.152939
R16419 GND.n1133 GND.n1132 0.152939
R16420 GND.n1134 GND.n1133 0.152939
R16421 GND.n1135 GND.n1134 0.152939
R16422 GND.n1140 GND.n1135 0.152939
R16423 GND.n1141 GND.n1140 0.152939
R16424 GND.n1142 GND.n1141 0.152939
R16425 GND.n1143 GND.n1142 0.152939
R16426 GND.n1148 GND.n1143 0.152939
R16427 GND.n1149 GND.n1148 0.152939
R16428 GND.n1150 GND.n1149 0.152939
R16429 GND.n1151 GND.n1150 0.152939
R16430 GND.n1156 GND.n1151 0.152939
R16431 GND.n1157 GND.n1156 0.152939
R16432 GND.n1158 GND.n1157 0.152939
R16433 GND.n1159 GND.n1158 0.152939
R16434 GND.n3542 GND.n1159 0.152939
R16435 GND.n3543 GND.n3542 0.152939
R16436 GND.n3543 GND.n3540 0.152939
R16437 GND.n3549 GND.n3540 0.152939
R16438 GND.n3550 GND.n3549 0.152939
R16439 GND.n3551 GND.n3550 0.152939
R16440 GND.n3552 GND.n3551 0.152939
R16441 GND.n3553 GND.n3552 0.152939
R16442 GND.n3556 GND.n3553 0.152939
R16443 GND.n3557 GND.n3556 0.152939
R16444 GND.n3558 GND.n3557 0.152939
R16445 GND.n3559 GND.n3558 0.152939
R16446 GND.n3562 GND.n3559 0.152939
R16447 GND.n3563 GND.n3562 0.152939
R16448 GND.n3564 GND.n3563 0.152939
R16449 GND.n3565 GND.n3564 0.152939
R16450 GND.n3568 GND.n3565 0.152939
R16451 GND.n3569 GND.n3568 0.152939
R16452 GND.n3570 GND.n3569 0.152939
R16453 GND.n3571 GND.n3570 0.152939
R16454 GND.n3574 GND.n3571 0.152939
R16455 GND.n3575 GND.n3574 0.152939
R16456 GND.n3576 GND.n3575 0.152939
R16457 GND.n5243 GND.n970 0.152939
R16458 GND.n975 GND.n970 0.152939
R16459 GND.n976 GND.n975 0.152939
R16460 GND.n977 GND.n976 0.152939
R16461 GND.n982 GND.n977 0.152939
R16462 GND.n983 GND.n982 0.152939
R16463 GND.n984 GND.n983 0.152939
R16464 GND.n985 GND.n984 0.152939
R16465 GND.n990 GND.n985 0.152939
R16466 GND.n991 GND.n990 0.152939
R16467 GND.n992 GND.n991 0.152939
R16468 GND.n993 GND.n992 0.152939
R16469 GND.n998 GND.n993 0.152939
R16470 GND.n999 GND.n998 0.152939
R16471 GND.n1000 GND.n999 0.152939
R16472 GND.n1001 GND.n1000 0.152939
R16473 GND.n1006 GND.n1001 0.152939
R16474 GND.n1007 GND.n1006 0.152939
R16475 GND.n1008 GND.n1007 0.152939
R16476 GND.n1009 GND.n1008 0.152939
R16477 GND.n1014 GND.n1009 0.152939
R16478 GND.n1015 GND.n1014 0.152939
R16479 GND.n1016 GND.n1015 0.152939
R16480 GND.n1017 GND.n1016 0.152939
R16481 GND.n1022 GND.n1017 0.152939
R16482 GND.n1023 GND.n1022 0.152939
R16483 GND.n1024 GND.n1023 0.152939
R16484 GND.n1025 GND.n1024 0.152939
R16485 GND.n1030 GND.n1025 0.152939
R16486 GND.n1031 GND.n1030 0.152939
R16487 GND.n1032 GND.n1031 0.152939
R16488 GND.n1033 GND.n1032 0.152939
R16489 GND.n1038 GND.n1033 0.152939
R16490 GND.n1039 GND.n1038 0.152939
R16491 GND.n1040 GND.n1039 0.152939
R16492 GND.n1041 GND.n1040 0.152939
R16493 GND.n1046 GND.n1041 0.152939
R16494 GND.n1047 GND.n1046 0.152939
R16495 GND.n1048 GND.n1047 0.152939
R16496 GND.n1049 GND.n1048 0.152939
R16497 GND.n1054 GND.n1049 0.152939
R16498 GND.n1055 GND.n1054 0.152939
R16499 GND.n1056 GND.n1055 0.152939
R16500 GND.n1057 GND.n1056 0.152939
R16501 GND.n1062 GND.n1057 0.152939
R16502 GND.n1063 GND.n1062 0.152939
R16503 GND.n1064 GND.n1063 0.152939
R16504 GND.n1065 GND.n1064 0.152939
R16505 GND.n1070 GND.n1065 0.152939
R16506 GND.n1071 GND.n1070 0.152939
R16507 GND.n1072 GND.n1071 0.152939
R16508 GND.n1073 GND.n1072 0.152939
R16509 GND.n1078 GND.n1073 0.152939
R16510 GND.n1079 GND.n1078 0.152939
R16511 GND.n5130 GND.n1079 0.152939
R16512 GND.n4822 GND.n4821 0.152939
R16513 GND.n4821 GND.n4820 0.152939
R16514 GND.n4820 GND.n4804 0.152939
R16515 GND.n4816 GND.n4804 0.152939
R16516 GND.n4816 GND.n4815 0.152939
R16517 GND.n4815 GND.n4814 0.152939
R16518 GND.n4814 GND.n4809 0.152939
R16519 GND.n4809 GND.n1400 0.152939
R16520 GND.n4803 GND.n1467 0.152939
R16521 GND.n4799 GND.n1467 0.152939
R16522 GND.n4799 GND.n4798 0.152939
R16523 GND.n4798 GND.n4797 0.152939
R16524 GND.n4797 GND.n1471 0.152939
R16525 GND.n4793 GND.n1471 0.152939
R16526 GND.n4793 GND.n4792 0.152939
R16527 GND.n4792 GND.n4791 0.152939
R16528 GND.n4791 GND.n1476 0.152939
R16529 GND.n4787 GND.n1476 0.152939
R16530 GND.n4787 GND.n4786 0.152939
R16531 GND.n4786 GND.n4785 0.152939
R16532 GND.n4785 GND.n1481 0.152939
R16533 GND.n4781 GND.n1481 0.152939
R16534 GND.n4781 GND.n4780 0.152939
R16535 GND.n4780 GND.n4779 0.152939
R16536 GND.n4779 GND.n1486 0.152939
R16537 GND.n4775 GND.n1486 0.152939
R16538 GND.n4775 GND.n4774 0.152939
R16539 GND.n4774 GND.n4773 0.152939
R16540 GND.n4773 GND.n1491 0.152939
R16541 GND.n4769 GND.n1491 0.152939
R16542 GND.n4769 GND.n4768 0.152939
R16543 GND.n4768 GND.n4767 0.152939
R16544 GND.n4767 GND.n1496 0.152939
R16545 GND.n4763 GND.n1496 0.152939
R16546 GND.n4763 GND.n4762 0.152939
R16547 GND.n4762 GND.n4761 0.152939
R16548 GND.n4761 GND.n1501 0.152939
R16549 GND.n4757 GND.n1501 0.152939
R16550 GND.n4757 GND.n4756 0.152939
R16551 GND.n4756 GND.n4755 0.152939
R16552 GND.n4755 GND.n1506 0.152939
R16553 GND.n4751 GND.n1506 0.152939
R16554 GND.n4751 GND.n4750 0.152939
R16555 GND.n4750 GND.n4749 0.152939
R16556 GND.n4749 GND.n1511 0.152939
R16557 GND.n4745 GND.n1511 0.152939
R16558 GND.n4745 GND.n4744 0.152939
R16559 GND.n4744 GND.n4743 0.152939
R16560 GND.n4743 GND.n1516 0.152939
R16561 GND.n4739 GND.n1516 0.152939
R16562 GND.n4739 GND.n4738 0.152939
R16563 GND.n4738 GND.n4737 0.152939
R16564 GND.n4737 GND.n1521 0.152939
R16565 GND.n4733 GND.n1521 0.152939
R16566 GND.n4733 GND.n4732 0.152939
R16567 GND.n4732 GND.n4731 0.152939
R16568 GND.n4731 GND.n1526 0.152939
R16569 GND.n4727 GND.n1526 0.152939
R16570 GND.n4727 GND.n4726 0.152939
R16571 GND.n4726 GND.n4725 0.152939
R16572 GND.n4725 GND.n1531 0.152939
R16573 GND.n4721 GND.n1531 0.152939
R16574 GND.n4721 GND.n4720 0.152939
R16575 GND.n4720 GND.n4719 0.152939
R16576 GND.n4719 GND.n1536 0.152939
R16577 GND.n4715 GND.n1536 0.152939
R16578 GND.n4715 GND.n4714 0.152939
R16579 GND.n4714 GND.n4713 0.152939
R16580 GND.n4713 GND.n1541 0.152939
R16581 GND.n4709 GND.n1541 0.152939
R16582 GND.n4709 GND.n4708 0.152939
R16583 GND.n4708 GND.n4707 0.152939
R16584 GND.n4707 GND.n1546 0.152939
R16585 GND.n4703 GND.n1546 0.152939
R16586 GND.n4703 GND.n4702 0.152939
R16587 GND.n4702 GND.n4701 0.152939
R16588 GND.n4701 GND.n1551 0.152939
R16589 GND.n1957 GND.n1956 0.152939
R16590 GND.n1965 GND.n1956 0.152939
R16591 GND.n1966 GND.n1965 0.152939
R16592 GND.n1967 GND.n1966 0.152939
R16593 GND.n1967 GND.n1952 0.152939
R16594 GND.n1975 GND.n1952 0.152939
R16595 GND.n1976 GND.n1975 0.152939
R16596 GND.n1977 GND.n1976 0.152939
R16597 GND.n3876 GND.n3875 0.152939
R16598 GND.n3876 GND.n2956 0.152939
R16599 GND.n3890 GND.n2956 0.152939
R16600 GND.n3891 GND.n3890 0.152939
R16601 GND.n3892 GND.n3891 0.152939
R16602 GND.n3892 GND.n2261 0.152939
R16603 GND.n3906 GND.n2261 0.152939
R16604 GND.n3907 GND.n3906 0.152939
R16605 GND.n3908 GND.n3907 0.152939
R16606 GND.n3908 GND.n2246 0.152939
R16607 GND.n3922 GND.n2246 0.152939
R16608 GND.n3923 GND.n3922 0.152939
R16609 GND.n3924 GND.n3923 0.152939
R16610 GND.n3924 GND.n2232 0.152939
R16611 GND.n3938 GND.n2232 0.152939
R16612 GND.n3939 GND.n3938 0.152939
R16613 GND.n3940 GND.n3939 0.152939
R16614 GND.n3940 GND.n2217 0.152939
R16615 GND.n3954 GND.n2217 0.152939
R16616 GND.n3955 GND.n3954 0.152939
R16617 GND.n3956 GND.n3955 0.152939
R16618 GND.n3956 GND.n2203 0.152939
R16619 GND.n3970 GND.n2203 0.152939
R16620 GND.n3971 GND.n3970 0.152939
R16621 GND.n3972 GND.n3971 0.152939
R16622 GND.n3972 GND.n2187 0.152939
R16623 GND.n3986 GND.n2187 0.152939
R16624 GND.n3987 GND.n3986 0.152939
R16625 GND.n3988 GND.n3987 0.152939
R16626 GND.n3988 GND.n2173 0.152939
R16627 GND.n4002 GND.n2173 0.152939
R16628 GND.n4003 GND.n4002 0.152939
R16629 GND.n4004 GND.n4003 0.152939
R16630 GND.n4004 GND.n2158 0.152939
R16631 GND.n4018 GND.n2158 0.152939
R16632 GND.n4019 GND.n4018 0.152939
R16633 GND.n4020 GND.n4019 0.152939
R16634 GND.n4020 GND.n2144 0.152939
R16635 GND.n4034 GND.n2144 0.152939
R16636 GND.n4035 GND.n4034 0.152939
R16637 GND.n4036 GND.n4035 0.152939
R16638 GND.n4036 GND.n2130 0.152939
R16639 GND.n4050 GND.n2130 0.152939
R16640 GND.n4051 GND.n4050 0.152939
R16641 GND.n4052 GND.n4051 0.152939
R16642 GND.n4052 GND.n2115 0.152939
R16643 GND.n4066 GND.n2115 0.152939
R16644 GND.n4067 GND.n4066 0.152939
R16645 GND.n4068 GND.n4067 0.152939
R16646 GND.n4068 GND.n2100 0.152939
R16647 GND.n4082 GND.n2100 0.152939
R16648 GND.n4083 GND.n4082 0.152939
R16649 GND.n4084 GND.n4083 0.152939
R16650 GND.n4084 GND.n2087 0.152939
R16651 GND.n4097 GND.n2087 0.152939
R16652 GND.n4098 GND.n4097 0.152939
R16653 GND.n4099 GND.n4098 0.152939
R16654 GND.n4099 GND.n2071 0.152939
R16655 GND.n4113 GND.n2071 0.152939
R16656 GND.n4114 GND.n4113 0.152939
R16657 GND.n4115 GND.n4114 0.152939
R16658 GND.n4115 GND.n2057 0.152939
R16659 GND.n4129 GND.n2057 0.152939
R16660 GND.n4130 GND.n4129 0.152939
R16661 GND.n4133 GND.n4130 0.152939
R16662 GND.n4133 GND.n4132 0.152939
R16663 GND.n4132 GND.n4131 0.152939
R16664 GND.n4131 GND.n2042 0.152939
R16665 GND.n4152 GND.n2042 0.152939
R16666 GND.n3712 GND.n3206 0.152939
R16667 GND.n3713 GND.n3712 0.152939
R16668 GND.n3714 GND.n3713 0.152939
R16669 GND.n3714 GND.n3057 0.152939
R16670 GND.n3769 GND.n3057 0.152939
R16671 GND.n3770 GND.n3769 0.152939
R16672 GND.n3772 GND.n3770 0.152939
R16673 GND.n3772 GND.n3771 0.152939
R16674 GND.n3771 GND.n3035 0.152939
R16675 GND.n3794 GND.n3035 0.152939
R16676 GND.n3795 GND.n3794 0.152939
R16677 GND.n3797 GND.n3795 0.152939
R16678 GND.n3797 GND.n3796 0.152939
R16679 GND.n3796 GND.n3011 0.152939
R16680 GND.n3818 GND.n3011 0.152939
R16681 GND.n3819 GND.n3818 0.152939
R16682 GND.n3821 GND.n3819 0.152939
R16683 GND.n3821 GND.n3820 0.152939
R16684 GND.n3820 GND.n2988 0.152939
R16685 GND.n3843 GND.n2988 0.152939
R16686 GND.n3844 GND.n3843 0.152939
R16687 GND.n3851 GND.n3844 0.152939
R16688 GND.n3851 GND.n3850 0.152939
R16689 GND.n3850 GND.n3849 0.152939
R16690 GND.n3849 GND.n3845 0.152939
R16691 GND.n3845 GND.n2968 0.152939
R16692 GND.n3873 GND.n2968 0.152939
R16693 GND.n4949 GND.n1299 0.152939
R16694 GND.n4945 GND.n1299 0.152939
R16695 GND.n4945 GND.n4944 0.152939
R16696 GND.n4944 GND.n4943 0.152939
R16697 GND.n4943 GND.n1303 0.152939
R16698 GND.n4939 GND.n1303 0.152939
R16699 GND.n4939 GND.n4938 0.152939
R16700 GND.n4938 GND.n4937 0.152939
R16701 GND.n4937 GND.n1308 0.152939
R16702 GND.n1313 GND.n1308 0.152939
R16703 GND.n4932 GND.n1313 0.152939
R16704 GND.n4932 GND.n4931 0.152939
R16705 GND.n4931 GND.n4930 0.152939
R16706 GND.n4930 GND.n1317 0.152939
R16707 GND.n4926 GND.n1317 0.152939
R16708 GND.n4926 GND.n4925 0.152939
R16709 GND.n4925 GND.n4924 0.152939
R16710 GND.n4924 GND.n1322 0.152939
R16711 GND.n4920 GND.n1322 0.152939
R16712 GND.n4920 GND.n4919 0.152939
R16713 GND.n4919 GND.n4918 0.152939
R16714 GND.n4908 GND.n1350 0.152939
R16715 GND.n4908 GND.n4907 0.152939
R16716 GND.n4907 GND.n4906 0.152939
R16717 GND.n4906 GND.n1351 0.152939
R16718 GND.n4902 GND.n1351 0.152939
R16719 GND.n4902 GND.n4901 0.152939
R16720 GND.n4901 GND.n4900 0.152939
R16721 GND.n4900 GND.n1358 0.152939
R16722 GND.n4896 GND.n1358 0.152939
R16723 GND.n4896 GND.n4895 0.152939
R16724 GND.n4895 GND.n4894 0.152939
R16725 GND.n4894 GND.n1366 0.152939
R16726 GND.n4889 GND.n1366 0.152939
R16727 GND.n4889 GND.n4888 0.152939
R16728 GND.n4888 GND.n4887 0.152939
R16729 GND.n4887 GND.n1376 0.152939
R16730 GND.n4883 GND.n1376 0.152939
R16731 GND.n4883 GND.n4882 0.152939
R16732 GND.n4882 GND.n4881 0.152939
R16733 GND.n4881 GND.n1384 0.152939
R16734 GND.n4877 GND.n1384 0.152939
R16735 GND.n4877 GND.n4876 0.152939
R16736 GND.n4876 GND.n4875 0.152939
R16737 GND.n4875 GND.n1392 0.152939
R16738 GND.n4871 GND.n1392 0.152939
R16739 GND.n3494 GND.n3306 0.152939
R16740 GND.n3502 GND.n3306 0.152939
R16741 GND.n3503 GND.n3502 0.152939
R16742 GND.n3504 GND.n3503 0.152939
R16743 GND.n3504 GND.n3302 0.152939
R16744 GND.n3512 GND.n3302 0.152939
R16745 GND.n3513 GND.n3512 0.152939
R16746 GND.n3515 GND.n3513 0.152939
R16747 GND.n3515 GND.n3514 0.152939
R16748 GND.n3514 GND.n3295 0.152939
R16749 GND.n3524 GND.n3295 0.152939
R16750 GND.n3525 GND.n3294 0.152939
R16751 GND.n3532 GND.n3294 0.152939
R16752 GND.n3533 GND.n3532 0.152939
R16753 GND.n3534 GND.n3533 0.152939
R16754 GND.n3534 GND.n3279 0.152939
R16755 GND.n3625 GND.n3279 0.152939
R16756 GND.n3626 GND.n3625 0.152939
R16757 GND.n3628 GND.n3626 0.152939
R16758 GND.n3628 GND.n3627 0.152939
R16759 GND.n3627 GND.n3255 0.152939
R16760 GND.n3649 GND.n3255 0.152939
R16761 GND.n3650 GND.n3649 0.152939
R16762 GND.n3652 GND.n3650 0.152939
R16763 GND.n3652 GND.n3651 0.152939
R16764 GND.n3651 GND.n3232 0.152939
R16765 GND.n3674 GND.n3232 0.152939
R16766 GND.n3675 GND.n3674 0.152939
R16767 GND.n3677 GND.n3675 0.152939
R16768 GND.n3677 GND.n3676 0.152939
R16769 GND.n3676 GND.n3210 0.152939
R16770 GND.n3697 GND.n3210 0.152939
R16771 GND.n3698 GND.n3697 0.152939
R16772 GND.n3699 GND.n3698 0.152939
R16773 GND.n3699 GND.n3208 0.152939
R16774 GND.n3705 GND.n3208 0.152939
R16775 GND.n3706 GND.n3705 0.152939
R16776 GND.n3708 GND.n3706 0.152939
R16777 GND.n4288 GND.n163 0.131598
R16778 GND.n3576 GND.n3069 0.131598
R16779 GND.n6331 GND.n161 0.0767195
R16780 GND.n6331 GND.n162 0.0767195
R16781 GND.n3761 GND.n3760 0.0767195
R16782 GND.n3760 GND.n3068 0.0767195
R16783 GND.n6339 GND.n148 0.0695946
R16784 GND.n6339 GND.n6338 0.0695946
R16785 GND.n3707 GND.n3206 0.0695946
R16786 GND.n3708 GND.n3707 0.0695946
R16787 GND.n4591 GND.n1659 0.063
R16788 GND.n4870 GND.n4869 0.063
R16789 GND.n4869 GND.n1400 0.0523293
R16790 GND.n1977 GND.n1659 0.0523293
R16791 GND.n4591 GND.n4590 0.046356
R16792 GND.n6163 GND.n6162 0.046356
R16793 GND.n3493 GND.n3492 0.046356
R16794 GND.n4870 GND.n1287 0.046356
R16795 GND.n4590 GND.n1661 0.0344674
R16796 GND.n4157 GND.n1661 0.0344674
R16797 GND.n4157 GND.n1686 0.0344674
R16798 GND.n1687 GND.n1686 0.0344674
R16799 GND.n1688 GND.n1687 0.0344674
R16800 GND.n4172 GND.n1688 0.0344674
R16801 GND.n4172 GND.n1707 0.0344674
R16802 GND.n1708 GND.n1707 0.0344674
R16803 GND.n1709 GND.n1708 0.0344674
R16804 GND.n4187 GND.n1709 0.0344674
R16805 GND.n4187 GND.n1728 0.0344674
R16806 GND.n1729 GND.n1728 0.0344674
R16807 GND.n1730 GND.n1729 0.0344674
R16808 GND.n4202 GND.n1730 0.0344674
R16809 GND.n4202 GND.n1749 0.0344674
R16810 GND.n1750 GND.n1749 0.0344674
R16811 GND.n1751 GND.n1750 0.0344674
R16812 GND.n4217 GND.n1751 0.0344674
R16813 GND.n4217 GND.n1770 0.0344674
R16814 GND.n1771 GND.n1770 0.0344674
R16815 GND.n1772 GND.n1771 0.0344674
R16816 GND.n4232 GND.n1772 0.0344674
R16817 GND.n4232 GND.n1789 0.0344674
R16818 GND.n1790 GND.n1789 0.0344674
R16819 GND.n1791 GND.n1790 0.0344674
R16820 GND.n4252 GND.n1791 0.0344674
R16821 GND.n4253 GND.n4252 0.0344674
R16822 GND.n4257 GND.n4253 0.0344674
R16823 GND.n4257 GND.n1896 0.0344674
R16824 GND.n4494 GND.n1896 0.0344674
R16825 GND.n4494 GND.n1897 0.0344674
R16826 GND.n1897 GND.n179 0.0344674
R16827 GND.n180 GND.n179 0.0344674
R16828 GND.n181 GND.n180 0.0344674
R16829 GND.n4268 GND.n181 0.0344674
R16830 GND.n4268 GND.n199 0.0344674
R16831 GND.n200 GND.n199 0.0344674
R16832 GND.n201 GND.n200 0.0344674
R16833 GND.n4346 GND.n201 0.0344674
R16834 GND.n4346 GND.n219 0.0344674
R16835 GND.n220 GND.n219 0.0344674
R16836 GND.n221 GND.n220 0.0344674
R16837 GND.n4340 GND.n221 0.0344674
R16838 GND.n4340 GND.n240 0.0344674
R16839 GND.n241 GND.n240 0.0344674
R16840 GND.n242 GND.n241 0.0344674
R16841 GND.n4335 GND.n242 0.0344674
R16842 GND.n4335 GND.n261 0.0344674
R16843 GND.n262 GND.n261 0.0344674
R16844 GND.n263 GND.n262 0.0344674
R16845 GND.n4386 GND.n263 0.0344674
R16846 GND.n4386 GND.n281 0.0344674
R16847 GND.n282 GND.n281 0.0344674
R16848 GND.n283 GND.n282 0.0344674
R16849 GND.n6162 GND.n283 0.0344674
R16850 GND.n3492 GND.n1182 0.0344674
R16851 GND.n5035 GND.n1182 0.0344674
R16852 GND.n5035 GND.n1183 0.0344674
R16853 GND.n5031 GND.n1183 0.0344674
R16854 GND.n5031 GND.n5030 0.0344674
R16855 GND.n5030 GND.n5029 0.0344674
R16856 GND.n5029 GND.n1191 0.0344674
R16857 GND.n5025 GND.n1191 0.0344674
R16858 GND.n5025 GND.n5024 0.0344674
R16859 GND.n5024 GND.n5023 0.0344674
R16860 GND.n5023 GND.n1199 0.0344674
R16861 GND.n5019 GND.n1199 0.0344674
R16862 GND.n5019 GND.n5018 0.0344674
R16863 GND.n5018 GND.n5017 0.0344674
R16864 GND.n5017 GND.n1207 0.0344674
R16865 GND.n5013 GND.n1207 0.0344674
R16866 GND.n5013 GND.n5012 0.0344674
R16867 GND.n5012 GND.n5011 0.0344674
R16868 GND.n5011 GND.n1215 0.0344674
R16869 GND.n5007 GND.n1215 0.0344674
R16870 GND.n5007 GND.n5006 0.0344674
R16871 GND.n5006 GND.n5005 0.0344674
R16872 GND.n5005 GND.n1223 0.0344674
R16873 GND.n5001 GND.n1223 0.0344674
R16874 GND.n5001 GND.n5000 0.0344674
R16875 GND.n5000 GND.n4999 0.0344674
R16876 GND.n4999 GND.n1231 0.0344674
R16877 GND.n4995 GND.n1231 0.0344674
R16878 GND.n4995 GND.n4994 0.0344674
R16879 GND.n4994 GND.n4993 0.0344674
R16880 GND.n4993 GND.n1239 0.0344674
R16881 GND.n4989 GND.n1239 0.0344674
R16882 GND.n4989 GND.n4988 0.0344674
R16883 GND.n4988 GND.n4987 0.0344674
R16884 GND.n4987 GND.n1247 0.0344674
R16885 GND.n4983 GND.n1247 0.0344674
R16886 GND.n4983 GND.n4982 0.0344674
R16887 GND.n4982 GND.n4981 0.0344674
R16888 GND.n4981 GND.n1255 0.0344674
R16889 GND.n4977 GND.n1255 0.0344674
R16890 GND.n4977 GND.n4976 0.0344674
R16891 GND.n4976 GND.n4975 0.0344674
R16892 GND.n4975 GND.n1263 0.0344674
R16893 GND.n4971 GND.n1263 0.0344674
R16894 GND.n4971 GND.n4970 0.0344674
R16895 GND.n4970 GND.n4969 0.0344674
R16896 GND.n4969 GND.n1271 0.0344674
R16897 GND.n4965 GND.n1271 0.0344674
R16898 GND.n4965 GND.n4964 0.0344674
R16899 GND.n4964 GND.n4963 0.0344674
R16900 GND.n4963 GND.n1279 0.0344674
R16901 GND.n4959 GND.n1279 0.0344674
R16902 GND.n4959 GND.n4958 0.0344674
R16903 GND.n4958 GND.n4957 0.0344674
R16904 GND.n4957 GND.n1287 0.0344674
R16905 GND.n2041 GND.n1923 0.0343753
R16906 GND.n4831 GND.n1444 0.0343753
R16907 GND.n1948 GND.n1947 0.0286165
R16908 GND.n1987 GND.n1985 0.0286165
R16909 GND.n1986 GND.n1944 0.0286165
R16910 GND.n1996 GND.n1995 0.0286165
R16911 GND.n1945 GND.n1940 0.0286165
R16912 GND.n2006 GND.n2004 0.0286165
R16913 GND.n2005 GND.n1937 0.0286165
R16914 GND.n2015 GND.n2014 0.0286165
R16915 GND.n1938 GND.n1933 0.0286165
R16916 GND.n2028 GND.n2026 0.0286165
R16917 GND.n2027 GND.n1927 0.0286165
R16918 GND.n2034 GND.n2033 0.0286165
R16919 GND.n4868 GND.n1401 0.0286165
R16920 GND.n4865 GND.n4864 0.0286165
R16921 GND.n4861 GND.n1406 0.0286165
R16922 GND.n4860 GND.n1413 0.0286165
R16923 GND.n4857 GND.n4856 0.0286165
R16924 GND.n4853 GND.n1417 0.0286165
R16925 GND.n4852 GND.n1424 0.0286165
R16926 GND.n4849 GND.n4848 0.0286165
R16927 GND.n4845 GND.n1428 0.0286165
R16928 GND.n4844 GND.n1434 0.0286165
R16929 GND.n4838 GND.n4837 0.0286165
R16930 GND.n4832 GND.n1438 0.0286165
R16931 GND.n1948 GND.n1659 0.0228577
R16932 GND.n4869 GND.n4868 0.0228577
R16933 GND.n3115 GND.n3069 0.0218415
R16934 GND.n1880 GND.n163 0.0218415
R16935 GND.n4153 GND.n2041 0.0113401
R16936 GND.n3874 GND.n1444 0.0113401
R16937 GND.n1985 GND.n1947 0.00625881
R16938 GND.n1987 GND.n1986 0.00625881
R16939 GND.n1996 GND.n1944 0.00625881
R16940 GND.n1995 GND.n1945 0.00625881
R16941 GND.n2004 GND.n1940 0.00625881
R16942 GND.n2006 GND.n2005 0.00625881
R16943 GND.n2015 GND.n1937 0.00625881
R16944 GND.n2014 GND.n1938 0.00625881
R16945 GND.n2026 GND.n1933 0.00625881
R16946 GND.n2028 GND.n2027 0.00625881
R16947 GND.n2034 GND.n1927 0.00625881
R16948 GND.n2033 GND.n1923 0.00625881
R16949 GND.n4865 GND.n1401 0.00625881
R16950 GND.n4864 GND.n1406 0.00625881
R16951 GND.n4861 GND.n4860 0.00625881
R16952 GND.n4857 GND.n1413 0.00625881
R16953 GND.n4856 GND.n1417 0.00625881
R16954 GND.n4853 GND.n4852 0.00625881
R16955 GND.n4849 GND.n1424 0.00625881
R16956 GND.n4848 GND.n1428 0.00625881
R16957 GND.n4845 GND.n4844 0.00625881
R16958 GND.n4838 GND.n1434 0.00625881
R16959 GND.n4837 GND.n1438 0.00625881
R16960 GND.n4832 GND.n4831 0.00625881
R16961 a_n1672_n179.n23 a_n1672_n179.n20 289.615
R16962 a_n1672_n179.n33 a_n1672_n179.n30 289.615
R16963 a_n1672_n179.n43 a_n1672_n179.n18 289.615
R16964 a_n1672_n179.n0 a_n1672_n179.n36 199.814
R16965 a_n1672_n179.n0 a_n1672_n179.n26 199.788
R16966 a_n1672_n179.n42 a_n1672_n179.n41 199.788
R16967 a_n1672_n179.n24 a_n1672_n179.n23 185
R16968 a_n1672_n179.n22 a_n1672_n179.n2 185
R16969 a_n1672_n179.n12 a_n1672_n179.n11 185
R16970 a_n1672_n179.n7 a_n1672_n179.n21 187.962
R16971 a_n1672_n179.n34 a_n1672_n179.n33 185
R16972 a_n1672_n179.n32 a_n1672_n179.n4 185
R16973 a_n1672_n179.n14 a_n1672_n179.n13 185
R16974 a_n1672_n179.n8 a_n1672_n179.n31 187.962
R16975 a_n1672_n179.n19 a_n1672_n179.n18 185
R16976 a_n1672_n179.n45 a_n1672_n179.n6 185
R16977 a_n1672_n179.n5 a_n1672_n179.n46 185
R16978 a_n1672_n179.n10 a_n1672_n179.n17 187.962
R16979 a_n1672_n179.n23 a_n1672_n179.n22 104.615
R16980 a_n1672_n179.n22 a_n1672_n179.n11 104.615
R16981 a_n1672_n179.n21 a_n1672_n179.n11 104.615
R16982 a_n1672_n179.n33 a_n1672_n179.n32 104.615
R16983 a_n1672_n179.n32 a_n1672_n179.n13 104.615
R16984 a_n1672_n179.n31 a_n1672_n179.n13 104.615
R16985 a_n1672_n179.n45 a_n1672_n179.n18 104.615
R16986 a_n1672_n179.n46 a_n1672_n179.n45 104.615
R16987 a_n1672_n179.n46 a_n1672_n179.n17 104.615
R16988 a_n1672_n179.n15 a_n1672_n179.t0 64.3005
R16989 a_n1672_n179.n15 a_n1672_n179.t4 64.3003
R16990 a_n1672_n179.n39 a_n1672_n179.t12 64.3003
R16991 a_n1672_n179.n16 a_n1672_n179.t5 64.3003
R16992 a_n1672_n179.n15 a_n1672_n179.n27 59.5063
R16993 a_n1672_n179.n29 a_n1672_n179.n28 59.5063
R16994 a_n1672_n179.n16 a_n1672_n179.n38 59.5061
R16995 a_n1672_n179.n16 a_n1672_n179.n37 59.5061
R16996 a_n1672_n179.n21 a_n1672_n179.t9 52.3082
R16997 a_n1672_n179.n31 a_n1672_n179.t8 52.3082
R16998 a_n1672_n179.t10 a_n1672_n179.n17 52.3082
R16999 a_n1672_n179.n7 a_n1672_n179.n12 4.42678
R17000 a_n1672_n179.n8 a_n1672_n179.n14 4.42678
R17001 a_n1672_n179.n10 a_n1672_n179.n5 4.42678
R17002 a_n1672_n179.n2 a_n1672_n179.n12 12.0247
R17003 a_n1672_n179.n4 a_n1672_n179.n14 12.0247
R17004 a_n1672_n179.n6 a_n1672_n179.n5 12.0247
R17005 a_n1672_n179.n24 a_n1672_n179.n2 11.249
R17006 a_n1672_n179.n34 a_n1672_n179.n4 11.249
R17007 a_n1672_n179.n6 a_n1672_n179.n19 11.249
R17008 a_n1672_n179.n0 a_n1672_n179.n29 10.8929
R17009 a_n1672_n179.n25 a_n1672_n179.n20 10.4732
R17010 a_n1672_n179.n35 a_n1672_n179.n30 10.4732
R17011 a_n1672_n179.n44 a_n1672_n179.n43 10.4732
R17012 a_n1672_n179.n40 a_n1672_n179.n15 10.3476
R17013 a_n1672_n179.n26 a_n1672_n179.n1 9.45567
R17014 a_n1672_n179.n36 a_n1672_n179.n3 9.45567
R17015 a_n1672_n179.n9 a_n1672_n179.n42 9.45567
R17016 a_n1672_n179.n1 a_n1672_n179.n25 9.3005
R17017 a_n1672_n179.n3 a_n1672_n179.n35 9.3005
R17018 a_n1672_n179.n9 a_n1672_n179.n44 9.3005
R17019 a_n1672_n179.n16 a_n1672_n179.n0 5.98757
R17020 a_n1672_n179.n40 a_n1672_n179.n39 5.44231
R17021 a_n1672_n179.n38 a_n1672_n179.t6 4.79469
R17022 a_n1672_n179.n38 a_n1672_n179.t2 4.79469
R17023 a_n1672_n179.n37 a_n1672_n179.t14 4.79469
R17024 a_n1672_n179.n37 a_n1672_n179.t11 4.79469
R17025 a_n1672_n179.n27 a_n1672_n179.t3 4.79469
R17026 a_n1672_n179.n27 a_n1672_n179.t7 4.79469
R17027 a_n1672_n179.n28 a_n1672_n179.t1 4.79469
R17028 a_n1672_n179.n28 a_n1672_n179.t13 4.79469
R17029 a_n1672_n179.n1 a_n1672_n179.t9 150.207
R17030 a_n1672_n179.n3 a_n1672_n179.t8 150.207
R17031 a_n1672_n179.t10 a_n1672_n179.n9 150.207
R17032 a_n1672_n179.n6 a_n1672_n179.n9 11.2399
R17033 a_n1672_n179.n4 a_n1672_n179.n3 11.2399
R17034 a_n1672_n179.n2 a_n1672_n179.n1 11.2399
R17035 a_n1672_n179.n41 a_n1672_n179.n0 4.48834
R17036 a_n1672_n179.n9 a_n1672_n179.n10 2.42091
R17037 a_n1672_n179.n8 a_n1672_n179.n3 2.42091
R17038 a_n1672_n179.n7 a_n1672_n179.n1 2.42091
R17039 a_n1672_n179.n26 a_n1672_n179.n20 3.49141
R17040 a_n1672_n179.n36 a_n1672_n179.n30 3.49141
R17041 a_n1672_n179.n43 a_n1672_n179.n42 3.49141
R17042 a_n1672_n179.n41 a_n1672_n179.n40 3.06829
R17043 a_n1672_n179.n39 a_n1672_n179.n16 2.96171
R17044 a_n1672_n179.n29 a_n1672_n179.n15 2.96171
R17045 a_n1672_n179.n25 a_n1672_n179.n24 2.71565
R17046 a_n1672_n179.n35 a_n1672_n179.n34 2.71565
R17047 a_n1672_n179.n44 a_n1672_n179.n19 2.71565
R17048 CS_BIAS.n114 CS_BIAS.n113 161.3
R17049 CS_BIAS.n112 CS_BIAS.n95 161.3
R17050 CS_BIAS.n111 CS_BIAS.n110 161.3
R17051 CS_BIAS.n109 CS_BIAS.n96 161.3
R17052 CS_BIAS.n108 CS_BIAS.n107 161.3
R17053 CS_BIAS.n106 CS_BIAS.n97 161.3
R17054 CS_BIAS.n105 CS_BIAS.n104 161.3
R17055 CS_BIAS.n103 CS_BIAS.n98 161.3
R17056 CS_BIAS.n102 CS_BIAS.n101 161.3
R17057 CS_BIAS.n79 CS_BIAS.n78 161.3
R17058 CS_BIAS.n80 CS_BIAS.n75 161.3
R17059 CS_BIAS.n82 CS_BIAS.n81 161.3
R17060 CS_BIAS.n83 CS_BIAS.n74 161.3
R17061 CS_BIAS.n85 CS_BIAS.n84 161.3
R17062 CS_BIAS.n86 CS_BIAS.n73 161.3
R17063 CS_BIAS.n88 CS_BIAS.n87 161.3
R17064 CS_BIAS.n89 CS_BIAS.n72 161.3
R17065 CS_BIAS.n91 CS_BIAS.n90 161.3
R17066 CS_BIAS.n56 CS_BIAS.n55 161.3
R17067 CS_BIAS.n57 CS_BIAS.n52 161.3
R17068 CS_BIAS.n59 CS_BIAS.n58 161.3
R17069 CS_BIAS.n60 CS_BIAS.n51 161.3
R17070 CS_BIAS.n62 CS_BIAS.n61 161.3
R17071 CS_BIAS.n63 CS_BIAS.n50 161.3
R17072 CS_BIAS.n65 CS_BIAS.n64 161.3
R17073 CS_BIAS.n66 CS_BIAS.n49 161.3
R17074 CS_BIAS.n68 CS_BIAS.n67 161.3
R17075 CS_BIAS.n13 CS_BIAS.n12 161.3
R17076 CS_BIAS.n14 CS_BIAS.n9 161.3
R17077 CS_BIAS.n16 CS_BIAS.n15 161.3
R17078 CS_BIAS.n17 CS_BIAS.n8 161.3
R17079 CS_BIAS.n19 CS_BIAS.n18 161.3
R17080 CS_BIAS.n20 CS_BIAS.n7 161.3
R17081 CS_BIAS.n22 CS_BIAS.n21 161.3
R17082 CS_BIAS.n23 CS_BIAS.n6 161.3
R17083 CS_BIAS.n25 CS_BIAS.n24 161.3
R17084 CS_BIAS.n34 CS_BIAS.n33 161.3
R17085 CS_BIAS.n35 CS_BIAS.n4 161.3
R17086 CS_BIAS.n37 CS_BIAS.n36 161.3
R17087 CS_BIAS.n38 CS_BIAS.n3 161.3
R17088 CS_BIAS.n40 CS_BIAS.n39 161.3
R17089 CS_BIAS.n41 CS_BIAS.n2 161.3
R17090 CS_BIAS.n43 CS_BIAS.n42 161.3
R17091 CS_BIAS.n44 CS_BIAS.n1 161.3
R17092 CS_BIAS.n46 CS_BIAS.n45 161.3
R17093 CS_BIAS.n231 CS_BIAS.n230 161.3
R17094 CS_BIAS.n229 CS_BIAS.n212 161.3
R17095 CS_BIAS.n228 CS_BIAS.n227 161.3
R17096 CS_BIAS.n226 CS_BIAS.n213 161.3
R17097 CS_BIAS.n225 CS_BIAS.n224 161.3
R17098 CS_BIAS.n223 CS_BIAS.n214 161.3
R17099 CS_BIAS.n222 CS_BIAS.n221 161.3
R17100 CS_BIAS.n220 CS_BIAS.n215 161.3
R17101 CS_BIAS.n219 CS_BIAS.n218 161.3
R17102 CS_BIAS.n208 CS_BIAS.n207 161.3
R17103 CS_BIAS.n206 CS_BIAS.n189 161.3
R17104 CS_BIAS.n205 CS_BIAS.n204 161.3
R17105 CS_BIAS.n203 CS_BIAS.n190 161.3
R17106 CS_BIAS.n202 CS_BIAS.n201 161.3
R17107 CS_BIAS.n200 CS_BIAS.n191 161.3
R17108 CS_BIAS.n199 CS_BIAS.n198 161.3
R17109 CS_BIAS.n197 CS_BIAS.n192 161.3
R17110 CS_BIAS.n196 CS_BIAS.n195 161.3
R17111 CS_BIAS.n185 CS_BIAS.n184 161.3
R17112 CS_BIAS.n183 CS_BIAS.n166 161.3
R17113 CS_BIAS.n182 CS_BIAS.n181 161.3
R17114 CS_BIAS.n180 CS_BIAS.n167 161.3
R17115 CS_BIAS.n179 CS_BIAS.n178 161.3
R17116 CS_BIAS.n177 CS_BIAS.n168 161.3
R17117 CS_BIAS.n176 CS_BIAS.n175 161.3
R17118 CS_BIAS.n174 CS_BIAS.n169 161.3
R17119 CS_BIAS.n173 CS_BIAS.n172 161.3
R17120 CS_BIAS.n142 CS_BIAS.n141 161.3
R17121 CS_BIAS.n140 CS_BIAS.n123 161.3
R17122 CS_BIAS.n139 CS_BIAS.n138 161.3
R17123 CS_BIAS.n137 CS_BIAS.n124 161.3
R17124 CS_BIAS.n136 CS_BIAS.n135 161.3
R17125 CS_BIAS.n134 CS_BIAS.n125 161.3
R17126 CS_BIAS.n133 CS_BIAS.n132 161.3
R17127 CS_BIAS.n131 CS_BIAS.n126 161.3
R17128 CS_BIAS.n130 CS_BIAS.n129 161.3
R17129 CS_BIAS.n163 CS_BIAS.n162 161.3
R17130 CS_BIAS.n161 CS_BIAS.n118 161.3
R17131 CS_BIAS.n160 CS_BIAS.n159 161.3
R17132 CS_BIAS.n158 CS_BIAS.n119 161.3
R17133 CS_BIAS.n157 CS_BIAS.n156 161.3
R17134 CS_BIAS.n155 CS_BIAS.n120 161.3
R17135 CS_BIAS.n154 CS_BIAS.n153 161.3
R17136 CS_BIAS.n152 CS_BIAS.n121 161.3
R17137 CS_BIAS.n151 CS_BIAS.n150 161.3
R17138 CS_BIAS.n146 CS_BIAS.t1 99.5328
R17139 CS_BIAS.n27 CS_BIAS.t9 97.9229
R17140 CS_BIAS.n29 CS_BIAS.n28 92.77
R17141 CS_BIAS.n145 CS_BIAS.n144 92.2334
R17142 CS_BIAS.n115 CS_BIAS.n94 55.4214
R17143 CS_BIAS.n92 CS_BIAS.n71 55.4214
R17144 CS_BIAS.n69 CS_BIAS.n48 55.4214
R17145 CS_BIAS.n26 CS_BIAS.n5 55.4214
R17146 CS_BIAS.n47 CS_BIAS.n0 55.4214
R17147 CS_BIAS.n232 CS_BIAS.n211 55.4214
R17148 CS_BIAS.n209 CS_BIAS.n188 55.4214
R17149 CS_BIAS.n186 CS_BIAS.n165 55.4214
R17150 CS_BIAS.n143 CS_BIAS.n122 55.4214
R17151 CS_BIAS.n164 CS_BIAS.n117 55.4214
R17152 CS_BIAS.n32 CS_BIAS.n31 51.1899
R17153 CS_BIAS.n149 CS_BIAS.n148 51.1899
R17154 CS_BIAS.n77 CS_BIAS.n76 51.1859
R17155 CS_BIAS.n54 CS_BIAS.n53 51.1859
R17156 CS_BIAS.n11 CS_BIAS.n10 51.1859
R17157 CS_BIAS.n217 CS_BIAS.n216 51.1859
R17158 CS_BIAS.n194 CS_BIAS.n193 51.1859
R17159 CS_BIAS.n171 CS_BIAS.n170 51.1859
R17160 CS_BIAS.n128 CS_BIAS.n127 51.1859
R17161 CS_BIAS.n100 CS_BIAS.n99 51.1859
R17162 CS_BIAS.n99 CS_BIAS.t12 50.4863
R17163 CS_BIAS.n216 CS_BIAS.t29 50.4863
R17164 CS_BIAS.n193 CS_BIAS.t16 50.4863
R17165 CS_BIAS.n170 CS_BIAS.t19 50.4863
R17166 CS_BIAS.n127 CS_BIAS.t0 50.4863
R17167 CS_BIAS.n76 CS_BIAS.t23 50.4861
R17168 CS_BIAS.n53 CS_BIAS.t26 50.4861
R17169 CS_BIAS.n10 CS_BIAS.t10 50.4861
R17170 CS_BIAS.n148 CS_BIAS.t15 50.4803
R17171 CS_BIAS.n31 CS_BIAS.t18 50.4801
R17172 CS_BIAS.n107 CS_BIAS.n106 41.5458
R17173 CS_BIAS.n84 CS_BIAS.n83 41.5458
R17174 CS_BIAS.n61 CS_BIAS.n60 41.5458
R17175 CS_BIAS.n18 CS_BIAS.n17 41.5458
R17176 CS_BIAS.n39 CS_BIAS.n38 41.5458
R17177 CS_BIAS.n224 CS_BIAS.n223 41.5458
R17178 CS_BIAS.n201 CS_BIAS.n200 41.5458
R17179 CS_BIAS.n178 CS_BIAS.n177 41.5458
R17180 CS_BIAS.n135 CS_BIAS.n134 41.5458
R17181 CS_BIAS.n156 CS_BIAS.n155 41.5458
R17182 CS_BIAS.n107 CS_BIAS.n96 39.6083
R17183 CS_BIAS.n84 CS_BIAS.n73 39.6083
R17184 CS_BIAS.n61 CS_BIAS.n50 39.6083
R17185 CS_BIAS.n18 CS_BIAS.n7 39.6083
R17186 CS_BIAS.n39 CS_BIAS.n2 39.6083
R17187 CS_BIAS.n224 CS_BIAS.n213 39.6083
R17188 CS_BIAS.n201 CS_BIAS.n190 39.6083
R17189 CS_BIAS.n178 CS_BIAS.n167 39.6083
R17190 CS_BIAS.n135 CS_BIAS.n124 39.6083
R17191 CS_BIAS.n156 CS_BIAS.n119 39.6083
R17192 CS_BIAS.n106 CS_BIAS.n105 24.5923
R17193 CS_BIAS.n105 CS_BIAS.n98 24.5923
R17194 CS_BIAS.n101 CS_BIAS.n98 24.5923
R17195 CS_BIAS.n101 CS_BIAS.n100 24.5923
R17196 CS_BIAS.n113 CS_BIAS.n112 24.5923
R17197 CS_BIAS.n112 CS_BIAS.n111 24.5923
R17198 CS_BIAS.n111 CS_BIAS.n96 24.5923
R17199 CS_BIAS.n90 CS_BIAS.n89 24.5923
R17200 CS_BIAS.n89 CS_BIAS.n88 24.5923
R17201 CS_BIAS.n88 CS_BIAS.n73 24.5923
R17202 CS_BIAS.n83 CS_BIAS.n82 24.5923
R17203 CS_BIAS.n82 CS_BIAS.n75 24.5923
R17204 CS_BIAS.n78 CS_BIAS.n75 24.5923
R17205 CS_BIAS.n78 CS_BIAS.n77 24.5923
R17206 CS_BIAS.n67 CS_BIAS.n66 24.5923
R17207 CS_BIAS.n66 CS_BIAS.n65 24.5923
R17208 CS_BIAS.n65 CS_BIAS.n50 24.5923
R17209 CS_BIAS.n60 CS_BIAS.n59 24.5923
R17210 CS_BIAS.n59 CS_BIAS.n52 24.5923
R17211 CS_BIAS.n55 CS_BIAS.n52 24.5923
R17212 CS_BIAS.n55 CS_BIAS.n54 24.5923
R17213 CS_BIAS.n24 CS_BIAS.n23 24.5923
R17214 CS_BIAS.n23 CS_BIAS.n22 24.5923
R17215 CS_BIAS.n22 CS_BIAS.n7 24.5923
R17216 CS_BIAS.n17 CS_BIAS.n16 24.5923
R17217 CS_BIAS.n16 CS_BIAS.n9 24.5923
R17218 CS_BIAS.n12 CS_BIAS.n9 24.5923
R17219 CS_BIAS.n12 CS_BIAS.n11 24.5923
R17220 CS_BIAS.n45 CS_BIAS.n44 24.5923
R17221 CS_BIAS.n44 CS_BIAS.n43 24.5923
R17222 CS_BIAS.n43 CS_BIAS.n2 24.5923
R17223 CS_BIAS.n38 CS_BIAS.n37 24.5923
R17224 CS_BIAS.n37 CS_BIAS.n4 24.5923
R17225 CS_BIAS.n33 CS_BIAS.n4 24.5923
R17226 CS_BIAS.n33 CS_BIAS.n32 24.5923
R17227 CS_BIAS.n218 CS_BIAS.n217 24.5923
R17228 CS_BIAS.n218 CS_BIAS.n215 24.5923
R17229 CS_BIAS.n222 CS_BIAS.n215 24.5923
R17230 CS_BIAS.n223 CS_BIAS.n222 24.5923
R17231 CS_BIAS.n228 CS_BIAS.n213 24.5923
R17232 CS_BIAS.n229 CS_BIAS.n228 24.5923
R17233 CS_BIAS.n230 CS_BIAS.n229 24.5923
R17234 CS_BIAS.n195 CS_BIAS.n194 24.5923
R17235 CS_BIAS.n195 CS_BIAS.n192 24.5923
R17236 CS_BIAS.n199 CS_BIAS.n192 24.5923
R17237 CS_BIAS.n200 CS_BIAS.n199 24.5923
R17238 CS_BIAS.n205 CS_BIAS.n190 24.5923
R17239 CS_BIAS.n206 CS_BIAS.n205 24.5923
R17240 CS_BIAS.n207 CS_BIAS.n206 24.5923
R17241 CS_BIAS.n172 CS_BIAS.n171 24.5923
R17242 CS_BIAS.n172 CS_BIAS.n169 24.5923
R17243 CS_BIAS.n176 CS_BIAS.n169 24.5923
R17244 CS_BIAS.n177 CS_BIAS.n176 24.5923
R17245 CS_BIAS.n182 CS_BIAS.n167 24.5923
R17246 CS_BIAS.n183 CS_BIAS.n182 24.5923
R17247 CS_BIAS.n184 CS_BIAS.n183 24.5923
R17248 CS_BIAS.n129 CS_BIAS.n128 24.5923
R17249 CS_BIAS.n129 CS_BIAS.n126 24.5923
R17250 CS_BIAS.n133 CS_BIAS.n126 24.5923
R17251 CS_BIAS.n134 CS_BIAS.n133 24.5923
R17252 CS_BIAS.n139 CS_BIAS.n124 24.5923
R17253 CS_BIAS.n140 CS_BIAS.n139 24.5923
R17254 CS_BIAS.n141 CS_BIAS.n140 24.5923
R17255 CS_BIAS.n160 CS_BIAS.n119 24.5923
R17256 CS_BIAS.n161 CS_BIAS.n160 24.5923
R17257 CS_BIAS.n162 CS_BIAS.n161 24.5923
R17258 CS_BIAS.n150 CS_BIAS.n149 24.5923
R17259 CS_BIAS.n150 CS_BIAS.n121 24.5923
R17260 CS_BIAS.n154 CS_BIAS.n121 24.5923
R17261 CS_BIAS.n155 CS_BIAS.n154 24.5923
R17262 CS_BIAS.n113 CS_BIAS.n94 23.6087
R17263 CS_BIAS.n90 CS_BIAS.n71 23.6087
R17264 CS_BIAS.n67 CS_BIAS.n48 23.6087
R17265 CS_BIAS.n24 CS_BIAS.n5 23.6087
R17266 CS_BIAS.n45 CS_BIAS.n0 23.6087
R17267 CS_BIAS.n230 CS_BIAS.n211 23.6087
R17268 CS_BIAS.n207 CS_BIAS.n188 23.6087
R17269 CS_BIAS.n184 CS_BIAS.n165 23.6087
R17270 CS_BIAS.n141 CS_BIAS.n122 23.6087
R17271 CS_BIAS.n162 CS_BIAS.n117 23.6087
R17272 CS_BIAS.n100 CS_BIAS.t13 18.0366
R17273 CS_BIAS.n94 CS_BIAS.t22 18.0366
R17274 CS_BIAS.n77 CS_BIAS.t25 18.0366
R17275 CS_BIAS.n71 CS_BIAS.t30 18.0366
R17276 CS_BIAS.n54 CS_BIAS.t27 18.0366
R17277 CS_BIAS.n48 CS_BIAS.t34 18.0366
R17278 CS_BIAS.n11 CS_BIAS.t2 18.0366
R17279 CS_BIAS.n5 CS_BIAS.t8 18.0366
R17280 CS_BIAS.n32 CS_BIAS.t14 18.0366
R17281 CS_BIAS.n0 CS_BIAS.t28 18.0366
R17282 CS_BIAS.n217 CS_BIAS.t31 18.0366
R17283 CS_BIAS.n211 CS_BIAS.t33 18.0366
R17284 CS_BIAS.n194 CS_BIAS.t17 18.0366
R17285 CS_BIAS.n188 CS_BIAS.t20 18.0366
R17286 CS_BIAS.n171 CS_BIAS.t21 18.0366
R17287 CS_BIAS.n165 CS_BIAS.t24 18.0366
R17288 CS_BIAS.n128 CS_BIAS.t4 18.0366
R17289 CS_BIAS.n122 CS_BIAS.t6 18.0366
R17290 CS_BIAS.n149 CS_BIAS.t35 18.0366
R17291 CS_BIAS.n117 CS_BIAS.t32 18.0366
R17292 CS_BIAS.n145 CS_BIAS.n143 13.0441
R17293 CS_BIAS.n27 CS_BIAS.n26 11.9708
R17294 CS_BIAS.n30 CS_BIAS.n29 9.50363
R17295 CS_BIAS.n147 CS_BIAS.n146 9.50363
R17296 CS_BIAS.n234 CS_BIAS.n116 8.50759
R17297 CS_BIAS.n70 CS_BIAS.n47 7.74971
R17298 CS_BIAS.n187 CS_BIAS.n164 7.74971
R17299 CS_BIAS.n234 CS_BIAS.n233 6.82906
R17300 CS_BIAS.n28 CS_BIAS.t3 5.69016
R17301 CS_BIAS.n28 CS_BIAS.t11 5.69016
R17302 CS_BIAS.n144 CS_BIAS.t5 5.69016
R17303 CS_BIAS.n144 CS_BIAS.t7 5.69016
R17304 CS_BIAS.n116 CS_BIAS.n115 5.38986
R17305 CS_BIAS.n93 CS_BIAS.n92 5.38986
R17306 CS_BIAS.n70 CS_BIAS.n69 5.38986
R17307 CS_BIAS.n233 CS_BIAS.n232 5.38986
R17308 CS_BIAS.n210 CS_BIAS.n209 5.38986
R17309 CS_BIAS.n187 CS_BIAS.n186 5.38986
R17310 CS_BIAS CS_BIAS.n234 4.39923
R17311 CS_BIAS.n116 CS_BIAS.n93 2.36035
R17312 CS_BIAS.n233 CS_BIAS.n210 2.36035
R17313 CS_BIAS.n93 CS_BIAS.n70 2.35656
R17314 CS_BIAS.n210 CS_BIAS.n187 2.35656
R17315 CS_BIAS.n29 CS_BIAS.n27 1.61041
R17316 CS_BIAS.n219 CS_BIAS.n216 1.44731
R17317 CS_BIAS.n196 CS_BIAS.n193 1.44731
R17318 CS_BIAS.n173 CS_BIAS.n170 1.44731
R17319 CS_BIAS.n130 CS_BIAS.n127 1.44731
R17320 CS_BIAS.n102 CS_BIAS.n99 1.44731
R17321 CS_BIAS.n79 CS_BIAS.n76 1.44731
R17322 CS_BIAS.n56 CS_BIAS.n53 1.44731
R17323 CS_BIAS.n13 CS_BIAS.n10 1.44731
R17324 CS_BIAS.n148 CS_BIAS.n147 1.24524
R17325 CS_BIAS.n31 CS_BIAS.n30 1.24523
R17326 CS_BIAS.n146 CS_BIAS.n145 0.537138
R17327 CS_BIAS.n115 CS_BIAS.n114 0.46582
R17328 CS_BIAS.n92 CS_BIAS.n91 0.46582
R17329 CS_BIAS.n69 CS_BIAS.n68 0.46582
R17330 CS_BIAS.n26 CS_BIAS.n25 0.46582
R17331 CS_BIAS.n47 CS_BIAS.n46 0.46582
R17332 CS_BIAS.n232 CS_BIAS.n231 0.46582
R17333 CS_BIAS.n209 CS_BIAS.n208 0.46582
R17334 CS_BIAS.n186 CS_BIAS.n185 0.46582
R17335 CS_BIAS.n143 CS_BIAS.n142 0.46582
R17336 CS_BIAS.n164 CS_BIAS.n163 0.46582
R17337 CS_BIAS.n114 CS_BIAS.n95 0.189894
R17338 CS_BIAS.n110 CS_BIAS.n95 0.189894
R17339 CS_BIAS.n110 CS_BIAS.n109 0.189894
R17340 CS_BIAS.n109 CS_BIAS.n108 0.189894
R17341 CS_BIAS.n108 CS_BIAS.n97 0.189894
R17342 CS_BIAS.n104 CS_BIAS.n97 0.189894
R17343 CS_BIAS.n104 CS_BIAS.n103 0.189894
R17344 CS_BIAS.n103 CS_BIAS.n102 0.189894
R17345 CS_BIAS.n91 CS_BIAS.n72 0.189894
R17346 CS_BIAS.n87 CS_BIAS.n72 0.189894
R17347 CS_BIAS.n87 CS_BIAS.n86 0.189894
R17348 CS_BIAS.n86 CS_BIAS.n85 0.189894
R17349 CS_BIAS.n85 CS_BIAS.n74 0.189894
R17350 CS_BIAS.n81 CS_BIAS.n74 0.189894
R17351 CS_BIAS.n81 CS_BIAS.n80 0.189894
R17352 CS_BIAS.n80 CS_BIAS.n79 0.189894
R17353 CS_BIAS.n68 CS_BIAS.n49 0.189894
R17354 CS_BIAS.n64 CS_BIAS.n49 0.189894
R17355 CS_BIAS.n64 CS_BIAS.n63 0.189894
R17356 CS_BIAS.n63 CS_BIAS.n62 0.189894
R17357 CS_BIAS.n62 CS_BIAS.n51 0.189894
R17358 CS_BIAS.n58 CS_BIAS.n51 0.189894
R17359 CS_BIAS.n58 CS_BIAS.n57 0.189894
R17360 CS_BIAS.n57 CS_BIAS.n56 0.189894
R17361 CS_BIAS.n25 CS_BIAS.n6 0.189894
R17362 CS_BIAS.n21 CS_BIAS.n6 0.189894
R17363 CS_BIAS.n21 CS_BIAS.n20 0.189894
R17364 CS_BIAS.n20 CS_BIAS.n19 0.189894
R17365 CS_BIAS.n19 CS_BIAS.n8 0.189894
R17366 CS_BIAS.n15 CS_BIAS.n8 0.189894
R17367 CS_BIAS.n15 CS_BIAS.n14 0.189894
R17368 CS_BIAS.n14 CS_BIAS.n13 0.189894
R17369 CS_BIAS.n46 CS_BIAS.n1 0.189894
R17370 CS_BIAS.n42 CS_BIAS.n1 0.189894
R17371 CS_BIAS.n42 CS_BIAS.n41 0.189894
R17372 CS_BIAS.n41 CS_BIAS.n40 0.189894
R17373 CS_BIAS.n40 CS_BIAS.n3 0.189894
R17374 CS_BIAS.n36 CS_BIAS.n3 0.189894
R17375 CS_BIAS.n36 CS_BIAS.n35 0.189894
R17376 CS_BIAS.n35 CS_BIAS.n34 0.189894
R17377 CS_BIAS.n220 CS_BIAS.n219 0.189894
R17378 CS_BIAS.n221 CS_BIAS.n220 0.189894
R17379 CS_BIAS.n221 CS_BIAS.n214 0.189894
R17380 CS_BIAS.n225 CS_BIAS.n214 0.189894
R17381 CS_BIAS.n226 CS_BIAS.n225 0.189894
R17382 CS_BIAS.n227 CS_BIAS.n226 0.189894
R17383 CS_BIAS.n227 CS_BIAS.n212 0.189894
R17384 CS_BIAS.n231 CS_BIAS.n212 0.189894
R17385 CS_BIAS.n197 CS_BIAS.n196 0.189894
R17386 CS_BIAS.n198 CS_BIAS.n197 0.189894
R17387 CS_BIAS.n198 CS_BIAS.n191 0.189894
R17388 CS_BIAS.n202 CS_BIAS.n191 0.189894
R17389 CS_BIAS.n203 CS_BIAS.n202 0.189894
R17390 CS_BIAS.n204 CS_BIAS.n203 0.189894
R17391 CS_BIAS.n204 CS_BIAS.n189 0.189894
R17392 CS_BIAS.n208 CS_BIAS.n189 0.189894
R17393 CS_BIAS.n174 CS_BIAS.n173 0.189894
R17394 CS_BIAS.n175 CS_BIAS.n174 0.189894
R17395 CS_BIAS.n175 CS_BIAS.n168 0.189894
R17396 CS_BIAS.n179 CS_BIAS.n168 0.189894
R17397 CS_BIAS.n180 CS_BIAS.n179 0.189894
R17398 CS_BIAS.n181 CS_BIAS.n180 0.189894
R17399 CS_BIAS.n181 CS_BIAS.n166 0.189894
R17400 CS_BIAS.n185 CS_BIAS.n166 0.189894
R17401 CS_BIAS.n131 CS_BIAS.n130 0.189894
R17402 CS_BIAS.n132 CS_BIAS.n131 0.189894
R17403 CS_BIAS.n132 CS_BIAS.n125 0.189894
R17404 CS_BIAS.n136 CS_BIAS.n125 0.189894
R17405 CS_BIAS.n137 CS_BIAS.n136 0.189894
R17406 CS_BIAS.n138 CS_BIAS.n137 0.189894
R17407 CS_BIAS.n138 CS_BIAS.n123 0.189894
R17408 CS_BIAS.n142 CS_BIAS.n123 0.189894
R17409 CS_BIAS.n152 CS_BIAS.n151 0.189894
R17410 CS_BIAS.n153 CS_BIAS.n152 0.189894
R17411 CS_BIAS.n153 CS_BIAS.n120 0.189894
R17412 CS_BIAS.n157 CS_BIAS.n120 0.189894
R17413 CS_BIAS.n158 CS_BIAS.n157 0.189894
R17414 CS_BIAS.n159 CS_BIAS.n158 0.189894
R17415 CS_BIAS.n159 CS_BIAS.n118 0.189894
R17416 CS_BIAS.n163 CS_BIAS.n118 0.189894
R17417 CS_BIAS.n34 CS_BIAS.n30 0.170955
R17418 CS_BIAS.n151 CS_BIAS.n147 0.170955
R17419 VOUT.n37 VOUT.n35 756.745
R17420 VOUT.n28 VOUT.n26 756.745
R17421 VOUT.n12 VOUT.n10 756.745
R17422 VOUT.n3 VOUT.n1 756.745
R17423 VOUT.n38 VOUT.n37 585
R17424 VOUT.n29 VOUT.n28 585
R17425 VOUT.n13 VOUT.n12 585
R17426 VOUT.n4 VOUT.n3 585
R17427 VOUT.t5 VOUT.n36 417.779
R17428 VOUT.t6 VOUT.n27 417.779
R17429 VOUT.t8 VOUT.n11 417.779
R17430 VOUT.t9 VOUT.n2 417.779
R17431 VOUT.n17 VOUT.n9 220.571
R17432 VOUT.n8 VOUT.n0 220.571
R17433 VOUT.n43 VOUT.n42 217.898
R17434 VOUT.n34 VOUT.n33 217.898
R17435 VOUT.n55 VOUT.t25 100.07
R17436 VOUT.n52 VOUT.t17 100.07
R17437 VOUT.n49 VOUT.t13 100.07
R17438 VOUT.n47 VOUT.t19 100.07
R17439 VOUT.n67 VOUT.t18 97.9229
R17440 VOUT.n64 VOUT.t31 97.9229
R17441 VOUT.n61 VOUT.t28 97.9229
R17442 VOUT.n59 VOUT.t32 97.9229
R17443 VOUT.n67 VOUT.n66 94.3799
R17444 VOUT.n64 VOUT.n63 94.3799
R17445 VOUT.n61 VOUT.n60 94.3799
R17446 VOUT.n59 VOUT.n58 94.3799
R17447 VOUT.n55 VOUT.n54 92.2334
R17448 VOUT.n52 VOUT.n51 92.2334
R17449 VOUT.n49 VOUT.n48 92.2334
R17450 VOUT.n47 VOUT.n46 92.2334
R17451 VOUT.n37 VOUT.t5 85.8723
R17452 VOUT.n28 VOUT.t6 85.8723
R17453 VOUT.n12 VOUT.t8 85.8723
R17454 VOUT.n3 VOUT.t9 85.8723
R17455 VOUT.n43 VOUT.n41 67.8275
R17456 VOUT.n34 VOUT.n32 67.8275
R17457 VOUT.n17 VOUT.n16 65.155
R17458 VOUT.n8 VOUT.n7 65.155
R17459 VOUT.n42 VOUT.t0 16.1721
R17460 VOUT.n42 VOUT.t3 16.1721
R17461 VOUT.n33 VOUT.t2 16.1721
R17462 VOUT.n33 VOUT.t11 16.1721
R17463 VOUT.n9 VOUT.t4 16.1721
R17464 VOUT.n9 VOUT.t1 16.1721
R17465 VOUT.n0 VOUT.t7 16.1721
R17466 VOUT.n0 VOUT.t10 16.1721
R17467 VOUT.n38 VOUT.n36 9.84608
R17468 VOUT.n29 VOUT.n27 9.84608
R17469 VOUT.n13 VOUT.n11 9.84608
R17470 VOUT.n4 VOUT.n2 9.84608
R17471 VOUT.n41 VOUT.n40 9.45567
R17472 VOUT.n32 VOUT.n31 9.45567
R17473 VOUT.n16 VOUT.n15 9.45567
R17474 VOUT.n7 VOUT.n6 9.45567
R17475 VOUT.n40 VOUT.n39 9.3005
R17476 VOUT.n31 VOUT.n30 9.3005
R17477 VOUT.n15 VOUT.n14 9.3005
R17478 VOUT.n6 VOUT.n5 9.3005
R17479 VOUT.n57 VOUT.n45 9.11273
R17480 VOUT.n41 VOUT.n35 8.14595
R17481 VOUT.n32 VOUT.n26 8.14595
R17482 VOUT.n16 VOUT.n10 8.14595
R17483 VOUT.n7 VOUT.n1 8.14595
R17484 VOUT.n50 VOUT.n47 7.40352
R17485 VOUT.n39 VOUT.n38 7.3702
R17486 VOUT.n30 VOUT.n29 7.3702
R17487 VOUT.n14 VOUT.n13 7.3702
R17488 VOUT.n5 VOUT.n4 7.3702
R17489 VOUT.n44 VOUT.n34 7.34964
R17490 VOUT.n45 VOUT.n44 6.47192
R17491 VOUT.n19 VOUT.n18 6.47192
R17492 VOUT.n62 VOUT.n59 6.33024
R17493 VOUT.n44 VOUT.n43 6.30222
R17494 VOUT.n56 VOUT.n55 6.03929
R17495 VOUT.n53 VOUT.n52 6.03929
R17496 VOUT.n50 VOUT.n49 6.03929
R17497 VOUT.n18 VOUT.n8 6.01343
R17498 VOUT.n39 VOUT.n35 5.81868
R17499 VOUT.n30 VOUT.n26 5.81868
R17500 VOUT.n14 VOUT.n10 5.81868
R17501 VOUT.n5 VOUT.n1 5.81868
R17502 VOUT.n54 VOUT.t34 5.69016
R17503 VOUT.n54 VOUT.t35 5.69016
R17504 VOUT.n51 VOUT.t22 5.69016
R17505 VOUT.n51 VOUT.t24 5.69016
R17506 VOUT.n48 VOUT.t20 5.69016
R17507 VOUT.n48 VOUT.t21 5.69016
R17508 VOUT.n46 VOUT.t33 5.69016
R17509 VOUT.n46 VOUT.t29 5.69016
R17510 VOUT.n66 VOUT.t16 5.69016
R17511 VOUT.n66 VOUT.t14 5.69016
R17512 VOUT.n63 VOUT.t30 5.69016
R17513 VOUT.n63 VOUT.t27 5.69016
R17514 VOUT.n60 VOUT.t26 5.69016
R17515 VOUT.n60 VOUT.t23 5.69016
R17516 VOUT.n58 VOUT.t12 5.69016
R17517 VOUT.n58 VOUT.t15 5.69016
R17518 VOUT.n18 VOUT.n17 4.96602
R17519 VOUT.n68 VOUT.n67 4.96602
R17520 VOUT.n65 VOUT.n64 4.96602
R17521 VOUT.n62 VOUT.n61 4.96602
R17522 VOUT.n70 VOUT.n19 4.7639
R17523 VOUT.n57 VOUT.n56 4.76287
R17524 VOUT.n69 VOUT.n68 4.76287
R17525 VOUT.n70 VOUT.n69 4.32982
R17526 VOUT.n25 VOUT 4.1083
R17527 VOUT.n45 VOUT.n19 3.93064
R17528 VOUT.n40 VOUT.n36 3.32369
R17529 VOUT.n31 VOUT.n27 3.32369
R17530 VOUT.n15 VOUT.n11 3.32369
R17531 VOUT.n6 VOUT.n2 3.32369
R17532 VOUT.n69 VOUT.n57 2.72587
R17533 VOUT.n56 VOUT.n53 1.36472
R17534 VOUT.n68 VOUT.n65 1.36472
R17535 VOUT.n53 VOUT.n50 1.36257
R17536 VOUT.n65 VOUT.n62 1.36257
R17537 VOUT.n70 VOUT.n25 0.40188
R17538 VOUT.n25 VOUT.n24 0.384144
R17539 VOUT.n23 VOUT.n22 0.104763
R17540 VOUT.n21 VOUT.n20 0.104763
R17541 VOUT.n22 VOUT.n21 0.0585126
R17542 VOUT.n24 VOUT.n20 0.0525046
R17543 VOUT.n20 VOUT.t38 0.0227451
R17544 VOUT.n23 VOUT.t39 0.0227451
R17545 VOUT.n21 VOUT.t36 0.022001
R17546 VOUT.n22 VOUT.t37 0.022001
R17547 VOUT.n24 VOUT.n23 0.0138602
R17548 VOUT VOUT.n70 0.0099
R17549 VP.n34 VP.t3 243.255
R17550 VP.n31 VP.n29 224.169
R17551 VP.n33 VP.n32 223.454
R17552 VP.n31 VP.n30 223.454
R17553 VP.n19 VP.n16 161.3
R17554 VP.n21 VP.n20 161.3
R17555 VP.n22 VP.n15 161.3
R17556 VP.n24 VP.n23 161.3
R17557 VP.n25 VP.n14 161.3
R17558 VP.n11 VP.n0 161.3
R17559 VP.n10 VP.n9 161.3
R17560 VP.n8 VP.n1 161.3
R17561 VP.n7 VP.n6 161.3
R17562 VP.n5 VP.n2 161.3
R17563 VP.n27 VP.n26 97.0549
R17564 VP.n13 VP.n12 97.0549
R17565 VP.n17 VP.t10 77.6701
R17566 VP.n3 VP.t7 77.6701
R17567 VP.n18 VP.n17 59.2585
R17568 VP.n4 VP.n3 59.2585
R17569 VP.n26 VP.t8 45.2428
R17570 VP.n18 VP.t11 45.2428
R17571 VP.n4 VP.t9 45.2428
R17572 VP.n12 VP.t12 45.2428
R17573 VP.n24 VP.n15 41.9503
R17574 VP.n10 VP.n1 41.9503
R17575 VP.n20 VP.n15 39.0365
R17576 VP.n6 VP.n1 39.0365
R17577 VP.n28 VP.n27 30.4489
R17578 VP.n25 VP.n24 24.4675
R17579 VP.n20 VP.n19 24.4675
R17580 VP.n6 VP.n5 24.4675
R17581 VP.n11 VP.n10 24.4675
R17582 VP.n32 VP.t1 19.8005
R17583 VP.n32 VP.t5 19.8005
R17584 VP.n30 VP.t0 19.8005
R17585 VP.n30 VP.t4 19.8005
R17586 VP.n29 VP.t2 19.8005
R17587 VP.n29 VP.t6 19.8005
R17588 VP.n26 VP.n25 13.702
R17589 VP.n12 VP.n11 13.702
R17590 VP VP.n35 12.7615
R17591 VP.n19 VP.n18 12.234
R17592 VP.n5 VP.n4 12.234
R17593 VP.n28 VP.n13 11.6232
R17594 VP.n17 VP.n16 9.58252
R17595 VP.n3 VP.n2 9.58252
R17596 VP.n35 VP.n34 4.80222
R17597 VP.n35 VP.n28 0.972091
R17598 VP.n33 VP.n31 0.716017
R17599 VP.n34 VP.n33 0.716017
R17600 VP.n27 VP.n14 0.278367
R17601 VP.n13 VP.n0 0.278367
R17602 VP.n23 VP.n14 0.189894
R17603 VP.n23 VP.n22 0.189894
R17604 VP.n22 VP.n21 0.189894
R17605 VP.n21 VP.n16 0.189894
R17606 VP.n7 VP.n2 0.189894
R17607 VP.n8 VP.n7 0.189894
R17608 VP.n9 VP.n8 0.189894
R17609 VP.n9 VP.n0 0.189894
R17610 VN.n30 VN.t3 243.97
R17611 VN.n30 VN.n29 223.454
R17612 VN.n32 VN.n31 223.454
R17613 VN.n34 VN.n33 223.454
R17614 VN.n25 VN.n14 161.3
R17615 VN.n24 VN.n23 161.3
R17616 VN.n22 VN.n15 161.3
R17617 VN.n21 VN.n20 161.3
R17618 VN.n19 VN.n16 161.3
R17619 VN.n5 VN.n2 161.3
R17620 VN.n7 VN.n6 161.3
R17621 VN.n8 VN.n1 161.3
R17622 VN.n10 VN.n9 161.3
R17623 VN.n11 VN.n0 161.3
R17624 VN.n27 VN.n26 97.0549
R17625 VN.n13 VN.n12 97.0549
R17626 VN.n17 VN.t10 77.6701
R17627 VN.n3 VN.t7 77.6701
R17628 VN.n18 VN.n17 59.2585
R17629 VN.n4 VN.n3 59.2585
R17630 VN.n18 VN.t12 45.2428
R17631 VN.n26 VN.t9 45.2428
R17632 VN.n12 VN.t11 45.2428
R17633 VN.n4 VN.t8 45.2428
R17634 VN.n24 VN.n15 41.9503
R17635 VN.n10 VN.n1 41.9503
R17636 VN.n20 VN.n15 39.0365
R17637 VN.n6 VN.n1 39.0365
R17638 VN.n28 VN.n27 30.233
R17639 VN.n20 VN.n19 24.4675
R17640 VN.n25 VN.n24 24.4675
R17641 VN.n11 VN.n10 24.4675
R17642 VN.n6 VN.n5 24.4675
R17643 VN.n29 VN.t5 19.8005
R17644 VN.n29 VN.t2 19.8005
R17645 VN.n31 VN.t6 19.8005
R17646 VN.n31 VN.t0 19.8005
R17647 VN.n33 VN.t4 19.8005
R17648 VN.n33 VN.t1 19.8005
R17649 VN VN.n35 15.515
R17650 VN.n26 VN.n25 13.702
R17651 VN.n12 VN.n11 13.702
R17652 VN.n19 VN.n18 12.234
R17653 VN.n5 VN.n4 12.234
R17654 VN.n28 VN.n13 11.4072
R17655 VN.n17 VN.n16 9.58252
R17656 VN.n3 VN.n2 9.58252
R17657 VN.n35 VN.n34 5.40567
R17658 VN.n35 VN.n28 1.188
R17659 VN.n34 VN.n32 0.716017
R17660 VN.n32 VN.n30 0.716017
R17661 VN.n27 VN.n14 0.278367
R17662 VN.n13 VN.n0 0.278367
R17663 VN.n21 VN.n16 0.189894
R17664 VN.n22 VN.n21 0.189894
R17665 VN.n23 VN.n22 0.189894
R17666 VN.n23 VN.n14 0.189894
R17667 VN.n9 VN.n0 0.189894
R17668 VN.n9 VN.n8 0.189894
R17669 VN.n8 VN.n7 0.189894
R17670 VN.n7 VN.n2 0.189894
R17671 a_n5082_9332.n7 a_n5082_9332.n5 127.225
R17672 a_n5082_9332.n10 a_n5082_9332.n8 126.522
R17673 a_n5082_9332.n10 a_n5082_9332.n9 126.035
R17674 a_n5082_9332.n7 a_n5082_9332.n6 126.034
R17675 a_n5082_9332.n2 a_n5082_9332.t5 106.963
R17676 a_n5082_9332.n0 a_n5082_9332.t3 105.775
R17677 a_n5082_9332.n0 a_n5082_9332.t1 105.775
R17678 a_n5082_9332.t7 a_n5082_9332.n12 105.775
R17679 a_n5082_9332.n4 a_n5082_9332.n3 98.1078
R17680 a_n5082_9332.n2 a_n5082_9332.n1 98.1078
R17681 a_n5082_9332.n11 a_n5082_9332.n10 15.4513
R17682 a_n5082_9332.n11 a_n5082_9332.n7 11.5663
R17683 a_n5082_9332.n3 a_n5082_9332.t6 7.66677
R17684 a_n5082_9332.n3 a_n5082_9332.t4 7.66677
R17685 a_n5082_9332.n1 a_n5082_9332.t0 7.66677
R17686 a_n5082_9332.n1 a_n5082_9332.t2 7.66677
R17687 a_n5082_9332.n6 a_n5082_9332.t13 7.66677
R17688 a_n5082_9332.n6 a_n5082_9332.t15 7.66677
R17689 a_n5082_9332.n5 a_n5082_9332.t10 7.66677
R17690 a_n5082_9332.n5 a_n5082_9332.t12 7.66677
R17691 a_n5082_9332.n9 a_n5082_9332.t11 7.66677
R17692 a_n5082_9332.n9 a_n5082_9332.t14 7.66677
R17693 a_n5082_9332.n8 a_n5082_9332.t8 7.66677
R17694 a_n5082_9332.n8 a_n5082_9332.t9 7.66677
R17695 a_n5082_9332.n12 a_n5082_9332.n11 5.59964
R17696 a_n5082_9332.n4 a_n5082_9332.n0 1.49727
R17697 a_n5082_9332.n0 a_n5082_9332.n2 1.19016
R17698 a_n5082_9332.n12 a_n5082_9332.n4 1.19016
C0 VOUT CS_BIAS 21.899302f
C1 VP VN 9.77428f
C2 VP CS_BIAS 0.324737f
C3 VP DIFFPAIR_BIAS 1.21e-19
C4 VN CS_BIAS 0.282762f
C5 VN DIFFPAIR_BIAS 1.21e-19
C6 a_5210_9332# VDD 1.13464f
C7 VDD VOUT 26.464499f
C8 VDD VN 0.094261f
C9 VOUT VP 3.76645f
C10 a_n5852_9332# VDD 1.13464f
C11 VOUT VN 0.918274f
C12 DIFFPAIR_BIAS GND 29.168999f
C13 CS_BIAS GND 0.111176p
C14 VN GND 31.555141f
C15 VP GND 28.357391f
C16 VOUT GND 72.67107f
C17 VDD GND 0.477464p
C18 a_5210_9332# GND 0.319159f
C19 a_n5852_9332# GND 0.319159f
C20 a_n5082_9332.n0 GND 1.85862f
C21 a_n5082_9332.t5 GND 0.669736f
C22 a_n5082_9332.t0 GND 0.085968f
C23 a_n5082_9332.t2 GND 0.085968f
C24 a_n5082_9332.n1 GND 0.470721f
C25 a_n5082_9332.n2 GND 2.01526f
C26 a_n5082_9332.t1 GND 0.6603f
C27 a_n5082_9332.t3 GND 0.6603f
C28 a_n5082_9332.t6 GND 0.085968f
C29 a_n5082_9332.t4 GND 0.085968f
C30 a_n5082_9332.n3 GND 0.470721f
C31 a_n5082_9332.n4 GND 1.17629f
C32 a_n5082_9332.t10 GND 0.085968f
C33 a_n5082_9332.t12 GND 0.085968f
C34 a_n5082_9332.n5 GND 0.577113f
C35 a_n5082_9332.t13 GND 0.085968f
C36 a_n5082_9332.t15 GND 0.085968f
C37 a_n5082_9332.n6 GND 0.566266f
C38 a_n5082_9332.n7 GND 3.9267f
C39 a_n5082_9332.t8 GND 0.085968f
C40 a_n5082_9332.t9 GND 0.085968f
C41 a_n5082_9332.n8 GND 0.575214f
C42 a_n5082_9332.t11 GND 0.085968f
C43 a_n5082_9332.t14 GND 0.085968f
C44 a_n5082_9332.n9 GND 0.566268f
C45 a_n5082_9332.n10 GND 8.518459f
C46 a_n5082_9332.n11 GND 3.08814f
C47 a_n5082_9332.n12 GND 1.50799f
C48 a_n5082_9332.t7 GND 0.6603f
C49 VN.n0 GND 0.02021f
C50 VN.t11 GND 0.358822f
C51 VN.n1 GND 0.012437f
C52 VN.n2 GND 0.130484f
C53 VN.t8 GND 0.358822f
C54 VN.t7 GND 0.453311f
C55 VN.n3 GND 0.178564f
C56 VN.n4 GND 0.183761f
C57 VN.n5 GND 0.021517f
C58 VN.n6 GND 0.030675f
C59 VN.n7 GND 0.015329f
C60 VN.n8 GND 0.015329f
C61 VN.n9 GND 0.015329f
C62 VN.n10 GND 0.030215f
C63 VN.n11 GND 0.022363f
C64 VN.n12 GND 0.190308f
C65 VN.n13 GND 0.19251f
C66 VN.n14 GND 0.02021f
C67 VN.t9 GND 0.358822f
C68 VN.n15 GND 0.012437f
C69 VN.n16 GND 0.130484f
C70 VN.t12 GND 0.358822f
C71 VN.t10 GND 0.453311f
C72 VN.n17 GND 0.178564f
C73 VN.n18 GND 0.183761f
C74 VN.n19 GND 0.021517f
C75 VN.n20 GND 0.030675f
C76 VN.n21 GND 0.015329f
C77 VN.n22 GND 0.015329f
C78 VN.n23 GND 0.015329f
C79 VN.n24 GND 0.030215f
C80 VN.n25 GND 0.022363f
C81 VN.n26 GND 0.190308f
C82 VN.n27 GND 0.460268f
C83 VN.n28 GND 0.648622f
C84 VN.t3 GND 0.026462f
C85 VN.t5 GND 0.004725f
C86 VN.t2 GND 0.004725f
C87 VN.n29 GND 0.015325f
C88 VN.n30 GND 0.118973f
C89 VN.t6 GND 0.004725f
C90 VN.t0 GND 0.004725f
C91 VN.n31 GND 0.015325f
C92 VN.n32 GND 0.0643f
C93 VN.t4 GND 0.004725f
C94 VN.t1 GND 0.004725f
C95 VN.n33 GND 0.015325f
C96 VN.n34 GND 0.089304f
C97 VN.n35 GND 2.26394f
C98 VP.n0 GND 0.030216f
C99 VP.t12 GND 0.53649f
C100 VP.n1 GND 0.018595f
C101 VP.n2 GND 0.195092f
C102 VP.t9 GND 0.53649f
C103 VP.t7 GND 0.677763f
C104 VP.n3 GND 0.266979f
C105 VP.n4 GND 0.274748f
C106 VP.n5 GND 0.032171f
C107 VP.n6 GND 0.045863f
C108 VP.n7 GND 0.022919f
C109 VP.n8 GND 0.022919f
C110 VP.n9 GND 0.022919f
C111 VP.n10 GND 0.045176f
C112 VP.n11 GND 0.033436f
C113 VP.n12 GND 0.284538f
C114 VP.n13 GND 0.293233f
C115 VP.n14 GND 0.030216f
C116 VP.t8 GND 0.53649f
C117 VP.n15 GND 0.018595f
C118 VP.n16 GND 0.195092f
C119 VP.t11 GND 0.53649f
C120 VP.t10 GND 0.677763f
C121 VP.n17 GND 0.266979f
C122 VP.n18 GND 0.274748f
C123 VP.n19 GND 0.032171f
C124 VP.n20 GND 0.045863f
C125 VP.n21 GND 0.022919f
C126 VP.n22 GND 0.022919f
C127 VP.n23 GND 0.022919f
C128 VP.n24 GND 0.045176f
C129 VP.n25 GND 0.033436f
C130 VP.n26 GND 0.284538f
C131 VP.n27 GND 0.69735f
C132 VP.n28 GND 0.979357f
C133 VP.t2 GND 0.007065f
C134 VP.t6 GND 0.007065f
C135 VP.n29 GND 0.023232f
C136 VP.t0 GND 0.007065f
C137 VP.t4 GND 0.007065f
C138 VP.n30 GND 0.022914f
C139 VP.n31 GND 0.195559f
C140 VP.t1 GND 0.007065f
C141 VP.t5 GND 0.007065f
C142 VP.n32 GND 0.022914f
C143 VP.n33 GND 0.096138f
C144 VP.t3 GND 0.039324f
C145 VP.n34 GND 0.106715f
C146 VP.n35 GND 2.14156f
C147 VOUT.t7 GND 0.008839f
C148 VOUT.t10 GND 0.008839f
C149 VOUT.n0 GND 0.047467f
C150 VOUT.n1 GND 0.006304f
C151 VOUT.n2 GND 0.016282f
C152 VOUT.t9 GND 0.016345f
C153 VOUT.n3 GND 0.015988f
C154 VOUT.n4 GND 0.00461f
C155 VOUT.n5 GND 0.00299f
C156 VOUT.n6 GND 0.038717f
C157 VOUT.n7 GND 0.016652f
C158 VOUT.n8 GND 0.734711f
C159 VOUT.t4 GND 0.008839f
C160 VOUT.t1 GND 0.008839f
C161 VOUT.n9 GND 0.047467f
C162 VOUT.n10 GND 0.006304f
C163 VOUT.n11 GND 0.016282f
C164 VOUT.t8 GND 0.016345f
C165 VOUT.n12 GND 0.015988f
C166 VOUT.n13 GND 0.00461f
C167 VOUT.n14 GND 0.00299f
C168 VOUT.n15 GND 0.038717f
C169 VOUT.n16 GND 0.016652f
C170 VOUT.n17 GND 0.719812f
C171 VOUT.n18 GND 0.543533f
C172 VOUT.n19 GND 6.52408f
C173 VOUT.t38 GND 9.118389f
C174 VOUT.n20 GND 6.58776f
C175 VOUT.t39 GND 9.118389f
C176 VOUT.t37 GND 9.28858f
C177 VOUT.t36 GND 9.28858f
C178 VOUT.n21 GND 7.38645f
C179 VOUT.n22 GND 7.38645f
C180 VOUT.n23 GND 3.21162f
C181 VOUT.n24 GND 7.45934f
C182 VOUT.n25 GND 1.75621f
C183 VOUT.n26 GND 0.006304f
C184 VOUT.n27 GND 0.016282f
C185 VOUT.t6 GND 0.016345f
C186 VOUT.n28 GND 0.015988f
C187 VOUT.n29 GND 0.00461f
C188 VOUT.n30 GND 0.00299f
C189 VOUT.n31 GND 0.038717f
C190 VOUT.n32 GND 0.024859f
C191 VOUT.t2 GND 0.008839f
C192 VOUT.t11 GND 0.008839f
C193 VOUT.n33 GND 0.041993f
C194 VOUT.n34 GND 0.699174f
C195 VOUT.n35 GND 0.006304f
C196 VOUT.n36 GND 0.016282f
C197 VOUT.t5 GND 0.016345f
C198 VOUT.n37 GND 0.015988f
C199 VOUT.n38 GND 0.00461f
C200 VOUT.n39 GND 0.00299f
C201 VOUT.n40 GND 0.038717f
C202 VOUT.n41 GND 0.024859f
C203 VOUT.t0 GND 0.008839f
C204 VOUT.t3 GND 0.008839f
C205 VOUT.n42 GND 0.041993f
C206 VOUT.n43 GND 0.681982f
C207 VOUT.n44 GND 0.611432f
C208 VOUT.n45 GND 8.72067f
C209 VOUT.t19 GND 0.163671f
C210 VOUT.t33 GND 0.015304f
C211 VOUT.t29 GND 0.015304f
C212 VOUT.n46 GND 0.126339f
C213 VOUT.n47 GND 0.621342f
C214 VOUT.t13 GND 0.163671f
C215 VOUT.t20 GND 0.015304f
C216 VOUT.t21 GND 0.015304f
C217 VOUT.n48 GND 0.126339f
C218 VOUT.n49 GND 0.59659f
C219 VOUT.n50 GND 0.334938f
C220 VOUT.t17 GND 0.163671f
C221 VOUT.t22 GND 0.015304f
C222 VOUT.t24 GND 0.015304f
C223 VOUT.n51 GND 0.126339f
C224 VOUT.n52 GND 0.59659f
C225 VOUT.n53 GND 0.225371f
C226 VOUT.t25 GND 0.163671f
C227 VOUT.t34 GND 0.015304f
C228 VOUT.t35 GND 0.015304f
C229 VOUT.n54 GND 0.126339f
C230 VOUT.n55 GND 0.59659f
C231 VOUT.n56 GND 0.373926f
C232 VOUT.n57 GND 8.08769f
C233 VOUT.t12 GND 0.015304f
C234 VOUT.t15 GND 0.015304f
C235 VOUT.n58 GND 0.134379f
C236 VOUT.t32 GND 0.159201f
C237 VOUT.n59 GND 0.642418f
C238 VOUT.t26 GND 0.015304f
C239 VOUT.t23 GND 0.015304f
C240 VOUT.n60 GND 0.134379f
C241 VOUT.t28 GND 0.159201f
C242 VOUT.n61 GND 0.619086f
C243 VOUT.n62 GND 0.284228f
C244 VOUT.t30 GND 0.015304f
C245 VOUT.t27 GND 0.015304f
C246 VOUT.n63 GND 0.134379f
C247 VOUT.t31 GND 0.159201f
C248 VOUT.n64 GND 0.619086f
C249 VOUT.n65 GND 0.199305f
C250 VOUT.t16 GND 0.015304f
C251 VOUT.t14 GND 0.015304f
C252 VOUT.n66 GND 0.134379f
C253 VOUT.t18 GND 0.159201f
C254 VOUT.n67 GND 0.619086f
C255 VOUT.n68 GND 0.34786f
C256 VOUT.n69 GND 5.68025f
C257 VOUT.n70 GND 4.73036f
C258 CS_BIAS.t28 GND 0.238609f
C259 CS_BIAS.n0 GND 0.119968f
C260 CS_BIAS.n1 GND 0.005819f
C261 CS_BIAS.n2 GND 0.011558f
C262 CS_BIAS.n3 GND 0.005819f
C263 CS_BIAS.n4 GND 0.010791f
C264 CS_BIAS.t8 GND 0.238609f
C265 CS_BIAS.n5 GND 0.119968f
C266 CS_BIAS.n6 GND 0.005819f
C267 CS_BIAS.n7 GND 0.011558f
C268 CS_BIAS.n8 GND 0.005819f
C269 CS_BIAS.n9 GND 0.010791f
C270 CS_BIAS.t10 GND 0.331048f
C271 CS_BIAS.n10 GND 0.138674f
C272 CS_BIAS.t2 GND 0.238609f
C273 CS_BIAS.n11 GND 0.118798f
C274 CS_BIAS.n12 GND 0.010791f
C275 CS_BIAS.n13 GND 0.077877f
C276 CS_BIAS.n14 GND 0.005819f
C277 CS_BIAS.n15 GND 0.005819f
C278 CS_BIAS.n16 GND 0.010791f
C279 CS_BIAS.n17 GND 0.011443f
C280 CS_BIAS.n18 GND 0.004707f
C281 CS_BIAS.n19 GND 0.005819f
C282 CS_BIAS.n20 GND 0.005819f
C283 CS_BIAS.n21 GND 0.005819f
C284 CS_BIAS.n22 GND 0.010791f
C285 CS_BIAS.n23 GND 0.010791f
C286 CS_BIAS.n24 GND 0.010578f
C287 CS_BIAS.n25 GND 0.012307f
C288 CS_BIAS.n26 GND 0.078057f
C289 CS_BIAS.t9 GND 0.064937f
C290 CS_BIAS.n27 GND 0.10283f
C291 CS_BIAS.t3 GND 0.006242f
C292 CS_BIAS.t11 GND 0.006242f
C293 CS_BIAS.n28 GND 0.052095f
C294 CS_BIAS.n29 GND 0.194122f
C295 CS_BIAS.n30 GND 0.119924f
C296 CS_BIAS.t14 GND 0.238609f
C297 CS_BIAS.t18 GND 0.331023f
C298 CS_BIAS.n31 GND 0.127051f
C299 CS_BIAS.n32 GND 0.118798f
C300 CS_BIAS.n33 GND 0.010791f
C301 CS_BIAS.n34 GND 0.005791f
C302 CS_BIAS.n35 GND 0.005819f
C303 CS_BIAS.n36 GND 0.005819f
C304 CS_BIAS.n37 GND 0.010791f
C305 CS_BIAS.n38 GND 0.011443f
C306 CS_BIAS.n39 GND 0.004707f
C307 CS_BIAS.n40 GND 0.005819f
C308 CS_BIAS.n41 GND 0.005819f
C309 CS_BIAS.n42 GND 0.005819f
C310 CS_BIAS.n43 GND 0.010791f
C311 CS_BIAS.n44 GND 0.010791f
C312 CS_BIAS.n45 GND 0.010578f
C313 CS_BIAS.n46 GND 0.012307f
C314 CS_BIAS.n47 GND 0.059904f
C315 CS_BIAS.t34 GND 0.238609f
C316 CS_BIAS.n48 GND 0.119968f
C317 CS_BIAS.n49 GND 0.005819f
C318 CS_BIAS.n50 GND 0.011558f
C319 CS_BIAS.n51 GND 0.005819f
C320 CS_BIAS.n52 GND 0.010791f
C321 CS_BIAS.t26 GND 0.331048f
C322 CS_BIAS.n53 GND 0.138674f
C323 CS_BIAS.t27 GND 0.238609f
C324 CS_BIAS.n54 GND 0.118798f
C325 CS_BIAS.n55 GND 0.010791f
C326 CS_BIAS.n56 GND 0.077877f
C327 CS_BIAS.n57 GND 0.005819f
C328 CS_BIAS.n58 GND 0.005819f
C329 CS_BIAS.n59 GND 0.010791f
C330 CS_BIAS.n60 GND 0.011443f
C331 CS_BIAS.n61 GND 0.004707f
C332 CS_BIAS.n62 GND 0.005819f
C333 CS_BIAS.n63 GND 0.005819f
C334 CS_BIAS.n64 GND 0.005819f
C335 CS_BIAS.n65 GND 0.010791f
C336 CS_BIAS.n66 GND 0.010791f
C337 CS_BIAS.n67 GND 0.010578f
C338 CS_BIAS.n68 GND 0.012307f
C339 CS_BIAS.n69 GND 0.051173f
C340 CS_BIAS.n70 GND 0.069745f
C341 CS_BIAS.t30 GND 0.238609f
C342 CS_BIAS.n71 GND 0.119968f
C343 CS_BIAS.n72 GND 0.005819f
C344 CS_BIAS.n73 GND 0.011558f
C345 CS_BIAS.n74 GND 0.005819f
C346 CS_BIAS.n75 GND 0.010791f
C347 CS_BIAS.t23 GND 0.331048f
C348 CS_BIAS.n76 GND 0.138674f
C349 CS_BIAS.t25 GND 0.238609f
C350 CS_BIAS.n77 GND 0.118798f
C351 CS_BIAS.n78 GND 0.010791f
C352 CS_BIAS.n79 GND 0.077877f
C353 CS_BIAS.n80 GND 0.005819f
C354 CS_BIAS.n81 GND 0.005819f
C355 CS_BIAS.n82 GND 0.010791f
C356 CS_BIAS.n83 GND 0.011443f
C357 CS_BIAS.n84 GND 0.004707f
C358 CS_BIAS.n85 GND 0.005819f
C359 CS_BIAS.n86 GND 0.005819f
C360 CS_BIAS.n87 GND 0.005819f
C361 CS_BIAS.n88 GND 0.010791f
C362 CS_BIAS.n89 GND 0.010791f
C363 CS_BIAS.n90 GND 0.010578f
C364 CS_BIAS.n91 GND 0.012307f
C365 CS_BIAS.n92 GND 0.051173f
C366 CS_BIAS.n93 GND 0.049804f
C367 CS_BIAS.t22 GND 0.238609f
C368 CS_BIAS.n94 GND 0.119968f
C369 CS_BIAS.n95 GND 0.005819f
C370 CS_BIAS.n96 GND 0.011558f
C371 CS_BIAS.n97 GND 0.005819f
C372 CS_BIAS.n98 GND 0.010791f
C373 CS_BIAS.t12 GND 0.331048f
C374 CS_BIAS.n99 GND 0.138674f
C375 CS_BIAS.t13 GND 0.238609f
C376 CS_BIAS.n100 GND 0.118798f
C377 CS_BIAS.n101 GND 0.010791f
C378 CS_BIAS.n102 GND 0.077877f
C379 CS_BIAS.n103 GND 0.005819f
C380 CS_BIAS.n104 GND 0.005819f
C381 CS_BIAS.n105 GND 0.010791f
C382 CS_BIAS.n106 GND 0.011443f
C383 CS_BIAS.n107 GND 0.004707f
C384 CS_BIAS.n108 GND 0.005819f
C385 CS_BIAS.n109 GND 0.005819f
C386 CS_BIAS.n110 GND 0.005819f
C387 CS_BIAS.n111 GND 0.010791f
C388 CS_BIAS.n112 GND 0.010791f
C389 CS_BIAS.n113 GND 0.010578f
C390 CS_BIAS.n114 GND 0.012307f
C391 CS_BIAS.n115 GND 0.051173f
C392 CS_BIAS.n116 GND 0.285063f
C393 CS_BIAS.t32 GND 0.238609f
C394 CS_BIAS.n117 GND 0.119968f
C395 CS_BIAS.n118 GND 0.005819f
C396 CS_BIAS.n119 GND 0.011558f
C397 CS_BIAS.n120 GND 0.005819f
C398 CS_BIAS.n121 GND 0.010791f
C399 CS_BIAS.t1 GND 0.066058f
C400 CS_BIAS.t6 GND 0.238609f
C401 CS_BIAS.n122 GND 0.119968f
C402 CS_BIAS.n123 GND 0.005819f
C403 CS_BIAS.n124 GND 0.011558f
C404 CS_BIAS.n125 GND 0.005819f
C405 CS_BIAS.n126 GND 0.010791f
C406 CS_BIAS.t0 GND 0.331048f
C407 CS_BIAS.n127 GND 0.138674f
C408 CS_BIAS.t4 GND 0.238609f
C409 CS_BIAS.n128 GND 0.118798f
C410 CS_BIAS.n129 GND 0.010791f
C411 CS_BIAS.n130 GND 0.077877f
C412 CS_BIAS.n131 GND 0.005819f
C413 CS_BIAS.n132 GND 0.005819f
C414 CS_BIAS.n133 GND 0.010791f
C415 CS_BIAS.n134 GND 0.011443f
C416 CS_BIAS.n135 GND 0.004707f
C417 CS_BIAS.n136 GND 0.005819f
C418 CS_BIAS.n137 GND 0.005819f
C419 CS_BIAS.n138 GND 0.005819f
C420 CS_BIAS.n139 GND 0.010791f
C421 CS_BIAS.n140 GND 0.010791f
C422 CS_BIAS.n141 GND 0.010578f
C423 CS_BIAS.n142 GND 0.012307f
C424 CS_BIAS.n143 GND 0.083549f
C425 CS_BIAS.t5 GND 0.006242f
C426 CS_BIAS.t7 GND 0.006242f
C427 CS_BIAS.n144 GND 0.051533f
C428 CS_BIAS.n145 GND 0.125118f
C429 CS_BIAS.n146 GND 0.165782f
C430 CS_BIAS.n147 GND 0.119923f
C431 CS_BIAS.t35 GND 0.238609f
C432 CS_BIAS.t15 GND 0.331024f
C433 CS_BIAS.n148 GND 0.12705f
C434 CS_BIAS.n149 GND 0.118798f
C435 CS_BIAS.n150 GND 0.010791f
C436 CS_BIAS.n151 GND 0.005791f
C437 CS_BIAS.n152 GND 0.005819f
C438 CS_BIAS.n153 GND 0.005819f
C439 CS_BIAS.n154 GND 0.010791f
C440 CS_BIAS.n155 GND 0.011443f
C441 CS_BIAS.n156 GND 0.004707f
C442 CS_BIAS.n157 GND 0.005819f
C443 CS_BIAS.n158 GND 0.005819f
C444 CS_BIAS.n159 GND 0.005819f
C445 CS_BIAS.n160 GND 0.010791f
C446 CS_BIAS.n161 GND 0.010791f
C447 CS_BIAS.n162 GND 0.010578f
C448 CS_BIAS.n163 GND 0.012307f
C449 CS_BIAS.n164 GND 0.059904f
C450 CS_BIAS.t24 GND 0.238609f
C451 CS_BIAS.n165 GND 0.119968f
C452 CS_BIAS.n166 GND 0.005819f
C453 CS_BIAS.n167 GND 0.011558f
C454 CS_BIAS.n168 GND 0.005819f
C455 CS_BIAS.n169 GND 0.010791f
C456 CS_BIAS.t19 GND 0.331048f
C457 CS_BIAS.n170 GND 0.138674f
C458 CS_BIAS.t21 GND 0.238609f
C459 CS_BIAS.n171 GND 0.118798f
C460 CS_BIAS.n172 GND 0.010791f
C461 CS_BIAS.n173 GND 0.077877f
C462 CS_BIAS.n174 GND 0.005819f
C463 CS_BIAS.n175 GND 0.005819f
C464 CS_BIAS.n176 GND 0.010791f
C465 CS_BIAS.n177 GND 0.011443f
C466 CS_BIAS.n178 GND 0.004707f
C467 CS_BIAS.n179 GND 0.005819f
C468 CS_BIAS.n180 GND 0.005819f
C469 CS_BIAS.n181 GND 0.005819f
C470 CS_BIAS.n182 GND 0.010791f
C471 CS_BIAS.n183 GND 0.010791f
C472 CS_BIAS.n184 GND 0.010578f
C473 CS_BIAS.n185 GND 0.012307f
C474 CS_BIAS.n186 GND 0.051173f
C475 CS_BIAS.n187 GND 0.069745f
C476 CS_BIAS.t20 GND 0.238609f
C477 CS_BIAS.n188 GND 0.119968f
C478 CS_BIAS.n189 GND 0.005819f
C479 CS_BIAS.n190 GND 0.011558f
C480 CS_BIAS.n191 GND 0.005819f
C481 CS_BIAS.n192 GND 0.010791f
C482 CS_BIAS.t16 GND 0.331048f
C483 CS_BIAS.n193 GND 0.138674f
C484 CS_BIAS.t17 GND 0.238609f
C485 CS_BIAS.n194 GND 0.118798f
C486 CS_BIAS.n195 GND 0.010791f
C487 CS_BIAS.n196 GND 0.077877f
C488 CS_BIAS.n197 GND 0.005819f
C489 CS_BIAS.n198 GND 0.005819f
C490 CS_BIAS.n199 GND 0.010791f
C491 CS_BIAS.n200 GND 0.011443f
C492 CS_BIAS.n201 GND 0.004707f
C493 CS_BIAS.n202 GND 0.005819f
C494 CS_BIAS.n203 GND 0.005819f
C495 CS_BIAS.n204 GND 0.005819f
C496 CS_BIAS.n205 GND 0.010791f
C497 CS_BIAS.n206 GND 0.010791f
C498 CS_BIAS.n207 GND 0.010578f
C499 CS_BIAS.n208 GND 0.012307f
C500 CS_BIAS.n209 GND 0.051173f
C501 CS_BIAS.n210 GND 0.049804f
C502 CS_BIAS.t33 GND 0.238609f
C503 CS_BIAS.n211 GND 0.119968f
C504 CS_BIAS.n212 GND 0.005819f
C505 CS_BIAS.n213 GND 0.011558f
C506 CS_BIAS.n214 GND 0.005819f
C507 CS_BIAS.n215 GND 0.010791f
C508 CS_BIAS.t29 GND 0.331048f
C509 CS_BIAS.n216 GND 0.138674f
C510 CS_BIAS.t31 GND 0.238609f
C511 CS_BIAS.n217 GND 0.118798f
C512 CS_BIAS.n218 GND 0.010791f
C513 CS_BIAS.n219 GND 0.077877f
C514 CS_BIAS.n220 GND 0.005819f
C515 CS_BIAS.n221 GND 0.005819f
C516 CS_BIAS.n222 GND 0.010791f
C517 CS_BIAS.n223 GND 0.011443f
C518 CS_BIAS.n224 GND 0.004707f
C519 CS_BIAS.n225 GND 0.005819f
C520 CS_BIAS.n226 GND 0.005819f
C521 CS_BIAS.n227 GND 0.005819f
C522 CS_BIAS.n228 GND 0.010791f
C523 CS_BIAS.n229 GND 0.010791f
C524 CS_BIAS.n230 GND 0.010578f
C525 CS_BIAS.n231 GND 0.012307f
C526 CS_BIAS.n232 GND 0.051173f
C527 CS_BIAS.n233 GND 0.099978f
C528 CS_BIAS.n234 GND 3.32642f
C529 a_n1672_n179.n0 GND 2.81788f
C530 a_n1672_n179.n1 GND 0.351236f
C531 a_n1672_n179.n2 GND 0.016932f
C532 a_n1672_n179.n3 GND 0.351236f
C533 a_n1672_n179.n4 GND 0.016932f
C534 a_n1672_n179.n5 GND 0.016932f
C535 a_n1672_n179.n6 GND 0.016932f
C536 a_n1672_n179.n7 GND 0.019355f
C537 a_n1672_n179.n8 GND 0.019355f
C538 a_n1672_n179.n9 GND 0.351236f
C539 a_n1672_n179.n10 GND 0.019355f
C540 a_n1672_n179.n11 GND 0.019439f
C541 a_n1672_n179.n12 GND 0.016932f
C542 a_n1672_n179.n13 GND 0.019439f
C543 a_n1672_n179.n14 GND 0.016932f
C544 a_n1672_n179.n15 GND 1.92784f
C545 a_n1672_n179.n16 GND 1.89762f
C546 a_n1672_n179.n17 GND 0.014889f
C547 a_n1672_n179.n18 GND 0.043178f
C548 a_n1672_n179.n19 GND 0.008708f
C549 a_n1672_n179.n20 GND 0.022132f
C550 a_n1672_n179.t9 GND 0.033312f
C551 a_n1672_n179.n21 GND 0.014889f
C552 a_n1672_n179.n22 GND 0.019439f
C553 a_n1672_n179.n23 GND 0.043178f
C554 a_n1672_n179.n24 GND 0.008708f
C555 a_n1672_n179.n25 GND 0.008224f
C556 a_n1672_n179.n26 GND 0.127465f
C557 a_n1672_n179.t4 GND 0.474871f
C558 a_n1672_n179.t3 GND 0.04995f
C559 a_n1672_n179.t7 GND 0.04995f
C560 a_n1672_n179.n27 GND 0.372881f
C561 a_n1672_n179.t0 GND 0.474872f
C562 a_n1672_n179.t1 GND 0.04995f
C563 a_n1672_n179.t13 GND 0.04995f
C564 a_n1672_n179.n28 GND 0.372881f
C565 a_n1672_n179.n29 GND 1.04976f
C566 a_n1672_n179.n30 GND 0.022132f
C567 a_n1672_n179.t8 GND 0.033312f
C568 a_n1672_n179.n31 GND 0.014889f
C569 a_n1672_n179.n32 GND 0.019439f
C570 a_n1672_n179.n33 GND 0.043178f
C571 a_n1672_n179.n34 GND 0.008708f
C572 a_n1672_n179.n35 GND 0.008224f
C573 a_n1672_n179.n36 GND 0.127486f
C574 a_n1672_n179.t14 GND 0.04995f
C575 a_n1672_n179.t11 GND 0.04995f
C576 a_n1672_n179.n37 GND 0.372879f
C577 a_n1672_n179.t5 GND 0.474871f
C578 a_n1672_n179.t6 GND 0.04995f
C579 a_n1672_n179.t2 GND 0.04995f
C580 a_n1672_n179.n38 GND 0.372879f
C581 a_n1672_n179.t12 GND 0.474871f
C582 a_n1672_n179.n39 GND 0.73144f
C583 a_n1672_n179.n40 GND 0.89511f
C584 a_n1672_n179.n41 GND 1.586f
C585 a_n1672_n179.n42 GND 0.127465f
C586 a_n1672_n179.n43 GND 0.022132f
C587 a_n1672_n179.n44 GND 0.008224f
C588 a_n1672_n179.n45 GND 0.019439f
C589 a_n1672_n179.n46 GND 0.019439f
C590 a_n1672_n179.t10 GND 0.033312f
C591 VDD.t90 GND 0.009941f
C592 VDD.t84 GND 0.009941f
C593 VDD.n0 GND 0.066737f
C594 VDD.t114 GND 0.009941f
C595 VDD.t108 GND 0.009941f
C596 VDD.n1 GND 0.065483f
C597 VDD.n2 GND 0.276336f
C598 VDD.t97 GND 0.009941f
C599 VDD.t92 GND 0.009941f
C600 VDD.n3 GND 0.065483f
C601 VDD.n4 GND 0.143472f
C602 VDD.t79 GND 0.009941f
C603 VDD.t110 GND 0.009941f
C604 VDD.n5 GND 0.065483f
C605 VDD.n6 GND 0.122827f
C606 VDD.t99 GND 0.009941f
C607 VDD.t106 GND 0.009941f
C608 VDD.n7 GND 0.066737f
C609 VDD.t95 GND 0.009941f
C610 VDD.t104 GND 0.009941f
C611 VDD.n8 GND 0.065483f
C612 VDD.n9 GND 0.276336f
C613 VDD.t87 GND 0.009941f
C614 VDD.t82 GND 0.009941f
C615 VDD.n10 GND 0.065483f
C616 VDD.n11 GND 0.143472f
C617 VDD.t101 GND 0.009941f
C618 VDD.t76 GND 0.009941f
C619 VDD.n12 GND 0.065483f
C620 VDD.n13 GND 0.122827f
C621 VDD.n14 GND 0.088064f
C622 VDD.n15 GND 1.7538f
C623 VDD.t68 GND 0.004713f
C624 VDD.t61 GND 0.004713f
C625 VDD.n16 GND 0.020974f
C626 VDD.n17 GND 0.003361f
C627 VDD.n18 GND 0.008681f
C628 VDD.t74 GND 0.008714f
C629 VDD.n19 GND 0.008524f
C630 VDD.n20 GND 0.002458f
C631 VDD.n21 GND 0.001594f
C632 VDD.n22 GND 0.020642f
C633 VDD.n23 GND 0.005467f
C634 VDD.n24 GND 0.36775f
C635 VDD.t67 GND 0.004713f
C636 VDD.t58 GND 0.004713f
C637 VDD.n25 GND 0.020974f
C638 VDD.n26 GND 0.003361f
C639 VDD.n27 GND 0.008681f
C640 VDD.t63 GND 0.008714f
C641 VDD.n28 GND 0.008524f
C642 VDD.n29 GND 0.002458f
C643 VDD.n30 GND 0.001594f
C644 VDD.n31 GND 0.020642f
C645 VDD.n32 GND 0.005467f
C646 VDD.n33 GND 0.359722f
C647 VDD.n34 GND 0.276087f
C648 VDD.n35 GND 0.004478f
C649 VDD.n36 GND 0.005826f
C650 VDD.n37 GND 0.004689f
C651 VDD.n38 GND 0.004689f
C652 VDD.n39 GND 0.005826f
C653 VDD.n40 GND 0.005826f
C654 VDD.t57 GND 0.196239f
C655 VDD.n41 GND 0.005826f
C656 VDD.n42 GND 0.005826f
C657 VDD.n43 GND 0.005826f
C658 VDD.n44 GND 0.392477f
C659 VDD.n45 GND 0.005826f
C660 VDD.n46 GND 0.005826f
C661 VDD.n47 GND 0.005826f
C662 VDD.n48 GND 0.005826f
C663 VDD.n49 GND 0.004689f
C664 VDD.n50 GND 0.005826f
C665 VDD.n51 GND 0.005826f
C666 VDD.n52 GND 0.005826f
C667 VDD.n53 GND 0.005826f
C668 VDD.n54 GND 0.392477f
C669 VDD.n55 GND 0.005826f
C670 VDD.n56 GND 0.005826f
C671 VDD.n57 GND 0.005826f
C672 VDD.n58 GND 0.005826f
C673 VDD.n59 GND 0.005826f
C674 VDD.n60 GND 0.004689f
C675 VDD.n61 GND 0.005826f
C676 VDD.n62 GND 0.005826f
C677 VDD.n63 GND 0.005826f
C678 VDD.n64 GND 0.005826f
C679 VDD.n65 GND 0.372853f
C680 VDD.n66 GND 0.005826f
C681 VDD.n67 GND 0.005826f
C682 VDD.n68 GND 0.005826f
C683 VDD.n69 GND 0.005826f
C684 VDD.n70 GND 0.005826f
C685 VDD.n71 GND 0.004689f
C686 VDD.n72 GND 0.005826f
C687 VDD.t62 GND 0.196239f
C688 VDD.n73 GND 0.005826f
C689 VDD.n74 GND 0.005826f
C690 VDD.n75 GND 0.005826f
C691 VDD.n76 GND 0.392477f
C692 VDD.n77 GND 0.005826f
C693 VDD.n78 GND 0.005826f
C694 VDD.n79 GND 0.005826f
C695 VDD.n80 GND 0.005826f
C696 VDD.n81 GND 0.005826f
C697 VDD.n82 GND 0.004689f
C698 VDD.n83 GND 0.005826f
C699 VDD.n84 GND 0.005826f
C700 VDD.n85 GND 0.005826f
C701 VDD.n86 GND 0.005826f
C702 VDD.n87 GND 0.392477f
C703 VDD.n88 GND 0.005826f
C704 VDD.n89 GND 0.005826f
C705 VDD.n90 GND 0.005826f
C706 VDD.n91 GND 0.005826f
C707 VDD.n92 GND 0.005826f
C708 VDD.n93 GND 0.004689f
C709 VDD.n94 GND 0.005826f
C710 VDD.n95 GND 0.005826f
C711 VDD.n96 GND 0.005826f
C712 VDD.n97 GND 0.005826f
C713 VDD.n98 GND 0.392477f
C714 VDD.n99 GND 0.005826f
C715 VDD.n100 GND 0.005826f
C716 VDD.n101 GND 0.005826f
C717 VDD.n102 GND 0.005826f
C718 VDD.n103 GND 0.005826f
C719 VDD.n104 GND 0.004689f
C720 VDD.n105 GND 0.005826f
C721 VDD.n106 GND 0.005826f
C722 VDD.n107 GND 0.005826f
C723 VDD.n108 GND 0.005826f
C724 VDD.t5 GND 0.196239f
C725 VDD.n109 GND 0.005826f
C726 VDD.n110 GND 0.005826f
C727 VDD.n111 GND 0.005826f
C728 VDD.n112 GND 0.005826f
C729 VDD.n113 GND 0.005826f
C730 VDD.n114 GND 0.004689f
C731 VDD.n115 GND 0.005826f
C732 VDD.n116 GND 0.298283f
C733 VDD.n117 GND 0.005826f
C734 VDD.n118 GND 0.005826f
C735 VDD.n119 GND 0.005826f
C736 VDD.n120 GND 0.392477f
C737 VDD.n121 GND 0.005826f
C738 VDD.n122 GND 0.005826f
C739 VDD.n123 GND 0.005826f
C740 VDD.n124 GND 0.005826f
C741 VDD.n125 GND 0.005826f
C742 VDD.n126 GND 0.003892f
C743 VDD.n127 GND 0.012127f
C744 VDD.n128 GND 0.005826f
C745 VDD.n129 GND 0.012127f
C746 VDD.n139 GND 0.005826f
C747 VDD.n140 GND 0.012127f
C748 VDD.n141 GND 0.012459f
C749 VDD.n142 GND 0.004689f
C750 VDD.n143 GND 0.005826f
C751 VDD.n144 GND 0.005826f
C752 VDD.n145 GND 0.005826f
C753 VDD.n146 GND 0.005826f
C754 VDD.n147 GND 0.005826f
C755 VDD.n148 GND 0.005826f
C756 VDD.n149 GND 0.005826f
C757 VDD.n150 GND 0.005826f
C758 VDD.n151 GND 0.005826f
C759 VDD.n152 GND 0.005826f
C760 VDD.n153 GND 0.005826f
C761 VDD.n154 GND 0.005826f
C762 VDD.n155 GND 0.005826f
C763 VDD.n156 GND 0.012459f
C764 VDD.n157 GND 0.002978f
C765 VDD.t7 GND 0.019391f
C766 VDD.t6 GND 0.032488f
C767 VDD.t4 GND 0.334077f
C768 VDD.n158 GND 0.060478f
C769 VDD.n159 GND 0.043121f
C770 VDD.n160 GND 0.005826f
C771 VDD.n161 GND 0.004689f
C772 VDD.n162 GND 0.005826f
C773 VDD.n163 GND 0.004689f
C774 VDD.n164 GND 0.005826f
C775 VDD.n165 GND 0.004689f
C776 VDD.n166 GND 0.005826f
C777 VDD.n167 GND 0.004689f
C778 VDD.n168 GND 0.005826f
C779 VDD.n169 GND 0.004689f
C780 VDD.n170 GND 0.005826f
C781 VDD.n171 GND 0.004689f
C782 VDD.n172 GND 0.005826f
C783 VDD.n173 GND 0.004689f
C784 VDD.n174 GND 0.005826f
C785 VDD.n175 GND 0.004689f
C786 VDD.n176 GND 0.005826f
C787 VDD.n177 GND 0.004689f
C788 VDD.n178 GND 0.005826f
C789 VDD.n179 GND 0.005826f
C790 VDD.n180 GND 0.392477f
C791 VDD.n181 GND 0.005826f
C792 VDD.n182 GND 0.004689f
C793 VDD.n183 GND 0.005826f
C794 VDD.n184 GND 0.004689f
C795 VDD.n185 GND 0.005826f
C796 VDD.n186 GND 0.392477f
C797 VDD.n187 GND 0.005826f
C798 VDD.n188 GND 0.005826f
C799 VDD.n189 GND 0.004689f
C800 VDD.n190 GND 0.005826f
C801 VDD.n191 GND 0.004689f
C802 VDD.n192 GND 0.005826f
C803 VDD.n193 GND 0.392477f
C804 VDD.n194 GND 0.005826f
C805 VDD.n195 GND 0.004689f
C806 VDD.n196 GND 0.005826f
C807 VDD.n197 GND 0.004689f
C808 VDD.n198 GND 0.005826f
C809 VDD.n199 GND 0.392477f
C810 VDD.n200 GND 0.005826f
C811 VDD.n201 GND 0.004689f
C812 VDD.n202 GND 0.005826f
C813 VDD.n203 GND 0.004689f
C814 VDD.n204 GND 0.005826f
C815 VDD.n205 GND 0.392477f
C816 VDD.n206 GND 0.005826f
C817 VDD.n207 GND 0.004689f
C818 VDD.n208 GND 0.005826f
C819 VDD.n209 GND 0.004689f
C820 VDD.n210 GND 0.005826f
C821 VDD.t66 GND 0.196239f
C822 VDD.n211 GND 0.005826f
C823 VDD.n212 GND 0.004689f
C824 VDD.n213 GND 0.005826f
C825 VDD.n214 GND 0.004689f
C826 VDD.n215 GND 0.005826f
C827 VDD.n216 GND 0.392477f
C828 VDD.n217 GND 0.215862f
C829 VDD.n218 GND 0.005826f
C830 VDD.n219 GND 0.004689f
C831 VDD.n220 GND 0.005826f
C832 VDD.n221 GND 0.004689f
C833 VDD.n222 GND 0.005826f
C834 VDD.n223 GND 0.392477f
C835 VDD.n224 GND 0.005826f
C836 VDD.n225 GND 0.004689f
C837 VDD.n226 GND 0.005826f
C838 VDD.n227 GND 0.004689f
C839 VDD.n228 GND 0.005826f
C840 VDD.n229 GND 0.392477f
C841 VDD.n230 GND 0.005826f
C842 VDD.n231 GND 0.004689f
C843 VDD.n232 GND 0.005826f
C844 VDD.n233 GND 0.004689f
C845 VDD.n234 GND 0.005826f
C846 VDD.n235 GND 0.392477f
C847 VDD.n236 GND 0.005826f
C848 VDD.n237 GND 0.004689f
C849 VDD.n238 GND 0.005826f
C850 VDD.n239 GND 0.004689f
C851 VDD.n240 GND 0.005826f
C852 VDD.n241 GND 0.392477f
C853 VDD.n242 GND 0.005826f
C854 VDD.n243 GND 0.004689f
C855 VDD.n244 GND 0.005826f
C856 VDD.n245 GND 0.004689f
C857 VDD.n246 GND 0.005826f
C858 VDD.n247 GND 0.392477f
C859 VDD.n248 GND 0.005826f
C860 VDD.n249 GND 0.004689f
C861 VDD.n250 GND 0.005826f
C862 VDD.n251 GND 0.004689f
C863 VDD.n252 GND 0.005826f
C864 VDD.n253 GND 0.290433f
C865 VDD.n254 GND 0.005826f
C866 VDD.n255 GND 0.004689f
C867 VDD.n256 GND 0.005826f
C868 VDD.n257 GND 0.004689f
C869 VDD.n258 GND 0.005826f
C870 VDD.n259 GND 0.392477f
C871 VDD.n260 GND 0.005826f
C872 VDD.n261 GND 0.004689f
C873 VDD.n262 GND 0.005826f
C874 VDD.n263 GND 0.004689f
C875 VDD.n264 GND 0.005826f
C876 VDD.n265 GND 0.392477f
C877 VDD.n266 GND 0.005826f
C878 VDD.n267 GND 0.004689f
C879 VDD.n268 GND 0.005826f
C880 VDD.n269 GND 0.004689f
C881 VDD.n270 GND 0.005826f
C882 VDD.n271 GND 0.392477f
C883 VDD.n272 GND 0.005826f
C884 VDD.n273 GND 0.004689f
C885 VDD.n274 GND 0.012459f
C886 VDD.n275 GND 0.012459f
C887 VDD.n276 GND 0.396402f
C888 VDD.n277 GND 0.009601f
C889 VDD.n298 GND 0.008926f
C890 VDD.n299 GND 0.003962f
C891 VDD.n300 GND 0.008926f
C892 VDD.t26 GND 0.064081f
C893 VDD.t25 GND 0.074164f
C894 VDD.t23 GND 0.279207f
C895 VDD.n301 GND 0.052604f
C896 VDD.n302 GND 0.035175f
C897 VDD.n303 GND 0.009395f
C898 VDD.n304 GND 0.003962f
C899 VDD.n305 GND 0.003962f
C900 VDD.n306 GND 0.188389f
C901 VDD.n307 GND 0.003962f
C902 VDD.n308 GND 0.003962f
C903 VDD.n309 GND 0.003962f
C904 VDD.n310 GND 0.003962f
C905 VDD.n311 GND 0.003962f
C906 VDD.n312 GND 0.266884f
C907 VDD.n313 GND 0.003962f
C908 VDD.n314 GND 0.003962f
C909 VDD.t98 GND 0.133442f
C910 VDD.n315 GND 0.003962f
C911 VDD.n316 GND 0.003962f
C912 VDD.n317 GND 0.003962f
C913 VDD.t29 GND 0.064081f
C914 VDD.t28 GND 0.074164f
C915 VDD.t27 GND 0.279207f
C916 VDD.n318 GND 0.052604f
C917 VDD.n319 GND 0.035175f
C918 VDD.n320 GND 0.003962f
C919 VDD.n321 GND 0.003962f
C920 VDD.n322 GND 0.266884f
C921 VDD.n323 GND 0.003962f
C922 VDD.n324 GND 0.003962f
C923 VDD.n325 GND 0.003962f
C924 VDD.n326 GND 0.003962f
C925 VDD.n327 GND 0.003962f
C926 VDD.n328 GND 0.266884f
C927 VDD.n329 GND 0.003962f
C928 VDD.n330 GND 0.003962f
C929 VDD.n331 GND 0.003962f
C930 VDD.n332 GND 0.003962f
C931 VDD.n333 GND 0.003962f
C932 VDD.n334 GND 0.003962f
C933 VDD.n335 GND 0.204088f
C934 VDD.n336 GND 0.003962f
C935 VDD.n337 GND 0.003962f
C936 VDD.n338 GND 0.003962f
C937 VDD.n339 GND 0.003962f
C938 VDD.n340 GND 0.003962f
C939 VDD.n341 GND 0.266884f
C940 VDD.n342 GND 0.003962f
C941 VDD.n343 GND 0.003962f
C942 VDD.t103 GND 0.133442f
C943 VDD.n344 GND 0.003962f
C944 VDD.n345 GND 0.003962f
C945 VDD.n346 GND 0.003962f
C946 VDD.n347 GND 0.266884f
C947 VDD.n348 GND 0.003962f
C948 VDD.n349 GND 0.003962f
C949 VDD.n350 GND 0.003962f
C950 VDD.n351 GND 0.003962f
C951 VDD.n352 GND 0.003962f
C952 VDD.n353 GND 0.176615f
C953 VDD.n354 GND 0.003962f
C954 VDD.n355 GND 0.003962f
C955 VDD.n356 GND 0.003962f
C956 VDD.n357 GND 0.003962f
C957 VDD.n358 GND 0.003962f
C958 VDD.n359 GND 0.219787f
C959 VDD.n360 GND 0.003962f
C960 VDD.n361 GND 0.003962f
C961 VDD.t77 GND 0.133442f
C962 VDD.n362 GND 0.003962f
C963 VDD.n363 GND 0.003962f
C964 VDD.n364 GND 0.003962f
C965 VDD.n365 GND 0.266884f
C966 VDD.n366 GND 0.003962f
C967 VDD.n367 GND 0.003962f
C968 VDD.t94 GND 0.133442f
C969 VDD.n368 GND 0.003962f
C970 VDD.n369 GND 0.003962f
C971 VDD.n370 GND 0.003962f
C972 VDD.n371 GND 0.266884f
C973 VDD.n372 GND 0.003962f
C974 VDD.n373 GND 0.003962f
C975 VDD.n374 GND 0.003962f
C976 VDD.n375 GND 0.003962f
C977 VDD.n376 GND 0.003962f
C978 VDD.n377 GND 0.192314f
C979 VDD.n378 GND 0.003962f
C980 VDD.n379 GND 0.003962f
C981 VDD.n380 GND 0.003962f
C982 VDD.n381 GND 0.003962f
C983 VDD.n382 GND 0.003962f
C984 VDD.n383 GND 0.266884f
C985 VDD.n384 GND 0.003962f
C986 VDD.n385 GND 0.003962f
C987 VDD.t111 GND 0.133442f
C988 VDD.n386 GND 0.003962f
C989 VDD.n387 GND 0.003962f
C990 VDD.n388 GND 0.003962f
C991 VDD.n389 GND 0.266884f
C992 VDD.n390 GND 0.003962f
C993 VDD.n391 GND 0.003962f
C994 VDD.n392 GND 0.003962f
C995 VDD.n393 GND 0.003962f
C996 VDD.n394 GND 0.003962f
C997 VDD.n395 GND 0.260997f
C998 VDD.n396 GND 0.003962f
C999 VDD.n397 GND 0.003962f
C1000 VDD.n398 GND 0.003962f
C1001 VDD.n399 GND 0.003962f
C1002 VDD.n400 GND 0.003962f
C1003 VDD.n401 GND 0.208013f
C1004 VDD.n402 GND 0.003962f
C1005 VDD.n403 GND 0.003962f
C1006 VDD.t81 GND 0.133442f
C1007 VDD.n404 GND 0.003962f
C1008 VDD.n405 GND 0.003962f
C1009 VDD.n406 GND 0.003962f
C1010 VDD.n407 GND 0.266884f
C1011 VDD.n408 GND 0.003962f
C1012 VDD.n409 GND 0.003962f
C1013 VDD.t102 GND 0.133442f
C1014 VDD.n410 GND 0.003962f
C1015 VDD.n411 GND 0.003962f
C1016 VDD.n412 GND 0.003962f
C1017 VDD.n413 GND 0.266884f
C1018 VDD.n414 GND 0.003962f
C1019 VDD.n415 GND 0.003962f
C1020 VDD.n416 GND 0.003962f
C1021 VDD.n417 GND 0.003962f
C1022 VDD.n418 GND 0.003962f
C1023 VDD.n419 GND 0.266884f
C1024 VDD.n420 GND 0.003962f
C1025 VDD.n421 GND 0.003962f
C1026 VDD.n422 GND 0.003962f
C1027 VDD.n423 GND 0.003962f
C1028 VDD.n424 GND 0.003962f
C1029 VDD.t86 GND 0.133442f
C1030 VDD.n425 GND 0.003962f
C1031 VDD.n426 GND 0.003962f
C1032 VDD.n427 GND 0.003962f
C1033 VDD.n428 GND 0.003962f
C1034 VDD.n429 GND 0.003962f
C1035 VDD.n430 GND 0.266884f
C1036 VDD.n431 GND 0.003962f
C1037 VDD.n432 GND 0.003962f
C1038 VDD.t88 GND 0.133442f
C1039 VDD.n433 GND 0.003962f
C1040 VDD.n434 GND 0.003962f
C1041 VDD.n435 GND 0.003962f
C1042 VDD.n436 GND 0.266884f
C1043 VDD.n437 GND 0.003962f
C1044 VDD.n438 GND 0.003962f
C1045 VDD.n439 GND 0.003962f
C1046 VDD.n440 GND 0.003962f
C1047 VDD.n441 GND 0.003962f
C1048 VDD.n442 GND 0.266884f
C1049 VDD.n443 GND 0.003962f
C1050 VDD.n444 GND 0.003962f
C1051 VDD.n445 GND 0.003962f
C1052 VDD.n446 GND 0.003962f
C1053 VDD.n447 GND 0.003962f
C1054 VDD.t75 GND 0.133442f
C1055 VDD.n448 GND 0.003962f
C1056 VDD.n449 GND 0.003962f
C1057 VDD.n450 GND 0.003962f
C1058 VDD.n451 GND 0.003962f
C1059 VDD.n452 GND 0.003962f
C1060 VDD.n453 GND 0.266884f
C1061 VDD.n454 GND 0.003962f
C1062 VDD.n455 GND 0.003962f
C1063 VDD.n456 GND 0.241373f
C1064 VDD.n457 GND 0.003962f
C1065 VDD.n458 GND 0.003962f
C1066 VDD.n459 GND 0.003962f
C1067 VDD.t16 GND 0.266884f
C1068 VDD.n460 GND 0.003962f
C1069 VDD.n461 GND 0.003962f
C1070 VDD.n462 GND 0.003962f
C1071 VDD.n463 GND 0.003962f
C1072 VDD.n464 GND 0.003962f
C1073 VDD.n465 GND 0.266884f
C1074 VDD.n466 GND 0.003962f
C1075 VDD.n467 GND 0.003962f
C1076 VDD.n468 GND 0.003962f
C1077 VDD.n469 GND 0.003962f
C1078 VDD.n470 GND 0.003962f
C1079 VDD.t100 GND 0.133442f
C1080 VDD.n471 GND 0.003962f
C1081 VDD.n472 GND 0.003962f
C1082 VDD.n473 GND 0.003962f
C1083 VDD.n474 GND 0.009601f
C1084 VDD.n475 GND 0.009601f
C1085 VDD.n476 GND 0.396402f
C1086 VDD.n477 GND 0.009601f
C1087 VDD.n498 GND 0.008926f
C1088 VDD.n499 GND 0.003962f
C1089 VDD.n500 GND 0.008926f
C1090 VDD.t45 GND 0.064081f
C1091 VDD.t44 GND 0.074164f
C1092 VDD.t43 GND 0.279207f
C1093 VDD.n501 GND 0.052604f
C1094 VDD.n502 GND 0.035175f
C1095 VDD.n503 GND 0.009395f
C1096 VDD.n504 GND 0.003962f
C1097 VDD.n505 GND 0.003962f
C1098 VDD.t109 GND 0.133442f
C1099 VDD.n506 GND 0.003962f
C1100 VDD.n507 GND 0.003962f
C1101 VDD.n508 GND 0.003962f
C1102 VDD.n509 GND 0.003962f
C1103 VDD.n510 GND 0.003962f
C1104 VDD.n511 GND 0.266884f
C1105 VDD.n512 GND 0.003962f
C1106 VDD.n513 GND 0.003962f
C1107 VDD.n514 GND 0.174652f
C1108 VDD.n515 GND 0.003962f
C1109 VDD.n516 GND 0.003962f
C1110 VDD.n517 GND 0.003962f
C1111 VDD.t42 GND 0.064081f
C1112 VDD.t41 GND 0.074164f
C1113 VDD.t39 GND 0.279207f
C1114 VDD.n518 GND 0.052604f
C1115 VDD.n519 GND 0.035175f
C1116 VDD.n520 GND 0.003962f
C1117 VDD.n521 GND 0.003962f
C1118 VDD.n522 GND 0.266884f
C1119 VDD.n523 GND 0.003962f
C1120 VDD.n524 GND 0.003962f
C1121 VDD.n525 GND 0.003962f
C1122 VDD.n526 GND 0.003962f
C1123 VDD.n527 GND 0.003962f
C1124 VDD.n528 GND 0.266884f
C1125 VDD.n529 GND 0.003962f
C1126 VDD.n530 GND 0.003962f
C1127 VDD.n531 GND 0.003962f
C1128 VDD.n532 GND 0.003962f
C1129 VDD.n533 GND 0.003962f
C1130 VDD.n534 GND 0.003962f
C1131 VDD.t78 GND 0.133442f
C1132 VDD.n535 GND 0.003962f
C1133 VDD.n536 GND 0.003962f
C1134 VDD.n537 GND 0.003962f
C1135 VDD.n538 GND 0.003962f
C1136 VDD.n539 GND 0.003962f
C1137 VDD.n540 GND 0.266884f
C1138 VDD.n541 GND 0.003962f
C1139 VDD.n542 GND 0.003962f
C1140 VDD.n543 GND 0.158953f
C1141 VDD.n544 GND 0.003962f
C1142 VDD.n545 GND 0.003962f
C1143 VDD.n546 GND 0.003962f
C1144 VDD.n547 GND 0.266884f
C1145 VDD.n548 GND 0.003962f
C1146 VDD.n549 GND 0.003962f
C1147 VDD.n550 GND 0.003962f
C1148 VDD.n551 GND 0.003962f
C1149 VDD.n552 GND 0.003962f
C1150 VDD.n553 GND 0.176615f
C1151 VDD.n554 GND 0.003962f
C1152 VDD.n555 GND 0.003962f
C1153 VDD.n556 GND 0.003962f
C1154 VDD.n557 GND 0.003962f
C1155 VDD.n558 GND 0.003962f
C1156 VDD.t91 GND 0.133442f
C1157 VDD.n559 GND 0.003962f
C1158 VDD.n560 GND 0.003962f
C1159 VDD.t112 GND 0.133442f
C1160 VDD.n561 GND 0.003962f
C1161 VDD.n562 GND 0.003962f
C1162 VDD.n563 GND 0.003962f
C1163 VDD.n564 GND 0.266884f
C1164 VDD.n565 GND 0.003962f
C1165 VDD.n566 GND 0.003962f
C1166 VDD.n567 GND 0.143254f
C1167 VDD.n568 GND 0.003962f
C1168 VDD.n569 GND 0.003962f
C1169 VDD.n570 GND 0.003962f
C1170 VDD.n571 GND 0.266884f
C1171 VDD.n572 GND 0.003962f
C1172 VDD.n573 GND 0.003962f
C1173 VDD.n574 GND 0.003962f
C1174 VDD.n575 GND 0.003962f
C1175 VDD.n576 GND 0.003962f
C1176 VDD.n577 GND 0.192314f
C1177 VDD.n578 GND 0.003962f
C1178 VDD.n579 GND 0.003962f
C1179 VDD.n580 GND 0.003962f
C1180 VDD.n581 GND 0.003962f
C1181 VDD.n582 GND 0.003962f
C1182 VDD.n583 GND 0.139329f
C1183 VDD.n584 GND 0.003962f
C1184 VDD.n585 GND 0.003962f
C1185 VDD.t93 GND 0.133442f
C1186 VDD.n586 GND 0.003962f
C1187 VDD.n587 GND 0.003962f
C1188 VDD.n588 GND 0.003962f
C1189 VDD.n589 GND 0.266884f
C1190 VDD.n590 GND 0.003962f
C1191 VDD.n591 GND 0.003962f
C1192 VDD.t96 GND 0.133442f
C1193 VDD.n592 GND 0.003962f
C1194 VDD.n593 GND 0.003962f
C1195 VDD.n594 GND 0.003962f
C1196 VDD.n595 GND 0.266884f
C1197 VDD.n596 GND 0.003962f
C1198 VDD.n597 GND 0.003962f
C1199 VDD.n598 GND 0.003962f
C1200 VDD.n599 GND 0.003962f
C1201 VDD.n600 GND 0.003962f
C1202 VDD.n601 GND 0.208013f
C1203 VDD.n602 GND 0.003962f
C1204 VDD.n603 GND 0.003962f
C1205 VDD.n604 GND 0.003962f
C1206 VDD.n605 GND 0.003962f
C1207 VDD.n606 GND 0.003962f
C1208 VDD.n607 GND 0.266884f
C1209 VDD.n608 GND 0.003962f
C1210 VDD.n609 GND 0.003962f
C1211 VDD.t85 GND 0.133442f
C1212 VDD.n610 GND 0.003962f
C1213 VDD.n611 GND 0.003962f
C1214 VDD.n612 GND 0.003962f
C1215 VDD.n613 GND 0.266884f
C1216 VDD.n614 GND 0.003962f
C1217 VDD.n615 GND 0.003962f
C1218 VDD.n616 GND 0.003962f
C1219 VDD.n617 GND 0.003962f
C1220 VDD.n618 GND 0.003962f
C1221 VDD.n619 GND 0.180539f
C1222 VDD.n620 GND 0.003962f
C1223 VDD.n621 GND 0.003962f
C1224 VDD.n622 GND 0.003962f
C1225 VDD.n623 GND 0.003962f
C1226 VDD.n624 GND 0.003962f
C1227 VDD.n625 GND 0.223712f
C1228 VDD.n626 GND 0.003962f
C1229 VDD.n627 GND 0.003962f
C1230 VDD.t107 GND 0.133442f
C1231 VDD.n628 GND 0.003962f
C1232 VDD.n629 GND 0.003962f
C1233 VDD.n630 GND 0.003962f
C1234 VDD.n631 GND 0.266884f
C1235 VDD.n632 GND 0.003962f
C1236 VDD.n633 GND 0.003962f
C1237 VDD.t80 GND 0.133442f
C1238 VDD.n634 GND 0.003962f
C1239 VDD.n635 GND 0.003962f
C1240 VDD.n636 GND 0.003962f
C1241 VDD.n637 GND 0.266884f
C1242 VDD.n638 GND 0.003962f
C1243 VDD.n639 GND 0.003962f
C1244 VDD.n640 GND 0.003962f
C1245 VDD.n641 GND 0.003962f
C1246 VDD.n642 GND 0.003962f
C1247 VDD.n643 GND 0.196239f
C1248 VDD.n644 GND 0.003962f
C1249 VDD.n645 GND 0.003962f
C1250 VDD.n646 GND 0.003962f
C1251 VDD.n647 GND 0.003962f
C1252 VDD.n648 GND 0.003962f
C1253 VDD.n649 GND 0.266884f
C1254 VDD.n650 GND 0.003962f
C1255 VDD.n651 GND 0.003962f
C1256 VDD.t113 GND 0.133442f
C1257 VDD.n652 GND 0.003962f
C1258 VDD.n653 GND 0.003962f
C1259 VDD.n654 GND 0.003962f
C1260 VDD.n655 GND 0.266884f
C1261 VDD.n656 GND 0.003962f
C1262 VDD.n657 GND 0.003962f
C1263 VDD.n658 GND 0.003962f
C1264 VDD.n659 GND 0.003962f
C1265 VDD.n660 GND 0.003962f
C1266 VDD.t50 GND 0.266884f
C1267 VDD.n661 GND 0.003962f
C1268 VDD.n662 GND 0.003962f
C1269 VDD.n663 GND 0.003962f
C1270 VDD.n664 GND 0.003962f
C1271 VDD.n665 GND 0.003962f
C1272 VDD.n666 GND 0.211938f
C1273 VDD.n667 GND 0.003962f
C1274 VDD.n668 GND 0.003962f
C1275 VDD.n669 GND 0.003962f
C1276 VDD.n670 GND 0.003962f
C1277 VDD.n671 GND 0.003962f
C1278 VDD.n672 GND 0.266884f
C1279 VDD.n673 GND 0.003962f
C1280 VDD.n674 GND 0.003962f
C1281 VDD.t83 GND 0.133442f
C1282 VDD.n675 GND 0.003962f
C1283 VDD.n676 GND 0.009601f
C1284 VDD.n677 GND 0.009601f
C1285 VDD.n678 GND 0.51022f
C1286 VDD.n688 GND 0.005826f
C1287 VDD.n689 GND 0.012127f
C1288 VDD.t32 GND 0.019391f
C1289 VDD.t31 GND 0.032488f
C1290 VDD.t30 GND 0.334077f
C1291 VDD.n690 GND 0.060478f
C1292 VDD.n691 GND 0.043121f
C1293 VDD.n692 GND 0.009566f
C1294 VDD.n693 GND 0.005826f
C1295 VDD.n694 GND 0.005826f
C1296 VDD.n695 GND 0.004689f
C1297 VDD.n696 GND 0.005826f
C1298 VDD.n697 GND 0.392477f
C1299 VDD.n698 GND 0.005826f
C1300 VDD.n699 GND 0.012127f
C1301 VDD.n700 GND 0.004689f
C1302 VDD.n701 GND 0.003892f
C1303 VDD.n702 GND 0.005826f
C1304 VDD.n703 GND 0.004689f
C1305 VDD.n704 GND 0.005826f
C1306 VDD.n705 GND 0.392477f
C1307 VDD.n706 GND 0.005826f
C1308 VDD.n707 GND 0.004689f
C1309 VDD.n708 GND 0.005826f
C1310 VDD.n709 GND 0.004689f
C1311 VDD.n710 GND 0.005826f
C1312 VDD.n711 GND 0.298283f
C1313 VDD.n712 GND 0.005826f
C1314 VDD.n713 GND 0.004689f
C1315 VDD.n714 GND 0.005826f
C1316 VDD.n715 GND 0.004689f
C1317 VDD.n716 GND 0.005826f
C1318 VDD.n717 GND 0.392477f
C1319 VDD.n718 GND 0.005826f
C1320 VDD.n719 GND 0.004689f
C1321 VDD.n720 GND 0.005826f
C1322 VDD.n721 GND 0.004689f
C1323 VDD.n722 GND 0.005826f
C1324 VDD.n723 GND 0.392477f
C1325 VDD.n724 GND 0.005826f
C1326 VDD.n725 GND 0.004689f
C1327 VDD.n726 GND 0.005826f
C1328 VDD.n727 GND 0.004689f
C1329 VDD.n728 GND 0.005826f
C1330 VDD.n729 GND 0.392477f
C1331 VDD.n730 GND 0.005826f
C1332 VDD.n731 GND 0.004689f
C1333 VDD.n732 GND 0.005826f
C1334 VDD.n733 GND 0.004689f
C1335 VDD.n734 GND 0.005826f
C1336 VDD.n735 GND 0.392477f
C1337 VDD.n736 GND 0.005826f
C1338 VDD.n737 GND 0.004689f
C1339 VDD.n738 GND 0.005826f
C1340 VDD.n739 GND 0.004689f
C1341 VDD.n740 GND 0.005826f
C1342 VDD.n741 GND 0.392477f
C1343 VDD.n742 GND 0.005826f
C1344 VDD.n743 GND 0.004689f
C1345 VDD.n744 GND 0.005826f
C1346 VDD.n745 GND 0.004689f
C1347 VDD.n746 GND 0.005826f
C1348 VDD.n747 GND 0.392477f
C1349 VDD.n748 GND 0.005826f
C1350 VDD.n749 GND 0.004689f
C1351 VDD.n750 GND 0.005826f
C1352 VDD.n751 GND 0.004689f
C1353 VDD.n752 GND 0.005826f
C1354 VDD.n753 GND 0.392477f
C1355 VDD.n754 GND 0.005826f
C1356 VDD.n755 GND 0.004689f
C1357 VDD.n756 GND 0.005826f
C1358 VDD.n757 GND 0.004689f
C1359 VDD.n758 GND 0.005826f
C1360 VDD.t59 GND 0.196239f
C1361 VDD.n759 GND 0.005826f
C1362 VDD.n760 GND 0.004689f
C1363 VDD.n761 GND 0.005826f
C1364 VDD.n762 GND 0.004689f
C1365 VDD.n763 GND 0.005826f
C1366 VDD.n764 GND 0.392477f
C1367 VDD.n765 GND 0.005826f
C1368 VDD.n766 GND 0.004689f
C1369 VDD.n767 GND 0.005826f
C1370 VDD.n768 GND 0.004689f
C1371 VDD.n769 GND 0.005826f
C1372 VDD.n770 GND 0.392477f
C1373 VDD.n771 GND 0.005826f
C1374 VDD.n772 GND 0.004689f
C1375 VDD.n773 GND 0.005826f
C1376 VDD.n774 GND 0.004689f
C1377 VDD.n775 GND 0.005826f
C1378 VDD.n776 GND 0.392477f
C1379 VDD.n777 GND 0.005826f
C1380 VDD.n778 GND 0.004689f
C1381 VDD.n779 GND 0.005826f
C1382 VDD.n780 GND 0.004689f
C1383 VDD.n781 GND 0.005826f
C1384 VDD.n782 GND 0.392477f
C1385 VDD.n783 GND 0.005826f
C1386 VDD.n784 GND 0.004689f
C1387 VDD.n785 GND 0.005826f
C1388 VDD.n786 GND 0.004689f
C1389 VDD.n787 GND 0.005826f
C1390 VDD.n788 GND 0.392477f
C1391 VDD.n789 GND 0.005826f
C1392 VDD.n790 GND 0.004689f
C1393 VDD.n791 GND 0.005826f
C1394 VDD.n792 GND 0.004689f
C1395 VDD.n793 GND 0.005826f
C1396 VDD.t64 GND 0.196239f
C1397 VDD.n794 GND 0.005826f
C1398 VDD.n795 GND 0.004689f
C1399 VDD.n796 GND 0.005826f
C1400 VDD.n797 GND 0.004689f
C1401 VDD.n798 GND 0.005826f
C1402 VDD.n799 GND 0.392477f
C1403 VDD.n800 GND 0.005826f
C1404 VDD.n801 GND 0.004689f
C1405 VDD.n802 GND 0.005826f
C1406 VDD.n803 GND 0.004689f
C1407 VDD.n804 GND 0.005826f
C1408 VDD.n805 GND 0.392477f
C1409 VDD.n806 GND 0.005826f
C1410 VDD.n807 GND 0.004689f
C1411 VDD.n808 GND 0.005826f
C1412 VDD.n809 GND 0.004689f
C1413 VDD.n810 GND 0.005826f
C1414 VDD.n811 GND 0.392477f
C1415 VDD.n812 GND 0.005826f
C1416 VDD.n813 GND 0.004689f
C1417 VDD.n814 GND 0.005826f
C1418 VDD.n815 GND 0.004689f
C1419 VDD.n816 GND 0.005826f
C1420 VDD.n817 GND 0.392477f
C1421 VDD.n818 GND 0.005826f
C1422 VDD.n819 GND 0.004689f
C1423 VDD.n820 GND 0.005826f
C1424 VDD.n821 GND 0.004689f
C1425 VDD.n822 GND 0.005826f
C1426 VDD.n823 GND 0.392477f
C1427 VDD.n824 GND 0.005826f
C1428 VDD.n825 GND 0.004689f
C1429 VDD.n826 GND 0.005826f
C1430 VDD.n827 GND 0.004689f
C1431 VDD.n828 GND 0.005826f
C1432 VDD.t70 GND 0.196239f
C1433 VDD.n829 GND 0.005826f
C1434 VDD.n830 GND 0.004689f
C1435 VDD.n831 GND 0.005826f
C1436 VDD.n832 GND 0.004689f
C1437 VDD.n833 GND 0.005826f
C1438 VDD.n834 GND 0.392477f
C1439 VDD.n835 GND 0.005826f
C1440 VDD.n836 GND 0.004689f
C1441 VDD.n837 GND 0.005826f
C1442 VDD.n838 GND 0.004689f
C1443 VDD.n839 GND 0.005826f
C1444 VDD.n840 GND 0.392477f
C1445 VDD.n841 GND 0.005826f
C1446 VDD.n842 GND 0.004689f
C1447 VDD.n843 GND 0.005826f
C1448 VDD.n844 GND 0.004689f
C1449 VDD.n845 GND 0.005826f
C1450 VDD.n846 GND 0.392477f
C1451 VDD.n847 GND 0.005826f
C1452 VDD.n848 GND 0.004689f
C1453 VDD.n849 GND 0.005826f
C1454 VDD.n850 GND 0.004689f
C1455 VDD.n851 GND 0.005826f
C1456 VDD.n852 GND 0.392477f
C1457 VDD.n853 GND 0.005826f
C1458 VDD.n854 GND 0.004689f
C1459 VDD.n855 GND 0.005826f
C1460 VDD.n856 GND 0.004689f
C1461 VDD.n857 GND 0.005826f
C1462 VDD.n858 GND 0.392477f
C1463 VDD.n859 GND 0.005826f
C1464 VDD.n860 GND 0.004689f
C1465 VDD.n861 GND 0.005826f
C1466 VDD.n862 GND 0.004689f
C1467 VDD.n863 GND 0.005826f
C1468 VDD.n864 GND 0.392477f
C1469 VDD.n865 GND 0.005826f
C1470 VDD.n866 GND 0.004689f
C1471 VDD.n867 GND 0.005826f
C1472 VDD.n868 GND 0.004689f
C1473 VDD.n869 GND 0.005826f
C1474 VDD.n870 GND 0.290433f
C1475 VDD.n871 GND 0.005826f
C1476 VDD.n872 GND 0.004689f
C1477 VDD.n873 GND 0.005826f
C1478 VDD.n874 GND 0.004689f
C1479 VDD.n875 GND 0.005826f
C1480 VDD.n876 GND 0.392477f
C1481 VDD.t9 GND 0.196239f
C1482 VDD.n877 GND 0.005826f
C1483 VDD.n878 GND 0.004689f
C1484 VDD.n879 GND 0.005826f
C1485 VDD.n880 GND 0.004689f
C1486 VDD.n881 GND 0.005826f
C1487 VDD.n882 GND 0.392477f
C1488 VDD.n883 GND 0.005826f
C1489 VDD.n884 GND 0.004689f
C1490 VDD.n885 GND 0.005826f
C1491 VDD.n886 GND 0.004689f
C1492 VDD.n887 GND 0.005826f
C1493 VDD.n888 GND 0.392477f
C1494 VDD.n889 GND 0.005826f
C1495 VDD.n890 GND 0.004689f
C1496 VDD.n891 GND 0.012459f
C1497 VDD.n892 GND 0.012459f
C1498 VDD.n893 GND 0.859525f
C1499 VDD.n894 GND 0.012459f
C1500 VDD.n895 GND 0.005826f
C1501 VDD.n897 GND 0.005826f
C1502 VDD.t47 GND 0.019391f
C1503 VDD.t48 GND 0.032488f
C1504 VDD.t46 GND 0.334077f
C1505 VDD.n898 GND 0.060478f
C1506 VDD.n899 GND 0.043121f
C1507 VDD.n900 GND 0.004689f
C1508 VDD.n901 GND 0.005826f
C1509 VDD.n902 GND 0.005826f
C1510 VDD.n903 GND 0.004689f
C1511 VDD.n905 GND 0.005826f
C1512 VDD.n906 GND 0.004689f
C1513 VDD.n907 GND 0.005826f
C1514 VDD.n908 GND 0.004689f
C1515 VDD.n909 GND 0.005826f
C1516 VDD.n910 GND 0.003118f
C1517 VDD.n911 GND 0.005826f
C1518 VDD.n912 GND 0.004689f
C1519 VDD.t10 GND 0.019391f
C1520 VDD.t11 GND 0.032488f
C1521 VDD.t8 GND 0.334077f
C1522 VDD.n913 GND 0.060478f
C1523 VDD.n914 GND 0.043121f
C1524 VDD.n915 GND 0.007221f
C1525 VDD.n916 GND 0.005826f
C1526 VDD.n917 GND 0.004689f
C1527 VDD.n918 GND 0.005826f
C1528 VDD.n919 GND 0.004689f
C1529 VDD.n920 GND 0.003892f
C1530 VDD.n922 GND 0.005826f
C1531 VDD.n923 GND 0.004689f
C1532 VDD.n924 GND 0.005826f
C1533 VDD.n925 GND 0.005826f
C1534 VDD.n926 GND 0.005826f
C1535 VDD.n927 GND 0.004689f
C1536 VDD.n928 GND 0.005826f
C1537 VDD.n930 GND 0.005826f
C1538 VDD.n932 GND 0.005826f
C1539 VDD.n933 GND 0.004689f
C1540 VDD.n934 GND 0.005826f
C1541 VDD.n935 GND 0.005826f
C1542 VDD.n936 GND 0.005826f
C1543 VDD.n937 GND 0.002368f
C1544 VDD.n938 GND 0.005826f
C1545 VDD.n940 GND 0.005826f
C1546 VDD.n942 GND 0.005826f
C1547 VDD.n943 GND 0.004689f
C1548 VDD.n944 GND 0.005826f
C1549 VDD.n945 GND 0.005826f
C1550 VDD.n946 GND 0.005826f
C1551 VDD.n947 GND 0.005826f
C1552 VDD.n948 GND 0.004689f
C1553 VDD.n949 GND 0.005826f
C1554 VDD.n951 GND 0.005826f
C1555 VDD.n952 GND 0.005826f
C1556 VDD.n954 GND 0.005826f
C1557 VDD.n955 GND 0.004689f
C1558 VDD.n956 GND 0.005826f
C1559 VDD.n957 GND 0.005826f
C1560 VDD.n958 GND 0.005826f
C1561 VDD.n959 GND 0.004056f
C1562 VDD.n960 GND 0.009566f
C1563 VDD.n961 GND 0.002978f
C1564 VDD.n962 GND 0.012459f
C1565 VDD.n963 GND 0.012127f
C1566 VDD.n964 GND 0.003892f
C1567 VDD.n965 GND 0.012127f
C1568 VDD.n966 GND 0.51022f
C1569 VDD.n967 GND 0.012127f
C1570 VDD.n968 GND 0.003892f
C1571 VDD.n969 GND 0.012127f
C1572 VDD.n970 GND 0.005826f
C1573 VDD.n971 GND 0.005826f
C1574 VDD.n972 GND 0.004689f
C1575 VDD.n973 GND 0.005826f
C1576 VDD.n974 GND 0.392477f
C1577 VDD.n975 GND 0.005826f
C1578 VDD.n976 GND 0.004689f
C1579 VDD.n977 GND 0.005826f
C1580 VDD.n978 GND 0.005826f
C1581 VDD.n979 GND 0.005826f
C1582 VDD.n980 GND 0.004689f
C1583 VDD.n981 GND 0.005826f
C1584 VDD.n982 GND 0.392477f
C1585 VDD.n983 GND 0.005826f
C1586 VDD.n984 GND 0.004689f
C1587 VDD.n985 GND 0.005826f
C1588 VDD.n986 GND 0.005826f
C1589 VDD.n987 GND 0.005826f
C1590 VDD.n988 GND 0.004689f
C1591 VDD.n989 GND 0.005826f
C1592 VDD.n990 GND 0.298283f
C1593 VDD.n991 GND 0.005826f
C1594 VDD.n992 GND 0.004689f
C1595 VDD.n993 GND 0.005826f
C1596 VDD.n994 GND 0.005826f
C1597 VDD.n995 GND 0.005826f
C1598 VDD.n996 GND 0.004689f
C1599 VDD.n997 GND 0.005826f
C1600 VDD.n998 GND 0.392477f
C1601 VDD.n999 GND 0.005826f
C1602 VDD.n1000 GND 0.004689f
C1603 VDD.n1001 GND 0.005826f
C1604 VDD.n1002 GND 0.005826f
C1605 VDD.n1003 GND 0.005826f
C1606 VDD.n1004 GND 0.004689f
C1607 VDD.n1005 GND 0.005826f
C1608 VDD.n1006 GND 0.392477f
C1609 VDD.n1007 GND 0.005826f
C1610 VDD.n1008 GND 0.004689f
C1611 VDD.n1009 GND 0.005826f
C1612 VDD.n1010 GND 0.005826f
C1613 VDD.n1011 GND 0.005826f
C1614 VDD.n1012 GND 0.004689f
C1615 VDD.n1013 GND 0.005826f
C1616 VDD.n1014 GND 0.392477f
C1617 VDD.n1015 GND 0.005826f
C1618 VDD.n1016 GND 0.004689f
C1619 VDD.n1017 GND 0.005826f
C1620 VDD.n1018 GND 0.005826f
C1621 VDD.n1019 GND 0.005826f
C1622 VDD.n1020 GND 0.004689f
C1623 VDD.n1021 GND 0.005826f
C1624 VDD.n1022 GND 0.392477f
C1625 VDD.n1023 GND 0.005826f
C1626 VDD.n1024 GND 0.004689f
C1627 VDD.n1025 GND 0.005826f
C1628 VDD.n1026 GND 0.005826f
C1629 VDD.n1027 GND 0.005826f
C1630 VDD.n1028 GND 0.004689f
C1631 VDD.n1029 GND 0.005826f
C1632 VDD.n1030 GND 0.392477f
C1633 VDD.n1031 GND 0.005826f
C1634 VDD.n1032 GND 0.004689f
C1635 VDD.n1033 GND 0.005826f
C1636 VDD.n1034 GND 0.005826f
C1637 VDD.n1035 GND 0.005826f
C1638 VDD.n1036 GND 0.004689f
C1639 VDD.n1037 GND 0.005826f
C1640 VDD.n1038 GND 0.392477f
C1641 VDD.n1039 GND 0.005826f
C1642 VDD.n1040 GND 0.004689f
C1643 VDD.n1041 GND 0.005826f
C1644 VDD.n1042 GND 0.005826f
C1645 VDD.n1043 GND 0.005826f
C1646 VDD.n1044 GND 0.004689f
C1647 VDD.n1045 GND 0.005826f
C1648 VDD.n1046 GND 0.215862f
C1649 VDD.n1047 GND 0.392477f
C1650 VDD.n1048 GND 0.005826f
C1651 VDD.n1049 GND 0.004689f
C1652 VDD.n1050 GND 0.005826f
C1653 VDD.n1051 GND 0.005826f
C1654 VDD.n1052 GND 0.005826f
C1655 VDD.n1053 GND 0.004689f
C1656 VDD.n1054 GND 0.005826f
C1657 VDD.n1055 GND 0.372853f
C1658 VDD.n1056 GND 0.005826f
C1659 VDD.n1057 GND 0.004689f
C1660 VDD.n1058 GND 0.005826f
C1661 VDD.n1059 GND 0.005826f
C1662 VDD.n1060 GND 0.005826f
C1663 VDD.n1061 GND 0.004689f
C1664 VDD.n1062 GND 0.005826f
C1665 VDD.n1063 GND 0.392477f
C1666 VDD.n1064 GND 0.005826f
C1667 VDD.n1065 GND 0.004689f
C1668 VDD.n1066 GND 0.005826f
C1669 VDD.n1067 GND 0.005826f
C1670 VDD.n1068 GND 0.005826f
C1671 VDD.n1069 GND 0.004689f
C1672 VDD.n1070 GND 0.005826f
C1673 VDD.n1071 GND 0.392477f
C1674 VDD.n1072 GND 0.005826f
C1675 VDD.n1073 GND 0.004689f
C1676 VDD.n1074 GND 0.005826f
C1677 VDD.n1075 GND 0.005826f
C1678 VDD.n1076 GND 0.005826f
C1679 VDD.n1077 GND 0.004689f
C1680 VDD.n1078 GND 0.005826f
C1681 VDD.n1079 GND 0.392477f
C1682 VDD.n1080 GND 0.005826f
C1683 VDD.n1081 GND 0.004689f
C1684 VDD.n1082 GND 0.005826f
C1685 VDD.n1083 GND 0.005826f
C1686 VDD.n1084 GND 0.005826f
C1687 VDD.n1085 GND 0.004689f
C1688 VDD.n1086 GND 0.005826f
C1689 VDD.n1087 GND 0.392477f
C1690 VDD.n1088 GND 0.005826f
C1691 VDD.n1089 GND 0.004689f
C1692 VDD.n1090 GND 0.005826f
C1693 VDD.n1091 GND 0.005826f
C1694 VDD.n1092 GND 0.005826f
C1695 VDD.n1093 GND 0.004689f
C1696 VDD.n1094 GND 0.005826f
C1697 VDD.n1095 GND 0.294358f
C1698 VDD.n1096 GND 0.392477f
C1699 VDD.n1097 GND 0.005826f
C1700 VDD.n1098 GND 0.004689f
C1701 VDD.n1099 GND 0.005826f
C1702 VDD.n1100 GND 0.004478f
C1703 VDD.n1101 GND 0.003361f
C1704 VDD.n1102 GND 0.008681f
C1705 VDD.t73 GND 0.008714f
C1706 VDD.n1103 GND 0.008524f
C1707 VDD.n1104 GND 0.002458f
C1708 VDD.n1105 GND 0.001594f
C1709 VDD.n1106 GND 0.020642f
C1710 VDD.n1107 GND 0.012681f
C1711 VDD.t72 GND 0.004713f
C1712 VDD.t69 GND 0.004713f
C1713 VDD.n1108 GND 0.017661f
C1714 VDD.n1109 GND 0.349151f
C1715 VDD.n1110 GND 0.003361f
C1716 VDD.n1111 GND 0.008681f
C1717 VDD.t60 GND 0.008714f
C1718 VDD.n1112 GND 0.008524f
C1719 VDD.n1113 GND 0.002458f
C1720 VDD.n1114 GND 0.001594f
C1721 VDD.n1115 GND 0.020642f
C1722 VDD.n1116 GND 0.012681f
C1723 VDD.t71 GND 0.004713f
C1724 VDD.t65 GND 0.004713f
C1725 VDD.n1117 GND 0.017661f
C1726 VDD.n1118 GND 0.340351f
C1727 VDD.n1119 GND 0.306254f
C1728 VDD.n1120 GND 2.34731f
C1729 VDD.n1121 GND 0.607017f
C1730 VDD.n1122 GND 0.004478f
C1731 VDD.n1123 GND 0.004689f
C1732 VDD.n1124 GND 0.005826f
C1733 VDD.n1125 GND 0.294358f
C1734 VDD.n1126 GND 0.005826f
C1735 VDD.n1127 GND 0.004689f
C1736 VDD.n1128 GND 0.005826f
C1737 VDD.n1129 GND 0.005826f
C1738 VDD.n1130 GND 0.005826f
C1739 VDD.n1131 GND 0.004689f
C1740 VDD.n1132 GND 0.005826f
C1741 VDD.n1133 GND 0.392477f
C1742 VDD.n1134 GND 0.005826f
C1743 VDD.n1135 GND 0.004689f
C1744 VDD.n1136 GND 0.005826f
C1745 VDD.n1137 GND 0.005826f
C1746 VDD.n1138 GND 0.005826f
C1747 VDD.n1139 GND 0.004689f
C1748 VDD.n1140 GND 0.005826f
C1749 VDD.n1141 GND 0.392477f
C1750 VDD.n1142 GND 0.005826f
C1751 VDD.n1143 GND 0.004689f
C1752 VDD.n1144 GND 0.005826f
C1753 VDD.n1145 GND 0.005826f
C1754 VDD.n1146 GND 0.005826f
C1755 VDD.n1147 GND 0.004689f
C1756 VDD.n1148 GND 0.005826f
C1757 VDD.n1149 GND 0.392477f
C1758 VDD.n1150 GND 0.005826f
C1759 VDD.n1151 GND 0.004689f
C1760 VDD.n1152 GND 0.005826f
C1761 VDD.n1153 GND 0.005826f
C1762 VDD.n1154 GND 0.005826f
C1763 VDD.n1155 GND 0.004689f
C1764 VDD.n1156 GND 0.005826f
C1765 VDD.n1157 GND 0.392477f
C1766 VDD.n1158 GND 0.005826f
C1767 VDD.n1159 GND 0.004689f
C1768 VDD.n1160 GND 0.005826f
C1769 VDD.n1161 GND 0.005826f
C1770 VDD.n1162 GND 0.005826f
C1771 VDD.n1163 GND 0.004689f
C1772 VDD.n1164 GND 0.005826f
C1773 VDD.n1165 GND 0.372853f
C1774 VDD.n1166 GND 0.392477f
C1775 VDD.n1167 GND 0.005826f
C1776 VDD.n1168 GND 0.004689f
C1777 VDD.n1169 GND 0.005826f
C1778 VDD.n1170 GND 0.005826f
C1779 VDD.n1171 GND 0.005826f
C1780 VDD.n1172 GND 0.004689f
C1781 VDD.n1173 GND 0.005826f
C1782 VDD.n1174 GND 0.215862f
C1783 VDD.n1175 GND 0.005826f
C1784 VDD.n1176 GND 0.004689f
C1785 VDD.n1177 GND 0.005826f
C1786 VDD.n1178 GND 0.005826f
C1787 VDD.n1179 GND 0.005826f
C1788 VDD.n1180 GND 0.004689f
C1789 VDD.n1181 GND 0.005826f
C1790 VDD.n1182 GND 0.392477f
C1791 VDD.n1183 GND 0.005826f
C1792 VDD.n1184 GND 0.004689f
C1793 VDD.n1185 GND 0.005826f
C1794 VDD.n1186 GND 0.005826f
C1795 VDD.n1187 GND 0.005826f
C1796 VDD.n1188 GND 0.004689f
C1797 VDD.n1189 GND 0.005826f
C1798 VDD.n1190 GND 0.392477f
C1799 VDD.n1191 GND 0.005826f
C1800 VDD.n1192 GND 0.004689f
C1801 VDD.n1193 GND 0.005826f
C1802 VDD.n1194 GND 0.005826f
C1803 VDD.n1195 GND 0.005826f
C1804 VDD.n1196 GND 0.004689f
C1805 VDD.n1197 GND 0.005826f
C1806 VDD.n1198 GND 0.392477f
C1807 VDD.n1199 GND 0.005826f
C1808 VDD.n1200 GND 0.004689f
C1809 VDD.n1201 GND 0.005826f
C1810 VDD.n1202 GND 0.005826f
C1811 VDD.n1203 GND 0.005826f
C1812 VDD.n1204 GND 0.004689f
C1813 VDD.n1205 GND 0.005826f
C1814 VDD.n1206 GND 0.392477f
C1815 VDD.n1207 GND 0.005826f
C1816 VDD.n1208 GND 0.004689f
C1817 VDD.n1209 GND 0.005826f
C1818 VDD.n1210 GND 0.005826f
C1819 VDD.n1211 GND 0.005826f
C1820 VDD.n1212 GND 0.004689f
C1821 VDD.n1213 GND 0.005826f
C1822 VDD.n1214 GND 0.392477f
C1823 VDD.n1215 GND 0.005826f
C1824 VDD.n1216 GND 0.004689f
C1825 VDD.n1217 GND 0.005826f
C1826 VDD.n1218 GND 0.005826f
C1827 VDD.n1219 GND 0.005826f
C1828 VDD.n1220 GND 0.004689f
C1829 VDD.n1221 GND 0.005826f
C1830 VDD.n1222 GND 0.392477f
C1831 VDD.n1223 GND 0.005826f
C1832 VDD.n1224 GND 0.004689f
C1833 VDD.n1225 GND 0.005826f
C1834 VDD.n1226 GND 0.005826f
C1835 VDD.n1227 GND 0.005826f
C1836 VDD.n1228 GND 0.004689f
C1837 VDD.n1229 GND 0.005826f
C1838 VDD.t1 GND 0.196239f
C1839 VDD.n1230 GND 0.290433f
C1840 VDD.n1231 GND 0.005826f
C1841 VDD.n1232 GND 0.004689f
C1842 VDD.n1233 GND 0.005826f
C1843 VDD.n1234 GND 0.005826f
C1844 VDD.n1235 GND 0.005826f
C1845 VDD.n1236 GND 0.004689f
C1846 VDD.n1237 GND 0.005826f
C1847 VDD.n1238 GND 0.392477f
C1848 VDD.n1239 GND 0.005826f
C1849 VDD.n1240 GND 0.004689f
C1850 VDD.n1241 GND 0.005826f
C1851 VDD.n1242 GND 0.005826f
C1852 VDD.n1243 GND 0.005826f
C1853 VDD.n1244 GND 0.005826f
C1854 VDD.n1245 GND 0.004689f
C1855 VDD.n1246 GND 0.005826f
C1856 VDD.n1247 GND 0.392477f
C1857 VDD.n1248 GND 0.005826f
C1858 VDD.n1249 GND 0.004689f
C1859 VDD.n1250 GND 0.005826f
C1860 VDD.n1251 GND 0.005826f
C1861 VDD.n1252 GND 0.005826f
C1862 VDD.n1253 GND 0.012459f
C1863 VDD.n1254 GND 0.005826f
C1864 VDD.n1255 GND 0.005826f
C1865 VDD.n1256 GND 0.004689f
C1866 VDD.n1257 GND 0.005826f
C1867 VDD.n1258 GND 0.005826f
C1868 VDD.n1259 GND 0.005826f
C1869 VDD.n1260 GND 0.005826f
C1870 VDD.n1261 GND 0.005826f
C1871 VDD.n1262 GND 0.002368f
C1872 VDD.n1263 GND 0.005826f
C1873 VDD.t3 GND 0.019391f
C1874 VDD.t2 GND 0.032488f
C1875 VDD.t0 GND 0.334077f
C1876 VDD.n1264 GND 0.060478f
C1877 VDD.n1265 GND 0.043121f
C1878 VDD.n1266 GND 0.007221f
C1879 VDD.n1267 GND 0.005826f
C1880 VDD.n1268 GND 0.005826f
C1881 VDD.n1269 GND 0.005826f
C1882 VDD.n1270 GND 0.005826f
C1883 VDD.n1271 GND 0.004689f
C1884 VDD.n1272 GND 0.005826f
C1885 VDD.n1273 GND 0.005826f
C1886 VDD.n1274 GND 0.005826f
C1887 VDD.n1275 GND 0.005826f
C1888 VDD.n1276 GND 0.005826f
C1889 VDD.n1277 GND 0.004689f
C1890 VDD.n1278 GND 0.005826f
C1891 VDD.n1279 GND 0.005826f
C1892 VDD.n1280 GND 0.004056f
C1893 VDD.n1281 GND 0.005826f
C1894 VDD.n1282 GND 0.005826f
C1895 VDD.n1283 GND 0.005826f
C1896 VDD.n1284 GND 0.004689f
C1897 VDD.n1285 GND 0.004689f
C1898 VDD.n1286 GND 0.004689f
C1899 VDD.n1287 GND 0.005826f
C1900 VDD.n1288 GND 0.005826f
C1901 VDD.n1289 GND 0.005826f
C1902 VDD.n1290 GND 0.004689f
C1903 VDD.n1291 GND 0.004689f
C1904 VDD.n1292 GND 0.003118f
C1905 VDD.n1293 GND 0.005826f
C1906 VDD.n1294 GND 0.005826f
C1907 VDD.n1295 GND 0.005826f
C1908 VDD.n1296 GND 0.004689f
C1909 VDD.n1297 GND 0.004689f
C1910 VDD.n1298 GND 0.004689f
C1911 VDD.n1299 GND 0.005826f
C1912 VDD.n1300 GND 0.005826f
C1913 VDD.n1301 GND 0.005826f
C1914 VDD.n1302 GND 0.004689f
C1915 VDD.n1303 GND 0.004689f
C1916 VDD.n1304 GND 0.003892f
C1917 VDD.n1305 GND 0.012459f
C1918 VDD.n1306 GND 0.012127f
C1919 VDD.n1307 GND 0.005826f
C1920 VDD.n1308 GND 0.004689f
C1921 VDD.n1309 GND 0.005826f
C1922 VDD.n1310 GND 0.392477f
C1923 VDD.n1311 GND 0.005826f
C1924 VDD.n1312 GND 0.004689f
C1925 VDD.n1313 GND 0.003892f
C1926 VDD.n1314 GND 0.012127f
C1927 VDD.n1315 GND 0.012459f
C1928 VDD.n1316 GND 0.002978f
C1929 VDD.n1317 GND 0.012459f
C1930 VDD.n1318 GND 2.50793f
C1931 VDD.t115 GND 3.70498f
C1932 VDD.t89 GND 2.00948f
C1933 VDD.n1319 GND 0.761405f
C1934 VDD.n1320 GND 0.008926f
C1935 VDD.n1321 GND 0.009601f
C1936 VDD.n1322 GND 0.003962f
C1937 VDD.n1323 GND 0.003059f
C1938 VDD.t51 GND 0.064081f
C1939 VDD.t52 GND 0.074164f
C1940 VDD.t49 GND 0.279207f
C1941 VDD.n1324 GND 0.052604f
C1942 VDD.n1325 GND 0.035175f
C1943 VDD.n1326 GND 0.005662f
C1944 VDD.n1327 GND 0.002884f
C1945 VDD.n1328 GND 0.003962f
C1946 VDD.n1329 GND 0.003962f
C1947 VDD.n1330 GND 0.003962f
C1948 VDD.n1331 GND 0.003962f
C1949 VDD.n1332 GND 0.003962f
C1950 VDD.n1333 GND 0.003962f
C1951 VDD.n1334 GND 0.003962f
C1952 VDD.n1335 GND 0.003962f
C1953 VDD.n1337 GND 0.003962f
C1954 VDD.n1339 GND 0.003962f
C1955 VDD.n1340 GND 0.003962f
C1956 VDD.n1341 GND 0.003962f
C1957 VDD.n1342 GND 0.003962f
C1958 VDD.n1343 GND 0.003962f
C1959 VDD.n1345 GND 0.003962f
C1960 VDD.n1347 GND 0.003962f
C1961 VDD.n1348 GND 0.003962f
C1962 VDD.n1349 GND 0.003962f
C1963 VDD.n1350 GND 0.003962f
C1964 VDD.n1351 GND 0.003962f
C1965 VDD.n1353 GND 0.003962f
C1966 VDD.n1355 GND 0.003962f
C1967 VDD.n1356 GND 0.612713f
C1968 VDD.n1357 GND 0.003962f
C1969 VDD.n1358 GND 0.003962f
C1970 VDD.n1359 GND 0.003962f
C1971 VDD.n1361 GND 0.003962f
C1972 VDD.n1363 GND 0.003962f
C1973 VDD.n1364 GND 0.003962f
C1974 VDD.n1365 GND 0.003962f
C1975 VDD.n1366 GND 0.003962f
C1976 VDD.n1367 GND 0.003962f
C1977 VDD.n1369 GND 0.003962f
C1978 VDD.n1370 GND 0.003962f
C1979 VDD.n1372 GND 0.003962f
C1980 VDD.n1373 GND 0.003962f
C1981 VDD.n1374 GND 0.009601f
C1982 VDD.n1375 GND 0.003962f
C1983 VDD.n1376 GND 0.003962f
C1984 VDD.n1377 GND 0.003962f
C1985 VDD.n1378 GND 0.003962f
C1986 VDD.n1379 GND 0.003962f
C1987 VDD.n1380 GND 0.003962f
C1988 VDD.n1381 GND 0.003962f
C1989 VDD.n1382 GND 0.003962f
C1990 VDD.n1383 GND 0.003962f
C1991 VDD.n1384 GND 0.003962f
C1992 VDD.n1385 GND 0.003962f
C1993 VDD.n1386 GND 0.003962f
C1994 VDD.n1387 GND 0.003962f
C1995 VDD.n1388 GND 0.003962f
C1996 VDD.n1389 GND 0.003962f
C1997 VDD.n1390 GND 0.003962f
C1998 VDD.n1391 GND 0.003962f
C1999 VDD.n1392 GND 0.003962f
C2000 VDD.n1393 GND 0.003962f
C2001 VDD.n1394 GND 0.003962f
C2002 VDD.n1395 GND 0.003962f
C2003 VDD.n1396 GND 0.003962f
C2004 VDD.n1397 GND 0.003962f
C2005 VDD.n1398 GND 0.003962f
C2006 VDD.n1399 GND 0.003962f
C2007 VDD.n1400 GND 0.003962f
C2008 VDD.n1401 GND 0.003962f
C2009 VDD.n1402 GND 0.003962f
C2010 VDD.n1403 GND 0.003962f
C2011 VDD.n1404 GND 0.003962f
C2012 VDD.n1405 GND 0.003962f
C2013 VDD.n1406 GND 0.003962f
C2014 VDD.n1407 GND 0.003962f
C2015 VDD.n1408 GND 0.003962f
C2016 VDD.n1409 GND 0.003962f
C2017 VDD.n1410 GND 0.003962f
C2018 VDD.n1411 GND 0.003962f
C2019 VDD.n1412 GND 0.003962f
C2020 VDD.n1413 GND 0.003962f
C2021 VDD.n1414 GND 0.003962f
C2022 VDD.n1415 GND 0.003962f
C2023 VDD.n1416 GND 0.003962f
C2024 VDD.n1417 GND 0.003962f
C2025 VDD.n1418 GND 0.003962f
C2026 VDD.n1419 GND 0.003962f
C2027 VDD.n1420 GND 0.003962f
C2028 VDD.n1421 GND 0.003962f
C2029 VDD.n1422 GND 0.003962f
C2030 VDD.n1423 GND 0.003962f
C2031 VDD.n1424 GND 0.003962f
C2032 VDD.n1425 GND 0.003962f
C2033 VDD.n1426 GND 0.003962f
C2034 VDD.n1427 GND 0.003962f
C2035 VDD.n1428 GND 0.003962f
C2036 VDD.n1429 GND 0.003962f
C2037 VDD.n1430 GND 0.003962f
C2038 VDD.n1431 GND 0.003962f
C2039 VDD.n1432 GND 0.003962f
C2040 VDD.n1433 GND 0.003962f
C2041 VDD.n1434 GND 0.003962f
C2042 VDD.n1435 GND 0.003962f
C2043 VDD.n1436 GND 0.003962f
C2044 VDD.n1437 GND 0.003962f
C2045 VDD.n1438 GND 0.003962f
C2046 VDD.n1439 GND 0.003962f
C2047 VDD.n1440 GND 0.003962f
C2048 VDD.n1441 GND 0.003962f
C2049 VDD.n1442 GND 0.003962f
C2050 VDD.n1443 GND 0.003962f
C2051 VDD.n1444 GND 0.003962f
C2052 VDD.n1445 GND 0.003962f
C2053 VDD.n1446 GND 0.003962f
C2054 VDD.n1447 GND 0.003962f
C2055 VDD.n1448 GND 0.003962f
C2056 VDD.n1449 GND 0.003962f
C2057 VDD.n1450 GND 0.008926f
C2058 VDD.n1451 GND 0.008926f
C2059 VDD.n1452 GND 0.009601f
C2060 VDD.n1453 GND 0.003962f
C2061 VDD.n1455 GND 0.003962f
C2062 VDD.n1456 GND 0.003962f
C2063 VDD.n1457 GND 0.003962f
C2064 VDD.n1458 GND 0.003962f
C2065 VDD.n1459 GND 0.003962f
C2066 VDD.n1460 GND 0.003962f
C2067 VDD.n1461 GND 0.002884f
C2068 VDD.n1462 GND 0.003962f
C2069 VDD.t54 GND 0.064081f
C2070 VDD.t55 GND 0.074164f
C2071 VDD.t53 GND 0.279207f
C2072 VDD.n1463 GND 0.052604f
C2073 VDD.n1464 GND 0.035175f
C2074 VDD.n1465 GND 0.005662f
C2075 VDD.n1466 GND 0.003962f
C2076 VDD.n1467 GND 0.003962f
C2077 VDD.n1468 GND 0.003962f
C2078 VDD.n1469 GND 0.003962f
C2079 VDD.n1470 GND 0.003962f
C2080 VDD.n1471 GND 0.003962f
C2081 VDD.n1472 GND 0.003962f
C2082 VDD.n1473 GND 0.003962f
C2083 VDD.n1474 GND 0.003962f
C2084 VDD.n1475 GND 0.003962f
C2085 VDD.n1476 GND 0.003962f
C2086 VDD.n1477 GND 0.003962f
C2087 VDD.n1478 GND 0.003962f
C2088 VDD.n1479 GND 0.003962f
C2089 VDD.n1480 GND 0.003962f
C2090 VDD.n1481 GND 0.003962f
C2091 VDD.n1482 GND 0.003962f
C2092 VDD.n1483 GND 0.003962f
C2093 VDD.n1484 GND 0.003962f
C2094 VDD.n1485 GND 0.003962f
C2095 VDD.n1486 GND 0.003962f
C2096 VDD.n1487 GND 0.003962f
C2097 VDD.n1488 GND 0.003962f
C2098 VDD.n1489 GND 0.003962f
C2099 VDD.n1490 GND 0.003962f
C2100 VDD.n1491 GND 0.003962f
C2101 VDD.n1492 GND 0.003962f
C2102 VDD.n1493 GND 0.003962f
C2103 VDD.n1494 GND 0.003962f
C2104 VDD.n1495 GND 0.003962f
C2105 VDD.n1496 GND 0.003962f
C2106 VDD.n1497 GND 0.003962f
C2107 VDD.n1498 GND 0.003962f
C2108 VDD.n1499 GND 0.003962f
C2109 VDD.n1500 GND 0.003962f
C2110 VDD.n1501 GND 0.003962f
C2111 VDD.n1502 GND 0.003962f
C2112 VDD.n1503 GND 0.003962f
C2113 VDD.n1504 GND 0.003962f
C2114 VDD.n1505 GND 0.003962f
C2115 VDD.n1506 GND 0.003962f
C2116 VDD.n1507 GND 0.003962f
C2117 VDD.n1508 GND 0.003962f
C2118 VDD.n1509 GND 0.003962f
C2119 VDD.n1510 GND 0.003962f
C2120 VDD.n1511 GND 0.003962f
C2121 VDD.n1512 GND 0.003962f
C2122 VDD.n1513 GND 0.003962f
C2123 VDD.n1514 GND 0.003962f
C2124 VDD.n1515 GND 0.003962f
C2125 VDD.n1516 GND 0.003962f
C2126 VDD.n1517 GND 0.003962f
C2127 VDD.n1518 GND 0.003962f
C2128 VDD.n1519 GND 0.003962f
C2129 VDD.n1520 GND 0.003962f
C2130 VDD.n1521 GND 0.003962f
C2131 VDD.n1522 GND 0.003962f
C2132 VDD.n1523 GND 0.003962f
C2133 VDD.n1524 GND 0.003962f
C2134 VDD.n1525 GND 0.003962f
C2135 VDD.n1526 GND 0.003962f
C2136 VDD.n1527 GND 0.003962f
C2137 VDD.n1528 GND 0.003962f
C2138 VDD.n1529 GND 0.003962f
C2139 VDD.n1530 GND 0.003962f
C2140 VDD.n1531 GND 0.003962f
C2141 VDD.n1532 GND 0.003962f
C2142 VDD.n1533 GND 0.003962f
C2143 VDD.n1534 GND 0.003962f
C2144 VDD.n1535 GND 0.003962f
C2145 VDD.n1536 GND 0.003962f
C2146 VDD.n1537 GND 0.003962f
C2147 VDD.n1538 GND 0.003962f
C2148 VDD.n1539 GND 0.003962f
C2149 VDD.n1540 GND 0.003962f
C2150 VDD.n1541 GND 0.003962f
C2151 VDD.n1542 GND 0.003962f
C2152 VDD.n1543 GND 0.003962f
C2153 VDD.n1544 GND 0.003962f
C2154 VDD.n1545 GND 0.003962f
C2155 VDD.n1546 GND 0.003962f
C2156 VDD.n1547 GND 0.003962f
C2157 VDD.n1548 GND 0.008926f
C2158 VDD.n1550 GND 0.009601f
C2159 VDD.n1551 GND 0.009601f
C2160 VDD.n1552 GND 0.003962f
C2161 VDD.n1553 GND 0.003059f
C2162 VDD.n1554 GND 0.003962f
C2163 VDD.n1556 GND 0.003962f
C2164 VDD.n1558 GND 0.003962f
C2165 VDD.n1559 GND 0.003962f
C2166 VDD.n1560 GND 0.003962f
C2167 VDD.n1561 GND 0.003962f
C2168 VDD.n1562 GND 0.003962f
C2169 VDD.n1564 GND 0.003962f
C2170 VDD.n1566 GND 0.003962f
C2171 VDD.n1567 GND 0.003962f
C2172 VDD.n1568 GND 0.003962f
C2173 VDD.n1569 GND 0.601061f
C2174 VDD.n1570 GND 0.003962f
C2175 VDD.n1572 GND 0.003962f
C2176 VDD.n1574 GND 0.003962f
C2177 VDD.n1575 GND 0.003962f
C2178 VDD.n1576 GND 0.003962f
C2179 VDD.n1577 GND 0.003962f
C2180 VDD.n1578 GND 0.003962f
C2181 VDD.n1580 GND 0.003962f
C2182 VDD.n1581 GND 0.003962f
C2183 VDD.n1582 GND 0.003962f
C2184 VDD.n1583 GND 0.003962f
C2185 VDD.n1584 GND 0.003962f
C2186 VDD.n1585 GND 0.003962f
C2187 VDD.n1587 GND 0.003962f
C2188 VDD.n1588 GND 0.003962f
C2189 VDD.n1589 GND 0.009601f
C2190 VDD.n1590 GND 0.008926f
C2191 VDD.n1591 GND 0.008926f
C2192 VDD.n1592 GND 0.396402f
C2193 VDD.n1593 GND 0.008926f
C2194 VDD.n1594 GND 0.008926f
C2195 VDD.n1595 GND 0.003962f
C2196 VDD.n1596 GND 0.003962f
C2197 VDD.n1597 GND 0.003962f
C2198 VDD.n1598 GND 0.188389f
C2199 VDD.n1599 GND 0.003962f
C2200 VDD.n1600 GND 0.003962f
C2201 VDD.n1601 GND 0.003962f
C2202 VDD.n1602 GND 0.003962f
C2203 VDD.n1603 GND 0.003962f
C2204 VDD.n1604 GND 0.266884f
C2205 VDD.n1605 GND 0.003962f
C2206 VDD.n1606 GND 0.003962f
C2207 VDD.n1607 GND 0.003962f
C2208 VDD.n1608 GND 0.003962f
C2209 VDD.n1609 GND 0.003962f
C2210 VDD.n1610 GND 0.266884f
C2211 VDD.n1611 GND 0.003962f
C2212 VDD.n1612 GND 0.003962f
C2213 VDD.n1613 GND 0.003962f
C2214 VDD.n1614 GND 0.003962f
C2215 VDD.n1615 GND 0.003962f
C2216 VDD.n1616 GND 0.266884f
C2217 VDD.n1617 GND 0.003962f
C2218 VDD.n1618 GND 0.003962f
C2219 VDD.n1619 GND 0.003962f
C2220 VDD.n1620 GND 0.003962f
C2221 VDD.n1621 GND 0.003962f
C2222 VDD.n1622 GND 0.204088f
C2223 VDD.n1623 GND 0.003962f
C2224 VDD.n1624 GND 0.003962f
C2225 VDD.n1625 GND 0.003962f
C2226 VDD.n1626 GND 0.003962f
C2227 VDD.n1627 GND 0.003962f
C2228 VDD.n1628 GND 0.266884f
C2229 VDD.n1629 GND 0.003962f
C2230 VDD.n1630 GND 0.003962f
C2231 VDD.n1631 GND 0.003962f
C2232 VDD.n1632 GND 0.003962f
C2233 VDD.n1633 GND 0.003962f
C2234 VDD.n1634 GND 0.266884f
C2235 VDD.n1635 GND 0.003962f
C2236 VDD.n1636 GND 0.003962f
C2237 VDD.n1637 GND 0.003962f
C2238 VDD.n1638 GND 0.003962f
C2239 VDD.n1639 GND 0.003962f
C2240 VDD.n1640 GND 0.176615f
C2241 VDD.n1641 GND 0.003962f
C2242 VDD.n1642 GND 0.003962f
C2243 VDD.n1643 GND 0.003962f
C2244 VDD.n1644 GND 0.003962f
C2245 VDD.n1645 GND 0.003962f
C2246 VDD.n1646 GND 0.219787f
C2247 VDD.n1647 GND 0.003962f
C2248 VDD.n1648 GND 0.003962f
C2249 VDD.n1649 GND 0.003962f
C2250 VDD.n1650 GND 0.003962f
C2251 VDD.n1651 GND 0.003962f
C2252 VDD.n1652 GND 0.266884f
C2253 VDD.n1653 GND 0.003962f
C2254 VDD.n1654 GND 0.003962f
C2255 VDD.n1655 GND 0.003962f
C2256 VDD.n1656 GND 0.003962f
C2257 VDD.n1657 GND 0.003962f
C2258 VDD.n1658 GND 0.266884f
C2259 VDD.n1659 GND 0.003962f
C2260 VDD.n1660 GND 0.003962f
C2261 VDD.n1661 GND 0.003962f
C2262 VDD.n1662 GND 0.003962f
C2263 VDD.n1663 GND 0.003962f
C2264 VDD.n1664 GND 0.192314f
C2265 VDD.n1665 GND 0.003962f
C2266 VDD.n1666 GND 0.003962f
C2267 VDD.n1667 GND 0.003962f
C2268 VDD.n1668 GND 0.003962f
C2269 VDD.n1669 GND 0.003962f
C2270 VDD.n1670 GND 0.266884f
C2271 VDD.n1671 GND 0.003962f
C2272 VDD.n1672 GND 0.003962f
C2273 VDD.n1673 GND 0.003962f
C2274 VDD.n1674 GND 0.003962f
C2275 VDD.n1675 GND 0.003962f
C2276 VDD.n1676 GND 0.266884f
C2277 VDD.n1677 GND 0.003962f
C2278 VDD.n1678 GND 0.003962f
C2279 VDD.n1679 GND 0.003962f
C2280 VDD.n1680 GND 0.003962f
C2281 VDD.n1681 GND 0.003962f
C2282 VDD.n1682 GND 0.260997f
C2283 VDD.n1683 GND 0.003962f
C2284 VDD.n1684 GND 0.003962f
C2285 VDD.n1685 GND 0.003962f
C2286 VDD.n1686 GND 0.003962f
C2287 VDD.n1687 GND 0.003962f
C2288 VDD.n1688 GND 0.208013f
C2289 VDD.n1689 GND 0.003962f
C2290 VDD.n1690 GND 0.003962f
C2291 VDD.n1691 GND 0.003962f
C2292 VDD.n1692 GND 0.003962f
C2293 VDD.n1693 GND 0.003962f
C2294 VDD.n1694 GND 0.266884f
C2295 VDD.n1695 GND 0.003962f
C2296 VDD.n1696 GND 0.003962f
C2297 VDD.n1697 GND 0.003962f
C2298 VDD.n1698 GND 0.003962f
C2299 VDD.n1699 GND 0.003962f
C2300 VDD.n1700 GND 0.266884f
C2301 VDD.n1701 GND 0.003962f
C2302 VDD.n1702 GND 0.003962f
C2303 VDD.n1703 GND 0.003962f
C2304 VDD.n1704 GND 0.003962f
C2305 VDD.n1705 GND 0.003962f
C2306 VDD.n1706 GND 0.266884f
C2307 VDD.n1707 GND 0.003962f
C2308 VDD.n1708 GND 0.003962f
C2309 VDD.n1709 GND 0.003962f
C2310 VDD.n1710 GND 0.003962f
C2311 VDD.n1711 GND 0.003962f
C2312 VDD.n1712 GND 0.2139f
C2313 VDD.n1713 GND 0.003962f
C2314 VDD.n1714 GND 0.003962f
C2315 VDD.n1715 GND 0.003962f
C2316 VDD.n1716 GND 0.003962f
C2317 VDD.n1717 GND 0.003962f
C2318 VDD.n1718 GND 0.266884f
C2319 VDD.n1719 GND 0.003962f
C2320 VDD.n1720 GND 0.003962f
C2321 VDD.n1721 GND 0.003962f
C2322 VDD.n1722 GND 0.003962f
C2323 VDD.n1723 GND 0.003962f
C2324 VDD.n1724 GND 0.266884f
C2325 VDD.n1725 GND 0.003962f
C2326 VDD.n1726 GND 0.003962f
C2327 VDD.n1727 GND 0.003962f
C2328 VDD.n1728 GND 0.003962f
C2329 VDD.n1729 GND 0.003962f
C2330 VDD.n1730 GND 0.266884f
C2331 VDD.n1731 GND 0.003962f
C2332 VDD.n1732 GND 0.003962f
C2333 VDD.n1733 GND 0.003962f
C2334 VDD.n1734 GND 0.003962f
C2335 VDD.n1735 GND 0.003962f
C2336 VDD.n1736 GND 0.241373f
C2337 VDD.n1737 GND 0.003962f
C2338 VDD.n1738 GND 0.003962f
C2339 VDD.n1739 GND 0.003962f
C2340 VDD.n1740 GND 0.003962f
C2341 VDD.n1741 GND 0.003962f
C2342 VDD.n1742 GND 0.003962f
C2343 VDD.n1743 GND 0.003962f
C2344 VDD.n1744 GND 0.266884f
C2345 VDD.n1745 GND 0.003962f
C2346 VDD.n1746 GND 0.003962f
C2347 VDD.n1747 GND 0.003962f
C2348 VDD.n1748 GND 0.003962f
C2349 VDD.n1749 GND 0.003962f
C2350 VDD.t40 GND 0.266884f
C2351 VDD.n1750 GND 0.003962f
C2352 VDD.n1751 GND 0.003962f
C2353 VDD.n1752 GND 0.003962f
C2354 VDD.n1753 GND 0.003962f
C2355 VDD.n1754 GND 0.003962f
C2356 VDD.n1755 GND 0.003962f
C2357 VDD.n1756 GND 0.003962f
C2358 VDD.n1757 GND 0.009395f
C2359 VDD.n1758 GND 0.008926f
C2360 VDD.n1759 GND 0.009601f
C2361 VDD.n1760 GND 0.009132f
C2362 VDD.n1761 GND 0.003962f
C2363 VDD.n1762 GND 0.003962f
C2364 VDD.n1763 GND 0.003962f
C2365 VDD.n1764 GND 0.003059f
C2366 VDD.n1765 GND 0.005662f
C2367 VDD.n1766 GND 0.002884f
C2368 VDD.n1767 GND 0.003962f
C2369 VDD.n1768 GND 0.003962f
C2370 VDD.n1769 GND 0.003962f
C2371 VDD.n1770 GND 0.003962f
C2372 VDD.n1771 GND 0.003962f
C2373 VDD.n1772 GND 0.003962f
C2374 VDD.n1773 GND 0.003962f
C2375 VDD.n1774 GND 0.003962f
C2376 VDD.n1775 GND 0.003962f
C2377 VDD.n1776 GND 0.003962f
C2378 VDD.n1777 GND 0.003962f
C2379 VDD.n1778 GND 0.003962f
C2380 VDD.n1779 GND 0.003962f
C2381 VDD.n1780 GND 0.003962f
C2382 VDD.n1781 GND 0.003962f
C2383 VDD.n1782 GND 0.003962f
C2384 VDD.n1783 GND 0.003962f
C2385 VDD.n1784 GND 0.003962f
C2386 VDD.n1785 GND 0.003962f
C2387 VDD.n1786 GND 0.003962f
C2388 VDD.n1787 GND 0.003962f
C2389 VDD.n1788 GND 0.003962f
C2390 VDD.n1789 GND 0.003962f
C2391 VDD.n1790 GND 0.003962f
C2392 VDD.n1791 GND 0.003962f
C2393 VDD.n1792 GND 0.003962f
C2394 VDD.n1793 GND 0.003962f
C2395 VDD.n1794 GND 0.003962f
C2396 VDD.n1795 GND 0.003962f
C2397 VDD.n1796 GND 0.003962f
C2398 VDD.n1797 GND 0.003962f
C2399 VDD.n1798 GND 0.003962f
C2400 VDD.n1799 GND 0.003962f
C2401 VDD.n1800 GND 0.009601f
C2402 VDD.n1801 GND 0.008926f
C2403 VDD.n1802 GND 0.008926f
C2404 VDD.n1803 GND 0.003962f
C2405 VDD.n1804 GND 0.003962f
C2406 VDD.n1805 GND 0.003962f
C2407 VDD.n1806 GND 0.003962f
C2408 VDD.n1807 GND 0.266884f
C2409 VDD.n1808 GND 0.003962f
C2410 VDD.n1809 GND 0.003962f
C2411 VDD.n1810 GND 0.003962f
C2412 VDD.n1811 GND 0.003962f
C2413 VDD.n1812 GND 0.003962f
C2414 VDD.n1813 GND 0.225674f
C2415 VDD.n1814 GND 0.003962f
C2416 VDD.n1815 GND 0.008926f
C2417 VDD.n1816 GND 0.009601f
C2418 VDD.n1817 GND 0.009132f
C2419 VDD.n1818 GND 0.003962f
C2420 VDD.n1819 GND 0.003962f
C2421 VDD.n1820 GND 0.003962f
C2422 VDD.n1821 GND 0.003059f
C2423 VDD.n1822 GND 0.005662f
C2424 VDD.n1823 GND 0.002884f
C2425 VDD.n1824 GND 0.003962f
C2426 VDD.n1825 GND 0.003962f
C2427 VDD.n1826 GND 0.003962f
C2428 VDD.n1827 GND 0.003962f
C2429 VDD.n1828 GND 0.003962f
C2430 VDD.n1829 GND 0.003962f
C2431 VDD.n1830 GND 0.003962f
C2432 VDD.n1831 GND 0.003962f
C2433 VDD.n1832 GND 0.003962f
C2434 VDD.n1833 GND 0.003962f
C2435 VDD.n1834 GND 0.003962f
C2436 VDD.n1835 GND 0.003962f
C2437 VDD.n1836 GND 0.003962f
C2438 VDD.n1837 GND 0.003962f
C2439 VDD.n1838 GND 0.003962f
C2440 VDD.n1839 GND 0.003962f
C2441 VDD.n1840 GND 0.003962f
C2442 VDD.n1841 GND 0.003962f
C2443 VDD.n1842 GND 0.003962f
C2444 VDD.n1843 GND 0.003962f
C2445 VDD.n1844 GND 0.003962f
C2446 VDD.n1845 GND 0.003962f
C2447 VDD.n1846 GND 0.003962f
C2448 VDD.n1847 GND 0.003962f
C2449 VDD.n1848 GND 0.003962f
C2450 VDD.n1849 GND 0.003962f
C2451 VDD.n1850 GND 0.003962f
C2452 VDD.n1851 GND 0.003962f
C2453 VDD.n1852 GND 0.003962f
C2454 VDD.n1853 GND 0.003962f
C2455 VDD.n1854 GND 0.003962f
C2456 VDD.n1855 GND 0.003962f
C2457 VDD.n1856 GND 0.009601f
C2458 VDD.n1857 GND 0.009601f
C2459 VDD.n1858 GND 1.68765f
C2460 VDD.n1859 GND 1.68765f
C2461 VDD.n1860 GND 0.008926f
C2462 VDD.n1861 GND 0.008926f
C2463 VDD.n1862 GND 0.225674f
C2464 VDD.n1863 GND 0.009601f
C2465 VDD.n1864 GND 0.003962f
C2466 VDD.n1866 GND 0.003962f
C2467 VDD.n1867 GND 0.003962f
C2468 VDD.n1868 GND 0.003962f
C2469 VDD.n1869 GND 0.003962f
C2470 VDD.n1870 GND 0.003962f
C2471 VDD.n1871 GND 0.003962f
C2472 VDD.n1872 GND 0.002884f
C2473 VDD.n1873 GND 0.003962f
C2474 VDD.t17 GND 0.064081f
C2475 VDD.t18 GND 0.074164f
C2476 VDD.t15 GND 0.279207f
C2477 VDD.n1874 GND 0.052604f
C2478 VDD.n1875 GND 0.035175f
C2479 VDD.n1876 GND 0.005662f
C2480 VDD.n1877 GND 0.003962f
C2481 VDD.n1878 GND 0.003962f
C2482 VDD.n1879 GND 0.003962f
C2483 VDD.n1880 GND 0.003962f
C2484 VDD.n1881 GND 0.003962f
C2485 VDD.n1882 GND 0.003962f
C2486 VDD.n1883 GND 0.003962f
C2487 VDD.n1884 GND 0.003962f
C2488 VDD.n1885 GND 0.003962f
C2489 VDD.n1886 GND 0.003962f
C2490 VDD.n1887 GND 0.003962f
C2491 VDD.n1888 GND 0.003962f
C2492 VDD.n1889 GND 0.003962f
C2493 VDD.n1890 GND 0.003962f
C2494 VDD.n1891 GND 0.003962f
C2495 VDD.n1892 GND 0.003962f
C2496 VDD.n1893 GND 0.003962f
C2497 VDD.n1894 GND 0.003962f
C2498 VDD.n1895 GND 0.003962f
C2499 VDD.n1896 GND 0.003962f
C2500 VDD.n1897 GND 0.003962f
C2501 VDD.n1898 GND 0.003962f
C2502 VDD.n1899 GND 0.003962f
C2503 VDD.n1900 GND 0.003962f
C2504 VDD.n1901 GND 0.003962f
C2505 VDD.n1902 GND 0.003962f
C2506 VDD.n1903 GND 0.003962f
C2507 VDD.n1904 GND 0.003962f
C2508 VDD.n1905 GND 0.003962f
C2509 VDD.n1906 GND 0.003962f
C2510 VDD.n1907 GND 0.003962f
C2511 VDD.n1908 GND 0.003962f
C2512 VDD.n1909 GND 0.003962f
C2513 VDD.n1910 GND 0.003962f
C2514 VDD.n1911 GND 0.003962f
C2515 VDD.n1912 GND 0.003962f
C2516 VDD.n1913 GND 0.003962f
C2517 VDD.n1914 GND 0.003962f
C2518 VDD.n1915 GND 0.003962f
C2519 VDD.n1916 GND 0.003962f
C2520 VDD.n1917 GND 0.003962f
C2521 VDD.n1918 GND 0.003962f
C2522 VDD.n1919 GND 0.003962f
C2523 VDD.n1920 GND 0.003962f
C2524 VDD.n1921 GND 0.003962f
C2525 VDD.n1922 GND 0.003962f
C2526 VDD.n1923 GND 0.003962f
C2527 VDD.n1924 GND 0.003962f
C2528 VDD.n1925 GND 0.003962f
C2529 VDD.n1926 GND 0.003962f
C2530 VDD.n1927 GND 0.003962f
C2531 VDD.n1928 GND 0.003962f
C2532 VDD.n1929 GND 0.003962f
C2533 VDD.n1930 GND 0.003962f
C2534 VDD.n1931 GND 0.003962f
C2535 VDD.n1932 GND 0.003962f
C2536 VDD.n1933 GND 0.003962f
C2537 VDD.n1934 GND 0.003962f
C2538 VDD.t37 GND 0.064081f
C2539 VDD.t38 GND 0.074164f
C2540 VDD.t36 GND 0.279207f
C2541 VDD.n1935 GND 0.052604f
C2542 VDD.n1936 GND 0.035175f
C2543 VDD.n1937 GND 0.003962f
C2544 VDD.n1938 GND 0.003962f
C2545 VDD.n1939 GND 0.003962f
C2546 VDD.n1940 GND 0.003962f
C2547 VDD.n1941 GND 0.003962f
C2548 VDD.n1942 GND 0.003962f
C2549 VDD.n1943 GND 0.003962f
C2550 VDD.n1945 GND 0.003962f
C2551 VDD.n1946 GND 0.003962f
C2552 VDD.n1947 GND 0.003962f
C2553 VDD.n1948 GND 0.003962f
C2554 VDD.n1950 GND 0.003962f
C2555 VDD.n1952 GND 0.003962f
C2556 VDD.n1953 GND 0.003962f
C2557 VDD.n1954 GND 0.003962f
C2558 VDD.n1955 GND 0.003962f
C2559 VDD.n1956 GND 0.003962f
C2560 VDD.n1958 GND 0.003962f
C2561 VDD.n1960 GND 0.003962f
C2562 VDD.n1961 GND 0.003962f
C2563 VDD.n1962 GND 0.003962f
C2564 VDD.n1963 GND 0.003962f
C2565 VDD.n1964 GND 0.003962f
C2566 VDD.n1966 GND 0.003962f
C2567 VDD.n1968 GND 0.003962f
C2568 VDD.n1969 GND 0.003962f
C2569 VDD.n1970 GND 0.003962f
C2570 VDD.n1971 GND 0.003962f
C2571 VDD.n1972 GND 0.003962f
C2572 VDD.n1974 GND 0.003962f
C2573 VDD.n1976 GND 0.003962f
C2574 VDD.n1977 GND 0.003962f
C2575 VDD.n1978 GND 0.002884f
C2576 VDD.n1979 GND 0.005662f
C2577 VDD.n1980 GND 0.003059f
C2578 VDD.n1981 GND 0.003962f
C2579 VDD.n1983 GND 0.003962f
C2580 VDD.n1984 GND 0.009601f
C2581 VDD.n1985 GND 0.009601f
C2582 VDD.n1986 GND 0.008926f
C2583 VDD.n1987 GND 0.003962f
C2584 VDD.n1988 GND 0.003962f
C2585 VDD.n1989 GND 0.003962f
C2586 VDD.n1990 GND 0.003962f
C2587 VDD.n1991 GND 0.003962f
C2588 VDD.n1992 GND 0.003962f
C2589 VDD.n1993 GND 0.003962f
C2590 VDD.n1994 GND 0.003962f
C2591 VDD.n1995 GND 0.003962f
C2592 VDD.n1996 GND 0.003962f
C2593 VDD.n1997 GND 0.003962f
C2594 VDD.n1998 GND 0.003962f
C2595 VDD.n1999 GND 0.003962f
C2596 VDD.n2000 GND 0.003962f
C2597 VDD.n2001 GND 0.003962f
C2598 VDD.n2002 GND 0.003962f
C2599 VDD.n2003 GND 0.003962f
C2600 VDD.n2004 GND 0.003962f
C2601 VDD.n2005 GND 0.003962f
C2602 VDD.n2006 GND 0.003962f
C2603 VDD.n2007 GND 0.003962f
C2604 VDD.n2008 GND 0.003962f
C2605 VDD.n2009 GND 0.003962f
C2606 VDD.n2010 GND 0.003962f
C2607 VDD.n2011 GND 0.003962f
C2608 VDD.n2012 GND 0.003962f
C2609 VDD.n2013 GND 0.003962f
C2610 VDD.n2014 GND 0.003962f
C2611 VDD.n2015 GND 0.003962f
C2612 VDD.n2016 GND 0.003962f
C2613 VDD.n2017 GND 0.003962f
C2614 VDD.n2018 GND 0.003962f
C2615 VDD.n2019 GND 0.003962f
C2616 VDD.n2020 GND 0.003962f
C2617 VDD.n2021 GND 0.003962f
C2618 VDD.n2022 GND 0.003962f
C2619 VDD.n2023 GND 0.003962f
C2620 VDD.n2024 GND 0.003962f
C2621 VDD.n2025 GND 0.003962f
C2622 VDD.n2026 GND 0.003962f
C2623 VDD.n2027 GND 0.003962f
C2624 VDD.n2028 GND 0.003962f
C2625 VDD.n2029 GND 0.003962f
C2626 VDD.n2030 GND 0.003962f
C2627 VDD.n2031 GND 0.003962f
C2628 VDD.n2032 GND 0.003962f
C2629 VDD.n2033 GND 0.003962f
C2630 VDD.n2034 GND 0.003962f
C2631 VDD.n2035 GND 0.003962f
C2632 VDD.n2036 GND 0.003962f
C2633 VDD.n2037 GND 0.003962f
C2634 VDD.n2038 GND 0.003962f
C2635 VDD.n2039 GND 0.003962f
C2636 VDD.n2040 GND 0.003962f
C2637 VDD.n2041 GND 0.003962f
C2638 VDD.n2042 GND 0.003962f
C2639 VDD.n2043 GND 0.003962f
C2640 VDD.n2044 GND 0.003962f
C2641 VDD.n2045 GND 0.003962f
C2642 VDD.n2046 GND 0.003962f
C2643 VDD.n2047 GND 0.003962f
C2644 VDD.n2048 GND 0.003962f
C2645 VDD.n2049 GND 0.003962f
C2646 VDD.n2050 GND 0.003962f
C2647 VDD.n2051 GND 0.003962f
C2648 VDD.n2052 GND 0.003962f
C2649 VDD.n2053 GND 0.003962f
C2650 VDD.n2054 GND 0.003962f
C2651 VDD.n2055 GND 0.003962f
C2652 VDD.n2056 GND 0.003962f
C2653 VDD.n2057 GND 0.003962f
C2654 VDD.n2058 GND 0.003962f
C2655 VDD.n2059 GND 0.003962f
C2656 VDD.n2060 GND 0.003962f
C2657 VDD.n2061 GND 0.003962f
C2658 VDD.n2062 GND 0.003962f
C2659 VDD.n2063 GND 0.2139f
C2660 VDD.n2064 GND 0.003962f
C2661 VDD.n2065 GND 0.003962f
C2662 VDD.n2066 GND 0.003962f
C2663 VDD.n2067 GND 0.003962f
C2664 VDD.n2068 GND 0.003962f
C2665 VDD.n2069 GND 0.003962f
C2666 VDD.n2070 GND 0.003962f
C2667 VDD.n2071 GND 0.003962f
C2668 VDD.n2072 GND 0.003962f
C2669 VDD.n2073 GND 0.003962f
C2670 VDD.n2074 GND 0.003962f
C2671 VDD.n2075 GND 0.003962f
C2672 VDD.n2076 GND 0.003962f
C2673 VDD.n2077 GND 0.003962f
C2674 VDD.n2078 GND 0.003962f
C2675 VDD.n2079 GND 0.003962f
C2676 VDD.n2080 GND 0.003962f
C2677 VDD.n2081 GND 0.003962f
C2678 VDD.n2082 GND 0.003962f
C2679 VDD.n2083 GND 0.003962f
C2680 VDD.n2084 GND 0.003962f
C2681 VDD.n2085 GND 0.003962f
C2682 VDD.n2086 GND 0.003962f
C2683 VDD.n2087 GND 0.003962f
C2684 VDD.n2088 GND 0.003962f
C2685 VDD.n2089 GND 0.003962f
C2686 VDD.n2090 GND 0.008926f
C2687 VDD.n2092 GND 0.009601f
C2688 VDD.n2093 GND 0.009601f
C2689 VDD.n2094 GND 0.003962f
C2690 VDD.n2095 GND 0.003059f
C2691 VDD.n2096 GND 0.003962f
C2692 VDD.n2098 GND 0.003962f
C2693 VDD.n2100 GND 0.003962f
C2694 VDD.n2101 GND 0.003962f
C2695 VDD.n2102 GND 0.003962f
C2696 VDD.n2103 GND 0.003962f
C2697 VDD.n2104 GND 0.003962f
C2698 VDD.n2106 GND 0.003962f
C2699 VDD.n2108 GND 0.003962f
C2700 VDD.n2109 GND 0.003962f
C2701 VDD.n2110 GND 0.003962f
C2702 VDD.n2111 GND 0.003962f
C2703 VDD.n2112 GND 0.003962f
C2704 VDD.n2114 GND 0.003962f
C2705 VDD.n2116 GND 0.003962f
C2706 VDD.n2117 GND 0.003962f
C2707 VDD.n2118 GND 0.003962f
C2708 VDD.n2119 GND 0.003962f
C2709 VDD.n2120 GND 0.003962f
C2710 VDD.n2122 GND 0.003962f
C2711 VDD.n2123 GND 0.003962f
C2712 VDD.n2124 GND 0.003962f
C2713 VDD.n2125 GND 0.003962f
C2714 VDD.n2126 GND 0.003962f
C2715 VDD.n2127 GND 0.003962f
C2716 VDD.n2129 GND 0.003962f
C2717 VDD.n2130 GND 0.003962f
C2718 VDD.n2131 GND 0.009601f
C2719 VDD.n2132 GND 0.008926f
C2720 VDD.n2133 GND 0.008926f
C2721 VDD.n2134 GND 0.396402f
C2722 VDD.n2135 GND 0.008926f
C2723 VDD.n2136 GND 0.008926f
C2724 VDD.n2137 GND 0.003962f
C2725 VDD.n2138 GND 0.003962f
C2726 VDD.n2139 GND 0.003962f
C2727 VDD.n2140 GND 0.174652f
C2728 VDD.n2141 GND 0.003962f
C2729 VDD.n2142 GND 0.003962f
C2730 VDD.n2143 GND 0.003962f
C2731 VDD.n2144 GND 0.003962f
C2732 VDD.n2145 GND 0.003962f
C2733 VDD.n2146 GND 0.266884f
C2734 VDD.n2147 GND 0.003962f
C2735 VDD.n2148 GND 0.003962f
C2736 VDD.n2149 GND 0.003962f
C2737 VDD.n2150 GND 0.003962f
C2738 VDD.n2151 GND 0.003962f
C2739 VDD.n2152 GND 0.266884f
C2740 VDD.n2153 GND 0.003962f
C2741 VDD.n2154 GND 0.003962f
C2742 VDD.n2155 GND 0.003962f
C2743 VDD.n2156 GND 0.003962f
C2744 VDD.n2157 GND 0.003962f
C2745 VDD.n2158 GND 0.266884f
C2746 VDD.n2159 GND 0.003962f
C2747 VDD.n2160 GND 0.003962f
C2748 VDD.n2161 GND 0.003962f
C2749 VDD.n2162 GND 0.003962f
C2750 VDD.n2163 GND 0.003962f
C2751 VDD.n2164 GND 0.158953f
C2752 VDD.n2165 GND 0.003962f
C2753 VDD.n2166 GND 0.003962f
C2754 VDD.n2167 GND 0.003962f
C2755 VDD.n2168 GND 0.003962f
C2756 VDD.n2169 GND 0.003962f
C2757 VDD.n2170 GND 0.266884f
C2758 VDD.n2171 GND 0.003962f
C2759 VDD.n2172 GND 0.003962f
C2760 VDD.n2173 GND 0.003962f
C2761 VDD.n2174 GND 0.003962f
C2762 VDD.n2175 GND 0.003962f
C2763 VDD.n2176 GND 0.266884f
C2764 VDD.n2177 GND 0.003962f
C2765 VDD.n2178 GND 0.003962f
C2766 VDD.n2179 GND 0.003962f
C2767 VDD.n2180 GND 0.003962f
C2768 VDD.n2181 GND 0.003962f
C2769 VDD.n2182 GND 0.176615f
C2770 VDD.n2183 GND 0.003962f
C2771 VDD.n2184 GND 0.003962f
C2772 VDD.n2185 GND 0.003962f
C2773 VDD.n2186 GND 0.003962f
C2774 VDD.n2187 GND 0.003962f
C2775 VDD.n2188 GND 0.143254f
C2776 VDD.n2189 GND 0.003962f
C2777 VDD.n2190 GND 0.003962f
C2778 VDD.n2191 GND 0.003962f
C2779 VDD.n2192 GND 0.003962f
C2780 VDD.n2193 GND 0.003962f
C2781 VDD.n2194 GND 0.266884f
C2782 VDD.n2195 GND 0.003962f
C2783 VDD.n2196 GND 0.003962f
C2784 VDD.n2197 GND 0.003962f
C2785 VDD.n2198 GND 0.003962f
C2786 VDD.n2199 GND 0.003962f
C2787 VDD.n2200 GND 0.266884f
C2788 VDD.n2201 GND 0.003962f
C2789 VDD.n2202 GND 0.003962f
C2790 VDD.n2203 GND 0.003962f
C2791 VDD.n2204 GND 0.003962f
C2792 VDD.n2205 GND 0.003962f
C2793 VDD.n2206 GND 0.192314f
C2794 VDD.n2207 GND 0.003962f
C2795 VDD.n2208 GND 0.003962f
C2796 VDD.n2209 GND 0.003962f
C2797 VDD.n2210 GND 0.003962f
C2798 VDD.n2211 GND 0.003962f
C2799 VDD.n2212 GND 0.139329f
C2800 VDD.n2213 GND 0.003962f
C2801 VDD.n2214 GND 0.003962f
C2802 VDD.n2215 GND 0.003962f
C2803 VDD.n2216 GND 0.003962f
C2804 VDD.n2217 GND 0.003962f
C2805 VDD.n2218 GND 0.266884f
C2806 VDD.n2219 GND 0.003962f
C2807 VDD.n2220 GND 0.003962f
C2808 VDD.n2221 GND 0.003962f
C2809 VDD.n2222 GND 0.003962f
C2810 VDD.n2223 GND 0.003962f
C2811 VDD.n2224 GND 0.266884f
C2812 VDD.n2225 GND 0.003962f
C2813 VDD.n2226 GND 0.003962f
C2814 VDD.n2227 GND 0.003962f
C2815 VDD.n2228 GND 0.003962f
C2816 VDD.n2229 GND 0.003962f
C2817 VDD.n2230 GND 0.208013f
C2818 VDD.n2231 GND 0.003962f
C2819 VDD.n2232 GND 0.003962f
C2820 VDD.n2233 GND 0.003962f
C2821 VDD.n2234 GND 0.003962f
C2822 VDD.n2235 GND 0.003962f
C2823 VDD.n2236 GND 0.266884f
C2824 VDD.n2237 GND 0.003962f
C2825 VDD.n2238 GND 0.003962f
C2826 VDD.n2239 GND 0.003962f
C2827 VDD.n2240 GND 0.003962f
C2828 VDD.n2241 GND 0.003962f
C2829 VDD.n2242 GND 0.266884f
C2830 VDD.n2243 GND 0.003962f
C2831 VDD.n2244 GND 0.003962f
C2832 VDD.n2245 GND 0.003962f
C2833 VDD.n2246 GND 0.003962f
C2834 VDD.n2247 GND 0.003962f
C2835 VDD.n2248 GND 0.180539f
C2836 VDD.n2249 GND 0.003962f
C2837 VDD.n2250 GND 0.003962f
C2838 VDD.n2251 GND 0.003962f
C2839 VDD.n2252 GND 0.003962f
C2840 VDD.n2253 GND 0.003962f
C2841 VDD.n2254 GND 0.223712f
C2842 VDD.n2255 GND 0.003962f
C2843 VDD.n2256 GND 0.003962f
C2844 VDD.n2257 GND 0.003962f
C2845 VDD.n2258 GND 0.003962f
C2846 VDD.n2259 GND 0.003962f
C2847 VDD.n2260 GND 0.266884f
C2848 VDD.n2261 GND 0.003962f
C2849 VDD.n2262 GND 0.003962f
C2850 VDD.n2263 GND 0.003962f
C2851 VDD.n2264 GND 0.003962f
C2852 VDD.n2265 GND 0.003962f
C2853 VDD.n2266 GND 0.266884f
C2854 VDD.n2267 GND 0.003962f
C2855 VDD.n2268 GND 0.003962f
C2856 VDD.n2269 GND 0.003962f
C2857 VDD.n2270 GND 0.003962f
C2858 VDD.n2271 GND 0.003962f
C2859 VDD.n2272 GND 0.196239f
C2860 VDD.n2273 GND 0.003962f
C2861 VDD.n2274 GND 0.003962f
C2862 VDD.n2275 GND 0.003962f
C2863 VDD.n2276 GND 0.003962f
C2864 VDD.n2277 GND 0.003962f
C2865 VDD.n2278 GND 0.266884f
C2866 VDD.n2279 GND 0.003962f
C2867 VDD.n2280 GND 0.003962f
C2868 VDD.n2281 GND 0.003962f
C2869 VDD.n2282 GND 0.003962f
C2870 VDD.n2283 GND 0.003962f
C2871 VDD.n2284 GND 0.003962f
C2872 VDD.n2285 GND 0.003962f
C2873 VDD.n2286 GND 0.266884f
C2874 VDD.n2287 GND 0.003962f
C2875 VDD.n2288 GND 0.003962f
C2876 VDD.n2289 GND 0.003962f
C2877 VDD.n2290 GND 0.003962f
C2878 VDD.n2291 GND 0.003962f
C2879 VDD.t24 GND 0.266884f
C2880 VDD.n2292 GND 0.003962f
C2881 VDD.n2293 GND 0.003962f
C2882 VDD.n2294 GND 0.003962f
C2883 VDD.n2295 GND 0.003962f
C2884 VDD.n2296 GND 0.003962f
C2885 VDD.n2297 GND 0.003962f
C2886 VDD.n2298 GND 0.003962f
C2887 VDD.n2299 GND 0.009395f
C2888 VDD.n2300 GND 0.008926f
C2889 VDD.n2301 GND 0.009601f
C2890 VDD.n2302 GND 0.009132f
C2891 VDD.n2303 GND 0.003962f
C2892 VDD.n2304 GND 0.003962f
C2893 VDD.n2305 GND 0.003962f
C2894 VDD.n2306 GND 0.003059f
C2895 VDD.n2307 GND 0.005662f
C2896 VDD.n2308 GND 0.002884f
C2897 VDD.n2309 GND 0.003962f
C2898 VDD.n2310 GND 0.003962f
C2899 VDD.n2311 GND 0.003962f
C2900 VDD.n2312 GND 0.003962f
C2901 VDD.n2313 GND 0.003962f
C2902 VDD.n2314 GND 0.003962f
C2903 VDD.n2315 GND 0.003962f
C2904 VDD.n2316 GND 0.003962f
C2905 VDD.n2317 GND 0.003962f
C2906 VDD.n2318 GND 0.003962f
C2907 VDD.n2319 GND 0.003962f
C2908 VDD.n2320 GND 0.003962f
C2909 VDD.n2321 GND 0.003962f
C2910 VDD.n2322 GND 0.003962f
C2911 VDD.n2323 GND -0.60479f
C2912 VDD.n2324 GND 0.003962f
C2913 VDD.n2325 GND 0.003962f
C2914 VDD.n2326 GND 0.003962f
C2915 VDD.n2327 GND 0.003962f
C2916 VDD.n2328 GND 0.003962f
C2917 VDD.n2329 GND 0.003962f
C2918 VDD.n2330 GND 0.003962f
C2919 VDD.n2331 GND 0.003962f
C2920 VDD.n2332 GND 0.003962f
C2921 VDD.n2333 GND 0.003962f
C2922 VDD.n2334 GND 0.003962f
C2923 VDD.n2335 GND 0.003962f
C2924 VDD.n2336 GND 0.003962f
C2925 VDD.n2337 GND 0.003962f
C2926 VDD.n2338 GND 0.003962f
C2927 VDD.n2339 GND 0.003962f
C2928 VDD.n2340 GND 0.003962f
C2929 VDD.n2341 GND 0.003962f
C2930 VDD.n2342 GND 0.009601f
C2931 VDD.n2343 GND 0.008926f
C2932 VDD.n2344 GND 0.008926f
C2933 VDD.n2345 GND 0.003962f
C2934 VDD.n2346 GND 0.003962f
C2935 VDD.n2347 GND 0.003962f
C2936 VDD.n2348 GND 0.003962f
C2937 VDD.n2349 GND 0.211938f
C2938 VDD.n2350 GND 0.003962f
C2939 VDD.n2351 GND 0.003962f
C2940 VDD.n2352 GND 0.003962f
C2941 VDD.n2353 GND 0.003962f
C2942 VDD.n2354 GND 0.003962f
C2943 VDD.n2355 GND 0.266884f
C2944 VDD.n2356 GND 0.003962f
C2945 VDD.n2357 GND 0.008926f
C2946 VDD.n2358 GND 0.009601f
C2947 VDD.n2359 GND 0.009132f
C2948 VDD.n2360 GND 0.003962f
C2949 VDD.n2361 GND 0.003962f
C2950 VDD.n2362 GND 0.003962f
C2951 VDD.n2363 GND 0.003059f
C2952 VDD.n2364 GND 0.005662f
C2953 VDD.n2365 GND 0.002884f
C2954 VDD.n2366 GND 0.003962f
C2955 VDD.n2367 GND 0.003962f
C2956 VDD.n2368 GND 0.003962f
C2957 VDD.n2369 GND 0.003962f
C2958 VDD.n2370 GND 0.003962f
C2959 VDD.n2371 GND 0.003962f
C2960 VDD.n2372 GND 0.003962f
C2961 VDD.n2373 GND 0.003962f
C2962 VDD.n2374 GND 0.003962f
C2963 VDD.n2375 GND 0.003962f
C2964 VDD.n2376 GND 0.003962f
C2965 VDD.n2377 GND 0.003962f
C2966 VDD.n2378 GND 0.003962f
C2967 VDD.n2379 GND 0.003962f
C2968 VDD.n2380 GND -0.593138f
C2969 VDD.n2381 GND 0.003962f
C2970 VDD.n2382 GND 0.003962f
C2971 VDD.n2383 GND 0.003962f
C2972 VDD.n2384 GND 0.003962f
C2973 VDD.n2385 GND 0.003962f
C2974 VDD.n2386 GND 0.003962f
C2975 VDD.n2387 GND 0.003962f
C2976 VDD.n2388 GND 0.003962f
C2977 VDD.n2389 GND 0.003962f
C2978 VDD.n2390 GND 0.003962f
C2979 VDD.n2391 GND 0.003962f
C2980 VDD.n2392 GND 0.003962f
C2981 VDD.n2393 GND 0.003962f
C2982 VDD.n2394 GND 0.003962f
C2983 VDD.n2395 GND 0.003962f
C2984 VDD.n2396 GND 0.003962f
C2985 VDD.n2397 GND 0.003962f
C2986 VDD.n2398 GND 0.009601f
C2987 VDD.n2399 GND 0.009601f
C2988 VDD.n2400 GND 0.761405f
C2989 VDD.t105 GND 2.00948f
C2990 VDD.t56 GND 3.70498f
C2991 VDD.n2401 GND 2.50793f
C2992 VDD.n2402 GND 0.012459f
C2993 VDD.n2403 GND 0.005826f
C2994 VDD.n2404 GND 0.004689f
C2995 VDD.n2406 GND 0.005826f
C2996 VDD.n2407 GND 0.005826f
C2997 VDD.n2408 GND 0.005826f
C2998 VDD.n2409 GND 0.004689f
C2999 VDD.n2410 GND 0.005826f
C3000 VDD.n2411 GND 0.005826f
C3001 VDD.n2412 GND 0.005826f
C3002 VDD.n2413 GND 0.005826f
C3003 VDD.t21 GND 0.019391f
C3004 VDD.t22 GND 0.032488f
C3005 VDD.t19 GND 0.334077f
C3006 VDD.n2414 GND 0.060478f
C3007 VDD.n2415 GND 0.043121f
C3008 VDD.n2416 GND 0.005826f
C3009 VDD.n2417 GND 0.004689f
C3010 VDD.n2418 GND 0.005826f
C3011 VDD.n2419 GND 0.005826f
C3012 VDD.n2420 GND 0.005826f
C3013 VDD.n2421 GND 0.005826f
C3014 VDD.n2422 GND 0.005826f
C3015 VDD.n2423 GND 0.004689f
C3016 VDD.n2424 GND 0.005826f
C3017 VDD.n2425 GND 0.005826f
C3018 VDD.n2426 GND 0.005826f
C3019 VDD.n2427 GND 0.005826f
C3020 VDD.n2429 GND 0.005826f
C3021 VDD.n2430 GND 0.002978f
C3022 VDD.n2432 GND 0.005826f
C3023 VDD.t34 GND 0.019391f
C3024 VDD.t35 GND 0.032488f
C3025 VDD.t33 GND 0.334077f
C3026 VDD.n2433 GND 0.060478f
C3027 VDD.n2434 GND 0.043121f
C3028 VDD.n2435 GND 0.009566f
C3029 VDD.n2436 GND 0.005826f
C3030 VDD.n2437 GND 0.005826f
C3031 VDD.n2438 GND 0.004056f
C3032 VDD.n2439 GND 0.004689f
C3033 VDD.n2440 GND 0.004689f
C3034 VDD.n2441 GND 0.005826f
C3035 VDD.n2443 GND 0.005826f
C3036 VDD.n2445 GND 0.005826f
C3037 VDD.n2446 GND 0.004689f
C3038 VDD.n2447 GND 0.004689f
C3039 VDD.n2448 GND 0.004689f
C3040 VDD.n2449 GND 0.005826f
C3041 VDD.n2451 GND 0.005826f
C3042 VDD.n2453 GND 0.005826f
C3043 VDD.n2454 GND 0.003118f
C3044 VDD.n2455 GND 0.007221f
C3045 VDD.n2456 GND 0.002368f
C3046 VDD.n2457 GND 0.004689f
C3047 VDD.n2458 GND 0.005826f
C3048 VDD.n2460 GND 0.005826f
C3049 VDD.n2461 GND 0.005826f
C3050 VDD.n2462 GND 0.004689f
C3051 VDD.n2463 GND 0.004689f
C3052 VDD.n2464 GND 0.005826f
C3053 VDD.n2465 GND 0.005826f
C3054 VDD.n2467 GND 0.005826f
C3055 VDD.n2468 GND 0.004689f
C3056 VDD.n2469 GND 0.003892f
C3057 VDD.n2470 GND 0.012459f
C3058 VDD.n2471 GND 0.012127f
C3059 VDD.n2472 GND 0.003892f
C3060 VDD.n2473 GND 0.012127f
C3061 VDD.n2474 GND 0.51022f
C3062 VDD.n2475 GND 0.012127f
C3063 VDD.n2476 GND 0.003892f
C3064 VDD.n2477 GND 0.012127f
C3065 VDD.n2478 GND 0.005826f
C3066 VDD.n2479 GND 0.005826f
C3067 VDD.n2480 GND 0.004689f
C3068 VDD.n2481 GND 0.005826f
C3069 VDD.n2482 GND 0.392477f
C3070 VDD.n2483 GND 0.005826f
C3071 VDD.n2484 GND 0.004689f
C3072 VDD.n2485 GND 0.005826f
C3073 VDD.n2486 GND 0.005826f
C3074 VDD.n2487 GND 0.005826f
C3075 VDD.n2488 GND 0.004689f
C3076 VDD.n2489 GND 0.005826f
C3077 VDD.n2490 GND 0.392477f
C3078 VDD.n2491 GND 0.005826f
C3079 VDD.n2492 GND 0.004689f
C3080 VDD.n2493 GND 0.005826f
C3081 VDD.n2494 GND 0.005826f
C3082 VDD.n2495 GND 0.005826f
C3083 VDD.n2496 GND 0.004689f
C3084 VDD.n2497 GND 0.005826f
C3085 VDD.t20 GND 0.196239f
C3086 VDD.n2498 GND 0.298283f
C3087 VDD.n2499 GND 0.005826f
C3088 VDD.n2500 GND 0.004689f
C3089 VDD.n2501 GND 0.005826f
C3090 VDD.n2502 GND 0.005826f
C3091 VDD.n2503 GND 0.005826f
C3092 VDD.n2504 GND 0.004689f
C3093 VDD.n2505 GND 0.005826f
C3094 VDD.n2506 GND 0.392477f
C3095 VDD.n2507 GND 0.005826f
C3096 VDD.n2508 GND 0.004689f
C3097 VDD.n2509 GND 0.005826f
C3098 VDD.n2510 GND 0.005826f
C3099 VDD.n2511 GND 0.005826f
C3100 VDD.n2512 GND 0.004689f
C3101 VDD.n2513 GND 0.005826f
C3102 VDD.n2514 GND 0.392477f
C3103 VDD.n2515 GND 0.005826f
C3104 VDD.n2516 GND 0.004689f
C3105 VDD.n2517 GND 0.005826f
C3106 VDD.n2518 GND 0.005826f
C3107 VDD.n2519 GND 0.005826f
C3108 VDD.n2520 GND 0.004689f
C3109 VDD.n2521 GND 0.005826f
C3110 VDD.n2522 GND 0.392477f
C3111 VDD.n2523 GND 0.005826f
C3112 VDD.n2524 GND 0.004689f
C3113 VDD.n2525 GND 0.005826f
C3114 VDD.n2526 GND 0.005826f
C3115 VDD.n2527 GND 0.005826f
C3116 VDD.n2528 GND 0.004689f
C3117 VDD.n2529 GND 0.005826f
C3118 VDD.n2530 GND 0.392477f
C3119 VDD.n2531 GND 0.005826f
C3120 VDD.n2532 GND 0.004689f
C3121 VDD.n2533 GND 0.005826f
C3122 VDD.n2534 GND 0.005826f
C3123 VDD.n2535 GND 0.005826f
C3124 VDD.n2536 GND 0.004689f
C3125 VDD.n2537 GND 0.005826f
C3126 VDD.n2538 GND 0.392477f
C3127 VDD.n2539 GND 0.005826f
C3128 VDD.n2540 GND 0.004689f
C3129 VDD.n2541 GND 0.005826f
C3130 VDD.n2542 GND 0.005826f
C3131 VDD.n2543 GND 0.005826f
C3132 VDD.n2544 GND 0.004689f
C3133 VDD.n2545 GND 0.005826f
C3134 VDD.n2546 GND 0.392477f
C3135 VDD.n2547 GND 0.005826f
C3136 VDD.n2548 GND 0.004689f
C3137 VDD.n2549 GND 0.005826f
C3138 VDD.n2550 GND 0.005826f
C3139 VDD.n2551 GND 0.005826f
C3140 VDD.n2552 GND 0.004689f
C3141 VDD.n2553 GND 0.005826f
C3142 VDD.n2554 GND 0.392477f
C3143 VDD.n2555 GND 0.005826f
C3144 VDD.n2556 GND 0.004689f
C3145 VDD.n2557 GND 0.005826f
C3146 VDD.n2558 GND 0.005826f
C3147 VDD.n2559 GND 0.005826f
C3148 VDD.n2560 GND 0.004689f
C3149 VDD.n2561 GND 0.005826f
C3150 VDD.n2562 GND 0.372853f
C3151 VDD.n2563 GND 0.005826f
C3152 VDD.n2564 GND 0.004689f
C3153 VDD.n2565 GND 0.005826f
C3154 VDD.n2566 GND 0.005826f
C3155 VDD.n2567 GND 0.005826f
C3156 VDD.n2568 GND 0.004689f
C3157 VDD.n2569 GND 0.005826f
C3158 VDD.n2570 GND 0.392477f
C3159 VDD.n2571 GND 0.005826f
C3160 VDD.n2572 GND 0.004689f
C3161 VDD.n2573 GND 0.005826f
C3162 VDD.n2574 GND 0.005826f
C3163 VDD.n2575 GND 0.005826f
C3164 VDD.n2576 GND 0.004689f
C3165 VDD.n2577 GND 0.005826f
C3166 VDD.n2578 GND 0.392477f
C3167 VDD.n2579 GND 0.005826f
C3168 VDD.n2580 GND 0.004689f
C3169 VDD.n2581 GND 0.005826f
C3170 VDD.n2582 GND 0.005826f
C3171 VDD.n2583 GND 0.005826f
C3172 VDD.n2584 GND 0.004689f
C3173 VDD.n2585 GND 0.005826f
C3174 VDD.n2586 GND 0.392477f
C3175 VDD.n2587 GND 0.005826f
C3176 VDD.n2588 GND 0.004689f
C3177 VDD.n2589 GND 0.005826f
C3178 VDD.n2590 GND 0.005826f
C3179 VDD.n2591 GND 0.005826f
C3180 VDD.n2592 GND 0.005826f
C3181 VDD.n2593 GND 0.005826f
C3182 VDD.n2594 GND 0.004689f
C3183 VDD.n2595 GND 0.004689f
C3184 VDD.n2596 GND 0.005826f
C3185 VDD.n2597 GND 0.392477f
C3186 VDD.n2598 GND 0.005826f
C3187 VDD.n2599 GND 0.004689f
C3188 VDD.n2600 GND 0.005826f
C3189 VDD.n2601 GND 0.005826f
C3190 VDD.n2602 GND 0.005826f
C3191 VDD.n2603 GND 0.004689f
C3192 VDD.n2604 GND 0.005826f
C3193 VDD.n2605 GND 0.392477f
C3194 VDD.n2606 GND 0.294358f
C3195 VDD.n2607 GND 0.005826f
C3196 VDD.n2608 GND 0.004689f
C3197 VDD.n2609 GND 0.004689f
C3198 VDD.n2610 GND 0.004689f
C3199 VDD.n2611 GND 0.005826f
C3200 VDD.n2612 GND 0.005826f
C3201 VDD.n2613 GND 0.005826f
C3202 VDD.n2614 GND 0.005826f
C3203 VDD.n2615 GND 0.004689f
C3204 VDD.n2616 GND 0.004689f
C3205 VDD.n2617 GND 0.004689f
C3206 VDD.n2618 GND 0.005826f
C3207 VDD.n2619 GND 0.005826f
C3208 VDD.n2620 GND 0.005826f
C3209 VDD.n2621 GND 0.005826f
C3210 VDD.n2622 GND 0.004689f
C3211 VDD.n2623 GND 0.004689f
C3212 VDD.n2624 GND 0.004689f
C3213 VDD.n2625 GND 0.005826f
C3214 VDD.n2626 GND 0.005826f
C3215 VDD.n2627 GND 0.005826f
C3216 VDD.n2628 GND 0.005826f
C3217 VDD.n2629 GND 0.004689f
C3218 VDD.n2630 GND 0.004689f
C3219 VDD.n2631 GND 0.004689f
C3220 VDD.n2632 GND 0.005826f
C3221 VDD.n2633 GND 0.005826f
C3222 VDD.n2634 GND 0.005826f
C3223 VDD.n2635 GND 0.005826f
C3224 VDD.n2636 GND 0.004689f
C3225 VDD.n2637 GND 0.004689f
C3226 VDD.n2638 GND 0.004689f
C3227 VDD.n2639 GND 0.005826f
C3228 VDD.n2640 GND 0.005826f
C3229 VDD.n2641 GND 0.005826f
C3230 VDD.n2642 GND 0.005826f
C3231 VDD.n2643 GND 0.004689f
C3232 VDD.n2644 GND 0.004689f
C3233 VDD.n2645 GND 0.004689f
C3234 VDD.n2646 GND 0.005826f
C3235 VDD.n2647 GND 0.005826f
C3236 VDD.n2648 GND 0.005826f
C3237 VDD.n2649 GND 0.005826f
C3238 VDD.n2650 GND 0.004689f
C3239 VDD.n2651 GND 0.004689f
C3240 VDD.n2652 GND 0.004689f
C3241 VDD.n2653 GND 0.005826f
C3242 VDD.n2654 GND 0.005826f
C3243 VDD.n2655 GND 0.005826f
C3244 VDD.n2656 GND 0.005826f
C3245 VDD.n2657 GND 0.004689f
C3246 VDD.n2658 GND 0.004689f
C3247 VDD.n2659 GND 0.004689f
C3248 VDD.n2660 GND 0.005826f
C3249 VDD.n2661 GND 0.005826f
C3250 VDD.n2662 GND 0.005826f
C3251 VDD.n2663 GND 0.005826f
C3252 VDD.n2664 GND 0.004689f
C3253 VDD.n2665 GND 0.004689f
C3254 VDD.n2666 GND 0.003892f
C3255 VDD.n2667 GND 0.012127f
C3256 VDD.n2668 GND 0.012459f
C3257 VDD.n2669 GND 0.005826f
C3258 VDD.n2670 GND 0.009566f
C3259 VDD.n2671 GND 0.005826f
C3260 VDD.n2672 GND 0.005826f
C3261 VDD.n2673 GND 0.004056f
C3262 VDD.n2674 GND 0.004689f
C3263 VDD.n2675 GND 0.005826f
C3264 VDD.n2676 GND 0.005826f
C3265 VDD.n2677 GND 0.004689f
C3266 VDD.n2678 GND 0.004689f
C3267 VDD.n2679 GND 0.005826f
C3268 VDD.n2680 GND 0.005826f
C3269 VDD.n2681 GND 0.004689f
C3270 VDD.n2682 GND 0.004689f
C3271 VDD.n2683 GND 0.005826f
C3272 VDD.n2684 GND 0.005826f
C3273 VDD.n2685 GND 0.004689f
C3274 VDD.n2686 GND 0.004689f
C3275 VDD.n2687 GND 0.005826f
C3276 VDD.n2688 GND 0.005826f
C3277 VDD.n2689 GND 0.003118f
C3278 VDD.t14 GND 0.019391f
C3279 VDD.t13 GND 0.032488f
C3280 VDD.t12 GND 0.334077f
C3281 VDD.n2690 GND 0.060478f
C3282 VDD.n2691 GND 0.043121f
C3283 VDD.n2692 GND 0.007221f
C3284 VDD.n2693 GND 0.002368f
C3285 VDD.n2694 GND 0.005826f
C3286 VDD.n2695 GND 0.005826f
C3287 VDD.n2696 GND 0.004689f
C3288 VDD.n2697 GND 0.004689f
C3289 VDD.n2698 GND 0.005826f
C3290 VDD.n2699 GND 0.005826f
C3291 VDD.n2700 GND 0.004689f
C3292 VDD.n2701 GND 0.005826f
C3293 VDD.n2702 GND 0.005826f
C3294 VDD.n2703 GND 0.004689f
C3295 VDD.n2704 GND 0.005826f
C3296 VDD.n2705 GND 0.005826f
C3297 VDD.n2706 GND 0.005826f
C3298 VDD.n2707 GND 0.004689f
C3299 VDD.n2708 GND 0.003892f
C3300 VDD.n2709 GND 0.012459f
C3301 VDD.n2710 GND 0.859525f
C3302 VDD.n2711 GND 0.51022f
C3303 VDD.n2712 GND 0.392477f
C3304 VDD.n2713 GND 0.005826f
C3305 VDD.n2714 GND 0.004689f
C3306 VDD.n2715 GND 0.004689f
C3307 VDD.n2716 GND 0.004689f
C3308 VDD.n2717 GND 0.005826f
C3309 VDD.n2718 GND 0.392477f
C3310 VDD.n2719 GND 0.392477f
C3311 VDD.n2720 GND 0.392477f
C3312 VDD.n2721 GND 0.005826f
C3313 VDD.n2722 GND 0.004689f
C3314 VDD.n2723 GND 0.004689f
C3315 VDD.n2724 GND 0.004689f
C3316 VDD.n2725 GND 0.005826f
C3317 VDD.n2726 GND 0.290433f
C3318 VDD.n2727 GND 0.392477f
C3319 VDD.n2728 GND 0.392477f
C3320 VDD.n2729 GND 0.005826f
C3321 VDD.n2730 GND 0.004689f
C3322 VDD.n2731 GND 0.004689f
C3323 VDD.n2732 GND 0.004689f
C3324 VDD.n2733 GND 0.005826f
C3325 VDD.n2734 GND 0.392477f
C3326 VDD.n2735 GND 0.392477f
C3327 VDD.n2736 GND 0.392477f
C3328 VDD.n2737 GND 0.005826f
C3329 VDD.n2738 GND 0.004689f
C3330 VDD.n2739 GND 0.004689f
C3331 VDD.n2740 GND 0.004689f
C3332 VDD.n2741 GND 0.005826f
C3333 VDD.n2742 GND 0.392477f
C3334 VDD.n2743 GND 0.392477f
C3335 VDD.n2744 GND 0.392477f
C3336 VDD.n2745 GND 0.005826f
C3337 VDD.n2746 GND 0.004689f
C3338 VDD.n2747 GND 0.004689f
C3339 VDD.n2748 GND 0.004689f
C3340 VDD.n2749 GND 0.005826f
C3341 VDD.n2750 GND 0.392477f
C3342 VDD.n2751 GND 0.392477f
C3343 VDD.n2752 GND 0.215862f
C3344 VDD.n2753 GND 0.005826f
C3345 VDD.n2754 GND 0.004689f
C3346 VDD.n2755 GND 0.004689f
C3347 VDD.n2756 GND 0.004689f
C3348 VDD.n2757 GND 0.005826f
C3349 VDD.n2758 GND 0.392477f
C3350 VDD.n2759 GND 0.392477f
C3351 VDD.n2760 GND 0.392477f
C3352 VDD.n2761 GND 0.005826f
C3353 VDD.n2762 GND 0.004689f
C3354 VDD.n2763 GND 0.004689f
C3355 VDD.n2764 GND 0.004689f
C3356 VDD.n2765 GND 0.005826f
C3357 VDD.n2766 GND 0.392477f
C3358 VDD.n2767 GND 0.392477f
C3359 VDD.n2768 GND 0.392477f
C3360 VDD.n2769 GND 0.005826f
C3361 VDD.n2770 GND 0.004689f
C3362 VDD.n2771 GND 0.004689f
C3363 VDD.n2772 GND 0.004689f
C3364 VDD.n2773 GND 0.005826f
C3365 VDD.n2774 GND 0.392477f
C3366 VDD.n2775 GND 0.392477f
C3367 VDD.n2776 GND 0.294358f
C3368 VDD.n2777 GND 0.005826f
C3369 VDD.n2778 GND 0.004689f
C3370 VDD.n2779 GND 0.004478f
C3371 VDD.n2780 GND 0.607017f
C3372 VDD.n2781 GND 2.34126f
C3373 a_n11986_8880.n0 GND 0.641477f
C3374 a_n11986_8880.n1 GND 0.26761f
C3375 a_n11986_8880.n2 GND 0.641477f
C3376 a_n11986_8880.n3 GND 0.26761f
C3377 a_n11986_8880.n4 GND 0.147859f
C3378 a_n11986_8880.n5 GND 0.546717f
C3379 a_n11986_8880.n6 GND 0.392023f
C3380 a_n11986_8880.n7 GND 0.147859f
C3381 a_n11986_8880.n8 GND 0.585968f
C3382 a_n11986_8880.n9 GND 0.392023f
C3383 a_n11986_8880.n10 GND 0.147859f
C3384 a_n11986_8880.n11 GND 0.546717f
C3385 a_n11986_8880.n12 GND 0.392023f
C3386 a_n11986_8880.n13 GND 0.147859f
C3387 a_n11986_8880.n14 GND 0.585968f
C3388 a_n11986_8880.n15 GND 0.392023f
C3389 a_n11986_8880.n16 GND 0.265688f
C3390 a_n11986_8880.n17 GND 0.265688f
C3391 a_n11986_8880.n18 GND 0.493618f
C3392 a_n11986_8880.n19 GND 0.147859f
C3393 a_n11986_8880.n20 GND 0.227534f
C3394 a_n11986_8880.n21 GND 0.245714f
C3395 a_n11986_8880.n22 GND 0.493618f
C3396 a_n11986_8880.n23 GND 0.147859f
C3397 a_n11986_8880.n24 GND 0.227534f
C3398 a_n11986_8880.n25 GND 0.245714f
C3399 a_n11986_8880.n26 GND 2.63641f
C3400 a_n11986_8880.n27 GND 0.133744f
C3401 a_n11986_8880.n28 GND 0.133744f
C3402 a_n11986_8880.t12 GND 0.048315f
C3403 a_n11986_8880.t10 GND 0.048315f
C3404 a_n11986_8880.t9 GND 0.048315f
C3405 a_n11986_8880.n29 GND 0.324348f
C3406 a_n11986_8880.t11 GND 0.048315f
C3407 a_n11986_8880.t6 GND 0.048315f
C3408 a_n11986_8880.n30 GND 0.318253f
C3409 a_n11986_8880.n31 GND 2.78493f
C3410 a_n11986_8880.t0 GND 0.503282f
C3411 a_n11986_8880.t5 GND 0.503281f
C3412 a_n11986_8880.t4 GND 0.047062f
C3413 a_n11986_8880.t2 GND 0.047062f
C3414 a_n11986_8880.n32 GND 0.398361f
C3415 a_n11986_8880.n33 GND 2.12942f
C3416 a_n11986_8880.t3 GND 0.047062f
C3417 a_n11986_8880.t1 GND 0.047062f
C3418 a_n11986_8880.n34 GND 0.397206f
C3419 a_n11986_8880.t24 GND 1.38852f
C3420 a_n11986_8880.t17 GND 1.65625f
C3421 a_n11986_8880.n35 GND 1.08316f
C3422 a_n11986_8880.t21 GND 1.01956f
C3423 a_n11986_8880.n36 GND 0.691096f
C3424 a_n11986_8880.t15 GND 1.38852f
C3425 a_n11986_8880.t16 GND 1.65625f
C3426 a_n11986_8880.n37 GND 1.08316f
C3427 a_n11986_8880.t18 GND 1.01956f
C3428 a_n11986_8880.n38 GND 0.691096f
C3429 a_n11986_8880.n39 GND 1.56439f
C3430 a_n11986_8880.t20 GND 1.38852f
C3431 a_n11986_8880.t22 GND 1.65624f
C3432 a_n11986_8880.n40 GND 1.08316f
C3433 a_n11986_8880.t25 GND 1.01956f
C3434 a_n11986_8880.n41 GND 0.617402f
C3435 a_n11986_8880.t19 GND 1.38852f
C3436 a_n11986_8880.t14 GND 1.65624f
C3437 a_n11986_8880.n42 GND 1.08316f
C3438 a_n11986_8880.t23 GND 1.01956f
C3439 a_n11986_8880.n43 GND 0.617402f
C3440 a_n11986_8880.n44 GND 1.3157f
C3441 a_n11986_8880.n45 GND 16.2876f
C3442 a_n11986_8880.n46 GND 3.17065f
C3443 a_n11986_8880.n47 GND 5.60394f
C3444 a_n11986_8880.t8 GND 0.048315f
C3445 a_n11986_8880.t7 GND 0.048315f
C3446 a_n11986_8880.n48 GND 0.318253f
C3447 a_n11986_8880.n49 GND 3.36656f
C3448 a_n11986_8880.n50 GND 0.324348f
C3449 a_n11986_8880.t13 GND 0.048315f
C3450 a_n3584_7550.n0 GND 2.69399f
C3451 a_n3584_7550.n1 GND 4.9628f
C3452 a_n3584_7550.n2 GND 2.36221f
C3453 a_n3584_7550.n3 GND 1.77427f
C3454 a_n3584_7550.t0 GND 74.3692f
C3455 a_n3584_7550.t3 GND 0.275118f
C3456 a_n3584_7550.t15 GND 0.035314f
C3457 a_n3584_7550.t11 GND 0.035314f
C3458 a_n3584_7550.n4 GND 0.193365f
C3459 a_n3584_7550.t8 GND 0.271241f
C3460 a_n3584_7550.t5 GND 0.275118f
C3461 a_n3584_7550.t12 GND 0.035314f
C3462 a_n3584_7550.t6 GND 0.035314f
C3463 a_n3584_7550.n5 GND 0.193365f
C3464 a_n3584_7550.t9 GND 0.271241f
C3465 a_n3584_7550.t4 GND 0.271241f
C3466 a_n3584_7550.t7 GND 0.035314f
C3467 a_n3584_7550.t14 GND 0.035314f
C3468 a_n3584_7550.n6 GND 0.193365f
C3469 a_n3584_7550.t13 GND 0.271241f
C3470 a_n3584_7550.t10 GND 0.271241f
C3471 a_n3584_7550.t16 GND 0.035314f
C3472 a_n3584_7550.t2 GND 0.035314f
C3473 a_n3584_7550.n7 GND 0.193365f
C3474 a_n3584_7550.t1 GND 0.275118f
C3475 a_n5004_9136.n0 GND 1.70425f
C3476 a_n5004_9136.n1 GND 3.80246f
C3477 a_n5004_9136.n2 GND 0.489851f
C3478 a_n5004_9136.n3 GND 2.19274f
C3479 a_n5004_9136.n4 GND 0.489851f
C3480 a_n5004_9136.n5 GND 0.724788f
C3481 a_n5004_9136.n6 GND 1.46795f
C3482 a_n5004_9136.n7 GND 0.48985f
C3483 a_n5004_9136.n8 GND 0.48985f
C3484 a_n5004_9136.n9 GND 1.67848f
C3485 a_n5004_9136.n10 GND 0.48985f
C3486 a_n5004_9136.n11 GND 1.7902f
C3487 a_n5004_9136.n12 GND 0.48985f
C3488 a_n5004_9136.n13 GND 1.55584f
C3489 a_n5004_9136.n14 GND 0.48985f
C3490 a_n5004_9136.n15 GND 0.48985f
C3491 a_n5004_9136.n16 GND 0.48985f
C3492 a_n5004_9136.n17 GND 0.48985f
C3493 a_n5004_9136.n18 GND 0.489851f
C3494 a_n5004_9136.n19 GND 0.489851f
C3495 a_n5004_9136.n20 GND 0.489851f
C3496 a_n5004_9136.n21 GND 0.489851f
C3497 a_n5004_9136.n22 GND 0.489851f
C3498 a_n5004_9136.n23 GND 1.29857f
C3499 a_n5004_9136.n24 GND 2.62277f
C3500 a_n5004_9136.n25 GND 2.54785f
C3501 a_n5004_9136.n26 GND 4.53977f
C3502 a_n5004_9136.n27 GND 0.142621f
C3503 a_n5004_9136.n28 GND 0.142621f
C3504 a_n5004_9136.n29 GND 0.142621f
C3505 a_n5004_9136.n30 GND 0.142621f
C3506 a_n5004_9136.n31 GND 0.142621f
C3507 a_n5004_9136.n32 GND 0.142621f
C3508 a_n5004_9136.n33 GND 0.142621f
C3509 a_n5004_9136.n34 GND 0.142621f
C3510 a_n5004_9136.n35 GND 0.498347f
C3511 a_n5004_9136.n36 GND 0.131227f
C3512 a_n5004_9136.t5 GND 0.050415f
C3513 a_n5004_9136.t28 GND 1.33325f
C3514 a_n5004_9136.t29 GND 1.0535f
C3515 a_n5004_9136.n37 GND 0.624399f
C3516 a_n5004_9136.t25 GND 1.0535f
C3517 a_n5004_9136.t44 GND 1.33325f
C3518 a_n5004_9136.t17 GND 0.403223f
C3519 a_n5004_9136.t7 GND 0.051758f
C3520 a_n5004_9136.t11 GND 0.051758f
C3521 a_n5004_9136.n38 GND 0.283404f
C3522 a_n5004_9136.t15 GND 0.397541f
C3523 a_n5004_9136.t30 GND 1.33325f
C3524 a_n5004_9136.t34 GND 1.0535f
C3525 a_n5004_9136.n39 GND 0.624397f
C3526 a_n5004_9136.t31 GND 1.0535f
C3527 a_n5004_9136.t36 GND 1.33325f
C3528 a_n5004_9136.t42 GND 1.28259f
C3529 a_n5004_9136.t40 GND 1.0535f
C3530 a_n5004_9136.n40 GND 0.535331f
C3531 a_n5004_9136.t45 GND 1.0535f
C3532 a_n5004_9136.t33 GND 1.33325f
C3533 a_n5004_9136.t26 GND 1.33325f
C3534 a_n5004_9136.t43 GND 1.0535f
C3535 a_n5004_9136.n41 GND 0.624397f
C3536 a_n5004_9136.t37 GND 1.0535f
C3537 a_n5004_9136.t35 GND 1.33325f
C3538 a_n5004_9136.t27 GND 1.33325f
C3539 a_n5004_9136.t23 GND 1.0535f
C3540 a_n5004_9136.n42 GND 0.624397f
C3541 a_n5004_9136.t41 GND 1.0535f
C3542 a_n5004_9136.t38 GND 1.33325f
C3543 a_n5004_9136.t32 GND 1.33325f
C3544 a_n5004_9136.t39 GND 1.0535f
C3545 a_n5004_9136.n43 GND 0.624399f
C3546 a_n5004_9136.t24 GND 1.0535f
C3547 a_n5004_9136.t22 GND 1.33325f
C3548 a_n5004_9136.t16 GND 1.33325f
C3549 a_n5004_9136.t6 GND 1.0535f
C3550 a_n5004_9136.n44 GND 0.624399f
C3551 a_n5004_9136.t10 GND 1.0535f
C3552 a_n5004_9136.t14 GND 1.33325f
C3553 a_n5004_9136.n45 GND 0.624397f
C3554 a_n5004_9136.n46 GND 0.624397f
C3555 a_n5004_9136.t20 GND 1.33325f
C3556 a_n5004_9136.t18 GND 1.0535f
C3557 a_n5004_9136.n47 GND 0.624399f
C3558 a_n5004_9136.t12 GND 1.0535f
C3559 a_n5004_9136.t8 GND 1.33325f
C3560 a_n5004_9136.n48 GND 0.624397f
C3561 a_n5004_9136.t9 GND 0.403223f
C3562 a_n5004_9136.t19 GND 0.051758f
C3563 a_n5004_9136.t13 GND 0.051758f
C3564 a_n5004_9136.n49 GND 0.283404f
C3565 a_n5004_9136.t21 GND 0.397542f
C3566 a_n5004_9136.n50 GND 0.624399f
C3567 a_n5004_9136.n51 GND 0.624399f
C3568 a_n5004_9136.n52 GND 0.624399f
C3569 a_n5004_9136.n53 GND 0.624399f
C3570 a_n5004_9136.n54 GND 0.624397f
C3571 a_n5004_9136.t3 GND 0.539141f
C3572 a_n5004_9136.t2 GND 0.050415f
C3573 a_n5004_9136.t4 GND 0.050415f
C3574 a_n5004_9136.n55 GND 0.426746f
C3575 a_n5004_9136.n56 GND 2.21146f
C3576 a_n5004_9136.t1 GND 0.536359f
C3577 a_n5004_9136.n57 GND 0.426747f
C3578 a_n5004_9136.t0 GND 0.050415f
.ends

