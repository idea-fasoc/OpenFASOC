* NGSPICE file created from diff_pair_sample_0600.ext - technology: sky130A

.subckt diff_pair_sample_0600 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t18 B.t0 sky130_fd_pr__nfet_01v8 ad=0.6666 pd=4.37 as=0.6666 ps=4.37 w=4.04 l=4
X1 VDD2.t8 VN.t1 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5756 pd=8.86 as=0.6666 ps=4.37 w=4.04 l=4
X2 VDD1.t9 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5756 pd=8.86 as=0.6666 ps=4.37 w=4.04 l=4
X3 VTAIL.t14 VN.t2 VDD2.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=0.6666 pd=4.37 as=0.6666 ps=4.37 w=4.04 l=4
X4 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=1.5756 pd=8.86 as=0 ps=0 w=4.04 l=4
X5 VDD2.t6 VN.t3 VTAIL.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=0.6666 pd=4.37 as=0.6666 ps=4.37 w=4.04 l=4
X6 VDD1.t8 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.6666 pd=4.37 as=0.6666 ps=4.37 w=4.04 l=4
X7 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=1.5756 pd=8.86 as=0 ps=0 w=4.04 l=4
X8 VTAIL.t17 VN.t4 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.6666 pd=4.37 as=0.6666 ps=4.37 w=4.04 l=4
X9 VDD2.t4 VN.t5 VTAIL.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=0.6666 pd=4.37 as=1.5756 ps=8.86 w=4.04 l=4
X10 VTAIL.t10 VN.t6 VDD2.t3 B.t8 sky130_fd_pr__nfet_01v8 ad=0.6666 pd=4.37 as=0.6666 ps=4.37 w=4.04 l=4
X11 VTAIL.t9 VN.t7 VDD2.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=0.6666 pd=4.37 as=0.6666 ps=4.37 w=4.04 l=4
X12 VTAIL.t8 VP.t2 VDD1.t7 B.t8 sky130_fd_pr__nfet_01v8 ad=0.6666 pd=4.37 as=0.6666 ps=4.37 w=4.04 l=4
X13 VTAIL.t7 VP.t3 VDD1.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=0.6666 pd=4.37 as=0.6666 ps=4.37 w=4.04 l=4
X14 VDD1.t5 VP.t4 VTAIL.t19 B.t9 sky130_fd_pr__nfet_01v8 ad=0.6666 pd=4.37 as=0.6666 ps=4.37 w=4.04 l=4
X15 VTAIL.t2 VP.t5 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.6666 pd=4.37 as=0.6666 ps=4.37 w=4.04 l=4
X16 VDD2.t1 VN.t8 VTAIL.t15 B.t5 sky130_fd_pr__nfet_01v8 ad=1.5756 pd=8.86 as=0.6666 ps=4.37 w=4.04 l=4
X17 VDD1.t3 VP.t6 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.6666 pd=4.37 as=1.5756 ps=8.86 w=4.04 l=4
X18 VDD1.t2 VP.t7 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.6666 pd=4.37 as=1.5756 ps=8.86 w=4.04 l=4
X19 VDD2.t0 VN.t9 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=0.6666 pd=4.37 as=1.5756 ps=8.86 w=4.04 l=4
X20 VTAIL.t6 VP.t8 VDD1.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=0.6666 pd=4.37 as=0.6666 ps=4.37 w=4.04 l=4
X21 VDD1.t0 VP.t9 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.5756 pd=8.86 as=0.6666 ps=4.37 w=4.04 l=4
X22 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=1.5756 pd=8.86 as=0 ps=0 w=4.04 l=4
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.5756 pd=8.86 as=0 ps=0 w=4.04 l=4
R0 VN.n113 VN.n58 161.3
R1 VN.n112 VN.n111 161.3
R2 VN.n110 VN.n59 161.3
R3 VN.n109 VN.n108 161.3
R4 VN.n107 VN.n60 161.3
R5 VN.n106 VN.n105 161.3
R6 VN.n104 VN.n61 161.3
R7 VN.n103 VN.n102 161.3
R8 VN.n100 VN.n62 161.3
R9 VN.n99 VN.n98 161.3
R10 VN.n97 VN.n63 161.3
R11 VN.n96 VN.n95 161.3
R12 VN.n94 VN.n64 161.3
R13 VN.n93 VN.n92 161.3
R14 VN.n91 VN.n65 161.3
R15 VN.n90 VN.n89 161.3
R16 VN.n88 VN.n66 161.3
R17 VN.n86 VN.n85 161.3
R18 VN.n84 VN.n67 161.3
R19 VN.n83 VN.n82 161.3
R20 VN.n81 VN.n68 161.3
R21 VN.n80 VN.n79 161.3
R22 VN.n78 VN.n69 161.3
R23 VN.n77 VN.n76 161.3
R24 VN.n75 VN.n70 161.3
R25 VN.n74 VN.n73 161.3
R26 VN.n55 VN.n0 161.3
R27 VN.n54 VN.n53 161.3
R28 VN.n52 VN.n1 161.3
R29 VN.n51 VN.n50 161.3
R30 VN.n49 VN.n2 161.3
R31 VN.n48 VN.n47 161.3
R32 VN.n46 VN.n3 161.3
R33 VN.n45 VN.n44 161.3
R34 VN.n42 VN.n4 161.3
R35 VN.n41 VN.n40 161.3
R36 VN.n39 VN.n5 161.3
R37 VN.n38 VN.n37 161.3
R38 VN.n36 VN.n6 161.3
R39 VN.n35 VN.n34 161.3
R40 VN.n33 VN.n7 161.3
R41 VN.n32 VN.n31 161.3
R42 VN.n30 VN.n8 161.3
R43 VN.n28 VN.n27 161.3
R44 VN.n26 VN.n9 161.3
R45 VN.n25 VN.n24 161.3
R46 VN.n23 VN.n10 161.3
R47 VN.n22 VN.n21 161.3
R48 VN.n20 VN.n11 161.3
R49 VN.n19 VN.n18 161.3
R50 VN.n17 VN.n12 161.3
R51 VN.n16 VN.n15 161.3
R52 VN.n14 VN.n13 71.3575
R53 VN.n72 VN.n71 71.3575
R54 VN.n57 VN.n56 62.2146
R55 VN.n115 VN.n114 62.2146
R56 VN.n14 VN.t1 56.6923
R57 VN.n72 VN.t9 56.6923
R58 VN.n50 VN.n49 56.5617
R59 VN.n108 VN.n107 56.5617
R60 VN VN.n115 54.9779
R61 VN.n23 VN.n22 48.8116
R62 VN.n36 VN.n35 48.8116
R63 VN.n81 VN.n80 48.8116
R64 VN.n94 VN.n93 48.8116
R65 VN.n22 VN.n11 32.3425
R66 VN.n37 VN.n36 32.3425
R67 VN.n80 VN.n69 32.3425
R68 VN.n95 VN.n94 32.3425
R69 VN.n17 VN.n16 24.5923
R70 VN.n18 VN.n17 24.5923
R71 VN.n18 VN.n11 24.5923
R72 VN.n24 VN.n23 24.5923
R73 VN.n24 VN.n9 24.5923
R74 VN.n28 VN.n9 24.5923
R75 VN.n31 VN.n30 24.5923
R76 VN.n31 VN.n7 24.5923
R77 VN.n35 VN.n7 24.5923
R78 VN.n37 VN.n5 24.5923
R79 VN.n41 VN.n5 24.5923
R80 VN.n42 VN.n41 24.5923
R81 VN.n44 VN.n3 24.5923
R82 VN.n48 VN.n3 24.5923
R83 VN.n49 VN.n48 24.5923
R84 VN.n50 VN.n1 24.5923
R85 VN.n54 VN.n1 24.5923
R86 VN.n55 VN.n54 24.5923
R87 VN.n76 VN.n69 24.5923
R88 VN.n76 VN.n75 24.5923
R89 VN.n75 VN.n74 24.5923
R90 VN.n93 VN.n65 24.5923
R91 VN.n89 VN.n65 24.5923
R92 VN.n89 VN.n88 24.5923
R93 VN.n86 VN.n67 24.5923
R94 VN.n82 VN.n67 24.5923
R95 VN.n82 VN.n81 24.5923
R96 VN.n107 VN.n106 24.5923
R97 VN.n106 VN.n61 24.5923
R98 VN.n102 VN.n61 24.5923
R99 VN.n100 VN.n99 24.5923
R100 VN.n99 VN.n63 24.5923
R101 VN.n95 VN.n63 24.5923
R102 VN.n113 VN.n112 24.5923
R103 VN.n112 VN.n59 24.5923
R104 VN.n108 VN.n59 24.5923
R105 VN.n13 VN.t7 24.3415
R106 VN.n29 VN.t0 24.3415
R107 VN.n43 VN.t6 24.3415
R108 VN.n56 VN.t5 24.3415
R109 VN.n71 VN.t2 24.3415
R110 VN.n87 VN.t3 24.3415
R111 VN.n101 VN.t4 24.3415
R112 VN.n114 VN.t8 24.3415
R113 VN.n44 VN.n43 20.6576
R114 VN.n102 VN.n101 20.6576
R115 VN.n56 VN.n55 20.1658
R116 VN.n114 VN.n113 20.1658
R117 VN.n29 VN.n28 12.2964
R118 VN.n30 VN.n29 12.2964
R119 VN.n88 VN.n87 12.2964
R120 VN.n87 VN.n86 12.2964
R121 VN.n16 VN.n13 3.93519
R122 VN.n43 VN.n42 3.93519
R123 VN.n74 VN.n71 3.93519
R124 VN.n101 VN.n100 3.93519
R125 VN.n73 VN.n72 2.6805
R126 VN.n15 VN.n14 2.6805
R127 VN.n115 VN.n58 0.417304
R128 VN.n57 VN.n0 0.417304
R129 VN VN.n57 0.394524
R130 VN.n111 VN.n58 0.189894
R131 VN.n111 VN.n110 0.189894
R132 VN.n110 VN.n109 0.189894
R133 VN.n109 VN.n60 0.189894
R134 VN.n105 VN.n60 0.189894
R135 VN.n105 VN.n104 0.189894
R136 VN.n104 VN.n103 0.189894
R137 VN.n103 VN.n62 0.189894
R138 VN.n98 VN.n62 0.189894
R139 VN.n98 VN.n97 0.189894
R140 VN.n97 VN.n96 0.189894
R141 VN.n96 VN.n64 0.189894
R142 VN.n92 VN.n64 0.189894
R143 VN.n92 VN.n91 0.189894
R144 VN.n91 VN.n90 0.189894
R145 VN.n90 VN.n66 0.189894
R146 VN.n85 VN.n66 0.189894
R147 VN.n85 VN.n84 0.189894
R148 VN.n84 VN.n83 0.189894
R149 VN.n83 VN.n68 0.189894
R150 VN.n79 VN.n68 0.189894
R151 VN.n79 VN.n78 0.189894
R152 VN.n78 VN.n77 0.189894
R153 VN.n77 VN.n70 0.189894
R154 VN.n73 VN.n70 0.189894
R155 VN.n15 VN.n12 0.189894
R156 VN.n19 VN.n12 0.189894
R157 VN.n20 VN.n19 0.189894
R158 VN.n21 VN.n20 0.189894
R159 VN.n21 VN.n10 0.189894
R160 VN.n25 VN.n10 0.189894
R161 VN.n26 VN.n25 0.189894
R162 VN.n27 VN.n26 0.189894
R163 VN.n27 VN.n8 0.189894
R164 VN.n32 VN.n8 0.189894
R165 VN.n33 VN.n32 0.189894
R166 VN.n34 VN.n33 0.189894
R167 VN.n34 VN.n6 0.189894
R168 VN.n38 VN.n6 0.189894
R169 VN.n39 VN.n38 0.189894
R170 VN.n40 VN.n39 0.189894
R171 VN.n40 VN.n4 0.189894
R172 VN.n45 VN.n4 0.189894
R173 VN.n46 VN.n45 0.189894
R174 VN.n47 VN.n46 0.189894
R175 VN.n47 VN.n2 0.189894
R176 VN.n51 VN.n2 0.189894
R177 VN.n52 VN.n51 0.189894
R178 VN.n53 VN.n52 0.189894
R179 VN.n53 VN.n0 0.189894
R180 VTAIL.n88 VTAIL.n74 289.615
R181 VTAIL.n16 VTAIL.n2 289.615
R182 VTAIL.n68 VTAIL.n54 289.615
R183 VTAIL.n44 VTAIL.n30 289.615
R184 VTAIL.n81 VTAIL.n80 185
R185 VTAIL.n78 VTAIL.n77 185
R186 VTAIL.n87 VTAIL.n86 185
R187 VTAIL.n89 VTAIL.n88 185
R188 VTAIL.n9 VTAIL.n8 185
R189 VTAIL.n6 VTAIL.n5 185
R190 VTAIL.n15 VTAIL.n14 185
R191 VTAIL.n17 VTAIL.n16 185
R192 VTAIL.n69 VTAIL.n68 185
R193 VTAIL.n67 VTAIL.n66 185
R194 VTAIL.n58 VTAIL.n57 185
R195 VTAIL.n61 VTAIL.n60 185
R196 VTAIL.n45 VTAIL.n44 185
R197 VTAIL.n43 VTAIL.n42 185
R198 VTAIL.n34 VTAIL.n33 185
R199 VTAIL.n37 VTAIL.n36 185
R200 VTAIL.t12 VTAIL.n79 147.888
R201 VTAIL.t4 VTAIL.n7 147.888
R202 VTAIL.t1 VTAIL.n59 147.888
R203 VTAIL.t11 VTAIL.n35 147.888
R204 VTAIL.n80 VTAIL.n77 104.615
R205 VTAIL.n87 VTAIL.n77 104.615
R206 VTAIL.n88 VTAIL.n87 104.615
R207 VTAIL.n8 VTAIL.n5 104.615
R208 VTAIL.n15 VTAIL.n5 104.615
R209 VTAIL.n16 VTAIL.n15 104.615
R210 VTAIL.n68 VTAIL.n67 104.615
R211 VTAIL.n67 VTAIL.n57 104.615
R212 VTAIL.n60 VTAIL.n57 104.615
R213 VTAIL.n44 VTAIL.n43 104.615
R214 VTAIL.n43 VTAIL.n33 104.615
R215 VTAIL.n36 VTAIL.n33 104.615
R216 VTAIL.n53 VTAIL.n52 60.6641
R217 VTAIL.n51 VTAIL.n50 60.6641
R218 VTAIL.n29 VTAIL.n28 60.6641
R219 VTAIL.n27 VTAIL.n26 60.6641
R220 VTAIL.n95 VTAIL.n94 60.664
R221 VTAIL.n1 VTAIL.n0 60.664
R222 VTAIL.n23 VTAIL.n22 60.664
R223 VTAIL.n25 VTAIL.n24 60.664
R224 VTAIL.n80 VTAIL.t12 52.3082
R225 VTAIL.n8 VTAIL.t4 52.3082
R226 VTAIL.n60 VTAIL.t1 52.3082
R227 VTAIL.n36 VTAIL.t11 52.3082
R228 VTAIL.n93 VTAIL.n92 36.0641
R229 VTAIL.n21 VTAIL.n20 36.0641
R230 VTAIL.n73 VTAIL.n72 36.0641
R231 VTAIL.n49 VTAIL.n48 36.0641
R232 VTAIL.n27 VTAIL.n25 23.3152
R233 VTAIL.n93 VTAIL.n73 19.5824
R234 VTAIL.n81 VTAIL.n79 15.6496
R235 VTAIL.n9 VTAIL.n7 15.6496
R236 VTAIL.n61 VTAIL.n59 15.6496
R237 VTAIL.n37 VTAIL.n35 15.6496
R238 VTAIL.n82 VTAIL.n78 12.8005
R239 VTAIL.n10 VTAIL.n6 12.8005
R240 VTAIL.n62 VTAIL.n58 12.8005
R241 VTAIL.n38 VTAIL.n34 12.8005
R242 VTAIL.n86 VTAIL.n85 12.0247
R243 VTAIL.n14 VTAIL.n13 12.0247
R244 VTAIL.n66 VTAIL.n65 12.0247
R245 VTAIL.n42 VTAIL.n41 12.0247
R246 VTAIL.n89 VTAIL.n76 11.249
R247 VTAIL.n17 VTAIL.n4 11.249
R248 VTAIL.n69 VTAIL.n56 11.249
R249 VTAIL.n45 VTAIL.n32 11.249
R250 VTAIL.n90 VTAIL.n74 10.4732
R251 VTAIL.n18 VTAIL.n2 10.4732
R252 VTAIL.n70 VTAIL.n54 10.4732
R253 VTAIL.n46 VTAIL.n30 10.4732
R254 VTAIL.n92 VTAIL.n91 9.45567
R255 VTAIL.n20 VTAIL.n19 9.45567
R256 VTAIL.n72 VTAIL.n71 9.45567
R257 VTAIL.n48 VTAIL.n47 9.45567
R258 VTAIL.n91 VTAIL.n90 9.3005
R259 VTAIL.n76 VTAIL.n75 9.3005
R260 VTAIL.n85 VTAIL.n84 9.3005
R261 VTAIL.n83 VTAIL.n82 9.3005
R262 VTAIL.n19 VTAIL.n18 9.3005
R263 VTAIL.n4 VTAIL.n3 9.3005
R264 VTAIL.n13 VTAIL.n12 9.3005
R265 VTAIL.n11 VTAIL.n10 9.3005
R266 VTAIL.n71 VTAIL.n70 9.3005
R267 VTAIL.n56 VTAIL.n55 9.3005
R268 VTAIL.n65 VTAIL.n64 9.3005
R269 VTAIL.n63 VTAIL.n62 9.3005
R270 VTAIL.n47 VTAIL.n46 9.3005
R271 VTAIL.n32 VTAIL.n31 9.3005
R272 VTAIL.n41 VTAIL.n40 9.3005
R273 VTAIL.n39 VTAIL.n38 9.3005
R274 VTAIL.n94 VTAIL.t18 4.90149
R275 VTAIL.n94 VTAIL.t10 4.90149
R276 VTAIL.n0 VTAIL.t13 4.90149
R277 VTAIL.n0 VTAIL.t9 4.90149
R278 VTAIL.n22 VTAIL.t19 4.90149
R279 VTAIL.n22 VTAIL.t6 4.90149
R280 VTAIL.n24 VTAIL.t5 4.90149
R281 VTAIL.n24 VTAIL.t2 4.90149
R282 VTAIL.n52 VTAIL.t0 4.90149
R283 VTAIL.n52 VTAIL.t8 4.90149
R284 VTAIL.n50 VTAIL.t3 4.90149
R285 VTAIL.n50 VTAIL.t7 4.90149
R286 VTAIL.n28 VTAIL.t16 4.90149
R287 VTAIL.n28 VTAIL.t14 4.90149
R288 VTAIL.n26 VTAIL.t15 4.90149
R289 VTAIL.n26 VTAIL.t17 4.90149
R290 VTAIL.n83 VTAIL.n79 4.40546
R291 VTAIL.n11 VTAIL.n7 4.40546
R292 VTAIL.n63 VTAIL.n59 4.40546
R293 VTAIL.n39 VTAIL.n35 4.40546
R294 VTAIL.n29 VTAIL.n27 3.73326
R295 VTAIL.n49 VTAIL.n29 3.73326
R296 VTAIL.n53 VTAIL.n51 3.73326
R297 VTAIL.n73 VTAIL.n53 3.73326
R298 VTAIL.n25 VTAIL.n23 3.73326
R299 VTAIL.n23 VTAIL.n21 3.73326
R300 VTAIL.n95 VTAIL.n93 3.73326
R301 VTAIL.n92 VTAIL.n74 3.49141
R302 VTAIL.n20 VTAIL.n2 3.49141
R303 VTAIL.n72 VTAIL.n54 3.49141
R304 VTAIL.n48 VTAIL.n30 3.49141
R305 VTAIL VTAIL.n1 2.85826
R306 VTAIL.n90 VTAIL.n89 2.71565
R307 VTAIL.n18 VTAIL.n17 2.71565
R308 VTAIL.n70 VTAIL.n69 2.71565
R309 VTAIL.n46 VTAIL.n45 2.71565
R310 VTAIL.n51 VTAIL.n49 2.33671
R311 VTAIL.n21 VTAIL.n1 2.33671
R312 VTAIL.n86 VTAIL.n76 1.93989
R313 VTAIL.n14 VTAIL.n4 1.93989
R314 VTAIL.n66 VTAIL.n56 1.93989
R315 VTAIL.n42 VTAIL.n32 1.93989
R316 VTAIL.n85 VTAIL.n78 1.16414
R317 VTAIL.n13 VTAIL.n6 1.16414
R318 VTAIL.n65 VTAIL.n58 1.16414
R319 VTAIL.n41 VTAIL.n34 1.16414
R320 VTAIL VTAIL.n95 0.8755
R321 VTAIL.n82 VTAIL.n81 0.388379
R322 VTAIL.n10 VTAIL.n9 0.388379
R323 VTAIL.n62 VTAIL.n61 0.388379
R324 VTAIL.n38 VTAIL.n37 0.388379
R325 VTAIL.n84 VTAIL.n83 0.155672
R326 VTAIL.n84 VTAIL.n75 0.155672
R327 VTAIL.n91 VTAIL.n75 0.155672
R328 VTAIL.n12 VTAIL.n11 0.155672
R329 VTAIL.n12 VTAIL.n3 0.155672
R330 VTAIL.n19 VTAIL.n3 0.155672
R331 VTAIL.n71 VTAIL.n55 0.155672
R332 VTAIL.n64 VTAIL.n55 0.155672
R333 VTAIL.n64 VTAIL.n63 0.155672
R334 VTAIL.n47 VTAIL.n31 0.155672
R335 VTAIL.n40 VTAIL.n31 0.155672
R336 VTAIL.n40 VTAIL.n39 0.155672
R337 VDD2.n37 VDD2.n23 289.615
R338 VDD2.n14 VDD2.n0 289.615
R339 VDD2.n38 VDD2.n37 185
R340 VDD2.n36 VDD2.n35 185
R341 VDD2.n27 VDD2.n26 185
R342 VDD2.n30 VDD2.n29 185
R343 VDD2.n7 VDD2.n6 185
R344 VDD2.n4 VDD2.n3 185
R345 VDD2.n13 VDD2.n12 185
R346 VDD2.n15 VDD2.n14 185
R347 VDD2.t1 VDD2.n28 147.888
R348 VDD2.t8 VDD2.n5 147.888
R349 VDD2.n37 VDD2.n36 104.615
R350 VDD2.n36 VDD2.n26 104.615
R351 VDD2.n29 VDD2.n26 104.615
R352 VDD2.n6 VDD2.n3 104.615
R353 VDD2.n13 VDD2.n3 104.615
R354 VDD2.n14 VDD2.n13 104.615
R355 VDD2.n22 VDD2.n21 80.087
R356 VDD2 VDD2.n45 80.0841
R357 VDD2.n44 VDD2.n43 77.3429
R358 VDD2.n20 VDD2.n19 77.3428
R359 VDD2.n20 VDD2.n18 56.4757
R360 VDD2.n42 VDD2.n41 52.7429
R361 VDD2.n29 VDD2.t1 52.3082
R362 VDD2.n6 VDD2.t8 52.3082
R363 VDD2.n42 VDD2.n22 44.9287
R364 VDD2.n30 VDD2.n28 15.6496
R365 VDD2.n7 VDD2.n5 15.6496
R366 VDD2.n31 VDD2.n27 12.8005
R367 VDD2.n8 VDD2.n4 12.8005
R368 VDD2.n35 VDD2.n34 12.0247
R369 VDD2.n12 VDD2.n11 12.0247
R370 VDD2.n38 VDD2.n25 11.249
R371 VDD2.n15 VDD2.n2 11.249
R372 VDD2.n39 VDD2.n23 10.4732
R373 VDD2.n16 VDD2.n0 10.4732
R374 VDD2.n41 VDD2.n40 9.45567
R375 VDD2.n18 VDD2.n17 9.45567
R376 VDD2.n40 VDD2.n39 9.3005
R377 VDD2.n25 VDD2.n24 9.3005
R378 VDD2.n34 VDD2.n33 9.3005
R379 VDD2.n32 VDD2.n31 9.3005
R380 VDD2.n17 VDD2.n16 9.3005
R381 VDD2.n2 VDD2.n1 9.3005
R382 VDD2.n11 VDD2.n10 9.3005
R383 VDD2.n9 VDD2.n8 9.3005
R384 VDD2.n45 VDD2.t7 4.90149
R385 VDD2.n45 VDD2.t0 4.90149
R386 VDD2.n43 VDD2.t5 4.90149
R387 VDD2.n43 VDD2.t6 4.90149
R388 VDD2.n21 VDD2.t3 4.90149
R389 VDD2.n21 VDD2.t4 4.90149
R390 VDD2.n19 VDD2.t2 4.90149
R391 VDD2.n19 VDD2.t9 4.90149
R392 VDD2.n32 VDD2.n28 4.40546
R393 VDD2.n9 VDD2.n5 4.40546
R394 VDD2.n44 VDD2.n42 3.73326
R395 VDD2.n41 VDD2.n23 3.49141
R396 VDD2.n18 VDD2.n0 3.49141
R397 VDD2.n39 VDD2.n38 2.71565
R398 VDD2.n16 VDD2.n15 2.71565
R399 VDD2.n35 VDD2.n25 1.93989
R400 VDD2.n12 VDD2.n2 1.93989
R401 VDD2.n34 VDD2.n27 1.16414
R402 VDD2.n11 VDD2.n4 1.16414
R403 VDD2 VDD2.n44 0.991879
R404 VDD2.n22 VDD2.n20 0.878344
R405 VDD2.n31 VDD2.n30 0.388379
R406 VDD2.n8 VDD2.n7 0.388379
R407 VDD2.n40 VDD2.n24 0.155672
R408 VDD2.n33 VDD2.n24 0.155672
R409 VDD2.n33 VDD2.n32 0.155672
R410 VDD2.n10 VDD2.n9 0.155672
R411 VDD2.n10 VDD2.n1 0.155672
R412 VDD2.n17 VDD2.n1 0.155672
R413 B.n917 B.n916 585
R414 B.n269 B.n176 585
R415 B.n268 B.n267 585
R416 B.n266 B.n265 585
R417 B.n264 B.n263 585
R418 B.n262 B.n261 585
R419 B.n260 B.n259 585
R420 B.n258 B.n257 585
R421 B.n256 B.n255 585
R422 B.n254 B.n253 585
R423 B.n252 B.n251 585
R424 B.n250 B.n249 585
R425 B.n248 B.n247 585
R426 B.n246 B.n245 585
R427 B.n244 B.n243 585
R428 B.n242 B.n241 585
R429 B.n240 B.n239 585
R430 B.n238 B.n237 585
R431 B.n236 B.n235 585
R432 B.n234 B.n233 585
R433 B.n232 B.n231 585
R434 B.n230 B.n229 585
R435 B.n228 B.n227 585
R436 B.n226 B.n225 585
R437 B.n224 B.n223 585
R438 B.n222 B.n221 585
R439 B.n220 B.n219 585
R440 B.n218 B.n217 585
R441 B.n216 B.n215 585
R442 B.n214 B.n213 585
R443 B.n212 B.n211 585
R444 B.n210 B.n209 585
R445 B.n208 B.n207 585
R446 B.n206 B.n205 585
R447 B.n204 B.n203 585
R448 B.n202 B.n201 585
R449 B.n200 B.n199 585
R450 B.n198 B.n197 585
R451 B.n196 B.n195 585
R452 B.n194 B.n193 585
R453 B.n192 B.n191 585
R454 B.n190 B.n189 585
R455 B.n188 B.n187 585
R456 B.n186 B.n185 585
R457 B.n184 B.n183 585
R458 B.n152 B.n151 585
R459 B.n915 B.n153 585
R460 B.n920 B.n153 585
R461 B.n914 B.n913 585
R462 B.n913 B.n149 585
R463 B.n912 B.n148 585
R464 B.n926 B.n148 585
R465 B.n911 B.n147 585
R466 B.n927 B.n147 585
R467 B.n910 B.n146 585
R468 B.n928 B.n146 585
R469 B.n909 B.n908 585
R470 B.n908 B.n142 585
R471 B.n907 B.n141 585
R472 B.n934 B.n141 585
R473 B.n906 B.n140 585
R474 B.n935 B.n140 585
R475 B.n905 B.n139 585
R476 B.n936 B.n139 585
R477 B.n904 B.n903 585
R478 B.n903 B.n138 585
R479 B.n902 B.n134 585
R480 B.n942 B.n134 585
R481 B.n901 B.n133 585
R482 B.n943 B.n133 585
R483 B.n900 B.n132 585
R484 B.n944 B.n132 585
R485 B.n899 B.n898 585
R486 B.n898 B.n128 585
R487 B.n897 B.n127 585
R488 B.n950 B.n127 585
R489 B.n896 B.n126 585
R490 B.n951 B.n126 585
R491 B.n895 B.n125 585
R492 B.n952 B.n125 585
R493 B.n894 B.n893 585
R494 B.n893 B.n121 585
R495 B.n892 B.n120 585
R496 B.n958 B.n120 585
R497 B.n891 B.n119 585
R498 B.n959 B.n119 585
R499 B.n890 B.n118 585
R500 B.n960 B.n118 585
R501 B.n889 B.n888 585
R502 B.n888 B.n114 585
R503 B.n887 B.n113 585
R504 B.n966 B.n113 585
R505 B.n886 B.n112 585
R506 B.n967 B.n112 585
R507 B.n885 B.n111 585
R508 B.n968 B.n111 585
R509 B.n884 B.n883 585
R510 B.n883 B.n110 585
R511 B.n882 B.n106 585
R512 B.n974 B.n106 585
R513 B.n881 B.n105 585
R514 B.n975 B.n105 585
R515 B.n880 B.n104 585
R516 B.n976 B.n104 585
R517 B.n879 B.n878 585
R518 B.n878 B.n100 585
R519 B.n877 B.n99 585
R520 B.n982 B.n99 585
R521 B.n876 B.n98 585
R522 B.n983 B.n98 585
R523 B.n875 B.n97 585
R524 B.n984 B.n97 585
R525 B.n874 B.n873 585
R526 B.n873 B.n93 585
R527 B.n872 B.n92 585
R528 B.n990 B.n92 585
R529 B.n871 B.n91 585
R530 B.n991 B.n91 585
R531 B.n870 B.n90 585
R532 B.n992 B.n90 585
R533 B.n869 B.n868 585
R534 B.n868 B.n86 585
R535 B.n867 B.n85 585
R536 B.n998 B.n85 585
R537 B.n866 B.n84 585
R538 B.n999 B.n84 585
R539 B.n865 B.n83 585
R540 B.n1000 B.n83 585
R541 B.n864 B.n863 585
R542 B.n863 B.n79 585
R543 B.n862 B.n78 585
R544 B.n1006 B.n78 585
R545 B.n861 B.n77 585
R546 B.n1007 B.n77 585
R547 B.n860 B.n76 585
R548 B.n1008 B.n76 585
R549 B.n859 B.n858 585
R550 B.n858 B.n72 585
R551 B.n857 B.n71 585
R552 B.n1014 B.n71 585
R553 B.n856 B.n70 585
R554 B.n1015 B.n70 585
R555 B.n855 B.n69 585
R556 B.n1016 B.n69 585
R557 B.n854 B.n853 585
R558 B.n853 B.n65 585
R559 B.n852 B.n64 585
R560 B.n1022 B.n64 585
R561 B.n851 B.n63 585
R562 B.n1023 B.n63 585
R563 B.n850 B.n62 585
R564 B.n1024 B.n62 585
R565 B.n849 B.n848 585
R566 B.n848 B.n58 585
R567 B.n847 B.n57 585
R568 B.n1030 B.n57 585
R569 B.n846 B.n56 585
R570 B.n1031 B.n56 585
R571 B.n845 B.n55 585
R572 B.n1032 B.n55 585
R573 B.n844 B.n843 585
R574 B.n843 B.n51 585
R575 B.n842 B.n50 585
R576 B.n1038 B.n50 585
R577 B.n841 B.n49 585
R578 B.n1039 B.n49 585
R579 B.n840 B.n48 585
R580 B.n1040 B.n48 585
R581 B.n839 B.n838 585
R582 B.n838 B.n44 585
R583 B.n837 B.n43 585
R584 B.n1046 B.n43 585
R585 B.n836 B.n42 585
R586 B.n1047 B.n42 585
R587 B.n835 B.n41 585
R588 B.n1048 B.n41 585
R589 B.n834 B.n833 585
R590 B.n833 B.n37 585
R591 B.n832 B.n36 585
R592 B.n1054 B.n36 585
R593 B.n831 B.n35 585
R594 B.n1055 B.n35 585
R595 B.n830 B.n34 585
R596 B.n1056 B.n34 585
R597 B.n829 B.n828 585
R598 B.n828 B.n30 585
R599 B.n827 B.n29 585
R600 B.n1062 B.n29 585
R601 B.n826 B.n28 585
R602 B.n1063 B.n28 585
R603 B.n825 B.n27 585
R604 B.n1064 B.n27 585
R605 B.n824 B.n823 585
R606 B.n823 B.n23 585
R607 B.n822 B.n22 585
R608 B.n1070 B.n22 585
R609 B.n821 B.n21 585
R610 B.n1071 B.n21 585
R611 B.n820 B.n20 585
R612 B.n1072 B.n20 585
R613 B.n819 B.n818 585
R614 B.n818 B.n16 585
R615 B.n817 B.n15 585
R616 B.n1078 B.n15 585
R617 B.n816 B.n14 585
R618 B.n1079 B.n14 585
R619 B.n815 B.n13 585
R620 B.n1080 B.n13 585
R621 B.n814 B.n813 585
R622 B.n813 B.n12 585
R623 B.n812 B.n811 585
R624 B.n812 B.n8 585
R625 B.n810 B.n7 585
R626 B.n1087 B.n7 585
R627 B.n809 B.n6 585
R628 B.n1088 B.n6 585
R629 B.n808 B.n5 585
R630 B.n1089 B.n5 585
R631 B.n807 B.n806 585
R632 B.n806 B.n4 585
R633 B.n805 B.n270 585
R634 B.n805 B.n804 585
R635 B.n795 B.n271 585
R636 B.n272 B.n271 585
R637 B.n797 B.n796 585
R638 B.n798 B.n797 585
R639 B.n794 B.n277 585
R640 B.n277 B.n276 585
R641 B.n793 B.n792 585
R642 B.n792 B.n791 585
R643 B.n279 B.n278 585
R644 B.n280 B.n279 585
R645 B.n784 B.n783 585
R646 B.n785 B.n784 585
R647 B.n782 B.n285 585
R648 B.n285 B.n284 585
R649 B.n781 B.n780 585
R650 B.n780 B.n779 585
R651 B.n287 B.n286 585
R652 B.n288 B.n287 585
R653 B.n772 B.n771 585
R654 B.n773 B.n772 585
R655 B.n770 B.n293 585
R656 B.n293 B.n292 585
R657 B.n769 B.n768 585
R658 B.n768 B.n767 585
R659 B.n295 B.n294 585
R660 B.n296 B.n295 585
R661 B.n760 B.n759 585
R662 B.n761 B.n760 585
R663 B.n758 B.n301 585
R664 B.n301 B.n300 585
R665 B.n757 B.n756 585
R666 B.n756 B.n755 585
R667 B.n303 B.n302 585
R668 B.n304 B.n303 585
R669 B.n748 B.n747 585
R670 B.n749 B.n748 585
R671 B.n746 B.n308 585
R672 B.n312 B.n308 585
R673 B.n745 B.n744 585
R674 B.n744 B.n743 585
R675 B.n310 B.n309 585
R676 B.n311 B.n310 585
R677 B.n736 B.n735 585
R678 B.n737 B.n736 585
R679 B.n734 B.n317 585
R680 B.n317 B.n316 585
R681 B.n733 B.n732 585
R682 B.n732 B.n731 585
R683 B.n319 B.n318 585
R684 B.n320 B.n319 585
R685 B.n724 B.n723 585
R686 B.n725 B.n724 585
R687 B.n722 B.n325 585
R688 B.n325 B.n324 585
R689 B.n721 B.n720 585
R690 B.n720 B.n719 585
R691 B.n327 B.n326 585
R692 B.n328 B.n327 585
R693 B.n712 B.n711 585
R694 B.n713 B.n712 585
R695 B.n710 B.n332 585
R696 B.n336 B.n332 585
R697 B.n709 B.n708 585
R698 B.n708 B.n707 585
R699 B.n334 B.n333 585
R700 B.n335 B.n334 585
R701 B.n700 B.n699 585
R702 B.n701 B.n700 585
R703 B.n698 B.n341 585
R704 B.n341 B.n340 585
R705 B.n697 B.n696 585
R706 B.n696 B.n695 585
R707 B.n343 B.n342 585
R708 B.n344 B.n343 585
R709 B.n688 B.n687 585
R710 B.n689 B.n688 585
R711 B.n686 B.n349 585
R712 B.n349 B.n348 585
R713 B.n685 B.n684 585
R714 B.n684 B.n683 585
R715 B.n351 B.n350 585
R716 B.n352 B.n351 585
R717 B.n676 B.n675 585
R718 B.n677 B.n676 585
R719 B.n674 B.n357 585
R720 B.n357 B.n356 585
R721 B.n673 B.n672 585
R722 B.n672 B.n671 585
R723 B.n359 B.n358 585
R724 B.n360 B.n359 585
R725 B.n664 B.n663 585
R726 B.n665 B.n664 585
R727 B.n662 B.n365 585
R728 B.n365 B.n364 585
R729 B.n661 B.n660 585
R730 B.n660 B.n659 585
R731 B.n367 B.n366 585
R732 B.n368 B.n367 585
R733 B.n652 B.n651 585
R734 B.n653 B.n652 585
R735 B.n650 B.n373 585
R736 B.n373 B.n372 585
R737 B.n649 B.n648 585
R738 B.n648 B.n647 585
R739 B.n375 B.n374 585
R740 B.n376 B.n375 585
R741 B.n640 B.n639 585
R742 B.n641 B.n640 585
R743 B.n638 B.n381 585
R744 B.n381 B.n380 585
R745 B.n637 B.n636 585
R746 B.n636 B.n635 585
R747 B.n383 B.n382 585
R748 B.n628 B.n383 585
R749 B.n627 B.n626 585
R750 B.n629 B.n627 585
R751 B.n625 B.n388 585
R752 B.n388 B.n387 585
R753 B.n624 B.n623 585
R754 B.n623 B.n622 585
R755 B.n390 B.n389 585
R756 B.n391 B.n390 585
R757 B.n615 B.n614 585
R758 B.n616 B.n615 585
R759 B.n613 B.n396 585
R760 B.n396 B.n395 585
R761 B.n612 B.n611 585
R762 B.n611 B.n610 585
R763 B.n398 B.n397 585
R764 B.n399 B.n398 585
R765 B.n603 B.n602 585
R766 B.n604 B.n603 585
R767 B.n601 B.n404 585
R768 B.n404 B.n403 585
R769 B.n600 B.n599 585
R770 B.n599 B.n598 585
R771 B.n406 B.n405 585
R772 B.n407 B.n406 585
R773 B.n591 B.n590 585
R774 B.n592 B.n591 585
R775 B.n589 B.n412 585
R776 B.n412 B.n411 585
R777 B.n588 B.n587 585
R778 B.n587 B.n586 585
R779 B.n414 B.n413 585
R780 B.n579 B.n414 585
R781 B.n578 B.n577 585
R782 B.n580 B.n578 585
R783 B.n576 B.n419 585
R784 B.n419 B.n418 585
R785 B.n575 B.n574 585
R786 B.n574 B.n573 585
R787 B.n421 B.n420 585
R788 B.n422 B.n421 585
R789 B.n566 B.n565 585
R790 B.n567 B.n566 585
R791 B.n564 B.n427 585
R792 B.n427 B.n426 585
R793 B.n563 B.n562 585
R794 B.n562 B.n561 585
R795 B.n429 B.n428 585
R796 B.n430 B.n429 585
R797 B.n554 B.n553 585
R798 B.n555 B.n554 585
R799 B.n433 B.n432 585
R800 B.n462 B.n460 585
R801 B.n463 B.n459 585
R802 B.n463 B.n434 585
R803 B.n466 B.n465 585
R804 B.n467 B.n458 585
R805 B.n469 B.n468 585
R806 B.n471 B.n457 585
R807 B.n474 B.n473 585
R808 B.n475 B.n456 585
R809 B.n477 B.n476 585
R810 B.n479 B.n455 585
R811 B.n482 B.n481 585
R812 B.n483 B.n454 585
R813 B.n485 B.n484 585
R814 B.n487 B.n453 585
R815 B.n490 B.n489 585
R816 B.n491 B.n452 585
R817 B.n496 B.n495 585
R818 B.n498 B.n451 585
R819 B.n501 B.n500 585
R820 B.n502 B.n450 585
R821 B.n504 B.n503 585
R822 B.n506 B.n449 585
R823 B.n509 B.n508 585
R824 B.n510 B.n448 585
R825 B.n512 B.n511 585
R826 B.n514 B.n447 585
R827 B.n517 B.n516 585
R828 B.n519 B.n444 585
R829 B.n521 B.n520 585
R830 B.n523 B.n443 585
R831 B.n526 B.n525 585
R832 B.n527 B.n442 585
R833 B.n529 B.n528 585
R834 B.n531 B.n441 585
R835 B.n534 B.n533 585
R836 B.n535 B.n440 585
R837 B.n537 B.n536 585
R838 B.n539 B.n439 585
R839 B.n542 B.n541 585
R840 B.n543 B.n438 585
R841 B.n545 B.n544 585
R842 B.n547 B.n437 585
R843 B.n548 B.n436 585
R844 B.n551 B.n550 585
R845 B.n552 B.n435 585
R846 B.n435 B.n434 585
R847 B.n557 B.n556 585
R848 B.n556 B.n555 585
R849 B.n558 B.n431 585
R850 B.n431 B.n430 585
R851 B.n560 B.n559 585
R852 B.n561 B.n560 585
R853 B.n425 B.n424 585
R854 B.n426 B.n425 585
R855 B.n569 B.n568 585
R856 B.n568 B.n567 585
R857 B.n570 B.n423 585
R858 B.n423 B.n422 585
R859 B.n572 B.n571 585
R860 B.n573 B.n572 585
R861 B.n417 B.n416 585
R862 B.n418 B.n417 585
R863 B.n582 B.n581 585
R864 B.n581 B.n580 585
R865 B.n583 B.n415 585
R866 B.n579 B.n415 585
R867 B.n585 B.n584 585
R868 B.n586 B.n585 585
R869 B.n410 B.n409 585
R870 B.n411 B.n410 585
R871 B.n594 B.n593 585
R872 B.n593 B.n592 585
R873 B.n595 B.n408 585
R874 B.n408 B.n407 585
R875 B.n597 B.n596 585
R876 B.n598 B.n597 585
R877 B.n402 B.n401 585
R878 B.n403 B.n402 585
R879 B.n606 B.n605 585
R880 B.n605 B.n604 585
R881 B.n607 B.n400 585
R882 B.n400 B.n399 585
R883 B.n609 B.n608 585
R884 B.n610 B.n609 585
R885 B.n394 B.n393 585
R886 B.n395 B.n394 585
R887 B.n618 B.n617 585
R888 B.n617 B.n616 585
R889 B.n619 B.n392 585
R890 B.n392 B.n391 585
R891 B.n621 B.n620 585
R892 B.n622 B.n621 585
R893 B.n386 B.n385 585
R894 B.n387 B.n386 585
R895 B.n631 B.n630 585
R896 B.n630 B.n629 585
R897 B.n632 B.n384 585
R898 B.n628 B.n384 585
R899 B.n634 B.n633 585
R900 B.n635 B.n634 585
R901 B.n379 B.n378 585
R902 B.n380 B.n379 585
R903 B.n643 B.n642 585
R904 B.n642 B.n641 585
R905 B.n644 B.n377 585
R906 B.n377 B.n376 585
R907 B.n646 B.n645 585
R908 B.n647 B.n646 585
R909 B.n371 B.n370 585
R910 B.n372 B.n371 585
R911 B.n655 B.n654 585
R912 B.n654 B.n653 585
R913 B.n656 B.n369 585
R914 B.n369 B.n368 585
R915 B.n658 B.n657 585
R916 B.n659 B.n658 585
R917 B.n363 B.n362 585
R918 B.n364 B.n363 585
R919 B.n667 B.n666 585
R920 B.n666 B.n665 585
R921 B.n668 B.n361 585
R922 B.n361 B.n360 585
R923 B.n670 B.n669 585
R924 B.n671 B.n670 585
R925 B.n355 B.n354 585
R926 B.n356 B.n355 585
R927 B.n679 B.n678 585
R928 B.n678 B.n677 585
R929 B.n680 B.n353 585
R930 B.n353 B.n352 585
R931 B.n682 B.n681 585
R932 B.n683 B.n682 585
R933 B.n347 B.n346 585
R934 B.n348 B.n347 585
R935 B.n691 B.n690 585
R936 B.n690 B.n689 585
R937 B.n692 B.n345 585
R938 B.n345 B.n344 585
R939 B.n694 B.n693 585
R940 B.n695 B.n694 585
R941 B.n339 B.n338 585
R942 B.n340 B.n339 585
R943 B.n703 B.n702 585
R944 B.n702 B.n701 585
R945 B.n704 B.n337 585
R946 B.n337 B.n335 585
R947 B.n706 B.n705 585
R948 B.n707 B.n706 585
R949 B.n331 B.n330 585
R950 B.n336 B.n331 585
R951 B.n715 B.n714 585
R952 B.n714 B.n713 585
R953 B.n716 B.n329 585
R954 B.n329 B.n328 585
R955 B.n718 B.n717 585
R956 B.n719 B.n718 585
R957 B.n323 B.n322 585
R958 B.n324 B.n323 585
R959 B.n727 B.n726 585
R960 B.n726 B.n725 585
R961 B.n728 B.n321 585
R962 B.n321 B.n320 585
R963 B.n730 B.n729 585
R964 B.n731 B.n730 585
R965 B.n315 B.n314 585
R966 B.n316 B.n315 585
R967 B.n739 B.n738 585
R968 B.n738 B.n737 585
R969 B.n740 B.n313 585
R970 B.n313 B.n311 585
R971 B.n742 B.n741 585
R972 B.n743 B.n742 585
R973 B.n307 B.n306 585
R974 B.n312 B.n307 585
R975 B.n751 B.n750 585
R976 B.n750 B.n749 585
R977 B.n752 B.n305 585
R978 B.n305 B.n304 585
R979 B.n754 B.n753 585
R980 B.n755 B.n754 585
R981 B.n299 B.n298 585
R982 B.n300 B.n299 585
R983 B.n763 B.n762 585
R984 B.n762 B.n761 585
R985 B.n764 B.n297 585
R986 B.n297 B.n296 585
R987 B.n766 B.n765 585
R988 B.n767 B.n766 585
R989 B.n291 B.n290 585
R990 B.n292 B.n291 585
R991 B.n775 B.n774 585
R992 B.n774 B.n773 585
R993 B.n776 B.n289 585
R994 B.n289 B.n288 585
R995 B.n778 B.n777 585
R996 B.n779 B.n778 585
R997 B.n283 B.n282 585
R998 B.n284 B.n283 585
R999 B.n787 B.n786 585
R1000 B.n786 B.n785 585
R1001 B.n788 B.n281 585
R1002 B.n281 B.n280 585
R1003 B.n790 B.n789 585
R1004 B.n791 B.n790 585
R1005 B.n275 B.n274 585
R1006 B.n276 B.n275 585
R1007 B.n800 B.n799 585
R1008 B.n799 B.n798 585
R1009 B.n801 B.n273 585
R1010 B.n273 B.n272 585
R1011 B.n803 B.n802 585
R1012 B.n804 B.n803 585
R1013 B.n3 B.n0 585
R1014 B.n4 B.n3 585
R1015 B.n1086 B.n1 585
R1016 B.n1087 B.n1086 585
R1017 B.n1085 B.n1084 585
R1018 B.n1085 B.n8 585
R1019 B.n1083 B.n9 585
R1020 B.n12 B.n9 585
R1021 B.n1082 B.n1081 585
R1022 B.n1081 B.n1080 585
R1023 B.n11 B.n10 585
R1024 B.n1079 B.n11 585
R1025 B.n1077 B.n1076 585
R1026 B.n1078 B.n1077 585
R1027 B.n1075 B.n17 585
R1028 B.n17 B.n16 585
R1029 B.n1074 B.n1073 585
R1030 B.n1073 B.n1072 585
R1031 B.n19 B.n18 585
R1032 B.n1071 B.n19 585
R1033 B.n1069 B.n1068 585
R1034 B.n1070 B.n1069 585
R1035 B.n1067 B.n24 585
R1036 B.n24 B.n23 585
R1037 B.n1066 B.n1065 585
R1038 B.n1065 B.n1064 585
R1039 B.n26 B.n25 585
R1040 B.n1063 B.n26 585
R1041 B.n1061 B.n1060 585
R1042 B.n1062 B.n1061 585
R1043 B.n1059 B.n31 585
R1044 B.n31 B.n30 585
R1045 B.n1058 B.n1057 585
R1046 B.n1057 B.n1056 585
R1047 B.n33 B.n32 585
R1048 B.n1055 B.n33 585
R1049 B.n1053 B.n1052 585
R1050 B.n1054 B.n1053 585
R1051 B.n1051 B.n38 585
R1052 B.n38 B.n37 585
R1053 B.n1050 B.n1049 585
R1054 B.n1049 B.n1048 585
R1055 B.n40 B.n39 585
R1056 B.n1047 B.n40 585
R1057 B.n1045 B.n1044 585
R1058 B.n1046 B.n1045 585
R1059 B.n1043 B.n45 585
R1060 B.n45 B.n44 585
R1061 B.n1042 B.n1041 585
R1062 B.n1041 B.n1040 585
R1063 B.n47 B.n46 585
R1064 B.n1039 B.n47 585
R1065 B.n1037 B.n1036 585
R1066 B.n1038 B.n1037 585
R1067 B.n1035 B.n52 585
R1068 B.n52 B.n51 585
R1069 B.n1034 B.n1033 585
R1070 B.n1033 B.n1032 585
R1071 B.n54 B.n53 585
R1072 B.n1031 B.n54 585
R1073 B.n1029 B.n1028 585
R1074 B.n1030 B.n1029 585
R1075 B.n1027 B.n59 585
R1076 B.n59 B.n58 585
R1077 B.n1026 B.n1025 585
R1078 B.n1025 B.n1024 585
R1079 B.n61 B.n60 585
R1080 B.n1023 B.n61 585
R1081 B.n1021 B.n1020 585
R1082 B.n1022 B.n1021 585
R1083 B.n1019 B.n66 585
R1084 B.n66 B.n65 585
R1085 B.n1018 B.n1017 585
R1086 B.n1017 B.n1016 585
R1087 B.n68 B.n67 585
R1088 B.n1015 B.n68 585
R1089 B.n1013 B.n1012 585
R1090 B.n1014 B.n1013 585
R1091 B.n1011 B.n73 585
R1092 B.n73 B.n72 585
R1093 B.n1010 B.n1009 585
R1094 B.n1009 B.n1008 585
R1095 B.n75 B.n74 585
R1096 B.n1007 B.n75 585
R1097 B.n1005 B.n1004 585
R1098 B.n1006 B.n1005 585
R1099 B.n1003 B.n80 585
R1100 B.n80 B.n79 585
R1101 B.n1002 B.n1001 585
R1102 B.n1001 B.n1000 585
R1103 B.n82 B.n81 585
R1104 B.n999 B.n82 585
R1105 B.n997 B.n996 585
R1106 B.n998 B.n997 585
R1107 B.n995 B.n87 585
R1108 B.n87 B.n86 585
R1109 B.n994 B.n993 585
R1110 B.n993 B.n992 585
R1111 B.n89 B.n88 585
R1112 B.n991 B.n89 585
R1113 B.n989 B.n988 585
R1114 B.n990 B.n989 585
R1115 B.n987 B.n94 585
R1116 B.n94 B.n93 585
R1117 B.n986 B.n985 585
R1118 B.n985 B.n984 585
R1119 B.n96 B.n95 585
R1120 B.n983 B.n96 585
R1121 B.n981 B.n980 585
R1122 B.n982 B.n981 585
R1123 B.n979 B.n101 585
R1124 B.n101 B.n100 585
R1125 B.n978 B.n977 585
R1126 B.n977 B.n976 585
R1127 B.n103 B.n102 585
R1128 B.n975 B.n103 585
R1129 B.n973 B.n972 585
R1130 B.n974 B.n973 585
R1131 B.n971 B.n107 585
R1132 B.n110 B.n107 585
R1133 B.n970 B.n969 585
R1134 B.n969 B.n968 585
R1135 B.n109 B.n108 585
R1136 B.n967 B.n109 585
R1137 B.n965 B.n964 585
R1138 B.n966 B.n965 585
R1139 B.n963 B.n115 585
R1140 B.n115 B.n114 585
R1141 B.n962 B.n961 585
R1142 B.n961 B.n960 585
R1143 B.n117 B.n116 585
R1144 B.n959 B.n117 585
R1145 B.n957 B.n956 585
R1146 B.n958 B.n957 585
R1147 B.n955 B.n122 585
R1148 B.n122 B.n121 585
R1149 B.n954 B.n953 585
R1150 B.n953 B.n952 585
R1151 B.n124 B.n123 585
R1152 B.n951 B.n124 585
R1153 B.n949 B.n948 585
R1154 B.n950 B.n949 585
R1155 B.n947 B.n129 585
R1156 B.n129 B.n128 585
R1157 B.n946 B.n945 585
R1158 B.n945 B.n944 585
R1159 B.n131 B.n130 585
R1160 B.n943 B.n131 585
R1161 B.n941 B.n940 585
R1162 B.n942 B.n941 585
R1163 B.n939 B.n135 585
R1164 B.n138 B.n135 585
R1165 B.n938 B.n937 585
R1166 B.n937 B.n936 585
R1167 B.n137 B.n136 585
R1168 B.n935 B.n137 585
R1169 B.n933 B.n932 585
R1170 B.n934 B.n933 585
R1171 B.n931 B.n143 585
R1172 B.n143 B.n142 585
R1173 B.n930 B.n929 585
R1174 B.n929 B.n928 585
R1175 B.n145 B.n144 585
R1176 B.n927 B.n145 585
R1177 B.n925 B.n924 585
R1178 B.n926 B.n925 585
R1179 B.n923 B.n150 585
R1180 B.n150 B.n149 585
R1181 B.n922 B.n921 585
R1182 B.n921 B.n920 585
R1183 B.n1090 B.n1089 585
R1184 B.n1088 B.n2 585
R1185 B.n921 B.n152 502.111
R1186 B.n917 B.n153 502.111
R1187 B.n554 B.n435 502.111
R1188 B.n556 B.n433 502.111
R1189 B.n919 B.n918 256.663
R1190 B.n919 B.n175 256.663
R1191 B.n919 B.n174 256.663
R1192 B.n919 B.n173 256.663
R1193 B.n919 B.n172 256.663
R1194 B.n919 B.n171 256.663
R1195 B.n919 B.n170 256.663
R1196 B.n919 B.n169 256.663
R1197 B.n919 B.n168 256.663
R1198 B.n919 B.n167 256.663
R1199 B.n919 B.n166 256.663
R1200 B.n919 B.n165 256.663
R1201 B.n919 B.n164 256.663
R1202 B.n919 B.n163 256.663
R1203 B.n919 B.n162 256.663
R1204 B.n919 B.n161 256.663
R1205 B.n919 B.n160 256.663
R1206 B.n919 B.n159 256.663
R1207 B.n919 B.n158 256.663
R1208 B.n919 B.n157 256.663
R1209 B.n919 B.n156 256.663
R1210 B.n919 B.n155 256.663
R1211 B.n919 B.n154 256.663
R1212 B.n461 B.n434 256.663
R1213 B.n464 B.n434 256.663
R1214 B.n470 B.n434 256.663
R1215 B.n472 B.n434 256.663
R1216 B.n478 B.n434 256.663
R1217 B.n480 B.n434 256.663
R1218 B.n486 B.n434 256.663
R1219 B.n488 B.n434 256.663
R1220 B.n497 B.n434 256.663
R1221 B.n499 B.n434 256.663
R1222 B.n505 B.n434 256.663
R1223 B.n507 B.n434 256.663
R1224 B.n513 B.n434 256.663
R1225 B.n515 B.n434 256.663
R1226 B.n522 B.n434 256.663
R1227 B.n524 B.n434 256.663
R1228 B.n530 B.n434 256.663
R1229 B.n532 B.n434 256.663
R1230 B.n538 B.n434 256.663
R1231 B.n540 B.n434 256.663
R1232 B.n546 B.n434 256.663
R1233 B.n549 B.n434 256.663
R1234 B.n1092 B.n1091 256.663
R1235 B.n180 B.t10 233.833
R1236 B.n177 B.t21 233.833
R1237 B.n445 B.t18 233.833
R1238 B.n492 B.t14 233.833
R1239 B.n177 B.t22 230.012
R1240 B.n445 B.t20 230.012
R1241 B.n180 B.t12 230.012
R1242 B.n492 B.t17 230.012
R1243 B.n185 B.n184 163.367
R1244 B.n189 B.n188 163.367
R1245 B.n193 B.n192 163.367
R1246 B.n197 B.n196 163.367
R1247 B.n201 B.n200 163.367
R1248 B.n205 B.n204 163.367
R1249 B.n209 B.n208 163.367
R1250 B.n213 B.n212 163.367
R1251 B.n217 B.n216 163.367
R1252 B.n221 B.n220 163.367
R1253 B.n225 B.n224 163.367
R1254 B.n229 B.n228 163.367
R1255 B.n233 B.n232 163.367
R1256 B.n237 B.n236 163.367
R1257 B.n241 B.n240 163.367
R1258 B.n245 B.n244 163.367
R1259 B.n249 B.n248 163.367
R1260 B.n253 B.n252 163.367
R1261 B.n257 B.n256 163.367
R1262 B.n261 B.n260 163.367
R1263 B.n265 B.n264 163.367
R1264 B.n267 B.n176 163.367
R1265 B.n554 B.n429 163.367
R1266 B.n562 B.n429 163.367
R1267 B.n562 B.n427 163.367
R1268 B.n566 B.n427 163.367
R1269 B.n566 B.n421 163.367
R1270 B.n574 B.n421 163.367
R1271 B.n574 B.n419 163.367
R1272 B.n578 B.n419 163.367
R1273 B.n578 B.n414 163.367
R1274 B.n587 B.n414 163.367
R1275 B.n587 B.n412 163.367
R1276 B.n591 B.n412 163.367
R1277 B.n591 B.n406 163.367
R1278 B.n599 B.n406 163.367
R1279 B.n599 B.n404 163.367
R1280 B.n603 B.n404 163.367
R1281 B.n603 B.n398 163.367
R1282 B.n611 B.n398 163.367
R1283 B.n611 B.n396 163.367
R1284 B.n615 B.n396 163.367
R1285 B.n615 B.n390 163.367
R1286 B.n623 B.n390 163.367
R1287 B.n623 B.n388 163.367
R1288 B.n627 B.n388 163.367
R1289 B.n627 B.n383 163.367
R1290 B.n636 B.n383 163.367
R1291 B.n636 B.n381 163.367
R1292 B.n640 B.n381 163.367
R1293 B.n640 B.n375 163.367
R1294 B.n648 B.n375 163.367
R1295 B.n648 B.n373 163.367
R1296 B.n652 B.n373 163.367
R1297 B.n652 B.n367 163.367
R1298 B.n660 B.n367 163.367
R1299 B.n660 B.n365 163.367
R1300 B.n664 B.n365 163.367
R1301 B.n664 B.n359 163.367
R1302 B.n672 B.n359 163.367
R1303 B.n672 B.n357 163.367
R1304 B.n676 B.n357 163.367
R1305 B.n676 B.n351 163.367
R1306 B.n684 B.n351 163.367
R1307 B.n684 B.n349 163.367
R1308 B.n688 B.n349 163.367
R1309 B.n688 B.n343 163.367
R1310 B.n696 B.n343 163.367
R1311 B.n696 B.n341 163.367
R1312 B.n700 B.n341 163.367
R1313 B.n700 B.n334 163.367
R1314 B.n708 B.n334 163.367
R1315 B.n708 B.n332 163.367
R1316 B.n712 B.n332 163.367
R1317 B.n712 B.n327 163.367
R1318 B.n720 B.n327 163.367
R1319 B.n720 B.n325 163.367
R1320 B.n724 B.n325 163.367
R1321 B.n724 B.n319 163.367
R1322 B.n732 B.n319 163.367
R1323 B.n732 B.n317 163.367
R1324 B.n736 B.n317 163.367
R1325 B.n736 B.n310 163.367
R1326 B.n744 B.n310 163.367
R1327 B.n744 B.n308 163.367
R1328 B.n748 B.n308 163.367
R1329 B.n748 B.n303 163.367
R1330 B.n756 B.n303 163.367
R1331 B.n756 B.n301 163.367
R1332 B.n760 B.n301 163.367
R1333 B.n760 B.n295 163.367
R1334 B.n768 B.n295 163.367
R1335 B.n768 B.n293 163.367
R1336 B.n772 B.n293 163.367
R1337 B.n772 B.n287 163.367
R1338 B.n780 B.n287 163.367
R1339 B.n780 B.n285 163.367
R1340 B.n784 B.n285 163.367
R1341 B.n784 B.n279 163.367
R1342 B.n792 B.n279 163.367
R1343 B.n792 B.n277 163.367
R1344 B.n797 B.n277 163.367
R1345 B.n797 B.n271 163.367
R1346 B.n805 B.n271 163.367
R1347 B.n806 B.n805 163.367
R1348 B.n806 B.n5 163.367
R1349 B.n6 B.n5 163.367
R1350 B.n7 B.n6 163.367
R1351 B.n812 B.n7 163.367
R1352 B.n813 B.n812 163.367
R1353 B.n813 B.n13 163.367
R1354 B.n14 B.n13 163.367
R1355 B.n15 B.n14 163.367
R1356 B.n818 B.n15 163.367
R1357 B.n818 B.n20 163.367
R1358 B.n21 B.n20 163.367
R1359 B.n22 B.n21 163.367
R1360 B.n823 B.n22 163.367
R1361 B.n823 B.n27 163.367
R1362 B.n28 B.n27 163.367
R1363 B.n29 B.n28 163.367
R1364 B.n828 B.n29 163.367
R1365 B.n828 B.n34 163.367
R1366 B.n35 B.n34 163.367
R1367 B.n36 B.n35 163.367
R1368 B.n833 B.n36 163.367
R1369 B.n833 B.n41 163.367
R1370 B.n42 B.n41 163.367
R1371 B.n43 B.n42 163.367
R1372 B.n838 B.n43 163.367
R1373 B.n838 B.n48 163.367
R1374 B.n49 B.n48 163.367
R1375 B.n50 B.n49 163.367
R1376 B.n843 B.n50 163.367
R1377 B.n843 B.n55 163.367
R1378 B.n56 B.n55 163.367
R1379 B.n57 B.n56 163.367
R1380 B.n848 B.n57 163.367
R1381 B.n848 B.n62 163.367
R1382 B.n63 B.n62 163.367
R1383 B.n64 B.n63 163.367
R1384 B.n853 B.n64 163.367
R1385 B.n853 B.n69 163.367
R1386 B.n70 B.n69 163.367
R1387 B.n71 B.n70 163.367
R1388 B.n858 B.n71 163.367
R1389 B.n858 B.n76 163.367
R1390 B.n77 B.n76 163.367
R1391 B.n78 B.n77 163.367
R1392 B.n863 B.n78 163.367
R1393 B.n863 B.n83 163.367
R1394 B.n84 B.n83 163.367
R1395 B.n85 B.n84 163.367
R1396 B.n868 B.n85 163.367
R1397 B.n868 B.n90 163.367
R1398 B.n91 B.n90 163.367
R1399 B.n92 B.n91 163.367
R1400 B.n873 B.n92 163.367
R1401 B.n873 B.n97 163.367
R1402 B.n98 B.n97 163.367
R1403 B.n99 B.n98 163.367
R1404 B.n878 B.n99 163.367
R1405 B.n878 B.n104 163.367
R1406 B.n105 B.n104 163.367
R1407 B.n106 B.n105 163.367
R1408 B.n883 B.n106 163.367
R1409 B.n883 B.n111 163.367
R1410 B.n112 B.n111 163.367
R1411 B.n113 B.n112 163.367
R1412 B.n888 B.n113 163.367
R1413 B.n888 B.n118 163.367
R1414 B.n119 B.n118 163.367
R1415 B.n120 B.n119 163.367
R1416 B.n893 B.n120 163.367
R1417 B.n893 B.n125 163.367
R1418 B.n126 B.n125 163.367
R1419 B.n127 B.n126 163.367
R1420 B.n898 B.n127 163.367
R1421 B.n898 B.n132 163.367
R1422 B.n133 B.n132 163.367
R1423 B.n134 B.n133 163.367
R1424 B.n903 B.n134 163.367
R1425 B.n903 B.n139 163.367
R1426 B.n140 B.n139 163.367
R1427 B.n141 B.n140 163.367
R1428 B.n908 B.n141 163.367
R1429 B.n908 B.n146 163.367
R1430 B.n147 B.n146 163.367
R1431 B.n148 B.n147 163.367
R1432 B.n913 B.n148 163.367
R1433 B.n913 B.n153 163.367
R1434 B.n463 B.n462 163.367
R1435 B.n465 B.n463 163.367
R1436 B.n469 B.n458 163.367
R1437 B.n473 B.n471 163.367
R1438 B.n477 B.n456 163.367
R1439 B.n481 B.n479 163.367
R1440 B.n485 B.n454 163.367
R1441 B.n489 B.n487 163.367
R1442 B.n496 B.n452 163.367
R1443 B.n500 B.n498 163.367
R1444 B.n504 B.n450 163.367
R1445 B.n508 B.n506 163.367
R1446 B.n512 B.n448 163.367
R1447 B.n516 B.n514 163.367
R1448 B.n521 B.n444 163.367
R1449 B.n525 B.n523 163.367
R1450 B.n529 B.n442 163.367
R1451 B.n533 B.n531 163.367
R1452 B.n537 B.n440 163.367
R1453 B.n541 B.n539 163.367
R1454 B.n545 B.n438 163.367
R1455 B.n548 B.n547 163.367
R1456 B.n550 B.n435 163.367
R1457 B.n556 B.n431 163.367
R1458 B.n560 B.n431 163.367
R1459 B.n560 B.n425 163.367
R1460 B.n568 B.n425 163.367
R1461 B.n568 B.n423 163.367
R1462 B.n572 B.n423 163.367
R1463 B.n572 B.n417 163.367
R1464 B.n581 B.n417 163.367
R1465 B.n581 B.n415 163.367
R1466 B.n585 B.n415 163.367
R1467 B.n585 B.n410 163.367
R1468 B.n593 B.n410 163.367
R1469 B.n593 B.n408 163.367
R1470 B.n597 B.n408 163.367
R1471 B.n597 B.n402 163.367
R1472 B.n605 B.n402 163.367
R1473 B.n605 B.n400 163.367
R1474 B.n609 B.n400 163.367
R1475 B.n609 B.n394 163.367
R1476 B.n617 B.n394 163.367
R1477 B.n617 B.n392 163.367
R1478 B.n621 B.n392 163.367
R1479 B.n621 B.n386 163.367
R1480 B.n630 B.n386 163.367
R1481 B.n630 B.n384 163.367
R1482 B.n634 B.n384 163.367
R1483 B.n634 B.n379 163.367
R1484 B.n642 B.n379 163.367
R1485 B.n642 B.n377 163.367
R1486 B.n646 B.n377 163.367
R1487 B.n646 B.n371 163.367
R1488 B.n654 B.n371 163.367
R1489 B.n654 B.n369 163.367
R1490 B.n658 B.n369 163.367
R1491 B.n658 B.n363 163.367
R1492 B.n666 B.n363 163.367
R1493 B.n666 B.n361 163.367
R1494 B.n670 B.n361 163.367
R1495 B.n670 B.n355 163.367
R1496 B.n678 B.n355 163.367
R1497 B.n678 B.n353 163.367
R1498 B.n682 B.n353 163.367
R1499 B.n682 B.n347 163.367
R1500 B.n690 B.n347 163.367
R1501 B.n690 B.n345 163.367
R1502 B.n694 B.n345 163.367
R1503 B.n694 B.n339 163.367
R1504 B.n702 B.n339 163.367
R1505 B.n702 B.n337 163.367
R1506 B.n706 B.n337 163.367
R1507 B.n706 B.n331 163.367
R1508 B.n714 B.n331 163.367
R1509 B.n714 B.n329 163.367
R1510 B.n718 B.n329 163.367
R1511 B.n718 B.n323 163.367
R1512 B.n726 B.n323 163.367
R1513 B.n726 B.n321 163.367
R1514 B.n730 B.n321 163.367
R1515 B.n730 B.n315 163.367
R1516 B.n738 B.n315 163.367
R1517 B.n738 B.n313 163.367
R1518 B.n742 B.n313 163.367
R1519 B.n742 B.n307 163.367
R1520 B.n750 B.n307 163.367
R1521 B.n750 B.n305 163.367
R1522 B.n754 B.n305 163.367
R1523 B.n754 B.n299 163.367
R1524 B.n762 B.n299 163.367
R1525 B.n762 B.n297 163.367
R1526 B.n766 B.n297 163.367
R1527 B.n766 B.n291 163.367
R1528 B.n774 B.n291 163.367
R1529 B.n774 B.n289 163.367
R1530 B.n778 B.n289 163.367
R1531 B.n778 B.n283 163.367
R1532 B.n786 B.n283 163.367
R1533 B.n786 B.n281 163.367
R1534 B.n790 B.n281 163.367
R1535 B.n790 B.n275 163.367
R1536 B.n799 B.n275 163.367
R1537 B.n799 B.n273 163.367
R1538 B.n803 B.n273 163.367
R1539 B.n803 B.n3 163.367
R1540 B.n1090 B.n3 163.367
R1541 B.n1086 B.n2 163.367
R1542 B.n1086 B.n1085 163.367
R1543 B.n1085 B.n9 163.367
R1544 B.n1081 B.n9 163.367
R1545 B.n1081 B.n11 163.367
R1546 B.n1077 B.n11 163.367
R1547 B.n1077 B.n17 163.367
R1548 B.n1073 B.n17 163.367
R1549 B.n1073 B.n19 163.367
R1550 B.n1069 B.n19 163.367
R1551 B.n1069 B.n24 163.367
R1552 B.n1065 B.n24 163.367
R1553 B.n1065 B.n26 163.367
R1554 B.n1061 B.n26 163.367
R1555 B.n1061 B.n31 163.367
R1556 B.n1057 B.n31 163.367
R1557 B.n1057 B.n33 163.367
R1558 B.n1053 B.n33 163.367
R1559 B.n1053 B.n38 163.367
R1560 B.n1049 B.n38 163.367
R1561 B.n1049 B.n40 163.367
R1562 B.n1045 B.n40 163.367
R1563 B.n1045 B.n45 163.367
R1564 B.n1041 B.n45 163.367
R1565 B.n1041 B.n47 163.367
R1566 B.n1037 B.n47 163.367
R1567 B.n1037 B.n52 163.367
R1568 B.n1033 B.n52 163.367
R1569 B.n1033 B.n54 163.367
R1570 B.n1029 B.n54 163.367
R1571 B.n1029 B.n59 163.367
R1572 B.n1025 B.n59 163.367
R1573 B.n1025 B.n61 163.367
R1574 B.n1021 B.n61 163.367
R1575 B.n1021 B.n66 163.367
R1576 B.n1017 B.n66 163.367
R1577 B.n1017 B.n68 163.367
R1578 B.n1013 B.n68 163.367
R1579 B.n1013 B.n73 163.367
R1580 B.n1009 B.n73 163.367
R1581 B.n1009 B.n75 163.367
R1582 B.n1005 B.n75 163.367
R1583 B.n1005 B.n80 163.367
R1584 B.n1001 B.n80 163.367
R1585 B.n1001 B.n82 163.367
R1586 B.n997 B.n82 163.367
R1587 B.n997 B.n87 163.367
R1588 B.n993 B.n87 163.367
R1589 B.n993 B.n89 163.367
R1590 B.n989 B.n89 163.367
R1591 B.n989 B.n94 163.367
R1592 B.n985 B.n94 163.367
R1593 B.n985 B.n96 163.367
R1594 B.n981 B.n96 163.367
R1595 B.n981 B.n101 163.367
R1596 B.n977 B.n101 163.367
R1597 B.n977 B.n103 163.367
R1598 B.n973 B.n103 163.367
R1599 B.n973 B.n107 163.367
R1600 B.n969 B.n107 163.367
R1601 B.n969 B.n109 163.367
R1602 B.n965 B.n109 163.367
R1603 B.n965 B.n115 163.367
R1604 B.n961 B.n115 163.367
R1605 B.n961 B.n117 163.367
R1606 B.n957 B.n117 163.367
R1607 B.n957 B.n122 163.367
R1608 B.n953 B.n122 163.367
R1609 B.n953 B.n124 163.367
R1610 B.n949 B.n124 163.367
R1611 B.n949 B.n129 163.367
R1612 B.n945 B.n129 163.367
R1613 B.n945 B.n131 163.367
R1614 B.n941 B.n131 163.367
R1615 B.n941 B.n135 163.367
R1616 B.n937 B.n135 163.367
R1617 B.n937 B.n137 163.367
R1618 B.n933 B.n137 163.367
R1619 B.n933 B.n143 163.367
R1620 B.n929 B.n143 163.367
R1621 B.n929 B.n145 163.367
R1622 B.n925 B.n145 163.367
R1623 B.n925 B.n150 163.367
R1624 B.n921 B.n150 163.367
R1625 B.n555 B.n434 147.612
R1626 B.n920 B.n919 147.612
R1627 B.n178 B.t23 146.036
R1628 B.n446 B.t19 146.036
R1629 B.n181 B.t13 146.036
R1630 B.n493 B.t16 146.036
R1631 B.n181 B.n180 83.9763
R1632 B.n178 B.n177 83.9763
R1633 B.n446 B.n445 83.9763
R1634 B.n493 B.n492 83.9763
R1635 B.n555 B.n430 80.3011
R1636 B.n561 B.n430 80.3011
R1637 B.n561 B.n426 80.3011
R1638 B.n567 B.n426 80.3011
R1639 B.n567 B.n422 80.3011
R1640 B.n573 B.n422 80.3011
R1641 B.n573 B.n418 80.3011
R1642 B.n580 B.n418 80.3011
R1643 B.n580 B.n579 80.3011
R1644 B.n586 B.n411 80.3011
R1645 B.n592 B.n411 80.3011
R1646 B.n592 B.n407 80.3011
R1647 B.n598 B.n407 80.3011
R1648 B.n598 B.n403 80.3011
R1649 B.n604 B.n403 80.3011
R1650 B.n604 B.n399 80.3011
R1651 B.n610 B.n399 80.3011
R1652 B.n610 B.n395 80.3011
R1653 B.n616 B.n395 80.3011
R1654 B.n616 B.n391 80.3011
R1655 B.n622 B.n391 80.3011
R1656 B.n622 B.n387 80.3011
R1657 B.n629 B.n387 80.3011
R1658 B.n629 B.n628 80.3011
R1659 B.n635 B.n380 80.3011
R1660 B.n641 B.n380 80.3011
R1661 B.n641 B.n376 80.3011
R1662 B.n647 B.n376 80.3011
R1663 B.n647 B.n372 80.3011
R1664 B.n653 B.n372 80.3011
R1665 B.n653 B.n368 80.3011
R1666 B.n659 B.n368 80.3011
R1667 B.n659 B.n364 80.3011
R1668 B.n665 B.n364 80.3011
R1669 B.n665 B.n360 80.3011
R1670 B.n671 B.n360 80.3011
R1671 B.n677 B.n356 80.3011
R1672 B.n677 B.n352 80.3011
R1673 B.n683 B.n352 80.3011
R1674 B.n683 B.n348 80.3011
R1675 B.n689 B.n348 80.3011
R1676 B.n689 B.n344 80.3011
R1677 B.n695 B.n344 80.3011
R1678 B.n695 B.n340 80.3011
R1679 B.n701 B.n340 80.3011
R1680 B.n701 B.n335 80.3011
R1681 B.n707 B.n335 80.3011
R1682 B.n707 B.n336 80.3011
R1683 B.n713 B.n328 80.3011
R1684 B.n719 B.n328 80.3011
R1685 B.n719 B.n324 80.3011
R1686 B.n725 B.n324 80.3011
R1687 B.n725 B.n320 80.3011
R1688 B.n731 B.n320 80.3011
R1689 B.n731 B.n316 80.3011
R1690 B.n737 B.n316 80.3011
R1691 B.n737 B.n311 80.3011
R1692 B.n743 B.n311 80.3011
R1693 B.n743 B.n312 80.3011
R1694 B.n749 B.n304 80.3011
R1695 B.n755 B.n304 80.3011
R1696 B.n755 B.n300 80.3011
R1697 B.n761 B.n300 80.3011
R1698 B.n761 B.n296 80.3011
R1699 B.n767 B.n296 80.3011
R1700 B.n767 B.n292 80.3011
R1701 B.n773 B.n292 80.3011
R1702 B.n773 B.n288 80.3011
R1703 B.n779 B.n288 80.3011
R1704 B.n779 B.n284 80.3011
R1705 B.n785 B.n284 80.3011
R1706 B.n791 B.n280 80.3011
R1707 B.n791 B.n276 80.3011
R1708 B.n798 B.n276 80.3011
R1709 B.n798 B.n272 80.3011
R1710 B.n804 B.n272 80.3011
R1711 B.n804 B.n4 80.3011
R1712 B.n1089 B.n4 80.3011
R1713 B.n1089 B.n1088 80.3011
R1714 B.n1088 B.n1087 80.3011
R1715 B.n1087 B.n8 80.3011
R1716 B.n12 B.n8 80.3011
R1717 B.n1080 B.n12 80.3011
R1718 B.n1080 B.n1079 80.3011
R1719 B.n1079 B.n1078 80.3011
R1720 B.n1078 B.n16 80.3011
R1721 B.n1072 B.n1071 80.3011
R1722 B.n1071 B.n1070 80.3011
R1723 B.n1070 B.n23 80.3011
R1724 B.n1064 B.n23 80.3011
R1725 B.n1064 B.n1063 80.3011
R1726 B.n1063 B.n1062 80.3011
R1727 B.n1062 B.n30 80.3011
R1728 B.n1056 B.n30 80.3011
R1729 B.n1056 B.n1055 80.3011
R1730 B.n1055 B.n1054 80.3011
R1731 B.n1054 B.n37 80.3011
R1732 B.n1048 B.n37 80.3011
R1733 B.n1047 B.n1046 80.3011
R1734 B.n1046 B.n44 80.3011
R1735 B.n1040 B.n44 80.3011
R1736 B.n1040 B.n1039 80.3011
R1737 B.n1039 B.n1038 80.3011
R1738 B.n1038 B.n51 80.3011
R1739 B.n1032 B.n51 80.3011
R1740 B.n1032 B.n1031 80.3011
R1741 B.n1031 B.n1030 80.3011
R1742 B.n1030 B.n58 80.3011
R1743 B.n1024 B.n58 80.3011
R1744 B.n1023 B.n1022 80.3011
R1745 B.n1022 B.n65 80.3011
R1746 B.n1016 B.n65 80.3011
R1747 B.n1016 B.n1015 80.3011
R1748 B.n1015 B.n1014 80.3011
R1749 B.n1014 B.n72 80.3011
R1750 B.n1008 B.n72 80.3011
R1751 B.n1008 B.n1007 80.3011
R1752 B.n1007 B.n1006 80.3011
R1753 B.n1006 B.n79 80.3011
R1754 B.n1000 B.n79 80.3011
R1755 B.n1000 B.n999 80.3011
R1756 B.n998 B.n86 80.3011
R1757 B.n992 B.n86 80.3011
R1758 B.n992 B.n991 80.3011
R1759 B.n991 B.n990 80.3011
R1760 B.n990 B.n93 80.3011
R1761 B.n984 B.n93 80.3011
R1762 B.n984 B.n983 80.3011
R1763 B.n983 B.n982 80.3011
R1764 B.n982 B.n100 80.3011
R1765 B.n976 B.n100 80.3011
R1766 B.n976 B.n975 80.3011
R1767 B.n975 B.n974 80.3011
R1768 B.n968 B.n110 80.3011
R1769 B.n968 B.n967 80.3011
R1770 B.n967 B.n966 80.3011
R1771 B.n966 B.n114 80.3011
R1772 B.n960 B.n114 80.3011
R1773 B.n960 B.n959 80.3011
R1774 B.n959 B.n958 80.3011
R1775 B.n958 B.n121 80.3011
R1776 B.n952 B.n121 80.3011
R1777 B.n952 B.n951 80.3011
R1778 B.n951 B.n950 80.3011
R1779 B.n950 B.n128 80.3011
R1780 B.n944 B.n128 80.3011
R1781 B.n944 B.n943 80.3011
R1782 B.n943 B.n942 80.3011
R1783 B.n936 B.n138 80.3011
R1784 B.n936 B.n935 80.3011
R1785 B.n935 B.n934 80.3011
R1786 B.n934 B.n142 80.3011
R1787 B.n928 B.n142 80.3011
R1788 B.n928 B.n927 80.3011
R1789 B.n927 B.n926 80.3011
R1790 B.n926 B.n149 80.3011
R1791 B.n920 B.n149 80.3011
R1792 B.n713 B.t9 75.5775
R1793 B.n1024 B.t0 75.5775
R1794 B.n154 B.n152 71.676
R1795 B.n185 B.n155 71.676
R1796 B.n189 B.n156 71.676
R1797 B.n193 B.n157 71.676
R1798 B.n197 B.n158 71.676
R1799 B.n201 B.n159 71.676
R1800 B.n205 B.n160 71.676
R1801 B.n209 B.n161 71.676
R1802 B.n213 B.n162 71.676
R1803 B.n217 B.n163 71.676
R1804 B.n221 B.n164 71.676
R1805 B.n225 B.n165 71.676
R1806 B.n229 B.n166 71.676
R1807 B.n233 B.n167 71.676
R1808 B.n237 B.n168 71.676
R1809 B.n241 B.n169 71.676
R1810 B.n245 B.n170 71.676
R1811 B.n249 B.n171 71.676
R1812 B.n253 B.n172 71.676
R1813 B.n257 B.n173 71.676
R1814 B.n261 B.n174 71.676
R1815 B.n265 B.n175 71.676
R1816 B.n918 B.n176 71.676
R1817 B.n918 B.n917 71.676
R1818 B.n267 B.n175 71.676
R1819 B.n264 B.n174 71.676
R1820 B.n260 B.n173 71.676
R1821 B.n256 B.n172 71.676
R1822 B.n252 B.n171 71.676
R1823 B.n248 B.n170 71.676
R1824 B.n244 B.n169 71.676
R1825 B.n240 B.n168 71.676
R1826 B.n236 B.n167 71.676
R1827 B.n232 B.n166 71.676
R1828 B.n228 B.n165 71.676
R1829 B.n224 B.n164 71.676
R1830 B.n220 B.n163 71.676
R1831 B.n216 B.n162 71.676
R1832 B.n212 B.n161 71.676
R1833 B.n208 B.n160 71.676
R1834 B.n204 B.n159 71.676
R1835 B.n200 B.n158 71.676
R1836 B.n196 B.n157 71.676
R1837 B.n192 B.n156 71.676
R1838 B.n188 B.n155 71.676
R1839 B.n184 B.n154 71.676
R1840 B.n461 B.n433 71.676
R1841 B.n465 B.n464 71.676
R1842 B.n470 B.n469 71.676
R1843 B.n473 B.n472 71.676
R1844 B.n478 B.n477 71.676
R1845 B.n481 B.n480 71.676
R1846 B.n486 B.n485 71.676
R1847 B.n489 B.n488 71.676
R1848 B.n497 B.n496 71.676
R1849 B.n500 B.n499 71.676
R1850 B.n505 B.n504 71.676
R1851 B.n508 B.n507 71.676
R1852 B.n513 B.n512 71.676
R1853 B.n516 B.n515 71.676
R1854 B.n522 B.n521 71.676
R1855 B.n525 B.n524 71.676
R1856 B.n530 B.n529 71.676
R1857 B.n533 B.n532 71.676
R1858 B.n538 B.n537 71.676
R1859 B.n541 B.n540 71.676
R1860 B.n546 B.n545 71.676
R1861 B.n549 B.n548 71.676
R1862 B.n462 B.n461 71.676
R1863 B.n464 B.n458 71.676
R1864 B.n471 B.n470 71.676
R1865 B.n472 B.n456 71.676
R1866 B.n479 B.n478 71.676
R1867 B.n480 B.n454 71.676
R1868 B.n487 B.n486 71.676
R1869 B.n488 B.n452 71.676
R1870 B.n498 B.n497 71.676
R1871 B.n499 B.n450 71.676
R1872 B.n506 B.n505 71.676
R1873 B.n507 B.n448 71.676
R1874 B.n514 B.n513 71.676
R1875 B.n515 B.n444 71.676
R1876 B.n523 B.n522 71.676
R1877 B.n524 B.n442 71.676
R1878 B.n531 B.n530 71.676
R1879 B.n532 B.n440 71.676
R1880 B.n539 B.n538 71.676
R1881 B.n540 B.n438 71.676
R1882 B.n547 B.n546 71.676
R1883 B.n550 B.n549 71.676
R1884 B.n1091 B.n1090 71.676
R1885 B.n1091 B.n2 71.676
R1886 B.n312 B.t6 63.7686
R1887 B.t7 B.n1047 63.7686
R1888 B.n182 B.n181 59.5399
R1889 B.n179 B.n178 59.5399
R1890 B.n518 B.n446 59.5399
R1891 B.n494 B.n493 59.5399
R1892 B.t2 B.n356 54.3215
R1893 B.n999 B.t8 54.3215
R1894 B.n579 B.t15 51.9597
R1895 B.n138 B.t11 51.9597
R1896 B.n628 B.t5 47.2361
R1897 B.n110 B.t1 47.2361
R1898 B.n785 B.t4 42.5126
R1899 B.n1072 B.t3 42.5126
R1900 B.t4 B.n280 37.789
R1901 B.t3 B.n16 37.789
R1902 B.n635 B.t5 33.0654
R1903 B.n974 B.t1 33.0654
R1904 B.n557 B.n432 32.6249
R1905 B.n553 B.n552 32.6249
R1906 B.n916 B.n915 32.6249
R1907 B.n922 B.n151 32.6249
R1908 B.n586 B.t15 28.3419
R1909 B.n942 B.t11 28.3419
R1910 B.n671 B.t2 25.9801
R1911 B.t8 B.n998 25.9801
R1912 B B.n1092 18.0485
R1913 B.n749 B.t6 16.533
R1914 B.n1048 B.t7 16.533
R1915 B.n558 B.n557 10.6151
R1916 B.n559 B.n558 10.6151
R1917 B.n559 B.n424 10.6151
R1918 B.n569 B.n424 10.6151
R1919 B.n570 B.n569 10.6151
R1920 B.n571 B.n570 10.6151
R1921 B.n571 B.n416 10.6151
R1922 B.n582 B.n416 10.6151
R1923 B.n583 B.n582 10.6151
R1924 B.n584 B.n583 10.6151
R1925 B.n584 B.n409 10.6151
R1926 B.n594 B.n409 10.6151
R1927 B.n595 B.n594 10.6151
R1928 B.n596 B.n595 10.6151
R1929 B.n596 B.n401 10.6151
R1930 B.n606 B.n401 10.6151
R1931 B.n607 B.n606 10.6151
R1932 B.n608 B.n607 10.6151
R1933 B.n608 B.n393 10.6151
R1934 B.n618 B.n393 10.6151
R1935 B.n619 B.n618 10.6151
R1936 B.n620 B.n619 10.6151
R1937 B.n620 B.n385 10.6151
R1938 B.n631 B.n385 10.6151
R1939 B.n632 B.n631 10.6151
R1940 B.n633 B.n632 10.6151
R1941 B.n633 B.n378 10.6151
R1942 B.n643 B.n378 10.6151
R1943 B.n644 B.n643 10.6151
R1944 B.n645 B.n644 10.6151
R1945 B.n645 B.n370 10.6151
R1946 B.n655 B.n370 10.6151
R1947 B.n656 B.n655 10.6151
R1948 B.n657 B.n656 10.6151
R1949 B.n657 B.n362 10.6151
R1950 B.n667 B.n362 10.6151
R1951 B.n668 B.n667 10.6151
R1952 B.n669 B.n668 10.6151
R1953 B.n669 B.n354 10.6151
R1954 B.n679 B.n354 10.6151
R1955 B.n680 B.n679 10.6151
R1956 B.n681 B.n680 10.6151
R1957 B.n681 B.n346 10.6151
R1958 B.n691 B.n346 10.6151
R1959 B.n692 B.n691 10.6151
R1960 B.n693 B.n692 10.6151
R1961 B.n693 B.n338 10.6151
R1962 B.n703 B.n338 10.6151
R1963 B.n704 B.n703 10.6151
R1964 B.n705 B.n704 10.6151
R1965 B.n705 B.n330 10.6151
R1966 B.n715 B.n330 10.6151
R1967 B.n716 B.n715 10.6151
R1968 B.n717 B.n716 10.6151
R1969 B.n717 B.n322 10.6151
R1970 B.n727 B.n322 10.6151
R1971 B.n728 B.n727 10.6151
R1972 B.n729 B.n728 10.6151
R1973 B.n729 B.n314 10.6151
R1974 B.n739 B.n314 10.6151
R1975 B.n740 B.n739 10.6151
R1976 B.n741 B.n740 10.6151
R1977 B.n741 B.n306 10.6151
R1978 B.n751 B.n306 10.6151
R1979 B.n752 B.n751 10.6151
R1980 B.n753 B.n752 10.6151
R1981 B.n753 B.n298 10.6151
R1982 B.n763 B.n298 10.6151
R1983 B.n764 B.n763 10.6151
R1984 B.n765 B.n764 10.6151
R1985 B.n765 B.n290 10.6151
R1986 B.n775 B.n290 10.6151
R1987 B.n776 B.n775 10.6151
R1988 B.n777 B.n776 10.6151
R1989 B.n777 B.n282 10.6151
R1990 B.n787 B.n282 10.6151
R1991 B.n788 B.n787 10.6151
R1992 B.n789 B.n788 10.6151
R1993 B.n789 B.n274 10.6151
R1994 B.n800 B.n274 10.6151
R1995 B.n801 B.n800 10.6151
R1996 B.n802 B.n801 10.6151
R1997 B.n802 B.n0 10.6151
R1998 B.n460 B.n432 10.6151
R1999 B.n460 B.n459 10.6151
R2000 B.n466 B.n459 10.6151
R2001 B.n467 B.n466 10.6151
R2002 B.n468 B.n467 10.6151
R2003 B.n468 B.n457 10.6151
R2004 B.n474 B.n457 10.6151
R2005 B.n475 B.n474 10.6151
R2006 B.n476 B.n475 10.6151
R2007 B.n476 B.n455 10.6151
R2008 B.n482 B.n455 10.6151
R2009 B.n483 B.n482 10.6151
R2010 B.n484 B.n483 10.6151
R2011 B.n484 B.n453 10.6151
R2012 B.n490 B.n453 10.6151
R2013 B.n491 B.n490 10.6151
R2014 B.n495 B.n491 10.6151
R2015 B.n501 B.n451 10.6151
R2016 B.n502 B.n501 10.6151
R2017 B.n503 B.n502 10.6151
R2018 B.n503 B.n449 10.6151
R2019 B.n509 B.n449 10.6151
R2020 B.n510 B.n509 10.6151
R2021 B.n511 B.n510 10.6151
R2022 B.n511 B.n447 10.6151
R2023 B.n517 B.n447 10.6151
R2024 B.n520 B.n519 10.6151
R2025 B.n520 B.n443 10.6151
R2026 B.n526 B.n443 10.6151
R2027 B.n527 B.n526 10.6151
R2028 B.n528 B.n527 10.6151
R2029 B.n528 B.n441 10.6151
R2030 B.n534 B.n441 10.6151
R2031 B.n535 B.n534 10.6151
R2032 B.n536 B.n535 10.6151
R2033 B.n536 B.n439 10.6151
R2034 B.n542 B.n439 10.6151
R2035 B.n543 B.n542 10.6151
R2036 B.n544 B.n543 10.6151
R2037 B.n544 B.n437 10.6151
R2038 B.n437 B.n436 10.6151
R2039 B.n551 B.n436 10.6151
R2040 B.n552 B.n551 10.6151
R2041 B.n553 B.n428 10.6151
R2042 B.n563 B.n428 10.6151
R2043 B.n564 B.n563 10.6151
R2044 B.n565 B.n564 10.6151
R2045 B.n565 B.n420 10.6151
R2046 B.n575 B.n420 10.6151
R2047 B.n576 B.n575 10.6151
R2048 B.n577 B.n576 10.6151
R2049 B.n577 B.n413 10.6151
R2050 B.n588 B.n413 10.6151
R2051 B.n589 B.n588 10.6151
R2052 B.n590 B.n589 10.6151
R2053 B.n590 B.n405 10.6151
R2054 B.n600 B.n405 10.6151
R2055 B.n601 B.n600 10.6151
R2056 B.n602 B.n601 10.6151
R2057 B.n602 B.n397 10.6151
R2058 B.n612 B.n397 10.6151
R2059 B.n613 B.n612 10.6151
R2060 B.n614 B.n613 10.6151
R2061 B.n614 B.n389 10.6151
R2062 B.n624 B.n389 10.6151
R2063 B.n625 B.n624 10.6151
R2064 B.n626 B.n625 10.6151
R2065 B.n626 B.n382 10.6151
R2066 B.n637 B.n382 10.6151
R2067 B.n638 B.n637 10.6151
R2068 B.n639 B.n638 10.6151
R2069 B.n639 B.n374 10.6151
R2070 B.n649 B.n374 10.6151
R2071 B.n650 B.n649 10.6151
R2072 B.n651 B.n650 10.6151
R2073 B.n651 B.n366 10.6151
R2074 B.n661 B.n366 10.6151
R2075 B.n662 B.n661 10.6151
R2076 B.n663 B.n662 10.6151
R2077 B.n663 B.n358 10.6151
R2078 B.n673 B.n358 10.6151
R2079 B.n674 B.n673 10.6151
R2080 B.n675 B.n674 10.6151
R2081 B.n675 B.n350 10.6151
R2082 B.n685 B.n350 10.6151
R2083 B.n686 B.n685 10.6151
R2084 B.n687 B.n686 10.6151
R2085 B.n687 B.n342 10.6151
R2086 B.n697 B.n342 10.6151
R2087 B.n698 B.n697 10.6151
R2088 B.n699 B.n698 10.6151
R2089 B.n699 B.n333 10.6151
R2090 B.n709 B.n333 10.6151
R2091 B.n710 B.n709 10.6151
R2092 B.n711 B.n710 10.6151
R2093 B.n711 B.n326 10.6151
R2094 B.n721 B.n326 10.6151
R2095 B.n722 B.n721 10.6151
R2096 B.n723 B.n722 10.6151
R2097 B.n723 B.n318 10.6151
R2098 B.n733 B.n318 10.6151
R2099 B.n734 B.n733 10.6151
R2100 B.n735 B.n734 10.6151
R2101 B.n735 B.n309 10.6151
R2102 B.n745 B.n309 10.6151
R2103 B.n746 B.n745 10.6151
R2104 B.n747 B.n746 10.6151
R2105 B.n747 B.n302 10.6151
R2106 B.n757 B.n302 10.6151
R2107 B.n758 B.n757 10.6151
R2108 B.n759 B.n758 10.6151
R2109 B.n759 B.n294 10.6151
R2110 B.n769 B.n294 10.6151
R2111 B.n770 B.n769 10.6151
R2112 B.n771 B.n770 10.6151
R2113 B.n771 B.n286 10.6151
R2114 B.n781 B.n286 10.6151
R2115 B.n782 B.n781 10.6151
R2116 B.n783 B.n782 10.6151
R2117 B.n783 B.n278 10.6151
R2118 B.n793 B.n278 10.6151
R2119 B.n794 B.n793 10.6151
R2120 B.n796 B.n794 10.6151
R2121 B.n796 B.n795 10.6151
R2122 B.n795 B.n270 10.6151
R2123 B.n807 B.n270 10.6151
R2124 B.n808 B.n807 10.6151
R2125 B.n809 B.n808 10.6151
R2126 B.n810 B.n809 10.6151
R2127 B.n811 B.n810 10.6151
R2128 B.n814 B.n811 10.6151
R2129 B.n815 B.n814 10.6151
R2130 B.n816 B.n815 10.6151
R2131 B.n817 B.n816 10.6151
R2132 B.n819 B.n817 10.6151
R2133 B.n820 B.n819 10.6151
R2134 B.n821 B.n820 10.6151
R2135 B.n822 B.n821 10.6151
R2136 B.n824 B.n822 10.6151
R2137 B.n825 B.n824 10.6151
R2138 B.n826 B.n825 10.6151
R2139 B.n827 B.n826 10.6151
R2140 B.n829 B.n827 10.6151
R2141 B.n830 B.n829 10.6151
R2142 B.n831 B.n830 10.6151
R2143 B.n832 B.n831 10.6151
R2144 B.n834 B.n832 10.6151
R2145 B.n835 B.n834 10.6151
R2146 B.n836 B.n835 10.6151
R2147 B.n837 B.n836 10.6151
R2148 B.n839 B.n837 10.6151
R2149 B.n840 B.n839 10.6151
R2150 B.n841 B.n840 10.6151
R2151 B.n842 B.n841 10.6151
R2152 B.n844 B.n842 10.6151
R2153 B.n845 B.n844 10.6151
R2154 B.n846 B.n845 10.6151
R2155 B.n847 B.n846 10.6151
R2156 B.n849 B.n847 10.6151
R2157 B.n850 B.n849 10.6151
R2158 B.n851 B.n850 10.6151
R2159 B.n852 B.n851 10.6151
R2160 B.n854 B.n852 10.6151
R2161 B.n855 B.n854 10.6151
R2162 B.n856 B.n855 10.6151
R2163 B.n857 B.n856 10.6151
R2164 B.n859 B.n857 10.6151
R2165 B.n860 B.n859 10.6151
R2166 B.n861 B.n860 10.6151
R2167 B.n862 B.n861 10.6151
R2168 B.n864 B.n862 10.6151
R2169 B.n865 B.n864 10.6151
R2170 B.n866 B.n865 10.6151
R2171 B.n867 B.n866 10.6151
R2172 B.n869 B.n867 10.6151
R2173 B.n870 B.n869 10.6151
R2174 B.n871 B.n870 10.6151
R2175 B.n872 B.n871 10.6151
R2176 B.n874 B.n872 10.6151
R2177 B.n875 B.n874 10.6151
R2178 B.n876 B.n875 10.6151
R2179 B.n877 B.n876 10.6151
R2180 B.n879 B.n877 10.6151
R2181 B.n880 B.n879 10.6151
R2182 B.n881 B.n880 10.6151
R2183 B.n882 B.n881 10.6151
R2184 B.n884 B.n882 10.6151
R2185 B.n885 B.n884 10.6151
R2186 B.n886 B.n885 10.6151
R2187 B.n887 B.n886 10.6151
R2188 B.n889 B.n887 10.6151
R2189 B.n890 B.n889 10.6151
R2190 B.n891 B.n890 10.6151
R2191 B.n892 B.n891 10.6151
R2192 B.n894 B.n892 10.6151
R2193 B.n895 B.n894 10.6151
R2194 B.n896 B.n895 10.6151
R2195 B.n897 B.n896 10.6151
R2196 B.n899 B.n897 10.6151
R2197 B.n900 B.n899 10.6151
R2198 B.n901 B.n900 10.6151
R2199 B.n902 B.n901 10.6151
R2200 B.n904 B.n902 10.6151
R2201 B.n905 B.n904 10.6151
R2202 B.n906 B.n905 10.6151
R2203 B.n907 B.n906 10.6151
R2204 B.n909 B.n907 10.6151
R2205 B.n910 B.n909 10.6151
R2206 B.n911 B.n910 10.6151
R2207 B.n912 B.n911 10.6151
R2208 B.n914 B.n912 10.6151
R2209 B.n915 B.n914 10.6151
R2210 B.n1084 B.n1 10.6151
R2211 B.n1084 B.n1083 10.6151
R2212 B.n1083 B.n1082 10.6151
R2213 B.n1082 B.n10 10.6151
R2214 B.n1076 B.n10 10.6151
R2215 B.n1076 B.n1075 10.6151
R2216 B.n1075 B.n1074 10.6151
R2217 B.n1074 B.n18 10.6151
R2218 B.n1068 B.n18 10.6151
R2219 B.n1068 B.n1067 10.6151
R2220 B.n1067 B.n1066 10.6151
R2221 B.n1066 B.n25 10.6151
R2222 B.n1060 B.n25 10.6151
R2223 B.n1060 B.n1059 10.6151
R2224 B.n1059 B.n1058 10.6151
R2225 B.n1058 B.n32 10.6151
R2226 B.n1052 B.n32 10.6151
R2227 B.n1052 B.n1051 10.6151
R2228 B.n1051 B.n1050 10.6151
R2229 B.n1050 B.n39 10.6151
R2230 B.n1044 B.n39 10.6151
R2231 B.n1044 B.n1043 10.6151
R2232 B.n1043 B.n1042 10.6151
R2233 B.n1042 B.n46 10.6151
R2234 B.n1036 B.n46 10.6151
R2235 B.n1036 B.n1035 10.6151
R2236 B.n1035 B.n1034 10.6151
R2237 B.n1034 B.n53 10.6151
R2238 B.n1028 B.n53 10.6151
R2239 B.n1028 B.n1027 10.6151
R2240 B.n1027 B.n1026 10.6151
R2241 B.n1026 B.n60 10.6151
R2242 B.n1020 B.n60 10.6151
R2243 B.n1020 B.n1019 10.6151
R2244 B.n1019 B.n1018 10.6151
R2245 B.n1018 B.n67 10.6151
R2246 B.n1012 B.n67 10.6151
R2247 B.n1012 B.n1011 10.6151
R2248 B.n1011 B.n1010 10.6151
R2249 B.n1010 B.n74 10.6151
R2250 B.n1004 B.n74 10.6151
R2251 B.n1004 B.n1003 10.6151
R2252 B.n1003 B.n1002 10.6151
R2253 B.n1002 B.n81 10.6151
R2254 B.n996 B.n81 10.6151
R2255 B.n996 B.n995 10.6151
R2256 B.n995 B.n994 10.6151
R2257 B.n994 B.n88 10.6151
R2258 B.n988 B.n88 10.6151
R2259 B.n988 B.n987 10.6151
R2260 B.n987 B.n986 10.6151
R2261 B.n986 B.n95 10.6151
R2262 B.n980 B.n95 10.6151
R2263 B.n980 B.n979 10.6151
R2264 B.n979 B.n978 10.6151
R2265 B.n978 B.n102 10.6151
R2266 B.n972 B.n102 10.6151
R2267 B.n972 B.n971 10.6151
R2268 B.n971 B.n970 10.6151
R2269 B.n970 B.n108 10.6151
R2270 B.n964 B.n108 10.6151
R2271 B.n964 B.n963 10.6151
R2272 B.n963 B.n962 10.6151
R2273 B.n962 B.n116 10.6151
R2274 B.n956 B.n116 10.6151
R2275 B.n956 B.n955 10.6151
R2276 B.n955 B.n954 10.6151
R2277 B.n954 B.n123 10.6151
R2278 B.n948 B.n123 10.6151
R2279 B.n948 B.n947 10.6151
R2280 B.n947 B.n946 10.6151
R2281 B.n946 B.n130 10.6151
R2282 B.n940 B.n130 10.6151
R2283 B.n940 B.n939 10.6151
R2284 B.n939 B.n938 10.6151
R2285 B.n938 B.n136 10.6151
R2286 B.n932 B.n136 10.6151
R2287 B.n932 B.n931 10.6151
R2288 B.n931 B.n930 10.6151
R2289 B.n930 B.n144 10.6151
R2290 B.n924 B.n144 10.6151
R2291 B.n924 B.n923 10.6151
R2292 B.n923 B.n922 10.6151
R2293 B.n183 B.n151 10.6151
R2294 B.n186 B.n183 10.6151
R2295 B.n187 B.n186 10.6151
R2296 B.n190 B.n187 10.6151
R2297 B.n191 B.n190 10.6151
R2298 B.n194 B.n191 10.6151
R2299 B.n195 B.n194 10.6151
R2300 B.n198 B.n195 10.6151
R2301 B.n199 B.n198 10.6151
R2302 B.n202 B.n199 10.6151
R2303 B.n203 B.n202 10.6151
R2304 B.n206 B.n203 10.6151
R2305 B.n207 B.n206 10.6151
R2306 B.n210 B.n207 10.6151
R2307 B.n211 B.n210 10.6151
R2308 B.n214 B.n211 10.6151
R2309 B.n215 B.n214 10.6151
R2310 B.n219 B.n218 10.6151
R2311 B.n222 B.n219 10.6151
R2312 B.n223 B.n222 10.6151
R2313 B.n226 B.n223 10.6151
R2314 B.n227 B.n226 10.6151
R2315 B.n230 B.n227 10.6151
R2316 B.n231 B.n230 10.6151
R2317 B.n234 B.n231 10.6151
R2318 B.n235 B.n234 10.6151
R2319 B.n239 B.n238 10.6151
R2320 B.n242 B.n239 10.6151
R2321 B.n243 B.n242 10.6151
R2322 B.n246 B.n243 10.6151
R2323 B.n247 B.n246 10.6151
R2324 B.n250 B.n247 10.6151
R2325 B.n251 B.n250 10.6151
R2326 B.n254 B.n251 10.6151
R2327 B.n255 B.n254 10.6151
R2328 B.n258 B.n255 10.6151
R2329 B.n259 B.n258 10.6151
R2330 B.n262 B.n259 10.6151
R2331 B.n263 B.n262 10.6151
R2332 B.n266 B.n263 10.6151
R2333 B.n268 B.n266 10.6151
R2334 B.n269 B.n268 10.6151
R2335 B.n916 B.n269 10.6151
R2336 B.n495 B.n494 9.36635
R2337 B.n519 B.n518 9.36635
R2338 B.n215 B.n182 9.36635
R2339 B.n238 B.n179 9.36635
R2340 B.n1092 B.n0 8.11757
R2341 B.n1092 B.n1 8.11757
R2342 B.n336 B.t9 4.72406
R2343 B.t0 B.n1023 4.72406
R2344 B.n494 B.n451 1.24928
R2345 B.n518 B.n517 1.24928
R2346 B.n218 B.n182 1.24928
R2347 B.n235 B.n179 1.24928
R2348 VP.n34 VP.n33 161.3
R2349 VP.n35 VP.n30 161.3
R2350 VP.n37 VP.n36 161.3
R2351 VP.n38 VP.n29 161.3
R2352 VP.n40 VP.n39 161.3
R2353 VP.n41 VP.n28 161.3
R2354 VP.n43 VP.n42 161.3
R2355 VP.n44 VP.n27 161.3
R2356 VP.n46 VP.n45 161.3
R2357 VP.n48 VP.n26 161.3
R2358 VP.n50 VP.n49 161.3
R2359 VP.n51 VP.n25 161.3
R2360 VP.n53 VP.n52 161.3
R2361 VP.n54 VP.n24 161.3
R2362 VP.n56 VP.n55 161.3
R2363 VP.n57 VP.n23 161.3
R2364 VP.n59 VP.n58 161.3
R2365 VP.n60 VP.n22 161.3
R2366 VP.n63 VP.n62 161.3
R2367 VP.n64 VP.n21 161.3
R2368 VP.n66 VP.n65 161.3
R2369 VP.n67 VP.n20 161.3
R2370 VP.n69 VP.n68 161.3
R2371 VP.n70 VP.n19 161.3
R2372 VP.n72 VP.n71 161.3
R2373 VP.n73 VP.n18 161.3
R2374 VP.n130 VP.n0 161.3
R2375 VP.n129 VP.n128 161.3
R2376 VP.n127 VP.n1 161.3
R2377 VP.n126 VP.n125 161.3
R2378 VP.n124 VP.n2 161.3
R2379 VP.n123 VP.n122 161.3
R2380 VP.n121 VP.n3 161.3
R2381 VP.n120 VP.n119 161.3
R2382 VP.n117 VP.n4 161.3
R2383 VP.n116 VP.n115 161.3
R2384 VP.n114 VP.n5 161.3
R2385 VP.n113 VP.n112 161.3
R2386 VP.n111 VP.n6 161.3
R2387 VP.n110 VP.n109 161.3
R2388 VP.n108 VP.n7 161.3
R2389 VP.n107 VP.n106 161.3
R2390 VP.n105 VP.n8 161.3
R2391 VP.n103 VP.n102 161.3
R2392 VP.n101 VP.n9 161.3
R2393 VP.n100 VP.n99 161.3
R2394 VP.n98 VP.n10 161.3
R2395 VP.n97 VP.n96 161.3
R2396 VP.n95 VP.n11 161.3
R2397 VP.n94 VP.n93 161.3
R2398 VP.n92 VP.n12 161.3
R2399 VP.n91 VP.n90 161.3
R2400 VP.n89 VP.n88 161.3
R2401 VP.n87 VP.n14 161.3
R2402 VP.n86 VP.n85 161.3
R2403 VP.n84 VP.n15 161.3
R2404 VP.n83 VP.n82 161.3
R2405 VP.n81 VP.n16 161.3
R2406 VP.n80 VP.n79 161.3
R2407 VP.n78 VP.n17 161.3
R2408 VP.n32 VP.n31 71.3575
R2409 VP.n77 VP.n76 62.2146
R2410 VP.n132 VP.n131 62.2146
R2411 VP.n75 VP.n74 62.2146
R2412 VP.n32 VP.t0 56.692
R2413 VP.n82 VP.n15 56.5617
R2414 VP.n125 VP.n124 56.5617
R2415 VP.n68 VP.n67 56.5617
R2416 VP.n77 VP.n75 54.9401
R2417 VP.n98 VP.n97 48.8116
R2418 VP.n111 VP.n110 48.8116
R2419 VP.n54 VP.n53 48.8116
R2420 VP.n41 VP.n40 48.8116
R2421 VP.n97 VP.n11 32.3425
R2422 VP.n112 VP.n111 32.3425
R2423 VP.n55 VP.n54 32.3425
R2424 VP.n40 VP.n29 32.3425
R2425 VP.n80 VP.n17 24.5923
R2426 VP.n81 VP.n80 24.5923
R2427 VP.n82 VP.n81 24.5923
R2428 VP.n86 VP.n15 24.5923
R2429 VP.n87 VP.n86 24.5923
R2430 VP.n88 VP.n87 24.5923
R2431 VP.n92 VP.n91 24.5923
R2432 VP.n93 VP.n92 24.5923
R2433 VP.n93 VP.n11 24.5923
R2434 VP.n99 VP.n98 24.5923
R2435 VP.n99 VP.n9 24.5923
R2436 VP.n103 VP.n9 24.5923
R2437 VP.n106 VP.n105 24.5923
R2438 VP.n106 VP.n7 24.5923
R2439 VP.n110 VP.n7 24.5923
R2440 VP.n112 VP.n5 24.5923
R2441 VP.n116 VP.n5 24.5923
R2442 VP.n117 VP.n116 24.5923
R2443 VP.n119 VP.n3 24.5923
R2444 VP.n123 VP.n3 24.5923
R2445 VP.n124 VP.n123 24.5923
R2446 VP.n125 VP.n1 24.5923
R2447 VP.n129 VP.n1 24.5923
R2448 VP.n130 VP.n129 24.5923
R2449 VP.n68 VP.n19 24.5923
R2450 VP.n72 VP.n19 24.5923
R2451 VP.n73 VP.n72 24.5923
R2452 VP.n55 VP.n23 24.5923
R2453 VP.n59 VP.n23 24.5923
R2454 VP.n60 VP.n59 24.5923
R2455 VP.n62 VP.n21 24.5923
R2456 VP.n66 VP.n21 24.5923
R2457 VP.n67 VP.n66 24.5923
R2458 VP.n42 VP.n41 24.5923
R2459 VP.n42 VP.n27 24.5923
R2460 VP.n46 VP.n27 24.5923
R2461 VP.n49 VP.n48 24.5923
R2462 VP.n49 VP.n25 24.5923
R2463 VP.n53 VP.n25 24.5923
R2464 VP.n35 VP.n34 24.5923
R2465 VP.n36 VP.n35 24.5923
R2466 VP.n36 VP.n29 24.5923
R2467 VP.n76 VP.t9 24.3415
R2468 VP.n13 VP.t5 24.3415
R2469 VP.n104 VP.t4 24.3415
R2470 VP.n118 VP.t8 24.3415
R2471 VP.n131 VP.t6 24.3415
R2472 VP.n74 VP.t7 24.3415
R2473 VP.n61 VP.t2 24.3415
R2474 VP.n47 VP.t1 24.3415
R2475 VP.n31 VP.t3 24.3415
R2476 VP.n88 VP.n13 20.6576
R2477 VP.n119 VP.n118 20.6576
R2478 VP.n62 VP.n61 20.6576
R2479 VP.n76 VP.n17 20.1658
R2480 VP.n131 VP.n130 20.1658
R2481 VP.n74 VP.n73 20.1658
R2482 VP.n104 VP.n103 12.2964
R2483 VP.n105 VP.n104 12.2964
R2484 VP.n47 VP.n46 12.2964
R2485 VP.n48 VP.n47 12.2964
R2486 VP.n91 VP.n13 3.93519
R2487 VP.n118 VP.n117 3.93519
R2488 VP.n61 VP.n60 3.93519
R2489 VP.n34 VP.n31 3.93519
R2490 VP.n33 VP.n32 2.68047
R2491 VP.n75 VP.n18 0.417304
R2492 VP.n78 VP.n77 0.417304
R2493 VP.n132 VP.n0 0.417304
R2494 VP VP.n132 0.394524
R2495 VP.n33 VP.n30 0.189894
R2496 VP.n37 VP.n30 0.189894
R2497 VP.n38 VP.n37 0.189894
R2498 VP.n39 VP.n38 0.189894
R2499 VP.n39 VP.n28 0.189894
R2500 VP.n43 VP.n28 0.189894
R2501 VP.n44 VP.n43 0.189894
R2502 VP.n45 VP.n44 0.189894
R2503 VP.n45 VP.n26 0.189894
R2504 VP.n50 VP.n26 0.189894
R2505 VP.n51 VP.n50 0.189894
R2506 VP.n52 VP.n51 0.189894
R2507 VP.n52 VP.n24 0.189894
R2508 VP.n56 VP.n24 0.189894
R2509 VP.n57 VP.n56 0.189894
R2510 VP.n58 VP.n57 0.189894
R2511 VP.n58 VP.n22 0.189894
R2512 VP.n63 VP.n22 0.189894
R2513 VP.n64 VP.n63 0.189894
R2514 VP.n65 VP.n64 0.189894
R2515 VP.n65 VP.n20 0.189894
R2516 VP.n69 VP.n20 0.189894
R2517 VP.n70 VP.n69 0.189894
R2518 VP.n71 VP.n70 0.189894
R2519 VP.n71 VP.n18 0.189894
R2520 VP.n79 VP.n78 0.189894
R2521 VP.n79 VP.n16 0.189894
R2522 VP.n83 VP.n16 0.189894
R2523 VP.n84 VP.n83 0.189894
R2524 VP.n85 VP.n84 0.189894
R2525 VP.n85 VP.n14 0.189894
R2526 VP.n89 VP.n14 0.189894
R2527 VP.n90 VP.n89 0.189894
R2528 VP.n90 VP.n12 0.189894
R2529 VP.n94 VP.n12 0.189894
R2530 VP.n95 VP.n94 0.189894
R2531 VP.n96 VP.n95 0.189894
R2532 VP.n96 VP.n10 0.189894
R2533 VP.n100 VP.n10 0.189894
R2534 VP.n101 VP.n100 0.189894
R2535 VP.n102 VP.n101 0.189894
R2536 VP.n102 VP.n8 0.189894
R2537 VP.n107 VP.n8 0.189894
R2538 VP.n108 VP.n107 0.189894
R2539 VP.n109 VP.n108 0.189894
R2540 VP.n109 VP.n6 0.189894
R2541 VP.n113 VP.n6 0.189894
R2542 VP.n114 VP.n113 0.189894
R2543 VP.n115 VP.n114 0.189894
R2544 VP.n115 VP.n4 0.189894
R2545 VP.n120 VP.n4 0.189894
R2546 VP.n121 VP.n120 0.189894
R2547 VP.n122 VP.n121 0.189894
R2548 VP.n122 VP.n2 0.189894
R2549 VP.n126 VP.n2 0.189894
R2550 VP.n127 VP.n126 0.189894
R2551 VP.n128 VP.n127 0.189894
R2552 VP.n128 VP.n0 0.189894
R2553 VDD1.n14 VDD1.n0 289.615
R2554 VDD1.n35 VDD1.n21 289.615
R2555 VDD1.n15 VDD1.n14 185
R2556 VDD1.n13 VDD1.n12 185
R2557 VDD1.n4 VDD1.n3 185
R2558 VDD1.n7 VDD1.n6 185
R2559 VDD1.n28 VDD1.n27 185
R2560 VDD1.n25 VDD1.n24 185
R2561 VDD1.n34 VDD1.n33 185
R2562 VDD1.n36 VDD1.n35 185
R2563 VDD1.t9 VDD1.n5 147.888
R2564 VDD1.t0 VDD1.n26 147.888
R2565 VDD1.n14 VDD1.n13 104.615
R2566 VDD1.n13 VDD1.n3 104.615
R2567 VDD1.n6 VDD1.n3 104.615
R2568 VDD1.n27 VDD1.n24 104.615
R2569 VDD1.n34 VDD1.n24 104.615
R2570 VDD1.n35 VDD1.n34 104.615
R2571 VDD1.n43 VDD1.n42 80.087
R2572 VDD1.n20 VDD1.n19 77.3429
R2573 VDD1.n45 VDD1.n44 77.3428
R2574 VDD1.n41 VDD1.n40 77.3428
R2575 VDD1.n20 VDD1.n18 56.4757
R2576 VDD1.n41 VDD1.n39 56.4757
R2577 VDD1.n6 VDD1.t9 52.3082
R2578 VDD1.n27 VDD1.t0 52.3082
R2579 VDD1.n45 VDD1.n43 47.378
R2580 VDD1.n7 VDD1.n5 15.6496
R2581 VDD1.n28 VDD1.n26 15.6496
R2582 VDD1.n8 VDD1.n4 12.8005
R2583 VDD1.n29 VDD1.n25 12.8005
R2584 VDD1.n12 VDD1.n11 12.0247
R2585 VDD1.n33 VDD1.n32 12.0247
R2586 VDD1.n15 VDD1.n2 11.249
R2587 VDD1.n36 VDD1.n23 11.249
R2588 VDD1.n16 VDD1.n0 10.4732
R2589 VDD1.n37 VDD1.n21 10.4732
R2590 VDD1.n18 VDD1.n17 9.45567
R2591 VDD1.n39 VDD1.n38 9.45567
R2592 VDD1.n17 VDD1.n16 9.3005
R2593 VDD1.n2 VDD1.n1 9.3005
R2594 VDD1.n11 VDD1.n10 9.3005
R2595 VDD1.n9 VDD1.n8 9.3005
R2596 VDD1.n38 VDD1.n37 9.3005
R2597 VDD1.n23 VDD1.n22 9.3005
R2598 VDD1.n32 VDD1.n31 9.3005
R2599 VDD1.n30 VDD1.n29 9.3005
R2600 VDD1.n44 VDD1.t7 4.90149
R2601 VDD1.n44 VDD1.t2 4.90149
R2602 VDD1.n19 VDD1.t6 4.90149
R2603 VDD1.n19 VDD1.t8 4.90149
R2604 VDD1.n42 VDD1.t1 4.90149
R2605 VDD1.n42 VDD1.t3 4.90149
R2606 VDD1.n40 VDD1.t4 4.90149
R2607 VDD1.n40 VDD1.t5 4.90149
R2608 VDD1.n9 VDD1.n5 4.40546
R2609 VDD1.n30 VDD1.n26 4.40546
R2610 VDD1.n18 VDD1.n0 3.49141
R2611 VDD1.n39 VDD1.n21 3.49141
R2612 VDD1 VDD1.n45 2.74188
R2613 VDD1.n16 VDD1.n15 2.71565
R2614 VDD1.n37 VDD1.n36 2.71565
R2615 VDD1.n12 VDD1.n2 1.93989
R2616 VDD1.n33 VDD1.n23 1.93989
R2617 VDD1.n11 VDD1.n4 1.16414
R2618 VDD1.n32 VDD1.n25 1.16414
R2619 VDD1 VDD1.n20 0.991879
R2620 VDD1.n43 VDD1.n41 0.878344
R2621 VDD1.n8 VDD1.n7 0.388379
R2622 VDD1.n29 VDD1.n28 0.388379
R2623 VDD1.n17 VDD1.n1 0.155672
R2624 VDD1.n10 VDD1.n1 0.155672
R2625 VDD1.n10 VDD1.n9 0.155672
R2626 VDD1.n31 VDD1.n30 0.155672
R2627 VDD1.n31 VDD1.n22 0.155672
R2628 VDD1.n38 VDD1.n22 0.155672
C0 VDD1 VN 0.161223f
C1 VDD1 VP 4.83061f
C2 VDD2 VN 4.22875f
C3 VDD2 VP 0.767091f
C4 VDD1 VTAIL 8.14611f
C5 VDD2 VTAIL 8.208679f
C6 VP VN 8.98743f
C7 VN VTAIL 6.20511f
C8 VP VTAIL 6.219471f
C9 VDD1 VDD2 3.08629f
C10 VDD2 B 7.56508f
C11 VDD1 B 7.449311f
C12 VTAIL B 5.350293f
C13 VN B 24.09261f
C14 VP B 22.533785f
C15 VDD1.n0 B 0.042457f
C16 VDD1.n1 B 0.029088f
C17 VDD1.n2 B 0.015631f
C18 VDD1.n3 B 0.036946f
C19 VDD1.n4 B 0.01655f
C20 VDD1.n5 B 0.113091f
C21 VDD1.t9 B 0.061636f
C22 VDD1.n6 B 0.027709f
C23 VDD1.n7 B 0.021745f
C24 VDD1.n8 B 0.015631f
C25 VDD1.n9 B 0.426397f
C26 VDD1.n10 B 0.029088f
C27 VDD1.n11 B 0.015631f
C28 VDD1.n12 B 0.01655f
C29 VDD1.n13 B 0.036946f
C30 VDD1.n14 B 0.082758f
C31 VDD1.n15 B 0.01655f
C32 VDD1.n16 B 0.015631f
C33 VDD1.n17 B 0.075184f
C34 VDD1.n18 B 0.093982f
C35 VDD1.t6 B 0.092866f
C36 VDD1.t8 B 0.092866f
C37 VDD1.n19 B 0.730037f
C38 VDD1.n20 B 1.05371f
C39 VDD1.n21 B 0.042457f
C40 VDD1.n22 B 0.029088f
C41 VDD1.n23 B 0.015631f
C42 VDD1.n24 B 0.036946f
C43 VDD1.n25 B 0.01655f
C44 VDD1.n26 B 0.113091f
C45 VDD1.t0 B 0.061636f
C46 VDD1.n27 B 0.027709f
C47 VDD1.n28 B 0.021745f
C48 VDD1.n29 B 0.015631f
C49 VDD1.n30 B 0.426397f
C50 VDD1.n31 B 0.029088f
C51 VDD1.n32 B 0.015631f
C52 VDD1.n33 B 0.01655f
C53 VDD1.n34 B 0.036946f
C54 VDD1.n35 B 0.082758f
C55 VDD1.n36 B 0.01655f
C56 VDD1.n37 B 0.015631f
C57 VDD1.n38 B 0.075184f
C58 VDD1.n39 B 0.093982f
C59 VDD1.t4 B 0.092866f
C60 VDD1.t5 B 0.092866f
C61 VDD1.n40 B 0.730034f
C62 VDD1.n41 B 1.04384f
C63 VDD1.t1 B 0.092866f
C64 VDD1.t3 B 0.092866f
C65 VDD1.n42 B 0.759045f
C66 VDD1.n43 B 3.83449f
C67 VDD1.t7 B 0.092866f
C68 VDD1.t2 B 0.092866f
C69 VDD1.n44 B 0.730034f
C70 VDD1.n45 B 3.6476f
C71 VP.n0 B 0.040708f
C72 VP.t6 B 0.899504f
C73 VP.n1 B 0.040144f
C74 VP.n2 B 0.021648f
C75 VP.n3 B 0.040144f
C76 VP.n4 B 0.021648f
C77 VP.t8 B 0.899504f
C78 VP.n5 B 0.040144f
C79 VP.n6 B 0.021648f
C80 VP.n7 B 0.040144f
C81 VP.n8 B 0.021648f
C82 VP.t4 B 0.899504f
C83 VP.n9 B 0.040144f
C84 VP.n10 B 0.021648f
C85 VP.n11 B 0.043374f
C86 VP.n12 B 0.021648f
C87 VP.t5 B 0.899504f
C88 VP.n13 B 0.346617f
C89 VP.n14 B 0.021648f
C90 VP.n15 B 0.031169f
C91 VP.n16 B 0.021648f
C92 VP.n17 B 0.036577f
C93 VP.n18 B 0.040708f
C94 VP.t7 B 0.899504f
C95 VP.n19 B 0.040144f
C96 VP.n20 B 0.021648f
C97 VP.n21 B 0.040144f
C98 VP.n22 B 0.021648f
C99 VP.t2 B 0.899504f
C100 VP.n23 B 0.040144f
C101 VP.n24 B 0.021648f
C102 VP.n25 B 0.040144f
C103 VP.n26 B 0.021648f
C104 VP.t1 B 0.899504f
C105 VP.n27 B 0.040144f
C106 VP.n28 B 0.021648f
C107 VP.n29 B 0.043374f
C108 VP.n30 B 0.021648f
C109 VP.t3 B 0.899504f
C110 VP.n31 B 0.418992f
C111 VP.t0 B 1.19448f
C112 VP.n32 B 0.429623f
C113 VP.n33 B 0.289413f
C114 VP.n34 B 0.023497f
C115 VP.n35 B 0.040144f
C116 VP.n36 B 0.040144f
C117 VP.n37 B 0.021648f
C118 VP.n38 B 0.021648f
C119 VP.n39 B 0.021648f
C120 VP.n40 B 0.019564f
C121 VP.n41 B 0.040144f
C122 VP.n42 B 0.040144f
C123 VP.n43 B 0.021648f
C124 VP.n44 B 0.021648f
C125 VP.n45 B 0.021648f
C126 VP.n46 B 0.030235f
C127 VP.n47 B 0.346617f
C128 VP.n48 B 0.030235f
C129 VP.n49 B 0.040144f
C130 VP.n50 B 0.021648f
C131 VP.n51 B 0.021648f
C132 VP.n52 B 0.021648f
C133 VP.n53 B 0.040144f
C134 VP.n54 B 0.019564f
C135 VP.n55 B 0.043374f
C136 VP.n56 B 0.021648f
C137 VP.n57 B 0.021648f
C138 VP.n58 B 0.021648f
C139 VP.n59 B 0.040144f
C140 VP.n60 B 0.023497f
C141 VP.n61 B 0.346617f
C142 VP.n62 B 0.036973f
C143 VP.n63 B 0.021648f
C144 VP.n64 B 0.021648f
C145 VP.n65 B 0.021648f
C146 VP.n66 B 0.040144f
C147 VP.n67 B 0.031169f
C148 VP.n68 B 0.031768f
C149 VP.n69 B 0.021648f
C150 VP.n70 B 0.021648f
C151 VP.n71 B 0.021648f
C152 VP.n72 B 0.040144f
C153 VP.n73 B 0.036577f
C154 VP.n74 B 0.441156f
C155 VP.n75 B 1.43587f
C156 VP.t9 B 0.899504f
C157 VP.n76 B 0.441156f
C158 VP.n77 B 1.45008f
C159 VP.n78 B 0.040708f
C160 VP.n79 B 0.021648f
C161 VP.n80 B 0.040144f
C162 VP.n81 B 0.040144f
C163 VP.n82 B 0.031768f
C164 VP.n83 B 0.021648f
C165 VP.n84 B 0.021648f
C166 VP.n85 B 0.021648f
C167 VP.n86 B 0.040144f
C168 VP.n87 B 0.040144f
C169 VP.n88 B 0.036973f
C170 VP.n89 B 0.021648f
C171 VP.n90 B 0.021648f
C172 VP.n91 B 0.023497f
C173 VP.n92 B 0.040144f
C174 VP.n93 B 0.040144f
C175 VP.n94 B 0.021648f
C176 VP.n95 B 0.021648f
C177 VP.n96 B 0.021648f
C178 VP.n97 B 0.019564f
C179 VP.n98 B 0.040144f
C180 VP.n99 B 0.040144f
C181 VP.n100 B 0.021648f
C182 VP.n101 B 0.021648f
C183 VP.n102 B 0.021648f
C184 VP.n103 B 0.030235f
C185 VP.n104 B 0.346617f
C186 VP.n105 B 0.030235f
C187 VP.n106 B 0.040144f
C188 VP.n107 B 0.021648f
C189 VP.n108 B 0.021648f
C190 VP.n109 B 0.021648f
C191 VP.n110 B 0.040144f
C192 VP.n111 B 0.019564f
C193 VP.n112 B 0.043374f
C194 VP.n113 B 0.021648f
C195 VP.n114 B 0.021648f
C196 VP.n115 B 0.021648f
C197 VP.n116 B 0.040144f
C198 VP.n117 B 0.023497f
C199 VP.n118 B 0.346617f
C200 VP.n119 B 0.036973f
C201 VP.n120 B 0.021648f
C202 VP.n121 B 0.021648f
C203 VP.n122 B 0.021648f
C204 VP.n123 B 0.040144f
C205 VP.n124 B 0.031169f
C206 VP.n125 B 0.031768f
C207 VP.n126 B 0.021648f
C208 VP.n127 B 0.021648f
C209 VP.n128 B 0.021648f
C210 VP.n129 B 0.040144f
C211 VP.n130 B 0.036577f
C212 VP.n131 B 0.441156f
C213 VP.n132 B 0.069389f
C214 VDD2.n0 B 0.041408f
C215 VDD2.n1 B 0.02837f
C216 VDD2.n2 B 0.015245f
C217 VDD2.n3 B 0.036033f
C218 VDD2.n4 B 0.016142f
C219 VDD2.n5 B 0.110297f
C220 VDD2.t8 B 0.060113f
C221 VDD2.n6 B 0.027025f
C222 VDD2.n7 B 0.021208f
C223 VDD2.n8 B 0.015245f
C224 VDD2.n9 B 0.415864f
C225 VDD2.n10 B 0.02837f
C226 VDD2.n11 B 0.015245f
C227 VDD2.n12 B 0.016142f
C228 VDD2.n13 B 0.036033f
C229 VDD2.n14 B 0.080714f
C230 VDD2.n15 B 0.016142f
C231 VDD2.n16 B 0.015245f
C232 VDD2.n17 B 0.073327f
C233 VDD2.n18 B 0.09166f
C234 VDD2.t2 B 0.090572f
C235 VDD2.t9 B 0.090572f
C236 VDD2.n19 B 0.712001f
C237 VDD2.n20 B 1.01806f
C238 VDD2.t3 B 0.090572f
C239 VDD2.t4 B 0.090572f
C240 VDD2.n21 B 0.740296f
C241 VDD2.n22 B 3.56278f
C242 VDD2.n23 B 0.041408f
C243 VDD2.n24 B 0.02837f
C244 VDD2.n25 B 0.015245f
C245 VDD2.n26 B 0.036033f
C246 VDD2.n27 B 0.016142f
C247 VDD2.n28 B 0.110297f
C248 VDD2.t1 B 0.060113f
C249 VDD2.n29 B 0.027025f
C250 VDD2.n30 B 0.021208f
C251 VDD2.n31 B 0.015245f
C252 VDD2.n32 B 0.415864f
C253 VDD2.n33 B 0.02837f
C254 VDD2.n34 B 0.015245f
C255 VDD2.n35 B 0.016142f
C256 VDD2.n36 B 0.036033f
C257 VDD2.n37 B 0.080714f
C258 VDD2.n38 B 0.016142f
C259 VDD2.n39 B 0.015245f
C260 VDD2.n40 B 0.073327f
C261 VDD2.n41 B 0.065203f
C262 VDD2.n42 B 3.20476f
C263 VDD2.t5 B 0.090572f
C264 VDD2.t6 B 0.090572f
C265 VDD2.n43 B 0.712004f
C266 VDD2.n44 B 0.653847f
C267 VDD2.t7 B 0.090572f
C268 VDD2.t0 B 0.090572f
C269 VDD2.n45 B 0.740251f
C270 VTAIL.t13 B 0.106714f
C271 VTAIL.t9 B 0.106714f
C272 VTAIL.n0 B 0.768733f
C273 VTAIL.n1 B 0.845715f
C274 VTAIL.n2 B 0.048788f
C275 VTAIL.n3 B 0.033426f
C276 VTAIL.n4 B 0.017962f
C277 VTAIL.n5 B 0.042455f
C278 VTAIL.n6 B 0.019018f
C279 VTAIL.n7 B 0.129955f
C280 VTAIL.t4 B 0.070827f
C281 VTAIL.n8 B 0.031841f
C282 VTAIL.n9 B 0.024987f
C283 VTAIL.n10 B 0.017962f
C284 VTAIL.n11 B 0.489981f
C285 VTAIL.n12 B 0.033426f
C286 VTAIL.n13 B 0.017962f
C287 VTAIL.n14 B 0.019018f
C288 VTAIL.n15 B 0.042455f
C289 VTAIL.n16 B 0.095099f
C290 VTAIL.n17 B 0.019018f
C291 VTAIL.n18 B 0.017962f
C292 VTAIL.n19 B 0.086396f
C293 VTAIL.n20 B 0.053806f
C294 VTAIL.n21 B 0.687385f
C295 VTAIL.t19 B 0.106714f
C296 VTAIL.t6 B 0.106714f
C297 VTAIL.n22 B 0.768733f
C298 VTAIL.n23 B 1.09038f
C299 VTAIL.t5 B 0.106714f
C300 VTAIL.t2 B 0.106714f
C301 VTAIL.n24 B 0.768733f
C302 VTAIL.n25 B 2.32159f
C303 VTAIL.t15 B 0.106714f
C304 VTAIL.t17 B 0.106714f
C305 VTAIL.n26 B 0.768738f
C306 VTAIL.n27 B 2.32159f
C307 VTAIL.t16 B 0.106714f
C308 VTAIL.t14 B 0.106714f
C309 VTAIL.n28 B 0.768738f
C310 VTAIL.n29 B 1.09037f
C311 VTAIL.n30 B 0.048788f
C312 VTAIL.n31 B 0.033426f
C313 VTAIL.n32 B 0.017962f
C314 VTAIL.n33 B 0.042455f
C315 VTAIL.n34 B 0.019018f
C316 VTAIL.n35 B 0.129955f
C317 VTAIL.t11 B 0.070827f
C318 VTAIL.n36 B 0.031841f
C319 VTAIL.n37 B 0.024987f
C320 VTAIL.n38 B 0.017962f
C321 VTAIL.n39 B 0.489981f
C322 VTAIL.n40 B 0.033426f
C323 VTAIL.n41 B 0.017962f
C324 VTAIL.n42 B 0.019018f
C325 VTAIL.n43 B 0.042455f
C326 VTAIL.n44 B 0.095099f
C327 VTAIL.n45 B 0.019018f
C328 VTAIL.n46 B 0.017962f
C329 VTAIL.n47 B 0.086396f
C330 VTAIL.n48 B 0.053806f
C331 VTAIL.n49 B 0.687385f
C332 VTAIL.t3 B 0.106714f
C333 VTAIL.t7 B 0.106714f
C334 VTAIL.n50 B 0.768738f
C335 VTAIL.n51 B 0.939954f
C336 VTAIL.t0 B 0.106714f
C337 VTAIL.t8 B 0.106714f
C338 VTAIL.n52 B 0.768738f
C339 VTAIL.n53 B 1.09037f
C340 VTAIL.n54 B 0.048788f
C341 VTAIL.n55 B 0.033426f
C342 VTAIL.n56 B 0.017962f
C343 VTAIL.n57 B 0.042455f
C344 VTAIL.n58 B 0.019018f
C345 VTAIL.n59 B 0.129955f
C346 VTAIL.t1 B 0.070827f
C347 VTAIL.n60 B 0.031841f
C348 VTAIL.n61 B 0.024987f
C349 VTAIL.n62 B 0.017962f
C350 VTAIL.n63 B 0.489981f
C351 VTAIL.n64 B 0.033426f
C352 VTAIL.n65 B 0.017962f
C353 VTAIL.n66 B 0.019018f
C354 VTAIL.n67 B 0.042455f
C355 VTAIL.n68 B 0.095099f
C356 VTAIL.n69 B 0.019018f
C357 VTAIL.n70 B 0.017962f
C358 VTAIL.n71 B 0.086396f
C359 VTAIL.n72 B 0.053806f
C360 VTAIL.n73 B 1.66697f
C361 VTAIL.n74 B 0.048788f
C362 VTAIL.n75 B 0.033426f
C363 VTAIL.n76 B 0.017962f
C364 VTAIL.n77 B 0.042455f
C365 VTAIL.n78 B 0.019018f
C366 VTAIL.n79 B 0.129955f
C367 VTAIL.t12 B 0.070827f
C368 VTAIL.n80 B 0.031841f
C369 VTAIL.n81 B 0.024987f
C370 VTAIL.n82 B 0.017962f
C371 VTAIL.n83 B 0.489981f
C372 VTAIL.n84 B 0.033426f
C373 VTAIL.n85 B 0.017962f
C374 VTAIL.n86 B 0.019018f
C375 VTAIL.n87 B 0.042455f
C376 VTAIL.n88 B 0.095099f
C377 VTAIL.n89 B 0.019018f
C378 VTAIL.n90 B 0.017962f
C379 VTAIL.n91 B 0.086396f
C380 VTAIL.n92 B 0.053806f
C381 VTAIL.n93 B 1.66697f
C382 VTAIL.t18 B 0.106714f
C383 VTAIL.t10 B 0.106714f
C384 VTAIL.n94 B 0.768733f
C385 VTAIL.n95 B 0.782577f
C386 VN.n0 B 0.039427f
C387 VN.t5 B 0.871194f
C388 VN.n1 B 0.038881f
C389 VN.n2 B 0.020967f
C390 VN.n3 B 0.038881f
C391 VN.n4 B 0.020967f
C392 VN.t6 B 0.871194f
C393 VN.n5 B 0.038881f
C394 VN.n6 B 0.020967f
C395 VN.n7 B 0.038881f
C396 VN.n8 B 0.020967f
C397 VN.t0 B 0.871194f
C398 VN.n9 B 0.038881f
C399 VN.n10 B 0.020967f
C400 VN.n11 B 0.042009f
C401 VN.n12 B 0.020967f
C402 VN.t7 B 0.871194f
C403 VN.n13 B 0.405805f
C404 VN.t1 B 1.15689f
C405 VN.n14 B 0.4161f
C406 VN.n15 B 0.280303f
C407 VN.n16 B 0.022757f
C408 VN.n17 B 0.038881f
C409 VN.n18 B 0.038881f
C410 VN.n19 B 0.020967f
C411 VN.n20 B 0.020967f
C412 VN.n21 B 0.020967f
C413 VN.n22 B 0.018948f
C414 VN.n23 B 0.038881f
C415 VN.n24 B 0.038881f
C416 VN.n25 B 0.020967f
C417 VN.n26 B 0.020967f
C418 VN.n27 B 0.020967f
C419 VN.n28 B 0.029284f
C420 VN.n29 B 0.335707f
C421 VN.n30 B 0.029284f
C422 VN.n31 B 0.038881f
C423 VN.n32 B 0.020967f
C424 VN.n33 B 0.020967f
C425 VN.n34 B 0.020967f
C426 VN.n35 B 0.038881f
C427 VN.n36 B 0.018948f
C428 VN.n37 B 0.042009f
C429 VN.n38 B 0.020967f
C430 VN.n39 B 0.020967f
C431 VN.n40 B 0.020967f
C432 VN.n41 B 0.038881f
C433 VN.n42 B 0.022757f
C434 VN.n43 B 0.335707f
C435 VN.n44 B 0.03581f
C436 VN.n45 B 0.020967f
C437 VN.n46 B 0.020967f
C438 VN.n47 B 0.020967f
C439 VN.n48 B 0.038881f
C440 VN.n49 B 0.030188f
C441 VN.n50 B 0.030768f
C442 VN.n51 B 0.020967f
C443 VN.n52 B 0.020967f
C444 VN.n53 B 0.020967f
C445 VN.n54 B 0.038881f
C446 VN.n55 B 0.035426f
C447 VN.n56 B 0.427271f
C448 VN.n57 B 0.067205f
C449 VN.n58 B 0.039427f
C450 VN.t8 B 0.871194f
C451 VN.n59 B 0.038881f
C452 VN.n60 B 0.020967f
C453 VN.n61 B 0.038881f
C454 VN.n62 B 0.020967f
C455 VN.t4 B 0.871194f
C456 VN.n63 B 0.038881f
C457 VN.n64 B 0.020967f
C458 VN.n65 B 0.038881f
C459 VN.n66 B 0.020967f
C460 VN.t3 B 0.871194f
C461 VN.n67 B 0.038881f
C462 VN.n68 B 0.020967f
C463 VN.n69 B 0.042009f
C464 VN.n70 B 0.020967f
C465 VN.t2 B 0.871194f
C466 VN.n71 B 0.405805f
C467 VN.t9 B 1.15689f
C468 VN.n72 B 0.4161f
C469 VN.n73 B 0.280303f
C470 VN.n74 B 0.022757f
C471 VN.n75 B 0.038881f
C472 VN.n76 B 0.038881f
C473 VN.n77 B 0.020967f
C474 VN.n78 B 0.020967f
C475 VN.n79 B 0.020967f
C476 VN.n80 B 0.018948f
C477 VN.n81 B 0.038881f
C478 VN.n82 B 0.038881f
C479 VN.n83 B 0.020967f
C480 VN.n84 B 0.020967f
C481 VN.n85 B 0.020967f
C482 VN.n86 B 0.029284f
C483 VN.n87 B 0.335707f
C484 VN.n88 B 0.029284f
C485 VN.n89 B 0.038881f
C486 VN.n90 B 0.020967f
C487 VN.n91 B 0.020967f
C488 VN.n92 B 0.020967f
C489 VN.n93 B 0.038881f
C490 VN.n94 B 0.018948f
C491 VN.n95 B 0.042009f
C492 VN.n96 B 0.020967f
C493 VN.n97 B 0.020967f
C494 VN.n98 B 0.020967f
C495 VN.n99 B 0.038881f
C496 VN.n100 B 0.022757f
C497 VN.n101 B 0.335707f
C498 VN.n102 B 0.03581f
C499 VN.n103 B 0.020967f
C500 VN.n104 B 0.020967f
C501 VN.n105 B 0.020967f
C502 VN.n106 B 0.038881f
C503 VN.n107 B 0.030188f
C504 VN.n108 B 0.030768f
C505 VN.n109 B 0.020967f
C506 VN.n110 B 0.020967f
C507 VN.n111 B 0.020967f
C508 VN.n112 B 0.038881f
C509 VN.n113 B 0.035426f
C510 VN.n114 B 0.427271f
C511 VN.n115 B 1.39578f
.ends

