* NGSPICE file created from diff_pair_sample_1307.ext - technology: sky130A

.subckt diff_pair_sample_1307 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t18 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=2.35785 pd=14.62 as=2.35785 ps=14.62 w=14.29 l=4
X1 VDD1.t9 VP.t0 VTAIL.t1 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=2.35785 pd=14.62 as=2.35785 ps=14.62 w=14.29 l=4
X2 VTAIL.t13 VN.t1 VDD2.t8 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=2.35785 pd=14.62 as=2.35785 ps=14.62 w=14.29 l=4
X3 VTAIL.t2 VP.t1 VDD1.t8 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=2.35785 pd=14.62 as=2.35785 ps=14.62 w=14.29 l=4
X4 VTAIL.t4 VP.t2 VDD1.t7 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=2.35785 pd=14.62 as=2.35785 ps=14.62 w=14.29 l=4
X5 VDD2.t7 VN.t2 VTAIL.t12 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=2.35785 pd=14.62 as=2.35785 ps=14.62 w=14.29 l=4
X6 VDD2.t6 VN.t3 VTAIL.t19 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=5.5731 pd=29.36 as=2.35785 ps=14.62 w=14.29 l=4
X7 VDD2.t5 VN.t4 VTAIL.t16 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=5.5731 pd=29.36 as=2.35785 ps=14.62 w=14.29 l=4
X8 VDD1.t6 VP.t3 VTAIL.t3 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=2.35785 pd=14.62 as=5.5731 ps=29.36 w=14.29 l=4
X9 B.t11 B.t9 B.t10 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=5.5731 pd=29.36 as=0 ps=0 w=14.29 l=4
X10 VDD2.t4 VN.t5 VTAIL.t11 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=2.35785 pd=14.62 as=5.5731 ps=29.36 w=14.29 l=4
X11 B.t8 B.t6 B.t7 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=5.5731 pd=29.36 as=0 ps=0 w=14.29 l=4
X12 VDD2.t3 VN.t6 VTAIL.t17 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=2.35785 pd=14.62 as=5.5731 ps=29.36 w=14.29 l=4
X13 VTAIL.t14 VN.t7 VDD2.t2 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=2.35785 pd=14.62 as=2.35785 ps=14.62 w=14.29 l=4
X14 VTAIL.t15 VN.t8 VDD2.t1 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=2.35785 pd=14.62 as=2.35785 ps=14.62 w=14.29 l=4
X15 B.t5 B.t3 B.t4 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=5.5731 pd=29.36 as=0 ps=0 w=14.29 l=4
X16 VDD1.t5 VP.t4 VTAIL.t7 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=2.35785 pd=14.62 as=2.35785 ps=14.62 w=14.29 l=4
X17 VTAIL.t5 VP.t5 VDD1.t4 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=2.35785 pd=14.62 as=2.35785 ps=14.62 w=14.29 l=4
X18 VDD1.t3 VP.t6 VTAIL.t9 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=2.35785 pd=14.62 as=5.5731 ps=29.36 w=14.29 l=4
X19 B.t2 B.t0 B.t1 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=5.5731 pd=29.36 as=0 ps=0 w=14.29 l=4
X20 VTAIL.t0 VP.t7 VDD1.t2 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=2.35785 pd=14.62 as=2.35785 ps=14.62 w=14.29 l=4
X21 VDD1.t1 VP.t8 VTAIL.t6 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=5.5731 pd=29.36 as=2.35785 ps=14.62 w=14.29 l=4
X22 VDD1.t0 VP.t9 VTAIL.t8 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=5.5731 pd=29.36 as=2.35785 ps=14.62 w=14.29 l=4
X23 VTAIL.t10 VN.t9 VDD2.t0 w_n6166_n3826# sky130_fd_pr__pfet_01v8 ad=2.35785 pd=14.62 as=2.35785 ps=14.62 w=14.29 l=4
R0 VN.n113 VN.n58 161.3
R1 VN.n112 VN.n111 161.3
R2 VN.n110 VN.n59 161.3
R3 VN.n109 VN.n108 161.3
R4 VN.n107 VN.n60 161.3
R5 VN.n106 VN.n105 161.3
R6 VN.n104 VN.n61 161.3
R7 VN.n103 VN.n102 161.3
R8 VN.n100 VN.n62 161.3
R9 VN.n99 VN.n98 161.3
R10 VN.n97 VN.n63 161.3
R11 VN.n96 VN.n95 161.3
R12 VN.n94 VN.n64 161.3
R13 VN.n93 VN.n92 161.3
R14 VN.n91 VN.n65 161.3
R15 VN.n90 VN.n89 161.3
R16 VN.n88 VN.n66 161.3
R17 VN.n86 VN.n85 161.3
R18 VN.n84 VN.n67 161.3
R19 VN.n83 VN.n82 161.3
R20 VN.n81 VN.n68 161.3
R21 VN.n80 VN.n79 161.3
R22 VN.n78 VN.n69 161.3
R23 VN.n77 VN.n76 161.3
R24 VN.n75 VN.n70 161.3
R25 VN.n74 VN.n73 161.3
R26 VN.n55 VN.n0 161.3
R27 VN.n54 VN.n53 161.3
R28 VN.n52 VN.n1 161.3
R29 VN.n51 VN.n50 161.3
R30 VN.n49 VN.n2 161.3
R31 VN.n48 VN.n47 161.3
R32 VN.n46 VN.n3 161.3
R33 VN.n45 VN.n44 161.3
R34 VN.n42 VN.n4 161.3
R35 VN.n41 VN.n40 161.3
R36 VN.n39 VN.n5 161.3
R37 VN.n38 VN.n37 161.3
R38 VN.n36 VN.n6 161.3
R39 VN.n35 VN.n34 161.3
R40 VN.n33 VN.n7 161.3
R41 VN.n32 VN.n31 161.3
R42 VN.n30 VN.n8 161.3
R43 VN.n28 VN.n27 161.3
R44 VN.n26 VN.n9 161.3
R45 VN.n25 VN.n24 161.3
R46 VN.n23 VN.n10 161.3
R47 VN.n22 VN.n21 161.3
R48 VN.n20 VN.n11 161.3
R49 VN.n19 VN.n18 161.3
R50 VN.n17 VN.n12 161.3
R51 VN.n16 VN.n15 161.3
R52 VN.n14 VN.t4 118.368
R53 VN.n72 VN.t5 118.368
R54 VN.n13 VN.t8 86.0978
R55 VN.n29 VN.t2 86.0978
R56 VN.n43 VN.t7 86.0978
R57 VN.n56 VN.t6 86.0978
R58 VN.n71 VN.t9 86.0978
R59 VN.n87 VN.t0 86.0978
R60 VN.n101 VN.t1 86.0978
R61 VN.n114 VN.t3 86.0978
R62 VN.n14 VN.n13 71.1462
R63 VN.n72 VN.n71 71.1462
R64 VN VN.n115 62.7428
R65 VN.n57 VN.n56 62.1188
R66 VN.n115 VN.n114 62.1188
R67 VN.n50 VN.n49 56.5193
R68 VN.n108 VN.n107 56.5193
R69 VN.n23 VN.n22 48.7492
R70 VN.n36 VN.n35 48.7492
R71 VN.n81 VN.n80 48.7492
R72 VN.n94 VN.n93 48.7492
R73 VN.n22 VN.n11 32.2376
R74 VN.n37 VN.n36 32.2376
R75 VN.n80 VN.n69 32.2376
R76 VN.n95 VN.n94 32.2376
R77 VN.n17 VN.n16 24.4675
R78 VN.n18 VN.n17 24.4675
R79 VN.n18 VN.n11 24.4675
R80 VN.n24 VN.n23 24.4675
R81 VN.n24 VN.n9 24.4675
R82 VN.n28 VN.n9 24.4675
R83 VN.n31 VN.n30 24.4675
R84 VN.n31 VN.n7 24.4675
R85 VN.n35 VN.n7 24.4675
R86 VN.n37 VN.n5 24.4675
R87 VN.n41 VN.n5 24.4675
R88 VN.n42 VN.n41 24.4675
R89 VN.n44 VN.n3 24.4675
R90 VN.n48 VN.n3 24.4675
R91 VN.n49 VN.n48 24.4675
R92 VN.n50 VN.n1 24.4675
R93 VN.n54 VN.n1 24.4675
R94 VN.n55 VN.n54 24.4675
R95 VN.n76 VN.n69 24.4675
R96 VN.n76 VN.n75 24.4675
R97 VN.n75 VN.n74 24.4675
R98 VN.n93 VN.n65 24.4675
R99 VN.n89 VN.n65 24.4675
R100 VN.n89 VN.n88 24.4675
R101 VN.n86 VN.n67 24.4675
R102 VN.n82 VN.n67 24.4675
R103 VN.n82 VN.n81 24.4675
R104 VN.n107 VN.n106 24.4675
R105 VN.n106 VN.n61 24.4675
R106 VN.n102 VN.n61 24.4675
R107 VN.n100 VN.n99 24.4675
R108 VN.n99 VN.n63 24.4675
R109 VN.n95 VN.n63 24.4675
R110 VN.n113 VN.n112 24.4675
R111 VN.n112 VN.n59 24.4675
R112 VN.n108 VN.n59 24.4675
R113 VN.n44 VN.n43 20.5528
R114 VN.n102 VN.n101 20.5528
R115 VN.n56 VN.n55 20.0634
R116 VN.n114 VN.n113 20.0634
R117 VN.n29 VN.n28 12.234
R118 VN.n30 VN.n29 12.234
R119 VN.n88 VN.n87 12.234
R120 VN.n87 VN.n86 12.234
R121 VN.n16 VN.n13 3.91522
R122 VN.n43 VN.n42 3.91522
R123 VN.n74 VN.n71 3.91522
R124 VN.n101 VN.n100 3.91522
R125 VN.n73 VN.n72 2.69184
R126 VN.n15 VN.n14 2.69184
R127 VN.n115 VN.n58 0.417535
R128 VN.n57 VN.n0 0.417535
R129 VN VN.n57 0.394291
R130 VN.n111 VN.n58 0.189894
R131 VN.n111 VN.n110 0.189894
R132 VN.n110 VN.n109 0.189894
R133 VN.n109 VN.n60 0.189894
R134 VN.n105 VN.n60 0.189894
R135 VN.n105 VN.n104 0.189894
R136 VN.n104 VN.n103 0.189894
R137 VN.n103 VN.n62 0.189894
R138 VN.n98 VN.n62 0.189894
R139 VN.n98 VN.n97 0.189894
R140 VN.n97 VN.n96 0.189894
R141 VN.n96 VN.n64 0.189894
R142 VN.n92 VN.n64 0.189894
R143 VN.n92 VN.n91 0.189894
R144 VN.n91 VN.n90 0.189894
R145 VN.n90 VN.n66 0.189894
R146 VN.n85 VN.n66 0.189894
R147 VN.n85 VN.n84 0.189894
R148 VN.n84 VN.n83 0.189894
R149 VN.n83 VN.n68 0.189894
R150 VN.n79 VN.n68 0.189894
R151 VN.n79 VN.n78 0.189894
R152 VN.n78 VN.n77 0.189894
R153 VN.n77 VN.n70 0.189894
R154 VN.n73 VN.n70 0.189894
R155 VN.n15 VN.n12 0.189894
R156 VN.n19 VN.n12 0.189894
R157 VN.n20 VN.n19 0.189894
R158 VN.n21 VN.n20 0.189894
R159 VN.n21 VN.n10 0.189894
R160 VN.n25 VN.n10 0.189894
R161 VN.n26 VN.n25 0.189894
R162 VN.n27 VN.n26 0.189894
R163 VN.n27 VN.n8 0.189894
R164 VN.n32 VN.n8 0.189894
R165 VN.n33 VN.n32 0.189894
R166 VN.n34 VN.n33 0.189894
R167 VN.n34 VN.n6 0.189894
R168 VN.n38 VN.n6 0.189894
R169 VN.n39 VN.n38 0.189894
R170 VN.n40 VN.n39 0.189894
R171 VN.n40 VN.n4 0.189894
R172 VN.n45 VN.n4 0.189894
R173 VN.n46 VN.n45 0.189894
R174 VN.n47 VN.n46 0.189894
R175 VN.n47 VN.n2 0.189894
R176 VN.n51 VN.n2 0.189894
R177 VN.n52 VN.n51 0.189894
R178 VN.n53 VN.n52 0.189894
R179 VN.n53 VN.n0 0.189894
R180 VTAIL.n11 VTAIL.t11 56.8323
R181 VTAIL.n17 VTAIL.t17 56.8322
R182 VTAIL.n2 VTAIL.t9 56.8322
R183 VTAIL.n16 VTAIL.t3 56.8322
R184 VTAIL.n15 VTAIL.n14 54.5577
R185 VTAIL.n13 VTAIL.n12 54.5577
R186 VTAIL.n10 VTAIL.n9 54.5577
R187 VTAIL.n8 VTAIL.n7 54.5577
R188 VTAIL.n19 VTAIL.n18 54.5575
R189 VTAIL.n1 VTAIL.n0 54.5575
R190 VTAIL.n4 VTAIL.n3 54.5575
R191 VTAIL.n6 VTAIL.n5 54.5575
R192 VTAIL.n8 VTAIL.n6 32.1514
R193 VTAIL.n17 VTAIL.n16 28.4186
R194 VTAIL.n10 VTAIL.n8 3.73326
R195 VTAIL.n11 VTAIL.n10 3.73326
R196 VTAIL.n15 VTAIL.n13 3.73326
R197 VTAIL.n16 VTAIL.n15 3.73326
R198 VTAIL.n6 VTAIL.n4 3.73326
R199 VTAIL.n4 VTAIL.n2 3.73326
R200 VTAIL.n19 VTAIL.n17 3.73326
R201 VTAIL VTAIL.n1 2.85826
R202 VTAIL.n13 VTAIL.n11 2.33671
R203 VTAIL.n2 VTAIL.n1 2.33671
R204 VTAIL.n18 VTAIL.t12 2.27517
R205 VTAIL.n18 VTAIL.t14 2.27517
R206 VTAIL.n0 VTAIL.t16 2.27517
R207 VTAIL.n0 VTAIL.t15 2.27517
R208 VTAIL.n3 VTAIL.t7 2.27517
R209 VTAIL.n3 VTAIL.t0 2.27517
R210 VTAIL.n5 VTAIL.t6 2.27517
R211 VTAIL.n5 VTAIL.t5 2.27517
R212 VTAIL.n14 VTAIL.t1 2.27517
R213 VTAIL.n14 VTAIL.t2 2.27517
R214 VTAIL.n12 VTAIL.t8 2.27517
R215 VTAIL.n12 VTAIL.t4 2.27517
R216 VTAIL.n9 VTAIL.t18 2.27517
R217 VTAIL.n9 VTAIL.t10 2.27517
R218 VTAIL.n7 VTAIL.t19 2.27517
R219 VTAIL.n7 VTAIL.t13 2.27517
R220 VTAIL VTAIL.n19 0.8755
R221 VDD2.n1 VDD2.t5 77.2438
R222 VDD2.n3 VDD2.n2 73.9805
R223 VDD2 VDD2.n7 73.9777
R224 VDD2.n4 VDD2.t6 73.5111
R225 VDD2.n6 VDD2.n5 71.2365
R226 VDD2.n1 VDD2.n0 71.2363
R227 VDD2.n4 VDD2.n3 53.7649
R228 VDD2.n6 VDD2.n4 3.73326
R229 VDD2.n7 VDD2.t0 2.27517
R230 VDD2.n7 VDD2.t4 2.27517
R231 VDD2.n5 VDD2.t8 2.27517
R232 VDD2.n5 VDD2.t9 2.27517
R233 VDD2.n2 VDD2.t2 2.27517
R234 VDD2.n2 VDD2.t3 2.27517
R235 VDD2.n0 VDD2.t1 2.27517
R236 VDD2.n0 VDD2.t7 2.27517
R237 VDD2 VDD2.n6 0.991879
R238 VDD2.n3 VDD2.n1 0.878344
R239 VP.n34 VP.n33 161.3
R240 VP.n35 VP.n30 161.3
R241 VP.n37 VP.n36 161.3
R242 VP.n38 VP.n29 161.3
R243 VP.n40 VP.n39 161.3
R244 VP.n41 VP.n28 161.3
R245 VP.n43 VP.n42 161.3
R246 VP.n44 VP.n27 161.3
R247 VP.n46 VP.n45 161.3
R248 VP.n48 VP.n26 161.3
R249 VP.n50 VP.n49 161.3
R250 VP.n51 VP.n25 161.3
R251 VP.n53 VP.n52 161.3
R252 VP.n54 VP.n24 161.3
R253 VP.n56 VP.n55 161.3
R254 VP.n57 VP.n23 161.3
R255 VP.n59 VP.n58 161.3
R256 VP.n60 VP.n22 161.3
R257 VP.n63 VP.n62 161.3
R258 VP.n64 VP.n21 161.3
R259 VP.n66 VP.n65 161.3
R260 VP.n67 VP.n20 161.3
R261 VP.n69 VP.n68 161.3
R262 VP.n70 VP.n19 161.3
R263 VP.n72 VP.n71 161.3
R264 VP.n73 VP.n18 161.3
R265 VP.n130 VP.n0 161.3
R266 VP.n129 VP.n128 161.3
R267 VP.n127 VP.n1 161.3
R268 VP.n126 VP.n125 161.3
R269 VP.n124 VP.n2 161.3
R270 VP.n123 VP.n122 161.3
R271 VP.n121 VP.n3 161.3
R272 VP.n120 VP.n119 161.3
R273 VP.n117 VP.n4 161.3
R274 VP.n116 VP.n115 161.3
R275 VP.n114 VP.n5 161.3
R276 VP.n113 VP.n112 161.3
R277 VP.n111 VP.n6 161.3
R278 VP.n110 VP.n109 161.3
R279 VP.n108 VP.n7 161.3
R280 VP.n107 VP.n106 161.3
R281 VP.n105 VP.n8 161.3
R282 VP.n103 VP.n102 161.3
R283 VP.n101 VP.n9 161.3
R284 VP.n100 VP.n99 161.3
R285 VP.n98 VP.n10 161.3
R286 VP.n97 VP.n96 161.3
R287 VP.n95 VP.n11 161.3
R288 VP.n94 VP.n93 161.3
R289 VP.n92 VP.n12 161.3
R290 VP.n91 VP.n90 161.3
R291 VP.n89 VP.n88 161.3
R292 VP.n87 VP.n14 161.3
R293 VP.n86 VP.n85 161.3
R294 VP.n84 VP.n15 161.3
R295 VP.n83 VP.n82 161.3
R296 VP.n81 VP.n16 161.3
R297 VP.n80 VP.n79 161.3
R298 VP.n78 VP.n17 161.3
R299 VP.n32 VP.t9 118.367
R300 VP.n76 VP.t8 86.0978
R301 VP.n13 VP.t5 86.0978
R302 VP.n104 VP.t4 86.0978
R303 VP.n118 VP.t7 86.0978
R304 VP.n131 VP.t6 86.0978
R305 VP.n74 VP.t3 86.0978
R306 VP.n61 VP.t1 86.0978
R307 VP.n47 VP.t0 86.0978
R308 VP.n31 VP.t2 86.0978
R309 VP.n32 VP.n31 71.1463
R310 VP.n77 VP.n75 62.7048
R311 VP.n77 VP.n76 62.1188
R312 VP.n132 VP.n131 62.1188
R313 VP.n75 VP.n74 62.1188
R314 VP.n82 VP.n15 56.5193
R315 VP.n125 VP.n124 56.5193
R316 VP.n68 VP.n67 56.5193
R317 VP.n98 VP.n97 48.7492
R318 VP.n111 VP.n110 48.7492
R319 VP.n54 VP.n53 48.7492
R320 VP.n41 VP.n40 48.7492
R321 VP.n97 VP.n11 32.2376
R322 VP.n112 VP.n111 32.2376
R323 VP.n55 VP.n54 32.2376
R324 VP.n40 VP.n29 32.2376
R325 VP.n80 VP.n17 24.4675
R326 VP.n81 VP.n80 24.4675
R327 VP.n82 VP.n81 24.4675
R328 VP.n86 VP.n15 24.4675
R329 VP.n87 VP.n86 24.4675
R330 VP.n88 VP.n87 24.4675
R331 VP.n92 VP.n91 24.4675
R332 VP.n93 VP.n92 24.4675
R333 VP.n93 VP.n11 24.4675
R334 VP.n99 VP.n98 24.4675
R335 VP.n99 VP.n9 24.4675
R336 VP.n103 VP.n9 24.4675
R337 VP.n106 VP.n105 24.4675
R338 VP.n106 VP.n7 24.4675
R339 VP.n110 VP.n7 24.4675
R340 VP.n112 VP.n5 24.4675
R341 VP.n116 VP.n5 24.4675
R342 VP.n117 VP.n116 24.4675
R343 VP.n119 VP.n3 24.4675
R344 VP.n123 VP.n3 24.4675
R345 VP.n124 VP.n123 24.4675
R346 VP.n125 VP.n1 24.4675
R347 VP.n129 VP.n1 24.4675
R348 VP.n130 VP.n129 24.4675
R349 VP.n68 VP.n19 24.4675
R350 VP.n72 VP.n19 24.4675
R351 VP.n73 VP.n72 24.4675
R352 VP.n55 VP.n23 24.4675
R353 VP.n59 VP.n23 24.4675
R354 VP.n60 VP.n59 24.4675
R355 VP.n62 VP.n21 24.4675
R356 VP.n66 VP.n21 24.4675
R357 VP.n67 VP.n66 24.4675
R358 VP.n42 VP.n41 24.4675
R359 VP.n42 VP.n27 24.4675
R360 VP.n46 VP.n27 24.4675
R361 VP.n49 VP.n48 24.4675
R362 VP.n49 VP.n25 24.4675
R363 VP.n53 VP.n25 24.4675
R364 VP.n35 VP.n34 24.4675
R365 VP.n36 VP.n35 24.4675
R366 VP.n36 VP.n29 24.4675
R367 VP.n88 VP.n13 20.5528
R368 VP.n119 VP.n118 20.5528
R369 VP.n62 VP.n61 20.5528
R370 VP.n76 VP.n17 20.0634
R371 VP.n131 VP.n130 20.0634
R372 VP.n74 VP.n73 20.0634
R373 VP.n104 VP.n103 12.234
R374 VP.n105 VP.n104 12.234
R375 VP.n47 VP.n46 12.234
R376 VP.n48 VP.n47 12.234
R377 VP.n91 VP.n13 3.91522
R378 VP.n118 VP.n117 3.91522
R379 VP.n61 VP.n60 3.91522
R380 VP.n34 VP.n31 3.91522
R381 VP.n33 VP.n32 2.69182
R382 VP.n75 VP.n18 0.417535
R383 VP.n78 VP.n77 0.417535
R384 VP.n132 VP.n0 0.417535
R385 VP VP.n132 0.394291
R386 VP.n33 VP.n30 0.189894
R387 VP.n37 VP.n30 0.189894
R388 VP.n38 VP.n37 0.189894
R389 VP.n39 VP.n38 0.189894
R390 VP.n39 VP.n28 0.189894
R391 VP.n43 VP.n28 0.189894
R392 VP.n44 VP.n43 0.189894
R393 VP.n45 VP.n44 0.189894
R394 VP.n45 VP.n26 0.189894
R395 VP.n50 VP.n26 0.189894
R396 VP.n51 VP.n50 0.189894
R397 VP.n52 VP.n51 0.189894
R398 VP.n52 VP.n24 0.189894
R399 VP.n56 VP.n24 0.189894
R400 VP.n57 VP.n56 0.189894
R401 VP.n58 VP.n57 0.189894
R402 VP.n58 VP.n22 0.189894
R403 VP.n63 VP.n22 0.189894
R404 VP.n64 VP.n63 0.189894
R405 VP.n65 VP.n64 0.189894
R406 VP.n65 VP.n20 0.189894
R407 VP.n69 VP.n20 0.189894
R408 VP.n70 VP.n69 0.189894
R409 VP.n71 VP.n70 0.189894
R410 VP.n71 VP.n18 0.189894
R411 VP.n79 VP.n78 0.189894
R412 VP.n79 VP.n16 0.189894
R413 VP.n83 VP.n16 0.189894
R414 VP.n84 VP.n83 0.189894
R415 VP.n85 VP.n84 0.189894
R416 VP.n85 VP.n14 0.189894
R417 VP.n89 VP.n14 0.189894
R418 VP.n90 VP.n89 0.189894
R419 VP.n90 VP.n12 0.189894
R420 VP.n94 VP.n12 0.189894
R421 VP.n95 VP.n94 0.189894
R422 VP.n96 VP.n95 0.189894
R423 VP.n96 VP.n10 0.189894
R424 VP.n100 VP.n10 0.189894
R425 VP.n101 VP.n100 0.189894
R426 VP.n102 VP.n101 0.189894
R427 VP.n102 VP.n8 0.189894
R428 VP.n107 VP.n8 0.189894
R429 VP.n108 VP.n107 0.189894
R430 VP.n109 VP.n108 0.189894
R431 VP.n109 VP.n6 0.189894
R432 VP.n113 VP.n6 0.189894
R433 VP.n114 VP.n113 0.189894
R434 VP.n115 VP.n114 0.189894
R435 VP.n115 VP.n4 0.189894
R436 VP.n120 VP.n4 0.189894
R437 VP.n121 VP.n120 0.189894
R438 VP.n122 VP.n121 0.189894
R439 VP.n122 VP.n2 0.189894
R440 VP.n126 VP.n2 0.189894
R441 VP.n127 VP.n126 0.189894
R442 VP.n128 VP.n127 0.189894
R443 VP.n128 VP.n0 0.189894
R444 VDD1.n1 VDD1.t0 77.2439
R445 VDD1.n3 VDD1.t1 77.2438
R446 VDD1.n5 VDD1.n4 73.9805
R447 VDD1.n1 VDD1.n0 71.2365
R448 VDD1.n7 VDD1.n6 71.2363
R449 VDD1.n3 VDD1.n2 71.2363
R450 VDD1.n7 VDD1.n5 56.2143
R451 VDD1 VDD1.n7 2.74188
R452 VDD1.n6 VDD1.t8 2.27517
R453 VDD1.n6 VDD1.t6 2.27517
R454 VDD1.n0 VDD1.t7 2.27517
R455 VDD1.n0 VDD1.t9 2.27517
R456 VDD1.n4 VDD1.t2 2.27517
R457 VDD1.n4 VDD1.t3 2.27517
R458 VDD1.n2 VDD1.t4 2.27517
R459 VDD1.n2 VDD1.t5 2.27517
R460 VDD1 VDD1.n1 0.991879
R461 VDD1.n5 VDD1.n3 0.878344
R462 B.n570 B.n569 585
R463 B.n568 B.n187 585
R464 B.n567 B.n566 585
R465 B.n565 B.n188 585
R466 B.n564 B.n563 585
R467 B.n562 B.n189 585
R468 B.n561 B.n560 585
R469 B.n559 B.n190 585
R470 B.n558 B.n557 585
R471 B.n556 B.n191 585
R472 B.n555 B.n554 585
R473 B.n553 B.n192 585
R474 B.n552 B.n551 585
R475 B.n550 B.n193 585
R476 B.n549 B.n548 585
R477 B.n547 B.n194 585
R478 B.n546 B.n545 585
R479 B.n544 B.n195 585
R480 B.n543 B.n542 585
R481 B.n541 B.n196 585
R482 B.n540 B.n539 585
R483 B.n538 B.n197 585
R484 B.n537 B.n536 585
R485 B.n535 B.n198 585
R486 B.n534 B.n533 585
R487 B.n532 B.n199 585
R488 B.n531 B.n530 585
R489 B.n529 B.n200 585
R490 B.n528 B.n527 585
R491 B.n526 B.n201 585
R492 B.n525 B.n524 585
R493 B.n523 B.n202 585
R494 B.n522 B.n521 585
R495 B.n520 B.n203 585
R496 B.n519 B.n518 585
R497 B.n517 B.n204 585
R498 B.n516 B.n515 585
R499 B.n514 B.n205 585
R500 B.n513 B.n512 585
R501 B.n511 B.n206 585
R502 B.n510 B.n509 585
R503 B.n508 B.n207 585
R504 B.n507 B.n506 585
R505 B.n505 B.n208 585
R506 B.n504 B.n503 585
R507 B.n502 B.n209 585
R508 B.n501 B.n500 585
R509 B.n499 B.n210 585
R510 B.n498 B.n497 585
R511 B.n493 B.n211 585
R512 B.n492 B.n491 585
R513 B.n490 B.n212 585
R514 B.n489 B.n488 585
R515 B.n487 B.n213 585
R516 B.n486 B.n485 585
R517 B.n484 B.n214 585
R518 B.n483 B.n482 585
R519 B.n481 B.n215 585
R520 B.n479 B.n478 585
R521 B.n477 B.n218 585
R522 B.n476 B.n475 585
R523 B.n474 B.n219 585
R524 B.n473 B.n472 585
R525 B.n471 B.n220 585
R526 B.n470 B.n469 585
R527 B.n468 B.n221 585
R528 B.n467 B.n466 585
R529 B.n465 B.n222 585
R530 B.n464 B.n463 585
R531 B.n462 B.n223 585
R532 B.n461 B.n460 585
R533 B.n459 B.n224 585
R534 B.n458 B.n457 585
R535 B.n456 B.n225 585
R536 B.n455 B.n454 585
R537 B.n453 B.n226 585
R538 B.n452 B.n451 585
R539 B.n450 B.n227 585
R540 B.n449 B.n448 585
R541 B.n447 B.n228 585
R542 B.n446 B.n445 585
R543 B.n444 B.n229 585
R544 B.n443 B.n442 585
R545 B.n441 B.n230 585
R546 B.n440 B.n439 585
R547 B.n438 B.n231 585
R548 B.n437 B.n436 585
R549 B.n435 B.n232 585
R550 B.n434 B.n433 585
R551 B.n432 B.n233 585
R552 B.n431 B.n430 585
R553 B.n429 B.n234 585
R554 B.n428 B.n427 585
R555 B.n426 B.n235 585
R556 B.n425 B.n424 585
R557 B.n423 B.n236 585
R558 B.n422 B.n421 585
R559 B.n420 B.n237 585
R560 B.n419 B.n418 585
R561 B.n417 B.n238 585
R562 B.n416 B.n415 585
R563 B.n414 B.n239 585
R564 B.n413 B.n412 585
R565 B.n411 B.n240 585
R566 B.n410 B.n409 585
R567 B.n408 B.n241 585
R568 B.n571 B.n186 585
R569 B.n573 B.n572 585
R570 B.n574 B.n185 585
R571 B.n576 B.n575 585
R572 B.n577 B.n184 585
R573 B.n579 B.n578 585
R574 B.n580 B.n183 585
R575 B.n582 B.n581 585
R576 B.n583 B.n182 585
R577 B.n585 B.n584 585
R578 B.n586 B.n181 585
R579 B.n588 B.n587 585
R580 B.n589 B.n180 585
R581 B.n591 B.n590 585
R582 B.n592 B.n179 585
R583 B.n594 B.n593 585
R584 B.n595 B.n178 585
R585 B.n597 B.n596 585
R586 B.n598 B.n177 585
R587 B.n600 B.n599 585
R588 B.n601 B.n176 585
R589 B.n603 B.n602 585
R590 B.n604 B.n175 585
R591 B.n606 B.n605 585
R592 B.n607 B.n174 585
R593 B.n609 B.n608 585
R594 B.n610 B.n173 585
R595 B.n612 B.n611 585
R596 B.n613 B.n172 585
R597 B.n615 B.n614 585
R598 B.n616 B.n171 585
R599 B.n618 B.n617 585
R600 B.n619 B.n170 585
R601 B.n621 B.n620 585
R602 B.n622 B.n169 585
R603 B.n624 B.n623 585
R604 B.n625 B.n168 585
R605 B.n627 B.n626 585
R606 B.n628 B.n167 585
R607 B.n630 B.n629 585
R608 B.n631 B.n166 585
R609 B.n633 B.n632 585
R610 B.n634 B.n165 585
R611 B.n636 B.n635 585
R612 B.n637 B.n164 585
R613 B.n639 B.n638 585
R614 B.n640 B.n163 585
R615 B.n642 B.n641 585
R616 B.n643 B.n162 585
R617 B.n645 B.n644 585
R618 B.n646 B.n161 585
R619 B.n648 B.n647 585
R620 B.n649 B.n160 585
R621 B.n651 B.n650 585
R622 B.n652 B.n159 585
R623 B.n654 B.n653 585
R624 B.n655 B.n158 585
R625 B.n657 B.n656 585
R626 B.n658 B.n157 585
R627 B.n660 B.n659 585
R628 B.n661 B.n156 585
R629 B.n663 B.n662 585
R630 B.n664 B.n155 585
R631 B.n666 B.n665 585
R632 B.n667 B.n154 585
R633 B.n669 B.n668 585
R634 B.n670 B.n153 585
R635 B.n672 B.n671 585
R636 B.n673 B.n152 585
R637 B.n675 B.n674 585
R638 B.n676 B.n151 585
R639 B.n678 B.n677 585
R640 B.n679 B.n150 585
R641 B.n681 B.n680 585
R642 B.n682 B.n149 585
R643 B.n684 B.n683 585
R644 B.n685 B.n148 585
R645 B.n687 B.n686 585
R646 B.n688 B.n147 585
R647 B.n690 B.n689 585
R648 B.n691 B.n146 585
R649 B.n693 B.n692 585
R650 B.n694 B.n145 585
R651 B.n696 B.n695 585
R652 B.n697 B.n144 585
R653 B.n699 B.n698 585
R654 B.n700 B.n143 585
R655 B.n702 B.n701 585
R656 B.n703 B.n142 585
R657 B.n705 B.n704 585
R658 B.n706 B.n141 585
R659 B.n708 B.n707 585
R660 B.n709 B.n140 585
R661 B.n711 B.n710 585
R662 B.n712 B.n139 585
R663 B.n714 B.n713 585
R664 B.n715 B.n138 585
R665 B.n717 B.n716 585
R666 B.n718 B.n137 585
R667 B.n720 B.n719 585
R668 B.n721 B.n136 585
R669 B.n723 B.n722 585
R670 B.n724 B.n135 585
R671 B.n726 B.n725 585
R672 B.n727 B.n134 585
R673 B.n729 B.n728 585
R674 B.n730 B.n133 585
R675 B.n732 B.n731 585
R676 B.n733 B.n132 585
R677 B.n735 B.n734 585
R678 B.n736 B.n131 585
R679 B.n738 B.n737 585
R680 B.n739 B.n130 585
R681 B.n741 B.n740 585
R682 B.n742 B.n129 585
R683 B.n744 B.n743 585
R684 B.n745 B.n128 585
R685 B.n747 B.n746 585
R686 B.n748 B.n127 585
R687 B.n750 B.n749 585
R688 B.n751 B.n126 585
R689 B.n753 B.n752 585
R690 B.n754 B.n125 585
R691 B.n756 B.n755 585
R692 B.n757 B.n124 585
R693 B.n759 B.n758 585
R694 B.n760 B.n123 585
R695 B.n762 B.n761 585
R696 B.n763 B.n122 585
R697 B.n765 B.n764 585
R698 B.n766 B.n121 585
R699 B.n768 B.n767 585
R700 B.n769 B.n120 585
R701 B.n771 B.n770 585
R702 B.n772 B.n119 585
R703 B.n774 B.n773 585
R704 B.n775 B.n118 585
R705 B.n777 B.n776 585
R706 B.n778 B.n117 585
R707 B.n780 B.n779 585
R708 B.n781 B.n116 585
R709 B.n783 B.n782 585
R710 B.n784 B.n115 585
R711 B.n786 B.n785 585
R712 B.n787 B.n114 585
R713 B.n789 B.n788 585
R714 B.n790 B.n113 585
R715 B.n792 B.n791 585
R716 B.n793 B.n112 585
R717 B.n795 B.n794 585
R718 B.n796 B.n111 585
R719 B.n798 B.n797 585
R720 B.n799 B.n110 585
R721 B.n801 B.n800 585
R722 B.n802 B.n109 585
R723 B.n804 B.n803 585
R724 B.n805 B.n108 585
R725 B.n807 B.n806 585
R726 B.n808 B.n107 585
R727 B.n810 B.n809 585
R728 B.n811 B.n106 585
R729 B.n813 B.n812 585
R730 B.n814 B.n105 585
R731 B.n816 B.n815 585
R732 B.n817 B.n104 585
R733 B.n819 B.n818 585
R734 B.n820 B.n103 585
R735 B.n822 B.n821 585
R736 B.n823 B.n102 585
R737 B.n825 B.n824 585
R738 B.n985 B.n44 585
R739 B.n984 B.n983 585
R740 B.n982 B.n45 585
R741 B.n981 B.n980 585
R742 B.n979 B.n46 585
R743 B.n978 B.n977 585
R744 B.n976 B.n47 585
R745 B.n975 B.n974 585
R746 B.n973 B.n48 585
R747 B.n972 B.n971 585
R748 B.n970 B.n49 585
R749 B.n969 B.n968 585
R750 B.n967 B.n50 585
R751 B.n966 B.n965 585
R752 B.n964 B.n51 585
R753 B.n963 B.n962 585
R754 B.n961 B.n52 585
R755 B.n960 B.n959 585
R756 B.n958 B.n53 585
R757 B.n957 B.n956 585
R758 B.n955 B.n54 585
R759 B.n954 B.n953 585
R760 B.n952 B.n55 585
R761 B.n951 B.n950 585
R762 B.n949 B.n56 585
R763 B.n948 B.n947 585
R764 B.n946 B.n57 585
R765 B.n945 B.n944 585
R766 B.n943 B.n58 585
R767 B.n942 B.n941 585
R768 B.n940 B.n59 585
R769 B.n939 B.n938 585
R770 B.n937 B.n60 585
R771 B.n936 B.n935 585
R772 B.n934 B.n61 585
R773 B.n933 B.n932 585
R774 B.n931 B.n62 585
R775 B.n930 B.n929 585
R776 B.n928 B.n63 585
R777 B.n927 B.n926 585
R778 B.n925 B.n64 585
R779 B.n924 B.n923 585
R780 B.n922 B.n65 585
R781 B.n921 B.n920 585
R782 B.n919 B.n66 585
R783 B.n918 B.n917 585
R784 B.n916 B.n67 585
R785 B.n915 B.n914 585
R786 B.n913 B.n912 585
R787 B.n911 B.n71 585
R788 B.n910 B.n909 585
R789 B.n908 B.n72 585
R790 B.n907 B.n906 585
R791 B.n905 B.n73 585
R792 B.n904 B.n903 585
R793 B.n902 B.n74 585
R794 B.n901 B.n900 585
R795 B.n899 B.n75 585
R796 B.n897 B.n896 585
R797 B.n895 B.n78 585
R798 B.n894 B.n893 585
R799 B.n892 B.n79 585
R800 B.n891 B.n890 585
R801 B.n889 B.n80 585
R802 B.n888 B.n887 585
R803 B.n886 B.n81 585
R804 B.n885 B.n884 585
R805 B.n883 B.n82 585
R806 B.n882 B.n881 585
R807 B.n880 B.n83 585
R808 B.n879 B.n878 585
R809 B.n877 B.n84 585
R810 B.n876 B.n875 585
R811 B.n874 B.n85 585
R812 B.n873 B.n872 585
R813 B.n871 B.n86 585
R814 B.n870 B.n869 585
R815 B.n868 B.n87 585
R816 B.n867 B.n866 585
R817 B.n865 B.n88 585
R818 B.n864 B.n863 585
R819 B.n862 B.n89 585
R820 B.n861 B.n860 585
R821 B.n859 B.n90 585
R822 B.n858 B.n857 585
R823 B.n856 B.n91 585
R824 B.n855 B.n854 585
R825 B.n853 B.n92 585
R826 B.n852 B.n851 585
R827 B.n850 B.n93 585
R828 B.n849 B.n848 585
R829 B.n847 B.n94 585
R830 B.n846 B.n845 585
R831 B.n844 B.n95 585
R832 B.n843 B.n842 585
R833 B.n841 B.n96 585
R834 B.n840 B.n839 585
R835 B.n838 B.n97 585
R836 B.n837 B.n836 585
R837 B.n835 B.n98 585
R838 B.n834 B.n833 585
R839 B.n832 B.n99 585
R840 B.n831 B.n830 585
R841 B.n829 B.n100 585
R842 B.n828 B.n827 585
R843 B.n826 B.n101 585
R844 B.n987 B.n986 585
R845 B.n988 B.n43 585
R846 B.n990 B.n989 585
R847 B.n991 B.n42 585
R848 B.n993 B.n992 585
R849 B.n994 B.n41 585
R850 B.n996 B.n995 585
R851 B.n997 B.n40 585
R852 B.n999 B.n998 585
R853 B.n1000 B.n39 585
R854 B.n1002 B.n1001 585
R855 B.n1003 B.n38 585
R856 B.n1005 B.n1004 585
R857 B.n1006 B.n37 585
R858 B.n1008 B.n1007 585
R859 B.n1009 B.n36 585
R860 B.n1011 B.n1010 585
R861 B.n1012 B.n35 585
R862 B.n1014 B.n1013 585
R863 B.n1015 B.n34 585
R864 B.n1017 B.n1016 585
R865 B.n1018 B.n33 585
R866 B.n1020 B.n1019 585
R867 B.n1021 B.n32 585
R868 B.n1023 B.n1022 585
R869 B.n1024 B.n31 585
R870 B.n1026 B.n1025 585
R871 B.n1027 B.n30 585
R872 B.n1029 B.n1028 585
R873 B.n1030 B.n29 585
R874 B.n1032 B.n1031 585
R875 B.n1033 B.n28 585
R876 B.n1035 B.n1034 585
R877 B.n1036 B.n27 585
R878 B.n1038 B.n1037 585
R879 B.n1039 B.n26 585
R880 B.n1041 B.n1040 585
R881 B.n1042 B.n25 585
R882 B.n1044 B.n1043 585
R883 B.n1045 B.n24 585
R884 B.n1047 B.n1046 585
R885 B.n1048 B.n23 585
R886 B.n1050 B.n1049 585
R887 B.n1051 B.n22 585
R888 B.n1053 B.n1052 585
R889 B.n1054 B.n21 585
R890 B.n1056 B.n1055 585
R891 B.n1057 B.n20 585
R892 B.n1059 B.n1058 585
R893 B.n1060 B.n19 585
R894 B.n1062 B.n1061 585
R895 B.n1063 B.n18 585
R896 B.n1065 B.n1064 585
R897 B.n1066 B.n17 585
R898 B.n1068 B.n1067 585
R899 B.n1069 B.n16 585
R900 B.n1071 B.n1070 585
R901 B.n1072 B.n15 585
R902 B.n1074 B.n1073 585
R903 B.n1075 B.n14 585
R904 B.n1077 B.n1076 585
R905 B.n1078 B.n13 585
R906 B.n1080 B.n1079 585
R907 B.n1081 B.n12 585
R908 B.n1083 B.n1082 585
R909 B.n1084 B.n11 585
R910 B.n1086 B.n1085 585
R911 B.n1087 B.n10 585
R912 B.n1089 B.n1088 585
R913 B.n1090 B.n9 585
R914 B.n1092 B.n1091 585
R915 B.n1093 B.n8 585
R916 B.n1095 B.n1094 585
R917 B.n1096 B.n7 585
R918 B.n1098 B.n1097 585
R919 B.n1099 B.n6 585
R920 B.n1101 B.n1100 585
R921 B.n1102 B.n5 585
R922 B.n1104 B.n1103 585
R923 B.n1105 B.n4 585
R924 B.n1107 B.n1106 585
R925 B.n1108 B.n3 585
R926 B.n1110 B.n1109 585
R927 B.n1111 B.n0 585
R928 B.n2 B.n1 585
R929 B.n284 B.n283 585
R930 B.n285 B.n282 585
R931 B.n287 B.n286 585
R932 B.n288 B.n281 585
R933 B.n290 B.n289 585
R934 B.n291 B.n280 585
R935 B.n293 B.n292 585
R936 B.n294 B.n279 585
R937 B.n296 B.n295 585
R938 B.n297 B.n278 585
R939 B.n299 B.n298 585
R940 B.n300 B.n277 585
R941 B.n302 B.n301 585
R942 B.n303 B.n276 585
R943 B.n305 B.n304 585
R944 B.n306 B.n275 585
R945 B.n308 B.n307 585
R946 B.n309 B.n274 585
R947 B.n311 B.n310 585
R948 B.n312 B.n273 585
R949 B.n314 B.n313 585
R950 B.n315 B.n272 585
R951 B.n317 B.n316 585
R952 B.n318 B.n271 585
R953 B.n320 B.n319 585
R954 B.n321 B.n270 585
R955 B.n323 B.n322 585
R956 B.n324 B.n269 585
R957 B.n326 B.n325 585
R958 B.n327 B.n268 585
R959 B.n329 B.n328 585
R960 B.n330 B.n267 585
R961 B.n332 B.n331 585
R962 B.n333 B.n266 585
R963 B.n335 B.n334 585
R964 B.n336 B.n265 585
R965 B.n338 B.n337 585
R966 B.n339 B.n264 585
R967 B.n341 B.n340 585
R968 B.n342 B.n263 585
R969 B.n344 B.n343 585
R970 B.n345 B.n262 585
R971 B.n347 B.n346 585
R972 B.n348 B.n261 585
R973 B.n350 B.n349 585
R974 B.n351 B.n260 585
R975 B.n353 B.n352 585
R976 B.n354 B.n259 585
R977 B.n356 B.n355 585
R978 B.n357 B.n258 585
R979 B.n359 B.n358 585
R980 B.n360 B.n257 585
R981 B.n362 B.n361 585
R982 B.n363 B.n256 585
R983 B.n365 B.n364 585
R984 B.n366 B.n255 585
R985 B.n368 B.n367 585
R986 B.n369 B.n254 585
R987 B.n371 B.n370 585
R988 B.n372 B.n253 585
R989 B.n374 B.n373 585
R990 B.n375 B.n252 585
R991 B.n377 B.n376 585
R992 B.n378 B.n251 585
R993 B.n380 B.n379 585
R994 B.n381 B.n250 585
R995 B.n383 B.n382 585
R996 B.n384 B.n249 585
R997 B.n386 B.n385 585
R998 B.n387 B.n248 585
R999 B.n389 B.n388 585
R1000 B.n390 B.n247 585
R1001 B.n392 B.n391 585
R1002 B.n393 B.n246 585
R1003 B.n395 B.n394 585
R1004 B.n396 B.n245 585
R1005 B.n398 B.n397 585
R1006 B.n399 B.n244 585
R1007 B.n401 B.n400 585
R1008 B.n402 B.n243 585
R1009 B.n404 B.n403 585
R1010 B.n405 B.n242 585
R1011 B.n407 B.n406 585
R1012 B.n406 B.n241 526.135
R1013 B.n571 B.n570 526.135
R1014 B.n824 B.n101 526.135
R1015 B.n986 B.n985 526.135
R1016 B.n216 B.t0 295.589
R1017 B.n494 B.t9 295.589
R1018 B.n76 B.t6 295.589
R1019 B.n68 B.t3 295.589
R1020 B.n1113 B.n1112 256.663
R1021 B.n1112 B.n1111 235.042
R1022 B.n1112 B.n2 235.042
R1023 B.n494 B.t10 190.839
R1024 B.n76 B.t8 190.839
R1025 B.n216 B.t1 190.821
R1026 B.n68 B.t5 190.821
R1027 B.n410 B.n241 163.367
R1028 B.n411 B.n410 163.367
R1029 B.n412 B.n411 163.367
R1030 B.n412 B.n239 163.367
R1031 B.n416 B.n239 163.367
R1032 B.n417 B.n416 163.367
R1033 B.n418 B.n417 163.367
R1034 B.n418 B.n237 163.367
R1035 B.n422 B.n237 163.367
R1036 B.n423 B.n422 163.367
R1037 B.n424 B.n423 163.367
R1038 B.n424 B.n235 163.367
R1039 B.n428 B.n235 163.367
R1040 B.n429 B.n428 163.367
R1041 B.n430 B.n429 163.367
R1042 B.n430 B.n233 163.367
R1043 B.n434 B.n233 163.367
R1044 B.n435 B.n434 163.367
R1045 B.n436 B.n435 163.367
R1046 B.n436 B.n231 163.367
R1047 B.n440 B.n231 163.367
R1048 B.n441 B.n440 163.367
R1049 B.n442 B.n441 163.367
R1050 B.n442 B.n229 163.367
R1051 B.n446 B.n229 163.367
R1052 B.n447 B.n446 163.367
R1053 B.n448 B.n447 163.367
R1054 B.n448 B.n227 163.367
R1055 B.n452 B.n227 163.367
R1056 B.n453 B.n452 163.367
R1057 B.n454 B.n453 163.367
R1058 B.n454 B.n225 163.367
R1059 B.n458 B.n225 163.367
R1060 B.n459 B.n458 163.367
R1061 B.n460 B.n459 163.367
R1062 B.n460 B.n223 163.367
R1063 B.n464 B.n223 163.367
R1064 B.n465 B.n464 163.367
R1065 B.n466 B.n465 163.367
R1066 B.n466 B.n221 163.367
R1067 B.n470 B.n221 163.367
R1068 B.n471 B.n470 163.367
R1069 B.n472 B.n471 163.367
R1070 B.n472 B.n219 163.367
R1071 B.n476 B.n219 163.367
R1072 B.n477 B.n476 163.367
R1073 B.n478 B.n477 163.367
R1074 B.n478 B.n215 163.367
R1075 B.n483 B.n215 163.367
R1076 B.n484 B.n483 163.367
R1077 B.n485 B.n484 163.367
R1078 B.n485 B.n213 163.367
R1079 B.n489 B.n213 163.367
R1080 B.n490 B.n489 163.367
R1081 B.n491 B.n490 163.367
R1082 B.n491 B.n211 163.367
R1083 B.n498 B.n211 163.367
R1084 B.n499 B.n498 163.367
R1085 B.n500 B.n499 163.367
R1086 B.n500 B.n209 163.367
R1087 B.n504 B.n209 163.367
R1088 B.n505 B.n504 163.367
R1089 B.n506 B.n505 163.367
R1090 B.n506 B.n207 163.367
R1091 B.n510 B.n207 163.367
R1092 B.n511 B.n510 163.367
R1093 B.n512 B.n511 163.367
R1094 B.n512 B.n205 163.367
R1095 B.n516 B.n205 163.367
R1096 B.n517 B.n516 163.367
R1097 B.n518 B.n517 163.367
R1098 B.n518 B.n203 163.367
R1099 B.n522 B.n203 163.367
R1100 B.n523 B.n522 163.367
R1101 B.n524 B.n523 163.367
R1102 B.n524 B.n201 163.367
R1103 B.n528 B.n201 163.367
R1104 B.n529 B.n528 163.367
R1105 B.n530 B.n529 163.367
R1106 B.n530 B.n199 163.367
R1107 B.n534 B.n199 163.367
R1108 B.n535 B.n534 163.367
R1109 B.n536 B.n535 163.367
R1110 B.n536 B.n197 163.367
R1111 B.n540 B.n197 163.367
R1112 B.n541 B.n540 163.367
R1113 B.n542 B.n541 163.367
R1114 B.n542 B.n195 163.367
R1115 B.n546 B.n195 163.367
R1116 B.n547 B.n546 163.367
R1117 B.n548 B.n547 163.367
R1118 B.n548 B.n193 163.367
R1119 B.n552 B.n193 163.367
R1120 B.n553 B.n552 163.367
R1121 B.n554 B.n553 163.367
R1122 B.n554 B.n191 163.367
R1123 B.n558 B.n191 163.367
R1124 B.n559 B.n558 163.367
R1125 B.n560 B.n559 163.367
R1126 B.n560 B.n189 163.367
R1127 B.n564 B.n189 163.367
R1128 B.n565 B.n564 163.367
R1129 B.n566 B.n565 163.367
R1130 B.n566 B.n187 163.367
R1131 B.n570 B.n187 163.367
R1132 B.n824 B.n823 163.367
R1133 B.n823 B.n822 163.367
R1134 B.n822 B.n103 163.367
R1135 B.n818 B.n103 163.367
R1136 B.n818 B.n817 163.367
R1137 B.n817 B.n816 163.367
R1138 B.n816 B.n105 163.367
R1139 B.n812 B.n105 163.367
R1140 B.n812 B.n811 163.367
R1141 B.n811 B.n810 163.367
R1142 B.n810 B.n107 163.367
R1143 B.n806 B.n107 163.367
R1144 B.n806 B.n805 163.367
R1145 B.n805 B.n804 163.367
R1146 B.n804 B.n109 163.367
R1147 B.n800 B.n109 163.367
R1148 B.n800 B.n799 163.367
R1149 B.n799 B.n798 163.367
R1150 B.n798 B.n111 163.367
R1151 B.n794 B.n111 163.367
R1152 B.n794 B.n793 163.367
R1153 B.n793 B.n792 163.367
R1154 B.n792 B.n113 163.367
R1155 B.n788 B.n113 163.367
R1156 B.n788 B.n787 163.367
R1157 B.n787 B.n786 163.367
R1158 B.n786 B.n115 163.367
R1159 B.n782 B.n115 163.367
R1160 B.n782 B.n781 163.367
R1161 B.n781 B.n780 163.367
R1162 B.n780 B.n117 163.367
R1163 B.n776 B.n117 163.367
R1164 B.n776 B.n775 163.367
R1165 B.n775 B.n774 163.367
R1166 B.n774 B.n119 163.367
R1167 B.n770 B.n119 163.367
R1168 B.n770 B.n769 163.367
R1169 B.n769 B.n768 163.367
R1170 B.n768 B.n121 163.367
R1171 B.n764 B.n121 163.367
R1172 B.n764 B.n763 163.367
R1173 B.n763 B.n762 163.367
R1174 B.n762 B.n123 163.367
R1175 B.n758 B.n123 163.367
R1176 B.n758 B.n757 163.367
R1177 B.n757 B.n756 163.367
R1178 B.n756 B.n125 163.367
R1179 B.n752 B.n125 163.367
R1180 B.n752 B.n751 163.367
R1181 B.n751 B.n750 163.367
R1182 B.n750 B.n127 163.367
R1183 B.n746 B.n127 163.367
R1184 B.n746 B.n745 163.367
R1185 B.n745 B.n744 163.367
R1186 B.n744 B.n129 163.367
R1187 B.n740 B.n129 163.367
R1188 B.n740 B.n739 163.367
R1189 B.n739 B.n738 163.367
R1190 B.n738 B.n131 163.367
R1191 B.n734 B.n131 163.367
R1192 B.n734 B.n733 163.367
R1193 B.n733 B.n732 163.367
R1194 B.n732 B.n133 163.367
R1195 B.n728 B.n133 163.367
R1196 B.n728 B.n727 163.367
R1197 B.n727 B.n726 163.367
R1198 B.n726 B.n135 163.367
R1199 B.n722 B.n135 163.367
R1200 B.n722 B.n721 163.367
R1201 B.n721 B.n720 163.367
R1202 B.n720 B.n137 163.367
R1203 B.n716 B.n137 163.367
R1204 B.n716 B.n715 163.367
R1205 B.n715 B.n714 163.367
R1206 B.n714 B.n139 163.367
R1207 B.n710 B.n139 163.367
R1208 B.n710 B.n709 163.367
R1209 B.n709 B.n708 163.367
R1210 B.n708 B.n141 163.367
R1211 B.n704 B.n141 163.367
R1212 B.n704 B.n703 163.367
R1213 B.n703 B.n702 163.367
R1214 B.n702 B.n143 163.367
R1215 B.n698 B.n143 163.367
R1216 B.n698 B.n697 163.367
R1217 B.n697 B.n696 163.367
R1218 B.n696 B.n145 163.367
R1219 B.n692 B.n145 163.367
R1220 B.n692 B.n691 163.367
R1221 B.n691 B.n690 163.367
R1222 B.n690 B.n147 163.367
R1223 B.n686 B.n147 163.367
R1224 B.n686 B.n685 163.367
R1225 B.n685 B.n684 163.367
R1226 B.n684 B.n149 163.367
R1227 B.n680 B.n149 163.367
R1228 B.n680 B.n679 163.367
R1229 B.n679 B.n678 163.367
R1230 B.n678 B.n151 163.367
R1231 B.n674 B.n151 163.367
R1232 B.n674 B.n673 163.367
R1233 B.n673 B.n672 163.367
R1234 B.n672 B.n153 163.367
R1235 B.n668 B.n153 163.367
R1236 B.n668 B.n667 163.367
R1237 B.n667 B.n666 163.367
R1238 B.n666 B.n155 163.367
R1239 B.n662 B.n155 163.367
R1240 B.n662 B.n661 163.367
R1241 B.n661 B.n660 163.367
R1242 B.n660 B.n157 163.367
R1243 B.n656 B.n157 163.367
R1244 B.n656 B.n655 163.367
R1245 B.n655 B.n654 163.367
R1246 B.n654 B.n159 163.367
R1247 B.n650 B.n159 163.367
R1248 B.n650 B.n649 163.367
R1249 B.n649 B.n648 163.367
R1250 B.n648 B.n161 163.367
R1251 B.n644 B.n161 163.367
R1252 B.n644 B.n643 163.367
R1253 B.n643 B.n642 163.367
R1254 B.n642 B.n163 163.367
R1255 B.n638 B.n163 163.367
R1256 B.n638 B.n637 163.367
R1257 B.n637 B.n636 163.367
R1258 B.n636 B.n165 163.367
R1259 B.n632 B.n165 163.367
R1260 B.n632 B.n631 163.367
R1261 B.n631 B.n630 163.367
R1262 B.n630 B.n167 163.367
R1263 B.n626 B.n167 163.367
R1264 B.n626 B.n625 163.367
R1265 B.n625 B.n624 163.367
R1266 B.n624 B.n169 163.367
R1267 B.n620 B.n169 163.367
R1268 B.n620 B.n619 163.367
R1269 B.n619 B.n618 163.367
R1270 B.n618 B.n171 163.367
R1271 B.n614 B.n171 163.367
R1272 B.n614 B.n613 163.367
R1273 B.n613 B.n612 163.367
R1274 B.n612 B.n173 163.367
R1275 B.n608 B.n173 163.367
R1276 B.n608 B.n607 163.367
R1277 B.n607 B.n606 163.367
R1278 B.n606 B.n175 163.367
R1279 B.n602 B.n175 163.367
R1280 B.n602 B.n601 163.367
R1281 B.n601 B.n600 163.367
R1282 B.n600 B.n177 163.367
R1283 B.n596 B.n177 163.367
R1284 B.n596 B.n595 163.367
R1285 B.n595 B.n594 163.367
R1286 B.n594 B.n179 163.367
R1287 B.n590 B.n179 163.367
R1288 B.n590 B.n589 163.367
R1289 B.n589 B.n588 163.367
R1290 B.n588 B.n181 163.367
R1291 B.n584 B.n181 163.367
R1292 B.n584 B.n583 163.367
R1293 B.n583 B.n582 163.367
R1294 B.n582 B.n183 163.367
R1295 B.n578 B.n183 163.367
R1296 B.n578 B.n577 163.367
R1297 B.n577 B.n576 163.367
R1298 B.n576 B.n185 163.367
R1299 B.n572 B.n185 163.367
R1300 B.n572 B.n571 163.367
R1301 B.n985 B.n984 163.367
R1302 B.n984 B.n45 163.367
R1303 B.n980 B.n45 163.367
R1304 B.n980 B.n979 163.367
R1305 B.n979 B.n978 163.367
R1306 B.n978 B.n47 163.367
R1307 B.n974 B.n47 163.367
R1308 B.n974 B.n973 163.367
R1309 B.n973 B.n972 163.367
R1310 B.n972 B.n49 163.367
R1311 B.n968 B.n49 163.367
R1312 B.n968 B.n967 163.367
R1313 B.n967 B.n966 163.367
R1314 B.n966 B.n51 163.367
R1315 B.n962 B.n51 163.367
R1316 B.n962 B.n961 163.367
R1317 B.n961 B.n960 163.367
R1318 B.n960 B.n53 163.367
R1319 B.n956 B.n53 163.367
R1320 B.n956 B.n955 163.367
R1321 B.n955 B.n954 163.367
R1322 B.n954 B.n55 163.367
R1323 B.n950 B.n55 163.367
R1324 B.n950 B.n949 163.367
R1325 B.n949 B.n948 163.367
R1326 B.n948 B.n57 163.367
R1327 B.n944 B.n57 163.367
R1328 B.n944 B.n943 163.367
R1329 B.n943 B.n942 163.367
R1330 B.n942 B.n59 163.367
R1331 B.n938 B.n59 163.367
R1332 B.n938 B.n937 163.367
R1333 B.n937 B.n936 163.367
R1334 B.n936 B.n61 163.367
R1335 B.n932 B.n61 163.367
R1336 B.n932 B.n931 163.367
R1337 B.n931 B.n930 163.367
R1338 B.n930 B.n63 163.367
R1339 B.n926 B.n63 163.367
R1340 B.n926 B.n925 163.367
R1341 B.n925 B.n924 163.367
R1342 B.n924 B.n65 163.367
R1343 B.n920 B.n65 163.367
R1344 B.n920 B.n919 163.367
R1345 B.n919 B.n918 163.367
R1346 B.n918 B.n67 163.367
R1347 B.n914 B.n67 163.367
R1348 B.n914 B.n913 163.367
R1349 B.n913 B.n71 163.367
R1350 B.n909 B.n71 163.367
R1351 B.n909 B.n908 163.367
R1352 B.n908 B.n907 163.367
R1353 B.n907 B.n73 163.367
R1354 B.n903 B.n73 163.367
R1355 B.n903 B.n902 163.367
R1356 B.n902 B.n901 163.367
R1357 B.n901 B.n75 163.367
R1358 B.n896 B.n75 163.367
R1359 B.n896 B.n895 163.367
R1360 B.n895 B.n894 163.367
R1361 B.n894 B.n79 163.367
R1362 B.n890 B.n79 163.367
R1363 B.n890 B.n889 163.367
R1364 B.n889 B.n888 163.367
R1365 B.n888 B.n81 163.367
R1366 B.n884 B.n81 163.367
R1367 B.n884 B.n883 163.367
R1368 B.n883 B.n882 163.367
R1369 B.n882 B.n83 163.367
R1370 B.n878 B.n83 163.367
R1371 B.n878 B.n877 163.367
R1372 B.n877 B.n876 163.367
R1373 B.n876 B.n85 163.367
R1374 B.n872 B.n85 163.367
R1375 B.n872 B.n871 163.367
R1376 B.n871 B.n870 163.367
R1377 B.n870 B.n87 163.367
R1378 B.n866 B.n87 163.367
R1379 B.n866 B.n865 163.367
R1380 B.n865 B.n864 163.367
R1381 B.n864 B.n89 163.367
R1382 B.n860 B.n89 163.367
R1383 B.n860 B.n859 163.367
R1384 B.n859 B.n858 163.367
R1385 B.n858 B.n91 163.367
R1386 B.n854 B.n91 163.367
R1387 B.n854 B.n853 163.367
R1388 B.n853 B.n852 163.367
R1389 B.n852 B.n93 163.367
R1390 B.n848 B.n93 163.367
R1391 B.n848 B.n847 163.367
R1392 B.n847 B.n846 163.367
R1393 B.n846 B.n95 163.367
R1394 B.n842 B.n95 163.367
R1395 B.n842 B.n841 163.367
R1396 B.n841 B.n840 163.367
R1397 B.n840 B.n97 163.367
R1398 B.n836 B.n97 163.367
R1399 B.n836 B.n835 163.367
R1400 B.n835 B.n834 163.367
R1401 B.n834 B.n99 163.367
R1402 B.n830 B.n99 163.367
R1403 B.n830 B.n829 163.367
R1404 B.n829 B.n828 163.367
R1405 B.n828 B.n101 163.367
R1406 B.n986 B.n43 163.367
R1407 B.n990 B.n43 163.367
R1408 B.n991 B.n990 163.367
R1409 B.n992 B.n991 163.367
R1410 B.n992 B.n41 163.367
R1411 B.n996 B.n41 163.367
R1412 B.n997 B.n996 163.367
R1413 B.n998 B.n997 163.367
R1414 B.n998 B.n39 163.367
R1415 B.n1002 B.n39 163.367
R1416 B.n1003 B.n1002 163.367
R1417 B.n1004 B.n1003 163.367
R1418 B.n1004 B.n37 163.367
R1419 B.n1008 B.n37 163.367
R1420 B.n1009 B.n1008 163.367
R1421 B.n1010 B.n1009 163.367
R1422 B.n1010 B.n35 163.367
R1423 B.n1014 B.n35 163.367
R1424 B.n1015 B.n1014 163.367
R1425 B.n1016 B.n1015 163.367
R1426 B.n1016 B.n33 163.367
R1427 B.n1020 B.n33 163.367
R1428 B.n1021 B.n1020 163.367
R1429 B.n1022 B.n1021 163.367
R1430 B.n1022 B.n31 163.367
R1431 B.n1026 B.n31 163.367
R1432 B.n1027 B.n1026 163.367
R1433 B.n1028 B.n1027 163.367
R1434 B.n1028 B.n29 163.367
R1435 B.n1032 B.n29 163.367
R1436 B.n1033 B.n1032 163.367
R1437 B.n1034 B.n1033 163.367
R1438 B.n1034 B.n27 163.367
R1439 B.n1038 B.n27 163.367
R1440 B.n1039 B.n1038 163.367
R1441 B.n1040 B.n1039 163.367
R1442 B.n1040 B.n25 163.367
R1443 B.n1044 B.n25 163.367
R1444 B.n1045 B.n1044 163.367
R1445 B.n1046 B.n1045 163.367
R1446 B.n1046 B.n23 163.367
R1447 B.n1050 B.n23 163.367
R1448 B.n1051 B.n1050 163.367
R1449 B.n1052 B.n1051 163.367
R1450 B.n1052 B.n21 163.367
R1451 B.n1056 B.n21 163.367
R1452 B.n1057 B.n1056 163.367
R1453 B.n1058 B.n1057 163.367
R1454 B.n1058 B.n19 163.367
R1455 B.n1062 B.n19 163.367
R1456 B.n1063 B.n1062 163.367
R1457 B.n1064 B.n1063 163.367
R1458 B.n1064 B.n17 163.367
R1459 B.n1068 B.n17 163.367
R1460 B.n1069 B.n1068 163.367
R1461 B.n1070 B.n1069 163.367
R1462 B.n1070 B.n15 163.367
R1463 B.n1074 B.n15 163.367
R1464 B.n1075 B.n1074 163.367
R1465 B.n1076 B.n1075 163.367
R1466 B.n1076 B.n13 163.367
R1467 B.n1080 B.n13 163.367
R1468 B.n1081 B.n1080 163.367
R1469 B.n1082 B.n1081 163.367
R1470 B.n1082 B.n11 163.367
R1471 B.n1086 B.n11 163.367
R1472 B.n1087 B.n1086 163.367
R1473 B.n1088 B.n1087 163.367
R1474 B.n1088 B.n9 163.367
R1475 B.n1092 B.n9 163.367
R1476 B.n1093 B.n1092 163.367
R1477 B.n1094 B.n1093 163.367
R1478 B.n1094 B.n7 163.367
R1479 B.n1098 B.n7 163.367
R1480 B.n1099 B.n1098 163.367
R1481 B.n1100 B.n1099 163.367
R1482 B.n1100 B.n5 163.367
R1483 B.n1104 B.n5 163.367
R1484 B.n1105 B.n1104 163.367
R1485 B.n1106 B.n1105 163.367
R1486 B.n1106 B.n3 163.367
R1487 B.n1110 B.n3 163.367
R1488 B.n1111 B.n1110 163.367
R1489 B.n284 B.n2 163.367
R1490 B.n285 B.n284 163.367
R1491 B.n286 B.n285 163.367
R1492 B.n286 B.n281 163.367
R1493 B.n290 B.n281 163.367
R1494 B.n291 B.n290 163.367
R1495 B.n292 B.n291 163.367
R1496 B.n292 B.n279 163.367
R1497 B.n296 B.n279 163.367
R1498 B.n297 B.n296 163.367
R1499 B.n298 B.n297 163.367
R1500 B.n298 B.n277 163.367
R1501 B.n302 B.n277 163.367
R1502 B.n303 B.n302 163.367
R1503 B.n304 B.n303 163.367
R1504 B.n304 B.n275 163.367
R1505 B.n308 B.n275 163.367
R1506 B.n309 B.n308 163.367
R1507 B.n310 B.n309 163.367
R1508 B.n310 B.n273 163.367
R1509 B.n314 B.n273 163.367
R1510 B.n315 B.n314 163.367
R1511 B.n316 B.n315 163.367
R1512 B.n316 B.n271 163.367
R1513 B.n320 B.n271 163.367
R1514 B.n321 B.n320 163.367
R1515 B.n322 B.n321 163.367
R1516 B.n322 B.n269 163.367
R1517 B.n326 B.n269 163.367
R1518 B.n327 B.n326 163.367
R1519 B.n328 B.n327 163.367
R1520 B.n328 B.n267 163.367
R1521 B.n332 B.n267 163.367
R1522 B.n333 B.n332 163.367
R1523 B.n334 B.n333 163.367
R1524 B.n334 B.n265 163.367
R1525 B.n338 B.n265 163.367
R1526 B.n339 B.n338 163.367
R1527 B.n340 B.n339 163.367
R1528 B.n340 B.n263 163.367
R1529 B.n344 B.n263 163.367
R1530 B.n345 B.n344 163.367
R1531 B.n346 B.n345 163.367
R1532 B.n346 B.n261 163.367
R1533 B.n350 B.n261 163.367
R1534 B.n351 B.n350 163.367
R1535 B.n352 B.n351 163.367
R1536 B.n352 B.n259 163.367
R1537 B.n356 B.n259 163.367
R1538 B.n357 B.n356 163.367
R1539 B.n358 B.n357 163.367
R1540 B.n358 B.n257 163.367
R1541 B.n362 B.n257 163.367
R1542 B.n363 B.n362 163.367
R1543 B.n364 B.n363 163.367
R1544 B.n364 B.n255 163.367
R1545 B.n368 B.n255 163.367
R1546 B.n369 B.n368 163.367
R1547 B.n370 B.n369 163.367
R1548 B.n370 B.n253 163.367
R1549 B.n374 B.n253 163.367
R1550 B.n375 B.n374 163.367
R1551 B.n376 B.n375 163.367
R1552 B.n376 B.n251 163.367
R1553 B.n380 B.n251 163.367
R1554 B.n381 B.n380 163.367
R1555 B.n382 B.n381 163.367
R1556 B.n382 B.n249 163.367
R1557 B.n386 B.n249 163.367
R1558 B.n387 B.n386 163.367
R1559 B.n388 B.n387 163.367
R1560 B.n388 B.n247 163.367
R1561 B.n392 B.n247 163.367
R1562 B.n393 B.n392 163.367
R1563 B.n394 B.n393 163.367
R1564 B.n394 B.n245 163.367
R1565 B.n398 B.n245 163.367
R1566 B.n399 B.n398 163.367
R1567 B.n400 B.n399 163.367
R1568 B.n400 B.n243 163.367
R1569 B.n404 B.n243 163.367
R1570 B.n405 B.n404 163.367
R1571 B.n406 B.n405 163.367
R1572 B.n495 B.t11 106.862
R1573 B.n77 B.t7 106.862
R1574 B.n217 B.t2 106.844
R1575 B.n69 B.t4 106.844
R1576 B.n217 B.n216 83.9763
R1577 B.n495 B.n494 83.9763
R1578 B.n77 B.n76 83.9763
R1579 B.n69 B.n68 83.9763
R1580 B.n480 B.n217 59.5399
R1581 B.n496 B.n495 59.5399
R1582 B.n898 B.n77 59.5399
R1583 B.n70 B.n69 59.5399
R1584 B.n987 B.n44 34.1859
R1585 B.n826 B.n825 34.1859
R1586 B.n569 B.n186 34.1859
R1587 B.n408 B.n407 34.1859
R1588 B B.n1113 18.0485
R1589 B.n988 B.n987 10.6151
R1590 B.n989 B.n988 10.6151
R1591 B.n989 B.n42 10.6151
R1592 B.n993 B.n42 10.6151
R1593 B.n994 B.n993 10.6151
R1594 B.n995 B.n994 10.6151
R1595 B.n995 B.n40 10.6151
R1596 B.n999 B.n40 10.6151
R1597 B.n1000 B.n999 10.6151
R1598 B.n1001 B.n1000 10.6151
R1599 B.n1001 B.n38 10.6151
R1600 B.n1005 B.n38 10.6151
R1601 B.n1006 B.n1005 10.6151
R1602 B.n1007 B.n1006 10.6151
R1603 B.n1007 B.n36 10.6151
R1604 B.n1011 B.n36 10.6151
R1605 B.n1012 B.n1011 10.6151
R1606 B.n1013 B.n1012 10.6151
R1607 B.n1013 B.n34 10.6151
R1608 B.n1017 B.n34 10.6151
R1609 B.n1018 B.n1017 10.6151
R1610 B.n1019 B.n1018 10.6151
R1611 B.n1019 B.n32 10.6151
R1612 B.n1023 B.n32 10.6151
R1613 B.n1024 B.n1023 10.6151
R1614 B.n1025 B.n1024 10.6151
R1615 B.n1025 B.n30 10.6151
R1616 B.n1029 B.n30 10.6151
R1617 B.n1030 B.n1029 10.6151
R1618 B.n1031 B.n1030 10.6151
R1619 B.n1031 B.n28 10.6151
R1620 B.n1035 B.n28 10.6151
R1621 B.n1036 B.n1035 10.6151
R1622 B.n1037 B.n1036 10.6151
R1623 B.n1037 B.n26 10.6151
R1624 B.n1041 B.n26 10.6151
R1625 B.n1042 B.n1041 10.6151
R1626 B.n1043 B.n1042 10.6151
R1627 B.n1043 B.n24 10.6151
R1628 B.n1047 B.n24 10.6151
R1629 B.n1048 B.n1047 10.6151
R1630 B.n1049 B.n1048 10.6151
R1631 B.n1049 B.n22 10.6151
R1632 B.n1053 B.n22 10.6151
R1633 B.n1054 B.n1053 10.6151
R1634 B.n1055 B.n1054 10.6151
R1635 B.n1055 B.n20 10.6151
R1636 B.n1059 B.n20 10.6151
R1637 B.n1060 B.n1059 10.6151
R1638 B.n1061 B.n1060 10.6151
R1639 B.n1061 B.n18 10.6151
R1640 B.n1065 B.n18 10.6151
R1641 B.n1066 B.n1065 10.6151
R1642 B.n1067 B.n1066 10.6151
R1643 B.n1067 B.n16 10.6151
R1644 B.n1071 B.n16 10.6151
R1645 B.n1072 B.n1071 10.6151
R1646 B.n1073 B.n1072 10.6151
R1647 B.n1073 B.n14 10.6151
R1648 B.n1077 B.n14 10.6151
R1649 B.n1078 B.n1077 10.6151
R1650 B.n1079 B.n1078 10.6151
R1651 B.n1079 B.n12 10.6151
R1652 B.n1083 B.n12 10.6151
R1653 B.n1084 B.n1083 10.6151
R1654 B.n1085 B.n1084 10.6151
R1655 B.n1085 B.n10 10.6151
R1656 B.n1089 B.n10 10.6151
R1657 B.n1090 B.n1089 10.6151
R1658 B.n1091 B.n1090 10.6151
R1659 B.n1091 B.n8 10.6151
R1660 B.n1095 B.n8 10.6151
R1661 B.n1096 B.n1095 10.6151
R1662 B.n1097 B.n1096 10.6151
R1663 B.n1097 B.n6 10.6151
R1664 B.n1101 B.n6 10.6151
R1665 B.n1102 B.n1101 10.6151
R1666 B.n1103 B.n1102 10.6151
R1667 B.n1103 B.n4 10.6151
R1668 B.n1107 B.n4 10.6151
R1669 B.n1108 B.n1107 10.6151
R1670 B.n1109 B.n1108 10.6151
R1671 B.n1109 B.n0 10.6151
R1672 B.n983 B.n44 10.6151
R1673 B.n983 B.n982 10.6151
R1674 B.n982 B.n981 10.6151
R1675 B.n981 B.n46 10.6151
R1676 B.n977 B.n46 10.6151
R1677 B.n977 B.n976 10.6151
R1678 B.n976 B.n975 10.6151
R1679 B.n975 B.n48 10.6151
R1680 B.n971 B.n48 10.6151
R1681 B.n971 B.n970 10.6151
R1682 B.n970 B.n969 10.6151
R1683 B.n969 B.n50 10.6151
R1684 B.n965 B.n50 10.6151
R1685 B.n965 B.n964 10.6151
R1686 B.n964 B.n963 10.6151
R1687 B.n963 B.n52 10.6151
R1688 B.n959 B.n52 10.6151
R1689 B.n959 B.n958 10.6151
R1690 B.n958 B.n957 10.6151
R1691 B.n957 B.n54 10.6151
R1692 B.n953 B.n54 10.6151
R1693 B.n953 B.n952 10.6151
R1694 B.n952 B.n951 10.6151
R1695 B.n951 B.n56 10.6151
R1696 B.n947 B.n56 10.6151
R1697 B.n947 B.n946 10.6151
R1698 B.n946 B.n945 10.6151
R1699 B.n945 B.n58 10.6151
R1700 B.n941 B.n58 10.6151
R1701 B.n941 B.n940 10.6151
R1702 B.n940 B.n939 10.6151
R1703 B.n939 B.n60 10.6151
R1704 B.n935 B.n60 10.6151
R1705 B.n935 B.n934 10.6151
R1706 B.n934 B.n933 10.6151
R1707 B.n933 B.n62 10.6151
R1708 B.n929 B.n62 10.6151
R1709 B.n929 B.n928 10.6151
R1710 B.n928 B.n927 10.6151
R1711 B.n927 B.n64 10.6151
R1712 B.n923 B.n64 10.6151
R1713 B.n923 B.n922 10.6151
R1714 B.n922 B.n921 10.6151
R1715 B.n921 B.n66 10.6151
R1716 B.n917 B.n66 10.6151
R1717 B.n917 B.n916 10.6151
R1718 B.n916 B.n915 10.6151
R1719 B.n912 B.n911 10.6151
R1720 B.n911 B.n910 10.6151
R1721 B.n910 B.n72 10.6151
R1722 B.n906 B.n72 10.6151
R1723 B.n906 B.n905 10.6151
R1724 B.n905 B.n904 10.6151
R1725 B.n904 B.n74 10.6151
R1726 B.n900 B.n74 10.6151
R1727 B.n900 B.n899 10.6151
R1728 B.n897 B.n78 10.6151
R1729 B.n893 B.n78 10.6151
R1730 B.n893 B.n892 10.6151
R1731 B.n892 B.n891 10.6151
R1732 B.n891 B.n80 10.6151
R1733 B.n887 B.n80 10.6151
R1734 B.n887 B.n886 10.6151
R1735 B.n886 B.n885 10.6151
R1736 B.n885 B.n82 10.6151
R1737 B.n881 B.n82 10.6151
R1738 B.n881 B.n880 10.6151
R1739 B.n880 B.n879 10.6151
R1740 B.n879 B.n84 10.6151
R1741 B.n875 B.n84 10.6151
R1742 B.n875 B.n874 10.6151
R1743 B.n874 B.n873 10.6151
R1744 B.n873 B.n86 10.6151
R1745 B.n869 B.n86 10.6151
R1746 B.n869 B.n868 10.6151
R1747 B.n868 B.n867 10.6151
R1748 B.n867 B.n88 10.6151
R1749 B.n863 B.n88 10.6151
R1750 B.n863 B.n862 10.6151
R1751 B.n862 B.n861 10.6151
R1752 B.n861 B.n90 10.6151
R1753 B.n857 B.n90 10.6151
R1754 B.n857 B.n856 10.6151
R1755 B.n856 B.n855 10.6151
R1756 B.n855 B.n92 10.6151
R1757 B.n851 B.n92 10.6151
R1758 B.n851 B.n850 10.6151
R1759 B.n850 B.n849 10.6151
R1760 B.n849 B.n94 10.6151
R1761 B.n845 B.n94 10.6151
R1762 B.n845 B.n844 10.6151
R1763 B.n844 B.n843 10.6151
R1764 B.n843 B.n96 10.6151
R1765 B.n839 B.n96 10.6151
R1766 B.n839 B.n838 10.6151
R1767 B.n838 B.n837 10.6151
R1768 B.n837 B.n98 10.6151
R1769 B.n833 B.n98 10.6151
R1770 B.n833 B.n832 10.6151
R1771 B.n832 B.n831 10.6151
R1772 B.n831 B.n100 10.6151
R1773 B.n827 B.n100 10.6151
R1774 B.n827 B.n826 10.6151
R1775 B.n825 B.n102 10.6151
R1776 B.n821 B.n102 10.6151
R1777 B.n821 B.n820 10.6151
R1778 B.n820 B.n819 10.6151
R1779 B.n819 B.n104 10.6151
R1780 B.n815 B.n104 10.6151
R1781 B.n815 B.n814 10.6151
R1782 B.n814 B.n813 10.6151
R1783 B.n813 B.n106 10.6151
R1784 B.n809 B.n106 10.6151
R1785 B.n809 B.n808 10.6151
R1786 B.n808 B.n807 10.6151
R1787 B.n807 B.n108 10.6151
R1788 B.n803 B.n108 10.6151
R1789 B.n803 B.n802 10.6151
R1790 B.n802 B.n801 10.6151
R1791 B.n801 B.n110 10.6151
R1792 B.n797 B.n110 10.6151
R1793 B.n797 B.n796 10.6151
R1794 B.n796 B.n795 10.6151
R1795 B.n795 B.n112 10.6151
R1796 B.n791 B.n112 10.6151
R1797 B.n791 B.n790 10.6151
R1798 B.n790 B.n789 10.6151
R1799 B.n789 B.n114 10.6151
R1800 B.n785 B.n114 10.6151
R1801 B.n785 B.n784 10.6151
R1802 B.n784 B.n783 10.6151
R1803 B.n783 B.n116 10.6151
R1804 B.n779 B.n116 10.6151
R1805 B.n779 B.n778 10.6151
R1806 B.n778 B.n777 10.6151
R1807 B.n777 B.n118 10.6151
R1808 B.n773 B.n118 10.6151
R1809 B.n773 B.n772 10.6151
R1810 B.n772 B.n771 10.6151
R1811 B.n771 B.n120 10.6151
R1812 B.n767 B.n120 10.6151
R1813 B.n767 B.n766 10.6151
R1814 B.n766 B.n765 10.6151
R1815 B.n765 B.n122 10.6151
R1816 B.n761 B.n122 10.6151
R1817 B.n761 B.n760 10.6151
R1818 B.n760 B.n759 10.6151
R1819 B.n759 B.n124 10.6151
R1820 B.n755 B.n124 10.6151
R1821 B.n755 B.n754 10.6151
R1822 B.n754 B.n753 10.6151
R1823 B.n753 B.n126 10.6151
R1824 B.n749 B.n126 10.6151
R1825 B.n749 B.n748 10.6151
R1826 B.n748 B.n747 10.6151
R1827 B.n747 B.n128 10.6151
R1828 B.n743 B.n128 10.6151
R1829 B.n743 B.n742 10.6151
R1830 B.n742 B.n741 10.6151
R1831 B.n741 B.n130 10.6151
R1832 B.n737 B.n130 10.6151
R1833 B.n737 B.n736 10.6151
R1834 B.n736 B.n735 10.6151
R1835 B.n735 B.n132 10.6151
R1836 B.n731 B.n132 10.6151
R1837 B.n731 B.n730 10.6151
R1838 B.n730 B.n729 10.6151
R1839 B.n729 B.n134 10.6151
R1840 B.n725 B.n134 10.6151
R1841 B.n725 B.n724 10.6151
R1842 B.n724 B.n723 10.6151
R1843 B.n723 B.n136 10.6151
R1844 B.n719 B.n136 10.6151
R1845 B.n719 B.n718 10.6151
R1846 B.n718 B.n717 10.6151
R1847 B.n717 B.n138 10.6151
R1848 B.n713 B.n138 10.6151
R1849 B.n713 B.n712 10.6151
R1850 B.n712 B.n711 10.6151
R1851 B.n711 B.n140 10.6151
R1852 B.n707 B.n140 10.6151
R1853 B.n707 B.n706 10.6151
R1854 B.n706 B.n705 10.6151
R1855 B.n705 B.n142 10.6151
R1856 B.n701 B.n142 10.6151
R1857 B.n701 B.n700 10.6151
R1858 B.n700 B.n699 10.6151
R1859 B.n699 B.n144 10.6151
R1860 B.n695 B.n144 10.6151
R1861 B.n695 B.n694 10.6151
R1862 B.n694 B.n693 10.6151
R1863 B.n693 B.n146 10.6151
R1864 B.n689 B.n146 10.6151
R1865 B.n689 B.n688 10.6151
R1866 B.n688 B.n687 10.6151
R1867 B.n687 B.n148 10.6151
R1868 B.n683 B.n148 10.6151
R1869 B.n683 B.n682 10.6151
R1870 B.n682 B.n681 10.6151
R1871 B.n681 B.n150 10.6151
R1872 B.n677 B.n150 10.6151
R1873 B.n677 B.n676 10.6151
R1874 B.n676 B.n675 10.6151
R1875 B.n675 B.n152 10.6151
R1876 B.n671 B.n152 10.6151
R1877 B.n671 B.n670 10.6151
R1878 B.n670 B.n669 10.6151
R1879 B.n669 B.n154 10.6151
R1880 B.n665 B.n154 10.6151
R1881 B.n665 B.n664 10.6151
R1882 B.n664 B.n663 10.6151
R1883 B.n663 B.n156 10.6151
R1884 B.n659 B.n156 10.6151
R1885 B.n659 B.n658 10.6151
R1886 B.n658 B.n657 10.6151
R1887 B.n657 B.n158 10.6151
R1888 B.n653 B.n158 10.6151
R1889 B.n653 B.n652 10.6151
R1890 B.n652 B.n651 10.6151
R1891 B.n651 B.n160 10.6151
R1892 B.n647 B.n160 10.6151
R1893 B.n647 B.n646 10.6151
R1894 B.n646 B.n645 10.6151
R1895 B.n645 B.n162 10.6151
R1896 B.n641 B.n162 10.6151
R1897 B.n641 B.n640 10.6151
R1898 B.n640 B.n639 10.6151
R1899 B.n639 B.n164 10.6151
R1900 B.n635 B.n164 10.6151
R1901 B.n635 B.n634 10.6151
R1902 B.n634 B.n633 10.6151
R1903 B.n633 B.n166 10.6151
R1904 B.n629 B.n166 10.6151
R1905 B.n629 B.n628 10.6151
R1906 B.n628 B.n627 10.6151
R1907 B.n627 B.n168 10.6151
R1908 B.n623 B.n168 10.6151
R1909 B.n623 B.n622 10.6151
R1910 B.n622 B.n621 10.6151
R1911 B.n621 B.n170 10.6151
R1912 B.n617 B.n170 10.6151
R1913 B.n617 B.n616 10.6151
R1914 B.n616 B.n615 10.6151
R1915 B.n615 B.n172 10.6151
R1916 B.n611 B.n172 10.6151
R1917 B.n611 B.n610 10.6151
R1918 B.n610 B.n609 10.6151
R1919 B.n609 B.n174 10.6151
R1920 B.n605 B.n174 10.6151
R1921 B.n605 B.n604 10.6151
R1922 B.n604 B.n603 10.6151
R1923 B.n603 B.n176 10.6151
R1924 B.n599 B.n176 10.6151
R1925 B.n599 B.n598 10.6151
R1926 B.n598 B.n597 10.6151
R1927 B.n597 B.n178 10.6151
R1928 B.n593 B.n178 10.6151
R1929 B.n593 B.n592 10.6151
R1930 B.n592 B.n591 10.6151
R1931 B.n591 B.n180 10.6151
R1932 B.n587 B.n180 10.6151
R1933 B.n587 B.n586 10.6151
R1934 B.n586 B.n585 10.6151
R1935 B.n585 B.n182 10.6151
R1936 B.n581 B.n182 10.6151
R1937 B.n581 B.n580 10.6151
R1938 B.n580 B.n579 10.6151
R1939 B.n579 B.n184 10.6151
R1940 B.n575 B.n184 10.6151
R1941 B.n575 B.n574 10.6151
R1942 B.n574 B.n573 10.6151
R1943 B.n573 B.n186 10.6151
R1944 B.n283 B.n1 10.6151
R1945 B.n283 B.n282 10.6151
R1946 B.n287 B.n282 10.6151
R1947 B.n288 B.n287 10.6151
R1948 B.n289 B.n288 10.6151
R1949 B.n289 B.n280 10.6151
R1950 B.n293 B.n280 10.6151
R1951 B.n294 B.n293 10.6151
R1952 B.n295 B.n294 10.6151
R1953 B.n295 B.n278 10.6151
R1954 B.n299 B.n278 10.6151
R1955 B.n300 B.n299 10.6151
R1956 B.n301 B.n300 10.6151
R1957 B.n301 B.n276 10.6151
R1958 B.n305 B.n276 10.6151
R1959 B.n306 B.n305 10.6151
R1960 B.n307 B.n306 10.6151
R1961 B.n307 B.n274 10.6151
R1962 B.n311 B.n274 10.6151
R1963 B.n312 B.n311 10.6151
R1964 B.n313 B.n312 10.6151
R1965 B.n313 B.n272 10.6151
R1966 B.n317 B.n272 10.6151
R1967 B.n318 B.n317 10.6151
R1968 B.n319 B.n318 10.6151
R1969 B.n319 B.n270 10.6151
R1970 B.n323 B.n270 10.6151
R1971 B.n324 B.n323 10.6151
R1972 B.n325 B.n324 10.6151
R1973 B.n325 B.n268 10.6151
R1974 B.n329 B.n268 10.6151
R1975 B.n330 B.n329 10.6151
R1976 B.n331 B.n330 10.6151
R1977 B.n331 B.n266 10.6151
R1978 B.n335 B.n266 10.6151
R1979 B.n336 B.n335 10.6151
R1980 B.n337 B.n336 10.6151
R1981 B.n337 B.n264 10.6151
R1982 B.n341 B.n264 10.6151
R1983 B.n342 B.n341 10.6151
R1984 B.n343 B.n342 10.6151
R1985 B.n343 B.n262 10.6151
R1986 B.n347 B.n262 10.6151
R1987 B.n348 B.n347 10.6151
R1988 B.n349 B.n348 10.6151
R1989 B.n349 B.n260 10.6151
R1990 B.n353 B.n260 10.6151
R1991 B.n354 B.n353 10.6151
R1992 B.n355 B.n354 10.6151
R1993 B.n355 B.n258 10.6151
R1994 B.n359 B.n258 10.6151
R1995 B.n360 B.n359 10.6151
R1996 B.n361 B.n360 10.6151
R1997 B.n361 B.n256 10.6151
R1998 B.n365 B.n256 10.6151
R1999 B.n366 B.n365 10.6151
R2000 B.n367 B.n366 10.6151
R2001 B.n367 B.n254 10.6151
R2002 B.n371 B.n254 10.6151
R2003 B.n372 B.n371 10.6151
R2004 B.n373 B.n372 10.6151
R2005 B.n373 B.n252 10.6151
R2006 B.n377 B.n252 10.6151
R2007 B.n378 B.n377 10.6151
R2008 B.n379 B.n378 10.6151
R2009 B.n379 B.n250 10.6151
R2010 B.n383 B.n250 10.6151
R2011 B.n384 B.n383 10.6151
R2012 B.n385 B.n384 10.6151
R2013 B.n385 B.n248 10.6151
R2014 B.n389 B.n248 10.6151
R2015 B.n390 B.n389 10.6151
R2016 B.n391 B.n390 10.6151
R2017 B.n391 B.n246 10.6151
R2018 B.n395 B.n246 10.6151
R2019 B.n396 B.n395 10.6151
R2020 B.n397 B.n396 10.6151
R2021 B.n397 B.n244 10.6151
R2022 B.n401 B.n244 10.6151
R2023 B.n402 B.n401 10.6151
R2024 B.n403 B.n402 10.6151
R2025 B.n403 B.n242 10.6151
R2026 B.n407 B.n242 10.6151
R2027 B.n409 B.n408 10.6151
R2028 B.n409 B.n240 10.6151
R2029 B.n413 B.n240 10.6151
R2030 B.n414 B.n413 10.6151
R2031 B.n415 B.n414 10.6151
R2032 B.n415 B.n238 10.6151
R2033 B.n419 B.n238 10.6151
R2034 B.n420 B.n419 10.6151
R2035 B.n421 B.n420 10.6151
R2036 B.n421 B.n236 10.6151
R2037 B.n425 B.n236 10.6151
R2038 B.n426 B.n425 10.6151
R2039 B.n427 B.n426 10.6151
R2040 B.n427 B.n234 10.6151
R2041 B.n431 B.n234 10.6151
R2042 B.n432 B.n431 10.6151
R2043 B.n433 B.n432 10.6151
R2044 B.n433 B.n232 10.6151
R2045 B.n437 B.n232 10.6151
R2046 B.n438 B.n437 10.6151
R2047 B.n439 B.n438 10.6151
R2048 B.n439 B.n230 10.6151
R2049 B.n443 B.n230 10.6151
R2050 B.n444 B.n443 10.6151
R2051 B.n445 B.n444 10.6151
R2052 B.n445 B.n228 10.6151
R2053 B.n449 B.n228 10.6151
R2054 B.n450 B.n449 10.6151
R2055 B.n451 B.n450 10.6151
R2056 B.n451 B.n226 10.6151
R2057 B.n455 B.n226 10.6151
R2058 B.n456 B.n455 10.6151
R2059 B.n457 B.n456 10.6151
R2060 B.n457 B.n224 10.6151
R2061 B.n461 B.n224 10.6151
R2062 B.n462 B.n461 10.6151
R2063 B.n463 B.n462 10.6151
R2064 B.n463 B.n222 10.6151
R2065 B.n467 B.n222 10.6151
R2066 B.n468 B.n467 10.6151
R2067 B.n469 B.n468 10.6151
R2068 B.n469 B.n220 10.6151
R2069 B.n473 B.n220 10.6151
R2070 B.n474 B.n473 10.6151
R2071 B.n475 B.n474 10.6151
R2072 B.n475 B.n218 10.6151
R2073 B.n479 B.n218 10.6151
R2074 B.n482 B.n481 10.6151
R2075 B.n482 B.n214 10.6151
R2076 B.n486 B.n214 10.6151
R2077 B.n487 B.n486 10.6151
R2078 B.n488 B.n487 10.6151
R2079 B.n488 B.n212 10.6151
R2080 B.n492 B.n212 10.6151
R2081 B.n493 B.n492 10.6151
R2082 B.n497 B.n493 10.6151
R2083 B.n501 B.n210 10.6151
R2084 B.n502 B.n501 10.6151
R2085 B.n503 B.n502 10.6151
R2086 B.n503 B.n208 10.6151
R2087 B.n507 B.n208 10.6151
R2088 B.n508 B.n507 10.6151
R2089 B.n509 B.n508 10.6151
R2090 B.n509 B.n206 10.6151
R2091 B.n513 B.n206 10.6151
R2092 B.n514 B.n513 10.6151
R2093 B.n515 B.n514 10.6151
R2094 B.n515 B.n204 10.6151
R2095 B.n519 B.n204 10.6151
R2096 B.n520 B.n519 10.6151
R2097 B.n521 B.n520 10.6151
R2098 B.n521 B.n202 10.6151
R2099 B.n525 B.n202 10.6151
R2100 B.n526 B.n525 10.6151
R2101 B.n527 B.n526 10.6151
R2102 B.n527 B.n200 10.6151
R2103 B.n531 B.n200 10.6151
R2104 B.n532 B.n531 10.6151
R2105 B.n533 B.n532 10.6151
R2106 B.n533 B.n198 10.6151
R2107 B.n537 B.n198 10.6151
R2108 B.n538 B.n537 10.6151
R2109 B.n539 B.n538 10.6151
R2110 B.n539 B.n196 10.6151
R2111 B.n543 B.n196 10.6151
R2112 B.n544 B.n543 10.6151
R2113 B.n545 B.n544 10.6151
R2114 B.n545 B.n194 10.6151
R2115 B.n549 B.n194 10.6151
R2116 B.n550 B.n549 10.6151
R2117 B.n551 B.n550 10.6151
R2118 B.n551 B.n192 10.6151
R2119 B.n555 B.n192 10.6151
R2120 B.n556 B.n555 10.6151
R2121 B.n557 B.n556 10.6151
R2122 B.n557 B.n190 10.6151
R2123 B.n561 B.n190 10.6151
R2124 B.n562 B.n561 10.6151
R2125 B.n563 B.n562 10.6151
R2126 B.n563 B.n188 10.6151
R2127 B.n567 B.n188 10.6151
R2128 B.n568 B.n567 10.6151
R2129 B.n569 B.n568 10.6151
R2130 B.n915 B.n70 9.36635
R2131 B.n898 B.n897 9.36635
R2132 B.n480 B.n479 9.36635
R2133 B.n496 B.n210 9.36635
R2134 B.n1113 B.n0 8.11757
R2135 B.n1113 B.n1 8.11757
R2136 B.n912 B.n70 1.24928
R2137 B.n899 B.n898 1.24928
R2138 B.n481 B.n480 1.24928
R2139 B.n497 B.n496 1.24928
C0 VP w_n6166_n3826# 14.467599f
C1 B w_n6166_n3826# 13.5423f
C2 VTAIL w_n6166_n3826# 3.71806f
C3 B VP 3.03129f
C4 VTAIL VP 14.679199f
C5 VDD1 w_n6166_n3826# 3.47095f
C6 B VTAIL 4.80106f
C7 VDD2 w_n6166_n3826# 3.68726f
C8 VDD1 VP 14.1342f
C9 B VDD1 3.20832f
C10 VDD2 VP 0.761612f
C11 VDD1 VTAIL 12.0321f
C12 B VDD2 3.38076f
C13 VDD2 VTAIL 12.093201f
C14 VDD2 VDD1 3.08704f
C15 VN w_n6166_n3826# 13.660501f
C16 VN VP 10.889299f
C17 VN B 1.66638f
C18 VN VTAIL 14.6642f
C19 VN VDD1 0.156594f
C20 VN VDD2 13.5327f
C21 VDD2 VSUBS 2.73339f
C22 VDD1 VSUBS 2.613298f
C23 VTAIL VSUBS 1.714535f
C24 VN VSUBS 10.121189f
C25 VP VSUBS 6.120035f
C26 B VSUBS 7.294182f
C27 w_n6166_n3826# VSUBS 0.289531p
C28 B.n0 VSUBS 0.00719f
C29 B.n1 VSUBS 0.00719f
C30 B.n2 VSUBS 0.010633f
C31 B.n3 VSUBS 0.008148f
C32 B.n4 VSUBS 0.008148f
C33 B.n5 VSUBS 0.008148f
C34 B.n6 VSUBS 0.008148f
C35 B.n7 VSUBS 0.008148f
C36 B.n8 VSUBS 0.008148f
C37 B.n9 VSUBS 0.008148f
C38 B.n10 VSUBS 0.008148f
C39 B.n11 VSUBS 0.008148f
C40 B.n12 VSUBS 0.008148f
C41 B.n13 VSUBS 0.008148f
C42 B.n14 VSUBS 0.008148f
C43 B.n15 VSUBS 0.008148f
C44 B.n16 VSUBS 0.008148f
C45 B.n17 VSUBS 0.008148f
C46 B.n18 VSUBS 0.008148f
C47 B.n19 VSUBS 0.008148f
C48 B.n20 VSUBS 0.008148f
C49 B.n21 VSUBS 0.008148f
C50 B.n22 VSUBS 0.008148f
C51 B.n23 VSUBS 0.008148f
C52 B.n24 VSUBS 0.008148f
C53 B.n25 VSUBS 0.008148f
C54 B.n26 VSUBS 0.008148f
C55 B.n27 VSUBS 0.008148f
C56 B.n28 VSUBS 0.008148f
C57 B.n29 VSUBS 0.008148f
C58 B.n30 VSUBS 0.008148f
C59 B.n31 VSUBS 0.008148f
C60 B.n32 VSUBS 0.008148f
C61 B.n33 VSUBS 0.008148f
C62 B.n34 VSUBS 0.008148f
C63 B.n35 VSUBS 0.008148f
C64 B.n36 VSUBS 0.008148f
C65 B.n37 VSUBS 0.008148f
C66 B.n38 VSUBS 0.008148f
C67 B.n39 VSUBS 0.008148f
C68 B.n40 VSUBS 0.008148f
C69 B.n41 VSUBS 0.008148f
C70 B.n42 VSUBS 0.008148f
C71 B.n43 VSUBS 0.008148f
C72 B.n44 VSUBS 0.02f
C73 B.n45 VSUBS 0.008148f
C74 B.n46 VSUBS 0.008148f
C75 B.n47 VSUBS 0.008148f
C76 B.n48 VSUBS 0.008148f
C77 B.n49 VSUBS 0.008148f
C78 B.n50 VSUBS 0.008148f
C79 B.n51 VSUBS 0.008148f
C80 B.n52 VSUBS 0.008148f
C81 B.n53 VSUBS 0.008148f
C82 B.n54 VSUBS 0.008148f
C83 B.n55 VSUBS 0.008148f
C84 B.n56 VSUBS 0.008148f
C85 B.n57 VSUBS 0.008148f
C86 B.n58 VSUBS 0.008148f
C87 B.n59 VSUBS 0.008148f
C88 B.n60 VSUBS 0.008148f
C89 B.n61 VSUBS 0.008148f
C90 B.n62 VSUBS 0.008148f
C91 B.n63 VSUBS 0.008148f
C92 B.n64 VSUBS 0.008148f
C93 B.n65 VSUBS 0.008148f
C94 B.n66 VSUBS 0.008148f
C95 B.n67 VSUBS 0.008148f
C96 B.t4 VSUBS 0.551386f
C97 B.t5 VSUBS 0.586116f
C98 B.t3 VSUBS 3.08333f
C99 B.n68 VSUBS 0.350186f
C100 B.n69 VSUBS 0.090539f
C101 B.n70 VSUBS 0.018879f
C102 B.n71 VSUBS 0.008148f
C103 B.n72 VSUBS 0.008148f
C104 B.n73 VSUBS 0.008148f
C105 B.n74 VSUBS 0.008148f
C106 B.n75 VSUBS 0.008148f
C107 B.t7 VSUBS 0.551371f
C108 B.t8 VSUBS 0.586104f
C109 B.t6 VSUBS 3.08333f
C110 B.n76 VSUBS 0.350197f
C111 B.n77 VSUBS 0.090554f
C112 B.n78 VSUBS 0.008148f
C113 B.n79 VSUBS 0.008148f
C114 B.n80 VSUBS 0.008148f
C115 B.n81 VSUBS 0.008148f
C116 B.n82 VSUBS 0.008148f
C117 B.n83 VSUBS 0.008148f
C118 B.n84 VSUBS 0.008148f
C119 B.n85 VSUBS 0.008148f
C120 B.n86 VSUBS 0.008148f
C121 B.n87 VSUBS 0.008148f
C122 B.n88 VSUBS 0.008148f
C123 B.n89 VSUBS 0.008148f
C124 B.n90 VSUBS 0.008148f
C125 B.n91 VSUBS 0.008148f
C126 B.n92 VSUBS 0.008148f
C127 B.n93 VSUBS 0.008148f
C128 B.n94 VSUBS 0.008148f
C129 B.n95 VSUBS 0.008148f
C130 B.n96 VSUBS 0.008148f
C131 B.n97 VSUBS 0.008148f
C132 B.n98 VSUBS 0.008148f
C133 B.n99 VSUBS 0.008148f
C134 B.n100 VSUBS 0.008148f
C135 B.n101 VSUBS 0.02f
C136 B.n102 VSUBS 0.008148f
C137 B.n103 VSUBS 0.008148f
C138 B.n104 VSUBS 0.008148f
C139 B.n105 VSUBS 0.008148f
C140 B.n106 VSUBS 0.008148f
C141 B.n107 VSUBS 0.008148f
C142 B.n108 VSUBS 0.008148f
C143 B.n109 VSUBS 0.008148f
C144 B.n110 VSUBS 0.008148f
C145 B.n111 VSUBS 0.008148f
C146 B.n112 VSUBS 0.008148f
C147 B.n113 VSUBS 0.008148f
C148 B.n114 VSUBS 0.008148f
C149 B.n115 VSUBS 0.008148f
C150 B.n116 VSUBS 0.008148f
C151 B.n117 VSUBS 0.008148f
C152 B.n118 VSUBS 0.008148f
C153 B.n119 VSUBS 0.008148f
C154 B.n120 VSUBS 0.008148f
C155 B.n121 VSUBS 0.008148f
C156 B.n122 VSUBS 0.008148f
C157 B.n123 VSUBS 0.008148f
C158 B.n124 VSUBS 0.008148f
C159 B.n125 VSUBS 0.008148f
C160 B.n126 VSUBS 0.008148f
C161 B.n127 VSUBS 0.008148f
C162 B.n128 VSUBS 0.008148f
C163 B.n129 VSUBS 0.008148f
C164 B.n130 VSUBS 0.008148f
C165 B.n131 VSUBS 0.008148f
C166 B.n132 VSUBS 0.008148f
C167 B.n133 VSUBS 0.008148f
C168 B.n134 VSUBS 0.008148f
C169 B.n135 VSUBS 0.008148f
C170 B.n136 VSUBS 0.008148f
C171 B.n137 VSUBS 0.008148f
C172 B.n138 VSUBS 0.008148f
C173 B.n139 VSUBS 0.008148f
C174 B.n140 VSUBS 0.008148f
C175 B.n141 VSUBS 0.008148f
C176 B.n142 VSUBS 0.008148f
C177 B.n143 VSUBS 0.008148f
C178 B.n144 VSUBS 0.008148f
C179 B.n145 VSUBS 0.008148f
C180 B.n146 VSUBS 0.008148f
C181 B.n147 VSUBS 0.008148f
C182 B.n148 VSUBS 0.008148f
C183 B.n149 VSUBS 0.008148f
C184 B.n150 VSUBS 0.008148f
C185 B.n151 VSUBS 0.008148f
C186 B.n152 VSUBS 0.008148f
C187 B.n153 VSUBS 0.008148f
C188 B.n154 VSUBS 0.008148f
C189 B.n155 VSUBS 0.008148f
C190 B.n156 VSUBS 0.008148f
C191 B.n157 VSUBS 0.008148f
C192 B.n158 VSUBS 0.008148f
C193 B.n159 VSUBS 0.008148f
C194 B.n160 VSUBS 0.008148f
C195 B.n161 VSUBS 0.008148f
C196 B.n162 VSUBS 0.008148f
C197 B.n163 VSUBS 0.008148f
C198 B.n164 VSUBS 0.008148f
C199 B.n165 VSUBS 0.008148f
C200 B.n166 VSUBS 0.008148f
C201 B.n167 VSUBS 0.008148f
C202 B.n168 VSUBS 0.008148f
C203 B.n169 VSUBS 0.008148f
C204 B.n170 VSUBS 0.008148f
C205 B.n171 VSUBS 0.008148f
C206 B.n172 VSUBS 0.008148f
C207 B.n173 VSUBS 0.008148f
C208 B.n174 VSUBS 0.008148f
C209 B.n175 VSUBS 0.008148f
C210 B.n176 VSUBS 0.008148f
C211 B.n177 VSUBS 0.008148f
C212 B.n178 VSUBS 0.008148f
C213 B.n179 VSUBS 0.008148f
C214 B.n180 VSUBS 0.008148f
C215 B.n181 VSUBS 0.008148f
C216 B.n182 VSUBS 0.008148f
C217 B.n183 VSUBS 0.008148f
C218 B.n184 VSUBS 0.008148f
C219 B.n185 VSUBS 0.008148f
C220 B.n186 VSUBS 0.020224f
C221 B.n187 VSUBS 0.008148f
C222 B.n188 VSUBS 0.008148f
C223 B.n189 VSUBS 0.008148f
C224 B.n190 VSUBS 0.008148f
C225 B.n191 VSUBS 0.008148f
C226 B.n192 VSUBS 0.008148f
C227 B.n193 VSUBS 0.008148f
C228 B.n194 VSUBS 0.008148f
C229 B.n195 VSUBS 0.008148f
C230 B.n196 VSUBS 0.008148f
C231 B.n197 VSUBS 0.008148f
C232 B.n198 VSUBS 0.008148f
C233 B.n199 VSUBS 0.008148f
C234 B.n200 VSUBS 0.008148f
C235 B.n201 VSUBS 0.008148f
C236 B.n202 VSUBS 0.008148f
C237 B.n203 VSUBS 0.008148f
C238 B.n204 VSUBS 0.008148f
C239 B.n205 VSUBS 0.008148f
C240 B.n206 VSUBS 0.008148f
C241 B.n207 VSUBS 0.008148f
C242 B.n208 VSUBS 0.008148f
C243 B.n209 VSUBS 0.008148f
C244 B.n210 VSUBS 0.007669f
C245 B.n211 VSUBS 0.008148f
C246 B.n212 VSUBS 0.008148f
C247 B.n213 VSUBS 0.008148f
C248 B.n214 VSUBS 0.008148f
C249 B.n215 VSUBS 0.008148f
C250 B.t2 VSUBS 0.551386f
C251 B.t1 VSUBS 0.586116f
C252 B.t0 VSUBS 3.08333f
C253 B.n216 VSUBS 0.350186f
C254 B.n217 VSUBS 0.090539f
C255 B.n218 VSUBS 0.008148f
C256 B.n219 VSUBS 0.008148f
C257 B.n220 VSUBS 0.008148f
C258 B.n221 VSUBS 0.008148f
C259 B.n222 VSUBS 0.008148f
C260 B.n223 VSUBS 0.008148f
C261 B.n224 VSUBS 0.008148f
C262 B.n225 VSUBS 0.008148f
C263 B.n226 VSUBS 0.008148f
C264 B.n227 VSUBS 0.008148f
C265 B.n228 VSUBS 0.008148f
C266 B.n229 VSUBS 0.008148f
C267 B.n230 VSUBS 0.008148f
C268 B.n231 VSUBS 0.008148f
C269 B.n232 VSUBS 0.008148f
C270 B.n233 VSUBS 0.008148f
C271 B.n234 VSUBS 0.008148f
C272 B.n235 VSUBS 0.008148f
C273 B.n236 VSUBS 0.008148f
C274 B.n237 VSUBS 0.008148f
C275 B.n238 VSUBS 0.008148f
C276 B.n239 VSUBS 0.008148f
C277 B.n240 VSUBS 0.008148f
C278 B.n241 VSUBS 0.02f
C279 B.n242 VSUBS 0.008148f
C280 B.n243 VSUBS 0.008148f
C281 B.n244 VSUBS 0.008148f
C282 B.n245 VSUBS 0.008148f
C283 B.n246 VSUBS 0.008148f
C284 B.n247 VSUBS 0.008148f
C285 B.n248 VSUBS 0.008148f
C286 B.n249 VSUBS 0.008148f
C287 B.n250 VSUBS 0.008148f
C288 B.n251 VSUBS 0.008148f
C289 B.n252 VSUBS 0.008148f
C290 B.n253 VSUBS 0.008148f
C291 B.n254 VSUBS 0.008148f
C292 B.n255 VSUBS 0.008148f
C293 B.n256 VSUBS 0.008148f
C294 B.n257 VSUBS 0.008148f
C295 B.n258 VSUBS 0.008148f
C296 B.n259 VSUBS 0.008148f
C297 B.n260 VSUBS 0.008148f
C298 B.n261 VSUBS 0.008148f
C299 B.n262 VSUBS 0.008148f
C300 B.n263 VSUBS 0.008148f
C301 B.n264 VSUBS 0.008148f
C302 B.n265 VSUBS 0.008148f
C303 B.n266 VSUBS 0.008148f
C304 B.n267 VSUBS 0.008148f
C305 B.n268 VSUBS 0.008148f
C306 B.n269 VSUBS 0.008148f
C307 B.n270 VSUBS 0.008148f
C308 B.n271 VSUBS 0.008148f
C309 B.n272 VSUBS 0.008148f
C310 B.n273 VSUBS 0.008148f
C311 B.n274 VSUBS 0.008148f
C312 B.n275 VSUBS 0.008148f
C313 B.n276 VSUBS 0.008148f
C314 B.n277 VSUBS 0.008148f
C315 B.n278 VSUBS 0.008148f
C316 B.n279 VSUBS 0.008148f
C317 B.n280 VSUBS 0.008148f
C318 B.n281 VSUBS 0.008148f
C319 B.n282 VSUBS 0.008148f
C320 B.n283 VSUBS 0.008148f
C321 B.n284 VSUBS 0.008148f
C322 B.n285 VSUBS 0.008148f
C323 B.n286 VSUBS 0.008148f
C324 B.n287 VSUBS 0.008148f
C325 B.n288 VSUBS 0.008148f
C326 B.n289 VSUBS 0.008148f
C327 B.n290 VSUBS 0.008148f
C328 B.n291 VSUBS 0.008148f
C329 B.n292 VSUBS 0.008148f
C330 B.n293 VSUBS 0.008148f
C331 B.n294 VSUBS 0.008148f
C332 B.n295 VSUBS 0.008148f
C333 B.n296 VSUBS 0.008148f
C334 B.n297 VSUBS 0.008148f
C335 B.n298 VSUBS 0.008148f
C336 B.n299 VSUBS 0.008148f
C337 B.n300 VSUBS 0.008148f
C338 B.n301 VSUBS 0.008148f
C339 B.n302 VSUBS 0.008148f
C340 B.n303 VSUBS 0.008148f
C341 B.n304 VSUBS 0.008148f
C342 B.n305 VSUBS 0.008148f
C343 B.n306 VSUBS 0.008148f
C344 B.n307 VSUBS 0.008148f
C345 B.n308 VSUBS 0.008148f
C346 B.n309 VSUBS 0.008148f
C347 B.n310 VSUBS 0.008148f
C348 B.n311 VSUBS 0.008148f
C349 B.n312 VSUBS 0.008148f
C350 B.n313 VSUBS 0.008148f
C351 B.n314 VSUBS 0.008148f
C352 B.n315 VSUBS 0.008148f
C353 B.n316 VSUBS 0.008148f
C354 B.n317 VSUBS 0.008148f
C355 B.n318 VSUBS 0.008148f
C356 B.n319 VSUBS 0.008148f
C357 B.n320 VSUBS 0.008148f
C358 B.n321 VSUBS 0.008148f
C359 B.n322 VSUBS 0.008148f
C360 B.n323 VSUBS 0.008148f
C361 B.n324 VSUBS 0.008148f
C362 B.n325 VSUBS 0.008148f
C363 B.n326 VSUBS 0.008148f
C364 B.n327 VSUBS 0.008148f
C365 B.n328 VSUBS 0.008148f
C366 B.n329 VSUBS 0.008148f
C367 B.n330 VSUBS 0.008148f
C368 B.n331 VSUBS 0.008148f
C369 B.n332 VSUBS 0.008148f
C370 B.n333 VSUBS 0.008148f
C371 B.n334 VSUBS 0.008148f
C372 B.n335 VSUBS 0.008148f
C373 B.n336 VSUBS 0.008148f
C374 B.n337 VSUBS 0.008148f
C375 B.n338 VSUBS 0.008148f
C376 B.n339 VSUBS 0.008148f
C377 B.n340 VSUBS 0.008148f
C378 B.n341 VSUBS 0.008148f
C379 B.n342 VSUBS 0.008148f
C380 B.n343 VSUBS 0.008148f
C381 B.n344 VSUBS 0.008148f
C382 B.n345 VSUBS 0.008148f
C383 B.n346 VSUBS 0.008148f
C384 B.n347 VSUBS 0.008148f
C385 B.n348 VSUBS 0.008148f
C386 B.n349 VSUBS 0.008148f
C387 B.n350 VSUBS 0.008148f
C388 B.n351 VSUBS 0.008148f
C389 B.n352 VSUBS 0.008148f
C390 B.n353 VSUBS 0.008148f
C391 B.n354 VSUBS 0.008148f
C392 B.n355 VSUBS 0.008148f
C393 B.n356 VSUBS 0.008148f
C394 B.n357 VSUBS 0.008148f
C395 B.n358 VSUBS 0.008148f
C396 B.n359 VSUBS 0.008148f
C397 B.n360 VSUBS 0.008148f
C398 B.n361 VSUBS 0.008148f
C399 B.n362 VSUBS 0.008148f
C400 B.n363 VSUBS 0.008148f
C401 B.n364 VSUBS 0.008148f
C402 B.n365 VSUBS 0.008148f
C403 B.n366 VSUBS 0.008148f
C404 B.n367 VSUBS 0.008148f
C405 B.n368 VSUBS 0.008148f
C406 B.n369 VSUBS 0.008148f
C407 B.n370 VSUBS 0.008148f
C408 B.n371 VSUBS 0.008148f
C409 B.n372 VSUBS 0.008148f
C410 B.n373 VSUBS 0.008148f
C411 B.n374 VSUBS 0.008148f
C412 B.n375 VSUBS 0.008148f
C413 B.n376 VSUBS 0.008148f
C414 B.n377 VSUBS 0.008148f
C415 B.n378 VSUBS 0.008148f
C416 B.n379 VSUBS 0.008148f
C417 B.n380 VSUBS 0.008148f
C418 B.n381 VSUBS 0.008148f
C419 B.n382 VSUBS 0.008148f
C420 B.n383 VSUBS 0.008148f
C421 B.n384 VSUBS 0.008148f
C422 B.n385 VSUBS 0.008148f
C423 B.n386 VSUBS 0.008148f
C424 B.n387 VSUBS 0.008148f
C425 B.n388 VSUBS 0.008148f
C426 B.n389 VSUBS 0.008148f
C427 B.n390 VSUBS 0.008148f
C428 B.n391 VSUBS 0.008148f
C429 B.n392 VSUBS 0.008148f
C430 B.n393 VSUBS 0.008148f
C431 B.n394 VSUBS 0.008148f
C432 B.n395 VSUBS 0.008148f
C433 B.n396 VSUBS 0.008148f
C434 B.n397 VSUBS 0.008148f
C435 B.n398 VSUBS 0.008148f
C436 B.n399 VSUBS 0.008148f
C437 B.n400 VSUBS 0.008148f
C438 B.n401 VSUBS 0.008148f
C439 B.n402 VSUBS 0.008148f
C440 B.n403 VSUBS 0.008148f
C441 B.n404 VSUBS 0.008148f
C442 B.n405 VSUBS 0.008148f
C443 B.n406 VSUBS 0.019304f
C444 B.n407 VSUBS 0.019304f
C445 B.n408 VSUBS 0.02f
C446 B.n409 VSUBS 0.008148f
C447 B.n410 VSUBS 0.008148f
C448 B.n411 VSUBS 0.008148f
C449 B.n412 VSUBS 0.008148f
C450 B.n413 VSUBS 0.008148f
C451 B.n414 VSUBS 0.008148f
C452 B.n415 VSUBS 0.008148f
C453 B.n416 VSUBS 0.008148f
C454 B.n417 VSUBS 0.008148f
C455 B.n418 VSUBS 0.008148f
C456 B.n419 VSUBS 0.008148f
C457 B.n420 VSUBS 0.008148f
C458 B.n421 VSUBS 0.008148f
C459 B.n422 VSUBS 0.008148f
C460 B.n423 VSUBS 0.008148f
C461 B.n424 VSUBS 0.008148f
C462 B.n425 VSUBS 0.008148f
C463 B.n426 VSUBS 0.008148f
C464 B.n427 VSUBS 0.008148f
C465 B.n428 VSUBS 0.008148f
C466 B.n429 VSUBS 0.008148f
C467 B.n430 VSUBS 0.008148f
C468 B.n431 VSUBS 0.008148f
C469 B.n432 VSUBS 0.008148f
C470 B.n433 VSUBS 0.008148f
C471 B.n434 VSUBS 0.008148f
C472 B.n435 VSUBS 0.008148f
C473 B.n436 VSUBS 0.008148f
C474 B.n437 VSUBS 0.008148f
C475 B.n438 VSUBS 0.008148f
C476 B.n439 VSUBS 0.008148f
C477 B.n440 VSUBS 0.008148f
C478 B.n441 VSUBS 0.008148f
C479 B.n442 VSUBS 0.008148f
C480 B.n443 VSUBS 0.008148f
C481 B.n444 VSUBS 0.008148f
C482 B.n445 VSUBS 0.008148f
C483 B.n446 VSUBS 0.008148f
C484 B.n447 VSUBS 0.008148f
C485 B.n448 VSUBS 0.008148f
C486 B.n449 VSUBS 0.008148f
C487 B.n450 VSUBS 0.008148f
C488 B.n451 VSUBS 0.008148f
C489 B.n452 VSUBS 0.008148f
C490 B.n453 VSUBS 0.008148f
C491 B.n454 VSUBS 0.008148f
C492 B.n455 VSUBS 0.008148f
C493 B.n456 VSUBS 0.008148f
C494 B.n457 VSUBS 0.008148f
C495 B.n458 VSUBS 0.008148f
C496 B.n459 VSUBS 0.008148f
C497 B.n460 VSUBS 0.008148f
C498 B.n461 VSUBS 0.008148f
C499 B.n462 VSUBS 0.008148f
C500 B.n463 VSUBS 0.008148f
C501 B.n464 VSUBS 0.008148f
C502 B.n465 VSUBS 0.008148f
C503 B.n466 VSUBS 0.008148f
C504 B.n467 VSUBS 0.008148f
C505 B.n468 VSUBS 0.008148f
C506 B.n469 VSUBS 0.008148f
C507 B.n470 VSUBS 0.008148f
C508 B.n471 VSUBS 0.008148f
C509 B.n472 VSUBS 0.008148f
C510 B.n473 VSUBS 0.008148f
C511 B.n474 VSUBS 0.008148f
C512 B.n475 VSUBS 0.008148f
C513 B.n476 VSUBS 0.008148f
C514 B.n477 VSUBS 0.008148f
C515 B.n478 VSUBS 0.008148f
C516 B.n479 VSUBS 0.007669f
C517 B.n480 VSUBS 0.018879f
C518 B.n481 VSUBS 0.004554f
C519 B.n482 VSUBS 0.008148f
C520 B.n483 VSUBS 0.008148f
C521 B.n484 VSUBS 0.008148f
C522 B.n485 VSUBS 0.008148f
C523 B.n486 VSUBS 0.008148f
C524 B.n487 VSUBS 0.008148f
C525 B.n488 VSUBS 0.008148f
C526 B.n489 VSUBS 0.008148f
C527 B.n490 VSUBS 0.008148f
C528 B.n491 VSUBS 0.008148f
C529 B.n492 VSUBS 0.008148f
C530 B.n493 VSUBS 0.008148f
C531 B.t11 VSUBS 0.551371f
C532 B.t10 VSUBS 0.586104f
C533 B.t9 VSUBS 3.08333f
C534 B.n494 VSUBS 0.350197f
C535 B.n495 VSUBS 0.090554f
C536 B.n496 VSUBS 0.018879f
C537 B.n497 VSUBS 0.004554f
C538 B.n498 VSUBS 0.008148f
C539 B.n499 VSUBS 0.008148f
C540 B.n500 VSUBS 0.008148f
C541 B.n501 VSUBS 0.008148f
C542 B.n502 VSUBS 0.008148f
C543 B.n503 VSUBS 0.008148f
C544 B.n504 VSUBS 0.008148f
C545 B.n505 VSUBS 0.008148f
C546 B.n506 VSUBS 0.008148f
C547 B.n507 VSUBS 0.008148f
C548 B.n508 VSUBS 0.008148f
C549 B.n509 VSUBS 0.008148f
C550 B.n510 VSUBS 0.008148f
C551 B.n511 VSUBS 0.008148f
C552 B.n512 VSUBS 0.008148f
C553 B.n513 VSUBS 0.008148f
C554 B.n514 VSUBS 0.008148f
C555 B.n515 VSUBS 0.008148f
C556 B.n516 VSUBS 0.008148f
C557 B.n517 VSUBS 0.008148f
C558 B.n518 VSUBS 0.008148f
C559 B.n519 VSUBS 0.008148f
C560 B.n520 VSUBS 0.008148f
C561 B.n521 VSUBS 0.008148f
C562 B.n522 VSUBS 0.008148f
C563 B.n523 VSUBS 0.008148f
C564 B.n524 VSUBS 0.008148f
C565 B.n525 VSUBS 0.008148f
C566 B.n526 VSUBS 0.008148f
C567 B.n527 VSUBS 0.008148f
C568 B.n528 VSUBS 0.008148f
C569 B.n529 VSUBS 0.008148f
C570 B.n530 VSUBS 0.008148f
C571 B.n531 VSUBS 0.008148f
C572 B.n532 VSUBS 0.008148f
C573 B.n533 VSUBS 0.008148f
C574 B.n534 VSUBS 0.008148f
C575 B.n535 VSUBS 0.008148f
C576 B.n536 VSUBS 0.008148f
C577 B.n537 VSUBS 0.008148f
C578 B.n538 VSUBS 0.008148f
C579 B.n539 VSUBS 0.008148f
C580 B.n540 VSUBS 0.008148f
C581 B.n541 VSUBS 0.008148f
C582 B.n542 VSUBS 0.008148f
C583 B.n543 VSUBS 0.008148f
C584 B.n544 VSUBS 0.008148f
C585 B.n545 VSUBS 0.008148f
C586 B.n546 VSUBS 0.008148f
C587 B.n547 VSUBS 0.008148f
C588 B.n548 VSUBS 0.008148f
C589 B.n549 VSUBS 0.008148f
C590 B.n550 VSUBS 0.008148f
C591 B.n551 VSUBS 0.008148f
C592 B.n552 VSUBS 0.008148f
C593 B.n553 VSUBS 0.008148f
C594 B.n554 VSUBS 0.008148f
C595 B.n555 VSUBS 0.008148f
C596 B.n556 VSUBS 0.008148f
C597 B.n557 VSUBS 0.008148f
C598 B.n558 VSUBS 0.008148f
C599 B.n559 VSUBS 0.008148f
C600 B.n560 VSUBS 0.008148f
C601 B.n561 VSUBS 0.008148f
C602 B.n562 VSUBS 0.008148f
C603 B.n563 VSUBS 0.008148f
C604 B.n564 VSUBS 0.008148f
C605 B.n565 VSUBS 0.008148f
C606 B.n566 VSUBS 0.008148f
C607 B.n567 VSUBS 0.008148f
C608 B.n568 VSUBS 0.008148f
C609 B.n569 VSUBS 0.01908f
C610 B.n570 VSUBS 0.02f
C611 B.n571 VSUBS 0.019304f
C612 B.n572 VSUBS 0.008148f
C613 B.n573 VSUBS 0.008148f
C614 B.n574 VSUBS 0.008148f
C615 B.n575 VSUBS 0.008148f
C616 B.n576 VSUBS 0.008148f
C617 B.n577 VSUBS 0.008148f
C618 B.n578 VSUBS 0.008148f
C619 B.n579 VSUBS 0.008148f
C620 B.n580 VSUBS 0.008148f
C621 B.n581 VSUBS 0.008148f
C622 B.n582 VSUBS 0.008148f
C623 B.n583 VSUBS 0.008148f
C624 B.n584 VSUBS 0.008148f
C625 B.n585 VSUBS 0.008148f
C626 B.n586 VSUBS 0.008148f
C627 B.n587 VSUBS 0.008148f
C628 B.n588 VSUBS 0.008148f
C629 B.n589 VSUBS 0.008148f
C630 B.n590 VSUBS 0.008148f
C631 B.n591 VSUBS 0.008148f
C632 B.n592 VSUBS 0.008148f
C633 B.n593 VSUBS 0.008148f
C634 B.n594 VSUBS 0.008148f
C635 B.n595 VSUBS 0.008148f
C636 B.n596 VSUBS 0.008148f
C637 B.n597 VSUBS 0.008148f
C638 B.n598 VSUBS 0.008148f
C639 B.n599 VSUBS 0.008148f
C640 B.n600 VSUBS 0.008148f
C641 B.n601 VSUBS 0.008148f
C642 B.n602 VSUBS 0.008148f
C643 B.n603 VSUBS 0.008148f
C644 B.n604 VSUBS 0.008148f
C645 B.n605 VSUBS 0.008148f
C646 B.n606 VSUBS 0.008148f
C647 B.n607 VSUBS 0.008148f
C648 B.n608 VSUBS 0.008148f
C649 B.n609 VSUBS 0.008148f
C650 B.n610 VSUBS 0.008148f
C651 B.n611 VSUBS 0.008148f
C652 B.n612 VSUBS 0.008148f
C653 B.n613 VSUBS 0.008148f
C654 B.n614 VSUBS 0.008148f
C655 B.n615 VSUBS 0.008148f
C656 B.n616 VSUBS 0.008148f
C657 B.n617 VSUBS 0.008148f
C658 B.n618 VSUBS 0.008148f
C659 B.n619 VSUBS 0.008148f
C660 B.n620 VSUBS 0.008148f
C661 B.n621 VSUBS 0.008148f
C662 B.n622 VSUBS 0.008148f
C663 B.n623 VSUBS 0.008148f
C664 B.n624 VSUBS 0.008148f
C665 B.n625 VSUBS 0.008148f
C666 B.n626 VSUBS 0.008148f
C667 B.n627 VSUBS 0.008148f
C668 B.n628 VSUBS 0.008148f
C669 B.n629 VSUBS 0.008148f
C670 B.n630 VSUBS 0.008148f
C671 B.n631 VSUBS 0.008148f
C672 B.n632 VSUBS 0.008148f
C673 B.n633 VSUBS 0.008148f
C674 B.n634 VSUBS 0.008148f
C675 B.n635 VSUBS 0.008148f
C676 B.n636 VSUBS 0.008148f
C677 B.n637 VSUBS 0.008148f
C678 B.n638 VSUBS 0.008148f
C679 B.n639 VSUBS 0.008148f
C680 B.n640 VSUBS 0.008148f
C681 B.n641 VSUBS 0.008148f
C682 B.n642 VSUBS 0.008148f
C683 B.n643 VSUBS 0.008148f
C684 B.n644 VSUBS 0.008148f
C685 B.n645 VSUBS 0.008148f
C686 B.n646 VSUBS 0.008148f
C687 B.n647 VSUBS 0.008148f
C688 B.n648 VSUBS 0.008148f
C689 B.n649 VSUBS 0.008148f
C690 B.n650 VSUBS 0.008148f
C691 B.n651 VSUBS 0.008148f
C692 B.n652 VSUBS 0.008148f
C693 B.n653 VSUBS 0.008148f
C694 B.n654 VSUBS 0.008148f
C695 B.n655 VSUBS 0.008148f
C696 B.n656 VSUBS 0.008148f
C697 B.n657 VSUBS 0.008148f
C698 B.n658 VSUBS 0.008148f
C699 B.n659 VSUBS 0.008148f
C700 B.n660 VSUBS 0.008148f
C701 B.n661 VSUBS 0.008148f
C702 B.n662 VSUBS 0.008148f
C703 B.n663 VSUBS 0.008148f
C704 B.n664 VSUBS 0.008148f
C705 B.n665 VSUBS 0.008148f
C706 B.n666 VSUBS 0.008148f
C707 B.n667 VSUBS 0.008148f
C708 B.n668 VSUBS 0.008148f
C709 B.n669 VSUBS 0.008148f
C710 B.n670 VSUBS 0.008148f
C711 B.n671 VSUBS 0.008148f
C712 B.n672 VSUBS 0.008148f
C713 B.n673 VSUBS 0.008148f
C714 B.n674 VSUBS 0.008148f
C715 B.n675 VSUBS 0.008148f
C716 B.n676 VSUBS 0.008148f
C717 B.n677 VSUBS 0.008148f
C718 B.n678 VSUBS 0.008148f
C719 B.n679 VSUBS 0.008148f
C720 B.n680 VSUBS 0.008148f
C721 B.n681 VSUBS 0.008148f
C722 B.n682 VSUBS 0.008148f
C723 B.n683 VSUBS 0.008148f
C724 B.n684 VSUBS 0.008148f
C725 B.n685 VSUBS 0.008148f
C726 B.n686 VSUBS 0.008148f
C727 B.n687 VSUBS 0.008148f
C728 B.n688 VSUBS 0.008148f
C729 B.n689 VSUBS 0.008148f
C730 B.n690 VSUBS 0.008148f
C731 B.n691 VSUBS 0.008148f
C732 B.n692 VSUBS 0.008148f
C733 B.n693 VSUBS 0.008148f
C734 B.n694 VSUBS 0.008148f
C735 B.n695 VSUBS 0.008148f
C736 B.n696 VSUBS 0.008148f
C737 B.n697 VSUBS 0.008148f
C738 B.n698 VSUBS 0.008148f
C739 B.n699 VSUBS 0.008148f
C740 B.n700 VSUBS 0.008148f
C741 B.n701 VSUBS 0.008148f
C742 B.n702 VSUBS 0.008148f
C743 B.n703 VSUBS 0.008148f
C744 B.n704 VSUBS 0.008148f
C745 B.n705 VSUBS 0.008148f
C746 B.n706 VSUBS 0.008148f
C747 B.n707 VSUBS 0.008148f
C748 B.n708 VSUBS 0.008148f
C749 B.n709 VSUBS 0.008148f
C750 B.n710 VSUBS 0.008148f
C751 B.n711 VSUBS 0.008148f
C752 B.n712 VSUBS 0.008148f
C753 B.n713 VSUBS 0.008148f
C754 B.n714 VSUBS 0.008148f
C755 B.n715 VSUBS 0.008148f
C756 B.n716 VSUBS 0.008148f
C757 B.n717 VSUBS 0.008148f
C758 B.n718 VSUBS 0.008148f
C759 B.n719 VSUBS 0.008148f
C760 B.n720 VSUBS 0.008148f
C761 B.n721 VSUBS 0.008148f
C762 B.n722 VSUBS 0.008148f
C763 B.n723 VSUBS 0.008148f
C764 B.n724 VSUBS 0.008148f
C765 B.n725 VSUBS 0.008148f
C766 B.n726 VSUBS 0.008148f
C767 B.n727 VSUBS 0.008148f
C768 B.n728 VSUBS 0.008148f
C769 B.n729 VSUBS 0.008148f
C770 B.n730 VSUBS 0.008148f
C771 B.n731 VSUBS 0.008148f
C772 B.n732 VSUBS 0.008148f
C773 B.n733 VSUBS 0.008148f
C774 B.n734 VSUBS 0.008148f
C775 B.n735 VSUBS 0.008148f
C776 B.n736 VSUBS 0.008148f
C777 B.n737 VSUBS 0.008148f
C778 B.n738 VSUBS 0.008148f
C779 B.n739 VSUBS 0.008148f
C780 B.n740 VSUBS 0.008148f
C781 B.n741 VSUBS 0.008148f
C782 B.n742 VSUBS 0.008148f
C783 B.n743 VSUBS 0.008148f
C784 B.n744 VSUBS 0.008148f
C785 B.n745 VSUBS 0.008148f
C786 B.n746 VSUBS 0.008148f
C787 B.n747 VSUBS 0.008148f
C788 B.n748 VSUBS 0.008148f
C789 B.n749 VSUBS 0.008148f
C790 B.n750 VSUBS 0.008148f
C791 B.n751 VSUBS 0.008148f
C792 B.n752 VSUBS 0.008148f
C793 B.n753 VSUBS 0.008148f
C794 B.n754 VSUBS 0.008148f
C795 B.n755 VSUBS 0.008148f
C796 B.n756 VSUBS 0.008148f
C797 B.n757 VSUBS 0.008148f
C798 B.n758 VSUBS 0.008148f
C799 B.n759 VSUBS 0.008148f
C800 B.n760 VSUBS 0.008148f
C801 B.n761 VSUBS 0.008148f
C802 B.n762 VSUBS 0.008148f
C803 B.n763 VSUBS 0.008148f
C804 B.n764 VSUBS 0.008148f
C805 B.n765 VSUBS 0.008148f
C806 B.n766 VSUBS 0.008148f
C807 B.n767 VSUBS 0.008148f
C808 B.n768 VSUBS 0.008148f
C809 B.n769 VSUBS 0.008148f
C810 B.n770 VSUBS 0.008148f
C811 B.n771 VSUBS 0.008148f
C812 B.n772 VSUBS 0.008148f
C813 B.n773 VSUBS 0.008148f
C814 B.n774 VSUBS 0.008148f
C815 B.n775 VSUBS 0.008148f
C816 B.n776 VSUBS 0.008148f
C817 B.n777 VSUBS 0.008148f
C818 B.n778 VSUBS 0.008148f
C819 B.n779 VSUBS 0.008148f
C820 B.n780 VSUBS 0.008148f
C821 B.n781 VSUBS 0.008148f
C822 B.n782 VSUBS 0.008148f
C823 B.n783 VSUBS 0.008148f
C824 B.n784 VSUBS 0.008148f
C825 B.n785 VSUBS 0.008148f
C826 B.n786 VSUBS 0.008148f
C827 B.n787 VSUBS 0.008148f
C828 B.n788 VSUBS 0.008148f
C829 B.n789 VSUBS 0.008148f
C830 B.n790 VSUBS 0.008148f
C831 B.n791 VSUBS 0.008148f
C832 B.n792 VSUBS 0.008148f
C833 B.n793 VSUBS 0.008148f
C834 B.n794 VSUBS 0.008148f
C835 B.n795 VSUBS 0.008148f
C836 B.n796 VSUBS 0.008148f
C837 B.n797 VSUBS 0.008148f
C838 B.n798 VSUBS 0.008148f
C839 B.n799 VSUBS 0.008148f
C840 B.n800 VSUBS 0.008148f
C841 B.n801 VSUBS 0.008148f
C842 B.n802 VSUBS 0.008148f
C843 B.n803 VSUBS 0.008148f
C844 B.n804 VSUBS 0.008148f
C845 B.n805 VSUBS 0.008148f
C846 B.n806 VSUBS 0.008148f
C847 B.n807 VSUBS 0.008148f
C848 B.n808 VSUBS 0.008148f
C849 B.n809 VSUBS 0.008148f
C850 B.n810 VSUBS 0.008148f
C851 B.n811 VSUBS 0.008148f
C852 B.n812 VSUBS 0.008148f
C853 B.n813 VSUBS 0.008148f
C854 B.n814 VSUBS 0.008148f
C855 B.n815 VSUBS 0.008148f
C856 B.n816 VSUBS 0.008148f
C857 B.n817 VSUBS 0.008148f
C858 B.n818 VSUBS 0.008148f
C859 B.n819 VSUBS 0.008148f
C860 B.n820 VSUBS 0.008148f
C861 B.n821 VSUBS 0.008148f
C862 B.n822 VSUBS 0.008148f
C863 B.n823 VSUBS 0.008148f
C864 B.n824 VSUBS 0.019304f
C865 B.n825 VSUBS 0.019304f
C866 B.n826 VSUBS 0.02f
C867 B.n827 VSUBS 0.008148f
C868 B.n828 VSUBS 0.008148f
C869 B.n829 VSUBS 0.008148f
C870 B.n830 VSUBS 0.008148f
C871 B.n831 VSUBS 0.008148f
C872 B.n832 VSUBS 0.008148f
C873 B.n833 VSUBS 0.008148f
C874 B.n834 VSUBS 0.008148f
C875 B.n835 VSUBS 0.008148f
C876 B.n836 VSUBS 0.008148f
C877 B.n837 VSUBS 0.008148f
C878 B.n838 VSUBS 0.008148f
C879 B.n839 VSUBS 0.008148f
C880 B.n840 VSUBS 0.008148f
C881 B.n841 VSUBS 0.008148f
C882 B.n842 VSUBS 0.008148f
C883 B.n843 VSUBS 0.008148f
C884 B.n844 VSUBS 0.008148f
C885 B.n845 VSUBS 0.008148f
C886 B.n846 VSUBS 0.008148f
C887 B.n847 VSUBS 0.008148f
C888 B.n848 VSUBS 0.008148f
C889 B.n849 VSUBS 0.008148f
C890 B.n850 VSUBS 0.008148f
C891 B.n851 VSUBS 0.008148f
C892 B.n852 VSUBS 0.008148f
C893 B.n853 VSUBS 0.008148f
C894 B.n854 VSUBS 0.008148f
C895 B.n855 VSUBS 0.008148f
C896 B.n856 VSUBS 0.008148f
C897 B.n857 VSUBS 0.008148f
C898 B.n858 VSUBS 0.008148f
C899 B.n859 VSUBS 0.008148f
C900 B.n860 VSUBS 0.008148f
C901 B.n861 VSUBS 0.008148f
C902 B.n862 VSUBS 0.008148f
C903 B.n863 VSUBS 0.008148f
C904 B.n864 VSUBS 0.008148f
C905 B.n865 VSUBS 0.008148f
C906 B.n866 VSUBS 0.008148f
C907 B.n867 VSUBS 0.008148f
C908 B.n868 VSUBS 0.008148f
C909 B.n869 VSUBS 0.008148f
C910 B.n870 VSUBS 0.008148f
C911 B.n871 VSUBS 0.008148f
C912 B.n872 VSUBS 0.008148f
C913 B.n873 VSUBS 0.008148f
C914 B.n874 VSUBS 0.008148f
C915 B.n875 VSUBS 0.008148f
C916 B.n876 VSUBS 0.008148f
C917 B.n877 VSUBS 0.008148f
C918 B.n878 VSUBS 0.008148f
C919 B.n879 VSUBS 0.008148f
C920 B.n880 VSUBS 0.008148f
C921 B.n881 VSUBS 0.008148f
C922 B.n882 VSUBS 0.008148f
C923 B.n883 VSUBS 0.008148f
C924 B.n884 VSUBS 0.008148f
C925 B.n885 VSUBS 0.008148f
C926 B.n886 VSUBS 0.008148f
C927 B.n887 VSUBS 0.008148f
C928 B.n888 VSUBS 0.008148f
C929 B.n889 VSUBS 0.008148f
C930 B.n890 VSUBS 0.008148f
C931 B.n891 VSUBS 0.008148f
C932 B.n892 VSUBS 0.008148f
C933 B.n893 VSUBS 0.008148f
C934 B.n894 VSUBS 0.008148f
C935 B.n895 VSUBS 0.008148f
C936 B.n896 VSUBS 0.008148f
C937 B.n897 VSUBS 0.007669f
C938 B.n898 VSUBS 0.018879f
C939 B.n899 VSUBS 0.004554f
C940 B.n900 VSUBS 0.008148f
C941 B.n901 VSUBS 0.008148f
C942 B.n902 VSUBS 0.008148f
C943 B.n903 VSUBS 0.008148f
C944 B.n904 VSUBS 0.008148f
C945 B.n905 VSUBS 0.008148f
C946 B.n906 VSUBS 0.008148f
C947 B.n907 VSUBS 0.008148f
C948 B.n908 VSUBS 0.008148f
C949 B.n909 VSUBS 0.008148f
C950 B.n910 VSUBS 0.008148f
C951 B.n911 VSUBS 0.008148f
C952 B.n912 VSUBS 0.004554f
C953 B.n913 VSUBS 0.008148f
C954 B.n914 VSUBS 0.008148f
C955 B.n915 VSUBS 0.007669f
C956 B.n916 VSUBS 0.008148f
C957 B.n917 VSUBS 0.008148f
C958 B.n918 VSUBS 0.008148f
C959 B.n919 VSUBS 0.008148f
C960 B.n920 VSUBS 0.008148f
C961 B.n921 VSUBS 0.008148f
C962 B.n922 VSUBS 0.008148f
C963 B.n923 VSUBS 0.008148f
C964 B.n924 VSUBS 0.008148f
C965 B.n925 VSUBS 0.008148f
C966 B.n926 VSUBS 0.008148f
C967 B.n927 VSUBS 0.008148f
C968 B.n928 VSUBS 0.008148f
C969 B.n929 VSUBS 0.008148f
C970 B.n930 VSUBS 0.008148f
C971 B.n931 VSUBS 0.008148f
C972 B.n932 VSUBS 0.008148f
C973 B.n933 VSUBS 0.008148f
C974 B.n934 VSUBS 0.008148f
C975 B.n935 VSUBS 0.008148f
C976 B.n936 VSUBS 0.008148f
C977 B.n937 VSUBS 0.008148f
C978 B.n938 VSUBS 0.008148f
C979 B.n939 VSUBS 0.008148f
C980 B.n940 VSUBS 0.008148f
C981 B.n941 VSUBS 0.008148f
C982 B.n942 VSUBS 0.008148f
C983 B.n943 VSUBS 0.008148f
C984 B.n944 VSUBS 0.008148f
C985 B.n945 VSUBS 0.008148f
C986 B.n946 VSUBS 0.008148f
C987 B.n947 VSUBS 0.008148f
C988 B.n948 VSUBS 0.008148f
C989 B.n949 VSUBS 0.008148f
C990 B.n950 VSUBS 0.008148f
C991 B.n951 VSUBS 0.008148f
C992 B.n952 VSUBS 0.008148f
C993 B.n953 VSUBS 0.008148f
C994 B.n954 VSUBS 0.008148f
C995 B.n955 VSUBS 0.008148f
C996 B.n956 VSUBS 0.008148f
C997 B.n957 VSUBS 0.008148f
C998 B.n958 VSUBS 0.008148f
C999 B.n959 VSUBS 0.008148f
C1000 B.n960 VSUBS 0.008148f
C1001 B.n961 VSUBS 0.008148f
C1002 B.n962 VSUBS 0.008148f
C1003 B.n963 VSUBS 0.008148f
C1004 B.n964 VSUBS 0.008148f
C1005 B.n965 VSUBS 0.008148f
C1006 B.n966 VSUBS 0.008148f
C1007 B.n967 VSUBS 0.008148f
C1008 B.n968 VSUBS 0.008148f
C1009 B.n969 VSUBS 0.008148f
C1010 B.n970 VSUBS 0.008148f
C1011 B.n971 VSUBS 0.008148f
C1012 B.n972 VSUBS 0.008148f
C1013 B.n973 VSUBS 0.008148f
C1014 B.n974 VSUBS 0.008148f
C1015 B.n975 VSUBS 0.008148f
C1016 B.n976 VSUBS 0.008148f
C1017 B.n977 VSUBS 0.008148f
C1018 B.n978 VSUBS 0.008148f
C1019 B.n979 VSUBS 0.008148f
C1020 B.n980 VSUBS 0.008148f
C1021 B.n981 VSUBS 0.008148f
C1022 B.n982 VSUBS 0.008148f
C1023 B.n983 VSUBS 0.008148f
C1024 B.n984 VSUBS 0.008148f
C1025 B.n985 VSUBS 0.02f
C1026 B.n986 VSUBS 0.019304f
C1027 B.n987 VSUBS 0.019304f
C1028 B.n988 VSUBS 0.008148f
C1029 B.n989 VSUBS 0.008148f
C1030 B.n990 VSUBS 0.008148f
C1031 B.n991 VSUBS 0.008148f
C1032 B.n992 VSUBS 0.008148f
C1033 B.n993 VSUBS 0.008148f
C1034 B.n994 VSUBS 0.008148f
C1035 B.n995 VSUBS 0.008148f
C1036 B.n996 VSUBS 0.008148f
C1037 B.n997 VSUBS 0.008148f
C1038 B.n998 VSUBS 0.008148f
C1039 B.n999 VSUBS 0.008148f
C1040 B.n1000 VSUBS 0.008148f
C1041 B.n1001 VSUBS 0.008148f
C1042 B.n1002 VSUBS 0.008148f
C1043 B.n1003 VSUBS 0.008148f
C1044 B.n1004 VSUBS 0.008148f
C1045 B.n1005 VSUBS 0.008148f
C1046 B.n1006 VSUBS 0.008148f
C1047 B.n1007 VSUBS 0.008148f
C1048 B.n1008 VSUBS 0.008148f
C1049 B.n1009 VSUBS 0.008148f
C1050 B.n1010 VSUBS 0.008148f
C1051 B.n1011 VSUBS 0.008148f
C1052 B.n1012 VSUBS 0.008148f
C1053 B.n1013 VSUBS 0.008148f
C1054 B.n1014 VSUBS 0.008148f
C1055 B.n1015 VSUBS 0.008148f
C1056 B.n1016 VSUBS 0.008148f
C1057 B.n1017 VSUBS 0.008148f
C1058 B.n1018 VSUBS 0.008148f
C1059 B.n1019 VSUBS 0.008148f
C1060 B.n1020 VSUBS 0.008148f
C1061 B.n1021 VSUBS 0.008148f
C1062 B.n1022 VSUBS 0.008148f
C1063 B.n1023 VSUBS 0.008148f
C1064 B.n1024 VSUBS 0.008148f
C1065 B.n1025 VSUBS 0.008148f
C1066 B.n1026 VSUBS 0.008148f
C1067 B.n1027 VSUBS 0.008148f
C1068 B.n1028 VSUBS 0.008148f
C1069 B.n1029 VSUBS 0.008148f
C1070 B.n1030 VSUBS 0.008148f
C1071 B.n1031 VSUBS 0.008148f
C1072 B.n1032 VSUBS 0.008148f
C1073 B.n1033 VSUBS 0.008148f
C1074 B.n1034 VSUBS 0.008148f
C1075 B.n1035 VSUBS 0.008148f
C1076 B.n1036 VSUBS 0.008148f
C1077 B.n1037 VSUBS 0.008148f
C1078 B.n1038 VSUBS 0.008148f
C1079 B.n1039 VSUBS 0.008148f
C1080 B.n1040 VSUBS 0.008148f
C1081 B.n1041 VSUBS 0.008148f
C1082 B.n1042 VSUBS 0.008148f
C1083 B.n1043 VSUBS 0.008148f
C1084 B.n1044 VSUBS 0.008148f
C1085 B.n1045 VSUBS 0.008148f
C1086 B.n1046 VSUBS 0.008148f
C1087 B.n1047 VSUBS 0.008148f
C1088 B.n1048 VSUBS 0.008148f
C1089 B.n1049 VSUBS 0.008148f
C1090 B.n1050 VSUBS 0.008148f
C1091 B.n1051 VSUBS 0.008148f
C1092 B.n1052 VSUBS 0.008148f
C1093 B.n1053 VSUBS 0.008148f
C1094 B.n1054 VSUBS 0.008148f
C1095 B.n1055 VSUBS 0.008148f
C1096 B.n1056 VSUBS 0.008148f
C1097 B.n1057 VSUBS 0.008148f
C1098 B.n1058 VSUBS 0.008148f
C1099 B.n1059 VSUBS 0.008148f
C1100 B.n1060 VSUBS 0.008148f
C1101 B.n1061 VSUBS 0.008148f
C1102 B.n1062 VSUBS 0.008148f
C1103 B.n1063 VSUBS 0.008148f
C1104 B.n1064 VSUBS 0.008148f
C1105 B.n1065 VSUBS 0.008148f
C1106 B.n1066 VSUBS 0.008148f
C1107 B.n1067 VSUBS 0.008148f
C1108 B.n1068 VSUBS 0.008148f
C1109 B.n1069 VSUBS 0.008148f
C1110 B.n1070 VSUBS 0.008148f
C1111 B.n1071 VSUBS 0.008148f
C1112 B.n1072 VSUBS 0.008148f
C1113 B.n1073 VSUBS 0.008148f
C1114 B.n1074 VSUBS 0.008148f
C1115 B.n1075 VSUBS 0.008148f
C1116 B.n1076 VSUBS 0.008148f
C1117 B.n1077 VSUBS 0.008148f
C1118 B.n1078 VSUBS 0.008148f
C1119 B.n1079 VSUBS 0.008148f
C1120 B.n1080 VSUBS 0.008148f
C1121 B.n1081 VSUBS 0.008148f
C1122 B.n1082 VSUBS 0.008148f
C1123 B.n1083 VSUBS 0.008148f
C1124 B.n1084 VSUBS 0.008148f
C1125 B.n1085 VSUBS 0.008148f
C1126 B.n1086 VSUBS 0.008148f
C1127 B.n1087 VSUBS 0.008148f
C1128 B.n1088 VSUBS 0.008148f
C1129 B.n1089 VSUBS 0.008148f
C1130 B.n1090 VSUBS 0.008148f
C1131 B.n1091 VSUBS 0.008148f
C1132 B.n1092 VSUBS 0.008148f
C1133 B.n1093 VSUBS 0.008148f
C1134 B.n1094 VSUBS 0.008148f
C1135 B.n1095 VSUBS 0.008148f
C1136 B.n1096 VSUBS 0.008148f
C1137 B.n1097 VSUBS 0.008148f
C1138 B.n1098 VSUBS 0.008148f
C1139 B.n1099 VSUBS 0.008148f
C1140 B.n1100 VSUBS 0.008148f
C1141 B.n1101 VSUBS 0.008148f
C1142 B.n1102 VSUBS 0.008148f
C1143 B.n1103 VSUBS 0.008148f
C1144 B.n1104 VSUBS 0.008148f
C1145 B.n1105 VSUBS 0.008148f
C1146 B.n1106 VSUBS 0.008148f
C1147 B.n1107 VSUBS 0.008148f
C1148 B.n1108 VSUBS 0.008148f
C1149 B.n1109 VSUBS 0.008148f
C1150 B.n1110 VSUBS 0.008148f
C1151 B.n1111 VSUBS 0.010633f
C1152 B.n1112 VSUBS 0.011327f
C1153 B.n1113 VSUBS 0.022525f
C1154 VDD1.t0 VSUBS 3.65796f
C1155 VDD1.t7 VSUBS 0.344024f
C1156 VDD1.t9 VSUBS 0.344024f
C1157 VDD1.n0 VSUBS 2.7726f
C1158 VDD1.n1 VSUBS 2.05205f
C1159 VDD1.t1 VSUBS 3.65794f
C1160 VDD1.t4 VSUBS 0.344024f
C1161 VDD1.t5 VSUBS 0.344024f
C1162 VDD1.n2 VSUBS 2.7726f
C1163 VDD1.n3 VSUBS 2.04173f
C1164 VDD1.t2 VSUBS 0.344024f
C1165 VDD1.t3 VSUBS 0.344024f
C1166 VDD1.n4 VSUBS 2.8181f
C1167 VDD1.n5 VSUBS 5.12364f
C1168 VDD1.t8 VSUBS 0.344024f
C1169 VDD1.t6 VSUBS 0.344024f
C1170 VDD1.n6 VSUBS 2.77259f
C1171 VDD1.n7 VSUBS 5.11217f
C1172 VP.n0 VSUBS 0.043351f
C1173 VP.t6 VSUBS 3.60572f
C1174 VP.n1 VSUBS 0.042953f
C1175 VP.n2 VSUBS 0.023047f
C1176 VP.n3 VSUBS 0.042953f
C1177 VP.n4 VSUBS 0.023047f
C1178 VP.t7 VSUBS 3.60572f
C1179 VP.n5 VSUBS 0.042953f
C1180 VP.n6 VSUBS 0.023047f
C1181 VP.n7 VSUBS 0.042953f
C1182 VP.n8 VSUBS 0.023047f
C1183 VP.t4 VSUBS 3.60572f
C1184 VP.n9 VSUBS 0.042953f
C1185 VP.n10 VSUBS 0.023047f
C1186 VP.n11 VSUBS 0.046429f
C1187 VP.n12 VSUBS 0.023047f
C1188 VP.t5 VSUBS 3.60572f
C1189 VP.n13 VSUBS 1.25182f
C1190 VP.n14 VSUBS 0.023047f
C1191 VP.n15 VSUBS 0.033325f
C1192 VP.n16 VSUBS 0.023047f
C1193 VP.n17 VSUBS 0.039136f
C1194 VP.n18 VSUBS 0.043351f
C1195 VP.t3 VSUBS 3.60572f
C1196 VP.n19 VSUBS 0.042953f
C1197 VP.n20 VSUBS 0.023047f
C1198 VP.n21 VSUBS 0.042953f
C1199 VP.n22 VSUBS 0.023047f
C1200 VP.t1 VSUBS 3.60572f
C1201 VP.n23 VSUBS 0.042953f
C1202 VP.n24 VSUBS 0.023047f
C1203 VP.n25 VSUBS 0.042953f
C1204 VP.n26 VSUBS 0.023047f
C1205 VP.t0 VSUBS 3.60572f
C1206 VP.n27 VSUBS 0.042953f
C1207 VP.n28 VSUBS 0.023047f
C1208 VP.n29 VSUBS 0.046429f
C1209 VP.n30 VSUBS 0.023047f
C1210 VP.t2 VSUBS 3.60572f
C1211 VP.n31 VSUBS 1.32941f
C1212 VP.t9 VSUBS 3.99675f
C1213 VP.n32 VSUBS 1.26473f
C1214 VP.n33 VSUBS 0.308421f
C1215 VP.n34 VSUBS 0.02514f
C1216 VP.n35 VSUBS 0.042953f
C1217 VP.n36 VSUBS 0.042953f
C1218 VP.n37 VSUBS 0.023047f
C1219 VP.n38 VSUBS 0.023047f
C1220 VP.n39 VSUBS 0.023047f
C1221 VP.n40 VSUBS 0.020863f
C1222 VP.n41 VSUBS 0.042953f
C1223 VP.n42 VSUBS 0.042953f
C1224 VP.n43 VSUBS 0.023047f
C1225 VP.n44 VSUBS 0.023047f
C1226 VP.n45 VSUBS 0.023047f
C1227 VP.n46 VSUBS 0.03235f
C1228 VP.n47 VSUBS 1.25182f
C1229 VP.n48 VSUBS 0.03235f
C1230 VP.n49 VSUBS 0.042953f
C1231 VP.n50 VSUBS 0.023047f
C1232 VP.n51 VSUBS 0.023047f
C1233 VP.n52 VSUBS 0.023047f
C1234 VP.n53 VSUBS 0.042953f
C1235 VP.n54 VSUBS 0.020863f
C1236 VP.n55 VSUBS 0.046429f
C1237 VP.n56 VSUBS 0.023047f
C1238 VP.n57 VSUBS 0.023047f
C1239 VP.n58 VSUBS 0.023047f
C1240 VP.n59 VSUBS 0.042953f
C1241 VP.n60 VSUBS 0.02514f
C1242 VP.n61 VSUBS 1.25182f
C1243 VP.n62 VSUBS 0.03956f
C1244 VP.n63 VSUBS 0.023047f
C1245 VP.n64 VSUBS 0.023047f
C1246 VP.n65 VSUBS 0.023047f
C1247 VP.n66 VSUBS 0.042953f
C1248 VP.n67 VSUBS 0.033325f
C1249 VP.n68 VSUBS 0.033967f
C1250 VP.n69 VSUBS 0.023047f
C1251 VP.n70 VSUBS 0.023047f
C1252 VP.n71 VSUBS 0.023047f
C1253 VP.n72 VSUBS 0.042953f
C1254 VP.n73 VSUBS 0.039136f
C1255 VP.n74 VSUBS 1.35316f
C1256 VP.n75 VSUBS 1.82103f
C1257 VP.t8 VSUBS 3.60572f
C1258 VP.n76 VSUBS 1.35316f
C1259 VP.n77 VSUBS 1.83424f
C1260 VP.n78 VSUBS 0.043351f
C1261 VP.n79 VSUBS 0.023047f
C1262 VP.n80 VSUBS 0.042953f
C1263 VP.n81 VSUBS 0.042953f
C1264 VP.n82 VSUBS 0.033967f
C1265 VP.n83 VSUBS 0.023047f
C1266 VP.n84 VSUBS 0.023047f
C1267 VP.n85 VSUBS 0.023047f
C1268 VP.n86 VSUBS 0.042953f
C1269 VP.n87 VSUBS 0.042953f
C1270 VP.n88 VSUBS 0.03956f
C1271 VP.n89 VSUBS 0.023047f
C1272 VP.n90 VSUBS 0.023047f
C1273 VP.n91 VSUBS 0.02514f
C1274 VP.n92 VSUBS 0.042953f
C1275 VP.n93 VSUBS 0.042953f
C1276 VP.n94 VSUBS 0.023047f
C1277 VP.n95 VSUBS 0.023047f
C1278 VP.n96 VSUBS 0.023047f
C1279 VP.n97 VSUBS 0.020863f
C1280 VP.n98 VSUBS 0.042953f
C1281 VP.n99 VSUBS 0.042953f
C1282 VP.n100 VSUBS 0.023047f
C1283 VP.n101 VSUBS 0.023047f
C1284 VP.n102 VSUBS 0.023047f
C1285 VP.n103 VSUBS 0.03235f
C1286 VP.n104 VSUBS 1.25182f
C1287 VP.n105 VSUBS 0.03235f
C1288 VP.n106 VSUBS 0.042953f
C1289 VP.n107 VSUBS 0.023047f
C1290 VP.n108 VSUBS 0.023047f
C1291 VP.n109 VSUBS 0.023047f
C1292 VP.n110 VSUBS 0.042953f
C1293 VP.n111 VSUBS 0.020863f
C1294 VP.n112 VSUBS 0.046429f
C1295 VP.n113 VSUBS 0.023047f
C1296 VP.n114 VSUBS 0.023047f
C1297 VP.n115 VSUBS 0.023047f
C1298 VP.n116 VSUBS 0.042953f
C1299 VP.n117 VSUBS 0.02514f
C1300 VP.n118 VSUBS 1.25182f
C1301 VP.n119 VSUBS 0.03956f
C1302 VP.n120 VSUBS 0.023047f
C1303 VP.n121 VSUBS 0.023047f
C1304 VP.n122 VSUBS 0.023047f
C1305 VP.n123 VSUBS 0.042953f
C1306 VP.n124 VSUBS 0.033325f
C1307 VP.n125 VSUBS 0.033967f
C1308 VP.n126 VSUBS 0.023047f
C1309 VP.n127 VSUBS 0.023047f
C1310 VP.n128 VSUBS 0.023047f
C1311 VP.n129 VSUBS 0.042953f
C1312 VP.n130 VSUBS 0.039136f
C1313 VP.n131 VSUBS 1.35316f
C1314 VP.n132 VSUBS 0.073971f
C1315 VDD2.t5 VSUBS 3.65922f
C1316 VDD2.t1 VSUBS 0.344144f
C1317 VDD2.t7 VSUBS 0.344144f
C1318 VDD2.n0 VSUBS 2.77357f
C1319 VDD2.n1 VSUBS 2.04244f
C1320 VDD2.t2 VSUBS 0.344144f
C1321 VDD2.t3 VSUBS 0.344144f
C1322 VDD2.n2 VSUBS 2.81909f
C1323 VDD2.n3 VSUBS 4.92348f
C1324 VDD2.t6 VSUBS 3.60794f
C1325 VDD2.n4 VSUBS 5.03835f
C1326 VDD2.t8 VSUBS 0.344144f
C1327 VDD2.t9 VSUBS 0.344144f
C1328 VDD2.n5 VSUBS 2.77357f
C1329 VDD2.n6 VSUBS 1.04247f
C1330 VDD2.t0 VSUBS 0.344144f
C1331 VDD2.t4 VSUBS 0.344144f
C1332 VDD2.n7 VSUBS 2.81901f
C1333 VTAIL.t16 VSUBS 0.330981f
C1334 VTAIL.t15 VSUBS 0.330981f
C1335 VTAIL.n0 VSUBS 2.49908f
C1336 VTAIL.n1 VSUBS 1.17553f
C1337 VTAIL.t9 VSUBS 3.27884f
C1338 VTAIL.n2 VSUBS 1.38109f
C1339 VTAIL.t7 VSUBS 0.330981f
C1340 VTAIL.t0 VSUBS 0.330981f
C1341 VTAIL.n3 VSUBS 2.49908f
C1342 VTAIL.n4 VSUBS 1.39007f
C1343 VTAIL.t6 VSUBS 0.330981f
C1344 VTAIL.t5 VSUBS 0.330981f
C1345 VTAIL.n5 VSUBS 2.49908f
C1346 VTAIL.n6 VSUBS 3.30419f
C1347 VTAIL.t19 VSUBS 0.330981f
C1348 VTAIL.t13 VSUBS 0.330981f
C1349 VTAIL.n7 VSUBS 2.49908f
C1350 VTAIL.n8 VSUBS 3.30419f
C1351 VTAIL.t18 VSUBS 0.330981f
C1352 VTAIL.t10 VSUBS 0.330981f
C1353 VTAIL.n9 VSUBS 2.49908f
C1354 VTAIL.n10 VSUBS 1.39006f
C1355 VTAIL.t11 VSUBS 3.27886f
C1356 VTAIL.n11 VSUBS 1.38106f
C1357 VTAIL.t8 VSUBS 0.330981f
C1358 VTAIL.t4 VSUBS 0.330981f
C1359 VTAIL.n12 VSUBS 2.49908f
C1360 VTAIL.n13 VSUBS 1.25817f
C1361 VTAIL.t1 VSUBS 0.330981f
C1362 VTAIL.t2 VSUBS 0.330981f
C1363 VTAIL.n14 VSUBS 2.49908f
C1364 VTAIL.n15 VSUBS 1.39006f
C1365 VTAIL.t3 VSUBS 3.27884f
C1366 VTAIL.n16 VSUBS 3.07458f
C1367 VTAIL.t17 VSUBS 3.27884f
C1368 VTAIL.n17 VSUBS 3.07458f
C1369 VTAIL.t12 VSUBS 0.330981f
C1370 VTAIL.t14 VSUBS 0.330981f
C1371 VTAIL.n18 VSUBS 2.49908f
C1372 VTAIL.n19 VSUBS 1.12017f
C1373 VN.n0 VSUBS 0.039994f
C1374 VN.t6 VSUBS 3.32647f
C1375 VN.n1 VSUBS 0.039627f
C1376 VN.n2 VSUBS 0.021262f
C1377 VN.n3 VSUBS 0.039627f
C1378 VN.n4 VSUBS 0.021262f
C1379 VN.t7 VSUBS 3.32647f
C1380 VN.n5 VSUBS 0.039627f
C1381 VN.n6 VSUBS 0.021262f
C1382 VN.n7 VSUBS 0.039627f
C1383 VN.n8 VSUBS 0.021262f
C1384 VN.t2 VSUBS 3.32647f
C1385 VN.n9 VSUBS 0.039627f
C1386 VN.n10 VSUBS 0.021262f
C1387 VN.n11 VSUBS 0.042833f
C1388 VN.n12 VSUBS 0.021262f
C1389 VN.t8 VSUBS 3.32647f
C1390 VN.n13 VSUBS 1.22645f
C1391 VN.t4 VSUBS 3.68722f
C1392 VN.n14 VSUBS 1.16678f
C1393 VN.n15 VSUBS 0.284534f
C1394 VN.n16 VSUBS 0.023193f
C1395 VN.n17 VSUBS 0.039627f
C1396 VN.n18 VSUBS 0.039627f
C1397 VN.n19 VSUBS 0.021262f
C1398 VN.n20 VSUBS 0.021262f
C1399 VN.n21 VSUBS 0.021262f
C1400 VN.n22 VSUBS 0.019248f
C1401 VN.n23 VSUBS 0.039627f
C1402 VN.n24 VSUBS 0.039627f
C1403 VN.n25 VSUBS 0.021262f
C1404 VN.n26 VSUBS 0.021262f
C1405 VN.n27 VSUBS 0.021262f
C1406 VN.n28 VSUBS 0.029845f
C1407 VN.n29 VSUBS 1.15487f
C1408 VN.n30 VSUBS 0.029845f
C1409 VN.n31 VSUBS 0.039627f
C1410 VN.n32 VSUBS 0.021262f
C1411 VN.n33 VSUBS 0.021262f
C1412 VN.n34 VSUBS 0.021262f
C1413 VN.n35 VSUBS 0.039627f
C1414 VN.n36 VSUBS 0.019248f
C1415 VN.n37 VSUBS 0.042833f
C1416 VN.n38 VSUBS 0.021262f
C1417 VN.n39 VSUBS 0.021262f
C1418 VN.n40 VSUBS 0.021262f
C1419 VN.n41 VSUBS 0.039627f
C1420 VN.n42 VSUBS 0.023193f
C1421 VN.n43 VSUBS 1.15487f
C1422 VN.n44 VSUBS 0.036497f
C1423 VN.n45 VSUBS 0.021262f
C1424 VN.n46 VSUBS 0.021262f
C1425 VN.n47 VSUBS 0.021262f
C1426 VN.n48 VSUBS 0.039627f
C1427 VN.n49 VSUBS 0.030744f
C1428 VN.n50 VSUBS 0.031337f
C1429 VN.n51 VSUBS 0.021262f
C1430 VN.n52 VSUBS 0.021262f
C1431 VN.n53 VSUBS 0.021262f
C1432 VN.n54 VSUBS 0.039627f
C1433 VN.n55 VSUBS 0.036105f
C1434 VN.n56 VSUBS 1.24836f
C1435 VN.n57 VSUBS 0.068242f
C1436 VN.n58 VSUBS 0.039994f
C1437 VN.t3 VSUBS 3.32647f
C1438 VN.n59 VSUBS 0.039627f
C1439 VN.n60 VSUBS 0.021262f
C1440 VN.n61 VSUBS 0.039627f
C1441 VN.n62 VSUBS 0.021262f
C1442 VN.t1 VSUBS 3.32647f
C1443 VN.n63 VSUBS 0.039627f
C1444 VN.n64 VSUBS 0.021262f
C1445 VN.n65 VSUBS 0.039627f
C1446 VN.n66 VSUBS 0.021262f
C1447 VN.t0 VSUBS 3.32647f
C1448 VN.n67 VSUBS 0.039627f
C1449 VN.n68 VSUBS 0.021262f
C1450 VN.n69 VSUBS 0.042833f
C1451 VN.n70 VSUBS 0.021262f
C1452 VN.t9 VSUBS 3.32647f
C1453 VN.n71 VSUBS 1.22645f
C1454 VN.t5 VSUBS 3.68722f
C1455 VN.n72 VSUBS 1.16678f
C1456 VN.n73 VSUBS 0.284534f
C1457 VN.n74 VSUBS 0.023193f
C1458 VN.n75 VSUBS 0.039627f
C1459 VN.n76 VSUBS 0.039627f
C1460 VN.n77 VSUBS 0.021262f
C1461 VN.n78 VSUBS 0.021262f
C1462 VN.n79 VSUBS 0.021262f
C1463 VN.n80 VSUBS 0.019248f
C1464 VN.n81 VSUBS 0.039627f
C1465 VN.n82 VSUBS 0.039627f
C1466 VN.n83 VSUBS 0.021262f
C1467 VN.n84 VSUBS 0.021262f
C1468 VN.n85 VSUBS 0.021262f
C1469 VN.n86 VSUBS 0.029845f
C1470 VN.n87 VSUBS 1.15487f
C1471 VN.n88 VSUBS 0.029845f
C1472 VN.n89 VSUBS 0.039627f
C1473 VN.n90 VSUBS 0.021262f
C1474 VN.n91 VSUBS 0.021262f
C1475 VN.n92 VSUBS 0.021262f
C1476 VN.n93 VSUBS 0.039627f
C1477 VN.n94 VSUBS 0.019248f
C1478 VN.n95 VSUBS 0.042833f
C1479 VN.n96 VSUBS 0.021262f
C1480 VN.n97 VSUBS 0.021262f
C1481 VN.n98 VSUBS 0.021262f
C1482 VN.n99 VSUBS 0.039627f
C1483 VN.n100 VSUBS 0.023193f
C1484 VN.n101 VSUBS 1.15487f
C1485 VN.n102 VSUBS 0.036497f
C1486 VN.n103 VSUBS 0.021262f
C1487 VN.n104 VSUBS 0.021262f
C1488 VN.n105 VSUBS 0.021262f
C1489 VN.n106 VSUBS 0.039627f
C1490 VN.n107 VSUBS 0.030744f
C1491 VN.n108 VSUBS 0.031337f
C1492 VN.n109 VSUBS 0.021262f
C1493 VN.n110 VSUBS 0.021262f
C1494 VN.n111 VSUBS 0.021262f
C1495 VN.n112 VSUBS 0.039627f
C1496 VN.n113 VSUBS 0.036105f
C1497 VN.n114 VSUBS 1.24836f
C1498 VN.n115 VSUBS 1.6847f
.ends

