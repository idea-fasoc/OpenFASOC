* NGSPICE file created from diff_pair_sample_0836.ext - technology: sky130A

.subckt diff_pair_sample_0836 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t9 VN.t0 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.4157 pd=8.91 as=1.4157 ps=8.91 w=8.58 l=0.64
X1 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=3.3462 pd=17.94 as=0 ps=0 w=8.58 l=0.64
X2 VDD1.t5 VP.t0 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=3.3462 pd=17.94 as=1.4157 ps=8.91 w=8.58 l=0.64
X3 VDD2.t5 VN.t1 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=3.3462 pd=17.94 as=1.4157 ps=8.91 w=8.58 l=0.64
X4 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=3.3462 pd=17.94 as=0 ps=0 w=8.58 l=0.64
X5 VDD1.t4 VP.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.3462 pd=17.94 as=1.4157 ps=8.91 w=8.58 l=0.64
X6 VDD2.t3 VN.t2 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=3.3462 pd=17.94 as=1.4157 ps=8.91 w=8.58 l=0.64
X7 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=3.3462 pd=17.94 as=0 ps=0 w=8.58 l=0.64
X8 VTAIL.t11 VP.t2 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.4157 pd=8.91 as=1.4157 ps=8.91 w=8.58 l=0.64
X9 VDD2.t2 VN.t3 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4157 pd=8.91 as=3.3462 ps=17.94 w=8.58 l=0.64
X10 VDD2.t0 VN.t4 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.4157 pd=8.91 as=3.3462 ps=17.94 w=8.58 l=0.64
X11 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.3462 pd=17.94 as=0 ps=0 w=8.58 l=0.64
X12 VTAIL.t0 VP.t3 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.4157 pd=8.91 as=1.4157 ps=8.91 w=8.58 l=0.64
X13 VTAIL.t4 VN.t5 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.4157 pd=8.91 as=1.4157 ps=8.91 w=8.58 l=0.64
X14 VDD1.t1 VP.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4157 pd=8.91 as=3.3462 ps=17.94 w=8.58 l=0.64
X15 VDD1.t0 VP.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.4157 pd=8.91 as=3.3462 ps=17.94 w=8.58 l=0.64
R0 VN.n0 VN.t1 411.291
R1 VN.n4 VN.t4 411.291
R2 VN.n1 VN.t5 384.471
R3 VN.n2 VN.t3 384.471
R4 VN.n5 VN.t0 384.471
R5 VN.n6 VN.t2 384.471
R6 VN.n3 VN.n2 161.3
R7 VN.n7 VN.n6 161.3
R8 VN.n2 VN.n1 48.2005
R9 VN.n6 VN.n5 48.2005
R10 VN.n7 VN.n4 45.1367
R11 VN.n3 VN.n0 45.1367
R12 VN VN.n7 38.885
R13 VN.n5 VN.n4 13.3799
R14 VN.n1 VN.n0 13.3799
R15 VN VN.n3 0.0516364
R16 VDD2.n87 VDD2.n47 289.615
R17 VDD2.n40 VDD2.n0 289.615
R18 VDD2.n88 VDD2.n87 185
R19 VDD2.n86 VDD2.n85 185
R20 VDD2.n84 VDD2.n50 185
R21 VDD2.n54 VDD2.n51 185
R22 VDD2.n79 VDD2.n78 185
R23 VDD2.n77 VDD2.n76 185
R24 VDD2.n56 VDD2.n55 185
R25 VDD2.n71 VDD2.n70 185
R26 VDD2.n69 VDD2.n68 185
R27 VDD2.n60 VDD2.n59 185
R28 VDD2.n63 VDD2.n62 185
R29 VDD2.n15 VDD2.n14 185
R30 VDD2.n12 VDD2.n11 185
R31 VDD2.n21 VDD2.n20 185
R32 VDD2.n23 VDD2.n22 185
R33 VDD2.n8 VDD2.n7 185
R34 VDD2.n29 VDD2.n28 185
R35 VDD2.n32 VDD2.n31 185
R36 VDD2.n30 VDD2.n4 185
R37 VDD2.n37 VDD2.n3 185
R38 VDD2.n39 VDD2.n38 185
R39 VDD2.n41 VDD2.n40 185
R40 VDD2.t3 VDD2.n61 149.524
R41 VDD2.t5 VDD2.n13 149.524
R42 VDD2.n87 VDD2.n86 104.615
R43 VDD2.n86 VDD2.n50 104.615
R44 VDD2.n54 VDD2.n50 104.615
R45 VDD2.n78 VDD2.n54 104.615
R46 VDD2.n78 VDD2.n77 104.615
R47 VDD2.n77 VDD2.n55 104.615
R48 VDD2.n70 VDD2.n55 104.615
R49 VDD2.n70 VDD2.n69 104.615
R50 VDD2.n69 VDD2.n59 104.615
R51 VDD2.n62 VDD2.n59 104.615
R52 VDD2.n14 VDD2.n11 104.615
R53 VDD2.n21 VDD2.n11 104.615
R54 VDD2.n22 VDD2.n21 104.615
R55 VDD2.n22 VDD2.n7 104.615
R56 VDD2.n29 VDD2.n7 104.615
R57 VDD2.n31 VDD2.n29 104.615
R58 VDD2.n31 VDD2.n30 104.615
R59 VDD2.n30 VDD2.n3 104.615
R60 VDD2.n39 VDD2.n3 104.615
R61 VDD2.n40 VDD2.n39 104.615
R62 VDD2.n46 VDD2.n45 64.7584
R63 VDD2 VDD2.n93 64.7555
R64 VDD2.n62 VDD2.t3 52.3082
R65 VDD2.n14 VDD2.t5 52.3082
R66 VDD2.n46 VDD2.n44 50.5996
R67 VDD2.n92 VDD2.n91 50.0278
R68 VDD2.n92 VDD2.n46 33.8295
R69 VDD2.n85 VDD2.n84 13.1884
R70 VDD2.n38 VDD2.n37 13.1884
R71 VDD2.n88 VDD2.n49 12.8005
R72 VDD2.n83 VDD2.n51 12.8005
R73 VDD2.n36 VDD2.n4 12.8005
R74 VDD2.n41 VDD2.n2 12.8005
R75 VDD2.n89 VDD2.n47 12.0247
R76 VDD2.n80 VDD2.n79 12.0247
R77 VDD2.n33 VDD2.n32 12.0247
R78 VDD2.n42 VDD2.n0 12.0247
R79 VDD2.n76 VDD2.n53 11.249
R80 VDD2.n28 VDD2.n6 11.249
R81 VDD2.n75 VDD2.n56 10.4732
R82 VDD2.n27 VDD2.n8 10.4732
R83 VDD2.n63 VDD2.n61 10.2747
R84 VDD2.n15 VDD2.n13 10.2747
R85 VDD2.n72 VDD2.n71 9.69747
R86 VDD2.n24 VDD2.n23 9.69747
R87 VDD2.n91 VDD2.n90 9.45567
R88 VDD2.n44 VDD2.n43 9.45567
R89 VDD2.n65 VDD2.n64 9.3005
R90 VDD2.n67 VDD2.n66 9.3005
R91 VDD2.n58 VDD2.n57 9.3005
R92 VDD2.n73 VDD2.n72 9.3005
R93 VDD2.n75 VDD2.n74 9.3005
R94 VDD2.n53 VDD2.n52 9.3005
R95 VDD2.n81 VDD2.n80 9.3005
R96 VDD2.n83 VDD2.n82 9.3005
R97 VDD2.n90 VDD2.n89 9.3005
R98 VDD2.n49 VDD2.n48 9.3005
R99 VDD2.n43 VDD2.n42 9.3005
R100 VDD2.n2 VDD2.n1 9.3005
R101 VDD2.n17 VDD2.n16 9.3005
R102 VDD2.n19 VDD2.n18 9.3005
R103 VDD2.n10 VDD2.n9 9.3005
R104 VDD2.n25 VDD2.n24 9.3005
R105 VDD2.n27 VDD2.n26 9.3005
R106 VDD2.n6 VDD2.n5 9.3005
R107 VDD2.n34 VDD2.n33 9.3005
R108 VDD2.n36 VDD2.n35 9.3005
R109 VDD2.n68 VDD2.n58 8.92171
R110 VDD2.n20 VDD2.n10 8.92171
R111 VDD2.n67 VDD2.n60 8.14595
R112 VDD2.n19 VDD2.n12 8.14595
R113 VDD2.n64 VDD2.n63 7.3702
R114 VDD2.n16 VDD2.n15 7.3702
R115 VDD2.n64 VDD2.n60 5.81868
R116 VDD2.n16 VDD2.n12 5.81868
R117 VDD2.n68 VDD2.n67 5.04292
R118 VDD2.n20 VDD2.n19 5.04292
R119 VDD2.n71 VDD2.n58 4.26717
R120 VDD2.n23 VDD2.n10 4.26717
R121 VDD2.n72 VDD2.n56 3.49141
R122 VDD2.n24 VDD2.n8 3.49141
R123 VDD2.n17 VDD2.n13 2.84303
R124 VDD2.n65 VDD2.n61 2.84303
R125 VDD2.n76 VDD2.n75 2.71565
R126 VDD2.n28 VDD2.n27 2.71565
R127 VDD2.n93 VDD2.t4 2.30819
R128 VDD2.n93 VDD2.t0 2.30819
R129 VDD2.n45 VDD2.t1 2.30819
R130 VDD2.n45 VDD2.t2 2.30819
R131 VDD2.n91 VDD2.n47 1.93989
R132 VDD2.n79 VDD2.n53 1.93989
R133 VDD2.n32 VDD2.n6 1.93989
R134 VDD2.n44 VDD2.n0 1.93989
R135 VDD2.n89 VDD2.n88 1.16414
R136 VDD2.n80 VDD2.n51 1.16414
R137 VDD2.n33 VDD2.n4 1.16414
R138 VDD2.n42 VDD2.n41 1.16414
R139 VDD2 VDD2.n92 0.685845
R140 VDD2.n85 VDD2.n49 0.388379
R141 VDD2.n84 VDD2.n83 0.388379
R142 VDD2.n37 VDD2.n36 0.388379
R143 VDD2.n38 VDD2.n2 0.388379
R144 VDD2.n90 VDD2.n48 0.155672
R145 VDD2.n82 VDD2.n48 0.155672
R146 VDD2.n82 VDD2.n81 0.155672
R147 VDD2.n81 VDD2.n52 0.155672
R148 VDD2.n74 VDD2.n52 0.155672
R149 VDD2.n74 VDD2.n73 0.155672
R150 VDD2.n73 VDD2.n57 0.155672
R151 VDD2.n66 VDD2.n57 0.155672
R152 VDD2.n66 VDD2.n65 0.155672
R153 VDD2.n18 VDD2.n17 0.155672
R154 VDD2.n18 VDD2.n9 0.155672
R155 VDD2.n25 VDD2.n9 0.155672
R156 VDD2.n26 VDD2.n25 0.155672
R157 VDD2.n26 VDD2.n5 0.155672
R158 VDD2.n34 VDD2.n5 0.155672
R159 VDD2.n35 VDD2.n34 0.155672
R160 VDD2.n35 VDD2.n1 0.155672
R161 VDD2.n43 VDD2.n1 0.155672
R162 VTAIL.n186 VTAIL.n146 289.615
R163 VTAIL.n42 VTAIL.n2 289.615
R164 VTAIL.n140 VTAIL.n100 289.615
R165 VTAIL.n92 VTAIL.n52 289.615
R166 VTAIL.n161 VTAIL.n160 185
R167 VTAIL.n158 VTAIL.n157 185
R168 VTAIL.n167 VTAIL.n166 185
R169 VTAIL.n169 VTAIL.n168 185
R170 VTAIL.n154 VTAIL.n153 185
R171 VTAIL.n175 VTAIL.n174 185
R172 VTAIL.n178 VTAIL.n177 185
R173 VTAIL.n176 VTAIL.n150 185
R174 VTAIL.n183 VTAIL.n149 185
R175 VTAIL.n185 VTAIL.n184 185
R176 VTAIL.n187 VTAIL.n186 185
R177 VTAIL.n17 VTAIL.n16 185
R178 VTAIL.n14 VTAIL.n13 185
R179 VTAIL.n23 VTAIL.n22 185
R180 VTAIL.n25 VTAIL.n24 185
R181 VTAIL.n10 VTAIL.n9 185
R182 VTAIL.n31 VTAIL.n30 185
R183 VTAIL.n34 VTAIL.n33 185
R184 VTAIL.n32 VTAIL.n6 185
R185 VTAIL.n39 VTAIL.n5 185
R186 VTAIL.n41 VTAIL.n40 185
R187 VTAIL.n43 VTAIL.n42 185
R188 VTAIL.n141 VTAIL.n140 185
R189 VTAIL.n139 VTAIL.n138 185
R190 VTAIL.n137 VTAIL.n103 185
R191 VTAIL.n107 VTAIL.n104 185
R192 VTAIL.n132 VTAIL.n131 185
R193 VTAIL.n130 VTAIL.n129 185
R194 VTAIL.n109 VTAIL.n108 185
R195 VTAIL.n124 VTAIL.n123 185
R196 VTAIL.n122 VTAIL.n121 185
R197 VTAIL.n113 VTAIL.n112 185
R198 VTAIL.n116 VTAIL.n115 185
R199 VTAIL.n93 VTAIL.n92 185
R200 VTAIL.n91 VTAIL.n90 185
R201 VTAIL.n89 VTAIL.n55 185
R202 VTAIL.n59 VTAIL.n56 185
R203 VTAIL.n84 VTAIL.n83 185
R204 VTAIL.n82 VTAIL.n81 185
R205 VTAIL.n61 VTAIL.n60 185
R206 VTAIL.n76 VTAIL.n75 185
R207 VTAIL.n74 VTAIL.n73 185
R208 VTAIL.n65 VTAIL.n64 185
R209 VTAIL.n68 VTAIL.n67 185
R210 VTAIL.t6 VTAIL.n159 149.524
R211 VTAIL.t2 VTAIL.n15 149.524
R212 VTAIL.t1 VTAIL.n114 149.524
R213 VTAIL.t5 VTAIL.n66 149.524
R214 VTAIL.n160 VTAIL.n157 104.615
R215 VTAIL.n167 VTAIL.n157 104.615
R216 VTAIL.n168 VTAIL.n167 104.615
R217 VTAIL.n168 VTAIL.n153 104.615
R218 VTAIL.n175 VTAIL.n153 104.615
R219 VTAIL.n177 VTAIL.n175 104.615
R220 VTAIL.n177 VTAIL.n176 104.615
R221 VTAIL.n176 VTAIL.n149 104.615
R222 VTAIL.n185 VTAIL.n149 104.615
R223 VTAIL.n186 VTAIL.n185 104.615
R224 VTAIL.n16 VTAIL.n13 104.615
R225 VTAIL.n23 VTAIL.n13 104.615
R226 VTAIL.n24 VTAIL.n23 104.615
R227 VTAIL.n24 VTAIL.n9 104.615
R228 VTAIL.n31 VTAIL.n9 104.615
R229 VTAIL.n33 VTAIL.n31 104.615
R230 VTAIL.n33 VTAIL.n32 104.615
R231 VTAIL.n32 VTAIL.n5 104.615
R232 VTAIL.n41 VTAIL.n5 104.615
R233 VTAIL.n42 VTAIL.n41 104.615
R234 VTAIL.n140 VTAIL.n139 104.615
R235 VTAIL.n139 VTAIL.n103 104.615
R236 VTAIL.n107 VTAIL.n103 104.615
R237 VTAIL.n131 VTAIL.n107 104.615
R238 VTAIL.n131 VTAIL.n130 104.615
R239 VTAIL.n130 VTAIL.n108 104.615
R240 VTAIL.n123 VTAIL.n108 104.615
R241 VTAIL.n123 VTAIL.n122 104.615
R242 VTAIL.n122 VTAIL.n112 104.615
R243 VTAIL.n115 VTAIL.n112 104.615
R244 VTAIL.n92 VTAIL.n91 104.615
R245 VTAIL.n91 VTAIL.n55 104.615
R246 VTAIL.n59 VTAIL.n55 104.615
R247 VTAIL.n83 VTAIL.n59 104.615
R248 VTAIL.n83 VTAIL.n82 104.615
R249 VTAIL.n82 VTAIL.n60 104.615
R250 VTAIL.n75 VTAIL.n60 104.615
R251 VTAIL.n75 VTAIL.n74 104.615
R252 VTAIL.n74 VTAIL.n64 104.615
R253 VTAIL.n67 VTAIL.n64 104.615
R254 VTAIL.n160 VTAIL.t6 52.3082
R255 VTAIL.n16 VTAIL.t2 52.3082
R256 VTAIL.n115 VTAIL.t1 52.3082
R257 VTAIL.n67 VTAIL.t5 52.3082
R258 VTAIL.n99 VTAIL.n98 47.926
R259 VTAIL.n51 VTAIL.n50 47.926
R260 VTAIL.n1 VTAIL.n0 47.9259
R261 VTAIL.n49 VTAIL.n48 47.9259
R262 VTAIL.n191 VTAIL.n190 33.349
R263 VTAIL.n47 VTAIL.n46 33.349
R264 VTAIL.n145 VTAIL.n144 33.349
R265 VTAIL.n97 VTAIL.n96 33.349
R266 VTAIL.n51 VTAIL.n49 21.4358
R267 VTAIL.n191 VTAIL.n145 20.5996
R268 VTAIL.n184 VTAIL.n183 13.1884
R269 VTAIL.n40 VTAIL.n39 13.1884
R270 VTAIL.n138 VTAIL.n137 13.1884
R271 VTAIL.n90 VTAIL.n89 13.1884
R272 VTAIL.n182 VTAIL.n150 12.8005
R273 VTAIL.n187 VTAIL.n148 12.8005
R274 VTAIL.n38 VTAIL.n6 12.8005
R275 VTAIL.n43 VTAIL.n4 12.8005
R276 VTAIL.n141 VTAIL.n102 12.8005
R277 VTAIL.n136 VTAIL.n104 12.8005
R278 VTAIL.n93 VTAIL.n54 12.8005
R279 VTAIL.n88 VTAIL.n56 12.8005
R280 VTAIL.n179 VTAIL.n178 12.0247
R281 VTAIL.n188 VTAIL.n146 12.0247
R282 VTAIL.n35 VTAIL.n34 12.0247
R283 VTAIL.n44 VTAIL.n2 12.0247
R284 VTAIL.n142 VTAIL.n100 12.0247
R285 VTAIL.n133 VTAIL.n132 12.0247
R286 VTAIL.n94 VTAIL.n52 12.0247
R287 VTAIL.n85 VTAIL.n84 12.0247
R288 VTAIL.n174 VTAIL.n152 11.249
R289 VTAIL.n30 VTAIL.n8 11.249
R290 VTAIL.n129 VTAIL.n106 11.249
R291 VTAIL.n81 VTAIL.n58 11.249
R292 VTAIL.n173 VTAIL.n154 10.4732
R293 VTAIL.n29 VTAIL.n10 10.4732
R294 VTAIL.n128 VTAIL.n109 10.4732
R295 VTAIL.n80 VTAIL.n61 10.4732
R296 VTAIL.n161 VTAIL.n159 10.2747
R297 VTAIL.n17 VTAIL.n15 10.2747
R298 VTAIL.n116 VTAIL.n114 10.2747
R299 VTAIL.n68 VTAIL.n66 10.2747
R300 VTAIL.n170 VTAIL.n169 9.69747
R301 VTAIL.n26 VTAIL.n25 9.69747
R302 VTAIL.n125 VTAIL.n124 9.69747
R303 VTAIL.n77 VTAIL.n76 9.69747
R304 VTAIL.n190 VTAIL.n189 9.45567
R305 VTAIL.n46 VTAIL.n45 9.45567
R306 VTAIL.n144 VTAIL.n143 9.45567
R307 VTAIL.n96 VTAIL.n95 9.45567
R308 VTAIL.n189 VTAIL.n188 9.3005
R309 VTAIL.n148 VTAIL.n147 9.3005
R310 VTAIL.n163 VTAIL.n162 9.3005
R311 VTAIL.n165 VTAIL.n164 9.3005
R312 VTAIL.n156 VTAIL.n155 9.3005
R313 VTAIL.n171 VTAIL.n170 9.3005
R314 VTAIL.n173 VTAIL.n172 9.3005
R315 VTAIL.n152 VTAIL.n151 9.3005
R316 VTAIL.n180 VTAIL.n179 9.3005
R317 VTAIL.n182 VTAIL.n181 9.3005
R318 VTAIL.n45 VTAIL.n44 9.3005
R319 VTAIL.n4 VTAIL.n3 9.3005
R320 VTAIL.n19 VTAIL.n18 9.3005
R321 VTAIL.n21 VTAIL.n20 9.3005
R322 VTAIL.n12 VTAIL.n11 9.3005
R323 VTAIL.n27 VTAIL.n26 9.3005
R324 VTAIL.n29 VTAIL.n28 9.3005
R325 VTAIL.n8 VTAIL.n7 9.3005
R326 VTAIL.n36 VTAIL.n35 9.3005
R327 VTAIL.n38 VTAIL.n37 9.3005
R328 VTAIL.n118 VTAIL.n117 9.3005
R329 VTAIL.n120 VTAIL.n119 9.3005
R330 VTAIL.n111 VTAIL.n110 9.3005
R331 VTAIL.n126 VTAIL.n125 9.3005
R332 VTAIL.n128 VTAIL.n127 9.3005
R333 VTAIL.n106 VTAIL.n105 9.3005
R334 VTAIL.n134 VTAIL.n133 9.3005
R335 VTAIL.n136 VTAIL.n135 9.3005
R336 VTAIL.n143 VTAIL.n142 9.3005
R337 VTAIL.n102 VTAIL.n101 9.3005
R338 VTAIL.n70 VTAIL.n69 9.3005
R339 VTAIL.n72 VTAIL.n71 9.3005
R340 VTAIL.n63 VTAIL.n62 9.3005
R341 VTAIL.n78 VTAIL.n77 9.3005
R342 VTAIL.n80 VTAIL.n79 9.3005
R343 VTAIL.n58 VTAIL.n57 9.3005
R344 VTAIL.n86 VTAIL.n85 9.3005
R345 VTAIL.n88 VTAIL.n87 9.3005
R346 VTAIL.n95 VTAIL.n94 9.3005
R347 VTAIL.n54 VTAIL.n53 9.3005
R348 VTAIL.n166 VTAIL.n156 8.92171
R349 VTAIL.n22 VTAIL.n12 8.92171
R350 VTAIL.n121 VTAIL.n111 8.92171
R351 VTAIL.n73 VTAIL.n63 8.92171
R352 VTAIL.n165 VTAIL.n158 8.14595
R353 VTAIL.n21 VTAIL.n14 8.14595
R354 VTAIL.n120 VTAIL.n113 8.14595
R355 VTAIL.n72 VTAIL.n65 8.14595
R356 VTAIL.n162 VTAIL.n161 7.3702
R357 VTAIL.n18 VTAIL.n17 7.3702
R358 VTAIL.n117 VTAIL.n116 7.3702
R359 VTAIL.n69 VTAIL.n68 7.3702
R360 VTAIL.n162 VTAIL.n158 5.81868
R361 VTAIL.n18 VTAIL.n14 5.81868
R362 VTAIL.n117 VTAIL.n113 5.81868
R363 VTAIL.n69 VTAIL.n65 5.81868
R364 VTAIL.n166 VTAIL.n165 5.04292
R365 VTAIL.n22 VTAIL.n21 5.04292
R366 VTAIL.n121 VTAIL.n120 5.04292
R367 VTAIL.n73 VTAIL.n72 5.04292
R368 VTAIL.n169 VTAIL.n156 4.26717
R369 VTAIL.n25 VTAIL.n12 4.26717
R370 VTAIL.n124 VTAIL.n111 4.26717
R371 VTAIL.n76 VTAIL.n63 4.26717
R372 VTAIL.n170 VTAIL.n154 3.49141
R373 VTAIL.n26 VTAIL.n10 3.49141
R374 VTAIL.n125 VTAIL.n109 3.49141
R375 VTAIL.n77 VTAIL.n61 3.49141
R376 VTAIL.n163 VTAIL.n159 2.84303
R377 VTAIL.n19 VTAIL.n15 2.84303
R378 VTAIL.n118 VTAIL.n114 2.84303
R379 VTAIL.n70 VTAIL.n66 2.84303
R380 VTAIL.n174 VTAIL.n173 2.71565
R381 VTAIL.n30 VTAIL.n29 2.71565
R382 VTAIL.n129 VTAIL.n128 2.71565
R383 VTAIL.n81 VTAIL.n80 2.71565
R384 VTAIL.n0 VTAIL.t8 2.30819
R385 VTAIL.n0 VTAIL.t4 2.30819
R386 VTAIL.n48 VTAIL.t3 2.30819
R387 VTAIL.n48 VTAIL.t0 2.30819
R388 VTAIL.n98 VTAIL.t10 2.30819
R389 VTAIL.n98 VTAIL.t11 2.30819
R390 VTAIL.n50 VTAIL.t7 2.30819
R391 VTAIL.n50 VTAIL.t9 2.30819
R392 VTAIL.n178 VTAIL.n152 1.93989
R393 VTAIL.n190 VTAIL.n146 1.93989
R394 VTAIL.n34 VTAIL.n8 1.93989
R395 VTAIL.n46 VTAIL.n2 1.93989
R396 VTAIL.n144 VTAIL.n100 1.93989
R397 VTAIL.n132 VTAIL.n106 1.93989
R398 VTAIL.n96 VTAIL.n52 1.93989
R399 VTAIL.n84 VTAIL.n58 1.93989
R400 VTAIL.n179 VTAIL.n150 1.16414
R401 VTAIL.n188 VTAIL.n187 1.16414
R402 VTAIL.n35 VTAIL.n6 1.16414
R403 VTAIL.n44 VTAIL.n43 1.16414
R404 VTAIL.n142 VTAIL.n141 1.16414
R405 VTAIL.n133 VTAIL.n104 1.16414
R406 VTAIL.n94 VTAIL.n93 1.16414
R407 VTAIL.n85 VTAIL.n56 1.16414
R408 VTAIL.n99 VTAIL.n97 0.888431
R409 VTAIL.n47 VTAIL.n1 0.888431
R410 VTAIL.n97 VTAIL.n51 0.836707
R411 VTAIL.n145 VTAIL.n99 0.836707
R412 VTAIL.n49 VTAIL.n47 0.836707
R413 VTAIL VTAIL.n191 0.569465
R414 VTAIL.n183 VTAIL.n182 0.388379
R415 VTAIL.n184 VTAIL.n148 0.388379
R416 VTAIL.n39 VTAIL.n38 0.388379
R417 VTAIL.n40 VTAIL.n4 0.388379
R418 VTAIL.n138 VTAIL.n102 0.388379
R419 VTAIL.n137 VTAIL.n136 0.388379
R420 VTAIL.n90 VTAIL.n54 0.388379
R421 VTAIL.n89 VTAIL.n88 0.388379
R422 VTAIL VTAIL.n1 0.267741
R423 VTAIL.n164 VTAIL.n163 0.155672
R424 VTAIL.n164 VTAIL.n155 0.155672
R425 VTAIL.n171 VTAIL.n155 0.155672
R426 VTAIL.n172 VTAIL.n171 0.155672
R427 VTAIL.n172 VTAIL.n151 0.155672
R428 VTAIL.n180 VTAIL.n151 0.155672
R429 VTAIL.n181 VTAIL.n180 0.155672
R430 VTAIL.n181 VTAIL.n147 0.155672
R431 VTAIL.n189 VTAIL.n147 0.155672
R432 VTAIL.n20 VTAIL.n19 0.155672
R433 VTAIL.n20 VTAIL.n11 0.155672
R434 VTAIL.n27 VTAIL.n11 0.155672
R435 VTAIL.n28 VTAIL.n27 0.155672
R436 VTAIL.n28 VTAIL.n7 0.155672
R437 VTAIL.n36 VTAIL.n7 0.155672
R438 VTAIL.n37 VTAIL.n36 0.155672
R439 VTAIL.n37 VTAIL.n3 0.155672
R440 VTAIL.n45 VTAIL.n3 0.155672
R441 VTAIL.n143 VTAIL.n101 0.155672
R442 VTAIL.n135 VTAIL.n101 0.155672
R443 VTAIL.n135 VTAIL.n134 0.155672
R444 VTAIL.n134 VTAIL.n105 0.155672
R445 VTAIL.n127 VTAIL.n105 0.155672
R446 VTAIL.n127 VTAIL.n126 0.155672
R447 VTAIL.n126 VTAIL.n110 0.155672
R448 VTAIL.n119 VTAIL.n110 0.155672
R449 VTAIL.n119 VTAIL.n118 0.155672
R450 VTAIL.n95 VTAIL.n53 0.155672
R451 VTAIL.n87 VTAIL.n53 0.155672
R452 VTAIL.n87 VTAIL.n86 0.155672
R453 VTAIL.n86 VTAIL.n57 0.155672
R454 VTAIL.n79 VTAIL.n57 0.155672
R455 VTAIL.n79 VTAIL.n78 0.155672
R456 VTAIL.n78 VTAIL.n62 0.155672
R457 VTAIL.n71 VTAIL.n62 0.155672
R458 VTAIL.n71 VTAIL.n70 0.155672
R459 B.n531 B.n530 585
R460 B.n532 B.n531 585
R461 B.n222 B.n76 585
R462 B.n221 B.n220 585
R463 B.n219 B.n218 585
R464 B.n217 B.n216 585
R465 B.n215 B.n214 585
R466 B.n213 B.n212 585
R467 B.n211 B.n210 585
R468 B.n209 B.n208 585
R469 B.n207 B.n206 585
R470 B.n205 B.n204 585
R471 B.n203 B.n202 585
R472 B.n201 B.n200 585
R473 B.n199 B.n198 585
R474 B.n197 B.n196 585
R475 B.n195 B.n194 585
R476 B.n193 B.n192 585
R477 B.n191 B.n190 585
R478 B.n189 B.n188 585
R479 B.n187 B.n186 585
R480 B.n185 B.n184 585
R481 B.n183 B.n182 585
R482 B.n181 B.n180 585
R483 B.n179 B.n178 585
R484 B.n177 B.n176 585
R485 B.n175 B.n174 585
R486 B.n173 B.n172 585
R487 B.n171 B.n170 585
R488 B.n169 B.n168 585
R489 B.n167 B.n166 585
R490 B.n165 B.n164 585
R491 B.n163 B.n162 585
R492 B.n160 B.n159 585
R493 B.n158 B.n157 585
R494 B.n156 B.n155 585
R495 B.n154 B.n153 585
R496 B.n152 B.n151 585
R497 B.n150 B.n149 585
R498 B.n148 B.n147 585
R499 B.n146 B.n145 585
R500 B.n144 B.n143 585
R501 B.n142 B.n141 585
R502 B.n140 B.n139 585
R503 B.n138 B.n137 585
R504 B.n136 B.n135 585
R505 B.n134 B.n133 585
R506 B.n132 B.n131 585
R507 B.n130 B.n129 585
R508 B.n128 B.n127 585
R509 B.n126 B.n125 585
R510 B.n124 B.n123 585
R511 B.n122 B.n121 585
R512 B.n120 B.n119 585
R513 B.n118 B.n117 585
R514 B.n116 B.n115 585
R515 B.n114 B.n113 585
R516 B.n112 B.n111 585
R517 B.n110 B.n109 585
R518 B.n108 B.n107 585
R519 B.n106 B.n105 585
R520 B.n104 B.n103 585
R521 B.n102 B.n101 585
R522 B.n100 B.n99 585
R523 B.n98 B.n97 585
R524 B.n96 B.n95 585
R525 B.n94 B.n93 585
R526 B.n92 B.n91 585
R527 B.n90 B.n89 585
R528 B.n88 B.n87 585
R529 B.n86 B.n85 585
R530 B.n84 B.n83 585
R531 B.n40 B.n39 585
R532 B.n535 B.n534 585
R533 B.n529 B.n77 585
R534 B.n77 B.n37 585
R535 B.n528 B.n36 585
R536 B.n539 B.n36 585
R537 B.n527 B.n35 585
R538 B.n540 B.n35 585
R539 B.n526 B.n34 585
R540 B.n541 B.n34 585
R541 B.n525 B.n524 585
R542 B.n524 B.n33 585
R543 B.n523 B.n29 585
R544 B.n547 B.n29 585
R545 B.n522 B.n28 585
R546 B.n548 B.n28 585
R547 B.n521 B.n27 585
R548 B.n549 B.n27 585
R549 B.n520 B.n519 585
R550 B.n519 B.n23 585
R551 B.n518 B.n22 585
R552 B.n555 B.n22 585
R553 B.n517 B.n21 585
R554 B.n556 B.n21 585
R555 B.n516 B.n20 585
R556 B.n557 B.n20 585
R557 B.n515 B.n514 585
R558 B.n514 B.n16 585
R559 B.n513 B.n15 585
R560 B.n563 B.n15 585
R561 B.n512 B.n14 585
R562 B.n564 B.n14 585
R563 B.n511 B.n13 585
R564 B.n565 B.n13 585
R565 B.n510 B.n509 585
R566 B.n509 B.n12 585
R567 B.n508 B.n507 585
R568 B.n508 B.n8 585
R569 B.n506 B.n7 585
R570 B.n572 B.n7 585
R571 B.n505 B.n6 585
R572 B.n573 B.n6 585
R573 B.n504 B.n5 585
R574 B.n574 B.n5 585
R575 B.n503 B.n502 585
R576 B.n502 B.n4 585
R577 B.n501 B.n223 585
R578 B.n501 B.n500 585
R579 B.n490 B.n224 585
R580 B.n493 B.n224 585
R581 B.n492 B.n491 585
R582 B.n494 B.n492 585
R583 B.n489 B.n229 585
R584 B.n229 B.n228 585
R585 B.n488 B.n487 585
R586 B.n487 B.n486 585
R587 B.n231 B.n230 585
R588 B.n232 B.n231 585
R589 B.n479 B.n478 585
R590 B.n480 B.n479 585
R591 B.n477 B.n236 585
R592 B.n240 B.n236 585
R593 B.n476 B.n475 585
R594 B.n475 B.n474 585
R595 B.n238 B.n237 585
R596 B.n239 B.n238 585
R597 B.n467 B.n466 585
R598 B.n468 B.n467 585
R599 B.n465 B.n245 585
R600 B.n245 B.n244 585
R601 B.n464 B.n463 585
R602 B.n463 B.n462 585
R603 B.n247 B.n246 585
R604 B.n455 B.n247 585
R605 B.n454 B.n453 585
R606 B.n456 B.n454 585
R607 B.n452 B.n252 585
R608 B.n252 B.n251 585
R609 B.n451 B.n450 585
R610 B.n450 B.n449 585
R611 B.n254 B.n253 585
R612 B.n255 B.n254 585
R613 B.n445 B.n444 585
R614 B.n258 B.n257 585
R615 B.n441 B.n440 585
R616 B.n442 B.n441 585
R617 B.n439 B.n294 585
R618 B.n438 B.n437 585
R619 B.n436 B.n435 585
R620 B.n434 B.n433 585
R621 B.n432 B.n431 585
R622 B.n430 B.n429 585
R623 B.n428 B.n427 585
R624 B.n426 B.n425 585
R625 B.n424 B.n423 585
R626 B.n422 B.n421 585
R627 B.n420 B.n419 585
R628 B.n418 B.n417 585
R629 B.n416 B.n415 585
R630 B.n414 B.n413 585
R631 B.n412 B.n411 585
R632 B.n410 B.n409 585
R633 B.n408 B.n407 585
R634 B.n406 B.n405 585
R635 B.n404 B.n403 585
R636 B.n402 B.n401 585
R637 B.n400 B.n399 585
R638 B.n398 B.n397 585
R639 B.n396 B.n395 585
R640 B.n394 B.n393 585
R641 B.n392 B.n391 585
R642 B.n390 B.n389 585
R643 B.n388 B.n387 585
R644 B.n386 B.n385 585
R645 B.n384 B.n383 585
R646 B.n381 B.n380 585
R647 B.n379 B.n378 585
R648 B.n377 B.n376 585
R649 B.n375 B.n374 585
R650 B.n373 B.n372 585
R651 B.n371 B.n370 585
R652 B.n369 B.n368 585
R653 B.n367 B.n366 585
R654 B.n365 B.n364 585
R655 B.n363 B.n362 585
R656 B.n361 B.n360 585
R657 B.n359 B.n358 585
R658 B.n357 B.n356 585
R659 B.n355 B.n354 585
R660 B.n353 B.n352 585
R661 B.n351 B.n350 585
R662 B.n349 B.n348 585
R663 B.n347 B.n346 585
R664 B.n345 B.n344 585
R665 B.n343 B.n342 585
R666 B.n341 B.n340 585
R667 B.n339 B.n338 585
R668 B.n337 B.n336 585
R669 B.n335 B.n334 585
R670 B.n333 B.n332 585
R671 B.n331 B.n330 585
R672 B.n329 B.n328 585
R673 B.n327 B.n326 585
R674 B.n325 B.n324 585
R675 B.n323 B.n322 585
R676 B.n321 B.n320 585
R677 B.n319 B.n318 585
R678 B.n317 B.n316 585
R679 B.n315 B.n314 585
R680 B.n313 B.n312 585
R681 B.n311 B.n310 585
R682 B.n309 B.n308 585
R683 B.n307 B.n306 585
R684 B.n305 B.n304 585
R685 B.n303 B.n302 585
R686 B.n301 B.n300 585
R687 B.n446 B.n256 585
R688 B.n256 B.n255 585
R689 B.n448 B.n447 585
R690 B.n449 B.n448 585
R691 B.n250 B.n249 585
R692 B.n251 B.n250 585
R693 B.n458 B.n457 585
R694 B.n457 B.n456 585
R695 B.n459 B.n248 585
R696 B.n455 B.n248 585
R697 B.n461 B.n460 585
R698 B.n462 B.n461 585
R699 B.n243 B.n242 585
R700 B.n244 B.n243 585
R701 B.n470 B.n469 585
R702 B.n469 B.n468 585
R703 B.n471 B.n241 585
R704 B.n241 B.n239 585
R705 B.n473 B.n472 585
R706 B.n474 B.n473 585
R707 B.n235 B.n234 585
R708 B.n240 B.n235 585
R709 B.n482 B.n481 585
R710 B.n481 B.n480 585
R711 B.n483 B.n233 585
R712 B.n233 B.n232 585
R713 B.n485 B.n484 585
R714 B.n486 B.n485 585
R715 B.n227 B.n226 585
R716 B.n228 B.n227 585
R717 B.n496 B.n495 585
R718 B.n495 B.n494 585
R719 B.n497 B.n225 585
R720 B.n493 B.n225 585
R721 B.n499 B.n498 585
R722 B.n500 B.n499 585
R723 B.n3 B.n0 585
R724 B.n4 B.n3 585
R725 B.n571 B.n1 585
R726 B.n572 B.n571 585
R727 B.n570 B.n569 585
R728 B.n570 B.n8 585
R729 B.n568 B.n9 585
R730 B.n12 B.n9 585
R731 B.n567 B.n566 585
R732 B.n566 B.n565 585
R733 B.n11 B.n10 585
R734 B.n564 B.n11 585
R735 B.n562 B.n561 585
R736 B.n563 B.n562 585
R737 B.n560 B.n17 585
R738 B.n17 B.n16 585
R739 B.n559 B.n558 585
R740 B.n558 B.n557 585
R741 B.n19 B.n18 585
R742 B.n556 B.n19 585
R743 B.n554 B.n553 585
R744 B.n555 B.n554 585
R745 B.n552 B.n24 585
R746 B.n24 B.n23 585
R747 B.n551 B.n550 585
R748 B.n550 B.n549 585
R749 B.n26 B.n25 585
R750 B.n548 B.n26 585
R751 B.n546 B.n545 585
R752 B.n547 B.n546 585
R753 B.n544 B.n30 585
R754 B.n33 B.n30 585
R755 B.n543 B.n542 585
R756 B.n542 B.n541 585
R757 B.n32 B.n31 585
R758 B.n540 B.n32 585
R759 B.n538 B.n537 585
R760 B.n539 B.n538 585
R761 B.n536 B.n38 585
R762 B.n38 B.n37 585
R763 B.n575 B.n574 585
R764 B.n573 B.n2 585
R765 B.n80 B.t6 526.862
R766 B.n78 B.t10 526.862
R767 B.n297 B.t17 526.862
R768 B.n295 B.t13 526.862
R769 B.n534 B.n38 478.086
R770 B.n531 B.n77 478.086
R771 B.n300 B.n254 478.086
R772 B.n444 B.n256 478.086
R773 B.n532 B.n75 256.663
R774 B.n532 B.n74 256.663
R775 B.n532 B.n73 256.663
R776 B.n532 B.n72 256.663
R777 B.n532 B.n71 256.663
R778 B.n532 B.n70 256.663
R779 B.n532 B.n69 256.663
R780 B.n532 B.n68 256.663
R781 B.n532 B.n67 256.663
R782 B.n532 B.n66 256.663
R783 B.n532 B.n65 256.663
R784 B.n532 B.n64 256.663
R785 B.n532 B.n63 256.663
R786 B.n532 B.n62 256.663
R787 B.n532 B.n61 256.663
R788 B.n532 B.n60 256.663
R789 B.n532 B.n59 256.663
R790 B.n532 B.n58 256.663
R791 B.n532 B.n57 256.663
R792 B.n532 B.n56 256.663
R793 B.n532 B.n55 256.663
R794 B.n532 B.n54 256.663
R795 B.n532 B.n53 256.663
R796 B.n532 B.n52 256.663
R797 B.n532 B.n51 256.663
R798 B.n532 B.n50 256.663
R799 B.n532 B.n49 256.663
R800 B.n532 B.n48 256.663
R801 B.n532 B.n47 256.663
R802 B.n532 B.n46 256.663
R803 B.n532 B.n45 256.663
R804 B.n532 B.n44 256.663
R805 B.n532 B.n43 256.663
R806 B.n532 B.n42 256.663
R807 B.n532 B.n41 256.663
R808 B.n533 B.n532 256.663
R809 B.n443 B.n442 256.663
R810 B.n442 B.n259 256.663
R811 B.n442 B.n260 256.663
R812 B.n442 B.n261 256.663
R813 B.n442 B.n262 256.663
R814 B.n442 B.n263 256.663
R815 B.n442 B.n264 256.663
R816 B.n442 B.n265 256.663
R817 B.n442 B.n266 256.663
R818 B.n442 B.n267 256.663
R819 B.n442 B.n268 256.663
R820 B.n442 B.n269 256.663
R821 B.n442 B.n270 256.663
R822 B.n442 B.n271 256.663
R823 B.n442 B.n272 256.663
R824 B.n442 B.n273 256.663
R825 B.n442 B.n274 256.663
R826 B.n442 B.n275 256.663
R827 B.n442 B.n276 256.663
R828 B.n442 B.n277 256.663
R829 B.n442 B.n278 256.663
R830 B.n442 B.n279 256.663
R831 B.n442 B.n280 256.663
R832 B.n442 B.n281 256.663
R833 B.n442 B.n282 256.663
R834 B.n442 B.n283 256.663
R835 B.n442 B.n284 256.663
R836 B.n442 B.n285 256.663
R837 B.n442 B.n286 256.663
R838 B.n442 B.n287 256.663
R839 B.n442 B.n288 256.663
R840 B.n442 B.n289 256.663
R841 B.n442 B.n290 256.663
R842 B.n442 B.n291 256.663
R843 B.n442 B.n292 256.663
R844 B.n442 B.n293 256.663
R845 B.n577 B.n576 256.663
R846 B.n78 B.t11 241.874
R847 B.n297 B.t19 241.874
R848 B.n80 B.t8 241.873
R849 B.n295 B.t16 241.873
R850 B.n79 B.t12 223.06
R851 B.n298 B.t18 223.06
R852 B.n81 B.t9 223.06
R853 B.n296 B.t15 223.06
R854 B.n83 B.n40 163.367
R855 B.n87 B.n86 163.367
R856 B.n91 B.n90 163.367
R857 B.n95 B.n94 163.367
R858 B.n99 B.n98 163.367
R859 B.n103 B.n102 163.367
R860 B.n107 B.n106 163.367
R861 B.n111 B.n110 163.367
R862 B.n115 B.n114 163.367
R863 B.n119 B.n118 163.367
R864 B.n123 B.n122 163.367
R865 B.n127 B.n126 163.367
R866 B.n131 B.n130 163.367
R867 B.n135 B.n134 163.367
R868 B.n139 B.n138 163.367
R869 B.n143 B.n142 163.367
R870 B.n147 B.n146 163.367
R871 B.n151 B.n150 163.367
R872 B.n155 B.n154 163.367
R873 B.n159 B.n158 163.367
R874 B.n164 B.n163 163.367
R875 B.n168 B.n167 163.367
R876 B.n172 B.n171 163.367
R877 B.n176 B.n175 163.367
R878 B.n180 B.n179 163.367
R879 B.n184 B.n183 163.367
R880 B.n188 B.n187 163.367
R881 B.n192 B.n191 163.367
R882 B.n196 B.n195 163.367
R883 B.n200 B.n199 163.367
R884 B.n204 B.n203 163.367
R885 B.n208 B.n207 163.367
R886 B.n212 B.n211 163.367
R887 B.n216 B.n215 163.367
R888 B.n220 B.n219 163.367
R889 B.n531 B.n76 163.367
R890 B.n450 B.n254 163.367
R891 B.n450 B.n252 163.367
R892 B.n454 B.n252 163.367
R893 B.n454 B.n247 163.367
R894 B.n463 B.n247 163.367
R895 B.n463 B.n245 163.367
R896 B.n467 B.n245 163.367
R897 B.n467 B.n238 163.367
R898 B.n475 B.n238 163.367
R899 B.n475 B.n236 163.367
R900 B.n479 B.n236 163.367
R901 B.n479 B.n231 163.367
R902 B.n487 B.n231 163.367
R903 B.n487 B.n229 163.367
R904 B.n492 B.n229 163.367
R905 B.n492 B.n224 163.367
R906 B.n501 B.n224 163.367
R907 B.n502 B.n501 163.367
R908 B.n502 B.n5 163.367
R909 B.n6 B.n5 163.367
R910 B.n7 B.n6 163.367
R911 B.n508 B.n7 163.367
R912 B.n509 B.n508 163.367
R913 B.n509 B.n13 163.367
R914 B.n14 B.n13 163.367
R915 B.n15 B.n14 163.367
R916 B.n514 B.n15 163.367
R917 B.n514 B.n20 163.367
R918 B.n21 B.n20 163.367
R919 B.n22 B.n21 163.367
R920 B.n519 B.n22 163.367
R921 B.n519 B.n27 163.367
R922 B.n28 B.n27 163.367
R923 B.n29 B.n28 163.367
R924 B.n524 B.n29 163.367
R925 B.n524 B.n34 163.367
R926 B.n35 B.n34 163.367
R927 B.n36 B.n35 163.367
R928 B.n77 B.n36 163.367
R929 B.n441 B.n258 163.367
R930 B.n441 B.n294 163.367
R931 B.n437 B.n436 163.367
R932 B.n433 B.n432 163.367
R933 B.n429 B.n428 163.367
R934 B.n425 B.n424 163.367
R935 B.n421 B.n420 163.367
R936 B.n417 B.n416 163.367
R937 B.n413 B.n412 163.367
R938 B.n409 B.n408 163.367
R939 B.n405 B.n404 163.367
R940 B.n401 B.n400 163.367
R941 B.n397 B.n396 163.367
R942 B.n393 B.n392 163.367
R943 B.n389 B.n388 163.367
R944 B.n385 B.n384 163.367
R945 B.n380 B.n379 163.367
R946 B.n376 B.n375 163.367
R947 B.n372 B.n371 163.367
R948 B.n368 B.n367 163.367
R949 B.n364 B.n363 163.367
R950 B.n360 B.n359 163.367
R951 B.n356 B.n355 163.367
R952 B.n352 B.n351 163.367
R953 B.n348 B.n347 163.367
R954 B.n344 B.n343 163.367
R955 B.n340 B.n339 163.367
R956 B.n336 B.n335 163.367
R957 B.n332 B.n331 163.367
R958 B.n328 B.n327 163.367
R959 B.n324 B.n323 163.367
R960 B.n320 B.n319 163.367
R961 B.n316 B.n315 163.367
R962 B.n312 B.n311 163.367
R963 B.n308 B.n307 163.367
R964 B.n304 B.n303 163.367
R965 B.n448 B.n256 163.367
R966 B.n448 B.n250 163.367
R967 B.n457 B.n250 163.367
R968 B.n457 B.n248 163.367
R969 B.n461 B.n248 163.367
R970 B.n461 B.n243 163.367
R971 B.n469 B.n243 163.367
R972 B.n469 B.n241 163.367
R973 B.n473 B.n241 163.367
R974 B.n473 B.n235 163.367
R975 B.n481 B.n235 163.367
R976 B.n481 B.n233 163.367
R977 B.n485 B.n233 163.367
R978 B.n485 B.n227 163.367
R979 B.n495 B.n227 163.367
R980 B.n495 B.n225 163.367
R981 B.n499 B.n225 163.367
R982 B.n499 B.n3 163.367
R983 B.n575 B.n3 163.367
R984 B.n571 B.n2 163.367
R985 B.n571 B.n570 163.367
R986 B.n570 B.n9 163.367
R987 B.n566 B.n9 163.367
R988 B.n566 B.n11 163.367
R989 B.n562 B.n11 163.367
R990 B.n562 B.n17 163.367
R991 B.n558 B.n17 163.367
R992 B.n558 B.n19 163.367
R993 B.n554 B.n19 163.367
R994 B.n554 B.n24 163.367
R995 B.n550 B.n24 163.367
R996 B.n550 B.n26 163.367
R997 B.n546 B.n26 163.367
R998 B.n546 B.n30 163.367
R999 B.n542 B.n30 163.367
R1000 B.n542 B.n32 163.367
R1001 B.n538 B.n32 163.367
R1002 B.n538 B.n38 163.367
R1003 B.n442 B.n255 99.2426
R1004 B.n532 B.n37 99.2426
R1005 B.n534 B.n533 71.676
R1006 B.n83 B.n41 71.676
R1007 B.n87 B.n42 71.676
R1008 B.n91 B.n43 71.676
R1009 B.n95 B.n44 71.676
R1010 B.n99 B.n45 71.676
R1011 B.n103 B.n46 71.676
R1012 B.n107 B.n47 71.676
R1013 B.n111 B.n48 71.676
R1014 B.n115 B.n49 71.676
R1015 B.n119 B.n50 71.676
R1016 B.n123 B.n51 71.676
R1017 B.n127 B.n52 71.676
R1018 B.n131 B.n53 71.676
R1019 B.n135 B.n54 71.676
R1020 B.n139 B.n55 71.676
R1021 B.n143 B.n56 71.676
R1022 B.n147 B.n57 71.676
R1023 B.n151 B.n58 71.676
R1024 B.n155 B.n59 71.676
R1025 B.n159 B.n60 71.676
R1026 B.n164 B.n61 71.676
R1027 B.n168 B.n62 71.676
R1028 B.n172 B.n63 71.676
R1029 B.n176 B.n64 71.676
R1030 B.n180 B.n65 71.676
R1031 B.n184 B.n66 71.676
R1032 B.n188 B.n67 71.676
R1033 B.n192 B.n68 71.676
R1034 B.n196 B.n69 71.676
R1035 B.n200 B.n70 71.676
R1036 B.n204 B.n71 71.676
R1037 B.n208 B.n72 71.676
R1038 B.n212 B.n73 71.676
R1039 B.n216 B.n74 71.676
R1040 B.n220 B.n75 71.676
R1041 B.n76 B.n75 71.676
R1042 B.n219 B.n74 71.676
R1043 B.n215 B.n73 71.676
R1044 B.n211 B.n72 71.676
R1045 B.n207 B.n71 71.676
R1046 B.n203 B.n70 71.676
R1047 B.n199 B.n69 71.676
R1048 B.n195 B.n68 71.676
R1049 B.n191 B.n67 71.676
R1050 B.n187 B.n66 71.676
R1051 B.n183 B.n65 71.676
R1052 B.n179 B.n64 71.676
R1053 B.n175 B.n63 71.676
R1054 B.n171 B.n62 71.676
R1055 B.n167 B.n61 71.676
R1056 B.n163 B.n60 71.676
R1057 B.n158 B.n59 71.676
R1058 B.n154 B.n58 71.676
R1059 B.n150 B.n57 71.676
R1060 B.n146 B.n56 71.676
R1061 B.n142 B.n55 71.676
R1062 B.n138 B.n54 71.676
R1063 B.n134 B.n53 71.676
R1064 B.n130 B.n52 71.676
R1065 B.n126 B.n51 71.676
R1066 B.n122 B.n50 71.676
R1067 B.n118 B.n49 71.676
R1068 B.n114 B.n48 71.676
R1069 B.n110 B.n47 71.676
R1070 B.n106 B.n46 71.676
R1071 B.n102 B.n45 71.676
R1072 B.n98 B.n44 71.676
R1073 B.n94 B.n43 71.676
R1074 B.n90 B.n42 71.676
R1075 B.n86 B.n41 71.676
R1076 B.n533 B.n40 71.676
R1077 B.n444 B.n443 71.676
R1078 B.n294 B.n259 71.676
R1079 B.n436 B.n260 71.676
R1080 B.n432 B.n261 71.676
R1081 B.n428 B.n262 71.676
R1082 B.n424 B.n263 71.676
R1083 B.n420 B.n264 71.676
R1084 B.n416 B.n265 71.676
R1085 B.n412 B.n266 71.676
R1086 B.n408 B.n267 71.676
R1087 B.n404 B.n268 71.676
R1088 B.n400 B.n269 71.676
R1089 B.n396 B.n270 71.676
R1090 B.n392 B.n271 71.676
R1091 B.n388 B.n272 71.676
R1092 B.n384 B.n273 71.676
R1093 B.n379 B.n274 71.676
R1094 B.n375 B.n275 71.676
R1095 B.n371 B.n276 71.676
R1096 B.n367 B.n277 71.676
R1097 B.n363 B.n278 71.676
R1098 B.n359 B.n279 71.676
R1099 B.n355 B.n280 71.676
R1100 B.n351 B.n281 71.676
R1101 B.n347 B.n282 71.676
R1102 B.n343 B.n283 71.676
R1103 B.n339 B.n284 71.676
R1104 B.n335 B.n285 71.676
R1105 B.n331 B.n286 71.676
R1106 B.n327 B.n287 71.676
R1107 B.n323 B.n288 71.676
R1108 B.n319 B.n289 71.676
R1109 B.n315 B.n290 71.676
R1110 B.n311 B.n291 71.676
R1111 B.n307 B.n292 71.676
R1112 B.n303 B.n293 71.676
R1113 B.n443 B.n258 71.676
R1114 B.n437 B.n259 71.676
R1115 B.n433 B.n260 71.676
R1116 B.n429 B.n261 71.676
R1117 B.n425 B.n262 71.676
R1118 B.n421 B.n263 71.676
R1119 B.n417 B.n264 71.676
R1120 B.n413 B.n265 71.676
R1121 B.n409 B.n266 71.676
R1122 B.n405 B.n267 71.676
R1123 B.n401 B.n268 71.676
R1124 B.n397 B.n269 71.676
R1125 B.n393 B.n270 71.676
R1126 B.n389 B.n271 71.676
R1127 B.n385 B.n272 71.676
R1128 B.n380 B.n273 71.676
R1129 B.n376 B.n274 71.676
R1130 B.n372 B.n275 71.676
R1131 B.n368 B.n276 71.676
R1132 B.n364 B.n277 71.676
R1133 B.n360 B.n278 71.676
R1134 B.n356 B.n279 71.676
R1135 B.n352 B.n280 71.676
R1136 B.n348 B.n281 71.676
R1137 B.n344 B.n282 71.676
R1138 B.n340 B.n283 71.676
R1139 B.n336 B.n284 71.676
R1140 B.n332 B.n285 71.676
R1141 B.n328 B.n286 71.676
R1142 B.n324 B.n287 71.676
R1143 B.n320 B.n288 71.676
R1144 B.n316 B.n289 71.676
R1145 B.n312 B.n290 71.676
R1146 B.n308 B.n291 71.676
R1147 B.n304 B.n292 71.676
R1148 B.n300 B.n293 71.676
R1149 B.n576 B.n575 71.676
R1150 B.n576 B.n2 71.676
R1151 B.n82 B.n81 59.5399
R1152 B.n161 B.n79 59.5399
R1153 B.n299 B.n298 59.5399
R1154 B.n382 B.n296 59.5399
R1155 B.n449 B.n255 53.9882
R1156 B.n449 B.n251 53.9882
R1157 B.n456 B.n251 53.9882
R1158 B.n456 B.n455 53.9882
R1159 B.n462 B.n244 53.9882
R1160 B.n468 B.n244 53.9882
R1161 B.n468 B.n239 53.9882
R1162 B.n474 B.n239 53.9882
R1163 B.n474 B.n240 53.9882
R1164 B.n480 B.n232 53.9882
R1165 B.n486 B.n232 53.9882
R1166 B.n494 B.n228 53.9882
R1167 B.n494 B.n493 53.9882
R1168 B.n500 B.n4 53.9882
R1169 B.n574 B.n4 53.9882
R1170 B.n574 B.n573 53.9882
R1171 B.n573 B.n572 53.9882
R1172 B.n572 B.n8 53.9882
R1173 B.n565 B.n12 53.9882
R1174 B.n565 B.n564 53.9882
R1175 B.n563 B.n16 53.9882
R1176 B.n557 B.n16 53.9882
R1177 B.n556 B.n555 53.9882
R1178 B.n555 B.n23 53.9882
R1179 B.n549 B.n23 53.9882
R1180 B.n549 B.n548 53.9882
R1181 B.n548 B.n547 53.9882
R1182 B.n541 B.n33 53.9882
R1183 B.n541 B.n540 53.9882
R1184 B.n540 B.n539 53.9882
R1185 B.n539 B.n37 53.9882
R1186 B.n240 B.t3 41.2852
R1187 B.t1 B.n556 41.2852
R1188 B.n455 B.t14 38.1095
R1189 B.n33 B.t7 38.1095
R1190 B.n486 B.t0 33.3459
R1191 B.t4 B.n563 33.3459
R1192 B.n446 B.n445 31.0639
R1193 B.n301 B.n253 31.0639
R1194 B.n530 B.n529 31.0639
R1195 B.n536 B.n535 31.0639
R1196 B.n500 B.t2 28.5822
R1197 B.t5 B.n8 28.5822
R1198 B.n493 B.t2 25.4065
R1199 B.n12 B.t5 25.4065
R1200 B.t0 B.n228 20.6429
R1201 B.n564 B.t4 20.6429
R1202 B.n81 B.n80 18.8126
R1203 B.n79 B.n78 18.8126
R1204 B.n298 B.n297 18.8126
R1205 B.n296 B.n295 18.8126
R1206 B B.n577 18.0485
R1207 B.n462 B.t14 15.8792
R1208 B.n547 B.t7 15.8792
R1209 B.n480 B.t3 12.7035
R1210 B.n557 B.t1 12.7035
R1211 B.n447 B.n446 10.6151
R1212 B.n447 B.n249 10.6151
R1213 B.n458 B.n249 10.6151
R1214 B.n459 B.n458 10.6151
R1215 B.n460 B.n459 10.6151
R1216 B.n460 B.n242 10.6151
R1217 B.n470 B.n242 10.6151
R1218 B.n471 B.n470 10.6151
R1219 B.n472 B.n471 10.6151
R1220 B.n472 B.n234 10.6151
R1221 B.n482 B.n234 10.6151
R1222 B.n483 B.n482 10.6151
R1223 B.n484 B.n483 10.6151
R1224 B.n484 B.n226 10.6151
R1225 B.n496 B.n226 10.6151
R1226 B.n497 B.n496 10.6151
R1227 B.n498 B.n497 10.6151
R1228 B.n498 B.n0 10.6151
R1229 B.n445 B.n257 10.6151
R1230 B.n440 B.n257 10.6151
R1231 B.n440 B.n439 10.6151
R1232 B.n439 B.n438 10.6151
R1233 B.n438 B.n435 10.6151
R1234 B.n435 B.n434 10.6151
R1235 B.n434 B.n431 10.6151
R1236 B.n431 B.n430 10.6151
R1237 B.n430 B.n427 10.6151
R1238 B.n427 B.n426 10.6151
R1239 B.n426 B.n423 10.6151
R1240 B.n423 B.n422 10.6151
R1241 B.n422 B.n419 10.6151
R1242 B.n419 B.n418 10.6151
R1243 B.n418 B.n415 10.6151
R1244 B.n415 B.n414 10.6151
R1245 B.n414 B.n411 10.6151
R1246 B.n411 B.n410 10.6151
R1247 B.n410 B.n407 10.6151
R1248 B.n407 B.n406 10.6151
R1249 B.n406 B.n403 10.6151
R1250 B.n403 B.n402 10.6151
R1251 B.n402 B.n399 10.6151
R1252 B.n399 B.n398 10.6151
R1253 B.n398 B.n395 10.6151
R1254 B.n395 B.n394 10.6151
R1255 B.n394 B.n391 10.6151
R1256 B.n391 B.n390 10.6151
R1257 B.n390 B.n387 10.6151
R1258 B.n387 B.n386 10.6151
R1259 B.n386 B.n383 10.6151
R1260 B.n381 B.n378 10.6151
R1261 B.n378 B.n377 10.6151
R1262 B.n377 B.n374 10.6151
R1263 B.n374 B.n373 10.6151
R1264 B.n373 B.n370 10.6151
R1265 B.n370 B.n369 10.6151
R1266 B.n369 B.n366 10.6151
R1267 B.n366 B.n365 10.6151
R1268 B.n362 B.n361 10.6151
R1269 B.n361 B.n358 10.6151
R1270 B.n358 B.n357 10.6151
R1271 B.n357 B.n354 10.6151
R1272 B.n354 B.n353 10.6151
R1273 B.n353 B.n350 10.6151
R1274 B.n350 B.n349 10.6151
R1275 B.n349 B.n346 10.6151
R1276 B.n346 B.n345 10.6151
R1277 B.n345 B.n342 10.6151
R1278 B.n342 B.n341 10.6151
R1279 B.n341 B.n338 10.6151
R1280 B.n338 B.n337 10.6151
R1281 B.n337 B.n334 10.6151
R1282 B.n334 B.n333 10.6151
R1283 B.n333 B.n330 10.6151
R1284 B.n330 B.n329 10.6151
R1285 B.n329 B.n326 10.6151
R1286 B.n326 B.n325 10.6151
R1287 B.n325 B.n322 10.6151
R1288 B.n322 B.n321 10.6151
R1289 B.n321 B.n318 10.6151
R1290 B.n318 B.n317 10.6151
R1291 B.n317 B.n314 10.6151
R1292 B.n314 B.n313 10.6151
R1293 B.n313 B.n310 10.6151
R1294 B.n310 B.n309 10.6151
R1295 B.n309 B.n306 10.6151
R1296 B.n306 B.n305 10.6151
R1297 B.n305 B.n302 10.6151
R1298 B.n302 B.n301 10.6151
R1299 B.n451 B.n253 10.6151
R1300 B.n452 B.n451 10.6151
R1301 B.n453 B.n452 10.6151
R1302 B.n453 B.n246 10.6151
R1303 B.n464 B.n246 10.6151
R1304 B.n465 B.n464 10.6151
R1305 B.n466 B.n465 10.6151
R1306 B.n466 B.n237 10.6151
R1307 B.n476 B.n237 10.6151
R1308 B.n477 B.n476 10.6151
R1309 B.n478 B.n477 10.6151
R1310 B.n478 B.n230 10.6151
R1311 B.n488 B.n230 10.6151
R1312 B.n489 B.n488 10.6151
R1313 B.n491 B.n489 10.6151
R1314 B.n491 B.n490 10.6151
R1315 B.n490 B.n223 10.6151
R1316 B.n503 B.n223 10.6151
R1317 B.n504 B.n503 10.6151
R1318 B.n505 B.n504 10.6151
R1319 B.n506 B.n505 10.6151
R1320 B.n507 B.n506 10.6151
R1321 B.n510 B.n507 10.6151
R1322 B.n511 B.n510 10.6151
R1323 B.n512 B.n511 10.6151
R1324 B.n513 B.n512 10.6151
R1325 B.n515 B.n513 10.6151
R1326 B.n516 B.n515 10.6151
R1327 B.n517 B.n516 10.6151
R1328 B.n518 B.n517 10.6151
R1329 B.n520 B.n518 10.6151
R1330 B.n521 B.n520 10.6151
R1331 B.n522 B.n521 10.6151
R1332 B.n523 B.n522 10.6151
R1333 B.n525 B.n523 10.6151
R1334 B.n526 B.n525 10.6151
R1335 B.n527 B.n526 10.6151
R1336 B.n528 B.n527 10.6151
R1337 B.n529 B.n528 10.6151
R1338 B.n569 B.n1 10.6151
R1339 B.n569 B.n568 10.6151
R1340 B.n568 B.n567 10.6151
R1341 B.n567 B.n10 10.6151
R1342 B.n561 B.n10 10.6151
R1343 B.n561 B.n560 10.6151
R1344 B.n560 B.n559 10.6151
R1345 B.n559 B.n18 10.6151
R1346 B.n553 B.n18 10.6151
R1347 B.n553 B.n552 10.6151
R1348 B.n552 B.n551 10.6151
R1349 B.n551 B.n25 10.6151
R1350 B.n545 B.n25 10.6151
R1351 B.n545 B.n544 10.6151
R1352 B.n544 B.n543 10.6151
R1353 B.n543 B.n31 10.6151
R1354 B.n537 B.n31 10.6151
R1355 B.n537 B.n536 10.6151
R1356 B.n535 B.n39 10.6151
R1357 B.n84 B.n39 10.6151
R1358 B.n85 B.n84 10.6151
R1359 B.n88 B.n85 10.6151
R1360 B.n89 B.n88 10.6151
R1361 B.n92 B.n89 10.6151
R1362 B.n93 B.n92 10.6151
R1363 B.n96 B.n93 10.6151
R1364 B.n97 B.n96 10.6151
R1365 B.n100 B.n97 10.6151
R1366 B.n101 B.n100 10.6151
R1367 B.n104 B.n101 10.6151
R1368 B.n105 B.n104 10.6151
R1369 B.n108 B.n105 10.6151
R1370 B.n109 B.n108 10.6151
R1371 B.n112 B.n109 10.6151
R1372 B.n113 B.n112 10.6151
R1373 B.n116 B.n113 10.6151
R1374 B.n117 B.n116 10.6151
R1375 B.n120 B.n117 10.6151
R1376 B.n121 B.n120 10.6151
R1377 B.n124 B.n121 10.6151
R1378 B.n125 B.n124 10.6151
R1379 B.n128 B.n125 10.6151
R1380 B.n129 B.n128 10.6151
R1381 B.n132 B.n129 10.6151
R1382 B.n133 B.n132 10.6151
R1383 B.n136 B.n133 10.6151
R1384 B.n137 B.n136 10.6151
R1385 B.n140 B.n137 10.6151
R1386 B.n141 B.n140 10.6151
R1387 B.n145 B.n144 10.6151
R1388 B.n148 B.n145 10.6151
R1389 B.n149 B.n148 10.6151
R1390 B.n152 B.n149 10.6151
R1391 B.n153 B.n152 10.6151
R1392 B.n156 B.n153 10.6151
R1393 B.n157 B.n156 10.6151
R1394 B.n160 B.n157 10.6151
R1395 B.n165 B.n162 10.6151
R1396 B.n166 B.n165 10.6151
R1397 B.n169 B.n166 10.6151
R1398 B.n170 B.n169 10.6151
R1399 B.n173 B.n170 10.6151
R1400 B.n174 B.n173 10.6151
R1401 B.n177 B.n174 10.6151
R1402 B.n178 B.n177 10.6151
R1403 B.n181 B.n178 10.6151
R1404 B.n182 B.n181 10.6151
R1405 B.n185 B.n182 10.6151
R1406 B.n186 B.n185 10.6151
R1407 B.n189 B.n186 10.6151
R1408 B.n190 B.n189 10.6151
R1409 B.n193 B.n190 10.6151
R1410 B.n194 B.n193 10.6151
R1411 B.n197 B.n194 10.6151
R1412 B.n198 B.n197 10.6151
R1413 B.n201 B.n198 10.6151
R1414 B.n202 B.n201 10.6151
R1415 B.n205 B.n202 10.6151
R1416 B.n206 B.n205 10.6151
R1417 B.n209 B.n206 10.6151
R1418 B.n210 B.n209 10.6151
R1419 B.n213 B.n210 10.6151
R1420 B.n214 B.n213 10.6151
R1421 B.n217 B.n214 10.6151
R1422 B.n218 B.n217 10.6151
R1423 B.n221 B.n218 10.6151
R1424 B.n222 B.n221 10.6151
R1425 B.n530 B.n222 10.6151
R1426 B.n577 B.n0 8.11757
R1427 B.n577 B.n1 8.11757
R1428 B.n382 B.n381 6.5566
R1429 B.n365 B.n299 6.5566
R1430 B.n144 B.n82 6.5566
R1431 B.n161 B.n160 6.5566
R1432 B.n383 B.n382 4.05904
R1433 B.n362 B.n299 4.05904
R1434 B.n141 B.n82 4.05904
R1435 B.n162 B.n161 4.05904
R1436 VP.n1 VP.t0 411.291
R1437 VP.n6 VP.t1 384.471
R1438 VP.n7 VP.t3 384.471
R1439 VP.n8 VP.t5 384.471
R1440 VP.n3 VP.t4 384.471
R1441 VP.n2 VP.t2 384.471
R1442 VP.n9 VP.n8 161.3
R1443 VP.n4 VP.n3 161.3
R1444 VP.n6 VP.n5 161.3
R1445 VP.n7 VP.n0 80.6037
R1446 VP.n7 VP.n6 48.2005
R1447 VP.n8 VP.n7 48.2005
R1448 VP.n3 VP.n2 48.2005
R1449 VP.n4 VP.n1 45.1367
R1450 VP.n5 VP.n4 38.5043
R1451 VP.n2 VP.n1 13.3799
R1452 VP.n5 VP.n0 0.285035
R1453 VP.n9 VP.n0 0.285035
R1454 VP VP.n9 0.0516364
R1455 VDD1.n40 VDD1.n0 289.615
R1456 VDD1.n85 VDD1.n45 289.615
R1457 VDD1.n41 VDD1.n40 185
R1458 VDD1.n39 VDD1.n38 185
R1459 VDD1.n37 VDD1.n3 185
R1460 VDD1.n7 VDD1.n4 185
R1461 VDD1.n32 VDD1.n31 185
R1462 VDD1.n30 VDD1.n29 185
R1463 VDD1.n9 VDD1.n8 185
R1464 VDD1.n24 VDD1.n23 185
R1465 VDD1.n22 VDD1.n21 185
R1466 VDD1.n13 VDD1.n12 185
R1467 VDD1.n16 VDD1.n15 185
R1468 VDD1.n60 VDD1.n59 185
R1469 VDD1.n57 VDD1.n56 185
R1470 VDD1.n66 VDD1.n65 185
R1471 VDD1.n68 VDD1.n67 185
R1472 VDD1.n53 VDD1.n52 185
R1473 VDD1.n74 VDD1.n73 185
R1474 VDD1.n77 VDD1.n76 185
R1475 VDD1.n75 VDD1.n49 185
R1476 VDD1.n82 VDD1.n48 185
R1477 VDD1.n84 VDD1.n83 185
R1478 VDD1.n86 VDD1.n85 185
R1479 VDD1.t5 VDD1.n14 149.524
R1480 VDD1.t4 VDD1.n58 149.524
R1481 VDD1.n40 VDD1.n39 104.615
R1482 VDD1.n39 VDD1.n3 104.615
R1483 VDD1.n7 VDD1.n3 104.615
R1484 VDD1.n31 VDD1.n7 104.615
R1485 VDD1.n31 VDD1.n30 104.615
R1486 VDD1.n30 VDD1.n8 104.615
R1487 VDD1.n23 VDD1.n8 104.615
R1488 VDD1.n23 VDD1.n22 104.615
R1489 VDD1.n22 VDD1.n12 104.615
R1490 VDD1.n15 VDD1.n12 104.615
R1491 VDD1.n59 VDD1.n56 104.615
R1492 VDD1.n66 VDD1.n56 104.615
R1493 VDD1.n67 VDD1.n66 104.615
R1494 VDD1.n67 VDD1.n52 104.615
R1495 VDD1.n74 VDD1.n52 104.615
R1496 VDD1.n76 VDD1.n74 104.615
R1497 VDD1.n76 VDD1.n75 104.615
R1498 VDD1.n75 VDD1.n48 104.615
R1499 VDD1.n84 VDD1.n48 104.615
R1500 VDD1.n85 VDD1.n84 104.615
R1501 VDD1.n91 VDD1.n90 64.7584
R1502 VDD1.n93 VDD1.n92 64.6046
R1503 VDD1.n15 VDD1.t5 52.3082
R1504 VDD1.n59 VDD1.t4 52.3082
R1505 VDD1 VDD1.n44 50.7131
R1506 VDD1.n91 VDD1.n89 50.5996
R1507 VDD1.n93 VDD1.n91 34.8306
R1508 VDD1.n38 VDD1.n37 13.1884
R1509 VDD1.n83 VDD1.n82 13.1884
R1510 VDD1.n41 VDD1.n2 12.8005
R1511 VDD1.n36 VDD1.n4 12.8005
R1512 VDD1.n81 VDD1.n49 12.8005
R1513 VDD1.n86 VDD1.n47 12.8005
R1514 VDD1.n42 VDD1.n0 12.0247
R1515 VDD1.n33 VDD1.n32 12.0247
R1516 VDD1.n78 VDD1.n77 12.0247
R1517 VDD1.n87 VDD1.n45 12.0247
R1518 VDD1.n29 VDD1.n6 11.249
R1519 VDD1.n73 VDD1.n51 11.249
R1520 VDD1.n28 VDD1.n9 10.4732
R1521 VDD1.n72 VDD1.n53 10.4732
R1522 VDD1.n16 VDD1.n14 10.2747
R1523 VDD1.n60 VDD1.n58 10.2747
R1524 VDD1.n25 VDD1.n24 9.69747
R1525 VDD1.n69 VDD1.n68 9.69747
R1526 VDD1.n44 VDD1.n43 9.45567
R1527 VDD1.n89 VDD1.n88 9.45567
R1528 VDD1.n18 VDD1.n17 9.3005
R1529 VDD1.n20 VDD1.n19 9.3005
R1530 VDD1.n11 VDD1.n10 9.3005
R1531 VDD1.n26 VDD1.n25 9.3005
R1532 VDD1.n28 VDD1.n27 9.3005
R1533 VDD1.n6 VDD1.n5 9.3005
R1534 VDD1.n34 VDD1.n33 9.3005
R1535 VDD1.n36 VDD1.n35 9.3005
R1536 VDD1.n43 VDD1.n42 9.3005
R1537 VDD1.n2 VDD1.n1 9.3005
R1538 VDD1.n88 VDD1.n87 9.3005
R1539 VDD1.n47 VDD1.n46 9.3005
R1540 VDD1.n62 VDD1.n61 9.3005
R1541 VDD1.n64 VDD1.n63 9.3005
R1542 VDD1.n55 VDD1.n54 9.3005
R1543 VDD1.n70 VDD1.n69 9.3005
R1544 VDD1.n72 VDD1.n71 9.3005
R1545 VDD1.n51 VDD1.n50 9.3005
R1546 VDD1.n79 VDD1.n78 9.3005
R1547 VDD1.n81 VDD1.n80 9.3005
R1548 VDD1.n21 VDD1.n11 8.92171
R1549 VDD1.n65 VDD1.n55 8.92171
R1550 VDD1.n20 VDD1.n13 8.14595
R1551 VDD1.n64 VDD1.n57 8.14595
R1552 VDD1.n17 VDD1.n16 7.3702
R1553 VDD1.n61 VDD1.n60 7.3702
R1554 VDD1.n17 VDD1.n13 5.81868
R1555 VDD1.n61 VDD1.n57 5.81868
R1556 VDD1.n21 VDD1.n20 5.04292
R1557 VDD1.n65 VDD1.n64 5.04292
R1558 VDD1.n24 VDD1.n11 4.26717
R1559 VDD1.n68 VDD1.n55 4.26717
R1560 VDD1.n25 VDD1.n9 3.49141
R1561 VDD1.n69 VDD1.n53 3.49141
R1562 VDD1.n62 VDD1.n58 2.84303
R1563 VDD1.n18 VDD1.n14 2.84303
R1564 VDD1.n29 VDD1.n28 2.71565
R1565 VDD1.n73 VDD1.n72 2.71565
R1566 VDD1.n92 VDD1.t3 2.30819
R1567 VDD1.n92 VDD1.t1 2.30819
R1568 VDD1.n90 VDD1.t2 2.30819
R1569 VDD1.n90 VDD1.t0 2.30819
R1570 VDD1.n44 VDD1.n0 1.93989
R1571 VDD1.n32 VDD1.n6 1.93989
R1572 VDD1.n77 VDD1.n51 1.93989
R1573 VDD1.n89 VDD1.n45 1.93989
R1574 VDD1.n42 VDD1.n41 1.16414
R1575 VDD1.n33 VDD1.n4 1.16414
R1576 VDD1.n78 VDD1.n49 1.16414
R1577 VDD1.n87 VDD1.n86 1.16414
R1578 VDD1.n38 VDD1.n2 0.388379
R1579 VDD1.n37 VDD1.n36 0.388379
R1580 VDD1.n82 VDD1.n81 0.388379
R1581 VDD1.n83 VDD1.n47 0.388379
R1582 VDD1.n43 VDD1.n1 0.155672
R1583 VDD1.n35 VDD1.n1 0.155672
R1584 VDD1.n35 VDD1.n34 0.155672
R1585 VDD1.n34 VDD1.n5 0.155672
R1586 VDD1.n27 VDD1.n5 0.155672
R1587 VDD1.n27 VDD1.n26 0.155672
R1588 VDD1.n26 VDD1.n10 0.155672
R1589 VDD1.n19 VDD1.n10 0.155672
R1590 VDD1.n19 VDD1.n18 0.155672
R1591 VDD1.n63 VDD1.n62 0.155672
R1592 VDD1.n63 VDD1.n54 0.155672
R1593 VDD1.n70 VDD1.n54 0.155672
R1594 VDD1.n71 VDD1.n70 0.155672
R1595 VDD1.n71 VDD1.n50 0.155672
R1596 VDD1.n79 VDD1.n50 0.155672
R1597 VDD1.n80 VDD1.n79 0.155672
R1598 VDD1.n80 VDD1.n46 0.155672
R1599 VDD1.n88 VDD1.n46 0.155672
R1600 VDD1 VDD1.n93 0.151362
C0 VDD2 VDD1 0.688699f
C1 VP VN 4.38233f
C2 VDD2 VN 3.05573f
C3 VDD1 VN 0.148449f
C4 VTAIL VP 2.87436f
C5 VTAIL VDD2 7.90334f
C6 VTAIL VDD1 7.86795f
C7 VTAIL VN 2.85988f
C8 VP VDD2 0.292426f
C9 VP VDD1 3.19631f
C10 VDD2 B 3.832656f
C11 VDD1 B 3.850971f
C12 VTAIL B 5.088089f
C13 VN B 7.18316f
C14 VP B 5.344308f
C15 VDD1.n0 B 0.031213f
C16 VDD1.n1 B 0.023806f
C17 VDD1.n2 B 0.012793f
C18 VDD1.n3 B 0.030237f
C19 VDD1.n4 B 0.013545f
C20 VDD1.n5 B 0.023806f
C21 VDD1.n6 B 0.012793f
C22 VDD1.n7 B 0.030237f
C23 VDD1.n8 B 0.030237f
C24 VDD1.n9 B 0.013545f
C25 VDD1.n10 B 0.023806f
C26 VDD1.n11 B 0.012793f
C27 VDD1.n12 B 0.030237f
C28 VDD1.n13 B 0.013545f
C29 VDD1.n14 B 0.140397f
C30 VDD1.t5 B 0.050637f
C31 VDD1.n15 B 0.022678f
C32 VDD1.n16 B 0.021375f
C33 VDD1.n17 B 0.012793f
C34 VDD1.n18 B 0.83884f
C35 VDD1.n19 B 0.023806f
C36 VDD1.n20 B 0.012793f
C37 VDD1.n21 B 0.013545f
C38 VDD1.n22 B 0.030237f
C39 VDD1.n23 B 0.030237f
C40 VDD1.n24 B 0.013545f
C41 VDD1.n25 B 0.012793f
C42 VDD1.n26 B 0.023806f
C43 VDD1.n27 B 0.023806f
C44 VDD1.n28 B 0.012793f
C45 VDD1.n29 B 0.013545f
C46 VDD1.n30 B 0.030237f
C47 VDD1.n31 B 0.030237f
C48 VDD1.n32 B 0.013545f
C49 VDD1.n33 B 0.012793f
C50 VDD1.n34 B 0.023806f
C51 VDD1.n35 B 0.023806f
C52 VDD1.n36 B 0.012793f
C53 VDD1.n37 B 0.013169f
C54 VDD1.n38 B 0.013169f
C55 VDD1.n39 B 0.030237f
C56 VDD1.n40 B 0.061481f
C57 VDD1.n41 B 0.013545f
C58 VDD1.n42 B 0.012793f
C59 VDD1.n43 B 0.056979f
C60 VDD1.n44 B 0.05182f
C61 VDD1.n45 B 0.031213f
C62 VDD1.n46 B 0.023806f
C63 VDD1.n47 B 0.012793f
C64 VDD1.n48 B 0.030237f
C65 VDD1.n49 B 0.013545f
C66 VDD1.n50 B 0.023806f
C67 VDD1.n51 B 0.012793f
C68 VDD1.n52 B 0.030237f
C69 VDD1.n53 B 0.013545f
C70 VDD1.n54 B 0.023806f
C71 VDD1.n55 B 0.012793f
C72 VDD1.n56 B 0.030237f
C73 VDD1.n57 B 0.013545f
C74 VDD1.n58 B 0.140397f
C75 VDD1.t4 B 0.050637f
C76 VDD1.n59 B 0.022678f
C77 VDD1.n60 B 0.021375f
C78 VDD1.n61 B 0.012793f
C79 VDD1.n62 B 0.83884f
C80 VDD1.n63 B 0.023806f
C81 VDD1.n64 B 0.012793f
C82 VDD1.n65 B 0.013545f
C83 VDD1.n66 B 0.030237f
C84 VDD1.n67 B 0.030237f
C85 VDD1.n68 B 0.013545f
C86 VDD1.n69 B 0.012793f
C87 VDD1.n70 B 0.023806f
C88 VDD1.n71 B 0.023806f
C89 VDD1.n72 B 0.012793f
C90 VDD1.n73 B 0.013545f
C91 VDD1.n74 B 0.030237f
C92 VDD1.n75 B 0.030237f
C93 VDD1.n76 B 0.030237f
C94 VDD1.n77 B 0.013545f
C95 VDD1.n78 B 0.012793f
C96 VDD1.n79 B 0.023806f
C97 VDD1.n80 B 0.023806f
C98 VDD1.n81 B 0.012793f
C99 VDD1.n82 B 0.013169f
C100 VDD1.n83 B 0.013169f
C101 VDD1.n84 B 0.030237f
C102 VDD1.n85 B 0.061481f
C103 VDD1.n86 B 0.013545f
C104 VDD1.n87 B 0.012793f
C105 VDD1.n88 B 0.056979f
C106 VDD1.n89 B 0.051512f
C107 VDD1.t2 B 0.161412f
C108 VDD1.t0 B 0.161412f
C109 VDD1.n90 B 1.40643f
C110 VDD1.n91 B 1.61041f
C111 VDD1.t3 B 0.161412f
C112 VDD1.t1 B 0.161412f
C113 VDD1.n92 B 1.40577f
C114 VDD1.n93 B 1.86846f
C115 VP.n0 B 0.065274f
C116 VP.t0 B 0.79453f
C117 VP.n1 B 0.309337f
C118 VP.t4 B 0.773016f
C119 VP.t2 B 0.773016f
C120 VP.n2 B 0.340898f
C121 VP.n3 B 0.329772f
C122 VP.n4 B 1.90648f
C123 VP.n5 B 1.80523f
C124 VP.t1 B 0.773016f
C125 VP.n6 B 0.329772f
C126 VP.t3 B 0.773016f
C127 VP.n7 B 0.340898f
C128 VP.t5 B 0.773016f
C129 VP.n8 B 0.329772f
C130 VP.n9 B 0.054393f
C131 VTAIL.t8 B 0.171763f
C132 VTAIL.t4 B 0.171763f
C133 VTAIL.n0 B 1.42698f
C134 VTAIL.n1 B 0.331691f
C135 VTAIL.n2 B 0.033215f
C136 VTAIL.n3 B 0.025333f
C137 VTAIL.n4 B 0.013613f
C138 VTAIL.n5 B 0.032176f
C139 VTAIL.n6 B 0.014414f
C140 VTAIL.n7 B 0.025333f
C141 VTAIL.n8 B 0.013613f
C142 VTAIL.n9 B 0.032176f
C143 VTAIL.n10 B 0.014414f
C144 VTAIL.n11 B 0.025333f
C145 VTAIL.n12 B 0.013613f
C146 VTAIL.n13 B 0.032176f
C147 VTAIL.n14 B 0.014414f
C148 VTAIL.n15 B 0.1494f
C149 VTAIL.t2 B 0.053884f
C150 VTAIL.n16 B 0.024132f
C151 VTAIL.n17 B 0.022746f
C152 VTAIL.n18 B 0.013613f
C153 VTAIL.n19 B 0.89263f
C154 VTAIL.n20 B 0.025333f
C155 VTAIL.n21 B 0.013613f
C156 VTAIL.n22 B 0.014414f
C157 VTAIL.n23 B 0.032176f
C158 VTAIL.n24 B 0.032176f
C159 VTAIL.n25 B 0.014414f
C160 VTAIL.n26 B 0.013613f
C161 VTAIL.n27 B 0.025333f
C162 VTAIL.n28 B 0.025333f
C163 VTAIL.n29 B 0.013613f
C164 VTAIL.n30 B 0.014414f
C165 VTAIL.n31 B 0.032176f
C166 VTAIL.n32 B 0.032176f
C167 VTAIL.n33 B 0.032176f
C168 VTAIL.n34 B 0.014414f
C169 VTAIL.n35 B 0.013613f
C170 VTAIL.n36 B 0.025333f
C171 VTAIL.n37 B 0.025333f
C172 VTAIL.n38 B 0.013613f
C173 VTAIL.n39 B 0.014013f
C174 VTAIL.n40 B 0.014013f
C175 VTAIL.n41 B 0.032176f
C176 VTAIL.n42 B 0.065424f
C177 VTAIL.n43 B 0.014414f
C178 VTAIL.n44 B 0.013613f
C179 VTAIL.n45 B 0.060633f
C180 VTAIL.n46 B 0.036235f
C181 VTAIL.n47 B 0.163549f
C182 VTAIL.t3 B 0.171763f
C183 VTAIL.t0 B 0.171763f
C184 VTAIL.n48 B 1.42698f
C185 VTAIL.n49 B 1.39006f
C186 VTAIL.t7 B 0.171763f
C187 VTAIL.t9 B 0.171763f
C188 VTAIL.n50 B 1.42699f
C189 VTAIL.n51 B 1.39005f
C190 VTAIL.n52 B 0.033215f
C191 VTAIL.n53 B 0.025333f
C192 VTAIL.n54 B 0.013613f
C193 VTAIL.n55 B 0.032176f
C194 VTAIL.n56 B 0.014414f
C195 VTAIL.n57 B 0.025333f
C196 VTAIL.n58 B 0.013613f
C197 VTAIL.n59 B 0.032176f
C198 VTAIL.n60 B 0.032176f
C199 VTAIL.n61 B 0.014414f
C200 VTAIL.n62 B 0.025333f
C201 VTAIL.n63 B 0.013613f
C202 VTAIL.n64 B 0.032176f
C203 VTAIL.n65 B 0.014414f
C204 VTAIL.n66 B 0.1494f
C205 VTAIL.t5 B 0.053884f
C206 VTAIL.n67 B 0.024132f
C207 VTAIL.n68 B 0.022746f
C208 VTAIL.n69 B 0.013613f
C209 VTAIL.n70 B 0.89263f
C210 VTAIL.n71 B 0.025333f
C211 VTAIL.n72 B 0.013613f
C212 VTAIL.n73 B 0.014414f
C213 VTAIL.n74 B 0.032176f
C214 VTAIL.n75 B 0.032176f
C215 VTAIL.n76 B 0.014414f
C216 VTAIL.n77 B 0.013613f
C217 VTAIL.n78 B 0.025333f
C218 VTAIL.n79 B 0.025333f
C219 VTAIL.n80 B 0.013613f
C220 VTAIL.n81 B 0.014414f
C221 VTAIL.n82 B 0.032176f
C222 VTAIL.n83 B 0.032176f
C223 VTAIL.n84 B 0.014414f
C224 VTAIL.n85 B 0.013613f
C225 VTAIL.n86 B 0.025333f
C226 VTAIL.n87 B 0.025333f
C227 VTAIL.n88 B 0.013613f
C228 VTAIL.n89 B 0.014013f
C229 VTAIL.n90 B 0.014013f
C230 VTAIL.n91 B 0.032176f
C231 VTAIL.n92 B 0.065424f
C232 VTAIL.n93 B 0.014414f
C233 VTAIL.n94 B 0.013613f
C234 VTAIL.n95 B 0.060633f
C235 VTAIL.n96 B 0.036235f
C236 VTAIL.n97 B 0.163549f
C237 VTAIL.t10 B 0.171763f
C238 VTAIL.t11 B 0.171763f
C239 VTAIL.n98 B 1.42699f
C240 VTAIL.n99 B 0.378126f
C241 VTAIL.n100 B 0.033215f
C242 VTAIL.n101 B 0.025333f
C243 VTAIL.n102 B 0.013613f
C244 VTAIL.n103 B 0.032176f
C245 VTAIL.n104 B 0.014414f
C246 VTAIL.n105 B 0.025333f
C247 VTAIL.n106 B 0.013613f
C248 VTAIL.n107 B 0.032176f
C249 VTAIL.n108 B 0.032176f
C250 VTAIL.n109 B 0.014414f
C251 VTAIL.n110 B 0.025333f
C252 VTAIL.n111 B 0.013613f
C253 VTAIL.n112 B 0.032176f
C254 VTAIL.n113 B 0.014414f
C255 VTAIL.n114 B 0.1494f
C256 VTAIL.t1 B 0.053884f
C257 VTAIL.n115 B 0.024132f
C258 VTAIL.n116 B 0.022746f
C259 VTAIL.n117 B 0.013613f
C260 VTAIL.n118 B 0.89263f
C261 VTAIL.n119 B 0.025333f
C262 VTAIL.n120 B 0.013613f
C263 VTAIL.n121 B 0.014414f
C264 VTAIL.n122 B 0.032176f
C265 VTAIL.n123 B 0.032176f
C266 VTAIL.n124 B 0.014414f
C267 VTAIL.n125 B 0.013613f
C268 VTAIL.n126 B 0.025333f
C269 VTAIL.n127 B 0.025333f
C270 VTAIL.n128 B 0.013613f
C271 VTAIL.n129 B 0.014414f
C272 VTAIL.n130 B 0.032176f
C273 VTAIL.n131 B 0.032176f
C274 VTAIL.n132 B 0.014414f
C275 VTAIL.n133 B 0.013613f
C276 VTAIL.n134 B 0.025333f
C277 VTAIL.n135 B 0.025333f
C278 VTAIL.n136 B 0.013613f
C279 VTAIL.n137 B 0.014013f
C280 VTAIL.n138 B 0.014013f
C281 VTAIL.n139 B 0.032176f
C282 VTAIL.n140 B 0.065424f
C283 VTAIL.n141 B 0.014414f
C284 VTAIL.n142 B 0.013613f
C285 VTAIL.n143 B 0.060633f
C286 VTAIL.n144 B 0.036235f
C287 VTAIL.n145 B 1.10722f
C288 VTAIL.n146 B 0.033215f
C289 VTAIL.n147 B 0.025333f
C290 VTAIL.n148 B 0.013613f
C291 VTAIL.n149 B 0.032176f
C292 VTAIL.n150 B 0.014414f
C293 VTAIL.n151 B 0.025333f
C294 VTAIL.n152 B 0.013613f
C295 VTAIL.n153 B 0.032176f
C296 VTAIL.n154 B 0.014414f
C297 VTAIL.n155 B 0.025333f
C298 VTAIL.n156 B 0.013613f
C299 VTAIL.n157 B 0.032176f
C300 VTAIL.n158 B 0.014414f
C301 VTAIL.n159 B 0.1494f
C302 VTAIL.t6 B 0.053884f
C303 VTAIL.n160 B 0.024132f
C304 VTAIL.n161 B 0.022746f
C305 VTAIL.n162 B 0.013613f
C306 VTAIL.n163 B 0.89263f
C307 VTAIL.n164 B 0.025333f
C308 VTAIL.n165 B 0.013613f
C309 VTAIL.n166 B 0.014414f
C310 VTAIL.n167 B 0.032176f
C311 VTAIL.n168 B 0.032176f
C312 VTAIL.n169 B 0.014414f
C313 VTAIL.n170 B 0.013613f
C314 VTAIL.n171 B 0.025333f
C315 VTAIL.n172 B 0.025333f
C316 VTAIL.n173 B 0.013613f
C317 VTAIL.n174 B 0.014414f
C318 VTAIL.n175 B 0.032176f
C319 VTAIL.n176 B 0.032176f
C320 VTAIL.n177 B 0.032176f
C321 VTAIL.n178 B 0.014414f
C322 VTAIL.n179 B 0.013613f
C323 VTAIL.n180 B 0.025333f
C324 VTAIL.n181 B 0.025333f
C325 VTAIL.n182 B 0.013613f
C326 VTAIL.n183 B 0.014013f
C327 VTAIL.n184 B 0.014013f
C328 VTAIL.n185 B 0.032176f
C329 VTAIL.n186 B 0.065424f
C330 VTAIL.n187 B 0.014414f
C331 VTAIL.n188 B 0.013613f
C332 VTAIL.n189 B 0.060633f
C333 VTAIL.n190 B 0.036235f
C334 VTAIL.n191 B 1.0854f
C335 VDD2.n0 B 0.031179f
C336 VDD2.n1 B 0.02378f
C337 VDD2.n2 B 0.012779f
C338 VDD2.n3 B 0.030204f
C339 VDD2.n4 B 0.01353f
C340 VDD2.n5 B 0.02378f
C341 VDD2.n6 B 0.012779f
C342 VDD2.n7 B 0.030204f
C343 VDD2.n8 B 0.01353f
C344 VDD2.n9 B 0.02378f
C345 VDD2.n10 B 0.012779f
C346 VDD2.n11 B 0.030204f
C347 VDD2.n12 B 0.01353f
C348 VDD2.n13 B 0.140243f
C349 VDD2.t5 B 0.050582f
C350 VDD2.n14 B 0.022653f
C351 VDD2.n15 B 0.021352f
C352 VDD2.n16 B 0.012779f
C353 VDD2.n17 B 0.83792f
C354 VDD2.n18 B 0.02378f
C355 VDD2.n19 B 0.012779f
C356 VDD2.n20 B 0.01353f
C357 VDD2.n21 B 0.030204f
C358 VDD2.n22 B 0.030204f
C359 VDD2.n23 B 0.01353f
C360 VDD2.n24 B 0.012779f
C361 VDD2.n25 B 0.02378f
C362 VDD2.n26 B 0.02378f
C363 VDD2.n27 B 0.012779f
C364 VDD2.n28 B 0.01353f
C365 VDD2.n29 B 0.030204f
C366 VDD2.n30 B 0.030204f
C367 VDD2.n31 B 0.030204f
C368 VDD2.n32 B 0.01353f
C369 VDD2.n33 B 0.012779f
C370 VDD2.n34 B 0.02378f
C371 VDD2.n35 B 0.02378f
C372 VDD2.n36 B 0.012779f
C373 VDD2.n37 B 0.013154f
C374 VDD2.n38 B 0.013154f
C375 VDD2.n39 B 0.030204f
C376 VDD2.n40 B 0.061414f
C377 VDD2.n41 B 0.01353f
C378 VDD2.n42 B 0.012779f
C379 VDD2.n43 B 0.056916f
C380 VDD2.n44 B 0.051455f
C381 VDD2.t1 B 0.161235f
C382 VDD2.t2 B 0.161235f
C383 VDD2.n45 B 1.40489f
C384 VDD2.n46 B 1.53776f
C385 VDD2.n47 B 0.031179f
C386 VDD2.n48 B 0.02378f
C387 VDD2.n49 B 0.012779f
C388 VDD2.n50 B 0.030204f
C389 VDD2.n51 B 0.01353f
C390 VDD2.n52 B 0.02378f
C391 VDD2.n53 B 0.012779f
C392 VDD2.n54 B 0.030204f
C393 VDD2.n55 B 0.030204f
C394 VDD2.n56 B 0.01353f
C395 VDD2.n57 B 0.02378f
C396 VDD2.n58 B 0.012779f
C397 VDD2.n59 B 0.030204f
C398 VDD2.n60 B 0.01353f
C399 VDD2.n61 B 0.140243f
C400 VDD2.t3 B 0.050582f
C401 VDD2.n62 B 0.022653f
C402 VDD2.n63 B 0.021352f
C403 VDD2.n64 B 0.012779f
C404 VDD2.n65 B 0.83792f
C405 VDD2.n66 B 0.02378f
C406 VDD2.n67 B 0.012779f
C407 VDD2.n68 B 0.01353f
C408 VDD2.n69 B 0.030204f
C409 VDD2.n70 B 0.030204f
C410 VDD2.n71 B 0.01353f
C411 VDD2.n72 B 0.012779f
C412 VDD2.n73 B 0.02378f
C413 VDD2.n74 B 0.02378f
C414 VDD2.n75 B 0.012779f
C415 VDD2.n76 B 0.01353f
C416 VDD2.n77 B 0.030204f
C417 VDD2.n78 B 0.030204f
C418 VDD2.n79 B 0.01353f
C419 VDD2.n80 B 0.012779f
C420 VDD2.n81 B 0.02378f
C421 VDD2.n82 B 0.02378f
C422 VDD2.n83 B 0.012779f
C423 VDD2.n84 B 0.013154f
C424 VDD2.n85 B 0.013154f
C425 VDD2.n86 B 0.030204f
C426 VDD2.n87 B 0.061414f
C427 VDD2.n88 B 0.01353f
C428 VDD2.n89 B 0.012779f
C429 VDD2.n90 B 0.056916f
C430 VDD2.n91 B 0.050419f
C431 VDD2.n92 B 1.67321f
C432 VDD2.t4 B 0.161235f
C433 VDD2.t0 B 0.161235f
C434 VDD2.n93 B 1.40487f
C435 VN.t1 B 0.781831f
C436 VN.n0 B 0.304393f
C437 VN.t5 B 0.76066f
C438 VN.n1 B 0.335449f
C439 VN.t3 B 0.76066f
C440 VN.n2 B 0.324501f
C441 VN.n3 B 0.198326f
C442 VN.t4 B 0.781831f
C443 VN.n4 B 0.304393f
C444 VN.t0 B 0.76066f
C445 VN.n5 B 0.335449f
C446 VN.t2 B 0.76066f
C447 VN.n6 B 0.324501f
C448 VN.n7 B 1.90786f
.ends

