* NGSPICE file created from diff_pair_sample_1500.ext - technology: sky130A

.subckt diff_pair_sample_1500 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 w_n1494_n4352# sky130_fd_pr__pfet_01v8 ad=6.591 pd=34.58 as=6.591 ps=34.58 w=16.9 l=0.98
X1 VDD2.t1 VN.t0 VTAIL.t0 w_n1494_n4352# sky130_fd_pr__pfet_01v8 ad=6.591 pd=34.58 as=6.591 ps=34.58 w=16.9 l=0.98
X2 B.t11 B.t9 B.t10 w_n1494_n4352# sky130_fd_pr__pfet_01v8 ad=6.591 pd=34.58 as=0 ps=0 w=16.9 l=0.98
X3 B.t8 B.t6 B.t7 w_n1494_n4352# sky130_fd_pr__pfet_01v8 ad=6.591 pd=34.58 as=0 ps=0 w=16.9 l=0.98
X4 VDD2.t0 VN.t1 VTAIL.t1 w_n1494_n4352# sky130_fd_pr__pfet_01v8 ad=6.591 pd=34.58 as=6.591 ps=34.58 w=16.9 l=0.98
X5 B.t5 B.t3 B.t4 w_n1494_n4352# sky130_fd_pr__pfet_01v8 ad=6.591 pd=34.58 as=0 ps=0 w=16.9 l=0.98
X6 VDD1.t0 VP.t1 VTAIL.t3 w_n1494_n4352# sky130_fd_pr__pfet_01v8 ad=6.591 pd=34.58 as=6.591 ps=34.58 w=16.9 l=0.98
X7 B.t2 B.t0 B.t1 w_n1494_n4352# sky130_fd_pr__pfet_01v8 ad=6.591 pd=34.58 as=0 ps=0 w=16.9 l=0.98
R0 VP.n0 VP.t0 661.074
R1 VP.n0 VP.t1 616.987
R2 VP VP.n0 0.0516364
R3 VTAIL.n370 VTAIL.n282 756.745
R4 VTAIL.n88 VTAIL.n0 756.745
R5 VTAIL.n276 VTAIL.n188 756.745
R6 VTAIL.n182 VTAIL.n94 756.745
R7 VTAIL.n313 VTAIL.n312 585
R8 VTAIL.n310 VTAIL.n309 585
R9 VTAIL.n319 VTAIL.n318 585
R10 VTAIL.n321 VTAIL.n320 585
R11 VTAIL.n306 VTAIL.n305 585
R12 VTAIL.n327 VTAIL.n326 585
R13 VTAIL.n329 VTAIL.n328 585
R14 VTAIL.n302 VTAIL.n301 585
R15 VTAIL.n335 VTAIL.n334 585
R16 VTAIL.n337 VTAIL.n336 585
R17 VTAIL.n298 VTAIL.n297 585
R18 VTAIL.n343 VTAIL.n342 585
R19 VTAIL.n345 VTAIL.n344 585
R20 VTAIL.n294 VTAIL.n293 585
R21 VTAIL.n351 VTAIL.n350 585
R22 VTAIL.n354 VTAIL.n353 585
R23 VTAIL.n352 VTAIL.n290 585
R24 VTAIL.n359 VTAIL.n289 585
R25 VTAIL.n361 VTAIL.n360 585
R26 VTAIL.n363 VTAIL.n362 585
R27 VTAIL.n286 VTAIL.n285 585
R28 VTAIL.n369 VTAIL.n368 585
R29 VTAIL.n371 VTAIL.n370 585
R30 VTAIL.n31 VTAIL.n30 585
R31 VTAIL.n28 VTAIL.n27 585
R32 VTAIL.n37 VTAIL.n36 585
R33 VTAIL.n39 VTAIL.n38 585
R34 VTAIL.n24 VTAIL.n23 585
R35 VTAIL.n45 VTAIL.n44 585
R36 VTAIL.n47 VTAIL.n46 585
R37 VTAIL.n20 VTAIL.n19 585
R38 VTAIL.n53 VTAIL.n52 585
R39 VTAIL.n55 VTAIL.n54 585
R40 VTAIL.n16 VTAIL.n15 585
R41 VTAIL.n61 VTAIL.n60 585
R42 VTAIL.n63 VTAIL.n62 585
R43 VTAIL.n12 VTAIL.n11 585
R44 VTAIL.n69 VTAIL.n68 585
R45 VTAIL.n72 VTAIL.n71 585
R46 VTAIL.n70 VTAIL.n8 585
R47 VTAIL.n77 VTAIL.n7 585
R48 VTAIL.n79 VTAIL.n78 585
R49 VTAIL.n81 VTAIL.n80 585
R50 VTAIL.n4 VTAIL.n3 585
R51 VTAIL.n87 VTAIL.n86 585
R52 VTAIL.n89 VTAIL.n88 585
R53 VTAIL.n277 VTAIL.n276 585
R54 VTAIL.n275 VTAIL.n274 585
R55 VTAIL.n192 VTAIL.n191 585
R56 VTAIL.n269 VTAIL.n268 585
R57 VTAIL.n267 VTAIL.n266 585
R58 VTAIL.n265 VTAIL.n195 585
R59 VTAIL.n199 VTAIL.n196 585
R60 VTAIL.n260 VTAIL.n259 585
R61 VTAIL.n258 VTAIL.n257 585
R62 VTAIL.n201 VTAIL.n200 585
R63 VTAIL.n252 VTAIL.n251 585
R64 VTAIL.n250 VTAIL.n249 585
R65 VTAIL.n205 VTAIL.n204 585
R66 VTAIL.n244 VTAIL.n243 585
R67 VTAIL.n242 VTAIL.n241 585
R68 VTAIL.n209 VTAIL.n208 585
R69 VTAIL.n236 VTAIL.n235 585
R70 VTAIL.n234 VTAIL.n233 585
R71 VTAIL.n213 VTAIL.n212 585
R72 VTAIL.n228 VTAIL.n227 585
R73 VTAIL.n226 VTAIL.n225 585
R74 VTAIL.n217 VTAIL.n216 585
R75 VTAIL.n220 VTAIL.n219 585
R76 VTAIL.n183 VTAIL.n182 585
R77 VTAIL.n181 VTAIL.n180 585
R78 VTAIL.n98 VTAIL.n97 585
R79 VTAIL.n175 VTAIL.n174 585
R80 VTAIL.n173 VTAIL.n172 585
R81 VTAIL.n171 VTAIL.n101 585
R82 VTAIL.n105 VTAIL.n102 585
R83 VTAIL.n166 VTAIL.n165 585
R84 VTAIL.n164 VTAIL.n163 585
R85 VTAIL.n107 VTAIL.n106 585
R86 VTAIL.n158 VTAIL.n157 585
R87 VTAIL.n156 VTAIL.n155 585
R88 VTAIL.n111 VTAIL.n110 585
R89 VTAIL.n150 VTAIL.n149 585
R90 VTAIL.n148 VTAIL.n147 585
R91 VTAIL.n115 VTAIL.n114 585
R92 VTAIL.n142 VTAIL.n141 585
R93 VTAIL.n140 VTAIL.n139 585
R94 VTAIL.n119 VTAIL.n118 585
R95 VTAIL.n134 VTAIL.n133 585
R96 VTAIL.n132 VTAIL.n131 585
R97 VTAIL.n123 VTAIL.n122 585
R98 VTAIL.n126 VTAIL.n125 585
R99 VTAIL.t2 VTAIL.n218 327.466
R100 VTAIL.t1 VTAIL.n124 327.466
R101 VTAIL.t0 VTAIL.n311 327.466
R102 VTAIL.t3 VTAIL.n29 327.466
R103 VTAIL.n312 VTAIL.n309 171.744
R104 VTAIL.n319 VTAIL.n309 171.744
R105 VTAIL.n320 VTAIL.n319 171.744
R106 VTAIL.n320 VTAIL.n305 171.744
R107 VTAIL.n327 VTAIL.n305 171.744
R108 VTAIL.n328 VTAIL.n327 171.744
R109 VTAIL.n328 VTAIL.n301 171.744
R110 VTAIL.n335 VTAIL.n301 171.744
R111 VTAIL.n336 VTAIL.n335 171.744
R112 VTAIL.n336 VTAIL.n297 171.744
R113 VTAIL.n343 VTAIL.n297 171.744
R114 VTAIL.n344 VTAIL.n343 171.744
R115 VTAIL.n344 VTAIL.n293 171.744
R116 VTAIL.n351 VTAIL.n293 171.744
R117 VTAIL.n353 VTAIL.n351 171.744
R118 VTAIL.n353 VTAIL.n352 171.744
R119 VTAIL.n352 VTAIL.n289 171.744
R120 VTAIL.n361 VTAIL.n289 171.744
R121 VTAIL.n362 VTAIL.n361 171.744
R122 VTAIL.n362 VTAIL.n285 171.744
R123 VTAIL.n369 VTAIL.n285 171.744
R124 VTAIL.n370 VTAIL.n369 171.744
R125 VTAIL.n30 VTAIL.n27 171.744
R126 VTAIL.n37 VTAIL.n27 171.744
R127 VTAIL.n38 VTAIL.n37 171.744
R128 VTAIL.n38 VTAIL.n23 171.744
R129 VTAIL.n45 VTAIL.n23 171.744
R130 VTAIL.n46 VTAIL.n45 171.744
R131 VTAIL.n46 VTAIL.n19 171.744
R132 VTAIL.n53 VTAIL.n19 171.744
R133 VTAIL.n54 VTAIL.n53 171.744
R134 VTAIL.n54 VTAIL.n15 171.744
R135 VTAIL.n61 VTAIL.n15 171.744
R136 VTAIL.n62 VTAIL.n61 171.744
R137 VTAIL.n62 VTAIL.n11 171.744
R138 VTAIL.n69 VTAIL.n11 171.744
R139 VTAIL.n71 VTAIL.n69 171.744
R140 VTAIL.n71 VTAIL.n70 171.744
R141 VTAIL.n70 VTAIL.n7 171.744
R142 VTAIL.n79 VTAIL.n7 171.744
R143 VTAIL.n80 VTAIL.n79 171.744
R144 VTAIL.n80 VTAIL.n3 171.744
R145 VTAIL.n87 VTAIL.n3 171.744
R146 VTAIL.n88 VTAIL.n87 171.744
R147 VTAIL.n276 VTAIL.n275 171.744
R148 VTAIL.n275 VTAIL.n191 171.744
R149 VTAIL.n268 VTAIL.n191 171.744
R150 VTAIL.n268 VTAIL.n267 171.744
R151 VTAIL.n267 VTAIL.n195 171.744
R152 VTAIL.n199 VTAIL.n195 171.744
R153 VTAIL.n259 VTAIL.n199 171.744
R154 VTAIL.n259 VTAIL.n258 171.744
R155 VTAIL.n258 VTAIL.n200 171.744
R156 VTAIL.n251 VTAIL.n200 171.744
R157 VTAIL.n251 VTAIL.n250 171.744
R158 VTAIL.n250 VTAIL.n204 171.744
R159 VTAIL.n243 VTAIL.n204 171.744
R160 VTAIL.n243 VTAIL.n242 171.744
R161 VTAIL.n242 VTAIL.n208 171.744
R162 VTAIL.n235 VTAIL.n208 171.744
R163 VTAIL.n235 VTAIL.n234 171.744
R164 VTAIL.n234 VTAIL.n212 171.744
R165 VTAIL.n227 VTAIL.n212 171.744
R166 VTAIL.n227 VTAIL.n226 171.744
R167 VTAIL.n226 VTAIL.n216 171.744
R168 VTAIL.n219 VTAIL.n216 171.744
R169 VTAIL.n182 VTAIL.n181 171.744
R170 VTAIL.n181 VTAIL.n97 171.744
R171 VTAIL.n174 VTAIL.n97 171.744
R172 VTAIL.n174 VTAIL.n173 171.744
R173 VTAIL.n173 VTAIL.n101 171.744
R174 VTAIL.n105 VTAIL.n101 171.744
R175 VTAIL.n165 VTAIL.n105 171.744
R176 VTAIL.n165 VTAIL.n164 171.744
R177 VTAIL.n164 VTAIL.n106 171.744
R178 VTAIL.n157 VTAIL.n106 171.744
R179 VTAIL.n157 VTAIL.n156 171.744
R180 VTAIL.n156 VTAIL.n110 171.744
R181 VTAIL.n149 VTAIL.n110 171.744
R182 VTAIL.n149 VTAIL.n148 171.744
R183 VTAIL.n148 VTAIL.n114 171.744
R184 VTAIL.n141 VTAIL.n114 171.744
R185 VTAIL.n141 VTAIL.n140 171.744
R186 VTAIL.n140 VTAIL.n118 171.744
R187 VTAIL.n133 VTAIL.n118 171.744
R188 VTAIL.n133 VTAIL.n132 171.744
R189 VTAIL.n132 VTAIL.n122 171.744
R190 VTAIL.n125 VTAIL.n122 171.744
R191 VTAIL.n312 VTAIL.t0 85.8723
R192 VTAIL.n30 VTAIL.t3 85.8723
R193 VTAIL.n219 VTAIL.t2 85.8723
R194 VTAIL.n125 VTAIL.t1 85.8723
R195 VTAIL.n375 VTAIL.n374 34.1247
R196 VTAIL.n93 VTAIL.n92 34.1247
R197 VTAIL.n281 VTAIL.n280 34.1247
R198 VTAIL.n187 VTAIL.n186 34.1247
R199 VTAIL.n187 VTAIL.n93 29.2117
R200 VTAIL.n375 VTAIL.n281 28.0824
R201 VTAIL.n313 VTAIL.n311 16.3895
R202 VTAIL.n31 VTAIL.n29 16.3895
R203 VTAIL.n220 VTAIL.n218 16.3895
R204 VTAIL.n126 VTAIL.n124 16.3895
R205 VTAIL.n360 VTAIL.n359 13.1884
R206 VTAIL.n78 VTAIL.n77 13.1884
R207 VTAIL.n266 VTAIL.n265 13.1884
R208 VTAIL.n172 VTAIL.n171 13.1884
R209 VTAIL.n314 VTAIL.n310 12.8005
R210 VTAIL.n358 VTAIL.n290 12.8005
R211 VTAIL.n363 VTAIL.n288 12.8005
R212 VTAIL.n32 VTAIL.n28 12.8005
R213 VTAIL.n76 VTAIL.n8 12.8005
R214 VTAIL.n81 VTAIL.n6 12.8005
R215 VTAIL.n269 VTAIL.n194 12.8005
R216 VTAIL.n264 VTAIL.n196 12.8005
R217 VTAIL.n221 VTAIL.n217 12.8005
R218 VTAIL.n175 VTAIL.n100 12.8005
R219 VTAIL.n170 VTAIL.n102 12.8005
R220 VTAIL.n127 VTAIL.n123 12.8005
R221 VTAIL.n318 VTAIL.n317 12.0247
R222 VTAIL.n355 VTAIL.n354 12.0247
R223 VTAIL.n364 VTAIL.n286 12.0247
R224 VTAIL.n36 VTAIL.n35 12.0247
R225 VTAIL.n73 VTAIL.n72 12.0247
R226 VTAIL.n82 VTAIL.n4 12.0247
R227 VTAIL.n270 VTAIL.n192 12.0247
R228 VTAIL.n261 VTAIL.n260 12.0247
R229 VTAIL.n225 VTAIL.n224 12.0247
R230 VTAIL.n176 VTAIL.n98 12.0247
R231 VTAIL.n167 VTAIL.n166 12.0247
R232 VTAIL.n131 VTAIL.n130 12.0247
R233 VTAIL.n321 VTAIL.n308 11.249
R234 VTAIL.n350 VTAIL.n292 11.249
R235 VTAIL.n368 VTAIL.n367 11.249
R236 VTAIL.n39 VTAIL.n26 11.249
R237 VTAIL.n68 VTAIL.n10 11.249
R238 VTAIL.n86 VTAIL.n85 11.249
R239 VTAIL.n274 VTAIL.n273 11.249
R240 VTAIL.n257 VTAIL.n198 11.249
R241 VTAIL.n228 VTAIL.n215 11.249
R242 VTAIL.n180 VTAIL.n179 11.249
R243 VTAIL.n163 VTAIL.n104 11.249
R244 VTAIL.n134 VTAIL.n121 11.249
R245 VTAIL.n322 VTAIL.n306 10.4732
R246 VTAIL.n349 VTAIL.n294 10.4732
R247 VTAIL.n371 VTAIL.n284 10.4732
R248 VTAIL.n40 VTAIL.n24 10.4732
R249 VTAIL.n67 VTAIL.n12 10.4732
R250 VTAIL.n89 VTAIL.n2 10.4732
R251 VTAIL.n277 VTAIL.n190 10.4732
R252 VTAIL.n256 VTAIL.n201 10.4732
R253 VTAIL.n229 VTAIL.n213 10.4732
R254 VTAIL.n183 VTAIL.n96 10.4732
R255 VTAIL.n162 VTAIL.n107 10.4732
R256 VTAIL.n135 VTAIL.n119 10.4732
R257 VTAIL.n326 VTAIL.n325 9.69747
R258 VTAIL.n346 VTAIL.n345 9.69747
R259 VTAIL.n372 VTAIL.n282 9.69747
R260 VTAIL.n44 VTAIL.n43 9.69747
R261 VTAIL.n64 VTAIL.n63 9.69747
R262 VTAIL.n90 VTAIL.n0 9.69747
R263 VTAIL.n278 VTAIL.n188 9.69747
R264 VTAIL.n253 VTAIL.n252 9.69747
R265 VTAIL.n233 VTAIL.n232 9.69747
R266 VTAIL.n184 VTAIL.n94 9.69747
R267 VTAIL.n159 VTAIL.n158 9.69747
R268 VTAIL.n139 VTAIL.n138 9.69747
R269 VTAIL.n374 VTAIL.n373 9.45567
R270 VTAIL.n92 VTAIL.n91 9.45567
R271 VTAIL.n280 VTAIL.n279 9.45567
R272 VTAIL.n186 VTAIL.n185 9.45567
R273 VTAIL.n373 VTAIL.n372 9.3005
R274 VTAIL.n284 VTAIL.n283 9.3005
R275 VTAIL.n367 VTAIL.n366 9.3005
R276 VTAIL.n365 VTAIL.n364 9.3005
R277 VTAIL.n288 VTAIL.n287 9.3005
R278 VTAIL.n333 VTAIL.n332 9.3005
R279 VTAIL.n331 VTAIL.n330 9.3005
R280 VTAIL.n304 VTAIL.n303 9.3005
R281 VTAIL.n325 VTAIL.n324 9.3005
R282 VTAIL.n323 VTAIL.n322 9.3005
R283 VTAIL.n308 VTAIL.n307 9.3005
R284 VTAIL.n317 VTAIL.n316 9.3005
R285 VTAIL.n315 VTAIL.n314 9.3005
R286 VTAIL.n300 VTAIL.n299 9.3005
R287 VTAIL.n339 VTAIL.n338 9.3005
R288 VTAIL.n341 VTAIL.n340 9.3005
R289 VTAIL.n296 VTAIL.n295 9.3005
R290 VTAIL.n347 VTAIL.n346 9.3005
R291 VTAIL.n349 VTAIL.n348 9.3005
R292 VTAIL.n292 VTAIL.n291 9.3005
R293 VTAIL.n356 VTAIL.n355 9.3005
R294 VTAIL.n358 VTAIL.n357 9.3005
R295 VTAIL.n91 VTAIL.n90 9.3005
R296 VTAIL.n2 VTAIL.n1 9.3005
R297 VTAIL.n85 VTAIL.n84 9.3005
R298 VTAIL.n83 VTAIL.n82 9.3005
R299 VTAIL.n6 VTAIL.n5 9.3005
R300 VTAIL.n51 VTAIL.n50 9.3005
R301 VTAIL.n49 VTAIL.n48 9.3005
R302 VTAIL.n22 VTAIL.n21 9.3005
R303 VTAIL.n43 VTAIL.n42 9.3005
R304 VTAIL.n41 VTAIL.n40 9.3005
R305 VTAIL.n26 VTAIL.n25 9.3005
R306 VTAIL.n35 VTAIL.n34 9.3005
R307 VTAIL.n33 VTAIL.n32 9.3005
R308 VTAIL.n18 VTAIL.n17 9.3005
R309 VTAIL.n57 VTAIL.n56 9.3005
R310 VTAIL.n59 VTAIL.n58 9.3005
R311 VTAIL.n14 VTAIL.n13 9.3005
R312 VTAIL.n65 VTAIL.n64 9.3005
R313 VTAIL.n67 VTAIL.n66 9.3005
R314 VTAIL.n10 VTAIL.n9 9.3005
R315 VTAIL.n74 VTAIL.n73 9.3005
R316 VTAIL.n76 VTAIL.n75 9.3005
R317 VTAIL.n246 VTAIL.n245 9.3005
R318 VTAIL.n248 VTAIL.n247 9.3005
R319 VTAIL.n203 VTAIL.n202 9.3005
R320 VTAIL.n254 VTAIL.n253 9.3005
R321 VTAIL.n256 VTAIL.n255 9.3005
R322 VTAIL.n198 VTAIL.n197 9.3005
R323 VTAIL.n262 VTAIL.n261 9.3005
R324 VTAIL.n264 VTAIL.n263 9.3005
R325 VTAIL.n279 VTAIL.n278 9.3005
R326 VTAIL.n190 VTAIL.n189 9.3005
R327 VTAIL.n273 VTAIL.n272 9.3005
R328 VTAIL.n271 VTAIL.n270 9.3005
R329 VTAIL.n194 VTAIL.n193 9.3005
R330 VTAIL.n207 VTAIL.n206 9.3005
R331 VTAIL.n240 VTAIL.n239 9.3005
R332 VTAIL.n238 VTAIL.n237 9.3005
R333 VTAIL.n211 VTAIL.n210 9.3005
R334 VTAIL.n232 VTAIL.n231 9.3005
R335 VTAIL.n230 VTAIL.n229 9.3005
R336 VTAIL.n215 VTAIL.n214 9.3005
R337 VTAIL.n224 VTAIL.n223 9.3005
R338 VTAIL.n222 VTAIL.n221 9.3005
R339 VTAIL.n152 VTAIL.n151 9.3005
R340 VTAIL.n154 VTAIL.n153 9.3005
R341 VTAIL.n109 VTAIL.n108 9.3005
R342 VTAIL.n160 VTAIL.n159 9.3005
R343 VTAIL.n162 VTAIL.n161 9.3005
R344 VTAIL.n104 VTAIL.n103 9.3005
R345 VTAIL.n168 VTAIL.n167 9.3005
R346 VTAIL.n170 VTAIL.n169 9.3005
R347 VTAIL.n185 VTAIL.n184 9.3005
R348 VTAIL.n96 VTAIL.n95 9.3005
R349 VTAIL.n179 VTAIL.n178 9.3005
R350 VTAIL.n177 VTAIL.n176 9.3005
R351 VTAIL.n100 VTAIL.n99 9.3005
R352 VTAIL.n113 VTAIL.n112 9.3005
R353 VTAIL.n146 VTAIL.n145 9.3005
R354 VTAIL.n144 VTAIL.n143 9.3005
R355 VTAIL.n117 VTAIL.n116 9.3005
R356 VTAIL.n138 VTAIL.n137 9.3005
R357 VTAIL.n136 VTAIL.n135 9.3005
R358 VTAIL.n121 VTAIL.n120 9.3005
R359 VTAIL.n130 VTAIL.n129 9.3005
R360 VTAIL.n128 VTAIL.n127 9.3005
R361 VTAIL.n329 VTAIL.n304 8.92171
R362 VTAIL.n342 VTAIL.n296 8.92171
R363 VTAIL.n47 VTAIL.n22 8.92171
R364 VTAIL.n60 VTAIL.n14 8.92171
R365 VTAIL.n249 VTAIL.n203 8.92171
R366 VTAIL.n236 VTAIL.n211 8.92171
R367 VTAIL.n155 VTAIL.n109 8.92171
R368 VTAIL.n142 VTAIL.n117 8.92171
R369 VTAIL.n330 VTAIL.n302 8.14595
R370 VTAIL.n341 VTAIL.n298 8.14595
R371 VTAIL.n48 VTAIL.n20 8.14595
R372 VTAIL.n59 VTAIL.n16 8.14595
R373 VTAIL.n248 VTAIL.n205 8.14595
R374 VTAIL.n237 VTAIL.n209 8.14595
R375 VTAIL.n154 VTAIL.n111 8.14595
R376 VTAIL.n143 VTAIL.n115 8.14595
R377 VTAIL.n334 VTAIL.n333 7.3702
R378 VTAIL.n338 VTAIL.n337 7.3702
R379 VTAIL.n52 VTAIL.n51 7.3702
R380 VTAIL.n56 VTAIL.n55 7.3702
R381 VTAIL.n245 VTAIL.n244 7.3702
R382 VTAIL.n241 VTAIL.n240 7.3702
R383 VTAIL.n151 VTAIL.n150 7.3702
R384 VTAIL.n147 VTAIL.n146 7.3702
R385 VTAIL.n334 VTAIL.n300 6.59444
R386 VTAIL.n337 VTAIL.n300 6.59444
R387 VTAIL.n52 VTAIL.n18 6.59444
R388 VTAIL.n55 VTAIL.n18 6.59444
R389 VTAIL.n244 VTAIL.n207 6.59444
R390 VTAIL.n241 VTAIL.n207 6.59444
R391 VTAIL.n150 VTAIL.n113 6.59444
R392 VTAIL.n147 VTAIL.n113 6.59444
R393 VTAIL.n333 VTAIL.n302 5.81868
R394 VTAIL.n338 VTAIL.n298 5.81868
R395 VTAIL.n51 VTAIL.n20 5.81868
R396 VTAIL.n56 VTAIL.n16 5.81868
R397 VTAIL.n245 VTAIL.n205 5.81868
R398 VTAIL.n240 VTAIL.n209 5.81868
R399 VTAIL.n151 VTAIL.n111 5.81868
R400 VTAIL.n146 VTAIL.n115 5.81868
R401 VTAIL.n330 VTAIL.n329 5.04292
R402 VTAIL.n342 VTAIL.n341 5.04292
R403 VTAIL.n48 VTAIL.n47 5.04292
R404 VTAIL.n60 VTAIL.n59 5.04292
R405 VTAIL.n249 VTAIL.n248 5.04292
R406 VTAIL.n237 VTAIL.n236 5.04292
R407 VTAIL.n155 VTAIL.n154 5.04292
R408 VTAIL.n143 VTAIL.n142 5.04292
R409 VTAIL.n326 VTAIL.n304 4.26717
R410 VTAIL.n345 VTAIL.n296 4.26717
R411 VTAIL.n374 VTAIL.n282 4.26717
R412 VTAIL.n44 VTAIL.n22 4.26717
R413 VTAIL.n63 VTAIL.n14 4.26717
R414 VTAIL.n92 VTAIL.n0 4.26717
R415 VTAIL.n280 VTAIL.n188 4.26717
R416 VTAIL.n252 VTAIL.n203 4.26717
R417 VTAIL.n233 VTAIL.n211 4.26717
R418 VTAIL.n186 VTAIL.n94 4.26717
R419 VTAIL.n158 VTAIL.n109 4.26717
R420 VTAIL.n139 VTAIL.n117 4.26717
R421 VTAIL.n315 VTAIL.n311 3.70982
R422 VTAIL.n33 VTAIL.n29 3.70982
R423 VTAIL.n222 VTAIL.n218 3.70982
R424 VTAIL.n128 VTAIL.n124 3.70982
R425 VTAIL.n325 VTAIL.n306 3.49141
R426 VTAIL.n346 VTAIL.n294 3.49141
R427 VTAIL.n372 VTAIL.n371 3.49141
R428 VTAIL.n43 VTAIL.n24 3.49141
R429 VTAIL.n64 VTAIL.n12 3.49141
R430 VTAIL.n90 VTAIL.n89 3.49141
R431 VTAIL.n278 VTAIL.n277 3.49141
R432 VTAIL.n253 VTAIL.n201 3.49141
R433 VTAIL.n232 VTAIL.n213 3.49141
R434 VTAIL.n184 VTAIL.n183 3.49141
R435 VTAIL.n159 VTAIL.n107 3.49141
R436 VTAIL.n138 VTAIL.n119 3.49141
R437 VTAIL.n322 VTAIL.n321 2.71565
R438 VTAIL.n350 VTAIL.n349 2.71565
R439 VTAIL.n368 VTAIL.n284 2.71565
R440 VTAIL.n40 VTAIL.n39 2.71565
R441 VTAIL.n68 VTAIL.n67 2.71565
R442 VTAIL.n86 VTAIL.n2 2.71565
R443 VTAIL.n274 VTAIL.n190 2.71565
R444 VTAIL.n257 VTAIL.n256 2.71565
R445 VTAIL.n229 VTAIL.n228 2.71565
R446 VTAIL.n180 VTAIL.n96 2.71565
R447 VTAIL.n163 VTAIL.n162 2.71565
R448 VTAIL.n135 VTAIL.n134 2.71565
R449 VTAIL.n318 VTAIL.n308 1.93989
R450 VTAIL.n354 VTAIL.n292 1.93989
R451 VTAIL.n367 VTAIL.n286 1.93989
R452 VTAIL.n36 VTAIL.n26 1.93989
R453 VTAIL.n72 VTAIL.n10 1.93989
R454 VTAIL.n85 VTAIL.n4 1.93989
R455 VTAIL.n273 VTAIL.n192 1.93989
R456 VTAIL.n260 VTAIL.n198 1.93989
R457 VTAIL.n225 VTAIL.n215 1.93989
R458 VTAIL.n179 VTAIL.n98 1.93989
R459 VTAIL.n166 VTAIL.n104 1.93989
R460 VTAIL.n131 VTAIL.n121 1.93989
R461 VTAIL.n317 VTAIL.n310 1.16414
R462 VTAIL.n355 VTAIL.n290 1.16414
R463 VTAIL.n364 VTAIL.n363 1.16414
R464 VTAIL.n35 VTAIL.n28 1.16414
R465 VTAIL.n73 VTAIL.n8 1.16414
R466 VTAIL.n82 VTAIL.n81 1.16414
R467 VTAIL.n270 VTAIL.n269 1.16414
R468 VTAIL.n261 VTAIL.n196 1.16414
R469 VTAIL.n224 VTAIL.n217 1.16414
R470 VTAIL.n176 VTAIL.n175 1.16414
R471 VTAIL.n167 VTAIL.n102 1.16414
R472 VTAIL.n130 VTAIL.n123 1.16414
R473 VTAIL.n281 VTAIL.n187 1.03498
R474 VTAIL VTAIL.n93 0.810845
R475 VTAIL.n314 VTAIL.n313 0.388379
R476 VTAIL.n359 VTAIL.n358 0.388379
R477 VTAIL.n360 VTAIL.n288 0.388379
R478 VTAIL.n32 VTAIL.n31 0.388379
R479 VTAIL.n77 VTAIL.n76 0.388379
R480 VTAIL.n78 VTAIL.n6 0.388379
R481 VTAIL.n266 VTAIL.n194 0.388379
R482 VTAIL.n265 VTAIL.n264 0.388379
R483 VTAIL.n221 VTAIL.n220 0.388379
R484 VTAIL.n172 VTAIL.n100 0.388379
R485 VTAIL.n171 VTAIL.n170 0.388379
R486 VTAIL.n127 VTAIL.n126 0.388379
R487 VTAIL VTAIL.n375 0.224638
R488 VTAIL.n316 VTAIL.n315 0.155672
R489 VTAIL.n316 VTAIL.n307 0.155672
R490 VTAIL.n323 VTAIL.n307 0.155672
R491 VTAIL.n324 VTAIL.n323 0.155672
R492 VTAIL.n324 VTAIL.n303 0.155672
R493 VTAIL.n331 VTAIL.n303 0.155672
R494 VTAIL.n332 VTAIL.n331 0.155672
R495 VTAIL.n332 VTAIL.n299 0.155672
R496 VTAIL.n339 VTAIL.n299 0.155672
R497 VTAIL.n340 VTAIL.n339 0.155672
R498 VTAIL.n340 VTAIL.n295 0.155672
R499 VTAIL.n347 VTAIL.n295 0.155672
R500 VTAIL.n348 VTAIL.n347 0.155672
R501 VTAIL.n348 VTAIL.n291 0.155672
R502 VTAIL.n356 VTAIL.n291 0.155672
R503 VTAIL.n357 VTAIL.n356 0.155672
R504 VTAIL.n357 VTAIL.n287 0.155672
R505 VTAIL.n365 VTAIL.n287 0.155672
R506 VTAIL.n366 VTAIL.n365 0.155672
R507 VTAIL.n366 VTAIL.n283 0.155672
R508 VTAIL.n373 VTAIL.n283 0.155672
R509 VTAIL.n34 VTAIL.n33 0.155672
R510 VTAIL.n34 VTAIL.n25 0.155672
R511 VTAIL.n41 VTAIL.n25 0.155672
R512 VTAIL.n42 VTAIL.n41 0.155672
R513 VTAIL.n42 VTAIL.n21 0.155672
R514 VTAIL.n49 VTAIL.n21 0.155672
R515 VTAIL.n50 VTAIL.n49 0.155672
R516 VTAIL.n50 VTAIL.n17 0.155672
R517 VTAIL.n57 VTAIL.n17 0.155672
R518 VTAIL.n58 VTAIL.n57 0.155672
R519 VTAIL.n58 VTAIL.n13 0.155672
R520 VTAIL.n65 VTAIL.n13 0.155672
R521 VTAIL.n66 VTAIL.n65 0.155672
R522 VTAIL.n66 VTAIL.n9 0.155672
R523 VTAIL.n74 VTAIL.n9 0.155672
R524 VTAIL.n75 VTAIL.n74 0.155672
R525 VTAIL.n75 VTAIL.n5 0.155672
R526 VTAIL.n83 VTAIL.n5 0.155672
R527 VTAIL.n84 VTAIL.n83 0.155672
R528 VTAIL.n84 VTAIL.n1 0.155672
R529 VTAIL.n91 VTAIL.n1 0.155672
R530 VTAIL.n279 VTAIL.n189 0.155672
R531 VTAIL.n272 VTAIL.n189 0.155672
R532 VTAIL.n272 VTAIL.n271 0.155672
R533 VTAIL.n271 VTAIL.n193 0.155672
R534 VTAIL.n263 VTAIL.n193 0.155672
R535 VTAIL.n263 VTAIL.n262 0.155672
R536 VTAIL.n262 VTAIL.n197 0.155672
R537 VTAIL.n255 VTAIL.n197 0.155672
R538 VTAIL.n255 VTAIL.n254 0.155672
R539 VTAIL.n254 VTAIL.n202 0.155672
R540 VTAIL.n247 VTAIL.n202 0.155672
R541 VTAIL.n247 VTAIL.n246 0.155672
R542 VTAIL.n246 VTAIL.n206 0.155672
R543 VTAIL.n239 VTAIL.n206 0.155672
R544 VTAIL.n239 VTAIL.n238 0.155672
R545 VTAIL.n238 VTAIL.n210 0.155672
R546 VTAIL.n231 VTAIL.n210 0.155672
R547 VTAIL.n231 VTAIL.n230 0.155672
R548 VTAIL.n230 VTAIL.n214 0.155672
R549 VTAIL.n223 VTAIL.n214 0.155672
R550 VTAIL.n223 VTAIL.n222 0.155672
R551 VTAIL.n185 VTAIL.n95 0.155672
R552 VTAIL.n178 VTAIL.n95 0.155672
R553 VTAIL.n178 VTAIL.n177 0.155672
R554 VTAIL.n177 VTAIL.n99 0.155672
R555 VTAIL.n169 VTAIL.n99 0.155672
R556 VTAIL.n169 VTAIL.n168 0.155672
R557 VTAIL.n168 VTAIL.n103 0.155672
R558 VTAIL.n161 VTAIL.n103 0.155672
R559 VTAIL.n161 VTAIL.n160 0.155672
R560 VTAIL.n160 VTAIL.n108 0.155672
R561 VTAIL.n153 VTAIL.n108 0.155672
R562 VTAIL.n153 VTAIL.n152 0.155672
R563 VTAIL.n152 VTAIL.n112 0.155672
R564 VTAIL.n145 VTAIL.n112 0.155672
R565 VTAIL.n145 VTAIL.n144 0.155672
R566 VTAIL.n144 VTAIL.n116 0.155672
R567 VTAIL.n137 VTAIL.n116 0.155672
R568 VTAIL.n137 VTAIL.n136 0.155672
R569 VTAIL.n136 VTAIL.n120 0.155672
R570 VTAIL.n129 VTAIL.n120 0.155672
R571 VTAIL.n129 VTAIL.n128 0.155672
R572 VDD1.n88 VDD1.n0 756.745
R573 VDD1.n181 VDD1.n93 756.745
R574 VDD1.n89 VDD1.n88 585
R575 VDD1.n87 VDD1.n86 585
R576 VDD1.n4 VDD1.n3 585
R577 VDD1.n81 VDD1.n80 585
R578 VDD1.n79 VDD1.n78 585
R579 VDD1.n77 VDD1.n7 585
R580 VDD1.n11 VDD1.n8 585
R581 VDD1.n72 VDD1.n71 585
R582 VDD1.n70 VDD1.n69 585
R583 VDD1.n13 VDD1.n12 585
R584 VDD1.n64 VDD1.n63 585
R585 VDD1.n62 VDD1.n61 585
R586 VDD1.n17 VDD1.n16 585
R587 VDD1.n56 VDD1.n55 585
R588 VDD1.n54 VDD1.n53 585
R589 VDD1.n21 VDD1.n20 585
R590 VDD1.n48 VDD1.n47 585
R591 VDD1.n46 VDD1.n45 585
R592 VDD1.n25 VDD1.n24 585
R593 VDD1.n40 VDD1.n39 585
R594 VDD1.n38 VDD1.n37 585
R595 VDD1.n29 VDD1.n28 585
R596 VDD1.n32 VDD1.n31 585
R597 VDD1.n124 VDD1.n123 585
R598 VDD1.n121 VDD1.n120 585
R599 VDD1.n130 VDD1.n129 585
R600 VDD1.n132 VDD1.n131 585
R601 VDD1.n117 VDD1.n116 585
R602 VDD1.n138 VDD1.n137 585
R603 VDD1.n140 VDD1.n139 585
R604 VDD1.n113 VDD1.n112 585
R605 VDD1.n146 VDD1.n145 585
R606 VDD1.n148 VDD1.n147 585
R607 VDD1.n109 VDD1.n108 585
R608 VDD1.n154 VDD1.n153 585
R609 VDD1.n156 VDD1.n155 585
R610 VDD1.n105 VDD1.n104 585
R611 VDD1.n162 VDD1.n161 585
R612 VDD1.n165 VDD1.n164 585
R613 VDD1.n163 VDD1.n101 585
R614 VDD1.n170 VDD1.n100 585
R615 VDD1.n172 VDD1.n171 585
R616 VDD1.n174 VDD1.n173 585
R617 VDD1.n97 VDD1.n96 585
R618 VDD1.n180 VDD1.n179 585
R619 VDD1.n182 VDD1.n181 585
R620 VDD1.t1 VDD1.n30 327.466
R621 VDD1.t0 VDD1.n122 327.466
R622 VDD1.n88 VDD1.n87 171.744
R623 VDD1.n87 VDD1.n3 171.744
R624 VDD1.n80 VDD1.n3 171.744
R625 VDD1.n80 VDD1.n79 171.744
R626 VDD1.n79 VDD1.n7 171.744
R627 VDD1.n11 VDD1.n7 171.744
R628 VDD1.n71 VDD1.n11 171.744
R629 VDD1.n71 VDD1.n70 171.744
R630 VDD1.n70 VDD1.n12 171.744
R631 VDD1.n63 VDD1.n12 171.744
R632 VDD1.n63 VDD1.n62 171.744
R633 VDD1.n62 VDD1.n16 171.744
R634 VDD1.n55 VDD1.n16 171.744
R635 VDD1.n55 VDD1.n54 171.744
R636 VDD1.n54 VDD1.n20 171.744
R637 VDD1.n47 VDD1.n20 171.744
R638 VDD1.n47 VDD1.n46 171.744
R639 VDD1.n46 VDD1.n24 171.744
R640 VDD1.n39 VDD1.n24 171.744
R641 VDD1.n39 VDD1.n38 171.744
R642 VDD1.n38 VDD1.n28 171.744
R643 VDD1.n31 VDD1.n28 171.744
R644 VDD1.n123 VDD1.n120 171.744
R645 VDD1.n130 VDD1.n120 171.744
R646 VDD1.n131 VDD1.n130 171.744
R647 VDD1.n131 VDD1.n116 171.744
R648 VDD1.n138 VDD1.n116 171.744
R649 VDD1.n139 VDD1.n138 171.744
R650 VDD1.n139 VDD1.n112 171.744
R651 VDD1.n146 VDD1.n112 171.744
R652 VDD1.n147 VDD1.n146 171.744
R653 VDD1.n147 VDD1.n108 171.744
R654 VDD1.n154 VDD1.n108 171.744
R655 VDD1.n155 VDD1.n154 171.744
R656 VDD1.n155 VDD1.n104 171.744
R657 VDD1.n162 VDD1.n104 171.744
R658 VDD1.n164 VDD1.n162 171.744
R659 VDD1.n164 VDD1.n163 171.744
R660 VDD1.n163 VDD1.n100 171.744
R661 VDD1.n172 VDD1.n100 171.744
R662 VDD1.n173 VDD1.n172 171.744
R663 VDD1.n173 VDD1.n96 171.744
R664 VDD1.n180 VDD1.n96 171.744
R665 VDD1.n181 VDD1.n180 171.744
R666 VDD1 VDD1.n185 92.115
R667 VDD1.n31 VDD1.t1 85.8723
R668 VDD1.n123 VDD1.t0 85.8723
R669 VDD1 VDD1.n92 51.144
R670 VDD1.n32 VDD1.n30 16.3895
R671 VDD1.n124 VDD1.n122 16.3895
R672 VDD1.n78 VDD1.n77 13.1884
R673 VDD1.n171 VDD1.n170 13.1884
R674 VDD1.n81 VDD1.n6 12.8005
R675 VDD1.n76 VDD1.n8 12.8005
R676 VDD1.n33 VDD1.n29 12.8005
R677 VDD1.n125 VDD1.n121 12.8005
R678 VDD1.n169 VDD1.n101 12.8005
R679 VDD1.n174 VDD1.n99 12.8005
R680 VDD1.n82 VDD1.n4 12.0247
R681 VDD1.n73 VDD1.n72 12.0247
R682 VDD1.n37 VDD1.n36 12.0247
R683 VDD1.n129 VDD1.n128 12.0247
R684 VDD1.n166 VDD1.n165 12.0247
R685 VDD1.n175 VDD1.n97 12.0247
R686 VDD1.n86 VDD1.n85 11.249
R687 VDD1.n69 VDD1.n10 11.249
R688 VDD1.n40 VDD1.n27 11.249
R689 VDD1.n132 VDD1.n119 11.249
R690 VDD1.n161 VDD1.n103 11.249
R691 VDD1.n179 VDD1.n178 11.249
R692 VDD1.n89 VDD1.n2 10.4732
R693 VDD1.n68 VDD1.n13 10.4732
R694 VDD1.n41 VDD1.n25 10.4732
R695 VDD1.n133 VDD1.n117 10.4732
R696 VDD1.n160 VDD1.n105 10.4732
R697 VDD1.n182 VDD1.n95 10.4732
R698 VDD1.n90 VDD1.n0 9.69747
R699 VDD1.n65 VDD1.n64 9.69747
R700 VDD1.n45 VDD1.n44 9.69747
R701 VDD1.n137 VDD1.n136 9.69747
R702 VDD1.n157 VDD1.n156 9.69747
R703 VDD1.n183 VDD1.n93 9.69747
R704 VDD1.n92 VDD1.n91 9.45567
R705 VDD1.n185 VDD1.n184 9.45567
R706 VDD1.n58 VDD1.n57 9.3005
R707 VDD1.n60 VDD1.n59 9.3005
R708 VDD1.n15 VDD1.n14 9.3005
R709 VDD1.n66 VDD1.n65 9.3005
R710 VDD1.n68 VDD1.n67 9.3005
R711 VDD1.n10 VDD1.n9 9.3005
R712 VDD1.n74 VDD1.n73 9.3005
R713 VDD1.n76 VDD1.n75 9.3005
R714 VDD1.n91 VDD1.n90 9.3005
R715 VDD1.n2 VDD1.n1 9.3005
R716 VDD1.n85 VDD1.n84 9.3005
R717 VDD1.n83 VDD1.n82 9.3005
R718 VDD1.n6 VDD1.n5 9.3005
R719 VDD1.n19 VDD1.n18 9.3005
R720 VDD1.n52 VDD1.n51 9.3005
R721 VDD1.n50 VDD1.n49 9.3005
R722 VDD1.n23 VDD1.n22 9.3005
R723 VDD1.n44 VDD1.n43 9.3005
R724 VDD1.n42 VDD1.n41 9.3005
R725 VDD1.n27 VDD1.n26 9.3005
R726 VDD1.n36 VDD1.n35 9.3005
R727 VDD1.n34 VDD1.n33 9.3005
R728 VDD1.n184 VDD1.n183 9.3005
R729 VDD1.n95 VDD1.n94 9.3005
R730 VDD1.n178 VDD1.n177 9.3005
R731 VDD1.n176 VDD1.n175 9.3005
R732 VDD1.n99 VDD1.n98 9.3005
R733 VDD1.n144 VDD1.n143 9.3005
R734 VDD1.n142 VDD1.n141 9.3005
R735 VDD1.n115 VDD1.n114 9.3005
R736 VDD1.n136 VDD1.n135 9.3005
R737 VDD1.n134 VDD1.n133 9.3005
R738 VDD1.n119 VDD1.n118 9.3005
R739 VDD1.n128 VDD1.n127 9.3005
R740 VDD1.n126 VDD1.n125 9.3005
R741 VDD1.n111 VDD1.n110 9.3005
R742 VDD1.n150 VDD1.n149 9.3005
R743 VDD1.n152 VDD1.n151 9.3005
R744 VDD1.n107 VDD1.n106 9.3005
R745 VDD1.n158 VDD1.n157 9.3005
R746 VDD1.n160 VDD1.n159 9.3005
R747 VDD1.n103 VDD1.n102 9.3005
R748 VDD1.n167 VDD1.n166 9.3005
R749 VDD1.n169 VDD1.n168 9.3005
R750 VDD1.n61 VDD1.n15 8.92171
R751 VDD1.n48 VDD1.n23 8.92171
R752 VDD1.n140 VDD1.n115 8.92171
R753 VDD1.n153 VDD1.n107 8.92171
R754 VDD1.n60 VDD1.n17 8.14595
R755 VDD1.n49 VDD1.n21 8.14595
R756 VDD1.n141 VDD1.n113 8.14595
R757 VDD1.n152 VDD1.n109 8.14595
R758 VDD1.n57 VDD1.n56 7.3702
R759 VDD1.n53 VDD1.n52 7.3702
R760 VDD1.n145 VDD1.n144 7.3702
R761 VDD1.n149 VDD1.n148 7.3702
R762 VDD1.n56 VDD1.n19 6.59444
R763 VDD1.n53 VDD1.n19 6.59444
R764 VDD1.n145 VDD1.n111 6.59444
R765 VDD1.n148 VDD1.n111 6.59444
R766 VDD1.n57 VDD1.n17 5.81868
R767 VDD1.n52 VDD1.n21 5.81868
R768 VDD1.n144 VDD1.n113 5.81868
R769 VDD1.n149 VDD1.n109 5.81868
R770 VDD1.n61 VDD1.n60 5.04292
R771 VDD1.n49 VDD1.n48 5.04292
R772 VDD1.n141 VDD1.n140 5.04292
R773 VDD1.n153 VDD1.n152 5.04292
R774 VDD1.n92 VDD1.n0 4.26717
R775 VDD1.n64 VDD1.n15 4.26717
R776 VDD1.n45 VDD1.n23 4.26717
R777 VDD1.n137 VDD1.n115 4.26717
R778 VDD1.n156 VDD1.n107 4.26717
R779 VDD1.n185 VDD1.n93 4.26717
R780 VDD1.n34 VDD1.n30 3.70982
R781 VDD1.n126 VDD1.n122 3.70982
R782 VDD1.n90 VDD1.n89 3.49141
R783 VDD1.n65 VDD1.n13 3.49141
R784 VDD1.n44 VDD1.n25 3.49141
R785 VDD1.n136 VDD1.n117 3.49141
R786 VDD1.n157 VDD1.n105 3.49141
R787 VDD1.n183 VDD1.n182 3.49141
R788 VDD1.n86 VDD1.n2 2.71565
R789 VDD1.n69 VDD1.n68 2.71565
R790 VDD1.n41 VDD1.n40 2.71565
R791 VDD1.n133 VDD1.n132 2.71565
R792 VDD1.n161 VDD1.n160 2.71565
R793 VDD1.n179 VDD1.n95 2.71565
R794 VDD1.n85 VDD1.n4 1.93989
R795 VDD1.n72 VDD1.n10 1.93989
R796 VDD1.n37 VDD1.n27 1.93989
R797 VDD1.n129 VDD1.n119 1.93989
R798 VDD1.n165 VDD1.n103 1.93989
R799 VDD1.n178 VDD1.n97 1.93989
R800 VDD1.n82 VDD1.n81 1.16414
R801 VDD1.n73 VDD1.n8 1.16414
R802 VDD1.n36 VDD1.n29 1.16414
R803 VDD1.n128 VDD1.n121 1.16414
R804 VDD1.n166 VDD1.n101 1.16414
R805 VDD1.n175 VDD1.n174 1.16414
R806 VDD1.n78 VDD1.n6 0.388379
R807 VDD1.n77 VDD1.n76 0.388379
R808 VDD1.n33 VDD1.n32 0.388379
R809 VDD1.n125 VDD1.n124 0.388379
R810 VDD1.n170 VDD1.n169 0.388379
R811 VDD1.n171 VDD1.n99 0.388379
R812 VDD1.n91 VDD1.n1 0.155672
R813 VDD1.n84 VDD1.n1 0.155672
R814 VDD1.n84 VDD1.n83 0.155672
R815 VDD1.n83 VDD1.n5 0.155672
R816 VDD1.n75 VDD1.n5 0.155672
R817 VDD1.n75 VDD1.n74 0.155672
R818 VDD1.n74 VDD1.n9 0.155672
R819 VDD1.n67 VDD1.n9 0.155672
R820 VDD1.n67 VDD1.n66 0.155672
R821 VDD1.n66 VDD1.n14 0.155672
R822 VDD1.n59 VDD1.n14 0.155672
R823 VDD1.n59 VDD1.n58 0.155672
R824 VDD1.n58 VDD1.n18 0.155672
R825 VDD1.n51 VDD1.n18 0.155672
R826 VDD1.n51 VDD1.n50 0.155672
R827 VDD1.n50 VDD1.n22 0.155672
R828 VDD1.n43 VDD1.n22 0.155672
R829 VDD1.n43 VDD1.n42 0.155672
R830 VDD1.n42 VDD1.n26 0.155672
R831 VDD1.n35 VDD1.n26 0.155672
R832 VDD1.n35 VDD1.n34 0.155672
R833 VDD1.n127 VDD1.n126 0.155672
R834 VDD1.n127 VDD1.n118 0.155672
R835 VDD1.n134 VDD1.n118 0.155672
R836 VDD1.n135 VDD1.n134 0.155672
R837 VDD1.n135 VDD1.n114 0.155672
R838 VDD1.n142 VDD1.n114 0.155672
R839 VDD1.n143 VDD1.n142 0.155672
R840 VDD1.n143 VDD1.n110 0.155672
R841 VDD1.n150 VDD1.n110 0.155672
R842 VDD1.n151 VDD1.n150 0.155672
R843 VDD1.n151 VDD1.n106 0.155672
R844 VDD1.n158 VDD1.n106 0.155672
R845 VDD1.n159 VDD1.n158 0.155672
R846 VDD1.n159 VDD1.n102 0.155672
R847 VDD1.n167 VDD1.n102 0.155672
R848 VDD1.n168 VDD1.n167 0.155672
R849 VDD1.n168 VDD1.n98 0.155672
R850 VDD1.n176 VDD1.n98 0.155672
R851 VDD1.n177 VDD1.n176 0.155672
R852 VDD1.n177 VDD1.n94 0.155672
R853 VDD1.n184 VDD1.n94 0.155672
R854 VN VN.t1 661.456
R855 VN VN.t0 617.038
R856 VDD2.n181 VDD2.n93 756.745
R857 VDD2.n88 VDD2.n0 756.745
R858 VDD2.n182 VDD2.n181 585
R859 VDD2.n180 VDD2.n179 585
R860 VDD2.n97 VDD2.n96 585
R861 VDD2.n174 VDD2.n173 585
R862 VDD2.n172 VDD2.n171 585
R863 VDD2.n170 VDD2.n100 585
R864 VDD2.n104 VDD2.n101 585
R865 VDD2.n165 VDD2.n164 585
R866 VDD2.n163 VDD2.n162 585
R867 VDD2.n106 VDD2.n105 585
R868 VDD2.n157 VDD2.n156 585
R869 VDD2.n155 VDD2.n154 585
R870 VDD2.n110 VDD2.n109 585
R871 VDD2.n149 VDD2.n148 585
R872 VDD2.n147 VDD2.n146 585
R873 VDD2.n114 VDD2.n113 585
R874 VDD2.n141 VDD2.n140 585
R875 VDD2.n139 VDD2.n138 585
R876 VDD2.n118 VDD2.n117 585
R877 VDD2.n133 VDD2.n132 585
R878 VDD2.n131 VDD2.n130 585
R879 VDD2.n122 VDD2.n121 585
R880 VDD2.n125 VDD2.n124 585
R881 VDD2.n31 VDD2.n30 585
R882 VDD2.n28 VDD2.n27 585
R883 VDD2.n37 VDD2.n36 585
R884 VDD2.n39 VDD2.n38 585
R885 VDD2.n24 VDD2.n23 585
R886 VDD2.n45 VDD2.n44 585
R887 VDD2.n47 VDD2.n46 585
R888 VDD2.n20 VDD2.n19 585
R889 VDD2.n53 VDD2.n52 585
R890 VDD2.n55 VDD2.n54 585
R891 VDD2.n16 VDD2.n15 585
R892 VDD2.n61 VDD2.n60 585
R893 VDD2.n63 VDD2.n62 585
R894 VDD2.n12 VDD2.n11 585
R895 VDD2.n69 VDD2.n68 585
R896 VDD2.n72 VDD2.n71 585
R897 VDD2.n70 VDD2.n8 585
R898 VDD2.n77 VDD2.n7 585
R899 VDD2.n79 VDD2.n78 585
R900 VDD2.n81 VDD2.n80 585
R901 VDD2.n4 VDD2.n3 585
R902 VDD2.n87 VDD2.n86 585
R903 VDD2.n89 VDD2.n88 585
R904 VDD2.t0 VDD2.n123 327.466
R905 VDD2.t1 VDD2.n29 327.466
R906 VDD2.n181 VDD2.n180 171.744
R907 VDD2.n180 VDD2.n96 171.744
R908 VDD2.n173 VDD2.n96 171.744
R909 VDD2.n173 VDD2.n172 171.744
R910 VDD2.n172 VDD2.n100 171.744
R911 VDD2.n104 VDD2.n100 171.744
R912 VDD2.n164 VDD2.n104 171.744
R913 VDD2.n164 VDD2.n163 171.744
R914 VDD2.n163 VDD2.n105 171.744
R915 VDD2.n156 VDD2.n105 171.744
R916 VDD2.n156 VDD2.n155 171.744
R917 VDD2.n155 VDD2.n109 171.744
R918 VDD2.n148 VDD2.n109 171.744
R919 VDD2.n148 VDD2.n147 171.744
R920 VDD2.n147 VDD2.n113 171.744
R921 VDD2.n140 VDD2.n113 171.744
R922 VDD2.n140 VDD2.n139 171.744
R923 VDD2.n139 VDD2.n117 171.744
R924 VDD2.n132 VDD2.n117 171.744
R925 VDD2.n132 VDD2.n131 171.744
R926 VDD2.n131 VDD2.n121 171.744
R927 VDD2.n124 VDD2.n121 171.744
R928 VDD2.n30 VDD2.n27 171.744
R929 VDD2.n37 VDD2.n27 171.744
R930 VDD2.n38 VDD2.n37 171.744
R931 VDD2.n38 VDD2.n23 171.744
R932 VDD2.n45 VDD2.n23 171.744
R933 VDD2.n46 VDD2.n45 171.744
R934 VDD2.n46 VDD2.n19 171.744
R935 VDD2.n53 VDD2.n19 171.744
R936 VDD2.n54 VDD2.n53 171.744
R937 VDD2.n54 VDD2.n15 171.744
R938 VDD2.n61 VDD2.n15 171.744
R939 VDD2.n62 VDD2.n61 171.744
R940 VDD2.n62 VDD2.n11 171.744
R941 VDD2.n69 VDD2.n11 171.744
R942 VDD2.n71 VDD2.n69 171.744
R943 VDD2.n71 VDD2.n70 171.744
R944 VDD2.n70 VDD2.n7 171.744
R945 VDD2.n79 VDD2.n7 171.744
R946 VDD2.n80 VDD2.n79 171.744
R947 VDD2.n80 VDD2.n3 171.744
R948 VDD2.n87 VDD2.n3 171.744
R949 VDD2.n88 VDD2.n87 171.744
R950 VDD2.n186 VDD2.n92 91.3078
R951 VDD2.n124 VDD2.t0 85.8723
R952 VDD2.n30 VDD2.t1 85.8723
R953 VDD2.n186 VDD2.n185 50.8035
R954 VDD2.n125 VDD2.n123 16.3895
R955 VDD2.n31 VDD2.n29 16.3895
R956 VDD2.n171 VDD2.n170 13.1884
R957 VDD2.n78 VDD2.n77 13.1884
R958 VDD2.n174 VDD2.n99 12.8005
R959 VDD2.n169 VDD2.n101 12.8005
R960 VDD2.n126 VDD2.n122 12.8005
R961 VDD2.n32 VDD2.n28 12.8005
R962 VDD2.n76 VDD2.n8 12.8005
R963 VDD2.n81 VDD2.n6 12.8005
R964 VDD2.n175 VDD2.n97 12.0247
R965 VDD2.n166 VDD2.n165 12.0247
R966 VDD2.n130 VDD2.n129 12.0247
R967 VDD2.n36 VDD2.n35 12.0247
R968 VDD2.n73 VDD2.n72 12.0247
R969 VDD2.n82 VDD2.n4 12.0247
R970 VDD2.n179 VDD2.n178 11.249
R971 VDD2.n162 VDD2.n103 11.249
R972 VDD2.n133 VDD2.n120 11.249
R973 VDD2.n39 VDD2.n26 11.249
R974 VDD2.n68 VDD2.n10 11.249
R975 VDD2.n86 VDD2.n85 11.249
R976 VDD2.n182 VDD2.n95 10.4732
R977 VDD2.n161 VDD2.n106 10.4732
R978 VDD2.n134 VDD2.n118 10.4732
R979 VDD2.n40 VDD2.n24 10.4732
R980 VDD2.n67 VDD2.n12 10.4732
R981 VDD2.n89 VDD2.n2 10.4732
R982 VDD2.n183 VDD2.n93 9.69747
R983 VDD2.n158 VDD2.n157 9.69747
R984 VDD2.n138 VDD2.n137 9.69747
R985 VDD2.n44 VDD2.n43 9.69747
R986 VDD2.n64 VDD2.n63 9.69747
R987 VDD2.n90 VDD2.n0 9.69747
R988 VDD2.n185 VDD2.n184 9.45567
R989 VDD2.n92 VDD2.n91 9.45567
R990 VDD2.n151 VDD2.n150 9.3005
R991 VDD2.n153 VDD2.n152 9.3005
R992 VDD2.n108 VDD2.n107 9.3005
R993 VDD2.n159 VDD2.n158 9.3005
R994 VDD2.n161 VDD2.n160 9.3005
R995 VDD2.n103 VDD2.n102 9.3005
R996 VDD2.n167 VDD2.n166 9.3005
R997 VDD2.n169 VDD2.n168 9.3005
R998 VDD2.n184 VDD2.n183 9.3005
R999 VDD2.n95 VDD2.n94 9.3005
R1000 VDD2.n178 VDD2.n177 9.3005
R1001 VDD2.n176 VDD2.n175 9.3005
R1002 VDD2.n99 VDD2.n98 9.3005
R1003 VDD2.n112 VDD2.n111 9.3005
R1004 VDD2.n145 VDD2.n144 9.3005
R1005 VDD2.n143 VDD2.n142 9.3005
R1006 VDD2.n116 VDD2.n115 9.3005
R1007 VDD2.n137 VDD2.n136 9.3005
R1008 VDD2.n135 VDD2.n134 9.3005
R1009 VDD2.n120 VDD2.n119 9.3005
R1010 VDD2.n129 VDD2.n128 9.3005
R1011 VDD2.n127 VDD2.n126 9.3005
R1012 VDD2.n91 VDD2.n90 9.3005
R1013 VDD2.n2 VDD2.n1 9.3005
R1014 VDD2.n85 VDD2.n84 9.3005
R1015 VDD2.n83 VDD2.n82 9.3005
R1016 VDD2.n6 VDD2.n5 9.3005
R1017 VDD2.n51 VDD2.n50 9.3005
R1018 VDD2.n49 VDD2.n48 9.3005
R1019 VDD2.n22 VDD2.n21 9.3005
R1020 VDD2.n43 VDD2.n42 9.3005
R1021 VDD2.n41 VDD2.n40 9.3005
R1022 VDD2.n26 VDD2.n25 9.3005
R1023 VDD2.n35 VDD2.n34 9.3005
R1024 VDD2.n33 VDD2.n32 9.3005
R1025 VDD2.n18 VDD2.n17 9.3005
R1026 VDD2.n57 VDD2.n56 9.3005
R1027 VDD2.n59 VDD2.n58 9.3005
R1028 VDD2.n14 VDD2.n13 9.3005
R1029 VDD2.n65 VDD2.n64 9.3005
R1030 VDD2.n67 VDD2.n66 9.3005
R1031 VDD2.n10 VDD2.n9 9.3005
R1032 VDD2.n74 VDD2.n73 9.3005
R1033 VDD2.n76 VDD2.n75 9.3005
R1034 VDD2.n154 VDD2.n108 8.92171
R1035 VDD2.n141 VDD2.n116 8.92171
R1036 VDD2.n47 VDD2.n22 8.92171
R1037 VDD2.n60 VDD2.n14 8.92171
R1038 VDD2.n153 VDD2.n110 8.14595
R1039 VDD2.n142 VDD2.n114 8.14595
R1040 VDD2.n48 VDD2.n20 8.14595
R1041 VDD2.n59 VDD2.n16 8.14595
R1042 VDD2.n150 VDD2.n149 7.3702
R1043 VDD2.n146 VDD2.n145 7.3702
R1044 VDD2.n52 VDD2.n51 7.3702
R1045 VDD2.n56 VDD2.n55 7.3702
R1046 VDD2.n149 VDD2.n112 6.59444
R1047 VDD2.n146 VDD2.n112 6.59444
R1048 VDD2.n52 VDD2.n18 6.59444
R1049 VDD2.n55 VDD2.n18 6.59444
R1050 VDD2.n150 VDD2.n110 5.81868
R1051 VDD2.n145 VDD2.n114 5.81868
R1052 VDD2.n51 VDD2.n20 5.81868
R1053 VDD2.n56 VDD2.n16 5.81868
R1054 VDD2.n154 VDD2.n153 5.04292
R1055 VDD2.n142 VDD2.n141 5.04292
R1056 VDD2.n48 VDD2.n47 5.04292
R1057 VDD2.n60 VDD2.n59 5.04292
R1058 VDD2.n185 VDD2.n93 4.26717
R1059 VDD2.n157 VDD2.n108 4.26717
R1060 VDD2.n138 VDD2.n116 4.26717
R1061 VDD2.n44 VDD2.n22 4.26717
R1062 VDD2.n63 VDD2.n14 4.26717
R1063 VDD2.n92 VDD2.n0 4.26717
R1064 VDD2.n127 VDD2.n123 3.70982
R1065 VDD2.n33 VDD2.n29 3.70982
R1066 VDD2.n183 VDD2.n182 3.49141
R1067 VDD2.n158 VDD2.n106 3.49141
R1068 VDD2.n137 VDD2.n118 3.49141
R1069 VDD2.n43 VDD2.n24 3.49141
R1070 VDD2.n64 VDD2.n12 3.49141
R1071 VDD2.n90 VDD2.n89 3.49141
R1072 VDD2.n179 VDD2.n95 2.71565
R1073 VDD2.n162 VDD2.n161 2.71565
R1074 VDD2.n134 VDD2.n133 2.71565
R1075 VDD2.n40 VDD2.n39 2.71565
R1076 VDD2.n68 VDD2.n67 2.71565
R1077 VDD2.n86 VDD2.n2 2.71565
R1078 VDD2.n178 VDD2.n97 1.93989
R1079 VDD2.n165 VDD2.n103 1.93989
R1080 VDD2.n130 VDD2.n120 1.93989
R1081 VDD2.n36 VDD2.n26 1.93989
R1082 VDD2.n72 VDD2.n10 1.93989
R1083 VDD2.n85 VDD2.n4 1.93989
R1084 VDD2.n175 VDD2.n174 1.16414
R1085 VDD2.n166 VDD2.n101 1.16414
R1086 VDD2.n129 VDD2.n122 1.16414
R1087 VDD2.n35 VDD2.n28 1.16414
R1088 VDD2.n73 VDD2.n8 1.16414
R1089 VDD2.n82 VDD2.n81 1.16414
R1090 VDD2.n171 VDD2.n99 0.388379
R1091 VDD2.n170 VDD2.n169 0.388379
R1092 VDD2.n126 VDD2.n125 0.388379
R1093 VDD2.n32 VDD2.n31 0.388379
R1094 VDD2.n77 VDD2.n76 0.388379
R1095 VDD2.n78 VDD2.n6 0.388379
R1096 VDD2 VDD2.n186 0.341017
R1097 VDD2.n184 VDD2.n94 0.155672
R1098 VDD2.n177 VDD2.n94 0.155672
R1099 VDD2.n177 VDD2.n176 0.155672
R1100 VDD2.n176 VDD2.n98 0.155672
R1101 VDD2.n168 VDD2.n98 0.155672
R1102 VDD2.n168 VDD2.n167 0.155672
R1103 VDD2.n167 VDD2.n102 0.155672
R1104 VDD2.n160 VDD2.n102 0.155672
R1105 VDD2.n160 VDD2.n159 0.155672
R1106 VDD2.n159 VDD2.n107 0.155672
R1107 VDD2.n152 VDD2.n107 0.155672
R1108 VDD2.n152 VDD2.n151 0.155672
R1109 VDD2.n151 VDD2.n111 0.155672
R1110 VDD2.n144 VDD2.n111 0.155672
R1111 VDD2.n144 VDD2.n143 0.155672
R1112 VDD2.n143 VDD2.n115 0.155672
R1113 VDD2.n136 VDD2.n115 0.155672
R1114 VDD2.n136 VDD2.n135 0.155672
R1115 VDD2.n135 VDD2.n119 0.155672
R1116 VDD2.n128 VDD2.n119 0.155672
R1117 VDD2.n128 VDD2.n127 0.155672
R1118 VDD2.n34 VDD2.n33 0.155672
R1119 VDD2.n34 VDD2.n25 0.155672
R1120 VDD2.n41 VDD2.n25 0.155672
R1121 VDD2.n42 VDD2.n41 0.155672
R1122 VDD2.n42 VDD2.n21 0.155672
R1123 VDD2.n49 VDD2.n21 0.155672
R1124 VDD2.n50 VDD2.n49 0.155672
R1125 VDD2.n50 VDD2.n17 0.155672
R1126 VDD2.n57 VDD2.n17 0.155672
R1127 VDD2.n58 VDD2.n57 0.155672
R1128 VDD2.n58 VDD2.n13 0.155672
R1129 VDD2.n65 VDD2.n13 0.155672
R1130 VDD2.n66 VDD2.n65 0.155672
R1131 VDD2.n66 VDD2.n9 0.155672
R1132 VDD2.n74 VDD2.n9 0.155672
R1133 VDD2.n75 VDD2.n74 0.155672
R1134 VDD2.n75 VDD2.n5 0.155672
R1135 VDD2.n83 VDD2.n5 0.155672
R1136 VDD2.n84 VDD2.n83 0.155672
R1137 VDD2.n84 VDD2.n1 0.155672
R1138 VDD2.n91 VDD2.n1 0.155672
R1139 B.n120 B.t0 618.39
R1140 B.n128 B.t3 618.39
R1141 B.n38 B.t9 618.39
R1142 B.n46 B.t6 618.39
R1143 B.n422 B.n75 585
R1144 B.n424 B.n423 585
R1145 B.n425 B.n74 585
R1146 B.n427 B.n426 585
R1147 B.n428 B.n73 585
R1148 B.n430 B.n429 585
R1149 B.n431 B.n72 585
R1150 B.n433 B.n432 585
R1151 B.n434 B.n71 585
R1152 B.n436 B.n435 585
R1153 B.n437 B.n70 585
R1154 B.n439 B.n438 585
R1155 B.n440 B.n69 585
R1156 B.n442 B.n441 585
R1157 B.n443 B.n68 585
R1158 B.n445 B.n444 585
R1159 B.n446 B.n67 585
R1160 B.n448 B.n447 585
R1161 B.n449 B.n66 585
R1162 B.n451 B.n450 585
R1163 B.n452 B.n65 585
R1164 B.n454 B.n453 585
R1165 B.n455 B.n64 585
R1166 B.n457 B.n456 585
R1167 B.n458 B.n63 585
R1168 B.n460 B.n459 585
R1169 B.n461 B.n62 585
R1170 B.n463 B.n462 585
R1171 B.n464 B.n61 585
R1172 B.n466 B.n465 585
R1173 B.n467 B.n60 585
R1174 B.n469 B.n468 585
R1175 B.n470 B.n59 585
R1176 B.n472 B.n471 585
R1177 B.n473 B.n58 585
R1178 B.n475 B.n474 585
R1179 B.n476 B.n57 585
R1180 B.n478 B.n477 585
R1181 B.n479 B.n56 585
R1182 B.n481 B.n480 585
R1183 B.n482 B.n55 585
R1184 B.n484 B.n483 585
R1185 B.n485 B.n54 585
R1186 B.n487 B.n486 585
R1187 B.n488 B.n53 585
R1188 B.n490 B.n489 585
R1189 B.n491 B.n52 585
R1190 B.n493 B.n492 585
R1191 B.n494 B.n51 585
R1192 B.n496 B.n495 585
R1193 B.n497 B.n50 585
R1194 B.n499 B.n498 585
R1195 B.n500 B.n49 585
R1196 B.n502 B.n501 585
R1197 B.n503 B.n48 585
R1198 B.n505 B.n504 585
R1199 B.n507 B.n45 585
R1200 B.n509 B.n508 585
R1201 B.n510 B.n44 585
R1202 B.n512 B.n511 585
R1203 B.n513 B.n43 585
R1204 B.n515 B.n514 585
R1205 B.n516 B.n42 585
R1206 B.n518 B.n517 585
R1207 B.n519 B.n41 585
R1208 B.n521 B.n520 585
R1209 B.n523 B.n522 585
R1210 B.n524 B.n37 585
R1211 B.n526 B.n525 585
R1212 B.n527 B.n36 585
R1213 B.n529 B.n528 585
R1214 B.n530 B.n35 585
R1215 B.n532 B.n531 585
R1216 B.n533 B.n34 585
R1217 B.n535 B.n534 585
R1218 B.n536 B.n33 585
R1219 B.n538 B.n537 585
R1220 B.n539 B.n32 585
R1221 B.n541 B.n540 585
R1222 B.n542 B.n31 585
R1223 B.n544 B.n543 585
R1224 B.n545 B.n30 585
R1225 B.n547 B.n546 585
R1226 B.n548 B.n29 585
R1227 B.n550 B.n549 585
R1228 B.n551 B.n28 585
R1229 B.n553 B.n552 585
R1230 B.n554 B.n27 585
R1231 B.n556 B.n555 585
R1232 B.n557 B.n26 585
R1233 B.n559 B.n558 585
R1234 B.n560 B.n25 585
R1235 B.n562 B.n561 585
R1236 B.n563 B.n24 585
R1237 B.n565 B.n564 585
R1238 B.n566 B.n23 585
R1239 B.n568 B.n567 585
R1240 B.n569 B.n22 585
R1241 B.n571 B.n570 585
R1242 B.n572 B.n21 585
R1243 B.n574 B.n573 585
R1244 B.n575 B.n20 585
R1245 B.n577 B.n576 585
R1246 B.n578 B.n19 585
R1247 B.n580 B.n579 585
R1248 B.n581 B.n18 585
R1249 B.n583 B.n582 585
R1250 B.n584 B.n17 585
R1251 B.n586 B.n585 585
R1252 B.n587 B.n16 585
R1253 B.n589 B.n588 585
R1254 B.n590 B.n15 585
R1255 B.n592 B.n591 585
R1256 B.n593 B.n14 585
R1257 B.n595 B.n594 585
R1258 B.n596 B.n13 585
R1259 B.n598 B.n597 585
R1260 B.n599 B.n12 585
R1261 B.n601 B.n600 585
R1262 B.n602 B.n11 585
R1263 B.n604 B.n603 585
R1264 B.n605 B.n10 585
R1265 B.n421 B.n420 585
R1266 B.n419 B.n76 585
R1267 B.n418 B.n417 585
R1268 B.n416 B.n77 585
R1269 B.n415 B.n414 585
R1270 B.n413 B.n78 585
R1271 B.n412 B.n411 585
R1272 B.n410 B.n79 585
R1273 B.n409 B.n408 585
R1274 B.n407 B.n80 585
R1275 B.n406 B.n405 585
R1276 B.n404 B.n81 585
R1277 B.n403 B.n402 585
R1278 B.n401 B.n82 585
R1279 B.n400 B.n399 585
R1280 B.n398 B.n83 585
R1281 B.n397 B.n396 585
R1282 B.n395 B.n84 585
R1283 B.n394 B.n393 585
R1284 B.n392 B.n85 585
R1285 B.n391 B.n390 585
R1286 B.n389 B.n86 585
R1287 B.n388 B.n387 585
R1288 B.n386 B.n87 585
R1289 B.n385 B.n384 585
R1290 B.n383 B.n88 585
R1291 B.n382 B.n381 585
R1292 B.n380 B.n89 585
R1293 B.n379 B.n378 585
R1294 B.n377 B.n90 585
R1295 B.n376 B.n375 585
R1296 B.n374 B.n91 585
R1297 B.n373 B.n372 585
R1298 B.n188 B.n157 585
R1299 B.n190 B.n189 585
R1300 B.n191 B.n156 585
R1301 B.n193 B.n192 585
R1302 B.n194 B.n155 585
R1303 B.n196 B.n195 585
R1304 B.n197 B.n154 585
R1305 B.n199 B.n198 585
R1306 B.n200 B.n153 585
R1307 B.n202 B.n201 585
R1308 B.n203 B.n152 585
R1309 B.n205 B.n204 585
R1310 B.n206 B.n151 585
R1311 B.n208 B.n207 585
R1312 B.n209 B.n150 585
R1313 B.n211 B.n210 585
R1314 B.n212 B.n149 585
R1315 B.n214 B.n213 585
R1316 B.n215 B.n148 585
R1317 B.n217 B.n216 585
R1318 B.n218 B.n147 585
R1319 B.n220 B.n219 585
R1320 B.n221 B.n146 585
R1321 B.n223 B.n222 585
R1322 B.n224 B.n145 585
R1323 B.n226 B.n225 585
R1324 B.n227 B.n144 585
R1325 B.n229 B.n228 585
R1326 B.n230 B.n143 585
R1327 B.n232 B.n231 585
R1328 B.n233 B.n142 585
R1329 B.n235 B.n234 585
R1330 B.n236 B.n141 585
R1331 B.n238 B.n237 585
R1332 B.n239 B.n140 585
R1333 B.n241 B.n240 585
R1334 B.n242 B.n139 585
R1335 B.n244 B.n243 585
R1336 B.n245 B.n138 585
R1337 B.n247 B.n246 585
R1338 B.n248 B.n137 585
R1339 B.n250 B.n249 585
R1340 B.n251 B.n136 585
R1341 B.n253 B.n252 585
R1342 B.n254 B.n135 585
R1343 B.n256 B.n255 585
R1344 B.n257 B.n134 585
R1345 B.n259 B.n258 585
R1346 B.n260 B.n133 585
R1347 B.n262 B.n261 585
R1348 B.n263 B.n132 585
R1349 B.n265 B.n264 585
R1350 B.n266 B.n131 585
R1351 B.n268 B.n267 585
R1352 B.n269 B.n130 585
R1353 B.n271 B.n270 585
R1354 B.n273 B.n127 585
R1355 B.n275 B.n274 585
R1356 B.n276 B.n126 585
R1357 B.n278 B.n277 585
R1358 B.n279 B.n125 585
R1359 B.n281 B.n280 585
R1360 B.n282 B.n124 585
R1361 B.n284 B.n283 585
R1362 B.n285 B.n123 585
R1363 B.n287 B.n286 585
R1364 B.n289 B.n288 585
R1365 B.n290 B.n119 585
R1366 B.n292 B.n291 585
R1367 B.n293 B.n118 585
R1368 B.n295 B.n294 585
R1369 B.n296 B.n117 585
R1370 B.n298 B.n297 585
R1371 B.n299 B.n116 585
R1372 B.n301 B.n300 585
R1373 B.n302 B.n115 585
R1374 B.n304 B.n303 585
R1375 B.n305 B.n114 585
R1376 B.n307 B.n306 585
R1377 B.n308 B.n113 585
R1378 B.n310 B.n309 585
R1379 B.n311 B.n112 585
R1380 B.n313 B.n312 585
R1381 B.n314 B.n111 585
R1382 B.n316 B.n315 585
R1383 B.n317 B.n110 585
R1384 B.n319 B.n318 585
R1385 B.n320 B.n109 585
R1386 B.n322 B.n321 585
R1387 B.n323 B.n108 585
R1388 B.n325 B.n324 585
R1389 B.n326 B.n107 585
R1390 B.n328 B.n327 585
R1391 B.n329 B.n106 585
R1392 B.n331 B.n330 585
R1393 B.n332 B.n105 585
R1394 B.n334 B.n333 585
R1395 B.n335 B.n104 585
R1396 B.n337 B.n336 585
R1397 B.n338 B.n103 585
R1398 B.n340 B.n339 585
R1399 B.n341 B.n102 585
R1400 B.n343 B.n342 585
R1401 B.n344 B.n101 585
R1402 B.n346 B.n345 585
R1403 B.n347 B.n100 585
R1404 B.n349 B.n348 585
R1405 B.n350 B.n99 585
R1406 B.n352 B.n351 585
R1407 B.n353 B.n98 585
R1408 B.n355 B.n354 585
R1409 B.n356 B.n97 585
R1410 B.n358 B.n357 585
R1411 B.n359 B.n96 585
R1412 B.n361 B.n360 585
R1413 B.n362 B.n95 585
R1414 B.n364 B.n363 585
R1415 B.n365 B.n94 585
R1416 B.n367 B.n366 585
R1417 B.n368 B.n93 585
R1418 B.n370 B.n369 585
R1419 B.n371 B.n92 585
R1420 B.n187 B.n186 585
R1421 B.n185 B.n158 585
R1422 B.n184 B.n183 585
R1423 B.n182 B.n159 585
R1424 B.n181 B.n180 585
R1425 B.n179 B.n160 585
R1426 B.n178 B.n177 585
R1427 B.n176 B.n161 585
R1428 B.n175 B.n174 585
R1429 B.n173 B.n162 585
R1430 B.n172 B.n171 585
R1431 B.n170 B.n163 585
R1432 B.n169 B.n168 585
R1433 B.n167 B.n164 585
R1434 B.n166 B.n165 585
R1435 B.n2 B.n0 585
R1436 B.n629 B.n1 585
R1437 B.n628 B.n627 585
R1438 B.n626 B.n3 585
R1439 B.n625 B.n624 585
R1440 B.n623 B.n4 585
R1441 B.n622 B.n621 585
R1442 B.n620 B.n5 585
R1443 B.n619 B.n618 585
R1444 B.n617 B.n6 585
R1445 B.n616 B.n615 585
R1446 B.n614 B.n7 585
R1447 B.n613 B.n612 585
R1448 B.n611 B.n8 585
R1449 B.n610 B.n609 585
R1450 B.n608 B.n9 585
R1451 B.n607 B.n606 585
R1452 B.n631 B.n630 585
R1453 B.n120 B.t2 489.387
R1454 B.n46 B.t7 489.387
R1455 B.n128 B.t5 489.387
R1456 B.n38 B.t10 489.387
R1457 B.n121 B.t1 463.981
R1458 B.n47 B.t8 463.981
R1459 B.n129 B.t4 463.981
R1460 B.n39 B.t11 463.981
R1461 B.n186 B.n157 449.257
R1462 B.n606 B.n605 449.257
R1463 B.n372 B.n371 449.257
R1464 B.n420 B.n75 449.257
R1465 B.n186 B.n185 163.367
R1466 B.n185 B.n184 163.367
R1467 B.n184 B.n159 163.367
R1468 B.n180 B.n159 163.367
R1469 B.n180 B.n179 163.367
R1470 B.n179 B.n178 163.367
R1471 B.n178 B.n161 163.367
R1472 B.n174 B.n161 163.367
R1473 B.n174 B.n173 163.367
R1474 B.n173 B.n172 163.367
R1475 B.n172 B.n163 163.367
R1476 B.n168 B.n163 163.367
R1477 B.n168 B.n167 163.367
R1478 B.n167 B.n166 163.367
R1479 B.n166 B.n2 163.367
R1480 B.n630 B.n2 163.367
R1481 B.n630 B.n629 163.367
R1482 B.n629 B.n628 163.367
R1483 B.n628 B.n3 163.367
R1484 B.n624 B.n3 163.367
R1485 B.n624 B.n623 163.367
R1486 B.n623 B.n622 163.367
R1487 B.n622 B.n5 163.367
R1488 B.n618 B.n5 163.367
R1489 B.n618 B.n617 163.367
R1490 B.n617 B.n616 163.367
R1491 B.n616 B.n7 163.367
R1492 B.n612 B.n7 163.367
R1493 B.n612 B.n611 163.367
R1494 B.n611 B.n610 163.367
R1495 B.n610 B.n9 163.367
R1496 B.n606 B.n9 163.367
R1497 B.n190 B.n157 163.367
R1498 B.n191 B.n190 163.367
R1499 B.n192 B.n191 163.367
R1500 B.n192 B.n155 163.367
R1501 B.n196 B.n155 163.367
R1502 B.n197 B.n196 163.367
R1503 B.n198 B.n197 163.367
R1504 B.n198 B.n153 163.367
R1505 B.n202 B.n153 163.367
R1506 B.n203 B.n202 163.367
R1507 B.n204 B.n203 163.367
R1508 B.n204 B.n151 163.367
R1509 B.n208 B.n151 163.367
R1510 B.n209 B.n208 163.367
R1511 B.n210 B.n209 163.367
R1512 B.n210 B.n149 163.367
R1513 B.n214 B.n149 163.367
R1514 B.n215 B.n214 163.367
R1515 B.n216 B.n215 163.367
R1516 B.n216 B.n147 163.367
R1517 B.n220 B.n147 163.367
R1518 B.n221 B.n220 163.367
R1519 B.n222 B.n221 163.367
R1520 B.n222 B.n145 163.367
R1521 B.n226 B.n145 163.367
R1522 B.n227 B.n226 163.367
R1523 B.n228 B.n227 163.367
R1524 B.n228 B.n143 163.367
R1525 B.n232 B.n143 163.367
R1526 B.n233 B.n232 163.367
R1527 B.n234 B.n233 163.367
R1528 B.n234 B.n141 163.367
R1529 B.n238 B.n141 163.367
R1530 B.n239 B.n238 163.367
R1531 B.n240 B.n239 163.367
R1532 B.n240 B.n139 163.367
R1533 B.n244 B.n139 163.367
R1534 B.n245 B.n244 163.367
R1535 B.n246 B.n245 163.367
R1536 B.n246 B.n137 163.367
R1537 B.n250 B.n137 163.367
R1538 B.n251 B.n250 163.367
R1539 B.n252 B.n251 163.367
R1540 B.n252 B.n135 163.367
R1541 B.n256 B.n135 163.367
R1542 B.n257 B.n256 163.367
R1543 B.n258 B.n257 163.367
R1544 B.n258 B.n133 163.367
R1545 B.n262 B.n133 163.367
R1546 B.n263 B.n262 163.367
R1547 B.n264 B.n263 163.367
R1548 B.n264 B.n131 163.367
R1549 B.n268 B.n131 163.367
R1550 B.n269 B.n268 163.367
R1551 B.n270 B.n269 163.367
R1552 B.n270 B.n127 163.367
R1553 B.n275 B.n127 163.367
R1554 B.n276 B.n275 163.367
R1555 B.n277 B.n276 163.367
R1556 B.n277 B.n125 163.367
R1557 B.n281 B.n125 163.367
R1558 B.n282 B.n281 163.367
R1559 B.n283 B.n282 163.367
R1560 B.n283 B.n123 163.367
R1561 B.n287 B.n123 163.367
R1562 B.n288 B.n287 163.367
R1563 B.n288 B.n119 163.367
R1564 B.n292 B.n119 163.367
R1565 B.n293 B.n292 163.367
R1566 B.n294 B.n293 163.367
R1567 B.n294 B.n117 163.367
R1568 B.n298 B.n117 163.367
R1569 B.n299 B.n298 163.367
R1570 B.n300 B.n299 163.367
R1571 B.n300 B.n115 163.367
R1572 B.n304 B.n115 163.367
R1573 B.n305 B.n304 163.367
R1574 B.n306 B.n305 163.367
R1575 B.n306 B.n113 163.367
R1576 B.n310 B.n113 163.367
R1577 B.n311 B.n310 163.367
R1578 B.n312 B.n311 163.367
R1579 B.n312 B.n111 163.367
R1580 B.n316 B.n111 163.367
R1581 B.n317 B.n316 163.367
R1582 B.n318 B.n317 163.367
R1583 B.n318 B.n109 163.367
R1584 B.n322 B.n109 163.367
R1585 B.n323 B.n322 163.367
R1586 B.n324 B.n323 163.367
R1587 B.n324 B.n107 163.367
R1588 B.n328 B.n107 163.367
R1589 B.n329 B.n328 163.367
R1590 B.n330 B.n329 163.367
R1591 B.n330 B.n105 163.367
R1592 B.n334 B.n105 163.367
R1593 B.n335 B.n334 163.367
R1594 B.n336 B.n335 163.367
R1595 B.n336 B.n103 163.367
R1596 B.n340 B.n103 163.367
R1597 B.n341 B.n340 163.367
R1598 B.n342 B.n341 163.367
R1599 B.n342 B.n101 163.367
R1600 B.n346 B.n101 163.367
R1601 B.n347 B.n346 163.367
R1602 B.n348 B.n347 163.367
R1603 B.n348 B.n99 163.367
R1604 B.n352 B.n99 163.367
R1605 B.n353 B.n352 163.367
R1606 B.n354 B.n353 163.367
R1607 B.n354 B.n97 163.367
R1608 B.n358 B.n97 163.367
R1609 B.n359 B.n358 163.367
R1610 B.n360 B.n359 163.367
R1611 B.n360 B.n95 163.367
R1612 B.n364 B.n95 163.367
R1613 B.n365 B.n364 163.367
R1614 B.n366 B.n365 163.367
R1615 B.n366 B.n93 163.367
R1616 B.n370 B.n93 163.367
R1617 B.n371 B.n370 163.367
R1618 B.n372 B.n91 163.367
R1619 B.n376 B.n91 163.367
R1620 B.n377 B.n376 163.367
R1621 B.n378 B.n377 163.367
R1622 B.n378 B.n89 163.367
R1623 B.n382 B.n89 163.367
R1624 B.n383 B.n382 163.367
R1625 B.n384 B.n383 163.367
R1626 B.n384 B.n87 163.367
R1627 B.n388 B.n87 163.367
R1628 B.n389 B.n388 163.367
R1629 B.n390 B.n389 163.367
R1630 B.n390 B.n85 163.367
R1631 B.n394 B.n85 163.367
R1632 B.n395 B.n394 163.367
R1633 B.n396 B.n395 163.367
R1634 B.n396 B.n83 163.367
R1635 B.n400 B.n83 163.367
R1636 B.n401 B.n400 163.367
R1637 B.n402 B.n401 163.367
R1638 B.n402 B.n81 163.367
R1639 B.n406 B.n81 163.367
R1640 B.n407 B.n406 163.367
R1641 B.n408 B.n407 163.367
R1642 B.n408 B.n79 163.367
R1643 B.n412 B.n79 163.367
R1644 B.n413 B.n412 163.367
R1645 B.n414 B.n413 163.367
R1646 B.n414 B.n77 163.367
R1647 B.n418 B.n77 163.367
R1648 B.n419 B.n418 163.367
R1649 B.n420 B.n419 163.367
R1650 B.n605 B.n604 163.367
R1651 B.n604 B.n11 163.367
R1652 B.n600 B.n11 163.367
R1653 B.n600 B.n599 163.367
R1654 B.n599 B.n598 163.367
R1655 B.n598 B.n13 163.367
R1656 B.n594 B.n13 163.367
R1657 B.n594 B.n593 163.367
R1658 B.n593 B.n592 163.367
R1659 B.n592 B.n15 163.367
R1660 B.n588 B.n15 163.367
R1661 B.n588 B.n587 163.367
R1662 B.n587 B.n586 163.367
R1663 B.n586 B.n17 163.367
R1664 B.n582 B.n17 163.367
R1665 B.n582 B.n581 163.367
R1666 B.n581 B.n580 163.367
R1667 B.n580 B.n19 163.367
R1668 B.n576 B.n19 163.367
R1669 B.n576 B.n575 163.367
R1670 B.n575 B.n574 163.367
R1671 B.n574 B.n21 163.367
R1672 B.n570 B.n21 163.367
R1673 B.n570 B.n569 163.367
R1674 B.n569 B.n568 163.367
R1675 B.n568 B.n23 163.367
R1676 B.n564 B.n23 163.367
R1677 B.n564 B.n563 163.367
R1678 B.n563 B.n562 163.367
R1679 B.n562 B.n25 163.367
R1680 B.n558 B.n25 163.367
R1681 B.n558 B.n557 163.367
R1682 B.n557 B.n556 163.367
R1683 B.n556 B.n27 163.367
R1684 B.n552 B.n27 163.367
R1685 B.n552 B.n551 163.367
R1686 B.n551 B.n550 163.367
R1687 B.n550 B.n29 163.367
R1688 B.n546 B.n29 163.367
R1689 B.n546 B.n545 163.367
R1690 B.n545 B.n544 163.367
R1691 B.n544 B.n31 163.367
R1692 B.n540 B.n31 163.367
R1693 B.n540 B.n539 163.367
R1694 B.n539 B.n538 163.367
R1695 B.n538 B.n33 163.367
R1696 B.n534 B.n33 163.367
R1697 B.n534 B.n533 163.367
R1698 B.n533 B.n532 163.367
R1699 B.n532 B.n35 163.367
R1700 B.n528 B.n35 163.367
R1701 B.n528 B.n527 163.367
R1702 B.n527 B.n526 163.367
R1703 B.n526 B.n37 163.367
R1704 B.n522 B.n37 163.367
R1705 B.n522 B.n521 163.367
R1706 B.n521 B.n41 163.367
R1707 B.n517 B.n41 163.367
R1708 B.n517 B.n516 163.367
R1709 B.n516 B.n515 163.367
R1710 B.n515 B.n43 163.367
R1711 B.n511 B.n43 163.367
R1712 B.n511 B.n510 163.367
R1713 B.n510 B.n509 163.367
R1714 B.n509 B.n45 163.367
R1715 B.n504 B.n45 163.367
R1716 B.n504 B.n503 163.367
R1717 B.n503 B.n502 163.367
R1718 B.n502 B.n49 163.367
R1719 B.n498 B.n49 163.367
R1720 B.n498 B.n497 163.367
R1721 B.n497 B.n496 163.367
R1722 B.n496 B.n51 163.367
R1723 B.n492 B.n51 163.367
R1724 B.n492 B.n491 163.367
R1725 B.n491 B.n490 163.367
R1726 B.n490 B.n53 163.367
R1727 B.n486 B.n53 163.367
R1728 B.n486 B.n485 163.367
R1729 B.n485 B.n484 163.367
R1730 B.n484 B.n55 163.367
R1731 B.n480 B.n55 163.367
R1732 B.n480 B.n479 163.367
R1733 B.n479 B.n478 163.367
R1734 B.n478 B.n57 163.367
R1735 B.n474 B.n57 163.367
R1736 B.n474 B.n473 163.367
R1737 B.n473 B.n472 163.367
R1738 B.n472 B.n59 163.367
R1739 B.n468 B.n59 163.367
R1740 B.n468 B.n467 163.367
R1741 B.n467 B.n466 163.367
R1742 B.n466 B.n61 163.367
R1743 B.n462 B.n61 163.367
R1744 B.n462 B.n461 163.367
R1745 B.n461 B.n460 163.367
R1746 B.n460 B.n63 163.367
R1747 B.n456 B.n63 163.367
R1748 B.n456 B.n455 163.367
R1749 B.n455 B.n454 163.367
R1750 B.n454 B.n65 163.367
R1751 B.n450 B.n65 163.367
R1752 B.n450 B.n449 163.367
R1753 B.n449 B.n448 163.367
R1754 B.n448 B.n67 163.367
R1755 B.n444 B.n67 163.367
R1756 B.n444 B.n443 163.367
R1757 B.n443 B.n442 163.367
R1758 B.n442 B.n69 163.367
R1759 B.n438 B.n69 163.367
R1760 B.n438 B.n437 163.367
R1761 B.n437 B.n436 163.367
R1762 B.n436 B.n71 163.367
R1763 B.n432 B.n71 163.367
R1764 B.n432 B.n431 163.367
R1765 B.n431 B.n430 163.367
R1766 B.n430 B.n73 163.367
R1767 B.n426 B.n73 163.367
R1768 B.n426 B.n425 163.367
R1769 B.n425 B.n424 163.367
R1770 B.n424 B.n75 163.367
R1771 B.n122 B.n121 59.5399
R1772 B.n272 B.n129 59.5399
R1773 B.n40 B.n39 59.5399
R1774 B.n506 B.n47 59.5399
R1775 B.n607 B.n10 29.1907
R1776 B.n373 B.n92 29.1907
R1777 B.n188 B.n187 29.1907
R1778 B.n422 B.n421 29.1907
R1779 B.n121 B.n120 25.4066
R1780 B.n129 B.n128 25.4066
R1781 B.n39 B.n38 25.4066
R1782 B.n47 B.n46 25.4066
R1783 B B.n631 18.0485
R1784 B.n603 B.n10 10.6151
R1785 B.n603 B.n602 10.6151
R1786 B.n602 B.n601 10.6151
R1787 B.n601 B.n12 10.6151
R1788 B.n597 B.n12 10.6151
R1789 B.n597 B.n596 10.6151
R1790 B.n596 B.n595 10.6151
R1791 B.n595 B.n14 10.6151
R1792 B.n591 B.n14 10.6151
R1793 B.n591 B.n590 10.6151
R1794 B.n590 B.n589 10.6151
R1795 B.n589 B.n16 10.6151
R1796 B.n585 B.n16 10.6151
R1797 B.n585 B.n584 10.6151
R1798 B.n584 B.n583 10.6151
R1799 B.n583 B.n18 10.6151
R1800 B.n579 B.n18 10.6151
R1801 B.n579 B.n578 10.6151
R1802 B.n578 B.n577 10.6151
R1803 B.n577 B.n20 10.6151
R1804 B.n573 B.n20 10.6151
R1805 B.n573 B.n572 10.6151
R1806 B.n572 B.n571 10.6151
R1807 B.n571 B.n22 10.6151
R1808 B.n567 B.n22 10.6151
R1809 B.n567 B.n566 10.6151
R1810 B.n566 B.n565 10.6151
R1811 B.n565 B.n24 10.6151
R1812 B.n561 B.n24 10.6151
R1813 B.n561 B.n560 10.6151
R1814 B.n560 B.n559 10.6151
R1815 B.n559 B.n26 10.6151
R1816 B.n555 B.n26 10.6151
R1817 B.n555 B.n554 10.6151
R1818 B.n554 B.n553 10.6151
R1819 B.n553 B.n28 10.6151
R1820 B.n549 B.n28 10.6151
R1821 B.n549 B.n548 10.6151
R1822 B.n548 B.n547 10.6151
R1823 B.n547 B.n30 10.6151
R1824 B.n543 B.n30 10.6151
R1825 B.n543 B.n542 10.6151
R1826 B.n542 B.n541 10.6151
R1827 B.n541 B.n32 10.6151
R1828 B.n537 B.n32 10.6151
R1829 B.n537 B.n536 10.6151
R1830 B.n536 B.n535 10.6151
R1831 B.n535 B.n34 10.6151
R1832 B.n531 B.n34 10.6151
R1833 B.n531 B.n530 10.6151
R1834 B.n530 B.n529 10.6151
R1835 B.n529 B.n36 10.6151
R1836 B.n525 B.n36 10.6151
R1837 B.n525 B.n524 10.6151
R1838 B.n524 B.n523 10.6151
R1839 B.n520 B.n519 10.6151
R1840 B.n519 B.n518 10.6151
R1841 B.n518 B.n42 10.6151
R1842 B.n514 B.n42 10.6151
R1843 B.n514 B.n513 10.6151
R1844 B.n513 B.n512 10.6151
R1845 B.n512 B.n44 10.6151
R1846 B.n508 B.n44 10.6151
R1847 B.n508 B.n507 10.6151
R1848 B.n505 B.n48 10.6151
R1849 B.n501 B.n48 10.6151
R1850 B.n501 B.n500 10.6151
R1851 B.n500 B.n499 10.6151
R1852 B.n499 B.n50 10.6151
R1853 B.n495 B.n50 10.6151
R1854 B.n495 B.n494 10.6151
R1855 B.n494 B.n493 10.6151
R1856 B.n493 B.n52 10.6151
R1857 B.n489 B.n52 10.6151
R1858 B.n489 B.n488 10.6151
R1859 B.n488 B.n487 10.6151
R1860 B.n487 B.n54 10.6151
R1861 B.n483 B.n54 10.6151
R1862 B.n483 B.n482 10.6151
R1863 B.n482 B.n481 10.6151
R1864 B.n481 B.n56 10.6151
R1865 B.n477 B.n56 10.6151
R1866 B.n477 B.n476 10.6151
R1867 B.n476 B.n475 10.6151
R1868 B.n475 B.n58 10.6151
R1869 B.n471 B.n58 10.6151
R1870 B.n471 B.n470 10.6151
R1871 B.n470 B.n469 10.6151
R1872 B.n469 B.n60 10.6151
R1873 B.n465 B.n60 10.6151
R1874 B.n465 B.n464 10.6151
R1875 B.n464 B.n463 10.6151
R1876 B.n463 B.n62 10.6151
R1877 B.n459 B.n62 10.6151
R1878 B.n459 B.n458 10.6151
R1879 B.n458 B.n457 10.6151
R1880 B.n457 B.n64 10.6151
R1881 B.n453 B.n64 10.6151
R1882 B.n453 B.n452 10.6151
R1883 B.n452 B.n451 10.6151
R1884 B.n451 B.n66 10.6151
R1885 B.n447 B.n66 10.6151
R1886 B.n447 B.n446 10.6151
R1887 B.n446 B.n445 10.6151
R1888 B.n445 B.n68 10.6151
R1889 B.n441 B.n68 10.6151
R1890 B.n441 B.n440 10.6151
R1891 B.n440 B.n439 10.6151
R1892 B.n439 B.n70 10.6151
R1893 B.n435 B.n70 10.6151
R1894 B.n435 B.n434 10.6151
R1895 B.n434 B.n433 10.6151
R1896 B.n433 B.n72 10.6151
R1897 B.n429 B.n72 10.6151
R1898 B.n429 B.n428 10.6151
R1899 B.n428 B.n427 10.6151
R1900 B.n427 B.n74 10.6151
R1901 B.n423 B.n74 10.6151
R1902 B.n423 B.n422 10.6151
R1903 B.n374 B.n373 10.6151
R1904 B.n375 B.n374 10.6151
R1905 B.n375 B.n90 10.6151
R1906 B.n379 B.n90 10.6151
R1907 B.n380 B.n379 10.6151
R1908 B.n381 B.n380 10.6151
R1909 B.n381 B.n88 10.6151
R1910 B.n385 B.n88 10.6151
R1911 B.n386 B.n385 10.6151
R1912 B.n387 B.n386 10.6151
R1913 B.n387 B.n86 10.6151
R1914 B.n391 B.n86 10.6151
R1915 B.n392 B.n391 10.6151
R1916 B.n393 B.n392 10.6151
R1917 B.n393 B.n84 10.6151
R1918 B.n397 B.n84 10.6151
R1919 B.n398 B.n397 10.6151
R1920 B.n399 B.n398 10.6151
R1921 B.n399 B.n82 10.6151
R1922 B.n403 B.n82 10.6151
R1923 B.n404 B.n403 10.6151
R1924 B.n405 B.n404 10.6151
R1925 B.n405 B.n80 10.6151
R1926 B.n409 B.n80 10.6151
R1927 B.n410 B.n409 10.6151
R1928 B.n411 B.n410 10.6151
R1929 B.n411 B.n78 10.6151
R1930 B.n415 B.n78 10.6151
R1931 B.n416 B.n415 10.6151
R1932 B.n417 B.n416 10.6151
R1933 B.n417 B.n76 10.6151
R1934 B.n421 B.n76 10.6151
R1935 B.n189 B.n188 10.6151
R1936 B.n189 B.n156 10.6151
R1937 B.n193 B.n156 10.6151
R1938 B.n194 B.n193 10.6151
R1939 B.n195 B.n194 10.6151
R1940 B.n195 B.n154 10.6151
R1941 B.n199 B.n154 10.6151
R1942 B.n200 B.n199 10.6151
R1943 B.n201 B.n200 10.6151
R1944 B.n201 B.n152 10.6151
R1945 B.n205 B.n152 10.6151
R1946 B.n206 B.n205 10.6151
R1947 B.n207 B.n206 10.6151
R1948 B.n207 B.n150 10.6151
R1949 B.n211 B.n150 10.6151
R1950 B.n212 B.n211 10.6151
R1951 B.n213 B.n212 10.6151
R1952 B.n213 B.n148 10.6151
R1953 B.n217 B.n148 10.6151
R1954 B.n218 B.n217 10.6151
R1955 B.n219 B.n218 10.6151
R1956 B.n219 B.n146 10.6151
R1957 B.n223 B.n146 10.6151
R1958 B.n224 B.n223 10.6151
R1959 B.n225 B.n224 10.6151
R1960 B.n225 B.n144 10.6151
R1961 B.n229 B.n144 10.6151
R1962 B.n230 B.n229 10.6151
R1963 B.n231 B.n230 10.6151
R1964 B.n231 B.n142 10.6151
R1965 B.n235 B.n142 10.6151
R1966 B.n236 B.n235 10.6151
R1967 B.n237 B.n236 10.6151
R1968 B.n237 B.n140 10.6151
R1969 B.n241 B.n140 10.6151
R1970 B.n242 B.n241 10.6151
R1971 B.n243 B.n242 10.6151
R1972 B.n243 B.n138 10.6151
R1973 B.n247 B.n138 10.6151
R1974 B.n248 B.n247 10.6151
R1975 B.n249 B.n248 10.6151
R1976 B.n249 B.n136 10.6151
R1977 B.n253 B.n136 10.6151
R1978 B.n254 B.n253 10.6151
R1979 B.n255 B.n254 10.6151
R1980 B.n255 B.n134 10.6151
R1981 B.n259 B.n134 10.6151
R1982 B.n260 B.n259 10.6151
R1983 B.n261 B.n260 10.6151
R1984 B.n261 B.n132 10.6151
R1985 B.n265 B.n132 10.6151
R1986 B.n266 B.n265 10.6151
R1987 B.n267 B.n266 10.6151
R1988 B.n267 B.n130 10.6151
R1989 B.n271 B.n130 10.6151
R1990 B.n274 B.n273 10.6151
R1991 B.n274 B.n126 10.6151
R1992 B.n278 B.n126 10.6151
R1993 B.n279 B.n278 10.6151
R1994 B.n280 B.n279 10.6151
R1995 B.n280 B.n124 10.6151
R1996 B.n284 B.n124 10.6151
R1997 B.n285 B.n284 10.6151
R1998 B.n286 B.n285 10.6151
R1999 B.n290 B.n289 10.6151
R2000 B.n291 B.n290 10.6151
R2001 B.n291 B.n118 10.6151
R2002 B.n295 B.n118 10.6151
R2003 B.n296 B.n295 10.6151
R2004 B.n297 B.n296 10.6151
R2005 B.n297 B.n116 10.6151
R2006 B.n301 B.n116 10.6151
R2007 B.n302 B.n301 10.6151
R2008 B.n303 B.n302 10.6151
R2009 B.n303 B.n114 10.6151
R2010 B.n307 B.n114 10.6151
R2011 B.n308 B.n307 10.6151
R2012 B.n309 B.n308 10.6151
R2013 B.n309 B.n112 10.6151
R2014 B.n313 B.n112 10.6151
R2015 B.n314 B.n313 10.6151
R2016 B.n315 B.n314 10.6151
R2017 B.n315 B.n110 10.6151
R2018 B.n319 B.n110 10.6151
R2019 B.n320 B.n319 10.6151
R2020 B.n321 B.n320 10.6151
R2021 B.n321 B.n108 10.6151
R2022 B.n325 B.n108 10.6151
R2023 B.n326 B.n325 10.6151
R2024 B.n327 B.n326 10.6151
R2025 B.n327 B.n106 10.6151
R2026 B.n331 B.n106 10.6151
R2027 B.n332 B.n331 10.6151
R2028 B.n333 B.n332 10.6151
R2029 B.n333 B.n104 10.6151
R2030 B.n337 B.n104 10.6151
R2031 B.n338 B.n337 10.6151
R2032 B.n339 B.n338 10.6151
R2033 B.n339 B.n102 10.6151
R2034 B.n343 B.n102 10.6151
R2035 B.n344 B.n343 10.6151
R2036 B.n345 B.n344 10.6151
R2037 B.n345 B.n100 10.6151
R2038 B.n349 B.n100 10.6151
R2039 B.n350 B.n349 10.6151
R2040 B.n351 B.n350 10.6151
R2041 B.n351 B.n98 10.6151
R2042 B.n355 B.n98 10.6151
R2043 B.n356 B.n355 10.6151
R2044 B.n357 B.n356 10.6151
R2045 B.n357 B.n96 10.6151
R2046 B.n361 B.n96 10.6151
R2047 B.n362 B.n361 10.6151
R2048 B.n363 B.n362 10.6151
R2049 B.n363 B.n94 10.6151
R2050 B.n367 B.n94 10.6151
R2051 B.n368 B.n367 10.6151
R2052 B.n369 B.n368 10.6151
R2053 B.n369 B.n92 10.6151
R2054 B.n187 B.n158 10.6151
R2055 B.n183 B.n158 10.6151
R2056 B.n183 B.n182 10.6151
R2057 B.n182 B.n181 10.6151
R2058 B.n181 B.n160 10.6151
R2059 B.n177 B.n160 10.6151
R2060 B.n177 B.n176 10.6151
R2061 B.n176 B.n175 10.6151
R2062 B.n175 B.n162 10.6151
R2063 B.n171 B.n162 10.6151
R2064 B.n171 B.n170 10.6151
R2065 B.n170 B.n169 10.6151
R2066 B.n169 B.n164 10.6151
R2067 B.n165 B.n164 10.6151
R2068 B.n165 B.n0 10.6151
R2069 B.n627 B.n1 10.6151
R2070 B.n627 B.n626 10.6151
R2071 B.n626 B.n625 10.6151
R2072 B.n625 B.n4 10.6151
R2073 B.n621 B.n4 10.6151
R2074 B.n621 B.n620 10.6151
R2075 B.n620 B.n619 10.6151
R2076 B.n619 B.n6 10.6151
R2077 B.n615 B.n6 10.6151
R2078 B.n615 B.n614 10.6151
R2079 B.n614 B.n613 10.6151
R2080 B.n613 B.n8 10.6151
R2081 B.n609 B.n8 10.6151
R2082 B.n609 B.n608 10.6151
R2083 B.n608 B.n607 10.6151
R2084 B.n523 B.n40 8.74196
R2085 B.n506 B.n505 8.74196
R2086 B.n272 B.n271 8.74196
R2087 B.n289 B.n122 8.74196
R2088 B.n631 B.n0 2.81026
R2089 B.n631 B.n1 2.81026
R2090 B.n520 B.n40 1.87367
R2091 B.n507 B.n506 1.87367
R2092 B.n273 B.n272 1.87367
R2093 B.n286 B.n122 1.87367
C0 VDD1 B 1.82827f
C1 B VN 0.83555f
C2 VDD1 w_n1494_n4352# 1.95869f
C3 VTAIL VDD2 6.9826f
C4 VP B 1.13618f
C5 w_n1494_n4352# VN 2.00701f
C6 VP w_n1494_n4352# 2.19382f
C7 VDD2 VDD1 0.491211f
C8 VDD2 VN 3.03308f
C9 VTAIL VDD1 6.94822f
C10 VP VDD2 0.26764f
C11 VTAIL VN 2.3552f
C12 B w_n1494_n4352# 8.436831f
C13 VTAIL VP 2.3699f
C14 VDD1 VN 0.14905f
C15 VDD2 B 1.84477f
C16 VP VDD1 3.14623f
C17 VTAIL B 3.80224f
C18 VDD2 w_n1494_n4352# 1.96615f
C19 VP VN 5.59341f
C20 VTAIL w_n1494_n4352# 3.65507f
C21 VDD2 VSUBS 0.929255f
C22 VDD1 VSUBS 3.7712f
C23 VTAIL VSUBS 0.981953f
C24 VN VSUBS 8.64411f
C25 VP VSUBS 1.378621f
C26 B VSUBS 3.115775f
C27 w_n1494_n4352# VSUBS 79.5824f
C28 B.n0 VSUBS 0.004169f
C29 B.n1 VSUBS 0.004169f
C30 B.n2 VSUBS 0.006593f
C31 B.n3 VSUBS 0.006593f
C32 B.n4 VSUBS 0.006593f
C33 B.n5 VSUBS 0.006593f
C34 B.n6 VSUBS 0.006593f
C35 B.n7 VSUBS 0.006593f
C36 B.n8 VSUBS 0.006593f
C37 B.n9 VSUBS 0.006593f
C38 B.n10 VSUBS 0.014721f
C39 B.n11 VSUBS 0.006593f
C40 B.n12 VSUBS 0.006593f
C41 B.n13 VSUBS 0.006593f
C42 B.n14 VSUBS 0.006593f
C43 B.n15 VSUBS 0.006593f
C44 B.n16 VSUBS 0.006593f
C45 B.n17 VSUBS 0.006593f
C46 B.n18 VSUBS 0.006593f
C47 B.n19 VSUBS 0.006593f
C48 B.n20 VSUBS 0.006593f
C49 B.n21 VSUBS 0.006593f
C50 B.n22 VSUBS 0.006593f
C51 B.n23 VSUBS 0.006593f
C52 B.n24 VSUBS 0.006593f
C53 B.n25 VSUBS 0.006593f
C54 B.n26 VSUBS 0.006593f
C55 B.n27 VSUBS 0.006593f
C56 B.n28 VSUBS 0.006593f
C57 B.n29 VSUBS 0.006593f
C58 B.n30 VSUBS 0.006593f
C59 B.n31 VSUBS 0.006593f
C60 B.n32 VSUBS 0.006593f
C61 B.n33 VSUBS 0.006593f
C62 B.n34 VSUBS 0.006593f
C63 B.n35 VSUBS 0.006593f
C64 B.n36 VSUBS 0.006593f
C65 B.n37 VSUBS 0.006593f
C66 B.t11 VSUBS 0.305816f
C67 B.t10 VSUBS 0.320417f
C68 B.t9 VSUBS 0.645107f
C69 B.n38 VSUBS 0.420184f
C70 B.n39 VSUBS 0.290644f
C71 B.n40 VSUBS 0.015275f
C72 B.n41 VSUBS 0.006593f
C73 B.n42 VSUBS 0.006593f
C74 B.n43 VSUBS 0.006593f
C75 B.n44 VSUBS 0.006593f
C76 B.n45 VSUBS 0.006593f
C77 B.t8 VSUBS 0.305819f
C78 B.t7 VSUBS 0.32042f
C79 B.t6 VSUBS 0.645107f
C80 B.n46 VSUBS 0.420181f
C81 B.n47 VSUBS 0.290641f
C82 B.n48 VSUBS 0.006593f
C83 B.n49 VSUBS 0.006593f
C84 B.n50 VSUBS 0.006593f
C85 B.n51 VSUBS 0.006593f
C86 B.n52 VSUBS 0.006593f
C87 B.n53 VSUBS 0.006593f
C88 B.n54 VSUBS 0.006593f
C89 B.n55 VSUBS 0.006593f
C90 B.n56 VSUBS 0.006593f
C91 B.n57 VSUBS 0.006593f
C92 B.n58 VSUBS 0.006593f
C93 B.n59 VSUBS 0.006593f
C94 B.n60 VSUBS 0.006593f
C95 B.n61 VSUBS 0.006593f
C96 B.n62 VSUBS 0.006593f
C97 B.n63 VSUBS 0.006593f
C98 B.n64 VSUBS 0.006593f
C99 B.n65 VSUBS 0.006593f
C100 B.n66 VSUBS 0.006593f
C101 B.n67 VSUBS 0.006593f
C102 B.n68 VSUBS 0.006593f
C103 B.n69 VSUBS 0.006593f
C104 B.n70 VSUBS 0.006593f
C105 B.n71 VSUBS 0.006593f
C106 B.n72 VSUBS 0.006593f
C107 B.n73 VSUBS 0.006593f
C108 B.n74 VSUBS 0.006593f
C109 B.n75 VSUBS 0.014721f
C110 B.n76 VSUBS 0.006593f
C111 B.n77 VSUBS 0.006593f
C112 B.n78 VSUBS 0.006593f
C113 B.n79 VSUBS 0.006593f
C114 B.n80 VSUBS 0.006593f
C115 B.n81 VSUBS 0.006593f
C116 B.n82 VSUBS 0.006593f
C117 B.n83 VSUBS 0.006593f
C118 B.n84 VSUBS 0.006593f
C119 B.n85 VSUBS 0.006593f
C120 B.n86 VSUBS 0.006593f
C121 B.n87 VSUBS 0.006593f
C122 B.n88 VSUBS 0.006593f
C123 B.n89 VSUBS 0.006593f
C124 B.n90 VSUBS 0.006593f
C125 B.n91 VSUBS 0.006593f
C126 B.n92 VSUBS 0.014721f
C127 B.n93 VSUBS 0.006593f
C128 B.n94 VSUBS 0.006593f
C129 B.n95 VSUBS 0.006593f
C130 B.n96 VSUBS 0.006593f
C131 B.n97 VSUBS 0.006593f
C132 B.n98 VSUBS 0.006593f
C133 B.n99 VSUBS 0.006593f
C134 B.n100 VSUBS 0.006593f
C135 B.n101 VSUBS 0.006593f
C136 B.n102 VSUBS 0.006593f
C137 B.n103 VSUBS 0.006593f
C138 B.n104 VSUBS 0.006593f
C139 B.n105 VSUBS 0.006593f
C140 B.n106 VSUBS 0.006593f
C141 B.n107 VSUBS 0.006593f
C142 B.n108 VSUBS 0.006593f
C143 B.n109 VSUBS 0.006593f
C144 B.n110 VSUBS 0.006593f
C145 B.n111 VSUBS 0.006593f
C146 B.n112 VSUBS 0.006593f
C147 B.n113 VSUBS 0.006593f
C148 B.n114 VSUBS 0.006593f
C149 B.n115 VSUBS 0.006593f
C150 B.n116 VSUBS 0.006593f
C151 B.n117 VSUBS 0.006593f
C152 B.n118 VSUBS 0.006593f
C153 B.n119 VSUBS 0.006593f
C154 B.t1 VSUBS 0.305819f
C155 B.t2 VSUBS 0.32042f
C156 B.t0 VSUBS 0.645107f
C157 B.n120 VSUBS 0.420181f
C158 B.n121 VSUBS 0.290641f
C159 B.n122 VSUBS 0.015275f
C160 B.n123 VSUBS 0.006593f
C161 B.n124 VSUBS 0.006593f
C162 B.n125 VSUBS 0.006593f
C163 B.n126 VSUBS 0.006593f
C164 B.n127 VSUBS 0.006593f
C165 B.t4 VSUBS 0.305816f
C166 B.t5 VSUBS 0.320417f
C167 B.t3 VSUBS 0.645107f
C168 B.n128 VSUBS 0.420184f
C169 B.n129 VSUBS 0.290644f
C170 B.n130 VSUBS 0.006593f
C171 B.n131 VSUBS 0.006593f
C172 B.n132 VSUBS 0.006593f
C173 B.n133 VSUBS 0.006593f
C174 B.n134 VSUBS 0.006593f
C175 B.n135 VSUBS 0.006593f
C176 B.n136 VSUBS 0.006593f
C177 B.n137 VSUBS 0.006593f
C178 B.n138 VSUBS 0.006593f
C179 B.n139 VSUBS 0.006593f
C180 B.n140 VSUBS 0.006593f
C181 B.n141 VSUBS 0.006593f
C182 B.n142 VSUBS 0.006593f
C183 B.n143 VSUBS 0.006593f
C184 B.n144 VSUBS 0.006593f
C185 B.n145 VSUBS 0.006593f
C186 B.n146 VSUBS 0.006593f
C187 B.n147 VSUBS 0.006593f
C188 B.n148 VSUBS 0.006593f
C189 B.n149 VSUBS 0.006593f
C190 B.n150 VSUBS 0.006593f
C191 B.n151 VSUBS 0.006593f
C192 B.n152 VSUBS 0.006593f
C193 B.n153 VSUBS 0.006593f
C194 B.n154 VSUBS 0.006593f
C195 B.n155 VSUBS 0.006593f
C196 B.n156 VSUBS 0.006593f
C197 B.n157 VSUBS 0.014721f
C198 B.n158 VSUBS 0.006593f
C199 B.n159 VSUBS 0.006593f
C200 B.n160 VSUBS 0.006593f
C201 B.n161 VSUBS 0.006593f
C202 B.n162 VSUBS 0.006593f
C203 B.n163 VSUBS 0.006593f
C204 B.n164 VSUBS 0.006593f
C205 B.n165 VSUBS 0.006593f
C206 B.n166 VSUBS 0.006593f
C207 B.n167 VSUBS 0.006593f
C208 B.n168 VSUBS 0.006593f
C209 B.n169 VSUBS 0.006593f
C210 B.n170 VSUBS 0.006593f
C211 B.n171 VSUBS 0.006593f
C212 B.n172 VSUBS 0.006593f
C213 B.n173 VSUBS 0.006593f
C214 B.n174 VSUBS 0.006593f
C215 B.n175 VSUBS 0.006593f
C216 B.n176 VSUBS 0.006593f
C217 B.n177 VSUBS 0.006593f
C218 B.n178 VSUBS 0.006593f
C219 B.n179 VSUBS 0.006593f
C220 B.n180 VSUBS 0.006593f
C221 B.n181 VSUBS 0.006593f
C222 B.n182 VSUBS 0.006593f
C223 B.n183 VSUBS 0.006593f
C224 B.n184 VSUBS 0.006593f
C225 B.n185 VSUBS 0.006593f
C226 B.n186 VSUBS 0.013977f
C227 B.n187 VSUBS 0.013977f
C228 B.n188 VSUBS 0.014721f
C229 B.n189 VSUBS 0.006593f
C230 B.n190 VSUBS 0.006593f
C231 B.n191 VSUBS 0.006593f
C232 B.n192 VSUBS 0.006593f
C233 B.n193 VSUBS 0.006593f
C234 B.n194 VSUBS 0.006593f
C235 B.n195 VSUBS 0.006593f
C236 B.n196 VSUBS 0.006593f
C237 B.n197 VSUBS 0.006593f
C238 B.n198 VSUBS 0.006593f
C239 B.n199 VSUBS 0.006593f
C240 B.n200 VSUBS 0.006593f
C241 B.n201 VSUBS 0.006593f
C242 B.n202 VSUBS 0.006593f
C243 B.n203 VSUBS 0.006593f
C244 B.n204 VSUBS 0.006593f
C245 B.n205 VSUBS 0.006593f
C246 B.n206 VSUBS 0.006593f
C247 B.n207 VSUBS 0.006593f
C248 B.n208 VSUBS 0.006593f
C249 B.n209 VSUBS 0.006593f
C250 B.n210 VSUBS 0.006593f
C251 B.n211 VSUBS 0.006593f
C252 B.n212 VSUBS 0.006593f
C253 B.n213 VSUBS 0.006593f
C254 B.n214 VSUBS 0.006593f
C255 B.n215 VSUBS 0.006593f
C256 B.n216 VSUBS 0.006593f
C257 B.n217 VSUBS 0.006593f
C258 B.n218 VSUBS 0.006593f
C259 B.n219 VSUBS 0.006593f
C260 B.n220 VSUBS 0.006593f
C261 B.n221 VSUBS 0.006593f
C262 B.n222 VSUBS 0.006593f
C263 B.n223 VSUBS 0.006593f
C264 B.n224 VSUBS 0.006593f
C265 B.n225 VSUBS 0.006593f
C266 B.n226 VSUBS 0.006593f
C267 B.n227 VSUBS 0.006593f
C268 B.n228 VSUBS 0.006593f
C269 B.n229 VSUBS 0.006593f
C270 B.n230 VSUBS 0.006593f
C271 B.n231 VSUBS 0.006593f
C272 B.n232 VSUBS 0.006593f
C273 B.n233 VSUBS 0.006593f
C274 B.n234 VSUBS 0.006593f
C275 B.n235 VSUBS 0.006593f
C276 B.n236 VSUBS 0.006593f
C277 B.n237 VSUBS 0.006593f
C278 B.n238 VSUBS 0.006593f
C279 B.n239 VSUBS 0.006593f
C280 B.n240 VSUBS 0.006593f
C281 B.n241 VSUBS 0.006593f
C282 B.n242 VSUBS 0.006593f
C283 B.n243 VSUBS 0.006593f
C284 B.n244 VSUBS 0.006593f
C285 B.n245 VSUBS 0.006593f
C286 B.n246 VSUBS 0.006593f
C287 B.n247 VSUBS 0.006593f
C288 B.n248 VSUBS 0.006593f
C289 B.n249 VSUBS 0.006593f
C290 B.n250 VSUBS 0.006593f
C291 B.n251 VSUBS 0.006593f
C292 B.n252 VSUBS 0.006593f
C293 B.n253 VSUBS 0.006593f
C294 B.n254 VSUBS 0.006593f
C295 B.n255 VSUBS 0.006593f
C296 B.n256 VSUBS 0.006593f
C297 B.n257 VSUBS 0.006593f
C298 B.n258 VSUBS 0.006593f
C299 B.n259 VSUBS 0.006593f
C300 B.n260 VSUBS 0.006593f
C301 B.n261 VSUBS 0.006593f
C302 B.n262 VSUBS 0.006593f
C303 B.n263 VSUBS 0.006593f
C304 B.n264 VSUBS 0.006593f
C305 B.n265 VSUBS 0.006593f
C306 B.n266 VSUBS 0.006593f
C307 B.n267 VSUBS 0.006593f
C308 B.n268 VSUBS 0.006593f
C309 B.n269 VSUBS 0.006593f
C310 B.n270 VSUBS 0.006593f
C311 B.n271 VSUBS 0.006011f
C312 B.n272 VSUBS 0.015275f
C313 B.n273 VSUBS 0.003878f
C314 B.n274 VSUBS 0.006593f
C315 B.n275 VSUBS 0.006593f
C316 B.n276 VSUBS 0.006593f
C317 B.n277 VSUBS 0.006593f
C318 B.n278 VSUBS 0.006593f
C319 B.n279 VSUBS 0.006593f
C320 B.n280 VSUBS 0.006593f
C321 B.n281 VSUBS 0.006593f
C322 B.n282 VSUBS 0.006593f
C323 B.n283 VSUBS 0.006593f
C324 B.n284 VSUBS 0.006593f
C325 B.n285 VSUBS 0.006593f
C326 B.n286 VSUBS 0.003878f
C327 B.n287 VSUBS 0.006593f
C328 B.n288 VSUBS 0.006593f
C329 B.n289 VSUBS 0.006011f
C330 B.n290 VSUBS 0.006593f
C331 B.n291 VSUBS 0.006593f
C332 B.n292 VSUBS 0.006593f
C333 B.n293 VSUBS 0.006593f
C334 B.n294 VSUBS 0.006593f
C335 B.n295 VSUBS 0.006593f
C336 B.n296 VSUBS 0.006593f
C337 B.n297 VSUBS 0.006593f
C338 B.n298 VSUBS 0.006593f
C339 B.n299 VSUBS 0.006593f
C340 B.n300 VSUBS 0.006593f
C341 B.n301 VSUBS 0.006593f
C342 B.n302 VSUBS 0.006593f
C343 B.n303 VSUBS 0.006593f
C344 B.n304 VSUBS 0.006593f
C345 B.n305 VSUBS 0.006593f
C346 B.n306 VSUBS 0.006593f
C347 B.n307 VSUBS 0.006593f
C348 B.n308 VSUBS 0.006593f
C349 B.n309 VSUBS 0.006593f
C350 B.n310 VSUBS 0.006593f
C351 B.n311 VSUBS 0.006593f
C352 B.n312 VSUBS 0.006593f
C353 B.n313 VSUBS 0.006593f
C354 B.n314 VSUBS 0.006593f
C355 B.n315 VSUBS 0.006593f
C356 B.n316 VSUBS 0.006593f
C357 B.n317 VSUBS 0.006593f
C358 B.n318 VSUBS 0.006593f
C359 B.n319 VSUBS 0.006593f
C360 B.n320 VSUBS 0.006593f
C361 B.n321 VSUBS 0.006593f
C362 B.n322 VSUBS 0.006593f
C363 B.n323 VSUBS 0.006593f
C364 B.n324 VSUBS 0.006593f
C365 B.n325 VSUBS 0.006593f
C366 B.n326 VSUBS 0.006593f
C367 B.n327 VSUBS 0.006593f
C368 B.n328 VSUBS 0.006593f
C369 B.n329 VSUBS 0.006593f
C370 B.n330 VSUBS 0.006593f
C371 B.n331 VSUBS 0.006593f
C372 B.n332 VSUBS 0.006593f
C373 B.n333 VSUBS 0.006593f
C374 B.n334 VSUBS 0.006593f
C375 B.n335 VSUBS 0.006593f
C376 B.n336 VSUBS 0.006593f
C377 B.n337 VSUBS 0.006593f
C378 B.n338 VSUBS 0.006593f
C379 B.n339 VSUBS 0.006593f
C380 B.n340 VSUBS 0.006593f
C381 B.n341 VSUBS 0.006593f
C382 B.n342 VSUBS 0.006593f
C383 B.n343 VSUBS 0.006593f
C384 B.n344 VSUBS 0.006593f
C385 B.n345 VSUBS 0.006593f
C386 B.n346 VSUBS 0.006593f
C387 B.n347 VSUBS 0.006593f
C388 B.n348 VSUBS 0.006593f
C389 B.n349 VSUBS 0.006593f
C390 B.n350 VSUBS 0.006593f
C391 B.n351 VSUBS 0.006593f
C392 B.n352 VSUBS 0.006593f
C393 B.n353 VSUBS 0.006593f
C394 B.n354 VSUBS 0.006593f
C395 B.n355 VSUBS 0.006593f
C396 B.n356 VSUBS 0.006593f
C397 B.n357 VSUBS 0.006593f
C398 B.n358 VSUBS 0.006593f
C399 B.n359 VSUBS 0.006593f
C400 B.n360 VSUBS 0.006593f
C401 B.n361 VSUBS 0.006593f
C402 B.n362 VSUBS 0.006593f
C403 B.n363 VSUBS 0.006593f
C404 B.n364 VSUBS 0.006593f
C405 B.n365 VSUBS 0.006593f
C406 B.n366 VSUBS 0.006593f
C407 B.n367 VSUBS 0.006593f
C408 B.n368 VSUBS 0.006593f
C409 B.n369 VSUBS 0.006593f
C410 B.n370 VSUBS 0.006593f
C411 B.n371 VSUBS 0.014721f
C412 B.n372 VSUBS 0.013977f
C413 B.n373 VSUBS 0.013977f
C414 B.n374 VSUBS 0.006593f
C415 B.n375 VSUBS 0.006593f
C416 B.n376 VSUBS 0.006593f
C417 B.n377 VSUBS 0.006593f
C418 B.n378 VSUBS 0.006593f
C419 B.n379 VSUBS 0.006593f
C420 B.n380 VSUBS 0.006593f
C421 B.n381 VSUBS 0.006593f
C422 B.n382 VSUBS 0.006593f
C423 B.n383 VSUBS 0.006593f
C424 B.n384 VSUBS 0.006593f
C425 B.n385 VSUBS 0.006593f
C426 B.n386 VSUBS 0.006593f
C427 B.n387 VSUBS 0.006593f
C428 B.n388 VSUBS 0.006593f
C429 B.n389 VSUBS 0.006593f
C430 B.n390 VSUBS 0.006593f
C431 B.n391 VSUBS 0.006593f
C432 B.n392 VSUBS 0.006593f
C433 B.n393 VSUBS 0.006593f
C434 B.n394 VSUBS 0.006593f
C435 B.n395 VSUBS 0.006593f
C436 B.n396 VSUBS 0.006593f
C437 B.n397 VSUBS 0.006593f
C438 B.n398 VSUBS 0.006593f
C439 B.n399 VSUBS 0.006593f
C440 B.n400 VSUBS 0.006593f
C441 B.n401 VSUBS 0.006593f
C442 B.n402 VSUBS 0.006593f
C443 B.n403 VSUBS 0.006593f
C444 B.n404 VSUBS 0.006593f
C445 B.n405 VSUBS 0.006593f
C446 B.n406 VSUBS 0.006593f
C447 B.n407 VSUBS 0.006593f
C448 B.n408 VSUBS 0.006593f
C449 B.n409 VSUBS 0.006593f
C450 B.n410 VSUBS 0.006593f
C451 B.n411 VSUBS 0.006593f
C452 B.n412 VSUBS 0.006593f
C453 B.n413 VSUBS 0.006593f
C454 B.n414 VSUBS 0.006593f
C455 B.n415 VSUBS 0.006593f
C456 B.n416 VSUBS 0.006593f
C457 B.n417 VSUBS 0.006593f
C458 B.n418 VSUBS 0.006593f
C459 B.n419 VSUBS 0.006593f
C460 B.n420 VSUBS 0.013977f
C461 B.n421 VSUBS 0.014848f
C462 B.n422 VSUBS 0.013849f
C463 B.n423 VSUBS 0.006593f
C464 B.n424 VSUBS 0.006593f
C465 B.n425 VSUBS 0.006593f
C466 B.n426 VSUBS 0.006593f
C467 B.n427 VSUBS 0.006593f
C468 B.n428 VSUBS 0.006593f
C469 B.n429 VSUBS 0.006593f
C470 B.n430 VSUBS 0.006593f
C471 B.n431 VSUBS 0.006593f
C472 B.n432 VSUBS 0.006593f
C473 B.n433 VSUBS 0.006593f
C474 B.n434 VSUBS 0.006593f
C475 B.n435 VSUBS 0.006593f
C476 B.n436 VSUBS 0.006593f
C477 B.n437 VSUBS 0.006593f
C478 B.n438 VSUBS 0.006593f
C479 B.n439 VSUBS 0.006593f
C480 B.n440 VSUBS 0.006593f
C481 B.n441 VSUBS 0.006593f
C482 B.n442 VSUBS 0.006593f
C483 B.n443 VSUBS 0.006593f
C484 B.n444 VSUBS 0.006593f
C485 B.n445 VSUBS 0.006593f
C486 B.n446 VSUBS 0.006593f
C487 B.n447 VSUBS 0.006593f
C488 B.n448 VSUBS 0.006593f
C489 B.n449 VSUBS 0.006593f
C490 B.n450 VSUBS 0.006593f
C491 B.n451 VSUBS 0.006593f
C492 B.n452 VSUBS 0.006593f
C493 B.n453 VSUBS 0.006593f
C494 B.n454 VSUBS 0.006593f
C495 B.n455 VSUBS 0.006593f
C496 B.n456 VSUBS 0.006593f
C497 B.n457 VSUBS 0.006593f
C498 B.n458 VSUBS 0.006593f
C499 B.n459 VSUBS 0.006593f
C500 B.n460 VSUBS 0.006593f
C501 B.n461 VSUBS 0.006593f
C502 B.n462 VSUBS 0.006593f
C503 B.n463 VSUBS 0.006593f
C504 B.n464 VSUBS 0.006593f
C505 B.n465 VSUBS 0.006593f
C506 B.n466 VSUBS 0.006593f
C507 B.n467 VSUBS 0.006593f
C508 B.n468 VSUBS 0.006593f
C509 B.n469 VSUBS 0.006593f
C510 B.n470 VSUBS 0.006593f
C511 B.n471 VSUBS 0.006593f
C512 B.n472 VSUBS 0.006593f
C513 B.n473 VSUBS 0.006593f
C514 B.n474 VSUBS 0.006593f
C515 B.n475 VSUBS 0.006593f
C516 B.n476 VSUBS 0.006593f
C517 B.n477 VSUBS 0.006593f
C518 B.n478 VSUBS 0.006593f
C519 B.n479 VSUBS 0.006593f
C520 B.n480 VSUBS 0.006593f
C521 B.n481 VSUBS 0.006593f
C522 B.n482 VSUBS 0.006593f
C523 B.n483 VSUBS 0.006593f
C524 B.n484 VSUBS 0.006593f
C525 B.n485 VSUBS 0.006593f
C526 B.n486 VSUBS 0.006593f
C527 B.n487 VSUBS 0.006593f
C528 B.n488 VSUBS 0.006593f
C529 B.n489 VSUBS 0.006593f
C530 B.n490 VSUBS 0.006593f
C531 B.n491 VSUBS 0.006593f
C532 B.n492 VSUBS 0.006593f
C533 B.n493 VSUBS 0.006593f
C534 B.n494 VSUBS 0.006593f
C535 B.n495 VSUBS 0.006593f
C536 B.n496 VSUBS 0.006593f
C537 B.n497 VSUBS 0.006593f
C538 B.n498 VSUBS 0.006593f
C539 B.n499 VSUBS 0.006593f
C540 B.n500 VSUBS 0.006593f
C541 B.n501 VSUBS 0.006593f
C542 B.n502 VSUBS 0.006593f
C543 B.n503 VSUBS 0.006593f
C544 B.n504 VSUBS 0.006593f
C545 B.n505 VSUBS 0.006011f
C546 B.n506 VSUBS 0.015275f
C547 B.n507 VSUBS 0.003878f
C548 B.n508 VSUBS 0.006593f
C549 B.n509 VSUBS 0.006593f
C550 B.n510 VSUBS 0.006593f
C551 B.n511 VSUBS 0.006593f
C552 B.n512 VSUBS 0.006593f
C553 B.n513 VSUBS 0.006593f
C554 B.n514 VSUBS 0.006593f
C555 B.n515 VSUBS 0.006593f
C556 B.n516 VSUBS 0.006593f
C557 B.n517 VSUBS 0.006593f
C558 B.n518 VSUBS 0.006593f
C559 B.n519 VSUBS 0.006593f
C560 B.n520 VSUBS 0.003878f
C561 B.n521 VSUBS 0.006593f
C562 B.n522 VSUBS 0.006593f
C563 B.n523 VSUBS 0.006011f
C564 B.n524 VSUBS 0.006593f
C565 B.n525 VSUBS 0.006593f
C566 B.n526 VSUBS 0.006593f
C567 B.n527 VSUBS 0.006593f
C568 B.n528 VSUBS 0.006593f
C569 B.n529 VSUBS 0.006593f
C570 B.n530 VSUBS 0.006593f
C571 B.n531 VSUBS 0.006593f
C572 B.n532 VSUBS 0.006593f
C573 B.n533 VSUBS 0.006593f
C574 B.n534 VSUBS 0.006593f
C575 B.n535 VSUBS 0.006593f
C576 B.n536 VSUBS 0.006593f
C577 B.n537 VSUBS 0.006593f
C578 B.n538 VSUBS 0.006593f
C579 B.n539 VSUBS 0.006593f
C580 B.n540 VSUBS 0.006593f
C581 B.n541 VSUBS 0.006593f
C582 B.n542 VSUBS 0.006593f
C583 B.n543 VSUBS 0.006593f
C584 B.n544 VSUBS 0.006593f
C585 B.n545 VSUBS 0.006593f
C586 B.n546 VSUBS 0.006593f
C587 B.n547 VSUBS 0.006593f
C588 B.n548 VSUBS 0.006593f
C589 B.n549 VSUBS 0.006593f
C590 B.n550 VSUBS 0.006593f
C591 B.n551 VSUBS 0.006593f
C592 B.n552 VSUBS 0.006593f
C593 B.n553 VSUBS 0.006593f
C594 B.n554 VSUBS 0.006593f
C595 B.n555 VSUBS 0.006593f
C596 B.n556 VSUBS 0.006593f
C597 B.n557 VSUBS 0.006593f
C598 B.n558 VSUBS 0.006593f
C599 B.n559 VSUBS 0.006593f
C600 B.n560 VSUBS 0.006593f
C601 B.n561 VSUBS 0.006593f
C602 B.n562 VSUBS 0.006593f
C603 B.n563 VSUBS 0.006593f
C604 B.n564 VSUBS 0.006593f
C605 B.n565 VSUBS 0.006593f
C606 B.n566 VSUBS 0.006593f
C607 B.n567 VSUBS 0.006593f
C608 B.n568 VSUBS 0.006593f
C609 B.n569 VSUBS 0.006593f
C610 B.n570 VSUBS 0.006593f
C611 B.n571 VSUBS 0.006593f
C612 B.n572 VSUBS 0.006593f
C613 B.n573 VSUBS 0.006593f
C614 B.n574 VSUBS 0.006593f
C615 B.n575 VSUBS 0.006593f
C616 B.n576 VSUBS 0.006593f
C617 B.n577 VSUBS 0.006593f
C618 B.n578 VSUBS 0.006593f
C619 B.n579 VSUBS 0.006593f
C620 B.n580 VSUBS 0.006593f
C621 B.n581 VSUBS 0.006593f
C622 B.n582 VSUBS 0.006593f
C623 B.n583 VSUBS 0.006593f
C624 B.n584 VSUBS 0.006593f
C625 B.n585 VSUBS 0.006593f
C626 B.n586 VSUBS 0.006593f
C627 B.n587 VSUBS 0.006593f
C628 B.n588 VSUBS 0.006593f
C629 B.n589 VSUBS 0.006593f
C630 B.n590 VSUBS 0.006593f
C631 B.n591 VSUBS 0.006593f
C632 B.n592 VSUBS 0.006593f
C633 B.n593 VSUBS 0.006593f
C634 B.n594 VSUBS 0.006593f
C635 B.n595 VSUBS 0.006593f
C636 B.n596 VSUBS 0.006593f
C637 B.n597 VSUBS 0.006593f
C638 B.n598 VSUBS 0.006593f
C639 B.n599 VSUBS 0.006593f
C640 B.n600 VSUBS 0.006593f
C641 B.n601 VSUBS 0.006593f
C642 B.n602 VSUBS 0.006593f
C643 B.n603 VSUBS 0.006593f
C644 B.n604 VSUBS 0.006593f
C645 B.n605 VSUBS 0.014721f
C646 B.n606 VSUBS 0.013977f
C647 B.n607 VSUBS 0.013977f
C648 B.n608 VSUBS 0.006593f
C649 B.n609 VSUBS 0.006593f
C650 B.n610 VSUBS 0.006593f
C651 B.n611 VSUBS 0.006593f
C652 B.n612 VSUBS 0.006593f
C653 B.n613 VSUBS 0.006593f
C654 B.n614 VSUBS 0.006593f
C655 B.n615 VSUBS 0.006593f
C656 B.n616 VSUBS 0.006593f
C657 B.n617 VSUBS 0.006593f
C658 B.n618 VSUBS 0.006593f
C659 B.n619 VSUBS 0.006593f
C660 B.n620 VSUBS 0.006593f
C661 B.n621 VSUBS 0.006593f
C662 B.n622 VSUBS 0.006593f
C663 B.n623 VSUBS 0.006593f
C664 B.n624 VSUBS 0.006593f
C665 B.n625 VSUBS 0.006593f
C666 B.n626 VSUBS 0.006593f
C667 B.n627 VSUBS 0.006593f
C668 B.n628 VSUBS 0.006593f
C669 B.n629 VSUBS 0.006593f
C670 B.n630 VSUBS 0.006593f
C671 B.n631 VSUBS 0.014928f
C672 VDD2.n0 VSUBS 0.022433f
C673 VDD2.n1 VSUBS 0.020337f
C674 VDD2.n2 VSUBS 0.010928f
C675 VDD2.n3 VSUBS 0.02583f
C676 VDD2.n4 VSUBS 0.011571f
C677 VDD2.n5 VSUBS 0.020337f
C678 VDD2.n6 VSUBS 0.010928f
C679 VDD2.n7 VSUBS 0.02583f
C680 VDD2.n8 VSUBS 0.011571f
C681 VDD2.n9 VSUBS 0.020337f
C682 VDD2.n10 VSUBS 0.010928f
C683 VDD2.n11 VSUBS 0.02583f
C684 VDD2.n12 VSUBS 0.011571f
C685 VDD2.n13 VSUBS 0.020337f
C686 VDD2.n14 VSUBS 0.010928f
C687 VDD2.n15 VSUBS 0.02583f
C688 VDD2.n16 VSUBS 0.011571f
C689 VDD2.n17 VSUBS 0.020337f
C690 VDD2.n18 VSUBS 0.010928f
C691 VDD2.n19 VSUBS 0.02583f
C692 VDD2.n20 VSUBS 0.011571f
C693 VDD2.n21 VSUBS 0.020337f
C694 VDD2.n22 VSUBS 0.010928f
C695 VDD2.n23 VSUBS 0.02583f
C696 VDD2.n24 VSUBS 0.011571f
C697 VDD2.n25 VSUBS 0.020337f
C698 VDD2.n26 VSUBS 0.010928f
C699 VDD2.n27 VSUBS 0.02583f
C700 VDD2.n28 VSUBS 0.011571f
C701 VDD2.n29 VSUBS 0.154752f
C702 VDD2.t1 VSUBS 0.055393f
C703 VDD2.n30 VSUBS 0.019372f
C704 VDD2.n31 VSUBS 0.016432f
C705 VDD2.n32 VSUBS 0.010928f
C706 VDD2.n33 VSUBS 1.47394f
C707 VDD2.n34 VSUBS 0.020337f
C708 VDD2.n35 VSUBS 0.010928f
C709 VDD2.n36 VSUBS 0.011571f
C710 VDD2.n37 VSUBS 0.02583f
C711 VDD2.n38 VSUBS 0.02583f
C712 VDD2.n39 VSUBS 0.011571f
C713 VDD2.n40 VSUBS 0.010928f
C714 VDD2.n41 VSUBS 0.020337f
C715 VDD2.n42 VSUBS 0.020337f
C716 VDD2.n43 VSUBS 0.010928f
C717 VDD2.n44 VSUBS 0.011571f
C718 VDD2.n45 VSUBS 0.02583f
C719 VDD2.n46 VSUBS 0.02583f
C720 VDD2.n47 VSUBS 0.011571f
C721 VDD2.n48 VSUBS 0.010928f
C722 VDD2.n49 VSUBS 0.020337f
C723 VDD2.n50 VSUBS 0.020337f
C724 VDD2.n51 VSUBS 0.010928f
C725 VDD2.n52 VSUBS 0.011571f
C726 VDD2.n53 VSUBS 0.02583f
C727 VDD2.n54 VSUBS 0.02583f
C728 VDD2.n55 VSUBS 0.011571f
C729 VDD2.n56 VSUBS 0.010928f
C730 VDD2.n57 VSUBS 0.020337f
C731 VDD2.n58 VSUBS 0.020337f
C732 VDD2.n59 VSUBS 0.010928f
C733 VDD2.n60 VSUBS 0.011571f
C734 VDD2.n61 VSUBS 0.02583f
C735 VDD2.n62 VSUBS 0.02583f
C736 VDD2.n63 VSUBS 0.011571f
C737 VDD2.n64 VSUBS 0.010928f
C738 VDD2.n65 VSUBS 0.020337f
C739 VDD2.n66 VSUBS 0.020337f
C740 VDD2.n67 VSUBS 0.010928f
C741 VDD2.n68 VSUBS 0.011571f
C742 VDD2.n69 VSUBS 0.02583f
C743 VDD2.n70 VSUBS 0.02583f
C744 VDD2.n71 VSUBS 0.02583f
C745 VDD2.n72 VSUBS 0.011571f
C746 VDD2.n73 VSUBS 0.010928f
C747 VDD2.n74 VSUBS 0.020337f
C748 VDD2.n75 VSUBS 0.020337f
C749 VDD2.n76 VSUBS 0.010928f
C750 VDD2.n77 VSUBS 0.011249f
C751 VDD2.n78 VSUBS 0.011249f
C752 VDD2.n79 VSUBS 0.02583f
C753 VDD2.n80 VSUBS 0.02583f
C754 VDD2.n81 VSUBS 0.011571f
C755 VDD2.n82 VSUBS 0.010928f
C756 VDD2.n83 VSUBS 0.020337f
C757 VDD2.n84 VSUBS 0.020337f
C758 VDD2.n85 VSUBS 0.010928f
C759 VDD2.n86 VSUBS 0.011571f
C760 VDD2.n87 VSUBS 0.02583f
C761 VDD2.n88 VSUBS 0.062829f
C762 VDD2.n89 VSUBS 0.011571f
C763 VDD2.n90 VSUBS 0.010928f
C764 VDD2.n91 VSUBS 0.049785f
C765 VDD2.n92 VSUBS 0.64314f
C766 VDD2.n93 VSUBS 0.022433f
C767 VDD2.n94 VSUBS 0.020337f
C768 VDD2.n95 VSUBS 0.010928f
C769 VDD2.n96 VSUBS 0.02583f
C770 VDD2.n97 VSUBS 0.011571f
C771 VDD2.n98 VSUBS 0.020337f
C772 VDD2.n99 VSUBS 0.010928f
C773 VDD2.n100 VSUBS 0.02583f
C774 VDD2.n101 VSUBS 0.011571f
C775 VDD2.n102 VSUBS 0.020337f
C776 VDD2.n103 VSUBS 0.010928f
C777 VDD2.n104 VSUBS 0.02583f
C778 VDD2.n105 VSUBS 0.02583f
C779 VDD2.n106 VSUBS 0.011571f
C780 VDD2.n107 VSUBS 0.020337f
C781 VDD2.n108 VSUBS 0.010928f
C782 VDD2.n109 VSUBS 0.02583f
C783 VDD2.n110 VSUBS 0.011571f
C784 VDD2.n111 VSUBS 0.020337f
C785 VDD2.n112 VSUBS 0.010928f
C786 VDD2.n113 VSUBS 0.02583f
C787 VDD2.n114 VSUBS 0.011571f
C788 VDD2.n115 VSUBS 0.020337f
C789 VDD2.n116 VSUBS 0.010928f
C790 VDD2.n117 VSUBS 0.02583f
C791 VDD2.n118 VSUBS 0.011571f
C792 VDD2.n119 VSUBS 0.020337f
C793 VDD2.n120 VSUBS 0.010928f
C794 VDD2.n121 VSUBS 0.02583f
C795 VDD2.n122 VSUBS 0.011571f
C796 VDD2.n123 VSUBS 0.154752f
C797 VDD2.t0 VSUBS 0.055393f
C798 VDD2.n124 VSUBS 0.019372f
C799 VDD2.n125 VSUBS 0.016432f
C800 VDD2.n126 VSUBS 0.010928f
C801 VDD2.n127 VSUBS 1.47394f
C802 VDD2.n128 VSUBS 0.020337f
C803 VDD2.n129 VSUBS 0.010928f
C804 VDD2.n130 VSUBS 0.011571f
C805 VDD2.n131 VSUBS 0.02583f
C806 VDD2.n132 VSUBS 0.02583f
C807 VDD2.n133 VSUBS 0.011571f
C808 VDD2.n134 VSUBS 0.010928f
C809 VDD2.n135 VSUBS 0.020337f
C810 VDD2.n136 VSUBS 0.020337f
C811 VDD2.n137 VSUBS 0.010928f
C812 VDD2.n138 VSUBS 0.011571f
C813 VDD2.n139 VSUBS 0.02583f
C814 VDD2.n140 VSUBS 0.02583f
C815 VDD2.n141 VSUBS 0.011571f
C816 VDD2.n142 VSUBS 0.010928f
C817 VDD2.n143 VSUBS 0.020337f
C818 VDD2.n144 VSUBS 0.020337f
C819 VDD2.n145 VSUBS 0.010928f
C820 VDD2.n146 VSUBS 0.011571f
C821 VDD2.n147 VSUBS 0.02583f
C822 VDD2.n148 VSUBS 0.02583f
C823 VDD2.n149 VSUBS 0.011571f
C824 VDD2.n150 VSUBS 0.010928f
C825 VDD2.n151 VSUBS 0.020337f
C826 VDD2.n152 VSUBS 0.020337f
C827 VDD2.n153 VSUBS 0.010928f
C828 VDD2.n154 VSUBS 0.011571f
C829 VDD2.n155 VSUBS 0.02583f
C830 VDD2.n156 VSUBS 0.02583f
C831 VDD2.n157 VSUBS 0.011571f
C832 VDD2.n158 VSUBS 0.010928f
C833 VDD2.n159 VSUBS 0.020337f
C834 VDD2.n160 VSUBS 0.020337f
C835 VDD2.n161 VSUBS 0.010928f
C836 VDD2.n162 VSUBS 0.011571f
C837 VDD2.n163 VSUBS 0.02583f
C838 VDD2.n164 VSUBS 0.02583f
C839 VDD2.n165 VSUBS 0.011571f
C840 VDD2.n166 VSUBS 0.010928f
C841 VDD2.n167 VSUBS 0.020337f
C842 VDD2.n168 VSUBS 0.020337f
C843 VDD2.n169 VSUBS 0.010928f
C844 VDD2.n170 VSUBS 0.011249f
C845 VDD2.n171 VSUBS 0.011249f
C846 VDD2.n172 VSUBS 0.02583f
C847 VDD2.n173 VSUBS 0.02583f
C848 VDD2.n174 VSUBS 0.011571f
C849 VDD2.n175 VSUBS 0.010928f
C850 VDD2.n176 VSUBS 0.020337f
C851 VDD2.n177 VSUBS 0.020337f
C852 VDD2.n178 VSUBS 0.010928f
C853 VDD2.n179 VSUBS 0.011571f
C854 VDD2.n180 VSUBS 0.02583f
C855 VDD2.n181 VSUBS 0.062829f
C856 VDD2.n182 VSUBS 0.011571f
C857 VDD2.n183 VSUBS 0.010928f
C858 VDD2.n184 VSUBS 0.049785f
C859 VDD2.n185 VSUBS 0.045714f
C860 VDD2.n186 VSUBS 2.65441f
C861 VN.t0 VSUBS 3.02973f
C862 VN.t1 VSUBS 3.26114f
C863 VDD1.n0 VSUBS 0.022266f
C864 VDD1.n1 VSUBS 0.020185f
C865 VDD1.n2 VSUBS 0.010847f
C866 VDD1.n3 VSUBS 0.025637f
C867 VDD1.n4 VSUBS 0.011485f
C868 VDD1.n5 VSUBS 0.020185f
C869 VDD1.n6 VSUBS 0.010847f
C870 VDD1.n7 VSUBS 0.025637f
C871 VDD1.n8 VSUBS 0.011485f
C872 VDD1.n9 VSUBS 0.020185f
C873 VDD1.n10 VSUBS 0.010847f
C874 VDD1.n11 VSUBS 0.025637f
C875 VDD1.n12 VSUBS 0.025637f
C876 VDD1.n13 VSUBS 0.011485f
C877 VDD1.n14 VSUBS 0.020185f
C878 VDD1.n15 VSUBS 0.010847f
C879 VDD1.n16 VSUBS 0.025637f
C880 VDD1.n17 VSUBS 0.011485f
C881 VDD1.n18 VSUBS 0.020185f
C882 VDD1.n19 VSUBS 0.010847f
C883 VDD1.n20 VSUBS 0.025637f
C884 VDD1.n21 VSUBS 0.011485f
C885 VDD1.n22 VSUBS 0.020185f
C886 VDD1.n23 VSUBS 0.010847f
C887 VDD1.n24 VSUBS 0.025637f
C888 VDD1.n25 VSUBS 0.011485f
C889 VDD1.n26 VSUBS 0.020185f
C890 VDD1.n27 VSUBS 0.010847f
C891 VDD1.n28 VSUBS 0.025637f
C892 VDD1.n29 VSUBS 0.011485f
C893 VDD1.n30 VSUBS 0.153598f
C894 VDD1.t1 VSUBS 0.054979f
C895 VDD1.n31 VSUBS 0.019228f
C896 VDD1.n32 VSUBS 0.016309f
C897 VDD1.n33 VSUBS 0.010847f
C898 VDD1.n34 VSUBS 1.46296f
C899 VDD1.n35 VSUBS 0.020185f
C900 VDD1.n36 VSUBS 0.010847f
C901 VDD1.n37 VSUBS 0.011485f
C902 VDD1.n38 VSUBS 0.025637f
C903 VDD1.n39 VSUBS 0.025637f
C904 VDD1.n40 VSUBS 0.011485f
C905 VDD1.n41 VSUBS 0.010847f
C906 VDD1.n42 VSUBS 0.020185f
C907 VDD1.n43 VSUBS 0.020185f
C908 VDD1.n44 VSUBS 0.010847f
C909 VDD1.n45 VSUBS 0.011485f
C910 VDD1.n46 VSUBS 0.025637f
C911 VDD1.n47 VSUBS 0.025637f
C912 VDD1.n48 VSUBS 0.011485f
C913 VDD1.n49 VSUBS 0.010847f
C914 VDD1.n50 VSUBS 0.020185f
C915 VDD1.n51 VSUBS 0.020185f
C916 VDD1.n52 VSUBS 0.010847f
C917 VDD1.n53 VSUBS 0.011485f
C918 VDD1.n54 VSUBS 0.025637f
C919 VDD1.n55 VSUBS 0.025637f
C920 VDD1.n56 VSUBS 0.011485f
C921 VDD1.n57 VSUBS 0.010847f
C922 VDD1.n58 VSUBS 0.020185f
C923 VDD1.n59 VSUBS 0.020185f
C924 VDD1.n60 VSUBS 0.010847f
C925 VDD1.n61 VSUBS 0.011485f
C926 VDD1.n62 VSUBS 0.025637f
C927 VDD1.n63 VSUBS 0.025637f
C928 VDD1.n64 VSUBS 0.011485f
C929 VDD1.n65 VSUBS 0.010847f
C930 VDD1.n66 VSUBS 0.020185f
C931 VDD1.n67 VSUBS 0.020185f
C932 VDD1.n68 VSUBS 0.010847f
C933 VDD1.n69 VSUBS 0.011485f
C934 VDD1.n70 VSUBS 0.025637f
C935 VDD1.n71 VSUBS 0.025637f
C936 VDD1.n72 VSUBS 0.011485f
C937 VDD1.n73 VSUBS 0.010847f
C938 VDD1.n74 VSUBS 0.020185f
C939 VDD1.n75 VSUBS 0.020185f
C940 VDD1.n76 VSUBS 0.010847f
C941 VDD1.n77 VSUBS 0.011165f
C942 VDD1.n78 VSUBS 0.011165f
C943 VDD1.n79 VSUBS 0.025637f
C944 VDD1.n80 VSUBS 0.025637f
C945 VDD1.n81 VSUBS 0.011485f
C946 VDD1.n82 VSUBS 0.010847f
C947 VDD1.n83 VSUBS 0.020185f
C948 VDD1.n84 VSUBS 0.020185f
C949 VDD1.n85 VSUBS 0.010847f
C950 VDD1.n86 VSUBS 0.011485f
C951 VDD1.n87 VSUBS 0.025637f
C952 VDD1.n88 VSUBS 0.06236f
C953 VDD1.n89 VSUBS 0.011485f
C954 VDD1.n90 VSUBS 0.010847f
C955 VDD1.n91 VSUBS 0.049414f
C956 VDD1.n92 VSUBS 0.04579f
C957 VDD1.n93 VSUBS 0.022266f
C958 VDD1.n94 VSUBS 0.020185f
C959 VDD1.n95 VSUBS 0.010847f
C960 VDD1.n96 VSUBS 0.025637f
C961 VDD1.n97 VSUBS 0.011485f
C962 VDD1.n98 VSUBS 0.020185f
C963 VDD1.n99 VSUBS 0.010847f
C964 VDD1.n100 VSUBS 0.025637f
C965 VDD1.n101 VSUBS 0.011485f
C966 VDD1.n102 VSUBS 0.020185f
C967 VDD1.n103 VSUBS 0.010847f
C968 VDD1.n104 VSUBS 0.025637f
C969 VDD1.n105 VSUBS 0.011485f
C970 VDD1.n106 VSUBS 0.020185f
C971 VDD1.n107 VSUBS 0.010847f
C972 VDD1.n108 VSUBS 0.025637f
C973 VDD1.n109 VSUBS 0.011485f
C974 VDD1.n110 VSUBS 0.020185f
C975 VDD1.n111 VSUBS 0.010847f
C976 VDD1.n112 VSUBS 0.025637f
C977 VDD1.n113 VSUBS 0.011485f
C978 VDD1.n114 VSUBS 0.020185f
C979 VDD1.n115 VSUBS 0.010847f
C980 VDD1.n116 VSUBS 0.025637f
C981 VDD1.n117 VSUBS 0.011485f
C982 VDD1.n118 VSUBS 0.020185f
C983 VDD1.n119 VSUBS 0.010847f
C984 VDD1.n120 VSUBS 0.025637f
C985 VDD1.n121 VSUBS 0.011485f
C986 VDD1.n122 VSUBS 0.153598f
C987 VDD1.t0 VSUBS 0.054979f
C988 VDD1.n123 VSUBS 0.019228f
C989 VDD1.n124 VSUBS 0.016309f
C990 VDD1.n125 VSUBS 0.010847f
C991 VDD1.n126 VSUBS 1.46296f
C992 VDD1.n127 VSUBS 0.020185f
C993 VDD1.n128 VSUBS 0.010847f
C994 VDD1.n129 VSUBS 0.011485f
C995 VDD1.n130 VSUBS 0.025637f
C996 VDD1.n131 VSUBS 0.025637f
C997 VDD1.n132 VSUBS 0.011485f
C998 VDD1.n133 VSUBS 0.010847f
C999 VDD1.n134 VSUBS 0.020185f
C1000 VDD1.n135 VSUBS 0.020185f
C1001 VDD1.n136 VSUBS 0.010847f
C1002 VDD1.n137 VSUBS 0.011485f
C1003 VDD1.n138 VSUBS 0.025637f
C1004 VDD1.n139 VSUBS 0.025637f
C1005 VDD1.n140 VSUBS 0.011485f
C1006 VDD1.n141 VSUBS 0.010847f
C1007 VDD1.n142 VSUBS 0.020185f
C1008 VDD1.n143 VSUBS 0.020185f
C1009 VDD1.n144 VSUBS 0.010847f
C1010 VDD1.n145 VSUBS 0.011485f
C1011 VDD1.n146 VSUBS 0.025637f
C1012 VDD1.n147 VSUBS 0.025637f
C1013 VDD1.n148 VSUBS 0.011485f
C1014 VDD1.n149 VSUBS 0.010847f
C1015 VDD1.n150 VSUBS 0.020185f
C1016 VDD1.n151 VSUBS 0.020185f
C1017 VDD1.n152 VSUBS 0.010847f
C1018 VDD1.n153 VSUBS 0.011485f
C1019 VDD1.n154 VSUBS 0.025637f
C1020 VDD1.n155 VSUBS 0.025637f
C1021 VDD1.n156 VSUBS 0.011485f
C1022 VDD1.n157 VSUBS 0.010847f
C1023 VDD1.n158 VSUBS 0.020185f
C1024 VDD1.n159 VSUBS 0.020185f
C1025 VDD1.n160 VSUBS 0.010847f
C1026 VDD1.n161 VSUBS 0.011485f
C1027 VDD1.n162 VSUBS 0.025637f
C1028 VDD1.n163 VSUBS 0.025637f
C1029 VDD1.n164 VSUBS 0.025637f
C1030 VDD1.n165 VSUBS 0.011485f
C1031 VDD1.n166 VSUBS 0.010847f
C1032 VDD1.n167 VSUBS 0.020185f
C1033 VDD1.n168 VSUBS 0.020185f
C1034 VDD1.n169 VSUBS 0.010847f
C1035 VDD1.n170 VSUBS 0.011165f
C1036 VDD1.n171 VSUBS 0.011165f
C1037 VDD1.n172 VSUBS 0.025637f
C1038 VDD1.n173 VSUBS 0.025637f
C1039 VDD1.n174 VSUBS 0.011485f
C1040 VDD1.n175 VSUBS 0.010847f
C1041 VDD1.n176 VSUBS 0.020185f
C1042 VDD1.n177 VSUBS 0.020185f
C1043 VDD1.n178 VSUBS 0.010847f
C1044 VDD1.n179 VSUBS 0.011485f
C1045 VDD1.n180 VSUBS 0.025637f
C1046 VDD1.n181 VSUBS 0.06236f
C1047 VDD1.n182 VSUBS 0.011485f
C1048 VDD1.n183 VSUBS 0.010847f
C1049 VDD1.n184 VSUBS 0.049414f
C1050 VDD1.n185 VSUBS 0.668762f
C1051 VTAIL.n0 VSUBS 0.030869f
C1052 VTAIL.n1 VSUBS 0.027985f
C1053 VTAIL.n2 VSUBS 0.015038f
C1054 VTAIL.n3 VSUBS 0.035544f
C1055 VTAIL.n4 VSUBS 0.015922f
C1056 VTAIL.n5 VSUBS 0.027985f
C1057 VTAIL.n6 VSUBS 0.015038f
C1058 VTAIL.n7 VSUBS 0.035544f
C1059 VTAIL.n8 VSUBS 0.015922f
C1060 VTAIL.n9 VSUBS 0.027985f
C1061 VTAIL.n10 VSUBS 0.015038f
C1062 VTAIL.n11 VSUBS 0.035544f
C1063 VTAIL.n12 VSUBS 0.015922f
C1064 VTAIL.n13 VSUBS 0.027985f
C1065 VTAIL.n14 VSUBS 0.015038f
C1066 VTAIL.n15 VSUBS 0.035544f
C1067 VTAIL.n16 VSUBS 0.015922f
C1068 VTAIL.n17 VSUBS 0.027985f
C1069 VTAIL.n18 VSUBS 0.015038f
C1070 VTAIL.n19 VSUBS 0.035544f
C1071 VTAIL.n20 VSUBS 0.015922f
C1072 VTAIL.n21 VSUBS 0.027985f
C1073 VTAIL.n22 VSUBS 0.015038f
C1074 VTAIL.n23 VSUBS 0.035544f
C1075 VTAIL.n24 VSUBS 0.015922f
C1076 VTAIL.n25 VSUBS 0.027985f
C1077 VTAIL.n26 VSUBS 0.015038f
C1078 VTAIL.n27 VSUBS 0.035544f
C1079 VTAIL.n28 VSUBS 0.015922f
C1080 VTAIL.n29 VSUBS 0.21295f
C1081 VTAIL.t3 VSUBS 0.076224f
C1082 VTAIL.n30 VSUBS 0.026658f
C1083 VTAIL.n31 VSUBS 0.022611f
C1084 VTAIL.n32 VSUBS 0.015038f
C1085 VTAIL.n33 VSUBS 2.02826f
C1086 VTAIL.n34 VSUBS 0.027985f
C1087 VTAIL.n35 VSUBS 0.015038f
C1088 VTAIL.n36 VSUBS 0.015922f
C1089 VTAIL.n37 VSUBS 0.035544f
C1090 VTAIL.n38 VSUBS 0.035544f
C1091 VTAIL.n39 VSUBS 0.015922f
C1092 VTAIL.n40 VSUBS 0.015038f
C1093 VTAIL.n41 VSUBS 0.027985f
C1094 VTAIL.n42 VSUBS 0.027985f
C1095 VTAIL.n43 VSUBS 0.015038f
C1096 VTAIL.n44 VSUBS 0.015922f
C1097 VTAIL.n45 VSUBS 0.035544f
C1098 VTAIL.n46 VSUBS 0.035544f
C1099 VTAIL.n47 VSUBS 0.015922f
C1100 VTAIL.n48 VSUBS 0.015038f
C1101 VTAIL.n49 VSUBS 0.027985f
C1102 VTAIL.n50 VSUBS 0.027985f
C1103 VTAIL.n51 VSUBS 0.015038f
C1104 VTAIL.n52 VSUBS 0.015922f
C1105 VTAIL.n53 VSUBS 0.035544f
C1106 VTAIL.n54 VSUBS 0.035544f
C1107 VTAIL.n55 VSUBS 0.015922f
C1108 VTAIL.n56 VSUBS 0.015038f
C1109 VTAIL.n57 VSUBS 0.027985f
C1110 VTAIL.n58 VSUBS 0.027985f
C1111 VTAIL.n59 VSUBS 0.015038f
C1112 VTAIL.n60 VSUBS 0.015922f
C1113 VTAIL.n61 VSUBS 0.035544f
C1114 VTAIL.n62 VSUBS 0.035544f
C1115 VTAIL.n63 VSUBS 0.015922f
C1116 VTAIL.n64 VSUBS 0.015038f
C1117 VTAIL.n65 VSUBS 0.027985f
C1118 VTAIL.n66 VSUBS 0.027985f
C1119 VTAIL.n67 VSUBS 0.015038f
C1120 VTAIL.n68 VSUBS 0.015922f
C1121 VTAIL.n69 VSUBS 0.035544f
C1122 VTAIL.n70 VSUBS 0.035544f
C1123 VTAIL.n71 VSUBS 0.035544f
C1124 VTAIL.n72 VSUBS 0.015922f
C1125 VTAIL.n73 VSUBS 0.015038f
C1126 VTAIL.n74 VSUBS 0.027985f
C1127 VTAIL.n75 VSUBS 0.027985f
C1128 VTAIL.n76 VSUBS 0.015038f
C1129 VTAIL.n77 VSUBS 0.01548f
C1130 VTAIL.n78 VSUBS 0.01548f
C1131 VTAIL.n79 VSUBS 0.035544f
C1132 VTAIL.n80 VSUBS 0.035544f
C1133 VTAIL.n81 VSUBS 0.015922f
C1134 VTAIL.n82 VSUBS 0.015038f
C1135 VTAIL.n83 VSUBS 0.027985f
C1136 VTAIL.n84 VSUBS 0.027985f
C1137 VTAIL.n85 VSUBS 0.015038f
C1138 VTAIL.n86 VSUBS 0.015922f
C1139 VTAIL.n87 VSUBS 0.035544f
C1140 VTAIL.n88 VSUBS 0.086457f
C1141 VTAIL.n89 VSUBS 0.015922f
C1142 VTAIL.n90 VSUBS 0.015038f
C1143 VTAIL.n91 VSUBS 0.068508f
C1144 VTAIL.n92 VSUBS 0.043611f
C1145 VTAIL.n93 VSUBS 1.99821f
C1146 VTAIL.n94 VSUBS 0.030869f
C1147 VTAIL.n95 VSUBS 0.027985f
C1148 VTAIL.n96 VSUBS 0.015038f
C1149 VTAIL.n97 VSUBS 0.035544f
C1150 VTAIL.n98 VSUBS 0.015922f
C1151 VTAIL.n99 VSUBS 0.027985f
C1152 VTAIL.n100 VSUBS 0.015038f
C1153 VTAIL.n101 VSUBS 0.035544f
C1154 VTAIL.n102 VSUBS 0.015922f
C1155 VTAIL.n103 VSUBS 0.027985f
C1156 VTAIL.n104 VSUBS 0.015038f
C1157 VTAIL.n105 VSUBS 0.035544f
C1158 VTAIL.n106 VSUBS 0.035544f
C1159 VTAIL.n107 VSUBS 0.015922f
C1160 VTAIL.n108 VSUBS 0.027985f
C1161 VTAIL.n109 VSUBS 0.015038f
C1162 VTAIL.n110 VSUBS 0.035544f
C1163 VTAIL.n111 VSUBS 0.015922f
C1164 VTAIL.n112 VSUBS 0.027985f
C1165 VTAIL.n113 VSUBS 0.015038f
C1166 VTAIL.n114 VSUBS 0.035544f
C1167 VTAIL.n115 VSUBS 0.015922f
C1168 VTAIL.n116 VSUBS 0.027985f
C1169 VTAIL.n117 VSUBS 0.015038f
C1170 VTAIL.n118 VSUBS 0.035544f
C1171 VTAIL.n119 VSUBS 0.015922f
C1172 VTAIL.n120 VSUBS 0.027985f
C1173 VTAIL.n121 VSUBS 0.015038f
C1174 VTAIL.n122 VSUBS 0.035544f
C1175 VTAIL.n123 VSUBS 0.015922f
C1176 VTAIL.n124 VSUBS 0.21295f
C1177 VTAIL.t1 VSUBS 0.076224f
C1178 VTAIL.n125 VSUBS 0.026658f
C1179 VTAIL.n126 VSUBS 0.022611f
C1180 VTAIL.n127 VSUBS 0.015038f
C1181 VTAIL.n128 VSUBS 2.02826f
C1182 VTAIL.n129 VSUBS 0.027985f
C1183 VTAIL.n130 VSUBS 0.015038f
C1184 VTAIL.n131 VSUBS 0.015922f
C1185 VTAIL.n132 VSUBS 0.035544f
C1186 VTAIL.n133 VSUBS 0.035544f
C1187 VTAIL.n134 VSUBS 0.015922f
C1188 VTAIL.n135 VSUBS 0.015038f
C1189 VTAIL.n136 VSUBS 0.027985f
C1190 VTAIL.n137 VSUBS 0.027985f
C1191 VTAIL.n138 VSUBS 0.015038f
C1192 VTAIL.n139 VSUBS 0.015922f
C1193 VTAIL.n140 VSUBS 0.035544f
C1194 VTAIL.n141 VSUBS 0.035544f
C1195 VTAIL.n142 VSUBS 0.015922f
C1196 VTAIL.n143 VSUBS 0.015038f
C1197 VTAIL.n144 VSUBS 0.027985f
C1198 VTAIL.n145 VSUBS 0.027985f
C1199 VTAIL.n146 VSUBS 0.015038f
C1200 VTAIL.n147 VSUBS 0.015922f
C1201 VTAIL.n148 VSUBS 0.035544f
C1202 VTAIL.n149 VSUBS 0.035544f
C1203 VTAIL.n150 VSUBS 0.015922f
C1204 VTAIL.n151 VSUBS 0.015038f
C1205 VTAIL.n152 VSUBS 0.027985f
C1206 VTAIL.n153 VSUBS 0.027985f
C1207 VTAIL.n154 VSUBS 0.015038f
C1208 VTAIL.n155 VSUBS 0.015922f
C1209 VTAIL.n156 VSUBS 0.035544f
C1210 VTAIL.n157 VSUBS 0.035544f
C1211 VTAIL.n158 VSUBS 0.015922f
C1212 VTAIL.n159 VSUBS 0.015038f
C1213 VTAIL.n160 VSUBS 0.027985f
C1214 VTAIL.n161 VSUBS 0.027985f
C1215 VTAIL.n162 VSUBS 0.015038f
C1216 VTAIL.n163 VSUBS 0.015922f
C1217 VTAIL.n164 VSUBS 0.035544f
C1218 VTAIL.n165 VSUBS 0.035544f
C1219 VTAIL.n166 VSUBS 0.015922f
C1220 VTAIL.n167 VSUBS 0.015038f
C1221 VTAIL.n168 VSUBS 0.027985f
C1222 VTAIL.n169 VSUBS 0.027985f
C1223 VTAIL.n170 VSUBS 0.015038f
C1224 VTAIL.n171 VSUBS 0.01548f
C1225 VTAIL.n172 VSUBS 0.01548f
C1226 VTAIL.n173 VSUBS 0.035544f
C1227 VTAIL.n174 VSUBS 0.035544f
C1228 VTAIL.n175 VSUBS 0.015922f
C1229 VTAIL.n176 VSUBS 0.015038f
C1230 VTAIL.n177 VSUBS 0.027985f
C1231 VTAIL.n178 VSUBS 0.027985f
C1232 VTAIL.n179 VSUBS 0.015038f
C1233 VTAIL.n180 VSUBS 0.015922f
C1234 VTAIL.n181 VSUBS 0.035544f
C1235 VTAIL.n182 VSUBS 0.086457f
C1236 VTAIL.n183 VSUBS 0.015922f
C1237 VTAIL.n184 VSUBS 0.015038f
C1238 VTAIL.n185 VSUBS 0.068508f
C1239 VTAIL.n186 VSUBS 0.043611f
C1240 VTAIL.n187 VSUBS 2.01843f
C1241 VTAIL.n188 VSUBS 0.030869f
C1242 VTAIL.n189 VSUBS 0.027985f
C1243 VTAIL.n190 VSUBS 0.015038f
C1244 VTAIL.n191 VSUBS 0.035544f
C1245 VTAIL.n192 VSUBS 0.015922f
C1246 VTAIL.n193 VSUBS 0.027985f
C1247 VTAIL.n194 VSUBS 0.015038f
C1248 VTAIL.n195 VSUBS 0.035544f
C1249 VTAIL.n196 VSUBS 0.015922f
C1250 VTAIL.n197 VSUBS 0.027985f
C1251 VTAIL.n198 VSUBS 0.015038f
C1252 VTAIL.n199 VSUBS 0.035544f
C1253 VTAIL.n200 VSUBS 0.035544f
C1254 VTAIL.n201 VSUBS 0.015922f
C1255 VTAIL.n202 VSUBS 0.027985f
C1256 VTAIL.n203 VSUBS 0.015038f
C1257 VTAIL.n204 VSUBS 0.035544f
C1258 VTAIL.n205 VSUBS 0.015922f
C1259 VTAIL.n206 VSUBS 0.027985f
C1260 VTAIL.n207 VSUBS 0.015038f
C1261 VTAIL.n208 VSUBS 0.035544f
C1262 VTAIL.n209 VSUBS 0.015922f
C1263 VTAIL.n210 VSUBS 0.027985f
C1264 VTAIL.n211 VSUBS 0.015038f
C1265 VTAIL.n212 VSUBS 0.035544f
C1266 VTAIL.n213 VSUBS 0.015922f
C1267 VTAIL.n214 VSUBS 0.027985f
C1268 VTAIL.n215 VSUBS 0.015038f
C1269 VTAIL.n216 VSUBS 0.035544f
C1270 VTAIL.n217 VSUBS 0.015922f
C1271 VTAIL.n218 VSUBS 0.21295f
C1272 VTAIL.t2 VSUBS 0.076224f
C1273 VTAIL.n219 VSUBS 0.026658f
C1274 VTAIL.n220 VSUBS 0.022611f
C1275 VTAIL.n221 VSUBS 0.015038f
C1276 VTAIL.n222 VSUBS 2.02826f
C1277 VTAIL.n223 VSUBS 0.027985f
C1278 VTAIL.n224 VSUBS 0.015038f
C1279 VTAIL.n225 VSUBS 0.015922f
C1280 VTAIL.n226 VSUBS 0.035544f
C1281 VTAIL.n227 VSUBS 0.035544f
C1282 VTAIL.n228 VSUBS 0.015922f
C1283 VTAIL.n229 VSUBS 0.015038f
C1284 VTAIL.n230 VSUBS 0.027985f
C1285 VTAIL.n231 VSUBS 0.027985f
C1286 VTAIL.n232 VSUBS 0.015038f
C1287 VTAIL.n233 VSUBS 0.015922f
C1288 VTAIL.n234 VSUBS 0.035544f
C1289 VTAIL.n235 VSUBS 0.035544f
C1290 VTAIL.n236 VSUBS 0.015922f
C1291 VTAIL.n237 VSUBS 0.015038f
C1292 VTAIL.n238 VSUBS 0.027985f
C1293 VTAIL.n239 VSUBS 0.027985f
C1294 VTAIL.n240 VSUBS 0.015038f
C1295 VTAIL.n241 VSUBS 0.015922f
C1296 VTAIL.n242 VSUBS 0.035544f
C1297 VTAIL.n243 VSUBS 0.035544f
C1298 VTAIL.n244 VSUBS 0.015922f
C1299 VTAIL.n245 VSUBS 0.015038f
C1300 VTAIL.n246 VSUBS 0.027985f
C1301 VTAIL.n247 VSUBS 0.027985f
C1302 VTAIL.n248 VSUBS 0.015038f
C1303 VTAIL.n249 VSUBS 0.015922f
C1304 VTAIL.n250 VSUBS 0.035544f
C1305 VTAIL.n251 VSUBS 0.035544f
C1306 VTAIL.n252 VSUBS 0.015922f
C1307 VTAIL.n253 VSUBS 0.015038f
C1308 VTAIL.n254 VSUBS 0.027985f
C1309 VTAIL.n255 VSUBS 0.027985f
C1310 VTAIL.n256 VSUBS 0.015038f
C1311 VTAIL.n257 VSUBS 0.015922f
C1312 VTAIL.n258 VSUBS 0.035544f
C1313 VTAIL.n259 VSUBS 0.035544f
C1314 VTAIL.n260 VSUBS 0.015922f
C1315 VTAIL.n261 VSUBS 0.015038f
C1316 VTAIL.n262 VSUBS 0.027985f
C1317 VTAIL.n263 VSUBS 0.027985f
C1318 VTAIL.n264 VSUBS 0.015038f
C1319 VTAIL.n265 VSUBS 0.01548f
C1320 VTAIL.n266 VSUBS 0.01548f
C1321 VTAIL.n267 VSUBS 0.035544f
C1322 VTAIL.n268 VSUBS 0.035544f
C1323 VTAIL.n269 VSUBS 0.015922f
C1324 VTAIL.n270 VSUBS 0.015038f
C1325 VTAIL.n271 VSUBS 0.027985f
C1326 VTAIL.n272 VSUBS 0.027985f
C1327 VTAIL.n273 VSUBS 0.015038f
C1328 VTAIL.n274 VSUBS 0.015922f
C1329 VTAIL.n275 VSUBS 0.035544f
C1330 VTAIL.n276 VSUBS 0.086457f
C1331 VTAIL.n277 VSUBS 0.015922f
C1332 VTAIL.n278 VSUBS 0.015038f
C1333 VTAIL.n279 VSUBS 0.068508f
C1334 VTAIL.n280 VSUBS 0.043611f
C1335 VTAIL.n281 VSUBS 1.91659f
C1336 VTAIL.n282 VSUBS 0.030869f
C1337 VTAIL.n283 VSUBS 0.027985f
C1338 VTAIL.n284 VSUBS 0.015038f
C1339 VTAIL.n285 VSUBS 0.035544f
C1340 VTAIL.n286 VSUBS 0.015922f
C1341 VTAIL.n287 VSUBS 0.027985f
C1342 VTAIL.n288 VSUBS 0.015038f
C1343 VTAIL.n289 VSUBS 0.035544f
C1344 VTAIL.n290 VSUBS 0.015922f
C1345 VTAIL.n291 VSUBS 0.027985f
C1346 VTAIL.n292 VSUBS 0.015038f
C1347 VTAIL.n293 VSUBS 0.035544f
C1348 VTAIL.n294 VSUBS 0.015922f
C1349 VTAIL.n295 VSUBS 0.027985f
C1350 VTAIL.n296 VSUBS 0.015038f
C1351 VTAIL.n297 VSUBS 0.035544f
C1352 VTAIL.n298 VSUBS 0.015922f
C1353 VTAIL.n299 VSUBS 0.027985f
C1354 VTAIL.n300 VSUBS 0.015038f
C1355 VTAIL.n301 VSUBS 0.035544f
C1356 VTAIL.n302 VSUBS 0.015922f
C1357 VTAIL.n303 VSUBS 0.027985f
C1358 VTAIL.n304 VSUBS 0.015038f
C1359 VTAIL.n305 VSUBS 0.035544f
C1360 VTAIL.n306 VSUBS 0.015922f
C1361 VTAIL.n307 VSUBS 0.027985f
C1362 VTAIL.n308 VSUBS 0.015038f
C1363 VTAIL.n309 VSUBS 0.035544f
C1364 VTAIL.n310 VSUBS 0.015922f
C1365 VTAIL.n311 VSUBS 0.21295f
C1366 VTAIL.t0 VSUBS 0.076224f
C1367 VTAIL.n312 VSUBS 0.026658f
C1368 VTAIL.n313 VSUBS 0.022611f
C1369 VTAIL.n314 VSUBS 0.015038f
C1370 VTAIL.n315 VSUBS 2.02826f
C1371 VTAIL.n316 VSUBS 0.027985f
C1372 VTAIL.n317 VSUBS 0.015038f
C1373 VTAIL.n318 VSUBS 0.015922f
C1374 VTAIL.n319 VSUBS 0.035544f
C1375 VTAIL.n320 VSUBS 0.035544f
C1376 VTAIL.n321 VSUBS 0.015922f
C1377 VTAIL.n322 VSUBS 0.015038f
C1378 VTAIL.n323 VSUBS 0.027985f
C1379 VTAIL.n324 VSUBS 0.027985f
C1380 VTAIL.n325 VSUBS 0.015038f
C1381 VTAIL.n326 VSUBS 0.015922f
C1382 VTAIL.n327 VSUBS 0.035544f
C1383 VTAIL.n328 VSUBS 0.035544f
C1384 VTAIL.n329 VSUBS 0.015922f
C1385 VTAIL.n330 VSUBS 0.015038f
C1386 VTAIL.n331 VSUBS 0.027985f
C1387 VTAIL.n332 VSUBS 0.027985f
C1388 VTAIL.n333 VSUBS 0.015038f
C1389 VTAIL.n334 VSUBS 0.015922f
C1390 VTAIL.n335 VSUBS 0.035544f
C1391 VTAIL.n336 VSUBS 0.035544f
C1392 VTAIL.n337 VSUBS 0.015922f
C1393 VTAIL.n338 VSUBS 0.015038f
C1394 VTAIL.n339 VSUBS 0.027985f
C1395 VTAIL.n340 VSUBS 0.027985f
C1396 VTAIL.n341 VSUBS 0.015038f
C1397 VTAIL.n342 VSUBS 0.015922f
C1398 VTAIL.n343 VSUBS 0.035544f
C1399 VTAIL.n344 VSUBS 0.035544f
C1400 VTAIL.n345 VSUBS 0.015922f
C1401 VTAIL.n346 VSUBS 0.015038f
C1402 VTAIL.n347 VSUBS 0.027985f
C1403 VTAIL.n348 VSUBS 0.027985f
C1404 VTAIL.n349 VSUBS 0.015038f
C1405 VTAIL.n350 VSUBS 0.015922f
C1406 VTAIL.n351 VSUBS 0.035544f
C1407 VTAIL.n352 VSUBS 0.035544f
C1408 VTAIL.n353 VSUBS 0.035544f
C1409 VTAIL.n354 VSUBS 0.015922f
C1410 VTAIL.n355 VSUBS 0.015038f
C1411 VTAIL.n356 VSUBS 0.027985f
C1412 VTAIL.n357 VSUBS 0.027985f
C1413 VTAIL.n358 VSUBS 0.015038f
C1414 VTAIL.n359 VSUBS 0.01548f
C1415 VTAIL.n360 VSUBS 0.01548f
C1416 VTAIL.n361 VSUBS 0.035544f
C1417 VTAIL.n362 VSUBS 0.035544f
C1418 VTAIL.n363 VSUBS 0.015922f
C1419 VTAIL.n364 VSUBS 0.015038f
C1420 VTAIL.n365 VSUBS 0.027985f
C1421 VTAIL.n366 VSUBS 0.027985f
C1422 VTAIL.n367 VSUBS 0.015038f
C1423 VTAIL.n368 VSUBS 0.015922f
C1424 VTAIL.n369 VSUBS 0.035544f
C1425 VTAIL.n370 VSUBS 0.086457f
C1426 VTAIL.n371 VSUBS 0.015922f
C1427 VTAIL.n372 VSUBS 0.015038f
C1428 VTAIL.n373 VSUBS 0.068508f
C1429 VTAIL.n374 VSUBS 0.043611f
C1430 VTAIL.n375 VSUBS 1.84352f
C1431 VP.t0 VSUBS 3.35318f
C1432 VP.t1 VSUBS 3.11939f
C1433 VP.n0 VSUBS 6.79593f
.ends

