* NGSPICE file created from diff_pair_sample_1748.ext - technology: sky130A

.subckt diff_pair_sample_1748 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=5.6394 pd=29.7 as=0 ps=0 w=14.46 l=0.57
X1 VDD1.t1 VP.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=5.6394 pd=29.7 as=5.6394 ps=29.7 w=14.46 l=0.57
X2 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.6394 pd=29.7 as=5.6394 ps=29.7 w=14.46 l=0.57
X3 VDD1.t0 VP.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=5.6394 pd=29.7 as=5.6394 ps=29.7 w=14.46 l=0.57
X4 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=5.6394 pd=29.7 as=0 ps=0 w=14.46 l=0.57
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.6394 pd=29.7 as=0 ps=0 w=14.46 l=0.57
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=5.6394 pd=29.7 as=0 ps=0 w=14.46 l=0.57
X7 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.6394 pd=29.7 as=5.6394 ps=29.7 w=14.46 l=0.57
R0 B.n86 B.t2 816.308
R1 B.n83 B.t13 816.308
R2 B.n381 B.t10 816.308
R3 B.n378 B.t6 816.308
R4 B.n656 B.n655 585
R5 B.n657 B.n656 585
R6 B.n299 B.n82 585
R7 B.n298 B.n297 585
R8 B.n296 B.n295 585
R9 B.n294 B.n293 585
R10 B.n292 B.n291 585
R11 B.n290 B.n289 585
R12 B.n288 B.n287 585
R13 B.n286 B.n285 585
R14 B.n284 B.n283 585
R15 B.n282 B.n281 585
R16 B.n280 B.n279 585
R17 B.n278 B.n277 585
R18 B.n276 B.n275 585
R19 B.n274 B.n273 585
R20 B.n272 B.n271 585
R21 B.n270 B.n269 585
R22 B.n268 B.n267 585
R23 B.n266 B.n265 585
R24 B.n264 B.n263 585
R25 B.n262 B.n261 585
R26 B.n260 B.n259 585
R27 B.n258 B.n257 585
R28 B.n256 B.n255 585
R29 B.n254 B.n253 585
R30 B.n252 B.n251 585
R31 B.n250 B.n249 585
R32 B.n248 B.n247 585
R33 B.n246 B.n245 585
R34 B.n244 B.n243 585
R35 B.n242 B.n241 585
R36 B.n240 B.n239 585
R37 B.n238 B.n237 585
R38 B.n236 B.n235 585
R39 B.n234 B.n233 585
R40 B.n232 B.n231 585
R41 B.n230 B.n229 585
R42 B.n228 B.n227 585
R43 B.n226 B.n225 585
R44 B.n224 B.n223 585
R45 B.n222 B.n221 585
R46 B.n220 B.n219 585
R47 B.n218 B.n217 585
R48 B.n216 B.n215 585
R49 B.n214 B.n213 585
R50 B.n212 B.n211 585
R51 B.n210 B.n209 585
R52 B.n208 B.n207 585
R53 B.n206 B.n205 585
R54 B.n204 B.n203 585
R55 B.n202 B.n201 585
R56 B.n200 B.n199 585
R57 B.n198 B.n197 585
R58 B.n196 B.n195 585
R59 B.n194 B.n193 585
R60 B.n192 B.n191 585
R61 B.n190 B.n189 585
R62 B.n188 B.n187 585
R63 B.n185 B.n184 585
R64 B.n183 B.n182 585
R65 B.n181 B.n180 585
R66 B.n179 B.n178 585
R67 B.n177 B.n176 585
R68 B.n175 B.n174 585
R69 B.n173 B.n172 585
R70 B.n171 B.n170 585
R71 B.n169 B.n168 585
R72 B.n167 B.n166 585
R73 B.n165 B.n164 585
R74 B.n163 B.n162 585
R75 B.n161 B.n160 585
R76 B.n159 B.n158 585
R77 B.n157 B.n156 585
R78 B.n155 B.n154 585
R79 B.n153 B.n152 585
R80 B.n151 B.n150 585
R81 B.n149 B.n148 585
R82 B.n147 B.n146 585
R83 B.n145 B.n144 585
R84 B.n143 B.n142 585
R85 B.n141 B.n140 585
R86 B.n139 B.n138 585
R87 B.n137 B.n136 585
R88 B.n135 B.n134 585
R89 B.n133 B.n132 585
R90 B.n131 B.n130 585
R91 B.n129 B.n128 585
R92 B.n127 B.n126 585
R93 B.n125 B.n124 585
R94 B.n123 B.n122 585
R95 B.n121 B.n120 585
R96 B.n119 B.n118 585
R97 B.n117 B.n116 585
R98 B.n115 B.n114 585
R99 B.n113 B.n112 585
R100 B.n111 B.n110 585
R101 B.n109 B.n108 585
R102 B.n107 B.n106 585
R103 B.n105 B.n104 585
R104 B.n103 B.n102 585
R105 B.n101 B.n100 585
R106 B.n99 B.n98 585
R107 B.n97 B.n96 585
R108 B.n95 B.n94 585
R109 B.n93 B.n92 585
R110 B.n91 B.n90 585
R111 B.n89 B.n88 585
R112 B.n654 B.n28 585
R113 B.n658 B.n28 585
R114 B.n653 B.n27 585
R115 B.n659 B.n27 585
R116 B.n652 B.n651 585
R117 B.n651 B.n23 585
R118 B.n650 B.n22 585
R119 B.n665 B.n22 585
R120 B.n649 B.n21 585
R121 B.n666 B.n21 585
R122 B.n648 B.n20 585
R123 B.n667 B.n20 585
R124 B.n647 B.n646 585
R125 B.n646 B.n16 585
R126 B.n645 B.n15 585
R127 B.n673 B.n15 585
R128 B.n644 B.n14 585
R129 B.n674 B.n14 585
R130 B.n643 B.n13 585
R131 B.n675 B.n13 585
R132 B.n642 B.n641 585
R133 B.n641 B.n12 585
R134 B.n640 B.n639 585
R135 B.n640 B.n8 585
R136 B.n638 B.n7 585
R137 B.n682 B.n7 585
R138 B.n637 B.n6 585
R139 B.n683 B.n6 585
R140 B.n636 B.n5 585
R141 B.n684 B.n5 585
R142 B.n635 B.n634 585
R143 B.n634 B.n4 585
R144 B.n633 B.n300 585
R145 B.n633 B.n632 585
R146 B.n622 B.n301 585
R147 B.n625 B.n301 585
R148 B.n624 B.n623 585
R149 B.n626 B.n624 585
R150 B.n621 B.n306 585
R151 B.n306 B.n305 585
R152 B.n620 B.n619 585
R153 B.n619 B.n618 585
R154 B.n308 B.n307 585
R155 B.n309 B.n308 585
R156 B.n611 B.n610 585
R157 B.n612 B.n611 585
R158 B.n609 B.n313 585
R159 B.n317 B.n313 585
R160 B.n608 B.n607 585
R161 B.n607 B.n606 585
R162 B.n315 B.n314 585
R163 B.n316 B.n315 585
R164 B.n599 B.n598 585
R165 B.n600 B.n599 585
R166 B.n597 B.n322 585
R167 B.n322 B.n321 585
R168 B.n591 B.n590 585
R169 B.n589 B.n377 585
R170 B.n588 B.n376 585
R171 B.n593 B.n376 585
R172 B.n587 B.n586 585
R173 B.n585 B.n584 585
R174 B.n583 B.n582 585
R175 B.n581 B.n580 585
R176 B.n579 B.n578 585
R177 B.n577 B.n576 585
R178 B.n575 B.n574 585
R179 B.n573 B.n572 585
R180 B.n571 B.n570 585
R181 B.n569 B.n568 585
R182 B.n567 B.n566 585
R183 B.n565 B.n564 585
R184 B.n563 B.n562 585
R185 B.n561 B.n560 585
R186 B.n559 B.n558 585
R187 B.n557 B.n556 585
R188 B.n555 B.n554 585
R189 B.n553 B.n552 585
R190 B.n551 B.n550 585
R191 B.n549 B.n548 585
R192 B.n547 B.n546 585
R193 B.n545 B.n544 585
R194 B.n543 B.n542 585
R195 B.n541 B.n540 585
R196 B.n539 B.n538 585
R197 B.n537 B.n536 585
R198 B.n535 B.n534 585
R199 B.n533 B.n532 585
R200 B.n531 B.n530 585
R201 B.n529 B.n528 585
R202 B.n527 B.n526 585
R203 B.n525 B.n524 585
R204 B.n523 B.n522 585
R205 B.n521 B.n520 585
R206 B.n519 B.n518 585
R207 B.n517 B.n516 585
R208 B.n515 B.n514 585
R209 B.n513 B.n512 585
R210 B.n511 B.n510 585
R211 B.n509 B.n508 585
R212 B.n507 B.n506 585
R213 B.n505 B.n504 585
R214 B.n503 B.n502 585
R215 B.n501 B.n500 585
R216 B.n499 B.n498 585
R217 B.n497 B.n496 585
R218 B.n495 B.n494 585
R219 B.n493 B.n492 585
R220 B.n491 B.n490 585
R221 B.n489 B.n488 585
R222 B.n487 B.n486 585
R223 B.n485 B.n484 585
R224 B.n483 B.n482 585
R225 B.n481 B.n480 585
R226 B.n479 B.n478 585
R227 B.n476 B.n475 585
R228 B.n474 B.n473 585
R229 B.n472 B.n471 585
R230 B.n470 B.n469 585
R231 B.n468 B.n467 585
R232 B.n466 B.n465 585
R233 B.n464 B.n463 585
R234 B.n462 B.n461 585
R235 B.n460 B.n459 585
R236 B.n458 B.n457 585
R237 B.n456 B.n455 585
R238 B.n454 B.n453 585
R239 B.n452 B.n451 585
R240 B.n450 B.n449 585
R241 B.n448 B.n447 585
R242 B.n446 B.n445 585
R243 B.n444 B.n443 585
R244 B.n442 B.n441 585
R245 B.n440 B.n439 585
R246 B.n438 B.n437 585
R247 B.n436 B.n435 585
R248 B.n434 B.n433 585
R249 B.n432 B.n431 585
R250 B.n430 B.n429 585
R251 B.n428 B.n427 585
R252 B.n426 B.n425 585
R253 B.n424 B.n423 585
R254 B.n422 B.n421 585
R255 B.n420 B.n419 585
R256 B.n418 B.n417 585
R257 B.n416 B.n415 585
R258 B.n414 B.n413 585
R259 B.n412 B.n411 585
R260 B.n410 B.n409 585
R261 B.n408 B.n407 585
R262 B.n406 B.n405 585
R263 B.n404 B.n403 585
R264 B.n402 B.n401 585
R265 B.n400 B.n399 585
R266 B.n398 B.n397 585
R267 B.n396 B.n395 585
R268 B.n394 B.n393 585
R269 B.n392 B.n391 585
R270 B.n390 B.n389 585
R271 B.n388 B.n387 585
R272 B.n386 B.n385 585
R273 B.n384 B.n383 585
R274 B.n324 B.n323 585
R275 B.n596 B.n595 585
R276 B.n320 B.n319 585
R277 B.n321 B.n320 585
R278 B.n602 B.n601 585
R279 B.n601 B.n600 585
R280 B.n603 B.n318 585
R281 B.n318 B.n316 585
R282 B.n605 B.n604 585
R283 B.n606 B.n605 585
R284 B.n312 B.n311 585
R285 B.n317 B.n312 585
R286 B.n614 B.n613 585
R287 B.n613 B.n612 585
R288 B.n615 B.n310 585
R289 B.n310 B.n309 585
R290 B.n617 B.n616 585
R291 B.n618 B.n617 585
R292 B.n304 B.n303 585
R293 B.n305 B.n304 585
R294 B.n628 B.n627 585
R295 B.n627 B.n626 585
R296 B.n629 B.n302 585
R297 B.n625 B.n302 585
R298 B.n631 B.n630 585
R299 B.n632 B.n631 585
R300 B.n3 B.n0 585
R301 B.n4 B.n3 585
R302 B.n681 B.n1 585
R303 B.n682 B.n681 585
R304 B.n680 B.n679 585
R305 B.n680 B.n8 585
R306 B.n678 B.n9 585
R307 B.n12 B.n9 585
R308 B.n677 B.n676 585
R309 B.n676 B.n675 585
R310 B.n11 B.n10 585
R311 B.n674 B.n11 585
R312 B.n672 B.n671 585
R313 B.n673 B.n672 585
R314 B.n670 B.n17 585
R315 B.n17 B.n16 585
R316 B.n669 B.n668 585
R317 B.n668 B.n667 585
R318 B.n19 B.n18 585
R319 B.n666 B.n19 585
R320 B.n664 B.n663 585
R321 B.n665 B.n664 585
R322 B.n662 B.n24 585
R323 B.n24 B.n23 585
R324 B.n661 B.n660 585
R325 B.n660 B.n659 585
R326 B.n26 B.n25 585
R327 B.n658 B.n26 585
R328 B.n685 B.n684 585
R329 B.n683 B.n2 585
R330 B.n88 B.n26 516.524
R331 B.n656 B.n28 516.524
R332 B.n595 B.n322 516.524
R333 B.n591 B.n320 516.524
R334 B.n657 B.n81 256.663
R335 B.n657 B.n80 256.663
R336 B.n657 B.n79 256.663
R337 B.n657 B.n78 256.663
R338 B.n657 B.n77 256.663
R339 B.n657 B.n76 256.663
R340 B.n657 B.n75 256.663
R341 B.n657 B.n74 256.663
R342 B.n657 B.n73 256.663
R343 B.n657 B.n72 256.663
R344 B.n657 B.n71 256.663
R345 B.n657 B.n70 256.663
R346 B.n657 B.n69 256.663
R347 B.n657 B.n68 256.663
R348 B.n657 B.n67 256.663
R349 B.n657 B.n66 256.663
R350 B.n657 B.n65 256.663
R351 B.n657 B.n64 256.663
R352 B.n657 B.n63 256.663
R353 B.n657 B.n62 256.663
R354 B.n657 B.n61 256.663
R355 B.n657 B.n60 256.663
R356 B.n657 B.n59 256.663
R357 B.n657 B.n58 256.663
R358 B.n657 B.n57 256.663
R359 B.n657 B.n56 256.663
R360 B.n657 B.n55 256.663
R361 B.n657 B.n54 256.663
R362 B.n657 B.n53 256.663
R363 B.n657 B.n52 256.663
R364 B.n657 B.n51 256.663
R365 B.n657 B.n50 256.663
R366 B.n657 B.n49 256.663
R367 B.n657 B.n48 256.663
R368 B.n657 B.n47 256.663
R369 B.n657 B.n46 256.663
R370 B.n657 B.n45 256.663
R371 B.n657 B.n44 256.663
R372 B.n657 B.n43 256.663
R373 B.n657 B.n42 256.663
R374 B.n657 B.n41 256.663
R375 B.n657 B.n40 256.663
R376 B.n657 B.n39 256.663
R377 B.n657 B.n38 256.663
R378 B.n657 B.n37 256.663
R379 B.n657 B.n36 256.663
R380 B.n657 B.n35 256.663
R381 B.n657 B.n34 256.663
R382 B.n657 B.n33 256.663
R383 B.n657 B.n32 256.663
R384 B.n657 B.n31 256.663
R385 B.n657 B.n30 256.663
R386 B.n657 B.n29 256.663
R387 B.n593 B.n592 256.663
R388 B.n593 B.n325 256.663
R389 B.n593 B.n326 256.663
R390 B.n593 B.n327 256.663
R391 B.n593 B.n328 256.663
R392 B.n593 B.n329 256.663
R393 B.n593 B.n330 256.663
R394 B.n593 B.n331 256.663
R395 B.n593 B.n332 256.663
R396 B.n593 B.n333 256.663
R397 B.n593 B.n334 256.663
R398 B.n593 B.n335 256.663
R399 B.n593 B.n336 256.663
R400 B.n593 B.n337 256.663
R401 B.n593 B.n338 256.663
R402 B.n593 B.n339 256.663
R403 B.n593 B.n340 256.663
R404 B.n593 B.n341 256.663
R405 B.n593 B.n342 256.663
R406 B.n593 B.n343 256.663
R407 B.n593 B.n344 256.663
R408 B.n593 B.n345 256.663
R409 B.n593 B.n346 256.663
R410 B.n593 B.n347 256.663
R411 B.n593 B.n348 256.663
R412 B.n593 B.n349 256.663
R413 B.n593 B.n350 256.663
R414 B.n593 B.n351 256.663
R415 B.n593 B.n352 256.663
R416 B.n593 B.n353 256.663
R417 B.n593 B.n354 256.663
R418 B.n593 B.n355 256.663
R419 B.n593 B.n356 256.663
R420 B.n593 B.n357 256.663
R421 B.n593 B.n358 256.663
R422 B.n593 B.n359 256.663
R423 B.n593 B.n360 256.663
R424 B.n593 B.n361 256.663
R425 B.n593 B.n362 256.663
R426 B.n593 B.n363 256.663
R427 B.n593 B.n364 256.663
R428 B.n593 B.n365 256.663
R429 B.n593 B.n366 256.663
R430 B.n593 B.n367 256.663
R431 B.n593 B.n368 256.663
R432 B.n593 B.n369 256.663
R433 B.n593 B.n370 256.663
R434 B.n593 B.n371 256.663
R435 B.n593 B.n372 256.663
R436 B.n593 B.n373 256.663
R437 B.n593 B.n374 256.663
R438 B.n593 B.n375 256.663
R439 B.n594 B.n593 256.663
R440 B.n687 B.n686 256.663
R441 B.n92 B.n91 163.367
R442 B.n96 B.n95 163.367
R443 B.n100 B.n99 163.367
R444 B.n104 B.n103 163.367
R445 B.n108 B.n107 163.367
R446 B.n112 B.n111 163.367
R447 B.n116 B.n115 163.367
R448 B.n120 B.n119 163.367
R449 B.n124 B.n123 163.367
R450 B.n128 B.n127 163.367
R451 B.n132 B.n131 163.367
R452 B.n136 B.n135 163.367
R453 B.n140 B.n139 163.367
R454 B.n144 B.n143 163.367
R455 B.n148 B.n147 163.367
R456 B.n152 B.n151 163.367
R457 B.n156 B.n155 163.367
R458 B.n160 B.n159 163.367
R459 B.n164 B.n163 163.367
R460 B.n168 B.n167 163.367
R461 B.n172 B.n171 163.367
R462 B.n176 B.n175 163.367
R463 B.n180 B.n179 163.367
R464 B.n184 B.n183 163.367
R465 B.n189 B.n188 163.367
R466 B.n193 B.n192 163.367
R467 B.n197 B.n196 163.367
R468 B.n201 B.n200 163.367
R469 B.n205 B.n204 163.367
R470 B.n209 B.n208 163.367
R471 B.n213 B.n212 163.367
R472 B.n217 B.n216 163.367
R473 B.n221 B.n220 163.367
R474 B.n225 B.n224 163.367
R475 B.n229 B.n228 163.367
R476 B.n233 B.n232 163.367
R477 B.n237 B.n236 163.367
R478 B.n241 B.n240 163.367
R479 B.n245 B.n244 163.367
R480 B.n249 B.n248 163.367
R481 B.n253 B.n252 163.367
R482 B.n257 B.n256 163.367
R483 B.n261 B.n260 163.367
R484 B.n265 B.n264 163.367
R485 B.n269 B.n268 163.367
R486 B.n273 B.n272 163.367
R487 B.n277 B.n276 163.367
R488 B.n281 B.n280 163.367
R489 B.n285 B.n284 163.367
R490 B.n289 B.n288 163.367
R491 B.n293 B.n292 163.367
R492 B.n297 B.n296 163.367
R493 B.n656 B.n82 163.367
R494 B.n599 B.n322 163.367
R495 B.n599 B.n315 163.367
R496 B.n607 B.n315 163.367
R497 B.n607 B.n313 163.367
R498 B.n611 B.n313 163.367
R499 B.n611 B.n308 163.367
R500 B.n619 B.n308 163.367
R501 B.n619 B.n306 163.367
R502 B.n624 B.n306 163.367
R503 B.n624 B.n301 163.367
R504 B.n633 B.n301 163.367
R505 B.n634 B.n633 163.367
R506 B.n634 B.n5 163.367
R507 B.n6 B.n5 163.367
R508 B.n7 B.n6 163.367
R509 B.n640 B.n7 163.367
R510 B.n641 B.n640 163.367
R511 B.n641 B.n13 163.367
R512 B.n14 B.n13 163.367
R513 B.n15 B.n14 163.367
R514 B.n646 B.n15 163.367
R515 B.n646 B.n20 163.367
R516 B.n21 B.n20 163.367
R517 B.n22 B.n21 163.367
R518 B.n651 B.n22 163.367
R519 B.n651 B.n27 163.367
R520 B.n28 B.n27 163.367
R521 B.n377 B.n376 163.367
R522 B.n586 B.n376 163.367
R523 B.n584 B.n583 163.367
R524 B.n580 B.n579 163.367
R525 B.n576 B.n575 163.367
R526 B.n572 B.n571 163.367
R527 B.n568 B.n567 163.367
R528 B.n564 B.n563 163.367
R529 B.n560 B.n559 163.367
R530 B.n556 B.n555 163.367
R531 B.n552 B.n551 163.367
R532 B.n548 B.n547 163.367
R533 B.n544 B.n543 163.367
R534 B.n540 B.n539 163.367
R535 B.n536 B.n535 163.367
R536 B.n532 B.n531 163.367
R537 B.n528 B.n527 163.367
R538 B.n524 B.n523 163.367
R539 B.n520 B.n519 163.367
R540 B.n516 B.n515 163.367
R541 B.n512 B.n511 163.367
R542 B.n508 B.n507 163.367
R543 B.n504 B.n503 163.367
R544 B.n500 B.n499 163.367
R545 B.n496 B.n495 163.367
R546 B.n492 B.n491 163.367
R547 B.n488 B.n487 163.367
R548 B.n484 B.n483 163.367
R549 B.n480 B.n479 163.367
R550 B.n475 B.n474 163.367
R551 B.n471 B.n470 163.367
R552 B.n467 B.n466 163.367
R553 B.n463 B.n462 163.367
R554 B.n459 B.n458 163.367
R555 B.n455 B.n454 163.367
R556 B.n451 B.n450 163.367
R557 B.n447 B.n446 163.367
R558 B.n443 B.n442 163.367
R559 B.n439 B.n438 163.367
R560 B.n435 B.n434 163.367
R561 B.n431 B.n430 163.367
R562 B.n427 B.n426 163.367
R563 B.n423 B.n422 163.367
R564 B.n419 B.n418 163.367
R565 B.n415 B.n414 163.367
R566 B.n411 B.n410 163.367
R567 B.n407 B.n406 163.367
R568 B.n403 B.n402 163.367
R569 B.n399 B.n398 163.367
R570 B.n395 B.n394 163.367
R571 B.n391 B.n390 163.367
R572 B.n387 B.n386 163.367
R573 B.n383 B.n324 163.367
R574 B.n601 B.n320 163.367
R575 B.n601 B.n318 163.367
R576 B.n605 B.n318 163.367
R577 B.n605 B.n312 163.367
R578 B.n613 B.n312 163.367
R579 B.n613 B.n310 163.367
R580 B.n617 B.n310 163.367
R581 B.n617 B.n304 163.367
R582 B.n627 B.n304 163.367
R583 B.n627 B.n302 163.367
R584 B.n631 B.n302 163.367
R585 B.n631 B.n3 163.367
R586 B.n685 B.n3 163.367
R587 B.n681 B.n2 163.367
R588 B.n681 B.n680 163.367
R589 B.n680 B.n9 163.367
R590 B.n676 B.n9 163.367
R591 B.n676 B.n11 163.367
R592 B.n672 B.n11 163.367
R593 B.n672 B.n17 163.367
R594 B.n668 B.n17 163.367
R595 B.n668 B.n19 163.367
R596 B.n664 B.n19 163.367
R597 B.n664 B.n24 163.367
R598 B.n660 B.n24 163.367
R599 B.n660 B.n26 163.367
R600 B.n83 B.t14 88.4581
R601 B.n381 B.t12 88.4581
R602 B.n86 B.t4 88.4394
R603 B.n378 B.t9 88.4394
R604 B.n88 B.n29 71.676
R605 B.n92 B.n30 71.676
R606 B.n96 B.n31 71.676
R607 B.n100 B.n32 71.676
R608 B.n104 B.n33 71.676
R609 B.n108 B.n34 71.676
R610 B.n112 B.n35 71.676
R611 B.n116 B.n36 71.676
R612 B.n120 B.n37 71.676
R613 B.n124 B.n38 71.676
R614 B.n128 B.n39 71.676
R615 B.n132 B.n40 71.676
R616 B.n136 B.n41 71.676
R617 B.n140 B.n42 71.676
R618 B.n144 B.n43 71.676
R619 B.n148 B.n44 71.676
R620 B.n152 B.n45 71.676
R621 B.n156 B.n46 71.676
R622 B.n160 B.n47 71.676
R623 B.n164 B.n48 71.676
R624 B.n168 B.n49 71.676
R625 B.n172 B.n50 71.676
R626 B.n176 B.n51 71.676
R627 B.n180 B.n52 71.676
R628 B.n184 B.n53 71.676
R629 B.n189 B.n54 71.676
R630 B.n193 B.n55 71.676
R631 B.n197 B.n56 71.676
R632 B.n201 B.n57 71.676
R633 B.n205 B.n58 71.676
R634 B.n209 B.n59 71.676
R635 B.n213 B.n60 71.676
R636 B.n217 B.n61 71.676
R637 B.n221 B.n62 71.676
R638 B.n225 B.n63 71.676
R639 B.n229 B.n64 71.676
R640 B.n233 B.n65 71.676
R641 B.n237 B.n66 71.676
R642 B.n241 B.n67 71.676
R643 B.n245 B.n68 71.676
R644 B.n249 B.n69 71.676
R645 B.n253 B.n70 71.676
R646 B.n257 B.n71 71.676
R647 B.n261 B.n72 71.676
R648 B.n265 B.n73 71.676
R649 B.n269 B.n74 71.676
R650 B.n273 B.n75 71.676
R651 B.n277 B.n76 71.676
R652 B.n281 B.n77 71.676
R653 B.n285 B.n78 71.676
R654 B.n289 B.n79 71.676
R655 B.n293 B.n80 71.676
R656 B.n297 B.n81 71.676
R657 B.n82 B.n81 71.676
R658 B.n296 B.n80 71.676
R659 B.n292 B.n79 71.676
R660 B.n288 B.n78 71.676
R661 B.n284 B.n77 71.676
R662 B.n280 B.n76 71.676
R663 B.n276 B.n75 71.676
R664 B.n272 B.n74 71.676
R665 B.n268 B.n73 71.676
R666 B.n264 B.n72 71.676
R667 B.n260 B.n71 71.676
R668 B.n256 B.n70 71.676
R669 B.n252 B.n69 71.676
R670 B.n248 B.n68 71.676
R671 B.n244 B.n67 71.676
R672 B.n240 B.n66 71.676
R673 B.n236 B.n65 71.676
R674 B.n232 B.n64 71.676
R675 B.n228 B.n63 71.676
R676 B.n224 B.n62 71.676
R677 B.n220 B.n61 71.676
R678 B.n216 B.n60 71.676
R679 B.n212 B.n59 71.676
R680 B.n208 B.n58 71.676
R681 B.n204 B.n57 71.676
R682 B.n200 B.n56 71.676
R683 B.n196 B.n55 71.676
R684 B.n192 B.n54 71.676
R685 B.n188 B.n53 71.676
R686 B.n183 B.n52 71.676
R687 B.n179 B.n51 71.676
R688 B.n175 B.n50 71.676
R689 B.n171 B.n49 71.676
R690 B.n167 B.n48 71.676
R691 B.n163 B.n47 71.676
R692 B.n159 B.n46 71.676
R693 B.n155 B.n45 71.676
R694 B.n151 B.n44 71.676
R695 B.n147 B.n43 71.676
R696 B.n143 B.n42 71.676
R697 B.n139 B.n41 71.676
R698 B.n135 B.n40 71.676
R699 B.n131 B.n39 71.676
R700 B.n127 B.n38 71.676
R701 B.n123 B.n37 71.676
R702 B.n119 B.n36 71.676
R703 B.n115 B.n35 71.676
R704 B.n111 B.n34 71.676
R705 B.n107 B.n33 71.676
R706 B.n103 B.n32 71.676
R707 B.n99 B.n31 71.676
R708 B.n95 B.n30 71.676
R709 B.n91 B.n29 71.676
R710 B.n592 B.n591 71.676
R711 B.n586 B.n325 71.676
R712 B.n583 B.n326 71.676
R713 B.n579 B.n327 71.676
R714 B.n575 B.n328 71.676
R715 B.n571 B.n329 71.676
R716 B.n567 B.n330 71.676
R717 B.n563 B.n331 71.676
R718 B.n559 B.n332 71.676
R719 B.n555 B.n333 71.676
R720 B.n551 B.n334 71.676
R721 B.n547 B.n335 71.676
R722 B.n543 B.n336 71.676
R723 B.n539 B.n337 71.676
R724 B.n535 B.n338 71.676
R725 B.n531 B.n339 71.676
R726 B.n527 B.n340 71.676
R727 B.n523 B.n341 71.676
R728 B.n519 B.n342 71.676
R729 B.n515 B.n343 71.676
R730 B.n511 B.n344 71.676
R731 B.n507 B.n345 71.676
R732 B.n503 B.n346 71.676
R733 B.n499 B.n347 71.676
R734 B.n495 B.n348 71.676
R735 B.n491 B.n349 71.676
R736 B.n487 B.n350 71.676
R737 B.n483 B.n351 71.676
R738 B.n479 B.n352 71.676
R739 B.n474 B.n353 71.676
R740 B.n470 B.n354 71.676
R741 B.n466 B.n355 71.676
R742 B.n462 B.n356 71.676
R743 B.n458 B.n357 71.676
R744 B.n454 B.n358 71.676
R745 B.n450 B.n359 71.676
R746 B.n446 B.n360 71.676
R747 B.n442 B.n361 71.676
R748 B.n438 B.n362 71.676
R749 B.n434 B.n363 71.676
R750 B.n430 B.n364 71.676
R751 B.n426 B.n365 71.676
R752 B.n422 B.n366 71.676
R753 B.n418 B.n367 71.676
R754 B.n414 B.n368 71.676
R755 B.n410 B.n369 71.676
R756 B.n406 B.n370 71.676
R757 B.n402 B.n371 71.676
R758 B.n398 B.n372 71.676
R759 B.n394 B.n373 71.676
R760 B.n390 B.n374 71.676
R761 B.n386 B.n375 71.676
R762 B.n594 B.n324 71.676
R763 B.n592 B.n377 71.676
R764 B.n584 B.n325 71.676
R765 B.n580 B.n326 71.676
R766 B.n576 B.n327 71.676
R767 B.n572 B.n328 71.676
R768 B.n568 B.n329 71.676
R769 B.n564 B.n330 71.676
R770 B.n560 B.n331 71.676
R771 B.n556 B.n332 71.676
R772 B.n552 B.n333 71.676
R773 B.n548 B.n334 71.676
R774 B.n544 B.n335 71.676
R775 B.n540 B.n336 71.676
R776 B.n536 B.n337 71.676
R777 B.n532 B.n338 71.676
R778 B.n528 B.n339 71.676
R779 B.n524 B.n340 71.676
R780 B.n520 B.n341 71.676
R781 B.n516 B.n342 71.676
R782 B.n512 B.n343 71.676
R783 B.n508 B.n344 71.676
R784 B.n504 B.n345 71.676
R785 B.n500 B.n346 71.676
R786 B.n496 B.n347 71.676
R787 B.n492 B.n348 71.676
R788 B.n488 B.n349 71.676
R789 B.n484 B.n350 71.676
R790 B.n480 B.n351 71.676
R791 B.n475 B.n352 71.676
R792 B.n471 B.n353 71.676
R793 B.n467 B.n354 71.676
R794 B.n463 B.n355 71.676
R795 B.n459 B.n356 71.676
R796 B.n455 B.n357 71.676
R797 B.n451 B.n358 71.676
R798 B.n447 B.n359 71.676
R799 B.n443 B.n360 71.676
R800 B.n439 B.n361 71.676
R801 B.n435 B.n362 71.676
R802 B.n431 B.n363 71.676
R803 B.n427 B.n364 71.676
R804 B.n423 B.n365 71.676
R805 B.n419 B.n366 71.676
R806 B.n415 B.n367 71.676
R807 B.n411 B.n368 71.676
R808 B.n407 B.n369 71.676
R809 B.n403 B.n370 71.676
R810 B.n399 B.n371 71.676
R811 B.n395 B.n372 71.676
R812 B.n391 B.n373 71.676
R813 B.n387 B.n374 71.676
R814 B.n383 B.n375 71.676
R815 B.n595 B.n594 71.676
R816 B.n686 B.n685 71.676
R817 B.n686 B.n2 71.676
R818 B.n84 B.t15 71.0036
R819 B.n382 B.t11 71.0036
R820 B.n87 B.t5 70.9849
R821 B.n379 B.t8 70.9849
R822 B.n593 B.n321 65.1486
R823 B.n658 B.n657 65.1486
R824 B.n186 B.n87 59.5399
R825 B.n85 B.n84 59.5399
R826 B.n477 B.n382 59.5399
R827 B.n380 B.n379 59.5399
R828 B.n600 B.n321 37.8643
R829 B.n600 B.n316 37.8643
R830 B.n606 B.n316 37.8643
R831 B.n606 B.n317 37.8643
R832 B.n612 B.n309 37.8643
R833 B.n618 B.n309 37.8643
R834 B.n618 B.n305 37.8643
R835 B.n626 B.n305 37.8643
R836 B.n626 B.n625 37.8643
R837 B.n632 B.n4 37.8643
R838 B.n684 B.n4 37.8643
R839 B.n684 B.n683 37.8643
R840 B.n683 B.n682 37.8643
R841 B.n682 B.n8 37.8643
R842 B.n675 B.n12 37.8643
R843 B.n675 B.n674 37.8643
R844 B.n674 B.n673 37.8643
R845 B.n673 B.n16 37.8643
R846 B.n667 B.n16 37.8643
R847 B.n666 B.n665 37.8643
R848 B.n665 B.n23 37.8643
R849 B.n659 B.n23 37.8643
R850 B.n659 B.n658 37.8643
R851 B.n590 B.n319 33.5615
R852 B.n597 B.n596 33.5615
R853 B.n655 B.n654 33.5615
R854 B.n89 B.n25 33.5615
R855 B.n317 B.t7 27.2847
R856 B.t3 B.n666 27.2847
R857 B.n625 B.t1 21.7165
R858 B.n12 B.t0 21.7165
R859 B B.n687 18.0485
R860 B.n87 B.n86 17.455
R861 B.n84 B.n83 17.455
R862 B.n382 B.n381 17.455
R863 B.n379 B.n378 17.455
R864 B.n632 B.t1 16.1483
R865 B.t0 B.n8 16.1483
R866 B.n602 B.n319 10.6151
R867 B.n603 B.n602 10.6151
R868 B.n604 B.n603 10.6151
R869 B.n604 B.n311 10.6151
R870 B.n614 B.n311 10.6151
R871 B.n615 B.n614 10.6151
R872 B.n616 B.n615 10.6151
R873 B.n616 B.n303 10.6151
R874 B.n628 B.n303 10.6151
R875 B.n629 B.n628 10.6151
R876 B.n630 B.n629 10.6151
R877 B.n630 B.n0 10.6151
R878 B.n590 B.n589 10.6151
R879 B.n589 B.n588 10.6151
R880 B.n588 B.n587 10.6151
R881 B.n587 B.n585 10.6151
R882 B.n585 B.n582 10.6151
R883 B.n582 B.n581 10.6151
R884 B.n581 B.n578 10.6151
R885 B.n578 B.n577 10.6151
R886 B.n577 B.n574 10.6151
R887 B.n574 B.n573 10.6151
R888 B.n573 B.n570 10.6151
R889 B.n570 B.n569 10.6151
R890 B.n569 B.n566 10.6151
R891 B.n566 B.n565 10.6151
R892 B.n565 B.n562 10.6151
R893 B.n562 B.n561 10.6151
R894 B.n561 B.n558 10.6151
R895 B.n558 B.n557 10.6151
R896 B.n557 B.n554 10.6151
R897 B.n554 B.n553 10.6151
R898 B.n553 B.n550 10.6151
R899 B.n550 B.n549 10.6151
R900 B.n549 B.n546 10.6151
R901 B.n546 B.n545 10.6151
R902 B.n545 B.n542 10.6151
R903 B.n542 B.n541 10.6151
R904 B.n541 B.n538 10.6151
R905 B.n538 B.n537 10.6151
R906 B.n537 B.n534 10.6151
R907 B.n534 B.n533 10.6151
R908 B.n533 B.n530 10.6151
R909 B.n530 B.n529 10.6151
R910 B.n529 B.n526 10.6151
R911 B.n526 B.n525 10.6151
R912 B.n525 B.n522 10.6151
R913 B.n522 B.n521 10.6151
R914 B.n521 B.n518 10.6151
R915 B.n518 B.n517 10.6151
R916 B.n517 B.n514 10.6151
R917 B.n514 B.n513 10.6151
R918 B.n513 B.n510 10.6151
R919 B.n510 B.n509 10.6151
R920 B.n509 B.n506 10.6151
R921 B.n506 B.n505 10.6151
R922 B.n505 B.n502 10.6151
R923 B.n502 B.n501 10.6151
R924 B.n501 B.n498 10.6151
R925 B.n498 B.n497 10.6151
R926 B.n494 B.n493 10.6151
R927 B.n493 B.n490 10.6151
R928 B.n490 B.n489 10.6151
R929 B.n489 B.n486 10.6151
R930 B.n486 B.n485 10.6151
R931 B.n485 B.n482 10.6151
R932 B.n482 B.n481 10.6151
R933 B.n481 B.n478 10.6151
R934 B.n476 B.n473 10.6151
R935 B.n473 B.n472 10.6151
R936 B.n472 B.n469 10.6151
R937 B.n469 B.n468 10.6151
R938 B.n468 B.n465 10.6151
R939 B.n465 B.n464 10.6151
R940 B.n464 B.n461 10.6151
R941 B.n461 B.n460 10.6151
R942 B.n460 B.n457 10.6151
R943 B.n457 B.n456 10.6151
R944 B.n456 B.n453 10.6151
R945 B.n453 B.n452 10.6151
R946 B.n452 B.n449 10.6151
R947 B.n449 B.n448 10.6151
R948 B.n448 B.n445 10.6151
R949 B.n445 B.n444 10.6151
R950 B.n444 B.n441 10.6151
R951 B.n441 B.n440 10.6151
R952 B.n440 B.n437 10.6151
R953 B.n437 B.n436 10.6151
R954 B.n436 B.n433 10.6151
R955 B.n433 B.n432 10.6151
R956 B.n432 B.n429 10.6151
R957 B.n429 B.n428 10.6151
R958 B.n428 B.n425 10.6151
R959 B.n425 B.n424 10.6151
R960 B.n424 B.n421 10.6151
R961 B.n421 B.n420 10.6151
R962 B.n420 B.n417 10.6151
R963 B.n417 B.n416 10.6151
R964 B.n416 B.n413 10.6151
R965 B.n413 B.n412 10.6151
R966 B.n412 B.n409 10.6151
R967 B.n409 B.n408 10.6151
R968 B.n408 B.n405 10.6151
R969 B.n405 B.n404 10.6151
R970 B.n404 B.n401 10.6151
R971 B.n401 B.n400 10.6151
R972 B.n400 B.n397 10.6151
R973 B.n397 B.n396 10.6151
R974 B.n396 B.n393 10.6151
R975 B.n393 B.n392 10.6151
R976 B.n392 B.n389 10.6151
R977 B.n389 B.n388 10.6151
R978 B.n388 B.n385 10.6151
R979 B.n385 B.n384 10.6151
R980 B.n384 B.n323 10.6151
R981 B.n596 B.n323 10.6151
R982 B.n598 B.n597 10.6151
R983 B.n598 B.n314 10.6151
R984 B.n608 B.n314 10.6151
R985 B.n609 B.n608 10.6151
R986 B.n610 B.n609 10.6151
R987 B.n610 B.n307 10.6151
R988 B.n620 B.n307 10.6151
R989 B.n621 B.n620 10.6151
R990 B.n623 B.n621 10.6151
R991 B.n623 B.n622 10.6151
R992 B.n622 B.n300 10.6151
R993 B.n635 B.n300 10.6151
R994 B.n636 B.n635 10.6151
R995 B.n637 B.n636 10.6151
R996 B.n638 B.n637 10.6151
R997 B.n639 B.n638 10.6151
R998 B.n642 B.n639 10.6151
R999 B.n643 B.n642 10.6151
R1000 B.n644 B.n643 10.6151
R1001 B.n645 B.n644 10.6151
R1002 B.n647 B.n645 10.6151
R1003 B.n648 B.n647 10.6151
R1004 B.n649 B.n648 10.6151
R1005 B.n650 B.n649 10.6151
R1006 B.n652 B.n650 10.6151
R1007 B.n653 B.n652 10.6151
R1008 B.n654 B.n653 10.6151
R1009 B.n679 B.n1 10.6151
R1010 B.n679 B.n678 10.6151
R1011 B.n678 B.n677 10.6151
R1012 B.n677 B.n10 10.6151
R1013 B.n671 B.n10 10.6151
R1014 B.n671 B.n670 10.6151
R1015 B.n670 B.n669 10.6151
R1016 B.n669 B.n18 10.6151
R1017 B.n663 B.n18 10.6151
R1018 B.n663 B.n662 10.6151
R1019 B.n662 B.n661 10.6151
R1020 B.n661 B.n25 10.6151
R1021 B.n90 B.n89 10.6151
R1022 B.n93 B.n90 10.6151
R1023 B.n94 B.n93 10.6151
R1024 B.n97 B.n94 10.6151
R1025 B.n98 B.n97 10.6151
R1026 B.n101 B.n98 10.6151
R1027 B.n102 B.n101 10.6151
R1028 B.n105 B.n102 10.6151
R1029 B.n106 B.n105 10.6151
R1030 B.n109 B.n106 10.6151
R1031 B.n110 B.n109 10.6151
R1032 B.n113 B.n110 10.6151
R1033 B.n114 B.n113 10.6151
R1034 B.n117 B.n114 10.6151
R1035 B.n118 B.n117 10.6151
R1036 B.n121 B.n118 10.6151
R1037 B.n122 B.n121 10.6151
R1038 B.n125 B.n122 10.6151
R1039 B.n126 B.n125 10.6151
R1040 B.n129 B.n126 10.6151
R1041 B.n130 B.n129 10.6151
R1042 B.n133 B.n130 10.6151
R1043 B.n134 B.n133 10.6151
R1044 B.n137 B.n134 10.6151
R1045 B.n138 B.n137 10.6151
R1046 B.n141 B.n138 10.6151
R1047 B.n142 B.n141 10.6151
R1048 B.n145 B.n142 10.6151
R1049 B.n146 B.n145 10.6151
R1050 B.n149 B.n146 10.6151
R1051 B.n150 B.n149 10.6151
R1052 B.n153 B.n150 10.6151
R1053 B.n154 B.n153 10.6151
R1054 B.n157 B.n154 10.6151
R1055 B.n158 B.n157 10.6151
R1056 B.n161 B.n158 10.6151
R1057 B.n162 B.n161 10.6151
R1058 B.n165 B.n162 10.6151
R1059 B.n166 B.n165 10.6151
R1060 B.n169 B.n166 10.6151
R1061 B.n170 B.n169 10.6151
R1062 B.n173 B.n170 10.6151
R1063 B.n174 B.n173 10.6151
R1064 B.n177 B.n174 10.6151
R1065 B.n178 B.n177 10.6151
R1066 B.n181 B.n178 10.6151
R1067 B.n182 B.n181 10.6151
R1068 B.n185 B.n182 10.6151
R1069 B.n190 B.n187 10.6151
R1070 B.n191 B.n190 10.6151
R1071 B.n194 B.n191 10.6151
R1072 B.n195 B.n194 10.6151
R1073 B.n198 B.n195 10.6151
R1074 B.n199 B.n198 10.6151
R1075 B.n202 B.n199 10.6151
R1076 B.n203 B.n202 10.6151
R1077 B.n207 B.n206 10.6151
R1078 B.n210 B.n207 10.6151
R1079 B.n211 B.n210 10.6151
R1080 B.n214 B.n211 10.6151
R1081 B.n215 B.n214 10.6151
R1082 B.n218 B.n215 10.6151
R1083 B.n219 B.n218 10.6151
R1084 B.n222 B.n219 10.6151
R1085 B.n223 B.n222 10.6151
R1086 B.n226 B.n223 10.6151
R1087 B.n227 B.n226 10.6151
R1088 B.n230 B.n227 10.6151
R1089 B.n231 B.n230 10.6151
R1090 B.n234 B.n231 10.6151
R1091 B.n235 B.n234 10.6151
R1092 B.n238 B.n235 10.6151
R1093 B.n239 B.n238 10.6151
R1094 B.n242 B.n239 10.6151
R1095 B.n243 B.n242 10.6151
R1096 B.n246 B.n243 10.6151
R1097 B.n247 B.n246 10.6151
R1098 B.n250 B.n247 10.6151
R1099 B.n251 B.n250 10.6151
R1100 B.n254 B.n251 10.6151
R1101 B.n255 B.n254 10.6151
R1102 B.n258 B.n255 10.6151
R1103 B.n259 B.n258 10.6151
R1104 B.n262 B.n259 10.6151
R1105 B.n263 B.n262 10.6151
R1106 B.n266 B.n263 10.6151
R1107 B.n267 B.n266 10.6151
R1108 B.n270 B.n267 10.6151
R1109 B.n271 B.n270 10.6151
R1110 B.n274 B.n271 10.6151
R1111 B.n275 B.n274 10.6151
R1112 B.n278 B.n275 10.6151
R1113 B.n279 B.n278 10.6151
R1114 B.n282 B.n279 10.6151
R1115 B.n283 B.n282 10.6151
R1116 B.n286 B.n283 10.6151
R1117 B.n287 B.n286 10.6151
R1118 B.n290 B.n287 10.6151
R1119 B.n291 B.n290 10.6151
R1120 B.n294 B.n291 10.6151
R1121 B.n295 B.n294 10.6151
R1122 B.n298 B.n295 10.6151
R1123 B.n299 B.n298 10.6151
R1124 B.n655 B.n299 10.6151
R1125 B.n612 B.t7 10.5801
R1126 B.n667 B.t3 10.5801
R1127 B.n687 B.n0 8.11757
R1128 B.n687 B.n1 8.11757
R1129 B.n494 B.n380 7.18099
R1130 B.n478 B.n477 7.18099
R1131 B.n187 B.n186 7.18099
R1132 B.n203 B.n85 7.18099
R1133 B.n497 B.n380 3.43465
R1134 B.n477 B.n476 3.43465
R1135 B.n186 B.n185 3.43465
R1136 B.n206 B.n85 3.43465
R1137 VP.n0 VP.t1 883.595
R1138 VP.n0 VP.t0 842.442
R1139 VP VP.n0 0.0516364
R1140 VTAIL.n1 VTAIL.t1 49.1472
R1141 VTAIL.n2 VTAIL.t3 49.1471
R1142 VTAIL.n3 VTAIL.t0 49.1471
R1143 VTAIL.n0 VTAIL.t2 49.1471
R1144 VTAIL.n1 VTAIL.n0 26.4014
R1145 VTAIL.n3 VTAIL.n2 25.6255
R1146 VTAIL.n2 VTAIL.n1 0.858259
R1147 VTAIL VTAIL.n0 0.722483
R1148 VTAIL VTAIL.n3 0.136276
R1149 VDD1 VDD1.t1 104.239
R1150 VDD1 VDD1.t0 66.0781
R1151 VN VN.t0 883.975
R1152 VN VN.t1 842.494
R1153 VDD2.n0 VDD2.t0 103.519
R1154 VDD2.n0 VDD2.t1 65.8259
R1155 VDD2 VDD2.n0 0.252655
C0 VDD2 VN 2.1716f
C1 VDD1 VTAIL 6.88745f
C2 VP VTAIL 1.54516f
C3 VDD2 VTAIL 6.9184f
C4 VDD1 VP 2.26759f
C5 VN VTAIL 1.53039f
C6 VDD2 VDD1 0.450707f
C7 VDD2 VP 0.249666f
C8 VDD1 VN 0.148196f
C9 VN VP 4.96057f
C10 VDD2 B 4.151219f
C11 VDD1 B 7.23344f
C12 VTAIL B 7.244626f
C13 VN B 8.745871f
C14 VP B 4.039763f
C15 VDD2.t0 B 3.34169f
C16 VDD2.t1 B 2.81778f
C17 VDD2.n0 B 2.89586f
C18 VN.t1 B 1.23283f
C19 VN.t0 B 1.3429f
C20 VDD1.t0 B 2.82521f
C21 VDD1.t1 B 3.37497f
C22 VTAIL.t2 B 2.19839f
C23 VTAIL.n0 B 1.26553f
C24 VTAIL.t1 B 2.19841f
C25 VTAIL.n1 B 1.27301f
C26 VTAIL.t3 B 2.19839f
C27 VTAIL.n2 B 1.2302f
C28 VTAIL.t0 B 2.19839f
C29 VTAIL.n3 B 1.19034f
C30 VP.t1 B 1.37218f
C31 VP.t0 B 1.262f
C32 VP.n0 B 4.65237f
.ends

