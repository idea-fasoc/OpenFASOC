* NGSPICE file created from diff_pair_sample_0557.ext - technology: sky130A

.subckt diff_pair_sample_0557 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1442_n3546# sky130_fd_pr__pfet_01v8 ad=5.0193 pd=26.52 as=0 ps=0 w=12.87 l=0.85
X1 B.t8 B.t6 B.t7 w_n1442_n3546# sky130_fd_pr__pfet_01v8 ad=5.0193 pd=26.52 as=0 ps=0 w=12.87 l=0.85
X2 B.t5 B.t3 B.t4 w_n1442_n3546# sky130_fd_pr__pfet_01v8 ad=5.0193 pd=26.52 as=0 ps=0 w=12.87 l=0.85
X3 B.t2 B.t0 B.t1 w_n1442_n3546# sky130_fd_pr__pfet_01v8 ad=5.0193 pd=26.52 as=0 ps=0 w=12.87 l=0.85
X4 VDD2.t1 VN.t0 VTAIL.t3 w_n1442_n3546# sky130_fd_pr__pfet_01v8 ad=5.0193 pd=26.52 as=5.0193 ps=26.52 w=12.87 l=0.85
X5 VDD2.t0 VN.t1 VTAIL.t2 w_n1442_n3546# sky130_fd_pr__pfet_01v8 ad=5.0193 pd=26.52 as=5.0193 ps=26.52 w=12.87 l=0.85
X6 VDD1.t1 VP.t0 VTAIL.t1 w_n1442_n3546# sky130_fd_pr__pfet_01v8 ad=5.0193 pd=26.52 as=5.0193 ps=26.52 w=12.87 l=0.85
X7 VDD1.t0 VP.t1 VTAIL.t0 w_n1442_n3546# sky130_fd_pr__pfet_01v8 ad=5.0193 pd=26.52 as=5.0193 ps=26.52 w=12.87 l=0.85
R0 B.n356 B.n63 585
R1 B.n358 B.n357 585
R2 B.n359 B.n62 585
R3 B.n361 B.n360 585
R4 B.n362 B.n61 585
R5 B.n364 B.n363 585
R6 B.n365 B.n60 585
R7 B.n367 B.n366 585
R8 B.n368 B.n59 585
R9 B.n370 B.n369 585
R10 B.n371 B.n58 585
R11 B.n373 B.n372 585
R12 B.n374 B.n57 585
R13 B.n376 B.n375 585
R14 B.n377 B.n56 585
R15 B.n379 B.n378 585
R16 B.n380 B.n55 585
R17 B.n382 B.n381 585
R18 B.n383 B.n54 585
R19 B.n385 B.n384 585
R20 B.n386 B.n53 585
R21 B.n388 B.n387 585
R22 B.n389 B.n52 585
R23 B.n391 B.n390 585
R24 B.n392 B.n51 585
R25 B.n394 B.n393 585
R26 B.n395 B.n50 585
R27 B.n397 B.n396 585
R28 B.n398 B.n49 585
R29 B.n400 B.n399 585
R30 B.n401 B.n48 585
R31 B.n403 B.n402 585
R32 B.n404 B.n47 585
R33 B.n406 B.n405 585
R34 B.n407 B.n46 585
R35 B.n409 B.n408 585
R36 B.n410 B.n45 585
R37 B.n412 B.n411 585
R38 B.n413 B.n44 585
R39 B.n415 B.n414 585
R40 B.n416 B.n43 585
R41 B.n418 B.n417 585
R42 B.n419 B.n39 585
R43 B.n421 B.n420 585
R44 B.n422 B.n38 585
R45 B.n424 B.n423 585
R46 B.n425 B.n37 585
R47 B.n427 B.n426 585
R48 B.n428 B.n36 585
R49 B.n430 B.n429 585
R50 B.n431 B.n35 585
R51 B.n433 B.n432 585
R52 B.n434 B.n34 585
R53 B.n436 B.n435 585
R54 B.n438 B.n31 585
R55 B.n440 B.n439 585
R56 B.n441 B.n30 585
R57 B.n443 B.n442 585
R58 B.n444 B.n29 585
R59 B.n446 B.n445 585
R60 B.n447 B.n28 585
R61 B.n449 B.n448 585
R62 B.n450 B.n27 585
R63 B.n452 B.n451 585
R64 B.n453 B.n26 585
R65 B.n455 B.n454 585
R66 B.n456 B.n25 585
R67 B.n458 B.n457 585
R68 B.n459 B.n24 585
R69 B.n461 B.n460 585
R70 B.n462 B.n23 585
R71 B.n464 B.n463 585
R72 B.n465 B.n22 585
R73 B.n467 B.n466 585
R74 B.n468 B.n21 585
R75 B.n470 B.n469 585
R76 B.n471 B.n20 585
R77 B.n473 B.n472 585
R78 B.n474 B.n19 585
R79 B.n476 B.n475 585
R80 B.n477 B.n18 585
R81 B.n479 B.n478 585
R82 B.n480 B.n17 585
R83 B.n482 B.n481 585
R84 B.n483 B.n16 585
R85 B.n485 B.n484 585
R86 B.n486 B.n15 585
R87 B.n488 B.n487 585
R88 B.n489 B.n14 585
R89 B.n491 B.n490 585
R90 B.n492 B.n13 585
R91 B.n494 B.n493 585
R92 B.n495 B.n12 585
R93 B.n497 B.n496 585
R94 B.n498 B.n11 585
R95 B.n500 B.n499 585
R96 B.n501 B.n10 585
R97 B.n503 B.n502 585
R98 B.n355 B.n354 585
R99 B.n353 B.n64 585
R100 B.n352 B.n351 585
R101 B.n350 B.n65 585
R102 B.n349 B.n348 585
R103 B.n347 B.n66 585
R104 B.n346 B.n345 585
R105 B.n344 B.n67 585
R106 B.n343 B.n342 585
R107 B.n341 B.n68 585
R108 B.n340 B.n339 585
R109 B.n338 B.n69 585
R110 B.n337 B.n336 585
R111 B.n335 B.n70 585
R112 B.n334 B.n333 585
R113 B.n332 B.n71 585
R114 B.n331 B.n330 585
R115 B.n329 B.n72 585
R116 B.n328 B.n327 585
R117 B.n326 B.n73 585
R118 B.n325 B.n324 585
R119 B.n323 B.n74 585
R120 B.n322 B.n321 585
R121 B.n320 B.n75 585
R122 B.n319 B.n318 585
R123 B.n317 B.n76 585
R124 B.n316 B.n315 585
R125 B.n314 B.n77 585
R126 B.n313 B.n312 585
R127 B.n311 B.n78 585
R128 B.n310 B.n309 585
R129 B.n161 B.n132 585
R130 B.n163 B.n162 585
R131 B.n164 B.n131 585
R132 B.n166 B.n165 585
R133 B.n167 B.n130 585
R134 B.n169 B.n168 585
R135 B.n170 B.n129 585
R136 B.n172 B.n171 585
R137 B.n173 B.n128 585
R138 B.n175 B.n174 585
R139 B.n176 B.n127 585
R140 B.n178 B.n177 585
R141 B.n179 B.n126 585
R142 B.n181 B.n180 585
R143 B.n182 B.n125 585
R144 B.n184 B.n183 585
R145 B.n185 B.n124 585
R146 B.n187 B.n186 585
R147 B.n188 B.n123 585
R148 B.n190 B.n189 585
R149 B.n191 B.n122 585
R150 B.n193 B.n192 585
R151 B.n194 B.n121 585
R152 B.n196 B.n195 585
R153 B.n197 B.n120 585
R154 B.n199 B.n198 585
R155 B.n200 B.n119 585
R156 B.n202 B.n201 585
R157 B.n203 B.n118 585
R158 B.n205 B.n204 585
R159 B.n206 B.n117 585
R160 B.n208 B.n207 585
R161 B.n209 B.n116 585
R162 B.n211 B.n210 585
R163 B.n212 B.n115 585
R164 B.n214 B.n213 585
R165 B.n215 B.n114 585
R166 B.n217 B.n216 585
R167 B.n218 B.n113 585
R168 B.n220 B.n219 585
R169 B.n221 B.n112 585
R170 B.n223 B.n222 585
R171 B.n224 B.n111 585
R172 B.n226 B.n225 585
R173 B.n228 B.n108 585
R174 B.n230 B.n229 585
R175 B.n231 B.n107 585
R176 B.n233 B.n232 585
R177 B.n234 B.n106 585
R178 B.n236 B.n235 585
R179 B.n237 B.n105 585
R180 B.n239 B.n238 585
R181 B.n240 B.n104 585
R182 B.n242 B.n241 585
R183 B.n244 B.n243 585
R184 B.n245 B.n100 585
R185 B.n247 B.n246 585
R186 B.n248 B.n99 585
R187 B.n250 B.n249 585
R188 B.n251 B.n98 585
R189 B.n253 B.n252 585
R190 B.n254 B.n97 585
R191 B.n256 B.n255 585
R192 B.n257 B.n96 585
R193 B.n259 B.n258 585
R194 B.n260 B.n95 585
R195 B.n262 B.n261 585
R196 B.n263 B.n94 585
R197 B.n265 B.n264 585
R198 B.n266 B.n93 585
R199 B.n268 B.n267 585
R200 B.n269 B.n92 585
R201 B.n271 B.n270 585
R202 B.n272 B.n91 585
R203 B.n274 B.n273 585
R204 B.n275 B.n90 585
R205 B.n277 B.n276 585
R206 B.n278 B.n89 585
R207 B.n280 B.n279 585
R208 B.n281 B.n88 585
R209 B.n283 B.n282 585
R210 B.n284 B.n87 585
R211 B.n286 B.n285 585
R212 B.n287 B.n86 585
R213 B.n289 B.n288 585
R214 B.n290 B.n85 585
R215 B.n292 B.n291 585
R216 B.n293 B.n84 585
R217 B.n295 B.n294 585
R218 B.n296 B.n83 585
R219 B.n298 B.n297 585
R220 B.n299 B.n82 585
R221 B.n301 B.n300 585
R222 B.n302 B.n81 585
R223 B.n304 B.n303 585
R224 B.n305 B.n80 585
R225 B.n307 B.n306 585
R226 B.n308 B.n79 585
R227 B.n160 B.n159 585
R228 B.n158 B.n133 585
R229 B.n157 B.n156 585
R230 B.n155 B.n134 585
R231 B.n154 B.n153 585
R232 B.n152 B.n135 585
R233 B.n151 B.n150 585
R234 B.n149 B.n136 585
R235 B.n148 B.n147 585
R236 B.n146 B.n137 585
R237 B.n145 B.n144 585
R238 B.n143 B.n138 585
R239 B.n142 B.n141 585
R240 B.n140 B.n139 585
R241 B.n2 B.n0 585
R242 B.n525 B.n1 585
R243 B.n524 B.n523 585
R244 B.n522 B.n3 585
R245 B.n521 B.n520 585
R246 B.n519 B.n4 585
R247 B.n518 B.n517 585
R248 B.n516 B.n5 585
R249 B.n515 B.n514 585
R250 B.n513 B.n6 585
R251 B.n512 B.n511 585
R252 B.n510 B.n7 585
R253 B.n509 B.n508 585
R254 B.n507 B.n8 585
R255 B.n506 B.n505 585
R256 B.n504 B.n9 585
R257 B.n527 B.n526 585
R258 B.n101 B.t0 566.692
R259 B.n109 B.t6 566.692
R260 B.n32 B.t3 566.692
R261 B.n40 B.t9 566.692
R262 B.n159 B.n132 511.721
R263 B.n502 B.n9 511.721
R264 B.n309 B.n308 511.721
R265 B.n356 B.n355 511.721
R266 B.n101 B.t2 414.346
R267 B.n40 B.t10 414.346
R268 B.n109 B.t8 414.346
R269 B.n32 B.t4 414.346
R270 B.n102 B.t1 391.462
R271 B.n41 B.t11 391.462
R272 B.n110 B.t7 391.462
R273 B.n33 B.t5 391.462
R274 B.n159 B.n158 163.367
R275 B.n158 B.n157 163.367
R276 B.n157 B.n134 163.367
R277 B.n153 B.n134 163.367
R278 B.n153 B.n152 163.367
R279 B.n152 B.n151 163.367
R280 B.n151 B.n136 163.367
R281 B.n147 B.n136 163.367
R282 B.n147 B.n146 163.367
R283 B.n146 B.n145 163.367
R284 B.n145 B.n138 163.367
R285 B.n141 B.n138 163.367
R286 B.n141 B.n140 163.367
R287 B.n140 B.n2 163.367
R288 B.n526 B.n2 163.367
R289 B.n526 B.n525 163.367
R290 B.n525 B.n524 163.367
R291 B.n524 B.n3 163.367
R292 B.n520 B.n3 163.367
R293 B.n520 B.n519 163.367
R294 B.n519 B.n518 163.367
R295 B.n518 B.n5 163.367
R296 B.n514 B.n5 163.367
R297 B.n514 B.n513 163.367
R298 B.n513 B.n512 163.367
R299 B.n512 B.n7 163.367
R300 B.n508 B.n7 163.367
R301 B.n508 B.n507 163.367
R302 B.n507 B.n506 163.367
R303 B.n506 B.n9 163.367
R304 B.n163 B.n132 163.367
R305 B.n164 B.n163 163.367
R306 B.n165 B.n164 163.367
R307 B.n165 B.n130 163.367
R308 B.n169 B.n130 163.367
R309 B.n170 B.n169 163.367
R310 B.n171 B.n170 163.367
R311 B.n171 B.n128 163.367
R312 B.n175 B.n128 163.367
R313 B.n176 B.n175 163.367
R314 B.n177 B.n176 163.367
R315 B.n177 B.n126 163.367
R316 B.n181 B.n126 163.367
R317 B.n182 B.n181 163.367
R318 B.n183 B.n182 163.367
R319 B.n183 B.n124 163.367
R320 B.n187 B.n124 163.367
R321 B.n188 B.n187 163.367
R322 B.n189 B.n188 163.367
R323 B.n189 B.n122 163.367
R324 B.n193 B.n122 163.367
R325 B.n194 B.n193 163.367
R326 B.n195 B.n194 163.367
R327 B.n195 B.n120 163.367
R328 B.n199 B.n120 163.367
R329 B.n200 B.n199 163.367
R330 B.n201 B.n200 163.367
R331 B.n201 B.n118 163.367
R332 B.n205 B.n118 163.367
R333 B.n206 B.n205 163.367
R334 B.n207 B.n206 163.367
R335 B.n207 B.n116 163.367
R336 B.n211 B.n116 163.367
R337 B.n212 B.n211 163.367
R338 B.n213 B.n212 163.367
R339 B.n213 B.n114 163.367
R340 B.n217 B.n114 163.367
R341 B.n218 B.n217 163.367
R342 B.n219 B.n218 163.367
R343 B.n219 B.n112 163.367
R344 B.n223 B.n112 163.367
R345 B.n224 B.n223 163.367
R346 B.n225 B.n224 163.367
R347 B.n225 B.n108 163.367
R348 B.n230 B.n108 163.367
R349 B.n231 B.n230 163.367
R350 B.n232 B.n231 163.367
R351 B.n232 B.n106 163.367
R352 B.n236 B.n106 163.367
R353 B.n237 B.n236 163.367
R354 B.n238 B.n237 163.367
R355 B.n238 B.n104 163.367
R356 B.n242 B.n104 163.367
R357 B.n243 B.n242 163.367
R358 B.n243 B.n100 163.367
R359 B.n247 B.n100 163.367
R360 B.n248 B.n247 163.367
R361 B.n249 B.n248 163.367
R362 B.n249 B.n98 163.367
R363 B.n253 B.n98 163.367
R364 B.n254 B.n253 163.367
R365 B.n255 B.n254 163.367
R366 B.n255 B.n96 163.367
R367 B.n259 B.n96 163.367
R368 B.n260 B.n259 163.367
R369 B.n261 B.n260 163.367
R370 B.n261 B.n94 163.367
R371 B.n265 B.n94 163.367
R372 B.n266 B.n265 163.367
R373 B.n267 B.n266 163.367
R374 B.n267 B.n92 163.367
R375 B.n271 B.n92 163.367
R376 B.n272 B.n271 163.367
R377 B.n273 B.n272 163.367
R378 B.n273 B.n90 163.367
R379 B.n277 B.n90 163.367
R380 B.n278 B.n277 163.367
R381 B.n279 B.n278 163.367
R382 B.n279 B.n88 163.367
R383 B.n283 B.n88 163.367
R384 B.n284 B.n283 163.367
R385 B.n285 B.n284 163.367
R386 B.n285 B.n86 163.367
R387 B.n289 B.n86 163.367
R388 B.n290 B.n289 163.367
R389 B.n291 B.n290 163.367
R390 B.n291 B.n84 163.367
R391 B.n295 B.n84 163.367
R392 B.n296 B.n295 163.367
R393 B.n297 B.n296 163.367
R394 B.n297 B.n82 163.367
R395 B.n301 B.n82 163.367
R396 B.n302 B.n301 163.367
R397 B.n303 B.n302 163.367
R398 B.n303 B.n80 163.367
R399 B.n307 B.n80 163.367
R400 B.n308 B.n307 163.367
R401 B.n309 B.n78 163.367
R402 B.n313 B.n78 163.367
R403 B.n314 B.n313 163.367
R404 B.n315 B.n314 163.367
R405 B.n315 B.n76 163.367
R406 B.n319 B.n76 163.367
R407 B.n320 B.n319 163.367
R408 B.n321 B.n320 163.367
R409 B.n321 B.n74 163.367
R410 B.n325 B.n74 163.367
R411 B.n326 B.n325 163.367
R412 B.n327 B.n326 163.367
R413 B.n327 B.n72 163.367
R414 B.n331 B.n72 163.367
R415 B.n332 B.n331 163.367
R416 B.n333 B.n332 163.367
R417 B.n333 B.n70 163.367
R418 B.n337 B.n70 163.367
R419 B.n338 B.n337 163.367
R420 B.n339 B.n338 163.367
R421 B.n339 B.n68 163.367
R422 B.n343 B.n68 163.367
R423 B.n344 B.n343 163.367
R424 B.n345 B.n344 163.367
R425 B.n345 B.n66 163.367
R426 B.n349 B.n66 163.367
R427 B.n350 B.n349 163.367
R428 B.n351 B.n350 163.367
R429 B.n351 B.n64 163.367
R430 B.n355 B.n64 163.367
R431 B.n502 B.n501 163.367
R432 B.n501 B.n500 163.367
R433 B.n500 B.n11 163.367
R434 B.n496 B.n11 163.367
R435 B.n496 B.n495 163.367
R436 B.n495 B.n494 163.367
R437 B.n494 B.n13 163.367
R438 B.n490 B.n13 163.367
R439 B.n490 B.n489 163.367
R440 B.n489 B.n488 163.367
R441 B.n488 B.n15 163.367
R442 B.n484 B.n15 163.367
R443 B.n484 B.n483 163.367
R444 B.n483 B.n482 163.367
R445 B.n482 B.n17 163.367
R446 B.n478 B.n17 163.367
R447 B.n478 B.n477 163.367
R448 B.n477 B.n476 163.367
R449 B.n476 B.n19 163.367
R450 B.n472 B.n19 163.367
R451 B.n472 B.n471 163.367
R452 B.n471 B.n470 163.367
R453 B.n470 B.n21 163.367
R454 B.n466 B.n21 163.367
R455 B.n466 B.n465 163.367
R456 B.n465 B.n464 163.367
R457 B.n464 B.n23 163.367
R458 B.n460 B.n23 163.367
R459 B.n460 B.n459 163.367
R460 B.n459 B.n458 163.367
R461 B.n458 B.n25 163.367
R462 B.n454 B.n25 163.367
R463 B.n454 B.n453 163.367
R464 B.n453 B.n452 163.367
R465 B.n452 B.n27 163.367
R466 B.n448 B.n27 163.367
R467 B.n448 B.n447 163.367
R468 B.n447 B.n446 163.367
R469 B.n446 B.n29 163.367
R470 B.n442 B.n29 163.367
R471 B.n442 B.n441 163.367
R472 B.n441 B.n440 163.367
R473 B.n440 B.n31 163.367
R474 B.n435 B.n31 163.367
R475 B.n435 B.n434 163.367
R476 B.n434 B.n433 163.367
R477 B.n433 B.n35 163.367
R478 B.n429 B.n35 163.367
R479 B.n429 B.n428 163.367
R480 B.n428 B.n427 163.367
R481 B.n427 B.n37 163.367
R482 B.n423 B.n37 163.367
R483 B.n423 B.n422 163.367
R484 B.n422 B.n421 163.367
R485 B.n421 B.n39 163.367
R486 B.n417 B.n39 163.367
R487 B.n417 B.n416 163.367
R488 B.n416 B.n415 163.367
R489 B.n415 B.n44 163.367
R490 B.n411 B.n44 163.367
R491 B.n411 B.n410 163.367
R492 B.n410 B.n409 163.367
R493 B.n409 B.n46 163.367
R494 B.n405 B.n46 163.367
R495 B.n405 B.n404 163.367
R496 B.n404 B.n403 163.367
R497 B.n403 B.n48 163.367
R498 B.n399 B.n48 163.367
R499 B.n399 B.n398 163.367
R500 B.n398 B.n397 163.367
R501 B.n397 B.n50 163.367
R502 B.n393 B.n50 163.367
R503 B.n393 B.n392 163.367
R504 B.n392 B.n391 163.367
R505 B.n391 B.n52 163.367
R506 B.n387 B.n52 163.367
R507 B.n387 B.n386 163.367
R508 B.n386 B.n385 163.367
R509 B.n385 B.n54 163.367
R510 B.n381 B.n54 163.367
R511 B.n381 B.n380 163.367
R512 B.n380 B.n379 163.367
R513 B.n379 B.n56 163.367
R514 B.n375 B.n56 163.367
R515 B.n375 B.n374 163.367
R516 B.n374 B.n373 163.367
R517 B.n373 B.n58 163.367
R518 B.n369 B.n58 163.367
R519 B.n369 B.n368 163.367
R520 B.n368 B.n367 163.367
R521 B.n367 B.n60 163.367
R522 B.n363 B.n60 163.367
R523 B.n363 B.n362 163.367
R524 B.n362 B.n361 163.367
R525 B.n361 B.n62 163.367
R526 B.n357 B.n62 163.367
R527 B.n357 B.n356 163.367
R528 B.n103 B.n102 59.5399
R529 B.n227 B.n110 59.5399
R530 B.n437 B.n33 59.5399
R531 B.n42 B.n41 59.5399
R532 B.n504 B.n503 33.2493
R533 B.n354 B.n63 33.2493
R534 B.n310 B.n79 33.2493
R535 B.n161 B.n160 33.2493
R536 B.n102 B.n101 22.8853
R537 B.n110 B.n109 22.8853
R538 B.n33 B.n32 22.8853
R539 B.n41 B.n40 22.8853
R540 B B.n527 18.0485
R541 B.n503 B.n10 10.6151
R542 B.n499 B.n10 10.6151
R543 B.n499 B.n498 10.6151
R544 B.n498 B.n497 10.6151
R545 B.n497 B.n12 10.6151
R546 B.n493 B.n12 10.6151
R547 B.n493 B.n492 10.6151
R548 B.n492 B.n491 10.6151
R549 B.n491 B.n14 10.6151
R550 B.n487 B.n14 10.6151
R551 B.n487 B.n486 10.6151
R552 B.n486 B.n485 10.6151
R553 B.n485 B.n16 10.6151
R554 B.n481 B.n16 10.6151
R555 B.n481 B.n480 10.6151
R556 B.n480 B.n479 10.6151
R557 B.n479 B.n18 10.6151
R558 B.n475 B.n18 10.6151
R559 B.n475 B.n474 10.6151
R560 B.n474 B.n473 10.6151
R561 B.n473 B.n20 10.6151
R562 B.n469 B.n20 10.6151
R563 B.n469 B.n468 10.6151
R564 B.n468 B.n467 10.6151
R565 B.n467 B.n22 10.6151
R566 B.n463 B.n22 10.6151
R567 B.n463 B.n462 10.6151
R568 B.n462 B.n461 10.6151
R569 B.n461 B.n24 10.6151
R570 B.n457 B.n24 10.6151
R571 B.n457 B.n456 10.6151
R572 B.n456 B.n455 10.6151
R573 B.n455 B.n26 10.6151
R574 B.n451 B.n26 10.6151
R575 B.n451 B.n450 10.6151
R576 B.n450 B.n449 10.6151
R577 B.n449 B.n28 10.6151
R578 B.n445 B.n28 10.6151
R579 B.n445 B.n444 10.6151
R580 B.n444 B.n443 10.6151
R581 B.n443 B.n30 10.6151
R582 B.n439 B.n30 10.6151
R583 B.n439 B.n438 10.6151
R584 B.n436 B.n34 10.6151
R585 B.n432 B.n34 10.6151
R586 B.n432 B.n431 10.6151
R587 B.n431 B.n430 10.6151
R588 B.n430 B.n36 10.6151
R589 B.n426 B.n36 10.6151
R590 B.n426 B.n425 10.6151
R591 B.n425 B.n424 10.6151
R592 B.n424 B.n38 10.6151
R593 B.n420 B.n419 10.6151
R594 B.n419 B.n418 10.6151
R595 B.n418 B.n43 10.6151
R596 B.n414 B.n43 10.6151
R597 B.n414 B.n413 10.6151
R598 B.n413 B.n412 10.6151
R599 B.n412 B.n45 10.6151
R600 B.n408 B.n45 10.6151
R601 B.n408 B.n407 10.6151
R602 B.n407 B.n406 10.6151
R603 B.n406 B.n47 10.6151
R604 B.n402 B.n47 10.6151
R605 B.n402 B.n401 10.6151
R606 B.n401 B.n400 10.6151
R607 B.n400 B.n49 10.6151
R608 B.n396 B.n49 10.6151
R609 B.n396 B.n395 10.6151
R610 B.n395 B.n394 10.6151
R611 B.n394 B.n51 10.6151
R612 B.n390 B.n51 10.6151
R613 B.n390 B.n389 10.6151
R614 B.n389 B.n388 10.6151
R615 B.n388 B.n53 10.6151
R616 B.n384 B.n53 10.6151
R617 B.n384 B.n383 10.6151
R618 B.n383 B.n382 10.6151
R619 B.n382 B.n55 10.6151
R620 B.n378 B.n55 10.6151
R621 B.n378 B.n377 10.6151
R622 B.n377 B.n376 10.6151
R623 B.n376 B.n57 10.6151
R624 B.n372 B.n57 10.6151
R625 B.n372 B.n371 10.6151
R626 B.n371 B.n370 10.6151
R627 B.n370 B.n59 10.6151
R628 B.n366 B.n59 10.6151
R629 B.n366 B.n365 10.6151
R630 B.n365 B.n364 10.6151
R631 B.n364 B.n61 10.6151
R632 B.n360 B.n61 10.6151
R633 B.n360 B.n359 10.6151
R634 B.n359 B.n358 10.6151
R635 B.n358 B.n63 10.6151
R636 B.n311 B.n310 10.6151
R637 B.n312 B.n311 10.6151
R638 B.n312 B.n77 10.6151
R639 B.n316 B.n77 10.6151
R640 B.n317 B.n316 10.6151
R641 B.n318 B.n317 10.6151
R642 B.n318 B.n75 10.6151
R643 B.n322 B.n75 10.6151
R644 B.n323 B.n322 10.6151
R645 B.n324 B.n323 10.6151
R646 B.n324 B.n73 10.6151
R647 B.n328 B.n73 10.6151
R648 B.n329 B.n328 10.6151
R649 B.n330 B.n329 10.6151
R650 B.n330 B.n71 10.6151
R651 B.n334 B.n71 10.6151
R652 B.n335 B.n334 10.6151
R653 B.n336 B.n335 10.6151
R654 B.n336 B.n69 10.6151
R655 B.n340 B.n69 10.6151
R656 B.n341 B.n340 10.6151
R657 B.n342 B.n341 10.6151
R658 B.n342 B.n67 10.6151
R659 B.n346 B.n67 10.6151
R660 B.n347 B.n346 10.6151
R661 B.n348 B.n347 10.6151
R662 B.n348 B.n65 10.6151
R663 B.n352 B.n65 10.6151
R664 B.n353 B.n352 10.6151
R665 B.n354 B.n353 10.6151
R666 B.n162 B.n161 10.6151
R667 B.n162 B.n131 10.6151
R668 B.n166 B.n131 10.6151
R669 B.n167 B.n166 10.6151
R670 B.n168 B.n167 10.6151
R671 B.n168 B.n129 10.6151
R672 B.n172 B.n129 10.6151
R673 B.n173 B.n172 10.6151
R674 B.n174 B.n173 10.6151
R675 B.n174 B.n127 10.6151
R676 B.n178 B.n127 10.6151
R677 B.n179 B.n178 10.6151
R678 B.n180 B.n179 10.6151
R679 B.n180 B.n125 10.6151
R680 B.n184 B.n125 10.6151
R681 B.n185 B.n184 10.6151
R682 B.n186 B.n185 10.6151
R683 B.n186 B.n123 10.6151
R684 B.n190 B.n123 10.6151
R685 B.n191 B.n190 10.6151
R686 B.n192 B.n191 10.6151
R687 B.n192 B.n121 10.6151
R688 B.n196 B.n121 10.6151
R689 B.n197 B.n196 10.6151
R690 B.n198 B.n197 10.6151
R691 B.n198 B.n119 10.6151
R692 B.n202 B.n119 10.6151
R693 B.n203 B.n202 10.6151
R694 B.n204 B.n203 10.6151
R695 B.n204 B.n117 10.6151
R696 B.n208 B.n117 10.6151
R697 B.n209 B.n208 10.6151
R698 B.n210 B.n209 10.6151
R699 B.n210 B.n115 10.6151
R700 B.n214 B.n115 10.6151
R701 B.n215 B.n214 10.6151
R702 B.n216 B.n215 10.6151
R703 B.n216 B.n113 10.6151
R704 B.n220 B.n113 10.6151
R705 B.n221 B.n220 10.6151
R706 B.n222 B.n221 10.6151
R707 B.n222 B.n111 10.6151
R708 B.n226 B.n111 10.6151
R709 B.n229 B.n228 10.6151
R710 B.n229 B.n107 10.6151
R711 B.n233 B.n107 10.6151
R712 B.n234 B.n233 10.6151
R713 B.n235 B.n234 10.6151
R714 B.n235 B.n105 10.6151
R715 B.n239 B.n105 10.6151
R716 B.n240 B.n239 10.6151
R717 B.n241 B.n240 10.6151
R718 B.n245 B.n244 10.6151
R719 B.n246 B.n245 10.6151
R720 B.n246 B.n99 10.6151
R721 B.n250 B.n99 10.6151
R722 B.n251 B.n250 10.6151
R723 B.n252 B.n251 10.6151
R724 B.n252 B.n97 10.6151
R725 B.n256 B.n97 10.6151
R726 B.n257 B.n256 10.6151
R727 B.n258 B.n257 10.6151
R728 B.n258 B.n95 10.6151
R729 B.n262 B.n95 10.6151
R730 B.n263 B.n262 10.6151
R731 B.n264 B.n263 10.6151
R732 B.n264 B.n93 10.6151
R733 B.n268 B.n93 10.6151
R734 B.n269 B.n268 10.6151
R735 B.n270 B.n269 10.6151
R736 B.n270 B.n91 10.6151
R737 B.n274 B.n91 10.6151
R738 B.n275 B.n274 10.6151
R739 B.n276 B.n275 10.6151
R740 B.n276 B.n89 10.6151
R741 B.n280 B.n89 10.6151
R742 B.n281 B.n280 10.6151
R743 B.n282 B.n281 10.6151
R744 B.n282 B.n87 10.6151
R745 B.n286 B.n87 10.6151
R746 B.n287 B.n286 10.6151
R747 B.n288 B.n287 10.6151
R748 B.n288 B.n85 10.6151
R749 B.n292 B.n85 10.6151
R750 B.n293 B.n292 10.6151
R751 B.n294 B.n293 10.6151
R752 B.n294 B.n83 10.6151
R753 B.n298 B.n83 10.6151
R754 B.n299 B.n298 10.6151
R755 B.n300 B.n299 10.6151
R756 B.n300 B.n81 10.6151
R757 B.n304 B.n81 10.6151
R758 B.n305 B.n304 10.6151
R759 B.n306 B.n305 10.6151
R760 B.n306 B.n79 10.6151
R761 B.n160 B.n133 10.6151
R762 B.n156 B.n133 10.6151
R763 B.n156 B.n155 10.6151
R764 B.n155 B.n154 10.6151
R765 B.n154 B.n135 10.6151
R766 B.n150 B.n135 10.6151
R767 B.n150 B.n149 10.6151
R768 B.n149 B.n148 10.6151
R769 B.n148 B.n137 10.6151
R770 B.n144 B.n137 10.6151
R771 B.n144 B.n143 10.6151
R772 B.n143 B.n142 10.6151
R773 B.n142 B.n139 10.6151
R774 B.n139 B.n0 10.6151
R775 B.n523 B.n1 10.6151
R776 B.n523 B.n522 10.6151
R777 B.n522 B.n521 10.6151
R778 B.n521 B.n4 10.6151
R779 B.n517 B.n4 10.6151
R780 B.n517 B.n516 10.6151
R781 B.n516 B.n515 10.6151
R782 B.n515 B.n6 10.6151
R783 B.n511 B.n6 10.6151
R784 B.n511 B.n510 10.6151
R785 B.n510 B.n509 10.6151
R786 B.n509 B.n8 10.6151
R787 B.n505 B.n8 10.6151
R788 B.n505 B.n504 10.6151
R789 B.n438 B.n437 8.74196
R790 B.n420 B.n42 8.74196
R791 B.n227 B.n226 8.74196
R792 B.n244 B.n103 8.74196
R793 B.n527 B.n0 2.81026
R794 B.n527 B.n1 2.81026
R795 B.n437 B.n436 1.87367
R796 B.n42 B.n38 1.87367
R797 B.n228 B.n227 1.87367
R798 B.n241 B.n103 1.87367
R799 VN VN.t1 613.771
R800 VN VN.t0 572.753
R801 VTAIL.n274 VTAIL.n210 756.745
R802 VTAIL.n64 VTAIL.n0 756.745
R803 VTAIL.n204 VTAIL.n140 756.745
R804 VTAIL.n134 VTAIL.n70 756.745
R805 VTAIL.n233 VTAIL.n232 585
R806 VTAIL.n230 VTAIL.n229 585
R807 VTAIL.n239 VTAIL.n238 585
R808 VTAIL.n241 VTAIL.n240 585
R809 VTAIL.n226 VTAIL.n225 585
R810 VTAIL.n247 VTAIL.n246 585
R811 VTAIL.n250 VTAIL.n249 585
R812 VTAIL.n248 VTAIL.n222 585
R813 VTAIL.n255 VTAIL.n221 585
R814 VTAIL.n257 VTAIL.n256 585
R815 VTAIL.n259 VTAIL.n258 585
R816 VTAIL.n218 VTAIL.n217 585
R817 VTAIL.n265 VTAIL.n264 585
R818 VTAIL.n267 VTAIL.n266 585
R819 VTAIL.n214 VTAIL.n213 585
R820 VTAIL.n273 VTAIL.n272 585
R821 VTAIL.n275 VTAIL.n274 585
R822 VTAIL.n23 VTAIL.n22 585
R823 VTAIL.n20 VTAIL.n19 585
R824 VTAIL.n29 VTAIL.n28 585
R825 VTAIL.n31 VTAIL.n30 585
R826 VTAIL.n16 VTAIL.n15 585
R827 VTAIL.n37 VTAIL.n36 585
R828 VTAIL.n40 VTAIL.n39 585
R829 VTAIL.n38 VTAIL.n12 585
R830 VTAIL.n45 VTAIL.n11 585
R831 VTAIL.n47 VTAIL.n46 585
R832 VTAIL.n49 VTAIL.n48 585
R833 VTAIL.n8 VTAIL.n7 585
R834 VTAIL.n55 VTAIL.n54 585
R835 VTAIL.n57 VTAIL.n56 585
R836 VTAIL.n4 VTAIL.n3 585
R837 VTAIL.n63 VTAIL.n62 585
R838 VTAIL.n65 VTAIL.n64 585
R839 VTAIL.n205 VTAIL.n204 585
R840 VTAIL.n203 VTAIL.n202 585
R841 VTAIL.n144 VTAIL.n143 585
R842 VTAIL.n197 VTAIL.n196 585
R843 VTAIL.n195 VTAIL.n194 585
R844 VTAIL.n148 VTAIL.n147 585
R845 VTAIL.n189 VTAIL.n188 585
R846 VTAIL.n187 VTAIL.n186 585
R847 VTAIL.n185 VTAIL.n151 585
R848 VTAIL.n155 VTAIL.n152 585
R849 VTAIL.n180 VTAIL.n179 585
R850 VTAIL.n178 VTAIL.n177 585
R851 VTAIL.n157 VTAIL.n156 585
R852 VTAIL.n172 VTAIL.n171 585
R853 VTAIL.n170 VTAIL.n169 585
R854 VTAIL.n161 VTAIL.n160 585
R855 VTAIL.n164 VTAIL.n163 585
R856 VTAIL.n135 VTAIL.n134 585
R857 VTAIL.n133 VTAIL.n132 585
R858 VTAIL.n74 VTAIL.n73 585
R859 VTAIL.n127 VTAIL.n126 585
R860 VTAIL.n125 VTAIL.n124 585
R861 VTAIL.n78 VTAIL.n77 585
R862 VTAIL.n119 VTAIL.n118 585
R863 VTAIL.n117 VTAIL.n116 585
R864 VTAIL.n115 VTAIL.n81 585
R865 VTAIL.n85 VTAIL.n82 585
R866 VTAIL.n110 VTAIL.n109 585
R867 VTAIL.n108 VTAIL.n107 585
R868 VTAIL.n87 VTAIL.n86 585
R869 VTAIL.n102 VTAIL.n101 585
R870 VTAIL.n100 VTAIL.n99 585
R871 VTAIL.n91 VTAIL.n90 585
R872 VTAIL.n94 VTAIL.n93 585
R873 VTAIL.t3 VTAIL.n231 329.036
R874 VTAIL.t0 VTAIL.n21 329.036
R875 VTAIL.t1 VTAIL.n162 329.036
R876 VTAIL.t2 VTAIL.n92 329.036
R877 VTAIL.n232 VTAIL.n229 171.744
R878 VTAIL.n239 VTAIL.n229 171.744
R879 VTAIL.n240 VTAIL.n239 171.744
R880 VTAIL.n240 VTAIL.n225 171.744
R881 VTAIL.n247 VTAIL.n225 171.744
R882 VTAIL.n249 VTAIL.n247 171.744
R883 VTAIL.n249 VTAIL.n248 171.744
R884 VTAIL.n248 VTAIL.n221 171.744
R885 VTAIL.n257 VTAIL.n221 171.744
R886 VTAIL.n258 VTAIL.n257 171.744
R887 VTAIL.n258 VTAIL.n217 171.744
R888 VTAIL.n265 VTAIL.n217 171.744
R889 VTAIL.n266 VTAIL.n265 171.744
R890 VTAIL.n266 VTAIL.n213 171.744
R891 VTAIL.n273 VTAIL.n213 171.744
R892 VTAIL.n274 VTAIL.n273 171.744
R893 VTAIL.n22 VTAIL.n19 171.744
R894 VTAIL.n29 VTAIL.n19 171.744
R895 VTAIL.n30 VTAIL.n29 171.744
R896 VTAIL.n30 VTAIL.n15 171.744
R897 VTAIL.n37 VTAIL.n15 171.744
R898 VTAIL.n39 VTAIL.n37 171.744
R899 VTAIL.n39 VTAIL.n38 171.744
R900 VTAIL.n38 VTAIL.n11 171.744
R901 VTAIL.n47 VTAIL.n11 171.744
R902 VTAIL.n48 VTAIL.n47 171.744
R903 VTAIL.n48 VTAIL.n7 171.744
R904 VTAIL.n55 VTAIL.n7 171.744
R905 VTAIL.n56 VTAIL.n55 171.744
R906 VTAIL.n56 VTAIL.n3 171.744
R907 VTAIL.n63 VTAIL.n3 171.744
R908 VTAIL.n64 VTAIL.n63 171.744
R909 VTAIL.n204 VTAIL.n203 171.744
R910 VTAIL.n203 VTAIL.n143 171.744
R911 VTAIL.n196 VTAIL.n143 171.744
R912 VTAIL.n196 VTAIL.n195 171.744
R913 VTAIL.n195 VTAIL.n147 171.744
R914 VTAIL.n188 VTAIL.n147 171.744
R915 VTAIL.n188 VTAIL.n187 171.744
R916 VTAIL.n187 VTAIL.n151 171.744
R917 VTAIL.n155 VTAIL.n151 171.744
R918 VTAIL.n179 VTAIL.n155 171.744
R919 VTAIL.n179 VTAIL.n178 171.744
R920 VTAIL.n178 VTAIL.n156 171.744
R921 VTAIL.n171 VTAIL.n156 171.744
R922 VTAIL.n171 VTAIL.n170 171.744
R923 VTAIL.n170 VTAIL.n160 171.744
R924 VTAIL.n163 VTAIL.n160 171.744
R925 VTAIL.n134 VTAIL.n133 171.744
R926 VTAIL.n133 VTAIL.n73 171.744
R927 VTAIL.n126 VTAIL.n73 171.744
R928 VTAIL.n126 VTAIL.n125 171.744
R929 VTAIL.n125 VTAIL.n77 171.744
R930 VTAIL.n118 VTAIL.n77 171.744
R931 VTAIL.n118 VTAIL.n117 171.744
R932 VTAIL.n117 VTAIL.n81 171.744
R933 VTAIL.n85 VTAIL.n81 171.744
R934 VTAIL.n109 VTAIL.n85 171.744
R935 VTAIL.n109 VTAIL.n108 171.744
R936 VTAIL.n108 VTAIL.n86 171.744
R937 VTAIL.n101 VTAIL.n86 171.744
R938 VTAIL.n101 VTAIL.n100 171.744
R939 VTAIL.n100 VTAIL.n90 171.744
R940 VTAIL.n93 VTAIL.n90 171.744
R941 VTAIL.n232 VTAIL.t3 85.8723
R942 VTAIL.n22 VTAIL.t0 85.8723
R943 VTAIL.n163 VTAIL.t1 85.8723
R944 VTAIL.n93 VTAIL.t2 85.8723
R945 VTAIL.n279 VTAIL.n278 32.7672
R946 VTAIL.n69 VTAIL.n68 32.7672
R947 VTAIL.n209 VTAIL.n208 32.7672
R948 VTAIL.n139 VTAIL.n138 32.7672
R949 VTAIL.n139 VTAIL.n69 25.5134
R950 VTAIL.n279 VTAIL.n209 24.4962
R951 VTAIL.n256 VTAIL.n255 13.1884
R952 VTAIL.n46 VTAIL.n45 13.1884
R953 VTAIL.n186 VTAIL.n185 13.1884
R954 VTAIL.n116 VTAIL.n115 13.1884
R955 VTAIL.n254 VTAIL.n222 12.8005
R956 VTAIL.n259 VTAIL.n220 12.8005
R957 VTAIL.n44 VTAIL.n12 12.8005
R958 VTAIL.n49 VTAIL.n10 12.8005
R959 VTAIL.n189 VTAIL.n150 12.8005
R960 VTAIL.n184 VTAIL.n152 12.8005
R961 VTAIL.n119 VTAIL.n80 12.8005
R962 VTAIL.n114 VTAIL.n82 12.8005
R963 VTAIL.n251 VTAIL.n250 12.0247
R964 VTAIL.n260 VTAIL.n218 12.0247
R965 VTAIL.n41 VTAIL.n40 12.0247
R966 VTAIL.n50 VTAIL.n8 12.0247
R967 VTAIL.n190 VTAIL.n148 12.0247
R968 VTAIL.n181 VTAIL.n180 12.0247
R969 VTAIL.n120 VTAIL.n78 12.0247
R970 VTAIL.n111 VTAIL.n110 12.0247
R971 VTAIL.n246 VTAIL.n224 11.249
R972 VTAIL.n264 VTAIL.n263 11.249
R973 VTAIL.n36 VTAIL.n14 11.249
R974 VTAIL.n54 VTAIL.n53 11.249
R975 VTAIL.n194 VTAIL.n193 11.249
R976 VTAIL.n177 VTAIL.n154 11.249
R977 VTAIL.n124 VTAIL.n123 11.249
R978 VTAIL.n107 VTAIL.n84 11.249
R979 VTAIL.n233 VTAIL.n231 10.7239
R980 VTAIL.n23 VTAIL.n21 10.7239
R981 VTAIL.n164 VTAIL.n162 10.7239
R982 VTAIL.n94 VTAIL.n92 10.7239
R983 VTAIL.n245 VTAIL.n226 10.4732
R984 VTAIL.n267 VTAIL.n216 10.4732
R985 VTAIL.n35 VTAIL.n16 10.4732
R986 VTAIL.n57 VTAIL.n6 10.4732
R987 VTAIL.n197 VTAIL.n146 10.4732
R988 VTAIL.n176 VTAIL.n157 10.4732
R989 VTAIL.n127 VTAIL.n76 10.4732
R990 VTAIL.n106 VTAIL.n87 10.4732
R991 VTAIL.n242 VTAIL.n241 9.69747
R992 VTAIL.n268 VTAIL.n214 9.69747
R993 VTAIL.n32 VTAIL.n31 9.69747
R994 VTAIL.n58 VTAIL.n4 9.69747
R995 VTAIL.n198 VTAIL.n144 9.69747
R996 VTAIL.n173 VTAIL.n172 9.69747
R997 VTAIL.n128 VTAIL.n74 9.69747
R998 VTAIL.n103 VTAIL.n102 9.69747
R999 VTAIL.n278 VTAIL.n277 9.45567
R1000 VTAIL.n68 VTAIL.n67 9.45567
R1001 VTAIL.n208 VTAIL.n207 9.45567
R1002 VTAIL.n138 VTAIL.n137 9.45567
R1003 VTAIL.n212 VTAIL.n211 9.3005
R1004 VTAIL.n271 VTAIL.n270 9.3005
R1005 VTAIL.n269 VTAIL.n268 9.3005
R1006 VTAIL.n216 VTAIL.n215 9.3005
R1007 VTAIL.n263 VTAIL.n262 9.3005
R1008 VTAIL.n261 VTAIL.n260 9.3005
R1009 VTAIL.n220 VTAIL.n219 9.3005
R1010 VTAIL.n235 VTAIL.n234 9.3005
R1011 VTAIL.n237 VTAIL.n236 9.3005
R1012 VTAIL.n228 VTAIL.n227 9.3005
R1013 VTAIL.n243 VTAIL.n242 9.3005
R1014 VTAIL.n245 VTAIL.n244 9.3005
R1015 VTAIL.n224 VTAIL.n223 9.3005
R1016 VTAIL.n252 VTAIL.n251 9.3005
R1017 VTAIL.n254 VTAIL.n253 9.3005
R1018 VTAIL.n277 VTAIL.n276 9.3005
R1019 VTAIL.n2 VTAIL.n1 9.3005
R1020 VTAIL.n61 VTAIL.n60 9.3005
R1021 VTAIL.n59 VTAIL.n58 9.3005
R1022 VTAIL.n6 VTAIL.n5 9.3005
R1023 VTAIL.n53 VTAIL.n52 9.3005
R1024 VTAIL.n51 VTAIL.n50 9.3005
R1025 VTAIL.n10 VTAIL.n9 9.3005
R1026 VTAIL.n25 VTAIL.n24 9.3005
R1027 VTAIL.n27 VTAIL.n26 9.3005
R1028 VTAIL.n18 VTAIL.n17 9.3005
R1029 VTAIL.n33 VTAIL.n32 9.3005
R1030 VTAIL.n35 VTAIL.n34 9.3005
R1031 VTAIL.n14 VTAIL.n13 9.3005
R1032 VTAIL.n42 VTAIL.n41 9.3005
R1033 VTAIL.n44 VTAIL.n43 9.3005
R1034 VTAIL.n67 VTAIL.n66 9.3005
R1035 VTAIL.n166 VTAIL.n165 9.3005
R1036 VTAIL.n168 VTAIL.n167 9.3005
R1037 VTAIL.n159 VTAIL.n158 9.3005
R1038 VTAIL.n174 VTAIL.n173 9.3005
R1039 VTAIL.n176 VTAIL.n175 9.3005
R1040 VTAIL.n154 VTAIL.n153 9.3005
R1041 VTAIL.n182 VTAIL.n181 9.3005
R1042 VTAIL.n184 VTAIL.n183 9.3005
R1043 VTAIL.n207 VTAIL.n206 9.3005
R1044 VTAIL.n142 VTAIL.n141 9.3005
R1045 VTAIL.n201 VTAIL.n200 9.3005
R1046 VTAIL.n199 VTAIL.n198 9.3005
R1047 VTAIL.n146 VTAIL.n145 9.3005
R1048 VTAIL.n193 VTAIL.n192 9.3005
R1049 VTAIL.n191 VTAIL.n190 9.3005
R1050 VTAIL.n150 VTAIL.n149 9.3005
R1051 VTAIL.n96 VTAIL.n95 9.3005
R1052 VTAIL.n98 VTAIL.n97 9.3005
R1053 VTAIL.n89 VTAIL.n88 9.3005
R1054 VTAIL.n104 VTAIL.n103 9.3005
R1055 VTAIL.n106 VTAIL.n105 9.3005
R1056 VTAIL.n84 VTAIL.n83 9.3005
R1057 VTAIL.n112 VTAIL.n111 9.3005
R1058 VTAIL.n114 VTAIL.n113 9.3005
R1059 VTAIL.n137 VTAIL.n136 9.3005
R1060 VTAIL.n72 VTAIL.n71 9.3005
R1061 VTAIL.n131 VTAIL.n130 9.3005
R1062 VTAIL.n129 VTAIL.n128 9.3005
R1063 VTAIL.n76 VTAIL.n75 9.3005
R1064 VTAIL.n123 VTAIL.n122 9.3005
R1065 VTAIL.n121 VTAIL.n120 9.3005
R1066 VTAIL.n80 VTAIL.n79 9.3005
R1067 VTAIL.n238 VTAIL.n228 8.92171
R1068 VTAIL.n272 VTAIL.n271 8.92171
R1069 VTAIL.n28 VTAIL.n18 8.92171
R1070 VTAIL.n62 VTAIL.n61 8.92171
R1071 VTAIL.n202 VTAIL.n201 8.92171
R1072 VTAIL.n169 VTAIL.n159 8.92171
R1073 VTAIL.n132 VTAIL.n131 8.92171
R1074 VTAIL.n99 VTAIL.n89 8.92171
R1075 VTAIL.n237 VTAIL.n230 8.14595
R1076 VTAIL.n275 VTAIL.n212 8.14595
R1077 VTAIL.n27 VTAIL.n20 8.14595
R1078 VTAIL.n65 VTAIL.n2 8.14595
R1079 VTAIL.n205 VTAIL.n142 8.14595
R1080 VTAIL.n168 VTAIL.n161 8.14595
R1081 VTAIL.n135 VTAIL.n72 8.14595
R1082 VTAIL.n98 VTAIL.n91 8.14595
R1083 VTAIL.n234 VTAIL.n233 7.3702
R1084 VTAIL.n276 VTAIL.n210 7.3702
R1085 VTAIL.n24 VTAIL.n23 7.3702
R1086 VTAIL.n66 VTAIL.n0 7.3702
R1087 VTAIL.n206 VTAIL.n140 7.3702
R1088 VTAIL.n165 VTAIL.n164 7.3702
R1089 VTAIL.n136 VTAIL.n70 7.3702
R1090 VTAIL.n95 VTAIL.n94 7.3702
R1091 VTAIL.n278 VTAIL.n210 6.59444
R1092 VTAIL.n68 VTAIL.n0 6.59444
R1093 VTAIL.n208 VTAIL.n140 6.59444
R1094 VTAIL.n138 VTAIL.n70 6.59444
R1095 VTAIL.n234 VTAIL.n230 5.81868
R1096 VTAIL.n276 VTAIL.n275 5.81868
R1097 VTAIL.n24 VTAIL.n20 5.81868
R1098 VTAIL.n66 VTAIL.n65 5.81868
R1099 VTAIL.n206 VTAIL.n205 5.81868
R1100 VTAIL.n165 VTAIL.n161 5.81868
R1101 VTAIL.n136 VTAIL.n135 5.81868
R1102 VTAIL.n95 VTAIL.n91 5.81868
R1103 VTAIL.n238 VTAIL.n237 5.04292
R1104 VTAIL.n272 VTAIL.n212 5.04292
R1105 VTAIL.n28 VTAIL.n27 5.04292
R1106 VTAIL.n62 VTAIL.n2 5.04292
R1107 VTAIL.n202 VTAIL.n142 5.04292
R1108 VTAIL.n169 VTAIL.n168 5.04292
R1109 VTAIL.n132 VTAIL.n72 5.04292
R1110 VTAIL.n99 VTAIL.n98 5.04292
R1111 VTAIL.n241 VTAIL.n228 4.26717
R1112 VTAIL.n271 VTAIL.n214 4.26717
R1113 VTAIL.n31 VTAIL.n18 4.26717
R1114 VTAIL.n61 VTAIL.n4 4.26717
R1115 VTAIL.n201 VTAIL.n144 4.26717
R1116 VTAIL.n172 VTAIL.n159 4.26717
R1117 VTAIL.n131 VTAIL.n74 4.26717
R1118 VTAIL.n102 VTAIL.n89 4.26717
R1119 VTAIL.n242 VTAIL.n226 3.49141
R1120 VTAIL.n268 VTAIL.n267 3.49141
R1121 VTAIL.n32 VTAIL.n16 3.49141
R1122 VTAIL.n58 VTAIL.n57 3.49141
R1123 VTAIL.n198 VTAIL.n197 3.49141
R1124 VTAIL.n173 VTAIL.n157 3.49141
R1125 VTAIL.n128 VTAIL.n127 3.49141
R1126 VTAIL.n103 VTAIL.n87 3.49141
R1127 VTAIL.n246 VTAIL.n245 2.71565
R1128 VTAIL.n264 VTAIL.n216 2.71565
R1129 VTAIL.n36 VTAIL.n35 2.71565
R1130 VTAIL.n54 VTAIL.n6 2.71565
R1131 VTAIL.n194 VTAIL.n146 2.71565
R1132 VTAIL.n177 VTAIL.n176 2.71565
R1133 VTAIL.n124 VTAIL.n76 2.71565
R1134 VTAIL.n107 VTAIL.n106 2.71565
R1135 VTAIL.n235 VTAIL.n231 2.41282
R1136 VTAIL.n25 VTAIL.n21 2.41282
R1137 VTAIL.n166 VTAIL.n162 2.41282
R1138 VTAIL.n96 VTAIL.n92 2.41282
R1139 VTAIL.n250 VTAIL.n224 1.93989
R1140 VTAIL.n263 VTAIL.n218 1.93989
R1141 VTAIL.n40 VTAIL.n14 1.93989
R1142 VTAIL.n53 VTAIL.n8 1.93989
R1143 VTAIL.n193 VTAIL.n148 1.93989
R1144 VTAIL.n180 VTAIL.n154 1.93989
R1145 VTAIL.n123 VTAIL.n78 1.93989
R1146 VTAIL.n110 VTAIL.n84 1.93989
R1147 VTAIL.n251 VTAIL.n222 1.16414
R1148 VTAIL.n260 VTAIL.n259 1.16414
R1149 VTAIL.n41 VTAIL.n12 1.16414
R1150 VTAIL.n50 VTAIL.n49 1.16414
R1151 VTAIL.n190 VTAIL.n189 1.16414
R1152 VTAIL.n181 VTAIL.n152 1.16414
R1153 VTAIL.n120 VTAIL.n119 1.16414
R1154 VTAIL.n111 VTAIL.n82 1.16414
R1155 VTAIL.n209 VTAIL.n139 0.978948
R1156 VTAIL VTAIL.n69 0.782828
R1157 VTAIL.n255 VTAIL.n254 0.388379
R1158 VTAIL.n256 VTAIL.n220 0.388379
R1159 VTAIL.n45 VTAIL.n44 0.388379
R1160 VTAIL.n46 VTAIL.n10 0.388379
R1161 VTAIL.n186 VTAIL.n150 0.388379
R1162 VTAIL.n185 VTAIL.n184 0.388379
R1163 VTAIL.n116 VTAIL.n80 0.388379
R1164 VTAIL.n115 VTAIL.n114 0.388379
R1165 VTAIL VTAIL.n279 0.196621
R1166 VTAIL.n236 VTAIL.n235 0.155672
R1167 VTAIL.n236 VTAIL.n227 0.155672
R1168 VTAIL.n243 VTAIL.n227 0.155672
R1169 VTAIL.n244 VTAIL.n243 0.155672
R1170 VTAIL.n244 VTAIL.n223 0.155672
R1171 VTAIL.n252 VTAIL.n223 0.155672
R1172 VTAIL.n253 VTAIL.n252 0.155672
R1173 VTAIL.n253 VTAIL.n219 0.155672
R1174 VTAIL.n261 VTAIL.n219 0.155672
R1175 VTAIL.n262 VTAIL.n261 0.155672
R1176 VTAIL.n262 VTAIL.n215 0.155672
R1177 VTAIL.n269 VTAIL.n215 0.155672
R1178 VTAIL.n270 VTAIL.n269 0.155672
R1179 VTAIL.n270 VTAIL.n211 0.155672
R1180 VTAIL.n277 VTAIL.n211 0.155672
R1181 VTAIL.n26 VTAIL.n25 0.155672
R1182 VTAIL.n26 VTAIL.n17 0.155672
R1183 VTAIL.n33 VTAIL.n17 0.155672
R1184 VTAIL.n34 VTAIL.n33 0.155672
R1185 VTAIL.n34 VTAIL.n13 0.155672
R1186 VTAIL.n42 VTAIL.n13 0.155672
R1187 VTAIL.n43 VTAIL.n42 0.155672
R1188 VTAIL.n43 VTAIL.n9 0.155672
R1189 VTAIL.n51 VTAIL.n9 0.155672
R1190 VTAIL.n52 VTAIL.n51 0.155672
R1191 VTAIL.n52 VTAIL.n5 0.155672
R1192 VTAIL.n59 VTAIL.n5 0.155672
R1193 VTAIL.n60 VTAIL.n59 0.155672
R1194 VTAIL.n60 VTAIL.n1 0.155672
R1195 VTAIL.n67 VTAIL.n1 0.155672
R1196 VTAIL.n207 VTAIL.n141 0.155672
R1197 VTAIL.n200 VTAIL.n141 0.155672
R1198 VTAIL.n200 VTAIL.n199 0.155672
R1199 VTAIL.n199 VTAIL.n145 0.155672
R1200 VTAIL.n192 VTAIL.n145 0.155672
R1201 VTAIL.n192 VTAIL.n191 0.155672
R1202 VTAIL.n191 VTAIL.n149 0.155672
R1203 VTAIL.n183 VTAIL.n149 0.155672
R1204 VTAIL.n183 VTAIL.n182 0.155672
R1205 VTAIL.n182 VTAIL.n153 0.155672
R1206 VTAIL.n175 VTAIL.n153 0.155672
R1207 VTAIL.n175 VTAIL.n174 0.155672
R1208 VTAIL.n174 VTAIL.n158 0.155672
R1209 VTAIL.n167 VTAIL.n158 0.155672
R1210 VTAIL.n167 VTAIL.n166 0.155672
R1211 VTAIL.n137 VTAIL.n71 0.155672
R1212 VTAIL.n130 VTAIL.n71 0.155672
R1213 VTAIL.n130 VTAIL.n129 0.155672
R1214 VTAIL.n129 VTAIL.n75 0.155672
R1215 VTAIL.n122 VTAIL.n75 0.155672
R1216 VTAIL.n122 VTAIL.n121 0.155672
R1217 VTAIL.n121 VTAIL.n79 0.155672
R1218 VTAIL.n113 VTAIL.n79 0.155672
R1219 VTAIL.n113 VTAIL.n112 0.155672
R1220 VTAIL.n112 VTAIL.n83 0.155672
R1221 VTAIL.n105 VTAIL.n83 0.155672
R1222 VTAIL.n105 VTAIL.n104 0.155672
R1223 VTAIL.n104 VTAIL.n88 0.155672
R1224 VTAIL.n97 VTAIL.n88 0.155672
R1225 VTAIL.n97 VTAIL.n96 0.155672
R1226 VDD2.n133 VDD2.n69 756.745
R1227 VDD2.n64 VDD2.n0 756.745
R1228 VDD2.n134 VDD2.n133 585
R1229 VDD2.n132 VDD2.n131 585
R1230 VDD2.n73 VDD2.n72 585
R1231 VDD2.n126 VDD2.n125 585
R1232 VDD2.n124 VDD2.n123 585
R1233 VDD2.n77 VDD2.n76 585
R1234 VDD2.n118 VDD2.n117 585
R1235 VDD2.n116 VDD2.n115 585
R1236 VDD2.n114 VDD2.n80 585
R1237 VDD2.n84 VDD2.n81 585
R1238 VDD2.n109 VDD2.n108 585
R1239 VDD2.n107 VDD2.n106 585
R1240 VDD2.n86 VDD2.n85 585
R1241 VDD2.n101 VDD2.n100 585
R1242 VDD2.n99 VDD2.n98 585
R1243 VDD2.n90 VDD2.n89 585
R1244 VDD2.n93 VDD2.n92 585
R1245 VDD2.n23 VDD2.n22 585
R1246 VDD2.n20 VDD2.n19 585
R1247 VDD2.n29 VDD2.n28 585
R1248 VDD2.n31 VDD2.n30 585
R1249 VDD2.n16 VDD2.n15 585
R1250 VDD2.n37 VDD2.n36 585
R1251 VDD2.n40 VDD2.n39 585
R1252 VDD2.n38 VDD2.n12 585
R1253 VDD2.n45 VDD2.n11 585
R1254 VDD2.n47 VDD2.n46 585
R1255 VDD2.n49 VDD2.n48 585
R1256 VDD2.n8 VDD2.n7 585
R1257 VDD2.n55 VDD2.n54 585
R1258 VDD2.n57 VDD2.n56 585
R1259 VDD2.n4 VDD2.n3 585
R1260 VDD2.n63 VDD2.n62 585
R1261 VDD2.n65 VDD2.n64 585
R1262 VDD2.t1 VDD2.n21 329.036
R1263 VDD2.t0 VDD2.n91 329.036
R1264 VDD2.n133 VDD2.n132 171.744
R1265 VDD2.n132 VDD2.n72 171.744
R1266 VDD2.n125 VDD2.n72 171.744
R1267 VDD2.n125 VDD2.n124 171.744
R1268 VDD2.n124 VDD2.n76 171.744
R1269 VDD2.n117 VDD2.n76 171.744
R1270 VDD2.n117 VDD2.n116 171.744
R1271 VDD2.n116 VDD2.n80 171.744
R1272 VDD2.n84 VDD2.n80 171.744
R1273 VDD2.n108 VDD2.n84 171.744
R1274 VDD2.n108 VDD2.n107 171.744
R1275 VDD2.n107 VDD2.n85 171.744
R1276 VDD2.n100 VDD2.n85 171.744
R1277 VDD2.n100 VDD2.n99 171.744
R1278 VDD2.n99 VDD2.n89 171.744
R1279 VDD2.n92 VDD2.n89 171.744
R1280 VDD2.n22 VDD2.n19 171.744
R1281 VDD2.n29 VDD2.n19 171.744
R1282 VDD2.n30 VDD2.n29 171.744
R1283 VDD2.n30 VDD2.n15 171.744
R1284 VDD2.n37 VDD2.n15 171.744
R1285 VDD2.n39 VDD2.n37 171.744
R1286 VDD2.n39 VDD2.n38 171.744
R1287 VDD2.n38 VDD2.n11 171.744
R1288 VDD2.n47 VDD2.n11 171.744
R1289 VDD2.n48 VDD2.n47 171.744
R1290 VDD2.n48 VDD2.n7 171.744
R1291 VDD2.n55 VDD2.n7 171.744
R1292 VDD2.n56 VDD2.n55 171.744
R1293 VDD2.n56 VDD2.n3 171.744
R1294 VDD2.n63 VDD2.n3 171.744
R1295 VDD2.n64 VDD2.n63 171.744
R1296 VDD2.n138 VDD2.n68 86.2519
R1297 VDD2.n92 VDD2.t0 85.8723
R1298 VDD2.n22 VDD2.t1 85.8723
R1299 VDD2.n138 VDD2.n137 49.446
R1300 VDD2.n115 VDD2.n114 13.1884
R1301 VDD2.n46 VDD2.n45 13.1884
R1302 VDD2.n118 VDD2.n79 12.8005
R1303 VDD2.n113 VDD2.n81 12.8005
R1304 VDD2.n44 VDD2.n12 12.8005
R1305 VDD2.n49 VDD2.n10 12.8005
R1306 VDD2.n119 VDD2.n77 12.0247
R1307 VDD2.n110 VDD2.n109 12.0247
R1308 VDD2.n41 VDD2.n40 12.0247
R1309 VDD2.n50 VDD2.n8 12.0247
R1310 VDD2.n123 VDD2.n122 11.249
R1311 VDD2.n106 VDD2.n83 11.249
R1312 VDD2.n36 VDD2.n14 11.249
R1313 VDD2.n54 VDD2.n53 11.249
R1314 VDD2.n93 VDD2.n91 10.7239
R1315 VDD2.n23 VDD2.n21 10.7239
R1316 VDD2.n126 VDD2.n75 10.4732
R1317 VDD2.n105 VDD2.n86 10.4732
R1318 VDD2.n35 VDD2.n16 10.4732
R1319 VDD2.n57 VDD2.n6 10.4732
R1320 VDD2.n127 VDD2.n73 9.69747
R1321 VDD2.n102 VDD2.n101 9.69747
R1322 VDD2.n32 VDD2.n31 9.69747
R1323 VDD2.n58 VDD2.n4 9.69747
R1324 VDD2.n137 VDD2.n136 9.45567
R1325 VDD2.n68 VDD2.n67 9.45567
R1326 VDD2.n95 VDD2.n94 9.3005
R1327 VDD2.n97 VDD2.n96 9.3005
R1328 VDD2.n88 VDD2.n87 9.3005
R1329 VDD2.n103 VDD2.n102 9.3005
R1330 VDD2.n105 VDD2.n104 9.3005
R1331 VDD2.n83 VDD2.n82 9.3005
R1332 VDD2.n111 VDD2.n110 9.3005
R1333 VDD2.n113 VDD2.n112 9.3005
R1334 VDD2.n136 VDD2.n135 9.3005
R1335 VDD2.n71 VDD2.n70 9.3005
R1336 VDD2.n130 VDD2.n129 9.3005
R1337 VDD2.n128 VDD2.n127 9.3005
R1338 VDD2.n75 VDD2.n74 9.3005
R1339 VDD2.n122 VDD2.n121 9.3005
R1340 VDD2.n120 VDD2.n119 9.3005
R1341 VDD2.n79 VDD2.n78 9.3005
R1342 VDD2.n2 VDD2.n1 9.3005
R1343 VDD2.n61 VDD2.n60 9.3005
R1344 VDD2.n59 VDD2.n58 9.3005
R1345 VDD2.n6 VDD2.n5 9.3005
R1346 VDD2.n53 VDD2.n52 9.3005
R1347 VDD2.n51 VDD2.n50 9.3005
R1348 VDD2.n10 VDD2.n9 9.3005
R1349 VDD2.n25 VDD2.n24 9.3005
R1350 VDD2.n27 VDD2.n26 9.3005
R1351 VDD2.n18 VDD2.n17 9.3005
R1352 VDD2.n33 VDD2.n32 9.3005
R1353 VDD2.n35 VDD2.n34 9.3005
R1354 VDD2.n14 VDD2.n13 9.3005
R1355 VDD2.n42 VDD2.n41 9.3005
R1356 VDD2.n44 VDD2.n43 9.3005
R1357 VDD2.n67 VDD2.n66 9.3005
R1358 VDD2.n131 VDD2.n130 8.92171
R1359 VDD2.n98 VDD2.n88 8.92171
R1360 VDD2.n28 VDD2.n18 8.92171
R1361 VDD2.n62 VDD2.n61 8.92171
R1362 VDD2.n134 VDD2.n71 8.14595
R1363 VDD2.n97 VDD2.n90 8.14595
R1364 VDD2.n27 VDD2.n20 8.14595
R1365 VDD2.n65 VDD2.n2 8.14595
R1366 VDD2.n135 VDD2.n69 7.3702
R1367 VDD2.n94 VDD2.n93 7.3702
R1368 VDD2.n24 VDD2.n23 7.3702
R1369 VDD2.n66 VDD2.n0 7.3702
R1370 VDD2.n137 VDD2.n69 6.59444
R1371 VDD2.n68 VDD2.n0 6.59444
R1372 VDD2.n135 VDD2.n134 5.81868
R1373 VDD2.n94 VDD2.n90 5.81868
R1374 VDD2.n24 VDD2.n20 5.81868
R1375 VDD2.n66 VDD2.n65 5.81868
R1376 VDD2.n131 VDD2.n71 5.04292
R1377 VDD2.n98 VDD2.n97 5.04292
R1378 VDD2.n28 VDD2.n27 5.04292
R1379 VDD2.n62 VDD2.n2 5.04292
R1380 VDD2.n130 VDD2.n73 4.26717
R1381 VDD2.n101 VDD2.n88 4.26717
R1382 VDD2.n31 VDD2.n18 4.26717
R1383 VDD2.n61 VDD2.n4 4.26717
R1384 VDD2.n127 VDD2.n126 3.49141
R1385 VDD2.n102 VDD2.n86 3.49141
R1386 VDD2.n32 VDD2.n16 3.49141
R1387 VDD2.n58 VDD2.n57 3.49141
R1388 VDD2.n123 VDD2.n75 2.71565
R1389 VDD2.n106 VDD2.n105 2.71565
R1390 VDD2.n36 VDD2.n35 2.71565
R1391 VDD2.n54 VDD2.n6 2.71565
R1392 VDD2.n95 VDD2.n91 2.41282
R1393 VDD2.n25 VDD2.n21 2.41282
R1394 VDD2.n122 VDD2.n77 1.93989
R1395 VDD2.n109 VDD2.n83 1.93989
R1396 VDD2.n40 VDD2.n14 1.93989
R1397 VDD2.n53 VDD2.n8 1.93989
R1398 VDD2.n119 VDD2.n118 1.16414
R1399 VDD2.n110 VDD2.n81 1.16414
R1400 VDD2.n41 VDD2.n12 1.16414
R1401 VDD2.n50 VDD2.n49 1.16414
R1402 VDD2.n115 VDD2.n79 0.388379
R1403 VDD2.n114 VDD2.n113 0.388379
R1404 VDD2.n45 VDD2.n44 0.388379
R1405 VDD2.n46 VDD2.n10 0.388379
R1406 VDD2 VDD2.n138 0.313
R1407 VDD2.n136 VDD2.n70 0.155672
R1408 VDD2.n129 VDD2.n70 0.155672
R1409 VDD2.n129 VDD2.n128 0.155672
R1410 VDD2.n128 VDD2.n74 0.155672
R1411 VDD2.n121 VDD2.n74 0.155672
R1412 VDD2.n121 VDD2.n120 0.155672
R1413 VDD2.n120 VDD2.n78 0.155672
R1414 VDD2.n112 VDD2.n78 0.155672
R1415 VDD2.n112 VDD2.n111 0.155672
R1416 VDD2.n111 VDD2.n82 0.155672
R1417 VDD2.n104 VDD2.n82 0.155672
R1418 VDD2.n104 VDD2.n103 0.155672
R1419 VDD2.n103 VDD2.n87 0.155672
R1420 VDD2.n96 VDD2.n87 0.155672
R1421 VDD2.n96 VDD2.n95 0.155672
R1422 VDD2.n26 VDD2.n25 0.155672
R1423 VDD2.n26 VDD2.n17 0.155672
R1424 VDD2.n33 VDD2.n17 0.155672
R1425 VDD2.n34 VDD2.n33 0.155672
R1426 VDD2.n34 VDD2.n13 0.155672
R1427 VDD2.n42 VDD2.n13 0.155672
R1428 VDD2.n43 VDD2.n42 0.155672
R1429 VDD2.n43 VDD2.n9 0.155672
R1430 VDD2.n51 VDD2.n9 0.155672
R1431 VDD2.n52 VDD2.n51 0.155672
R1432 VDD2.n52 VDD2.n5 0.155672
R1433 VDD2.n59 VDD2.n5 0.155672
R1434 VDD2.n60 VDD2.n59 0.155672
R1435 VDD2.n60 VDD2.n1 0.155672
R1436 VDD2.n67 VDD2.n1 0.155672
R1437 VP.n0 VP.t0 613.391
R1438 VP.n0 VP.t1 572.702
R1439 VP VP.n0 0.0516364
R1440 VDD1.n64 VDD1.n0 756.745
R1441 VDD1.n133 VDD1.n69 756.745
R1442 VDD1.n65 VDD1.n64 585
R1443 VDD1.n63 VDD1.n62 585
R1444 VDD1.n4 VDD1.n3 585
R1445 VDD1.n57 VDD1.n56 585
R1446 VDD1.n55 VDD1.n54 585
R1447 VDD1.n8 VDD1.n7 585
R1448 VDD1.n49 VDD1.n48 585
R1449 VDD1.n47 VDD1.n46 585
R1450 VDD1.n45 VDD1.n11 585
R1451 VDD1.n15 VDD1.n12 585
R1452 VDD1.n40 VDD1.n39 585
R1453 VDD1.n38 VDD1.n37 585
R1454 VDD1.n17 VDD1.n16 585
R1455 VDD1.n32 VDD1.n31 585
R1456 VDD1.n30 VDD1.n29 585
R1457 VDD1.n21 VDD1.n20 585
R1458 VDD1.n24 VDD1.n23 585
R1459 VDD1.n92 VDD1.n91 585
R1460 VDD1.n89 VDD1.n88 585
R1461 VDD1.n98 VDD1.n97 585
R1462 VDD1.n100 VDD1.n99 585
R1463 VDD1.n85 VDD1.n84 585
R1464 VDD1.n106 VDD1.n105 585
R1465 VDD1.n109 VDD1.n108 585
R1466 VDD1.n107 VDD1.n81 585
R1467 VDD1.n114 VDD1.n80 585
R1468 VDD1.n116 VDD1.n115 585
R1469 VDD1.n118 VDD1.n117 585
R1470 VDD1.n77 VDD1.n76 585
R1471 VDD1.n124 VDD1.n123 585
R1472 VDD1.n126 VDD1.n125 585
R1473 VDD1.n73 VDD1.n72 585
R1474 VDD1.n132 VDD1.n131 585
R1475 VDD1.n134 VDD1.n133 585
R1476 VDD1.t0 VDD1.n90 329.036
R1477 VDD1.t1 VDD1.n22 329.036
R1478 VDD1.n64 VDD1.n63 171.744
R1479 VDD1.n63 VDD1.n3 171.744
R1480 VDD1.n56 VDD1.n3 171.744
R1481 VDD1.n56 VDD1.n55 171.744
R1482 VDD1.n55 VDD1.n7 171.744
R1483 VDD1.n48 VDD1.n7 171.744
R1484 VDD1.n48 VDD1.n47 171.744
R1485 VDD1.n47 VDD1.n11 171.744
R1486 VDD1.n15 VDD1.n11 171.744
R1487 VDD1.n39 VDD1.n15 171.744
R1488 VDD1.n39 VDD1.n38 171.744
R1489 VDD1.n38 VDD1.n16 171.744
R1490 VDD1.n31 VDD1.n16 171.744
R1491 VDD1.n31 VDD1.n30 171.744
R1492 VDD1.n30 VDD1.n20 171.744
R1493 VDD1.n23 VDD1.n20 171.744
R1494 VDD1.n91 VDD1.n88 171.744
R1495 VDD1.n98 VDD1.n88 171.744
R1496 VDD1.n99 VDD1.n98 171.744
R1497 VDD1.n99 VDD1.n84 171.744
R1498 VDD1.n106 VDD1.n84 171.744
R1499 VDD1.n108 VDD1.n106 171.744
R1500 VDD1.n108 VDD1.n107 171.744
R1501 VDD1.n107 VDD1.n80 171.744
R1502 VDD1.n116 VDD1.n80 171.744
R1503 VDD1.n117 VDD1.n116 171.744
R1504 VDD1.n117 VDD1.n76 171.744
R1505 VDD1.n124 VDD1.n76 171.744
R1506 VDD1.n125 VDD1.n124 171.744
R1507 VDD1.n125 VDD1.n72 171.744
R1508 VDD1.n132 VDD1.n72 171.744
R1509 VDD1.n133 VDD1.n132 171.744
R1510 VDD1 VDD1.n137 87.0311
R1511 VDD1.n23 VDD1.t1 85.8723
R1512 VDD1.n91 VDD1.t0 85.8723
R1513 VDD1 VDD1.n68 49.7585
R1514 VDD1.n46 VDD1.n45 13.1884
R1515 VDD1.n115 VDD1.n114 13.1884
R1516 VDD1.n49 VDD1.n10 12.8005
R1517 VDD1.n44 VDD1.n12 12.8005
R1518 VDD1.n113 VDD1.n81 12.8005
R1519 VDD1.n118 VDD1.n79 12.8005
R1520 VDD1.n50 VDD1.n8 12.0247
R1521 VDD1.n41 VDD1.n40 12.0247
R1522 VDD1.n110 VDD1.n109 12.0247
R1523 VDD1.n119 VDD1.n77 12.0247
R1524 VDD1.n54 VDD1.n53 11.249
R1525 VDD1.n37 VDD1.n14 11.249
R1526 VDD1.n105 VDD1.n83 11.249
R1527 VDD1.n123 VDD1.n122 11.249
R1528 VDD1.n24 VDD1.n22 10.7239
R1529 VDD1.n92 VDD1.n90 10.7239
R1530 VDD1.n57 VDD1.n6 10.4732
R1531 VDD1.n36 VDD1.n17 10.4732
R1532 VDD1.n104 VDD1.n85 10.4732
R1533 VDD1.n126 VDD1.n75 10.4732
R1534 VDD1.n58 VDD1.n4 9.69747
R1535 VDD1.n33 VDD1.n32 9.69747
R1536 VDD1.n101 VDD1.n100 9.69747
R1537 VDD1.n127 VDD1.n73 9.69747
R1538 VDD1.n68 VDD1.n67 9.45567
R1539 VDD1.n137 VDD1.n136 9.45567
R1540 VDD1.n26 VDD1.n25 9.3005
R1541 VDD1.n28 VDD1.n27 9.3005
R1542 VDD1.n19 VDD1.n18 9.3005
R1543 VDD1.n34 VDD1.n33 9.3005
R1544 VDD1.n36 VDD1.n35 9.3005
R1545 VDD1.n14 VDD1.n13 9.3005
R1546 VDD1.n42 VDD1.n41 9.3005
R1547 VDD1.n44 VDD1.n43 9.3005
R1548 VDD1.n67 VDD1.n66 9.3005
R1549 VDD1.n2 VDD1.n1 9.3005
R1550 VDD1.n61 VDD1.n60 9.3005
R1551 VDD1.n59 VDD1.n58 9.3005
R1552 VDD1.n6 VDD1.n5 9.3005
R1553 VDD1.n53 VDD1.n52 9.3005
R1554 VDD1.n51 VDD1.n50 9.3005
R1555 VDD1.n10 VDD1.n9 9.3005
R1556 VDD1.n71 VDD1.n70 9.3005
R1557 VDD1.n130 VDD1.n129 9.3005
R1558 VDD1.n128 VDD1.n127 9.3005
R1559 VDD1.n75 VDD1.n74 9.3005
R1560 VDD1.n122 VDD1.n121 9.3005
R1561 VDD1.n120 VDD1.n119 9.3005
R1562 VDD1.n79 VDD1.n78 9.3005
R1563 VDD1.n94 VDD1.n93 9.3005
R1564 VDD1.n96 VDD1.n95 9.3005
R1565 VDD1.n87 VDD1.n86 9.3005
R1566 VDD1.n102 VDD1.n101 9.3005
R1567 VDD1.n104 VDD1.n103 9.3005
R1568 VDD1.n83 VDD1.n82 9.3005
R1569 VDD1.n111 VDD1.n110 9.3005
R1570 VDD1.n113 VDD1.n112 9.3005
R1571 VDD1.n136 VDD1.n135 9.3005
R1572 VDD1.n62 VDD1.n61 8.92171
R1573 VDD1.n29 VDD1.n19 8.92171
R1574 VDD1.n97 VDD1.n87 8.92171
R1575 VDD1.n131 VDD1.n130 8.92171
R1576 VDD1.n65 VDD1.n2 8.14595
R1577 VDD1.n28 VDD1.n21 8.14595
R1578 VDD1.n96 VDD1.n89 8.14595
R1579 VDD1.n134 VDD1.n71 8.14595
R1580 VDD1.n66 VDD1.n0 7.3702
R1581 VDD1.n25 VDD1.n24 7.3702
R1582 VDD1.n93 VDD1.n92 7.3702
R1583 VDD1.n135 VDD1.n69 7.3702
R1584 VDD1.n68 VDD1.n0 6.59444
R1585 VDD1.n137 VDD1.n69 6.59444
R1586 VDD1.n66 VDD1.n65 5.81868
R1587 VDD1.n25 VDD1.n21 5.81868
R1588 VDD1.n93 VDD1.n89 5.81868
R1589 VDD1.n135 VDD1.n134 5.81868
R1590 VDD1.n62 VDD1.n2 5.04292
R1591 VDD1.n29 VDD1.n28 5.04292
R1592 VDD1.n97 VDD1.n96 5.04292
R1593 VDD1.n131 VDD1.n71 5.04292
R1594 VDD1.n61 VDD1.n4 4.26717
R1595 VDD1.n32 VDD1.n19 4.26717
R1596 VDD1.n100 VDD1.n87 4.26717
R1597 VDD1.n130 VDD1.n73 4.26717
R1598 VDD1.n58 VDD1.n57 3.49141
R1599 VDD1.n33 VDD1.n17 3.49141
R1600 VDD1.n101 VDD1.n85 3.49141
R1601 VDD1.n127 VDD1.n126 3.49141
R1602 VDD1.n54 VDD1.n6 2.71565
R1603 VDD1.n37 VDD1.n36 2.71565
R1604 VDD1.n105 VDD1.n104 2.71565
R1605 VDD1.n123 VDD1.n75 2.71565
R1606 VDD1.n26 VDD1.n22 2.41282
R1607 VDD1.n94 VDD1.n90 2.41282
R1608 VDD1.n53 VDD1.n8 1.93989
R1609 VDD1.n40 VDD1.n14 1.93989
R1610 VDD1.n109 VDD1.n83 1.93989
R1611 VDD1.n122 VDD1.n77 1.93989
R1612 VDD1.n50 VDD1.n49 1.16414
R1613 VDD1.n41 VDD1.n12 1.16414
R1614 VDD1.n110 VDD1.n81 1.16414
R1615 VDD1.n119 VDD1.n118 1.16414
R1616 VDD1.n46 VDD1.n10 0.388379
R1617 VDD1.n45 VDD1.n44 0.388379
R1618 VDD1.n114 VDD1.n113 0.388379
R1619 VDD1.n115 VDD1.n79 0.388379
R1620 VDD1.n67 VDD1.n1 0.155672
R1621 VDD1.n60 VDD1.n1 0.155672
R1622 VDD1.n60 VDD1.n59 0.155672
R1623 VDD1.n59 VDD1.n5 0.155672
R1624 VDD1.n52 VDD1.n5 0.155672
R1625 VDD1.n52 VDD1.n51 0.155672
R1626 VDD1.n51 VDD1.n9 0.155672
R1627 VDD1.n43 VDD1.n9 0.155672
R1628 VDD1.n43 VDD1.n42 0.155672
R1629 VDD1.n42 VDD1.n13 0.155672
R1630 VDD1.n35 VDD1.n13 0.155672
R1631 VDD1.n35 VDD1.n34 0.155672
R1632 VDD1.n34 VDD1.n18 0.155672
R1633 VDD1.n27 VDD1.n18 0.155672
R1634 VDD1.n27 VDD1.n26 0.155672
R1635 VDD1.n95 VDD1.n94 0.155672
R1636 VDD1.n95 VDD1.n86 0.155672
R1637 VDD1.n102 VDD1.n86 0.155672
R1638 VDD1.n103 VDD1.n102 0.155672
R1639 VDD1.n103 VDD1.n82 0.155672
R1640 VDD1.n111 VDD1.n82 0.155672
R1641 VDD1.n112 VDD1.n111 0.155672
R1642 VDD1.n112 VDD1.n78 0.155672
R1643 VDD1.n120 VDD1.n78 0.155672
R1644 VDD1.n121 VDD1.n120 0.155672
R1645 VDD1.n121 VDD1.n74 0.155672
R1646 VDD1.n128 VDD1.n74 0.155672
R1647 VDD1.n129 VDD1.n128 0.155672
R1648 VDD1.n129 VDD1.n70 0.155672
R1649 VDD1.n136 VDD1.n70 0.155672
C0 B w_n1442_n3546# 7.16612f
C1 VDD2 VDD1 0.47705f
C2 VDD2 VTAIL 5.78325f
C3 VDD2 VN 2.25949f
C4 VDD1 w_n1442_n3546# 1.65169f
C5 VTAIL w_n1442_n3546# 3.0297f
C6 VN w_n1442_n3546# 1.8545f
C7 B VP 1.05226f
C8 VP VDD1 2.36779f
C9 VTAIL VP 1.75256f
C10 VDD2 w_n1442_n3546# 1.65786f
C11 VP VN 4.79063f
C12 VDD2 VP 0.261355f
C13 VP w_n1442_n3546# 2.03441f
C14 B VDD1 1.50632f
C15 VTAIL B 2.9761f
C16 B VN 0.763505f
C17 VTAIL VDD1 5.74828f
C18 VDD1 VN 0.148657f
C19 VTAIL VN 1.73796f
C20 VDD2 B 1.52188f
C21 VDD2 VSUBS 0.788114f
C22 VDD1 VSUBS 3.30444f
C23 VTAIL VSUBS 0.804615f
C24 VN VSUBS 5.76138f
C25 VP VSUBS 1.187585f
C26 B VSUBS 2.680149f
C27 w_n1442_n3546# VSUBS 62.865395f
C28 VDD1.n0 VSUBS 0.023147f
C29 VDD1.n1 VSUBS 0.020588f
C30 VDD1.n2 VSUBS 0.011063f
C31 VDD1.n3 VSUBS 0.026149f
C32 VDD1.n4 VSUBS 0.011714f
C33 VDD1.n5 VSUBS 0.020588f
C34 VDD1.n6 VSUBS 0.011063f
C35 VDD1.n7 VSUBS 0.026149f
C36 VDD1.n8 VSUBS 0.011714f
C37 VDD1.n9 VSUBS 0.020588f
C38 VDD1.n10 VSUBS 0.011063f
C39 VDD1.n11 VSUBS 0.026149f
C40 VDD1.n12 VSUBS 0.011714f
C41 VDD1.n13 VSUBS 0.020588f
C42 VDD1.n14 VSUBS 0.011063f
C43 VDD1.n15 VSUBS 0.026149f
C44 VDD1.n16 VSUBS 0.026149f
C45 VDD1.n17 VSUBS 0.011714f
C46 VDD1.n18 VSUBS 0.020588f
C47 VDD1.n19 VSUBS 0.011063f
C48 VDD1.n20 VSUBS 0.026149f
C49 VDD1.n21 VSUBS 0.011714f
C50 VDD1.n22 VSUBS 0.170242f
C51 VDD1.t1 VSUBS 0.056409f
C52 VDD1.n23 VSUBS 0.019612f
C53 VDD1.n24 VSUBS 0.019671f
C54 VDD1.n25 VSUBS 0.011063f
C55 VDD1.n26 VSUBS 1.09005f
C56 VDD1.n27 VSUBS 0.020588f
C57 VDD1.n28 VSUBS 0.011063f
C58 VDD1.n29 VSUBS 0.011714f
C59 VDD1.n30 VSUBS 0.026149f
C60 VDD1.n31 VSUBS 0.026149f
C61 VDD1.n32 VSUBS 0.011714f
C62 VDD1.n33 VSUBS 0.011063f
C63 VDD1.n34 VSUBS 0.020588f
C64 VDD1.n35 VSUBS 0.020588f
C65 VDD1.n36 VSUBS 0.011063f
C66 VDD1.n37 VSUBS 0.011714f
C67 VDD1.n38 VSUBS 0.026149f
C68 VDD1.n39 VSUBS 0.026149f
C69 VDD1.n40 VSUBS 0.011714f
C70 VDD1.n41 VSUBS 0.011063f
C71 VDD1.n42 VSUBS 0.020588f
C72 VDD1.n43 VSUBS 0.020588f
C73 VDD1.n44 VSUBS 0.011063f
C74 VDD1.n45 VSUBS 0.011389f
C75 VDD1.n46 VSUBS 0.011389f
C76 VDD1.n47 VSUBS 0.026149f
C77 VDD1.n48 VSUBS 0.026149f
C78 VDD1.n49 VSUBS 0.011714f
C79 VDD1.n50 VSUBS 0.011063f
C80 VDD1.n51 VSUBS 0.020588f
C81 VDD1.n52 VSUBS 0.020588f
C82 VDD1.n53 VSUBS 0.011063f
C83 VDD1.n54 VSUBS 0.011714f
C84 VDD1.n55 VSUBS 0.026149f
C85 VDD1.n56 VSUBS 0.026149f
C86 VDD1.n57 VSUBS 0.011714f
C87 VDD1.n58 VSUBS 0.011063f
C88 VDD1.n59 VSUBS 0.020588f
C89 VDD1.n60 VSUBS 0.020588f
C90 VDD1.n61 VSUBS 0.011063f
C91 VDD1.n62 VSUBS 0.011714f
C92 VDD1.n63 VSUBS 0.026149f
C93 VDD1.n64 VSUBS 0.065092f
C94 VDD1.n65 VSUBS 0.011714f
C95 VDD1.n66 VSUBS 0.011063f
C96 VDD1.n67 VSUBS 0.048432f
C97 VDD1.n68 VSUBS 0.047431f
C98 VDD1.n69 VSUBS 0.023147f
C99 VDD1.n70 VSUBS 0.020588f
C100 VDD1.n71 VSUBS 0.011063f
C101 VDD1.n72 VSUBS 0.026149f
C102 VDD1.n73 VSUBS 0.011714f
C103 VDD1.n74 VSUBS 0.020588f
C104 VDD1.n75 VSUBS 0.011063f
C105 VDD1.n76 VSUBS 0.026149f
C106 VDD1.n77 VSUBS 0.011714f
C107 VDD1.n78 VSUBS 0.020588f
C108 VDD1.n79 VSUBS 0.011063f
C109 VDD1.n80 VSUBS 0.026149f
C110 VDD1.n81 VSUBS 0.011714f
C111 VDD1.n82 VSUBS 0.020588f
C112 VDD1.n83 VSUBS 0.011063f
C113 VDD1.n84 VSUBS 0.026149f
C114 VDD1.n85 VSUBS 0.011714f
C115 VDD1.n86 VSUBS 0.020588f
C116 VDD1.n87 VSUBS 0.011063f
C117 VDD1.n88 VSUBS 0.026149f
C118 VDD1.n89 VSUBS 0.011714f
C119 VDD1.n90 VSUBS 0.170242f
C120 VDD1.t0 VSUBS 0.056409f
C121 VDD1.n91 VSUBS 0.019612f
C122 VDD1.n92 VSUBS 0.019671f
C123 VDD1.n93 VSUBS 0.011063f
C124 VDD1.n94 VSUBS 1.09005f
C125 VDD1.n95 VSUBS 0.020588f
C126 VDD1.n96 VSUBS 0.011063f
C127 VDD1.n97 VSUBS 0.011714f
C128 VDD1.n98 VSUBS 0.026149f
C129 VDD1.n99 VSUBS 0.026149f
C130 VDD1.n100 VSUBS 0.011714f
C131 VDD1.n101 VSUBS 0.011063f
C132 VDD1.n102 VSUBS 0.020588f
C133 VDD1.n103 VSUBS 0.020588f
C134 VDD1.n104 VSUBS 0.011063f
C135 VDD1.n105 VSUBS 0.011714f
C136 VDD1.n106 VSUBS 0.026149f
C137 VDD1.n107 VSUBS 0.026149f
C138 VDD1.n108 VSUBS 0.026149f
C139 VDD1.n109 VSUBS 0.011714f
C140 VDD1.n110 VSUBS 0.011063f
C141 VDD1.n111 VSUBS 0.020588f
C142 VDD1.n112 VSUBS 0.020588f
C143 VDD1.n113 VSUBS 0.011063f
C144 VDD1.n114 VSUBS 0.011389f
C145 VDD1.n115 VSUBS 0.011389f
C146 VDD1.n116 VSUBS 0.026149f
C147 VDD1.n117 VSUBS 0.026149f
C148 VDD1.n118 VSUBS 0.011714f
C149 VDD1.n119 VSUBS 0.011063f
C150 VDD1.n120 VSUBS 0.020588f
C151 VDD1.n121 VSUBS 0.020588f
C152 VDD1.n122 VSUBS 0.011063f
C153 VDD1.n123 VSUBS 0.011714f
C154 VDD1.n124 VSUBS 0.026149f
C155 VDD1.n125 VSUBS 0.026149f
C156 VDD1.n126 VSUBS 0.011714f
C157 VDD1.n127 VSUBS 0.011063f
C158 VDD1.n128 VSUBS 0.020588f
C159 VDD1.n129 VSUBS 0.020588f
C160 VDD1.n130 VSUBS 0.011063f
C161 VDD1.n131 VSUBS 0.011714f
C162 VDD1.n132 VSUBS 0.026149f
C163 VDD1.n133 VSUBS 0.065092f
C164 VDD1.n134 VSUBS 0.011714f
C165 VDD1.n135 VSUBS 0.011063f
C166 VDD1.n136 VSUBS 0.048432f
C167 VDD1.n137 VSUBS 0.564597f
C168 VP.t0 VSUBS 2.09158f
C169 VP.t1 VSUBS 1.91512f
C170 VP.n0 VSUBS 5.16888f
C171 VDD2.n0 VSUBS 0.023366f
C172 VDD2.n1 VSUBS 0.020783f
C173 VDD2.n2 VSUBS 0.011168f
C174 VDD2.n3 VSUBS 0.026397f
C175 VDD2.n4 VSUBS 0.011825f
C176 VDD2.n5 VSUBS 0.020783f
C177 VDD2.n6 VSUBS 0.011168f
C178 VDD2.n7 VSUBS 0.026397f
C179 VDD2.n8 VSUBS 0.011825f
C180 VDD2.n9 VSUBS 0.020783f
C181 VDD2.n10 VSUBS 0.011168f
C182 VDD2.n11 VSUBS 0.026397f
C183 VDD2.n12 VSUBS 0.011825f
C184 VDD2.n13 VSUBS 0.020783f
C185 VDD2.n14 VSUBS 0.011168f
C186 VDD2.n15 VSUBS 0.026397f
C187 VDD2.n16 VSUBS 0.011825f
C188 VDD2.n17 VSUBS 0.020783f
C189 VDD2.n18 VSUBS 0.011168f
C190 VDD2.n19 VSUBS 0.026397f
C191 VDD2.n20 VSUBS 0.011825f
C192 VDD2.n21 VSUBS 0.171856f
C193 VDD2.t1 VSUBS 0.056943f
C194 VDD2.n22 VSUBS 0.019798f
C195 VDD2.n23 VSUBS 0.019857f
C196 VDD2.n24 VSUBS 0.011168f
C197 VDD2.n25 VSUBS 1.10038f
C198 VDD2.n26 VSUBS 0.020783f
C199 VDD2.n27 VSUBS 0.011168f
C200 VDD2.n28 VSUBS 0.011825f
C201 VDD2.n29 VSUBS 0.026397f
C202 VDD2.n30 VSUBS 0.026397f
C203 VDD2.n31 VSUBS 0.011825f
C204 VDD2.n32 VSUBS 0.011168f
C205 VDD2.n33 VSUBS 0.020783f
C206 VDD2.n34 VSUBS 0.020783f
C207 VDD2.n35 VSUBS 0.011168f
C208 VDD2.n36 VSUBS 0.011825f
C209 VDD2.n37 VSUBS 0.026397f
C210 VDD2.n38 VSUBS 0.026397f
C211 VDD2.n39 VSUBS 0.026397f
C212 VDD2.n40 VSUBS 0.011825f
C213 VDD2.n41 VSUBS 0.011168f
C214 VDD2.n42 VSUBS 0.020783f
C215 VDD2.n43 VSUBS 0.020783f
C216 VDD2.n44 VSUBS 0.011168f
C217 VDD2.n45 VSUBS 0.011497f
C218 VDD2.n46 VSUBS 0.011497f
C219 VDD2.n47 VSUBS 0.026397f
C220 VDD2.n48 VSUBS 0.026397f
C221 VDD2.n49 VSUBS 0.011825f
C222 VDD2.n50 VSUBS 0.011168f
C223 VDD2.n51 VSUBS 0.020783f
C224 VDD2.n52 VSUBS 0.020783f
C225 VDD2.n53 VSUBS 0.011168f
C226 VDD2.n54 VSUBS 0.011825f
C227 VDD2.n55 VSUBS 0.026397f
C228 VDD2.n56 VSUBS 0.026397f
C229 VDD2.n57 VSUBS 0.011825f
C230 VDD2.n58 VSUBS 0.011168f
C231 VDD2.n59 VSUBS 0.020783f
C232 VDD2.n60 VSUBS 0.020783f
C233 VDD2.n61 VSUBS 0.011168f
C234 VDD2.n62 VSUBS 0.011825f
C235 VDD2.n63 VSUBS 0.026397f
C236 VDD2.n64 VSUBS 0.065709f
C237 VDD2.n65 VSUBS 0.011825f
C238 VDD2.n66 VSUBS 0.011168f
C239 VDD2.n67 VSUBS 0.048891f
C240 VDD2.n68 VSUBS 0.540996f
C241 VDD2.n69 VSUBS 0.023366f
C242 VDD2.n70 VSUBS 0.020783f
C243 VDD2.n71 VSUBS 0.011168f
C244 VDD2.n72 VSUBS 0.026397f
C245 VDD2.n73 VSUBS 0.011825f
C246 VDD2.n74 VSUBS 0.020783f
C247 VDD2.n75 VSUBS 0.011168f
C248 VDD2.n76 VSUBS 0.026397f
C249 VDD2.n77 VSUBS 0.011825f
C250 VDD2.n78 VSUBS 0.020783f
C251 VDD2.n79 VSUBS 0.011168f
C252 VDD2.n80 VSUBS 0.026397f
C253 VDD2.n81 VSUBS 0.011825f
C254 VDD2.n82 VSUBS 0.020783f
C255 VDD2.n83 VSUBS 0.011168f
C256 VDD2.n84 VSUBS 0.026397f
C257 VDD2.n85 VSUBS 0.026397f
C258 VDD2.n86 VSUBS 0.011825f
C259 VDD2.n87 VSUBS 0.020783f
C260 VDD2.n88 VSUBS 0.011168f
C261 VDD2.n89 VSUBS 0.026397f
C262 VDD2.n90 VSUBS 0.011825f
C263 VDD2.n91 VSUBS 0.171856f
C264 VDD2.t0 VSUBS 0.056943f
C265 VDD2.n92 VSUBS 0.019798f
C266 VDD2.n93 VSUBS 0.019857f
C267 VDD2.n94 VSUBS 0.011168f
C268 VDD2.n95 VSUBS 1.10038f
C269 VDD2.n96 VSUBS 0.020783f
C270 VDD2.n97 VSUBS 0.011168f
C271 VDD2.n98 VSUBS 0.011825f
C272 VDD2.n99 VSUBS 0.026397f
C273 VDD2.n100 VSUBS 0.026397f
C274 VDD2.n101 VSUBS 0.011825f
C275 VDD2.n102 VSUBS 0.011168f
C276 VDD2.n103 VSUBS 0.020783f
C277 VDD2.n104 VSUBS 0.020783f
C278 VDD2.n105 VSUBS 0.011168f
C279 VDD2.n106 VSUBS 0.011825f
C280 VDD2.n107 VSUBS 0.026397f
C281 VDD2.n108 VSUBS 0.026397f
C282 VDD2.n109 VSUBS 0.011825f
C283 VDD2.n110 VSUBS 0.011168f
C284 VDD2.n111 VSUBS 0.020783f
C285 VDD2.n112 VSUBS 0.020783f
C286 VDD2.n113 VSUBS 0.011168f
C287 VDD2.n114 VSUBS 0.011497f
C288 VDD2.n115 VSUBS 0.011497f
C289 VDD2.n116 VSUBS 0.026397f
C290 VDD2.n117 VSUBS 0.026397f
C291 VDD2.n118 VSUBS 0.011825f
C292 VDD2.n119 VSUBS 0.011168f
C293 VDD2.n120 VSUBS 0.020783f
C294 VDD2.n121 VSUBS 0.020783f
C295 VDD2.n122 VSUBS 0.011168f
C296 VDD2.n123 VSUBS 0.011825f
C297 VDD2.n124 VSUBS 0.026397f
C298 VDD2.n125 VSUBS 0.026397f
C299 VDD2.n126 VSUBS 0.011825f
C300 VDD2.n127 VSUBS 0.011168f
C301 VDD2.n128 VSUBS 0.020783f
C302 VDD2.n129 VSUBS 0.020783f
C303 VDD2.n130 VSUBS 0.011168f
C304 VDD2.n131 VSUBS 0.011825f
C305 VDD2.n132 VSUBS 0.026397f
C306 VDD2.n133 VSUBS 0.065709f
C307 VDD2.n134 VSUBS 0.011825f
C308 VDD2.n135 VSUBS 0.011168f
C309 VDD2.n136 VSUBS 0.048891f
C310 VDD2.n137 VSUBS 0.047495f
C311 VDD2.n138 VSUBS 2.33403f
C312 VTAIL.n0 VSUBS 0.026856f
C313 VTAIL.n1 VSUBS 0.023887f
C314 VTAIL.n2 VSUBS 0.012836f
C315 VTAIL.n3 VSUBS 0.030339f
C316 VTAIL.n4 VSUBS 0.013591f
C317 VTAIL.n5 VSUBS 0.023887f
C318 VTAIL.n6 VSUBS 0.012836f
C319 VTAIL.n7 VSUBS 0.030339f
C320 VTAIL.n8 VSUBS 0.013591f
C321 VTAIL.n9 VSUBS 0.023887f
C322 VTAIL.n10 VSUBS 0.012836f
C323 VTAIL.n11 VSUBS 0.030339f
C324 VTAIL.n12 VSUBS 0.013591f
C325 VTAIL.n13 VSUBS 0.023887f
C326 VTAIL.n14 VSUBS 0.012836f
C327 VTAIL.n15 VSUBS 0.030339f
C328 VTAIL.n16 VSUBS 0.013591f
C329 VTAIL.n17 VSUBS 0.023887f
C330 VTAIL.n18 VSUBS 0.012836f
C331 VTAIL.n19 VSUBS 0.030339f
C332 VTAIL.n20 VSUBS 0.013591f
C333 VTAIL.n21 VSUBS 0.197521f
C334 VTAIL.t0 VSUBS 0.065447f
C335 VTAIL.n22 VSUBS 0.022755f
C336 VTAIL.n23 VSUBS 0.022823f
C337 VTAIL.n24 VSUBS 0.012836f
C338 VTAIL.n25 VSUBS 1.26471f
C339 VTAIL.n26 VSUBS 0.023887f
C340 VTAIL.n27 VSUBS 0.012836f
C341 VTAIL.n28 VSUBS 0.013591f
C342 VTAIL.n29 VSUBS 0.030339f
C343 VTAIL.n30 VSUBS 0.030339f
C344 VTAIL.n31 VSUBS 0.013591f
C345 VTAIL.n32 VSUBS 0.012836f
C346 VTAIL.n33 VSUBS 0.023887f
C347 VTAIL.n34 VSUBS 0.023887f
C348 VTAIL.n35 VSUBS 0.012836f
C349 VTAIL.n36 VSUBS 0.013591f
C350 VTAIL.n37 VSUBS 0.030339f
C351 VTAIL.n38 VSUBS 0.030339f
C352 VTAIL.n39 VSUBS 0.030339f
C353 VTAIL.n40 VSUBS 0.013591f
C354 VTAIL.n41 VSUBS 0.012836f
C355 VTAIL.n42 VSUBS 0.023887f
C356 VTAIL.n43 VSUBS 0.023887f
C357 VTAIL.n44 VSUBS 0.012836f
C358 VTAIL.n45 VSUBS 0.013213f
C359 VTAIL.n46 VSUBS 0.013213f
C360 VTAIL.n47 VSUBS 0.030339f
C361 VTAIL.n48 VSUBS 0.030339f
C362 VTAIL.n49 VSUBS 0.013591f
C363 VTAIL.n50 VSUBS 0.012836f
C364 VTAIL.n51 VSUBS 0.023887f
C365 VTAIL.n52 VSUBS 0.023887f
C366 VTAIL.n53 VSUBS 0.012836f
C367 VTAIL.n54 VSUBS 0.013591f
C368 VTAIL.n55 VSUBS 0.030339f
C369 VTAIL.n56 VSUBS 0.030339f
C370 VTAIL.n57 VSUBS 0.013591f
C371 VTAIL.n58 VSUBS 0.012836f
C372 VTAIL.n59 VSUBS 0.023887f
C373 VTAIL.n60 VSUBS 0.023887f
C374 VTAIL.n61 VSUBS 0.012836f
C375 VTAIL.n62 VSUBS 0.013591f
C376 VTAIL.n63 VSUBS 0.030339f
C377 VTAIL.n64 VSUBS 0.075523f
C378 VTAIL.n65 VSUBS 0.013591f
C379 VTAIL.n66 VSUBS 0.012836f
C380 VTAIL.n67 VSUBS 0.056193f
C381 VTAIL.n68 VSUBS 0.038102f
C382 VTAIL.n69 VSUBS 1.41754f
C383 VTAIL.n70 VSUBS 0.026856f
C384 VTAIL.n71 VSUBS 0.023887f
C385 VTAIL.n72 VSUBS 0.012836f
C386 VTAIL.n73 VSUBS 0.030339f
C387 VTAIL.n74 VSUBS 0.013591f
C388 VTAIL.n75 VSUBS 0.023887f
C389 VTAIL.n76 VSUBS 0.012836f
C390 VTAIL.n77 VSUBS 0.030339f
C391 VTAIL.n78 VSUBS 0.013591f
C392 VTAIL.n79 VSUBS 0.023887f
C393 VTAIL.n80 VSUBS 0.012836f
C394 VTAIL.n81 VSUBS 0.030339f
C395 VTAIL.n82 VSUBS 0.013591f
C396 VTAIL.n83 VSUBS 0.023887f
C397 VTAIL.n84 VSUBS 0.012836f
C398 VTAIL.n85 VSUBS 0.030339f
C399 VTAIL.n86 VSUBS 0.030339f
C400 VTAIL.n87 VSUBS 0.013591f
C401 VTAIL.n88 VSUBS 0.023887f
C402 VTAIL.n89 VSUBS 0.012836f
C403 VTAIL.n90 VSUBS 0.030339f
C404 VTAIL.n91 VSUBS 0.013591f
C405 VTAIL.n92 VSUBS 0.197521f
C406 VTAIL.t2 VSUBS 0.065447f
C407 VTAIL.n93 VSUBS 0.022755f
C408 VTAIL.n94 VSUBS 0.022823f
C409 VTAIL.n95 VSUBS 0.012836f
C410 VTAIL.n96 VSUBS 1.26471f
C411 VTAIL.n97 VSUBS 0.023887f
C412 VTAIL.n98 VSUBS 0.012836f
C413 VTAIL.n99 VSUBS 0.013591f
C414 VTAIL.n100 VSUBS 0.030339f
C415 VTAIL.n101 VSUBS 0.030339f
C416 VTAIL.n102 VSUBS 0.013591f
C417 VTAIL.n103 VSUBS 0.012836f
C418 VTAIL.n104 VSUBS 0.023887f
C419 VTAIL.n105 VSUBS 0.023887f
C420 VTAIL.n106 VSUBS 0.012836f
C421 VTAIL.n107 VSUBS 0.013591f
C422 VTAIL.n108 VSUBS 0.030339f
C423 VTAIL.n109 VSUBS 0.030339f
C424 VTAIL.n110 VSUBS 0.013591f
C425 VTAIL.n111 VSUBS 0.012836f
C426 VTAIL.n112 VSUBS 0.023887f
C427 VTAIL.n113 VSUBS 0.023887f
C428 VTAIL.n114 VSUBS 0.012836f
C429 VTAIL.n115 VSUBS 0.013213f
C430 VTAIL.n116 VSUBS 0.013213f
C431 VTAIL.n117 VSUBS 0.030339f
C432 VTAIL.n118 VSUBS 0.030339f
C433 VTAIL.n119 VSUBS 0.013591f
C434 VTAIL.n120 VSUBS 0.012836f
C435 VTAIL.n121 VSUBS 0.023887f
C436 VTAIL.n122 VSUBS 0.023887f
C437 VTAIL.n123 VSUBS 0.012836f
C438 VTAIL.n124 VSUBS 0.013591f
C439 VTAIL.n125 VSUBS 0.030339f
C440 VTAIL.n126 VSUBS 0.030339f
C441 VTAIL.n127 VSUBS 0.013591f
C442 VTAIL.n128 VSUBS 0.012836f
C443 VTAIL.n129 VSUBS 0.023887f
C444 VTAIL.n130 VSUBS 0.023887f
C445 VTAIL.n131 VSUBS 0.012836f
C446 VTAIL.n132 VSUBS 0.013591f
C447 VTAIL.n133 VSUBS 0.030339f
C448 VTAIL.n134 VSUBS 0.075523f
C449 VTAIL.n135 VSUBS 0.013591f
C450 VTAIL.n136 VSUBS 0.012836f
C451 VTAIL.n137 VSUBS 0.056193f
C452 VTAIL.n138 VSUBS 0.038102f
C453 VTAIL.n139 VSUBS 1.43263f
C454 VTAIL.n140 VSUBS 0.026856f
C455 VTAIL.n141 VSUBS 0.023887f
C456 VTAIL.n142 VSUBS 0.012836f
C457 VTAIL.n143 VSUBS 0.030339f
C458 VTAIL.n144 VSUBS 0.013591f
C459 VTAIL.n145 VSUBS 0.023887f
C460 VTAIL.n146 VSUBS 0.012836f
C461 VTAIL.n147 VSUBS 0.030339f
C462 VTAIL.n148 VSUBS 0.013591f
C463 VTAIL.n149 VSUBS 0.023887f
C464 VTAIL.n150 VSUBS 0.012836f
C465 VTAIL.n151 VSUBS 0.030339f
C466 VTAIL.n152 VSUBS 0.013591f
C467 VTAIL.n153 VSUBS 0.023887f
C468 VTAIL.n154 VSUBS 0.012836f
C469 VTAIL.n155 VSUBS 0.030339f
C470 VTAIL.n156 VSUBS 0.030339f
C471 VTAIL.n157 VSUBS 0.013591f
C472 VTAIL.n158 VSUBS 0.023887f
C473 VTAIL.n159 VSUBS 0.012836f
C474 VTAIL.n160 VSUBS 0.030339f
C475 VTAIL.n161 VSUBS 0.013591f
C476 VTAIL.n162 VSUBS 0.197521f
C477 VTAIL.t1 VSUBS 0.065447f
C478 VTAIL.n163 VSUBS 0.022755f
C479 VTAIL.n164 VSUBS 0.022823f
C480 VTAIL.n165 VSUBS 0.012836f
C481 VTAIL.n166 VSUBS 1.26471f
C482 VTAIL.n167 VSUBS 0.023887f
C483 VTAIL.n168 VSUBS 0.012836f
C484 VTAIL.n169 VSUBS 0.013591f
C485 VTAIL.n170 VSUBS 0.030339f
C486 VTAIL.n171 VSUBS 0.030339f
C487 VTAIL.n172 VSUBS 0.013591f
C488 VTAIL.n173 VSUBS 0.012836f
C489 VTAIL.n174 VSUBS 0.023887f
C490 VTAIL.n175 VSUBS 0.023887f
C491 VTAIL.n176 VSUBS 0.012836f
C492 VTAIL.n177 VSUBS 0.013591f
C493 VTAIL.n178 VSUBS 0.030339f
C494 VTAIL.n179 VSUBS 0.030339f
C495 VTAIL.n180 VSUBS 0.013591f
C496 VTAIL.n181 VSUBS 0.012836f
C497 VTAIL.n182 VSUBS 0.023887f
C498 VTAIL.n183 VSUBS 0.023887f
C499 VTAIL.n184 VSUBS 0.012836f
C500 VTAIL.n185 VSUBS 0.013213f
C501 VTAIL.n186 VSUBS 0.013213f
C502 VTAIL.n187 VSUBS 0.030339f
C503 VTAIL.n188 VSUBS 0.030339f
C504 VTAIL.n189 VSUBS 0.013591f
C505 VTAIL.n190 VSUBS 0.012836f
C506 VTAIL.n191 VSUBS 0.023887f
C507 VTAIL.n192 VSUBS 0.023887f
C508 VTAIL.n193 VSUBS 0.012836f
C509 VTAIL.n194 VSUBS 0.013591f
C510 VTAIL.n195 VSUBS 0.030339f
C511 VTAIL.n196 VSUBS 0.030339f
C512 VTAIL.n197 VSUBS 0.013591f
C513 VTAIL.n198 VSUBS 0.012836f
C514 VTAIL.n199 VSUBS 0.023887f
C515 VTAIL.n200 VSUBS 0.023887f
C516 VTAIL.n201 VSUBS 0.012836f
C517 VTAIL.n202 VSUBS 0.013591f
C518 VTAIL.n203 VSUBS 0.030339f
C519 VTAIL.n204 VSUBS 0.075523f
C520 VTAIL.n205 VSUBS 0.013591f
C521 VTAIL.n206 VSUBS 0.012836f
C522 VTAIL.n207 VSUBS 0.056193f
C523 VTAIL.n208 VSUBS 0.038102f
C524 VTAIL.n209 VSUBS 1.35433f
C525 VTAIL.n210 VSUBS 0.026856f
C526 VTAIL.n211 VSUBS 0.023887f
C527 VTAIL.n212 VSUBS 0.012836f
C528 VTAIL.n213 VSUBS 0.030339f
C529 VTAIL.n214 VSUBS 0.013591f
C530 VTAIL.n215 VSUBS 0.023887f
C531 VTAIL.n216 VSUBS 0.012836f
C532 VTAIL.n217 VSUBS 0.030339f
C533 VTAIL.n218 VSUBS 0.013591f
C534 VTAIL.n219 VSUBS 0.023887f
C535 VTAIL.n220 VSUBS 0.012836f
C536 VTAIL.n221 VSUBS 0.030339f
C537 VTAIL.n222 VSUBS 0.013591f
C538 VTAIL.n223 VSUBS 0.023887f
C539 VTAIL.n224 VSUBS 0.012836f
C540 VTAIL.n225 VSUBS 0.030339f
C541 VTAIL.n226 VSUBS 0.013591f
C542 VTAIL.n227 VSUBS 0.023887f
C543 VTAIL.n228 VSUBS 0.012836f
C544 VTAIL.n229 VSUBS 0.030339f
C545 VTAIL.n230 VSUBS 0.013591f
C546 VTAIL.n231 VSUBS 0.197521f
C547 VTAIL.t3 VSUBS 0.065447f
C548 VTAIL.n232 VSUBS 0.022755f
C549 VTAIL.n233 VSUBS 0.022823f
C550 VTAIL.n234 VSUBS 0.012836f
C551 VTAIL.n235 VSUBS 1.26471f
C552 VTAIL.n236 VSUBS 0.023887f
C553 VTAIL.n237 VSUBS 0.012836f
C554 VTAIL.n238 VSUBS 0.013591f
C555 VTAIL.n239 VSUBS 0.030339f
C556 VTAIL.n240 VSUBS 0.030339f
C557 VTAIL.n241 VSUBS 0.013591f
C558 VTAIL.n242 VSUBS 0.012836f
C559 VTAIL.n243 VSUBS 0.023887f
C560 VTAIL.n244 VSUBS 0.023887f
C561 VTAIL.n245 VSUBS 0.012836f
C562 VTAIL.n246 VSUBS 0.013591f
C563 VTAIL.n247 VSUBS 0.030339f
C564 VTAIL.n248 VSUBS 0.030339f
C565 VTAIL.n249 VSUBS 0.030339f
C566 VTAIL.n250 VSUBS 0.013591f
C567 VTAIL.n251 VSUBS 0.012836f
C568 VTAIL.n252 VSUBS 0.023887f
C569 VTAIL.n253 VSUBS 0.023887f
C570 VTAIL.n254 VSUBS 0.012836f
C571 VTAIL.n255 VSUBS 0.013213f
C572 VTAIL.n256 VSUBS 0.013213f
C573 VTAIL.n257 VSUBS 0.030339f
C574 VTAIL.n258 VSUBS 0.030339f
C575 VTAIL.n259 VSUBS 0.013591f
C576 VTAIL.n260 VSUBS 0.012836f
C577 VTAIL.n261 VSUBS 0.023887f
C578 VTAIL.n262 VSUBS 0.023887f
C579 VTAIL.n263 VSUBS 0.012836f
C580 VTAIL.n264 VSUBS 0.013591f
C581 VTAIL.n265 VSUBS 0.030339f
C582 VTAIL.n266 VSUBS 0.030339f
C583 VTAIL.n267 VSUBS 0.013591f
C584 VTAIL.n268 VSUBS 0.012836f
C585 VTAIL.n269 VSUBS 0.023887f
C586 VTAIL.n270 VSUBS 0.023887f
C587 VTAIL.n271 VSUBS 0.012836f
C588 VTAIL.n272 VSUBS 0.013591f
C589 VTAIL.n273 VSUBS 0.030339f
C590 VTAIL.n274 VSUBS 0.075523f
C591 VTAIL.n275 VSUBS 0.013591f
C592 VTAIL.n276 VSUBS 0.012836f
C593 VTAIL.n277 VSUBS 0.056193f
C594 VTAIL.n278 VSUBS 0.038102f
C595 VTAIL.n279 VSUBS 1.29412f
C596 VN.t0 VSUBS 1.4656f
C597 VN.t1 VSUBS 1.60365f
C598 B.n0 VSUBS 0.004541f
C599 B.n1 VSUBS 0.004541f
C600 B.n2 VSUBS 0.007181f
C601 B.n3 VSUBS 0.007181f
C602 B.n4 VSUBS 0.007181f
C603 B.n5 VSUBS 0.007181f
C604 B.n6 VSUBS 0.007181f
C605 B.n7 VSUBS 0.007181f
C606 B.n8 VSUBS 0.007181f
C607 B.n9 VSUBS 0.016584f
C608 B.n10 VSUBS 0.007181f
C609 B.n11 VSUBS 0.007181f
C610 B.n12 VSUBS 0.007181f
C611 B.n13 VSUBS 0.007181f
C612 B.n14 VSUBS 0.007181f
C613 B.n15 VSUBS 0.007181f
C614 B.n16 VSUBS 0.007181f
C615 B.n17 VSUBS 0.007181f
C616 B.n18 VSUBS 0.007181f
C617 B.n19 VSUBS 0.007181f
C618 B.n20 VSUBS 0.007181f
C619 B.n21 VSUBS 0.007181f
C620 B.n22 VSUBS 0.007181f
C621 B.n23 VSUBS 0.007181f
C622 B.n24 VSUBS 0.007181f
C623 B.n25 VSUBS 0.007181f
C624 B.n26 VSUBS 0.007181f
C625 B.n27 VSUBS 0.007181f
C626 B.n28 VSUBS 0.007181f
C627 B.n29 VSUBS 0.007181f
C628 B.n30 VSUBS 0.007181f
C629 B.n31 VSUBS 0.007181f
C630 B.t5 VSUBS 0.236692f
C631 B.t4 VSUBS 0.250649f
C632 B.t3 VSUBS 0.467207f
C633 B.n32 VSUBS 0.350671f
C634 B.n33 VSUBS 0.262937f
C635 B.n34 VSUBS 0.007181f
C636 B.n35 VSUBS 0.007181f
C637 B.n36 VSUBS 0.007181f
C638 B.n37 VSUBS 0.007181f
C639 B.n38 VSUBS 0.004224f
C640 B.n39 VSUBS 0.007181f
C641 B.t11 VSUBS 0.236696f
C642 B.t10 VSUBS 0.250652f
C643 B.t9 VSUBS 0.467207f
C644 B.n40 VSUBS 0.350668f
C645 B.n41 VSUBS 0.262933f
C646 B.n42 VSUBS 0.016637f
C647 B.n43 VSUBS 0.007181f
C648 B.n44 VSUBS 0.007181f
C649 B.n45 VSUBS 0.007181f
C650 B.n46 VSUBS 0.007181f
C651 B.n47 VSUBS 0.007181f
C652 B.n48 VSUBS 0.007181f
C653 B.n49 VSUBS 0.007181f
C654 B.n50 VSUBS 0.007181f
C655 B.n51 VSUBS 0.007181f
C656 B.n52 VSUBS 0.007181f
C657 B.n53 VSUBS 0.007181f
C658 B.n54 VSUBS 0.007181f
C659 B.n55 VSUBS 0.007181f
C660 B.n56 VSUBS 0.007181f
C661 B.n57 VSUBS 0.007181f
C662 B.n58 VSUBS 0.007181f
C663 B.n59 VSUBS 0.007181f
C664 B.n60 VSUBS 0.007181f
C665 B.n61 VSUBS 0.007181f
C666 B.n62 VSUBS 0.007181f
C667 B.n63 VSUBS 0.016584f
C668 B.n64 VSUBS 0.007181f
C669 B.n65 VSUBS 0.007181f
C670 B.n66 VSUBS 0.007181f
C671 B.n67 VSUBS 0.007181f
C672 B.n68 VSUBS 0.007181f
C673 B.n69 VSUBS 0.007181f
C674 B.n70 VSUBS 0.007181f
C675 B.n71 VSUBS 0.007181f
C676 B.n72 VSUBS 0.007181f
C677 B.n73 VSUBS 0.007181f
C678 B.n74 VSUBS 0.007181f
C679 B.n75 VSUBS 0.007181f
C680 B.n76 VSUBS 0.007181f
C681 B.n77 VSUBS 0.007181f
C682 B.n78 VSUBS 0.007181f
C683 B.n79 VSUBS 0.017418f
C684 B.n80 VSUBS 0.007181f
C685 B.n81 VSUBS 0.007181f
C686 B.n82 VSUBS 0.007181f
C687 B.n83 VSUBS 0.007181f
C688 B.n84 VSUBS 0.007181f
C689 B.n85 VSUBS 0.007181f
C690 B.n86 VSUBS 0.007181f
C691 B.n87 VSUBS 0.007181f
C692 B.n88 VSUBS 0.007181f
C693 B.n89 VSUBS 0.007181f
C694 B.n90 VSUBS 0.007181f
C695 B.n91 VSUBS 0.007181f
C696 B.n92 VSUBS 0.007181f
C697 B.n93 VSUBS 0.007181f
C698 B.n94 VSUBS 0.007181f
C699 B.n95 VSUBS 0.007181f
C700 B.n96 VSUBS 0.007181f
C701 B.n97 VSUBS 0.007181f
C702 B.n98 VSUBS 0.007181f
C703 B.n99 VSUBS 0.007181f
C704 B.n100 VSUBS 0.007181f
C705 B.t1 VSUBS 0.236696f
C706 B.t2 VSUBS 0.250652f
C707 B.t0 VSUBS 0.467207f
C708 B.n101 VSUBS 0.350668f
C709 B.n102 VSUBS 0.262933f
C710 B.n103 VSUBS 0.016637f
C711 B.n104 VSUBS 0.007181f
C712 B.n105 VSUBS 0.007181f
C713 B.n106 VSUBS 0.007181f
C714 B.n107 VSUBS 0.007181f
C715 B.n108 VSUBS 0.007181f
C716 B.t7 VSUBS 0.236692f
C717 B.t8 VSUBS 0.250649f
C718 B.t6 VSUBS 0.467207f
C719 B.n109 VSUBS 0.350671f
C720 B.n110 VSUBS 0.262937f
C721 B.n111 VSUBS 0.007181f
C722 B.n112 VSUBS 0.007181f
C723 B.n113 VSUBS 0.007181f
C724 B.n114 VSUBS 0.007181f
C725 B.n115 VSUBS 0.007181f
C726 B.n116 VSUBS 0.007181f
C727 B.n117 VSUBS 0.007181f
C728 B.n118 VSUBS 0.007181f
C729 B.n119 VSUBS 0.007181f
C730 B.n120 VSUBS 0.007181f
C731 B.n121 VSUBS 0.007181f
C732 B.n122 VSUBS 0.007181f
C733 B.n123 VSUBS 0.007181f
C734 B.n124 VSUBS 0.007181f
C735 B.n125 VSUBS 0.007181f
C736 B.n126 VSUBS 0.007181f
C737 B.n127 VSUBS 0.007181f
C738 B.n128 VSUBS 0.007181f
C739 B.n129 VSUBS 0.007181f
C740 B.n130 VSUBS 0.007181f
C741 B.n131 VSUBS 0.007181f
C742 B.n132 VSUBS 0.017418f
C743 B.n133 VSUBS 0.007181f
C744 B.n134 VSUBS 0.007181f
C745 B.n135 VSUBS 0.007181f
C746 B.n136 VSUBS 0.007181f
C747 B.n137 VSUBS 0.007181f
C748 B.n138 VSUBS 0.007181f
C749 B.n139 VSUBS 0.007181f
C750 B.n140 VSUBS 0.007181f
C751 B.n141 VSUBS 0.007181f
C752 B.n142 VSUBS 0.007181f
C753 B.n143 VSUBS 0.007181f
C754 B.n144 VSUBS 0.007181f
C755 B.n145 VSUBS 0.007181f
C756 B.n146 VSUBS 0.007181f
C757 B.n147 VSUBS 0.007181f
C758 B.n148 VSUBS 0.007181f
C759 B.n149 VSUBS 0.007181f
C760 B.n150 VSUBS 0.007181f
C761 B.n151 VSUBS 0.007181f
C762 B.n152 VSUBS 0.007181f
C763 B.n153 VSUBS 0.007181f
C764 B.n154 VSUBS 0.007181f
C765 B.n155 VSUBS 0.007181f
C766 B.n156 VSUBS 0.007181f
C767 B.n157 VSUBS 0.007181f
C768 B.n158 VSUBS 0.007181f
C769 B.n159 VSUBS 0.016584f
C770 B.n160 VSUBS 0.016584f
C771 B.n161 VSUBS 0.017418f
C772 B.n162 VSUBS 0.007181f
C773 B.n163 VSUBS 0.007181f
C774 B.n164 VSUBS 0.007181f
C775 B.n165 VSUBS 0.007181f
C776 B.n166 VSUBS 0.007181f
C777 B.n167 VSUBS 0.007181f
C778 B.n168 VSUBS 0.007181f
C779 B.n169 VSUBS 0.007181f
C780 B.n170 VSUBS 0.007181f
C781 B.n171 VSUBS 0.007181f
C782 B.n172 VSUBS 0.007181f
C783 B.n173 VSUBS 0.007181f
C784 B.n174 VSUBS 0.007181f
C785 B.n175 VSUBS 0.007181f
C786 B.n176 VSUBS 0.007181f
C787 B.n177 VSUBS 0.007181f
C788 B.n178 VSUBS 0.007181f
C789 B.n179 VSUBS 0.007181f
C790 B.n180 VSUBS 0.007181f
C791 B.n181 VSUBS 0.007181f
C792 B.n182 VSUBS 0.007181f
C793 B.n183 VSUBS 0.007181f
C794 B.n184 VSUBS 0.007181f
C795 B.n185 VSUBS 0.007181f
C796 B.n186 VSUBS 0.007181f
C797 B.n187 VSUBS 0.007181f
C798 B.n188 VSUBS 0.007181f
C799 B.n189 VSUBS 0.007181f
C800 B.n190 VSUBS 0.007181f
C801 B.n191 VSUBS 0.007181f
C802 B.n192 VSUBS 0.007181f
C803 B.n193 VSUBS 0.007181f
C804 B.n194 VSUBS 0.007181f
C805 B.n195 VSUBS 0.007181f
C806 B.n196 VSUBS 0.007181f
C807 B.n197 VSUBS 0.007181f
C808 B.n198 VSUBS 0.007181f
C809 B.n199 VSUBS 0.007181f
C810 B.n200 VSUBS 0.007181f
C811 B.n201 VSUBS 0.007181f
C812 B.n202 VSUBS 0.007181f
C813 B.n203 VSUBS 0.007181f
C814 B.n204 VSUBS 0.007181f
C815 B.n205 VSUBS 0.007181f
C816 B.n206 VSUBS 0.007181f
C817 B.n207 VSUBS 0.007181f
C818 B.n208 VSUBS 0.007181f
C819 B.n209 VSUBS 0.007181f
C820 B.n210 VSUBS 0.007181f
C821 B.n211 VSUBS 0.007181f
C822 B.n212 VSUBS 0.007181f
C823 B.n213 VSUBS 0.007181f
C824 B.n214 VSUBS 0.007181f
C825 B.n215 VSUBS 0.007181f
C826 B.n216 VSUBS 0.007181f
C827 B.n217 VSUBS 0.007181f
C828 B.n218 VSUBS 0.007181f
C829 B.n219 VSUBS 0.007181f
C830 B.n220 VSUBS 0.007181f
C831 B.n221 VSUBS 0.007181f
C832 B.n222 VSUBS 0.007181f
C833 B.n223 VSUBS 0.007181f
C834 B.n224 VSUBS 0.007181f
C835 B.n225 VSUBS 0.007181f
C836 B.n226 VSUBS 0.006547f
C837 B.n227 VSUBS 0.016637f
C838 B.n228 VSUBS 0.004224f
C839 B.n229 VSUBS 0.007181f
C840 B.n230 VSUBS 0.007181f
C841 B.n231 VSUBS 0.007181f
C842 B.n232 VSUBS 0.007181f
C843 B.n233 VSUBS 0.007181f
C844 B.n234 VSUBS 0.007181f
C845 B.n235 VSUBS 0.007181f
C846 B.n236 VSUBS 0.007181f
C847 B.n237 VSUBS 0.007181f
C848 B.n238 VSUBS 0.007181f
C849 B.n239 VSUBS 0.007181f
C850 B.n240 VSUBS 0.007181f
C851 B.n241 VSUBS 0.004224f
C852 B.n242 VSUBS 0.007181f
C853 B.n243 VSUBS 0.007181f
C854 B.n244 VSUBS 0.006547f
C855 B.n245 VSUBS 0.007181f
C856 B.n246 VSUBS 0.007181f
C857 B.n247 VSUBS 0.007181f
C858 B.n248 VSUBS 0.007181f
C859 B.n249 VSUBS 0.007181f
C860 B.n250 VSUBS 0.007181f
C861 B.n251 VSUBS 0.007181f
C862 B.n252 VSUBS 0.007181f
C863 B.n253 VSUBS 0.007181f
C864 B.n254 VSUBS 0.007181f
C865 B.n255 VSUBS 0.007181f
C866 B.n256 VSUBS 0.007181f
C867 B.n257 VSUBS 0.007181f
C868 B.n258 VSUBS 0.007181f
C869 B.n259 VSUBS 0.007181f
C870 B.n260 VSUBS 0.007181f
C871 B.n261 VSUBS 0.007181f
C872 B.n262 VSUBS 0.007181f
C873 B.n263 VSUBS 0.007181f
C874 B.n264 VSUBS 0.007181f
C875 B.n265 VSUBS 0.007181f
C876 B.n266 VSUBS 0.007181f
C877 B.n267 VSUBS 0.007181f
C878 B.n268 VSUBS 0.007181f
C879 B.n269 VSUBS 0.007181f
C880 B.n270 VSUBS 0.007181f
C881 B.n271 VSUBS 0.007181f
C882 B.n272 VSUBS 0.007181f
C883 B.n273 VSUBS 0.007181f
C884 B.n274 VSUBS 0.007181f
C885 B.n275 VSUBS 0.007181f
C886 B.n276 VSUBS 0.007181f
C887 B.n277 VSUBS 0.007181f
C888 B.n278 VSUBS 0.007181f
C889 B.n279 VSUBS 0.007181f
C890 B.n280 VSUBS 0.007181f
C891 B.n281 VSUBS 0.007181f
C892 B.n282 VSUBS 0.007181f
C893 B.n283 VSUBS 0.007181f
C894 B.n284 VSUBS 0.007181f
C895 B.n285 VSUBS 0.007181f
C896 B.n286 VSUBS 0.007181f
C897 B.n287 VSUBS 0.007181f
C898 B.n288 VSUBS 0.007181f
C899 B.n289 VSUBS 0.007181f
C900 B.n290 VSUBS 0.007181f
C901 B.n291 VSUBS 0.007181f
C902 B.n292 VSUBS 0.007181f
C903 B.n293 VSUBS 0.007181f
C904 B.n294 VSUBS 0.007181f
C905 B.n295 VSUBS 0.007181f
C906 B.n296 VSUBS 0.007181f
C907 B.n297 VSUBS 0.007181f
C908 B.n298 VSUBS 0.007181f
C909 B.n299 VSUBS 0.007181f
C910 B.n300 VSUBS 0.007181f
C911 B.n301 VSUBS 0.007181f
C912 B.n302 VSUBS 0.007181f
C913 B.n303 VSUBS 0.007181f
C914 B.n304 VSUBS 0.007181f
C915 B.n305 VSUBS 0.007181f
C916 B.n306 VSUBS 0.007181f
C917 B.n307 VSUBS 0.007181f
C918 B.n308 VSUBS 0.017418f
C919 B.n309 VSUBS 0.016584f
C920 B.n310 VSUBS 0.016584f
C921 B.n311 VSUBS 0.007181f
C922 B.n312 VSUBS 0.007181f
C923 B.n313 VSUBS 0.007181f
C924 B.n314 VSUBS 0.007181f
C925 B.n315 VSUBS 0.007181f
C926 B.n316 VSUBS 0.007181f
C927 B.n317 VSUBS 0.007181f
C928 B.n318 VSUBS 0.007181f
C929 B.n319 VSUBS 0.007181f
C930 B.n320 VSUBS 0.007181f
C931 B.n321 VSUBS 0.007181f
C932 B.n322 VSUBS 0.007181f
C933 B.n323 VSUBS 0.007181f
C934 B.n324 VSUBS 0.007181f
C935 B.n325 VSUBS 0.007181f
C936 B.n326 VSUBS 0.007181f
C937 B.n327 VSUBS 0.007181f
C938 B.n328 VSUBS 0.007181f
C939 B.n329 VSUBS 0.007181f
C940 B.n330 VSUBS 0.007181f
C941 B.n331 VSUBS 0.007181f
C942 B.n332 VSUBS 0.007181f
C943 B.n333 VSUBS 0.007181f
C944 B.n334 VSUBS 0.007181f
C945 B.n335 VSUBS 0.007181f
C946 B.n336 VSUBS 0.007181f
C947 B.n337 VSUBS 0.007181f
C948 B.n338 VSUBS 0.007181f
C949 B.n339 VSUBS 0.007181f
C950 B.n340 VSUBS 0.007181f
C951 B.n341 VSUBS 0.007181f
C952 B.n342 VSUBS 0.007181f
C953 B.n343 VSUBS 0.007181f
C954 B.n344 VSUBS 0.007181f
C955 B.n345 VSUBS 0.007181f
C956 B.n346 VSUBS 0.007181f
C957 B.n347 VSUBS 0.007181f
C958 B.n348 VSUBS 0.007181f
C959 B.n349 VSUBS 0.007181f
C960 B.n350 VSUBS 0.007181f
C961 B.n351 VSUBS 0.007181f
C962 B.n352 VSUBS 0.007181f
C963 B.n353 VSUBS 0.007181f
C964 B.n354 VSUBS 0.017418f
C965 B.n355 VSUBS 0.016584f
C966 B.n356 VSUBS 0.017418f
C967 B.n357 VSUBS 0.007181f
C968 B.n358 VSUBS 0.007181f
C969 B.n359 VSUBS 0.007181f
C970 B.n360 VSUBS 0.007181f
C971 B.n361 VSUBS 0.007181f
C972 B.n362 VSUBS 0.007181f
C973 B.n363 VSUBS 0.007181f
C974 B.n364 VSUBS 0.007181f
C975 B.n365 VSUBS 0.007181f
C976 B.n366 VSUBS 0.007181f
C977 B.n367 VSUBS 0.007181f
C978 B.n368 VSUBS 0.007181f
C979 B.n369 VSUBS 0.007181f
C980 B.n370 VSUBS 0.007181f
C981 B.n371 VSUBS 0.007181f
C982 B.n372 VSUBS 0.007181f
C983 B.n373 VSUBS 0.007181f
C984 B.n374 VSUBS 0.007181f
C985 B.n375 VSUBS 0.007181f
C986 B.n376 VSUBS 0.007181f
C987 B.n377 VSUBS 0.007181f
C988 B.n378 VSUBS 0.007181f
C989 B.n379 VSUBS 0.007181f
C990 B.n380 VSUBS 0.007181f
C991 B.n381 VSUBS 0.007181f
C992 B.n382 VSUBS 0.007181f
C993 B.n383 VSUBS 0.007181f
C994 B.n384 VSUBS 0.007181f
C995 B.n385 VSUBS 0.007181f
C996 B.n386 VSUBS 0.007181f
C997 B.n387 VSUBS 0.007181f
C998 B.n388 VSUBS 0.007181f
C999 B.n389 VSUBS 0.007181f
C1000 B.n390 VSUBS 0.007181f
C1001 B.n391 VSUBS 0.007181f
C1002 B.n392 VSUBS 0.007181f
C1003 B.n393 VSUBS 0.007181f
C1004 B.n394 VSUBS 0.007181f
C1005 B.n395 VSUBS 0.007181f
C1006 B.n396 VSUBS 0.007181f
C1007 B.n397 VSUBS 0.007181f
C1008 B.n398 VSUBS 0.007181f
C1009 B.n399 VSUBS 0.007181f
C1010 B.n400 VSUBS 0.007181f
C1011 B.n401 VSUBS 0.007181f
C1012 B.n402 VSUBS 0.007181f
C1013 B.n403 VSUBS 0.007181f
C1014 B.n404 VSUBS 0.007181f
C1015 B.n405 VSUBS 0.007181f
C1016 B.n406 VSUBS 0.007181f
C1017 B.n407 VSUBS 0.007181f
C1018 B.n408 VSUBS 0.007181f
C1019 B.n409 VSUBS 0.007181f
C1020 B.n410 VSUBS 0.007181f
C1021 B.n411 VSUBS 0.007181f
C1022 B.n412 VSUBS 0.007181f
C1023 B.n413 VSUBS 0.007181f
C1024 B.n414 VSUBS 0.007181f
C1025 B.n415 VSUBS 0.007181f
C1026 B.n416 VSUBS 0.007181f
C1027 B.n417 VSUBS 0.007181f
C1028 B.n418 VSUBS 0.007181f
C1029 B.n419 VSUBS 0.007181f
C1030 B.n420 VSUBS 0.006547f
C1031 B.n421 VSUBS 0.007181f
C1032 B.n422 VSUBS 0.007181f
C1033 B.n423 VSUBS 0.007181f
C1034 B.n424 VSUBS 0.007181f
C1035 B.n425 VSUBS 0.007181f
C1036 B.n426 VSUBS 0.007181f
C1037 B.n427 VSUBS 0.007181f
C1038 B.n428 VSUBS 0.007181f
C1039 B.n429 VSUBS 0.007181f
C1040 B.n430 VSUBS 0.007181f
C1041 B.n431 VSUBS 0.007181f
C1042 B.n432 VSUBS 0.007181f
C1043 B.n433 VSUBS 0.007181f
C1044 B.n434 VSUBS 0.007181f
C1045 B.n435 VSUBS 0.007181f
C1046 B.n436 VSUBS 0.004224f
C1047 B.n437 VSUBS 0.016637f
C1048 B.n438 VSUBS 0.006547f
C1049 B.n439 VSUBS 0.007181f
C1050 B.n440 VSUBS 0.007181f
C1051 B.n441 VSUBS 0.007181f
C1052 B.n442 VSUBS 0.007181f
C1053 B.n443 VSUBS 0.007181f
C1054 B.n444 VSUBS 0.007181f
C1055 B.n445 VSUBS 0.007181f
C1056 B.n446 VSUBS 0.007181f
C1057 B.n447 VSUBS 0.007181f
C1058 B.n448 VSUBS 0.007181f
C1059 B.n449 VSUBS 0.007181f
C1060 B.n450 VSUBS 0.007181f
C1061 B.n451 VSUBS 0.007181f
C1062 B.n452 VSUBS 0.007181f
C1063 B.n453 VSUBS 0.007181f
C1064 B.n454 VSUBS 0.007181f
C1065 B.n455 VSUBS 0.007181f
C1066 B.n456 VSUBS 0.007181f
C1067 B.n457 VSUBS 0.007181f
C1068 B.n458 VSUBS 0.007181f
C1069 B.n459 VSUBS 0.007181f
C1070 B.n460 VSUBS 0.007181f
C1071 B.n461 VSUBS 0.007181f
C1072 B.n462 VSUBS 0.007181f
C1073 B.n463 VSUBS 0.007181f
C1074 B.n464 VSUBS 0.007181f
C1075 B.n465 VSUBS 0.007181f
C1076 B.n466 VSUBS 0.007181f
C1077 B.n467 VSUBS 0.007181f
C1078 B.n468 VSUBS 0.007181f
C1079 B.n469 VSUBS 0.007181f
C1080 B.n470 VSUBS 0.007181f
C1081 B.n471 VSUBS 0.007181f
C1082 B.n472 VSUBS 0.007181f
C1083 B.n473 VSUBS 0.007181f
C1084 B.n474 VSUBS 0.007181f
C1085 B.n475 VSUBS 0.007181f
C1086 B.n476 VSUBS 0.007181f
C1087 B.n477 VSUBS 0.007181f
C1088 B.n478 VSUBS 0.007181f
C1089 B.n479 VSUBS 0.007181f
C1090 B.n480 VSUBS 0.007181f
C1091 B.n481 VSUBS 0.007181f
C1092 B.n482 VSUBS 0.007181f
C1093 B.n483 VSUBS 0.007181f
C1094 B.n484 VSUBS 0.007181f
C1095 B.n485 VSUBS 0.007181f
C1096 B.n486 VSUBS 0.007181f
C1097 B.n487 VSUBS 0.007181f
C1098 B.n488 VSUBS 0.007181f
C1099 B.n489 VSUBS 0.007181f
C1100 B.n490 VSUBS 0.007181f
C1101 B.n491 VSUBS 0.007181f
C1102 B.n492 VSUBS 0.007181f
C1103 B.n493 VSUBS 0.007181f
C1104 B.n494 VSUBS 0.007181f
C1105 B.n495 VSUBS 0.007181f
C1106 B.n496 VSUBS 0.007181f
C1107 B.n497 VSUBS 0.007181f
C1108 B.n498 VSUBS 0.007181f
C1109 B.n499 VSUBS 0.007181f
C1110 B.n500 VSUBS 0.007181f
C1111 B.n501 VSUBS 0.007181f
C1112 B.n502 VSUBS 0.017418f
C1113 B.n503 VSUBS 0.017418f
C1114 B.n504 VSUBS 0.016584f
C1115 B.n505 VSUBS 0.007181f
C1116 B.n506 VSUBS 0.007181f
C1117 B.n507 VSUBS 0.007181f
C1118 B.n508 VSUBS 0.007181f
C1119 B.n509 VSUBS 0.007181f
C1120 B.n510 VSUBS 0.007181f
C1121 B.n511 VSUBS 0.007181f
C1122 B.n512 VSUBS 0.007181f
C1123 B.n513 VSUBS 0.007181f
C1124 B.n514 VSUBS 0.007181f
C1125 B.n515 VSUBS 0.007181f
C1126 B.n516 VSUBS 0.007181f
C1127 B.n517 VSUBS 0.007181f
C1128 B.n518 VSUBS 0.007181f
C1129 B.n519 VSUBS 0.007181f
C1130 B.n520 VSUBS 0.007181f
C1131 B.n521 VSUBS 0.007181f
C1132 B.n522 VSUBS 0.007181f
C1133 B.n523 VSUBS 0.007181f
C1134 B.n524 VSUBS 0.007181f
C1135 B.n525 VSUBS 0.007181f
C1136 B.n526 VSUBS 0.007181f
C1137 B.n527 VSUBS 0.016259f
.ends

