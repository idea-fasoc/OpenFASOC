* NGSPICE file created from diff_pair_sample_0067.ext - technology: sky130A

.subckt diff_pair_sample_0067 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t14 w_n1850_n3600# sky130_fd_pr__pfet_01v8 ad=2.1714 pd=13.49 as=2.1714 ps=13.49 w=13.16 l=0.55
X1 VTAIL.t13 VP.t1 VDD1.t6 w_n1850_n3600# sky130_fd_pr__pfet_01v8 ad=5.1324 pd=27.1 as=2.1714 ps=13.49 w=13.16 l=0.55
X2 VDD1.t5 VP.t2 VTAIL.t8 w_n1850_n3600# sky130_fd_pr__pfet_01v8 ad=2.1714 pd=13.49 as=5.1324 ps=27.1 w=13.16 l=0.55
X3 VTAIL.t11 VP.t3 VDD1.t4 w_n1850_n3600# sky130_fd_pr__pfet_01v8 ad=2.1714 pd=13.49 as=2.1714 ps=13.49 w=13.16 l=0.55
X4 VDD2.t7 VN.t0 VTAIL.t4 w_n1850_n3600# sky130_fd_pr__pfet_01v8 ad=2.1714 pd=13.49 as=5.1324 ps=27.1 w=13.16 l=0.55
X5 VDD2.t6 VN.t1 VTAIL.t7 w_n1850_n3600# sky130_fd_pr__pfet_01v8 ad=2.1714 pd=13.49 as=2.1714 ps=13.49 w=13.16 l=0.55
X6 VTAIL.t12 VP.t4 VDD1.t3 w_n1850_n3600# sky130_fd_pr__pfet_01v8 ad=2.1714 pd=13.49 as=2.1714 ps=13.49 w=13.16 l=0.55
X7 VDD2.t5 VN.t2 VTAIL.t1 w_n1850_n3600# sky130_fd_pr__pfet_01v8 ad=2.1714 pd=13.49 as=5.1324 ps=27.1 w=13.16 l=0.55
X8 VDD1.t2 VP.t5 VTAIL.t9 w_n1850_n3600# sky130_fd_pr__pfet_01v8 ad=2.1714 pd=13.49 as=2.1714 ps=13.49 w=13.16 l=0.55
X9 B.t11 B.t9 B.t10 w_n1850_n3600# sky130_fd_pr__pfet_01v8 ad=5.1324 pd=27.1 as=0 ps=0 w=13.16 l=0.55
X10 VTAIL.t0 VN.t3 VDD2.t4 w_n1850_n3600# sky130_fd_pr__pfet_01v8 ad=5.1324 pd=27.1 as=2.1714 ps=13.49 w=13.16 l=0.55
X11 VDD2.t3 VN.t4 VTAIL.t2 w_n1850_n3600# sky130_fd_pr__pfet_01v8 ad=2.1714 pd=13.49 as=2.1714 ps=13.49 w=13.16 l=0.55
X12 VDD1.t1 VP.t6 VTAIL.t15 w_n1850_n3600# sky130_fd_pr__pfet_01v8 ad=2.1714 pd=13.49 as=5.1324 ps=27.1 w=13.16 l=0.55
X13 B.t8 B.t6 B.t7 w_n1850_n3600# sky130_fd_pr__pfet_01v8 ad=5.1324 pd=27.1 as=0 ps=0 w=13.16 l=0.55
X14 VTAIL.t3 VN.t5 VDD2.t2 w_n1850_n3600# sky130_fd_pr__pfet_01v8 ad=2.1714 pd=13.49 as=2.1714 ps=13.49 w=13.16 l=0.55
X15 B.t5 B.t3 B.t4 w_n1850_n3600# sky130_fd_pr__pfet_01v8 ad=5.1324 pd=27.1 as=0 ps=0 w=13.16 l=0.55
X16 VTAIL.t10 VP.t7 VDD1.t0 w_n1850_n3600# sky130_fd_pr__pfet_01v8 ad=5.1324 pd=27.1 as=2.1714 ps=13.49 w=13.16 l=0.55
X17 VTAIL.t5 VN.t6 VDD2.t1 w_n1850_n3600# sky130_fd_pr__pfet_01v8 ad=5.1324 pd=27.1 as=2.1714 ps=13.49 w=13.16 l=0.55
X18 VTAIL.t6 VN.t7 VDD2.t0 w_n1850_n3600# sky130_fd_pr__pfet_01v8 ad=2.1714 pd=13.49 as=2.1714 ps=13.49 w=13.16 l=0.55
X19 B.t2 B.t0 B.t1 w_n1850_n3600# sky130_fd_pr__pfet_01v8 ad=5.1324 pd=27.1 as=0 ps=0 w=13.16 l=0.55
R0 VP.n4 VP.t7 673.793
R1 VP.n11 VP.t1 648.072
R2 VP.n1 VP.t5 648.072
R3 VP.n16 VP.t4 648.072
R4 VP.n18 VP.t6 648.072
R5 VP.n8 VP.t2 648.072
R6 VP.n6 VP.t3 648.072
R7 VP.n5 VP.t0 648.072
R8 VP.n19 VP.n18 161.3
R9 VP.n6 VP.n3 161.3
R10 VP.n7 VP.n2 161.3
R11 VP.n9 VP.n8 161.3
R12 VP.n17 VP.n0 161.3
R13 VP.n16 VP.n15 161.3
R14 VP.n14 VP.n1 161.3
R15 VP.n13 VP.n12 161.3
R16 VP.n11 VP.n10 161.3
R17 VP.n16 VP.n1 48.2005
R18 VP.n6 VP.n5 48.2005
R19 VP.n4 VP.n3 45.029
R20 VP.n12 VP.n11 43.0884
R21 VP.n18 VP.n17 43.0884
R22 VP.n8 VP.n7 43.0884
R23 VP.n10 VP.n9 42.152
R24 VP.n5 VP.n4 15.1442
R25 VP.n12 VP.n1 5.11262
R26 VP.n17 VP.n16 5.11262
R27 VP.n7 VP.n6 5.11262
R28 VP.n3 VP.n2 0.189894
R29 VP.n9 VP.n2 0.189894
R30 VP.n13 VP.n10 0.189894
R31 VP.n14 VP.n13 0.189894
R32 VP.n15 VP.n14 0.189894
R33 VP.n15 VP.n0 0.189894
R34 VP.n19 VP.n0 0.189894
R35 VP VP.n19 0.0516364
R36 VTAIL.n11 VTAIL.t10 57.6501
R37 VTAIL.n10 VTAIL.t1 57.6501
R38 VTAIL.n7 VTAIL.t5 57.6501
R39 VTAIL.n15 VTAIL.t4 57.6499
R40 VTAIL.n2 VTAIL.t0 57.6499
R41 VTAIL.n3 VTAIL.t15 57.6499
R42 VTAIL.n6 VTAIL.t13 57.6499
R43 VTAIL.n14 VTAIL.t8 57.6499
R44 VTAIL.n13 VTAIL.n12 55.1801
R45 VTAIL.n9 VTAIL.n8 55.1801
R46 VTAIL.n1 VTAIL.n0 55.1801
R47 VTAIL.n5 VTAIL.n4 55.1801
R48 VTAIL.n15 VTAIL.n14 24.4703
R49 VTAIL.n7 VTAIL.n6 24.4703
R50 VTAIL.n0 VTAIL.t7 2.47048
R51 VTAIL.n0 VTAIL.t6 2.47048
R52 VTAIL.n4 VTAIL.t9 2.47048
R53 VTAIL.n4 VTAIL.t12 2.47048
R54 VTAIL.n12 VTAIL.t14 2.47048
R55 VTAIL.n12 VTAIL.t11 2.47048
R56 VTAIL.n8 VTAIL.t2 2.47048
R57 VTAIL.n8 VTAIL.t3 2.47048
R58 VTAIL.n9 VTAIL.n7 0.759121
R59 VTAIL.n10 VTAIL.n9 0.759121
R60 VTAIL.n13 VTAIL.n11 0.759121
R61 VTAIL.n14 VTAIL.n13 0.759121
R62 VTAIL.n6 VTAIL.n5 0.759121
R63 VTAIL.n5 VTAIL.n3 0.759121
R64 VTAIL.n2 VTAIL.n1 0.759121
R65 VTAIL VTAIL.n15 0.700931
R66 VTAIL.n11 VTAIL.n10 0.470328
R67 VTAIL.n3 VTAIL.n2 0.470328
R68 VTAIL VTAIL.n1 0.0586897
R69 VDD1 VDD1.n0 72.2964
R70 VDD1.n3 VDD1.n2 72.1828
R71 VDD1.n3 VDD1.n1 72.1828
R72 VDD1.n5 VDD1.n4 71.8587
R73 VDD1.n5 VDD1.n3 39.0569
R74 VDD1.n4 VDD1.t4 2.47048
R75 VDD1.n4 VDD1.t5 2.47048
R76 VDD1.n0 VDD1.t0 2.47048
R77 VDD1.n0 VDD1.t7 2.47048
R78 VDD1.n2 VDD1.t3 2.47048
R79 VDD1.n2 VDD1.t1 2.47048
R80 VDD1.n1 VDD1.t6 2.47048
R81 VDD1.n1 VDD1.t2 2.47048
R82 VDD1 VDD1.n5 0.321621
R83 VN.n2 VN.t3 673.793
R84 VN.n10 VN.t2 673.793
R85 VN.n1 VN.t1 648.072
R86 VN.n4 VN.t7 648.072
R87 VN.n6 VN.t0 648.072
R88 VN.n9 VN.t5 648.072
R89 VN.n12 VN.t4 648.072
R90 VN.n14 VN.t6 648.072
R91 VN.n7 VN.n6 161.3
R92 VN.n15 VN.n14 161.3
R93 VN.n13 VN.n8 161.3
R94 VN.n12 VN.n11 161.3
R95 VN.n5 VN.n0 161.3
R96 VN.n4 VN.n3 161.3
R97 VN.n4 VN.n1 48.2005
R98 VN.n12 VN.n9 48.2005
R99 VN.n11 VN.n10 45.029
R100 VN.n3 VN.n2 45.029
R101 VN.n6 VN.n5 43.0884
R102 VN.n14 VN.n13 43.0884
R103 VN VN.n15 42.5327
R104 VN.n2 VN.n1 15.1442
R105 VN.n10 VN.n9 15.1442
R106 VN.n5 VN.n4 5.11262
R107 VN.n13 VN.n12 5.11262
R108 VN.n15 VN.n8 0.189894
R109 VN.n11 VN.n8 0.189894
R110 VN.n3 VN.n0 0.189894
R111 VN.n7 VN.n0 0.189894
R112 VN VN.n7 0.0516364
R113 VDD2.n2 VDD2.n1 72.1828
R114 VDD2.n2 VDD2.n0 72.1828
R115 VDD2 VDD2.n5 72.1799
R116 VDD2.n4 VDD2.n3 71.8589
R117 VDD2.n4 VDD2.n2 38.4739
R118 VDD2.n5 VDD2.t2 2.47048
R119 VDD2.n5 VDD2.t5 2.47048
R120 VDD2.n3 VDD2.t1 2.47048
R121 VDD2.n3 VDD2.t3 2.47048
R122 VDD2.n1 VDD2.t0 2.47048
R123 VDD2.n1 VDD2.t7 2.47048
R124 VDD2.n0 VDD2.t4 2.47048
R125 VDD2.n0 VDD2.t6 2.47048
R126 VDD2 VDD2.n4 0.438
R127 B.n112 B.t9 781.96
R128 B.n118 B.t3 781.96
R129 B.n36 B.t0 781.96
R130 B.n42 B.t6 781.96
R131 B.n400 B.n399 585
R132 B.n401 B.n66 585
R133 B.n403 B.n402 585
R134 B.n404 B.n65 585
R135 B.n406 B.n405 585
R136 B.n407 B.n64 585
R137 B.n409 B.n408 585
R138 B.n410 B.n63 585
R139 B.n412 B.n411 585
R140 B.n413 B.n62 585
R141 B.n415 B.n414 585
R142 B.n416 B.n61 585
R143 B.n418 B.n417 585
R144 B.n419 B.n60 585
R145 B.n421 B.n420 585
R146 B.n422 B.n59 585
R147 B.n424 B.n423 585
R148 B.n425 B.n58 585
R149 B.n427 B.n426 585
R150 B.n428 B.n57 585
R151 B.n430 B.n429 585
R152 B.n431 B.n56 585
R153 B.n433 B.n432 585
R154 B.n434 B.n55 585
R155 B.n436 B.n435 585
R156 B.n437 B.n54 585
R157 B.n439 B.n438 585
R158 B.n440 B.n53 585
R159 B.n442 B.n441 585
R160 B.n443 B.n52 585
R161 B.n445 B.n444 585
R162 B.n446 B.n51 585
R163 B.n448 B.n447 585
R164 B.n449 B.n50 585
R165 B.n451 B.n450 585
R166 B.n452 B.n49 585
R167 B.n454 B.n453 585
R168 B.n455 B.n48 585
R169 B.n457 B.n456 585
R170 B.n458 B.n47 585
R171 B.n460 B.n459 585
R172 B.n461 B.n46 585
R173 B.n463 B.n462 585
R174 B.n464 B.n45 585
R175 B.n466 B.n465 585
R176 B.n468 B.n467 585
R177 B.n469 B.n41 585
R178 B.n471 B.n470 585
R179 B.n472 B.n40 585
R180 B.n474 B.n473 585
R181 B.n475 B.n39 585
R182 B.n477 B.n476 585
R183 B.n478 B.n38 585
R184 B.n480 B.n479 585
R185 B.n481 B.n35 585
R186 B.n484 B.n483 585
R187 B.n485 B.n34 585
R188 B.n487 B.n486 585
R189 B.n488 B.n33 585
R190 B.n490 B.n489 585
R191 B.n491 B.n32 585
R192 B.n493 B.n492 585
R193 B.n494 B.n31 585
R194 B.n496 B.n495 585
R195 B.n497 B.n30 585
R196 B.n499 B.n498 585
R197 B.n500 B.n29 585
R198 B.n502 B.n501 585
R199 B.n503 B.n28 585
R200 B.n505 B.n504 585
R201 B.n506 B.n27 585
R202 B.n508 B.n507 585
R203 B.n509 B.n26 585
R204 B.n511 B.n510 585
R205 B.n512 B.n25 585
R206 B.n514 B.n513 585
R207 B.n515 B.n24 585
R208 B.n517 B.n516 585
R209 B.n518 B.n23 585
R210 B.n520 B.n519 585
R211 B.n521 B.n22 585
R212 B.n523 B.n522 585
R213 B.n524 B.n21 585
R214 B.n526 B.n525 585
R215 B.n527 B.n20 585
R216 B.n529 B.n528 585
R217 B.n530 B.n19 585
R218 B.n532 B.n531 585
R219 B.n533 B.n18 585
R220 B.n535 B.n534 585
R221 B.n536 B.n17 585
R222 B.n538 B.n537 585
R223 B.n539 B.n16 585
R224 B.n541 B.n540 585
R225 B.n542 B.n15 585
R226 B.n544 B.n543 585
R227 B.n545 B.n14 585
R228 B.n547 B.n546 585
R229 B.n548 B.n13 585
R230 B.n550 B.n549 585
R231 B.n398 B.n67 585
R232 B.n397 B.n396 585
R233 B.n395 B.n68 585
R234 B.n394 B.n393 585
R235 B.n392 B.n69 585
R236 B.n391 B.n390 585
R237 B.n389 B.n70 585
R238 B.n388 B.n387 585
R239 B.n386 B.n71 585
R240 B.n385 B.n384 585
R241 B.n383 B.n72 585
R242 B.n382 B.n381 585
R243 B.n380 B.n73 585
R244 B.n379 B.n378 585
R245 B.n377 B.n74 585
R246 B.n376 B.n375 585
R247 B.n374 B.n75 585
R248 B.n373 B.n372 585
R249 B.n371 B.n76 585
R250 B.n370 B.n369 585
R251 B.n368 B.n77 585
R252 B.n367 B.n366 585
R253 B.n365 B.n78 585
R254 B.n364 B.n363 585
R255 B.n362 B.n79 585
R256 B.n361 B.n360 585
R257 B.n359 B.n80 585
R258 B.n358 B.n357 585
R259 B.n356 B.n81 585
R260 B.n355 B.n354 585
R261 B.n353 B.n82 585
R262 B.n352 B.n351 585
R263 B.n350 B.n83 585
R264 B.n349 B.n348 585
R265 B.n347 B.n84 585
R266 B.n346 B.n345 585
R267 B.n344 B.n85 585
R268 B.n343 B.n342 585
R269 B.n341 B.n86 585
R270 B.n340 B.n339 585
R271 B.n338 B.n87 585
R272 B.n337 B.n336 585
R273 B.n335 B.n88 585
R274 B.n184 B.n183 585
R275 B.n185 B.n142 585
R276 B.n187 B.n186 585
R277 B.n188 B.n141 585
R278 B.n190 B.n189 585
R279 B.n191 B.n140 585
R280 B.n193 B.n192 585
R281 B.n194 B.n139 585
R282 B.n196 B.n195 585
R283 B.n197 B.n138 585
R284 B.n199 B.n198 585
R285 B.n200 B.n137 585
R286 B.n202 B.n201 585
R287 B.n203 B.n136 585
R288 B.n205 B.n204 585
R289 B.n206 B.n135 585
R290 B.n208 B.n207 585
R291 B.n209 B.n134 585
R292 B.n211 B.n210 585
R293 B.n212 B.n133 585
R294 B.n214 B.n213 585
R295 B.n215 B.n132 585
R296 B.n217 B.n216 585
R297 B.n218 B.n131 585
R298 B.n220 B.n219 585
R299 B.n221 B.n130 585
R300 B.n223 B.n222 585
R301 B.n224 B.n129 585
R302 B.n226 B.n225 585
R303 B.n227 B.n128 585
R304 B.n229 B.n228 585
R305 B.n230 B.n127 585
R306 B.n232 B.n231 585
R307 B.n233 B.n126 585
R308 B.n235 B.n234 585
R309 B.n236 B.n125 585
R310 B.n238 B.n237 585
R311 B.n239 B.n124 585
R312 B.n241 B.n240 585
R313 B.n242 B.n123 585
R314 B.n244 B.n243 585
R315 B.n245 B.n122 585
R316 B.n247 B.n246 585
R317 B.n248 B.n121 585
R318 B.n250 B.n249 585
R319 B.n252 B.n251 585
R320 B.n253 B.n117 585
R321 B.n255 B.n254 585
R322 B.n256 B.n116 585
R323 B.n258 B.n257 585
R324 B.n259 B.n115 585
R325 B.n261 B.n260 585
R326 B.n262 B.n114 585
R327 B.n264 B.n263 585
R328 B.n265 B.n111 585
R329 B.n268 B.n267 585
R330 B.n269 B.n110 585
R331 B.n271 B.n270 585
R332 B.n272 B.n109 585
R333 B.n274 B.n273 585
R334 B.n275 B.n108 585
R335 B.n277 B.n276 585
R336 B.n278 B.n107 585
R337 B.n280 B.n279 585
R338 B.n281 B.n106 585
R339 B.n283 B.n282 585
R340 B.n284 B.n105 585
R341 B.n286 B.n285 585
R342 B.n287 B.n104 585
R343 B.n289 B.n288 585
R344 B.n290 B.n103 585
R345 B.n292 B.n291 585
R346 B.n293 B.n102 585
R347 B.n295 B.n294 585
R348 B.n296 B.n101 585
R349 B.n298 B.n297 585
R350 B.n299 B.n100 585
R351 B.n301 B.n300 585
R352 B.n302 B.n99 585
R353 B.n304 B.n303 585
R354 B.n305 B.n98 585
R355 B.n307 B.n306 585
R356 B.n308 B.n97 585
R357 B.n310 B.n309 585
R358 B.n311 B.n96 585
R359 B.n313 B.n312 585
R360 B.n314 B.n95 585
R361 B.n316 B.n315 585
R362 B.n317 B.n94 585
R363 B.n319 B.n318 585
R364 B.n320 B.n93 585
R365 B.n322 B.n321 585
R366 B.n323 B.n92 585
R367 B.n325 B.n324 585
R368 B.n326 B.n91 585
R369 B.n328 B.n327 585
R370 B.n329 B.n90 585
R371 B.n331 B.n330 585
R372 B.n332 B.n89 585
R373 B.n334 B.n333 585
R374 B.n182 B.n143 585
R375 B.n181 B.n180 585
R376 B.n179 B.n144 585
R377 B.n178 B.n177 585
R378 B.n176 B.n145 585
R379 B.n175 B.n174 585
R380 B.n173 B.n146 585
R381 B.n172 B.n171 585
R382 B.n170 B.n147 585
R383 B.n169 B.n168 585
R384 B.n167 B.n148 585
R385 B.n166 B.n165 585
R386 B.n164 B.n149 585
R387 B.n163 B.n162 585
R388 B.n161 B.n150 585
R389 B.n160 B.n159 585
R390 B.n158 B.n151 585
R391 B.n157 B.n156 585
R392 B.n155 B.n152 585
R393 B.n154 B.n153 585
R394 B.n2 B.n0 585
R395 B.n581 B.n1 585
R396 B.n580 B.n579 585
R397 B.n578 B.n3 585
R398 B.n577 B.n576 585
R399 B.n575 B.n4 585
R400 B.n574 B.n573 585
R401 B.n572 B.n5 585
R402 B.n571 B.n570 585
R403 B.n569 B.n6 585
R404 B.n568 B.n567 585
R405 B.n566 B.n7 585
R406 B.n565 B.n564 585
R407 B.n563 B.n8 585
R408 B.n562 B.n561 585
R409 B.n560 B.n9 585
R410 B.n559 B.n558 585
R411 B.n557 B.n10 585
R412 B.n556 B.n555 585
R413 B.n554 B.n11 585
R414 B.n553 B.n552 585
R415 B.n551 B.n12 585
R416 B.n583 B.n582 585
R417 B.n184 B.n143 478.086
R418 B.n551 B.n550 478.086
R419 B.n335 B.n334 478.086
R420 B.n400 B.n67 478.086
R421 B.n180 B.n143 163.367
R422 B.n180 B.n179 163.367
R423 B.n179 B.n178 163.367
R424 B.n178 B.n145 163.367
R425 B.n174 B.n145 163.367
R426 B.n174 B.n173 163.367
R427 B.n173 B.n172 163.367
R428 B.n172 B.n147 163.367
R429 B.n168 B.n147 163.367
R430 B.n168 B.n167 163.367
R431 B.n167 B.n166 163.367
R432 B.n166 B.n149 163.367
R433 B.n162 B.n149 163.367
R434 B.n162 B.n161 163.367
R435 B.n161 B.n160 163.367
R436 B.n160 B.n151 163.367
R437 B.n156 B.n151 163.367
R438 B.n156 B.n155 163.367
R439 B.n155 B.n154 163.367
R440 B.n154 B.n2 163.367
R441 B.n582 B.n2 163.367
R442 B.n582 B.n581 163.367
R443 B.n581 B.n580 163.367
R444 B.n580 B.n3 163.367
R445 B.n576 B.n3 163.367
R446 B.n576 B.n575 163.367
R447 B.n575 B.n574 163.367
R448 B.n574 B.n5 163.367
R449 B.n570 B.n5 163.367
R450 B.n570 B.n569 163.367
R451 B.n569 B.n568 163.367
R452 B.n568 B.n7 163.367
R453 B.n564 B.n7 163.367
R454 B.n564 B.n563 163.367
R455 B.n563 B.n562 163.367
R456 B.n562 B.n9 163.367
R457 B.n558 B.n9 163.367
R458 B.n558 B.n557 163.367
R459 B.n557 B.n556 163.367
R460 B.n556 B.n11 163.367
R461 B.n552 B.n11 163.367
R462 B.n552 B.n551 163.367
R463 B.n185 B.n184 163.367
R464 B.n186 B.n185 163.367
R465 B.n186 B.n141 163.367
R466 B.n190 B.n141 163.367
R467 B.n191 B.n190 163.367
R468 B.n192 B.n191 163.367
R469 B.n192 B.n139 163.367
R470 B.n196 B.n139 163.367
R471 B.n197 B.n196 163.367
R472 B.n198 B.n197 163.367
R473 B.n198 B.n137 163.367
R474 B.n202 B.n137 163.367
R475 B.n203 B.n202 163.367
R476 B.n204 B.n203 163.367
R477 B.n204 B.n135 163.367
R478 B.n208 B.n135 163.367
R479 B.n209 B.n208 163.367
R480 B.n210 B.n209 163.367
R481 B.n210 B.n133 163.367
R482 B.n214 B.n133 163.367
R483 B.n215 B.n214 163.367
R484 B.n216 B.n215 163.367
R485 B.n216 B.n131 163.367
R486 B.n220 B.n131 163.367
R487 B.n221 B.n220 163.367
R488 B.n222 B.n221 163.367
R489 B.n222 B.n129 163.367
R490 B.n226 B.n129 163.367
R491 B.n227 B.n226 163.367
R492 B.n228 B.n227 163.367
R493 B.n228 B.n127 163.367
R494 B.n232 B.n127 163.367
R495 B.n233 B.n232 163.367
R496 B.n234 B.n233 163.367
R497 B.n234 B.n125 163.367
R498 B.n238 B.n125 163.367
R499 B.n239 B.n238 163.367
R500 B.n240 B.n239 163.367
R501 B.n240 B.n123 163.367
R502 B.n244 B.n123 163.367
R503 B.n245 B.n244 163.367
R504 B.n246 B.n245 163.367
R505 B.n246 B.n121 163.367
R506 B.n250 B.n121 163.367
R507 B.n251 B.n250 163.367
R508 B.n251 B.n117 163.367
R509 B.n255 B.n117 163.367
R510 B.n256 B.n255 163.367
R511 B.n257 B.n256 163.367
R512 B.n257 B.n115 163.367
R513 B.n261 B.n115 163.367
R514 B.n262 B.n261 163.367
R515 B.n263 B.n262 163.367
R516 B.n263 B.n111 163.367
R517 B.n268 B.n111 163.367
R518 B.n269 B.n268 163.367
R519 B.n270 B.n269 163.367
R520 B.n270 B.n109 163.367
R521 B.n274 B.n109 163.367
R522 B.n275 B.n274 163.367
R523 B.n276 B.n275 163.367
R524 B.n276 B.n107 163.367
R525 B.n280 B.n107 163.367
R526 B.n281 B.n280 163.367
R527 B.n282 B.n281 163.367
R528 B.n282 B.n105 163.367
R529 B.n286 B.n105 163.367
R530 B.n287 B.n286 163.367
R531 B.n288 B.n287 163.367
R532 B.n288 B.n103 163.367
R533 B.n292 B.n103 163.367
R534 B.n293 B.n292 163.367
R535 B.n294 B.n293 163.367
R536 B.n294 B.n101 163.367
R537 B.n298 B.n101 163.367
R538 B.n299 B.n298 163.367
R539 B.n300 B.n299 163.367
R540 B.n300 B.n99 163.367
R541 B.n304 B.n99 163.367
R542 B.n305 B.n304 163.367
R543 B.n306 B.n305 163.367
R544 B.n306 B.n97 163.367
R545 B.n310 B.n97 163.367
R546 B.n311 B.n310 163.367
R547 B.n312 B.n311 163.367
R548 B.n312 B.n95 163.367
R549 B.n316 B.n95 163.367
R550 B.n317 B.n316 163.367
R551 B.n318 B.n317 163.367
R552 B.n318 B.n93 163.367
R553 B.n322 B.n93 163.367
R554 B.n323 B.n322 163.367
R555 B.n324 B.n323 163.367
R556 B.n324 B.n91 163.367
R557 B.n328 B.n91 163.367
R558 B.n329 B.n328 163.367
R559 B.n330 B.n329 163.367
R560 B.n330 B.n89 163.367
R561 B.n334 B.n89 163.367
R562 B.n336 B.n335 163.367
R563 B.n336 B.n87 163.367
R564 B.n340 B.n87 163.367
R565 B.n341 B.n340 163.367
R566 B.n342 B.n341 163.367
R567 B.n342 B.n85 163.367
R568 B.n346 B.n85 163.367
R569 B.n347 B.n346 163.367
R570 B.n348 B.n347 163.367
R571 B.n348 B.n83 163.367
R572 B.n352 B.n83 163.367
R573 B.n353 B.n352 163.367
R574 B.n354 B.n353 163.367
R575 B.n354 B.n81 163.367
R576 B.n358 B.n81 163.367
R577 B.n359 B.n358 163.367
R578 B.n360 B.n359 163.367
R579 B.n360 B.n79 163.367
R580 B.n364 B.n79 163.367
R581 B.n365 B.n364 163.367
R582 B.n366 B.n365 163.367
R583 B.n366 B.n77 163.367
R584 B.n370 B.n77 163.367
R585 B.n371 B.n370 163.367
R586 B.n372 B.n371 163.367
R587 B.n372 B.n75 163.367
R588 B.n376 B.n75 163.367
R589 B.n377 B.n376 163.367
R590 B.n378 B.n377 163.367
R591 B.n378 B.n73 163.367
R592 B.n382 B.n73 163.367
R593 B.n383 B.n382 163.367
R594 B.n384 B.n383 163.367
R595 B.n384 B.n71 163.367
R596 B.n388 B.n71 163.367
R597 B.n389 B.n388 163.367
R598 B.n390 B.n389 163.367
R599 B.n390 B.n69 163.367
R600 B.n394 B.n69 163.367
R601 B.n395 B.n394 163.367
R602 B.n396 B.n395 163.367
R603 B.n396 B.n67 163.367
R604 B.n550 B.n13 163.367
R605 B.n546 B.n13 163.367
R606 B.n546 B.n545 163.367
R607 B.n545 B.n544 163.367
R608 B.n544 B.n15 163.367
R609 B.n540 B.n15 163.367
R610 B.n540 B.n539 163.367
R611 B.n539 B.n538 163.367
R612 B.n538 B.n17 163.367
R613 B.n534 B.n17 163.367
R614 B.n534 B.n533 163.367
R615 B.n533 B.n532 163.367
R616 B.n532 B.n19 163.367
R617 B.n528 B.n19 163.367
R618 B.n528 B.n527 163.367
R619 B.n527 B.n526 163.367
R620 B.n526 B.n21 163.367
R621 B.n522 B.n21 163.367
R622 B.n522 B.n521 163.367
R623 B.n521 B.n520 163.367
R624 B.n520 B.n23 163.367
R625 B.n516 B.n23 163.367
R626 B.n516 B.n515 163.367
R627 B.n515 B.n514 163.367
R628 B.n514 B.n25 163.367
R629 B.n510 B.n25 163.367
R630 B.n510 B.n509 163.367
R631 B.n509 B.n508 163.367
R632 B.n508 B.n27 163.367
R633 B.n504 B.n27 163.367
R634 B.n504 B.n503 163.367
R635 B.n503 B.n502 163.367
R636 B.n502 B.n29 163.367
R637 B.n498 B.n29 163.367
R638 B.n498 B.n497 163.367
R639 B.n497 B.n496 163.367
R640 B.n496 B.n31 163.367
R641 B.n492 B.n31 163.367
R642 B.n492 B.n491 163.367
R643 B.n491 B.n490 163.367
R644 B.n490 B.n33 163.367
R645 B.n486 B.n33 163.367
R646 B.n486 B.n485 163.367
R647 B.n485 B.n484 163.367
R648 B.n484 B.n35 163.367
R649 B.n479 B.n35 163.367
R650 B.n479 B.n478 163.367
R651 B.n478 B.n477 163.367
R652 B.n477 B.n39 163.367
R653 B.n473 B.n39 163.367
R654 B.n473 B.n472 163.367
R655 B.n472 B.n471 163.367
R656 B.n471 B.n41 163.367
R657 B.n467 B.n41 163.367
R658 B.n467 B.n466 163.367
R659 B.n466 B.n45 163.367
R660 B.n462 B.n45 163.367
R661 B.n462 B.n461 163.367
R662 B.n461 B.n460 163.367
R663 B.n460 B.n47 163.367
R664 B.n456 B.n47 163.367
R665 B.n456 B.n455 163.367
R666 B.n455 B.n454 163.367
R667 B.n454 B.n49 163.367
R668 B.n450 B.n49 163.367
R669 B.n450 B.n449 163.367
R670 B.n449 B.n448 163.367
R671 B.n448 B.n51 163.367
R672 B.n444 B.n51 163.367
R673 B.n444 B.n443 163.367
R674 B.n443 B.n442 163.367
R675 B.n442 B.n53 163.367
R676 B.n438 B.n53 163.367
R677 B.n438 B.n437 163.367
R678 B.n437 B.n436 163.367
R679 B.n436 B.n55 163.367
R680 B.n432 B.n55 163.367
R681 B.n432 B.n431 163.367
R682 B.n431 B.n430 163.367
R683 B.n430 B.n57 163.367
R684 B.n426 B.n57 163.367
R685 B.n426 B.n425 163.367
R686 B.n425 B.n424 163.367
R687 B.n424 B.n59 163.367
R688 B.n420 B.n59 163.367
R689 B.n420 B.n419 163.367
R690 B.n419 B.n418 163.367
R691 B.n418 B.n61 163.367
R692 B.n414 B.n61 163.367
R693 B.n414 B.n413 163.367
R694 B.n413 B.n412 163.367
R695 B.n412 B.n63 163.367
R696 B.n408 B.n63 163.367
R697 B.n408 B.n407 163.367
R698 B.n407 B.n406 163.367
R699 B.n406 B.n65 163.367
R700 B.n402 B.n65 163.367
R701 B.n402 B.n401 163.367
R702 B.n401 B.n400 163.367
R703 B.n112 B.t11 128.584
R704 B.n42 B.t7 128.584
R705 B.n118 B.t5 128.569
R706 B.n36 B.t1 128.569
R707 B.n113 B.t10 111.519
R708 B.n43 B.t8 111.519
R709 B.n119 B.t4 111.502
R710 B.n37 B.t2 111.502
R711 B.n266 B.n113 59.5399
R712 B.n120 B.n119 59.5399
R713 B.n482 B.n37 59.5399
R714 B.n44 B.n43 59.5399
R715 B.n549 B.n12 31.0639
R716 B.n399 B.n398 31.0639
R717 B.n333 B.n88 31.0639
R718 B.n183 B.n182 31.0639
R719 B B.n583 18.0485
R720 B.n113 B.n112 17.0672
R721 B.n119 B.n118 17.0672
R722 B.n37 B.n36 17.0672
R723 B.n43 B.n42 17.0672
R724 B.n549 B.n548 10.6151
R725 B.n548 B.n547 10.6151
R726 B.n547 B.n14 10.6151
R727 B.n543 B.n14 10.6151
R728 B.n543 B.n542 10.6151
R729 B.n542 B.n541 10.6151
R730 B.n541 B.n16 10.6151
R731 B.n537 B.n16 10.6151
R732 B.n537 B.n536 10.6151
R733 B.n536 B.n535 10.6151
R734 B.n535 B.n18 10.6151
R735 B.n531 B.n18 10.6151
R736 B.n531 B.n530 10.6151
R737 B.n530 B.n529 10.6151
R738 B.n529 B.n20 10.6151
R739 B.n525 B.n20 10.6151
R740 B.n525 B.n524 10.6151
R741 B.n524 B.n523 10.6151
R742 B.n523 B.n22 10.6151
R743 B.n519 B.n22 10.6151
R744 B.n519 B.n518 10.6151
R745 B.n518 B.n517 10.6151
R746 B.n517 B.n24 10.6151
R747 B.n513 B.n24 10.6151
R748 B.n513 B.n512 10.6151
R749 B.n512 B.n511 10.6151
R750 B.n511 B.n26 10.6151
R751 B.n507 B.n26 10.6151
R752 B.n507 B.n506 10.6151
R753 B.n506 B.n505 10.6151
R754 B.n505 B.n28 10.6151
R755 B.n501 B.n28 10.6151
R756 B.n501 B.n500 10.6151
R757 B.n500 B.n499 10.6151
R758 B.n499 B.n30 10.6151
R759 B.n495 B.n30 10.6151
R760 B.n495 B.n494 10.6151
R761 B.n494 B.n493 10.6151
R762 B.n493 B.n32 10.6151
R763 B.n489 B.n32 10.6151
R764 B.n489 B.n488 10.6151
R765 B.n488 B.n487 10.6151
R766 B.n487 B.n34 10.6151
R767 B.n483 B.n34 10.6151
R768 B.n481 B.n480 10.6151
R769 B.n480 B.n38 10.6151
R770 B.n476 B.n38 10.6151
R771 B.n476 B.n475 10.6151
R772 B.n475 B.n474 10.6151
R773 B.n474 B.n40 10.6151
R774 B.n470 B.n40 10.6151
R775 B.n470 B.n469 10.6151
R776 B.n469 B.n468 10.6151
R777 B.n465 B.n464 10.6151
R778 B.n464 B.n463 10.6151
R779 B.n463 B.n46 10.6151
R780 B.n459 B.n46 10.6151
R781 B.n459 B.n458 10.6151
R782 B.n458 B.n457 10.6151
R783 B.n457 B.n48 10.6151
R784 B.n453 B.n48 10.6151
R785 B.n453 B.n452 10.6151
R786 B.n452 B.n451 10.6151
R787 B.n451 B.n50 10.6151
R788 B.n447 B.n50 10.6151
R789 B.n447 B.n446 10.6151
R790 B.n446 B.n445 10.6151
R791 B.n445 B.n52 10.6151
R792 B.n441 B.n52 10.6151
R793 B.n441 B.n440 10.6151
R794 B.n440 B.n439 10.6151
R795 B.n439 B.n54 10.6151
R796 B.n435 B.n54 10.6151
R797 B.n435 B.n434 10.6151
R798 B.n434 B.n433 10.6151
R799 B.n433 B.n56 10.6151
R800 B.n429 B.n56 10.6151
R801 B.n429 B.n428 10.6151
R802 B.n428 B.n427 10.6151
R803 B.n427 B.n58 10.6151
R804 B.n423 B.n58 10.6151
R805 B.n423 B.n422 10.6151
R806 B.n422 B.n421 10.6151
R807 B.n421 B.n60 10.6151
R808 B.n417 B.n60 10.6151
R809 B.n417 B.n416 10.6151
R810 B.n416 B.n415 10.6151
R811 B.n415 B.n62 10.6151
R812 B.n411 B.n62 10.6151
R813 B.n411 B.n410 10.6151
R814 B.n410 B.n409 10.6151
R815 B.n409 B.n64 10.6151
R816 B.n405 B.n64 10.6151
R817 B.n405 B.n404 10.6151
R818 B.n404 B.n403 10.6151
R819 B.n403 B.n66 10.6151
R820 B.n399 B.n66 10.6151
R821 B.n337 B.n88 10.6151
R822 B.n338 B.n337 10.6151
R823 B.n339 B.n338 10.6151
R824 B.n339 B.n86 10.6151
R825 B.n343 B.n86 10.6151
R826 B.n344 B.n343 10.6151
R827 B.n345 B.n344 10.6151
R828 B.n345 B.n84 10.6151
R829 B.n349 B.n84 10.6151
R830 B.n350 B.n349 10.6151
R831 B.n351 B.n350 10.6151
R832 B.n351 B.n82 10.6151
R833 B.n355 B.n82 10.6151
R834 B.n356 B.n355 10.6151
R835 B.n357 B.n356 10.6151
R836 B.n357 B.n80 10.6151
R837 B.n361 B.n80 10.6151
R838 B.n362 B.n361 10.6151
R839 B.n363 B.n362 10.6151
R840 B.n363 B.n78 10.6151
R841 B.n367 B.n78 10.6151
R842 B.n368 B.n367 10.6151
R843 B.n369 B.n368 10.6151
R844 B.n369 B.n76 10.6151
R845 B.n373 B.n76 10.6151
R846 B.n374 B.n373 10.6151
R847 B.n375 B.n374 10.6151
R848 B.n375 B.n74 10.6151
R849 B.n379 B.n74 10.6151
R850 B.n380 B.n379 10.6151
R851 B.n381 B.n380 10.6151
R852 B.n381 B.n72 10.6151
R853 B.n385 B.n72 10.6151
R854 B.n386 B.n385 10.6151
R855 B.n387 B.n386 10.6151
R856 B.n387 B.n70 10.6151
R857 B.n391 B.n70 10.6151
R858 B.n392 B.n391 10.6151
R859 B.n393 B.n392 10.6151
R860 B.n393 B.n68 10.6151
R861 B.n397 B.n68 10.6151
R862 B.n398 B.n397 10.6151
R863 B.n183 B.n142 10.6151
R864 B.n187 B.n142 10.6151
R865 B.n188 B.n187 10.6151
R866 B.n189 B.n188 10.6151
R867 B.n189 B.n140 10.6151
R868 B.n193 B.n140 10.6151
R869 B.n194 B.n193 10.6151
R870 B.n195 B.n194 10.6151
R871 B.n195 B.n138 10.6151
R872 B.n199 B.n138 10.6151
R873 B.n200 B.n199 10.6151
R874 B.n201 B.n200 10.6151
R875 B.n201 B.n136 10.6151
R876 B.n205 B.n136 10.6151
R877 B.n206 B.n205 10.6151
R878 B.n207 B.n206 10.6151
R879 B.n207 B.n134 10.6151
R880 B.n211 B.n134 10.6151
R881 B.n212 B.n211 10.6151
R882 B.n213 B.n212 10.6151
R883 B.n213 B.n132 10.6151
R884 B.n217 B.n132 10.6151
R885 B.n218 B.n217 10.6151
R886 B.n219 B.n218 10.6151
R887 B.n219 B.n130 10.6151
R888 B.n223 B.n130 10.6151
R889 B.n224 B.n223 10.6151
R890 B.n225 B.n224 10.6151
R891 B.n225 B.n128 10.6151
R892 B.n229 B.n128 10.6151
R893 B.n230 B.n229 10.6151
R894 B.n231 B.n230 10.6151
R895 B.n231 B.n126 10.6151
R896 B.n235 B.n126 10.6151
R897 B.n236 B.n235 10.6151
R898 B.n237 B.n236 10.6151
R899 B.n237 B.n124 10.6151
R900 B.n241 B.n124 10.6151
R901 B.n242 B.n241 10.6151
R902 B.n243 B.n242 10.6151
R903 B.n243 B.n122 10.6151
R904 B.n247 B.n122 10.6151
R905 B.n248 B.n247 10.6151
R906 B.n249 B.n248 10.6151
R907 B.n253 B.n252 10.6151
R908 B.n254 B.n253 10.6151
R909 B.n254 B.n116 10.6151
R910 B.n258 B.n116 10.6151
R911 B.n259 B.n258 10.6151
R912 B.n260 B.n259 10.6151
R913 B.n260 B.n114 10.6151
R914 B.n264 B.n114 10.6151
R915 B.n265 B.n264 10.6151
R916 B.n267 B.n110 10.6151
R917 B.n271 B.n110 10.6151
R918 B.n272 B.n271 10.6151
R919 B.n273 B.n272 10.6151
R920 B.n273 B.n108 10.6151
R921 B.n277 B.n108 10.6151
R922 B.n278 B.n277 10.6151
R923 B.n279 B.n278 10.6151
R924 B.n279 B.n106 10.6151
R925 B.n283 B.n106 10.6151
R926 B.n284 B.n283 10.6151
R927 B.n285 B.n284 10.6151
R928 B.n285 B.n104 10.6151
R929 B.n289 B.n104 10.6151
R930 B.n290 B.n289 10.6151
R931 B.n291 B.n290 10.6151
R932 B.n291 B.n102 10.6151
R933 B.n295 B.n102 10.6151
R934 B.n296 B.n295 10.6151
R935 B.n297 B.n296 10.6151
R936 B.n297 B.n100 10.6151
R937 B.n301 B.n100 10.6151
R938 B.n302 B.n301 10.6151
R939 B.n303 B.n302 10.6151
R940 B.n303 B.n98 10.6151
R941 B.n307 B.n98 10.6151
R942 B.n308 B.n307 10.6151
R943 B.n309 B.n308 10.6151
R944 B.n309 B.n96 10.6151
R945 B.n313 B.n96 10.6151
R946 B.n314 B.n313 10.6151
R947 B.n315 B.n314 10.6151
R948 B.n315 B.n94 10.6151
R949 B.n319 B.n94 10.6151
R950 B.n320 B.n319 10.6151
R951 B.n321 B.n320 10.6151
R952 B.n321 B.n92 10.6151
R953 B.n325 B.n92 10.6151
R954 B.n326 B.n325 10.6151
R955 B.n327 B.n326 10.6151
R956 B.n327 B.n90 10.6151
R957 B.n331 B.n90 10.6151
R958 B.n332 B.n331 10.6151
R959 B.n333 B.n332 10.6151
R960 B.n182 B.n181 10.6151
R961 B.n181 B.n144 10.6151
R962 B.n177 B.n144 10.6151
R963 B.n177 B.n176 10.6151
R964 B.n176 B.n175 10.6151
R965 B.n175 B.n146 10.6151
R966 B.n171 B.n146 10.6151
R967 B.n171 B.n170 10.6151
R968 B.n170 B.n169 10.6151
R969 B.n169 B.n148 10.6151
R970 B.n165 B.n148 10.6151
R971 B.n165 B.n164 10.6151
R972 B.n164 B.n163 10.6151
R973 B.n163 B.n150 10.6151
R974 B.n159 B.n150 10.6151
R975 B.n159 B.n158 10.6151
R976 B.n158 B.n157 10.6151
R977 B.n157 B.n152 10.6151
R978 B.n153 B.n152 10.6151
R979 B.n153 B.n0 10.6151
R980 B.n579 B.n1 10.6151
R981 B.n579 B.n578 10.6151
R982 B.n578 B.n577 10.6151
R983 B.n577 B.n4 10.6151
R984 B.n573 B.n4 10.6151
R985 B.n573 B.n572 10.6151
R986 B.n572 B.n571 10.6151
R987 B.n571 B.n6 10.6151
R988 B.n567 B.n6 10.6151
R989 B.n567 B.n566 10.6151
R990 B.n566 B.n565 10.6151
R991 B.n565 B.n8 10.6151
R992 B.n561 B.n8 10.6151
R993 B.n561 B.n560 10.6151
R994 B.n560 B.n559 10.6151
R995 B.n559 B.n10 10.6151
R996 B.n555 B.n10 10.6151
R997 B.n555 B.n554 10.6151
R998 B.n554 B.n553 10.6151
R999 B.n553 B.n12 10.6151
R1000 B.n483 B.n482 9.36635
R1001 B.n465 B.n44 9.36635
R1002 B.n249 B.n120 9.36635
R1003 B.n267 B.n266 9.36635
R1004 B.n583 B.n0 2.81026
R1005 B.n583 B.n1 2.81026
R1006 B.n482 B.n481 1.24928
R1007 B.n468 B.n44 1.24928
R1008 B.n252 B.n120 1.24928
R1009 B.n266 B.n265 1.24928
C0 VN VP 5.370029f
C1 VDD2 VP 0.301758f
C2 w_n1850_n3600# VP 3.44927f
C3 VP VDD1 5.41756f
C4 VTAIL VN 4.91262f
C5 VDD2 VTAIL 13.415901f
C6 VTAIL w_n1850_n3600# 4.529f
C7 VTAIL VDD1 13.3752f
C8 B VP 1.14294f
C9 VDD2 VN 5.26441f
C10 w_n1850_n3600# VN 3.21515f
C11 VN VDD1 0.148251f
C12 VTAIL B 4.02001f
C13 VDD2 w_n1850_n3600# 1.29945f
C14 VDD2 VDD1 0.751778f
C15 w_n1850_n3600# VDD1 1.27082f
C16 VTAIL VP 4.92672f
C17 B VN 0.761393f
C18 VDD2 B 1.08748f
C19 B w_n1850_n3600# 7.30457f
C20 B VDD1 1.05545f
C21 VDD2 VSUBS 1.373825f
C22 VDD1 VSUBS 1.652923f
C23 VTAIL VSUBS 0.885753f
C24 VN VSUBS 4.67942f
C25 VP VSUBS 1.534175f
C26 B VSUBS 2.80997f
C27 w_n1850_n3600# VSUBS 81.851395f
C28 B.n0 VSUBS 0.005186f
C29 B.n1 VSUBS 0.005186f
C30 B.n2 VSUBS 0.008202f
C31 B.n3 VSUBS 0.008202f
C32 B.n4 VSUBS 0.008202f
C33 B.n5 VSUBS 0.008202f
C34 B.n6 VSUBS 0.008202f
C35 B.n7 VSUBS 0.008202f
C36 B.n8 VSUBS 0.008202f
C37 B.n9 VSUBS 0.008202f
C38 B.n10 VSUBS 0.008202f
C39 B.n11 VSUBS 0.008202f
C40 B.n12 VSUBS 0.017891f
C41 B.n13 VSUBS 0.008202f
C42 B.n14 VSUBS 0.008202f
C43 B.n15 VSUBS 0.008202f
C44 B.n16 VSUBS 0.008202f
C45 B.n17 VSUBS 0.008202f
C46 B.n18 VSUBS 0.008202f
C47 B.n19 VSUBS 0.008202f
C48 B.n20 VSUBS 0.008202f
C49 B.n21 VSUBS 0.008202f
C50 B.n22 VSUBS 0.008202f
C51 B.n23 VSUBS 0.008202f
C52 B.n24 VSUBS 0.008202f
C53 B.n25 VSUBS 0.008202f
C54 B.n26 VSUBS 0.008202f
C55 B.n27 VSUBS 0.008202f
C56 B.n28 VSUBS 0.008202f
C57 B.n29 VSUBS 0.008202f
C58 B.n30 VSUBS 0.008202f
C59 B.n31 VSUBS 0.008202f
C60 B.n32 VSUBS 0.008202f
C61 B.n33 VSUBS 0.008202f
C62 B.n34 VSUBS 0.008202f
C63 B.n35 VSUBS 0.008202f
C64 B.t2 VSUBS 0.507252f
C65 B.t1 VSUBS 0.515555f
C66 B.t0 VSUBS 0.342555f
C67 B.n36 VSUBS 0.152491f
C68 B.n37 VSUBS 0.074248f
C69 B.n38 VSUBS 0.008202f
C70 B.n39 VSUBS 0.008202f
C71 B.n40 VSUBS 0.008202f
C72 B.n41 VSUBS 0.008202f
C73 B.t8 VSUBS 0.507241f
C74 B.t7 VSUBS 0.515545f
C75 B.t6 VSUBS 0.342555f
C76 B.n42 VSUBS 0.152502f
C77 B.n43 VSUBS 0.074259f
C78 B.n44 VSUBS 0.019002f
C79 B.n45 VSUBS 0.008202f
C80 B.n46 VSUBS 0.008202f
C81 B.n47 VSUBS 0.008202f
C82 B.n48 VSUBS 0.008202f
C83 B.n49 VSUBS 0.008202f
C84 B.n50 VSUBS 0.008202f
C85 B.n51 VSUBS 0.008202f
C86 B.n52 VSUBS 0.008202f
C87 B.n53 VSUBS 0.008202f
C88 B.n54 VSUBS 0.008202f
C89 B.n55 VSUBS 0.008202f
C90 B.n56 VSUBS 0.008202f
C91 B.n57 VSUBS 0.008202f
C92 B.n58 VSUBS 0.008202f
C93 B.n59 VSUBS 0.008202f
C94 B.n60 VSUBS 0.008202f
C95 B.n61 VSUBS 0.008202f
C96 B.n62 VSUBS 0.008202f
C97 B.n63 VSUBS 0.008202f
C98 B.n64 VSUBS 0.008202f
C99 B.n65 VSUBS 0.008202f
C100 B.n66 VSUBS 0.008202f
C101 B.n67 VSUBS 0.017891f
C102 B.n68 VSUBS 0.008202f
C103 B.n69 VSUBS 0.008202f
C104 B.n70 VSUBS 0.008202f
C105 B.n71 VSUBS 0.008202f
C106 B.n72 VSUBS 0.008202f
C107 B.n73 VSUBS 0.008202f
C108 B.n74 VSUBS 0.008202f
C109 B.n75 VSUBS 0.008202f
C110 B.n76 VSUBS 0.008202f
C111 B.n77 VSUBS 0.008202f
C112 B.n78 VSUBS 0.008202f
C113 B.n79 VSUBS 0.008202f
C114 B.n80 VSUBS 0.008202f
C115 B.n81 VSUBS 0.008202f
C116 B.n82 VSUBS 0.008202f
C117 B.n83 VSUBS 0.008202f
C118 B.n84 VSUBS 0.008202f
C119 B.n85 VSUBS 0.008202f
C120 B.n86 VSUBS 0.008202f
C121 B.n87 VSUBS 0.008202f
C122 B.n88 VSUBS 0.017891f
C123 B.n89 VSUBS 0.008202f
C124 B.n90 VSUBS 0.008202f
C125 B.n91 VSUBS 0.008202f
C126 B.n92 VSUBS 0.008202f
C127 B.n93 VSUBS 0.008202f
C128 B.n94 VSUBS 0.008202f
C129 B.n95 VSUBS 0.008202f
C130 B.n96 VSUBS 0.008202f
C131 B.n97 VSUBS 0.008202f
C132 B.n98 VSUBS 0.008202f
C133 B.n99 VSUBS 0.008202f
C134 B.n100 VSUBS 0.008202f
C135 B.n101 VSUBS 0.008202f
C136 B.n102 VSUBS 0.008202f
C137 B.n103 VSUBS 0.008202f
C138 B.n104 VSUBS 0.008202f
C139 B.n105 VSUBS 0.008202f
C140 B.n106 VSUBS 0.008202f
C141 B.n107 VSUBS 0.008202f
C142 B.n108 VSUBS 0.008202f
C143 B.n109 VSUBS 0.008202f
C144 B.n110 VSUBS 0.008202f
C145 B.n111 VSUBS 0.008202f
C146 B.t10 VSUBS 0.507241f
C147 B.t11 VSUBS 0.515545f
C148 B.t9 VSUBS 0.342555f
C149 B.n112 VSUBS 0.152502f
C150 B.n113 VSUBS 0.074259f
C151 B.n114 VSUBS 0.008202f
C152 B.n115 VSUBS 0.008202f
C153 B.n116 VSUBS 0.008202f
C154 B.n117 VSUBS 0.008202f
C155 B.t4 VSUBS 0.507252f
C156 B.t5 VSUBS 0.515555f
C157 B.t3 VSUBS 0.342555f
C158 B.n118 VSUBS 0.152491f
C159 B.n119 VSUBS 0.074248f
C160 B.n120 VSUBS 0.019002f
C161 B.n121 VSUBS 0.008202f
C162 B.n122 VSUBS 0.008202f
C163 B.n123 VSUBS 0.008202f
C164 B.n124 VSUBS 0.008202f
C165 B.n125 VSUBS 0.008202f
C166 B.n126 VSUBS 0.008202f
C167 B.n127 VSUBS 0.008202f
C168 B.n128 VSUBS 0.008202f
C169 B.n129 VSUBS 0.008202f
C170 B.n130 VSUBS 0.008202f
C171 B.n131 VSUBS 0.008202f
C172 B.n132 VSUBS 0.008202f
C173 B.n133 VSUBS 0.008202f
C174 B.n134 VSUBS 0.008202f
C175 B.n135 VSUBS 0.008202f
C176 B.n136 VSUBS 0.008202f
C177 B.n137 VSUBS 0.008202f
C178 B.n138 VSUBS 0.008202f
C179 B.n139 VSUBS 0.008202f
C180 B.n140 VSUBS 0.008202f
C181 B.n141 VSUBS 0.008202f
C182 B.n142 VSUBS 0.008202f
C183 B.n143 VSUBS 0.017891f
C184 B.n144 VSUBS 0.008202f
C185 B.n145 VSUBS 0.008202f
C186 B.n146 VSUBS 0.008202f
C187 B.n147 VSUBS 0.008202f
C188 B.n148 VSUBS 0.008202f
C189 B.n149 VSUBS 0.008202f
C190 B.n150 VSUBS 0.008202f
C191 B.n151 VSUBS 0.008202f
C192 B.n152 VSUBS 0.008202f
C193 B.n153 VSUBS 0.008202f
C194 B.n154 VSUBS 0.008202f
C195 B.n155 VSUBS 0.008202f
C196 B.n156 VSUBS 0.008202f
C197 B.n157 VSUBS 0.008202f
C198 B.n158 VSUBS 0.008202f
C199 B.n159 VSUBS 0.008202f
C200 B.n160 VSUBS 0.008202f
C201 B.n161 VSUBS 0.008202f
C202 B.n162 VSUBS 0.008202f
C203 B.n163 VSUBS 0.008202f
C204 B.n164 VSUBS 0.008202f
C205 B.n165 VSUBS 0.008202f
C206 B.n166 VSUBS 0.008202f
C207 B.n167 VSUBS 0.008202f
C208 B.n168 VSUBS 0.008202f
C209 B.n169 VSUBS 0.008202f
C210 B.n170 VSUBS 0.008202f
C211 B.n171 VSUBS 0.008202f
C212 B.n172 VSUBS 0.008202f
C213 B.n173 VSUBS 0.008202f
C214 B.n174 VSUBS 0.008202f
C215 B.n175 VSUBS 0.008202f
C216 B.n176 VSUBS 0.008202f
C217 B.n177 VSUBS 0.008202f
C218 B.n178 VSUBS 0.008202f
C219 B.n179 VSUBS 0.008202f
C220 B.n180 VSUBS 0.008202f
C221 B.n181 VSUBS 0.008202f
C222 B.n182 VSUBS 0.017891f
C223 B.n183 VSUBS 0.019258f
C224 B.n184 VSUBS 0.019258f
C225 B.n185 VSUBS 0.008202f
C226 B.n186 VSUBS 0.008202f
C227 B.n187 VSUBS 0.008202f
C228 B.n188 VSUBS 0.008202f
C229 B.n189 VSUBS 0.008202f
C230 B.n190 VSUBS 0.008202f
C231 B.n191 VSUBS 0.008202f
C232 B.n192 VSUBS 0.008202f
C233 B.n193 VSUBS 0.008202f
C234 B.n194 VSUBS 0.008202f
C235 B.n195 VSUBS 0.008202f
C236 B.n196 VSUBS 0.008202f
C237 B.n197 VSUBS 0.008202f
C238 B.n198 VSUBS 0.008202f
C239 B.n199 VSUBS 0.008202f
C240 B.n200 VSUBS 0.008202f
C241 B.n201 VSUBS 0.008202f
C242 B.n202 VSUBS 0.008202f
C243 B.n203 VSUBS 0.008202f
C244 B.n204 VSUBS 0.008202f
C245 B.n205 VSUBS 0.008202f
C246 B.n206 VSUBS 0.008202f
C247 B.n207 VSUBS 0.008202f
C248 B.n208 VSUBS 0.008202f
C249 B.n209 VSUBS 0.008202f
C250 B.n210 VSUBS 0.008202f
C251 B.n211 VSUBS 0.008202f
C252 B.n212 VSUBS 0.008202f
C253 B.n213 VSUBS 0.008202f
C254 B.n214 VSUBS 0.008202f
C255 B.n215 VSUBS 0.008202f
C256 B.n216 VSUBS 0.008202f
C257 B.n217 VSUBS 0.008202f
C258 B.n218 VSUBS 0.008202f
C259 B.n219 VSUBS 0.008202f
C260 B.n220 VSUBS 0.008202f
C261 B.n221 VSUBS 0.008202f
C262 B.n222 VSUBS 0.008202f
C263 B.n223 VSUBS 0.008202f
C264 B.n224 VSUBS 0.008202f
C265 B.n225 VSUBS 0.008202f
C266 B.n226 VSUBS 0.008202f
C267 B.n227 VSUBS 0.008202f
C268 B.n228 VSUBS 0.008202f
C269 B.n229 VSUBS 0.008202f
C270 B.n230 VSUBS 0.008202f
C271 B.n231 VSUBS 0.008202f
C272 B.n232 VSUBS 0.008202f
C273 B.n233 VSUBS 0.008202f
C274 B.n234 VSUBS 0.008202f
C275 B.n235 VSUBS 0.008202f
C276 B.n236 VSUBS 0.008202f
C277 B.n237 VSUBS 0.008202f
C278 B.n238 VSUBS 0.008202f
C279 B.n239 VSUBS 0.008202f
C280 B.n240 VSUBS 0.008202f
C281 B.n241 VSUBS 0.008202f
C282 B.n242 VSUBS 0.008202f
C283 B.n243 VSUBS 0.008202f
C284 B.n244 VSUBS 0.008202f
C285 B.n245 VSUBS 0.008202f
C286 B.n246 VSUBS 0.008202f
C287 B.n247 VSUBS 0.008202f
C288 B.n248 VSUBS 0.008202f
C289 B.n249 VSUBS 0.007719f
C290 B.n250 VSUBS 0.008202f
C291 B.n251 VSUBS 0.008202f
C292 B.n252 VSUBS 0.004583f
C293 B.n253 VSUBS 0.008202f
C294 B.n254 VSUBS 0.008202f
C295 B.n255 VSUBS 0.008202f
C296 B.n256 VSUBS 0.008202f
C297 B.n257 VSUBS 0.008202f
C298 B.n258 VSUBS 0.008202f
C299 B.n259 VSUBS 0.008202f
C300 B.n260 VSUBS 0.008202f
C301 B.n261 VSUBS 0.008202f
C302 B.n262 VSUBS 0.008202f
C303 B.n263 VSUBS 0.008202f
C304 B.n264 VSUBS 0.008202f
C305 B.n265 VSUBS 0.004583f
C306 B.n266 VSUBS 0.019002f
C307 B.n267 VSUBS 0.007719f
C308 B.n268 VSUBS 0.008202f
C309 B.n269 VSUBS 0.008202f
C310 B.n270 VSUBS 0.008202f
C311 B.n271 VSUBS 0.008202f
C312 B.n272 VSUBS 0.008202f
C313 B.n273 VSUBS 0.008202f
C314 B.n274 VSUBS 0.008202f
C315 B.n275 VSUBS 0.008202f
C316 B.n276 VSUBS 0.008202f
C317 B.n277 VSUBS 0.008202f
C318 B.n278 VSUBS 0.008202f
C319 B.n279 VSUBS 0.008202f
C320 B.n280 VSUBS 0.008202f
C321 B.n281 VSUBS 0.008202f
C322 B.n282 VSUBS 0.008202f
C323 B.n283 VSUBS 0.008202f
C324 B.n284 VSUBS 0.008202f
C325 B.n285 VSUBS 0.008202f
C326 B.n286 VSUBS 0.008202f
C327 B.n287 VSUBS 0.008202f
C328 B.n288 VSUBS 0.008202f
C329 B.n289 VSUBS 0.008202f
C330 B.n290 VSUBS 0.008202f
C331 B.n291 VSUBS 0.008202f
C332 B.n292 VSUBS 0.008202f
C333 B.n293 VSUBS 0.008202f
C334 B.n294 VSUBS 0.008202f
C335 B.n295 VSUBS 0.008202f
C336 B.n296 VSUBS 0.008202f
C337 B.n297 VSUBS 0.008202f
C338 B.n298 VSUBS 0.008202f
C339 B.n299 VSUBS 0.008202f
C340 B.n300 VSUBS 0.008202f
C341 B.n301 VSUBS 0.008202f
C342 B.n302 VSUBS 0.008202f
C343 B.n303 VSUBS 0.008202f
C344 B.n304 VSUBS 0.008202f
C345 B.n305 VSUBS 0.008202f
C346 B.n306 VSUBS 0.008202f
C347 B.n307 VSUBS 0.008202f
C348 B.n308 VSUBS 0.008202f
C349 B.n309 VSUBS 0.008202f
C350 B.n310 VSUBS 0.008202f
C351 B.n311 VSUBS 0.008202f
C352 B.n312 VSUBS 0.008202f
C353 B.n313 VSUBS 0.008202f
C354 B.n314 VSUBS 0.008202f
C355 B.n315 VSUBS 0.008202f
C356 B.n316 VSUBS 0.008202f
C357 B.n317 VSUBS 0.008202f
C358 B.n318 VSUBS 0.008202f
C359 B.n319 VSUBS 0.008202f
C360 B.n320 VSUBS 0.008202f
C361 B.n321 VSUBS 0.008202f
C362 B.n322 VSUBS 0.008202f
C363 B.n323 VSUBS 0.008202f
C364 B.n324 VSUBS 0.008202f
C365 B.n325 VSUBS 0.008202f
C366 B.n326 VSUBS 0.008202f
C367 B.n327 VSUBS 0.008202f
C368 B.n328 VSUBS 0.008202f
C369 B.n329 VSUBS 0.008202f
C370 B.n330 VSUBS 0.008202f
C371 B.n331 VSUBS 0.008202f
C372 B.n332 VSUBS 0.008202f
C373 B.n333 VSUBS 0.019258f
C374 B.n334 VSUBS 0.019258f
C375 B.n335 VSUBS 0.017891f
C376 B.n336 VSUBS 0.008202f
C377 B.n337 VSUBS 0.008202f
C378 B.n338 VSUBS 0.008202f
C379 B.n339 VSUBS 0.008202f
C380 B.n340 VSUBS 0.008202f
C381 B.n341 VSUBS 0.008202f
C382 B.n342 VSUBS 0.008202f
C383 B.n343 VSUBS 0.008202f
C384 B.n344 VSUBS 0.008202f
C385 B.n345 VSUBS 0.008202f
C386 B.n346 VSUBS 0.008202f
C387 B.n347 VSUBS 0.008202f
C388 B.n348 VSUBS 0.008202f
C389 B.n349 VSUBS 0.008202f
C390 B.n350 VSUBS 0.008202f
C391 B.n351 VSUBS 0.008202f
C392 B.n352 VSUBS 0.008202f
C393 B.n353 VSUBS 0.008202f
C394 B.n354 VSUBS 0.008202f
C395 B.n355 VSUBS 0.008202f
C396 B.n356 VSUBS 0.008202f
C397 B.n357 VSUBS 0.008202f
C398 B.n358 VSUBS 0.008202f
C399 B.n359 VSUBS 0.008202f
C400 B.n360 VSUBS 0.008202f
C401 B.n361 VSUBS 0.008202f
C402 B.n362 VSUBS 0.008202f
C403 B.n363 VSUBS 0.008202f
C404 B.n364 VSUBS 0.008202f
C405 B.n365 VSUBS 0.008202f
C406 B.n366 VSUBS 0.008202f
C407 B.n367 VSUBS 0.008202f
C408 B.n368 VSUBS 0.008202f
C409 B.n369 VSUBS 0.008202f
C410 B.n370 VSUBS 0.008202f
C411 B.n371 VSUBS 0.008202f
C412 B.n372 VSUBS 0.008202f
C413 B.n373 VSUBS 0.008202f
C414 B.n374 VSUBS 0.008202f
C415 B.n375 VSUBS 0.008202f
C416 B.n376 VSUBS 0.008202f
C417 B.n377 VSUBS 0.008202f
C418 B.n378 VSUBS 0.008202f
C419 B.n379 VSUBS 0.008202f
C420 B.n380 VSUBS 0.008202f
C421 B.n381 VSUBS 0.008202f
C422 B.n382 VSUBS 0.008202f
C423 B.n383 VSUBS 0.008202f
C424 B.n384 VSUBS 0.008202f
C425 B.n385 VSUBS 0.008202f
C426 B.n386 VSUBS 0.008202f
C427 B.n387 VSUBS 0.008202f
C428 B.n388 VSUBS 0.008202f
C429 B.n389 VSUBS 0.008202f
C430 B.n390 VSUBS 0.008202f
C431 B.n391 VSUBS 0.008202f
C432 B.n392 VSUBS 0.008202f
C433 B.n393 VSUBS 0.008202f
C434 B.n394 VSUBS 0.008202f
C435 B.n395 VSUBS 0.008202f
C436 B.n396 VSUBS 0.008202f
C437 B.n397 VSUBS 0.008202f
C438 B.n398 VSUBS 0.01891f
C439 B.n399 VSUBS 0.018239f
C440 B.n400 VSUBS 0.019258f
C441 B.n401 VSUBS 0.008202f
C442 B.n402 VSUBS 0.008202f
C443 B.n403 VSUBS 0.008202f
C444 B.n404 VSUBS 0.008202f
C445 B.n405 VSUBS 0.008202f
C446 B.n406 VSUBS 0.008202f
C447 B.n407 VSUBS 0.008202f
C448 B.n408 VSUBS 0.008202f
C449 B.n409 VSUBS 0.008202f
C450 B.n410 VSUBS 0.008202f
C451 B.n411 VSUBS 0.008202f
C452 B.n412 VSUBS 0.008202f
C453 B.n413 VSUBS 0.008202f
C454 B.n414 VSUBS 0.008202f
C455 B.n415 VSUBS 0.008202f
C456 B.n416 VSUBS 0.008202f
C457 B.n417 VSUBS 0.008202f
C458 B.n418 VSUBS 0.008202f
C459 B.n419 VSUBS 0.008202f
C460 B.n420 VSUBS 0.008202f
C461 B.n421 VSUBS 0.008202f
C462 B.n422 VSUBS 0.008202f
C463 B.n423 VSUBS 0.008202f
C464 B.n424 VSUBS 0.008202f
C465 B.n425 VSUBS 0.008202f
C466 B.n426 VSUBS 0.008202f
C467 B.n427 VSUBS 0.008202f
C468 B.n428 VSUBS 0.008202f
C469 B.n429 VSUBS 0.008202f
C470 B.n430 VSUBS 0.008202f
C471 B.n431 VSUBS 0.008202f
C472 B.n432 VSUBS 0.008202f
C473 B.n433 VSUBS 0.008202f
C474 B.n434 VSUBS 0.008202f
C475 B.n435 VSUBS 0.008202f
C476 B.n436 VSUBS 0.008202f
C477 B.n437 VSUBS 0.008202f
C478 B.n438 VSUBS 0.008202f
C479 B.n439 VSUBS 0.008202f
C480 B.n440 VSUBS 0.008202f
C481 B.n441 VSUBS 0.008202f
C482 B.n442 VSUBS 0.008202f
C483 B.n443 VSUBS 0.008202f
C484 B.n444 VSUBS 0.008202f
C485 B.n445 VSUBS 0.008202f
C486 B.n446 VSUBS 0.008202f
C487 B.n447 VSUBS 0.008202f
C488 B.n448 VSUBS 0.008202f
C489 B.n449 VSUBS 0.008202f
C490 B.n450 VSUBS 0.008202f
C491 B.n451 VSUBS 0.008202f
C492 B.n452 VSUBS 0.008202f
C493 B.n453 VSUBS 0.008202f
C494 B.n454 VSUBS 0.008202f
C495 B.n455 VSUBS 0.008202f
C496 B.n456 VSUBS 0.008202f
C497 B.n457 VSUBS 0.008202f
C498 B.n458 VSUBS 0.008202f
C499 B.n459 VSUBS 0.008202f
C500 B.n460 VSUBS 0.008202f
C501 B.n461 VSUBS 0.008202f
C502 B.n462 VSUBS 0.008202f
C503 B.n463 VSUBS 0.008202f
C504 B.n464 VSUBS 0.008202f
C505 B.n465 VSUBS 0.007719f
C506 B.n466 VSUBS 0.008202f
C507 B.n467 VSUBS 0.008202f
C508 B.n468 VSUBS 0.004583f
C509 B.n469 VSUBS 0.008202f
C510 B.n470 VSUBS 0.008202f
C511 B.n471 VSUBS 0.008202f
C512 B.n472 VSUBS 0.008202f
C513 B.n473 VSUBS 0.008202f
C514 B.n474 VSUBS 0.008202f
C515 B.n475 VSUBS 0.008202f
C516 B.n476 VSUBS 0.008202f
C517 B.n477 VSUBS 0.008202f
C518 B.n478 VSUBS 0.008202f
C519 B.n479 VSUBS 0.008202f
C520 B.n480 VSUBS 0.008202f
C521 B.n481 VSUBS 0.004583f
C522 B.n482 VSUBS 0.019002f
C523 B.n483 VSUBS 0.007719f
C524 B.n484 VSUBS 0.008202f
C525 B.n485 VSUBS 0.008202f
C526 B.n486 VSUBS 0.008202f
C527 B.n487 VSUBS 0.008202f
C528 B.n488 VSUBS 0.008202f
C529 B.n489 VSUBS 0.008202f
C530 B.n490 VSUBS 0.008202f
C531 B.n491 VSUBS 0.008202f
C532 B.n492 VSUBS 0.008202f
C533 B.n493 VSUBS 0.008202f
C534 B.n494 VSUBS 0.008202f
C535 B.n495 VSUBS 0.008202f
C536 B.n496 VSUBS 0.008202f
C537 B.n497 VSUBS 0.008202f
C538 B.n498 VSUBS 0.008202f
C539 B.n499 VSUBS 0.008202f
C540 B.n500 VSUBS 0.008202f
C541 B.n501 VSUBS 0.008202f
C542 B.n502 VSUBS 0.008202f
C543 B.n503 VSUBS 0.008202f
C544 B.n504 VSUBS 0.008202f
C545 B.n505 VSUBS 0.008202f
C546 B.n506 VSUBS 0.008202f
C547 B.n507 VSUBS 0.008202f
C548 B.n508 VSUBS 0.008202f
C549 B.n509 VSUBS 0.008202f
C550 B.n510 VSUBS 0.008202f
C551 B.n511 VSUBS 0.008202f
C552 B.n512 VSUBS 0.008202f
C553 B.n513 VSUBS 0.008202f
C554 B.n514 VSUBS 0.008202f
C555 B.n515 VSUBS 0.008202f
C556 B.n516 VSUBS 0.008202f
C557 B.n517 VSUBS 0.008202f
C558 B.n518 VSUBS 0.008202f
C559 B.n519 VSUBS 0.008202f
C560 B.n520 VSUBS 0.008202f
C561 B.n521 VSUBS 0.008202f
C562 B.n522 VSUBS 0.008202f
C563 B.n523 VSUBS 0.008202f
C564 B.n524 VSUBS 0.008202f
C565 B.n525 VSUBS 0.008202f
C566 B.n526 VSUBS 0.008202f
C567 B.n527 VSUBS 0.008202f
C568 B.n528 VSUBS 0.008202f
C569 B.n529 VSUBS 0.008202f
C570 B.n530 VSUBS 0.008202f
C571 B.n531 VSUBS 0.008202f
C572 B.n532 VSUBS 0.008202f
C573 B.n533 VSUBS 0.008202f
C574 B.n534 VSUBS 0.008202f
C575 B.n535 VSUBS 0.008202f
C576 B.n536 VSUBS 0.008202f
C577 B.n537 VSUBS 0.008202f
C578 B.n538 VSUBS 0.008202f
C579 B.n539 VSUBS 0.008202f
C580 B.n540 VSUBS 0.008202f
C581 B.n541 VSUBS 0.008202f
C582 B.n542 VSUBS 0.008202f
C583 B.n543 VSUBS 0.008202f
C584 B.n544 VSUBS 0.008202f
C585 B.n545 VSUBS 0.008202f
C586 B.n546 VSUBS 0.008202f
C587 B.n547 VSUBS 0.008202f
C588 B.n548 VSUBS 0.008202f
C589 B.n549 VSUBS 0.019258f
C590 B.n550 VSUBS 0.019258f
C591 B.n551 VSUBS 0.017891f
C592 B.n552 VSUBS 0.008202f
C593 B.n553 VSUBS 0.008202f
C594 B.n554 VSUBS 0.008202f
C595 B.n555 VSUBS 0.008202f
C596 B.n556 VSUBS 0.008202f
C597 B.n557 VSUBS 0.008202f
C598 B.n558 VSUBS 0.008202f
C599 B.n559 VSUBS 0.008202f
C600 B.n560 VSUBS 0.008202f
C601 B.n561 VSUBS 0.008202f
C602 B.n562 VSUBS 0.008202f
C603 B.n563 VSUBS 0.008202f
C604 B.n564 VSUBS 0.008202f
C605 B.n565 VSUBS 0.008202f
C606 B.n566 VSUBS 0.008202f
C607 B.n567 VSUBS 0.008202f
C608 B.n568 VSUBS 0.008202f
C609 B.n569 VSUBS 0.008202f
C610 B.n570 VSUBS 0.008202f
C611 B.n571 VSUBS 0.008202f
C612 B.n572 VSUBS 0.008202f
C613 B.n573 VSUBS 0.008202f
C614 B.n574 VSUBS 0.008202f
C615 B.n575 VSUBS 0.008202f
C616 B.n576 VSUBS 0.008202f
C617 B.n577 VSUBS 0.008202f
C618 B.n578 VSUBS 0.008202f
C619 B.n579 VSUBS 0.008202f
C620 B.n580 VSUBS 0.008202f
C621 B.n581 VSUBS 0.008202f
C622 B.n582 VSUBS 0.008202f
C623 B.n583 VSUBS 0.018571f
C624 VDD2.t4 VSUBS 0.299053f
C625 VDD2.t6 VSUBS 0.299053f
C626 VDD2.n0 VSUBS 2.36812f
C627 VDD2.t0 VSUBS 0.299053f
C628 VDD2.t7 VSUBS 0.299053f
C629 VDD2.n1 VSUBS 2.36812f
C630 VDD2.n2 VSUBS 3.1106f
C631 VDD2.t1 VSUBS 0.299053f
C632 VDD2.t3 VSUBS 0.299053f
C633 VDD2.n3 VSUBS 2.36513f
C634 VDD2.n4 VSUBS 2.99497f
C635 VDD2.t2 VSUBS 0.299053f
C636 VDD2.t5 VSUBS 0.299053f
C637 VDD2.n5 VSUBS 2.36808f
C638 VN.n0 VSUBS 0.057557f
C639 VN.t1 VSUBS 1.18612f
C640 VN.n1 VSUBS 0.481478f
C641 VN.t3 VSUBS 1.20405f
C642 VN.n2 VSUBS 0.454698f
C643 VN.n3 VSUBS 0.235817f
C644 VN.t7 VSUBS 1.18612f
C645 VN.n4 VSUBS 0.471186f
C646 VN.n5 VSUBS 0.013061f
C647 VN.t0 VSUBS 1.18612f
C648 VN.n6 VSUBS 0.468702f
C649 VN.n7 VSUBS 0.044604f
C650 VN.n8 VSUBS 0.057557f
C651 VN.t5 VSUBS 1.18612f
C652 VN.n9 VSUBS 0.481478f
C653 VN.t4 VSUBS 1.18612f
C654 VN.t2 VSUBS 1.20405f
C655 VN.n10 VSUBS 0.454698f
C656 VN.n11 VSUBS 0.235817f
C657 VN.n12 VSUBS 0.471186f
C658 VN.n13 VSUBS 0.013061f
C659 VN.t6 VSUBS 1.18612f
C660 VN.n14 VSUBS 0.468702f
C661 VN.n15 VSUBS 2.42779f
C662 VDD1.t0 VSUBS 0.298954f
C663 VDD1.t7 VSUBS 0.298954f
C664 VDD1.n0 VSUBS 2.36844f
C665 VDD1.t6 VSUBS 0.298954f
C666 VDD1.t2 VSUBS 0.298954f
C667 VDD1.n1 VSUBS 2.36734f
C668 VDD1.t3 VSUBS 0.298954f
C669 VDD1.t1 VSUBS 0.298954f
C670 VDD1.n2 VSUBS 2.36734f
C671 VDD1.n3 VSUBS 3.17098f
C672 VDD1.t4 VSUBS 0.298954f
C673 VDD1.t5 VSUBS 0.298954f
C674 VDD1.n4 VSUBS 2.36434f
C675 VDD1.n5 VSUBS 3.02797f
C676 VTAIL.t7 VSUBS 0.265393f
C677 VTAIL.t6 VSUBS 0.265393f
C678 VTAIL.n0 VSUBS 1.95189f
C679 VTAIL.n1 VSUBS 0.670777f
C680 VTAIL.t0 VSUBS 2.57242f
C681 VTAIL.n2 VSUBS 0.8079f
C682 VTAIL.t15 VSUBS 2.57242f
C683 VTAIL.n3 VSUBS 0.8079f
C684 VTAIL.t9 VSUBS 0.265393f
C685 VTAIL.t12 VSUBS 0.265393f
C686 VTAIL.n4 VSUBS 1.95189f
C687 VTAIL.n5 VSUBS 0.728374f
C688 VTAIL.t13 VSUBS 2.57242f
C689 VTAIL.n6 VSUBS 2.1112f
C690 VTAIL.t5 VSUBS 2.57243f
C691 VTAIL.n7 VSUBS 2.11119f
C692 VTAIL.t2 VSUBS 0.265393f
C693 VTAIL.t3 VSUBS 0.265393f
C694 VTAIL.n8 VSUBS 1.9519f
C695 VTAIL.n9 VSUBS 0.72837f
C696 VTAIL.t1 VSUBS 2.57243f
C697 VTAIL.n10 VSUBS 0.807891f
C698 VTAIL.t10 VSUBS 2.57243f
C699 VTAIL.n11 VSUBS 0.807891f
C700 VTAIL.t14 VSUBS 0.265393f
C701 VTAIL.t11 VSUBS 0.265393f
C702 VTAIL.n12 VSUBS 1.9519f
C703 VTAIL.n13 VSUBS 0.72837f
C704 VTAIL.t8 VSUBS 2.57242f
C705 VTAIL.n14 VSUBS 2.1112f
C706 VTAIL.t4 VSUBS 2.57242f
C707 VTAIL.n15 VSUBS 2.10642f
C708 VP.n0 VSUBS 0.058728f
C709 VP.t5 VSUBS 1.21026f
C710 VP.n1 VSUBS 0.480774f
C711 VP.n2 VSUBS 0.058728f
C712 VP.t2 VSUBS 1.21026f
C713 VP.t3 VSUBS 1.21026f
C714 VP.n3 VSUBS 0.240616f
C715 VP.t0 VSUBS 1.21026f
C716 VP.t7 VSUBS 1.22855f
C717 VP.n4 VSUBS 0.46395f
C718 VP.n5 VSUBS 0.491275f
C719 VP.n6 VSUBS 0.480774f
C720 VP.n7 VSUBS 0.013326f
C721 VP.n8 VSUBS 0.47824f
C722 VP.n9 VSUBS 2.43865f
C723 VP.n10 VSUBS 2.48888f
C724 VP.t1 VSUBS 1.21026f
C725 VP.n11 VSUBS 0.47824f
C726 VP.n12 VSUBS 0.013326f
C727 VP.n13 VSUBS 0.058728f
C728 VP.n14 VSUBS 0.058728f
C729 VP.n15 VSUBS 0.058728f
C730 VP.t4 VSUBS 1.21026f
C731 VP.n16 VSUBS 0.480774f
C732 VP.n17 VSUBS 0.013326f
C733 VP.t6 VSUBS 1.21026f
C734 VP.n18 VSUBS 0.47824f
C735 VP.n19 VSUBS 0.045512f
.ends

