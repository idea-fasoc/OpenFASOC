* NGSPICE file created from diff_pair_sample_1652.ext - technology: sky130A

.subckt diff_pair_sample_1652 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.8381 pd=11.47 as=1.8381 ps=11.47 w=11.14 l=0.75
X1 VDD2.t6 VN.t1 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8381 pd=11.47 as=4.3446 ps=23.06 w=11.14 l=0.75
X2 VTAIL.t8 VN.t2 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=4.3446 pd=23.06 as=1.8381 ps=11.47 w=11.14 l=0.75
X3 VTAIL.t7 VN.t3 VDD2.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=1.8381 pd=11.47 as=1.8381 ps=11.47 w=11.14 l=0.75
X4 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=4.3446 pd=23.06 as=0 ps=0 w=11.14 l=0.75
X5 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=4.3446 pd=23.06 as=0 ps=0 w=11.14 l=0.75
X6 VDD1.t7 VP.t0 VTAIL.t15 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8381 pd=11.47 as=1.8381 ps=11.47 w=11.14 l=0.75
X7 VTAIL.t14 VP.t1 VDD1.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=1.8381 pd=11.47 as=1.8381 ps=11.47 w=11.14 l=0.75
X8 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=4.3446 pd=23.06 as=0 ps=0 w=11.14 l=0.75
X9 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.3446 pd=23.06 as=0 ps=0 w=11.14 l=0.75
X10 VTAIL.t2 VP.t2 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=4.3446 pd=23.06 as=1.8381 ps=11.47 w=11.14 l=0.75
X11 VTAIL.t13 VP.t3 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=1.8381 pd=11.47 as=1.8381 ps=11.47 w=11.14 l=0.75
X12 VDD2.t3 VN.t4 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=1.8381 pd=11.47 as=4.3446 ps=23.06 w=11.14 l=0.75
X13 VTAIL.t9 VN.t5 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=4.3446 pd=23.06 as=1.8381 ps=11.47 w=11.14 l=0.75
X14 VDD1.t3 VP.t4 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=1.8381 pd=11.47 as=4.3446 ps=23.06 w=11.14 l=0.75
X15 VDD2.t1 VN.t6 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8381 pd=11.47 as=1.8381 ps=11.47 w=11.14 l=0.75
X16 VDD1.t2 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8381 pd=11.47 as=4.3446 ps=23.06 w=11.14 l=0.75
X17 VTAIL.t4 VN.t7 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=1.8381 pd=11.47 as=1.8381 ps=11.47 w=11.14 l=0.75
X18 VTAIL.t1 VP.t6 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.3446 pd=23.06 as=1.8381 ps=11.47 w=11.14 l=0.75
X19 VDD1.t0 VP.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.8381 pd=11.47 as=1.8381 ps=11.47 w=11.14 l=0.75
R0 VN.n3 VN.t5 435.01
R1 VN.n13 VN.t4 435.01
R2 VN.n2 VN.t6 410.986
R3 VN.n6 VN.t3 410.986
R4 VN.n8 VN.t1 410.986
R5 VN.n12 VN.t7 410.986
R6 VN.n16 VN.t0 410.986
R7 VN.n18 VN.t2 410.986
R8 VN.n9 VN.n8 161.3
R9 VN.n19 VN.n18 161.3
R10 VN.n17 VN.n10 161.3
R11 VN.n16 VN.n15 161.3
R12 VN.n14 VN.n11 161.3
R13 VN.n7 VN.n0 161.3
R14 VN.n6 VN.n5 161.3
R15 VN.n4 VN.n1 161.3
R16 VN.n14 VN.n13 44.92
R17 VN.n4 VN.n3 44.92
R18 VN VN.n19 42.0251
R19 VN.n8 VN.n7 35.7853
R20 VN.n18 VN.n17 35.7853
R21 VN.n2 VN.n1 24.1005
R22 VN.n6 VN.n1 24.1005
R23 VN.n16 VN.n11 24.1005
R24 VN.n12 VN.n11 24.1005
R25 VN.n3 VN.n2 17.5118
R26 VN.n13 VN.n12 17.5118
R27 VN.n7 VN.n6 12.4157
R28 VN.n17 VN.n16 12.4157
R29 VN.n19 VN.n10 0.189894
R30 VN.n15 VN.n10 0.189894
R31 VN.n15 VN.n14 0.189894
R32 VN.n5 VN.n4 0.189894
R33 VN.n5 VN.n0 0.189894
R34 VN.n9 VN.n0 0.189894
R35 VN VN.n9 0.0516364
R36 VTAIL.n11 VTAIL.t1 49.2471
R37 VTAIL.n10 VTAIL.t10 49.2471
R38 VTAIL.n7 VTAIL.t8 49.2471
R39 VTAIL.n15 VTAIL.t11 49.247
R40 VTAIL.n2 VTAIL.t9 49.247
R41 VTAIL.n3 VTAIL.t12 49.247
R42 VTAIL.n6 VTAIL.t2 49.247
R43 VTAIL.n14 VTAIL.t3 49.247
R44 VTAIL.n13 VTAIL.n12 47.4697
R45 VTAIL.n9 VTAIL.n8 47.4697
R46 VTAIL.n1 VTAIL.n0 47.4695
R47 VTAIL.n5 VTAIL.n4 47.4695
R48 VTAIL.n15 VTAIL.n14 22.9014
R49 VTAIL.n7 VTAIL.n6 22.9014
R50 VTAIL.n0 VTAIL.t5 1.77788
R51 VTAIL.n0 VTAIL.t7 1.77788
R52 VTAIL.n4 VTAIL.t0 1.77788
R53 VTAIL.n4 VTAIL.t14 1.77788
R54 VTAIL.n12 VTAIL.t15 1.77788
R55 VTAIL.n12 VTAIL.t13 1.77788
R56 VTAIL.n8 VTAIL.t6 1.77788
R57 VTAIL.n8 VTAIL.t4 1.77788
R58 VTAIL.n9 VTAIL.n7 0.931535
R59 VTAIL.n10 VTAIL.n9 0.931535
R60 VTAIL.n13 VTAIL.n11 0.931535
R61 VTAIL.n14 VTAIL.n13 0.931535
R62 VTAIL.n6 VTAIL.n5 0.931535
R63 VTAIL.n5 VTAIL.n3 0.931535
R64 VTAIL.n2 VTAIL.n1 0.931535
R65 VTAIL VTAIL.n15 0.873345
R66 VTAIL.n11 VTAIL.n10 0.470328
R67 VTAIL.n3 VTAIL.n2 0.470328
R68 VTAIL VTAIL.n1 0.0586897
R69 VDD2.n2 VDD2.n1 64.5585
R70 VDD2.n2 VDD2.n0 64.5585
R71 VDD2 VDD2.n5 64.5557
R72 VDD2.n4 VDD2.n3 64.1485
R73 VDD2.n4 VDD2.n2 37.5084
R74 VDD2.n5 VDD2.t0 1.77788
R75 VDD2.n5 VDD2.t3 1.77788
R76 VDD2.n3 VDD2.t5 1.77788
R77 VDD2.n3 VDD2.t7 1.77788
R78 VDD2.n1 VDD2.t4 1.77788
R79 VDD2.n1 VDD2.t6 1.77788
R80 VDD2.n0 VDD2.t2 1.77788
R81 VDD2.n0 VDD2.t1 1.77788
R82 VDD2 VDD2.n4 0.524207
R83 B.n644 B.n643 585
R84 B.n268 B.n91 585
R85 B.n267 B.n266 585
R86 B.n265 B.n264 585
R87 B.n263 B.n262 585
R88 B.n261 B.n260 585
R89 B.n259 B.n258 585
R90 B.n257 B.n256 585
R91 B.n255 B.n254 585
R92 B.n253 B.n252 585
R93 B.n251 B.n250 585
R94 B.n249 B.n248 585
R95 B.n247 B.n246 585
R96 B.n245 B.n244 585
R97 B.n243 B.n242 585
R98 B.n241 B.n240 585
R99 B.n239 B.n238 585
R100 B.n237 B.n236 585
R101 B.n235 B.n234 585
R102 B.n233 B.n232 585
R103 B.n231 B.n230 585
R104 B.n229 B.n228 585
R105 B.n227 B.n226 585
R106 B.n225 B.n224 585
R107 B.n223 B.n222 585
R108 B.n221 B.n220 585
R109 B.n219 B.n218 585
R110 B.n217 B.n216 585
R111 B.n215 B.n214 585
R112 B.n213 B.n212 585
R113 B.n211 B.n210 585
R114 B.n209 B.n208 585
R115 B.n207 B.n206 585
R116 B.n205 B.n204 585
R117 B.n203 B.n202 585
R118 B.n201 B.n200 585
R119 B.n199 B.n198 585
R120 B.n197 B.n196 585
R121 B.n195 B.n194 585
R122 B.n192 B.n191 585
R123 B.n190 B.n189 585
R124 B.n188 B.n187 585
R125 B.n186 B.n185 585
R126 B.n184 B.n183 585
R127 B.n182 B.n181 585
R128 B.n180 B.n179 585
R129 B.n178 B.n177 585
R130 B.n176 B.n175 585
R131 B.n174 B.n173 585
R132 B.n171 B.n170 585
R133 B.n169 B.n168 585
R134 B.n167 B.n166 585
R135 B.n165 B.n164 585
R136 B.n163 B.n162 585
R137 B.n161 B.n160 585
R138 B.n159 B.n158 585
R139 B.n157 B.n156 585
R140 B.n155 B.n154 585
R141 B.n153 B.n152 585
R142 B.n151 B.n150 585
R143 B.n149 B.n148 585
R144 B.n147 B.n146 585
R145 B.n145 B.n144 585
R146 B.n143 B.n142 585
R147 B.n141 B.n140 585
R148 B.n139 B.n138 585
R149 B.n137 B.n136 585
R150 B.n135 B.n134 585
R151 B.n133 B.n132 585
R152 B.n131 B.n130 585
R153 B.n129 B.n128 585
R154 B.n127 B.n126 585
R155 B.n125 B.n124 585
R156 B.n123 B.n122 585
R157 B.n121 B.n120 585
R158 B.n119 B.n118 585
R159 B.n117 B.n116 585
R160 B.n115 B.n114 585
R161 B.n113 B.n112 585
R162 B.n111 B.n110 585
R163 B.n109 B.n108 585
R164 B.n107 B.n106 585
R165 B.n105 B.n104 585
R166 B.n103 B.n102 585
R167 B.n101 B.n100 585
R168 B.n99 B.n98 585
R169 B.n97 B.n96 585
R170 B.n46 B.n45 585
R171 B.n642 B.n47 585
R172 B.n647 B.n47 585
R173 B.n641 B.n640 585
R174 B.n640 B.n43 585
R175 B.n639 B.n42 585
R176 B.n653 B.n42 585
R177 B.n638 B.n41 585
R178 B.n654 B.n41 585
R179 B.n637 B.n40 585
R180 B.n655 B.n40 585
R181 B.n636 B.n635 585
R182 B.n635 B.n36 585
R183 B.n634 B.n35 585
R184 B.n661 B.n35 585
R185 B.n633 B.n34 585
R186 B.n662 B.n34 585
R187 B.n632 B.n33 585
R188 B.n663 B.n33 585
R189 B.n631 B.n630 585
R190 B.n630 B.n29 585
R191 B.n629 B.n28 585
R192 B.n669 B.n28 585
R193 B.n628 B.n27 585
R194 B.n670 B.n27 585
R195 B.n627 B.n26 585
R196 B.n671 B.n26 585
R197 B.n626 B.n625 585
R198 B.n625 B.n22 585
R199 B.n624 B.n21 585
R200 B.n677 B.n21 585
R201 B.n623 B.n20 585
R202 B.n678 B.n20 585
R203 B.n622 B.n19 585
R204 B.n679 B.n19 585
R205 B.n621 B.n620 585
R206 B.n620 B.n18 585
R207 B.n619 B.n14 585
R208 B.n685 B.n14 585
R209 B.n618 B.n13 585
R210 B.n686 B.n13 585
R211 B.n617 B.n12 585
R212 B.n687 B.n12 585
R213 B.n616 B.n615 585
R214 B.n615 B.n8 585
R215 B.n614 B.n7 585
R216 B.n693 B.n7 585
R217 B.n613 B.n6 585
R218 B.n694 B.n6 585
R219 B.n612 B.n5 585
R220 B.n695 B.n5 585
R221 B.n611 B.n610 585
R222 B.n610 B.n4 585
R223 B.n609 B.n269 585
R224 B.n609 B.n608 585
R225 B.n599 B.n270 585
R226 B.n271 B.n270 585
R227 B.n601 B.n600 585
R228 B.n602 B.n601 585
R229 B.n598 B.n276 585
R230 B.n276 B.n275 585
R231 B.n597 B.n596 585
R232 B.n596 B.n595 585
R233 B.n278 B.n277 585
R234 B.n588 B.n278 585
R235 B.n587 B.n586 585
R236 B.n589 B.n587 585
R237 B.n585 B.n283 585
R238 B.n283 B.n282 585
R239 B.n584 B.n583 585
R240 B.n583 B.n582 585
R241 B.n285 B.n284 585
R242 B.n286 B.n285 585
R243 B.n575 B.n574 585
R244 B.n576 B.n575 585
R245 B.n573 B.n290 585
R246 B.n294 B.n290 585
R247 B.n572 B.n571 585
R248 B.n571 B.n570 585
R249 B.n292 B.n291 585
R250 B.n293 B.n292 585
R251 B.n563 B.n562 585
R252 B.n564 B.n563 585
R253 B.n561 B.n299 585
R254 B.n299 B.n298 585
R255 B.n560 B.n559 585
R256 B.n559 B.n558 585
R257 B.n301 B.n300 585
R258 B.n302 B.n301 585
R259 B.n551 B.n550 585
R260 B.n552 B.n551 585
R261 B.n549 B.n307 585
R262 B.n307 B.n306 585
R263 B.n548 B.n547 585
R264 B.n547 B.n546 585
R265 B.n309 B.n308 585
R266 B.n310 B.n309 585
R267 B.n539 B.n538 585
R268 B.n540 B.n539 585
R269 B.n313 B.n312 585
R270 B.n366 B.n365 585
R271 B.n367 B.n363 585
R272 B.n363 B.n314 585
R273 B.n369 B.n368 585
R274 B.n371 B.n362 585
R275 B.n374 B.n373 585
R276 B.n375 B.n361 585
R277 B.n377 B.n376 585
R278 B.n379 B.n360 585
R279 B.n382 B.n381 585
R280 B.n383 B.n359 585
R281 B.n385 B.n384 585
R282 B.n387 B.n358 585
R283 B.n390 B.n389 585
R284 B.n391 B.n357 585
R285 B.n393 B.n392 585
R286 B.n395 B.n356 585
R287 B.n398 B.n397 585
R288 B.n399 B.n355 585
R289 B.n401 B.n400 585
R290 B.n403 B.n354 585
R291 B.n406 B.n405 585
R292 B.n407 B.n353 585
R293 B.n409 B.n408 585
R294 B.n411 B.n352 585
R295 B.n414 B.n413 585
R296 B.n415 B.n351 585
R297 B.n417 B.n416 585
R298 B.n419 B.n350 585
R299 B.n422 B.n421 585
R300 B.n423 B.n349 585
R301 B.n425 B.n424 585
R302 B.n427 B.n348 585
R303 B.n430 B.n429 585
R304 B.n431 B.n347 585
R305 B.n433 B.n432 585
R306 B.n435 B.n346 585
R307 B.n438 B.n437 585
R308 B.n439 B.n343 585
R309 B.n442 B.n441 585
R310 B.n444 B.n342 585
R311 B.n447 B.n446 585
R312 B.n448 B.n341 585
R313 B.n450 B.n449 585
R314 B.n452 B.n340 585
R315 B.n455 B.n454 585
R316 B.n456 B.n339 585
R317 B.n458 B.n457 585
R318 B.n460 B.n338 585
R319 B.n463 B.n462 585
R320 B.n464 B.n334 585
R321 B.n466 B.n465 585
R322 B.n468 B.n333 585
R323 B.n471 B.n470 585
R324 B.n472 B.n332 585
R325 B.n474 B.n473 585
R326 B.n476 B.n331 585
R327 B.n479 B.n478 585
R328 B.n480 B.n330 585
R329 B.n482 B.n481 585
R330 B.n484 B.n329 585
R331 B.n487 B.n486 585
R332 B.n488 B.n328 585
R333 B.n490 B.n489 585
R334 B.n492 B.n327 585
R335 B.n495 B.n494 585
R336 B.n496 B.n326 585
R337 B.n498 B.n497 585
R338 B.n500 B.n325 585
R339 B.n503 B.n502 585
R340 B.n504 B.n324 585
R341 B.n506 B.n505 585
R342 B.n508 B.n323 585
R343 B.n511 B.n510 585
R344 B.n512 B.n322 585
R345 B.n514 B.n513 585
R346 B.n516 B.n321 585
R347 B.n519 B.n518 585
R348 B.n520 B.n320 585
R349 B.n522 B.n521 585
R350 B.n524 B.n319 585
R351 B.n527 B.n526 585
R352 B.n528 B.n318 585
R353 B.n530 B.n529 585
R354 B.n532 B.n317 585
R355 B.n533 B.n316 585
R356 B.n536 B.n535 585
R357 B.n537 B.n315 585
R358 B.n315 B.n314 585
R359 B.n542 B.n541 585
R360 B.n541 B.n540 585
R361 B.n543 B.n311 585
R362 B.n311 B.n310 585
R363 B.n545 B.n544 585
R364 B.n546 B.n545 585
R365 B.n305 B.n304 585
R366 B.n306 B.n305 585
R367 B.n554 B.n553 585
R368 B.n553 B.n552 585
R369 B.n555 B.n303 585
R370 B.n303 B.n302 585
R371 B.n557 B.n556 585
R372 B.n558 B.n557 585
R373 B.n297 B.n296 585
R374 B.n298 B.n297 585
R375 B.n566 B.n565 585
R376 B.n565 B.n564 585
R377 B.n567 B.n295 585
R378 B.n295 B.n293 585
R379 B.n569 B.n568 585
R380 B.n570 B.n569 585
R381 B.n289 B.n288 585
R382 B.n294 B.n289 585
R383 B.n578 B.n577 585
R384 B.n577 B.n576 585
R385 B.n579 B.n287 585
R386 B.n287 B.n286 585
R387 B.n581 B.n580 585
R388 B.n582 B.n581 585
R389 B.n281 B.n280 585
R390 B.n282 B.n281 585
R391 B.n591 B.n590 585
R392 B.n590 B.n589 585
R393 B.n592 B.n279 585
R394 B.n588 B.n279 585
R395 B.n594 B.n593 585
R396 B.n595 B.n594 585
R397 B.n274 B.n273 585
R398 B.n275 B.n274 585
R399 B.n604 B.n603 585
R400 B.n603 B.n602 585
R401 B.n605 B.n272 585
R402 B.n272 B.n271 585
R403 B.n607 B.n606 585
R404 B.n608 B.n607 585
R405 B.n2 B.n0 585
R406 B.n4 B.n2 585
R407 B.n3 B.n1 585
R408 B.n694 B.n3 585
R409 B.n692 B.n691 585
R410 B.n693 B.n692 585
R411 B.n690 B.n9 585
R412 B.n9 B.n8 585
R413 B.n689 B.n688 585
R414 B.n688 B.n687 585
R415 B.n11 B.n10 585
R416 B.n686 B.n11 585
R417 B.n684 B.n683 585
R418 B.n685 B.n684 585
R419 B.n682 B.n15 585
R420 B.n18 B.n15 585
R421 B.n681 B.n680 585
R422 B.n680 B.n679 585
R423 B.n17 B.n16 585
R424 B.n678 B.n17 585
R425 B.n676 B.n675 585
R426 B.n677 B.n676 585
R427 B.n674 B.n23 585
R428 B.n23 B.n22 585
R429 B.n673 B.n672 585
R430 B.n672 B.n671 585
R431 B.n25 B.n24 585
R432 B.n670 B.n25 585
R433 B.n668 B.n667 585
R434 B.n669 B.n668 585
R435 B.n666 B.n30 585
R436 B.n30 B.n29 585
R437 B.n665 B.n664 585
R438 B.n664 B.n663 585
R439 B.n32 B.n31 585
R440 B.n662 B.n32 585
R441 B.n660 B.n659 585
R442 B.n661 B.n660 585
R443 B.n658 B.n37 585
R444 B.n37 B.n36 585
R445 B.n657 B.n656 585
R446 B.n656 B.n655 585
R447 B.n39 B.n38 585
R448 B.n654 B.n39 585
R449 B.n652 B.n651 585
R450 B.n653 B.n652 585
R451 B.n650 B.n44 585
R452 B.n44 B.n43 585
R453 B.n649 B.n648 585
R454 B.n648 B.n647 585
R455 B.n697 B.n696 585
R456 B.n696 B.n695 585
R457 B.n335 B.t15 560.356
R458 B.n344 B.t19 560.356
R459 B.n94 B.t12 560.356
R460 B.n92 B.t8 560.356
R461 B.n541 B.n313 478.086
R462 B.n648 B.n46 478.086
R463 B.n539 B.n315 478.086
R464 B.n644 B.n47 478.086
R465 B.n646 B.n645 256.663
R466 B.n646 B.n90 256.663
R467 B.n646 B.n89 256.663
R468 B.n646 B.n88 256.663
R469 B.n646 B.n87 256.663
R470 B.n646 B.n86 256.663
R471 B.n646 B.n85 256.663
R472 B.n646 B.n84 256.663
R473 B.n646 B.n83 256.663
R474 B.n646 B.n82 256.663
R475 B.n646 B.n81 256.663
R476 B.n646 B.n80 256.663
R477 B.n646 B.n79 256.663
R478 B.n646 B.n78 256.663
R479 B.n646 B.n77 256.663
R480 B.n646 B.n76 256.663
R481 B.n646 B.n75 256.663
R482 B.n646 B.n74 256.663
R483 B.n646 B.n73 256.663
R484 B.n646 B.n72 256.663
R485 B.n646 B.n71 256.663
R486 B.n646 B.n70 256.663
R487 B.n646 B.n69 256.663
R488 B.n646 B.n68 256.663
R489 B.n646 B.n67 256.663
R490 B.n646 B.n66 256.663
R491 B.n646 B.n65 256.663
R492 B.n646 B.n64 256.663
R493 B.n646 B.n63 256.663
R494 B.n646 B.n62 256.663
R495 B.n646 B.n61 256.663
R496 B.n646 B.n60 256.663
R497 B.n646 B.n59 256.663
R498 B.n646 B.n58 256.663
R499 B.n646 B.n57 256.663
R500 B.n646 B.n56 256.663
R501 B.n646 B.n55 256.663
R502 B.n646 B.n54 256.663
R503 B.n646 B.n53 256.663
R504 B.n646 B.n52 256.663
R505 B.n646 B.n51 256.663
R506 B.n646 B.n50 256.663
R507 B.n646 B.n49 256.663
R508 B.n646 B.n48 256.663
R509 B.n364 B.n314 256.663
R510 B.n370 B.n314 256.663
R511 B.n372 B.n314 256.663
R512 B.n378 B.n314 256.663
R513 B.n380 B.n314 256.663
R514 B.n386 B.n314 256.663
R515 B.n388 B.n314 256.663
R516 B.n394 B.n314 256.663
R517 B.n396 B.n314 256.663
R518 B.n402 B.n314 256.663
R519 B.n404 B.n314 256.663
R520 B.n410 B.n314 256.663
R521 B.n412 B.n314 256.663
R522 B.n418 B.n314 256.663
R523 B.n420 B.n314 256.663
R524 B.n426 B.n314 256.663
R525 B.n428 B.n314 256.663
R526 B.n434 B.n314 256.663
R527 B.n436 B.n314 256.663
R528 B.n443 B.n314 256.663
R529 B.n445 B.n314 256.663
R530 B.n451 B.n314 256.663
R531 B.n453 B.n314 256.663
R532 B.n459 B.n314 256.663
R533 B.n461 B.n314 256.663
R534 B.n467 B.n314 256.663
R535 B.n469 B.n314 256.663
R536 B.n475 B.n314 256.663
R537 B.n477 B.n314 256.663
R538 B.n483 B.n314 256.663
R539 B.n485 B.n314 256.663
R540 B.n491 B.n314 256.663
R541 B.n493 B.n314 256.663
R542 B.n499 B.n314 256.663
R543 B.n501 B.n314 256.663
R544 B.n507 B.n314 256.663
R545 B.n509 B.n314 256.663
R546 B.n515 B.n314 256.663
R547 B.n517 B.n314 256.663
R548 B.n523 B.n314 256.663
R549 B.n525 B.n314 256.663
R550 B.n531 B.n314 256.663
R551 B.n534 B.n314 256.663
R552 B.n541 B.n311 163.367
R553 B.n545 B.n311 163.367
R554 B.n545 B.n305 163.367
R555 B.n553 B.n305 163.367
R556 B.n553 B.n303 163.367
R557 B.n557 B.n303 163.367
R558 B.n557 B.n297 163.367
R559 B.n565 B.n297 163.367
R560 B.n565 B.n295 163.367
R561 B.n569 B.n295 163.367
R562 B.n569 B.n289 163.367
R563 B.n577 B.n289 163.367
R564 B.n577 B.n287 163.367
R565 B.n581 B.n287 163.367
R566 B.n581 B.n281 163.367
R567 B.n590 B.n281 163.367
R568 B.n590 B.n279 163.367
R569 B.n594 B.n279 163.367
R570 B.n594 B.n274 163.367
R571 B.n603 B.n274 163.367
R572 B.n603 B.n272 163.367
R573 B.n607 B.n272 163.367
R574 B.n607 B.n2 163.367
R575 B.n696 B.n2 163.367
R576 B.n696 B.n3 163.367
R577 B.n692 B.n3 163.367
R578 B.n692 B.n9 163.367
R579 B.n688 B.n9 163.367
R580 B.n688 B.n11 163.367
R581 B.n684 B.n11 163.367
R582 B.n684 B.n15 163.367
R583 B.n680 B.n15 163.367
R584 B.n680 B.n17 163.367
R585 B.n676 B.n17 163.367
R586 B.n676 B.n23 163.367
R587 B.n672 B.n23 163.367
R588 B.n672 B.n25 163.367
R589 B.n668 B.n25 163.367
R590 B.n668 B.n30 163.367
R591 B.n664 B.n30 163.367
R592 B.n664 B.n32 163.367
R593 B.n660 B.n32 163.367
R594 B.n660 B.n37 163.367
R595 B.n656 B.n37 163.367
R596 B.n656 B.n39 163.367
R597 B.n652 B.n39 163.367
R598 B.n652 B.n44 163.367
R599 B.n648 B.n44 163.367
R600 B.n365 B.n363 163.367
R601 B.n369 B.n363 163.367
R602 B.n373 B.n371 163.367
R603 B.n377 B.n361 163.367
R604 B.n381 B.n379 163.367
R605 B.n385 B.n359 163.367
R606 B.n389 B.n387 163.367
R607 B.n393 B.n357 163.367
R608 B.n397 B.n395 163.367
R609 B.n401 B.n355 163.367
R610 B.n405 B.n403 163.367
R611 B.n409 B.n353 163.367
R612 B.n413 B.n411 163.367
R613 B.n417 B.n351 163.367
R614 B.n421 B.n419 163.367
R615 B.n425 B.n349 163.367
R616 B.n429 B.n427 163.367
R617 B.n433 B.n347 163.367
R618 B.n437 B.n435 163.367
R619 B.n442 B.n343 163.367
R620 B.n446 B.n444 163.367
R621 B.n450 B.n341 163.367
R622 B.n454 B.n452 163.367
R623 B.n458 B.n339 163.367
R624 B.n462 B.n460 163.367
R625 B.n466 B.n334 163.367
R626 B.n470 B.n468 163.367
R627 B.n474 B.n332 163.367
R628 B.n478 B.n476 163.367
R629 B.n482 B.n330 163.367
R630 B.n486 B.n484 163.367
R631 B.n490 B.n328 163.367
R632 B.n494 B.n492 163.367
R633 B.n498 B.n326 163.367
R634 B.n502 B.n500 163.367
R635 B.n506 B.n324 163.367
R636 B.n510 B.n508 163.367
R637 B.n514 B.n322 163.367
R638 B.n518 B.n516 163.367
R639 B.n522 B.n320 163.367
R640 B.n526 B.n524 163.367
R641 B.n530 B.n318 163.367
R642 B.n533 B.n532 163.367
R643 B.n535 B.n315 163.367
R644 B.n539 B.n309 163.367
R645 B.n547 B.n309 163.367
R646 B.n547 B.n307 163.367
R647 B.n551 B.n307 163.367
R648 B.n551 B.n301 163.367
R649 B.n559 B.n301 163.367
R650 B.n559 B.n299 163.367
R651 B.n563 B.n299 163.367
R652 B.n563 B.n292 163.367
R653 B.n571 B.n292 163.367
R654 B.n571 B.n290 163.367
R655 B.n575 B.n290 163.367
R656 B.n575 B.n285 163.367
R657 B.n583 B.n285 163.367
R658 B.n583 B.n283 163.367
R659 B.n587 B.n283 163.367
R660 B.n587 B.n278 163.367
R661 B.n596 B.n278 163.367
R662 B.n596 B.n276 163.367
R663 B.n601 B.n276 163.367
R664 B.n601 B.n270 163.367
R665 B.n609 B.n270 163.367
R666 B.n610 B.n609 163.367
R667 B.n610 B.n5 163.367
R668 B.n6 B.n5 163.367
R669 B.n7 B.n6 163.367
R670 B.n615 B.n7 163.367
R671 B.n615 B.n12 163.367
R672 B.n13 B.n12 163.367
R673 B.n14 B.n13 163.367
R674 B.n620 B.n14 163.367
R675 B.n620 B.n19 163.367
R676 B.n20 B.n19 163.367
R677 B.n21 B.n20 163.367
R678 B.n625 B.n21 163.367
R679 B.n625 B.n26 163.367
R680 B.n27 B.n26 163.367
R681 B.n28 B.n27 163.367
R682 B.n630 B.n28 163.367
R683 B.n630 B.n33 163.367
R684 B.n34 B.n33 163.367
R685 B.n35 B.n34 163.367
R686 B.n635 B.n35 163.367
R687 B.n635 B.n40 163.367
R688 B.n41 B.n40 163.367
R689 B.n42 B.n41 163.367
R690 B.n640 B.n42 163.367
R691 B.n640 B.n47 163.367
R692 B.n98 B.n97 163.367
R693 B.n102 B.n101 163.367
R694 B.n106 B.n105 163.367
R695 B.n110 B.n109 163.367
R696 B.n114 B.n113 163.367
R697 B.n118 B.n117 163.367
R698 B.n122 B.n121 163.367
R699 B.n126 B.n125 163.367
R700 B.n130 B.n129 163.367
R701 B.n134 B.n133 163.367
R702 B.n138 B.n137 163.367
R703 B.n142 B.n141 163.367
R704 B.n146 B.n145 163.367
R705 B.n150 B.n149 163.367
R706 B.n154 B.n153 163.367
R707 B.n158 B.n157 163.367
R708 B.n162 B.n161 163.367
R709 B.n166 B.n165 163.367
R710 B.n170 B.n169 163.367
R711 B.n175 B.n174 163.367
R712 B.n179 B.n178 163.367
R713 B.n183 B.n182 163.367
R714 B.n187 B.n186 163.367
R715 B.n191 B.n190 163.367
R716 B.n196 B.n195 163.367
R717 B.n200 B.n199 163.367
R718 B.n204 B.n203 163.367
R719 B.n208 B.n207 163.367
R720 B.n212 B.n211 163.367
R721 B.n216 B.n215 163.367
R722 B.n220 B.n219 163.367
R723 B.n224 B.n223 163.367
R724 B.n228 B.n227 163.367
R725 B.n232 B.n231 163.367
R726 B.n236 B.n235 163.367
R727 B.n240 B.n239 163.367
R728 B.n244 B.n243 163.367
R729 B.n248 B.n247 163.367
R730 B.n252 B.n251 163.367
R731 B.n256 B.n255 163.367
R732 B.n260 B.n259 163.367
R733 B.n264 B.n263 163.367
R734 B.n266 B.n91 163.367
R735 B.n335 B.t18 93.9037
R736 B.n92 B.t10 93.9037
R737 B.n344 B.t21 93.8899
R738 B.n94 B.t13 93.8899
R739 B.n540 B.n314 82.4251
R740 B.n647 B.n646 82.4251
R741 B.n336 B.t17 72.9582
R742 B.n93 B.t11 72.9582
R743 B.n345 B.t20 72.9445
R744 B.n95 B.t14 72.9445
R745 B.n364 B.n313 71.676
R746 B.n370 B.n369 71.676
R747 B.n373 B.n372 71.676
R748 B.n378 B.n377 71.676
R749 B.n381 B.n380 71.676
R750 B.n386 B.n385 71.676
R751 B.n389 B.n388 71.676
R752 B.n394 B.n393 71.676
R753 B.n397 B.n396 71.676
R754 B.n402 B.n401 71.676
R755 B.n405 B.n404 71.676
R756 B.n410 B.n409 71.676
R757 B.n413 B.n412 71.676
R758 B.n418 B.n417 71.676
R759 B.n421 B.n420 71.676
R760 B.n426 B.n425 71.676
R761 B.n429 B.n428 71.676
R762 B.n434 B.n433 71.676
R763 B.n437 B.n436 71.676
R764 B.n443 B.n442 71.676
R765 B.n446 B.n445 71.676
R766 B.n451 B.n450 71.676
R767 B.n454 B.n453 71.676
R768 B.n459 B.n458 71.676
R769 B.n462 B.n461 71.676
R770 B.n467 B.n466 71.676
R771 B.n470 B.n469 71.676
R772 B.n475 B.n474 71.676
R773 B.n478 B.n477 71.676
R774 B.n483 B.n482 71.676
R775 B.n486 B.n485 71.676
R776 B.n491 B.n490 71.676
R777 B.n494 B.n493 71.676
R778 B.n499 B.n498 71.676
R779 B.n502 B.n501 71.676
R780 B.n507 B.n506 71.676
R781 B.n510 B.n509 71.676
R782 B.n515 B.n514 71.676
R783 B.n518 B.n517 71.676
R784 B.n523 B.n522 71.676
R785 B.n526 B.n525 71.676
R786 B.n531 B.n530 71.676
R787 B.n534 B.n533 71.676
R788 B.n48 B.n46 71.676
R789 B.n98 B.n49 71.676
R790 B.n102 B.n50 71.676
R791 B.n106 B.n51 71.676
R792 B.n110 B.n52 71.676
R793 B.n114 B.n53 71.676
R794 B.n118 B.n54 71.676
R795 B.n122 B.n55 71.676
R796 B.n126 B.n56 71.676
R797 B.n130 B.n57 71.676
R798 B.n134 B.n58 71.676
R799 B.n138 B.n59 71.676
R800 B.n142 B.n60 71.676
R801 B.n146 B.n61 71.676
R802 B.n150 B.n62 71.676
R803 B.n154 B.n63 71.676
R804 B.n158 B.n64 71.676
R805 B.n162 B.n65 71.676
R806 B.n166 B.n66 71.676
R807 B.n170 B.n67 71.676
R808 B.n175 B.n68 71.676
R809 B.n179 B.n69 71.676
R810 B.n183 B.n70 71.676
R811 B.n187 B.n71 71.676
R812 B.n191 B.n72 71.676
R813 B.n196 B.n73 71.676
R814 B.n200 B.n74 71.676
R815 B.n204 B.n75 71.676
R816 B.n208 B.n76 71.676
R817 B.n212 B.n77 71.676
R818 B.n216 B.n78 71.676
R819 B.n220 B.n79 71.676
R820 B.n224 B.n80 71.676
R821 B.n228 B.n81 71.676
R822 B.n232 B.n82 71.676
R823 B.n236 B.n83 71.676
R824 B.n240 B.n84 71.676
R825 B.n244 B.n85 71.676
R826 B.n248 B.n86 71.676
R827 B.n252 B.n87 71.676
R828 B.n256 B.n88 71.676
R829 B.n260 B.n89 71.676
R830 B.n264 B.n90 71.676
R831 B.n645 B.n91 71.676
R832 B.n645 B.n644 71.676
R833 B.n266 B.n90 71.676
R834 B.n263 B.n89 71.676
R835 B.n259 B.n88 71.676
R836 B.n255 B.n87 71.676
R837 B.n251 B.n86 71.676
R838 B.n247 B.n85 71.676
R839 B.n243 B.n84 71.676
R840 B.n239 B.n83 71.676
R841 B.n235 B.n82 71.676
R842 B.n231 B.n81 71.676
R843 B.n227 B.n80 71.676
R844 B.n223 B.n79 71.676
R845 B.n219 B.n78 71.676
R846 B.n215 B.n77 71.676
R847 B.n211 B.n76 71.676
R848 B.n207 B.n75 71.676
R849 B.n203 B.n74 71.676
R850 B.n199 B.n73 71.676
R851 B.n195 B.n72 71.676
R852 B.n190 B.n71 71.676
R853 B.n186 B.n70 71.676
R854 B.n182 B.n69 71.676
R855 B.n178 B.n68 71.676
R856 B.n174 B.n67 71.676
R857 B.n169 B.n66 71.676
R858 B.n165 B.n65 71.676
R859 B.n161 B.n64 71.676
R860 B.n157 B.n63 71.676
R861 B.n153 B.n62 71.676
R862 B.n149 B.n61 71.676
R863 B.n145 B.n60 71.676
R864 B.n141 B.n59 71.676
R865 B.n137 B.n58 71.676
R866 B.n133 B.n57 71.676
R867 B.n129 B.n56 71.676
R868 B.n125 B.n55 71.676
R869 B.n121 B.n54 71.676
R870 B.n117 B.n53 71.676
R871 B.n113 B.n52 71.676
R872 B.n109 B.n51 71.676
R873 B.n105 B.n50 71.676
R874 B.n101 B.n49 71.676
R875 B.n97 B.n48 71.676
R876 B.n365 B.n364 71.676
R877 B.n371 B.n370 71.676
R878 B.n372 B.n361 71.676
R879 B.n379 B.n378 71.676
R880 B.n380 B.n359 71.676
R881 B.n387 B.n386 71.676
R882 B.n388 B.n357 71.676
R883 B.n395 B.n394 71.676
R884 B.n396 B.n355 71.676
R885 B.n403 B.n402 71.676
R886 B.n404 B.n353 71.676
R887 B.n411 B.n410 71.676
R888 B.n412 B.n351 71.676
R889 B.n419 B.n418 71.676
R890 B.n420 B.n349 71.676
R891 B.n427 B.n426 71.676
R892 B.n428 B.n347 71.676
R893 B.n435 B.n434 71.676
R894 B.n436 B.n343 71.676
R895 B.n444 B.n443 71.676
R896 B.n445 B.n341 71.676
R897 B.n452 B.n451 71.676
R898 B.n453 B.n339 71.676
R899 B.n460 B.n459 71.676
R900 B.n461 B.n334 71.676
R901 B.n468 B.n467 71.676
R902 B.n469 B.n332 71.676
R903 B.n476 B.n475 71.676
R904 B.n477 B.n330 71.676
R905 B.n484 B.n483 71.676
R906 B.n485 B.n328 71.676
R907 B.n492 B.n491 71.676
R908 B.n493 B.n326 71.676
R909 B.n500 B.n499 71.676
R910 B.n501 B.n324 71.676
R911 B.n508 B.n507 71.676
R912 B.n509 B.n322 71.676
R913 B.n516 B.n515 71.676
R914 B.n517 B.n320 71.676
R915 B.n524 B.n523 71.676
R916 B.n525 B.n318 71.676
R917 B.n532 B.n531 71.676
R918 B.n535 B.n534 71.676
R919 B.n337 B.n336 59.5399
R920 B.n440 B.n345 59.5399
R921 B.n172 B.n95 59.5399
R922 B.n193 B.n93 59.5399
R923 B.n540 B.n310 45.5686
R924 B.n546 B.n310 45.5686
R925 B.n546 B.n306 45.5686
R926 B.n552 B.n306 45.5686
R927 B.n558 B.n302 45.5686
R928 B.n558 B.n298 45.5686
R929 B.n564 B.n298 45.5686
R930 B.n564 B.n293 45.5686
R931 B.n570 B.n293 45.5686
R932 B.n570 B.n294 45.5686
R933 B.n576 B.n286 45.5686
R934 B.n582 B.n286 45.5686
R935 B.n589 B.n282 45.5686
R936 B.n589 B.n588 45.5686
R937 B.n595 B.n275 45.5686
R938 B.n602 B.n275 45.5686
R939 B.n608 B.n271 45.5686
R940 B.n608 B.n4 45.5686
R941 B.n695 B.n4 45.5686
R942 B.n695 B.n694 45.5686
R943 B.n694 B.n693 45.5686
R944 B.n693 B.n8 45.5686
R945 B.n687 B.n686 45.5686
R946 B.n686 B.n685 45.5686
R947 B.n679 B.n18 45.5686
R948 B.n679 B.n678 45.5686
R949 B.n677 B.n22 45.5686
R950 B.n671 B.n22 45.5686
R951 B.n670 B.n669 45.5686
R952 B.n669 B.n29 45.5686
R953 B.n663 B.n29 45.5686
R954 B.n663 B.n662 45.5686
R955 B.n662 B.n661 45.5686
R956 B.n661 B.n36 45.5686
R957 B.n655 B.n654 45.5686
R958 B.n654 B.n653 45.5686
R959 B.n653 B.n43 45.5686
R960 B.n647 B.n43 45.5686
R961 B.n552 B.t16 40.8777
R962 B.n655 B.t9 40.8777
R963 B.n602 B.t6 36.857
R964 B.n687 B.t1 36.857
R965 B.n576 B.t2 32.8363
R966 B.n671 B.t3 32.8363
R967 B.n649 B.n45 31.0639
R968 B.n643 B.n642 31.0639
R969 B.n538 B.n537 31.0639
R970 B.n542 B.n312 31.0639
R971 B.n588 B.t4 28.8156
R972 B.n18 B.t5 28.8156
R973 B.t0 B.n282 24.7949
R974 B.n678 B.t7 24.7949
R975 B.n336 B.n335 20.946
R976 B.n345 B.n344 20.946
R977 B.n95 B.n94 20.946
R978 B.n93 B.n92 20.946
R979 B.n582 B.t0 20.7742
R980 B.t7 B.n677 20.7742
R981 B B.n697 18.0485
R982 B.n595 B.t4 16.7535
R983 B.n685 B.t5 16.7535
R984 B.n294 B.t2 12.7328
R985 B.t3 B.n670 12.7328
R986 B.n96 B.n45 10.6151
R987 B.n99 B.n96 10.6151
R988 B.n100 B.n99 10.6151
R989 B.n103 B.n100 10.6151
R990 B.n104 B.n103 10.6151
R991 B.n107 B.n104 10.6151
R992 B.n108 B.n107 10.6151
R993 B.n111 B.n108 10.6151
R994 B.n112 B.n111 10.6151
R995 B.n115 B.n112 10.6151
R996 B.n116 B.n115 10.6151
R997 B.n119 B.n116 10.6151
R998 B.n120 B.n119 10.6151
R999 B.n123 B.n120 10.6151
R1000 B.n124 B.n123 10.6151
R1001 B.n127 B.n124 10.6151
R1002 B.n128 B.n127 10.6151
R1003 B.n131 B.n128 10.6151
R1004 B.n132 B.n131 10.6151
R1005 B.n135 B.n132 10.6151
R1006 B.n136 B.n135 10.6151
R1007 B.n139 B.n136 10.6151
R1008 B.n140 B.n139 10.6151
R1009 B.n143 B.n140 10.6151
R1010 B.n144 B.n143 10.6151
R1011 B.n147 B.n144 10.6151
R1012 B.n148 B.n147 10.6151
R1013 B.n151 B.n148 10.6151
R1014 B.n152 B.n151 10.6151
R1015 B.n155 B.n152 10.6151
R1016 B.n156 B.n155 10.6151
R1017 B.n159 B.n156 10.6151
R1018 B.n160 B.n159 10.6151
R1019 B.n163 B.n160 10.6151
R1020 B.n164 B.n163 10.6151
R1021 B.n167 B.n164 10.6151
R1022 B.n168 B.n167 10.6151
R1023 B.n171 B.n168 10.6151
R1024 B.n176 B.n173 10.6151
R1025 B.n177 B.n176 10.6151
R1026 B.n180 B.n177 10.6151
R1027 B.n181 B.n180 10.6151
R1028 B.n184 B.n181 10.6151
R1029 B.n185 B.n184 10.6151
R1030 B.n188 B.n185 10.6151
R1031 B.n189 B.n188 10.6151
R1032 B.n192 B.n189 10.6151
R1033 B.n197 B.n194 10.6151
R1034 B.n198 B.n197 10.6151
R1035 B.n201 B.n198 10.6151
R1036 B.n202 B.n201 10.6151
R1037 B.n205 B.n202 10.6151
R1038 B.n206 B.n205 10.6151
R1039 B.n209 B.n206 10.6151
R1040 B.n210 B.n209 10.6151
R1041 B.n213 B.n210 10.6151
R1042 B.n214 B.n213 10.6151
R1043 B.n217 B.n214 10.6151
R1044 B.n218 B.n217 10.6151
R1045 B.n221 B.n218 10.6151
R1046 B.n222 B.n221 10.6151
R1047 B.n225 B.n222 10.6151
R1048 B.n226 B.n225 10.6151
R1049 B.n229 B.n226 10.6151
R1050 B.n230 B.n229 10.6151
R1051 B.n233 B.n230 10.6151
R1052 B.n234 B.n233 10.6151
R1053 B.n237 B.n234 10.6151
R1054 B.n238 B.n237 10.6151
R1055 B.n241 B.n238 10.6151
R1056 B.n242 B.n241 10.6151
R1057 B.n245 B.n242 10.6151
R1058 B.n246 B.n245 10.6151
R1059 B.n249 B.n246 10.6151
R1060 B.n250 B.n249 10.6151
R1061 B.n253 B.n250 10.6151
R1062 B.n254 B.n253 10.6151
R1063 B.n257 B.n254 10.6151
R1064 B.n258 B.n257 10.6151
R1065 B.n261 B.n258 10.6151
R1066 B.n262 B.n261 10.6151
R1067 B.n265 B.n262 10.6151
R1068 B.n267 B.n265 10.6151
R1069 B.n268 B.n267 10.6151
R1070 B.n643 B.n268 10.6151
R1071 B.n538 B.n308 10.6151
R1072 B.n548 B.n308 10.6151
R1073 B.n549 B.n548 10.6151
R1074 B.n550 B.n549 10.6151
R1075 B.n550 B.n300 10.6151
R1076 B.n560 B.n300 10.6151
R1077 B.n561 B.n560 10.6151
R1078 B.n562 B.n561 10.6151
R1079 B.n562 B.n291 10.6151
R1080 B.n572 B.n291 10.6151
R1081 B.n573 B.n572 10.6151
R1082 B.n574 B.n573 10.6151
R1083 B.n574 B.n284 10.6151
R1084 B.n584 B.n284 10.6151
R1085 B.n585 B.n584 10.6151
R1086 B.n586 B.n585 10.6151
R1087 B.n586 B.n277 10.6151
R1088 B.n597 B.n277 10.6151
R1089 B.n598 B.n597 10.6151
R1090 B.n600 B.n598 10.6151
R1091 B.n600 B.n599 10.6151
R1092 B.n599 B.n269 10.6151
R1093 B.n611 B.n269 10.6151
R1094 B.n612 B.n611 10.6151
R1095 B.n613 B.n612 10.6151
R1096 B.n614 B.n613 10.6151
R1097 B.n616 B.n614 10.6151
R1098 B.n617 B.n616 10.6151
R1099 B.n618 B.n617 10.6151
R1100 B.n619 B.n618 10.6151
R1101 B.n621 B.n619 10.6151
R1102 B.n622 B.n621 10.6151
R1103 B.n623 B.n622 10.6151
R1104 B.n624 B.n623 10.6151
R1105 B.n626 B.n624 10.6151
R1106 B.n627 B.n626 10.6151
R1107 B.n628 B.n627 10.6151
R1108 B.n629 B.n628 10.6151
R1109 B.n631 B.n629 10.6151
R1110 B.n632 B.n631 10.6151
R1111 B.n633 B.n632 10.6151
R1112 B.n634 B.n633 10.6151
R1113 B.n636 B.n634 10.6151
R1114 B.n637 B.n636 10.6151
R1115 B.n638 B.n637 10.6151
R1116 B.n639 B.n638 10.6151
R1117 B.n641 B.n639 10.6151
R1118 B.n642 B.n641 10.6151
R1119 B.n366 B.n312 10.6151
R1120 B.n367 B.n366 10.6151
R1121 B.n368 B.n367 10.6151
R1122 B.n368 B.n362 10.6151
R1123 B.n374 B.n362 10.6151
R1124 B.n375 B.n374 10.6151
R1125 B.n376 B.n375 10.6151
R1126 B.n376 B.n360 10.6151
R1127 B.n382 B.n360 10.6151
R1128 B.n383 B.n382 10.6151
R1129 B.n384 B.n383 10.6151
R1130 B.n384 B.n358 10.6151
R1131 B.n390 B.n358 10.6151
R1132 B.n391 B.n390 10.6151
R1133 B.n392 B.n391 10.6151
R1134 B.n392 B.n356 10.6151
R1135 B.n398 B.n356 10.6151
R1136 B.n399 B.n398 10.6151
R1137 B.n400 B.n399 10.6151
R1138 B.n400 B.n354 10.6151
R1139 B.n406 B.n354 10.6151
R1140 B.n407 B.n406 10.6151
R1141 B.n408 B.n407 10.6151
R1142 B.n408 B.n352 10.6151
R1143 B.n414 B.n352 10.6151
R1144 B.n415 B.n414 10.6151
R1145 B.n416 B.n415 10.6151
R1146 B.n416 B.n350 10.6151
R1147 B.n422 B.n350 10.6151
R1148 B.n423 B.n422 10.6151
R1149 B.n424 B.n423 10.6151
R1150 B.n424 B.n348 10.6151
R1151 B.n430 B.n348 10.6151
R1152 B.n431 B.n430 10.6151
R1153 B.n432 B.n431 10.6151
R1154 B.n432 B.n346 10.6151
R1155 B.n438 B.n346 10.6151
R1156 B.n439 B.n438 10.6151
R1157 B.n441 B.n342 10.6151
R1158 B.n447 B.n342 10.6151
R1159 B.n448 B.n447 10.6151
R1160 B.n449 B.n448 10.6151
R1161 B.n449 B.n340 10.6151
R1162 B.n455 B.n340 10.6151
R1163 B.n456 B.n455 10.6151
R1164 B.n457 B.n456 10.6151
R1165 B.n457 B.n338 10.6151
R1166 B.n464 B.n463 10.6151
R1167 B.n465 B.n464 10.6151
R1168 B.n465 B.n333 10.6151
R1169 B.n471 B.n333 10.6151
R1170 B.n472 B.n471 10.6151
R1171 B.n473 B.n472 10.6151
R1172 B.n473 B.n331 10.6151
R1173 B.n479 B.n331 10.6151
R1174 B.n480 B.n479 10.6151
R1175 B.n481 B.n480 10.6151
R1176 B.n481 B.n329 10.6151
R1177 B.n487 B.n329 10.6151
R1178 B.n488 B.n487 10.6151
R1179 B.n489 B.n488 10.6151
R1180 B.n489 B.n327 10.6151
R1181 B.n495 B.n327 10.6151
R1182 B.n496 B.n495 10.6151
R1183 B.n497 B.n496 10.6151
R1184 B.n497 B.n325 10.6151
R1185 B.n503 B.n325 10.6151
R1186 B.n504 B.n503 10.6151
R1187 B.n505 B.n504 10.6151
R1188 B.n505 B.n323 10.6151
R1189 B.n511 B.n323 10.6151
R1190 B.n512 B.n511 10.6151
R1191 B.n513 B.n512 10.6151
R1192 B.n513 B.n321 10.6151
R1193 B.n519 B.n321 10.6151
R1194 B.n520 B.n519 10.6151
R1195 B.n521 B.n520 10.6151
R1196 B.n521 B.n319 10.6151
R1197 B.n527 B.n319 10.6151
R1198 B.n528 B.n527 10.6151
R1199 B.n529 B.n528 10.6151
R1200 B.n529 B.n317 10.6151
R1201 B.n317 B.n316 10.6151
R1202 B.n536 B.n316 10.6151
R1203 B.n537 B.n536 10.6151
R1204 B.n543 B.n542 10.6151
R1205 B.n544 B.n543 10.6151
R1206 B.n544 B.n304 10.6151
R1207 B.n554 B.n304 10.6151
R1208 B.n555 B.n554 10.6151
R1209 B.n556 B.n555 10.6151
R1210 B.n556 B.n296 10.6151
R1211 B.n566 B.n296 10.6151
R1212 B.n567 B.n566 10.6151
R1213 B.n568 B.n567 10.6151
R1214 B.n568 B.n288 10.6151
R1215 B.n578 B.n288 10.6151
R1216 B.n579 B.n578 10.6151
R1217 B.n580 B.n579 10.6151
R1218 B.n580 B.n280 10.6151
R1219 B.n591 B.n280 10.6151
R1220 B.n592 B.n591 10.6151
R1221 B.n593 B.n592 10.6151
R1222 B.n593 B.n273 10.6151
R1223 B.n604 B.n273 10.6151
R1224 B.n605 B.n604 10.6151
R1225 B.n606 B.n605 10.6151
R1226 B.n606 B.n0 10.6151
R1227 B.n691 B.n1 10.6151
R1228 B.n691 B.n690 10.6151
R1229 B.n690 B.n689 10.6151
R1230 B.n689 B.n10 10.6151
R1231 B.n683 B.n10 10.6151
R1232 B.n683 B.n682 10.6151
R1233 B.n682 B.n681 10.6151
R1234 B.n681 B.n16 10.6151
R1235 B.n675 B.n16 10.6151
R1236 B.n675 B.n674 10.6151
R1237 B.n674 B.n673 10.6151
R1238 B.n673 B.n24 10.6151
R1239 B.n667 B.n24 10.6151
R1240 B.n667 B.n666 10.6151
R1241 B.n666 B.n665 10.6151
R1242 B.n665 B.n31 10.6151
R1243 B.n659 B.n31 10.6151
R1244 B.n659 B.n658 10.6151
R1245 B.n658 B.n657 10.6151
R1246 B.n657 B.n38 10.6151
R1247 B.n651 B.n38 10.6151
R1248 B.n651 B.n650 10.6151
R1249 B.n650 B.n649 10.6151
R1250 B.n172 B.n171 9.36635
R1251 B.n194 B.n193 9.36635
R1252 B.n440 B.n439 9.36635
R1253 B.n463 B.n337 9.36635
R1254 B.t6 B.n271 8.71204
R1255 B.t1 B.n8 8.71204
R1256 B.t16 B.n302 4.69133
R1257 B.t9 B.n36 4.69133
R1258 B.n697 B.n0 2.81026
R1259 B.n697 B.n1 2.81026
R1260 B.n173 B.n172 1.24928
R1261 B.n193 B.n192 1.24928
R1262 B.n441 B.n440 1.24928
R1263 B.n338 B.n337 1.24928
R1264 VP.n6 VP.t6 435.01
R1265 VP.n14 VP.t2 410.986
R1266 VP.n16 VP.t7 410.986
R1267 VP.n20 VP.t1 410.986
R1268 VP.n22 VP.t4 410.986
R1269 VP.n11 VP.t5 410.986
R1270 VP.n9 VP.t3 410.986
R1271 VP.n5 VP.t0 410.986
R1272 VP.n23 VP.n22 161.3
R1273 VP.n8 VP.n7 161.3
R1274 VP.n9 VP.n4 161.3
R1275 VP.n10 VP.n3 161.3
R1276 VP.n12 VP.n11 161.3
R1277 VP.n21 VP.n0 161.3
R1278 VP.n20 VP.n19 161.3
R1279 VP.n18 VP.n1 161.3
R1280 VP.n17 VP.n16 161.3
R1281 VP.n15 VP.n2 161.3
R1282 VP.n14 VP.n13 161.3
R1283 VP.n7 VP.n6 44.92
R1284 VP.n13 VP.n12 41.6444
R1285 VP.n15 VP.n14 35.7853
R1286 VP.n22 VP.n21 35.7853
R1287 VP.n11 VP.n10 35.7853
R1288 VP.n16 VP.n1 24.1005
R1289 VP.n20 VP.n1 24.1005
R1290 VP.n8 VP.n5 24.1005
R1291 VP.n9 VP.n8 24.1005
R1292 VP.n6 VP.n5 17.5118
R1293 VP.n16 VP.n15 12.4157
R1294 VP.n21 VP.n20 12.4157
R1295 VP.n10 VP.n9 12.4157
R1296 VP.n7 VP.n4 0.189894
R1297 VP.n4 VP.n3 0.189894
R1298 VP.n12 VP.n3 0.189894
R1299 VP.n13 VP.n2 0.189894
R1300 VP.n17 VP.n2 0.189894
R1301 VP.n18 VP.n17 0.189894
R1302 VP.n19 VP.n18 0.189894
R1303 VP.n19 VP.n0 0.189894
R1304 VP.n23 VP.n0 0.189894
R1305 VP VP.n23 0.0516364
R1306 VDD1 VDD1.n0 64.6722
R1307 VDD1.n3 VDD1.n2 64.5585
R1308 VDD1.n3 VDD1.n1 64.5585
R1309 VDD1.n5 VDD1.n4 64.1484
R1310 VDD1.n5 VDD1.n3 38.0914
R1311 VDD1.n4 VDD1.t4 1.77788
R1312 VDD1.n4 VDD1.t2 1.77788
R1313 VDD1.n0 VDD1.t1 1.77788
R1314 VDD1.n0 VDD1.t7 1.77788
R1315 VDD1.n2 VDD1.t6 1.77788
R1316 VDD1.n2 VDD1.t3 1.77788
R1317 VDD1.n1 VDD1.t5 1.77788
R1318 VDD1.n1 VDD1.t0 1.77788
R1319 VDD1 VDD1.n5 0.407828
C0 VN VDD2 5.325799f
C1 VTAIL VP 5.15136f
C2 VDD1 VP 5.49976f
C3 VN VP 5.24185f
C4 VDD1 VTAIL 10.1338f
C5 VDD2 VP 0.322204f
C6 VN VTAIL 5.13725f
C7 VDD2 VTAIL 10.175799f
C8 VN VDD1 0.147776f
C9 VDD2 VDD1 0.849097f
C10 VDD2 B 3.468691f
C11 VDD1 B 3.707688f
C12 VTAIL B 8.507095f
C13 VN B 8.63903f
C14 VP B 6.770648f
C15 VDD1.t1 B 0.237545f
C16 VDD1.t7 B 0.237545f
C17 VDD1.n0 B 2.11166f
C18 VDD1.t5 B 0.237545f
C19 VDD1.t0 B 0.237545f
C20 VDD1.n1 B 2.11098f
C21 VDD1.t6 B 0.237545f
C22 VDD1.t3 B 0.237545f
C23 VDD1.n2 B 2.11098f
C24 VDD1.n3 B 2.37311f
C25 VDD1.t4 B 0.237545f
C26 VDD1.t2 B 0.237545f
C27 VDD1.n4 B 2.10876f
C28 VDD1.n5 B 2.44856f
C29 VP.n0 B 0.043685f
C30 VP.n1 B 0.009913f
C31 VP.n2 B 0.043685f
C32 VP.n3 B 0.043685f
C33 VP.t5 B 1.04275f
C34 VP.t3 B 1.04275f
C35 VP.n4 B 0.043685f
C36 VP.t0 B 1.04275f
C37 VP.n5 B 0.425008f
C38 VP.t6 B 1.06599f
C39 VP.n6 B 0.401285f
C40 VP.n7 B 0.187001f
C41 VP.n8 B 0.009913f
C42 VP.n9 B 0.419411f
C43 VP.n10 B 0.009913f
C44 VP.n11 B 0.419276f
C45 VP.n12 B 1.77778f
C46 VP.n13 B 1.81538f
C47 VP.t2 B 1.04275f
C48 VP.n14 B 0.419276f
C49 VP.n15 B 0.009913f
C50 VP.t7 B 1.04275f
C51 VP.n16 B 0.419411f
C52 VP.n17 B 0.043685f
C53 VP.n18 B 0.043685f
C54 VP.n19 B 0.043685f
C55 VP.t1 B 1.04275f
C56 VP.n20 B 0.419411f
C57 VP.n21 B 0.009913f
C58 VP.t4 B 1.04275f
C59 VP.n22 B 0.419276f
C60 VP.n23 B 0.033854f
C61 VDD2.t2 B 0.23754f
C62 VDD2.t1 B 0.23754f
C63 VDD2.n0 B 2.11093f
C64 VDD2.t4 B 0.23754f
C65 VDD2.t6 B 0.23754f
C66 VDD2.n1 B 2.11093f
C67 VDD2.n2 B 2.31547f
C68 VDD2.t5 B 0.23754f
C69 VDD2.t7 B 0.23754f
C70 VDD2.n3 B 2.10872f
C71 VDD2.n4 B 2.41654f
C72 VDD2.t0 B 0.23754f
C73 VDD2.t3 B 0.23754f
C74 VDD2.n5 B 2.1109f
C75 VTAIL.t5 B 0.176519f
C76 VTAIL.t7 B 0.176519f
C77 VTAIL.n0 B 1.51087f
C78 VTAIL.n1 B 0.256421f
C79 VTAIL.t9 B 1.92675f
C80 VTAIL.n2 B 0.348555f
C81 VTAIL.t12 B 1.92675f
C82 VTAIL.n3 B 0.348555f
C83 VTAIL.t0 B 0.176519f
C84 VTAIL.t14 B 0.176519f
C85 VTAIL.n4 B 1.51087f
C86 VTAIL.n5 B 0.312817f
C87 VTAIL.t2 B 1.92675f
C88 VTAIL.n6 B 1.27123f
C89 VTAIL.t8 B 1.92676f
C90 VTAIL.n7 B 1.27121f
C91 VTAIL.t6 B 0.176519f
C92 VTAIL.t4 B 0.176519f
C93 VTAIL.n8 B 1.51087f
C94 VTAIL.n9 B 0.312812f
C95 VTAIL.t10 B 1.92676f
C96 VTAIL.n10 B 0.348543f
C97 VTAIL.t1 B 1.92676f
C98 VTAIL.n11 B 0.348543f
C99 VTAIL.t15 B 0.176519f
C100 VTAIL.t13 B 0.176519f
C101 VTAIL.n12 B 1.51087f
C102 VTAIL.n13 B 0.312812f
C103 VTAIL.t3 B 1.92675f
C104 VTAIL.n14 B 1.27123f
C105 VTAIL.t11 B 1.92675f
C106 VTAIL.n15 B 1.26747f
C107 VN.n0 B 0.042695f
C108 VN.n1 B 0.009688f
C109 VN.t5 B 1.04186f
C110 VN.t6 B 1.01914f
C111 VN.n2 B 0.415384f
C112 VN.n3 B 0.392199f
C113 VN.n4 B 0.182767f
C114 VN.n5 B 0.042695f
C115 VN.t3 B 1.01914f
C116 VN.n6 B 0.409914f
C117 VN.n7 B 0.009688f
C118 VN.t1 B 1.01914f
C119 VN.n8 B 0.409783f
C120 VN.n9 B 0.033087f
C121 VN.n10 B 0.042695f
C122 VN.n11 B 0.009688f
C123 VN.t0 B 1.01914f
C124 VN.t4 B 1.04186f
C125 VN.t7 B 1.01914f
C126 VN.n12 B 0.415384f
C127 VN.n13 B 0.392199f
C128 VN.n14 B 0.182767f
C129 VN.n15 B 0.042695f
C130 VN.n16 B 0.409914f
C131 VN.n17 B 0.009688f
C132 VN.t2 B 1.01914f
C133 VN.n18 B 0.409783f
C134 VN.n19 B 1.76557f
.ends

