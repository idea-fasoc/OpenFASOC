* NGSPICE file created from diff_pair_sample_0256.ext - technology: sky130A

.subckt diff_pair_sample_0256 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=1.09725 pd=6.98 as=1.09725 ps=6.98 w=6.65 l=2.64
X1 VTAIL.t10 VN.t1 VDD2.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.5935 pd=14.08 as=1.09725 ps=6.98 w=6.65 l=2.64
X2 VDD1.t7 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.09725 pd=6.98 as=2.5935 ps=14.08 w=6.65 l=2.64
X3 VDD1.t6 VP.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.09725 pd=6.98 as=2.5935 ps=14.08 w=6.65 l=2.64
X4 VTAIL.t6 VP.t2 VDD1.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=2.5935 pd=14.08 as=1.09725 ps=6.98 w=6.65 l=2.64
X5 VTAIL.t0 VP.t3 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.09725 pd=6.98 as=1.09725 ps=6.98 w=6.65 l=2.64
X6 VTAIL.t14 VN.t2 VDD2.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=2.5935 pd=14.08 as=1.09725 ps=6.98 w=6.65 l=2.64
X7 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=2.5935 pd=14.08 as=0 ps=0 w=6.65 l=2.64
X8 VDD2.t4 VN.t3 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=1.09725 pd=6.98 as=1.09725 ps=6.98 w=6.65 l=2.64
X9 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=2.5935 pd=14.08 as=0 ps=0 w=6.65 l=2.64
X10 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=2.5935 pd=14.08 as=0 ps=0 w=6.65 l=2.64
X11 VTAIL.t7 VP.t4 VDD1.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=1.09725 pd=6.98 as=1.09725 ps=6.98 w=6.65 l=2.64
X12 VDD1.t2 VP.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.09725 pd=6.98 as=1.09725 ps=6.98 w=6.65 l=2.64
X13 VDD2.t3 VN.t4 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=1.09725 pd=6.98 as=2.5935 ps=14.08 w=6.65 l=2.64
X14 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.5935 pd=14.08 as=0 ps=0 w=6.65 l=2.64
X15 VTAIL.t15 VN.t5 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.09725 pd=6.98 as=1.09725 ps=6.98 w=6.65 l=2.64
X16 VTAIL.t13 VN.t6 VDD2.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=1.09725 pd=6.98 as=1.09725 ps=6.98 w=6.65 l=2.64
X17 VDD2.t0 VN.t7 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=1.09725 pd=6.98 as=2.5935 ps=14.08 w=6.65 l=2.64
X18 VTAIL.t3 VP.t6 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=2.5935 pd=14.08 as=1.09725 ps=6.98 w=6.65 l=2.64
X19 VDD1.t0 VP.t7 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.09725 pd=6.98 as=1.09725 ps=6.98 w=6.65 l=2.64
R0 VN.n55 VN.n29 161.3
R1 VN.n54 VN.n53 161.3
R2 VN.n52 VN.n30 161.3
R3 VN.n51 VN.n50 161.3
R4 VN.n49 VN.n31 161.3
R5 VN.n48 VN.n47 161.3
R6 VN.n46 VN.n45 161.3
R7 VN.n44 VN.n33 161.3
R8 VN.n43 VN.n42 161.3
R9 VN.n41 VN.n34 161.3
R10 VN.n40 VN.n39 161.3
R11 VN.n38 VN.n35 161.3
R12 VN.n26 VN.n0 161.3
R13 VN.n25 VN.n24 161.3
R14 VN.n23 VN.n1 161.3
R15 VN.n22 VN.n21 161.3
R16 VN.n20 VN.n2 161.3
R17 VN.n19 VN.n18 161.3
R18 VN.n17 VN.n16 161.3
R19 VN.n15 VN.n4 161.3
R20 VN.n14 VN.n13 161.3
R21 VN.n12 VN.n5 161.3
R22 VN.n11 VN.n10 161.3
R23 VN.n9 VN.n6 161.3
R24 VN.n28 VN.n27 100.725
R25 VN.n57 VN.n56 100.725
R26 VN.n7 VN.t1 94.3223
R27 VN.n36 VN.t4 94.3223
R28 VN.n8 VN.n7 60.9555
R29 VN.n37 VN.n36 60.9555
R30 VN.n8 VN.t3 60.7069
R31 VN.n3 VN.t5 60.7069
R32 VN.n27 VN.t7 60.7069
R33 VN.n37 VN.t6 60.7069
R34 VN.n32 VN.t0 60.7069
R35 VN.n56 VN.t2 60.7069
R36 VN.n14 VN.n5 56.5193
R37 VN.n21 VN.n1 56.5193
R38 VN.n43 VN.n34 56.5193
R39 VN.n50 VN.n30 56.5193
R40 VN VN.n57 47.3391
R41 VN.n10 VN.n9 24.4675
R42 VN.n10 VN.n5 24.4675
R43 VN.n15 VN.n14 24.4675
R44 VN.n16 VN.n15 24.4675
R45 VN.n20 VN.n19 24.4675
R46 VN.n21 VN.n20 24.4675
R47 VN.n25 VN.n1 24.4675
R48 VN.n26 VN.n25 24.4675
R49 VN.n39 VN.n34 24.4675
R50 VN.n39 VN.n38 24.4675
R51 VN.n50 VN.n49 24.4675
R52 VN.n49 VN.n48 24.4675
R53 VN.n45 VN.n44 24.4675
R54 VN.n44 VN.n43 24.4675
R55 VN.n55 VN.n54 24.4675
R56 VN.n54 VN.n30 24.4675
R57 VN.n19 VN.n3 12.968
R58 VN.n48 VN.n32 12.968
R59 VN.n9 VN.n8 11.5
R60 VN.n16 VN.n3 11.5
R61 VN.n38 VN.n37 11.5
R62 VN.n45 VN.n32 11.5
R63 VN.n27 VN.n26 10.032
R64 VN.n56 VN.n55 10.032
R65 VN.n36 VN.n35 6.848
R66 VN.n7 VN.n6 6.848
R67 VN.n57 VN.n29 0.278367
R68 VN.n28 VN.n0 0.278367
R69 VN.n53 VN.n29 0.189894
R70 VN.n53 VN.n52 0.189894
R71 VN.n52 VN.n51 0.189894
R72 VN.n51 VN.n31 0.189894
R73 VN.n47 VN.n31 0.189894
R74 VN.n47 VN.n46 0.189894
R75 VN.n46 VN.n33 0.189894
R76 VN.n42 VN.n33 0.189894
R77 VN.n42 VN.n41 0.189894
R78 VN.n41 VN.n40 0.189894
R79 VN.n40 VN.n35 0.189894
R80 VN.n11 VN.n6 0.189894
R81 VN.n12 VN.n11 0.189894
R82 VN.n13 VN.n12 0.189894
R83 VN.n13 VN.n4 0.189894
R84 VN.n17 VN.n4 0.189894
R85 VN.n18 VN.n17 0.189894
R86 VN.n18 VN.n2 0.189894
R87 VN.n22 VN.n2 0.189894
R88 VN.n23 VN.n22 0.189894
R89 VN.n24 VN.n23 0.189894
R90 VN.n24 VN.n0 0.189894
R91 VN VN.n28 0.153454
R92 VTAIL.n290 VTAIL.n260 289.615
R93 VTAIL.n32 VTAIL.n2 289.615
R94 VTAIL.n68 VTAIL.n38 289.615
R95 VTAIL.n106 VTAIL.n76 289.615
R96 VTAIL.n254 VTAIL.n224 289.615
R97 VTAIL.n216 VTAIL.n186 289.615
R98 VTAIL.n180 VTAIL.n150 289.615
R99 VTAIL.n142 VTAIL.n112 289.615
R100 VTAIL.n273 VTAIL.n272 185
R101 VTAIL.n275 VTAIL.n274 185
R102 VTAIL.n268 VTAIL.n267 185
R103 VTAIL.n281 VTAIL.n280 185
R104 VTAIL.n283 VTAIL.n282 185
R105 VTAIL.n264 VTAIL.n263 185
R106 VTAIL.n289 VTAIL.n288 185
R107 VTAIL.n291 VTAIL.n290 185
R108 VTAIL.n15 VTAIL.n14 185
R109 VTAIL.n17 VTAIL.n16 185
R110 VTAIL.n10 VTAIL.n9 185
R111 VTAIL.n23 VTAIL.n22 185
R112 VTAIL.n25 VTAIL.n24 185
R113 VTAIL.n6 VTAIL.n5 185
R114 VTAIL.n31 VTAIL.n30 185
R115 VTAIL.n33 VTAIL.n32 185
R116 VTAIL.n51 VTAIL.n50 185
R117 VTAIL.n53 VTAIL.n52 185
R118 VTAIL.n46 VTAIL.n45 185
R119 VTAIL.n59 VTAIL.n58 185
R120 VTAIL.n61 VTAIL.n60 185
R121 VTAIL.n42 VTAIL.n41 185
R122 VTAIL.n67 VTAIL.n66 185
R123 VTAIL.n69 VTAIL.n68 185
R124 VTAIL.n89 VTAIL.n88 185
R125 VTAIL.n91 VTAIL.n90 185
R126 VTAIL.n84 VTAIL.n83 185
R127 VTAIL.n97 VTAIL.n96 185
R128 VTAIL.n99 VTAIL.n98 185
R129 VTAIL.n80 VTAIL.n79 185
R130 VTAIL.n105 VTAIL.n104 185
R131 VTAIL.n107 VTAIL.n106 185
R132 VTAIL.n255 VTAIL.n254 185
R133 VTAIL.n253 VTAIL.n252 185
R134 VTAIL.n228 VTAIL.n227 185
R135 VTAIL.n247 VTAIL.n246 185
R136 VTAIL.n245 VTAIL.n244 185
R137 VTAIL.n232 VTAIL.n231 185
R138 VTAIL.n239 VTAIL.n238 185
R139 VTAIL.n237 VTAIL.n236 185
R140 VTAIL.n217 VTAIL.n216 185
R141 VTAIL.n215 VTAIL.n214 185
R142 VTAIL.n190 VTAIL.n189 185
R143 VTAIL.n209 VTAIL.n208 185
R144 VTAIL.n207 VTAIL.n206 185
R145 VTAIL.n194 VTAIL.n193 185
R146 VTAIL.n201 VTAIL.n200 185
R147 VTAIL.n199 VTAIL.n198 185
R148 VTAIL.n181 VTAIL.n180 185
R149 VTAIL.n179 VTAIL.n178 185
R150 VTAIL.n154 VTAIL.n153 185
R151 VTAIL.n173 VTAIL.n172 185
R152 VTAIL.n171 VTAIL.n170 185
R153 VTAIL.n158 VTAIL.n157 185
R154 VTAIL.n165 VTAIL.n164 185
R155 VTAIL.n163 VTAIL.n162 185
R156 VTAIL.n143 VTAIL.n142 185
R157 VTAIL.n141 VTAIL.n140 185
R158 VTAIL.n116 VTAIL.n115 185
R159 VTAIL.n135 VTAIL.n134 185
R160 VTAIL.n133 VTAIL.n132 185
R161 VTAIL.n120 VTAIL.n119 185
R162 VTAIL.n127 VTAIL.n126 185
R163 VTAIL.n125 VTAIL.n124 185
R164 VTAIL.n271 VTAIL.t8 147.659
R165 VTAIL.n13 VTAIL.t10 147.659
R166 VTAIL.n49 VTAIL.t4 147.659
R167 VTAIL.n87 VTAIL.t6 147.659
R168 VTAIL.n235 VTAIL.t2 147.659
R169 VTAIL.n197 VTAIL.t3 147.659
R170 VTAIL.n161 VTAIL.t9 147.659
R171 VTAIL.n123 VTAIL.t14 147.659
R172 VTAIL.n274 VTAIL.n273 104.615
R173 VTAIL.n274 VTAIL.n267 104.615
R174 VTAIL.n281 VTAIL.n267 104.615
R175 VTAIL.n282 VTAIL.n281 104.615
R176 VTAIL.n282 VTAIL.n263 104.615
R177 VTAIL.n289 VTAIL.n263 104.615
R178 VTAIL.n290 VTAIL.n289 104.615
R179 VTAIL.n16 VTAIL.n15 104.615
R180 VTAIL.n16 VTAIL.n9 104.615
R181 VTAIL.n23 VTAIL.n9 104.615
R182 VTAIL.n24 VTAIL.n23 104.615
R183 VTAIL.n24 VTAIL.n5 104.615
R184 VTAIL.n31 VTAIL.n5 104.615
R185 VTAIL.n32 VTAIL.n31 104.615
R186 VTAIL.n52 VTAIL.n51 104.615
R187 VTAIL.n52 VTAIL.n45 104.615
R188 VTAIL.n59 VTAIL.n45 104.615
R189 VTAIL.n60 VTAIL.n59 104.615
R190 VTAIL.n60 VTAIL.n41 104.615
R191 VTAIL.n67 VTAIL.n41 104.615
R192 VTAIL.n68 VTAIL.n67 104.615
R193 VTAIL.n90 VTAIL.n89 104.615
R194 VTAIL.n90 VTAIL.n83 104.615
R195 VTAIL.n97 VTAIL.n83 104.615
R196 VTAIL.n98 VTAIL.n97 104.615
R197 VTAIL.n98 VTAIL.n79 104.615
R198 VTAIL.n105 VTAIL.n79 104.615
R199 VTAIL.n106 VTAIL.n105 104.615
R200 VTAIL.n254 VTAIL.n253 104.615
R201 VTAIL.n253 VTAIL.n227 104.615
R202 VTAIL.n246 VTAIL.n227 104.615
R203 VTAIL.n246 VTAIL.n245 104.615
R204 VTAIL.n245 VTAIL.n231 104.615
R205 VTAIL.n238 VTAIL.n231 104.615
R206 VTAIL.n238 VTAIL.n237 104.615
R207 VTAIL.n216 VTAIL.n215 104.615
R208 VTAIL.n215 VTAIL.n189 104.615
R209 VTAIL.n208 VTAIL.n189 104.615
R210 VTAIL.n208 VTAIL.n207 104.615
R211 VTAIL.n207 VTAIL.n193 104.615
R212 VTAIL.n200 VTAIL.n193 104.615
R213 VTAIL.n200 VTAIL.n199 104.615
R214 VTAIL.n180 VTAIL.n179 104.615
R215 VTAIL.n179 VTAIL.n153 104.615
R216 VTAIL.n172 VTAIL.n153 104.615
R217 VTAIL.n172 VTAIL.n171 104.615
R218 VTAIL.n171 VTAIL.n157 104.615
R219 VTAIL.n164 VTAIL.n157 104.615
R220 VTAIL.n164 VTAIL.n163 104.615
R221 VTAIL.n142 VTAIL.n141 104.615
R222 VTAIL.n141 VTAIL.n115 104.615
R223 VTAIL.n134 VTAIL.n115 104.615
R224 VTAIL.n134 VTAIL.n133 104.615
R225 VTAIL.n133 VTAIL.n119 104.615
R226 VTAIL.n126 VTAIL.n119 104.615
R227 VTAIL.n126 VTAIL.n125 104.615
R228 VTAIL.n273 VTAIL.t8 52.3082
R229 VTAIL.n15 VTAIL.t10 52.3082
R230 VTAIL.n51 VTAIL.t4 52.3082
R231 VTAIL.n89 VTAIL.t6 52.3082
R232 VTAIL.n237 VTAIL.t2 52.3082
R233 VTAIL.n199 VTAIL.t3 52.3082
R234 VTAIL.n163 VTAIL.t9 52.3082
R235 VTAIL.n125 VTAIL.t14 52.3082
R236 VTAIL.n223 VTAIL.n222 48.0378
R237 VTAIL.n149 VTAIL.n148 48.0378
R238 VTAIL.n1 VTAIL.n0 48.0376
R239 VTAIL.n75 VTAIL.n74 48.0376
R240 VTAIL.n295 VTAIL.n294 30.8278
R241 VTAIL.n37 VTAIL.n36 30.8278
R242 VTAIL.n73 VTAIL.n72 30.8278
R243 VTAIL.n111 VTAIL.n110 30.8278
R244 VTAIL.n259 VTAIL.n258 30.8278
R245 VTAIL.n221 VTAIL.n220 30.8278
R246 VTAIL.n185 VTAIL.n184 30.8278
R247 VTAIL.n147 VTAIL.n146 30.8278
R248 VTAIL.n295 VTAIL.n259 20.66
R249 VTAIL.n147 VTAIL.n111 20.66
R250 VTAIL.n272 VTAIL.n271 15.6676
R251 VTAIL.n14 VTAIL.n13 15.6676
R252 VTAIL.n50 VTAIL.n49 15.6676
R253 VTAIL.n88 VTAIL.n87 15.6676
R254 VTAIL.n236 VTAIL.n235 15.6676
R255 VTAIL.n198 VTAIL.n197 15.6676
R256 VTAIL.n162 VTAIL.n161 15.6676
R257 VTAIL.n124 VTAIL.n123 15.6676
R258 VTAIL.n275 VTAIL.n270 12.8005
R259 VTAIL.n17 VTAIL.n12 12.8005
R260 VTAIL.n53 VTAIL.n48 12.8005
R261 VTAIL.n91 VTAIL.n86 12.8005
R262 VTAIL.n239 VTAIL.n234 12.8005
R263 VTAIL.n201 VTAIL.n196 12.8005
R264 VTAIL.n165 VTAIL.n160 12.8005
R265 VTAIL.n127 VTAIL.n122 12.8005
R266 VTAIL.n276 VTAIL.n268 12.0247
R267 VTAIL.n18 VTAIL.n10 12.0247
R268 VTAIL.n54 VTAIL.n46 12.0247
R269 VTAIL.n92 VTAIL.n84 12.0247
R270 VTAIL.n240 VTAIL.n232 12.0247
R271 VTAIL.n202 VTAIL.n194 12.0247
R272 VTAIL.n166 VTAIL.n158 12.0247
R273 VTAIL.n128 VTAIL.n120 12.0247
R274 VTAIL.n280 VTAIL.n279 11.249
R275 VTAIL.n22 VTAIL.n21 11.249
R276 VTAIL.n58 VTAIL.n57 11.249
R277 VTAIL.n96 VTAIL.n95 11.249
R278 VTAIL.n244 VTAIL.n243 11.249
R279 VTAIL.n206 VTAIL.n205 11.249
R280 VTAIL.n170 VTAIL.n169 11.249
R281 VTAIL.n132 VTAIL.n131 11.249
R282 VTAIL.n283 VTAIL.n266 10.4732
R283 VTAIL.n25 VTAIL.n8 10.4732
R284 VTAIL.n61 VTAIL.n44 10.4732
R285 VTAIL.n99 VTAIL.n82 10.4732
R286 VTAIL.n247 VTAIL.n230 10.4732
R287 VTAIL.n209 VTAIL.n192 10.4732
R288 VTAIL.n173 VTAIL.n156 10.4732
R289 VTAIL.n135 VTAIL.n118 10.4732
R290 VTAIL.n284 VTAIL.n264 9.69747
R291 VTAIL.n26 VTAIL.n6 9.69747
R292 VTAIL.n62 VTAIL.n42 9.69747
R293 VTAIL.n100 VTAIL.n80 9.69747
R294 VTAIL.n248 VTAIL.n228 9.69747
R295 VTAIL.n210 VTAIL.n190 9.69747
R296 VTAIL.n174 VTAIL.n154 9.69747
R297 VTAIL.n136 VTAIL.n116 9.69747
R298 VTAIL.n294 VTAIL.n293 9.45567
R299 VTAIL.n36 VTAIL.n35 9.45567
R300 VTAIL.n72 VTAIL.n71 9.45567
R301 VTAIL.n110 VTAIL.n109 9.45567
R302 VTAIL.n258 VTAIL.n257 9.45567
R303 VTAIL.n220 VTAIL.n219 9.45567
R304 VTAIL.n184 VTAIL.n183 9.45567
R305 VTAIL.n146 VTAIL.n145 9.45567
R306 VTAIL.n262 VTAIL.n261 9.3005
R307 VTAIL.n287 VTAIL.n286 9.3005
R308 VTAIL.n285 VTAIL.n284 9.3005
R309 VTAIL.n266 VTAIL.n265 9.3005
R310 VTAIL.n279 VTAIL.n278 9.3005
R311 VTAIL.n277 VTAIL.n276 9.3005
R312 VTAIL.n270 VTAIL.n269 9.3005
R313 VTAIL.n293 VTAIL.n292 9.3005
R314 VTAIL.n4 VTAIL.n3 9.3005
R315 VTAIL.n29 VTAIL.n28 9.3005
R316 VTAIL.n27 VTAIL.n26 9.3005
R317 VTAIL.n8 VTAIL.n7 9.3005
R318 VTAIL.n21 VTAIL.n20 9.3005
R319 VTAIL.n19 VTAIL.n18 9.3005
R320 VTAIL.n12 VTAIL.n11 9.3005
R321 VTAIL.n35 VTAIL.n34 9.3005
R322 VTAIL.n40 VTAIL.n39 9.3005
R323 VTAIL.n65 VTAIL.n64 9.3005
R324 VTAIL.n63 VTAIL.n62 9.3005
R325 VTAIL.n44 VTAIL.n43 9.3005
R326 VTAIL.n57 VTAIL.n56 9.3005
R327 VTAIL.n55 VTAIL.n54 9.3005
R328 VTAIL.n48 VTAIL.n47 9.3005
R329 VTAIL.n71 VTAIL.n70 9.3005
R330 VTAIL.n78 VTAIL.n77 9.3005
R331 VTAIL.n103 VTAIL.n102 9.3005
R332 VTAIL.n101 VTAIL.n100 9.3005
R333 VTAIL.n82 VTAIL.n81 9.3005
R334 VTAIL.n95 VTAIL.n94 9.3005
R335 VTAIL.n93 VTAIL.n92 9.3005
R336 VTAIL.n86 VTAIL.n85 9.3005
R337 VTAIL.n109 VTAIL.n108 9.3005
R338 VTAIL.n257 VTAIL.n256 9.3005
R339 VTAIL.n226 VTAIL.n225 9.3005
R340 VTAIL.n251 VTAIL.n250 9.3005
R341 VTAIL.n249 VTAIL.n248 9.3005
R342 VTAIL.n230 VTAIL.n229 9.3005
R343 VTAIL.n243 VTAIL.n242 9.3005
R344 VTAIL.n241 VTAIL.n240 9.3005
R345 VTAIL.n234 VTAIL.n233 9.3005
R346 VTAIL.n219 VTAIL.n218 9.3005
R347 VTAIL.n188 VTAIL.n187 9.3005
R348 VTAIL.n213 VTAIL.n212 9.3005
R349 VTAIL.n211 VTAIL.n210 9.3005
R350 VTAIL.n192 VTAIL.n191 9.3005
R351 VTAIL.n205 VTAIL.n204 9.3005
R352 VTAIL.n203 VTAIL.n202 9.3005
R353 VTAIL.n196 VTAIL.n195 9.3005
R354 VTAIL.n183 VTAIL.n182 9.3005
R355 VTAIL.n152 VTAIL.n151 9.3005
R356 VTAIL.n177 VTAIL.n176 9.3005
R357 VTAIL.n175 VTAIL.n174 9.3005
R358 VTAIL.n156 VTAIL.n155 9.3005
R359 VTAIL.n169 VTAIL.n168 9.3005
R360 VTAIL.n167 VTAIL.n166 9.3005
R361 VTAIL.n160 VTAIL.n159 9.3005
R362 VTAIL.n145 VTAIL.n144 9.3005
R363 VTAIL.n114 VTAIL.n113 9.3005
R364 VTAIL.n139 VTAIL.n138 9.3005
R365 VTAIL.n137 VTAIL.n136 9.3005
R366 VTAIL.n118 VTAIL.n117 9.3005
R367 VTAIL.n131 VTAIL.n130 9.3005
R368 VTAIL.n129 VTAIL.n128 9.3005
R369 VTAIL.n122 VTAIL.n121 9.3005
R370 VTAIL.n288 VTAIL.n287 8.92171
R371 VTAIL.n30 VTAIL.n29 8.92171
R372 VTAIL.n66 VTAIL.n65 8.92171
R373 VTAIL.n104 VTAIL.n103 8.92171
R374 VTAIL.n252 VTAIL.n251 8.92171
R375 VTAIL.n214 VTAIL.n213 8.92171
R376 VTAIL.n178 VTAIL.n177 8.92171
R377 VTAIL.n140 VTAIL.n139 8.92171
R378 VTAIL.n291 VTAIL.n262 8.14595
R379 VTAIL.n33 VTAIL.n4 8.14595
R380 VTAIL.n69 VTAIL.n40 8.14595
R381 VTAIL.n107 VTAIL.n78 8.14595
R382 VTAIL.n255 VTAIL.n226 8.14595
R383 VTAIL.n217 VTAIL.n188 8.14595
R384 VTAIL.n181 VTAIL.n152 8.14595
R385 VTAIL.n143 VTAIL.n114 8.14595
R386 VTAIL.n292 VTAIL.n260 7.3702
R387 VTAIL.n34 VTAIL.n2 7.3702
R388 VTAIL.n70 VTAIL.n38 7.3702
R389 VTAIL.n108 VTAIL.n76 7.3702
R390 VTAIL.n256 VTAIL.n224 7.3702
R391 VTAIL.n218 VTAIL.n186 7.3702
R392 VTAIL.n182 VTAIL.n150 7.3702
R393 VTAIL.n144 VTAIL.n112 7.3702
R394 VTAIL.n294 VTAIL.n260 6.59444
R395 VTAIL.n36 VTAIL.n2 6.59444
R396 VTAIL.n72 VTAIL.n38 6.59444
R397 VTAIL.n110 VTAIL.n76 6.59444
R398 VTAIL.n258 VTAIL.n224 6.59444
R399 VTAIL.n220 VTAIL.n186 6.59444
R400 VTAIL.n184 VTAIL.n150 6.59444
R401 VTAIL.n146 VTAIL.n112 6.59444
R402 VTAIL.n292 VTAIL.n291 5.81868
R403 VTAIL.n34 VTAIL.n33 5.81868
R404 VTAIL.n70 VTAIL.n69 5.81868
R405 VTAIL.n108 VTAIL.n107 5.81868
R406 VTAIL.n256 VTAIL.n255 5.81868
R407 VTAIL.n218 VTAIL.n217 5.81868
R408 VTAIL.n182 VTAIL.n181 5.81868
R409 VTAIL.n144 VTAIL.n143 5.81868
R410 VTAIL.n288 VTAIL.n262 5.04292
R411 VTAIL.n30 VTAIL.n4 5.04292
R412 VTAIL.n66 VTAIL.n40 5.04292
R413 VTAIL.n104 VTAIL.n78 5.04292
R414 VTAIL.n252 VTAIL.n226 5.04292
R415 VTAIL.n214 VTAIL.n188 5.04292
R416 VTAIL.n178 VTAIL.n152 5.04292
R417 VTAIL.n140 VTAIL.n114 5.04292
R418 VTAIL.n271 VTAIL.n269 4.38571
R419 VTAIL.n13 VTAIL.n11 4.38571
R420 VTAIL.n49 VTAIL.n47 4.38571
R421 VTAIL.n87 VTAIL.n85 4.38571
R422 VTAIL.n235 VTAIL.n233 4.38571
R423 VTAIL.n197 VTAIL.n195 4.38571
R424 VTAIL.n161 VTAIL.n159 4.38571
R425 VTAIL.n123 VTAIL.n121 4.38571
R426 VTAIL.n287 VTAIL.n264 4.26717
R427 VTAIL.n29 VTAIL.n6 4.26717
R428 VTAIL.n65 VTAIL.n42 4.26717
R429 VTAIL.n103 VTAIL.n80 4.26717
R430 VTAIL.n251 VTAIL.n228 4.26717
R431 VTAIL.n213 VTAIL.n190 4.26717
R432 VTAIL.n177 VTAIL.n154 4.26717
R433 VTAIL.n139 VTAIL.n116 4.26717
R434 VTAIL.n284 VTAIL.n283 3.49141
R435 VTAIL.n26 VTAIL.n25 3.49141
R436 VTAIL.n62 VTAIL.n61 3.49141
R437 VTAIL.n100 VTAIL.n99 3.49141
R438 VTAIL.n248 VTAIL.n247 3.49141
R439 VTAIL.n210 VTAIL.n209 3.49141
R440 VTAIL.n174 VTAIL.n173 3.49141
R441 VTAIL.n136 VTAIL.n135 3.49141
R442 VTAIL.n0 VTAIL.t12 2.97794
R443 VTAIL.n0 VTAIL.t15 2.97794
R444 VTAIL.n74 VTAIL.t1 2.97794
R445 VTAIL.n74 VTAIL.t7 2.97794
R446 VTAIL.n222 VTAIL.t5 2.97794
R447 VTAIL.n222 VTAIL.t0 2.97794
R448 VTAIL.n148 VTAIL.t11 2.97794
R449 VTAIL.n148 VTAIL.t13 2.97794
R450 VTAIL.n280 VTAIL.n266 2.71565
R451 VTAIL.n22 VTAIL.n8 2.71565
R452 VTAIL.n58 VTAIL.n44 2.71565
R453 VTAIL.n96 VTAIL.n82 2.71565
R454 VTAIL.n244 VTAIL.n230 2.71565
R455 VTAIL.n206 VTAIL.n192 2.71565
R456 VTAIL.n170 VTAIL.n156 2.71565
R457 VTAIL.n132 VTAIL.n118 2.71565
R458 VTAIL.n149 VTAIL.n147 2.56084
R459 VTAIL.n185 VTAIL.n149 2.56084
R460 VTAIL.n223 VTAIL.n221 2.56084
R461 VTAIL.n259 VTAIL.n223 2.56084
R462 VTAIL.n111 VTAIL.n75 2.56084
R463 VTAIL.n75 VTAIL.n73 2.56084
R464 VTAIL.n37 VTAIL.n1 2.56084
R465 VTAIL VTAIL.n295 2.50266
R466 VTAIL.n279 VTAIL.n268 1.93989
R467 VTAIL.n21 VTAIL.n10 1.93989
R468 VTAIL.n57 VTAIL.n46 1.93989
R469 VTAIL.n95 VTAIL.n84 1.93989
R470 VTAIL.n243 VTAIL.n232 1.93989
R471 VTAIL.n205 VTAIL.n194 1.93989
R472 VTAIL.n169 VTAIL.n158 1.93989
R473 VTAIL.n131 VTAIL.n120 1.93989
R474 VTAIL.n276 VTAIL.n275 1.16414
R475 VTAIL.n18 VTAIL.n17 1.16414
R476 VTAIL.n54 VTAIL.n53 1.16414
R477 VTAIL.n92 VTAIL.n91 1.16414
R478 VTAIL.n240 VTAIL.n239 1.16414
R479 VTAIL.n202 VTAIL.n201 1.16414
R480 VTAIL.n166 VTAIL.n165 1.16414
R481 VTAIL.n128 VTAIL.n127 1.16414
R482 VTAIL.n221 VTAIL.n185 0.470328
R483 VTAIL.n73 VTAIL.n37 0.470328
R484 VTAIL.n272 VTAIL.n270 0.388379
R485 VTAIL.n14 VTAIL.n12 0.388379
R486 VTAIL.n50 VTAIL.n48 0.388379
R487 VTAIL.n88 VTAIL.n86 0.388379
R488 VTAIL.n236 VTAIL.n234 0.388379
R489 VTAIL.n198 VTAIL.n196 0.388379
R490 VTAIL.n162 VTAIL.n160 0.388379
R491 VTAIL.n124 VTAIL.n122 0.388379
R492 VTAIL.n277 VTAIL.n269 0.155672
R493 VTAIL.n278 VTAIL.n277 0.155672
R494 VTAIL.n278 VTAIL.n265 0.155672
R495 VTAIL.n285 VTAIL.n265 0.155672
R496 VTAIL.n286 VTAIL.n285 0.155672
R497 VTAIL.n286 VTAIL.n261 0.155672
R498 VTAIL.n293 VTAIL.n261 0.155672
R499 VTAIL.n19 VTAIL.n11 0.155672
R500 VTAIL.n20 VTAIL.n19 0.155672
R501 VTAIL.n20 VTAIL.n7 0.155672
R502 VTAIL.n27 VTAIL.n7 0.155672
R503 VTAIL.n28 VTAIL.n27 0.155672
R504 VTAIL.n28 VTAIL.n3 0.155672
R505 VTAIL.n35 VTAIL.n3 0.155672
R506 VTAIL.n55 VTAIL.n47 0.155672
R507 VTAIL.n56 VTAIL.n55 0.155672
R508 VTAIL.n56 VTAIL.n43 0.155672
R509 VTAIL.n63 VTAIL.n43 0.155672
R510 VTAIL.n64 VTAIL.n63 0.155672
R511 VTAIL.n64 VTAIL.n39 0.155672
R512 VTAIL.n71 VTAIL.n39 0.155672
R513 VTAIL.n93 VTAIL.n85 0.155672
R514 VTAIL.n94 VTAIL.n93 0.155672
R515 VTAIL.n94 VTAIL.n81 0.155672
R516 VTAIL.n101 VTAIL.n81 0.155672
R517 VTAIL.n102 VTAIL.n101 0.155672
R518 VTAIL.n102 VTAIL.n77 0.155672
R519 VTAIL.n109 VTAIL.n77 0.155672
R520 VTAIL.n257 VTAIL.n225 0.155672
R521 VTAIL.n250 VTAIL.n225 0.155672
R522 VTAIL.n250 VTAIL.n249 0.155672
R523 VTAIL.n249 VTAIL.n229 0.155672
R524 VTAIL.n242 VTAIL.n229 0.155672
R525 VTAIL.n242 VTAIL.n241 0.155672
R526 VTAIL.n241 VTAIL.n233 0.155672
R527 VTAIL.n219 VTAIL.n187 0.155672
R528 VTAIL.n212 VTAIL.n187 0.155672
R529 VTAIL.n212 VTAIL.n211 0.155672
R530 VTAIL.n211 VTAIL.n191 0.155672
R531 VTAIL.n204 VTAIL.n191 0.155672
R532 VTAIL.n204 VTAIL.n203 0.155672
R533 VTAIL.n203 VTAIL.n195 0.155672
R534 VTAIL.n183 VTAIL.n151 0.155672
R535 VTAIL.n176 VTAIL.n151 0.155672
R536 VTAIL.n176 VTAIL.n175 0.155672
R537 VTAIL.n175 VTAIL.n155 0.155672
R538 VTAIL.n168 VTAIL.n155 0.155672
R539 VTAIL.n168 VTAIL.n167 0.155672
R540 VTAIL.n167 VTAIL.n159 0.155672
R541 VTAIL.n145 VTAIL.n113 0.155672
R542 VTAIL.n138 VTAIL.n113 0.155672
R543 VTAIL.n138 VTAIL.n137 0.155672
R544 VTAIL.n137 VTAIL.n117 0.155672
R545 VTAIL.n130 VTAIL.n117 0.155672
R546 VTAIL.n130 VTAIL.n129 0.155672
R547 VTAIL.n129 VTAIL.n121 0.155672
R548 VTAIL VTAIL.n1 0.0586897
R549 VDD2.n2 VDD2.n1 65.9412
R550 VDD2.n2 VDD2.n0 65.9412
R551 VDD2 VDD2.n5 65.9384
R552 VDD2.n4 VDD2.n3 64.7165
R553 VDD2.n4 VDD2.n2 40.9696
R554 VDD2.n5 VDD2.t1 2.97794
R555 VDD2.n5 VDD2.t3 2.97794
R556 VDD2.n3 VDD2.t5 2.97794
R557 VDD2.n3 VDD2.t7 2.97794
R558 VDD2.n1 VDD2.t2 2.97794
R559 VDD2.n1 VDD2.t0 2.97794
R560 VDD2.n0 VDD2.t6 2.97794
R561 VDD2.n0 VDD2.t4 2.97794
R562 VDD2 VDD2.n4 1.33886
R563 B.n727 B.n726 585
R564 B.n728 B.n727 585
R565 B.n248 B.n126 585
R566 B.n247 B.n246 585
R567 B.n245 B.n244 585
R568 B.n243 B.n242 585
R569 B.n241 B.n240 585
R570 B.n239 B.n238 585
R571 B.n237 B.n236 585
R572 B.n235 B.n234 585
R573 B.n233 B.n232 585
R574 B.n231 B.n230 585
R575 B.n229 B.n228 585
R576 B.n227 B.n226 585
R577 B.n225 B.n224 585
R578 B.n223 B.n222 585
R579 B.n221 B.n220 585
R580 B.n219 B.n218 585
R581 B.n217 B.n216 585
R582 B.n215 B.n214 585
R583 B.n213 B.n212 585
R584 B.n211 B.n210 585
R585 B.n209 B.n208 585
R586 B.n207 B.n206 585
R587 B.n205 B.n204 585
R588 B.n203 B.n202 585
R589 B.n201 B.n200 585
R590 B.n198 B.n197 585
R591 B.n196 B.n195 585
R592 B.n194 B.n193 585
R593 B.n192 B.n191 585
R594 B.n190 B.n189 585
R595 B.n188 B.n187 585
R596 B.n186 B.n185 585
R597 B.n184 B.n183 585
R598 B.n182 B.n181 585
R599 B.n180 B.n179 585
R600 B.n178 B.n177 585
R601 B.n176 B.n175 585
R602 B.n174 B.n173 585
R603 B.n172 B.n171 585
R604 B.n170 B.n169 585
R605 B.n168 B.n167 585
R606 B.n166 B.n165 585
R607 B.n164 B.n163 585
R608 B.n162 B.n161 585
R609 B.n160 B.n159 585
R610 B.n158 B.n157 585
R611 B.n156 B.n155 585
R612 B.n154 B.n153 585
R613 B.n152 B.n151 585
R614 B.n150 B.n149 585
R615 B.n148 B.n147 585
R616 B.n146 B.n145 585
R617 B.n144 B.n143 585
R618 B.n142 B.n141 585
R619 B.n140 B.n139 585
R620 B.n138 B.n137 585
R621 B.n136 B.n135 585
R622 B.n134 B.n133 585
R623 B.n96 B.n95 585
R624 B.n731 B.n730 585
R625 B.n725 B.n127 585
R626 B.n127 B.n93 585
R627 B.n724 B.n92 585
R628 B.n735 B.n92 585
R629 B.n723 B.n91 585
R630 B.n736 B.n91 585
R631 B.n722 B.n90 585
R632 B.n737 B.n90 585
R633 B.n721 B.n720 585
R634 B.n720 B.n86 585
R635 B.n719 B.n85 585
R636 B.n743 B.n85 585
R637 B.n718 B.n84 585
R638 B.n744 B.n84 585
R639 B.n717 B.n83 585
R640 B.n745 B.n83 585
R641 B.n716 B.n715 585
R642 B.n715 B.n79 585
R643 B.n714 B.n78 585
R644 B.n751 B.n78 585
R645 B.n713 B.n77 585
R646 B.n752 B.n77 585
R647 B.n712 B.n76 585
R648 B.n753 B.n76 585
R649 B.n711 B.n710 585
R650 B.n710 B.n72 585
R651 B.n709 B.n71 585
R652 B.n759 B.n71 585
R653 B.n708 B.n70 585
R654 B.n760 B.n70 585
R655 B.n707 B.n69 585
R656 B.n761 B.n69 585
R657 B.n706 B.n705 585
R658 B.n705 B.n65 585
R659 B.n704 B.n64 585
R660 B.n767 B.n64 585
R661 B.n703 B.n63 585
R662 B.n768 B.n63 585
R663 B.n702 B.n62 585
R664 B.n769 B.n62 585
R665 B.n701 B.n700 585
R666 B.n700 B.n58 585
R667 B.n699 B.n57 585
R668 B.n775 B.n57 585
R669 B.n698 B.n56 585
R670 B.n776 B.n56 585
R671 B.n697 B.n55 585
R672 B.n777 B.n55 585
R673 B.n696 B.n695 585
R674 B.n695 B.n51 585
R675 B.n694 B.n50 585
R676 B.n783 B.n50 585
R677 B.n693 B.n49 585
R678 B.n784 B.n49 585
R679 B.n692 B.n48 585
R680 B.n785 B.n48 585
R681 B.n691 B.n690 585
R682 B.n690 B.n47 585
R683 B.n689 B.n43 585
R684 B.n791 B.n43 585
R685 B.n688 B.n42 585
R686 B.n792 B.n42 585
R687 B.n687 B.n41 585
R688 B.n793 B.n41 585
R689 B.n686 B.n685 585
R690 B.n685 B.n37 585
R691 B.n684 B.n36 585
R692 B.n799 B.n36 585
R693 B.n683 B.n35 585
R694 B.n800 B.n35 585
R695 B.n682 B.n34 585
R696 B.n801 B.n34 585
R697 B.n681 B.n680 585
R698 B.n680 B.n33 585
R699 B.n679 B.n29 585
R700 B.n807 B.n29 585
R701 B.n678 B.n28 585
R702 B.n808 B.n28 585
R703 B.n677 B.n27 585
R704 B.n809 B.n27 585
R705 B.n676 B.n675 585
R706 B.n675 B.n23 585
R707 B.n674 B.n22 585
R708 B.n815 B.n22 585
R709 B.n673 B.n21 585
R710 B.n816 B.n21 585
R711 B.n672 B.n20 585
R712 B.n817 B.n20 585
R713 B.n671 B.n670 585
R714 B.n670 B.n16 585
R715 B.n669 B.n15 585
R716 B.n823 B.n15 585
R717 B.n668 B.n14 585
R718 B.n824 B.n14 585
R719 B.n667 B.n13 585
R720 B.n825 B.n13 585
R721 B.n666 B.n665 585
R722 B.n665 B.n12 585
R723 B.n664 B.n663 585
R724 B.n664 B.n8 585
R725 B.n662 B.n7 585
R726 B.n832 B.n7 585
R727 B.n661 B.n6 585
R728 B.n833 B.n6 585
R729 B.n660 B.n5 585
R730 B.n834 B.n5 585
R731 B.n659 B.n658 585
R732 B.n658 B.n4 585
R733 B.n657 B.n249 585
R734 B.n657 B.n656 585
R735 B.n647 B.n250 585
R736 B.n251 B.n250 585
R737 B.n649 B.n648 585
R738 B.n650 B.n649 585
R739 B.n646 B.n256 585
R740 B.n256 B.n255 585
R741 B.n645 B.n644 585
R742 B.n644 B.n643 585
R743 B.n258 B.n257 585
R744 B.n259 B.n258 585
R745 B.n636 B.n635 585
R746 B.n637 B.n636 585
R747 B.n634 B.n264 585
R748 B.n264 B.n263 585
R749 B.n633 B.n632 585
R750 B.n632 B.n631 585
R751 B.n266 B.n265 585
R752 B.n267 B.n266 585
R753 B.n624 B.n623 585
R754 B.n625 B.n624 585
R755 B.n622 B.n272 585
R756 B.n272 B.n271 585
R757 B.n621 B.n620 585
R758 B.n620 B.n619 585
R759 B.n274 B.n273 585
R760 B.n612 B.n274 585
R761 B.n611 B.n610 585
R762 B.n613 B.n611 585
R763 B.n609 B.n279 585
R764 B.n279 B.n278 585
R765 B.n608 B.n607 585
R766 B.n607 B.n606 585
R767 B.n281 B.n280 585
R768 B.n282 B.n281 585
R769 B.n599 B.n598 585
R770 B.n600 B.n599 585
R771 B.n597 B.n287 585
R772 B.n287 B.n286 585
R773 B.n596 B.n595 585
R774 B.n595 B.n594 585
R775 B.n289 B.n288 585
R776 B.n587 B.n289 585
R777 B.n586 B.n585 585
R778 B.n588 B.n586 585
R779 B.n584 B.n294 585
R780 B.n294 B.n293 585
R781 B.n583 B.n582 585
R782 B.n582 B.n581 585
R783 B.n296 B.n295 585
R784 B.n297 B.n296 585
R785 B.n574 B.n573 585
R786 B.n575 B.n574 585
R787 B.n572 B.n302 585
R788 B.n302 B.n301 585
R789 B.n571 B.n570 585
R790 B.n570 B.n569 585
R791 B.n304 B.n303 585
R792 B.n305 B.n304 585
R793 B.n562 B.n561 585
R794 B.n563 B.n562 585
R795 B.n560 B.n310 585
R796 B.n310 B.n309 585
R797 B.n559 B.n558 585
R798 B.n558 B.n557 585
R799 B.n312 B.n311 585
R800 B.n313 B.n312 585
R801 B.n550 B.n549 585
R802 B.n551 B.n550 585
R803 B.n548 B.n318 585
R804 B.n318 B.n317 585
R805 B.n547 B.n546 585
R806 B.n546 B.n545 585
R807 B.n320 B.n319 585
R808 B.n321 B.n320 585
R809 B.n538 B.n537 585
R810 B.n539 B.n538 585
R811 B.n536 B.n326 585
R812 B.n326 B.n325 585
R813 B.n535 B.n534 585
R814 B.n534 B.n533 585
R815 B.n328 B.n327 585
R816 B.n329 B.n328 585
R817 B.n526 B.n525 585
R818 B.n527 B.n526 585
R819 B.n524 B.n334 585
R820 B.n334 B.n333 585
R821 B.n523 B.n522 585
R822 B.n522 B.n521 585
R823 B.n336 B.n335 585
R824 B.n337 B.n336 585
R825 B.n514 B.n513 585
R826 B.n515 B.n514 585
R827 B.n512 B.n342 585
R828 B.n342 B.n341 585
R829 B.n511 B.n510 585
R830 B.n510 B.n509 585
R831 B.n344 B.n343 585
R832 B.n345 B.n344 585
R833 B.n505 B.n504 585
R834 B.n348 B.n347 585
R835 B.n501 B.n500 585
R836 B.n502 B.n501 585
R837 B.n499 B.n378 585
R838 B.n498 B.n497 585
R839 B.n496 B.n495 585
R840 B.n494 B.n493 585
R841 B.n492 B.n491 585
R842 B.n490 B.n489 585
R843 B.n488 B.n487 585
R844 B.n486 B.n485 585
R845 B.n484 B.n483 585
R846 B.n482 B.n481 585
R847 B.n480 B.n479 585
R848 B.n478 B.n477 585
R849 B.n476 B.n475 585
R850 B.n474 B.n473 585
R851 B.n472 B.n471 585
R852 B.n470 B.n469 585
R853 B.n468 B.n467 585
R854 B.n466 B.n465 585
R855 B.n464 B.n463 585
R856 B.n462 B.n461 585
R857 B.n460 B.n459 585
R858 B.n458 B.n457 585
R859 B.n456 B.n455 585
R860 B.n453 B.n452 585
R861 B.n451 B.n450 585
R862 B.n449 B.n448 585
R863 B.n447 B.n446 585
R864 B.n445 B.n444 585
R865 B.n443 B.n442 585
R866 B.n441 B.n440 585
R867 B.n439 B.n438 585
R868 B.n437 B.n436 585
R869 B.n435 B.n434 585
R870 B.n433 B.n432 585
R871 B.n431 B.n430 585
R872 B.n429 B.n428 585
R873 B.n427 B.n426 585
R874 B.n425 B.n424 585
R875 B.n423 B.n422 585
R876 B.n421 B.n420 585
R877 B.n419 B.n418 585
R878 B.n417 B.n416 585
R879 B.n415 B.n414 585
R880 B.n413 B.n412 585
R881 B.n411 B.n410 585
R882 B.n409 B.n408 585
R883 B.n407 B.n406 585
R884 B.n405 B.n404 585
R885 B.n403 B.n402 585
R886 B.n401 B.n400 585
R887 B.n399 B.n398 585
R888 B.n397 B.n396 585
R889 B.n395 B.n394 585
R890 B.n393 B.n392 585
R891 B.n391 B.n390 585
R892 B.n389 B.n388 585
R893 B.n387 B.n386 585
R894 B.n385 B.n384 585
R895 B.n506 B.n346 585
R896 B.n346 B.n345 585
R897 B.n508 B.n507 585
R898 B.n509 B.n508 585
R899 B.n340 B.n339 585
R900 B.n341 B.n340 585
R901 B.n517 B.n516 585
R902 B.n516 B.n515 585
R903 B.n518 B.n338 585
R904 B.n338 B.n337 585
R905 B.n520 B.n519 585
R906 B.n521 B.n520 585
R907 B.n332 B.n331 585
R908 B.n333 B.n332 585
R909 B.n529 B.n528 585
R910 B.n528 B.n527 585
R911 B.n530 B.n330 585
R912 B.n330 B.n329 585
R913 B.n532 B.n531 585
R914 B.n533 B.n532 585
R915 B.n324 B.n323 585
R916 B.n325 B.n324 585
R917 B.n541 B.n540 585
R918 B.n540 B.n539 585
R919 B.n542 B.n322 585
R920 B.n322 B.n321 585
R921 B.n544 B.n543 585
R922 B.n545 B.n544 585
R923 B.n316 B.n315 585
R924 B.n317 B.n316 585
R925 B.n553 B.n552 585
R926 B.n552 B.n551 585
R927 B.n554 B.n314 585
R928 B.n314 B.n313 585
R929 B.n556 B.n555 585
R930 B.n557 B.n556 585
R931 B.n308 B.n307 585
R932 B.n309 B.n308 585
R933 B.n565 B.n564 585
R934 B.n564 B.n563 585
R935 B.n566 B.n306 585
R936 B.n306 B.n305 585
R937 B.n568 B.n567 585
R938 B.n569 B.n568 585
R939 B.n300 B.n299 585
R940 B.n301 B.n300 585
R941 B.n577 B.n576 585
R942 B.n576 B.n575 585
R943 B.n578 B.n298 585
R944 B.n298 B.n297 585
R945 B.n580 B.n579 585
R946 B.n581 B.n580 585
R947 B.n292 B.n291 585
R948 B.n293 B.n292 585
R949 B.n590 B.n589 585
R950 B.n589 B.n588 585
R951 B.n591 B.n290 585
R952 B.n587 B.n290 585
R953 B.n593 B.n592 585
R954 B.n594 B.n593 585
R955 B.n285 B.n284 585
R956 B.n286 B.n285 585
R957 B.n602 B.n601 585
R958 B.n601 B.n600 585
R959 B.n603 B.n283 585
R960 B.n283 B.n282 585
R961 B.n605 B.n604 585
R962 B.n606 B.n605 585
R963 B.n277 B.n276 585
R964 B.n278 B.n277 585
R965 B.n615 B.n614 585
R966 B.n614 B.n613 585
R967 B.n616 B.n275 585
R968 B.n612 B.n275 585
R969 B.n618 B.n617 585
R970 B.n619 B.n618 585
R971 B.n270 B.n269 585
R972 B.n271 B.n270 585
R973 B.n627 B.n626 585
R974 B.n626 B.n625 585
R975 B.n628 B.n268 585
R976 B.n268 B.n267 585
R977 B.n630 B.n629 585
R978 B.n631 B.n630 585
R979 B.n262 B.n261 585
R980 B.n263 B.n262 585
R981 B.n639 B.n638 585
R982 B.n638 B.n637 585
R983 B.n640 B.n260 585
R984 B.n260 B.n259 585
R985 B.n642 B.n641 585
R986 B.n643 B.n642 585
R987 B.n254 B.n253 585
R988 B.n255 B.n254 585
R989 B.n652 B.n651 585
R990 B.n651 B.n650 585
R991 B.n653 B.n252 585
R992 B.n252 B.n251 585
R993 B.n655 B.n654 585
R994 B.n656 B.n655 585
R995 B.n3 B.n0 585
R996 B.n4 B.n3 585
R997 B.n831 B.n1 585
R998 B.n832 B.n831 585
R999 B.n830 B.n829 585
R1000 B.n830 B.n8 585
R1001 B.n828 B.n9 585
R1002 B.n12 B.n9 585
R1003 B.n827 B.n826 585
R1004 B.n826 B.n825 585
R1005 B.n11 B.n10 585
R1006 B.n824 B.n11 585
R1007 B.n822 B.n821 585
R1008 B.n823 B.n822 585
R1009 B.n820 B.n17 585
R1010 B.n17 B.n16 585
R1011 B.n819 B.n818 585
R1012 B.n818 B.n817 585
R1013 B.n19 B.n18 585
R1014 B.n816 B.n19 585
R1015 B.n814 B.n813 585
R1016 B.n815 B.n814 585
R1017 B.n812 B.n24 585
R1018 B.n24 B.n23 585
R1019 B.n811 B.n810 585
R1020 B.n810 B.n809 585
R1021 B.n26 B.n25 585
R1022 B.n808 B.n26 585
R1023 B.n806 B.n805 585
R1024 B.n807 B.n806 585
R1025 B.n804 B.n30 585
R1026 B.n33 B.n30 585
R1027 B.n803 B.n802 585
R1028 B.n802 B.n801 585
R1029 B.n32 B.n31 585
R1030 B.n800 B.n32 585
R1031 B.n798 B.n797 585
R1032 B.n799 B.n798 585
R1033 B.n796 B.n38 585
R1034 B.n38 B.n37 585
R1035 B.n795 B.n794 585
R1036 B.n794 B.n793 585
R1037 B.n40 B.n39 585
R1038 B.n792 B.n40 585
R1039 B.n790 B.n789 585
R1040 B.n791 B.n790 585
R1041 B.n788 B.n44 585
R1042 B.n47 B.n44 585
R1043 B.n787 B.n786 585
R1044 B.n786 B.n785 585
R1045 B.n46 B.n45 585
R1046 B.n784 B.n46 585
R1047 B.n782 B.n781 585
R1048 B.n783 B.n782 585
R1049 B.n780 B.n52 585
R1050 B.n52 B.n51 585
R1051 B.n779 B.n778 585
R1052 B.n778 B.n777 585
R1053 B.n54 B.n53 585
R1054 B.n776 B.n54 585
R1055 B.n774 B.n773 585
R1056 B.n775 B.n774 585
R1057 B.n772 B.n59 585
R1058 B.n59 B.n58 585
R1059 B.n771 B.n770 585
R1060 B.n770 B.n769 585
R1061 B.n61 B.n60 585
R1062 B.n768 B.n61 585
R1063 B.n766 B.n765 585
R1064 B.n767 B.n766 585
R1065 B.n764 B.n66 585
R1066 B.n66 B.n65 585
R1067 B.n763 B.n762 585
R1068 B.n762 B.n761 585
R1069 B.n68 B.n67 585
R1070 B.n760 B.n68 585
R1071 B.n758 B.n757 585
R1072 B.n759 B.n758 585
R1073 B.n756 B.n73 585
R1074 B.n73 B.n72 585
R1075 B.n755 B.n754 585
R1076 B.n754 B.n753 585
R1077 B.n75 B.n74 585
R1078 B.n752 B.n75 585
R1079 B.n750 B.n749 585
R1080 B.n751 B.n750 585
R1081 B.n748 B.n80 585
R1082 B.n80 B.n79 585
R1083 B.n747 B.n746 585
R1084 B.n746 B.n745 585
R1085 B.n82 B.n81 585
R1086 B.n744 B.n82 585
R1087 B.n742 B.n741 585
R1088 B.n743 B.n742 585
R1089 B.n740 B.n87 585
R1090 B.n87 B.n86 585
R1091 B.n739 B.n738 585
R1092 B.n738 B.n737 585
R1093 B.n89 B.n88 585
R1094 B.n736 B.n89 585
R1095 B.n734 B.n733 585
R1096 B.n735 B.n734 585
R1097 B.n732 B.n94 585
R1098 B.n94 B.n93 585
R1099 B.n835 B.n834 585
R1100 B.n833 B.n2 585
R1101 B.n730 B.n94 574.183
R1102 B.n727 B.n127 574.183
R1103 B.n384 B.n344 574.183
R1104 B.n504 B.n346 574.183
R1105 B.n130 B.t12 268.813
R1106 B.n128 B.t19 268.813
R1107 B.n381 B.t16 268.813
R1108 B.n379 B.t8 268.813
R1109 B.n728 B.n125 256.663
R1110 B.n728 B.n124 256.663
R1111 B.n728 B.n123 256.663
R1112 B.n728 B.n122 256.663
R1113 B.n728 B.n121 256.663
R1114 B.n728 B.n120 256.663
R1115 B.n728 B.n119 256.663
R1116 B.n728 B.n118 256.663
R1117 B.n728 B.n117 256.663
R1118 B.n728 B.n116 256.663
R1119 B.n728 B.n115 256.663
R1120 B.n728 B.n114 256.663
R1121 B.n728 B.n113 256.663
R1122 B.n728 B.n112 256.663
R1123 B.n728 B.n111 256.663
R1124 B.n728 B.n110 256.663
R1125 B.n728 B.n109 256.663
R1126 B.n728 B.n108 256.663
R1127 B.n728 B.n107 256.663
R1128 B.n728 B.n106 256.663
R1129 B.n728 B.n105 256.663
R1130 B.n728 B.n104 256.663
R1131 B.n728 B.n103 256.663
R1132 B.n728 B.n102 256.663
R1133 B.n728 B.n101 256.663
R1134 B.n728 B.n100 256.663
R1135 B.n728 B.n99 256.663
R1136 B.n728 B.n98 256.663
R1137 B.n728 B.n97 256.663
R1138 B.n729 B.n728 256.663
R1139 B.n503 B.n502 256.663
R1140 B.n502 B.n349 256.663
R1141 B.n502 B.n350 256.663
R1142 B.n502 B.n351 256.663
R1143 B.n502 B.n352 256.663
R1144 B.n502 B.n353 256.663
R1145 B.n502 B.n354 256.663
R1146 B.n502 B.n355 256.663
R1147 B.n502 B.n356 256.663
R1148 B.n502 B.n357 256.663
R1149 B.n502 B.n358 256.663
R1150 B.n502 B.n359 256.663
R1151 B.n502 B.n360 256.663
R1152 B.n502 B.n361 256.663
R1153 B.n502 B.n362 256.663
R1154 B.n502 B.n363 256.663
R1155 B.n502 B.n364 256.663
R1156 B.n502 B.n365 256.663
R1157 B.n502 B.n366 256.663
R1158 B.n502 B.n367 256.663
R1159 B.n502 B.n368 256.663
R1160 B.n502 B.n369 256.663
R1161 B.n502 B.n370 256.663
R1162 B.n502 B.n371 256.663
R1163 B.n502 B.n372 256.663
R1164 B.n502 B.n373 256.663
R1165 B.n502 B.n374 256.663
R1166 B.n502 B.n375 256.663
R1167 B.n502 B.n376 256.663
R1168 B.n502 B.n377 256.663
R1169 B.n837 B.n836 256.663
R1170 B.n128 B.t20 247.683
R1171 B.n381 B.t18 247.683
R1172 B.n130 B.t14 247.683
R1173 B.n379 B.t11 247.683
R1174 B.n129 B.t21 190.083
R1175 B.n382 B.t17 190.083
R1176 B.n131 B.t15 190.083
R1177 B.n380 B.t10 190.083
R1178 B.n133 B.n96 163.367
R1179 B.n137 B.n136 163.367
R1180 B.n141 B.n140 163.367
R1181 B.n145 B.n144 163.367
R1182 B.n149 B.n148 163.367
R1183 B.n153 B.n152 163.367
R1184 B.n157 B.n156 163.367
R1185 B.n161 B.n160 163.367
R1186 B.n165 B.n164 163.367
R1187 B.n169 B.n168 163.367
R1188 B.n173 B.n172 163.367
R1189 B.n177 B.n176 163.367
R1190 B.n181 B.n180 163.367
R1191 B.n185 B.n184 163.367
R1192 B.n189 B.n188 163.367
R1193 B.n193 B.n192 163.367
R1194 B.n197 B.n196 163.367
R1195 B.n202 B.n201 163.367
R1196 B.n206 B.n205 163.367
R1197 B.n210 B.n209 163.367
R1198 B.n214 B.n213 163.367
R1199 B.n218 B.n217 163.367
R1200 B.n222 B.n221 163.367
R1201 B.n226 B.n225 163.367
R1202 B.n230 B.n229 163.367
R1203 B.n234 B.n233 163.367
R1204 B.n238 B.n237 163.367
R1205 B.n242 B.n241 163.367
R1206 B.n246 B.n245 163.367
R1207 B.n727 B.n126 163.367
R1208 B.n510 B.n344 163.367
R1209 B.n510 B.n342 163.367
R1210 B.n514 B.n342 163.367
R1211 B.n514 B.n336 163.367
R1212 B.n522 B.n336 163.367
R1213 B.n522 B.n334 163.367
R1214 B.n526 B.n334 163.367
R1215 B.n526 B.n328 163.367
R1216 B.n534 B.n328 163.367
R1217 B.n534 B.n326 163.367
R1218 B.n538 B.n326 163.367
R1219 B.n538 B.n320 163.367
R1220 B.n546 B.n320 163.367
R1221 B.n546 B.n318 163.367
R1222 B.n550 B.n318 163.367
R1223 B.n550 B.n312 163.367
R1224 B.n558 B.n312 163.367
R1225 B.n558 B.n310 163.367
R1226 B.n562 B.n310 163.367
R1227 B.n562 B.n304 163.367
R1228 B.n570 B.n304 163.367
R1229 B.n570 B.n302 163.367
R1230 B.n574 B.n302 163.367
R1231 B.n574 B.n296 163.367
R1232 B.n582 B.n296 163.367
R1233 B.n582 B.n294 163.367
R1234 B.n586 B.n294 163.367
R1235 B.n586 B.n289 163.367
R1236 B.n595 B.n289 163.367
R1237 B.n595 B.n287 163.367
R1238 B.n599 B.n287 163.367
R1239 B.n599 B.n281 163.367
R1240 B.n607 B.n281 163.367
R1241 B.n607 B.n279 163.367
R1242 B.n611 B.n279 163.367
R1243 B.n611 B.n274 163.367
R1244 B.n620 B.n274 163.367
R1245 B.n620 B.n272 163.367
R1246 B.n624 B.n272 163.367
R1247 B.n624 B.n266 163.367
R1248 B.n632 B.n266 163.367
R1249 B.n632 B.n264 163.367
R1250 B.n636 B.n264 163.367
R1251 B.n636 B.n258 163.367
R1252 B.n644 B.n258 163.367
R1253 B.n644 B.n256 163.367
R1254 B.n649 B.n256 163.367
R1255 B.n649 B.n250 163.367
R1256 B.n657 B.n250 163.367
R1257 B.n658 B.n657 163.367
R1258 B.n658 B.n5 163.367
R1259 B.n6 B.n5 163.367
R1260 B.n7 B.n6 163.367
R1261 B.n664 B.n7 163.367
R1262 B.n665 B.n664 163.367
R1263 B.n665 B.n13 163.367
R1264 B.n14 B.n13 163.367
R1265 B.n15 B.n14 163.367
R1266 B.n670 B.n15 163.367
R1267 B.n670 B.n20 163.367
R1268 B.n21 B.n20 163.367
R1269 B.n22 B.n21 163.367
R1270 B.n675 B.n22 163.367
R1271 B.n675 B.n27 163.367
R1272 B.n28 B.n27 163.367
R1273 B.n29 B.n28 163.367
R1274 B.n680 B.n29 163.367
R1275 B.n680 B.n34 163.367
R1276 B.n35 B.n34 163.367
R1277 B.n36 B.n35 163.367
R1278 B.n685 B.n36 163.367
R1279 B.n685 B.n41 163.367
R1280 B.n42 B.n41 163.367
R1281 B.n43 B.n42 163.367
R1282 B.n690 B.n43 163.367
R1283 B.n690 B.n48 163.367
R1284 B.n49 B.n48 163.367
R1285 B.n50 B.n49 163.367
R1286 B.n695 B.n50 163.367
R1287 B.n695 B.n55 163.367
R1288 B.n56 B.n55 163.367
R1289 B.n57 B.n56 163.367
R1290 B.n700 B.n57 163.367
R1291 B.n700 B.n62 163.367
R1292 B.n63 B.n62 163.367
R1293 B.n64 B.n63 163.367
R1294 B.n705 B.n64 163.367
R1295 B.n705 B.n69 163.367
R1296 B.n70 B.n69 163.367
R1297 B.n71 B.n70 163.367
R1298 B.n710 B.n71 163.367
R1299 B.n710 B.n76 163.367
R1300 B.n77 B.n76 163.367
R1301 B.n78 B.n77 163.367
R1302 B.n715 B.n78 163.367
R1303 B.n715 B.n83 163.367
R1304 B.n84 B.n83 163.367
R1305 B.n85 B.n84 163.367
R1306 B.n720 B.n85 163.367
R1307 B.n720 B.n90 163.367
R1308 B.n91 B.n90 163.367
R1309 B.n92 B.n91 163.367
R1310 B.n127 B.n92 163.367
R1311 B.n501 B.n348 163.367
R1312 B.n501 B.n378 163.367
R1313 B.n497 B.n496 163.367
R1314 B.n493 B.n492 163.367
R1315 B.n489 B.n488 163.367
R1316 B.n485 B.n484 163.367
R1317 B.n481 B.n480 163.367
R1318 B.n477 B.n476 163.367
R1319 B.n473 B.n472 163.367
R1320 B.n469 B.n468 163.367
R1321 B.n465 B.n464 163.367
R1322 B.n461 B.n460 163.367
R1323 B.n457 B.n456 163.367
R1324 B.n452 B.n451 163.367
R1325 B.n448 B.n447 163.367
R1326 B.n444 B.n443 163.367
R1327 B.n440 B.n439 163.367
R1328 B.n436 B.n435 163.367
R1329 B.n432 B.n431 163.367
R1330 B.n428 B.n427 163.367
R1331 B.n424 B.n423 163.367
R1332 B.n420 B.n419 163.367
R1333 B.n416 B.n415 163.367
R1334 B.n412 B.n411 163.367
R1335 B.n408 B.n407 163.367
R1336 B.n404 B.n403 163.367
R1337 B.n400 B.n399 163.367
R1338 B.n396 B.n395 163.367
R1339 B.n392 B.n391 163.367
R1340 B.n388 B.n387 163.367
R1341 B.n508 B.n346 163.367
R1342 B.n508 B.n340 163.367
R1343 B.n516 B.n340 163.367
R1344 B.n516 B.n338 163.367
R1345 B.n520 B.n338 163.367
R1346 B.n520 B.n332 163.367
R1347 B.n528 B.n332 163.367
R1348 B.n528 B.n330 163.367
R1349 B.n532 B.n330 163.367
R1350 B.n532 B.n324 163.367
R1351 B.n540 B.n324 163.367
R1352 B.n540 B.n322 163.367
R1353 B.n544 B.n322 163.367
R1354 B.n544 B.n316 163.367
R1355 B.n552 B.n316 163.367
R1356 B.n552 B.n314 163.367
R1357 B.n556 B.n314 163.367
R1358 B.n556 B.n308 163.367
R1359 B.n564 B.n308 163.367
R1360 B.n564 B.n306 163.367
R1361 B.n568 B.n306 163.367
R1362 B.n568 B.n300 163.367
R1363 B.n576 B.n300 163.367
R1364 B.n576 B.n298 163.367
R1365 B.n580 B.n298 163.367
R1366 B.n580 B.n292 163.367
R1367 B.n589 B.n292 163.367
R1368 B.n589 B.n290 163.367
R1369 B.n593 B.n290 163.367
R1370 B.n593 B.n285 163.367
R1371 B.n601 B.n285 163.367
R1372 B.n601 B.n283 163.367
R1373 B.n605 B.n283 163.367
R1374 B.n605 B.n277 163.367
R1375 B.n614 B.n277 163.367
R1376 B.n614 B.n275 163.367
R1377 B.n618 B.n275 163.367
R1378 B.n618 B.n270 163.367
R1379 B.n626 B.n270 163.367
R1380 B.n626 B.n268 163.367
R1381 B.n630 B.n268 163.367
R1382 B.n630 B.n262 163.367
R1383 B.n638 B.n262 163.367
R1384 B.n638 B.n260 163.367
R1385 B.n642 B.n260 163.367
R1386 B.n642 B.n254 163.367
R1387 B.n651 B.n254 163.367
R1388 B.n651 B.n252 163.367
R1389 B.n655 B.n252 163.367
R1390 B.n655 B.n3 163.367
R1391 B.n835 B.n3 163.367
R1392 B.n831 B.n2 163.367
R1393 B.n831 B.n830 163.367
R1394 B.n830 B.n9 163.367
R1395 B.n826 B.n9 163.367
R1396 B.n826 B.n11 163.367
R1397 B.n822 B.n11 163.367
R1398 B.n822 B.n17 163.367
R1399 B.n818 B.n17 163.367
R1400 B.n818 B.n19 163.367
R1401 B.n814 B.n19 163.367
R1402 B.n814 B.n24 163.367
R1403 B.n810 B.n24 163.367
R1404 B.n810 B.n26 163.367
R1405 B.n806 B.n26 163.367
R1406 B.n806 B.n30 163.367
R1407 B.n802 B.n30 163.367
R1408 B.n802 B.n32 163.367
R1409 B.n798 B.n32 163.367
R1410 B.n798 B.n38 163.367
R1411 B.n794 B.n38 163.367
R1412 B.n794 B.n40 163.367
R1413 B.n790 B.n40 163.367
R1414 B.n790 B.n44 163.367
R1415 B.n786 B.n44 163.367
R1416 B.n786 B.n46 163.367
R1417 B.n782 B.n46 163.367
R1418 B.n782 B.n52 163.367
R1419 B.n778 B.n52 163.367
R1420 B.n778 B.n54 163.367
R1421 B.n774 B.n54 163.367
R1422 B.n774 B.n59 163.367
R1423 B.n770 B.n59 163.367
R1424 B.n770 B.n61 163.367
R1425 B.n766 B.n61 163.367
R1426 B.n766 B.n66 163.367
R1427 B.n762 B.n66 163.367
R1428 B.n762 B.n68 163.367
R1429 B.n758 B.n68 163.367
R1430 B.n758 B.n73 163.367
R1431 B.n754 B.n73 163.367
R1432 B.n754 B.n75 163.367
R1433 B.n750 B.n75 163.367
R1434 B.n750 B.n80 163.367
R1435 B.n746 B.n80 163.367
R1436 B.n746 B.n82 163.367
R1437 B.n742 B.n82 163.367
R1438 B.n742 B.n87 163.367
R1439 B.n738 B.n87 163.367
R1440 B.n738 B.n89 163.367
R1441 B.n734 B.n89 163.367
R1442 B.n734 B.n94 163.367
R1443 B.n502 B.n345 131.909
R1444 B.n728 B.n93 131.909
R1445 B.n730 B.n729 71.676
R1446 B.n133 B.n97 71.676
R1447 B.n137 B.n98 71.676
R1448 B.n141 B.n99 71.676
R1449 B.n145 B.n100 71.676
R1450 B.n149 B.n101 71.676
R1451 B.n153 B.n102 71.676
R1452 B.n157 B.n103 71.676
R1453 B.n161 B.n104 71.676
R1454 B.n165 B.n105 71.676
R1455 B.n169 B.n106 71.676
R1456 B.n173 B.n107 71.676
R1457 B.n177 B.n108 71.676
R1458 B.n181 B.n109 71.676
R1459 B.n185 B.n110 71.676
R1460 B.n189 B.n111 71.676
R1461 B.n193 B.n112 71.676
R1462 B.n197 B.n113 71.676
R1463 B.n202 B.n114 71.676
R1464 B.n206 B.n115 71.676
R1465 B.n210 B.n116 71.676
R1466 B.n214 B.n117 71.676
R1467 B.n218 B.n118 71.676
R1468 B.n222 B.n119 71.676
R1469 B.n226 B.n120 71.676
R1470 B.n230 B.n121 71.676
R1471 B.n234 B.n122 71.676
R1472 B.n238 B.n123 71.676
R1473 B.n242 B.n124 71.676
R1474 B.n246 B.n125 71.676
R1475 B.n126 B.n125 71.676
R1476 B.n245 B.n124 71.676
R1477 B.n241 B.n123 71.676
R1478 B.n237 B.n122 71.676
R1479 B.n233 B.n121 71.676
R1480 B.n229 B.n120 71.676
R1481 B.n225 B.n119 71.676
R1482 B.n221 B.n118 71.676
R1483 B.n217 B.n117 71.676
R1484 B.n213 B.n116 71.676
R1485 B.n209 B.n115 71.676
R1486 B.n205 B.n114 71.676
R1487 B.n201 B.n113 71.676
R1488 B.n196 B.n112 71.676
R1489 B.n192 B.n111 71.676
R1490 B.n188 B.n110 71.676
R1491 B.n184 B.n109 71.676
R1492 B.n180 B.n108 71.676
R1493 B.n176 B.n107 71.676
R1494 B.n172 B.n106 71.676
R1495 B.n168 B.n105 71.676
R1496 B.n164 B.n104 71.676
R1497 B.n160 B.n103 71.676
R1498 B.n156 B.n102 71.676
R1499 B.n152 B.n101 71.676
R1500 B.n148 B.n100 71.676
R1501 B.n144 B.n99 71.676
R1502 B.n140 B.n98 71.676
R1503 B.n136 B.n97 71.676
R1504 B.n729 B.n96 71.676
R1505 B.n504 B.n503 71.676
R1506 B.n378 B.n349 71.676
R1507 B.n496 B.n350 71.676
R1508 B.n492 B.n351 71.676
R1509 B.n488 B.n352 71.676
R1510 B.n484 B.n353 71.676
R1511 B.n480 B.n354 71.676
R1512 B.n476 B.n355 71.676
R1513 B.n472 B.n356 71.676
R1514 B.n468 B.n357 71.676
R1515 B.n464 B.n358 71.676
R1516 B.n460 B.n359 71.676
R1517 B.n456 B.n360 71.676
R1518 B.n451 B.n361 71.676
R1519 B.n447 B.n362 71.676
R1520 B.n443 B.n363 71.676
R1521 B.n439 B.n364 71.676
R1522 B.n435 B.n365 71.676
R1523 B.n431 B.n366 71.676
R1524 B.n427 B.n367 71.676
R1525 B.n423 B.n368 71.676
R1526 B.n419 B.n369 71.676
R1527 B.n415 B.n370 71.676
R1528 B.n411 B.n371 71.676
R1529 B.n407 B.n372 71.676
R1530 B.n403 B.n373 71.676
R1531 B.n399 B.n374 71.676
R1532 B.n395 B.n375 71.676
R1533 B.n391 B.n376 71.676
R1534 B.n387 B.n377 71.676
R1535 B.n503 B.n348 71.676
R1536 B.n497 B.n349 71.676
R1537 B.n493 B.n350 71.676
R1538 B.n489 B.n351 71.676
R1539 B.n485 B.n352 71.676
R1540 B.n481 B.n353 71.676
R1541 B.n477 B.n354 71.676
R1542 B.n473 B.n355 71.676
R1543 B.n469 B.n356 71.676
R1544 B.n465 B.n357 71.676
R1545 B.n461 B.n358 71.676
R1546 B.n457 B.n359 71.676
R1547 B.n452 B.n360 71.676
R1548 B.n448 B.n361 71.676
R1549 B.n444 B.n362 71.676
R1550 B.n440 B.n363 71.676
R1551 B.n436 B.n364 71.676
R1552 B.n432 B.n365 71.676
R1553 B.n428 B.n366 71.676
R1554 B.n424 B.n367 71.676
R1555 B.n420 B.n368 71.676
R1556 B.n416 B.n369 71.676
R1557 B.n412 B.n370 71.676
R1558 B.n408 B.n371 71.676
R1559 B.n404 B.n372 71.676
R1560 B.n400 B.n373 71.676
R1561 B.n396 B.n374 71.676
R1562 B.n392 B.n375 71.676
R1563 B.n388 B.n376 71.676
R1564 B.n384 B.n377 71.676
R1565 B.n836 B.n835 71.676
R1566 B.n836 B.n2 71.676
R1567 B.n509 B.n345 62.7259
R1568 B.n509 B.n341 62.7259
R1569 B.n515 B.n341 62.7259
R1570 B.n515 B.n337 62.7259
R1571 B.n521 B.n337 62.7259
R1572 B.n521 B.n333 62.7259
R1573 B.n527 B.n333 62.7259
R1574 B.n533 B.n329 62.7259
R1575 B.n533 B.n325 62.7259
R1576 B.n539 B.n325 62.7259
R1577 B.n539 B.n321 62.7259
R1578 B.n545 B.n321 62.7259
R1579 B.n545 B.n317 62.7259
R1580 B.n551 B.n317 62.7259
R1581 B.n551 B.n313 62.7259
R1582 B.n557 B.n313 62.7259
R1583 B.n557 B.n309 62.7259
R1584 B.n563 B.n309 62.7259
R1585 B.n569 B.n305 62.7259
R1586 B.n569 B.n301 62.7259
R1587 B.n575 B.n301 62.7259
R1588 B.n575 B.n297 62.7259
R1589 B.n581 B.n297 62.7259
R1590 B.n581 B.n293 62.7259
R1591 B.n588 B.n293 62.7259
R1592 B.n588 B.n587 62.7259
R1593 B.n594 B.n286 62.7259
R1594 B.n600 B.n286 62.7259
R1595 B.n600 B.n282 62.7259
R1596 B.n606 B.n282 62.7259
R1597 B.n606 B.n278 62.7259
R1598 B.n613 B.n278 62.7259
R1599 B.n613 B.n612 62.7259
R1600 B.n619 B.n271 62.7259
R1601 B.n625 B.n271 62.7259
R1602 B.n625 B.n267 62.7259
R1603 B.n631 B.n267 62.7259
R1604 B.n631 B.n263 62.7259
R1605 B.n637 B.n263 62.7259
R1606 B.n637 B.n259 62.7259
R1607 B.n643 B.n259 62.7259
R1608 B.n650 B.n255 62.7259
R1609 B.n650 B.n251 62.7259
R1610 B.n656 B.n251 62.7259
R1611 B.n656 B.n4 62.7259
R1612 B.n834 B.n4 62.7259
R1613 B.n834 B.n833 62.7259
R1614 B.n833 B.n832 62.7259
R1615 B.n832 B.n8 62.7259
R1616 B.n12 B.n8 62.7259
R1617 B.n825 B.n12 62.7259
R1618 B.n825 B.n824 62.7259
R1619 B.n823 B.n16 62.7259
R1620 B.n817 B.n16 62.7259
R1621 B.n817 B.n816 62.7259
R1622 B.n816 B.n815 62.7259
R1623 B.n815 B.n23 62.7259
R1624 B.n809 B.n23 62.7259
R1625 B.n809 B.n808 62.7259
R1626 B.n808 B.n807 62.7259
R1627 B.n801 B.n33 62.7259
R1628 B.n801 B.n800 62.7259
R1629 B.n800 B.n799 62.7259
R1630 B.n799 B.n37 62.7259
R1631 B.n793 B.n37 62.7259
R1632 B.n793 B.n792 62.7259
R1633 B.n792 B.n791 62.7259
R1634 B.n785 B.n47 62.7259
R1635 B.n785 B.n784 62.7259
R1636 B.n784 B.n783 62.7259
R1637 B.n783 B.n51 62.7259
R1638 B.n777 B.n51 62.7259
R1639 B.n777 B.n776 62.7259
R1640 B.n776 B.n775 62.7259
R1641 B.n775 B.n58 62.7259
R1642 B.n769 B.n768 62.7259
R1643 B.n768 B.n767 62.7259
R1644 B.n767 B.n65 62.7259
R1645 B.n761 B.n65 62.7259
R1646 B.n761 B.n760 62.7259
R1647 B.n760 B.n759 62.7259
R1648 B.n759 B.n72 62.7259
R1649 B.n753 B.n72 62.7259
R1650 B.n753 B.n752 62.7259
R1651 B.n752 B.n751 62.7259
R1652 B.n751 B.n79 62.7259
R1653 B.n745 B.n744 62.7259
R1654 B.n744 B.n743 62.7259
R1655 B.n743 B.n86 62.7259
R1656 B.n737 B.n86 62.7259
R1657 B.n737 B.n736 62.7259
R1658 B.n736 B.n735 62.7259
R1659 B.n735 B.n93 62.7259
R1660 B.n132 B.n131 59.5399
R1661 B.n199 B.n129 59.5399
R1662 B.n383 B.n382 59.5399
R1663 B.n454 B.n380 59.5399
R1664 B.n594 B.t1 59.0361
R1665 B.n791 B.t0 59.0361
R1666 B.n131 B.n130 57.6005
R1667 B.n129 B.n128 57.6005
R1668 B.n382 B.n381 57.6005
R1669 B.n380 B.n379 57.6005
R1670 B.n612 B.t7 49.8118
R1671 B.n33 B.t5 49.8118
R1672 B.t6 B.n305 42.4324
R1673 B.t2 B.n58 42.4324
R1674 B.t9 B.n329 38.7426
R1675 B.t13 B.n79 38.7426
R1676 B.n506 B.n505 37.3078
R1677 B.n385 B.n343 37.3078
R1678 B.n726 B.n725 37.3078
R1679 B.n732 B.n731 37.3078
R1680 B.n643 B.t4 33.208
R1681 B.t3 B.n823 33.208
R1682 B.t4 B.n255 29.5183
R1683 B.n824 B.t3 29.5183
R1684 B.n527 B.t9 23.9837
R1685 B.n745 B.t13 23.9837
R1686 B.n563 B.t6 20.294
R1687 B.n769 B.t2 20.294
R1688 B B.n837 18.0485
R1689 B.n619 B.t7 12.9145
R1690 B.n807 B.t5 12.9145
R1691 B.n507 B.n506 10.6151
R1692 B.n507 B.n339 10.6151
R1693 B.n517 B.n339 10.6151
R1694 B.n518 B.n517 10.6151
R1695 B.n519 B.n518 10.6151
R1696 B.n519 B.n331 10.6151
R1697 B.n529 B.n331 10.6151
R1698 B.n530 B.n529 10.6151
R1699 B.n531 B.n530 10.6151
R1700 B.n531 B.n323 10.6151
R1701 B.n541 B.n323 10.6151
R1702 B.n542 B.n541 10.6151
R1703 B.n543 B.n542 10.6151
R1704 B.n543 B.n315 10.6151
R1705 B.n553 B.n315 10.6151
R1706 B.n554 B.n553 10.6151
R1707 B.n555 B.n554 10.6151
R1708 B.n555 B.n307 10.6151
R1709 B.n565 B.n307 10.6151
R1710 B.n566 B.n565 10.6151
R1711 B.n567 B.n566 10.6151
R1712 B.n567 B.n299 10.6151
R1713 B.n577 B.n299 10.6151
R1714 B.n578 B.n577 10.6151
R1715 B.n579 B.n578 10.6151
R1716 B.n579 B.n291 10.6151
R1717 B.n590 B.n291 10.6151
R1718 B.n591 B.n590 10.6151
R1719 B.n592 B.n591 10.6151
R1720 B.n592 B.n284 10.6151
R1721 B.n602 B.n284 10.6151
R1722 B.n603 B.n602 10.6151
R1723 B.n604 B.n603 10.6151
R1724 B.n604 B.n276 10.6151
R1725 B.n615 B.n276 10.6151
R1726 B.n616 B.n615 10.6151
R1727 B.n617 B.n616 10.6151
R1728 B.n617 B.n269 10.6151
R1729 B.n627 B.n269 10.6151
R1730 B.n628 B.n627 10.6151
R1731 B.n629 B.n628 10.6151
R1732 B.n629 B.n261 10.6151
R1733 B.n639 B.n261 10.6151
R1734 B.n640 B.n639 10.6151
R1735 B.n641 B.n640 10.6151
R1736 B.n641 B.n253 10.6151
R1737 B.n652 B.n253 10.6151
R1738 B.n653 B.n652 10.6151
R1739 B.n654 B.n653 10.6151
R1740 B.n654 B.n0 10.6151
R1741 B.n505 B.n347 10.6151
R1742 B.n500 B.n347 10.6151
R1743 B.n500 B.n499 10.6151
R1744 B.n499 B.n498 10.6151
R1745 B.n498 B.n495 10.6151
R1746 B.n495 B.n494 10.6151
R1747 B.n494 B.n491 10.6151
R1748 B.n491 B.n490 10.6151
R1749 B.n490 B.n487 10.6151
R1750 B.n487 B.n486 10.6151
R1751 B.n486 B.n483 10.6151
R1752 B.n483 B.n482 10.6151
R1753 B.n482 B.n479 10.6151
R1754 B.n479 B.n478 10.6151
R1755 B.n478 B.n475 10.6151
R1756 B.n475 B.n474 10.6151
R1757 B.n474 B.n471 10.6151
R1758 B.n471 B.n470 10.6151
R1759 B.n470 B.n467 10.6151
R1760 B.n467 B.n466 10.6151
R1761 B.n466 B.n463 10.6151
R1762 B.n463 B.n462 10.6151
R1763 B.n462 B.n459 10.6151
R1764 B.n459 B.n458 10.6151
R1765 B.n458 B.n455 10.6151
R1766 B.n453 B.n450 10.6151
R1767 B.n450 B.n449 10.6151
R1768 B.n449 B.n446 10.6151
R1769 B.n446 B.n445 10.6151
R1770 B.n445 B.n442 10.6151
R1771 B.n442 B.n441 10.6151
R1772 B.n441 B.n438 10.6151
R1773 B.n438 B.n437 10.6151
R1774 B.n434 B.n433 10.6151
R1775 B.n433 B.n430 10.6151
R1776 B.n430 B.n429 10.6151
R1777 B.n429 B.n426 10.6151
R1778 B.n426 B.n425 10.6151
R1779 B.n425 B.n422 10.6151
R1780 B.n422 B.n421 10.6151
R1781 B.n421 B.n418 10.6151
R1782 B.n418 B.n417 10.6151
R1783 B.n417 B.n414 10.6151
R1784 B.n414 B.n413 10.6151
R1785 B.n413 B.n410 10.6151
R1786 B.n410 B.n409 10.6151
R1787 B.n409 B.n406 10.6151
R1788 B.n406 B.n405 10.6151
R1789 B.n405 B.n402 10.6151
R1790 B.n402 B.n401 10.6151
R1791 B.n401 B.n398 10.6151
R1792 B.n398 B.n397 10.6151
R1793 B.n397 B.n394 10.6151
R1794 B.n394 B.n393 10.6151
R1795 B.n393 B.n390 10.6151
R1796 B.n390 B.n389 10.6151
R1797 B.n389 B.n386 10.6151
R1798 B.n386 B.n385 10.6151
R1799 B.n511 B.n343 10.6151
R1800 B.n512 B.n511 10.6151
R1801 B.n513 B.n512 10.6151
R1802 B.n513 B.n335 10.6151
R1803 B.n523 B.n335 10.6151
R1804 B.n524 B.n523 10.6151
R1805 B.n525 B.n524 10.6151
R1806 B.n525 B.n327 10.6151
R1807 B.n535 B.n327 10.6151
R1808 B.n536 B.n535 10.6151
R1809 B.n537 B.n536 10.6151
R1810 B.n537 B.n319 10.6151
R1811 B.n547 B.n319 10.6151
R1812 B.n548 B.n547 10.6151
R1813 B.n549 B.n548 10.6151
R1814 B.n549 B.n311 10.6151
R1815 B.n559 B.n311 10.6151
R1816 B.n560 B.n559 10.6151
R1817 B.n561 B.n560 10.6151
R1818 B.n561 B.n303 10.6151
R1819 B.n571 B.n303 10.6151
R1820 B.n572 B.n571 10.6151
R1821 B.n573 B.n572 10.6151
R1822 B.n573 B.n295 10.6151
R1823 B.n583 B.n295 10.6151
R1824 B.n584 B.n583 10.6151
R1825 B.n585 B.n584 10.6151
R1826 B.n585 B.n288 10.6151
R1827 B.n596 B.n288 10.6151
R1828 B.n597 B.n596 10.6151
R1829 B.n598 B.n597 10.6151
R1830 B.n598 B.n280 10.6151
R1831 B.n608 B.n280 10.6151
R1832 B.n609 B.n608 10.6151
R1833 B.n610 B.n609 10.6151
R1834 B.n610 B.n273 10.6151
R1835 B.n621 B.n273 10.6151
R1836 B.n622 B.n621 10.6151
R1837 B.n623 B.n622 10.6151
R1838 B.n623 B.n265 10.6151
R1839 B.n633 B.n265 10.6151
R1840 B.n634 B.n633 10.6151
R1841 B.n635 B.n634 10.6151
R1842 B.n635 B.n257 10.6151
R1843 B.n645 B.n257 10.6151
R1844 B.n646 B.n645 10.6151
R1845 B.n648 B.n646 10.6151
R1846 B.n648 B.n647 10.6151
R1847 B.n647 B.n249 10.6151
R1848 B.n659 B.n249 10.6151
R1849 B.n660 B.n659 10.6151
R1850 B.n661 B.n660 10.6151
R1851 B.n662 B.n661 10.6151
R1852 B.n663 B.n662 10.6151
R1853 B.n666 B.n663 10.6151
R1854 B.n667 B.n666 10.6151
R1855 B.n668 B.n667 10.6151
R1856 B.n669 B.n668 10.6151
R1857 B.n671 B.n669 10.6151
R1858 B.n672 B.n671 10.6151
R1859 B.n673 B.n672 10.6151
R1860 B.n674 B.n673 10.6151
R1861 B.n676 B.n674 10.6151
R1862 B.n677 B.n676 10.6151
R1863 B.n678 B.n677 10.6151
R1864 B.n679 B.n678 10.6151
R1865 B.n681 B.n679 10.6151
R1866 B.n682 B.n681 10.6151
R1867 B.n683 B.n682 10.6151
R1868 B.n684 B.n683 10.6151
R1869 B.n686 B.n684 10.6151
R1870 B.n687 B.n686 10.6151
R1871 B.n688 B.n687 10.6151
R1872 B.n689 B.n688 10.6151
R1873 B.n691 B.n689 10.6151
R1874 B.n692 B.n691 10.6151
R1875 B.n693 B.n692 10.6151
R1876 B.n694 B.n693 10.6151
R1877 B.n696 B.n694 10.6151
R1878 B.n697 B.n696 10.6151
R1879 B.n698 B.n697 10.6151
R1880 B.n699 B.n698 10.6151
R1881 B.n701 B.n699 10.6151
R1882 B.n702 B.n701 10.6151
R1883 B.n703 B.n702 10.6151
R1884 B.n704 B.n703 10.6151
R1885 B.n706 B.n704 10.6151
R1886 B.n707 B.n706 10.6151
R1887 B.n708 B.n707 10.6151
R1888 B.n709 B.n708 10.6151
R1889 B.n711 B.n709 10.6151
R1890 B.n712 B.n711 10.6151
R1891 B.n713 B.n712 10.6151
R1892 B.n714 B.n713 10.6151
R1893 B.n716 B.n714 10.6151
R1894 B.n717 B.n716 10.6151
R1895 B.n718 B.n717 10.6151
R1896 B.n719 B.n718 10.6151
R1897 B.n721 B.n719 10.6151
R1898 B.n722 B.n721 10.6151
R1899 B.n723 B.n722 10.6151
R1900 B.n724 B.n723 10.6151
R1901 B.n725 B.n724 10.6151
R1902 B.n829 B.n1 10.6151
R1903 B.n829 B.n828 10.6151
R1904 B.n828 B.n827 10.6151
R1905 B.n827 B.n10 10.6151
R1906 B.n821 B.n10 10.6151
R1907 B.n821 B.n820 10.6151
R1908 B.n820 B.n819 10.6151
R1909 B.n819 B.n18 10.6151
R1910 B.n813 B.n18 10.6151
R1911 B.n813 B.n812 10.6151
R1912 B.n812 B.n811 10.6151
R1913 B.n811 B.n25 10.6151
R1914 B.n805 B.n25 10.6151
R1915 B.n805 B.n804 10.6151
R1916 B.n804 B.n803 10.6151
R1917 B.n803 B.n31 10.6151
R1918 B.n797 B.n31 10.6151
R1919 B.n797 B.n796 10.6151
R1920 B.n796 B.n795 10.6151
R1921 B.n795 B.n39 10.6151
R1922 B.n789 B.n39 10.6151
R1923 B.n789 B.n788 10.6151
R1924 B.n788 B.n787 10.6151
R1925 B.n787 B.n45 10.6151
R1926 B.n781 B.n45 10.6151
R1927 B.n781 B.n780 10.6151
R1928 B.n780 B.n779 10.6151
R1929 B.n779 B.n53 10.6151
R1930 B.n773 B.n53 10.6151
R1931 B.n773 B.n772 10.6151
R1932 B.n772 B.n771 10.6151
R1933 B.n771 B.n60 10.6151
R1934 B.n765 B.n60 10.6151
R1935 B.n765 B.n764 10.6151
R1936 B.n764 B.n763 10.6151
R1937 B.n763 B.n67 10.6151
R1938 B.n757 B.n67 10.6151
R1939 B.n757 B.n756 10.6151
R1940 B.n756 B.n755 10.6151
R1941 B.n755 B.n74 10.6151
R1942 B.n749 B.n74 10.6151
R1943 B.n749 B.n748 10.6151
R1944 B.n748 B.n747 10.6151
R1945 B.n747 B.n81 10.6151
R1946 B.n741 B.n81 10.6151
R1947 B.n741 B.n740 10.6151
R1948 B.n740 B.n739 10.6151
R1949 B.n739 B.n88 10.6151
R1950 B.n733 B.n88 10.6151
R1951 B.n733 B.n732 10.6151
R1952 B.n731 B.n95 10.6151
R1953 B.n134 B.n95 10.6151
R1954 B.n135 B.n134 10.6151
R1955 B.n138 B.n135 10.6151
R1956 B.n139 B.n138 10.6151
R1957 B.n142 B.n139 10.6151
R1958 B.n143 B.n142 10.6151
R1959 B.n146 B.n143 10.6151
R1960 B.n147 B.n146 10.6151
R1961 B.n150 B.n147 10.6151
R1962 B.n151 B.n150 10.6151
R1963 B.n154 B.n151 10.6151
R1964 B.n155 B.n154 10.6151
R1965 B.n158 B.n155 10.6151
R1966 B.n159 B.n158 10.6151
R1967 B.n162 B.n159 10.6151
R1968 B.n163 B.n162 10.6151
R1969 B.n166 B.n163 10.6151
R1970 B.n167 B.n166 10.6151
R1971 B.n170 B.n167 10.6151
R1972 B.n171 B.n170 10.6151
R1973 B.n174 B.n171 10.6151
R1974 B.n175 B.n174 10.6151
R1975 B.n178 B.n175 10.6151
R1976 B.n179 B.n178 10.6151
R1977 B.n183 B.n182 10.6151
R1978 B.n186 B.n183 10.6151
R1979 B.n187 B.n186 10.6151
R1980 B.n190 B.n187 10.6151
R1981 B.n191 B.n190 10.6151
R1982 B.n194 B.n191 10.6151
R1983 B.n195 B.n194 10.6151
R1984 B.n198 B.n195 10.6151
R1985 B.n203 B.n200 10.6151
R1986 B.n204 B.n203 10.6151
R1987 B.n207 B.n204 10.6151
R1988 B.n208 B.n207 10.6151
R1989 B.n211 B.n208 10.6151
R1990 B.n212 B.n211 10.6151
R1991 B.n215 B.n212 10.6151
R1992 B.n216 B.n215 10.6151
R1993 B.n219 B.n216 10.6151
R1994 B.n220 B.n219 10.6151
R1995 B.n223 B.n220 10.6151
R1996 B.n224 B.n223 10.6151
R1997 B.n227 B.n224 10.6151
R1998 B.n228 B.n227 10.6151
R1999 B.n231 B.n228 10.6151
R2000 B.n232 B.n231 10.6151
R2001 B.n235 B.n232 10.6151
R2002 B.n236 B.n235 10.6151
R2003 B.n239 B.n236 10.6151
R2004 B.n240 B.n239 10.6151
R2005 B.n243 B.n240 10.6151
R2006 B.n244 B.n243 10.6151
R2007 B.n247 B.n244 10.6151
R2008 B.n248 B.n247 10.6151
R2009 B.n726 B.n248 10.6151
R2010 B.n837 B.n0 8.11757
R2011 B.n837 B.n1 8.11757
R2012 B.n454 B.n453 6.5566
R2013 B.n437 B.n383 6.5566
R2014 B.n182 B.n132 6.5566
R2015 B.n199 B.n198 6.5566
R2016 B.n455 B.n454 4.05904
R2017 B.n434 B.n383 4.05904
R2018 B.n179 B.n132 4.05904
R2019 B.n200 B.n199 4.05904
R2020 B.n587 B.t1 3.69023
R2021 B.n47 B.t0 3.69023
R2022 VP.n19 VP.n16 161.3
R2023 VP.n21 VP.n20 161.3
R2024 VP.n22 VP.n15 161.3
R2025 VP.n24 VP.n23 161.3
R2026 VP.n25 VP.n14 161.3
R2027 VP.n27 VP.n26 161.3
R2028 VP.n29 VP.n28 161.3
R2029 VP.n30 VP.n12 161.3
R2030 VP.n32 VP.n31 161.3
R2031 VP.n33 VP.n11 161.3
R2032 VP.n35 VP.n34 161.3
R2033 VP.n36 VP.n10 161.3
R2034 VP.n68 VP.n0 161.3
R2035 VP.n67 VP.n66 161.3
R2036 VP.n65 VP.n1 161.3
R2037 VP.n64 VP.n63 161.3
R2038 VP.n62 VP.n2 161.3
R2039 VP.n61 VP.n60 161.3
R2040 VP.n59 VP.n58 161.3
R2041 VP.n57 VP.n4 161.3
R2042 VP.n56 VP.n55 161.3
R2043 VP.n54 VP.n5 161.3
R2044 VP.n53 VP.n52 161.3
R2045 VP.n51 VP.n6 161.3
R2046 VP.n49 VP.n48 161.3
R2047 VP.n47 VP.n7 161.3
R2048 VP.n46 VP.n45 161.3
R2049 VP.n44 VP.n8 161.3
R2050 VP.n43 VP.n42 161.3
R2051 VP.n41 VP.n9 161.3
R2052 VP.n40 VP.n39 100.725
R2053 VP.n70 VP.n69 100.725
R2054 VP.n38 VP.n37 100.725
R2055 VP.n17 VP.t6 94.3223
R2056 VP.n18 VP.n17 60.9555
R2057 VP.n39 VP.t2 60.7069
R2058 VP.n50 VP.t5 60.7069
R2059 VP.n3 VP.t4 60.7069
R2060 VP.n69 VP.t1 60.7069
R2061 VP.n37 VP.t0 60.7069
R2062 VP.n13 VP.t3 60.7069
R2063 VP.n18 VP.t7 60.7069
R2064 VP.n45 VP.n44 56.5193
R2065 VP.n56 VP.n5 56.5193
R2066 VP.n63 VP.n1 56.5193
R2067 VP.n31 VP.n11 56.5193
R2068 VP.n24 VP.n15 56.5193
R2069 VP.n40 VP.n38 47.0602
R2070 VP.n43 VP.n9 24.4675
R2071 VP.n44 VP.n43 24.4675
R2072 VP.n45 VP.n7 24.4675
R2073 VP.n49 VP.n7 24.4675
R2074 VP.n52 VP.n51 24.4675
R2075 VP.n52 VP.n5 24.4675
R2076 VP.n57 VP.n56 24.4675
R2077 VP.n58 VP.n57 24.4675
R2078 VP.n62 VP.n61 24.4675
R2079 VP.n63 VP.n62 24.4675
R2080 VP.n67 VP.n1 24.4675
R2081 VP.n68 VP.n67 24.4675
R2082 VP.n35 VP.n11 24.4675
R2083 VP.n36 VP.n35 24.4675
R2084 VP.n25 VP.n24 24.4675
R2085 VP.n26 VP.n25 24.4675
R2086 VP.n30 VP.n29 24.4675
R2087 VP.n31 VP.n30 24.4675
R2088 VP.n20 VP.n19 24.4675
R2089 VP.n20 VP.n15 24.4675
R2090 VP.n50 VP.n49 12.968
R2091 VP.n61 VP.n3 12.968
R2092 VP.n29 VP.n13 12.968
R2093 VP.n51 VP.n50 11.5
R2094 VP.n58 VP.n3 11.5
R2095 VP.n26 VP.n13 11.5
R2096 VP.n19 VP.n18 11.5
R2097 VP.n39 VP.n9 10.032
R2098 VP.n69 VP.n68 10.032
R2099 VP.n37 VP.n36 10.032
R2100 VP.n17 VP.n16 6.848
R2101 VP.n38 VP.n10 0.278367
R2102 VP.n41 VP.n40 0.278367
R2103 VP.n70 VP.n0 0.278367
R2104 VP.n21 VP.n16 0.189894
R2105 VP.n22 VP.n21 0.189894
R2106 VP.n23 VP.n22 0.189894
R2107 VP.n23 VP.n14 0.189894
R2108 VP.n27 VP.n14 0.189894
R2109 VP.n28 VP.n27 0.189894
R2110 VP.n28 VP.n12 0.189894
R2111 VP.n32 VP.n12 0.189894
R2112 VP.n33 VP.n32 0.189894
R2113 VP.n34 VP.n33 0.189894
R2114 VP.n34 VP.n10 0.189894
R2115 VP.n42 VP.n41 0.189894
R2116 VP.n42 VP.n8 0.189894
R2117 VP.n46 VP.n8 0.189894
R2118 VP.n47 VP.n46 0.189894
R2119 VP.n48 VP.n47 0.189894
R2120 VP.n48 VP.n6 0.189894
R2121 VP.n53 VP.n6 0.189894
R2122 VP.n54 VP.n53 0.189894
R2123 VP.n55 VP.n54 0.189894
R2124 VP.n55 VP.n4 0.189894
R2125 VP.n59 VP.n4 0.189894
R2126 VP.n60 VP.n59 0.189894
R2127 VP.n60 VP.n2 0.189894
R2128 VP.n64 VP.n2 0.189894
R2129 VP.n65 VP.n64 0.189894
R2130 VP.n66 VP.n65 0.189894
R2131 VP.n66 VP.n0 0.189894
R2132 VP VP.n70 0.153454
R2133 VDD1 VDD1.n0 66.0549
R2134 VDD1.n3 VDD1.n2 65.9412
R2135 VDD1.n3 VDD1.n1 65.9412
R2136 VDD1.n5 VDD1.n4 64.7164
R2137 VDD1.n5 VDD1.n3 41.5526
R2138 VDD1.n4 VDD1.t4 2.97794
R2139 VDD1.n4 VDD1.t7 2.97794
R2140 VDD1.n0 VDD1.t1 2.97794
R2141 VDD1.n0 VDD1.t0 2.97794
R2142 VDD1.n2 VDD1.t3 2.97794
R2143 VDD1.n2 VDD1.t6 2.97794
R2144 VDD1.n1 VDD1.t5 2.97794
R2145 VDD1.n1 VDD1.t2 2.97794
R2146 VDD1 VDD1.n5 1.22248
C0 VP VTAIL 5.86057f
C1 VDD2 VTAIL 6.35609f
C2 VP VDD2 0.524035f
C3 VDD1 VN 0.151908f
C4 VTAIL VN 5.84647f
C5 VDD1 VTAIL 6.3014f
C6 VP VN 6.71891f
C7 VDD1 VP 5.40058f
C8 VDD2 VN 5.02987f
C9 VDD1 VDD2 1.79895f
C10 VDD2 B 4.968823f
C11 VDD1 B 5.41399f
C12 VTAIL B 6.940331f
C13 VN B 15.04896f
C14 VP B 13.684029f
C15 VDD1.t1 B 0.129783f
C16 VDD1.t0 B 0.129783f
C17 VDD1.n0 B 1.10526f
C18 VDD1.t5 B 0.129783f
C19 VDD1.t2 B 0.129783f
C20 VDD1.n1 B 1.10421f
C21 VDD1.t3 B 0.129783f
C22 VDD1.t6 B 0.129783f
C23 VDD1.n2 B 1.10421f
C24 VDD1.n3 B 2.98642f
C25 VDD1.t4 B 0.129783f
C26 VDD1.t7 B 0.129783f
C27 VDD1.n4 B 1.09465f
C28 VDD1.n5 B 2.55055f
C29 VP.n0 B 0.03259f
C30 VP.t1 B 1.15523f
C31 VP.n1 B 0.038152f
C32 VP.n2 B 0.024719f
C33 VP.t4 B 1.15523f
C34 VP.n3 B 0.428142f
C35 VP.n4 B 0.024719f
C36 VP.n5 B 0.036086f
C37 VP.n6 B 0.024719f
C38 VP.t5 B 1.15523f
C39 VP.n7 B 0.046071f
C40 VP.n8 B 0.024719f
C41 VP.n9 B 0.03265f
C42 VP.n10 B 0.03259f
C43 VP.t0 B 1.15523f
C44 VP.n11 B 0.038152f
C45 VP.n12 B 0.024719f
C46 VP.t3 B 1.15523f
C47 VP.n13 B 0.428142f
C48 VP.n14 B 0.024719f
C49 VP.n15 B 0.036086f
C50 VP.n16 B 0.239947f
C51 VP.t7 B 1.15523f
C52 VP.t6 B 1.3631f
C53 VP.n17 B 0.480154f
C54 VP.n18 B 0.499343f
C55 VP.n19 B 0.034015f
C56 VP.n20 B 0.046071f
C57 VP.n21 B 0.024719f
C58 VP.n22 B 0.024719f
C59 VP.n23 B 0.024719f
C60 VP.n24 B 0.036086f
C61 VP.n25 B 0.046071f
C62 VP.n26 B 0.034015f
C63 VP.n27 B 0.024719f
C64 VP.n28 B 0.024719f
C65 VP.n29 B 0.035379f
C66 VP.n30 B 0.046071f
C67 VP.n31 B 0.034019f
C68 VP.n32 B 0.024719f
C69 VP.n33 B 0.024719f
C70 VP.n34 B 0.024719f
C71 VP.n35 B 0.046071f
C72 VP.n36 B 0.03265f
C73 VP.n37 B 0.5125f
C74 VP.n38 B 1.2572f
C75 VP.t2 B 1.15523f
C76 VP.n39 B 0.5125f
C77 VP.n40 B 1.27609f
C78 VP.n41 B 0.03259f
C79 VP.n42 B 0.024719f
C80 VP.n43 B 0.046071f
C81 VP.n44 B 0.038152f
C82 VP.n45 B 0.034019f
C83 VP.n46 B 0.024719f
C84 VP.n47 B 0.024719f
C85 VP.n48 B 0.024719f
C86 VP.n49 B 0.035379f
C87 VP.n50 B 0.428142f
C88 VP.n51 B 0.034015f
C89 VP.n52 B 0.046071f
C90 VP.n53 B 0.024719f
C91 VP.n54 B 0.024719f
C92 VP.n55 B 0.024719f
C93 VP.n56 B 0.036086f
C94 VP.n57 B 0.046071f
C95 VP.n58 B 0.034015f
C96 VP.n59 B 0.024719f
C97 VP.n60 B 0.024719f
C98 VP.n61 B 0.035379f
C99 VP.n62 B 0.046071f
C100 VP.n63 B 0.034019f
C101 VP.n64 B 0.024719f
C102 VP.n65 B 0.024719f
C103 VP.n66 B 0.024719f
C104 VP.n67 B 0.046071f
C105 VP.n68 B 0.03265f
C106 VP.n69 B 0.5125f
C107 VP.n70 B 0.040496f
C108 VDD2.t6 B 0.127448f
C109 VDD2.t4 B 0.127448f
C110 VDD2.n0 B 1.08436f
C111 VDD2.t2 B 0.127448f
C112 VDD2.t0 B 0.127448f
C113 VDD2.n1 B 1.08436f
C114 VDD2.n2 B 2.88205f
C115 VDD2.t5 B 0.127448f
C116 VDD2.t7 B 0.127448f
C117 VDD2.n3 B 1.07497f
C118 VDD2.n4 B 2.47484f
C119 VDD2.t1 B 0.127448f
C120 VDD2.t3 B 0.127448f
C121 VDD2.n5 B 1.08432f
C122 VTAIL.t12 B 0.119809f
C123 VTAIL.t15 B 0.119809f
C124 VTAIL.n0 B 0.946943f
C125 VTAIL.n1 B 0.412446f
C126 VTAIL.n2 B 0.031584f
C127 VTAIL.n3 B 0.022799f
C128 VTAIL.n4 B 0.012251f
C129 VTAIL.n5 B 0.028957f
C130 VTAIL.n6 B 0.012972f
C131 VTAIL.n7 B 0.022799f
C132 VTAIL.n8 B 0.012251f
C133 VTAIL.n9 B 0.028957f
C134 VTAIL.n10 B 0.012972f
C135 VTAIL.n11 B 0.610638f
C136 VTAIL.n12 B 0.012251f
C137 VTAIL.t10 B 0.047166f
C138 VTAIL.n13 B 0.101116f
C139 VTAIL.n14 B 0.017106f
C140 VTAIL.n15 B 0.021718f
C141 VTAIL.n16 B 0.028957f
C142 VTAIL.n17 B 0.012972f
C143 VTAIL.n18 B 0.012251f
C144 VTAIL.n19 B 0.022799f
C145 VTAIL.n20 B 0.022799f
C146 VTAIL.n21 B 0.012251f
C147 VTAIL.n22 B 0.012972f
C148 VTAIL.n23 B 0.028957f
C149 VTAIL.n24 B 0.028957f
C150 VTAIL.n25 B 0.012972f
C151 VTAIL.n26 B 0.012251f
C152 VTAIL.n27 B 0.022799f
C153 VTAIL.n28 B 0.022799f
C154 VTAIL.n29 B 0.012251f
C155 VTAIL.n30 B 0.012972f
C156 VTAIL.n31 B 0.028957f
C157 VTAIL.n32 B 0.061871f
C158 VTAIL.n33 B 0.012972f
C159 VTAIL.n34 B 0.012251f
C160 VTAIL.n35 B 0.050518f
C161 VTAIL.n36 B 0.034467f
C162 VTAIL.n37 B 0.240848f
C163 VTAIL.n38 B 0.031584f
C164 VTAIL.n39 B 0.022799f
C165 VTAIL.n40 B 0.012251f
C166 VTAIL.n41 B 0.028957f
C167 VTAIL.n42 B 0.012972f
C168 VTAIL.n43 B 0.022799f
C169 VTAIL.n44 B 0.012251f
C170 VTAIL.n45 B 0.028957f
C171 VTAIL.n46 B 0.012972f
C172 VTAIL.n47 B 0.610638f
C173 VTAIL.n48 B 0.012251f
C174 VTAIL.t4 B 0.047166f
C175 VTAIL.n49 B 0.101116f
C176 VTAIL.n50 B 0.017106f
C177 VTAIL.n51 B 0.021718f
C178 VTAIL.n52 B 0.028957f
C179 VTAIL.n53 B 0.012972f
C180 VTAIL.n54 B 0.012251f
C181 VTAIL.n55 B 0.022799f
C182 VTAIL.n56 B 0.022799f
C183 VTAIL.n57 B 0.012251f
C184 VTAIL.n58 B 0.012972f
C185 VTAIL.n59 B 0.028957f
C186 VTAIL.n60 B 0.028957f
C187 VTAIL.n61 B 0.012972f
C188 VTAIL.n62 B 0.012251f
C189 VTAIL.n63 B 0.022799f
C190 VTAIL.n64 B 0.022799f
C191 VTAIL.n65 B 0.012251f
C192 VTAIL.n66 B 0.012972f
C193 VTAIL.n67 B 0.028957f
C194 VTAIL.n68 B 0.061871f
C195 VTAIL.n69 B 0.012972f
C196 VTAIL.n70 B 0.012251f
C197 VTAIL.n71 B 0.050518f
C198 VTAIL.n72 B 0.034467f
C199 VTAIL.n73 B 0.240848f
C200 VTAIL.t1 B 0.119809f
C201 VTAIL.t7 B 0.119809f
C202 VTAIL.n74 B 0.946943f
C203 VTAIL.n75 B 0.596262f
C204 VTAIL.n76 B 0.031584f
C205 VTAIL.n77 B 0.022799f
C206 VTAIL.n78 B 0.012251f
C207 VTAIL.n79 B 0.028957f
C208 VTAIL.n80 B 0.012972f
C209 VTAIL.n81 B 0.022799f
C210 VTAIL.n82 B 0.012251f
C211 VTAIL.n83 B 0.028957f
C212 VTAIL.n84 B 0.012972f
C213 VTAIL.n85 B 0.610638f
C214 VTAIL.n86 B 0.012251f
C215 VTAIL.t6 B 0.047166f
C216 VTAIL.n87 B 0.101116f
C217 VTAIL.n88 B 0.017106f
C218 VTAIL.n89 B 0.021718f
C219 VTAIL.n90 B 0.028957f
C220 VTAIL.n91 B 0.012972f
C221 VTAIL.n92 B 0.012251f
C222 VTAIL.n93 B 0.022799f
C223 VTAIL.n94 B 0.022799f
C224 VTAIL.n95 B 0.012251f
C225 VTAIL.n96 B 0.012972f
C226 VTAIL.n97 B 0.028957f
C227 VTAIL.n98 B 0.028957f
C228 VTAIL.n99 B 0.012972f
C229 VTAIL.n100 B 0.012251f
C230 VTAIL.n101 B 0.022799f
C231 VTAIL.n102 B 0.022799f
C232 VTAIL.n103 B 0.012251f
C233 VTAIL.n104 B 0.012972f
C234 VTAIL.n105 B 0.028957f
C235 VTAIL.n106 B 0.061871f
C236 VTAIL.n107 B 0.012972f
C237 VTAIL.n108 B 0.012251f
C238 VTAIL.n109 B 0.050518f
C239 VTAIL.n110 B 0.034467f
C240 VTAIL.n111 B 1.12527f
C241 VTAIL.n112 B 0.031584f
C242 VTAIL.n113 B 0.022799f
C243 VTAIL.n114 B 0.012251f
C244 VTAIL.n115 B 0.028957f
C245 VTAIL.n116 B 0.012972f
C246 VTAIL.n117 B 0.022799f
C247 VTAIL.n118 B 0.012251f
C248 VTAIL.n119 B 0.028957f
C249 VTAIL.n120 B 0.012972f
C250 VTAIL.n121 B 0.610638f
C251 VTAIL.n122 B 0.012251f
C252 VTAIL.t14 B 0.047166f
C253 VTAIL.n123 B 0.101116f
C254 VTAIL.n124 B 0.017106f
C255 VTAIL.n125 B 0.021718f
C256 VTAIL.n126 B 0.028957f
C257 VTAIL.n127 B 0.012972f
C258 VTAIL.n128 B 0.012251f
C259 VTAIL.n129 B 0.022799f
C260 VTAIL.n130 B 0.022799f
C261 VTAIL.n131 B 0.012251f
C262 VTAIL.n132 B 0.012972f
C263 VTAIL.n133 B 0.028957f
C264 VTAIL.n134 B 0.028957f
C265 VTAIL.n135 B 0.012972f
C266 VTAIL.n136 B 0.012251f
C267 VTAIL.n137 B 0.022799f
C268 VTAIL.n138 B 0.022799f
C269 VTAIL.n139 B 0.012251f
C270 VTAIL.n140 B 0.012972f
C271 VTAIL.n141 B 0.028957f
C272 VTAIL.n142 B 0.061871f
C273 VTAIL.n143 B 0.012972f
C274 VTAIL.n144 B 0.012251f
C275 VTAIL.n145 B 0.050518f
C276 VTAIL.n146 B 0.034467f
C277 VTAIL.n147 B 1.12527f
C278 VTAIL.t11 B 0.119809f
C279 VTAIL.t13 B 0.119809f
C280 VTAIL.n148 B 0.94695f
C281 VTAIL.n149 B 0.596255f
C282 VTAIL.n150 B 0.031584f
C283 VTAIL.n151 B 0.022799f
C284 VTAIL.n152 B 0.012251f
C285 VTAIL.n153 B 0.028957f
C286 VTAIL.n154 B 0.012972f
C287 VTAIL.n155 B 0.022799f
C288 VTAIL.n156 B 0.012251f
C289 VTAIL.n157 B 0.028957f
C290 VTAIL.n158 B 0.012972f
C291 VTAIL.n159 B 0.610638f
C292 VTAIL.n160 B 0.012251f
C293 VTAIL.t9 B 0.047166f
C294 VTAIL.n161 B 0.101116f
C295 VTAIL.n162 B 0.017106f
C296 VTAIL.n163 B 0.021718f
C297 VTAIL.n164 B 0.028957f
C298 VTAIL.n165 B 0.012972f
C299 VTAIL.n166 B 0.012251f
C300 VTAIL.n167 B 0.022799f
C301 VTAIL.n168 B 0.022799f
C302 VTAIL.n169 B 0.012251f
C303 VTAIL.n170 B 0.012972f
C304 VTAIL.n171 B 0.028957f
C305 VTAIL.n172 B 0.028957f
C306 VTAIL.n173 B 0.012972f
C307 VTAIL.n174 B 0.012251f
C308 VTAIL.n175 B 0.022799f
C309 VTAIL.n176 B 0.022799f
C310 VTAIL.n177 B 0.012251f
C311 VTAIL.n178 B 0.012972f
C312 VTAIL.n179 B 0.028957f
C313 VTAIL.n180 B 0.061871f
C314 VTAIL.n181 B 0.012972f
C315 VTAIL.n182 B 0.012251f
C316 VTAIL.n183 B 0.050518f
C317 VTAIL.n184 B 0.034467f
C318 VTAIL.n185 B 0.240848f
C319 VTAIL.n186 B 0.031584f
C320 VTAIL.n187 B 0.022799f
C321 VTAIL.n188 B 0.012251f
C322 VTAIL.n189 B 0.028957f
C323 VTAIL.n190 B 0.012972f
C324 VTAIL.n191 B 0.022799f
C325 VTAIL.n192 B 0.012251f
C326 VTAIL.n193 B 0.028957f
C327 VTAIL.n194 B 0.012972f
C328 VTAIL.n195 B 0.610638f
C329 VTAIL.n196 B 0.012251f
C330 VTAIL.t3 B 0.047166f
C331 VTAIL.n197 B 0.101116f
C332 VTAIL.n198 B 0.017106f
C333 VTAIL.n199 B 0.021718f
C334 VTAIL.n200 B 0.028957f
C335 VTAIL.n201 B 0.012972f
C336 VTAIL.n202 B 0.012251f
C337 VTAIL.n203 B 0.022799f
C338 VTAIL.n204 B 0.022799f
C339 VTAIL.n205 B 0.012251f
C340 VTAIL.n206 B 0.012972f
C341 VTAIL.n207 B 0.028957f
C342 VTAIL.n208 B 0.028957f
C343 VTAIL.n209 B 0.012972f
C344 VTAIL.n210 B 0.012251f
C345 VTAIL.n211 B 0.022799f
C346 VTAIL.n212 B 0.022799f
C347 VTAIL.n213 B 0.012251f
C348 VTAIL.n214 B 0.012972f
C349 VTAIL.n215 B 0.028957f
C350 VTAIL.n216 B 0.061871f
C351 VTAIL.n217 B 0.012972f
C352 VTAIL.n218 B 0.012251f
C353 VTAIL.n219 B 0.050518f
C354 VTAIL.n220 B 0.034467f
C355 VTAIL.n221 B 0.240848f
C356 VTAIL.t5 B 0.119809f
C357 VTAIL.t0 B 0.119809f
C358 VTAIL.n222 B 0.94695f
C359 VTAIL.n223 B 0.596255f
C360 VTAIL.n224 B 0.031584f
C361 VTAIL.n225 B 0.022799f
C362 VTAIL.n226 B 0.012251f
C363 VTAIL.n227 B 0.028957f
C364 VTAIL.n228 B 0.012972f
C365 VTAIL.n229 B 0.022799f
C366 VTAIL.n230 B 0.012251f
C367 VTAIL.n231 B 0.028957f
C368 VTAIL.n232 B 0.012972f
C369 VTAIL.n233 B 0.610638f
C370 VTAIL.n234 B 0.012251f
C371 VTAIL.t2 B 0.047166f
C372 VTAIL.n235 B 0.101116f
C373 VTAIL.n236 B 0.017106f
C374 VTAIL.n237 B 0.021718f
C375 VTAIL.n238 B 0.028957f
C376 VTAIL.n239 B 0.012972f
C377 VTAIL.n240 B 0.012251f
C378 VTAIL.n241 B 0.022799f
C379 VTAIL.n242 B 0.022799f
C380 VTAIL.n243 B 0.012251f
C381 VTAIL.n244 B 0.012972f
C382 VTAIL.n245 B 0.028957f
C383 VTAIL.n246 B 0.028957f
C384 VTAIL.n247 B 0.012972f
C385 VTAIL.n248 B 0.012251f
C386 VTAIL.n249 B 0.022799f
C387 VTAIL.n250 B 0.022799f
C388 VTAIL.n251 B 0.012251f
C389 VTAIL.n252 B 0.012972f
C390 VTAIL.n253 B 0.028957f
C391 VTAIL.n254 B 0.061871f
C392 VTAIL.n255 B 0.012972f
C393 VTAIL.n256 B 0.012251f
C394 VTAIL.n257 B 0.050518f
C395 VTAIL.n258 B 0.034467f
C396 VTAIL.n259 B 1.12527f
C397 VTAIL.n260 B 0.031584f
C398 VTAIL.n261 B 0.022799f
C399 VTAIL.n262 B 0.012251f
C400 VTAIL.n263 B 0.028957f
C401 VTAIL.n264 B 0.012972f
C402 VTAIL.n265 B 0.022799f
C403 VTAIL.n266 B 0.012251f
C404 VTAIL.n267 B 0.028957f
C405 VTAIL.n268 B 0.012972f
C406 VTAIL.n269 B 0.610638f
C407 VTAIL.n270 B 0.012251f
C408 VTAIL.t8 B 0.047166f
C409 VTAIL.n271 B 0.101116f
C410 VTAIL.n272 B 0.017106f
C411 VTAIL.n273 B 0.021718f
C412 VTAIL.n274 B 0.028957f
C413 VTAIL.n275 B 0.012972f
C414 VTAIL.n276 B 0.012251f
C415 VTAIL.n277 B 0.022799f
C416 VTAIL.n278 B 0.022799f
C417 VTAIL.n279 B 0.012251f
C418 VTAIL.n280 B 0.012972f
C419 VTAIL.n281 B 0.028957f
C420 VTAIL.n282 B 0.028957f
C421 VTAIL.n283 B 0.012972f
C422 VTAIL.n284 B 0.012251f
C423 VTAIL.n285 B 0.022799f
C424 VTAIL.n286 B 0.022799f
C425 VTAIL.n287 B 0.012251f
C426 VTAIL.n288 B 0.012972f
C427 VTAIL.n289 B 0.028957f
C428 VTAIL.n290 B 0.061871f
C429 VTAIL.n291 B 0.012972f
C430 VTAIL.n292 B 0.012251f
C431 VTAIL.n293 B 0.050518f
C432 VTAIL.n294 B 0.034467f
C433 VTAIL.n295 B 1.12099f
C434 VN.n0 B 0.031624f
C435 VN.t7 B 1.12098f
C436 VN.n1 B 0.037021f
C437 VN.n2 B 0.023986f
C438 VN.t5 B 1.12098f
C439 VN.n3 B 0.415447f
C440 VN.n4 B 0.023986f
C441 VN.n5 B 0.035016f
C442 VN.n6 B 0.232833f
C443 VN.t3 B 1.12098f
C444 VN.t1 B 1.32269f
C445 VN.n7 B 0.465917f
C446 VN.n8 B 0.484537f
C447 VN.n9 B 0.033006f
C448 VN.n10 B 0.044705f
C449 VN.n11 B 0.023986f
C450 VN.n12 B 0.023986f
C451 VN.n13 B 0.023986f
C452 VN.n14 B 0.035016f
C453 VN.n15 B 0.044705f
C454 VN.n16 B 0.033006f
C455 VN.n17 B 0.023986f
C456 VN.n18 B 0.023986f
C457 VN.n19 B 0.03433f
C458 VN.n20 B 0.044705f
C459 VN.n21 B 0.033011f
C460 VN.n22 B 0.023986f
C461 VN.n23 B 0.023986f
C462 VN.n24 B 0.023986f
C463 VN.n25 B 0.044705f
C464 VN.n26 B 0.031682f
C465 VN.n27 B 0.497304f
C466 VN.n28 B 0.039295f
C467 VN.n29 B 0.031624f
C468 VN.t2 B 1.12098f
C469 VN.n30 B 0.037021f
C470 VN.n31 B 0.023986f
C471 VN.t0 B 1.12098f
C472 VN.n32 B 0.415447f
C473 VN.n33 B 0.023986f
C474 VN.n34 B 0.035016f
C475 VN.n35 B 0.232833f
C476 VN.t6 B 1.12098f
C477 VN.t4 B 1.32269f
C478 VN.n36 B 0.465917f
C479 VN.n37 B 0.484537f
C480 VN.n38 B 0.033006f
C481 VN.n39 B 0.044705f
C482 VN.n40 B 0.023986f
C483 VN.n41 B 0.023986f
C484 VN.n42 B 0.023986f
C485 VN.n43 B 0.035016f
C486 VN.n44 B 0.044705f
C487 VN.n45 B 0.033006f
C488 VN.n46 B 0.023986f
C489 VN.n47 B 0.023986f
C490 VN.n48 B 0.03433f
C491 VN.n49 B 0.044705f
C492 VN.n50 B 0.033011f
C493 VN.n51 B 0.023986f
C494 VN.n52 B 0.023986f
C495 VN.n53 B 0.023986f
C496 VN.n54 B 0.044705f
C497 VN.n55 B 0.031682f
C498 VN.n56 B 0.497304f
C499 VN.n57 B 1.23294f
.ends

