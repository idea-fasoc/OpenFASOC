* NGSPICE file created from diff_pair_sample_1512.ext - technology: sky130A

.subckt diff_pair_sample_1512 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=2.0553 pd=11.32 as=0 ps=0 w=5.27 l=0.37
X1 VDD1.t9 VP.t0 VTAIL.t15 B.t8 sky130_fd_pr__nfet_01v8 ad=0.86955 pd=5.6 as=2.0553 ps=11.32 w=5.27 l=0.37
X2 VDD1.t8 VP.t1 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=0.37
X3 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=2.0553 pd=11.32 as=0 ps=0 w=5.27 l=0.37
X4 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=2.0553 pd=11.32 as=0 ps=0 w=5.27 l=0.37
X5 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.0553 pd=11.32 as=0 ps=0 w=5.27 l=0.37
X6 VTAIL.t11 VP.t2 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=0.37
X7 VDD2.t9 VN.t0 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=0.37
X8 VDD1.t6 VP.t3 VTAIL.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=0.37
X9 VTAIL.t1 VN.t1 VDD2.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=0.37
X10 VTAIL.t13 VP.t4 VDD1.t5 B.t9 sky130_fd_pr__nfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=0.37
X11 VDD1.t4 VP.t5 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=2.0553 pd=11.32 as=0.86955 ps=5.6 w=5.27 l=0.37
X12 VDD2.t7 VN.t2 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=0.37
X13 VDD2.t6 VN.t3 VTAIL.t17 B.t8 sky130_fd_pr__nfet_01v8 ad=0.86955 pd=5.6 as=2.0553 ps=11.32 w=5.27 l=0.37
X14 VDD1.t3 VP.t6 VTAIL.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=0.86955 pd=5.6 as=2.0553 ps=11.32 w=5.27 l=0.37
X15 VTAIL.t18 VN.t4 VDD2.t5 B.t9 sky130_fd_pr__nfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=0.37
X16 VDD1.t2 VP.t7 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.0553 pd=11.32 as=0.86955 ps=5.6 w=5.27 l=0.37
X17 VDD2.t4 VN.t5 VTAIL.t19 B.t7 sky130_fd_pr__nfet_01v8 ad=2.0553 pd=11.32 as=0.86955 ps=5.6 w=5.27 l=0.37
X18 VDD2.t3 VN.t6 VTAIL.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=0.86955 pd=5.6 as=2.0553 ps=11.32 w=5.27 l=0.37
X19 VDD2.t2 VN.t7 VTAIL.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=2.0553 pd=11.32 as=0.86955 ps=5.6 w=5.27 l=0.37
X20 VTAIL.t6 VN.t8 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=0.37
X21 VTAIL.t2 VN.t9 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=0.37
X22 VTAIL.t9 VP.t8 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=0.37
X23 VTAIL.t16 VP.t9 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=0.37
R0 B.n441 B.n440 585
R1 B.n442 B.n441 585
R2 B.n175 B.n68 585
R3 B.n174 B.n173 585
R4 B.n172 B.n171 585
R5 B.n170 B.n169 585
R6 B.n168 B.n167 585
R7 B.n166 B.n165 585
R8 B.n164 B.n163 585
R9 B.n162 B.n161 585
R10 B.n160 B.n159 585
R11 B.n158 B.n157 585
R12 B.n156 B.n155 585
R13 B.n154 B.n153 585
R14 B.n152 B.n151 585
R15 B.n150 B.n149 585
R16 B.n148 B.n147 585
R17 B.n146 B.n145 585
R18 B.n144 B.n143 585
R19 B.n142 B.n141 585
R20 B.n140 B.n139 585
R21 B.n138 B.n137 585
R22 B.n136 B.n135 585
R23 B.n133 B.n132 585
R24 B.n131 B.n130 585
R25 B.n129 B.n128 585
R26 B.n127 B.n126 585
R27 B.n125 B.n124 585
R28 B.n123 B.n122 585
R29 B.n121 B.n120 585
R30 B.n119 B.n118 585
R31 B.n117 B.n116 585
R32 B.n115 B.n114 585
R33 B.n113 B.n112 585
R34 B.n111 B.n110 585
R35 B.n109 B.n108 585
R36 B.n107 B.n106 585
R37 B.n105 B.n104 585
R38 B.n103 B.n102 585
R39 B.n101 B.n100 585
R40 B.n99 B.n98 585
R41 B.n97 B.n96 585
R42 B.n95 B.n94 585
R43 B.n93 B.n92 585
R44 B.n91 B.n90 585
R45 B.n89 B.n88 585
R46 B.n87 B.n86 585
R47 B.n85 B.n84 585
R48 B.n83 B.n82 585
R49 B.n81 B.n80 585
R50 B.n79 B.n78 585
R51 B.n77 B.n76 585
R52 B.n75 B.n74 585
R53 B.n40 B.n39 585
R54 B.n439 B.n41 585
R55 B.n443 B.n41 585
R56 B.n438 B.n437 585
R57 B.n437 B.n37 585
R58 B.n436 B.n36 585
R59 B.n449 B.n36 585
R60 B.n435 B.n35 585
R61 B.n450 B.n35 585
R62 B.n434 B.n34 585
R63 B.n451 B.n34 585
R64 B.n433 B.n432 585
R65 B.n432 B.n30 585
R66 B.n431 B.n29 585
R67 B.n457 B.n29 585
R68 B.n430 B.n28 585
R69 B.n458 B.n28 585
R70 B.n429 B.n27 585
R71 B.n459 B.n27 585
R72 B.n428 B.n427 585
R73 B.n427 B.n26 585
R74 B.n426 B.n22 585
R75 B.n465 B.n22 585
R76 B.n425 B.n21 585
R77 B.n466 B.n21 585
R78 B.n424 B.n20 585
R79 B.n467 B.n20 585
R80 B.n423 B.n422 585
R81 B.n422 B.n19 585
R82 B.n421 B.n15 585
R83 B.n473 B.n15 585
R84 B.n420 B.n14 585
R85 B.n474 B.n14 585
R86 B.n419 B.n13 585
R87 B.n475 B.n13 585
R88 B.n418 B.n417 585
R89 B.n417 B.n12 585
R90 B.n416 B.n415 585
R91 B.n416 B.n8 585
R92 B.n414 B.n7 585
R93 B.n482 B.n7 585
R94 B.n413 B.n6 585
R95 B.n483 B.n6 585
R96 B.n412 B.n5 585
R97 B.n484 B.n5 585
R98 B.n411 B.n410 585
R99 B.n410 B.n4 585
R100 B.n409 B.n176 585
R101 B.n409 B.n408 585
R102 B.n398 B.n177 585
R103 B.n401 B.n177 585
R104 B.n400 B.n399 585
R105 B.n402 B.n400 585
R106 B.n397 B.n181 585
R107 B.n184 B.n181 585
R108 B.n396 B.n395 585
R109 B.n395 B.n394 585
R110 B.n183 B.n182 585
R111 B.n387 B.n183 585
R112 B.n386 B.n385 585
R113 B.n388 B.n386 585
R114 B.n384 B.n188 585
R115 B.n191 B.n188 585
R116 B.n383 B.n382 585
R117 B.n382 B.n381 585
R118 B.n190 B.n189 585
R119 B.n374 B.n190 585
R120 B.n373 B.n372 585
R121 B.n375 B.n373 585
R122 B.n371 B.n196 585
R123 B.n196 B.n195 585
R124 B.n370 B.n369 585
R125 B.n369 B.n368 585
R126 B.n198 B.n197 585
R127 B.n199 B.n198 585
R128 B.n361 B.n360 585
R129 B.n362 B.n361 585
R130 B.n359 B.n204 585
R131 B.n204 B.n203 585
R132 B.n358 B.n357 585
R133 B.n357 B.n356 585
R134 B.n206 B.n205 585
R135 B.n207 B.n206 585
R136 B.n349 B.n348 585
R137 B.n350 B.n349 585
R138 B.n210 B.n209 585
R139 B.n243 B.n241 585
R140 B.n244 B.n240 585
R141 B.n244 B.n211 585
R142 B.n247 B.n246 585
R143 B.n248 B.n239 585
R144 B.n250 B.n249 585
R145 B.n252 B.n238 585
R146 B.n255 B.n254 585
R147 B.n256 B.n237 585
R148 B.n258 B.n257 585
R149 B.n260 B.n236 585
R150 B.n263 B.n262 585
R151 B.n264 B.n235 585
R152 B.n266 B.n265 585
R153 B.n268 B.n234 585
R154 B.n271 B.n270 585
R155 B.n272 B.n233 585
R156 B.n274 B.n273 585
R157 B.n276 B.n232 585
R158 B.n279 B.n278 585
R159 B.n280 B.n231 585
R160 B.n285 B.n284 585
R161 B.n287 B.n230 585
R162 B.n290 B.n289 585
R163 B.n291 B.n229 585
R164 B.n293 B.n292 585
R165 B.n295 B.n228 585
R166 B.n298 B.n297 585
R167 B.n299 B.n227 585
R168 B.n301 B.n300 585
R169 B.n303 B.n226 585
R170 B.n306 B.n305 585
R171 B.n307 B.n222 585
R172 B.n309 B.n308 585
R173 B.n311 B.n221 585
R174 B.n314 B.n313 585
R175 B.n315 B.n220 585
R176 B.n317 B.n316 585
R177 B.n319 B.n219 585
R178 B.n322 B.n321 585
R179 B.n323 B.n218 585
R180 B.n325 B.n324 585
R181 B.n327 B.n217 585
R182 B.n330 B.n329 585
R183 B.n331 B.n216 585
R184 B.n333 B.n332 585
R185 B.n335 B.n215 585
R186 B.n338 B.n337 585
R187 B.n339 B.n214 585
R188 B.n341 B.n340 585
R189 B.n343 B.n213 585
R190 B.n346 B.n345 585
R191 B.n347 B.n212 585
R192 B.n352 B.n351 585
R193 B.n351 B.n350 585
R194 B.n353 B.n208 585
R195 B.n208 B.n207 585
R196 B.n355 B.n354 585
R197 B.n356 B.n355 585
R198 B.n202 B.n201 585
R199 B.n203 B.n202 585
R200 B.n364 B.n363 585
R201 B.n363 B.n362 585
R202 B.n365 B.n200 585
R203 B.n200 B.n199 585
R204 B.n367 B.n366 585
R205 B.n368 B.n367 585
R206 B.n194 B.n193 585
R207 B.n195 B.n194 585
R208 B.n377 B.n376 585
R209 B.n376 B.n375 585
R210 B.n378 B.n192 585
R211 B.n374 B.n192 585
R212 B.n380 B.n379 585
R213 B.n381 B.n380 585
R214 B.n187 B.n186 585
R215 B.n191 B.n187 585
R216 B.n390 B.n389 585
R217 B.n389 B.n388 585
R218 B.n391 B.n185 585
R219 B.n387 B.n185 585
R220 B.n393 B.n392 585
R221 B.n394 B.n393 585
R222 B.n180 B.n179 585
R223 B.n184 B.n180 585
R224 B.n404 B.n403 585
R225 B.n403 B.n402 585
R226 B.n405 B.n178 585
R227 B.n401 B.n178 585
R228 B.n407 B.n406 585
R229 B.n408 B.n407 585
R230 B.n3 B.n0 585
R231 B.n4 B.n3 585
R232 B.n481 B.n1 585
R233 B.n482 B.n481 585
R234 B.n480 B.n479 585
R235 B.n480 B.n8 585
R236 B.n478 B.n9 585
R237 B.n12 B.n9 585
R238 B.n477 B.n476 585
R239 B.n476 B.n475 585
R240 B.n11 B.n10 585
R241 B.n474 B.n11 585
R242 B.n472 B.n471 585
R243 B.n473 B.n472 585
R244 B.n470 B.n16 585
R245 B.n19 B.n16 585
R246 B.n469 B.n468 585
R247 B.n468 B.n467 585
R248 B.n18 B.n17 585
R249 B.n466 B.n18 585
R250 B.n464 B.n463 585
R251 B.n465 B.n464 585
R252 B.n462 B.n23 585
R253 B.n26 B.n23 585
R254 B.n461 B.n460 585
R255 B.n460 B.n459 585
R256 B.n25 B.n24 585
R257 B.n458 B.n25 585
R258 B.n456 B.n455 585
R259 B.n457 B.n456 585
R260 B.n454 B.n31 585
R261 B.n31 B.n30 585
R262 B.n453 B.n452 585
R263 B.n452 B.n451 585
R264 B.n33 B.n32 585
R265 B.n450 B.n33 585
R266 B.n448 B.n447 585
R267 B.n449 B.n448 585
R268 B.n446 B.n38 585
R269 B.n38 B.n37 585
R270 B.n445 B.n444 585
R271 B.n444 B.n443 585
R272 B.n485 B.n484 585
R273 B.n483 B.n2 585
R274 B.n71 B.t17 553.904
R275 B.n69 B.t21 553.904
R276 B.n223 B.t14 553.904
R277 B.n281 B.t10 553.904
R278 B.n444 B.n40 511.721
R279 B.n441 B.n41 511.721
R280 B.n349 B.n212 511.721
R281 B.n351 B.n210 511.721
R282 B.n442 B.n67 256.663
R283 B.n442 B.n66 256.663
R284 B.n442 B.n65 256.663
R285 B.n442 B.n64 256.663
R286 B.n442 B.n63 256.663
R287 B.n442 B.n62 256.663
R288 B.n442 B.n61 256.663
R289 B.n442 B.n60 256.663
R290 B.n442 B.n59 256.663
R291 B.n442 B.n58 256.663
R292 B.n442 B.n57 256.663
R293 B.n442 B.n56 256.663
R294 B.n442 B.n55 256.663
R295 B.n442 B.n54 256.663
R296 B.n442 B.n53 256.663
R297 B.n442 B.n52 256.663
R298 B.n442 B.n51 256.663
R299 B.n442 B.n50 256.663
R300 B.n442 B.n49 256.663
R301 B.n442 B.n48 256.663
R302 B.n442 B.n47 256.663
R303 B.n442 B.n46 256.663
R304 B.n442 B.n45 256.663
R305 B.n442 B.n44 256.663
R306 B.n442 B.n43 256.663
R307 B.n442 B.n42 256.663
R308 B.n242 B.n211 256.663
R309 B.n245 B.n211 256.663
R310 B.n251 B.n211 256.663
R311 B.n253 B.n211 256.663
R312 B.n259 B.n211 256.663
R313 B.n261 B.n211 256.663
R314 B.n267 B.n211 256.663
R315 B.n269 B.n211 256.663
R316 B.n275 B.n211 256.663
R317 B.n277 B.n211 256.663
R318 B.n286 B.n211 256.663
R319 B.n288 B.n211 256.663
R320 B.n294 B.n211 256.663
R321 B.n296 B.n211 256.663
R322 B.n302 B.n211 256.663
R323 B.n304 B.n211 256.663
R324 B.n310 B.n211 256.663
R325 B.n312 B.n211 256.663
R326 B.n318 B.n211 256.663
R327 B.n320 B.n211 256.663
R328 B.n326 B.n211 256.663
R329 B.n328 B.n211 256.663
R330 B.n334 B.n211 256.663
R331 B.n336 B.n211 256.663
R332 B.n342 B.n211 256.663
R333 B.n344 B.n211 256.663
R334 B.n487 B.n486 256.663
R335 B.n69 B.t22 179.956
R336 B.n223 B.t16 179.956
R337 B.n71 B.t19 179.956
R338 B.n281 B.t13 179.956
R339 B.n70 B.t23 166.38
R340 B.n224 B.t15 166.38
R341 B.n72 B.t20 166.38
R342 B.n282 B.t12 166.38
R343 B.n76 B.n75 163.367
R344 B.n80 B.n79 163.367
R345 B.n84 B.n83 163.367
R346 B.n88 B.n87 163.367
R347 B.n92 B.n91 163.367
R348 B.n96 B.n95 163.367
R349 B.n100 B.n99 163.367
R350 B.n104 B.n103 163.367
R351 B.n108 B.n107 163.367
R352 B.n112 B.n111 163.367
R353 B.n116 B.n115 163.367
R354 B.n120 B.n119 163.367
R355 B.n124 B.n123 163.367
R356 B.n128 B.n127 163.367
R357 B.n132 B.n131 163.367
R358 B.n137 B.n136 163.367
R359 B.n141 B.n140 163.367
R360 B.n145 B.n144 163.367
R361 B.n149 B.n148 163.367
R362 B.n153 B.n152 163.367
R363 B.n157 B.n156 163.367
R364 B.n161 B.n160 163.367
R365 B.n165 B.n164 163.367
R366 B.n169 B.n168 163.367
R367 B.n173 B.n172 163.367
R368 B.n441 B.n68 163.367
R369 B.n349 B.n206 163.367
R370 B.n357 B.n206 163.367
R371 B.n357 B.n204 163.367
R372 B.n361 B.n204 163.367
R373 B.n361 B.n198 163.367
R374 B.n369 B.n198 163.367
R375 B.n369 B.n196 163.367
R376 B.n373 B.n196 163.367
R377 B.n373 B.n190 163.367
R378 B.n382 B.n190 163.367
R379 B.n382 B.n188 163.367
R380 B.n386 B.n188 163.367
R381 B.n386 B.n183 163.367
R382 B.n395 B.n183 163.367
R383 B.n395 B.n181 163.367
R384 B.n400 B.n181 163.367
R385 B.n400 B.n177 163.367
R386 B.n409 B.n177 163.367
R387 B.n410 B.n409 163.367
R388 B.n410 B.n5 163.367
R389 B.n6 B.n5 163.367
R390 B.n7 B.n6 163.367
R391 B.n416 B.n7 163.367
R392 B.n417 B.n416 163.367
R393 B.n417 B.n13 163.367
R394 B.n14 B.n13 163.367
R395 B.n15 B.n14 163.367
R396 B.n422 B.n15 163.367
R397 B.n422 B.n20 163.367
R398 B.n21 B.n20 163.367
R399 B.n22 B.n21 163.367
R400 B.n427 B.n22 163.367
R401 B.n427 B.n27 163.367
R402 B.n28 B.n27 163.367
R403 B.n29 B.n28 163.367
R404 B.n432 B.n29 163.367
R405 B.n432 B.n34 163.367
R406 B.n35 B.n34 163.367
R407 B.n36 B.n35 163.367
R408 B.n437 B.n36 163.367
R409 B.n437 B.n41 163.367
R410 B.n244 B.n243 163.367
R411 B.n246 B.n244 163.367
R412 B.n250 B.n239 163.367
R413 B.n254 B.n252 163.367
R414 B.n258 B.n237 163.367
R415 B.n262 B.n260 163.367
R416 B.n266 B.n235 163.367
R417 B.n270 B.n268 163.367
R418 B.n274 B.n233 163.367
R419 B.n278 B.n276 163.367
R420 B.n285 B.n231 163.367
R421 B.n289 B.n287 163.367
R422 B.n293 B.n229 163.367
R423 B.n297 B.n295 163.367
R424 B.n301 B.n227 163.367
R425 B.n305 B.n303 163.367
R426 B.n309 B.n222 163.367
R427 B.n313 B.n311 163.367
R428 B.n317 B.n220 163.367
R429 B.n321 B.n319 163.367
R430 B.n325 B.n218 163.367
R431 B.n329 B.n327 163.367
R432 B.n333 B.n216 163.367
R433 B.n337 B.n335 163.367
R434 B.n341 B.n214 163.367
R435 B.n345 B.n343 163.367
R436 B.n351 B.n208 163.367
R437 B.n355 B.n208 163.367
R438 B.n355 B.n202 163.367
R439 B.n363 B.n202 163.367
R440 B.n363 B.n200 163.367
R441 B.n367 B.n200 163.367
R442 B.n367 B.n194 163.367
R443 B.n376 B.n194 163.367
R444 B.n376 B.n192 163.367
R445 B.n380 B.n192 163.367
R446 B.n380 B.n187 163.367
R447 B.n389 B.n187 163.367
R448 B.n389 B.n185 163.367
R449 B.n393 B.n185 163.367
R450 B.n393 B.n180 163.367
R451 B.n403 B.n180 163.367
R452 B.n403 B.n178 163.367
R453 B.n407 B.n178 163.367
R454 B.n407 B.n3 163.367
R455 B.n485 B.n3 163.367
R456 B.n481 B.n2 163.367
R457 B.n481 B.n480 163.367
R458 B.n480 B.n9 163.367
R459 B.n476 B.n9 163.367
R460 B.n476 B.n11 163.367
R461 B.n472 B.n11 163.367
R462 B.n472 B.n16 163.367
R463 B.n468 B.n16 163.367
R464 B.n468 B.n18 163.367
R465 B.n464 B.n18 163.367
R466 B.n464 B.n23 163.367
R467 B.n460 B.n23 163.367
R468 B.n460 B.n25 163.367
R469 B.n456 B.n25 163.367
R470 B.n456 B.n31 163.367
R471 B.n452 B.n31 163.367
R472 B.n452 B.n33 163.367
R473 B.n448 B.n33 163.367
R474 B.n448 B.n38 163.367
R475 B.n444 B.n38 163.367
R476 B.n350 B.n211 126.222
R477 B.n443 B.n442 126.222
R478 B.n42 B.n40 71.676
R479 B.n76 B.n43 71.676
R480 B.n80 B.n44 71.676
R481 B.n84 B.n45 71.676
R482 B.n88 B.n46 71.676
R483 B.n92 B.n47 71.676
R484 B.n96 B.n48 71.676
R485 B.n100 B.n49 71.676
R486 B.n104 B.n50 71.676
R487 B.n108 B.n51 71.676
R488 B.n112 B.n52 71.676
R489 B.n116 B.n53 71.676
R490 B.n120 B.n54 71.676
R491 B.n124 B.n55 71.676
R492 B.n128 B.n56 71.676
R493 B.n132 B.n57 71.676
R494 B.n137 B.n58 71.676
R495 B.n141 B.n59 71.676
R496 B.n145 B.n60 71.676
R497 B.n149 B.n61 71.676
R498 B.n153 B.n62 71.676
R499 B.n157 B.n63 71.676
R500 B.n161 B.n64 71.676
R501 B.n165 B.n65 71.676
R502 B.n169 B.n66 71.676
R503 B.n173 B.n67 71.676
R504 B.n68 B.n67 71.676
R505 B.n172 B.n66 71.676
R506 B.n168 B.n65 71.676
R507 B.n164 B.n64 71.676
R508 B.n160 B.n63 71.676
R509 B.n156 B.n62 71.676
R510 B.n152 B.n61 71.676
R511 B.n148 B.n60 71.676
R512 B.n144 B.n59 71.676
R513 B.n140 B.n58 71.676
R514 B.n136 B.n57 71.676
R515 B.n131 B.n56 71.676
R516 B.n127 B.n55 71.676
R517 B.n123 B.n54 71.676
R518 B.n119 B.n53 71.676
R519 B.n115 B.n52 71.676
R520 B.n111 B.n51 71.676
R521 B.n107 B.n50 71.676
R522 B.n103 B.n49 71.676
R523 B.n99 B.n48 71.676
R524 B.n95 B.n47 71.676
R525 B.n91 B.n46 71.676
R526 B.n87 B.n45 71.676
R527 B.n83 B.n44 71.676
R528 B.n79 B.n43 71.676
R529 B.n75 B.n42 71.676
R530 B.n242 B.n210 71.676
R531 B.n246 B.n245 71.676
R532 B.n251 B.n250 71.676
R533 B.n254 B.n253 71.676
R534 B.n259 B.n258 71.676
R535 B.n262 B.n261 71.676
R536 B.n267 B.n266 71.676
R537 B.n270 B.n269 71.676
R538 B.n275 B.n274 71.676
R539 B.n278 B.n277 71.676
R540 B.n286 B.n285 71.676
R541 B.n289 B.n288 71.676
R542 B.n294 B.n293 71.676
R543 B.n297 B.n296 71.676
R544 B.n302 B.n301 71.676
R545 B.n305 B.n304 71.676
R546 B.n310 B.n309 71.676
R547 B.n313 B.n312 71.676
R548 B.n318 B.n317 71.676
R549 B.n321 B.n320 71.676
R550 B.n326 B.n325 71.676
R551 B.n329 B.n328 71.676
R552 B.n334 B.n333 71.676
R553 B.n337 B.n336 71.676
R554 B.n342 B.n341 71.676
R555 B.n345 B.n344 71.676
R556 B.n243 B.n242 71.676
R557 B.n245 B.n239 71.676
R558 B.n252 B.n251 71.676
R559 B.n253 B.n237 71.676
R560 B.n260 B.n259 71.676
R561 B.n261 B.n235 71.676
R562 B.n268 B.n267 71.676
R563 B.n269 B.n233 71.676
R564 B.n276 B.n275 71.676
R565 B.n277 B.n231 71.676
R566 B.n287 B.n286 71.676
R567 B.n288 B.n229 71.676
R568 B.n295 B.n294 71.676
R569 B.n296 B.n227 71.676
R570 B.n303 B.n302 71.676
R571 B.n304 B.n222 71.676
R572 B.n311 B.n310 71.676
R573 B.n312 B.n220 71.676
R574 B.n319 B.n318 71.676
R575 B.n320 B.n218 71.676
R576 B.n327 B.n326 71.676
R577 B.n328 B.n216 71.676
R578 B.n335 B.n334 71.676
R579 B.n336 B.n214 71.676
R580 B.n343 B.n342 71.676
R581 B.n344 B.n212 71.676
R582 B.n486 B.n485 71.676
R583 B.n486 B.n2 71.676
R584 B.n350 B.n207 70.9346
R585 B.n356 B.n207 70.9346
R586 B.n356 B.n203 70.9346
R587 B.n362 B.n203 70.9346
R588 B.n368 B.n199 70.9346
R589 B.n368 B.n195 70.9346
R590 B.n375 B.n195 70.9346
R591 B.n375 B.n374 70.9346
R592 B.n381 B.n191 70.9346
R593 B.n388 B.n387 70.9346
R594 B.n394 B.n184 70.9346
R595 B.n402 B.n401 70.9346
R596 B.n408 B.n4 70.9346
R597 B.n484 B.n4 70.9346
R598 B.n484 B.n483 70.9346
R599 B.n483 B.n482 70.9346
R600 B.n482 B.n8 70.9346
R601 B.n475 B.n12 70.9346
R602 B.n474 B.n473 70.9346
R603 B.n467 B.n19 70.9346
R604 B.n466 B.n465 70.9346
R605 B.n459 B.n26 70.9346
R606 B.n459 B.n458 70.9346
R607 B.n458 B.n457 70.9346
R608 B.n457 B.n30 70.9346
R609 B.n451 B.n450 70.9346
R610 B.n450 B.n449 70.9346
R611 B.n449 B.n37 70.9346
R612 B.n443 B.n37 70.9346
R613 B.n401 B.t8 61.5463
R614 B.n12 B.t7 61.5463
R615 B.n73 B.n72 59.5399
R616 B.n134 B.n70 59.5399
R617 B.n225 B.n224 59.5399
R618 B.n283 B.n282 59.5399
R619 B.n184 B.t2 57.3737
R620 B.t9 B.n474 57.3737
R621 B.n387 B.t1 53.2011
R622 B.n19 B.t0 53.2011
R623 B.n191 B.t3 49.0285
R624 B.t4 B.n466 49.0285
R625 B.t11 B.n199 44.8559
R626 B.n374 B.t5 44.8559
R627 B.n26 B.t6 44.8559
R628 B.t18 B.n30 44.8559
R629 B.n352 B.n209 33.2493
R630 B.n348 B.n347 33.2493
R631 B.n440 B.n439 33.2493
R632 B.n445 B.n39 33.2493
R633 B.n362 B.t11 26.0792
R634 B.n381 B.t5 26.0792
R635 B.n465 B.t6 26.0792
R636 B.n451 B.t18 26.0792
R637 B.n388 B.t3 21.9066
R638 B.n467 B.t4 21.9066
R639 B B.n487 18.0485
R640 B.n394 B.t1 17.734
R641 B.n473 B.t0 17.734
R642 B.n72 B.n71 13.5763
R643 B.n70 B.n69 13.5763
R644 B.n224 B.n223 13.5763
R645 B.n282 B.n281 13.5763
R646 B.n402 B.t2 13.5614
R647 B.n475 B.t9 13.5614
R648 B.n353 B.n352 10.6151
R649 B.n354 B.n353 10.6151
R650 B.n354 B.n201 10.6151
R651 B.n364 B.n201 10.6151
R652 B.n365 B.n364 10.6151
R653 B.n366 B.n365 10.6151
R654 B.n366 B.n193 10.6151
R655 B.n377 B.n193 10.6151
R656 B.n378 B.n377 10.6151
R657 B.n379 B.n378 10.6151
R658 B.n379 B.n186 10.6151
R659 B.n390 B.n186 10.6151
R660 B.n391 B.n390 10.6151
R661 B.n392 B.n391 10.6151
R662 B.n392 B.n179 10.6151
R663 B.n404 B.n179 10.6151
R664 B.n405 B.n404 10.6151
R665 B.n406 B.n405 10.6151
R666 B.n406 B.n0 10.6151
R667 B.n241 B.n209 10.6151
R668 B.n241 B.n240 10.6151
R669 B.n247 B.n240 10.6151
R670 B.n248 B.n247 10.6151
R671 B.n249 B.n248 10.6151
R672 B.n249 B.n238 10.6151
R673 B.n255 B.n238 10.6151
R674 B.n256 B.n255 10.6151
R675 B.n257 B.n256 10.6151
R676 B.n257 B.n236 10.6151
R677 B.n263 B.n236 10.6151
R678 B.n264 B.n263 10.6151
R679 B.n265 B.n264 10.6151
R680 B.n265 B.n234 10.6151
R681 B.n271 B.n234 10.6151
R682 B.n272 B.n271 10.6151
R683 B.n273 B.n272 10.6151
R684 B.n273 B.n232 10.6151
R685 B.n279 B.n232 10.6151
R686 B.n280 B.n279 10.6151
R687 B.n284 B.n280 10.6151
R688 B.n290 B.n230 10.6151
R689 B.n291 B.n290 10.6151
R690 B.n292 B.n291 10.6151
R691 B.n292 B.n228 10.6151
R692 B.n298 B.n228 10.6151
R693 B.n299 B.n298 10.6151
R694 B.n300 B.n299 10.6151
R695 B.n300 B.n226 10.6151
R696 B.n307 B.n306 10.6151
R697 B.n308 B.n307 10.6151
R698 B.n308 B.n221 10.6151
R699 B.n314 B.n221 10.6151
R700 B.n315 B.n314 10.6151
R701 B.n316 B.n315 10.6151
R702 B.n316 B.n219 10.6151
R703 B.n322 B.n219 10.6151
R704 B.n323 B.n322 10.6151
R705 B.n324 B.n323 10.6151
R706 B.n324 B.n217 10.6151
R707 B.n330 B.n217 10.6151
R708 B.n331 B.n330 10.6151
R709 B.n332 B.n331 10.6151
R710 B.n332 B.n215 10.6151
R711 B.n338 B.n215 10.6151
R712 B.n339 B.n338 10.6151
R713 B.n340 B.n339 10.6151
R714 B.n340 B.n213 10.6151
R715 B.n346 B.n213 10.6151
R716 B.n347 B.n346 10.6151
R717 B.n348 B.n205 10.6151
R718 B.n358 B.n205 10.6151
R719 B.n359 B.n358 10.6151
R720 B.n360 B.n359 10.6151
R721 B.n360 B.n197 10.6151
R722 B.n370 B.n197 10.6151
R723 B.n371 B.n370 10.6151
R724 B.n372 B.n371 10.6151
R725 B.n372 B.n189 10.6151
R726 B.n383 B.n189 10.6151
R727 B.n384 B.n383 10.6151
R728 B.n385 B.n384 10.6151
R729 B.n385 B.n182 10.6151
R730 B.n396 B.n182 10.6151
R731 B.n397 B.n396 10.6151
R732 B.n399 B.n397 10.6151
R733 B.n399 B.n398 10.6151
R734 B.n398 B.n176 10.6151
R735 B.n411 B.n176 10.6151
R736 B.n412 B.n411 10.6151
R737 B.n413 B.n412 10.6151
R738 B.n414 B.n413 10.6151
R739 B.n415 B.n414 10.6151
R740 B.n418 B.n415 10.6151
R741 B.n419 B.n418 10.6151
R742 B.n420 B.n419 10.6151
R743 B.n421 B.n420 10.6151
R744 B.n423 B.n421 10.6151
R745 B.n424 B.n423 10.6151
R746 B.n425 B.n424 10.6151
R747 B.n426 B.n425 10.6151
R748 B.n428 B.n426 10.6151
R749 B.n429 B.n428 10.6151
R750 B.n430 B.n429 10.6151
R751 B.n431 B.n430 10.6151
R752 B.n433 B.n431 10.6151
R753 B.n434 B.n433 10.6151
R754 B.n435 B.n434 10.6151
R755 B.n436 B.n435 10.6151
R756 B.n438 B.n436 10.6151
R757 B.n439 B.n438 10.6151
R758 B.n479 B.n1 10.6151
R759 B.n479 B.n478 10.6151
R760 B.n478 B.n477 10.6151
R761 B.n477 B.n10 10.6151
R762 B.n471 B.n10 10.6151
R763 B.n471 B.n470 10.6151
R764 B.n470 B.n469 10.6151
R765 B.n469 B.n17 10.6151
R766 B.n463 B.n17 10.6151
R767 B.n463 B.n462 10.6151
R768 B.n462 B.n461 10.6151
R769 B.n461 B.n24 10.6151
R770 B.n455 B.n24 10.6151
R771 B.n455 B.n454 10.6151
R772 B.n454 B.n453 10.6151
R773 B.n453 B.n32 10.6151
R774 B.n447 B.n32 10.6151
R775 B.n447 B.n446 10.6151
R776 B.n446 B.n445 10.6151
R777 B.n74 B.n39 10.6151
R778 B.n77 B.n74 10.6151
R779 B.n78 B.n77 10.6151
R780 B.n81 B.n78 10.6151
R781 B.n82 B.n81 10.6151
R782 B.n85 B.n82 10.6151
R783 B.n86 B.n85 10.6151
R784 B.n89 B.n86 10.6151
R785 B.n90 B.n89 10.6151
R786 B.n93 B.n90 10.6151
R787 B.n94 B.n93 10.6151
R788 B.n97 B.n94 10.6151
R789 B.n98 B.n97 10.6151
R790 B.n101 B.n98 10.6151
R791 B.n102 B.n101 10.6151
R792 B.n105 B.n102 10.6151
R793 B.n106 B.n105 10.6151
R794 B.n109 B.n106 10.6151
R795 B.n110 B.n109 10.6151
R796 B.n113 B.n110 10.6151
R797 B.n114 B.n113 10.6151
R798 B.n118 B.n117 10.6151
R799 B.n121 B.n118 10.6151
R800 B.n122 B.n121 10.6151
R801 B.n125 B.n122 10.6151
R802 B.n126 B.n125 10.6151
R803 B.n129 B.n126 10.6151
R804 B.n130 B.n129 10.6151
R805 B.n133 B.n130 10.6151
R806 B.n138 B.n135 10.6151
R807 B.n139 B.n138 10.6151
R808 B.n142 B.n139 10.6151
R809 B.n143 B.n142 10.6151
R810 B.n146 B.n143 10.6151
R811 B.n147 B.n146 10.6151
R812 B.n150 B.n147 10.6151
R813 B.n151 B.n150 10.6151
R814 B.n154 B.n151 10.6151
R815 B.n155 B.n154 10.6151
R816 B.n158 B.n155 10.6151
R817 B.n159 B.n158 10.6151
R818 B.n162 B.n159 10.6151
R819 B.n163 B.n162 10.6151
R820 B.n166 B.n163 10.6151
R821 B.n167 B.n166 10.6151
R822 B.n170 B.n167 10.6151
R823 B.n171 B.n170 10.6151
R824 B.n174 B.n171 10.6151
R825 B.n175 B.n174 10.6151
R826 B.n440 B.n175 10.6151
R827 B.n408 B.t8 9.38884
R828 B.t7 B.n8 9.38884
R829 B.n487 B.n0 8.11757
R830 B.n487 B.n1 8.11757
R831 B.n283 B.n230 6.5566
R832 B.n226 B.n225 6.5566
R833 B.n117 B.n73 6.5566
R834 B.n134 B.n133 6.5566
R835 B.n284 B.n283 4.05904
R836 B.n306 B.n225 4.05904
R837 B.n114 B.n73 4.05904
R838 B.n135 B.n134 4.05904
R839 VP.n5 VP.t7 471.065
R840 VP.n15 VP.t5 450.084
R841 VP.n16 VP.t2 450.084
R842 VP.n1 VP.t3 450.084
R843 VP.n21 VP.t8 450.084
R844 VP.n22 VP.t0 450.084
R845 VP.n12 VP.t6 450.084
R846 VP.n11 VP.t9 450.084
R847 VP.n4 VP.t1 450.084
R848 VP.n6 VP.t4 450.084
R849 VP.n23 VP.n22 161.3
R850 VP.n8 VP.n7 161.3
R851 VP.n10 VP.n9 161.3
R852 VP.n11 VP.n3 161.3
R853 VP.n13 VP.n12 161.3
R854 VP.n21 VP.n0 161.3
R855 VP.n20 VP.n19 161.3
R856 VP.n18 VP.n17 161.3
R857 VP.n16 VP.n2 161.3
R858 VP.n15 VP.n14 161.3
R859 VP.n8 VP.n5 70.4033
R860 VP.n16 VP.n15 48.2005
R861 VP.n22 VP.n21 48.2005
R862 VP.n12 VP.n11 48.2005
R863 VP.n17 VP.n16 38.7066
R864 VP.n21 VP.n20 38.7066
R865 VP.n11 VP.n10 38.7066
R866 VP.n7 VP.n6 38.7066
R867 VP.n14 VP.n13 35.8793
R868 VP.n6 VP.n5 20.9576
R869 VP.n17 VP.n1 9.49444
R870 VP.n20 VP.n1 9.49444
R871 VP.n10 VP.n4 9.49444
R872 VP.n7 VP.n4 9.49444
R873 VP.n9 VP.n8 0.189894
R874 VP.n9 VP.n3 0.189894
R875 VP.n13 VP.n3 0.189894
R876 VP.n14 VP.n2 0.189894
R877 VP.n18 VP.n2 0.189894
R878 VP.n19 VP.n18 0.189894
R879 VP.n19 VP.n0 0.189894
R880 VP.n23 VP.n0 0.189894
R881 VP VP.n23 0.0516364
R882 VTAIL.n120 VTAIL.n98 289.615
R883 VTAIL.n24 VTAIL.n2 289.615
R884 VTAIL.n92 VTAIL.n70 289.615
R885 VTAIL.n60 VTAIL.n38 289.615
R886 VTAIL.n106 VTAIL.n105 185
R887 VTAIL.n111 VTAIL.n110 185
R888 VTAIL.n113 VTAIL.n112 185
R889 VTAIL.n102 VTAIL.n101 185
R890 VTAIL.n119 VTAIL.n118 185
R891 VTAIL.n121 VTAIL.n120 185
R892 VTAIL.n10 VTAIL.n9 185
R893 VTAIL.n15 VTAIL.n14 185
R894 VTAIL.n17 VTAIL.n16 185
R895 VTAIL.n6 VTAIL.n5 185
R896 VTAIL.n23 VTAIL.n22 185
R897 VTAIL.n25 VTAIL.n24 185
R898 VTAIL.n93 VTAIL.n92 185
R899 VTAIL.n91 VTAIL.n90 185
R900 VTAIL.n74 VTAIL.n73 185
R901 VTAIL.n85 VTAIL.n84 185
R902 VTAIL.n83 VTAIL.n82 185
R903 VTAIL.n78 VTAIL.n77 185
R904 VTAIL.n61 VTAIL.n60 185
R905 VTAIL.n59 VTAIL.n58 185
R906 VTAIL.n42 VTAIL.n41 185
R907 VTAIL.n53 VTAIL.n52 185
R908 VTAIL.n51 VTAIL.n50 185
R909 VTAIL.n46 VTAIL.n45 185
R910 VTAIL.n107 VTAIL.t4 147.672
R911 VTAIL.n11 VTAIL.t15 147.672
R912 VTAIL.n79 VTAIL.t8 147.672
R913 VTAIL.n47 VTAIL.t17 147.672
R914 VTAIL.n111 VTAIL.n105 104.615
R915 VTAIL.n112 VTAIL.n111 104.615
R916 VTAIL.n112 VTAIL.n101 104.615
R917 VTAIL.n119 VTAIL.n101 104.615
R918 VTAIL.n120 VTAIL.n119 104.615
R919 VTAIL.n15 VTAIL.n9 104.615
R920 VTAIL.n16 VTAIL.n15 104.615
R921 VTAIL.n16 VTAIL.n5 104.615
R922 VTAIL.n23 VTAIL.n5 104.615
R923 VTAIL.n24 VTAIL.n23 104.615
R924 VTAIL.n92 VTAIL.n91 104.615
R925 VTAIL.n91 VTAIL.n73 104.615
R926 VTAIL.n84 VTAIL.n73 104.615
R927 VTAIL.n84 VTAIL.n83 104.615
R928 VTAIL.n83 VTAIL.n77 104.615
R929 VTAIL.n60 VTAIL.n59 104.615
R930 VTAIL.n59 VTAIL.n41 104.615
R931 VTAIL.n52 VTAIL.n41 104.615
R932 VTAIL.n52 VTAIL.n51 104.615
R933 VTAIL.n51 VTAIL.n45 104.615
R934 VTAIL.t4 VTAIL.n105 52.3082
R935 VTAIL.t15 VTAIL.n9 52.3082
R936 VTAIL.t8 VTAIL.n77 52.3082
R937 VTAIL.t17 VTAIL.n45 52.3082
R938 VTAIL.n69 VTAIL.n68 51.7825
R939 VTAIL.n67 VTAIL.n66 51.7825
R940 VTAIL.n37 VTAIL.n36 51.7825
R941 VTAIL.n35 VTAIL.n34 51.7825
R942 VTAIL.n127 VTAIL.n126 51.7824
R943 VTAIL.n1 VTAIL.n0 51.7824
R944 VTAIL.n31 VTAIL.n30 51.7824
R945 VTAIL.n33 VTAIL.n32 51.7824
R946 VTAIL.n125 VTAIL.n124 31.9914
R947 VTAIL.n29 VTAIL.n28 31.9914
R948 VTAIL.n97 VTAIL.n96 31.9914
R949 VTAIL.n65 VTAIL.n64 31.9914
R950 VTAIL.n35 VTAIL.n33 18.1169
R951 VTAIL.n125 VTAIL.n97 17.5134
R952 VTAIL.n107 VTAIL.n106 15.6666
R953 VTAIL.n11 VTAIL.n10 15.6666
R954 VTAIL.n79 VTAIL.n78 15.6666
R955 VTAIL.n47 VTAIL.n46 15.6666
R956 VTAIL.n110 VTAIL.n109 12.8005
R957 VTAIL.n14 VTAIL.n13 12.8005
R958 VTAIL.n82 VTAIL.n81 12.8005
R959 VTAIL.n50 VTAIL.n49 12.8005
R960 VTAIL.n113 VTAIL.n104 12.0247
R961 VTAIL.n17 VTAIL.n8 12.0247
R962 VTAIL.n85 VTAIL.n76 12.0247
R963 VTAIL.n53 VTAIL.n44 12.0247
R964 VTAIL.n114 VTAIL.n102 11.249
R965 VTAIL.n18 VTAIL.n6 11.249
R966 VTAIL.n86 VTAIL.n74 11.249
R967 VTAIL.n54 VTAIL.n42 11.249
R968 VTAIL.n118 VTAIL.n117 10.4732
R969 VTAIL.n22 VTAIL.n21 10.4732
R970 VTAIL.n90 VTAIL.n89 10.4732
R971 VTAIL.n58 VTAIL.n57 10.4732
R972 VTAIL.n121 VTAIL.n100 9.69747
R973 VTAIL.n25 VTAIL.n4 9.69747
R974 VTAIL.n93 VTAIL.n72 9.69747
R975 VTAIL.n61 VTAIL.n40 9.69747
R976 VTAIL.n124 VTAIL.n123 9.45567
R977 VTAIL.n28 VTAIL.n27 9.45567
R978 VTAIL.n96 VTAIL.n95 9.45567
R979 VTAIL.n64 VTAIL.n63 9.45567
R980 VTAIL.n123 VTAIL.n122 9.3005
R981 VTAIL.n100 VTAIL.n99 9.3005
R982 VTAIL.n117 VTAIL.n116 9.3005
R983 VTAIL.n115 VTAIL.n114 9.3005
R984 VTAIL.n104 VTAIL.n103 9.3005
R985 VTAIL.n109 VTAIL.n108 9.3005
R986 VTAIL.n27 VTAIL.n26 9.3005
R987 VTAIL.n4 VTAIL.n3 9.3005
R988 VTAIL.n21 VTAIL.n20 9.3005
R989 VTAIL.n19 VTAIL.n18 9.3005
R990 VTAIL.n8 VTAIL.n7 9.3005
R991 VTAIL.n13 VTAIL.n12 9.3005
R992 VTAIL.n95 VTAIL.n94 9.3005
R993 VTAIL.n72 VTAIL.n71 9.3005
R994 VTAIL.n89 VTAIL.n88 9.3005
R995 VTAIL.n87 VTAIL.n86 9.3005
R996 VTAIL.n76 VTAIL.n75 9.3005
R997 VTAIL.n81 VTAIL.n80 9.3005
R998 VTAIL.n63 VTAIL.n62 9.3005
R999 VTAIL.n40 VTAIL.n39 9.3005
R1000 VTAIL.n57 VTAIL.n56 9.3005
R1001 VTAIL.n55 VTAIL.n54 9.3005
R1002 VTAIL.n44 VTAIL.n43 9.3005
R1003 VTAIL.n49 VTAIL.n48 9.3005
R1004 VTAIL.n122 VTAIL.n98 8.92171
R1005 VTAIL.n26 VTAIL.n2 8.92171
R1006 VTAIL.n94 VTAIL.n70 8.92171
R1007 VTAIL.n62 VTAIL.n38 8.92171
R1008 VTAIL.n124 VTAIL.n98 5.04292
R1009 VTAIL.n28 VTAIL.n2 5.04292
R1010 VTAIL.n96 VTAIL.n70 5.04292
R1011 VTAIL.n64 VTAIL.n38 5.04292
R1012 VTAIL.n108 VTAIL.n107 4.38687
R1013 VTAIL.n12 VTAIL.n11 4.38687
R1014 VTAIL.n80 VTAIL.n79 4.38687
R1015 VTAIL.n48 VTAIL.n47 4.38687
R1016 VTAIL.n122 VTAIL.n121 4.26717
R1017 VTAIL.n26 VTAIL.n25 4.26717
R1018 VTAIL.n94 VTAIL.n93 4.26717
R1019 VTAIL.n62 VTAIL.n61 4.26717
R1020 VTAIL.n126 VTAIL.t5 3.75762
R1021 VTAIL.n126 VTAIL.t6 3.75762
R1022 VTAIL.n0 VTAIL.t19 3.75762
R1023 VTAIL.n0 VTAIL.t18 3.75762
R1024 VTAIL.n30 VTAIL.t12 3.75762
R1025 VTAIL.n30 VTAIL.t9 3.75762
R1026 VTAIL.n32 VTAIL.t10 3.75762
R1027 VTAIL.n32 VTAIL.t11 3.75762
R1028 VTAIL.n68 VTAIL.t14 3.75762
R1029 VTAIL.n68 VTAIL.t16 3.75762
R1030 VTAIL.n66 VTAIL.t7 3.75762
R1031 VTAIL.n66 VTAIL.t13 3.75762
R1032 VTAIL.n36 VTAIL.t0 3.75762
R1033 VTAIL.n36 VTAIL.t1 3.75762
R1034 VTAIL.n34 VTAIL.t3 3.75762
R1035 VTAIL.n34 VTAIL.t2 3.75762
R1036 VTAIL.n118 VTAIL.n100 3.49141
R1037 VTAIL.n22 VTAIL.n4 3.49141
R1038 VTAIL.n90 VTAIL.n72 3.49141
R1039 VTAIL.n58 VTAIL.n40 3.49141
R1040 VTAIL.n117 VTAIL.n102 2.71565
R1041 VTAIL.n21 VTAIL.n6 2.71565
R1042 VTAIL.n89 VTAIL.n74 2.71565
R1043 VTAIL.n57 VTAIL.n42 2.71565
R1044 VTAIL.n114 VTAIL.n113 1.93989
R1045 VTAIL.n18 VTAIL.n17 1.93989
R1046 VTAIL.n86 VTAIL.n85 1.93989
R1047 VTAIL.n54 VTAIL.n53 1.93989
R1048 VTAIL.n110 VTAIL.n104 1.16414
R1049 VTAIL.n14 VTAIL.n8 1.16414
R1050 VTAIL.n82 VTAIL.n76 1.16414
R1051 VTAIL.n50 VTAIL.n44 1.16414
R1052 VTAIL.n67 VTAIL.n65 0.772052
R1053 VTAIL.n29 VTAIL.n1 0.772052
R1054 VTAIL.n37 VTAIL.n35 0.603948
R1055 VTAIL.n65 VTAIL.n37 0.603948
R1056 VTAIL.n69 VTAIL.n67 0.603948
R1057 VTAIL.n97 VTAIL.n69 0.603948
R1058 VTAIL.n33 VTAIL.n31 0.603948
R1059 VTAIL.n31 VTAIL.n29 0.603948
R1060 VTAIL.n127 VTAIL.n125 0.603948
R1061 VTAIL VTAIL.n1 0.511276
R1062 VTAIL.n109 VTAIL.n106 0.388379
R1063 VTAIL.n13 VTAIL.n10 0.388379
R1064 VTAIL.n81 VTAIL.n78 0.388379
R1065 VTAIL.n49 VTAIL.n46 0.388379
R1066 VTAIL.n108 VTAIL.n103 0.155672
R1067 VTAIL.n115 VTAIL.n103 0.155672
R1068 VTAIL.n116 VTAIL.n115 0.155672
R1069 VTAIL.n116 VTAIL.n99 0.155672
R1070 VTAIL.n123 VTAIL.n99 0.155672
R1071 VTAIL.n12 VTAIL.n7 0.155672
R1072 VTAIL.n19 VTAIL.n7 0.155672
R1073 VTAIL.n20 VTAIL.n19 0.155672
R1074 VTAIL.n20 VTAIL.n3 0.155672
R1075 VTAIL.n27 VTAIL.n3 0.155672
R1076 VTAIL.n95 VTAIL.n71 0.155672
R1077 VTAIL.n88 VTAIL.n71 0.155672
R1078 VTAIL.n88 VTAIL.n87 0.155672
R1079 VTAIL.n87 VTAIL.n75 0.155672
R1080 VTAIL.n80 VTAIL.n75 0.155672
R1081 VTAIL.n63 VTAIL.n39 0.155672
R1082 VTAIL.n56 VTAIL.n39 0.155672
R1083 VTAIL.n56 VTAIL.n55 0.155672
R1084 VTAIL.n55 VTAIL.n43 0.155672
R1085 VTAIL.n48 VTAIL.n43 0.155672
R1086 VTAIL VTAIL.n127 0.0931724
R1087 VDD1.n22 VDD1.n0 289.615
R1088 VDD1.n51 VDD1.n29 289.615
R1089 VDD1.n23 VDD1.n22 185
R1090 VDD1.n21 VDD1.n20 185
R1091 VDD1.n4 VDD1.n3 185
R1092 VDD1.n15 VDD1.n14 185
R1093 VDD1.n13 VDD1.n12 185
R1094 VDD1.n8 VDD1.n7 185
R1095 VDD1.n37 VDD1.n36 185
R1096 VDD1.n42 VDD1.n41 185
R1097 VDD1.n44 VDD1.n43 185
R1098 VDD1.n33 VDD1.n32 185
R1099 VDD1.n50 VDD1.n49 185
R1100 VDD1.n52 VDD1.n51 185
R1101 VDD1.n9 VDD1.t2 147.672
R1102 VDD1.n38 VDD1.t4 147.672
R1103 VDD1.n22 VDD1.n21 104.615
R1104 VDD1.n21 VDD1.n3 104.615
R1105 VDD1.n14 VDD1.n3 104.615
R1106 VDD1.n14 VDD1.n13 104.615
R1107 VDD1.n13 VDD1.n7 104.615
R1108 VDD1.n42 VDD1.n36 104.615
R1109 VDD1.n43 VDD1.n42 104.615
R1110 VDD1.n43 VDD1.n32 104.615
R1111 VDD1.n50 VDD1.n32 104.615
R1112 VDD1.n51 VDD1.n50 104.615
R1113 VDD1.n59 VDD1.n58 68.8584
R1114 VDD1.n28 VDD1.n27 68.4613
R1115 VDD1.n61 VDD1.n60 68.4612
R1116 VDD1.n57 VDD1.n56 68.4612
R1117 VDD1.t2 VDD1.n7 52.3082
R1118 VDD1.t4 VDD1.n36 52.3082
R1119 VDD1.n28 VDD1.n26 49.2736
R1120 VDD1.n57 VDD1.n55 49.2736
R1121 VDD1.n61 VDD1.n59 32.0095
R1122 VDD1.n9 VDD1.n8 15.6666
R1123 VDD1.n38 VDD1.n37 15.6666
R1124 VDD1.n12 VDD1.n11 12.8005
R1125 VDD1.n41 VDD1.n40 12.8005
R1126 VDD1.n15 VDD1.n6 12.0247
R1127 VDD1.n44 VDD1.n35 12.0247
R1128 VDD1.n16 VDD1.n4 11.249
R1129 VDD1.n45 VDD1.n33 11.249
R1130 VDD1.n20 VDD1.n19 10.4732
R1131 VDD1.n49 VDD1.n48 10.4732
R1132 VDD1.n23 VDD1.n2 9.69747
R1133 VDD1.n52 VDD1.n31 9.69747
R1134 VDD1.n26 VDD1.n25 9.45567
R1135 VDD1.n55 VDD1.n54 9.45567
R1136 VDD1.n25 VDD1.n24 9.3005
R1137 VDD1.n2 VDD1.n1 9.3005
R1138 VDD1.n19 VDD1.n18 9.3005
R1139 VDD1.n17 VDD1.n16 9.3005
R1140 VDD1.n6 VDD1.n5 9.3005
R1141 VDD1.n11 VDD1.n10 9.3005
R1142 VDD1.n54 VDD1.n53 9.3005
R1143 VDD1.n31 VDD1.n30 9.3005
R1144 VDD1.n48 VDD1.n47 9.3005
R1145 VDD1.n46 VDD1.n45 9.3005
R1146 VDD1.n35 VDD1.n34 9.3005
R1147 VDD1.n40 VDD1.n39 9.3005
R1148 VDD1.n24 VDD1.n0 8.92171
R1149 VDD1.n53 VDD1.n29 8.92171
R1150 VDD1.n26 VDD1.n0 5.04292
R1151 VDD1.n55 VDD1.n29 5.04292
R1152 VDD1.n10 VDD1.n9 4.38687
R1153 VDD1.n39 VDD1.n38 4.38687
R1154 VDD1.n24 VDD1.n23 4.26717
R1155 VDD1.n53 VDD1.n52 4.26717
R1156 VDD1.n60 VDD1.t0 3.75762
R1157 VDD1.n60 VDD1.t3 3.75762
R1158 VDD1.n27 VDD1.t5 3.75762
R1159 VDD1.n27 VDD1.t8 3.75762
R1160 VDD1.n58 VDD1.t1 3.75762
R1161 VDD1.n58 VDD1.t9 3.75762
R1162 VDD1.n56 VDD1.t7 3.75762
R1163 VDD1.n56 VDD1.t6 3.75762
R1164 VDD1.n20 VDD1.n2 3.49141
R1165 VDD1.n49 VDD1.n31 3.49141
R1166 VDD1.n19 VDD1.n4 2.71565
R1167 VDD1.n48 VDD1.n33 2.71565
R1168 VDD1.n16 VDD1.n15 1.93989
R1169 VDD1.n45 VDD1.n44 1.93989
R1170 VDD1.n12 VDD1.n6 1.16414
R1171 VDD1.n41 VDD1.n35 1.16414
R1172 VDD1 VDD1.n61 0.394897
R1173 VDD1.n11 VDD1.n8 0.388379
R1174 VDD1.n40 VDD1.n37 0.388379
R1175 VDD1 VDD1.n28 0.209552
R1176 VDD1.n25 VDD1.n1 0.155672
R1177 VDD1.n18 VDD1.n1 0.155672
R1178 VDD1.n18 VDD1.n17 0.155672
R1179 VDD1.n17 VDD1.n5 0.155672
R1180 VDD1.n10 VDD1.n5 0.155672
R1181 VDD1.n39 VDD1.n34 0.155672
R1182 VDD1.n46 VDD1.n34 0.155672
R1183 VDD1.n47 VDD1.n46 0.155672
R1184 VDD1.n47 VDD1.n30 0.155672
R1185 VDD1.n54 VDD1.n30 0.155672
R1186 VDD1.n59 VDD1.n57 0.096016
R1187 VN.n2 VN.t5 471.065
R1188 VN.n13 VN.t3 471.065
R1189 VN.n3 VN.t4 450.084
R1190 VN.n1 VN.t2 450.084
R1191 VN.n8 VN.t8 450.084
R1192 VN.n9 VN.t6 450.084
R1193 VN.n14 VN.t1 450.084
R1194 VN.n12 VN.t0 450.084
R1195 VN.n19 VN.t9 450.084
R1196 VN.n20 VN.t7 450.084
R1197 VN.n10 VN.n9 161.3
R1198 VN.n21 VN.n20 161.3
R1199 VN.n19 VN.n11 161.3
R1200 VN.n18 VN.n17 161.3
R1201 VN.n16 VN.n15 161.3
R1202 VN.n8 VN.n0 161.3
R1203 VN.n7 VN.n6 161.3
R1204 VN.n5 VN.n4 161.3
R1205 VN.n16 VN.n13 70.4033
R1206 VN.n5 VN.n2 70.4033
R1207 VN.n9 VN.n8 48.2005
R1208 VN.n20 VN.n19 48.2005
R1209 VN.n4 VN.n3 38.7066
R1210 VN.n8 VN.n7 38.7066
R1211 VN.n15 VN.n14 38.7066
R1212 VN.n19 VN.n18 38.7066
R1213 VN VN.n21 36.26
R1214 VN.n14 VN.n13 20.9576
R1215 VN.n3 VN.n2 20.9576
R1216 VN.n4 VN.n1 9.49444
R1217 VN.n7 VN.n1 9.49444
R1218 VN.n15 VN.n12 9.49444
R1219 VN.n18 VN.n12 9.49444
R1220 VN.n21 VN.n11 0.189894
R1221 VN.n17 VN.n11 0.189894
R1222 VN.n17 VN.n16 0.189894
R1223 VN.n6 VN.n5 0.189894
R1224 VN.n6 VN.n0 0.189894
R1225 VN.n10 VN.n0 0.189894
R1226 VN VN.n10 0.0516364
R1227 VDD2.n53 VDD2.n31 289.615
R1228 VDD2.n22 VDD2.n0 289.615
R1229 VDD2.n54 VDD2.n53 185
R1230 VDD2.n52 VDD2.n51 185
R1231 VDD2.n35 VDD2.n34 185
R1232 VDD2.n46 VDD2.n45 185
R1233 VDD2.n44 VDD2.n43 185
R1234 VDD2.n39 VDD2.n38 185
R1235 VDD2.n8 VDD2.n7 185
R1236 VDD2.n13 VDD2.n12 185
R1237 VDD2.n15 VDD2.n14 185
R1238 VDD2.n4 VDD2.n3 185
R1239 VDD2.n21 VDD2.n20 185
R1240 VDD2.n23 VDD2.n22 185
R1241 VDD2.n40 VDD2.t2 147.672
R1242 VDD2.n9 VDD2.t4 147.672
R1243 VDD2.n53 VDD2.n52 104.615
R1244 VDD2.n52 VDD2.n34 104.615
R1245 VDD2.n45 VDD2.n34 104.615
R1246 VDD2.n45 VDD2.n44 104.615
R1247 VDD2.n44 VDD2.n38 104.615
R1248 VDD2.n13 VDD2.n7 104.615
R1249 VDD2.n14 VDD2.n13 104.615
R1250 VDD2.n14 VDD2.n3 104.615
R1251 VDD2.n21 VDD2.n3 104.615
R1252 VDD2.n22 VDD2.n21 104.615
R1253 VDD2.n30 VDD2.n29 68.8584
R1254 VDD2 VDD2.n61 68.8556
R1255 VDD2.n60 VDD2.n59 68.4613
R1256 VDD2.n28 VDD2.n27 68.4612
R1257 VDD2.t2 VDD2.n38 52.3082
R1258 VDD2.t4 VDD2.n7 52.3082
R1259 VDD2.n28 VDD2.n26 49.2736
R1260 VDD2.n58 VDD2.n57 48.6702
R1261 VDD2.n58 VDD2.n30 31.1248
R1262 VDD2.n40 VDD2.n39 15.6666
R1263 VDD2.n9 VDD2.n8 15.6666
R1264 VDD2.n43 VDD2.n42 12.8005
R1265 VDD2.n12 VDD2.n11 12.8005
R1266 VDD2.n46 VDD2.n37 12.0247
R1267 VDD2.n15 VDD2.n6 12.0247
R1268 VDD2.n47 VDD2.n35 11.249
R1269 VDD2.n16 VDD2.n4 11.249
R1270 VDD2.n51 VDD2.n50 10.4732
R1271 VDD2.n20 VDD2.n19 10.4732
R1272 VDD2.n54 VDD2.n33 9.69747
R1273 VDD2.n23 VDD2.n2 9.69747
R1274 VDD2.n57 VDD2.n56 9.45567
R1275 VDD2.n26 VDD2.n25 9.45567
R1276 VDD2.n56 VDD2.n55 9.3005
R1277 VDD2.n33 VDD2.n32 9.3005
R1278 VDD2.n50 VDD2.n49 9.3005
R1279 VDD2.n48 VDD2.n47 9.3005
R1280 VDD2.n37 VDD2.n36 9.3005
R1281 VDD2.n42 VDD2.n41 9.3005
R1282 VDD2.n25 VDD2.n24 9.3005
R1283 VDD2.n2 VDD2.n1 9.3005
R1284 VDD2.n19 VDD2.n18 9.3005
R1285 VDD2.n17 VDD2.n16 9.3005
R1286 VDD2.n6 VDD2.n5 9.3005
R1287 VDD2.n11 VDD2.n10 9.3005
R1288 VDD2.n55 VDD2.n31 8.92171
R1289 VDD2.n24 VDD2.n0 8.92171
R1290 VDD2.n57 VDD2.n31 5.04292
R1291 VDD2.n26 VDD2.n0 5.04292
R1292 VDD2.n41 VDD2.n40 4.38687
R1293 VDD2.n10 VDD2.n9 4.38687
R1294 VDD2.n55 VDD2.n54 4.26717
R1295 VDD2.n24 VDD2.n23 4.26717
R1296 VDD2.n61 VDD2.t8 3.75762
R1297 VDD2.n61 VDD2.t6 3.75762
R1298 VDD2.n59 VDD2.t0 3.75762
R1299 VDD2.n59 VDD2.t9 3.75762
R1300 VDD2.n29 VDD2.t1 3.75762
R1301 VDD2.n29 VDD2.t3 3.75762
R1302 VDD2.n27 VDD2.t5 3.75762
R1303 VDD2.n27 VDD2.t7 3.75762
R1304 VDD2.n51 VDD2.n33 3.49141
R1305 VDD2.n20 VDD2.n2 3.49141
R1306 VDD2.n50 VDD2.n35 2.71565
R1307 VDD2.n19 VDD2.n4 2.71565
R1308 VDD2.n47 VDD2.n46 1.93989
R1309 VDD2.n16 VDD2.n15 1.93989
R1310 VDD2.n43 VDD2.n37 1.16414
R1311 VDD2.n12 VDD2.n6 1.16414
R1312 VDD2.n60 VDD2.n58 0.603948
R1313 VDD2.n42 VDD2.n39 0.388379
R1314 VDD2.n11 VDD2.n8 0.388379
R1315 VDD2 VDD2.n60 0.209552
R1316 VDD2.n56 VDD2.n32 0.155672
R1317 VDD2.n49 VDD2.n32 0.155672
R1318 VDD2.n49 VDD2.n48 0.155672
R1319 VDD2.n48 VDD2.n36 0.155672
R1320 VDD2.n41 VDD2.n36 0.155672
R1321 VDD2.n10 VDD2.n5 0.155672
R1322 VDD2.n17 VDD2.n5 0.155672
R1323 VDD2.n18 VDD2.n17 0.155672
R1324 VDD2.n18 VDD2.n1 0.155672
R1325 VDD2.n25 VDD2.n1 0.155672
R1326 VDD2.n30 VDD2.n28 0.096016
C0 VN VDD1 0.148262f
C1 VDD2 VDD1 0.766256f
C2 VDD1 VP 2.37754f
C3 VTAIL VDD1 9.56184f
C4 VN VDD2 2.22976f
C5 VN VP 3.8675f
C6 VTAIL VN 2.21095f
C7 VDD2 VP 0.302458f
C8 VTAIL VDD2 9.59692f
C9 VTAIL VP 2.22533f
C10 VDD2 B 3.393386f
C11 VDD1 B 3.285943f
C12 VTAIL B 3.673477f
C13 VN B 7.13342f
C14 VP B 5.381966f
C15 VDD2.n0 B 0.038078f
C16 VDD2.n1 B 0.027756f
C17 VDD2.n2 B 0.014915f
C18 VDD2.n3 B 0.035254f
C19 VDD2.n4 B 0.015792f
C20 VDD2.n5 B 0.027756f
C21 VDD2.n6 B 0.014915f
C22 VDD2.n7 B 0.02644f
C23 VDD2.n8 B 0.02082f
C24 VDD2.t4 B 0.057543f
C25 VDD2.n9 B 0.113988f
C26 VDD2.n10 B 0.567133f
C27 VDD2.n11 B 0.014915f
C28 VDD2.n12 B 0.015792f
C29 VDD2.n13 B 0.035254f
C30 VDD2.n14 B 0.035254f
C31 VDD2.n15 B 0.015792f
C32 VDD2.n16 B 0.014915f
C33 VDD2.n17 B 0.027756f
C34 VDD2.n18 B 0.027756f
C35 VDD2.n19 B 0.014915f
C36 VDD2.n20 B 0.015792f
C37 VDD2.n21 B 0.035254f
C38 VDD2.n22 B 0.074662f
C39 VDD2.n23 B 0.015792f
C40 VDD2.n24 B 0.014915f
C41 VDD2.n25 B 0.063778f
C42 VDD2.n26 B 0.062076f
C43 VDD2.t5 B 0.115592f
C44 VDD2.t7 B 0.115592f
C45 VDD2.n27 B 0.948097f
C46 VDD2.n28 B 0.397538f
C47 VDD2.t1 B 0.115592f
C48 VDD2.t3 B 0.115592f
C49 VDD2.n29 B 0.949971f
C50 VDD2.n30 B 1.46859f
C51 VDD2.n31 B 0.038078f
C52 VDD2.n32 B 0.027756f
C53 VDD2.n33 B 0.014915f
C54 VDD2.n34 B 0.035254f
C55 VDD2.n35 B 0.015792f
C56 VDD2.n36 B 0.027756f
C57 VDD2.n37 B 0.014915f
C58 VDD2.n38 B 0.02644f
C59 VDD2.n39 B 0.02082f
C60 VDD2.t2 B 0.057543f
C61 VDD2.n40 B 0.113988f
C62 VDD2.n41 B 0.567133f
C63 VDD2.n42 B 0.014915f
C64 VDD2.n43 B 0.015792f
C65 VDD2.n44 B 0.035254f
C66 VDD2.n45 B 0.035254f
C67 VDD2.n46 B 0.015792f
C68 VDD2.n47 B 0.014915f
C69 VDD2.n48 B 0.027756f
C70 VDD2.n49 B 0.027756f
C71 VDD2.n50 B 0.014915f
C72 VDD2.n51 B 0.015792f
C73 VDD2.n52 B 0.035254f
C74 VDD2.n53 B 0.074662f
C75 VDD2.n54 B 0.015792f
C76 VDD2.n55 B 0.014915f
C77 VDD2.n56 B 0.063778f
C78 VDD2.n57 B 0.060763f
C79 VDD2.n58 B 1.6543f
C80 VDD2.t0 B 0.115592f
C81 VDD2.t9 B 0.115592f
C82 VDD2.n59 B 0.948102f
C83 VDD2.n60 B 0.295064f
C84 VDD2.t8 B 0.115592f
C85 VDD2.t6 B 0.115592f
C86 VDD2.n61 B 0.949947f
C87 VN.n0 B 0.051343f
C88 VN.t2 B 0.291921f
C89 VN.n1 B 0.138452f
C90 VN.t5 B 0.298426f
C91 VN.n2 B 0.139839f
C92 VN.t4 B 0.291921f
C93 VN.n3 B 0.154376f
C94 VN.n4 B 0.011651f
C95 VN.n5 B 0.159052f
C96 VN.n6 B 0.051343f
C97 VN.n7 B 0.011651f
C98 VN.t8 B 0.291921f
C99 VN.n8 B 0.154376f
C100 VN.t6 B 0.291921f
C101 VN.n9 B 0.145988f
C102 VN.n10 B 0.039789f
C103 VN.n11 B 0.051343f
C104 VN.t0 B 0.291921f
C105 VN.n12 B 0.138452f
C106 VN.t3 B 0.298426f
C107 VN.n13 B 0.139839f
C108 VN.t1 B 0.291921f
C109 VN.n14 B 0.154376f
C110 VN.n15 B 0.011651f
C111 VN.n16 B 0.159052f
C112 VN.n17 B 0.051343f
C113 VN.n18 B 0.011651f
C114 VN.t9 B 0.291921f
C115 VN.n19 B 0.154376f
C116 VN.t7 B 0.291921f
C117 VN.n20 B 0.145988f
C118 VN.n21 B 1.63808f
C119 VDD1.n0 B 0.03839f
C120 VDD1.n1 B 0.027984f
C121 VDD1.n2 B 0.015037f
C122 VDD1.n3 B 0.035542f
C123 VDD1.n4 B 0.015922f
C124 VDD1.n5 B 0.027984f
C125 VDD1.n6 B 0.015037f
C126 VDD1.n7 B 0.026657f
C127 VDD1.n8 B 0.020991f
C128 VDD1.t2 B 0.058015f
C129 VDD1.n9 B 0.114921f
C130 VDD1.n10 B 0.571778f
C131 VDD1.n11 B 0.015037f
C132 VDD1.n12 B 0.015922f
C133 VDD1.n13 B 0.035542f
C134 VDD1.n14 B 0.035542f
C135 VDD1.n15 B 0.015922f
C136 VDD1.n16 B 0.015037f
C137 VDD1.n17 B 0.027984f
C138 VDD1.n18 B 0.027984f
C139 VDD1.n19 B 0.015037f
C140 VDD1.n20 B 0.015922f
C141 VDD1.n21 B 0.035542f
C142 VDD1.n22 B 0.075274f
C143 VDD1.n23 B 0.015922f
C144 VDD1.n24 B 0.015037f
C145 VDD1.n25 B 0.064301f
C146 VDD1.n26 B 0.062584f
C147 VDD1.t5 B 0.116538f
C148 VDD1.t8 B 0.116538f
C149 VDD1.n27 B 0.955867f
C150 VDD1.n28 B 0.404235f
C151 VDD1.n29 B 0.03839f
C152 VDD1.n30 B 0.027984f
C153 VDD1.n31 B 0.015037f
C154 VDD1.n32 B 0.035542f
C155 VDD1.n33 B 0.015922f
C156 VDD1.n34 B 0.027984f
C157 VDD1.n35 B 0.015037f
C158 VDD1.n36 B 0.026657f
C159 VDD1.n37 B 0.020991f
C160 VDD1.t4 B 0.058015f
C161 VDD1.n38 B 0.114921f
C162 VDD1.n39 B 0.571778f
C163 VDD1.n40 B 0.015037f
C164 VDD1.n41 B 0.015922f
C165 VDD1.n42 B 0.035542f
C166 VDD1.n43 B 0.035542f
C167 VDD1.n44 B 0.015922f
C168 VDD1.n45 B 0.015037f
C169 VDD1.n46 B 0.027984f
C170 VDD1.n47 B 0.027984f
C171 VDD1.n48 B 0.015037f
C172 VDD1.n49 B 0.015922f
C173 VDD1.n50 B 0.035542f
C174 VDD1.n51 B 0.075274f
C175 VDD1.n52 B 0.015922f
C176 VDD1.n53 B 0.015037f
C177 VDD1.n54 B 0.064301f
C178 VDD1.n55 B 0.062584f
C179 VDD1.t7 B 0.116538f
C180 VDD1.t6 B 0.116538f
C181 VDD1.n56 B 0.955862f
C182 VDD1.n57 B 0.400794f
C183 VDD1.t1 B 0.116538f
C184 VDD1.t9 B 0.116538f
C185 VDD1.n58 B 0.957751f
C186 VDD1.n59 B 1.55607f
C187 VDD1.t0 B 0.116538f
C188 VDD1.t3 B 0.116538f
C189 VDD1.n60 B 0.955863f
C190 VDD1.n61 B 1.91315f
C191 VTAIL.t19 B 0.12807f
C192 VTAIL.t18 B 0.12807f
C193 VTAIL.n0 B 0.972966f
C194 VTAIL.n1 B 0.409161f
C195 VTAIL.n2 B 0.042188f
C196 VTAIL.n3 B 0.030753f
C197 VTAIL.n4 B 0.016525f
C198 VTAIL.n5 B 0.03906f
C199 VTAIL.n6 B 0.017497f
C200 VTAIL.n7 B 0.030753f
C201 VTAIL.n8 B 0.016525f
C202 VTAIL.n9 B 0.029295f
C203 VTAIL.n10 B 0.023068f
C204 VTAIL.t15 B 0.063755f
C205 VTAIL.n11 B 0.126293f
C206 VTAIL.n12 B 0.628357f
C207 VTAIL.n13 B 0.016525f
C208 VTAIL.n14 B 0.017497f
C209 VTAIL.n15 B 0.03906f
C210 VTAIL.n16 B 0.03906f
C211 VTAIL.n17 B 0.017497f
C212 VTAIL.n18 B 0.016525f
C213 VTAIL.n19 B 0.030753f
C214 VTAIL.n20 B 0.030753f
C215 VTAIL.n21 B 0.016525f
C216 VTAIL.n22 B 0.017497f
C217 VTAIL.n23 B 0.03906f
C218 VTAIL.n24 B 0.082723f
C219 VTAIL.n25 B 0.017497f
C220 VTAIL.n26 B 0.016525f
C221 VTAIL.n27 B 0.070663f
C222 VTAIL.n28 B 0.046085f
C223 VTAIL.n29 B 0.16228f
C224 VTAIL.t12 B 0.12807f
C225 VTAIL.t9 B 0.12807f
C226 VTAIL.n30 B 0.972966f
C227 VTAIL.n31 B 0.401686f
C228 VTAIL.t10 B 0.12807f
C229 VTAIL.t11 B 0.12807f
C230 VTAIL.n32 B 0.972966f
C231 VTAIL.n33 B 1.32941f
C232 VTAIL.t3 B 0.12807f
C233 VTAIL.t2 B 0.12807f
C234 VTAIL.n34 B 0.972973f
C235 VTAIL.n35 B 1.3294f
C236 VTAIL.t0 B 0.12807f
C237 VTAIL.t1 B 0.12807f
C238 VTAIL.n36 B 0.972973f
C239 VTAIL.n37 B 0.401679f
C240 VTAIL.n38 B 0.042188f
C241 VTAIL.n39 B 0.030753f
C242 VTAIL.n40 B 0.016525f
C243 VTAIL.n41 B 0.03906f
C244 VTAIL.n42 B 0.017497f
C245 VTAIL.n43 B 0.030753f
C246 VTAIL.n44 B 0.016525f
C247 VTAIL.n45 B 0.029295f
C248 VTAIL.n46 B 0.023068f
C249 VTAIL.t17 B 0.063755f
C250 VTAIL.n47 B 0.126293f
C251 VTAIL.n48 B 0.628357f
C252 VTAIL.n49 B 0.016525f
C253 VTAIL.n50 B 0.017497f
C254 VTAIL.n51 B 0.03906f
C255 VTAIL.n52 B 0.03906f
C256 VTAIL.n53 B 0.017497f
C257 VTAIL.n54 B 0.016525f
C258 VTAIL.n55 B 0.030753f
C259 VTAIL.n56 B 0.030753f
C260 VTAIL.n57 B 0.016525f
C261 VTAIL.n58 B 0.017497f
C262 VTAIL.n59 B 0.03906f
C263 VTAIL.n60 B 0.082723f
C264 VTAIL.n61 B 0.017497f
C265 VTAIL.n62 B 0.016525f
C266 VTAIL.n63 B 0.070663f
C267 VTAIL.n64 B 0.046085f
C268 VTAIL.n65 B 0.16228f
C269 VTAIL.t7 B 0.12807f
C270 VTAIL.t13 B 0.12807f
C271 VTAIL.n66 B 0.972973f
C272 VTAIL.n67 B 0.418337f
C273 VTAIL.t14 B 0.12807f
C274 VTAIL.t16 B 0.12807f
C275 VTAIL.n68 B 0.972973f
C276 VTAIL.n69 B 0.401679f
C277 VTAIL.n70 B 0.042188f
C278 VTAIL.n71 B 0.030753f
C279 VTAIL.n72 B 0.016525f
C280 VTAIL.n73 B 0.03906f
C281 VTAIL.n74 B 0.017497f
C282 VTAIL.n75 B 0.030753f
C283 VTAIL.n76 B 0.016525f
C284 VTAIL.n77 B 0.029295f
C285 VTAIL.n78 B 0.023068f
C286 VTAIL.t8 B 0.063755f
C287 VTAIL.n79 B 0.126293f
C288 VTAIL.n80 B 0.628357f
C289 VTAIL.n81 B 0.016525f
C290 VTAIL.n82 B 0.017497f
C291 VTAIL.n83 B 0.03906f
C292 VTAIL.n84 B 0.03906f
C293 VTAIL.n85 B 0.017497f
C294 VTAIL.n86 B 0.016525f
C295 VTAIL.n87 B 0.030753f
C296 VTAIL.n88 B 0.030753f
C297 VTAIL.n89 B 0.016525f
C298 VTAIL.n90 B 0.017497f
C299 VTAIL.n91 B 0.03906f
C300 VTAIL.n92 B 0.082723f
C301 VTAIL.n93 B 0.017497f
C302 VTAIL.n94 B 0.016525f
C303 VTAIL.n95 B 0.070663f
C304 VTAIL.n96 B 0.046085f
C305 VTAIL.n97 B 1.01355f
C306 VTAIL.n98 B 0.042188f
C307 VTAIL.n99 B 0.030753f
C308 VTAIL.n100 B 0.016525f
C309 VTAIL.n101 B 0.03906f
C310 VTAIL.n102 B 0.017497f
C311 VTAIL.n103 B 0.030753f
C312 VTAIL.n104 B 0.016525f
C313 VTAIL.n105 B 0.029295f
C314 VTAIL.n106 B 0.023068f
C315 VTAIL.t4 B 0.063755f
C316 VTAIL.n107 B 0.126293f
C317 VTAIL.n108 B 0.628357f
C318 VTAIL.n109 B 0.016525f
C319 VTAIL.n110 B 0.017497f
C320 VTAIL.n111 B 0.03906f
C321 VTAIL.n112 B 0.03906f
C322 VTAIL.n113 B 0.017497f
C323 VTAIL.n114 B 0.016525f
C324 VTAIL.n115 B 0.030753f
C325 VTAIL.n116 B 0.030753f
C326 VTAIL.n117 B 0.016525f
C327 VTAIL.n118 B 0.017497f
C328 VTAIL.n119 B 0.03906f
C329 VTAIL.n120 B 0.082723f
C330 VTAIL.n121 B 0.017497f
C331 VTAIL.n122 B 0.016525f
C332 VTAIL.n123 B 0.070663f
C333 VTAIL.n124 B 0.046085f
C334 VTAIL.n125 B 1.01355f
C335 VTAIL.t5 B 0.12807f
C336 VTAIL.t6 B 0.12807f
C337 VTAIL.n126 B 0.972966f
C338 VTAIL.n127 B 0.351072f
C339 VP.n0 B 0.053041f
C340 VP.t3 B 0.301577f
C341 VP.n1 B 0.143032f
C342 VP.n2 B 0.053041f
C343 VP.n3 B 0.053041f
C344 VP.t6 B 0.301577f
C345 VP.t9 B 0.301577f
C346 VP.t1 B 0.301577f
C347 VP.n4 B 0.143032f
C348 VP.t7 B 0.308298f
C349 VP.n5 B 0.144465f
C350 VP.t4 B 0.301577f
C351 VP.n6 B 0.159483f
C352 VP.n7 B 0.012036f
C353 VP.n8 B 0.164313f
C354 VP.n9 B 0.053041f
C355 VP.n10 B 0.012036f
C356 VP.n11 B 0.159483f
C357 VP.n12 B 0.150817f
C358 VP.n13 B 1.65707f
C359 VP.n14 B 1.71022f
C360 VP.t5 B 0.301577f
C361 VP.n15 B 0.150817f
C362 VP.t2 B 0.301577f
C363 VP.n16 B 0.159483f
C364 VP.n17 B 0.012036f
C365 VP.n18 B 0.053041f
C366 VP.n19 B 0.053041f
C367 VP.n20 B 0.012036f
C368 VP.t8 B 0.301577f
C369 VP.n21 B 0.159483f
C370 VP.t0 B 0.301577f
C371 VP.n22 B 0.150817f
C372 VP.n23 B 0.041105f
.ends

