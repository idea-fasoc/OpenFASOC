* NGSPICE file created from diff_pair_sample_1493.ext - technology: sky130A

.subckt diff_pair_sample_1493 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t19 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=3.12015 pd=19.24 as=3.12015 ps=19.24 w=18.91 l=0.2
X1 VTAIL.t2 VP.t0 VDD1.t9 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=3.12015 pd=19.24 as=3.12015 ps=19.24 w=18.91 l=0.2
X2 VDD2.t8 VN.t1 VTAIL.t16 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=7.3749 pd=38.6 as=3.12015 ps=19.24 w=18.91 l=0.2
X3 VTAIL.t17 VN.t2 VDD2.t7 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=3.12015 pd=19.24 as=3.12015 ps=19.24 w=18.91 l=0.2
X4 VTAIL.t11 VN.t3 VDD2.t6 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=3.12015 pd=19.24 as=3.12015 ps=19.24 w=18.91 l=0.2
X5 VTAIL.t12 VN.t4 VDD2.t5 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=3.12015 pd=19.24 as=3.12015 ps=19.24 w=18.91 l=0.2
X6 VDD1.t8 VP.t1 VTAIL.t7 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=7.3749 pd=38.6 as=3.12015 ps=19.24 w=18.91 l=0.2
X7 VDD2.t4 VN.t5 VTAIL.t10 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=3.12015 pd=19.24 as=7.3749 ps=38.6 w=18.91 l=0.2
X8 B.t11 B.t9 B.t10 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=7.3749 pd=38.6 as=0 ps=0 w=18.91 l=0.2
X9 VDD2.t3 VN.t6 VTAIL.t18 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=3.12015 pd=19.24 as=7.3749 ps=38.6 w=18.91 l=0.2
X10 VDD2.t2 VN.t7 VTAIL.t15 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=7.3749 pd=38.6 as=3.12015 ps=19.24 w=18.91 l=0.2
X11 B.t8 B.t6 B.t7 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=7.3749 pd=38.6 as=0 ps=0 w=18.91 l=0.2
X12 VDD1.t7 VP.t2 VTAIL.t9 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=3.12015 pd=19.24 as=7.3749 ps=38.6 w=18.91 l=0.2
X13 VTAIL.t6 VP.t3 VDD1.t6 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=3.12015 pd=19.24 as=3.12015 ps=19.24 w=18.91 l=0.2
X14 VTAIL.t0 VP.t4 VDD1.t5 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=3.12015 pd=19.24 as=3.12015 ps=19.24 w=18.91 l=0.2
X15 VTAIL.t14 VN.t8 VDD2.t1 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=3.12015 pd=19.24 as=3.12015 ps=19.24 w=18.91 l=0.2
X16 B.t5 B.t3 B.t4 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=7.3749 pd=38.6 as=0 ps=0 w=18.91 l=0.2
X17 VDD1.t4 VP.t5 VTAIL.t8 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=7.3749 pd=38.6 as=3.12015 ps=19.24 w=18.91 l=0.2
X18 VDD1.t3 VP.t6 VTAIL.t1 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=3.12015 pd=19.24 as=7.3749 ps=38.6 w=18.91 l=0.2
X19 VDD1.t2 VP.t7 VTAIL.t4 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=3.12015 pd=19.24 as=3.12015 ps=19.24 w=18.91 l=0.2
X20 VDD1.t1 VP.t8 VTAIL.t5 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=3.12015 pd=19.24 as=3.12015 ps=19.24 w=18.91 l=0.2
X21 B.t2 B.t0 B.t1 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=7.3749 pd=38.6 as=0 ps=0 w=18.91 l=0.2
X22 VTAIL.t3 VP.t9 VDD1.t0 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=3.12015 pd=19.24 as=3.12015 ps=19.24 w=18.91 l=0.2
X23 VDD2.t0 VN.t9 VTAIL.t13 w_n1606_n4750# sky130_fd_pr__pfet_01v8 ad=3.12015 pd=19.24 as=3.12015 ps=19.24 w=18.91 l=0.2
R0 VN.n8 VN.t5 2481.79
R1 VN.n2 VN.t1 2481.79
R2 VN.n18 VN.t7 2481.79
R3 VN.n12 VN.t6 2481.79
R4 VN.n7 VN.t2 2436.51
R5 VN.n5 VN.t0 2436.51
R6 VN.n1 VN.t3 2436.51
R7 VN.n17 VN.t8 2436.51
R8 VN.n15 VN.t9 2436.51
R9 VN.n11 VN.t4 2436.51
R10 VN.n13 VN.n12 161.489
R11 VN.n3 VN.n2 161.489
R12 VN.n9 VN.n8 161.3
R13 VN.n19 VN.n18 161.3
R14 VN.n16 VN.n10 161.3
R15 VN.n14 VN.n13 161.3
R16 VN.n6 VN.n0 161.3
R17 VN.n4 VN.n3 161.3
R18 VN VN.n19 45.7486
R19 VN.n4 VN.n1 40.8975
R20 VN.n7 VN.n6 40.8975
R21 VN.n17 VN.n16 40.8975
R22 VN.n14 VN.n11 40.8975
R23 VN.n5 VN.n4 36.5157
R24 VN.n6 VN.n5 36.5157
R25 VN.n16 VN.n15 36.5157
R26 VN.n15 VN.n14 36.5157
R27 VN.n2 VN.n1 32.1338
R28 VN.n8 VN.n7 32.1338
R29 VN.n18 VN.n17 32.1338
R30 VN.n12 VN.n11 32.1338
R31 VN.n19 VN.n10 0.189894
R32 VN.n13 VN.n10 0.189894
R33 VN.n3 VN.n0 0.189894
R34 VN.n9 VN.n0 0.189894
R35 VN VN.n9 0.0516364
R36 VTAIL.n432 VTAIL.n332 756.745
R37 VTAIL.n102 VTAIL.n2 756.745
R38 VTAIL.n326 VTAIL.n226 756.745
R39 VTAIL.n216 VTAIL.n116 756.745
R40 VTAIL.n367 VTAIL.n366 585
R41 VTAIL.n364 VTAIL.n363 585
R42 VTAIL.n373 VTAIL.n372 585
R43 VTAIL.n375 VTAIL.n374 585
R44 VTAIL.n360 VTAIL.n359 585
R45 VTAIL.n381 VTAIL.n380 585
R46 VTAIL.n383 VTAIL.n382 585
R47 VTAIL.n356 VTAIL.n355 585
R48 VTAIL.n389 VTAIL.n388 585
R49 VTAIL.n391 VTAIL.n390 585
R50 VTAIL.n352 VTAIL.n351 585
R51 VTAIL.n397 VTAIL.n396 585
R52 VTAIL.n399 VTAIL.n398 585
R53 VTAIL.n348 VTAIL.n347 585
R54 VTAIL.n405 VTAIL.n404 585
R55 VTAIL.n408 VTAIL.n407 585
R56 VTAIL.n406 VTAIL.n344 585
R57 VTAIL.n413 VTAIL.n343 585
R58 VTAIL.n415 VTAIL.n414 585
R59 VTAIL.n417 VTAIL.n416 585
R60 VTAIL.n340 VTAIL.n339 585
R61 VTAIL.n423 VTAIL.n422 585
R62 VTAIL.n425 VTAIL.n424 585
R63 VTAIL.n336 VTAIL.n335 585
R64 VTAIL.n431 VTAIL.n430 585
R65 VTAIL.n433 VTAIL.n432 585
R66 VTAIL.n37 VTAIL.n36 585
R67 VTAIL.n34 VTAIL.n33 585
R68 VTAIL.n43 VTAIL.n42 585
R69 VTAIL.n45 VTAIL.n44 585
R70 VTAIL.n30 VTAIL.n29 585
R71 VTAIL.n51 VTAIL.n50 585
R72 VTAIL.n53 VTAIL.n52 585
R73 VTAIL.n26 VTAIL.n25 585
R74 VTAIL.n59 VTAIL.n58 585
R75 VTAIL.n61 VTAIL.n60 585
R76 VTAIL.n22 VTAIL.n21 585
R77 VTAIL.n67 VTAIL.n66 585
R78 VTAIL.n69 VTAIL.n68 585
R79 VTAIL.n18 VTAIL.n17 585
R80 VTAIL.n75 VTAIL.n74 585
R81 VTAIL.n78 VTAIL.n77 585
R82 VTAIL.n76 VTAIL.n14 585
R83 VTAIL.n83 VTAIL.n13 585
R84 VTAIL.n85 VTAIL.n84 585
R85 VTAIL.n87 VTAIL.n86 585
R86 VTAIL.n10 VTAIL.n9 585
R87 VTAIL.n93 VTAIL.n92 585
R88 VTAIL.n95 VTAIL.n94 585
R89 VTAIL.n6 VTAIL.n5 585
R90 VTAIL.n101 VTAIL.n100 585
R91 VTAIL.n103 VTAIL.n102 585
R92 VTAIL.n327 VTAIL.n326 585
R93 VTAIL.n325 VTAIL.n324 585
R94 VTAIL.n230 VTAIL.n229 585
R95 VTAIL.n319 VTAIL.n318 585
R96 VTAIL.n317 VTAIL.n316 585
R97 VTAIL.n234 VTAIL.n233 585
R98 VTAIL.n311 VTAIL.n310 585
R99 VTAIL.n309 VTAIL.n308 585
R100 VTAIL.n307 VTAIL.n237 585
R101 VTAIL.n241 VTAIL.n238 585
R102 VTAIL.n302 VTAIL.n301 585
R103 VTAIL.n300 VTAIL.n299 585
R104 VTAIL.n243 VTAIL.n242 585
R105 VTAIL.n294 VTAIL.n293 585
R106 VTAIL.n292 VTAIL.n291 585
R107 VTAIL.n247 VTAIL.n246 585
R108 VTAIL.n286 VTAIL.n285 585
R109 VTAIL.n284 VTAIL.n283 585
R110 VTAIL.n251 VTAIL.n250 585
R111 VTAIL.n278 VTAIL.n277 585
R112 VTAIL.n276 VTAIL.n275 585
R113 VTAIL.n255 VTAIL.n254 585
R114 VTAIL.n270 VTAIL.n269 585
R115 VTAIL.n268 VTAIL.n267 585
R116 VTAIL.n259 VTAIL.n258 585
R117 VTAIL.n262 VTAIL.n261 585
R118 VTAIL.n217 VTAIL.n216 585
R119 VTAIL.n215 VTAIL.n214 585
R120 VTAIL.n120 VTAIL.n119 585
R121 VTAIL.n209 VTAIL.n208 585
R122 VTAIL.n207 VTAIL.n206 585
R123 VTAIL.n124 VTAIL.n123 585
R124 VTAIL.n201 VTAIL.n200 585
R125 VTAIL.n199 VTAIL.n198 585
R126 VTAIL.n197 VTAIL.n127 585
R127 VTAIL.n131 VTAIL.n128 585
R128 VTAIL.n192 VTAIL.n191 585
R129 VTAIL.n190 VTAIL.n189 585
R130 VTAIL.n133 VTAIL.n132 585
R131 VTAIL.n184 VTAIL.n183 585
R132 VTAIL.n182 VTAIL.n181 585
R133 VTAIL.n137 VTAIL.n136 585
R134 VTAIL.n176 VTAIL.n175 585
R135 VTAIL.n174 VTAIL.n173 585
R136 VTAIL.n141 VTAIL.n140 585
R137 VTAIL.n168 VTAIL.n167 585
R138 VTAIL.n166 VTAIL.n165 585
R139 VTAIL.n145 VTAIL.n144 585
R140 VTAIL.n160 VTAIL.n159 585
R141 VTAIL.n158 VTAIL.n157 585
R142 VTAIL.n149 VTAIL.n148 585
R143 VTAIL.n152 VTAIL.n151 585
R144 VTAIL.t9 VTAIL.n260 327.466
R145 VTAIL.t18 VTAIL.n150 327.466
R146 VTAIL.t10 VTAIL.n365 327.466
R147 VTAIL.t1 VTAIL.n35 327.466
R148 VTAIL.n366 VTAIL.n363 171.744
R149 VTAIL.n373 VTAIL.n363 171.744
R150 VTAIL.n374 VTAIL.n373 171.744
R151 VTAIL.n374 VTAIL.n359 171.744
R152 VTAIL.n381 VTAIL.n359 171.744
R153 VTAIL.n382 VTAIL.n381 171.744
R154 VTAIL.n382 VTAIL.n355 171.744
R155 VTAIL.n389 VTAIL.n355 171.744
R156 VTAIL.n390 VTAIL.n389 171.744
R157 VTAIL.n390 VTAIL.n351 171.744
R158 VTAIL.n397 VTAIL.n351 171.744
R159 VTAIL.n398 VTAIL.n397 171.744
R160 VTAIL.n398 VTAIL.n347 171.744
R161 VTAIL.n405 VTAIL.n347 171.744
R162 VTAIL.n407 VTAIL.n405 171.744
R163 VTAIL.n407 VTAIL.n406 171.744
R164 VTAIL.n406 VTAIL.n343 171.744
R165 VTAIL.n415 VTAIL.n343 171.744
R166 VTAIL.n416 VTAIL.n415 171.744
R167 VTAIL.n416 VTAIL.n339 171.744
R168 VTAIL.n423 VTAIL.n339 171.744
R169 VTAIL.n424 VTAIL.n423 171.744
R170 VTAIL.n424 VTAIL.n335 171.744
R171 VTAIL.n431 VTAIL.n335 171.744
R172 VTAIL.n432 VTAIL.n431 171.744
R173 VTAIL.n36 VTAIL.n33 171.744
R174 VTAIL.n43 VTAIL.n33 171.744
R175 VTAIL.n44 VTAIL.n43 171.744
R176 VTAIL.n44 VTAIL.n29 171.744
R177 VTAIL.n51 VTAIL.n29 171.744
R178 VTAIL.n52 VTAIL.n51 171.744
R179 VTAIL.n52 VTAIL.n25 171.744
R180 VTAIL.n59 VTAIL.n25 171.744
R181 VTAIL.n60 VTAIL.n59 171.744
R182 VTAIL.n60 VTAIL.n21 171.744
R183 VTAIL.n67 VTAIL.n21 171.744
R184 VTAIL.n68 VTAIL.n67 171.744
R185 VTAIL.n68 VTAIL.n17 171.744
R186 VTAIL.n75 VTAIL.n17 171.744
R187 VTAIL.n77 VTAIL.n75 171.744
R188 VTAIL.n77 VTAIL.n76 171.744
R189 VTAIL.n76 VTAIL.n13 171.744
R190 VTAIL.n85 VTAIL.n13 171.744
R191 VTAIL.n86 VTAIL.n85 171.744
R192 VTAIL.n86 VTAIL.n9 171.744
R193 VTAIL.n93 VTAIL.n9 171.744
R194 VTAIL.n94 VTAIL.n93 171.744
R195 VTAIL.n94 VTAIL.n5 171.744
R196 VTAIL.n101 VTAIL.n5 171.744
R197 VTAIL.n102 VTAIL.n101 171.744
R198 VTAIL.n326 VTAIL.n325 171.744
R199 VTAIL.n325 VTAIL.n229 171.744
R200 VTAIL.n318 VTAIL.n229 171.744
R201 VTAIL.n318 VTAIL.n317 171.744
R202 VTAIL.n317 VTAIL.n233 171.744
R203 VTAIL.n310 VTAIL.n233 171.744
R204 VTAIL.n310 VTAIL.n309 171.744
R205 VTAIL.n309 VTAIL.n237 171.744
R206 VTAIL.n241 VTAIL.n237 171.744
R207 VTAIL.n301 VTAIL.n241 171.744
R208 VTAIL.n301 VTAIL.n300 171.744
R209 VTAIL.n300 VTAIL.n242 171.744
R210 VTAIL.n293 VTAIL.n242 171.744
R211 VTAIL.n293 VTAIL.n292 171.744
R212 VTAIL.n292 VTAIL.n246 171.744
R213 VTAIL.n285 VTAIL.n246 171.744
R214 VTAIL.n285 VTAIL.n284 171.744
R215 VTAIL.n284 VTAIL.n250 171.744
R216 VTAIL.n277 VTAIL.n250 171.744
R217 VTAIL.n277 VTAIL.n276 171.744
R218 VTAIL.n276 VTAIL.n254 171.744
R219 VTAIL.n269 VTAIL.n254 171.744
R220 VTAIL.n269 VTAIL.n268 171.744
R221 VTAIL.n268 VTAIL.n258 171.744
R222 VTAIL.n261 VTAIL.n258 171.744
R223 VTAIL.n216 VTAIL.n215 171.744
R224 VTAIL.n215 VTAIL.n119 171.744
R225 VTAIL.n208 VTAIL.n119 171.744
R226 VTAIL.n208 VTAIL.n207 171.744
R227 VTAIL.n207 VTAIL.n123 171.744
R228 VTAIL.n200 VTAIL.n123 171.744
R229 VTAIL.n200 VTAIL.n199 171.744
R230 VTAIL.n199 VTAIL.n127 171.744
R231 VTAIL.n131 VTAIL.n127 171.744
R232 VTAIL.n191 VTAIL.n131 171.744
R233 VTAIL.n191 VTAIL.n190 171.744
R234 VTAIL.n190 VTAIL.n132 171.744
R235 VTAIL.n183 VTAIL.n132 171.744
R236 VTAIL.n183 VTAIL.n182 171.744
R237 VTAIL.n182 VTAIL.n136 171.744
R238 VTAIL.n175 VTAIL.n136 171.744
R239 VTAIL.n175 VTAIL.n174 171.744
R240 VTAIL.n174 VTAIL.n140 171.744
R241 VTAIL.n167 VTAIL.n140 171.744
R242 VTAIL.n167 VTAIL.n166 171.744
R243 VTAIL.n166 VTAIL.n144 171.744
R244 VTAIL.n159 VTAIL.n144 171.744
R245 VTAIL.n159 VTAIL.n158 171.744
R246 VTAIL.n158 VTAIL.n148 171.744
R247 VTAIL.n151 VTAIL.n148 171.744
R248 VTAIL.n366 VTAIL.t10 85.8723
R249 VTAIL.n36 VTAIL.t1 85.8723
R250 VTAIL.n261 VTAIL.t9 85.8723
R251 VTAIL.n151 VTAIL.t18 85.8723
R252 VTAIL.n439 VTAIL.n438 50.7364
R253 VTAIL.n1 VTAIL.n0 50.7364
R254 VTAIL.n109 VTAIL.n108 50.7364
R255 VTAIL.n111 VTAIL.n110 50.7364
R256 VTAIL.n225 VTAIL.n224 50.7364
R257 VTAIL.n223 VTAIL.n222 50.7364
R258 VTAIL.n115 VTAIL.n114 50.7364
R259 VTAIL.n113 VTAIL.n112 50.7364
R260 VTAIL.n437 VTAIL.n436 31.2157
R261 VTAIL.n107 VTAIL.n106 31.2157
R262 VTAIL.n331 VTAIL.n330 31.2157
R263 VTAIL.n221 VTAIL.n220 31.2157
R264 VTAIL.n113 VTAIL.n111 29.5824
R265 VTAIL.n437 VTAIL.n331 29.1255
R266 VTAIL.n367 VTAIL.n365 16.3895
R267 VTAIL.n37 VTAIL.n35 16.3895
R268 VTAIL.n262 VTAIL.n260 16.3895
R269 VTAIL.n152 VTAIL.n150 16.3895
R270 VTAIL.n414 VTAIL.n413 13.1884
R271 VTAIL.n84 VTAIL.n83 13.1884
R272 VTAIL.n308 VTAIL.n307 13.1884
R273 VTAIL.n198 VTAIL.n197 13.1884
R274 VTAIL.n368 VTAIL.n364 12.8005
R275 VTAIL.n412 VTAIL.n344 12.8005
R276 VTAIL.n417 VTAIL.n342 12.8005
R277 VTAIL.n38 VTAIL.n34 12.8005
R278 VTAIL.n82 VTAIL.n14 12.8005
R279 VTAIL.n87 VTAIL.n12 12.8005
R280 VTAIL.n311 VTAIL.n236 12.8005
R281 VTAIL.n306 VTAIL.n238 12.8005
R282 VTAIL.n263 VTAIL.n259 12.8005
R283 VTAIL.n201 VTAIL.n126 12.8005
R284 VTAIL.n196 VTAIL.n128 12.8005
R285 VTAIL.n153 VTAIL.n149 12.8005
R286 VTAIL.n372 VTAIL.n371 12.0247
R287 VTAIL.n409 VTAIL.n408 12.0247
R288 VTAIL.n418 VTAIL.n340 12.0247
R289 VTAIL.n42 VTAIL.n41 12.0247
R290 VTAIL.n79 VTAIL.n78 12.0247
R291 VTAIL.n88 VTAIL.n10 12.0247
R292 VTAIL.n312 VTAIL.n234 12.0247
R293 VTAIL.n303 VTAIL.n302 12.0247
R294 VTAIL.n267 VTAIL.n266 12.0247
R295 VTAIL.n202 VTAIL.n124 12.0247
R296 VTAIL.n193 VTAIL.n192 12.0247
R297 VTAIL.n157 VTAIL.n156 12.0247
R298 VTAIL.n375 VTAIL.n362 11.249
R299 VTAIL.n404 VTAIL.n346 11.249
R300 VTAIL.n422 VTAIL.n421 11.249
R301 VTAIL.n45 VTAIL.n32 11.249
R302 VTAIL.n74 VTAIL.n16 11.249
R303 VTAIL.n92 VTAIL.n91 11.249
R304 VTAIL.n316 VTAIL.n315 11.249
R305 VTAIL.n299 VTAIL.n240 11.249
R306 VTAIL.n270 VTAIL.n257 11.249
R307 VTAIL.n206 VTAIL.n205 11.249
R308 VTAIL.n189 VTAIL.n130 11.249
R309 VTAIL.n160 VTAIL.n147 11.249
R310 VTAIL.n376 VTAIL.n360 10.4732
R311 VTAIL.n403 VTAIL.n348 10.4732
R312 VTAIL.n425 VTAIL.n338 10.4732
R313 VTAIL.n46 VTAIL.n30 10.4732
R314 VTAIL.n73 VTAIL.n18 10.4732
R315 VTAIL.n95 VTAIL.n8 10.4732
R316 VTAIL.n319 VTAIL.n232 10.4732
R317 VTAIL.n298 VTAIL.n243 10.4732
R318 VTAIL.n271 VTAIL.n255 10.4732
R319 VTAIL.n209 VTAIL.n122 10.4732
R320 VTAIL.n188 VTAIL.n133 10.4732
R321 VTAIL.n161 VTAIL.n145 10.4732
R322 VTAIL.n380 VTAIL.n379 9.69747
R323 VTAIL.n400 VTAIL.n399 9.69747
R324 VTAIL.n426 VTAIL.n336 9.69747
R325 VTAIL.n50 VTAIL.n49 9.69747
R326 VTAIL.n70 VTAIL.n69 9.69747
R327 VTAIL.n96 VTAIL.n6 9.69747
R328 VTAIL.n320 VTAIL.n230 9.69747
R329 VTAIL.n295 VTAIL.n294 9.69747
R330 VTAIL.n275 VTAIL.n274 9.69747
R331 VTAIL.n210 VTAIL.n120 9.69747
R332 VTAIL.n185 VTAIL.n184 9.69747
R333 VTAIL.n165 VTAIL.n164 9.69747
R334 VTAIL.n436 VTAIL.n435 9.45567
R335 VTAIL.n106 VTAIL.n105 9.45567
R336 VTAIL.n330 VTAIL.n329 9.45567
R337 VTAIL.n220 VTAIL.n219 9.45567
R338 VTAIL.n334 VTAIL.n333 9.3005
R339 VTAIL.n429 VTAIL.n428 9.3005
R340 VTAIL.n427 VTAIL.n426 9.3005
R341 VTAIL.n338 VTAIL.n337 9.3005
R342 VTAIL.n421 VTAIL.n420 9.3005
R343 VTAIL.n419 VTAIL.n418 9.3005
R344 VTAIL.n342 VTAIL.n341 9.3005
R345 VTAIL.n387 VTAIL.n386 9.3005
R346 VTAIL.n385 VTAIL.n384 9.3005
R347 VTAIL.n358 VTAIL.n357 9.3005
R348 VTAIL.n379 VTAIL.n378 9.3005
R349 VTAIL.n377 VTAIL.n376 9.3005
R350 VTAIL.n362 VTAIL.n361 9.3005
R351 VTAIL.n371 VTAIL.n370 9.3005
R352 VTAIL.n369 VTAIL.n368 9.3005
R353 VTAIL.n354 VTAIL.n353 9.3005
R354 VTAIL.n393 VTAIL.n392 9.3005
R355 VTAIL.n395 VTAIL.n394 9.3005
R356 VTAIL.n350 VTAIL.n349 9.3005
R357 VTAIL.n401 VTAIL.n400 9.3005
R358 VTAIL.n403 VTAIL.n402 9.3005
R359 VTAIL.n346 VTAIL.n345 9.3005
R360 VTAIL.n410 VTAIL.n409 9.3005
R361 VTAIL.n412 VTAIL.n411 9.3005
R362 VTAIL.n435 VTAIL.n434 9.3005
R363 VTAIL.n4 VTAIL.n3 9.3005
R364 VTAIL.n99 VTAIL.n98 9.3005
R365 VTAIL.n97 VTAIL.n96 9.3005
R366 VTAIL.n8 VTAIL.n7 9.3005
R367 VTAIL.n91 VTAIL.n90 9.3005
R368 VTAIL.n89 VTAIL.n88 9.3005
R369 VTAIL.n12 VTAIL.n11 9.3005
R370 VTAIL.n57 VTAIL.n56 9.3005
R371 VTAIL.n55 VTAIL.n54 9.3005
R372 VTAIL.n28 VTAIL.n27 9.3005
R373 VTAIL.n49 VTAIL.n48 9.3005
R374 VTAIL.n47 VTAIL.n46 9.3005
R375 VTAIL.n32 VTAIL.n31 9.3005
R376 VTAIL.n41 VTAIL.n40 9.3005
R377 VTAIL.n39 VTAIL.n38 9.3005
R378 VTAIL.n24 VTAIL.n23 9.3005
R379 VTAIL.n63 VTAIL.n62 9.3005
R380 VTAIL.n65 VTAIL.n64 9.3005
R381 VTAIL.n20 VTAIL.n19 9.3005
R382 VTAIL.n71 VTAIL.n70 9.3005
R383 VTAIL.n73 VTAIL.n72 9.3005
R384 VTAIL.n16 VTAIL.n15 9.3005
R385 VTAIL.n80 VTAIL.n79 9.3005
R386 VTAIL.n82 VTAIL.n81 9.3005
R387 VTAIL.n105 VTAIL.n104 9.3005
R388 VTAIL.n288 VTAIL.n287 9.3005
R389 VTAIL.n290 VTAIL.n289 9.3005
R390 VTAIL.n245 VTAIL.n244 9.3005
R391 VTAIL.n296 VTAIL.n295 9.3005
R392 VTAIL.n298 VTAIL.n297 9.3005
R393 VTAIL.n240 VTAIL.n239 9.3005
R394 VTAIL.n304 VTAIL.n303 9.3005
R395 VTAIL.n306 VTAIL.n305 9.3005
R396 VTAIL.n329 VTAIL.n328 9.3005
R397 VTAIL.n228 VTAIL.n227 9.3005
R398 VTAIL.n323 VTAIL.n322 9.3005
R399 VTAIL.n321 VTAIL.n320 9.3005
R400 VTAIL.n232 VTAIL.n231 9.3005
R401 VTAIL.n315 VTAIL.n314 9.3005
R402 VTAIL.n313 VTAIL.n312 9.3005
R403 VTAIL.n236 VTAIL.n235 9.3005
R404 VTAIL.n249 VTAIL.n248 9.3005
R405 VTAIL.n282 VTAIL.n281 9.3005
R406 VTAIL.n280 VTAIL.n279 9.3005
R407 VTAIL.n253 VTAIL.n252 9.3005
R408 VTAIL.n274 VTAIL.n273 9.3005
R409 VTAIL.n272 VTAIL.n271 9.3005
R410 VTAIL.n257 VTAIL.n256 9.3005
R411 VTAIL.n266 VTAIL.n265 9.3005
R412 VTAIL.n264 VTAIL.n263 9.3005
R413 VTAIL.n178 VTAIL.n177 9.3005
R414 VTAIL.n180 VTAIL.n179 9.3005
R415 VTAIL.n135 VTAIL.n134 9.3005
R416 VTAIL.n186 VTAIL.n185 9.3005
R417 VTAIL.n188 VTAIL.n187 9.3005
R418 VTAIL.n130 VTAIL.n129 9.3005
R419 VTAIL.n194 VTAIL.n193 9.3005
R420 VTAIL.n196 VTAIL.n195 9.3005
R421 VTAIL.n219 VTAIL.n218 9.3005
R422 VTAIL.n118 VTAIL.n117 9.3005
R423 VTAIL.n213 VTAIL.n212 9.3005
R424 VTAIL.n211 VTAIL.n210 9.3005
R425 VTAIL.n122 VTAIL.n121 9.3005
R426 VTAIL.n205 VTAIL.n204 9.3005
R427 VTAIL.n203 VTAIL.n202 9.3005
R428 VTAIL.n126 VTAIL.n125 9.3005
R429 VTAIL.n139 VTAIL.n138 9.3005
R430 VTAIL.n172 VTAIL.n171 9.3005
R431 VTAIL.n170 VTAIL.n169 9.3005
R432 VTAIL.n143 VTAIL.n142 9.3005
R433 VTAIL.n164 VTAIL.n163 9.3005
R434 VTAIL.n162 VTAIL.n161 9.3005
R435 VTAIL.n147 VTAIL.n146 9.3005
R436 VTAIL.n156 VTAIL.n155 9.3005
R437 VTAIL.n154 VTAIL.n153 9.3005
R438 VTAIL.n383 VTAIL.n358 8.92171
R439 VTAIL.n396 VTAIL.n350 8.92171
R440 VTAIL.n430 VTAIL.n429 8.92171
R441 VTAIL.n53 VTAIL.n28 8.92171
R442 VTAIL.n66 VTAIL.n20 8.92171
R443 VTAIL.n100 VTAIL.n99 8.92171
R444 VTAIL.n324 VTAIL.n323 8.92171
R445 VTAIL.n291 VTAIL.n245 8.92171
R446 VTAIL.n278 VTAIL.n253 8.92171
R447 VTAIL.n214 VTAIL.n213 8.92171
R448 VTAIL.n181 VTAIL.n135 8.92171
R449 VTAIL.n168 VTAIL.n143 8.92171
R450 VTAIL.n384 VTAIL.n356 8.14595
R451 VTAIL.n395 VTAIL.n352 8.14595
R452 VTAIL.n433 VTAIL.n334 8.14595
R453 VTAIL.n54 VTAIL.n26 8.14595
R454 VTAIL.n65 VTAIL.n22 8.14595
R455 VTAIL.n103 VTAIL.n4 8.14595
R456 VTAIL.n327 VTAIL.n228 8.14595
R457 VTAIL.n290 VTAIL.n247 8.14595
R458 VTAIL.n279 VTAIL.n251 8.14595
R459 VTAIL.n217 VTAIL.n118 8.14595
R460 VTAIL.n180 VTAIL.n137 8.14595
R461 VTAIL.n169 VTAIL.n141 8.14595
R462 VTAIL.n388 VTAIL.n387 7.3702
R463 VTAIL.n392 VTAIL.n391 7.3702
R464 VTAIL.n434 VTAIL.n332 7.3702
R465 VTAIL.n58 VTAIL.n57 7.3702
R466 VTAIL.n62 VTAIL.n61 7.3702
R467 VTAIL.n104 VTAIL.n2 7.3702
R468 VTAIL.n328 VTAIL.n226 7.3702
R469 VTAIL.n287 VTAIL.n286 7.3702
R470 VTAIL.n283 VTAIL.n282 7.3702
R471 VTAIL.n218 VTAIL.n116 7.3702
R472 VTAIL.n177 VTAIL.n176 7.3702
R473 VTAIL.n173 VTAIL.n172 7.3702
R474 VTAIL.n388 VTAIL.n354 6.59444
R475 VTAIL.n391 VTAIL.n354 6.59444
R476 VTAIL.n436 VTAIL.n332 6.59444
R477 VTAIL.n58 VTAIL.n24 6.59444
R478 VTAIL.n61 VTAIL.n24 6.59444
R479 VTAIL.n106 VTAIL.n2 6.59444
R480 VTAIL.n330 VTAIL.n226 6.59444
R481 VTAIL.n286 VTAIL.n249 6.59444
R482 VTAIL.n283 VTAIL.n249 6.59444
R483 VTAIL.n220 VTAIL.n116 6.59444
R484 VTAIL.n176 VTAIL.n139 6.59444
R485 VTAIL.n173 VTAIL.n139 6.59444
R486 VTAIL.n387 VTAIL.n356 5.81868
R487 VTAIL.n392 VTAIL.n352 5.81868
R488 VTAIL.n434 VTAIL.n433 5.81868
R489 VTAIL.n57 VTAIL.n26 5.81868
R490 VTAIL.n62 VTAIL.n22 5.81868
R491 VTAIL.n104 VTAIL.n103 5.81868
R492 VTAIL.n328 VTAIL.n327 5.81868
R493 VTAIL.n287 VTAIL.n247 5.81868
R494 VTAIL.n282 VTAIL.n251 5.81868
R495 VTAIL.n218 VTAIL.n217 5.81868
R496 VTAIL.n177 VTAIL.n137 5.81868
R497 VTAIL.n172 VTAIL.n141 5.81868
R498 VTAIL.n384 VTAIL.n383 5.04292
R499 VTAIL.n396 VTAIL.n395 5.04292
R500 VTAIL.n430 VTAIL.n334 5.04292
R501 VTAIL.n54 VTAIL.n53 5.04292
R502 VTAIL.n66 VTAIL.n65 5.04292
R503 VTAIL.n100 VTAIL.n4 5.04292
R504 VTAIL.n324 VTAIL.n228 5.04292
R505 VTAIL.n291 VTAIL.n290 5.04292
R506 VTAIL.n279 VTAIL.n278 5.04292
R507 VTAIL.n214 VTAIL.n118 5.04292
R508 VTAIL.n181 VTAIL.n180 5.04292
R509 VTAIL.n169 VTAIL.n168 5.04292
R510 VTAIL.n380 VTAIL.n358 4.26717
R511 VTAIL.n399 VTAIL.n350 4.26717
R512 VTAIL.n429 VTAIL.n336 4.26717
R513 VTAIL.n50 VTAIL.n28 4.26717
R514 VTAIL.n69 VTAIL.n20 4.26717
R515 VTAIL.n99 VTAIL.n6 4.26717
R516 VTAIL.n323 VTAIL.n230 4.26717
R517 VTAIL.n294 VTAIL.n245 4.26717
R518 VTAIL.n275 VTAIL.n253 4.26717
R519 VTAIL.n213 VTAIL.n120 4.26717
R520 VTAIL.n184 VTAIL.n135 4.26717
R521 VTAIL.n165 VTAIL.n143 4.26717
R522 VTAIL.n369 VTAIL.n365 3.70982
R523 VTAIL.n39 VTAIL.n35 3.70982
R524 VTAIL.n264 VTAIL.n260 3.70982
R525 VTAIL.n154 VTAIL.n150 3.70982
R526 VTAIL.n379 VTAIL.n360 3.49141
R527 VTAIL.n400 VTAIL.n348 3.49141
R528 VTAIL.n426 VTAIL.n425 3.49141
R529 VTAIL.n49 VTAIL.n30 3.49141
R530 VTAIL.n70 VTAIL.n18 3.49141
R531 VTAIL.n96 VTAIL.n95 3.49141
R532 VTAIL.n320 VTAIL.n319 3.49141
R533 VTAIL.n295 VTAIL.n243 3.49141
R534 VTAIL.n274 VTAIL.n255 3.49141
R535 VTAIL.n210 VTAIL.n209 3.49141
R536 VTAIL.n185 VTAIL.n133 3.49141
R537 VTAIL.n164 VTAIL.n145 3.49141
R538 VTAIL.n376 VTAIL.n375 2.71565
R539 VTAIL.n404 VTAIL.n403 2.71565
R540 VTAIL.n422 VTAIL.n338 2.71565
R541 VTAIL.n46 VTAIL.n45 2.71565
R542 VTAIL.n74 VTAIL.n73 2.71565
R543 VTAIL.n92 VTAIL.n8 2.71565
R544 VTAIL.n316 VTAIL.n232 2.71565
R545 VTAIL.n299 VTAIL.n298 2.71565
R546 VTAIL.n271 VTAIL.n270 2.71565
R547 VTAIL.n206 VTAIL.n122 2.71565
R548 VTAIL.n189 VTAIL.n188 2.71565
R549 VTAIL.n161 VTAIL.n160 2.71565
R550 VTAIL.n372 VTAIL.n362 1.93989
R551 VTAIL.n408 VTAIL.n346 1.93989
R552 VTAIL.n421 VTAIL.n340 1.93989
R553 VTAIL.n42 VTAIL.n32 1.93989
R554 VTAIL.n78 VTAIL.n16 1.93989
R555 VTAIL.n91 VTAIL.n10 1.93989
R556 VTAIL.n315 VTAIL.n234 1.93989
R557 VTAIL.n302 VTAIL.n240 1.93989
R558 VTAIL.n267 VTAIL.n257 1.93989
R559 VTAIL.n205 VTAIL.n124 1.93989
R560 VTAIL.n192 VTAIL.n130 1.93989
R561 VTAIL.n157 VTAIL.n147 1.93989
R562 VTAIL.n438 VTAIL.t19 1.71943
R563 VTAIL.n438 VTAIL.t17 1.71943
R564 VTAIL.n0 VTAIL.t16 1.71943
R565 VTAIL.n0 VTAIL.t11 1.71943
R566 VTAIL.n108 VTAIL.t4 1.71943
R567 VTAIL.n108 VTAIL.t3 1.71943
R568 VTAIL.n110 VTAIL.t8 1.71943
R569 VTAIL.n110 VTAIL.t0 1.71943
R570 VTAIL.n224 VTAIL.t5 1.71943
R571 VTAIL.n224 VTAIL.t6 1.71943
R572 VTAIL.n222 VTAIL.t7 1.71943
R573 VTAIL.n222 VTAIL.t2 1.71943
R574 VTAIL.n114 VTAIL.t13 1.71943
R575 VTAIL.n114 VTAIL.t12 1.71943
R576 VTAIL.n112 VTAIL.t15 1.71943
R577 VTAIL.n112 VTAIL.t14 1.71943
R578 VTAIL.n371 VTAIL.n364 1.16414
R579 VTAIL.n409 VTAIL.n344 1.16414
R580 VTAIL.n418 VTAIL.n417 1.16414
R581 VTAIL.n41 VTAIL.n34 1.16414
R582 VTAIL.n79 VTAIL.n14 1.16414
R583 VTAIL.n88 VTAIL.n87 1.16414
R584 VTAIL.n312 VTAIL.n311 1.16414
R585 VTAIL.n303 VTAIL.n238 1.16414
R586 VTAIL.n266 VTAIL.n259 1.16414
R587 VTAIL.n202 VTAIL.n201 1.16414
R588 VTAIL.n193 VTAIL.n128 1.16414
R589 VTAIL.n156 VTAIL.n149 1.16414
R590 VTAIL.n223 VTAIL.n221 0.698776
R591 VTAIL.n107 VTAIL.n1 0.698776
R592 VTAIL.n115 VTAIL.n113 0.457397
R593 VTAIL.n221 VTAIL.n115 0.457397
R594 VTAIL.n225 VTAIL.n223 0.457397
R595 VTAIL.n331 VTAIL.n225 0.457397
R596 VTAIL.n111 VTAIL.n109 0.457397
R597 VTAIL.n109 VTAIL.n107 0.457397
R598 VTAIL.n439 VTAIL.n437 0.457397
R599 VTAIL VTAIL.n1 0.401362
R600 VTAIL.n368 VTAIL.n367 0.388379
R601 VTAIL.n413 VTAIL.n412 0.388379
R602 VTAIL.n414 VTAIL.n342 0.388379
R603 VTAIL.n38 VTAIL.n37 0.388379
R604 VTAIL.n83 VTAIL.n82 0.388379
R605 VTAIL.n84 VTAIL.n12 0.388379
R606 VTAIL.n308 VTAIL.n236 0.388379
R607 VTAIL.n307 VTAIL.n306 0.388379
R608 VTAIL.n263 VTAIL.n262 0.388379
R609 VTAIL.n198 VTAIL.n126 0.388379
R610 VTAIL.n197 VTAIL.n196 0.388379
R611 VTAIL.n153 VTAIL.n152 0.388379
R612 VTAIL.n370 VTAIL.n369 0.155672
R613 VTAIL.n370 VTAIL.n361 0.155672
R614 VTAIL.n377 VTAIL.n361 0.155672
R615 VTAIL.n378 VTAIL.n377 0.155672
R616 VTAIL.n378 VTAIL.n357 0.155672
R617 VTAIL.n385 VTAIL.n357 0.155672
R618 VTAIL.n386 VTAIL.n385 0.155672
R619 VTAIL.n386 VTAIL.n353 0.155672
R620 VTAIL.n393 VTAIL.n353 0.155672
R621 VTAIL.n394 VTAIL.n393 0.155672
R622 VTAIL.n394 VTAIL.n349 0.155672
R623 VTAIL.n401 VTAIL.n349 0.155672
R624 VTAIL.n402 VTAIL.n401 0.155672
R625 VTAIL.n402 VTAIL.n345 0.155672
R626 VTAIL.n410 VTAIL.n345 0.155672
R627 VTAIL.n411 VTAIL.n410 0.155672
R628 VTAIL.n411 VTAIL.n341 0.155672
R629 VTAIL.n419 VTAIL.n341 0.155672
R630 VTAIL.n420 VTAIL.n419 0.155672
R631 VTAIL.n420 VTAIL.n337 0.155672
R632 VTAIL.n427 VTAIL.n337 0.155672
R633 VTAIL.n428 VTAIL.n427 0.155672
R634 VTAIL.n428 VTAIL.n333 0.155672
R635 VTAIL.n435 VTAIL.n333 0.155672
R636 VTAIL.n40 VTAIL.n39 0.155672
R637 VTAIL.n40 VTAIL.n31 0.155672
R638 VTAIL.n47 VTAIL.n31 0.155672
R639 VTAIL.n48 VTAIL.n47 0.155672
R640 VTAIL.n48 VTAIL.n27 0.155672
R641 VTAIL.n55 VTAIL.n27 0.155672
R642 VTAIL.n56 VTAIL.n55 0.155672
R643 VTAIL.n56 VTAIL.n23 0.155672
R644 VTAIL.n63 VTAIL.n23 0.155672
R645 VTAIL.n64 VTAIL.n63 0.155672
R646 VTAIL.n64 VTAIL.n19 0.155672
R647 VTAIL.n71 VTAIL.n19 0.155672
R648 VTAIL.n72 VTAIL.n71 0.155672
R649 VTAIL.n72 VTAIL.n15 0.155672
R650 VTAIL.n80 VTAIL.n15 0.155672
R651 VTAIL.n81 VTAIL.n80 0.155672
R652 VTAIL.n81 VTAIL.n11 0.155672
R653 VTAIL.n89 VTAIL.n11 0.155672
R654 VTAIL.n90 VTAIL.n89 0.155672
R655 VTAIL.n90 VTAIL.n7 0.155672
R656 VTAIL.n97 VTAIL.n7 0.155672
R657 VTAIL.n98 VTAIL.n97 0.155672
R658 VTAIL.n98 VTAIL.n3 0.155672
R659 VTAIL.n105 VTAIL.n3 0.155672
R660 VTAIL.n329 VTAIL.n227 0.155672
R661 VTAIL.n322 VTAIL.n227 0.155672
R662 VTAIL.n322 VTAIL.n321 0.155672
R663 VTAIL.n321 VTAIL.n231 0.155672
R664 VTAIL.n314 VTAIL.n231 0.155672
R665 VTAIL.n314 VTAIL.n313 0.155672
R666 VTAIL.n313 VTAIL.n235 0.155672
R667 VTAIL.n305 VTAIL.n235 0.155672
R668 VTAIL.n305 VTAIL.n304 0.155672
R669 VTAIL.n304 VTAIL.n239 0.155672
R670 VTAIL.n297 VTAIL.n239 0.155672
R671 VTAIL.n297 VTAIL.n296 0.155672
R672 VTAIL.n296 VTAIL.n244 0.155672
R673 VTAIL.n289 VTAIL.n244 0.155672
R674 VTAIL.n289 VTAIL.n288 0.155672
R675 VTAIL.n288 VTAIL.n248 0.155672
R676 VTAIL.n281 VTAIL.n248 0.155672
R677 VTAIL.n281 VTAIL.n280 0.155672
R678 VTAIL.n280 VTAIL.n252 0.155672
R679 VTAIL.n273 VTAIL.n252 0.155672
R680 VTAIL.n273 VTAIL.n272 0.155672
R681 VTAIL.n272 VTAIL.n256 0.155672
R682 VTAIL.n265 VTAIL.n256 0.155672
R683 VTAIL.n265 VTAIL.n264 0.155672
R684 VTAIL.n219 VTAIL.n117 0.155672
R685 VTAIL.n212 VTAIL.n117 0.155672
R686 VTAIL.n212 VTAIL.n211 0.155672
R687 VTAIL.n211 VTAIL.n121 0.155672
R688 VTAIL.n204 VTAIL.n121 0.155672
R689 VTAIL.n204 VTAIL.n203 0.155672
R690 VTAIL.n203 VTAIL.n125 0.155672
R691 VTAIL.n195 VTAIL.n125 0.155672
R692 VTAIL.n195 VTAIL.n194 0.155672
R693 VTAIL.n194 VTAIL.n129 0.155672
R694 VTAIL.n187 VTAIL.n129 0.155672
R695 VTAIL.n187 VTAIL.n186 0.155672
R696 VTAIL.n186 VTAIL.n134 0.155672
R697 VTAIL.n179 VTAIL.n134 0.155672
R698 VTAIL.n179 VTAIL.n178 0.155672
R699 VTAIL.n178 VTAIL.n138 0.155672
R700 VTAIL.n171 VTAIL.n138 0.155672
R701 VTAIL.n171 VTAIL.n170 0.155672
R702 VTAIL.n170 VTAIL.n142 0.155672
R703 VTAIL.n163 VTAIL.n142 0.155672
R704 VTAIL.n163 VTAIL.n162 0.155672
R705 VTAIL.n162 VTAIL.n146 0.155672
R706 VTAIL.n155 VTAIL.n146 0.155672
R707 VTAIL.n155 VTAIL.n154 0.155672
R708 VTAIL VTAIL.n439 0.0565345
R709 VDD2.n209 VDD2.n109 756.745
R710 VDD2.n100 VDD2.n0 756.745
R711 VDD2.n210 VDD2.n209 585
R712 VDD2.n208 VDD2.n207 585
R713 VDD2.n113 VDD2.n112 585
R714 VDD2.n202 VDD2.n201 585
R715 VDD2.n200 VDD2.n199 585
R716 VDD2.n117 VDD2.n116 585
R717 VDD2.n194 VDD2.n193 585
R718 VDD2.n192 VDD2.n191 585
R719 VDD2.n190 VDD2.n120 585
R720 VDD2.n124 VDD2.n121 585
R721 VDD2.n185 VDD2.n184 585
R722 VDD2.n183 VDD2.n182 585
R723 VDD2.n126 VDD2.n125 585
R724 VDD2.n177 VDD2.n176 585
R725 VDD2.n175 VDD2.n174 585
R726 VDD2.n130 VDD2.n129 585
R727 VDD2.n169 VDD2.n168 585
R728 VDD2.n167 VDD2.n166 585
R729 VDD2.n134 VDD2.n133 585
R730 VDD2.n161 VDD2.n160 585
R731 VDD2.n159 VDD2.n158 585
R732 VDD2.n138 VDD2.n137 585
R733 VDD2.n153 VDD2.n152 585
R734 VDD2.n151 VDD2.n150 585
R735 VDD2.n142 VDD2.n141 585
R736 VDD2.n145 VDD2.n144 585
R737 VDD2.n35 VDD2.n34 585
R738 VDD2.n32 VDD2.n31 585
R739 VDD2.n41 VDD2.n40 585
R740 VDD2.n43 VDD2.n42 585
R741 VDD2.n28 VDD2.n27 585
R742 VDD2.n49 VDD2.n48 585
R743 VDD2.n51 VDD2.n50 585
R744 VDD2.n24 VDD2.n23 585
R745 VDD2.n57 VDD2.n56 585
R746 VDD2.n59 VDD2.n58 585
R747 VDD2.n20 VDD2.n19 585
R748 VDD2.n65 VDD2.n64 585
R749 VDD2.n67 VDD2.n66 585
R750 VDD2.n16 VDD2.n15 585
R751 VDD2.n73 VDD2.n72 585
R752 VDD2.n76 VDD2.n75 585
R753 VDD2.n74 VDD2.n12 585
R754 VDD2.n81 VDD2.n11 585
R755 VDD2.n83 VDD2.n82 585
R756 VDD2.n85 VDD2.n84 585
R757 VDD2.n8 VDD2.n7 585
R758 VDD2.n91 VDD2.n90 585
R759 VDD2.n93 VDD2.n92 585
R760 VDD2.n4 VDD2.n3 585
R761 VDD2.n99 VDD2.n98 585
R762 VDD2.n101 VDD2.n100 585
R763 VDD2.t2 VDD2.n143 327.466
R764 VDD2.t8 VDD2.n33 327.466
R765 VDD2.n209 VDD2.n208 171.744
R766 VDD2.n208 VDD2.n112 171.744
R767 VDD2.n201 VDD2.n112 171.744
R768 VDD2.n201 VDD2.n200 171.744
R769 VDD2.n200 VDD2.n116 171.744
R770 VDD2.n193 VDD2.n116 171.744
R771 VDD2.n193 VDD2.n192 171.744
R772 VDD2.n192 VDD2.n120 171.744
R773 VDD2.n124 VDD2.n120 171.744
R774 VDD2.n184 VDD2.n124 171.744
R775 VDD2.n184 VDD2.n183 171.744
R776 VDD2.n183 VDD2.n125 171.744
R777 VDD2.n176 VDD2.n125 171.744
R778 VDD2.n176 VDD2.n175 171.744
R779 VDD2.n175 VDD2.n129 171.744
R780 VDD2.n168 VDD2.n129 171.744
R781 VDD2.n168 VDD2.n167 171.744
R782 VDD2.n167 VDD2.n133 171.744
R783 VDD2.n160 VDD2.n133 171.744
R784 VDD2.n160 VDD2.n159 171.744
R785 VDD2.n159 VDD2.n137 171.744
R786 VDD2.n152 VDD2.n137 171.744
R787 VDD2.n152 VDD2.n151 171.744
R788 VDD2.n151 VDD2.n141 171.744
R789 VDD2.n144 VDD2.n141 171.744
R790 VDD2.n34 VDD2.n31 171.744
R791 VDD2.n41 VDD2.n31 171.744
R792 VDD2.n42 VDD2.n41 171.744
R793 VDD2.n42 VDD2.n27 171.744
R794 VDD2.n49 VDD2.n27 171.744
R795 VDD2.n50 VDD2.n49 171.744
R796 VDD2.n50 VDD2.n23 171.744
R797 VDD2.n57 VDD2.n23 171.744
R798 VDD2.n58 VDD2.n57 171.744
R799 VDD2.n58 VDD2.n19 171.744
R800 VDD2.n65 VDD2.n19 171.744
R801 VDD2.n66 VDD2.n65 171.744
R802 VDD2.n66 VDD2.n15 171.744
R803 VDD2.n73 VDD2.n15 171.744
R804 VDD2.n75 VDD2.n73 171.744
R805 VDD2.n75 VDD2.n74 171.744
R806 VDD2.n74 VDD2.n11 171.744
R807 VDD2.n83 VDD2.n11 171.744
R808 VDD2.n84 VDD2.n83 171.744
R809 VDD2.n84 VDD2.n7 171.744
R810 VDD2.n91 VDD2.n7 171.744
R811 VDD2.n92 VDD2.n91 171.744
R812 VDD2.n92 VDD2.n3 171.744
R813 VDD2.n99 VDD2.n3 171.744
R814 VDD2.n100 VDD2.n99 171.744
R815 VDD2.n144 VDD2.t2 85.8723
R816 VDD2.n34 VDD2.t8 85.8723
R817 VDD2.n108 VDD2.n107 67.7026
R818 VDD2 VDD2.n217 67.6995
R819 VDD2.n106 VDD2.n105 67.4152
R820 VDD2.n216 VDD2.n215 67.4152
R821 VDD2.n106 VDD2.n104 48.3513
R822 VDD2.n214 VDD2.n213 47.8944
R823 VDD2.n214 VDD2.n108 42.1873
R824 VDD2.n145 VDD2.n143 16.3895
R825 VDD2.n35 VDD2.n33 16.3895
R826 VDD2.n191 VDD2.n190 13.1884
R827 VDD2.n82 VDD2.n81 13.1884
R828 VDD2.n194 VDD2.n119 12.8005
R829 VDD2.n189 VDD2.n121 12.8005
R830 VDD2.n146 VDD2.n142 12.8005
R831 VDD2.n36 VDD2.n32 12.8005
R832 VDD2.n80 VDD2.n12 12.8005
R833 VDD2.n85 VDD2.n10 12.8005
R834 VDD2.n195 VDD2.n117 12.0247
R835 VDD2.n186 VDD2.n185 12.0247
R836 VDD2.n150 VDD2.n149 12.0247
R837 VDD2.n40 VDD2.n39 12.0247
R838 VDD2.n77 VDD2.n76 12.0247
R839 VDD2.n86 VDD2.n8 12.0247
R840 VDD2.n199 VDD2.n198 11.249
R841 VDD2.n182 VDD2.n123 11.249
R842 VDD2.n153 VDD2.n140 11.249
R843 VDD2.n43 VDD2.n30 11.249
R844 VDD2.n72 VDD2.n14 11.249
R845 VDD2.n90 VDD2.n89 11.249
R846 VDD2.n202 VDD2.n115 10.4732
R847 VDD2.n181 VDD2.n126 10.4732
R848 VDD2.n154 VDD2.n138 10.4732
R849 VDD2.n44 VDD2.n28 10.4732
R850 VDD2.n71 VDD2.n16 10.4732
R851 VDD2.n93 VDD2.n6 10.4732
R852 VDD2.n203 VDD2.n113 9.69747
R853 VDD2.n178 VDD2.n177 9.69747
R854 VDD2.n158 VDD2.n157 9.69747
R855 VDD2.n48 VDD2.n47 9.69747
R856 VDD2.n68 VDD2.n67 9.69747
R857 VDD2.n94 VDD2.n4 9.69747
R858 VDD2.n213 VDD2.n212 9.45567
R859 VDD2.n104 VDD2.n103 9.45567
R860 VDD2.n171 VDD2.n170 9.3005
R861 VDD2.n173 VDD2.n172 9.3005
R862 VDD2.n128 VDD2.n127 9.3005
R863 VDD2.n179 VDD2.n178 9.3005
R864 VDD2.n181 VDD2.n180 9.3005
R865 VDD2.n123 VDD2.n122 9.3005
R866 VDD2.n187 VDD2.n186 9.3005
R867 VDD2.n189 VDD2.n188 9.3005
R868 VDD2.n212 VDD2.n211 9.3005
R869 VDD2.n111 VDD2.n110 9.3005
R870 VDD2.n206 VDD2.n205 9.3005
R871 VDD2.n204 VDD2.n203 9.3005
R872 VDD2.n115 VDD2.n114 9.3005
R873 VDD2.n198 VDD2.n197 9.3005
R874 VDD2.n196 VDD2.n195 9.3005
R875 VDD2.n119 VDD2.n118 9.3005
R876 VDD2.n132 VDD2.n131 9.3005
R877 VDD2.n165 VDD2.n164 9.3005
R878 VDD2.n163 VDD2.n162 9.3005
R879 VDD2.n136 VDD2.n135 9.3005
R880 VDD2.n157 VDD2.n156 9.3005
R881 VDD2.n155 VDD2.n154 9.3005
R882 VDD2.n140 VDD2.n139 9.3005
R883 VDD2.n149 VDD2.n148 9.3005
R884 VDD2.n147 VDD2.n146 9.3005
R885 VDD2.n2 VDD2.n1 9.3005
R886 VDD2.n97 VDD2.n96 9.3005
R887 VDD2.n95 VDD2.n94 9.3005
R888 VDD2.n6 VDD2.n5 9.3005
R889 VDD2.n89 VDD2.n88 9.3005
R890 VDD2.n87 VDD2.n86 9.3005
R891 VDD2.n10 VDD2.n9 9.3005
R892 VDD2.n55 VDD2.n54 9.3005
R893 VDD2.n53 VDD2.n52 9.3005
R894 VDD2.n26 VDD2.n25 9.3005
R895 VDD2.n47 VDD2.n46 9.3005
R896 VDD2.n45 VDD2.n44 9.3005
R897 VDD2.n30 VDD2.n29 9.3005
R898 VDD2.n39 VDD2.n38 9.3005
R899 VDD2.n37 VDD2.n36 9.3005
R900 VDD2.n22 VDD2.n21 9.3005
R901 VDD2.n61 VDD2.n60 9.3005
R902 VDD2.n63 VDD2.n62 9.3005
R903 VDD2.n18 VDD2.n17 9.3005
R904 VDD2.n69 VDD2.n68 9.3005
R905 VDD2.n71 VDD2.n70 9.3005
R906 VDD2.n14 VDD2.n13 9.3005
R907 VDD2.n78 VDD2.n77 9.3005
R908 VDD2.n80 VDD2.n79 9.3005
R909 VDD2.n103 VDD2.n102 9.3005
R910 VDD2.n207 VDD2.n206 8.92171
R911 VDD2.n174 VDD2.n128 8.92171
R912 VDD2.n161 VDD2.n136 8.92171
R913 VDD2.n51 VDD2.n26 8.92171
R914 VDD2.n64 VDD2.n18 8.92171
R915 VDD2.n98 VDD2.n97 8.92171
R916 VDD2.n210 VDD2.n111 8.14595
R917 VDD2.n173 VDD2.n130 8.14595
R918 VDD2.n162 VDD2.n134 8.14595
R919 VDD2.n52 VDD2.n24 8.14595
R920 VDD2.n63 VDD2.n20 8.14595
R921 VDD2.n101 VDD2.n2 8.14595
R922 VDD2.n211 VDD2.n109 7.3702
R923 VDD2.n170 VDD2.n169 7.3702
R924 VDD2.n166 VDD2.n165 7.3702
R925 VDD2.n56 VDD2.n55 7.3702
R926 VDD2.n60 VDD2.n59 7.3702
R927 VDD2.n102 VDD2.n0 7.3702
R928 VDD2.n213 VDD2.n109 6.59444
R929 VDD2.n169 VDD2.n132 6.59444
R930 VDD2.n166 VDD2.n132 6.59444
R931 VDD2.n56 VDD2.n22 6.59444
R932 VDD2.n59 VDD2.n22 6.59444
R933 VDD2.n104 VDD2.n0 6.59444
R934 VDD2.n211 VDD2.n210 5.81868
R935 VDD2.n170 VDD2.n130 5.81868
R936 VDD2.n165 VDD2.n134 5.81868
R937 VDD2.n55 VDD2.n24 5.81868
R938 VDD2.n60 VDD2.n20 5.81868
R939 VDD2.n102 VDD2.n101 5.81868
R940 VDD2.n207 VDD2.n111 5.04292
R941 VDD2.n174 VDD2.n173 5.04292
R942 VDD2.n162 VDD2.n161 5.04292
R943 VDD2.n52 VDD2.n51 5.04292
R944 VDD2.n64 VDD2.n63 5.04292
R945 VDD2.n98 VDD2.n2 5.04292
R946 VDD2.n206 VDD2.n113 4.26717
R947 VDD2.n177 VDD2.n128 4.26717
R948 VDD2.n158 VDD2.n136 4.26717
R949 VDD2.n48 VDD2.n26 4.26717
R950 VDD2.n67 VDD2.n18 4.26717
R951 VDD2.n97 VDD2.n4 4.26717
R952 VDD2.n147 VDD2.n143 3.70982
R953 VDD2.n37 VDD2.n33 3.70982
R954 VDD2.n203 VDD2.n202 3.49141
R955 VDD2.n178 VDD2.n126 3.49141
R956 VDD2.n157 VDD2.n138 3.49141
R957 VDD2.n47 VDD2.n28 3.49141
R958 VDD2.n68 VDD2.n16 3.49141
R959 VDD2.n94 VDD2.n93 3.49141
R960 VDD2.n199 VDD2.n115 2.71565
R961 VDD2.n182 VDD2.n181 2.71565
R962 VDD2.n154 VDD2.n153 2.71565
R963 VDD2.n44 VDD2.n43 2.71565
R964 VDD2.n72 VDD2.n71 2.71565
R965 VDD2.n90 VDD2.n6 2.71565
R966 VDD2.n198 VDD2.n117 1.93989
R967 VDD2.n185 VDD2.n123 1.93989
R968 VDD2.n150 VDD2.n140 1.93989
R969 VDD2.n40 VDD2.n30 1.93989
R970 VDD2.n76 VDD2.n14 1.93989
R971 VDD2.n89 VDD2.n8 1.93989
R972 VDD2.n217 VDD2.t5 1.71943
R973 VDD2.n217 VDD2.t3 1.71943
R974 VDD2.n215 VDD2.t1 1.71943
R975 VDD2.n215 VDD2.t0 1.71943
R976 VDD2.n107 VDD2.t7 1.71943
R977 VDD2.n107 VDD2.t4 1.71943
R978 VDD2.n105 VDD2.t6 1.71943
R979 VDD2.n105 VDD2.t9 1.71943
R980 VDD2.n195 VDD2.n194 1.16414
R981 VDD2.n186 VDD2.n121 1.16414
R982 VDD2.n149 VDD2.n142 1.16414
R983 VDD2.n39 VDD2.n32 1.16414
R984 VDD2.n77 VDD2.n12 1.16414
R985 VDD2.n86 VDD2.n85 1.16414
R986 VDD2.n216 VDD2.n214 0.457397
R987 VDD2.n191 VDD2.n119 0.388379
R988 VDD2.n190 VDD2.n189 0.388379
R989 VDD2.n146 VDD2.n145 0.388379
R990 VDD2.n36 VDD2.n35 0.388379
R991 VDD2.n81 VDD2.n80 0.388379
R992 VDD2.n82 VDD2.n10 0.388379
R993 VDD2 VDD2.n216 0.172914
R994 VDD2.n212 VDD2.n110 0.155672
R995 VDD2.n205 VDD2.n110 0.155672
R996 VDD2.n205 VDD2.n204 0.155672
R997 VDD2.n204 VDD2.n114 0.155672
R998 VDD2.n197 VDD2.n114 0.155672
R999 VDD2.n197 VDD2.n196 0.155672
R1000 VDD2.n196 VDD2.n118 0.155672
R1001 VDD2.n188 VDD2.n118 0.155672
R1002 VDD2.n188 VDD2.n187 0.155672
R1003 VDD2.n187 VDD2.n122 0.155672
R1004 VDD2.n180 VDD2.n122 0.155672
R1005 VDD2.n180 VDD2.n179 0.155672
R1006 VDD2.n179 VDD2.n127 0.155672
R1007 VDD2.n172 VDD2.n127 0.155672
R1008 VDD2.n172 VDD2.n171 0.155672
R1009 VDD2.n171 VDD2.n131 0.155672
R1010 VDD2.n164 VDD2.n131 0.155672
R1011 VDD2.n164 VDD2.n163 0.155672
R1012 VDD2.n163 VDD2.n135 0.155672
R1013 VDD2.n156 VDD2.n135 0.155672
R1014 VDD2.n156 VDD2.n155 0.155672
R1015 VDD2.n155 VDD2.n139 0.155672
R1016 VDD2.n148 VDD2.n139 0.155672
R1017 VDD2.n148 VDD2.n147 0.155672
R1018 VDD2.n38 VDD2.n37 0.155672
R1019 VDD2.n38 VDD2.n29 0.155672
R1020 VDD2.n45 VDD2.n29 0.155672
R1021 VDD2.n46 VDD2.n45 0.155672
R1022 VDD2.n46 VDD2.n25 0.155672
R1023 VDD2.n53 VDD2.n25 0.155672
R1024 VDD2.n54 VDD2.n53 0.155672
R1025 VDD2.n54 VDD2.n21 0.155672
R1026 VDD2.n61 VDD2.n21 0.155672
R1027 VDD2.n62 VDD2.n61 0.155672
R1028 VDD2.n62 VDD2.n17 0.155672
R1029 VDD2.n69 VDD2.n17 0.155672
R1030 VDD2.n70 VDD2.n69 0.155672
R1031 VDD2.n70 VDD2.n13 0.155672
R1032 VDD2.n78 VDD2.n13 0.155672
R1033 VDD2.n79 VDD2.n78 0.155672
R1034 VDD2.n79 VDD2.n9 0.155672
R1035 VDD2.n87 VDD2.n9 0.155672
R1036 VDD2.n88 VDD2.n87 0.155672
R1037 VDD2.n88 VDD2.n5 0.155672
R1038 VDD2.n95 VDD2.n5 0.155672
R1039 VDD2.n96 VDD2.n95 0.155672
R1040 VDD2.n96 VDD2.n1 0.155672
R1041 VDD2.n103 VDD2.n1 0.155672
R1042 VDD2.n108 VDD2.n106 0.0593781
R1043 VP.n19 VP.t6 2481.79
R1044 VP.n12 VP.t5 2481.79
R1045 VP.n4 VP.t1 2481.79
R1046 VP.n10 VP.t2 2481.79
R1047 VP.n18 VP.t9 2436.51
R1048 VP.n16 VP.t7 2436.51
R1049 VP.n1 VP.t4 2436.51
R1050 VP.n3 VP.t0 2436.51
R1051 VP.n7 VP.t8 2436.51
R1052 VP.n9 VP.t3 2436.51
R1053 VP.n5 VP.n4 161.489
R1054 VP.n20 VP.n19 161.3
R1055 VP.n6 VP.n5 161.3
R1056 VP.n8 VP.n2 161.3
R1057 VP.n11 VP.n10 161.3
R1058 VP.n17 VP.n0 161.3
R1059 VP.n15 VP.n14 161.3
R1060 VP.n13 VP.n12 161.3
R1061 VP.n13 VP.n11 45.3679
R1062 VP.n15 VP.n1 40.8975
R1063 VP.n18 VP.n17 40.8975
R1064 VP.n6 VP.n3 40.8975
R1065 VP.n9 VP.n8 40.8975
R1066 VP.n16 VP.n15 36.5157
R1067 VP.n17 VP.n16 36.5157
R1068 VP.n7 VP.n6 36.5157
R1069 VP.n8 VP.n7 36.5157
R1070 VP.n12 VP.n1 32.1338
R1071 VP.n19 VP.n18 32.1338
R1072 VP.n4 VP.n3 32.1338
R1073 VP.n10 VP.n9 32.1338
R1074 VP.n5 VP.n2 0.189894
R1075 VP.n11 VP.n2 0.189894
R1076 VP.n14 VP.n13 0.189894
R1077 VP.n14 VP.n0 0.189894
R1078 VP.n20 VP.n0 0.189894
R1079 VP VP.n20 0.0516364
R1080 VDD1.n100 VDD1.n0 756.745
R1081 VDD1.n207 VDD1.n107 756.745
R1082 VDD1.n101 VDD1.n100 585
R1083 VDD1.n99 VDD1.n98 585
R1084 VDD1.n4 VDD1.n3 585
R1085 VDD1.n93 VDD1.n92 585
R1086 VDD1.n91 VDD1.n90 585
R1087 VDD1.n8 VDD1.n7 585
R1088 VDD1.n85 VDD1.n84 585
R1089 VDD1.n83 VDD1.n82 585
R1090 VDD1.n81 VDD1.n11 585
R1091 VDD1.n15 VDD1.n12 585
R1092 VDD1.n76 VDD1.n75 585
R1093 VDD1.n74 VDD1.n73 585
R1094 VDD1.n17 VDD1.n16 585
R1095 VDD1.n68 VDD1.n67 585
R1096 VDD1.n66 VDD1.n65 585
R1097 VDD1.n21 VDD1.n20 585
R1098 VDD1.n60 VDD1.n59 585
R1099 VDD1.n58 VDD1.n57 585
R1100 VDD1.n25 VDD1.n24 585
R1101 VDD1.n52 VDD1.n51 585
R1102 VDD1.n50 VDD1.n49 585
R1103 VDD1.n29 VDD1.n28 585
R1104 VDD1.n44 VDD1.n43 585
R1105 VDD1.n42 VDD1.n41 585
R1106 VDD1.n33 VDD1.n32 585
R1107 VDD1.n36 VDD1.n35 585
R1108 VDD1.n142 VDD1.n141 585
R1109 VDD1.n139 VDD1.n138 585
R1110 VDD1.n148 VDD1.n147 585
R1111 VDD1.n150 VDD1.n149 585
R1112 VDD1.n135 VDD1.n134 585
R1113 VDD1.n156 VDD1.n155 585
R1114 VDD1.n158 VDD1.n157 585
R1115 VDD1.n131 VDD1.n130 585
R1116 VDD1.n164 VDD1.n163 585
R1117 VDD1.n166 VDD1.n165 585
R1118 VDD1.n127 VDD1.n126 585
R1119 VDD1.n172 VDD1.n171 585
R1120 VDD1.n174 VDD1.n173 585
R1121 VDD1.n123 VDD1.n122 585
R1122 VDD1.n180 VDD1.n179 585
R1123 VDD1.n183 VDD1.n182 585
R1124 VDD1.n181 VDD1.n119 585
R1125 VDD1.n188 VDD1.n118 585
R1126 VDD1.n190 VDD1.n189 585
R1127 VDD1.n192 VDD1.n191 585
R1128 VDD1.n115 VDD1.n114 585
R1129 VDD1.n198 VDD1.n197 585
R1130 VDD1.n200 VDD1.n199 585
R1131 VDD1.n111 VDD1.n110 585
R1132 VDD1.n206 VDD1.n205 585
R1133 VDD1.n208 VDD1.n207 585
R1134 VDD1.t8 VDD1.n34 327.466
R1135 VDD1.t4 VDD1.n140 327.466
R1136 VDD1.n100 VDD1.n99 171.744
R1137 VDD1.n99 VDD1.n3 171.744
R1138 VDD1.n92 VDD1.n3 171.744
R1139 VDD1.n92 VDD1.n91 171.744
R1140 VDD1.n91 VDD1.n7 171.744
R1141 VDD1.n84 VDD1.n7 171.744
R1142 VDD1.n84 VDD1.n83 171.744
R1143 VDD1.n83 VDD1.n11 171.744
R1144 VDD1.n15 VDD1.n11 171.744
R1145 VDD1.n75 VDD1.n15 171.744
R1146 VDD1.n75 VDD1.n74 171.744
R1147 VDD1.n74 VDD1.n16 171.744
R1148 VDD1.n67 VDD1.n16 171.744
R1149 VDD1.n67 VDD1.n66 171.744
R1150 VDD1.n66 VDD1.n20 171.744
R1151 VDD1.n59 VDD1.n20 171.744
R1152 VDD1.n59 VDD1.n58 171.744
R1153 VDD1.n58 VDD1.n24 171.744
R1154 VDD1.n51 VDD1.n24 171.744
R1155 VDD1.n51 VDD1.n50 171.744
R1156 VDD1.n50 VDD1.n28 171.744
R1157 VDD1.n43 VDD1.n28 171.744
R1158 VDD1.n43 VDD1.n42 171.744
R1159 VDD1.n42 VDD1.n32 171.744
R1160 VDD1.n35 VDD1.n32 171.744
R1161 VDD1.n141 VDD1.n138 171.744
R1162 VDD1.n148 VDD1.n138 171.744
R1163 VDD1.n149 VDD1.n148 171.744
R1164 VDD1.n149 VDD1.n134 171.744
R1165 VDD1.n156 VDD1.n134 171.744
R1166 VDD1.n157 VDD1.n156 171.744
R1167 VDD1.n157 VDD1.n130 171.744
R1168 VDD1.n164 VDD1.n130 171.744
R1169 VDD1.n165 VDD1.n164 171.744
R1170 VDD1.n165 VDD1.n126 171.744
R1171 VDD1.n172 VDD1.n126 171.744
R1172 VDD1.n173 VDD1.n172 171.744
R1173 VDD1.n173 VDD1.n122 171.744
R1174 VDD1.n180 VDD1.n122 171.744
R1175 VDD1.n182 VDD1.n180 171.744
R1176 VDD1.n182 VDD1.n181 171.744
R1177 VDD1.n181 VDD1.n118 171.744
R1178 VDD1.n190 VDD1.n118 171.744
R1179 VDD1.n191 VDD1.n190 171.744
R1180 VDD1.n191 VDD1.n114 171.744
R1181 VDD1.n198 VDD1.n114 171.744
R1182 VDD1.n199 VDD1.n198 171.744
R1183 VDD1.n199 VDD1.n110 171.744
R1184 VDD1.n206 VDD1.n110 171.744
R1185 VDD1.n207 VDD1.n206 171.744
R1186 VDD1.n35 VDD1.t8 85.8723
R1187 VDD1.n141 VDD1.t4 85.8723
R1188 VDD1.n215 VDD1.n214 67.7026
R1189 VDD1.n213 VDD1.n212 67.4152
R1190 VDD1.n106 VDD1.n105 67.4152
R1191 VDD1.n217 VDD1.n216 67.415
R1192 VDD1.n106 VDD1.n104 48.3513
R1193 VDD1.n213 VDD1.n211 48.3513
R1194 VDD1.n217 VDD1.n215 42.9987
R1195 VDD1.n36 VDD1.n34 16.3895
R1196 VDD1.n142 VDD1.n140 16.3895
R1197 VDD1.n82 VDD1.n81 13.1884
R1198 VDD1.n189 VDD1.n188 13.1884
R1199 VDD1.n85 VDD1.n10 12.8005
R1200 VDD1.n80 VDD1.n12 12.8005
R1201 VDD1.n37 VDD1.n33 12.8005
R1202 VDD1.n143 VDD1.n139 12.8005
R1203 VDD1.n187 VDD1.n119 12.8005
R1204 VDD1.n192 VDD1.n117 12.8005
R1205 VDD1.n86 VDD1.n8 12.0247
R1206 VDD1.n77 VDD1.n76 12.0247
R1207 VDD1.n41 VDD1.n40 12.0247
R1208 VDD1.n147 VDD1.n146 12.0247
R1209 VDD1.n184 VDD1.n183 12.0247
R1210 VDD1.n193 VDD1.n115 12.0247
R1211 VDD1.n90 VDD1.n89 11.249
R1212 VDD1.n73 VDD1.n14 11.249
R1213 VDD1.n44 VDD1.n31 11.249
R1214 VDD1.n150 VDD1.n137 11.249
R1215 VDD1.n179 VDD1.n121 11.249
R1216 VDD1.n197 VDD1.n196 11.249
R1217 VDD1.n93 VDD1.n6 10.4732
R1218 VDD1.n72 VDD1.n17 10.4732
R1219 VDD1.n45 VDD1.n29 10.4732
R1220 VDD1.n151 VDD1.n135 10.4732
R1221 VDD1.n178 VDD1.n123 10.4732
R1222 VDD1.n200 VDD1.n113 10.4732
R1223 VDD1.n94 VDD1.n4 9.69747
R1224 VDD1.n69 VDD1.n68 9.69747
R1225 VDD1.n49 VDD1.n48 9.69747
R1226 VDD1.n155 VDD1.n154 9.69747
R1227 VDD1.n175 VDD1.n174 9.69747
R1228 VDD1.n201 VDD1.n111 9.69747
R1229 VDD1.n104 VDD1.n103 9.45567
R1230 VDD1.n211 VDD1.n210 9.45567
R1231 VDD1.n62 VDD1.n61 9.3005
R1232 VDD1.n64 VDD1.n63 9.3005
R1233 VDD1.n19 VDD1.n18 9.3005
R1234 VDD1.n70 VDD1.n69 9.3005
R1235 VDD1.n72 VDD1.n71 9.3005
R1236 VDD1.n14 VDD1.n13 9.3005
R1237 VDD1.n78 VDD1.n77 9.3005
R1238 VDD1.n80 VDD1.n79 9.3005
R1239 VDD1.n103 VDD1.n102 9.3005
R1240 VDD1.n2 VDD1.n1 9.3005
R1241 VDD1.n97 VDD1.n96 9.3005
R1242 VDD1.n95 VDD1.n94 9.3005
R1243 VDD1.n6 VDD1.n5 9.3005
R1244 VDD1.n89 VDD1.n88 9.3005
R1245 VDD1.n87 VDD1.n86 9.3005
R1246 VDD1.n10 VDD1.n9 9.3005
R1247 VDD1.n23 VDD1.n22 9.3005
R1248 VDD1.n56 VDD1.n55 9.3005
R1249 VDD1.n54 VDD1.n53 9.3005
R1250 VDD1.n27 VDD1.n26 9.3005
R1251 VDD1.n48 VDD1.n47 9.3005
R1252 VDD1.n46 VDD1.n45 9.3005
R1253 VDD1.n31 VDD1.n30 9.3005
R1254 VDD1.n40 VDD1.n39 9.3005
R1255 VDD1.n38 VDD1.n37 9.3005
R1256 VDD1.n109 VDD1.n108 9.3005
R1257 VDD1.n204 VDD1.n203 9.3005
R1258 VDD1.n202 VDD1.n201 9.3005
R1259 VDD1.n113 VDD1.n112 9.3005
R1260 VDD1.n196 VDD1.n195 9.3005
R1261 VDD1.n194 VDD1.n193 9.3005
R1262 VDD1.n117 VDD1.n116 9.3005
R1263 VDD1.n162 VDD1.n161 9.3005
R1264 VDD1.n160 VDD1.n159 9.3005
R1265 VDD1.n133 VDD1.n132 9.3005
R1266 VDD1.n154 VDD1.n153 9.3005
R1267 VDD1.n152 VDD1.n151 9.3005
R1268 VDD1.n137 VDD1.n136 9.3005
R1269 VDD1.n146 VDD1.n145 9.3005
R1270 VDD1.n144 VDD1.n143 9.3005
R1271 VDD1.n129 VDD1.n128 9.3005
R1272 VDD1.n168 VDD1.n167 9.3005
R1273 VDD1.n170 VDD1.n169 9.3005
R1274 VDD1.n125 VDD1.n124 9.3005
R1275 VDD1.n176 VDD1.n175 9.3005
R1276 VDD1.n178 VDD1.n177 9.3005
R1277 VDD1.n121 VDD1.n120 9.3005
R1278 VDD1.n185 VDD1.n184 9.3005
R1279 VDD1.n187 VDD1.n186 9.3005
R1280 VDD1.n210 VDD1.n209 9.3005
R1281 VDD1.n98 VDD1.n97 8.92171
R1282 VDD1.n65 VDD1.n19 8.92171
R1283 VDD1.n52 VDD1.n27 8.92171
R1284 VDD1.n158 VDD1.n133 8.92171
R1285 VDD1.n171 VDD1.n125 8.92171
R1286 VDD1.n205 VDD1.n204 8.92171
R1287 VDD1.n101 VDD1.n2 8.14595
R1288 VDD1.n64 VDD1.n21 8.14595
R1289 VDD1.n53 VDD1.n25 8.14595
R1290 VDD1.n159 VDD1.n131 8.14595
R1291 VDD1.n170 VDD1.n127 8.14595
R1292 VDD1.n208 VDD1.n109 8.14595
R1293 VDD1.n102 VDD1.n0 7.3702
R1294 VDD1.n61 VDD1.n60 7.3702
R1295 VDD1.n57 VDD1.n56 7.3702
R1296 VDD1.n163 VDD1.n162 7.3702
R1297 VDD1.n167 VDD1.n166 7.3702
R1298 VDD1.n209 VDD1.n107 7.3702
R1299 VDD1.n104 VDD1.n0 6.59444
R1300 VDD1.n60 VDD1.n23 6.59444
R1301 VDD1.n57 VDD1.n23 6.59444
R1302 VDD1.n163 VDD1.n129 6.59444
R1303 VDD1.n166 VDD1.n129 6.59444
R1304 VDD1.n211 VDD1.n107 6.59444
R1305 VDD1.n102 VDD1.n101 5.81868
R1306 VDD1.n61 VDD1.n21 5.81868
R1307 VDD1.n56 VDD1.n25 5.81868
R1308 VDD1.n162 VDD1.n131 5.81868
R1309 VDD1.n167 VDD1.n127 5.81868
R1310 VDD1.n209 VDD1.n208 5.81868
R1311 VDD1.n98 VDD1.n2 5.04292
R1312 VDD1.n65 VDD1.n64 5.04292
R1313 VDD1.n53 VDD1.n52 5.04292
R1314 VDD1.n159 VDD1.n158 5.04292
R1315 VDD1.n171 VDD1.n170 5.04292
R1316 VDD1.n205 VDD1.n109 5.04292
R1317 VDD1.n97 VDD1.n4 4.26717
R1318 VDD1.n68 VDD1.n19 4.26717
R1319 VDD1.n49 VDD1.n27 4.26717
R1320 VDD1.n155 VDD1.n133 4.26717
R1321 VDD1.n174 VDD1.n125 4.26717
R1322 VDD1.n204 VDD1.n111 4.26717
R1323 VDD1.n38 VDD1.n34 3.70982
R1324 VDD1.n144 VDD1.n140 3.70982
R1325 VDD1.n94 VDD1.n93 3.49141
R1326 VDD1.n69 VDD1.n17 3.49141
R1327 VDD1.n48 VDD1.n29 3.49141
R1328 VDD1.n154 VDD1.n135 3.49141
R1329 VDD1.n175 VDD1.n123 3.49141
R1330 VDD1.n201 VDD1.n200 3.49141
R1331 VDD1.n90 VDD1.n6 2.71565
R1332 VDD1.n73 VDD1.n72 2.71565
R1333 VDD1.n45 VDD1.n44 2.71565
R1334 VDD1.n151 VDD1.n150 2.71565
R1335 VDD1.n179 VDD1.n178 2.71565
R1336 VDD1.n197 VDD1.n113 2.71565
R1337 VDD1.n89 VDD1.n8 1.93989
R1338 VDD1.n76 VDD1.n14 1.93989
R1339 VDD1.n41 VDD1.n31 1.93989
R1340 VDD1.n147 VDD1.n137 1.93989
R1341 VDD1.n183 VDD1.n121 1.93989
R1342 VDD1.n196 VDD1.n115 1.93989
R1343 VDD1.n216 VDD1.t6 1.71943
R1344 VDD1.n216 VDD1.t7 1.71943
R1345 VDD1.n105 VDD1.t9 1.71943
R1346 VDD1.n105 VDD1.t1 1.71943
R1347 VDD1.n214 VDD1.t0 1.71943
R1348 VDD1.n214 VDD1.t3 1.71943
R1349 VDD1.n212 VDD1.t5 1.71943
R1350 VDD1.n212 VDD1.t2 1.71943
R1351 VDD1.n86 VDD1.n85 1.16414
R1352 VDD1.n77 VDD1.n12 1.16414
R1353 VDD1.n40 VDD1.n33 1.16414
R1354 VDD1.n146 VDD1.n139 1.16414
R1355 VDD1.n184 VDD1.n119 1.16414
R1356 VDD1.n193 VDD1.n192 1.16414
R1357 VDD1.n82 VDD1.n10 0.388379
R1358 VDD1.n81 VDD1.n80 0.388379
R1359 VDD1.n37 VDD1.n36 0.388379
R1360 VDD1.n143 VDD1.n142 0.388379
R1361 VDD1.n188 VDD1.n187 0.388379
R1362 VDD1.n189 VDD1.n117 0.388379
R1363 VDD1 VDD1.n217 0.284983
R1364 VDD1 VDD1.n106 0.172914
R1365 VDD1.n103 VDD1.n1 0.155672
R1366 VDD1.n96 VDD1.n1 0.155672
R1367 VDD1.n96 VDD1.n95 0.155672
R1368 VDD1.n95 VDD1.n5 0.155672
R1369 VDD1.n88 VDD1.n5 0.155672
R1370 VDD1.n88 VDD1.n87 0.155672
R1371 VDD1.n87 VDD1.n9 0.155672
R1372 VDD1.n79 VDD1.n9 0.155672
R1373 VDD1.n79 VDD1.n78 0.155672
R1374 VDD1.n78 VDD1.n13 0.155672
R1375 VDD1.n71 VDD1.n13 0.155672
R1376 VDD1.n71 VDD1.n70 0.155672
R1377 VDD1.n70 VDD1.n18 0.155672
R1378 VDD1.n63 VDD1.n18 0.155672
R1379 VDD1.n63 VDD1.n62 0.155672
R1380 VDD1.n62 VDD1.n22 0.155672
R1381 VDD1.n55 VDD1.n22 0.155672
R1382 VDD1.n55 VDD1.n54 0.155672
R1383 VDD1.n54 VDD1.n26 0.155672
R1384 VDD1.n47 VDD1.n26 0.155672
R1385 VDD1.n47 VDD1.n46 0.155672
R1386 VDD1.n46 VDD1.n30 0.155672
R1387 VDD1.n39 VDD1.n30 0.155672
R1388 VDD1.n39 VDD1.n38 0.155672
R1389 VDD1.n145 VDD1.n144 0.155672
R1390 VDD1.n145 VDD1.n136 0.155672
R1391 VDD1.n152 VDD1.n136 0.155672
R1392 VDD1.n153 VDD1.n152 0.155672
R1393 VDD1.n153 VDD1.n132 0.155672
R1394 VDD1.n160 VDD1.n132 0.155672
R1395 VDD1.n161 VDD1.n160 0.155672
R1396 VDD1.n161 VDD1.n128 0.155672
R1397 VDD1.n168 VDD1.n128 0.155672
R1398 VDD1.n169 VDD1.n168 0.155672
R1399 VDD1.n169 VDD1.n124 0.155672
R1400 VDD1.n176 VDD1.n124 0.155672
R1401 VDD1.n177 VDD1.n176 0.155672
R1402 VDD1.n177 VDD1.n120 0.155672
R1403 VDD1.n185 VDD1.n120 0.155672
R1404 VDD1.n186 VDD1.n185 0.155672
R1405 VDD1.n186 VDD1.n116 0.155672
R1406 VDD1.n194 VDD1.n116 0.155672
R1407 VDD1.n195 VDD1.n194 0.155672
R1408 VDD1.n195 VDD1.n112 0.155672
R1409 VDD1.n202 VDD1.n112 0.155672
R1410 VDD1.n203 VDD1.n202 0.155672
R1411 VDD1.n203 VDD1.n108 0.155672
R1412 VDD1.n210 VDD1.n108 0.155672
R1413 VDD1.n215 VDD1.n213 0.0593781
R1414 B.n136 B.t0 2515
R1415 B.n306 B.t9 2515
R1416 B.n48 B.t6 2515
R1417 B.n42 B.t3 2515
R1418 B.n403 B.n402 585
R1419 B.n401 B.n100 585
R1420 B.n400 B.n399 585
R1421 B.n398 B.n101 585
R1422 B.n397 B.n396 585
R1423 B.n395 B.n102 585
R1424 B.n394 B.n393 585
R1425 B.n392 B.n103 585
R1426 B.n391 B.n390 585
R1427 B.n389 B.n104 585
R1428 B.n388 B.n387 585
R1429 B.n386 B.n105 585
R1430 B.n385 B.n384 585
R1431 B.n383 B.n106 585
R1432 B.n382 B.n381 585
R1433 B.n380 B.n107 585
R1434 B.n379 B.n378 585
R1435 B.n377 B.n108 585
R1436 B.n376 B.n375 585
R1437 B.n374 B.n109 585
R1438 B.n373 B.n372 585
R1439 B.n371 B.n110 585
R1440 B.n370 B.n369 585
R1441 B.n368 B.n111 585
R1442 B.n367 B.n366 585
R1443 B.n365 B.n112 585
R1444 B.n364 B.n363 585
R1445 B.n362 B.n113 585
R1446 B.n361 B.n360 585
R1447 B.n359 B.n114 585
R1448 B.n358 B.n357 585
R1449 B.n356 B.n115 585
R1450 B.n355 B.n354 585
R1451 B.n353 B.n116 585
R1452 B.n352 B.n351 585
R1453 B.n350 B.n117 585
R1454 B.n349 B.n348 585
R1455 B.n347 B.n118 585
R1456 B.n346 B.n345 585
R1457 B.n344 B.n119 585
R1458 B.n343 B.n342 585
R1459 B.n341 B.n120 585
R1460 B.n340 B.n339 585
R1461 B.n338 B.n121 585
R1462 B.n337 B.n336 585
R1463 B.n335 B.n122 585
R1464 B.n334 B.n333 585
R1465 B.n332 B.n123 585
R1466 B.n331 B.n330 585
R1467 B.n329 B.n124 585
R1468 B.n328 B.n327 585
R1469 B.n326 B.n125 585
R1470 B.n325 B.n324 585
R1471 B.n323 B.n126 585
R1472 B.n322 B.n321 585
R1473 B.n320 B.n127 585
R1474 B.n319 B.n318 585
R1475 B.n317 B.n128 585
R1476 B.n316 B.n315 585
R1477 B.n314 B.n129 585
R1478 B.n313 B.n312 585
R1479 B.n311 B.n130 585
R1480 B.n310 B.n309 585
R1481 B.n305 B.n131 585
R1482 B.n304 B.n303 585
R1483 B.n302 B.n132 585
R1484 B.n301 B.n300 585
R1485 B.n299 B.n133 585
R1486 B.n298 B.n297 585
R1487 B.n296 B.n134 585
R1488 B.n295 B.n294 585
R1489 B.n292 B.n135 585
R1490 B.n291 B.n290 585
R1491 B.n289 B.n138 585
R1492 B.n288 B.n287 585
R1493 B.n286 B.n139 585
R1494 B.n285 B.n284 585
R1495 B.n283 B.n140 585
R1496 B.n282 B.n281 585
R1497 B.n280 B.n141 585
R1498 B.n279 B.n278 585
R1499 B.n277 B.n142 585
R1500 B.n276 B.n275 585
R1501 B.n274 B.n143 585
R1502 B.n273 B.n272 585
R1503 B.n271 B.n144 585
R1504 B.n270 B.n269 585
R1505 B.n268 B.n145 585
R1506 B.n267 B.n266 585
R1507 B.n265 B.n146 585
R1508 B.n264 B.n263 585
R1509 B.n262 B.n147 585
R1510 B.n261 B.n260 585
R1511 B.n259 B.n148 585
R1512 B.n258 B.n257 585
R1513 B.n256 B.n149 585
R1514 B.n255 B.n254 585
R1515 B.n253 B.n150 585
R1516 B.n252 B.n251 585
R1517 B.n250 B.n151 585
R1518 B.n249 B.n248 585
R1519 B.n247 B.n152 585
R1520 B.n246 B.n245 585
R1521 B.n244 B.n153 585
R1522 B.n243 B.n242 585
R1523 B.n241 B.n154 585
R1524 B.n240 B.n239 585
R1525 B.n238 B.n155 585
R1526 B.n237 B.n236 585
R1527 B.n235 B.n156 585
R1528 B.n234 B.n233 585
R1529 B.n232 B.n157 585
R1530 B.n231 B.n230 585
R1531 B.n229 B.n158 585
R1532 B.n228 B.n227 585
R1533 B.n226 B.n159 585
R1534 B.n225 B.n224 585
R1535 B.n223 B.n160 585
R1536 B.n222 B.n221 585
R1537 B.n220 B.n161 585
R1538 B.n219 B.n218 585
R1539 B.n217 B.n162 585
R1540 B.n216 B.n215 585
R1541 B.n214 B.n163 585
R1542 B.n213 B.n212 585
R1543 B.n211 B.n164 585
R1544 B.n210 B.n209 585
R1545 B.n208 B.n165 585
R1546 B.n207 B.n206 585
R1547 B.n205 B.n166 585
R1548 B.n204 B.n203 585
R1549 B.n202 B.n167 585
R1550 B.n201 B.n200 585
R1551 B.n404 B.n99 585
R1552 B.n406 B.n405 585
R1553 B.n407 B.n98 585
R1554 B.n409 B.n408 585
R1555 B.n410 B.n97 585
R1556 B.n412 B.n411 585
R1557 B.n413 B.n96 585
R1558 B.n415 B.n414 585
R1559 B.n416 B.n95 585
R1560 B.n418 B.n417 585
R1561 B.n419 B.n94 585
R1562 B.n421 B.n420 585
R1563 B.n422 B.n93 585
R1564 B.n424 B.n423 585
R1565 B.n425 B.n92 585
R1566 B.n427 B.n426 585
R1567 B.n428 B.n91 585
R1568 B.n430 B.n429 585
R1569 B.n431 B.n90 585
R1570 B.n433 B.n432 585
R1571 B.n434 B.n89 585
R1572 B.n436 B.n435 585
R1573 B.n437 B.n88 585
R1574 B.n439 B.n438 585
R1575 B.n440 B.n87 585
R1576 B.n442 B.n441 585
R1577 B.n443 B.n86 585
R1578 B.n445 B.n444 585
R1579 B.n446 B.n85 585
R1580 B.n448 B.n447 585
R1581 B.n449 B.n84 585
R1582 B.n451 B.n450 585
R1583 B.n452 B.n83 585
R1584 B.n454 B.n453 585
R1585 B.n455 B.n82 585
R1586 B.n457 B.n456 585
R1587 B.n658 B.n657 585
R1588 B.n656 B.n11 585
R1589 B.n655 B.n654 585
R1590 B.n653 B.n12 585
R1591 B.n652 B.n651 585
R1592 B.n650 B.n13 585
R1593 B.n649 B.n648 585
R1594 B.n647 B.n14 585
R1595 B.n646 B.n645 585
R1596 B.n644 B.n15 585
R1597 B.n643 B.n642 585
R1598 B.n641 B.n16 585
R1599 B.n640 B.n639 585
R1600 B.n638 B.n17 585
R1601 B.n637 B.n636 585
R1602 B.n635 B.n18 585
R1603 B.n634 B.n633 585
R1604 B.n632 B.n19 585
R1605 B.n631 B.n630 585
R1606 B.n629 B.n20 585
R1607 B.n628 B.n627 585
R1608 B.n626 B.n21 585
R1609 B.n625 B.n624 585
R1610 B.n623 B.n22 585
R1611 B.n622 B.n621 585
R1612 B.n620 B.n23 585
R1613 B.n619 B.n618 585
R1614 B.n617 B.n24 585
R1615 B.n616 B.n615 585
R1616 B.n614 B.n25 585
R1617 B.n613 B.n612 585
R1618 B.n611 B.n26 585
R1619 B.n610 B.n609 585
R1620 B.n608 B.n27 585
R1621 B.n607 B.n606 585
R1622 B.n605 B.n28 585
R1623 B.n604 B.n603 585
R1624 B.n602 B.n29 585
R1625 B.n601 B.n600 585
R1626 B.n599 B.n30 585
R1627 B.n598 B.n597 585
R1628 B.n596 B.n31 585
R1629 B.n595 B.n594 585
R1630 B.n593 B.n32 585
R1631 B.n592 B.n591 585
R1632 B.n590 B.n33 585
R1633 B.n589 B.n588 585
R1634 B.n587 B.n34 585
R1635 B.n586 B.n585 585
R1636 B.n584 B.n35 585
R1637 B.n583 B.n582 585
R1638 B.n581 B.n36 585
R1639 B.n580 B.n579 585
R1640 B.n578 B.n37 585
R1641 B.n577 B.n576 585
R1642 B.n575 B.n38 585
R1643 B.n574 B.n573 585
R1644 B.n572 B.n39 585
R1645 B.n571 B.n570 585
R1646 B.n569 B.n40 585
R1647 B.n568 B.n567 585
R1648 B.n566 B.n41 585
R1649 B.n564 B.n563 585
R1650 B.n562 B.n44 585
R1651 B.n561 B.n560 585
R1652 B.n559 B.n45 585
R1653 B.n558 B.n557 585
R1654 B.n556 B.n46 585
R1655 B.n555 B.n554 585
R1656 B.n553 B.n47 585
R1657 B.n552 B.n551 585
R1658 B.n550 B.n549 585
R1659 B.n548 B.n51 585
R1660 B.n547 B.n546 585
R1661 B.n545 B.n52 585
R1662 B.n544 B.n543 585
R1663 B.n542 B.n53 585
R1664 B.n541 B.n540 585
R1665 B.n539 B.n54 585
R1666 B.n538 B.n537 585
R1667 B.n536 B.n55 585
R1668 B.n535 B.n534 585
R1669 B.n533 B.n56 585
R1670 B.n532 B.n531 585
R1671 B.n530 B.n57 585
R1672 B.n529 B.n528 585
R1673 B.n527 B.n58 585
R1674 B.n526 B.n525 585
R1675 B.n524 B.n59 585
R1676 B.n523 B.n522 585
R1677 B.n521 B.n60 585
R1678 B.n520 B.n519 585
R1679 B.n518 B.n61 585
R1680 B.n517 B.n516 585
R1681 B.n515 B.n62 585
R1682 B.n514 B.n513 585
R1683 B.n512 B.n63 585
R1684 B.n511 B.n510 585
R1685 B.n509 B.n64 585
R1686 B.n508 B.n507 585
R1687 B.n506 B.n65 585
R1688 B.n505 B.n504 585
R1689 B.n503 B.n66 585
R1690 B.n502 B.n501 585
R1691 B.n500 B.n67 585
R1692 B.n499 B.n498 585
R1693 B.n497 B.n68 585
R1694 B.n496 B.n495 585
R1695 B.n494 B.n69 585
R1696 B.n493 B.n492 585
R1697 B.n491 B.n70 585
R1698 B.n490 B.n489 585
R1699 B.n488 B.n71 585
R1700 B.n487 B.n486 585
R1701 B.n485 B.n72 585
R1702 B.n484 B.n483 585
R1703 B.n482 B.n73 585
R1704 B.n481 B.n480 585
R1705 B.n479 B.n74 585
R1706 B.n478 B.n477 585
R1707 B.n476 B.n75 585
R1708 B.n475 B.n474 585
R1709 B.n473 B.n76 585
R1710 B.n472 B.n471 585
R1711 B.n470 B.n77 585
R1712 B.n469 B.n468 585
R1713 B.n467 B.n78 585
R1714 B.n466 B.n465 585
R1715 B.n464 B.n79 585
R1716 B.n463 B.n462 585
R1717 B.n461 B.n80 585
R1718 B.n460 B.n459 585
R1719 B.n458 B.n81 585
R1720 B.n659 B.n10 585
R1721 B.n661 B.n660 585
R1722 B.n662 B.n9 585
R1723 B.n664 B.n663 585
R1724 B.n665 B.n8 585
R1725 B.n667 B.n666 585
R1726 B.n668 B.n7 585
R1727 B.n670 B.n669 585
R1728 B.n671 B.n6 585
R1729 B.n673 B.n672 585
R1730 B.n674 B.n5 585
R1731 B.n676 B.n675 585
R1732 B.n677 B.n4 585
R1733 B.n679 B.n678 585
R1734 B.n680 B.n3 585
R1735 B.n682 B.n681 585
R1736 B.n683 B.n0 585
R1737 B.n2 B.n1 585
R1738 B.n177 B.n176 585
R1739 B.n178 B.n175 585
R1740 B.n180 B.n179 585
R1741 B.n181 B.n174 585
R1742 B.n183 B.n182 585
R1743 B.n184 B.n173 585
R1744 B.n186 B.n185 585
R1745 B.n187 B.n172 585
R1746 B.n189 B.n188 585
R1747 B.n190 B.n171 585
R1748 B.n192 B.n191 585
R1749 B.n193 B.n170 585
R1750 B.n195 B.n194 585
R1751 B.n196 B.n169 585
R1752 B.n198 B.n197 585
R1753 B.n199 B.n168 585
R1754 B.n200 B.n199 530.939
R1755 B.n402 B.n99 530.939
R1756 B.n456 B.n81 530.939
R1757 B.n659 B.n658 530.939
R1758 B.n306 B.t10 510.423
R1759 B.n48 B.t8 510.423
R1760 B.n136 B.t1 510.423
R1761 B.n42 B.t5 510.423
R1762 B.n307 B.t11 500.144
R1763 B.n49 B.t7 500.144
R1764 B.n137 B.t2 500.144
R1765 B.n43 B.t4 500.144
R1766 B.n685 B.n684 256.663
R1767 B.n684 B.n683 235.042
R1768 B.n684 B.n2 235.042
R1769 B.n200 B.n167 163.367
R1770 B.n204 B.n167 163.367
R1771 B.n205 B.n204 163.367
R1772 B.n206 B.n205 163.367
R1773 B.n206 B.n165 163.367
R1774 B.n210 B.n165 163.367
R1775 B.n211 B.n210 163.367
R1776 B.n212 B.n211 163.367
R1777 B.n212 B.n163 163.367
R1778 B.n216 B.n163 163.367
R1779 B.n217 B.n216 163.367
R1780 B.n218 B.n217 163.367
R1781 B.n218 B.n161 163.367
R1782 B.n222 B.n161 163.367
R1783 B.n223 B.n222 163.367
R1784 B.n224 B.n223 163.367
R1785 B.n224 B.n159 163.367
R1786 B.n228 B.n159 163.367
R1787 B.n229 B.n228 163.367
R1788 B.n230 B.n229 163.367
R1789 B.n230 B.n157 163.367
R1790 B.n234 B.n157 163.367
R1791 B.n235 B.n234 163.367
R1792 B.n236 B.n235 163.367
R1793 B.n236 B.n155 163.367
R1794 B.n240 B.n155 163.367
R1795 B.n241 B.n240 163.367
R1796 B.n242 B.n241 163.367
R1797 B.n242 B.n153 163.367
R1798 B.n246 B.n153 163.367
R1799 B.n247 B.n246 163.367
R1800 B.n248 B.n247 163.367
R1801 B.n248 B.n151 163.367
R1802 B.n252 B.n151 163.367
R1803 B.n253 B.n252 163.367
R1804 B.n254 B.n253 163.367
R1805 B.n254 B.n149 163.367
R1806 B.n258 B.n149 163.367
R1807 B.n259 B.n258 163.367
R1808 B.n260 B.n259 163.367
R1809 B.n260 B.n147 163.367
R1810 B.n264 B.n147 163.367
R1811 B.n265 B.n264 163.367
R1812 B.n266 B.n265 163.367
R1813 B.n266 B.n145 163.367
R1814 B.n270 B.n145 163.367
R1815 B.n271 B.n270 163.367
R1816 B.n272 B.n271 163.367
R1817 B.n272 B.n143 163.367
R1818 B.n276 B.n143 163.367
R1819 B.n277 B.n276 163.367
R1820 B.n278 B.n277 163.367
R1821 B.n278 B.n141 163.367
R1822 B.n282 B.n141 163.367
R1823 B.n283 B.n282 163.367
R1824 B.n284 B.n283 163.367
R1825 B.n284 B.n139 163.367
R1826 B.n288 B.n139 163.367
R1827 B.n289 B.n288 163.367
R1828 B.n290 B.n289 163.367
R1829 B.n290 B.n135 163.367
R1830 B.n295 B.n135 163.367
R1831 B.n296 B.n295 163.367
R1832 B.n297 B.n296 163.367
R1833 B.n297 B.n133 163.367
R1834 B.n301 B.n133 163.367
R1835 B.n302 B.n301 163.367
R1836 B.n303 B.n302 163.367
R1837 B.n303 B.n131 163.367
R1838 B.n310 B.n131 163.367
R1839 B.n311 B.n310 163.367
R1840 B.n312 B.n311 163.367
R1841 B.n312 B.n129 163.367
R1842 B.n316 B.n129 163.367
R1843 B.n317 B.n316 163.367
R1844 B.n318 B.n317 163.367
R1845 B.n318 B.n127 163.367
R1846 B.n322 B.n127 163.367
R1847 B.n323 B.n322 163.367
R1848 B.n324 B.n323 163.367
R1849 B.n324 B.n125 163.367
R1850 B.n328 B.n125 163.367
R1851 B.n329 B.n328 163.367
R1852 B.n330 B.n329 163.367
R1853 B.n330 B.n123 163.367
R1854 B.n334 B.n123 163.367
R1855 B.n335 B.n334 163.367
R1856 B.n336 B.n335 163.367
R1857 B.n336 B.n121 163.367
R1858 B.n340 B.n121 163.367
R1859 B.n341 B.n340 163.367
R1860 B.n342 B.n341 163.367
R1861 B.n342 B.n119 163.367
R1862 B.n346 B.n119 163.367
R1863 B.n347 B.n346 163.367
R1864 B.n348 B.n347 163.367
R1865 B.n348 B.n117 163.367
R1866 B.n352 B.n117 163.367
R1867 B.n353 B.n352 163.367
R1868 B.n354 B.n353 163.367
R1869 B.n354 B.n115 163.367
R1870 B.n358 B.n115 163.367
R1871 B.n359 B.n358 163.367
R1872 B.n360 B.n359 163.367
R1873 B.n360 B.n113 163.367
R1874 B.n364 B.n113 163.367
R1875 B.n365 B.n364 163.367
R1876 B.n366 B.n365 163.367
R1877 B.n366 B.n111 163.367
R1878 B.n370 B.n111 163.367
R1879 B.n371 B.n370 163.367
R1880 B.n372 B.n371 163.367
R1881 B.n372 B.n109 163.367
R1882 B.n376 B.n109 163.367
R1883 B.n377 B.n376 163.367
R1884 B.n378 B.n377 163.367
R1885 B.n378 B.n107 163.367
R1886 B.n382 B.n107 163.367
R1887 B.n383 B.n382 163.367
R1888 B.n384 B.n383 163.367
R1889 B.n384 B.n105 163.367
R1890 B.n388 B.n105 163.367
R1891 B.n389 B.n388 163.367
R1892 B.n390 B.n389 163.367
R1893 B.n390 B.n103 163.367
R1894 B.n394 B.n103 163.367
R1895 B.n395 B.n394 163.367
R1896 B.n396 B.n395 163.367
R1897 B.n396 B.n101 163.367
R1898 B.n400 B.n101 163.367
R1899 B.n401 B.n400 163.367
R1900 B.n402 B.n401 163.367
R1901 B.n456 B.n455 163.367
R1902 B.n455 B.n454 163.367
R1903 B.n454 B.n83 163.367
R1904 B.n450 B.n83 163.367
R1905 B.n450 B.n449 163.367
R1906 B.n449 B.n448 163.367
R1907 B.n448 B.n85 163.367
R1908 B.n444 B.n85 163.367
R1909 B.n444 B.n443 163.367
R1910 B.n443 B.n442 163.367
R1911 B.n442 B.n87 163.367
R1912 B.n438 B.n87 163.367
R1913 B.n438 B.n437 163.367
R1914 B.n437 B.n436 163.367
R1915 B.n436 B.n89 163.367
R1916 B.n432 B.n89 163.367
R1917 B.n432 B.n431 163.367
R1918 B.n431 B.n430 163.367
R1919 B.n430 B.n91 163.367
R1920 B.n426 B.n91 163.367
R1921 B.n426 B.n425 163.367
R1922 B.n425 B.n424 163.367
R1923 B.n424 B.n93 163.367
R1924 B.n420 B.n93 163.367
R1925 B.n420 B.n419 163.367
R1926 B.n419 B.n418 163.367
R1927 B.n418 B.n95 163.367
R1928 B.n414 B.n95 163.367
R1929 B.n414 B.n413 163.367
R1930 B.n413 B.n412 163.367
R1931 B.n412 B.n97 163.367
R1932 B.n408 B.n97 163.367
R1933 B.n408 B.n407 163.367
R1934 B.n407 B.n406 163.367
R1935 B.n406 B.n99 163.367
R1936 B.n658 B.n11 163.367
R1937 B.n654 B.n11 163.367
R1938 B.n654 B.n653 163.367
R1939 B.n653 B.n652 163.367
R1940 B.n652 B.n13 163.367
R1941 B.n648 B.n13 163.367
R1942 B.n648 B.n647 163.367
R1943 B.n647 B.n646 163.367
R1944 B.n646 B.n15 163.367
R1945 B.n642 B.n15 163.367
R1946 B.n642 B.n641 163.367
R1947 B.n641 B.n640 163.367
R1948 B.n640 B.n17 163.367
R1949 B.n636 B.n17 163.367
R1950 B.n636 B.n635 163.367
R1951 B.n635 B.n634 163.367
R1952 B.n634 B.n19 163.367
R1953 B.n630 B.n19 163.367
R1954 B.n630 B.n629 163.367
R1955 B.n629 B.n628 163.367
R1956 B.n628 B.n21 163.367
R1957 B.n624 B.n21 163.367
R1958 B.n624 B.n623 163.367
R1959 B.n623 B.n622 163.367
R1960 B.n622 B.n23 163.367
R1961 B.n618 B.n23 163.367
R1962 B.n618 B.n617 163.367
R1963 B.n617 B.n616 163.367
R1964 B.n616 B.n25 163.367
R1965 B.n612 B.n25 163.367
R1966 B.n612 B.n611 163.367
R1967 B.n611 B.n610 163.367
R1968 B.n610 B.n27 163.367
R1969 B.n606 B.n27 163.367
R1970 B.n606 B.n605 163.367
R1971 B.n605 B.n604 163.367
R1972 B.n604 B.n29 163.367
R1973 B.n600 B.n29 163.367
R1974 B.n600 B.n599 163.367
R1975 B.n599 B.n598 163.367
R1976 B.n598 B.n31 163.367
R1977 B.n594 B.n31 163.367
R1978 B.n594 B.n593 163.367
R1979 B.n593 B.n592 163.367
R1980 B.n592 B.n33 163.367
R1981 B.n588 B.n33 163.367
R1982 B.n588 B.n587 163.367
R1983 B.n587 B.n586 163.367
R1984 B.n586 B.n35 163.367
R1985 B.n582 B.n35 163.367
R1986 B.n582 B.n581 163.367
R1987 B.n581 B.n580 163.367
R1988 B.n580 B.n37 163.367
R1989 B.n576 B.n37 163.367
R1990 B.n576 B.n575 163.367
R1991 B.n575 B.n574 163.367
R1992 B.n574 B.n39 163.367
R1993 B.n570 B.n39 163.367
R1994 B.n570 B.n569 163.367
R1995 B.n569 B.n568 163.367
R1996 B.n568 B.n41 163.367
R1997 B.n563 B.n41 163.367
R1998 B.n563 B.n562 163.367
R1999 B.n562 B.n561 163.367
R2000 B.n561 B.n45 163.367
R2001 B.n557 B.n45 163.367
R2002 B.n557 B.n556 163.367
R2003 B.n556 B.n555 163.367
R2004 B.n555 B.n47 163.367
R2005 B.n551 B.n47 163.367
R2006 B.n551 B.n550 163.367
R2007 B.n550 B.n51 163.367
R2008 B.n546 B.n51 163.367
R2009 B.n546 B.n545 163.367
R2010 B.n545 B.n544 163.367
R2011 B.n544 B.n53 163.367
R2012 B.n540 B.n53 163.367
R2013 B.n540 B.n539 163.367
R2014 B.n539 B.n538 163.367
R2015 B.n538 B.n55 163.367
R2016 B.n534 B.n55 163.367
R2017 B.n534 B.n533 163.367
R2018 B.n533 B.n532 163.367
R2019 B.n532 B.n57 163.367
R2020 B.n528 B.n57 163.367
R2021 B.n528 B.n527 163.367
R2022 B.n527 B.n526 163.367
R2023 B.n526 B.n59 163.367
R2024 B.n522 B.n59 163.367
R2025 B.n522 B.n521 163.367
R2026 B.n521 B.n520 163.367
R2027 B.n520 B.n61 163.367
R2028 B.n516 B.n61 163.367
R2029 B.n516 B.n515 163.367
R2030 B.n515 B.n514 163.367
R2031 B.n514 B.n63 163.367
R2032 B.n510 B.n63 163.367
R2033 B.n510 B.n509 163.367
R2034 B.n509 B.n508 163.367
R2035 B.n508 B.n65 163.367
R2036 B.n504 B.n65 163.367
R2037 B.n504 B.n503 163.367
R2038 B.n503 B.n502 163.367
R2039 B.n502 B.n67 163.367
R2040 B.n498 B.n67 163.367
R2041 B.n498 B.n497 163.367
R2042 B.n497 B.n496 163.367
R2043 B.n496 B.n69 163.367
R2044 B.n492 B.n69 163.367
R2045 B.n492 B.n491 163.367
R2046 B.n491 B.n490 163.367
R2047 B.n490 B.n71 163.367
R2048 B.n486 B.n71 163.367
R2049 B.n486 B.n485 163.367
R2050 B.n485 B.n484 163.367
R2051 B.n484 B.n73 163.367
R2052 B.n480 B.n73 163.367
R2053 B.n480 B.n479 163.367
R2054 B.n479 B.n478 163.367
R2055 B.n478 B.n75 163.367
R2056 B.n474 B.n75 163.367
R2057 B.n474 B.n473 163.367
R2058 B.n473 B.n472 163.367
R2059 B.n472 B.n77 163.367
R2060 B.n468 B.n77 163.367
R2061 B.n468 B.n467 163.367
R2062 B.n467 B.n466 163.367
R2063 B.n466 B.n79 163.367
R2064 B.n462 B.n79 163.367
R2065 B.n462 B.n461 163.367
R2066 B.n461 B.n460 163.367
R2067 B.n460 B.n81 163.367
R2068 B.n660 B.n659 163.367
R2069 B.n660 B.n9 163.367
R2070 B.n664 B.n9 163.367
R2071 B.n665 B.n664 163.367
R2072 B.n666 B.n665 163.367
R2073 B.n666 B.n7 163.367
R2074 B.n670 B.n7 163.367
R2075 B.n671 B.n670 163.367
R2076 B.n672 B.n671 163.367
R2077 B.n672 B.n5 163.367
R2078 B.n676 B.n5 163.367
R2079 B.n677 B.n676 163.367
R2080 B.n678 B.n677 163.367
R2081 B.n678 B.n3 163.367
R2082 B.n682 B.n3 163.367
R2083 B.n683 B.n682 163.367
R2084 B.n176 B.n2 163.367
R2085 B.n176 B.n175 163.367
R2086 B.n180 B.n175 163.367
R2087 B.n181 B.n180 163.367
R2088 B.n182 B.n181 163.367
R2089 B.n182 B.n173 163.367
R2090 B.n186 B.n173 163.367
R2091 B.n187 B.n186 163.367
R2092 B.n188 B.n187 163.367
R2093 B.n188 B.n171 163.367
R2094 B.n192 B.n171 163.367
R2095 B.n193 B.n192 163.367
R2096 B.n194 B.n193 163.367
R2097 B.n194 B.n169 163.367
R2098 B.n198 B.n169 163.367
R2099 B.n199 B.n198 163.367
R2100 B.n293 B.n137 59.5399
R2101 B.n308 B.n307 59.5399
R2102 B.n50 B.n49 59.5399
R2103 B.n565 B.n43 59.5399
R2104 B.n657 B.n10 34.4981
R2105 B.n458 B.n457 34.4981
R2106 B.n404 B.n403 34.4981
R2107 B.n201 B.n168 34.4981
R2108 B B.n685 18.0485
R2109 B.n661 B.n10 10.6151
R2110 B.n662 B.n661 10.6151
R2111 B.n663 B.n662 10.6151
R2112 B.n663 B.n8 10.6151
R2113 B.n667 B.n8 10.6151
R2114 B.n668 B.n667 10.6151
R2115 B.n669 B.n668 10.6151
R2116 B.n669 B.n6 10.6151
R2117 B.n673 B.n6 10.6151
R2118 B.n674 B.n673 10.6151
R2119 B.n675 B.n674 10.6151
R2120 B.n675 B.n4 10.6151
R2121 B.n679 B.n4 10.6151
R2122 B.n680 B.n679 10.6151
R2123 B.n681 B.n680 10.6151
R2124 B.n681 B.n0 10.6151
R2125 B.n657 B.n656 10.6151
R2126 B.n656 B.n655 10.6151
R2127 B.n655 B.n12 10.6151
R2128 B.n651 B.n12 10.6151
R2129 B.n651 B.n650 10.6151
R2130 B.n650 B.n649 10.6151
R2131 B.n649 B.n14 10.6151
R2132 B.n645 B.n14 10.6151
R2133 B.n645 B.n644 10.6151
R2134 B.n644 B.n643 10.6151
R2135 B.n643 B.n16 10.6151
R2136 B.n639 B.n16 10.6151
R2137 B.n639 B.n638 10.6151
R2138 B.n638 B.n637 10.6151
R2139 B.n637 B.n18 10.6151
R2140 B.n633 B.n18 10.6151
R2141 B.n633 B.n632 10.6151
R2142 B.n632 B.n631 10.6151
R2143 B.n631 B.n20 10.6151
R2144 B.n627 B.n20 10.6151
R2145 B.n627 B.n626 10.6151
R2146 B.n626 B.n625 10.6151
R2147 B.n625 B.n22 10.6151
R2148 B.n621 B.n22 10.6151
R2149 B.n621 B.n620 10.6151
R2150 B.n620 B.n619 10.6151
R2151 B.n619 B.n24 10.6151
R2152 B.n615 B.n24 10.6151
R2153 B.n615 B.n614 10.6151
R2154 B.n614 B.n613 10.6151
R2155 B.n613 B.n26 10.6151
R2156 B.n609 B.n26 10.6151
R2157 B.n609 B.n608 10.6151
R2158 B.n608 B.n607 10.6151
R2159 B.n607 B.n28 10.6151
R2160 B.n603 B.n28 10.6151
R2161 B.n603 B.n602 10.6151
R2162 B.n602 B.n601 10.6151
R2163 B.n601 B.n30 10.6151
R2164 B.n597 B.n30 10.6151
R2165 B.n597 B.n596 10.6151
R2166 B.n596 B.n595 10.6151
R2167 B.n595 B.n32 10.6151
R2168 B.n591 B.n32 10.6151
R2169 B.n591 B.n590 10.6151
R2170 B.n590 B.n589 10.6151
R2171 B.n589 B.n34 10.6151
R2172 B.n585 B.n34 10.6151
R2173 B.n585 B.n584 10.6151
R2174 B.n584 B.n583 10.6151
R2175 B.n583 B.n36 10.6151
R2176 B.n579 B.n36 10.6151
R2177 B.n579 B.n578 10.6151
R2178 B.n578 B.n577 10.6151
R2179 B.n577 B.n38 10.6151
R2180 B.n573 B.n38 10.6151
R2181 B.n573 B.n572 10.6151
R2182 B.n572 B.n571 10.6151
R2183 B.n571 B.n40 10.6151
R2184 B.n567 B.n40 10.6151
R2185 B.n567 B.n566 10.6151
R2186 B.n564 B.n44 10.6151
R2187 B.n560 B.n44 10.6151
R2188 B.n560 B.n559 10.6151
R2189 B.n559 B.n558 10.6151
R2190 B.n558 B.n46 10.6151
R2191 B.n554 B.n46 10.6151
R2192 B.n554 B.n553 10.6151
R2193 B.n553 B.n552 10.6151
R2194 B.n549 B.n548 10.6151
R2195 B.n548 B.n547 10.6151
R2196 B.n547 B.n52 10.6151
R2197 B.n543 B.n52 10.6151
R2198 B.n543 B.n542 10.6151
R2199 B.n542 B.n541 10.6151
R2200 B.n541 B.n54 10.6151
R2201 B.n537 B.n54 10.6151
R2202 B.n537 B.n536 10.6151
R2203 B.n536 B.n535 10.6151
R2204 B.n535 B.n56 10.6151
R2205 B.n531 B.n56 10.6151
R2206 B.n531 B.n530 10.6151
R2207 B.n530 B.n529 10.6151
R2208 B.n529 B.n58 10.6151
R2209 B.n525 B.n58 10.6151
R2210 B.n525 B.n524 10.6151
R2211 B.n524 B.n523 10.6151
R2212 B.n523 B.n60 10.6151
R2213 B.n519 B.n60 10.6151
R2214 B.n519 B.n518 10.6151
R2215 B.n518 B.n517 10.6151
R2216 B.n517 B.n62 10.6151
R2217 B.n513 B.n62 10.6151
R2218 B.n513 B.n512 10.6151
R2219 B.n512 B.n511 10.6151
R2220 B.n511 B.n64 10.6151
R2221 B.n507 B.n64 10.6151
R2222 B.n507 B.n506 10.6151
R2223 B.n506 B.n505 10.6151
R2224 B.n505 B.n66 10.6151
R2225 B.n501 B.n66 10.6151
R2226 B.n501 B.n500 10.6151
R2227 B.n500 B.n499 10.6151
R2228 B.n499 B.n68 10.6151
R2229 B.n495 B.n68 10.6151
R2230 B.n495 B.n494 10.6151
R2231 B.n494 B.n493 10.6151
R2232 B.n493 B.n70 10.6151
R2233 B.n489 B.n70 10.6151
R2234 B.n489 B.n488 10.6151
R2235 B.n488 B.n487 10.6151
R2236 B.n487 B.n72 10.6151
R2237 B.n483 B.n72 10.6151
R2238 B.n483 B.n482 10.6151
R2239 B.n482 B.n481 10.6151
R2240 B.n481 B.n74 10.6151
R2241 B.n477 B.n74 10.6151
R2242 B.n477 B.n476 10.6151
R2243 B.n476 B.n475 10.6151
R2244 B.n475 B.n76 10.6151
R2245 B.n471 B.n76 10.6151
R2246 B.n471 B.n470 10.6151
R2247 B.n470 B.n469 10.6151
R2248 B.n469 B.n78 10.6151
R2249 B.n465 B.n78 10.6151
R2250 B.n465 B.n464 10.6151
R2251 B.n464 B.n463 10.6151
R2252 B.n463 B.n80 10.6151
R2253 B.n459 B.n80 10.6151
R2254 B.n459 B.n458 10.6151
R2255 B.n457 B.n82 10.6151
R2256 B.n453 B.n82 10.6151
R2257 B.n453 B.n452 10.6151
R2258 B.n452 B.n451 10.6151
R2259 B.n451 B.n84 10.6151
R2260 B.n447 B.n84 10.6151
R2261 B.n447 B.n446 10.6151
R2262 B.n446 B.n445 10.6151
R2263 B.n445 B.n86 10.6151
R2264 B.n441 B.n86 10.6151
R2265 B.n441 B.n440 10.6151
R2266 B.n440 B.n439 10.6151
R2267 B.n439 B.n88 10.6151
R2268 B.n435 B.n88 10.6151
R2269 B.n435 B.n434 10.6151
R2270 B.n434 B.n433 10.6151
R2271 B.n433 B.n90 10.6151
R2272 B.n429 B.n90 10.6151
R2273 B.n429 B.n428 10.6151
R2274 B.n428 B.n427 10.6151
R2275 B.n427 B.n92 10.6151
R2276 B.n423 B.n92 10.6151
R2277 B.n423 B.n422 10.6151
R2278 B.n422 B.n421 10.6151
R2279 B.n421 B.n94 10.6151
R2280 B.n417 B.n94 10.6151
R2281 B.n417 B.n416 10.6151
R2282 B.n416 B.n415 10.6151
R2283 B.n415 B.n96 10.6151
R2284 B.n411 B.n96 10.6151
R2285 B.n411 B.n410 10.6151
R2286 B.n410 B.n409 10.6151
R2287 B.n409 B.n98 10.6151
R2288 B.n405 B.n98 10.6151
R2289 B.n405 B.n404 10.6151
R2290 B.n177 B.n1 10.6151
R2291 B.n178 B.n177 10.6151
R2292 B.n179 B.n178 10.6151
R2293 B.n179 B.n174 10.6151
R2294 B.n183 B.n174 10.6151
R2295 B.n184 B.n183 10.6151
R2296 B.n185 B.n184 10.6151
R2297 B.n185 B.n172 10.6151
R2298 B.n189 B.n172 10.6151
R2299 B.n190 B.n189 10.6151
R2300 B.n191 B.n190 10.6151
R2301 B.n191 B.n170 10.6151
R2302 B.n195 B.n170 10.6151
R2303 B.n196 B.n195 10.6151
R2304 B.n197 B.n196 10.6151
R2305 B.n197 B.n168 10.6151
R2306 B.n202 B.n201 10.6151
R2307 B.n203 B.n202 10.6151
R2308 B.n203 B.n166 10.6151
R2309 B.n207 B.n166 10.6151
R2310 B.n208 B.n207 10.6151
R2311 B.n209 B.n208 10.6151
R2312 B.n209 B.n164 10.6151
R2313 B.n213 B.n164 10.6151
R2314 B.n214 B.n213 10.6151
R2315 B.n215 B.n214 10.6151
R2316 B.n215 B.n162 10.6151
R2317 B.n219 B.n162 10.6151
R2318 B.n220 B.n219 10.6151
R2319 B.n221 B.n220 10.6151
R2320 B.n221 B.n160 10.6151
R2321 B.n225 B.n160 10.6151
R2322 B.n226 B.n225 10.6151
R2323 B.n227 B.n226 10.6151
R2324 B.n227 B.n158 10.6151
R2325 B.n231 B.n158 10.6151
R2326 B.n232 B.n231 10.6151
R2327 B.n233 B.n232 10.6151
R2328 B.n233 B.n156 10.6151
R2329 B.n237 B.n156 10.6151
R2330 B.n238 B.n237 10.6151
R2331 B.n239 B.n238 10.6151
R2332 B.n239 B.n154 10.6151
R2333 B.n243 B.n154 10.6151
R2334 B.n244 B.n243 10.6151
R2335 B.n245 B.n244 10.6151
R2336 B.n245 B.n152 10.6151
R2337 B.n249 B.n152 10.6151
R2338 B.n250 B.n249 10.6151
R2339 B.n251 B.n250 10.6151
R2340 B.n251 B.n150 10.6151
R2341 B.n255 B.n150 10.6151
R2342 B.n256 B.n255 10.6151
R2343 B.n257 B.n256 10.6151
R2344 B.n257 B.n148 10.6151
R2345 B.n261 B.n148 10.6151
R2346 B.n262 B.n261 10.6151
R2347 B.n263 B.n262 10.6151
R2348 B.n263 B.n146 10.6151
R2349 B.n267 B.n146 10.6151
R2350 B.n268 B.n267 10.6151
R2351 B.n269 B.n268 10.6151
R2352 B.n269 B.n144 10.6151
R2353 B.n273 B.n144 10.6151
R2354 B.n274 B.n273 10.6151
R2355 B.n275 B.n274 10.6151
R2356 B.n275 B.n142 10.6151
R2357 B.n279 B.n142 10.6151
R2358 B.n280 B.n279 10.6151
R2359 B.n281 B.n280 10.6151
R2360 B.n281 B.n140 10.6151
R2361 B.n285 B.n140 10.6151
R2362 B.n286 B.n285 10.6151
R2363 B.n287 B.n286 10.6151
R2364 B.n287 B.n138 10.6151
R2365 B.n291 B.n138 10.6151
R2366 B.n292 B.n291 10.6151
R2367 B.n294 B.n134 10.6151
R2368 B.n298 B.n134 10.6151
R2369 B.n299 B.n298 10.6151
R2370 B.n300 B.n299 10.6151
R2371 B.n300 B.n132 10.6151
R2372 B.n304 B.n132 10.6151
R2373 B.n305 B.n304 10.6151
R2374 B.n309 B.n305 10.6151
R2375 B.n313 B.n130 10.6151
R2376 B.n314 B.n313 10.6151
R2377 B.n315 B.n314 10.6151
R2378 B.n315 B.n128 10.6151
R2379 B.n319 B.n128 10.6151
R2380 B.n320 B.n319 10.6151
R2381 B.n321 B.n320 10.6151
R2382 B.n321 B.n126 10.6151
R2383 B.n325 B.n126 10.6151
R2384 B.n326 B.n325 10.6151
R2385 B.n327 B.n326 10.6151
R2386 B.n327 B.n124 10.6151
R2387 B.n331 B.n124 10.6151
R2388 B.n332 B.n331 10.6151
R2389 B.n333 B.n332 10.6151
R2390 B.n333 B.n122 10.6151
R2391 B.n337 B.n122 10.6151
R2392 B.n338 B.n337 10.6151
R2393 B.n339 B.n338 10.6151
R2394 B.n339 B.n120 10.6151
R2395 B.n343 B.n120 10.6151
R2396 B.n344 B.n343 10.6151
R2397 B.n345 B.n344 10.6151
R2398 B.n345 B.n118 10.6151
R2399 B.n349 B.n118 10.6151
R2400 B.n350 B.n349 10.6151
R2401 B.n351 B.n350 10.6151
R2402 B.n351 B.n116 10.6151
R2403 B.n355 B.n116 10.6151
R2404 B.n356 B.n355 10.6151
R2405 B.n357 B.n356 10.6151
R2406 B.n357 B.n114 10.6151
R2407 B.n361 B.n114 10.6151
R2408 B.n362 B.n361 10.6151
R2409 B.n363 B.n362 10.6151
R2410 B.n363 B.n112 10.6151
R2411 B.n367 B.n112 10.6151
R2412 B.n368 B.n367 10.6151
R2413 B.n369 B.n368 10.6151
R2414 B.n369 B.n110 10.6151
R2415 B.n373 B.n110 10.6151
R2416 B.n374 B.n373 10.6151
R2417 B.n375 B.n374 10.6151
R2418 B.n375 B.n108 10.6151
R2419 B.n379 B.n108 10.6151
R2420 B.n380 B.n379 10.6151
R2421 B.n381 B.n380 10.6151
R2422 B.n381 B.n106 10.6151
R2423 B.n385 B.n106 10.6151
R2424 B.n386 B.n385 10.6151
R2425 B.n387 B.n386 10.6151
R2426 B.n387 B.n104 10.6151
R2427 B.n391 B.n104 10.6151
R2428 B.n392 B.n391 10.6151
R2429 B.n393 B.n392 10.6151
R2430 B.n393 B.n102 10.6151
R2431 B.n397 B.n102 10.6151
R2432 B.n398 B.n397 10.6151
R2433 B.n399 B.n398 10.6151
R2434 B.n399 B.n100 10.6151
R2435 B.n403 B.n100 10.6151
R2436 B.n137 B.n136 10.2793
R2437 B.n307 B.n306 10.2793
R2438 B.n49 B.n48 10.2793
R2439 B.n43 B.n42 10.2793
R2440 B.n685 B.n0 8.11757
R2441 B.n685 B.n1 8.11757
R2442 B.n565 B.n564 6.5566
R2443 B.n552 B.n50 6.5566
R2444 B.n294 B.n293 6.5566
R2445 B.n309 B.n308 6.5566
R2446 B.n566 B.n565 4.05904
R2447 B.n549 B.n50 4.05904
R2448 B.n293 B.n292 4.05904
R2449 B.n308 B.n130 4.05904
C0 w_n1606_n4750# VDD1 2.32508f
C1 VN VDD1 0.1475f
C2 w_n1606_n4750# VDD2 2.34413f
C3 VN VDD2 4.60493f
C4 VP VTAIL 3.85755f
C5 B VP 1.07482f
C6 B VTAIL 3.4607f
C7 VP VDD1 4.72811f
C8 VP VDD2 0.279016f
C9 VTAIL VDD1 37.8639f
C10 B VDD1 1.95915f
C11 VTAIL VDD2 37.887104f
C12 B VDD2 1.9844f
C13 w_n1606_n4750# VN 2.8416f
C14 VDD1 VDD2 0.666425f
C15 w_n1606_n4750# VP 3.04328f
C16 VP VN 6.14025f
C17 w_n1606_n4750# VTAIL 4.18898f
C18 w_n1606_n4750# B 8.512799f
C19 VN VTAIL 3.84234f
C20 B VN 0.748914f
C21 VDD2 VSUBS 1.792666f
C22 VDD1 VSUBS 1.192799f
C23 VTAIL VSUBS 0.593063f
C24 VN VSUBS 5.31311f
C25 VP VSUBS 1.451569f
C26 B VSUBS 2.968809f
C27 w_n1606_n4750# VSUBS 93.2187f
C28 B.n0 VSUBS 0.006538f
C29 B.n1 VSUBS 0.006538f
C30 B.n2 VSUBS 0.009669f
C31 B.n3 VSUBS 0.00741f
C32 B.n4 VSUBS 0.00741f
C33 B.n5 VSUBS 0.00741f
C34 B.n6 VSUBS 0.00741f
C35 B.n7 VSUBS 0.00741f
C36 B.n8 VSUBS 0.00741f
C37 B.n9 VSUBS 0.00741f
C38 B.n10 VSUBS 0.017767f
C39 B.n11 VSUBS 0.00741f
C40 B.n12 VSUBS 0.00741f
C41 B.n13 VSUBS 0.00741f
C42 B.n14 VSUBS 0.00741f
C43 B.n15 VSUBS 0.00741f
C44 B.n16 VSUBS 0.00741f
C45 B.n17 VSUBS 0.00741f
C46 B.n18 VSUBS 0.00741f
C47 B.n19 VSUBS 0.00741f
C48 B.n20 VSUBS 0.00741f
C49 B.n21 VSUBS 0.00741f
C50 B.n22 VSUBS 0.00741f
C51 B.n23 VSUBS 0.00741f
C52 B.n24 VSUBS 0.00741f
C53 B.n25 VSUBS 0.00741f
C54 B.n26 VSUBS 0.00741f
C55 B.n27 VSUBS 0.00741f
C56 B.n28 VSUBS 0.00741f
C57 B.n29 VSUBS 0.00741f
C58 B.n30 VSUBS 0.00741f
C59 B.n31 VSUBS 0.00741f
C60 B.n32 VSUBS 0.00741f
C61 B.n33 VSUBS 0.00741f
C62 B.n34 VSUBS 0.00741f
C63 B.n35 VSUBS 0.00741f
C64 B.n36 VSUBS 0.00741f
C65 B.n37 VSUBS 0.00741f
C66 B.n38 VSUBS 0.00741f
C67 B.n39 VSUBS 0.00741f
C68 B.n40 VSUBS 0.00741f
C69 B.n41 VSUBS 0.00741f
C70 B.t4 VSUBS 0.395074f
C71 B.t5 VSUBS 0.401886f
C72 B.t3 VSUBS 0.153421f
C73 B.n42 VSUBS 0.389482f
C74 B.n43 VSUBS 0.348814f
C75 B.n44 VSUBS 0.00741f
C76 B.n45 VSUBS 0.00741f
C77 B.n46 VSUBS 0.00741f
C78 B.n47 VSUBS 0.00741f
C79 B.t7 VSUBS 0.395078f
C80 B.t8 VSUBS 0.401889f
C81 B.t6 VSUBS 0.153421f
C82 B.n48 VSUBS 0.389479f
C83 B.n49 VSUBS 0.34881f
C84 B.n50 VSUBS 0.017168f
C85 B.n51 VSUBS 0.00741f
C86 B.n52 VSUBS 0.00741f
C87 B.n53 VSUBS 0.00741f
C88 B.n54 VSUBS 0.00741f
C89 B.n55 VSUBS 0.00741f
C90 B.n56 VSUBS 0.00741f
C91 B.n57 VSUBS 0.00741f
C92 B.n58 VSUBS 0.00741f
C93 B.n59 VSUBS 0.00741f
C94 B.n60 VSUBS 0.00741f
C95 B.n61 VSUBS 0.00741f
C96 B.n62 VSUBS 0.00741f
C97 B.n63 VSUBS 0.00741f
C98 B.n64 VSUBS 0.00741f
C99 B.n65 VSUBS 0.00741f
C100 B.n66 VSUBS 0.00741f
C101 B.n67 VSUBS 0.00741f
C102 B.n68 VSUBS 0.00741f
C103 B.n69 VSUBS 0.00741f
C104 B.n70 VSUBS 0.00741f
C105 B.n71 VSUBS 0.00741f
C106 B.n72 VSUBS 0.00741f
C107 B.n73 VSUBS 0.00741f
C108 B.n74 VSUBS 0.00741f
C109 B.n75 VSUBS 0.00741f
C110 B.n76 VSUBS 0.00741f
C111 B.n77 VSUBS 0.00741f
C112 B.n78 VSUBS 0.00741f
C113 B.n79 VSUBS 0.00741f
C114 B.n80 VSUBS 0.00741f
C115 B.n81 VSUBS 0.018192f
C116 B.n82 VSUBS 0.00741f
C117 B.n83 VSUBS 0.00741f
C118 B.n84 VSUBS 0.00741f
C119 B.n85 VSUBS 0.00741f
C120 B.n86 VSUBS 0.00741f
C121 B.n87 VSUBS 0.00741f
C122 B.n88 VSUBS 0.00741f
C123 B.n89 VSUBS 0.00741f
C124 B.n90 VSUBS 0.00741f
C125 B.n91 VSUBS 0.00741f
C126 B.n92 VSUBS 0.00741f
C127 B.n93 VSUBS 0.00741f
C128 B.n94 VSUBS 0.00741f
C129 B.n95 VSUBS 0.00741f
C130 B.n96 VSUBS 0.00741f
C131 B.n97 VSUBS 0.00741f
C132 B.n98 VSUBS 0.00741f
C133 B.n99 VSUBS 0.017767f
C134 B.n100 VSUBS 0.00741f
C135 B.n101 VSUBS 0.00741f
C136 B.n102 VSUBS 0.00741f
C137 B.n103 VSUBS 0.00741f
C138 B.n104 VSUBS 0.00741f
C139 B.n105 VSUBS 0.00741f
C140 B.n106 VSUBS 0.00741f
C141 B.n107 VSUBS 0.00741f
C142 B.n108 VSUBS 0.00741f
C143 B.n109 VSUBS 0.00741f
C144 B.n110 VSUBS 0.00741f
C145 B.n111 VSUBS 0.00741f
C146 B.n112 VSUBS 0.00741f
C147 B.n113 VSUBS 0.00741f
C148 B.n114 VSUBS 0.00741f
C149 B.n115 VSUBS 0.00741f
C150 B.n116 VSUBS 0.00741f
C151 B.n117 VSUBS 0.00741f
C152 B.n118 VSUBS 0.00741f
C153 B.n119 VSUBS 0.00741f
C154 B.n120 VSUBS 0.00741f
C155 B.n121 VSUBS 0.00741f
C156 B.n122 VSUBS 0.00741f
C157 B.n123 VSUBS 0.00741f
C158 B.n124 VSUBS 0.00741f
C159 B.n125 VSUBS 0.00741f
C160 B.n126 VSUBS 0.00741f
C161 B.n127 VSUBS 0.00741f
C162 B.n128 VSUBS 0.00741f
C163 B.n129 VSUBS 0.00741f
C164 B.n130 VSUBS 0.005121f
C165 B.n131 VSUBS 0.00741f
C166 B.n132 VSUBS 0.00741f
C167 B.n133 VSUBS 0.00741f
C168 B.n134 VSUBS 0.00741f
C169 B.n135 VSUBS 0.00741f
C170 B.t2 VSUBS 0.395074f
C171 B.t1 VSUBS 0.401886f
C172 B.t0 VSUBS 0.153421f
C173 B.n136 VSUBS 0.389482f
C174 B.n137 VSUBS 0.348814f
C175 B.n138 VSUBS 0.00741f
C176 B.n139 VSUBS 0.00741f
C177 B.n140 VSUBS 0.00741f
C178 B.n141 VSUBS 0.00741f
C179 B.n142 VSUBS 0.00741f
C180 B.n143 VSUBS 0.00741f
C181 B.n144 VSUBS 0.00741f
C182 B.n145 VSUBS 0.00741f
C183 B.n146 VSUBS 0.00741f
C184 B.n147 VSUBS 0.00741f
C185 B.n148 VSUBS 0.00741f
C186 B.n149 VSUBS 0.00741f
C187 B.n150 VSUBS 0.00741f
C188 B.n151 VSUBS 0.00741f
C189 B.n152 VSUBS 0.00741f
C190 B.n153 VSUBS 0.00741f
C191 B.n154 VSUBS 0.00741f
C192 B.n155 VSUBS 0.00741f
C193 B.n156 VSUBS 0.00741f
C194 B.n157 VSUBS 0.00741f
C195 B.n158 VSUBS 0.00741f
C196 B.n159 VSUBS 0.00741f
C197 B.n160 VSUBS 0.00741f
C198 B.n161 VSUBS 0.00741f
C199 B.n162 VSUBS 0.00741f
C200 B.n163 VSUBS 0.00741f
C201 B.n164 VSUBS 0.00741f
C202 B.n165 VSUBS 0.00741f
C203 B.n166 VSUBS 0.00741f
C204 B.n167 VSUBS 0.00741f
C205 B.n168 VSUBS 0.017767f
C206 B.n169 VSUBS 0.00741f
C207 B.n170 VSUBS 0.00741f
C208 B.n171 VSUBS 0.00741f
C209 B.n172 VSUBS 0.00741f
C210 B.n173 VSUBS 0.00741f
C211 B.n174 VSUBS 0.00741f
C212 B.n175 VSUBS 0.00741f
C213 B.n176 VSUBS 0.00741f
C214 B.n177 VSUBS 0.00741f
C215 B.n178 VSUBS 0.00741f
C216 B.n179 VSUBS 0.00741f
C217 B.n180 VSUBS 0.00741f
C218 B.n181 VSUBS 0.00741f
C219 B.n182 VSUBS 0.00741f
C220 B.n183 VSUBS 0.00741f
C221 B.n184 VSUBS 0.00741f
C222 B.n185 VSUBS 0.00741f
C223 B.n186 VSUBS 0.00741f
C224 B.n187 VSUBS 0.00741f
C225 B.n188 VSUBS 0.00741f
C226 B.n189 VSUBS 0.00741f
C227 B.n190 VSUBS 0.00741f
C228 B.n191 VSUBS 0.00741f
C229 B.n192 VSUBS 0.00741f
C230 B.n193 VSUBS 0.00741f
C231 B.n194 VSUBS 0.00741f
C232 B.n195 VSUBS 0.00741f
C233 B.n196 VSUBS 0.00741f
C234 B.n197 VSUBS 0.00741f
C235 B.n198 VSUBS 0.00741f
C236 B.n199 VSUBS 0.017767f
C237 B.n200 VSUBS 0.018192f
C238 B.n201 VSUBS 0.018192f
C239 B.n202 VSUBS 0.00741f
C240 B.n203 VSUBS 0.00741f
C241 B.n204 VSUBS 0.00741f
C242 B.n205 VSUBS 0.00741f
C243 B.n206 VSUBS 0.00741f
C244 B.n207 VSUBS 0.00741f
C245 B.n208 VSUBS 0.00741f
C246 B.n209 VSUBS 0.00741f
C247 B.n210 VSUBS 0.00741f
C248 B.n211 VSUBS 0.00741f
C249 B.n212 VSUBS 0.00741f
C250 B.n213 VSUBS 0.00741f
C251 B.n214 VSUBS 0.00741f
C252 B.n215 VSUBS 0.00741f
C253 B.n216 VSUBS 0.00741f
C254 B.n217 VSUBS 0.00741f
C255 B.n218 VSUBS 0.00741f
C256 B.n219 VSUBS 0.00741f
C257 B.n220 VSUBS 0.00741f
C258 B.n221 VSUBS 0.00741f
C259 B.n222 VSUBS 0.00741f
C260 B.n223 VSUBS 0.00741f
C261 B.n224 VSUBS 0.00741f
C262 B.n225 VSUBS 0.00741f
C263 B.n226 VSUBS 0.00741f
C264 B.n227 VSUBS 0.00741f
C265 B.n228 VSUBS 0.00741f
C266 B.n229 VSUBS 0.00741f
C267 B.n230 VSUBS 0.00741f
C268 B.n231 VSUBS 0.00741f
C269 B.n232 VSUBS 0.00741f
C270 B.n233 VSUBS 0.00741f
C271 B.n234 VSUBS 0.00741f
C272 B.n235 VSUBS 0.00741f
C273 B.n236 VSUBS 0.00741f
C274 B.n237 VSUBS 0.00741f
C275 B.n238 VSUBS 0.00741f
C276 B.n239 VSUBS 0.00741f
C277 B.n240 VSUBS 0.00741f
C278 B.n241 VSUBS 0.00741f
C279 B.n242 VSUBS 0.00741f
C280 B.n243 VSUBS 0.00741f
C281 B.n244 VSUBS 0.00741f
C282 B.n245 VSUBS 0.00741f
C283 B.n246 VSUBS 0.00741f
C284 B.n247 VSUBS 0.00741f
C285 B.n248 VSUBS 0.00741f
C286 B.n249 VSUBS 0.00741f
C287 B.n250 VSUBS 0.00741f
C288 B.n251 VSUBS 0.00741f
C289 B.n252 VSUBS 0.00741f
C290 B.n253 VSUBS 0.00741f
C291 B.n254 VSUBS 0.00741f
C292 B.n255 VSUBS 0.00741f
C293 B.n256 VSUBS 0.00741f
C294 B.n257 VSUBS 0.00741f
C295 B.n258 VSUBS 0.00741f
C296 B.n259 VSUBS 0.00741f
C297 B.n260 VSUBS 0.00741f
C298 B.n261 VSUBS 0.00741f
C299 B.n262 VSUBS 0.00741f
C300 B.n263 VSUBS 0.00741f
C301 B.n264 VSUBS 0.00741f
C302 B.n265 VSUBS 0.00741f
C303 B.n266 VSUBS 0.00741f
C304 B.n267 VSUBS 0.00741f
C305 B.n268 VSUBS 0.00741f
C306 B.n269 VSUBS 0.00741f
C307 B.n270 VSUBS 0.00741f
C308 B.n271 VSUBS 0.00741f
C309 B.n272 VSUBS 0.00741f
C310 B.n273 VSUBS 0.00741f
C311 B.n274 VSUBS 0.00741f
C312 B.n275 VSUBS 0.00741f
C313 B.n276 VSUBS 0.00741f
C314 B.n277 VSUBS 0.00741f
C315 B.n278 VSUBS 0.00741f
C316 B.n279 VSUBS 0.00741f
C317 B.n280 VSUBS 0.00741f
C318 B.n281 VSUBS 0.00741f
C319 B.n282 VSUBS 0.00741f
C320 B.n283 VSUBS 0.00741f
C321 B.n284 VSUBS 0.00741f
C322 B.n285 VSUBS 0.00741f
C323 B.n286 VSUBS 0.00741f
C324 B.n287 VSUBS 0.00741f
C325 B.n288 VSUBS 0.00741f
C326 B.n289 VSUBS 0.00741f
C327 B.n290 VSUBS 0.00741f
C328 B.n291 VSUBS 0.00741f
C329 B.n292 VSUBS 0.005121f
C330 B.n293 VSUBS 0.017168f
C331 B.n294 VSUBS 0.005993f
C332 B.n295 VSUBS 0.00741f
C333 B.n296 VSUBS 0.00741f
C334 B.n297 VSUBS 0.00741f
C335 B.n298 VSUBS 0.00741f
C336 B.n299 VSUBS 0.00741f
C337 B.n300 VSUBS 0.00741f
C338 B.n301 VSUBS 0.00741f
C339 B.n302 VSUBS 0.00741f
C340 B.n303 VSUBS 0.00741f
C341 B.n304 VSUBS 0.00741f
C342 B.n305 VSUBS 0.00741f
C343 B.t11 VSUBS 0.395078f
C344 B.t10 VSUBS 0.401889f
C345 B.t9 VSUBS 0.153421f
C346 B.n306 VSUBS 0.389479f
C347 B.n307 VSUBS 0.34881f
C348 B.n308 VSUBS 0.017168f
C349 B.n309 VSUBS 0.005993f
C350 B.n310 VSUBS 0.00741f
C351 B.n311 VSUBS 0.00741f
C352 B.n312 VSUBS 0.00741f
C353 B.n313 VSUBS 0.00741f
C354 B.n314 VSUBS 0.00741f
C355 B.n315 VSUBS 0.00741f
C356 B.n316 VSUBS 0.00741f
C357 B.n317 VSUBS 0.00741f
C358 B.n318 VSUBS 0.00741f
C359 B.n319 VSUBS 0.00741f
C360 B.n320 VSUBS 0.00741f
C361 B.n321 VSUBS 0.00741f
C362 B.n322 VSUBS 0.00741f
C363 B.n323 VSUBS 0.00741f
C364 B.n324 VSUBS 0.00741f
C365 B.n325 VSUBS 0.00741f
C366 B.n326 VSUBS 0.00741f
C367 B.n327 VSUBS 0.00741f
C368 B.n328 VSUBS 0.00741f
C369 B.n329 VSUBS 0.00741f
C370 B.n330 VSUBS 0.00741f
C371 B.n331 VSUBS 0.00741f
C372 B.n332 VSUBS 0.00741f
C373 B.n333 VSUBS 0.00741f
C374 B.n334 VSUBS 0.00741f
C375 B.n335 VSUBS 0.00741f
C376 B.n336 VSUBS 0.00741f
C377 B.n337 VSUBS 0.00741f
C378 B.n338 VSUBS 0.00741f
C379 B.n339 VSUBS 0.00741f
C380 B.n340 VSUBS 0.00741f
C381 B.n341 VSUBS 0.00741f
C382 B.n342 VSUBS 0.00741f
C383 B.n343 VSUBS 0.00741f
C384 B.n344 VSUBS 0.00741f
C385 B.n345 VSUBS 0.00741f
C386 B.n346 VSUBS 0.00741f
C387 B.n347 VSUBS 0.00741f
C388 B.n348 VSUBS 0.00741f
C389 B.n349 VSUBS 0.00741f
C390 B.n350 VSUBS 0.00741f
C391 B.n351 VSUBS 0.00741f
C392 B.n352 VSUBS 0.00741f
C393 B.n353 VSUBS 0.00741f
C394 B.n354 VSUBS 0.00741f
C395 B.n355 VSUBS 0.00741f
C396 B.n356 VSUBS 0.00741f
C397 B.n357 VSUBS 0.00741f
C398 B.n358 VSUBS 0.00741f
C399 B.n359 VSUBS 0.00741f
C400 B.n360 VSUBS 0.00741f
C401 B.n361 VSUBS 0.00741f
C402 B.n362 VSUBS 0.00741f
C403 B.n363 VSUBS 0.00741f
C404 B.n364 VSUBS 0.00741f
C405 B.n365 VSUBS 0.00741f
C406 B.n366 VSUBS 0.00741f
C407 B.n367 VSUBS 0.00741f
C408 B.n368 VSUBS 0.00741f
C409 B.n369 VSUBS 0.00741f
C410 B.n370 VSUBS 0.00741f
C411 B.n371 VSUBS 0.00741f
C412 B.n372 VSUBS 0.00741f
C413 B.n373 VSUBS 0.00741f
C414 B.n374 VSUBS 0.00741f
C415 B.n375 VSUBS 0.00741f
C416 B.n376 VSUBS 0.00741f
C417 B.n377 VSUBS 0.00741f
C418 B.n378 VSUBS 0.00741f
C419 B.n379 VSUBS 0.00741f
C420 B.n380 VSUBS 0.00741f
C421 B.n381 VSUBS 0.00741f
C422 B.n382 VSUBS 0.00741f
C423 B.n383 VSUBS 0.00741f
C424 B.n384 VSUBS 0.00741f
C425 B.n385 VSUBS 0.00741f
C426 B.n386 VSUBS 0.00741f
C427 B.n387 VSUBS 0.00741f
C428 B.n388 VSUBS 0.00741f
C429 B.n389 VSUBS 0.00741f
C430 B.n390 VSUBS 0.00741f
C431 B.n391 VSUBS 0.00741f
C432 B.n392 VSUBS 0.00741f
C433 B.n393 VSUBS 0.00741f
C434 B.n394 VSUBS 0.00741f
C435 B.n395 VSUBS 0.00741f
C436 B.n396 VSUBS 0.00741f
C437 B.n397 VSUBS 0.00741f
C438 B.n398 VSUBS 0.00741f
C439 B.n399 VSUBS 0.00741f
C440 B.n400 VSUBS 0.00741f
C441 B.n401 VSUBS 0.00741f
C442 B.n402 VSUBS 0.018192f
C443 B.n403 VSUBS 0.017363f
C444 B.n404 VSUBS 0.018596f
C445 B.n405 VSUBS 0.00741f
C446 B.n406 VSUBS 0.00741f
C447 B.n407 VSUBS 0.00741f
C448 B.n408 VSUBS 0.00741f
C449 B.n409 VSUBS 0.00741f
C450 B.n410 VSUBS 0.00741f
C451 B.n411 VSUBS 0.00741f
C452 B.n412 VSUBS 0.00741f
C453 B.n413 VSUBS 0.00741f
C454 B.n414 VSUBS 0.00741f
C455 B.n415 VSUBS 0.00741f
C456 B.n416 VSUBS 0.00741f
C457 B.n417 VSUBS 0.00741f
C458 B.n418 VSUBS 0.00741f
C459 B.n419 VSUBS 0.00741f
C460 B.n420 VSUBS 0.00741f
C461 B.n421 VSUBS 0.00741f
C462 B.n422 VSUBS 0.00741f
C463 B.n423 VSUBS 0.00741f
C464 B.n424 VSUBS 0.00741f
C465 B.n425 VSUBS 0.00741f
C466 B.n426 VSUBS 0.00741f
C467 B.n427 VSUBS 0.00741f
C468 B.n428 VSUBS 0.00741f
C469 B.n429 VSUBS 0.00741f
C470 B.n430 VSUBS 0.00741f
C471 B.n431 VSUBS 0.00741f
C472 B.n432 VSUBS 0.00741f
C473 B.n433 VSUBS 0.00741f
C474 B.n434 VSUBS 0.00741f
C475 B.n435 VSUBS 0.00741f
C476 B.n436 VSUBS 0.00741f
C477 B.n437 VSUBS 0.00741f
C478 B.n438 VSUBS 0.00741f
C479 B.n439 VSUBS 0.00741f
C480 B.n440 VSUBS 0.00741f
C481 B.n441 VSUBS 0.00741f
C482 B.n442 VSUBS 0.00741f
C483 B.n443 VSUBS 0.00741f
C484 B.n444 VSUBS 0.00741f
C485 B.n445 VSUBS 0.00741f
C486 B.n446 VSUBS 0.00741f
C487 B.n447 VSUBS 0.00741f
C488 B.n448 VSUBS 0.00741f
C489 B.n449 VSUBS 0.00741f
C490 B.n450 VSUBS 0.00741f
C491 B.n451 VSUBS 0.00741f
C492 B.n452 VSUBS 0.00741f
C493 B.n453 VSUBS 0.00741f
C494 B.n454 VSUBS 0.00741f
C495 B.n455 VSUBS 0.00741f
C496 B.n456 VSUBS 0.017767f
C497 B.n457 VSUBS 0.017767f
C498 B.n458 VSUBS 0.018192f
C499 B.n459 VSUBS 0.00741f
C500 B.n460 VSUBS 0.00741f
C501 B.n461 VSUBS 0.00741f
C502 B.n462 VSUBS 0.00741f
C503 B.n463 VSUBS 0.00741f
C504 B.n464 VSUBS 0.00741f
C505 B.n465 VSUBS 0.00741f
C506 B.n466 VSUBS 0.00741f
C507 B.n467 VSUBS 0.00741f
C508 B.n468 VSUBS 0.00741f
C509 B.n469 VSUBS 0.00741f
C510 B.n470 VSUBS 0.00741f
C511 B.n471 VSUBS 0.00741f
C512 B.n472 VSUBS 0.00741f
C513 B.n473 VSUBS 0.00741f
C514 B.n474 VSUBS 0.00741f
C515 B.n475 VSUBS 0.00741f
C516 B.n476 VSUBS 0.00741f
C517 B.n477 VSUBS 0.00741f
C518 B.n478 VSUBS 0.00741f
C519 B.n479 VSUBS 0.00741f
C520 B.n480 VSUBS 0.00741f
C521 B.n481 VSUBS 0.00741f
C522 B.n482 VSUBS 0.00741f
C523 B.n483 VSUBS 0.00741f
C524 B.n484 VSUBS 0.00741f
C525 B.n485 VSUBS 0.00741f
C526 B.n486 VSUBS 0.00741f
C527 B.n487 VSUBS 0.00741f
C528 B.n488 VSUBS 0.00741f
C529 B.n489 VSUBS 0.00741f
C530 B.n490 VSUBS 0.00741f
C531 B.n491 VSUBS 0.00741f
C532 B.n492 VSUBS 0.00741f
C533 B.n493 VSUBS 0.00741f
C534 B.n494 VSUBS 0.00741f
C535 B.n495 VSUBS 0.00741f
C536 B.n496 VSUBS 0.00741f
C537 B.n497 VSUBS 0.00741f
C538 B.n498 VSUBS 0.00741f
C539 B.n499 VSUBS 0.00741f
C540 B.n500 VSUBS 0.00741f
C541 B.n501 VSUBS 0.00741f
C542 B.n502 VSUBS 0.00741f
C543 B.n503 VSUBS 0.00741f
C544 B.n504 VSUBS 0.00741f
C545 B.n505 VSUBS 0.00741f
C546 B.n506 VSUBS 0.00741f
C547 B.n507 VSUBS 0.00741f
C548 B.n508 VSUBS 0.00741f
C549 B.n509 VSUBS 0.00741f
C550 B.n510 VSUBS 0.00741f
C551 B.n511 VSUBS 0.00741f
C552 B.n512 VSUBS 0.00741f
C553 B.n513 VSUBS 0.00741f
C554 B.n514 VSUBS 0.00741f
C555 B.n515 VSUBS 0.00741f
C556 B.n516 VSUBS 0.00741f
C557 B.n517 VSUBS 0.00741f
C558 B.n518 VSUBS 0.00741f
C559 B.n519 VSUBS 0.00741f
C560 B.n520 VSUBS 0.00741f
C561 B.n521 VSUBS 0.00741f
C562 B.n522 VSUBS 0.00741f
C563 B.n523 VSUBS 0.00741f
C564 B.n524 VSUBS 0.00741f
C565 B.n525 VSUBS 0.00741f
C566 B.n526 VSUBS 0.00741f
C567 B.n527 VSUBS 0.00741f
C568 B.n528 VSUBS 0.00741f
C569 B.n529 VSUBS 0.00741f
C570 B.n530 VSUBS 0.00741f
C571 B.n531 VSUBS 0.00741f
C572 B.n532 VSUBS 0.00741f
C573 B.n533 VSUBS 0.00741f
C574 B.n534 VSUBS 0.00741f
C575 B.n535 VSUBS 0.00741f
C576 B.n536 VSUBS 0.00741f
C577 B.n537 VSUBS 0.00741f
C578 B.n538 VSUBS 0.00741f
C579 B.n539 VSUBS 0.00741f
C580 B.n540 VSUBS 0.00741f
C581 B.n541 VSUBS 0.00741f
C582 B.n542 VSUBS 0.00741f
C583 B.n543 VSUBS 0.00741f
C584 B.n544 VSUBS 0.00741f
C585 B.n545 VSUBS 0.00741f
C586 B.n546 VSUBS 0.00741f
C587 B.n547 VSUBS 0.00741f
C588 B.n548 VSUBS 0.00741f
C589 B.n549 VSUBS 0.005121f
C590 B.n550 VSUBS 0.00741f
C591 B.n551 VSUBS 0.00741f
C592 B.n552 VSUBS 0.005993f
C593 B.n553 VSUBS 0.00741f
C594 B.n554 VSUBS 0.00741f
C595 B.n555 VSUBS 0.00741f
C596 B.n556 VSUBS 0.00741f
C597 B.n557 VSUBS 0.00741f
C598 B.n558 VSUBS 0.00741f
C599 B.n559 VSUBS 0.00741f
C600 B.n560 VSUBS 0.00741f
C601 B.n561 VSUBS 0.00741f
C602 B.n562 VSUBS 0.00741f
C603 B.n563 VSUBS 0.00741f
C604 B.n564 VSUBS 0.005993f
C605 B.n565 VSUBS 0.017168f
C606 B.n566 VSUBS 0.005121f
C607 B.n567 VSUBS 0.00741f
C608 B.n568 VSUBS 0.00741f
C609 B.n569 VSUBS 0.00741f
C610 B.n570 VSUBS 0.00741f
C611 B.n571 VSUBS 0.00741f
C612 B.n572 VSUBS 0.00741f
C613 B.n573 VSUBS 0.00741f
C614 B.n574 VSUBS 0.00741f
C615 B.n575 VSUBS 0.00741f
C616 B.n576 VSUBS 0.00741f
C617 B.n577 VSUBS 0.00741f
C618 B.n578 VSUBS 0.00741f
C619 B.n579 VSUBS 0.00741f
C620 B.n580 VSUBS 0.00741f
C621 B.n581 VSUBS 0.00741f
C622 B.n582 VSUBS 0.00741f
C623 B.n583 VSUBS 0.00741f
C624 B.n584 VSUBS 0.00741f
C625 B.n585 VSUBS 0.00741f
C626 B.n586 VSUBS 0.00741f
C627 B.n587 VSUBS 0.00741f
C628 B.n588 VSUBS 0.00741f
C629 B.n589 VSUBS 0.00741f
C630 B.n590 VSUBS 0.00741f
C631 B.n591 VSUBS 0.00741f
C632 B.n592 VSUBS 0.00741f
C633 B.n593 VSUBS 0.00741f
C634 B.n594 VSUBS 0.00741f
C635 B.n595 VSUBS 0.00741f
C636 B.n596 VSUBS 0.00741f
C637 B.n597 VSUBS 0.00741f
C638 B.n598 VSUBS 0.00741f
C639 B.n599 VSUBS 0.00741f
C640 B.n600 VSUBS 0.00741f
C641 B.n601 VSUBS 0.00741f
C642 B.n602 VSUBS 0.00741f
C643 B.n603 VSUBS 0.00741f
C644 B.n604 VSUBS 0.00741f
C645 B.n605 VSUBS 0.00741f
C646 B.n606 VSUBS 0.00741f
C647 B.n607 VSUBS 0.00741f
C648 B.n608 VSUBS 0.00741f
C649 B.n609 VSUBS 0.00741f
C650 B.n610 VSUBS 0.00741f
C651 B.n611 VSUBS 0.00741f
C652 B.n612 VSUBS 0.00741f
C653 B.n613 VSUBS 0.00741f
C654 B.n614 VSUBS 0.00741f
C655 B.n615 VSUBS 0.00741f
C656 B.n616 VSUBS 0.00741f
C657 B.n617 VSUBS 0.00741f
C658 B.n618 VSUBS 0.00741f
C659 B.n619 VSUBS 0.00741f
C660 B.n620 VSUBS 0.00741f
C661 B.n621 VSUBS 0.00741f
C662 B.n622 VSUBS 0.00741f
C663 B.n623 VSUBS 0.00741f
C664 B.n624 VSUBS 0.00741f
C665 B.n625 VSUBS 0.00741f
C666 B.n626 VSUBS 0.00741f
C667 B.n627 VSUBS 0.00741f
C668 B.n628 VSUBS 0.00741f
C669 B.n629 VSUBS 0.00741f
C670 B.n630 VSUBS 0.00741f
C671 B.n631 VSUBS 0.00741f
C672 B.n632 VSUBS 0.00741f
C673 B.n633 VSUBS 0.00741f
C674 B.n634 VSUBS 0.00741f
C675 B.n635 VSUBS 0.00741f
C676 B.n636 VSUBS 0.00741f
C677 B.n637 VSUBS 0.00741f
C678 B.n638 VSUBS 0.00741f
C679 B.n639 VSUBS 0.00741f
C680 B.n640 VSUBS 0.00741f
C681 B.n641 VSUBS 0.00741f
C682 B.n642 VSUBS 0.00741f
C683 B.n643 VSUBS 0.00741f
C684 B.n644 VSUBS 0.00741f
C685 B.n645 VSUBS 0.00741f
C686 B.n646 VSUBS 0.00741f
C687 B.n647 VSUBS 0.00741f
C688 B.n648 VSUBS 0.00741f
C689 B.n649 VSUBS 0.00741f
C690 B.n650 VSUBS 0.00741f
C691 B.n651 VSUBS 0.00741f
C692 B.n652 VSUBS 0.00741f
C693 B.n653 VSUBS 0.00741f
C694 B.n654 VSUBS 0.00741f
C695 B.n655 VSUBS 0.00741f
C696 B.n656 VSUBS 0.00741f
C697 B.n657 VSUBS 0.018192f
C698 B.n658 VSUBS 0.018192f
C699 B.n659 VSUBS 0.017767f
C700 B.n660 VSUBS 0.00741f
C701 B.n661 VSUBS 0.00741f
C702 B.n662 VSUBS 0.00741f
C703 B.n663 VSUBS 0.00741f
C704 B.n664 VSUBS 0.00741f
C705 B.n665 VSUBS 0.00741f
C706 B.n666 VSUBS 0.00741f
C707 B.n667 VSUBS 0.00741f
C708 B.n668 VSUBS 0.00741f
C709 B.n669 VSUBS 0.00741f
C710 B.n670 VSUBS 0.00741f
C711 B.n671 VSUBS 0.00741f
C712 B.n672 VSUBS 0.00741f
C713 B.n673 VSUBS 0.00741f
C714 B.n674 VSUBS 0.00741f
C715 B.n675 VSUBS 0.00741f
C716 B.n676 VSUBS 0.00741f
C717 B.n677 VSUBS 0.00741f
C718 B.n678 VSUBS 0.00741f
C719 B.n679 VSUBS 0.00741f
C720 B.n680 VSUBS 0.00741f
C721 B.n681 VSUBS 0.00741f
C722 B.n682 VSUBS 0.00741f
C723 B.n683 VSUBS 0.009669f
C724 B.n684 VSUBS 0.0103f
C725 B.n685 VSUBS 0.020483f
C726 VDD1.n0 VSUBS 0.038986f
C727 VDD1.n1 VSUBS 0.035755f
C728 VDD1.n2 VSUBS 0.019213f
C729 VDD1.n3 VSUBS 0.045412f
C730 VDD1.n4 VSUBS 0.020343f
C731 VDD1.n5 VSUBS 0.035755f
C732 VDD1.n6 VSUBS 0.019213f
C733 VDD1.n7 VSUBS 0.045412f
C734 VDD1.n8 VSUBS 0.020343f
C735 VDD1.n9 VSUBS 0.035755f
C736 VDD1.n10 VSUBS 0.019213f
C737 VDD1.n11 VSUBS 0.045412f
C738 VDD1.n12 VSUBS 0.020343f
C739 VDD1.n13 VSUBS 0.035755f
C740 VDD1.n14 VSUBS 0.019213f
C741 VDD1.n15 VSUBS 0.045412f
C742 VDD1.n16 VSUBS 0.045412f
C743 VDD1.n17 VSUBS 0.020343f
C744 VDD1.n18 VSUBS 0.035755f
C745 VDD1.n19 VSUBS 0.019213f
C746 VDD1.n20 VSUBS 0.045412f
C747 VDD1.n21 VSUBS 0.020343f
C748 VDD1.n22 VSUBS 0.035755f
C749 VDD1.n23 VSUBS 0.019213f
C750 VDD1.n24 VSUBS 0.045412f
C751 VDD1.n25 VSUBS 0.020343f
C752 VDD1.n26 VSUBS 0.035755f
C753 VDD1.n27 VSUBS 0.019213f
C754 VDD1.n28 VSUBS 0.045412f
C755 VDD1.n29 VSUBS 0.020343f
C756 VDD1.n30 VSUBS 0.035755f
C757 VDD1.n31 VSUBS 0.019213f
C758 VDD1.n32 VSUBS 0.045412f
C759 VDD1.n33 VSUBS 0.020343f
C760 VDD1.n34 VSUBS 0.293274f
C761 VDD1.t8 VSUBS 0.097567f
C762 VDD1.n35 VSUBS 0.034059f
C763 VDD1.n36 VSUBS 0.028889f
C764 VDD1.n37 VSUBS 0.019213f
C765 VDD1.n38 VSUBS 2.91766f
C766 VDD1.n39 VSUBS 0.035755f
C767 VDD1.n40 VSUBS 0.019213f
C768 VDD1.n41 VSUBS 0.020343f
C769 VDD1.n42 VSUBS 0.045412f
C770 VDD1.n43 VSUBS 0.045412f
C771 VDD1.n44 VSUBS 0.020343f
C772 VDD1.n45 VSUBS 0.019213f
C773 VDD1.n46 VSUBS 0.035755f
C774 VDD1.n47 VSUBS 0.035755f
C775 VDD1.n48 VSUBS 0.019213f
C776 VDD1.n49 VSUBS 0.020343f
C777 VDD1.n50 VSUBS 0.045412f
C778 VDD1.n51 VSUBS 0.045412f
C779 VDD1.n52 VSUBS 0.020343f
C780 VDD1.n53 VSUBS 0.019213f
C781 VDD1.n54 VSUBS 0.035755f
C782 VDD1.n55 VSUBS 0.035755f
C783 VDD1.n56 VSUBS 0.019213f
C784 VDD1.n57 VSUBS 0.020343f
C785 VDD1.n58 VSUBS 0.045412f
C786 VDD1.n59 VSUBS 0.045412f
C787 VDD1.n60 VSUBS 0.020343f
C788 VDD1.n61 VSUBS 0.019213f
C789 VDD1.n62 VSUBS 0.035755f
C790 VDD1.n63 VSUBS 0.035755f
C791 VDD1.n64 VSUBS 0.019213f
C792 VDD1.n65 VSUBS 0.020343f
C793 VDD1.n66 VSUBS 0.045412f
C794 VDD1.n67 VSUBS 0.045412f
C795 VDD1.n68 VSUBS 0.020343f
C796 VDD1.n69 VSUBS 0.019213f
C797 VDD1.n70 VSUBS 0.035755f
C798 VDD1.n71 VSUBS 0.035755f
C799 VDD1.n72 VSUBS 0.019213f
C800 VDD1.n73 VSUBS 0.020343f
C801 VDD1.n74 VSUBS 0.045412f
C802 VDD1.n75 VSUBS 0.045412f
C803 VDD1.n76 VSUBS 0.020343f
C804 VDD1.n77 VSUBS 0.019213f
C805 VDD1.n78 VSUBS 0.035755f
C806 VDD1.n79 VSUBS 0.035755f
C807 VDD1.n80 VSUBS 0.019213f
C808 VDD1.n81 VSUBS 0.019778f
C809 VDD1.n82 VSUBS 0.019778f
C810 VDD1.n83 VSUBS 0.045412f
C811 VDD1.n84 VSUBS 0.045412f
C812 VDD1.n85 VSUBS 0.020343f
C813 VDD1.n86 VSUBS 0.019213f
C814 VDD1.n87 VSUBS 0.035755f
C815 VDD1.n88 VSUBS 0.035755f
C816 VDD1.n89 VSUBS 0.019213f
C817 VDD1.n90 VSUBS 0.020343f
C818 VDD1.n91 VSUBS 0.045412f
C819 VDD1.n92 VSUBS 0.045412f
C820 VDD1.n93 VSUBS 0.020343f
C821 VDD1.n94 VSUBS 0.019213f
C822 VDD1.n95 VSUBS 0.035755f
C823 VDD1.n96 VSUBS 0.035755f
C824 VDD1.n97 VSUBS 0.019213f
C825 VDD1.n98 VSUBS 0.020343f
C826 VDD1.n99 VSUBS 0.045412f
C827 VDD1.n100 VSUBS 0.108913f
C828 VDD1.n101 VSUBS 0.020343f
C829 VDD1.n102 VSUBS 0.019213f
C830 VDD1.n103 VSUBS 0.080203f
C831 VDD1.n104 VSUBS 0.080492f
C832 VDD1.t9 VSUBS 0.53429f
C833 VDD1.t1 VSUBS 0.53429f
C834 VDD1.n105 VSUBS 4.4567f
C835 VDD1.n106 VSUBS 0.909588f
C836 VDD1.n107 VSUBS 0.038986f
C837 VDD1.n108 VSUBS 0.035755f
C838 VDD1.n109 VSUBS 0.019213f
C839 VDD1.n110 VSUBS 0.045412f
C840 VDD1.n111 VSUBS 0.020343f
C841 VDD1.n112 VSUBS 0.035755f
C842 VDD1.n113 VSUBS 0.019213f
C843 VDD1.n114 VSUBS 0.045412f
C844 VDD1.n115 VSUBS 0.020343f
C845 VDD1.n116 VSUBS 0.035755f
C846 VDD1.n117 VSUBS 0.019213f
C847 VDD1.n118 VSUBS 0.045412f
C848 VDD1.n119 VSUBS 0.020343f
C849 VDD1.n120 VSUBS 0.035755f
C850 VDD1.n121 VSUBS 0.019213f
C851 VDD1.n122 VSUBS 0.045412f
C852 VDD1.n123 VSUBS 0.020343f
C853 VDD1.n124 VSUBS 0.035755f
C854 VDD1.n125 VSUBS 0.019213f
C855 VDD1.n126 VSUBS 0.045412f
C856 VDD1.n127 VSUBS 0.020343f
C857 VDD1.n128 VSUBS 0.035755f
C858 VDD1.n129 VSUBS 0.019213f
C859 VDD1.n130 VSUBS 0.045412f
C860 VDD1.n131 VSUBS 0.020343f
C861 VDD1.n132 VSUBS 0.035755f
C862 VDD1.n133 VSUBS 0.019213f
C863 VDD1.n134 VSUBS 0.045412f
C864 VDD1.n135 VSUBS 0.020343f
C865 VDD1.n136 VSUBS 0.035755f
C866 VDD1.n137 VSUBS 0.019213f
C867 VDD1.n138 VSUBS 0.045412f
C868 VDD1.n139 VSUBS 0.020343f
C869 VDD1.n140 VSUBS 0.293274f
C870 VDD1.t4 VSUBS 0.097567f
C871 VDD1.n141 VSUBS 0.034059f
C872 VDD1.n142 VSUBS 0.028889f
C873 VDD1.n143 VSUBS 0.019213f
C874 VDD1.n144 VSUBS 2.91766f
C875 VDD1.n145 VSUBS 0.035755f
C876 VDD1.n146 VSUBS 0.019213f
C877 VDD1.n147 VSUBS 0.020343f
C878 VDD1.n148 VSUBS 0.045412f
C879 VDD1.n149 VSUBS 0.045412f
C880 VDD1.n150 VSUBS 0.020343f
C881 VDD1.n151 VSUBS 0.019213f
C882 VDD1.n152 VSUBS 0.035755f
C883 VDD1.n153 VSUBS 0.035755f
C884 VDD1.n154 VSUBS 0.019213f
C885 VDD1.n155 VSUBS 0.020343f
C886 VDD1.n156 VSUBS 0.045412f
C887 VDD1.n157 VSUBS 0.045412f
C888 VDD1.n158 VSUBS 0.020343f
C889 VDD1.n159 VSUBS 0.019213f
C890 VDD1.n160 VSUBS 0.035755f
C891 VDD1.n161 VSUBS 0.035755f
C892 VDD1.n162 VSUBS 0.019213f
C893 VDD1.n163 VSUBS 0.020343f
C894 VDD1.n164 VSUBS 0.045412f
C895 VDD1.n165 VSUBS 0.045412f
C896 VDD1.n166 VSUBS 0.020343f
C897 VDD1.n167 VSUBS 0.019213f
C898 VDD1.n168 VSUBS 0.035755f
C899 VDD1.n169 VSUBS 0.035755f
C900 VDD1.n170 VSUBS 0.019213f
C901 VDD1.n171 VSUBS 0.020343f
C902 VDD1.n172 VSUBS 0.045412f
C903 VDD1.n173 VSUBS 0.045412f
C904 VDD1.n174 VSUBS 0.020343f
C905 VDD1.n175 VSUBS 0.019213f
C906 VDD1.n176 VSUBS 0.035755f
C907 VDD1.n177 VSUBS 0.035755f
C908 VDD1.n178 VSUBS 0.019213f
C909 VDD1.n179 VSUBS 0.020343f
C910 VDD1.n180 VSUBS 0.045412f
C911 VDD1.n181 VSUBS 0.045412f
C912 VDD1.n182 VSUBS 0.045412f
C913 VDD1.n183 VSUBS 0.020343f
C914 VDD1.n184 VSUBS 0.019213f
C915 VDD1.n185 VSUBS 0.035755f
C916 VDD1.n186 VSUBS 0.035755f
C917 VDD1.n187 VSUBS 0.019213f
C918 VDD1.n188 VSUBS 0.019778f
C919 VDD1.n189 VSUBS 0.019778f
C920 VDD1.n190 VSUBS 0.045412f
C921 VDD1.n191 VSUBS 0.045412f
C922 VDD1.n192 VSUBS 0.020343f
C923 VDD1.n193 VSUBS 0.019213f
C924 VDD1.n194 VSUBS 0.035755f
C925 VDD1.n195 VSUBS 0.035755f
C926 VDD1.n196 VSUBS 0.019213f
C927 VDD1.n197 VSUBS 0.020343f
C928 VDD1.n198 VSUBS 0.045412f
C929 VDD1.n199 VSUBS 0.045412f
C930 VDD1.n200 VSUBS 0.020343f
C931 VDD1.n201 VSUBS 0.019213f
C932 VDD1.n202 VSUBS 0.035755f
C933 VDD1.n203 VSUBS 0.035755f
C934 VDD1.n204 VSUBS 0.019213f
C935 VDD1.n205 VSUBS 0.020343f
C936 VDD1.n206 VSUBS 0.045412f
C937 VDD1.n207 VSUBS 0.108913f
C938 VDD1.n208 VSUBS 0.020343f
C939 VDD1.n209 VSUBS 0.019213f
C940 VDD1.n210 VSUBS 0.080203f
C941 VDD1.n211 VSUBS 0.080492f
C942 VDD1.t5 VSUBS 0.53429f
C943 VDD1.t2 VSUBS 0.53429f
C944 VDD1.n212 VSUBS 4.45669f
C945 VDD1.n213 VSUBS 0.910598f
C946 VDD1.t0 VSUBS 0.53429f
C947 VDD1.t3 VSUBS 0.53429f
C948 VDD1.n214 VSUBS 4.46017f
C949 VDD1.n215 VSUBS 3.46f
C950 VDD1.t6 VSUBS 0.53429f
C951 VDD1.t7 VSUBS 0.53429f
C952 VDD1.n216 VSUBS 4.45668f
C953 VDD1.n217 VSUBS 4.30248f
C954 VP.n0 VSUBS 0.070511f
C955 VP.t9 VSUBS 0.75143f
C956 VP.t7 VSUBS 0.75143f
C957 VP.t4 VSUBS 0.75143f
C958 VP.n1 VSUBS 0.28811f
C959 VP.n2 VSUBS 0.070511f
C960 VP.t3 VSUBS 0.75143f
C961 VP.t8 VSUBS 0.75143f
C962 VP.t0 VSUBS 0.75143f
C963 VP.n3 VSUBS 0.28811f
C964 VP.t1 VSUBS 0.756694f
C965 VP.n4 VSUBS 0.308074f
C966 VP.n5 VSUBS 0.154835f
C967 VP.n6 VSUBS 0.024695f
C968 VP.n7 VSUBS 0.28811f
C969 VP.n8 VSUBS 0.024695f
C970 VP.n9 VSUBS 0.28811f
C971 VP.t2 VSUBS 0.756694f
C972 VP.n10 VSUBS 0.307975f
C973 VP.n11 VSUBS 3.29927f
C974 VP.t5 VSUBS 0.756694f
C975 VP.n12 VSUBS 0.307975f
C976 VP.n13 VSUBS 3.35514f
C977 VP.n14 VSUBS 0.070511f
C978 VP.n15 VSUBS 0.024695f
C979 VP.n16 VSUBS 0.28811f
C980 VP.n17 VSUBS 0.024695f
C981 VP.n18 VSUBS 0.28811f
C982 VP.t6 VSUBS 0.756694f
C983 VP.n19 VSUBS 0.307975f
C984 VP.n20 VSUBS 0.054644f
C985 VDD2.n0 VSUBS 0.039014f
C986 VDD2.n1 VSUBS 0.03578f
C987 VDD2.n2 VSUBS 0.019227f
C988 VDD2.n3 VSUBS 0.045445f
C989 VDD2.n4 VSUBS 0.020358f
C990 VDD2.n5 VSUBS 0.03578f
C991 VDD2.n6 VSUBS 0.019227f
C992 VDD2.n7 VSUBS 0.045445f
C993 VDD2.n8 VSUBS 0.020358f
C994 VDD2.n9 VSUBS 0.03578f
C995 VDD2.n10 VSUBS 0.019227f
C996 VDD2.n11 VSUBS 0.045445f
C997 VDD2.n12 VSUBS 0.020358f
C998 VDD2.n13 VSUBS 0.03578f
C999 VDD2.n14 VSUBS 0.019227f
C1000 VDD2.n15 VSUBS 0.045445f
C1001 VDD2.n16 VSUBS 0.020358f
C1002 VDD2.n17 VSUBS 0.03578f
C1003 VDD2.n18 VSUBS 0.019227f
C1004 VDD2.n19 VSUBS 0.045445f
C1005 VDD2.n20 VSUBS 0.020358f
C1006 VDD2.n21 VSUBS 0.03578f
C1007 VDD2.n22 VSUBS 0.019227f
C1008 VDD2.n23 VSUBS 0.045445f
C1009 VDD2.n24 VSUBS 0.020358f
C1010 VDD2.n25 VSUBS 0.03578f
C1011 VDD2.n26 VSUBS 0.019227f
C1012 VDD2.n27 VSUBS 0.045445f
C1013 VDD2.n28 VSUBS 0.020358f
C1014 VDD2.n29 VSUBS 0.03578f
C1015 VDD2.n30 VSUBS 0.019227f
C1016 VDD2.n31 VSUBS 0.045445f
C1017 VDD2.n32 VSUBS 0.020358f
C1018 VDD2.n33 VSUBS 0.293484f
C1019 VDD2.t8 VSUBS 0.097636f
C1020 VDD2.n34 VSUBS 0.034084f
C1021 VDD2.n35 VSUBS 0.02891f
C1022 VDD2.n36 VSUBS 0.019227f
C1023 VDD2.n37 VSUBS 2.91975f
C1024 VDD2.n38 VSUBS 0.03578f
C1025 VDD2.n39 VSUBS 0.019227f
C1026 VDD2.n40 VSUBS 0.020358f
C1027 VDD2.n41 VSUBS 0.045445f
C1028 VDD2.n42 VSUBS 0.045445f
C1029 VDD2.n43 VSUBS 0.020358f
C1030 VDD2.n44 VSUBS 0.019227f
C1031 VDD2.n45 VSUBS 0.03578f
C1032 VDD2.n46 VSUBS 0.03578f
C1033 VDD2.n47 VSUBS 0.019227f
C1034 VDD2.n48 VSUBS 0.020358f
C1035 VDD2.n49 VSUBS 0.045445f
C1036 VDD2.n50 VSUBS 0.045445f
C1037 VDD2.n51 VSUBS 0.020358f
C1038 VDD2.n52 VSUBS 0.019227f
C1039 VDD2.n53 VSUBS 0.03578f
C1040 VDD2.n54 VSUBS 0.03578f
C1041 VDD2.n55 VSUBS 0.019227f
C1042 VDD2.n56 VSUBS 0.020358f
C1043 VDD2.n57 VSUBS 0.045445f
C1044 VDD2.n58 VSUBS 0.045445f
C1045 VDD2.n59 VSUBS 0.020358f
C1046 VDD2.n60 VSUBS 0.019227f
C1047 VDD2.n61 VSUBS 0.03578f
C1048 VDD2.n62 VSUBS 0.03578f
C1049 VDD2.n63 VSUBS 0.019227f
C1050 VDD2.n64 VSUBS 0.020358f
C1051 VDD2.n65 VSUBS 0.045445f
C1052 VDD2.n66 VSUBS 0.045445f
C1053 VDD2.n67 VSUBS 0.020358f
C1054 VDD2.n68 VSUBS 0.019227f
C1055 VDD2.n69 VSUBS 0.03578f
C1056 VDD2.n70 VSUBS 0.03578f
C1057 VDD2.n71 VSUBS 0.019227f
C1058 VDD2.n72 VSUBS 0.020358f
C1059 VDD2.n73 VSUBS 0.045445f
C1060 VDD2.n74 VSUBS 0.045445f
C1061 VDD2.n75 VSUBS 0.045445f
C1062 VDD2.n76 VSUBS 0.020358f
C1063 VDD2.n77 VSUBS 0.019227f
C1064 VDD2.n78 VSUBS 0.03578f
C1065 VDD2.n79 VSUBS 0.03578f
C1066 VDD2.n80 VSUBS 0.019227f
C1067 VDD2.n81 VSUBS 0.019792f
C1068 VDD2.n82 VSUBS 0.019792f
C1069 VDD2.n83 VSUBS 0.045445f
C1070 VDD2.n84 VSUBS 0.045445f
C1071 VDD2.n85 VSUBS 0.020358f
C1072 VDD2.n86 VSUBS 0.019227f
C1073 VDD2.n87 VSUBS 0.03578f
C1074 VDD2.n88 VSUBS 0.03578f
C1075 VDD2.n89 VSUBS 0.019227f
C1076 VDD2.n90 VSUBS 0.020358f
C1077 VDD2.n91 VSUBS 0.045445f
C1078 VDD2.n92 VSUBS 0.045445f
C1079 VDD2.n93 VSUBS 0.020358f
C1080 VDD2.n94 VSUBS 0.019227f
C1081 VDD2.n95 VSUBS 0.03578f
C1082 VDD2.n96 VSUBS 0.03578f
C1083 VDD2.n97 VSUBS 0.019227f
C1084 VDD2.n98 VSUBS 0.020358f
C1085 VDD2.n99 VSUBS 0.045445f
C1086 VDD2.n100 VSUBS 0.108991f
C1087 VDD2.n101 VSUBS 0.020358f
C1088 VDD2.n102 VSUBS 0.019227f
C1089 VDD2.n103 VSUBS 0.08026f
C1090 VDD2.n104 VSUBS 0.08055f
C1091 VDD2.t6 VSUBS 0.534673f
C1092 VDD2.t9 VSUBS 0.534673f
C1093 VDD2.n105 VSUBS 4.45988f
C1094 VDD2.n106 VSUBS 0.91125f
C1095 VDD2.t7 VSUBS 0.534673f
C1096 VDD2.t4 VSUBS 0.534673f
C1097 VDD2.n107 VSUBS 4.46337f
C1098 VDD2.n108 VSUBS 3.36754f
C1099 VDD2.n109 VSUBS 0.039014f
C1100 VDD2.n110 VSUBS 0.03578f
C1101 VDD2.n111 VSUBS 0.019227f
C1102 VDD2.n112 VSUBS 0.045445f
C1103 VDD2.n113 VSUBS 0.020358f
C1104 VDD2.n114 VSUBS 0.03578f
C1105 VDD2.n115 VSUBS 0.019227f
C1106 VDD2.n116 VSUBS 0.045445f
C1107 VDD2.n117 VSUBS 0.020358f
C1108 VDD2.n118 VSUBS 0.03578f
C1109 VDD2.n119 VSUBS 0.019227f
C1110 VDD2.n120 VSUBS 0.045445f
C1111 VDD2.n121 VSUBS 0.020358f
C1112 VDD2.n122 VSUBS 0.03578f
C1113 VDD2.n123 VSUBS 0.019227f
C1114 VDD2.n124 VSUBS 0.045445f
C1115 VDD2.n125 VSUBS 0.045445f
C1116 VDD2.n126 VSUBS 0.020358f
C1117 VDD2.n127 VSUBS 0.03578f
C1118 VDD2.n128 VSUBS 0.019227f
C1119 VDD2.n129 VSUBS 0.045445f
C1120 VDD2.n130 VSUBS 0.020358f
C1121 VDD2.n131 VSUBS 0.03578f
C1122 VDD2.n132 VSUBS 0.019227f
C1123 VDD2.n133 VSUBS 0.045445f
C1124 VDD2.n134 VSUBS 0.020358f
C1125 VDD2.n135 VSUBS 0.03578f
C1126 VDD2.n136 VSUBS 0.019227f
C1127 VDD2.n137 VSUBS 0.045445f
C1128 VDD2.n138 VSUBS 0.020358f
C1129 VDD2.n139 VSUBS 0.03578f
C1130 VDD2.n140 VSUBS 0.019227f
C1131 VDD2.n141 VSUBS 0.045445f
C1132 VDD2.n142 VSUBS 0.020358f
C1133 VDD2.n143 VSUBS 0.293484f
C1134 VDD2.t2 VSUBS 0.097636f
C1135 VDD2.n144 VSUBS 0.034084f
C1136 VDD2.n145 VSUBS 0.02891f
C1137 VDD2.n146 VSUBS 0.019227f
C1138 VDD2.n147 VSUBS 2.91975f
C1139 VDD2.n148 VSUBS 0.03578f
C1140 VDD2.n149 VSUBS 0.019227f
C1141 VDD2.n150 VSUBS 0.020358f
C1142 VDD2.n151 VSUBS 0.045445f
C1143 VDD2.n152 VSUBS 0.045445f
C1144 VDD2.n153 VSUBS 0.020358f
C1145 VDD2.n154 VSUBS 0.019227f
C1146 VDD2.n155 VSUBS 0.03578f
C1147 VDD2.n156 VSUBS 0.03578f
C1148 VDD2.n157 VSUBS 0.019227f
C1149 VDD2.n158 VSUBS 0.020358f
C1150 VDD2.n159 VSUBS 0.045445f
C1151 VDD2.n160 VSUBS 0.045445f
C1152 VDD2.n161 VSUBS 0.020358f
C1153 VDD2.n162 VSUBS 0.019227f
C1154 VDD2.n163 VSUBS 0.03578f
C1155 VDD2.n164 VSUBS 0.03578f
C1156 VDD2.n165 VSUBS 0.019227f
C1157 VDD2.n166 VSUBS 0.020358f
C1158 VDD2.n167 VSUBS 0.045445f
C1159 VDD2.n168 VSUBS 0.045445f
C1160 VDD2.n169 VSUBS 0.020358f
C1161 VDD2.n170 VSUBS 0.019227f
C1162 VDD2.n171 VSUBS 0.03578f
C1163 VDD2.n172 VSUBS 0.03578f
C1164 VDD2.n173 VSUBS 0.019227f
C1165 VDD2.n174 VSUBS 0.020358f
C1166 VDD2.n175 VSUBS 0.045445f
C1167 VDD2.n176 VSUBS 0.045445f
C1168 VDD2.n177 VSUBS 0.020358f
C1169 VDD2.n178 VSUBS 0.019227f
C1170 VDD2.n179 VSUBS 0.03578f
C1171 VDD2.n180 VSUBS 0.03578f
C1172 VDD2.n181 VSUBS 0.019227f
C1173 VDD2.n182 VSUBS 0.020358f
C1174 VDD2.n183 VSUBS 0.045445f
C1175 VDD2.n184 VSUBS 0.045445f
C1176 VDD2.n185 VSUBS 0.020358f
C1177 VDD2.n186 VSUBS 0.019227f
C1178 VDD2.n187 VSUBS 0.03578f
C1179 VDD2.n188 VSUBS 0.03578f
C1180 VDD2.n189 VSUBS 0.019227f
C1181 VDD2.n190 VSUBS 0.019792f
C1182 VDD2.n191 VSUBS 0.019792f
C1183 VDD2.n192 VSUBS 0.045445f
C1184 VDD2.n193 VSUBS 0.045445f
C1185 VDD2.n194 VSUBS 0.020358f
C1186 VDD2.n195 VSUBS 0.019227f
C1187 VDD2.n196 VSUBS 0.03578f
C1188 VDD2.n197 VSUBS 0.03578f
C1189 VDD2.n198 VSUBS 0.019227f
C1190 VDD2.n199 VSUBS 0.020358f
C1191 VDD2.n200 VSUBS 0.045445f
C1192 VDD2.n201 VSUBS 0.045445f
C1193 VDD2.n202 VSUBS 0.020358f
C1194 VDD2.n203 VSUBS 0.019227f
C1195 VDD2.n204 VSUBS 0.03578f
C1196 VDD2.n205 VSUBS 0.03578f
C1197 VDD2.n206 VSUBS 0.019227f
C1198 VDD2.n207 VSUBS 0.020358f
C1199 VDD2.n208 VSUBS 0.045445f
C1200 VDD2.n209 VSUBS 0.108991f
C1201 VDD2.n210 VSUBS 0.020358f
C1202 VDD2.n211 VSUBS 0.019227f
C1203 VDD2.n212 VSUBS 0.08026f
C1204 VDD2.n213 VSUBS 0.079415f
C1205 VDD2.n214 VSUBS 3.56998f
C1206 VDD2.t1 VSUBS 0.534673f
C1207 VDD2.t0 VSUBS 0.534673f
C1208 VDD2.n215 VSUBS 4.45989f
C1209 VDD2.n216 VSUBS 0.7912f
C1210 VDD2.t5 VSUBS 0.534673f
C1211 VDD2.t3 VSUBS 0.534673f
C1212 VDD2.n217 VSUBS 4.46331f
C1213 VTAIL.t16 VSUBS 0.561199f
C1214 VTAIL.t11 VSUBS 0.561199f
C1215 VTAIL.n0 VSUBS 4.43552f
C1216 VTAIL.n1 VSUBS 1.08189f
C1217 VTAIL.n2 VSUBS 0.040949f
C1218 VTAIL.n3 VSUBS 0.037555f
C1219 VTAIL.n4 VSUBS 0.020181f
C1220 VTAIL.n5 VSUBS 0.0477f
C1221 VTAIL.n6 VSUBS 0.021368f
C1222 VTAIL.n7 VSUBS 0.037555f
C1223 VTAIL.n8 VSUBS 0.020181f
C1224 VTAIL.n9 VSUBS 0.0477f
C1225 VTAIL.n10 VSUBS 0.021368f
C1226 VTAIL.n11 VSUBS 0.037555f
C1227 VTAIL.n12 VSUBS 0.020181f
C1228 VTAIL.n13 VSUBS 0.0477f
C1229 VTAIL.n14 VSUBS 0.021368f
C1230 VTAIL.n15 VSUBS 0.037555f
C1231 VTAIL.n16 VSUBS 0.020181f
C1232 VTAIL.n17 VSUBS 0.0477f
C1233 VTAIL.n18 VSUBS 0.021368f
C1234 VTAIL.n19 VSUBS 0.037555f
C1235 VTAIL.n20 VSUBS 0.020181f
C1236 VTAIL.n21 VSUBS 0.0477f
C1237 VTAIL.n22 VSUBS 0.021368f
C1238 VTAIL.n23 VSUBS 0.037555f
C1239 VTAIL.n24 VSUBS 0.020181f
C1240 VTAIL.n25 VSUBS 0.0477f
C1241 VTAIL.n26 VSUBS 0.021368f
C1242 VTAIL.n27 VSUBS 0.037555f
C1243 VTAIL.n28 VSUBS 0.020181f
C1244 VTAIL.n29 VSUBS 0.0477f
C1245 VTAIL.n30 VSUBS 0.021368f
C1246 VTAIL.n31 VSUBS 0.037555f
C1247 VTAIL.n32 VSUBS 0.020181f
C1248 VTAIL.n33 VSUBS 0.0477f
C1249 VTAIL.n34 VSUBS 0.021368f
C1250 VTAIL.n35 VSUBS 0.308044f
C1251 VTAIL.t1 VSUBS 0.10248f
C1252 VTAIL.n36 VSUBS 0.035775f
C1253 VTAIL.n37 VSUBS 0.030344f
C1254 VTAIL.n38 VSUBS 0.020181f
C1255 VTAIL.n39 VSUBS 3.0646f
C1256 VTAIL.n40 VSUBS 0.037555f
C1257 VTAIL.n41 VSUBS 0.020181f
C1258 VTAIL.n42 VSUBS 0.021368f
C1259 VTAIL.n43 VSUBS 0.0477f
C1260 VTAIL.n44 VSUBS 0.0477f
C1261 VTAIL.n45 VSUBS 0.021368f
C1262 VTAIL.n46 VSUBS 0.020181f
C1263 VTAIL.n47 VSUBS 0.037555f
C1264 VTAIL.n48 VSUBS 0.037555f
C1265 VTAIL.n49 VSUBS 0.020181f
C1266 VTAIL.n50 VSUBS 0.021368f
C1267 VTAIL.n51 VSUBS 0.0477f
C1268 VTAIL.n52 VSUBS 0.0477f
C1269 VTAIL.n53 VSUBS 0.021368f
C1270 VTAIL.n54 VSUBS 0.020181f
C1271 VTAIL.n55 VSUBS 0.037555f
C1272 VTAIL.n56 VSUBS 0.037555f
C1273 VTAIL.n57 VSUBS 0.020181f
C1274 VTAIL.n58 VSUBS 0.021368f
C1275 VTAIL.n59 VSUBS 0.0477f
C1276 VTAIL.n60 VSUBS 0.0477f
C1277 VTAIL.n61 VSUBS 0.021368f
C1278 VTAIL.n62 VSUBS 0.020181f
C1279 VTAIL.n63 VSUBS 0.037555f
C1280 VTAIL.n64 VSUBS 0.037555f
C1281 VTAIL.n65 VSUBS 0.020181f
C1282 VTAIL.n66 VSUBS 0.021368f
C1283 VTAIL.n67 VSUBS 0.0477f
C1284 VTAIL.n68 VSUBS 0.0477f
C1285 VTAIL.n69 VSUBS 0.021368f
C1286 VTAIL.n70 VSUBS 0.020181f
C1287 VTAIL.n71 VSUBS 0.037555f
C1288 VTAIL.n72 VSUBS 0.037555f
C1289 VTAIL.n73 VSUBS 0.020181f
C1290 VTAIL.n74 VSUBS 0.021368f
C1291 VTAIL.n75 VSUBS 0.0477f
C1292 VTAIL.n76 VSUBS 0.0477f
C1293 VTAIL.n77 VSUBS 0.0477f
C1294 VTAIL.n78 VSUBS 0.021368f
C1295 VTAIL.n79 VSUBS 0.020181f
C1296 VTAIL.n80 VSUBS 0.037555f
C1297 VTAIL.n81 VSUBS 0.037555f
C1298 VTAIL.n82 VSUBS 0.020181f
C1299 VTAIL.n83 VSUBS 0.020774f
C1300 VTAIL.n84 VSUBS 0.020774f
C1301 VTAIL.n85 VSUBS 0.0477f
C1302 VTAIL.n86 VSUBS 0.0477f
C1303 VTAIL.n87 VSUBS 0.021368f
C1304 VTAIL.n88 VSUBS 0.020181f
C1305 VTAIL.n89 VSUBS 0.037555f
C1306 VTAIL.n90 VSUBS 0.037555f
C1307 VTAIL.n91 VSUBS 0.020181f
C1308 VTAIL.n92 VSUBS 0.021368f
C1309 VTAIL.n93 VSUBS 0.0477f
C1310 VTAIL.n94 VSUBS 0.0477f
C1311 VTAIL.n95 VSUBS 0.021368f
C1312 VTAIL.n96 VSUBS 0.020181f
C1313 VTAIL.n97 VSUBS 0.037555f
C1314 VTAIL.n98 VSUBS 0.037555f
C1315 VTAIL.n99 VSUBS 0.020181f
C1316 VTAIL.n100 VSUBS 0.021368f
C1317 VTAIL.n101 VSUBS 0.0477f
C1318 VTAIL.n102 VSUBS 0.114398f
C1319 VTAIL.n103 VSUBS 0.021368f
C1320 VTAIL.n104 VSUBS 0.020181f
C1321 VTAIL.n105 VSUBS 0.084242f
C1322 VTAIL.n106 VSUBS 0.057402f
C1323 VTAIL.n107 VSUBS 0.170418f
C1324 VTAIL.t4 VSUBS 0.561199f
C1325 VTAIL.t3 VSUBS 0.561199f
C1326 VTAIL.n108 VSUBS 4.43552f
C1327 VTAIL.n109 VSUBS 1.05947f
C1328 VTAIL.t8 VSUBS 0.561199f
C1329 VTAIL.t0 VSUBS 0.561199f
C1330 VTAIL.n110 VSUBS 4.43552f
C1331 VTAIL.n111 VSUBS 3.5976f
C1332 VTAIL.t15 VSUBS 0.561199f
C1333 VTAIL.t14 VSUBS 0.561199f
C1334 VTAIL.n112 VSUBS 4.43554f
C1335 VTAIL.n113 VSUBS 3.59758f
C1336 VTAIL.t13 VSUBS 0.561199f
C1337 VTAIL.t12 VSUBS 0.561199f
C1338 VTAIL.n114 VSUBS 4.43554f
C1339 VTAIL.n115 VSUBS 1.05945f
C1340 VTAIL.n116 VSUBS 0.040949f
C1341 VTAIL.n117 VSUBS 0.037555f
C1342 VTAIL.n118 VSUBS 0.020181f
C1343 VTAIL.n119 VSUBS 0.0477f
C1344 VTAIL.n120 VSUBS 0.021368f
C1345 VTAIL.n121 VSUBS 0.037555f
C1346 VTAIL.n122 VSUBS 0.020181f
C1347 VTAIL.n123 VSUBS 0.0477f
C1348 VTAIL.n124 VSUBS 0.021368f
C1349 VTAIL.n125 VSUBS 0.037555f
C1350 VTAIL.n126 VSUBS 0.020181f
C1351 VTAIL.n127 VSUBS 0.0477f
C1352 VTAIL.n128 VSUBS 0.021368f
C1353 VTAIL.n129 VSUBS 0.037555f
C1354 VTAIL.n130 VSUBS 0.020181f
C1355 VTAIL.n131 VSUBS 0.0477f
C1356 VTAIL.n132 VSUBS 0.0477f
C1357 VTAIL.n133 VSUBS 0.021368f
C1358 VTAIL.n134 VSUBS 0.037555f
C1359 VTAIL.n135 VSUBS 0.020181f
C1360 VTAIL.n136 VSUBS 0.0477f
C1361 VTAIL.n137 VSUBS 0.021368f
C1362 VTAIL.n138 VSUBS 0.037555f
C1363 VTAIL.n139 VSUBS 0.020181f
C1364 VTAIL.n140 VSUBS 0.0477f
C1365 VTAIL.n141 VSUBS 0.021368f
C1366 VTAIL.n142 VSUBS 0.037555f
C1367 VTAIL.n143 VSUBS 0.020181f
C1368 VTAIL.n144 VSUBS 0.0477f
C1369 VTAIL.n145 VSUBS 0.021368f
C1370 VTAIL.n146 VSUBS 0.037555f
C1371 VTAIL.n147 VSUBS 0.020181f
C1372 VTAIL.n148 VSUBS 0.0477f
C1373 VTAIL.n149 VSUBS 0.021368f
C1374 VTAIL.n150 VSUBS 0.308044f
C1375 VTAIL.t18 VSUBS 0.10248f
C1376 VTAIL.n151 VSUBS 0.035775f
C1377 VTAIL.n152 VSUBS 0.030344f
C1378 VTAIL.n153 VSUBS 0.020181f
C1379 VTAIL.n154 VSUBS 3.0646f
C1380 VTAIL.n155 VSUBS 0.037555f
C1381 VTAIL.n156 VSUBS 0.020181f
C1382 VTAIL.n157 VSUBS 0.021368f
C1383 VTAIL.n158 VSUBS 0.0477f
C1384 VTAIL.n159 VSUBS 0.0477f
C1385 VTAIL.n160 VSUBS 0.021368f
C1386 VTAIL.n161 VSUBS 0.020181f
C1387 VTAIL.n162 VSUBS 0.037555f
C1388 VTAIL.n163 VSUBS 0.037555f
C1389 VTAIL.n164 VSUBS 0.020181f
C1390 VTAIL.n165 VSUBS 0.021368f
C1391 VTAIL.n166 VSUBS 0.0477f
C1392 VTAIL.n167 VSUBS 0.0477f
C1393 VTAIL.n168 VSUBS 0.021368f
C1394 VTAIL.n169 VSUBS 0.020181f
C1395 VTAIL.n170 VSUBS 0.037555f
C1396 VTAIL.n171 VSUBS 0.037555f
C1397 VTAIL.n172 VSUBS 0.020181f
C1398 VTAIL.n173 VSUBS 0.021368f
C1399 VTAIL.n174 VSUBS 0.0477f
C1400 VTAIL.n175 VSUBS 0.0477f
C1401 VTAIL.n176 VSUBS 0.021368f
C1402 VTAIL.n177 VSUBS 0.020181f
C1403 VTAIL.n178 VSUBS 0.037555f
C1404 VTAIL.n179 VSUBS 0.037555f
C1405 VTAIL.n180 VSUBS 0.020181f
C1406 VTAIL.n181 VSUBS 0.021368f
C1407 VTAIL.n182 VSUBS 0.0477f
C1408 VTAIL.n183 VSUBS 0.0477f
C1409 VTAIL.n184 VSUBS 0.021368f
C1410 VTAIL.n185 VSUBS 0.020181f
C1411 VTAIL.n186 VSUBS 0.037555f
C1412 VTAIL.n187 VSUBS 0.037555f
C1413 VTAIL.n188 VSUBS 0.020181f
C1414 VTAIL.n189 VSUBS 0.021368f
C1415 VTAIL.n190 VSUBS 0.0477f
C1416 VTAIL.n191 VSUBS 0.0477f
C1417 VTAIL.n192 VSUBS 0.021368f
C1418 VTAIL.n193 VSUBS 0.020181f
C1419 VTAIL.n194 VSUBS 0.037555f
C1420 VTAIL.n195 VSUBS 0.037555f
C1421 VTAIL.n196 VSUBS 0.020181f
C1422 VTAIL.n197 VSUBS 0.020774f
C1423 VTAIL.n198 VSUBS 0.020774f
C1424 VTAIL.n199 VSUBS 0.0477f
C1425 VTAIL.n200 VSUBS 0.0477f
C1426 VTAIL.n201 VSUBS 0.021368f
C1427 VTAIL.n202 VSUBS 0.020181f
C1428 VTAIL.n203 VSUBS 0.037555f
C1429 VTAIL.n204 VSUBS 0.037555f
C1430 VTAIL.n205 VSUBS 0.020181f
C1431 VTAIL.n206 VSUBS 0.021368f
C1432 VTAIL.n207 VSUBS 0.0477f
C1433 VTAIL.n208 VSUBS 0.0477f
C1434 VTAIL.n209 VSUBS 0.021368f
C1435 VTAIL.n210 VSUBS 0.020181f
C1436 VTAIL.n211 VSUBS 0.037555f
C1437 VTAIL.n212 VSUBS 0.037555f
C1438 VTAIL.n213 VSUBS 0.020181f
C1439 VTAIL.n214 VSUBS 0.021368f
C1440 VTAIL.n215 VSUBS 0.0477f
C1441 VTAIL.n216 VSUBS 0.114398f
C1442 VTAIL.n217 VSUBS 0.021368f
C1443 VTAIL.n218 VSUBS 0.020181f
C1444 VTAIL.n219 VSUBS 0.084242f
C1445 VTAIL.n220 VSUBS 0.057402f
C1446 VTAIL.n221 VSUBS 0.170418f
C1447 VTAIL.t7 VSUBS 0.561199f
C1448 VTAIL.t2 VSUBS 0.561199f
C1449 VTAIL.n222 VSUBS 4.43554f
C1450 VTAIL.n223 VSUBS 1.08866f
C1451 VTAIL.t5 VSUBS 0.561199f
C1452 VTAIL.t6 VSUBS 0.561199f
C1453 VTAIL.n224 VSUBS 4.43554f
C1454 VTAIL.n225 VSUBS 1.05945f
C1455 VTAIL.n226 VSUBS 0.040949f
C1456 VTAIL.n227 VSUBS 0.037555f
C1457 VTAIL.n228 VSUBS 0.020181f
C1458 VTAIL.n229 VSUBS 0.0477f
C1459 VTAIL.n230 VSUBS 0.021368f
C1460 VTAIL.n231 VSUBS 0.037555f
C1461 VTAIL.n232 VSUBS 0.020181f
C1462 VTAIL.n233 VSUBS 0.0477f
C1463 VTAIL.n234 VSUBS 0.021368f
C1464 VTAIL.n235 VSUBS 0.037555f
C1465 VTAIL.n236 VSUBS 0.020181f
C1466 VTAIL.n237 VSUBS 0.0477f
C1467 VTAIL.n238 VSUBS 0.021368f
C1468 VTAIL.n239 VSUBS 0.037555f
C1469 VTAIL.n240 VSUBS 0.020181f
C1470 VTAIL.n241 VSUBS 0.0477f
C1471 VTAIL.n242 VSUBS 0.0477f
C1472 VTAIL.n243 VSUBS 0.021368f
C1473 VTAIL.n244 VSUBS 0.037555f
C1474 VTAIL.n245 VSUBS 0.020181f
C1475 VTAIL.n246 VSUBS 0.0477f
C1476 VTAIL.n247 VSUBS 0.021368f
C1477 VTAIL.n248 VSUBS 0.037555f
C1478 VTAIL.n249 VSUBS 0.020181f
C1479 VTAIL.n250 VSUBS 0.0477f
C1480 VTAIL.n251 VSUBS 0.021368f
C1481 VTAIL.n252 VSUBS 0.037555f
C1482 VTAIL.n253 VSUBS 0.020181f
C1483 VTAIL.n254 VSUBS 0.0477f
C1484 VTAIL.n255 VSUBS 0.021368f
C1485 VTAIL.n256 VSUBS 0.037555f
C1486 VTAIL.n257 VSUBS 0.020181f
C1487 VTAIL.n258 VSUBS 0.0477f
C1488 VTAIL.n259 VSUBS 0.021368f
C1489 VTAIL.n260 VSUBS 0.308044f
C1490 VTAIL.t9 VSUBS 0.10248f
C1491 VTAIL.n261 VSUBS 0.035775f
C1492 VTAIL.n262 VSUBS 0.030344f
C1493 VTAIL.n263 VSUBS 0.020181f
C1494 VTAIL.n264 VSUBS 3.0646f
C1495 VTAIL.n265 VSUBS 0.037555f
C1496 VTAIL.n266 VSUBS 0.020181f
C1497 VTAIL.n267 VSUBS 0.021368f
C1498 VTAIL.n268 VSUBS 0.0477f
C1499 VTAIL.n269 VSUBS 0.0477f
C1500 VTAIL.n270 VSUBS 0.021368f
C1501 VTAIL.n271 VSUBS 0.020181f
C1502 VTAIL.n272 VSUBS 0.037555f
C1503 VTAIL.n273 VSUBS 0.037555f
C1504 VTAIL.n274 VSUBS 0.020181f
C1505 VTAIL.n275 VSUBS 0.021368f
C1506 VTAIL.n276 VSUBS 0.0477f
C1507 VTAIL.n277 VSUBS 0.0477f
C1508 VTAIL.n278 VSUBS 0.021368f
C1509 VTAIL.n279 VSUBS 0.020181f
C1510 VTAIL.n280 VSUBS 0.037555f
C1511 VTAIL.n281 VSUBS 0.037555f
C1512 VTAIL.n282 VSUBS 0.020181f
C1513 VTAIL.n283 VSUBS 0.021368f
C1514 VTAIL.n284 VSUBS 0.0477f
C1515 VTAIL.n285 VSUBS 0.0477f
C1516 VTAIL.n286 VSUBS 0.021368f
C1517 VTAIL.n287 VSUBS 0.020181f
C1518 VTAIL.n288 VSUBS 0.037555f
C1519 VTAIL.n289 VSUBS 0.037555f
C1520 VTAIL.n290 VSUBS 0.020181f
C1521 VTAIL.n291 VSUBS 0.021368f
C1522 VTAIL.n292 VSUBS 0.0477f
C1523 VTAIL.n293 VSUBS 0.0477f
C1524 VTAIL.n294 VSUBS 0.021368f
C1525 VTAIL.n295 VSUBS 0.020181f
C1526 VTAIL.n296 VSUBS 0.037555f
C1527 VTAIL.n297 VSUBS 0.037555f
C1528 VTAIL.n298 VSUBS 0.020181f
C1529 VTAIL.n299 VSUBS 0.021368f
C1530 VTAIL.n300 VSUBS 0.0477f
C1531 VTAIL.n301 VSUBS 0.0477f
C1532 VTAIL.n302 VSUBS 0.021368f
C1533 VTAIL.n303 VSUBS 0.020181f
C1534 VTAIL.n304 VSUBS 0.037555f
C1535 VTAIL.n305 VSUBS 0.037555f
C1536 VTAIL.n306 VSUBS 0.020181f
C1537 VTAIL.n307 VSUBS 0.020774f
C1538 VTAIL.n308 VSUBS 0.020774f
C1539 VTAIL.n309 VSUBS 0.0477f
C1540 VTAIL.n310 VSUBS 0.0477f
C1541 VTAIL.n311 VSUBS 0.021368f
C1542 VTAIL.n312 VSUBS 0.020181f
C1543 VTAIL.n313 VSUBS 0.037555f
C1544 VTAIL.n314 VSUBS 0.037555f
C1545 VTAIL.n315 VSUBS 0.020181f
C1546 VTAIL.n316 VSUBS 0.021368f
C1547 VTAIL.n317 VSUBS 0.0477f
C1548 VTAIL.n318 VSUBS 0.0477f
C1549 VTAIL.n319 VSUBS 0.021368f
C1550 VTAIL.n320 VSUBS 0.020181f
C1551 VTAIL.n321 VSUBS 0.037555f
C1552 VTAIL.n322 VSUBS 0.037555f
C1553 VTAIL.n323 VSUBS 0.020181f
C1554 VTAIL.n324 VSUBS 0.021368f
C1555 VTAIL.n325 VSUBS 0.0477f
C1556 VTAIL.n326 VSUBS 0.114398f
C1557 VTAIL.n327 VSUBS 0.021368f
C1558 VTAIL.n328 VSUBS 0.020181f
C1559 VTAIL.n329 VSUBS 0.084242f
C1560 VTAIL.n330 VSUBS 0.057402f
C1561 VTAIL.n331 VSUBS 2.62405f
C1562 VTAIL.n332 VSUBS 0.040949f
C1563 VTAIL.n333 VSUBS 0.037555f
C1564 VTAIL.n334 VSUBS 0.020181f
C1565 VTAIL.n335 VSUBS 0.0477f
C1566 VTAIL.n336 VSUBS 0.021368f
C1567 VTAIL.n337 VSUBS 0.037555f
C1568 VTAIL.n338 VSUBS 0.020181f
C1569 VTAIL.n339 VSUBS 0.0477f
C1570 VTAIL.n340 VSUBS 0.021368f
C1571 VTAIL.n341 VSUBS 0.037555f
C1572 VTAIL.n342 VSUBS 0.020181f
C1573 VTAIL.n343 VSUBS 0.0477f
C1574 VTAIL.n344 VSUBS 0.021368f
C1575 VTAIL.n345 VSUBS 0.037555f
C1576 VTAIL.n346 VSUBS 0.020181f
C1577 VTAIL.n347 VSUBS 0.0477f
C1578 VTAIL.n348 VSUBS 0.021368f
C1579 VTAIL.n349 VSUBS 0.037555f
C1580 VTAIL.n350 VSUBS 0.020181f
C1581 VTAIL.n351 VSUBS 0.0477f
C1582 VTAIL.n352 VSUBS 0.021368f
C1583 VTAIL.n353 VSUBS 0.037555f
C1584 VTAIL.n354 VSUBS 0.020181f
C1585 VTAIL.n355 VSUBS 0.0477f
C1586 VTAIL.n356 VSUBS 0.021368f
C1587 VTAIL.n357 VSUBS 0.037555f
C1588 VTAIL.n358 VSUBS 0.020181f
C1589 VTAIL.n359 VSUBS 0.0477f
C1590 VTAIL.n360 VSUBS 0.021368f
C1591 VTAIL.n361 VSUBS 0.037555f
C1592 VTAIL.n362 VSUBS 0.020181f
C1593 VTAIL.n363 VSUBS 0.0477f
C1594 VTAIL.n364 VSUBS 0.021368f
C1595 VTAIL.n365 VSUBS 0.308044f
C1596 VTAIL.t10 VSUBS 0.10248f
C1597 VTAIL.n366 VSUBS 0.035775f
C1598 VTAIL.n367 VSUBS 0.030344f
C1599 VTAIL.n368 VSUBS 0.020181f
C1600 VTAIL.n369 VSUBS 3.0646f
C1601 VTAIL.n370 VSUBS 0.037555f
C1602 VTAIL.n371 VSUBS 0.020181f
C1603 VTAIL.n372 VSUBS 0.021368f
C1604 VTAIL.n373 VSUBS 0.0477f
C1605 VTAIL.n374 VSUBS 0.0477f
C1606 VTAIL.n375 VSUBS 0.021368f
C1607 VTAIL.n376 VSUBS 0.020181f
C1608 VTAIL.n377 VSUBS 0.037555f
C1609 VTAIL.n378 VSUBS 0.037555f
C1610 VTAIL.n379 VSUBS 0.020181f
C1611 VTAIL.n380 VSUBS 0.021368f
C1612 VTAIL.n381 VSUBS 0.0477f
C1613 VTAIL.n382 VSUBS 0.0477f
C1614 VTAIL.n383 VSUBS 0.021368f
C1615 VTAIL.n384 VSUBS 0.020181f
C1616 VTAIL.n385 VSUBS 0.037555f
C1617 VTAIL.n386 VSUBS 0.037555f
C1618 VTAIL.n387 VSUBS 0.020181f
C1619 VTAIL.n388 VSUBS 0.021368f
C1620 VTAIL.n389 VSUBS 0.0477f
C1621 VTAIL.n390 VSUBS 0.0477f
C1622 VTAIL.n391 VSUBS 0.021368f
C1623 VTAIL.n392 VSUBS 0.020181f
C1624 VTAIL.n393 VSUBS 0.037555f
C1625 VTAIL.n394 VSUBS 0.037555f
C1626 VTAIL.n395 VSUBS 0.020181f
C1627 VTAIL.n396 VSUBS 0.021368f
C1628 VTAIL.n397 VSUBS 0.0477f
C1629 VTAIL.n398 VSUBS 0.0477f
C1630 VTAIL.n399 VSUBS 0.021368f
C1631 VTAIL.n400 VSUBS 0.020181f
C1632 VTAIL.n401 VSUBS 0.037555f
C1633 VTAIL.n402 VSUBS 0.037555f
C1634 VTAIL.n403 VSUBS 0.020181f
C1635 VTAIL.n404 VSUBS 0.021368f
C1636 VTAIL.n405 VSUBS 0.0477f
C1637 VTAIL.n406 VSUBS 0.0477f
C1638 VTAIL.n407 VSUBS 0.0477f
C1639 VTAIL.n408 VSUBS 0.021368f
C1640 VTAIL.n409 VSUBS 0.020181f
C1641 VTAIL.n410 VSUBS 0.037555f
C1642 VTAIL.n411 VSUBS 0.037555f
C1643 VTAIL.n412 VSUBS 0.020181f
C1644 VTAIL.n413 VSUBS 0.020774f
C1645 VTAIL.n414 VSUBS 0.020774f
C1646 VTAIL.n415 VSUBS 0.0477f
C1647 VTAIL.n416 VSUBS 0.0477f
C1648 VTAIL.n417 VSUBS 0.021368f
C1649 VTAIL.n418 VSUBS 0.020181f
C1650 VTAIL.n419 VSUBS 0.037555f
C1651 VTAIL.n420 VSUBS 0.037555f
C1652 VTAIL.n421 VSUBS 0.020181f
C1653 VTAIL.n422 VSUBS 0.021368f
C1654 VTAIL.n423 VSUBS 0.0477f
C1655 VTAIL.n424 VSUBS 0.0477f
C1656 VTAIL.n425 VSUBS 0.021368f
C1657 VTAIL.n426 VSUBS 0.020181f
C1658 VTAIL.n427 VSUBS 0.037555f
C1659 VTAIL.n428 VSUBS 0.037555f
C1660 VTAIL.n429 VSUBS 0.020181f
C1661 VTAIL.n430 VSUBS 0.021368f
C1662 VTAIL.n431 VSUBS 0.0477f
C1663 VTAIL.n432 VSUBS 0.114398f
C1664 VTAIL.n433 VSUBS 0.021368f
C1665 VTAIL.n434 VSUBS 0.020181f
C1666 VTAIL.n435 VSUBS 0.084242f
C1667 VTAIL.n436 VSUBS 0.057402f
C1668 VTAIL.n437 VSUBS 2.62405f
C1669 VTAIL.t19 VSUBS 0.561199f
C1670 VTAIL.t17 VSUBS 0.561199f
C1671 VTAIL.n438 VSUBS 4.43552f
C1672 VTAIL.n439 VSUBS 1.01096f
C1673 VN.n0 VSUBS 0.068534f
C1674 VN.t2 VSUBS 0.730359f
C1675 VN.t0 VSUBS 0.730359f
C1676 VN.t3 VSUBS 0.730359f
C1677 VN.n1 VSUBS 0.280031f
C1678 VN.t1 VSUBS 0.735475f
C1679 VN.n2 VSUBS 0.299435f
C1680 VN.n3 VSUBS 0.150493f
C1681 VN.n4 VSUBS 0.024003f
C1682 VN.n5 VSUBS 0.280031f
C1683 VN.n6 VSUBS 0.024003f
C1684 VN.n7 VSUBS 0.280031f
C1685 VN.t5 VSUBS 0.735475f
C1686 VN.n8 VSUBS 0.299339f
C1687 VN.n9 VSUBS 0.053111f
C1688 VN.n10 VSUBS 0.068534f
C1689 VN.t7 VSUBS 0.735475f
C1690 VN.t8 VSUBS 0.730359f
C1691 VN.t9 VSUBS 0.730359f
C1692 VN.t4 VSUBS 0.730359f
C1693 VN.n11 VSUBS 0.280031f
C1694 VN.t6 VSUBS 0.735475f
C1695 VN.n12 VSUBS 0.299435f
C1696 VN.n13 VSUBS 0.150493f
C1697 VN.n14 VSUBS 0.024003f
C1698 VN.n15 VSUBS 0.280031f
C1699 VN.n16 VSUBS 0.024003f
C1700 VN.n17 VSUBS 0.280031f
C1701 VN.n18 VSUBS 0.299339f
C1702 VN.n19 VSUBS 3.25154f
.ends

