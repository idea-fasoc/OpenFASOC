* NGSPICE file created from diff_pair_sample_1681.ext - technology: sky130A

.subckt diff_pair_sample_1681 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=5.8149 pd=30.6 as=5.8149 ps=30.6 w=14.91 l=1.03
X1 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.8149 pd=30.6 as=5.8149 ps=30.6 w=14.91 l=1.03
X2 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=5.8149 pd=30.6 as=0 ps=0 w=14.91 l=1.03
X3 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=5.8149 pd=30.6 as=0 ps=0 w=14.91 l=1.03
X4 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.8149 pd=30.6 as=5.8149 ps=30.6 w=14.91 l=1.03
X5 VDD1.t0 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=5.8149 pd=30.6 as=5.8149 ps=30.6 w=14.91 l=1.03
X6 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=5.8149 pd=30.6 as=0 ps=0 w=14.91 l=1.03
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=5.8149 pd=30.6 as=0 ps=0 w=14.91 l=1.03
R0 VP.n0 VP.t1 591.25
R1 VP.n0 VP.t0 548.538
R2 VP VP.n0 0.0516364
R3 VTAIL.n322 VTAIL.n246 289.615
R4 VTAIL.n76 VTAIL.n0 289.615
R5 VTAIL.n240 VTAIL.n164 289.615
R6 VTAIL.n158 VTAIL.n82 289.615
R7 VTAIL.n273 VTAIL.n272 185
R8 VTAIL.n270 VTAIL.n269 185
R9 VTAIL.n279 VTAIL.n278 185
R10 VTAIL.n281 VTAIL.n280 185
R11 VTAIL.n266 VTAIL.n265 185
R12 VTAIL.n287 VTAIL.n286 185
R13 VTAIL.n290 VTAIL.n289 185
R14 VTAIL.n288 VTAIL.n262 185
R15 VTAIL.n295 VTAIL.n261 185
R16 VTAIL.n297 VTAIL.n296 185
R17 VTAIL.n299 VTAIL.n298 185
R18 VTAIL.n258 VTAIL.n257 185
R19 VTAIL.n305 VTAIL.n304 185
R20 VTAIL.n307 VTAIL.n306 185
R21 VTAIL.n254 VTAIL.n253 185
R22 VTAIL.n313 VTAIL.n312 185
R23 VTAIL.n315 VTAIL.n314 185
R24 VTAIL.n250 VTAIL.n249 185
R25 VTAIL.n321 VTAIL.n320 185
R26 VTAIL.n323 VTAIL.n322 185
R27 VTAIL.n27 VTAIL.n26 185
R28 VTAIL.n24 VTAIL.n23 185
R29 VTAIL.n33 VTAIL.n32 185
R30 VTAIL.n35 VTAIL.n34 185
R31 VTAIL.n20 VTAIL.n19 185
R32 VTAIL.n41 VTAIL.n40 185
R33 VTAIL.n44 VTAIL.n43 185
R34 VTAIL.n42 VTAIL.n16 185
R35 VTAIL.n49 VTAIL.n15 185
R36 VTAIL.n51 VTAIL.n50 185
R37 VTAIL.n53 VTAIL.n52 185
R38 VTAIL.n12 VTAIL.n11 185
R39 VTAIL.n59 VTAIL.n58 185
R40 VTAIL.n61 VTAIL.n60 185
R41 VTAIL.n8 VTAIL.n7 185
R42 VTAIL.n67 VTAIL.n66 185
R43 VTAIL.n69 VTAIL.n68 185
R44 VTAIL.n4 VTAIL.n3 185
R45 VTAIL.n75 VTAIL.n74 185
R46 VTAIL.n77 VTAIL.n76 185
R47 VTAIL.n241 VTAIL.n240 185
R48 VTAIL.n239 VTAIL.n238 185
R49 VTAIL.n168 VTAIL.n167 185
R50 VTAIL.n233 VTAIL.n232 185
R51 VTAIL.n231 VTAIL.n230 185
R52 VTAIL.n172 VTAIL.n171 185
R53 VTAIL.n225 VTAIL.n224 185
R54 VTAIL.n223 VTAIL.n222 185
R55 VTAIL.n176 VTAIL.n175 185
R56 VTAIL.n217 VTAIL.n216 185
R57 VTAIL.n215 VTAIL.n214 185
R58 VTAIL.n213 VTAIL.n179 185
R59 VTAIL.n183 VTAIL.n180 185
R60 VTAIL.n208 VTAIL.n207 185
R61 VTAIL.n206 VTAIL.n205 185
R62 VTAIL.n185 VTAIL.n184 185
R63 VTAIL.n200 VTAIL.n199 185
R64 VTAIL.n198 VTAIL.n197 185
R65 VTAIL.n189 VTAIL.n188 185
R66 VTAIL.n192 VTAIL.n191 185
R67 VTAIL.n159 VTAIL.n158 185
R68 VTAIL.n157 VTAIL.n156 185
R69 VTAIL.n86 VTAIL.n85 185
R70 VTAIL.n151 VTAIL.n150 185
R71 VTAIL.n149 VTAIL.n148 185
R72 VTAIL.n90 VTAIL.n89 185
R73 VTAIL.n143 VTAIL.n142 185
R74 VTAIL.n141 VTAIL.n140 185
R75 VTAIL.n94 VTAIL.n93 185
R76 VTAIL.n135 VTAIL.n134 185
R77 VTAIL.n133 VTAIL.n132 185
R78 VTAIL.n131 VTAIL.n97 185
R79 VTAIL.n101 VTAIL.n98 185
R80 VTAIL.n126 VTAIL.n125 185
R81 VTAIL.n124 VTAIL.n123 185
R82 VTAIL.n103 VTAIL.n102 185
R83 VTAIL.n118 VTAIL.n117 185
R84 VTAIL.n116 VTAIL.n115 185
R85 VTAIL.n107 VTAIL.n106 185
R86 VTAIL.n110 VTAIL.n109 185
R87 VTAIL.t1 VTAIL.n271 149.524
R88 VTAIL.t2 VTAIL.n25 149.524
R89 VTAIL.t3 VTAIL.n190 149.524
R90 VTAIL.t0 VTAIL.n108 149.524
R91 VTAIL.n272 VTAIL.n269 104.615
R92 VTAIL.n279 VTAIL.n269 104.615
R93 VTAIL.n280 VTAIL.n279 104.615
R94 VTAIL.n280 VTAIL.n265 104.615
R95 VTAIL.n287 VTAIL.n265 104.615
R96 VTAIL.n289 VTAIL.n287 104.615
R97 VTAIL.n289 VTAIL.n288 104.615
R98 VTAIL.n288 VTAIL.n261 104.615
R99 VTAIL.n297 VTAIL.n261 104.615
R100 VTAIL.n298 VTAIL.n297 104.615
R101 VTAIL.n298 VTAIL.n257 104.615
R102 VTAIL.n305 VTAIL.n257 104.615
R103 VTAIL.n306 VTAIL.n305 104.615
R104 VTAIL.n306 VTAIL.n253 104.615
R105 VTAIL.n313 VTAIL.n253 104.615
R106 VTAIL.n314 VTAIL.n313 104.615
R107 VTAIL.n314 VTAIL.n249 104.615
R108 VTAIL.n321 VTAIL.n249 104.615
R109 VTAIL.n322 VTAIL.n321 104.615
R110 VTAIL.n26 VTAIL.n23 104.615
R111 VTAIL.n33 VTAIL.n23 104.615
R112 VTAIL.n34 VTAIL.n33 104.615
R113 VTAIL.n34 VTAIL.n19 104.615
R114 VTAIL.n41 VTAIL.n19 104.615
R115 VTAIL.n43 VTAIL.n41 104.615
R116 VTAIL.n43 VTAIL.n42 104.615
R117 VTAIL.n42 VTAIL.n15 104.615
R118 VTAIL.n51 VTAIL.n15 104.615
R119 VTAIL.n52 VTAIL.n51 104.615
R120 VTAIL.n52 VTAIL.n11 104.615
R121 VTAIL.n59 VTAIL.n11 104.615
R122 VTAIL.n60 VTAIL.n59 104.615
R123 VTAIL.n60 VTAIL.n7 104.615
R124 VTAIL.n67 VTAIL.n7 104.615
R125 VTAIL.n68 VTAIL.n67 104.615
R126 VTAIL.n68 VTAIL.n3 104.615
R127 VTAIL.n75 VTAIL.n3 104.615
R128 VTAIL.n76 VTAIL.n75 104.615
R129 VTAIL.n240 VTAIL.n239 104.615
R130 VTAIL.n239 VTAIL.n167 104.615
R131 VTAIL.n232 VTAIL.n167 104.615
R132 VTAIL.n232 VTAIL.n231 104.615
R133 VTAIL.n231 VTAIL.n171 104.615
R134 VTAIL.n224 VTAIL.n171 104.615
R135 VTAIL.n224 VTAIL.n223 104.615
R136 VTAIL.n223 VTAIL.n175 104.615
R137 VTAIL.n216 VTAIL.n175 104.615
R138 VTAIL.n216 VTAIL.n215 104.615
R139 VTAIL.n215 VTAIL.n179 104.615
R140 VTAIL.n183 VTAIL.n179 104.615
R141 VTAIL.n207 VTAIL.n183 104.615
R142 VTAIL.n207 VTAIL.n206 104.615
R143 VTAIL.n206 VTAIL.n184 104.615
R144 VTAIL.n199 VTAIL.n184 104.615
R145 VTAIL.n199 VTAIL.n198 104.615
R146 VTAIL.n198 VTAIL.n188 104.615
R147 VTAIL.n191 VTAIL.n188 104.615
R148 VTAIL.n158 VTAIL.n157 104.615
R149 VTAIL.n157 VTAIL.n85 104.615
R150 VTAIL.n150 VTAIL.n85 104.615
R151 VTAIL.n150 VTAIL.n149 104.615
R152 VTAIL.n149 VTAIL.n89 104.615
R153 VTAIL.n142 VTAIL.n89 104.615
R154 VTAIL.n142 VTAIL.n141 104.615
R155 VTAIL.n141 VTAIL.n93 104.615
R156 VTAIL.n134 VTAIL.n93 104.615
R157 VTAIL.n134 VTAIL.n133 104.615
R158 VTAIL.n133 VTAIL.n97 104.615
R159 VTAIL.n101 VTAIL.n97 104.615
R160 VTAIL.n125 VTAIL.n101 104.615
R161 VTAIL.n125 VTAIL.n124 104.615
R162 VTAIL.n124 VTAIL.n102 104.615
R163 VTAIL.n117 VTAIL.n102 104.615
R164 VTAIL.n117 VTAIL.n116 104.615
R165 VTAIL.n116 VTAIL.n106 104.615
R166 VTAIL.n109 VTAIL.n106 104.615
R167 VTAIL.n272 VTAIL.t1 52.3082
R168 VTAIL.n26 VTAIL.t2 52.3082
R169 VTAIL.n191 VTAIL.t3 52.3082
R170 VTAIL.n109 VTAIL.t0 52.3082
R171 VTAIL.n327 VTAIL.n326 30.4399
R172 VTAIL.n81 VTAIL.n80 30.4399
R173 VTAIL.n245 VTAIL.n244 30.4399
R174 VTAIL.n163 VTAIL.n162 30.4399
R175 VTAIL.n163 VTAIL.n81 27.5824
R176 VTAIL.n327 VTAIL.n245 26.41
R177 VTAIL.n296 VTAIL.n295 13.1884
R178 VTAIL.n50 VTAIL.n49 13.1884
R179 VTAIL.n214 VTAIL.n213 13.1884
R180 VTAIL.n132 VTAIL.n131 13.1884
R181 VTAIL.n294 VTAIL.n262 12.8005
R182 VTAIL.n299 VTAIL.n260 12.8005
R183 VTAIL.n48 VTAIL.n16 12.8005
R184 VTAIL.n53 VTAIL.n14 12.8005
R185 VTAIL.n217 VTAIL.n178 12.8005
R186 VTAIL.n212 VTAIL.n180 12.8005
R187 VTAIL.n135 VTAIL.n96 12.8005
R188 VTAIL.n130 VTAIL.n98 12.8005
R189 VTAIL.n291 VTAIL.n290 12.0247
R190 VTAIL.n300 VTAIL.n258 12.0247
R191 VTAIL.n45 VTAIL.n44 12.0247
R192 VTAIL.n54 VTAIL.n12 12.0247
R193 VTAIL.n218 VTAIL.n176 12.0247
R194 VTAIL.n209 VTAIL.n208 12.0247
R195 VTAIL.n136 VTAIL.n94 12.0247
R196 VTAIL.n127 VTAIL.n126 12.0247
R197 VTAIL.n286 VTAIL.n264 11.249
R198 VTAIL.n304 VTAIL.n303 11.249
R199 VTAIL.n40 VTAIL.n18 11.249
R200 VTAIL.n58 VTAIL.n57 11.249
R201 VTAIL.n222 VTAIL.n221 11.249
R202 VTAIL.n205 VTAIL.n182 11.249
R203 VTAIL.n140 VTAIL.n139 11.249
R204 VTAIL.n123 VTAIL.n100 11.249
R205 VTAIL.n285 VTAIL.n266 10.4732
R206 VTAIL.n307 VTAIL.n256 10.4732
R207 VTAIL.n39 VTAIL.n20 10.4732
R208 VTAIL.n61 VTAIL.n10 10.4732
R209 VTAIL.n225 VTAIL.n174 10.4732
R210 VTAIL.n204 VTAIL.n185 10.4732
R211 VTAIL.n143 VTAIL.n92 10.4732
R212 VTAIL.n122 VTAIL.n103 10.4732
R213 VTAIL.n273 VTAIL.n271 10.2747
R214 VTAIL.n27 VTAIL.n25 10.2747
R215 VTAIL.n192 VTAIL.n190 10.2747
R216 VTAIL.n110 VTAIL.n108 10.2747
R217 VTAIL.n282 VTAIL.n281 9.69747
R218 VTAIL.n308 VTAIL.n254 9.69747
R219 VTAIL.n36 VTAIL.n35 9.69747
R220 VTAIL.n62 VTAIL.n8 9.69747
R221 VTAIL.n226 VTAIL.n172 9.69747
R222 VTAIL.n201 VTAIL.n200 9.69747
R223 VTAIL.n144 VTAIL.n90 9.69747
R224 VTAIL.n119 VTAIL.n118 9.69747
R225 VTAIL.n326 VTAIL.n325 9.45567
R226 VTAIL.n80 VTAIL.n79 9.45567
R227 VTAIL.n244 VTAIL.n243 9.45567
R228 VTAIL.n162 VTAIL.n161 9.45567
R229 VTAIL.n319 VTAIL.n318 9.3005
R230 VTAIL.n248 VTAIL.n247 9.3005
R231 VTAIL.n325 VTAIL.n324 9.3005
R232 VTAIL.n252 VTAIL.n251 9.3005
R233 VTAIL.n311 VTAIL.n310 9.3005
R234 VTAIL.n309 VTAIL.n308 9.3005
R235 VTAIL.n256 VTAIL.n255 9.3005
R236 VTAIL.n303 VTAIL.n302 9.3005
R237 VTAIL.n301 VTAIL.n300 9.3005
R238 VTAIL.n260 VTAIL.n259 9.3005
R239 VTAIL.n275 VTAIL.n274 9.3005
R240 VTAIL.n277 VTAIL.n276 9.3005
R241 VTAIL.n268 VTAIL.n267 9.3005
R242 VTAIL.n283 VTAIL.n282 9.3005
R243 VTAIL.n285 VTAIL.n284 9.3005
R244 VTAIL.n264 VTAIL.n263 9.3005
R245 VTAIL.n292 VTAIL.n291 9.3005
R246 VTAIL.n294 VTAIL.n293 9.3005
R247 VTAIL.n317 VTAIL.n316 9.3005
R248 VTAIL.n73 VTAIL.n72 9.3005
R249 VTAIL.n2 VTAIL.n1 9.3005
R250 VTAIL.n79 VTAIL.n78 9.3005
R251 VTAIL.n6 VTAIL.n5 9.3005
R252 VTAIL.n65 VTAIL.n64 9.3005
R253 VTAIL.n63 VTAIL.n62 9.3005
R254 VTAIL.n10 VTAIL.n9 9.3005
R255 VTAIL.n57 VTAIL.n56 9.3005
R256 VTAIL.n55 VTAIL.n54 9.3005
R257 VTAIL.n14 VTAIL.n13 9.3005
R258 VTAIL.n29 VTAIL.n28 9.3005
R259 VTAIL.n31 VTAIL.n30 9.3005
R260 VTAIL.n22 VTAIL.n21 9.3005
R261 VTAIL.n37 VTAIL.n36 9.3005
R262 VTAIL.n39 VTAIL.n38 9.3005
R263 VTAIL.n18 VTAIL.n17 9.3005
R264 VTAIL.n46 VTAIL.n45 9.3005
R265 VTAIL.n48 VTAIL.n47 9.3005
R266 VTAIL.n71 VTAIL.n70 9.3005
R267 VTAIL.n166 VTAIL.n165 9.3005
R268 VTAIL.n237 VTAIL.n236 9.3005
R269 VTAIL.n235 VTAIL.n234 9.3005
R270 VTAIL.n170 VTAIL.n169 9.3005
R271 VTAIL.n229 VTAIL.n228 9.3005
R272 VTAIL.n227 VTAIL.n226 9.3005
R273 VTAIL.n174 VTAIL.n173 9.3005
R274 VTAIL.n221 VTAIL.n220 9.3005
R275 VTAIL.n219 VTAIL.n218 9.3005
R276 VTAIL.n178 VTAIL.n177 9.3005
R277 VTAIL.n212 VTAIL.n211 9.3005
R278 VTAIL.n210 VTAIL.n209 9.3005
R279 VTAIL.n182 VTAIL.n181 9.3005
R280 VTAIL.n204 VTAIL.n203 9.3005
R281 VTAIL.n202 VTAIL.n201 9.3005
R282 VTAIL.n187 VTAIL.n186 9.3005
R283 VTAIL.n196 VTAIL.n195 9.3005
R284 VTAIL.n194 VTAIL.n193 9.3005
R285 VTAIL.n243 VTAIL.n242 9.3005
R286 VTAIL.n112 VTAIL.n111 9.3005
R287 VTAIL.n114 VTAIL.n113 9.3005
R288 VTAIL.n105 VTAIL.n104 9.3005
R289 VTAIL.n120 VTAIL.n119 9.3005
R290 VTAIL.n122 VTAIL.n121 9.3005
R291 VTAIL.n100 VTAIL.n99 9.3005
R292 VTAIL.n128 VTAIL.n127 9.3005
R293 VTAIL.n130 VTAIL.n129 9.3005
R294 VTAIL.n84 VTAIL.n83 9.3005
R295 VTAIL.n161 VTAIL.n160 9.3005
R296 VTAIL.n155 VTAIL.n154 9.3005
R297 VTAIL.n153 VTAIL.n152 9.3005
R298 VTAIL.n88 VTAIL.n87 9.3005
R299 VTAIL.n147 VTAIL.n146 9.3005
R300 VTAIL.n145 VTAIL.n144 9.3005
R301 VTAIL.n92 VTAIL.n91 9.3005
R302 VTAIL.n139 VTAIL.n138 9.3005
R303 VTAIL.n137 VTAIL.n136 9.3005
R304 VTAIL.n96 VTAIL.n95 9.3005
R305 VTAIL.n278 VTAIL.n268 8.92171
R306 VTAIL.n312 VTAIL.n311 8.92171
R307 VTAIL.n326 VTAIL.n246 8.92171
R308 VTAIL.n32 VTAIL.n22 8.92171
R309 VTAIL.n66 VTAIL.n65 8.92171
R310 VTAIL.n80 VTAIL.n0 8.92171
R311 VTAIL.n244 VTAIL.n164 8.92171
R312 VTAIL.n230 VTAIL.n229 8.92171
R313 VTAIL.n197 VTAIL.n187 8.92171
R314 VTAIL.n162 VTAIL.n82 8.92171
R315 VTAIL.n148 VTAIL.n147 8.92171
R316 VTAIL.n115 VTAIL.n105 8.92171
R317 VTAIL.n277 VTAIL.n270 8.14595
R318 VTAIL.n315 VTAIL.n252 8.14595
R319 VTAIL.n324 VTAIL.n323 8.14595
R320 VTAIL.n31 VTAIL.n24 8.14595
R321 VTAIL.n69 VTAIL.n6 8.14595
R322 VTAIL.n78 VTAIL.n77 8.14595
R323 VTAIL.n242 VTAIL.n241 8.14595
R324 VTAIL.n233 VTAIL.n170 8.14595
R325 VTAIL.n196 VTAIL.n189 8.14595
R326 VTAIL.n160 VTAIL.n159 8.14595
R327 VTAIL.n151 VTAIL.n88 8.14595
R328 VTAIL.n114 VTAIL.n107 8.14595
R329 VTAIL.n274 VTAIL.n273 7.3702
R330 VTAIL.n316 VTAIL.n250 7.3702
R331 VTAIL.n320 VTAIL.n248 7.3702
R332 VTAIL.n28 VTAIL.n27 7.3702
R333 VTAIL.n70 VTAIL.n4 7.3702
R334 VTAIL.n74 VTAIL.n2 7.3702
R335 VTAIL.n238 VTAIL.n166 7.3702
R336 VTAIL.n234 VTAIL.n168 7.3702
R337 VTAIL.n193 VTAIL.n192 7.3702
R338 VTAIL.n156 VTAIL.n84 7.3702
R339 VTAIL.n152 VTAIL.n86 7.3702
R340 VTAIL.n111 VTAIL.n110 7.3702
R341 VTAIL.n319 VTAIL.n250 6.59444
R342 VTAIL.n320 VTAIL.n319 6.59444
R343 VTAIL.n73 VTAIL.n4 6.59444
R344 VTAIL.n74 VTAIL.n73 6.59444
R345 VTAIL.n238 VTAIL.n237 6.59444
R346 VTAIL.n237 VTAIL.n168 6.59444
R347 VTAIL.n156 VTAIL.n155 6.59444
R348 VTAIL.n155 VTAIL.n86 6.59444
R349 VTAIL.n274 VTAIL.n270 5.81868
R350 VTAIL.n316 VTAIL.n315 5.81868
R351 VTAIL.n323 VTAIL.n248 5.81868
R352 VTAIL.n28 VTAIL.n24 5.81868
R353 VTAIL.n70 VTAIL.n69 5.81868
R354 VTAIL.n77 VTAIL.n2 5.81868
R355 VTAIL.n241 VTAIL.n166 5.81868
R356 VTAIL.n234 VTAIL.n233 5.81868
R357 VTAIL.n193 VTAIL.n189 5.81868
R358 VTAIL.n159 VTAIL.n84 5.81868
R359 VTAIL.n152 VTAIL.n151 5.81868
R360 VTAIL.n111 VTAIL.n107 5.81868
R361 VTAIL.n278 VTAIL.n277 5.04292
R362 VTAIL.n312 VTAIL.n252 5.04292
R363 VTAIL.n324 VTAIL.n246 5.04292
R364 VTAIL.n32 VTAIL.n31 5.04292
R365 VTAIL.n66 VTAIL.n6 5.04292
R366 VTAIL.n78 VTAIL.n0 5.04292
R367 VTAIL.n242 VTAIL.n164 5.04292
R368 VTAIL.n230 VTAIL.n170 5.04292
R369 VTAIL.n197 VTAIL.n196 5.04292
R370 VTAIL.n160 VTAIL.n82 5.04292
R371 VTAIL.n148 VTAIL.n88 5.04292
R372 VTAIL.n115 VTAIL.n114 5.04292
R373 VTAIL.n281 VTAIL.n268 4.26717
R374 VTAIL.n311 VTAIL.n254 4.26717
R375 VTAIL.n35 VTAIL.n22 4.26717
R376 VTAIL.n65 VTAIL.n8 4.26717
R377 VTAIL.n229 VTAIL.n172 4.26717
R378 VTAIL.n200 VTAIL.n187 4.26717
R379 VTAIL.n147 VTAIL.n90 4.26717
R380 VTAIL.n118 VTAIL.n105 4.26717
R381 VTAIL.n282 VTAIL.n266 3.49141
R382 VTAIL.n308 VTAIL.n307 3.49141
R383 VTAIL.n36 VTAIL.n20 3.49141
R384 VTAIL.n62 VTAIL.n61 3.49141
R385 VTAIL.n226 VTAIL.n225 3.49141
R386 VTAIL.n201 VTAIL.n185 3.49141
R387 VTAIL.n144 VTAIL.n143 3.49141
R388 VTAIL.n119 VTAIL.n103 3.49141
R389 VTAIL.n275 VTAIL.n271 2.84303
R390 VTAIL.n29 VTAIL.n25 2.84303
R391 VTAIL.n194 VTAIL.n190 2.84303
R392 VTAIL.n112 VTAIL.n108 2.84303
R393 VTAIL.n286 VTAIL.n285 2.71565
R394 VTAIL.n304 VTAIL.n256 2.71565
R395 VTAIL.n40 VTAIL.n39 2.71565
R396 VTAIL.n58 VTAIL.n10 2.71565
R397 VTAIL.n222 VTAIL.n174 2.71565
R398 VTAIL.n205 VTAIL.n204 2.71565
R399 VTAIL.n140 VTAIL.n92 2.71565
R400 VTAIL.n123 VTAIL.n122 2.71565
R401 VTAIL.n290 VTAIL.n264 1.93989
R402 VTAIL.n303 VTAIL.n258 1.93989
R403 VTAIL.n44 VTAIL.n18 1.93989
R404 VTAIL.n57 VTAIL.n12 1.93989
R405 VTAIL.n221 VTAIL.n176 1.93989
R406 VTAIL.n208 VTAIL.n182 1.93989
R407 VTAIL.n139 VTAIL.n94 1.93989
R408 VTAIL.n126 VTAIL.n100 1.93989
R409 VTAIL.n291 VTAIL.n262 1.16414
R410 VTAIL.n300 VTAIL.n299 1.16414
R411 VTAIL.n45 VTAIL.n16 1.16414
R412 VTAIL.n54 VTAIL.n53 1.16414
R413 VTAIL.n218 VTAIL.n217 1.16414
R414 VTAIL.n209 VTAIL.n180 1.16414
R415 VTAIL.n136 VTAIL.n135 1.16414
R416 VTAIL.n127 VTAIL.n98 1.16414
R417 VTAIL.n245 VTAIL.n163 1.05653
R418 VTAIL VTAIL.n81 0.821621
R419 VTAIL.n295 VTAIL.n294 0.388379
R420 VTAIL.n296 VTAIL.n260 0.388379
R421 VTAIL.n49 VTAIL.n48 0.388379
R422 VTAIL.n50 VTAIL.n14 0.388379
R423 VTAIL.n214 VTAIL.n178 0.388379
R424 VTAIL.n213 VTAIL.n212 0.388379
R425 VTAIL.n132 VTAIL.n96 0.388379
R426 VTAIL.n131 VTAIL.n130 0.388379
R427 VTAIL VTAIL.n327 0.235414
R428 VTAIL.n276 VTAIL.n275 0.155672
R429 VTAIL.n276 VTAIL.n267 0.155672
R430 VTAIL.n283 VTAIL.n267 0.155672
R431 VTAIL.n284 VTAIL.n283 0.155672
R432 VTAIL.n284 VTAIL.n263 0.155672
R433 VTAIL.n292 VTAIL.n263 0.155672
R434 VTAIL.n293 VTAIL.n292 0.155672
R435 VTAIL.n293 VTAIL.n259 0.155672
R436 VTAIL.n301 VTAIL.n259 0.155672
R437 VTAIL.n302 VTAIL.n301 0.155672
R438 VTAIL.n302 VTAIL.n255 0.155672
R439 VTAIL.n309 VTAIL.n255 0.155672
R440 VTAIL.n310 VTAIL.n309 0.155672
R441 VTAIL.n310 VTAIL.n251 0.155672
R442 VTAIL.n317 VTAIL.n251 0.155672
R443 VTAIL.n318 VTAIL.n317 0.155672
R444 VTAIL.n318 VTAIL.n247 0.155672
R445 VTAIL.n325 VTAIL.n247 0.155672
R446 VTAIL.n30 VTAIL.n29 0.155672
R447 VTAIL.n30 VTAIL.n21 0.155672
R448 VTAIL.n37 VTAIL.n21 0.155672
R449 VTAIL.n38 VTAIL.n37 0.155672
R450 VTAIL.n38 VTAIL.n17 0.155672
R451 VTAIL.n46 VTAIL.n17 0.155672
R452 VTAIL.n47 VTAIL.n46 0.155672
R453 VTAIL.n47 VTAIL.n13 0.155672
R454 VTAIL.n55 VTAIL.n13 0.155672
R455 VTAIL.n56 VTAIL.n55 0.155672
R456 VTAIL.n56 VTAIL.n9 0.155672
R457 VTAIL.n63 VTAIL.n9 0.155672
R458 VTAIL.n64 VTAIL.n63 0.155672
R459 VTAIL.n64 VTAIL.n5 0.155672
R460 VTAIL.n71 VTAIL.n5 0.155672
R461 VTAIL.n72 VTAIL.n71 0.155672
R462 VTAIL.n72 VTAIL.n1 0.155672
R463 VTAIL.n79 VTAIL.n1 0.155672
R464 VTAIL.n243 VTAIL.n165 0.155672
R465 VTAIL.n236 VTAIL.n165 0.155672
R466 VTAIL.n236 VTAIL.n235 0.155672
R467 VTAIL.n235 VTAIL.n169 0.155672
R468 VTAIL.n228 VTAIL.n169 0.155672
R469 VTAIL.n228 VTAIL.n227 0.155672
R470 VTAIL.n227 VTAIL.n173 0.155672
R471 VTAIL.n220 VTAIL.n173 0.155672
R472 VTAIL.n220 VTAIL.n219 0.155672
R473 VTAIL.n219 VTAIL.n177 0.155672
R474 VTAIL.n211 VTAIL.n177 0.155672
R475 VTAIL.n211 VTAIL.n210 0.155672
R476 VTAIL.n210 VTAIL.n181 0.155672
R477 VTAIL.n203 VTAIL.n181 0.155672
R478 VTAIL.n203 VTAIL.n202 0.155672
R479 VTAIL.n202 VTAIL.n186 0.155672
R480 VTAIL.n195 VTAIL.n186 0.155672
R481 VTAIL.n195 VTAIL.n194 0.155672
R482 VTAIL.n161 VTAIL.n83 0.155672
R483 VTAIL.n154 VTAIL.n83 0.155672
R484 VTAIL.n154 VTAIL.n153 0.155672
R485 VTAIL.n153 VTAIL.n87 0.155672
R486 VTAIL.n146 VTAIL.n87 0.155672
R487 VTAIL.n146 VTAIL.n145 0.155672
R488 VTAIL.n145 VTAIL.n91 0.155672
R489 VTAIL.n138 VTAIL.n91 0.155672
R490 VTAIL.n138 VTAIL.n137 0.155672
R491 VTAIL.n137 VTAIL.n95 0.155672
R492 VTAIL.n129 VTAIL.n95 0.155672
R493 VTAIL.n129 VTAIL.n128 0.155672
R494 VTAIL.n128 VTAIL.n99 0.155672
R495 VTAIL.n121 VTAIL.n99 0.155672
R496 VTAIL.n121 VTAIL.n120 0.155672
R497 VTAIL.n120 VTAIL.n104 0.155672
R498 VTAIL.n113 VTAIL.n104 0.155672
R499 VTAIL.n113 VTAIL.n112 0.155672
R500 VDD1.n76 VDD1.n0 289.615
R501 VDD1.n157 VDD1.n81 289.615
R502 VDD1.n77 VDD1.n76 185
R503 VDD1.n75 VDD1.n74 185
R504 VDD1.n4 VDD1.n3 185
R505 VDD1.n69 VDD1.n68 185
R506 VDD1.n67 VDD1.n66 185
R507 VDD1.n8 VDD1.n7 185
R508 VDD1.n61 VDD1.n60 185
R509 VDD1.n59 VDD1.n58 185
R510 VDD1.n12 VDD1.n11 185
R511 VDD1.n53 VDD1.n52 185
R512 VDD1.n51 VDD1.n50 185
R513 VDD1.n49 VDD1.n15 185
R514 VDD1.n19 VDD1.n16 185
R515 VDD1.n44 VDD1.n43 185
R516 VDD1.n42 VDD1.n41 185
R517 VDD1.n21 VDD1.n20 185
R518 VDD1.n36 VDD1.n35 185
R519 VDD1.n34 VDD1.n33 185
R520 VDD1.n25 VDD1.n24 185
R521 VDD1.n28 VDD1.n27 185
R522 VDD1.n108 VDD1.n107 185
R523 VDD1.n105 VDD1.n104 185
R524 VDD1.n114 VDD1.n113 185
R525 VDD1.n116 VDD1.n115 185
R526 VDD1.n101 VDD1.n100 185
R527 VDD1.n122 VDD1.n121 185
R528 VDD1.n125 VDD1.n124 185
R529 VDD1.n123 VDD1.n97 185
R530 VDD1.n130 VDD1.n96 185
R531 VDD1.n132 VDD1.n131 185
R532 VDD1.n134 VDD1.n133 185
R533 VDD1.n93 VDD1.n92 185
R534 VDD1.n140 VDD1.n139 185
R535 VDD1.n142 VDD1.n141 185
R536 VDD1.n89 VDD1.n88 185
R537 VDD1.n148 VDD1.n147 185
R538 VDD1.n150 VDD1.n149 185
R539 VDD1.n85 VDD1.n84 185
R540 VDD1.n156 VDD1.n155 185
R541 VDD1.n158 VDD1.n157 185
R542 VDD1.t0 VDD1.n26 149.524
R543 VDD1.t1 VDD1.n106 149.524
R544 VDD1.n76 VDD1.n75 104.615
R545 VDD1.n75 VDD1.n3 104.615
R546 VDD1.n68 VDD1.n3 104.615
R547 VDD1.n68 VDD1.n67 104.615
R548 VDD1.n67 VDD1.n7 104.615
R549 VDD1.n60 VDD1.n7 104.615
R550 VDD1.n60 VDD1.n59 104.615
R551 VDD1.n59 VDD1.n11 104.615
R552 VDD1.n52 VDD1.n11 104.615
R553 VDD1.n52 VDD1.n51 104.615
R554 VDD1.n51 VDD1.n15 104.615
R555 VDD1.n19 VDD1.n15 104.615
R556 VDD1.n43 VDD1.n19 104.615
R557 VDD1.n43 VDD1.n42 104.615
R558 VDD1.n42 VDD1.n20 104.615
R559 VDD1.n35 VDD1.n20 104.615
R560 VDD1.n35 VDD1.n34 104.615
R561 VDD1.n34 VDD1.n24 104.615
R562 VDD1.n27 VDD1.n24 104.615
R563 VDD1.n107 VDD1.n104 104.615
R564 VDD1.n114 VDD1.n104 104.615
R565 VDD1.n115 VDD1.n114 104.615
R566 VDD1.n115 VDD1.n100 104.615
R567 VDD1.n122 VDD1.n100 104.615
R568 VDD1.n124 VDD1.n122 104.615
R569 VDD1.n124 VDD1.n123 104.615
R570 VDD1.n123 VDD1.n96 104.615
R571 VDD1.n132 VDD1.n96 104.615
R572 VDD1.n133 VDD1.n132 104.615
R573 VDD1.n133 VDD1.n92 104.615
R574 VDD1.n140 VDD1.n92 104.615
R575 VDD1.n141 VDD1.n140 104.615
R576 VDD1.n141 VDD1.n88 104.615
R577 VDD1.n148 VDD1.n88 104.615
R578 VDD1.n149 VDD1.n148 104.615
R579 VDD1.n149 VDD1.n84 104.615
R580 VDD1.n156 VDD1.n84 104.615
R581 VDD1.n157 VDD1.n156 104.615
R582 VDD1 VDD1.n161 86.8116
R583 VDD1.n27 VDD1.t0 52.3082
R584 VDD1.n107 VDD1.t1 52.3082
R585 VDD1 VDD1.n80 47.47
R586 VDD1.n50 VDD1.n49 13.1884
R587 VDD1.n131 VDD1.n130 13.1884
R588 VDD1.n53 VDD1.n14 12.8005
R589 VDD1.n48 VDD1.n16 12.8005
R590 VDD1.n129 VDD1.n97 12.8005
R591 VDD1.n134 VDD1.n95 12.8005
R592 VDD1.n54 VDD1.n12 12.0247
R593 VDD1.n45 VDD1.n44 12.0247
R594 VDD1.n126 VDD1.n125 12.0247
R595 VDD1.n135 VDD1.n93 12.0247
R596 VDD1.n58 VDD1.n57 11.249
R597 VDD1.n41 VDD1.n18 11.249
R598 VDD1.n121 VDD1.n99 11.249
R599 VDD1.n139 VDD1.n138 11.249
R600 VDD1.n61 VDD1.n10 10.4732
R601 VDD1.n40 VDD1.n21 10.4732
R602 VDD1.n120 VDD1.n101 10.4732
R603 VDD1.n142 VDD1.n91 10.4732
R604 VDD1.n28 VDD1.n26 10.2747
R605 VDD1.n108 VDD1.n106 10.2747
R606 VDD1.n62 VDD1.n8 9.69747
R607 VDD1.n37 VDD1.n36 9.69747
R608 VDD1.n117 VDD1.n116 9.69747
R609 VDD1.n143 VDD1.n89 9.69747
R610 VDD1.n80 VDD1.n79 9.45567
R611 VDD1.n161 VDD1.n160 9.45567
R612 VDD1.n2 VDD1.n1 9.3005
R613 VDD1.n73 VDD1.n72 9.3005
R614 VDD1.n71 VDD1.n70 9.3005
R615 VDD1.n6 VDD1.n5 9.3005
R616 VDD1.n65 VDD1.n64 9.3005
R617 VDD1.n63 VDD1.n62 9.3005
R618 VDD1.n10 VDD1.n9 9.3005
R619 VDD1.n57 VDD1.n56 9.3005
R620 VDD1.n55 VDD1.n54 9.3005
R621 VDD1.n14 VDD1.n13 9.3005
R622 VDD1.n48 VDD1.n47 9.3005
R623 VDD1.n46 VDD1.n45 9.3005
R624 VDD1.n18 VDD1.n17 9.3005
R625 VDD1.n40 VDD1.n39 9.3005
R626 VDD1.n38 VDD1.n37 9.3005
R627 VDD1.n23 VDD1.n22 9.3005
R628 VDD1.n32 VDD1.n31 9.3005
R629 VDD1.n30 VDD1.n29 9.3005
R630 VDD1.n79 VDD1.n78 9.3005
R631 VDD1.n154 VDD1.n153 9.3005
R632 VDD1.n83 VDD1.n82 9.3005
R633 VDD1.n160 VDD1.n159 9.3005
R634 VDD1.n87 VDD1.n86 9.3005
R635 VDD1.n146 VDD1.n145 9.3005
R636 VDD1.n144 VDD1.n143 9.3005
R637 VDD1.n91 VDD1.n90 9.3005
R638 VDD1.n138 VDD1.n137 9.3005
R639 VDD1.n136 VDD1.n135 9.3005
R640 VDD1.n95 VDD1.n94 9.3005
R641 VDD1.n110 VDD1.n109 9.3005
R642 VDD1.n112 VDD1.n111 9.3005
R643 VDD1.n103 VDD1.n102 9.3005
R644 VDD1.n118 VDD1.n117 9.3005
R645 VDD1.n120 VDD1.n119 9.3005
R646 VDD1.n99 VDD1.n98 9.3005
R647 VDD1.n127 VDD1.n126 9.3005
R648 VDD1.n129 VDD1.n128 9.3005
R649 VDD1.n152 VDD1.n151 9.3005
R650 VDD1.n80 VDD1.n0 8.92171
R651 VDD1.n66 VDD1.n65 8.92171
R652 VDD1.n33 VDD1.n23 8.92171
R653 VDD1.n113 VDD1.n103 8.92171
R654 VDD1.n147 VDD1.n146 8.92171
R655 VDD1.n161 VDD1.n81 8.92171
R656 VDD1.n78 VDD1.n77 8.14595
R657 VDD1.n69 VDD1.n6 8.14595
R658 VDD1.n32 VDD1.n25 8.14595
R659 VDD1.n112 VDD1.n105 8.14595
R660 VDD1.n150 VDD1.n87 8.14595
R661 VDD1.n159 VDD1.n158 8.14595
R662 VDD1.n74 VDD1.n2 7.3702
R663 VDD1.n70 VDD1.n4 7.3702
R664 VDD1.n29 VDD1.n28 7.3702
R665 VDD1.n109 VDD1.n108 7.3702
R666 VDD1.n151 VDD1.n85 7.3702
R667 VDD1.n155 VDD1.n83 7.3702
R668 VDD1.n74 VDD1.n73 6.59444
R669 VDD1.n73 VDD1.n4 6.59444
R670 VDD1.n154 VDD1.n85 6.59444
R671 VDD1.n155 VDD1.n154 6.59444
R672 VDD1.n77 VDD1.n2 5.81868
R673 VDD1.n70 VDD1.n69 5.81868
R674 VDD1.n29 VDD1.n25 5.81868
R675 VDD1.n109 VDD1.n105 5.81868
R676 VDD1.n151 VDD1.n150 5.81868
R677 VDD1.n158 VDD1.n83 5.81868
R678 VDD1.n78 VDD1.n0 5.04292
R679 VDD1.n66 VDD1.n6 5.04292
R680 VDD1.n33 VDD1.n32 5.04292
R681 VDD1.n113 VDD1.n112 5.04292
R682 VDD1.n147 VDD1.n87 5.04292
R683 VDD1.n159 VDD1.n81 5.04292
R684 VDD1.n65 VDD1.n8 4.26717
R685 VDD1.n36 VDD1.n23 4.26717
R686 VDD1.n116 VDD1.n103 4.26717
R687 VDD1.n146 VDD1.n89 4.26717
R688 VDD1.n62 VDD1.n61 3.49141
R689 VDD1.n37 VDD1.n21 3.49141
R690 VDD1.n117 VDD1.n101 3.49141
R691 VDD1.n143 VDD1.n142 3.49141
R692 VDD1.n110 VDD1.n106 2.84303
R693 VDD1.n30 VDD1.n26 2.84303
R694 VDD1.n58 VDD1.n10 2.71565
R695 VDD1.n41 VDD1.n40 2.71565
R696 VDD1.n121 VDD1.n120 2.71565
R697 VDD1.n139 VDD1.n91 2.71565
R698 VDD1.n57 VDD1.n12 1.93989
R699 VDD1.n44 VDD1.n18 1.93989
R700 VDD1.n125 VDD1.n99 1.93989
R701 VDD1.n138 VDD1.n93 1.93989
R702 VDD1.n54 VDD1.n53 1.16414
R703 VDD1.n45 VDD1.n16 1.16414
R704 VDD1.n126 VDD1.n97 1.16414
R705 VDD1.n135 VDD1.n134 1.16414
R706 VDD1.n50 VDD1.n14 0.388379
R707 VDD1.n49 VDD1.n48 0.388379
R708 VDD1.n130 VDD1.n129 0.388379
R709 VDD1.n131 VDD1.n95 0.388379
R710 VDD1.n79 VDD1.n1 0.155672
R711 VDD1.n72 VDD1.n1 0.155672
R712 VDD1.n72 VDD1.n71 0.155672
R713 VDD1.n71 VDD1.n5 0.155672
R714 VDD1.n64 VDD1.n5 0.155672
R715 VDD1.n64 VDD1.n63 0.155672
R716 VDD1.n63 VDD1.n9 0.155672
R717 VDD1.n56 VDD1.n9 0.155672
R718 VDD1.n56 VDD1.n55 0.155672
R719 VDD1.n55 VDD1.n13 0.155672
R720 VDD1.n47 VDD1.n13 0.155672
R721 VDD1.n47 VDD1.n46 0.155672
R722 VDD1.n46 VDD1.n17 0.155672
R723 VDD1.n39 VDD1.n17 0.155672
R724 VDD1.n39 VDD1.n38 0.155672
R725 VDD1.n38 VDD1.n22 0.155672
R726 VDD1.n31 VDD1.n22 0.155672
R727 VDD1.n31 VDD1.n30 0.155672
R728 VDD1.n111 VDD1.n110 0.155672
R729 VDD1.n111 VDD1.n102 0.155672
R730 VDD1.n118 VDD1.n102 0.155672
R731 VDD1.n119 VDD1.n118 0.155672
R732 VDD1.n119 VDD1.n98 0.155672
R733 VDD1.n127 VDD1.n98 0.155672
R734 VDD1.n128 VDD1.n127 0.155672
R735 VDD1.n128 VDD1.n94 0.155672
R736 VDD1.n136 VDD1.n94 0.155672
R737 VDD1.n137 VDD1.n136 0.155672
R738 VDD1.n137 VDD1.n90 0.155672
R739 VDD1.n144 VDD1.n90 0.155672
R740 VDD1.n145 VDD1.n144 0.155672
R741 VDD1.n145 VDD1.n86 0.155672
R742 VDD1.n152 VDD1.n86 0.155672
R743 VDD1.n153 VDD1.n152 0.155672
R744 VDD1.n153 VDD1.n82 0.155672
R745 VDD1.n160 VDD1.n82 0.155672
R746 B.n690 B.n689 585
R747 B.n309 B.n88 585
R748 B.n308 B.n307 585
R749 B.n306 B.n305 585
R750 B.n304 B.n303 585
R751 B.n302 B.n301 585
R752 B.n300 B.n299 585
R753 B.n298 B.n297 585
R754 B.n296 B.n295 585
R755 B.n294 B.n293 585
R756 B.n292 B.n291 585
R757 B.n290 B.n289 585
R758 B.n288 B.n287 585
R759 B.n286 B.n285 585
R760 B.n284 B.n283 585
R761 B.n282 B.n281 585
R762 B.n280 B.n279 585
R763 B.n278 B.n277 585
R764 B.n276 B.n275 585
R765 B.n274 B.n273 585
R766 B.n272 B.n271 585
R767 B.n270 B.n269 585
R768 B.n268 B.n267 585
R769 B.n266 B.n265 585
R770 B.n264 B.n263 585
R771 B.n262 B.n261 585
R772 B.n260 B.n259 585
R773 B.n258 B.n257 585
R774 B.n256 B.n255 585
R775 B.n254 B.n253 585
R776 B.n252 B.n251 585
R777 B.n250 B.n249 585
R778 B.n248 B.n247 585
R779 B.n246 B.n245 585
R780 B.n244 B.n243 585
R781 B.n242 B.n241 585
R782 B.n240 B.n239 585
R783 B.n238 B.n237 585
R784 B.n236 B.n235 585
R785 B.n234 B.n233 585
R786 B.n232 B.n231 585
R787 B.n230 B.n229 585
R788 B.n228 B.n227 585
R789 B.n226 B.n225 585
R790 B.n224 B.n223 585
R791 B.n222 B.n221 585
R792 B.n220 B.n219 585
R793 B.n218 B.n217 585
R794 B.n216 B.n215 585
R795 B.n214 B.n213 585
R796 B.n212 B.n211 585
R797 B.n210 B.n209 585
R798 B.n208 B.n207 585
R799 B.n206 B.n205 585
R800 B.n204 B.n203 585
R801 B.n202 B.n201 585
R802 B.n200 B.n199 585
R803 B.n198 B.n197 585
R804 B.n196 B.n195 585
R805 B.n194 B.n193 585
R806 B.n192 B.n191 585
R807 B.n190 B.n189 585
R808 B.n188 B.n187 585
R809 B.n186 B.n185 585
R810 B.n184 B.n183 585
R811 B.n182 B.n181 585
R812 B.n180 B.n179 585
R813 B.n178 B.n177 585
R814 B.n176 B.n175 585
R815 B.n174 B.n173 585
R816 B.n172 B.n171 585
R817 B.n170 B.n169 585
R818 B.n168 B.n167 585
R819 B.n166 B.n165 585
R820 B.n164 B.n163 585
R821 B.n162 B.n161 585
R822 B.n160 B.n159 585
R823 B.n158 B.n157 585
R824 B.n156 B.n155 585
R825 B.n154 B.n153 585
R826 B.n152 B.n151 585
R827 B.n150 B.n149 585
R828 B.n148 B.n147 585
R829 B.n146 B.n145 585
R830 B.n144 B.n143 585
R831 B.n142 B.n141 585
R832 B.n140 B.n139 585
R833 B.n138 B.n137 585
R834 B.n136 B.n135 585
R835 B.n134 B.n133 585
R836 B.n132 B.n131 585
R837 B.n130 B.n129 585
R838 B.n128 B.n127 585
R839 B.n126 B.n125 585
R840 B.n124 B.n123 585
R841 B.n122 B.n121 585
R842 B.n120 B.n119 585
R843 B.n118 B.n117 585
R844 B.n116 B.n115 585
R845 B.n114 B.n113 585
R846 B.n112 B.n111 585
R847 B.n110 B.n109 585
R848 B.n108 B.n107 585
R849 B.n106 B.n105 585
R850 B.n104 B.n103 585
R851 B.n102 B.n101 585
R852 B.n100 B.n99 585
R853 B.n98 B.n97 585
R854 B.n96 B.n95 585
R855 B.n32 B.n31 585
R856 B.n688 B.n33 585
R857 B.n693 B.n33 585
R858 B.n687 B.n686 585
R859 B.n686 B.n29 585
R860 B.n685 B.n28 585
R861 B.n699 B.n28 585
R862 B.n684 B.n27 585
R863 B.n700 B.n27 585
R864 B.n683 B.n26 585
R865 B.n701 B.n26 585
R866 B.n682 B.n681 585
R867 B.n681 B.n25 585
R868 B.n680 B.n21 585
R869 B.n707 B.n21 585
R870 B.n679 B.n20 585
R871 B.n708 B.n20 585
R872 B.n678 B.n19 585
R873 B.n709 B.n19 585
R874 B.n677 B.n676 585
R875 B.n676 B.n15 585
R876 B.n675 B.n14 585
R877 B.n715 B.n14 585
R878 B.n674 B.n13 585
R879 B.n716 B.n13 585
R880 B.n673 B.n12 585
R881 B.n717 B.n12 585
R882 B.n672 B.n671 585
R883 B.n671 B.n8 585
R884 B.n670 B.n7 585
R885 B.n723 B.n7 585
R886 B.n669 B.n6 585
R887 B.n724 B.n6 585
R888 B.n668 B.n5 585
R889 B.n725 B.n5 585
R890 B.n667 B.n666 585
R891 B.n666 B.n4 585
R892 B.n665 B.n310 585
R893 B.n665 B.n664 585
R894 B.n655 B.n311 585
R895 B.n312 B.n311 585
R896 B.n657 B.n656 585
R897 B.n658 B.n657 585
R898 B.n654 B.n317 585
R899 B.n317 B.n316 585
R900 B.n653 B.n652 585
R901 B.n652 B.n651 585
R902 B.n319 B.n318 585
R903 B.n320 B.n319 585
R904 B.n644 B.n643 585
R905 B.n645 B.n644 585
R906 B.n642 B.n325 585
R907 B.n325 B.n324 585
R908 B.n641 B.n640 585
R909 B.n640 B.n639 585
R910 B.n327 B.n326 585
R911 B.n632 B.n327 585
R912 B.n631 B.n630 585
R913 B.n633 B.n631 585
R914 B.n629 B.n332 585
R915 B.n332 B.n331 585
R916 B.n628 B.n627 585
R917 B.n627 B.n626 585
R918 B.n334 B.n333 585
R919 B.n335 B.n334 585
R920 B.n619 B.n618 585
R921 B.n620 B.n619 585
R922 B.n338 B.n337 585
R923 B.n399 B.n397 585
R924 B.n400 B.n396 585
R925 B.n400 B.n339 585
R926 B.n403 B.n402 585
R927 B.n404 B.n395 585
R928 B.n406 B.n405 585
R929 B.n408 B.n394 585
R930 B.n411 B.n410 585
R931 B.n412 B.n393 585
R932 B.n414 B.n413 585
R933 B.n416 B.n392 585
R934 B.n419 B.n418 585
R935 B.n420 B.n391 585
R936 B.n422 B.n421 585
R937 B.n424 B.n390 585
R938 B.n427 B.n426 585
R939 B.n428 B.n389 585
R940 B.n430 B.n429 585
R941 B.n432 B.n388 585
R942 B.n435 B.n434 585
R943 B.n436 B.n387 585
R944 B.n438 B.n437 585
R945 B.n440 B.n386 585
R946 B.n443 B.n442 585
R947 B.n444 B.n385 585
R948 B.n446 B.n445 585
R949 B.n448 B.n384 585
R950 B.n451 B.n450 585
R951 B.n452 B.n383 585
R952 B.n454 B.n453 585
R953 B.n456 B.n382 585
R954 B.n459 B.n458 585
R955 B.n460 B.n381 585
R956 B.n462 B.n461 585
R957 B.n464 B.n380 585
R958 B.n467 B.n466 585
R959 B.n468 B.n379 585
R960 B.n470 B.n469 585
R961 B.n472 B.n378 585
R962 B.n475 B.n474 585
R963 B.n476 B.n377 585
R964 B.n478 B.n477 585
R965 B.n480 B.n376 585
R966 B.n483 B.n482 585
R967 B.n484 B.n375 585
R968 B.n486 B.n485 585
R969 B.n488 B.n374 585
R970 B.n491 B.n490 585
R971 B.n492 B.n373 585
R972 B.n497 B.n496 585
R973 B.n499 B.n372 585
R974 B.n502 B.n501 585
R975 B.n503 B.n371 585
R976 B.n505 B.n504 585
R977 B.n507 B.n370 585
R978 B.n510 B.n509 585
R979 B.n511 B.n369 585
R980 B.n513 B.n512 585
R981 B.n515 B.n368 585
R982 B.n518 B.n517 585
R983 B.n520 B.n365 585
R984 B.n522 B.n521 585
R985 B.n524 B.n364 585
R986 B.n527 B.n526 585
R987 B.n528 B.n363 585
R988 B.n530 B.n529 585
R989 B.n532 B.n362 585
R990 B.n535 B.n534 585
R991 B.n536 B.n361 585
R992 B.n538 B.n537 585
R993 B.n540 B.n360 585
R994 B.n543 B.n542 585
R995 B.n544 B.n359 585
R996 B.n546 B.n545 585
R997 B.n548 B.n358 585
R998 B.n551 B.n550 585
R999 B.n552 B.n357 585
R1000 B.n554 B.n553 585
R1001 B.n556 B.n356 585
R1002 B.n559 B.n558 585
R1003 B.n560 B.n355 585
R1004 B.n562 B.n561 585
R1005 B.n564 B.n354 585
R1006 B.n567 B.n566 585
R1007 B.n568 B.n353 585
R1008 B.n570 B.n569 585
R1009 B.n572 B.n352 585
R1010 B.n575 B.n574 585
R1011 B.n576 B.n351 585
R1012 B.n578 B.n577 585
R1013 B.n580 B.n350 585
R1014 B.n583 B.n582 585
R1015 B.n584 B.n349 585
R1016 B.n586 B.n585 585
R1017 B.n588 B.n348 585
R1018 B.n591 B.n590 585
R1019 B.n592 B.n347 585
R1020 B.n594 B.n593 585
R1021 B.n596 B.n346 585
R1022 B.n599 B.n598 585
R1023 B.n600 B.n345 585
R1024 B.n602 B.n601 585
R1025 B.n604 B.n344 585
R1026 B.n607 B.n606 585
R1027 B.n608 B.n343 585
R1028 B.n610 B.n609 585
R1029 B.n612 B.n342 585
R1030 B.n613 B.n341 585
R1031 B.n616 B.n615 585
R1032 B.n617 B.n340 585
R1033 B.n340 B.n339 585
R1034 B.n622 B.n621 585
R1035 B.n621 B.n620 585
R1036 B.n623 B.n336 585
R1037 B.n336 B.n335 585
R1038 B.n625 B.n624 585
R1039 B.n626 B.n625 585
R1040 B.n330 B.n329 585
R1041 B.n331 B.n330 585
R1042 B.n635 B.n634 585
R1043 B.n634 B.n633 585
R1044 B.n636 B.n328 585
R1045 B.n632 B.n328 585
R1046 B.n638 B.n637 585
R1047 B.n639 B.n638 585
R1048 B.n323 B.n322 585
R1049 B.n324 B.n323 585
R1050 B.n647 B.n646 585
R1051 B.n646 B.n645 585
R1052 B.n648 B.n321 585
R1053 B.n321 B.n320 585
R1054 B.n650 B.n649 585
R1055 B.n651 B.n650 585
R1056 B.n315 B.n314 585
R1057 B.n316 B.n315 585
R1058 B.n660 B.n659 585
R1059 B.n659 B.n658 585
R1060 B.n661 B.n313 585
R1061 B.n313 B.n312 585
R1062 B.n663 B.n662 585
R1063 B.n664 B.n663 585
R1064 B.n2 B.n0 585
R1065 B.n4 B.n2 585
R1066 B.n3 B.n1 585
R1067 B.n724 B.n3 585
R1068 B.n722 B.n721 585
R1069 B.n723 B.n722 585
R1070 B.n720 B.n9 585
R1071 B.n9 B.n8 585
R1072 B.n719 B.n718 585
R1073 B.n718 B.n717 585
R1074 B.n11 B.n10 585
R1075 B.n716 B.n11 585
R1076 B.n714 B.n713 585
R1077 B.n715 B.n714 585
R1078 B.n712 B.n16 585
R1079 B.n16 B.n15 585
R1080 B.n711 B.n710 585
R1081 B.n710 B.n709 585
R1082 B.n18 B.n17 585
R1083 B.n708 B.n18 585
R1084 B.n706 B.n705 585
R1085 B.n707 B.n706 585
R1086 B.n704 B.n22 585
R1087 B.n25 B.n22 585
R1088 B.n703 B.n702 585
R1089 B.n702 B.n701 585
R1090 B.n24 B.n23 585
R1091 B.n700 B.n24 585
R1092 B.n698 B.n697 585
R1093 B.n699 B.n698 585
R1094 B.n696 B.n30 585
R1095 B.n30 B.n29 585
R1096 B.n695 B.n694 585
R1097 B.n694 B.n693 585
R1098 B.n727 B.n726 585
R1099 B.n726 B.n725 585
R1100 B.n366 B.t2 551.991
R1101 B.n493 B.t6 551.991
R1102 B.n92 B.t9 551.991
R1103 B.n89 B.t13 551.991
R1104 B.n621 B.n338 521.33
R1105 B.n694 B.n32 521.33
R1106 B.n619 B.n340 521.33
R1107 B.n690 B.n33 521.33
R1108 B.n366 B.t5 358.918
R1109 B.n89 B.t14 358.918
R1110 B.n493 B.t8 358.918
R1111 B.n92 B.t11 358.918
R1112 B.n367 B.t4 332.543
R1113 B.n90 B.t15 332.543
R1114 B.n494 B.t7 332.543
R1115 B.n93 B.t12 332.543
R1116 B.n692 B.n691 256.663
R1117 B.n692 B.n87 256.663
R1118 B.n692 B.n86 256.663
R1119 B.n692 B.n85 256.663
R1120 B.n692 B.n84 256.663
R1121 B.n692 B.n83 256.663
R1122 B.n692 B.n82 256.663
R1123 B.n692 B.n81 256.663
R1124 B.n692 B.n80 256.663
R1125 B.n692 B.n79 256.663
R1126 B.n692 B.n78 256.663
R1127 B.n692 B.n77 256.663
R1128 B.n692 B.n76 256.663
R1129 B.n692 B.n75 256.663
R1130 B.n692 B.n74 256.663
R1131 B.n692 B.n73 256.663
R1132 B.n692 B.n72 256.663
R1133 B.n692 B.n71 256.663
R1134 B.n692 B.n70 256.663
R1135 B.n692 B.n69 256.663
R1136 B.n692 B.n68 256.663
R1137 B.n692 B.n67 256.663
R1138 B.n692 B.n66 256.663
R1139 B.n692 B.n65 256.663
R1140 B.n692 B.n64 256.663
R1141 B.n692 B.n63 256.663
R1142 B.n692 B.n62 256.663
R1143 B.n692 B.n61 256.663
R1144 B.n692 B.n60 256.663
R1145 B.n692 B.n59 256.663
R1146 B.n692 B.n58 256.663
R1147 B.n692 B.n57 256.663
R1148 B.n692 B.n56 256.663
R1149 B.n692 B.n55 256.663
R1150 B.n692 B.n54 256.663
R1151 B.n692 B.n53 256.663
R1152 B.n692 B.n52 256.663
R1153 B.n692 B.n51 256.663
R1154 B.n692 B.n50 256.663
R1155 B.n692 B.n49 256.663
R1156 B.n692 B.n48 256.663
R1157 B.n692 B.n47 256.663
R1158 B.n692 B.n46 256.663
R1159 B.n692 B.n45 256.663
R1160 B.n692 B.n44 256.663
R1161 B.n692 B.n43 256.663
R1162 B.n692 B.n42 256.663
R1163 B.n692 B.n41 256.663
R1164 B.n692 B.n40 256.663
R1165 B.n692 B.n39 256.663
R1166 B.n692 B.n38 256.663
R1167 B.n692 B.n37 256.663
R1168 B.n692 B.n36 256.663
R1169 B.n692 B.n35 256.663
R1170 B.n692 B.n34 256.663
R1171 B.n398 B.n339 256.663
R1172 B.n401 B.n339 256.663
R1173 B.n407 B.n339 256.663
R1174 B.n409 B.n339 256.663
R1175 B.n415 B.n339 256.663
R1176 B.n417 B.n339 256.663
R1177 B.n423 B.n339 256.663
R1178 B.n425 B.n339 256.663
R1179 B.n431 B.n339 256.663
R1180 B.n433 B.n339 256.663
R1181 B.n439 B.n339 256.663
R1182 B.n441 B.n339 256.663
R1183 B.n447 B.n339 256.663
R1184 B.n449 B.n339 256.663
R1185 B.n455 B.n339 256.663
R1186 B.n457 B.n339 256.663
R1187 B.n463 B.n339 256.663
R1188 B.n465 B.n339 256.663
R1189 B.n471 B.n339 256.663
R1190 B.n473 B.n339 256.663
R1191 B.n479 B.n339 256.663
R1192 B.n481 B.n339 256.663
R1193 B.n487 B.n339 256.663
R1194 B.n489 B.n339 256.663
R1195 B.n498 B.n339 256.663
R1196 B.n500 B.n339 256.663
R1197 B.n506 B.n339 256.663
R1198 B.n508 B.n339 256.663
R1199 B.n514 B.n339 256.663
R1200 B.n516 B.n339 256.663
R1201 B.n523 B.n339 256.663
R1202 B.n525 B.n339 256.663
R1203 B.n531 B.n339 256.663
R1204 B.n533 B.n339 256.663
R1205 B.n539 B.n339 256.663
R1206 B.n541 B.n339 256.663
R1207 B.n547 B.n339 256.663
R1208 B.n549 B.n339 256.663
R1209 B.n555 B.n339 256.663
R1210 B.n557 B.n339 256.663
R1211 B.n563 B.n339 256.663
R1212 B.n565 B.n339 256.663
R1213 B.n571 B.n339 256.663
R1214 B.n573 B.n339 256.663
R1215 B.n579 B.n339 256.663
R1216 B.n581 B.n339 256.663
R1217 B.n587 B.n339 256.663
R1218 B.n589 B.n339 256.663
R1219 B.n595 B.n339 256.663
R1220 B.n597 B.n339 256.663
R1221 B.n603 B.n339 256.663
R1222 B.n605 B.n339 256.663
R1223 B.n611 B.n339 256.663
R1224 B.n614 B.n339 256.663
R1225 B.n621 B.n336 163.367
R1226 B.n625 B.n336 163.367
R1227 B.n625 B.n330 163.367
R1228 B.n634 B.n330 163.367
R1229 B.n634 B.n328 163.367
R1230 B.n638 B.n328 163.367
R1231 B.n638 B.n323 163.367
R1232 B.n646 B.n323 163.367
R1233 B.n646 B.n321 163.367
R1234 B.n650 B.n321 163.367
R1235 B.n650 B.n315 163.367
R1236 B.n659 B.n315 163.367
R1237 B.n659 B.n313 163.367
R1238 B.n663 B.n313 163.367
R1239 B.n663 B.n2 163.367
R1240 B.n726 B.n2 163.367
R1241 B.n726 B.n3 163.367
R1242 B.n722 B.n3 163.367
R1243 B.n722 B.n9 163.367
R1244 B.n718 B.n9 163.367
R1245 B.n718 B.n11 163.367
R1246 B.n714 B.n11 163.367
R1247 B.n714 B.n16 163.367
R1248 B.n710 B.n16 163.367
R1249 B.n710 B.n18 163.367
R1250 B.n706 B.n18 163.367
R1251 B.n706 B.n22 163.367
R1252 B.n702 B.n22 163.367
R1253 B.n702 B.n24 163.367
R1254 B.n698 B.n24 163.367
R1255 B.n698 B.n30 163.367
R1256 B.n694 B.n30 163.367
R1257 B.n400 B.n399 163.367
R1258 B.n402 B.n400 163.367
R1259 B.n406 B.n395 163.367
R1260 B.n410 B.n408 163.367
R1261 B.n414 B.n393 163.367
R1262 B.n418 B.n416 163.367
R1263 B.n422 B.n391 163.367
R1264 B.n426 B.n424 163.367
R1265 B.n430 B.n389 163.367
R1266 B.n434 B.n432 163.367
R1267 B.n438 B.n387 163.367
R1268 B.n442 B.n440 163.367
R1269 B.n446 B.n385 163.367
R1270 B.n450 B.n448 163.367
R1271 B.n454 B.n383 163.367
R1272 B.n458 B.n456 163.367
R1273 B.n462 B.n381 163.367
R1274 B.n466 B.n464 163.367
R1275 B.n470 B.n379 163.367
R1276 B.n474 B.n472 163.367
R1277 B.n478 B.n377 163.367
R1278 B.n482 B.n480 163.367
R1279 B.n486 B.n375 163.367
R1280 B.n490 B.n488 163.367
R1281 B.n497 B.n373 163.367
R1282 B.n501 B.n499 163.367
R1283 B.n505 B.n371 163.367
R1284 B.n509 B.n507 163.367
R1285 B.n513 B.n369 163.367
R1286 B.n517 B.n515 163.367
R1287 B.n522 B.n365 163.367
R1288 B.n526 B.n524 163.367
R1289 B.n530 B.n363 163.367
R1290 B.n534 B.n532 163.367
R1291 B.n538 B.n361 163.367
R1292 B.n542 B.n540 163.367
R1293 B.n546 B.n359 163.367
R1294 B.n550 B.n548 163.367
R1295 B.n554 B.n357 163.367
R1296 B.n558 B.n556 163.367
R1297 B.n562 B.n355 163.367
R1298 B.n566 B.n564 163.367
R1299 B.n570 B.n353 163.367
R1300 B.n574 B.n572 163.367
R1301 B.n578 B.n351 163.367
R1302 B.n582 B.n580 163.367
R1303 B.n586 B.n349 163.367
R1304 B.n590 B.n588 163.367
R1305 B.n594 B.n347 163.367
R1306 B.n598 B.n596 163.367
R1307 B.n602 B.n345 163.367
R1308 B.n606 B.n604 163.367
R1309 B.n610 B.n343 163.367
R1310 B.n613 B.n612 163.367
R1311 B.n615 B.n340 163.367
R1312 B.n619 B.n334 163.367
R1313 B.n627 B.n334 163.367
R1314 B.n627 B.n332 163.367
R1315 B.n631 B.n332 163.367
R1316 B.n631 B.n327 163.367
R1317 B.n640 B.n327 163.367
R1318 B.n640 B.n325 163.367
R1319 B.n644 B.n325 163.367
R1320 B.n644 B.n319 163.367
R1321 B.n652 B.n319 163.367
R1322 B.n652 B.n317 163.367
R1323 B.n657 B.n317 163.367
R1324 B.n657 B.n311 163.367
R1325 B.n665 B.n311 163.367
R1326 B.n666 B.n665 163.367
R1327 B.n666 B.n5 163.367
R1328 B.n6 B.n5 163.367
R1329 B.n7 B.n6 163.367
R1330 B.n671 B.n7 163.367
R1331 B.n671 B.n12 163.367
R1332 B.n13 B.n12 163.367
R1333 B.n14 B.n13 163.367
R1334 B.n676 B.n14 163.367
R1335 B.n676 B.n19 163.367
R1336 B.n20 B.n19 163.367
R1337 B.n21 B.n20 163.367
R1338 B.n681 B.n21 163.367
R1339 B.n681 B.n26 163.367
R1340 B.n27 B.n26 163.367
R1341 B.n28 B.n27 163.367
R1342 B.n686 B.n28 163.367
R1343 B.n686 B.n33 163.367
R1344 B.n97 B.n96 163.367
R1345 B.n101 B.n100 163.367
R1346 B.n105 B.n104 163.367
R1347 B.n109 B.n108 163.367
R1348 B.n113 B.n112 163.367
R1349 B.n117 B.n116 163.367
R1350 B.n121 B.n120 163.367
R1351 B.n125 B.n124 163.367
R1352 B.n129 B.n128 163.367
R1353 B.n133 B.n132 163.367
R1354 B.n137 B.n136 163.367
R1355 B.n141 B.n140 163.367
R1356 B.n145 B.n144 163.367
R1357 B.n149 B.n148 163.367
R1358 B.n153 B.n152 163.367
R1359 B.n157 B.n156 163.367
R1360 B.n161 B.n160 163.367
R1361 B.n165 B.n164 163.367
R1362 B.n169 B.n168 163.367
R1363 B.n173 B.n172 163.367
R1364 B.n177 B.n176 163.367
R1365 B.n181 B.n180 163.367
R1366 B.n185 B.n184 163.367
R1367 B.n189 B.n188 163.367
R1368 B.n193 B.n192 163.367
R1369 B.n197 B.n196 163.367
R1370 B.n201 B.n200 163.367
R1371 B.n205 B.n204 163.367
R1372 B.n209 B.n208 163.367
R1373 B.n213 B.n212 163.367
R1374 B.n217 B.n216 163.367
R1375 B.n221 B.n220 163.367
R1376 B.n225 B.n224 163.367
R1377 B.n229 B.n228 163.367
R1378 B.n233 B.n232 163.367
R1379 B.n237 B.n236 163.367
R1380 B.n241 B.n240 163.367
R1381 B.n245 B.n244 163.367
R1382 B.n249 B.n248 163.367
R1383 B.n253 B.n252 163.367
R1384 B.n257 B.n256 163.367
R1385 B.n261 B.n260 163.367
R1386 B.n265 B.n264 163.367
R1387 B.n269 B.n268 163.367
R1388 B.n273 B.n272 163.367
R1389 B.n277 B.n276 163.367
R1390 B.n281 B.n280 163.367
R1391 B.n285 B.n284 163.367
R1392 B.n289 B.n288 163.367
R1393 B.n293 B.n292 163.367
R1394 B.n297 B.n296 163.367
R1395 B.n301 B.n300 163.367
R1396 B.n305 B.n304 163.367
R1397 B.n307 B.n88 163.367
R1398 B.n398 B.n338 71.676
R1399 B.n402 B.n401 71.676
R1400 B.n407 B.n406 71.676
R1401 B.n410 B.n409 71.676
R1402 B.n415 B.n414 71.676
R1403 B.n418 B.n417 71.676
R1404 B.n423 B.n422 71.676
R1405 B.n426 B.n425 71.676
R1406 B.n431 B.n430 71.676
R1407 B.n434 B.n433 71.676
R1408 B.n439 B.n438 71.676
R1409 B.n442 B.n441 71.676
R1410 B.n447 B.n446 71.676
R1411 B.n450 B.n449 71.676
R1412 B.n455 B.n454 71.676
R1413 B.n458 B.n457 71.676
R1414 B.n463 B.n462 71.676
R1415 B.n466 B.n465 71.676
R1416 B.n471 B.n470 71.676
R1417 B.n474 B.n473 71.676
R1418 B.n479 B.n478 71.676
R1419 B.n482 B.n481 71.676
R1420 B.n487 B.n486 71.676
R1421 B.n490 B.n489 71.676
R1422 B.n498 B.n497 71.676
R1423 B.n501 B.n500 71.676
R1424 B.n506 B.n505 71.676
R1425 B.n509 B.n508 71.676
R1426 B.n514 B.n513 71.676
R1427 B.n517 B.n516 71.676
R1428 B.n523 B.n522 71.676
R1429 B.n526 B.n525 71.676
R1430 B.n531 B.n530 71.676
R1431 B.n534 B.n533 71.676
R1432 B.n539 B.n538 71.676
R1433 B.n542 B.n541 71.676
R1434 B.n547 B.n546 71.676
R1435 B.n550 B.n549 71.676
R1436 B.n555 B.n554 71.676
R1437 B.n558 B.n557 71.676
R1438 B.n563 B.n562 71.676
R1439 B.n566 B.n565 71.676
R1440 B.n571 B.n570 71.676
R1441 B.n574 B.n573 71.676
R1442 B.n579 B.n578 71.676
R1443 B.n582 B.n581 71.676
R1444 B.n587 B.n586 71.676
R1445 B.n590 B.n589 71.676
R1446 B.n595 B.n594 71.676
R1447 B.n598 B.n597 71.676
R1448 B.n603 B.n602 71.676
R1449 B.n606 B.n605 71.676
R1450 B.n611 B.n610 71.676
R1451 B.n614 B.n613 71.676
R1452 B.n34 B.n32 71.676
R1453 B.n97 B.n35 71.676
R1454 B.n101 B.n36 71.676
R1455 B.n105 B.n37 71.676
R1456 B.n109 B.n38 71.676
R1457 B.n113 B.n39 71.676
R1458 B.n117 B.n40 71.676
R1459 B.n121 B.n41 71.676
R1460 B.n125 B.n42 71.676
R1461 B.n129 B.n43 71.676
R1462 B.n133 B.n44 71.676
R1463 B.n137 B.n45 71.676
R1464 B.n141 B.n46 71.676
R1465 B.n145 B.n47 71.676
R1466 B.n149 B.n48 71.676
R1467 B.n153 B.n49 71.676
R1468 B.n157 B.n50 71.676
R1469 B.n161 B.n51 71.676
R1470 B.n165 B.n52 71.676
R1471 B.n169 B.n53 71.676
R1472 B.n173 B.n54 71.676
R1473 B.n177 B.n55 71.676
R1474 B.n181 B.n56 71.676
R1475 B.n185 B.n57 71.676
R1476 B.n189 B.n58 71.676
R1477 B.n193 B.n59 71.676
R1478 B.n197 B.n60 71.676
R1479 B.n201 B.n61 71.676
R1480 B.n205 B.n62 71.676
R1481 B.n209 B.n63 71.676
R1482 B.n213 B.n64 71.676
R1483 B.n217 B.n65 71.676
R1484 B.n221 B.n66 71.676
R1485 B.n225 B.n67 71.676
R1486 B.n229 B.n68 71.676
R1487 B.n233 B.n69 71.676
R1488 B.n237 B.n70 71.676
R1489 B.n241 B.n71 71.676
R1490 B.n245 B.n72 71.676
R1491 B.n249 B.n73 71.676
R1492 B.n253 B.n74 71.676
R1493 B.n257 B.n75 71.676
R1494 B.n261 B.n76 71.676
R1495 B.n265 B.n77 71.676
R1496 B.n269 B.n78 71.676
R1497 B.n273 B.n79 71.676
R1498 B.n277 B.n80 71.676
R1499 B.n281 B.n81 71.676
R1500 B.n285 B.n82 71.676
R1501 B.n289 B.n83 71.676
R1502 B.n293 B.n84 71.676
R1503 B.n297 B.n85 71.676
R1504 B.n301 B.n86 71.676
R1505 B.n305 B.n87 71.676
R1506 B.n691 B.n88 71.676
R1507 B.n691 B.n690 71.676
R1508 B.n307 B.n87 71.676
R1509 B.n304 B.n86 71.676
R1510 B.n300 B.n85 71.676
R1511 B.n296 B.n84 71.676
R1512 B.n292 B.n83 71.676
R1513 B.n288 B.n82 71.676
R1514 B.n284 B.n81 71.676
R1515 B.n280 B.n80 71.676
R1516 B.n276 B.n79 71.676
R1517 B.n272 B.n78 71.676
R1518 B.n268 B.n77 71.676
R1519 B.n264 B.n76 71.676
R1520 B.n260 B.n75 71.676
R1521 B.n256 B.n74 71.676
R1522 B.n252 B.n73 71.676
R1523 B.n248 B.n72 71.676
R1524 B.n244 B.n71 71.676
R1525 B.n240 B.n70 71.676
R1526 B.n236 B.n69 71.676
R1527 B.n232 B.n68 71.676
R1528 B.n228 B.n67 71.676
R1529 B.n224 B.n66 71.676
R1530 B.n220 B.n65 71.676
R1531 B.n216 B.n64 71.676
R1532 B.n212 B.n63 71.676
R1533 B.n208 B.n62 71.676
R1534 B.n204 B.n61 71.676
R1535 B.n200 B.n60 71.676
R1536 B.n196 B.n59 71.676
R1537 B.n192 B.n58 71.676
R1538 B.n188 B.n57 71.676
R1539 B.n184 B.n56 71.676
R1540 B.n180 B.n55 71.676
R1541 B.n176 B.n54 71.676
R1542 B.n172 B.n53 71.676
R1543 B.n168 B.n52 71.676
R1544 B.n164 B.n51 71.676
R1545 B.n160 B.n50 71.676
R1546 B.n156 B.n49 71.676
R1547 B.n152 B.n48 71.676
R1548 B.n148 B.n47 71.676
R1549 B.n144 B.n46 71.676
R1550 B.n140 B.n45 71.676
R1551 B.n136 B.n44 71.676
R1552 B.n132 B.n43 71.676
R1553 B.n128 B.n42 71.676
R1554 B.n124 B.n41 71.676
R1555 B.n120 B.n40 71.676
R1556 B.n116 B.n39 71.676
R1557 B.n112 B.n38 71.676
R1558 B.n108 B.n37 71.676
R1559 B.n104 B.n36 71.676
R1560 B.n100 B.n35 71.676
R1561 B.n96 B.n34 71.676
R1562 B.n399 B.n398 71.676
R1563 B.n401 B.n395 71.676
R1564 B.n408 B.n407 71.676
R1565 B.n409 B.n393 71.676
R1566 B.n416 B.n415 71.676
R1567 B.n417 B.n391 71.676
R1568 B.n424 B.n423 71.676
R1569 B.n425 B.n389 71.676
R1570 B.n432 B.n431 71.676
R1571 B.n433 B.n387 71.676
R1572 B.n440 B.n439 71.676
R1573 B.n441 B.n385 71.676
R1574 B.n448 B.n447 71.676
R1575 B.n449 B.n383 71.676
R1576 B.n456 B.n455 71.676
R1577 B.n457 B.n381 71.676
R1578 B.n464 B.n463 71.676
R1579 B.n465 B.n379 71.676
R1580 B.n472 B.n471 71.676
R1581 B.n473 B.n377 71.676
R1582 B.n480 B.n479 71.676
R1583 B.n481 B.n375 71.676
R1584 B.n488 B.n487 71.676
R1585 B.n489 B.n373 71.676
R1586 B.n499 B.n498 71.676
R1587 B.n500 B.n371 71.676
R1588 B.n507 B.n506 71.676
R1589 B.n508 B.n369 71.676
R1590 B.n515 B.n514 71.676
R1591 B.n516 B.n365 71.676
R1592 B.n524 B.n523 71.676
R1593 B.n525 B.n363 71.676
R1594 B.n532 B.n531 71.676
R1595 B.n533 B.n361 71.676
R1596 B.n540 B.n539 71.676
R1597 B.n541 B.n359 71.676
R1598 B.n548 B.n547 71.676
R1599 B.n549 B.n357 71.676
R1600 B.n556 B.n555 71.676
R1601 B.n557 B.n355 71.676
R1602 B.n564 B.n563 71.676
R1603 B.n565 B.n353 71.676
R1604 B.n572 B.n571 71.676
R1605 B.n573 B.n351 71.676
R1606 B.n580 B.n579 71.676
R1607 B.n581 B.n349 71.676
R1608 B.n588 B.n587 71.676
R1609 B.n589 B.n347 71.676
R1610 B.n596 B.n595 71.676
R1611 B.n597 B.n345 71.676
R1612 B.n604 B.n603 71.676
R1613 B.n605 B.n343 71.676
R1614 B.n612 B.n611 71.676
R1615 B.n615 B.n614 71.676
R1616 B.n620 B.n339 71.3195
R1617 B.n693 B.n692 71.3195
R1618 B.n519 B.n367 59.5399
R1619 B.n495 B.n494 59.5399
R1620 B.n94 B.n93 59.5399
R1621 B.n91 B.n90 59.5399
R1622 B.n620 B.n335 37.021
R1623 B.n626 B.n335 37.021
R1624 B.n626 B.n331 37.021
R1625 B.n633 B.n331 37.021
R1626 B.n633 B.n632 37.021
R1627 B.n639 B.n324 37.021
R1628 B.n645 B.n324 37.021
R1629 B.n645 B.n320 37.021
R1630 B.n651 B.n320 37.021
R1631 B.n651 B.n316 37.021
R1632 B.n658 B.n316 37.021
R1633 B.n664 B.n312 37.021
R1634 B.n664 B.n4 37.021
R1635 B.n725 B.n4 37.021
R1636 B.n725 B.n724 37.021
R1637 B.n724 B.n723 37.021
R1638 B.n723 B.n8 37.021
R1639 B.n717 B.n716 37.021
R1640 B.n716 B.n715 37.021
R1641 B.n715 B.n15 37.021
R1642 B.n709 B.n15 37.021
R1643 B.n709 B.n708 37.021
R1644 B.n708 B.n707 37.021
R1645 B.n701 B.n25 37.021
R1646 B.n701 B.n700 37.021
R1647 B.n700 B.n699 37.021
R1648 B.n699 B.n29 37.021
R1649 B.n693 B.n29 37.021
R1650 B.n695 B.n31 33.8737
R1651 B.n689 B.n688 33.8737
R1652 B.n618 B.n617 33.8737
R1653 B.n622 B.n337 33.8737
R1654 B.n639 B.t3 29.9436
R1655 B.n707 B.t10 29.9436
R1656 B.n367 B.n366 26.3763
R1657 B.n494 B.n493 26.3763
R1658 B.n93 B.n92 26.3763
R1659 B.n90 B.n89 26.3763
R1660 B.t0 B.n312 22.3217
R1661 B.t1 B.n8 22.3217
R1662 B B.n727 18.0485
R1663 B.n658 B.t0 14.6998
R1664 B.n717 B.t1 14.6998
R1665 B.n95 B.n31 10.6151
R1666 B.n98 B.n95 10.6151
R1667 B.n99 B.n98 10.6151
R1668 B.n102 B.n99 10.6151
R1669 B.n103 B.n102 10.6151
R1670 B.n106 B.n103 10.6151
R1671 B.n107 B.n106 10.6151
R1672 B.n110 B.n107 10.6151
R1673 B.n111 B.n110 10.6151
R1674 B.n114 B.n111 10.6151
R1675 B.n115 B.n114 10.6151
R1676 B.n118 B.n115 10.6151
R1677 B.n119 B.n118 10.6151
R1678 B.n122 B.n119 10.6151
R1679 B.n123 B.n122 10.6151
R1680 B.n126 B.n123 10.6151
R1681 B.n127 B.n126 10.6151
R1682 B.n130 B.n127 10.6151
R1683 B.n131 B.n130 10.6151
R1684 B.n134 B.n131 10.6151
R1685 B.n135 B.n134 10.6151
R1686 B.n138 B.n135 10.6151
R1687 B.n139 B.n138 10.6151
R1688 B.n142 B.n139 10.6151
R1689 B.n143 B.n142 10.6151
R1690 B.n146 B.n143 10.6151
R1691 B.n147 B.n146 10.6151
R1692 B.n150 B.n147 10.6151
R1693 B.n151 B.n150 10.6151
R1694 B.n154 B.n151 10.6151
R1695 B.n155 B.n154 10.6151
R1696 B.n158 B.n155 10.6151
R1697 B.n159 B.n158 10.6151
R1698 B.n162 B.n159 10.6151
R1699 B.n163 B.n162 10.6151
R1700 B.n166 B.n163 10.6151
R1701 B.n167 B.n166 10.6151
R1702 B.n170 B.n167 10.6151
R1703 B.n171 B.n170 10.6151
R1704 B.n174 B.n171 10.6151
R1705 B.n175 B.n174 10.6151
R1706 B.n178 B.n175 10.6151
R1707 B.n179 B.n178 10.6151
R1708 B.n182 B.n179 10.6151
R1709 B.n183 B.n182 10.6151
R1710 B.n186 B.n183 10.6151
R1711 B.n187 B.n186 10.6151
R1712 B.n190 B.n187 10.6151
R1713 B.n191 B.n190 10.6151
R1714 B.n195 B.n194 10.6151
R1715 B.n198 B.n195 10.6151
R1716 B.n199 B.n198 10.6151
R1717 B.n202 B.n199 10.6151
R1718 B.n203 B.n202 10.6151
R1719 B.n206 B.n203 10.6151
R1720 B.n207 B.n206 10.6151
R1721 B.n210 B.n207 10.6151
R1722 B.n211 B.n210 10.6151
R1723 B.n215 B.n214 10.6151
R1724 B.n218 B.n215 10.6151
R1725 B.n219 B.n218 10.6151
R1726 B.n222 B.n219 10.6151
R1727 B.n223 B.n222 10.6151
R1728 B.n226 B.n223 10.6151
R1729 B.n227 B.n226 10.6151
R1730 B.n230 B.n227 10.6151
R1731 B.n231 B.n230 10.6151
R1732 B.n234 B.n231 10.6151
R1733 B.n235 B.n234 10.6151
R1734 B.n238 B.n235 10.6151
R1735 B.n239 B.n238 10.6151
R1736 B.n242 B.n239 10.6151
R1737 B.n243 B.n242 10.6151
R1738 B.n246 B.n243 10.6151
R1739 B.n247 B.n246 10.6151
R1740 B.n250 B.n247 10.6151
R1741 B.n251 B.n250 10.6151
R1742 B.n254 B.n251 10.6151
R1743 B.n255 B.n254 10.6151
R1744 B.n258 B.n255 10.6151
R1745 B.n259 B.n258 10.6151
R1746 B.n262 B.n259 10.6151
R1747 B.n263 B.n262 10.6151
R1748 B.n266 B.n263 10.6151
R1749 B.n267 B.n266 10.6151
R1750 B.n270 B.n267 10.6151
R1751 B.n271 B.n270 10.6151
R1752 B.n274 B.n271 10.6151
R1753 B.n275 B.n274 10.6151
R1754 B.n278 B.n275 10.6151
R1755 B.n279 B.n278 10.6151
R1756 B.n282 B.n279 10.6151
R1757 B.n283 B.n282 10.6151
R1758 B.n286 B.n283 10.6151
R1759 B.n287 B.n286 10.6151
R1760 B.n290 B.n287 10.6151
R1761 B.n291 B.n290 10.6151
R1762 B.n294 B.n291 10.6151
R1763 B.n295 B.n294 10.6151
R1764 B.n298 B.n295 10.6151
R1765 B.n299 B.n298 10.6151
R1766 B.n302 B.n299 10.6151
R1767 B.n303 B.n302 10.6151
R1768 B.n306 B.n303 10.6151
R1769 B.n308 B.n306 10.6151
R1770 B.n309 B.n308 10.6151
R1771 B.n689 B.n309 10.6151
R1772 B.n618 B.n333 10.6151
R1773 B.n628 B.n333 10.6151
R1774 B.n629 B.n628 10.6151
R1775 B.n630 B.n629 10.6151
R1776 B.n630 B.n326 10.6151
R1777 B.n641 B.n326 10.6151
R1778 B.n642 B.n641 10.6151
R1779 B.n643 B.n642 10.6151
R1780 B.n643 B.n318 10.6151
R1781 B.n653 B.n318 10.6151
R1782 B.n654 B.n653 10.6151
R1783 B.n656 B.n654 10.6151
R1784 B.n656 B.n655 10.6151
R1785 B.n655 B.n310 10.6151
R1786 B.n667 B.n310 10.6151
R1787 B.n668 B.n667 10.6151
R1788 B.n669 B.n668 10.6151
R1789 B.n670 B.n669 10.6151
R1790 B.n672 B.n670 10.6151
R1791 B.n673 B.n672 10.6151
R1792 B.n674 B.n673 10.6151
R1793 B.n675 B.n674 10.6151
R1794 B.n677 B.n675 10.6151
R1795 B.n678 B.n677 10.6151
R1796 B.n679 B.n678 10.6151
R1797 B.n680 B.n679 10.6151
R1798 B.n682 B.n680 10.6151
R1799 B.n683 B.n682 10.6151
R1800 B.n684 B.n683 10.6151
R1801 B.n685 B.n684 10.6151
R1802 B.n687 B.n685 10.6151
R1803 B.n688 B.n687 10.6151
R1804 B.n397 B.n337 10.6151
R1805 B.n397 B.n396 10.6151
R1806 B.n403 B.n396 10.6151
R1807 B.n404 B.n403 10.6151
R1808 B.n405 B.n404 10.6151
R1809 B.n405 B.n394 10.6151
R1810 B.n411 B.n394 10.6151
R1811 B.n412 B.n411 10.6151
R1812 B.n413 B.n412 10.6151
R1813 B.n413 B.n392 10.6151
R1814 B.n419 B.n392 10.6151
R1815 B.n420 B.n419 10.6151
R1816 B.n421 B.n420 10.6151
R1817 B.n421 B.n390 10.6151
R1818 B.n427 B.n390 10.6151
R1819 B.n428 B.n427 10.6151
R1820 B.n429 B.n428 10.6151
R1821 B.n429 B.n388 10.6151
R1822 B.n435 B.n388 10.6151
R1823 B.n436 B.n435 10.6151
R1824 B.n437 B.n436 10.6151
R1825 B.n437 B.n386 10.6151
R1826 B.n443 B.n386 10.6151
R1827 B.n444 B.n443 10.6151
R1828 B.n445 B.n444 10.6151
R1829 B.n445 B.n384 10.6151
R1830 B.n451 B.n384 10.6151
R1831 B.n452 B.n451 10.6151
R1832 B.n453 B.n452 10.6151
R1833 B.n453 B.n382 10.6151
R1834 B.n459 B.n382 10.6151
R1835 B.n460 B.n459 10.6151
R1836 B.n461 B.n460 10.6151
R1837 B.n461 B.n380 10.6151
R1838 B.n467 B.n380 10.6151
R1839 B.n468 B.n467 10.6151
R1840 B.n469 B.n468 10.6151
R1841 B.n469 B.n378 10.6151
R1842 B.n475 B.n378 10.6151
R1843 B.n476 B.n475 10.6151
R1844 B.n477 B.n476 10.6151
R1845 B.n477 B.n376 10.6151
R1846 B.n483 B.n376 10.6151
R1847 B.n484 B.n483 10.6151
R1848 B.n485 B.n484 10.6151
R1849 B.n485 B.n374 10.6151
R1850 B.n491 B.n374 10.6151
R1851 B.n492 B.n491 10.6151
R1852 B.n496 B.n492 10.6151
R1853 B.n502 B.n372 10.6151
R1854 B.n503 B.n502 10.6151
R1855 B.n504 B.n503 10.6151
R1856 B.n504 B.n370 10.6151
R1857 B.n510 B.n370 10.6151
R1858 B.n511 B.n510 10.6151
R1859 B.n512 B.n511 10.6151
R1860 B.n512 B.n368 10.6151
R1861 B.n518 B.n368 10.6151
R1862 B.n521 B.n520 10.6151
R1863 B.n521 B.n364 10.6151
R1864 B.n527 B.n364 10.6151
R1865 B.n528 B.n527 10.6151
R1866 B.n529 B.n528 10.6151
R1867 B.n529 B.n362 10.6151
R1868 B.n535 B.n362 10.6151
R1869 B.n536 B.n535 10.6151
R1870 B.n537 B.n536 10.6151
R1871 B.n537 B.n360 10.6151
R1872 B.n543 B.n360 10.6151
R1873 B.n544 B.n543 10.6151
R1874 B.n545 B.n544 10.6151
R1875 B.n545 B.n358 10.6151
R1876 B.n551 B.n358 10.6151
R1877 B.n552 B.n551 10.6151
R1878 B.n553 B.n552 10.6151
R1879 B.n553 B.n356 10.6151
R1880 B.n559 B.n356 10.6151
R1881 B.n560 B.n559 10.6151
R1882 B.n561 B.n560 10.6151
R1883 B.n561 B.n354 10.6151
R1884 B.n567 B.n354 10.6151
R1885 B.n568 B.n567 10.6151
R1886 B.n569 B.n568 10.6151
R1887 B.n569 B.n352 10.6151
R1888 B.n575 B.n352 10.6151
R1889 B.n576 B.n575 10.6151
R1890 B.n577 B.n576 10.6151
R1891 B.n577 B.n350 10.6151
R1892 B.n583 B.n350 10.6151
R1893 B.n584 B.n583 10.6151
R1894 B.n585 B.n584 10.6151
R1895 B.n585 B.n348 10.6151
R1896 B.n591 B.n348 10.6151
R1897 B.n592 B.n591 10.6151
R1898 B.n593 B.n592 10.6151
R1899 B.n593 B.n346 10.6151
R1900 B.n599 B.n346 10.6151
R1901 B.n600 B.n599 10.6151
R1902 B.n601 B.n600 10.6151
R1903 B.n601 B.n344 10.6151
R1904 B.n607 B.n344 10.6151
R1905 B.n608 B.n607 10.6151
R1906 B.n609 B.n608 10.6151
R1907 B.n609 B.n342 10.6151
R1908 B.n342 B.n341 10.6151
R1909 B.n616 B.n341 10.6151
R1910 B.n617 B.n616 10.6151
R1911 B.n623 B.n622 10.6151
R1912 B.n624 B.n623 10.6151
R1913 B.n624 B.n329 10.6151
R1914 B.n635 B.n329 10.6151
R1915 B.n636 B.n635 10.6151
R1916 B.n637 B.n636 10.6151
R1917 B.n637 B.n322 10.6151
R1918 B.n647 B.n322 10.6151
R1919 B.n648 B.n647 10.6151
R1920 B.n649 B.n648 10.6151
R1921 B.n649 B.n314 10.6151
R1922 B.n660 B.n314 10.6151
R1923 B.n661 B.n660 10.6151
R1924 B.n662 B.n661 10.6151
R1925 B.n662 B.n0 10.6151
R1926 B.n721 B.n1 10.6151
R1927 B.n721 B.n720 10.6151
R1928 B.n720 B.n719 10.6151
R1929 B.n719 B.n10 10.6151
R1930 B.n713 B.n10 10.6151
R1931 B.n713 B.n712 10.6151
R1932 B.n712 B.n711 10.6151
R1933 B.n711 B.n17 10.6151
R1934 B.n705 B.n17 10.6151
R1935 B.n705 B.n704 10.6151
R1936 B.n704 B.n703 10.6151
R1937 B.n703 B.n23 10.6151
R1938 B.n697 B.n23 10.6151
R1939 B.n697 B.n696 10.6151
R1940 B.n696 B.n695 10.6151
R1941 B.n191 B.n94 8.74196
R1942 B.n214 B.n91 8.74196
R1943 B.n496 B.n495 8.74196
R1944 B.n520 B.n519 8.74196
R1945 B.n632 B.t3 7.07796
R1946 B.n25 B.t10 7.07796
R1947 B.n727 B.n0 2.81026
R1948 B.n727 B.n1 2.81026
R1949 B.n194 B.n94 1.87367
R1950 B.n211 B.n91 1.87367
R1951 B.n495 B.n372 1.87367
R1952 B.n519 B.n518 1.87367
R1953 VN VN.t0 591.631
R1954 VN VN.t1 548.59
R1955 VDD2.n157 VDD2.n81 289.615
R1956 VDD2.n76 VDD2.n0 289.615
R1957 VDD2.n158 VDD2.n157 185
R1958 VDD2.n156 VDD2.n155 185
R1959 VDD2.n85 VDD2.n84 185
R1960 VDD2.n150 VDD2.n149 185
R1961 VDD2.n148 VDD2.n147 185
R1962 VDD2.n89 VDD2.n88 185
R1963 VDD2.n142 VDD2.n141 185
R1964 VDD2.n140 VDD2.n139 185
R1965 VDD2.n93 VDD2.n92 185
R1966 VDD2.n134 VDD2.n133 185
R1967 VDD2.n132 VDD2.n131 185
R1968 VDD2.n130 VDD2.n96 185
R1969 VDD2.n100 VDD2.n97 185
R1970 VDD2.n125 VDD2.n124 185
R1971 VDD2.n123 VDD2.n122 185
R1972 VDD2.n102 VDD2.n101 185
R1973 VDD2.n117 VDD2.n116 185
R1974 VDD2.n115 VDD2.n114 185
R1975 VDD2.n106 VDD2.n105 185
R1976 VDD2.n109 VDD2.n108 185
R1977 VDD2.n27 VDD2.n26 185
R1978 VDD2.n24 VDD2.n23 185
R1979 VDD2.n33 VDD2.n32 185
R1980 VDD2.n35 VDD2.n34 185
R1981 VDD2.n20 VDD2.n19 185
R1982 VDD2.n41 VDD2.n40 185
R1983 VDD2.n44 VDD2.n43 185
R1984 VDD2.n42 VDD2.n16 185
R1985 VDD2.n49 VDD2.n15 185
R1986 VDD2.n51 VDD2.n50 185
R1987 VDD2.n53 VDD2.n52 185
R1988 VDD2.n12 VDD2.n11 185
R1989 VDD2.n59 VDD2.n58 185
R1990 VDD2.n61 VDD2.n60 185
R1991 VDD2.n8 VDD2.n7 185
R1992 VDD2.n67 VDD2.n66 185
R1993 VDD2.n69 VDD2.n68 185
R1994 VDD2.n4 VDD2.n3 185
R1995 VDD2.n75 VDD2.n74 185
R1996 VDD2.n77 VDD2.n76 185
R1997 VDD2.t1 VDD2.n107 149.524
R1998 VDD2.t0 VDD2.n25 149.524
R1999 VDD2.n157 VDD2.n156 104.615
R2000 VDD2.n156 VDD2.n84 104.615
R2001 VDD2.n149 VDD2.n84 104.615
R2002 VDD2.n149 VDD2.n148 104.615
R2003 VDD2.n148 VDD2.n88 104.615
R2004 VDD2.n141 VDD2.n88 104.615
R2005 VDD2.n141 VDD2.n140 104.615
R2006 VDD2.n140 VDD2.n92 104.615
R2007 VDD2.n133 VDD2.n92 104.615
R2008 VDD2.n133 VDD2.n132 104.615
R2009 VDD2.n132 VDD2.n96 104.615
R2010 VDD2.n100 VDD2.n96 104.615
R2011 VDD2.n124 VDD2.n100 104.615
R2012 VDD2.n124 VDD2.n123 104.615
R2013 VDD2.n123 VDD2.n101 104.615
R2014 VDD2.n116 VDD2.n101 104.615
R2015 VDD2.n116 VDD2.n115 104.615
R2016 VDD2.n115 VDD2.n105 104.615
R2017 VDD2.n108 VDD2.n105 104.615
R2018 VDD2.n26 VDD2.n23 104.615
R2019 VDD2.n33 VDD2.n23 104.615
R2020 VDD2.n34 VDD2.n33 104.615
R2021 VDD2.n34 VDD2.n19 104.615
R2022 VDD2.n41 VDD2.n19 104.615
R2023 VDD2.n43 VDD2.n41 104.615
R2024 VDD2.n43 VDD2.n42 104.615
R2025 VDD2.n42 VDD2.n15 104.615
R2026 VDD2.n51 VDD2.n15 104.615
R2027 VDD2.n52 VDD2.n51 104.615
R2028 VDD2.n52 VDD2.n11 104.615
R2029 VDD2.n59 VDD2.n11 104.615
R2030 VDD2.n60 VDD2.n59 104.615
R2031 VDD2.n60 VDD2.n7 104.615
R2032 VDD2.n67 VDD2.n7 104.615
R2033 VDD2.n68 VDD2.n67 104.615
R2034 VDD2.n68 VDD2.n3 104.615
R2035 VDD2.n75 VDD2.n3 104.615
R2036 VDD2.n76 VDD2.n75 104.615
R2037 VDD2.n162 VDD2.n80 85.9937
R2038 VDD2.n108 VDD2.t1 52.3082
R2039 VDD2.n26 VDD2.t0 52.3082
R2040 VDD2.n162 VDD2.n161 47.1187
R2041 VDD2.n131 VDD2.n130 13.1884
R2042 VDD2.n50 VDD2.n49 13.1884
R2043 VDD2.n134 VDD2.n95 12.8005
R2044 VDD2.n129 VDD2.n97 12.8005
R2045 VDD2.n48 VDD2.n16 12.8005
R2046 VDD2.n53 VDD2.n14 12.8005
R2047 VDD2.n135 VDD2.n93 12.0247
R2048 VDD2.n126 VDD2.n125 12.0247
R2049 VDD2.n45 VDD2.n44 12.0247
R2050 VDD2.n54 VDD2.n12 12.0247
R2051 VDD2.n139 VDD2.n138 11.249
R2052 VDD2.n122 VDD2.n99 11.249
R2053 VDD2.n40 VDD2.n18 11.249
R2054 VDD2.n58 VDD2.n57 11.249
R2055 VDD2.n142 VDD2.n91 10.4732
R2056 VDD2.n121 VDD2.n102 10.4732
R2057 VDD2.n39 VDD2.n20 10.4732
R2058 VDD2.n61 VDD2.n10 10.4732
R2059 VDD2.n109 VDD2.n107 10.2747
R2060 VDD2.n27 VDD2.n25 10.2747
R2061 VDD2.n143 VDD2.n89 9.69747
R2062 VDD2.n118 VDD2.n117 9.69747
R2063 VDD2.n36 VDD2.n35 9.69747
R2064 VDD2.n62 VDD2.n8 9.69747
R2065 VDD2.n161 VDD2.n160 9.45567
R2066 VDD2.n80 VDD2.n79 9.45567
R2067 VDD2.n83 VDD2.n82 9.3005
R2068 VDD2.n154 VDD2.n153 9.3005
R2069 VDD2.n152 VDD2.n151 9.3005
R2070 VDD2.n87 VDD2.n86 9.3005
R2071 VDD2.n146 VDD2.n145 9.3005
R2072 VDD2.n144 VDD2.n143 9.3005
R2073 VDD2.n91 VDD2.n90 9.3005
R2074 VDD2.n138 VDD2.n137 9.3005
R2075 VDD2.n136 VDD2.n135 9.3005
R2076 VDD2.n95 VDD2.n94 9.3005
R2077 VDD2.n129 VDD2.n128 9.3005
R2078 VDD2.n127 VDD2.n126 9.3005
R2079 VDD2.n99 VDD2.n98 9.3005
R2080 VDD2.n121 VDD2.n120 9.3005
R2081 VDD2.n119 VDD2.n118 9.3005
R2082 VDD2.n104 VDD2.n103 9.3005
R2083 VDD2.n113 VDD2.n112 9.3005
R2084 VDD2.n111 VDD2.n110 9.3005
R2085 VDD2.n160 VDD2.n159 9.3005
R2086 VDD2.n73 VDD2.n72 9.3005
R2087 VDD2.n2 VDD2.n1 9.3005
R2088 VDD2.n79 VDD2.n78 9.3005
R2089 VDD2.n6 VDD2.n5 9.3005
R2090 VDD2.n65 VDD2.n64 9.3005
R2091 VDD2.n63 VDD2.n62 9.3005
R2092 VDD2.n10 VDD2.n9 9.3005
R2093 VDD2.n57 VDD2.n56 9.3005
R2094 VDD2.n55 VDD2.n54 9.3005
R2095 VDD2.n14 VDD2.n13 9.3005
R2096 VDD2.n29 VDD2.n28 9.3005
R2097 VDD2.n31 VDD2.n30 9.3005
R2098 VDD2.n22 VDD2.n21 9.3005
R2099 VDD2.n37 VDD2.n36 9.3005
R2100 VDD2.n39 VDD2.n38 9.3005
R2101 VDD2.n18 VDD2.n17 9.3005
R2102 VDD2.n46 VDD2.n45 9.3005
R2103 VDD2.n48 VDD2.n47 9.3005
R2104 VDD2.n71 VDD2.n70 9.3005
R2105 VDD2.n161 VDD2.n81 8.92171
R2106 VDD2.n147 VDD2.n146 8.92171
R2107 VDD2.n114 VDD2.n104 8.92171
R2108 VDD2.n32 VDD2.n22 8.92171
R2109 VDD2.n66 VDD2.n65 8.92171
R2110 VDD2.n80 VDD2.n0 8.92171
R2111 VDD2.n159 VDD2.n158 8.14595
R2112 VDD2.n150 VDD2.n87 8.14595
R2113 VDD2.n113 VDD2.n106 8.14595
R2114 VDD2.n31 VDD2.n24 8.14595
R2115 VDD2.n69 VDD2.n6 8.14595
R2116 VDD2.n78 VDD2.n77 8.14595
R2117 VDD2.n155 VDD2.n83 7.3702
R2118 VDD2.n151 VDD2.n85 7.3702
R2119 VDD2.n110 VDD2.n109 7.3702
R2120 VDD2.n28 VDD2.n27 7.3702
R2121 VDD2.n70 VDD2.n4 7.3702
R2122 VDD2.n74 VDD2.n2 7.3702
R2123 VDD2.n155 VDD2.n154 6.59444
R2124 VDD2.n154 VDD2.n85 6.59444
R2125 VDD2.n73 VDD2.n4 6.59444
R2126 VDD2.n74 VDD2.n73 6.59444
R2127 VDD2.n158 VDD2.n83 5.81868
R2128 VDD2.n151 VDD2.n150 5.81868
R2129 VDD2.n110 VDD2.n106 5.81868
R2130 VDD2.n28 VDD2.n24 5.81868
R2131 VDD2.n70 VDD2.n69 5.81868
R2132 VDD2.n77 VDD2.n2 5.81868
R2133 VDD2.n159 VDD2.n81 5.04292
R2134 VDD2.n147 VDD2.n87 5.04292
R2135 VDD2.n114 VDD2.n113 5.04292
R2136 VDD2.n32 VDD2.n31 5.04292
R2137 VDD2.n66 VDD2.n6 5.04292
R2138 VDD2.n78 VDD2.n0 5.04292
R2139 VDD2.n146 VDD2.n89 4.26717
R2140 VDD2.n117 VDD2.n104 4.26717
R2141 VDD2.n35 VDD2.n22 4.26717
R2142 VDD2.n65 VDD2.n8 4.26717
R2143 VDD2.n143 VDD2.n142 3.49141
R2144 VDD2.n118 VDD2.n102 3.49141
R2145 VDD2.n36 VDD2.n20 3.49141
R2146 VDD2.n62 VDD2.n61 3.49141
R2147 VDD2.n29 VDD2.n25 2.84303
R2148 VDD2.n111 VDD2.n107 2.84303
R2149 VDD2.n139 VDD2.n91 2.71565
R2150 VDD2.n122 VDD2.n121 2.71565
R2151 VDD2.n40 VDD2.n39 2.71565
R2152 VDD2.n58 VDD2.n10 2.71565
R2153 VDD2.n138 VDD2.n93 1.93989
R2154 VDD2.n125 VDD2.n99 1.93989
R2155 VDD2.n44 VDD2.n18 1.93989
R2156 VDD2.n57 VDD2.n12 1.93989
R2157 VDD2.n135 VDD2.n134 1.16414
R2158 VDD2.n126 VDD2.n97 1.16414
R2159 VDD2.n45 VDD2.n16 1.16414
R2160 VDD2.n54 VDD2.n53 1.16414
R2161 VDD2.n131 VDD2.n95 0.388379
R2162 VDD2.n130 VDD2.n129 0.388379
R2163 VDD2.n49 VDD2.n48 0.388379
R2164 VDD2.n50 VDD2.n14 0.388379
R2165 VDD2 VDD2.n162 0.351793
R2166 VDD2.n160 VDD2.n82 0.155672
R2167 VDD2.n153 VDD2.n82 0.155672
R2168 VDD2.n153 VDD2.n152 0.155672
R2169 VDD2.n152 VDD2.n86 0.155672
R2170 VDD2.n145 VDD2.n86 0.155672
R2171 VDD2.n145 VDD2.n144 0.155672
R2172 VDD2.n144 VDD2.n90 0.155672
R2173 VDD2.n137 VDD2.n90 0.155672
R2174 VDD2.n137 VDD2.n136 0.155672
R2175 VDD2.n136 VDD2.n94 0.155672
R2176 VDD2.n128 VDD2.n94 0.155672
R2177 VDD2.n128 VDD2.n127 0.155672
R2178 VDD2.n127 VDD2.n98 0.155672
R2179 VDD2.n120 VDD2.n98 0.155672
R2180 VDD2.n120 VDD2.n119 0.155672
R2181 VDD2.n119 VDD2.n103 0.155672
R2182 VDD2.n112 VDD2.n103 0.155672
R2183 VDD2.n112 VDD2.n111 0.155672
R2184 VDD2.n30 VDD2.n29 0.155672
R2185 VDD2.n30 VDD2.n21 0.155672
R2186 VDD2.n37 VDD2.n21 0.155672
R2187 VDD2.n38 VDD2.n37 0.155672
R2188 VDD2.n38 VDD2.n17 0.155672
R2189 VDD2.n46 VDD2.n17 0.155672
R2190 VDD2.n47 VDD2.n46 0.155672
R2191 VDD2.n47 VDD2.n13 0.155672
R2192 VDD2.n55 VDD2.n13 0.155672
R2193 VDD2.n56 VDD2.n55 0.155672
R2194 VDD2.n56 VDD2.n9 0.155672
R2195 VDD2.n63 VDD2.n9 0.155672
R2196 VDD2.n64 VDD2.n63 0.155672
R2197 VDD2.n64 VDD2.n5 0.155672
R2198 VDD2.n71 VDD2.n5 0.155672
R2199 VDD2.n72 VDD2.n71 0.155672
R2200 VDD2.n72 VDD2.n1 0.155672
R2201 VDD2.n79 VDD2.n1 0.155672
C0 VN VP 5.24966f
C1 VDD1 VN 0.148739f
C2 VN VDD2 2.74607f
C3 VP VTAIL 2.17628f
C4 VDD1 VTAIL 6.23291f
C5 VDD2 VTAIL 6.26876f
C6 VDD1 VP 2.8617f
C7 VP VDD2 0.26911f
C8 VN VTAIL 2.16167f
C9 VDD1 VDD2 0.495903f
C10 VDD2 B 4.400015f
C11 VDD1 B 7.05838f
C12 VTAIL B 7.673086f
C13 VN B 9.8992f
C14 VP B 4.627516f
C15 VDD2.n0 B 0.029529f
C16 VDD2.n1 B 0.020326f
C17 VDD2.n2 B 0.010922f
C18 VDD2.n3 B 0.025816f
C19 VDD2.n4 B 0.011565f
C20 VDD2.n5 B 0.020326f
C21 VDD2.n6 B 0.010922f
C22 VDD2.n7 B 0.025816f
C23 VDD2.n8 B 0.011565f
C24 VDD2.n9 B 0.020326f
C25 VDD2.n10 B 0.010922f
C26 VDD2.n11 B 0.025816f
C27 VDD2.n12 B 0.011565f
C28 VDD2.n13 B 0.020326f
C29 VDD2.n14 B 0.010922f
C30 VDD2.n15 B 0.025816f
C31 VDD2.n16 B 0.011565f
C32 VDD2.n17 B 0.020326f
C33 VDD2.n18 B 0.010922f
C34 VDD2.n19 B 0.025816f
C35 VDD2.n20 B 0.011565f
C36 VDD2.n21 B 0.020326f
C37 VDD2.n22 B 0.010922f
C38 VDD2.n23 B 0.025816f
C39 VDD2.n24 B 0.011565f
C40 VDD2.n25 B 0.169253f
C41 VDD2.t0 B 0.04392f
C42 VDD2.n26 B 0.019362f
C43 VDD2.n27 B 0.01825f
C44 VDD2.n28 B 0.010922f
C45 VDD2.n29 B 1.28847f
C46 VDD2.n30 B 0.020326f
C47 VDD2.n31 B 0.010922f
C48 VDD2.n32 B 0.011565f
C49 VDD2.n33 B 0.025816f
C50 VDD2.n34 B 0.025816f
C51 VDD2.n35 B 0.011565f
C52 VDD2.n36 B 0.010922f
C53 VDD2.n37 B 0.020326f
C54 VDD2.n38 B 0.020326f
C55 VDD2.n39 B 0.010922f
C56 VDD2.n40 B 0.011565f
C57 VDD2.n41 B 0.025816f
C58 VDD2.n42 B 0.025816f
C59 VDD2.n43 B 0.025816f
C60 VDD2.n44 B 0.011565f
C61 VDD2.n45 B 0.010922f
C62 VDD2.n46 B 0.020326f
C63 VDD2.n47 B 0.020326f
C64 VDD2.n48 B 0.010922f
C65 VDD2.n49 B 0.011243f
C66 VDD2.n50 B 0.011243f
C67 VDD2.n51 B 0.025816f
C68 VDD2.n52 B 0.025816f
C69 VDD2.n53 B 0.011565f
C70 VDD2.n54 B 0.010922f
C71 VDD2.n55 B 0.020326f
C72 VDD2.n56 B 0.020326f
C73 VDD2.n57 B 0.010922f
C74 VDD2.n58 B 0.011565f
C75 VDD2.n59 B 0.025816f
C76 VDD2.n60 B 0.025816f
C77 VDD2.n61 B 0.011565f
C78 VDD2.n62 B 0.010922f
C79 VDD2.n63 B 0.020326f
C80 VDD2.n64 B 0.020326f
C81 VDD2.n65 B 0.010922f
C82 VDD2.n66 B 0.011565f
C83 VDD2.n67 B 0.025816f
C84 VDD2.n68 B 0.025816f
C85 VDD2.n69 B 0.011565f
C86 VDD2.n70 B 0.010922f
C87 VDD2.n71 B 0.020326f
C88 VDD2.n72 B 0.020326f
C89 VDD2.n73 B 0.010922f
C90 VDD2.n74 B 0.011565f
C91 VDD2.n75 B 0.025816f
C92 VDD2.n76 B 0.057585f
C93 VDD2.n77 B 0.011565f
C94 VDD2.n78 B 0.010922f
C95 VDD2.n79 B 0.044483f
C96 VDD2.n80 B 0.610148f
C97 VDD2.n81 B 0.029529f
C98 VDD2.n82 B 0.020326f
C99 VDD2.n83 B 0.010922f
C100 VDD2.n84 B 0.025816f
C101 VDD2.n85 B 0.011565f
C102 VDD2.n86 B 0.020326f
C103 VDD2.n87 B 0.010922f
C104 VDD2.n88 B 0.025816f
C105 VDD2.n89 B 0.011565f
C106 VDD2.n90 B 0.020326f
C107 VDD2.n91 B 0.010922f
C108 VDD2.n92 B 0.025816f
C109 VDD2.n93 B 0.011565f
C110 VDD2.n94 B 0.020326f
C111 VDD2.n95 B 0.010922f
C112 VDD2.n96 B 0.025816f
C113 VDD2.n97 B 0.011565f
C114 VDD2.n98 B 0.020326f
C115 VDD2.n99 B 0.010922f
C116 VDD2.n100 B 0.025816f
C117 VDD2.n101 B 0.025816f
C118 VDD2.n102 B 0.011565f
C119 VDD2.n103 B 0.020326f
C120 VDD2.n104 B 0.010922f
C121 VDD2.n105 B 0.025816f
C122 VDD2.n106 B 0.011565f
C123 VDD2.n107 B 0.169253f
C124 VDD2.t1 B 0.04392f
C125 VDD2.n108 B 0.019362f
C126 VDD2.n109 B 0.01825f
C127 VDD2.n110 B 0.010922f
C128 VDD2.n111 B 1.28847f
C129 VDD2.n112 B 0.020326f
C130 VDD2.n113 B 0.010922f
C131 VDD2.n114 B 0.011565f
C132 VDD2.n115 B 0.025816f
C133 VDD2.n116 B 0.025816f
C134 VDD2.n117 B 0.011565f
C135 VDD2.n118 B 0.010922f
C136 VDD2.n119 B 0.020326f
C137 VDD2.n120 B 0.020326f
C138 VDD2.n121 B 0.010922f
C139 VDD2.n122 B 0.011565f
C140 VDD2.n123 B 0.025816f
C141 VDD2.n124 B 0.025816f
C142 VDD2.n125 B 0.011565f
C143 VDD2.n126 B 0.010922f
C144 VDD2.n127 B 0.020326f
C145 VDD2.n128 B 0.020326f
C146 VDD2.n129 B 0.010922f
C147 VDD2.n130 B 0.011243f
C148 VDD2.n131 B 0.011243f
C149 VDD2.n132 B 0.025816f
C150 VDD2.n133 B 0.025816f
C151 VDD2.n134 B 0.011565f
C152 VDD2.n135 B 0.010922f
C153 VDD2.n136 B 0.020326f
C154 VDD2.n137 B 0.020326f
C155 VDD2.n138 B 0.010922f
C156 VDD2.n139 B 0.011565f
C157 VDD2.n140 B 0.025816f
C158 VDD2.n141 B 0.025816f
C159 VDD2.n142 B 0.011565f
C160 VDD2.n143 B 0.010922f
C161 VDD2.n144 B 0.020326f
C162 VDD2.n145 B 0.020326f
C163 VDD2.n146 B 0.010922f
C164 VDD2.n147 B 0.011565f
C165 VDD2.n148 B 0.025816f
C166 VDD2.n149 B 0.025816f
C167 VDD2.n150 B 0.011565f
C168 VDD2.n151 B 0.010922f
C169 VDD2.n152 B 0.020326f
C170 VDD2.n153 B 0.020326f
C171 VDD2.n154 B 0.010922f
C172 VDD2.n155 B 0.011565f
C173 VDD2.n156 B 0.025816f
C174 VDD2.n157 B 0.057585f
C175 VDD2.n158 B 0.011565f
C176 VDD2.n159 B 0.010922f
C177 VDD2.n160 B 0.044483f
C178 VDD2.n161 B 0.046372f
C179 VDD2.n162 B 2.46615f
C180 VN.t1 B 2.35361f
C181 VN.t0 B 2.54829f
C182 VDD1.n0 B 0.029611f
C183 VDD1.n1 B 0.020382f
C184 VDD1.n2 B 0.010952f
C185 VDD1.n3 B 0.025887f
C186 VDD1.n4 B 0.011596f
C187 VDD1.n5 B 0.020382f
C188 VDD1.n6 B 0.010952f
C189 VDD1.n7 B 0.025887f
C190 VDD1.n8 B 0.011596f
C191 VDD1.n9 B 0.020382f
C192 VDD1.n10 B 0.010952f
C193 VDD1.n11 B 0.025887f
C194 VDD1.n12 B 0.011596f
C195 VDD1.n13 B 0.020382f
C196 VDD1.n14 B 0.010952f
C197 VDD1.n15 B 0.025887f
C198 VDD1.n16 B 0.011596f
C199 VDD1.n17 B 0.020382f
C200 VDD1.n18 B 0.010952f
C201 VDD1.n19 B 0.025887f
C202 VDD1.n20 B 0.025887f
C203 VDD1.n21 B 0.011596f
C204 VDD1.n22 B 0.020382f
C205 VDD1.n23 B 0.010952f
C206 VDD1.n24 B 0.025887f
C207 VDD1.n25 B 0.011596f
C208 VDD1.n26 B 0.169718f
C209 VDD1.t0 B 0.04404f
C210 VDD1.n27 B 0.019415f
C211 VDD1.n28 B 0.0183f
C212 VDD1.n29 B 0.010952f
C213 VDD1.n30 B 1.29201f
C214 VDD1.n31 B 0.020382f
C215 VDD1.n32 B 0.010952f
C216 VDD1.n33 B 0.011596f
C217 VDD1.n34 B 0.025887f
C218 VDD1.n35 B 0.025887f
C219 VDD1.n36 B 0.011596f
C220 VDD1.n37 B 0.010952f
C221 VDD1.n38 B 0.020382f
C222 VDD1.n39 B 0.020382f
C223 VDD1.n40 B 0.010952f
C224 VDD1.n41 B 0.011596f
C225 VDD1.n42 B 0.025887f
C226 VDD1.n43 B 0.025887f
C227 VDD1.n44 B 0.011596f
C228 VDD1.n45 B 0.010952f
C229 VDD1.n46 B 0.020382f
C230 VDD1.n47 B 0.020382f
C231 VDD1.n48 B 0.010952f
C232 VDD1.n49 B 0.011274f
C233 VDD1.n50 B 0.011274f
C234 VDD1.n51 B 0.025887f
C235 VDD1.n52 B 0.025887f
C236 VDD1.n53 B 0.011596f
C237 VDD1.n54 B 0.010952f
C238 VDD1.n55 B 0.020382f
C239 VDD1.n56 B 0.020382f
C240 VDD1.n57 B 0.010952f
C241 VDD1.n58 B 0.011596f
C242 VDD1.n59 B 0.025887f
C243 VDD1.n60 B 0.025887f
C244 VDD1.n61 B 0.011596f
C245 VDD1.n62 B 0.010952f
C246 VDD1.n63 B 0.020382f
C247 VDD1.n64 B 0.020382f
C248 VDD1.n65 B 0.010952f
C249 VDD1.n66 B 0.011596f
C250 VDD1.n67 B 0.025887f
C251 VDD1.n68 B 0.025887f
C252 VDD1.n69 B 0.011596f
C253 VDD1.n70 B 0.010952f
C254 VDD1.n71 B 0.020382f
C255 VDD1.n72 B 0.020382f
C256 VDD1.n73 B 0.010952f
C257 VDD1.n74 B 0.011596f
C258 VDD1.n75 B 0.025887f
C259 VDD1.n76 B 0.057743f
C260 VDD1.n77 B 0.011596f
C261 VDD1.n78 B 0.010952f
C262 VDD1.n79 B 0.044605f
C263 VDD1.n80 B 0.04695f
C264 VDD1.n81 B 0.029611f
C265 VDD1.n82 B 0.020382f
C266 VDD1.n83 B 0.010952f
C267 VDD1.n84 B 0.025887f
C268 VDD1.n85 B 0.011596f
C269 VDD1.n86 B 0.020382f
C270 VDD1.n87 B 0.010952f
C271 VDD1.n88 B 0.025887f
C272 VDD1.n89 B 0.011596f
C273 VDD1.n90 B 0.020382f
C274 VDD1.n91 B 0.010952f
C275 VDD1.n92 B 0.025887f
C276 VDD1.n93 B 0.011596f
C277 VDD1.n94 B 0.020382f
C278 VDD1.n95 B 0.010952f
C279 VDD1.n96 B 0.025887f
C280 VDD1.n97 B 0.011596f
C281 VDD1.n98 B 0.020382f
C282 VDD1.n99 B 0.010952f
C283 VDD1.n100 B 0.025887f
C284 VDD1.n101 B 0.011596f
C285 VDD1.n102 B 0.020382f
C286 VDD1.n103 B 0.010952f
C287 VDD1.n104 B 0.025887f
C288 VDD1.n105 B 0.011596f
C289 VDD1.n106 B 0.169718f
C290 VDD1.t1 B 0.04404f
C291 VDD1.n107 B 0.019415f
C292 VDD1.n108 B 0.0183f
C293 VDD1.n109 B 0.010952f
C294 VDD1.n110 B 1.29201f
C295 VDD1.n111 B 0.020382f
C296 VDD1.n112 B 0.010952f
C297 VDD1.n113 B 0.011596f
C298 VDD1.n114 B 0.025887f
C299 VDD1.n115 B 0.025887f
C300 VDD1.n116 B 0.011596f
C301 VDD1.n117 B 0.010952f
C302 VDD1.n118 B 0.020382f
C303 VDD1.n119 B 0.020382f
C304 VDD1.n120 B 0.010952f
C305 VDD1.n121 B 0.011596f
C306 VDD1.n122 B 0.025887f
C307 VDD1.n123 B 0.025887f
C308 VDD1.n124 B 0.025887f
C309 VDD1.n125 B 0.011596f
C310 VDD1.n126 B 0.010952f
C311 VDD1.n127 B 0.020382f
C312 VDD1.n128 B 0.020382f
C313 VDD1.n129 B 0.010952f
C314 VDD1.n130 B 0.011274f
C315 VDD1.n131 B 0.011274f
C316 VDD1.n132 B 0.025887f
C317 VDD1.n133 B 0.025887f
C318 VDD1.n134 B 0.011596f
C319 VDD1.n135 B 0.010952f
C320 VDD1.n136 B 0.020382f
C321 VDD1.n137 B 0.020382f
C322 VDD1.n138 B 0.010952f
C323 VDD1.n139 B 0.011596f
C324 VDD1.n140 B 0.025887f
C325 VDD1.n141 B 0.025887f
C326 VDD1.n142 B 0.011596f
C327 VDD1.n143 B 0.010952f
C328 VDD1.n144 B 0.020382f
C329 VDD1.n145 B 0.020382f
C330 VDD1.n146 B 0.010952f
C331 VDD1.n147 B 0.011596f
C332 VDD1.n148 B 0.025887f
C333 VDD1.n149 B 0.025887f
C334 VDD1.n150 B 0.011596f
C335 VDD1.n151 B 0.010952f
C336 VDD1.n152 B 0.020382f
C337 VDD1.n153 B 0.020382f
C338 VDD1.n154 B 0.010952f
C339 VDD1.n155 B 0.011596f
C340 VDD1.n156 B 0.025887f
C341 VDD1.n157 B 0.057743f
C342 VDD1.n158 B 0.011596f
C343 VDD1.n159 B 0.010952f
C344 VDD1.n160 B 0.044605f
C345 VDD1.n161 B 0.643031f
C346 VTAIL.n0 B 0.029291f
C347 VTAIL.n1 B 0.020162f
C348 VTAIL.n2 B 0.010834f
C349 VTAIL.n3 B 0.025608f
C350 VTAIL.n4 B 0.011471f
C351 VTAIL.n5 B 0.020162f
C352 VTAIL.n6 B 0.010834f
C353 VTAIL.n7 B 0.025608f
C354 VTAIL.n8 B 0.011471f
C355 VTAIL.n9 B 0.020162f
C356 VTAIL.n10 B 0.010834f
C357 VTAIL.n11 B 0.025608f
C358 VTAIL.n12 B 0.011471f
C359 VTAIL.n13 B 0.020162f
C360 VTAIL.n14 B 0.010834f
C361 VTAIL.n15 B 0.025608f
C362 VTAIL.n16 B 0.011471f
C363 VTAIL.n17 B 0.020162f
C364 VTAIL.n18 B 0.010834f
C365 VTAIL.n19 B 0.025608f
C366 VTAIL.n20 B 0.011471f
C367 VTAIL.n21 B 0.020162f
C368 VTAIL.n22 B 0.010834f
C369 VTAIL.n23 B 0.025608f
C370 VTAIL.n24 B 0.011471f
C371 VTAIL.n25 B 0.167889f
C372 VTAIL.t2 B 0.043566f
C373 VTAIL.n26 B 0.019206f
C374 VTAIL.n27 B 0.018103f
C375 VTAIL.n28 B 0.010834f
C376 VTAIL.n29 B 1.27809f
C377 VTAIL.n30 B 0.020162f
C378 VTAIL.n31 B 0.010834f
C379 VTAIL.n32 B 0.011471f
C380 VTAIL.n33 B 0.025608f
C381 VTAIL.n34 B 0.025608f
C382 VTAIL.n35 B 0.011471f
C383 VTAIL.n36 B 0.010834f
C384 VTAIL.n37 B 0.020162f
C385 VTAIL.n38 B 0.020162f
C386 VTAIL.n39 B 0.010834f
C387 VTAIL.n40 B 0.011471f
C388 VTAIL.n41 B 0.025608f
C389 VTAIL.n42 B 0.025608f
C390 VTAIL.n43 B 0.025608f
C391 VTAIL.n44 B 0.011471f
C392 VTAIL.n45 B 0.010834f
C393 VTAIL.n46 B 0.020162f
C394 VTAIL.n47 B 0.020162f
C395 VTAIL.n48 B 0.010834f
C396 VTAIL.n49 B 0.011153f
C397 VTAIL.n50 B 0.011153f
C398 VTAIL.n51 B 0.025608f
C399 VTAIL.n52 B 0.025608f
C400 VTAIL.n53 B 0.011471f
C401 VTAIL.n54 B 0.010834f
C402 VTAIL.n55 B 0.020162f
C403 VTAIL.n56 B 0.020162f
C404 VTAIL.n57 B 0.010834f
C405 VTAIL.n58 B 0.011471f
C406 VTAIL.n59 B 0.025608f
C407 VTAIL.n60 B 0.025608f
C408 VTAIL.n61 B 0.011471f
C409 VTAIL.n62 B 0.010834f
C410 VTAIL.n63 B 0.020162f
C411 VTAIL.n64 B 0.020162f
C412 VTAIL.n65 B 0.010834f
C413 VTAIL.n66 B 0.011471f
C414 VTAIL.n67 B 0.025608f
C415 VTAIL.n68 B 0.025608f
C416 VTAIL.n69 B 0.011471f
C417 VTAIL.n70 B 0.010834f
C418 VTAIL.n71 B 0.020162f
C419 VTAIL.n72 B 0.020162f
C420 VTAIL.n73 B 0.010834f
C421 VTAIL.n74 B 0.011471f
C422 VTAIL.n75 B 0.025608f
C423 VTAIL.n76 B 0.05712f
C424 VTAIL.n77 B 0.011471f
C425 VTAIL.n78 B 0.010834f
C426 VTAIL.n79 B 0.044124f
C427 VTAIL.n80 B 0.032056f
C428 VTAIL.n81 B 1.33153f
C429 VTAIL.n82 B 0.029291f
C430 VTAIL.n83 B 0.020162f
C431 VTAIL.n84 B 0.010834f
C432 VTAIL.n85 B 0.025608f
C433 VTAIL.n86 B 0.011471f
C434 VTAIL.n87 B 0.020162f
C435 VTAIL.n88 B 0.010834f
C436 VTAIL.n89 B 0.025608f
C437 VTAIL.n90 B 0.011471f
C438 VTAIL.n91 B 0.020162f
C439 VTAIL.n92 B 0.010834f
C440 VTAIL.n93 B 0.025608f
C441 VTAIL.n94 B 0.011471f
C442 VTAIL.n95 B 0.020162f
C443 VTAIL.n96 B 0.010834f
C444 VTAIL.n97 B 0.025608f
C445 VTAIL.n98 B 0.011471f
C446 VTAIL.n99 B 0.020162f
C447 VTAIL.n100 B 0.010834f
C448 VTAIL.n101 B 0.025608f
C449 VTAIL.n102 B 0.025608f
C450 VTAIL.n103 B 0.011471f
C451 VTAIL.n104 B 0.020162f
C452 VTAIL.n105 B 0.010834f
C453 VTAIL.n106 B 0.025608f
C454 VTAIL.n107 B 0.011471f
C455 VTAIL.n108 B 0.167889f
C456 VTAIL.t0 B 0.043566f
C457 VTAIL.n109 B 0.019206f
C458 VTAIL.n110 B 0.018103f
C459 VTAIL.n111 B 0.010834f
C460 VTAIL.n112 B 1.27809f
C461 VTAIL.n113 B 0.020162f
C462 VTAIL.n114 B 0.010834f
C463 VTAIL.n115 B 0.011471f
C464 VTAIL.n116 B 0.025608f
C465 VTAIL.n117 B 0.025608f
C466 VTAIL.n118 B 0.011471f
C467 VTAIL.n119 B 0.010834f
C468 VTAIL.n120 B 0.020162f
C469 VTAIL.n121 B 0.020162f
C470 VTAIL.n122 B 0.010834f
C471 VTAIL.n123 B 0.011471f
C472 VTAIL.n124 B 0.025608f
C473 VTAIL.n125 B 0.025608f
C474 VTAIL.n126 B 0.011471f
C475 VTAIL.n127 B 0.010834f
C476 VTAIL.n128 B 0.020162f
C477 VTAIL.n129 B 0.020162f
C478 VTAIL.n130 B 0.010834f
C479 VTAIL.n131 B 0.011153f
C480 VTAIL.n132 B 0.011153f
C481 VTAIL.n133 B 0.025608f
C482 VTAIL.n134 B 0.025608f
C483 VTAIL.n135 B 0.011471f
C484 VTAIL.n136 B 0.010834f
C485 VTAIL.n137 B 0.020162f
C486 VTAIL.n138 B 0.020162f
C487 VTAIL.n139 B 0.010834f
C488 VTAIL.n140 B 0.011471f
C489 VTAIL.n141 B 0.025608f
C490 VTAIL.n142 B 0.025608f
C491 VTAIL.n143 B 0.011471f
C492 VTAIL.n144 B 0.010834f
C493 VTAIL.n145 B 0.020162f
C494 VTAIL.n146 B 0.020162f
C495 VTAIL.n147 B 0.010834f
C496 VTAIL.n148 B 0.011471f
C497 VTAIL.n149 B 0.025608f
C498 VTAIL.n150 B 0.025608f
C499 VTAIL.n151 B 0.011471f
C500 VTAIL.n152 B 0.010834f
C501 VTAIL.n153 B 0.020162f
C502 VTAIL.n154 B 0.020162f
C503 VTAIL.n155 B 0.010834f
C504 VTAIL.n156 B 0.011471f
C505 VTAIL.n157 B 0.025608f
C506 VTAIL.n158 B 0.05712f
C507 VTAIL.n159 B 0.011471f
C508 VTAIL.n160 B 0.010834f
C509 VTAIL.n161 B 0.044124f
C510 VTAIL.n162 B 0.032056f
C511 VTAIL.n163 B 1.34679f
C512 VTAIL.n164 B 0.029291f
C513 VTAIL.n165 B 0.020162f
C514 VTAIL.n166 B 0.010834f
C515 VTAIL.n167 B 0.025608f
C516 VTAIL.n168 B 0.011471f
C517 VTAIL.n169 B 0.020162f
C518 VTAIL.n170 B 0.010834f
C519 VTAIL.n171 B 0.025608f
C520 VTAIL.n172 B 0.011471f
C521 VTAIL.n173 B 0.020162f
C522 VTAIL.n174 B 0.010834f
C523 VTAIL.n175 B 0.025608f
C524 VTAIL.n176 B 0.011471f
C525 VTAIL.n177 B 0.020162f
C526 VTAIL.n178 B 0.010834f
C527 VTAIL.n179 B 0.025608f
C528 VTAIL.n180 B 0.011471f
C529 VTAIL.n181 B 0.020162f
C530 VTAIL.n182 B 0.010834f
C531 VTAIL.n183 B 0.025608f
C532 VTAIL.n184 B 0.025608f
C533 VTAIL.n185 B 0.011471f
C534 VTAIL.n186 B 0.020162f
C535 VTAIL.n187 B 0.010834f
C536 VTAIL.n188 B 0.025608f
C537 VTAIL.n189 B 0.011471f
C538 VTAIL.n190 B 0.167889f
C539 VTAIL.t3 B 0.043566f
C540 VTAIL.n191 B 0.019206f
C541 VTAIL.n192 B 0.018103f
C542 VTAIL.n193 B 0.010834f
C543 VTAIL.n194 B 1.27809f
C544 VTAIL.n195 B 0.020162f
C545 VTAIL.n196 B 0.010834f
C546 VTAIL.n197 B 0.011471f
C547 VTAIL.n198 B 0.025608f
C548 VTAIL.n199 B 0.025608f
C549 VTAIL.n200 B 0.011471f
C550 VTAIL.n201 B 0.010834f
C551 VTAIL.n202 B 0.020162f
C552 VTAIL.n203 B 0.020162f
C553 VTAIL.n204 B 0.010834f
C554 VTAIL.n205 B 0.011471f
C555 VTAIL.n206 B 0.025608f
C556 VTAIL.n207 B 0.025608f
C557 VTAIL.n208 B 0.011471f
C558 VTAIL.n209 B 0.010834f
C559 VTAIL.n210 B 0.020162f
C560 VTAIL.n211 B 0.020162f
C561 VTAIL.n212 B 0.010834f
C562 VTAIL.n213 B 0.011153f
C563 VTAIL.n214 B 0.011153f
C564 VTAIL.n215 B 0.025608f
C565 VTAIL.n216 B 0.025608f
C566 VTAIL.n217 B 0.011471f
C567 VTAIL.n218 B 0.010834f
C568 VTAIL.n219 B 0.020162f
C569 VTAIL.n220 B 0.020162f
C570 VTAIL.n221 B 0.010834f
C571 VTAIL.n222 B 0.011471f
C572 VTAIL.n223 B 0.025608f
C573 VTAIL.n224 B 0.025608f
C574 VTAIL.n225 B 0.011471f
C575 VTAIL.n226 B 0.010834f
C576 VTAIL.n227 B 0.020162f
C577 VTAIL.n228 B 0.020162f
C578 VTAIL.n229 B 0.010834f
C579 VTAIL.n230 B 0.011471f
C580 VTAIL.n231 B 0.025608f
C581 VTAIL.n232 B 0.025608f
C582 VTAIL.n233 B 0.011471f
C583 VTAIL.n234 B 0.010834f
C584 VTAIL.n235 B 0.020162f
C585 VTAIL.n236 B 0.020162f
C586 VTAIL.n237 B 0.010834f
C587 VTAIL.n238 B 0.011471f
C588 VTAIL.n239 B 0.025608f
C589 VTAIL.n240 B 0.05712f
C590 VTAIL.n241 B 0.011471f
C591 VTAIL.n242 B 0.010834f
C592 VTAIL.n243 B 0.044124f
C593 VTAIL.n244 B 0.032056f
C594 VTAIL.n245 B 1.27062f
C595 VTAIL.n246 B 0.029291f
C596 VTAIL.n247 B 0.020162f
C597 VTAIL.n248 B 0.010834f
C598 VTAIL.n249 B 0.025608f
C599 VTAIL.n250 B 0.011471f
C600 VTAIL.n251 B 0.020162f
C601 VTAIL.n252 B 0.010834f
C602 VTAIL.n253 B 0.025608f
C603 VTAIL.n254 B 0.011471f
C604 VTAIL.n255 B 0.020162f
C605 VTAIL.n256 B 0.010834f
C606 VTAIL.n257 B 0.025608f
C607 VTAIL.n258 B 0.011471f
C608 VTAIL.n259 B 0.020162f
C609 VTAIL.n260 B 0.010834f
C610 VTAIL.n261 B 0.025608f
C611 VTAIL.n262 B 0.011471f
C612 VTAIL.n263 B 0.020162f
C613 VTAIL.n264 B 0.010834f
C614 VTAIL.n265 B 0.025608f
C615 VTAIL.n266 B 0.011471f
C616 VTAIL.n267 B 0.020162f
C617 VTAIL.n268 B 0.010834f
C618 VTAIL.n269 B 0.025608f
C619 VTAIL.n270 B 0.011471f
C620 VTAIL.n271 B 0.167889f
C621 VTAIL.t1 B 0.043566f
C622 VTAIL.n272 B 0.019206f
C623 VTAIL.n273 B 0.018103f
C624 VTAIL.n274 B 0.010834f
C625 VTAIL.n275 B 1.27809f
C626 VTAIL.n276 B 0.020162f
C627 VTAIL.n277 B 0.010834f
C628 VTAIL.n278 B 0.011471f
C629 VTAIL.n279 B 0.025608f
C630 VTAIL.n280 B 0.025608f
C631 VTAIL.n281 B 0.011471f
C632 VTAIL.n282 B 0.010834f
C633 VTAIL.n283 B 0.020162f
C634 VTAIL.n284 B 0.020162f
C635 VTAIL.n285 B 0.010834f
C636 VTAIL.n286 B 0.011471f
C637 VTAIL.n287 B 0.025608f
C638 VTAIL.n288 B 0.025608f
C639 VTAIL.n289 B 0.025608f
C640 VTAIL.n290 B 0.011471f
C641 VTAIL.n291 B 0.010834f
C642 VTAIL.n292 B 0.020162f
C643 VTAIL.n293 B 0.020162f
C644 VTAIL.n294 B 0.010834f
C645 VTAIL.n295 B 0.011153f
C646 VTAIL.n296 B 0.011153f
C647 VTAIL.n297 B 0.025608f
C648 VTAIL.n298 B 0.025608f
C649 VTAIL.n299 B 0.011471f
C650 VTAIL.n300 B 0.010834f
C651 VTAIL.n301 B 0.020162f
C652 VTAIL.n302 B 0.020162f
C653 VTAIL.n303 B 0.010834f
C654 VTAIL.n304 B 0.011471f
C655 VTAIL.n305 B 0.025608f
C656 VTAIL.n306 B 0.025608f
C657 VTAIL.n307 B 0.011471f
C658 VTAIL.n308 B 0.010834f
C659 VTAIL.n309 B 0.020162f
C660 VTAIL.n310 B 0.020162f
C661 VTAIL.n311 B 0.010834f
C662 VTAIL.n312 B 0.011471f
C663 VTAIL.n313 B 0.025608f
C664 VTAIL.n314 B 0.025608f
C665 VTAIL.n315 B 0.011471f
C666 VTAIL.n316 B 0.010834f
C667 VTAIL.n317 B 0.020162f
C668 VTAIL.n318 B 0.020162f
C669 VTAIL.n319 B 0.010834f
C670 VTAIL.n320 B 0.011471f
C671 VTAIL.n321 B 0.025608f
C672 VTAIL.n322 B 0.05712f
C673 VTAIL.n323 B 0.011471f
C674 VTAIL.n324 B 0.010834f
C675 VTAIL.n325 B 0.044124f
C676 VTAIL.n326 B 0.032056f
C677 VTAIL.n327 B 1.21728f
C678 VP.t1 B 2.61241f
C679 VP.t0 B 2.41647f
C680 VP.n0 B 5.24365f
.ends

