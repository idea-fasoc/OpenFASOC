* NGSPICE file created from diff_pair_sample_1270.ext - technology: sky130A

.subckt diff_pair_sample_1270 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t0 w_n1730_n3340# sky130_fd_pr__pfet_01v8 ad=1.9569 pd=12.19 as=1.9569 ps=12.19 w=11.86 l=0.62
X1 VDD1.t5 VP.t0 VTAIL.t2 w_n1730_n3340# sky130_fd_pr__pfet_01v8 ad=4.6254 pd=24.5 as=1.9569 ps=12.19 w=11.86 l=0.62
X2 VDD1.t4 VP.t1 VTAIL.t1 w_n1730_n3340# sky130_fd_pr__pfet_01v8 ad=1.9569 pd=12.19 as=4.6254 ps=24.5 w=11.86 l=0.62
X3 VTAIL.t3 VP.t2 VDD1.t3 w_n1730_n3340# sky130_fd_pr__pfet_01v8 ad=1.9569 pd=12.19 as=1.9569 ps=12.19 w=11.86 l=0.62
X4 VDD1.t2 VP.t3 VTAIL.t5 w_n1730_n3340# sky130_fd_pr__pfet_01v8 ad=4.6254 pd=24.5 as=1.9569 ps=12.19 w=11.86 l=0.62
X5 B.t11 B.t9 B.t10 w_n1730_n3340# sky130_fd_pr__pfet_01v8 ad=4.6254 pd=24.5 as=0 ps=0 w=11.86 l=0.62
X6 VDD2.t3 VN.t1 VTAIL.t10 w_n1730_n3340# sky130_fd_pr__pfet_01v8 ad=1.9569 pd=12.19 as=4.6254 ps=24.5 w=11.86 l=0.62
X7 VDD1.t1 VP.t4 VTAIL.t0 w_n1730_n3340# sky130_fd_pr__pfet_01v8 ad=1.9569 pd=12.19 as=4.6254 ps=24.5 w=11.86 l=0.62
X8 B.t8 B.t6 B.t7 w_n1730_n3340# sky130_fd_pr__pfet_01v8 ad=4.6254 pd=24.5 as=0 ps=0 w=11.86 l=0.62
X9 VDD2.t4 VN.t2 VTAIL.t9 w_n1730_n3340# sky130_fd_pr__pfet_01v8 ad=4.6254 pd=24.5 as=1.9569 ps=12.19 w=11.86 l=0.62
X10 VDD2.t2 VN.t3 VTAIL.t8 w_n1730_n3340# sky130_fd_pr__pfet_01v8 ad=4.6254 pd=24.5 as=1.9569 ps=12.19 w=11.86 l=0.62
X11 VTAIL.t7 VN.t4 VDD2.t1 w_n1730_n3340# sky130_fd_pr__pfet_01v8 ad=1.9569 pd=12.19 as=1.9569 ps=12.19 w=11.86 l=0.62
X12 VTAIL.t4 VP.t5 VDD1.t0 w_n1730_n3340# sky130_fd_pr__pfet_01v8 ad=1.9569 pd=12.19 as=1.9569 ps=12.19 w=11.86 l=0.62
X13 B.t5 B.t3 B.t4 w_n1730_n3340# sky130_fd_pr__pfet_01v8 ad=4.6254 pd=24.5 as=0 ps=0 w=11.86 l=0.62
X14 VDD2.t5 VN.t5 VTAIL.t6 w_n1730_n3340# sky130_fd_pr__pfet_01v8 ad=1.9569 pd=12.19 as=4.6254 ps=24.5 w=11.86 l=0.62
X15 B.t2 B.t0 B.t1 w_n1730_n3340# sky130_fd_pr__pfet_01v8 ad=4.6254 pd=24.5 as=0 ps=0 w=11.86 l=0.62
R0 VN.n0 VN.t3 551.191
R1 VN.n4 VN.t1 551.191
R2 VN.n1 VN.t4 524.37
R3 VN.n2 VN.t5 524.37
R4 VN.n5 VN.t0 524.37
R5 VN.n6 VN.t2 524.37
R6 VN.n3 VN.n2 161.3
R7 VN.n7 VN.n6 161.3
R8 VN.n2 VN.n1 48.2005
R9 VN.n6 VN.n5 48.2005
R10 VN.n7 VN.n4 45.1367
R11 VN.n3 VN.n0 45.1367
R12 VN VN.n7 41.2713
R13 VN.n5 VN.n4 13.3799
R14 VN.n1 VN.n0 13.3799
R15 VN VN.n3 0.0516364
R16 VDD2.n1 VDD2.t2 79.5337
R17 VDD2.n2 VDD2.t4 78.9751
R18 VDD2.n1 VDD2.n0 76.3835
R19 VDD2 VDD2.n3 76.3807
R20 VDD2.n2 VDD2.n1 36.6011
R21 VDD2.n3 VDD2.t0 2.74123
R22 VDD2.n3 VDD2.t3 2.74123
R23 VDD2.n0 VDD2.t1 2.74123
R24 VDD2.n0 VDD2.t5 2.74123
R25 VDD2 VDD2.n2 0.672914
R26 VTAIL.n7 VTAIL.t10 62.2963
R27 VTAIL.n11 VTAIL.t6 62.296
R28 VTAIL.n2 VTAIL.t1 62.296
R29 VTAIL.n10 VTAIL.t0 62.296
R30 VTAIL.n9 VTAIL.n8 59.5555
R31 VTAIL.n6 VTAIL.n5 59.5555
R32 VTAIL.n1 VTAIL.n0 59.5553
R33 VTAIL.n4 VTAIL.n3 59.5553
R34 VTAIL.n6 VTAIL.n4 24.2289
R35 VTAIL.n11 VTAIL.n10 23.41
R36 VTAIL.n0 VTAIL.t8 2.74123
R37 VTAIL.n0 VTAIL.t7 2.74123
R38 VTAIL.n3 VTAIL.t5 2.74123
R39 VTAIL.n3 VTAIL.t3 2.74123
R40 VTAIL.n8 VTAIL.t2 2.74123
R41 VTAIL.n8 VTAIL.t4 2.74123
R42 VTAIL.n5 VTAIL.t9 2.74123
R43 VTAIL.n5 VTAIL.t11 2.74123
R44 VTAIL.n9 VTAIL.n7 0.87981
R45 VTAIL.n2 VTAIL.n1 0.87981
R46 VTAIL.n7 VTAIL.n6 0.819465
R47 VTAIL.n10 VTAIL.n9 0.819465
R48 VTAIL.n4 VTAIL.n2 0.819465
R49 VTAIL VTAIL.n11 0.556535
R50 VTAIL VTAIL.n1 0.263431
R51 VP.n1 VP.t0 551.191
R52 VP.n6 VP.t3 524.37
R53 VP.n7 VP.t2 524.37
R54 VP.n8 VP.t1 524.37
R55 VP.n3 VP.t4 524.37
R56 VP.n2 VP.t5 524.37
R57 VP.n9 VP.n8 161.3
R58 VP.n4 VP.n3 161.3
R59 VP.n6 VP.n5 161.3
R60 VP.n7 VP.n0 80.6037
R61 VP.n7 VP.n6 48.2005
R62 VP.n8 VP.n7 48.2005
R63 VP.n3 VP.n2 48.2005
R64 VP.n4 VP.n1 45.1367
R65 VP.n5 VP.n4 40.8907
R66 VP.n2 VP.n1 13.3799
R67 VP.n5 VP.n0 0.285035
R68 VP.n9 VP.n0 0.285035
R69 VP VP.n9 0.0516364
R70 VDD1 VDD1.t5 79.6475
R71 VDD1.n1 VDD1.t2 79.5337
R72 VDD1.n1 VDD1.n0 76.3835
R73 VDD1.n3 VDD1.n2 76.2341
R74 VDD1.n3 VDD1.n1 37.5936
R75 VDD1.n2 VDD1.t0 2.74123
R76 VDD1.n2 VDD1.t1 2.74123
R77 VDD1.n0 VDD1.t3 2.74123
R78 VDD1.n0 VDD1.t4 2.74123
R79 VDD1 VDD1.n3 0.147052
R80 B.n102 B.t9 665.086
R81 B.n110 B.t0 665.086
R82 B.n32 B.t6 665.086
R83 B.n40 B.t3 665.086
R84 B.n367 B.n366 585
R85 B.n368 B.n61 585
R86 B.n370 B.n369 585
R87 B.n371 B.n60 585
R88 B.n373 B.n372 585
R89 B.n374 B.n59 585
R90 B.n376 B.n375 585
R91 B.n377 B.n58 585
R92 B.n379 B.n378 585
R93 B.n380 B.n57 585
R94 B.n382 B.n381 585
R95 B.n383 B.n56 585
R96 B.n385 B.n384 585
R97 B.n386 B.n55 585
R98 B.n388 B.n387 585
R99 B.n389 B.n54 585
R100 B.n391 B.n390 585
R101 B.n392 B.n53 585
R102 B.n394 B.n393 585
R103 B.n395 B.n52 585
R104 B.n397 B.n396 585
R105 B.n398 B.n51 585
R106 B.n400 B.n399 585
R107 B.n401 B.n50 585
R108 B.n403 B.n402 585
R109 B.n404 B.n49 585
R110 B.n406 B.n405 585
R111 B.n407 B.n48 585
R112 B.n409 B.n408 585
R113 B.n410 B.n47 585
R114 B.n412 B.n411 585
R115 B.n413 B.n46 585
R116 B.n415 B.n414 585
R117 B.n416 B.n45 585
R118 B.n418 B.n417 585
R119 B.n419 B.n44 585
R120 B.n421 B.n420 585
R121 B.n422 B.n43 585
R122 B.n424 B.n423 585
R123 B.n425 B.n42 585
R124 B.n427 B.n426 585
R125 B.n429 B.n39 585
R126 B.n431 B.n430 585
R127 B.n432 B.n38 585
R128 B.n434 B.n433 585
R129 B.n435 B.n37 585
R130 B.n437 B.n436 585
R131 B.n438 B.n36 585
R132 B.n440 B.n439 585
R133 B.n441 B.n35 585
R134 B.n443 B.n442 585
R135 B.n445 B.n444 585
R136 B.n446 B.n31 585
R137 B.n448 B.n447 585
R138 B.n449 B.n30 585
R139 B.n451 B.n450 585
R140 B.n452 B.n29 585
R141 B.n454 B.n453 585
R142 B.n455 B.n28 585
R143 B.n457 B.n456 585
R144 B.n458 B.n27 585
R145 B.n460 B.n459 585
R146 B.n461 B.n26 585
R147 B.n463 B.n462 585
R148 B.n464 B.n25 585
R149 B.n466 B.n465 585
R150 B.n467 B.n24 585
R151 B.n469 B.n468 585
R152 B.n470 B.n23 585
R153 B.n472 B.n471 585
R154 B.n473 B.n22 585
R155 B.n475 B.n474 585
R156 B.n476 B.n21 585
R157 B.n478 B.n477 585
R158 B.n479 B.n20 585
R159 B.n481 B.n480 585
R160 B.n482 B.n19 585
R161 B.n484 B.n483 585
R162 B.n485 B.n18 585
R163 B.n487 B.n486 585
R164 B.n488 B.n17 585
R165 B.n490 B.n489 585
R166 B.n491 B.n16 585
R167 B.n493 B.n492 585
R168 B.n494 B.n15 585
R169 B.n496 B.n495 585
R170 B.n497 B.n14 585
R171 B.n499 B.n498 585
R172 B.n500 B.n13 585
R173 B.n502 B.n501 585
R174 B.n503 B.n12 585
R175 B.n505 B.n504 585
R176 B.n365 B.n62 585
R177 B.n364 B.n363 585
R178 B.n362 B.n63 585
R179 B.n361 B.n360 585
R180 B.n359 B.n64 585
R181 B.n358 B.n357 585
R182 B.n356 B.n65 585
R183 B.n355 B.n354 585
R184 B.n353 B.n66 585
R185 B.n352 B.n351 585
R186 B.n350 B.n67 585
R187 B.n349 B.n348 585
R188 B.n347 B.n68 585
R189 B.n346 B.n345 585
R190 B.n344 B.n69 585
R191 B.n343 B.n342 585
R192 B.n341 B.n70 585
R193 B.n340 B.n339 585
R194 B.n338 B.n71 585
R195 B.n337 B.n336 585
R196 B.n335 B.n72 585
R197 B.n334 B.n333 585
R198 B.n332 B.n73 585
R199 B.n331 B.n330 585
R200 B.n329 B.n74 585
R201 B.n328 B.n327 585
R202 B.n326 B.n75 585
R203 B.n325 B.n324 585
R204 B.n323 B.n76 585
R205 B.n322 B.n321 585
R206 B.n320 B.n77 585
R207 B.n319 B.n318 585
R208 B.n317 B.n78 585
R209 B.n316 B.n315 585
R210 B.n314 B.n79 585
R211 B.n313 B.n312 585
R212 B.n311 B.n80 585
R213 B.n310 B.n309 585
R214 B.n308 B.n81 585
R215 B.n169 B.n168 585
R216 B.n170 B.n131 585
R217 B.n172 B.n171 585
R218 B.n173 B.n130 585
R219 B.n175 B.n174 585
R220 B.n176 B.n129 585
R221 B.n178 B.n177 585
R222 B.n179 B.n128 585
R223 B.n181 B.n180 585
R224 B.n182 B.n127 585
R225 B.n184 B.n183 585
R226 B.n185 B.n126 585
R227 B.n187 B.n186 585
R228 B.n188 B.n125 585
R229 B.n190 B.n189 585
R230 B.n191 B.n124 585
R231 B.n193 B.n192 585
R232 B.n194 B.n123 585
R233 B.n196 B.n195 585
R234 B.n197 B.n122 585
R235 B.n199 B.n198 585
R236 B.n200 B.n121 585
R237 B.n202 B.n201 585
R238 B.n203 B.n120 585
R239 B.n205 B.n204 585
R240 B.n206 B.n119 585
R241 B.n208 B.n207 585
R242 B.n209 B.n118 585
R243 B.n211 B.n210 585
R244 B.n212 B.n117 585
R245 B.n214 B.n213 585
R246 B.n215 B.n116 585
R247 B.n217 B.n216 585
R248 B.n218 B.n115 585
R249 B.n220 B.n219 585
R250 B.n221 B.n114 585
R251 B.n223 B.n222 585
R252 B.n224 B.n113 585
R253 B.n226 B.n225 585
R254 B.n227 B.n112 585
R255 B.n229 B.n228 585
R256 B.n231 B.n109 585
R257 B.n233 B.n232 585
R258 B.n234 B.n108 585
R259 B.n236 B.n235 585
R260 B.n237 B.n107 585
R261 B.n239 B.n238 585
R262 B.n240 B.n106 585
R263 B.n242 B.n241 585
R264 B.n243 B.n105 585
R265 B.n245 B.n244 585
R266 B.n247 B.n246 585
R267 B.n248 B.n101 585
R268 B.n250 B.n249 585
R269 B.n251 B.n100 585
R270 B.n253 B.n252 585
R271 B.n254 B.n99 585
R272 B.n256 B.n255 585
R273 B.n257 B.n98 585
R274 B.n259 B.n258 585
R275 B.n260 B.n97 585
R276 B.n262 B.n261 585
R277 B.n263 B.n96 585
R278 B.n265 B.n264 585
R279 B.n266 B.n95 585
R280 B.n268 B.n267 585
R281 B.n269 B.n94 585
R282 B.n271 B.n270 585
R283 B.n272 B.n93 585
R284 B.n274 B.n273 585
R285 B.n275 B.n92 585
R286 B.n277 B.n276 585
R287 B.n278 B.n91 585
R288 B.n280 B.n279 585
R289 B.n281 B.n90 585
R290 B.n283 B.n282 585
R291 B.n284 B.n89 585
R292 B.n286 B.n285 585
R293 B.n287 B.n88 585
R294 B.n289 B.n288 585
R295 B.n290 B.n87 585
R296 B.n292 B.n291 585
R297 B.n293 B.n86 585
R298 B.n295 B.n294 585
R299 B.n296 B.n85 585
R300 B.n298 B.n297 585
R301 B.n299 B.n84 585
R302 B.n301 B.n300 585
R303 B.n302 B.n83 585
R304 B.n304 B.n303 585
R305 B.n305 B.n82 585
R306 B.n307 B.n306 585
R307 B.n167 B.n132 585
R308 B.n166 B.n165 585
R309 B.n164 B.n133 585
R310 B.n163 B.n162 585
R311 B.n161 B.n134 585
R312 B.n160 B.n159 585
R313 B.n158 B.n135 585
R314 B.n157 B.n156 585
R315 B.n155 B.n136 585
R316 B.n154 B.n153 585
R317 B.n152 B.n137 585
R318 B.n151 B.n150 585
R319 B.n149 B.n138 585
R320 B.n148 B.n147 585
R321 B.n146 B.n139 585
R322 B.n145 B.n144 585
R323 B.n143 B.n140 585
R324 B.n142 B.n141 585
R325 B.n2 B.n0 585
R326 B.n533 B.n1 585
R327 B.n532 B.n531 585
R328 B.n530 B.n3 585
R329 B.n529 B.n528 585
R330 B.n527 B.n4 585
R331 B.n526 B.n525 585
R332 B.n524 B.n5 585
R333 B.n523 B.n522 585
R334 B.n521 B.n6 585
R335 B.n520 B.n519 585
R336 B.n518 B.n7 585
R337 B.n517 B.n516 585
R338 B.n515 B.n8 585
R339 B.n514 B.n513 585
R340 B.n512 B.n9 585
R341 B.n511 B.n510 585
R342 B.n509 B.n10 585
R343 B.n508 B.n507 585
R344 B.n506 B.n11 585
R345 B.n535 B.n534 585
R346 B.n168 B.n167 545.355
R347 B.n504 B.n11 545.355
R348 B.n306 B.n81 545.355
R349 B.n366 B.n365 545.355
R350 B.n167 B.n166 163.367
R351 B.n166 B.n133 163.367
R352 B.n162 B.n133 163.367
R353 B.n162 B.n161 163.367
R354 B.n161 B.n160 163.367
R355 B.n160 B.n135 163.367
R356 B.n156 B.n135 163.367
R357 B.n156 B.n155 163.367
R358 B.n155 B.n154 163.367
R359 B.n154 B.n137 163.367
R360 B.n150 B.n137 163.367
R361 B.n150 B.n149 163.367
R362 B.n149 B.n148 163.367
R363 B.n148 B.n139 163.367
R364 B.n144 B.n139 163.367
R365 B.n144 B.n143 163.367
R366 B.n143 B.n142 163.367
R367 B.n142 B.n2 163.367
R368 B.n534 B.n2 163.367
R369 B.n534 B.n533 163.367
R370 B.n533 B.n532 163.367
R371 B.n532 B.n3 163.367
R372 B.n528 B.n3 163.367
R373 B.n528 B.n527 163.367
R374 B.n527 B.n526 163.367
R375 B.n526 B.n5 163.367
R376 B.n522 B.n5 163.367
R377 B.n522 B.n521 163.367
R378 B.n521 B.n520 163.367
R379 B.n520 B.n7 163.367
R380 B.n516 B.n7 163.367
R381 B.n516 B.n515 163.367
R382 B.n515 B.n514 163.367
R383 B.n514 B.n9 163.367
R384 B.n510 B.n9 163.367
R385 B.n510 B.n509 163.367
R386 B.n509 B.n508 163.367
R387 B.n508 B.n11 163.367
R388 B.n168 B.n131 163.367
R389 B.n172 B.n131 163.367
R390 B.n173 B.n172 163.367
R391 B.n174 B.n173 163.367
R392 B.n174 B.n129 163.367
R393 B.n178 B.n129 163.367
R394 B.n179 B.n178 163.367
R395 B.n180 B.n179 163.367
R396 B.n180 B.n127 163.367
R397 B.n184 B.n127 163.367
R398 B.n185 B.n184 163.367
R399 B.n186 B.n185 163.367
R400 B.n186 B.n125 163.367
R401 B.n190 B.n125 163.367
R402 B.n191 B.n190 163.367
R403 B.n192 B.n191 163.367
R404 B.n192 B.n123 163.367
R405 B.n196 B.n123 163.367
R406 B.n197 B.n196 163.367
R407 B.n198 B.n197 163.367
R408 B.n198 B.n121 163.367
R409 B.n202 B.n121 163.367
R410 B.n203 B.n202 163.367
R411 B.n204 B.n203 163.367
R412 B.n204 B.n119 163.367
R413 B.n208 B.n119 163.367
R414 B.n209 B.n208 163.367
R415 B.n210 B.n209 163.367
R416 B.n210 B.n117 163.367
R417 B.n214 B.n117 163.367
R418 B.n215 B.n214 163.367
R419 B.n216 B.n215 163.367
R420 B.n216 B.n115 163.367
R421 B.n220 B.n115 163.367
R422 B.n221 B.n220 163.367
R423 B.n222 B.n221 163.367
R424 B.n222 B.n113 163.367
R425 B.n226 B.n113 163.367
R426 B.n227 B.n226 163.367
R427 B.n228 B.n227 163.367
R428 B.n228 B.n109 163.367
R429 B.n233 B.n109 163.367
R430 B.n234 B.n233 163.367
R431 B.n235 B.n234 163.367
R432 B.n235 B.n107 163.367
R433 B.n239 B.n107 163.367
R434 B.n240 B.n239 163.367
R435 B.n241 B.n240 163.367
R436 B.n241 B.n105 163.367
R437 B.n245 B.n105 163.367
R438 B.n246 B.n245 163.367
R439 B.n246 B.n101 163.367
R440 B.n250 B.n101 163.367
R441 B.n251 B.n250 163.367
R442 B.n252 B.n251 163.367
R443 B.n252 B.n99 163.367
R444 B.n256 B.n99 163.367
R445 B.n257 B.n256 163.367
R446 B.n258 B.n257 163.367
R447 B.n258 B.n97 163.367
R448 B.n262 B.n97 163.367
R449 B.n263 B.n262 163.367
R450 B.n264 B.n263 163.367
R451 B.n264 B.n95 163.367
R452 B.n268 B.n95 163.367
R453 B.n269 B.n268 163.367
R454 B.n270 B.n269 163.367
R455 B.n270 B.n93 163.367
R456 B.n274 B.n93 163.367
R457 B.n275 B.n274 163.367
R458 B.n276 B.n275 163.367
R459 B.n276 B.n91 163.367
R460 B.n280 B.n91 163.367
R461 B.n281 B.n280 163.367
R462 B.n282 B.n281 163.367
R463 B.n282 B.n89 163.367
R464 B.n286 B.n89 163.367
R465 B.n287 B.n286 163.367
R466 B.n288 B.n287 163.367
R467 B.n288 B.n87 163.367
R468 B.n292 B.n87 163.367
R469 B.n293 B.n292 163.367
R470 B.n294 B.n293 163.367
R471 B.n294 B.n85 163.367
R472 B.n298 B.n85 163.367
R473 B.n299 B.n298 163.367
R474 B.n300 B.n299 163.367
R475 B.n300 B.n83 163.367
R476 B.n304 B.n83 163.367
R477 B.n305 B.n304 163.367
R478 B.n306 B.n305 163.367
R479 B.n310 B.n81 163.367
R480 B.n311 B.n310 163.367
R481 B.n312 B.n311 163.367
R482 B.n312 B.n79 163.367
R483 B.n316 B.n79 163.367
R484 B.n317 B.n316 163.367
R485 B.n318 B.n317 163.367
R486 B.n318 B.n77 163.367
R487 B.n322 B.n77 163.367
R488 B.n323 B.n322 163.367
R489 B.n324 B.n323 163.367
R490 B.n324 B.n75 163.367
R491 B.n328 B.n75 163.367
R492 B.n329 B.n328 163.367
R493 B.n330 B.n329 163.367
R494 B.n330 B.n73 163.367
R495 B.n334 B.n73 163.367
R496 B.n335 B.n334 163.367
R497 B.n336 B.n335 163.367
R498 B.n336 B.n71 163.367
R499 B.n340 B.n71 163.367
R500 B.n341 B.n340 163.367
R501 B.n342 B.n341 163.367
R502 B.n342 B.n69 163.367
R503 B.n346 B.n69 163.367
R504 B.n347 B.n346 163.367
R505 B.n348 B.n347 163.367
R506 B.n348 B.n67 163.367
R507 B.n352 B.n67 163.367
R508 B.n353 B.n352 163.367
R509 B.n354 B.n353 163.367
R510 B.n354 B.n65 163.367
R511 B.n358 B.n65 163.367
R512 B.n359 B.n358 163.367
R513 B.n360 B.n359 163.367
R514 B.n360 B.n63 163.367
R515 B.n364 B.n63 163.367
R516 B.n365 B.n364 163.367
R517 B.n504 B.n503 163.367
R518 B.n503 B.n502 163.367
R519 B.n502 B.n13 163.367
R520 B.n498 B.n13 163.367
R521 B.n498 B.n497 163.367
R522 B.n497 B.n496 163.367
R523 B.n496 B.n15 163.367
R524 B.n492 B.n15 163.367
R525 B.n492 B.n491 163.367
R526 B.n491 B.n490 163.367
R527 B.n490 B.n17 163.367
R528 B.n486 B.n17 163.367
R529 B.n486 B.n485 163.367
R530 B.n485 B.n484 163.367
R531 B.n484 B.n19 163.367
R532 B.n480 B.n19 163.367
R533 B.n480 B.n479 163.367
R534 B.n479 B.n478 163.367
R535 B.n478 B.n21 163.367
R536 B.n474 B.n21 163.367
R537 B.n474 B.n473 163.367
R538 B.n473 B.n472 163.367
R539 B.n472 B.n23 163.367
R540 B.n468 B.n23 163.367
R541 B.n468 B.n467 163.367
R542 B.n467 B.n466 163.367
R543 B.n466 B.n25 163.367
R544 B.n462 B.n25 163.367
R545 B.n462 B.n461 163.367
R546 B.n461 B.n460 163.367
R547 B.n460 B.n27 163.367
R548 B.n456 B.n27 163.367
R549 B.n456 B.n455 163.367
R550 B.n455 B.n454 163.367
R551 B.n454 B.n29 163.367
R552 B.n450 B.n29 163.367
R553 B.n450 B.n449 163.367
R554 B.n449 B.n448 163.367
R555 B.n448 B.n31 163.367
R556 B.n444 B.n31 163.367
R557 B.n444 B.n443 163.367
R558 B.n443 B.n35 163.367
R559 B.n439 B.n35 163.367
R560 B.n439 B.n438 163.367
R561 B.n438 B.n437 163.367
R562 B.n437 B.n37 163.367
R563 B.n433 B.n37 163.367
R564 B.n433 B.n432 163.367
R565 B.n432 B.n431 163.367
R566 B.n431 B.n39 163.367
R567 B.n426 B.n39 163.367
R568 B.n426 B.n425 163.367
R569 B.n425 B.n424 163.367
R570 B.n424 B.n43 163.367
R571 B.n420 B.n43 163.367
R572 B.n420 B.n419 163.367
R573 B.n419 B.n418 163.367
R574 B.n418 B.n45 163.367
R575 B.n414 B.n45 163.367
R576 B.n414 B.n413 163.367
R577 B.n413 B.n412 163.367
R578 B.n412 B.n47 163.367
R579 B.n408 B.n47 163.367
R580 B.n408 B.n407 163.367
R581 B.n407 B.n406 163.367
R582 B.n406 B.n49 163.367
R583 B.n402 B.n49 163.367
R584 B.n402 B.n401 163.367
R585 B.n401 B.n400 163.367
R586 B.n400 B.n51 163.367
R587 B.n396 B.n51 163.367
R588 B.n396 B.n395 163.367
R589 B.n395 B.n394 163.367
R590 B.n394 B.n53 163.367
R591 B.n390 B.n53 163.367
R592 B.n390 B.n389 163.367
R593 B.n389 B.n388 163.367
R594 B.n388 B.n55 163.367
R595 B.n384 B.n55 163.367
R596 B.n384 B.n383 163.367
R597 B.n383 B.n382 163.367
R598 B.n382 B.n57 163.367
R599 B.n378 B.n57 163.367
R600 B.n378 B.n377 163.367
R601 B.n377 B.n376 163.367
R602 B.n376 B.n59 163.367
R603 B.n372 B.n59 163.367
R604 B.n372 B.n371 163.367
R605 B.n371 B.n370 163.367
R606 B.n370 B.n61 163.367
R607 B.n366 B.n61 163.367
R608 B.n102 B.t11 131.381
R609 B.n40 B.t4 131.381
R610 B.n110 B.t2 131.367
R611 B.n32 B.t7 131.367
R612 B.n103 B.t10 112.957
R613 B.n41 B.t5 112.957
R614 B.n111 B.t1 112.942
R615 B.n33 B.t8 112.942
R616 B.n104 B.n103 59.5399
R617 B.n230 B.n111 59.5399
R618 B.n34 B.n33 59.5399
R619 B.n428 B.n41 59.5399
R620 B.n506 B.n505 35.4346
R621 B.n367 B.n62 35.4346
R622 B.n308 B.n307 35.4346
R623 B.n169 B.n132 35.4346
R624 B.n103 B.n102 18.4247
R625 B.n111 B.n110 18.4247
R626 B.n33 B.n32 18.4247
R627 B.n41 B.n40 18.4247
R628 B B.n535 18.0485
R629 B.n505 B.n12 10.6151
R630 B.n501 B.n12 10.6151
R631 B.n501 B.n500 10.6151
R632 B.n500 B.n499 10.6151
R633 B.n499 B.n14 10.6151
R634 B.n495 B.n14 10.6151
R635 B.n495 B.n494 10.6151
R636 B.n494 B.n493 10.6151
R637 B.n493 B.n16 10.6151
R638 B.n489 B.n16 10.6151
R639 B.n489 B.n488 10.6151
R640 B.n488 B.n487 10.6151
R641 B.n487 B.n18 10.6151
R642 B.n483 B.n18 10.6151
R643 B.n483 B.n482 10.6151
R644 B.n482 B.n481 10.6151
R645 B.n481 B.n20 10.6151
R646 B.n477 B.n20 10.6151
R647 B.n477 B.n476 10.6151
R648 B.n476 B.n475 10.6151
R649 B.n475 B.n22 10.6151
R650 B.n471 B.n22 10.6151
R651 B.n471 B.n470 10.6151
R652 B.n470 B.n469 10.6151
R653 B.n469 B.n24 10.6151
R654 B.n465 B.n24 10.6151
R655 B.n465 B.n464 10.6151
R656 B.n464 B.n463 10.6151
R657 B.n463 B.n26 10.6151
R658 B.n459 B.n26 10.6151
R659 B.n459 B.n458 10.6151
R660 B.n458 B.n457 10.6151
R661 B.n457 B.n28 10.6151
R662 B.n453 B.n28 10.6151
R663 B.n453 B.n452 10.6151
R664 B.n452 B.n451 10.6151
R665 B.n451 B.n30 10.6151
R666 B.n447 B.n30 10.6151
R667 B.n447 B.n446 10.6151
R668 B.n446 B.n445 10.6151
R669 B.n442 B.n441 10.6151
R670 B.n441 B.n440 10.6151
R671 B.n440 B.n36 10.6151
R672 B.n436 B.n36 10.6151
R673 B.n436 B.n435 10.6151
R674 B.n435 B.n434 10.6151
R675 B.n434 B.n38 10.6151
R676 B.n430 B.n38 10.6151
R677 B.n430 B.n429 10.6151
R678 B.n427 B.n42 10.6151
R679 B.n423 B.n42 10.6151
R680 B.n423 B.n422 10.6151
R681 B.n422 B.n421 10.6151
R682 B.n421 B.n44 10.6151
R683 B.n417 B.n44 10.6151
R684 B.n417 B.n416 10.6151
R685 B.n416 B.n415 10.6151
R686 B.n415 B.n46 10.6151
R687 B.n411 B.n46 10.6151
R688 B.n411 B.n410 10.6151
R689 B.n410 B.n409 10.6151
R690 B.n409 B.n48 10.6151
R691 B.n405 B.n48 10.6151
R692 B.n405 B.n404 10.6151
R693 B.n404 B.n403 10.6151
R694 B.n403 B.n50 10.6151
R695 B.n399 B.n50 10.6151
R696 B.n399 B.n398 10.6151
R697 B.n398 B.n397 10.6151
R698 B.n397 B.n52 10.6151
R699 B.n393 B.n52 10.6151
R700 B.n393 B.n392 10.6151
R701 B.n392 B.n391 10.6151
R702 B.n391 B.n54 10.6151
R703 B.n387 B.n54 10.6151
R704 B.n387 B.n386 10.6151
R705 B.n386 B.n385 10.6151
R706 B.n385 B.n56 10.6151
R707 B.n381 B.n56 10.6151
R708 B.n381 B.n380 10.6151
R709 B.n380 B.n379 10.6151
R710 B.n379 B.n58 10.6151
R711 B.n375 B.n58 10.6151
R712 B.n375 B.n374 10.6151
R713 B.n374 B.n373 10.6151
R714 B.n373 B.n60 10.6151
R715 B.n369 B.n60 10.6151
R716 B.n369 B.n368 10.6151
R717 B.n368 B.n367 10.6151
R718 B.n309 B.n308 10.6151
R719 B.n309 B.n80 10.6151
R720 B.n313 B.n80 10.6151
R721 B.n314 B.n313 10.6151
R722 B.n315 B.n314 10.6151
R723 B.n315 B.n78 10.6151
R724 B.n319 B.n78 10.6151
R725 B.n320 B.n319 10.6151
R726 B.n321 B.n320 10.6151
R727 B.n321 B.n76 10.6151
R728 B.n325 B.n76 10.6151
R729 B.n326 B.n325 10.6151
R730 B.n327 B.n326 10.6151
R731 B.n327 B.n74 10.6151
R732 B.n331 B.n74 10.6151
R733 B.n332 B.n331 10.6151
R734 B.n333 B.n332 10.6151
R735 B.n333 B.n72 10.6151
R736 B.n337 B.n72 10.6151
R737 B.n338 B.n337 10.6151
R738 B.n339 B.n338 10.6151
R739 B.n339 B.n70 10.6151
R740 B.n343 B.n70 10.6151
R741 B.n344 B.n343 10.6151
R742 B.n345 B.n344 10.6151
R743 B.n345 B.n68 10.6151
R744 B.n349 B.n68 10.6151
R745 B.n350 B.n349 10.6151
R746 B.n351 B.n350 10.6151
R747 B.n351 B.n66 10.6151
R748 B.n355 B.n66 10.6151
R749 B.n356 B.n355 10.6151
R750 B.n357 B.n356 10.6151
R751 B.n357 B.n64 10.6151
R752 B.n361 B.n64 10.6151
R753 B.n362 B.n361 10.6151
R754 B.n363 B.n362 10.6151
R755 B.n363 B.n62 10.6151
R756 B.n170 B.n169 10.6151
R757 B.n171 B.n170 10.6151
R758 B.n171 B.n130 10.6151
R759 B.n175 B.n130 10.6151
R760 B.n176 B.n175 10.6151
R761 B.n177 B.n176 10.6151
R762 B.n177 B.n128 10.6151
R763 B.n181 B.n128 10.6151
R764 B.n182 B.n181 10.6151
R765 B.n183 B.n182 10.6151
R766 B.n183 B.n126 10.6151
R767 B.n187 B.n126 10.6151
R768 B.n188 B.n187 10.6151
R769 B.n189 B.n188 10.6151
R770 B.n189 B.n124 10.6151
R771 B.n193 B.n124 10.6151
R772 B.n194 B.n193 10.6151
R773 B.n195 B.n194 10.6151
R774 B.n195 B.n122 10.6151
R775 B.n199 B.n122 10.6151
R776 B.n200 B.n199 10.6151
R777 B.n201 B.n200 10.6151
R778 B.n201 B.n120 10.6151
R779 B.n205 B.n120 10.6151
R780 B.n206 B.n205 10.6151
R781 B.n207 B.n206 10.6151
R782 B.n207 B.n118 10.6151
R783 B.n211 B.n118 10.6151
R784 B.n212 B.n211 10.6151
R785 B.n213 B.n212 10.6151
R786 B.n213 B.n116 10.6151
R787 B.n217 B.n116 10.6151
R788 B.n218 B.n217 10.6151
R789 B.n219 B.n218 10.6151
R790 B.n219 B.n114 10.6151
R791 B.n223 B.n114 10.6151
R792 B.n224 B.n223 10.6151
R793 B.n225 B.n224 10.6151
R794 B.n225 B.n112 10.6151
R795 B.n229 B.n112 10.6151
R796 B.n232 B.n231 10.6151
R797 B.n232 B.n108 10.6151
R798 B.n236 B.n108 10.6151
R799 B.n237 B.n236 10.6151
R800 B.n238 B.n237 10.6151
R801 B.n238 B.n106 10.6151
R802 B.n242 B.n106 10.6151
R803 B.n243 B.n242 10.6151
R804 B.n244 B.n243 10.6151
R805 B.n248 B.n247 10.6151
R806 B.n249 B.n248 10.6151
R807 B.n249 B.n100 10.6151
R808 B.n253 B.n100 10.6151
R809 B.n254 B.n253 10.6151
R810 B.n255 B.n254 10.6151
R811 B.n255 B.n98 10.6151
R812 B.n259 B.n98 10.6151
R813 B.n260 B.n259 10.6151
R814 B.n261 B.n260 10.6151
R815 B.n261 B.n96 10.6151
R816 B.n265 B.n96 10.6151
R817 B.n266 B.n265 10.6151
R818 B.n267 B.n266 10.6151
R819 B.n267 B.n94 10.6151
R820 B.n271 B.n94 10.6151
R821 B.n272 B.n271 10.6151
R822 B.n273 B.n272 10.6151
R823 B.n273 B.n92 10.6151
R824 B.n277 B.n92 10.6151
R825 B.n278 B.n277 10.6151
R826 B.n279 B.n278 10.6151
R827 B.n279 B.n90 10.6151
R828 B.n283 B.n90 10.6151
R829 B.n284 B.n283 10.6151
R830 B.n285 B.n284 10.6151
R831 B.n285 B.n88 10.6151
R832 B.n289 B.n88 10.6151
R833 B.n290 B.n289 10.6151
R834 B.n291 B.n290 10.6151
R835 B.n291 B.n86 10.6151
R836 B.n295 B.n86 10.6151
R837 B.n296 B.n295 10.6151
R838 B.n297 B.n296 10.6151
R839 B.n297 B.n84 10.6151
R840 B.n301 B.n84 10.6151
R841 B.n302 B.n301 10.6151
R842 B.n303 B.n302 10.6151
R843 B.n303 B.n82 10.6151
R844 B.n307 B.n82 10.6151
R845 B.n165 B.n132 10.6151
R846 B.n165 B.n164 10.6151
R847 B.n164 B.n163 10.6151
R848 B.n163 B.n134 10.6151
R849 B.n159 B.n134 10.6151
R850 B.n159 B.n158 10.6151
R851 B.n158 B.n157 10.6151
R852 B.n157 B.n136 10.6151
R853 B.n153 B.n136 10.6151
R854 B.n153 B.n152 10.6151
R855 B.n152 B.n151 10.6151
R856 B.n151 B.n138 10.6151
R857 B.n147 B.n138 10.6151
R858 B.n147 B.n146 10.6151
R859 B.n146 B.n145 10.6151
R860 B.n145 B.n140 10.6151
R861 B.n141 B.n140 10.6151
R862 B.n141 B.n0 10.6151
R863 B.n531 B.n1 10.6151
R864 B.n531 B.n530 10.6151
R865 B.n530 B.n529 10.6151
R866 B.n529 B.n4 10.6151
R867 B.n525 B.n4 10.6151
R868 B.n525 B.n524 10.6151
R869 B.n524 B.n523 10.6151
R870 B.n523 B.n6 10.6151
R871 B.n519 B.n6 10.6151
R872 B.n519 B.n518 10.6151
R873 B.n518 B.n517 10.6151
R874 B.n517 B.n8 10.6151
R875 B.n513 B.n8 10.6151
R876 B.n513 B.n512 10.6151
R877 B.n512 B.n511 10.6151
R878 B.n511 B.n10 10.6151
R879 B.n507 B.n10 10.6151
R880 B.n507 B.n506 10.6151
R881 B.n445 B.n34 9.36635
R882 B.n428 B.n427 9.36635
R883 B.n230 B.n229 9.36635
R884 B.n247 B.n104 9.36635
R885 B.n535 B.n0 2.81026
R886 B.n535 B.n1 2.81026
R887 B.n442 B.n34 1.24928
R888 B.n429 B.n428 1.24928
R889 B.n231 B.n230 1.24928
R890 B.n244 B.n104 1.24928
C0 VDD1 VN 0.148421f
C1 VN VP 4.97131f
C2 VDD1 VDD2 0.682489f
C3 VP VDD2 0.291251f
C4 VDD1 B 1.52466f
C5 VDD1 w_n1730_n3340# 1.77961f
C6 VP B 1.10171f
C7 w_n1730_n3340# VP 3.00088f
C8 VDD1 VTAIL 10.3005f
C9 VTAIL VP 3.71536f
C10 VN VDD2 4.03372f
C11 VN B 0.747457f
C12 w_n1730_n3340# VN 2.78273f
C13 VDD2 B 1.55175f
C14 w_n1730_n3340# VDD2 1.80118f
C15 VTAIL VN 3.70073f
C16 w_n1730_n3340# B 6.90407f
C17 VTAIL VDD2 10.333799f
C18 VTAIL B 2.62943f
C19 w_n1730_n3340# VTAIL 2.92579f
C20 VDD1 VP 4.17196f
C21 VDD2 VSUBS 1.296957f
C22 VDD1 VSUBS 1.591414f
C23 VTAIL VSUBS 0.723231f
C24 VN VSUBS 4.41918f
C25 VP VSUBS 1.410725f
C26 B VSUBS 2.66262f
C27 w_n1730_n3340# VSUBS 71.1445f
C28 B.n0 VSUBS 0.004681f
C29 B.n1 VSUBS 0.004681f
C30 B.n2 VSUBS 0.007403f
C31 B.n3 VSUBS 0.007403f
C32 B.n4 VSUBS 0.007403f
C33 B.n5 VSUBS 0.007403f
C34 B.n6 VSUBS 0.007403f
C35 B.n7 VSUBS 0.007403f
C36 B.n8 VSUBS 0.007403f
C37 B.n9 VSUBS 0.007403f
C38 B.n10 VSUBS 0.007403f
C39 B.n11 VSUBS 0.017709f
C40 B.n12 VSUBS 0.007403f
C41 B.n13 VSUBS 0.007403f
C42 B.n14 VSUBS 0.007403f
C43 B.n15 VSUBS 0.007403f
C44 B.n16 VSUBS 0.007403f
C45 B.n17 VSUBS 0.007403f
C46 B.n18 VSUBS 0.007403f
C47 B.n19 VSUBS 0.007403f
C48 B.n20 VSUBS 0.007403f
C49 B.n21 VSUBS 0.007403f
C50 B.n22 VSUBS 0.007403f
C51 B.n23 VSUBS 0.007403f
C52 B.n24 VSUBS 0.007403f
C53 B.n25 VSUBS 0.007403f
C54 B.n26 VSUBS 0.007403f
C55 B.n27 VSUBS 0.007403f
C56 B.n28 VSUBS 0.007403f
C57 B.n29 VSUBS 0.007403f
C58 B.n30 VSUBS 0.007403f
C59 B.n31 VSUBS 0.007403f
C60 B.t8 VSUBS 0.408215f
C61 B.t7 VSUBS 0.416165f
C62 B.t6 VSUBS 0.318363f
C63 B.n32 VSUBS 0.134956f
C64 B.n33 VSUBS 0.06724f
C65 B.n34 VSUBS 0.017151f
C66 B.n35 VSUBS 0.007403f
C67 B.n36 VSUBS 0.007403f
C68 B.n37 VSUBS 0.007403f
C69 B.n38 VSUBS 0.007403f
C70 B.n39 VSUBS 0.007403f
C71 B.t5 VSUBS 0.408208f
C72 B.t4 VSUBS 0.416158f
C73 B.t3 VSUBS 0.318363f
C74 B.n40 VSUBS 0.134963f
C75 B.n41 VSUBS 0.067248f
C76 B.n42 VSUBS 0.007403f
C77 B.n43 VSUBS 0.007403f
C78 B.n44 VSUBS 0.007403f
C79 B.n45 VSUBS 0.007403f
C80 B.n46 VSUBS 0.007403f
C81 B.n47 VSUBS 0.007403f
C82 B.n48 VSUBS 0.007403f
C83 B.n49 VSUBS 0.007403f
C84 B.n50 VSUBS 0.007403f
C85 B.n51 VSUBS 0.007403f
C86 B.n52 VSUBS 0.007403f
C87 B.n53 VSUBS 0.007403f
C88 B.n54 VSUBS 0.007403f
C89 B.n55 VSUBS 0.007403f
C90 B.n56 VSUBS 0.007403f
C91 B.n57 VSUBS 0.007403f
C92 B.n58 VSUBS 0.007403f
C93 B.n59 VSUBS 0.007403f
C94 B.n60 VSUBS 0.007403f
C95 B.n61 VSUBS 0.007403f
C96 B.n62 VSUBS 0.018515f
C97 B.n63 VSUBS 0.007403f
C98 B.n64 VSUBS 0.007403f
C99 B.n65 VSUBS 0.007403f
C100 B.n66 VSUBS 0.007403f
C101 B.n67 VSUBS 0.007403f
C102 B.n68 VSUBS 0.007403f
C103 B.n69 VSUBS 0.007403f
C104 B.n70 VSUBS 0.007403f
C105 B.n71 VSUBS 0.007403f
C106 B.n72 VSUBS 0.007403f
C107 B.n73 VSUBS 0.007403f
C108 B.n74 VSUBS 0.007403f
C109 B.n75 VSUBS 0.007403f
C110 B.n76 VSUBS 0.007403f
C111 B.n77 VSUBS 0.007403f
C112 B.n78 VSUBS 0.007403f
C113 B.n79 VSUBS 0.007403f
C114 B.n80 VSUBS 0.007403f
C115 B.n81 VSUBS 0.017709f
C116 B.n82 VSUBS 0.007403f
C117 B.n83 VSUBS 0.007403f
C118 B.n84 VSUBS 0.007403f
C119 B.n85 VSUBS 0.007403f
C120 B.n86 VSUBS 0.007403f
C121 B.n87 VSUBS 0.007403f
C122 B.n88 VSUBS 0.007403f
C123 B.n89 VSUBS 0.007403f
C124 B.n90 VSUBS 0.007403f
C125 B.n91 VSUBS 0.007403f
C126 B.n92 VSUBS 0.007403f
C127 B.n93 VSUBS 0.007403f
C128 B.n94 VSUBS 0.007403f
C129 B.n95 VSUBS 0.007403f
C130 B.n96 VSUBS 0.007403f
C131 B.n97 VSUBS 0.007403f
C132 B.n98 VSUBS 0.007403f
C133 B.n99 VSUBS 0.007403f
C134 B.n100 VSUBS 0.007403f
C135 B.n101 VSUBS 0.007403f
C136 B.t10 VSUBS 0.408208f
C137 B.t11 VSUBS 0.416158f
C138 B.t9 VSUBS 0.318363f
C139 B.n102 VSUBS 0.134963f
C140 B.n103 VSUBS 0.067248f
C141 B.n104 VSUBS 0.017151f
C142 B.n105 VSUBS 0.007403f
C143 B.n106 VSUBS 0.007403f
C144 B.n107 VSUBS 0.007403f
C145 B.n108 VSUBS 0.007403f
C146 B.n109 VSUBS 0.007403f
C147 B.t1 VSUBS 0.408215f
C148 B.t2 VSUBS 0.416165f
C149 B.t0 VSUBS 0.318363f
C150 B.n110 VSUBS 0.134956f
C151 B.n111 VSUBS 0.06724f
C152 B.n112 VSUBS 0.007403f
C153 B.n113 VSUBS 0.007403f
C154 B.n114 VSUBS 0.007403f
C155 B.n115 VSUBS 0.007403f
C156 B.n116 VSUBS 0.007403f
C157 B.n117 VSUBS 0.007403f
C158 B.n118 VSUBS 0.007403f
C159 B.n119 VSUBS 0.007403f
C160 B.n120 VSUBS 0.007403f
C161 B.n121 VSUBS 0.007403f
C162 B.n122 VSUBS 0.007403f
C163 B.n123 VSUBS 0.007403f
C164 B.n124 VSUBS 0.007403f
C165 B.n125 VSUBS 0.007403f
C166 B.n126 VSUBS 0.007403f
C167 B.n127 VSUBS 0.007403f
C168 B.n128 VSUBS 0.007403f
C169 B.n129 VSUBS 0.007403f
C170 B.n130 VSUBS 0.007403f
C171 B.n131 VSUBS 0.007403f
C172 B.n132 VSUBS 0.017709f
C173 B.n133 VSUBS 0.007403f
C174 B.n134 VSUBS 0.007403f
C175 B.n135 VSUBS 0.007403f
C176 B.n136 VSUBS 0.007403f
C177 B.n137 VSUBS 0.007403f
C178 B.n138 VSUBS 0.007403f
C179 B.n139 VSUBS 0.007403f
C180 B.n140 VSUBS 0.007403f
C181 B.n141 VSUBS 0.007403f
C182 B.n142 VSUBS 0.007403f
C183 B.n143 VSUBS 0.007403f
C184 B.n144 VSUBS 0.007403f
C185 B.n145 VSUBS 0.007403f
C186 B.n146 VSUBS 0.007403f
C187 B.n147 VSUBS 0.007403f
C188 B.n148 VSUBS 0.007403f
C189 B.n149 VSUBS 0.007403f
C190 B.n150 VSUBS 0.007403f
C191 B.n151 VSUBS 0.007403f
C192 B.n152 VSUBS 0.007403f
C193 B.n153 VSUBS 0.007403f
C194 B.n154 VSUBS 0.007403f
C195 B.n155 VSUBS 0.007403f
C196 B.n156 VSUBS 0.007403f
C197 B.n157 VSUBS 0.007403f
C198 B.n158 VSUBS 0.007403f
C199 B.n159 VSUBS 0.007403f
C200 B.n160 VSUBS 0.007403f
C201 B.n161 VSUBS 0.007403f
C202 B.n162 VSUBS 0.007403f
C203 B.n163 VSUBS 0.007403f
C204 B.n164 VSUBS 0.007403f
C205 B.n165 VSUBS 0.007403f
C206 B.n166 VSUBS 0.007403f
C207 B.n167 VSUBS 0.017709f
C208 B.n168 VSUBS 0.018869f
C209 B.n169 VSUBS 0.018869f
C210 B.n170 VSUBS 0.007403f
C211 B.n171 VSUBS 0.007403f
C212 B.n172 VSUBS 0.007403f
C213 B.n173 VSUBS 0.007403f
C214 B.n174 VSUBS 0.007403f
C215 B.n175 VSUBS 0.007403f
C216 B.n176 VSUBS 0.007403f
C217 B.n177 VSUBS 0.007403f
C218 B.n178 VSUBS 0.007403f
C219 B.n179 VSUBS 0.007403f
C220 B.n180 VSUBS 0.007403f
C221 B.n181 VSUBS 0.007403f
C222 B.n182 VSUBS 0.007403f
C223 B.n183 VSUBS 0.007403f
C224 B.n184 VSUBS 0.007403f
C225 B.n185 VSUBS 0.007403f
C226 B.n186 VSUBS 0.007403f
C227 B.n187 VSUBS 0.007403f
C228 B.n188 VSUBS 0.007403f
C229 B.n189 VSUBS 0.007403f
C230 B.n190 VSUBS 0.007403f
C231 B.n191 VSUBS 0.007403f
C232 B.n192 VSUBS 0.007403f
C233 B.n193 VSUBS 0.007403f
C234 B.n194 VSUBS 0.007403f
C235 B.n195 VSUBS 0.007403f
C236 B.n196 VSUBS 0.007403f
C237 B.n197 VSUBS 0.007403f
C238 B.n198 VSUBS 0.007403f
C239 B.n199 VSUBS 0.007403f
C240 B.n200 VSUBS 0.007403f
C241 B.n201 VSUBS 0.007403f
C242 B.n202 VSUBS 0.007403f
C243 B.n203 VSUBS 0.007403f
C244 B.n204 VSUBS 0.007403f
C245 B.n205 VSUBS 0.007403f
C246 B.n206 VSUBS 0.007403f
C247 B.n207 VSUBS 0.007403f
C248 B.n208 VSUBS 0.007403f
C249 B.n209 VSUBS 0.007403f
C250 B.n210 VSUBS 0.007403f
C251 B.n211 VSUBS 0.007403f
C252 B.n212 VSUBS 0.007403f
C253 B.n213 VSUBS 0.007403f
C254 B.n214 VSUBS 0.007403f
C255 B.n215 VSUBS 0.007403f
C256 B.n216 VSUBS 0.007403f
C257 B.n217 VSUBS 0.007403f
C258 B.n218 VSUBS 0.007403f
C259 B.n219 VSUBS 0.007403f
C260 B.n220 VSUBS 0.007403f
C261 B.n221 VSUBS 0.007403f
C262 B.n222 VSUBS 0.007403f
C263 B.n223 VSUBS 0.007403f
C264 B.n224 VSUBS 0.007403f
C265 B.n225 VSUBS 0.007403f
C266 B.n226 VSUBS 0.007403f
C267 B.n227 VSUBS 0.007403f
C268 B.n228 VSUBS 0.007403f
C269 B.n229 VSUBS 0.006967f
C270 B.n230 VSUBS 0.017151f
C271 B.n231 VSUBS 0.004137f
C272 B.n232 VSUBS 0.007403f
C273 B.n233 VSUBS 0.007403f
C274 B.n234 VSUBS 0.007403f
C275 B.n235 VSUBS 0.007403f
C276 B.n236 VSUBS 0.007403f
C277 B.n237 VSUBS 0.007403f
C278 B.n238 VSUBS 0.007403f
C279 B.n239 VSUBS 0.007403f
C280 B.n240 VSUBS 0.007403f
C281 B.n241 VSUBS 0.007403f
C282 B.n242 VSUBS 0.007403f
C283 B.n243 VSUBS 0.007403f
C284 B.n244 VSUBS 0.004137f
C285 B.n245 VSUBS 0.007403f
C286 B.n246 VSUBS 0.007403f
C287 B.n247 VSUBS 0.006967f
C288 B.n248 VSUBS 0.007403f
C289 B.n249 VSUBS 0.007403f
C290 B.n250 VSUBS 0.007403f
C291 B.n251 VSUBS 0.007403f
C292 B.n252 VSUBS 0.007403f
C293 B.n253 VSUBS 0.007403f
C294 B.n254 VSUBS 0.007403f
C295 B.n255 VSUBS 0.007403f
C296 B.n256 VSUBS 0.007403f
C297 B.n257 VSUBS 0.007403f
C298 B.n258 VSUBS 0.007403f
C299 B.n259 VSUBS 0.007403f
C300 B.n260 VSUBS 0.007403f
C301 B.n261 VSUBS 0.007403f
C302 B.n262 VSUBS 0.007403f
C303 B.n263 VSUBS 0.007403f
C304 B.n264 VSUBS 0.007403f
C305 B.n265 VSUBS 0.007403f
C306 B.n266 VSUBS 0.007403f
C307 B.n267 VSUBS 0.007403f
C308 B.n268 VSUBS 0.007403f
C309 B.n269 VSUBS 0.007403f
C310 B.n270 VSUBS 0.007403f
C311 B.n271 VSUBS 0.007403f
C312 B.n272 VSUBS 0.007403f
C313 B.n273 VSUBS 0.007403f
C314 B.n274 VSUBS 0.007403f
C315 B.n275 VSUBS 0.007403f
C316 B.n276 VSUBS 0.007403f
C317 B.n277 VSUBS 0.007403f
C318 B.n278 VSUBS 0.007403f
C319 B.n279 VSUBS 0.007403f
C320 B.n280 VSUBS 0.007403f
C321 B.n281 VSUBS 0.007403f
C322 B.n282 VSUBS 0.007403f
C323 B.n283 VSUBS 0.007403f
C324 B.n284 VSUBS 0.007403f
C325 B.n285 VSUBS 0.007403f
C326 B.n286 VSUBS 0.007403f
C327 B.n287 VSUBS 0.007403f
C328 B.n288 VSUBS 0.007403f
C329 B.n289 VSUBS 0.007403f
C330 B.n290 VSUBS 0.007403f
C331 B.n291 VSUBS 0.007403f
C332 B.n292 VSUBS 0.007403f
C333 B.n293 VSUBS 0.007403f
C334 B.n294 VSUBS 0.007403f
C335 B.n295 VSUBS 0.007403f
C336 B.n296 VSUBS 0.007403f
C337 B.n297 VSUBS 0.007403f
C338 B.n298 VSUBS 0.007403f
C339 B.n299 VSUBS 0.007403f
C340 B.n300 VSUBS 0.007403f
C341 B.n301 VSUBS 0.007403f
C342 B.n302 VSUBS 0.007403f
C343 B.n303 VSUBS 0.007403f
C344 B.n304 VSUBS 0.007403f
C345 B.n305 VSUBS 0.007403f
C346 B.n306 VSUBS 0.018869f
C347 B.n307 VSUBS 0.018869f
C348 B.n308 VSUBS 0.017709f
C349 B.n309 VSUBS 0.007403f
C350 B.n310 VSUBS 0.007403f
C351 B.n311 VSUBS 0.007403f
C352 B.n312 VSUBS 0.007403f
C353 B.n313 VSUBS 0.007403f
C354 B.n314 VSUBS 0.007403f
C355 B.n315 VSUBS 0.007403f
C356 B.n316 VSUBS 0.007403f
C357 B.n317 VSUBS 0.007403f
C358 B.n318 VSUBS 0.007403f
C359 B.n319 VSUBS 0.007403f
C360 B.n320 VSUBS 0.007403f
C361 B.n321 VSUBS 0.007403f
C362 B.n322 VSUBS 0.007403f
C363 B.n323 VSUBS 0.007403f
C364 B.n324 VSUBS 0.007403f
C365 B.n325 VSUBS 0.007403f
C366 B.n326 VSUBS 0.007403f
C367 B.n327 VSUBS 0.007403f
C368 B.n328 VSUBS 0.007403f
C369 B.n329 VSUBS 0.007403f
C370 B.n330 VSUBS 0.007403f
C371 B.n331 VSUBS 0.007403f
C372 B.n332 VSUBS 0.007403f
C373 B.n333 VSUBS 0.007403f
C374 B.n334 VSUBS 0.007403f
C375 B.n335 VSUBS 0.007403f
C376 B.n336 VSUBS 0.007403f
C377 B.n337 VSUBS 0.007403f
C378 B.n338 VSUBS 0.007403f
C379 B.n339 VSUBS 0.007403f
C380 B.n340 VSUBS 0.007403f
C381 B.n341 VSUBS 0.007403f
C382 B.n342 VSUBS 0.007403f
C383 B.n343 VSUBS 0.007403f
C384 B.n344 VSUBS 0.007403f
C385 B.n345 VSUBS 0.007403f
C386 B.n346 VSUBS 0.007403f
C387 B.n347 VSUBS 0.007403f
C388 B.n348 VSUBS 0.007403f
C389 B.n349 VSUBS 0.007403f
C390 B.n350 VSUBS 0.007403f
C391 B.n351 VSUBS 0.007403f
C392 B.n352 VSUBS 0.007403f
C393 B.n353 VSUBS 0.007403f
C394 B.n354 VSUBS 0.007403f
C395 B.n355 VSUBS 0.007403f
C396 B.n356 VSUBS 0.007403f
C397 B.n357 VSUBS 0.007403f
C398 B.n358 VSUBS 0.007403f
C399 B.n359 VSUBS 0.007403f
C400 B.n360 VSUBS 0.007403f
C401 B.n361 VSUBS 0.007403f
C402 B.n362 VSUBS 0.007403f
C403 B.n363 VSUBS 0.007403f
C404 B.n364 VSUBS 0.007403f
C405 B.n365 VSUBS 0.017709f
C406 B.n366 VSUBS 0.018869f
C407 B.n367 VSUBS 0.018063f
C408 B.n368 VSUBS 0.007403f
C409 B.n369 VSUBS 0.007403f
C410 B.n370 VSUBS 0.007403f
C411 B.n371 VSUBS 0.007403f
C412 B.n372 VSUBS 0.007403f
C413 B.n373 VSUBS 0.007403f
C414 B.n374 VSUBS 0.007403f
C415 B.n375 VSUBS 0.007403f
C416 B.n376 VSUBS 0.007403f
C417 B.n377 VSUBS 0.007403f
C418 B.n378 VSUBS 0.007403f
C419 B.n379 VSUBS 0.007403f
C420 B.n380 VSUBS 0.007403f
C421 B.n381 VSUBS 0.007403f
C422 B.n382 VSUBS 0.007403f
C423 B.n383 VSUBS 0.007403f
C424 B.n384 VSUBS 0.007403f
C425 B.n385 VSUBS 0.007403f
C426 B.n386 VSUBS 0.007403f
C427 B.n387 VSUBS 0.007403f
C428 B.n388 VSUBS 0.007403f
C429 B.n389 VSUBS 0.007403f
C430 B.n390 VSUBS 0.007403f
C431 B.n391 VSUBS 0.007403f
C432 B.n392 VSUBS 0.007403f
C433 B.n393 VSUBS 0.007403f
C434 B.n394 VSUBS 0.007403f
C435 B.n395 VSUBS 0.007403f
C436 B.n396 VSUBS 0.007403f
C437 B.n397 VSUBS 0.007403f
C438 B.n398 VSUBS 0.007403f
C439 B.n399 VSUBS 0.007403f
C440 B.n400 VSUBS 0.007403f
C441 B.n401 VSUBS 0.007403f
C442 B.n402 VSUBS 0.007403f
C443 B.n403 VSUBS 0.007403f
C444 B.n404 VSUBS 0.007403f
C445 B.n405 VSUBS 0.007403f
C446 B.n406 VSUBS 0.007403f
C447 B.n407 VSUBS 0.007403f
C448 B.n408 VSUBS 0.007403f
C449 B.n409 VSUBS 0.007403f
C450 B.n410 VSUBS 0.007403f
C451 B.n411 VSUBS 0.007403f
C452 B.n412 VSUBS 0.007403f
C453 B.n413 VSUBS 0.007403f
C454 B.n414 VSUBS 0.007403f
C455 B.n415 VSUBS 0.007403f
C456 B.n416 VSUBS 0.007403f
C457 B.n417 VSUBS 0.007403f
C458 B.n418 VSUBS 0.007403f
C459 B.n419 VSUBS 0.007403f
C460 B.n420 VSUBS 0.007403f
C461 B.n421 VSUBS 0.007403f
C462 B.n422 VSUBS 0.007403f
C463 B.n423 VSUBS 0.007403f
C464 B.n424 VSUBS 0.007403f
C465 B.n425 VSUBS 0.007403f
C466 B.n426 VSUBS 0.007403f
C467 B.n427 VSUBS 0.006967f
C468 B.n428 VSUBS 0.017151f
C469 B.n429 VSUBS 0.004137f
C470 B.n430 VSUBS 0.007403f
C471 B.n431 VSUBS 0.007403f
C472 B.n432 VSUBS 0.007403f
C473 B.n433 VSUBS 0.007403f
C474 B.n434 VSUBS 0.007403f
C475 B.n435 VSUBS 0.007403f
C476 B.n436 VSUBS 0.007403f
C477 B.n437 VSUBS 0.007403f
C478 B.n438 VSUBS 0.007403f
C479 B.n439 VSUBS 0.007403f
C480 B.n440 VSUBS 0.007403f
C481 B.n441 VSUBS 0.007403f
C482 B.n442 VSUBS 0.004137f
C483 B.n443 VSUBS 0.007403f
C484 B.n444 VSUBS 0.007403f
C485 B.n445 VSUBS 0.006967f
C486 B.n446 VSUBS 0.007403f
C487 B.n447 VSUBS 0.007403f
C488 B.n448 VSUBS 0.007403f
C489 B.n449 VSUBS 0.007403f
C490 B.n450 VSUBS 0.007403f
C491 B.n451 VSUBS 0.007403f
C492 B.n452 VSUBS 0.007403f
C493 B.n453 VSUBS 0.007403f
C494 B.n454 VSUBS 0.007403f
C495 B.n455 VSUBS 0.007403f
C496 B.n456 VSUBS 0.007403f
C497 B.n457 VSUBS 0.007403f
C498 B.n458 VSUBS 0.007403f
C499 B.n459 VSUBS 0.007403f
C500 B.n460 VSUBS 0.007403f
C501 B.n461 VSUBS 0.007403f
C502 B.n462 VSUBS 0.007403f
C503 B.n463 VSUBS 0.007403f
C504 B.n464 VSUBS 0.007403f
C505 B.n465 VSUBS 0.007403f
C506 B.n466 VSUBS 0.007403f
C507 B.n467 VSUBS 0.007403f
C508 B.n468 VSUBS 0.007403f
C509 B.n469 VSUBS 0.007403f
C510 B.n470 VSUBS 0.007403f
C511 B.n471 VSUBS 0.007403f
C512 B.n472 VSUBS 0.007403f
C513 B.n473 VSUBS 0.007403f
C514 B.n474 VSUBS 0.007403f
C515 B.n475 VSUBS 0.007403f
C516 B.n476 VSUBS 0.007403f
C517 B.n477 VSUBS 0.007403f
C518 B.n478 VSUBS 0.007403f
C519 B.n479 VSUBS 0.007403f
C520 B.n480 VSUBS 0.007403f
C521 B.n481 VSUBS 0.007403f
C522 B.n482 VSUBS 0.007403f
C523 B.n483 VSUBS 0.007403f
C524 B.n484 VSUBS 0.007403f
C525 B.n485 VSUBS 0.007403f
C526 B.n486 VSUBS 0.007403f
C527 B.n487 VSUBS 0.007403f
C528 B.n488 VSUBS 0.007403f
C529 B.n489 VSUBS 0.007403f
C530 B.n490 VSUBS 0.007403f
C531 B.n491 VSUBS 0.007403f
C532 B.n492 VSUBS 0.007403f
C533 B.n493 VSUBS 0.007403f
C534 B.n494 VSUBS 0.007403f
C535 B.n495 VSUBS 0.007403f
C536 B.n496 VSUBS 0.007403f
C537 B.n497 VSUBS 0.007403f
C538 B.n498 VSUBS 0.007403f
C539 B.n499 VSUBS 0.007403f
C540 B.n500 VSUBS 0.007403f
C541 B.n501 VSUBS 0.007403f
C542 B.n502 VSUBS 0.007403f
C543 B.n503 VSUBS 0.007403f
C544 B.n504 VSUBS 0.018869f
C545 B.n505 VSUBS 0.018869f
C546 B.n506 VSUBS 0.017709f
C547 B.n507 VSUBS 0.007403f
C548 B.n508 VSUBS 0.007403f
C549 B.n509 VSUBS 0.007403f
C550 B.n510 VSUBS 0.007403f
C551 B.n511 VSUBS 0.007403f
C552 B.n512 VSUBS 0.007403f
C553 B.n513 VSUBS 0.007403f
C554 B.n514 VSUBS 0.007403f
C555 B.n515 VSUBS 0.007403f
C556 B.n516 VSUBS 0.007403f
C557 B.n517 VSUBS 0.007403f
C558 B.n518 VSUBS 0.007403f
C559 B.n519 VSUBS 0.007403f
C560 B.n520 VSUBS 0.007403f
C561 B.n521 VSUBS 0.007403f
C562 B.n522 VSUBS 0.007403f
C563 B.n523 VSUBS 0.007403f
C564 B.n524 VSUBS 0.007403f
C565 B.n525 VSUBS 0.007403f
C566 B.n526 VSUBS 0.007403f
C567 B.n527 VSUBS 0.007403f
C568 B.n528 VSUBS 0.007403f
C569 B.n529 VSUBS 0.007403f
C570 B.n530 VSUBS 0.007403f
C571 B.n531 VSUBS 0.007403f
C572 B.n532 VSUBS 0.007403f
C573 B.n533 VSUBS 0.007403f
C574 B.n534 VSUBS 0.007403f
C575 B.n535 VSUBS 0.016762f
C576 VDD1.t5 VSUBS 2.29094f
C577 VDD1.t2 VSUBS 2.29007f
C578 VDD1.t3 VSUBS 0.223902f
C579 VDD1.t4 VSUBS 0.223902f
C580 VDD1.n0 VSUBS 1.7506f
C581 VDD1.n1 VSUBS 2.52156f
C582 VDD1.t0 VSUBS 0.223902f
C583 VDD1.t1 VSUBS 0.223902f
C584 VDD1.n2 VSUBS 1.74956f
C585 VDD1.n3 VSUBS 2.36629f
C586 VP.n0 VSUBS 0.080403f
C587 VP.t0 VSUBS 1.2914f
C588 VP.n1 VSUBS 0.485229f
C589 VP.t4 VSUBS 1.26664f
C590 VP.t5 VSUBS 1.26664f
C591 VP.n2 VSUBS 0.522383f
C592 VP.n3 VSUBS 0.508678f
C593 VP.n4 VSUBS 2.5824f
C594 VP.n5 VSUBS 2.4566f
C595 VP.t3 VSUBS 1.26664f
C596 VP.n6 VSUBS 0.508678f
C597 VP.t2 VSUBS 1.26664f
C598 VP.n7 VSUBS 0.522383f
C599 VP.t1 VSUBS 1.26664f
C600 VP.n8 VSUBS 0.508678f
C601 VP.n9 VSUBS 0.067f
C602 VTAIL.t8 VSUBS 0.276742f
C603 VTAIL.t7 VSUBS 0.276742f
C604 VTAIL.n0 VSUBS 2.01114f
C605 VTAIL.n1 VSUBS 0.765784f
C606 VTAIL.t1 VSUBS 2.65638f
C607 VTAIL.n2 VSUBS 0.9282f
C608 VTAIL.t5 VSUBS 0.276742f
C609 VTAIL.t3 VSUBS 0.276742f
C610 VTAIL.n3 VSUBS 2.01114f
C611 VTAIL.n4 VSUBS 2.26476f
C612 VTAIL.t9 VSUBS 0.276742f
C613 VTAIL.t11 VSUBS 0.276742f
C614 VTAIL.n5 VSUBS 2.01115f
C615 VTAIL.n6 VSUBS 2.26476f
C616 VTAIL.t10 VSUBS 2.65638f
C617 VTAIL.n7 VSUBS 0.928192f
C618 VTAIL.t2 VSUBS 0.276742f
C619 VTAIL.t4 VSUBS 0.276742f
C620 VTAIL.n8 VSUBS 2.01115f
C621 VTAIL.n9 VSUBS 0.818681f
C622 VTAIL.t0 VSUBS 2.65638f
C623 VTAIL.n10 VSUBS 2.29635f
C624 VTAIL.t6 VSUBS 2.65638f
C625 VTAIL.n11 VSUBS 2.27134f
C626 VDD2.t2 VSUBS 2.27231f
C627 VDD2.t1 VSUBS 0.222165f
C628 VDD2.t5 VSUBS 0.222165f
C629 VDD2.n0 VSUBS 1.73702f
C630 VDD2.n1 VSUBS 2.43068f
C631 VDD2.t4 VSUBS 2.26834f
C632 VDD2.n2 VSUBS 2.38288f
C633 VDD2.t0 VSUBS 0.222165f
C634 VDD2.t3 VSUBS 0.222165f
C635 VDD2.n3 VSUBS 1.73699f
C636 VN.t3 VSUBS 1.25223f
C637 VN.n0 VSUBS 0.47051f
C638 VN.t4 VSUBS 1.22822f
C639 VN.n1 VSUBS 0.506537f
C640 VN.t5 VSUBS 1.22822f
C641 VN.n2 VSUBS 0.493247f
C642 VN.n3 VSUBS 0.238583f
C643 VN.t1 VSUBS 1.25223f
C644 VN.n4 VSUBS 0.47051f
C645 VN.t0 VSUBS 1.22822f
C646 VN.n5 VSUBS 0.506537f
C647 VN.t2 VSUBS 1.22822f
C648 VN.n6 VSUBS 0.493247f
C649 VN.n7 VSUBS 2.54258f
.ends

