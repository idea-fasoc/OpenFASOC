* NGSPICE file created from tg_sample_0002.ext - technology: sky130A

.subckt tg_sample_0002 VIN VGN VGP VSS VCC VOUT
X0 VOUT.t1 VGP.t0 VIN.t1 VCC.t1 sky130_fd_pr__pfet_01v8 ad=0.66 pd=4.33 as=1.56 ps=8.78 w=4 l=0.18
X1 VIN.t0 VGP.t1 VOUT.t0 VCC.t0 sky130_fd_pr__pfet_01v8 ad=1.56 pd=8.78 as=0.66 ps=4.33 w=4 l=0.18
X2 VCC.t9 VCC.t6 VCC.t8 VCC.t7 sky130_fd_pr__pfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=0.18
X3 VSS.t8 VSS.t5 VSS.t7 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.18
X4 VOUT.t2 VGN.t0 VIN.t2 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.78 ps=4.78 w=2 l=0.18
X5 VIN.t3 VGN.t1 VOUT.t3 VSS.t9 sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0.33 ps=2.33 w=2 l=0.18
X6 VSS.t4 VSS.t1 VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.78 pd=4.78 as=0 ps=0 w=2 l=0.18
X7 VCC.t5 VCC.t2 VCC.t4 VCC.t3 sky130_fd_pr__pfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=0.18
R0 VGP.n0 VGP.t0 746.857
R1 VGP.n0 VGP.t1 746.857
R2 VGP VGP.n0 161.381
R3 VIN.n14 VIN.n0 756.745
R4 VIN.n33 VIN.n19 756.745
R5 VIN.n7 VIN.n6 585
R6 VIN.n4 VIN.n3 585
R7 VIN.n13 VIN.n12 585
R8 VIN.n15 VIN.n14 585
R9 VIN.n26 VIN.n25 585
R10 VIN.n23 VIN.n22 585
R11 VIN.n32 VIN.n31 585
R12 VIN.n34 VIN.n33 585
R13 VIN.t1 VIN.n5 330.707
R14 VIN.t0 VIN.n24 330.707
R15 VIN.n41 VIN.n39 289.615
R16 VIN.n48 VIN.n46 289.615
R17 VIN.n42 VIN.n41 185
R18 VIN.n49 VIN.n48 185
R19 VIN.n6 VIN.n3 171.744
R20 VIN.n13 VIN.n3 171.744
R21 VIN.n14 VIN.n13 171.744
R22 VIN.n25 VIN.n22 171.744
R23 VIN.n32 VIN.n22 171.744
R24 VIN.n33 VIN.n32 171.744
R25 VIN.t2 VIN.n40 167.117
R26 VIN.t3 VIN.n47 167.117
R27 VIN.n6 VIN.t1 85.8723
R28 VIN.n25 VIN.t0 85.8723
R29 VIN.n41 VIN.t2 52.3082
R30 VIN.n48 VIN.t3 52.3082
R31 VIN.n38 VIN.n18 35.728
R32 VIN.n38 VIN.n37 35.2884
R33 VIN.n53 VIN.n45 31.8492
R34 VIN.n53 VIN.n52 31.4096
R35 VIN.n7 VIN.n5 16.3201
R36 VIN.n26 VIN.n24 16.3201
R37 VIN.n8 VIN.n4 12.8005
R38 VIN.n27 VIN.n23 12.8005
R39 VIN.n12 VIN.n11 12.0247
R40 VIN.n31 VIN.n30 12.0247
R41 VIN VIN.n38 11.3669
R42 VIN.n15 VIN.n2 11.249
R43 VIN.n34 VIN.n21 11.249
R44 VIN.n16 VIN.n0 10.4732
R45 VIN.n35 VIN.n19 10.4732
R46 VIN.n42 VIN.n40 9.71174
R47 VIN.n49 VIN.n47 9.71174
R48 VIN.n45 VIN.n44 9.45567
R49 VIN.n52 VIN.n51 9.45567
R50 VIN.n18 VIN.n17 9.45567
R51 VIN.n37 VIN.n36 9.45567
R52 VIN.n44 VIN.n43 9.3005
R53 VIN.n51 VIN.n50 9.3005
R54 VIN.n17 VIN.n16 9.3005
R55 VIN.n2 VIN.n1 9.3005
R56 VIN.n11 VIN.n10 9.3005
R57 VIN.n9 VIN.n8 9.3005
R58 VIN.n36 VIN.n35 9.3005
R59 VIN.n21 VIN.n20 9.3005
R60 VIN.n30 VIN.n29 9.3005
R61 VIN.n28 VIN.n27 9.3005
R62 VIN.n45 VIN.n39 8.14595
R63 VIN.n52 VIN.n46 8.14595
R64 VIN.n43 VIN.n42 7.3702
R65 VIN.n50 VIN.n49 7.3702
R66 VIN.n43 VIN.n39 5.81868
R67 VIN.n50 VIN.n46 5.81868
R68 VIN.n9 VIN.n5 3.78097
R69 VIN.n28 VIN.n24 3.78097
R70 VIN.n18 VIN.n0 3.49141
R71 VIN.n37 VIN.n19 3.49141
R72 VIN.n44 VIN.n40 3.44771
R73 VIN.n51 VIN.n47 3.44771
R74 VIN.n16 VIN.n15 2.71565
R75 VIN.n35 VIN.n34 2.71565
R76 VIN.n12 VIN.n2 1.93989
R77 VIN.n31 VIN.n21 1.93989
R78 VIN.n11 VIN.n4 1.16414
R79 VIN.n30 VIN.n23 1.16414
R80 VIN.n8 VIN.n7 0.388379
R81 VIN.n27 VIN.n26 0.388379
R82 VIN.n10 VIN.n9 0.155672
R83 VIN.n10 VIN.n1 0.155672
R84 VIN.n17 VIN.n1 0.155672
R85 VIN.n29 VIN.n28 0.155672
R86 VIN.n29 VIN.n20 0.155672
R87 VIN.n36 VIN.n20 0.155672
R88 VIN VIN.n53 0.00481034
R89 VOUT VOUT.n0 117.01
R90 VOUT VOUT.n1 111.775
R91 VOUT.n1 VOUT.t3 9.9005
R92 VOUT.n1 VOUT.t2 9.9005
R93 VOUT.n0 VOUT.t0 8.12675
R94 VOUT.n0 VOUT.t1 8.12675
R95 VCC.n118 VCC.t2 778.601
R96 VCC.n44 VCC.t6 778.601
R97 VCC.n158 VCC.n9 370.245
R98 VCC.n156 VCC.n12 370.245
R99 VCC.n79 VCC.n30 370.245
R100 VCC.n76 VCC.n29 370.245
R101 VCC.n118 VCC.t4 245.52
R102 VCC.n44 VCC.t9 245.52
R103 VCC.n119 VCC.t5 235.63
R104 VCC.n45 VCC.t8 235.63
R105 VCC.n156 VCC.n155 185
R106 VCC.n157 VCC.n156 185
R107 VCC.n13 VCC.n11 185
R108 VCC.n103 VCC.n11 185
R109 VCC.n106 VCC.n105 185
R110 VCC.n105 VCC.n104 185
R111 VCC.n16 VCC.n15 185
R112 VCC.n102 VCC.n16 185
R113 VCC.n100 VCC.n99 185
R114 VCC.n101 VCC.n100 185
R115 VCC.n19 VCC.n18 185
R116 VCC.n18 VCC.n17 185
R117 VCC.n95 VCC.n94 185
R118 VCC.n94 VCC.n93 185
R119 VCC.n22 VCC.n21 185
R120 VCC.n23 VCC.n22 185
R121 VCC.n84 VCC.n83 185
R122 VCC.n85 VCC.n84 185
R123 VCC.n31 VCC.n30 185
R124 VCC.n41 VCC.n30 185
R125 VCC.n29 VCC.n28 185
R126 VCC.n41 VCC.n29 185
R127 VCC.n87 VCC.n86 185
R128 VCC.n86 VCC.n85 185
R129 VCC.n26 VCC.n24 185
R130 VCC.n24 VCC.n23 185
R131 VCC.n92 VCC.n91 185
R132 VCC.n93 VCC.n92 185
R133 VCC.n25 VCC.n2 185
R134 VCC.n25 VCC.n17 185
R135 VCC.n165 VCC.n3 185
R136 VCC.n101 VCC.n3 185
R137 VCC.n164 VCC.n4 185
R138 VCC.n102 VCC.n4 185
R139 VCC.n163 VCC.n5 185
R140 VCC.n104 VCC.n5 185
R141 VCC.n8 VCC.n6 185
R142 VCC.n103 VCC.n8 185
R143 VCC.n159 VCC.n158 185
R144 VCC.n158 VCC.n157 185
R145 VCC.n153 VCC.n12 185
R146 VCC.n152 VCC.n151 185
R147 VCC.n149 VCC.n109 185
R148 VCC.n147 VCC.n146 185
R149 VCC.n145 VCC.n110 185
R150 VCC.n144 VCC.n143 185
R151 VCC.n141 VCC.n111 185
R152 VCC.n139 VCC.n138 185
R153 VCC.n137 VCC.n112 185
R154 VCC.n136 VCC.n135 185
R155 VCC.n133 VCC.n113 185
R156 VCC.n131 VCC.n130 185
R157 VCC.n129 VCC.n114 185
R158 VCC.n128 VCC.n127 185
R159 VCC.n125 VCC.n115 185
R160 VCC.n123 VCC.n122 185
R161 VCC.n120 VCC.n117 185
R162 VCC.n9 VCC.n7 185
R163 VCC.n76 VCC.n75 185
R164 VCC.n74 VCC.n43 185
R165 VCC.n72 VCC.n42 185
R166 VCC.n78 VCC.n42 185
R167 VCC.n71 VCC.n70 185
R168 VCC.n69 VCC.n68 185
R169 VCC.n67 VCC.n66 185
R170 VCC.n65 VCC.n64 185
R171 VCC.n63 VCC.n62 185
R172 VCC.n61 VCC.n60 185
R173 VCC.n59 VCC.n58 185
R174 VCC.n57 VCC.n56 185
R175 VCC.n55 VCC.n54 185
R176 VCC.n53 VCC.n52 185
R177 VCC.n51 VCC.n50 185
R178 VCC.n49 VCC.n48 185
R179 VCC.n47 VCC.n46 185
R180 VCC.n33 VCC.n32 185
R181 VCC.n80 VCC.n79 185
R182 VCC.n79 VCC.n78 185
R183 VCC.n84 VCC.n30 146.341
R184 VCC.n84 VCC.n22 146.341
R185 VCC.n94 VCC.n22 146.341
R186 VCC.n94 VCC.n18 146.341
R187 VCC.n100 VCC.n18 146.341
R188 VCC.n100 VCC.n16 146.341
R189 VCC.n105 VCC.n16 146.341
R190 VCC.n105 VCC.n11 146.341
R191 VCC.n156 VCC.n11 146.341
R192 VCC.n86 VCC.n29 146.341
R193 VCC.n86 VCC.n24 146.341
R194 VCC.n92 VCC.n24 146.341
R195 VCC.n92 VCC.n25 146.341
R196 VCC.n25 VCC.n3 146.341
R197 VCC.n4 VCC.n3 146.341
R198 VCC.n5 VCC.n4 146.341
R199 VCC.n8 VCC.n5 146.341
R200 VCC.n158 VCC.n8 146.341
R201 VCC.n123 VCC.n117 99.5127
R202 VCC.n127 VCC.n125 99.5127
R203 VCC.n131 VCC.n114 99.5127
R204 VCC.n135 VCC.n133 99.5127
R205 VCC.n139 VCC.n112 99.5127
R206 VCC.n143 VCC.n141 99.5127
R207 VCC.n147 VCC.n110 99.5127
R208 VCC.n151 VCC.n149 99.5127
R209 VCC.n43 VCC.n42 99.5127
R210 VCC.n70 VCC.n42 99.5127
R211 VCC.n68 VCC.n67 99.5127
R212 VCC.n64 VCC.n63 99.5127
R213 VCC.n60 VCC.n59 99.5127
R214 VCC.n56 VCC.n55 99.5127
R215 VCC.n52 VCC.n51 99.5127
R216 VCC.n48 VCC.n47 99.5127
R217 VCC.n79 VCC.n33 99.5127
R218 VCC.n78 VCC.n41 96.0548
R219 VCC.n157 VCC.n10 96.0548
R220 VCC.n150 VCC.n10 72.8958
R221 VCC.n148 VCC.n10 72.8958
R222 VCC.n142 VCC.n10 72.8958
R223 VCC.n140 VCC.n10 72.8958
R224 VCC.n134 VCC.n10 72.8958
R225 VCC.n132 VCC.n10 72.8958
R226 VCC.n126 VCC.n10 72.8958
R227 VCC.n124 VCC.n10 72.8958
R228 VCC.n116 VCC.n10 72.8958
R229 VCC.n78 VCC.n77 72.8958
R230 VCC.n78 VCC.n34 72.8958
R231 VCC.n78 VCC.n35 72.8958
R232 VCC.n78 VCC.n36 72.8958
R233 VCC.n78 VCC.n37 72.8958
R234 VCC.n78 VCC.n38 72.8958
R235 VCC.n78 VCC.n39 72.8958
R236 VCC.n78 VCC.n40 72.8958
R237 VCC.n85 VCC.n23 58.5702
R238 VCC.n93 VCC.n23 58.5702
R239 VCC.n101 VCC.n17 58.5702
R240 VCC.n104 VCC.n102 58.5702
R241 VCC.n104 VCC.n103 58.5702
R242 VCC.n93 VCC.t0 57.9845
R243 VCC.n102 VCC.t1 57.9845
R244 VCC.n41 VCC.t7 46.2705
R245 VCC.n157 VCC.t3 46.2705
R246 VCC.n117 VCC.n116 39.2114
R247 VCC.n125 VCC.n124 39.2114
R248 VCC.n126 VCC.n114 39.2114
R249 VCC.n133 VCC.n132 39.2114
R250 VCC.n134 VCC.n112 39.2114
R251 VCC.n141 VCC.n140 39.2114
R252 VCC.n142 VCC.n110 39.2114
R253 VCC.n149 VCC.n148 39.2114
R254 VCC.n150 VCC.n12 39.2114
R255 VCC.n77 VCC.n76 39.2114
R256 VCC.n70 VCC.n34 39.2114
R257 VCC.n67 VCC.n35 39.2114
R258 VCC.n63 VCC.n36 39.2114
R259 VCC.n59 VCC.n37 39.2114
R260 VCC.n55 VCC.n38 39.2114
R261 VCC.n51 VCC.n39 39.2114
R262 VCC.n47 VCC.n40 39.2114
R263 VCC.n151 VCC.n150 39.2114
R264 VCC.n148 VCC.n147 39.2114
R265 VCC.n143 VCC.n142 39.2114
R266 VCC.n140 VCC.n139 39.2114
R267 VCC.n135 VCC.n134 39.2114
R268 VCC.n132 VCC.n131 39.2114
R269 VCC.n127 VCC.n126 39.2114
R270 VCC.n124 VCC.n123 39.2114
R271 VCC.n116 VCC.n9 39.2114
R272 VCC.n77 VCC.n43 39.2114
R273 VCC.n68 VCC.n34 39.2114
R274 VCC.n64 VCC.n35 39.2114
R275 VCC.n60 VCC.n36 39.2114
R276 VCC.n56 VCC.n37 39.2114
R277 VCC.n52 VCC.n38 39.2114
R278 VCC.n48 VCC.n39 39.2114
R279 VCC.n40 VCC.n33 39.2114
R280 VCC.n160 VCC.n7 29.8432
R281 VCC.n154 VCC.n153 29.8432
R282 VCC.n75 VCC.n27 29.8432
R283 VCC.n81 VCC.n80 29.8432
R284 VCC.n121 VCC.n119 29.2853
R285 VCC.n73 VCC.n45 29.2853
R286 VCC.n83 VCC.n31 19.3944
R287 VCC.n83 VCC.n21 19.3944
R288 VCC.n95 VCC.n21 19.3944
R289 VCC.n95 VCC.n19 19.3944
R290 VCC.n99 VCC.n19 19.3944
R291 VCC.n99 VCC.n15 19.3944
R292 VCC.n106 VCC.n15 19.3944
R293 VCC.n106 VCC.n13 19.3944
R294 VCC.n155 VCC.n13 19.3944
R295 VCC.n87 VCC.n28 19.3944
R296 VCC.n87 VCC.n26 19.3944
R297 VCC.n91 VCC.n26 19.3944
R298 VCC.n91 VCC.n2 19.3944
R299 VCC.n165 VCC.n2 19.3944
R300 VCC.n165 VCC.n164 19.3944
R301 VCC.n164 VCC.n163 19.3944
R302 VCC.n163 VCC.n6 19.3944
R303 VCC.n159 VCC.n6 19.3944
R304 VCC.n85 VCC.t7 12.3001
R305 VCC.n103 VCC.t3 12.3001
R306 VCC.n120 VCC.n7 10.6151
R307 VCC.n122 VCC.n115 10.6151
R308 VCC.n128 VCC.n115 10.6151
R309 VCC.n129 VCC.n128 10.6151
R310 VCC.n130 VCC.n129 10.6151
R311 VCC.n130 VCC.n113 10.6151
R312 VCC.n136 VCC.n113 10.6151
R313 VCC.n137 VCC.n136 10.6151
R314 VCC.n138 VCC.n137 10.6151
R315 VCC.n138 VCC.n111 10.6151
R316 VCC.n144 VCC.n111 10.6151
R317 VCC.n145 VCC.n144 10.6151
R318 VCC.n146 VCC.n145 10.6151
R319 VCC.n146 VCC.n109 10.6151
R320 VCC.n152 VCC.n109 10.6151
R321 VCC.n153 VCC.n152 10.6151
R322 VCC.n75 VCC.n74 10.6151
R323 VCC.n72 VCC.n71 10.6151
R324 VCC.n71 VCC.n69 10.6151
R325 VCC.n69 VCC.n66 10.6151
R326 VCC.n66 VCC.n65 10.6151
R327 VCC.n65 VCC.n62 10.6151
R328 VCC.n62 VCC.n61 10.6151
R329 VCC.n61 VCC.n58 10.6151
R330 VCC.n58 VCC.n57 10.6151
R331 VCC.n57 VCC.n54 10.6151
R332 VCC.n54 VCC.n53 10.6151
R333 VCC.n53 VCC.n50 10.6151
R334 VCC.n50 VCC.n49 10.6151
R335 VCC.n49 VCC.n46 10.6151
R336 VCC.n46 VCC.n32 10.6151
R337 VCC.n80 VCC.n32 10.6151
R338 VCC.n119 VCC.n118 9.89141
R339 VCC.n45 VCC.n44 9.89141
R340 VCC.n164 VCC.n0 9.3005
R341 VCC.n163 VCC.n162 9.3005
R342 VCC.n161 VCC.n6 9.3005
R343 VCC.n160 VCC.n159 9.3005
R344 VCC.n83 VCC.n82 9.3005
R345 VCC.n21 VCC.n20 9.3005
R346 VCC.n96 VCC.n95 9.3005
R347 VCC.n97 VCC.n19 9.3005
R348 VCC.n99 VCC.n98 9.3005
R349 VCC.n15 VCC.n14 9.3005
R350 VCC.n107 VCC.n106 9.3005
R351 VCC.n108 VCC.n13 9.3005
R352 VCC.n155 VCC.n154 9.3005
R353 VCC.n81 VCC.n31 9.3005
R354 VCC.n28 VCC.n27 9.3005
R355 VCC.n88 VCC.n87 9.3005
R356 VCC.n89 VCC.n26 9.3005
R357 VCC.n91 VCC.n90 9.3005
R358 VCC.n2 VCC.n1 9.3005
R359 VCC VCC.n165 9.3005
R360 VCC.n121 VCC.n120 6.4005
R361 VCC.n74 VCC.n73 6.4005
R362 VCC.n122 VCC.n121 4.21513
R363 VCC.n73 VCC.n72 4.21513
R364 VCC.t0 VCC.n17 0.586197
R365 VCC.t1 VCC.n101 0.586197
R366 VCC VCC.n0 0.152939
R367 VCC.n162 VCC.n0 0.152939
R368 VCC.n162 VCC.n161 0.152939
R369 VCC.n161 VCC.n160 0.152939
R370 VCC.n82 VCC.n81 0.152939
R371 VCC.n82 VCC.n20 0.152939
R372 VCC.n96 VCC.n20 0.152939
R373 VCC.n97 VCC.n96 0.152939
R374 VCC.n98 VCC.n97 0.152939
R375 VCC.n98 VCC.n14 0.152939
R376 VCC.n107 VCC.n14 0.152939
R377 VCC.n108 VCC.n107 0.152939
R378 VCC.n154 VCC.n108 0.152939
R379 VCC.n88 VCC.n27 0.152939
R380 VCC.n89 VCC.n88 0.152939
R381 VCC.n90 VCC.n89 0.152939
R382 VCC.n90 VCC.n1 0.152939
R383 VCC VCC.n1 0.1255
R384 VSS.n314 VSS.n313 5367.03
R385 VSS.n352 VSS.n55 5367.03
R386 VSS.n314 VSS.n72 2953.02
R387 VSS.n322 VSS.n72 2953.02
R388 VSS.n323 VSS.n322 2953.02
R389 VSS.n324 VSS.n323 2953.02
R390 VSS.n324 VSS.n66 2953.02
R391 VSS.n332 VSS.n66 2953.02
R392 VSS.n333 VSS.n332 2953.02
R393 VSS.n334 VSS.n333 2953.02
R394 VSS.n334 VSS.n60 2953.02
R395 VSS.n343 VSS.n60 2953.02
R396 VSS.n344 VSS.n343 2953.02
R397 VSS.n345 VSS.n344 2953.02
R398 VSS.n345 VSS.n55 2953.02
R399 VSS.n313 VSS.n312 1719.54
R400 VSS.n312 VSS.n77 1719.54
R401 VSS.n306 VSS.n77 1719.54
R402 VSS.n306 VSS.n305 1719.54
R403 VSS.n305 VSS.n304 1719.54
R404 VSS.n304 VSS.n81 1719.54
R405 VSS.n298 VSS.n81 1719.54
R406 VSS.n298 VSS.n297 1719.54
R407 VSS.n297 VSS.n296 1719.54
R408 VSS.n296 VSS.n85 1719.54
R409 VSS.n290 VSS.n85 1719.54
R410 VSS.n290 VSS.n289 1719.54
R411 VSS.n289 VSS.n288 1719.54
R412 VSS.n288 VSS.n89 1719.54
R413 VSS.n282 VSS.n89 1719.54
R414 VSS.n282 VSS.n281 1719.54
R415 VSS.n281 VSS.n280 1719.54
R416 VSS.n280 VSS.n93 1719.54
R417 VSS.n274 VSS.n93 1719.54
R418 VSS.n274 VSS.n273 1719.54
R419 VSS.n273 VSS.n272 1719.54
R420 VSS.n272 VSS.n97 1719.54
R421 VSS.n353 VSS.n352 1719.54
R422 VSS.n354 VSS.n353 1719.54
R423 VSS.n354 VSS.n51 1719.54
R424 VSS.n360 VSS.n51 1719.54
R425 VSS.n361 VSS.n360 1719.54
R426 VSS.n362 VSS.n361 1719.54
R427 VSS.n362 VSS.n47 1719.54
R428 VSS.n368 VSS.n47 1719.54
R429 VSS.n369 VSS.n368 1719.54
R430 VSS.n370 VSS.n369 1719.54
R431 VSS.n370 VSS.n43 1719.54
R432 VSS.n376 VSS.n43 1719.54
R433 VSS.n377 VSS.n376 1719.54
R434 VSS.n378 VSS.n377 1719.54
R435 VSS.n378 VSS.n39 1719.54
R436 VSS.n384 VSS.n39 1719.54
R437 VSS.n385 VSS.n384 1719.54
R438 VSS.n386 VSS.n385 1719.54
R439 VSS.n386 VSS.n35 1719.54
R440 VSS.n393 VSS.n35 1719.54
R441 VSS.n394 VSS.n393 1719.54
R442 VSS.n395 VSS.n394 1719.54
R443 VSS.n110 VSS.n97 1668.97
R444 VSS.n395 VSS.n17 1668.97
R445 VSS.n315 VSS.n76 660.672
R446 VSS.n351 VSS.n56 660.672
R447 VSS.n438 VSS.n19 660.672
R448 VSS.n228 VSS.n109 660.672
R449 VSS.n224 VSS.n123 660.672
R450 VSS.n200 VSS.n199 660.672
R451 VSS.n474 VSS.n13 660.672
R452 VSS.n476 VSS.n9 660.672
R453 VSS.n76 VSS.n75 585
R454 VSS.n313 VSS.n76 585
R455 VSS.n311 VSS.n310 585
R456 VSS.n312 VSS.n311 585
R457 VSS.n309 VSS.n78 585
R458 VSS.n78 VSS.n77 585
R459 VSS.n308 VSS.n307 585
R460 VSS.n307 VSS.n306 585
R461 VSS.n80 VSS.n79 585
R462 VSS.n305 VSS.n80 585
R463 VSS.n303 VSS.n302 585
R464 VSS.n304 VSS.n303 585
R465 VSS.n301 VSS.n82 585
R466 VSS.n82 VSS.n81 585
R467 VSS.n300 VSS.n299 585
R468 VSS.n299 VSS.n298 585
R469 VSS.n84 VSS.n83 585
R470 VSS.n297 VSS.n84 585
R471 VSS.n295 VSS.n294 585
R472 VSS.n296 VSS.n295 585
R473 VSS.n293 VSS.n86 585
R474 VSS.n86 VSS.n85 585
R475 VSS.n292 VSS.n291 585
R476 VSS.n291 VSS.n290 585
R477 VSS.n88 VSS.n87 585
R478 VSS.n289 VSS.n88 585
R479 VSS.n287 VSS.n286 585
R480 VSS.n288 VSS.n287 585
R481 VSS.n285 VSS.n90 585
R482 VSS.n90 VSS.n89 585
R483 VSS.n284 VSS.n283 585
R484 VSS.n283 VSS.n282 585
R485 VSS.n92 VSS.n91 585
R486 VSS.n281 VSS.n92 585
R487 VSS.n279 VSS.n278 585
R488 VSS.n280 VSS.n279 585
R489 VSS.n277 VSS.n94 585
R490 VSS.n94 VSS.n93 585
R491 VSS.n276 VSS.n275 585
R492 VSS.n275 VSS.n274 585
R493 VSS.n96 VSS.n95 585
R494 VSS.n273 VSS.n96 585
R495 VSS.n271 VSS.n270 585
R496 VSS.n272 VSS.n271 585
R497 VSS.n269 VSS.n98 585
R498 VSS.n98 VSS.n97 585
R499 VSS.n316 VSS.n315 585
R500 VSS.n315 VSS.n314 585
R501 VSS.n74 VSS.n73 585
R502 VSS.n73 VSS.n72 585
R503 VSS.n321 VSS.n320 585
R504 VSS.n322 VSS.n321 585
R505 VSS.n71 VSS.n70 585
R506 VSS.n323 VSS.n71 585
R507 VSS.n326 VSS.n325 585
R508 VSS.n325 VSS.n324 585
R509 VSS.n68 VSS.n67 585
R510 VSS.n67 VSS.n66 585
R511 VSS.n331 VSS.n330 585
R512 VSS.n332 VSS.n331 585
R513 VSS.n65 VSS.n64 585
R514 VSS.n333 VSS.n65 585
R515 VSS.n336 VSS.n335 585
R516 VSS.n335 VSS.n334 585
R517 VSS.n62 VSS.n61 585
R518 VSS.n61 VSS.n60 585
R519 VSS.n342 VSS.n341 585
R520 VSS.n343 VSS.n342 585
R521 VSS.n59 VSS.n58 585
R522 VSS.n344 VSS.n59 585
R523 VSS.n347 VSS.n346 585
R524 VSS.n346 VSS.n345 585
R525 VSS.n348 VSS.n56 585
R526 VSS.n56 VSS.n55 585
R527 VSS.n396 VSS.n33 585
R528 VSS.n396 VSS.n395 585
R529 VSS.n390 VSS.n34 585
R530 VSS.n394 VSS.n34 585
R531 VSS.n392 VSS.n391 585
R532 VSS.n393 VSS.n392 585
R533 VSS.n389 VSS.n36 585
R534 VSS.n36 VSS.n35 585
R535 VSS.n388 VSS.n387 585
R536 VSS.n387 VSS.n386 585
R537 VSS.n38 VSS.n37 585
R538 VSS.n385 VSS.n38 585
R539 VSS.n383 VSS.n382 585
R540 VSS.n384 VSS.n383 585
R541 VSS.n381 VSS.n40 585
R542 VSS.n40 VSS.n39 585
R543 VSS.n380 VSS.n379 585
R544 VSS.n379 VSS.n378 585
R545 VSS.n42 VSS.n41 585
R546 VSS.n377 VSS.n42 585
R547 VSS.n375 VSS.n374 585
R548 VSS.n376 VSS.n375 585
R549 VSS.n373 VSS.n44 585
R550 VSS.n44 VSS.n43 585
R551 VSS.n372 VSS.n371 585
R552 VSS.n371 VSS.n370 585
R553 VSS.n46 VSS.n45 585
R554 VSS.n369 VSS.n46 585
R555 VSS.n367 VSS.n366 585
R556 VSS.n368 VSS.n367 585
R557 VSS.n365 VSS.n48 585
R558 VSS.n48 VSS.n47 585
R559 VSS.n364 VSS.n363 585
R560 VSS.n363 VSS.n362 585
R561 VSS.n50 VSS.n49 585
R562 VSS.n361 VSS.n50 585
R563 VSS.n359 VSS.n358 585
R564 VSS.n360 VSS.n359 585
R565 VSS.n357 VSS.n52 585
R566 VSS.n52 VSS.n51 585
R567 VSS.n356 VSS.n355 585
R568 VSS.n355 VSS.n354 585
R569 VSS.n54 VSS.n53 585
R570 VSS.n353 VSS.n54 585
R571 VSS.n351 VSS.n350 585
R572 VSS.n352 VSS.n351 585
R573 VSS.n268 VSS.n267 585
R574 VSS.n100 VSS.n99 585
R575 VSS.n264 VSS.n263 585
R576 VSS.n265 VSS.n264 585
R577 VSS.n262 VSS.n111 585
R578 VSS.n261 VSS.n260 585
R579 VSS.n259 VSS.n258 585
R580 VSS.n257 VSS.n256 585
R581 VSS.n255 VSS.n254 585
R582 VSS.n253 VSS.n252 585
R583 VSS.n251 VSS.n250 585
R584 VSS.n249 VSS.n248 585
R585 VSS.n247 VSS.n246 585
R586 VSS.n245 VSS.n244 585
R587 VSS.n243 VSS.n242 585
R588 VSS.n241 VSS.n240 585
R589 VSS.n239 VSS.n238 585
R590 VSS.n237 VSS.n236 585
R591 VSS.n235 VSS.n234 585
R592 VSS.n233 VSS.n232 585
R593 VSS.n231 VSS.n109 585
R594 VSS.n265 VSS.n109 585
R595 VSS.n435 VSS.n19 585
R596 VSS.n434 VSS.n433 585
R597 VSS.n23 VSS.n22 585
R598 VSS.n429 VSS.n428 585
R599 VSS.n427 VSS.n32 585
R600 VSS.n426 VSS.n425 585
R601 VSS.n424 VSS.n423 585
R602 VSS.n422 VSS.n421 585
R603 VSS.n420 VSS.n419 585
R604 VSS.n418 VSS.n417 585
R605 VSS.n416 VSS.n415 585
R606 VSS.n414 VSS.n413 585
R607 VSS.n412 VSS.n411 585
R608 VSS.n410 VSS.n409 585
R609 VSS.n408 VSS.n407 585
R610 VSS.n406 VSS.n405 585
R611 VSS.n404 VSS.n403 585
R612 VSS.n402 VSS.n401 585
R613 VSS.n400 VSS.n399 585
R614 VSS.n398 VSS.n397 585
R615 VSS.n438 VSS.n437 585
R616 VSS.n439 VSS.n438 585
R617 VSS.n20 VSS.n18 585
R618 VSS.n18 VSS.n10 585
R619 VSS.n175 VSS.n11 585
R620 VSS.n475 VSS.n11 585
R621 VSS.n176 VSS.n152 585
R622 VSS.n152 VSS.n150 585
R623 VSS.n178 VSS.n177 585
R624 VSS.n179 VSS.n178 585
R625 VSS.n153 VSS.n151 585
R626 VSS.n151 VSS.n149 585
R627 VSS.n169 VSS.n168 585
R628 VSS.n168 VSS.n167 585
R629 VSS.n157 VSS.n156 585
R630 VSS.n166 VSS.n157 585
R631 VSS.n135 VSS.n134 585
R632 VSS.n138 VSS.n135 585
R633 VSS.n194 VSS.n193 585
R634 VSS.n193 VSS.n192 585
R635 VSS.n195 VSS.n130 585
R636 VSS.n136 VSS.n130 585
R637 VSS.n197 VSS.n196 585
R638 VSS.n198 VSS.n197 585
R639 VSS.n114 VSS.n113 585
R640 VSS.n120 VSS.n114 585
R641 VSS.n229 VSS.n228 585
R642 VSS.n228 VSS.n227 585
R643 VSS.n474 VSS.n473 585
R644 VSS.n475 VSS.n474 585
R645 VSS.n14 VSS.n12 585
R646 VSS.n150 VSS.n12 585
R647 VSS.n181 VSS.n180 585
R648 VSS.n180 VSS.n179 585
R649 VSS.n184 VSS.n148 585
R650 VSS.n149 VSS.n148 585
R651 VSS.n185 VSS.n147 585
R652 VSS.n167 VSS.n147 585
R653 VSS.n186 VSS.n146 585
R654 VSS.n166 VSS.n146 585
R655 VSS.n143 VSS.n140 585
R656 VSS.n140 VSS.n138 585
R657 VSS.n191 VSS.n190 585
R658 VSS.n192 VSS.n191 585
R659 VSS.n142 VSS.n139 585
R660 VSS.n139 VSS.n136 585
R661 VSS.n141 VSS.n123 585
R662 VSS.n198 VSS.n123 585
R663 VSS.n477 VSS.n476 585
R664 VSS.n476 VSS.n475 585
R665 VSS.n8 VSS.n6 585
R666 VSS.n150 VSS.n8 585
R667 VSS.n481 VSS.n5 585
R668 VSS.n179 VSS.n5 585
R669 VSS.n482 VSS.n4 585
R670 VSS.n149 VSS.n4 585
R671 VSS.n483 VSS.n3 585
R672 VSS.n167 VSS.n3 585
R673 VSS.n165 VSS.n2 585
R674 VSS.n166 VSS.n165 585
R675 VSS.n164 VSS.n163 585
R676 VSS.n164 VSS.n138 585
R677 VSS.n158 VSS.n137 585
R678 VSS.n192 VSS.n137 585
R679 VSS.n159 VSS.n128 585
R680 VSS.n136 VSS.n128 585
R681 VSS.n199 VSS.n129 585
R682 VSS.n199 VSS.n198 585
R683 VSS.n9 VSS.n7 585
R684 VSS.n451 VSS.n448 585
R685 VSS.n453 VSS.n452 585
R686 VSS.n455 VSS.n445 585
R687 VSS.n457 VSS.n456 585
R688 VSS.n459 VSS.n443 585
R689 VSS.n461 VSS.n460 585
R690 VSS.n462 VSS.n442 585
R691 VSS.n464 VSS.n463 585
R692 VSS.n466 VSS.n441 585
R693 VSS.n467 VSS.n16 585
R694 VSS.n470 VSS.n469 585
R695 VSS.n471 VSS.n13 585
R696 VSS.n440 VSS.n13 585
R697 VSS.n224 VSS.n223 585
R698 VSS.n222 VSS.n122 585
R699 VSS.n221 VSS.n121 585
R700 VSS.n226 VSS.n121 585
R701 VSS.n220 VSS.n219 585
R702 VSS.n218 VSS.n217 585
R703 VSS.n216 VSS.n215 585
R704 VSS.n214 VSS.n213 585
R705 VSS.n212 VSS.n211 585
R706 VSS.n210 VSS.n209 585
R707 VSS.n208 VSS.n207 585
R708 VSS.n205 VSS.n204 585
R709 VSS.n203 VSS.n202 585
R710 VSS.n201 VSS.n200 585
R711 VSS.n446 VSS.t5 510.822
R712 VSS.n125 VSS.t1 510.822
R713 VSS.n227 VSS.n110 450.832
R714 VSS.n439 VSS.n17 450.832
R715 VSS.n198 VSS.n120 292.748
R716 VSS.n192 VSS.n136 292.748
R717 VSS.n192 VSS.n138 292.748
R718 VSS.n167 VSS.n166 292.748
R719 VSS.n179 VSS.n149 292.748
R720 VSS.n179 VSS.n150 292.748
R721 VSS.n475 VSS.n10 292.748
R722 VSS.t9 VSS.n138 289.82
R723 VSS.t0 VSS.n149 289.82
R724 VSS.n226 VSS.n120 263.474
R725 VSS.n440 VSS.n10 263.474
R726 VSS.n266 VSS.n265 256.663
R727 VSS.n265 VSS.n101 256.663
R728 VSS.n265 VSS.n102 256.663
R729 VSS.n265 VSS.n103 256.663
R730 VSS.n265 VSS.n104 256.663
R731 VSS.n265 VSS.n105 256.663
R732 VSS.n265 VSS.n106 256.663
R733 VSS.n265 VSS.n107 256.663
R734 VSS.n265 VSS.n108 256.663
R735 VSS.n432 VSS.n431 256.663
R736 VSS.n431 VSS.n430 256.663
R737 VSS.n431 VSS.n31 256.663
R738 VSS.n431 VSS.n30 256.663
R739 VSS.n431 VSS.n29 256.663
R740 VSS.n431 VSS.n28 256.663
R741 VSS.n431 VSS.n27 256.663
R742 VSS.n431 VSS.n26 256.663
R743 VSS.n431 VSS.n25 256.663
R744 VSS.n431 VSS.n24 256.663
R745 VSS.n450 VSS.n440 256.663
R746 VSS.n449 VSS.n440 256.663
R747 VSS.n458 VSS.n440 256.663
R748 VSS.n444 VSS.n440 256.663
R749 VSS.n465 VSS.n440 256.663
R750 VSS.n468 VSS.n440 256.663
R751 VSS.n226 VSS.n225 256.663
R752 VSS.n226 VSS.n115 256.663
R753 VSS.n226 VSS.n116 256.663
R754 VSS.n226 VSS.n117 256.663
R755 VSS.n226 VSS.n118 256.663
R756 VSS.n226 VSS.n119 256.663
R757 VSS.n315 VSS.n73 240.244
R758 VSS.n321 VSS.n73 240.244
R759 VSS.n321 VSS.n71 240.244
R760 VSS.n325 VSS.n71 240.244
R761 VSS.n325 VSS.n67 240.244
R762 VSS.n331 VSS.n67 240.244
R763 VSS.n331 VSS.n65 240.244
R764 VSS.n335 VSS.n65 240.244
R765 VSS.n335 VSS.n61 240.244
R766 VSS.n342 VSS.n61 240.244
R767 VSS.n342 VSS.n59 240.244
R768 VSS.n346 VSS.n59 240.244
R769 VSS.n346 VSS.n56 240.244
R770 VSS.n228 VSS.n114 240.244
R771 VSS.n197 VSS.n114 240.244
R772 VSS.n197 VSS.n130 240.244
R773 VSS.n193 VSS.n130 240.244
R774 VSS.n193 VSS.n135 240.244
R775 VSS.n157 VSS.n135 240.244
R776 VSS.n168 VSS.n157 240.244
R777 VSS.n168 VSS.n151 240.244
R778 VSS.n178 VSS.n151 240.244
R779 VSS.n178 VSS.n152 240.244
R780 VSS.n152 VSS.n11 240.244
R781 VSS.n18 VSS.n11 240.244
R782 VSS.n438 VSS.n18 240.244
R783 VSS.n139 VSS.n123 240.244
R784 VSS.n191 VSS.n139 240.244
R785 VSS.n191 VSS.n140 240.244
R786 VSS.n146 VSS.n140 240.244
R787 VSS.n147 VSS.n146 240.244
R788 VSS.n148 VSS.n147 240.244
R789 VSS.n180 VSS.n148 240.244
R790 VSS.n180 VSS.n12 240.244
R791 VSS.n474 VSS.n12 240.244
R792 VSS.n199 VSS.n128 240.244
R793 VSS.n137 VSS.n128 240.244
R794 VSS.n164 VSS.n137 240.244
R795 VSS.n165 VSS.n164 240.244
R796 VSS.n165 VSS.n3 240.244
R797 VSS.n4 VSS.n3 240.244
R798 VSS.n5 VSS.n4 240.244
R799 VSS.n8 VSS.n5 240.244
R800 VSS.n476 VSS.n8 240.244
R801 VSS.n198 VSS.t2 231.272
R802 VSS.n475 VSS.t6 231.272
R803 VSS.n351 VSS.n54 163.367
R804 VSS.n355 VSS.n54 163.367
R805 VSS.n355 VSS.n52 163.367
R806 VSS.n359 VSS.n52 163.367
R807 VSS.n359 VSS.n50 163.367
R808 VSS.n363 VSS.n50 163.367
R809 VSS.n363 VSS.n48 163.367
R810 VSS.n367 VSS.n48 163.367
R811 VSS.n367 VSS.n46 163.367
R812 VSS.n371 VSS.n46 163.367
R813 VSS.n371 VSS.n44 163.367
R814 VSS.n375 VSS.n44 163.367
R815 VSS.n375 VSS.n42 163.367
R816 VSS.n379 VSS.n42 163.367
R817 VSS.n379 VSS.n40 163.367
R818 VSS.n383 VSS.n40 163.367
R819 VSS.n383 VSS.n38 163.367
R820 VSS.n387 VSS.n38 163.367
R821 VSS.n387 VSS.n36 163.367
R822 VSS.n392 VSS.n36 163.367
R823 VSS.n392 VSS.n34 163.367
R824 VSS.n396 VSS.n34 163.367
R825 VSS.n397 VSS.n396 163.367
R826 VSS.n401 VSS.n400 163.367
R827 VSS.n405 VSS.n404 163.367
R828 VSS.n409 VSS.n408 163.367
R829 VSS.n413 VSS.n412 163.367
R830 VSS.n417 VSS.n416 163.367
R831 VSS.n421 VSS.n420 163.367
R832 VSS.n425 VSS.n424 163.367
R833 VSS.n429 VSS.n32 163.367
R834 VSS.n433 VSS.n23 163.367
R835 VSS.n311 VSS.n76 163.367
R836 VSS.n311 VSS.n78 163.367
R837 VSS.n307 VSS.n78 163.367
R838 VSS.n307 VSS.n80 163.367
R839 VSS.n303 VSS.n80 163.367
R840 VSS.n303 VSS.n82 163.367
R841 VSS.n299 VSS.n82 163.367
R842 VSS.n299 VSS.n84 163.367
R843 VSS.n295 VSS.n84 163.367
R844 VSS.n295 VSS.n86 163.367
R845 VSS.n291 VSS.n86 163.367
R846 VSS.n291 VSS.n88 163.367
R847 VSS.n287 VSS.n88 163.367
R848 VSS.n287 VSS.n90 163.367
R849 VSS.n283 VSS.n90 163.367
R850 VSS.n283 VSS.n92 163.367
R851 VSS.n279 VSS.n92 163.367
R852 VSS.n279 VSS.n94 163.367
R853 VSS.n275 VSS.n94 163.367
R854 VSS.n275 VSS.n96 163.367
R855 VSS.n271 VSS.n96 163.367
R856 VSS.n271 VSS.n98 163.367
R857 VSS.n267 VSS.n98 163.367
R858 VSS.n264 VSS.n100 163.367
R859 VSS.n264 VSS.n111 163.367
R860 VSS.n260 VSS.n259 163.367
R861 VSS.n256 VSS.n255 163.367
R862 VSS.n252 VSS.n251 163.367
R863 VSS.n248 VSS.n247 163.367
R864 VSS.n244 VSS.n243 163.367
R865 VSS.n240 VSS.n239 163.367
R866 VSS.n236 VSS.n235 163.367
R867 VSS.n232 VSS.n109 163.367
R868 VSS.n122 VSS.n121 163.367
R869 VSS.n219 VSS.n121 163.367
R870 VSS.n217 VSS.n216 163.367
R871 VSS.n213 VSS.n212 163.367
R872 VSS.n209 VSS.n208 163.367
R873 VSS.n204 VSS.n203 163.367
R874 VSS.n469 VSS.n13 163.367
R875 VSS.n467 VSS.n466 163.367
R876 VSS.n464 VSS.n442 163.367
R877 VSS.n460 VSS.n459 163.367
R878 VSS.n457 VSS.n445 163.367
R879 VSS.n452 VSS.n451 163.367
R880 VSS.n446 VSS.t7 132.91
R881 VSS.n125 VSS.t4 132.91
R882 VSS.n447 VSS.t8 123.019
R883 VSS.n126 VSS.t3 123.019
R884 VSS.n400 VSS.n24 71.676
R885 VSS.n404 VSS.n25 71.676
R886 VSS.n408 VSS.n26 71.676
R887 VSS.n412 VSS.n27 71.676
R888 VSS.n416 VSS.n28 71.676
R889 VSS.n420 VSS.n29 71.676
R890 VSS.n424 VSS.n30 71.676
R891 VSS.n32 VSS.n31 71.676
R892 VSS.n430 VSS.n23 71.676
R893 VSS.n432 VSS.n19 71.676
R894 VSS.n267 VSS.n266 71.676
R895 VSS.n111 VSS.n101 71.676
R896 VSS.n259 VSS.n102 71.676
R897 VSS.n255 VSS.n103 71.676
R898 VSS.n251 VSS.n104 71.676
R899 VSS.n247 VSS.n105 71.676
R900 VSS.n243 VSS.n106 71.676
R901 VSS.n239 VSS.n107 71.676
R902 VSS.n235 VSS.n108 71.676
R903 VSS.n266 VSS.n100 71.676
R904 VSS.n260 VSS.n101 71.676
R905 VSS.n256 VSS.n102 71.676
R906 VSS.n252 VSS.n103 71.676
R907 VSS.n248 VSS.n104 71.676
R908 VSS.n244 VSS.n105 71.676
R909 VSS.n240 VSS.n106 71.676
R910 VSS.n236 VSS.n107 71.676
R911 VSS.n232 VSS.n108 71.676
R912 VSS.n433 VSS.n432 71.676
R913 VSS.n430 VSS.n429 71.676
R914 VSS.n425 VSS.n31 71.676
R915 VSS.n421 VSS.n30 71.676
R916 VSS.n417 VSS.n29 71.676
R917 VSS.n413 VSS.n28 71.676
R918 VSS.n409 VSS.n27 71.676
R919 VSS.n405 VSS.n26 71.676
R920 VSS.n401 VSS.n25 71.676
R921 VSS.n397 VSS.n24 71.676
R922 VSS.n225 VSS.n224 71.676
R923 VSS.n219 VSS.n115 71.676
R924 VSS.n216 VSS.n116 71.676
R925 VSS.n212 VSS.n117 71.676
R926 VSS.n208 VSS.n118 71.676
R927 VSS.n203 VSS.n119 71.676
R928 VSS.n468 VSS.n467 71.676
R929 VSS.n465 VSS.n464 71.676
R930 VSS.n460 VSS.n444 71.676
R931 VSS.n458 VSS.n457 71.676
R932 VSS.n452 VSS.n449 71.676
R933 VSS.n450 VSS.n9 71.676
R934 VSS.n451 VSS.n450 71.676
R935 VSS.n449 VSS.n445 71.676
R936 VSS.n459 VSS.n458 71.676
R937 VSS.n444 VSS.n442 71.676
R938 VSS.n466 VSS.n465 71.676
R939 VSS.n469 VSS.n468 71.676
R940 VSS.n225 VSS.n122 71.676
R941 VSS.n217 VSS.n115 71.676
R942 VSS.n213 VSS.n116 71.676
R943 VSS.n209 VSS.n117 71.676
R944 VSS.n204 VSS.n118 71.676
R945 VSS.n200 VSS.n119 71.676
R946 VSS.n136 VSS.t2 61.4775
R947 VSS.n150 VSS.t6 61.4775
R948 VSS.n265 VSS.n110 58.5501
R949 VSS.n431 VSS.n17 58.5501
R950 VSS.n454 VSS.n447 34.3278
R951 VSS.n206 VSS.n126 34.3278
R952 VSS.n350 VSS.n349 31.7316
R953 VSS.n436 VSS.n435 31.7316
R954 VSS.n317 VSS.n75 31.7316
R955 VSS.n231 VSS.n230 31.7316
R956 VSS.n227 VSS.n226 29.2753
R957 VSS.n440 VSS.n439 29.2753
R958 VSS.n472 VSS.n471 29.2584
R959 VSS.n478 VSS.n7 29.2584
R960 VSS.n223 VSS.n124 29.2584
R961 VSS.n201 VSS.n127 29.2584
R962 VSS.n316 VSS.n74 19.3944
R963 VSS.n320 VSS.n74 19.3944
R964 VSS.n320 VSS.n70 19.3944
R965 VSS.n326 VSS.n70 19.3944
R966 VSS.n326 VSS.n68 19.3944
R967 VSS.n330 VSS.n68 19.3944
R968 VSS.n330 VSS.n64 19.3944
R969 VSS.n336 VSS.n64 19.3944
R970 VSS.n336 VSS.n62 19.3944
R971 VSS.n341 VSS.n62 19.3944
R972 VSS.n341 VSS.n58 19.3944
R973 VSS.n347 VSS.n58 19.3944
R974 VSS.n348 VSS.n347 19.3944
R975 VSS.n229 VSS.n113 19.3944
R976 VSS.n196 VSS.n113 19.3944
R977 VSS.n196 VSS.n195 19.3944
R978 VSS.n195 VSS.n194 19.3944
R979 VSS.n194 VSS.n134 19.3944
R980 VSS.n156 VSS.n134 19.3944
R981 VSS.n169 VSS.n156 19.3944
R982 VSS.n169 VSS.n153 19.3944
R983 VSS.n177 VSS.n153 19.3944
R984 VSS.n177 VSS.n176 19.3944
R985 VSS.n176 VSS.n175 19.3944
R986 VSS.n175 VSS.n20 19.3944
R987 VSS.n437 VSS.n20 19.3944
R988 VSS.n142 VSS.n141 19.3944
R989 VSS.n190 VSS.n142 19.3944
R990 VSS.n190 VSS.n143 19.3944
R991 VSS.n186 VSS.n143 19.3944
R992 VSS.n186 VSS.n185 19.3944
R993 VSS.n185 VSS.n184 19.3944
R994 VSS.n184 VSS.n181 19.3944
R995 VSS.n181 VSS.n14 19.3944
R996 VSS.n473 VSS.n14 19.3944
R997 VSS.n159 VSS.n129 19.3944
R998 VSS.n159 VSS.n158 19.3944
R999 VSS.n163 VSS.n158 19.3944
R1000 VSS.n163 VSS.n2 19.3944
R1001 VSS.n483 VSS.n2 19.3944
R1002 VSS.n483 VSS.n482 19.3944
R1003 VSS.n482 VSS.n481 19.3944
R1004 VSS.n481 VSS.n6 19.3944
R1005 VSS.n477 VSS.n6 19.3944
R1006 VSS.n350 VSS.n53 10.6151
R1007 VSS.n356 VSS.n53 10.6151
R1008 VSS.n357 VSS.n356 10.6151
R1009 VSS.n358 VSS.n357 10.6151
R1010 VSS.n358 VSS.n49 10.6151
R1011 VSS.n364 VSS.n49 10.6151
R1012 VSS.n365 VSS.n364 10.6151
R1013 VSS.n366 VSS.n365 10.6151
R1014 VSS.n366 VSS.n45 10.6151
R1015 VSS.n372 VSS.n45 10.6151
R1016 VSS.n373 VSS.n372 10.6151
R1017 VSS.n374 VSS.n373 10.6151
R1018 VSS.n374 VSS.n41 10.6151
R1019 VSS.n380 VSS.n41 10.6151
R1020 VSS.n381 VSS.n380 10.6151
R1021 VSS.n382 VSS.n381 10.6151
R1022 VSS.n382 VSS.n37 10.6151
R1023 VSS.n388 VSS.n37 10.6151
R1024 VSS.n389 VSS.n388 10.6151
R1025 VSS.n391 VSS.n389 10.6151
R1026 VSS.n391 VSS.n390 10.6151
R1027 VSS.n390 VSS.n33 10.6151
R1028 VSS.n398 VSS.n33 10.6151
R1029 VSS.n399 VSS.n398 10.6151
R1030 VSS.n402 VSS.n399 10.6151
R1031 VSS.n403 VSS.n402 10.6151
R1032 VSS.n406 VSS.n403 10.6151
R1033 VSS.n407 VSS.n406 10.6151
R1034 VSS.n410 VSS.n407 10.6151
R1035 VSS.n411 VSS.n410 10.6151
R1036 VSS.n414 VSS.n411 10.6151
R1037 VSS.n415 VSS.n414 10.6151
R1038 VSS.n418 VSS.n415 10.6151
R1039 VSS.n419 VSS.n418 10.6151
R1040 VSS.n422 VSS.n419 10.6151
R1041 VSS.n423 VSS.n422 10.6151
R1042 VSS.n426 VSS.n423 10.6151
R1043 VSS.n427 VSS.n426 10.6151
R1044 VSS.n428 VSS.n427 10.6151
R1045 VSS.n428 VSS.n22 10.6151
R1046 VSS.n434 VSS.n22 10.6151
R1047 VSS.n435 VSS.n434 10.6151
R1048 VSS.n310 VSS.n75 10.6151
R1049 VSS.n310 VSS.n309 10.6151
R1050 VSS.n309 VSS.n308 10.6151
R1051 VSS.n308 VSS.n79 10.6151
R1052 VSS.n302 VSS.n79 10.6151
R1053 VSS.n302 VSS.n301 10.6151
R1054 VSS.n301 VSS.n300 10.6151
R1055 VSS.n300 VSS.n83 10.6151
R1056 VSS.n294 VSS.n83 10.6151
R1057 VSS.n294 VSS.n293 10.6151
R1058 VSS.n293 VSS.n292 10.6151
R1059 VSS.n292 VSS.n87 10.6151
R1060 VSS.n286 VSS.n87 10.6151
R1061 VSS.n286 VSS.n285 10.6151
R1062 VSS.n285 VSS.n284 10.6151
R1063 VSS.n284 VSS.n91 10.6151
R1064 VSS.n278 VSS.n91 10.6151
R1065 VSS.n278 VSS.n277 10.6151
R1066 VSS.n277 VSS.n276 10.6151
R1067 VSS.n276 VSS.n95 10.6151
R1068 VSS.n270 VSS.n95 10.6151
R1069 VSS.n270 VSS.n269 10.6151
R1070 VSS.n269 VSS.n268 10.6151
R1071 VSS.n268 VSS.n99 10.6151
R1072 VSS.n263 VSS.n99 10.6151
R1073 VSS.n263 VSS.n262 10.6151
R1074 VSS.n262 VSS.n261 10.6151
R1075 VSS.n261 VSS.n258 10.6151
R1076 VSS.n258 VSS.n257 10.6151
R1077 VSS.n257 VSS.n254 10.6151
R1078 VSS.n254 VSS.n253 10.6151
R1079 VSS.n253 VSS.n250 10.6151
R1080 VSS.n250 VSS.n249 10.6151
R1081 VSS.n249 VSS.n246 10.6151
R1082 VSS.n246 VSS.n245 10.6151
R1083 VSS.n245 VSS.n242 10.6151
R1084 VSS.n242 VSS.n241 10.6151
R1085 VSS.n241 VSS.n238 10.6151
R1086 VSS.n238 VSS.n237 10.6151
R1087 VSS.n237 VSS.n234 10.6151
R1088 VSS.n234 VSS.n233 10.6151
R1089 VSS.n233 VSS.n231 10.6151
R1090 VSS.n471 VSS.n470 10.6151
R1091 VSS.n470 VSS.n16 10.6151
R1092 VSS.n441 VSS.n16 10.6151
R1093 VSS.n463 VSS.n441 10.6151
R1094 VSS.n463 VSS.n462 10.6151
R1095 VSS.n462 VSS.n461 10.6151
R1096 VSS.n461 VSS.n443 10.6151
R1097 VSS.n456 VSS.n443 10.6151
R1098 VSS.n456 VSS.n455 10.6151
R1099 VSS.n453 VSS.n448 10.6151
R1100 VSS.n448 VSS.n7 10.6151
R1101 VSS.n223 VSS.n222 10.6151
R1102 VSS.n222 VSS.n221 10.6151
R1103 VSS.n221 VSS.n220 10.6151
R1104 VSS.n220 VSS.n218 10.6151
R1105 VSS.n218 VSS.n215 10.6151
R1106 VSS.n215 VSS.n214 10.6151
R1107 VSS.n214 VSS.n211 10.6151
R1108 VSS.n211 VSS.n210 10.6151
R1109 VSS.n210 VSS.n207 10.6151
R1110 VSS.n205 VSS.n202 10.6151
R1111 VSS.n202 VSS.n201 10.6151
R1112 VSS.n455 VSS.n454 10.1468
R1113 VSS.n207 VSS.n206 10.1468
R1114 VSS.n447 VSS.n446 9.89141
R1115 VSS.n126 VSS.n125 9.89141
R1116 VSS.n113 VSS.n112 9.3005
R1117 VSS.n196 VSS.n131 9.3005
R1118 VSS.n195 VSS.n132 9.3005
R1119 VSS.n194 VSS.n133 9.3005
R1120 VSS.n154 VSS.n134 9.3005
R1121 VSS.n156 VSS.n155 9.3005
R1122 VSS.n170 VSS.n169 9.3005
R1123 VSS.n171 VSS.n153 9.3005
R1124 VSS.n177 VSS.n172 9.3005
R1125 VSS.n176 VSS.n173 9.3005
R1126 VSS.n175 VSS.n174 9.3005
R1127 VSS.n21 VSS.n20 9.3005
R1128 VSS.n437 VSS.n436 9.3005
R1129 VSS.n230 VSS.n229 9.3005
R1130 VSS.n317 VSS.n316 9.3005
R1131 VSS.n318 VSS.n74 9.3005
R1132 VSS.n320 VSS.n319 9.3005
R1133 VSS.n70 VSS.n69 9.3005
R1134 VSS.n327 VSS.n326 9.3005
R1135 VSS.n328 VSS.n68 9.3005
R1136 VSS.n330 VSS.n329 9.3005
R1137 VSS.n64 VSS.n63 9.3005
R1138 VSS.n337 VSS.n336 9.3005
R1139 VSS.n338 VSS.n62 9.3005
R1140 VSS.n341 VSS.n340 9.3005
R1141 VSS.n339 VSS.n58 9.3005
R1142 VSS.n347 VSS.n57 9.3005
R1143 VSS.n349 VSS.n348 9.3005
R1144 VSS.n482 VSS.n0 9.3005
R1145 VSS.n481 VSS.n480 9.3005
R1146 VSS.n479 VSS.n6 9.3005
R1147 VSS.n478 VSS.n477 9.3005
R1148 VSS.n144 VSS.n142 9.3005
R1149 VSS.n190 VSS.n189 9.3005
R1150 VSS.n188 VSS.n143 9.3005
R1151 VSS.n187 VSS.n186 9.3005
R1152 VSS.n185 VSS.n145 9.3005
R1153 VSS.n184 VSS.n183 9.3005
R1154 VSS.n182 VSS.n181 9.3005
R1155 VSS.n15 VSS.n14 9.3005
R1156 VSS.n473 VSS.n472 9.3005
R1157 VSS.n141 VSS.n124 9.3005
R1158 VSS.n160 VSS.n159 9.3005
R1159 VSS.n161 VSS.n158 9.3005
R1160 VSS.n163 VSS.n162 9.3005
R1161 VSS.n2 VSS.n1 9.3005
R1162 VSS.n129 VSS.n127 9.3005
R1163 VSS VSS.n483 9.3005
R1164 VSS.n166 VSS.t9 2.92798
R1165 VSS.n167 VSS.t0 2.92798
R1166 VSS.n454 VSS.n453 0.468793
R1167 VSS.n206 VSS.n205 0.468793
R1168 VSS.n230 VSS.n112 0.152939
R1169 VSS.n131 VSS.n112 0.152939
R1170 VSS.n132 VSS.n131 0.152939
R1171 VSS.n133 VSS.n132 0.152939
R1172 VSS.n154 VSS.n133 0.152939
R1173 VSS.n155 VSS.n154 0.152939
R1174 VSS.n170 VSS.n155 0.152939
R1175 VSS.n171 VSS.n170 0.152939
R1176 VSS.n172 VSS.n171 0.152939
R1177 VSS.n173 VSS.n172 0.152939
R1178 VSS.n174 VSS.n173 0.152939
R1179 VSS.n174 VSS.n21 0.152939
R1180 VSS.n436 VSS.n21 0.152939
R1181 VSS.n318 VSS.n317 0.152939
R1182 VSS.n319 VSS.n318 0.152939
R1183 VSS.n319 VSS.n69 0.152939
R1184 VSS.n327 VSS.n69 0.152939
R1185 VSS.n328 VSS.n327 0.152939
R1186 VSS.n329 VSS.n328 0.152939
R1187 VSS.n329 VSS.n63 0.152939
R1188 VSS.n337 VSS.n63 0.152939
R1189 VSS.n338 VSS.n337 0.152939
R1190 VSS.n340 VSS.n338 0.152939
R1191 VSS.n340 VSS.n339 0.152939
R1192 VSS.n339 VSS.n57 0.152939
R1193 VSS.n349 VSS.n57 0.152939
R1194 VSS VSS.n0 0.152939
R1195 VSS.n480 VSS.n0 0.152939
R1196 VSS.n480 VSS.n479 0.152939
R1197 VSS.n479 VSS.n478 0.152939
R1198 VSS.n144 VSS.n124 0.152939
R1199 VSS.n189 VSS.n144 0.152939
R1200 VSS.n189 VSS.n188 0.152939
R1201 VSS.n188 VSS.n187 0.152939
R1202 VSS.n187 VSS.n145 0.152939
R1203 VSS.n183 VSS.n145 0.152939
R1204 VSS.n183 VSS.n182 0.152939
R1205 VSS.n182 VSS.n15 0.152939
R1206 VSS.n472 VSS.n15 0.152939
R1207 VSS.n160 VSS.n127 0.152939
R1208 VSS.n161 VSS.n160 0.152939
R1209 VSS.n162 VSS.n161 0.152939
R1210 VSS.n162 VSS.n1 0.152939
R1211 VSS VSS.n1 0.1255
R1212 VGN.n0 VGN.t1 479.079
R1213 VGN.n0 VGN.t0 479.079
R1214 VGN VGN.n0 161.381
C0 VOUT VGN 0.101313f
C1 VOUT VIN 2.7367f
C2 VCC VOUT 0.45657f
C3 VOUT VGP 0.163715f
C4 VGN VIN 0.101199f
C5 VCC VGN 0.001688f
C6 VCC VIN 0.936093f
C7 VGN VGP 0.00144f
C8 VGP VIN 0.163012f
C9 VCC VGP 0.446573f
C10 VGN VSS 0.492795f
C11 VOUT VSS 1.976219f
C12 VIN VSS 1.195349f
C13 VGP VSS 0.06621f
C14 VCC VSS 8.669099f
C15 VOUT.t0 VSS 0.101912f
C16 VOUT.t1 VSS 0.101912f
C17 VOUT.n0 VSS 0.597439f
C18 VOUT.t3 VSS 0.050956f
C19 VOUT.t2 VSS 0.050956f
C20 VOUT.n1 VSS 0.381558f
C21 VIN.n0 VSS 0.020271f
C22 VIN.n1 VSS 0.018236f
C23 VIN.n2 VSS 0.009799f
C24 VIN.n3 VSS 0.023162f
C25 VIN.n4 VSS 0.010376f
C26 VIN.n5 VSS 0.071238f
C27 VIN.t1 VSS 0.051491f
C28 VIN.n6 VSS 0.017372f
C29 VIN.n7 VSS 0.014569f
C30 VIN.n8 VSS 0.009799f
C31 VIN.n9 VSS 0.249664f
C32 VIN.n10 VSS 0.018236f
C33 VIN.n11 VSS 0.009799f
C34 VIN.n12 VSS 0.010376f
C35 VIN.n13 VSS 0.023162f
C36 VIN.n14 VSS 0.056867f
C37 VIN.n15 VSS 0.010376f
C38 VIN.n16 VSS 0.009799f
C39 VIN.n17 VSS 0.046138f
C40 VIN.n18 VSS 0.029378f
C41 VIN.n19 VSS 0.020271f
C42 VIN.n20 VSS 0.018236f
C43 VIN.n21 VSS 0.009799f
C44 VIN.n22 VSS 0.023162f
C45 VIN.n23 VSS 0.010376f
C46 VIN.n24 VSS 0.071238f
C47 VIN.t0 VSS 0.051491f
C48 VIN.n25 VSS 0.017372f
C49 VIN.n26 VSS 0.014569f
C50 VIN.n27 VSS 0.009799f
C51 VIN.n28 VSS 0.249664f
C52 VIN.n29 VSS 0.018236f
C53 VIN.n30 VSS 0.009799f
C54 VIN.n31 VSS 0.010376f
C55 VIN.n32 VSS 0.023162f
C56 VIN.n33 VSS 0.056867f
C57 VIN.n34 VSS 0.010376f
C58 VIN.n35 VSS 0.009799f
C59 VIN.n36 VSS 0.046138f
C60 VIN.n37 VSS 0.028751f
C61 VIN.n38 VSS 0.283185f
C62 VIN.n39 VSS 0.026617f
C63 VIN.n40 VSS 0.058893f
C64 VIN.t2 VSS 0.044196f
C65 VIN.n41 VSS 0.046092f
C66 VIN.n42 VSS 0.014858f
C67 VIN.n43 VSS 0.009799f
C68 VIN.n44 VSS 0.129815f
C69 VIN.n45 VSS 0.029844f
C70 VIN.n46 VSS 0.026617f
C71 VIN.n47 VSS 0.058893f
C72 VIN.t3 VSS 0.044196f
C73 VIN.n48 VSS 0.046092f
C74 VIN.n49 VSS 0.014858f
C75 VIN.n50 VSS 0.009799f
C76 VIN.n51 VSS 0.129815f
C77 VIN.n52 VSS 0.029178f
C78 VIN.n53 VSS 0.088629f
.ends

