* NGSPICE file created from diff_pair_sample_1487.ext - technology: sky130A

.subckt diff_pair_sample_1487 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t0 w_n2050_n2038# sky130_fd_pr__pfet_01v8 ad=0.88275 pd=5.68 as=0.88275 ps=5.68 w=5.35 l=1.02
X1 VDD2.t5 VN.t0 VTAIL.t1 w_n2050_n2038# sky130_fd_pr__pfet_01v8 ad=0.88275 pd=5.68 as=2.0865 ps=11.48 w=5.35 l=1.02
X2 VDD1.t5 VP.t1 VTAIL.t10 w_n2050_n2038# sky130_fd_pr__pfet_01v8 ad=2.0865 pd=11.48 as=0.88275 ps=5.68 w=5.35 l=1.02
X3 B.t11 B.t9 B.t10 w_n2050_n2038# sky130_fd_pr__pfet_01v8 ad=2.0865 pd=11.48 as=0 ps=0 w=5.35 l=1.02
X4 VTAIL.t9 VP.t2 VDD1.t3 w_n2050_n2038# sky130_fd_pr__pfet_01v8 ad=0.88275 pd=5.68 as=0.88275 ps=5.68 w=5.35 l=1.02
X5 VTAIL.t0 VN.t1 VDD2.t4 w_n2050_n2038# sky130_fd_pr__pfet_01v8 ad=0.88275 pd=5.68 as=0.88275 ps=5.68 w=5.35 l=1.02
X6 B.t8 B.t6 B.t7 w_n2050_n2038# sky130_fd_pr__pfet_01v8 ad=2.0865 pd=11.48 as=0 ps=0 w=5.35 l=1.02
X7 B.t5 B.t3 B.t4 w_n2050_n2038# sky130_fd_pr__pfet_01v8 ad=2.0865 pd=11.48 as=0 ps=0 w=5.35 l=1.02
X8 B.t2 B.t0 B.t1 w_n2050_n2038# sky130_fd_pr__pfet_01v8 ad=2.0865 pd=11.48 as=0 ps=0 w=5.35 l=1.02
X9 VDD2.t3 VN.t2 VTAIL.t2 w_n2050_n2038# sky130_fd_pr__pfet_01v8 ad=0.88275 pd=5.68 as=2.0865 ps=11.48 w=5.35 l=1.02
X10 VDD1.t1 VP.t3 VTAIL.t8 w_n2050_n2038# sky130_fd_pr__pfet_01v8 ad=2.0865 pd=11.48 as=0.88275 ps=5.68 w=5.35 l=1.02
X11 VDD2.t2 VN.t3 VTAIL.t4 w_n2050_n2038# sky130_fd_pr__pfet_01v8 ad=2.0865 pd=11.48 as=0.88275 ps=5.68 w=5.35 l=1.02
X12 VDD1.t4 VP.t4 VTAIL.t7 w_n2050_n2038# sky130_fd_pr__pfet_01v8 ad=0.88275 pd=5.68 as=2.0865 ps=11.48 w=5.35 l=1.02
X13 VDD1.t2 VP.t5 VTAIL.t6 w_n2050_n2038# sky130_fd_pr__pfet_01v8 ad=0.88275 pd=5.68 as=2.0865 ps=11.48 w=5.35 l=1.02
X14 VDD2.t1 VN.t4 VTAIL.t5 w_n2050_n2038# sky130_fd_pr__pfet_01v8 ad=2.0865 pd=11.48 as=0.88275 ps=5.68 w=5.35 l=1.02
X15 VTAIL.t3 VN.t5 VDD2.t0 w_n2050_n2038# sky130_fd_pr__pfet_01v8 ad=0.88275 pd=5.68 as=0.88275 ps=5.68 w=5.35 l=1.02
R0 VP.n3 VP.t3 187.69
R1 VP.n8 VP.t1 165.156
R2 VP.n14 VP.t4 165.156
R3 VP.n6 VP.t5 165.156
R4 VP.n5 VP.n2 161.3
R5 VP.n13 VP.n0 161.3
R6 VP.n12 VP.n11 161.3
R7 VP.n10 VP.n1 161.3
R8 VP.n12 VP.t0 126.407
R9 VP.n4 VP.t2 126.407
R10 VP.n7 VP.n6 80.6037
R11 VP.n15 VP.n14 80.6037
R12 VP.n9 VP.n8 80.6037
R13 VP.n8 VP.n1 48.6898
R14 VP.n14 VP.n13 48.6898
R15 VP.n6 VP.n5 48.6898
R16 VP.n9 VP.n7 37.5506
R17 VP.n4 VP.n3 32.2015
R18 VP.n3 VP.n2 28.3725
R19 VP.n12 VP.n1 24.4675
R20 VP.n13 VP.n12 24.4675
R21 VP.n5 VP.n4 24.4675
R22 VP.n7 VP.n2 0.285035
R23 VP.n10 VP.n9 0.285035
R24 VP.n15 VP.n0 0.285035
R25 VP.n11 VP.n10 0.189894
R26 VP.n11 VP.n0 0.189894
R27 VP VP.n15 0.146778
R28 VDD1.n22 VDD1.n0 756.745
R29 VDD1.n49 VDD1.n27 756.745
R30 VDD1.n23 VDD1.n22 585
R31 VDD1.n21 VDD1.n20 585
R32 VDD1.n4 VDD1.n3 585
R33 VDD1.n15 VDD1.n14 585
R34 VDD1.n13 VDD1.n12 585
R35 VDD1.n8 VDD1.n7 585
R36 VDD1.n35 VDD1.n34 585
R37 VDD1.n40 VDD1.n39 585
R38 VDD1.n42 VDD1.n41 585
R39 VDD1.n31 VDD1.n30 585
R40 VDD1.n48 VDD1.n47 585
R41 VDD1.n50 VDD1.n49 585
R42 VDD1.n9 VDD1.t1 327.856
R43 VDD1.n36 VDD1.t5 327.856
R44 VDD1.n22 VDD1.n21 171.744
R45 VDD1.n21 VDD1.n3 171.744
R46 VDD1.n14 VDD1.n3 171.744
R47 VDD1.n14 VDD1.n13 171.744
R48 VDD1.n13 VDD1.n7 171.744
R49 VDD1.n40 VDD1.n34 171.744
R50 VDD1.n41 VDD1.n40 171.744
R51 VDD1.n41 VDD1.n30 171.744
R52 VDD1.n48 VDD1.n30 171.744
R53 VDD1.n49 VDD1.n48 171.744
R54 VDD1.n55 VDD1.n54 98.9239
R55 VDD1.n57 VDD1.n56 98.6883
R56 VDD1.t1 VDD1.n7 85.8723
R57 VDD1.t5 VDD1.n34 85.8723
R58 VDD1 VDD1.n26 51.1527
R59 VDD1.n55 VDD1.n53 51.0392
R60 VDD1.n57 VDD1.n55 33.2746
R61 VDD1.n9 VDD1.n8 16.381
R62 VDD1.n36 VDD1.n35 16.381
R63 VDD1.n12 VDD1.n11 12.8005
R64 VDD1.n39 VDD1.n38 12.8005
R65 VDD1.n15 VDD1.n6 12.0247
R66 VDD1.n42 VDD1.n33 12.0247
R67 VDD1.n16 VDD1.n4 11.249
R68 VDD1.n43 VDD1.n31 11.249
R69 VDD1.n20 VDD1.n19 10.4732
R70 VDD1.n47 VDD1.n46 10.4732
R71 VDD1.n23 VDD1.n2 9.69747
R72 VDD1.n50 VDD1.n29 9.69747
R73 VDD1.n26 VDD1.n25 9.45567
R74 VDD1.n53 VDD1.n52 9.45567
R75 VDD1.n25 VDD1.n24 9.3005
R76 VDD1.n2 VDD1.n1 9.3005
R77 VDD1.n19 VDD1.n18 9.3005
R78 VDD1.n17 VDD1.n16 9.3005
R79 VDD1.n6 VDD1.n5 9.3005
R80 VDD1.n11 VDD1.n10 9.3005
R81 VDD1.n52 VDD1.n51 9.3005
R82 VDD1.n29 VDD1.n28 9.3005
R83 VDD1.n46 VDD1.n45 9.3005
R84 VDD1.n44 VDD1.n43 9.3005
R85 VDD1.n33 VDD1.n32 9.3005
R86 VDD1.n38 VDD1.n37 9.3005
R87 VDD1.n24 VDD1.n0 8.92171
R88 VDD1.n51 VDD1.n27 8.92171
R89 VDD1.n56 VDD1.t3 6.0762
R90 VDD1.n56 VDD1.t2 6.0762
R91 VDD1.n54 VDD1.t0 6.0762
R92 VDD1.n54 VDD1.t4 6.0762
R93 VDD1.n26 VDD1.n0 5.04292
R94 VDD1.n53 VDD1.n27 5.04292
R95 VDD1.n24 VDD1.n23 4.26717
R96 VDD1.n51 VDD1.n50 4.26717
R97 VDD1.n10 VDD1.n9 3.71853
R98 VDD1.n37 VDD1.n36 3.71853
R99 VDD1.n20 VDD1.n2 3.49141
R100 VDD1.n47 VDD1.n29 3.49141
R101 VDD1.n19 VDD1.n4 2.71565
R102 VDD1.n46 VDD1.n31 2.71565
R103 VDD1.n16 VDD1.n15 1.93989
R104 VDD1.n43 VDD1.n42 1.93989
R105 VDD1.n12 VDD1.n6 1.16414
R106 VDD1.n39 VDD1.n33 1.16414
R107 VDD1.n11 VDD1.n8 0.388379
R108 VDD1.n38 VDD1.n35 0.388379
R109 VDD1 VDD1.n57 0.233259
R110 VDD1.n25 VDD1.n1 0.155672
R111 VDD1.n18 VDD1.n1 0.155672
R112 VDD1.n18 VDD1.n17 0.155672
R113 VDD1.n17 VDD1.n5 0.155672
R114 VDD1.n10 VDD1.n5 0.155672
R115 VDD1.n37 VDD1.n32 0.155672
R116 VDD1.n44 VDD1.n32 0.155672
R117 VDD1.n45 VDD1.n44 0.155672
R118 VDD1.n45 VDD1.n28 0.155672
R119 VDD1.n52 VDD1.n28 0.155672
R120 VTAIL.n114 VTAIL.n92 756.745
R121 VTAIL.n24 VTAIL.n2 756.745
R122 VTAIL.n86 VTAIL.n64 756.745
R123 VTAIL.n56 VTAIL.n34 756.745
R124 VTAIL.n100 VTAIL.n99 585
R125 VTAIL.n105 VTAIL.n104 585
R126 VTAIL.n107 VTAIL.n106 585
R127 VTAIL.n96 VTAIL.n95 585
R128 VTAIL.n113 VTAIL.n112 585
R129 VTAIL.n115 VTAIL.n114 585
R130 VTAIL.n10 VTAIL.n9 585
R131 VTAIL.n15 VTAIL.n14 585
R132 VTAIL.n17 VTAIL.n16 585
R133 VTAIL.n6 VTAIL.n5 585
R134 VTAIL.n23 VTAIL.n22 585
R135 VTAIL.n25 VTAIL.n24 585
R136 VTAIL.n87 VTAIL.n86 585
R137 VTAIL.n85 VTAIL.n84 585
R138 VTAIL.n68 VTAIL.n67 585
R139 VTAIL.n79 VTAIL.n78 585
R140 VTAIL.n77 VTAIL.n76 585
R141 VTAIL.n72 VTAIL.n71 585
R142 VTAIL.n57 VTAIL.n56 585
R143 VTAIL.n55 VTAIL.n54 585
R144 VTAIL.n38 VTAIL.n37 585
R145 VTAIL.n49 VTAIL.n48 585
R146 VTAIL.n47 VTAIL.n46 585
R147 VTAIL.n42 VTAIL.n41 585
R148 VTAIL.n101 VTAIL.t1 327.856
R149 VTAIL.n11 VTAIL.t7 327.856
R150 VTAIL.n73 VTAIL.t6 327.856
R151 VTAIL.n43 VTAIL.t2 327.856
R152 VTAIL.n105 VTAIL.n99 171.744
R153 VTAIL.n106 VTAIL.n105 171.744
R154 VTAIL.n106 VTAIL.n95 171.744
R155 VTAIL.n113 VTAIL.n95 171.744
R156 VTAIL.n114 VTAIL.n113 171.744
R157 VTAIL.n15 VTAIL.n9 171.744
R158 VTAIL.n16 VTAIL.n15 171.744
R159 VTAIL.n16 VTAIL.n5 171.744
R160 VTAIL.n23 VTAIL.n5 171.744
R161 VTAIL.n24 VTAIL.n23 171.744
R162 VTAIL.n86 VTAIL.n85 171.744
R163 VTAIL.n85 VTAIL.n67 171.744
R164 VTAIL.n78 VTAIL.n67 171.744
R165 VTAIL.n78 VTAIL.n77 171.744
R166 VTAIL.n77 VTAIL.n71 171.744
R167 VTAIL.n56 VTAIL.n55 171.744
R168 VTAIL.n55 VTAIL.n37 171.744
R169 VTAIL.n48 VTAIL.n37 171.744
R170 VTAIL.n48 VTAIL.n47 171.744
R171 VTAIL.n47 VTAIL.n41 171.744
R172 VTAIL.t1 VTAIL.n99 85.8723
R173 VTAIL.t7 VTAIL.n9 85.8723
R174 VTAIL.t6 VTAIL.n71 85.8723
R175 VTAIL.t2 VTAIL.n41 85.8723
R176 VTAIL.n63 VTAIL.n62 82.0097
R177 VTAIL.n33 VTAIL.n32 82.0097
R178 VTAIL.n1 VTAIL.n0 82.0096
R179 VTAIL.n31 VTAIL.n30 82.0096
R180 VTAIL.n119 VTAIL.n118 33.5429
R181 VTAIL.n29 VTAIL.n28 33.5429
R182 VTAIL.n91 VTAIL.n90 33.5429
R183 VTAIL.n61 VTAIL.n60 33.5429
R184 VTAIL.n33 VTAIL.n31 19.3065
R185 VTAIL.n119 VTAIL.n91 18.1427
R186 VTAIL.n101 VTAIL.n100 16.381
R187 VTAIL.n11 VTAIL.n10 16.381
R188 VTAIL.n73 VTAIL.n72 16.381
R189 VTAIL.n43 VTAIL.n42 16.381
R190 VTAIL.n104 VTAIL.n103 12.8005
R191 VTAIL.n14 VTAIL.n13 12.8005
R192 VTAIL.n76 VTAIL.n75 12.8005
R193 VTAIL.n46 VTAIL.n45 12.8005
R194 VTAIL.n107 VTAIL.n98 12.0247
R195 VTAIL.n17 VTAIL.n8 12.0247
R196 VTAIL.n79 VTAIL.n70 12.0247
R197 VTAIL.n49 VTAIL.n40 12.0247
R198 VTAIL.n108 VTAIL.n96 11.249
R199 VTAIL.n18 VTAIL.n6 11.249
R200 VTAIL.n80 VTAIL.n68 11.249
R201 VTAIL.n50 VTAIL.n38 11.249
R202 VTAIL.n112 VTAIL.n111 10.4732
R203 VTAIL.n22 VTAIL.n21 10.4732
R204 VTAIL.n84 VTAIL.n83 10.4732
R205 VTAIL.n54 VTAIL.n53 10.4732
R206 VTAIL.n115 VTAIL.n94 9.69747
R207 VTAIL.n25 VTAIL.n4 9.69747
R208 VTAIL.n87 VTAIL.n66 9.69747
R209 VTAIL.n57 VTAIL.n36 9.69747
R210 VTAIL.n118 VTAIL.n117 9.45567
R211 VTAIL.n28 VTAIL.n27 9.45567
R212 VTAIL.n90 VTAIL.n89 9.45567
R213 VTAIL.n60 VTAIL.n59 9.45567
R214 VTAIL.n117 VTAIL.n116 9.3005
R215 VTAIL.n94 VTAIL.n93 9.3005
R216 VTAIL.n111 VTAIL.n110 9.3005
R217 VTAIL.n109 VTAIL.n108 9.3005
R218 VTAIL.n98 VTAIL.n97 9.3005
R219 VTAIL.n103 VTAIL.n102 9.3005
R220 VTAIL.n27 VTAIL.n26 9.3005
R221 VTAIL.n4 VTAIL.n3 9.3005
R222 VTAIL.n21 VTAIL.n20 9.3005
R223 VTAIL.n19 VTAIL.n18 9.3005
R224 VTAIL.n8 VTAIL.n7 9.3005
R225 VTAIL.n13 VTAIL.n12 9.3005
R226 VTAIL.n89 VTAIL.n88 9.3005
R227 VTAIL.n66 VTAIL.n65 9.3005
R228 VTAIL.n83 VTAIL.n82 9.3005
R229 VTAIL.n81 VTAIL.n80 9.3005
R230 VTAIL.n70 VTAIL.n69 9.3005
R231 VTAIL.n75 VTAIL.n74 9.3005
R232 VTAIL.n59 VTAIL.n58 9.3005
R233 VTAIL.n36 VTAIL.n35 9.3005
R234 VTAIL.n53 VTAIL.n52 9.3005
R235 VTAIL.n51 VTAIL.n50 9.3005
R236 VTAIL.n40 VTAIL.n39 9.3005
R237 VTAIL.n45 VTAIL.n44 9.3005
R238 VTAIL.n116 VTAIL.n92 8.92171
R239 VTAIL.n26 VTAIL.n2 8.92171
R240 VTAIL.n88 VTAIL.n64 8.92171
R241 VTAIL.n58 VTAIL.n34 8.92171
R242 VTAIL.n0 VTAIL.t4 6.0762
R243 VTAIL.n0 VTAIL.t3 6.0762
R244 VTAIL.n30 VTAIL.t10 6.0762
R245 VTAIL.n30 VTAIL.t11 6.0762
R246 VTAIL.n62 VTAIL.t8 6.0762
R247 VTAIL.n62 VTAIL.t9 6.0762
R248 VTAIL.n32 VTAIL.t5 6.0762
R249 VTAIL.n32 VTAIL.t0 6.0762
R250 VTAIL.n118 VTAIL.n92 5.04292
R251 VTAIL.n28 VTAIL.n2 5.04292
R252 VTAIL.n90 VTAIL.n64 5.04292
R253 VTAIL.n60 VTAIL.n34 5.04292
R254 VTAIL.n116 VTAIL.n115 4.26717
R255 VTAIL.n26 VTAIL.n25 4.26717
R256 VTAIL.n88 VTAIL.n87 4.26717
R257 VTAIL.n58 VTAIL.n57 4.26717
R258 VTAIL.n74 VTAIL.n73 3.71853
R259 VTAIL.n44 VTAIL.n43 3.71853
R260 VTAIL.n102 VTAIL.n101 3.71853
R261 VTAIL.n12 VTAIL.n11 3.71853
R262 VTAIL.n112 VTAIL.n94 3.49141
R263 VTAIL.n22 VTAIL.n4 3.49141
R264 VTAIL.n84 VTAIL.n66 3.49141
R265 VTAIL.n54 VTAIL.n36 3.49141
R266 VTAIL.n111 VTAIL.n96 2.71565
R267 VTAIL.n21 VTAIL.n6 2.71565
R268 VTAIL.n83 VTAIL.n68 2.71565
R269 VTAIL.n53 VTAIL.n38 2.71565
R270 VTAIL.n108 VTAIL.n107 1.93989
R271 VTAIL.n18 VTAIL.n17 1.93989
R272 VTAIL.n80 VTAIL.n79 1.93989
R273 VTAIL.n50 VTAIL.n49 1.93989
R274 VTAIL.n61 VTAIL.n33 1.16429
R275 VTAIL.n91 VTAIL.n63 1.16429
R276 VTAIL.n31 VTAIL.n29 1.16429
R277 VTAIL.n104 VTAIL.n98 1.16414
R278 VTAIL.n14 VTAIL.n8 1.16414
R279 VTAIL.n76 VTAIL.n70 1.16414
R280 VTAIL.n46 VTAIL.n40 1.16414
R281 VTAIL.n63 VTAIL.n61 1.05222
R282 VTAIL.n29 VTAIL.n1 1.05222
R283 VTAIL VTAIL.n119 0.815155
R284 VTAIL.n103 VTAIL.n100 0.388379
R285 VTAIL.n13 VTAIL.n10 0.388379
R286 VTAIL.n75 VTAIL.n72 0.388379
R287 VTAIL.n45 VTAIL.n42 0.388379
R288 VTAIL VTAIL.n1 0.349638
R289 VTAIL.n102 VTAIL.n97 0.155672
R290 VTAIL.n109 VTAIL.n97 0.155672
R291 VTAIL.n110 VTAIL.n109 0.155672
R292 VTAIL.n110 VTAIL.n93 0.155672
R293 VTAIL.n117 VTAIL.n93 0.155672
R294 VTAIL.n12 VTAIL.n7 0.155672
R295 VTAIL.n19 VTAIL.n7 0.155672
R296 VTAIL.n20 VTAIL.n19 0.155672
R297 VTAIL.n20 VTAIL.n3 0.155672
R298 VTAIL.n27 VTAIL.n3 0.155672
R299 VTAIL.n89 VTAIL.n65 0.155672
R300 VTAIL.n82 VTAIL.n65 0.155672
R301 VTAIL.n82 VTAIL.n81 0.155672
R302 VTAIL.n81 VTAIL.n69 0.155672
R303 VTAIL.n74 VTAIL.n69 0.155672
R304 VTAIL.n59 VTAIL.n35 0.155672
R305 VTAIL.n52 VTAIL.n35 0.155672
R306 VTAIL.n52 VTAIL.n51 0.155672
R307 VTAIL.n51 VTAIL.n39 0.155672
R308 VTAIL.n44 VTAIL.n39 0.155672
R309 VN.n1 VN.t3 187.69
R310 VN.n7 VN.t2 187.69
R311 VN.n4 VN.t0 165.156
R312 VN.n10 VN.t4 165.156
R313 VN.n9 VN.n6 161.3
R314 VN.n3 VN.n0 161.3
R315 VN.n2 VN.t5 126.407
R316 VN.n8 VN.t1 126.407
R317 VN.n11 VN.n10 80.6037
R318 VN.n5 VN.n4 80.6037
R319 VN.n4 VN.n3 48.6898
R320 VN.n10 VN.n9 48.6898
R321 VN VN.n11 37.8362
R322 VN.n2 VN.n1 32.2015
R323 VN.n8 VN.n7 32.2015
R324 VN.n7 VN.n6 28.3725
R325 VN.n1 VN.n0 28.3725
R326 VN.n3 VN.n2 24.4675
R327 VN.n9 VN.n8 24.4675
R328 VN.n11 VN.n6 0.285035
R329 VN.n5 VN.n0 0.285035
R330 VN VN.n5 0.146778
R331 VDD2.n51 VDD2.n29 756.745
R332 VDD2.n22 VDD2.n0 756.745
R333 VDD2.n52 VDD2.n51 585
R334 VDD2.n50 VDD2.n49 585
R335 VDD2.n33 VDD2.n32 585
R336 VDD2.n44 VDD2.n43 585
R337 VDD2.n42 VDD2.n41 585
R338 VDD2.n37 VDD2.n36 585
R339 VDD2.n8 VDD2.n7 585
R340 VDD2.n13 VDD2.n12 585
R341 VDD2.n15 VDD2.n14 585
R342 VDD2.n4 VDD2.n3 585
R343 VDD2.n21 VDD2.n20 585
R344 VDD2.n23 VDD2.n22 585
R345 VDD2.n38 VDD2.t1 327.856
R346 VDD2.n9 VDD2.t2 327.856
R347 VDD2.n51 VDD2.n50 171.744
R348 VDD2.n50 VDD2.n32 171.744
R349 VDD2.n43 VDD2.n32 171.744
R350 VDD2.n43 VDD2.n42 171.744
R351 VDD2.n42 VDD2.n36 171.744
R352 VDD2.n13 VDD2.n7 171.744
R353 VDD2.n14 VDD2.n13 171.744
R354 VDD2.n14 VDD2.n3 171.744
R355 VDD2.n21 VDD2.n3 171.744
R356 VDD2.n22 VDD2.n21 171.744
R357 VDD2.n28 VDD2.n27 98.9239
R358 VDD2 VDD2.n57 98.9211
R359 VDD2.t1 VDD2.n36 85.8723
R360 VDD2.t2 VDD2.n7 85.8723
R361 VDD2.n28 VDD2.n26 51.0392
R362 VDD2.n56 VDD2.n55 50.2217
R363 VDD2.n56 VDD2.n28 32.1097
R364 VDD2.n38 VDD2.n37 16.381
R365 VDD2.n9 VDD2.n8 16.381
R366 VDD2.n41 VDD2.n40 12.8005
R367 VDD2.n12 VDD2.n11 12.8005
R368 VDD2.n44 VDD2.n35 12.0247
R369 VDD2.n15 VDD2.n6 12.0247
R370 VDD2.n45 VDD2.n33 11.249
R371 VDD2.n16 VDD2.n4 11.249
R372 VDD2.n49 VDD2.n48 10.4732
R373 VDD2.n20 VDD2.n19 10.4732
R374 VDD2.n52 VDD2.n31 9.69747
R375 VDD2.n23 VDD2.n2 9.69747
R376 VDD2.n55 VDD2.n54 9.45567
R377 VDD2.n26 VDD2.n25 9.45567
R378 VDD2.n54 VDD2.n53 9.3005
R379 VDD2.n31 VDD2.n30 9.3005
R380 VDD2.n48 VDD2.n47 9.3005
R381 VDD2.n46 VDD2.n45 9.3005
R382 VDD2.n35 VDD2.n34 9.3005
R383 VDD2.n40 VDD2.n39 9.3005
R384 VDD2.n25 VDD2.n24 9.3005
R385 VDD2.n2 VDD2.n1 9.3005
R386 VDD2.n19 VDD2.n18 9.3005
R387 VDD2.n17 VDD2.n16 9.3005
R388 VDD2.n6 VDD2.n5 9.3005
R389 VDD2.n11 VDD2.n10 9.3005
R390 VDD2.n53 VDD2.n29 8.92171
R391 VDD2.n24 VDD2.n0 8.92171
R392 VDD2.n57 VDD2.t4 6.0762
R393 VDD2.n57 VDD2.t3 6.0762
R394 VDD2.n27 VDD2.t0 6.0762
R395 VDD2.n27 VDD2.t5 6.0762
R396 VDD2.n55 VDD2.n29 5.04292
R397 VDD2.n26 VDD2.n0 5.04292
R398 VDD2.n53 VDD2.n52 4.26717
R399 VDD2.n24 VDD2.n23 4.26717
R400 VDD2.n39 VDD2.n38 3.71853
R401 VDD2.n10 VDD2.n9 3.71853
R402 VDD2.n49 VDD2.n31 3.49141
R403 VDD2.n20 VDD2.n2 3.49141
R404 VDD2.n48 VDD2.n33 2.71565
R405 VDD2.n19 VDD2.n4 2.71565
R406 VDD2.n45 VDD2.n44 1.93989
R407 VDD2.n16 VDD2.n15 1.93989
R408 VDD2.n41 VDD2.n35 1.16414
R409 VDD2.n12 VDD2.n6 1.16414
R410 VDD2 VDD2.n56 0.931535
R411 VDD2.n40 VDD2.n37 0.388379
R412 VDD2.n11 VDD2.n8 0.388379
R413 VDD2.n54 VDD2.n30 0.155672
R414 VDD2.n47 VDD2.n30 0.155672
R415 VDD2.n47 VDD2.n46 0.155672
R416 VDD2.n46 VDD2.n34 0.155672
R417 VDD2.n39 VDD2.n34 0.155672
R418 VDD2.n10 VDD2.n5 0.155672
R419 VDD2.n17 VDD2.n5 0.155672
R420 VDD2.n18 VDD2.n17 0.155672
R421 VDD2.n18 VDD2.n1 0.155672
R422 VDD2.n25 VDD2.n1 0.155672
R423 B.n304 B.n45 585
R424 B.n306 B.n305 585
R425 B.n307 B.n44 585
R426 B.n309 B.n308 585
R427 B.n310 B.n43 585
R428 B.n312 B.n311 585
R429 B.n313 B.n42 585
R430 B.n315 B.n314 585
R431 B.n316 B.n41 585
R432 B.n318 B.n317 585
R433 B.n319 B.n40 585
R434 B.n321 B.n320 585
R435 B.n322 B.n39 585
R436 B.n324 B.n323 585
R437 B.n325 B.n38 585
R438 B.n327 B.n326 585
R439 B.n328 B.n37 585
R440 B.n330 B.n329 585
R441 B.n331 B.n36 585
R442 B.n333 B.n332 585
R443 B.n334 B.n35 585
R444 B.n336 B.n335 585
R445 B.n338 B.n337 585
R446 B.n339 B.n31 585
R447 B.n341 B.n340 585
R448 B.n342 B.n30 585
R449 B.n344 B.n343 585
R450 B.n345 B.n29 585
R451 B.n347 B.n346 585
R452 B.n348 B.n28 585
R453 B.n350 B.n349 585
R454 B.n351 B.n25 585
R455 B.n354 B.n353 585
R456 B.n355 B.n24 585
R457 B.n357 B.n356 585
R458 B.n358 B.n23 585
R459 B.n360 B.n359 585
R460 B.n361 B.n22 585
R461 B.n363 B.n362 585
R462 B.n364 B.n21 585
R463 B.n366 B.n365 585
R464 B.n367 B.n20 585
R465 B.n369 B.n368 585
R466 B.n370 B.n19 585
R467 B.n372 B.n371 585
R468 B.n373 B.n18 585
R469 B.n375 B.n374 585
R470 B.n376 B.n17 585
R471 B.n378 B.n377 585
R472 B.n379 B.n16 585
R473 B.n381 B.n380 585
R474 B.n382 B.n15 585
R475 B.n384 B.n383 585
R476 B.n385 B.n14 585
R477 B.n303 B.n302 585
R478 B.n301 B.n46 585
R479 B.n300 B.n299 585
R480 B.n298 B.n47 585
R481 B.n297 B.n296 585
R482 B.n295 B.n48 585
R483 B.n294 B.n293 585
R484 B.n292 B.n49 585
R485 B.n291 B.n290 585
R486 B.n289 B.n50 585
R487 B.n288 B.n287 585
R488 B.n286 B.n51 585
R489 B.n285 B.n284 585
R490 B.n283 B.n52 585
R491 B.n282 B.n281 585
R492 B.n280 B.n53 585
R493 B.n279 B.n278 585
R494 B.n277 B.n54 585
R495 B.n276 B.n275 585
R496 B.n274 B.n55 585
R497 B.n273 B.n272 585
R498 B.n271 B.n56 585
R499 B.n270 B.n269 585
R500 B.n268 B.n57 585
R501 B.n267 B.n266 585
R502 B.n265 B.n58 585
R503 B.n264 B.n263 585
R504 B.n262 B.n59 585
R505 B.n261 B.n260 585
R506 B.n259 B.n60 585
R507 B.n258 B.n257 585
R508 B.n256 B.n61 585
R509 B.n255 B.n254 585
R510 B.n253 B.n62 585
R511 B.n252 B.n251 585
R512 B.n250 B.n63 585
R513 B.n249 B.n248 585
R514 B.n247 B.n64 585
R515 B.n246 B.n245 585
R516 B.n244 B.n65 585
R517 B.n243 B.n242 585
R518 B.n241 B.n66 585
R519 B.n240 B.n239 585
R520 B.n238 B.n67 585
R521 B.n237 B.n236 585
R522 B.n235 B.n68 585
R523 B.n234 B.n233 585
R524 B.n232 B.n69 585
R525 B.n231 B.n230 585
R526 B.n148 B.n101 585
R527 B.n150 B.n149 585
R528 B.n151 B.n100 585
R529 B.n153 B.n152 585
R530 B.n154 B.n99 585
R531 B.n156 B.n155 585
R532 B.n157 B.n98 585
R533 B.n159 B.n158 585
R534 B.n160 B.n97 585
R535 B.n162 B.n161 585
R536 B.n163 B.n96 585
R537 B.n165 B.n164 585
R538 B.n166 B.n95 585
R539 B.n168 B.n167 585
R540 B.n169 B.n94 585
R541 B.n171 B.n170 585
R542 B.n172 B.n93 585
R543 B.n174 B.n173 585
R544 B.n175 B.n92 585
R545 B.n177 B.n176 585
R546 B.n178 B.n91 585
R547 B.n180 B.n179 585
R548 B.n182 B.n181 585
R549 B.n183 B.n87 585
R550 B.n185 B.n184 585
R551 B.n186 B.n86 585
R552 B.n188 B.n187 585
R553 B.n189 B.n85 585
R554 B.n191 B.n190 585
R555 B.n192 B.n84 585
R556 B.n194 B.n193 585
R557 B.n195 B.n81 585
R558 B.n198 B.n197 585
R559 B.n199 B.n80 585
R560 B.n201 B.n200 585
R561 B.n202 B.n79 585
R562 B.n204 B.n203 585
R563 B.n205 B.n78 585
R564 B.n207 B.n206 585
R565 B.n208 B.n77 585
R566 B.n210 B.n209 585
R567 B.n211 B.n76 585
R568 B.n213 B.n212 585
R569 B.n214 B.n75 585
R570 B.n216 B.n215 585
R571 B.n217 B.n74 585
R572 B.n219 B.n218 585
R573 B.n220 B.n73 585
R574 B.n222 B.n221 585
R575 B.n223 B.n72 585
R576 B.n225 B.n224 585
R577 B.n226 B.n71 585
R578 B.n228 B.n227 585
R579 B.n229 B.n70 585
R580 B.n147 B.n146 585
R581 B.n145 B.n102 585
R582 B.n144 B.n143 585
R583 B.n142 B.n103 585
R584 B.n141 B.n140 585
R585 B.n139 B.n104 585
R586 B.n138 B.n137 585
R587 B.n136 B.n105 585
R588 B.n135 B.n134 585
R589 B.n133 B.n106 585
R590 B.n132 B.n131 585
R591 B.n130 B.n107 585
R592 B.n129 B.n128 585
R593 B.n127 B.n108 585
R594 B.n126 B.n125 585
R595 B.n124 B.n109 585
R596 B.n123 B.n122 585
R597 B.n121 B.n110 585
R598 B.n120 B.n119 585
R599 B.n118 B.n111 585
R600 B.n117 B.n116 585
R601 B.n115 B.n112 585
R602 B.n114 B.n113 585
R603 B.n2 B.n0 585
R604 B.n421 B.n1 585
R605 B.n420 B.n419 585
R606 B.n418 B.n3 585
R607 B.n417 B.n416 585
R608 B.n415 B.n4 585
R609 B.n414 B.n413 585
R610 B.n412 B.n5 585
R611 B.n411 B.n410 585
R612 B.n409 B.n6 585
R613 B.n408 B.n407 585
R614 B.n406 B.n7 585
R615 B.n405 B.n404 585
R616 B.n403 B.n8 585
R617 B.n402 B.n401 585
R618 B.n400 B.n9 585
R619 B.n399 B.n398 585
R620 B.n397 B.n10 585
R621 B.n396 B.n395 585
R622 B.n394 B.n11 585
R623 B.n393 B.n392 585
R624 B.n391 B.n12 585
R625 B.n390 B.n389 585
R626 B.n388 B.n13 585
R627 B.n387 B.n386 585
R628 B.n423 B.n422 585
R629 B.n146 B.n101 473.281
R630 B.n386 B.n385 473.281
R631 B.n230 B.n229 473.281
R632 B.n302 B.n45 473.281
R633 B.n82 B.t6 329.466
R634 B.n88 B.t3 329.466
R635 B.n26 B.t9 329.466
R636 B.n32 B.t0 329.466
R637 B.n82 B.t8 283.188
R638 B.n32 B.t1 283.188
R639 B.n88 B.t5 283.188
R640 B.n26 B.t10 283.188
R641 B.n83 B.t7 257.005
R642 B.n33 B.t2 257.005
R643 B.n89 B.t4 257.005
R644 B.n27 B.t11 257.005
R645 B.n146 B.n145 163.367
R646 B.n145 B.n144 163.367
R647 B.n144 B.n103 163.367
R648 B.n140 B.n103 163.367
R649 B.n140 B.n139 163.367
R650 B.n139 B.n138 163.367
R651 B.n138 B.n105 163.367
R652 B.n134 B.n105 163.367
R653 B.n134 B.n133 163.367
R654 B.n133 B.n132 163.367
R655 B.n132 B.n107 163.367
R656 B.n128 B.n107 163.367
R657 B.n128 B.n127 163.367
R658 B.n127 B.n126 163.367
R659 B.n126 B.n109 163.367
R660 B.n122 B.n109 163.367
R661 B.n122 B.n121 163.367
R662 B.n121 B.n120 163.367
R663 B.n120 B.n111 163.367
R664 B.n116 B.n111 163.367
R665 B.n116 B.n115 163.367
R666 B.n115 B.n114 163.367
R667 B.n114 B.n2 163.367
R668 B.n422 B.n2 163.367
R669 B.n422 B.n421 163.367
R670 B.n421 B.n420 163.367
R671 B.n420 B.n3 163.367
R672 B.n416 B.n3 163.367
R673 B.n416 B.n415 163.367
R674 B.n415 B.n414 163.367
R675 B.n414 B.n5 163.367
R676 B.n410 B.n5 163.367
R677 B.n410 B.n409 163.367
R678 B.n409 B.n408 163.367
R679 B.n408 B.n7 163.367
R680 B.n404 B.n7 163.367
R681 B.n404 B.n403 163.367
R682 B.n403 B.n402 163.367
R683 B.n402 B.n9 163.367
R684 B.n398 B.n9 163.367
R685 B.n398 B.n397 163.367
R686 B.n397 B.n396 163.367
R687 B.n396 B.n11 163.367
R688 B.n392 B.n11 163.367
R689 B.n392 B.n391 163.367
R690 B.n391 B.n390 163.367
R691 B.n390 B.n13 163.367
R692 B.n386 B.n13 163.367
R693 B.n150 B.n101 163.367
R694 B.n151 B.n150 163.367
R695 B.n152 B.n151 163.367
R696 B.n152 B.n99 163.367
R697 B.n156 B.n99 163.367
R698 B.n157 B.n156 163.367
R699 B.n158 B.n157 163.367
R700 B.n158 B.n97 163.367
R701 B.n162 B.n97 163.367
R702 B.n163 B.n162 163.367
R703 B.n164 B.n163 163.367
R704 B.n164 B.n95 163.367
R705 B.n168 B.n95 163.367
R706 B.n169 B.n168 163.367
R707 B.n170 B.n169 163.367
R708 B.n170 B.n93 163.367
R709 B.n174 B.n93 163.367
R710 B.n175 B.n174 163.367
R711 B.n176 B.n175 163.367
R712 B.n176 B.n91 163.367
R713 B.n180 B.n91 163.367
R714 B.n181 B.n180 163.367
R715 B.n181 B.n87 163.367
R716 B.n185 B.n87 163.367
R717 B.n186 B.n185 163.367
R718 B.n187 B.n186 163.367
R719 B.n187 B.n85 163.367
R720 B.n191 B.n85 163.367
R721 B.n192 B.n191 163.367
R722 B.n193 B.n192 163.367
R723 B.n193 B.n81 163.367
R724 B.n198 B.n81 163.367
R725 B.n199 B.n198 163.367
R726 B.n200 B.n199 163.367
R727 B.n200 B.n79 163.367
R728 B.n204 B.n79 163.367
R729 B.n205 B.n204 163.367
R730 B.n206 B.n205 163.367
R731 B.n206 B.n77 163.367
R732 B.n210 B.n77 163.367
R733 B.n211 B.n210 163.367
R734 B.n212 B.n211 163.367
R735 B.n212 B.n75 163.367
R736 B.n216 B.n75 163.367
R737 B.n217 B.n216 163.367
R738 B.n218 B.n217 163.367
R739 B.n218 B.n73 163.367
R740 B.n222 B.n73 163.367
R741 B.n223 B.n222 163.367
R742 B.n224 B.n223 163.367
R743 B.n224 B.n71 163.367
R744 B.n228 B.n71 163.367
R745 B.n229 B.n228 163.367
R746 B.n230 B.n69 163.367
R747 B.n234 B.n69 163.367
R748 B.n235 B.n234 163.367
R749 B.n236 B.n235 163.367
R750 B.n236 B.n67 163.367
R751 B.n240 B.n67 163.367
R752 B.n241 B.n240 163.367
R753 B.n242 B.n241 163.367
R754 B.n242 B.n65 163.367
R755 B.n246 B.n65 163.367
R756 B.n247 B.n246 163.367
R757 B.n248 B.n247 163.367
R758 B.n248 B.n63 163.367
R759 B.n252 B.n63 163.367
R760 B.n253 B.n252 163.367
R761 B.n254 B.n253 163.367
R762 B.n254 B.n61 163.367
R763 B.n258 B.n61 163.367
R764 B.n259 B.n258 163.367
R765 B.n260 B.n259 163.367
R766 B.n260 B.n59 163.367
R767 B.n264 B.n59 163.367
R768 B.n265 B.n264 163.367
R769 B.n266 B.n265 163.367
R770 B.n266 B.n57 163.367
R771 B.n270 B.n57 163.367
R772 B.n271 B.n270 163.367
R773 B.n272 B.n271 163.367
R774 B.n272 B.n55 163.367
R775 B.n276 B.n55 163.367
R776 B.n277 B.n276 163.367
R777 B.n278 B.n277 163.367
R778 B.n278 B.n53 163.367
R779 B.n282 B.n53 163.367
R780 B.n283 B.n282 163.367
R781 B.n284 B.n283 163.367
R782 B.n284 B.n51 163.367
R783 B.n288 B.n51 163.367
R784 B.n289 B.n288 163.367
R785 B.n290 B.n289 163.367
R786 B.n290 B.n49 163.367
R787 B.n294 B.n49 163.367
R788 B.n295 B.n294 163.367
R789 B.n296 B.n295 163.367
R790 B.n296 B.n47 163.367
R791 B.n300 B.n47 163.367
R792 B.n301 B.n300 163.367
R793 B.n302 B.n301 163.367
R794 B.n385 B.n384 163.367
R795 B.n384 B.n15 163.367
R796 B.n380 B.n15 163.367
R797 B.n380 B.n379 163.367
R798 B.n379 B.n378 163.367
R799 B.n378 B.n17 163.367
R800 B.n374 B.n17 163.367
R801 B.n374 B.n373 163.367
R802 B.n373 B.n372 163.367
R803 B.n372 B.n19 163.367
R804 B.n368 B.n19 163.367
R805 B.n368 B.n367 163.367
R806 B.n367 B.n366 163.367
R807 B.n366 B.n21 163.367
R808 B.n362 B.n21 163.367
R809 B.n362 B.n361 163.367
R810 B.n361 B.n360 163.367
R811 B.n360 B.n23 163.367
R812 B.n356 B.n23 163.367
R813 B.n356 B.n355 163.367
R814 B.n355 B.n354 163.367
R815 B.n354 B.n25 163.367
R816 B.n349 B.n25 163.367
R817 B.n349 B.n348 163.367
R818 B.n348 B.n347 163.367
R819 B.n347 B.n29 163.367
R820 B.n343 B.n29 163.367
R821 B.n343 B.n342 163.367
R822 B.n342 B.n341 163.367
R823 B.n341 B.n31 163.367
R824 B.n337 B.n31 163.367
R825 B.n337 B.n336 163.367
R826 B.n336 B.n35 163.367
R827 B.n332 B.n35 163.367
R828 B.n332 B.n331 163.367
R829 B.n331 B.n330 163.367
R830 B.n330 B.n37 163.367
R831 B.n326 B.n37 163.367
R832 B.n326 B.n325 163.367
R833 B.n325 B.n324 163.367
R834 B.n324 B.n39 163.367
R835 B.n320 B.n39 163.367
R836 B.n320 B.n319 163.367
R837 B.n319 B.n318 163.367
R838 B.n318 B.n41 163.367
R839 B.n314 B.n41 163.367
R840 B.n314 B.n313 163.367
R841 B.n313 B.n312 163.367
R842 B.n312 B.n43 163.367
R843 B.n308 B.n43 163.367
R844 B.n308 B.n307 163.367
R845 B.n307 B.n306 163.367
R846 B.n306 B.n45 163.367
R847 B.n196 B.n83 59.5399
R848 B.n90 B.n89 59.5399
R849 B.n352 B.n27 59.5399
R850 B.n34 B.n33 59.5399
R851 B.n387 B.n14 30.7517
R852 B.n304 B.n303 30.7517
R853 B.n231 B.n70 30.7517
R854 B.n148 B.n147 30.7517
R855 B.n83 B.n82 26.1823
R856 B.n89 B.n88 26.1823
R857 B.n27 B.n26 26.1823
R858 B.n33 B.n32 26.1823
R859 B B.n423 18.0485
R860 B.n383 B.n14 10.6151
R861 B.n383 B.n382 10.6151
R862 B.n382 B.n381 10.6151
R863 B.n381 B.n16 10.6151
R864 B.n377 B.n16 10.6151
R865 B.n377 B.n376 10.6151
R866 B.n376 B.n375 10.6151
R867 B.n375 B.n18 10.6151
R868 B.n371 B.n18 10.6151
R869 B.n371 B.n370 10.6151
R870 B.n370 B.n369 10.6151
R871 B.n369 B.n20 10.6151
R872 B.n365 B.n20 10.6151
R873 B.n365 B.n364 10.6151
R874 B.n364 B.n363 10.6151
R875 B.n363 B.n22 10.6151
R876 B.n359 B.n22 10.6151
R877 B.n359 B.n358 10.6151
R878 B.n358 B.n357 10.6151
R879 B.n357 B.n24 10.6151
R880 B.n353 B.n24 10.6151
R881 B.n351 B.n350 10.6151
R882 B.n350 B.n28 10.6151
R883 B.n346 B.n28 10.6151
R884 B.n346 B.n345 10.6151
R885 B.n345 B.n344 10.6151
R886 B.n344 B.n30 10.6151
R887 B.n340 B.n30 10.6151
R888 B.n340 B.n339 10.6151
R889 B.n339 B.n338 10.6151
R890 B.n335 B.n334 10.6151
R891 B.n334 B.n333 10.6151
R892 B.n333 B.n36 10.6151
R893 B.n329 B.n36 10.6151
R894 B.n329 B.n328 10.6151
R895 B.n328 B.n327 10.6151
R896 B.n327 B.n38 10.6151
R897 B.n323 B.n38 10.6151
R898 B.n323 B.n322 10.6151
R899 B.n322 B.n321 10.6151
R900 B.n321 B.n40 10.6151
R901 B.n317 B.n40 10.6151
R902 B.n317 B.n316 10.6151
R903 B.n316 B.n315 10.6151
R904 B.n315 B.n42 10.6151
R905 B.n311 B.n42 10.6151
R906 B.n311 B.n310 10.6151
R907 B.n310 B.n309 10.6151
R908 B.n309 B.n44 10.6151
R909 B.n305 B.n44 10.6151
R910 B.n305 B.n304 10.6151
R911 B.n232 B.n231 10.6151
R912 B.n233 B.n232 10.6151
R913 B.n233 B.n68 10.6151
R914 B.n237 B.n68 10.6151
R915 B.n238 B.n237 10.6151
R916 B.n239 B.n238 10.6151
R917 B.n239 B.n66 10.6151
R918 B.n243 B.n66 10.6151
R919 B.n244 B.n243 10.6151
R920 B.n245 B.n244 10.6151
R921 B.n245 B.n64 10.6151
R922 B.n249 B.n64 10.6151
R923 B.n250 B.n249 10.6151
R924 B.n251 B.n250 10.6151
R925 B.n251 B.n62 10.6151
R926 B.n255 B.n62 10.6151
R927 B.n256 B.n255 10.6151
R928 B.n257 B.n256 10.6151
R929 B.n257 B.n60 10.6151
R930 B.n261 B.n60 10.6151
R931 B.n262 B.n261 10.6151
R932 B.n263 B.n262 10.6151
R933 B.n263 B.n58 10.6151
R934 B.n267 B.n58 10.6151
R935 B.n268 B.n267 10.6151
R936 B.n269 B.n268 10.6151
R937 B.n269 B.n56 10.6151
R938 B.n273 B.n56 10.6151
R939 B.n274 B.n273 10.6151
R940 B.n275 B.n274 10.6151
R941 B.n275 B.n54 10.6151
R942 B.n279 B.n54 10.6151
R943 B.n280 B.n279 10.6151
R944 B.n281 B.n280 10.6151
R945 B.n281 B.n52 10.6151
R946 B.n285 B.n52 10.6151
R947 B.n286 B.n285 10.6151
R948 B.n287 B.n286 10.6151
R949 B.n287 B.n50 10.6151
R950 B.n291 B.n50 10.6151
R951 B.n292 B.n291 10.6151
R952 B.n293 B.n292 10.6151
R953 B.n293 B.n48 10.6151
R954 B.n297 B.n48 10.6151
R955 B.n298 B.n297 10.6151
R956 B.n299 B.n298 10.6151
R957 B.n299 B.n46 10.6151
R958 B.n303 B.n46 10.6151
R959 B.n149 B.n148 10.6151
R960 B.n149 B.n100 10.6151
R961 B.n153 B.n100 10.6151
R962 B.n154 B.n153 10.6151
R963 B.n155 B.n154 10.6151
R964 B.n155 B.n98 10.6151
R965 B.n159 B.n98 10.6151
R966 B.n160 B.n159 10.6151
R967 B.n161 B.n160 10.6151
R968 B.n161 B.n96 10.6151
R969 B.n165 B.n96 10.6151
R970 B.n166 B.n165 10.6151
R971 B.n167 B.n166 10.6151
R972 B.n167 B.n94 10.6151
R973 B.n171 B.n94 10.6151
R974 B.n172 B.n171 10.6151
R975 B.n173 B.n172 10.6151
R976 B.n173 B.n92 10.6151
R977 B.n177 B.n92 10.6151
R978 B.n178 B.n177 10.6151
R979 B.n179 B.n178 10.6151
R980 B.n183 B.n182 10.6151
R981 B.n184 B.n183 10.6151
R982 B.n184 B.n86 10.6151
R983 B.n188 B.n86 10.6151
R984 B.n189 B.n188 10.6151
R985 B.n190 B.n189 10.6151
R986 B.n190 B.n84 10.6151
R987 B.n194 B.n84 10.6151
R988 B.n195 B.n194 10.6151
R989 B.n197 B.n80 10.6151
R990 B.n201 B.n80 10.6151
R991 B.n202 B.n201 10.6151
R992 B.n203 B.n202 10.6151
R993 B.n203 B.n78 10.6151
R994 B.n207 B.n78 10.6151
R995 B.n208 B.n207 10.6151
R996 B.n209 B.n208 10.6151
R997 B.n209 B.n76 10.6151
R998 B.n213 B.n76 10.6151
R999 B.n214 B.n213 10.6151
R1000 B.n215 B.n214 10.6151
R1001 B.n215 B.n74 10.6151
R1002 B.n219 B.n74 10.6151
R1003 B.n220 B.n219 10.6151
R1004 B.n221 B.n220 10.6151
R1005 B.n221 B.n72 10.6151
R1006 B.n225 B.n72 10.6151
R1007 B.n226 B.n225 10.6151
R1008 B.n227 B.n226 10.6151
R1009 B.n227 B.n70 10.6151
R1010 B.n147 B.n102 10.6151
R1011 B.n143 B.n102 10.6151
R1012 B.n143 B.n142 10.6151
R1013 B.n142 B.n141 10.6151
R1014 B.n141 B.n104 10.6151
R1015 B.n137 B.n104 10.6151
R1016 B.n137 B.n136 10.6151
R1017 B.n136 B.n135 10.6151
R1018 B.n135 B.n106 10.6151
R1019 B.n131 B.n106 10.6151
R1020 B.n131 B.n130 10.6151
R1021 B.n130 B.n129 10.6151
R1022 B.n129 B.n108 10.6151
R1023 B.n125 B.n108 10.6151
R1024 B.n125 B.n124 10.6151
R1025 B.n124 B.n123 10.6151
R1026 B.n123 B.n110 10.6151
R1027 B.n119 B.n110 10.6151
R1028 B.n119 B.n118 10.6151
R1029 B.n118 B.n117 10.6151
R1030 B.n117 B.n112 10.6151
R1031 B.n113 B.n112 10.6151
R1032 B.n113 B.n0 10.6151
R1033 B.n419 B.n1 10.6151
R1034 B.n419 B.n418 10.6151
R1035 B.n418 B.n417 10.6151
R1036 B.n417 B.n4 10.6151
R1037 B.n413 B.n4 10.6151
R1038 B.n413 B.n412 10.6151
R1039 B.n412 B.n411 10.6151
R1040 B.n411 B.n6 10.6151
R1041 B.n407 B.n6 10.6151
R1042 B.n407 B.n406 10.6151
R1043 B.n406 B.n405 10.6151
R1044 B.n405 B.n8 10.6151
R1045 B.n401 B.n8 10.6151
R1046 B.n401 B.n400 10.6151
R1047 B.n400 B.n399 10.6151
R1048 B.n399 B.n10 10.6151
R1049 B.n395 B.n10 10.6151
R1050 B.n395 B.n394 10.6151
R1051 B.n394 B.n393 10.6151
R1052 B.n393 B.n12 10.6151
R1053 B.n389 B.n12 10.6151
R1054 B.n389 B.n388 10.6151
R1055 B.n388 B.n387 10.6151
R1056 B.n353 B.n352 9.36635
R1057 B.n335 B.n34 9.36635
R1058 B.n179 B.n90 9.36635
R1059 B.n197 B.n196 9.36635
R1060 B.n423 B.n0 2.81026
R1061 B.n423 B.n1 2.81026
R1062 B.n352 B.n351 1.24928
R1063 B.n338 B.n34 1.24928
R1064 B.n182 B.n90 1.24928
R1065 B.n196 B.n195 1.24928
C0 B VTAIL 1.64798f
C1 VDD1 VTAIL 5.07741f
C2 VP w_n2050_n2038# 3.64087f
C3 VP VN 4.16236f
C4 w_n2050_n2038# VN 3.3803f
C5 B VDD2 1.19832f
C6 VDD1 VDD2 0.826704f
C7 VP VTAIL 2.61138f
C8 VDD1 B 1.1617f
C9 w_n2050_n2038# VTAIL 1.90035f
C10 VTAIL VN 2.59709f
C11 VP VDD2 0.327701f
C12 w_n2050_n2038# VDD2 1.44787f
C13 VDD2 VN 2.4793f
C14 B VP 1.17785f
C15 B w_n2050_n2038# 5.63436f
C16 B VN 0.750656f
C17 VDD1 VP 2.65231f
C18 VDD1 w_n2050_n2038# 1.41382f
C19 VDD1 VN 0.14864f
C20 VTAIL VDD2 5.11785f
C21 VDD2 VSUBS 1.066937f
C22 VDD1 VSUBS 1.017476f
C23 VTAIL VSUBS 0.459998f
C24 VN VSUBS 4.167429f
C25 VP VSUBS 1.404639f
C26 B VSUBS 2.430558f
C27 w_n2050_n2038# VSUBS 52.275f
C28 B.n0 VSUBS 0.004175f
C29 B.n1 VSUBS 0.004175f
C30 B.n2 VSUBS 0.006602f
C31 B.n3 VSUBS 0.006602f
C32 B.n4 VSUBS 0.006602f
C33 B.n5 VSUBS 0.006602f
C34 B.n6 VSUBS 0.006602f
C35 B.n7 VSUBS 0.006602f
C36 B.n8 VSUBS 0.006602f
C37 B.n9 VSUBS 0.006602f
C38 B.n10 VSUBS 0.006602f
C39 B.n11 VSUBS 0.006602f
C40 B.n12 VSUBS 0.006602f
C41 B.n13 VSUBS 0.006602f
C42 B.n14 VSUBS 0.01535f
C43 B.n15 VSUBS 0.006602f
C44 B.n16 VSUBS 0.006602f
C45 B.n17 VSUBS 0.006602f
C46 B.n18 VSUBS 0.006602f
C47 B.n19 VSUBS 0.006602f
C48 B.n20 VSUBS 0.006602f
C49 B.n21 VSUBS 0.006602f
C50 B.n22 VSUBS 0.006602f
C51 B.n23 VSUBS 0.006602f
C52 B.n24 VSUBS 0.006602f
C53 B.n25 VSUBS 0.006602f
C54 B.t11 VSUBS 0.074102f
C55 B.t10 VSUBS 0.085205f
C56 B.t9 VSUBS 0.231322f
C57 B.n26 VSUBS 0.151841f
C58 B.n27 VSUBS 0.129518f
C59 B.n28 VSUBS 0.006602f
C60 B.n29 VSUBS 0.006602f
C61 B.n30 VSUBS 0.006602f
C62 B.n31 VSUBS 0.006602f
C63 B.t2 VSUBS 0.074103f
C64 B.t1 VSUBS 0.085207f
C65 B.t0 VSUBS 0.231322f
C66 B.n32 VSUBS 0.15184f
C67 B.n33 VSUBS 0.129517f
C68 B.n34 VSUBS 0.015297f
C69 B.n35 VSUBS 0.006602f
C70 B.n36 VSUBS 0.006602f
C71 B.n37 VSUBS 0.006602f
C72 B.n38 VSUBS 0.006602f
C73 B.n39 VSUBS 0.006602f
C74 B.n40 VSUBS 0.006602f
C75 B.n41 VSUBS 0.006602f
C76 B.n42 VSUBS 0.006602f
C77 B.n43 VSUBS 0.006602f
C78 B.n44 VSUBS 0.006602f
C79 B.n45 VSUBS 0.01535f
C80 B.n46 VSUBS 0.006602f
C81 B.n47 VSUBS 0.006602f
C82 B.n48 VSUBS 0.006602f
C83 B.n49 VSUBS 0.006602f
C84 B.n50 VSUBS 0.006602f
C85 B.n51 VSUBS 0.006602f
C86 B.n52 VSUBS 0.006602f
C87 B.n53 VSUBS 0.006602f
C88 B.n54 VSUBS 0.006602f
C89 B.n55 VSUBS 0.006602f
C90 B.n56 VSUBS 0.006602f
C91 B.n57 VSUBS 0.006602f
C92 B.n58 VSUBS 0.006602f
C93 B.n59 VSUBS 0.006602f
C94 B.n60 VSUBS 0.006602f
C95 B.n61 VSUBS 0.006602f
C96 B.n62 VSUBS 0.006602f
C97 B.n63 VSUBS 0.006602f
C98 B.n64 VSUBS 0.006602f
C99 B.n65 VSUBS 0.006602f
C100 B.n66 VSUBS 0.006602f
C101 B.n67 VSUBS 0.006602f
C102 B.n68 VSUBS 0.006602f
C103 B.n69 VSUBS 0.006602f
C104 B.n70 VSUBS 0.01535f
C105 B.n71 VSUBS 0.006602f
C106 B.n72 VSUBS 0.006602f
C107 B.n73 VSUBS 0.006602f
C108 B.n74 VSUBS 0.006602f
C109 B.n75 VSUBS 0.006602f
C110 B.n76 VSUBS 0.006602f
C111 B.n77 VSUBS 0.006602f
C112 B.n78 VSUBS 0.006602f
C113 B.n79 VSUBS 0.006602f
C114 B.n80 VSUBS 0.006602f
C115 B.n81 VSUBS 0.006602f
C116 B.t7 VSUBS 0.074103f
C117 B.t8 VSUBS 0.085207f
C118 B.t6 VSUBS 0.231322f
C119 B.n82 VSUBS 0.15184f
C120 B.n83 VSUBS 0.129517f
C121 B.n84 VSUBS 0.006602f
C122 B.n85 VSUBS 0.006602f
C123 B.n86 VSUBS 0.006602f
C124 B.n87 VSUBS 0.006602f
C125 B.t4 VSUBS 0.074102f
C126 B.t5 VSUBS 0.085205f
C127 B.t3 VSUBS 0.231322f
C128 B.n88 VSUBS 0.151841f
C129 B.n89 VSUBS 0.129518f
C130 B.n90 VSUBS 0.015297f
C131 B.n91 VSUBS 0.006602f
C132 B.n92 VSUBS 0.006602f
C133 B.n93 VSUBS 0.006602f
C134 B.n94 VSUBS 0.006602f
C135 B.n95 VSUBS 0.006602f
C136 B.n96 VSUBS 0.006602f
C137 B.n97 VSUBS 0.006602f
C138 B.n98 VSUBS 0.006602f
C139 B.n99 VSUBS 0.006602f
C140 B.n100 VSUBS 0.006602f
C141 B.n101 VSUBS 0.01535f
C142 B.n102 VSUBS 0.006602f
C143 B.n103 VSUBS 0.006602f
C144 B.n104 VSUBS 0.006602f
C145 B.n105 VSUBS 0.006602f
C146 B.n106 VSUBS 0.006602f
C147 B.n107 VSUBS 0.006602f
C148 B.n108 VSUBS 0.006602f
C149 B.n109 VSUBS 0.006602f
C150 B.n110 VSUBS 0.006602f
C151 B.n111 VSUBS 0.006602f
C152 B.n112 VSUBS 0.006602f
C153 B.n113 VSUBS 0.006602f
C154 B.n114 VSUBS 0.006602f
C155 B.n115 VSUBS 0.006602f
C156 B.n116 VSUBS 0.006602f
C157 B.n117 VSUBS 0.006602f
C158 B.n118 VSUBS 0.006602f
C159 B.n119 VSUBS 0.006602f
C160 B.n120 VSUBS 0.006602f
C161 B.n121 VSUBS 0.006602f
C162 B.n122 VSUBS 0.006602f
C163 B.n123 VSUBS 0.006602f
C164 B.n124 VSUBS 0.006602f
C165 B.n125 VSUBS 0.006602f
C166 B.n126 VSUBS 0.006602f
C167 B.n127 VSUBS 0.006602f
C168 B.n128 VSUBS 0.006602f
C169 B.n129 VSUBS 0.006602f
C170 B.n130 VSUBS 0.006602f
C171 B.n131 VSUBS 0.006602f
C172 B.n132 VSUBS 0.006602f
C173 B.n133 VSUBS 0.006602f
C174 B.n134 VSUBS 0.006602f
C175 B.n135 VSUBS 0.006602f
C176 B.n136 VSUBS 0.006602f
C177 B.n137 VSUBS 0.006602f
C178 B.n138 VSUBS 0.006602f
C179 B.n139 VSUBS 0.006602f
C180 B.n140 VSUBS 0.006602f
C181 B.n141 VSUBS 0.006602f
C182 B.n142 VSUBS 0.006602f
C183 B.n143 VSUBS 0.006602f
C184 B.n144 VSUBS 0.006602f
C185 B.n145 VSUBS 0.006602f
C186 B.n146 VSUBS 0.01436f
C187 B.n147 VSUBS 0.01436f
C188 B.n148 VSUBS 0.01535f
C189 B.n149 VSUBS 0.006602f
C190 B.n150 VSUBS 0.006602f
C191 B.n151 VSUBS 0.006602f
C192 B.n152 VSUBS 0.006602f
C193 B.n153 VSUBS 0.006602f
C194 B.n154 VSUBS 0.006602f
C195 B.n155 VSUBS 0.006602f
C196 B.n156 VSUBS 0.006602f
C197 B.n157 VSUBS 0.006602f
C198 B.n158 VSUBS 0.006602f
C199 B.n159 VSUBS 0.006602f
C200 B.n160 VSUBS 0.006602f
C201 B.n161 VSUBS 0.006602f
C202 B.n162 VSUBS 0.006602f
C203 B.n163 VSUBS 0.006602f
C204 B.n164 VSUBS 0.006602f
C205 B.n165 VSUBS 0.006602f
C206 B.n166 VSUBS 0.006602f
C207 B.n167 VSUBS 0.006602f
C208 B.n168 VSUBS 0.006602f
C209 B.n169 VSUBS 0.006602f
C210 B.n170 VSUBS 0.006602f
C211 B.n171 VSUBS 0.006602f
C212 B.n172 VSUBS 0.006602f
C213 B.n173 VSUBS 0.006602f
C214 B.n174 VSUBS 0.006602f
C215 B.n175 VSUBS 0.006602f
C216 B.n176 VSUBS 0.006602f
C217 B.n177 VSUBS 0.006602f
C218 B.n178 VSUBS 0.006602f
C219 B.n179 VSUBS 0.006214f
C220 B.n180 VSUBS 0.006602f
C221 B.n181 VSUBS 0.006602f
C222 B.n182 VSUBS 0.00369f
C223 B.n183 VSUBS 0.006602f
C224 B.n184 VSUBS 0.006602f
C225 B.n185 VSUBS 0.006602f
C226 B.n186 VSUBS 0.006602f
C227 B.n187 VSUBS 0.006602f
C228 B.n188 VSUBS 0.006602f
C229 B.n189 VSUBS 0.006602f
C230 B.n190 VSUBS 0.006602f
C231 B.n191 VSUBS 0.006602f
C232 B.n192 VSUBS 0.006602f
C233 B.n193 VSUBS 0.006602f
C234 B.n194 VSUBS 0.006602f
C235 B.n195 VSUBS 0.00369f
C236 B.n196 VSUBS 0.015297f
C237 B.n197 VSUBS 0.006214f
C238 B.n198 VSUBS 0.006602f
C239 B.n199 VSUBS 0.006602f
C240 B.n200 VSUBS 0.006602f
C241 B.n201 VSUBS 0.006602f
C242 B.n202 VSUBS 0.006602f
C243 B.n203 VSUBS 0.006602f
C244 B.n204 VSUBS 0.006602f
C245 B.n205 VSUBS 0.006602f
C246 B.n206 VSUBS 0.006602f
C247 B.n207 VSUBS 0.006602f
C248 B.n208 VSUBS 0.006602f
C249 B.n209 VSUBS 0.006602f
C250 B.n210 VSUBS 0.006602f
C251 B.n211 VSUBS 0.006602f
C252 B.n212 VSUBS 0.006602f
C253 B.n213 VSUBS 0.006602f
C254 B.n214 VSUBS 0.006602f
C255 B.n215 VSUBS 0.006602f
C256 B.n216 VSUBS 0.006602f
C257 B.n217 VSUBS 0.006602f
C258 B.n218 VSUBS 0.006602f
C259 B.n219 VSUBS 0.006602f
C260 B.n220 VSUBS 0.006602f
C261 B.n221 VSUBS 0.006602f
C262 B.n222 VSUBS 0.006602f
C263 B.n223 VSUBS 0.006602f
C264 B.n224 VSUBS 0.006602f
C265 B.n225 VSUBS 0.006602f
C266 B.n226 VSUBS 0.006602f
C267 B.n227 VSUBS 0.006602f
C268 B.n228 VSUBS 0.006602f
C269 B.n229 VSUBS 0.01535f
C270 B.n230 VSUBS 0.01436f
C271 B.n231 VSUBS 0.01436f
C272 B.n232 VSUBS 0.006602f
C273 B.n233 VSUBS 0.006602f
C274 B.n234 VSUBS 0.006602f
C275 B.n235 VSUBS 0.006602f
C276 B.n236 VSUBS 0.006602f
C277 B.n237 VSUBS 0.006602f
C278 B.n238 VSUBS 0.006602f
C279 B.n239 VSUBS 0.006602f
C280 B.n240 VSUBS 0.006602f
C281 B.n241 VSUBS 0.006602f
C282 B.n242 VSUBS 0.006602f
C283 B.n243 VSUBS 0.006602f
C284 B.n244 VSUBS 0.006602f
C285 B.n245 VSUBS 0.006602f
C286 B.n246 VSUBS 0.006602f
C287 B.n247 VSUBS 0.006602f
C288 B.n248 VSUBS 0.006602f
C289 B.n249 VSUBS 0.006602f
C290 B.n250 VSUBS 0.006602f
C291 B.n251 VSUBS 0.006602f
C292 B.n252 VSUBS 0.006602f
C293 B.n253 VSUBS 0.006602f
C294 B.n254 VSUBS 0.006602f
C295 B.n255 VSUBS 0.006602f
C296 B.n256 VSUBS 0.006602f
C297 B.n257 VSUBS 0.006602f
C298 B.n258 VSUBS 0.006602f
C299 B.n259 VSUBS 0.006602f
C300 B.n260 VSUBS 0.006602f
C301 B.n261 VSUBS 0.006602f
C302 B.n262 VSUBS 0.006602f
C303 B.n263 VSUBS 0.006602f
C304 B.n264 VSUBS 0.006602f
C305 B.n265 VSUBS 0.006602f
C306 B.n266 VSUBS 0.006602f
C307 B.n267 VSUBS 0.006602f
C308 B.n268 VSUBS 0.006602f
C309 B.n269 VSUBS 0.006602f
C310 B.n270 VSUBS 0.006602f
C311 B.n271 VSUBS 0.006602f
C312 B.n272 VSUBS 0.006602f
C313 B.n273 VSUBS 0.006602f
C314 B.n274 VSUBS 0.006602f
C315 B.n275 VSUBS 0.006602f
C316 B.n276 VSUBS 0.006602f
C317 B.n277 VSUBS 0.006602f
C318 B.n278 VSUBS 0.006602f
C319 B.n279 VSUBS 0.006602f
C320 B.n280 VSUBS 0.006602f
C321 B.n281 VSUBS 0.006602f
C322 B.n282 VSUBS 0.006602f
C323 B.n283 VSUBS 0.006602f
C324 B.n284 VSUBS 0.006602f
C325 B.n285 VSUBS 0.006602f
C326 B.n286 VSUBS 0.006602f
C327 B.n287 VSUBS 0.006602f
C328 B.n288 VSUBS 0.006602f
C329 B.n289 VSUBS 0.006602f
C330 B.n290 VSUBS 0.006602f
C331 B.n291 VSUBS 0.006602f
C332 B.n292 VSUBS 0.006602f
C333 B.n293 VSUBS 0.006602f
C334 B.n294 VSUBS 0.006602f
C335 B.n295 VSUBS 0.006602f
C336 B.n296 VSUBS 0.006602f
C337 B.n297 VSUBS 0.006602f
C338 B.n298 VSUBS 0.006602f
C339 B.n299 VSUBS 0.006602f
C340 B.n300 VSUBS 0.006602f
C341 B.n301 VSUBS 0.006602f
C342 B.n302 VSUBS 0.01436f
C343 B.n303 VSUBS 0.015189f
C344 B.n304 VSUBS 0.014522f
C345 B.n305 VSUBS 0.006602f
C346 B.n306 VSUBS 0.006602f
C347 B.n307 VSUBS 0.006602f
C348 B.n308 VSUBS 0.006602f
C349 B.n309 VSUBS 0.006602f
C350 B.n310 VSUBS 0.006602f
C351 B.n311 VSUBS 0.006602f
C352 B.n312 VSUBS 0.006602f
C353 B.n313 VSUBS 0.006602f
C354 B.n314 VSUBS 0.006602f
C355 B.n315 VSUBS 0.006602f
C356 B.n316 VSUBS 0.006602f
C357 B.n317 VSUBS 0.006602f
C358 B.n318 VSUBS 0.006602f
C359 B.n319 VSUBS 0.006602f
C360 B.n320 VSUBS 0.006602f
C361 B.n321 VSUBS 0.006602f
C362 B.n322 VSUBS 0.006602f
C363 B.n323 VSUBS 0.006602f
C364 B.n324 VSUBS 0.006602f
C365 B.n325 VSUBS 0.006602f
C366 B.n326 VSUBS 0.006602f
C367 B.n327 VSUBS 0.006602f
C368 B.n328 VSUBS 0.006602f
C369 B.n329 VSUBS 0.006602f
C370 B.n330 VSUBS 0.006602f
C371 B.n331 VSUBS 0.006602f
C372 B.n332 VSUBS 0.006602f
C373 B.n333 VSUBS 0.006602f
C374 B.n334 VSUBS 0.006602f
C375 B.n335 VSUBS 0.006214f
C376 B.n336 VSUBS 0.006602f
C377 B.n337 VSUBS 0.006602f
C378 B.n338 VSUBS 0.00369f
C379 B.n339 VSUBS 0.006602f
C380 B.n340 VSUBS 0.006602f
C381 B.n341 VSUBS 0.006602f
C382 B.n342 VSUBS 0.006602f
C383 B.n343 VSUBS 0.006602f
C384 B.n344 VSUBS 0.006602f
C385 B.n345 VSUBS 0.006602f
C386 B.n346 VSUBS 0.006602f
C387 B.n347 VSUBS 0.006602f
C388 B.n348 VSUBS 0.006602f
C389 B.n349 VSUBS 0.006602f
C390 B.n350 VSUBS 0.006602f
C391 B.n351 VSUBS 0.00369f
C392 B.n352 VSUBS 0.015297f
C393 B.n353 VSUBS 0.006214f
C394 B.n354 VSUBS 0.006602f
C395 B.n355 VSUBS 0.006602f
C396 B.n356 VSUBS 0.006602f
C397 B.n357 VSUBS 0.006602f
C398 B.n358 VSUBS 0.006602f
C399 B.n359 VSUBS 0.006602f
C400 B.n360 VSUBS 0.006602f
C401 B.n361 VSUBS 0.006602f
C402 B.n362 VSUBS 0.006602f
C403 B.n363 VSUBS 0.006602f
C404 B.n364 VSUBS 0.006602f
C405 B.n365 VSUBS 0.006602f
C406 B.n366 VSUBS 0.006602f
C407 B.n367 VSUBS 0.006602f
C408 B.n368 VSUBS 0.006602f
C409 B.n369 VSUBS 0.006602f
C410 B.n370 VSUBS 0.006602f
C411 B.n371 VSUBS 0.006602f
C412 B.n372 VSUBS 0.006602f
C413 B.n373 VSUBS 0.006602f
C414 B.n374 VSUBS 0.006602f
C415 B.n375 VSUBS 0.006602f
C416 B.n376 VSUBS 0.006602f
C417 B.n377 VSUBS 0.006602f
C418 B.n378 VSUBS 0.006602f
C419 B.n379 VSUBS 0.006602f
C420 B.n380 VSUBS 0.006602f
C421 B.n381 VSUBS 0.006602f
C422 B.n382 VSUBS 0.006602f
C423 B.n383 VSUBS 0.006602f
C424 B.n384 VSUBS 0.006602f
C425 B.n385 VSUBS 0.01535f
C426 B.n386 VSUBS 0.01436f
C427 B.n387 VSUBS 0.01436f
C428 B.n388 VSUBS 0.006602f
C429 B.n389 VSUBS 0.006602f
C430 B.n390 VSUBS 0.006602f
C431 B.n391 VSUBS 0.006602f
C432 B.n392 VSUBS 0.006602f
C433 B.n393 VSUBS 0.006602f
C434 B.n394 VSUBS 0.006602f
C435 B.n395 VSUBS 0.006602f
C436 B.n396 VSUBS 0.006602f
C437 B.n397 VSUBS 0.006602f
C438 B.n398 VSUBS 0.006602f
C439 B.n399 VSUBS 0.006602f
C440 B.n400 VSUBS 0.006602f
C441 B.n401 VSUBS 0.006602f
C442 B.n402 VSUBS 0.006602f
C443 B.n403 VSUBS 0.006602f
C444 B.n404 VSUBS 0.006602f
C445 B.n405 VSUBS 0.006602f
C446 B.n406 VSUBS 0.006602f
C447 B.n407 VSUBS 0.006602f
C448 B.n408 VSUBS 0.006602f
C449 B.n409 VSUBS 0.006602f
C450 B.n410 VSUBS 0.006602f
C451 B.n411 VSUBS 0.006602f
C452 B.n412 VSUBS 0.006602f
C453 B.n413 VSUBS 0.006602f
C454 B.n414 VSUBS 0.006602f
C455 B.n415 VSUBS 0.006602f
C456 B.n416 VSUBS 0.006602f
C457 B.n417 VSUBS 0.006602f
C458 B.n418 VSUBS 0.006602f
C459 B.n419 VSUBS 0.006602f
C460 B.n420 VSUBS 0.006602f
C461 B.n421 VSUBS 0.006602f
C462 B.n422 VSUBS 0.006602f
C463 B.n423 VSUBS 0.01495f
C464 VDD2.n0 VSUBS 0.025007f
C465 VDD2.n1 VSUBS 0.022583f
C466 VDD2.n2 VSUBS 0.012135f
C467 VDD2.n3 VSUBS 0.028683f
C468 VDD2.n4 VSUBS 0.012849f
C469 VDD2.n5 VSUBS 0.022583f
C470 VDD2.n6 VSUBS 0.012135f
C471 VDD2.n7 VSUBS 0.021512f
C472 VDD2.n8 VSUBS 0.01822f
C473 VDD2.t2 VSUBS 0.061998f
C474 VDD2.n9 VSUBS 0.095946f
C475 VDD2.n10 VSUBS 0.450505f
C476 VDD2.n11 VSUBS 0.012135f
C477 VDD2.n12 VSUBS 0.012849f
C478 VDD2.n13 VSUBS 0.028683f
C479 VDD2.n14 VSUBS 0.028683f
C480 VDD2.n15 VSUBS 0.012849f
C481 VDD2.n16 VSUBS 0.012135f
C482 VDD2.n17 VSUBS 0.022583f
C483 VDD2.n18 VSUBS 0.022583f
C484 VDD2.n19 VSUBS 0.012135f
C485 VDD2.n20 VSUBS 0.012849f
C486 VDD2.n21 VSUBS 0.028683f
C487 VDD2.n22 VSUBS 0.070095f
C488 VDD2.n23 VSUBS 0.012849f
C489 VDD2.n24 VSUBS 0.012135f
C490 VDD2.n25 VSUBS 0.054359f
C491 VDD2.n26 VSUBS 0.052601f
C492 VDD2.t0 VSUBS 0.095475f
C493 VDD2.t5 VSUBS 0.095475f
C494 VDD2.n27 VSUBS 0.614171f
C495 VDD2.n28 VSUBS 1.61085f
C496 VDD2.n29 VSUBS 0.025007f
C497 VDD2.n30 VSUBS 0.022583f
C498 VDD2.n31 VSUBS 0.012135f
C499 VDD2.n32 VSUBS 0.028683f
C500 VDD2.n33 VSUBS 0.012849f
C501 VDD2.n34 VSUBS 0.022583f
C502 VDD2.n35 VSUBS 0.012135f
C503 VDD2.n36 VSUBS 0.021512f
C504 VDD2.n37 VSUBS 0.01822f
C505 VDD2.t1 VSUBS 0.061998f
C506 VDD2.n38 VSUBS 0.095946f
C507 VDD2.n39 VSUBS 0.450505f
C508 VDD2.n40 VSUBS 0.012135f
C509 VDD2.n41 VSUBS 0.012849f
C510 VDD2.n42 VSUBS 0.028683f
C511 VDD2.n43 VSUBS 0.028683f
C512 VDD2.n44 VSUBS 0.012849f
C513 VDD2.n45 VSUBS 0.012135f
C514 VDD2.n46 VSUBS 0.022583f
C515 VDD2.n47 VSUBS 0.022583f
C516 VDD2.n48 VSUBS 0.012135f
C517 VDD2.n49 VSUBS 0.012849f
C518 VDD2.n50 VSUBS 0.028683f
C519 VDD2.n51 VSUBS 0.070095f
C520 VDD2.n52 VSUBS 0.012849f
C521 VDD2.n53 VSUBS 0.012135f
C522 VDD2.n54 VSUBS 0.054359f
C523 VDD2.n55 VSUBS 0.050921f
C524 VDD2.n56 VSUBS 1.44871f
C525 VDD2.t4 VSUBS 0.095475f
C526 VDD2.t3 VSUBS 0.095475f
C527 VDD2.n57 VSUBS 0.614152f
C528 VN.n0 VSUBS 0.308719f
C529 VN.t5 VSUBS 0.81635f
C530 VN.t3 VSUBS 0.958463f
C531 VN.n1 VSUBS 0.410833f
C532 VN.n2 VSUBS 0.431585f
C533 VN.n3 VSUBS 0.067267f
C534 VN.t0 VSUBS 0.905307f
C535 VN.n4 VSUBS 0.429336f
C536 VN.n5 VSUBS 0.053315f
C537 VN.n6 VSUBS 0.308719f
C538 VN.t1 VSUBS 0.81635f
C539 VN.t2 VSUBS 0.958463f
C540 VN.n7 VSUBS 0.410833f
C541 VN.n8 VSUBS 0.431585f
C542 VN.n9 VSUBS 0.067267f
C543 VN.t4 VSUBS 0.905307f
C544 VN.n10 VSUBS 0.429336f
C545 VN.n11 VSUBS 1.98749f
C546 VTAIL.t4 VSUBS 0.110149f
C547 VTAIL.t3 VSUBS 0.110149f
C548 VTAIL.n0 VSUBS 0.625502f
C549 VTAIL.n1 VSUBS 0.571071f
C550 VTAIL.n2 VSUBS 0.02885f
C551 VTAIL.n3 VSUBS 0.026054f
C552 VTAIL.n4 VSUBS 0.014f
C553 VTAIL.n5 VSUBS 0.033092f
C554 VTAIL.n6 VSUBS 0.014824f
C555 VTAIL.n7 VSUBS 0.026054f
C556 VTAIL.n8 VSUBS 0.014f
C557 VTAIL.n9 VSUBS 0.024819f
C558 VTAIL.n10 VSUBS 0.02102f
C559 VTAIL.t7 VSUBS 0.071527f
C560 VTAIL.n11 VSUBS 0.110692f
C561 VTAIL.n12 VSUBS 0.519747f
C562 VTAIL.n13 VSUBS 0.014f
C563 VTAIL.n14 VSUBS 0.014824f
C564 VTAIL.n15 VSUBS 0.033092f
C565 VTAIL.n16 VSUBS 0.033092f
C566 VTAIL.n17 VSUBS 0.014824f
C567 VTAIL.n18 VSUBS 0.014f
C568 VTAIL.n19 VSUBS 0.026054f
C569 VTAIL.n20 VSUBS 0.026054f
C570 VTAIL.n21 VSUBS 0.014f
C571 VTAIL.n22 VSUBS 0.014824f
C572 VTAIL.n23 VSUBS 0.033092f
C573 VTAIL.n24 VSUBS 0.080869f
C574 VTAIL.n25 VSUBS 0.014824f
C575 VTAIL.n26 VSUBS 0.014f
C576 VTAIL.n27 VSUBS 0.062714f
C577 VTAIL.n28 VSUBS 0.040777f
C578 VTAIL.n29 VSUBS 0.209656f
C579 VTAIL.t10 VSUBS 0.110149f
C580 VTAIL.t11 VSUBS 0.110149f
C581 VTAIL.n30 VSUBS 0.625502f
C582 VTAIL.n31 VSUBS 1.48768f
C583 VTAIL.t5 VSUBS 0.110149f
C584 VTAIL.t0 VSUBS 0.110149f
C585 VTAIL.n32 VSUBS 0.625507f
C586 VTAIL.n33 VSUBS 1.48767f
C587 VTAIL.n34 VSUBS 0.02885f
C588 VTAIL.n35 VSUBS 0.026054f
C589 VTAIL.n36 VSUBS 0.014f
C590 VTAIL.n37 VSUBS 0.033092f
C591 VTAIL.n38 VSUBS 0.014824f
C592 VTAIL.n39 VSUBS 0.026054f
C593 VTAIL.n40 VSUBS 0.014f
C594 VTAIL.n41 VSUBS 0.024819f
C595 VTAIL.n42 VSUBS 0.02102f
C596 VTAIL.t2 VSUBS 0.071527f
C597 VTAIL.n43 VSUBS 0.110692f
C598 VTAIL.n44 VSUBS 0.519747f
C599 VTAIL.n45 VSUBS 0.014f
C600 VTAIL.n46 VSUBS 0.014824f
C601 VTAIL.n47 VSUBS 0.033092f
C602 VTAIL.n48 VSUBS 0.033092f
C603 VTAIL.n49 VSUBS 0.014824f
C604 VTAIL.n50 VSUBS 0.014f
C605 VTAIL.n51 VSUBS 0.026054f
C606 VTAIL.n52 VSUBS 0.026054f
C607 VTAIL.n53 VSUBS 0.014f
C608 VTAIL.n54 VSUBS 0.014824f
C609 VTAIL.n55 VSUBS 0.033092f
C610 VTAIL.n56 VSUBS 0.080869f
C611 VTAIL.n57 VSUBS 0.014824f
C612 VTAIL.n58 VSUBS 0.014f
C613 VTAIL.n59 VSUBS 0.062714f
C614 VTAIL.n60 VSUBS 0.040777f
C615 VTAIL.n61 VSUBS 0.209656f
C616 VTAIL.t8 VSUBS 0.110149f
C617 VTAIL.t9 VSUBS 0.110149f
C618 VTAIL.n62 VSUBS 0.625507f
C619 VTAIL.n63 VSUBS 0.639459f
C620 VTAIL.n64 VSUBS 0.02885f
C621 VTAIL.n65 VSUBS 0.026054f
C622 VTAIL.n66 VSUBS 0.014f
C623 VTAIL.n67 VSUBS 0.033092f
C624 VTAIL.n68 VSUBS 0.014824f
C625 VTAIL.n69 VSUBS 0.026054f
C626 VTAIL.n70 VSUBS 0.014f
C627 VTAIL.n71 VSUBS 0.024819f
C628 VTAIL.n72 VSUBS 0.02102f
C629 VTAIL.t6 VSUBS 0.071527f
C630 VTAIL.n73 VSUBS 0.110692f
C631 VTAIL.n74 VSUBS 0.519747f
C632 VTAIL.n75 VSUBS 0.014f
C633 VTAIL.n76 VSUBS 0.014824f
C634 VTAIL.n77 VSUBS 0.033092f
C635 VTAIL.n78 VSUBS 0.033092f
C636 VTAIL.n79 VSUBS 0.014824f
C637 VTAIL.n80 VSUBS 0.014f
C638 VTAIL.n81 VSUBS 0.026054f
C639 VTAIL.n82 VSUBS 0.026054f
C640 VTAIL.n83 VSUBS 0.014f
C641 VTAIL.n84 VSUBS 0.014824f
C642 VTAIL.n85 VSUBS 0.033092f
C643 VTAIL.n86 VSUBS 0.080869f
C644 VTAIL.n87 VSUBS 0.014824f
C645 VTAIL.n88 VSUBS 0.014f
C646 VTAIL.n89 VSUBS 0.062714f
C647 VTAIL.n90 VSUBS 0.040777f
C648 VTAIL.n91 VSUBS 0.960168f
C649 VTAIL.n92 VSUBS 0.02885f
C650 VTAIL.n93 VSUBS 0.026054f
C651 VTAIL.n94 VSUBS 0.014f
C652 VTAIL.n95 VSUBS 0.033092f
C653 VTAIL.n96 VSUBS 0.014824f
C654 VTAIL.n97 VSUBS 0.026054f
C655 VTAIL.n98 VSUBS 0.014f
C656 VTAIL.n99 VSUBS 0.024819f
C657 VTAIL.n100 VSUBS 0.02102f
C658 VTAIL.t1 VSUBS 0.071527f
C659 VTAIL.n101 VSUBS 0.110692f
C660 VTAIL.n102 VSUBS 0.519747f
C661 VTAIL.n103 VSUBS 0.014f
C662 VTAIL.n104 VSUBS 0.014824f
C663 VTAIL.n105 VSUBS 0.033092f
C664 VTAIL.n106 VSUBS 0.033092f
C665 VTAIL.n107 VSUBS 0.014824f
C666 VTAIL.n108 VSUBS 0.014f
C667 VTAIL.n109 VSUBS 0.026054f
C668 VTAIL.n110 VSUBS 0.026054f
C669 VTAIL.n111 VSUBS 0.014f
C670 VTAIL.n112 VSUBS 0.014824f
C671 VTAIL.n113 VSUBS 0.033092f
C672 VTAIL.n114 VSUBS 0.080869f
C673 VTAIL.n115 VSUBS 0.014824f
C674 VTAIL.n116 VSUBS 0.014f
C675 VTAIL.n117 VSUBS 0.062714f
C676 VTAIL.n118 VSUBS 0.040777f
C677 VTAIL.n119 VSUBS 0.930857f
C678 VDD1.n0 VSUBS 0.025386f
C679 VDD1.n1 VSUBS 0.022926f
C680 VDD1.n2 VSUBS 0.012319f
C681 VDD1.n3 VSUBS 0.029118f
C682 VDD1.n4 VSUBS 0.013044f
C683 VDD1.n5 VSUBS 0.022926f
C684 VDD1.n6 VSUBS 0.012319f
C685 VDD1.n7 VSUBS 0.021839f
C686 VDD1.n8 VSUBS 0.018496f
C687 VDD1.t1 VSUBS 0.062939f
C688 VDD1.n9 VSUBS 0.097401f
C689 VDD1.n10 VSUBS 0.457341f
C690 VDD1.n11 VSUBS 0.012319f
C691 VDD1.n12 VSUBS 0.013044f
C692 VDD1.n13 VSUBS 0.029118f
C693 VDD1.n14 VSUBS 0.029118f
C694 VDD1.n15 VSUBS 0.013044f
C695 VDD1.n16 VSUBS 0.012319f
C696 VDD1.n17 VSUBS 0.022926f
C697 VDD1.n18 VSUBS 0.022926f
C698 VDD1.n19 VSUBS 0.012319f
C699 VDD1.n20 VSUBS 0.013044f
C700 VDD1.n21 VSUBS 0.029118f
C701 VDD1.n22 VSUBS 0.071159f
C702 VDD1.n23 VSUBS 0.013044f
C703 VDD1.n24 VSUBS 0.012319f
C704 VDD1.n25 VSUBS 0.055184f
C705 VDD1.n26 VSUBS 0.053772f
C706 VDD1.n27 VSUBS 0.025386f
C707 VDD1.n28 VSUBS 0.022926f
C708 VDD1.n29 VSUBS 0.012319f
C709 VDD1.n30 VSUBS 0.029118f
C710 VDD1.n31 VSUBS 0.013044f
C711 VDD1.n32 VSUBS 0.022926f
C712 VDD1.n33 VSUBS 0.012319f
C713 VDD1.n34 VSUBS 0.021839f
C714 VDD1.n35 VSUBS 0.018496f
C715 VDD1.t5 VSUBS 0.062939f
C716 VDD1.n36 VSUBS 0.097401f
C717 VDD1.n37 VSUBS 0.457341f
C718 VDD1.n38 VSUBS 0.012319f
C719 VDD1.n39 VSUBS 0.013044f
C720 VDD1.n40 VSUBS 0.029118f
C721 VDD1.n41 VSUBS 0.029118f
C722 VDD1.n42 VSUBS 0.013044f
C723 VDD1.n43 VSUBS 0.012319f
C724 VDD1.n44 VSUBS 0.022926f
C725 VDD1.n45 VSUBS 0.022926f
C726 VDD1.n46 VSUBS 0.012319f
C727 VDD1.n47 VSUBS 0.013044f
C728 VDD1.n48 VSUBS 0.029118f
C729 VDD1.n49 VSUBS 0.071159f
C730 VDD1.n50 VSUBS 0.013044f
C731 VDD1.n51 VSUBS 0.012319f
C732 VDD1.n52 VSUBS 0.055184f
C733 VDD1.n53 VSUBS 0.053399f
C734 VDD1.t0 VSUBS 0.096924f
C735 VDD1.t4 VSUBS 0.096924f
C736 VDD1.n54 VSUBS 0.623491f
C737 VDD1.n55 VSUBS 1.70957f
C738 VDD1.t3 VSUBS 0.096924f
C739 VDD1.t2 VSUBS 0.096924f
C740 VDD1.n56 VSUBS 0.622364f
C741 VDD1.n57 VSUBS 1.83753f
C742 VP.n0 VSUBS 0.078852f
C743 VP.t0 VSUBS 0.847401f
C744 VP.n1 VSUBS 0.069826f
C745 VP.n2 VSUBS 0.320462f
C746 VP.t5 VSUBS 0.939743f
C747 VP.t2 VSUBS 0.847401f
C748 VP.t3 VSUBS 0.994919f
C749 VP.n3 VSUBS 0.426459f
C750 VP.n4 VSUBS 0.448001f
C751 VP.n5 VSUBS 0.069826f
C752 VP.n6 VSUBS 0.445666f
C753 VP.n7 VSUBS 2.02924f
C754 VP.t1 VSUBS 0.939743f
C755 VP.n8 VSUBS 0.445666f
C756 VP.n9 VSUBS 2.08581f
C757 VP.n10 VSUBS 0.078852f
C758 VP.n11 VSUBS 0.059093f
C759 VP.n12 VSUBS 0.411369f
C760 VP.n13 VSUBS 0.069826f
C761 VP.t4 VSUBS 0.939743f
C762 VP.n14 VSUBS 0.445666f
C763 VP.n15 VSUBS 0.055342f
.ends

