* NGSPICE file created from diff_pair_sample_0070.ext - technology: sky130A

.subckt diff_pair_sample_0070 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t9 w_n3170_n1092# sky130_fd_pr__pfet_01v8 ad=0.2418 pd=2.02 as=0.1023 ps=0.95 w=0.62 l=2.42
X1 B.t11 B.t9 B.t10 w_n3170_n1092# sky130_fd_pr__pfet_01v8 ad=0.2418 pd=2.02 as=0 ps=0 w=0.62 l=2.42
X2 VTAIL.t6 VP.t1 VDD1.t4 w_n3170_n1092# sky130_fd_pr__pfet_01v8 ad=0.1023 pd=0.95 as=0.1023 ps=0.95 w=0.62 l=2.42
X3 VDD2.t5 VN.t0 VTAIL.t3 w_n3170_n1092# sky130_fd_pr__pfet_01v8 ad=0.2418 pd=2.02 as=0.1023 ps=0.95 w=0.62 l=2.42
X4 VTAIL.t5 VN.t1 VDD2.t4 w_n3170_n1092# sky130_fd_pr__pfet_01v8 ad=0.1023 pd=0.95 as=0.1023 ps=0.95 w=0.62 l=2.42
X5 VDD2.t3 VN.t2 VTAIL.t1 w_n3170_n1092# sky130_fd_pr__pfet_01v8 ad=0.1023 pd=0.95 as=0.2418 ps=2.02 w=0.62 l=2.42
X6 VDD2.t2 VN.t3 VTAIL.t2 w_n3170_n1092# sky130_fd_pr__pfet_01v8 ad=0.1023 pd=0.95 as=0.2418 ps=2.02 w=0.62 l=2.42
X7 B.t8 B.t6 B.t7 w_n3170_n1092# sky130_fd_pr__pfet_01v8 ad=0.2418 pd=2.02 as=0 ps=0 w=0.62 l=2.42
X8 VDD1.t3 VP.t2 VTAIL.t11 w_n3170_n1092# sky130_fd_pr__pfet_01v8 ad=0.1023 pd=0.95 as=0.2418 ps=2.02 w=0.62 l=2.42
X9 B.t5 B.t3 B.t4 w_n3170_n1092# sky130_fd_pr__pfet_01v8 ad=0.2418 pd=2.02 as=0 ps=0 w=0.62 l=2.42
X10 VTAIL.t4 VN.t4 VDD2.t1 w_n3170_n1092# sky130_fd_pr__pfet_01v8 ad=0.1023 pd=0.95 as=0.1023 ps=0.95 w=0.62 l=2.42
X11 VDD1.t2 VP.t3 VTAIL.t8 w_n3170_n1092# sky130_fd_pr__pfet_01v8 ad=0.1023 pd=0.95 as=0.2418 ps=2.02 w=0.62 l=2.42
X12 VTAIL.t7 VP.t4 VDD1.t1 w_n3170_n1092# sky130_fd_pr__pfet_01v8 ad=0.1023 pd=0.95 as=0.1023 ps=0.95 w=0.62 l=2.42
X13 VDD1.t0 VP.t5 VTAIL.t10 w_n3170_n1092# sky130_fd_pr__pfet_01v8 ad=0.2418 pd=2.02 as=0.1023 ps=0.95 w=0.62 l=2.42
X14 B.t2 B.t0 B.t1 w_n3170_n1092# sky130_fd_pr__pfet_01v8 ad=0.2418 pd=2.02 as=0 ps=0 w=0.62 l=2.42
X15 VDD2.t0 VN.t5 VTAIL.t0 w_n3170_n1092# sky130_fd_pr__pfet_01v8 ad=0.2418 pd=2.02 as=0.1023 ps=0.95 w=0.62 l=2.42
R0 VP.n11 VP.n8 161.3
R1 VP.n13 VP.n12 161.3
R2 VP.n14 VP.n7 161.3
R3 VP.n16 VP.n15 161.3
R4 VP.n17 VP.n6 161.3
R5 VP.n37 VP.n0 161.3
R6 VP.n36 VP.n35 161.3
R7 VP.n34 VP.n1 161.3
R8 VP.n33 VP.n32 161.3
R9 VP.n31 VP.n2 161.3
R10 VP.n30 VP.n29 161.3
R11 VP.n28 VP.n3 161.3
R12 VP.n27 VP.n26 161.3
R13 VP.n25 VP.n4 161.3
R14 VP.n24 VP.n23 161.3
R15 VP.n22 VP.n5 161.3
R16 VP.n21 VP.n20 98.4345
R17 VP.n39 VP.n38 98.4345
R18 VP.n19 VP.n18 98.4345
R19 VP.n26 VP.n25 52.5823
R20 VP.n32 VP.n1 52.5823
R21 VP.n12 VP.n7 52.5823
R22 VP.n10 VP.n9 47.9004
R23 VP.n9 VP.t0 40.4735
R24 VP.n21 VP.n19 39.3594
R25 VP.n25 VP.n24 28.2389
R26 VP.n36 VP.n1 28.2389
R27 VP.n16 VP.n7 28.2389
R28 VP.n24 VP.n5 24.3439
R29 VP.n26 VP.n3 24.3439
R30 VP.n30 VP.n3 24.3439
R31 VP.n31 VP.n30 24.3439
R32 VP.n32 VP.n31 24.3439
R33 VP.n37 VP.n36 24.3439
R34 VP.n17 VP.n16 24.3439
R35 VP.n11 VP.n10 24.3439
R36 VP.n12 VP.n11 24.3439
R37 VP.n20 VP.n5 12.1722
R38 VP.n38 VP.n37 12.1722
R39 VP.n18 VP.n17 12.1722
R40 VP.n9 VP.n8 6.7099
R41 VP.n30 VP.t4 6.17488
R42 VP.n20 VP.t5 6.17488
R43 VP.n38 VP.t2 6.17488
R44 VP.n10 VP.t1 6.17488
R45 VP.n18 VP.t3 6.17488
R46 VP.n19 VP.n6 0.278398
R47 VP.n22 VP.n21 0.278398
R48 VP.n39 VP.n0 0.278398
R49 VP.n13 VP.n8 0.189894
R50 VP.n14 VP.n13 0.189894
R51 VP.n15 VP.n14 0.189894
R52 VP.n15 VP.n6 0.189894
R53 VP.n23 VP.n22 0.189894
R54 VP.n23 VP.n4 0.189894
R55 VP.n27 VP.n4 0.189894
R56 VP.n28 VP.n27 0.189894
R57 VP.n29 VP.n28 0.189894
R58 VP.n29 VP.n2 0.189894
R59 VP.n33 VP.n2 0.189894
R60 VP.n34 VP.n33 0.189894
R61 VP.n35 VP.n34 0.189894
R62 VP.n35 VP.n0 0.189894
R63 VP VP.n39 0.153422
R64 VTAIL.n11 VTAIL.t1 670
R65 VTAIL.n2 VTAIL.t11 670
R66 VTAIL.n10 VTAIL.t8 670
R67 VTAIL.n7 VTAIL.t2 670
R68 VTAIL.n1 VTAIL.n0 617.573
R69 VTAIL.n4 VTAIL.n3 617.573
R70 VTAIL.n9 VTAIL.n8 617.573
R71 VTAIL.n6 VTAIL.n5 617.573
R72 VTAIL.n0 VTAIL.t0 52.4279
R73 VTAIL.n0 VTAIL.t5 52.4279
R74 VTAIL.n3 VTAIL.t10 52.4279
R75 VTAIL.n3 VTAIL.t7 52.4279
R76 VTAIL.n8 VTAIL.t9 52.4279
R77 VTAIL.n8 VTAIL.t6 52.4279
R78 VTAIL.n5 VTAIL.t3 52.4279
R79 VTAIL.n5 VTAIL.t4 52.4279
R80 VTAIL.n6 VTAIL.n4 17.6427
R81 VTAIL.n11 VTAIL.n10 15.2721
R82 VTAIL.n7 VTAIL.n6 2.37119
R83 VTAIL.n10 VTAIL.n9 2.37119
R84 VTAIL.n4 VTAIL.n2 2.37119
R85 VTAIL VTAIL.n11 1.72033
R86 VTAIL.n9 VTAIL.n7 1.65567
R87 VTAIL.n2 VTAIL.n1 1.65567
R88 VTAIL VTAIL.n1 0.651362
R89 VDD1 VDD1.t5 688.515
R90 VDD1.n1 VDD1.t0 688.403
R91 VDD1.n1 VDD1.n0 634.789
R92 VDD1.n3 VDD1.n2 634.253
R93 VDD1.n2 VDD1.t4 52.4279
R94 VDD1.n2 VDD1.t2 52.4279
R95 VDD1.n0 VDD1.t1 52.4279
R96 VDD1.n0 VDD1.t3 52.4279
R97 VDD1.n3 VDD1.n1 33.7229
R98 VDD1 VDD1.n3 0.534983
R99 B.n90 B.t10 712.482
R100 B.n200 B.t7 712.482
R101 B.n34 B.t5 712.482
R102 B.n26 B.t2 712.482
R103 B.n91 B.t11 659.149
R104 B.n201 B.t8 659.149
R105 B.n35 B.t4 659.149
R106 B.n27 B.t1 659.149
R107 B.n216 B.n215 585
R108 B.n214 B.n81 585
R109 B.n213 B.n212 585
R110 B.n211 B.n82 585
R111 B.n210 B.n209 585
R112 B.n208 B.n83 585
R113 B.n207 B.n206 585
R114 B.n205 B.n84 585
R115 B.n204 B.n203 585
R116 B.n199 B.n85 585
R117 B.n198 B.n197 585
R118 B.n196 B.n86 585
R119 B.n195 B.n194 585
R120 B.n193 B.n87 585
R121 B.n192 B.n191 585
R122 B.n190 B.n88 585
R123 B.n189 B.n188 585
R124 B.n187 B.n89 585
R125 B.n185 B.n184 585
R126 B.n183 B.n92 585
R127 B.n182 B.n181 585
R128 B.n180 B.n93 585
R129 B.n179 B.n178 585
R130 B.n177 B.n94 585
R131 B.n176 B.n175 585
R132 B.n174 B.n95 585
R133 B.n217 B.n80 585
R134 B.n219 B.n218 585
R135 B.n220 B.n79 585
R136 B.n222 B.n221 585
R137 B.n223 B.n78 585
R138 B.n225 B.n224 585
R139 B.n226 B.n77 585
R140 B.n228 B.n227 585
R141 B.n229 B.n76 585
R142 B.n231 B.n230 585
R143 B.n232 B.n75 585
R144 B.n234 B.n233 585
R145 B.n235 B.n74 585
R146 B.n237 B.n236 585
R147 B.n238 B.n73 585
R148 B.n240 B.n239 585
R149 B.n241 B.n72 585
R150 B.n243 B.n242 585
R151 B.n244 B.n71 585
R152 B.n246 B.n245 585
R153 B.n247 B.n70 585
R154 B.n249 B.n248 585
R155 B.n250 B.n69 585
R156 B.n252 B.n251 585
R157 B.n253 B.n68 585
R158 B.n255 B.n254 585
R159 B.n256 B.n67 585
R160 B.n258 B.n257 585
R161 B.n259 B.n66 585
R162 B.n261 B.n260 585
R163 B.n262 B.n65 585
R164 B.n264 B.n263 585
R165 B.n265 B.n64 585
R166 B.n267 B.n266 585
R167 B.n268 B.n63 585
R168 B.n270 B.n269 585
R169 B.n271 B.n62 585
R170 B.n273 B.n272 585
R171 B.n274 B.n61 585
R172 B.n276 B.n275 585
R173 B.n277 B.n60 585
R174 B.n279 B.n278 585
R175 B.n280 B.n59 585
R176 B.n282 B.n281 585
R177 B.n283 B.n58 585
R178 B.n285 B.n284 585
R179 B.n286 B.n57 585
R180 B.n288 B.n287 585
R181 B.n289 B.n56 585
R182 B.n291 B.n290 585
R183 B.n292 B.n55 585
R184 B.n294 B.n293 585
R185 B.n295 B.n54 585
R186 B.n297 B.n296 585
R187 B.n298 B.n53 585
R188 B.n300 B.n299 585
R189 B.n301 B.n52 585
R190 B.n303 B.n302 585
R191 B.n304 B.n51 585
R192 B.n306 B.n305 585
R193 B.n307 B.n50 585
R194 B.n309 B.n308 585
R195 B.n310 B.n49 585
R196 B.n312 B.n311 585
R197 B.n313 B.n48 585
R198 B.n315 B.n314 585
R199 B.n316 B.n47 585
R200 B.n318 B.n317 585
R201 B.n319 B.n46 585
R202 B.n321 B.n320 585
R203 B.n322 B.n45 585
R204 B.n324 B.n323 585
R205 B.n325 B.n44 585
R206 B.n327 B.n326 585
R207 B.n328 B.n43 585
R208 B.n330 B.n329 585
R209 B.n331 B.n42 585
R210 B.n333 B.n332 585
R211 B.n334 B.n41 585
R212 B.n336 B.n335 585
R213 B.n337 B.n40 585
R214 B.n339 B.n338 585
R215 B.n379 B.n22 585
R216 B.n378 B.n377 585
R217 B.n376 B.n23 585
R218 B.n375 B.n374 585
R219 B.n373 B.n24 585
R220 B.n372 B.n371 585
R221 B.n370 B.n25 585
R222 B.n369 B.n368 585
R223 B.n367 B.n366 585
R224 B.n365 B.n29 585
R225 B.n364 B.n363 585
R226 B.n362 B.n30 585
R227 B.n361 B.n360 585
R228 B.n359 B.n31 585
R229 B.n358 B.n357 585
R230 B.n356 B.n32 585
R231 B.n355 B.n354 585
R232 B.n353 B.n33 585
R233 B.n351 B.n350 585
R234 B.n349 B.n36 585
R235 B.n348 B.n347 585
R236 B.n346 B.n37 585
R237 B.n345 B.n344 585
R238 B.n343 B.n38 585
R239 B.n342 B.n341 585
R240 B.n340 B.n39 585
R241 B.n381 B.n380 585
R242 B.n382 B.n21 585
R243 B.n384 B.n383 585
R244 B.n385 B.n20 585
R245 B.n387 B.n386 585
R246 B.n388 B.n19 585
R247 B.n390 B.n389 585
R248 B.n391 B.n18 585
R249 B.n393 B.n392 585
R250 B.n394 B.n17 585
R251 B.n396 B.n395 585
R252 B.n397 B.n16 585
R253 B.n399 B.n398 585
R254 B.n400 B.n15 585
R255 B.n402 B.n401 585
R256 B.n403 B.n14 585
R257 B.n405 B.n404 585
R258 B.n406 B.n13 585
R259 B.n408 B.n407 585
R260 B.n409 B.n12 585
R261 B.n411 B.n410 585
R262 B.n412 B.n11 585
R263 B.n414 B.n413 585
R264 B.n415 B.n10 585
R265 B.n417 B.n416 585
R266 B.n418 B.n9 585
R267 B.n420 B.n419 585
R268 B.n421 B.n8 585
R269 B.n423 B.n422 585
R270 B.n424 B.n7 585
R271 B.n426 B.n425 585
R272 B.n427 B.n6 585
R273 B.n429 B.n428 585
R274 B.n430 B.n5 585
R275 B.n432 B.n431 585
R276 B.n433 B.n4 585
R277 B.n435 B.n434 585
R278 B.n436 B.n3 585
R279 B.n438 B.n437 585
R280 B.n439 B.n0 585
R281 B.n2 B.n1 585
R282 B.n116 B.n115 585
R283 B.n117 B.n114 585
R284 B.n119 B.n118 585
R285 B.n120 B.n113 585
R286 B.n122 B.n121 585
R287 B.n123 B.n112 585
R288 B.n125 B.n124 585
R289 B.n126 B.n111 585
R290 B.n128 B.n127 585
R291 B.n129 B.n110 585
R292 B.n131 B.n130 585
R293 B.n132 B.n109 585
R294 B.n134 B.n133 585
R295 B.n135 B.n108 585
R296 B.n137 B.n136 585
R297 B.n138 B.n107 585
R298 B.n140 B.n139 585
R299 B.n141 B.n106 585
R300 B.n143 B.n142 585
R301 B.n144 B.n105 585
R302 B.n146 B.n145 585
R303 B.n147 B.n104 585
R304 B.n149 B.n148 585
R305 B.n150 B.n103 585
R306 B.n152 B.n151 585
R307 B.n153 B.n102 585
R308 B.n155 B.n154 585
R309 B.n156 B.n101 585
R310 B.n158 B.n157 585
R311 B.n159 B.n100 585
R312 B.n161 B.n160 585
R313 B.n162 B.n99 585
R314 B.n164 B.n163 585
R315 B.n165 B.n98 585
R316 B.n167 B.n166 585
R317 B.n168 B.n97 585
R318 B.n170 B.n169 585
R319 B.n171 B.n96 585
R320 B.n173 B.n172 585
R321 B.n172 B.n95 482.89
R322 B.n217 B.n216 482.89
R323 B.n338 B.n39 482.89
R324 B.n380 B.n379 482.89
R325 B.n441 B.n440 256.663
R326 B.n440 B.n439 235.042
R327 B.n440 B.n2 235.042
R328 B.n90 B.t9 209.119
R329 B.n200 B.t6 209.119
R330 B.n34 B.t3 209.119
R331 B.n26 B.t0 209.119
R332 B.n176 B.n95 163.367
R333 B.n177 B.n176 163.367
R334 B.n178 B.n177 163.367
R335 B.n178 B.n93 163.367
R336 B.n182 B.n93 163.367
R337 B.n183 B.n182 163.367
R338 B.n184 B.n183 163.367
R339 B.n184 B.n89 163.367
R340 B.n189 B.n89 163.367
R341 B.n190 B.n189 163.367
R342 B.n191 B.n190 163.367
R343 B.n191 B.n87 163.367
R344 B.n195 B.n87 163.367
R345 B.n196 B.n195 163.367
R346 B.n197 B.n196 163.367
R347 B.n197 B.n85 163.367
R348 B.n204 B.n85 163.367
R349 B.n205 B.n204 163.367
R350 B.n206 B.n205 163.367
R351 B.n206 B.n83 163.367
R352 B.n210 B.n83 163.367
R353 B.n211 B.n210 163.367
R354 B.n212 B.n211 163.367
R355 B.n212 B.n81 163.367
R356 B.n216 B.n81 163.367
R357 B.n338 B.n337 163.367
R358 B.n337 B.n336 163.367
R359 B.n336 B.n41 163.367
R360 B.n332 B.n41 163.367
R361 B.n332 B.n331 163.367
R362 B.n331 B.n330 163.367
R363 B.n330 B.n43 163.367
R364 B.n326 B.n43 163.367
R365 B.n326 B.n325 163.367
R366 B.n325 B.n324 163.367
R367 B.n324 B.n45 163.367
R368 B.n320 B.n45 163.367
R369 B.n320 B.n319 163.367
R370 B.n319 B.n318 163.367
R371 B.n318 B.n47 163.367
R372 B.n314 B.n47 163.367
R373 B.n314 B.n313 163.367
R374 B.n313 B.n312 163.367
R375 B.n312 B.n49 163.367
R376 B.n308 B.n49 163.367
R377 B.n308 B.n307 163.367
R378 B.n307 B.n306 163.367
R379 B.n306 B.n51 163.367
R380 B.n302 B.n51 163.367
R381 B.n302 B.n301 163.367
R382 B.n301 B.n300 163.367
R383 B.n300 B.n53 163.367
R384 B.n296 B.n53 163.367
R385 B.n296 B.n295 163.367
R386 B.n295 B.n294 163.367
R387 B.n294 B.n55 163.367
R388 B.n290 B.n55 163.367
R389 B.n290 B.n289 163.367
R390 B.n289 B.n288 163.367
R391 B.n288 B.n57 163.367
R392 B.n284 B.n57 163.367
R393 B.n284 B.n283 163.367
R394 B.n283 B.n282 163.367
R395 B.n282 B.n59 163.367
R396 B.n278 B.n59 163.367
R397 B.n278 B.n277 163.367
R398 B.n277 B.n276 163.367
R399 B.n276 B.n61 163.367
R400 B.n272 B.n61 163.367
R401 B.n272 B.n271 163.367
R402 B.n271 B.n270 163.367
R403 B.n270 B.n63 163.367
R404 B.n266 B.n63 163.367
R405 B.n266 B.n265 163.367
R406 B.n265 B.n264 163.367
R407 B.n264 B.n65 163.367
R408 B.n260 B.n65 163.367
R409 B.n260 B.n259 163.367
R410 B.n259 B.n258 163.367
R411 B.n258 B.n67 163.367
R412 B.n254 B.n67 163.367
R413 B.n254 B.n253 163.367
R414 B.n253 B.n252 163.367
R415 B.n252 B.n69 163.367
R416 B.n248 B.n69 163.367
R417 B.n248 B.n247 163.367
R418 B.n247 B.n246 163.367
R419 B.n246 B.n71 163.367
R420 B.n242 B.n71 163.367
R421 B.n242 B.n241 163.367
R422 B.n241 B.n240 163.367
R423 B.n240 B.n73 163.367
R424 B.n236 B.n73 163.367
R425 B.n236 B.n235 163.367
R426 B.n235 B.n234 163.367
R427 B.n234 B.n75 163.367
R428 B.n230 B.n75 163.367
R429 B.n230 B.n229 163.367
R430 B.n229 B.n228 163.367
R431 B.n228 B.n77 163.367
R432 B.n224 B.n77 163.367
R433 B.n224 B.n223 163.367
R434 B.n223 B.n222 163.367
R435 B.n222 B.n79 163.367
R436 B.n218 B.n79 163.367
R437 B.n218 B.n217 163.367
R438 B.n379 B.n378 163.367
R439 B.n378 B.n23 163.367
R440 B.n374 B.n23 163.367
R441 B.n374 B.n373 163.367
R442 B.n373 B.n372 163.367
R443 B.n372 B.n25 163.367
R444 B.n368 B.n25 163.367
R445 B.n368 B.n367 163.367
R446 B.n367 B.n29 163.367
R447 B.n363 B.n29 163.367
R448 B.n363 B.n362 163.367
R449 B.n362 B.n361 163.367
R450 B.n361 B.n31 163.367
R451 B.n357 B.n31 163.367
R452 B.n357 B.n356 163.367
R453 B.n356 B.n355 163.367
R454 B.n355 B.n33 163.367
R455 B.n350 B.n33 163.367
R456 B.n350 B.n349 163.367
R457 B.n349 B.n348 163.367
R458 B.n348 B.n37 163.367
R459 B.n344 B.n37 163.367
R460 B.n344 B.n343 163.367
R461 B.n343 B.n342 163.367
R462 B.n342 B.n39 163.367
R463 B.n380 B.n21 163.367
R464 B.n384 B.n21 163.367
R465 B.n385 B.n384 163.367
R466 B.n386 B.n385 163.367
R467 B.n386 B.n19 163.367
R468 B.n390 B.n19 163.367
R469 B.n391 B.n390 163.367
R470 B.n392 B.n391 163.367
R471 B.n392 B.n17 163.367
R472 B.n396 B.n17 163.367
R473 B.n397 B.n396 163.367
R474 B.n398 B.n397 163.367
R475 B.n398 B.n15 163.367
R476 B.n402 B.n15 163.367
R477 B.n403 B.n402 163.367
R478 B.n404 B.n403 163.367
R479 B.n404 B.n13 163.367
R480 B.n408 B.n13 163.367
R481 B.n409 B.n408 163.367
R482 B.n410 B.n409 163.367
R483 B.n410 B.n11 163.367
R484 B.n414 B.n11 163.367
R485 B.n415 B.n414 163.367
R486 B.n416 B.n415 163.367
R487 B.n416 B.n9 163.367
R488 B.n420 B.n9 163.367
R489 B.n421 B.n420 163.367
R490 B.n422 B.n421 163.367
R491 B.n422 B.n7 163.367
R492 B.n426 B.n7 163.367
R493 B.n427 B.n426 163.367
R494 B.n428 B.n427 163.367
R495 B.n428 B.n5 163.367
R496 B.n432 B.n5 163.367
R497 B.n433 B.n432 163.367
R498 B.n434 B.n433 163.367
R499 B.n434 B.n3 163.367
R500 B.n438 B.n3 163.367
R501 B.n439 B.n438 163.367
R502 B.n116 B.n2 163.367
R503 B.n117 B.n116 163.367
R504 B.n118 B.n117 163.367
R505 B.n118 B.n113 163.367
R506 B.n122 B.n113 163.367
R507 B.n123 B.n122 163.367
R508 B.n124 B.n123 163.367
R509 B.n124 B.n111 163.367
R510 B.n128 B.n111 163.367
R511 B.n129 B.n128 163.367
R512 B.n130 B.n129 163.367
R513 B.n130 B.n109 163.367
R514 B.n134 B.n109 163.367
R515 B.n135 B.n134 163.367
R516 B.n136 B.n135 163.367
R517 B.n136 B.n107 163.367
R518 B.n140 B.n107 163.367
R519 B.n141 B.n140 163.367
R520 B.n142 B.n141 163.367
R521 B.n142 B.n105 163.367
R522 B.n146 B.n105 163.367
R523 B.n147 B.n146 163.367
R524 B.n148 B.n147 163.367
R525 B.n148 B.n103 163.367
R526 B.n152 B.n103 163.367
R527 B.n153 B.n152 163.367
R528 B.n154 B.n153 163.367
R529 B.n154 B.n101 163.367
R530 B.n158 B.n101 163.367
R531 B.n159 B.n158 163.367
R532 B.n160 B.n159 163.367
R533 B.n160 B.n99 163.367
R534 B.n164 B.n99 163.367
R535 B.n165 B.n164 163.367
R536 B.n166 B.n165 163.367
R537 B.n166 B.n97 163.367
R538 B.n170 B.n97 163.367
R539 B.n171 B.n170 163.367
R540 B.n172 B.n171 163.367
R541 B.n186 B.n91 59.5399
R542 B.n202 B.n201 59.5399
R543 B.n352 B.n35 59.5399
R544 B.n28 B.n27 59.5399
R545 B.n91 B.n90 53.3338
R546 B.n201 B.n200 53.3338
R547 B.n35 B.n34 53.3338
R548 B.n27 B.n26 53.3338
R549 B.n381 B.n22 31.3761
R550 B.n340 B.n339 31.3761
R551 B.n215 B.n80 31.3761
R552 B.n174 B.n173 31.3761
R553 B B.n441 18.0485
R554 B.n382 B.n381 10.6151
R555 B.n383 B.n382 10.6151
R556 B.n383 B.n20 10.6151
R557 B.n387 B.n20 10.6151
R558 B.n388 B.n387 10.6151
R559 B.n389 B.n388 10.6151
R560 B.n389 B.n18 10.6151
R561 B.n393 B.n18 10.6151
R562 B.n394 B.n393 10.6151
R563 B.n395 B.n394 10.6151
R564 B.n395 B.n16 10.6151
R565 B.n399 B.n16 10.6151
R566 B.n400 B.n399 10.6151
R567 B.n401 B.n400 10.6151
R568 B.n401 B.n14 10.6151
R569 B.n405 B.n14 10.6151
R570 B.n406 B.n405 10.6151
R571 B.n407 B.n406 10.6151
R572 B.n407 B.n12 10.6151
R573 B.n411 B.n12 10.6151
R574 B.n412 B.n411 10.6151
R575 B.n413 B.n412 10.6151
R576 B.n413 B.n10 10.6151
R577 B.n417 B.n10 10.6151
R578 B.n418 B.n417 10.6151
R579 B.n419 B.n418 10.6151
R580 B.n419 B.n8 10.6151
R581 B.n423 B.n8 10.6151
R582 B.n424 B.n423 10.6151
R583 B.n425 B.n424 10.6151
R584 B.n425 B.n6 10.6151
R585 B.n429 B.n6 10.6151
R586 B.n430 B.n429 10.6151
R587 B.n431 B.n430 10.6151
R588 B.n431 B.n4 10.6151
R589 B.n435 B.n4 10.6151
R590 B.n436 B.n435 10.6151
R591 B.n437 B.n436 10.6151
R592 B.n437 B.n0 10.6151
R593 B.n377 B.n22 10.6151
R594 B.n377 B.n376 10.6151
R595 B.n376 B.n375 10.6151
R596 B.n375 B.n24 10.6151
R597 B.n371 B.n24 10.6151
R598 B.n371 B.n370 10.6151
R599 B.n370 B.n369 10.6151
R600 B.n366 B.n365 10.6151
R601 B.n365 B.n364 10.6151
R602 B.n364 B.n30 10.6151
R603 B.n360 B.n30 10.6151
R604 B.n360 B.n359 10.6151
R605 B.n359 B.n358 10.6151
R606 B.n358 B.n32 10.6151
R607 B.n354 B.n32 10.6151
R608 B.n354 B.n353 10.6151
R609 B.n351 B.n36 10.6151
R610 B.n347 B.n36 10.6151
R611 B.n347 B.n346 10.6151
R612 B.n346 B.n345 10.6151
R613 B.n345 B.n38 10.6151
R614 B.n341 B.n38 10.6151
R615 B.n341 B.n340 10.6151
R616 B.n339 B.n40 10.6151
R617 B.n335 B.n40 10.6151
R618 B.n335 B.n334 10.6151
R619 B.n334 B.n333 10.6151
R620 B.n333 B.n42 10.6151
R621 B.n329 B.n42 10.6151
R622 B.n329 B.n328 10.6151
R623 B.n328 B.n327 10.6151
R624 B.n327 B.n44 10.6151
R625 B.n323 B.n44 10.6151
R626 B.n323 B.n322 10.6151
R627 B.n322 B.n321 10.6151
R628 B.n321 B.n46 10.6151
R629 B.n317 B.n46 10.6151
R630 B.n317 B.n316 10.6151
R631 B.n316 B.n315 10.6151
R632 B.n315 B.n48 10.6151
R633 B.n311 B.n48 10.6151
R634 B.n311 B.n310 10.6151
R635 B.n310 B.n309 10.6151
R636 B.n309 B.n50 10.6151
R637 B.n305 B.n50 10.6151
R638 B.n305 B.n304 10.6151
R639 B.n304 B.n303 10.6151
R640 B.n303 B.n52 10.6151
R641 B.n299 B.n52 10.6151
R642 B.n299 B.n298 10.6151
R643 B.n298 B.n297 10.6151
R644 B.n297 B.n54 10.6151
R645 B.n293 B.n54 10.6151
R646 B.n293 B.n292 10.6151
R647 B.n292 B.n291 10.6151
R648 B.n291 B.n56 10.6151
R649 B.n287 B.n56 10.6151
R650 B.n287 B.n286 10.6151
R651 B.n286 B.n285 10.6151
R652 B.n285 B.n58 10.6151
R653 B.n281 B.n58 10.6151
R654 B.n281 B.n280 10.6151
R655 B.n280 B.n279 10.6151
R656 B.n279 B.n60 10.6151
R657 B.n275 B.n60 10.6151
R658 B.n275 B.n274 10.6151
R659 B.n274 B.n273 10.6151
R660 B.n273 B.n62 10.6151
R661 B.n269 B.n62 10.6151
R662 B.n269 B.n268 10.6151
R663 B.n268 B.n267 10.6151
R664 B.n267 B.n64 10.6151
R665 B.n263 B.n64 10.6151
R666 B.n263 B.n262 10.6151
R667 B.n262 B.n261 10.6151
R668 B.n261 B.n66 10.6151
R669 B.n257 B.n66 10.6151
R670 B.n257 B.n256 10.6151
R671 B.n256 B.n255 10.6151
R672 B.n255 B.n68 10.6151
R673 B.n251 B.n68 10.6151
R674 B.n251 B.n250 10.6151
R675 B.n250 B.n249 10.6151
R676 B.n249 B.n70 10.6151
R677 B.n245 B.n70 10.6151
R678 B.n245 B.n244 10.6151
R679 B.n244 B.n243 10.6151
R680 B.n243 B.n72 10.6151
R681 B.n239 B.n72 10.6151
R682 B.n239 B.n238 10.6151
R683 B.n238 B.n237 10.6151
R684 B.n237 B.n74 10.6151
R685 B.n233 B.n74 10.6151
R686 B.n233 B.n232 10.6151
R687 B.n232 B.n231 10.6151
R688 B.n231 B.n76 10.6151
R689 B.n227 B.n76 10.6151
R690 B.n227 B.n226 10.6151
R691 B.n226 B.n225 10.6151
R692 B.n225 B.n78 10.6151
R693 B.n221 B.n78 10.6151
R694 B.n221 B.n220 10.6151
R695 B.n220 B.n219 10.6151
R696 B.n219 B.n80 10.6151
R697 B.n115 B.n1 10.6151
R698 B.n115 B.n114 10.6151
R699 B.n119 B.n114 10.6151
R700 B.n120 B.n119 10.6151
R701 B.n121 B.n120 10.6151
R702 B.n121 B.n112 10.6151
R703 B.n125 B.n112 10.6151
R704 B.n126 B.n125 10.6151
R705 B.n127 B.n126 10.6151
R706 B.n127 B.n110 10.6151
R707 B.n131 B.n110 10.6151
R708 B.n132 B.n131 10.6151
R709 B.n133 B.n132 10.6151
R710 B.n133 B.n108 10.6151
R711 B.n137 B.n108 10.6151
R712 B.n138 B.n137 10.6151
R713 B.n139 B.n138 10.6151
R714 B.n139 B.n106 10.6151
R715 B.n143 B.n106 10.6151
R716 B.n144 B.n143 10.6151
R717 B.n145 B.n144 10.6151
R718 B.n145 B.n104 10.6151
R719 B.n149 B.n104 10.6151
R720 B.n150 B.n149 10.6151
R721 B.n151 B.n150 10.6151
R722 B.n151 B.n102 10.6151
R723 B.n155 B.n102 10.6151
R724 B.n156 B.n155 10.6151
R725 B.n157 B.n156 10.6151
R726 B.n157 B.n100 10.6151
R727 B.n161 B.n100 10.6151
R728 B.n162 B.n161 10.6151
R729 B.n163 B.n162 10.6151
R730 B.n163 B.n98 10.6151
R731 B.n167 B.n98 10.6151
R732 B.n168 B.n167 10.6151
R733 B.n169 B.n168 10.6151
R734 B.n169 B.n96 10.6151
R735 B.n173 B.n96 10.6151
R736 B.n175 B.n174 10.6151
R737 B.n175 B.n94 10.6151
R738 B.n179 B.n94 10.6151
R739 B.n180 B.n179 10.6151
R740 B.n181 B.n180 10.6151
R741 B.n181 B.n92 10.6151
R742 B.n185 B.n92 10.6151
R743 B.n188 B.n187 10.6151
R744 B.n188 B.n88 10.6151
R745 B.n192 B.n88 10.6151
R746 B.n193 B.n192 10.6151
R747 B.n194 B.n193 10.6151
R748 B.n194 B.n86 10.6151
R749 B.n198 B.n86 10.6151
R750 B.n199 B.n198 10.6151
R751 B.n203 B.n199 10.6151
R752 B.n207 B.n84 10.6151
R753 B.n208 B.n207 10.6151
R754 B.n209 B.n208 10.6151
R755 B.n209 B.n82 10.6151
R756 B.n213 B.n82 10.6151
R757 B.n214 B.n213 10.6151
R758 B.n215 B.n214 10.6151
R759 B.n369 B.n28 9.36635
R760 B.n352 B.n351 9.36635
R761 B.n186 B.n185 9.36635
R762 B.n202 B.n84 9.36635
R763 B.n441 B.n0 8.11757
R764 B.n441 B.n1 8.11757
R765 B.n366 B.n28 1.24928
R766 B.n353 B.n352 1.24928
R767 B.n187 B.n186 1.24928
R768 B.n203 B.n202 1.24928
R769 VN.n25 VN.n14 161.3
R770 VN.n24 VN.n23 161.3
R771 VN.n22 VN.n15 161.3
R772 VN.n21 VN.n20 161.3
R773 VN.n19 VN.n16 161.3
R774 VN.n11 VN.n0 161.3
R775 VN.n10 VN.n9 161.3
R776 VN.n8 VN.n1 161.3
R777 VN.n7 VN.n6 161.3
R778 VN.n5 VN.n2 161.3
R779 VN.n13 VN.n12 98.4345
R780 VN.n27 VN.n26 98.4345
R781 VN.n6 VN.n1 52.5823
R782 VN.n20 VN.n15 52.5823
R783 VN.n4 VN.n3 47.9004
R784 VN.n18 VN.n17 47.9004
R785 VN.n3 VN.t5 40.4735
R786 VN.n17 VN.t3 40.4735
R787 VN VN.n27 39.6383
R788 VN.n10 VN.n1 28.2389
R789 VN.n24 VN.n15 28.2389
R790 VN.n5 VN.n4 24.3439
R791 VN.n6 VN.n5 24.3439
R792 VN.n11 VN.n10 24.3439
R793 VN.n20 VN.n19 24.3439
R794 VN.n19 VN.n18 24.3439
R795 VN.n25 VN.n24 24.3439
R796 VN.n12 VN.n11 12.1722
R797 VN.n26 VN.n25 12.1722
R798 VN.n17 VN.n16 6.7099
R799 VN.n3 VN.n2 6.7099
R800 VN.n4 VN.t1 6.17488
R801 VN.n12 VN.t2 6.17488
R802 VN.n18 VN.t4 6.17488
R803 VN.n26 VN.t0 6.17488
R804 VN.n27 VN.n14 0.278398
R805 VN.n13 VN.n0 0.278398
R806 VN.n23 VN.n14 0.189894
R807 VN.n23 VN.n22 0.189894
R808 VN.n22 VN.n21 0.189894
R809 VN.n21 VN.n16 0.189894
R810 VN.n7 VN.n2 0.189894
R811 VN.n8 VN.n7 0.189894
R812 VN.n9 VN.n8 0.189894
R813 VN.n9 VN.n0 0.189894
R814 VN VN.n13 0.153422
R815 VDD2.n1 VDD2.t0 688.403
R816 VDD2.n2 VDD2.t5 686.679
R817 VDD2.n1 VDD2.n0 634.789
R818 VDD2 VDD2.n3 634.787
R819 VDD2.n3 VDD2.t1 52.4279
R820 VDD2.n3 VDD2.t2 52.4279
R821 VDD2.n0 VDD2.t4 52.4279
R822 VDD2.n0 VDD2.t3 52.4279
R823 VDD2.n2 VDD2.n1 31.9545
R824 VDD2 VDD2.n2 1.83671
C0 VDD2 VDD1 1.33554f
C1 B VN 0.927951f
C2 VDD2 VTAIL 3.51104f
C3 VDD2 VP 0.45219f
C4 w_n3170_n1092# VN 5.75555f
C5 w_n3170_n1092# B 6.32164f
C6 VDD1 VN 0.158599f
C7 VDD1 B 1.15061f
C8 VTAIL VN 1.72224f
C9 VP VN 4.65917f
C10 VTAIL B 0.922389f
C11 VP B 1.60896f
C12 VDD1 w_n3170_n1092# 1.44295f
C13 VTAIL w_n3170_n1092# 1.2678f
C14 VP w_n3170_n1092# 6.15576f
C15 VDD2 VN 0.71242f
C16 VDD2 B 1.22112f
C17 VDD2 w_n3170_n1092# 1.52098f
C18 VDD1 VTAIL 3.45879f
C19 VDD1 VP 1.00253f
C20 VTAIL VP 1.73636f
C21 VDD2 VSUBS 0.925222f
C22 VDD1 VSUBS 1.333602f
C23 VTAIL VSUBS 0.438717f
C24 VN VSUBS 5.61161f
C25 VP VSUBS 2.194645f
C26 B VSUBS 3.288243f
C27 w_n3170_n1092# VSUBS 44.849197f
C28 VDD2.t0 VSUBS 0.04781f
C29 VDD2.t4 VSUBS 0.010238f
C30 VDD2.t3 VSUBS 0.010238f
C31 VDD2.n0 VSUBS 0.022716f
C32 VDD2.n1 VSUBS 1.53007f
C33 VDD2.t5 VSUBS 0.047349f
C34 VDD2.n2 VSUBS 1.36883f
C35 VDD2.t1 VSUBS 0.010238f
C36 VDD2.t2 VSUBS 0.010238f
C37 VDD2.n3 VSUBS 0.022714f
C38 VN.n0 VSUBS 0.076828f
C39 VN.t2 VSUBS 0.113288f
C40 VN.n1 VSUBS 0.06011f
C41 VN.n2 VSUBS 0.552827f
C42 VN.t1 VSUBS 0.113288f
C43 VN.t5 VSUBS 0.524501f
C44 VN.n3 VSUBS 0.280479f
C45 VN.n4 VSUBS 0.329363f
C46 VN.n5 VSUBS 0.109146f
C47 VN.n6 VSUBS 0.104516f
C48 VN.n7 VSUBS 0.058271f
C49 VN.n8 VSUBS 0.058271f
C50 VN.n9 VSUBS 0.058271f
C51 VN.n10 VSUBS 0.11539f
C52 VN.n11 VSUBS 0.082201f
C53 VN.n12 VSUBS 0.325174f
C54 VN.n13 VSUBS 0.088338f
C55 VN.n14 VSUBS 0.076828f
C56 VN.t0 VSUBS 0.113288f
C57 VN.n15 VSUBS 0.06011f
C58 VN.n16 VSUBS 0.552827f
C59 VN.t4 VSUBS 0.113288f
C60 VN.t3 VSUBS 0.524501f
C61 VN.n17 VSUBS 0.280479f
C62 VN.n18 VSUBS 0.329363f
C63 VN.n19 VSUBS 0.109146f
C64 VN.n20 VSUBS 0.104516f
C65 VN.n21 VSUBS 0.058271f
C66 VN.n22 VSUBS 0.058271f
C67 VN.n23 VSUBS 0.058271f
C68 VN.n24 VSUBS 0.11539f
C69 VN.n25 VSUBS 0.082201f
C70 VN.n26 VSUBS 0.325174f
C71 VN.n27 VSUBS 2.25325f
C72 B.n0 VSUBS 0.009702f
C73 B.n1 VSUBS 0.009702f
C74 B.n2 VSUBS 0.014349f
C75 B.n3 VSUBS 0.010996f
C76 B.n4 VSUBS 0.010996f
C77 B.n5 VSUBS 0.010996f
C78 B.n6 VSUBS 0.010996f
C79 B.n7 VSUBS 0.010996f
C80 B.n8 VSUBS 0.010996f
C81 B.n9 VSUBS 0.010996f
C82 B.n10 VSUBS 0.010996f
C83 B.n11 VSUBS 0.010996f
C84 B.n12 VSUBS 0.010996f
C85 B.n13 VSUBS 0.010996f
C86 B.n14 VSUBS 0.010996f
C87 B.n15 VSUBS 0.010996f
C88 B.n16 VSUBS 0.010996f
C89 B.n17 VSUBS 0.010996f
C90 B.n18 VSUBS 0.010996f
C91 B.n19 VSUBS 0.010996f
C92 B.n20 VSUBS 0.010996f
C93 B.n21 VSUBS 0.010996f
C94 B.n22 VSUBS 0.025741f
C95 B.n23 VSUBS 0.010996f
C96 B.n24 VSUBS 0.010996f
C97 B.n25 VSUBS 0.010996f
C98 B.t1 VSUBS 0.018383f
C99 B.t2 VSUBS 0.021792f
C100 B.t0 VSUBS 0.120801f
C101 B.n26 VSUBS 0.084055f
C102 B.n27 VSUBS 0.061212f
C103 B.n28 VSUBS 0.025477f
C104 B.n29 VSUBS 0.010996f
C105 B.n30 VSUBS 0.010996f
C106 B.n31 VSUBS 0.010996f
C107 B.n32 VSUBS 0.010996f
C108 B.n33 VSUBS 0.010996f
C109 B.t4 VSUBS 0.018383f
C110 B.t5 VSUBS 0.021792f
C111 B.t3 VSUBS 0.120801f
C112 B.n34 VSUBS 0.084055f
C113 B.n35 VSUBS 0.061212f
C114 B.n36 VSUBS 0.010996f
C115 B.n37 VSUBS 0.010996f
C116 B.n38 VSUBS 0.010996f
C117 B.n39 VSUBS 0.025741f
C118 B.n40 VSUBS 0.010996f
C119 B.n41 VSUBS 0.010996f
C120 B.n42 VSUBS 0.010996f
C121 B.n43 VSUBS 0.010996f
C122 B.n44 VSUBS 0.010996f
C123 B.n45 VSUBS 0.010996f
C124 B.n46 VSUBS 0.010996f
C125 B.n47 VSUBS 0.010996f
C126 B.n48 VSUBS 0.010996f
C127 B.n49 VSUBS 0.010996f
C128 B.n50 VSUBS 0.010996f
C129 B.n51 VSUBS 0.010996f
C130 B.n52 VSUBS 0.010996f
C131 B.n53 VSUBS 0.010996f
C132 B.n54 VSUBS 0.010996f
C133 B.n55 VSUBS 0.010996f
C134 B.n56 VSUBS 0.010996f
C135 B.n57 VSUBS 0.010996f
C136 B.n58 VSUBS 0.010996f
C137 B.n59 VSUBS 0.010996f
C138 B.n60 VSUBS 0.010996f
C139 B.n61 VSUBS 0.010996f
C140 B.n62 VSUBS 0.010996f
C141 B.n63 VSUBS 0.010996f
C142 B.n64 VSUBS 0.010996f
C143 B.n65 VSUBS 0.010996f
C144 B.n66 VSUBS 0.010996f
C145 B.n67 VSUBS 0.010996f
C146 B.n68 VSUBS 0.010996f
C147 B.n69 VSUBS 0.010996f
C148 B.n70 VSUBS 0.010996f
C149 B.n71 VSUBS 0.010996f
C150 B.n72 VSUBS 0.010996f
C151 B.n73 VSUBS 0.010996f
C152 B.n74 VSUBS 0.010996f
C153 B.n75 VSUBS 0.010996f
C154 B.n76 VSUBS 0.010996f
C155 B.n77 VSUBS 0.010996f
C156 B.n78 VSUBS 0.010996f
C157 B.n79 VSUBS 0.010996f
C158 B.n80 VSUBS 0.025741f
C159 B.n81 VSUBS 0.010996f
C160 B.n82 VSUBS 0.010996f
C161 B.n83 VSUBS 0.010996f
C162 B.n84 VSUBS 0.010349f
C163 B.n85 VSUBS 0.010996f
C164 B.n86 VSUBS 0.010996f
C165 B.n87 VSUBS 0.010996f
C166 B.n88 VSUBS 0.010996f
C167 B.n89 VSUBS 0.010996f
C168 B.t11 VSUBS 0.018383f
C169 B.t10 VSUBS 0.021792f
C170 B.t9 VSUBS 0.120801f
C171 B.n90 VSUBS 0.084055f
C172 B.n91 VSUBS 0.061212f
C173 B.n92 VSUBS 0.010996f
C174 B.n93 VSUBS 0.010996f
C175 B.n94 VSUBS 0.010996f
C176 B.n95 VSUBS 0.025741f
C177 B.n96 VSUBS 0.010996f
C178 B.n97 VSUBS 0.010996f
C179 B.n98 VSUBS 0.010996f
C180 B.n99 VSUBS 0.010996f
C181 B.n100 VSUBS 0.010996f
C182 B.n101 VSUBS 0.010996f
C183 B.n102 VSUBS 0.010996f
C184 B.n103 VSUBS 0.010996f
C185 B.n104 VSUBS 0.010996f
C186 B.n105 VSUBS 0.010996f
C187 B.n106 VSUBS 0.010996f
C188 B.n107 VSUBS 0.010996f
C189 B.n108 VSUBS 0.010996f
C190 B.n109 VSUBS 0.010996f
C191 B.n110 VSUBS 0.010996f
C192 B.n111 VSUBS 0.010996f
C193 B.n112 VSUBS 0.010996f
C194 B.n113 VSUBS 0.010996f
C195 B.n114 VSUBS 0.010996f
C196 B.n115 VSUBS 0.010996f
C197 B.n116 VSUBS 0.010996f
C198 B.n117 VSUBS 0.010996f
C199 B.n118 VSUBS 0.010996f
C200 B.n119 VSUBS 0.010996f
C201 B.n120 VSUBS 0.010996f
C202 B.n121 VSUBS 0.010996f
C203 B.n122 VSUBS 0.010996f
C204 B.n123 VSUBS 0.010996f
C205 B.n124 VSUBS 0.010996f
C206 B.n125 VSUBS 0.010996f
C207 B.n126 VSUBS 0.010996f
C208 B.n127 VSUBS 0.010996f
C209 B.n128 VSUBS 0.010996f
C210 B.n129 VSUBS 0.010996f
C211 B.n130 VSUBS 0.010996f
C212 B.n131 VSUBS 0.010996f
C213 B.n132 VSUBS 0.010996f
C214 B.n133 VSUBS 0.010996f
C215 B.n134 VSUBS 0.010996f
C216 B.n135 VSUBS 0.010996f
C217 B.n136 VSUBS 0.010996f
C218 B.n137 VSUBS 0.010996f
C219 B.n138 VSUBS 0.010996f
C220 B.n139 VSUBS 0.010996f
C221 B.n140 VSUBS 0.010996f
C222 B.n141 VSUBS 0.010996f
C223 B.n142 VSUBS 0.010996f
C224 B.n143 VSUBS 0.010996f
C225 B.n144 VSUBS 0.010996f
C226 B.n145 VSUBS 0.010996f
C227 B.n146 VSUBS 0.010996f
C228 B.n147 VSUBS 0.010996f
C229 B.n148 VSUBS 0.010996f
C230 B.n149 VSUBS 0.010996f
C231 B.n150 VSUBS 0.010996f
C232 B.n151 VSUBS 0.010996f
C233 B.n152 VSUBS 0.010996f
C234 B.n153 VSUBS 0.010996f
C235 B.n154 VSUBS 0.010996f
C236 B.n155 VSUBS 0.010996f
C237 B.n156 VSUBS 0.010996f
C238 B.n157 VSUBS 0.010996f
C239 B.n158 VSUBS 0.010996f
C240 B.n159 VSUBS 0.010996f
C241 B.n160 VSUBS 0.010996f
C242 B.n161 VSUBS 0.010996f
C243 B.n162 VSUBS 0.010996f
C244 B.n163 VSUBS 0.010996f
C245 B.n164 VSUBS 0.010996f
C246 B.n165 VSUBS 0.010996f
C247 B.n166 VSUBS 0.010996f
C248 B.n167 VSUBS 0.010996f
C249 B.n168 VSUBS 0.010996f
C250 B.n169 VSUBS 0.010996f
C251 B.n170 VSUBS 0.010996f
C252 B.n171 VSUBS 0.010996f
C253 B.n172 VSUBS 0.024388f
C254 B.n173 VSUBS 0.024388f
C255 B.n174 VSUBS 0.025741f
C256 B.n175 VSUBS 0.010996f
C257 B.n176 VSUBS 0.010996f
C258 B.n177 VSUBS 0.010996f
C259 B.n178 VSUBS 0.010996f
C260 B.n179 VSUBS 0.010996f
C261 B.n180 VSUBS 0.010996f
C262 B.n181 VSUBS 0.010996f
C263 B.n182 VSUBS 0.010996f
C264 B.n183 VSUBS 0.010996f
C265 B.n184 VSUBS 0.010996f
C266 B.n185 VSUBS 0.010349f
C267 B.n186 VSUBS 0.025477f
C268 B.n187 VSUBS 0.006145f
C269 B.n188 VSUBS 0.010996f
C270 B.n189 VSUBS 0.010996f
C271 B.n190 VSUBS 0.010996f
C272 B.n191 VSUBS 0.010996f
C273 B.n192 VSUBS 0.010996f
C274 B.n193 VSUBS 0.010996f
C275 B.n194 VSUBS 0.010996f
C276 B.n195 VSUBS 0.010996f
C277 B.n196 VSUBS 0.010996f
C278 B.n197 VSUBS 0.010996f
C279 B.n198 VSUBS 0.010996f
C280 B.n199 VSUBS 0.010996f
C281 B.t8 VSUBS 0.018383f
C282 B.t7 VSUBS 0.021792f
C283 B.t6 VSUBS 0.120801f
C284 B.n200 VSUBS 0.084055f
C285 B.n201 VSUBS 0.061212f
C286 B.n202 VSUBS 0.025477f
C287 B.n203 VSUBS 0.006145f
C288 B.n204 VSUBS 0.010996f
C289 B.n205 VSUBS 0.010996f
C290 B.n206 VSUBS 0.010996f
C291 B.n207 VSUBS 0.010996f
C292 B.n208 VSUBS 0.010996f
C293 B.n209 VSUBS 0.010996f
C294 B.n210 VSUBS 0.010996f
C295 B.n211 VSUBS 0.010996f
C296 B.n212 VSUBS 0.010996f
C297 B.n213 VSUBS 0.010996f
C298 B.n214 VSUBS 0.010996f
C299 B.n215 VSUBS 0.024388f
C300 B.n216 VSUBS 0.025741f
C301 B.n217 VSUBS 0.024388f
C302 B.n218 VSUBS 0.010996f
C303 B.n219 VSUBS 0.010996f
C304 B.n220 VSUBS 0.010996f
C305 B.n221 VSUBS 0.010996f
C306 B.n222 VSUBS 0.010996f
C307 B.n223 VSUBS 0.010996f
C308 B.n224 VSUBS 0.010996f
C309 B.n225 VSUBS 0.010996f
C310 B.n226 VSUBS 0.010996f
C311 B.n227 VSUBS 0.010996f
C312 B.n228 VSUBS 0.010996f
C313 B.n229 VSUBS 0.010996f
C314 B.n230 VSUBS 0.010996f
C315 B.n231 VSUBS 0.010996f
C316 B.n232 VSUBS 0.010996f
C317 B.n233 VSUBS 0.010996f
C318 B.n234 VSUBS 0.010996f
C319 B.n235 VSUBS 0.010996f
C320 B.n236 VSUBS 0.010996f
C321 B.n237 VSUBS 0.010996f
C322 B.n238 VSUBS 0.010996f
C323 B.n239 VSUBS 0.010996f
C324 B.n240 VSUBS 0.010996f
C325 B.n241 VSUBS 0.010996f
C326 B.n242 VSUBS 0.010996f
C327 B.n243 VSUBS 0.010996f
C328 B.n244 VSUBS 0.010996f
C329 B.n245 VSUBS 0.010996f
C330 B.n246 VSUBS 0.010996f
C331 B.n247 VSUBS 0.010996f
C332 B.n248 VSUBS 0.010996f
C333 B.n249 VSUBS 0.010996f
C334 B.n250 VSUBS 0.010996f
C335 B.n251 VSUBS 0.010996f
C336 B.n252 VSUBS 0.010996f
C337 B.n253 VSUBS 0.010996f
C338 B.n254 VSUBS 0.010996f
C339 B.n255 VSUBS 0.010996f
C340 B.n256 VSUBS 0.010996f
C341 B.n257 VSUBS 0.010996f
C342 B.n258 VSUBS 0.010996f
C343 B.n259 VSUBS 0.010996f
C344 B.n260 VSUBS 0.010996f
C345 B.n261 VSUBS 0.010996f
C346 B.n262 VSUBS 0.010996f
C347 B.n263 VSUBS 0.010996f
C348 B.n264 VSUBS 0.010996f
C349 B.n265 VSUBS 0.010996f
C350 B.n266 VSUBS 0.010996f
C351 B.n267 VSUBS 0.010996f
C352 B.n268 VSUBS 0.010996f
C353 B.n269 VSUBS 0.010996f
C354 B.n270 VSUBS 0.010996f
C355 B.n271 VSUBS 0.010996f
C356 B.n272 VSUBS 0.010996f
C357 B.n273 VSUBS 0.010996f
C358 B.n274 VSUBS 0.010996f
C359 B.n275 VSUBS 0.010996f
C360 B.n276 VSUBS 0.010996f
C361 B.n277 VSUBS 0.010996f
C362 B.n278 VSUBS 0.010996f
C363 B.n279 VSUBS 0.010996f
C364 B.n280 VSUBS 0.010996f
C365 B.n281 VSUBS 0.010996f
C366 B.n282 VSUBS 0.010996f
C367 B.n283 VSUBS 0.010996f
C368 B.n284 VSUBS 0.010996f
C369 B.n285 VSUBS 0.010996f
C370 B.n286 VSUBS 0.010996f
C371 B.n287 VSUBS 0.010996f
C372 B.n288 VSUBS 0.010996f
C373 B.n289 VSUBS 0.010996f
C374 B.n290 VSUBS 0.010996f
C375 B.n291 VSUBS 0.010996f
C376 B.n292 VSUBS 0.010996f
C377 B.n293 VSUBS 0.010996f
C378 B.n294 VSUBS 0.010996f
C379 B.n295 VSUBS 0.010996f
C380 B.n296 VSUBS 0.010996f
C381 B.n297 VSUBS 0.010996f
C382 B.n298 VSUBS 0.010996f
C383 B.n299 VSUBS 0.010996f
C384 B.n300 VSUBS 0.010996f
C385 B.n301 VSUBS 0.010996f
C386 B.n302 VSUBS 0.010996f
C387 B.n303 VSUBS 0.010996f
C388 B.n304 VSUBS 0.010996f
C389 B.n305 VSUBS 0.010996f
C390 B.n306 VSUBS 0.010996f
C391 B.n307 VSUBS 0.010996f
C392 B.n308 VSUBS 0.010996f
C393 B.n309 VSUBS 0.010996f
C394 B.n310 VSUBS 0.010996f
C395 B.n311 VSUBS 0.010996f
C396 B.n312 VSUBS 0.010996f
C397 B.n313 VSUBS 0.010996f
C398 B.n314 VSUBS 0.010996f
C399 B.n315 VSUBS 0.010996f
C400 B.n316 VSUBS 0.010996f
C401 B.n317 VSUBS 0.010996f
C402 B.n318 VSUBS 0.010996f
C403 B.n319 VSUBS 0.010996f
C404 B.n320 VSUBS 0.010996f
C405 B.n321 VSUBS 0.010996f
C406 B.n322 VSUBS 0.010996f
C407 B.n323 VSUBS 0.010996f
C408 B.n324 VSUBS 0.010996f
C409 B.n325 VSUBS 0.010996f
C410 B.n326 VSUBS 0.010996f
C411 B.n327 VSUBS 0.010996f
C412 B.n328 VSUBS 0.010996f
C413 B.n329 VSUBS 0.010996f
C414 B.n330 VSUBS 0.010996f
C415 B.n331 VSUBS 0.010996f
C416 B.n332 VSUBS 0.010996f
C417 B.n333 VSUBS 0.010996f
C418 B.n334 VSUBS 0.010996f
C419 B.n335 VSUBS 0.010996f
C420 B.n336 VSUBS 0.010996f
C421 B.n337 VSUBS 0.010996f
C422 B.n338 VSUBS 0.024388f
C423 B.n339 VSUBS 0.024388f
C424 B.n340 VSUBS 0.025741f
C425 B.n341 VSUBS 0.010996f
C426 B.n342 VSUBS 0.010996f
C427 B.n343 VSUBS 0.010996f
C428 B.n344 VSUBS 0.010996f
C429 B.n345 VSUBS 0.010996f
C430 B.n346 VSUBS 0.010996f
C431 B.n347 VSUBS 0.010996f
C432 B.n348 VSUBS 0.010996f
C433 B.n349 VSUBS 0.010996f
C434 B.n350 VSUBS 0.010996f
C435 B.n351 VSUBS 0.010349f
C436 B.n352 VSUBS 0.025477f
C437 B.n353 VSUBS 0.006145f
C438 B.n354 VSUBS 0.010996f
C439 B.n355 VSUBS 0.010996f
C440 B.n356 VSUBS 0.010996f
C441 B.n357 VSUBS 0.010996f
C442 B.n358 VSUBS 0.010996f
C443 B.n359 VSUBS 0.010996f
C444 B.n360 VSUBS 0.010996f
C445 B.n361 VSUBS 0.010996f
C446 B.n362 VSUBS 0.010996f
C447 B.n363 VSUBS 0.010996f
C448 B.n364 VSUBS 0.010996f
C449 B.n365 VSUBS 0.010996f
C450 B.n366 VSUBS 0.006145f
C451 B.n367 VSUBS 0.010996f
C452 B.n368 VSUBS 0.010996f
C453 B.n369 VSUBS 0.010349f
C454 B.n370 VSUBS 0.010996f
C455 B.n371 VSUBS 0.010996f
C456 B.n372 VSUBS 0.010996f
C457 B.n373 VSUBS 0.010996f
C458 B.n374 VSUBS 0.010996f
C459 B.n375 VSUBS 0.010996f
C460 B.n376 VSUBS 0.010996f
C461 B.n377 VSUBS 0.010996f
C462 B.n378 VSUBS 0.010996f
C463 B.n379 VSUBS 0.025741f
C464 B.n380 VSUBS 0.024388f
C465 B.n381 VSUBS 0.024388f
C466 B.n382 VSUBS 0.010996f
C467 B.n383 VSUBS 0.010996f
C468 B.n384 VSUBS 0.010996f
C469 B.n385 VSUBS 0.010996f
C470 B.n386 VSUBS 0.010996f
C471 B.n387 VSUBS 0.010996f
C472 B.n388 VSUBS 0.010996f
C473 B.n389 VSUBS 0.010996f
C474 B.n390 VSUBS 0.010996f
C475 B.n391 VSUBS 0.010996f
C476 B.n392 VSUBS 0.010996f
C477 B.n393 VSUBS 0.010996f
C478 B.n394 VSUBS 0.010996f
C479 B.n395 VSUBS 0.010996f
C480 B.n396 VSUBS 0.010996f
C481 B.n397 VSUBS 0.010996f
C482 B.n398 VSUBS 0.010996f
C483 B.n399 VSUBS 0.010996f
C484 B.n400 VSUBS 0.010996f
C485 B.n401 VSUBS 0.010996f
C486 B.n402 VSUBS 0.010996f
C487 B.n403 VSUBS 0.010996f
C488 B.n404 VSUBS 0.010996f
C489 B.n405 VSUBS 0.010996f
C490 B.n406 VSUBS 0.010996f
C491 B.n407 VSUBS 0.010996f
C492 B.n408 VSUBS 0.010996f
C493 B.n409 VSUBS 0.010996f
C494 B.n410 VSUBS 0.010996f
C495 B.n411 VSUBS 0.010996f
C496 B.n412 VSUBS 0.010996f
C497 B.n413 VSUBS 0.010996f
C498 B.n414 VSUBS 0.010996f
C499 B.n415 VSUBS 0.010996f
C500 B.n416 VSUBS 0.010996f
C501 B.n417 VSUBS 0.010996f
C502 B.n418 VSUBS 0.010996f
C503 B.n419 VSUBS 0.010996f
C504 B.n420 VSUBS 0.010996f
C505 B.n421 VSUBS 0.010996f
C506 B.n422 VSUBS 0.010996f
C507 B.n423 VSUBS 0.010996f
C508 B.n424 VSUBS 0.010996f
C509 B.n425 VSUBS 0.010996f
C510 B.n426 VSUBS 0.010996f
C511 B.n427 VSUBS 0.010996f
C512 B.n428 VSUBS 0.010996f
C513 B.n429 VSUBS 0.010996f
C514 B.n430 VSUBS 0.010996f
C515 B.n431 VSUBS 0.010996f
C516 B.n432 VSUBS 0.010996f
C517 B.n433 VSUBS 0.010996f
C518 B.n434 VSUBS 0.010996f
C519 B.n435 VSUBS 0.010996f
C520 B.n436 VSUBS 0.010996f
C521 B.n437 VSUBS 0.010996f
C522 B.n438 VSUBS 0.010996f
C523 B.n439 VSUBS 0.014349f
C524 B.n440 VSUBS 0.015286f
C525 B.n441 VSUBS 0.030397f
C526 VDD1.t5 VSUBS 0.046827f
C527 VDD1.t0 VSUBS 0.046778f
C528 VDD1.t1 VSUBS 0.010017f
C529 VDD1.t3 VSUBS 0.010017f
C530 VDD1.n0 VSUBS 0.022225f
C531 VDD1.n1 VSUBS 1.58463f
C532 VDD1.t4 VSUBS 0.010017f
C533 VDD1.t2 VSUBS 0.010017f
C534 VDD1.n2 VSUBS 0.022009f
C535 VDD1.n3 VSUBS 1.39466f
C536 VTAIL.t0 VSUBS 0.015733f
C537 VTAIL.t5 VSUBS 0.015733f
C538 VTAIL.n0 VSUBS 0.032403f
C539 VTAIL.n1 VSUBS 0.283363f
C540 VTAIL.t11 VSUBS 0.070649f
C541 VTAIL.n2 VSUBS 0.465978f
C542 VTAIL.t10 VSUBS 0.015733f
C543 VTAIL.t7 VSUBS 0.015733f
C544 VTAIL.n3 VSUBS 0.032403f
C545 VTAIL.n4 VSUBS 1.27215f
C546 VTAIL.t3 VSUBS 0.015733f
C547 VTAIL.t4 VSUBS 0.015733f
C548 VTAIL.n5 VSUBS 0.032403f
C549 VTAIL.n6 VSUBS 1.27215f
C550 VTAIL.t2 VSUBS 0.070649f
C551 VTAIL.n7 VSUBS 0.465978f
C552 VTAIL.t9 VSUBS 0.015733f
C553 VTAIL.t6 VSUBS 0.015733f
C554 VTAIL.n8 VSUBS 0.032403f
C555 VTAIL.n9 VSUBS 0.461316f
C556 VTAIL.t8 VSUBS 0.070649f
C557 VTAIL.n10 VSUBS 1.03152f
C558 VTAIL.t1 VSUBS 0.070649f
C559 VTAIL.n11 VSUBS 0.964172f
C560 VP.n0 VSUBS 0.080382f
C561 VP.t2 VSUBS 0.118528f
C562 VP.n1 VSUBS 0.062891f
C563 VP.n2 VSUBS 0.060966f
C564 VP.t4 VSUBS 0.118528f
C565 VP.n3 VSUBS 0.114195f
C566 VP.n4 VSUBS 0.060966f
C567 VP.n5 VSUBS 0.086004f
C568 VP.n6 VSUBS 0.080382f
C569 VP.t3 VSUBS 0.118528f
C570 VP.n7 VSUBS 0.062891f
C571 VP.n8 VSUBS 0.578399f
C572 VP.t1 VSUBS 0.118528f
C573 VP.t0 VSUBS 0.548763f
C574 VP.n9 VSUBS 0.293453f
C575 VP.n10 VSUBS 0.344599f
C576 VP.n11 VSUBS 0.114195f
C577 VP.n12 VSUBS 0.10935f
C578 VP.n13 VSUBS 0.060966f
C579 VP.n14 VSUBS 0.060966f
C580 VP.n15 VSUBS 0.060966f
C581 VP.n16 VSUBS 0.120727f
C582 VP.n17 VSUBS 0.086004f
C583 VP.n18 VSUBS 0.340215f
C584 VP.n19 VSUBS 2.32331f
C585 VP.t5 VSUBS 0.118528f
C586 VP.n20 VSUBS 0.340215f
C587 VP.n21 VSUBS 2.37883f
C588 VP.n22 VSUBS 0.080382f
C589 VP.n23 VSUBS 0.060966f
C590 VP.n24 VSUBS 0.120727f
C591 VP.n25 VSUBS 0.062891f
C592 VP.n26 VSUBS 0.10935f
C593 VP.n27 VSUBS 0.060966f
C594 VP.n28 VSUBS 0.060966f
C595 VP.n29 VSUBS 0.060966f
C596 VP.n30 VSUBS 0.199645f
C597 VP.n31 VSUBS 0.114195f
C598 VP.n32 VSUBS 0.10935f
C599 VP.n33 VSUBS 0.060966f
C600 VP.n34 VSUBS 0.060966f
C601 VP.n35 VSUBS 0.060966f
C602 VP.n36 VSUBS 0.120727f
C603 VP.n37 VSUBS 0.086004f
C604 VP.n38 VSUBS 0.340215f
C605 VP.n39 VSUBS 0.092425f
.ends

