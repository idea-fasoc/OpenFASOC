* NGSPICE file created from diff_pair_sample_0730.ext - technology: sky130A

.subckt diff_pair_sample_0730 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t0 w_n3250_n2194# sky130_fd_pr__pfet_01v8 ad=1.01145 pd=6.46 as=1.01145 ps=6.46 w=6.13 l=1.95
X1 B.t11 B.t9 B.t10 w_n3250_n2194# sky130_fd_pr__pfet_01v8 ad=2.3907 pd=13.04 as=0 ps=0 w=6.13 l=1.95
X2 VDD1.t7 VP.t0 VTAIL.t7 w_n3250_n2194# sky130_fd_pr__pfet_01v8 ad=1.01145 pd=6.46 as=2.3907 ps=13.04 w=6.13 l=1.95
X3 VTAIL.t14 VN.t1 VDD2.t1 w_n3250_n2194# sky130_fd_pr__pfet_01v8 ad=1.01145 pd=6.46 as=1.01145 ps=6.46 w=6.13 l=1.95
X4 VTAIL.t6 VP.t1 VDD1.t6 w_n3250_n2194# sky130_fd_pr__pfet_01v8 ad=2.3907 pd=13.04 as=1.01145 ps=6.46 w=6.13 l=1.95
X5 B.t8 B.t6 B.t7 w_n3250_n2194# sky130_fd_pr__pfet_01v8 ad=2.3907 pd=13.04 as=0 ps=0 w=6.13 l=1.95
X6 VDD2.t6 VN.t2 VTAIL.t13 w_n3250_n2194# sky130_fd_pr__pfet_01v8 ad=1.01145 pd=6.46 as=2.3907 ps=13.04 w=6.13 l=1.95
X7 VTAIL.t5 VP.t2 VDD1.t5 w_n3250_n2194# sky130_fd_pr__pfet_01v8 ad=1.01145 pd=6.46 as=1.01145 ps=6.46 w=6.13 l=1.95
X8 B.t5 B.t3 B.t4 w_n3250_n2194# sky130_fd_pr__pfet_01v8 ad=2.3907 pd=13.04 as=0 ps=0 w=6.13 l=1.95
X9 B.t2 B.t0 B.t1 w_n3250_n2194# sky130_fd_pr__pfet_01v8 ad=2.3907 pd=13.04 as=0 ps=0 w=6.13 l=1.95
X10 VDD2.t5 VN.t3 VTAIL.t12 w_n3250_n2194# sky130_fd_pr__pfet_01v8 ad=1.01145 pd=6.46 as=1.01145 ps=6.46 w=6.13 l=1.95
X11 VTAIL.t2 VP.t3 VDD1.t4 w_n3250_n2194# sky130_fd_pr__pfet_01v8 ad=2.3907 pd=13.04 as=1.01145 ps=6.46 w=6.13 l=1.95
X12 VTAIL.t4 VP.t4 VDD1.t3 w_n3250_n2194# sky130_fd_pr__pfet_01v8 ad=1.01145 pd=6.46 as=1.01145 ps=6.46 w=6.13 l=1.95
X13 VTAIL.t11 VN.t4 VDD2.t7 w_n3250_n2194# sky130_fd_pr__pfet_01v8 ad=2.3907 pd=13.04 as=1.01145 ps=6.46 w=6.13 l=1.95
X14 VDD1.t2 VP.t5 VTAIL.t0 w_n3250_n2194# sky130_fd_pr__pfet_01v8 ad=1.01145 pd=6.46 as=2.3907 ps=13.04 w=6.13 l=1.95
X15 VDD2.t2 VN.t5 VTAIL.t10 w_n3250_n2194# sky130_fd_pr__pfet_01v8 ad=1.01145 pd=6.46 as=1.01145 ps=6.46 w=6.13 l=1.95
X16 VDD2.t3 VN.t6 VTAIL.t9 w_n3250_n2194# sky130_fd_pr__pfet_01v8 ad=1.01145 pd=6.46 as=2.3907 ps=13.04 w=6.13 l=1.95
X17 VDD1.t1 VP.t6 VTAIL.t1 w_n3250_n2194# sky130_fd_pr__pfet_01v8 ad=1.01145 pd=6.46 as=1.01145 ps=6.46 w=6.13 l=1.95
X18 VDD1.t0 VP.t7 VTAIL.t3 w_n3250_n2194# sky130_fd_pr__pfet_01v8 ad=1.01145 pd=6.46 as=1.01145 ps=6.46 w=6.13 l=1.95
X19 VTAIL.t8 VN.t7 VDD2.t4 w_n3250_n2194# sky130_fd_pr__pfet_01v8 ad=2.3907 pd=13.04 as=1.01145 ps=6.46 w=6.13 l=1.95
R0 VN.n43 VN.n23 161.3
R1 VN.n42 VN.n41 161.3
R2 VN.n40 VN.n24 161.3
R3 VN.n39 VN.n38 161.3
R4 VN.n36 VN.n25 161.3
R5 VN.n35 VN.n34 161.3
R6 VN.n33 VN.n26 161.3
R7 VN.n32 VN.n31 161.3
R8 VN.n30 VN.n27 161.3
R9 VN.n20 VN.n0 161.3
R10 VN.n19 VN.n18 161.3
R11 VN.n17 VN.n1 161.3
R12 VN.n16 VN.n15 161.3
R13 VN.n13 VN.n2 161.3
R14 VN.n12 VN.n11 161.3
R15 VN.n10 VN.n3 161.3
R16 VN.n9 VN.n8 161.3
R17 VN.n7 VN.n4 161.3
R18 VN.n5 VN.t7 106.222
R19 VN.n28 VN.t2 106.222
R20 VN.n22 VN.n21 90.2042
R21 VN.n45 VN.n44 90.2042
R22 VN.n6 VN.t3 75.761
R23 VN.n14 VN.t1 75.761
R24 VN.n21 VN.t6 75.761
R25 VN.n29 VN.t0 75.761
R26 VN.n37 VN.t5 75.761
R27 VN.n44 VN.t4 75.761
R28 VN.n6 VN.n5 63.0337
R29 VN.n29 VN.n28 63.0337
R30 VN.n19 VN.n1 56.5193
R31 VN.n42 VN.n24 56.5193
R32 VN VN.n45 43.7103
R33 VN.n8 VN.n3 40.4934
R34 VN.n12 VN.n3 40.4934
R35 VN.n31 VN.n26 40.4934
R36 VN.n35 VN.n26 40.4934
R37 VN.n8 VN.n7 24.4675
R38 VN.n13 VN.n12 24.4675
R39 VN.n15 VN.n1 24.4675
R40 VN.n20 VN.n19 24.4675
R41 VN.n31 VN.n30 24.4675
R42 VN.n38 VN.n24 24.4675
R43 VN.n36 VN.n35 24.4675
R44 VN.n43 VN.n42 24.4675
R45 VN.n21 VN.n20 20.5528
R46 VN.n44 VN.n43 20.5528
R47 VN.n15 VN.n14 17.6167
R48 VN.n38 VN.n37 17.6167
R49 VN.n28 VN.n27 13.2264
R50 VN.n5 VN.n4 13.2264
R51 VN.n7 VN.n6 6.85126
R52 VN.n14 VN.n13 6.85126
R53 VN.n30 VN.n29 6.85126
R54 VN.n37 VN.n36 6.85126
R55 VN.n45 VN.n23 0.278367
R56 VN.n22 VN.n0 0.278367
R57 VN.n41 VN.n23 0.189894
R58 VN.n41 VN.n40 0.189894
R59 VN.n40 VN.n39 0.189894
R60 VN.n39 VN.n25 0.189894
R61 VN.n34 VN.n25 0.189894
R62 VN.n34 VN.n33 0.189894
R63 VN.n33 VN.n32 0.189894
R64 VN.n32 VN.n27 0.189894
R65 VN.n9 VN.n4 0.189894
R66 VN.n10 VN.n9 0.189894
R67 VN.n11 VN.n10 0.189894
R68 VN.n11 VN.n2 0.189894
R69 VN.n16 VN.n2 0.189894
R70 VN.n17 VN.n16 0.189894
R71 VN.n18 VN.n17 0.189894
R72 VN.n18 VN.n0 0.189894
R73 VN VN.n22 0.153454
R74 VDD2.n2 VDD2.n1 93.0733
R75 VDD2.n2 VDD2.n0 93.0733
R76 VDD2 VDD2.n5 93.0696
R77 VDD2.n4 VDD2.n3 92.146
R78 VDD2.n4 VDD2.n2 37.8446
R79 VDD2.n5 VDD2.t0 5.30311
R80 VDD2.n5 VDD2.t6 5.30311
R81 VDD2.n3 VDD2.t7 5.30311
R82 VDD2.n3 VDD2.t2 5.30311
R83 VDD2.n1 VDD2.t1 5.30311
R84 VDD2.n1 VDD2.t3 5.30311
R85 VDD2.n0 VDD2.t4 5.30311
R86 VDD2.n0 VDD2.t5 5.30311
R87 VDD2 VDD2.n4 1.04145
R88 VTAIL.n11 VTAIL.t6 80.7699
R89 VTAIL.n10 VTAIL.t13 80.7699
R90 VTAIL.n7 VTAIL.t11 80.7699
R91 VTAIL.n15 VTAIL.t9 80.7689
R92 VTAIL.n2 VTAIL.t8 80.7689
R93 VTAIL.n3 VTAIL.t0 80.7689
R94 VTAIL.n6 VTAIL.t2 80.7689
R95 VTAIL.n14 VTAIL.t7 80.7689
R96 VTAIL.n13 VTAIL.n12 75.4673
R97 VTAIL.n9 VTAIL.n8 75.4673
R98 VTAIL.n1 VTAIL.n0 75.4671
R99 VTAIL.n5 VTAIL.n4 75.4671
R100 VTAIL.n15 VTAIL.n14 19.6169
R101 VTAIL.n7 VTAIL.n6 19.6169
R102 VTAIL.n0 VTAIL.t12 5.30311
R103 VTAIL.n0 VTAIL.t14 5.30311
R104 VTAIL.n4 VTAIL.t1 5.30311
R105 VTAIL.n4 VTAIL.t5 5.30311
R106 VTAIL.n12 VTAIL.t3 5.30311
R107 VTAIL.n12 VTAIL.t4 5.30311
R108 VTAIL.n8 VTAIL.t10 5.30311
R109 VTAIL.n8 VTAIL.t15 5.30311
R110 VTAIL.n9 VTAIL.n7 1.96602
R111 VTAIL.n10 VTAIL.n9 1.96602
R112 VTAIL.n13 VTAIL.n11 1.96602
R113 VTAIL.n14 VTAIL.n13 1.96602
R114 VTAIL.n6 VTAIL.n5 1.96602
R115 VTAIL.n5 VTAIL.n3 1.96602
R116 VTAIL.n2 VTAIL.n1 1.96602
R117 VTAIL VTAIL.n15 1.90783
R118 VTAIL.n11 VTAIL.n10 0.470328
R119 VTAIL.n3 VTAIL.n2 0.470328
R120 VTAIL VTAIL.n1 0.0586897
R121 B.n300 B.n299 585
R122 B.n298 B.n99 585
R123 B.n297 B.n296 585
R124 B.n295 B.n100 585
R125 B.n294 B.n293 585
R126 B.n292 B.n101 585
R127 B.n291 B.n290 585
R128 B.n289 B.n102 585
R129 B.n288 B.n287 585
R130 B.n286 B.n103 585
R131 B.n285 B.n284 585
R132 B.n283 B.n104 585
R133 B.n282 B.n281 585
R134 B.n280 B.n105 585
R135 B.n279 B.n278 585
R136 B.n277 B.n106 585
R137 B.n276 B.n275 585
R138 B.n274 B.n107 585
R139 B.n273 B.n272 585
R140 B.n271 B.n108 585
R141 B.n270 B.n269 585
R142 B.n268 B.n109 585
R143 B.n267 B.n266 585
R144 B.n265 B.n110 585
R145 B.n263 B.n262 585
R146 B.n261 B.n113 585
R147 B.n260 B.n259 585
R148 B.n258 B.n114 585
R149 B.n257 B.n256 585
R150 B.n255 B.n115 585
R151 B.n254 B.n253 585
R152 B.n252 B.n116 585
R153 B.n251 B.n250 585
R154 B.n249 B.n117 585
R155 B.n248 B.n247 585
R156 B.n243 B.n118 585
R157 B.n242 B.n241 585
R158 B.n240 B.n119 585
R159 B.n239 B.n238 585
R160 B.n237 B.n120 585
R161 B.n236 B.n235 585
R162 B.n234 B.n121 585
R163 B.n233 B.n232 585
R164 B.n231 B.n122 585
R165 B.n230 B.n229 585
R166 B.n228 B.n123 585
R167 B.n227 B.n226 585
R168 B.n225 B.n124 585
R169 B.n224 B.n223 585
R170 B.n222 B.n125 585
R171 B.n221 B.n220 585
R172 B.n219 B.n126 585
R173 B.n218 B.n217 585
R174 B.n216 B.n127 585
R175 B.n215 B.n214 585
R176 B.n213 B.n128 585
R177 B.n212 B.n211 585
R178 B.n210 B.n129 585
R179 B.n301 B.n98 585
R180 B.n303 B.n302 585
R181 B.n304 B.n97 585
R182 B.n306 B.n305 585
R183 B.n307 B.n96 585
R184 B.n309 B.n308 585
R185 B.n310 B.n95 585
R186 B.n312 B.n311 585
R187 B.n313 B.n94 585
R188 B.n315 B.n314 585
R189 B.n316 B.n93 585
R190 B.n318 B.n317 585
R191 B.n319 B.n92 585
R192 B.n321 B.n320 585
R193 B.n322 B.n91 585
R194 B.n324 B.n323 585
R195 B.n325 B.n90 585
R196 B.n327 B.n326 585
R197 B.n328 B.n89 585
R198 B.n330 B.n329 585
R199 B.n331 B.n88 585
R200 B.n333 B.n332 585
R201 B.n334 B.n87 585
R202 B.n336 B.n335 585
R203 B.n337 B.n86 585
R204 B.n339 B.n338 585
R205 B.n340 B.n85 585
R206 B.n342 B.n341 585
R207 B.n343 B.n84 585
R208 B.n345 B.n344 585
R209 B.n346 B.n83 585
R210 B.n348 B.n347 585
R211 B.n349 B.n82 585
R212 B.n351 B.n350 585
R213 B.n352 B.n81 585
R214 B.n354 B.n353 585
R215 B.n355 B.n80 585
R216 B.n357 B.n356 585
R217 B.n358 B.n79 585
R218 B.n360 B.n359 585
R219 B.n361 B.n78 585
R220 B.n363 B.n362 585
R221 B.n364 B.n77 585
R222 B.n366 B.n365 585
R223 B.n367 B.n76 585
R224 B.n369 B.n368 585
R225 B.n370 B.n75 585
R226 B.n372 B.n371 585
R227 B.n373 B.n74 585
R228 B.n375 B.n374 585
R229 B.n376 B.n73 585
R230 B.n378 B.n377 585
R231 B.n379 B.n72 585
R232 B.n381 B.n380 585
R233 B.n382 B.n71 585
R234 B.n384 B.n383 585
R235 B.n385 B.n70 585
R236 B.n387 B.n386 585
R237 B.n388 B.n69 585
R238 B.n390 B.n389 585
R239 B.n391 B.n68 585
R240 B.n393 B.n392 585
R241 B.n394 B.n67 585
R242 B.n396 B.n395 585
R243 B.n397 B.n66 585
R244 B.n399 B.n398 585
R245 B.n400 B.n65 585
R246 B.n402 B.n401 585
R247 B.n403 B.n64 585
R248 B.n405 B.n404 585
R249 B.n406 B.n63 585
R250 B.n408 B.n407 585
R251 B.n409 B.n62 585
R252 B.n411 B.n410 585
R253 B.n412 B.n61 585
R254 B.n414 B.n413 585
R255 B.n415 B.n60 585
R256 B.n417 B.n416 585
R257 B.n418 B.n59 585
R258 B.n420 B.n419 585
R259 B.n421 B.n58 585
R260 B.n423 B.n422 585
R261 B.n424 B.n57 585
R262 B.n426 B.n425 585
R263 B.n514 B.n513 585
R264 B.n512 B.n23 585
R265 B.n511 B.n510 585
R266 B.n509 B.n24 585
R267 B.n508 B.n507 585
R268 B.n506 B.n25 585
R269 B.n505 B.n504 585
R270 B.n503 B.n26 585
R271 B.n502 B.n501 585
R272 B.n500 B.n27 585
R273 B.n499 B.n498 585
R274 B.n497 B.n28 585
R275 B.n496 B.n495 585
R276 B.n494 B.n29 585
R277 B.n493 B.n492 585
R278 B.n491 B.n30 585
R279 B.n490 B.n489 585
R280 B.n488 B.n31 585
R281 B.n487 B.n486 585
R282 B.n485 B.n32 585
R283 B.n484 B.n483 585
R284 B.n482 B.n33 585
R285 B.n481 B.n480 585
R286 B.n479 B.n34 585
R287 B.n478 B.n477 585
R288 B.n476 B.n35 585
R289 B.n475 B.n474 585
R290 B.n473 B.n39 585
R291 B.n472 B.n471 585
R292 B.n470 B.n40 585
R293 B.n469 B.n468 585
R294 B.n467 B.n41 585
R295 B.n466 B.n465 585
R296 B.n464 B.n42 585
R297 B.n462 B.n461 585
R298 B.n460 B.n45 585
R299 B.n459 B.n458 585
R300 B.n457 B.n46 585
R301 B.n456 B.n455 585
R302 B.n454 B.n47 585
R303 B.n453 B.n452 585
R304 B.n451 B.n48 585
R305 B.n450 B.n449 585
R306 B.n448 B.n49 585
R307 B.n447 B.n446 585
R308 B.n445 B.n50 585
R309 B.n444 B.n443 585
R310 B.n442 B.n51 585
R311 B.n441 B.n440 585
R312 B.n439 B.n52 585
R313 B.n438 B.n437 585
R314 B.n436 B.n53 585
R315 B.n435 B.n434 585
R316 B.n433 B.n54 585
R317 B.n432 B.n431 585
R318 B.n430 B.n55 585
R319 B.n429 B.n428 585
R320 B.n427 B.n56 585
R321 B.n515 B.n22 585
R322 B.n517 B.n516 585
R323 B.n518 B.n21 585
R324 B.n520 B.n519 585
R325 B.n521 B.n20 585
R326 B.n523 B.n522 585
R327 B.n524 B.n19 585
R328 B.n526 B.n525 585
R329 B.n527 B.n18 585
R330 B.n529 B.n528 585
R331 B.n530 B.n17 585
R332 B.n532 B.n531 585
R333 B.n533 B.n16 585
R334 B.n535 B.n534 585
R335 B.n536 B.n15 585
R336 B.n538 B.n537 585
R337 B.n539 B.n14 585
R338 B.n541 B.n540 585
R339 B.n542 B.n13 585
R340 B.n544 B.n543 585
R341 B.n545 B.n12 585
R342 B.n547 B.n546 585
R343 B.n548 B.n11 585
R344 B.n550 B.n549 585
R345 B.n551 B.n10 585
R346 B.n553 B.n552 585
R347 B.n554 B.n9 585
R348 B.n556 B.n555 585
R349 B.n557 B.n8 585
R350 B.n559 B.n558 585
R351 B.n560 B.n7 585
R352 B.n562 B.n561 585
R353 B.n563 B.n6 585
R354 B.n565 B.n564 585
R355 B.n566 B.n5 585
R356 B.n568 B.n567 585
R357 B.n569 B.n4 585
R358 B.n571 B.n570 585
R359 B.n572 B.n3 585
R360 B.n574 B.n573 585
R361 B.n575 B.n0 585
R362 B.n2 B.n1 585
R363 B.n150 B.n149 585
R364 B.n152 B.n151 585
R365 B.n153 B.n148 585
R366 B.n155 B.n154 585
R367 B.n156 B.n147 585
R368 B.n158 B.n157 585
R369 B.n159 B.n146 585
R370 B.n161 B.n160 585
R371 B.n162 B.n145 585
R372 B.n164 B.n163 585
R373 B.n165 B.n144 585
R374 B.n167 B.n166 585
R375 B.n168 B.n143 585
R376 B.n170 B.n169 585
R377 B.n171 B.n142 585
R378 B.n173 B.n172 585
R379 B.n174 B.n141 585
R380 B.n176 B.n175 585
R381 B.n177 B.n140 585
R382 B.n179 B.n178 585
R383 B.n180 B.n139 585
R384 B.n182 B.n181 585
R385 B.n183 B.n138 585
R386 B.n185 B.n184 585
R387 B.n186 B.n137 585
R388 B.n188 B.n187 585
R389 B.n189 B.n136 585
R390 B.n191 B.n190 585
R391 B.n192 B.n135 585
R392 B.n194 B.n193 585
R393 B.n195 B.n134 585
R394 B.n197 B.n196 585
R395 B.n198 B.n133 585
R396 B.n200 B.n199 585
R397 B.n201 B.n132 585
R398 B.n203 B.n202 585
R399 B.n204 B.n131 585
R400 B.n206 B.n205 585
R401 B.n207 B.n130 585
R402 B.n209 B.n208 585
R403 B.n210 B.n209 545.355
R404 B.n299 B.n98 545.355
R405 B.n425 B.n56 545.355
R406 B.n515 B.n514 545.355
R407 B.n244 B.t6 282.558
R408 B.n111 B.t3 282.558
R409 B.n43 B.t9 282.558
R410 B.n36 B.t0 282.558
R411 B.n577 B.n576 256.663
R412 B.n576 B.n575 235.042
R413 B.n576 B.n2 235.042
R414 B.n211 B.n210 163.367
R415 B.n211 B.n128 163.367
R416 B.n215 B.n128 163.367
R417 B.n216 B.n215 163.367
R418 B.n217 B.n216 163.367
R419 B.n217 B.n126 163.367
R420 B.n221 B.n126 163.367
R421 B.n222 B.n221 163.367
R422 B.n223 B.n222 163.367
R423 B.n223 B.n124 163.367
R424 B.n227 B.n124 163.367
R425 B.n228 B.n227 163.367
R426 B.n229 B.n228 163.367
R427 B.n229 B.n122 163.367
R428 B.n233 B.n122 163.367
R429 B.n234 B.n233 163.367
R430 B.n235 B.n234 163.367
R431 B.n235 B.n120 163.367
R432 B.n239 B.n120 163.367
R433 B.n240 B.n239 163.367
R434 B.n241 B.n240 163.367
R435 B.n241 B.n118 163.367
R436 B.n248 B.n118 163.367
R437 B.n249 B.n248 163.367
R438 B.n250 B.n249 163.367
R439 B.n250 B.n116 163.367
R440 B.n254 B.n116 163.367
R441 B.n255 B.n254 163.367
R442 B.n256 B.n255 163.367
R443 B.n256 B.n114 163.367
R444 B.n260 B.n114 163.367
R445 B.n261 B.n260 163.367
R446 B.n262 B.n261 163.367
R447 B.n262 B.n110 163.367
R448 B.n267 B.n110 163.367
R449 B.n268 B.n267 163.367
R450 B.n269 B.n268 163.367
R451 B.n269 B.n108 163.367
R452 B.n273 B.n108 163.367
R453 B.n274 B.n273 163.367
R454 B.n275 B.n274 163.367
R455 B.n275 B.n106 163.367
R456 B.n279 B.n106 163.367
R457 B.n280 B.n279 163.367
R458 B.n281 B.n280 163.367
R459 B.n281 B.n104 163.367
R460 B.n285 B.n104 163.367
R461 B.n286 B.n285 163.367
R462 B.n287 B.n286 163.367
R463 B.n287 B.n102 163.367
R464 B.n291 B.n102 163.367
R465 B.n292 B.n291 163.367
R466 B.n293 B.n292 163.367
R467 B.n293 B.n100 163.367
R468 B.n297 B.n100 163.367
R469 B.n298 B.n297 163.367
R470 B.n299 B.n298 163.367
R471 B.n425 B.n424 163.367
R472 B.n424 B.n423 163.367
R473 B.n423 B.n58 163.367
R474 B.n419 B.n58 163.367
R475 B.n419 B.n418 163.367
R476 B.n418 B.n417 163.367
R477 B.n417 B.n60 163.367
R478 B.n413 B.n60 163.367
R479 B.n413 B.n412 163.367
R480 B.n412 B.n411 163.367
R481 B.n411 B.n62 163.367
R482 B.n407 B.n62 163.367
R483 B.n407 B.n406 163.367
R484 B.n406 B.n405 163.367
R485 B.n405 B.n64 163.367
R486 B.n401 B.n64 163.367
R487 B.n401 B.n400 163.367
R488 B.n400 B.n399 163.367
R489 B.n399 B.n66 163.367
R490 B.n395 B.n66 163.367
R491 B.n395 B.n394 163.367
R492 B.n394 B.n393 163.367
R493 B.n393 B.n68 163.367
R494 B.n389 B.n68 163.367
R495 B.n389 B.n388 163.367
R496 B.n388 B.n387 163.367
R497 B.n387 B.n70 163.367
R498 B.n383 B.n70 163.367
R499 B.n383 B.n382 163.367
R500 B.n382 B.n381 163.367
R501 B.n381 B.n72 163.367
R502 B.n377 B.n72 163.367
R503 B.n377 B.n376 163.367
R504 B.n376 B.n375 163.367
R505 B.n375 B.n74 163.367
R506 B.n371 B.n74 163.367
R507 B.n371 B.n370 163.367
R508 B.n370 B.n369 163.367
R509 B.n369 B.n76 163.367
R510 B.n365 B.n76 163.367
R511 B.n365 B.n364 163.367
R512 B.n364 B.n363 163.367
R513 B.n363 B.n78 163.367
R514 B.n359 B.n78 163.367
R515 B.n359 B.n358 163.367
R516 B.n358 B.n357 163.367
R517 B.n357 B.n80 163.367
R518 B.n353 B.n80 163.367
R519 B.n353 B.n352 163.367
R520 B.n352 B.n351 163.367
R521 B.n351 B.n82 163.367
R522 B.n347 B.n82 163.367
R523 B.n347 B.n346 163.367
R524 B.n346 B.n345 163.367
R525 B.n345 B.n84 163.367
R526 B.n341 B.n84 163.367
R527 B.n341 B.n340 163.367
R528 B.n340 B.n339 163.367
R529 B.n339 B.n86 163.367
R530 B.n335 B.n86 163.367
R531 B.n335 B.n334 163.367
R532 B.n334 B.n333 163.367
R533 B.n333 B.n88 163.367
R534 B.n329 B.n88 163.367
R535 B.n329 B.n328 163.367
R536 B.n328 B.n327 163.367
R537 B.n327 B.n90 163.367
R538 B.n323 B.n90 163.367
R539 B.n323 B.n322 163.367
R540 B.n322 B.n321 163.367
R541 B.n321 B.n92 163.367
R542 B.n317 B.n92 163.367
R543 B.n317 B.n316 163.367
R544 B.n316 B.n315 163.367
R545 B.n315 B.n94 163.367
R546 B.n311 B.n94 163.367
R547 B.n311 B.n310 163.367
R548 B.n310 B.n309 163.367
R549 B.n309 B.n96 163.367
R550 B.n305 B.n96 163.367
R551 B.n305 B.n304 163.367
R552 B.n304 B.n303 163.367
R553 B.n303 B.n98 163.367
R554 B.n514 B.n23 163.367
R555 B.n510 B.n23 163.367
R556 B.n510 B.n509 163.367
R557 B.n509 B.n508 163.367
R558 B.n508 B.n25 163.367
R559 B.n504 B.n25 163.367
R560 B.n504 B.n503 163.367
R561 B.n503 B.n502 163.367
R562 B.n502 B.n27 163.367
R563 B.n498 B.n27 163.367
R564 B.n498 B.n497 163.367
R565 B.n497 B.n496 163.367
R566 B.n496 B.n29 163.367
R567 B.n492 B.n29 163.367
R568 B.n492 B.n491 163.367
R569 B.n491 B.n490 163.367
R570 B.n490 B.n31 163.367
R571 B.n486 B.n31 163.367
R572 B.n486 B.n485 163.367
R573 B.n485 B.n484 163.367
R574 B.n484 B.n33 163.367
R575 B.n480 B.n33 163.367
R576 B.n480 B.n479 163.367
R577 B.n479 B.n478 163.367
R578 B.n478 B.n35 163.367
R579 B.n474 B.n35 163.367
R580 B.n474 B.n473 163.367
R581 B.n473 B.n472 163.367
R582 B.n472 B.n40 163.367
R583 B.n468 B.n40 163.367
R584 B.n468 B.n467 163.367
R585 B.n467 B.n466 163.367
R586 B.n466 B.n42 163.367
R587 B.n461 B.n42 163.367
R588 B.n461 B.n460 163.367
R589 B.n460 B.n459 163.367
R590 B.n459 B.n46 163.367
R591 B.n455 B.n46 163.367
R592 B.n455 B.n454 163.367
R593 B.n454 B.n453 163.367
R594 B.n453 B.n48 163.367
R595 B.n449 B.n48 163.367
R596 B.n449 B.n448 163.367
R597 B.n448 B.n447 163.367
R598 B.n447 B.n50 163.367
R599 B.n443 B.n50 163.367
R600 B.n443 B.n442 163.367
R601 B.n442 B.n441 163.367
R602 B.n441 B.n52 163.367
R603 B.n437 B.n52 163.367
R604 B.n437 B.n436 163.367
R605 B.n436 B.n435 163.367
R606 B.n435 B.n54 163.367
R607 B.n431 B.n54 163.367
R608 B.n431 B.n430 163.367
R609 B.n430 B.n429 163.367
R610 B.n429 B.n56 163.367
R611 B.n516 B.n515 163.367
R612 B.n516 B.n21 163.367
R613 B.n520 B.n21 163.367
R614 B.n521 B.n520 163.367
R615 B.n522 B.n521 163.367
R616 B.n522 B.n19 163.367
R617 B.n526 B.n19 163.367
R618 B.n527 B.n526 163.367
R619 B.n528 B.n527 163.367
R620 B.n528 B.n17 163.367
R621 B.n532 B.n17 163.367
R622 B.n533 B.n532 163.367
R623 B.n534 B.n533 163.367
R624 B.n534 B.n15 163.367
R625 B.n538 B.n15 163.367
R626 B.n539 B.n538 163.367
R627 B.n540 B.n539 163.367
R628 B.n540 B.n13 163.367
R629 B.n544 B.n13 163.367
R630 B.n545 B.n544 163.367
R631 B.n546 B.n545 163.367
R632 B.n546 B.n11 163.367
R633 B.n550 B.n11 163.367
R634 B.n551 B.n550 163.367
R635 B.n552 B.n551 163.367
R636 B.n552 B.n9 163.367
R637 B.n556 B.n9 163.367
R638 B.n557 B.n556 163.367
R639 B.n558 B.n557 163.367
R640 B.n558 B.n7 163.367
R641 B.n562 B.n7 163.367
R642 B.n563 B.n562 163.367
R643 B.n564 B.n563 163.367
R644 B.n564 B.n5 163.367
R645 B.n568 B.n5 163.367
R646 B.n569 B.n568 163.367
R647 B.n570 B.n569 163.367
R648 B.n570 B.n3 163.367
R649 B.n574 B.n3 163.367
R650 B.n575 B.n574 163.367
R651 B.n150 B.n2 163.367
R652 B.n151 B.n150 163.367
R653 B.n151 B.n148 163.367
R654 B.n155 B.n148 163.367
R655 B.n156 B.n155 163.367
R656 B.n157 B.n156 163.367
R657 B.n157 B.n146 163.367
R658 B.n161 B.n146 163.367
R659 B.n162 B.n161 163.367
R660 B.n163 B.n162 163.367
R661 B.n163 B.n144 163.367
R662 B.n167 B.n144 163.367
R663 B.n168 B.n167 163.367
R664 B.n169 B.n168 163.367
R665 B.n169 B.n142 163.367
R666 B.n173 B.n142 163.367
R667 B.n174 B.n173 163.367
R668 B.n175 B.n174 163.367
R669 B.n175 B.n140 163.367
R670 B.n179 B.n140 163.367
R671 B.n180 B.n179 163.367
R672 B.n181 B.n180 163.367
R673 B.n181 B.n138 163.367
R674 B.n185 B.n138 163.367
R675 B.n186 B.n185 163.367
R676 B.n187 B.n186 163.367
R677 B.n187 B.n136 163.367
R678 B.n191 B.n136 163.367
R679 B.n192 B.n191 163.367
R680 B.n193 B.n192 163.367
R681 B.n193 B.n134 163.367
R682 B.n197 B.n134 163.367
R683 B.n198 B.n197 163.367
R684 B.n199 B.n198 163.367
R685 B.n199 B.n132 163.367
R686 B.n203 B.n132 163.367
R687 B.n204 B.n203 163.367
R688 B.n205 B.n204 163.367
R689 B.n205 B.n130 163.367
R690 B.n209 B.n130 163.367
R691 B.n111 B.t4 155.177
R692 B.n43 B.t11 155.177
R693 B.n244 B.t7 155.171
R694 B.n36 B.t2 155.171
R695 B.n112 B.t5 110.959
R696 B.n44 B.t10 110.959
R697 B.n245 B.t8 110.951
R698 B.n37 B.t1 110.951
R699 B.n246 B.n245 59.5399
R700 B.n264 B.n112 59.5399
R701 B.n463 B.n44 59.5399
R702 B.n38 B.n37 59.5399
R703 B.n245 B.n244 44.2187
R704 B.n112 B.n111 44.2187
R705 B.n44 B.n43 44.2187
R706 B.n37 B.n36 44.2187
R707 B.n513 B.n22 35.4346
R708 B.n427 B.n426 35.4346
R709 B.n208 B.n129 35.4346
R710 B.n301 B.n300 35.4346
R711 B B.n577 18.0485
R712 B.n517 B.n22 10.6151
R713 B.n518 B.n517 10.6151
R714 B.n519 B.n518 10.6151
R715 B.n519 B.n20 10.6151
R716 B.n523 B.n20 10.6151
R717 B.n524 B.n523 10.6151
R718 B.n525 B.n524 10.6151
R719 B.n525 B.n18 10.6151
R720 B.n529 B.n18 10.6151
R721 B.n530 B.n529 10.6151
R722 B.n531 B.n530 10.6151
R723 B.n531 B.n16 10.6151
R724 B.n535 B.n16 10.6151
R725 B.n536 B.n535 10.6151
R726 B.n537 B.n536 10.6151
R727 B.n537 B.n14 10.6151
R728 B.n541 B.n14 10.6151
R729 B.n542 B.n541 10.6151
R730 B.n543 B.n542 10.6151
R731 B.n543 B.n12 10.6151
R732 B.n547 B.n12 10.6151
R733 B.n548 B.n547 10.6151
R734 B.n549 B.n548 10.6151
R735 B.n549 B.n10 10.6151
R736 B.n553 B.n10 10.6151
R737 B.n554 B.n553 10.6151
R738 B.n555 B.n554 10.6151
R739 B.n555 B.n8 10.6151
R740 B.n559 B.n8 10.6151
R741 B.n560 B.n559 10.6151
R742 B.n561 B.n560 10.6151
R743 B.n561 B.n6 10.6151
R744 B.n565 B.n6 10.6151
R745 B.n566 B.n565 10.6151
R746 B.n567 B.n566 10.6151
R747 B.n567 B.n4 10.6151
R748 B.n571 B.n4 10.6151
R749 B.n572 B.n571 10.6151
R750 B.n573 B.n572 10.6151
R751 B.n573 B.n0 10.6151
R752 B.n513 B.n512 10.6151
R753 B.n512 B.n511 10.6151
R754 B.n511 B.n24 10.6151
R755 B.n507 B.n24 10.6151
R756 B.n507 B.n506 10.6151
R757 B.n506 B.n505 10.6151
R758 B.n505 B.n26 10.6151
R759 B.n501 B.n26 10.6151
R760 B.n501 B.n500 10.6151
R761 B.n500 B.n499 10.6151
R762 B.n499 B.n28 10.6151
R763 B.n495 B.n28 10.6151
R764 B.n495 B.n494 10.6151
R765 B.n494 B.n493 10.6151
R766 B.n493 B.n30 10.6151
R767 B.n489 B.n30 10.6151
R768 B.n489 B.n488 10.6151
R769 B.n488 B.n487 10.6151
R770 B.n487 B.n32 10.6151
R771 B.n483 B.n32 10.6151
R772 B.n483 B.n482 10.6151
R773 B.n482 B.n481 10.6151
R774 B.n481 B.n34 10.6151
R775 B.n477 B.n476 10.6151
R776 B.n476 B.n475 10.6151
R777 B.n475 B.n39 10.6151
R778 B.n471 B.n39 10.6151
R779 B.n471 B.n470 10.6151
R780 B.n470 B.n469 10.6151
R781 B.n469 B.n41 10.6151
R782 B.n465 B.n41 10.6151
R783 B.n465 B.n464 10.6151
R784 B.n462 B.n45 10.6151
R785 B.n458 B.n45 10.6151
R786 B.n458 B.n457 10.6151
R787 B.n457 B.n456 10.6151
R788 B.n456 B.n47 10.6151
R789 B.n452 B.n47 10.6151
R790 B.n452 B.n451 10.6151
R791 B.n451 B.n450 10.6151
R792 B.n450 B.n49 10.6151
R793 B.n446 B.n49 10.6151
R794 B.n446 B.n445 10.6151
R795 B.n445 B.n444 10.6151
R796 B.n444 B.n51 10.6151
R797 B.n440 B.n51 10.6151
R798 B.n440 B.n439 10.6151
R799 B.n439 B.n438 10.6151
R800 B.n438 B.n53 10.6151
R801 B.n434 B.n53 10.6151
R802 B.n434 B.n433 10.6151
R803 B.n433 B.n432 10.6151
R804 B.n432 B.n55 10.6151
R805 B.n428 B.n55 10.6151
R806 B.n428 B.n427 10.6151
R807 B.n426 B.n57 10.6151
R808 B.n422 B.n57 10.6151
R809 B.n422 B.n421 10.6151
R810 B.n421 B.n420 10.6151
R811 B.n420 B.n59 10.6151
R812 B.n416 B.n59 10.6151
R813 B.n416 B.n415 10.6151
R814 B.n415 B.n414 10.6151
R815 B.n414 B.n61 10.6151
R816 B.n410 B.n61 10.6151
R817 B.n410 B.n409 10.6151
R818 B.n409 B.n408 10.6151
R819 B.n408 B.n63 10.6151
R820 B.n404 B.n63 10.6151
R821 B.n404 B.n403 10.6151
R822 B.n403 B.n402 10.6151
R823 B.n402 B.n65 10.6151
R824 B.n398 B.n65 10.6151
R825 B.n398 B.n397 10.6151
R826 B.n397 B.n396 10.6151
R827 B.n396 B.n67 10.6151
R828 B.n392 B.n67 10.6151
R829 B.n392 B.n391 10.6151
R830 B.n391 B.n390 10.6151
R831 B.n390 B.n69 10.6151
R832 B.n386 B.n69 10.6151
R833 B.n386 B.n385 10.6151
R834 B.n385 B.n384 10.6151
R835 B.n384 B.n71 10.6151
R836 B.n380 B.n71 10.6151
R837 B.n380 B.n379 10.6151
R838 B.n379 B.n378 10.6151
R839 B.n378 B.n73 10.6151
R840 B.n374 B.n73 10.6151
R841 B.n374 B.n373 10.6151
R842 B.n373 B.n372 10.6151
R843 B.n372 B.n75 10.6151
R844 B.n368 B.n75 10.6151
R845 B.n368 B.n367 10.6151
R846 B.n367 B.n366 10.6151
R847 B.n366 B.n77 10.6151
R848 B.n362 B.n77 10.6151
R849 B.n362 B.n361 10.6151
R850 B.n361 B.n360 10.6151
R851 B.n360 B.n79 10.6151
R852 B.n356 B.n79 10.6151
R853 B.n356 B.n355 10.6151
R854 B.n355 B.n354 10.6151
R855 B.n354 B.n81 10.6151
R856 B.n350 B.n81 10.6151
R857 B.n350 B.n349 10.6151
R858 B.n349 B.n348 10.6151
R859 B.n348 B.n83 10.6151
R860 B.n344 B.n83 10.6151
R861 B.n344 B.n343 10.6151
R862 B.n343 B.n342 10.6151
R863 B.n342 B.n85 10.6151
R864 B.n338 B.n85 10.6151
R865 B.n338 B.n337 10.6151
R866 B.n337 B.n336 10.6151
R867 B.n336 B.n87 10.6151
R868 B.n332 B.n87 10.6151
R869 B.n332 B.n331 10.6151
R870 B.n331 B.n330 10.6151
R871 B.n330 B.n89 10.6151
R872 B.n326 B.n89 10.6151
R873 B.n326 B.n325 10.6151
R874 B.n325 B.n324 10.6151
R875 B.n324 B.n91 10.6151
R876 B.n320 B.n91 10.6151
R877 B.n320 B.n319 10.6151
R878 B.n319 B.n318 10.6151
R879 B.n318 B.n93 10.6151
R880 B.n314 B.n93 10.6151
R881 B.n314 B.n313 10.6151
R882 B.n313 B.n312 10.6151
R883 B.n312 B.n95 10.6151
R884 B.n308 B.n95 10.6151
R885 B.n308 B.n307 10.6151
R886 B.n307 B.n306 10.6151
R887 B.n306 B.n97 10.6151
R888 B.n302 B.n97 10.6151
R889 B.n302 B.n301 10.6151
R890 B.n149 B.n1 10.6151
R891 B.n152 B.n149 10.6151
R892 B.n153 B.n152 10.6151
R893 B.n154 B.n153 10.6151
R894 B.n154 B.n147 10.6151
R895 B.n158 B.n147 10.6151
R896 B.n159 B.n158 10.6151
R897 B.n160 B.n159 10.6151
R898 B.n160 B.n145 10.6151
R899 B.n164 B.n145 10.6151
R900 B.n165 B.n164 10.6151
R901 B.n166 B.n165 10.6151
R902 B.n166 B.n143 10.6151
R903 B.n170 B.n143 10.6151
R904 B.n171 B.n170 10.6151
R905 B.n172 B.n171 10.6151
R906 B.n172 B.n141 10.6151
R907 B.n176 B.n141 10.6151
R908 B.n177 B.n176 10.6151
R909 B.n178 B.n177 10.6151
R910 B.n178 B.n139 10.6151
R911 B.n182 B.n139 10.6151
R912 B.n183 B.n182 10.6151
R913 B.n184 B.n183 10.6151
R914 B.n184 B.n137 10.6151
R915 B.n188 B.n137 10.6151
R916 B.n189 B.n188 10.6151
R917 B.n190 B.n189 10.6151
R918 B.n190 B.n135 10.6151
R919 B.n194 B.n135 10.6151
R920 B.n195 B.n194 10.6151
R921 B.n196 B.n195 10.6151
R922 B.n196 B.n133 10.6151
R923 B.n200 B.n133 10.6151
R924 B.n201 B.n200 10.6151
R925 B.n202 B.n201 10.6151
R926 B.n202 B.n131 10.6151
R927 B.n206 B.n131 10.6151
R928 B.n207 B.n206 10.6151
R929 B.n208 B.n207 10.6151
R930 B.n212 B.n129 10.6151
R931 B.n213 B.n212 10.6151
R932 B.n214 B.n213 10.6151
R933 B.n214 B.n127 10.6151
R934 B.n218 B.n127 10.6151
R935 B.n219 B.n218 10.6151
R936 B.n220 B.n219 10.6151
R937 B.n220 B.n125 10.6151
R938 B.n224 B.n125 10.6151
R939 B.n225 B.n224 10.6151
R940 B.n226 B.n225 10.6151
R941 B.n226 B.n123 10.6151
R942 B.n230 B.n123 10.6151
R943 B.n231 B.n230 10.6151
R944 B.n232 B.n231 10.6151
R945 B.n232 B.n121 10.6151
R946 B.n236 B.n121 10.6151
R947 B.n237 B.n236 10.6151
R948 B.n238 B.n237 10.6151
R949 B.n238 B.n119 10.6151
R950 B.n242 B.n119 10.6151
R951 B.n243 B.n242 10.6151
R952 B.n247 B.n243 10.6151
R953 B.n251 B.n117 10.6151
R954 B.n252 B.n251 10.6151
R955 B.n253 B.n252 10.6151
R956 B.n253 B.n115 10.6151
R957 B.n257 B.n115 10.6151
R958 B.n258 B.n257 10.6151
R959 B.n259 B.n258 10.6151
R960 B.n259 B.n113 10.6151
R961 B.n263 B.n113 10.6151
R962 B.n266 B.n265 10.6151
R963 B.n266 B.n109 10.6151
R964 B.n270 B.n109 10.6151
R965 B.n271 B.n270 10.6151
R966 B.n272 B.n271 10.6151
R967 B.n272 B.n107 10.6151
R968 B.n276 B.n107 10.6151
R969 B.n277 B.n276 10.6151
R970 B.n278 B.n277 10.6151
R971 B.n278 B.n105 10.6151
R972 B.n282 B.n105 10.6151
R973 B.n283 B.n282 10.6151
R974 B.n284 B.n283 10.6151
R975 B.n284 B.n103 10.6151
R976 B.n288 B.n103 10.6151
R977 B.n289 B.n288 10.6151
R978 B.n290 B.n289 10.6151
R979 B.n290 B.n101 10.6151
R980 B.n294 B.n101 10.6151
R981 B.n295 B.n294 10.6151
R982 B.n296 B.n295 10.6151
R983 B.n296 B.n99 10.6151
R984 B.n300 B.n99 10.6151
R985 B.n38 B.n34 9.36635
R986 B.n463 B.n462 9.36635
R987 B.n247 B.n246 9.36635
R988 B.n265 B.n264 9.36635
R989 B.n577 B.n0 8.11757
R990 B.n577 B.n1 8.11757
R991 B.n477 B.n38 1.24928
R992 B.n464 B.n463 1.24928
R993 B.n246 B.n117 1.24928
R994 B.n264 B.n263 1.24928
R995 VP.n14 VP.n11 161.3
R996 VP.n16 VP.n15 161.3
R997 VP.n17 VP.n10 161.3
R998 VP.n19 VP.n18 161.3
R999 VP.n20 VP.n9 161.3
R1000 VP.n23 VP.n22 161.3
R1001 VP.n24 VP.n8 161.3
R1002 VP.n26 VP.n25 161.3
R1003 VP.n27 VP.n7 161.3
R1004 VP.n52 VP.n0 161.3
R1005 VP.n51 VP.n50 161.3
R1006 VP.n49 VP.n1 161.3
R1007 VP.n48 VP.n47 161.3
R1008 VP.n45 VP.n2 161.3
R1009 VP.n44 VP.n43 161.3
R1010 VP.n42 VP.n3 161.3
R1011 VP.n41 VP.n40 161.3
R1012 VP.n39 VP.n4 161.3
R1013 VP.n37 VP.n36 161.3
R1014 VP.n35 VP.n5 161.3
R1015 VP.n34 VP.n33 161.3
R1016 VP.n32 VP.n6 161.3
R1017 VP.n12 VP.t1 106.222
R1018 VP.n31 VP.n30 90.2042
R1019 VP.n54 VP.n53 90.2042
R1020 VP.n29 VP.n28 90.2042
R1021 VP.n31 VP.t3 75.761
R1022 VP.n38 VP.t6 75.761
R1023 VP.n46 VP.t2 75.761
R1024 VP.n53 VP.t5 75.761
R1025 VP.n28 VP.t0 75.761
R1026 VP.n21 VP.t4 75.761
R1027 VP.n13 VP.t7 75.761
R1028 VP.n13 VP.n12 63.0337
R1029 VP.n33 VP.n5 56.5193
R1030 VP.n51 VP.n1 56.5193
R1031 VP.n26 VP.n8 56.5193
R1032 VP.n30 VP.n29 43.4314
R1033 VP.n40 VP.n3 40.4934
R1034 VP.n44 VP.n3 40.4934
R1035 VP.n19 VP.n10 40.4934
R1036 VP.n15 VP.n10 40.4934
R1037 VP.n33 VP.n32 24.4675
R1038 VP.n37 VP.n5 24.4675
R1039 VP.n40 VP.n39 24.4675
R1040 VP.n45 VP.n44 24.4675
R1041 VP.n47 VP.n1 24.4675
R1042 VP.n52 VP.n51 24.4675
R1043 VP.n27 VP.n26 24.4675
R1044 VP.n20 VP.n19 24.4675
R1045 VP.n22 VP.n8 24.4675
R1046 VP.n15 VP.n14 24.4675
R1047 VP.n32 VP.n31 20.5528
R1048 VP.n53 VP.n52 20.5528
R1049 VP.n28 VP.n27 20.5528
R1050 VP.n38 VP.n37 17.6167
R1051 VP.n47 VP.n46 17.6167
R1052 VP.n22 VP.n21 17.6167
R1053 VP.n12 VP.n11 13.2264
R1054 VP.n39 VP.n38 6.85126
R1055 VP.n46 VP.n45 6.85126
R1056 VP.n21 VP.n20 6.85126
R1057 VP.n14 VP.n13 6.85126
R1058 VP.n29 VP.n7 0.278367
R1059 VP.n30 VP.n6 0.278367
R1060 VP.n54 VP.n0 0.278367
R1061 VP.n16 VP.n11 0.189894
R1062 VP.n17 VP.n16 0.189894
R1063 VP.n18 VP.n17 0.189894
R1064 VP.n18 VP.n9 0.189894
R1065 VP.n23 VP.n9 0.189894
R1066 VP.n24 VP.n23 0.189894
R1067 VP.n25 VP.n24 0.189894
R1068 VP.n25 VP.n7 0.189894
R1069 VP.n34 VP.n6 0.189894
R1070 VP.n35 VP.n34 0.189894
R1071 VP.n36 VP.n35 0.189894
R1072 VP.n36 VP.n4 0.189894
R1073 VP.n41 VP.n4 0.189894
R1074 VP.n42 VP.n41 0.189894
R1075 VP.n43 VP.n42 0.189894
R1076 VP.n43 VP.n2 0.189894
R1077 VP.n48 VP.n2 0.189894
R1078 VP.n49 VP.n48 0.189894
R1079 VP.n50 VP.n49 0.189894
R1080 VP.n50 VP.n0 0.189894
R1081 VP VP.n54 0.153454
R1082 VDD1 VDD1.n0 93.187
R1083 VDD1.n3 VDD1.n2 93.0733
R1084 VDD1.n3 VDD1.n1 93.0733
R1085 VDD1.n5 VDD1.n4 92.145
R1086 VDD1.n5 VDD1.n3 38.4276
R1087 VDD1.n4 VDD1.t3 5.30311
R1088 VDD1.n4 VDD1.t7 5.30311
R1089 VDD1.n0 VDD1.t6 5.30311
R1090 VDD1.n0 VDD1.t0 5.30311
R1091 VDD1.n2 VDD1.t5 5.30311
R1092 VDD1.n2 VDD1.t2 5.30311
R1093 VDD1.n1 VDD1.t4 5.30311
R1094 VDD1.n1 VDD1.t1 5.30311
R1095 VDD1 VDD1.n5 0.925069
C0 VN VDD2 4.37231f
C1 B VTAIL 2.81322f
C2 VDD1 B 1.29405f
C3 VDD1 VTAIL 5.80023f
C4 w_n3250_n2194# VP 6.75088f
C5 B VDD2 1.36963f
C6 VDD2 VTAIL 5.85029f
C7 VDD1 VDD2 1.43976f
C8 VN VP 5.78259f
C9 B VP 1.70242f
C10 VP VTAIL 4.96278f
C11 VDD1 VP 4.67119f
C12 VDD2 VP 0.450588f
C13 VN w_n3250_n2194# 6.33088f
C14 B w_n3250_n2194# 7.48172f
C15 w_n3250_n2194# VTAIL 2.80718f
C16 VDD1 w_n3250_n2194# 1.58696f
C17 w_n3250_n2194# VDD2 1.6744f
C18 VN B 1.00182f
C19 VN VTAIL 4.94867f
C20 VDD1 VN 0.150637f
C21 VDD2 VSUBS 1.411722f
C22 VDD1 VSUBS 1.944491f
C23 VTAIL VSUBS 0.661811f
C24 VN VSUBS 5.62367f
C25 VP VSUBS 2.562262f
C26 B VSUBS 3.780173f
C27 w_n3250_n2194# VSUBS 88.959f
C28 VDD1.t6 VSUBS 0.12074f
C29 VDD1.t0 VSUBS 0.12074f
C30 VDD1.n0 VSUBS 0.828599f
C31 VDD1.t4 VSUBS 0.12074f
C32 VDD1.t1 VSUBS 0.12074f
C33 VDD1.n1 VSUBS 0.827736f
C34 VDD1.t5 VSUBS 0.12074f
C35 VDD1.t2 VSUBS 0.12074f
C36 VDD1.n2 VSUBS 0.827736f
C37 VDD1.n3 VSUBS 2.95854f
C38 VDD1.t3 VSUBS 0.12074f
C39 VDD1.t7 VSUBS 0.12074f
C40 VDD1.n4 VSUBS 0.821418f
C41 VDD1.n5 VSUBS 2.47701f
C42 VP.n0 VSUBS 0.056196f
C43 VP.t5 VSUBS 1.35025f
C44 VP.n1 VSUBS 0.065788f
C45 VP.n2 VSUBS 0.042625f
C46 VP.t2 VSUBS 1.35025f
C47 VP.n3 VSUBS 0.034458f
C48 VP.n4 VSUBS 0.042625f
C49 VP.t6 VSUBS 1.35025f
C50 VP.n5 VSUBS 0.065788f
C51 VP.n6 VSUBS 0.056196f
C52 VP.t3 VSUBS 1.35025f
C53 VP.n7 VSUBS 0.056196f
C54 VP.t0 VSUBS 1.35025f
C55 VP.n8 VSUBS 0.065788f
C56 VP.n9 VSUBS 0.042625f
C57 VP.t4 VSUBS 1.35025f
C58 VP.n10 VSUBS 0.034458f
C59 VP.n11 VSUBS 0.317204f
C60 VP.t7 VSUBS 1.35025f
C61 VP.t1 VSUBS 1.55684f
C62 VP.n12 VSUBS 0.620179f
C63 VP.n13 VSUBS 0.60715f
C64 VP.n14 VSUBS 0.051203f
C65 VP.n15 VSUBS 0.084716f
C66 VP.n16 VSUBS 0.042625f
C67 VP.n17 VSUBS 0.042625f
C68 VP.n18 VSUBS 0.042625f
C69 VP.n19 VSUBS 0.084716f
C70 VP.n20 VSUBS 0.051203f
C71 VP.n21 VSUBS 0.515185f
C72 VP.n22 VSUBS 0.06846f
C73 VP.n23 VSUBS 0.042625f
C74 VP.n24 VSUBS 0.042625f
C75 VP.n25 VSUBS 0.042625f
C76 VP.n26 VSUBS 0.058661f
C77 VP.n27 VSUBS 0.073166f
C78 VP.n28 VSUBS 0.644543f
C79 VP.n29 VSUBS 1.89357f
C80 VP.n30 VSUBS 1.92885f
C81 VP.n31 VSUBS 0.644543f
C82 VP.n32 VSUBS 0.073166f
C83 VP.n33 VSUBS 0.058661f
C84 VP.n34 VSUBS 0.042625f
C85 VP.n35 VSUBS 0.042625f
C86 VP.n36 VSUBS 0.042625f
C87 VP.n37 VSUBS 0.06846f
C88 VP.n38 VSUBS 0.515185f
C89 VP.n39 VSUBS 0.051203f
C90 VP.n40 VSUBS 0.084716f
C91 VP.n41 VSUBS 0.042625f
C92 VP.n42 VSUBS 0.042625f
C93 VP.n43 VSUBS 0.042625f
C94 VP.n44 VSUBS 0.084716f
C95 VP.n45 VSUBS 0.051203f
C96 VP.n46 VSUBS 0.515185f
C97 VP.n47 VSUBS 0.06846f
C98 VP.n48 VSUBS 0.042625f
C99 VP.n49 VSUBS 0.042625f
C100 VP.n50 VSUBS 0.042625f
C101 VP.n51 VSUBS 0.058661f
C102 VP.n52 VSUBS 0.073166f
C103 VP.n53 VSUBS 0.644543f
C104 VP.n54 VSUBS 0.050465f
C105 B.n0 VSUBS 0.007358f
C106 B.n1 VSUBS 0.007358f
C107 B.n2 VSUBS 0.010882f
C108 B.n3 VSUBS 0.008339f
C109 B.n4 VSUBS 0.008339f
C110 B.n5 VSUBS 0.008339f
C111 B.n6 VSUBS 0.008339f
C112 B.n7 VSUBS 0.008339f
C113 B.n8 VSUBS 0.008339f
C114 B.n9 VSUBS 0.008339f
C115 B.n10 VSUBS 0.008339f
C116 B.n11 VSUBS 0.008339f
C117 B.n12 VSUBS 0.008339f
C118 B.n13 VSUBS 0.008339f
C119 B.n14 VSUBS 0.008339f
C120 B.n15 VSUBS 0.008339f
C121 B.n16 VSUBS 0.008339f
C122 B.n17 VSUBS 0.008339f
C123 B.n18 VSUBS 0.008339f
C124 B.n19 VSUBS 0.008339f
C125 B.n20 VSUBS 0.008339f
C126 B.n21 VSUBS 0.008339f
C127 B.n22 VSUBS 0.02017f
C128 B.n23 VSUBS 0.008339f
C129 B.n24 VSUBS 0.008339f
C130 B.n25 VSUBS 0.008339f
C131 B.n26 VSUBS 0.008339f
C132 B.n27 VSUBS 0.008339f
C133 B.n28 VSUBS 0.008339f
C134 B.n29 VSUBS 0.008339f
C135 B.n30 VSUBS 0.008339f
C136 B.n31 VSUBS 0.008339f
C137 B.n32 VSUBS 0.008339f
C138 B.n33 VSUBS 0.008339f
C139 B.n34 VSUBS 0.007848f
C140 B.n35 VSUBS 0.008339f
C141 B.t1 VSUBS 0.214266f
C142 B.t2 VSUBS 0.233987f
C143 B.t0 VSUBS 0.66245f
C144 B.n36 VSUBS 0.131118f
C145 B.n37 VSUBS 0.081097f
C146 B.n38 VSUBS 0.019321f
C147 B.n39 VSUBS 0.008339f
C148 B.n40 VSUBS 0.008339f
C149 B.n41 VSUBS 0.008339f
C150 B.n42 VSUBS 0.008339f
C151 B.t10 VSUBS 0.214266f
C152 B.t11 VSUBS 0.233986f
C153 B.t9 VSUBS 0.66245f
C154 B.n43 VSUBS 0.13112f
C155 B.n44 VSUBS 0.081098f
C156 B.n45 VSUBS 0.008339f
C157 B.n46 VSUBS 0.008339f
C158 B.n47 VSUBS 0.008339f
C159 B.n48 VSUBS 0.008339f
C160 B.n49 VSUBS 0.008339f
C161 B.n50 VSUBS 0.008339f
C162 B.n51 VSUBS 0.008339f
C163 B.n52 VSUBS 0.008339f
C164 B.n53 VSUBS 0.008339f
C165 B.n54 VSUBS 0.008339f
C166 B.n55 VSUBS 0.008339f
C167 B.n56 VSUBS 0.021034f
C168 B.n57 VSUBS 0.008339f
C169 B.n58 VSUBS 0.008339f
C170 B.n59 VSUBS 0.008339f
C171 B.n60 VSUBS 0.008339f
C172 B.n61 VSUBS 0.008339f
C173 B.n62 VSUBS 0.008339f
C174 B.n63 VSUBS 0.008339f
C175 B.n64 VSUBS 0.008339f
C176 B.n65 VSUBS 0.008339f
C177 B.n66 VSUBS 0.008339f
C178 B.n67 VSUBS 0.008339f
C179 B.n68 VSUBS 0.008339f
C180 B.n69 VSUBS 0.008339f
C181 B.n70 VSUBS 0.008339f
C182 B.n71 VSUBS 0.008339f
C183 B.n72 VSUBS 0.008339f
C184 B.n73 VSUBS 0.008339f
C185 B.n74 VSUBS 0.008339f
C186 B.n75 VSUBS 0.008339f
C187 B.n76 VSUBS 0.008339f
C188 B.n77 VSUBS 0.008339f
C189 B.n78 VSUBS 0.008339f
C190 B.n79 VSUBS 0.008339f
C191 B.n80 VSUBS 0.008339f
C192 B.n81 VSUBS 0.008339f
C193 B.n82 VSUBS 0.008339f
C194 B.n83 VSUBS 0.008339f
C195 B.n84 VSUBS 0.008339f
C196 B.n85 VSUBS 0.008339f
C197 B.n86 VSUBS 0.008339f
C198 B.n87 VSUBS 0.008339f
C199 B.n88 VSUBS 0.008339f
C200 B.n89 VSUBS 0.008339f
C201 B.n90 VSUBS 0.008339f
C202 B.n91 VSUBS 0.008339f
C203 B.n92 VSUBS 0.008339f
C204 B.n93 VSUBS 0.008339f
C205 B.n94 VSUBS 0.008339f
C206 B.n95 VSUBS 0.008339f
C207 B.n96 VSUBS 0.008339f
C208 B.n97 VSUBS 0.008339f
C209 B.n98 VSUBS 0.02017f
C210 B.n99 VSUBS 0.008339f
C211 B.n100 VSUBS 0.008339f
C212 B.n101 VSUBS 0.008339f
C213 B.n102 VSUBS 0.008339f
C214 B.n103 VSUBS 0.008339f
C215 B.n104 VSUBS 0.008339f
C216 B.n105 VSUBS 0.008339f
C217 B.n106 VSUBS 0.008339f
C218 B.n107 VSUBS 0.008339f
C219 B.n108 VSUBS 0.008339f
C220 B.n109 VSUBS 0.008339f
C221 B.n110 VSUBS 0.008339f
C222 B.t5 VSUBS 0.214266f
C223 B.t4 VSUBS 0.233986f
C224 B.t3 VSUBS 0.66245f
C225 B.n111 VSUBS 0.13112f
C226 B.n112 VSUBS 0.081098f
C227 B.n113 VSUBS 0.008339f
C228 B.n114 VSUBS 0.008339f
C229 B.n115 VSUBS 0.008339f
C230 B.n116 VSUBS 0.008339f
C231 B.n117 VSUBS 0.00466f
C232 B.n118 VSUBS 0.008339f
C233 B.n119 VSUBS 0.008339f
C234 B.n120 VSUBS 0.008339f
C235 B.n121 VSUBS 0.008339f
C236 B.n122 VSUBS 0.008339f
C237 B.n123 VSUBS 0.008339f
C238 B.n124 VSUBS 0.008339f
C239 B.n125 VSUBS 0.008339f
C240 B.n126 VSUBS 0.008339f
C241 B.n127 VSUBS 0.008339f
C242 B.n128 VSUBS 0.008339f
C243 B.n129 VSUBS 0.021034f
C244 B.n130 VSUBS 0.008339f
C245 B.n131 VSUBS 0.008339f
C246 B.n132 VSUBS 0.008339f
C247 B.n133 VSUBS 0.008339f
C248 B.n134 VSUBS 0.008339f
C249 B.n135 VSUBS 0.008339f
C250 B.n136 VSUBS 0.008339f
C251 B.n137 VSUBS 0.008339f
C252 B.n138 VSUBS 0.008339f
C253 B.n139 VSUBS 0.008339f
C254 B.n140 VSUBS 0.008339f
C255 B.n141 VSUBS 0.008339f
C256 B.n142 VSUBS 0.008339f
C257 B.n143 VSUBS 0.008339f
C258 B.n144 VSUBS 0.008339f
C259 B.n145 VSUBS 0.008339f
C260 B.n146 VSUBS 0.008339f
C261 B.n147 VSUBS 0.008339f
C262 B.n148 VSUBS 0.008339f
C263 B.n149 VSUBS 0.008339f
C264 B.n150 VSUBS 0.008339f
C265 B.n151 VSUBS 0.008339f
C266 B.n152 VSUBS 0.008339f
C267 B.n153 VSUBS 0.008339f
C268 B.n154 VSUBS 0.008339f
C269 B.n155 VSUBS 0.008339f
C270 B.n156 VSUBS 0.008339f
C271 B.n157 VSUBS 0.008339f
C272 B.n158 VSUBS 0.008339f
C273 B.n159 VSUBS 0.008339f
C274 B.n160 VSUBS 0.008339f
C275 B.n161 VSUBS 0.008339f
C276 B.n162 VSUBS 0.008339f
C277 B.n163 VSUBS 0.008339f
C278 B.n164 VSUBS 0.008339f
C279 B.n165 VSUBS 0.008339f
C280 B.n166 VSUBS 0.008339f
C281 B.n167 VSUBS 0.008339f
C282 B.n168 VSUBS 0.008339f
C283 B.n169 VSUBS 0.008339f
C284 B.n170 VSUBS 0.008339f
C285 B.n171 VSUBS 0.008339f
C286 B.n172 VSUBS 0.008339f
C287 B.n173 VSUBS 0.008339f
C288 B.n174 VSUBS 0.008339f
C289 B.n175 VSUBS 0.008339f
C290 B.n176 VSUBS 0.008339f
C291 B.n177 VSUBS 0.008339f
C292 B.n178 VSUBS 0.008339f
C293 B.n179 VSUBS 0.008339f
C294 B.n180 VSUBS 0.008339f
C295 B.n181 VSUBS 0.008339f
C296 B.n182 VSUBS 0.008339f
C297 B.n183 VSUBS 0.008339f
C298 B.n184 VSUBS 0.008339f
C299 B.n185 VSUBS 0.008339f
C300 B.n186 VSUBS 0.008339f
C301 B.n187 VSUBS 0.008339f
C302 B.n188 VSUBS 0.008339f
C303 B.n189 VSUBS 0.008339f
C304 B.n190 VSUBS 0.008339f
C305 B.n191 VSUBS 0.008339f
C306 B.n192 VSUBS 0.008339f
C307 B.n193 VSUBS 0.008339f
C308 B.n194 VSUBS 0.008339f
C309 B.n195 VSUBS 0.008339f
C310 B.n196 VSUBS 0.008339f
C311 B.n197 VSUBS 0.008339f
C312 B.n198 VSUBS 0.008339f
C313 B.n199 VSUBS 0.008339f
C314 B.n200 VSUBS 0.008339f
C315 B.n201 VSUBS 0.008339f
C316 B.n202 VSUBS 0.008339f
C317 B.n203 VSUBS 0.008339f
C318 B.n204 VSUBS 0.008339f
C319 B.n205 VSUBS 0.008339f
C320 B.n206 VSUBS 0.008339f
C321 B.n207 VSUBS 0.008339f
C322 B.n208 VSUBS 0.02017f
C323 B.n209 VSUBS 0.02017f
C324 B.n210 VSUBS 0.021034f
C325 B.n211 VSUBS 0.008339f
C326 B.n212 VSUBS 0.008339f
C327 B.n213 VSUBS 0.008339f
C328 B.n214 VSUBS 0.008339f
C329 B.n215 VSUBS 0.008339f
C330 B.n216 VSUBS 0.008339f
C331 B.n217 VSUBS 0.008339f
C332 B.n218 VSUBS 0.008339f
C333 B.n219 VSUBS 0.008339f
C334 B.n220 VSUBS 0.008339f
C335 B.n221 VSUBS 0.008339f
C336 B.n222 VSUBS 0.008339f
C337 B.n223 VSUBS 0.008339f
C338 B.n224 VSUBS 0.008339f
C339 B.n225 VSUBS 0.008339f
C340 B.n226 VSUBS 0.008339f
C341 B.n227 VSUBS 0.008339f
C342 B.n228 VSUBS 0.008339f
C343 B.n229 VSUBS 0.008339f
C344 B.n230 VSUBS 0.008339f
C345 B.n231 VSUBS 0.008339f
C346 B.n232 VSUBS 0.008339f
C347 B.n233 VSUBS 0.008339f
C348 B.n234 VSUBS 0.008339f
C349 B.n235 VSUBS 0.008339f
C350 B.n236 VSUBS 0.008339f
C351 B.n237 VSUBS 0.008339f
C352 B.n238 VSUBS 0.008339f
C353 B.n239 VSUBS 0.008339f
C354 B.n240 VSUBS 0.008339f
C355 B.n241 VSUBS 0.008339f
C356 B.n242 VSUBS 0.008339f
C357 B.n243 VSUBS 0.008339f
C358 B.t8 VSUBS 0.214266f
C359 B.t7 VSUBS 0.233987f
C360 B.t6 VSUBS 0.66245f
C361 B.n244 VSUBS 0.131118f
C362 B.n245 VSUBS 0.081097f
C363 B.n246 VSUBS 0.019321f
C364 B.n247 VSUBS 0.007848f
C365 B.n248 VSUBS 0.008339f
C366 B.n249 VSUBS 0.008339f
C367 B.n250 VSUBS 0.008339f
C368 B.n251 VSUBS 0.008339f
C369 B.n252 VSUBS 0.008339f
C370 B.n253 VSUBS 0.008339f
C371 B.n254 VSUBS 0.008339f
C372 B.n255 VSUBS 0.008339f
C373 B.n256 VSUBS 0.008339f
C374 B.n257 VSUBS 0.008339f
C375 B.n258 VSUBS 0.008339f
C376 B.n259 VSUBS 0.008339f
C377 B.n260 VSUBS 0.008339f
C378 B.n261 VSUBS 0.008339f
C379 B.n262 VSUBS 0.008339f
C380 B.n263 VSUBS 0.00466f
C381 B.n264 VSUBS 0.019321f
C382 B.n265 VSUBS 0.007848f
C383 B.n266 VSUBS 0.008339f
C384 B.n267 VSUBS 0.008339f
C385 B.n268 VSUBS 0.008339f
C386 B.n269 VSUBS 0.008339f
C387 B.n270 VSUBS 0.008339f
C388 B.n271 VSUBS 0.008339f
C389 B.n272 VSUBS 0.008339f
C390 B.n273 VSUBS 0.008339f
C391 B.n274 VSUBS 0.008339f
C392 B.n275 VSUBS 0.008339f
C393 B.n276 VSUBS 0.008339f
C394 B.n277 VSUBS 0.008339f
C395 B.n278 VSUBS 0.008339f
C396 B.n279 VSUBS 0.008339f
C397 B.n280 VSUBS 0.008339f
C398 B.n281 VSUBS 0.008339f
C399 B.n282 VSUBS 0.008339f
C400 B.n283 VSUBS 0.008339f
C401 B.n284 VSUBS 0.008339f
C402 B.n285 VSUBS 0.008339f
C403 B.n286 VSUBS 0.008339f
C404 B.n287 VSUBS 0.008339f
C405 B.n288 VSUBS 0.008339f
C406 B.n289 VSUBS 0.008339f
C407 B.n290 VSUBS 0.008339f
C408 B.n291 VSUBS 0.008339f
C409 B.n292 VSUBS 0.008339f
C410 B.n293 VSUBS 0.008339f
C411 B.n294 VSUBS 0.008339f
C412 B.n295 VSUBS 0.008339f
C413 B.n296 VSUBS 0.008339f
C414 B.n297 VSUBS 0.008339f
C415 B.n298 VSUBS 0.008339f
C416 B.n299 VSUBS 0.021034f
C417 B.n300 VSUBS 0.020126f
C418 B.n301 VSUBS 0.021079f
C419 B.n302 VSUBS 0.008339f
C420 B.n303 VSUBS 0.008339f
C421 B.n304 VSUBS 0.008339f
C422 B.n305 VSUBS 0.008339f
C423 B.n306 VSUBS 0.008339f
C424 B.n307 VSUBS 0.008339f
C425 B.n308 VSUBS 0.008339f
C426 B.n309 VSUBS 0.008339f
C427 B.n310 VSUBS 0.008339f
C428 B.n311 VSUBS 0.008339f
C429 B.n312 VSUBS 0.008339f
C430 B.n313 VSUBS 0.008339f
C431 B.n314 VSUBS 0.008339f
C432 B.n315 VSUBS 0.008339f
C433 B.n316 VSUBS 0.008339f
C434 B.n317 VSUBS 0.008339f
C435 B.n318 VSUBS 0.008339f
C436 B.n319 VSUBS 0.008339f
C437 B.n320 VSUBS 0.008339f
C438 B.n321 VSUBS 0.008339f
C439 B.n322 VSUBS 0.008339f
C440 B.n323 VSUBS 0.008339f
C441 B.n324 VSUBS 0.008339f
C442 B.n325 VSUBS 0.008339f
C443 B.n326 VSUBS 0.008339f
C444 B.n327 VSUBS 0.008339f
C445 B.n328 VSUBS 0.008339f
C446 B.n329 VSUBS 0.008339f
C447 B.n330 VSUBS 0.008339f
C448 B.n331 VSUBS 0.008339f
C449 B.n332 VSUBS 0.008339f
C450 B.n333 VSUBS 0.008339f
C451 B.n334 VSUBS 0.008339f
C452 B.n335 VSUBS 0.008339f
C453 B.n336 VSUBS 0.008339f
C454 B.n337 VSUBS 0.008339f
C455 B.n338 VSUBS 0.008339f
C456 B.n339 VSUBS 0.008339f
C457 B.n340 VSUBS 0.008339f
C458 B.n341 VSUBS 0.008339f
C459 B.n342 VSUBS 0.008339f
C460 B.n343 VSUBS 0.008339f
C461 B.n344 VSUBS 0.008339f
C462 B.n345 VSUBS 0.008339f
C463 B.n346 VSUBS 0.008339f
C464 B.n347 VSUBS 0.008339f
C465 B.n348 VSUBS 0.008339f
C466 B.n349 VSUBS 0.008339f
C467 B.n350 VSUBS 0.008339f
C468 B.n351 VSUBS 0.008339f
C469 B.n352 VSUBS 0.008339f
C470 B.n353 VSUBS 0.008339f
C471 B.n354 VSUBS 0.008339f
C472 B.n355 VSUBS 0.008339f
C473 B.n356 VSUBS 0.008339f
C474 B.n357 VSUBS 0.008339f
C475 B.n358 VSUBS 0.008339f
C476 B.n359 VSUBS 0.008339f
C477 B.n360 VSUBS 0.008339f
C478 B.n361 VSUBS 0.008339f
C479 B.n362 VSUBS 0.008339f
C480 B.n363 VSUBS 0.008339f
C481 B.n364 VSUBS 0.008339f
C482 B.n365 VSUBS 0.008339f
C483 B.n366 VSUBS 0.008339f
C484 B.n367 VSUBS 0.008339f
C485 B.n368 VSUBS 0.008339f
C486 B.n369 VSUBS 0.008339f
C487 B.n370 VSUBS 0.008339f
C488 B.n371 VSUBS 0.008339f
C489 B.n372 VSUBS 0.008339f
C490 B.n373 VSUBS 0.008339f
C491 B.n374 VSUBS 0.008339f
C492 B.n375 VSUBS 0.008339f
C493 B.n376 VSUBS 0.008339f
C494 B.n377 VSUBS 0.008339f
C495 B.n378 VSUBS 0.008339f
C496 B.n379 VSUBS 0.008339f
C497 B.n380 VSUBS 0.008339f
C498 B.n381 VSUBS 0.008339f
C499 B.n382 VSUBS 0.008339f
C500 B.n383 VSUBS 0.008339f
C501 B.n384 VSUBS 0.008339f
C502 B.n385 VSUBS 0.008339f
C503 B.n386 VSUBS 0.008339f
C504 B.n387 VSUBS 0.008339f
C505 B.n388 VSUBS 0.008339f
C506 B.n389 VSUBS 0.008339f
C507 B.n390 VSUBS 0.008339f
C508 B.n391 VSUBS 0.008339f
C509 B.n392 VSUBS 0.008339f
C510 B.n393 VSUBS 0.008339f
C511 B.n394 VSUBS 0.008339f
C512 B.n395 VSUBS 0.008339f
C513 B.n396 VSUBS 0.008339f
C514 B.n397 VSUBS 0.008339f
C515 B.n398 VSUBS 0.008339f
C516 B.n399 VSUBS 0.008339f
C517 B.n400 VSUBS 0.008339f
C518 B.n401 VSUBS 0.008339f
C519 B.n402 VSUBS 0.008339f
C520 B.n403 VSUBS 0.008339f
C521 B.n404 VSUBS 0.008339f
C522 B.n405 VSUBS 0.008339f
C523 B.n406 VSUBS 0.008339f
C524 B.n407 VSUBS 0.008339f
C525 B.n408 VSUBS 0.008339f
C526 B.n409 VSUBS 0.008339f
C527 B.n410 VSUBS 0.008339f
C528 B.n411 VSUBS 0.008339f
C529 B.n412 VSUBS 0.008339f
C530 B.n413 VSUBS 0.008339f
C531 B.n414 VSUBS 0.008339f
C532 B.n415 VSUBS 0.008339f
C533 B.n416 VSUBS 0.008339f
C534 B.n417 VSUBS 0.008339f
C535 B.n418 VSUBS 0.008339f
C536 B.n419 VSUBS 0.008339f
C537 B.n420 VSUBS 0.008339f
C538 B.n421 VSUBS 0.008339f
C539 B.n422 VSUBS 0.008339f
C540 B.n423 VSUBS 0.008339f
C541 B.n424 VSUBS 0.008339f
C542 B.n425 VSUBS 0.02017f
C543 B.n426 VSUBS 0.02017f
C544 B.n427 VSUBS 0.021034f
C545 B.n428 VSUBS 0.008339f
C546 B.n429 VSUBS 0.008339f
C547 B.n430 VSUBS 0.008339f
C548 B.n431 VSUBS 0.008339f
C549 B.n432 VSUBS 0.008339f
C550 B.n433 VSUBS 0.008339f
C551 B.n434 VSUBS 0.008339f
C552 B.n435 VSUBS 0.008339f
C553 B.n436 VSUBS 0.008339f
C554 B.n437 VSUBS 0.008339f
C555 B.n438 VSUBS 0.008339f
C556 B.n439 VSUBS 0.008339f
C557 B.n440 VSUBS 0.008339f
C558 B.n441 VSUBS 0.008339f
C559 B.n442 VSUBS 0.008339f
C560 B.n443 VSUBS 0.008339f
C561 B.n444 VSUBS 0.008339f
C562 B.n445 VSUBS 0.008339f
C563 B.n446 VSUBS 0.008339f
C564 B.n447 VSUBS 0.008339f
C565 B.n448 VSUBS 0.008339f
C566 B.n449 VSUBS 0.008339f
C567 B.n450 VSUBS 0.008339f
C568 B.n451 VSUBS 0.008339f
C569 B.n452 VSUBS 0.008339f
C570 B.n453 VSUBS 0.008339f
C571 B.n454 VSUBS 0.008339f
C572 B.n455 VSUBS 0.008339f
C573 B.n456 VSUBS 0.008339f
C574 B.n457 VSUBS 0.008339f
C575 B.n458 VSUBS 0.008339f
C576 B.n459 VSUBS 0.008339f
C577 B.n460 VSUBS 0.008339f
C578 B.n461 VSUBS 0.008339f
C579 B.n462 VSUBS 0.007848f
C580 B.n463 VSUBS 0.019321f
C581 B.n464 VSUBS 0.00466f
C582 B.n465 VSUBS 0.008339f
C583 B.n466 VSUBS 0.008339f
C584 B.n467 VSUBS 0.008339f
C585 B.n468 VSUBS 0.008339f
C586 B.n469 VSUBS 0.008339f
C587 B.n470 VSUBS 0.008339f
C588 B.n471 VSUBS 0.008339f
C589 B.n472 VSUBS 0.008339f
C590 B.n473 VSUBS 0.008339f
C591 B.n474 VSUBS 0.008339f
C592 B.n475 VSUBS 0.008339f
C593 B.n476 VSUBS 0.008339f
C594 B.n477 VSUBS 0.00466f
C595 B.n478 VSUBS 0.008339f
C596 B.n479 VSUBS 0.008339f
C597 B.n480 VSUBS 0.008339f
C598 B.n481 VSUBS 0.008339f
C599 B.n482 VSUBS 0.008339f
C600 B.n483 VSUBS 0.008339f
C601 B.n484 VSUBS 0.008339f
C602 B.n485 VSUBS 0.008339f
C603 B.n486 VSUBS 0.008339f
C604 B.n487 VSUBS 0.008339f
C605 B.n488 VSUBS 0.008339f
C606 B.n489 VSUBS 0.008339f
C607 B.n490 VSUBS 0.008339f
C608 B.n491 VSUBS 0.008339f
C609 B.n492 VSUBS 0.008339f
C610 B.n493 VSUBS 0.008339f
C611 B.n494 VSUBS 0.008339f
C612 B.n495 VSUBS 0.008339f
C613 B.n496 VSUBS 0.008339f
C614 B.n497 VSUBS 0.008339f
C615 B.n498 VSUBS 0.008339f
C616 B.n499 VSUBS 0.008339f
C617 B.n500 VSUBS 0.008339f
C618 B.n501 VSUBS 0.008339f
C619 B.n502 VSUBS 0.008339f
C620 B.n503 VSUBS 0.008339f
C621 B.n504 VSUBS 0.008339f
C622 B.n505 VSUBS 0.008339f
C623 B.n506 VSUBS 0.008339f
C624 B.n507 VSUBS 0.008339f
C625 B.n508 VSUBS 0.008339f
C626 B.n509 VSUBS 0.008339f
C627 B.n510 VSUBS 0.008339f
C628 B.n511 VSUBS 0.008339f
C629 B.n512 VSUBS 0.008339f
C630 B.n513 VSUBS 0.021034f
C631 B.n514 VSUBS 0.021034f
C632 B.n515 VSUBS 0.02017f
C633 B.n516 VSUBS 0.008339f
C634 B.n517 VSUBS 0.008339f
C635 B.n518 VSUBS 0.008339f
C636 B.n519 VSUBS 0.008339f
C637 B.n520 VSUBS 0.008339f
C638 B.n521 VSUBS 0.008339f
C639 B.n522 VSUBS 0.008339f
C640 B.n523 VSUBS 0.008339f
C641 B.n524 VSUBS 0.008339f
C642 B.n525 VSUBS 0.008339f
C643 B.n526 VSUBS 0.008339f
C644 B.n527 VSUBS 0.008339f
C645 B.n528 VSUBS 0.008339f
C646 B.n529 VSUBS 0.008339f
C647 B.n530 VSUBS 0.008339f
C648 B.n531 VSUBS 0.008339f
C649 B.n532 VSUBS 0.008339f
C650 B.n533 VSUBS 0.008339f
C651 B.n534 VSUBS 0.008339f
C652 B.n535 VSUBS 0.008339f
C653 B.n536 VSUBS 0.008339f
C654 B.n537 VSUBS 0.008339f
C655 B.n538 VSUBS 0.008339f
C656 B.n539 VSUBS 0.008339f
C657 B.n540 VSUBS 0.008339f
C658 B.n541 VSUBS 0.008339f
C659 B.n542 VSUBS 0.008339f
C660 B.n543 VSUBS 0.008339f
C661 B.n544 VSUBS 0.008339f
C662 B.n545 VSUBS 0.008339f
C663 B.n546 VSUBS 0.008339f
C664 B.n547 VSUBS 0.008339f
C665 B.n548 VSUBS 0.008339f
C666 B.n549 VSUBS 0.008339f
C667 B.n550 VSUBS 0.008339f
C668 B.n551 VSUBS 0.008339f
C669 B.n552 VSUBS 0.008339f
C670 B.n553 VSUBS 0.008339f
C671 B.n554 VSUBS 0.008339f
C672 B.n555 VSUBS 0.008339f
C673 B.n556 VSUBS 0.008339f
C674 B.n557 VSUBS 0.008339f
C675 B.n558 VSUBS 0.008339f
C676 B.n559 VSUBS 0.008339f
C677 B.n560 VSUBS 0.008339f
C678 B.n561 VSUBS 0.008339f
C679 B.n562 VSUBS 0.008339f
C680 B.n563 VSUBS 0.008339f
C681 B.n564 VSUBS 0.008339f
C682 B.n565 VSUBS 0.008339f
C683 B.n566 VSUBS 0.008339f
C684 B.n567 VSUBS 0.008339f
C685 B.n568 VSUBS 0.008339f
C686 B.n569 VSUBS 0.008339f
C687 B.n570 VSUBS 0.008339f
C688 B.n571 VSUBS 0.008339f
C689 B.n572 VSUBS 0.008339f
C690 B.n573 VSUBS 0.008339f
C691 B.n574 VSUBS 0.008339f
C692 B.n575 VSUBS 0.010882f
C693 B.n576 VSUBS 0.011592f
C694 B.n577 VSUBS 0.023052f
C695 VTAIL.t12 VSUBS 0.136264f
C696 VTAIL.t14 VSUBS 0.136264f
C697 VTAIL.n0 VSUBS 0.830728f
C698 VTAIL.n1 VSUBS 0.682619f
C699 VTAIL.t8 VSUBS 1.13237f
C700 VTAIL.n2 VSUBS 0.78992f
C701 VTAIL.t0 VSUBS 1.13237f
C702 VTAIL.n3 VSUBS 0.78992f
C703 VTAIL.t1 VSUBS 0.136264f
C704 VTAIL.t5 VSUBS 0.136264f
C705 VTAIL.n4 VSUBS 0.830728f
C706 VTAIL.n5 VSUBS 0.8555f
C707 VTAIL.t2 VSUBS 1.13237f
C708 VTAIL.n6 VSUBS 1.78659f
C709 VTAIL.t11 VSUBS 1.13237f
C710 VTAIL.n7 VSUBS 1.78658f
C711 VTAIL.t10 VSUBS 0.136264f
C712 VTAIL.t15 VSUBS 0.136264f
C713 VTAIL.n8 VSUBS 0.830733f
C714 VTAIL.n9 VSUBS 0.855495f
C715 VTAIL.t13 VSUBS 1.13237f
C716 VTAIL.n10 VSUBS 0.789915f
C717 VTAIL.t6 VSUBS 1.13237f
C718 VTAIL.n11 VSUBS 0.789915f
C719 VTAIL.t3 VSUBS 0.136264f
C720 VTAIL.t4 VSUBS 0.136264f
C721 VTAIL.n12 VSUBS 0.830733f
C722 VTAIL.n13 VSUBS 0.855495f
C723 VTAIL.t7 VSUBS 1.13236f
C724 VTAIL.n14 VSUBS 1.78659f
C725 VTAIL.t9 VSUBS 1.13237f
C726 VTAIL.n15 VSUBS 1.78132f
C727 VDD2.t4 VSUBS 0.119488f
C728 VDD2.t5 VSUBS 0.119488f
C729 VDD2.n0 VSUBS 0.819152f
C730 VDD2.t1 VSUBS 0.119488f
C731 VDD2.t3 VSUBS 0.119488f
C732 VDD2.n1 VSUBS 0.819152f
C733 VDD2.n2 VSUBS 2.87591f
C734 VDD2.t7 VSUBS 0.119488f
C735 VDD2.t2 VSUBS 0.119488f
C736 VDD2.n3 VSUBS 0.812904f
C737 VDD2.n4 VSUBS 2.42141f
C738 VDD2.t0 VSUBS 0.119488f
C739 VDD2.t6 VSUBS 0.119488f
C740 VDD2.n5 VSUBS 0.819123f
C741 VN.n0 VSUBS 0.053784f
C742 VN.t6 VSUBS 1.29228f
C743 VN.n1 VSUBS 0.062963f
C744 VN.n2 VSUBS 0.040795f
C745 VN.t1 VSUBS 1.29228f
C746 VN.n3 VSUBS 0.032979f
C747 VN.n4 VSUBS 0.303587f
C748 VN.t3 VSUBS 1.29228f
C749 VN.t7 VSUBS 1.49f
C750 VN.n5 VSUBS 0.593554f
C751 VN.n6 VSUBS 0.581085f
C752 VN.n7 VSUBS 0.049005f
C753 VN.n8 VSUBS 0.081079f
C754 VN.n9 VSUBS 0.040795f
C755 VN.n10 VSUBS 0.040795f
C756 VN.n11 VSUBS 0.040795f
C757 VN.n12 VSUBS 0.081079f
C758 VN.n13 VSUBS 0.049005f
C759 VN.n14 VSUBS 0.493068f
C760 VN.n15 VSUBS 0.065521f
C761 VN.n16 VSUBS 0.040795f
C762 VN.n17 VSUBS 0.040795f
C763 VN.n18 VSUBS 0.040795f
C764 VN.n19 VSUBS 0.056143f
C765 VN.n20 VSUBS 0.070025f
C766 VN.n21 VSUBS 0.616873f
C767 VN.n22 VSUBS 0.048298f
C768 VN.n23 VSUBS 0.053784f
C769 VN.t4 VSUBS 1.29228f
C770 VN.n24 VSUBS 0.062963f
C771 VN.n25 VSUBS 0.040795f
C772 VN.t5 VSUBS 1.29228f
C773 VN.n26 VSUBS 0.032979f
C774 VN.n27 VSUBS 0.303587f
C775 VN.t0 VSUBS 1.29228f
C776 VN.t2 VSUBS 1.49f
C777 VN.n28 VSUBS 0.593554f
C778 VN.n29 VSUBS 0.581085f
C779 VN.n30 VSUBS 0.049005f
C780 VN.n31 VSUBS 0.081079f
C781 VN.n32 VSUBS 0.040795f
C782 VN.n33 VSUBS 0.040795f
C783 VN.n34 VSUBS 0.040795f
C784 VN.n35 VSUBS 0.081079f
C785 VN.n36 VSUBS 0.049005f
C786 VN.n37 VSUBS 0.493068f
C787 VN.n38 VSUBS 0.065521f
C788 VN.n39 VSUBS 0.040795f
C789 VN.n40 VSUBS 0.040795f
C790 VN.n41 VSUBS 0.040795f
C791 VN.n42 VSUBS 0.056143f
C792 VN.n43 VSUBS 0.070025f
C793 VN.n44 VSUBS 0.616873f
C794 VN.n45 VSUBS 1.83473f
.ends

