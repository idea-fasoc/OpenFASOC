* NGSPICE file created from diff_pair_sample_0811.ext - technology: sky130A

.subckt diff_pair_sample_0811 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t4 w_n2098_n2784# sky130_fd_pr__pfet_01v8 ad=1.4982 pd=9.41 as=3.5412 ps=18.94 w=9.08 l=1.08
X1 VDD2.t5 VN.t0 VTAIL.t2 w_n2098_n2784# sky130_fd_pr__pfet_01v8 ad=1.4982 pd=9.41 as=3.5412 ps=18.94 w=9.08 l=1.08
X2 VDD2.t4 VN.t1 VTAIL.t1 w_n2098_n2784# sky130_fd_pr__pfet_01v8 ad=3.5412 pd=18.94 as=1.4982 ps=9.41 w=9.08 l=1.08
X3 VDD2.t3 VN.t2 VTAIL.t0 w_n2098_n2784# sky130_fd_pr__pfet_01v8 ad=3.5412 pd=18.94 as=1.4982 ps=9.41 w=9.08 l=1.08
X4 VDD2.t2 VN.t3 VTAIL.t11 w_n2098_n2784# sky130_fd_pr__pfet_01v8 ad=1.4982 pd=9.41 as=3.5412 ps=18.94 w=9.08 l=1.08
X5 VTAIL.t10 VN.t4 VDD2.t1 w_n2098_n2784# sky130_fd_pr__pfet_01v8 ad=1.4982 pd=9.41 as=1.4982 ps=9.41 w=9.08 l=1.08
X6 VDD1.t4 VP.t1 VTAIL.t7 w_n2098_n2784# sky130_fd_pr__pfet_01v8 ad=1.4982 pd=9.41 as=3.5412 ps=18.94 w=9.08 l=1.08
X7 VTAIL.t5 VP.t2 VDD1.t3 w_n2098_n2784# sky130_fd_pr__pfet_01v8 ad=1.4982 pd=9.41 as=1.4982 ps=9.41 w=9.08 l=1.08
X8 VDD1.t2 VP.t3 VTAIL.t3 w_n2098_n2784# sky130_fd_pr__pfet_01v8 ad=3.5412 pd=18.94 as=1.4982 ps=9.41 w=9.08 l=1.08
X9 VDD1.t1 VP.t4 VTAIL.t6 w_n2098_n2784# sky130_fd_pr__pfet_01v8 ad=3.5412 pd=18.94 as=1.4982 ps=9.41 w=9.08 l=1.08
X10 B.t11 B.t9 B.t10 w_n2098_n2784# sky130_fd_pr__pfet_01v8 ad=3.5412 pd=18.94 as=0 ps=0 w=9.08 l=1.08
X11 B.t8 B.t6 B.t7 w_n2098_n2784# sky130_fd_pr__pfet_01v8 ad=3.5412 pd=18.94 as=0 ps=0 w=9.08 l=1.08
X12 B.t5 B.t3 B.t4 w_n2098_n2784# sky130_fd_pr__pfet_01v8 ad=3.5412 pd=18.94 as=0 ps=0 w=9.08 l=1.08
X13 VTAIL.t8 VP.t5 VDD1.t0 w_n2098_n2784# sky130_fd_pr__pfet_01v8 ad=1.4982 pd=9.41 as=1.4982 ps=9.41 w=9.08 l=1.08
X14 B.t2 B.t0 B.t1 w_n2098_n2784# sky130_fd_pr__pfet_01v8 ad=3.5412 pd=18.94 as=0 ps=0 w=9.08 l=1.08
X15 VTAIL.t9 VN.t5 VDD2.t0 w_n2098_n2784# sky130_fd_pr__pfet_01v8 ad=1.4982 pd=9.41 as=1.4982 ps=9.41 w=9.08 l=1.08
R0 VP.n3 VP.t3 261.94
R1 VP.n8 VP.t4 238.993
R2 VP.n14 VP.t0 238.993
R3 VP.n6 VP.t1 238.993
R4 VP.n12 VP.t5 202.619
R5 VP.n4 VP.t2 202.619
R6 VP.n5 VP.n2 161.3
R7 VP.n13 VP.n0 161.3
R8 VP.n12 VP.n11 161.3
R9 VP.n10 VP.n1 161.3
R10 VP.n7 VP.n6 80.6037
R11 VP.n15 VP.n14 80.6037
R12 VP.n9 VP.n8 80.6037
R13 VP.n8 VP.n1 50.1678
R14 VP.n14 VP.n13 50.1678
R15 VP.n6 VP.n5 50.1678
R16 VP.n9 VP.n7 40.6718
R17 VP.n4 VP.n3 32.6313
R18 VP.n3 VP.n2 28.168
R19 VP.n12 VP.n1 24.5923
R20 VP.n13 VP.n12 24.5923
R21 VP.n5 VP.n4 24.5923
R22 VP.n7 VP.n2 0.285035
R23 VP.n10 VP.n9 0.285035
R24 VP.n15 VP.n0 0.285035
R25 VP.n11 VP.n10 0.189894
R26 VP.n11 VP.n0 0.189894
R27 VP VP.n15 0.146778
R28 VTAIL.n7 VTAIL.t11 70.1854
R29 VTAIL.n11 VTAIL.t2 70.1851
R30 VTAIL.n2 VTAIL.t4 70.1851
R31 VTAIL.n10 VTAIL.t7 70.1851
R32 VTAIL.n9 VTAIL.n8 66.6055
R33 VTAIL.n6 VTAIL.n5 66.6055
R34 VTAIL.n1 VTAIL.n0 66.6053
R35 VTAIL.n4 VTAIL.n3 66.6053
R36 VTAIL.n6 VTAIL.n4 22.6255
R37 VTAIL.n11 VTAIL.n10 21.41
R38 VTAIL.n0 VTAIL.t0 3.58035
R39 VTAIL.n0 VTAIL.t9 3.58035
R40 VTAIL.n3 VTAIL.t6 3.58035
R41 VTAIL.n3 VTAIL.t8 3.58035
R42 VTAIL.n8 VTAIL.t3 3.58035
R43 VTAIL.n8 VTAIL.t5 3.58035
R44 VTAIL.n5 VTAIL.t1 3.58035
R45 VTAIL.n5 VTAIL.t10 3.58035
R46 VTAIL.n7 VTAIL.n6 1.21602
R47 VTAIL.n10 VTAIL.n9 1.21602
R48 VTAIL.n4 VTAIL.n2 1.21602
R49 VTAIL.n9 VTAIL.n7 1.07809
R50 VTAIL.n2 VTAIL.n1 1.07809
R51 VTAIL VTAIL.n11 0.853948
R52 VTAIL VTAIL.n1 0.362569
R53 VDD1 VDD1.t2 87.834
R54 VDD1.n1 VDD1.t1 87.7202
R55 VDD1.n1 VDD1.n0 83.5326
R56 VDD1.n3 VDD1.n2 83.2841
R57 VDD1.n3 VDD1.n1 36.6841
R58 VDD1.n2 VDD1.t3 3.58035
R59 VDD1.n2 VDD1.t4 3.58035
R60 VDD1.n0 VDD1.t0 3.58035
R61 VDD1.n0 VDD1.t5 3.58035
R62 VDD1 VDD1.n3 0.24619
R63 VN.n1 VN.t2 261.94
R64 VN.n7 VN.t3 261.94
R65 VN.n4 VN.t0 238.993
R66 VN.n10 VN.t1 238.993
R67 VN.n2 VN.t5 202.619
R68 VN.n8 VN.t4 202.619
R69 VN.n9 VN.n6 161.3
R70 VN.n3 VN.n0 161.3
R71 VN.n11 VN.n10 80.6037
R72 VN.n5 VN.n4 80.6037
R73 VN.n4 VN.n3 50.1678
R74 VN.n10 VN.n9 50.1678
R75 VN VN.n11 40.9574
R76 VN.n2 VN.n1 32.6313
R77 VN.n8 VN.n7 32.6313
R78 VN.n7 VN.n6 28.168
R79 VN.n1 VN.n0 28.168
R80 VN.n3 VN.n2 24.5923
R81 VN.n9 VN.n8 24.5923
R82 VN.n11 VN.n6 0.285035
R83 VN.n5 VN.n0 0.285035
R84 VN VN.n5 0.146778
R85 VDD2.n1 VDD2.t3 87.7202
R86 VDD2.n2 VDD2.t4 86.8642
R87 VDD2.n1 VDD2.n0 83.5326
R88 VDD2 VDD2.n3 83.5298
R89 VDD2.n2 VDD2.n1 35.4933
R90 VDD2.n3 VDD2.t1 3.58035
R91 VDD2.n3 VDD2.t2 3.58035
R92 VDD2.n0 VDD2.t0 3.58035
R93 VDD2.n0 VDD2.t5 3.58035
R94 VDD2 VDD2.n2 0.970328
R95 B.n285 B.n82 585
R96 B.n284 B.n283 585
R97 B.n282 B.n83 585
R98 B.n281 B.n280 585
R99 B.n279 B.n84 585
R100 B.n278 B.n277 585
R101 B.n276 B.n85 585
R102 B.n275 B.n274 585
R103 B.n273 B.n86 585
R104 B.n272 B.n271 585
R105 B.n270 B.n87 585
R106 B.n269 B.n268 585
R107 B.n267 B.n88 585
R108 B.n266 B.n265 585
R109 B.n264 B.n89 585
R110 B.n263 B.n262 585
R111 B.n261 B.n90 585
R112 B.n260 B.n259 585
R113 B.n258 B.n91 585
R114 B.n257 B.n256 585
R115 B.n255 B.n92 585
R116 B.n254 B.n253 585
R117 B.n252 B.n93 585
R118 B.n251 B.n250 585
R119 B.n249 B.n94 585
R120 B.n248 B.n247 585
R121 B.n246 B.n95 585
R122 B.n245 B.n244 585
R123 B.n243 B.n96 585
R124 B.n242 B.n241 585
R125 B.n240 B.n97 585
R126 B.n239 B.n238 585
R127 B.n237 B.n98 585
R128 B.n235 B.n234 585
R129 B.n233 B.n101 585
R130 B.n232 B.n231 585
R131 B.n230 B.n102 585
R132 B.n229 B.n228 585
R133 B.n227 B.n103 585
R134 B.n226 B.n225 585
R135 B.n224 B.n104 585
R136 B.n223 B.n222 585
R137 B.n221 B.n105 585
R138 B.n220 B.n219 585
R139 B.n215 B.n106 585
R140 B.n214 B.n213 585
R141 B.n212 B.n107 585
R142 B.n211 B.n210 585
R143 B.n209 B.n108 585
R144 B.n208 B.n207 585
R145 B.n206 B.n109 585
R146 B.n205 B.n204 585
R147 B.n203 B.n110 585
R148 B.n202 B.n201 585
R149 B.n200 B.n111 585
R150 B.n199 B.n198 585
R151 B.n197 B.n112 585
R152 B.n196 B.n195 585
R153 B.n194 B.n113 585
R154 B.n193 B.n192 585
R155 B.n191 B.n114 585
R156 B.n190 B.n189 585
R157 B.n188 B.n115 585
R158 B.n187 B.n186 585
R159 B.n185 B.n116 585
R160 B.n184 B.n183 585
R161 B.n182 B.n117 585
R162 B.n181 B.n180 585
R163 B.n179 B.n118 585
R164 B.n178 B.n177 585
R165 B.n176 B.n119 585
R166 B.n175 B.n174 585
R167 B.n173 B.n120 585
R168 B.n172 B.n171 585
R169 B.n170 B.n121 585
R170 B.n169 B.n168 585
R171 B.n287 B.n286 585
R172 B.n288 B.n81 585
R173 B.n290 B.n289 585
R174 B.n291 B.n80 585
R175 B.n293 B.n292 585
R176 B.n294 B.n79 585
R177 B.n296 B.n295 585
R178 B.n297 B.n78 585
R179 B.n299 B.n298 585
R180 B.n300 B.n77 585
R181 B.n302 B.n301 585
R182 B.n303 B.n76 585
R183 B.n305 B.n304 585
R184 B.n306 B.n75 585
R185 B.n308 B.n307 585
R186 B.n309 B.n74 585
R187 B.n311 B.n310 585
R188 B.n312 B.n73 585
R189 B.n314 B.n313 585
R190 B.n315 B.n72 585
R191 B.n317 B.n316 585
R192 B.n318 B.n71 585
R193 B.n320 B.n319 585
R194 B.n321 B.n70 585
R195 B.n323 B.n322 585
R196 B.n324 B.n69 585
R197 B.n326 B.n325 585
R198 B.n327 B.n68 585
R199 B.n329 B.n328 585
R200 B.n330 B.n67 585
R201 B.n332 B.n331 585
R202 B.n333 B.n66 585
R203 B.n335 B.n334 585
R204 B.n336 B.n65 585
R205 B.n338 B.n337 585
R206 B.n339 B.n64 585
R207 B.n341 B.n340 585
R208 B.n342 B.n63 585
R209 B.n344 B.n343 585
R210 B.n345 B.n62 585
R211 B.n347 B.n346 585
R212 B.n348 B.n61 585
R213 B.n350 B.n349 585
R214 B.n351 B.n60 585
R215 B.n353 B.n352 585
R216 B.n354 B.n59 585
R217 B.n356 B.n355 585
R218 B.n357 B.n58 585
R219 B.n359 B.n358 585
R220 B.n360 B.n57 585
R221 B.n475 B.n14 585
R222 B.n474 B.n473 585
R223 B.n472 B.n15 585
R224 B.n471 B.n470 585
R225 B.n469 B.n16 585
R226 B.n468 B.n467 585
R227 B.n466 B.n17 585
R228 B.n465 B.n464 585
R229 B.n463 B.n18 585
R230 B.n462 B.n461 585
R231 B.n460 B.n19 585
R232 B.n459 B.n458 585
R233 B.n457 B.n20 585
R234 B.n456 B.n455 585
R235 B.n454 B.n21 585
R236 B.n453 B.n452 585
R237 B.n451 B.n22 585
R238 B.n450 B.n449 585
R239 B.n448 B.n23 585
R240 B.n447 B.n446 585
R241 B.n445 B.n24 585
R242 B.n444 B.n443 585
R243 B.n442 B.n25 585
R244 B.n441 B.n440 585
R245 B.n439 B.n26 585
R246 B.n438 B.n437 585
R247 B.n436 B.n27 585
R248 B.n435 B.n434 585
R249 B.n433 B.n28 585
R250 B.n432 B.n431 585
R251 B.n430 B.n29 585
R252 B.n429 B.n428 585
R253 B.n427 B.n30 585
R254 B.n426 B.n425 585
R255 B.n424 B.n31 585
R256 B.n423 B.n422 585
R257 B.n421 B.n35 585
R258 B.n420 B.n419 585
R259 B.n418 B.n36 585
R260 B.n417 B.n416 585
R261 B.n415 B.n37 585
R262 B.n414 B.n413 585
R263 B.n412 B.n38 585
R264 B.n410 B.n409 585
R265 B.n408 B.n41 585
R266 B.n407 B.n406 585
R267 B.n405 B.n42 585
R268 B.n404 B.n403 585
R269 B.n402 B.n43 585
R270 B.n401 B.n400 585
R271 B.n399 B.n44 585
R272 B.n398 B.n397 585
R273 B.n396 B.n45 585
R274 B.n395 B.n394 585
R275 B.n393 B.n46 585
R276 B.n392 B.n391 585
R277 B.n390 B.n47 585
R278 B.n389 B.n388 585
R279 B.n387 B.n48 585
R280 B.n386 B.n385 585
R281 B.n384 B.n49 585
R282 B.n383 B.n382 585
R283 B.n381 B.n50 585
R284 B.n380 B.n379 585
R285 B.n378 B.n51 585
R286 B.n377 B.n376 585
R287 B.n375 B.n52 585
R288 B.n374 B.n373 585
R289 B.n372 B.n53 585
R290 B.n371 B.n370 585
R291 B.n369 B.n54 585
R292 B.n368 B.n367 585
R293 B.n366 B.n55 585
R294 B.n365 B.n364 585
R295 B.n363 B.n56 585
R296 B.n362 B.n361 585
R297 B.n477 B.n476 585
R298 B.n478 B.n13 585
R299 B.n480 B.n479 585
R300 B.n481 B.n12 585
R301 B.n483 B.n482 585
R302 B.n484 B.n11 585
R303 B.n486 B.n485 585
R304 B.n487 B.n10 585
R305 B.n489 B.n488 585
R306 B.n490 B.n9 585
R307 B.n492 B.n491 585
R308 B.n493 B.n8 585
R309 B.n495 B.n494 585
R310 B.n496 B.n7 585
R311 B.n498 B.n497 585
R312 B.n499 B.n6 585
R313 B.n501 B.n500 585
R314 B.n502 B.n5 585
R315 B.n504 B.n503 585
R316 B.n505 B.n4 585
R317 B.n507 B.n506 585
R318 B.n508 B.n3 585
R319 B.n510 B.n509 585
R320 B.n511 B.n0 585
R321 B.n2 B.n1 585
R322 B.n134 B.n133 585
R323 B.n136 B.n135 585
R324 B.n137 B.n132 585
R325 B.n139 B.n138 585
R326 B.n140 B.n131 585
R327 B.n142 B.n141 585
R328 B.n143 B.n130 585
R329 B.n145 B.n144 585
R330 B.n146 B.n129 585
R331 B.n148 B.n147 585
R332 B.n149 B.n128 585
R333 B.n151 B.n150 585
R334 B.n152 B.n127 585
R335 B.n154 B.n153 585
R336 B.n155 B.n126 585
R337 B.n157 B.n156 585
R338 B.n158 B.n125 585
R339 B.n160 B.n159 585
R340 B.n161 B.n124 585
R341 B.n163 B.n162 585
R342 B.n164 B.n123 585
R343 B.n166 B.n165 585
R344 B.n167 B.n122 585
R345 B.n169 B.n122 502.111
R346 B.n287 B.n82 502.111
R347 B.n361 B.n360 502.111
R348 B.n476 B.n475 502.111
R349 B.n216 B.t9 406.058
R350 B.n99 B.t6 406.058
R351 B.n39 B.t3 406.058
R352 B.n32 B.t0 406.058
R353 B.n513 B.n512 256.663
R354 B.n512 B.n511 235.042
R355 B.n512 B.n2 235.042
R356 B.n170 B.n169 163.367
R357 B.n171 B.n170 163.367
R358 B.n171 B.n120 163.367
R359 B.n175 B.n120 163.367
R360 B.n176 B.n175 163.367
R361 B.n177 B.n176 163.367
R362 B.n177 B.n118 163.367
R363 B.n181 B.n118 163.367
R364 B.n182 B.n181 163.367
R365 B.n183 B.n182 163.367
R366 B.n183 B.n116 163.367
R367 B.n187 B.n116 163.367
R368 B.n188 B.n187 163.367
R369 B.n189 B.n188 163.367
R370 B.n189 B.n114 163.367
R371 B.n193 B.n114 163.367
R372 B.n194 B.n193 163.367
R373 B.n195 B.n194 163.367
R374 B.n195 B.n112 163.367
R375 B.n199 B.n112 163.367
R376 B.n200 B.n199 163.367
R377 B.n201 B.n200 163.367
R378 B.n201 B.n110 163.367
R379 B.n205 B.n110 163.367
R380 B.n206 B.n205 163.367
R381 B.n207 B.n206 163.367
R382 B.n207 B.n108 163.367
R383 B.n211 B.n108 163.367
R384 B.n212 B.n211 163.367
R385 B.n213 B.n212 163.367
R386 B.n213 B.n106 163.367
R387 B.n220 B.n106 163.367
R388 B.n221 B.n220 163.367
R389 B.n222 B.n221 163.367
R390 B.n222 B.n104 163.367
R391 B.n226 B.n104 163.367
R392 B.n227 B.n226 163.367
R393 B.n228 B.n227 163.367
R394 B.n228 B.n102 163.367
R395 B.n232 B.n102 163.367
R396 B.n233 B.n232 163.367
R397 B.n234 B.n233 163.367
R398 B.n234 B.n98 163.367
R399 B.n239 B.n98 163.367
R400 B.n240 B.n239 163.367
R401 B.n241 B.n240 163.367
R402 B.n241 B.n96 163.367
R403 B.n245 B.n96 163.367
R404 B.n246 B.n245 163.367
R405 B.n247 B.n246 163.367
R406 B.n247 B.n94 163.367
R407 B.n251 B.n94 163.367
R408 B.n252 B.n251 163.367
R409 B.n253 B.n252 163.367
R410 B.n253 B.n92 163.367
R411 B.n257 B.n92 163.367
R412 B.n258 B.n257 163.367
R413 B.n259 B.n258 163.367
R414 B.n259 B.n90 163.367
R415 B.n263 B.n90 163.367
R416 B.n264 B.n263 163.367
R417 B.n265 B.n264 163.367
R418 B.n265 B.n88 163.367
R419 B.n269 B.n88 163.367
R420 B.n270 B.n269 163.367
R421 B.n271 B.n270 163.367
R422 B.n271 B.n86 163.367
R423 B.n275 B.n86 163.367
R424 B.n276 B.n275 163.367
R425 B.n277 B.n276 163.367
R426 B.n277 B.n84 163.367
R427 B.n281 B.n84 163.367
R428 B.n282 B.n281 163.367
R429 B.n283 B.n282 163.367
R430 B.n283 B.n82 163.367
R431 B.n360 B.n359 163.367
R432 B.n359 B.n58 163.367
R433 B.n355 B.n58 163.367
R434 B.n355 B.n354 163.367
R435 B.n354 B.n353 163.367
R436 B.n353 B.n60 163.367
R437 B.n349 B.n60 163.367
R438 B.n349 B.n348 163.367
R439 B.n348 B.n347 163.367
R440 B.n347 B.n62 163.367
R441 B.n343 B.n62 163.367
R442 B.n343 B.n342 163.367
R443 B.n342 B.n341 163.367
R444 B.n341 B.n64 163.367
R445 B.n337 B.n64 163.367
R446 B.n337 B.n336 163.367
R447 B.n336 B.n335 163.367
R448 B.n335 B.n66 163.367
R449 B.n331 B.n66 163.367
R450 B.n331 B.n330 163.367
R451 B.n330 B.n329 163.367
R452 B.n329 B.n68 163.367
R453 B.n325 B.n68 163.367
R454 B.n325 B.n324 163.367
R455 B.n324 B.n323 163.367
R456 B.n323 B.n70 163.367
R457 B.n319 B.n70 163.367
R458 B.n319 B.n318 163.367
R459 B.n318 B.n317 163.367
R460 B.n317 B.n72 163.367
R461 B.n313 B.n72 163.367
R462 B.n313 B.n312 163.367
R463 B.n312 B.n311 163.367
R464 B.n311 B.n74 163.367
R465 B.n307 B.n74 163.367
R466 B.n307 B.n306 163.367
R467 B.n306 B.n305 163.367
R468 B.n305 B.n76 163.367
R469 B.n301 B.n76 163.367
R470 B.n301 B.n300 163.367
R471 B.n300 B.n299 163.367
R472 B.n299 B.n78 163.367
R473 B.n295 B.n78 163.367
R474 B.n295 B.n294 163.367
R475 B.n294 B.n293 163.367
R476 B.n293 B.n80 163.367
R477 B.n289 B.n80 163.367
R478 B.n289 B.n288 163.367
R479 B.n288 B.n287 163.367
R480 B.n475 B.n474 163.367
R481 B.n474 B.n15 163.367
R482 B.n470 B.n15 163.367
R483 B.n470 B.n469 163.367
R484 B.n469 B.n468 163.367
R485 B.n468 B.n17 163.367
R486 B.n464 B.n17 163.367
R487 B.n464 B.n463 163.367
R488 B.n463 B.n462 163.367
R489 B.n462 B.n19 163.367
R490 B.n458 B.n19 163.367
R491 B.n458 B.n457 163.367
R492 B.n457 B.n456 163.367
R493 B.n456 B.n21 163.367
R494 B.n452 B.n21 163.367
R495 B.n452 B.n451 163.367
R496 B.n451 B.n450 163.367
R497 B.n450 B.n23 163.367
R498 B.n446 B.n23 163.367
R499 B.n446 B.n445 163.367
R500 B.n445 B.n444 163.367
R501 B.n444 B.n25 163.367
R502 B.n440 B.n25 163.367
R503 B.n440 B.n439 163.367
R504 B.n439 B.n438 163.367
R505 B.n438 B.n27 163.367
R506 B.n434 B.n27 163.367
R507 B.n434 B.n433 163.367
R508 B.n433 B.n432 163.367
R509 B.n432 B.n29 163.367
R510 B.n428 B.n29 163.367
R511 B.n428 B.n427 163.367
R512 B.n427 B.n426 163.367
R513 B.n426 B.n31 163.367
R514 B.n422 B.n31 163.367
R515 B.n422 B.n421 163.367
R516 B.n421 B.n420 163.367
R517 B.n420 B.n36 163.367
R518 B.n416 B.n36 163.367
R519 B.n416 B.n415 163.367
R520 B.n415 B.n414 163.367
R521 B.n414 B.n38 163.367
R522 B.n409 B.n38 163.367
R523 B.n409 B.n408 163.367
R524 B.n408 B.n407 163.367
R525 B.n407 B.n42 163.367
R526 B.n403 B.n42 163.367
R527 B.n403 B.n402 163.367
R528 B.n402 B.n401 163.367
R529 B.n401 B.n44 163.367
R530 B.n397 B.n44 163.367
R531 B.n397 B.n396 163.367
R532 B.n396 B.n395 163.367
R533 B.n395 B.n46 163.367
R534 B.n391 B.n46 163.367
R535 B.n391 B.n390 163.367
R536 B.n390 B.n389 163.367
R537 B.n389 B.n48 163.367
R538 B.n385 B.n48 163.367
R539 B.n385 B.n384 163.367
R540 B.n384 B.n383 163.367
R541 B.n383 B.n50 163.367
R542 B.n379 B.n50 163.367
R543 B.n379 B.n378 163.367
R544 B.n378 B.n377 163.367
R545 B.n377 B.n52 163.367
R546 B.n373 B.n52 163.367
R547 B.n373 B.n372 163.367
R548 B.n372 B.n371 163.367
R549 B.n371 B.n54 163.367
R550 B.n367 B.n54 163.367
R551 B.n367 B.n366 163.367
R552 B.n366 B.n365 163.367
R553 B.n365 B.n56 163.367
R554 B.n361 B.n56 163.367
R555 B.n476 B.n13 163.367
R556 B.n480 B.n13 163.367
R557 B.n481 B.n480 163.367
R558 B.n482 B.n481 163.367
R559 B.n482 B.n11 163.367
R560 B.n486 B.n11 163.367
R561 B.n487 B.n486 163.367
R562 B.n488 B.n487 163.367
R563 B.n488 B.n9 163.367
R564 B.n492 B.n9 163.367
R565 B.n493 B.n492 163.367
R566 B.n494 B.n493 163.367
R567 B.n494 B.n7 163.367
R568 B.n498 B.n7 163.367
R569 B.n499 B.n498 163.367
R570 B.n500 B.n499 163.367
R571 B.n500 B.n5 163.367
R572 B.n504 B.n5 163.367
R573 B.n505 B.n504 163.367
R574 B.n506 B.n505 163.367
R575 B.n506 B.n3 163.367
R576 B.n510 B.n3 163.367
R577 B.n511 B.n510 163.367
R578 B.n134 B.n2 163.367
R579 B.n135 B.n134 163.367
R580 B.n135 B.n132 163.367
R581 B.n139 B.n132 163.367
R582 B.n140 B.n139 163.367
R583 B.n141 B.n140 163.367
R584 B.n141 B.n130 163.367
R585 B.n145 B.n130 163.367
R586 B.n146 B.n145 163.367
R587 B.n147 B.n146 163.367
R588 B.n147 B.n128 163.367
R589 B.n151 B.n128 163.367
R590 B.n152 B.n151 163.367
R591 B.n153 B.n152 163.367
R592 B.n153 B.n126 163.367
R593 B.n157 B.n126 163.367
R594 B.n158 B.n157 163.367
R595 B.n159 B.n158 163.367
R596 B.n159 B.n124 163.367
R597 B.n163 B.n124 163.367
R598 B.n164 B.n163 163.367
R599 B.n165 B.n164 163.367
R600 B.n165 B.n122 163.367
R601 B.n99 B.t7 140.062
R602 B.n39 B.t5 140.062
R603 B.n216 B.t10 140.053
R604 B.n32 B.t2 140.053
R605 B.n100 B.t8 112.716
R606 B.n40 B.t4 112.716
R607 B.n217 B.t11 112.707
R608 B.n33 B.t1 112.707
R609 B.n218 B.n217 59.5399
R610 B.n236 B.n100 59.5399
R611 B.n411 B.n40 59.5399
R612 B.n34 B.n33 59.5399
R613 B.n477 B.n14 32.6249
R614 B.n362 B.n57 32.6249
R615 B.n286 B.n285 32.6249
R616 B.n168 B.n167 32.6249
R617 B.n217 B.n216 27.346
R618 B.n100 B.n99 27.346
R619 B.n40 B.n39 27.346
R620 B.n33 B.n32 27.346
R621 B B.n513 18.0485
R622 B.n478 B.n477 10.6151
R623 B.n479 B.n478 10.6151
R624 B.n479 B.n12 10.6151
R625 B.n483 B.n12 10.6151
R626 B.n484 B.n483 10.6151
R627 B.n485 B.n484 10.6151
R628 B.n485 B.n10 10.6151
R629 B.n489 B.n10 10.6151
R630 B.n490 B.n489 10.6151
R631 B.n491 B.n490 10.6151
R632 B.n491 B.n8 10.6151
R633 B.n495 B.n8 10.6151
R634 B.n496 B.n495 10.6151
R635 B.n497 B.n496 10.6151
R636 B.n497 B.n6 10.6151
R637 B.n501 B.n6 10.6151
R638 B.n502 B.n501 10.6151
R639 B.n503 B.n502 10.6151
R640 B.n503 B.n4 10.6151
R641 B.n507 B.n4 10.6151
R642 B.n508 B.n507 10.6151
R643 B.n509 B.n508 10.6151
R644 B.n509 B.n0 10.6151
R645 B.n473 B.n14 10.6151
R646 B.n473 B.n472 10.6151
R647 B.n472 B.n471 10.6151
R648 B.n471 B.n16 10.6151
R649 B.n467 B.n16 10.6151
R650 B.n467 B.n466 10.6151
R651 B.n466 B.n465 10.6151
R652 B.n465 B.n18 10.6151
R653 B.n461 B.n18 10.6151
R654 B.n461 B.n460 10.6151
R655 B.n460 B.n459 10.6151
R656 B.n459 B.n20 10.6151
R657 B.n455 B.n20 10.6151
R658 B.n455 B.n454 10.6151
R659 B.n454 B.n453 10.6151
R660 B.n453 B.n22 10.6151
R661 B.n449 B.n22 10.6151
R662 B.n449 B.n448 10.6151
R663 B.n448 B.n447 10.6151
R664 B.n447 B.n24 10.6151
R665 B.n443 B.n24 10.6151
R666 B.n443 B.n442 10.6151
R667 B.n442 B.n441 10.6151
R668 B.n441 B.n26 10.6151
R669 B.n437 B.n26 10.6151
R670 B.n437 B.n436 10.6151
R671 B.n436 B.n435 10.6151
R672 B.n435 B.n28 10.6151
R673 B.n431 B.n28 10.6151
R674 B.n431 B.n430 10.6151
R675 B.n430 B.n429 10.6151
R676 B.n429 B.n30 10.6151
R677 B.n425 B.n424 10.6151
R678 B.n424 B.n423 10.6151
R679 B.n423 B.n35 10.6151
R680 B.n419 B.n35 10.6151
R681 B.n419 B.n418 10.6151
R682 B.n418 B.n417 10.6151
R683 B.n417 B.n37 10.6151
R684 B.n413 B.n37 10.6151
R685 B.n413 B.n412 10.6151
R686 B.n410 B.n41 10.6151
R687 B.n406 B.n41 10.6151
R688 B.n406 B.n405 10.6151
R689 B.n405 B.n404 10.6151
R690 B.n404 B.n43 10.6151
R691 B.n400 B.n43 10.6151
R692 B.n400 B.n399 10.6151
R693 B.n399 B.n398 10.6151
R694 B.n398 B.n45 10.6151
R695 B.n394 B.n45 10.6151
R696 B.n394 B.n393 10.6151
R697 B.n393 B.n392 10.6151
R698 B.n392 B.n47 10.6151
R699 B.n388 B.n47 10.6151
R700 B.n388 B.n387 10.6151
R701 B.n387 B.n386 10.6151
R702 B.n386 B.n49 10.6151
R703 B.n382 B.n49 10.6151
R704 B.n382 B.n381 10.6151
R705 B.n381 B.n380 10.6151
R706 B.n380 B.n51 10.6151
R707 B.n376 B.n51 10.6151
R708 B.n376 B.n375 10.6151
R709 B.n375 B.n374 10.6151
R710 B.n374 B.n53 10.6151
R711 B.n370 B.n53 10.6151
R712 B.n370 B.n369 10.6151
R713 B.n369 B.n368 10.6151
R714 B.n368 B.n55 10.6151
R715 B.n364 B.n55 10.6151
R716 B.n364 B.n363 10.6151
R717 B.n363 B.n362 10.6151
R718 B.n358 B.n57 10.6151
R719 B.n358 B.n357 10.6151
R720 B.n357 B.n356 10.6151
R721 B.n356 B.n59 10.6151
R722 B.n352 B.n59 10.6151
R723 B.n352 B.n351 10.6151
R724 B.n351 B.n350 10.6151
R725 B.n350 B.n61 10.6151
R726 B.n346 B.n61 10.6151
R727 B.n346 B.n345 10.6151
R728 B.n345 B.n344 10.6151
R729 B.n344 B.n63 10.6151
R730 B.n340 B.n63 10.6151
R731 B.n340 B.n339 10.6151
R732 B.n339 B.n338 10.6151
R733 B.n338 B.n65 10.6151
R734 B.n334 B.n65 10.6151
R735 B.n334 B.n333 10.6151
R736 B.n333 B.n332 10.6151
R737 B.n332 B.n67 10.6151
R738 B.n328 B.n67 10.6151
R739 B.n328 B.n327 10.6151
R740 B.n327 B.n326 10.6151
R741 B.n326 B.n69 10.6151
R742 B.n322 B.n69 10.6151
R743 B.n322 B.n321 10.6151
R744 B.n321 B.n320 10.6151
R745 B.n320 B.n71 10.6151
R746 B.n316 B.n71 10.6151
R747 B.n316 B.n315 10.6151
R748 B.n315 B.n314 10.6151
R749 B.n314 B.n73 10.6151
R750 B.n310 B.n73 10.6151
R751 B.n310 B.n309 10.6151
R752 B.n309 B.n308 10.6151
R753 B.n308 B.n75 10.6151
R754 B.n304 B.n75 10.6151
R755 B.n304 B.n303 10.6151
R756 B.n303 B.n302 10.6151
R757 B.n302 B.n77 10.6151
R758 B.n298 B.n77 10.6151
R759 B.n298 B.n297 10.6151
R760 B.n297 B.n296 10.6151
R761 B.n296 B.n79 10.6151
R762 B.n292 B.n79 10.6151
R763 B.n292 B.n291 10.6151
R764 B.n291 B.n290 10.6151
R765 B.n290 B.n81 10.6151
R766 B.n286 B.n81 10.6151
R767 B.n133 B.n1 10.6151
R768 B.n136 B.n133 10.6151
R769 B.n137 B.n136 10.6151
R770 B.n138 B.n137 10.6151
R771 B.n138 B.n131 10.6151
R772 B.n142 B.n131 10.6151
R773 B.n143 B.n142 10.6151
R774 B.n144 B.n143 10.6151
R775 B.n144 B.n129 10.6151
R776 B.n148 B.n129 10.6151
R777 B.n149 B.n148 10.6151
R778 B.n150 B.n149 10.6151
R779 B.n150 B.n127 10.6151
R780 B.n154 B.n127 10.6151
R781 B.n155 B.n154 10.6151
R782 B.n156 B.n155 10.6151
R783 B.n156 B.n125 10.6151
R784 B.n160 B.n125 10.6151
R785 B.n161 B.n160 10.6151
R786 B.n162 B.n161 10.6151
R787 B.n162 B.n123 10.6151
R788 B.n166 B.n123 10.6151
R789 B.n167 B.n166 10.6151
R790 B.n168 B.n121 10.6151
R791 B.n172 B.n121 10.6151
R792 B.n173 B.n172 10.6151
R793 B.n174 B.n173 10.6151
R794 B.n174 B.n119 10.6151
R795 B.n178 B.n119 10.6151
R796 B.n179 B.n178 10.6151
R797 B.n180 B.n179 10.6151
R798 B.n180 B.n117 10.6151
R799 B.n184 B.n117 10.6151
R800 B.n185 B.n184 10.6151
R801 B.n186 B.n185 10.6151
R802 B.n186 B.n115 10.6151
R803 B.n190 B.n115 10.6151
R804 B.n191 B.n190 10.6151
R805 B.n192 B.n191 10.6151
R806 B.n192 B.n113 10.6151
R807 B.n196 B.n113 10.6151
R808 B.n197 B.n196 10.6151
R809 B.n198 B.n197 10.6151
R810 B.n198 B.n111 10.6151
R811 B.n202 B.n111 10.6151
R812 B.n203 B.n202 10.6151
R813 B.n204 B.n203 10.6151
R814 B.n204 B.n109 10.6151
R815 B.n208 B.n109 10.6151
R816 B.n209 B.n208 10.6151
R817 B.n210 B.n209 10.6151
R818 B.n210 B.n107 10.6151
R819 B.n214 B.n107 10.6151
R820 B.n215 B.n214 10.6151
R821 B.n219 B.n215 10.6151
R822 B.n223 B.n105 10.6151
R823 B.n224 B.n223 10.6151
R824 B.n225 B.n224 10.6151
R825 B.n225 B.n103 10.6151
R826 B.n229 B.n103 10.6151
R827 B.n230 B.n229 10.6151
R828 B.n231 B.n230 10.6151
R829 B.n231 B.n101 10.6151
R830 B.n235 B.n101 10.6151
R831 B.n238 B.n237 10.6151
R832 B.n238 B.n97 10.6151
R833 B.n242 B.n97 10.6151
R834 B.n243 B.n242 10.6151
R835 B.n244 B.n243 10.6151
R836 B.n244 B.n95 10.6151
R837 B.n248 B.n95 10.6151
R838 B.n249 B.n248 10.6151
R839 B.n250 B.n249 10.6151
R840 B.n250 B.n93 10.6151
R841 B.n254 B.n93 10.6151
R842 B.n255 B.n254 10.6151
R843 B.n256 B.n255 10.6151
R844 B.n256 B.n91 10.6151
R845 B.n260 B.n91 10.6151
R846 B.n261 B.n260 10.6151
R847 B.n262 B.n261 10.6151
R848 B.n262 B.n89 10.6151
R849 B.n266 B.n89 10.6151
R850 B.n267 B.n266 10.6151
R851 B.n268 B.n267 10.6151
R852 B.n268 B.n87 10.6151
R853 B.n272 B.n87 10.6151
R854 B.n273 B.n272 10.6151
R855 B.n274 B.n273 10.6151
R856 B.n274 B.n85 10.6151
R857 B.n278 B.n85 10.6151
R858 B.n279 B.n278 10.6151
R859 B.n280 B.n279 10.6151
R860 B.n280 B.n83 10.6151
R861 B.n284 B.n83 10.6151
R862 B.n285 B.n284 10.6151
R863 B.n34 B.n30 9.36635
R864 B.n411 B.n410 9.36635
R865 B.n219 B.n218 9.36635
R866 B.n237 B.n236 9.36635
R867 B.n513 B.n0 8.11757
R868 B.n513 B.n1 8.11757
R869 B.n425 B.n34 1.24928
R870 B.n412 B.n411 1.24928
R871 B.n218 B.n105 1.24928
R872 B.n236 B.n235 1.24928
C0 VP w_n2098_n2784# 3.81158f
C1 VDD2 VDD1 0.849792f
C2 VTAIL VDD1 7.04417f
C3 VP VDD1 4.22949f
C4 VDD2 B 1.49396f
C5 w_n2098_n2784# VN 3.54457f
C6 B VTAIL 2.39186f
C7 VP B 1.25169f
C8 VN VDD1 0.149055f
C9 VDD2 VTAIL 7.08341f
C10 w_n2098_n2784# VDD1 1.70194f
C11 VP VDD2 0.329701f
C12 VP VTAIL 3.97771f
C13 VN B 0.81355f
C14 w_n2098_n2784# B 6.75885f
C15 VDD2 VN 4.05205f
C16 VDD2 w_n2098_n2784# 1.73806f
C17 B VDD1 1.45605f
C18 VN VTAIL 3.96331f
C19 w_n2098_n2784# VTAIL 2.4764f
C20 VP VN 4.90527f
C21 VDD2 VSUBS 1.240255f
C22 VDD1 VSUBS 1.560142f
C23 VTAIL VSUBS 0.772206f
C24 VN VSUBS 4.45129f
C25 VP VSUBS 1.6752f
C26 B VSUBS 2.889476f
C27 w_n2098_n2784# VSUBS 72.2803f
C28 B.n0 VSUBS 0.006648f
C29 B.n1 VSUBS 0.006648f
C30 B.n2 VSUBS 0.009832f
C31 B.n3 VSUBS 0.007534f
C32 B.n4 VSUBS 0.007534f
C33 B.n5 VSUBS 0.007534f
C34 B.n6 VSUBS 0.007534f
C35 B.n7 VSUBS 0.007534f
C36 B.n8 VSUBS 0.007534f
C37 B.n9 VSUBS 0.007534f
C38 B.n10 VSUBS 0.007534f
C39 B.n11 VSUBS 0.007534f
C40 B.n12 VSUBS 0.007534f
C41 B.n13 VSUBS 0.007534f
C42 B.n14 VSUBS 0.018323f
C43 B.n15 VSUBS 0.007534f
C44 B.n16 VSUBS 0.007534f
C45 B.n17 VSUBS 0.007534f
C46 B.n18 VSUBS 0.007534f
C47 B.n19 VSUBS 0.007534f
C48 B.n20 VSUBS 0.007534f
C49 B.n21 VSUBS 0.007534f
C50 B.n22 VSUBS 0.007534f
C51 B.n23 VSUBS 0.007534f
C52 B.n24 VSUBS 0.007534f
C53 B.n25 VSUBS 0.007534f
C54 B.n26 VSUBS 0.007534f
C55 B.n27 VSUBS 0.007534f
C56 B.n28 VSUBS 0.007534f
C57 B.n29 VSUBS 0.007534f
C58 B.n30 VSUBS 0.007091f
C59 B.n31 VSUBS 0.007534f
C60 B.t1 VSUBS 0.307538f
C61 B.t2 VSUBS 0.319154f
C62 B.t0 VSUBS 0.458724f
C63 B.n32 VSUBS 0.137628f
C64 B.n33 VSUBS 0.07024f
C65 B.n34 VSUBS 0.017456f
C66 B.n35 VSUBS 0.007534f
C67 B.n36 VSUBS 0.007534f
C68 B.n37 VSUBS 0.007534f
C69 B.n38 VSUBS 0.007534f
C70 B.t4 VSUBS 0.307535f
C71 B.t5 VSUBS 0.319151f
C72 B.t3 VSUBS 0.458724f
C73 B.n39 VSUBS 0.137632f
C74 B.n40 VSUBS 0.070244f
C75 B.n41 VSUBS 0.007534f
C76 B.n42 VSUBS 0.007534f
C77 B.n43 VSUBS 0.007534f
C78 B.n44 VSUBS 0.007534f
C79 B.n45 VSUBS 0.007534f
C80 B.n46 VSUBS 0.007534f
C81 B.n47 VSUBS 0.007534f
C82 B.n48 VSUBS 0.007534f
C83 B.n49 VSUBS 0.007534f
C84 B.n50 VSUBS 0.007534f
C85 B.n51 VSUBS 0.007534f
C86 B.n52 VSUBS 0.007534f
C87 B.n53 VSUBS 0.007534f
C88 B.n54 VSUBS 0.007534f
C89 B.n55 VSUBS 0.007534f
C90 B.n56 VSUBS 0.007534f
C91 B.n57 VSUBS 0.016911f
C92 B.n58 VSUBS 0.007534f
C93 B.n59 VSUBS 0.007534f
C94 B.n60 VSUBS 0.007534f
C95 B.n61 VSUBS 0.007534f
C96 B.n62 VSUBS 0.007534f
C97 B.n63 VSUBS 0.007534f
C98 B.n64 VSUBS 0.007534f
C99 B.n65 VSUBS 0.007534f
C100 B.n66 VSUBS 0.007534f
C101 B.n67 VSUBS 0.007534f
C102 B.n68 VSUBS 0.007534f
C103 B.n69 VSUBS 0.007534f
C104 B.n70 VSUBS 0.007534f
C105 B.n71 VSUBS 0.007534f
C106 B.n72 VSUBS 0.007534f
C107 B.n73 VSUBS 0.007534f
C108 B.n74 VSUBS 0.007534f
C109 B.n75 VSUBS 0.007534f
C110 B.n76 VSUBS 0.007534f
C111 B.n77 VSUBS 0.007534f
C112 B.n78 VSUBS 0.007534f
C113 B.n79 VSUBS 0.007534f
C114 B.n80 VSUBS 0.007534f
C115 B.n81 VSUBS 0.007534f
C116 B.n82 VSUBS 0.018323f
C117 B.n83 VSUBS 0.007534f
C118 B.n84 VSUBS 0.007534f
C119 B.n85 VSUBS 0.007534f
C120 B.n86 VSUBS 0.007534f
C121 B.n87 VSUBS 0.007534f
C122 B.n88 VSUBS 0.007534f
C123 B.n89 VSUBS 0.007534f
C124 B.n90 VSUBS 0.007534f
C125 B.n91 VSUBS 0.007534f
C126 B.n92 VSUBS 0.007534f
C127 B.n93 VSUBS 0.007534f
C128 B.n94 VSUBS 0.007534f
C129 B.n95 VSUBS 0.007534f
C130 B.n96 VSUBS 0.007534f
C131 B.n97 VSUBS 0.007534f
C132 B.n98 VSUBS 0.007534f
C133 B.t8 VSUBS 0.307535f
C134 B.t7 VSUBS 0.319151f
C135 B.t6 VSUBS 0.458724f
C136 B.n99 VSUBS 0.137632f
C137 B.n100 VSUBS 0.070244f
C138 B.n101 VSUBS 0.007534f
C139 B.n102 VSUBS 0.007534f
C140 B.n103 VSUBS 0.007534f
C141 B.n104 VSUBS 0.007534f
C142 B.n105 VSUBS 0.00421f
C143 B.n106 VSUBS 0.007534f
C144 B.n107 VSUBS 0.007534f
C145 B.n108 VSUBS 0.007534f
C146 B.n109 VSUBS 0.007534f
C147 B.n110 VSUBS 0.007534f
C148 B.n111 VSUBS 0.007534f
C149 B.n112 VSUBS 0.007534f
C150 B.n113 VSUBS 0.007534f
C151 B.n114 VSUBS 0.007534f
C152 B.n115 VSUBS 0.007534f
C153 B.n116 VSUBS 0.007534f
C154 B.n117 VSUBS 0.007534f
C155 B.n118 VSUBS 0.007534f
C156 B.n119 VSUBS 0.007534f
C157 B.n120 VSUBS 0.007534f
C158 B.n121 VSUBS 0.007534f
C159 B.n122 VSUBS 0.016911f
C160 B.n123 VSUBS 0.007534f
C161 B.n124 VSUBS 0.007534f
C162 B.n125 VSUBS 0.007534f
C163 B.n126 VSUBS 0.007534f
C164 B.n127 VSUBS 0.007534f
C165 B.n128 VSUBS 0.007534f
C166 B.n129 VSUBS 0.007534f
C167 B.n130 VSUBS 0.007534f
C168 B.n131 VSUBS 0.007534f
C169 B.n132 VSUBS 0.007534f
C170 B.n133 VSUBS 0.007534f
C171 B.n134 VSUBS 0.007534f
C172 B.n135 VSUBS 0.007534f
C173 B.n136 VSUBS 0.007534f
C174 B.n137 VSUBS 0.007534f
C175 B.n138 VSUBS 0.007534f
C176 B.n139 VSUBS 0.007534f
C177 B.n140 VSUBS 0.007534f
C178 B.n141 VSUBS 0.007534f
C179 B.n142 VSUBS 0.007534f
C180 B.n143 VSUBS 0.007534f
C181 B.n144 VSUBS 0.007534f
C182 B.n145 VSUBS 0.007534f
C183 B.n146 VSUBS 0.007534f
C184 B.n147 VSUBS 0.007534f
C185 B.n148 VSUBS 0.007534f
C186 B.n149 VSUBS 0.007534f
C187 B.n150 VSUBS 0.007534f
C188 B.n151 VSUBS 0.007534f
C189 B.n152 VSUBS 0.007534f
C190 B.n153 VSUBS 0.007534f
C191 B.n154 VSUBS 0.007534f
C192 B.n155 VSUBS 0.007534f
C193 B.n156 VSUBS 0.007534f
C194 B.n157 VSUBS 0.007534f
C195 B.n158 VSUBS 0.007534f
C196 B.n159 VSUBS 0.007534f
C197 B.n160 VSUBS 0.007534f
C198 B.n161 VSUBS 0.007534f
C199 B.n162 VSUBS 0.007534f
C200 B.n163 VSUBS 0.007534f
C201 B.n164 VSUBS 0.007534f
C202 B.n165 VSUBS 0.007534f
C203 B.n166 VSUBS 0.007534f
C204 B.n167 VSUBS 0.016911f
C205 B.n168 VSUBS 0.018323f
C206 B.n169 VSUBS 0.018323f
C207 B.n170 VSUBS 0.007534f
C208 B.n171 VSUBS 0.007534f
C209 B.n172 VSUBS 0.007534f
C210 B.n173 VSUBS 0.007534f
C211 B.n174 VSUBS 0.007534f
C212 B.n175 VSUBS 0.007534f
C213 B.n176 VSUBS 0.007534f
C214 B.n177 VSUBS 0.007534f
C215 B.n178 VSUBS 0.007534f
C216 B.n179 VSUBS 0.007534f
C217 B.n180 VSUBS 0.007534f
C218 B.n181 VSUBS 0.007534f
C219 B.n182 VSUBS 0.007534f
C220 B.n183 VSUBS 0.007534f
C221 B.n184 VSUBS 0.007534f
C222 B.n185 VSUBS 0.007534f
C223 B.n186 VSUBS 0.007534f
C224 B.n187 VSUBS 0.007534f
C225 B.n188 VSUBS 0.007534f
C226 B.n189 VSUBS 0.007534f
C227 B.n190 VSUBS 0.007534f
C228 B.n191 VSUBS 0.007534f
C229 B.n192 VSUBS 0.007534f
C230 B.n193 VSUBS 0.007534f
C231 B.n194 VSUBS 0.007534f
C232 B.n195 VSUBS 0.007534f
C233 B.n196 VSUBS 0.007534f
C234 B.n197 VSUBS 0.007534f
C235 B.n198 VSUBS 0.007534f
C236 B.n199 VSUBS 0.007534f
C237 B.n200 VSUBS 0.007534f
C238 B.n201 VSUBS 0.007534f
C239 B.n202 VSUBS 0.007534f
C240 B.n203 VSUBS 0.007534f
C241 B.n204 VSUBS 0.007534f
C242 B.n205 VSUBS 0.007534f
C243 B.n206 VSUBS 0.007534f
C244 B.n207 VSUBS 0.007534f
C245 B.n208 VSUBS 0.007534f
C246 B.n209 VSUBS 0.007534f
C247 B.n210 VSUBS 0.007534f
C248 B.n211 VSUBS 0.007534f
C249 B.n212 VSUBS 0.007534f
C250 B.n213 VSUBS 0.007534f
C251 B.n214 VSUBS 0.007534f
C252 B.n215 VSUBS 0.007534f
C253 B.t11 VSUBS 0.307538f
C254 B.t10 VSUBS 0.319154f
C255 B.t9 VSUBS 0.458724f
C256 B.n216 VSUBS 0.137628f
C257 B.n217 VSUBS 0.07024f
C258 B.n218 VSUBS 0.017456f
C259 B.n219 VSUBS 0.007091f
C260 B.n220 VSUBS 0.007534f
C261 B.n221 VSUBS 0.007534f
C262 B.n222 VSUBS 0.007534f
C263 B.n223 VSUBS 0.007534f
C264 B.n224 VSUBS 0.007534f
C265 B.n225 VSUBS 0.007534f
C266 B.n226 VSUBS 0.007534f
C267 B.n227 VSUBS 0.007534f
C268 B.n228 VSUBS 0.007534f
C269 B.n229 VSUBS 0.007534f
C270 B.n230 VSUBS 0.007534f
C271 B.n231 VSUBS 0.007534f
C272 B.n232 VSUBS 0.007534f
C273 B.n233 VSUBS 0.007534f
C274 B.n234 VSUBS 0.007534f
C275 B.n235 VSUBS 0.00421f
C276 B.n236 VSUBS 0.017456f
C277 B.n237 VSUBS 0.007091f
C278 B.n238 VSUBS 0.007534f
C279 B.n239 VSUBS 0.007534f
C280 B.n240 VSUBS 0.007534f
C281 B.n241 VSUBS 0.007534f
C282 B.n242 VSUBS 0.007534f
C283 B.n243 VSUBS 0.007534f
C284 B.n244 VSUBS 0.007534f
C285 B.n245 VSUBS 0.007534f
C286 B.n246 VSUBS 0.007534f
C287 B.n247 VSUBS 0.007534f
C288 B.n248 VSUBS 0.007534f
C289 B.n249 VSUBS 0.007534f
C290 B.n250 VSUBS 0.007534f
C291 B.n251 VSUBS 0.007534f
C292 B.n252 VSUBS 0.007534f
C293 B.n253 VSUBS 0.007534f
C294 B.n254 VSUBS 0.007534f
C295 B.n255 VSUBS 0.007534f
C296 B.n256 VSUBS 0.007534f
C297 B.n257 VSUBS 0.007534f
C298 B.n258 VSUBS 0.007534f
C299 B.n259 VSUBS 0.007534f
C300 B.n260 VSUBS 0.007534f
C301 B.n261 VSUBS 0.007534f
C302 B.n262 VSUBS 0.007534f
C303 B.n263 VSUBS 0.007534f
C304 B.n264 VSUBS 0.007534f
C305 B.n265 VSUBS 0.007534f
C306 B.n266 VSUBS 0.007534f
C307 B.n267 VSUBS 0.007534f
C308 B.n268 VSUBS 0.007534f
C309 B.n269 VSUBS 0.007534f
C310 B.n270 VSUBS 0.007534f
C311 B.n271 VSUBS 0.007534f
C312 B.n272 VSUBS 0.007534f
C313 B.n273 VSUBS 0.007534f
C314 B.n274 VSUBS 0.007534f
C315 B.n275 VSUBS 0.007534f
C316 B.n276 VSUBS 0.007534f
C317 B.n277 VSUBS 0.007534f
C318 B.n278 VSUBS 0.007534f
C319 B.n279 VSUBS 0.007534f
C320 B.n280 VSUBS 0.007534f
C321 B.n281 VSUBS 0.007534f
C322 B.n282 VSUBS 0.007534f
C323 B.n283 VSUBS 0.007534f
C324 B.n284 VSUBS 0.007534f
C325 B.n285 VSUBS 0.017432f
C326 B.n286 VSUBS 0.017802f
C327 B.n287 VSUBS 0.016911f
C328 B.n288 VSUBS 0.007534f
C329 B.n289 VSUBS 0.007534f
C330 B.n290 VSUBS 0.007534f
C331 B.n291 VSUBS 0.007534f
C332 B.n292 VSUBS 0.007534f
C333 B.n293 VSUBS 0.007534f
C334 B.n294 VSUBS 0.007534f
C335 B.n295 VSUBS 0.007534f
C336 B.n296 VSUBS 0.007534f
C337 B.n297 VSUBS 0.007534f
C338 B.n298 VSUBS 0.007534f
C339 B.n299 VSUBS 0.007534f
C340 B.n300 VSUBS 0.007534f
C341 B.n301 VSUBS 0.007534f
C342 B.n302 VSUBS 0.007534f
C343 B.n303 VSUBS 0.007534f
C344 B.n304 VSUBS 0.007534f
C345 B.n305 VSUBS 0.007534f
C346 B.n306 VSUBS 0.007534f
C347 B.n307 VSUBS 0.007534f
C348 B.n308 VSUBS 0.007534f
C349 B.n309 VSUBS 0.007534f
C350 B.n310 VSUBS 0.007534f
C351 B.n311 VSUBS 0.007534f
C352 B.n312 VSUBS 0.007534f
C353 B.n313 VSUBS 0.007534f
C354 B.n314 VSUBS 0.007534f
C355 B.n315 VSUBS 0.007534f
C356 B.n316 VSUBS 0.007534f
C357 B.n317 VSUBS 0.007534f
C358 B.n318 VSUBS 0.007534f
C359 B.n319 VSUBS 0.007534f
C360 B.n320 VSUBS 0.007534f
C361 B.n321 VSUBS 0.007534f
C362 B.n322 VSUBS 0.007534f
C363 B.n323 VSUBS 0.007534f
C364 B.n324 VSUBS 0.007534f
C365 B.n325 VSUBS 0.007534f
C366 B.n326 VSUBS 0.007534f
C367 B.n327 VSUBS 0.007534f
C368 B.n328 VSUBS 0.007534f
C369 B.n329 VSUBS 0.007534f
C370 B.n330 VSUBS 0.007534f
C371 B.n331 VSUBS 0.007534f
C372 B.n332 VSUBS 0.007534f
C373 B.n333 VSUBS 0.007534f
C374 B.n334 VSUBS 0.007534f
C375 B.n335 VSUBS 0.007534f
C376 B.n336 VSUBS 0.007534f
C377 B.n337 VSUBS 0.007534f
C378 B.n338 VSUBS 0.007534f
C379 B.n339 VSUBS 0.007534f
C380 B.n340 VSUBS 0.007534f
C381 B.n341 VSUBS 0.007534f
C382 B.n342 VSUBS 0.007534f
C383 B.n343 VSUBS 0.007534f
C384 B.n344 VSUBS 0.007534f
C385 B.n345 VSUBS 0.007534f
C386 B.n346 VSUBS 0.007534f
C387 B.n347 VSUBS 0.007534f
C388 B.n348 VSUBS 0.007534f
C389 B.n349 VSUBS 0.007534f
C390 B.n350 VSUBS 0.007534f
C391 B.n351 VSUBS 0.007534f
C392 B.n352 VSUBS 0.007534f
C393 B.n353 VSUBS 0.007534f
C394 B.n354 VSUBS 0.007534f
C395 B.n355 VSUBS 0.007534f
C396 B.n356 VSUBS 0.007534f
C397 B.n357 VSUBS 0.007534f
C398 B.n358 VSUBS 0.007534f
C399 B.n359 VSUBS 0.007534f
C400 B.n360 VSUBS 0.016911f
C401 B.n361 VSUBS 0.018323f
C402 B.n362 VSUBS 0.018323f
C403 B.n363 VSUBS 0.007534f
C404 B.n364 VSUBS 0.007534f
C405 B.n365 VSUBS 0.007534f
C406 B.n366 VSUBS 0.007534f
C407 B.n367 VSUBS 0.007534f
C408 B.n368 VSUBS 0.007534f
C409 B.n369 VSUBS 0.007534f
C410 B.n370 VSUBS 0.007534f
C411 B.n371 VSUBS 0.007534f
C412 B.n372 VSUBS 0.007534f
C413 B.n373 VSUBS 0.007534f
C414 B.n374 VSUBS 0.007534f
C415 B.n375 VSUBS 0.007534f
C416 B.n376 VSUBS 0.007534f
C417 B.n377 VSUBS 0.007534f
C418 B.n378 VSUBS 0.007534f
C419 B.n379 VSUBS 0.007534f
C420 B.n380 VSUBS 0.007534f
C421 B.n381 VSUBS 0.007534f
C422 B.n382 VSUBS 0.007534f
C423 B.n383 VSUBS 0.007534f
C424 B.n384 VSUBS 0.007534f
C425 B.n385 VSUBS 0.007534f
C426 B.n386 VSUBS 0.007534f
C427 B.n387 VSUBS 0.007534f
C428 B.n388 VSUBS 0.007534f
C429 B.n389 VSUBS 0.007534f
C430 B.n390 VSUBS 0.007534f
C431 B.n391 VSUBS 0.007534f
C432 B.n392 VSUBS 0.007534f
C433 B.n393 VSUBS 0.007534f
C434 B.n394 VSUBS 0.007534f
C435 B.n395 VSUBS 0.007534f
C436 B.n396 VSUBS 0.007534f
C437 B.n397 VSUBS 0.007534f
C438 B.n398 VSUBS 0.007534f
C439 B.n399 VSUBS 0.007534f
C440 B.n400 VSUBS 0.007534f
C441 B.n401 VSUBS 0.007534f
C442 B.n402 VSUBS 0.007534f
C443 B.n403 VSUBS 0.007534f
C444 B.n404 VSUBS 0.007534f
C445 B.n405 VSUBS 0.007534f
C446 B.n406 VSUBS 0.007534f
C447 B.n407 VSUBS 0.007534f
C448 B.n408 VSUBS 0.007534f
C449 B.n409 VSUBS 0.007534f
C450 B.n410 VSUBS 0.007091f
C451 B.n411 VSUBS 0.017456f
C452 B.n412 VSUBS 0.00421f
C453 B.n413 VSUBS 0.007534f
C454 B.n414 VSUBS 0.007534f
C455 B.n415 VSUBS 0.007534f
C456 B.n416 VSUBS 0.007534f
C457 B.n417 VSUBS 0.007534f
C458 B.n418 VSUBS 0.007534f
C459 B.n419 VSUBS 0.007534f
C460 B.n420 VSUBS 0.007534f
C461 B.n421 VSUBS 0.007534f
C462 B.n422 VSUBS 0.007534f
C463 B.n423 VSUBS 0.007534f
C464 B.n424 VSUBS 0.007534f
C465 B.n425 VSUBS 0.00421f
C466 B.n426 VSUBS 0.007534f
C467 B.n427 VSUBS 0.007534f
C468 B.n428 VSUBS 0.007534f
C469 B.n429 VSUBS 0.007534f
C470 B.n430 VSUBS 0.007534f
C471 B.n431 VSUBS 0.007534f
C472 B.n432 VSUBS 0.007534f
C473 B.n433 VSUBS 0.007534f
C474 B.n434 VSUBS 0.007534f
C475 B.n435 VSUBS 0.007534f
C476 B.n436 VSUBS 0.007534f
C477 B.n437 VSUBS 0.007534f
C478 B.n438 VSUBS 0.007534f
C479 B.n439 VSUBS 0.007534f
C480 B.n440 VSUBS 0.007534f
C481 B.n441 VSUBS 0.007534f
C482 B.n442 VSUBS 0.007534f
C483 B.n443 VSUBS 0.007534f
C484 B.n444 VSUBS 0.007534f
C485 B.n445 VSUBS 0.007534f
C486 B.n446 VSUBS 0.007534f
C487 B.n447 VSUBS 0.007534f
C488 B.n448 VSUBS 0.007534f
C489 B.n449 VSUBS 0.007534f
C490 B.n450 VSUBS 0.007534f
C491 B.n451 VSUBS 0.007534f
C492 B.n452 VSUBS 0.007534f
C493 B.n453 VSUBS 0.007534f
C494 B.n454 VSUBS 0.007534f
C495 B.n455 VSUBS 0.007534f
C496 B.n456 VSUBS 0.007534f
C497 B.n457 VSUBS 0.007534f
C498 B.n458 VSUBS 0.007534f
C499 B.n459 VSUBS 0.007534f
C500 B.n460 VSUBS 0.007534f
C501 B.n461 VSUBS 0.007534f
C502 B.n462 VSUBS 0.007534f
C503 B.n463 VSUBS 0.007534f
C504 B.n464 VSUBS 0.007534f
C505 B.n465 VSUBS 0.007534f
C506 B.n466 VSUBS 0.007534f
C507 B.n467 VSUBS 0.007534f
C508 B.n468 VSUBS 0.007534f
C509 B.n469 VSUBS 0.007534f
C510 B.n470 VSUBS 0.007534f
C511 B.n471 VSUBS 0.007534f
C512 B.n472 VSUBS 0.007534f
C513 B.n473 VSUBS 0.007534f
C514 B.n474 VSUBS 0.007534f
C515 B.n475 VSUBS 0.018323f
C516 B.n476 VSUBS 0.016911f
C517 B.n477 VSUBS 0.016911f
C518 B.n478 VSUBS 0.007534f
C519 B.n479 VSUBS 0.007534f
C520 B.n480 VSUBS 0.007534f
C521 B.n481 VSUBS 0.007534f
C522 B.n482 VSUBS 0.007534f
C523 B.n483 VSUBS 0.007534f
C524 B.n484 VSUBS 0.007534f
C525 B.n485 VSUBS 0.007534f
C526 B.n486 VSUBS 0.007534f
C527 B.n487 VSUBS 0.007534f
C528 B.n488 VSUBS 0.007534f
C529 B.n489 VSUBS 0.007534f
C530 B.n490 VSUBS 0.007534f
C531 B.n491 VSUBS 0.007534f
C532 B.n492 VSUBS 0.007534f
C533 B.n493 VSUBS 0.007534f
C534 B.n494 VSUBS 0.007534f
C535 B.n495 VSUBS 0.007534f
C536 B.n496 VSUBS 0.007534f
C537 B.n497 VSUBS 0.007534f
C538 B.n498 VSUBS 0.007534f
C539 B.n499 VSUBS 0.007534f
C540 B.n500 VSUBS 0.007534f
C541 B.n501 VSUBS 0.007534f
C542 B.n502 VSUBS 0.007534f
C543 B.n503 VSUBS 0.007534f
C544 B.n504 VSUBS 0.007534f
C545 B.n505 VSUBS 0.007534f
C546 B.n506 VSUBS 0.007534f
C547 B.n507 VSUBS 0.007534f
C548 B.n508 VSUBS 0.007534f
C549 B.n509 VSUBS 0.007534f
C550 B.n510 VSUBS 0.007534f
C551 B.n511 VSUBS 0.009832f
C552 B.n512 VSUBS 0.010473f
C553 B.n513 VSUBS 0.020827f
C554 VDD2.t3 VSUBS 1.58366f
C555 VDD2.t0 VSUBS 0.160921f
C556 VDD2.t5 VSUBS 0.160921f
C557 VDD2.n0 VSUBS 1.20214f
C558 VDD2.n1 VSUBS 2.26625f
C559 VDD2.t4 VSUBS 1.57859f
C560 VDD2.n2 VSUBS 2.13495f
C561 VDD2.t1 VSUBS 0.160921f
C562 VDD2.t2 VSUBS 0.160921f
C563 VDD2.n3 VSUBS 1.20212f
C564 VN.n0 VSUBS 0.275062f
C565 VN.t5 VSUBS 1.31627f
C566 VN.t2 VSUBS 1.45022f
C567 VN.n1 VSUBS 0.563468f
C568 VN.n2 VSUBS 0.581327f
C569 VN.n3 VSUBS 0.063544f
C570 VN.t0 VSUBS 1.39803f
C571 VN.n4 VSUBS 0.583337f
C572 VN.n5 VSUBS 0.046565f
C573 VN.n6 VSUBS 0.275062f
C574 VN.t4 VSUBS 1.31627f
C575 VN.t3 VSUBS 1.45022f
C576 VN.n7 VSUBS 0.563468f
C577 VN.n8 VSUBS 0.581327f
C578 VN.n9 VSUBS 0.063544f
C579 VN.t1 VSUBS 1.39803f
C580 VN.n10 VSUBS 0.583337f
C581 VN.n11 VSUBS 1.98982f
C582 VDD1.t2 VSUBS 1.57278f
C583 VDD1.t1 VSUBS 1.57203f
C584 VDD1.t0 VSUBS 0.15974f
C585 VDD1.t5 VSUBS 0.15974f
C586 VDD1.n0 VSUBS 1.19332f
C587 VDD1.n1 VSUBS 2.32499f
C588 VDD1.t3 VSUBS 0.15974f
C589 VDD1.t4 VSUBS 0.15974f
C590 VDD1.n2 VSUBS 1.19183f
C591 VDD1.n3 VSUBS 2.10089f
C592 VTAIL.t0 VSUBS 0.211661f
C593 VTAIL.t9 VSUBS 0.211661f
C594 VTAIL.n0 VSUBS 1.45295f
C595 VTAIL.n1 VSUBS 0.732837f
C596 VTAIL.t4 VSUBS 1.93745f
C597 VTAIL.n2 VSUBS 0.906715f
C598 VTAIL.t6 VSUBS 0.211661f
C599 VTAIL.t8 VSUBS 0.211661f
C600 VTAIL.n3 VSUBS 1.45295f
C601 VTAIL.n4 VSUBS 2.08733f
C602 VTAIL.t1 VSUBS 0.211661f
C603 VTAIL.t10 VSUBS 0.211661f
C604 VTAIL.n5 VSUBS 1.45296f
C605 VTAIL.n6 VSUBS 2.08732f
C606 VTAIL.t11 VSUBS 1.93746f
C607 VTAIL.n7 VSUBS 0.90671f
C608 VTAIL.t3 VSUBS 0.211661f
C609 VTAIL.t5 VSUBS 0.211661f
C610 VTAIL.n8 VSUBS 1.45296f
C611 VTAIL.n9 VSUBS 0.813953f
C612 VTAIL.t7 VSUBS 1.93745f
C613 VTAIL.n10 VSUBS 2.06455f
C614 VTAIL.t2 VSUBS 1.93745f
C615 VTAIL.n11 VSUBS 2.03013f
C616 VP.n0 VSUBS 0.068243f
C617 VP.t5 VSUBS 1.35391f
C618 VP.n1 VSUBS 0.065361f
C619 VP.n2 VSUBS 0.282929f
C620 VP.t1 VSUBS 1.43801f
C621 VP.t2 VSUBS 1.35391f
C622 VP.t3 VSUBS 1.4917f
C623 VP.n3 VSUBS 0.579583f
C624 VP.n4 VSUBS 0.597952f
C625 VP.n5 VSUBS 0.065361f
C626 VP.n6 VSUBS 0.60002f
C627 VP.n7 VSUBS 2.01787f
C628 VP.t4 VSUBS 1.43801f
C629 VP.n8 VSUBS 0.60002f
C630 VP.n9 VSUBS 2.0632f
C631 VP.n10 VSUBS 0.068243f
C632 VP.n11 VSUBS 0.051143f
C633 VP.n12 VSUBS 0.563341f
C634 VP.n13 VSUBS 0.065361f
C635 VP.t0 VSUBS 1.43801f
C636 VP.n14 VSUBS 0.60002f
C637 VP.n15 VSUBS 0.047897f
.ends

