* NGSPICE file created from diff_pair_sample_0726.ext - technology: sky130A

.subckt diff_pair_sample_0726 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t12 VN.t0 VDD2.t6 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=1.58895 ps=9.96 w=9.63 l=3.05
X1 VTAIL.t11 VN.t1 VDD2.t8 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=1.58895 ps=9.96 w=9.63 l=3.05
X2 VDD2.t2 VN.t2 VTAIL.t10 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=3.7557 pd=20.04 as=1.58895 ps=9.96 w=9.63 l=3.05
X3 VDD1.t9 VP.t0 VTAIL.t2 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=3.7557 pd=20.04 as=1.58895 ps=9.96 w=9.63 l=3.05
X4 VDD2.t3 VN.t3 VTAIL.t9 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=3.7557 ps=20.04 w=9.63 l=3.05
X5 VDD1.t8 VP.t1 VTAIL.t1 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=3.7557 ps=20.04 w=9.63 l=3.05
X6 B.t11 B.t9 B.t10 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=3.7557 pd=20.04 as=0 ps=0 w=9.63 l=3.05
X7 VTAIL.t8 VN.t4 VDD2.t5 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=1.58895 ps=9.96 w=9.63 l=3.05
X8 VDD1.t7 VP.t2 VTAIL.t13 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=1.58895 ps=9.96 w=9.63 l=3.05
X9 VDD2.t1 VN.t5 VTAIL.t7 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=1.58895 ps=9.96 w=9.63 l=3.05
X10 VDD2.t9 VN.t6 VTAIL.t6 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=3.7557 ps=20.04 w=9.63 l=3.05
X11 B.t8 B.t6 B.t7 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=3.7557 pd=20.04 as=0 ps=0 w=9.63 l=3.05
X12 VTAIL.t18 VP.t3 VDD1.t6 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=1.58895 ps=9.96 w=9.63 l=3.05
X13 VTAIL.t5 VN.t7 VDD2.t0 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=1.58895 ps=9.96 w=9.63 l=3.05
X14 VDD1.t5 VP.t4 VTAIL.t15 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=1.58895 ps=9.96 w=9.63 l=3.05
X15 B.t5 B.t3 B.t4 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=3.7557 pd=20.04 as=0 ps=0 w=9.63 l=3.05
X16 VDD2.t7 VN.t8 VTAIL.t4 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=1.58895 ps=9.96 w=9.63 l=3.05
X17 VDD1.t4 VP.t5 VTAIL.t17 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=3.7557 ps=20.04 w=9.63 l=3.05
X18 VDD1.t3 VP.t6 VTAIL.t0 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=3.7557 pd=20.04 as=1.58895 ps=9.96 w=9.63 l=3.05
X19 VTAIL.t14 VP.t7 VDD1.t2 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=1.58895 ps=9.96 w=9.63 l=3.05
X20 VDD2.t4 VN.t9 VTAIL.t3 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=3.7557 pd=20.04 as=1.58895 ps=9.96 w=9.63 l=3.05
X21 B.t2 B.t0 B.t1 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=3.7557 pd=20.04 as=0 ps=0 w=9.63 l=3.05
X22 VTAIL.t19 VP.t8 VDD1.t1 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=1.58895 ps=9.96 w=9.63 l=3.05
X23 VTAIL.t16 VP.t9 VDD1.t0 w_n5026_n2894# sky130_fd_pr__pfet_01v8 ad=1.58895 pd=9.96 as=1.58895 ps=9.96 w=9.63 l=3.05
R0 VN.n93 VN.n48 161.3
R1 VN.n92 VN.n91 161.3
R2 VN.n90 VN.n49 161.3
R3 VN.n89 VN.n88 161.3
R4 VN.n87 VN.n50 161.3
R5 VN.n86 VN.n85 161.3
R6 VN.n84 VN.n51 161.3
R7 VN.n83 VN.n82 161.3
R8 VN.n81 VN.n52 161.3
R9 VN.n80 VN.n79 161.3
R10 VN.n78 VN.n54 161.3
R11 VN.n77 VN.n76 161.3
R12 VN.n75 VN.n55 161.3
R13 VN.n74 VN.n73 161.3
R14 VN.n72 VN.n71 161.3
R15 VN.n70 VN.n57 161.3
R16 VN.n69 VN.n68 161.3
R17 VN.n67 VN.n58 161.3
R18 VN.n66 VN.n65 161.3
R19 VN.n64 VN.n59 161.3
R20 VN.n63 VN.n62 161.3
R21 VN.n45 VN.n0 161.3
R22 VN.n44 VN.n43 161.3
R23 VN.n42 VN.n1 161.3
R24 VN.n41 VN.n40 161.3
R25 VN.n39 VN.n2 161.3
R26 VN.n38 VN.n37 161.3
R27 VN.n36 VN.n3 161.3
R28 VN.n35 VN.n34 161.3
R29 VN.n32 VN.n4 161.3
R30 VN.n31 VN.n30 161.3
R31 VN.n29 VN.n5 161.3
R32 VN.n28 VN.n27 161.3
R33 VN.n26 VN.n6 161.3
R34 VN.n25 VN.n24 161.3
R35 VN.n23 VN.n22 161.3
R36 VN.n21 VN.n8 161.3
R37 VN.n20 VN.n19 161.3
R38 VN.n18 VN.n9 161.3
R39 VN.n17 VN.n16 161.3
R40 VN.n15 VN.n10 161.3
R41 VN.n14 VN.n13 161.3
R42 VN.n47 VN.n46 110.267
R43 VN.n95 VN.n94 110.267
R44 VN.n12 VN.t2 108.037
R45 VN.n61 VN.t6 108.037
R46 VN.n11 VN.t7 76.0933
R47 VN.n7 VN.t5 76.0933
R48 VN.n33 VN.t4 76.0933
R49 VN.n46 VN.t3 76.0933
R50 VN.n60 VN.t0 76.0933
R51 VN.n56 VN.t8 76.0933
R52 VN.n53 VN.t1 76.0933
R53 VN.n94 VN.t9 76.0933
R54 VN.n12 VN.n11 67.6363
R55 VN.n61 VN.n60 67.6363
R56 VN.n40 VN.n39 56.5193
R57 VN.n88 VN.n87 56.5193
R58 VN VN.n95 54.0285
R59 VN.n20 VN.n9 46.321
R60 VN.n27 VN.n5 46.321
R61 VN.n69 VN.n58 46.321
R62 VN.n76 VN.n54 46.321
R63 VN.n16 VN.n9 34.6658
R64 VN.n31 VN.n5 34.6658
R65 VN.n65 VN.n58 34.6658
R66 VN.n80 VN.n54 34.6658
R67 VN.n15 VN.n14 24.4675
R68 VN.n16 VN.n15 24.4675
R69 VN.n21 VN.n20 24.4675
R70 VN.n22 VN.n21 24.4675
R71 VN.n26 VN.n25 24.4675
R72 VN.n27 VN.n26 24.4675
R73 VN.n32 VN.n31 24.4675
R74 VN.n34 VN.n32 24.4675
R75 VN.n38 VN.n3 24.4675
R76 VN.n39 VN.n38 24.4675
R77 VN.n40 VN.n1 24.4675
R78 VN.n44 VN.n1 24.4675
R79 VN.n45 VN.n44 24.4675
R80 VN.n65 VN.n64 24.4675
R81 VN.n64 VN.n63 24.4675
R82 VN.n76 VN.n75 24.4675
R83 VN.n75 VN.n74 24.4675
R84 VN.n71 VN.n70 24.4675
R85 VN.n70 VN.n69 24.4675
R86 VN.n87 VN.n86 24.4675
R87 VN.n86 VN.n51 24.4675
R88 VN.n82 VN.n81 24.4675
R89 VN.n81 VN.n80 24.4675
R90 VN.n93 VN.n92 24.4675
R91 VN.n92 VN.n49 24.4675
R92 VN.n88 VN.n49 24.4675
R93 VN.n33 VN.n3 18.1061
R94 VN.n53 VN.n51 18.1061
R95 VN.n22 VN.n7 12.234
R96 VN.n25 VN.n7 12.234
R97 VN.n74 VN.n56 12.234
R98 VN.n71 VN.n56 12.234
R99 VN.n14 VN.n11 6.36192
R100 VN.n34 VN.n33 6.36192
R101 VN.n63 VN.n60 6.36192
R102 VN.n82 VN.n53 6.36192
R103 VN.n62 VN.n61 5.21216
R104 VN.n13 VN.n12 5.21216
R105 VN.n46 VN.n45 0.48984
R106 VN.n94 VN.n93 0.48984
R107 VN.n95 VN.n48 0.278367
R108 VN.n47 VN.n0 0.278367
R109 VN.n91 VN.n48 0.189894
R110 VN.n91 VN.n90 0.189894
R111 VN.n90 VN.n89 0.189894
R112 VN.n89 VN.n50 0.189894
R113 VN.n85 VN.n50 0.189894
R114 VN.n85 VN.n84 0.189894
R115 VN.n84 VN.n83 0.189894
R116 VN.n83 VN.n52 0.189894
R117 VN.n79 VN.n52 0.189894
R118 VN.n79 VN.n78 0.189894
R119 VN.n78 VN.n77 0.189894
R120 VN.n77 VN.n55 0.189894
R121 VN.n73 VN.n55 0.189894
R122 VN.n73 VN.n72 0.189894
R123 VN.n72 VN.n57 0.189894
R124 VN.n68 VN.n57 0.189894
R125 VN.n68 VN.n67 0.189894
R126 VN.n67 VN.n66 0.189894
R127 VN.n66 VN.n59 0.189894
R128 VN.n62 VN.n59 0.189894
R129 VN.n13 VN.n10 0.189894
R130 VN.n17 VN.n10 0.189894
R131 VN.n18 VN.n17 0.189894
R132 VN.n19 VN.n18 0.189894
R133 VN.n19 VN.n8 0.189894
R134 VN.n23 VN.n8 0.189894
R135 VN.n24 VN.n23 0.189894
R136 VN.n24 VN.n6 0.189894
R137 VN.n28 VN.n6 0.189894
R138 VN.n29 VN.n28 0.189894
R139 VN.n30 VN.n29 0.189894
R140 VN.n30 VN.n4 0.189894
R141 VN.n35 VN.n4 0.189894
R142 VN.n36 VN.n35 0.189894
R143 VN.n37 VN.n36 0.189894
R144 VN.n37 VN.n2 0.189894
R145 VN.n41 VN.n2 0.189894
R146 VN.n42 VN.n41 0.189894
R147 VN.n43 VN.n42 0.189894
R148 VN.n43 VN.n0 0.189894
R149 VN VN.n47 0.153454
R150 VDD2.n1 VDD2.t2 84.6912
R151 VDD2.n4 VDD2.t4 81.7775
R152 VDD2.n3 VDD2.n2 80.5319
R153 VDD2 VDD2.n7 80.5292
R154 VDD2.n6 VDD2.n5 78.4022
R155 VDD2.n1 VDD2.n0 78.4019
R156 VDD2.n4 VDD2.n3 45.8575
R157 VDD2.n7 VDD2.t6 3.37589
R158 VDD2.n7 VDD2.t9 3.37589
R159 VDD2.n5 VDD2.t8 3.37589
R160 VDD2.n5 VDD2.t7 3.37589
R161 VDD2.n2 VDD2.t5 3.37589
R162 VDD2.n2 VDD2.t3 3.37589
R163 VDD2.n0 VDD2.t0 3.37589
R164 VDD2.n0 VDD2.t1 3.37589
R165 VDD2.n6 VDD2.n4 2.91429
R166 VDD2 VDD2.n6 0.787138
R167 VDD2.n3 VDD2.n1 0.673602
R168 VTAIL.n11 VTAIL.t6 65.0987
R169 VTAIL.n17 VTAIL.t9 65.0986
R170 VTAIL.n2 VTAIL.t17 65.0986
R171 VTAIL.n16 VTAIL.t1 65.0986
R172 VTAIL.n15 VTAIL.n14 61.7234
R173 VTAIL.n13 VTAIL.n12 61.7234
R174 VTAIL.n10 VTAIL.n9 61.7234
R175 VTAIL.n8 VTAIL.n7 61.7234
R176 VTAIL.n19 VTAIL.n18 61.7232
R177 VTAIL.n1 VTAIL.n0 61.7232
R178 VTAIL.n4 VTAIL.n3 61.7232
R179 VTAIL.n6 VTAIL.n5 61.7232
R180 VTAIL.n8 VTAIL.n6 26.4962
R181 VTAIL.n17 VTAIL.n16 23.5824
R182 VTAIL.n18 VTAIL.t7 3.37589
R183 VTAIL.n18 VTAIL.t8 3.37589
R184 VTAIL.n0 VTAIL.t10 3.37589
R185 VTAIL.n0 VTAIL.t5 3.37589
R186 VTAIL.n3 VTAIL.t15 3.37589
R187 VTAIL.n3 VTAIL.t16 3.37589
R188 VTAIL.n5 VTAIL.t0 3.37589
R189 VTAIL.n5 VTAIL.t18 3.37589
R190 VTAIL.n14 VTAIL.t13 3.37589
R191 VTAIL.n14 VTAIL.t14 3.37589
R192 VTAIL.n12 VTAIL.t2 3.37589
R193 VTAIL.n12 VTAIL.t19 3.37589
R194 VTAIL.n9 VTAIL.t4 3.37589
R195 VTAIL.n9 VTAIL.t12 3.37589
R196 VTAIL.n7 VTAIL.t3 3.37589
R197 VTAIL.n7 VTAIL.t11 3.37589
R198 VTAIL.n10 VTAIL.n8 2.91429
R199 VTAIL.n11 VTAIL.n10 2.91429
R200 VTAIL.n15 VTAIL.n13 2.91429
R201 VTAIL.n16 VTAIL.n15 2.91429
R202 VTAIL.n6 VTAIL.n4 2.91429
R203 VTAIL.n4 VTAIL.n2 2.91429
R204 VTAIL.n19 VTAIL.n17 2.91429
R205 VTAIL VTAIL.n1 2.24403
R206 VTAIL.n13 VTAIL.n11 1.92722
R207 VTAIL.n2 VTAIL.n1 1.92722
R208 VTAIL VTAIL.n19 0.670759
R209 VP.n30 VP.n29 161.3
R210 VP.n31 VP.n26 161.3
R211 VP.n33 VP.n32 161.3
R212 VP.n34 VP.n25 161.3
R213 VP.n36 VP.n35 161.3
R214 VP.n37 VP.n24 161.3
R215 VP.n39 VP.n38 161.3
R216 VP.n41 VP.n40 161.3
R217 VP.n42 VP.n22 161.3
R218 VP.n44 VP.n43 161.3
R219 VP.n45 VP.n21 161.3
R220 VP.n47 VP.n46 161.3
R221 VP.n48 VP.n20 161.3
R222 VP.n51 VP.n50 161.3
R223 VP.n52 VP.n19 161.3
R224 VP.n54 VP.n53 161.3
R225 VP.n55 VP.n18 161.3
R226 VP.n57 VP.n56 161.3
R227 VP.n58 VP.n17 161.3
R228 VP.n60 VP.n59 161.3
R229 VP.n61 VP.n16 161.3
R230 VP.n108 VP.n0 161.3
R231 VP.n107 VP.n106 161.3
R232 VP.n105 VP.n1 161.3
R233 VP.n104 VP.n103 161.3
R234 VP.n102 VP.n2 161.3
R235 VP.n101 VP.n100 161.3
R236 VP.n99 VP.n3 161.3
R237 VP.n98 VP.n97 161.3
R238 VP.n95 VP.n4 161.3
R239 VP.n94 VP.n93 161.3
R240 VP.n92 VP.n5 161.3
R241 VP.n91 VP.n90 161.3
R242 VP.n89 VP.n6 161.3
R243 VP.n88 VP.n87 161.3
R244 VP.n86 VP.n85 161.3
R245 VP.n84 VP.n8 161.3
R246 VP.n83 VP.n82 161.3
R247 VP.n81 VP.n9 161.3
R248 VP.n80 VP.n79 161.3
R249 VP.n78 VP.n10 161.3
R250 VP.n77 VP.n76 161.3
R251 VP.n75 VP.n74 161.3
R252 VP.n73 VP.n12 161.3
R253 VP.n72 VP.n71 161.3
R254 VP.n70 VP.n13 161.3
R255 VP.n69 VP.n68 161.3
R256 VP.n67 VP.n14 161.3
R257 VP.n66 VP.n65 161.3
R258 VP.n64 VP.n15 110.267
R259 VP.n110 VP.n109 110.267
R260 VP.n63 VP.n62 110.267
R261 VP.n28 VP.t0 108.037
R262 VP.n15 VP.t6 76.0933
R263 VP.n11 VP.t3 76.0933
R264 VP.n7 VP.t4 76.0933
R265 VP.n96 VP.t9 76.0933
R266 VP.n109 VP.t5 76.0933
R267 VP.n62 VP.t1 76.0933
R268 VP.n49 VP.t7 76.0933
R269 VP.n23 VP.t2 76.0933
R270 VP.n27 VP.t8 76.0933
R271 VP.n28 VP.n27 67.6363
R272 VP.n72 VP.n13 56.5193
R273 VP.n56 VP.n55 56.5193
R274 VP.n103 VP.n102 56.5193
R275 VP.n64 VP.n63 53.7496
R276 VP.n83 VP.n9 46.321
R277 VP.n90 VP.n5 46.321
R278 VP.n43 VP.n21 46.321
R279 VP.n36 VP.n25 46.321
R280 VP.n79 VP.n9 34.6658
R281 VP.n94 VP.n5 34.6658
R282 VP.n47 VP.n21 34.6658
R283 VP.n32 VP.n25 34.6658
R284 VP.n67 VP.n66 24.4675
R285 VP.n68 VP.n67 24.4675
R286 VP.n68 VP.n13 24.4675
R287 VP.n73 VP.n72 24.4675
R288 VP.n74 VP.n73 24.4675
R289 VP.n78 VP.n77 24.4675
R290 VP.n79 VP.n78 24.4675
R291 VP.n84 VP.n83 24.4675
R292 VP.n85 VP.n84 24.4675
R293 VP.n89 VP.n88 24.4675
R294 VP.n90 VP.n89 24.4675
R295 VP.n95 VP.n94 24.4675
R296 VP.n97 VP.n95 24.4675
R297 VP.n101 VP.n3 24.4675
R298 VP.n102 VP.n101 24.4675
R299 VP.n103 VP.n1 24.4675
R300 VP.n107 VP.n1 24.4675
R301 VP.n108 VP.n107 24.4675
R302 VP.n56 VP.n17 24.4675
R303 VP.n60 VP.n17 24.4675
R304 VP.n61 VP.n60 24.4675
R305 VP.n48 VP.n47 24.4675
R306 VP.n50 VP.n48 24.4675
R307 VP.n54 VP.n19 24.4675
R308 VP.n55 VP.n54 24.4675
R309 VP.n37 VP.n36 24.4675
R310 VP.n38 VP.n37 24.4675
R311 VP.n42 VP.n41 24.4675
R312 VP.n43 VP.n42 24.4675
R313 VP.n31 VP.n30 24.4675
R314 VP.n32 VP.n31 24.4675
R315 VP.n74 VP.n11 18.1061
R316 VP.n96 VP.n3 18.1061
R317 VP.n49 VP.n19 18.1061
R318 VP.n85 VP.n7 12.234
R319 VP.n88 VP.n7 12.234
R320 VP.n38 VP.n23 12.234
R321 VP.n41 VP.n23 12.234
R322 VP.n77 VP.n11 6.36192
R323 VP.n97 VP.n96 6.36192
R324 VP.n50 VP.n49 6.36192
R325 VP.n30 VP.n27 6.36192
R326 VP.n29 VP.n28 5.21216
R327 VP.n66 VP.n15 0.48984
R328 VP.n109 VP.n108 0.48984
R329 VP.n62 VP.n61 0.48984
R330 VP.n63 VP.n16 0.278367
R331 VP.n65 VP.n64 0.278367
R332 VP.n110 VP.n0 0.278367
R333 VP.n29 VP.n26 0.189894
R334 VP.n33 VP.n26 0.189894
R335 VP.n34 VP.n33 0.189894
R336 VP.n35 VP.n34 0.189894
R337 VP.n35 VP.n24 0.189894
R338 VP.n39 VP.n24 0.189894
R339 VP.n40 VP.n39 0.189894
R340 VP.n40 VP.n22 0.189894
R341 VP.n44 VP.n22 0.189894
R342 VP.n45 VP.n44 0.189894
R343 VP.n46 VP.n45 0.189894
R344 VP.n46 VP.n20 0.189894
R345 VP.n51 VP.n20 0.189894
R346 VP.n52 VP.n51 0.189894
R347 VP.n53 VP.n52 0.189894
R348 VP.n53 VP.n18 0.189894
R349 VP.n57 VP.n18 0.189894
R350 VP.n58 VP.n57 0.189894
R351 VP.n59 VP.n58 0.189894
R352 VP.n59 VP.n16 0.189894
R353 VP.n65 VP.n14 0.189894
R354 VP.n69 VP.n14 0.189894
R355 VP.n70 VP.n69 0.189894
R356 VP.n71 VP.n70 0.189894
R357 VP.n71 VP.n12 0.189894
R358 VP.n75 VP.n12 0.189894
R359 VP.n76 VP.n75 0.189894
R360 VP.n76 VP.n10 0.189894
R361 VP.n80 VP.n10 0.189894
R362 VP.n81 VP.n80 0.189894
R363 VP.n82 VP.n81 0.189894
R364 VP.n82 VP.n8 0.189894
R365 VP.n86 VP.n8 0.189894
R366 VP.n87 VP.n86 0.189894
R367 VP.n87 VP.n6 0.189894
R368 VP.n91 VP.n6 0.189894
R369 VP.n92 VP.n91 0.189894
R370 VP.n93 VP.n92 0.189894
R371 VP.n93 VP.n4 0.189894
R372 VP.n98 VP.n4 0.189894
R373 VP.n99 VP.n98 0.189894
R374 VP.n100 VP.n99 0.189894
R375 VP.n100 VP.n2 0.189894
R376 VP.n104 VP.n2 0.189894
R377 VP.n105 VP.n104 0.189894
R378 VP.n106 VP.n105 0.189894
R379 VP.n106 VP.n0 0.189894
R380 VP VP.n110 0.153454
R381 VDD1.n1 VDD1.t9 84.6913
R382 VDD1.n3 VDD1.t3 84.6912
R383 VDD1.n5 VDD1.n4 80.5319
R384 VDD1.n1 VDD1.n0 78.4022
R385 VDD1.n7 VDD1.n6 78.402
R386 VDD1.n3 VDD1.n2 78.4019
R387 VDD1.n7 VDD1.n5 47.8974
R388 VDD1.n6 VDD1.t2 3.37589
R389 VDD1.n6 VDD1.t8 3.37589
R390 VDD1.n0 VDD1.t1 3.37589
R391 VDD1.n0 VDD1.t7 3.37589
R392 VDD1.n4 VDD1.t0 3.37589
R393 VDD1.n4 VDD1.t4 3.37589
R394 VDD1.n2 VDD1.t6 3.37589
R395 VDD1.n2 VDD1.t5 3.37589
R396 VDD1 VDD1.n7 2.12766
R397 VDD1 VDD1.n1 0.787138
R398 VDD1.n5 VDD1.n3 0.673602
R399 B.n442 B.n147 585
R400 B.n441 B.n440 585
R401 B.n439 B.n148 585
R402 B.n438 B.n437 585
R403 B.n436 B.n149 585
R404 B.n435 B.n434 585
R405 B.n433 B.n150 585
R406 B.n432 B.n431 585
R407 B.n430 B.n151 585
R408 B.n429 B.n428 585
R409 B.n427 B.n152 585
R410 B.n426 B.n425 585
R411 B.n424 B.n153 585
R412 B.n423 B.n422 585
R413 B.n421 B.n154 585
R414 B.n420 B.n419 585
R415 B.n418 B.n155 585
R416 B.n417 B.n416 585
R417 B.n415 B.n156 585
R418 B.n414 B.n413 585
R419 B.n412 B.n157 585
R420 B.n411 B.n410 585
R421 B.n409 B.n158 585
R422 B.n408 B.n407 585
R423 B.n406 B.n159 585
R424 B.n405 B.n404 585
R425 B.n403 B.n160 585
R426 B.n402 B.n401 585
R427 B.n400 B.n161 585
R428 B.n399 B.n398 585
R429 B.n397 B.n162 585
R430 B.n396 B.n395 585
R431 B.n394 B.n163 585
R432 B.n393 B.n392 585
R433 B.n391 B.n164 585
R434 B.n390 B.n389 585
R435 B.n385 B.n165 585
R436 B.n384 B.n383 585
R437 B.n382 B.n166 585
R438 B.n381 B.n380 585
R439 B.n379 B.n167 585
R440 B.n378 B.n377 585
R441 B.n376 B.n168 585
R442 B.n375 B.n374 585
R443 B.n372 B.n169 585
R444 B.n371 B.n370 585
R445 B.n369 B.n172 585
R446 B.n368 B.n367 585
R447 B.n366 B.n173 585
R448 B.n365 B.n364 585
R449 B.n363 B.n174 585
R450 B.n362 B.n361 585
R451 B.n360 B.n175 585
R452 B.n359 B.n358 585
R453 B.n357 B.n176 585
R454 B.n356 B.n355 585
R455 B.n354 B.n177 585
R456 B.n353 B.n352 585
R457 B.n351 B.n178 585
R458 B.n350 B.n349 585
R459 B.n348 B.n179 585
R460 B.n347 B.n346 585
R461 B.n345 B.n180 585
R462 B.n344 B.n343 585
R463 B.n342 B.n181 585
R464 B.n341 B.n340 585
R465 B.n339 B.n182 585
R466 B.n338 B.n337 585
R467 B.n336 B.n183 585
R468 B.n335 B.n334 585
R469 B.n333 B.n184 585
R470 B.n332 B.n331 585
R471 B.n330 B.n185 585
R472 B.n329 B.n328 585
R473 B.n327 B.n186 585
R474 B.n326 B.n325 585
R475 B.n324 B.n187 585
R476 B.n323 B.n322 585
R477 B.n321 B.n188 585
R478 B.n444 B.n443 585
R479 B.n445 B.n146 585
R480 B.n447 B.n446 585
R481 B.n448 B.n145 585
R482 B.n450 B.n449 585
R483 B.n451 B.n144 585
R484 B.n453 B.n452 585
R485 B.n454 B.n143 585
R486 B.n456 B.n455 585
R487 B.n457 B.n142 585
R488 B.n459 B.n458 585
R489 B.n460 B.n141 585
R490 B.n462 B.n461 585
R491 B.n463 B.n140 585
R492 B.n465 B.n464 585
R493 B.n466 B.n139 585
R494 B.n468 B.n467 585
R495 B.n469 B.n138 585
R496 B.n471 B.n470 585
R497 B.n472 B.n137 585
R498 B.n474 B.n473 585
R499 B.n475 B.n136 585
R500 B.n477 B.n476 585
R501 B.n478 B.n135 585
R502 B.n480 B.n479 585
R503 B.n481 B.n134 585
R504 B.n483 B.n482 585
R505 B.n484 B.n133 585
R506 B.n486 B.n485 585
R507 B.n487 B.n132 585
R508 B.n489 B.n488 585
R509 B.n490 B.n131 585
R510 B.n492 B.n491 585
R511 B.n493 B.n130 585
R512 B.n495 B.n494 585
R513 B.n496 B.n129 585
R514 B.n498 B.n497 585
R515 B.n499 B.n128 585
R516 B.n501 B.n500 585
R517 B.n502 B.n127 585
R518 B.n504 B.n503 585
R519 B.n505 B.n126 585
R520 B.n507 B.n506 585
R521 B.n508 B.n125 585
R522 B.n510 B.n509 585
R523 B.n511 B.n124 585
R524 B.n513 B.n512 585
R525 B.n514 B.n123 585
R526 B.n516 B.n515 585
R527 B.n517 B.n122 585
R528 B.n519 B.n518 585
R529 B.n520 B.n121 585
R530 B.n522 B.n521 585
R531 B.n523 B.n120 585
R532 B.n525 B.n524 585
R533 B.n526 B.n119 585
R534 B.n528 B.n527 585
R535 B.n529 B.n118 585
R536 B.n531 B.n530 585
R537 B.n532 B.n117 585
R538 B.n534 B.n533 585
R539 B.n535 B.n116 585
R540 B.n537 B.n536 585
R541 B.n538 B.n115 585
R542 B.n540 B.n539 585
R543 B.n541 B.n114 585
R544 B.n543 B.n542 585
R545 B.n544 B.n113 585
R546 B.n546 B.n545 585
R547 B.n547 B.n112 585
R548 B.n549 B.n548 585
R549 B.n550 B.n111 585
R550 B.n552 B.n551 585
R551 B.n553 B.n110 585
R552 B.n555 B.n554 585
R553 B.n556 B.n109 585
R554 B.n558 B.n557 585
R555 B.n559 B.n108 585
R556 B.n561 B.n560 585
R557 B.n562 B.n107 585
R558 B.n564 B.n563 585
R559 B.n565 B.n106 585
R560 B.n567 B.n566 585
R561 B.n568 B.n105 585
R562 B.n570 B.n569 585
R563 B.n571 B.n104 585
R564 B.n573 B.n572 585
R565 B.n574 B.n103 585
R566 B.n576 B.n575 585
R567 B.n577 B.n102 585
R568 B.n579 B.n578 585
R569 B.n580 B.n101 585
R570 B.n582 B.n581 585
R571 B.n583 B.n100 585
R572 B.n585 B.n584 585
R573 B.n586 B.n99 585
R574 B.n588 B.n587 585
R575 B.n589 B.n98 585
R576 B.n591 B.n590 585
R577 B.n592 B.n97 585
R578 B.n594 B.n593 585
R579 B.n595 B.n96 585
R580 B.n597 B.n596 585
R581 B.n598 B.n95 585
R582 B.n600 B.n599 585
R583 B.n601 B.n94 585
R584 B.n603 B.n602 585
R585 B.n604 B.n93 585
R586 B.n606 B.n605 585
R587 B.n607 B.n92 585
R588 B.n609 B.n608 585
R589 B.n610 B.n91 585
R590 B.n612 B.n611 585
R591 B.n613 B.n90 585
R592 B.n615 B.n614 585
R593 B.n616 B.n89 585
R594 B.n618 B.n617 585
R595 B.n619 B.n88 585
R596 B.n621 B.n620 585
R597 B.n622 B.n87 585
R598 B.n624 B.n623 585
R599 B.n625 B.n86 585
R600 B.n627 B.n626 585
R601 B.n628 B.n85 585
R602 B.n630 B.n629 585
R603 B.n631 B.n84 585
R604 B.n633 B.n632 585
R605 B.n634 B.n83 585
R606 B.n636 B.n635 585
R607 B.n637 B.n82 585
R608 B.n639 B.n638 585
R609 B.n640 B.n81 585
R610 B.n642 B.n641 585
R611 B.n643 B.n80 585
R612 B.n645 B.n644 585
R613 B.n646 B.n79 585
R614 B.n767 B.n766 585
R615 B.n765 B.n36 585
R616 B.n764 B.n763 585
R617 B.n762 B.n37 585
R618 B.n761 B.n760 585
R619 B.n759 B.n38 585
R620 B.n758 B.n757 585
R621 B.n756 B.n39 585
R622 B.n755 B.n754 585
R623 B.n753 B.n40 585
R624 B.n752 B.n751 585
R625 B.n750 B.n41 585
R626 B.n749 B.n748 585
R627 B.n747 B.n42 585
R628 B.n746 B.n745 585
R629 B.n744 B.n43 585
R630 B.n743 B.n742 585
R631 B.n741 B.n44 585
R632 B.n740 B.n739 585
R633 B.n738 B.n45 585
R634 B.n737 B.n736 585
R635 B.n735 B.n46 585
R636 B.n734 B.n733 585
R637 B.n732 B.n47 585
R638 B.n731 B.n730 585
R639 B.n729 B.n48 585
R640 B.n728 B.n727 585
R641 B.n726 B.n49 585
R642 B.n725 B.n724 585
R643 B.n723 B.n50 585
R644 B.n722 B.n721 585
R645 B.n720 B.n51 585
R646 B.n719 B.n718 585
R647 B.n717 B.n52 585
R648 B.n716 B.n715 585
R649 B.n713 B.n53 585
R650 B.n712 B.n711 585
R651 B.n710 B.n56 585
R652 B.n709 B.n708 585
R653 B.n707 B.n57 585
R654 B.n706 B.n705 585
R655 B.n704 B.n58 585
R656 B.n703 B.n702 585
R657 B.n701 B.n59 585
R658 B.n699 B.n698 585
R659 B.n697 B.n62 585
R660 B.n696 B.n695 585
R661 B.n694 B.n63 585
R662 B.n693 B.n692 585
R663 B.n691 B.n64 585
R664 B.n690 B.n689 585
R665 B.n688 B.n65 585
R666 B.n687 B.n686 585
R667 B.n685 B.n66 585
R668 B.n684 B.n683 585
R669 B.n682 B.n67 585
R670 B.n681 B.n680 585
R671 B.n679 B.n68 585
R672 B.n678 B.n677 585
R673 B.n676 B.n69 585
R674 B.n675 B.n674 585
R675 B.n673 B.n70 585
R676 B.n672 B.n671 585
R677 B.n670 B.n71 585
R678 B.n669 B.n668 585
R679 B.n667 B.n72 585
R680 B.n666 B.n665 585
R681 B.n664 B.n73 585
R682 B.n663 B.n662 585
R683 B.n661 B.n74 585
R684 B.n660 B.n659 585
R685 B.n658 B.n75 585
R686 B.n657 B.n656 585
R687 B.n655 B.n76 585
R688 B.n654 B.n653 585
R689 B.n652 B.n77 585
R690 B.n651 B.n650 585
R691 B.n649 B.n78 585
R692 B.n648 B.n647 585
R693 B.n768 B.n35 585
R694 B.n770 B.n769 585
R695 B.n771 B.n34 585
R696 B.n773 B.n772 585
R697 B.n774 B.n33 585
R698 B.n776 B.n775 585
R699 B.n777 B.n32 585
R700 B.n779 B.n778 585
R701 B.n780 B.n31 585
R702 B.n782 B.n781 585
R703 B.n783 B.n30 585
R704 B.n785 B.n784 585
R705 B.n786 B.n29 585
R706 B.n788 B.n787 585
R707 B.n789 B.n28 585
R708 B.n791 B.n790 585
R709 B.n792 B.n27 585
R710 B.n794 B.n793 585
R711 B.n795 B.n26 585
R712 B.n797 B.n796 585
R713 B.n798 B.n25 585
R714 B.n800 B.n799 585
R715 B.n801 B.n24 585
R716 B.n803 B.n802 585
R717 B.n804 B.n23 585
R718 B.n806 B.n805 585
R719 B.n807 B.n22 585
R720 B.n809 B.n808 585
R721 B.n810 B.n21 585
R722 B.n812 B.n811 585
R723 B.n813 B.n20 585
R724 B.n815 B.n814 585
R725 B.n816 B.n19 585
R726 B.n818 B.n817 585
R727 B.n819 B.n18 585
R728 B.n821 B.n820 585
R729 B.n822 B.n17 585
R730 B.n824 B.n823 585
R731 B.n825 B.n16 585
R732 B.n827 B.n826 585
R733 B.n828 B.n15 585
R734 B.n830 B.n829 585
R735 B.n831 B.n14 585
R736 B.n833 B.n832 585
R737 B.n834 B.n13 585
R738 B.n836 B.n835 585
R739 B.n837 B.n12 585
R740 B.n839 B.n838 585
R741 B.n840 B.n11 585
R742 B.n842 B.n841 585
R743 B.n843 B.n10 585
R744 B.n845 B.n844 585
R745 B.n846 B.n9 585
R746 B.n848 B.n847 585
R747 B.n849 B.n8 585
R748 B.n851 B.n850 585
R749 B.n852 B.n7 585
R750 B.n854 B.n853 585
R751 B.n855 B.n6 585
R752 B.n857 B.n856 585
R753 B.n858 B.n5 585
R754 B.n860 B.n859 585
R755 B.n861 B.n4 585
R756 B.n863 B.n862 585
R757 B.n864 B.n3 585
R758 B.n866 B.n865 585
R759 B.n867 B.n0 585
R760 B.n2 B.n1 585
R761 B.n222 B.n221 585
R762 B.n224 B.n223 585
R763 B.n225 B.n220 585
R764 B.n227 B.n226 585
R765 B.n228 B.n219 585
R766 B.n230 B.n229 585
R767 B.n231 B.n218 585
R768 B.n233 B.n232 585
R769 B.n234 B.n217 585
R770 B.n236 B.n235 585
R771 B.n237 B.n216 585
R772 B.n239 B.n238 585
R773 B.n240 B.n215 585
R774 B.n242 B.n241 585
R775 B.n243 B.n214 585
R776 B.n245 B.n244 585
R777 B.n246 B.n213 585
R778 B.n248 B.n247 585
R779 B.n249 B.n212 585
R780 B.n251 B.n250 585
R781 B.n252 B.n211 585
R782 B.n254 B.n253 585
R783 B.n255 B.n210 585
R784 B.n257 B.n256 585
R785 B.n258 B.n209 585
R786 B.n260 B.n259 585
R787 B.n261 B.n208 585
R788 B.n263 B.n262 585
R789 B.n264 B.n207 585
R790 B.n266 B.n265 585
R791 B.n267 B.n206 585
R792 B.n269 B.n268 585
R793 B.n270 B.n205 585
R794 B.n272 B.n271 585
R795 B.n273 B.n204 585
R796 B.n275 B.n274 585
R797 B.n276 B.n203 585
R798 B.n278 B.n277 585
R799 B.n279 B.n202 585
R800 B.n281 B.n280 585
R801 B.n282 B.n201 585
R802 B.n284 B.n283 585
R803 B.n285 B.n200 585
R804 B.n287 B.n286 585
R805 B.n288 B.n199 585
R806 B.n290 B.n289 585
R807 B.n291 B.n198 585
R808 B.n293 B.n292 585
R809 B.n294 B.n197 585
R810 B.n296 B.n295 585
R811 B.n297 B.n196 585
R812 B.n299 B.n298 585
R813 B.n300 B.n195 585
R814 B.n302 B.n301 585
R815 B.n303 B.n194 585
R816 B.n305 B.n304 585
R817 B.n306 B.n193 585
R818 B.n308 B.n307 585
R819 B.n309 B.n192 585
R820 B.n311 B.n310 585
R821 B.n312 B.n191 585
R822 B.n314 B.n313 585
R823 B.n315 B.n190 585
R824 B.n317 B.n316 585
R825 B.n318 B.n189 585
R826 B.n320 B.n319 585
R827 B.n321 B.n320 530.939
R828 B.n444 B.n147 530.939
R829 B.n648 B.n79 530.939
R830 B.n766 B.n35 530.939
R831 B.n170 B.t9 284.731
R832 B.n386 B.t6 284.731
R833 B.n60 B.t3 284.731
R834 B.n54 B.t0 284.731
R835 B.n869 B.n868 256.663
R836 B.n868 B.n867 235.042
R837 B.n868 B.n2 235.042
R838 B.n386 B.t7 175.5
R839 B.n60 B.t5 175.5
R840 B.n170 B.t10 175.488
R841 B.n54 B.t2 175.488
R842 B.n322 B.n321 163.367
R843 B.n322 B.n187 163.367
R844 B.n326 B.n187 163.367
R845 B.n327 B.n326 163.367
R846 B.n328 B.n327 163.367
R847 B.n328 B.n185 163.367
R848 B.n332 B.n185 163.367
R849 B.n333 B.n332 163.367
R850 B.n334 B.n333 163.367
R851 B.n334 B.n183 163.367
R852 B.n338 B.n183 163.367
R853 B.n339 B.n338 163.367
R854 B.n340 B.n339 163.367
R855 B.n340 B.n181 163.367
R856 B.n344 B.n181 163.367
R857 B.n345 B.n344 163.367
R858 B.n346 B.n345 163.367
R859 B.n346 B.n179 163.367
R860 B.n350 B.n179 163.367
R861 B.n351 B.n350 163.367
R862 B.n352 B.n351 163.367
R863 B.n352 B.n177 163.367
R864 B.n356 B.n177 163.367
R865 B.n357 B.n356 163.367
R866 B.n358 B.n357 163.367
R867 B.n358 B.n175 163.367
R868 B.n362 B.n175 163.367
R869 B.n363 B.n362 163.367
R870 B.n364 B.n363 163.367
R871 B.n364 B.n173 163.367
R872 B.n368 B.n173 163.367
R873 B.n369 B.n368 163.367
R874 B.n370 B.n369 163.367
R875 B.n370 B.n169 163.367
R876 B.n375 B.n169 163.367
R877 B.n376 B.n375 163.367
R878 B.n377 B.n376 163.367
R879 B.n377 B.n167 163.367
R880 B.n381 B.n167 163.367
R881 B.n382 B.n381 163.367
R882 B.n383 B.n382 163.367
R883 B.n383 B.n165 163.367
R884 B.n390 B.n165 163.367
R885 B.n391 B.n390 163.367
R886 B.n392 B.n391 163.367
R887 B.n392 B.n163 163.367
R888 B.n396 B.n163 163.367
R889 B.n397 B.n396 163.367
R890 B.n398 B.n397 163.367
R891 B.n398 B.n161 163.367
R892 B.n402 B.n161 163.367
R893 B.n403 B.n402 163.367
R894 B.n404 B.n403 163.367
R895 B.n404 B.n159 163.367
R896 B.n408 B.n159 163.367
R897 B.n409 B.n408 163.367
R898 B.n410 B.n409 163.367
R899 B.n410 B.n157 163.367
R900 B.n414 B.n157 163.367
R901 B.n415 B.n414 163.367
R902 B.n416 B.n415 163.367
R903 B.n416 B.n155 163.367
R904 B.n420 B.n155 163.367
R905 B.n421 B.n420 163.367
R906 B.n422 B.n421 163.367
R907 B.n422 B.n153 163.367
R908 B.n426 B.n153 163.367
R909 B.n427 B.n426 163.367
R910 B.n428 B.n427 163.367
R911 B.n428 B.n151 163.367
R912 B.n432 B.n151 163.367
R913 B.n433 B.n432 163.367
R914 B.n434 B.n433 163.367
R915 B.n434 B.n149 163.367
R916 B.n438 B.n149 163.367
R917 B.n439 B.n438 163.367
R918 B.n440 B.n439 163.367
R919 B.n440 B.n147 163.367
R920 B.n644 B.n79 163.367
R921 B.n644 B.n643 163.367
R922 B.n643 B.n642 163.367
R923 B.n642 B.n81 163.367
R924 B.n638 B.n81 163.367
R925 B.n638 B.n637 163.367
R926 B.n637 B.n636 163.367
R927 B.n636 B.n83 163.367
R928 B.n632 B.n83 163.367
R929 B.n632 B.n631 163.367
R930 B.n631 B.n630 163.367
R931 B.n630 B.n85 163.367
R932 B.n626 B.n85 163.367
R933 B.n626 B.n625 163.367
R934 B.n625 B.n624 163.367
R935 B.n624 B.n87 163.367
R936 B.n620 B.n87 163.367
R937 B.n620 B.n619 163.367
R938 B.n619 B.n618 163.367
R939 B.n618 B.n89 163.367
R940 B.n614 B.n89 163.367
R941 B.n614 B.n613 163.367
R942 B.n613 B.n612 163.367
R943 B.n612 B.n91 163.367
R944 B.n608 B.n91 163.367
R945 B.n608 B.n607 163.367
R946 B.n607 B.n606 163.367
R947 B.n606 B.n93 163.367
R948 B.n602 B.n93 163.367
R949 B.n602 B.n601 163.367
R950 B.n601 B.n600 163.367
R951 B.n600 B.n95 163.367
R952 B.n596 B.n95 163.367
R953 B.n596 B.n595 163.367
R954 B.n595 B.n594 163.367
R955 B.n594 B.n97 163.367
R956 B.n590 B.n97 163.367
R957 B.n590 B.n589 163.367
R958 B.n589 B.n588 163.367
R959 B.n588 B.n99 163.367
R960 B.n584 B.n99 163.367
R961 B.n584 B.n583 163.367
R962 B.n583 B.n582 163.367
R963 B.n582 B.n101 163.367
R964 B.n578 B.n101 163.367
R965 B.n578 B.n577 163.367
R966 B.n577 B.n576 163.367
R967 B.n576 B.n103 163.367
R968 B.n572 B.n103 163.367
R969 B.n572 B.n571 163.367
R970 B.n571 B.n570 163.367
R971 B.n570 B.n105 163.367
R972 B.n566 B.n105 163.367
R973 B.n566 B.n565 163.367
R974 B.n565 B.n564 163.367
R975 B.n564 B.n107 163.367
R976 B.n560 B.n107 163.367
R977 B.n560 B.n559 163.367
R978 B.n559 B.n558 163.367
R979 B.n558 B.n109 163.367
R980 B.n554 B.n109 163.367
R981 B.n554 B.n553 163.367
R982 B.n553 B.n552 163.367
R983 B.n552 B.n111 163.367
R984 B.n548 B.n111 163.367
R985 B.n548 B.n547 163.367
R986 B.n547 B.n546 163.367
R987 B.n546 B.n113 163.367
R988 B.n542 B.n113 163.367
R989 B.n542 B.n541 163.367
R990 B.n541 B.n540 163.367
R991 B.n540 B.n115 163.367
R992 B.n536 B.n115 163.367
R993 B.n536 B.n535 163.367
R994 B.n535 B.n534 163.367
R995 B.n534 B.n117 163.367
R996 B.n530 B.n117 163.367
R997 B.n530 B.n529 163.367
R998 B.n529 B.n528 163.367
R999 B.n528 B.n119 163.367
R1000 B.n524 B.n119 163.367
R1001 B.n524 B.n523 163.367
R1002 B.n523 B.n522 163.367
R1003 B.n522 B.n121 163.367
R1004 B.n518 B.n121 163.367
R1005 B.n518 B.n517 163.367
R1006 B.n517 B.n516 163.367
R1007 B.n516 B.n123 163.367
R1008 B.n512 B.n123 163.367
R1009 B.n512 B.n511 163.367
R1010 B.n511 B.n510 163.367
R1011 B.n510 B.n125 163.367
R1012 B.n506 B.n125 163.367
R1013 B.n506 B.n505 163.367
R1014 B.n505 B.n504 163.367
R1015 B.n504 B.n127 163.367
R1016 B.n500 B.n127 163.367
R1017 B.n500 B.n499 163.367
R1018 B.n499 B.n498 163.367
R1019 B.n498 B.n129 163.367
R1020 B.n494 B.n129 163.367
R1021 B.n494 B.n493 163.367
R1022 B.n493 B.n492 163.367
R1023 B.n492 B.n131 163.367
R1024 B.n488 B.n131 163.367
R1025 B.n488 B.n487 163.367
R1026 B.n487 B.n486 163.367
R1027 B.n486 B.n133 163.367
R1028 B.n482 B.n133 163.367
R1029 B.n482 B.n481 163.367
R1030 B.n481 B.n480 163.367
R1031 B.n480 B.n135 163.367
R1032 B.n476 B.n135 163.367
R1033 B.n476 B.n475 163.367
R1034 B.n475 B.n474 163.367
R1035 B.n474 B.n137 163.367
R1036 B.n470 B.n137 163.367
R1037 B.n470 B.n469 163.367
R1038 B.n469 B.n468 163.367
R1039 B.n468 B.n139 163.367
R1040 B.n464 B.n139 163.367
R1041 B.n464 B.n463 163.367
R1042 B.n463 B.n462 163.367
R1043 B.n462 B.n141 163.367
R1044 B.n458 B.n141 163.367
R1045 B.n458 B.n457 163.367
R1046 B.n457 B.n456 163.367
R1047 B.n456 B.n143 163.367
R1048 B.n452 B.n143 163.367
R1049 B.n452 B.n451 163.367
R1050 B.n451 B.n450 163.367
R1051 B.n450 B.n145 163.367
R1052 B.n446 B.n145 163.367
R1053 B.n446 B.n445 163.367
R1054 B.n445 B.n444 163.367
R1055 B.n766 B.n765 163.367
R1056 B.n765 B.n764 163.367
R1057 B.n764 B.n37 163.367
R1058 B.n760 B.n37 163.367
R1059 B.n760 B.n759 163.367
R1060 B.n759 B.n758 163.367
R1061 B.n758 B.n39 163.367
R1062 B.n754 B.n39 163.367
R1063 B.n754 B.n753 163.367
R1064 B.n753 B.n752 163.367
R1065 B.n752 B.n41 163.367
R1066 B.n748 B.n41 163.367
R1067 B.n748 B.n747 163.367
R1068 B.n747 B.n746 163.367
R1069 B.n746 B.n43 163.367
R1070 B.n742 B.n43 163.367
R1071 B.n742 B.n741 163.367
R1072 B.n741 B.n740 163.367
R1073 B.n740 B.n45 163.367
R1074 B.n736 B.n45 163.367
R1075 B.n736 B.n735 163.367
R1076 B.n735 B.n734 163.367
R1077 B.n734 B.n47 163.367
R1078 B.n730 B.n47 163.367
R1079 B.n730 B.n729 163.367
R1080 B.n729 B.n728 163.367
R1081 B.n728 B.n49 163.367
R1082 B.n724 B.n49 163.367
R1083 B.n724 B.n723 163.367
R1084 B.n723 B.n722 163.367
R1085 B.n722 B.n51 163.367
R1086 B.n718 B.n51 163.367
R1087 B.n718 B.n717 163.367
R1088 B.n717 B.n716 163.367
R1089 B.n716 B.n53 163.367
R1090 B.n711 B.n53 163.367
R1091 B.n711 B.n710 163.367
R1092 B.n710 B.n709 163.367
R1093 B.n709 B.n57 163.367
R1094 B.n705 B.n57 163.367
R1095 B.n705 B.n704 163.367
R1096 B.n704 B.n703 163.367
R1097 B.n703 B.n59 163.367
R1098 B.n698 B.n59 163.367
R1099 B.n698 B.n697 163.367
R1100 B.n697 B.n696 163.367
R1101 B.n696 B.n63 163.367
R1102 B.n692 B.n63 163.367
R1103 B.n692 B.n691 163.367
R1104 B.n691 B.n690 163.367
R1105 B.n690 B.n65 163.367
R1106 B.n686 B.n65 163.367
R1107 B.n686 B.n685 163.367
R1108 B.n685 B.n684 163.367
R1109 B.n684 B.n67 163.367
R1110 B.n680 B.n67 163.367
R1111 B.n680 B.n679 163.367
R1112 B.n679 B.n678 163.367
R1113 B.n678 B.n69 163.367
R1114 B.n674 B.n69 163.367
R1115 B.n674 B.n673 163.367
R1116 B.n673 B.n672 163.367
R1117 B.n672 B.n71 163.367
R1118 B.n668 B.n71 163.367
R1119 B.n668 B.n667 163.367
R1120 B.n667 B.n666 163.367
R1121 B.n666 B.n73 163.367
R1122 B.n662 B.n73 163.367
R1123 B.n662 B.n661 163.367
R1124 B.n661 B.n660 163.367
R1125 B.n660 B.n75 163.367
R1126 B.n656 B.n75 163.367
R1127 B.n656 B.n655 163.367
R1128 B.n655 B.n654 163.367
R1129 B.n654 B.n77 163.367
R1130 B.n650 B.n77 163.367
R1131 B.n650 B.n649 163.367
R1132 B.n649 B.n648 163.367
R1133 B.n770 B.n35 163.367
R1134 B.n771 B.n770 163.367
R1135 B.n772 B.n771 163.367
R1136 B.n772 B.n33 163.367
R1137 B.n776 B.n33 163.367
R1138 B.n777 B.n776 163.367
R1139 B.n778 B.n777 163.367
R1140 B.n778 B.n31 163.367
R1141 B.n782 B.n31 163.367
R1142 B.n783 B.n782 163.367
R1143 B.n784 B.n783 163.367
R1144 B.n784 B.n29 163.367
R1145 B.n788 B.n29 163.367
R1146 B.n789 B.n788 163.367
R1147 B.n790 B.n789 163.367
R1148 B.n790 B.n27 163.367
R1149 B.n794 B.n27 163.367
R1150 B.n795 B.n794 163.367
R1151 B.n796 B.n795 163.367
R1152 B.n796 B.n25 163.367
R1153 B.n800 B.n25 163.367
R1154 B.n801 B.n800 163.367
R1155 B.n802 B.n801 163.367
R1156 B.n802 B.n23 163.367
R1157 B.n806 B.n23 163.367
R1158 B.n807 B.n806 163.367
R1159 B.n808 B.n807 163.367
R1160 B.n808 B.n21 163.367
R1161 B.n812 B.n21 163.367
R1162 B.n813 B.n812 163.367
R1163 B.n814 B.n813 163.367
R1164 B.n814 B.n19 163.367
R1165 B.n818 B.n19 163.367
R1166 B.n819 B.n818 163.367
R1167 B.n820 B.n819 163.367
R1168 B.n820 B.n17 163.367
R1169 B.n824 B.n17 163.367
R1170 B.n825 B.n824 163.367
R1171 B.n826 B.n825 163.367
R1172 B.n826 B.n15 163.367
R1173 B.n830 B.n15 163.367
R1174 B.n831 B.n830 163.367
R1175 B.n832 B.n831 163.367
R1176 B.n832 B.n13 163.367
R1177 B.n836 B.n13 163.367
R1178 B.n837 B.n836 163.367
R1179 B.n838 B.n837 163.367
R1180 B.n838 B.n11 163.367
R1181 B.n842 B.n11 163.367
R1182 B.n843 B.n842 163.367
R1183 B.n844 B.n843 163.367
R1184 B.n844 B.n9 163.367
R1185 B.n848 B.n9 163.367
R1186 B.n849 B.n848 163.367
R1187 B.n850 B.n849 163.367
R1188 B.n850 B.n7 163.367
R1189 B.n854 B.n7 163.367
R1190 B.n855 B.n854 163.367
R1191 B.n856 B.n855 163.367
R1192 B.n856 B.n5 163.367
R1193 B.n860 B.n5 163.367
R1194 B.n861 B.n860 163.367
R1195 B.n862 B.n861 163.367
R1196 B.n862 B.n3 163.367
R1197 B.n866 B.n3 163.367
R1198 B.n867 B.n866 163.367
R1199 B.n221 B.n2 163.367
R1200 B.n224 B.n221 163.367
R1201 B.n225 B.n224 163.367
R1202 B.n226 B.n225 163.367
R1203 B.n226 B.n219 163.367
R1204 B.n230 B.n219 163.367
R1205 B.n231 B.n230 163.367
R1206 B.n232 B.n231 163.367
R1207 B.n232 B.n217 163.367
R1208 B.n236 B.n217 163.367
R1209 B.n237 B.n236 163.367
R1210 B.n238 B.n237 163.367
R1211 B.n238 B.n215 163.367
R1212 B.n242 B.n215 163.367
R1213 B.n243 B.n242 163.367
R1214 B.n244 B.n243 163.367
R1215 B.n244 B.n213 163.367
R1216 B.n248 B.n213 163.367
R1217 B.n249 B.n248 163.367
R1218 B.n250 B.n249 163.367
R1219 B.n250 B.n211 163.367
R1220 B.n254 B.n211 163.367
R1221 B.n255 B.n254 163.367
R1222 B.n256 B.n255 163.367
R1223 B.n256 B.n209 163.367
R1224 B.n260 B.n209 163.367
R1225 B.n261 B.n260 163.367
R1226 B.n262 B.n261 163.367
R1227 B.n262 B.n207 163.367
R1228 B.n266 B.n207 163.367
R1229 B.n267 B.n266 163.367
R1230 B.n268 B.n267 163.367
R1231 B.n268 B.n205 163.367
R1232 B.n272 B.n205 163.367
R1233 B.n273 B.n272 163.367
R1234 B.n274 B.n273 163.367
R1235 B.n274 B.n203 163.367
R1236 B.n278 B.n203 163.367
R1237 B.n279 B.n278 163.367
R1238 B.n280 B.n279 163.367
R1239 B.n280 B.n201 163.367
R1240 B.n284 B.n201 163.367
R1241 B.n285 B.n284 163.367
R1242 B.n286 B.n285 163.367
R1243 B.n286 B.n199 163.367
R1244 B.n290 B.n199 163.367
R1245 B.n291 B.n290 163.367
R1246 B.n292 B.n291 163.367
R1247 B.n292 B.n197 163.367
R1248 B.n296 B.n197 163.367
R1249 B.n297 B.n296 163.367
R1250 B.n298 B.n297 163.367
R1251 B.n298 B.n195 163.367
R1252 B.n302 B.n195 163.367
R1253 B.n303 B.n302 163.367
R1254 B.n304 B.n303 163.367
R1255 B.n304 B.n193 163.367
R1256 B.n308 B.n193 163.367
R1257 B.n309 B.n308 163.367
R1258 B.n310 B.n309 163.367
R1259 B.n310 B.n191 163.367
R1260 B.n314 B.n191 163.367
R1261 B.n315 B.n314 163.367
R1262 B.n316 B.n315 163.367
R1263 B.n316 B.n189 163.367
R1264 B.n320 B.n189 163.367
R1265 B.n387 B.t8 109.948
R1266 B.n61 B.t4 109.948
R1267 B.n171 B.t11 109.938
R1268 B.n55 B.t1 109.938
R1269 B.n171 B.n170 65.552
R1270 B.n387 B.n386 65.552
R1271 B.n61 B.n60 65.552
R1272 B.n55 B.n54 65.552
R1273 B.n373 B.n171 59.5399
R1274 B.n388 B.n387 59.5399
R1275 B.n700 B.n61 59.5399
R1276 B.n714 B.n55 59.5399
R1277 B.n768 B.n767 34.4981
R1278 B.n647 B.n646 34.4981
R1279 B.n443 B.n442 34.4981
R1280 B.n319 B.n188 34.4981
R1281 B B.n869 18.0485
R1282 B.n769 B.n768 10.6151
R1283 B.n769 B.n34 10.6151
R1284 B.n773 B.n34 10.6151
R1285 B.n774 B.n773 10.6151
R1286 B.n775 B.n774 10.6151
R1287 B.n775 B.n32 10.6151
R1288 B.n779 B.n32 10.6151
R1289 B.n780 B.n779 10.6151
R1290 B.n781 B.n780 10.6151
R1291 B.n781 B.n30 10.6151
R1292 B.n785 B.n30 10.6151
R1293 B.n786 B.n785 10.6151
R1294 B.n787 B.n786 10.6151
R1295 B.n787 B.n28 10.6151
R1296 B.n791 B.n28 10.6151
R1297 B.n792 B.n791 10.6151
R1298 B.n793 B.n792 10.6151
R1299 B.n793 B.n26 10.6151
R1300 B.n797 B.n26 10.6151
R1301 B.n798 B.n797 10.6151
R1302 B.n799 B.n798 10.6151
R1303 B.n799 B.n24 10.6151
R1304 B.n803 B.n24 10.6151
R1305 B.n804 B.n803 10.6151
R1306 B.n805 B.n804 10.6151
R1307 B.n805 B.n22 10.6151
R1308 B.n809 B.n22 10.6151
R1309 B.n810 B.n809 10.6151
R1310 B.n811 B.n810 10.6151
R1311 B.n811 B.n20 10.6151
R1312 B.n815 B.n20 10.6151
R1313 B.n816 B.n815 10.6151
R1314 B.n817 B.n816 10.6151
R1315 B.n817 B.n18 10.6151
R1316 B.n821 B.n18 10.6151
R1317 B.n822 B.n821 10.6151
R1318 B.n823 B.n822 10.6151
R1319 B.n823 B.n16 10.6151
R1320 B.n827 B.n16 10.6151
R1321 B.n828 B.n827 10.6151
R1322 B.n829 B.n828 10.6151
R1323 B.n829 B.n14 10.6151
R1324 B.n833 B.n14 10.6151
R1325 B.n834 B.n833 10.6151
R1326 B.n835 B.n834 10.6151
R1327 B.n835 B.n12 10.6151
R1328 B.n839 B.n12 10.6151
R1329 B.n840 B.n839 10.6151
R1330 B.n841 B.n840 10.6151
R1331 B.n841 B.n10 10.6151
R1332 B.n845 B.n10 10.6151
R1333 B.n846 B.n845 10.6151
R1334 B.n847 B.n846 10.6151
R1335 B.n847 B.n8 10.6151
R1336 B.n851 B.n8 10.6151
R1337 B.n852 B.n851 10.6151
R1338 B.n853 B.n852 10.6151
R1339 B.n853 B.n6 10.6151
R1340 B.n857 B.n6 10.6151
R1341 B.n858 B.n857 10.6151
R1342 B.n859 B.n858 10.6151
R1343 B.n859 B.n4 10.6151
R1344 B.n863 B.n4 10.6151
R1345 B.n864 B.n863 10.6151
R1346 B.n865 B.n864 10.6151
R1347 B.n865 B.n0 10.6151
R1348 B.n767 B.n36 10.6151
R1349 B.n763 B.n36 10.6151
R1350 B.n763 B.n762 10.6151
R1351 B.n762 B.n761 10.6151
R1352 B.n761 B.n38 10.6151
R1353 B.n757 B.n38 10.6151
R1354 B.n757 B.n756 10.6151
R1355 B.n756 B.n755 10.6151
R1356 B.n755 B.n40 10.6151
R1357 B.n751 B.n40 10.6151
R1358 B.n751 B.n750 10.6151
R1359 B.n750 B.n749 10.6151
R1360 B.n749 B.n42 10.6151
R1361 B.n745 B.n42 10.6151
R1362 B.n745 B.n744 10.6151
R1363 B.n744 B.n743 10.6151
R1364 B.n743 B.n44 10.6151
R1365 B.n739 B.n44 10.6151
R1366 B.n739 B.n738 10.6151
R1367 B.n738 B.n737 10.6151
R1368 B.n737 B.n46 10.6151
R1369 B.n733 B.n46 10.6151
R1370 B.n733 B.n732 10.6151
R1371 B.n732 B.n731 10.6151
R1372 B.n731 B.n48 10.6151
R1373 B.n727 B.n48 10.6151
R1374 B.n727 B.n726 10.6151
R1375 B.n726 B.n725 10.6151
R1376 B.n725 B.n50 10.6151
R1377 B.n721 B.n50 10.6151
R1378 B.n721 B.n720 10.6151
R1379 B.n720 B.n719 10.6151
R1380 B.n719 B.n52 10.6151
R1381 B.n715 B.n52 10.6151
R1382 B.n713 B.n712 10.6151
R1383 B.n712 B.n56 10.6151
R1384 B.n708 B.n56 10.6151
R1385 B.n708 B.n707 10.6151
R1386 B.n707 B.n706 10.6151
R1387 B.n706 B.n58 10.6151
R1388 B.n702 B.n58 10.6151
R1389 B.n702 B.n701 10.6151
R1390 B.n699 B.n62 10.6151
R1391 B.n695 B.n62 10.6151
R1392 B.n695 B.n694 10.6151
R1393 B.n694 B.n693 10.6151
R1394 B.n693 B.n64 10.6151
R1395 B.n689 B.n64 10.6151
R1396 B.n689 B.n688 10.6151
R1397 B.n688 B.n687 10.6151
R1398 B.n687 B.n66 10.6151
R1399 B.n683 B.n66 10.6151
R1400 B.n683 B.n682 10.6151
R1401 B.n682 B.n681 10.6151
R1402 B.n681 B.n68 10.6151
R1403 B.n677 B.n68 10.6151
R1404 B.n677 B.n676 10.6151
R1405 B.n676 B.n675 10.6151
R1406 B.n675 B.n70 10.6151
R1407 B.n671 B.n70 10.6151
R1408 B.n671 B.n670 10.6151
R1409 B.n670 B.n669 10.6151
R1410 B.n669 B.n72 10.6151
R1411 B.n665 B.n72 10.6151
R1412 B.n665 B.n664 10.6151
R1413 B.n664 B.n663 10.6151
R1414 B.n663 B.n74 10.6151
R1415 B.n659 B.n74 10.6151
R1416 B.n659 B.n658 10.6151
R1417 B.n658 B.n657 10.6151
R1418 B.n657 B.n76 10.6151
R1419 B.n653 B.n76 10.6151
R1420 B.n653 B.n652 10.6151
R1421 B.n652 B.n651 10.6151
R1422 B.n651 B.n78 10.6151
R1423 B.n647 B.n78 10.6151
R1424 B.n646 B.n645 10.6151
R1425 B.n645 B.n80 10.6151
R1426 B.n641 B.n80 10.6151
R1427 B.n641 B.n640 10.6151
R1428 B.n640 B.n639 10.6151
R1429 B.n639 B.n82 10.6151
R1430 B.n635 B.n82 10.6151
R1431 B.n635 B.n634 10.6151
R1432 B.n634 B.n633 10.6151
R1433 B.n633 B.n84 10.6151
R1434 B.n629 B.n84 10.6151
R1435 B.n629 B.n628 10.6151
R1436 B.n628 B.n627 10.6151
R1437 B.n627 B.n86 10.6151
R1438 B.n623 B.n86 10.6151
R1439 B.n623 B.n622 10.6151
R1440 B.n622 B.n621 10.6151
R1441 B.n621 B.n88 10.6151
R1442 B.n617 B.n88 10.6151
R1443 B.n617 B.n616 10.6151
R1444 B.n616 B.n615 10.6151
R1445 B.n615 B.n90 10.6151
R1446 B.n611 B.n90 10.6151
R1447 B.n611 B.n610 10.6151
R1448 B.n610 B.n609 10.6151
R1449 B.n609 B.n92 10.6151
R1450 B.n605 B.n92 10.6151
R1451 B.n605 B.n604 10.6151
R1452 B.n604 B.n603 10.6151
R1453 B.n603 B.n94 10.6151
R1454 B.n599 B.n94 10.6151
R1455 B.n599 B.n598 10.6151
R1456 B.n598 B.n597 10.6151
R1457 B.n597 B.n96 10.6151
R1458 B.n593 B.n96 10.6151
R1459 B.n593 B.n592 10.6151
R1460 B.n592 B.n591 10.6151
R1461 B.n591 B.n98 10.6151
R1462 B.n587 B.n98 10.6151
R1463 B.n587 B.n586 10.6151
R1464 B.n586 B.n585 10.6151
R1465 B.n585 B.n100 10.6151
R1466 B.n581 B.n100 10.6151
R1467 B.n581 B.n580 10.6151
R1468 B.n580 B.n579 10.6151
R1469 B.n579 B.n102 10.6151
R1470 B.n575 B.n102 10.6151
R1471 B.n575 B.n574 10.6151
R1472 B.n574 B.n573 10.6151
R1473 B.n573 B.n104 10.6151
R1474 B.n569 B.n104 10.6151
R1475 B.n569 B.n568 10.6151
R1476 B.n568 B.n567 10.6151
R1477 B.n567 B.n106 10.6151
R1478 B.n563 B.n106 10.6151
R1479 B.n563 B.n562 10.6151
R1480 B.n562 B.n561 10.6151
R1481 B.n561 B.n108 10.6151
R1482 B.n557 B.n108 10.6151
R1483 B.n557 B.n556 10.6151
R1484 B.n556 B.n555 10.6151
R1485 B.n555 B.n110 10.6151
R1486 B.n551 B.n110 10.6151
R1487 B.n551 B.n550 10.6151
R1488 B.n550 B.n549 10.6151
R1489 B.n549 B.n112 10.6151
R1490 B.n545 B.n112 10.6151
R1491 B.n545 B.n544 10.6151
R1492 B.n544 B.n543 10.6151
R1493 B.n543 B.n114 10.6151
R1494 B.n539 B.n114 10.6151
R1495 B.n539 B.n538 10.6151
R1496 B.n538 B.n537 10.6151
R1497 B.n537 B.n116 10.6151
R1498 B.n533 B.n116 10.6151
R1499 B.n533 B.n532 10.6151
R1500 B.n532 B.n531 10.6151
R1501 B.n531 B.n118 10.6151
R1502 B.n527 B.n118 10.6151
R1503 B.n527 B.n526 10.6151
R1504 B.n526 B.n525 10.6151
R1505 B.n525 B.n120 10.6151
R1506 B.n521 B.n120 10.6151
R1507 B.n521 B.n520 10.6151
R1508 B.n520 B.n519 10.6151
R1509 B.n519 B.n122 10.6151
R1510 B.n515 B.n122 10.6151
R1511 B.n515 B.n514 10.6151
R1512 B.n514 B.n513 10.6151
R1513 B.n513 B.n124 10.6151
R1514 B.n509 B.n124 10.6151
R1515 B.n509 B.n508 10.6151
R1516 B.n508 B.n507 10.6151
R1517 B.n507 B.n126 10.6151
R1518 B.n503 B.n126 10.6151
R1519 B.n503 B.n502 10.6151
R1520 B.n502 B.n501 10.6151
R1521 B.n501 B.n128 10.6151
R1522 B.n497 B.n128 10.6151
R1523 B.n497 B.n496 10.6151
R1524 B.n496 B.n495 10.6151
R1525 B.n495 B.n130 10.6151
R1526 B.n491 B.n130 10.6151
R1527 B.n491 B.n490 10.6151
R1528 B.n490 B.n489 10.6151
R1529 B.n489 B.n132 10.6151
R1530 B.n485 B.n132 10.6151
R1531 B.n485 B.n484 10.6151
R1532 B.n484 B.n483 10.6151
R1533 B.n483 B.n134 10.6151
R1534 B.n479 B.n134 10.6151
R1535 B.n479 B.n478 10.6151
R1536 B.n478 B.n477 10.6151
R1537 B.n477 B.n136 10.6151
R1538 B.n473 B.n136 10.6151
R1539 B.n473 B.n472 10.6151
R1540 B.n472 B.n471 10.6151
R1541 B.n471 B.n138 10.6151
R1542 B.n467 B.n138 10.6151
R1543 B.n467 B.n466 10.6151
R1544 B.n466 B.n465 10.6151
R1545 B.n465 B.n140 10.6151
R1546 B.n461 B.n140 10.6151
R1547 B.n461 B.n460 10.6151
R1548 B.n460 B.n459 10.6151
R1549 B.n459 B.n142 10.6151
R1550 B.n455 B.n142 10.6151
R1551 B.n455 B.n454 10.6151
R1552 B.n454 B.n453 10.6151
R1553 B.n453 B.n144 10.6151
R1554 B.n449 B.n144 10.6151
R1555 B.n449 B.n448 10.6151
R1556 B.n448 B.n447 10.6151
R1557 B.n447 B.n146 10.6151
R1558 B.n443 B.n146 10.6151
R1559 B.n222 B.n1 10.6151
R1560 B.n223 B.n222 10.6151
R1561 B.n223 B.n220 10.6151
R1562 B.n227 B.n220 10.6151
R1563 B.n228 B.n227 10.6151
R1564 B.n229 B.n228 10.6151
R1565 B.n229 B.n218 10.6151
R1566 B.n233 B.n218 10.6151
R1567 B.n234 B.n233 10.6151
R1568 B.n235 B.n234 10.6151
R1569 B.n235 B.n216 10.6151
R1570 B.n239 B.n216 10.6151
R1571 B.n240 B.n239 10.6151
R1572 B.n241 B.n240 10.6151
R1573 B.n241 B.n214 10.6151
R1574 B.n245 B.n214 10.6151
R1575 B.n246 B.n245 10.6151
R1576 B.n247 B.n246 10.6151
R1577 B.n247 B.n212 10.6151
R1578 B.n251 B.n212 10.6151
R1579 B.n252 B.n251 10.6151
R1580 B.n253 B.n252 10.6151
R1581 B.n253 B.n210 10.6151
R1582 B.n257 B.n210 10.6151
R1583 B.n258 B.n257 10.6151
R1584 B.n259 B.n258 10.6151
R1585 B.n259 B.n208 10.6151
R1586 B.n263 B.n208 10.6151
R1587 B.n264 B.n263 10.6151
R1588 B.n265 B.n264 10.6151
R1589 B.n265 B.n206 10.6151
R1590 B.n269 B.n206 10.6151
R1591 B.n270 B.n269 10.6151
R1592 B.n271 B.n270 10.6151
R1593 B.n271 B.n204 10.6151
R1594 B.n275 B.n204 10.6151
R1595 B.n276 B.n275 10.6151
R1596 B.n277 B.n276 10.6151
R1597 B.n277 B.n202 10.6151
R1598 B.n281 B.n202 10.6151
R1599 B.n282 B.n281 10.6151
R1600 B.n283 B.n282 10.6151
R1601 B.n283 B.n200 10.6151
R1602 B.n287 B.n200 10.6151
R1603 B.n288 B.n287 10.6151
R1604 B.n289 B.n288 10.6151
R1605 B.n289 B.n198 10.6151
R1606 B.n293 B.n198 10.6151
R1607 B.n294 B.n293 10.6151
R1608 B.n295 B.n294 10.6151
R1609 B.n295 B.n196 10.6151
R1610 B.n299 B.n196 10.6151
R1611 B.n300 B.n299 10.6151
R1612 B.n301 B.n300 10.6151
R1613 B.n301 B.n194 10.6151
R1614 B.n305 B.n194 10.6151
R1615 B.n306 B.n305 10.6151
R1616 B.n307 B.n306 10.6151
R1617 B.n307 B.n192 10.6151
R1618 B.n311 B.n192 10.6151
R1619 B.n312 B.n311 10.6151
R1620 B.n313 B.n312 10.6151
R1621 B.n313 B.n190 10.6151
R1622 B.n317 B.n190 10.6151
R1623 B.n318 B.n317 10.6151
R1624 B.n319 B.n318 10.6151
R1625 B.n323 B.n188 10.6151
R1626 B.n324 B.n323 10.6151
R1627 B.n325 B.n324 10.6151
R1628 B.n325 B.n186 10.6151
R1629 B.n329 B.n186 10.6151
R1630 B.n330 B.n329 10.6151
R1631 B.n331 B.n330 10.6151
R1632 B.n331 B.n184 10.6151
R1633 B.n335 B.n184 10.6151
R1634 B.n336 B.n335 10.6151
R1635 B.n337 B.n336 10.6151
R1636 B.n337 B.n182 10.6151
R1637 B.n341 B.n182 10.6151
R1638 B.n342 B.n341 10.6151
R1639 B.n343 B.n342 10.6151
R1640 B.n343 B.n180 10.6151
R1641 B.n347 B.n180 10.6151
R1642 B.n348 B.n347 10.6151
R1643 B.n349 B.n348 10.6151
R1644 B.n349 B.n178 10.6151
R1645 B.n353 B.n178 10.6151
R1646 B.n354 B.n353 10.6151
R1647 B.n355 B.n354 10.6151
R1648 B.n355 B.n176 10.6151
R1649 B.n359 B.n176 10.6151
R1650 B.n360 B.n359 10.6151
R1651 B.n361 B.n360 10.6151
R1652 B.n361 B.n174 10.6151
R1653 B.n365 B.n174 10.6151
R1654 B.n366 B.n365 10.6151
R1655 B.n367 B.n366 10.6151
R1656 B.n367 B.n172 10.6151
R1657 B.n371 B.n172 10.6151
R1658 B.n372 B.n371 10.6151
R1659 B.n374 B.n168 10.6151
R1660 B.n378 B.n168 10.6151
R1661 B.n379 B.n378 10.6151
R1662 B.n380 B.n379 10.6151
R1663 B.n380 B.n166 10.6151
R1664 B.n384 B.n166 10.6151
R1665 B.n385 B.n384 10.6151
R1666 B.n389 B.n385 10.6151
R1667 B.n393 B.n164 10.6151
R1668 B.n394 B.n393 10.6151
R1669 B.n395 B.n394 10.6151
R1670 B.n395 B.n162 10.6151
R1671 B.n399 B.n162 10.6151
R1672 B.n400 B.n399 10.6151
R1673 B.n401 B.n400 10.6151
R1674 B.n401 B.n160 10.6151
R1675 B.n405 B.n160 10.6151
R1676 B.n406 B.n405 10.6151
R1677 B.n407 B.n406 10.6151
R1678 B.n407 B.n158 10.6151
R1679 B.n411 B.n158 10.6151
R1680 B.n412 B.n411 10.6151
R1681 B.n413 B.n412 10.6151
R1682 B.n413 B.n156 10.6151
R1683 B.n417 B.n156 10.6151
R1684 B.n418 B.n417 10.6151
R1685 B.n419 B.n418 10.6151
R1686 B.n419 B.n154 10.6151
R1687 B.n423 B.n154 10.6151
R1688 B.n424 B.n423 10.6151
R1689 B.n425 B.n424 10.6151
R1690 B.n425 B.n152 10.6151
R1691 B.n429 B.n152 10.6151
R1692 B.n430 B.n429 10.6151
R1693 B.n431 B.n430 10.6151
R1694 B.n431 B.n150 10.6151
R1695 B.n435 B.n150 10.6151
R1696 B.n436 B.n435 10.6151
R1697 B.n437 B.n436 10.6151
R1698 B.n437 B.n148 10.6151
R1699 B.n441 B.n148 10.6151
R1700 B.n442 B.n441 10.6151
R1701 B.n869 B.n0 8.11757
R1702 B.n869 B.n1 8.11757
R1703 B.n714 B.n713 6.5566
R1704 B.n701 B.n700 6.5566
R1705 B.n374 B.n373 6.5566
R1706 B.n389 B.n388 6.5566
R1707 B.n715 B.n714 4.05904
R1708 B.n700 B.n699 4.05904
R1709 B.n373 B.n372 4.05904
R1710 B.n388 B.n164 4.05904
C0 VP w_n5026_n2894# 11.4922f
C1 VTAIL VN 9.867599f
C2 VTAIL VDD1 9.53527f
C3 VTAIL B 3.36424f
C4 VN VDD1 0.154361f
C5 VN B 1.36995f
C6 VTAIL w_n5026_n2894# 2.94762f
C7 VN w_n5026_n2894# 10.8365f
C8 VDD1 B 2.46707f
C9 VDD1 w_n5026_n2894# 2.7962f
C10 B w_n5026_n2894# 10.6392f
C11 VP VDD2 0.640793f
C12 VTAIL VDD2 9.59013f
C13 VN VDD2 8.922629f
C14 VTAIL VP 9.88183f
C15 VN VP 8.62108f
C16 VDD1 VDD2 2.46704f
C17 VDD2 B 2.60251f
C18 VDD2 w_n5026_n2894# 2.96314f
C19 VP VDD1 9.40555f
C20 VP B 2.47511f
C21 VDD2 VSUBS 2.3022f
C22 VDD1 VSUBS 2.088703f
C23 VTAIL VSUBS 1.337378f
C24 VN VSUBS 8.368141f
C25 VP VSUBS 4.716497f
C26 B VSUBS 5.72582f
C27 w_n5026_n2894# VSUBS 0.17979p
C28 B.n0 VSUBS 0.008737f
C29 B.n1 VSUBS 0.008737f
C30 B.n2 VSUBS 0.012922f
C31 B.n3 VSUBS 0.009902f
C32 B.n4 VSUBS 0.009902f
C33 B.n5 VSUBS 0.009902f
C34 B.n6 VSUBS 0.009902f
C35 B.n7 VSUBS 0.009902f
C36 B.n8 VSUBS 0.009902f
C37 B.n9 VSUBS 0.009902f
C38 B.n10 VSUBS 0.009902f
C39 B.n11 VSUBS 0.009902f
C40 B.n12 VSUBS 0.009902f
C41 B.n13 VSUBS 0.009902f
C42 B.n14 VSUBS 0.009902f
C43 B.n15 VSUBS 0.009902f
C44 B.n16 VSUBS 0.009902f
C45 B.n17 VSUBS 0.009902f
C46 B.n18 VSUBS 0.009902f
C47 B.n19 VSUBS 0.009902f
C48 B.n20 VSUBS 0.009902f
C49 B.n21 VSUBS 0.009902f
C50 B.n22 VSUBS 0.009902f
C51 B.n23 VSUBS 0.009902f
C52 B.n24 VSUBS 0.009902f
C53 B.n25 VSUBS 0.009902f
C54 B.n26 VSUBS 0.009902f
C55 B.n27 VSUBS 0.009902f
C56 B.n28 VSUBS 0.009902f
C57 B.n29 VSUBS 0.009902f
C58 B.n30 VSUBS 0.009902f
C59 B.n31 VSUBS 0.009902f
C60 B.n32 VSUBS 0.009902f
C61 B.n33 VSUBS 0.009902f
C62 B.n34 VSUBS 0.009902f
C63 B.n35 VSUBS 0.023204f
C64 B.n36 VSUBS 0.009902f
C65 B.n37 VSUBS 0.009902f
C66 B.n38 VSUBS 0.009902f
C67 B.n39 VSUBS 0.009902f
C68 B.n40 VSUBS 0.009902f
C69 B.n41 VSUBS 0.009902f
C70 B.n42 VSUBS 0.009902f
C71 B.n43 VSUBS 0.009902f
C72 B.n44 VSUBS 0.009902f
C73 B.n45 VSUBS 0.009902f
C74 B.n46 VSUBS 0.009902f
C75 B.n47 VSUBS 0.009902f
C76 B.n48 VSUBS 0.009902f
C77 B.n49 VSUBS 0.009902f
C78 B.n50 VSUBS 0.009902f
C79 B.n51 VSUBS 0.009902f
C80 B.n52 VSUBS 0.009902f
C81 B.n53 VSUBS 0.009902f
C82 B.t1 VSUBS 0.432287f
C83 B.t2 VSUBS 0.465825f
C84 B.t0 VSUBS 1.93593f
C85 B.n54 VSUBS 0.254098f
C86 B.n55 VSUBS 0.103908f
C87 B.n56 VSUBS 0.009902f
C88 B.n57 VSUBS 0.009902f
C89 B.n58 VSUBS 0.009902f
C90 B.n59 VSUBS 0.009902f
C91 B.t4 VSUBS 0.432282f
C92 B.t5 VSUBS 0.465819f
C93 B.t3 VSUBS 1.93593f
C94 B.n60 VSUBS 0.254103f
C95 B.n61 VSUBS 0.103913f
C96 B.n62 VSUBS 0.009902f
C97 B.n63 VSUBS 0.009902f
C98 B.n64 VSUBS 0.009902f
C99 B.n65 VSUBS 0.009902f
C100 B.n66 VSUBS 0.009902f
C101 B.n67 VSUBS 0.009902f
C102 B.n68 VSUBS 0.009902f
C103 B.n69 VSUBS 0.009902f
C104 B.n70 VSUBS 0.009902f
C105 B.n71 VSUBS 0.009902f
C106 B.n72 VSUBS 0.009902f
C107 B.n73 VSUBS 0.009902f
C108 B.n74 VSUBS 0.009902f
C109 B.n75 VSUBS 0.009902f
C110 B.n76 VSUBS 0.009902f
C111 B.n77 VSUBS 0.009902f
C112 B.n78 VSUBS 0.009902f
C113 B.n79 VSUBS 0.023204f
C114 B.n80 VSUBS 0.009902f
C115 B.n81 VSUBS 0.009902f
C116 B.n82 VSUBS 0.009902f
C117 B.n83 VSUBS 0.009902f
C118 B.n84 VSUBS 0.009902f
C119 B.n85 VSUBS 0.009902f
C120 B.n86 VSUBS 0.009902f
C121 B.n87 VSUBS 0.009902f
C122 B.n88 VSUBS 0.009902f
C123 B.n89 VSUBS 0.009902f
C124 B.n90 VSUBS 0.009902f
C125 B.n91 VSUBS 0.009902f
C126 B.n92 VSUBS 0.009902f
C127 B.n93 VSUBS 0.009902f
C128 B.n94 VSUBS 0.009902f
C129 B.n95 VSUBS 0.009902f
C130 B.n96 VSUBS 0.009902f
C131 B.n97 VSUBS 0.009902f
C132 B.n98 VSUBS 0.009902f
C133 B.n99 VSUBS 0.009902f
C134 B.n100 VSUBS 0.009902f
C135 B.n101 VSUBS 0.009902f
C136 B.n102 VSUBS 0.009902f
C137 B.n103 VSUBS 0.009902f
C138 B.n104 VSUBS 0.009902f
C139 B.n105 VSUBS 0.009902f
C140 B.n106 VSUBS 0.009902f
C141 B.n107 VSUBS 0.009902f
C142 B.n108 VSUBS 0.009902f
C143 B.n109 VSUBS 0.009902f
C144 B.n110 VSUBS 0.009902f
C145 B.n111 VSUBS 0.009902f
C146 B.n112 VSUBS 0.009902f
C147 B.n113 VSUBS 0.009902f
C148 B.n114 VSUBS 0.009902f
C149 B.n115 VSUBS 0.009902f
C150 B.n116 VSUBS 0.009902f
C151 B.n117 VSUBS 0.009902f
C152 B.n118 VSUBS 0.009902f
C153 B.n119 VSUBS 0.009902f
C154 B.n120 VSUBS 0.009902f
C155 B.n121 VSUBS 0.009902f
C156 B.n122 VSUBS 0.009902f
C157 B.n123 VSUBS 0.009902f
C158 B.n124 VSUBS 0.009902f
C159 B.n125 VSUBS 0.009902f
C160 B.n126 VSUBS 0.009902f
C161 B.n127 VSUBS 0.009902f
C162 B.n128 VSUBS 0.009902f
C163 B.n129 VSUBS 0.009902f
C164 B.n130 VSUBS 0.009902f
C165 B.n131 VSUBS 0.009902f
C166 B.n132 VSUBS 0.009902f
C167 B.n133 VSUBS 0.009902f
C168 B.n134 VSUBS 0.009902f
C169 B.n135 VSUBS 0.009902f
C170 B.n136 VSUBS 0.009902f
C171 B.n137 VSUBS 0.009902f
C172 B.n138 VSUBS 0.009902f
C173 B.n139 VSUBS 0.009902f
C174 B.n140 VSUBS 0.009902f
C175 B.n141 VSUBS 0.009902f
C176 B.n142 VSUBS 0.009902f
C177 B.n143 VSUBS 0.009902f
C178 B.n144 VSUBS 0.009902f
C179 B.n145 VSUBS 0.009902f
C180 B.n146 VSUBS 0.009902f
C181 B.n147 VSUBS 0.024852f
C182 B.n148 VSUBS 0.009902f
C183 B.n149 VSUBS 0.009902f
C184 B.n150 VSUBS 0.009902f
C185 B.n151 VSUBS 0.009902f
C186 B.n152 VSUBS 0.009902f
C187 B.n153 VSUBS 0.009902f
C188 B.n154 VSUBS 0.009902f
C189 B.n155 VSUBS 0.009902f
C190 B.n156 VSUBS 0.009902f
C191 B.n157 VSUBS 0.009902f
C192 B.n158 VSUBS 0.009902f
C193 B.n159 VSUBS 0.009902f
C194 B.n160 VSUBS 0.009902f
C195 B.n161 VSUBS 0.009902f
C196 B.n162 VSUBS 0.009902f
C197 B.n163 VSUBS 0.009902f
C198 B.n164 VSUBS 0.006844f
C199 B.n165 VSUBS 0.009902f
C200 B.n166 VSUBS 0.009902f
C201 B.n167 VSUBS 0.009902f
C202 B.n168 VSUBS 0.009902f
C203 B.n169 VSUBS 0.009902f
C204 B.t11 VSUBS 0.432287f
C205 B.t10 VSUBS 0.465825f
C206 B.t9 VSUBS 1.93593f
C207 B.n170 VSUBS 0.254098f
C208 B.n171 VSUBS 0.103908f
C209 B.n172 VSUBS 0.009902f
C210 B.n173 VSUBS 0.009902f
C211 B.n174 VSUBS 0.009902f
C212 B.n175 VSUBS 0.009902f
C213 B.n176 VSUBS 0.009902f
C214 B.n177 VSUBS 0.009902f
C215 B.n178 VSUBS 0.009902f
C216 B.n179 VSUBS 0.009902f
C217 B.n180 VSUBS 0.009902f
C218 B.n181 VSUBS 0.009902f
C219 B.n182 VSUBS 0.009902f
C220 B.n183 VSUBS 0.009902f
C221 B.n184 VSUBS 0.009902f
C222 B.n185 VSUBS 0.009902f
C223 B.n186 VSUBS 0.009902f
C224 B.n187 VSUBS 0.009902f
C225 B.n188 VSUBS 0.024852f
C226 B.n189 VSUBS 0.009902f
C227 B.n190 VSUBS 0.009902f
C228 B.n191 VSUBS 0.009902f
C229 B.n192 VSUBS 0.009902f
C230 B.n193 VSUBS 0.009902f
C231 B.n194 VSUBS 0.009902f
C232 B.n195 VSUBS 0.009902f
C233 B.n196 VSUBS 0.009902f
C234 B.n197 VSUBS 0.009902f
C235 B.n198 VSUBS 0.009902f
C236 B.n199 VSUBS 0.009902f
C237 B.n200 VSUBS 0.009902f
C238 B.n201 VSUBS 0.009902f
C239 B.n202 VSUBS 0.009902f
C240 B.n203 VSUBS 0.009902f
C241 B.n204 VSUBS 0.009902f
C242 B.n205 VSUBS 0.009902f
C243 B.n206 VSUBS 0.009902f
C244 B.n207 VSUBS 0.009902f
C245 B.n208 VSUBS 0.009902f
C246 B.n209 VSUBS 0.009902f
C247 B.n210 VSUBS 0.009902f
C248 B.n211 VSUBS 0.009902f
C249 B.n212 VSUBS 0.009902f
C250 B.n213 VSUBS 0.009902f
C251 B.n214 VSUBS 0.009902f
C252 B.n215 VSUBS 0.009902f
C253 B.n216 VSUBS 0.009902f
C254 B.n217 VSUBS 0.009902f
C255 B.n218 VSUBS 0.009902f
C256 B.n219 VSUBS 0.009902f
C257 B.n220 VSUBS 0.009902f
C258 B.n221 VSUBS 0.009902f
C259 B.n222 VSUBS 0.009902f
C260 B.n223 VSUBS 0.009902f
C261 B.n224 VSUBS 0.009902f
C262 B.n225 VSUBS 0.009902f
C263 B.n226 VSUBS 0.009902f
C264 B.n227 VSUBS 0.009902f
C265 B.n228 VSUBS 0.009902f
C266 B.n229 VSUBS 0.009902f
C267 B.n230 VSUBS 0.009902f
C268 B.n231 VSUBS 0.009902f
C269 B.n232 VSUBS 0.009902f
C270 B.n233 VSUBS 0.009902f
C271 B.n234 VSUBS 0.009902f
C272 B.n235 VSUBS 0.009902f
C273 B.n236 VSUBS 0.009902f
C274 B.n237 VSUBS 0.009902f
C275 B.n238 VSUBS 0.009902f
C276 B.n239 VSUBS 0.009902f
C277 B.n240 VSUBS 0.009902f
C278 B.n241 VSUBS 0.009902f
C279 B.n242 VSUBS 0.009902f
C280 B.n243 VSUBS 0.009902f
C281 B.n244 VSUBS 0.009902f
C282 B.n245 VSUBS 0.009902f
C283 B.n246 VSUBS 0.009902f
C284 B.n247 VSUBS 0.009902f
C285 B.n248 VSUBS 0.009902f
C286 B.n249 VSUBS 0.009902f
C287 B.n250 VSUBS 0.009902f
C288 B.n251 VSUBS 0.009902f
C289 B.n252 VSUBS 0.009902f
C290 B.n253 VSUBS 0.009902f
C291 B.n254 VSUBS 0.009902f
C292 B.n255 VSUBS 0.009902f
C293 B.n256 VSUBS 0.009902f
C294 B.n257 VSUBS 0.009902f
C295 B.n258 VSUBS 0.009902f
C296 B.n259 VSUBS 0.009902f
C297 B.n260 VSUBS 0.009902f
C298 B.n261 VSUBS 0.009902f
C299 B.n262 VSUBS 0.009902f
C300 B.n263 VSUBS 0.009902f
C301 B.n264 VSUBS 0.009902f
C302 B.n265 VSUBS 0.009902f
C303 B.n266 VSUBS 0.009902f
C304 B.n267 VSUBS 0.009902f
C305 B.n268 VSUBS 0.009902f
C306 B.n269 VSUBS 0.009902f
C307 B.n270 VSUBS 0.009902f
C308 B.n271 VSUBS 0.009902f
C309 B.n272 VSUBS 0.009902f
C310 B.n273 VSUBS 0.009902f
C311 B.n274 VSUBS 0.009902f
C312 B.n275 VSUBS 0.009902f
C313 B.n276 VSUBS 0.009902f
C314 B.n277 VSUBS 0.009902f
C315 B.n278 VSUBS 0.009902f
C316 B.n279 VSUBS 0.009902f
C317 B.n280 VSUBS 0.009902f
C318 B.n281 VSUBS 0.009902f
C319 B.n282 VSUBS 0.009902f
C320 B.n283 VSUBS 0.009902f
C321 B.n284 VSUBS 0.009902f
C322 B.n285 VSUBS 0.009902f
C323 B.n286 VSUBS 0.009902f
C324 B.n287 VSUBS 0.009902f
C325 B.n288 VSUBS 0.009902f
C326 B.n289 VSUBS 0.009902f
C327 B.n290 VSUBS 0.009902f
C328 B.n291 VSUBS 0.009902f
C329 B.n292 VSUBS 0.009902f
C330 B.n293 VSUBS 0.009902f
C331 B.n294 VSUBS 0.009902f
C332 B.n295 VSUBS 0.009902f
C333 B.n296 VSUBS 0.009902f
C334 B.n297 VSUBS 0.009902f
C335 B.n298 VSUBS 0.009902f
C336 B.n299 VSUBS 0.009902f
C337 B.n300 VSUBS 0.009902f
C338 B.n301 VSUBS 0.009902f
C339 B.n302 VSUBS 0.009902f
C340 B.n303 VSUBS 0.009902f
C341 B.n304 VSUBS 0.009902f
C342 B.n305 VSUBS 0.009902f
C343 B.n306 VSUBS 0.009902f
C344 B.n307 VSUBS 0.009902f
C345 B.n308 VSUBS 0.009902f
C346 B.n309 VSUBS 0.009902f
C347 B.n310 VSUBS 0.009902f
C348 B.n311 VSUBS 0.009902f
C349 B.n312 VSUBS 0.009902f
C350 B.n313 VSUBS 0.009902f
C351 B.n314 VSUBS 0.009902f
C352 B.n315 VSUBS 0.009902f
C353 B.n316 VSUBS 0.009902f
C354 B.n317 VSUBS 0.009902f
C355 B.n318 VSUBS 0.009902f
C356 B.n319 VSUBS 0.023204f
C357 B.n320 VSUBS 0.023204f
C358 B.n321 VSUBS 0.024852f
C359 B.n322 VSUBS 0.009902f
C360 B.n323 VSUBS 0.009902f
C361 B.n324 VSUBS 0.009902f
C362 B.n325 VSUBS 0.009902f
C363 B.n326 VSUBS 0.009902f
C364 B.n327 VSUBS 0.009902f
C365 B.n328 VSUBS 0.009902f
C366 B.n329 VSUBS 0.009902f
C367 B.n330 VSUBS 0.009902f
C368 B.n331 VSUBS 0.009902f
C369 B.n332 VSUBS 0.009902f
C370 B.n333 VSUBS 0.009902f
C371 B.n334 VSUBS 0.009902f
C372 B.n335 VSUBS 0.009902f
C373 B.n336 VSUBS 0.009902f
C374 B.n337 VSUBS 0.009902f
C375 B.n338 VSUBS 0.009902f
C376 B.n339 VSUBS 0.009902f
C377 B.n340 VSUBS 0.009902f
C378 B.n341 VSUBS 0.009902f
C379 B.n342 VSUBS 0.009902f
C380 B.n343 VSUBS 0.009902f
C381 B.n344 VSUBS 0.009902f
C382 B.n345 VSUBS 0.009902f
C383 B.n346 VSUBS 0.009902f
C384 B.n347 VSUBS 0.009902f
C385 B.n348 VSUBS 0.009902f
C386 B.n349 VSUBS 0.009902f
C387 B.n350 VSUBS 0.009902f
C388 B.n351 VSUBS 0.009902f
C389 B.n352 VSUBS 0.009902f
C390 B.n353 VSUBS 0.009902f
C391 B.n354 VSUBS 0.009902f
C392 B.n355 VSUBS 0.009902f
C393 B.n356 VSUBS 0.009902f
C394 B.n357 VSUBS 0.009902f
C395 B.n358 VSUBS 0.009902f
C396 B.n359 VSUBS 0.009902f
C397 B.n360 VSUBS 0.009902f
C398 B.n361 VSUBS 0.009902f
C399 B.n362 VSUBS 0.009902f
C400 B.n363 VSUBS 0.009902f
C401 B.n364 VSUBS 0.009902f
C402 B.n365 VSUBS 0.009902f
C403 B.n366 VSUBS 0.009902f
C404 B.n367 VSUBS 0.009902f
C405 B.n368 VSUBS 0.009902f
C406 B.n369 VSUBS 0.009902f
C407 B.n370 VSUBS 0.009902f
C408 B.n371 VSUBS 0.009902f
C409 B.n372 VSUBS 0.006844f
C410 B.n373 VSUBS 0.022943f
C411 B.n374 VSUBS 0.008009f
C412 B.n375 VSUBS 0.009902f
C413 B.n376 VSUBS 0.009902f
C414 B.n377 VSUBS 0.009902f
C415 B.n378 VSUBS 0.009902f
C416 B.n379 VSUBS 0.009902f
C417 B.n380 VSUBS 0.009902f
C418 B.n381 VSUBS 0.009902f
C419 B.n382 VSUBS 0.009902f
C420 B.n383 VSUBS 0.009902f
C421 B.n384 VSUBS 0.009902f
C422 B.n385 VSUBS 0.009902f
C423 B.t8 VSUBS 0.432282f
C424 B.t7 VSUBS 0.465819f
C425 B.t6 VSUBS 1.93593f
C426 B.n386 VSUBS 0.254103f
C427 B.n387 VSUBS 0.103913f
C428 B.n388 VSUBS 0.022943f
C429 B.n389 VSUBS 0.008009f
C430 B.n390 VSUBS 0.009902f
C431 B.n391 VSUBS 0.009902f
C432 B.n392 VSUBS 0.009902f
C433 B.n393 VSUBS 0.009902f
C434 B.n394 VSUBS 0.009902f
C435 B.n395 VSUBS 0.009902f
C436 B.n396 VSUBS 0.009902f
C437 B.n397 VSUBS 0.009902f
C438 B.n398 VSUBS 0.009902f
C439 B.n399 VSUBS 0.009902f
C440 B.n400 VSUBS 0.009902f
C441 B.n401 VSUBS 0.009902f
C442 B.n402 VSUBS 0.009902f
C443 B.n403 VSUBS 0.009902f
C444 B.n404 VSUBS 0.009902f
C445 B.n405 VSUBS 0.009902f
C446 B.n406 VSUBS 0.009902f
C447 B.n407 VSUBS 0.009902f
C448 B.n408 VSUBS 0.009902f
C449 B.n409 VSUBS 0.009902f
C450 B.n410 VSUBS 0.009902f
C451 B.n411 VSUBS 0.009902f
C452 B.n412 VSUBS 0.009902f
C453 B.n413 VSUBS 0.009902f
C454 B.n414 VSUBS 0.009902f
C455 B.n415 VSUBS 0.009902f
C456 B.n416 VSUBS 0.009902f
C457 B.n417 VSUBS 0.009902f
C458 B.n418 VSUBS 0.009902f
C459 B.n419 VSUBS 0.009902f
C460 B.n420 VSUBS 0.009902f
C461 B.n421 VSUBS 0.009902f
C462 B.n422 VSUBS 0.009902f
C463 B.n423 VSUBS 0.009902f
C464 B.n424 VSUBS 0.009902f
C465 B.n425 VSUBS 0.009902f
C466 B.n426 VSUBS 0.009902f
C467 B.n427 VSUBS 0.009902f
C468 B.n428 VSUBS 0.009902f
C469 B.n429 VSUBS 0.009902f
C470 B.n430 VSUBS 0.009902f
C471 B.n431 VSUBS 0.009902f
C472 B.n432 VSUBS 0.009902f
C473 B.n433 VSUBS 0.009902f
C474 B.n434 VSUBS 0.009902f
C475 B.n435 VSUBS 0.009902f
C476 B.n436 VSUBS 0.009902f
C477 B.n437 VSUBS 0.009902f
C478 B.n438 VSUBS 0.009902f
C479 B.n439 VSUBS 0.009902f
C480 B.n440 VSUBS 0.009902f
C481 B.n441 VSUBS 0.009902f
C482 B.n442 VSUBS 0.023744f
C483 B.n443 VSUBS 0.024312f
C484 B.n444 VSUBS 0.023204f
C485 B.n445 VSUBS 0.009902f
C486 B.n446 VSUBS 0.009902f
C487 B.n447 VSUBS 0.009902f
C488 B.n448 VSUBS 0.009902f
C489 B.n449 VSUBS 0.009902f
C490 B.n450 VSUBS 0.009902f
C491 B.n451 VSUBS 0.009902f
C492 B.n452 VSUBS 0.009902f
C493 B.n453 VSUBS 0.009902f
C494 B.n454 VSUBS 0.009902f
C495 B.n455 VSUBS 0.009902f
C496 B.n456 VSUBS 0.009902f
C497 B.n457 VSUBS 0.009902f
C498 B.n458 VSUBS 0.009902f
C499 B.n459 VSUBS 0.009902f
C500 B.n460 VSUBS 0.009902f
C501 B.n461 VSUBS 0.009902f
C502 B.n462 VSUBS 0.009902f
C503 B.n463 VSUBS 0.009902f
C504 B.n464 VSUBS 0.009902f
C505 B.n465 VSUBS 0.009902f
C506 B.n466 VSUBS 0.009902f
C507 B.n467 VSUBS 0.009902f
C508 B.n468 VSUBS 0.009902f
C509 B.n469 VSUBS 0.009902f
C510 B.n470 VSUBS 0.009902f
C511 B.n471 VSUBS 0.009902f
C512 B.n472 VSUBS 0.009902f
C513 B.n473 VSUBS 0.009902f
C514 B.n474 VSUBS 0.009902f
C515 B.n475 VSUBS 0.009902f
C516 B.n476 VSUBS 0.009902f
C517 B.n477 VSUBS 0.009902f
C518 B.n478 VSUBS 0.009902f
C519 B.n479 VSUBS 0.009902f
C520 B.n480 VSUBS 0.009902f
C521 B.n481 VSUBS 0.009902f
C522 B.n482 VSUBS 0.009902f
C523 B.n483 VSUBS 0.009902f
C524 B.n484 VSUBS 0.009902f
C525 B.n485 VSUBS 0.009902f
C526 B.n486 VSUBS 0.009902f
C527 B.n487 VSUBS 0.009902f
C528 B.n488 VSUBS 0.009902f
C529 B.n489 VSUBS 0.009902f
C530 B.n490 VSUBS 0.009902f
C531 B.n491 VSUBS 0.009902f
C532 B.n492 VSUBS 0.009902f
C533 B.n493 VSUBS 0.009902f
C534 B.n494 VSUBS 0.009902f
C535 B.n495 VSUBS 0.009902f
C536 B.n496 VSUBS 0.009902f
C537 B.n497 VSUBS 0.009902f
C538 B.n498 VSUBS 0.009902f
C539 B.n499 VSUBS 0.009902f
C540 B.n500 VSUBS 0.009902f
C541 B.n501 VSUBS 0.009902f
C542 B.n502 VSUBS 0.009902f
C543 B.n503 VSUBS 0.009902f
C544 B.n504 VSUBS 0.009902f
C545 B.n505 VSUBS 0.009902f
C546 B.n506 VSUBS 0.009902f
C547 B.n507 VSUBS 0.009902f
C548 B.n508 VSUBS 0.009902f
C549 B.n509 VSUBS 0.009902f
C550 B.n510 VSUBS 0.009902f
C551 B.n511 VSUBS 0.009902f
C552 B.n512 VSUBS 0.009902f
C553 B.n513 VSUBS 0.009902f
C554 B.n514 VSUBS 0.009902f
C555 B.n515 VSUBS 0.009902f
C556 B.n516 VSUBS 0.009902f
C557 B.n517 VSUBS 0.009902f
C558 B.n518 VSUBS 0.009902f
C559 B.n519 VSUBS 0.009902f
C560 B.n520 VSUBS 0.009902f
C561 B.n521 VSUBS 0.009902f
C562 B.n522 VSUBS 0.009902f
C563 B.n523 VSUBS 0.009902f
C564 B.n524 VSUBS 0.009902f
C565 B.n525 VSUBS 0.009902f
C566 B.n526 VSUBS 0.009902f
C567 B.n527 VSUBS 0.009902f
C568 B.n528 VSUBS 0.009902f
C569 B.n529 VSUBS 0.009902f
C570 B.n530 VSUBS 0.009902f
C571 B.n531 VSUBS 0.009902f
C572 B.n532 VSUBS 0.009902f
C573 B.n533 VSUBS 0.009902f
C574 B.n534 VSUBS 0.009902f
C575 B.n535 VSUBS 0.009902f
C576 B.n536 VSUBS 0.009902f
C577 B.n537 VSUBS 0.009902f
C578 B.n538 VSUBS 0.009902f
C579 B.n539 VSUBS 0.009902f
C580 B.n540 VSUBS 0.009902f
C581 B.n541 VSUBS 0.009902f
C582 B.n542 VSUBS 0.009902f
C583 B.n543 VSUBS 0.009902f
C584 B.n544 VSUBS 0.009902f
C585 B.n545 VSUBS 0.009902f
C586 B.n546 VSUBS 0.009902f
C587 B.n547 VSUBS 0.009902f
C588 B.n548 VSUBS 0.009902f
C589 B.n549 VSUBS 0.009902f
C590 B.n550 VSUBS 0.009902f
C591 B.n551 VSUBS 0.009902f
C592 B.n552 VSUBS 0.009902f
C593 B.n553 VSUBS 0.009902f
C594 B.n554 VSUBS 0.009902f
C595 B.n555 VSUBS 0.009902f
C596 B.n556 VSUBS 0.009902f
C597 B.n557 VSUBS 0.009902f
C598 B.n558 VSUBS 0.009902f
C599 B.n559 VSUBS 0.009902f
C600 B.n560 VSUBS 0.009902f
C601 B.n561 VSUBS 0.009902f
C602 B.n562 VSUBS 0.009902f
C603 B.n563 VSUBS 0.009902f
C604 B.n564 VSUBS 0.009902f
C605 B.n565 VSUBS 0.009902f
C606 B.n566 VSUBS 0.009902f
C607 B.n567 VSUBS 0.009902f
C608 B.n568 VSUBS 0.009902f
C609 B.n569 VSUBS 0.009902f
C610 B.n570 VSUBS 0.009902f
C611 B.n571 VSUBS 0.009902f
C612 B.n572 VSUBS 0.009902f
C613 B.n573 VSUBS 0.009902f
C614 B.n574 VSUBS 0.009902f
C615 B.n575 VSUBS 0.009902f
C616 B.n576 VSUBS 0.009902f
C617 B.n577 VSUBS 0.009902f
C618 B.n578 VSUBS 0.009902f
C619 B.n579 VSUBS 0.009902f
C620 B.n580 VSUBS 0.009902f
C621 B.n581 VSUBS 0.009902f
C622 B.n582 VSUBS 0.009902f
C623 B.n583 VSUBS 0.009902f
C624 B.n584 VSUBS 0.009902f
C625 B.n585 VSUBS 0.009902f
C626 B.n586 VSUBS 0.009902f
C627 B.n587 VSUBS 0.009902f
C628 B.n588 VSUBS 0.009902f
C629 B.n589 VSUBS 0.009902f
C630 B.n590 VSUBS 0.009902f
C631 B.n591 VSUBS 0.009902f
C632 B.n592 VSUBS 0.009902f
C633 B.n593 VSUBS 0.009902f
C634 B.n594 VSUBS 0.009902f
C635 B.n595 VSUBS 0.009902f
C636 B.n596 VSUBS 0.009902f
C637 B.n597 VSUBS 0.009902f
C638 B.n598 VSUBS 0.009902f
C639 B.n599 VSUBS 0.009902f
C640 B.n600 VSUBS 0.009902f
C641 B.n601 VSUBS 0.009902f
C642 B.n602 VSUBS 0.009902f
C643 B.n603 VSUBS 0.009902f
C644 B.n604 VSUBS 0.009902f
C645 B.n605 VSUBS 0.009902f
C646 B.n606 VSUBS 0.009902f
C647 B.n607 VSUBS 0.009902f
C648 B.n608 VSUBS 0.009902f
C649 B.n609 VSUBS 0.009902f
C650 B.n610 VSUBS 0.009902f
C651 B.n611 VSUBS 0.009902f
C652 B.n612 VSUBS 0.009902f
C653 B.n613 VSUBS 0.009902f
C654 B.n614 VSUBS 0.009902f
C655 B.n615 VSUBS 0.009902f
C656 B.n616 VSUBS 0.009902f
C657 B.n617 VSUBS 0.009902f
C658 B.n618 VSUBS 0.009902f
C659 B.n619 VSUBS 0.009902f
C660 B.n620 VSUBS 0.009902f
C661 B.n621 VSUBS 0.009902f
C662 B.n622 VSUBS 0.009902f
C663 B.n623 VSUBS 0.009902f
C664 B.n624 VSUBS 0.009902f
C665 B.n625 VSUBS 0.009902f
C666 B.n626 VSUBS 0.009902f
C667 B.n627 VSUBS 0.009902f
C668 B.n628 VSUBS 0.009902f
C669 B.n629 VSUBS 0.009902f
C670 B.n630 VSUBS 0.009902f
C671 B.n631 VSUBS 0.009902f
C672 B.n632 VSUBS 0.009902f
C673 B.n633 VSUBS 0.009902f
C674 B.n634 VSUBS 0.009902f
C675 B.n635 VSUBS 0.009902f
C676 B.n636 VSUBS 0.009902f
C677 B.n637 VSUBS 0.009902f
C678 B.n638 VSUBS 0.009902f
C679 B.n639 VSUBS 0.009902f
C680 B.n640 VSUBS 0.009902f
C681 B.n641 VSUBS 0.009902f
C682 B.n642 VSUBS 0.009902f
C683 B.n643 VSUBS 0.009902f
C684 B.n644 VSUBS 0.009902f
C685 B.n645 VSUBS 0.009902f
C686 B.n646 VSUBS 0.023204f
C687 B.n647 VSUBS 0.024852f
C688 B.n648 VSUBS 0.024852f
C689 B.n649 VSUBS 0.009902f
C690 B.n650 VSUBS 0.009902f
C691 B.n651 VSUBS 0.009902f
C692 B.n652 VSUBS 0.009902f
C693 B.n653 VSUBS 0.009902f
C694 B.n654 VSUBS 0.009902f
C695 B.n655 VSUBS 0.009902f
C696 B.n656 VSUBS 0.009902f
C697 B.n657 VSUBS 0.009902f
C698 B.n658 VSUBS 0.009902f
C699 B.n659 VSUBS 0.009902f
C700 B.n660 VSUBS 0.009902f
C701 B.n661 VSUBS 0.009902f
C702 B.n662 VSUBS 0.009902f
C703 B.n663 VSUBS 0.009902f
C704 B.n664 VSUBS 0.009902f
C705 B.n665 VSUBS 0.009902f
C706 B.n666 VSUBS 0.009902f
C707 B.n667 VSUBS 0.009902f
C708 B.n668 VSUBS 0.009902f
C709 B.n669 VSUBS 0.009902f
C710 B.n670 VSUBS 0.009902f
C711 B.n671 VSUBS 0.009902f
C712 B.n672 VSUBS 0.009902f
C713 B.n673 VSUBS 0.009902f
C714 B.n674 VSUBS 0.009902f
C715 B.n675 VSUBS 0.009902f
C716 B.n676 VSUBS 0.009902f
C717 B.n677 VSUBS 0.009902f
C718 B.n678 VSUBS 0.009902f
C719 B.n679 VSUBS 0.009902f
C720 B.n680 VSUBS 0.009902f
C721 B.n681 VSUBS 0.009902f
C722 B.n682 VSUBS 0.009902f
C723 B.n683 VSUBS 0.009902f
C724 B.n684 VSUBS 0.009902f
C725 B.n685 VSUBS 0.009902f
C726 B.n686 VSUBS 0.009902f
C727 B.n687 VSUBS 0.009902f
C728 B.n688 VSUBS 0.009902f
C729 B.n689 VSUBS 0.009902f
C730 B.n690 VSUBS 0.009902f
C731 B.n691 VSUBS 0.009902f
C732 B.n692 VSUBS 0.009902f
C733 B.n693 VSUBS 0.009902f
C734 B.n694 VSUBS 0.009902f
C735 B.n695 VSUBS 0.009902f
C736 B.n696 VSUBS 0.009902f
C737 B.n697 VSUBS 0.009902f
C738 B.n698 VSUBS 0.009902f
C739 B.n699 VSUBS 0.006844f
C740 B.n700 VSUBS 0.022943f
C741 B.n701 VSUBS 0.008009f
C742 B.n702 VSUBS 0.009902f
C743 B.n703 VSUBS 0.009902f
C744 B.n704 VSUBS 0.009902f
C745 B.n705 VSUBS 0.009902f
C746 B.n706 VSUBS 0.009902f
C747 B.n707 VSUBS 0.009902f
C748 B.n708 VSUBS 0.009902f
C749 B.n709 VSUBS 0.009902f
C750 B.n710 VSUBS 0.009902f
C751 B.n711 VSUBS 0.009902f
C752 B.n712 VSUBS 0.009902f
C753 B.n713 VSUBS 0.008009f
C754 B.n714 VSUBS 0.022943f
C755 B.n715 VSUBS 0.006844f
C756 B.n716 VSUBS 0.009902f
C757 B.n717 VSUBS 0.009902f
C758 B.n718 VSUBS 0.009902f
C759 B.n719 VSUBS 0.009902f
C760 B.n720 VSUBS 0.009902f
C761 B.n721 VSUBS 0.009902f
C762 B.n722 VSUBS 0.009902f
C763 B.n723 VSUBS 0.009902f
C764 B.n724 VSUBS 0.009902f
C765 B.n725 VSUBS 0.009902f
C766 B.n726 VSUBS 0.009902f
C767 B.n727 VSUBS 0.009902f
C768 B.n728 VSUBS 0.009902f
C769 B.n729 VSUBS 0.009902f
C770 B.n730 VSUBS 0.009902f
C771 B.n731 VSUBS 0.009902f
C772 B.n732 VSUBS 0.009902f
C773 B.n733 VSUBS 0.009902f
C774 B.n734 VSUBS 0.009902f
C775 B.n735 VSUBS 0.009902f
C776 B.n736 VSUBS 0.009902f
C777 B.n737 VSUBS 0.009902f
C778 B.n738 VSUBS 0.009902f
C779 B.n739 VSUBS 0.009902f
C780 B.n740 VSUBS 0.009902f
C781 B.n741 VSUBS 0.009902f
C782 B.n742 VSUBS 0.009902f
C783 B.n743 VSUBS 0.009902f
C784 B.n744 VSUBS 0.009902f
C785 B.n745 VSUBS 0.009902f
C786 B.n746 VSUBS 0.009902f
C787 B.n747 VSUBS 0.009902f
C788 B.n748 VSUBS 0.009902f
C789 B.n749 VSUBS 0.009902f
C790 B.n750 VSUBS 0.009902f
C791 B.n751 VSUBS 0.009902f
C792 B.n752 VSUBS 0.009902f
C793 B.n753 VSUBS 0.009902f
C794 B.n754 VSUBS 0.009902f
C795 B.n755 VSUBS 0.009902f
C796 B.n756 VSUBS 0.009902f
C797 B.n757 VSUBS 0.009902f
C798 B.n758 VSUBS 0.009902f
C799 B.n759 VSUBS 0.009902f
C800 B.n760 VSUBS 0.009902f
C801 B.n761 VSUBS 0.009902f
C802 B.n762 VSUBS 0.009902f
C803 B.n763 VSUBS 0.009902f
C804 B.n764 VSUBS 0.009902f
C805 B.n765 VSUBS 0.009902f
C806 B.n766 VSUBS 0.024852f
C807 B.n767 VSUBS 0.024852f
C808 B.n768 VSUBS 0.023204f
C809 B.n769 VSUBS 0.009902f
C810 B.n770 VSUBS 0.009902f
C811 B.n771 VSUBS 0.009902f
C812 B.n772 VSUBS 0.009902f
C813 B.n773 VSUBS 0.009902f
C814 B.n774 VSUBS 0.009902f
C815 B.n775 VSUBS 0.009902f
C816 B.n776 VSUBS 0.009902f
C817 B.n777 VSUBS 0.009902f
C818 B.n778 VSUBS 0.009902f
C819 B.n779 VSUBS 0.009902f
C820 B.n780 VSUBS 0.009902f
C821 B.n781 VSUBS 0.009902f
C822 B.n782 VSUBS 0.009902f
C823 B.n783 VSUBS 0.009902f
C824 B.n784 VSUBS 0.009902f
C825 B.n785 VSUBS 0.009902f
C826 B.n786 VSUBS 0.009902f
C827 B.n787 VSUBS 0.009902f
C828 B.n788 VSUBS 0.009902f
C829 B.n789 VSUBS 0.009902f
C830 B.n790 VSUBS 0.009902f
C831 B.n791 VSUBS 0.009902f
C832 B.n792 VSUBS 0.009902f
C833 B.n793 VSUBS 0.009902f
C834 B.n794 VSUBS 0.009902f
C835 B.n795 VSUBS 0.009902f
C836 B.n796 VSUBS 0.009902f
C837 B.n797 VSUBS 0.009902f
C838 B.n798 VSUBS 0.009902f
C839 B.n799 VSUBS 0.009902f
C840 B.n800 VSUBS 0.009902f
C841 B.n801 VSUBS 0.009902f
C842 B.n802 VSUBS 0.009902f
C843 B.n803 VSUBS 0.009902f
C844 B.n804 VSUBS 0.009902f
C845 B.n805 VSUBS 0.009902f
C846 B.n806 VSUBS 0.009902f
C847 B.n807 VSUBS 0.009902f
C848 B.n808 VSUBS 0.009902f
C849 B.n809 VSUBS 0.009902f
C850 B.n810 VSUBS 0.009902f
C851 B.n811 VSUBS 0.009902f
C852 B.n812 VSUBS 0.009902f
C853 B.n813 VSUBS 0.009902f
C854 B.n814 VSUBS 0.009902f
C855 B.n815 VSUBS 0.009902f
C856 B.n816 VSUBS 0.009902f
C857 B.n817 VSUBS 0.009902f
C858 B.n818 VSUBS 0.009902f
C859 B.n819 VSUBS 0.009902f
C860 B.n820 VSUBS 0.009902f
C861 B.n821 VSUBS 0.009902f
C862 B.n822 VSUBS 0.009902f
C863 B.n823 VSUBS 0.009902f
C864 B.n824 VSUBS 0.009902f
C865 B.n825 VSUBS 0.009902f
C866 B.n826 VSUBS 0.009902f
C867 B.n827 VSUBS 0.009902f
C868 B.n828 VSUBS 0.009902f
C869 B.n829 VSUBS 0.009902f
C870 B.n830 VSUBS 0.009902f
C871 B.n831 VSUBS 0.009902f
C872 B.n832 VSUBS 0.009902f
C873 B.n833 VSUBS 0.009902f
C874 B.n834 VSUBS 0.009902f
C875 B.n835 VSUBS 0.009902f
C876 B.n836 VSUBS 0.009902f
C877 B.n837 VSUBS 0.009902f
C878 B.n838 VSUBS 0.009902f
C879 B.n839 VSUBS 0.009902f
C880 B.n840 VSUBS 0.009902f
C881 B.n841 VSUBS 0.009902f
C882 B.n842 VSUBS 0.009902f
C883 B.n843 VSUBS 0.009902f
C884 B.n844 VSUBS 0.009902f
C885 B.n845 VSUBS 0.009902f
C886 B.n846 VSUBS 0.009902f
C887 B.n847 VSUBS 0.009902f
C888 B.n848 VSUBS 0.009902f
C889 B.n849 VSUBS 0.009902f
C890 B.n850 VSUBS 0.009902f
C891 B.n851 VSUBS 0.009902f
C892 B.n852 VSUBS 0.009902f
C893 B.n853 VSUBS 0.009902f
C894 B.n854 VSUBS 0.009902f
C895 B.n855 VSUBS 0.009902f
C896 B.n856 VSUBS 0.009902f
C897 B.n857 VSUBS 0.009902f
C898 B.n858 VSUBS 0.009902f
C899 B.n859 VSUBS 0.009902f
C900 B.n860 VSUBS 0.009902f
C901 B.n861 VSUBS 0.009902f
C902 B.n862 VSUBS 0.009902f
C903 B.n863 VSUBS 0.009902f
C904 B.n864 VSUBS 0.009902f
C905 B.n865 VSUBS 0.009902f
C906 B.n866 VSUBS 0.009902f
C907 B.n867 VSUBS 0.012922f
C908 B.n868 VSUBS 0.013765f
C909 B.n869 VSUBS 0.027374f
C910 VDD1.t9 VSUBS 2.41229f
C911 VDD1.t1 VSUBS 0.241522f
C912 VDD1.t7 VSUBS 0.241522f
C913 VDD1.n0 VSUBS 1.81226f
C914 VDD1.n1 VSUBS 1.8811f
C915 VDD1.t3 VSUBS 2.41227f
C916 VDD1.t6 VSUBS 0.241522f
C917 VDD1.t5 VSUBS 0.241522f
C918 VDD1.n2 VSUBS 1.81225f
C919 VDD1.n3 VSUBS 1.8706f
C920 VDD1.t0 VSUBS 0.241522f
C921 VDD1.t4 VSUBS 0.241522f
C922 VDD1.n4 VSUBS 1.84123f
C923 VDD1.n5 VSUBS 4.27481f
C924 VDD1.t2 VSUBS 0.241522f
C925 VDD1.t8 VSUBS 0.241522f
C926 VDD1.n6 VSUBS 1.81225f
C927 VDD1.n7 VSUBS 4.34079f
C928 VP.n0 VSUBS 0.04033f
C929 VP.t5 VSUBS 2.4308f
C930 VP.n1 VSUBS 0.057012f
C931 VP.n2 VSUBS 0.03059f
C932 VP.n3 VSUBS 0.049694f
C933 VP.n4 VSUBS 0.03059f
C934 VP.n5 VSUBS 0.026174f
C935 VP.n6 VSUBS 0.03059f
C936 VP.t4 VSUBS 2.4308f
C937 VP.n7 VSUBS 0.867466f
C938 VP.n8 VSUBS 0.03059f
C939 VP.n9 VSUBS 0.026174f
C940 VP.n10 VSUBS 0.03059f
C941 VP.t3 VSUBS 2.4308f
C942 VP.n11 VSUBS 0.867466f
C943 VP.n12 VSUBS 0.03059f
C944 VP.n13 VSUBS 0.038689f
C945 VP.n14 VSUBS 0.03059f
C946 VP.t6 VSUBS 2.4308f
C947 VP.n15 VSUBS 0.972182f
C948 VP.n16 VSUBS 0.04033f
C949 VP.t1 VSUBS 2.4308f
C950 VP.n17 VSUBS 0.057012f
C951 VP.n18 VSUBS 0.03059f
C952 VP.n19 VSUBS 0.049694f
C953 VP.n20 VSUBS 0.03059f
C954 VP.n21 VSUBS 0.026174f
C955 VP.n22 VSUBS 0.03059f
C956 VP.t2 VSUBS 2.4308f
C957 VP.n23 VSUBS 0.867466f
C958 VP.n24 VSUBS 0.03059f
C959 VP.n25 VSUBS 0.026174f
C960 VP.n26 VSUBS 0.03059f
C961 VP.t8 VSUBS 2.4308f
C962 VP.n27 VSUBS 0.959405f
C963 VP.t0 VSUBS 2.75052f
C964 VP.n28 VSUBS 0.92784f
C965 VP.n29 VSUBS 0.329641f
C966 VP.n30 VSUBS 0.036183f
C967 VP.n31 VSUBS 0.057012f
C968 VP.n32 VSUBS 0.061813f
C969 VP.n33 VSUBS 0.03059f
C970 VP.n34 VSUBS 0.03059f
C971 VP.n35 VSUBS 0.03059f
C972 VP.n36 VSUBS 0.058338f
C973 VP.n37 VSUBS 0.057012f
C974 VP.n38 VSUBS 0.042939f
C975 VP.n39 VSUBS 0.03059f
C976 VP.n40 VSUBS 0.03059f
C977 VP.n41 VSUBS 0.042939f
C978 VP.n42 VSUBS 0.057012f
C979 VP.n43 VSUBS 0.058338f
C980 VP.n44 VSUBS 0.03059f
C981 VP.n45 VSUBS 0.03059f
C982 VP.n46 VSUBS 0.03059f
C983 VP.n47 VSUBS 0.061813f
C984 VP.n48 VSUBS 0.057012f
C985 VP.t7 VSUBS 2.4308f
C986 VP.n49 VSUBS 0.867466f
C987 VP.n50 VSUBS 0.036183f
C988 VP.n51 VSUBS 0.03059f
C989 VP.n52 VSUBS 0.03059f
C990 VP.n53 VSUBS 0.03059f
C991 VP.n54 VSUBS 0.057012f
C992 VP.n55 VSUBS 0.050623f
C993 VP.n56 VSUBS 0.038689f
C994 VP.n57 VSUBS 0.03059f
C995 VP.n58 VSUBS 0.03059f
C996 VP.n59 VSUBS 0.03059f
C997 VP.n60 VSUBS 0.057012f
C998 VP.n61 VSUBS 0.029428f
C999 VP.n62 VSUBS 0.972182f
C1000 VP.n63 VSUBS 1.90209f
C1001 VP.n64 VSUBS 1.92255f
C1002 VP.n65 VSUBS 0.04033f
C1003 VP.n66 VSUBS 0.029428f
C1004 VP.n67 VSUBS 0.057012f
C1005 VP.n68 VSUBS 0.057012f
C1006 VP.n69 VSUBS 0.03059f
C1007 VP.n70 VSUBS 0.03059f
C1008 VP.n71 VSUBS 0.03059f
C1009 VP.n72 VSUBS 0.050623f
C1010 VP.n73 VSUBS 0.057012f
C1011 VP.n74 VSUBS 0.049694f
C1012 VP.n75 VSUBS 0.03059f
C1013 VP.n76 VSUBS 0.03059f
C1014 VP.n77 VSUBS 0.036183f
C1015 VP.n78 VSUBS 0.057012f
C1016 VP.n79 VSUBS 0.061813f
C1017 VP.n80 VSUBS 0.03059f
C1018 VP.n81 VSUBS 0.03059f
C1019 VP.n82 VSUBS 0.03059f
C1020 VP.n83 VSUBS 0.058338f
C1021 VP.n84 VSUBS 0.057012f
C1022 VP.n85 VSUBS 0.042939f
C1023 VP.n86 VSUBS 0.03059f
C1024 VP.n87 VSUBS 0.03059f
C1025 VP.n88 VSUBS 0.042939f
C1026 VP.n89 VSUBS 0.057012f
C1027 VP.n90 VSUBS 0.058338f
C1028 VP.n91 VSUBS 0.03059f
C1029 VP.n92 VSUBS 0.03059f
C1030 VP.n93 VSUBS 0.03059f
C1031 VP.n94 VSUBS 0.061813f
C1032 VP.n95 VSUBS 0.057012f
C1033 VP.t9 VSUBS 2.4308f
C1034 VP.n96 VSUBS 0.867466f
C1035 VP.n97 VSUBS 0.036183f
C1036 VP.n98 VSUBS 0.03059f
C1037 VP.n99 VSUBS 0.03059f
C1038 VP.n100 VSUBS 0.03059f
C1039 VP.n101 VSUBS 0.057012f
C1040 VP.n102 VSUBS 0.050623f
C1041 VP.n103 VSUBS 0.038689f
C1042 VP.n104 VSUBS 0.03059f
C1043 VP.n105 VSUBS 0.03059f
C1044 VP.n106 VSUBS 0.03059f
C1045 VP.n107 VSUBS 0.057012f
C1046 VP.n108 VSUBS 0.029428f
C1047 VP.n109 VSUBS 0.972182f
C1048 VP.n110 VSUBS 0.061797f
C1049 VTAIL.t10 VSUBS 0.232311f
C1050 VTAIL.t5 VSUBS 0.232311f
C1051 VTAIL.n0 VSUBS 1.59743f
C1052 VTAIL.n1 VSUBS 1.05944f
C1053 VTAIL.t17 VSUBS 2.12737f
C1054 VTAIL.n2 VSUBS 1.22901f
C1055 VTAIL.t15 VSUBS 0.232311f
C1056 VTAIL.t16 VSUBS 0.232311f
C1057 VTAIL.n3 VSUBS 1.59743f
C1058 VTAIL.n4 VSUBS 1.22246f
C1059 VTAIL.t0 VSUBS 0.232311f
C1060 VTAIL.t18 VSUBS 0.232311f
C1061 VTAIL.n5 VSUBS 1.59743f
C1062 VTAIL.n6 VSUBS 2.74037f
C1063 VTAIL.t3 VSUBS 0.232311f
C1064 VTAIL.t11 VSUBS 0.232311f
C1065 VTAIL.n7 VSUBS 1.59744f
C1066 VTAIL.n8 VSUBS 2.74036f
C1067 VTAIL.t4 VSUBS 0.232311f
C1068 VTAIL.t12 VSUBS 0.232311f
C1069 VTAIL.n9 VSUBS 1.59744f
C1070 VTAIL.n10 VSUBS 1.22246f
C1071 VTAIL.t6 VSUBS 2.12738f
C1072 VTAIL.n11 VSUBS 1.22899f
C1073 VTAIL.t2 VSUBS 0.232311f
C1074 VTAIL.t19 VSUBS 0.232311f
C1075 VTAIL.n12 VSUBS 1.59744f
C1076 VTAIL.n13 VSUBS 1.12536f
C1077 VTAIL.t13 VSUBS 0.232311f
C1078 VTAIL.t14 VSUBS 0.232311f
C1079 VTAIL.n14 VSUBS 1.59744f
C1080 VTAIL.n15 VSUBS 1.22246f
C1081 VTAIL.t1 VSUBS 2.12737f
C1082 VTAIL.n16 VSUBS 2.55739f
C1083 VTAIL.t9 VSUBS 2.12737f
C1084 VTAIL.n17 VSUBS 2.55739f
C1085 VTAIL.t7 VSUBS 0.232311f
C1086 VTAIL.t8 VSUBS 0.232311f
C1087 VTAIL.n18 VSUBS 1.59743f
C1088 VTAIL.n19 VSUBS 1.00178f
C1089 VDD2.t2 VSUBS 2.41384f
C1090 VDD2.t0 VSUBS 0.241678f
C1091 VDD2.t1 VSUBS 0.241678f
C1092 VDD2.n0 VSUBS 1.81342f
C1093 VDD2.n1 VSUBS 1.87181f
C1094 VDD2.t5 VSUBS 0.241678f
C1095 VDD2.t3 VSUBS 0.241678f
C1096 VDD2.n2 VSUBS 1.84242f
C1097 VDD2.n3 VSUBS 4.10554f
C1098 VDD2.t4 VSUBS 2.38048f
C1099 VDD2.n4 VSUBS 4.27274f
C1100 VDD2.t8 VSUBS 0.241678f
C1101 VDD2.t7 VSUBS 0.241678f
C1102 VDD2.n5 VSUBS 1.81343f
C1103 VDD2.n6 VSUBS 0.945662f
C1104 VDD2.t6 VSUBS 0.241678f
C1105 VDD2.t9 VSUBS 0.241678f
C1106 VDD2.n7 VSUBS 1.84236f
C1107 VN.n0 VSUBS 0.036731f
C1108 VN.t3 VSUBS 2.21388f
C1109 VN.n1 VSUBS 0.051925f
C1110 VN.n2 VSUBS 0.02786f
C1111 VN.n3 VSUBS 0.045259f
C1112 VN.n4 VSUBS 0.02786f
C1113 VN.n5 VSUBS 0.023838f
C1114 VN.n6 VSUBS 0.02786f
C1115 VN.t5 VSUBS 2.21388f
C1116 VN.n7 VSUBS 0.790053f
C1117 VN.n8 VSUBS 0.02786f
C1118 VN.n9 VSUBS 0.023838f
C1119 VN.n10 VSUBS 0.02786f
C1120 VN.t7 VSUBS 2.21388f
C1121 VN.n11 VSUBS 0.873787f
C1122 VN.t2 VSUBS 2.50506f
C1123 VN.n12 VSUBS 0.84504f
C1124 VN.n13 VSUBS 0.300224f
C1125 VN.n14 VSUBS 0.032954f
C1126 VN.n15 VSUBS 0.051925f
C1127 VN.n16 VSUBS 0.056297f
C1128 VN.n17 VSUBS 0.02786f
C1129 VN.n18 VSUBS 0.02786f
C1130 VN.n19 VSUBS 0.02786f
C1131 VN.n20 VSUBS 0.053132f
C1132 VN.n21 VSUBS 0.051925f
C1133 VN.n22 VSUBS 0.039107f
C1134 VN.n23 VSUBS 0.02786f
C1135 VN.n24 VSUBS 0.02786f
C1136 VN.n25 VSUBS 0.039107f
C1137 VN.n26 VSUBS 0.051925f
C1138 VN.n27 VSUBS 0.053132f
C1139 VN.n28 VSUBS 0.02786f
C1140 VN.n29 VSUBS 0.02786f
C1141 VN.n30 VSUBS 0.02786f
C1142 VN.n31 VSUBS 0.056297f
C1143 VN.n32 VSUBS 0.051925f
C1144 VN.t4 VSUBS 2.21388f
C1145 VN.n33 VSUBS 0.790053f
C1146 VN.n34 VSUBS 0.032954f
C1147 VN.n35 VSUBS 0.02786f
C1148 VN.n36 VSUBS 0.02786f
C1149 VN.n37 VSUBS 0.02786f
C1150 VN.n38 VSUBS 0.051925f
C1151 VN.n39 VSUBS 0.046106f
C1152 VN.n40 VSUBS 0.035237f
C1153 VN.n41 VSUBS 0.02786f
C1154 VN.n42 VSUBS 0.02786f
C1155 VN.n43 VSUBS 0.02786f
C1156 VN.n44 VSUBS 0.051925f
C1157 VN.n45 VSUBS 0.026802f
C1158 VN.n46 VSUBS 0.885425f
C1159 VN.n47 VSUBS 0.056283f
C1160 VN.n48 VSUBS 0.036731f
C1161 VN.t9 VSUBS 2.21388f
C1162 VN.n49 VSUBS 0.051925f
C1163 VN.n50 VSUBS 0.02786f
C1164 VN.n51 VSUBS 0.045259f
C1165 VN.n52 VSUBS 0.02786f
C1166 VN.t1 VSUBS 2.21388f
C1167 VN.n53 VSUBS 0.790053f
C1168 VN.n54 VSUBS 0.023838f
C1169 VN.n55 VSUBS 0.02786f
C1170 VN.t8 VSUBS 2.21388f
C1171 VN.n56 VSUBS 0.790053f
C1172 VN.n57 VSUBS 0.02786f
C1173 VN.n58 VSUBS 0.023838f
C1174 VN.n59 VSUBS 0.02786f
C1175 VN.t0 VSUBS 2.21388f
C1176 VN.n60 VSUBS 0.873787f
C1177 VN.t6 VSUBS 2.50506f
C1178 VN.n61 VSUBS 0.84504f
C1179 VN.n62 VSUBS 0.300224f
C1180 VN.n63 VSUBS 0.032954f
C1181 VN.n64 VSUBS 0.051925f
C1182 VN.n65 VSUBS 0.056297f
C1183 VN.n66 VSUBS 0.02786f
C1184 VN.n67 VSUBS 0.02786f
C1185 VN.n68 VSUBS 0.02786f
C1186 VN.n69 VSUBS 0.053132f
C1187 VN.n70 VSUBS 0.051925f
C1188 VN.n71 VSUBS 0.039107f
C1189 VN.n72 VSUBS 0.02786f
C1190 VN.n73 VSUBS 0.02786f
C1191 VN.n74 VSUBS 0.039107f
C1192 VN.n75 VSUBS 0.051925f
C1193 VN.n76 VSUBS 0.053132f
C1194 VN.n77 VSUBS 0.02786f
C1195 VN.n78 VSUBS 0.02786f
C1196 VN.n79 VSUBS 0.02786f
C1197 VN.n80 VSUBS 0.056297f
C1198 VN.n81 VSUBS 0.051925f
C1199 VN.n82 VSUBS 0.032954f
C1200 VN.n83 VSUBS 0.02786f
C1201 VN.n84 VSUBS 0.02786f
C1202 VN.n85 VSUBS 0.02786f
C1203 VN.n86 VSUBS 0.051925f
C1204 VN.n87 VSUBS 0.046106f
C1205 VN.n88 VSUBS 0.035237f
C1206 VN.n89 VSUBS 0.02786f
C1207 VN.n90 VSUBS 0.02786f
C1208 VN.n91 VSUBS 0.02786f
C1209 VN.n92 VSUBS 0.051925f
C1210 VN.n93 VSUBS 0.026802f
C1211 VN.n94 VSUBS 0.885425f
C1212 VN.n95 VSUBS 1.74715f
.ends

