* NGSPICE file created from diff_pair_sample_0532.ext - technology: sky130A

.subckt diff_pair_sample_0532 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2122_n1998# sky130_fd_pr__pfet_01v8 ad=2.0085 pd=11.08 as=0 ps=0 w=5.15 l=1.11
X1 B.t8 B.t6 B.t7 w_n2122_n1998# sky130_fd_pr__pfet_01v8 ad=2.0085 pd=11.08 as=0 ps=0 w=5.15 l=1.11
X2 VDD1.t5 VP.t0 VTAIL.t9 w_n2122_n1998# sky130_fd_pr__pfet_01v8 ad=2.0085 pd=11.08 as=0.84975 ps=5.48 w=5.15 l=1.11
X3 VDD2.t5 VN.t0 VTAIL.t2 w_n2122_n1998# sky130_fd_pr__pfet_01v8 ad=0.84975 pd=5.48 as=2.0085 ps=11.08 w=5.15 l=1.11
X4 VTAIL.t3 VN.t1 VDD2.t4 w_n2122_n1998# sky130_fd_pr__pfet_01v8 ad=0.84975 pd=5.48 as=0.84975 ps=5.48 w=5.15 l=1.11
X5 VTAIL.t7 VP.t1 VDD1.t4 w_n2122_n1998# sky130_fd_pr__pfet_01v8 ad=0.84975 pd=5.48 as=0.84975 ps=5.48 w=5.15 l=1.11
X6 VDD2.t3 VN.t2 VTAIL.t4 w_n2122_n1998# sky130_fd_pr__pfet_01v8 ad=0.84975 pd=5.48 as=2.0085 ps=11.08 w=5.15 l=1.11
X7 VTAIL.t1 VN.t3 VDD2.t2 w_n2122_n1998# sky130_fd_pr__pfet_01v8 ad=0.84975 pd=5.48 as=0.84975 ps=5.48 w=5.15 l=1.11
X8 VDD2.t1 VN.t4 VTAIL.t5 w_n2122_n1998# sky130_fd_pr__pfet_01v8 ad=2.0085 pd=11.08 as=0.84975 ps=5.48 w=5.15 l=1.11
X9 B.t5 B.t3 B.t4 w_n2122_n1998# sky130_fd_pr__pfet_01v8 ad=2.0085 pd=11.08 as=0 ps=0 w=5.15 l=1.11
X10 VTAIL.t6 VP.t2 VDD1.t3 w_n2122_n1998# sky130_fd_pr__pfet_01v8 ad=0.84975 pd=5.48 as=0.84975 ps=5.48 w=5.15 l=1.11
X11 VDD1.t2 VP.t3 VTAIL.t8 w_n2122_n1998# sky130_fd_pr__pfet_01v8 ad=2.0085 pd=11.08 as=0.84975 ps=5.48 w=5.15 l=1.11
X12 VDD1.t1 VP.t4 VTAIL.t11 w_n2122_n1998# sky130_fd_pr__pfet_01v8 ad=0.84975 pd=5.48 as=2.0085 ps=11.08 w=5.15 l=1.11
X13 B.t2 B.t0 B.t1 w_n2122_n1998# sky130_fd_pr__pfet_01v8 ad=2.0085 pd=11.08 as=0 ps=0 w=5.15 l=1.11
X14 VDD1.t0 VP.t5 VTAIL.t10 w_n2122_n1998# sky130_fd_pr__pfet_01v8 ad=0.84975 pd=5.48 as=2.0085 ps=11.08 w=5.15 l=1.11
X15 VDD2.t0 VN.t5 VTAIL.t0 w_n2122_n1998# sky130_fd_pr__pfet_01v8 ad=2.0085 pd=11.08 as=0.84975 ps=5.48 w=5.15 l=1.11
R0 B.n306 B.n305 585
R1 B.n307 B.n44 585
R2 B.n309 B.n308 585
R3 B.n310 B.n43 585
R4 B.n312 B.n311 585
R5 B.n313 B.n42 585
R6 B.n315 B.n314 585
R7 B.n316 B.n41 585
R8 B.n318 B.n317 585
R9 B.n319 B.n40 585
R10 B.n321 B.n320 585
R11 B.n322 B.n39 585
R12 B.n324 B.n323 585
R13 B.n325 B.n38 585
R14 B.n327 B.n326 585
R15 B.n328 B.n37 585
R16 B.n330 B.n329 585
R17 B.n331 B.n36 585
R18 B.n333 B.n332 585
R19 B.n334 B.n35 585
R20 B.n336 B.n335 585
R21 B.n338 B.n337 585
R22 B.n339 B.n31 585
R23 B.n341 B.n340 585
R24 B.n342 B.n30 585
R25 B.n344 B.n343 585
R26 B.n345 B.n29 585
R27 B.n347 B.n346 585
R28 B.n348 B.n28 585
R29 B.n350 B.n349 585
R30 B.n351 B.n25 585
R31 B.n354 B.n353 585
R32 B.n355 B.n24 585
R33 B.n357 B.n356 585
R34 B.n358 B.n23 585
R35 B.n360 B.n359 585
R36 B.n361 B.n22 585
R37 B.n363 B.n362 585
R38 B.n364 B.n21 585
R39 B.n366 B.n365 585
R40 B.n367 B.n20 585
R41 B.n369 B.n368 585
R42 B.n370 B.n19 585
R43 B.n372 B.n371 585
R44 B.n373 B.n18 585
R45 B.n375 B.n374 585
R46 B.n376 B.n17 585
R47 B.n378 B.n377 585
R48 B.n379 B.n16 585
R49 B.n381 B.n380 585
R50 B.n382 B.n15 585
R51 B.n384 B.n383 585
R52 B.n304 B.n45 585
R53 B.n303 B.n302 585
R54 B.n301 B.n46 585
R55 B.n300 B.n299 585
R56 B.n298 B.n47 585
R57 B.n297 B.n296 585
R58 B.n295 B.n48 585
R59 B.n294 B.n293 585
R60 B.n292 B.n49 585
R61 B.n291 B.n290 585
R62 B.n289 B.n50 585
R63 B.n288 B.n287 585
R64 B.n286 B.n51 585
R65 B.n285 B.n284 585
R66 B.n283 B.n52 585
R67 B.n282 B.n281 585
R68 B.n280 B.n53 585
R69 B.n279 B.n278 585
R70 B.n277 B.n54 585
R71 B.n276 B.n275 585
R72 B.n274 B.n55 585
R73 B.n273 B.n272 585
R74 B.n271 B.n56 585
R75 B.n270 B.n269 585
R76 B.n268 B.n57 585
R77 B.n267 B.n266 585
R78 B.n265 B.n58 585
R79 B.n264 B.n263 585
R80 B.n262 B.n59 585
R81 B.n261 B.n260 585
R82 B.n259 B.n60 585
R83 B.n258 B.n257 585
R84 B.n256 B.n61 585
R85 B.n255 B.n254 585
R86 B.n253 B.n62 585
R87 B.n252 B.n251 585
R88 B.n250 B.n63 585
R89 B.n249 B.n248 585
R90 B.n247 B.n64 585
R91 B.n246 B.n245 585
R92 B.n244 B.n65 585
R93 B.n243 B.n242 585
R94 B.n241 B.n66 585
R95 B.n240 B.n239 585
R96 B.n238 B.n67 585
R97 B.n237 B.n236 585
R98 B.n235 B.n68 585
R99 B.n234 B.n233 585
R100 B.n232 B.n69 585
R101 B.n231 B.n230 585
R102 B.n229 B.n70 585
R103 B.n150 B.n149 585
R104 B.n151 B.n100 585
R105 B.n153 B.n152 585
R106 B.n154 B.n99 585
R107 B.n156 B.n155 585
R108 B.n157 B.n98 585
R109 B.n159 B.n158 585
R110 B.n160 B.n97 585
R111 B.n162 B.n161 585
R112 B.n163 B.n96 585
R113 B.n165 B.n164 585
R114 B.n166 B.n95 585
R115 B.n168 B.n167 585
R116 B.n169 B.n94 585
R117 B.n171 B.n170 585
R118 B.n172 B.n93 585
R119 B.n174 B.n173 585
R120 B.n175 B.n92 585
R121 B.n177 B.n176 585
R122 B.n178 B.n91 585
R123 B.n180 B.n179 585
R124 B.n182 B.n181 585
R125 B.n183 B.n87 585
R126 B.n185 B.n184 585
R127 B.n186 B.n86 585
R128 B.n188 B.n187 585
R129 B.n189 B.n85 585
R130 B.n191 B.n190 585
R131 B.n192 B.n84 585
R132 B.n194 B.n193 585
R133 B.n195 B.n81 585
R134 B.n198 B.n197 585
R135 B.n199 B.n80 585
R136 B.n201 B.n200 585
R137 B.n202 B.n79 585
R138 B.n204 B.n203 585
R139 B.n205 B.n78 585
R140 B.n207 B.n206 585
R141 B.n208 B.n77 585
R142 B.n210 B.n209 585
R143 B.n211 B.n76 585
R144 B.n213 B.n212 585
R145 B.n214 B.n75 585
R146 B.n216 B.n215 585
R147 B.n217 B.n74 585
R148 B.n219 B.n218 585
R149 B.n220 B.n73 585
R150 B.n222 B.n221 585
R151 B.n223 B.n72 585
R152 B.n225 B.n224 585
R153 B.n226 B.n71 585
R154 B.n228 B.n227 585
R155 B.n148 B.n101 585
R156 B.n147 B.n146 585
R157 B.n145 B.n102 585
R158 B.n144 B.n143 585
R159 B.n142 B.n103 585
R160 B.n141 B.n140 585
R161 B.n139 B.n104 585
R162 B.n138 B.n137 585
R163 B.n136 B.n105 585
R164 B.n135 B.n134 585
R165 B.n133 B.n106 585
R166 B.n132 B.n131 585
R167 B.n130 B.n107 585
R168 B.n129 B.n128 585
R169 B.n127 B.n108 585
R170 B.n126 B.n125 585
R171 B.n124 B.n109 585
R172 B.n123 B.n122 585
R173 B.n121 B.n110 585
R174 B.n120 B.n119 585
R175 B.n118 B.n111 585
R176 B.n117 B.n116 585
R177 B.n115 B.n112 585
R178 B.n114 B.n113 585
R179 B.n2 B.n0 585
R180 B.n421 B.n1 585
R181 B.n420 B.n419 585
R182 B.n418 B.n3 585
R183 B.n417 B.n416 585
R184 B.n415 B.n4 585
R185 B.n414 B.n413 585
R186 B.n412 B.n5 585
R187 B.n411 B.n410 585
R188 B.n409 B.n6 585
R189 B.n408 B.n407 585
R190 B.n406 B.n7 585
R191 B.n405 B.n404 585
R192 B.n403 B.n8 585
R193 B.n402 B.n401 585
R194 B.n400 B.n9 585
R195 B.n399 B.n398 585
R196 B.n397 B.n10 585
R197 B.n396 B.n395 585
R198 B.n394 B.n11 585
R199 B.n393 B.n392 585
R200 B.n391 B.n12 585
R201 B.n390 B.n389 585
R202 B.n388 B.n13 585
R203 B.n387 B.n386 585
R204 B.n385 B.n14 585
R205 B.n423 B.n422 585
R206 B.n150 B.n101 550.159
R207 B.n385 B.n384 550.159
R208 B.n229 B.n228 550.159
R209 B.n306 B.n45 550.159
R210 B.n82 B.t3 315.435
R211 B.n88 B.t6 315.435
R212 B.n26 B.t9 315.435
R213 B.n32 B.t0 315.435
R214 B.n82 B.t5 281.055
R215 B.n32 B.t1 281.055
R216 B.n88 B.t8 281.055
R217 B.n26 B.t10 281.055
R218 B.n83 B.t4 253.127
R219 B.n33 B.t2 253.127
R220 B.n89 B.t7 253.127
R221 B.n27 B.t11 253.127
R222 B.n146 B.n101 163.367
R223 B.n146 B.n145 163.367
R224 B.n145 B.n144 163.367
R225 B.n144 B.n103 163.367
R226 B.n140 B.n103 163.367
R227 B.n140 B.n139 163.367
R228 B.n139 B.n138 163.367
R229 B.n138 B.n105 163.367
R230 B.n134 B.n105 163.367
R231 B.n134 B.n133 163.367
R232 B.n133 B.n132 163.367
R233 B.n132 B.n107 163.367
R234 B.n128 B.n107 163.367
R235 B.n128 B.n127 163.367
R236 B.n127 B.n126 163.367
R237 B.n126 B.n109 163.367
R238 B.n122 B.n109 163.367
R239 B.n122 B.n121 163.367
R240 B.n121 B.n120 163.367
R241 B.n120 B.n111 163.367
R242 B.n116 B.n111 163.367
R243 B.n116 B.n115 163.367
R244 B.n115 B.n114 163.367
R245 B.n114 B.n2 163.367
R246 B.n422 B.n2 163.367
R247 B.n422 B.n421 163.367
R248 B.n421 B.n420 163.367
R249 B.n420 B.n3 163.367
R250 B.n416 B.n3 163.367
R251 B.n416 B.n415 163.367
R252 B.n415 B.n414 163.367
R253 B.n414 B.n5 163.367
R254 B.n410 B.n5 163.367
R255 B.n410 B.n409 163.367
R256 B.n409 B.n408 163.367
R257 B.n408 B.n7 163.367
R258 B.n404 B.n7 163.367
R259 B.n404 B.n403 163.367
R260 B.n403 B.n402 163.367
R261 B.n402 B.n9 163.367
R262 B.n398 B.n9 163.367
R263 B.n398 B.n397 163.367
R264 B.n397 B.n396 163.367
R265 B.n396 B.n11 163.367
R266 B.n392 B.n11 163.367
R267 B.n392 B.n391 163.367
R268 B.n391 B.n390 163.367
R269 B.n390 B.n13 163.367
R270 B.n386 B.n13 163.367
R271 B.n386 B.n385 163.367
R272 B.n151 B.n150 163.367
R273 B.n152 B.n151 163.367
R274 B.n152 B.n99 163.367
R275 B.n156 B.n99 163.367
R276 B.n157 B.n156 163.367
R277 B.n158 B.n157 163.367
R278 B.n158 B.n97 163.367
R279 B.n162 B.n97 163.367
R280 B.n163 B.n162 163.367
R281 B.n164 B.n163 163.367
R282 B.n164 B.n95 163.367
R283 B.n168 B.n95 163.367
R284 B.n169 B.n168 163.367
R285 B.n170 B.n169 163.367
R286 B.n170 B.n93 163.367
R287 B.n174 B.n93 163.367
R288 B.n175 B.n174 163.367
R289 B.n176 B.n175 163.367
R290 B.n176 B.n91 163.367
R291 B.n180 B.n91 163.367
R292 B.n181 B.n180 163.367
R293 B.n181 B.n87 163.367
R294 B.n185 B.n87 163.367
R295 B.n186 B.n185 163.367
R296 B.n187 B.n186 163.367
R297 B.n187 B.n85 163.367
R298 B.n191 B.n85 163.367
R299 B.n192 B.n191 163.367
R300 B.n193 B.n192 163.367
R301 B.n193 B.n81 163.367
R302 B.n198 B.n81 163.367
R303 B.n199 B.n198 163.367
R304 B.n200 B.n199 163.367
R305 B.n200 B.n79 163.367
R306 B.n204 B.n79 163.367
R307 B.n205 B.n204 163.367
R308 B.n206 B.n205 163.367
R309 B.n206 B.n77 163.367
R310 B.n210 B.n77 163.367
R311 B.n211 B.n210 163.367
R312 B.n212 B.n211 163.367
R313 B.n212 B.n75 163.367
R314 B.n216 B.n75 163.367
R315 B.n217 B.n216 163.367
R316 B.n218 B.n217 163.367
R317 B.n218 B.n73 163.367
R318 B.n222 B.n73 163.367
R319 B.n223 B.n222 163.367
R320 B.n224 B.n223 163.367
R321 B.n224 B.n71 163.367
R322 B.n228 B.n71 163.367
R323 B.n230 B.n229 163.367
R324 B.n230 B.n69 163.367
R325 B.n234 B.n69 163.367
R326 B.n235 B.n234 163.367
R327 B.n236 B.n235 163.367
R328 B.n236 B.n67 163.367
R329 B.n240 B.n67 163.367
R330 B.n241 B.n240 163.367
R331 B.n242 B.n241 163.367
R332 B.n242 B.n65 163.367
R333 B.n246 B.n65 163.367
R334 B.n247 B.n246 163.367
R335 B.n248 B.n247 163.367
R336 B.n248 B.n63 163.367
R337 B.n252 B.n63 163.367
R338 B.n253 B.n252 163.367
R339 B.n254 B.n253 163.367
R340 B.n254 B.n61 163.367
R341 B.n258 B.n61 163.367
R342 B.n259 B.n258 163.367
R343 B.n260 B.n259 163.367
R344 B.n260 B.n59 163.367
R345 B.n264 B.n59 163.367
R346 B.n265 B.n264 163.367
R347 B.n266 B.n265 163.367
R348 B.n266 B.n57 163.367
R349 B.n270 B.n57 163.367
R350 B.n271 B.n270 163.367
R351 B.n272 B.n271 163.367
R352 B.n272 B.n55 163.367
R353 B.n276 B.n55 163.367
R354 B.n277 B.n276 163.367
R355 B.n278 B.n277 163.367
R356 B.n278 B.n53 163.367
R357 B.n282 B.n53 163.367
R358 B.n283 B.n282 163.367
R359 B.n284 B.n283 163.367
R360 B.n284 B.n51 163.367
R361 B.n288 B.n51 163.367
R362 B.n289 B.n288 163.367
R363 B.n290 B.n289 163.367
R364 B.n290 B.n49 163.367
R365 B.n294 B.n49 163.367
R366 B.n295 B.n294 163.367
R367 B.n296 B.n295 163.367
R368 B.n296 B.n47 163.367
R369 B.n300 B.n47 163.367
R370 B.n301 B.n300 163.367
R371 B.n302 B.n301 163.367
R372 B.n302 B.n45 163.367
R373 B.n384 B.n15 163.367
R374 B.n380 B.n15 163.367
R375 B.n380 B.n379 163.367
R376 B.n379 B.n378 163.367
R377 B.n378 B.n17 163.367
R378 B.n374 B.n17 163.367
R379 B.n374 B.n373 163.367
R380 B.n373 B.n372 163.367
R381 B.n372 B.n19 163.367
R382 B.n368 B.n19 163.367
R383 B.n368 B.n367 163.367
R384 B.n367 B.n366 163.367
R385 B.n366 B.n21 163.367
R386 B.n362 B.n21 163.367
R387 B.n362 B.n361 163.367
R388 B.n361 B.n360 163.367
R389 B.n360 B.n23 163.367
R390 B.n356 B.n23 163.367
R391 B.n356 B.n355 163.367
R392 B.n355 B.n354 163.367
R393 B.n354 B.n25 163.367
R394 B.n349 B.n25 163.367
R395 B.n349 B.n348 163.367
R396 B.n348 B.n347 163.367
R397 B.n347 B.n29 163.367
R398 B.n343 B.n29 163.367
R399 B.n343 B.n342 163.367
R400 B.n342 B.n341 163.367
R401 B.n341 B.n31 163.367
R402 B.n337 B.n31 163.367
R403 B.n337 B.n336 163.367
R404 B.n336 B.n35 163.367
R405 B.n332 B.n35 163.367
R406 B.n332 B.n331 163.367
R407 B.n331 B.n330 163.367
R408 B.n330 B.n37 163.367
R409 B.n326 B.n37 163.367
R410 B.n326 B.n325 163.367
R411 B.n325 B.n324 163.367
R412 B.n324 B.n39 163.367
R413 B.n320 B.n39 163.367
R414 B.n320 B.n319 163.367
R415 B.n319 B.n318 163.367
R416 B.n318 B.n41 163.367
R417 B.n314 B.n41 163.367
R418 B.n314 B.n313 163.367
R419 B.n313 B.n312 163.367
R420 B.n312 B.n43 163.367
R421 B.n308 B.n43 163.367
R422 B.n308 B.n307 163.367
R423 B.n307 B.n306 163.367
R424 B.n196 B.n83 59.5399
R425 B.n90 B.n89 59.5399
R426 B.n352 B.n27 59.5399
R427 B.n34 B.n33 59.5399
R428 B.n383 B.n14 35.7468
R429 B.n305 B.n304 35.7468
R430 B.n227 B.n70 35.7468
R431 B.n149 B.n148 35.7468
R432 B.n83 B.n82 27.9278
R433 B.n89 B.n88 27.9278
R434 B.n27 B.n26 27.9278
R435 B.n33 B.n32 27.9278
R436 B B.n423 18.0485
R437 B.n383 B.n382 10.6151
R438 B.n382 B.n381 10.6151
R439 B.n381 B.n16 10.6151
R440 B.n377 B.n16 10.6151
R441 B.n377 B.n376 10.6151
R442 B.n376 B.n375 10.6151
R443 B.n375 B.n18 10.6151
R444 B.n371 B.n18 10.6151
R445 B.n371 B.n370 10.6151
R446 B.n370 B.n369 10.6151
R447 B.n369 B.n20 10.6151
R448 B.n365 B.n20 10.6151
R449 B.n365 B.n364 10.6151
R450 B.n364 B.n363 10.6151
R451 B.n363 B.n22 10.6151
R452 B.n359 B.n22 10.6151
R453 B.n359 B.n358 10.6151
R454 B.n358 B.n357 10.6151
R455 B.n357 B.n24 10.6151
R456 B.n353 B.n24 10.6151
R457 B.n351 B.n350 10.6151
R458 B.n350 B.n28 10.6151
R459 B.n346 B.n28 10.6151
R460 B.n346 B.n345 10.6151
R461 B.n345 B.n344 10.6151
R462 B.n344 B.n30 10.6151
R463 B.n340 B.n30 10.6151
R464 B.n340 B.n339 10.6151
R465 B.n339 B.n338 10.6151
R466 B.n335 B.n334 10.6151
R467 B.n334 B.n333 10.6151
R468 B.n333 B.n36 10.6151
R469 B.n329 B.n36 10.6151
R470 B.n329 B.n328 10.6151
R471 B.n328 B.n327 10.6151
R472 B.n327 B.n38 10.6151
R473 B.n323 B.n38 10.6151
R474 B.n323 B.n322 10.6151
R475 B.n322 B.n321 10.6151
R476 B.n321 B.n40 10.6151
R477 B.n317 B.n40 10.6151
R478 B.n317 B.n316 10.6151
R479 B.n316 B.n315 10.6151
R480 B.n315 B.n42 10.6151
R481 B.n311 B.n42 10.6151
R482 B.n311 B.n310 10.6151
R483 B.n310 B.n309 10.6151
R484 B.n309 B.n44 10.6151
R485 B.n305 B.n44 10.6151
R486 B.n231 B.n70 10.6151
R487 B.n232 B.n231 10.6151
R488 B.n233 B.n232 10.6151
R489 B.n233 B.n68 10.6151
R490 B.n237 B.n68 10.6151
R491 B.n238 B.n237 10.6151
R492 B.n239 B.n238 10.6151
R493 B.n239 B.n66 10.6151
R494 B.n243 B.n66 10.6151
R495 B.n244 B.n243 10.6151
R496 B.n245 B.n244 10.6151
R497 B.n245 B.n64 10.6151
R498 B.n249 B.n64 10.6151
R499 B.n250 B.n249 10.6151
R500 B.n251 B.n250 10.6151
R501 B.n251 B.n62 10.6151
R502 B.n255 B.n62 10.6151
R503 B.n256 B.n255 10.6151
R504 B.n257 B.n256 10.6151
R505 B.n257 B.n60 10.6151
R506 B.n261 B.n60 10.6151
R507 B.n262 B.n261 10.6151
R508 B.n263 B.n262 10.6151
R509 B.n263 B.n58 10.6151
R510 B.n267 B.n58 10.6151
R511 B.n268 B.n267 10.6151
R512 B.n269 B.n268 10.6151
R513 B.n269 B.n56 10.6151
R514 B.n273 B.n56 10.6151
R515 B.n274 B.n273 10.6151
R516 B.n275 B.n274 10.6151
R517 B.n275 B.n54 10.6151
R518 B.n279 B.n54 10.6151
R519 B.n280 B.n279 10.6151
R520 B.n281 B.n280 10.6151
R521 B.n281 B.n52 10.6151
R522 B.n285 B.n52 10.6151
R523 B.n286 B.n285 10.6151
R524 B.n287 B.n286 10.6151
R525 B.n287 B.n50 10.6151
R526 B.n291 B.n50 10.6151
R527 B.n292 B.n291 10.6151
R528 B.n293 B.n292 10.6151
R529 B.n293 B.n48 10.6151
R530 B.n297 B.n48 10.6151
R531 B.n298 B.n297 10.6151
R532 B.n299 B.n298 10.6151
R533 B.n299 B.n46 10.6151
R534 B.n303 B.n46 10.6151
R535 B.n304 B.n303 10.6151
R536 B.n149 B.n100 10.6151
R537 B.n153 B.n100 10.6151
R538 B.n154 B.n153 10.6151
R539 B.n155 B.n154 10.6151
R540 B.n155 B.n98 10.6151
R541 B.n159 B.n98 10.6151
R542 B.n160 B.n159 10.6151
R543 B.n161 B.n160 10.6151
R544 B.n161 B.n96 10.6151
R545 B.n165 B.n96 10.6151
R546 B.n166 B.n165 10.6151
R547 B.n167 B.n166 10.6151
R548 B.n167 B.n94 10.6151
R549 B.n171 B.n94 10.6151
R550 B.n172 B.n171 10.6151
R551 B.n173 B.n172 10.6151
R552 B.n173 B.n92 10.6151
R553 B.n177 B.n92 10.6151
R554 B.n178 B.n177 10.6151
R555 B.n179 B.n178 10.6151
R556 B.n183 B.n182 10.6151
R557 B.n184 B.n183 10.6151
R558 B.n184 B.n86 10.6151
R559 B.n188 B.n86 10.6151
R560 B.n189 B.n188 10.6151
R561 B.n190 B.n189 10.6151
R562 B.n190 B.n84 10.6151
R563 B.n194 B.n84 10.6151
R564 B.n195 B.n194 10.6151
R565 B.n197 B.n80 10.6151
R566 B.n201 B.n80 10.6151
R567 B.n202 B.n201 10.6151
R568 B.n203 B.n202 10.6151
R569 B.n203 B.n78 10.6151
R570 B.n207 B.n78 10.6151
R571 B.n208 B.n207 10.6151
R572 B.n209 B.n208 10.6151
R573 B.n209 B.n76 10.6151
R574 B.n213 B.n76 10.6151
R575 B.n214 B.n213 10.6151
R576 B.n215 B.n214 10.6151
R577 B.n215 B.n74 10.6151
R578 B.n219 B.n74 10.6151
R579 B.n220 B.n219 10.6151
R580 B.n221 B.n220 10.6151
R581 B.n221 B.n72 10.6151
R582 B.n225 B.n72 10.6151
R583 B.n226 B.n225 10.6151
R584 B.n227 B.n226 10.6151
R585 B.n148 B.n147 10.6151
R586 B.n147 B.n102 10.6151
R587 B.n143 B.n102 10.6151
R588 B.n143 B.n142 10.6151
R589 B.n142 B.n141 10.6151
R590 B.n141 B.n104 10.6151
R591 B.n137 B.n104 10.6151
R592 B.n137 B.n136 10.6151
R593 B.n136 B.n135 10.6151
R594 B.n135 B.n106 10.6151
R595 B.n131 B.n106 10.6151
R596 B.n131 B.n130 10.6151
R597 B.n130 B.n129 10.6151
R598 B.n129 B.n108 10.6151
R599 B.n125 B.n108 10.6151
R600 B.n125 B.n124 10.6151
R601 B.n124 B.n123 10.6151
R602 B.n123 B.n110 10.6151
R603 B.n119 B.n110 10.6151
R604 B.n119 B.n118 10.6151
R605 B.n118 B.n117 10.6151
R606 B.n117 B.n112 10.6151
R607 B.n113 B.n112 10.6151
R608 B.n113 B.n0 10.6151
R609 B.n419 B.n1 10.6151
R610 B.n419 B.n418 10.6151
R611 B.n418 B.n417 10.6151
R612 B.n417 B.n4 10.6151
R613 B.n413 B.n4 10.6151
R614 B.n413 B.n412 10.6151
R615 B.n412 B.n411 10.6151
R616 B.n411 B.n6 10.6151
R617 B.n407 B.n6 10.6151
R618 B.n407 B.n406 10.6151
R619 B.n406 B.n405 10.6151
R620 B.n405 B.n8 10.6151
R621 B.n401 B.n8 10.6151
R622 B.n401 B.n400 10.6151
R623 B.n400 B.n399 10.6151
R624 B.n399 B.n10 10.6151
R625 B.n395 B.n10 10.6151
R626 B.n395 B.n394 10.6151
R627 B.n394 B.n393 10.6151
R628 B.n393 B.n12 10.6151
R629 B.n389 B.n12 10.6151
R630 B.n389 B.n388 10.6151
R631 B.n388 B.n387 10.6151
R632 B.n387 B.n14 10.6151
R633 B.n353 B.n352 9.36635
R634 B.n335 B.n34 9.36635
R635 B.n179 B.n90 9.36635
R636 B.n197 B.n196 9.36635
R637 B.n423 B.n0 2.81026
R638 B.n423 B.n1 2.81026
R639 B.n352 B.n351 1.24928
R640 B.n338 B.n34 1.24928
R641 B.n182 B.n90 1.24928
R642 B.n196 B.n195 1.24928
R643 VP.n3 VP.t3 170.547
R644 VP.n5 VP.n2 161.3
R645 VP.n13 VP.n0 161.3
R646 VP.n12 VP.n11 161.3
R647 VP.n10 VP.n1 161.3
R648 VP.n8 VP.t0 147.423
R649 VP.n14 VP.t5 147.423
R650 VP.n6 VP.t4 147.423
R651 VP.n12 VP.t1 111.816
R652 VP.n4 VP.t2 111.816
R653 VP.n7 VP.n6 80.6037
R654 VP.n15 VP.n14 80.6037
R655 VP.n9 VP.n8 80.6037
R656 VP.n8 VP.n1 50.8919
R657 VP.n14 VP.n13 50.8919
R658 VP.n6 VP.n5 50.8919
R659 VP.n9 VP.n7 37.8423
R660 VP.n4 VP.n3 32.7474
R661 VP.n3 VP.n2 28.089
R662 VP.n12 VP.n1 24.4675
R663 VP.n13 VP.n12 24.4675
R664 VP.n5 VP.n4 24.4675
R665 VP.n7 VP.n2 0.285035
R666 VP.n10 VP.n9 0.285035
R667 VP.n15 VP.n0 0.285035
R668 VP.n11 VP.n10 0.189894
R669 VP.n11 VP.n0 0.189894
R670 VP VP.n15 0.146778
R671 VTAIL.n110 VTAIL.n109 756.745
R672 VTAIL.n26 VTAIL.n25 756.745
R673 VTAIL.n84 VTAIL.n83 756.745
R674 VTAIL.n56 VTAIL.n55 756.745
R675 VTAIL.n95 VTAIL.n94 585
R676 VTAIL.n92 VTAIL.n91 585
R677 VTAIL.n101 VTAIL.n100 585
R678 VTAIL.n103 VTAIL.n102 585
R679 VTAIL.n88 VTAIL.n87 585
R680 VTAIL.n109 VTAIL.n108 585
R681 VTAIL.n11 VTAIL.n10 585
R682 VTAIL.n8 VTAIL.n7 585
R683 VTAIL.n17 VTAIL.n16 585
R684 VTAIL.n19 VTAIL.n18 585
R685 VTAIL.n4 VTAIL.n3 585
R686 VTAIL.n25 VTAIL.n24 585
R687 VTAIL.n83 VTAIL.n82 585
R688 VTAIL.n62 VTAIL.n61 585
R689 VTAIL.n77 VTAIL.n76 585
R690 VTAIL.n75 VTAIL.n74 585
R691 VTAIL.n66 VTAIL.n65 585
R692 VTAIL.n69 VTAIL.n68 585
R693 VTAIL.n55 VTAIL.n54 585
R694 VTAIL.n34 VTAIL.n33 585
R695 VTAIL.n49 VTAIL.n48 585
R696 VTAIL.n47 VTAIL.n46 585
R697 VTAIL.n38 VTAIL.n37 585
R698 VTAIL.n41 VTAIL.n40 585
R699 VTAIL.t11 VTAIL.n67 329.435
R700 VTAIL.t2 VTAIL.n93 329.435
R701 VTAIL.t10 VTAIL.n9 329.435
R702 VTAIL.t4 VTAIL.n39 329.435
R703 VTAIL.n94 VTAIL.n91 171.744
R704 VTAIL.n101 VTAIL.n91 171.744
R705 VTAIL.n102 VTAIL.n101 171.744
R706 VTAIL.n102 VTAIL.n87 171.744
R707 VTAIL.n109 VTAIL.n87 171.744
R708 VTAIL.n10 VTAIL.n7 171.744
R709 VTAIL.n17 VTAIL.n7 171.744
R710 VTAIL.n18 VTAIL.n17 171.744
R711 VTAIL.n18 VTAIL.n3 171.744
R712 VTAIL.n25 VTAIL.n3 171.744
R713 VTAIL.n83 VTAIL.n61 171.744
R714 VTAIL.n76 VTAIL.n61 171.744
R715 VTAIL.n76 VTAIL.n75 171.744
R716 VTAIL.n75 VTAIL.n65 171.744
R717 VTAIL.n68 VTAIL.n65 171.744
R718 VTAIL.n55 VTAIL.n33 171.744
R719 VTAIL.n48 VTAIL.n33 171.744
R720 VTAIL.n48 VTAIL.n47 171.744
R721 VTAIL.n47 VTAIL.n37 171.744
R722 VTAIL.n40 VTAIL.n37 171.744
R723 VTAIL.n94 VTAIL.t2 85.8723
R724 VTAIL.n10 VTAIL.t10 85.8723
R725 VTAIL.n68 VTAIL.t11 85.8723
R726 VTAIL.n40 VTAIL.t4 85.8723
R727 VTAIL.n59 VTAIL.n58 84.2808
R728 VTAIL.n31 VTAIL.n30 84.2808
R729 VTAIL.n1 VTAIL.n0 84.2807
R730 VTAIL.n29 VTAIL.n28 84.2807
R731 VTAIL.n111 VTAIL.n110 34.7066
R732 VTAIL.n27 VTAIL.n26 34.7066
R733 VTAIL.n85 VTAIL.n84 34.7066
R734 VTAIL.n57 VTAIL.n56 34.7066
R735 VTAIL.n31 VTAIL.n29 19.2893
R736 VTAIL.n111 VTAIL.n85 18.0479
R737 VTAIL.n108 VTAIL.n86 11.249
R738 VTAIL.n24 VTAIL.n2 11.249
R739 VTAIL.n82 VTAIL.n60 11.249
R740 VTAIL.n54 VTAIL.n32 11.249
R741 VTAIL.n95 VTAIL.n93 10.7185
R742 VTAIL.n11 VTAIL.n9 10.7185
R743 VTAIL.n69 VTAIL.n67 10.7185
R744 VTAIL.n41 VTAIL.n39 10.7185
R745 VTAIL.n107 VTAIL.n88 10.4732
R746 VTAIL.n23 VTAIL.n4 10.4732
R747 VTAIL.n81 VTAIL.n62 10.4732
R748 VTAIL.n53 VTAIL.n34 10.4732
R749 VTAIL.n104 VTAIL.n103 9.69747
R750 VTAIL.n20 VTAIL.n19 9.69747
R751 VTAIL.n78 VTAIL.n77 9.69747
R752 VTAIL.n50 VTAIL.n49 9.69747
R753 VTAIL.n106 VTAIL.n86 9.45567
R754 VTAIL.n22 VTAIL.n2 9.45567
R755 VTAIL.n80 VTAIL.n60 9.45567
R756 VTAIL.n52 VTAIL.n32 9.45567
R757 VTAIL.n97 VTAIL.n96 9.3005
R758 VTAIL.n99 VTAIL.n98 9.3005
R759 VTAIL.n90 VTAIL.n89 9.3005
R760 VTAIL.n105 VTAIL.n104 9.3005
R761 VTAIL.n107 VTAIL.n106 9.3005
R762 VTAIL.n13 VTAIL.n12 9.3005
R763 VTAIL.n15 VTAIL.n14 9.3005
R764 VTAIL.n6 VTAIL.n5 9.3005
R765 VTAIL.n21 VTAIL.n20 9.3005
R766 VTAIL.n23 VTAIL.n22 9.3005
R767 VTAIL.n81 VTAIL.n80 9.3005
R768 VTAIL.n79 VTAIL.n78 9.3005
R769 VTAIL.n64 VTAIL.n63 9.3005
R770 VTAIL.n73 VTAIL.n72 9.3005
R771 VTAIL.n71 VTAIL.n70 9.3005
R772 VTAIL.n45 VTAIL.n44 9.3005
R773 VTAIL.n36 VTAIL.n35 9.3005
R774 VTAIL.n51 VTAIL.n50 9.3005
R775 VTAIL.n53 VTAIL.n52 9.3005
R776 VTAIL.n43 VTAIL.n42 9.3005
R777 VTAIL.n100 VTAIL.n90 8.92171
R778 VTAIL.n16 VTAIL.n6 8.92171
R779 VTAIL.n74 VTAIL.n64 8.92171
R780 VTAIL.n46 VTAIL.n36 8.92171
R781 VTAIL.n99 VTAIL.n92 8.14595
R782 VTAIL.n15 VTAIL.n8 8.14595
R783 VTAIL.n73 VTAIL.n66 8.14595
R784 VTAIL.n45 VTAIL.n38 8.14595
R785 VTAIL.n96 VTAIL.n95 7.3702
R786 VTAIL.n12 VTAIL.n11 7.3702
R787 VTAIL.n70 VTAIL.n69 7.3702
R788 VTAIL.n42 VTAIL.n41 7.3702
R789 VTAIL.n0 VTAIL.t0 6.31215
R790 VTAIL.n0 VTAIL.t3 6.31215
R791 VTAIL.n28 VTAIL.t9 6.31215
R792 VTAIL.n28 VTAIL.t7 6.31215
R793 VTAIL.n58 VTAIL.t8 6.31215
R794 VTAIL.n58 VTAIL.t6 6.31215
R795 VTAIL.n30 VTAIL.t5 6.31215
R796 VTAIL.n30 VTAIL.t1 6.31215
R797 VTAIL.n96 VTAIL.n92 5.81868
R798 VTAIL.n12 VTAIL.n8 5.81868
R799 VTAIL.n70 VTAIL.n66 5.81868
R800 VTAIL.n42 VTAIL.n38 5.81868
R801 VTAIL.n100 VTAIL.n99 5.04292
R802 VTAIL.n16 VTAIL.n15 5.04292
R803 VTAIL.n74 VTAIL.n73 5.04292
R804 VTAIL.n46 VTAIL.n45 5.04292
R805 VTAIL.n103 VTAIL.n90 4.26717
R806 VTAIL.n19 VTAIL.n6 4.26717
R807 VTAIL.n77 VTAIL.n64 4.26717
R808 VTAIL.n49 VTAIL.n36 4.26717
R809 VTAIL.n104 VTAIL.n88 3.49141
R810 VTAIL.n20 VTAIL.n4 3.49141
R811 VTAIL.n78 VTAIL.n62 3.49141
R812 VTAIL.n50 VTAIL.n34 3.49141
R813 VTAIL.n108 VTAIL.n107 2.71565
R814 VTAIL.n24 VTAIL.n23 2.71565
R815 VTAIL.n82 VTAIL.n81 2.71565
R816 VTAIL.n54 VTAIL.n53 2.71565
R817 VTAIL.n97 VTAIL.n93 2.41827
R818 VTAIL.n13 VTAIL.n9 2.41827
R819 VTAIL.n71 VTAIL.n67 2.41827
R820 VTAIL.n43 VTAIL.n39 2.41827
R821 VTAIL.n110 VTAIL.n86 1.93989
R822 VTAIL.n26 VTAIL.n2 1.93989
R823 VTAIL.n84 VTAIL.n60 1.93989
R824 VTAIL.n56 VTAIL.n32 1.93989
R825 VTAIL.n57 VTAIL.n31 1.24188
R826 VTAIL.n85 VTAIL.n59 1.24188
R827 VTAIL.n29 VTAIL.n27 1.24188
R828 VTAIL.n59 VTAIL.n57 1.09102
R829 VTAIL.n27 VTAIL.n1 1.09102
R830 VTAIL VTAIL.n111 0.873345
R831 VTAIL VTAIL.n1 0.369034
R832 VTAIL.n98 VTAIL.n97 0.155672
R833 VTAIL.n98 VTAIL.n89 0.155672
R834 VTAIL.n105 VTAIL.n89 0.155672
R835 VTAIL.n106 VTAIL.n105 0.155672
R836 VTAIL.n14 VTAIL.n13 0.155672
R837 VTAIL.n14 VTAIL.n5 0.155672
R838 VTAIL.n21 VTAIL.n5 0.155672
R839 VTAIL.n22 VTAIL.n21 0.155672
R840 VTAIL.n80 VTAIL.n79 0.155672
R841 VTAIL.n79 VTAIL.n63 0.155672
R842 VTAIL.n72 VTAIL.n63 0.155672
R843 VTAIL.n72 VTAIL.n71 0.155672
R844 VTAIL.n52 VTAIL.n51 0.155672
R845 VTAIL.n51 VTAIL.n35 0.155672
R846 VTAIL.n44 VTAIL.n35 0.155672
R847 VTAIL.n44 VTAIL.n43 0.155672
R848 VDD1.n24 VDD1.n23 756.745
R849 VDD1.n49 VDD1.n48 756.745
R850 VDD1.n23 VDD1.n22 585
R851 VDD1.n2 VDD1.n1 585
R852 VDD1.n17 VDD1.n16 585
R853 VDD1.n15 VDD1.n14 585
R854 VDD1.n6 VDD1.n5 585
R855 VDD1.n9 VDD1.n8 585
R856 VDD1.n34 VDD1.n33 585
R857 VDD1.n31 VDD1.n30 585
R858 VDD1.n40 VDD1.n39 585
R859 VDD1.n42 VDD1.n41 585
R860 VDD1.n27 VDD1.n26 585
R861 VDD1.n48 VDD1.n47 585
R862 VDD1.t2 VDD1.n7 329.435
R863 VDD1.t5 VDD1.n32 329.435
R864 VDD1.n23 VDD1.n1 171.744
R865 VDD1.n16 VDD1.n1 171.744
R866 VDD1.n16 VDD1.n15 171.744
R867 VDD1.n15 VDD1.n5 171.744
R868 VDD1.n8 VDD1.n5 171.744
R869 VDD1.n33 VDD1.n30 171.744
R870 VDD1.n40 VDD1.n30 171.744
R871 VDD1.n41 VDD1.n40 171.744
R872 VDD1.n41 VDD1.n26 171.744
R873 VDD1.n48 VDD1.n26 171.744
R874 VDD1.n51 VDD1.n50 101.215
R875 VDD1.n53 VDD1.n52 100.959
R876 VDD1.n8 VDD1.t2 85.8723
R877 VDD1.n33 VDD1.t5 85.8723
R878 VDD1 VDD1.n24 52.3746
R879 VDD1.n51 VDD1.n49 52.261
R880 VDD1.n53 VDD1.n51 33.3931
R881 VDD1.n22 VDD1.n0 11.249
R882 VDD1.n47 VDD1.n25 11.249
R883 VDD1.n9 VDD1.n7 10.7185
R884 VDD1.n34 VDD1.n32 10.7185
R885 VDD1.n21 VDD1.n2 10.4732
R886 VDD1.n46 VDD1.n27 10.4732
R887 VDD1.n18 VDD1.n17 9.69747
R888 VDD1.n43 VDD1.n42 9.69747
R889 VDD1.n20 VDD1.n0 9.45567
R890 VDD1.n45 VDD1.n25 9.45567
R891 VDD1.n13 VDD1.n12 9.3005
R892 VDD1.n4 VDD1.n3 9.3005
R893 VDD1.n19 VDD1.n18 9.3005
R894 VDD1.n21 VDD1.n20 9.3005
R895 VDD1.n11 VDD1.n10 9.3005
R896 VDD1.n36 VDD1.n35 9.3005
R897 VDD1.n38 VDD1.n37 9.3005
R898 VDD1.n29 VDD1.n28 9.3005
R899 VDD1.n44 VDD1.n43 9.3005
R900 VDD1.n46 VDD1.n45 9.3005
R901 VDD1.n14 VDD1.n4 8.92171
R902 VDD1.n39 VDD1.n29 8.92171
R903 VDD1.n13 VDD1.n6 8.14595
R904 VDD1.n38 VDD1.n31 8.14595
R905 VDD1.n10 VDD1.n9 7.3702
R906 VDD1.n35 VDD1.n34 7.3702
R907 VDD1.n52 VDD1.t3 6.31215
R908 VDD1.n52 VDD1.t1 6.31215
R909 VDD1.n50 VDD1.t4 6.31215
R910 VDD1.n50 VDD1.t0 6.31215
R911 VDD1.n10 VDD1.n6 5.81868
R912 VDD1.n35 VDD1.n31 5.81868
R913 VDD1.n14 VDD1.n13 5.04292
R914 VDD1.n39 VDD1.n38 5.04292
R915 VDD1.n17 VDD1.n4 4.26717
R916 VDD1.n42 VDD1.n29 4.26717
R917 VDD1.n18 VDD1.n2 3.49141
R918 VDD1.n43 VDD1.n27 3.49141
R919 VDD1.n22 VDD1.n21 2.71565
R920 VDD1.n47 VDD1.n46 2.71565
R921 VDD1.n11 VDD1.n7 2.41827
R922 VDD1.n36 VDD1.n32 2.41827
R923 VDD1.n24 VDD1.n0 1.93989
R924 VDD1.n49 VDD1.n25 1.93989
R925 VDD1 VDD1.n53 0.252655
R926 VDD1.n20 VDD1.n19 0.155672
R927 VDD1.n19 VDD1.n3 0.155672
R928 VDD1.n12 VDD1.n3 0.155672
R929 VDD1.n12 VDD1.n11 0.155672
R930 VDD1.n37 VDD1.n36 0.155672
R931 VDD1.n37 VDD1.n28 0.155672
R932 VDD1.n44 VDD1.n28 0.155672
R933 VDD1.n45 VDD1.n44 0.155672
R934 VN.n1 VN.t5 170.547
R935 VN.n7 VN.t2 170.547
R936 VN.n9 VN.n6 161.3
R937 VN.n3 VN.n0 161.3
R938 VN.n4 VN.t0 147.423
R939 VN.n10 VN.t4 147.423
R940 VN.n2 VN.t1 111.816
R941 VN.n8 VN.t3 111.816
R942 VN.n11 VN.n10 80.6037
R943 VN.n5 VN.n4 80.6037
R944 VN.n4 VN.n3 50.8919
R945 VN.n10 VN.n9 50.8919
R946 VN VN.n11 38.1278
R947 VN.n2 VN.n1 32.7474
R948 VN.n8 VN.n7 32.7474
R949 VN.n7 VN.n6 28.089
R950 VN.n1 VN.n0 28.089
R951 VN.n3 VN.n2 24.4675
R952 VN.n9 VN.n8 24.4675
R953 VN.n11 VN.n6 0.285035
R954 VN.n5 VN.n0 0.285035
R955 VN VN.n5 0.146778
R956 VDD2.n51 VDD2.n50 756.745
R957 VDD2.n24 VDD2.n23 756.745
R958 VDD2.n50 VDD2.n49 585
R959 VDD2.n29 VDD2.n28 585
R960 VDD2.n44 VDD2.n43 585
R961 VDD2.n42 VDD2.n41 585
R962 VDD2.n33 VDD2.n32 585
R963 VDD2.n36 VDD2.n35 585
R964 VDD2.n9 VDD2.n8 585
R965 VDD2.n6 VDD2.n5 585
R966 VDD2.n15 VDD2.n14 585
R967 VDD2.n17 VDD2.n16 585
R968 VDD2.n2 VDD2.n1 585
R969 VDD2.n23 VDD2.n22 585
R970 VDD2.t1 VDD2.n34 329.435
R971 VDD2.t0 VDD2.n7 329.435
R972 VDD2.n50 VDD2.n28 171.744
R973 VDD2.n43 VDD2.n28 171.744
R974 VDD2.n43 VDD2.n42 171.744
R975 VDD2.n42 VDD2.n32 171.744
R976 VDD2.n35 VDD2.n32 171.744
R977 VDD2.n8 VDD2.n5 171.744
R978 VDD2.n15 VDD2.n5 171.744
R979 VDD2.n16 VDD2.n15 171.744
R980 VDD2.n16 VDD2.n1 171.744
R981 VDD2.n23 VDD2.n1 171.744
R982 VDD2.n26 VDD2.n25 101.215
R983 VDD2 VDD2.n53 101.21
R984 VDD2.n35 VDD2.t1 85.8723
R985 VDD2.n8 VDD2.t0 85.8723
R986 VDD2.n26 VDD2.n24 52.261
R987 VDD2.n52 VDD2.n51 51.3853
R988 VDD2.n52 VDD2.n26 32.1894
R989 VDD2.n49 VDD2.n27 11.249
R990 VDD2.n22 VDD2.n0 11.249
R991 VDD2.n36 VDD2.n34 10.7185
R992 VDD2.n9 VDD2.n7 10.7185
R993 VDD2.n48 VDD2.n29 10.4732
R994 VDD2.n21 VDD2.n2 10.4732
R995 VDD2.n45 VDD2.n44 9.69747
R996 VDD2.n18 VDD2.n17 9.69747
R997 VDD2.n47 VDD2.n27 9.45567
R998 VDD2.n20 VDD2.n0 9.45567
R999 VDD2.n40 VDD2.n39 9.3005
R1000 VDD2.n31 VDD2.n30 9.3005
R1001 VDD2.n46 VDD2.n45 9.3005
R1002 VDD2.n48 VDD2.n47 9.3005
R1003 VDD2.n38 VDD2.n37 9.3005
R1004 VDD2.n11 VDD2.n10 9.3005
R1005 VDD2.n13 VDD2.n12 9.3005
R1006 VDD2.n4 VDD2.n3 9.3005
R1007 VDD2.n19 VDD2.n18 9.3005
R1008 VDD2.n21 VDD2.n20 9.3005
R1009 VDD2.n41 VDD2.n31 8.92171
R1010 VDD2.n14 VDD2.n4 8.92171
R1011 VDD2.n40 VDD2.n33 8.14595
R1012 VDD2.n13 VDD2.n6 8.14595
R1013 VDD2.n37 VDD2.n36 7.3702
R1014 VDD2.n10 VDD2.n9 7.3702
R1015 VDD2.n53 VDD2.t2 6.31215
R1016 VDD2.n53 VDD2.t3 6.31215
R1017 VDD2.n25 VDD2.t4 6.31215
R1018 VDD2.n25 VDD2.t5 6.31215
R1019 VDD2.n37 VDD2.n33 5.81868
R1020 VDD2.n10 VDD2.n6 5.81868
R1021 VDD2.n41 VDD2.n40 5.04292
R1022 VDD2.n14 VDD2.n13 5.04292
R1023 VDD2.n44 VDD2.n31 4.26717
R1024 VDD2.n17 VDD2.n4 4.26717
R1025 VDD2.n45 VDD2.n29 3.49141
R1026 VDD2.n18 VDD2.n2 3.49141
R1027 VDD2.n49 VDD2.n48 2.71565
R1028 VDD2.n22 VDD2.n21 2.71565
R1029 VDD2.n38 VDD2.n34 2.41827
R1030 VDD2.n11 VDD2.n7 2.41827
R1031 VDD2.n51 VDD2.n27 1.93989
R1032 VDD2.n24 VDD2.n0 1.93989
R1033 VDD2 VDD2.n52 0.989724
R1034 VDD2.n47 VDD2.n46 0.155672
R1035 VDD2.n46 VDD2.n30 0.155672
R1036 VDD2.n39 VDD2.n30 0.155672
R1037 VDD2.n39 VDD2.n38 0.155672
R1038 VDD2.n12 VDD2.n11 0.155672
R1039 VDD2.n12 VDD2.n3 0.155672
R1040 VDD2.n19 VDD2.n3 0.155672
R1041 VDD2.n20 VDD2.n19 0.155672
C0 VN B 0.779332f
C1 VDD1 B 1.1706f
C2 VDD2 B 1.2093f
C3 B VP 1.22291f
C4 VDD1 VN 0.148764f
C5 VDD2 VN 2.47509f
C6 VN VP 4.20838f
C7 VDD2 VDD1 0.860047f
C8 VDD1 VP 2.65566f
C9 w_n2122_n1998# VTAIL 1.86758f
C10 VDD2 VP 0.335424f
C11 B VTAIL 1.64364f
C12 w_n2122_n1998# B 5.70219f
C13 VN VTAIL 2.63347f
C14 VDD1 VTAIL 4.91841f
C15 VDD2 VTAIL 4.95966f
C16 VTAIL VP 2.64774f
C17 w_n2122_n1998# VN 3.52293f
C18 VDD1 w_n2122_n1998# 1.42469f
C19 VDD2 w_n2122_n1998# 1.46146f
C20 w_n2122_n1998# VP 3.79304f
C21 VDD2 VSUBS 1.062168f
C22 VDD1 VSUBS 1.038218f
C23 VTAIL VSUBS 0.46178f
C24 VN VSUBS 4.20063f
C25 VP VSUBS 1.45101f
C26 B VSUBS 2.464779f
C27 w_n2122_n1998# VSUBS 53.0924f
C28 VDD2.n0 VSUBS 0.012789f
C29 VDD2.n1 VSUBS 0.028776f
C30 VDD2.n2 VSUBS 0.01289f
C31 VDD2.n3 VSUBS 0.022656f
C32 VDD2.n4 VSUBS 0.012174f
C33 VDD2.n5 VSUBS 0.028776f
C34 VDD2.n6 VSUBS 0.01289f
C35 VDD2.n7 VSUBS 0.108853f
C36 VDD2.t0 VSUBS 0.06224f
C37 VDD2.n8 VSUBS 0.021582f
C38 VDD2.n9 VSUBS 0.02162f
C39 VDD2.n10 VSUBS 0.012174f
C40 VDD2.n11 VSUBS 0.431831f
C41 VDD2.n12 VSUBS 0.022656f
C42 VDD2.n13 VSUBS 0.012174f
C43 VDD2.n14 VSUBS 0.01289f
C44 VDD2.n15 VSUBS 0.028776f
C45 VDD2.n16 VSUBS 0.028776f
C46 VDD2.n17 VSUBS 0.01289f
C47 VDD2.n18 VSUBS 0.012174f
C48 VDD2.n19 VSUBS 0.022656f
C49 VDD2.n20 VSUBS 0.059486f
C50 VDD2.n21 VSUBS 0.012174f
C51 VDD2.n22 VSUBS 0.01289f
C52 VDD2.n23 VSUBS 0.063779f
C53 VDD2.n24 VSUBS 0.060901f
C54 VDD2.t4 VSUBS 0.092202f
C55 VDD2.t5 VSUBS 0.092202f
C56 VDD2.n25 VSUBS 0.601162f
C57 VDD2.n26 VSUBS 1.62291f
C58 VDD2.n27 VSUBS 0.012789f
C59 VDD2.n28 VSUBS 0.028776f
C60 VDD2.n29 VSUBS 0.01289f
C61 VDD2.n30 VSUBS 0.022656f
C62 VDD2.n31 VSUBS 0.012174f
C63 VDD2.n32 VSUBS 0.028776f
C64 VDD2.n33 VSUBS 0.01289f
C65 VDD2.n34 VSUBS 0.108853f
C66 VDD2.t1 VSUBS 0.06224f
C67 VDD2.n35 VSUBS 0.021582f
C68 VDD2.n36 VSUBS 0.02162f
C69 VDD2.n37 VSUBS 0.012174f
C70 VDD2.n38 VSUBS 0.431831f
C71 VDD2.n39 VSUBS 0.022656f
C72 VDD2.n40 VSUBS 0.012174f
C73 VDD2.n41 VSUBS 0.01289f
C74 VDD2.n42 VSUBS 0.028776f
C75 VDD2.n43 VSUBS 0.028776f
C76 VDD2.n44 VSUBS 0.01289f
C77 VDD2.n45 VSUBS 0.012174f
C78 VDD2.n46 VSUBS 0.022656f
C79 VDD2.n47 VSUBS 0.059486f
C80 VDD2.n48 VSUBS 0.012174f
C81 VDD2.n49 VSUBS 0.01289f
C82 VDD2.n50 VSUBS 0.063779f
C83 VDD2.n51 VSUBS 0.05905f
C84 VDD2.n52 VSUBS 1.46228f
C85 VDD2.t2 VSUBS 0.092202f
C86 VDD2.t3 VSUBS 0.092202f
C87 VDD2.n53 VSUBS 0.601143f
C88 VN.n0 VSUBS 0.308666f
C89 VN.t1 VSUBS 0.82783f
C90 VN.t5 VSUBS 0.983569f
C91 VN.n1 VSUBS 0.416839f
C92 VN.n2 VSUBS 0.43733f
C93 VN.n3 VSUBS 0.073664f
C94 VN.t0 VSUBS 0.921785f
C95 VN.n4 VSUBS 0.441529f
C96 VN.n5 VSUBS 0.051744f
C97 VN.n6 VSUBS 0.308666f
C98 VN.t3 VSUBS 0.82783f
C99 VN.t2 VSUBS 0.983569f
C100 VN.n7 VSUBS 0.416839f
C101 VN.n8 VSUBS 0.43733f
C102 VN.n9 VSUBS 0.073664f
C103 VN.t4 VSUBS 0.921785f
C104 VN.n10 VSUBS 0.441529f
C105 VN.n11 VSUBS 1.95531f
C106 VDD1.n0 VSUBS 0.012816f
C107 VDD1.n1 VSUBS 0.028837f
C108 VDD1.n2 VSUBS 0.012918f
C109 VDD1.n3 VSUBS 0.022705f
C110 VDD1.n4 VSUBS 0.0122f
C111 VDD1.n5 VSUBS 0.028837f
C112 VDD1.n6 VSUBS 0.012918f
C113 VDD1.n7 VSUBS 0.109088f
C114 VDD1.t2 VSUBS 0.062374f
C115 VDD1.n8 VSUBS 0.021628f
C116 VDD1.n9 VSUBS 0.021667f
C117 VDD1.n10 VSUBS 0.0122f
C118 VDD1.n11 VSUBS 0.43276f
C119 VDD1.n12 VSUBS 0.022705f
C120 VDD1.n13 VSUBS 0.0122f
C121 VDD1.n14 VSUBS 0.012918f
C122 VDD1.n15 VSUBS 0.028837f
C123 VDD1.n16 VSUBS 0.028837f
C124 VDD1.n17 VSUBS 0.012918f
C125 VDD1.n18 VSUBS 0.0122f
C126 VDD1.n19 VSUBS 0.022705f
C127 VDD1.n20 VSUBS 0.059614f
C128 VDD1.n21 VSUBS 0.0122f
C129 VDD1.n22 VSUBS 0.012918f
C130 VDD1.n23 VSUBS 0.063916f
C131 VDD1.n24 VSUBS 0.061413f
C132 VDD1.n25 VSUBS 0.012816f
C133 VDD1.n26 VSUBS 0.028837f
C134 VDD1.n27 VSUBS 0.012918f
C135 VDD1.n28 VSUBS 0.022705f
C136 VDD1.n29 VSUBS 0.0122f
C137 VDD1.n30 VSUBS 0.028837f
C138 VDD1.n31 VSUBS 0.012918f
C139 VDD1.n32 VSUBS 0.109088f
C140 VDD1.t5 VSUBS 0.062374f
C141 VDD1.n33 VSUBS 0.021628f
C142 VDD1.n34 VSUBS 0.021667f
C143 VDD1.n35 VSUBS 0.0122f
C144 VDD1.n36 VSUBS 0.43276f
C145 VDD1.n37 VSUBS 0.022705f
C146 VDD1.n38 VSUBS 0.0122f
C147 VDD1.n39 VSUBS 0.012918f
C148 VDD1.n40 VSUBS 0.028837f
C149 VDD1.n41 VSUBS 0.028837f
C150 VDD1.n42 VSUBS 0.012918f
C151 VDD1.n43 VSUBS 0.0122f
C152 VDD1.n44 VSUBS 0.022705f
C153 VDD1.n45 VSUBS 0.059614f
C154 VDD1.n46 VSUBS 0.0122f
C155 VDD1.n47 VSUBS 0.012918f
C156 VDD1.n48 VSUBS 0.063916f
C157 VDD1.n49 VSUBS 0.061032f
C158 VDD1.t4 VSUBS 0.092401f
C159 VDD1.t0 VSUBS 0.092401f
C160 VDD1.n50 VSUBS 0.602456f
C161 VDD1.n51 VSUBS 1.7016f
C162 VDD1.t3 VSUBS 0.092401f
C163 VDD1.t1 VSUBS 0.092401f
C164 VDD1.n52 VSUBS 0.601305f
C165 VDD1.n53 VSUBS 1.80977f
C166 VTAIL.t0 VSUBS 0.106348f
C167 VTAIL.t3 VSUBS 0.106348f
C168 VTAIL.n0 VSUBS 0.616601f
C169 VTAIL.n1 VSUBS 0.549151f
C170 VTAIL.n2 VSUBS 0.014751f
C171 VTAIL.n3 VSUBS 0.03319f
C172 VTAIL.n4 VSUBS 0.014868f
C173 VTAIL.n5 VSUBS 0.026132f
C174 VTAIL.n6 VSUBS 0.014042f
C175 VTAIL.n7 VSUBS 0.03319f
C176 VTAIL.n8 VSUBS 0.014868f
C177 VTAIL.n9 VSUBS 0.125554f
C178 VTAIL.t10 VSUBS 0.071789f
C179 VTAIL.n10 VSUBS 0.024893f
C180 VTAIL.n11 VSUBS 0.024937f
C181 VTAIL.n12 VSUBS 0.014042f
C182 VTAIL.n13 VSUBS 0.498084f
C183 VTAIL.n14 VSUBS 0.026132f
C184 VTAIL.n15 VSUBS 0.014042f
C185 VTAIL.n16 VSUBS 0.014868f
C186 VTAIL.n17 VSUBS 0.03319f
C187 VTAIL.n18 VSUBS 0.03319f
C188 VTAIL.n19 VSUBS 0.014868f
C189 VTAIL.n20 VSUBS 0.014042f
C190 VTAIL.n21 VSUBS 0.026132f
C191 VTAIL.n22 VSUBS 0.068613f
C192 VTAIL.n23 VSUBS 0.014042f
C193 VTAIL.n24 VSUBS 0.014868f
C194 VTAIL.n25 VSUBS 0.073564f
C195 VTAIL.n26 VSUBS 0.0501f
C196 VTAIL.n27 VSUBS 0.221294f
C197 VTAIL.t9 VSUBS 0.106348f
C198 VTAIL.t7 VSUBS 0.106348f
C199 VTAIL.n28 VSUBS 0.616601f
C200 VTAIL.n29 VSUBS 1.46868f
C201 VTAIL.t5 VSUBS 0.106348f
C202 VTAIL.t1 VSUBS 0.106348f
C203 VTAIL.n30 VSUBS 0.616604f
C204 VTAIL.n31 VSUBS 1.46867f
C205 VTAIL.n32 VSUBS 0.014751f
C206 VTAIL.n33 VSUBS 0.03319f
C207 VTAIL.n34 VSUBS 0.014868f
C208 VTAIL.n35 VSUBS 0.026132f
C209 VTAIL.n36 VSUBS 0.014042f
C210 VTAIL.n37 VSUBS 0.03319f
C211 VTAIL.n38 VSUBS 0.014868f
C212 VTAIL.n39 VSUBS 0.125554f
C213 VTAIL.t4 VSUBS 0.071789f
C214 VTAIL.n40 VSUBS 0.024893f
C215 VTAIL.n41 VSUBS 0.024937f
C216 VTAIL.n42 VSUBS 0.014042f
C217 VTAIL.n43 VSUBS 0.498084f
C218 VTAIL.n44 VSUBS 0.026132f
C219 VTAIL.n45 VSUBS 0.014042f
C220 VTAIL.n46 VSUBS 0.014868f
C221 VTAIL.n47 VSUBS 0.03319f
C222 VTAIL.n48 VSUBS 0.03319f
C223 VTAIL.n49 VSUBS 0.014868f
C224 VTAIL.n50 VSUBS 0.014042f
C225 VTAIL.n51 VSUBS 0.026132f
C226 VTAIL.n52 VSUBS 0.068613f
C227 VTAIL.n53 VSUBS 0.014042f
C228 VTAIL.n54 VSUBS 0.014868f
C229 VTAIL.n55 VSUBS 0.073564f
C230 VTAIL.n56 VSUBS 0.0501f
C231 VTAIL.n57 VSUBS 0.221294f
C232 VTAIL.t8 VSUBS 0.106348f
C233 VTAIL.t6 VSUBS 0.106348f
C234 VTAIL.n58 VSUBS 0.616604f
C235 VTAIL.n59 VSUBS 0.622643f
C236 VTAIL.n60 VSUBS 0.014751f
C237 VTAIL.n61 VSUBS 0.03319f
C238 VTAIL.n62 VSUBS 0.014868f
C239 VTAIL.n63 VSUBS 0.026132f
C240 VTAIL.n64 VSUBS 0.014042f
C241 VTAIL.n65 VSUBS 0.03319f
C242 VTAIL.n66 VSUBS 0.014868f
C243 VTAIL.n67 VSUBS 0.125554f
C244 VTAIL.t11 VSUBS 0.071789f
C245 VTAIL.n68 VSUBS 0.024893f
C246 VTAIL.n69 VSUBS 0.024937f
C247 VTAIL.n70 VSUBS 0.014042f
C248 VTAIL.n71 VSUBS 0.498084f
C249 VTAIL.n72 VSUBS 0.026132f
C250 VTAIL.n73 VSUBS 0.014042f
C251 VTAIL.n74 VSUBS 0.014868f
C252 VTAIL.n75 VSUBS 0.03319f
C253 VTAIL.n76 VSUBS 0.03319f
C254 VTAIL.n77 VSUBS 0.014868f
C255 VTAIL.n78 VSUBS 0.014042f
C256 VTAIL.n79 VSUBS 0.026132f
C257 VTAIL.n80 VSUBS 0.068613f
C258 VTAIL.n81 VSUBS 0.014042f
C259 VTAIL.n82 VSUBS 0.014868f
C260 VTAIL.n83 VSUBS 0.073564f
C261 VTAIL.n84 VSUBS 0.0501f
C262 VTAIL.n85 VSUBS 0.962798f
C263 VTAIL.n86 VSUBS 0.014751f
C264 VTAIL.n87 VSUBS 0.03319f
C265 VTAIL.n88 VSUBS 0.014868f
C266 VTAIL.n89 VSUBS 0.026132f
C267 VTAIL.n90 VSUBS 0.014042f
C268 VTAIL.n91 VSUBS 0.03319f
C269 VTAIL.n92 VSUBS 0.014868f
C270 VTAIL.n93 VSUBS 0.125554f
C271 VTAIL.t2 VSUBS 0.071789f
C272 VTAIL.n94 VSUBS 0.024893f
C273 VTAIL.n95 VSUBS 0.024937f
C274 VTAIL.n96 VSUBS 0.014042f
C275 VTAIL.n97 VSUBS 0.498084f
C276 VTAIL.n98 VSUBS 0.026132f
C277 VTAIL.n99 VSUBS 0.014042f
C278 VTAIL.n100 VSUBS 0.014868f
C279 VTAIL.n101 VSUBS 0.03319f
C280 VTAIL.n102 VSUBS 0.03319f
C281 VTAIL.n103 VSUBS 0.014868f
C282 VTAIL.n104 VSUBS 0.014042f
C283 VTAIL.n105 VSUBS 0.026132f
C284 VTAIL.n106 VSUBS 0.068613f
C285 VTAIL.n107 VSUBS 0.014042f
C286 VTAIL.n108 VSUBS 0.014868f
C287 VTAIL.n109 VSUBS 0.073564f
C288 VTAIL.n110 VSUBS 0.0501f
C289 VTAIL.n111 VSUBS 0.931766f
C290 VP.n0 VSUBS 0.077072f
C291 VP.t1 VSUBS 0.865419f
C292 VP.n1 VSUBS 0.077009f
C293 VP.n2 VSUBS 0.322682f
C294 VP.t4 VSUBS 0.963639f
C295 VP.t2 VSUBS 0.865419f
C296 VP.t3 VSUBS 1.02823f
C297 VP.n3 VSUBS 0.435766f
C298 VP.n4 VSUBS 0.457187f
C299 VP.n5 VSUBS 0.077009f
C300 VP.n6 VSUBS 0.461577f
C301 VP.n7 VSUBS 2.01106f
C302 VP.t0 VSUBS 0.963639f
C303 VP.n8 VSUBS 0.461577f
C304 VP.n9 VSUBS 2.06593f
C305 VP.n10 VSUBS 0.077072f
C306 VP.n11 VSUBS 0.057759f
C307 VP.n12 VSUBS 0.416084f
C308 VP.n13 VSUBS 0.077009f
C309 VP.t5 VSUBS 0.963639f
C310 VP.n14 VSUBS 0.461577f
C311 VP.n15 VSUBS 0.054093f
C312 B.n0 VSUBS 0.004231f
C313 B.n1 VSUBS 0.004231f
C314 B.n2 VSUBS 0.00669f
C315 B.n3 VSUBS 0.00669f
C316 B.n4 VSUBS 0.00669f
C317 B.n5 VSUBS 0.00669f
C318 B.n6 VSUBS 0.00669f
C319 B.n7 VSUBS 0.00669f
C320 B.n8 VSUBS 0.00669f
C321 B.n9 VSUBS 0.00669f
C322 B.n10 VSUBS 0.00669f
C323 B.n11 VSUBS 0.00669f
C324 B.n12 VSUBS 0.00669f
C325 B.n13 VSUBS 0.00669f
C326 B.n14 VSUBS 0.016407f
C327 B.n15 VSUBS 0.00669f
C328 B.n16 VSUBS 0.00669f
C329 B.n17 VSUBS 0.00669f
C330 B.n18 VSUBS 0.00669f
C331 B.n19 VSUBS 0.00669f
C332 B.n20 VSUBS 0.00669f
C333 B.n21 VSUBS 0.00669f
C334 B.n22 VSUBS 0.00669f
C335 B.n23 VSUBS 0.00669f
C336 B.n24 VSUBS 0.00669f
C337 B.n25 VSUBS 0.00669f
C338 B.t11 VSUBS 0.071524f
C339 B.t10 VSUBS 0.083319f
C340 B.t9 VSUBS 0.247726f
C341 B.n26 VSUBS 0.150174f
C342 B.n27 VSUBS 0.128253f
C343 B.n28 VSUBS 0.00669f
C344 B.n29 VSUBS 0.00669f
C345 B.n30 VSUBS 0.00669f
C346 B.n31 VSUBS 0.00669f
C347 B.t2 VSUBS 0.071525f
C348 B.t1 VSUBS 0.083321f
C349 B.t0 VSUBS 0.247726f
C350 B.n32 VSUBS 0.150173f
C351 B.n33 VSUBS 0.128252f
C352 B.n34 VSUBS 0.015501f
C353 B.n35 VSUBS 0.00669f
C354 B.n36 VSUBS 0.00669f
C355 B.n37 VSUBS 0.00669f
C356 B.n38 VSUBS 0.00669f
C357 B.n39 VSUBS 0.00669f
C358 B.n40 VSUBS 0.00669f
C359 B.n41 VSUBS 0.00669f
C360 B.n42 VSUBS 0.00669f
C361 B.n43 VSUBS 0.00669f
C362 B.n44 VSUBS 0.00669f
C363 B.n45 VSUBS 0.016407f
C364 B.n46 VSUBS 0.00669f
C365 B.n47 VSUBS 0.00669f
C366 B.n48 VSUBS 0.00669f
C367 B.n49 VSUBS 0.00669f
C368 B.n50 VSUBS 0.00669f
C369 B.n51 VSUBS 0.00669f
C370 B.n52 VSUBS 0.00669f
C371 B.n53 VSUBS 0.00669f
C372 B.n54 VSUBS 0.00669f
C373 B.n55 VSUBS 0.00669f
C374 B.n56 VSUBS 0.00669f
C375 B.n57 VSUBS 0.00669f
C376 B.n58 VSUBS 0.00669f
C377 B.n59 VSUBS 0.00669f
C378 B.n60 VSUBS 0.00669f
C379 B.n61 VSUBS 0.00669f
C380 B.n62 VSUBS 0.00669f
C381 B.n63 VSUBS 0.00669f
C382 B.n64 VSUBS 0.00669f
C383 B.n65 VSUBS 0.00669f
C384 B.n66 VSUBS 0.00669f
C385 B.n67 VSUBS 0.00669f
C386 B.n68 VSUBS 0.00669f
C387 B.n69 VSUBS 0.00669f
C388 B.n70 VSUBS 0.016407f
C389 B.n71 VSUBS 0.00669f
C390 B.n72 VSUBS 0.00669f
C391 B.n73 VSUBS 0.00669f
C392 B.n74 VSUBS 0.00669f
C393 B.n75 VSUBS 0.00669f
C394 B.n76 VSUBS 0.00669f
C395 B.n77 VSUBS 0.00669f
C396 B.n78 VSUBS 0.00669f
C397 B.n79 VSUBS 0.00669f
C398 B.n80 VSUBS 0.00669f
C399 B.n81 VSUBS 0.00669f
C400 B.t4 VSUBS 0.071525f
C401 B.t5 VSUBS 0.083321f
C402 B.t3 VSUBS 0.247726f
C403 B.n82 VSUBS 0.150173f
C404 B.n83 VSUBS 0.128252f
C405 B.n84 VSUBS 0.00669f
C406 B.n85 VSUBS 0.00669f
C407 B.n86 VSUBS 0.00669f
C408 B.n87 VSUBS 0.00669f
C409 B.t7 VSUBS 0.071524f
C410 B.t8 VSUBS 0.083319f
C411 B.t6 VSUBS 0.247726f
C412 B.n88 VSUBS 0.150174f
C413 B.n89 VSUBS 0.128253f
C414 B.n90 VSUBS 0.015501f
C415 B.n91 VSUBS 0.00669f
C416 B.n92 VSUBS 0.00669f
C417 B.n93 VSUBS 0.00669f
C418 B.n94 VSUBS 0.00669f
C419 B.n95 VSUBS 0.00669f
C420 B.n96 VSUBS 0.00669f
C421 B.n97 VSUBS 0.00669f
C422 B.n98 VSUBS 0.00669f
C423 B.n99 VSUBS 0.00669f
C424 B.n100 VSUBS 0.00669f
C425 B.n101 VSUBS 0.016407f
C426 B.n102 VSUBS 0.00669f
C427 B.n103 VSUBS 0.00669f
C428 B.n104 VSUBS 0.00669f
C429 B.n105 VSUBS 0.00669f
C430 B.n106 VSUBS 0.00669f
C431 B.n107 VSUBS 0.00669f
C432 B.n108 VSUBS 0.00669f
C433 B.n109 VSUBS 0.00669f
C434 B.n110 VSUBS 0.00669f
C435 B.n111 VSUBS 0.00669f
C436 B.n112 VSUBS 0.00669f
C437 B.n113 VSUBS 0.00669f
C438 B.n114 VSUBS 0.00669f
C439 B.n115 VSUBS 0.00669f
C440 B.n116 VSUBS 0.00669f
C441 B.n117 VSUBS 0.00669f
C442 B.n118 VSUBS 0.00669f
C443 B.n119 VSUBS 0.00669f
C444 B.n120 VSUBS 0.00669f
C445 B.n121 VSUBS 0.00669f
C446 B.n122 VSUBS 0.00669f
C447 B.n123 VSUBS 0.00669f
C448 B.n124 VSUBS 0.00669f
C449 B.n125 VSUBS 0.00669f
C450 B.n126 VSUBS 0.00669f
C451 B.n127 VSUBS 0.00669f
C452 B.n128 VSUBS 0.00669f
C453 B.n129 VSUBS 0.00669f
C454 B.n130 VSUBS 0.00669f
C455 B.n131 VSUBS 0.00669f
C456 B.n132 VSUBS 0.00669f
C457 B.n133 VSUBS 0.00669f
C458 B.n134 VSUBS 0.00669f
C459 B.n135 VSUBS 0.00669f
C460 B.n136 VSUBS 0.00669f
C461 B.n137 VSUBS 0.00669f
C462 B.n138 VSUBS 0.00669f
C463 B.n139 VSUBS 0.00669f
C464 B.n140 VSUBS 0.00669f
C465 B.n141 VSUBS 0.00669f
C466 B.n142 VSUBS 0.00669f
C467 B.n143 VSUBS 0.00669f
C468 B.n144 VSUBS 0.00669f
C469 B.n145 VSUBS 0.00669f
C470 B.n146 VSUBS 0.00669f
C471 B.n147 VSUBS 0.00669f
C472 B.n148 VSUBS 0.016407f
C473 B.n149 VSUBS 0.016848f
C474 B.n150 VSUBS 0.016848f
C475 B.n151 VSUBS 0.00669f
C476 B.n152 VSUBS 0.00669f
C477 B.n153 VSUBS 0.00669f
C478 B.n154 VSUBS 0.00669f
C479 B.n155 VSUBS 0.00669f
C480 B.n156 VSUBS 0.00669f
C481 B.n157 VSUBS 0.00669f
C482 B.n158 VSUBS 0.00669f
C483 B.n159 VSUBS 0.00669f
C484 B.n160 VSUBS 0.00669f
C485 B.n161 VSUBS 0.00669f
C486 B.n162 VSUBS 0.00669f
C487 B.n163 VSUBS 0.00669f
C488 B.n164 VSUBS 0.00669f
C489 B.n165 VSUBS 0.00669f
C490 B.n166 VSUBS 0.00669f
C491 B.n167 VSUBS 0.00669f
C492 B.n168 VSUBS 0.00669f
C493 B.n169 VSUBS 0.00669f
C494 B.n170 VSUBS 0.00669f
C495 B.n171 VSUBS 0.00669f
C496 B.n172 VSUBS 0.00669f
C497 B.n173 VSUBS 0.00669f
C498 B.n174 VSUBS 0.00669f
C499 B.n175 VSUBS 0.00669f
C500 B.n176 VSUBS 0.00669f
C501 B.n177 VSUBS 0.00669f
C502 B.n178 VSUBS 0.00669f
C503 B.n179 VSUBS 0.006297f
C504 B.n180 VSUBS 0.00669f
C505 B.n181 VSUBS 0.00669f
C506 B.n182 VSUBS 0.003739f
C507 B.n183 VSUBS 0.00669f
C508 B.n184 VSUBS 0.00669f
C509 B.n185 VSUBS 0.00669f
C510 B.n186 VSUBS 0.00669f
C511 B.n187 VSUBS 0.00669f
C512 B.n188 VSUBS 0.00669f
C513 B.n189 VSUBS 0.00669f
C514 B.n190 VSUBS 0.00669f
C515 B.n191 VSUBS 0.00669f
C516 B.n192 VSUBS 0.00669f
C517 B.n193 VSUBS 0.00669f
C518 B.n194 VSUBS 0.00669f
C519 B.n195 VSUBS 0.003739f
C520 B.n196 VSUBS 0.015501f
C521 B.n197 VSUBS 0.006297f
C522 B.n198 VSUBS 0.00669f
C523 B.n199 VSUBS 0.00669f
C524 B.n200 VSUBS 0.00669f
C525 B.n201 VSUBS 0.00669f
C526 B.n202 VSUBS 0.00669f
C527 B.n203 VSUBS 0.00669f
C528 B.n204 VSUBS 0.00669f
C529 B.n205 VSUBS 0.00669f
C530 B.n206 VSUBS 0.00669f
C531 B.n207 VSUBS 0.00669f
C532 B.n208 VSUBS 0.00669f
C533 B.n209 VSUBS 0.00669f
C534 B.n210 VSUBS 0.00669f
C535 B.n211 VSUBS 0.00669f
C536 B.n212 VSUBS 0.00669f
C537 B.n213 VSUBS 0.00669f
C538 B.n214 VSUBS 0.00669f
C539 B.n215 VSUBS 0.00669f
C540 B.n216 VSUBS 0.00669f
C541 B.n217 VSUBS 0.00669f
C542 B.n218 VSUBS 0.00669f
C543 B.n219 VSUBS 0.00669f
C544 B.n220 VSUBS 0.00669f
C545 B.n221 VSUBS 0.00669f
C546 B.n222 VSUBS 0.00669f
C547 B.n223 VSUBS 0.00669f
C548 B.n224 VSUBS 0.00669f
C549 B.n225 VSUBS 0.00669f
C550 B.n226 VSUBS 0.00669f
C551 B.n227 VSUBS 0.016848f
C552 B.n228 VSUBS 0.016848f
C553 B.n229 VSUBS 0.016407f
C554 B.n230 VSUBS 0.00669f
C555 B.n231 VSUBS 0.00669f
C556 B.n232 VSUBS 0.00669f
C557 B.n233 VSUBS 0.00669f
C558 B.n234 VSUBS 0.00669f
C559 B.n235 VSUBS 0.00669f
C560 B.n236 VSUBS 0.00669f
C561 B.n237 VSUBS 0.00669f
C562 B.n238 VSUBS 0.00669f
C563 B.n239 VSUBS 0.00669f
C564 B.n240 VSUBS 0.00669f
C565 B.n241 VSUBS 0.00669f
C566 B.n242 VSUBS 0.00669f
C567 B.n243 VSUBS 0.00669f
C568 B.n244 VSUBS 0.00669f
C569 B.n245 VSUBS 0.00669f
C570 B.n246 VSUBS 0.00669f
C571 B.n247 VSUBS 0.00669f
C572 B.n248 VSUBS 0.00669f
C573 B.n249 VSUBS 0.00669f
C574 B.n250 VSUBS 0.00669f
C575 B.n251 VSUBS 0.00669f
C576 B.n252 VSUBS 0.00669f
C577 B.n253 VSUBS 0.00669f
C578 B.n254 VSUBS 0.00669f
C579 B.n255 VSUBS 0.00669f
C580 B.n256 VSUBS 0.00669f
C581 B.n257 VSUBS 0.00669f
C582 B.n258 VSUBS 0.00669f
C583 B.n259 VSUBS 0.00669f
C584 B.n260 VSUBS 0.00669f
C585 B.n261 VSUBS 0.00669f
C586 B.n262 VSUBS 0.00669f
C587 B.n263 VSUBS 0.00669f
C588 B.n264 VSUBS 0.00669f
C589 B.n265 VSUBS 0.00669f
C590 B.n266 VSUBS 0.00669f
C591 B.n267 VSUBS 0.00669f
C592 B.n268 VSUBS 0.00669f
C593 B.n269 VSUBS 0.00669f
C594 B.n270 VSUBS 0.00669f
C595 B.n271 VSUBS 0.00669f
C596 B.n272 VSUBS 0.00669f
C597 B.n273 VSUBS 0.00669f
C598 B.n274 VSUBS 0.00669f
C599 B.n275 VSUBS 0.00669f
C600 B.n276 VSUBS 0.00669f
C601 B.n277 VSUBS 0.00669f
C602 B.n278 VSUBS 0.00669f
C603 B.n279 VSUBS 0.00669f
C604 B.n280 VSUBS 0.00669f
C605 B.n281 VSUBS 0.00669f
C606 B.n282 VSUBS 0.00669f
C607 B.n283 VSUBS 0.00669f
C608 B.n284 VSUBS 0.00669f
C609 B.n285 VSUBS 0.00669f
C610 B.n286 VSUBS 0.00669f
C611 B.n287 VSUBS 0.00669f
C612 B.n288 VSUBS 0.00669f
C613 B.n289 VSUBS 0.00669f
C614 B.n290 VSUBS 0.00669f
C615 B.n291 VSUBS 0.00669f
C616 B.n292 VSUBS 0.00669f
C617 B.n293 VSUBS 0.00669f
C618 B.n294 VSUBS 0.00669f
C619 B.n295 VSUBS 0.00669f
C620 B.n296 VSUBS 0.00669f
C621 B.n297 VSUBS 0.00669f
C622 B.n298 VSUBS 0.00669f
C623 B.n299 VSUBS 0.00669f
C624 B.n300 VSUBS 0.00669f
C625 B.n301 VSUBS 0.00669f
C626 B.n302 VSUBS 0.00669f
C627 B.n303 VSUBS 0.00669f
C628 B.n304 VSUBS 0.017129f
C629 B.n305 VSUBS 0.016125f
C630 B.n306 VSUBS 0.016848f
C631 B.n307 VSUBS 0.00669f
C632 B.n308 VSUBS 0.00669f
C633 B.n309 VSUBS 0.00669f
C634 B.n310 VSUBS 0.00669f
C635 B.n311 VSUBS 0.00669f
C636 B.n312 VSUBS 0.00669f
C637 B.n313 VSUBS 0.00669f
C638 B.n314 VSUBS 0.00669f
C639 B.n315 VSUBS 0.00669f
C640 B.n316 VSUBS 0.00669f
C641 B.n317 VSUBS 0.00669f
C642 B.n318 VSUBS 0.00669f
C643 B.n319 VSUBS 0.00669f
C644 B.n320 VSUBS 0.00669f
C645 B.n321 VSUBS 0.00669f
C646 B.n322 VSUBS 0.00669f
C647 B.n323 VSUBS 0.00669f
C648 B.n324 VSUBS 0.00669f
C649 B.n325 VSUBS 0.00669f
C650 B.n326 VSUBS 0.00669f
C651 B.n327 VSUBS 0.00669f
C652 B.n328 VSUBS 0.00669f
C653 B.n329 VSUBS 0.00669f
C654 B.n330 VSUBS 0.00669f
C655 B.n331 VSUBS 0.00669f
C656 B.n332 VSUBS 0.00669f
C657 B.n333 VSUBS 0.00669f
C658 B.n334 VSUBS 0.00669f
C659 B.n335 VSUBS 0.006297f
C660 B.n336 VSUBS 0.00669f
C661 B.n337 VSUBS 0.00669f
C662 B.n338 VSUBS 0.003739f
C663 B.n339 VSUBS 0.00669f
C664 B.n340 VSUBS 0.00669f
C665 B.n341 VSUBS 0.00669f
C666 B.n342 VSUBS 0.00669f
C667 B.n343 VSUBS 0.00669f
C668 B.n344 VSUBS 0.00669f
C669 B.n345 VSUBS 0.00669f
C670 B.n346 VSUBS 0.00669f
C671 B.n347 VSUBS 0.00669f
C672 B.n348 VSUBS 0.00669f
C673 B.n349 VSUBS 0.00669f
C674 B.n350 VSUBS 0.00669f
C675 B.n351 VSUBS 0.003739f
C676 B.n352 VSUBS 0.015501f
C677 B.n353 VSUBS 0.006297f
C678 B.n354 VSUBS 0.00669f
C679 B.n355 VSUBS 0.00669f
C680 B.n356 VSUBS 0.00669f
C681 B.n357 VSUBS 0.00669f
C682 B.n358 VSUBS 0.00669f
C683 B.n359 VSUBS 0.00669f
C684 B.n360 VSUBS 0.00669f
C685 B.n361 VSUBS 0.00669f
C686 B.n362 VSUBS 0.00669f
C687 B.n363 VSUBS 0.00669f
C688 B.n364 VSUBS 0.00669f
C689 B.n365 VSUBS 0.00669f
C690 B.n366 VSUBS 0.00669f
C691 B.n367 VSUBS 0.00669f
C692 B.n368 VSUBS 0.00669f
C693 B.n369 VSUBS 0.00669f
C694 B.n370 VSUBS 0.00669f
C695 B.n371 VSUBS 0.00669f
C696 B.n372 VSUBS 0.00669f
C697 B.n373 VSUBS 0.00669f
C698 B.n374 VSUBS 0.00669f
C699 B.n375 VSUBS 0.00669f
C700 B.n376 VSUBS 0.00669f
C701 B.n377 VSUBS 0.00669f
C702 B.n378 VSUBS 0.00669f
C703 B.n379 VSUBS 0.00669f
C704 B.n380 VSUBS 0.00669f
C705 B.n381 VSUBS 0.00669f
C706 B.n382 VSUBS 0.00669f
C707 B.n383 VSUBS 0.016848f
C708 B.n384 VSUBS 0.016848f
C709 B.n385 VSUBS 0.016407f
C710 B.n386 VSUBS 0.00669f
C711 B.n387 VSUBS 0.00669f
C712 B.n388 VSUBS 0.00669f
C713 B.n389 VSUBS 0.00669f
C714 B.n390 VSUBS 0.00669f
C715 B.n391 VSUBS 0.00669f
C716 B.n392 VSUBS 0.00669f
C717 B.n393 VSUBS 0.00669f
C718 B.n394 VSUBS 0.00669f
C719 B.n395 VSUBS 0.00669f
C720 B.n396 VSUBS 0.00669f
C721 B.n397 VSUBS 0.00669f
C722 B.n398 VSUBS 0.00669f
C723 B.n399 VSUBS 0.00669f
C724 B.n400 VSUBS 0.00669f
C725 B.n401 VSUBS 0.00669f
C726 B.n402 VSUBS 0.00669f
C727 B.n403 VSUBS 0.00669f
C728 B.n404 VSUBS 0.00669f
C729 B.n405 VSUBS 0.00669f
C730 B.n406 VSUBS 0.00669f
C731 B.n407 VSUBS 0.00669f
C732 B.n408 VSUBS 0.00669f
C733 B.n409 VSUBS 0.00669f
C734 B.n410 VSUBS 0.00669f
C735 B.n411 VSUBS 0.00669f
C736 B.n412 VSUBS 0.00669f
C737 B.n413 VSUBS 0.00669f
C738 B.n414 VSUBS 0.00669f
C739 B.n415 VSUBS 0.00669f
C740 B.n416 VSUBS 0.00669f
C741 B.n417 VSUBS 0.00669f
C742 B.n418 VSUBS 0.00669f
C743 B.n419 VSUBS 0.00669f
C744 B.n420 VSUBS 0.00669f
C745 B.n421 VSUBS 0.00669f
C746 B.n422 VSUBS 0.00669f
C747 B.n423 VSUBS 0.015149f
.ends

