* NGSPICE file created from diff_pair_sample_0518.ext - technology: sky130A

.subckt diff_pair_sample_0518 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t4 w_n2518_n2914# sky130_fd_pr__pfet_01v8 ad=1.60545 pd=10.06 as=3.7947 ps=20.24 w=9.73 l=2.25
X1 B.t11 B.t9 B.t10 w_n2518_n2914# sky130_fd_pr__pfet_01v8 ad=3.7947 pd=20.24 as=0 ps=0 w=9.73 l=2.25
X2 VDD1.t2 VP.t1 VTAIL.t6 w_n2518_n2914# sky130_fd_pr__pfet_01v8 ad=1.60545 pd=10.06 as=3.7947 ps=20.24 w=9.73 l=2.25
X3 VDD2.t3 VN.t0 VTAIL.t0 w_n2518_n2914# sky130_fd_pr__pfet_01v8 ad=1.60545 pd=10.06 as=3.7947 ps=20.24 w=9.73 l=2.25
X4 VTAIL.t7 VP.t2 VDD1.t1 w_n2518_n2914# sky130_fd_pr__pfet_01v8 ad=3.7947 pd=20.24 as=1.60545 ps=10.06 w=9.73 l=2.25
X5 B.t8 B.t6 B.t7 w_n2518_n2914# sky130_fd_pr__pfet_01v8 ad=3.7947 pd=20.24 as=0 ps=0 w=9.73 l=2.25
X6 VDD2.t2 VN.t1 VTAIL.t1 w_n2518_n2914# sky130_fd_pr__pfet_01v8 ad=1.60545 pd=10.06 as=3.7947 ps=20.24 w=9.73 l=2.25
X7 B.t5 B.t3 B.t4 w_n2518_n2914# sky130_fd_pr__pfet_01v8 ad=3.7947 pd=20.24 as=0 ps=0 w=9.73 l=2.25
X8 VTAIL.t2 VN.t2 VDD2.t1 w_n2518_n2914# sky130_fd_pr__pfet_01v8 ad=3.7947 pd=20.24 as=1.60545 ps=10.06 w=9.73 l=2.25
X9 B.t2 B.t0 B.t1 w_n2518_n2914# sky130_fd_pr__pfet_01v8 ad=3.7947 pd=20.24 as=0 ps=0 w=9.73 l=2.25
X10 VTAIL.t3 VN.t3 VDD2.t0 w_n2518_n2914# sky130_fd_pr__pfet_01v8 ad=3.7947 pd=20.24 as=1.60545 ps=10.06 w=9.73 l=2.25
X11 VTAIL.t5 VP.t3 VDD1.t0 w_n2518_n2914# sky130_fd_pr__pfet_01v8 ad=3.7947 pd=20.24 as=1.60545 ps=10.06 w=9.73 l=2.25
R0 VP.n12 VP.n0 161.3
R1 VP.n11 VP.n10 161.3
R2 VP.n9 VP.n1 161.3
R3 VP.n8 VP.n7 161.3
R4 VP.n6 VP.n2 161.3
R5 VP.n3 VP.t3 140.242
R6 VP.n3 VP.t1 139.596
R7 VP.n5 VP.t2 104.219
R8 VP.n13 VP.t0 104.219
R9 VP.n5 VP.n4 96.5656
R10 VP.n14 VP.n13 96.5656
R11 VP.n4 VP.n3 49.1784
R12 VP.n7 VP.n1 40.4934
R13 VP.n11 VP.n1 40.4934
R14 VP.n7 VP.n6 24.4675
R15 VP.n12 VP.n11 24.4675
R16 VP.n6 VP.n5 14.1914
R17 VP.n13 VP.n12 14.1914
R18 VP.n4 VP.n2 0.278367
R19 VP.n14 VP.n0 0.278367
R20 VP.n8 VP.n2 0.189894
R21 VP.n9 VP.n8 0.189894
R22 VP.n10 VP.n9 0.189894
R23 VP.n10 VP.n0 0.189894
R24 VP VP.n14 0.153454
R25 VTAIL.n5 VTAIL.t5 67.0034
R26 VTAIL.n4 VTAIL.t0 67.0034
R27 VTAIL.n3 VTAIL.t2 67.0034
R28 VTAIL.n7 VTAIL.t1 67.0033
R29 VTAIL.n0 VTAIL.t3 67.0033
R30 VTAIL.n1 VTAIL.t4 67.0033
R31 VTAIL.n2 VTAIL.t7 67.0033
R32 VTAIL.n6 VTAIL.t6 67.0033
R33 VTAIL.n7 VTAIL.n6 22.9789
R34 VTAIL.n3 VTAIL.n2 22.9789
R35 VTAIL.n4 VTAIL.n3 2.22464
R36 VTAIL.n6 VTAIL.n5 2.22464
R37 VTAIL.n2 VTAIL.n1 2.22464
R38 VTAIL VTAIL.n0 1.17076
R39 VTAIL VTAIL.n7 1.05438
R40 VTAIL.n5 VTAIL.n4 0.470328
R41 VTAIL.n1 VTAIL.n0 0.470328
R42 VDD1 VDD1.n1 119.641
R43 VDD1 VDD1.n0 80.3996
R44 VDD1.n0 VDD1.t0 3.3412
R45 VDD1.n0 VDD1.t2 3.3412
R46 VDD1.n1 VDD1.t1 3.3412
R47 VDD1.n1 VDD1.t3 3.3412
R48 B.n412 B.n411 585
R49 B.n413 B.n60 585
R50 B.n415 B.n414 585
R51 B.n416 B.n59 585
R52 B.n418 B.n417 585
R53 B.n419 B.n58 585
R54 B.n421 B.n420 585
R55 B.n422 B.n57 585
R56 B.n424 B.n423 585
R57 B.n425 B.n56 585
R58 B.n427 B.n426 585
R59 B.n428 B.n55 585
R60 B.n430 B.n429 585
R61 B.n431 B.n54 585
R62 B.n433 B.n432 585
R63 B.n434 B.n53 585
R64 B.n436 B.n435 585
R65 B.n437 B.n52 585
R66 B.n439 B.n438 585
R67 B.n440 B.n51 585
R68 B.n442 B.n441 585
R69 B.n443 B.n50 585
R70 B.n445 B.n444 585
R71 B.n446 B.n49 585
R72 B.n448 B.n447 585
R73 B.n449 B.n48 585
R74 B.n451 B.n450 585
R75 B.n452 B.n47 585
R76 B.n454 B.n453 585
R77 B.n455 B.n46 585
R78 B.n457 B.n456 585
R79 B.n458 B.n45 585
R80 B.n460 B.n459 585
R81 B.n461 B.n44 585
R82 B.n463 B.n462 585
R83 B.n465 B.n41 585
R84 B.n467 B.n466 585
R85 B.n468 B.n40 585
R86 B.n470 B.n469 585
R87 B.n471 B.n39 585
R88 B.n473 B.n472 585
R89 B.n474 B.n38 585
R90 B.n476 B.n475 585
R91 B.n477 B.n35 585
R92 B.n480 B.n479 585
R93 B.n481 B.n34 585
R94 B.n483 B.n482 585
R95 B.n484 B.n33 585
R96 B.n486 B.n485 585
R97 B.n487 B.n32 585
R98 B.n489 B.n488 585
R99 B.n490 B.n31 585
R100 B.n492 B.n491 585
R101 B.n493 B.n30 585
R102 B.n495 B.n494 585
R103 B.n496 B.n29 585
R104 B.n498 B.n497 585
R105 B.n499 B.n28 585
R106 B.n501 B.n500 585
R107 B.n502 B.n27 585
R108 B.n504 B.n503 585
R109 B.n505 B.n26 585
R110 B.n507 B.n506 585
R111 B.n508 B.n25 585
R112 B.n510 B.n509 585
R113 B.n511 B.n24 585
R114 B.n513 B.n512 585
R115 B.n514 B.n23 585
R116 B.n516 B.n515 585
R117 B.n517 B.n22 585
R118 B.n519 B.n518 585
R119 B.n520 B.n21 585
R120 B.n522 B.n521 585
R121 B.n523 B.n20 585
R122 B.n525 B.n524 585
R123 B.n526 B.n19 585
R124 B.n528 B.n527 585
R125 B.n529 B.n18 585
R126 B.n531 B.n530 585
R127 B.n410 B.n61 585
R128 B.n409 B.n408 585
R129 B.n407 B.n62 585
R130 B.n406 B.n405 585
R131 B.n404 B.n63 585
R132 B.n403 B.n402 585
R133 B.n401 B.n64 585
R134 B.n400 B.n399 585
R135 B.n398 B.n65 585
R136 B.n397 B.n396 585
R137 B.n395 B.n66 585
R138 B.n394 B.n393 585
R139 B.n392 B.n67 585
R140 B.n391 B.n390 585
R141 B.n389 B.n68 585
R142 B.n388 B.n387 585
R143 B.n386 B.n69 585
R144 B.n385 B.n384 585
R145 B.n383 B.n70 585
R146 B.n382 B.n381 585
R147 B.n380 B.n71 585
R148 B.n379 B.n378 585
R149 B.n377 B.n72 585
R150 B.n376 B.n375 585
R151 B.n374 B.n73 585
R152 B.n373 B.n372 585
R153 B.n371 B.n74 585
R154 B.n370 B.n369 585
R155 B.n368 B.n75 585
R156 B.n367 B.n366 585
R157 B.n365 B.n76 585
R158 B.n364 B.n363 585
R159 B.n362 B.n77 585
R160 B.n361 B.n360 585
R161 B.n359 B.n78 585
R162 B.n358 B.n357 585
R163 B.n356 B.n79 585
R164 B.n355 B.n354 585
R165 B.n353 B.n80 585
R166 B.n352 B.n351 585
R167 B.n350 B.n81 585
R168 B.n349 B.n348 585
R169 B.n347 B.n82 585
R170 B.n346 B.n345 585
R171 B.n344 B.n83 585
R172 B.n343 B.n342 585
R173 B.n341 B.n84 585
R174 B.n340 B.n339 585
R175 B.n338 B.n85 585
R176 B.n337 B.n336 585
R177 B.n335 B.n86 585
R178 B.n334 B.n333 585
R179 B.n332 B.n87 585
R180 B.n331 B.n330 585
R181 B.n329 B.n88 585
R182 B.n328 B.n327 585
R183 B.n326 B.n89 585
R184 B.n325 B.n324 585
R185 B.n323 B.n90 585
R186 B.n322 B.n321 585
R187 B.n320 B.n91 585
R188 B.n319 B.n318 585
R189 B.n317 B.n92 585
R190 B.n197 B.n136 585
R191 B.n199 B.n198 585
R192 B.n200 B.n135 585
R193 B.n202 B.n201 585
R194 B.n203 B.n134 585
R195 B.n205 B.n204 585
R196 B.n206 B.n133 585
R197 B.n208 B.n207 585
R198 B.n209 B.n132 585
R199 B.n211 B.n210 585
R200 B.n212 B.n131 585
R201 B.n214 B.n213 585
R202 B.n215 B.n130 585
R203 B.n217 B.n216 585
R204 B.n218 B.n129 585
R205 B.n220 B.n219 585
R206 B.n221 B.n128 585
R207 B.n223 B.n222 585
R208 B.n224 B.n127 585
R209 B.n226 B.n225 585
R210 B.n227 B.n126 585
R211 B.n229 B.n228 585
R212 B.n230 B.n125 585
R213 B.n232 B.n231 585
R214 B.n233 B.n124 585
R215 B.n235 B.n234 585
R216 B.n236 B.n123 585
R217 B.n238 B.n237 585
R218 B.n239 B.n122 585
R219 B.n241 B.n240 585
R220 B.n242 B.n121 585
R221 B.n244 B.n243 585
R222 B.n245 B.n120 585
R223 B.n247 B.n246 585
R224 B.n248 B.n117 585
R225 B.n251 B.n250 585
R226 B.n252 B.n116 585
R227 B.n254 B.n253 585
R228 B.n255 B.n115 585
R229 B.n257 B.n256 585
R230 B.n258 B.n114 585
R231 B.n260 B.n259 585
R232 B.n261 B.n113 585
R233 B.n263 B.n262 585
R234 B.n265 B.n264 585
R235 B.n266 B.n109 585
R236 B.n268 B.n267 585
R237 B.n269 B.n108 585
R238 B.n271 B.n270 585
R239 B.n272 B.n107 585
R240 B.n274 B.n273 585
R241 B.n275 B.n106 585
R242 B.n277 B.n276 585
R243 B.n278 B.n105 585
R244 B.n280 B.n279 585
R245 B.n281 B.n104 585
R246 B.n283 B.n282 585
R247 B.n284 B.n103 585
R248 B.n286 B.n285 585
R249 B.n287 B.n102 585
R250 B.n289 B.n288 585
R251 B.n290 B.n101 585
R252 B.n292 B.n291 585
R253 B.n293 B.n100 585
R254 B.n295 B.n294 585
R255 B.n296 B.n99 585
R256 B.n298 B.n297 585
R257 B.n299 B.n98 585
R258 B.n301 B.n300 585
R259 B.n302 B.n97 585
R260 B.n304 B.n303 585
R261 B.n305 B.n96 585
R262 B.n307 B.n306 585
R263 B.n308 B.n95 585
R264 B.n310 B.n309 585
R265 B.n311 B.n94 585
R266 B.n313 B.n312 585
R267 B.n314 B.n93 585
R268 B.n316 B.n315 585
R269 B.n196 B.n195 585
R270 B.n194 B.n137 585
R271 B.n193 B.n192 585
R272 B.n191 B.n138 585
R273 B.n190 B.n189 585
R274 B.n188 B.n139 585
R275 B.n187 B.n186 585
R276 B.n185 B.n140 585
R277 B.n184 B.n183 585
R278 B.n182 B.n141 585
R279 B.n181 B.n180 585
R280 B.n179 B.n142 585
R281 B.n178 B.n177 585
R282 B.n176 B.n143 585
R283 B.n175 B.n174 585
R284 B.n173 B.n144 585
R285 B.n172 B.n171 585
R286 B.n170 B.n145 585
R287 B.n169 B.n168 585
R288 B.n167 B.n146 585
R289 B.n166 B.n165 585
R290 B.n164 B.n147 585
R291 B.n163 B.n162 585
R292 B.n161 B.n148 585
R293 B.n160 B.n159 585
R294 B.n158 B.n149 585
R295 B.n157 B.n156 585
R296 B.n155 B.n150 585
R297 B.n154 B.n153 585
R298 B.n152 B.n151 585
R299 B.n2 B.n0 585
R300 B.n577 B.n1 585
R301 B.n576 B.n575 585
R302 B.n574 B.n3 585
R303 B.n573 B.n572 585
R304 B.n571 B.n4 585
R305 B.n570 B.n569 585
R306 B.n568 B.n5 585
R307 B.n567 B.n566 585
R308 B.n565 B.n6 585
R309 B.n564 B.n563 585
R310 B.n562 B.n7 585
R311 B.n561 B.n560 585
R312 B.n559 B.n8 585
R313 B.n558 B.n557 585
R314 B.n556 B.n9 585
R315 B.n555 B.n554 585
R316 B.n553 B.n10 585
R317 B.n552 B.n551 585
R318 B.n550 B.n11 585
R319 B.n549 B.n548 585
R320 B.n547 B.n12 585
R321 B.n546 B.n545 585
R322 B.n544 B.n13 585
R323 B.n543 B.n542 585
R324 B.n541 B.n14 585
R325 B.n540 B.n539 585
R326 B.n538 B.n15 585
R327 B.n537 B.n536 585
R328 B.n535 B.n16 585
R329 B.n534 B.n533 585
R330 B.n532 B.n17 585
R331 B.n579 B.n578 585
R332 B.n197 B.n196 516.524
R333 B.n530 B.n17 516.524
R334 B.n317 B.n316 516.524
R335 B.n412 B.n61 516.524
R336 B.n110 B.t6 311.67
R337 B.n118 B.t3 311.67
R338 B.n36 B.t9 311.67
R339 B.n42 B.t0 311.67
R340 B.n196 B.n137 163.367
R341 B.n192 B.n137 163.367
R342 B.n192 B.n191 163.367
R343 B.n191 B.n190 163.367
R344 B.n190 B.n139 163.367
R345 B.n186 B.n139 163.367
R346 B.n186 B.n185 163.367
R347 B.n185 B.n184 163.367
R348 B.n184 B.n141 163.367
R349 B.n180 B.n141 163.367
R350 B.n180 B.n179 163.367
R351 B.n179 B.n178 163.367
R352 B.n178 B.n143 163.367
R353 B.n174 B.n143 163.367
R354 B.n174 B.n173 163.367
R355 B.n173 B.n172 163.367
R356 B.n172 B.n145 163.367
R357 B.n168 B.n145 163.367
R358 B.n168 B.n167 163.367
R359 B.n167 B.n166 163.367
R360 B.n166 B.n147 163.367
R361 B.n162 B.n147 163.367
R362 B.n162 B.n161 163.367
R363 B.n161 B.n160 163.367
R364 B.n160 B.n149 163.367
R365 B.n156 B.n149 163.367
R366 B.n156 B.n155 163.367
R367 B.n155 B.n154 163.367
R368 B.n154 B.n151 163.367
R369 B.n151 B.n2 163.367
R370 B.n578 B.n2 163.367
R371 B.n578 B.n577 163.367
R372 B.n577 B.n576 163.367
R373 B.n576 B.n3 163.367
R374 B.n572 B.n3 163.367
R375 B.n572 B.n571 163.367
R376 B.n571 B.n570 163.367
R377 B.n570 B.n5 163.367
R378 B.n566 B.n5 163.367
R379 B.n566 B.n565 163.367
R380 B.n565 B.n564 163.367
R381 B.n564 B.n7 163.367
R382 B.n560 B.n7 163.367
R383 B.n560 B.n559 163.367
R384 B.n559 B.n558 163.367
R385 B.n558 B.n9 163.367
R386 B.n554 B.n9 163.367
R387 B.n554 B.n553 163.367
R388 B.n553 B.n552 163.367
R389 B.n552 B.n11 163.367
R390 B.n548 B.n11 163.367
R391 B.n548 B.n547 163.367
R392 B.n547 B.n546 163.367
R393 B.n546 B.n13 163.367
R394 B.n542 B.n13 163.367
R395 B.n542 B.n541 163.367
R396 B.n541 B.n540 163.367
R397 B.n540 B.n15 163.367
R398 B.n536 B.n15 163.367
R399 B.n536 B.n535 163.367
R400 B.n535 B.n534 163.367
R401 B.n534 B.n17 163.367
R402 B.n198 B.n197 163.367
R403 B.n198 B.n135 163.367
R404 B.n202 B.n135 163.367
R405 B.n203 B.n202 163.367
R406 B.n204 B.n203 163.367
R407 B.n204 B.n133 163.367
R408 B.n208 B.n133 163.367
R409 B.n209 B.n208 163.367
R410 B.n210 B.n209 163.367
R411 B.n210 B.n131 163.367
R412 B.n214 B.n131 163.367
R413 B.n215 B.n214 163.367
R414 B.n216 B.n215 163.367
R415 B.n216 B.n129 163.367
R416 B.n220 B.n129 163.367
R417 B.n221 B.n220 163.367
R418 B.n222 B.n221 163.367
R419 B.n222 B.n127 163.367
R420 B.n226 B.n127 163.367
R421 B.n227 B.n226 163.367
R422 B.n228 B.n227 163.367
R423 B.n228 B.n125 163.367
R424 B.n232 B.n125 163.367
R425 B.n233 B.n232 163.367
R426 B.n234 B.n233 163.367
R427 B.n234 B.n123 163.367
R428 B.n238 B.n123 163.367
R429 B.n239 B.n238 163.367
R430 B.n240 B.n239 163.367
R431 B.n240 B.n121 163.367
R432 B.n244 B.n121 163.367
R433 B.n245 B.n244 163.367
R434 B.n246 B.n245 163.367
R435 B.n246 B.n117 163.367
R436 B.n251 B.n117 163.367
R437 B.n252 B.n251 163.367
R438 B.n253 B.n252 163.367
R439 B.n253 B.n115 163.367
R440 B.n257 B.n115 163.367
R441 B.n258 B.n257 163.367
R442 B.n259 B.n258 163.367
R443 B.n259 B.n113 163.367
R444 B.n263 B.n113 163.367
R445 B.n264 B.n263 163.367
R446 B.n264 B.n109 163.367
R447 B.n268 B.n109 163.367
R448 B.n269 B.n268 163.367
R449 B.n270 B.n269 163.367
R450 B.n270 B.n107 163.367
R451 B.n274 B.n107 163.367
R452 B.n275 B.n274 163.367
R453 B.n276 B.n275 163.367
R454 B.n276 B.n105 163.367
R455 B.n280 B.n105 163.367
R456 B.n281 B.n280 163.367
R457 B.n282 B.n281 163.367
R458 B.n282 B.n103 163.367
R459 B.n286 B.n103 163.367
R460 B.n287 B.n286 163.367
R461 B.n288 B.n287 163.367
R462 B.n288 B.n101 163.367
R463 B.n292 B.n101 163.367
R464 B.n293 B.n292 163.367
R465 B.n294 B.n293 163.367
R466 B.n294 B.n99 163.367
R467 B.n298 B.n99 163.367
R468 B.n299 B.n298 163.367
R469 B.n300 B.n299 163.367
R470 B.n300 B.n97 163.367
R471 B.n304 B.n97 163.367
R472 B.n305 B.n304 163.367
R473 B.n306 B.n305 163.367
R474 B.n306 B.n95 163.367
R475 B.n310 B.n95 163.367
R476 B.n311 B.n310 163.367
R477 B.n312 B.n311 163.367
R478 B.n312 B.n93 163.367
R479 B.n316 B.n93 163.367
R480 B.n318 B.n317 163.367
R481 B.n318 B.n91 163.367
R482 B.n322 B.n91 163.367
R483 B.n323 B.n322 163.367
R484 B.n324 B.n323 163.367
R485 B.n324 B.n89 163.367
R486 B.n328 B.n89 163.367
R487 B.n329 B.n328 163.367
R488 B.n330 B.n329 163.367
R489 B.n330 B.n87 163.367
R490 B.n334 B.n87 163.367
R491 B.n335 B.n334 163.367
R492 B.n336 B.n335 163.367
R493 B.n336 B.n85 163.367
R494 B.n340 B.n85 163.367
R495 B.n341 B.n340 163.367
R496 B.n342 B.n341 163.367
R497 B.n342 B.n83 163.367
R498 B.n346 B.n83 163.367
R499 B.n347 B.n346 163.367
R500 B.n348 B.n347 163.367
R501 B.n348 B.n81 163.367
R502 B.n352 B.n81 163.367
R503 B.n353 B.n352 163.367
R504 B.n354 B.n353 163.367
R505 B.n354 B.n79 163.367
R506 B.n358 B.n79 163.367
R507 B.n359 B.n358 163.367
R508 B.n360 B.n359 163.367
R509 B.n360 B.n77 163.367
R510 B.n364 B.n77 163.367
R511 B.n365 B.n364 163.367
R512 B.n366 B.n365 163.367
R513 B.n366 B.n75 163.367
R514 B.n370 B.n75 163.367
R515 B.n371 B.n370 163.367
R516 B.n372 B.n371 163.367
R517 B.n372 B.n73 163.367
R518 B.n376 B.n73 163.367
R519 B.n377 B.n376 163.367
R520 B.n378 B.n377 163.367
R521 B.n378 B.n71 163.367
R522 B.n382 B.n71 163.367
R523 B.n383 B.n382 163.367
R524 B.n384 B.n383 163.367
R525 B.n384 B.n69 163.367
R526 B.n388 B.n69 163.367
R527 B.n389 B.n388 163.367
R528 B.n390 B.n389 163.367
R529 B.n390 B.n67 163.367
R530 B.n394 B.n67 163.367
R531 B.n395 B.n394 163.367
R532 B.n396 B.n395 163.367
R533 B.n396 B.n65 163.367
R534 B.n400 B.n65 163.367
R535 B.n401 B.n400 163.367
R536 B.n402 B.n401 163.367
R537 B.n402 B.n63 163.367
R538 B.n406 B.n63 163.367
R539 B.n407 B.n406 163.367
R540 B.n408 B.n407 163.367
R541 B.n408 B.n61 163.367
R542 B.n530 B.n529 163.367
R543 B.n529 B.n528 163.367
R544 B.n528 B.n19 163.367
R545 B.n524 B.n19 163.367
R546 B.n524 B.n523 163.367
R547 B.n523 B.n522 163.367
R548 B.n522 B.n21 163.367
R549 B.n518 B.n21 163.367
R550 B.n518 B.n517 163.367
R551 B.n517 B.n516 163.367
R552 B.n516 B.n23 163.367
R553 B.n512 B.n23 163.367
R554 B.n512 B.n511 163.367
R555 B.n511 B.n510 163.367
R556 B.n510 B.n25 163.367
R557 B.n506 B.n25 163.367
R558 B.n506 B.n505 163.367
R559 B.n505 B.n504 163.367
R560 B.n504 B.n27 163.367
R561 B.n500 B.n27 163.367
R562 B.n500 B.n499 163.367
R563 B.n499 B.n498 163.367
R564 B.n498 B.n29 163.367
R565 B.n494 B.n29 163.367
R566 B.n494 B.n493 163.367
R567 B.n493 B.n492 163.367
R568 B.n492 B.n31 163.367
R569 B.n488 B.n31 163.367
R570 B.n488 B.n487 163.367
R571 B.n487 B.n486 163.367
R572 B.n486 B.n33 163.367
R573 B.n482 B.n33 163.367
R574 B.n482 B.n481 163.367
R575 B.n481 B.n480 163.367
R576 B.n480 B.n35 163.367
R577 B.n475 B.n35 163.367
R578 B.n475 B.n474 163.367
R579 B.n474 B.n473 163.367
R580 B.n473 B.n39 163.367
R581 B.n469 B.n39 163.367
R582 B.n469 B.n468 163.367
R583 B.n468 B.n467 163.367
R584 B.n467 B.n41 163.367
R585 B.n462 B.n41 163.367
R586 B.n462 B.n461 163.367
R587 B.n461 B.n460 163.367
R588 B.n460 B.n45 163.367
R589 B.n456 B.n45 163.367
R590 B.n456 B.n455 163.367
R591 B.n455 B.n454 163.367
R592 B.n454 B.n47 163.367
R593 B.n450 B.n47 163.367
R594 B.n450 B.n449 163.367
R595 B.n449 B.n448 163.367
R596 B.n448 B.n49 163.367
R597 B.n444 B.n49 163.367
R598 B.n444 B.n443 163.367
R599 B.n443 B.n442 163.367
R600 B.n442 B.n51 163.367
R601 B.n438 B.n51 163.367
R602 B.n438 B.n437 163.367
R603 B.n437 B.n436 163.367
R604 B.n436 B.n53 163.367
R605 B.n432 B.n53 163.367
R606 B.n432 B.n431 163.367
R607 B.n431 B.n430 163.367
R608 B.n430 B.n55 163.367
R609 B.n426 B.n55 163.367
R610 B.n426 B.n425 163.367
R611 B.n425 B.n424 163.367
R612 B.n424 B.n57 163.367
R613 B.n420 B.n57 163.367
R614 B.n420 B.n419 163.367
R615 B.n419 B.n418 163.367
R616 B.n418 B.n59 163.367
R617 B.n414 B.n59 163.367
R618 B.n414 B.n413 163.367
R619 B.n413 B.n412 163.367
R620 B.n110 B.t8 161.889
R621 B.n42 B.t1 161.889
R622 B.n118 B.t5 161.879
R623 B.n36 B.t10 161.879
R624 B.n111 B.t7 111.853
R625 B.n43 B.t2 111.853
R626 B.n119 B.t4 111.841
R627 B.n37 B.t11 111.841
R628 B.n112 B.n111 59.5399
R629 B.n249 B.n119 59.5399
R630 B.n478 B.n37 59.5399
R631 B.n464 B.n43 59.5399
R632 B.n111 B.n110 50.0369
R633 B.n119 B.n118 50.0369
R634 B.n37 B.n36 50.0369
R635 B.n43 B.n42 50.0369
R636 B.n532 B.n531 33.5615
R637 B.n411 B.n410 33.5615
R638 B.n315 B.n92 33.5615
R639 B.n195 B.n136 33.5615
R640 B B.n579 18.0485
R641 B.n531 B.n18 10.6151
R642 B.n527 B.n18 10.6151
R643 B.n527 B.n526 10.6151
R644 B.n526 B.n525 10.6151
R645 B.n525 B.n20 10.6151
R646 B.n521 B.n20 10.6151
R647 B.n521 B.n520 10.6151
R648 B.n520 B.n519 10.6151
R649 B.n519 B.n22 10.6151
R650 B.n515 B.n22 10.6151
R651 B.n515 B.n514 10.6151
R652 B.n514 B.n513 10.6151
R653 B.n513 B.n24 10.6151
R654 B.n509 B.n24 10.6151
R655 B.n509 B.n508 10.6151
R656 B.n508 B.n507 10.6151
R657 B.n507 B.n26 10.6151
R658 B.n503 B.n26 10.6151
R659 B.n503 B.n502 10.6151
R660 B.n502 B.n501 10.6151
R661 B.n501 B.n28 10.6151
R662 B.n497 B.n28 10.6151
R663 B.n497 B.n496 10.6151
R664 B.n496 B.n495 10.6151
R665 B.n495 B.n30 10.6151
R666 B.n491 B.n30 10.6151
R667 B.n491 B.n490 10.6151
R668 B.n490 B.n489 10.6151
R669 B.n489 B.n32 10.6151
R670 B.n485 B.n32 10.6151
R671 B.n485 B.n484 10.6151
R672 B.n484 B.n483 10.6151
R673 B.n483 B.n34 10.6151
R674 B.n479 B.n34 10.6151
R675 B.n477 B.n476 10.6151
R676 B.n476 B.n38 10.6151
R677 B.n472 B.n38 10.6151
R678 B.n472 B.n471 10.6151
R679 B.n471 B.n470 10.6151
R680 B.n470 B.n40 10.6151
R681 B.n466 B.n40 10.6151
R682 B.n466 B.n465 10.6151
R683 B.n463 B.n44 10.6151
R684 B.n459 B.n44 10.6151
R685 B.n459 B.n458 10.6151
R686 B.n458 B.n457 10.6151
R687 B.n457 B.n46 10.6151
R688 B.n453 B.n46 10.6151
R689 B.n453 B.n452 10.6151
R690 B.n452 B.n451 10.6151
R691 B.n451 B.n48 10.6151
R692 B.n447 B.n48 10.6151
R693 B.n447 B.n446 10.6151
R694 B.n446 B.n445 10.6151
R695 B.n445 B.n50 10.6151
R696 B.n441 B.n50 10.6151
R697 B.n441 B.n440 10.6151
R698 B.n440 B.n439 10.6151
R699 B.n439 B.n52 10.6151
R700 B.n435 B.n52 10.6151
R701 B.n435 B.n434 10.6151
R702 B.n434 B.n433 10.6151
R703 B.n433 B.n54 10.6151
R704 B.n429 B.n54 10.6151
R705 B.n429 B.n428 10.6151
R706 B.n428 B.n427 10.6151
R707 B.n427 B.n56 10.6151
R708 B.n423 B.n56 10.6151
R709 B.n423 B.n422 10.6151
R710 B.n422 B.n421 10.6151
R711 B.n421 B.n58 10.6151
R712 B.n417 B.n58 10.6151
R713 B.n417 B.n416 10.6151
R714 B.n416 B.n415 10.6151
R715 B.n415 B.n60 10.6151
R716 B.n411 B.n60 10.6151
R717 B.n319 B.n92 10.6151
R718 B.n320 B.n319 10.6151
R719 B.n321 B.n320 10.6151
R720 B.n321 B.n90 10.6151
R721 B.n325 B.n90 10.6151
R722 B.n326 B.n325 10.6151
R723 B.n327 B.n326 10.6151
R724 B.n327 B.n88 10.6151
R725 B.n331 B.n88 10.6151
R726 B.n332 B.n331 10.6151
R727 B.n333 B.n332 10.6151
R728 B.n333 B.n86 10.6151
R729 B.n337 B.n86 10.6151
R730 B.n338 B.n337 10.6151
R731 B.n339 B.n338 10.6151
R732 B.n339 B.n84 10.6151
R733 B.n343 B.n84 10.6151
R734 B.n344 B.n343 10.6151
R735 B.n345 B.n344 10.6151
R736 B.n345 B.n82 10.6151
R737 B.n349 B.n82 10.6151
R738 B.n350 B.n349 10.6151
R739 B.n351 B.n350 10.6151
R740 B.n351 B.n80 10.6151
R741 B.n355 B.n80 10.6151
R742 B.n356 B.n355 10.6151
R743 B.n357 B.n356 10.6151
R744 B.n357 B.n78 10.6151
R745 B.n361 B.n78 10.6151
R746 B.n362 B.n361 10.6151
R747 B.n363 B.n362 10.6151
R748 B.n363 B.n76 10.6151
R749 B.n367 B.n76 10.6151
R750 B.n368 B.n367 10.6151
R751 B.n369 B.n368 10.6151
R752 B.n369 B.n74 10.6151
R753 B.n373 B.n74 10.6151
R754 B.n374 B.n373 10.6151
R755 B.n375 B.n374 10.6151
R756 B.n375 B.n72 10.6151
R757 B.n379 B.n72 10.6151
R758 B.n380 B.n379 10.6151
R759 B.n381 B.n380 10.6151
R760 B.n381 B.n70 10.6151
R761 B.n385 B.n70 10.6151
R762 B.n386 B.n385 10.6151
R763 B.n387 B.n386 10.6151
R764 B.n387 B.n68 10.6151
R765 B.n391 B.n68 10.6151
R766 B.n392 B.n391 10.6151
R767 B.n393 B.n392 10.6151
R768 B.n393 B.n66 10.6151
R769 B.n397 B.n66 10.6151
R770 B.n398 B.n397 10.6151
R771 B.n399 B.n398 10.6151
R772 B.n399 B.n64 10.6151
R773 B.n403 B.n64 10.6151
R774 B.n404 B.n403 10.6151
R775 B.n405 B.n404 10.6151
R776 B.n405 B.n62 10.6151
R777 B.n409 B.n62 10.6151
R778 B.n410 B.n409 10.6151
R779 B.n199 B.n136 10.6151
R780 B.n200 B.n199 10.6151
R781 B.n201 B.n200 10.6151
R782 B.n201 B.n134 10.6151
R783 B.n205 B.n134 10.6151
R784 B.n206 B.n205 10.6151
R785 B.n207 B.n206 10.6151
R786 B.n207 B.n132 10.6151
R787 B.n211 B.n132 10.6151
R788 B.n212 B.n211 10.6151
R789 B.n213 B.n212 10.6151
R790 B.n213 B.n130 10.6151
R791 B.n217 B.n130 10.6151
R792 B.n218 B.n217 10.6151
R793 B.n219 B.n218 10.6151
R794 B.n219 B.n128 10.6151
R795 B.n223 B.n128 10.6151
R796 B.n224 B.n223 10.6151
R797 B.n225 B.n224 10.6151
R798 B.n225 B.n126 10.6151
R799 B.n229 B.n126 10.6151
R800 B.n230 B.n229 10.6151
R801 B.n231 B.n230 10.6151
R802 B.n231 B.n124 10.6151
R803 B.n235 B.n124 10.6151
R804 B.n236 B.n235 10.6151
R805 B.n237 B.n236 10.6151
R806 B.n237 B.n122 10.6151
R807 B.n241 B.n122 10.6151
R808 B.n242 B.n241 10.6151
R809 B.n243 B.n242 10.6151
R810 B.n243 B.n120 10.6151
R811 B.n247 B.n120 10.6151
R812 B.n248 B.n247 10.6151
R813 B.n250 B.n116 10.6151
R814 B.n254 B.n116 10.6151
R815 B.n255 B.n254 10.6151
R816 B.n256 B.n255 10.6151
R817 B.n256 B.n114 10.6151
R818 B.n260 B.n114 10.6151
R819 B.n261 B.n260 10.6151
R820 B.n262 B.n261 10.6151
R821 B.n266 B.n265 10.6151
R822 B.n267 B.n266 10.6151
R823 B.n267 B.n108 10.6151
R824 B.n271 B.n108 10.6151
R825 B.n272 B.n271 10.6151
R826 B.n273 B.n272 10.6151
R827 B.n273 B.n106 10.6151
R828 B.n277 B.n106 10.6151
R829 B.n278 B.n277 10.6151
R830 B.n279 B.n278 10.6151
R831 B.n279 B.n104 10.6151
R832 B.n283 B.n104 10.6151
R833 B.n284 B.n283 10.6151
R834 B.n285 B.n284 10.6151
R835 B.n285 B.n102 10.6151
R836 B.n289 B.n102 10.6151
R837 B.n290 B.n289 10.6151
R838 B.n291 B.n290 10.6151
R839 B.n291 B.n100 10.6151
R840 B.n295 B.n100 10.6151
R841 B.n296 B.n295 10.6151
R842 B.n297 B.n296 10.6151
R843 B.n297 B.n98 10.6151
R844 B.n301 B.n98 10.6151
R845 B.n302 B.n301 10.6151
R846 B.n303 B.n302 10.6151
R847 B.n303 B.n96 10.6151
R848 B.n307 B.n96 10.6151
R849 B.n308 B.n307 10.6151
R850 B.n309 B.n308 10.6151
R851 B.n309 B.n94 10.6151
R852 B.n313 B.n94 10.6151
R853 B.n314 B.n313 10.6151
R854 B.n315 B.n314 10.6151
R855 B.n195 B.n194 10.6151
R856 B.n194 B.n193 10.6151
R857 B.n193 B.n138 10.6151
R858 B.n189 B.n138 10.6151
R859 B.n189 B.n188 10.6151
R860 B.n188 B.n187 10.6151
R861 B.n187 B.n140 10.6151
R862 B.n183 B.n140 10.6151
R863 B.n183 B.n182 10.6151
R864 B.n182 B.n181 10.6151
R865 B.n181 B.n142 10.6151
R866 B.n177 B.n142 10.6151
R867 B.n177 B.n176 10.6151
R868 B.n176 B.n175 10.6151
R869 B.n175 B.n144 10.6151
R870 B.n171 B.n144 10.6151
R871 B.n171 B.n170 10.6151
R872 B.n170 B.n169 10.6151
R873 B.n169 B.n146 10.6151
R874 B.n165 B.n146 10.6151
R875 B.n165 B.n164 10.6151
R876 B.n164 B.n163 10.6151
R877 B.n163 B.n148 10.6151
R878 B.n159 B.n148 10.6151
R879 B.n159 B.n158 10.6151
R880 B.n158 B.n157 10.6151
R881 B.n157 B.n150 10.6151
R882 B.n153 B.n150 10.6151
R883 B.n153 B.n152 10.6151
R884 B.n152 B.n0 10.6151
R885 B.n575 B.n1 10.6151
R886 B.n575 B.n574 10.6151
R887 B.n574 B.n573 10.6151
R888 B.n573 B.n4 10.6151
R889 B.n569 B.n4 10.6151
R890 B.n569 B.n568 10.6151
R891 B.n568 B.n567 10.6151
R892 B.n567 B.n6 10.6151
R893 B.n563 B.n6 10.6151
R894 B.n563 B.n562 10.6151
R895 B.n562 B.n561 10.6151
R896 B.n561 B.n8 10.6151
R897 B.n557 B.n8 10.6151
R898 B.n557 B.n556 10.6151
R899 B.n556 B.n555 10.6151
R900 B.n555 B.n10 10.6151
R901 B.n551 B.n10 10.6151
R902 B.n551 B.n550 10.6151
R903 B.n550 B.n549 10.6151
R904 B.n549 B.n12 10.6151
R905 B.n545 B.n12 10.6151
R906 B.n545 B.n544 10.6151
R907 B.n544 B.n543 10.6151
R908 B.n543 B.n14 10.6151
R909 B.n539 B.n14 10.6151
R910 B.n539 B.n538 10.6151
R911 B.n538 B.n537 10.6151
R912 B.n537 B.n16 10.6151
R913 B.n533 B.n16 10.6151
R914 B.n533 B.n532 10.6151
R915 B.n478 B.n477 6.5566
R916 B.n465 B.n464 6.5566
R917 B.n250 B.n249 6.5566
R918 B.n262 B.n112 6.5566
R919 B.n479 B.n478 4.05904
R920 B.n464 B.n463 4.05904
R921 B.n249 B.n248 4.05904
R922 B.n265 B.n112 4.05904
R923 B.n579 B.n0 2.81026
R924 B.n579 B.n1 2.81026
R925 VN.n0 VN.t3 140.242
R926 VN.n1 VN.t0 140.242
R927 VN.n0 VN.t1 139.596
R928 VN.n1 VN.t2 139.596
R929 VN VN.n1 49.4572
R930 VN VN.n0 5.70346
R931 VDD2.n2 VDD2.n0 119.117
R932 VDD2.n2 VDD2.n1 80.3414
R933 VDD2.n1 VDD2.t1 3.3412
R934 VDD2.n1 VDD2.t3 3.3412
R935 VDD2.n0 VDD2.t0 3.3412
R936 VDD2.n0 VDD2.t2 3.3412
R937 VDD2 VDD2.n2 0.0586897
C0 VDD2 VTAIL 4.85315f
C1 VDD2 VP 0.371863f
C2 VN VTAIL 3.76391f
C3 VN VP 5.5198f
C4 VDD1 VTAIL 4.80128f
C5 VDD1 VP 4.03166f
C6 VTAIL w_n2518_n2914# 3.45507f
C7 B VTAIL 4.05392f
C8 VP w_n2518_n2914# 4.48617f
C9 B VP 1.54969f
C10 VDD2 VN 3.80896f
C11 VDD2 VDD1 0.944436f
C12 VDD2 w_n2518_n2914# 1.37012f
C13 VDD2 B 1.18659f
C14 VDD1 VN 0.148512f
C15 VN w_n2518_n2914# 4.16335f
C16 B VN 1.01562f
C17 VDD1 w_n2518_n2914# 1.32184f
C18 VDD1 B 1.14019f
C19 B w_n2518_n2914# 8.17926f
C20 VP VTAIL 3.77801f
C21 VDD2 VSUBS 0.829262f
C22 VDD1 VSUBS 5.212046f
C23 VTAIL VSUBS 1.063947f
C24 VN VSUBS 5.23404f
C25 VP VSUBS 2.020309f
C26 B VSUBS 3.77762f
C27 w_n2518_n2914# VSUBS 90.67821f
C28 VDD2.t0 VSUBS 0.207929f
C29 VDD2.t2 VSUBS 0.207929f
C30 VDD2.n0 VSUBS 2.144f
C31 VDD2.t1 VSUBS 0.207929f
C32 VDD2.t3 VSUBS 0.207929f
C33 VDD2.n1 VSUBS 1.56906f
C34 VDD2.n2 VSUBS 3.95559f
C35 VN.t3 VSUBS 2.49586f
C36 VN.t1 VSUBS 2.49121f
C37 VN.n0 VSUBS 1.64062f
C38 VN.t0 VSUBS 2.49586f
C39 VN.t2 VSUBS 2.49121f
C40 VN.n1 VSUBS 3.41604f
C41 B.n0 VSUBS 0.004656f
C42 B.n1 VSUBS 0.004656f
C43 B.n2 VSUBS 0.007363f
C44 B.n3 VSUBS 0.007363f
C45 B.n4 VSUBS 0.007363f
C46 B.n5 VSUBS 0.007363f
C47 B.n6 VSUBS 0.007363f
C48 B.n7 VSUBS 0.007363f
C49 B.n8 VSUBS 0.007363f
C50 B.n9 VSUBS 0.007363f
C51 B.n10 VSUBS 0.007363f
C52 B.n11 VSUBS 0.007363f
C53 B.n12 VSUBS 0.007363f
C54 B.n13 VSUBS 0.007363f
C55 B.n14 VSUBS 0.007363f
C56 B.n15 VSUBS 0.007363f
C57 B.n16 VSUBS 0.007363f
C58 B.n17 VSUBS 0.017386f
C59 B.n18 VSUBS 0.007363f
C60 B.n19 VSUBS 0.007363f
C61 B.n20 VSUBS 0.007363f
C62 B.n21 VSUBS 0.007363f
C63 B.n22 VSUBS 0.007363f
C64 B.n23 VSUBS 0.007363f
C65 B.n24 VSUBS 0.007363f
C66 B.n25 VSUBS 0.007363f
C67 B.n26 VSUBS 0.007363f
C68 B.n27 VSUBS 0.007363f
C69 B.n28 VSUBS 0.007363f
C70 B.n29 VSUBS 0.007363f
C71 B.n30 VSUBS 0.007363f
C72 B.n31 VSUBS 0.007363f
C73 B.n32 VSUBS 0.007363f
C74 B.n33 VSUBS 0.007363f
C75 B.n34 VSUBS 0.007363f
C76 B.n35 VSUBS 0.007363f
C77 B.t11 VSUBS 0.325206f
C78 B.t10 VSUBS 0.344771f
C79 B.t9 VSUBS 1.05218f
C80 B.n36 VSUBS 0.176121f
C81 B.n37 VSUBS 0.073798f
C82 B.n38 VSUBS 0.007363f
C83 B.n39 VSUBS 0.007363f
C84 B.n40 VSUBS 0.007363f
C85 B.n41 VSUBS 0.007363f
C86 B.t2 VSUBS 0.325202f
C87 B.t1 VSUBS 0.344767f
C88 B.t0 VSUBS 1.05218f
C89 B.n42 VSUBS 0.176125f
C90 B.n43 VSUBS 0.073802f
C91 B.n44 VSUBS 0.007363f
C92 B.n45 VSUBS 0.007363f
C93 B.n46 VSUBS 0.007363f
C94 B.n47 VSUBS 0.007363f
C95 B.n48 VSUBS 0.007363f
C96 B.n49 VSUBS 0.007363f
C97 B.n50 VSUBS 0.007363f
C98 B.n51 VSUBS 0.007363f
C99 B.n52 VSUBS 0.007363f
C100 B.n53 VSUBS 0.007363f
C101 B.n54 VSUBS 0.007363f
C102 B.n55 VSUBS 0.007363f
C103 B.n56 VSUBS 0.007363f
C104 B.n57 VSUBS 0.007363f
C105 B.n58 VSUBS 0.007363f
C106 B.n59 VSUBS 0.007363f
C107 B.n60 VSUBS 0.007363f
C108 B.n61 VSUBS 0.017386f
C109 B.n62 VSUBS 0.007363f
C110 B.n63 VSUBS 0.007363f
C111 B.n64 VSUBS 0.007363f
C112 B.n65 VSUBS 0.007363f
C113 B.n66 VSUBS 0.007363f
C114 B.n67 VSUBS 0.007363f
C115 B.n68 VSUBS 0.007363f
C116 B.n69 VSUBS 0.007363f
C117 B.n70 VSUBS 0.007363f
C118 B.n71 VSUBS 0.007363f
C119 B.n72 VSUBS 0.007363f
C120 B.n73 VSUBS 0.007363f
C121 B.n74 VSUBS 0.007363f
C122 B.n75 VSUBS 0.007363f
C123 B.n76 VSUBS 0.007363f
C124 B.n77 VSUBS 0.007363f
C125 B.n78 VSUBS 0.007363f
C126 B.n79 VSUBS 0.007363f
C127 B.n80 VSUBS 0.007363f
C128 B.n81 VSUBS 0.007363f
C129 B.n82 VSUBS 0.007363f
C130 B.n83 VSUBS 0.007363f
C131 B.n84 VSUBS 0.007363f
C132 B.n85 VSUBS 0.007363f
C133 B.n86 VSUBS 0.007363f
C134 B.n87 VSUBS 0.007363f
C135 B.n88 VSUBS 0.007363f
C136 B.n89 VSUBS 0.007363f
C137 B.n90 VSUBS 0.007363f
C138 B.n91 VSUBS 0.007363f
C139 B.n92 VSUBS 0.017386f
C140 B.n93 VSUBS 0.007363f
C141 B.n94 VSUBS 0.007363f
C142 B.n95 VSUBS 0.007363f
C143 B.n96 VSUBS 0.007363f
C144 B.n97 VSUBS 0.007363f
C145 B.n98 VSUBS 0.007363f
C146 B.n99 VSUBS 0.007363f
C147 B.n100 VSUBS 0.007363f
C148 B.n101 VSUBS 0.007363f
C149 B.n102 VSUBS 0.007363f
C150 B.n103 VSUBS 0.007363f
C151 B.n104 VSUBS 0.007363f
C152 B.n105 VSUBS 0.007363f
C153 B.n106 VSUBS 0.007363f
C154 B.n107 VSUBS 0.007363f
C155 B.n108 VSUBS 0.007363f
C156 B.n109 VSUBS 0.007363f
C157 B.t7 VSUBS 0.325202f
C158 B.t8 VSUBS 0.344767f
C159 B.t6 VSUBS 1.05218f
C160 B.n110 VSUBS 0.176125f
C161 B.n111 VSUBS 0.073802f
C162 B.n112 VSUBS 0.017059f
C163 B.n113 VSUBS 0.007363f
C164 B.n114 VSUBS 0.007363f
C165 B.n115 VSUBS 0.007363f
C166 B.n116 VSUBS 0.007363f
C167 B.n117 VSUBS 0.007363f
C168 B.t4 VSUBS 0.325206f
C169 B.t5 VSUBS 0.344771f
C170 B.t3 VSUBS 1.05218f
C171 B.n118 VSUBS 0.176121f
C172 B.n119 VSUBS 0.073798f
C173 B.n120 VSUBS 0.007363f
C174 B.n121 VSUBS 0.007363f
C175 B.n122 VSUBS 0.007363f
C176 B.n123 VSUBS 0.007363f
C177 B.n124 VSUBS 0.007363f
C178 B.n125 VSUBS 0.007363f
C179 B.n126 VSUBS 0.007363f
C180 B.n127 VSUBS 0.007363f
C181 B.n128 VSUBS 0.007363f
C182 B.n129 VSUBS 0.007363f
C183 B.n130 VSUBS 0.007363f
C184 B.n131 VSUBS 0.007363f
C185 B.n132 VSUBS 0.007363f
C186 B.n133 VSUBS 0.007363f
C187 B.n134 VSUBS 0.007363f
C188 B.n135 VSUBS 0.007363f
C189 B.n136 VSUBS 0.017696f
C190 B.n137 VSUBS 0.007363f
C191 B.n138 VSUBS 0.007363f
C192 B.n139 VSUBS 0.007363f
C193 B.n140 VSUBS 0.007363f
C194 B.n141 VSUBS 0.007363f
C195 B.n142 VSUBS 0.007363f
C196 B.n143 VSUBS 0.007363f
C197 B.n144 VSUBS 0.007363f
C198 B.n145 VSUBS 0.007363f
C199 B.n146 VSUBS 0.007363f
C200 B.n147 VSUBS 0.007363f
C201 B.n148 VSUBS 0.007363f
C202 B.n149 VSUBS 0.007363f
C203 B.n150 VSUBS 0.007363f
C204 B.n151 VSUBS 0.007363f
C205 B.n152 VSUBS 0.007363f
C206 B.n153 VSUBS 0.007363f
C207 B.n154 VSUBS 0.007363f
C208 B.n155 VSUBS 0.007363f
C209 B.n156 VSUBS 0.007363f
C210 B.n157 VSUBS 0.007363f
C211 B.n158 VSUBS 0.007363f
C212 B.n159 VSUBS 0.007363f
C213 B.n160 VSUBS 0.007363f
C214 B.n161 VSUBS 0.007363f
C215 B.n162 VSUBS 0.007363f
C216 B.n163 VSUBS 0.007363f
C217 B.n164 VSUBS 0.007363f
C218 B.n165 VSUBS 0.007363f
C219 B.n166 VSUBS 0.007363f
C220 B.n167 VSUBS 0.007363f
C221 B.n168 VSUBS 0.007363f
C222 B.n169 VSUBS 0.007363f
C223 B.n170 VSUBS 0.007363f
C224 B.n171 VSUBS 0.007363f
C225 B.n172 VSUBS 0.007363f
C226 B.n173 VSUBS 0.007363f
C227 B.n174 VSUBS 0.007363f
C228 B.n175 VSUBS 0.007363f
C229 B.n176 VSUBS 0.007363f
C230 B.n177 VSUBS 0.007363f
C231 B.n178 VSUBS 0.007363f
C232 B.n179 VSUBS 0.007363f
C233 B.n180 VSUBS 0.007363f
C234 B.n181 VSUBS 0.007363f
C235 B.n182 VSUBS 0.007363f
C236 B.n183 VSUBS 0.007363f
C237 B.n184 VSUBS 0.007363f
C238 B.n185 VSUBS 0.007363f
C239 B.n186 VSUBS 0.007363f
C240 B.n187 VSUBS 0.007363f
C241 B.n188 VSUBS 0.007363f
C242 B.n189 VSUBS 0.007363f
C243 B.n190 VSUBS 0.007363f
C244 B.n191 VSUBS 0.007363f
C245 B.n192 VSUBS 0.007363f
C246 B.n193 VSUBS 0.007363f
C247 B.n194 VSUBS 0.007363f
C248 B.n195 VSUBS 0.017386f
C249 B.n196 VSUBS 0.017386f
C250 B.n197 VSUBS 0.017696f
C251 B.n198 VSUBS 0.007363f
C252 B.n199 VSUBS 0.007363f
C253 B.n200 VSUBS 0.007363f
C254 B.n201 VSUBS 0.007363f
C255 B.n202 VSUBS 0.007363f
C256 B.n203 VSUBS 0.007363f
C257 B.n204 VSUBS 0.007363f
C258 B.n205 VSUBS 0.007363f
C259 B.n206 VSUBS 0.007363f
C260 B.n207 VSUBS 0.007363f
C261 B.n208 VSUBS 0.007363f
C262 B.n209 VSUBS 0.007363f
C263 B.n210 VSUBS 0.007363f
C264 B.n211 VSUBS 0.007363f
C265 B.n212 VSUBS 0.007363f
C266 B.n213 VSUBS 0.007363f
C267 B.n214 VSUBS 0.007363f
C268 B.n215 VSUBS 0.007363f
C269 B.n216 VSUBS 0.007363f
C270 B.n217 VSUBS 0.007363f
C271 B.n218 VSUBS 0.007363f
C272 B.n219 VSUBS 0.007363f
C273 B.n220 VSUBS 0.007363f
C274 B.n221 VSUBS 0.007363f
C275 B.n222 VSUBS 0.007363f
C276 B.n223 VSUBS 0.007363f
C277 B.n224 VSUBS 0.007363f
C278 B.n225 VSUBS 0.007363f
C279 B.n226 VSUBS 0.007363f
C280 B.n227 VSUBS 0.007363f
C281 B.n228 VSUBS 0.007363f
C282 B.n229 VSUBS 0.007363f
C283 B.n230 VSUBS 0.007363f
C284 B.n231 VSUBS 0.007363f
C285 B.n232 VSUBS 0.007363f
C286 B.n233 VSUBS 0.007363f
C287 B.n234 VSUBS 0.007363f
C288 B.n235 VSUBS 0.007363f
C289 B.n236 VSUBS 0.007363f
C290 B.n237 VSUBS 0.007363f
C291 B.n238 VSUBS 0.007363f
C292 B.n239 VSUBS 0.007363f
C293 B.n240 VSUBS 0.007363f
C294 B.n241 VSUBS 0.007363f
C295 B.n242 VSUBS 0.007363f
C296 B.n243 VSUBS 0.007363f
C297 B.n244 VSUBS 0.007363f
C298 B.n245 VSUBS 0.007363f
C299 B.n246 VSUBS 0.007363f
C300 B.n247 VSUBS 0.007363f
C301 B.n248 VSUBS 0.005089f
C302 B.n249 VSUBS 0.017059f
C303 B.n250 VSUBS 0.005955f
C304 B.n251 VSUBS 0.007363f
C305 B.n252 VSUBS 0.007363f
C306 B.n253 VSUBS 0.007363f
C307 B.n254 VSUBS 0.007363f
C308 B.n255 VSUBS 0.007363f
C309 B.n256 VSUBS 0.007363f
C310 B.n257 VSUBS 0.007363f
C311 B.n258 VSUBS 0.007363f
C312 B.n259 VSUBS 0.007363f
C313 B.n260 VSUBS 0.007363f
C314 B.n261 VSUBS 0.007363f
C315 B.n262 VSUBS 0.005955f
C316 B.n263 VSUBS 0.007363f
C317 B.n264 VSUBS 0.007363f
C318 B.n265 VSUBS 0.005089f
C319 B.n266 VSUBS 0.007363f
C320 B.n267 VSUBS 0.007363f
C321 B.n268 VSUBS 0.007363f
C322 B.n269 VSUBS 0.007363f
C323 B.n270 VSUBS 0.007363f
C324 B.n271 VSUBS 0.007363f
C325 B.n272 VSUBS 0.007363f
C326 B.n273 VSUBS 0.007363f
C327 B.n274 VSUBS 0.007363f
C328 B.n275 VSUBS 0.007363f
C329 B.n276 VSUBS 0.007363f
C330 B.n277 VSUBS 0.007363f
C331 B.n278 VSUBS 0.007363f
C332 B.n279 VSUBS 0.007363f
C333 B.n280 VSUBS 0.007363f
C334 B.n281 VSUBS 0.007363f
C335 B.n282 VSUBS 0.007363f
C336 B.n283 VSUBS 0.007363f
C337 B.n284 VSUBS 0.007363f
C338 B.n285 VSUBS 0.007363f
C339 B.n286 VSUBS 0.007363f
C340 B.n287 VSUBS 0.007363f
C341 B.n288 VSUBS 0.007363f
C342 B.n289 VSUBS 0.007363f
C343 B.n290 VSUBS 0.007363f
C344 B.n291 VSUBS 0.007363f
C345 B.n292 VSUBS 0.007363f
C346 B.n293 VSUBS 0.007363f
C347 B.n294 VSUBS 0.007363f
C348 B.n295 VSUBS 0.007363f
C349 B.n296 VSUBS 0.007363f
C350 B.n297 VSUBS 0.007363f
C351 B.n298 VSUBS 0.007363f
C352 B.n299 VSUBS 0.007363f
C353 B.n300 VSUBS 0.007363f
C354 B.n301 VSUBS 0.007363f
C355 B.n302 VSUBS 0.007363f
C356 B.n303 VSUBS 0.007363f
C357 B.n304 VSUBS 0.007363f
C358 B.n305 VSUBS 0.007363f
C359 B.n306 VSUBS 0.007363f
C360 B.n307 VSUBS 0.007363f
C361 B.n308 VSUBS 0.007363f
C362 B.n309 VSUBS 0.007363f
C363 B.n310 VSUBS 0.007363f
C364 B.n311 VSUBS 0.007363f
C365 B.n312 VSUBS 0.007363f
C366 B.n313 VSUBS 0.007363f
C367 B.n314 VSUBS 0.007363f
C368 B.n315 VSUBS 0.017696f
C369 B.n316 VSUBS 0.017696f
C370 B.n317 VSUBS 0.017386f
C371 B.n318 VSUBS 0.007363f
C372 B.n319 VSUBS 0.007363f
C373 B.n320 VSUBS 0.007363f
C374 B.n321 VSUBS 0.007363f
C375 B.n322 VSUBS 0.007363f
C376 B.n323 VSUBS 0.007363f
C377 B.n324 VSUBS 0.007363f
C378 B.n325 VSUBS 0.007363f
C379 B.n326 VSUBS 0.007363f
C380 B.n327 VSUBS 0.007363f
C381 B.n328 VSUBS 0.007363f
C382 B.n329 VSUBS 0.007363f
C383 B.n330 VSUBS 0.007363f
C384 B.n331 VSUBS 0.007363f
C385 B.n332 VSUBS 0.007363f
C386 B.n333 VSUBS 0.007363f
C387 B.n334 VSUBS 0.007363f
C388 B.n335 VSUBS 0.007363f
C389 B.n336 VSUBS 0.007363f
C390 B.n337 VSUBS 0.007363f
C391 B.n338 VSUBS 0.007363f
C392 B.n339 VSUBS 0.007363f
C393 B.n340 VSUBS 0.007363f
C394 B.n341 VSUBS 0.007363f
C395 B.n342 VSUBS 0.007363f
C396 B.n343 VSUBS 0.007363f
C397 B.n344 VSUBS 0.007363f
C398 B.n345 VSUBS 0.007363f
C399 B.n346 VSUBS 0.007363f
C400 B.n347 VSUBS 0.007363f
C401 B.n348 VSUBS 0.007363f
C402 B.n349 VSUBS 0.007363f
C403 B.n350 VSUBS 0.007363f
C404 B.n351 VSUBS 0.007363f
C405 B.n352 VSUBS 0.007363f
C406 B.n353 VSUBS 0.007363f
C407 B.n354 VSUBS 0.007363f
C408 B.n355 VSUBS 0.007363f
C409 B.n356 VSUBS 0.007363f
C410 B.n357 VSUBS 0.007363f
C411 B.n358 VSUBS 0.007363f
C412 B.n359 VSUBS 0.007363f
C413 B.n360 VSUBS 0.007363f
C414 B.n361 VSUBS 0.007363f
C415 B.n362 VSUBS 0.007363f
C416 B.n363 VSUBS 0.007363f
C417 B.n364 VSUBS 0.007363f
C418 B.n365 VSUBS 0.007363f
C419 B.n366 VSUBS 0.007363f
C420 B.n367 VSUBS 0.007363f
C421 B.n368 VSUBS 0.007363f
C422 B.n369 VSUBS 0.007363f
C423 B.n370 VSUBS 0.007363f
C424 B.n371 VSUBS 0.007363f
C425 B.n372 VSUBS 0.007363f
C426 B.n373 VSUBS 0.007363f
C427 B.n374 VSUBS 0.007363f
C428 B.n375 VSUBS 0.007363f
C429 B.n376 VSUBS 0.007363f
C430 B.n377 VSUBS 0.007363f
C431 B.n378 VSUBS 0.007363f
C432 B.n379 VSUBS 0.007363f
C433 B.n380 VSUBS 0.007363f
C434 B.n381 VSUBS 0.007363f
C435 B.n382 VSUBS 0.007363f
C436 B.n383 VSUBS 0.007363f
C437 B.n384 VSUBS 0.007363f
C438 B.n385 VSUBS 0.007363f
C439 B.n386 VSUBS 0.007363f
C440 B.n387 VSUBS 0.007363f
C441 B.n388 VSUBS 0.007363f
C442 B.n389 VSUBS 0.007363f
C443 B.n390 VSUBS 0.007363f
C444 B.n391 VSUBS 0.007363f
C445 B.n392 VSUBS 0.007363f
C446 B.n393 VSUBS 0.007363f
C447 B.n394 VSUBS 0.007363f
C448 B.n395 VSUBS 0.007363f
C449 B.n396 VSUBS 0.007363f
C450 B.n397 VSUBS 0.007363f
C451 B.n398 VSUBS 0.007363f
C452 B.n399 VSUBS 0.007363f
C453 B.n400 VSUBS 0.007363f
C454 B.n401 VSUBS 0.007363f
C455 B.n402 VSUBS 0.007363f
C456 B.n403 VSUBS 0.007363f
C457 B.n404 VSUBS 0.007363f
C458 B.n405 VSUBS 0.007363f
C459 B.n406 VSUBS 0.007363f
C460 B.n407 VSUBS 0.007363f
C461 B.n408 VSUBS 0.007363f
C462 B.n409 VSUBS 0.007363f
C463 B.n410 VSUBS 0.018233f
C464 B.n411 VSUBS 0.016849f
C465 B.n412 VSUBS 0.017696f
C466 B.n413 VSUBS 0.007363f
C467 B.n414 VSUBS 0.007363f
C468 B.n415 VSUBS 0.007363f
C469 B.n416 VSUBS 0.007363f
C470 B.n417 VSUBS 0.007363f
C471 B.n418 VSUBS 0.007363f
C472 B.n419 VSUBS 0.007363f
C473 B.n420 VSUBS 0.007363f
C474 B.n421 VSUBS 0.007363f
C475 B.n422 VSUBS 0.007363f
C476 B.n423 VSUBS 0.007363f
C477 B.n424 VSUBS 0.007363f
C478 B.n425 VSUBS 0.007363f
C479 B.n426 VSUBS 0.007363f
C480 B.n427 VSUBS 0.007363f
C481 B.n428 VSUBS 0.007363f
C482 B.n429 VSUBS 0.007363f
C483 B.n430 VSUBS 0.007363f
C484 B.n431 VSUBS 0.007363f
C485 B.n432 VSUBS 0.007363f
C486 B.n433 VSUBS 0.007363f
C487 B.n434 VSUBS 0.007363f
C488 B.n435 VSUBS 0.007363f
C489 B.n436 VSUBS 0.007363f
C490 B.n437 VSUBS 0.007363f
C491 B.n438 VSUBS 0.007363f
C492 B.n439 VSUBS 0.007363f
C493 B.n440 VSUBS 0.007363f
C494 B.n441 VSUBS 0.007363f
C495 B.n442 VSUBS 0.007363f
C496 B.n443 VSUBS 0.007363f
C497 B.n444 VSUBS 0.007363f
C498 B.n445 VSUBS 0.007363f
C499 B.n446 VSUBS 0.007363f
C500 B.n447 VSUBS 0.007363f
C501 B.n448 VSUBS 0.007363f
C502 B.n449 VSUBS 0.007363f
C503 B.n450 VSUBS 0.007363f
C504 B.n451 VSUBS 0.007363f
C505 B.n452 VSUBS 0.007363f
C506 B.n453 VSUBS 0.007363f
C507 B.n454 VSUBS 0.007363f
C508 B.n455 VSUBS 0.007363f
C509 B.n456 VSUBS 0.007363f
C510 B.n457 VSUBS 0.007363f
C511 B.n458 VSUBS 0.007363f
C512 B.n459 VSUBS 0.007363f
C513 B.n460 VSUBS 0.007363f
C514 B.n461 VSUBS 0.007363f
C515 B.n462 VSUBS 0.007363f
C516 B.n463 VSUBS 0.005089f
C517 B.n464 VSUBS 0.017059f
C518 B.n465 VSUBS 0.005955f
C519 B.n466 VSUBS 0.007363f
C520 B.n467 VSUBS 0.007363f
C521 B.n468 VSUBS 0.007363f
C522 B.n469 VSUBS 0.007363f
C523 B.n470 VSUBS 0.007363f
C524 B.n471 VSUBS 0.007363f
C525 B.n472 VSUBS 0.007363f
C526 B.n473 VSUBS 0.007363f
C527 B.n474 VSUBS 0.007363f
C528 B.n475 VSUBS 0.007363f
C529 B.n476 VSUBS 0.007363f
C530 B.n477 VSUBS 0.005955f
C531 B.n478 VSUBS 0.017059f
C532 B.n479 VSUBS 0.005089f
C533 B.n480 VSUBS 0.007363f
C534 B.n481 VSUBS 0.007363f
C535 B.n482 VSUBS 0.007363f
C536 B.n483 VSUBS 0.007363f
C537 B.n484 VSUBS 0.007363f
C538 B.n485 VSUBS 0.007363f
C539 B.n486 VSUBS 0.007363f
C540 B.n487 VSUBS 0.007363f
C541 B.n488 VSUBS 0.007363f
C542 B.n489 VSUBS 0.007363f
C543 B.n490 VSUBS 0.007363f
C544 B.n491 VSUBS 0.007363f
C545 B.n492 VSUBS 0.007363f
C546 B.n493 VSUBS 0.007363f
C547 B.n494 VSUBS 0.007363f
C548 B.n495 VSUBS 0.007363f
C549 B.n496 VSUBS 0.007363f
C550 B.n497 VSUBS 0.007363f
C551 B.n498 VSUBS 0.007363f
C552 B.n499 VSUBS 0.007363f
C553 B.n500 VSUBS 0.007363f
C554 B.n501 VSUBS 0.007363f
C555 B.n502 VSUBS 0.007363f
C556 B.n503 VSUBS 0.007363f
C557 B.n504 VSUBS 0.007363f
C558 B.n505 VSUBS 0.007363f
C559 B.n506 VSUBS 0.007363f
C560 B.n507 VSUBS 0.007363f
C561 B.n508 VSUBS 0.007363f
C562 B.n509 VSUBS 0.007363f
C563 B.n510 VSUBS 0.007363f
C564 B.n511 VSUBS 0.007363f
C565 B.n512 VSUBS 0.007363f
C566 B.n513 VSUBS 0.007363f
C567 B.n514 VSUBS 0.007363f
C568 B.n515 VSUBS 0.007363f
C569 B.n516 VSUBS 0.007363f
C570 B.n517 VSUBS 0.007363f
C571 B.n518 VSUBS 0.007363f
C572 B.n519 VSUBS 0.007363f
C573 B.n520 VSUBS 0.007363f
C574 B.n521 VSUBS 0.007363f
C575 B.n522 VSUBS 0.007363f
C576 B.n523 VSUBS 0.007363f
C577 B.n524 VSUBS 0.007363f
C578 B.n525 VSUBS 0.007363f
C579 B.n526 VSUBS 0.007363f
C580 B.n527 VSUBS 0.007363f
C581 B.n528 VSUBS 0.007363f
C582 B.n529 VSUBS 0.007363f
C583 B.n530 VSUBS 0.017696f
C584 B.n531 VSUBS 0.017696f
C585 B.n532 VSUBS 0.017386f
C586 B.n533 VSUBS 0.007363f
C587 B.n534 VSUBS 0.007363f
C588 B.n535 VSUBS 0.007363f
C589 B.n536 VSUBS 0.007363f
C590 B.n537 VSUBS 0.007363f
C591 B.n538 VSUBS 0.007363f
C592 B.n539 VSUBS 0.007363f
C593 B.n540 VSUBS 0.007363f
C594 B.n541 VSUBS 0.007363f
C595 B.n542 VSUBS 0.007363f
C596 B.n543 VSUBS 0.007363f
C597 B.n544 VSUBS 0.007363f
C598 B.n545 VSUBS 0.007363f
C599 B.n546 VSUBS 0.007363f
C600 B.n547 VSUBS 0.007363f
C601 B.n548 VSUBS 0.007363f
C602 B.n549 VSUBS 0.007363f
C603 B.n550 VSUBS 0.007363f
C604 B.n551 VSUBS 0.007363f
C605 B.n552 VSUBS 0.007363f
C606 B.n553 VSUBS 0.007363f
C607 B.n554 VSUBS 0.007363f
C608 B.n555 VSUBS 0.007363f
C609 B.n556 VSUBS 0.007363f
C610 B.n557 VSUBS 0.007363f
C611 B.n558 VSUBS 0.007363f
C612 B.n559 VSUBS 0.007363f
C613 B.n560 VSUBS 0.007363f
C614 B.n561 VSUBS 0.007363f
C615 B.n562 VSUBS 0.007363f
C616 B.n563 VSUBS 0.007363f
C617 B.n564 VSUBS 0.007363f
C618 B.n565 VSUBS 0.007363f
C619 B.n566 VSUBS 0.007363f
C620 B.n567 VSUBS 0.007363f
C621 B.n568 VSUBS 0.007363f
C622 B.n569 VSUBS 0.007363f
C623 B.n570 VSUBS 0.007363f
C624 B.n571 VSUBS 0.007363f
C625 B.n572 VSUBS 0.007363f
C626 B.n573 VSUBS 0.007363f
C627 B.n574 VSUBS 0.007363f
C628 B.n575 VSUBS 0.007363f
C629 B.n576 VSUBS 0.007363f
C630 B.n577 VSUBS 0.007363f
C631 B.n578 VSUBS 0.007363f
C632 B.n579 VSUBS 0.016672f
C633 VDD1.t0 VSUBS 0.207932f
C634 VDD1.t2 VSUBS 0.207932f
C635 VDD1.n0 VSUBS 1.56958f
C636 VDD1.t1 VSUBS 0.207932f
C637 VDD1.t3 VSUBS 0.207932f
C638 VDD1.n1 VSUBS 2.16707f
C639 VTAIL.t3 VSUBS 1.74029f
C640 VTAIL.n0 VSUBS 0.722726f
C641 VTAIL.t4 VSUBS 1.74029f
C642 VTAIL.n1 VSUBS 0.805866f
C643 VTAIL.t7 VSUBS 1.74029f
C644 VTAIL.n2 VSUBS 1.93855f
C645 VTAIL.t2 VSUBS 1.7403f
C646 VTAIL.n3 VSUBS 1.93854f
C647 VTAIL.t0 VSUBS 1.7403f
C648 VTAIL.n4 VSUBS 0.805854f
C649 VTAIL.t5 VSUBS 1.7403f
C650 VTAIL.n5 VSUBS 0.805854f
C651 VTAIL.t6 VSUBS 1.74029f
C652 VTAIL.n6 VSUBS 1.93855f
C653 VTAIL.t1 VSUBS 1.74029f
C654 VTAIL.n7 VSUBS 1.84623f
C655 VP.n0 VSUBS 0.051281f
C656 VP.t0 VSUBS 2.30467f
C657 VP.n1 VSUBS 0.031444f
C658 VP.n2 VSUBS 0.051281f
C659 VP.t2 VSUBS 2.30467f
C660 VP.t1 VSUBS 2.57108f
C661 VP.t3 VSUBS 2.57588f
C662 VP.n3 VSUBS 3.50527f
C663 VP.n4 VSUBS 2.0137f
C664 VP.n5 VSUBS 0.952068f
C665 VP.n6 VSUBS 0.057461f
C666 VP.n7 VSUBS 0.077307f
C667 VP.n8 VSUBS 0.038897f
C668 VP.n9 VSUBS 0.038897f
C669 VP.n10 VSUBS 0.038897f
C670 VP.n11 VSUBS 0.077307f
C671 VP.n12 VSUBS 0.057461f
C672 VP.n13 VSUBS 0.952068f
C673 VP.n14 VSUBS 0.055208f
.ends

