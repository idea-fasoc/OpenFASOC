* NGSPICE file created from diff_pair_sample_1366.ext - technology: sky130A

.subckt diff_pair_sample_1366 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t4 VP.t0 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.4329 pd=3 as=0.18315 ps=1.44 w=1.11 l=1.5
X1 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=0.4329 pd=3 as=0 ps=0 w=1.11 l=1.5
X2 VDD1.t1 VP.t1 VTAIL.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.18315 pd=1.44 as=0.4329 ps=3 w=1.11 l=1.5
X3 VDD2.t3 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.18315 pd=1.44 as=0.4329 ps=3 w=1.11 l=1.5
X4 VDD1.t0 VP.t2 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.18315 pd=1.44 as=0.4329 ps=3 w=1.11 l=1.5
X5 VTAIL.t5 VN.t1 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=0.4329 pd=3 as=0.18315 ps=1.44 w=1.11 l=1.5
X6 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=0.4329 pd=3 as=0 ps=0 w=1.11 l=1.5
X7 VTAIL.t1 VP.t3 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4329 pd=3 as=0.18315 ps=1.44 w=1.11 l=1.5
X8 VDD2.t1 VN.t2 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.18315 pd=1.44 as=0.4329 ps=3 w=1.11 l=1.5
X9 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=0.4329 pd=3 as=0 ps=0 w=1.11 l=1.5
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.4329 pd=3 as=0 ps=0 w=1.11 l=1.5
X11 VTAIL.t7 VN.t3 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4329 pd=3 as=0.18315 ps=1.44 w=1.11 l=1.5
R0 VP.n4 VP.n3 177.694
R1 VP.n12 VP.n11 177.694
R2 VP.n10 VP.n0 161.3
R3 VP.n9 VP.n8 161.3
R4 VP.n7 VP.n1 161.3
R5 VP.n6 VP.n5 161.3
R6 VP.n9 VP.n1 56.5193
R7 VP.n2 VP.t3 54.1947
R8 VP.n2 VP.t2 53.8783
R9 VP.n3 VP.n2 47.6345
R10 VP.n5 VP.n1 24.4675
R11 VP.n10 VP.n9 24.4675
R12 VP.n4 VP.t0 17.8345
R13 VP.n11 VP.t1 17.8345
R14 VP.n5 VP.n4 8.07461
R15 VP.n11 VP.n10 8.07461
R16 VP.n6 VP.n3 0.189894
R17 VP.n7 VP.n6 0.189894
R18 VP.n8 VP.n7 0.189894
R19 VP.n8 VP.n0 0.189894
R20 VP.n12 VP.n0 0.189894
R21 VP VP.n12 0.0516364
R22 VDD1 VDD1.n1 176.362
R23 VDD1 VDD1.n0 146.49
R24 VDD1.n0 VDD1.t2 17.8383
R25 VDD1.n0 VDD1.t0 17.8383
R26 VDD1.n1 VDD1.t3 17.8383
R27 VDD1.n1 VDD1.t1 17.8383
R28 VTAIL.n7 VTAIL.t0 155.916
R29 VTAIL.n0 VTAIL.t7 155.916
R30 VTAIL.n1 VTAIL.t3 155.916
R31 VTAIL.n2 VTAIL.t4 155.916
R32 VTAIL.n6 VTAIL.t2 155.916
R33 VTAIL.n5 VTAIL.t1 155.916
R34 VTAIL.n4 VTAIL.t6 155.916
R35 VTAIL.n3 VTAIL.t5 155.916
R36 VTAIL.n7 VTAIL.n6 14.9014
R37 VTAIL.n3 VTAIL.n2 14.9014
R38 VTAIL.n4 VTAIL.n3 1.57809
R39 VTAIL.n6 VTAIL.n5 1.57809
R40 VTAIL.n2 VTAIL.n1 1.57809
R41 VTAIL VTAIL.n0 0.847483
R42 VTAIL VTAIL.n7 0.731103
R43 VTAIL.n5 VTAIL.n4 0.470328
R44 VTAIL.n1 VTAIL.n0 0.470328
R45 B.n350 B.n349 585
R46 B.n351 B.n350 585
R47 B.n121 B.n62 585
R48 B.n120 B.n119 585
R49 B.n118 B.n117 585
R50 B.n116 B.n115 585
R51 B.n114 B.n113 585
R52 B.n112 B.n111 585
R53 B.n110 B.n109 585
R54 B.n108 B.n107 585
R55 B.n106 B.n105 585
R56 B.n103 B.n102 585
R57 B.n101 B.n100 585
R58 B.n99 B.n98 585
R59 B.n97 B.n96 585
R60 B.n95 B.n94 585
R61 B.n93 B.n92 585
R62 B.n91 B.n90 585
R63 B.n89 B.n88 585
R64 B.n87 B.n86 585
R65 B.n85 B.n84 585
R66 B.n83 B.n82 585
R67 B.n81 B.n80 585
R68 B.n79 B.n78 585
R69 B.n77 B.n76 585
R70 B.n75 B.n74 585
R71 B.n73 B.n72 585
R72 B.n71 B.n70 585
R73 B.n69 B.n68 585
R74 B.n46 B.n45 585
R75 B.n348 B.n47 585
R76 B.n352 B.n47 585
R77 B.n347 B.n346 585
R78 B.n346 B.n43 585
R79 B.n345 B.n42 585
R80 B.n358 B.n42 585
R81 B.n344 B.n41 585
R82 B.n359 B.n41 585
R83 B.n343 B.n40 585
R84 B.n360 B.n40 585
R85 B.n342 B.n341 585
R86 B.n341 B.n39 585
R87 B.n340 B.n35 585
R88 B.n366 B.n35 585
R89 B.n339 B.n34 585
R90 B.n367 B.n34 585
R91 B.n338 B.n33 585
R92 B.n368 B.n33 585
R93 B.n337 B.n336 585
R94 B.n336 B.n29 585
R95 B.n335 B.n28 585
R96 B.n374 B.n28 585
R97 B.n334 B.n27 585
R98 B.n375 B.n27 585
R99 B.n333 B.n26 585
R100 B.n376 B.n26 585
R101 B.n332 B.n331 585
R102 B.n331 B.n22 585
R103 B.n330 B.n21 585
R104 B.n382 B.n21 585
R105 B.n329 B.n20 585
R106 B.n383 B.n20 585
R107 B.n328 B.n19 585
R108 B.n384 B.n19 585
R109 B.n327 B.n326 585
R110 B.n326 B.n15 585
R111 B.n325 B.n14 585
R112 B.n390 B.n14 585
R113 B.n324 B.n13 585
R114 B.n391 B.n13 585
R115 B.n323 B.n12 585
R116 B.n392 B.n12 585
R117 B.n322 B.n321 585
R118 B.n321 B.n8 585
R119 B.n320 B.n7 585
R120 B.n398 B.n7 585
R121 B.n319 B.n6 585
R122 B.n399 B.n6 585
R123 B.n318 B.n5 585
R124 B.n400 B.n5 585
R125 B.n317 B.n316 585
R126 B.n316 B.n4 585
R127 B.n315 B.n122 585
R128 B.n315 B.n314 585
R129 B.n305 B.n123 585
R130 B.n124 B.n123 585
R131 B.n307 B.n306 585
R132 B.n308 B.n307 585
R133 B.n304 B.n128 585
R134 B.n132 B.n128 585
R135 B.n303 B.n302 585
R136 B.n302 B.n301 585
R137 B.n130 B.n129 585
R138 B.n131 B.n130 585
R139 B.n294 B.n293 585
R140 B.n295 B.n294 585
R141 B.n292 B.n137 585
R142 B.n137 B.n136 585
R143 B.n291 B.n290 585
R144 B.n290 B.n289 585
R145 B.n139 B.n138 585
R146 B.n140 B.n139 585
R147 B.n282 B.n281 585
R148 B.n283 B.n282 585
R149 B.n280 B.n145 585
R150 B.n145 B.n144 585
R151 B.n279 B.n278 585
R152 B.n278 B.n277 585
R153 B.n147 B.n146 585
R154 B.n148 B.n147 585
R155 B.n270 B.n269 585
R156 B.n271 B.n270 585
R157 B.n268 B.n153 585
R158 B.n153 B.n152 585
R159 B.n267 B.n266 585
R160 B.n266 B.n265 585
R161 B.n155 B.n154 585
R162 B.n258 B.n155 585
R163 B.n257 B.n256 585
R164 B.n259 B.n257 585
R165 B.n255 B.n160 585
R166 B.n160 B.n159 585
R167 B.n254 B.n253 585
R168 B.n253 B.n252 585
R169 B.n162 B.n161 585
R170 B.n163 B.n162 585
R171 B.n245 B.n244 585
R172 B.n246 B.n245 585
R173 B.n166 B.n165 585
R174 B.n187 B.n185 585
R175 B.n188 B.n184 585
R176 B.n188 B.n167 585
R177 B.n191 B.n190 585
R178 B.n192 B.n183 585
R179 B.n194 B.n193 585
R180 B.n196 B.n182 585
R181 B.n199 B.n198 585
R182 B.n200 B.n181 585
R183 B.n205 B.n204 585
R184 B.n207 B.n180 585
R185 B.n210 B.n209 585
R186 B.n211 B.n179 585
R187 B.n213 B.n212 585
R188 B.n215 B.n178 585
R189 B.n218 B.n217 585
R190 B.n219 B.n177 585
R191 B.n221 B.n220 585
R192 B.n223 B.n176 585
R193 B.n226 B.n225 585
R194 B.n227 B.n172 585
R195 B.n229 B.n228 585
R196 B.n231 B.n171 585
R197 B.n234 B.n233 585
R198 B.n235 B.n170 585
R199 B.n237 B.n236 585
R200 B.n239 B.n169 585
R201 B.n242 B.n241 585
R202 B.n243 B.n168 585
R203 B.n248 B.n247 585
R204 B.n247 B.n246 585
R205 B.n249 B.n164 585
R206 B.n164 B.n163 585
R207 B.n251 B.n250 585
R208 B.n252 B.n251 585
R209 B.n158 B.n157 585
R210 B.n159 B.n158 585
R211 B.n261 B.n260 585
R212 B.n260 B.n259 585
R213 B.n262 B.n156 585
R214 B.n258 B.n156 585
R215 B.n264 B.n263 585
R216 B.n265 B.n264 585
R217 B.n151 B.n150 585
R218 B.n152 B.n151 585
R219 B.n273 B.n272 585
R220 B.n272 B.n271 585
R221 B.n274 B.n149 585
R222 B.n149 B.n148 585
R223 B.n276 B.n275 585
R224 B.n277 B.n276 585
R225 B.n143 B.n142 585
R226 B.n144 B.n143 585
R227 B.n285 B.n284 585
R228 B.n284 B.n283 585
R229 B.n286 B.n141 585
R230 B.n141 B.n140 585
R231 B.n288 B.n287 585
R232 B.n289 B.n288 585
R233 B.n135 B.n134 585
R234 B.n136 B.n135 585
R235 B.n297 B.n296 585
R236 B.n296 B.n295 585
R237 B.n298 B.n133 585
R238 B.n133 B.n131 585
R239 B.n300 B.n299 585
R240 B.n301 B.n300 585
R241 B.n127 B.n126 585
R242 B.n132 B.n127 585
R243 B.n310 B.n309 585
R244 B.n309 B.n308 585
R245 B.n311 B.n125 585
R246 B.n125 B.n124 585
R247 B.n313 B.n312 585
R248 B.n314 B.n313 585
R249 B.n2 B.n0 585
R250 B.n4 B.n2 585
R251 B.n3 B.n1 585
R252 B.n399 B.n3 585
R253 B.n397 B.n396 585
R254 B.n398 B.n397 585
R255 B.n395 B.n9 585
R256 B.n9 B.n8 585
R257 B.n394 B.n393 585
R258 B.n393 B.n392 585
R259 B.n11 B.n10 585
R260 B.n391 B.n11 585
R261 B.n389 B.n388 585
R262 B.n390 B.n389 585
R263 B.n387 B.n16 585
R264 B.n16 B.n15 585
R265 B.n386 B.n385 585
R266 B.n385 B.n384 585
R267 B.n18 B.n17 585
R268 B.n383 B.n18 585
R269 B.n381 B.n380 585
R270 B.n382 B.n381 585
R271 B.n379 B.n23 585
R272 B.n23 B.n22 585
R273 B.n378 B.n377 585
R274 B.n377 B.n376 585
R275 B.n25 B.n24 585
R276 B.n375 B.n25 585
R277 B.n373 B.n372 585
R278 B.n374 B.n373 585
R279 B.n371 B.n30 585
R280 B.n30 B.n29 585
R281 B.n370 B.n369 585
R282 B.n369 B.n368 585
R283 B.n32 B.n31 585
R284 B.n367 B.n32 585
R285 B.n365 B.n364 585
R286 B.n366 B.n365 585
R287 B.n363 B.n36 585
R288 B.n39 B.n36 585
R289 B.n362 B.n361 585
R290 B.n361 B.n360 585
R291 B.n38 B.n37 585
R292 B.n359 B.n38 585
R293 B.n357 B.n356 585
R294 B.n358 B.n357 585
R295 B.n355 B.n44 585
R296 B.n44 B.n43 585
R297 B.n354 B.n353 585
R298 B.n353 B.n352 585
R299 B.n402 B.n401 585
R300 B.n401 B.n400 585
R301 B.n247 B.n166 521.33
R302 B.n353 B.n46 521.33
R303 B.n245 B.n168 521.33
R304 B.n350 B.n47 521.33
R305 B.n351 B.n61 256.663
R306 B.n351 B.n60 256.663
R307 B.n351 B.n59 256.663
R308 B.n351 B.n58 256.663
R309 B.n351 B.n57 256.663
R310 B.n351 B.n56 256.663
R311 B.n351 B.n55 256.663
R312 B.n351 B.n54 256.663
R313 B.n351 B.n53 256.663
R314 B.n351 B.n52 256.663
R315 B.n351 B.n51 256.663
R316 B.n351 B.n50 256.663
R317 B.n351 B.n49 256.663
R318 B.n351 B.n48 256.663
R319 B.n186 B.n167 256.663
R320 B.n189 B.n167 256.663
R321 B.n195 B.n167 256.663
R322 B.n197 B.n167 256.663
R323 B.n206 B.n167 256.663
R324 B.n208 B.n167 256.663
R325 B.n214 B.n167 256.663
R326 B.n216 B.n167 256.663
R327 B.n222 B.n167 256.663
R328 B.n224 B.n167 256.663
R329 B.n230 B.n167 256.663
R330 B.n232 B.n167 256.663
R331 B.n238 B.n167 256.663
R332 B.n240 B.n167 256.663
R333 B.n246 B.n167 242.913
R334 B.n352 B.n351 242.913
R335 B.n173 B.t8 223.274
R336 B.n201 B.t4 223.274
R337 B.n65 B.t11 223.274
R338 B.n63 B.t15 223.274
R339 B.n201 B.t7 181.984
R340 B.n65 B.t13 181.984
R341 B.n173 B.t10 181.984
R342 B.n63 B.t16 181.984
R343 B.n247 B.n164 163.367
R344 B.n251 B.n164 163.367
R345 B.n251 B.n158 163.367
R346 B.n260 B.n158 163.367
R347 B.n260 B.n156 163.367
R348 B.n264 B.n156 163.367
R349 B.n264 B.n151 163.367
R350 B.n272 B.n151 163.367
R351 B.n272 B.n149 163.367
R352 B.n276 B.n149 163.367
R353 B.n276 B.n143 163.367
R354 B.n284 B.n143 163.367
R355 B.n284 B.n141 163.367
R356 B.n288 B.n141 163.367
R357 B.n288 B.n135 163.367
R358 B.n296 B.n135 163.367
R359 B.n296 B.n133 163.367
R360 B.n300 B.n133 163.367
R361 B.n300 B.n127 163.367
R362 B.n309 B.n127 163.367
R363 B.n309 B.n125 163.367
R364 B.n313 B.n125 163.367
R365 B.n313 B.n2 163.367
R366 B.n401 B.n2 163.367
R367 B.n401 B.n3 163.367
R368 B.n397 B.n3 163.367
R369 B.n397 B.n9 163.367
R370 B.n393 B.n9 163.367
R371 B.n393 B.n11 163.367
R372 B.n389 B.n11 163.367
R373 B.n389 B.n16 163.367
R374 B.n385 B.n16 163.367
R375 B.n385 B.n18 163.367
R376 B.n381 B.n18 163.367
R377 B.n381 B.n23 163.367
R378 B.n377 B.n23 163.367
R379 B.n377 B.n25 163.367
R380 B.n373 B.n25 163.367
R381 B.n373 B.n30 163.367
R382 B.n369 B.n30 163.367
R383 B.n369 B.n32 163.367
R384 B.n365 B.n32 163.367
R385 B.n365 B.n36 163.367
R386 B.n361 B.n36 163.367
R387 B.n361 B.n38 163.367
R388 B.n357 B.n38 163.367
R389 B.n357 B.n44 163.367
R390 B.n353 B.n44 163.367
R391 B.n188 B.n187 163.367
R392 B.n190 B.n188 163.367
R393 B.n194 B.n183 163.367
R394 B.n198 B.n196 163.367
R395 B.n205 B.n181 163.367
R396 B.n209 B.n207 163.367
R397 B.n213 B.n179 163.367
R398 B.n217 B.n215 163.367
R399 B.n221 B.n177 163.367
R400 B.n225 B.n223 163.367
R401 B.n229 B.n172 163.367
R402 B.n233 B.n231 163.367
R403 B.n237 B.n170 163.367
R404 B.n241 B.n239 163.367
R405 B.n245 B.n162 163.367
R406 B.n253 B.n162 163.367
R407 B.n253 B.n160 163.367
R408 B.n257 B.n160 163.367
R409 B.n257 B.n155 163.367
R410 B.n266 B.n155 163.367
R411 B.n266 B.n153 163.367
R412 B.n270 B.n153 163.367
R413 B.n270 B.n147 163.367
R414 B.n278 B.n147 163.367
R415 B.n278 B.n145 163.367
R416 B.n282 B.n145 163.367
R417 B.n282 B.n139 163.367
R418 B.n290 B.n139 163.367
R419 B.n290 B.n137 163.367
R420 B.n294 B.n137 163.367
R421 B.n294 B.n130 163.367
R422 B.n302 B.n130 163.367
R423 B.n302 B.n128 163.367
R424 B.n307 B.n128 163.367
R425 B.n307 B.n123 163.367
R426 B.n315 B.n123 163.367
R427 B.n316 B.n315 163.367
R428 B.n316 B.n5 163.367
R429 B.n6 B.n5 163.367
R430 B.n7 B.n6 163.367
R431 B.n321 B.n7 163.367
R432 B.n321 B.n12 163.367
R433 B.n13 B.n12 163.367
R434 B.n14 B.n13 163.367
R435 B.n326 B.n14 163.367
R436 B.n326 B.n19 163.367
R437 B.n20 B.n19 163.367
R438 B.n21 B.n20 163.367
R439 B.n331 B.n21 163.367
R440 B.n331 B.n26 163.367
R441 B.n27 B.n26 163.367
R442 B.n28 B.n27 163.367
R443 B.n336 B.n28 163.367
R444 B.n336 B.n33 163.367
R445 B.n34 B.n33 163.367
R446 B.n35 B.n34 163.367
R447 B.n341 B.n35 163.367
R448 B.n341 B.n40 163.367
R449 B.n41 B.n40 163.367
R450 B.n42 B.n41 163.367
R451 B.n346 B.n42 163.367
R452 B.n346 B.n47 163.367
R453 B.n70 B.n69 163.367
R454 B.n74 B.n73 163.367
R455 B.n78 B.n77 163.367
R456 B.n82 B.n81 163.367
R457 B.n86 B.n85 163.367
R458 B.n90 B.n89 163.367
R459 B.n94 B.n93 163.367
R460 B.n98 B.n97 163.367
R461 B.n102 B.n101 163.367
R462 B.n107 B.n106 163.367
R463 B.n111 B.n110 163.367
R464 B.n115 B.n114 163.367
R465 B.n119 B.n118 163.367
R466 B.n350 B.n62 163.367
R467 B.n174 B.t9 146.494
R468 B.n202 B.t6 146.494
R469 B.n66 B.t14 146.494
R470 B.n64 B.t17 146.494
R471 B.n246 B.n163 117.15
R472 B.n252 B.n163 117.15
R473 B.n252 B.n159 117.15
R474 B.n259 B.n159 117.15
R475 B.n259 B.n258 117.15
R476 B.n265 B.n152 117.15
R477 B.n271 B.n152 117.15
R478 B.n271 B.n148 117.15
R479 B.n277 B.n148 117.15
R480 B.n277 B.n144 117.15
R481 B.n283 B.n144 117.15
R482 B.n283 B.n140 117.15
R483 B.n289 B.n140 117.15
R484 B.n295 B.n136 117.15
R485 B.n295 B.n131 117.15
R486 B.n301 B.n131 117.15
R487 B.n301 B.n132 117.15
R488 B.n308 B.n124 117.15
R489 B.n314 B.n124 117.15
R490 B.n314 B.n4 117.15
R491 B.n400 B.n4 117.15
R492 B.n400 B.n399 117.15
R493 B.n399 B.n398 117.15
R494 B.n398 B.n8 117.15
R495 B.n392 B.n8 117.15
R496 B.n391 B.n390 117.15
R497 B.n390 B.n15 117.15
R498 B.n384 B.n15 117.15
R499 B.n384 B.n383 117.15
R500 B.n382 B.n22 117.15
R501 B.n376 B.n22 117.15
R502 B.n376 B.n375 117.15
R503 B.n375 B.n374 117.15
R504 B.n374 B.n29 117.15
R505 B.n368 B.n29 117.15
R506 B.n368 B.n367 117.15
R507 B.n367 B.n366 117.15
R508 B.n360 B.n39 117.15
R509 B.n360 B.n359 117.15
R510 B.n359 B.n358 117.15
R511 B.n358 B.n43 117.15
R512 B.n352 B.n43 117.15
R513 B.n258 B.t5 86.1399
R514 B.n39 B.t12 86.1399
R515 B.n132 B.t2 82.6943
R516 B.t1 B.n391 82.6943
R517 B.t3 B.n136 79.2487
R518 B.n383 B.t0 79.2487
R519 B.n186 B.n166 71.676
R520 B.n190 B.n189 71.676
R521 B.n195 B.n194 71.676
R522 B.n198 B.n197 71.676
R523 B.n206 B.n205 71.676
R524 B.n209 B.n208 71.676
R525 B.n214 B.n213 71.676
R526 B.n217 B.n216 71.676
R527 B.n222 B.n221 71.676
R528 B.n225 B.n224 71.676
R529 B.n230 B.n229 71.676
R530 B.n233 B.n232 71.676
R531 B.n238 B.n237 71.676
R532 B.n241 B.n240 71.676
R533 B.n48 B.n46 71.676
R534 B.n70 B.n49 71.676
R535 B.n74 B.n50 71.676
R536 B.n78 B.n51 71.676
R537 B.n82 B.n52 71.676
R538 B.n86 B.n53 71.676
R539 B.n90 B.n54 71.676
R540 B.n94 B.n55 71.676
R541 B.n98 B.n56 71.676
R542 B.n102 B.n57 71.676
R543 B.n107 B.n58 71.676
R544 B.n111 B.n59 71.676
R545 B.n115 B.n60 71.676
R546 B.n119 B.n61 71.676
R547 B.n62 B.n61 71.676
R548 B.n118 B.n60 71.676
R549 B.n114 B.n59 71.676
R550 B.n110 B.n58 71.676
R551 B.n106 B.n57 71.676
R552 B.n101 B.n56 71.676
R553 B.n97 B.n55 71.676
R554 B.n93 B.n54 71.676
R555 B.n89 B.n53 71.676
R556 B.n85 B.n52 71.676
R557 B.n81 B.n51 71.676
R558 B.n77 B.n50 71.676
R559 B.n73 B.n49 71.676
R560 B.n69 B.n48 71.676
R561 B.n187 B.n186 71.676
R562 B.n189 B.n183 71.676
R563 B.n196 B.n195 71.676
R564 B.n197 B.n181 71.676
R565 B.n207 B.n206 71.676
R566 B.n208 B.n179 71.676
R567 B.n215 B.n214 71.676
R568 B.n216 B.n177 71.676
R569 B.n223 B.n222 71.676
R570 B.n224 B.n172 71.676
R571 B.n231 B.n230 71.676
R572 B.n232 B.n170 71.676
R573 B.n239 B.n238 71.676
R574 B.n240 B.n168 71.676
R575 B.n175 B.n174 59.5399
R576 B.n203 B.n202 59.5399
R577 B.n67 B.n66 59.5399
R578 B.n104 B.n64 59.5399
R579 B.n289 B.t3 37.9018
R580 B.t0 B.n382 37.9018
R581 B.n174 B.n173 35.4914
R582 B.n202 B.n201 35.4914
R583 B.n66 B.n65 35.4914
R584 B.n64 B.n63 35.4914
R585 B.n308 B.t2 34.4563
R586 B.n392 B.t1 34.4563
R587 B.n354 B.n45 33.8737
R588 B.n349 B.n348 33.8737
R589 B.n244 B.n243 33.8737
R590 B.n248 B.n165 33.8737
R591 B.n265 B.t5 31.0107
R592 B.n366 B.t12 31.0107
R593 B B.n402 18.0485
R594 B.n68 B.n45 10.6151
R595 B.n71 B.n68 10.6151
R596 B.n72 B.n71 10.6151
R597 B.n75 B.n72 10.6151
R598 B.n76 B.n75 10.6151
R599 B.n79 B.n76 10.6151
R600 B.n80 B.n79 10.6151
R601 B.n83 B.n80 10.6151
R602 B.n84 B.n83 10.6151
R603 B.n88 B.n87 10.6151
R604 B.n91 B.n88 10.6151
R605 B.n92 B.n91 10.6151
R606 B.n95 B.n92 10.6151
R607 B.n96 B.n95 10.6151
R608 B.n99 B.n96 10.6151
R609 B.n100 B.n99 10.6151
R610 B.n103 B.n100 10.6151
R611 B.n108 B.n105 10.6151
R612 B.n109 B.n108 10.6151
R613 B.n112 B.n109 10.6151
R614 B.n113 B.n112 10.6151
R615 B.n116 B.n113 10.6151
R616 B.n117 B.n116 10.6151
R617 B.n120 B.n117 10.6151
R618 B.n121 B.n120 10.6151
R619 B.n349 B.n121 10.6151
R620 B.n244 B.n161 10.6151
R621 B.n254 B.n161 10.6151
R622 B.n255 B.n254 10.6151
R623 B.n256 B.n255 10.6151
R624 B.n256 B.n154 10.6151
R625 B.n267 B.n154 10.6151
R626 B.n268 B.n267 10.6151
R627 B.n269 B.n268 10.6151
R628 B.n269 B.n146 10.6151
R629 B.n279 B.n146 10.6151
R630 B.n280 B.n279 10.6151
R631 B.n281 B.n280 10.6151
R632 B.n281 B.n138 10.6151
R633 B.n291 B.n138 10.6151
R634 B.n292 B.n291 10.6151
R635 B.n293 B.n292 10.6151
R636 B.n293 B.n129 10.6151
R637 B.n303 B.n129 10.6151
R638 B.n304 B.n303 10.6151
R639 B.n306 B.n304 10.6151
R640 B.n306 B.n305 10.6151
R641 B.n305 B.n122 10.6151
R642 B.n317 B.n122 10.6151
R643 B.n318 B.n317 10.6151
R644 B.n319 B.n318 10.6151
R645 B.n320 B.n319 10.6151
R646 B.n322 B.n320 10.6151
R647 B.n323 B.n322 10.6151
R648 B.n324 B.n323 10.6151
R649 B.n325 B.n324 10.6151
R650 B.n327 B.n325 10.6151
R651 B.n328 B.n327 10.6151
R652 B.n329 B.n328 10.6151
R653 B.n330 B.n329 10.6151
R654 B.n332 B.n330 10.6151
R655 B.n333 B.n332 10.6151
R656 B.n334 B.n333 10.6151
R657 B.n335 B.n334 10.6151
R658 B.n337 B.n335 10.6151
R659 B.n338 B.n337 10.6151
R660 B.n339 B.n338 10.6151
R661 B.n340 B.n339 10.6151
R662 B.n342 B.n340 10.6151
R663 B.n343 B.n342 10.6151
R664 B.n344 B.n343 10.6151
R665 B.n345 B.n344 10.6151
R666 B.n347 B.n345 10.6151
R667 B.n348 B.n347 10.6151
R668 B.n185 B.n165 10.6151
R669 B.n185 B.n184 10.6151
R670 B.n191 B.n184 10.6151
R671 B.n192 B.n191 10.6151
R672 B.n193 B.n192 10.6151
R673 B.n193 B.n182 10.6151
R674 B.n199 B.n182 10.6151
R675 B.n200 B.n199 10.6151
R676 B.n204 B.n200 10.6151
R677 B.n210 B.n180 10.6151
R678 B.n211 B.n210 10.6151
R679 B.n212 B.n211 10.6151
R680 B.n212 B.n178 10.6151
R681 B.n218 B.n178 10.6151
R682 B.n219 B.n218 10.6151
R683 B.n220 B.n219 10.6151
R684 B.n220 B.n176 10.6151
R685 B.n227 B.n226 10.6151
R686 B.n228 B.n227 10.6151
R687 B.n228 B.n171 10.6151
R688 B.n234 B.n171 10.6151
R689 B.n235 B.n234 10.6151
R690 B.n236 B.n235 10.6151
R691 B.n236 B.n169 10.6151
R692 B.n242 B.n169 10.6151
R693 B.n243 B.n242 10.6151
R694 B.n249 B.n248 10.6151
R695 B.n250 B.n249 10.6151
R696 B.n250 B.n157 10.6151
R697 B.n261 B.n157 10.6151
R698 B.n262 B.n261 10.6151
R699 B.n263 B.n262 10.6151
R700 B.n263 B.n150 10.6151
R701 B.n273 B.n150 10.6151
R702 B.n274 B.n273 10.6151
R703 B.n275 B.n274 10.6151
R704 B.n275 B.n142 10.6151
R705 B.n285 B.n142 10.6151
R706 B.n286 B.n285 10.6151
R707 B.n287 B.n286 10.6151
R708 B.n287 B.n134 10.6151
R709 B.n297 B.n134 10.6151
R710 B.n298 B.n297 10.6151
R711 B.n299 B.n298 10.6151
R712 B.n299 B.n126 10.6151
R713 B.n310 B.n126 10.6151
R714 B.n311 B.n310 10.6151
R715 B.n312 B.n311 10.6151
R716 B.n312 B.n0 10.6151
R717 B.n396 B.n1 10.6151
R718 B.n396 B.n395 10.6151
R719 B.n395 B.n394 10.6151
R720 B.n394 B.n10 10.6151
R721 B.n388 B.n10 10.6151
R722 B.n388 B.n387 10.6151
R723 B.n387 B.n386 10.6151
R724 B.n386 B.n17 10.6151
R725 B.n380 B.n17 10.6151
R726 B.n380 B.n379 10.6151
R727 B.n379 B.n378 10.6151
R728 B.n378 B.n24 10.6151
R729 B.n372 B.n24 10.6151
R730 B.n372 B.n371 10.6151
R731 B.n371 B.n370 10.6151
R732 B.n370 B.n31 10.6151
R733 B.n364 B.n31 10.6151
R734 B.n364 B.n363 10.6151
R735 B.n363 B.n362 10.6151
R736 B.n362 B.n37 10.6151
R737 B.n356 B.n37 10.6151
R738 B.n356 B.n355 10.6151
R739 B.n355 B.n354 10.6151
R740 B.n87 B.n67 6.5566
R741 B.n104 B.n103 6.5566
R742 B.n203 B.n180 6.5566
R743 B.n176 B.n175 6.5566
R744 B.n84 B.n67 4.05904
R745 B.n105 B.n104 4.05904
R746 B.n204 B.n203 4.05904
R747 B.n226 B.n175 4.05904
R748 B.n402 B.n0 2.81026
R749 B.n402 B.n1 2.81026
R750 VN.n0 VN.t3 54.1947
R751 VN.n1 VN.t2 54.1947
R752 VN.n0 VN.t0 53.8783
R753 VN.n1 VN.t1 53.8783
R754 VN VN.n1 48.0152
R755 VN VN.n0 13.0644
R756 VDD2.n2 VDD2.n0 175.837
R757 VDD2.n2 VDD2.n1 146.433
R758 VDD2.n1 VDD2.t2 17.8383
R759 VDD2.n1 VDD2.t1 17.8383
R760 VDD2.n0 VDD2.t0 17.8383
R761 VDD2.n0 VDD2.t3 17.8383
R762 VDD2 VDD2.n2 0.0586897
C0 VDD2 VTAIL 2.29856f
C1 VP VTAIL 1.07235f
C2 VP VDD2 0.332437f
C3 VDD1 VN 0.154969f
C4 VN VTAIL 1.05824f
C5 VDD1 VTAIL 2.25173f
C6 VN VDD2 0.666079f
C7 VDD1 VDD2 0.760223f
C8 VP VN 3.39138f
C9 VDD1 VP 0.841798f
C10 VDD2 B 2.263277f
C11 VDD1 B 4.28432f
C12 VTAIL B 2.667789f
C13 VN B 7.13941f
C14 VP B 5.637148f
C15 VDD2.t0 B 0.018938f
C16 VDD2.t3 B 0.018938f
C17 VDD2.n0 B 0.212517f
C18 VDD2.t2 B 0.018938f
C19 VDD2.t1 B 0.018938f
C20 VDD2.n1 B 0.097039f
C21 VDD2.n2 B 1.8003f
C22 VN.t3 B 0.227898f
C23 VN.t0 B 0.226816f
C24 VN.n0 B 0.172265f
C25 VN.t2 B 0.227898f
C26 VN.t1 B 0.226816f
C27 VN.n1 B 0.942139f
C28 VTAIL.t7 B 0.103889f
C29 VTAIL.n0 B 0.220698f
C30 VTAIL.t3 B 0.103889f
C31 VTAIL.n1 B 0.267963f
C32 VTAIL.t4 B 0.103889f
C33 VTAIL.n2 B 0.674258f
C34 VTAIL.t5 B 0.103889f
C35 VTAIL.n3 B 0.674258f
C36 VTAIL.t6 B 0.103889f
C37 VTAIL.n4 B 0.267963f
C38 VTAIL.t1 B 0.103889f
C39 VTAIL.n5 B 0.267963f
C40 VTAIL.t2 B 0.103889f
C41 VTAIL.n6 B 0.674258f
C42 VTAIL.t0 B 0.103889f
C43 VTAIL.n7 B 0.619464f
C44 VDD1.t2 B 0.018303f
C45 VDD1.t0 B 0.018303f
C46 VDD1.n0 B 0.093887f
C47 VDD1.t3 B 0.018303f
C48 VDD1.t1 B 0.018303f
C49 VDD1.n1 B 0.214321f
C50 VP.n0 B 0.030288f
C51 VP.t1 B 0.098886f
C52 VP.n1 B 0.044215f
C53 VP.t3 B 0.230752f
C54 VP.t2 B 0.229656f
C55 VP.n2 B 0.936975f
C56 VP.n3 B 1.20808f
C57 VP.t0 B 0.098886f
C58 VP.n4 B 0.134563f
C59 VP.n5 B 0.037775f
C60 VP.n6 B 0.030288f
C61 VP.n7 B 0.030288f
C62 VP.n8 B 0.030288f
C63 VP.n9 B 0.044215f
C64 VP.n10 B 0.037775f
C65 VP.n11 B 0.134563f
C66 VP.n12 B 0.029528f
.ends

