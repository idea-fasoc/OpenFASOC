* NGSPICE file created from diff_pair_sample_0647.ext - technology: sky130A

.subckt diff_pair_sample_0647 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 w_n2614_n4262# sky130_fd_pr__pfet_01v8 ad=6.4233 pd=33.72 as=6.4233 ps=33.72 w=16.47 l=3.78
X1 B.t11 B.t9 B.t10 w_n2614_n4262# sky130_fd_pr__pfet_01v8 ad=6.4233 pd=33.72 as=0 ps=0 w=16.47 l=3.78
X2 VDD2.t1 VN.t0 VTAIL.t0 w_n2614_n4262# sky130_fd_pr__pfet_01v8 ad=6.4233 pd=33.72 as=6.4233 ps=33.72 w=16.47 l=3.78
X3 B.t8 B.t6 B.t7 w_n2614_n4262# sky130_fd_pr__pfet_01v8 ad=6.4233 pd=33.72 as=0 ps=0 w=16.47 l=3.78
X4 VDD2.t0 VN.t1 VTAIL.t1 w_n2614_n4262# sky130_fd_pr__pfet_01v8 ad=6.4233 pd=33.72 as=6.4233 ps=33.72 w=16.47 l=3.78
X5 B.t5 B.t3 B.t4 w_n2614_n4262# sky130_fd_pr__pfet_01v8 ad=6.4233 pd=33.72 as=0 ps=0 w=16.47 l=3.78
X6 VDD1.t0 VP.t1 VTAIL.t2 w_n2614_n4262# sky130_fd_pr__pfet_01v8 ad=6.4233 pd=33.72 as=6.4233 ps=33.72 w=16.47 l=3.78
X7 B.t2 B.t0 B.t1 w_n2614_n4262# sky130_fd_pr__pfet_01v8 ad=6.4233 pd=33.72 as=0 ps=0 w=16.47 l=3.78
R0 VP.n0 VP.t0 191.216
R1 VP.n0 VP.t1 140.044
R2 VP VP.n0 0.621237
R3 VTAIL.n1 VTAIL.t0 55.4681
R4 VTAIL.n3 VTAIL.t1 55.4678
R5 VTAIL.n0 VTAIL.t2 55.4678
R6 VTAIL.n2 VTAIL.t3 55.4678
R7 VTAIL.n1 VTAIL.n0 33.6514
R8 VTAIL.n3 VTAIL.n2 30.1083
R9 VTAIL.n2 VTAIL.n1 2.24188
R10 VTAIL VTAIL.n0 1.41429
R11 VTAIL VTAIL.n3 0.828086
R12 VDD1 VDD1.t0 118.501
R13 VDD1 VDD1.t1 73.0906
R14 B.n420 B.n115 585
R15 B.n419 B.n418 585
R16 B.n417 B.n116 585
R17 B.n416 B.n415 585
R18 B.n414 B.n117 585
R19 B.n413 B.n412 585
R20 B.n411 B.n118 585
R21 B.n410 B.n409 585
R22 B.n408 B.n119 585
R23 B.n407 B.n406 585
R24 B.n405 B.n120 585
R25 B.n404 B.n403 585
R26 B.n402 B.n121 585
R27 B.n401 B.n400 585
R28 B.n399 B.n122 585
R29 B.n398 B.n397 585
R30 B.n396 B.n123 585
R31 B.n395 B.n394 585
R32 B.n393 B.n124 585
R33 B.n392 B.n391 585
R34 B.n390 B.n125 585
R35 B.n389 B.n388 585
R36 B.n387 B.n126 585
R37 B.n386 B.n385 585
R38 B.n384 B.n127 585
R39 B.n383 B.n382 585
R40 B.n381 B.n128 585
R41 B.n380 B.n379 585
R42 B.n378 B.n129 585
R43 B.n377 B.n376 585
R44 B.n375 B.n130 585
R45 B.n374 B.n373 585
R46 B.n372 B.n131 585
R47 B.n371 B.n370 585
R48 B.n369 B.n132 585
R49 B.n368 B.n367 585
R50 B.n366 B.n133 585
R51 B.n365 B.n364 585
R52 B.n363 B.n134 585
R53 B.n362 B.n361 585
R54 B.n360 B.n135 585
R55 B.n359 B.n358 585
R56 B.n357 B.n136 585
R57 B.n356 B.n355 585
R58 B.n354 B.n137 585
R59 B.n353 B.n352 585
R60 B.n351 B.n138 585
R61 B.n350 B.n349 585
R62 B.n348 B.n139 585
R63 B.n347 B.n346 585
R64 B.n345 B.n140 585
R65 B.n344 B.n343 585
R66 B.n342 B.n141 585
R67 B.n341 B.n340 585
R68 B.n339 B.n142 585
R69 B.n338 B.n337 585
R70 B.n333 B.n143 585
R71 B.n332 B.n331 585
R72 B.n330 B.n144 585
R73 B.n329 B.n328 585
R74 B.n327 B.n145 585
R75 B.n326 B.n325 585
R76 B.n324 B.n146 585
R77 B.n323 B.n322 585
R78 B.n320 B.n147 585
R79 B.n319 B.n318 585
R80 B.n317 B.n150 585
R81 B.n316 B.n315 585
R82 B.n314 B.n151 585
R83 B.n313 B.n312 585
R84 B.n311 B.n152 585
R85 B.n310 B.n309 585
R86 B.n308 B.n153 585
R87 B.n307 B.n306 585
R88 B.n305 B.n154 585
R89 B.n304 B.n303 585
R90 B.n302 B.n155 585
R91 B.n301 B.n300 585
R92 B.n299 B.n156 585
R93 B.n298 B.n297 585
R94 B.n296 B.n157 585
R95 B.n295 B.n294 585
R96 B.n293 B.n158 585
R97 B.n292 B.n291 585
R98 B.n290 B.n159 585
R99 B.n289 B.n288 585
R100 B.n287 B.n160 585
R101 B.n286 B.n285 585
R102 B.n284 B.n161 585
R103 B.n283 B.n282 585
R104 B.n281 B.n162 585
R105 B.n280 B.n279 585
R106 B.n278 B.n163 585
R107 B.n277 B.n276 585
R108 B.n275 B.n164 585
R109 B.n274 B.n273 585
R110 B.n272 B.n165 585
R111 B.n271 B.n270 585
R112 B.n269 B.n166 585
R113 B.n268 B.n267 585
R114 B.n266 B.n167 585
R115 B.n265 B.n264 585
R116 B.n263 B.n168 585
R117 B.n262 B.n261 585
R118 B.n260 B.n169 585
R119 B.n259 B.n258 585
R120 B.n257 B.n170 585
R121 B.n256 B.n255 585
R122 B.n254 B.n171 585
R123 B.n253 B.n252 585
R124 B.n251 B.n172 585
R125 B.n250 B.n249 585
R126 B.n248 B.n173 585
R127 B.n247 B.n246 585
R128 B.n245 B.n174 585
R129 B.n244 B.n243 585
R130 B.n242 B.n175 585
R131 B.n241 B.n240 585
R132 B.n239 B.n176 585
R133 B.n422 B.n421 585
R134 B.n423 B.n114 585
R135 B.n425 B.n424 585
R136 B.n426 B.n113 585
R137 B.n428 B.n427 585
R138 B.n429 B.n112 585
R139 B.n431 B.n430 585
R140 B.n432 B.n111 585
R141 B.n434 B.n433 585
R142 B.n435 B.n110 585
R143 B.n437 B.n436 585
R144 B.n438 B.n109 585
R145 B.n440 B.n439 585
R146 B.n441 B.n108 585
R147 B.n443 B.n442 585
R148 B.n444 B.n107 585
R149 B.n446 B.n445 585
R150 B.n447 B.n106 585
R151 B.n449 B.n448 585
R152 B.n450 B.n105 585
R153 B.n452 B.n451 585
R154 B.n453 B.n104 585
R155 B.n455 B.n454 585
R156 B.n456 B.n103 585
R157 B.n458 B.n457 585
R158 B.n459 B.n102 585
R159 B.n461 B.n460 585
R160 B.n462 B.n101 585
R161 B.n464 B.n463 585
R162 B.n465 B.n100 585
R163 B.n467 B.n466 585
R164 B.n468 B.n99 585
R165 B.n470 B.n469 585
R166 B.n471 B.n98 585
R167 B.n473 B.n472 585
R168 B.n474 B.n97 585
R169 B.n476 B.n475 585
R170 B.n477 B.n96 585
R171 B.n479 B.n478 585
R172 B.n480 B.n95 585
R173 B.n482 B.n481 585
R174 B.n483 B.n94 585
R175 B.n485 B.n484 585
R176 B.n486 B.n93 585
R177 B.n488 B.n487 585
R178 B.n489 B.n92 585
R179 B.n491 B.n490 585
R180 B.n492 B.n91 585
R181 B.n494 B.n493 585
R182 B.n495 B.n90 585
R183 B.n497 B.n496 585
R184 B.n498 B.n89 585
R185 B.n500 B.n499 585
R186 B.n501 B.n88 585
R187 B.n503 B.n502 585
R188 B.n504 B.n87 585
R189 B.n506 B.n505 585
R190 B.n507 B.n86 585
R191 B.n509 B.n508 585
R192 B.n510 B.n85 585
R193 B.n512 B.n511 585
R194 B.n513 B.n84 585
R195 B.n515 B.n514 585
R196 B.n516 B.n83 585
R197 B.n518 B.n517 585
R198 B.n519 B.n82 585
R199 B.n699 B.n18 585
R200 B.n698 B.n697 585
R201 B.n696 B.n19 585
R202 B.n695 B.n694 585
R203 B.n693 B.n20 585
R204 B.n692 B.n691 585
R205 B.n690 B.n21 585
R206 B.n689 B.n688 585
R207 B.n687 B.n22 585
R208 B.n686 B.n685 585
R209 B.n684 B.n23 585
R210 B.n683 B.n682 585
R211 B.n681 B.n24 585
R212 B.n680 B.n679 585
R213 B.n678 B.n25 585
R214 B.n677 B.n676 585
R215 B.n675 B.n26 585
R216 B.n674 B.n673 585
R217 B.n672 B.n27 585
R218 B.n671 B.n670 585
R219 B.n669 B.n28 585
R220 B.n668 B.n667 585
R221 B.n666 B.n29 585
R222 B.n665 B.n664 585
R223 B.n663 B.n30 585
R224 B.n662 B.n661 585
R225 B.n660 B.n31 585
R226 B.n659 B.n658 585
R227 B.n657 B.n32 585
R228 B.n656 B.n655 585
R229 B.n654 B.n33 585
R230 B.n653 B.n652 585
R231 B.n651 B.n34 585
R232 B.n650 B.n649 585
R233 B.n648 B.n35 585
R234 B.n647 B.n646 585
R235 B.n645 B.n36 585
R236 B.n644 B.n643 585
R237 B.n642 B.n37 585
R238 B.n641 B.n640 585
R239 B.n639 B.n38 585
R240 B.n638 B.n637 585
R241 B.n636 B.n39 585
R242 B.n635 B.n634 585
R243 B.n633 B.n40 585
R244 B.n632 B.n631 585
R245 B.n630 B.n41 585
R246 B.n629 B.n628 585
R247 B.n627 B.n42 585
R248 B.n626 B.n625 585
R249 B.n624 B.n43 585
R250 B.n623 B.n622 585
R251 B.n621 B.n44 585
R252 B.n620 B.n619 585
R253 B.n618 B.n45 585
R254 B.n616 B.n615 585
R255 B.n614 B.n48 585
R256 B.n613 B.n612 585
R257 B.n611 B.n49 585
R258 B.n610 B.n609 585
R259 B.n608 B.n50 585
R260 B.n607 B.n606 585
R261 B.n605 B.n51 585
R262 B.n604 B.n603 585
R263 B.n602 B.n601 585
R264 B.n600 B.n55 585
R265 B.n599 B.n598 585
R266 B.n597 B.n56 585
R267 B.n596 B.n595 585
R268 B.n594 B.n57 585
R269 B.n593 B.n592 585
R270 B.n591 B.n58 585
R271 B.n590 B.n589 585
R272 B.n588 B.n59 585
R273 B.n587 B.n586 585
R274 B.n585 B.n60 585
R275 B.n584 B.n583 585
R276 B.n582 B.n61 585
R277 B.n581 B.n580 585
R278 B.n579 B.n62 585
R279 B.n578 B.n577 585
R280 B.n576 B.n63 585
R281 B.n575 B.n574 585
R282 B.n573 B.n64 585
R283 B.n572 B.n571 585
R284 B.n570 B.n65 585
R285 B.n569 B.n568 585
R286 B.n567 B.n66 585
R287 B.n566 B.n565 585
R288 B.n564 B.n67 585
R289 B.n563 B.n562 585
R290 B.n561 B.n68 585
R291 B.n560 B.n559 585
R292 B.n558 B.n69 585
R293 B.n557 B.n556 585
R294 B.n555 B.n70 585
R295 B.n554 B.n553 585
R296 B.n552 B.n71 585
R297 B.n551 B.n550 585
R298 B.n549 B.n72 585
R299 B.n548 B.n547 585
R300 B.n546 B.n73 585
R301 B.n545 B.n544 585
R302 B.n543 B.n74 585
R303 B.n542 B.n541 585
R304 B.n540 B.n75 585
R305 B.n539 B.n538 585
R306 B.n537 B.n76 585
R307 B.n536 B.n535 585
R308 B.n534 B.n77 585
R309 B.n533 B.n532 585
R310 B.n531 B.n78 585
R311 B.n530 B.n529 585
R312 B.n528 B.n79 585
R313 B.n527 B.n526 585
R314 B.n525 B.n80 585
R315 B.n524 B.n523 585
R316 B.n522 B.n81 585
R317 B.n521 B.n520 585
R318 B.n701 B.n700 585
R319 B.n702 B.n17 585
R320 B.n704 B.n703 585
R321 B.n705 B.n16 585
R322 B.n707 B.n706 585
R323 B.n708 B.n15 585
R324 B.n710 B.n709 585
R325 B.n711 B.n14 585
R326 B.n713 B.n712 585
R327 B.n714 B.n13 585
R328 B.n716 B.n715 585
R329 B.n717 B.n12 585
R330 B.n719 B.n718 585
R331 B.n720 B.n11 585
R332 B.n722 B.n721 585
R333 B.n723 B.n10 585
R334 B.n725 B.n724 585
R335 B.n726 B.n9 585
R336 B.n728 B.n727 585
R337 B.n729 B.n8 585
R338 B.n731 B.n730 585
R339 B.n732 B.n7 585
R340 B.n734 B.n733 585
R341 B.n735 B.n6 585
R342 B.n737 B.n736 585
R343 B.n738 B.n5 585
R344 B.n740 B.n739 585
R345 B.n741 B.n4 585
R346 B.n743 B.n742 585
R347 B.n744 B.n3 585
R348 B.n746 B.n745 585
R349 B.n747 B.n0 585
R350 B.n2 B.n1 585
R351 B.n193 B.n192 585
R352 B.n194 B.n191 585
R353 B.n196 B.n195 585
R354 B.n197 B.n190 585
R355 B.n199 B.n198 585
R356 B.n200 B.n189 585
R357 B.n202 B.n201 585
R358 B.n203 B.n188 585
R359 B.n205 B.n204 585
R360 B.n206 B.n187 585
R361 B.n208 B.n207 585
R362 B.n209 B.n186 585
R363 B.n211 B.n210 585
R364 B.n212 B.n185 585
R365 B.n214 B.n213 585
R366 B.n215 B.n184 585
R367 B.n217 B.n216 585
R368 B.n218 B.n183 585
R369 B.n220 B.n219 585
R370 B.n221 B.n182 585
R371 B.n223 B.n222 585
R372 B.n224 B.n181 585
R373 B.n226 B.n225 585
R374 B.n227 B.n180 585
R375 B.n229 B.n228 585
R376 B.n230 B.n179 585
R377 B.n232 B.n231 585
R378 B.n233 B.n178 585
R379 B.n235 B.n234 585
R380 B.n236 B.n177 585
R381 B.n238 B.n237 585
R382 B.n239 B.n238 473.281
R383 B.n422 B.n115 473.281
R384 B.n520 B.n519 473.281
R385 B.n700 B.n699 473.281
R386 B.n148 B.t9 314.336
R387 B.n334 B.t0 314.336
R388 B.n52 B.t3 314.336
R389 B.n46 B.t6 314.336
R390 B.n749 B.n748 256.663
R391 B.n748 B.n747 235.042
R392 B.n748 B.n2 235.042
R393 B.n334 B.t1 188.988
R394 B.n52 B.t5 188.988
R395 B.n148 B.t10 188.966
R396 B.n46 B.t8 188.966
R397 B.n240 B.n239 163.367
R398 B.n240 B.n175 163.367
R399 B.n244 B.n175 163.367
R400 B.n245 B.n244 163.367
R401 B.n246 B.n245 163.367
R402 B.n246 B.n173 163.367
R403 B.n250 B.n173 163.367
R404 B.n251 B.n250 163.367
R405 B.n252 B.n251 163.367
R406 B.n252 B.n171 163.367
R407 B.n256 B.n171 163.367
R408 B.n257 B.n256 163.367
R409 B.n258 B.n257 163.367
R410 B.n258 B.n169 163.367
R411 B.n262 B.n169 163.367
R412 B.n263 B.n262 163.367
R413 B.n264 B.n263 163.367
R414 B.n264 B.n167 163.367
R415 B.n268 B.n167 163.367
R416 B.n269 B.n268 163.367
R417 B.n270 B.n269 163.367
R418 B.n270 B.n165 163.367
R419 B.n274 B.n165 163.367
R420 B.n275 B.n274 163.367
R421 B.n276 B.n275 163.367
R422 B.n276 B.n163 163.367
R423 B.n280 B.n163 163.367
R424 B.n281 B.n280 163.367
R425 B.n282 B.n281 163.367
R426 B.n282 B.n161 163.367
R427 B.n286 B.n161 163.367
R428 B.n287 B.n286 163.367
R429 B.n288 B.n287 163.367
R430 B.n288 B.n159 163.367
R431 B.n292 B.n159 163.367
R432 B.n293 B.n292 163.367
R433 B.n294 B.n293 163.367
R434 B.n294 B.n157 163.367
R435 B.n298 B.n157 163.367
R436 B.n299 B.n298 163.367
R437 B.n300 B.n299 163.367
R438 B.n300 B.n155 163.367
R439 B.n304 B.n155 163.367
R440 B.n305 B.n304 163.367
R441 B.n306 B.n305 163.367
R442 B.n306 B.n153 163.367
R443 B.n310 B.n153 163.367
R444 B.n311 B.n310 163.367
R445 B.n312 B.n311 163.367
R446 B.n312 B.n151 163.367
R447 B.n316 B.n151 163.367
R448 B.n317 B.n316 163.367
R449 B.n318 B.n317 163.367
R450 B.n318 B.n147 163.367
R451 B.n323 B.n147 163.367
R452 B.n324 B.n323 163.367
R453 B.n325 B.n324 163.367
R454 B.n325 B.n145 163.367
R455 B.n329 B.n145 163.367
R456 B.n330 B.n329 163.367
R457 B.n331 B.n330 163.367
R458 B.n331 B.n143 163.367
R459 B.n338 B.n143 163.367
R460 B.n339 B.n338 163.367
R461 B.n340 B.n339 163.367
R462 B.n340 B.n141 163.367
R463 B.n344 B.n141 163.367
R464 B.n345 B.n344 163.367
R465 B.n346 B.n345 163.367
R466 B.n346 B.n139 163.367
R467 B.n350 B.n139 163.367
R468 B.n351 B.n350 163.367
R469 B.n352 B.n351 163.367
R470 B.n352 B.n137 163.367
R471 B.n356 B.n137 163.367
R472 B.n357 B.n356 163.367
R473 B.n358 B.n357 163.367
R474 B.n358 B.n135 163.367
R475 B.n362 B.n135 163.367
R476 B.n363 B.n362 163.367
R477 B.n364 B.n363 163.367
R478 B.n364 B.n133 163.367
R479 B.n368 B.n133 163.367
R480 B.n369 B.n368 163.367
R481 B.n370 B.n369 163.367
R482 B.n370 B.n131 163.367
R483 B.n374 B.n131 163.367
R484 B.n375 B.n374 163.367
R485 B.n376 B.n375 163.367
R486 B.n376 B.n129 163.367
R487 B.n380 B.n129 163.367
R488 B.n381 B.n380 163.367
R489 B.n382 B.n381 163.367
R490 B.n382 B.n127 163.367
R491 B.n386 B.n127 163.367
R492 B.n387 B.n386 163.367
R493 B.n388 B.n387 163.367
R494 B.n388 B.n125 163.367
R495 B.n392 B.n125 163.367
R496 B.n393 B.n392 163.367
R497 B.n394 B.n393 163.367
R498 B.n394 B.n123 163.367
R499 B.n398 B.n123 163.367
R500 B.n399 B.n398 163.367
R501 B.n400 B.n399 163.367
R502 B.n400 B.n121 163.367
R503 B.n404 B.n121 163.367
R504 B.n405 B.n404 163.367
R505 B.n406 B.n405 163.367
R506 B.n406 B.n119 163.367
R507 B.n410 B.n119 163.367
R508 B.n411 B.n410 163.367
R509 B.n412 B.n411 163.367
R510 B.n412 B.n117 163.367
R511 B.n416 B.n117 163.367
R512 B.n417 B.n416 163.367
R513 B.n418 B.n417 163.367
R514 B.n418 B.n115 163.367
R515 B.n519 B.n518 163.367
R516 B.n518 B.n83 163.367
R517 B.n514 B.n83 163.367
R518 B.n514 B.n513 163.367
R519 B.n513 B.n512 163.367
R520 B.n512 B.n85 163.367
R521 B.n508 B.n85 163.367
R522 B.n508 B.n507 163.367
R523 B.n507 B.n506 163.367
R524 B.n506 B.n87 163.367
R525 B.n502 B.n87 163.367
R526 B.n502 B.n501 163.367
R527 B.n501 B.n500 163.367
R528 B.n500 B.n89 163.367
R529 B.n496 B.n89 163.367
R530 B.n496 B.n495 163.367
R531 B.n495 B.n494 163.367
R532 B.n494 B.n91 163.367
R533 B.n490 B.n91 163.367
R534 B.n490 B.n489 163.367
R535 B.n489 B.n488 163.367
R536 B.n488 B.n93 163.367
R537 B.n484 B.n93 163.367
R538 B.n484 B.n483 163.367
R539 B.n483 B.n482 163.367
R540 B.n482 B.n95 163.367
R541 B.n478 B.n95 163.367
R542 B.n478 B.n477 163.367
R543 B.n477 B.n476 163.367
R544 B.n476 B.n97 163.367
R545 B.n472 B.n97 163.367
R546 B.n472 B.n471 163.367
R547 B.n471 B.n470 163.367
R548 B.n470 B.n99 163.367
R549 B.n466 B.n99 163.367
R550 B.n466 B.n465 163.367
R551 B.n465 B.n464 163.367
R552 B.n464 B.n101 163.367
R553 B.n460 B.n101 163.367
R554 B.n460 B.n459 163.367
R555 B.n459 B.n458 163.367
R556 B.n458 B.n103 163.367
R557 B.n454 B.n103 163.367
R558 B.n454 B.n453 163.367
R559 B.n453 B.n452 163.367
R560 B.n452 B.n105 163.367
R561 B.n448 B.n105 163.367
R562 B.n448 B.n447 163.367
R563 B.n447 B.n446 163.367
R564 B.n446 B.n107 163.367
R565 B.n442 B.n107 163.367
R566 B.n442 B.n441 163.367
R567 B.n441 B.n440 163.367
R568 B.n440 B.n109 163.367
R569 B.n436 B.n109 163.367
R570 B.n436 B.n435 163.367
R571 B.n435 B.n434 163.367
R572 B.n434 B.n111 163.367
R573 B.n430 B.n111 163.367
R574 B.n430 B.n429 163.367
R575 B.n429 B.n428 163.367
R576 B.n428 B.n113 163.367
R577 B.n424 B.n113 163.367
R578 B.n424 B.n423 163.367
R579 B.n423 B.n422 163.367
R580 B.n699 B.n698 163.367
R581 B.n698 B.n19 163.367
R582 B.n694 B.n19 163.367
R583 B.n694 B.n693 163.367
R584 B.n693 B.n692 163.367
R585 B.n692 B.n21 163.367
R586 B.n688 B.n21 163.367
R587 B.n688 B.n687 163.367
R588 B.n687 B.n686 163.367
R589 B.n686 B.n23 163.367
R590 B.n682 B.n23 163.367
R591 B.n682 B.n681 163.367
R592 B.n681 B.n680 163.367
R593 B.n680 B.n25 163.367
R594 B.n676 B.n25 163.367
R595 B.n676 B.n675 163.367
R596 B.n675 B.n674 163.367
R597 B.n674 B.n27 163.367
R598 B.n670 B.n27 163.367
R599 B.n670 B.n669 163.367
R600 B.n669 B.n668 163.367
R601 B.n668 B.n29 163.367
R602 B.n664 B.n29 163.367
R603 B.n664 B.n663 163.367
R604 B.n663 B.n662 163.367
R605 B.n662 B.n31 163.367
R606 B.n658 B.n31 163.367
R607 B.n658 B.n657 163.367
R608 B.n657 B.n656 163.367
R609 B.n656 B.n33 163.367
R610 B.n652 B.n33 163.367
R611 B.n652 B.n651 163.367
R612 B.n651 B.n650 163.367
R613 B.n650 B.n35 163.367
R614 B.n646 B.n35 163.367
R615 B.n646 B.n645 163.367
R616 B.n645 B.n644 163.367
R617 B.n644 B.n37 163.367
R618 B.n640 B.n37 163.367
R619 B.n640 B.n639 163.367
R620 B.n639 B.n638 163.367
R621 B.n638 B.n39 163.367
R622 B.n634 B.n39 163.367
R623 B.n634 B.n633 163.367
R624 B.n633 B.n632 163.367
R625 B.n632 B.n41 163.367
R626 B.n628 B.n41 163.367
R627 B.n628 B.n627 163.367
R628 B.n627 B.n626 163.367
R629 B.n626 B.n43 163.367
R630 B.n622 B.n43 163.367
R631 B.n622 B.n621 163.367
R632 B.n621 B.n620 163.367
R633 B.n620 B.n45 163.367
R634 B.n615 B.n45 163.367
R635 B.n615 B.n614 163.367
R636 B.n614 B.n613 163.367
R637 B.n613 B.n49 163.367
R638 B.n609 B.n49 163.367
R639 B.n609 B.n608 163.367
R640 B.n608 B.n607 163.367
R641 B.n607 B.n51 163.367
R642 B.n603 B.n51 163.367
R643 B.n603 B.n602 163.367
R644 B.n602 B.n55 163.367
R645 B.n598 B.n55 163.367
R646 B.n598 B.n597 163.367
R647 B.n597 B.n596 163.367
R648 B.n596 B.n57 163.367
R649 B.n592 B.n57 163.367
R650 B.n592 B.n591 163.367
R651 B.n591 B.n590 163.367
R652 B.n590 B.n59 163.367
R653 B.n586 B.n59 163.367
R654 B.n586 B.n585 163.367
R655 B.n585 B.n584 163.367
R656 B.n584 B.n61 163.367
R657 B.n580 B.n61 163.367
R658 B.n580 B.n579 163.367
R659 B.n579 B.n578 163.367
R660 B.n578 B.n63 163.367
R661 B.n574 B.n63 163.367
R662 B.n574 B.n573 163.367
R663 B.n573 B.n572 163.367
R664 B.n572 B.n65 163.367
R665 B.n568 B.n65 163.367
R666 B.n568 B.n567 163.367
R667 B.n567 B.n566 163.367
R668 B.n566 B.n67 163.367
R669 B.n562 B.n67 163.367
R670 B.n562 B.n561 163.367
R671 B.n561 B.n560 163.367
R672 B.n560 B.n69 163.367
R673 B.n556 B.n69 163.367
R674 B.n556 B.n555 163.367
R675 B.n555 B.n554 163.367
R676 B.n554 B.n71 163.367
R677 B.n550 B.n71 163.367
R678 B.n550 B.n549 163.367
R679 B.n549 B.n548 163.367
R680 B.n548 B.n73 163.367
R681 B.n544 B.n73 163.367
R682 B.n544 B.n543 163.367
R683 B.n543 B.n542 163.367
R684 B.n542 B.n75 163.367
R685 B.n538 B.n75 163.367
R686 B.n538 B.n537 163.367
R687 B.n537 B.n536 163.367
R688 B.n536 B.n77 163.367
R689 B.n532 B.n77 163.367
R690 B.n532 B.n531 163.367
R691 B.n531 B.n530 163.367
R692 B.n530 B.n79 163.367
R693 B.n526 B.n79 163.367
R694 B.n526 B.n525 163.367
R695 B.n525 B.n524 163.367
R696 B.n524 B.n81 163.367
R697 B.n520 B.n81 163.367
R698 B.n700 B.n17 163.367
R699 B.n704 B.n17 163.367
R700 B.n705 B.n704 163.367
R701 B.n706 B.n705 163.367
R702 B.n706 B.n15 163.367
R703 B.n710 B.n15 163.367
R704 B.n711 B.n710 163.367
R705 B.n712 B.n711 163.367
R706 B.n712 B.n13 163.367
R707 B.n716 B.n13 163.367
R708 B.n717 B.n716 163.367
R709 B.n718 B.n717 163.367
R710 B.n718 B.n11 163.367
R711 B.n722 B.n11 163.367
R712 B.n723 B.n722 163.367
R713 B.n724 B.n723 163.367
R714 B.n724 B.n9 163.367
R715 B.n728 B.n9 163.367
R716 B.n729 B.n728 163.367
R717 B.n730 B.n729 163.367
R718 B.n730 B.n7 163.367
R719 B.n734 B.n7 163.367
R720 B.n735 B.n734 163.367
R721 B.n736 B.n735 163.367
R722 B.n736 B.n5 163.367
R723 B.n740 B.n5 163.367
R724 B.n741 B.n740 163.367
R725 B.n742 B.n741 163.367
R726 B.n742 B.n3 163.367
R727 B.n746 B.n3 163.367
R728 B.n747 B.n746 163.367
R729 B.n192 B.n2 163.367
R730 B.n192 B.n191 163.367
R731 B.n196 B.n191 163.367
R732 B.n197 B.n196 163.367
R733 B.n198 B.n197 163.367
R734 B.n198 B.n189 163.367
R735 B.n202 B.n189 163.367
R736 B.n203 B.n202 163.367
R737 B.n204 B.n203 163.367
R738 B.n204 B.n187 163.367
R739 B.n208 B.n187 163.367
R740 B.n209 B.n208 163.367
R741 B.n210 B.n209 163.367
R742 B.n210 B.n185 163.367
R743 B.n214 B.n185 163.367
R744 B.n215 B.n214 163.367
R745 B.n216 B.n215 163.367
R746 B.n216 B.n183 163.367
R747 B.n220 B.n183 163.367
R748 B.n221 B.n220 163.367
R749 B.n222 B.n221 163.367
R750 B.n222 B.n181 163.367
R751 B.n226 B.n181 163.367
R752 B.n227 B.n226 163.367
R753 B.n228 B.n227 163.367
R754 B.n228 B.n179 163.367
R755 B.n232 B.n179 163.367
R756 B.n233 B.n232 163.367
R757 B.n234 B.n233 163.367
R758 B.n234 B.n177 163.367
R759 B.n238 B.n177 163.367
R760 B.n335 B.t2 109.278
R761 B.n53 B.t4 109.278
R762 B.n149 B.t11 109.257
R763 B.n47 B.t7 109.257
R764 B.n149 B.n148 79.7096
R765 B.n335 B.n334 79.7096
R766 B.n53 B.n52 79.7096
R767 B.n47 B.n46 79.7096
R768 B.n321 B.n149 59.5399
R769 B.n336 B.n335 59.5399
R770 B.n54 B.n53 59.5399
R771 B.n617 B.n47 59.5399
R772 B.n701 B.n18 30.7517
R773 B.n521 B.n82 30.7517
R774 B.n421 B.n420 30.7517
R775 B.n237 B.n176 30.7517
R776 B B.n749 18.0485
R777 B.n702 B.n701 10.6151
R778 B.n703 B.n702 10.6151
R779 B.n703 B.n16 10.6151
R780 B.n707 B.n16 10.6151
R781 B.n708 B.n707 10.6151
R782 B.n709 B.n708 10.6151
R783 B.n709 B.n14 10.6151
R784 B.n713 B.n14 10.6151
R785 B.n714 B.n713 10.6151
R786 B.n715 B.n714 10.6151
R787 B.n715 B.n12 10.6151
R788 B.n719 B.n12 10.6151
R789 B.n720 B.n719 10.6151
R790 B.n721 B.n720 10.6151
R791 B.n721 B.n10 10.6151
R792 B.n725 B.n10 10.6151
R793 B.n726 B.n725 10.6151
R794 B.n727 B.n726 10.6151
R795 B.n727 B.n8 10.6151
R796 B.n731 B.n8 10.6151
R797 B.n732 B.n731 10.6151
R798 B.n733 B.n732 10.6151
R799 B.n733 B.n6 10.6151
R800 B.n737 B.n6 10.6151
R801 B.n738 B.n737 10.6151
R802 B.n739 B.n738 10.6151
R803 B.n739 B.n4 10.6151
R804 B.n743 B.n4 10.6151
R805 B.n744 B.n743 10.6151
R806 B.n745 B.n744 10.6151
R807 B.n745 B.n0 10.6151
R808 B.n697 B.n18 10.6151
R809 B.n697 B.n696 10.6151
R810 B.n696 B.n695 10.6151
R811 B.n695 B.n20 10.6151
R812 B.n691 B.n20 10.6151
R813 B.n691 B.n690 10.6151
R814 B.n690 B.n689 10.6151
R815 B.n689 B.n22 10.6151
R816 B.n685 B.n22 10.6151
R817 B.n685 B.n684 10.6151
R818 B.n684 B.n683 10.6151
R819 B.n683 B.n24 10.6151
R820 B.n679 B.n24 10.6151
R821 B.n679 B.n678 10.6151
R822 B.n678 B.n677 10.6151
R823 B.n677 B.n26 10.6151
R824 B.n673 B.n26 10.6151
R825 B.n673 B.n672 10.6151
R826 B.n672 B.n671 10.6151
R827 B.n671 B.n28 10.6151
R828 B.n667 B.n28 10.6151
R829 B.n667 B.n666 10.6151
R830 B.n666 B.n665 10.6151
R831 B.n665 B.n30 10.6151
R832 B.n661 B.n30 10.6151
R833 B.n661 B.n660 10.6151
R834 B.n660 B.n659 10.6151
R835 B.n659 B.n32 10.6151
R836 B.n655 B.n32 10.6151
R837 B.n655 B.n654 10.6151
R838 B.n654 B.n653 10.6151
R839 B.n653 B.n34 10.6151
R840 B.n649 B.n34 10.6151
R841 B.n649 B.n648 10.6151
R842 B.n648 B.n647 10.6151
R843 B.n647 B.n36 10.6151
R844 B.n643 B.n36 10.6151
R845 B.n643 B.n642 10.6151
R846 B.n642 B.n641 10.6151
R847 B.n641 B.n38 10.6151
R848 B.n637 B.n38 10.6151
R849 B.n637 B.n636 10.6151
R850 B.n636 B.n635 10.6151
R851 B.n635 B.n40 10.6151
R852 B.n631 B.n40 10.6151
R853 B.n631 B.n630 10.6151
R854 B.n630 B.n629 10.6151
R855 B.n629 B.n42 10.6151
R856 B.n625 B.n42 10.6151
R857 B.n625 B.n624 10.6151
R858 B.n624 B.n623 10.6151
R859 B.n623 B.n44 10.6151
R860 B.n619 B.n44 10.6151
R861 B.n619 B.n618 10.6151
R862 B.n616 B.n48 10.6151
R863 B.n612 B.n48 10.6151
R864 B.n612 B.n611 10.6151
R865 B.n611 B.n610 10.6151
R866 B.n610 B.n50 10.6151
R867 B.n606 B.n50 10.6151
R868 B.n606 B.n605 10.6151
R869 B.n605 B.n604 10.6151
R870 B.n601 B.n600 10.6151
R871 B.n600 B.n599 10.6151
R872 B.n599 B.n56 10.6151
R873 B.n595 B.n56 10.6151
R874 B.n595 B.n594 10.6151
R875 B.n594 B.n593 10.6151
R876 B.n593 B.n58 10.6151
R877 B.n589 B.n58 10.6151
R878 B.n589 B.n588 10.6151
R879 B.n588 B.n587 10.6151
R880 B.n587 B.n60 10.6151
R881 B.n583 B.n60 10.6151
R882 B.n583 B.n582 10.6151
R883 B.n582 B.n581 10.6151
R884 B.n581 B.n62 10.6151
R885 B.n577 B.n62 10.6151
R886 B.n577 B.n576 10.6151
R887 B.n576 B.n575 10.6151
R888 B.n575 B.n64 10.6151
R889 B.n571 B.n64 10.6151
R890 B.n571 B.n570 10.6151
R891 B.n570 B.n569 10.6151
R892 B.n569 B.n66 10.6151
R893 B.n565 B.n66 10.6151
R894 B.n565 B.n564 10.6151
R895 B.n564 B.n563 10.6151
R896 B.n563 B.n68 10.6151
R897 B.n559 B.n68 10.6151
R898 B.n559 B.n558 10.6151
R899 B.n558 B.n557 10.6151
R900 B.n557 B.n70 10.6151
R901 B.n553 B.n70 10.6151
R902 B.n553 B.n552 10.6151
R903 B.n552 B.n551 10.6151
R904 B.n551 B.n72 10.6151
R905 B.n547 B.n72 10.6151
R906 B.n547 B.n546 10.6151
R907 B.n546 B.n545 10.6151
R908 B.n545 B.n74 10.6151
R909 B.n541 B.n74 10.6151
R910 B.n541 B.n540 10.6151
R911 B.n540 B.n539 10.6151
R912 B.n539 B.n76 10.6151
R913 B.n535 B.n76 10.6151
R914 B.n535 B.n534 10.6151
R915 B.n534 B.n533 10.6151
R916 B.n533 B.n78 10.6151
R917 B.n529 B.n78 10.6151
R918 B.n529 B.n528 10.6151
R919 B.n528 B.n527 10.6151
R920 B.n527 B.n80 10.6151
R921 B.n523 B.n80 10.6151
R922 B.n523 B.n522 10.6151
R923 B.n522 B.n521 10.6151
R924 B.n517 B.n82 10.6151
R925 B.n517 B.n516 10.6151
R926 B.n516 B.n515 10.6151
R927 B.n515 B.n84 10.6151
R928 B.n511 B.n84 10.6151
R929 B.n511 B.n510 10.6151
R930 B.n510 B.n509 10.6151
R931 B.n509 B.n86 10.6151
R932 B.n505 B.n86 10.6151
R933 B.n505 B.n504 10.6151
R934 B.n504 B.n503 10.6151
R935 B.n503 B.n88 10.6151
R936 B.n499 B.n88 10.6151
R937 B.n499 B.n498 10.6151
R938 B.n498 B.n497 10.6151
R939 B.n497 B.n90 10.6151
R940 B.n493 B.n90 10.6151
R941 B.n493 B.n492 10.6151
R942 B.n492 B.n491 10.6151
R943 B.n491 B.n92 10.6151
R944 B.n487 B.n92 10.6151
R945 B.n487 B.n486 10.6151
R946 B.n486 B.n485 10.6151
R947 B.n485 B.n94 10.6151
R948 B.n481 B.n94 10.6151
R949 B.n481 B.n480 10.6151
R950 B.n480 B.n479 10.6151
R951 B.n479 B.n96 10.6151
R952 B.n475 B.n96 10.6151
R953 B.n475 B.n474 10.6151
R954 B.n474 B.n473 10.6151
R955 B.n473 B.n98 10.6151
R956 B.n469 B.n98 10.6151
R957 B.n469 B.n468 10.6151
R958 B.n468 B.n467 10.6151
R959 B.n467 B.n100 10.6151
R960 B.n463 B.n100 10.6151
R961 B.n463 B.n462 10.6151
R962 B.n462 B.n461 10.6151
R963 B.n461 B.n102 10.6151
R964 B.n457 B.n102 10.6151
R965 B.n457 B.n456 10.6151
R966 B.n456 B.n455 10.6151
R967 B.n455 B.n104 10.6151
R968 B.n451 B.n104 10.6151
R969 B.n451 B.n450 10.6151
R970 B.n450 B.n449 10.6151
R971 B.n449 B.n106 10.6151
R972 B.n445 B.n106 10.6151
R973 B.n445 B.n444 10.6151
R974 B.n444 B.n443 10.6151
R975 B.n443 B.n108 10.6151
R976 B.n439 B.n108 10.6151
R977 B.n439 B.n438 10.6151
R978 B.n438 B.n437 10.6151
R979 B.n437 B.n110 10.6151
R980 B.n433 B.n110 10.6151
R981 B.n433 B.n432 10.6151
R982 B.n432 B.n431 10.6151
R983 B.n431 B.n112 10.6151
R984 B.n427 B.n112 10.6151
R985 B.n427 B.n426 10.6151
R986 B.n426 B.n425 10.6151
R987 B.n425 B.n114 10.6151
R988 B.n421 B.n114 10.6151
R989 B.n193 B.n1 10.6151
R990 B.n194 B.n193 10.6151
R991 B.n195 B.n194 10.6151
R992 B.n195 B.n190 10.6151
R993 B.n199 B.n190 10.6151
R994 B.n200 B.n199 10.6151
R995 B.n201 B.n200 10.6151
R996 B.n201 B.n188 10.6151
R997 B.n205 B.n188 10.6151
R998 B.n206 B.n205 10.6151
R999 B.n207 B.n206 10.6151
R1000 B.n207 B.n186 10.6151
R1001 B.n211 B.n186 10.6151
R1002 B.n212 B.n211 10.6151
R1003 B.n213 B.n212 10.6151
R1004 B.n213 B.n184 10.6151
R1005 B.n217 B.n184 10.6151
R1006 B.n218 B.n217 10.6151
R1007 B.n219 B.n218 10.6151
R1008 B.n219 B.n182 10.6151
R1009 B.n223 B.n182 10.6151
R1010 B.n224 B.n223 10.6151
R1011 B.n225 B.n224 10.6151
R1012 B.n225 B.n180 10.6151
R1013 B.n229 B.n180 10.6151
R1014 B.n230 B.n229 10.6151
R1015 B.n231 B.n230 10.6151
R1016 B.n231 B.n178 10.6151
R1017 B.n235 B.n178 10.6151
R1018 B.n236 B.n235 10.6151
R1019 B.n237 B.n236 10.6151
R1020 B.n241 B.n176 10.6151
R1021 B.n242 B.n241 10.6151
R1022 B.n243 B.n242 10.6151
R1023 B.n243 B.n174 10.6151
R1024 B.n247 B.n174 10.6151
R1025 B.n248 B.n247 10.6151
R1026 B.n249 B.n248 10.6151
R1027 B.n249 B.n172 10.6151
R1028 B.n253 B.n172 10.6151
R1029 B.n254 B.n253 10.6151
R1030 B.n255 B.n254 10.6151
R1031 B.n255 B.n170 10.6151
R1032 B.n259 B.n170 10.6151
R1033 B.n260 B.n259 10.6151
R1034 B.n261 B.n260 10.6151
R1035 B.n261 B.n168 10.6151
R1036 B.n265 B.n168 10.6151
R1037 B.n266 B.n265 10.6151
R1038 B.n267 B.n266 10.6151
R1039 B.n267 B.n166 10.6151
R1040 B.n271 B.n166 10.6151
R1041 B.n272 B.n271 10.6151
R1042 B.n273 B.n272 10.6151
R1043 B.n273 B.n164 10.6151
R1044 B.n277 B.n164 10.6151
R1045 B.n278 B.n277 10.6151
R1046 B.n279 B.n278 10.6151
R1047 B.n279 B.n162 10.6151
R1048 B.n283 B.n162 10.6151
R1049 B.n284 B.n283 10.6151
R1050 B.n285 B.n284 10.6151
R1051 B.n285 B.n160 10.6151
R1052 B.n289 B.n160 10.6151
R1053 B.n290 B.n289 10.6151
R1054 B.n291 B.n290 10.6151
R1055 B.n291 B.n158 10.6151
R1056 B.n295 B.n158 10.6151
R1057 B.n296 B.n295 10.6151
R1058 B.n297 B.n296 10.6151
R1059 B.n297 B.n156 10.6151
R1060 B.n301 B.n156 10.6151
R1061 B.n302 B.n301 10.6151
R1062 B.n303 B.n302 10.6151
R1063 B.n303 B.n154 10.6151
R1064 B.n307 B.n154 10.6151
R1065 B.n308 B.n307 10.6151
R1066 B.n309 B.n308 10.6151
R1067 B.n309 B.n152 10.6151
R1068 B.n313 B.n152 10.6151
R1069 B.n314 B.n313 10.6151
R1070 B.n315 B.n314 10.6151
R1071 B.n315 B.n150 10.6151
R1072 B.n319 B.n150 10.6151
R1073 B.n320 B.n319 10.6151
R1074 B.n322 B.n146 10.6151
R1075 B.n326 B.n146 10.6151
R1076 B.n327 B.n326 10.6151
R1077 B.n328 B.n327 10.6151
R1078 B.n328 B.n144 10.6151
R1079 B.n332 B.n144 10.6151
R1080 B.n333 B.n332 10.6151
R1081 B.n337 B.n333 10.6151
R1082 B.n341 B.n142 10.6151
R1083 B.n342 B.n341 10.6151
R1084 B.n343 B.n342 10.6151
R1085 B.n343 B.n140 10.6151
R1086 B.n347 B.n140 10.6151
R1087 B.n348 B.n347 10.6151
R1088 B.n349 B.n348 10.6151
R1089 B.n349 B.n138 10.6151
R1090 B.n353 B.n138 10.6151
R1091 B.n354 B.n353 10.6151
R1092 B.n355 B.n354 10.6151
R1093 B.n355 B.n136 10.6151
R1094 B.n359 B.n136 10.6151
R1095 B.n360 B.n359 10.6151
R1096 B.n361 B.n360 10.6151
R1097 B.n361 B.n134 10.6151
R1098 B.n365 B.n134 10.6151
R1099 B.n366 B.n365 10.6151
R1100 B.n367 B.n366 10.6151
R1101 B.n367 B.n132 10.6151
R1102 B.n371 B.n132 10.6151
R1103 B.n372 B.n371 10.6151
R1104 B.n373 B.n372 10.6151
R1105 B.n373 B.n130 10.6151
R1106 B.n377 B.n130 10.6151
R1107 B.n378 B.n377 10.6151
R1108 B.n379 B.n378 10.6151
R1109 B.n379 B.n128 10.6151
R1110 B.n383 B.n128 10.6151
R1111 B.n384 B.n383 10.6151
R1112 B.n385 B.n384 10.6151
R1113 B.n385 B.n126 10.6151
R1114 B.n389 B.n126 10.6151
R1115 B.n390 B.n389 10.6151
R1116 B.n391 B.n390 10.6151
R1117 B.n391 B.n124 10.6151
R1118 B.n395 B.n124 10.6151
R1119 B.n396 B.n395 10.6151
R1120 B.n397 B.n396 10.6151
R1121 B.n397 B.n122 10.6151
R1122 B.n401 B.n122 10.6151
R1123 B.n402 B.n401 10.6151
R1124 B.n403 B.n402 10.6151
R1125 B.n403 B.n120 10.6151
R1126 B.n407 B.n120 10.6151
R1127 B.n408 B.n407 10.6151
R1128 B.n409 B.n408 10.6151
R1129 B.n409 B.n118 10.6151
R1130 B.n413 B.n118 10.6151
R1131 B.n414 B.n413 10.6151
R1132 B.n415 B.n414 10.6151
R1133 B.n415 B.n116 10.6151
R1134 B.n419 B.n116 10.6151
R1135 B.n420 B.n419 10.6151
R1136 B.n749 B.n0 8.11757
R1137 B.n749 B.n1 8.11757
R1138 B.n617 B.n616 6.5566
R1139 B.n604 B.n54 6.5566
R1140 B.n322 B.n321 6.5566
R1141 B.n337 B.n336 6.5566
R1142 B.n618 B.n617 4.05904
R1143 B.n601 B.n54 4.05904
R1144 B.n321 B.n320 4.05904
R1145 B.n336 B.n142 4.05904
R1146 VN VN.t0 191.03
R1147 VN VN.t1 140.666
R1148 VDD2.n0 VDD2.t0 117.091
R1149 VDD2.n0 VDD2.t1 72.1466
R1150 VDD2 VDD2.n0 0.944465
C0 B VP 1.85702f
C1 VN VTAIL 3.43612f
C2 VN VDD2 3.91142f
C3 VDD2 VTAIL 6.48115f
C4 B w_n2614_n4262# 11.336901f
C5 VN VDD1 0.148664f
C6 VTAIL VDD1 6.42237f
C7 VDD2 VDD1 0.805775f
C8 VN VP 6.83977f
C9 VP VTAIL 3.451f
C10 VP VDD2 0.382292f
C11 VN w_n2614_n4262# 3.81134f
C12 VTAIL w_n2614_n4262# 3.37657f
C13 VDD2 w_n2614_n4262# 2.25654f
C14 VP VDD1 4.14302f
C15 VDD1 w_n2614_n4262# 2.21613f
C16 B VN 1.30068f
C17 B VTAIL 5.15207f
C18 B VDD2 2.26238f
C19 VP w_n2614_n4262# 4.14685f
C20 B VDD1 2.22172f
C21 VDD2 VSUBS 1.218371f
C22 VDD1 VSUBS 7.04745f
C23 VTAIL VSUBS 1.29806f
C24 VN VSUBS 9.05042f
C25 VP VSUBS 2.193225f
C26 B VSUBS 5.152896f
C27 w_n2614_n4262# VSUBS 0.136419p
C28 VDD2.t0 VSUBS 5.14334f
C29 VDD2.t1 VSUBS 4.04013f
C30 VDD2.n0 VSUBS 5.56131f
C31 VN.t1 VSUBS 5.52005f
C32 VN.t0 VSUBS 6.42158f
C33 B.n0 VSUBS 0.005629f
C34 B.n1 VSUBS 0.005629f
C35 B.n2 VSUBS 0.008325f
C36 B.n3 VSUBS 0.00638f
C37 B.n4 VSUBS 0.00638f
C38 B.n5 VSUBS 0.00638f
C39 B.n6 VSUBS 0.00638f
C40 B.n7 VSUBS 0.00638f
C41 B.n8 VSUBS 0.00638f
C42 B.n9 VSUBS 0.00638f
C43 B.n10 VSUBS 0.00638f
C44 B.n11 VSUBS 0.00638f
C45 B.n12 VSUBS 0.00638f
C46 B.n13 VSUBS 0.00638f
C47 B.n14 VSUBS 0.00638f
C48 B.n15 VSUBS 0.00638f
C49 B.n16 VSUBS 0.00638f
C50 B.n17 VSUBS 0.00638f
C51 B.n18 VSUBS 0.01456f
C52 B.n19 VSUBS 0.00638f
C53 B.n20 VSUBS 0.00638f
C54 B.n21 VSUBS 0.00638f
C55 B.n22 VSUBS 0.00638f
C56 B.n23 VSUBS 0.00638f
C57 B.n24 VSUBS 0.00638f
C58 B.n25 VSUBS 0.00638f
C59 B.n26 VSUBS 0.00638f
C60 B.n27 VSUBS 0.00638f
C61 B.n28 VSUBS 0.00638f
C62 B.n29 VSUBS 0.00638f
C63 B.n30 VSUBS 0.00638f
C64 B.n31 VSUBS 0.00638f
C65 B.n32 VSUBS 0.00638f
C66 B.n33 VSUBS 0.00638f
C67 B.n34 VSUBS 0.00638f
C68 B.n35 VSUBS 0.00638f
C69 B.n36 VSUBS 0.00638f
C70 B.n37 VSUBS 0.00638f
C71 B.n38 VSUBS 0.00638f
C72 B.n39 VSUBS 0.00638f
C73 B.n40 VSUBS 0.00638f
C74 B.n41 VSUBS 0.00638f
C75 B.n42 VSUBS 0.00638f
C76 B.n43 VSUBS 0.00638f
C77 B.n44 VSUBS 0.00638f
C78 B.n45 VSUBS 0.00638f
C79 B.t7 VSUBS 0.503482f
C80 B.t8 VSUBS 0.529221f
C81 B.t6 VSUBS 2.5987f
C82 B.n46 VSUBS 0.32186f
C83 B.n47 VSUBS 0.070119f
C84 B.n48 VSUBS 0.00638f
C85 B.n49 VSUBS 0.00638f
C86 B.n50 VSUBS 0.00638f
C87 B.n51 VSUBS 0.00638f
C88 B.t4 VSUBS 0.503465f
C89 B.t5 VSUBS 0.529209f
C90 B.t3 VSUBS 2.5987f
C91 B.n52 VSUBS 0.321872f
C92 B.n53 VSUBS 0.070136f
C93 B.n54 VSUBS 0.014781f
C94 B.n55 VSUBS 0.00638f
C95 B.n56 VSUBS 0.00638f
C96 B.n57 VSUBS 0.00638f
C97 B.n58 VSUBS 0.00638f
C98 B.n59 VSUBS 0.00638f
C99 B.n60 VSUBS 0.00638f
C100 B.n61 VSUBS 0.00638f
C101 B.n62 VSUBS 0.00638f
C102 B.n63 VSUBS 0.00638f
C103 B.n64 VSUBS 0.00638f
C104 B.n65 VSUBS 0.00638f
C105 B.n66 VSUBS 0.00638f
C106 B.n67 VSUBS 0.00638f
C107 B.n68 VSUBS 0.00638f
C108 B.n69 VSUBS 0.00638f
C109 B.n70 VSUBS 0.00638f
C110 B.n71 VSUBS 0.00638f
C111 B.n72 VSUBS 0.00638f
C112 B.n73 VSUBS 0.00638f
C113 B.n74 VSUBS 0.00638f
C114 B.n75 VSUBS 0.00638f
C115 B.n76 VSUBS 0.00638f
C116 B.n77 VSUBS 0.00638f
C117 B.n78 VSUBS 0.00638f
C118 B.n79 VSUBS 0.00638f
C119 B.n80 VSUBS 0.00638f
C120 B.n81 VSUBS 0.00638f
C121 B.n82 VSUBS 0.01415f
C122 B.n83 VSUBS 0.00638f
C123 B.n84 VSUBS 0.00638f
C124 B.n85 VSUBS 0.00638f
C125 B.n86 VSUBS 0.00638f
C126 B.n87 VSUBS 0.00638f
C127 B.n88 VSUBS 0.00638f
C128 B.n89 VSUBS 0.00638f
C129 B.n90 VSUBS 0.00638f
C130 B.n91 VSUBS 0.00638f
C131 B.n92 VSUBS 0.00638f
C132 B.n93 VSUBS 0.00638f
C133 B.n94 VSUBS 0.00638f
C134 B.n95 VSUBS 0.00638f
C135 B.n96 VSUBS 0.00638f
C136 B.n97 VSUBS 0.00638f
C137 B.n98 VSUBS 0.00638f
C138 B.n99 VSUBS 0.00638f
C139 B.n100 VSUBS 0.00638f
C140 B.n101 VSUBS 0.00638f
C141 B.n102 VSUBS 0.00638f
C142 B.n103 VSUBS 0.00638f
C143 B.n104 VSUBS 0.00638f
C144 B.n105 VSUBS 0.00638f
C145 B.n106 VSUBS 0.00638f
C146 B.n107 VSUBS 0.00638f
C147 B.n108 VSUBS 0.00638f
C148 B.n109 VSUBS 0.00638f
C149 B.n110 VSUBS 0.00638f
C150 B.n111 VSUBS 0.00638f
C151 B.n112 VSUBS 0.00638f
C152 B.n113 VSUBS 0.00638f
C153 B.n114 VSUBS 0.00638f
C154 B.n115 VSUBS 0.01456f
C155 B.n116 VSUBS 0.00638f
C156 B.n117 VSUBS 0.00638f
C157 B.n118 VSUBS 0.00638f
C158 B.n119 VSUBS 0.00638f
C159 B.n120 VSUBS 0.00638f
C160 B.n121 VSUBS 0.00638f
C161 B.n122 VSUBS 0.00638f
C162 B.n123 VSUBS 0.00638f
C163 B.n124 VSUBS 0.00638f
C164 B.n125 VSUBS 0.00638f
C165 B.n126 VSUBS 0.00638f
C166 B.n127 VSUBS 0.00638f
C167 B.n128 VSUBS 0.00638f
C168 B.n129 VSUBS 0.00638f
C169 B.n130 VSUBS 0.00638f
C170 B.n131 VSUBS 0.00638f
C171 B.n132 VSUBS 0.00638f
C172 B.n133 VSUBS 0.00638f
C173 B.n134 VSUBS 0.00638f
C174 B.n135 VSUBS 0.00638f
C175 B.n136 VSUBS 0.00638f
C176 B.n137 VSUBS 0.00638f
C177 B.n138 VSUBS 0.00638f
C178 B.n139 VSUBS 0.00638f
C179 B.n140 VSUBS 0.00638f
C180 B.n141 VSUBS 0.00638f
C181 B.n142 VSUBS 0.00441f
C182 B.n143 VSUBS 0.00638f
C183 B.n144 VSUBS 0.00638f
C184 B.n145 VSUBS 0.00638f
C185 B.n146 VSUBS 0.00638f
C186 B.n147 VSUBS 0.00638f
C187 B.t11 VSUBS 0.503482f
C188 B.t10 VSUBS 0.529221f
C189 B.t9 VSUBS 2.5987f
C190 B.n148 VSUBS 0.32186f
C191 B.n149 VSUBS 0.070119f
C192 B.n150 VSUBS 0.00638f
C193 B.n151 VSUBS 0.00638f
C194 B.n152 VSUBS 0.00638f
C195 B.n153 VSUBS 0.00638f
C196 B.n154 VSUBS 0.00638f
C197 B.n155 VSUBS 0.00638f
C198 B.n156 VSUBS 0.00638f
C199 B.n157 VSUBS 0.00638f
C200 B.n158 VSUBS 0.00638f
C201 B.n159 VSUBS 0.00638f
C202 B.n160 VSUBS 0.00638f
C203 B.n161 VSUBS 0.00638f
C204 B.n162 VSUBS 0.00638f
C205 B.n163 VSUBS 0.00638f
C206 B.n164 VSUBS 0.00638f
C207 B.n165 VSUBS 0.00638f
C208 B.n166 VSUBS 0.00638f
C209 B.n167 VSUBS 0.00638f
C210 B.n168 VSUBS 0.00638f
C211 B.n169 VSUBS 0.00638f
C212 B.n170 VSUBS 0.00638f
C213 B.n171 VSUBS 0.00638f
C214 B.n172 VSUBS 0.00638f
C215 B.n173 VSUBS 0.00638f
C216 B.n174 VSUBS 0.00638f
C217 B.n175 VSUBS 0.00638f
C218 B.n176 VSUBS 0.01456f
C219 B.n177 VSUBS 0.00638f
C220 B.n178 VSUBS 0.00638f
C221 B.n179 VSUBS 0.00638f
C222 B.n180 VSUBS 0.00638f
C223 B.n181 VSUBS 0.00638f
C224 B.n182 VSUBS 0.00638f
C225 B.n183 VSUBS 0.00638f
C226 B.n184 VSUBS 0.00638f
C227 B.n185 VSUBS 0.00638f
C228 B.n186 VSUBS 0.00638f
C229 B.n187 VSUBS 0.00638f
C230 B.n188 VSUBS 0.00638f
C231 B.n189 VSUBS 0.00638f
C232 B.n190 VSUBS 0.00638f
C233 B.n191 VSUBS 0.00638f
C234 B.n192 VSUBS 0.00638f
C235 B.n193 VSUBS 0.00638f
C236 B.n194 VSUBS 0.00638f
C237 B.n195 VSUBS 0.00638f
C238 B.n196 VSUBS 0.00638f
C239 B.n197 VSUBS 0.00638f
C240 B.n198 VSUBS 0.00638f
C241 B.n199 VSUBS 0.00638f
C242 B.n200 VSUBS 0.00638f
C243 B.n201 VSUBS 0.00638f
C244 B.n202 VSUBS 0.00638f
C245 B.n203 VSUBS 0.00638f
C246 B.n204 VSUBS 0.00638f
C247 B.n205 VSUBS 0.00638f
C248 B.n206 VSUBS 0.00638f
C249 B.n207 VSUBS 0.00638f
C250 B.n208 VSUBS 0.00638f
C251 B.n209 VSUBS 0.00638f
C252 B.n210 VSUBS 0.00638f
C253 B.n211 VSUBS 0.00638f
C254 B.n212 VSUBS 0.00638f
C255 B.n213 VSUBS 0.00638f
C256 B.n214 VSUBS 0.00638f
C257 B.n215 VSUBS 0.00638f
C258 B.n216 VSUBS 0.00638f
C259 B.n217 VSUBS 0.00638f
C260 B.n218 VSUBS 0.00638f
C261 B.n219 VSUBS 0.00638f
C262 B.n220 VSUBS 0.00638f
C263 B.n221 VSUBS 0.00638f
C264 B.n222 VSUBS 0.00638f
C265 B.n223 VSUBS 0.00638f
C266 B.n224 VSUBS 0.00638f
C267 B.n225 VSUBS 0.00638f
C268 B.n226 VSUBS 0.00638f
C269 B.n227 VSUBS 0.00638f
C270 B.n228 VSUBS 0.00638f
C271 B.n229 VSUBS 0.00638f
C272 B.n230 VSUBS 0.00638f
C273 B.n231 VSUBS 0.00638f
C274 B.n232 VSUBS 0.00638f
C275 B.n233 VSUBS 0.00638f
C276 B.n234 VSUBS 0.00638f
C277 B.n235 VSUBS 0.00638f
C278 B.n236 VSUBS 0.00638f
C279 B.n237 VSUBS 0.01415f
C280 B.n238 VSUBS 0.01415f
C281 B.n239 VSUBS 0.01456f
C282 B.n240 VSUBS 0.00638f
C283 B.n241 VSUBS 0.00638f
C284 B.n242 VSUBS 0.00638f
C285 B.n243 VSUBS 0.00638f
C286 B.n244 VSUBS 0.00638f
C287 B.n245 VSUBS 0.00638f
C288 B.n246 VSUBS 0.00638f
C289 B.n247 VSUBS 0.00638f
C290 B.n248 VSUBS 0.00638f
C291 B.n249 VSUBS 0.00638f
C292 B.n250 VSUBS 0.00638f
C293 B.n251 VSUBS 0.00638f
C294 B.n252 VSUBS 0.00638f
C295 B.n253 VSUBS 0.00638f
C296 B.n254 VSUBS 0.00638f
C297 B.n255 VSUBS 0.00638f
C298 B.n256 VSUBS 0.00638f
C299 B.n257 VSUBS 0.00638f
C300 B.n258 VSUBS 0.00638f
C301 B.n259 VSUBS 0.00638f
C302 B.n260 VSUBS 0.00638f
C303 B.n261 VSUBS 0.00638f
C304 B.n262 VSUBS 0.00638f
C305 B.n263 VSUBS 0.00638f
C306 B.n264 VSUBS 0.00638f
C307 B.n265 VSUBS 0.00638f
C308 B.n266 VSUBS 0.00638f
C309 B.n267 VSUBS 0.00638f
C310 B.n268 VSUBS 0.00638f
C311 B.n269 VSUBS 0.00638f
C312 B.n270 VSUBS 0.00638f
C313 B.n271 VSUBS 0.00638f
C314 B.n272 VSUBS 0.00638f
C315 B.n273 VSUBS 0.00638f
C316 B.n274 VSUBS 0.00638f
C317 B.n275 VSUBS 0.00638f
C318 B.n276 VSUBS 0.00638f
C319 B.n277 VSUBS 0.00638f
C320 B.n278 VSUBS 0.00638f
C321 B.n279 VSUBS 0.00638f
C322 B.n280 VSUBS 0.00638f
C323 B.n281 VSUBS 0.00638f
C324 B.n282 VSUBS 0.00638f
C325 B.n283 VSUBS 0.00638f
C326 B.n284 VSUBS 0.00638f
C327 B.n285 VSUBS 0.00638f
C328 B.n286 VSUBS 0.00638f
C329 B.n287 VSUBS 0.00638f
C330 B.n288 VSUBS 0.00638f
C331 B.n289 VSUBS 0.00638f
C332 B.n290 VSUBS 0.00638f
C333 B.n291 VSUBS 0.00638f
C334 B.n292 VSUBS 0.00638f
C335 B.n293 VSUBS 0.00638f
C336 B.n294 VSUBS 0.00638f
C337 B.n295 VSUBS 0.00638f
C338 B.n296 VSUBS 0.00638f
C339 B.n297 VSUBS 0.00638f
C340 B.n298 VSUBS 0.00638f
C341 B.n299 VSUBS 0.00638f
C342 B.n300 VSUBS 0.00638f
C343 B.n301 VSUBS 0.00638f
C344 B.n302 VSUBS 0.00638f
C345 B.n303 VSUBS 0.00638f
C346 B.n304 VSUBS 0.00638f
C347 B.n305 VSUBS 0.00638f
C348 B.n306 VSUBS 0.00638f
C349 B.n307 VSUBS 0.00638f
C350 B.n308 VSUBS 0.00638f
C351 B.n309 VSUBS 0.00638f
C352 B.n310 VSUBS 0.00638f
C353 B.n311 VSUBS 0.00638f
C354 B.n312 VSUBS 0.00638f
C355 B.n313 VSUBS 0.00638f
C356 B.n314 VSUBS 0.00638f
C357 B.n315 VSUBS 0.00638f
C358 B.n316 VSUBS 0.00638f
C359 B.n317 VSUBS 0.00638f
C360 B.n318 VSUBS 0.00638f
C361 B.n319 VSUBS 0.00638f
C362 B.n320 VSUBS 0.00441f
C363 B.n321 VSUBS 0.014781f
C364 B.n322 VSUBS 0.00516f
C365 B.n323 VSUBS 0.00638f
C366 B.n324 VSUBS 0.00638f
C367 B.n325 VSUBS 0.00638f
C368 B.n326 VSUBS 0.00638f
C369 B.n327 VSUBS 0.00638f
C370 B.n328 VSUBS 0.00638f
C371 B.n329 VSUBS 0.00638f
C372 B.n330 VSUBS 0.00638f
C373 B.n331 VSUBS 0.00638f
C374 B.n332 VSUBS 0.00638f
C375 B.n333 VSUBS 0.00638f
C376 B.t2 VSUBS 0.503465f
C377 B.t1 VSUBS 0.529209f
C378 B.t0 VSUBS 2.5987f
C379 B.n334 VSUBS 0.321872f
C380 B.n335 VSUBS 0.070136f
C381 B.n336 VSUBS 0.014781f
C382 B.n337 VSUBS 0.00516f
C383 B.n338 VSUBS 0.00638f
C384 B.n339 VSUBS 0.00638f
C385 B.n340 VSUBS 0.00638f
C386 B.n341 VSUBS 0.00638f
C387 B.n342 VSUBS 0.00638f
C388 B.n343 VSUBS 0.00638f
C389 B.n344 VSUBS 0.00638f
C390 B.n345 VSUBS 0.00638f
C391 B.n346 VSUBS 0.00638f
C392 B.n347 VSUBS 0.00638f
C393 B.n348 VSUBS 0.00638f
C394 B.n349 VSUBS 0.00638f
C395 B.n350 VSUBS 0.00638f
C396 B.n351 VSUBS 0.00638f
C397 B.n352 VSUBS 0.00638f
C398 B.n353 VSUBS 0.00638f
C399 B.n354 VSUBS 0.00638f
C400 B.n355 VSUBS 0.00638f
C401 B.n356 VSUBS 0.00638f
C402 B.n357 VSUBS 0.00638f
C403 B.n358 VSUBS 0.00638f
C404 B.n359 VSUBS 0.00638f
C405 B.n360 VSUBS 0.00638f
C406 B.n361 VSUBS 0.00638f
C407 B.n362 VSUBS 0.00638f
C408 B.n363 VSUBS 0.00638f
C409 B.n364 VSUBS 0.00638f
C410 B.n365 VSUBS 0.00638f
C411 B.n366 VSUBS 0.00638f
C412 B.n367 VSUBS 0.00638f
C413 B.n368 VSUBS 0.00638f
C414 B.n369 VSUBS 0.00638f
C415 B.n370 VSUBS 0.00638f
C416 B.n371 VSUBS 0.00638f
C417 B.n372 VSUBS 0.00638f
C418 B.n373 VSUBS 0.00638f
C419 B.n374 VSUBS 0.00638f
C420 B.n375 VSUBS 0.00638f
C421 B.n376 VSUBS 0.00638f
C422 B.n377 VSUBS 0.00638f
C423 B.n378 VSUBS 0.00638f
C424 B.n379 VSUBS 0.00638f
C425 B.n380 VSUBS 0.00638f
C426 B.n381 VSUBS 0.00638f
C427 B.n382 VSUBS 0.00638f
C428 B.n383 VSUBS 0.00638f
C429 B.n384 VSUBS 0.00638f
C430 B.n385 VSUBS 0.00638f
C431 B.n386 VSUBS 0.00638f
C432 B.n387 VSUBS 0.00638f
C433 B.n388 VSUBS 0.00638f
C434 B.n389 VSUBS 0.00638f
C435 B.n390 VSUBS 0.00638f
C436 B.n391 VSUBS 0.00638f
C437 B.n392 VSUBS 0.00638f
C438 B.n393 VSUBS 0.00638f
C439 B.n394 VSUBS 0.00638f
C440 B.n395 VSUBS 0.00638f
C441 B.n396 VSUBS 0.00638f
C442 B.n397 VSUBS 0.00638f
C443 B.n398 VSUBS 0.00638f
C444 B.n399 VSUBS 0.00638f
C445 B.n400 VSUBS 0.00638f
C446 B.n401 VSUBS 0.00638f
C447 B.n402 VSUBS 0.00638f
C448 B.n403 VSUBS 0.00638f
C449 B.n404 VSUBS 0.00638f
C450 B.n405 VSUBS 0.00638f
C451 B.n406 VSUBS 0.00638f
C452 B.n407 VSUBS 0.00638f
C453 B.n408 VSUBS 0.00638f
C454 B.n409 VSUBS 0.00638f
C455 B.n410 VSUBS 0.00638f
C456 B.n411 VSUBS 0.00638f
C457 B.n412 VSUBS 0.00638f
C458 B.n413 VSUBS 0.00638f
C459 B.n414 VSUBS 0.00638f
C460 B.n415 VSUBS 0.00638f
C461 B.n416 VSUBS 0.00638f
C462 B.n417 VSUBS 0.00638f
C463 B.n418 VSUBS 0.00638f
C464 B.n419 VSUBS 0.00638f
C465 B.n420 VSUBS 0.013759f
C466 B.n421 VSUBS 0.01495f
C467 B.n422 VSUBS 0.01415f
C468 B.n423 VSUBS 0.00638f
C469 B.n424 VSUBS 0.00638f
C470 B.n425 VSUBS 0.00638f
C471 B.n426 VSUBS 0.00638f
C472 B.n427 VSUBS 0.00638f
C473 B.n428 VSUBS 0.00638f
C474 B.n429 VSUBS 0.00638f
C475 B.n430 VSUBS 0.00638f
C476 B.n431 VSUBS 0.00638f
C477 B.n432 VSUBS 0.00638f
C478 B.n433 VSUBS 0.00638f
C479 B.n434 VSUBS 0.00638f
C480 B.n435 VSUBS 0.00638f
C481 B.n436 VSUBS 0.00638f
C482 B.n437 VSUBS 0.00638f
C483 B.n438 VSUBS 0.00638f
C484 B.n439 VSUBS 0.00638f
C485 B.n440 VSUBS 0.00638f
C486 B.n441 VSUBS 0.00638f
C487 B.n442 VSUBS 0.00638f
C488 B.n443 VSUBS 0.00638f
C489 B.n444 VSUBS 0.00638f
C490 B.n445 VSUBS 0.00638f
C491 B.n446 VSUBS 0.00638f
C492 B.n447 VSUBS 0.00638f
C493 B.n448 VSUBS 0.00638f
C494 B.n449 VSUBS 0.00638f
C495 B.n450 VSUBS 0.00638f
C496 B.n451 VSUBS 0.00638f
C497 B.n452 VSUBS 0.00638f
C498 B.n453 VSUBS 0.00638f
C499 B.n454 VSUBS 0.00638f
C500 B.n455 VSUBS 0.00638f
C501 B.n456 VSUBS 0.00638f
C502 B.n457 VSUBS 0.00638f
C503 B.n458 VSUBS 0.00638f
C504 B.n459 VSUBS 0.00638f
C505 B.n460 VSUBS 0.00638f
C506 B.n461 VSUBS 0.00638f
C507 B.n462 VSUBS 0.00638f
C508 B.n463 VSUBS 0.00638f
C509 B.n464 VSUBS 0.00638f
C510 B.n465 VSUBS 0.00638f
C511 B.n466 VSUBS 0.00638f
C512 B.n467 VSUBS 0.00638f
C513 B.n468 VSUBS 0.00638f
C514 B.n469 VSUBS 0.00638f
C515 B.n470 VSUBS 0.00638f
C516 B.n471 VSUBS 0.00638f
C517 B.n472 VSUBS 0.00638f
C518 B.n473 VSUBS 0.00638f
C519 B.n474 VSUBS 0.00638f
C520 B.n475 VSUBS 0.00638f
C521 B.n476 VSUBS 0.00638f
C522 B.n477 VSUBS 0.00638f
C523 B.n478 VSUBS 0.00638f
C524 B.n479 VSUBS 0.00638f
C525 B.n480 VSUBS 0.00638f
C526 B.n481 VSUBS 0.00638f
C527 B.n482 VSUBS 0.00638f
C528 B.n483 VSUBS 0.00638f
C529 B.n484 VSUBS 0.00638f
C530 B.n485 VSUBS 0.00638f
C531 B.n486 VSUBS 0.00638f
C532 B.n487 VSUBS 0.00638f
C533 B.n488 VSUBS 0.00638f
C534 B.n489 VSUBS 0.00638f
C535 B.n490 VSUBS 0.00638f
C536 B.n491 VSUBS 0.00638f
C537 B.n492 VSUBS 0.00638f
C538 B.n493 VSUBS 0.00638f
C539 B.n494 VSUBS 0.00638f
C540 B.n495 VSUBS 0.00638f
C541 B.n496 VSUBS 0.00638f
C542 B.n497 VSUBS 0.00638f
C543 B.n498 VSUBS 0.00638f
C544 B.n499 VSUBS 0.00638f
C545 B.n500 VSUBS 0.00638f
C546 B.n501 VSUBS 0.00638f
C547 B.n502 VSUBS 0.00638f
C548 B.n503 VSUBS 0.00638f
C549 B.n504 VSUBS 0.00638f
C550 B.n505 VSUBS 0.00638f
C551 B.n506 VSUBS 0.00638f
C552 B.n507 VSUBS 0.00638f
C553 B.n508 VSUBS 0.00638f
C554 B.n509 VSUBS 0.00638f
C555 B.n510 VSUBS 0.00638f
C556 B.n511 VSUBS 0.00638f
C557 B.n512 VSUBS 0.00638f
C558 B.n513 VSUBS 0.00638f
C559 B.n514 VSUBS 0.00638f
C560 B.n515 VSUBS 0.00638f
C561 B.n516 VSUBS 0.00638f
C562 B.n517 VSUBS 0.00638f
C563 B.n518 VSUBS 0.00638f
C564 B.n519 VSUBS 0.01415f
C565 B.n520 VSUBS 0.01456f
C566 B.n521 VSUBS 0.01456f
C567 B.n522 VSUBS 0.00638f
C568 B.n523 VSUBS 0.00638f
C569 B.n524 VSUBS 0.00638f
C570 B.n525 VSUBS 0.00638f
C571 B.n526 VSUBS 0.00638f
C572 B.n527 VSUBS 0.00638f
C573 B.n528 VSUBS 0.00638f
C574 B.n529 VSUBS 0.00638f
C575 B.n530 VSUBS 0.00638f
C576 B.n531 VSUBS 0.00638f
C577 B.n532 VSUBS 0.00638f
C578 B.n533 VSUBS 0.00638f
C579 B.n534 VSUBS 0.00638f
C580 B.n535 VSUBS 0.00638f
C581 B.n536 VSUBS 0.00638f
C582 B.n537 VSUBS 0.00638f
C583 B.n538 VSUBS 0.00638f
C584 B.n539 VSUBS 0.00638f
C585 B.n540 VSUBS 0.00638f
C586 B.n541 VSUBS 0.00638f
C587 B.n542 VSUBS 0.00638f
C588 B.n543 VSUBS 0.00638f
C589 B.n544 VSUBS 0.00638f
C590 B.n545 VSUBS 0.00638f
C591 B.n546 VSUBS 0.00638f
C592 B.n547 VSUBS 0.00638f
C593 B.n548 VSUBS 0.00638f
C594 B.n549 VSUBS 0.00638f
C595 B.n550 VSUBS 0.00638f
C596 B.n551 VSUBS 0.00638f
C597 B.n552 VSUBS 0.00638f
C598 B.n553 VSUBS 0.00638f
C599 B.n554 VSUBS 0.00638f
C600 B.n555 VSUBS 0.00638f
C601 B.n556 VSUBS 0.00638f
C602 B.n557 VSUBS 0.00638f
C603 B.n558 VSUBS 0.00638f
C604 B.n559 VSUBS 0.00638f
C605 B.n560 VSUBS 0.00638f
C606 B.n561 VSUBS 0.00638f
C607 B.n562 VSUBS 0.00638f
C608 B.n563 VSUBS 0.00638f
C609 B.n564 VSUBS 0.00638f
C610 B.n565 VSUBS 0.00638f
C611 B.n566 VSUBS 0.00638f
C612 B.n567 VSUBS 0.00638f
C613 B.n568 VSUBS 0.00638f
C614 B.n569 VSUBS 0.00638f
C615 B.n570 VSUBS 0.00638f
C616 B.n571 VSUBS 0.00638f
C617 B.n572 VSUBS 0.00638f
C618 B.n573 VSUBS 0.00638f
C619 B.n574 VSUBS 0.00638f
C620 B.n575 VSUBS 0.00638f
C621 B.n576 VSUBS 0.00638f
C622 B.n577 VSUBS 0.00638f
C623 B.n578 VSUBS 0.00638f
C624 B.n579 VSUBS 0.00638f
C625 B.n580 VSUBS 0.00638f
C626 B.n581 VSUBS 0.00638f
C627 B.n582 VSUBS 0.00638f
C628 B.n583 VSUBS 0.00638f
C629 B.n584 VSUBS 0.00638f
C630 B.n585 VSUBS 0.00638f
C631 B.n586 VSUBS 0.00638f
C632 B.n587 VSUBS 0.00638f
C633 B.n588 VSUBS 0.00638f
C634 B.n589 VSUBS 0.00638f
C635 B.n590 VSUBS 0.00638f
C636 B.n591 VSUBS 0.00638f
C637 B.n592 VSUBS 0.00638f
C638 B.n593 VSUBS 0.00638f
C639 B.n594 VSUBS 0.00638f
C640 B.n595 VSUBS 0.00638f
C641 B.n596 VSUBS 0.00638f
C642 B.n597 VSUBS 0.00638f
C643 B.n598 VSUBS 0.00638f
C644 B.n599 VSUBS 0.00638f
C645 B.n600 VSUBS 0.00638f
C646 B.n601 VSUBS 0.00441f
C647 B.n602 VSUBS 0.00638f
C648 B.n603 VSUBS 0.00638f
C649 B.n604 VSUBS 0.00516f
C650 B.n605 VSUBS 0.00638f
C651 B.n606 VSUBS 0.00638f
C652 B.n607 VSUBS 0.00638f
C653 B.n608 VSUBS 0.00638f
C654 B.n609 VSUBS 0.00638f
C655 B.n610 VSUBS 0.00638f
C656 B.n611 VSUBS 0.00638f
C657 B.n612 VSUBS 0.00638f
C658 B.n613 VSUBS 0.00638f
C659 B.n614 VSUBS 0.00638f
C660 B.n615 VSUBS 0.00638f
C661 B.n616 VSUBS 0.00516f
C662 B.n617 VSUBS 0.014781f
C663 B.n618 VSUBS 0.00441f
C664 B.n619 VSUBS 0.00638f
C665 B.n620 VSUBS 0.00638f
C666 B.n621 VSUBS 0.00638f
C667 B.n622 VSUBS 0.00638f
C668 B.n623 VSUBS 0.00638f
C669 B.n624 VSUBS 0.00638f
C670 B.n625 VSUBS 0.00638f
C671 B.n626 VSUBS 0.00638f
C672 B.n627 VSUBS 0.00638f
C673 B.n628 VSUBS 0.00638f
C674 B.n629 VSUBS 0.00638f
C675 B.n630 VSUBS 0.00638f
C676 B.n631 VSUBS 0.00638f
C677 B.n632 VSUBS 0.00638f
C678 B.n633 VSUBS 0.00638f
C679 B.n634 VSUBS 0.00638f
C680 B.n635 VSUBS 0.00638f
C681 B.n636 VSUBS 0.00638f
C682 B.n637 VSUBS 0.00638f
C683 B.n638 VSUBS 0.00638f
C684 B.n639 VSUBS 0.00638f
C685 B.n640 VSUBS 0.00638f
C686 B.n641 VSUBS 0.00638f
C687 B.n642 VSUBS 0.00638f
C688 B.n643 VSUBS 0.00638f
C689 B.n644 VSUBS 0.00638f
C690 B.n645 VSUBS 0.00638f
C691 B.n646 VSUBS 0.00638f
C692 B.n647 VSUBS 0.00638f
C693 B.n648 VSUBS 0.00638f
C694 B.n649 VSUBS 0.00638f
C695 B.n650 VSUBS 0.00638f
C696 B.n651 VSUBS 0.00638f
C697 B.n652 VSUBS 0.00638f
C698 B.n653 VSUBS 0.00638f
C699 B.n654 VSUBS 0.00638f
C700 B.n655 VSUBS 0.00638f
C701 B.n656 VSUBS 0.00638f
C702 B.n657 VSUBS 0.00638f
C703 B.n658 VSUBS 0.00638f
C704 B.n659 VSUBS 0.00638f
C705 B.n660 VSUBS 0.00638f
C706 B.n661 VSUBS 0.00638f
C707 B.n662 VSUBS 0.00638f
C708 B.n663 VSUBS 0.00638f
C709 B.n664 VSUBS 0.00638f
C710 B.n665 VSUBS 0.00638f
C711 B.n666 VSUBS 0.00638f
C712 B.n667 VSUBS 0.00638f
C713 B.n668 VSUBS 0.00638f
C714 B.n669 VSUBS 0.00638f
C715 B.n670 VSUBS 0.00638f
C716 B.n671 VSUBS 0.00638f
C717 B.n672 VSUBS 0.00638f
C718 B.n673 VSUBS 0.00638f
C719 B.n674 VSUBS 0.00638f
C720 B.n675 VSUBS 0.00638f
C721 B.n676 VSUBS 0.00638f
C722 B.n677 VSUBS 0.00638f
C723 B.n678 VSUBS 0.00638f
C724 B.n679 VSUBS 0.00638f
C725 B.n680 VSUBS 0.00638f
C726 B.n681 VSUBS 0.00638f
C727 B.n682 VSUBS 0.00638f
C728 B.n683 VSUBS 0.00638f
C729 B.n684 VSUBS 0.00638f
C730 B.n685 VSUBS 0.00638f
C731 B.n686 VSUBS 0.00638f
C732 B.n687 VSUBS 0.00638f
C733 B.n688 VSUBS 0.00638f
C734 B.n689 VSUBS 0.00638f
C735 B.n690 VSUBS 0.00638f
C736 B.n691 VSUBS 0.00638f
C737 B.n692 VSUBS 0.00638f
C738 B.n693 VSUBS 0.00638f
C739 B.n694 VSUBS 0.00638f
C740 B.n695 VSUBS 0.00638f
C741 B.n696 VSUBS 0.00638f
C742 B.n697 VSUBS 0.00638f
C743 B.n698 VSUBS 0.00638f
C744 B.n699 VSUBS 0.01456f
C745 B.n700 VSUBS 0.01415f
C746 B.n701 VSUBS 0.01415f
C747 B.n702 VSUBS 0.00638f
C748 B.n703 VSUBS 0.00638f
C749 B.n704 VSUBS 0.00638f
C750 B.n705 VSUBS 0.00638f
C751 B.n706 VSUBS 0.00638f
C752 B.n707 VSUBS 0.00638f
C753 B.n708 VSUBS 0.00638f
C754 B.n709 VSUBS 0.00638f
C755 B.n710 VSUBS 0.00638f
C756 B.n711 VSUBS 0.00638f
C757 B.n712 VSUBS 0.00638f
C758 B.n713 VSUBS 0.00638f
C759 B.n714 VSUBS 0.00638f
C760 B.n715 VSUBS 0.00638f
C761 B.n716 VSUBS 0.00638f
C762 B.n717 VSUBS 0.00638f
C763 B.n718 VSUBS 0.00638f
C764 B.n719 VSUBS 0.00638f
C765 B.n720 VSUBS 0.00638f
C766 B.n721 VSUBS 0.00638f
C767 B.n722 VSUBS 0.00638f
C768 B.n723 VSUBS 0.00638f
C769 B.n724 VSUBS 0.00638f
C770 B.n725 VSUBS 0.00638f
C771 B.n726 VSUBS 0.00638f
C772 B.n727 VSUBS 0.00638f
C773 B.n728 VSUBS 0.00638f
C774 B.n729 VSUBS 0.00638f
C775 B.n730 VSUBS 0.00638f
C776 B.n731 VSUBS 0.00638f
C777 B.n732 VSUBS 0.00638f
C778 B.n733 VSUBS 0.00638f
C779 B.n734 VSUBS 0.00638f
C780 B.n735 VSUBS 0.00638f
C781 B.n736 VSUBS 0.00638f
C782 B.n737 VSUBS 0.00638f
C783 B.n738 VSUBS 0.00638f
C784 B.n739 VSUBS 0.00638f
C785 B.n740 VSUBS 0.00638f
C786 B.n741 VSUBS 0.00638f
C787 B.n742 VSUBS 0.00638f
C788 B.n743 VSUBS 0.00638f
C789 B.n744 VSUBS 0.00638f
C790 B.n745 VSUBS 0.00638f
C791 B.n746 VSUBS 0.00638f
C792 B.n747 VSUBS 0.008325f
C793 B.n748 VSUBS 0.008869f
C794 B.n749 VSUBS 0.017636f
C795 VDD1.t1 VSUBS 3.99444f
C796 VDD1.t0 VSUBS 5.13876f
C797 VTAIL.t2 VSUBS 3.84124f
C798 VTAIL.n0 VSUBS 3.34719f
C799 VTAIL.t0 VSUBS 3.84125f
C800 VTAIL.n1 VSUBS 3.42472f
C801 VTAIL.t3 VSUBS 3.84124f
C802 VTAIL.n2 VSUBS 3.09279f
C803 VTAIL.t1 VSUBS 3.84124f
C804 VTAIL.n3 VSUBS 2.96034f
C805 VP.t0 VSUBS 6.6548f
C806 VP.t1 VSUBS 5.71041f
C807 VP.n0 VSUBS 6.00626f
.ends

