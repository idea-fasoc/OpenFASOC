* NGSPICE file created from diff_pair_sample_0678.ext - technology: sky130A

.subckt diff_pair_sample_0678 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=2.028 pd=11.18 as=0 ps=0 w=5.2 l=1.22
X1 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=2.028 pd=11.18 as=0 ps=0 w=5.2 l=1.22
X2 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.028 pd=11.18 as=0 ps=0 w=5.2 l=1.22
X3 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.028 pd=11.18 as=0 ps=0 w=5.2 l=1.22
X4 VDD1.t1 VP.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.028 pd=11.18 as=2.028 ps=11.18 w=5.2 l=1.22
X5 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.028 pd=11.18 as=2.028 ps=11.18 w=5.2 l=1.22
X6 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.028 pd=11.18 as=2.028 ps=11.18 w=5.2 l=1.22
X7 VDD1.t0 VP.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.028 pd=11.18 as=2.028 ps=11.18 w=5.2 l=1.22
R0 B.n415 B.n414 585
R1 B.n416 B.n415 585
R2 B.n170 B.n61 585
R3 B.n169 B.n168 585
R4 B.n167 B.n166 585
R5 B.n165 B.n164 585
R6 B.n163 B.n162 585
R7 B.n161 B.n160 585
R8 B.n159 B.n158 585
R9 B.n157 B.n156 585
R10 B.n155 B.n154 585
R11 B.n153 B.n152 585
R12 B.n151 B.n150 585
R13 B.n149 B.n148 585
R14 B.n147 B.n146 585
R15 B.n145 B.n144 585
R16 B.n143 B.n142 585
R17 B.n141 B.n140 585
R18 B.n139 B.n138 585
R19 B.n137 B.n136 585
R20 B.n135 B.n134 585
R21 B.n133 B.n132 585
R22 B.n131 B.n130 585
R23 B.n128 B.n127 585
R24 B.n126 B.n125 585
R25 B.n124 B.n123 585
R26 B.n122 B.n121 585
R27 B.n120 B.n119 585
R28 B.n118 B.n117 585
R29 B.n116 B.n115 585
R30 B.n114 B.n113 585
R31 B.n112 B.n111 585
R32 B.n110 B.n109 585
R33 B.n108 B.n107 585
R34 B.n106 B.n105 585
R35 B.n104 B.n103 585
R36 B.n102 B.n101 585
R37 B.n100 B.n99 585
R38 B.n98 B.n97 585
R39 B.n96 B.n95 585
R40 B.n94 B.n93 585
R41 B.n92 B.n91 585
R42 B.n90 B.n89 585
R43 B.n88 B.n87 585
R44 B.n86 B.n85 585
R45 B.n84 B.n83 585
R46 B.n82 B.n81 585
R47 B.n80 B.n79 585
R48 B.n78 B.n77 585
R49 B.n76 B.n75 585
R50 B.n74 B.n73 585
R51 B.n72 B.n71 585
R52 B.n70 B.n69 585
R53 B.n68 B.n67 585
R54 B.n413 B.n34 585
R55 B.n417 B.n34 585
R56 B.n412 B.n33 585
R57 B.n418 B.n33 585
R58 B.n411 B.n410 585
R59 B.n410 B.n29 585
R60 B.n409 B.n28 585
R61 B.n424 B.n28 585
R62 B.n408 B.n27 585
R63 B.n425 B.n27 585
R64 B.n407 B.n26 585
R65 B.n426 B.n26 585
R66 B.n406 B.n405 585
R67 B.n405 B.n22 585
R68 B.n404 B.n21 585
R69 B.n432 B.n21 585
R70 B.n403 B.n20 585
R71 B.n433 B.n20 585
R72 B.n402 B.n19 585
R73 B.n434 B.n19 585
R74 B.n401 B.n400 585
R75 B.n400 B.n15 585
R76 B.n399 B.n14 585
R77 B.n440 B.n14 585
R78 B.n398 B.n13 585
R79 B.n441 B.n13 585
R80 B.n397 B.n12 585
R81 B.n442 B.n12 585
R82 B.n396 B.n395 585
R83 B.n395 B.n8 585
R84 B.n394 B.n7 585
R85 B.n448 B.n7 585
R86 B.n393 B.n6 585
R87 B.n449 B.n6 585
R88 B.n392 B.n5 585
R89 B.n450 B.n5 585
R90 B.n391 B.n390 585
R91 B.n390 B.n4 585
R92 B.n389 B.n171 585
R93 B.n389 B.n388 585
R94 B.n379 B.n172 585
R95 B.n173 B.n172 585
R96 B.n381 B.n380 585
R97 B.n382 B.n381 585
R98 B.n378 B.n178 585
R99 B.n178 B.n177 585
R100 B.n377 B.n376 585
R101 B.n376 B.n375 585
R102 B.n180 B.n179 585
R103 B.n181 B.n180 585
R104 B.n368 B.n367 585
R105 B.n369 B.n368 585
R106 B.n366 B.n186 585
R107 B.n186 B.n185 585
R108 B.n365 B.n364 585
R109 B.n364 B.n363 585
R110 B.n188 B.n187 585
R111 B.n189 B.n188 585
R112 B.n356 B.n355 585
R113 B.n357 B.n356 585
R114 B.n354 B.n194 585
R115 B.n194 B.n193 585
R116 B.n353 B.n352 585
R117 B.n352 B.n351 585
R118 B.n196 B.n195 585
R119 B.n197 B.n196 585
R120 B.n344 B.n343 585
R121 B.n345 B.n344 585
R122 B.n342 B.n202 585
R123 B.n202 B.n201 585
R124 B.n336 B.n335 585
R125 B.n334 B.n230 585
R126 B.n333 B.n229 585
R127 B.n338 B.n229 585
R128 B.n332 B.n331 585
R129 B.n330 B.n329 585
R130 B.n328 B.n327 585
R131 B.n326 B.n325 585
R132 B.n324 B.n323 585
R133 B.n322 B.n321 585
R134 B.n320 B.n319 585
R135 B.n318 B.n317 585
R136 B.n316 B.n315 585
R137 B.n314 B.n313 585
R138 B.n312 B.n311 585
R139 B.n310 B.n309 585
R140 B.n308 B.n307 585
R141 B.n306 B.n305 585
R142 B.n304 B.n303 585
R143 B.n302 B.n301 585
R144 B.n300 B.n299 585
R145 B.n298 B.n297 585
R146 B.n296 B.n295 585
R147 B.n293 B.n292 585
R148 B.n291 B.n290 585
R149 B.n289 B.n288 585
R150 B.n287 B.n286 585
R151 B.n285 B.n284 585
R152 B.n283 B.n282 585
R153 B.n281 B.n280 585
R154 B.n279 B.n278 585
R155 B.n277 B.n276 585
R156 B.n275 B.n274 585
R157 B.n273 B.n272 585
R158 B.n271 B.n270 585
R159 B.n269 B.n268 585
R160 B.n267 B.n266 585
R161 B.n265 B.n264 585
R162 B.n263 B.n262 585
R163 B.n261 B.n260 585
R164 B.n259 B.n258 585
R165 B.n257 B.n256 585
R166 B.n255 B.n254 585
R167 B.n253 B.n252 585
R168 B.n251 B.n250 585
R169 B.n249 B.n248 585
R170 B.n247 B.n246 585
R171 B.n245 B.n244 585
R172 B.n243 B.n242 585
R173 B.n241 B.n240 585
R174 B.n239 B.n238 585
R175 B.n237 B.n236 585
R176 B.n204 B.n203 585
R177 B.n341 B.n340 585
R178 B.n200 B.n199 585
R179 B.n201 B.n200 585
R180 B.n347 B.n346 585
R181 B.n346 B.n345 585
R182 B.n348 B.n198 585
R183 B.n198 B.n197 585
R184 B.n350 B.n349 585
R185 B.n351 B.n350 585
R186 B.n192 B.n191 585
R187 B.n193 B.n192 585
R188 B.n359 B.n358 585
R189 B.n358 B.n357 585
R190 B.n360 B.n190 585
R191 B.n190 B.n189 585
R192 B.n362 B.n361 585
R193 B.n363 B.n362 585
R194 B.n184 B.n183 585
R195 B.n185 B.n184 585
R196 B.n371 B.n370 585
R197 B.n370 B.n369 585
R198 B.n372 B.n182 585
R199 B.n182 B.n181 585
R200 B.n374 B.n373 585
R201 B.n375 B.n374 585
R202 B.n176 B.n175 585
R203 B.n177 B.n176 585
R204 B.n384 B.n383 585
R205 B.n383 B.n382 585
R206 B.n385 B.n174 585
R207 B.n174 B.n173 585
R208 B.n387 B.n386 585
R209 B.n388 B.n387 585
R210 B.n2 B.n0 585
R211 B.n4 B.n2 585
R212 B.n3 B.n1 585
R213 B.n449 B.n3 585
R214 B.n447 B.n446 585
R215 B.n448 B.n447 585
R216 B.n445 B.n9 585
R217 B.n9 B.n8 585
R218 B.n444 B.n443 585
R219 B.n443 B.n442 585
R220 B.n11 B.n10 585
R221 B.n441 B.n11 585
R222 B.n439 B.n438 585
R223 B.n440 B.n439 585
R224 B.n437 B.n16 585
R225 B.n16 B.n15 585
R226 B.n436 B.n435 585
R227 B.n435 B.n434 585
R228 B.n18 B.n17 585
R229 B.n433 B.n18 585
R230 B.n431 B.n430 585
R231 B.n432 B.n431 585
R232 B.n429 B.n23 585
R233 B.n23 B.n22 585
R234 B.n428 B.n427 585
R235 B.n427 B.n426 585
R236 B.n25 B.n24 585
R237 B.n425 B.n25 585
R238 B.n423 B.n422 585
R239 B.n424 B.n423 585
R240 B.n421 B.n30 585
R241 B.n30 B.n29 585
R242 B.n420 B.n419 585
R243 B.n419 B.n418 585
R244 B.n32 B.n31 585
R245 B.n417 B.n32 585
R246 B.n452 B.n451 585
R247 B.n451 B.n450 585
R248 B.n336 B.n200 521.33
R249 B.n67 B.n32 521.33
R250 B.n340 B.n202 521.33
R251 B.n415 B.n34 521.33
R252 B.n233 B.t9 306.942
R253 B.n231 B.t13 306.942
R254 B.n64 B.t6 306.942
R255 B.n62 B.t2 306.942
R256 B.n416 B.n60 256.663
R257 B.n416 B.n59 256.663
R258 B.n416 B.n58 256.663
R259 B.n416 B.n57 256.663
R260 B.n416 B.n56 256.663
R261 B.n416 B.n55 256.663
R262 B.n416 B.n54 256.663
R263 B.n416 B.n53 256.663
R264 B.n416 B.n52 256.663
R265 B.n416 B.n51 256.663
R266 B.n416 B.n50 256.663
R267 B.n416 B.n49 256.663
R268 B.n416 B.n48 256.663
R269 B.n416 B.n47 256.663
R270 B.n416 B.n46 256.663
R271 B.n416 B.n45 256.663
R272 B.n416 B.n44 256.663
R273 B.n416 B.n43 256.663
R274 B.n416 B.n42 256.663
R275 B.n416 B.n41 256.663
R276 B.n416 B.n40 256.663
R277 B.n416 B.n39 256.663
R278 B.n416 B.n38 256.663
R279 B.n416 B.n37 256.663
R280 B.n416 B.n36 256.663
R281 B.n416 B.n35 256.663
R282 B.n338 B.n337 256.663
R283 B.n338 B.n205 256.663
R284 B.n338 B.n206 256.663
R285 B.n338 B.n207 256.663
R286 B.n338 B.n208 256.663
R287 B.n338 B.n209 256.663
R288 B.n338 B.n210 256.663
R289 B.n338 B.n211 256.663
R290 B.n338 B.n212 256.663
R291 B.n338 B.n213 256.663
R292 B.n338 B.n214 256.663
R293 B.n338 B.n215 256.663
R294 B.n338 B.n216 256.663
R295 B.n338 B.n217 256.663
R296 B.n338 B.n218 256.663
R297 B.n338 B.n219 256.663
R298 B.n338 B.n220 256.663
R299 B.n338 B.n221 256.663
R300 B.n338 B.n222 256.663
R301 B.n338 B.n223 256.663
R302 B.n338 B.n224 256.663
R303 B.n338 B.n225 256.663
R304 B.n338 B.n226 256.663
R305 B.n338 B.n227 256.663
R306 B.n338 B.n228 256.663
R307 B.n339 B.n338 256.663
R308 B.n233 B.t12 195.083
R309 B.n62 B.t4 195.083
R310 B.n231 B.t15 195.083
R311 B.n64 B.t7 195.083
R312 B.n234 B.t11 165.023
R313 B.n63 B.t5 165.023
R314 B.n232 B.t14 165.023
R315 B.n65 B.t8 165.023
R316 B.n346 B.n200 163.367
R317 B.n346 B.n198 163.367
R318 B.n350 B.n198 163.367
R319 B.n350 B.n192 163.367
R320 B.n358 B.n192 163.367
R321 B.n358 B.n190 163.367
R322 B.n362 B.n190 163.367
R323 B.n362 B.n184 163.367
R324 B.n370 B.n184 163.367
R325 B.n370 B.n182 163.367
R326 B.n374 B.n182 163.367
R327 B.n374 B.n176 163.367
R328 B.n383 B.n176 163.367
R329 B.n383 B.n174 163.367
R330 B.n387 B.n174 163.367
R331 B.n387 B.n2 163.367
R332 B.n451 B.n2 163.367
R333 B.n451 B.n3 163.367
R334 B.n447 B.n3 163.367
R335 B.n447 B.n9 163.367
R336 B.n443 B.n9 163.367
R337 B.n443 B.n11 163.367
R338 B.n439 B.n11 163.367
R339 B.n439 B.n16 163.367
R340 B.n435 B.n16 163.367
R341 B.n435 B.n18 163.367
R342 B.n431 B.n18 163.367
R343 B.n431 B.n23 163.367
R344 B.n427 B.n23 163.367
R345 B.n427 B.n25 163.367
R346 B.n423 B.n25 163.367
R347 B.n423 B.n30 163.367
R348 B.n419 B.n30 163.367
R349 B.n419 B.n32 163.367
R350 B.n230 B.n229 163.367
R351 B.n331 B.n229 163.367
R352 B.n329 B.n328 163.367
R353 B.n325 B.n324 163.367
R354 B.n321 B.n320 163.367
R355 B.n317 B.n316 163.367
R356 B.n313 B.n312 163.367
R357 B.n309 B.n308 163.367
R358 B.n305 B.n304 163.367
R359 B.n301 B.n300 163.367
R360 B.n297 B.n296 163.367
R361 B.n292 B.n291 163.367
R362 B.n288 B.n287 163.367
R363 B.n284 B.n283 163.367
R364 B.n280 B.n279 163.367
R365 B.n276 B.n275 163.367
R366 B.n272 B.n271 163.367
R367 B.n268 B.n267 163.367
R368 B.n264 B.n263 163.367
R369 B.n260 B.n259 163.367
R370 B.n256 B.n255 163.367
R371 B.n252 B.n251 163.367
R372 B.n248 B.n247 163.367
R373 B.n244 B.n243 163.367
R374 B.n240 B.n239 163.367
R375 B.n236 B.n204 163.367
R376 B.n344 B.n202 163.367
R377 B.n344 B.n196 163.367
R378 B.n352 B.n196 163.367
R379 B.n352 B.n194 163.367
R380 B.n356 B.n194 163.367
R381 B.n356 B.n188 163.367
R382 B.n364 B.n188 163.367
R383 B.n364 B.n186 163.367
R384 B.n368 B.n186 163.367
R385 B.n368 B.n180 163.367
R386 B.n376 B.n180 163.367
R387 B.n376 B.n178 163.367
R388 B.n381 B.n178 163.367
R389 B.n381 B.n172 163.367
R390 B.n389 B.n172 163.367
R391 B.n390 B.n389 163.367
R392 B.n390 B.n5 163.367
R393 B.n6 B.n5 163.367
R394 B.n7 B.n6 163.367
R395 B.n395 B.n7 163.367
R396 B.n395 B.n12 163.367
R397 B.n13 B.n12 163.367
R398 B.n14 B.n13 163.367
R399 B.n400 B.n14 163.367
R400 B.n400 B.n19 163.367
R401 B.n20 B.n19 163.367
R402 B.n21 B.n20 163.367
R403 B.n405 B.n21 163.367
R404 B.n405 B.n26 163.367
R405 B.n27 B.n26 163.367
R406 B.n28 B.n27 163.367
R407 B.n410 B.n28 163.367
R408 B.n410 B.n33 163.367
R409 B.n34 B.n33 163.367
R410 B.n71 B.n70 163.367
R411 B.n75 B.n74 163.367
R412 B.n79 B.n78 163.367
R413 B.n83 B.n82 163.367
R414 B.n87 B.n86 163.367
R415 B.n91 B.n90 163.367
R416 B.n95 B.n94 163.367
R417 B.n99 B.n98 163.367
R418 B.n103 B.n102 163.367
R419 B.n107 B.n106 163.367
R420 B.n111 B.n110 163.367
R421 B.n115 B.n114 163.367
R422 B.n119 B.n118 163.367
R423 B.n123 B.n122 163.367
R424 B.n127 B.n126 163.367
R425 B.n132 B.n131 163.367
R426 B.n136 B.n135 163.367
R427 B.n140 B.n139 163.367
R428 B.n144 B.n143 163.367
R429 B.n148 B.n147 163.367
R430 B.n152 B.n151 163.367
R431 B.n156 B.n155 163.367
R432 B.n160 B.n159 163.367
R433 B.n164 B.n163 163.367
R434 B.n168 B.n167 163.367
R435 B.n415 B.n61 163.367
R436 B.n338 B.n201 145.968
R437 B.n417 B.n416 145.968
R438 B.n337 B.n336 71.676
R439 B.n331 B.n205 71.676
R440 B.n328 B.n206 71.676
R441 B.n324 B.n207 71.676
R442 B.n320 B.n208 71.676
R443 B.n316 B.n209 71.676
R444 B.n312 B.n210 71.676
R445 B.n308 B.n211 71.676
R446 B.n304 B.n212 71.676
R447 B.n300 B.n213 71.676
R448 B.n296 B.n214 71.676
R449 B.n291 B.n215 71.676
R450 B.n287 B.n216 71.676
R451 B.n283 B.n217 71.676
R452 B.n279 B.n218 71.676
R453 B.n275 B.n219 71.676
R454 B.n271 B.n220 71.676
R455 B.n267 B.n221 71.676
R456 B.n263 B.n222 71.676
R457 B.n259 B.n223 71.676
R458 B.n255 B.n224 71.676
R459 B.n251 B.n225 71.676
R460 B.n247 B.n226 71.676
R461 B.n243 B.n227 71.676
R462 B.n239 B.n228 71.676
R463 B.n339 B.n204 71.676
R464 B.n67 B.n35 71.676
R465 B.n71 B.n36 71.676
R466 B.n75 B.n37 71.676
R467 B.n79 B.n38 71.676
R468 B.n83 B.n39 71.676
R469 B.n87 B.n40 71.676
R470 B.n91 B.n41 71.676
R471 B.n95 B.n42 71.676
R472 B.n99 B.n43 71.676
R473 B.n103 B.n44 71.676
R474 B.n107 B.n45 71.676
R475 B.n111 B.n46 71.676
R476 B.n115 B.n47 71.676
R477 B.n119 B.n48 71.676
R478 B.n123 B.n49 71.676
R479 B.n127 B.n50 71.676
R480 B.n132 B.n51 71.676
R481 B.n136 B.n52 71.676
R482 B.n140 B.n53 71.676
R483 B.n144 B.n54 71.676
R484 B.n148 B.n55 71.676
R485 B.n152 B.n56 71.676
R486 B.n156 B.n57 71.676
R487 B.n160 B.n58 71.676
R488 B.n164 B.n59 71.676
R489 B.n168 B.n60 71.676
R490 B.n61 B.n60 71.676
R491 B.n167 B.n59 71.676
R492 B.n163 B.n58 71.676
R493 B.n159 B.n57 71.676
R494 B.n155 B.n56 71.676
R495 B.n151 B.n55 71.676
R496 B.n147 B.n54 71.676
R497 B.n143 B.n53 71.676
R498 B.n139 B.n52 71.676
R499 B.n135 B.n51 71.676
R500 B.n131 B.n50 71.676
R501 B.n126 B.n49 71.676
R502 B.n122 B.n48 71.676
R503 B.n118 B.n47 71.676
R504 B.n114 B.n46 71.676
R505 B.n110 B.n45 71.676
R506 B.n106 B.n44 71.676
R507 B.n102 B.n43 71.676
R508 B.n98 B.n42 71.676
R509 B.n94 B.n41 71.676
R510 B.n90 B.n40 71.676
R511 B.n86 B.n39 71.676
R512 B.n82 B.n38 71.676
R513 B.n78 B.n37 71.676
R514 B.n74 B.n36 71.676
R515 B.n70 B.n35 71.676
R516 B.n337 B.n230 71.676
R517 B.n329 B.n205 71.676
R518 B.n325 B.n206 71.676
R519 B.n321 B.n207 71.676
R520 B.n317 B.n208 71.676
R521 B.n313 B.n209 71.676
R522 B.n309 B.n210 71.676
R523 B.n305 B.n211 71.676
R524 B.n301 B.n212 71.676
R525 B.n297 B.n213 71.676
R526 B.n292 B.n214 71.676
R527 B.n288 B.n215 71.676
R528 B.n284 B.n216 71.676
R529 B.n280 B.n217 71.676
R530 B.n276 B.n218 71.676
R531 B.n272 B.n219 71.676
R532 B.n268 B.n220 71.676
R533 B.n264 B.n221 71.676
R534 B.n260 B.n222 71.676
R535 B.n256 B.n223 71.676
R536 B.n252 B.n224 71.676
R537 B.n248 B.n225 71.676
R538 B.n244 B.n226 71.676
R539 B.n240 B.n227 71.676
R540 B.n236 B.n228 71.676
R541 B.n340 B.n339 71.676
R542 B.n345 B.n201 71.4086
R543 B.n345 B.n197 71.4086
R544 B.n351 B.n197 71.4086
R545 B.n351 B.n193 71.4086
R546 B.n357 B.n193 71.4086
R547 B.n363 B.n189 71.4086
R548 B.n363 B.n185 71.4086
R549 B.n369 B.n185 71.4086
R550 B.n369 B.n181 71.4086
R551 B.n375 B.n181 71.4086
R552 B.n375 B.n177 71.4086
R553 B.n382 B.n177 71.4086
R554 B.n388 B.n173 71.4086
R555 B.n388 B.n4 71.4086
R556 B.n450 B.n4 71.4086
R557 B.n450 B.n449 71.4086
R558 B.n449 B.n448 71.4086
R559 B.n448 B.n8 71.4086
R560 B.n442 B.n441 71.4086
R561 B.n441 B.n440 71.4086
R562 B.n440 B.n15 71.4086
R563 B.n434 B.n15 71.4086
R564 B.n434 B.n433 71.4086
R565 B.n433 B.n432 71.4086
R566 B.n432 B.n22 71.4086
R567 B.n426 B.n425 71.4086
R568 B.n425 B.n424 71.4086
R569 B.n424 B.n29 71.4086
R570 B.n418 B.n29 71.4086
R571 B.n418 B.n417 71.4086
R572 B.t0 B.n173 63.0077
R573 B.t1 B.n8 63.0077
R574 B.n235 B.n234 59.5399
R575 B.n294 B.n232 59.5399
R576 B.n66 B.n65 59.5399
R577 B.n129 B.n63 59.5399
R578 B.t10 B.n189 46.2057
R579 B.t3 B.n22 46.2057
R580 B.n68 B.n31 33.8737
R581 B.n414 B.n413 33.8737
R582 B.n342 B.n341 33.8737
R583 B.n335 B.n199 33.8737
R584 B.n234 B.n233 30.0611
R585 B.n232 B.n231 30.0611
R586 B.n65 B.n64 30.0611
R587 B.n63 B.n62 30.0611
R588 B.n357 B.t10 25.2034
R589 B.n426 B.t3 25.2034
R590 B B.n452 18.0485
R591 B.n69 B.n68 10.6151
R592 B.n72 B.n69 10.6151
R593 B.n73 B.n72 10.6151
R594 B.n76 B.n73 10.6151
R595 B.n77 B.n76 10.6151
R596 B.n80 B.n77 10.6151
R597 B.n81 B.n80 10.6151
R598 B.n84 B.n81 10.6151
R599 B.n85 B.n84 10.6151
R600 B.n88 B.n85 10.6151
R601 B.n89 B.n88 10.6151
R602 B.n92 B.n89 10.6151
R603 B.n93 B.n92 10.6151
R604 B.n96 B.n93 10.6151
R605 B.n97 B.n96 10.6151
R606 B.n100 B.n97 10.6151
R607 B.n101 B.n100 10.6151
R608 B.n104 B.n101 10.6151
R609 B.n105 B.n104 10.6151
R610 B.n108 B.n105 10.6151
R611 B.n109 B.n108 10.6151
R612 B.n113 B.n112 10.6151
R613 B.n116 B.n113 10.6151
R614 B.n117 B.n116 10.6151
R615 B.n120 B.n117 10.6151
R616 B.n121 B.n120 10.6151
R617 B.n124 B.n121 10.6151
R618 B.n125 B.n124 10.6151
R619 B.n128 B.n125 10.6151
R620 B.n133 B.n130 10.6151
R621 B.n134 B.n133 10.6151
R622 B.n137 B.n134 10.6151
R623 B.n138 B.n137 10.6151
R624 B.n141 B.n138 10.6151
R625 B.n142 B.n141 10.6151
R626 B.n145 B.n142 10.6151
R627 B.n146 B.n145 10.6151
R628 B.n149 B.n146 10.6151
R629 B.n150 B.n149 10.6151
R630 B.n153 B.n150 10.6151
R631 B.n154 B.n153 10.6151
R632 B.n157 B.n154 10.6151
R633 B.n158 B.n157 10.6151
R634 B.n161 B.n158 10.6151
R635 B.n162 B.n161 10.6151
R636 B.n165 B.n162 10.6151
R637 B.n166 B.n165 10.6151
R638 B.n169 B.n166 10.6151
R639 B.n170 B.n169 10.6151
R640 B.n414 B.n170 10.6151
R641 B.n343 B.n342 10.6151
R642 B.n343 B.n195 10.6151
R643 B.n353 B.n195 10.6151
R644 B.n354 B.n353 10.6151
R645 B.n355 B.n354 10.6151
R646 B.n355 B.n187 10.6151
R647 B.n365 B.n187 10.6151
R648 B.n366 B.n365 10.6151
R649 B.n367 B.n366 10.6151
R650 B.n367 B.n179 10.6151
R651 B.n377 B.n179 10.6151
R652 B.n378 B.n377 10.6151
R653 B.n380 B.n378 10.6151
R654 B.n380 B.n379 10.6151
R655 B.n379 B.n171 10.6151
R656 B.n391 B.n171 10.6151
R657 B.n392 B.n391 10.6151
R658 B.n393 B.n392 10.6151
R659 B.n394 B.n393 10.6151
R660 B.n396 B.n394 10.6151
R661 B.n397 B.n396 10.6151
R662 B.n398 B.n397 10.6151
R663 B.n399 B.n398 10.6151
R664 B.n401 B.n399 10.6151
R665 B.n402 B.n401 10.6151
R666 B.n403 B.n402 10.6151
R667 B.n404 B.n403 10.6151
R668 B.n406 B.n404 10.6151
R669 B.n407 B.n406 10.6151
R670 B.n408 B.n407 10.6151
R671 B.n409 B.n408 10.6151
R672 B.n411 B.n409 10.6151
R673 B.n412 B.n411 10.6151
R674 B.n413 B.n412 10.6151
R675 B.n335 B.n334 10.6151
R676 B.n334 B.n333 10.6151
R677 B.n333 B.n332 10.6151
R678 B.n332 B.n330 10.6151
R679 B.n330 B.n327 10.6151
R680 B.n327 B.n326 10.6151
R681 B.n326 B.n323 10.6151
R682 B.n323 B.n322 10.6151
R683 B.n322 B.n319 10.6151
R684 B.n319 B.n318 10.6151
R685 B.n318 B.n315 10.6151
R686 B.n315 B.n314 10.6151
R687 B.n314 B.n311 10.6151
R688 B.n311 B.n310 10.6151
R689 B.n310 B.n307 10.6151
R690 B.n307 B.n306 10.6151
R691 B.n306 B.n303 10.6151
R692 B.n303 B.n302 10.6151
R693 B.n302 B.n299 10.6151
R694 B.n299 B.n298 10.6151
R695 B.n298 B.n295 10.6151
R696 B.n293 B.n290 10.6151
R697 B.n290 B.n289 10.6151
R698 B.n289 B.n286 10.6151
R699 B.n286 B.n285 10.6151
R700 B.n285 B.n282 10.6151
R701 B.n282 B.n281 10.6151
R702 B.n281 B.n278 10.6151
R703 B.n278 B.n277 10.6151
R704 B.n274 B.n273 10.6151
R705 B.n273 B.n270 10.6151
R706 B.n270 B.n269 10.6151
R707 B.n269 B.n266 10.6151
R708 B.n266 B.n265 10.6151
R709 B.n265 B.n262 10.6151
R710 B.n262 B.n261 10.6151
R711 B.n261 B.n258 10.6151
R712 B.n258 B.n257 10.6151
R713 B.n257 B.n254 10.6151
R714 B.n254 B.n253 10.6151
R715 B.n253 B.n250 10.6151
R716 B.n250 B.n249 10.6151
R717 B.n249 B.n246 10.6151
R718 B.n246 B.n245 10.6151
R719 B.n245 B.n242 10.6151
R720 B.n242 B.n241 10.6151
R721 B.n241 B.n238 10.6151
R722 B.n238 B.n237 10.6151
R723 B.n237 B.n203 10.6151
R724 B.n341 B.n203 10.6151
R725 B.n347 B.n199 10.6151
R726 B.n348 B.n347 10.6151
R727 B.n349 B.n348 10.6151
R728 B.n349 B.n191 10.6151
R729 B.n359 B.n191 10.6151
R730 B.n360 B.n359 10.6151
R731 B.n361 B.n360 10.6151
R732 B.n361 B.n183 10.6151
R733 B.n371 B.n183 10.6151
R734 B.n372 B.n371 10.6151
R735 B.n373 B.n372 10.6151
R736 B.n373 B.n175 10.6151
R737 B.n384 B.n175 10.6151
R738 B.n385 B.n384 10.6151
R739 B.n386 B.n385 10.6151
R740 B.n386 B.n0 10.6151
R741 B.n446 B.n1 10.6151
R742 B.n446 B.n445 10.6151
R743 B.n445 B.n444 10.6151
R744 B.n444 B.n10 10.6151
R745 B.n438 B.n10 10.6151
R746 B.n438 B.n437 10.6151
R747 B.n437 B.n436 10.6151
R748 B.n436 B.n17 10.6151
R749 B.n430 B.n17 10.6151
R750 B.n430 B.n429 10.6151
R751 B.n429 B.n428 10.6151
R752 B.n428 B.n24 10.6151
R753 B.n422 B.n24 10.6151
R754 B.n422 B.n421 10.6151
R755 B.n421 B.n420 10.6151
R756 B.n420 B.n31 10.6151
R757 B.n382 B.t0 8.40146
R758 B.n442 B.t1 8.40146
R759 B.n112 B.n66 6.5566
R760 B.n129 B.n128 6.5566
R761 B.n294 B.n293 6.5566
R762 B.n277 B.n235 6.5566
R763 B.n109 B.n66 4.05904
R764 B.n130 B.n129 4.05904
R765 B.n295 B.n294 4.05904
R766 B.n274 B.n235 4.05904
R767 B.n452 B.n0 2.81026
R768 B.n452 B.n1 2.81026
R769 VP.n0 VP.t0 251.369
R770 VP.n0 VP.t1 215.524
R771 VP VP.n0 0.146778
R772 VTAIL.n106 VTAIL.n84 289.615
R773 VTAIL.n22 VTAIL.n0 289.615
R774 VTAIL.n78 VTAIL.n56 289.615
R775 VTAIL.n50 VTAIL.n28 289.615
R776 VTAIL.n92 VTAIL.n91 185
R777 VTAIL.n97 VTAIL.n96 185
R778 VTAIL.n99 VTAIL.n98 185
R779 VTAIL.n88 VTAIL.n87 185
R780 VTAIL.n105 VTAIL.n104 185
R781 VTAIL.n107 VTAIL.n106 185
R782 VTAIL.n8 VTAIL.n7 185
R783 VTAIL.n13 VTAIL.n12 185
R784 VTAIL.n15 VTAIL.n14 185
R785 VTAIL.n4 VTAIL.n3 185
R786 VTAIL.n21 VTAIL.n20 185
R787 VTAIL.n23 VTAIL.n22 185
R788 VTAIL.n79 VTAIL.n78 185
R789 VTAIL.n77 VTAIL.n76 185
R790 VTAIL.n60 VTAIL.n59 185
R791 VTAIL.n71 VTAIL.n70 185
R792 VTAIL.n69 VTAIL.n68 185
R793 VTAIL.n64 VTAIL.n63 185
R794 VTAIL.n51 VTAIL.n50 185
R795 VTAIL.n49 VTAIL.n48 185
R796 VTAIL.n32 VTAIL.n31 185
R797 VTAIL.n43 VTAIL.n42 185
R798 VTAIL.n41 VTAIL.n40 185
R799 VTAIL.n36 VTAIL.n35 185
R800 VTAIL.n93 VTAIL.t1 147.672
R801 VTAIL.n9 VTAIL.t2 147.672
R802 VTAIL.n65 VTAIL.t3 147.672
R803 VTAIL.n37 VTAIL.t0 147.672
R804 VTAIL.n97 VTAIL.n91 104.615
R805 VTAIL.n98 VTAIL.n97 104.615
R806 VTAIL.n98 VTAIL.n87 104.615
R807 VTAIL.n105 VTAIL.n87 104.615
R808 VTAIL.n106 VTAIL.n105 104.615
R809 VTAIL.n13 VTAIL.n7 104.615
R810 VTAIL.n14 VTAIL.n13 104.615
R811 VTAIL.n14 VTAIL.n3 104.615
R812 VTAIL.n21 VTAIL.n3 104.615
R813 VTAIL.n22 VTAIL.n21 104.615
R814 VTAIL.n78 VTAIL.n77 104.615
R815 VTAIL.n77 VTAIL.n59 104.615
R816 VTAIL.n70 VTAIL.n59 104.615
R817 VTAIL.n70 VTAIL.n69 104.615
R818 VTAIL.n69 VTAIL.n63 104.615
R819 VTAIL.n50 VTAIL.n49 104.615
R820 VTAIL.n49 VTAIL.n31 104.615
R821 VTAIL.n42 VTAIL.n31 104.615
R822 VTAIL.n42 VTAIL.n41 104.615
R823 VTAIL.n41 VTAIL.n35 104.615
R824 VTAIL.t1 VTAIL.n91 52.3082
R825 VTAIL.t2 VTAIL.n7 52.3082
R826 VTAIL.t3 VTAIL.n63 52.3082
R827 VTAIL.t0 VTAIL.n35 52.3082
R828 VTAIL.n111 VTAIL.n110 30.6338
R829 VTAIL.n27 VTAIL.n26 30.6338
R830 VTAIL.n83 VTAIL.n82 30.6338
R831 VTAIL.n55 VTAIL.n54 30.6338
R832 VTAIL.n55 VTAIL.n27 19.5221
R833 VTAIL.n111 VTAIL.n83 18.1858
R834 VTAIL.n93 VTAIL.n92 15.6666
R835 VTAIL.n9 VTAIL.n8 15.6666
R836 VTAIL.n65 VTAIL.n64 15.6666
R837 VTAIL.n37 VTAIL.n36 15.6666
R838 VTAIL.n96 VTAIL.n95 12.8005
R839 VTAIL.n12 VTAIL.n11 12.8005
R840 VTAIL.n68 VTAIL.n67 12.8005
R841 VTAIL.n40 VTAIL.n39 12.8005
R842 VTAIL.n99 VTAIL.n90 12.0247
R843 VTAIL.n15 VTAIL.n6 12.0247
R844 VTAIL.n71 VTAIL.n62 12.0247
R845 VTAIL.n43 VTAIL.n34 12.0247
R846 VTAIL.n100 VTAIL.n88 11.249
R847 VTAIL.n16 VTAIL.n4 11.249
R848 VTAIL.n72 VTAIL.n60 11.249
R849 VTAIL.n44 VTAIL.n32 11.249
R850 VTAIL.n104 VTAIL.n103 10.4732
R851 VTAIL.n20 VTAIL.n19 10.4732
R852 VTAIL.n76 VTAIL.n75 10.4732
R853 VTAIL.n48 VTAIL.n47 10.4732
R854 VTAIL.n107 VTAIL.n86 9.69747
R855 VTAIL.n23 VTAIL.n2 9.69747
R856 VTAIL.n79 VTAIL.n58 9.69747
R857 VTAIL.n51 VTAIL.n30 9.69747
R858 VTAIL.n110 VTAIL.n109 9.45567
R859 VTAIL.n26 VTAIL.n25 9.45567
R860 VTAIL.n82 VTAIL.n81 9.45567
R861 VTAIL.n54 VTAIL.n53 9.45567
R862 VTAIL.n109 VTAIL.n108 9.3005
R863 VTAIL.n86 VTAIL.n85 9.3005
R864 VTAIL.n103 VTAIL.n102 9.3005
R865 VTAIL.n101 VTAIL.n100 9.3005
R866 VTAIL.n90 VTAIL.n89 9.3005
R867 VTAIL.n95 VTAIL.n94 9.3005
R868 VTAIL.n25 VTAIL.n24 9.3005
R869 VTAIL.n2 VTAIL.n1 9.3005
R870 VTAIL.n19 VTAIL.n18 9.3005
R871 VTAIL.n17 VTAIL.n16 9.3005
R872 VTAIL.n6 VTAIL.n5 9.3005
R873 VTAIL.n11 VTAIL.n10 9.3005
R874 VTAIL.n81 VTAIL.n80 9.3005
R875 VTAIL.n58 VTAIL.n57 9.3005
R876 VTAIL.n75 VTAIL.n74 9.3005
R877 VTAIL.n73 VTAIL.n72 9.3005
R878 VTAIL.n62 VTAIL.n61 9.3005
R879 VTAIL.n67 VTAIL.n66 9.3005
R880 VTAIL.n53 VTAIL.n52 9.3005
R881 VTAIL.n30 VTAIL.n29 9.3005
R882 VTAIL.n47 VTAIL.n46 9.3005
R883 VTAIL.n45 VTAIL.n44 9.3005
R884 VTAIL.n34 VTAIL.n33 9.3005
R885 VTAIL.n39 VTAIL.n38 9.3005
R886 VTAIL.n108 VTAIL.n84 8.92171
R887 VTAIL.n24 VTAIL.n0 8.92171
R888 VTAIL.n80 VTAIL.n56 8.92171
R889 VTAIL.n52 VTAIL.n28 8.92171
R890 VTAIL.n110 VTAIL.n84 5.04292
R891 VTAIL.n26 VTAIL.n0 5.04292
R892 VTAIL.n82 VTAIL.n56 5.04292
R893 VTAIL.n54 VTAIL.n28 5.04292
R894 VTAIL.n94 VTAIL.n93 4.38687
R895 VTAIL.n10 VTAIL.n9 4.38687
R896 VTAIL.n66 VTAIL.n65 4.38687
R897 VTAIL.n38 VTAIL.n37 4.38687
R898 VTAIL.n108 VTAIL.n107 4.26717
R899 VTAIL.n24 VTAIL.n23 4.26717
R900 VTAIL.n80 VTAIL.n79 4.26717
R901 VTAIL.n52 VTAIL.n51 4.26717
R902 VTAIL.n104 VTAIL.n86 3.49141
R903 VTAIL.n20 VTAIL.n2 3.49141
R904 VTAIL.n76 VTAIL.n58 3.49141
R905 VTAIL.n48 VTAIL.n30 3.49141
R906 VTAIL.n103 VTAIL.n88 2.71565
R907 VTAIL.n19 VTAIL.n4 2.71565
R908 VTAIL.n75 VTAIL.n60 2.71565
R909 VTAIL.n47 VTAIL.n32 2.71565
R910 VTAIL.n100 VTAIL.n99 1.93989
R911 VTAIL.n16 VTAIL.n15 1.93989
R912 VTAIL.n72 VTAIL.n71 1.93989
R913 VTAIL.n44 VTAIL.n43 1.93989
R914 VTAIL.n96 VTAIL.n90 1.16414
R915 VTAIL.n12 VTAIL.n6 1.16414
R916 VTAIL.n68 VTAIL.n62 1.16414
R917 VTAIL.n40 VTAIL.n34 1.16414
R918 VTAIL.n83 VTAIL.n55 1.13843
R919 VTAIL VTAIL.n27 0.862569
R920 VTAIL.n95 VTAIL.n92 0.388379
R921 VTAIL.n11 VTAIL.n8 0.388379
R922 VTAIL.n67 VTAIL.n64 0.388379
R923 VTAIL.n39 VTAIL.n36 0.388379
R924 VTAIL VTAIL.n111 0.276362
R925 VTAIL.n94 VTAIL.n89 0.155672
R926 VTAIL.n101 VTAIL.n89 0.155672
R927 VTAIL.n102 VTAIL.n101 0.155672
R928 VTAIL.n102 VTAIL.n85 0.155672
R929 VTAIL.n109 VTAIL.n85 0.155672
R930 VTAIL.n10 VTAIL.n5 0.155672
R931 VTAIL.n17 VTAIL.n5 0.155672
R932 VTAIL.n18 VTAIL.n17 0.155672
R933 VTAIL.n18 VTAIL.n1 0.155672
R934 VTAIL.n25 VTAIL.n1 0.155672
R935 VTAIL.n81 VTAIL.n57 0.155672
R936 VTAIL.n74 VTAIL.n57 0.155672
R937 VTAIL.n74 VTAIL.n73 0.155672
R938 VTAIL.n73 VTAIL.n61 0.155672
R939 VTAIL.n66 VTAIL.n61 0.155672
R940 VTAIL.n53 VTAIL.n29 0.155672
R941 VTAIL.n46 VTAIL.n29 0.155672
R942 VTAIL.n46 VTAIL.n45 0.155672
R943 VTAIL.n45 VTAIL.n33 0.155672
R944 VTAIL.n38 VTAIL.n33 0.155672
R945 VDD1.n22 VDD1.n0 289.615
R946 VDD1.n49 VDD1.n27 289.615
R947 VDD1.n23 VDD1.n22 185
R948 VDD1.n21 VDD1.n20 185
R949 VDD1.n4 VDD1.n3 185
R950 VDD1.n15 VDD1.n14 185
R951 VDD1.n13 VDD1.n12 185
R952 VDD1.n8 VDD1.n7 185
R953 VDD1.n35 VDD1.n34 185
R954 VDD1.n40 VDD1.n39 185
R955 VDD1.n42 VDD1.n41 185
R956 VDD1.n31 VDD1.n30 185
R957 VDD1.n48 VDD1.n47 185
R958 VDD1.n50 VDD1.n49 185
R959 VDD1.n9 VDD1.t1 147.672
R960 VDD1.n36 VDD1.t0 147.672
R961 VDD1.n22 VDD1.n21 104.615
R962 VDD1.n21 VDD1.n3 104.615
R963 VDD1.n14 VDD1.n3 104.615
R964 VDD1.n14 VDD1.n13 104.615
R965 VDD1.n13 VDD1.n7 104.615
R966 VDD1.n40 VDD1.n34 104.615
R967 VDD1.n41 VDD1.n40 104.615
R968 VDD1.n41 VDD1.n30 104.615
R969 VDD1.n48 VDD1.n30 104.615
R970 VDD1.n49 VDD1.n48 104.615
R971 VDD1 VDD1.n53 78.9861
R972 VDD1.t1 VDD1.n7 52.3082
R973 VDD1.t0 VDD1.n34 52.3082
R974 VDD1 VDD1.n26 47.7049
R975 VDD1.n9 VDD1.n8 15.6666
R976 VDD1.n36 VDD1.n35 15.6666
R977 VDD1.n12 VDD1.n11 12.8005
R978 VDD1.n39 VDD1.n38 12.8005
R979 VDD1.n15 VDD1.n6 12.0247
R980 VDD1.n42 VDD1.n33 12.0247
R981 VDD1.n16 VDD1.n4 11.249
R982 VDD1.n43 VDD1.n31 11.249
R983 VDD1.n20 VDD1.n19 10.4732
R984 VDD1.n47 VDD1.n46 10.4732
R985 VDD1.n23 VDD1.n2 9.69747
R986 VDD1.n50 VDD1.n29 9.69747
R987 VDD1.n26 VDD1.n25 9.45567
R988 VDD1.n53 VDD1.n52 9.45567
R989 VDD1.n25 VDD1.n24 9.3005
R990 VDD1.n2 VDD1.n1 9.3005
R991 VDD1.n19 VDD1.n18 9.3005
R992 VDD1.n17 VDD1.n16 9.3005
R993 VDD1.n6 VDD1.n5 9.3005
R994 VDD1.n11 VDD1.n10 9.3005
R995 VDD1.n52 VDD1.n51 9.3005
R996 VDD1.n29 VDD1.n28 9.3005
R997 VDD1.n46 VDD1.n45 9.3005
R998 VDD1.n44 VDD1.n43 9.3005
R999 VDD1.n33 VDD1.n32 9.3005
R1000 VDD1.n38 VDD1.n37 9.3005
R1001 VDD1.n24 VDD1.n0 8.92171
R1002 VDD1.n51 VDD1.n27 8.92171
R1003 VDD1.n26 VDD1.n0 5.04292
R1004 VDD1.n53 VDD1.n27 5.04292
R1005 VDD1.n10 VDD1.n9 4.38687
R1006 VDD1.n37 VDD1.n36 4.38687
R1007 VDD1.n24 VDD1.n23 4.26717
R1008 VDD1.n51 VDD1.n50 4.26717
R1009 VDD1.n20 VDD1.n2 3.49141
R1010 VDD1.n47 VDD1.n29 3.49141
R1011 VDD1.n19 VDD1.n4 2.71565
R1012 VDD1.n46 VDD1.n31 2.71565
R1013 VDD1.n16 VDD1.n15 1.93989
R1014 VDD1.n43 VDD1.n42 1.93989
R1015 VDD1.n12 VDD1.n6 1.16414
R1016 VDD1.n39 VDD1.n33 1.16414
R1017 VDD1.n11 VDD1.n8 0.388379
R1018 VDD1.n38 VDD1.n35 0.388379
R1019 VDD1.n25 VDD1.n1 0.155672
R1020 VDD1.n18 VDD1.n1 0.155672
R1021 VDD1.n18 VDD1.n17 0.155672
R1022 VDD1.n17 VDD1.n5 0.155672
R1023 VDD1.n10 VDD1.n5 0.155672
R1024 VDD1.n37 VDD1.n32 0.155672
R1025 VDD1.n44 VDD1.n32 0.155672
R1026 VDD1.n45 VDD1.n44 0.155672
R1027 VDD1.n45 VDD1.n28 0.155672
R1028 VDD1.n52 VDD1.n28 0.155672
R1029 VN VN.t1 251.655
R1030 VN VN.t0 215.671
R1031 VDD2.n49 VDD2.n27 289.615
R1032 VDD2.n22 VDD2.n0 289.615
R1033 VDD2.n50 VDD2.n49 185
R1034 VDD2.n48 VDD2.n47 185
R1035 VDD2.n31 VDD2.n30 185
R1036 VDD2.n42 VDD2.n41 185
R1037 VDD2.n40 VDD2.n39 185
R1038 VDD2.n35 VDD2.n34 185
R1039 VDD2.n8 VDD2.n7 185
R1040 VDD2.n13 VDD2.n12 185
R1041 VDD2.n15 VDD2.n14 185
R1042 VDD2.n4 VDD2.n3 185
R1043 VDD2.n21 VDD2.n20 185
R1044 VDD2.n23 VDD2.n22 185
R1045 VDD2.n36 VDD2.t0 147.672
R1046 VDD2.n9 VDD2.t1 147.672
R1047 VDD2.n49 VDD2.n48 104.615
R1048 VDD2.n48 VDD2.n30 104.615
R1049 VDD2.n41 VDD2.n30 104.615
R1050 VDD2.n41 VDD2.n40 104.615
R1051 VDD2.n40 VDD2.n34 104.615
R1052 VDD2.n13 VDD2.n7 104.615
R1053 VDD2.n14 VDD2.n13 104.615
R1054 VDD2.n14 VDD2.n3 104.615
R1055 VDD2.n21 VDD2.n3 104.615
R1056 VDD2.n22 VDD2.n21 104.615
R1057 VDD2.n54 VDD2.n26 78.1272
R1058 VDD2.t0 VDD2.n34 52.3082
R1059 VDD2.t1 VDD2.n7 52.3082
R1060 VDD2.n54 VDD2.n53 47.3126
R1061 VDD2.n36 VDD2.n35 15.6666
R1062 VDD2.n9 VDD2.n8 15.6666
R1063 VDD2.n39 VDD2.n38 12.8005
R1064 VDD2.n12 VDD2.n11 12.8005
R1065 VDD2.n42 VDD2.n33 12.0247
R1066 VDD2.n15 VDD2.n6 12.0247
R1067 VDD2.n43 VDD2.n31 11.249
R1068 VDD2.n16 VDD2.n4 11.249
R1069 VDD2.n47 VDD2.n46 10.4732
R1070 VDD2.n20 VDD2.n19 10.4732
R1071 VDD2.n50 VDD2.n29 9.69747
R1072 VDD2.n23 VDD2.n2 9.69747
R1073 VDD2.n53 VDD2.n52 9.45567
R1074 VDD2.n26 VDD2.n25 9.45567
R1075 VDD2.n52 VDD2.n51 9.3005
R1076 VDD2.n29 VDD2.n28 9.3005
R1077 VDD2.n46 VDD2.n45 9.3005
R1078 VDD2.n44 VDD2.n43 9.3005
R1079 VDD2.n33 VDD2.n32 9.3005
R1080 VDD2.n38 VDD2.n37 9.3005
R1081 VDD2.n25 VDD2.n24 9.3005
R1082 VDD2.n2 VDD2.n1 9.3005
R1083 VDD2.n19 VDD2.n18 9.3005
R1084 VDD2.n17 VDD2.n16 9.3005
R1085 VDD2.n6 VDD2.n5 9.3005
R1086 VDD2.n11 VDD2.n10 9.3005
R1087 VDD2.n51 VDD2.n27 8.92171
R1088 VDD2.n24 VDD2.n0 8.92171
R1089 VDD2.n53 VDD2.n27 5.04292
R1090 VDD2.n26 VDD2.n0 5.04292
R1091 VDD2.n37 VDD2.n36 4.38687
R1092 VDD2.n10 VDD2.n9 4.38687
R1093 VDD2.n51 VDD2.n50 4.26717
R1094 VDD2.n24 VDD2.n23 4.26717
R1095 VDD2.n47 VDD2.n29 3.49141
R1096 VDD2.n20 VDD2.n2 3.49141
R1097 VDD2.n46 VDD2.n31 2.71565
R1098 VDD2.n19 VDD2.n4 2.71565
R1099 VDD2.n43 VDD2.n42 1.93989
R1100 VDD2.n16 VDD2.n15 1.93989
R1101 VDD2.n39 VDD2.n33 1.16414
R1102 VDD2.n12 VDD2.n6 1.16414
R1103 VDD2 VDD2.n54 0.392741
R1104 VDD2.n38 VDD2.n35 0.388379
R1105 VDD2.n11 VDD2.n8 0.388379
R1106 VDD2.n52 VDD2.n28 0.155672
R1107 VDD2.n45 VDD2.n28 0.155672
R1108 VDD2.n45 VDD2.n44 0.155672
R1109 VDD2.n44 VDD2.n32 0.155672
R1110 VDD2.n37 VDD2.n32 0.155672
R1111 VDD2.n10 VDD2.n5 0.155672
R1112 VDD2.n17 VDD2.n5 0.155672
R1113 VDD2.n18 VDD2.n17 0.155672
R1114 VDD2.n18 VDD2.n1 0.155672
R1115 VDD2.n25 VDD2.n1 0.155672
C0 VDD1 VTAIL 3.03416f
C1 VN VP 3.54835f
C2 VDD2 VP 0.27873f
C3 VTAIL VP 1.09548f
C4 VDD1 VP 1.29064f
C5 VN VDD2 1.16541f
C6 VN VTAIL 1.08122f
C7 VDD2 VTAIL 3.07604f
C8 VN VDD1 0.147823f
C9 VDD1 VDD2 0.513985f
C10 VDD2 B 2.691209f
C11 VDD1 B 4.05843f
C12 VTAIL B 3.854955f
C13 VN B 6.29709f
C14 VP B 4.132893f
C15 VDD2.n0 B 0.020205f
C16 VDD2.n1 B 0.015253f
C17 VDD2.n2 B 0.008196f
C18 VDD2.n3 B 0.019374f
C19 VDD2.n4 B 0.008679f
C20 VDD2.n5 B 0.015253f
C21 VDD2.n6 B 0.008196f
C22 VDD2.n7 B 0.01453f
C23 VDD2.n8 B 0.011441f
C24 VDD2.t1 B 0.031591f
C25 VDD2.n9 B 0.062316f
C26 VDD2.n10 B 0.306856f
C27 VDD2.n11 B 0.008196f
C28 VDD2.n12 B 0.008679f
C29 VDD2.n13 B 0.019374f
C30 VDD2.n14 B 0.019374f
C31 VDD2.n15 B 0.008679f
C32 VDD2.n16 B 0.008196f
C33 VDD2.n17 B 0.015253f
C34 VDD2.n18 B 0.015253f
C35 VDD2.n19 B 0.008196f
C36 VDD2.n20 B 0.008679f
C37 VDD2.n21 B 0.019374f
C38 VDD2.n22 B 0.039756f
C39 VDD2.n23 B 0.008679f
C40 VDD2.n24 B 0.008196f
C41 VDD2.n25 B 0.03359f
C42 VDD2.n26 B 0.266959f
C43 VDD2.n27 B 0.020205f
C44 VDD2.n28 B 0.015253f
C45 VDD2.n29 B 0.008196f
C46 VDD2.n30 B 0.019374f
C47 VDD2.n31 B 0.008679f
C48 VDD2.n32 B 0.015253f
C49 VDD2.n33 B 0.008196f
C50 VDD2.n34 B 0.01453f
C51 VDD2.n35 B 0.011441f
C52 VDD2.t0 B 0.031591f
C53 VDD2.n36 B 0.062316f
C54 VDD2.n37 B 0.306856f
C55 VDD2.n38 B 0.008196f
C56 VDD2.n39 B 0.008679f
C57 VDD2.n40 B 0.019374f
C58 VDD2.n41 B 0.019374f
C59 VDD2.n42 B 0.008679f
C60 VDD2.n43 B 0.008196f
C61 VDD2.n44 B 0.015253f
C62 VDD2.n45 B 0.015253f
C63 VDD2.n46 B 0.008196f
C64 VDD2.n47 B 0.008679f
C65 VDD2.n48 B 0.019374f
C66 VDD2.n49 B 0.039756f
C67 VDD2.n50 B 0.008679f
C68 VDD2.n51 B 0.008196f
C69 VDD2.n52 B 0.03359f
C70 VDD2.n53 B 0.032515f
C71 VDD2.n54 B 1.24525f
C72 VN.t0 B 0.63013f
C73 VN.t1 B 0.788185f
C74 VDD1.n0 B 0.019204f
C75 VDD1.n1 B 0.014498f
C76 VDD1.n2 B 0.00779f
C77 VDD1.n3 B 0.018414f
C78 VDD1.n4 B 0.008249f
C79 VDD1.n5 B 0.014498f
C80 VDD1.n6 B 0.00779f
C81 VDD1.n7 B 0.01381f
C82 VDD1.n8 B 0.010875f
C83 VDD1.t1 B 0.030027f
C84 VDD1.n9 B 0.05923f
C85 VDD1.n10 B 0.291657f
C86 VDD1.n11 B 0.00779f
C87 VDD1.n12 B 0.008249f
C88 VDD1.n13 B 0.018414f
C89 VDD1.n14 B 0.018414f
C90 VDD1.n15 B 0.008249f
C91 VDD1.n16 B 0.00779f
C92 VDD1.n17 B 0.014498f
C93 VDD1.n18 B 0.014498f
C94 VDD1.n19 B 0.00779f
C95 VDD1.n20 B 0.008249f
C96 VDD1.n21 B 0.018414f
C97 VDD1.n22 B 0.037787f
C98 VDD1.n23 B 0.008249f
C99 VDD1.n24 B 0.00779f
C100 VDD1.n25 B 0.031927f
C101 VDD1.n26 B 0.031277f
C102 VDD1.n27 B 0.019204f
C103 VDD1.n28 B 0.014498f
C104 VDD1.n29 B 0.00779f
C105 VDD1.n30 B 0.018414f
C106 VDD1.n31 B 0.008249f
C107 VDD1.n32 B 0.014498f
C108 VDD1.n33 B 0.00779f
C109 VDD1.n34 B 0.01381f
C110 VDD1.n35 B 0.010875f
C111 VDD1.t0 B 0.030027f
C112 VDD1.n36 B 0.05923f
C113 VDD1.n37 B 0.291657f
C114 VDD1.n38 B 0.00779f
C115 VDD1.n39 B 0.008249f
C116 VDD1.n40 B 0.018414f
C117 VDD1.n41 B 0.018414f
C118 VDD1.n42 B 0.008249f
C119 VDD1.n43 B 0.00779f
C120 VDD1.n44 B 0.014498f
C121 VDD1.n45 B 0.014498f
C122 VDD1.n46 B 0.00779f
C123 VDD1.n47 B 0.008249f
C124 VDD1.n48 B 0.018414f
C125 VDD1.n49 B 0.037787f
C126 VDD1.n50 B 0.008249f
C127 VDD1.n51 B 0.00779f
C128 VDD1.n52 B 0.031927f
C129 VDD1.n53 B 0.272881f
C130 VTAIL.n0 B 0.022534f
C131 VTAIL.n1 B 0.017011f
C132 VTAIL.n2 B 0.009141f
C133 VTAIL.n3 B 0.021607f
C134 VTAIL.n4 B 0.009679f
C135 VTAIL.n5 B 0.017011f
C136 VTAIL.n6 B 0.009141f
C137 VTAIL.n7 B 0.016205f
C138 VTAIL.n8 B 0.01276f
C139 VTAIL.t2 B 0.035233f
C140 VTAIL.n9 B 0.069499f
C141 VTAIL.n10 B 0.342226f
C142 VTAIL.n11 B 0.009141f
C143 VTAIL.n12 B 0.009679f
C144 VTAIL.n13 B 0.021607f
C145 VTAIL.n14 B 0.021607f
C146 VTAIL.n15 B 0.009679f
C147 VTAIL.n16 B 0.009141f
C148 VTAIL.n17 B 0.017011f
C149 VTAIL.n18 B 0.017011f
C150 VTAIL.n19 B 0.009141f
C151 VTAIL.n20 B 0.009679f
C152 VTAIL.n21 B 0.021607f
C153 VTAIL.n22 B 0.044339f
C154 VTAIL.n23 B 0.009679f
C155 VTAIL.n24 B 0.009141f
C156 VTAIL.n25 B 0.037462f
C157 VTAIL.n26 B 0.024501f
C158 VTAIL.n27 B 0.684027f
C159 VTAIL.n28 B 0.022534f
C160 VTAIL.n29 B 0.017011f
C161 VTAIL.n30 B 0.009141f
C162 VTAIL.n31 B 0.021607f
C163 VTAIL.n32 B 0.009679f
C164 VTAIL.n33 B 0.017011f
C165 VTAIL.n34 B 0.009141f
C166 VTAIL.n35 B 0.016205f
C167 VTAIL.n36 B 0.01276f
C168 VTAIL.t0 B 0.035233f
C169 VTAIL.n37 B 0.069499f
C170 VTAIL.n38 B 0.342226f
C171 VTAIL.n39 B 0.009141f
C172 VTAIL.n40 B 0.009679f
C173 VTAIL.n41 B 0.021607f
C174 VTAIL.n42 B 0.021607f
C175 VTAIL.n43 B 0.009679f
C176 VTAIL.n44 B 0.009141f
C177 VTAIL.n45 B 0.017011f
C178 VTAIL.n46 B 0.017011f
C179 VTAIL.n47 B 0.009141f
C180 VTAIL.n48 B 0.009679f
C181 VTAIL.n49 B 0.021607f
C182 VTAIL.n50 B 0.044339f
C183 VTAIL.n51 B 0.009679f
C184 VTAIL.n52 B 0.009141f
C185 VTAIL.n53 B 0.037462f
C186 VTAIL.n54 B 0.024501f
C187 VTAIL.n55 B 0.699148f
C188 VTAIL.n56 B 0.022534f
C189 VTAIL.n57 B 0.017011f
C190 VTAIL.n58 B 0.009141f
C191 VTAIL.n59 B 0.021607f
C192 VTAIL.n60 B 0.009679f
C193 VTAIL.n61 B 0.017011f
C194 VTAIL.n62 B 0.009141f
C195 VTAIL.n63 B 0.016205f
C196 VTAIL.n64 B 0.01276f
C197 VTAIL.t3 B 0.035233f
C198 VTAIL.n65 B 0.069499f
C199 VTAIL.n66 B 0.342226f
C200 VTAIL.n67 B 0.009141f
C201 VTAIL.n68 B 0.009679f
C202 VTAIL.n69 B 0.021607f
C203 VTAIL.n70 B 0.021607f
C204 VTAIL.n71 B 0.009679f
C205 VTAIL.n72 B 0.009141f
C206 VTAIL.n73 B 0.017011f
C207 VTAIL.n74 B 0.017011f
C208 VTAIL.n75 B 0.009141f
C209 VTAIL.n76 B 0.009679f
C210 VTAIL.n77 B 0.021607f
C211 VTAIL.n78 B 0.044339f
C212 VTAIL.n79 B 0.009679f
C213 VTAIL.n80 B 0.009141f
C214 VTAIL.n81 B 0.037462f
C215 VTAIL.n82 B 0.024501f
C216 VTAIL.n83 B 0.625904f
C217 VTAIL.n84 B 0.022534f
C218 VTAIL.n85 B 0.017011f
C219 VTAIL.n86 B 0.009141f
C220 VTAIL.n87 B 0.021607f
C221 VTAIL.n88 B 0.009679f
C222 VTAIL.n89 B 0.017011f
C223 VTAIL.n90 B 0.009141f
C224 VTAIL.n91 B 0.016205f
C225 VTAIL.n92 B 0.01276f
C226 VTAIL.t1 B 0.035233f
C227 VTAIL.n93 B 0.069499f
C228 VTAIL.n94 B 0.342226f
C229 VTAIL.n95 B 0.009141f
C230 VTAIL.n96 B 0.009679f
C231 VTAIL.n97 B 0.021607f
C232 VTAIL.n98 B 0.021607f
C233 VTAIL.n99 B 0.009679f
C234 VTAIL.n100 B 0.009141f
C235 VTAIL.n101 B 0.017011f
C236 VTAIL.n102 B 0.017011f
C237 VTAIL.n103 B 0.009141f
C238 VTAIL.n104 B 0.009679f
C239 VTAIL.n105 B 0.021607f
C240 VTAIL.n106 B 0.044339f
C241 VTAIL.n107 B 0.009679f
C242 VTAIL.n108 B 0.009141f
C243 VTAIL.n109 B 0.037462f
C244 VTAIL.n110 B 0.024501f
C245 VTAIL.n111 B 0.57865f
C246 VP.t0 B 0.793976f
C247 VP.t1 B 0.637427f
C248 VP.n0 B 2.0432f
.ends

