* NGSPICE file created from diff_pair_sample_1212.ext - technology: sky130A

.subckt diff_pair_sample_1212 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 w_n1782_n3040# sky130_fd_pr__pfet_01v8 ad=4.0404 pd=21.5 as=4.0404 ps=21.5 w=10.36 l=1.7
X1 VDD2.t1 VN.t0 VTAIL.t0 w_n1782_n3040# sky130_fd_pr__pfet_01v8 ad=4.0404 pd=21.5 as=4.0404 ps=21.5 w=10.36 l=1.7
X2 B.t11 B.t9 B.t10 w_n1782_n3040# sky130_fd_pr__pfet_01v8 ad=4.0404 pd=21.5 as=0 ps=0 w=10.36 l=1.7
X3 VDD1.t0 VP.t1 VTAIL.t1 w_n1782_n3040# sky130_fd_pr__pfet_01v8 ad=4.0404 pd=21.5 as=4.0404 ps=21.5 w=10.36 l=1.7
X4 VDD2.t0 VN.t1 VTAIL.t3 w_n1782_n3040# sky130_fd_pr__pfet_01v8 ad=4.0404 pd=21.5 as=4.0404 ps=21.5 w=10.36 l=1.7
X5 B.t8 B.t6 B.t7 w_n1782_n3040# sky130_fd_pr__pfet_01v8 ad=4.0404 pd=21.5 as=0 ps=0 w=10.36 l=1.7
X6 B.t5 B.t3 B.t4 w_n1782_n3040# sky130_fd_pr__pfet_01v8 ad=4.0404 pd=21.5 as=0 ps=0 w=10.36 l=1.7
X7 B.t2 B.t0 B.t1 w_n1782_n3040# sky130_fd_pr__pfet_01v8 ad=4.0404 pd=21.5 as=0 ps=0 w=10.36 l=1.7
R0 VP.n0 VP.t1 246.781
R1 VP.n0 VP.t0 205.755
R2 VP VP.n0 0.241678
R3 VTAIL.n1 VTAIL.t3 63.7032
R4 VTAIL.n2 VTAIL.t1 63.703
R5 VTAIL.n3 VTAIL.t0 63.703
R6 VTAIL.n0 VTAIL.t2 63.703
R7 VTAIL.n1 VTAIL.n0 24.7979
R8 VTAIL.n3 VTAIL.n2 23.0479
R9 VTAIL.n2 VTAIL.n1 1.34533
R10 VTAIL VTAIL.n0 0.966017
R11 VTAIL VTAIL.n3 0.37981
R12 VDD1 VDD1.t1 117.434
R13 VDD1 VDD1.t0 80.8775
R14 VN VN.t1 246.974
R15 VN VN.t0 205.995
R16 VDD2.n0 VDD2.t1 116.472
R17 VDD2.n0 VDD2.t0 80.3818
R18 VDD2 VDD2.n0 0.49619
R19 B.n351 B.n58 585
R20 B.n353 B.n352 585
R21 B.n354 B.n57 585
R22 B.n356 B.n355 585
R23 B.n357 B.n56 585
R24 B.n359 B.n358 585
R25 B.n360 B.n55 585
R26 B.n362 B.n361 585
R27 B.n363 B.n54 585
R28 B.n365 B.n364 585
R29 B.n366 B.n53 585
R30 B.n368 B.n367 585
R31 B.n369 B.n52 585
R32 B.n371 B.n370 585
R33 B.n372 B.n51 585
R34 B.n374 B.n373 585
R35 B.n375 B.n50 585
R36 B.n377 B.n376 585
R37 B.n378 B.n49 585
R38 B.n380 B.n379 585
R39 B.n381 B.n48 585
R40 B.n383 B.n382 585
R41 B.n384 B.n47 585
R42 B.n386 B.n385 585
R43 B.n387 B.n46 585
R44 B.n389 B.n388 585
R45 B.n390 B.n45 585
R46 B.n392 B.n391 585
R47 B.n393 B.n44 585
R48 B.n395 B.n394 585
R49 B.n396 B.n43 585
R50 B.n398 B.n397 585
R51 B.n399 B.n42 585
R52 B.n401 B.n400 585
R53 B.n402 B.n41 585
R54 B.n404 B.n403 585
R55 B.n405 B.n38 585
R56 B.n408 B.n407 585
R57 B.n409 B.n37 585
R58 B.n411 B.n410 585
R59 B.n412 B.n36 585
R60 B.n414 B.n413 585
R61 B.n415 B.n35 585
R62 B.n417 B.n416 585
R63 B.n418 B.n31 585
R64 B.n420 B.n419 585
R65 B.n421 B.n30 585
R66 B.n423 B.n422 585
R67 B.n424 B.n29 585
R68 B.n426 B.n425 585
R69 B.n427 B.n28 585
R70 B.n429 B.n428 585
R71 B.n430 B.n27 585
R72 B.n432 B.n431 585
R73 B.n433 B.n26 585
R74 B.n435 B.n434 585
R75 B.n436 B.n25 585
R76 B.n438 B.n437 585
R77 B.n439 B.n24 585
R78 B.n441 B.n440 585
R79 B.n442 B.n23 585
R80 B.n444 B.n443 585
R81 B.n445 B.n22 585
R82 B.n447 B.n446 585
R83 B.n448 B.n21 585
R84 B.n450 B.n449 585
R85 B.n451 B.n20 585
R86 B.n453 B.n452 585
R87 B.n454 B.n19 585
R88 B.n456 B.n455 585
R89 B.n457 B.n18 585
R90 B.n459 B.n458 585
R91 B.n460 B.n17 585
R92 B.n462 B.n461 585
R93 B.n463 B.n16 585
R94 B.n465 B.n464 585
R95 B.n466 B.n15 585
R96 B.n468 B.n467 585
R97 B.n469 B.n14 585
R98 B.n471 B.n470 585
R99 B.n472 B.n13 585
R100 B.n474 B.n473 585
R101 B.n475 B.n12 585
R102 B.n350 B.n349 585
R103 B.n348 B.n59 585
R104 B.n347 B.n346 585
R105 B.n345 B.n60 585
R106 B.n344 B.n343 585
R107 B.n342 B.n61 585
R108 B.n341 B.n340 585
R109 B.n339 B.n62 585
R110 B.n338 B.n337 585
R111 B.n336 B.n63 585
R112 B.n335 B.n334 585
R113 B.n333 B.n64 585
R114 B.n332 B.n331 585
R115 B.n330 B.n65 585
R116 B.n329 B.n328 585
R117 B.n327 B.n66 585
R118 B.n326 B.n325 585
R119 B.n324 B.n67 585
R120 B.n323 B.n322 585
R121 B.n321 B.n68 585
R122 B.n320 B.n319 585
R123 B.n318 B.n69 585
R124 B.n317 B.n316 585
R125 B.n315 B.n70 585
R126 B.n314 B.n313 585
R127 B.n312 B.n71 585
R128 B.n311 B.n310 585
R129 B.n309 B.n72 585
R130 B.n308 B.n307 585
R131 B.n306 B.n73 585
R132 B.n305 B.n304 585
R133 B.n303 B.n74 585
R134 B.n302 B.n301 585
R135 B.n300 B.n75 585
R136 B.n299 B.n298 585
R137 B.n297 B.n76 585
R138 B.n296 B.n295 585
R139 B.n294 B.n77 585
R140 B.n293 B.n292 585
R141 B.n291 B.n78 585
R142 B.n290 B.n289 585
R143 B.n161 B.n122 585
R144 B.n163 B.n162 585
R145 B.n164 B.n121 585
R146 B.n166 B.n165 585
R147 B.n167 B.n120 585
R148 B.n169 B.n168 585
R149 B.n170 B.n119 585
R150 B.n172 B.n171 585
R151 B.n173 B.n118 585
R152 B.n175 B.n174 585
R153 B.n176 B.n117 585
R154 B.n178 B.n177 585
R155 B.n179 B.n116 585
R156 B.n181 B.n180 585
R157 B.n182 B.n115 585
R158 B.n184 B.n183 585
R159 B.n185 B.n114 585
R160 B.n187 B.n186 585
R161 B.n188 B.n113 585
R162 B.n190 B.n189 585
R163 B.n191 B.n112 585
R164 B.n193 B.n192 585
R165 B.n194 B.n111 585
R166 B.n196 B.n195 585
R167 B.n197 B.n110 585
R168 B.n199 B.n198 585
R169 B.n200 B.n109 585
R170 B.n202 B.n201 585
R171 B.n203 B.n108 585
R172 B.n205 B.n204 585
R173 B.n206 B.n107 585
R174 B.n208 B.n207 585
R175 B.n209 B.n106 585
R176 B.n211 B.n210 585
R177 B.n212 B.n105 585
R178 B.n214 B.n213 585
R179 B.n215 B.n102 585
R180 B.n218 B.n217 585
R181 B.n219 B.n101 585
R182 B.n221 B.n220 585
R183 B.n222 B.n100 585
R184 B.n224 B.n223 585
R185 B.n225 B.n99 585
R186 B.n227 B.n226 585
R187 B.n228 B.n98 585
R188 B.n233 B.n232 585
R189 B.n234 B.n97 585
R190 B.n236 B.n235 585
R191 B.n237 B.n96 585
R192 B.n239 B.n238 585
R193 B.n240 B.n95 585
R194 B.n242 B.n241 585
R195 B.n243 B.n94 585
R196 B.n245 B.n244 585
R197 B.n246 B.n93 585
R198 B.n248 B.n247 585
R199 B.n249 B.n92 585
R200 B.n251 B.n250 585
R201 B.n252 B.n91 585
R202 B.n254 B.n253 585
R203 B.n255 B.n90 585
R204 B.n257 B.n256 585
R205 B.n258 B.n89 585
R206 B.n260 B.n259 585
R207 B.n261 B.n88 585
R208 B.n263 B.n262 585
R209 B.n264 B.n87 585
R210 B.n266 B.n265 585
R211 B.n267 B.n86 585
R212 B.n269 B.n268 585
R213 B.n270 B.n85 585
R214 B.n272 B.n271 585
R215 B.n273 B.n84 585
R216 B.n275 B.n274 585
R217 B.n276 B.n83 585
R218 B.n278 B.n277 585
R219 B.n279 B.n82 585
R220 B.n281 B.n280 585
R221 B.n282 B.n81 585
R222 B.n284 B.n283 585
R223 B.n285 B.n80 585
R224 B.n287 B.n286 585
R225 B.n288 B.n79 585
R226 B.n160 B.n159 585
R227 B.n158 B.n123 585
R228 B.n157 B.n156 585
R229 B.n155 B.n124 585
R230 B.n154 B.n153 585
R231 B.n152 B.n125 585
R232 B.n151 B.n150 585
R233 B.n149 B.n126 585
R234 B.n148 B.n147 585
R235 B.n146 B.n127 585
R236 B.n145 B.n144 585
R237 B.n143 B.n128 585
R238 B.n142 B.n141 585
R239 B.n140 B.n129 585
R240 B.n139 B.n138 585
R241 B.n137 B.n130 585
R242 B.n136 B.n135 585
R243 B.n134 B.n131 585
R244 B.n133 B.n132 585
R245 B.n2 B.n0 585
R246 B.n505 B.n1 585
R247 B.n504 B.n503 585
R248 B.n502 B.n3 585
R249 B.n501 B.n500 585
R250 B.n499 B.n4 585
R251 B.n498 B.n497 585
R252 B.n496 B.n5 585
R253 B.n495 B.n494 585
R254 B.n493 B.n6 585
R255 B.n492 B.n491 585
R256 B.n490 B.n7 585
R257 B.n489 B.n488 585
R258 B.n487 B.n8 585
R259 B.n486 B.n485 585
R260 B.n484 B.n9 585
R261 B.n483 B.n482 585
R262 B.n481 B.n10 585
R263 B.n480 B.n479 585
R264 B.n478 B.n11 585
R265 B.n477 B.n476 585
R266 B.n507 B.n506 585
R267 B.n159 B.n122 521.33
R268 B.n476 B.n475 521.33
R269 B.n289 B.n288 521.33
R270 B.n349 B.n58 521.33
R271 B.n229 B.t0 352.983
R272 B.n103 B.t6 352.983
R273 B.n32 B.t3 352.983
R274 B.n39 B.t9 352.983
R275 B.n159 B.n158 163.367
R276 B.n158 B.n157 163.367
R277 B.n157 B.n124 163.367
R278 B.n153 B.n124 163.367
R279 B.n153 B.n152 163.367
R280 B.n152 B.n151 163.367
R281 B.n151 B.n126 163.367
R282 B.n147 B.n126 163.367
R283 B.n147 B.n146 163.367
R284 B.n146 B.n145 163.367
R285 B.n145 B.n128 163.367
R286 B.n141 B.n128 163.367
R287 B.n141 B.n140 163.367
R288 B.n140 B.n139 163.367
R289 B.n139 B.n130 163.367
R290 B.n135 B.n130 163.367
R291 B.n135 B.n134 163.367
R292 B.n134 B.n133 163.367
R293 B.n133 B.n2 163.367
R294 B.n506 B.n2 163.367
R295 B.n506 B.n505 163.367
R296 B.n505 B.n504 163.367
R297 B.n504 B.n3 163.367
R298 B.n500 B.n3 163.367
R299 B.n500 B.n499 163.367
R300 B.n499 B.n498 163.367
R301 B.n498 B.n5 163.367
R302 B.n494 B.n5 163.367
R303 B.n494 B.n493 163.367
R304 B.n493 B.n492 163.367
R305 B.n492 B.n7 163.367
R306 B.n488 B.n7 163.367
R307 B.n488 B.n487 163.367
R308 B.n487 B.n486 163.367
R309 B.n486 B.n9 163.367
R310 B.n482 B.n9 163.367
R311 B.n482 B.n481 163.367
R312 B.n481 B.n480 163.367
R313 B.n480 B.n11 163.367
R314 B.n476 B.n11 163.367
R315 B.n163 B.n122 163.367
R316 B.n164 B.n163 163.367
R317 B.n165 B.n164 163.367
R318 B.n165 B.n120 163.367
R319 B.n169 B.n120 163.367
R320 B.n170 B.n169 163.367
R321 B.n171 B.n170 163.367
R322 B.n171 B.n118 163.367
R323 B.n175 B.n118 163.367
R324 B.n176 B.n175 163.367
R325 B.n177 B.n176 163.367
R326 B.n177 B.n116 163.367
R327 B.n181 B.n116 163.367
R328 B.n182 B.n181 163.367
R329 B.n183 B.n182 163.367
R330 B.n183 B.n114 163.367
R331 B.n187 B.n114 163.367
R332 B.n188 B.n187 163.367
R333 B.n189 B.n188 163.367
R334 B.n189 B.n112 163.367
R335 B.n193 B.n112 163.367
R336 B.n194 B.n193 163.367
R337 B.n195 B.n194 163.367
R338 B.n195 B.n110 163.367
R339 B.n199 B.n110 163.367
R340 B.n200 B.n199 163.367
R341 B.n201 B.n200 163.367
R342 B.n201 B.n108 163.367
R343 B.n205 B.n108 163.367
R344 B.n206 B.n205 163.367
R345 B.n207 B.n206 163.367
R346 B.n207 B.n106 163.367
R347 B.n211 B.n106 163.367
R348 B.n212 B.n211 163.367
R349 B.n213 B.n212 163.367
R350 B.n213 B.n102 163.367
R351 B.n218 B.n102 163.367
R352 B.n219 B.n218 163.367
R353 B.n220 B.n219 163.367
R354 B.n220 B.n100 163.367
R355 B.n224 B.n100 163.367
R356 B.n225 B.n224 163.367
R357 B.n226 B.n225 163.367
R358 B.n226 B.n98 163.367
R359 B.n233 B.n98 163.367
R360 B.n234 B.n233 163.367
R361 B.n235 B.n234 163.367
R362 B.n235 B.n96 163.367
R363 B.n239 B.n96 163.367
R364 B.n240 B.n239 163.367
R365 B.n241 B.n240 163.367
R366 B.n241 B.n94 163.367
R367 B.n245 B.n94 163.367
R368 B.n246 B.n245 163.367
R369 B.n247 B.n246 163.367
R370 B.n247 B.n92 163.367
R371 B.n251 B.n92 163.367
R372 B.n252 B.n251 163.367
R373 B.n253 B.n252 163.367
R374 B.n253 B.n90 163.367
R375 B.n257 B.n90 163.367
R376 B.n258 B.n257 163.367
R377 B.n259 B.n258 163.367
R378 B.n259 B.n88 163.367
R379 B.n263 B.n88 163.367
R380 B.n264 B.n263 163.367
R381 B.n265 B.n264 163.367
R382 B.n265 B.n86 163.367
R383 B.n269 B.n86 163.367
R384 B.n270 B.n269 163.367
R385 B.n271 B.n270 163.367
R386 B.n271 B.n84 163.367
R387 B.n275 B.n84 163.367
R388 B.n276 B.n275 163.367
R389 B.n277 B.n276 163.367
R390 B.n277 B.n82 163.367
R391 B.n281 B.n82 163.367
R392 B.n282 B.n281 163.367
R393 B.n283 B.n282 163.367
R394 B.n283 B.n80 163.367
R395 B.n287 B.n80 163.367
R396 B.n288 B.n287 163.367
R397 B.n289 B.n78 163.367
R398 B.n293 B.n78 163.367
R399 B.n294 B.n293 163.367
R400 B.n295 B.n294 163.367
R401 B.n295 B.n76 163.367
R402 B.n299 B.n76 163.367
R403 B.n300 B.n299 163.367
R404 B.n301 B.n300 163.367
R405 B.n301 B.n74 163.367
R406 B.n305 B.n74 163.367
R407 B.n306 B.n305 163.367
R408 B.n307 B.n306 163.367
R409 B.n307 B.n72 163.367
R410 B.n311 B.n72 163.367
R411 B.n312 B.n311 163.367
R412 B.n313 B.n312 163.367
R413 B.n313 B.n70 163.367
R414 B.n317 B.n70 163.367
R415 B.n318 B.n317 163.367
R416 B.n319 B.n318 163.367
R417 B.n319 B.n68 163.367
R418 B.n323 B.n68 163.367
R419 B.n324 B.n323 163.367
R420 B.n325 B.n324 163.367
R421 B.n325 B.n66 163.367
R422 B.n329 B.n66 163.367
R423 B.n330 B.n329 163.367
R424 B.n331 B.n330 163.367
R425 B.n331 B.n64 163.367
R426 B.n335 B.n64 163.367
R427 B.n336 B.n335 163.367
R428 B.n337 B.n336 163.367
R429 B.n337 B.n62 163.367
R430 B.n341 B.n62 163.367
R431 B.n342 B.n341 163.367
R432 B.n343 B.n342 163.367
R433 B.n343 B.n60 163.367
R434 B.n347 B.n60 163.367
R435 B.n348 B.n347 163.367
R436 B.n349 B.n348 163.367
R437 B.n475 B.n474 163.367
R438 B.n474 B.n13 163.367
R439 B.n470 B.n13 163.367
R440 B.n470 B.n469 163.367
R441 B.n469 B.n468 163.367
R442 B.n468 B.n15 163.367
R443 B.n464 B.n15 163.367
R444 B.n464 B.n463 163.367
R445 B.n463 B.n462 163.367
R446 B.n462 B.n17 163.367
R447 B.n458 B.n17 163.367
R448 B.n458 B.n457 163.367
R449 B.n457 B.n456 163.367
R450 B.n456 B.n19 163.367
R451 B.n452 B.n19 163.367
R452 B.n452 B.n451 163.367
R453 B.n451 B.n450 163.367
R454 B.n450 B.n21 163.367
R455 B.n446 B.n21 163.367
R456 B.n446 B.n445 163.367
R457 B.n445 B.n444 163.367
R458 B.n444 B.n23 163.367
R459 B.n440 B.n23 163.367
R460 B.n440 B.n439 163.367
R461 B.n439 B.n438 163.367
R462 B.n438 B.n25 163.367
R463 B.n434 B.n25 163.367
R464 B.n434 B.n433 163.367
R465 B.n433 B.n432 163.367
R466 B.n432 B.n27 163.367
R467 B.n428 B.n27 163.367
R468 B.n428 B.n427 163.367
R469 B.n427 B.n426 163.367
R470 B.n426 B.n29 163.367
R471 B.n422 B.n29 163.367
R472 B.n422 B.n421 163.367
R473 B.n421 B.n420 163.367
R474 B.n420 B.n31 163.367
R475 B.n416 B.n31 163.367
R476 B.n416 B.n415 163.367
R477 B.n415 B.n414 163.367
R478 B.n414 B.n36 163.367
R479 B.n410 B.n36 163.367
R480 B.n410 B.n409 163.367
R481 B.n409 B.n408 163.367
R482 B.n408 B.n38 163.367
R483 B.n403 B.n38 163.367
R484 B.n403 B.n402 163.367
R485 B.n402 B.n401 163.367
R486 B.n401 B.n42 163.367
R487 B.n397 B.n42 163.367
R488 B.n397 B.n396 163.367
R489 B.n396 B.n395 163.367
R490 B.n395 B.n44 163.367
R491 B.n391 B.n44 163.367
R492 B.n391 B.n390 163.367
R493 B.n390 B.n389 163.367
R494 B.n389 B.n46 163.367
R495 B.n385 B.n46 163.367
R496 B.n385 B.n384 163.367
R497 B.n384 B.n383 163.367
R498 B.n383 B.n48 163.367
R499 B.n379 B.n48 163.367
R500 B.n379 B.n378 163.367
R501 B.n378 B.n377 163.367
R502 B.n377 B.n50 163.367
R503 B.n373 B.n50 163.367
R504 B.n373 B.n372 163.367
R505 B.n372 B.n371 163.367
R506 B.n371 B.n52 163.367
R507 B.n367 B.n52 163.367
R508 B.n367 B.n366 163.367
R509 B.n366 B.n365 163.367
R510 B.n365 B.n54 163.367
R511 B.n361 B.n54 163.367
R512 B.n361 B.n360 163.367
R513 B.n360 B.n359 163.367
R514 B.n359 B.n56 163.367
R515 B.n355 B.n56 163.367
R516 B.n355 B.n354 163.367
R517 B.n354 B.n353 163.367
R518 B.n353 B.n58 163.367
R519 B.n229 B.t2 150.026
R520 B.n39 B.t10 150.026
R521 B.n103 B.t8 150.014
R522 B.n32 B.t4 150.014
R523 B.n230 B.t1 110.656
R524 B.n40 B.t11 110.656
R525 B.n104 B.t7 110.644
R526 B.n33 B.t5 110.644
R527 B.n231 B.n230 59.5399
R528 B.n216 B.n104 59.5399
R529 B.n34 B.n33 59.5399
R530 B.n406 B.n40 59.5399
R531 B.n230 B.n229 39.3702
R532 B.n104 B.n103 39.3702
R533 B.n33 B.n32 39.3702
R534 B.n40 B.n39 39.3702
R535 B.n477 B.n12 33.8737
R536 B.n351 B.n350 33.8737
R537 B.n290 B.n79 33.8737
R538 B.n161 B.n160 33.8737
R539 B B.n507 18.0485
R540 B.n473 B.n12 10.6151
R541 B.n473 B.n472 10.6151
R542 B.n472 B.n471 10.6151
R543 B.n471 B.n14 10.6151
R544 B.n467 B.n14 10.6151
R545 B.n467 B.n466 10.6151
R546 B.n466 B.n465 10.6151
R547 B.n465 B.n16 10.6151
R548 B.n461 B.n16 10.6151
R549 B.n461 B.n460 10.6151
R550 B.n460 B.n459 10.6151
R551 B.n459 B.n18 10.6151
R552 B.n455 B.n18 10.6151
R553 B.n455 B.n454 10.6151
R554 B.n454 B.n453 10.6151
R555 B.n453 B.n20 10.6151
R556 B.n449 B.n20 10.6151
R557 B.n449 B.n448 10.6151
R558 B.n448 B.n447 10.6151
R559 B.n447 B.n22 10.6151
R560 B.n443 B.n22 10.6151
R561 B.n443 B.n442 10.6151
R562 B.n442 B.n441 10.6151
R563 B.n441 B.n24 10.6151
R564 B.n437 B.n24 10.6151
R565 B.n437 B.n436 10.6151
R566 B.n436 B.n435 10.6151
R567 B.n435 B.n26 10.6151
R568 B.n431 B.n26 10.6151
R569 B.n431 B.n430 10.6151
R570 B.n430 B.n429 10.6151
R571 B.n429 B.n28 10.6151
R572 B.n425 B.n28 10.6151
R573 B.n425 B.n424 10.6151
R574 B.n424 B.n423 10.6151
R575 B.n423 B.n30 10.6151
R576 B.n419 B.n418 10.6151
R577 B.n418 B.n417 10.6151
R578 B.n417 B.n35 10.6151
R579 B.n413 B.n35 10.6151
R580 B.n413 B.n412 10.6151
R581 B.n412 B.n411 10.6151
R582 B.n411 B.n37 10.6151
R583 B.n407 B.n37 10.6151
R584 B.n405 B.n404 10.6151
R585 B.n404 B.n41 10.6151
R586 B.n400 B.n41 10.6151
R587 B.n400 B.n399 10.6151
R588 B.n399 B.n398 10.6151
R589 B.n398 B.n43 10.6151
R590 B.n394 B.n43 10.6151
R591 B.n394 B.n393 10.6151
R592 B.n393 B.n392 10.6151
R593 B.n392 B.n45 10.6151
R594 B.n388 B.n45 10.6151
R595 B.n388 B.n387 10.6151
R596 B.n387 B.n386 10.6151
R597 B.n386 B.n47 10.6151
R598 B.n382 B.n47 10.6151
R599 B.n382 B.n381 10.6151
R600 B.n381 B.n380 10.6151
R601 B.n380 B.n49 10.6151
R602 B.n376 B.n49 10.6151
R603 B.n376 B.n375 10.6151
R604 B.n375 B.n374 10.6151
R605 B.n374 B.n51 10.6151
R606 B.n370 B.n51 10.6151
R607 B.n370 B.n369 10.6151
R608 B.n369 B.n368 10.6151
R609 B.n368 B.n53 10.6151
R610 B.n364 B.n53 10.6151
R611 B.n364 B.n363 10.6151
R612 B.n363 B.n362 10.6151
R613 B.n362 B.n55 10.6151
R614 B.n358 B.n55 10.6151
R615 B.n358 B.n357 10.6151
R616 B.n357 B.n356 10.6151
R617 B.n356 B.n57 10.6151
R618 B.n352 B.n57 10.6151
R619 B.n352 B.n351 10.6151
R620 B.n291 B.n290 10.6151
R621 B.n292 B.n291 10.6151
R622 B.n292 B.n77 10.6151
R623 B.n296 B.n77 10.6151
R624 B.n297 B.n296 10.6151
R625 B.n298 B.n297 10.6151
R626 B.n298 B.n75 10.6151
R627 B.n302 B.n75 10.6151
R628 B.n303 B.n302 10.6151
R629 B.n304 B.n303 10.6151
R630 B.n304 B.n73 10.6151
R631 B.n308 B.n73 10.6151
R632 B.n309 B.n308 10.6151
R633 B.n310 B.n309 10.6151
R634 B.n310 B.n71 10.6151
R635 B.n314 B.n71 10.6151
R636 B.n315 B.n314 10.6151
R637 B.n316 B.n315 10.6151
R638 B.n316 B.n69 10.6151
R639 B.n320 B.n69 10.6151
R640 B.n321 B.n320 10.6151
R641 B.n322 B.n321 10.6151
R642 B.n322 B.n67 10.6151
R643 B.n326 B.n67 10.6151
R644 B.n327 B.n326 10.6151
R645 B.n328 B.n327 10.6151
R646 B.n328 B.n65 10.6151
R647 B.n332 B.n65 10.6151
R648 B.n333 B.n332 10.6151
R649 B.n334 B.n333 10.6151
R650 B.n334 B.n63 10.6151
R651 B.n338 B.n63 10.6151
R652 B.n339 B.n338 10.6151
R653 B.n340 B.n339 10.6151
R654 B.n340 B.n61 10.6151
R655 B.n344 B.n61 10.6151
R656 B.n345 B.n344 10.6151
R657 B.n346 B.n345 10.6151
R658 B.n346 B.n59 10.6151
R659 B.n350 B.n59 10.6151
R660 B.n162 B.n161 10.6151
R661 B.n162 B.n121 10.6151
R662 B.n166 B.n121 10.6151
R663 B.n167 B.n166 10.6151
R664 B.n168 B.n167 10.6151
R665 B.n168 B.n119 10.6151
R666 B.n172 B.n119 10.6151
R667 B.n173 B.n172 10.6151
R668 B.n174 B.n173 10.6151
R669 B.n174 B.n117 10.6151
R670 B.n178 B.n117 10.6151
R671 B.n179 B.n178 10.6151
R672 B.n180 B.n179 10.6151
R673 B.n180 B.n115 10.6151
R674 B.n184 B.n115 10.6151
R675 B.n185 B.n184 10.6151
R676 B.n186 B.n185 10.6151
R677 B.n186 B.n113 10.6151
R678 B.n190 B.n113 10.6151
R679 B.n191 B.n190 10.6151
R680 B.n192 B.n191 10.6151
R681 B.n192 B.n111 10.6151
R682 B.n196 B.n111 10.6151
R683 B.n197 B.n196 10.6151
R684 B.n198 B.n197 10.6151
R685 B.n198 B.n109 10.6151
R686 B.n202 B.n109 10.6151
R687 B.n203 B.n202 10.6151
R688 B.n204 B.n203 10.6151
R689 B.n204 B.n107 10.6151
R690 B.n208 B.n107 10.6151
R691 B.n209 B.n208 10.6151
R692 B.n210 B.n209 10.6151
R693 B.n210 B.n105 10.6151
R694 B.n214 B.n105 10.6151
R695 B.n215 B.n214 10.6151
R696 B.n217 B.n101 10.6151
R697 B.n221 B.n101 10.6151
R698 B.n222 B.n221 10.6151
R699 B.n223 B.n222 10.6151
R700 B.n223 B.n99 10.6151
R701 B.n227 B.n99 10.6151
R702 B.n228 B.n227 10.6151
R703 B.n232 B.n228 10.6151
R704 B.n236 B.n97 10.6151
R705 B.n237 B.n236 10.6151
R706 B.n238 B.n237 10.6151
R707 B.n238 B.n95 10.6151
R708 B.n242 B.n95 10.6151
R709 B.n243 B.n242 10.6151
R710 B.n244 B.n243 10.6151
R711 B.n244 B.n93 10.6151
R712 B.n248 B.n93 10.6151
R713 B.n249 B.n248 10.6151
R714 B.n250 B.n249 10.6151
R715 B.n250 B.n91 10.6151
R716 B.n254 B.n91 10.6151
R717 B.n255 B.n254 10.6151
R718 B.n256 B.n255 10.6151
R719 B.n256 B.n89 10.6151
R720 B.n260 B.n89 10.6151
R721 B.n261 B.n260 10.6151
R722 B.n262 B.n261 10.6151
R723 B.n262 B.n87 10.6151
R724 B.n266 B.n87 10.6151
R725 B.n267 B.n266 10.6151
R726 B.n268 B.n267 10.6151
R727 B.n268 B.n85 10.6151
R728 B.n272 B.n85 10.6151
R729 B.n273 B.n272 10.6151
R730 B.n274 B.n273 10.6151
R731 B.n274 B.n83 10.6151
R732 B.n278 B.n83 10.6151
R733 B.n279 B.n278 10.6151
R734 B.n280 B.n279 10.6151
R735 B.n280 B.n81 10.6151
R736 B.n284 B.n81 10.6151
R737 B.n285 B.n284 10.6151
R738 B.n286 B.n285 10.6151
R739 B.n286 B.n79 10.6151
R740 B.n160 B.n123 10.6151
R741 B.n156 B.n123 10.6151
R742 B.n156 B.n155 10.6151
R743 B.n155 B.n154 10.6151
R744 B.n154 B.n125 10.6151
R745 B.n150 B.n125 10.6151
R746 B.n150 B.n149 10.6151
R747 B.n149 B.n148 10.6151
R748 B.n148 B.n127 10.6151
R749 B.n144 B.n127 10.6151
R750 B.n144 B.n143 10.6151
R751 B.n143 B.n142 10.6151
R752 B.n142 B.n129 10.6151
R753 B.n138 B.n129 10.6151
R754 B.n138 B.n137 10.6151
R755 B.n137 B.n136 10.6151
R756 B.n136 B.n131 10.6151
R757 B.n132 B.n131 10.6151
R758 B.n132 B.n0 10.6151
R759 B.n503 B.n1 10.6151
R760 B.n503 B.n502 10.6151
R761 B.n502 B.n501 10.6151
R762 B.n501 B.n4 10.6151
R763 B.n497 B.n4 10.6151
R764 B.n497 B.n496 10.6151
R765 B.n496 B.n495 10.6151
R766 B.n495 B.n6 10.6151
R767 B.n491 B.n6 10.6151
R768 B.n491 B.n490 10.6151
R769 B.n490 B.n489 10.6151
R770 B.n489 B.n8 10.6151
R771 B.n485 B.n8 10.6151
R772 B.n485 B.n484 10.6151
R773 B.n484 B.n483 10.6151
R774 B.n483 B.n10 10.6151
R775 B.n479 B.n10 10.6151
R776 B.n479 B.n478 10.6151
R777 B.n478 B.n477 10.6151
R778 B.n419 B.n34 6.5566
R779 B.n407 B.n406 6.5566
R780 B.n217 B.n216 6.5566
R781 B.n232 B.n231 6.5566
R782 B.n34 B.n30 4.05904
R783 B.n406 B.n405 4.05904
R784 B.n216 B.n215 4.05904
R785 B.n231 B.n97 4.05904
R786 B.n507 B.n0 2.81026
R787 B.n507 B.n1 2.81026
C0 VTAIL w_n1782_n3040# 2.54009f
C1 VDD1 VN 0.148043f
C2 w_n1782_n3040# B 7.37659f
C3 VDD1 VP 2.39686f
C4 VDD1 VDD2 0.568488f
C5 VTAIL VN 1.92766f
C6 VTAIL VP 1.94201f
C7 VTAIL VDD2 4.60437f
C8 VN B 0.881556f
C9 VN w_n1782_n3040# 2.3574f
C10 VP B 1.24794f
C11 VDD2 B 1.47484f
C12 VTAIL VDD1 4.56053f
C13 VP w_n1782_n3040# 2.58246f
C14 VDD2 w_n1782_n3040# 1.57944f
C15 VDD1 B 1.45272f
C16 VDD1 w_n1782_n3040# 1.56436f
C17 VP VN 4.72956f
C18 VDD2 VN 2.25215f
C19 VTAIL B 2.91796f
C20 VDD2 VP 0.295512f
C21 VDD2 VSUBS 0.766056f
C22 VDD1 VSUBS 4.048916f
C23 VTAIL VSUBS 0.813816f
C24 VN VSUBS 6.480761f
C25 VP VSUBS 1.354053f
C26 B VSUBS 3.088511f
C27 w_n1782_n3040# VSUBS 66.8678f
C28 B.n0 VSUBS 0.004352f
C29 B.n1 VSUBS 0.004352f
C30 B.n2 VSUBS 0.006881f
C31 B.n3 VSUBS 0.006881f
C32 B.n4 VSUBS 0.006881f
C33 B.n5 VSUBS 0.006881f
C34 B.n6 VSUBS 0.006881f
C35 B.n7 VSUBS 0.006881f
C36 B.n8 VSUBS 0.006881f
C37 B.n9 VSUBS 0.006881f
C38 B.n10 VSUBS 0.006881f
C39 B.n11 VSUBS 0.006881f
C40 B.n12 VSUBS 0.016849f
C41 B.n13 VSUBS 0.006881f
C42 B.n14 VSUBS 0.006881f
C43 B.n15 VSUBS 0.006881f
C44 B.n16 VSUBS 0.006881f
C45 B.n17 VSUBS 0.006881f
C46 B.n18 VSUBS 0.006881f
C47 B.n19 VSUBS 0.006881f
C48 B.n20 VSUBS 0.006881f
C49 B.n21 VSUBS 0.006881f
C50 B.n22 VSUBS 0.006881f
C51 B.n23 VSUBS 0.006881f
C52 B.n24 VSUBS 0.006881f
C53 B.n25 VSUBS 0.006881f
C54 B.n26 VSUBS 0.006881f
C55 B.n27 VSUBS 0.006881f
C56 B.n28 VSUBS 0.006881f
C57 B.n29 VSUBS 0.006881f
C58 B.n30 VSUBS 0.004756f
C59 B.n31 VSUBS 0.006881f
C60 B.t5 VSUBS 0.326285f
C61 B.t4 VSUBS 0.341236f
C62 B.t3 VSUBS 0.772365f
C63 B.n32 VSUBS 0.160982f
C64 B.n33 VSUBS 0.066782f
C65 B.n34 VSUBS 0.015944f
C66 B.n35 VSUBS 0.006881f
C67 B.n36 VSUBS 0.006881f
C68 B.n37 VSUBS 0.006881f
C69 B.n38 VSUBS 0.006881f
C70 B.t11 VSUBS 0.32628f
C71 B.t10 VSUBS 0.341231f
C72 B.t9 VSUBS 0.772365f
C73 B.n39 VSUBS 0.160987f
C74 B.n40 VSUBS 0.066787f
C75 B.n41 VSUBS 0.006881f
C76 B.n42 VSUBS 0.006881f
C77 B.n43 VSUBS 0.006881f
C78 B.n44 VSUBS 0.006881f
C79 B.n45 VSUBS 0.006881f
C80 B.n46 VSUBS 0.006881f
C81 B.n47 VSUBS 0.006881f
C82 B.n48 VSUBS 0.006881f
C83 B.n49 VSUBS 0.006881f
C84 B.n50 VSUBS 0.006881f
C85 B.n51 VSUBS 0.006881f
C86 B.n52 VSUBS 0.006881f
C87 B.n53 VSUBS 0.006881f
C88 B.n54 VSUBS 0.006881f
C89 B.n55 VSUBS 0.006881f
C90 B.n56 VSUBS 0.006881f
C91 B.n57 VSUBS 0.006881f
C92 B.n58 VSUBS 0.016849f
C93 B.n59 VSUBS 0.006881f
C94 B.n60 VSUBS 0.006881f
C95 B.n61 VSUBS 0.006881f
C96 B.n62 VSUBS 0.006881f
C97 B.n63 VSUBS 0.006881f
C98 B.n64 VSUBS 0.006881f
C99 B.n65 VSUBS 0.006881f
C100 B.n66 VSUBS 0.006881f
C101 B.n67 VSUBS 0.006881f
C102 B.n68 VSUBS 0.006881f
C103 B.n69 VSUBS 0.006881f
C104 B.n70 VSUBS 0.006881f
C105 B.n71 VSUBS 0.006881f
C106 B.n72 VSUBS 0.006881f
C107 B.n73 VSUBS 0.006881f
C108 B.n74 VSUBS 0.006881f
C109 B.n75 VSUBS 0.006881f
C110 B.n76 VSUBS 0.006881f
C111 B.n77 VSUBS 0.006881f
C112 B.n78 VSUBS 0.006881f
C113 B.n79 VSUBS 0.016849f
C114 B.n80 VSUBS 0.006881f
C115 B.n81 VSUBS 0.006881f
C116 B.n82 VSUBS 0.006881f
C117 B.n83 VSUBS 0.006881f
C118 B.n84 VSUBS 0.006881f
C119 B.n85 VSUBS 0.006881f
C120 B.n86 VSUBS 0.006881f
C121 B.n87 VSUBS 0.006881f
C122 B.n88 VSUBS 0.006881f
C123 B.n89 VSUBS 0.006881f
C124 B.n90 VSUBS 0.006881f
C125 B.n91 VSUBS 0.006881f
C126 B.n92 VSUBS 0.006881f
C127 B.n93 VSUBS 0.006881f
C128 B.n94 VSUBS 0.006881f
C129 B.n95 VSUBS 0.006881f
C130 B.n96 VSUBS 0.006881f
C131 B.n97 VSUBS 0.004756f
C132 B.n98 VSUBS 0.006881f
C133 B.n99 VSUBS 0.006881f
C134 B.n100 VSUBS 0.006881f
C135 B.n101 VSUBS 0.006881f
C136 B.n102 VSUBS 0.006881f
C137 B.t7 VSUBS 0.326285f
C138 B.t8 VSUBS 0.341236f
C139 B.t6 VSUBS 0.772365f
C140 B.n103 VSUBS 0.160982f
C141 B.n104 VSUBS 0.066782f
C142 B.n105 VSUBS 0.006881f
C143 B.n106 VSUBS 0.006881f
C144 B.n107 VSUBS 0.006881f
C145 B.n108 VSUBS 0.006881f
C146 B.n109 VSUBS 0.006881f
C147 B.n110 VSUBS 0.006881f
C148 B.n111 VSUBS 0.006881f
C149 B.n112 VSUBS 0.006881f
C150 B.n113 VSUBS 0.006881f
C151 B.n114 VSUBS 0.006881f
C152 B.n115 VSUBS 0.006881f
C153 B.n116 VSUBS 0.006881f
C154 B.n117 VSUBS 0.006881f
C155 B.n118 VSUBS 0.006881f
C156 B.n119 VSUBS 0.006881f
C157 B.n120 VSUBS 0.006881f
C158 B.n121 VSUBS 0.006881f
C159 B.n122 VSUBS 0.016849f
C160 B.n123 VSUBS 0.006881f
C161 B.n124 VSUBS 0.006881f
C162 B.n125 VSUBS 0.006881f
C163 B.n126 VSUBS 0.006881f
C164 B.n127 VSUBS 0.006881f
C165 B.n128 VSUBS 0.006881f
C166 B.n129 VSUBS 0.006881f
C167 B.n130 VSUBS 0.006881f
C168 B.n131 VSUBS 0.006881f
C169 B.n132 VSUBS 0.006881f
C170 B.n133 VSUBS 0.006881f
C171 B.n134 VSUBS 0.006881f
C172 B.n135 VSUBS 0.006881f
C173 B.n136 VSUBS 0.006881f
C174 B.n137 VSUBS 0.006881f
C175 B.n138 VSUBS 0.006881f
C176 B.n139 VSUBS 0.006881f
C177 B.n140 VSUBS 0.006881f
C178 B.n141 VSUBS 0.006881f
C179 B.n142 VSUBS 0.006881f
C180 B.n143 VSUBS 0.006881f
C181 B.n144 VSUBS 0.006881f
C182 B.n145 VSUBS 0.006881f
C183 B.n146 VSUBS 0.006881f
C184 B.n147 VSUBS 0.006881f
C185 B.n148 VSUBS 0.006881f
C186 B.n149 VSUBS 0.006881f
C187 B.n150 VSUBS 0.006881f
C188 B.n151 VSUBS 0.006881f
C189 B.n152 VSUBS 0.006881f
C190 B.n153 VSUBS 0.006881f
C191 B.n154 VSUBS 0.006881f
C192 B.n155 VSUBS 0.006881f
C193 B.n156 VSUBS 0.006881f
C194 B.n157 VSUBS 0.006881f
C195 B.n158 VSUBS 0.006881f
C196 B.n159 VSUBS 0.016142f
C197 B.n160 VSUBS 0.016142f
C198 B.n161 VSUBS 0.016849f
C199 B.n162 VSUBS 0.006881f
C200 B.n163 VSUBS 0.006881f
C201 B.n164 VSUBS 0.006881f
C202 B.n165 VSUBS 0.006881f
C203 B.n166 VSUBS 0.006881f
C204 B.n167 VSUBS 0.006881f
C205 B.n168 VSUBS 0.006881f
C206 B.n169 VSUBS 0.006881f
C207 B.n170 VSUBS 0.006881f
C208 B.n171 VSUBS 0.006881f
C209 B.n172 VSUBS 0.006881f
C210 B.n173 VSUBS 0.006881f
C211 B.n174 VSUBS 0.006881f
C212 B.n175 VSUBS 0.006881f
C213 B.n176 VSUBS 0.006881f
C214 B.n177 VSUBS 0.006881f
C215 B.n178 VSUBS 0.006881f
C216 B.n179 VSUBS 0.006881f
C217 B.n180 VSUBS 0.006881f
C218 B.n181 VSUBS 0.006881f
C219 B.n182 VSUBS 0.006881f
C220 B.n183 VSUBS 0.006881f
C221 B.n184 VSUBS 0.006881f
C222 B.n185 VSUBS 0.006881f
C223 B.n186 VSUBS 0.006881f
C224 B.n187 VSUBS 0.006881f
C225 B.n188 VSUBS 0.006881f
C226 B.n189 VSUBS 0.006881f
C227 B.n190 VSUBS 0.006881f
C228 B.n191 VSUBS 0.006881f
C229 B.n192 VSUBS 0.006881f
C230 B.n193 VSUBS 0.006881f
C231 B.n194 VSUBS 0.006881f
C232 B.n195 VSUBS 0.006881f
C233 B.n196 VSUBS 0.006881f
C234 B.n197 VSUBS 0.006881f
C235 B.n198 VSUBS 0.006881f
C236 B.n199 VSUBS 0.006881f
C237 B.n200 VSUBS 0.006881f
C238 B.n201 VSUBS 0.006881f
C239 B.n202 VSUBS 0.006881f
C240 B.n203 VSUBS 0.006881f
C241 B.n204 VSUBS 0.006881f
C242 B.n205 VSUBS 0.006881f
C243 B.n206 VSUBS 0.006881f
C244 B.n207 VSUBS 0.006881f
C245 B.n208 VSUBS 0.006881f
C246 B.n209 VSUBS 0.006881f
C247 B.n210 VSUBS 0.006881f
C248 B.n211 VSUBS 0.006881f
C249 B.n212 VSUBS 0.006881f
C250 B.n213 VSUBS 0.006881f
C251 B.n214 VSUBS 0.006881f
C252 B.n215 VSUBS 0.004756f
C253 B.n216 VSUBS 0.015944f
C254 B.n217 VSUBS 0.005566f
C255 B.n218 VSUBS 0.006881f
C256 B.n219 VSUBS 0.006881f
C257 B.n220 VSUBS 0.006881f
C258 B.n221 VSUBS 0.006881f
C259 B.n222 VSUBS 0.006881f
C260 B.n223 VSUBS 0.006881f
C261 B.n224 VSUBS 0.006881f
C262 B.n225 VSUBS 0.006881f
C263 B.n226 VSUBS 0.006881f
C264 B.n227 VSUBS 0.006881f
C265 B.n228 VSUBS 0.006881f
C266 B.t1 VSUBS 0.32628f
C267 B.t2 VSUBS 0.341231f
C268 B.t0 VSUBS 0.772365f
C269 B.n229 VSUBS 0.160987f
C270 B.n230 VSUBS 0.066787f
C271 B.n231 VSUBS 0.015944f
C272 B.n232 VSUBS 0.005566f
C273 B.n233 VSUBS 0.006881f
C274 B.n234 VSUBS 0.006881f
C275 B.n235 VSUBS 0.006881f
C276 B.n236 VSUBS 0.006881f
C277 B.n237 VSUBS 0.006881f
C278 B.n238 VSUBS 0.006881f
C279 B.n239 VSUBS 0.006881f
C280 B.n240 VSUBS 0.006881f
C281 B.n241 VSUBS 0.006881f
C282 B.n242 VSUBS 0.006881f
C283 B.n243 VSUBS 0.006881f
C284 B.n244 VSUBS 0.006881f
C285 B.n245 VSUBS 0.006881f
C286 B.n246 VSUBS 0.006881f
C287 B.n247 VSUBS 0.006881f
C288 B.n248 VSUBS 0.006881f
C289 B.n249 VSUBS 0.006881f
C290 B.n250 VSUBS 0.006881f
C291 B.n251 VSUBS 0.006881f
C292 B.n252 VSUBS 0.006881f
C293 B.n253 VSUBS 0.006881f
C294 B.n254 VSUBS 0.006881f
C295 B.n255 VSUBS 0.006881f
C296 B.n256 VSUBS 0.006881f
C297 B.n257 VSUBS 0.006881f
C298 B.n258 VSUBS 0.006881f
C299 B.n259 VSUBS 0.006881f
C300 B.n260 VSUBS 0.006881f
C301 B.n261 VSUBS 0.006881f
C302 B.n262 VSUBS 0.006881f
C303 B.n263 VSUBS 0.006881f
C304 B.n264 VSUBS 0.006881f
C305 B.n265 VSUBS 0.006881f
C306 B.n266 VSUBS 0.006881f
C307 B.n267 VSUBS 0.006881f
C308 B.n268 VSUBS 0.006881f
C309 B.n269 VSUBS 0.006881f
C310 B.n270 VSUBS 0.006881f
C311 B.n271 VSUBS 0.006881f
C312 B.n272 VSUBS 0.006881f
C313 B.n273 VSUBS 0.006881f
C314 B.n274 VSUBS 0.006881f
C315 B.n275 VSUBS 0.006881f
C316 B.n276 VSUBS 0.006881f
C317 B.n277 VSUBS 0.006881f
C318 B.n278 VSUBS 0.006881f
C319 B.n279 VSUBS 0.006881f
C320 B.n280 VSUBS 0.006881f
C321 B.n281 VSUBS 0.006881f
C322 B.n282 VSUBS 0.006881f
C323 B.n283 VSUBS 0.006881f
C324 B.n284 VSUBS 0.006881f
C325 B.n285 VSUBS 0.006881f
C326 B.n286 VSUBS 0.006881f
C327 B.n287 VSUBS 0.006881f
C328 B.n288 VSUBS 0.016849f
C329 B.n289 VSUBS 0.016142f
C330 B.n290 VSUBS 0.016142f
C331 B.n291 VSUBS 0.006881f
C332 B.n292 VSUBS 0.006881f
C333 B.n293 VSUBS 0.006881f
C334 B.n294 VSUBS 0.006881f
C335 B.n295 VSUBS 0.006881f
C336 B.n296 VSUBS 0.006881f
C337 B.n297 VSUBS 0.006881f
C338 B.n298 VSUBS 0.006881f
C339 B.n299 VSUBS 0.006881f
C340 B.n300 VSUBS 0.006881f
C341 B.n301 VSUBS 0.006881f
C342 B.n302 VSUBS 0.006881f
C343 B.n303 VSUBS 0.006881f
C344 B.n304 VSUBS 0.006881f
C345 B.n305 VSUBS 0.006881f
C346 B.n306 VSUBS 0.006881f
C347 B.n307 VSUBS 0.006881f
C348 B.n308 VSUBS 0.006881f
C349 B.n309 VSUBS 0.006881f
C350 B.n310 VSUBS 0.006881f
C351 B.n311 VSUBS 0.006881f
C352 B.n312 VSUBS 0.006881f
C353 B.n313 VSUBS 0.006881f
C354 B.n314 VSUBS 0.006881f
C355 B.n315 VSUBS 0.006881f
C356 B.n316 VSUBS 0.006881f
C357 B.n317 VSUBS 0.006881f
C358 B.n318 VSUBS 0.006881f
C359 B.n319 VSUBS 0.006881f
C360 B.n320 VSUBS 0.006881f
C361 B.n321 VSUBS 0.006881f
C362 B.n322 VSUBS 0.006881f
C363 B.n323 VSUBS 0.006881f
C364 B.n324 VSUBS 0.006881f
C365 B.n325 VSUBS 0.006881f
C366 B.n326 VSUBS 0.006881f
C367 B.n327 VSUBS 0.006881f
C368 B.n328 VSUBS 0.006881f
C369 B.n329 VSUBS 0.006881f
C370 B.n330 VSUBS 0.006881f
C371 B.n331 VSUBS 0.006881f
C372 B.n332 VSUBS 0.006881f
C373 B.n333 VSUBS 0.006881f
C374 B.n334 VSUBS 0.006881f
C375 B.n335 VSUBS 0.006881f
C376 B.n336 VSUBS 0.006881f
C377 B.n337 VSUBS 0.006881f
C378 B.n338 VSUBS 0.006881f
C379 B.n339 VSUBS 0.006881f
C380 B.n340 VSUBS 0.006881f
C381 B.n341 VSUBS 0.006881f
C382 B.n342 VSUBS 0.006881f
C383 B.n343 VSUBS 0.006881f
C384 B.n344 VSUBS 0.006881f
C385 B.n345 VSUBS 0.006881f
C386 B.n346 VSUBS 0.006881f
C387 B.n347 VSUBS 0.006881f
C388 B.n348 VSUBS 0.006881f
C389 B.n349 VSUBS 0.016142f
C390 B.n350 VSUBS 0.016926f
C391 B.n351 VSUBS 0.016065f
C392 B.n352 VSUBS 0.006881f
C393 B.n353 VSUBS 0.006881f
C394 B.n354 VSUBS 0.006881f
C395 B.n355 VSUBS 0.006881f
C396 B.n356 VSUBS 0.006881f
C397 B.n357 VSUBS 0.006881f
C398 B.n358 VSUBS 0.006881f
C399 B.n359 VSUBS 0.006881f
C400 B.n360 VSUBS 0.006881f
C401 B.n361 VSUBS 0.006881f
C402 B.n362 VSUBS 0.006881f
C403 B.n363 VSUBS 0.006881f
C404 B.n364 VSUBS 0.006881f
C405 B.n365 VSUBS 0.006881f
C406 B.n366 VSUBS 0.006881f
C407 B.n367 VSUBS 0.006881f
C408 B.n368 VSUBS 0.006881f
C409 B.n369 VSUBS 0.006881f
C410 B.n370 VSUBS 0.006881f
C411 B.n371 VSUBS 0.006881f
C412 B.n372 VSUBS 0.006881f
C413 B.n373 VSUBS 0.006881f
C414 B.n374 VSUBS 0.006881f
C415 B.n375 VSUBS 0.006881f
C416 B.n376 VSUBS 0.006881f
C417 B.n377 VSUBS 0.006881f
C418 B.n378 VSUBS 0.006881f
C419 B.n379 VSUBS 0.006881f
C420 B.n380 VSUBS 0.006881f
C421 B.n381 VSUBS 0.006881f
C422 B.n382 VSUBS 0.006881f
C423 B.n383 VSUBS 0.006881f
C424 B.n384 VSUBS 0.006881f
C425 B.n385 VSUBS 0.006881f
C426 B.n386 VSUBS 0.006881f
C427 B.n387 VSUBS 0.006881f
C428 B.n388 VSUBS 0.006881f
C429 B.n389 VSUBS 0.006881f
C430 B.n390 VSUBS 0.006881f
C431 B.n391 VSUBS 0.006881f
C432 B.n392 VSUBS 0.006881f
C433 B.n393 VSUBS 0.006881f
C434 B.n394 VSUBS 0.006881f
C435 B.n395 VSUBS 0.006881f
C436 B.n396 VSUBS 0.006881f
C437 B.n397 VSUBS 0.006881f
C438 B.n398 VSUBS 0.006881f
C439 B.n399 VSUBS 0.006881f
C440 B.n400 VSUBS 0.006881f
C441 B.n401 VSUBS 0.006881f
C442 B.n402 VSUBS 0.006881f
C443 B.n403 VSUBS 0.006881f
C444 B.n404 VSUBS 0.006881f
C445 B.n405 VSUBS 0.004756f
C446 B.n406 VSUBS 0.015944f
C447 B.n407 VSUBS 0.005566f
C448 B.n408 VSUBS 0.006881f
C449 B.n409 VSUBS 0.006881f
C450 B.n410 VSUBS 0.006881f
C451 B.n411 VSUBS 0.006881f
C452 B.n412 VSUBS 0.006881f
C453 B.n413 VSUBS 0.006881f
C454 B.n414 VSUBS 0.006881f
C455 B.n415 VSUBS 0.006881f
C456 B.n416 VSUBS 0.006881f
C457 B.n417 VSUBS 0.006881f
C458 B.n418 VSUBS 0.006881f
C459 B.n419 VSUBS 0.005566f
C460 B.n420 VSUBS 0.006881f
C461 B.n421 VSUBS 0.006881f
C462 B.n422 VSUBS 0.006881f
C463 B.n423 VSUBS 0.006881f
C464 B.n424 VSUBS 0.006881f
C465 B.n425 VSUBS 0.006881f
C466 B.n426 VSUBS 0.006881f
C467 B.n427 VSUBS 0.006881f
C468 B.n428 VSUBS 0.006881f
C469 B.n429 VSUBS 0.006881f
C470 B.n430 VSUBS 0.006881f
C471 B.n431 VSUBS 0.006881f
C472 B.n432 VSUBS 0.006881f
C473 B.n433 VSUBS 0.006881f
C474 B.n434 VSUBS 0.006881f
C475 B.n435 VSUBS 0.006881f
C476 B.n436 VSUBS 0.006881f
C477 B.n437 VSUBS 0.006881f
C478 B.n438 VSUBS 0.006881f
C479 B.n439 VSUBS 0.006881f
C480 B.n440 VSUBS 0.006881f
C481 B.n441 VSUBS 0.006881f
C482 B.n442 VSUBS 0.006881f
C483 B.n443 VSUBS 0.006881f
C484 B.n444 VSUBS 0.006881f
C485 B.n445 VSUBS 0.006881f
C486 B.n446 VSUBS 0.006881f
C487 B.n447 VSUBS 0.006881f
C488 B.n448 VSUBS 0.006881f
C489 B.n449 VSUBS 0.006881f
C490 B.n450 VSUBS 0.006881f
C491 B.n451 VSUBS 0.006881f
C492 B.n452 VSUBS 0.006881f
C493 B.n453 VSUBS 0.006881f
C494 B.n454 VSUBS 0.006881f
C495 B.n455 VSUBS 0.006881f
C496 B.n456 VSUBS 0.006881f
C497 B.n457 VSUBS 0.006881f
C498 B.n458 VSUBS 0.006881f
C499 B.n459 VSUBS 0.006881f
C500 B.n460 VSUBS 0.006881f
C501 B.n461 VSUBS 0.006881f
C502 B.n462 VSUBS 0.006881f
C503 B.n463 VSUBS 0.006881f
C504 B.n464 VSUBS 0.006881f
C505 B.n465 VSUBS 0.006881f
C506 B.n466 VSUBS 0.006881f
C507 B.n467 VSUBS 0.006881f
C508 B.n468 VSUBS 0.006881f
C509 B.n469 VSUBS 0.006881f
C510 B.n470 VSUBS 0.006881f
C511 B.n471 VSUBS 0.006881f
C512 B.n472 VSUBS 0.006881f
C513 B.n473 VSUBS 0.006881f
C514 B.n474 VSUBS 0.006881f
C515 B.n475 VSUBS 0.016849f
C516 B.n476 VSUBS 0.016142f
C517 B.n477 VSUBS 0.016142f
C518 B.n478 VSUBS 0.006881f
C519 B.n479 VSUBS 0.006881f
C520 B.n480 VSUBS 0.006881f
C521 B.n481 VSUBS 0.006881f
C522 B.n482 VSUBS 0.006881f
C523 B.n483 VSUBS 0.006881f
C524 B.n484 VSUBS 0.006881f
C525 B.n485 VSUBS 0.006881f
C526 B.n486 VSUBS 0.006881f
C527 B.n487 VSUBS 0.006881f
C528 B.n488 VSUBS 0.006881f
C529 B.n489 VSUBS 0.006881f
C530 B.n490 VSUBS 0.006881f
C531 B.n491 VSUBS 0.006881f
C532 B.n492 VSUBS 0.006881f
C533 B.n493 VSUBS 0.006881f
C534 B.n494 VSUBS 0.006881f
C535 B.n495 VSUBS 0.006881f
C536 B.n496 VSUBS 0.006881f
C537 B.n497 VSUBS 0.006881f
C538 B.n498 VSUBS 0.006881f
C539 B.n499 VSUBS 0.006881f
C540 B.n500 VSUBS 0.006881f
C541 B.n501 VSUBS 0.006881f
C542 B.n502 VSUBS 0.006881f
C543 B.n503 VSUBS 0.006881f
C544 B.n504 VSUBS 0.006881f
C545 B.n505 VSUBS 0.006881f
C546 B.n506 VSUBS 0.006881f
C547 B.n507 VSUBS 0.015582f
C548 VDD2.t1 VSUBS 2.12932f
C549 VDD2.t0 VSUBS 1.66829f
C550 VDD2.n0 VSUBS 3.01159f
C551 VN.t0 VSUBS 2.25457f
C552 VN.t1 VSUBS 2.65727f
C553 VDD1.t0 VSUBS 1.67706f
C554 VDD1.t1 VSUBS 2.16418f
C555 VTAIL.t2 VSUBS 1.77602f
C556 VTAIL.n0 VSUBS 1.91121f
C557 VTAIL.t3 VSUBS 1.77603f
C558 VTAIL.n1 VSUBS 1.9397f
C559 VTAIL.t1 VSUBS 1.77602f
C560 VTAIL.n2 VSUBS 1.80825f
C561 VTAIL.t0 VSUBS 1.77602f
C562 VTAIL.n3 VSUBS 1.73572f
C563 VP.t1 VSUBS 2.75429f
C564 VP.t0 VSUBS 2.34018f
C565 VP.n0 VSUBS 4.5432f
.ends

