* NGSPICE file created from diff_pair_sample_0079.ext - technology: sky130A

.subckt diff_pair_sample_0079 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=2.2935 pd=14.23 as=5.421 ps=28.58 w=13.9 l=1.82
X1 VDD1.t4 VP.t1 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=5.421 pd=28.58 as=2.2935 ps=14.23 w=13.9 l=1.82
X2 VDD2.t5 VN.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=5.421 pd=28.58 as=2.2935 ps=14.23 w=13.9 l=1.82
X3 VTAIL.t9 VP.t2 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=2.2935 pd=14.23 as=2.2935 ps=14.23 w=13.9 l=1.82
X4 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=5.421 pd=28.58 as=0 ps=0 w=13.9 l=1.82
X5 VTAIL.t6 VP.t3 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.2935 pd=14.23 as=2.2935 ps=14.23 w=13.9 l=1.82
X6 VDD1.t1 VP.t4 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=5.421 pd=28.58 as=2.2935 ps=14.23 w=13.9 l=1.82
X7 VDD1.t0 VP.t5 VTAIL.t8 B.t19 sky130_fd_pr__nfet_01v8 ad=2.2935 pd=14.23 as=5.421 ps=28.58 w=13.9 l=1.82
X8 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=5.421 pd=28.58 as=0 ps=0 w=13.9 l=1.82
X9 B.t11 B.t9 B.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=5.421 pd=28.58 as=0 ps=0 w=13.9 l=1.82
X10 VDD2.t4 VN.t1 VTAIL.t11 B.t19 sky130_fd_pr__nfet_01v8 ad=2.2935 pd=14.23 as=5.421 ps=28.58 w=13.9 l=1.82
X11 VTAIL.t3 VN.t2 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.2935 pd=14.23 as=2.2935 ps=14.23 w=13.9 l=1.82
X12 VDD2.t2 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.2935 pd=14.23 as=5.421 ps=28.58 w=13.9 l=1.82
X13 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=5.421 pd=28.58 as=0 ps=0 w=13.9 l=1.82
X14 VTAIL.t0 VN.t4 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.2935 pd=14.23 as=2.2935 ps=14.23 w=13.9 l=1.82
X15 VDD2.t0 VN.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.421 pd=28.58 as=2.2935 ps=14.23 w=13.9 l=1.82
R0 VP.n6 VP.t1 214.252
R1 VP.n17 VP.t4 184.06
R2 VP.n24 VP.t3 184.06
R3 VP.n31 VP.t5 184.06
R4 VP.n14 VP.t0 184.06
R5 VP.n7 VP.t2 184.06
R6 VP.n9 VP.n8 161.3
R7 VP.n10 VP.n5 161.3
R8 VP.n12 VP.n11 161.3
R9 VP.n13 VP.n4 161.3
R10 VP.n30 VP.n0 161.3
R11 VP.n29 VP.n28 161.3
R12 VP.n27 VP.n1 161.3
R13 VP.n26 VP.n25 161.3
R14 VP.n23 VP.n2 161.3
R15 VP.n22 VP.n21 161.3
R16 VP.n20 VP.n3 161.3
R17 VP.n19 VP.n18 161.3
R18 VP.n17 VP.n16 91.1314
R19 VP.n32 VP.n31 91.1314
R20 VP.n15 VP.n14 91.1314
R21 VP.n7 VP.n6 57.3616
R22 VP.n22 VP.n3 56.4773
R23 VP.n29 VP.n1 56.4773
R24 VP.n12 VP.n5 56.4773
R25 VP.n16 VP.n15 47.0336
R26 VP.n18 VP.n3 24.3439
R27 VP.n23 VP.n22 24.3439
R28 VP.n25 VP.n1 24.3439
R29 VP.n30 VP.n29 24.3439
R30 VP.n13 VP.n12 24.3439
R31 VP.n8 VP.n5 24.3439
R32 VP.n18 VP.n17 19.4752
R33 VP.n31 VP.n30 19.4752
R34 VP.n14 VP.n13 19.4752
R35 VP.n9 VP.n6 13.3877
R36 VP.n24 VP.n23 12.1722
R37 VP.n25 VP.n24 12.1722
R38 VP.n8 VP.n7 12.1722
R39 VP.n15 VP.n4 0.278398
R40 VP.n19 VP.n16 0.278398
R41 VP.n32 VP.n0 0.278398
R42 VP.n10 VP.n9 0.189894
R43 VP.n11 VP.n10 0.189894
R44 VP.n11 VP.n4 0.189894
R45 VP.n20 VP.n19 0.189894
R46 VP.n21 VP.n20 0.189894
R47 VP.n21 VP.n2 0.189894
R48 VP.n26 VP.n2 0.189894
R49 VP.n27 VP.n26 0.189894
R50 VP.n28 VP.n27 0.189894
R51 VP.n28 VP.n0 0.189894
R52 VP VP.n32 0.153422
R53 VTAIL.n10 VTAIL.t10 45.8461
R54 VTAIL.n7 VTAIL.t11 45.8461
R55 VTAIL.n11 VTAIL.t2 45.8459
R56 VTAIL.n2 VTAIL.t8 45.8459
R57 VTAIL.n9 VTAIL.n8 44.4216
R58 VTAIL.n6 VTAIL.n5 44.4216
R59 VTAIL.n1 VTAIL.n0 44.4216
R60 VTAIL.n4 VTAIL.n3 44.4216
R61 VTAIL.n6 VTAIL.n4 28.0565
R62 VTAIL.n11 VTAIL.n10 26.2031
R63 VTAIL.n7 VTAIL.n6 1.85395
R64 VTAIL.n10 VTAIL.n9 1.85395
R65 VTAIL.n4 VTAIL.n2 1.85395
R66 VTAIL.n0 VTAIL.t1 1.42496
R67 VTAIL.n0 VTAIL.t0 1.42496
R68 VTAIL.n3 VTAIL.t7 1.42496
R69 VTAIL.n3 VTAIL.t6 1.42496
R70 VTAIL.n8 VTAIL.t5 1.42496
R71 VTAIL.n8 VTAIL.t9 1.42496
R72 VTAIL.n5 VTAIL.t4 1.42496
R73 VTAIL.n5 VTAIL.t3 1.42496
R74 VTAIL.n9 VTAIL.n7 1.39705
R75 VTAIL.n2 VTAIL.n1 1.39705
R76 VTAIL VTAIL.n11 1.3324
R77 VTAIL VTAIL.n1 0.522052
R78 VDD1 VDD1.t4 63.9731
R79 VDD1.n1 VDD1.t1 63.8595
R80 VDD1.n1 VDD1.n0 61.5084
R81 VDD1.n3 VDD1.n2 61.1004
R82 VDD1.n3 VDD1.n1 43.2315
R83 VDD1.n2 VDD1.t3 1.42496
R84 VDD1.n2 VDD1.t5 1.42496
R85 VDD1.n0 VDD1.t2 1.42496
R86 VDD1.n0 VDD1.t0 1.42496
R87 VDD1 VDD1.n3 0.405672
R88 B.n800 B.n799 585
R89 B.n326 B.n115 585
R90 B.n325 B.n324 585
R91 B.n323 B.n322 585
R92 B.n321 B.n320 585
R93 B.n319 B.n318 585
R94 B.n317 B.n316 585
R95 B.n315 B.n314 585
R96 B.n313 B.n312 585
R97 B.n311 B.n310 585
R98 B.n309 B.n308 585
R99 B.n307 B.n306 585
R100 B.n305 B.n304 585
R101 B.n303 B.n302 585
R102 B.n301 B.n300 585
R103 B.n299 B.n298 585
R104 B.n297 B.n296 585
R105 B.n295 B.n294 585
R106 B.n293 B.n292 585
R107 B.n291 B.n290 585
R108 B.n289 B.n288 585
R109 B.n287 B.n286 585
R110 B.n285 B.n284 585
R111 B.n283 B.n282 585
R112 B.n281 B.n280 585
R113 B.n279 B.n278 585
R114 B.n277 B.n276 585
R115 B.n275 B.n274 585
R116 B.n273 B.n272 585
R117 B.n271 B.n270 585
R118 B.n269 B.n268 585
R119 B.n267 B.n266 585
R120 B.n265 B.n264 585
R121 B.n263 B.n262 585
R122 B.n261 B.n260 585
R123 B.n259 B.n258 585
R124 B.n257 B.n256 585
R125 B.n255 B.n254 585
R126 B.n253 B.n252 585
R127 B.n251 B.n250 585
R128 B.n249 B.n248 585
R129 B.n247 B.n246 585
R130 B.n245 B.n244 585
R131 B.n243 B.n242 585
R132 B.n241 B.n240 585
R133 B.n239 B.n238 585
R134 B.n237 B.n236 585
R135 B.n234 B.n233 585
R136 B.n232 B.n231 585
R137 B.n230 B.n229 585
R138 B.n228 B.n227 585
R139 B.n226 B.n225 585
R140 B.n224 B.n223 585
R141 B.n222 B.n221 585
R142 B.n220 B.n219 585
R143 B.n218 B.n217 585
R144 B.n216 B.n215 585
R145 B.n213 B.n212 585
R146 B.n211 B.n210 585
R147 B.n209 B.n208 585
R148 B.n207 B.n206 585
R149 B.n205 B.n204 585
R150 B.n203 B.n202 585
R151 B.n201 B.n200 585
R152 B.n199 B.n198 585
R153 B.n197 B.n196 585
R154 B.n195 B.n194 585
R155 B.n193 B.n192 585
R156 B.n191 B.n190 585
R157 B.n189 B.n188 585
R158 B.n187 B.n186 585
R159 B.n185 B.n184 585
R160 B.n183 B.n182 585
R161 B.n181 B.n180 585
R162 B.n179 B.n178 585
R163 B.n177 B.n176 585
R164 B.n175 B.n174 585
R165 B.n173 B.n172 585
R166 B.n171 B.n170 585
R167 B.n169 B.n168 585
R168 B.n167 B.n166 585
R169 B.n165 B.n164 585
R170 B.n163 B.n162 585
R171 B.n161 B.n160 585
R172 B.n159 B.n158 585
R173 B.n157 B.n156 585
R174 B.n155 B.n154 585
R175 B.n153 B.n152 585
R176 B.n151 B.n150 585
R177 B.n149 B.n148 585
R178 B.n147 B.n146 585
R179 B.n145 B.n144 585
R180 B.n143 B.n142 585
R181 B.n141 B.n140 585
R182 B.n139 B.n138 585
R183 B.n137 B.n136 585
R184 B.n135 B.n134 585
R185 B.n133 B.n132 585
R186 B.n131 B.n130 585
R187 B.n129 B.n128 585
R188 B.n127 B.n126 585
R189 B.n125 B.n124 585
R190 B.n123 B.n122 585
R191 B.n121 B.n120 585
R192 B.n798 B.n63 585
R193 B.n803 B.n63 585
R194 B.n797 B.n62 585
R195 B.n804 B.n62 585
R196 B.n796 B.n795 585
R197 B.n795 B.n58 585
R198 B.n794 B.n57 585
R199 B.n810 B.n57 585
R200 B.n793 B.n56 585
R201 B.n811 B.n56 585
R202 B.n792 B.n55 585
R203 B.n812 B.n55 585
R204 B.n791 B.n790 585
R205 B.n790 B.n54 585
R206 B.n789 B.n50 585
R207 B.n818 B.n50 585
R208 B.n788 B.n49 585
R209 B.n819 B.n49 585
R210 B.n787 B.n48 585
R211 B.n820 B.n48 585
R212 B.n786 B.n785 585
R213 B.n785 B.n44 585
R214 B.n784 B.n43 585
R215 B.n826 B.n43 585
R216 B.n783 B.n42 585
R217 B.n827 B.n42 585
R218 B.n782 B.n41 585
R219 B.n828 B.n41 585
R220 B.n781 B.n780 585
R221 B.n780 B.n37 585
R222 B.n779 B.n36 585
R223 B.n834 B.n36 585
R224 B.n778 B.n35 585
R225 B.n835 B.n35 585
R226 B.n777 B.n34 585
R227 B.n836 B.n34 585
R228 B.n776 B.n775 585
R229 B.n775 B.n30 585
R230 B.n774 B.n29 585
R231 B.n842 B.n29 585
R232 B.n773 B.n28 585
R233 B.n843 B.n28 585
R234 B.n772 B.n27 585
R235 B.n844 B.n27 585
R236 B.n771 B.n770 585
R237 B.n770 B.n26 585
R238 B.n769 B.n22 585
R239 B.n850 B.n22 585
R240 B.n768 B.n21 585
R241 B.n851 B.n21 585
R242 B.n767 B.n20 585
R243 B.n852 B.n20 585
R244 B.n766 B.n765 585
R245 B.n765 B.n16 585
R246 B.n764 B.n15 585
R247 B.n858 B.n15 585
R248 B.n763 B.n14 585
R249 B.n859 B.n14 585
R250 B.n762 B.n13 585
R251 B.n860 B.n13 585
R252 B.n761 B.n760 585
R253 B.n760 B.n12 585
R254 B.n759 B.n758 585
R255 B.n759 B.n8 585
R256 B.n757 B.n7 585
R257 B.n867 B.n7 585
R258 B.n756 B.n6 585
R259 B.n868 B.n6 585
R260 B.n755 B.n5 585
R261 B.n869 B.n5 585
R262 B.n754 B.n753 585
R263 B.n753 B.n4 585
R264 B.n752 B.n327 585
R265 B.n752 B.n751 585
R266 B.n742 B.n328 585
R267 B.n329 B.n328 585
R268 B.n744 B.n743 585
R269 B.n745 B.n744 585
R270 B.n741 B.n333 585
R271 B.n337 B.n333 585
R272 B.n740 B.n739 585
R273 B.n739 B.n738 585
R274 B.n335 B.n334 585
R275 B.n336 B.n335 585
R276 B.n731 B.n730 585
R277 B.n732 B.n731 585
R278 B.n729 B.n342 585
R279 B.n342 B.n341 585
R280 B.n728 B.n727 585
R281 B.n727 B.n726 585
R282 B.n344 B.n343 585
R283 B.n719 B.n344 585
R284 B.n718 B.n717 585
R285 B.n720 B.n718 585
R286 B.n716 B.n349 585
R287 B.n349 B.n348 585
R288 B.n715 B.n714 585
R289 B.n714 B.n713 585
R290 B.n351 B.n350 585
R291 B.n352 B.n351 585
R292 B.n706 B.n705 585
R293 B.n707 B.n706 585
R294 B.n704 B.n356 585
R295 B.n360 B.n356 585
R296 B.n703 B.n702 585
R297 B.n702 B.n701 585
R298 B.n358 B.n357 585
R299 B.n359 B.n358 585
R300 B.n694 B.n693 585
R301 B.n695 B.n694 585
R302 B.n692 B.n365 585
R303 B.n365 B.n364 585
R304 B.n691 B.n690 585
R305 B.n690 B.n689 585
R306 B.n367 B.n366 585
R307 B.n368 B.n367 585
R308 B.n682 B.n681 585
R309 B.n683 B.n682 585
R310 B.n680 B.n373 585
R311 B.n373 B.n372 585
R312 B.n679 B.n678 585
R313 B.n678 B.n677 585
R314 B.n375 B.n374 585
R315 B.n670 B.n375 585
R316 B.n669 B.n668 585
R317 B.n671 B.n669 585
R318 B.n667 B.n380 585
R319 B.n380 B.n379 585
R320 B.n666 B.n665 585
R321 B.n665 B.n664 585
R322 B.n382 B.n381 585
R323 B.n383 B.n382 585
R324 B.n657 B.n656 585
R325 B.n658 B.n657 585
R326 B.n655 B.n388 585
R327 B.n388 B.n387 585
R328 B.n650 B.n649 585
R329 B.n648 B.n442 585
R330 B.n647 B.n441 585
R331 B.n652 B.n441 585
R332 B.n646 B.n645 585
R333 B.n644 B.n643 585
R334 B.n642 B.n641 585
R335 B.n640 B.n639 585
R336 B.n638 B.n637 585
R337 B.n636 B.n635 585
R338 B.n634 B.n633 585
R339 B.n632 B.n631 585
R340 B.n630 B.n629 585
R341 B.n628 B.n627 585
R342 B.n626 B.n625 585
R343 B.n624 B.n623 585
R344 B.n622 B.n621 585
R345 B.n620 B.n619 585
R346 B.n618 B.n617 585
R347 B.n616 B.n615 585
R348 B.n614 B.n613 585
R349 B.n612 B.n611 585
R350 B.n610 B.n609 585
R351 B.n608 B.n607 585
R352 B.n606 B.n605 585
R353 B.n604 B.n603 585
R354 B.n602 B.n601 585
R355 B.n600 B.n599 585
R356 B.n598 B.n597 585
R357 B.n596 B.n595 585
R358 B.n594 B.n593 585
R359 B.n592 B.n591 585
R360 B.n590 B.n589 585
R361 B.n588 B.n587 585
R362 B.n586 B.n585 585
R363 B.n584 B.n583 585
R364 B.n582 B.n581 585
R365 B.n580 B.n579 585
R366 B.n578 B.n577 585
R367 B.n576 B.n575 585
R368 B.n574 B.n573 585
R369 B.n572 B.n571 585
R370 B.n570 B.n569 585
R371 B.n568 B.n567 585
R372 B.n566 B.n565 585
R373 B.n564 B.n563 585
R374 B.n562 B.n561 585
R375 B.n560 B.n559 585
R376 B.n558 B.n557 585
R377 B.n556 B.n555 585
R378 B.n554 B.n553 585
R379 B.n552 B.n551 585
R380 B.n550 B.n549 585
R381 B.n548 B.n547 585
R382 B.n546 B.n545 585
R383 B.n544 B.n543 585
R384 B.n542 B.n541 585
R385 B.n540 B.n539 585
R386 B.n538 B.n537 585
R387 B.n536 B.n535 585
R388 B.n534 B.n533 585
R389 B.n532 B.n531 585
R390 B.n530 B.n529 585
R391 B.n528 B.n527 585
R392 B.n526 B.n525 585
R393 B.n524 B.n523 585
R394 B.n522 B.n521 585
R395 B.n520 B.n519 585
R396 B.n518 B.n517 585
R397 B.n516 B.n515 585
R398 B.n514 B.n513 585
R399 B.n512 B.n511 585
R400 B.n510 B.n509 585
R401 B.n508 B.n507 585
R402 B.n506 B.n505 585
R403 B.n504 B.n503 585
R404 B.n502 B.n501 585
R405 B.n500 B.n499 585
R406 B.n498 B.n497 585
R407 B.n496 B.n495 585
R408 B.n494 B.n493 585
R409 B.n492 B.n491 585
R410 B.n490 B.n489 585
R411 B.n488 B.n487 585
R412 B.n486 B.n485 585
R413 B.n484 B.n483 585
R414 B.n482 B.n481 585
R415 B.n480 B.n479 585
R416 B.n478 B.n477 585
R417 B.n476 B.n475 585
R418 B.n474 B.n473 585
R419 B.n472 B.n471 585
R420 B.n470 B.n469 585
R421 B.n468 B.n467 585
R422 B.n466 B.n465 585
R423 B.n464 B.n463 585
R424 B.n462 B.n461 585
R425 B.n460 B.n459 585
R426 B.n458 B.n457 585
R427 B.n456 B.n455 585
R428 B.n454 B.n453 585
R429 B.n452 B.n451 585
R430 B.n450 B.n449 585
R431 B.n390 B.n389 585
R432 B.n654 B.n653 585
R433 B.n653 B.n652 585
R434 B.n386 B.n385 585
R435 B.n387 B.n386 585
R436 B.n660 B.n659 585
R437 B.n659 B.n658 585
R438 B.n661 B.n384 585
R439 B.n384 B.n383 585
R440 B.n663 B.n662 585
R441 B.n664 B.n663 585
R442 B.n378 B.n377 585
R443 B.n379 B.n378 585
R444 B.n673 B.n672 585
R445 B.n672 B.n671 585
R446 B.n674 B.n376 585
R447 B.n670 B.n376 585
R448 B.n676 B.n675 585
R449 B.n677 B.n676 585
R450 B.n371 B.n370 585
R451 B.n372 B.n371 585
R452 B.n685 B.n684 585
R453 B.n684 B.n683 585
R454 B.n686 B.n369 585
R455 B.n369 B.n368 585
R456 B.n688 B.n687 585
R457 B.n689 B.n688 585
R458 B.n363 B.n362 585
R459 B.n364 B.n363 585
R460 B.n697 B.n696 585
R461 B.n696 B.n695 585
R462 B.n698 B.n361 585
R463 B.n361 B.n359 585
R464 B.n700 B.n699 585
R465 B.n701 B.n700 585
R466 B.n355 B.n354 585
R467 B.n360 B.n355 585
R468 B.n709 B.n708 585
R469 B.n708 B.n707 585
R470 B.n710 B.n353 585
R471 B.n353 B.n352 585
R472 B.n712 B.n711 585
R473 B.n713 B.n712 585
R474 B.n347 B.n346 585
R475 B.n348 B.n347 585
R476 B.n722 B.n721 585
R477 B.n721 B.n720 585
R478 B.n723 B.n345 585
R479 B.n719 B.n345 585
R480 B.n725 B.n724 585
R481 B.n726 B.n725 585
R482 B.n340 B.n339 585
R483 B.n341 B.n340 585
R484 B.n734 B.n733 585
R485 B.n733 B.n732 585
R486 B.n735 B.n338 585
R487 B.n338 B.n336 585
R488 B.n737 B.n736 585
R489 B.n738 B.n737 585
R490 B.n332 B.n331 585
R491 B.n337 B.n332 585
R492 B.n747 B.n746 585
R493 B.n746 B.n745 585
R494 B.n748 B.n330 585
R495 B.n330 B.n329 585
R496 B.n750 B.n749 585
R497 B.n751 B.n750 585
R498 B.n3 B.n0 585
R499 B.n4 B.n3 585
R500 B.n866 B.n1 585
R501 B.n867 B.n866 585
R502 B.n865 B.n864 585
R503 B.n865 B.n8 585
R504 B.n863 B.n9 585
R505 B.n12 B.n9 585
R506 B.n862 B.n861 585
R507 B.n861 B.n860 585
R508 B.n11 B.n10 585
R509 B.n859 B.n11 585
R510 B.n857 B.n856 585
R511 B.n858 B.n857 585
R512 B.n855 B.n17 585
R513 B.n17 B.n16 585
R514 B.n854 B.n853 585
R515 B.n853 B.n852 585
R516 B.n19 B.n18 585
R517 B.n851 B.n19 585
R518 B.n849 B.n848 585
R519 B.n850 B.n849 585
R520 B.n847 B.n23 585
R521 B.n26 B.n23 585
R522 B.n846 B.n845 585
R523 B.n845 B.n844 585
R524 B.n25 B.n24 585
R525 B.n843 B.n25 585
R526 B.n841 B.n840 585
R527 B.n842 B.n841 585
R528 B.n839 B.n31 585
R529 B.n31 B.n30 585
R530 B.n838 B.n837 585
R531 B.n837 B.n836 585
R532 B.n33 B.n32 585
R533 B.n835 B.n33 585
R534 B.n833 B.n832 585
R535 B.n834 B.n833 585
R536 B.n831 B.n38 585
R537 B.n38 B.n37 585
R538 B.n830 B.n829 585
R539 B.n829 B.n828 585
R540 B.n40 B.n39 585
R541 B.n827 B.n40 585
R542 B.n825 B.n824 585
R543 B.n826 B.n825 585
R544 B.n823 B.n45 585
R545 B.n45 B.n44 585
R546 B.n822 B.n821 585
R547 B.n821 B.n820 585
R548 B.n47 B.n46 585
R549 B.n819 B.n47 585
R550 B.n817 B.n816 585
R551 B.n818 B.n817 585
R552 B.n815 B.n51 585
R553 B.n54 B.n51 585
R554 B.n814 B.n813 585
R555 B.n813 B.n812 585
R556 B.n53 B.n52 585
R557 B.n811 B.n53 585
R558 B.n809 B.n808 585
R559 B.n810 B.n809 585
R560 B.n807 B.n59 585
R561 B.n59 B.n58 585
R562 B.n806 B.n805 585
R563 B.n805 B.n804 585
R564 B.n61 B.n60 585
R565 B.n803 B.n61 585
R566 B.n870 B.n869 585
R567 B.n868 B.n2 585
R568 B.n120 B.n61 482.89
R569 B.n800 B.n63 482.89
R570 B.n653 B.n388 482.89
R571 B.n650 B.n386 482.89
R572 B.n118 B.t9 390.522
R573 B.n116 B.t5 390.522
R574 B.n446 B.t16 390.522
R575 B.n443 B.t12 390.522
R576 B.n802 B.n801 256.663
R577 B.n802 B.n114 256.663
R578 B.n802 B.n113 256.663
R579 B.n802 B.n112 256.663
R580 B.n802 B.n111 256.663
R581 B.n802 B.n110 256.663
R582 B.n802 B.n109 256.663
R583 B.n802 B.n108 256.663
R584 B.n802 B.n107 256.663
R585 B.n802 B.n106 256.663
R586 B.n802 B.n105 256.663
R587 B.n802 B.n104 256.663
R588 B.n802 B.n103 256.663
R589 B.n802 B.n102 256.663
R590 B.n802 B.n101 256.663
R591 B.n802 B.n100 256.663
R592 B.n802 B.n99 256.663
R593 B.n802 B.n98 256.663
R594 B.n802 B.n97 256.663
R595 B.n802 B.n96 256.663
R596 B.n802 B.n95 256.663
R597 B.n802 B.n94 256.663
R598 B.n802 B.n93 256.663
R599 B.n802 B.n92 256.663
R600 B.n802 B.n91 256.663
R601 B.n802 B.n90 256.663
R602 B.n802 B.n89 256.663
R603 B.n802 B.n88 256.663
R604 B.n802 B.n87 256.663
R605 B.n802 B.n86 256.663
R606 B.n802 B.n85 256.663
R607 B.n802 B.n84 256.663
R608 B.n802 B.n83 256.663
R609 B.n802 B.n82 256.663
R610 B.n802 B.n81 256.663
R611 B.n802 B.n80 256.663
R612 B.n802 B.n79 256.663
R613 B.n802 B.n78 256.663
R614 B.n802 B.n77 256.663
R615 B.n802 B.n76 256.663
R616 B.n802 B.n75 256.663
R617 B.n802 B.n74 256.663
R618 B.n802 B.n73 256.663
R619 B.n802 B.n72 256.663
R620 B.n802 B.n71 256.663
R621 B.n802 B.n70 256.663
R622 B.n802 B.n69 256.663
R623 B.n802 B.n68 256.663
R624 B.n802 B.n67 256.663
R625 B.n802 B.n66 256.663
R626 B.n802 B.n65 256.663
R627 B.n802 B.n64 256.663
R628 B.n652 B.n651 256.663
R629 B.n652 B.n391 256.663
R630 B.n652 B.n392 256.663
R631 B.n652 B.n393 256.663
R632 B.n652 B.n394 256.663
R633 B.n652 B.n395 256.663
R634 B.n652 B.n396 256.663
R635 B.n652 B.n397 256.663
R636 B.n652 B.n398 256.663
R637 B.n652 B.n399 256.663
R638 B.n652 B.n400 256.663
R639 B.n652 B.n401 256.663
R640 B.n652 B.n402 256.663
R641 B.n652 B.n403 256.663
R642 B.n652 B.n404 256.663
R643 B.n652 B.n405 256.663
R644 B.n652 B.n406 256.663
R645 B.n652 B.n407 256.663
R646 B.n652 B.n408 256.663
R647 B.n652 B.n409 256.663
R648 B.n652 B.n410 256.663
R649 B.n652 B.n411 256.663
R650 B.n652 B.n412 256.663
R651 B.n652 B.n413 256.663
R652 B.n652 B.n414 256.663
R653 B.n652 B.n415 256.663
R654 B.n652 B.n416 256.663
R655 B.n652 B.n417 256.663
R656 B.n652 B.n418 256.663
R657 B.n652 B.n419 256.663
R658 B.n652 B.n420 256.663
R659 B.n652 B.n421 256.663
R660 B.n652 B.n422 256.663
R661 B.n652 B.n423 256.663
R662 B.n652 B.n424 256.663
R663 B.n652 B.n425 256.663
R664 B.n652 B.n426 256.663
R665 B.n652 B.n427 256.663
R666 B.n652 B.n428 256.663
R667 B.n652 B.n429 256.663
R668 B.n652 B.n430 256.663
R669 B.n652 B.n431 256.663
R670 B.n652 B.n432 256.663
R671 B.n652 B.n433 256.663
R672 B.n652 B.n434 256.663
R673 B.n652 B.n435 256.663
R674 B.n652 B.n436 256.663
R675 B.n652 B.n437 256.663
R676 B.n652 B.n438 256.663
R677 B.n652 B.n439 256.663
R678 B.n652 B.n440 256.663
R679 B.n872 B.n871 256.663
R680 B.n124 B.n123 163.367
R681 B.n128 B.n127 163.367
R682 B.n132 B.n131 163.367
R683 B.n136 B.n135 163.367
R684 B.n140 B.n139 163.367
R685 B.n144 B.n143 163.367
R686 B.n148 B.n147 163.367
R687 B.n152 B.n151 163.367
R688 B.n156 B.n155 163.367
R689 B.n160 B.n159 163.367
R690 B.n164 B.n163 163.367
R691 B.n168 B.n167 163.367
R692 B.n172 B.n171 163.367
R693 B.n176 B.n175 163.367
R694 B.n180 B.n179 163.367
R695 B.n184 B.n183 163.367
R696 B.n188 B.n187 163.367
R697 B.n192 B.n191 163.367
R698 B.n196 B.n195 163.367
R699 B.n200 B.n199 163.367
R700 B.n204 B.n203 163.367
R701 B.n208 B.n207 163.367
R702 B.n212 B.n211 163.367
R703 B.n217 B.n216 163.367
R704 B.n221 B.n220 163.367
R705 B.n225 B.n224 163.367
R706 B.n229 B.n228 163.367
R707 B.n233 B.n232 163.367
R708 B.n238 B.n237 163.367
R709 B.n242 B.n241 163.367
R710 B.n246 B.n245 163.367
R711 B.n250 B.n249 163.367
R712 B.n254 B.n253 163.367
R713 B.n258 B.n257 163.367
R714 B.n262 B.n261 163.367
R715 B.n266 B.n265 163.367
R716 B.n270 B.n269 163.367
R717 B.n274 B.n273 163.367
R718 B.n278 B.n277 163.367
R719 B.n282 B.n281 163.367
R720 B.n286 B.n285 163.367
R721 B.n290 B.n289 163.367
R722 B.n294 B.n293 163.367
R723 B.n298 B.n297 163.367
R724 B.n302 B.n301 163.367
R725 B.n306 B.n305 163.367
R726 B.n310 B.n309 163.367
R727 B.n314 B.n313 163.367
R728 B.n318 B.n317 163.367
R729 B.n322 B.n321 163.367
R730 B.n324 B.n115 163.367
R731 B.n657 B.n388 163.367
R732 B.n657 B.n382 163.367
R733 B.n665 B.n382 163.367
R734 B.n665 B.n380 163.367
R735 B.n669 B.n380 163.367
R736 B.n669 B.n375 163.367
R737 B.n678 B.n375 163.367
R738 B.n678 B.n373 163.367
R739 B.n682 B.n373 163.367
R740 B.n682 B.n367 163.367
R741 B.n690 B.n367 163.367
R742 B.n690 B.n365 163.367
R743 B.n694 B.n365 163.367
R744 B.n694 B.n358 163.367
R745 B.n702 B.n358 163.367
R746 B.n702 B.n356 163.367
R747 B.n706 B.n356 163.367
R748 B.n706 B.n351 163.367
R749 B.n714 B.n351 163.367
R750 B.n714 B.n349 163.367
R751 B.n718 B.n349 163.367
R752 B.n718 B.n344 163.367
R753 B.n727 B.n344 163.367
R754 B.n727 B.n342 163.367
R755 B.n731 B.n342 163.367
R756 B.n731 B.n335 163.367
R757 B.n739 B.n335 163.367
R758 B.n739 B.n333 163.367
R759 B.n744 B.n333 163.367
R760 B.n744 B.n328 163.367
R761 B.n752 B.n328 163.367
R762 B.n753 B.n752 163.367
R763 B.n753 B.n5 163.367
R764 B.n6 B.n5 163.367
R765 B.n7 B.n6 163.367
R766 B.n759 B.n7 163.367
R767 B.n760 B.n759 163.367
R768 B.n760 B.n13 163.367
R769 B.n14 B.n13 163.367
R770 B.n15 B.n14 163.367
R771 B.n765 B.n15 163.367
R772 B.n765 B.n20 163.367
R773 B.n21 B.n20 163.367
R774 B.n22 B.n21 163.367
R775 B.n770 B.n22 163.367
R776 B.n770 B.n27 163.367
R777 B.n28 B.n27 163.367
R778 B.n29 B.n28 163.367
R779 B.n775 B.n29 163.367
R780 B.n775 B.n34 163.367
R781 B.n35 B.n34 163.367
R782 B.n36 B.n35 163.367
R783 B.n780 B.n36 163.367
R784 B.n780 B.n41 163.367
R785 B.n42 B.n41 163.367
R786 B.n43 B.n42 163.367
R787 B.n785 B.n43 163.367
R788 B.n785 B.n48 163.367
R789 B.n49 B.n48 163.367
R790 B.n50 B.n49 163.367
R791 B.n790 B.n50 163.367
R792 B.n790 B.n55 163.367
R793 B.n56 B.n55 163.367
R794 B.n57 B.n56 163.367
R795 B.n795 B.n57 163.367
R796 B.n795 B.n62 163.367
R797 B.n63 B.n62 163.367
R798 B.n442 B.n441 163.367
R799 B.n645 B.n441 163.367
R800 B.n643 B.n642 163.367
R801 B.n639 B.n638 163.367
R802 B.n635 B.n634 163.367
R803 B.n631 B.n630 163.367
R804 B.n627 B.n626 163.367
R805 B.n623 B.n622 163.367
R806 B.n619 B.n618 163.367
R807 B.n615 B.n614 163.367
R808 B.n611 B.n610 163.367
R809 B.n607 B.n606 163.367
R810 B.n603 B.n602 163.367
R811 B.n599 B.n598 163.367
R812 B.n595 B.n594 163.367
R813 B.n591 B.n590 163.367
R814 B.n587 B.n586 163.367
R815 B.n583 B.n582 163.367
R816 B.n579 B.n578 163.367
R817 B.n575 B.n574 163.367
R818 B.n571 B.n570 163.367
R819 B.n567 B.n566 163.367
R820 B.n563 B.n562 163.367
R821 B.n559 B.n558 163.367
R822 B.n555 B.n554 163.367
R823 B.n551 B.n550 163.367
R824 B.n547 B.n546 163.367
R825 B.n543 B.n542 163.367
R826 B.n539 B.n538 163.367
R827 B.n535 B.n534 163.367
R828 B.n531 B.n530 163.367
R829 B.n527 B.n526 163.367
R830 B.n523 B.n522 163.367
R831 B.n519 B.n518 163.367
R832 B.n515 B.n514 163.367
R833 B.n511 B.n510 163.367
R834 B.n507 B.n506 163.367
R835 B.n503 B.n502 163.367
R836 B.n499 B.n498 163.367
R837 B.n495 B.n494 163.367
R838 B.n491 B.n490 163.367
R839 B.n487 B.n486 163.367
R840 B.n483 B.n482 163.367
R841 B.n479 B.n478 163.367
R842 B.n475 B.n474 163.367
R843 B.n471 B.n470 163.367
R844 B.n467 B.n466 163.367
R845 B.n463 B.n462 163.367
R846 B.n459 B.n458 163.367
R847 B.n455 B.n454 163.367
R848 B.n451 B.n450 163.367
R849 B.n653 B.n390 163.367
R850 B.n659 B.n386 163.367
R851 B.n659 B.n384 163.367
R852 B.n663 B.n384 163.367
R853 B.n663 B.n378 163.367
R854 B.n672 B.n378 163.367
R855 B.n672 B.n376 163.367
R856 B.n676 B.n376 163.367
R857 B.n676 B.n371 163.367
R858 B.n684 B.n371 163.367
R859 B.n684 B.n369 163.367
R860 B.n688 B.n369 163.367
R861 B.n688 B.n363 163.367
R862 B.n696 B.n363 163.367
R863 B.n696 B.n361 163.367
R864 B.n700 B.n361 163.367
R865 B.n700 B.n355 163.367
R866 B.n708 B.n355 163.367
R867 B.n708 B.n353 163.367
R868 B.n712 B.n353 163.367
R869 B.n712 B.n347 163.367
R870 B.n721 B.n347 163.367
R871 B.n721 B.n345 163.367
R872 B.n725 B.n345 163.367
R873 B.n725 B.n340 163.367
R874 B.n733 B.n340 163.367
R875 B.n733 B.n338 163.367
R876 B.n737 B.n338 163.367
R877 B.n737 B.n332 163.367
R878 B.n746 B.n332 163.367
R879 B.n746 B.n330 163.367
R880 B.n750 B.n330 163.367
R881 B.n750 B.n3 163.367
R882 B.n870 B.n3 163.367
R883 B.n866 B.n2 163.367
R884 B.n866 B.n865 163.367
R885 B.n865 B.n9 163.367
R886 B.n861 B.n9 163.367
R887 B.n861 B.n11 163.367
R888 B.n857 B.n11 163.367
R889 B.n857 B.n17 163.367
R890 B.n853 B.n17 163.367
R891 B.n853 B.n19 163.367
R892 B.n849 B.n19 163.367
R893 B.n849 B.n23 163.367
R894 B.n845 B.n23 163.367
R895 B.n845 B.n25 163.367
R896 B.n841 B.n25 163.367
R897 B.n841 B.n31 163.367
R898 B.n837 B.n31 163.367
R899 B.n837 B.n33 163.367
R900 B.n833 B.n33 163.367
R901 B.n833 B.n38 163.367
R902 B.n829 B.n38 163.367
R903 B.n829 B.n40 163.367
R904 B.n825 B.n40 163.367
R905 B.n825 B.n45 163.367
R906 B.n821 B.n45 163.367
R907 B.n821 B.n47 163.367
R908 B.n817 B.n47 163.367
R909 B.n817 B.n51 163.367
R910 B.n813 B.n51 163.367
R911 B.n813 B.n53 163.367
R912 B.n809 B.n53 163.367
R913 B.n809 B.n59 163.367
R914 B.n805 B.n59 163.367
R915 B.n805 B.n61 163.367
R916 B.n116 B.t7 115.082
R917 B.n446 B.t18 115.082
R918 B.n118 B.t10 115.064
R919 B.n443 B.t15 115.064
R920 B.n117 B.t8 73.385
R921 B.n447 B.t17 73.385
R922 B.n119 B.t11 73.3673
R923 B.n444 B.t14 73.3673
R924 B.n120 B.n64 71.676
R925 B.n124 B.n65 71.676
R926 B.n128 B.n66 71.676
R927 B.n132 B.n67 71.676
R928 B.n136 B.n68 71.676
R929 B.n140 B.n69 71.676
R930 B.n144 B.n70 71.676
R931 B.n148 B.n71 71.676
R932 B.n152 B.n72 71.676
R933 B.n156 B.n73 71.676
R934 B.n160 B.n74 71.676
R935 B.n164 B.n75 71.676
R936 B.n168 B.n76 71.676
R937 B.n172 B.n77 71.676
R938 B.n176 B.n78 71.676
R939 B.n180 B.n79 71.676
R940 B.n184 B.n80 71.676
R941 B.n188 B.n81 71.676
R942 B.n192 B.n82 71.676
R943 B.n196 B.n83 71.676
R944 B.n200 B.n84 71.676
R945 B.n204 B.n85 71.676
R946 B.n208 B.n86 71.676
R947 B.n212 B.n87 71.676
R948 B.n217 B.n88 71.676
R949 B.n221 B.n89 71.676
R950 B.n225 B.n90 71.676
R951 B.n229 B.n91 71.676
R952 B.n233 B.n92 71.676
R953 B.n238 B.n93 71.676
R954 B.n242 B.n94 71.676
R955 B.n246 B.n95 71.676
R956 B.n250 B.n96 71.676
R957 B.n254 B.n97 71.676
R958 B.n258 B.n98 71.676
R959 B.n262 B.n99 71.676
R960 B.n266 B.n100 71.676
R961 B.n270 B.n101 71.676
R962 B.n274 B.n102 71.676
R963 B.n278 B.n103 71.676
R964 B.n282 B.n104 71.676
R965 B.n286 B.n105 71.676
R966 B.n290 B.n106 71.676
R967 B.n294 B.n107 71.676
R968 B.n298 B.n108 71.676
R969 B.n302 B.n109 71.676
R970 B.n306 B.n110 71.676
R971 B.n310 B.n111 71.676
R972 B.n314 B.n112 71.676
R973 B.n318 B.n113 71.676
R974 B.n322 B.n114 71.676
R975 B.n801 B.n115 71.676
R976 B.n801 B.n800 71.676
R977 B.n324 B.n114 71.676
R978 B.n321 B.n113 71.676
R979 B.n317 B.n112 71.676
R980 B.n313 B.n111 71.676
R981 B.n309 B.n110 71.676
R982 B.n305 B.n109 71.676
R983 B.n301 B.n108 71.676
R984 B.n297 B.n107 71.676
R985 B.n293 B.n106 71.676
R986 B.n289 B.n105 71.676
R987 B.n285 B.n104 71.676
R988 B.n281 B.n103 71.676
R989 B.n277 B.n102 71.676
R990 B.n273 B.n101 71.676
R991 B.n269 B.n100 71.676
R992 B.n265 B.n99 71.676
R993 B.n261 B.n98 71.676
R994 B.n257 B.n97 71.676
R995 B.n253 B.n96 71.676
R996 B.n249 B.n95 71.676
R997 B.n245 B.n94 71.676
R998 B.n241 B.n93 71.676
R999 B.n237 B.n92 71.676
R1000 B.n232 B.n91 71.676
R1001 B.n228 B.n90 71.676
R1002 B.n224 B.n89 71.676
R1003 B.n220 B.n88 71.676
R1004 B.n216 B.n87 71.676
R1005 B.n211 B.n86 71.676
R1006 B.n207 B.n85 71.676
R1007 B.n203 B.n84 71.676
R1008 B.n199 B.n83 71.676
R1009 B.n195 B.n82 71.676
R1010 B.n191 B.n81 71.676
R1011 B.n187 B.n80 71.676
R1012 B.n183 B.n79 71.676
R1013 B.n179 B.n78 71.676
R1014 B.n175 B.n77 71.676
R1015 B.n171 B.n76 71.676
R1016 B.n167 B.n75 71.676
R1017 B.n163 B.n74 71.676
R1018 B.n159 B.n73 71.676
R1019 B.n155 B.n72 71.676
R1020 B.n151 B.n71 71.676
R1021 B.n147 B.n70 71.676
R1022 B.n143 B.n69 71.676
R1023 B.n139 B.n68 71.676
R1024 B.n135 B.n67 71.676
R1025 B.n131 B.n66 71.676
R1026 B.n127 B.n65 71.676
R1027 B.n123 B.n64 71.676
R1028 B.n651 B.n650 71.676
R1029 B.n645 B.n391 71.676
R1030 B.n642 B.n392 71.676
R1031 B.n638 B.n393 71.676
R1032 B.n634 B.n394 71.676
R1033 B.n630 B.n395 71.676
R1034 B.n626 B.n396 71.676
R1035 B.n622 B.n397 71.676
R1036 B.n618 B.n398 71.676
R1037 B.n614 B.n399 71.676
R1038 B.n610 B.n400 71.676
R1039 B.n606 B.n401 71.676
R1040 B.n602 B.n402 71.676
R1041 B.n598 B.n403 71.676
R1042 B.n594 B.n404 71.676
R1043 B.n590 B.n405 71.676
R1044 B.n586 B.n406 71.676
R1045 B.n582 B.n407 71.676
R1046 B.n578 B.n408 71.676
R1047 B.n574 B.n409 71.676
R1048 B.n570 B.n410 71.676
R1049 B.n566 B.n411 71.676
R1050 B.n562 B.n412 71.676
R1051 B.n558 B.n413 71.676
R1052 B.n554 B.n414 71.676
R1053 B.n550 B.n415 71.676
R1054 B.n546 B.n416 71.676
R1055 B.n542 B.n417 71.676
R1056 B.n538 B.n418 71.676
R1057 B.n534 B.n419 71.676
R1058 B.n530 B.n420 71.676
R1059 B.n526 B.n421 71.676
R1060 B.n522 B.n422 71.676
R1061 B.n518 B.n423 71.676
R1062 B.n514 B.n424 71.676
R1063 B.n510 B.n425 71.676
R1064 B.n506 B.n426 71.676
R1065 B.n502 B.n427 71.676
R1066 B.n498 B.n428 71.676
R1067 B.n494 B.n429 71.676
R1068 B.n490 B.n430 71.676
R1069 B.n486 B.n431 71.676
R1070 B.n482 B.n432 71.676
R1071 B.n478 B.n433 71.676
R1072 B.n474 B.n434 71.676
R1073 B.n470 B.n435 71.676
R1074 B.n466 B.n436 71.676
R1075 B.n462 B.n437 71.676
R1076 B.n458 B.n438 71.676
R1077 B.n454 B.n439 71.676
R1078 B.n450 B.n440 71.676
R1079 B.n651 B.n442 71.676
R1080 B.n643 B.n391 71.676
R1081 B.n639 B.n392 71.676
R1082 B.n635 B.n393 71.676
R1083 B.n631 B.n394 71.676
R1084 B.n627 B.n395 71.676
R1085 B.n623 B.n396 71.676
R1086 B.n619 B.n397 71.676
R1087 B.n615 B.n398 71.676
R1088 B.n611 B.n399 71.676
R1089 B.n607 B.n400 71.676
R1090 B.n603 B.n401 71.676
R1091 B.n599 B.n402 71.676
R1092 B.n595 B.n403 71.676
R1093 B.n591 B.n404 71.676
R1094 B.n587 B.n405 71.676
R1095 B.n583 B.n406 71.676
R1096 B.n579 B.n407 71.676
R1097 B.n575 B.n408 71.676
R1098 B.n571 B.n409 71.676
R1099 B.n567 B.n410 71.676
R1100 B.n563 B.n411 71.676
R1101 B.n559 B.n412 71.676
R1102 B.n555 B.n413 71.676
R1103 B.n551 B.n414 71.676
R1104 B.n547 B.n415 71.676
R1105 B.n543 B.n416 71.676
R1106 B.n539 B.n417 71.676
R1107 B.n535 B.n418 71.676
R1108 B.n531 B.n419 71.676
R1109 B.n527 B.n420 71.676
R1110 B.n523 B.n421 71.676
R1111 B.n519 B.n422 71.676
R1112 B.n515 B.n423 71.676
R1113 B.n511 B.n424 71.676
R1114 B.n507 B.n425 71.676
R1115 B.n503 B.n426 71.676
R1116 B.n499 B.n427 71.676
R1117 B.n495 B.n428 71.676
R1118 B.n491 B.n429 71.676
R1119 B.n487 B.n430 71.676
R1120 B.n483 B.n431 71.676
R1121 B.n479 B.n432 71.676
R1122 B.n475 B.n433 71.676
R1123 B.n471 B.n434 71.676
R1124 B.n467 B.n435 71.676
R1125 B.n463 B.n436 71.676
R1126 B.n459 B.n437 71.676
R1127 B.n455 B.n438 71.676
R1128 B.n451 B.n439 71.676
R1129 B.n440 B.n390 71.676
R1130 B.n871 B.n870 71.676
R1131 B.n871 B.n2 71.676
R1132 B.n652 B.n387 67.1191
R1133 B.n803 B.n802 67.1191
R1134 B.n214 B.n119 59.5399
R1135 B.n235 B.n117 59.5399
R1136 B.n448 B.n447 59.5399
R1137 B.n445 B.n444 59.5399
R1138 B.n119 B.n118 41.6975
R1139 B.n117 B.n116 41.6975
R1140 B.n447 B.n446 41.6975
R1141 B.n444 B.n443 41.6975
R1142 B.n658 B.n387 39.0096
R1143 B.n658 B.n383 39.0096
R1144 B.n664 B.n383 39.0096
R1145 B.n664 B.n379 39.0096
R1146 B.n671 B.n379 39.0096
R1147 B.n671 B.n670 39.0096
R1148 B.n677 B.n372 39.0096
R1149 B.n683 B.n372 39.0096
R1150 B.n683 B.n368 39.0096
R1151 B.n689 B.n368 39.0096
R1152 B.n689 B.n364 39.0096
R1153 B.n695 B.n364 39.0096
R1154 B.n695 B.n359 39.0096
R1155 B.n701 B.n359 39.0096
R1156 B.n701 B.n360 39.0096
R1157 B.n707 B.n352 39.0096
R1158 B.n713 B.n352 39.0096
R1159 B.n713 B.n348 39.0096
R1160 B.n720 B.n348 39.0096
R1161 B.n720 B.n719 39.0096
R1162 B.n726 B.n341 39.0096
R1163 B.n732 B.n341 39.0096
R1164 B.n732 B.n336 39.0096
R1165 B.n738 B.n336 39.0096
R1166 B.n738 B.n337 39.0096
R1167 B.n745 B.n329 39.0096
R1168 B.n751 B.n329 39.0096
R1169 B.n751 B.n4 39.0096
R1170 B.n869 B.n4 39.0096
R1171 B.n869 B.n868 39.0096
R1172 B.n868 B.n867 39.0096
R1173 B.n867 B.n8 39.0096
R1174 B.n12 B.n8 39.0096
R1175 B.n860 B.n12 39.0096
R1176 B.n859 B.n858 39.0096
R1177 B.n858 B.n16 39.0096
R1178 B.n852 B.n16 39.0096
R1179 B.n852 B.n851 39.0096
R1180 B.n851 B.n850 39.0096
R1181 B.n844 B.n26 39.0096
R1182 B.n844 B.n843 39.0096
R1183 B.n843 B.n842 39.0096
R1184 B.n842 B.n30 39.0096
R1185 B.n836 B.n30 39.0096
R1186 B.n835 B.n834 39.0096
R1187 B.n834 B.n37 39.0096
R1188 B.n828 B.n37 39.0096
R1189 B.n828 B.n827 39.0096
R1190 B.n827 B.n826 39.0096
R1191 B.n826 B.n44 39.0096
R1192 B.n820 B.n44 39.0096
R1193 B.n820 B.n819 39.0096
R1194 B.n819 B.n818 39.0096
R1195 B.n812 B.n54 39.0096
R1196 B.n812 B.n811 39.0096
R1197 B.n811 B.n810 39.0096
R1198 B.n810 B.n58 39.0096
R1199 B.n804 B.n58 39.0096
R1200 B.n804 B.n803 39.0096
R1201 B.n707 B.t4 35.5676
R1202 B.n836 B.t2 35.5676
R1203 B.n649 B.n385 31.3761
R1204 B.n655 B.n654 31.3761
R1205 B.n799 B.n798 31.3761
R1206 B.n121 B.n60 31.3761
R1207 B.n337 B.t19 28.6837
R1208 B.t1 B.n859 28.6837
R1209 B.n726 B.t3 22.947
R1210 B.n850 B.t0 22.947
R1211 B.n670 B.t13 21.7997
R1212 B.n54 B.t6 21.7997
R1213 B B.n872 18.0485
R1214 B.n677 B.t13 17.2104
R1215 B.n818 B.t6 17.2104
R1216 B.n719 B.t3 16.0631
R1217 B.n26 B.t0 16.0631
R1218 B.n660 B.n385 10.6151
R1219 B.n661 B.n660 10.6151
R1220 B.n662 B.n661 10.6151
R1221 B.n662 B.n377 10.6151
R1222 B.n673 B.n377 10.6151
R1223 B.n674 B.n673 10.6151
R1224 B.n675 B.n674 10.6151
R1225 B.n675 B.n370 10.6151
R1226 B.n685 B.n370 10.6151
R1227 B.n686 B.n685 10.6151
R1228 B.n687 B.n686 10.6151
R1229 B.n687 B.n362 10.6151
R1230 B.n697 B.n362 10.6151
R1231 B.n698 B.n697 10.6151
R1232 B.n699 B.n698 10.6151
R1233 B.n699 B.n354 10.6151
R1234 B.n709 B.n354 10.6151
R1235 B.n710 B.n709 10.6151
R1236 B.n711 B.n710 10.6151
R1237 B.n711 B.n346 10.6151
R1238 B.n722 B.n346 10.6151
R1239 B.n723 B.n722 10.6151
R1240 B.n724 B.n723 10.6151
R1241 B.n724 B.n339 10.6151
R1242 B.n734 B.n339 10.6151
R1243 B.n735 B.n734 10.6151
R1244 B.n736 B.n735 10.6151
R1245 B.n736 B.n331 10.6151
R1246 B.n747 B.n331 10.6151
R1247 B.n748 B.n747 10.6151
R1248 B.n749 B.n748 10.6151
R1249 B.n749 B.n0 10.6151
R1250 B.n649 B.n648 10.6151
R1251 B.n648 B.n647 10.6151
R1252 B.n647 B.n646 10.6151
R1253 B.n646 B.n644 10.6151
R1254 B.n644 B.n641 10.6151
R1255 B.n641 B.n640 10.6151
R1256 B.n640 B.n637 10.6151
R1257 B.n637 B.n636 10.6151
R1258 B.n636 B.n633 10.6151
R1259 B.n633 B.n632 10.6151
R1260 B.n632 B.n629 10.6151
R1261 B.n629 B.n628 10.6151
R1262 B.n628 B.n625 10.6151
R1263 B.n625 B.n624 10.6151
R1264 B.n624 B.n621 10.6151
R1265 B.n621 B.n620 10.6151
R1266 B.n620 B.n617 10.6151
R1267 B.n617 B.n616 10.6151
R1268 B.n616 B.n613 10.6151
R1269 B.n613 B.n612 10.6151
R1270 B.n612 B.n609 10.6151
R1271 B.n609 B.n608 10.6151
R1272 B.n608 B.n605 10.6151
R1273 B.n605 B.n604 10.6151
R1274 B.n604 B.n601 10.6151
R1275 B.n601 B.n600 10.6151
R1276 B.n600 B.n597 10.6151
R1277 B.n597 B.n596 10.6151
R1278 B.n596 B.n593 10.6151
R1279 B.n593 B.n592 10.6151
R1280 B.n592 B.n589 10.6151
R1281 B.n589 B.n588 10.6151
R1282 B.n588 B.n585 10.6151
R1283 B.n585 B.n584 10.6151
R1284 B.n584 B.n581 10.6151
R1285 B.n581 B.n580 10.6151
R1286 B.n580 B.n577 10.6151
R1287 B.n577 B.n576 10.6151
R1288 B.n576 B.n573 10.6151
R1289 B.n573 B.n572 10.6151
R1290 B.n572 B.n569 10.6151
R1291 B.n569 B.n568 10.6151
R1292 B.n568 B.n565 10.6151
R1293 B.n565 B.n564 10.6151
R1294 B.n564 B.n561 10.6151
R1295 B.n561 B.n560 10.6151
R1296 B.n557 B.n556 10.6151
R1297 B.n556 B.n553 10.6151
R1298 B.n553 B.n552 10.6151
R1299 B.n552 B.n549 10.6151
R1300 B.n549 B.n548 10.6151
R1301 B.n548 B.n545 10.6151
R1302 B.n545 B.n544 10.6151
R1303 B.n544 B.n541 10.6151
R1304 B.n541 B.n540 10.6151
R1305 B.n537 B.n536 10.6151
R1306 B.n536 B.n533 10.6151
R1307 B.n533 B.n532 10.6151
R1308 B.n532 B.n529 10.6151
R1309 B.n529 B.n528 10.6151
R1310 B.n528 B.n525 10.6151
R1311 B.n525 B.n524 10.6151
R1312 B.n524 B.n521 10.6151
R1313 B.n521 B.n520 10.6151
R1314 B.n520 B.n517 10.6151
R1315 B.n517 B.n516 10.6151
R1316 B.n516 B.n513 10.6151
R1317 B.n513 B.n512 10.6151
R1318 B.n512 B.n509 10.6151
R1319 B.n509 B.n508 10.6151
R1320 B.n508 B.n505 10.6151
R1321 B.n505 B.n504 10.6151
R1322 B.n504 B.n501 10.6151
R1323 B.n501 B.n500 10.6151
R1324 B.n500 B.n497 10.6151
R1325 B.n497 B.n496 10.6151
R1326 B.n496 B.n493 10.6151
R1327 B.n493 B.n492 10.6151
R1328 B.n492 B.n489 10.6151
R1329 B.n489 B.n488 10.6151
R1330 B.n488 B.n485 10.6151
R1331 B.n485 B.n484 10.6151
R1332 B.n484 B.n481 10.6151
R1333 B.n481 B.n480 10.6151
R1334 B.n480 B.n477 10.6151
R1335 B.n477 B.n476 10.6151
R1336 B.n476 B.n473 10.6151
R1337 B.n473 B.n472 10.6151
R1338 B.n472 B.n469 10.6151
R1339 B.n469 B.n468 10.6151
R1340 B.n468 B.n465 10.6151
R1341 B.n465 B.n464 10.6151
R1342 B.n464 B.n461 10.6151
R1343 B.n461 B.n460 10.6151
R1344 B.n460 B.n457 10.6151
R1345 B.n457 B.n456 10.6151
R1346 B.n456 B.n453 10.6151
R1347 B.n453 B.n452 10.6151
R1348 B.n452 B.n449 10.6151
R1349 B.n449 B.n389 10.6151
R1350 B.n654 B.n389 10.6151
R1351 B.n656 B.n655 10.6151
R1352 B.n656 B.n381 10.6151
R1353 B.n666 B.n381 10.6151
R1354 B.n667 B.n666 10.6151
R1355 B.n668 B.n667 10.6151
R1356 B.n668 B.n374 10.6151
R1357 B.n679 B.n374 10.6151
R1358 B.n680 B.n679 10.6151
R1359 B.n681 B.n680 10.6151
R1360 B.n681 B.n366 10.6151
R1361 B.n691 B.n366 10.6151
R1362 B.n692 B.n691 10.6151
R1363 B.n693 B.n692 10.6151
R1364 B.n693 B.n357 10.6151
R1365 B.n703 B.n357 10.6151
R1366 B.n704 B.n703 10.6151
R1367 B.n705 B.n704 10.6151
R1368 B.n705 B.n350 10.6151
R1369 B.n715 B.n350 10.6151
R1370 B.n716 B.n715 10.6151
R1371 B.n717 B.n716 10.6151
R1372 B.n717 B.n343 10.6151
R1373 B.n728 B.n343 10.6151
R1374 B.n729 B.n728 10.6151
R1375 B.n730 B.n729 10.6151
R1376 B.n730 B.n334 10.6151
R1377 B.n740 B.n334 10.6151
R1378 B.n741 B.n740 10.6151
R1379 B.n743 B.n741 10.6151
R1380 B.n743 B.n742 10.6151
R1381 B.n742 B.n327 10.6151
R1382 B.n754 B.n327 10.6151
R1383 B.n755 B.n754 10.6151
R1384 B.n756 B.n755 10.6151
R1385 B.n757 B.n756 10.6151
R1386 B.n758 B.n757 10.6151
R1387 B.n761 B.n758 10.6151
R1388 B.n762 B.n761 10.6151
R1389 B.n763 B.n762 10.6151
R1390 B.n764 B.n763 10.6151
R1391 B.n766 B.n764 10.6151
R1392 B.n767 B.n766 10.6151
R1393 B.n768 B.n767 10.6151
R1394 B.n769 B.n768 10.6151
R1395 B.n771 B.n769 10.6151
R1396 B.n772 B.n771 10.6151
R1397 B.n773 B.n772 10.6151
R1398 B.n774 B.n773 10.6151
R1399 B.n776 B.n774 10.6151
R1400 B.n777 B.n776 10.6151
R1401 B.n778 B.n777 10.6151
R1402 B.n779 B.n778 10.6151
R1403 B.n781 B.n779 10.6151
R1404 B.n782 B.n781 10.6151
R1405 B.n783 B.n782 10.6151
R1406 B.n784 B.n783 10.6151
R1407 B.n786 B.n784 10.6151
R1408 B.n787 B.n786 10.6151
R1409 B.n788 B.n787 10.6151
R1410 B.n789 B.n788 10.6151
R1411 B.n791 B.n789 10.6151
R1412 B.n792 B.n791 10.6151
R1413 B.n793 B.n792 10.6151
R1414 B.n794 B.n793 10.6151
R1415 B.n796 B.n794 10.6151
R1416 B.n797 B.n796 10.6151
R1417 B.n798 B.n797 10.6151
R1418 B.n864 B.n1 10.6151
R1419 B.n864 B.n863 10.6151
R1420 B.n863 B.n862 10.6151
R1421 B.n862 B.n10 10.6151
R1422 B.n856 B.n10 10.6151
R1423 B.n856 B.n855 10.6151
R1424 B.n855 B.n854 10.6151
R1425 B.n854 B.n18 10.6151
R1426 B.n848 B.n18 10.6151
R1427 B.n848 B.n847 10.6151
R1428 B.n847 B.n846 10.6151
R1429 B.n846 B.n24 10.6151
R1430 B.n840 B.n24 10.6151
R1431 B.n840 B.n839 10.6151
R1432 B.n839 B.n838 10.6151
R1433 B.n838 B.n32 10.6151
R1434 B.n832 B.n32 10.6151
R1435 B.n832 B.n831 10.6151
R1436 B.n831 B.n830 10.6151
R1437 B.n830 B.n39 10.6151
R1438 B.n824 B.n39 10.6151
R1439 B.n824 B.n823 10.6151
R1440 B.n823 B.n822 10.6151
R1441 B.n822 B.n46 10.6151
R1442 B.n816 B.n46 10.6151
R1443 B.n816 B.n815 10.6151
R1444 B.n815 B.n814 10.6151
R1445 B.n814 B.n52 10.6151
R1446 B.n808 B.n52 10.6151
R1447 B.n808 B.n807 10.6151
R1448 B.n807 B.n806 10.6151
R1449 B.n806 B.n60 10.6151
R1450 B.n122 B.n121 10.6151
R1451 B.n125 B.n122 10.6151
R1452 B.n126 B.n125 10.6151
R1453 B.n129 B.n126 10.6151
R1454 B.n130 B.n129 10.6151
R1455 B.n133 B.n130 10.6151
R1456 B.n134 B.n133 10.6151
R1457 B.n137 B.n134 10.6151
R1458 B.n138 B.n137 10.6151
R1459 B.n141 B.n138 10.6151
R1460 B.n142 B.n141 10.6151
R1461 B.n145 B.n142 10.6151
R1462 B.n146 B.n145 10.6151
R1463 B.n149 B.n146 10.6151
R1464 B.n150 B.n149 10.6151
R1465 B.n153 B.n150 10.6151
R1466 B.n154 B.n153 10.6151
R1467 B.n157 B.n154 10.6151
R1468 B.n158 B.n157 10.6151
R1469 B.n161 B.n158 10.6151
R1470 B.n162 B.n161 10.6151
R1471 B.n165 B.n162 10.6151
R1472 B.n166 B.n165 10.6151
R1473 B.n169 B.n166 10.6151
R1474 B.n170 B.n169 10.6151
R1475 B.n173 B.n170 10.6151
R1476 B.n174 B.n173 10.6151
R1477 B.n177 B.n174 10.6151
R1478 B.n178 B.n177 10.6151
R1479 B.n181 B.n178 10.6151
R1480 B.n182 B.n181 10.6151
R1481 B.n185 B.n182 10.6151
R1482 B.n186 B.n185 10.6151
R1483 B.n189 B.n186 10.6151
R1484 B.n190 B.n189 10.6151
R1485 B.n193 B.n190 10.6151
R1486 B.n194 B.n193 10.6151
R1487 B.n197 B.n194 10.6151
R1488 B.n198 B.n197 10.6151
R1489 B.n201 B.n198 10.6151
R1490 B.n202 B.n201 10.6151
R1491 B.n205 B.n202 10.6151
R1492 B.n206 B.n205 10.6151
R1493 B.n209 B.n206 10.6151
R1494 B.n210 B.n209 10.6151
R1495 B.n213 B.n210 10.6151
R1496 B.n218 B.n215 10.6151
R1497 B.n219 B.n218 10.6151
R1498 B.n222 B.n219 10.6151
R1499 B.n223 B.n222 10.6151
R1500 B.n226 B.n223 10.6151
R1501 B.n227 B.n226 10.6151
R1502 B.n230 B.n227 10.6151
R1503 B.n231 B.n230 10.6151
R1504 B.n234 B.n231 10.6151
R1505 B.n239 B.n236 10.6151
R1506 B.n240 B.n239 10.6151
R1507 B.n243 B.n240 10.6151
R1508 B.n244 B.n243 10.6151
R1509 B.n247 B.n244 10.6151
R1510 B.n248 B.n247 10.6151
R1511 B.n251 B.n248 10.6151
R1512 B.n252 B.n251 10.6151
R1513 B.n255 B.n252 10.6151
R1514 B.n256 B.n255 10.6151
R1515 B.n259 B.n256 10.6151
R1516 B.n260 B.n259 10.6151
R1517 B.n263 B.n260 10.6151
R1518 B.n264 B.n263 10.6151
R1519 B.n267 B.n264 10.6151
R1520 B.n268 B.n267 10.6151
R1521 B.n271 B.n268 10.6151
R1522 B.n272 B.n271 10.6151
R1523 B.n275 B.n272 10.6151
R1524 B.n276 B.n275 10.6151
R1525 B.n279 B.n276 10.6151
R1526 B.n280 B.n279 10.6151
R1527 B.n283 B.n280 10.6151
R1528 B.n284 B.n283 10.6151
R1529 B.n287 B.n284 10.6151
R1530 B.n288 B.n287 10.6151
R1531 B.n291 B.n288 10.6151
R1532 B.n292 B.n291 10.6151
R1533 B.n295 B.n292 10.6151
R1534 B.n296 B.n295 10.6151
R1535 B.n299 B.n296 10.6151
R1536 B.n300 B.n299 10.6151
R1537 B.n303 B.n300 10.6151
R1538 B.n304 B.n303 10.6151
R1539 B.n307 B.n304 10.6151
R1540 B.n308 B.n307 10.6151
R1541 B.n311 B.n308 10.6151
R1542 B.n312 B.n311 10.6151
R1543 B.n315 B.n312 10.6151
R1544 B.n316 B.n315 10.6151
R1545 B.n319 B.n316 10.6151
R1546 B.n320 B.n319 10.6151
R1547 B.n323 B.n320 10.6151
R1548 B.n325 B.n323 10.6151
R1549 B.n326 B.n325 10.6151
R1550 B.n799 B.n326 10.6151
R1551 B.n745 B.t19 10.3264
R1552 B.n860 B.t1 10.3264
R1553 B.n560 B.n445 9.36635
R1554 B.n537 B.n448 9.36635
R1555 B.n214 B.n213 9.36635
R1556 B.n236 B.n235 9.36635
R1557 B.n872 B.n0 8.11757
R1558 B.n872 B.n1 8.11757
R1559 B.n360 B.t4 3.44248
R1560 B.t2 B.n835 3.44248
R1561 B.n557 B.n445 1.24928
R1562 B.n540 B.n448 1.24928
R1563 B.n215 B.n214 1.24928
R1564 B.n235 B.n234 1.24928
R1565 VN.n2 VN.t5 214.252
R1566 VN.n14 VN.t1 214.252
R1567 VN.n3 VN.t4 184.06
R1568 VN.n10 VN.t3 184.06
R1569 VN.n15 VN.t2 184.06
R1570 VN.n22 VN.t0 184.06
R1571 VN.n21 VN.n12 161.3
R1572 VN.n20 VN.n19 161.3
R1573 VN.n18 VN.n13 161.3
R1574 VN.n17 VN.n16 161.3
R1575 VN.n9 VN.n0 161.3
R1576 VN.n8 VN.n7 161.3
R1577 VN.n6 VN.n1 161.3
R1578 VN.n5 VN.n4 161.3
R1579 VN.n11 VN.n10 91.1314
R1580 VN.n23 VN.n22 91.1314
R1581 VN.n3 VN.n2 57.3616
R1582 VN.n15 VN.n14 57.3616
R1583 VN.n8 VN.n1 56.4773
R1584 VN.n20 VN.n13 56.4773
R1585 VN VN.n23 47.3125
R1586 VN.n4 VN.n1 24.3439
R1587 VN.n9 VN.n8 24.3439
R1588 VN.n16 VN.n13 24.3439
R1589 VN.n21 VN.n20 24.3439
R1590 VN.n10 VN.n9 19.4752
R1591 VN.n22 VN.n21 19.4752
R1592 VN.n17 VN.n14 13.3877
R1593 VN.n5 VN.n2 13.3877
R1594 VN.n4 VN.n3 12.1722
R1595 VN.n16 VN.n15 12.1722
R1596 VN.n23 VN.n12 0.278398
R1597 VN.n11 VN.n0 0.278398
R1598 VN.n19 VN.n12 0.189894
R1599 VN.n19 VN.n18 0.189894
R1600 VN.n18 VN.n17 0.189894
R1601 VN.n6 VN.n5 0.189894
R1602 VN.n7 VN.n6 0.189894
R1603 VN.n7 VN.n0 0.189894
R1604 VN VN.n11 0.153422
R1605 VDD2.n1 VDD2.t0 63.8595
R1606 VDD2.n2 VDD2.t5 62.5248
R1607 VDD2.n1 VDD2.n0 61.5084
R1608 VDD2 VDD2.n3 61.5056
R1609 VDD2.n2 VDD2.n1 41.7218
R1610 VDD2 VDD2.n2 1.44878
R1611 VDD2.n3 VDD2.t3 1.42496
R1612 VDD2.n3 VDD2.t4 1.42496
R1613 VDD2.n0 VDD2.t1 1.42496
R1614 VDD2.n0 VDD2.t2 1.42496
C0 VDD2 VTAIL 8.628611f
C1 VP VN 6.52936f
C2 VDD1 VN 0.149411f
C3 VTAIL VN 7.03114f
C4 VP VDD1 7.36883f
C5 VP VTAIL 7.04555f
C6 VDD1 VTAIL 8.58467f
C7 VDD2 VN 7.12998f
C8 VP VDD2 0.392186f
C9 VDD2 VDD1 1.1291f
C10 VDD2 B 5.70362f
C11 VDD1 B 5.992865f
C12 VTAIL B 8.028408f
C13 VN B 10.85442f
C14 VP B 9.297828f
C15 VDD2.t0 B 2.70506f
C16 VDD2.t1 B 0.235317f
C17 VDD2.t2 B 0.235317f
C18 VDD2.n0 B 2.11593f
C19 VDD2.n1 B 2.31048f
C20 VDD2.t5 B 2.69799f
C21 VDD2.n2 B 2.34319f
C22 VDD2.t3 B 0.235317f
C23 VDD2.t4 B 0.235317f
C24 VDD2.n3 B 2.1159f
C25 VN.n0 B 0.037606f
C26 VN.t3 B 1.97363f
C27 VN.n1 B 0.047821f
C28 VN.t5 B 2.09062f
C29 VN.n2 B 0.776338f
C30 VN.t4 B 1.97363f
C31 VN.n3 B 0.764521f
C32 VN.n4 B 0.040236f
C33 VN.n5 B 0.208857f
C34 VN.n6 B 0.028522f
C35 VN.n7 B 0.028522f
C36 VN.n8 B 0.035815f
C37 VN.n9 B 0.048149f
C38 VN.n10 B 0.780161f
C39 VN.n11 B 0.033951f
C40 VN.n12 B 0.037606f
C41 VN.t0 B 1.97363f
C42 VN.n13 B 0.047821f
C43 VN.t1 B 2.09062f
C44 VN.n14 B 0.776338f
C45 VN.t2 B 1.97363f
C46 VN.n15 B 0.764521f
C47 VN.n16 B 0.040236f
C48 VN.n17 B 0.208857f
C49 VN.n18 B 0.028522f
C50 VN.n19 B 0.028522f
C51 VN.n20 B 0.035815f
C52 VN.n21 B 0.048149f
C53 VN.n22 B 0.780161f
C54 VN.n23 B 1.45013f
C55 VDD1.t4 B 2.7437f
C56 VDD1.t1 B 2.74292f
C57 VDD1.t2 B 0.238611f
C58 VDD1.t0 B 0.238611f
C59 VDD1.n0 B 2.14554f
C60 VDD1.n1 B 2.43433f
C61 VDD1.t3 B 0.238611f
C62 VDD1.t5 B 0.238611f
C63 VDD1.n2 B 2.14322f
C64 VDD1.n3 B 2.36323f
C65 VTAIL.t1 B 0.251306f
C66 VTAIL.t0 B 0.251306f
C67 VTAIL.n0 B 2.18671f
C68 VTAIL.n1 B 0.373022f
C69 VTAIL.t8 B 2.79065f
C70 VTAIL.n2 B 0.552654f
C71 VTAIL.t7 B 0.251306f
C72 VTAIL.t6 B 0.251306f
C73 VTAIL.n3 B 2.18671f
C74 VTAIL.n4 B 1.83569f
C75 VTAIL.t4 B 0.251306f
C76 VTAIL.t3 B 0.251306f
C77 VTAIL.n5 B 2.18671f
C78 VTAIL.n6 B 1.83569f
C79 VTAIL.t11 B 2.79067f
C80 VTAIL.n7 B 0.552637f
C81 VTAIL.t5 B 0.251306f
C82 VTAIL.t9 B 0.251306f
C83 VTAIL.n8 B 2.18671f
C84 VTAIL.n9 B 0.471212f
C85 VTAIL.t10 B 2.79066f
C86 VTAIL.n10 B 1.78048f
C87 VTAIL.t2 B 2.79065f
C88 VTAIL.n11 B 1.74205f
C89 VP.n0 B 0.038228f
C90 VP.t5 B 2.00628f
C91 VP.n1 B 0.048612f
C92 VP.n2 B 0.028994f
C93 VP.t3 B 2.00628f
C94 VP.n3 B 0.036408f
C95 VP.n4 B 0.038228f
C96 VP.t0 B 2.00628f
C97 VP.n5 B 0.048612f
C98 VP.t1 B 2.1252f
C99 VP.n6 B 0.78918f
C100 VP.t2 B 2.00628f
C101 VP.n7 B 0.777168f
C102 VP.n8 B 0.040901f
C103 VP.n9 B 0.212312f
C104 VP.n10 B 0.028994f
C105 VP.n11 B 0.028994f
C106 VP.n12 B 0.036408f
C107 VP.n13 B 0.048945f
C108 VP.n14 B 0.793066f
C109 VP.n15 B 1.45838f
C110 VP.n16 B 1.48048f
C111 VP.t4 B 2.00628f
C112 VP.n17 B 0.793066f
C113 VP.n18 B 0.048945f
C114 VP.n19 B 0.038228f
C115 VP.n20 B 0.028994f
C116 VP.n21 B 0.028994f
C117 VP.n22 B 0.048612f
C118 VP.n23 B 0.040901f
C119 VP.n24 B 0.712006f
C120 VP.n25 B 0.040901f
C121 VP.n26 B 0.028994f
C122 VP.n27 B 0.028994f
C123 VP.n28 B 0.028994f
C124 VP.n29 B 0.036408f
C125 VP.n30 B 0.048945f
C126 VP.n31 B 0.793066f
C127 VP.n32 B 0.034512f
.ends

