* NGSPICE file created from diff_pair_sample_1400.ext - technology: sky130A

.subckt diff_pair_sample_1400 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=2.7495 pd=14.88 as=0 ps=0 w=7.05 l=3.48
X1 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=2.7495 pd=14.88 as=0 ps=0 w=7.05 l=3.48
X2 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7495 pd=14.88 as=0 ps=0 w=7.05 l=3.48
X3 VDD1.t1 VP.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7495 pd=14.88 as=2.7495 ps=14.88 w=7.05 l=3.48
X4 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7495 pd=14.88 as=2.7495 ps=14.88 w=7.05 l=3.48
X5 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.7495 pd=14.88 as=2.7495 ps=14.88 w=7.05 l=3.48
X6 VDD1.t0 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.7495 pd=14.88 as=2.7495 ps=14.88 w=7.05 l=3.48
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.7495 pd=14.88 as=0 ps=0 w=7.05 l=3.48
R0 B.n450 B.n449 585
R1 B.n452 B.n95 585
R2 B.n455 B.n454 585
R3 B.n456 B.n94 585
R4 B.n458 B.n457 585
R5 B.n460 B.n93 585
R6 B.n463 B.n462 585
R7 B.n464 B.n92 585
R8 B.n466 B.n465 585
R9 B.n468 B.n91 585
R10 B.n471 B.n470 585
R11 B.n472 B.n90 585
R12 B.n474 B.n473 585
R13 B.n476 B.n89 585
R14 B.n479 B.n478 585
R15 B.n480 B.n88 585
R16 B.n482 B.n481 585
R17 B.n484 B.n87 585
R18 B.n487 B.n486 585
R19 B.n488 B.n86 585
R20 B.n490 B.n489 585
R21 B.n492 B.n85 585
R22 B.n495 B.n494 585
R23 B.n496 B.n84 585
R24 B.n498 B.n497 585
R25 B.n500 B.n83 585
R26 B.n503 B.n502 585
R27 B.n505 B.n80 585
R28 B.n507 B.n506 585
R29 B.n509 B.n79 585
R30 B.n512 B.n511 585
R31 B.n513 B.n78 585
R32 B.n515 B.n514 585
R33 B.n517 B.n77 585
R34 B.n520 B.n519 585
R35 B.n521 B.n73 585
R36 B.n523 B.n522 585
R37 B.n525 B.n72 585
R38 B.n528 B.n527 585
R39 B.n529 B.n71 585
R40 B.n531 B.n530 585
R41 B.n533 B.n70 585
R42 B.n536 B.n535 585
R43 B.n537 B.n69 585
R44 B.n539 B.n538 585
R45 B.n541 B.n68 585
R46 B.n544 B.n543 585
R47 B.n545 B.n67 585
R48 B.n547 B.n546 585
R49 B.n549 B.n66 585
R50 B.n552 B.n551 585
R51 B.n553 B.n65 585
R52 B.n555 B.n554 585
R53 B.n557 B.n64 585
R54 B.n560 B.n559 585
R55 B.n561 B.n63 585
R56 B.n563 B.n562 585
R57 B.n565 B.n62 585
R58 B.n568 B.n567 585
R59 B.n569 B.n61 585
R60 B.n571 B.n570 585
R61 B.n573 B.n60 585
R62 B.n576 B.n575 585
R63 B.n577 B.n59 585
R64 B.n448 B.n57 585
R65 B.n580 B.n57 585
R66 B.n447 B.n56 585
R67 B.n581 B.n56 585
R68 B.n446 B.n55 585
R69 B.n582 B.n55 585
R70 B.n445 B.n444 585
R71 B.n444 B.n51 585
R72 B.n443 B.n50 585
R73 B.n588 B.n50 585
R74 B.n442 B.n49 585
R75 B.n589 B.n49 585
R76 B.n441 B.n48 585
R77 B.n590 B.n48 585
R78 B.n440 B.n439 585
R79 B.n439 B.n44 585
R80 B.n438 B.n43 585
R81 B.n596 B.n43 585
R82 B.n437 B.n42 585
R83 B.n597 B.n42 585
R84 B.n436 B.n41 585
R85 B.n598 B.n41 585
R86 B.n435 B.n434 585
R87 B.n434 B.n37 585
R88 B.n433 B.n36 585
R89 B.n604 B.n36 585
R90 B.n432 B.n35 585
R91 B.n605 B.n35 585
R92 B.n431 B.n34 585
R93 B.n606 B.n34 585
R94 B.n430 B.n429 585
R95 B.n429 B.n30 585
R96 B.n428 B.n29 585
R97 B.n612 B.n29 585
R98 B.n427 B.n28 585
R99 B.n613 B.n28 585
R100 B.n426 B.n27 585
R101 B.n614 B.n27 585
R102 B.n425 B.n424 585
R103 B.n424 B.n23 585
R104 B.n423 B.n22 585
R105 B.n620 B.n22 585
R106 B.n422 B.n21 585
R107 B.n621 B.n21 585
R108 B.n421 B.n20 585
R109 B.n622 B.n20 585
R110 B.n420 B.n419 585
R111 B.n419 B.n19 585
R112 B.n418 B.n15 585
R113 B.n628 B.n15 585
R114 B.n417 B.n14 585
R115 B.n629 B.n14 585
R116 B.n416 B.n13 585
R117 B.n630 B.n13 585
R118 B.n415 B.n414 585
R119 B.n414 B.n12 585
R120 B.n413 B.n412 585
R121 B.n413 B.n8 585
R122 B.n411 B.n7 585
R123 B.n637 B.n7 585
R124 B.n410 B.n6 585
R125 B.n638 B.n6 585
R126 B.n409 B.n5 585
R127 B.n639 B.n5 585
R128 B.n408 B.n407 585
R129 B.n407 B.n4 585
R130 B.n406 B.n96 585
R131 B.n406 B.n405 585
R132 B.n396 B.n97 585
R133 B.n98 B.n97 585
R134 B.n398 B.n397 585
R135 B.n399 B.n398 585
R136 B.n395 B.n103 585
R137 B.n103 B.n102 585
R138 B.n394 B.n393 585
R139 B.n393 B.n392 585
R140 B.n105 B.n104 585
R141 B.n385 B.n105 585
R142 B.n384 B.n383 585
R143 B.n386 B.n384 585
R144 B.n382 B.n110 585
R145 B.n110 B.n109 585
R146 B.n381 B.n380 585
R147 B.n380 B.n379 585
R148 B.n112 B.n111 585
R149 B.n113 B.n112 585
R150 B.n372 B.n371 585
R151 B.n373 B.n372 585
R152 B.n370 B.n118 585
R153 B.n118 B.n117 585
R154 B.n369 B.n368 585
R155 B.n368 B.n367 585
R156 B.n120 B.n119 585
R157 B.n121 B.n120 585
R158 B.n360 B.n359 585
R159 B.n361 B.n360 585
R160 B.n358 B.n126 585
R161 B.n126 B.n125 585
R162 B.n357 B.n356 585
R163 B.n356 B.n355 585
R164 B.n128 B.n127 585
R165 B.n129 B.n128 585
R166 B.n348 B.n347 585
R167 B.n349 B.n348 585
R168 B.n346 B.n134 585
R169 B.n134 B.n133 585
R170 B.n345 B.n344 585
R171 B.n344 B.n343 585
R172 B.n136 B.n135 585
R173 B.n137 B.n136 585
R174 B.n336 B.n335 585
R175 B.n337 B.n336 585
R176 B.n334 B.n142 585
R177 B.n142 B.n141 585
R178 B.n333 B.n332 585
R179 B.n332 B.n331 585
R180 B.n144 B.n143 585
R181 B.n145 B.n144 585
R182 B.n324 B.n323 585
R183 B.n325 B.n324 585
R184 B.n322 B.n150 585
R185 B.n150 B.n149 585
R186 B.n321 B.n320 585
R187 B.n320 B.n319 585
R188 B.n316 B.n154 585
R189 B.n315 B.n314 585
R190 B.n312 B.n155 585
R191 B.n312 B.n153 585
R192 B.n311 B.n310 585
R193 B.n309 B.n308 585
R194 B.n307 B.n157 585
R195 B.n305 B.n304 585
R196 B.n303 B.n158 585
R197 B.n302 B.n301 585
R198 B.n299 B.n159 585
R199 B.n297 B.n296 585
R200 B.n295 B.n160 585
R201 B.n294 B.n293 585
R202 B.n291 B.n161 585
R203 B.n289 B.n288 585
R204 B.n287 B.n162 585
R205 B.n286 B.n285 585
R206 B.n283 B.n163 585
R207 B.n281 B.n280 585
R208 B.n279 B.n164 585
R209 B.n278 B.n277 585
R210 B.n275 B.n165 585
R211 B.n273 B.n272 585
R212 B.n271 B.n166 585
R213 B.n270 B.n269 585
R214 B.n267 B.n167 585
R215 B.n265 B.n264 585
R216 B.n262 B.n168 585
R217 B.n261 B.n260 585
R218 B.n258 B.n171 585
R219 B.n256 B.n255 585
R220 B.n254 B.n172 585
R221 B.n253 B.n252 585
R222 B.n250 B.n173 585
R223 B.n248 B.n247 585
R224 B.n246 B.n174 585
R225 B.n245 B.n244 585
R226 B.n242 B.n241 585
R227 B.n240 B.n239 585
R228 B.n238 B.n179 585
R229 B.n236 B.n235 585
R230 B.n234 B.n180 585
R231 B.n233 B.n232 585
R232 B.n230 B.n181 585
R233 B.n228 B.n227 585
R234 B.n226 B.n182 585
R235 B.n225 B.n224 585
R236 B.n222 B.n183 585
R237 B.n220 B.n219 585
R238 B.n218 B.n184 585
R239 B.n217 B.n216 585
R240 B.n214 B.n185 585
R241 B.n212 B.n211 585
R242 B.n210 B.n186 585
R243 B.n209 B.n208 585
R244 B.n206 B.n187 585
R245 B.n204 B.n203 585
R246 B.n202 B.n188 585
R247 B.n201 B.n200 585
R248 B.n198 B.n189 585
R249 B.n196 B.n195 585
R250 B.n194 B.n190 585
R251 B.n193 B.n192 585
R252 B.n152 B.n151 585
R253 B.n153 B.n152 585
R254 B.n318 B.n317 585
R255 B.n319 B.n318 585
R256 B.n148 B.n147 585
R257 B.n149 B.n148 585
R258 B.n327 B.n326 585
R259 B.n326 B.n325 585
R260 B.n328 B.n146 585
R261 B.n146 B.n145 585
R262 B.n330 B.n329 585
R263 B.n331 B.n330 585
R264 B.n140 B.n139 585
R265 B.n141 B.n140 585
R266 B.n339 B.n338 585
R267 B.n338 B.n337 585
R268 B.n340 B.n138 585
R269 B.n138 B.n137 585
R270 B.n342 B.n341 585
R271 B.n343 B.n342 585
R272 B.n132 B.n131 585
R273 B.n133 B.n132 585
R274 B.n351 B.n350 585
R275 B.n350 B.n349 585
R276 B.n352 B.n130 585
R277 B.n130 B.n129 585
R278 B.n354 B.n353 585
R279 B.n355 B.n354 585
R280 B.n124 B.n123 585
R281 B.n125 B.n124 585
R282 B.n363 B.n362 585
R283 B.n362 B.n361 585
R284 B.n364 B.n122 585
R285 B.n122 B.n121 585
R286 B.n366 B.n365 585
R287 B.n367 B.n366 585
R288 B.n116 B.n115 585
R289 B.n117 B.n116 585
R290 B.n375 B.n374 585
R291 B.n374 B.n373 585
R292 B.n376 B.n114 585
R293 B.n114 B.n113 585
R294 B.n378 B.n377 585
R295 B.n379 B.n378 585
R296 B.n108 B.n107 585
R297 B.n109 B.n108 585
R298 B.n388 B.n387 585
R299 B.n387 B.n386 585
R300 B.n389 B.n106 585
R301 B.n385 B.n106 585
R302 B.n391 B.n390 585
R303 B.n392 B.n391 585
R304 B.n101 B.n100 585
R305 B.n102 B.n101 585
R306 B.n401 B.n400 585
R307 B.n400 B.n399 585
R308 B.n402 B.n99 585
R309 B.n99 B.n98 585
R310 B.n404 B.n403 585
R311 B.n405 B.n404 585
R312 B.n3 B.n0 585
R313 B.n4 B.n3 585
R314 B.n636 B.n1 585
R315 B.n637 B.n636 585
R316 B.n635 B.n634 585
R317 B.n635 B.n8 585
R318 B.n633 B.n9 585
R319 B.n12 B.n9 585
R320 B.n632 B.n631 585
R321 B.n631 B.n630 585
R322 B.n11 B.n10 585
R323 B.n629 B.n11 585
R324 B.n627 B.n626 585
R325 B.n628 B.n627 585
R326 B.n625 B.n16 585
R327 B.n19 B.n16 585
R328 B.n624 B.n623 585
R329 B.n623 B.n622 585
R330 B.n18 B.n17 585
R331 B.n621 B.n18 585
R332 B.n619 B.n618 585
R333 B.n620 B.n619 585
R334 B.n617 B.n24 585
R335 B.n24 B.n23 585
R336 B.n616 B.n615 585
R337 B.n615 B.n614 585
R338 B.n26 B.n25 585
R339 B.n613 B.n26 585
R340 B.n611 B.n610 585
R341 B.n612 B.n611 585
R342 B.n609 B.n31 585
R343 B.n31 B.n30 585
R344 B.n608 B.n607 585
R345 B.n607 B.n606 585
R346 B.n33 B.n32 585
R347 B.n605 B.n33 585
R348 B.n603 B.n602 585
R349 B.n604 B.n603 585
R350 B.n601 B.n38 585
R351 B.n38 B.n37 585
R352 B.n600 B.n599 585
R353 B.n599 B.n598 585
R354 B.n40 B.n39 585
R355 B.n597 B.n40 585
R356 B.n595 B.n594 585
R357 B.n596 B.n595 585
R358 B.n593 B.n45 585
R359 B.n45 B.n44 585
R360 B.n592 B.n591 585
R361 B.n591 B.n590 585
R362 B.n47 B.n46 585
R363 B.n589 B.n47 585
R364 B.n587 B.n586 585
R365 B.n588 B.n587 585
R366 B.n585 B.n52 585
R367 B.n52 B.n51 585
R368 B.n584 B.n583 585
R369 B.n583 B.n582 585
R370 B.n54 B.n53 585
R371 B.n581 B.n54 585
R372 B.n579 B.n578 585
R373 B.n580 B.n579 585
R374 B.n640 B.n639 585
R375 B.n638 B.n2 585
R376 B.n579 B.n59 478.086
R377 B.n450 B.n57 478.086
R378 B.n320 B.n152 478.086
R379 B.n318 B.n154 478.086
R380 B.n74 B.t9 257.899
R381 B.n81 B.t13 257.899
R382 B.n175 B.t2 257.899
R383 B.n169 B.t6 257.899
R384 B.n451 B.n58 256.663
R385 B.n453 B.n58 256.663
R386 B.n459 B.n58 256.663
R387 B.n461 B.n58 256.663
R388 B.n467 B.n58 256.663
R389 B.n469 B.n58 256.663
R390 B.n475 B.n58 256.663
R391 B.n477 B.n58 256.663
R392 B.n483 B.n58 256.663
R393 B.n485 B.n58 256.663
R394 B.n491 B.n58 256.663
R395 B.n493 B.n58 256.663
R396 B.n499 B.n58 256.663
R397 B.n501 B.n58 256.663
R398 B.n508 B.n58 256.663
R399 B.n510 B.n58 256.663
R400 B.n516 B.n58 256.663
R401 B.n518 B.n58 256.663
R402 B.n524 B.n58 256.663
R403 B.n526 B.n58 256.663
R404 B.n532 B.n58 256.663
R405 B.n534 B.n58 256.663
R406 B.n540 B.n58 256.663
R407 B.n542 B.n58 256.663
R408 B.n548 B.n58 256.663
R409 B.n550 B.n58 256.663
R410 B.n556 B.n58 256.663
R411 B.n558 B.n58 256.663
R412 B.n564 B.n58 256.663
R413 B.n566 B.n58 256.663
R414 B.n572 B.n58 256.663
R415 B.n574 B.n58 256.663
R416 B.n313 B.n153 256.663
R417 B.n156 B.n153 256.663
R418 B.n306 B.n153 256.663
R419 B.n300 B.n153 256.663
R420 B.n298 B.n153 256.663
R421 B.n292 B.n153 256.663
R422 B.n290 B.n153 256.663
R423 B.n284 B.n153 256.663
R424 B.n282 B.n153 256.663
R425 B.n276 B.n153 256.663
R426 B.n274 B.n153 256.663
R427 B.n268 B.n153 256.663
R428 B.n266 B.n153 256.663
R429 B.n259 B.n153 256.663
R430 B.n257 B.n153 256.663
R431 B.n251 B.n153 256.663
R432 B.n249 B.n153 256.663
R433 B.n243 B.n153 256.663
R434 B.n178 B.n153 256.663
R435 B.n237 B.n153 256.663
R436 B.n231 B.n153 256.663
R437 B.n229 B.n153 256.663
R438 B.n223 B.n153 256.663
R439 B.n221 B.n153 256.663
R440 B.n215 B.n153 256.663
R441 B.n213 B.n153 256.663
R442 B.n207 B.n153 256.663
R443 B.n205 B.n153 256.663
R444 B.n199 B.n153 256.663
R445 B.n197 B.n153 256.663
R446 B.n191 B.n153 256.663
R447 B.n642 B.n641 256.663
R448 B.n575 B.n573 163.367
R449 B.n571 B.n61 163.367
R450 B.n567 B.n565 163.367
R451 B.n563 B.n63 163.367
R452 B.n559 B.n557 163.367
R453 B.n555 B.n65 163.367
R454 B.n551 B.n549 163.367
R455 B.n547 B.n67 163.367
R456 B.n543 B.n541 163.367
R457 B.n539 B.n69 163.367
R458 B.n535 B.n533 163.367
R459 B.n531 B.n71 163.367
R460 B.n527 B.n525 163.367
R461 B.n523 B.n73 163.367
R462 B.n519 B.n517 163.367
R463 B.n515 B.n78 163.367
R464 B.n511 B.n509 163.367
R465 B.n507 B.n80 163.367
R466 B.n502 B.n500 163.367
R467 B.n498 B.n84 163.367
R468 B.n494 B.n492 163.367
R469 B.n490 B.n86 163.367
R470 B.n486 B.n484 163.367
R471 B.n482 B.n88 163.367
R472 B.n478 B.n476 163.367
R473 B.n474 B.n90 163.367
R474 B.n470 B.n468 163.367
R475 B.n466 B.n92 163.367
R476 B.n462 B.n460 163.367
R477 B.n458 B.n94 163.367
R478 B.n454 B.n452 163.367
R479 B.n320 B.n150 163.367
R480 B.n324 B.n150 163.367
R481 B.n324 B.n144 163.367
R482 B.n332 B.n144 163.367
R483 B.n332 B.n142 163.367
R484 B.n336 B.n142 163.367
R485 B.n336 B.n136 163.367
R486 B.n344 B.n136 163.367
R487 B.n344 B.n134 163.367
R488 B.n348 B.n134 163.367
R489 B.n348 B.n128 163.367
R490 B.n356 B.n128 163.367
R491 B.n356 B.n126 163.367
R492 B.n360 B.n126 163.367
R493 B.n360 B.n120 163.367
R494 B.n368 B.n120 163.367
R495 B.n368 B.n118 163.367
R496 B.n372 B.n118 163.367
R497 B.n372 B.n112 163.367
R498 B.n380 B.n112 163.367
R499 B.n380 B.n110 163.367
R500 B.n384 B.n110 163.367
R501 B.n384 B.n105 163.367
R502 B.n393 B.n105 163.367
R503 B.n393 B.n103 163.367
R504 B.n398 B.n103 163.367
R505 B.n398 B.n97 163.367
R506 B.n406 B.n97 163.367
R507 B.n407 B.n406 163.367
R508 B.n407 B.n5 163.367
R509 B.n6 B.n5 163.367
R510 B.n7 B.n6 163.367
R511 B.n413 B.n7 163.367
R512 B.n414 B.n413 163.367
R513 B.n414 B.n13 163.367
R514 B.n14 B.n13 163.367
R515 B.n15 B.n14 163.367
R516 B.n419 B.n15 163.367
R517 B.n419 B.n20 163.367
R518 B.n21 B.n20 163.367
R519 B.n22 B.n21 163.367
R520 B.n424 B.n22 163.367
R521 B.n424 B.n27 163.367
R522 B.n28 B.n27 163.367
R523 B.n29 B.n28 163.367
R524 B.n429 B.n29 163.367
R525 B.n429 B.n34 163.367
R526 B.n35 B.n34 163.367
R527 B.n36 B.n35 163.367
R528 B.n434 B.n36 163.367
R529 B.n434 B.n41 163.367
R530 B.n42 B.n41 163.367
R531 B.n43 B.n42 163.367
R532 B.n439 B.n43 163.367
R533 B.n439 B.n48 163.367
R534 B.n49 B.n48 163.367
R535 B.n50 B.n49 163.367
R536 B.n444 B.n50 163.367
R537 B.n444 B.n55 163.367
R538 B.n56 B.n55 163.367
R539 B.n57 B.n56 163.367
R540 B.n314 B.n312 163.367
R541 B.n312 B.n311 163.367
R542 B.n308 B.n307 163.367
R543 B.n305 B.n158 163.367
R544 B.n301 B.n299 163.367
R545 B.n297 B.n160 163.367
R546 B.n293 B.n291 163.367
R547 B.n289 B.n162 163.367
R548 B.n285 B.n283 163.367
R549 B.n281 B.n164 163.367
R550 B.n277 B.n275 163.367
R551 B.n273 B.n166 163.367
R552 B.n269 B.n267 163.367
R553 B.n265 B.n168 163.367
R554 B.n260 B.n258 163.367
R555 B.n256 B.n172 163.367
R556 B.n252 B.n250 163.367
R557 B.n248 B.n174 163.367
R558 B.n244 B.n242 163.367
R559 B.n239 B.n238 163.367
R560 B.n236 B.n180 163.367
R561 B.n232 B.n230 163.367
R562 B.n228 B.n182 163.367
R563 B.n224 B.n222 163.367
R564 B.n220 B.n184 163.367
R565 B.n216 B.n214 163.367
R566 B.n212 B.n186 163.367
R567 B.n208 B.n206 163.367
R568 B.n204 B.n188 163.367
R569 B.n200 B.n198 163.367
R570 B.n196 B.n190 163.367
R571 B.n192 B.n152 163.367
R572 B.n318 B.n148 163.367
R573 B.n326 B.n148 163.367
R574 B.n326 B.n146 163.367
R575 B.n330 B.n146 163.367
R576 B.n330 B.n140 163.367
R577 B.n338 B.n140 163.367
R578 B.n338 B.n138 163.367
R579 B.n342 B.n138 163.367
R580 B.n342 B.n132 163.367
R581 B.n350 B.n132 163.367
R582 B.n350 B.n130 163.367
R583 B.n354 B.n130 163.367
R584 B.n354 B.n124 163.367
R585 B.n362 B.n124 163.367
R586 B.n362 B.n122 163.367
R587 B.n366 B.n122 163.367
R588 B.n366 B.n116 163.367
R589 B.n374 B.n116 163.367
R590 B.n374 B.n114 163.367
R591 B.n378 B.n114 163.367
R592 B.n378 B.n108 163.367
R593 B.n387 B.n108 163.367
R594 B.n387 B.n106 163.367
R595 B.n391 B.n106 163.367
R596 B.n391 B.n101 163.367
R597 B.n400 B.n101 163.367
R598 B.n400 B.n99 163.367
R599 B.n404 B.n99 163.367
R600 B.n404 B.n3 163.367
R601 B.n640 B.n3 163.367
R602 B.n636 B.n2 163.367
R603 B.n636 B.n635 163.367
R604 B.n635 B.n9 163.367
R605 B.n631 B.n9 163.367
R606 B.n631 B.n11 163.367
R607 B.n627 B.n11 163.367
R608 B.n627 B.n16 163.367
R609 B.n623 B.n16 163.367
R610 B.n623 B.n18 163.367
R611 B.n619 B.n18 163.367
R612 B.n619 B.n24 163.367
R613 B.n615 B.n24 163.367
R614 B.n615 B.n26 163.367
R615 B.n611 B.n26 163.367
R616 B.n611 B.n31 163.367
R617 B.n607 B.n31 163.367
R618 B.n607 B.n33 163.367
R619 B.n603 B.n33 163.367
R620 B.n603 B.n38 163.367
R621 B.n599 B.n38 163.367
R622 B.n599 B.n40 163.367
R623 B.n595 B.n40 163.367
R624 B.n595 B.n45 163.367
R625 B.n591 B.n45 163.367
R626 B.n591 B.n47 163.367
R627 B.n587 B.n47 163.367
R628 B.n587 B.n52 163.367
R629 B.n583 B.n52 163.367
R630 B.n583 B.n54 163.367
R631 B.n579 B.n54 163.367
R632 B.n81 B.t14 147.685
R633 B.n175 B.t5 147.685
R634 B.n74 B.t11 147.677
R635 B.n169 B.t8 147.677
R636 B.n319 B.n153 111.562
R637 B.n580 B.n58 111.562
R638 B.n75 B.n74 73.8914
R639 B.n82 B.n81 73.8914
R640 B.n176 B.n175 73.8914
R641 B.n170 B.n169 73.8914
R642 B.n82 B.t15 73.7934
R643 B.n176 B.t4 73.7934
R644 B.n75 B.t12 73.7857
R645 B.n170 B.t7 73.7857
R646 B.n574 B.n59 71.676
R647 B.n573 B.n572 71.676
R648 B.n566 B.n61 71.676
R649 B.n565 B.n564 71.676
R650 B.n558 B.n63 71.676
R651 B.n557 B.n556 71.676
R652 B.n550 B.n65 71.676
R653 B.n549 B.n548 71.676
R654 B.n542 B.n67 71.676
R655 B.n541 B.n540 71.676
R656 B.n534 B.n69 71.676
R657 B.n533 B.n532 71.676
R658 B.n526 B.n71 71.676
R659 B.n525 B.n524 71.676
R660 B.n518 B.n73 71.676
R661 B.n517 B.n516 71.676
R662 B.n510 B.n78 71.676
R663 B.n509 B.n508 71.676
R664 B.n501 B.n80 71.676
R665 B.n500 B.n499 71.676
R666 B.n493 B.n84 71.676
R667 B.n492 B.n491 71.676
R668 B.n485 B.n86 71.676
R669 B.n484 B.n483 71.676
R670 B.n477 B.n88 71.676
R671 B.n476 B.n475 71.676
R672 B.n469 B.n90 71.676
R673 B.n468 B.n467 71.676
R674 B.n461 B.n92 71.676
R675 B.n460 B.n459 71.676
R676 B.n453 B.n94 71.676
R677 B.n452 B.n451 71.676
R678 B.n451 B.n450 71.676
R679 B.n454 B.n453 71.676
R680 B.n459 B.n458 71.676
R681 B.n462 B.n461 71.676
R682 B.n467 B.n466 71.676
R683 B.n470 B.n469 71.676
R684 B.n475 B.n474 71.676
R685 B.n478 B.n477 71.676
R686 B.n483 B.n482 71.676
R687 B.n486 B.n485 71.676
R688 B.n491 B.n490 71.676
R689 B.n494 B.n493 71.676
R690 B.n499 B.n498 71.676
R691 B.n502 B.n501 71.676
R692 B.n508 B.n507 71.676
R693 B.n511 B.n510 71.676
R694 B.n516 B.n515 71.676
R695 B.n519 B.n518 71.676
R696 B.n524 B.n523 71.676
R697 B.n527 B.n526 71.676
R698 B.n532 B.n531 71.676
R699 B.n535 B.n534 71.676
R700 B.n540 B.n539 71.676
R701 B.n543 B.n542 71.676
R702 B.n548 B.n547 71.676
R703 B.n551 B.n550 71.676
R704 B.n556 B.n555 71.676
R705 B.n559 B.n558 71.676
R706 B.n564 B.n563 71.676
R707 B.n567 B.n566 71.676
R708 B.n572 B.n571 71.676
R709 B.n575 B.n574 71.676
R710 B.n313 B.n154 71.676
R711 B.n311 B.n156 71.676
R712 B.n307 B.n306 71.676
R713 B.n300 B.n158 71.676
R714 B.n299 B.n298 71.676
R715 B.n292 B.n160 71.676
R716 B.n291 B.n290 71.676
R717 B.n284 B.n162 71.676
R718 B.n283 B.n282 71.676
R719 B.n276 B.n164 71.676
R720 B.n275 B.n274 71.676
R721 B.n268 B.n166 71.676
R722 B.n267 B.n266 71.676
R723 B.n259 B.n168 71.676
R724 B.n258 B.n257 71.676
R725 B.n251 B.n172 71.676
R726 B.n250 B.n249 71.676
R727 B.n243 B.n174 71.676
R728 B.n242 B.n178 71.676
R729 B.n238 B.n237 71.676
R730 B.n231 B.n180 71.676
R731 B.n230 B.n229 71.676
R732 B.n223 B.n182 71.676
R733 B.n222 B.n221 71.676
R734 B.n215 B.n184 71.676
R735 B.n214 B.n213 71.676
R736 B.n207 B.n186 71.676
R737 B.n206 B.n205 71.676
R738 B.n199 B.n188 71.676
R739 B.n198 B.n197 71.676
R740 B.n191 B.n190 71.676
R741 B.n314 B.n313 71.676
R742 B.n308 B.n156 71.676
R743 B.n306 B.n305 71.676
R744 B.n301 B.n300 71.676
R745 B.n298 B.n297 71.676
R746 B.n293 B.n292 71.676
R747 B.n290 B.n289 71.676
R748 B.n285 B.n284 71.676
R749 B.n282 B.n281 71.676
R750 B.n277 B.n276 71.676
R751 B.n274 B.n273 71.676
R752 B.n269 B.n268 71.676
R753 B.n266 B.n265 71.676
R754 B.n260 B.n259 71.676
R755 B.n257 B.n256 71.676
R756 B.n252 B.n251 71.676
R757 B.n249 B.n248 71.676
R758 B.n244 B.n243 71.676
R759 B.n239 B.n178 71.676
R760 B.n237 B.n236 71.676
R761 B.n232 B.n231 71.676
R762 B.n229 B.n228 71.676
R763 B.n224 B.n223 71.676
R764 B.n221 B.n220 71.676
R765 B.n216 B.n215 71.676
R766 B.n213 B.n212 71.676
R767 B.n208 B.n207 71.676
R768 B.n205 B.n204 71.676
R769 B.n200 B.n199 71.676
R770 B.n197 B.n196 71.676
R771 B.n192 B.n191 71.676
R772 B.n641 B.n640 71.676
R773 B.n641 B.n2 71.676
R774 B.n319 B.n149 60.6902
R775 B.n325 B.n149 60.6902
R776 B.n325 B.n145 60.6902
R777 B.n331 B.n145 60.6902
R778 B.n331 B.n141 60.6902
R779 B.n337 B.n141 60.6902
R780 B.n337 B.n137 60.6902
R781 B.n343 B.n137 60.6902
R782 B.n349 B.n133 60.6902
R783 B.n349 B.n129 60.6902
R784 B.n355 B.n129 60.6902
R785 B.n355 B.n125 60.6902
R786 B.n361 B.n125 60.6902
R787 B.n361 B.n121 60.6902
R788 B.n367 B.n121 60.6902
R789 B.n367 B.n117 60.6902
R790 B.n373 B.n117 60.6902
R791 B.n373 B.n113 60.6902
R792 B.n379 B.n113 60.6902
R793 B.n379 B.n109 60.6902
R794 B.n386 B.n109 60.6902
R795 B.n386 B.n385 60.6902
R796 B.n392 B.n102 60.6902
R797 B.n399 B.n102 60.6902
R798 B.n399 B.n98 60.6902
R799 B.n405 B.n98 60.6902
R800 B.n405 B.n4 60.6902
R801 B.n639 B.n4 60.6902
R802 B.n639 B.n638 60.6902
R803 B.n638 B.n637 60.6902
R804 B.n637 B.n8 60.6902
R805 B.n12 B.n8 60.6902
R806 B.n630 B.n12 60.6902
R807 B.n630 B.n629 60.6902
R808 B.n629 B.n628 60.6902
R809 B.n622 B.n19 60.6902
R810 B.n622 B.n621 60.6902
R811 B.n621 B.n620 60.6902
R812 B.n620 B.n23 60.6902
R813 B.n614 B.n23 60.6902
R814 B.n614 B.n613 60.6902
R815 B.n613 B.n612 60.6902
R816 B.n612 B.n30 60.6902
R817 B.n606 B.n30 60.6902
R818 B.n606 B.n605 60.6902
R819 B.n605 B.n604 60.6902
R820 B.n604 B.n37 60.6902
R821 B.n598 B.n37 60.6902
R822 B.n598 B.n597 60.6902
R823 B.n596 B.n44 60.6902
R824 B.n590 B.n44 60.6902
R825 B.n590 B.n589 60.6902
R826 B.n589 B.n588 60.6902
R827 B.n588 B.n51 60.6902
R828 B.n582 B.n51 60.6902
R829 B.n582 B.n581 60.6902
R830 B.n581 B.n580 60.6902
R831 B.n76 B.n75 59.5399
R832 B.n504 B.n82 59.5399
R833 B.n177 B.n176 59.5399
R834 B.n263 B.n170 59.5399
R835 B.n343 B.t3 53.5502
R836 B.t10 B.n596 53.5502
R837 B.n392 B.t0 42.8403
R838 B.n628 B.t1 42.8403
R839 B.n317 B.n316 31.0639
R840 B.n321 B.n151 31.0639
R841 B.n449 B.n448 31.0639
R842 B.n578 B.n577 31.0639
R843 B B.n642 18.0485
R844 B.n385 B.t0 17.8504
R845 B.n19 B.t1 17.8504
R846 B.n317 B.n147 10.6151
R847 B.n327 B.n147 10.6151
R848 B.n328 B.n327 10.6151
R849 B.n329 B.n328 10.6151
R850 B.n329 B.n139 10.6151
R851 B.n339 B.n139 10.6151
R852 B.n340 B.n339 10.6151
R853 B.n341 B.n340 10.6151
R854 B.n341 B.n131 10.6151
R855 B.n351 B.n131 10.6151
R856 B.n352 B.n351 10.6151
R857 B.n353 B.n352 10.6151
R858 B.n353 B.n123 10.6151
R859 B.n363 B.n123 10.6151
R860 B.n364 B.n363 10.6151
R861 B.n365 B.n364 10.6151
R862 B.n365 B.n115 10.6151
R863 B.n375 B.n115 10.6151
R864 B.n376 B.n375 10.6151
R865 B.n377 B.n376 10.6151
R866 B.n377 B.n107 10.6151
R867 B.n388 B.n107 10.6151
R868 B.n389 B.n388 10.6151
R869 B.n390 B.n389 10.6151
R870 B.n390 B.n100 10.6151
R871 B.n401 B.n100 10.6151
R872 B.n402 B.n401 10.6151
R873 B.n403 B.n402 10.6151
R874 B.n403 B.n0 10.6151
R875 B.n316 B.n315 10.6151
R876 B.n315 B.n155 10.6151
R877 B.n310 B.n155 10.6151
R878 B.n310 B.n309 10.6151
R879 B.n309 B.n157 10.6151
R880 B.n304 B.n157 10.6151
R881 B.n304 B.n303 10.6151
R882 B.n303 B.n302 10.6151
R883 B.n302 B.n159 10.6151
R884 B.n296 B.n159 10.6151
R885 B.n296 B.n295 10.6151
R886 B.n295 B.n294 10.6151
R887 B.n294 B.n161 10.6151
R888 B.n288 B.n161 10.6151
R889 B.n288 B.n287 10.6151
R890 B.n287 B.n286 10.6151
R891 B.n286 B.n163 10.6151
R892 B.n280 B.n163 10.6151
R893 B.n280 B.n279 10.6151
R894 B.n279 B.n278 10.6151
R895 B.n278 B.n165 10.6151
R896 B.n272 B.n165 10.6151
R897 B.n272 B.n271 10.6151
R898 B.n271 B.n270 10.6151
R899 B.n270 B.n167 10.6151
R900 B.n264 B.n167 10.6151
R901 B.n262 B.n261 10.6151
R902 B.n261 B.n171 10.6151
R903 B.n255 B.n171 10.6151
R904 B.n255 B.n254 10.6151
R905 B.n254 B.n253 10.6151
R906 B.n253 B.n173 10.6151
R907 B.n247 B.n173 10.6151
R908 B.n247 B.n246 10.6151
R909 B.n246 B.n245 10.6151
R910 B.n241 B.n240 10.6151
R911 B.n240 B.n179 10.6151
R912 B.n235 B.n179 10.6151
R913 B.n235 B.n234 10.6151
R914 B.n234 B.n233 10.6151
R915 B.n233 B.n181 10.6151
R916 B.n227 B.n181 10.6151
R917 B.n227 B.n226 10.6151
R918 B.n226 B.n225 10.6151
R919 B.n225 B.n183 10.6151
R920 B.n219 B.n183 10.6151
R921 B.n219 B.n218 10.6151
R922 B.n218 B.n217 10.6151
R923 B.n217 B.n185 10.6151
R924 B.n211 B.n185 10.6151
R925 B.n211 B.n210 10.6151
R926 B.n210 B.n209 10.6151
R927 B.n209 B.n187 10.6151
R928 B.n203 B.n187 10.6151
R929 B.n203 B.n202 10.6151
R930 B.n202 B.n201 10.6151
R931 B.n201 B.n189 10.6151
R932 B.n195 B.n189 10.6151
R933 B.n195 B.n194 10.6151
R934 B.n194 B.n193 10.6151
R935 B.n193 B.n151 10.6151
R936 B.n322 B.n321 10.6151
R937 B.n323 B.n322 10.6151
R938 B.n323 B.n143 10.6151
R939 B.n333 B.n143 10.6151
R940 B.n334 B.n333 10.6151
R941 B.n335 B.n334 10.6151
R942 B.n335 B.n135 10.6151
R943 B.n345 B.n135 10.6151
R944 B.n346 B.n345 10.6151
R945 B.n347 B.n346 10.6151
R946 B.n347 B.n127 10.6151
R947 B.n357 B.n127 10.6151
R948 B.n358 B.n357 10.6151
R949 B.n359 B.n358 10.6151
R950 B.n359 B.n119 10.6151
R951 B.n369 B.n119 10.6151
R952 B.n370 B.n369 10.6151
R953 B.n371 B.n370 10.6151
R954 B.n371 B.n111 10.6151
R955 B.n381 B.n111 10.6151
R956 B.n382 B.n381 10.6151
R957 B.n383 B.n382 10.6151
R958 B.n383 B.n104 10.6151
R959 B.n394 B.n104 10.6151
R960 B.n395 B.n394 10.6151
R961 B.n397 B.n395 10.6151
R962 B.n397 B.n396 10.6151
R963 B.n396 B.n96 10.6151
R964 B.n408 B.n96 10.6151
R965 B.n409 B.n408 10.6151
R966 B.n410 B.n409 10.6151
R967 B.n411 B.n410 10.6151
R968 B.n412 B.n411 10.6151
R969 B.n415 B.n412 10.6151
R970 B.n416 B.n415 10.6151
R971 B.n417 B.n416 10.6151
R972 B.n418 B.n417 10.6151
R973 B.n420 B.n418 10.6151
R974 B.n421 B.n420 10.6151
R975 B.n422 B.n421 10.6151
R976 B.n423 B.n422 10.6151
R977 B.n425 B.n423 10.6151
R978 B.n426 B.n425 10.6151
R979 B.n427 B.n426 10.6151
R980 B.n428 B.n427 10.6151
R981 B.n430 B.n428 10.6151
R982 B.n431 B.n430 10.6151
R983 B.n432 B.n431 10.6151
R984 B.n433 B.n432 10.6151
R985 B.n435 B.n433 10.6151
R986 B.n436 B.n435 10.6151
R987 B.n437 B.n436 10.6151
R988 B.n438 B.n437 10.6151
R989 B.n440 B.n438 10.6151
R990 B.n441 B.n440 10.6151
R991 B.n442 B.n441 10.6151
R992 B.n443 B.n442 10.6151
R993 B.n445 B.n443 10.6151
R994 B.n446 B.n445 10.6151
R995 B.n447 B.n446 10.6151
R996 B.n448 B.n447 10.6151
R997 B.n634 B.n1 10.6151
R998 B.n634 B.n633 10.6151
R999 B.n633 B.n632 10.6151
R1000 B.n632 B.n10 10.6151
R1001 B.n626 B.n10 10.6151
R1002 B.n626 B.n625 10.6151
R1003 B.n625 B.n624 10.6151
R1004 B.n624 B.n17 10.6151
R1005 B.n618 B.n17 10.6151
R1006 B.n618 B.n617 10.6151
R1007 B.n617 B.n616 10.6151
R1008 B.n616 B.n25 10.6151
R1009 B.n610 B.n25 10.6151
R1010 B.n610 B.n609 10.6151
R1011 B.n609 B.n608 10.6151
R1012 B.n608 B.n32 10.6151
R1013 B.n602 B.n32 10.6151
R1014 B.n602 B.n601 10.6151
R1015 B.n601 B.n600 10.6151
R1016 B.n600 B.n39 10.6151
R1017 B.n594 B.n39 10.6151
R1018 B.n594 B.n593 10.6151
R1019 B.n593 B.n592 10.6151
R1020 B.n592 B.n46 10.6151
R1021 B.n586 B.n46 10.6151
R1022 B.n586 B.n585 10.6151
R1023 B.n585 B.n584 10.6151
R1024 B.n584 B.n53 10.6151
R1025 B.n578 B.n53 10.6151
R1026 B.n577 B.n576 10.6151
R1027 B.n576 B.n60 10.6151
R1028 B.n570 B.n60 10.6151
R1029 B.n570 B.n569 10.6151
R1030 B.n569 B.n568 10.6151
R1031 B.n568 B.n62 10.6151
R1032 B.n562 B.n62 10.6151
R1033 B.n562 B.n561 10.6151
R1034 B.n561 B.n560 10.6151
R1035 B.n560 B.n64 10.6151
R1036 B.n554 B.n64 10.6151
R1037 B.n554 B.n553 10.6151
R1038 B.n553 B.n552 10.6151
R1039 B.n552 B.n66 10.6151
R1040 B.n546 B.n66 10.6151
R1041 B.n546 B.n545 10.6151
R1042 B.n545 B.n544 10.6151
R1043 B.n544 B.n68 10.6151
R1044 B.n538 B.n68 10.6151
R1045 B.n538 B.n537 10.6151
R1046 B.n537 B.n536 10.6151
R1047 B.n536 B.n70 10.6151
R1048 B.n530 B.n70 10.6151
R1049 B.n530 B.n529 10.6151
R1050 B.n529 B.n528 10.6151
R1051 B.n528 B.n72 10.6151
R1052 B.n522 B.n521 10.6151
R1053 B.n521 B.n520 10.6151
R1054 B.n520 B.n77 10.6151
R1055 B.n514 B.n77 10.6151
R1056 B.n514 B.n513 10.6151
R1057 B.n513 B.n512 10.6151
R1058 B.n512 B.n79 10.6151
R1059 B.n506 B.n79 10.6151
R1060 B.n506 B.n505 10.6151
R1061 B.n503 B.n83 10.6151
R1062 B.n497 B.n83 10.6151
R1063 B.n497 B.n496 10.6151
R1064 B.n496 B.n495 10.6151
R1065 B.n495 B.n85 10.6151
R1066 B.n489 B.n85 10.6151
R1067 B.n489 B.n488 10.6151
R1068 B.n488 B.n487 10.6151
R1069 B.n487 B.n87 10.6151
R1070 B.n481 B.n87 10.6151
R1071 B.n481 B.n480 10.6151
R1072 B.n480 B.n479 10.6151
R1073 B.n479 B.n89 10.6151
R1074 B.n473 B.n89 10.6151
R1075 B.n473 B.n472 10.6151
R1076 B.n472 B.n471 10.6151
R1077 B.n471 B.n91 10.6151
R1078 B.n465 B.n91 10.6151
R1079 B.n465 B.n464 10.6151
R1080 B.n464 B.n463 10.6151
R1081 B.n463 B.n93 10.6151
R1082 B.n457 B.n93 10.6151
R1083 B.n457 B.n456 10.6151
R1084 B.n456 B.n455 10.6151
R1085 B.n455 B.n95 10.6151
R1086 B.n449 B.n95 10.6151
R1087 B.n264 B.n263 9.36635
R1088 B.n241 B.n177 9.36635
R1089 B.n76 B.n72 9.36635
R1090 B.n504 B.n503 9.36635
R1091 B.n642 B.n0 8.11757
R1092 B.n642 B.n1 8.11757
R1093 B.t3 B.n133 7.14046
R1094 B.n597 B.t10 7.14046
R1095 B.n263 B.n262 1.24928
R1096 B.n245 B.n177 1.24928
R1097 B.n522 B.n76 1.24928
R1098 B.n505 B.n504 1.24928
R1099 VP.n0 VP.t1 130.851
R1100 VP.n0 VP.t0 87.6115
R1101 VP VP.n0 0.52637
R1102 VTAIL.n1 VTAIL.t0 51.1591
R1103 VTAIL.n3 VTAIL.t1 51.1589
R1104 VTAIL.n0 VTAIL.t2 51.1589
R1105 VTAIL.n2 VTAIL.t3 51.1589
R1106 VTAIL.n1 VTAIL.n0 25.0134
R1107 VTAIL.n3 VTAIL.n2 21.7289
R1108 VTAIL.n2 VTAIL.n1 2.11257
R1109 VTAIL VTAIL.n0 1.34964
R1110 VTAIL VTAIL.n3 0.763431
R1111 VDD1 VDD1.t1 105.49
R1112 VDD1 VDD1.t0 68.717
R1113 VN VN.t1 130.758
R1114 VN VN.t0 88.1374
R1115 VDD2.n0 VDD2.t1 104.144
R1116 VDD2.n0 VDD2.t0 67.8377
R1117 VDD2 VDD2.n0 0.87981
C0 VTAIL VDD2 4.0458f
C1 VDD1 VDD2 0.781677f
C2 VTAIL VDD1 3.98768f
C3 VN VP 4.95104f
C4 VP VDD2 0.369731f
C5 VTAIL VP 1.87263f
C6 VP VDD1 2.02291f
C7 VN VDD2 1.80321f
C8 VTAIL VN 1.85845f
C9 VN VDD1 0.148526f
C10 VDD2 B 3.800073f
C11 VDD1 B 6.83915f
C12 VTAIL B 5.477263f
C13 VN B 9.02887f
C14 VP B 7.028025f
C15 VDD2.t1 B 1.17916f
C16 VDD2.t0 B 0.866734f
C17 VDD2.n0 B 1.83661f
C18 VN.t0 B 1.33272f
C19 VN.t1 B 1.7109f
C20 VDD1.t0 B 1.28681f
C21 VDD1.t1 B 1.78456f
C22 VTAIL.t2 B 0.906219f
C23 VTAIL.n0 B 1.13903f
C24 VTAIL.t0 B 0.906223f
C25 VTAIL.n1 B 1.17828f
C26 VTAIL.t3 B 0.906219f
C27 VTAIL.n2 B 1.00928f
C28 VTAIL.t1 B 0.906219f
C29 VTAIL.n3 B 0.939851f
C30 VP.t1 B 2.40619f
C31 VP.t0 B 1.87115f
C32 VP.n0 B 2.63537f
.ends

