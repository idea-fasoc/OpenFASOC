* NGSPICE file created from diff_pair_sample_0124.ext - technology: sky130A

.subckt diff_pair_sample_0124 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=3.0624 pd=18.89 as=3.0624 ps=18.89 w=18.56 l=2.47
X1 VDD1.t5 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.0624 pd=18.89 as=7.2384 ps=37.9 w=18.56 l=2.47
X2 VDD1.t4 VP.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.0624 pd=18.89 as=7.2384 ps=37.9 w=18.56 l=2.47
X3 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=7.2384 pd=37.9 as=0 ps=0 w=18.56 l=2.47
X4 VDD1.t3 VP.t2 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=7.2384 pd=37.9 as=3.0624 ps=18.89 w=18.56 l=2.47
X5 VDD2.t0 VN.t1 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=3.0624 pd=18.89 as=7.2384 ps=37.9 w=18.56 l=2.47
X6 VTAIL.t1 VP.t3 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=3.0624 pd=18.89 as=3.0624 ps=18.89 w=18.56 l=2.47
X7 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=7.2384 pd=37.9 as=0 ps=0 w=18.56 l=2.47
X8 VDD2.t1 VN.t2 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=3.0624 pd=18.89 as=7.2384 ps=37.9 w=18.56 l=2.47
X9 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.2384 pd=37.9 as=0 ps=0 w=18.56 l=2.47
X10 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.2384 pd=37.9 as=0 ps=0 w=18.56 l=2.47
X11 VTAIL.t8 VN.t3 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.0624 pd=18.89 as=3.0624 ps=18.89 w=18.56 l=2.47
X12 VTAIL.t0 VP.t4 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=3.0624 pd=18.89 as=3.0624 ps=18.89 w=18.56 l=2.47
X13 VDD2.t5 VN.t4 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=7.2384 pd=37.9 as=3.0624 ps=18.89 w=18.56 l=2.47
X14 VDD2.t4 VN.t5 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=7.2384 pd=37.9 as=3.0624 ps=18.89 w=18.56 l=2.47
X15 VDD1.t0 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=7.2384 pd=37.9 as=3.0624 ps=18.89 w=18.56 l=2.47
R0 VN.n3 VN.t5 216.238
R1 VN.n17 VN.t2 216.238
R2 VN.n4 VN.t0 181.093
R3 VN.n12 VN.t1 181.093
R4 VN.n18 VN.t3 181.093
R5 VN.n26 VN.t4 181.093
R6 VN.n25 VN.n14 161.3
R7 VN.n24 VN.n23 161.3
R8 VN.n22 VN.n15 161.3
R9 VN.n21 VN.n20 161.3
R10 VN.n19 VN.n16 161.3
R11 VN.n11 VN.n0 161.3
R12 VN.n10 VN.n9 161.3
R13 VN.n8 VN.n1 161.3
R14 VN.n7 VN.n6 161.3
R15 VN.n5 VN.n2 161.3
R16 VN.n13 VN.n12 96.1531
R17 VN.n27 VN.n26 96.1531
R18 VN VN.n27 53.4755
R19 VN.n6 VN.n1 50.2647
R20 VN.n20 VN.n15 50.2647
R21 VN.n4 VN.n3 48.1821
R22 VN.n18 VN.n17 48.1821
R23 VN.n10 VN.n1 30.8893
R24 VN.n24 VN.n15 30.8893
R25 VN.n5 VN.n4 24.5923
R26 VN.n6 VN.n5 24.5923
R27 VN.n11 VN.n10 24.5923
R28 VN.n20 VN.n19 24.5923
R29 VN.n19 VN.n18 24.5923
R30 VN.n25 VN.n24 24.5923
R31 VN.n12 VN.n11 14.7556
R32 VN.n26 VN.n25 14.7556
R33 VN.n17 VN.n16 6.50797
R34 VN.n3 VN.n2 6.50797
R35 VN.n27 VN.n14 0.278335
R36 VN.n13 VN.n0 0.278335
R37 VN.n23 VN.n14 0.189894
R38 VN.n23 VN.n22 0.189894
R39 VN.n22 VN.n21 0.189894
R40 VN.n21 VN.n16 0.189894
R41 VN.n7 VN.n2 0.189894
R42 VN.n8 VN.n7 0.189894
R43 VN.n9 VN.n8 0.189894
R44 VN.n9 VN.n0 0.189894
R45 VN VN.n13 0.153485
R46 VDD2.n1 VDD2.t4 62.6799
R47 VDD2.n2 VDD2.t5 60.9251
R48 VDD2.n1 VDD2.n0 60.4062
R49 VDD2 VDD2.n3 60.4034
R50 VDD2.n2 VDD2.n1 47.5601
R51 VDD2 VDD2.n2 1.86903
R52 VDD2.n3 VDD2.t3 1.06731
R53 VDD2.n3 VDD2.t1 1.06731
R54 VDD2.n0 VDD2.t2 1.06731
R55 VDD2.n0 VDD2.t0 1.06731
R56 VTAIL.n7 VTAIL.t9 44.2463
R57 VTAIL.n11 VTAIL.t10 44.2462
R58 VTAIL.n2 VTAIL.t2 44.2462
R59 VTAIL.n10 VTAIL.t4 44.2462
R60 VTAIL.n9 VTAIL.n8 43.1795
R61 VTAIL.n6 VTAIL.n5 43.1795
R62 VTAIL.n1 VTAIL.n0 43.1793
R63 VTAIL.n4 VTAIL.n3 43.1793
R64 VTAIL.n6 VTAIL.n4 33.1945
R65 VTAIL.n11 VTAIL.n10 30.7807
R66 VTAIL.n7 VTAIL.n6 2.41429
R67 VTAIL.n10 VTAIL.n9 2.41429
R68 VTAIL.n4 VTAIL.n2 2.41429
R69 VTAIL VTAIL.n11 1.75266
R70 VTAIL.n9 VTAIL.n7 1.67722
R71 VTAIL.n2 VTAIL.n1 1.67722
R72 VTAIL.n0 VTAIL.t6 1.06731
R73 VTAIL.n0 VTAIL.t11 1.06731
R74 VTAIL.n3 VTAIL.t5 1.06731
R75 VTAIL.n3 VTAIL.t1 1.06731
R76 VTAIL.n8 VTAIL.t3 1.06731
R77 VTAIL.n8 VTAIL.t0 1.06731
R78 VTAIL.n5 VTAIL.t7 1.06731
R79 VTAIL.n5 VTAIL.t8 1.06731
R80 VTAIL VTAIL.n1 0.662138
R81 B.n997 B.n996 585
R82 B.n998 B.n997 585
R83 B.n407 B.n142 585
R84 B.n406 B.n405 585
R85 B.n404 B.n403 585
R86 B.n402 B.n401 585
R87 B.n400 B.n399 585
R88 B.n398 B.n397 585
R89 B.n396 B.n395 585
R90 B.n394 B.n393 585
R91 B.n392 B.n391 585
R92 B.n390 B.n389 585
R93 B.n388 B.n387 585
R94 B.n386 B.n385 585
R95 B.n384 B.n383 585
R96 B.n382 B.n381 585
R97 B.n380 B.n379 585
R98 B.n378 B.n377 585
R99 B.n376 B.n375 585
R100 B.n374 B.n373 585
R101 B.n372 B.n371 585
R102 B.n370 B.n369 585
R103 B.n368 B.n367 585
R104 B.n366 B.n365 585
R105 B.n364 B.n363 585
R106 B.n362 B.n361 585
R107 B.n360 B.n359 585
R108 B.n358 B.n357 585
R109 B.n356 B.n355 585
R110 B.n354 B.n353 585
R111 B.n352 B.n351 585
R112 B.n350 B.n349 585
R113 B.n348 B.n347 585
R114 B.n346 B.n345 585
R115 B.n344 B.n343 585
R116 B.n342 B.n341 585
R117 B.n340 B.n339 585
R118 B.n338 B.n337 585
R119 B.n336 B.n335 585
R120 B.n334 B.n333 585
R121 B.n332 B.n331 585
R122 B.n330 B.n329 585
R123 B.n328 B.n327 585
R124 B.n326 B.n325 585
R125 B.n324 B.n323 585
R126 B.n322 B.n321 585
R127 B.n320 B.n319 585
R128 B.n318 B.n317 585
R129 B.n316 B.n315 585
R130 B.n314 B.n313 585
R131 B.n312 B.n311 585
R132 B.n310 B.n309 585
R133 B.n308 B.n307 585
R134 B.n306 B.n305 585
R135 B.n304 B.n303 585
R136 B.n302 B.n301 585
R137 B.n300 B.n299 585
R138 B.n298 B.n297 585
R139 B.n296 B.n295 585
R140 B.n294 B.n293 585
R141 B.n292 B.n291 585
R142 B.n290 B.n289 585
R143 B.n288 B.n287 585
R144 B.n286 B.n285 585
R145 B.n284 B.n283 585
R146 B.n282 B.n281 585
R147 B.n280 B.n279 585
R148 B.n278 B.n277 585
R149 B.n276 B.n275 585
R150 B.n274 B.n273 585
R151 B.n272 B.n271 585
R152 B.n269 B.n268 585
R153 B.n267 B.n266 585
R154 B.n265 B.n264 585
R155 B.n263 B.n262 585
R156 B.n261 B.n260 585
R157 B.n259 B.n258 585
R158 B.n257 B.n256 585
R159 B.n255 B.n254 585
R160 B.n253 B.n252 585
R161 B.n251 B.n250 585
R162 B.n249 B.n248 585
R163 B.n247 B.n246 585
R164 B.n245 B.n244 585
R165 B.n243 B.n242 585
R166 B.n241 B.n240 585
R167 B.n239 B.n238 585
R168 B.n237 B.n236 585
R169 B.n235 B.n234 585
R170 B.n233 B.n232 585
R171 B.n231 B.n230 585
R172 B.n229 B.n228 585
R173 B.n227 B.n226 585
R174 B.n225 B.n224 585
R175 B.n223 B.n222 585
R176 B.n221 B.n220 585
R177 B.n219 B.n218 585
R178 B.n217 B.n216 585
R179 B.n215 B.n214 585
R180 B.n213 B.n212 585
R181 B.n211 B.n210 585
R182 B.n209 B.n208 585
R183 B.n207 B.n206 585
R184 B.n205 B.n204 585
R185 B.n203 B.n202 585
R186 B.n201 B.n200 585
R187 B.n199 B.n198 585
R188 B.n197 B.n196 585
R189 B.n195 B.n194 585
R190 B.n193 B.n192 585
R191 B.n191 B.n190 585
R192 B.n189 B.n188 585
R193 B.n187 B.n186 585
R194 B.n185 B.n184 585
R195 B.n183 B.n182 585
R196 B.n181 B.n180 585
R197 B.n179 B.n178 585
R198 B.n177 B.n176 585
R199 B.n175 B.n174 585
R200 B.n173 B.n172 585
R201 B.n171 B.n170 585
R202 B.n169 B.n168 585
R203 B.n167 B.n166 585
R204 B.n165 B.n164 585
R205 B.n163 B.n162 585
R206 B.n161 B.n160 585
R207 B.n159 B.n158 585
R208 B.n157 B.n156 585
R209 B.n155 B.n154 585
R210 B.n153 B.n152 585
R211 B.n151 B.n150 585
R212 B.n149 B.n148 585
R213 B.n995 B.n76 585
R214 B.n999 B.n76 585
R215 B.n994 B.n75 585
R216 B.n1000 B.n75 585
R217 B.n993 B.n992 585
R218 B.n992 B.n71 585
R219 B.n991 B.n70 585
R220 B.n1006 B.n70 585
R221 B.n990 B.n69 585
R222 B.n1007 B.n69 585
R223 B.n989 B.n68 585
R224 B.n1008 B.n68 585
R225 B.n988 B.n987 585
R226 B.n987 B.n64 585
R227 B.n986 B.n63 585
R228 B.n1014 B.n63 585
R229 B.n985 B.n62 585
R230 B.n1015 B.n62 585
R231 B.n984 B.n61 585
R232 B.n1016 B.n61 585
R233 B.n983 B.n982 585
R234 B.n982 B.n57 585
R235 B.n981 B.n56 585
R236 B.n1022 B.n56 585
R237 B.n980 B.n55 585
R238 B.n1023 B.n55 585
R239 B.n979 B.n54 585
R240 B.n1024 B.n54 585
R241 B.n978 B.n977 585
R242 B.n977 B.n50 585
R243 B.n976 B.n49 585
R244 B.n1030 B.n49 585
R245 B.n975 B.n48 585
R246 B.n1031 B.n48 585
R247 B.n974 B.n47 585
R248 B.n1032 B.n47 585
R249 B.n973 B.n972 585
R250 B.n972 B.n46 585
R251 B.n971 B.n42 585
R252 B.n1038 B.n42 585
R253 B.n970 B.n41 585
R254 B.n1039 B.n41 585
R255 B.n969 B.n40 585
R256 B.n1040 B.n40 585
R257 B.n968 B.n967 585
R258 B.n967 B.n36 585
R259 B.n966 B.n35 585
R260 B.n1046 B.n35 585
R261 B.n965 B.n34 585
R262 B.n1047 B.n34 585
R263 B.n964 B.n33 585
R264 B.n1048 B.n33 585
R265 B.n963 B.n962 585
R266 B.n962 B.n29 585
R267 B.n961 B.n28 585
R268 B.n1054 B.n28 585
R269 B.n960 B.n27 585
R270 B.n1055 B.n27 585
R271 B.n959 B.n26 585
R272 B.n1056 B.n26 585
R273 B.n958 B.n957 585
R274 B.n957 B.n22 585
R275 B.n956 B.n21 585
R276 B.n1062 B.n21 585
R277 B.n955 B.n20 585
R278 B.n1063 B.n20 585
R279 B.n954 B.n19 585
R280 B.n1064 B.n19 585
R281 B.n953 B.n952 585
R282 B.n952 B.n15 585
R283 B.n951 B.n14 585
R284 B.n1070 B.n14 585
R285 B.n950 B.n13 585
R286 B.n1071 B.n13 585
R287 B.n949 B.n12 585
R288 B.n1072 B.n12 585
R289 B.n948 B.n947 585
R290 B.n947 B.n8 585
R291 B.n946 B.n7 585
R292 B.n1078 B.n7 585
R293 B.n945 B.n6 585
R294 B.n1079 B.n6 585
R295 B.n944 B.n5 585
R296 B.n1080 B.n5 585
R297 B.n943 B.n942 585
R298 B.n942 B.n4 585
R299 B.n941 B.n408 585
R300 B.n941 B.n940 585
R301 B.n931 B.n409 585
R302 B.n410 B.n409 585
R303 B.n933 B.n932 585
R304 B.n934 B.n933 585
R305 B.n930 B.n415 585
R306 B.n415 B.n414 585
R307 B.n929 B.n928 585
R308 B.n928 B.n927 585
R309 B.n417 B.n416 585
R310 B.n418 B.n417 585
R311 B.n920 B.n919 585
R312 B.n921 B.n920 585
R313 B.n918 B.n423 585
R314 B.n423 B.n422 585
R315 B.n917 B.n916 585
R316 B.n916 B.n915 585
R317 B.n425 B.n424 585
R318 B.n426 B.n425 585
R319 B.n908 B.n907 585
R320 B.n909 B.n908 585
R321 B.n906 B.n431 585
R322 B.n431 B.n430 585
R323 B.n905 B.n904 585
R324 B.n904 B.n903 585
R325 B.n433 B.n432 585
R326 B.n434 B.n433 585
R327 B.n896 B.n895 585
R328 B.n897 B.n896 585
R329 B.n894 B.n439 585
R330 B.n439 B.n438 585
R331 B.n893 B.n892 585
R332 B.n892 B.n891 585
R333 B.n441 B.n440 585
R334 B.n442 B.n441 585
R335 B.n884 B.n883 585
R336 B.n885 B.n884 585
R337 B.n882 B.n447 585
R338 B.n447 B.n446 585
R339 B.n881 B.n880 585
R340 B.n880 B.n879 585
R341 B.n449 B.n448 585
R342 B.n872 B.n449 585
R343 B.n871 B.n870 585
R344 B.n873 B.n871 585
R345 B.n869 B.n454 585
R346 B.n454 B.n453 585
R347 B.n868 B.n867 585
R348 B.n867 B.n866 585
R349 B.n456 B.n455 585
R350 B.n457 B.n456 585
R351 B.n859 B.n858 585
R352 B.n860 B.n859 585
R353 B.n857 B.n462 585
R354 B.n462 B.n461 585
R355 B.n856 B.n855 585
R356 B.n855 B.n854 585
R357 B.n464 B.n463 585
R358 B.n465 B.n464 585
R359 B.n847 B.n846 585
R360 B.n848 B.n847 585
R361 B.n845 B.n470 585
R362 B.n470 B.n469 585
R363 B.n844 B.n843 585
R364 B.n843 B.n842 585
R365 B.n472 B.n471 585
R366 B.n473 B.n472 585
R367 B.n835 B.n834 585
R368 B.n836 B.n835 585
R369 B.n833 B.n478 585
R370 B.n478 B.n477 585
R371 B.n832 B.n831 585
R372 B.n831 B.n830 585
R373 B.n480 B.n479 585
R374 B.n481 B.n480 585
R375 B.n823 B.n822 585
R376 B.n824 B.n823 585
R377 B.n821 B.n486 585
R378 B.n486 B.n485 585
R379 B.n815 B.n814 585
R380 B.n813 B.n553 585
R381 B.n812 B.n552 585
R382 B.n817 B.n552 585
R383 B.n811 B.n810 585
R384 B.n809 B.n808 585
R385 B.n807 B.n806 585
R386 B.n805 B.n804 585
R387 B.n803 B.n802 585
R388 B.n801 B.n800 585
R389 B.n799 B.n798 585
R390 B.n797 B.n796 585
R391 B.n795 B.n794 585
R392 B.n793 B.n792 585
R393 B.n791 B.n790 585
R394 B.n789 B.n788 585
R395 B.n787 B.n786 585
R396 B.n785 B.n784 585
R397 B.n783 B.n782 585
R398 B.n781 B.n780 585
R399 B.n779 B.n778 585
R400 B.n777 B.n776 585
R401 B.n775 B.n774 585
R402 B.n773 B.n772 585
R403 B.n771 B.n770 585
R404 B.n769 B.n768 585
R405 B.n767 B.n766 585
R406 B.n765 B.n764 585
R407 B.n763 B.n762 585
R408 B.n761 B.n760 585
R409 B.n759 B.n758 585
R410 B.n757 B.n756 585
R411 B.n755 B.n754 585
R412 B.n753 B.n752 585
R413 B.n751 B.n750 585
R414 B.n749 B.n748 585
R415 B.n747 B.n746 585
R416 B.n745 B.n744 585
R417 B.n743 B.n742 585
R418 B.n741 B.n740 585
R419 B.n739 B.n738 585
R420 B.n737 B.n736 585
R421 B.n735 B.n734 585
R422 B.n733 B.n732 585
R423 B.n731 B.n730 585
R424 B.n729 B.n728 585
R425 B.n727 B.n726 585
R426 B.n725 B.n724 585
R427 B.n723 B.n722 585
R428 B.n721 B.n720 585
R429 B.n719 B.n718 585
R430 B.n717 B.n716 585
R431 B.n715 B.n714 585
R432 B.n713 B.n712 585
R433 B.n711 B.n710 585
R434 B.n709 B.n708 585
R435 B.n707 B.n706 585
R436 B.n705 B.n704 585
R437 B.n703 B.n702 585
R438 B.n701 B.n700 585
R439 B.n699 B.n698 585
R440 B.n697 B.n696 585
R441 B.n695 B.n694 585
R442 B.n693 B.n692 585
R443 B.n691 B.n690 585
R444 B.n689 B.n688 585
R445 B.n687 B.n686 585
R446 B.n685 B.n684 585
R447 B.n683 B.n682 585
R448 B.n681 B.n680 585
R449 B.n679 B.n678 585
R450 B.n676 B.n675 585
R451 B.n674 B.n673 585
R452 B.n672 B.n671 585
R453 B.n670 B.n669 585
R454 B.n668 B.n667 585
R455 B.n666 B.n665 585
R456 B.n664 B.n663 585
R457 B.n662 B.n661 585
R458 B.n660 B.n659 585
R459 B.n658 B.n657 585
R460 B.n656 B.n655 585
R461 B.n654 B.n653 585
R462 B.n652 B.n651 585
R463 B.n650 B.n649 585
R464 B.n648 B.n647 585
R465 B.n646 B.n645 585
R466 B.n644 B.n643 585
R467 B.n642 B.n641 585
R468 B.n640 B.n639 585
R469 B.n638 B.n637 585
R470 B.n636 B.n635 585
R471 B.n634 B.n633 585
R472 B.n632 B.n631 585
R473 B.n630 B.n629 585
R474 B.n628 B.n627 585
R475 B.n626 B.n625 585
R476 B.n624 B.n623 585
R477 B.n622 B.n621 585
R478 B.n620 B.n619 585
R479 B.n618 B.n617 585
R480 B.n616 B.n615 585
R481 B.n614 B.n613 585
R482 B.n612 B.n611 585
R483 B.n610 B.n609 585
R484 B.n608 B.n607 585
R485 B.n606 B.n605 585
R486 B.n604 B.n603 585
R487 B.n602 B.n601 585
R488 B.n600 B.n599 585
R489 B.n598 B.n597 585
R490 B.n596 B.n595 585
R491 B.n594 B.n593 585
R492 B.n592 B.n591 585
R493 B.n590 B.n589 585
R494 B.n588 B.n587 585
R495 B.n586 B.n585 585
R496 B.n584 B.n583 585
R497 B.n582 B.n581 585
R498 B.n580 B.n579 585
R499 B.n578 B.n577 585
R500 B.n576 B.n575 585
R501 B.n574 B.n573 585
R502 B.n572 B.n571 585
R503 B.n570 B.n569 585
R504 B.n568 B.n567 585
R505 B.n566 B.n565 585
R506 B.n564 B.n563 585
R507 B.n562 B.n561 585
R508 B.n560 B.n559 585
R509 B.n488 B.n487 585
R510 B.n820 B.n819 585
R511 B.n484 B.n483 585
R512 B.n485 B.n484 585
R513 B.n826 B.n825 585
R514 B.n825 B.n824 585
R515 B.n827 B.n482 585
R516 B.n482 B.n481 585
R517 B.n829 B.n828 585
R518 B.n830 B.n829 585
R519 B.n476 B.n475 585
R520 B.n477 B.n476 585
R521 B.n838 B.n837 585
R522 B.n837 B.n836 585
R523 B.n839 B.n474 585
R524 B.n474 B.n473 585
R525 B.n841 B.n840 585
R526 B.n842 B.n841 585
R527 B.n468 B.n467 585
R528 B.n469 B.n468 585
R529 B.n850 B.n849 585
R530 B.n849 B.n848 585
R531 B.n851 B.n466 585
R532 B.n466 B.n465 585
R533 B.n853 B.n852 585
R534 B.n854 B.n853 585
R535 B.n460 B.n459 585
R536 B.n461 B.n460 585
R537 B.n862 B.n861 585
R538 B.n861 B.n860 585
R539 B.n863 B.n458 585
R540 B.n458 B.n457 585
R541 B.n865 B.n864 585
R542 B.n866 B.n865 585
R543 B.n452 B.n451 585
R544 B.n453 B.n452 585
R545 B.n875 B.n874 585
R546 B.n874 B.n873 585
R547 B.n876 B.n450 585
R548 B.n872 B.n450 585
R549 B.n878 B.n877 585
R550 B.n879 B.n878 585
R551 B.n445 B.n444 585
R552 B.n446 B.n445 585
R553 B.n887 B.n886 585
R554 B.n886 B.n885 585
R555 B.n888 B.n443 585
R556 B.n443 B.n442 585
R557 B.n890 B.n889 585
R558 B.n891 B.n890 585
R559 B.n437 B.n436 585
R560 B.n438 B.n437 585
R561 B.n899 B.n898 585
R562 B.n898 B.n897 585
R563 B.n900 B.n435 585
R564 B.n435 B.n434 585
R565 B.n902 B.n901 585
R566 B.n903 B.n902 585
R567 B.n429 B.n428 585
R568 B.n430 B.n429 585
R569 B.n911 B.n910 585
R570 B.n910 B.n909 585
R571 B.n912 B.n427 585
R572 B.n427 B.n426 585
R573 B.n914 B.n913 585
R574 B.n915 B.n914 585
R575 B.n421 B.n420 585
R576 B.n422 B.n421 585
R577 B.n923 B.n922 585
R578 B.n922 B.n921 585
R579 B.n924 B.n419 585
R580 B.n419 B.n418 585
R581 B.n926 B.n925 585
R582 B.n927 B.n926 585
R583 B.n413 B.n412 585
R584 B.n414 B.n413 585
R585 B.n936 B.n935 585
R586 B.n935 B.n934 585
R587 B.n937 B.n411 585
R588 B.n411 B.n410 585
R589 B.n939 B.n938 585
R590 B.n940 B.n939 585
R591 B.n2 B.n0 585
R592 B.n4 B.n2 585
R593 B.n3 B.n1 585
R594 B.n1079 B.n3 585
R595 B.n1077 B.n1076 585
R596 B.n1078 B.n1077 585
R597 B.n1075 B.n9 585
R598 B.n9 B.n8 585
R599 B.n1074 B.n1073 585
R600 B.n1073 B.n1072 585
R601 B.n11 B.n10 585
R602 B.n1071 B.n11 585
R603 B.n1069 B.n1068 585
R604 B.n1070 B.n1069 585
R605 B.n1067 B.n16 585
R606 B.n16 B.n15 585
R607 B.n1066 B.n1065 585
R608 B.n1065 B.n1064 585
R609 B.n18 B.n17 585
R610 B.n1063 B.n18 585
R611 B.n1061 B.n1060 585
R612 B.n1062 B.n1061 585
R613 B.n1059 B.n23 585
R614 B.n23 B.n22 585
R615 B.n1058 B.n1057 585
R616 B.n1057 B.n1056 585
R617 B.n25 B.n24 585
R618 B.n1055 B.n25 585
R619 B.n1053 B.n1052 585
R620 B.n1054 B.n1053 585
R621 B.n1051 B.n30 585
R622 B.n30 B.n29 585
R623 B.n1050 B.n1049 585
R624 B.n1049 B.n1048 585
R625 B.n32 B.n31 585
R626 B.n1047 B.n32 585
R627 B.n1045 B.n1044 585
R628 B.n1046 B.n1045 585
R629 B.n1043 B.n37 585
R630 B.n37 B.n36 585
R631 B.n1042 B.n1041 585
R632 B.n1041 B.n1040 585
R633 B.n39 B.n38 585
R634 B.n1039 B.n39 585
R635 B.n1037 B.n1036 585
R636 B.n1038 B.n1037 585
R637 B.n1035 B.n43 585
R638 B.n46 B.n43 585
R639 B.n1034 B.n1033 585
R640 B.n1033 B.n1032 585
R641 B.n45 B.n44 585
R642 B.n1031 B.n45 585
R643 B.n1029 B.n1028 585
R644 B.n1030 B.n1029 585
R645 B.n1027 B.n51 585
R646 B.n51 B.n50 585
R647 B.n1026 B.n1025 585
R648 B.n1025 B.n1024 585
R649 B.n53 B.n52 585
R650 B.n1023 B.n53 585
R651 B.n1021 B.n1020 585
R652 B.n1022 B.n1021 585
R653 B.n1019 B.n58 585
R654 B.n58 B.n57 585
R655 B.n1018 B.n1017 585
R656 B.n1017 B.n1016 585
R657 B.n60 B.n59 585
R658 B.n1015 B.n60 585
R659 B.n1013 B.n1012 585
R660 B.n1014 B.n1013 585
R661 B.n1011 B.n65 585
R662 B.n65 B.n64 585
R663 B.n1010 B.n1009 585
R664 B.n1009 B.n1008 585
R665 B.n67 B.n66 585
R666 B.n1007 B.n67 585
R667 B.n1005 B.n1004 585
R668 B.n1006 B.n1005 585
R669 B.n1003 B.n72 585
R670 B.n72 B.n71 585
R671 B.n1002 B.n1001 585
R672 B.n1001 B.n1000 585
R673 B.n74 B.n73 585
R674 B.n999 B.n74 585
R675 B.n1082 B.n1081 585
R676 B.n1081 B.n1080 585
R677 B.n815 B.n484 540.549
R678 B.n148 B.n74 540.549
R679 B.n819 B.n486 540.549
R680 B.n997 B.n76 540.549
R681 B.n557 B.t10 388.933
R682 B.n554 B.t17 388.933
R683 B.n146 B.t14 388.933
R684 B.n143 B.t6 388.933
R685 B.n998 B.n141 256.663
R686 B.n998 B.n140 256.663
R687 B.n998 B.n139 256.663
R688 B.n998 B.n138 256.663
R689 B.n998 B.n137 256.663
R690 B.n998 B.n136 256.663
R691 B.n998 B.n135 256.663
R692 B.n998 B.n134 256.663
R693 B.n998 B.n133 256.663
R694 B.n998 B.n132 256.663
R695 B.n998 B.n131 256.663
R696 B.n998 B.n130 256.663
R697 B.n998 B.n129 256.663
R698 B.n998 B.n128 256.663
R699 B.n998 B.n127 256.663
R700 B.n998 B.n126 256.663
R701 B.n998 B.n125 256.663
R702 B.n998 B.n124 256.663
R703 B.n998 B.n123 256.663
R704 B.n998 B.n122 256.663
R705 B.n998 B.n121 256.663
R706 B.n998 B.n120 256.663
R707 B.n998 B.n119 256.663
R708 B.n998 B.n118 256.663
R709 B.n998 B.n117 256.663
R710 B.n998 B.n116 256.663
R711 B.n998 B.n115 256.663
R712 B.n998 B.n114 256.663
R713 B.n998 B.n113 256.663
R714 B.n998 B.n112 256.663
R715 B.n998 B.n111 256.663
R716 B.n998 B.n110 256.663
R717 B.n998 B.n109 256.663
R718 B.n998 B.n108 256.663
R719 B.n998 B.n107 256.663
R720 B.n998 B.n106 256.663
R721 B.n998 B.n105 256.663
R722 B.n998 B.n104 256.663
R723 B.n998 B.n103 256.663
R724 B.n998 B.n102 256.663
R725 B.n998 B.n101 256.663
R726 B.n998 B.n100 256.663
R727 B.n998 B.n99 256.663
R728 B.n998 B.n98 256.663
R729 B.n998 B.n97 256.663
R730 B.n998 B.n96 256.663
R731 B.n998 B.n95 256.663
R732 B.n998 B.n94 256.663
R733 B.n998 B.n93 256.663
R734 B.n998 B.n92 256.663
R735 B.n998 B.n91 256.663
R736 B.n998 B.n90 256.663
R737 B.n998 B.n89 256.663
R738 B.n998 B.n88 256.663
R739 B.n998 B.n87 256.663
R740 B.n998 B.n86 256.663
R741 B.n998 B.n85 256.663
R742 B.n998 B.n84 256.663
R743 B.n998 B.n83 256.663
R744 B.n998 B.n82 256.663
R745 B.n998 B.n81 256.663
R746 B.n998 B.n80 256.663
R747 B.n998 B.n79 256.663
R748 B.n998 B.n78 256.663
R749 B.n998 B.n77 256.663
R750 B.n817 B.n816 256.663
R751 B.n817 B.n489 256.663
R752 B.n817 B.n490 256.663
R753 B.n817 B.n491 256.663
R754 B.n817 B.n492 256.663
R755 B.n817 B.n493 256.663
R756 B.n817 B.n494 256.663
R757 B.n817 B.n495 256.663
R758 B.n817 B.n496 256.663
R759 B.n817 B.n497 256.663
R760 B.n817 B.n498 256.663
R761 B.n817 B.n499 256.663
R762 B.n817 B.n500 256.663
R763 B.n817 B.n501 256.663
R764 B.n817 B.n502 256.663
R765 B.n817 B.n503 256.663
R766 B.n817 B.n504 256.663
R767 B.n817 B.n505 256.663
R768 B.n817 B.n506 256.663
R769 B.n817 B.n507 256.663
R770 B.n817 B.n508 256.663
R771 B.n817 B.n509 256.663
R772 B.n817 B.n510 256.663
R773 B.n817 B.n511 256.663
R774 B.n817 B.n512 256.663
R775 B.n817 B.n513 256.663
R776 B.n817 B.n514 256.663
R777 B.n817 B.n515 256.663
R778 B.n817 B.n516 256.663
R779 B.n817 B.n517 256.663
R780 B.n817 B.n518 256.663
R781 B.n817 B.n519 256.663
R782 B.n817 B.n520 256.663
R783 B.n817 B.n521 256.663
R784 B.n817 B.n522 256.663
R785 B.n817 B.n523 256.663
R786 B.n817 B.n524 256.663
R787 B.n817 B.n525 256.663
R788 B.n817 B.n526 256.663
R789 B.n817 B.n527 256.663
R790 B.n817 B.n528 256.663
R791 B.n817 B.n529 256.663
R792 B.n817 B.n530 256.663
R793 B.n817 B.n531 256.663
R794 B.n817 B.n532 256.663
R795 B.n817 B.n533 256.663
R796 B.n817 B.n534 256.663
R797 B.n817 B.n535 256.663
R798 B.n817 B.n536 256.663
R799 B.n817 B.n537 256.663
R800 B.n817 B.n538 256.663
R801 B.n817 B.n539 256.663
R802 B.n817 B.n540 256.663
R803 B.n817 B.n541 256.663
R804 B.n817 B.n542 256.663
R805 B.n817 B.n543 256.663
R806 B.n817 B.n544 256.663
R807 B.n817 B.n545 256.663
R808 B.n817 B.n546 256.663
R809 B.n817 B.n547 256.663
R810 B.n817 B.n548 256.663
R811 B.n817 B.n549 256.663
R812 B.n817 B.n550 256.663
R813 B.n817 B.n551 256.663
R814 B.n818 B.n817 256.663
R815 B.n825 B.n484 163.367
R816 B.n825 B.n482 163.367
R817 B.n829 B.n482 163.367
R818 B.n829 B.n476 163.367
R819 B.n837 B.n476 163.367
R820 B.n837 B.n474 163.367
R821 B.n841 B.n474 163.367
R822 B.n841 B.n468 163.367
R823 B.n849 B.n468 163.367
R824 B.n849 B.n466 163.367
R825 B.n853 B.n466 163.367
R826 B.n853 B.n460 163.367
R827 B.n861 B.n460 163.367
R828 B.n861 B.n458 163.367
R829 B.n865 B.n458 163.367
R830 B.n865 B.n452 163.367
R831 B.n874 B.n452 163.367
R832 B.n874 B.n450 163.367
R833 B.n878 B.n450 163.367
R834 B.n878 B.n445 163.367
R835 B.n886 B.n445 163.367
R836 B.n886 B.n443 163.367
R837 B.n890 B.n443 163.367
R838 B.n890 B.n437 163.367
R839 B.n898 B.n437 163.367
R840 B.n898 B.n435 163.367
R841 B.n902 B.n435 163.367
R842 B.n902 B.n429 163.367
R843 B.n910 B.n429 163.367
R844 B.n910 B.n427 163.367
R845 B.n914 B.n427 163.367
R846 B.n914 B.n421 163.367
R847 B.n922 B.n421 163.367
R848 B.n922 B.n419 163.367
R849 B.n926 B.n419 163.367
R850 B.n926 B.n413 163.367
R851 B.n935 B.n413 163.367
R852 B.n935 B.n411 163.367
R853 B.n939 B.n411 163.367
R854 B.n939 B.n2 163.367
R855 B.n1081 B.n2 163.367
R856 B.n1081 B.n3 163.367
R857 B.n1077 B.n3 163.367
R858 B.n1077 B.n9 163.367
R859 B.n1073 B.n9 163.367
R860 B.n1073 B.n11 163.367
R861 B.n1069 B.n11 163.367
R862 B.n1069 B.n16 163.367
R863 B.n1065 B.n16 163.367
R864 B.n1065 B.n18 163.367
R865 B.n1061 B.n18 163.367
R866 B.n1061 B.n23 163.367
R867 B.n1057 B.n23 163.367
R868 B.n1057 B.n25 163.367
R869 B.n1053 B.n25 163.367
R870 B.n1053 B.n30 163.367
R871 B.n1049 B.n30 163.367
R872 B.n1049 B.n32 163.367
R873 B.n1045 B.n32 163.367
R874 B.n1045 B.n37 163.367
R875 B.n1041 B.n37 163.367
R876 B.n1041 B.n39 163.367
R877 B.n1037 B.n39 163.367
R878 B.n1037 B.n43 163.367
R879 B.n1033 B.n43 163.367
R880 B.n1033 B.n45 163.367
R881 B.n1029 B.n45 163.367
R882 B.n1029 B.n51 163.367
R883 B.n1025 B.n51 163.367
R884 B.n1025 B.n53 163.367
R885 B.n1021 B.n53 163.367
R886 B.n1021 B.n58 163.367
R887 B.n1017 B.n58 163.367
R888 B.n1017 B.n60 163.367
R889 B.n1013 B.n60 163.367
R890 B.n1013 B.n65 163.367
R891 B.n1009 B.n65 163.367
R892 B.n1009 B.n67 163.367
R893 B.n1005 B.n67 163.367
R894 B.n1005 B.n72 163.367
R895 B.n1001 B.n72 163.367
R896 B.n1001 B.n74 163.367
R897 B.n553 B.n552 163.367
R898 B.n810 B.n552 163.367
R899 B.n808 B.n807 163.367
R900 B.n804 B.n803 163.367
R901 B.n800 B.n799 163.367
R902 B.n796 B.n795 163.367
R903 B.n792 B.n791 163.367
R904 B.n788 B.n787 163.367
R905 B.n784 B.n783 163.367
R906 B.n780 B.n779 163.367
R907 B.n776 B.n775 163.367
R908 B.n772 B.n771 163.367
R909 B.n768 B.n767 163.367
R910 B.n764 B.n763 163.367
R911 B.n760 B.n759 163.367
R912 B.n756 B.n755 163.367
R913 B.n752 B.n751 163.367
R914 B.n748 B.n747 163.367
R915 B.n744 B.n743 163.367
R916 B.n740 B.n739 163.367
R917 B.n736 B.n735 163.367
R918 B.n732 B.n731 163.367
R919 B.n728 B.n727 163.367
R920 B.n724 B.n723 163.367
R921 B.n720 B.n719 163.367
R922 B.n716 B.n715 163.367
R923 B.n712 B.n711 163.367
R924 B.n708 B.n707 163.367
R925 B.n704 B.n703 163.367
R926 B.n700 B.n699 163.367
R927 B.n696 B.n695 163.367
R928 B.n692 B.n691 163.367
R929 B.n688 B.n687 163.367
R930 B.n684 B.n683 163.367
R931 B.n680 B.n679 163.367
R932 B.n675 B.n674 163.367
R933 B.n671 B.n670 163.367
R934 B.n667 B.n666 163.367
R935 B.n663 B.n662 163.367
R936 B.n659 B.n658 163.367
R937 B.n655 B.n654 163.367
R938 B.n651 B.n650 163.367
R939 B.n647 B.n646 163.367
R940 B.n643 B.n642 163.367
R941 B.n639 B.n638 163.367
R942 B.n635 B.n634 163.367
R943 B.n631 B.n630 163.367
R944 B.n627 B.n626 163.367
R945 B.n623 B.n622 163.367
R946 B.n619 B.n618 163.367
R947 B.n615 B.n614 163.367
R948 B.n611 B.n610 163.367
R949 B.n607 B.n606 163.367
R950 B.n603 B.n602 163.367
R951 B.n599 B.n598 163.367
R952 B.n595 B.n594 163.367
R953 B.n591 B.n590 163.367
R954 B.n587 B.n586 163.367
R955 B.n583 B.n582 163.367
R956 B.n579 B.n578 163.367
R957 B.n575 B.n574 163.367
R958 B.n571 B.n570 163.367
R959 B.n567 B.n566 163.367
R960 B.n563 B.n562 163.367
R961 B.n559 B.n488 163.367
R962 B.n823 B.n486 163.367
R963 B.n823 B.n480 163.367
R964 B.n831 B.n480 163.367
R965 B.n831 B.n478 163.367
R966 B.n835 B.n478 163.367
R967 B.n835 B.n472 163.367
R968 B.n843 B.n472 163.367
R969 B.n843 B.n470 163.367
R970 B.n847 B.n470 163.367
R971 B.n847 B.n464 163.367
R972 B.n855 B.n464 163.367
R973 B.n855 B.n462 163.367
R974 B.n859 B.n462 163.367
R975 B.n859 B.n456 163.367
R976 B.n867 B.n456 163.367
R977 B.n867 B.n454 163.367
R978 B.n871 B.n454 163.367
R979 B.n871 B.n449 163.367
R980 B.n880 B.n449 163.367
R981 B.n880 B.n447 163.367
R982 B.n884 B.n447 163.367
R983 B.n884 B.n441 163.367
R984 B.n892 B.n441 163.367
R985 B.n892 B.n439 163.367
R986 B.n896 B.n439 163.367
R987 B.n896 B.n433 163.367
R988 B.n904 B.n433 163.367
R989 B.n904 B.n431 163.367
R990 B.n908 B.n431 163.367
R991 B.n908 B.n425 163.367
R992 B.n916 B.n425 163.367
R993 B.n916 B.n423 163.367
R994 B.n920 B.n423 163.367
R995 B.n920 B.n417 163.367
R996 B.n928 B.n417 163.367
R997 B.n928 B.n415 163.367
R998 B.n933 B.n415 163.367
R999 B.n933 B.n409 163.367
R1000 B.n941 B.n409 163.367
R1001 B.n942 B.n941 163.367
R1002 B.n942 B.n5 163.367
R1003 B.n6 B.n5 163.367
R1004 B.n7 B.n6 163.367
R1005 B.n947 B.n7 163.367
R1006 B.n947 B.n12 163.367
R1007 B.n13 B.n12 163.367
R1008 B.n14 B.n13 163.367
R1009 B.n952 B.n14 163.367
R1010 B.n952 B.n19 163.367
R1011 B.n20 B.n19 163.367
R1012 B.n21 B.n20 163.367
R1013 B.n957 B.n21 163.367
R1014 B.n957 B.n26 163.367
R1015 B.n27 B.n26 163.367
R1016 B.n28 B.n27 163.367
R1017 B.n962 B.n28 163.367
R1018 B.n962 B.n33 163.367
R1019 B.n34 B.n33 163.367
R1020 B.n35 B.n34 163.367
R1021 B.n967 B.n35 163.367
R1022 B.n967 B.n40 163.367
R1023 B.n41 B.n40 163.367
R1024 B.n42 B.n41 163.367
R1025 B.n972 B.n42 163.367
R1026 B.n972 B.n47 163.367
R1027 B.n48 B.n47 163.367
R1028 B.n49 B.n48 163.367
R1029 B.n977 B.n49 163.367
R1030 B.n977 B.n54 163.367
R1031 B.n55 B.n54 163.367
R1032 B.n56 B.n55 163.367
R1033 B.n982 B.n56 163.367
R1034 B.n982 B.n61 163.367
R1035 B.n62 B.n61 163.367
R1036 B.n63 B.n62 163.367
R1037 B.n987 B.n63 163.367
R1038 B.n987 B.n68 163.367
R1039 B.n69 B.n68 163.367
R1040 B.n70 B.n69 163.367
R1041 B.n992 B.n70 163.367
R1042 B.n992 B.n75 163.367
R1043 B.n76 B.n75 163.367
R1044 B.n152 B.n151 163.367
R1045 B.n156 B.n155 163.367
R1046 B.n160 B.n159 163.367
R1047 B.n164 B.n163 163.367
R1048 B.n168 B.n167 163.367
R1049 B.n172 B.n171 163.367
R1050 B.n176 B.n175 163.367
R1051 B.n180 B.n179 163.367
R1052 B.n184 B.n183 163.367
R1053 B.n188 B.n187 163.367
R1054 B.n192 B.n191 163.367
R1055 B.n196 B.n195 163.367
R1056 B.n200 B.n199 163.367
R1057 B.n204 B.n203 163.367
R1058 B.n208 B.n207 163.367
R1059 B.n212 B.n211 163.367
R1060 B.n216 B.n215 163.367
R1061 B.n220 B.n219 163.367
R1062 B.n224 B.n223 163.367
R1063 B.n228 B.n227 163.367
R1064 B.n232 B.n231 163.367
R1065 B.n236 B.n235 163.367
R1066 B.n240 B.n239 163.367
R1067 B.n244 B.n243 163.367
R1068 B.n248 B.n247 163.367
R1069 B.n252 B.n251 163.367
R1070 B.n256 B.n255 163.367
R1071 B.n260 B.n259 163.367
R1072 B.n264 B.n263 163.367
R1073 B.n268 B.n267 163.367
R1074 B.n273 B.n272 163.367
R1075 B.n277 B.n276 163.367
R1076 B.n281 B.n280 163.367
R1077 B.n285 B.n284 163.367
R1078 B.n289 B.n288 163.367
R1079 B.n293 B.n292 163.367
R1080 B.n297 B.n296 163.367
R1081 B.n301 B.n300 163.367
R1082 B.n305 B.n304 163.367
R1083 B.n309 B.n308 163.367
R1084 B.n313 B.n312 163.367
R1085 B.n317 B.n316 163.367
R1086 B.n321 B.n320 163.367
R1087 B.n325 B.n324 163.367
R1088 B.n329 B.n328 163.367
R1089 B.n333 B.n332 163.367
R1090 B.n337 B.n336 163.367
R1091 B.n341 B.n340 163.367
R1092 B.n345 B.n344 163.367
R1093 B.n349 B.n348 163.367
R1094 B.n353 B.n352 163.367
R1095 B.n357 B.n356 163.367
R1096 B.n361 B.n360 163.367
R1097 B.n365 B.n364 163.367
R1098 B.n369 B.n368 163.367
R1099 B.n373 B.n372 163.367
R1100 B.n377 B.n376 163.367
R1101 B.n381 B.n380 163.367
R1102 B.n385 B.n384 163.367
R1103 B.n389 B.n388 163.367
R1104 B.n393 B.n392 163.367
R1105 B.n397 B.n396 163.367
R1106 B.n401 B.n400 163.367
R1107 B.n405 B.n404 163.367
R1108 B.n997 B.n142 163.367
R1109 B.n557 B.t13 125.398
R1110 B.n143 B.t8 125.398
R1111 B.n554 B.t19 125.374
R1112 B.n146 B.t15 125.374
R1113 B.n816 B.n815 71.676
R1114 B.n810 B.n489 71.676
R1115 B.n807 B.n490 71.676
R1116 B.n803 B.n491 71.676
R1117 B.n799 B.n492 71.676
R1118 B.n795 B.n493 71.676
R1119 B.n791 B.n494 71.676
R1120 B.n787 B.n495 71.676
R1121 B.n783 B.n496 71.676
R1122 B.n779 B.n497 71.676
R1123 B.n775 B.n498 71.676
R1124 B.n771 B.n499 71.676
R1125 B.n767 B.n500 71.676
R1126 B.n763 B.n501 71.676
R1127 B.n759 B.n502 71.676
R1128 B.n755 B.n503 71.676
R1129 B.n751 B.n504 71.676
R1130 B.n747 B.n505 71.676
R1131 B.n743 B.n506 71.676
R1132 B.n739 B.n507 71.676
R1133 B.n735 B.n508 71.676
R1134 B.n731 B.n509 71.676
R1135 B.n727 B.n510 71.676
R1136 B.n723 B.n511 71.676
R1137 B.n719 B.n512 71.676
R1138 B.n715 B.n513 71.676
R1139 B.n711 B.n514 71.676
R1140 B.n707 B.n515 71.676
R1141 B.n703 B.n516 71.676
R1142 B.n699 B.n517 71.676
R1143 B.n695 B.n518 71.676
R1144 B.n691 B.n519 71.676
R1145 B.n687 B.n520 71.676
R1146 B.n683 B.n521 71.676
R1147 B.n679 B.n522 71.676
R1148 B.n674 B.n523 71.676
R1149 B.n670 B.n524 71.676
R1150 B.n666 B.n525 71.676
R1151 B.n662 B.n526 71.676
R1152 B.n658 B.n527 71.676
R1153 B.n654 B.n528 71.676
R1154 B.n650 B.n529 71.676
R1155 B.n646 B.n530 71.676
R1156 B.n642 B.n531 71.676
R1157 B.n638 B.n532 71.676
R1158 B.n634 B.n533 71.676
R1159 B.n630 B.n534 71.676
R1160 B.n626 B.n535 71.676
R1161 B.n622 B.n536 71.676
R1162 B.n618 B.n537 71.676
R1163 B.n614 B.n538 71.676
R1164 B.n610 B.n539 71.676
R1165 B.n606 B.n540 71.676
R1166 B.n602 B.n541 71.676
R1167 B.n598 B.n542 71.676
R1168 B.n594 B.n543 71.676
R1169 B.n590 B.n544 71.676
R1170 B.n586 B.n545 71.676
R1171 B.n582 B.n546 71.676
R1172 B.n578 B.n547 71.676
R1173 B.n574 B.n548 71.676
R1174 B.n570 B.n549 71.676
R1175 B.n566 B.n550 71.676
R1176 B.n562 B.n551 71.676
R1177 B.n818 B.n488 71.676
R1178 B.n148 B.n77 71.676
R1179 B.n152 B.n78 71.676
R1180 B.n156 B.n79 71.676
R1181 B.n160 B.n80 71.676
R1182 B.n164 B.n81 71.676
R1183 B.n168 B.n82 71.676
R1184 B.n172 B.n83 71.676
R1185 B.n176 B.n84 71.676
R1186 B.n180 B.n85 71.676
R1187 B.n184 B.n86 71.676
R1188 B.n188 B.n87 71.676
R1189 B.n192 B.n88 71.676
R1190 B.n196 B.n89 71.676
R1191 B.n200 B.n90 71.676
R1192 B.n204 B.n91 71.676
R1193 B.n208 B.n92 71.676
R1194 B.n212 B.n93 71.676
R1195 B.n216 B.n94 71.676
R1196 B.n220 B.n95 71.676
R1197 B.n224 B.n96 71.676
R1198 B.n228 B.n97 71.676
R1199 B.n232 B.n98 71.676
R1200 B.n236 B.n99 71.676
R1201 B.n240 B.n100 71.676
R1202 B.n244 B.n101 71.676
R1203 B.n248 B.n102 71.676
R1204 B.n252 B.n103 71.676
R1205 B.n256 B.n104 71.676
R1206 B.n260 B.n105 71.676
R1207 B.n264 B.n106 71.676
R1208 B.n268 B.n107 71.676
R1209 B.n273 B.n108 71.676
R1210 B.n277 B.n109 71.676
R1211 B.n281 B.n110 71.676
R1212 B.n285 B.n111 71.676
R1213 B.n289 B.n112 71.676
R1214 B.n293 B.n113 71.676
R1215 B.n297 B.n114 71.676
R1216 B.n301 B.n115 71.676
R1217 B.n305 B.n116 71.676
R1218 B.n309 B.n117 71.676
R1219 B.n313 B.n118 71.676
R1220 B.n317 B.n119 71.676
R1221 B.n321 B.n120 71.676
R1222 B.n325 B.n121 71.676
R1223 B.n329 B.n122 71.676
R1224 B.n333 B.n123 71.676
R1225 B.n337 B.n124 71.676
R1226 B.n341 B.n125 71.676
R1227 B.n345 B.n126 71.676
R1228 B.n349 B.n127 71.676
R1229 B.n353 B.n128 71.676
R1230 B.n357 B.n129 71.676
R1231 B.n361 B.n130 71.676
R1232 B.n365 B.n131 71.676
R1233 B.n369 B.n132 71.676
R1234 B.n373 B.n133 71.676
R1235 B.n377 B.n134 71.676
R1236 B.n381 B.n135 71.676
R1237 B.n385 B.n136 71.676
R1238 B.n389 B.n137 71.676
R1239 B.n393 B.n138 71.676
R1240 B.n397 B.n139 71.676
R1241 B.n401 B.n140 71.676
R1242 B.n405 B.n141 71.676
R1243 B.n142 B.n141 71.676
R1244 B.n404 B.n140 71.676
R1245 B.n400 B.n139 71.676
R1246 B.n396 B.n138 71.676
R1247 B.n392 B.n137 71.676
R1248 B.n388 B.n136 71.676
R1249 B.n384 B.n135 71.676
R1250 B.n380 B.n134 71.676
R1251 B.n376 B.n133 71.676
R1252 B.n372 B.n132 71.676
R1253 B.n368 B.n131 71.676
R1254 B.n364 B.n130 71.676
R1255 B.n360 B.n129 71.676
R1256 B.n356 B.n128 71.676
R1257 B.n352 B.n127 71.676
R1258 B.n348 B.n126 71.676
R1259 B.n344 B.n125 71.676
R1260 B.n340 B.n124 71.676
R1261 B.n336 B.n123 71.676
R1262 B.n332 B.n122 71.676
R1263 B.n328 B.n121 71.676
R1264 B.n324 B.n120 71.676
R1265 B.n320 B.n119 71.676
R1266 B.n316 B.n118 71.676
R1267 B.n312 B.n117 71.676
R1268 B.n308 B.n116 71.676
R1269 B.n304 B.n115 71.676
R1270 B.n300 B.n114 71.676
R1271 B.n296 B.n113 71.676
R1272 B.n292 B.n112 71.676
R1273 B.n288 B.n111 71.676
R1274 B.n284 B.n110 71.676
R1275 B.n280 B.n109 71.676
R1276 B.n276 B.n108 71.676
R1277 B.n272 B.n107 71.676
R1278 B.n267 B.n106 71.676
R1279 B.n263 B.n105 71.676
R1280 B.n259 B.n104 71.676
R1281 B.n255 B.n103 71.676
R1282 B.n251 B.n102 71.676
R1283 B.n247 B.n101 71.676
R1284 B.n243 B.n100 71.676
R1285 B.n239 B.n99 71.676
R1286 B.n235 B.n98 71.676
R1287 B.n231 B.n97 71.676
R1288 B.n227 B.n96 71.676
R1289 B.n223 B.n95 71.676
R1290 B.n219 B.n94 71.676
R1291 B.n215 B.n93 71.676
R1292 B.n211 B.n92 71.676
R1293 B.n207 B.n91 71.676
R1294 B.n203 B.n90 71.676
R1295 B.n199 B.n89 71.676
R1296 B.n195 B.n88 71.676
R1297 B.n191 B.n87 71.676
R1298 B.n187 B.n86 71.676
R1299 B.n183 B.n85 71.676
R1300 B.n179 B.n84 71.676
R1301 B.n175 B.n83 71.676
R1302 B.n171 B.n82 71.676
R1303 B.n167 B.n81 71.676
R1304 B.n163 B.n80 71.676
R1305 B.n159 B.n79 71.676
R1306 B.n155 B.n78 71.676
R1307 B.n151 B.n77 71.676
R1308 B.n816 B.n553 71.676
R1309 B.n808 B.n489 71.676
R1310 B.n804 B.n490 71.676
R1311 B.n800 B.n491 71.676
R1312 B.n796 B.n492 71.676
R1313 B.n792 B.n493 71.676
R1314 B.n788 B.n494 71.676
R1315 B.n784 B.n495 71.676
R1316 B.n780 B.n496 71.676
R1317 B.n776 B.n497 71.676
R1318 B.n772 B.n498 71.676
R1319 B.n768 B.n499 71.676
R1320 B.n764 B.n500 71.676
R1321 B.n760 B.n501 71.676
R1322 B.n756 B.n502 71.676
R1323 B.n752 B.n503 71.676
R1324 B.n748 B.n504 71.676
R1325 B.n744 B.n505 71.676
R1326 B.n740 B.n506 71.676
R1327 B.n736 B.n507 71.676
R1328 B.n732 B.n508 71.676
R1329 B.n728 B.n509 71.676
R1330 B.n724 B.n510 71.676
R1331 B.n720 B.n511 71.676
R1332 B.n716 B.n512 71.676
R1333 B.n712 B.n513 71.676
R1334 B.n708 B.n514 71.676
R1335 B.n704 B.n515 71.676
R1336 B.n700 B.n516 71.676
R1337 B.n696 B.n517 71.676
R1338 B.n692 B.n518 71.676
R1339 B.n688 B.n519 71.676
R1340 B.n684 B.n520 71.676
R1341 B.n680 B.n521 71.676
R1342 B.n675 B.n522 71.676
R1343 B.n671 B.n523 71.676
R1344 B.n667 B.n524 71.676
R1345 B.n663 B.n525 71.676
R1346 B.n659 B.n526 71.676
R1347 B.n655 B.n527 71.676
R1348 B.n651 B.n528 71.676
R1349 B.n647 B.n529 71.676
R1350 B.n643 B.n530 71.676
R1351 B.n639 B.n531 71.676
R1352 B.n635 B.n532 71.676
R1353 B.n631 B.n533 71.676
R1354 B.n627 B.n534 71.676
R1355 B.n623 B.n535 71.676
R1356 B.n619 B.n536 71.676
R1357 B.n615 B.n537 71.676
R1358 B.n611 B.n538 71.676
R1359 B.n607 B.n539 71.676
R1360 B.n603 B.n540 71.676
R1361 B.n599 B.n541 71.676
R1362 B.n595 B.n542 71.676
R1363 B.n591 B.n543 71.676
R1364 B.n587 B.n544 71.676
R1365 B.n583 B.n545 71.676
R1366 B.n579 B.n546 71.676
R1367 B.n575 B.n547 71.676
R1368 B.n571 B.n548 71.676
R1369 B.n567 B.n549 71.676
R1370 B.n563 B.n550 71.676
R1371 B.n559 B.n551 71.676
R1372 B.n819 B.n818 71.676
R1373 B.n558 B.t12 71.095
R1374 B.n144 B.t9 71.095
R1375 B.n555 B.t18 71.0703
R1376 B.n147 B.t16 71.0703
R1377 B.n677 B.n558 59.5399
R1378 B.n556 B.n555 59.5399
R1379 B.n270 B.n147 59.5399
R1380 B.n145 B.n144 59.5399
R1381 B.n817 B.n485 58.6118
R1382 B.n999 B.n998 58.6118
R1383 B.n558 B.n557 54.3035
R1384 B.n555 B.n554 54.3035
R1385 B.n147 B.n146 54.3035
R1386 B.n144 B.n143 54.3035
R1387 B.n149 B.n73 35.1225
R1388 B.n996 B.n995 35.1225
R1389 B.n821 B.n820 35.1225
R1390 B.n814 B.n483 35.1225
R1391 B.n824 B.n485 31.3829
R1392 B.n824 B.n481 31.3829
R1393 B.n830 B.n481 31.3829
R1394 B.n830 B.n477 31.3829
R1395 B.n836 B.n477 31.3829
R1396 B.n836 B.n473 31.3829
R1397 B.n842 B.n473 31.3829
R1398 B.n848 B.n469 31.3829
R1399 B.n848 B.n465 31.3829
R1400 B.n854 B.n465 31.3829
R1401 B.n854 B.n461 31.3829
R1402 B.n860 B.n461 31.3829
R1403 B.n860 B.n457 31.3829
R1404 B.n866 B.n457 31.3829
R1405 B.n866 B.n453 31.3829
R1406 B.n873 B.n453 31.3829
R1407 B.n873 B.n872 31.3829
R1408 B.n879 B.n446 31.3829
R1409 B.n885 B.n446 31.3829
R1410 B.n885 B.n442 31.3829
R1411 B.n891 B.n442 31.3829
R1412 B.n891 B.n438 31.3829
R1413 B.n897 B.n438 31.3829
R1414 B.n897 B.n434 31.3829
R1415 B.n903 B.n434 31.3829
R1416 B.n909 B.n430 31.3829
R1417 B.n909 B.n426 31.3829
R1418 B.n915 B.n426 31.3829
R1419 B.n915 B.n422 31.3829
R1420 B.n921 B.n422 31.3829
R1421 B.n921 B.n418 31.3829
R1422 B.n927 B.n418 31.3829
R1423 B.n934 B.n414 31.3829
R1424 B.n934 B.n410 31.3829
R1425 B.n940 B.n410 31.3829
R1426 B.n940 B.n4 31.3829
R1427 B.n1080 B.n4 31.3829
R1428 B.n1080 B.n1079 31.3829
R1429 B.n1079 B.n1078 31.3829
R1430 B.n1078 B.n8 31.3829
R1431 B.n1072 B.n8 31.3829
R1432 B.n1072 B.n1071 31.3829
R1433 B.n1070 B.n15 31.3829
R1434 B.n1064 B.n15 31.3829
R1435 B.n1064 B.n1063 31.3829
R1436 B.n1063 B.n1062 31.3829
R1437 B.n1062 B.n22 31.3829
R1438 B.n1056 B.n22 31.3829
R1439 B.n1056 B.n1055 31.3829
R1440 B.n1054 B.n29 31.3829
R1441 B.n1048 B.n29 31.3829
R1442 B.n1048 B.n1047 31.3829
R1443 B.n1047 B.n1046 31.3829
R1444 B.n1046 B.n36 31.3829
R1445 B.n1040 B.n36 31.3829
R1446 B.n1040 B.n1039 31.3829
R1447 B.n1039 B.n1038 31.3829
R1448 B.n1032 B.n46 31.3829
R1449 B.n1032 B.n1031 31.3829
R1450 B.n1031 B.n1030 31.3829
R1451 B.n1030 B.n50 31.3829
R1452 B.n1024 B.n50 31.3829
R1453 B.n1024 B.n1023 31.3829
R1454 B.n1023 B.n1022 31.3829
R1455 B.n1022 B.n57 31.3829
R1456 B.n1016 B.n57 31.3829
R1457 B.n1016 B.n1015 31.3829
R1458 B.n1014 B.n64 31.3829
R1459 B.n1008 B.n64 31.3829
R1460 B.n1008 B.n1007 31.3829
R1461 B.n1007 B.n1006 31.3829
R1462 B.n1006 B.n71 31.3829
R1463 B.n1000 B.n71 31.3829
R1464 B.n1000 B.n999 31.3829
R1465 B.t1 B.n430 29.9984
R1466 B.n1055 B.t0 29.9984
R1467 B.n872 B.t5 25.3833
R1468 B.n46 B.t4 25.3833
R1469 B.t2 B.n414 22.6143
R1470 B.n1071 B.t3 22.6143
R1471 B.t11 B.n469 19.8453
R1472 B.n1015 B.t7 19.8453
R1473 B B.n1082 18.0485
R1474 B.n842 B.t11 11.5382
R1475 B.t7 B.n1014 11.5382
R1476 B.n150 B.n149 10.6151
R1477 B.n153 B.n150 10.6151
R1478 B.n154 B.n153 10.6151
R1479 B.n157 B.n154 10.6151
R1480 B.n158 B.n157 10.6151
R1481 B.n161 B.n158 10.6151
R1482 B.n162 B.n161 10.6151
R1483 B.n165 B.n162 10.6151
R1484 B.n166 B.n165 10.6151
R1485 B.n169 B.n166 10.6151
R1486 B.n170 B.n169 10.6151
R1487 B.n173 B.n170 10.6151
R1488 B.n174 B.n173 10.6151
R1489 B.n177 B.n174 10.6151
R1490 B.n178 B.n177 10.6151
R1491 B.n181 B.n178 10.6151
R1492 B.n182 B.n181 10.6151
R1493 B.n185 B.n182 10.6151
R1494 B.n186 B.n185 10.6151
R1495 B.n189 B.n186 10.6151
R1496 B.n190 B.n189 10.6151
R1497 B.n193 B.n190 10.6151
R1498 B.n194 B.n193 10.6151
R1499 B.n197 B.n194 10.6151
R1500 B.n198 B.n197 10.6151
R1501 B.n201 B.n198 10.6151
R1502 B.n202 B.n201 10.6151
R1503 B.n205 B.n202 10.6151
R1504 B.n206 B.n205 10.6151
R1505 B.n209 B.n206 10.6151
R1506 B.n210 B.n209 10.6151
R1507 B.n213 B.n210 10.6151
R1508 B.n214 B.n213 10.6151
R1509 B.n217 B.n214 10.6151
R1510 B.n218 B.n217 10.6151
R1511 B.n221 B.n218 10.6151
R1512 B.n222 B.n221 10.6151
R1513 B.n225 B.n222 10.6151
R1514 B.n226 B.n225 10.6151
R1515 B.n229 B.n226 10.6151
R1516 B.n230 B.n229 10.6151
R1517 B.n233 B.n230 10.6151
R1518 B.n234 B.n233 10.6151
R1519 B.n237 B.n234 10.6151
R1520 B.n238 B.n237 10.6151
R1521 B.n241 B.n238 10.6151
R1522 B.n242 B.n241 10.6151
R1523 B.n245 B.n242 10.6151
R1524 B.n246 B.n245 10.6151
R1525 B.n249 B.n246 10.6151
R1526 B.n250 B.n249 10.6151
R1527 B.n253 B.n250 10.6151
R1528 B.n254 B.n253 10.6151
R1529 B.n257 B.n254 10.6151
R1530 B.n258 B.n257 10.6151
R1531 B.n261 B.n258 10.6151
R1532 B.n262 B.n261 10.6151
R1533 B.n265 B.n262 10.6151
R1534 B.n266 B.n265 10.6151
R1535 B.n269 B.n266 10.6151
R1536 B.n274 B.n271 10.6151
R1537 B.n275 B.n274 10.6151
R1538 B.n278 B.n275 10.6151
R1539 B.n279 B.n278 10.6151
R1540 B.n282 B.n279 10.6151
R1541 B.n283 B.n282 10.6151
R1542 B.n286 B.n283 10.6151
R1543 B.n287 B.n286 10.6151
R1544 B.n291 B.n290 10.6151
R1545 B.n294 B.n291 10.6151
R1546 B.n295 B.n294 10.6151
R1547 B.n298 B.n295 10.6151
R1548 B.n299 B.n298 10.6151
R1549 B.n302 B.n299 10.6151
R1550 B.n303 B.n302 10.6151
R1551 B.n306 B.n303 10.6151
R1552 B.n307 B.n306 10.6151
R1553 B.n310 B.n307 10.6151
R1554 B.n311 B.n310 10.6151
R1555 B.n314 B.n311 10.6151
R1556 B.n315 B.n314 10.6151
R1557 B.n318 B.n315 10.6151
R1558 B.n319 B.n318 10.6151
R1559 B.n322 B.n319 10.6151
R1560 B.n323 B.n322 10.6151
R1561 B.n326 B.n323 10.6151
R1562 B.n327 B.n326 10.6151
R1563 B.n330 B.n327 10.6151
R1564 B.n331 B.n330 10.6151
R1565 B.n334 B.n331 10.6151
R1566 B.n335 B.n334 10.6151
R1567 B.n338 B.n335 10.6151
R1568 B.n339 B.n338 10.6151
R1569 B.n342 B.n339 10.6151
R1570 B.n343 B.n342 10.6151
R1571 B.n346 B.n343 10.6151
R1572 B.n347 B.n346 10.6151
R1573 B.n350 B.n347 10.6151
R1574 B.n351 B.n350 10.6151
R1575 B.n354 B.n351 10.6151
R1576 B.n355 B.n354 10.6151
R1577 B.n358 B.n355 10.6151
R1578 B.n359 B.n358 10.6151
R1579 B.n362 B.n359 10.6151
R1580 B.n363 B.n362 10.6151
R1581 B.n366 B.n363 10.6151
R1582 B.n367 B.n366 10.6151
R1583 B.n370 B.n367 10.6151
R1584 B.n371 B.n370 10.6151
R1585 B.n374 B.n371 10.6151
R1586 B.n375 B.n374 10.6151
R1587 B.n378 B.n375 10.6151
R1588 B.n379 B.n378 10.6151
R1589 B.n382 B.n379 10.6151
R1590 B.n383 B.n382 10.6151
R1591 B.n386 B.n383 10.6151
R1592 B.n387 B.n386 10.6151
R1593 B.n390 B.n387 10.6151
R1594 B.n391 B.n390 10.6151
R1595 B.n394 B.n391 10.6151
R1596 B.n395 B.n394 10.6151
R1597 B.n398 B.n395 10.6151
R1598 B.n399 B.n398 10.6151
R1599 B.n402 B.n399 10.6151
R1600 B.n403 B.n402 10.6151
R1601 B.n406 B.n403 10.6151
R1602 B.n407 B.n406 10.6151
R1603 B.n996 B.n407 10.6151
R1604 B.n822 B.n821 10.6151
R1605 B.n822 B.n479 10.6151
R1606 B.n832 B.n479 10.6151
R1607 B.n833 B.n832 10.6151
R1608 B.n834 B.n833 10.6151
R1609 B.n834 B.n471 10.6151
R1610 B.n844 B.n471 10.6151
R1611 B.n845 B.n844 10.6151
R1612 B.n846 B.n845 10.6151
R1613 B.n846 B.n463 10.6151
R1614 B.n856 B.n463 10.6151
R1615 B.n857 B.n856 10.6151
R1616 B.n858 B.n857 10.6151
R1617 B.n858 B.n455 10.6151
R1618 B.n868 B.n455 10.6151
R1619 B.n869 B.n868 10.6151
R1620 B.n870 B.n869 10.6151
R1621 B.n870 B.n448 10.6151
R1622 B.n881 B.n448 10.6151
R1623 B.n882 B.n881 10.6151
R1624 B.n883 B.n882 10.6151
R1625 B.n883 B.n440 10.6151
R1626 B.n893 B.n440 10.6151
R1627 B.n894 B.n893 10.6151
R1628 B.n895 B.n894 10.6151
R1629 B.n895 B.n432 10.6151
R1630 B.n905 B.n432 10.6151
R1631 B.n906 B.n905 10.6151
R1632 B.n907 B.n906 10.6151
R1633 B.n907 B.n424 10.6151
R1634 B.n917 B.n424 10.6151
R1635 B.n918 B.n917 10.6151
R1636 B.n919 B.n918 10.6151
R1637 B.n919 B.n416 10.6151
R1638 B.n929 B.n416 10.6151
R1639 B.n930 B.n929 10.6151
R1640 B.n932 B.n930 10.6151
R1641 B.n932 B.n931 10.6151
R1642 B.n931 B.n408 10.6151
R1643 B.n943 B.n408 10.6151
R1644 B.n944 B.n943 10.6151
R1645 B.n945 B.n944 10.6151
R1646 B.n946 B.n945 10.6151
R1647 B.n948 B.n946 10.6151
R1648 B.n949 B.n948 10.6151
R1649 B.n950 B.n949 10.6151
R1650 B.n951 B.n950 10.6151
R1651 B.n953 B.n951 10.6151
R1652 B.n954 B.n953 10.6151
R1653 B.n955 B.n954 10.6151
R1654 B.n956 B.n955 10.6151
R1655 B.n958 B.n956 10.6151
R1656 B.n959 B.n958 10.6151
R1657 B.n960 B.n959 10.6151
R1658 B.n961 B.n960 10.6151
R1659 B.n963 B.n961 10.6151
R1660 B.n964 B.n963 10.6151
R1661 B.n965 B.n964 10.6151
R1662 B.n966 B.n965 10.6151
R1663 B.n968 B.n966 10.6151
R1664 B.n969 B.n968 10.6151
R1665 B.n970 B.n969 10.6151
R1666 B.n971 B.n970 10.6151
R1667 B.n973 B.n971 10.6151
R1668 B.n974 B.n973 10.6151
R1669 B.n975 B.n974 10.6151
R1670 B.n976 B.n975 10.6151
R1671 B.n978 B.n976 10.6151
R1672 B.n979 B.n978 10.6151
R1673 B.n980 B.n979 10.6151
R1674 B.n981 B.n980 10.6151
R1675 B.n983 B.n981 10.6151
R1676 B.n984 B.n983 10.6151
R1677 B.n985 B.n984 10.6151
R1678 B.n986 B.n985 10.6151
R1679 B.n988 B.n986 10.6151
R1680 B.n989 B.n988 10.6151
R1681 B.n990 B.n989 10.6151
R1682 B.n991 B.n990 10.6151
R1683 B.n993 B.n991 10.6151
R1684 B.n994 B.n993 10.6151
R1685 B.n995 B.n994 10.6151
R1686 B.n814 B.n813 10.6151
R1687 B.n813 B.n812 10.6151
R1688 B.n812 B.n811 10.6151
R1689 B.n811 B.n809 10.6151
R1690 B.n809 B.n806 10.6151
R1691 B.n806 B.n805 10.6151
R1692 B.n805 B.n802 10.6151
R1693 B.n802 B.n801 10.6151
R1694 B.n801 B.n798 10.6151
R1695 B.n798 B.n797 10.6151
R1696 B.n797 B.n794 10.6151
R1697 B.n794 B.n793 10.6151
R1698 B.n793 B.n790 10.6151
R1699 B.n790 B.n789 10.6151
R1700 B.n789 B.n786 10.6151
R1701 B.n786 B.n785 10.6151
R1702 B.n785 B.n782 10.6151
R1703 B.n782 B.n781 10.6151
R1704 B.n781 B.n778 10.6151
R1705 B.n778 B.n777 10.6151
R1706 B.n777 B.n774 10.6151
R1707 B.n774 B.n773 10.6151
R1708 B.n773 B.n770 10.6151
R1709 B.n770 B.n769 10.6151
R1710 B.n769 B.n766 10.6151
R1711 B.n766 B.n765 10.6151
R1712 B.n765 B.n762 10.6151
R1713 B.n762 B.n761 10.6151
R1714 B.n761 B.n758 10.6151
R1715 B.n758 B.n757 10.6151
R1716 B.n757 B.n754 10.6151
R1717 B.n754 B.n753 10.6151
R1718 B.n753 B.n750 10.6151
R1719 B.n750 B.n749 10.6151
R1720 B.n749 B.n746 10.6151
R1721 B.n746 B.n745 10.6151
R1722 B.n745 B.n742 10.6151
R1723 B.n742 B.n741 10.6151
R1724 B.n741 B.n738 10.6151
R1725 B.n738 B.n737 10.6151
R1726 B.n737 B.n734 10.6151
R1727 B.n734 B.n733 10.6151
R1728 B.n733 B.n730 10.6151
R1729 B.n730 B.n729 10.6151
R1730 B.n729 B.n726 10.6151
R1731 B.n726 B.n725 10.6151
R1732 B.n725 B.n722 10.6151
R1733 B.n722 B.n721 10.6151
R1734 B.n721 B.n718 10.6151
R1735 B.n718 B.n717 10.6151
R1736 B.n717 B.n714 10.6151
R1737 B.n714 B.n713 10.6151
R1738 B.n713 B.n710 10.6151
R1739 B.n710 B.n709 10.6151
R1740 B.n709 B.n706 10.6151
R1741 B.n706 B.n705 10.6151
R1742 B.n705 B.n702 10.6151
R1743 B.n702 B.n701 10.6151
R1744 B.n701 B.n698 10.6151
R1745 B.n698 B.n697 10.6151
R1746 B.n694 B.n693 10.6151
R1747 B.n693 B.n690 10.6151
R1748 B.n690 B.n689 10.6151
R1749 B.n689 B.n686 10.6151
R1750 B.n686 B.n685 10.6151
R1751 B.n685 B.n682 10.6151
R1752 B.n682 B.n681 10.6151
R1753 B.n681 B.n678 10.6151
R1754 B.n676 B.n673 10.6151
R1755 B.n673 B.n672 10.6151
R1756 B.n672 B.n669 10.6151
R1757 B.n669 B.n668 10.6151
R1758 B.n668 B.n665 10.6151
R1759 B.n665 B.n664 10.6151
R1760 B.n664 B.n661 10.6151
R1761 B.n661 B.n660 10.6151
R1762 B.n660 B.n657 10.6151
R1763 B.n657 B.n656 10.6151
R1764 B.n656 B.n653 10.6151
R1765 B.n653 B.n652 10.6151
R1766 B.n652 B.n649 10.6151
R1767 B.n649 B.n648 10.6151
R1768 B.n648 B.n645 10.6151
R1769 B.n645 B.n644 10.6151
R1770 B.n644 B.n641 10.6151
R1771 B.n641 B.n640 10.6151
R1772 B.n640 B.n637 10.6151
R1773 B.n637 B.n636 10.6151
R1774 B.n636 B.n633 10.6151
R1775 B.n633 B.n632 10.6151
R1776 B.n632 B.n629 10.6151
R1777 B.n629 B.n628 10.6151
R1778 B.n628 B.n625 10.6151
R1779 B.n625 B.n624 10.6151
R1780 B.n624 B.n621 10.6151
R1781 B.n621 B.n620 10.6151
R1782 B.n620 B.n617 10.6151
R1783 B.n617 B.n616 10.6151
R1784 B.n616 B.n613 10.6151
R1785 B.n613 B.n612 10.6151
R1786 B.n612 B.n609 10.6151
R1787 B.n609 B.n608 10.6151
R1788 B.n608 B.n605 10.6151
R1789 B.n605 B.n604 10.6151
R1790 B.n604 B.n601 10.6151
R1791 B.n601 B.n600 10.6151
R1792 B.n600 B.n597 10.6151
R1793 B.n597 B.n596 10.6151
R1794 B.n596 B.n593 10.6151
R1795 B.n593 B.n592 10.6151
R1796 B.n592 B.n589 10.6151
R1797 B.n589 B.n588 10.6151
R1798 B.n588 B.n585 10.6151
R1799 B.n585 B.n584 10.6151
R1800 B.n584 B.n581 10.6151
R1801 B.n581 B.n580 10.6151
R1802 B.n580 B.n577 10.6151
R1803 B.n577 B.n576 10.6151
R1804 B.n576 B.n573 10.6151
R1805 B.n573 B.n572 10.6151
R1806 B.n572 B.n569 10.6151
R1807 B.n569 B.n568 10.6151
R1808 B.n568 B.n565 10.6151
R1809 B.n565 B.n564 10.6151
R1810 B.n564 B.n561 10.6151
R1811 B.n561 B.n560 10.6151
R1812 B.n560 B.n487 10.6151
R1813 B.n820 B.n487 10.6151
R1814 B.n826 B.n483 10.6151
R1815 B.n827 B.n826 10.6151
R1816 B.n828 B.n827 10.6151
R1817 B.n828 B.n475 10.6151
R1818 B.n838 B.n475 10.6151
R1819 B.n839 B.n838 10.6151
R1820 B.n840 B.n839 10.6151
R1821 B.n840 B.n467 10.6151
R1822 B.n850 B.n467 10.6151
R1823 B.n851 B.n850 10.6151
R1824 B.n852 B.n851 10.6151
R1825 B.n852 B.n459 10.6151
R1826 B.n862 B.n459 10.6151
R1827 B.n863 B.n862 10.6151
R1828 B.n864 B.n863 10.6151
R1829 B.n864 B.n451 10.6151
R1830 B.n875 B.n451 10.6151
R1831 B.n876 B.n875 10.6151
R1832 B.n877 B.n876 10.6151
R1833 B.n877 B.n444 10.6151
R1834 B.n887 B.n444 10.6151
R1835 B.n888 B.n887 10.6151
R1836 B.n889 B.n888 10.6151
R1837 B.n889 B.n436 10.6151
R1838 B.n899 B.n436 10.6151
R1839 B.n900 B.n899 10.6151
R1840 B.n901 B.n900 10.6151
R1841 B.n901 B.n428 10.6151
R1842 B.n911 B.n428 10.6151
R1843 B.n912 B.n911 10.6151
R1844 B.n913 B.n912 10.6151
R1845 B.n913 B.n420 10.6151
R1846 B.n923 B.n420 10.6151
R1847 B.n924 B.n923 10.6151
R1848 B.n925 B.n924 10.6151
R1849 B.n925 B.n412 10.6151
R1850 B.n936 B.n412 10.6151
R1851 B.n937 B.n936 10.6151
R1852 B.n938 B.n937 10.6151
R1853 B.n938 B.n0 10.6151
R1854 B.n1076 B.n1 10.6151
R1855 B.n1076 B.n1075 10.6151
R1856 B.n1075 B.n1074 10.6151
R1857 B.n1074 B.n10 10.6151
R1858 B.n1068 B.n10 10.6151
R1859 B.n1068 B.n1067 10.6151
R1860 B.n1067 B.n1066 10.6151
R1861 B.n1066 B.n17 10.6151
R1862 B.n1060 B.n17 10.6151
R1863 B.n1060 B.n1059 10.6151
R1864 B.n1059 B.n1058 10.6151
R1865 B.n1058 B.n24 10.6151
R1866 B.n1052 B.n24 10.6151
R1867 B.n1052 B.n1051 10.6151
R1868 B.n1051 B.n1050 10.6151
R1869 B.n1050 B.n31 10.6151
R1870 B.n1044 B.n31 10.6151
R1871 B.n1044 B.n1043 10.6151
R1872 B.n1043 B.n1042 10.6151
R1873 B.n1042 B.n38 10.6151
R1874 B.n1036 B.n38 10.6151
R1875 B.n1036 B.n1035 10.6151
R1876 B.n1035 B.n1034 10.6151
R1877 B.n1034 B.n44 10.6151
R1878 B.n1028 B.n44 10.6151
R1879 B.n1028 B.n1027 10.6151
R1880 B.n1027 B.n1026 10.6151
R1881 B.n1026 B.n52 10.6151
R1882 B.n1020 B.n52 10.6151
R1883 B.n1020 B.n1019 10.6151
R1884 B.n1019 B.n1018 10.6151
R1885 B.n1018 B.n59 10.6151
R1886 B.n1012 B.n59 10.6151
R1887 B.n1012 B.n1011 10.6151
R1888 B.n1011 B.n1010 10.6151
R1889 B.n1010 B.n66 10.6151
R1890 B.n1004 B.n66 10.6151
R1891 B.n1004 B.n1003 10.6151
R1892 B.n1003 B.n1002 10.6151
R1893 B.n1002 B.n73 10.6151
R1894 B.n927 B.t2 8.76912
R1895 B.t3 B.n1070 8.76912
R1896 B.n271 B.n270 6.5566
R1897 B.n287 B.n145 6.5566
R1898 B.n694 B.n556 6.5566
R1899 B.n678 B.n677 6.5566
R1900 B.n879 B.t5 6.00008
R1901 B.n1038 B.t4 6.00008
R1902 B.n270 B.n269 4.05904
R1903 B.n290 B.n145 4.05904
R1904 B.n697 B.n556 4.05904
R1905 B.n677 B.n676 4.05904
R1906 B.n1082 B.n0 2.81026
R1907 B.n1082 B.n1 2.81026
R1908 B.n903 B.t1 1.38502
R1909 B.t0 B.n1054 1.38502
R1910 VP.n9 VP.t5 216.238
R1911 VP.n30 VP.t3 181.093
R1912 VP.n20 VP.t2 181.093
R1913 VP.n38 VP.t0 181.093
R1914 VP.n10 VP.t4 181.093
R1915 VP.n18 VP.t1 181.093
R1916 VP.n11 VP.n8 161.3
R1917 VP.n13 VP.n12 161.3
R1918 VP.n14 VP.n7 161.3
R1919 VP.n16 VP.n15 161.3
R1920 VP.n17 VP.n6 161.3
R1921 VP.n37 VP.n0 161.3
R1922 VP.n36 VP.n35 161.3
R1923 VP.n34 VP.n1 161.3
R1924 VP.n33 VP.n32 161.3
R1925 VP.n31 VP.n2 161.3
R1926 VP.n30 VP.n29 161.3
R1927 VP.n28 VP.n3 161.3
R1928 VP.n27 VP.n26 161.3
R1929 VP.n25 VP.n4 161.3
R1930 VP.n24 VP.n23 161.3
R1931 VP.n22 VP.n5 161.3
R1932 VP.n21 VP.n20 96.1531
R1933 VP.n39 VP.n38 96.1531
R1934 VP.n19 VP.n18 96.1531
R1935 VP.n21 VP.n19 53.1966
R1936 VP.n26 VP.n25 50.2647
R1937 VP.n32 VP.n1 50.2647
R1938 VP.n12 VP.n7 50.2647
R1939 VP.n10 VP.n9 48.1821
R1940 VP.n25 VP.n24 30.8893
R1941 VP.n36 VP.n1 30.8893
R1942 VP.n16 VP.n7 30.8893
R1943 VP.n24 VP.n5 24.5923
R1944 VP.n26 VP.n3 24.5923
R1945 VP.n30 VP.n3 24.5923
R1946 VP.n31 VP.n30 24.5923
R1947 VP.n32 VP.n31 24.5923
R1948 VP.n37 VP.n36 24.5923
R1949 VP.n17 VP.n16 24.5923
R1950 VP.n11 VP.n10 24.5923
R1951 VP.n12 VP.n11 24.5923
R1952 VP.n20 VP.n5 14.7556
R1953 VP.n38 VP.n37 14.7556
R1954 VP.n18 VP.n17 14.7556
R1955 VP.n9 VP.n8 6.50797
R1956 VP.n19 VP.n6 0.278335
R1957 VP.n22 VP.n21 0.278335
R1958 VP.n39 VP.n0 0.278335
R1959 VP.n13 VP.n8 0.189894
R1960 VP.n14 VP.n13 0.189894
R1961 VP.n15 VP.n14 0.189894
R1962 VP.n15 VP.n6 0.189894
R1963 VP.n23 VP.n22 0.189894
R1964 VP.n23 VP.n4 0.189894
R1965 VP.n27 VP.n4 0.189894
R1966 VP.n28 VP.n27 0.189894
R1967 VP.n29 VP.n28 0.189894
R1968 VP.n29 VP.n2 0.189894
R1969 VP.n33 VP.n2 0.189894
R1970 VP.n34 VP.n33 0.189894
R1971 VP.n35 VP.n34 0.189894
R1972 VP.n35 VP.n0 0.189894
R1973 VP VP.n39 0.153485
R1974 VDD1 VDD1.t0 62.7936
R1975 VDD1.n1 VDD1.t3 62.6799
R1976 VDD1.n1 VDD1.n0 60.4062
R1977 VDD1.n3 VDD1.n2 59.8581
R1978 VDD1.n3 VDD1.n1 49.35
R1979 VDD1.n2 VDD1.t1 1.06731
R1980 VDD1.n2 VDD1.t4 1.06731
R1981 VDD1.n0 VDD1.t2 1.06731
R1982 VDD1.n0 VDD1.t5 1.06731
R1983 VDD1 VDD1.n3 0.545759
C0 VN VP 8.00807f
C1 VDD2 VDD1 1.35685f
C2 VDD2 VTAIL 10.1858f
C3 VDD1 VP 10.3833f
C4 VTAIL VP 9.94159f
C5 VDD1 VN 0.150851f
C6 VN VTAIL 9.927191f
C7 VDD1 VTAIL 10.1376f
C8 VDD2 VP 0.448137f
C9 VDD2 VN 10.090401f
C10 VDD2 B 7.05935f
C11 VDD1 B 7.377079f
C12 VTAIL B 10.34212f
C13 VN B 13.073319f
C14 VP B 11.554001f
C15 VDD1.t0 B 3.66138f
C16 VDD1.t3 B 3.6605f
C17 VDD1.t2 B 0.313203f
C18 VDD1.t5 B 0.313203f
C19 VDD1.n0 B 2.85904f
C20 VDD1.n1 B 2.90094f
C21 VDD1.t1 B 0.313203f
C22 VDD1.t4 B 0.313203f
C23 VDD1.n2 B 2.85547f
C24 VDD1.n3 B 2.77926f
C25 VP.n0 B 0.03062f
C26 VP.t0 B 2.93038f
C27 VP.n1 B 0.021899f
C28 VP.n2 B 0.023226f
C29 VP.t3 B 2.93038f
C30 VP.n3 B 0.043071f
C31 VP.n4 B 0.023226f
C32 VP.n5 B 0.034566f
C33 VP.n6 B 0.03062f
C34 VP.t1 B 2.93038f
C35 VP.n7 B 0.021899f
C36 VP.n8 B 0.221227f
C37 VP.t4 B 2.93038f
C38 VP.t5 B 3.11853f
C39 VP.n9 B 1.05429f
C40 VP.n10 B 1.09304f
C41 VP.n11 B 0.043071f
C42 VP.n12 B 0.042419f
C43 VP.n13 B 0.023226f
C44 VP.n14 B 0.023226f
C45 VP.n15 B 0.023226f
C46 VP.n16 B 0.046279f
C47 VP.n17 B 0.034566f
C48 VP.n18 B 1.09556f
C49 VP.n19 B 1.41018f
C50 VP.t2 B 2.93038f
C51 VP.n20 B 1.09556f
C52 VP.n21 B 1.42592f
C53 VP.n22 B 0.03062f
C54 VP.n23 B 0.023226f
C55 VP.n24 B 0.046279f
C56 VP.n25 B 0.021899f
C57 VP.n26 B 0.042419f
C58 VP.n27 B 0.023226f
C59 VP.n28 B 0.023226f
C60 VP.n29 B 0.023226f
C61 VP.n30 B 1.03773f
C62 VP.n31 B 0.043071f
C63 VP.n32 B 0.042419f
C64 VP.n33 B 0.023226f
C65 VP.n34 B 0.023226f
C66 VP.n35 B 0.023226f
C67 VP.n36 B 0.046279f
C68 VP.n37 B 0.034566f
C69 VP.n38 B 1.09556f
C70 VP.n39 B 0.033902f
C71 VTAIL.t6 B 0.327775f
C72 VTAIL.t11 B 0.327775f
C73 VTAIL.n0 B 2.9176f
C74 VTAIL.n1 B 0.396109f
C75 VTAIL.t2 B 3.72753f
C76 VTAIL.n2 B 0.60629f
C77 VTAIL.t5 B 0.327775f
C78 VTAIL.t1 B 0.327775f
C79 VTAIL.n3 B 2.9176f
C80 VTAIL.n4 B 2.20494f
C81 VTAIL.t7 B 0.327775f
C82 VTAIL.t8 B 0.327775f
C83 VTAIL.n5 B 2.91761f
C84 VTAIL.n6 B 2.20493f
C85 VTAIL.t9 B 3.72755f
C86 VTAIL.n7 B 0.606268f
C87 VTAIL.t3 B 0.327775f
C88 VTAIL.t0 B 0.327775f
C89 VTAIL.n8 B 2.91761f
C90 VTAIL.n9 B 0.52228f
C91 VTAIL.t4 B 3.72753f
C92 VTAIL.n10 B 2.11512f
C93 VTAIL.t10 B 3.72753f
C94 VTAIL.n11 B 2.06748f
C95 VDD2.t4 B 3.63879f
C96 VDD2.t2 B 0.311345f
C97 VDD2.t0 B 0.311345f
C98 VDD2.n0 B 2.84208f
C99 VDD2.n1 B 2.77769f
C100 VDD2.t5 B 3.62855f
C101 VDD2.n2 B 2.77494f
C102 VDD2.t3 B 0.311345f
C103 VDD2.t1 B 0.311345f
C104 VDD2.n3 B 2.84205f
C105 VN.n0 B 0.03026f
C106 VN.t1 B 2.89598f
C107 VN.n1 B 0.021642f
C108 VN.n2 B 0.21863f
C109 VN.t0 B 2.89598f
C110 VN.t5 B 3.08191f
C111 VN.n3 B 1.04192f
C112 VN.n4 B 1.08021f
C113 VN.n5 B 0.042565f
C114 VN.n6 B 0.041921f
C115 VN.n7 B 0.022954f
C116 VN.n8 B 0.022954f
C117 VN.n9 B 0.022954f
C118 VN.n10 B 0.045735f
C119 VN.n11 B 0.03416f
C120 VN.n12 B 1.0827f
C121 VN.n13 B 0.033504f
C122 VN.n14 B 0.03026f
C123 VN.t4 B 2.89598f
C124 VN.n15 B 0.021642f
C125 VN.n16 B 0.21863f
C126 VN.t3 B 2.89598f
C127 VN.t2 B 3.08191f
C128 VN.n17 B 1.04192f
C129 VN.n18 B 1.08021f
C130 VN.n19 B 0.042565f
C131 VN.n20 B 0.041921f
C132 VN.n21 B 0.022954f
C133 VN.n22 B 0.022954f
C134 VN.n23 B 0.022954f
C135 VN.n24 B 0.045735f
C136 VN.n25 B 0.03416f
C137 VN.n26 B 1.0827f
C138 VN.n27 B 1.40583f
.ends

