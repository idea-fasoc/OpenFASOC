* NGSPICE file created from diff_pair_sample_0573.ext - technology: sky130A

.subckt diff_pair_sample_0573 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2212_n1208# sky130_fd_pr__pfet_01v8 ad=0.468 pd=3.18 as=0 ps=0 w=1.2 l=1.74
X1 VTAIL.t7 VN.t0 VDD2.t2 w_n2212_n1208# sky130_fd_pr__pfet_01v8 ad=0.468 pd=3.18 as=0.198 ps=1.53 w=1.2 l=1.74
X2 VDD1.t3 VP.t0 VTAIL.t1 w_n2212_n1208# sky130_fd_pr__pfet_01v8 ad=0.198 pd=1.53 as=0.468 ps=3.18 w=1.2 l=1.74
X3 VDD2.t1 VN.t1 VTAIL.t6 w_n2212_n1208# sky130_fd_pr__pfet_01v8 ad=0.198 pd=1.53 as=0.468 ps=3.18 w=1.2 l=1.74
X4 B.t8 B.t6 B.t7 w_n2212_n1208# sky130_fd_pr__pfet_01v8 ad=0.468 pd=3.18 as=0 ps=0 w=1.2 l=1.74
X5 VTAIL.t2 VP.t1 VDD1.t2 w_n2212_n1208# sky130_fd_pr__pfet_01v8 ad=0.468 pd=3.18 as=0.198 ps=1.53 w=1.2 l=1.74
X6 B.t5 B.t3 B.t4 w_n2212_n1208# sky130_fd_pr__pfet_01v8 ad=0.468 pd=3.18 as=0 ps=0 w=1.2 l=1.74
X7 VTAIL.t5 VN.t2 VDD2.t3 w_n2212_n1208# sky130_fd_pr__pfet_01v8 ad=0.468 pd=3.18 as=0.198 ps=1.53 w=1.2 l=1.74
X8 VDD2.t0 VN.t3 VTAIL.t4 w_n2212_n1208# sky130_fd_pr__pfet_01v8 ad=0.198 pd=1.53 as=0.468 ps=3.18 w=1.2 l=1.74
X9 VTAIL.t3 VP.t2 VDD1.t1 w_n2212_n1208# sky130_fd_pr__pfet_01v8 ad=0.468 pd=3.18 as=0.198 ps=1.53 w=1.2 l=1.74
X10 VDD1.t0 VP.t3 VTAIL.t0 w_n2212_n1208# sky130_fd_pr__pfet_01v8 ad=0.198 pd=1.53 as=0.468 ps=3.18 w=1.2 l=1.74
X11 B.t2 B.t0 B.t1 w_n2212_n1208# sky130_fd_pr__pfet_01v8 ad=0.468 pd=3.18 as=0 ps=0 w=1.2 l=1.74
R0 B.n174 B.n61 585
R1 B.n173 B.n172 585
R2 B.n171 B.n62 585
R3 B.n170 B.n169 585
R4 B.n168 B.n63 585
R5 B.n167 B.n166 585
R6 B.n165 B.n64 585
R7 B.n164 B.n163 585
R8 B.n162 B.n65 585
R9 B.n161 B.n160 585
R10 B.n159 B.n158 585
R11 B.n157 B.n69 585
R12 B.n156 B.n155 585
R13 B.n154 B.n70 585
R14 B.n153 B.n152 585
R15 B.n151 B.n71 585
R16 B.n150 B.n149 585
R17 B.n148 B.n72 585
R18 B.n147 B.n146 585
R19 B.n144 B.n73 585
R20 B.n143 B.n142 585
R21 B.n141 B.n76 585
R22 B.n140 B.n139 585
R23 B.n138 B.n77 585
R24 B.n137 B.n136 585
R25 B.n135 B.n78 585
R26 B.n134 B.n133 585
R27 B.n132 B.n79 585
R28 B.n131 B.n130 585
R29 B.n176 B.n175 585
R30 B.n177 B.n60 585
R31 B.n179 B.n178 585
R32 B.n180 B.n59 585
R33 B.n182 B.n181 585
R34 B.n183 B.n58 585
R35 B.n185 B.n184 585
R36 B.n186 B.n57 585
R37 B.n188 B.n187 585
R38 B.n189 B.n56 585
R39 B.n191 B.n190 585
R40 B.n192 B.n55 585
R41 B.n194 B.n193 585
R42 B.n195 B.n54 585
R43 B.n197 B.n196 585
R44 B.n198 B.n53 585
R45 B.n200 B.n199 585
R46 B.n201 B.n52 585
R47 B.n203 B.n202 585
R48 B.n204 B.n51 585
R49 B.n206 B.n205 585
R50 B.n207 B.n50 585
R51 B.n209 B.n208 585
R52 B.n210 B.n49 585
R53 B.n212 B.n211 585
R54 B.n213 B.n48 585
R55 B.n215 B.n214 585
R56 B.n216 B.n47 585
R57 B.n218 B.n217 585
R58 B.n219 B.n46 585
R59 B.n221 B.n220 585
R60 B.n222 B.n45 585
R61 B.n224 B.n223 585
R62 B.n225 B.n44 585
R63 B.n227 B.n226 585
R64 B.n228 B.n43 585
R65 B.n230 B.n229 585
R66 B.n231 B.n42 585
R67 B.n233 B.n232 585
R68 B.n234 B.n41 585
R69 B.n236 B.n235 585
R70 B.n237 B.n40 585
R71 B.n239 B.n238 585
R72 B.n240 B.n39 585
R73 B.n242 B.n241 585
R74 B.n243 B.n38 585
R75 B.n245 B.n244 585
R76 B.n246 B.n37 585
R77 B.n248 B.n247 585
R78 B.n249 B.n36 585
R79 B.n251 B.n250 585
R80 B.n252 B.n35 585
R81 B.n254 B.n253 585
R82 B.n255 B.n34 585
R83 B.n300 B.n15 585
R84 B.n299 B.n298 585
R85 B.n297 B.n16 585
R86 B.n296 B.n295 585
R87 B.n294 B.n17 585
R88 B.n293 B.n292 585
R89 B.n291 B.n18 585
R90 B.n290 B.n289 585
R91 B.n288 B.n19 585
R92 B.n287 B.n286 585
R93 B.n285 B.n284 585
R94 B.n283 B.n23 585
R95 B.n282 B.n281 585
R96 B.n280 B.n24 585
R97 B.n279 B.n278 585
R98 B.n277 B.n25 585
R99 B.n276 B.n275 585
R100 B.n274 B.n26 585
R101 B.n273 B.n272 585
R102 B.n270 B.n27 585
R103 B.n269 B.n268 585
R104 B.n267 B.n30 585
R105 B.n266 B.n265 585
R106 B.n264 B.n31 585
R107 B.n263 B.n262 585
R108 B.n261 B.n32 585
R109 B.n260 B.n259 585
R110 B.n258 B.n33 585
R111 B.n257 B.n256 585
R112 B.n302 B.n301 585
R113 B.n303 B.n14 585
R114 B.n305 B.n304 585
R115 B.n306 B.n13 585
R116 B.n308 B.n307 585
R117 B.n309 B.n12 585
R118 B.n311 B.n310 585
R119 B.n312 B.n11 585
R120 B.n314 B.n313 585
R121 B.n315 B.n10 585
R122 B.n317 B.n316 585
R123 B.n318 B.n9 585
R124 B.n320 B.n319 585
R125 B.n321 B.n8 585
R126 B.n323 B.n322 585
R127 B.n324 B.n7 585
R128 B.n326 B.n325 585
R129 B.n327 B.n6 585
R130 B.n329 B.n328 585
R131 B.n330 B.n5 585
R132 B.n332 B.n331 585
R133 B.n333 B.n4 585
R134 B.n335 B.n334 585
R135 B.n336 B.n3 585
R136 B.n338 B.n337 585
R137 B.n339 B.n0 585
R138 B.n2 B.n1 585
R139 B.n93 B.n92 585
R140 B.n95 B.n94 585
R141 B.n96 B.n91 585
R142 B.n98 B.n97 585
R143 B.n99 B.n90 585
R144 B.n101 B.n100 585
R145 B.n102 B.n89 585
R146 B.n104 B.n103 585
R147 B.n105 B.n88 585
R148 B.n107 B.n106 585
R149 B.n108 B.n87 585
R150 B.n110 B.n109 585
R151 B.n111 B.n86 585
R152 B.n113 B.n112 585
R153 B.n114 B.n85 585
R154 B.n116 B.n115 585
R155 B.n117 B.n84 585
R156 B.n119 B.n118 585
R157 B.n120 B.n83 585
R158 B.n122 B.n121 585
R159 B.n123 B.n82 585
R160 B.n125 B.n124 585
R161 B.n126 B.n81 585
R162 B.n128 B.n127 585
R163 B.n129 B.n80 585
R164 B.n130 B.n129 502.111
R165 B.n176 B.n61 502.111
R166 B.n256 B.n255 502.111
R167 B.n302 B.n15 502.111
R168 B.n74 B.t10 405.224
R169 B.n66 B.t1 405.224
R170 B.n28 B.t5 405.224
R171 B.n20 B.t8 405.224
R172 B.n75 B.t11 365.079
R173 B.n67 B.t2 365.079
R174 B.n29 B.t4 365.079
R175 B.n21 B.t7 365.079
R176 B.n341 B.n340 256.663
R177 B.n340 B.n339 235.042
R178 B.n340 B.n2 235.042
R179 B.n74 B.t9 222.856
R180 B.n66 B.t0 222.856
R181 B.n28 B.t3 222.856
R182 B.n20 B.t6 222.856
R183 B.n130 B.n79 163.367
R184 B.n134 B.n79 163.367
R185 B.n135 B.n134 163.367
R186 B.n136 B.n135 163.367
R187 B.n136 B.n77 163.367
R188 B.n140 B.n77 163.367
R189 B.n141 B.n140 163.367
R190 B.n142 B.n141 163.367
R191 B.n142 B.n73 163.367
R192 B.n147 B.n73 163.367
R193 B.n148 B.n147 163.367
R194 B.n149 B.n148 163.367
R195 B.n149 B.n71 163.367
R196 B.n153 B.n71 163.367
R197 B.n154 B.n153 163.367
R198 B.n155 B.n154 163.367
R199 B.n155 B.n69 163.367
R200 B.n159 B.n69 163.367
R201 B.n160 B.n159 163.367
R202 B.n160 B.n65 163.367
R203 B.n164 B.n65 163.367
R204 B.n165 B.n164 163.367
R205 B.n166 B.n165 163.367
R206 B.n166 B.n63 163.367
R207 B.n170 B.n63 163.367
R208 B.n171 B.n170 163.367
R209 B.n172 B.n171 163.367
R210 B.n172 B.n61 163.367
R211 B.n255 B.n254 163.367
R212 B.n254 B.n35 163.367
R213 B.n250 B.n35 163.367
R214 B.n250 B.n249 163.367
R215 B.n249 B.n248 163.367
R216 B.n248 B.n37 163.367
R217 B.n244 B.n37 163.367
R218 B.n244 B.n243 163.367
R219 B.n243 B.n242 163.367
R220 B.n242 B.n39 163.367
R221 B.n238 B.n39 163.367
R222 B.n238 B.n237 163.367
R223 B.n237 B.n236 163.367
R224 B.n236 B.n41 163.367
R225 B.n232 B.n41 163.367
R226 B.n232 B.n231 163.367
R227 B.n231 B.n230 163.367
R228 B.n230 B.n43 163.367
R229 B.n226 B.n43 163.367
R230 B.n226 B.n225 163.367
R231 B.n225 B.n224 163.367
R232 B.n224 B.n45 163.367
R233 B.n220 B.n45 163.367
R234 B.n220 B.n219 163.367
R235 B.n219 B.n218 163.367
R236 B.n218 B.n47 163.367
R237 B.n214 B.n47 163.367
R238 B.n214 B.n213 163.367
R239 B.n213 B.n212 163.367
R240 B.n212 B.n49 163.367
R241 B.n208 B.n49 163.367
R242 B.n208 B.n207 163.367
R243 B.n207 B.n206 163.367
R244 B.n206 B.n51 163.367
R245 B.n202 B.n51 163.367
R246 B.n202 B.n201 163.367
R247 B.n201 B.n200 163.367
R248 B.n200 B.n53 163.367
R249 B.n196 B.n53 163.367
R250 B.n196 B.n195 163.367
R251 B.n195 B.n194 163.367
R252 B.n194 B.n55 163.367
R253 B.n190 B.n55 163.367
R254 B.n190 B.n189 163.367
R255 B.n189 B.n188 163.367
R256 B.n188 B.n57 163.367
R257 B.n184 B.n57 163.367
R258 B.n184 B.n183 163.367
R259 B.n183 B.n182 163.367
R260 B.n182 B.n59 163.367
R261 B.n178 B.n59 163.367
R262 B.n178 B.n177 163.367
R263 B.n177 B.n176 163.367
R264 B.n298 B.n15 163.367
R265 B.n298 B.n297 163.367
R266 B.n297 B.n296 163.367
R267 B.n296 B.n17 163.367
R268 B.n292 B.n17 163.367
R269 B.n292 B.n291 163.367
R270 B.n291 B.n290 163.367
R271 B.n290 B.n19 163.367
R272 B.n286 B.n19 163.367
R273 B.n286 B.n285 163.367
R274 B.n285 B.n23 163.367
R275 B.n281 B.n23 163.367
R276 B.n281 B.n280 163.367
R277 B.n280 B.n279 163.367
R278 B.n279 B.n25 163.367
R279 B.n275 B.n25 163.367
R280 B.n275 B.n274 163.367
R281 B.n274 B.n273 163.367
R282 B.n273 B.n27 163.367
R283 B.n268 B.n27 163.367
R284 B.n268 B.n267 163.367
R285 B.n267 B.n266 163.367
R286 B.n266 B.n31 163.367
R287 B.n262 B.n31 163.367
R288 B.n262 B.n261 163.367
R289 B.n261 B.n260 163.367
R290 B.n260 B.n33 163.367
R291 B.n256 B.n33 163.367
R292 B.n303 B.n302 163.367
R293 B.n304 B.n303 163.367
R294 B.n304 B.n13 163.367
R295 B.n308 B.n13 163.367
R296 B.n309 B.n308 163.367
R297 B.n310 B.n309 163.367
R298 B.n310 B.n11 163.367
R299 B.n314 B.n11 163.367
R300 B.n315 B.n314 163.367
R301 B.n316 B.n315 163.367
R302 B.n316 B.n9 163.367
R303 B.n320 B.n9 163.367
R304 B.n321 B.n320 163.367
R305 B.n322 B.n321 163.367
R306 B.n322 B.n7 163.367
R307 B.n326 B.n7 163.367
R308 B.n327 B.n326 163.367
R309 B.n328 B.n327 163.367
R310 B.n328 B.n5 163.367
R311 B.n332 B.n5 163.367
R312 B.n333 B.n332 163.367
R313 B.n334 B.n333 163.367
R314 B.n334 B.n3 163.367
R315 B.n338 B.n3 163.367
R316 B.n339 B.n338 163.367
R317 B.n93 B.n2 163.367
R318 B.n94 B.n93 163.367
R319 B.n94 B.n91 163.367
R320 B.n98 B.n91 163.367
R321 B.n99 B.n98 163.367
R322 B.n100 B.n99 163.367
R323 B.n100 B.n89 163.367
R324 B.n104 B.n89 163.367
R325 B.n105 B.n104 163.367
R326 B.n106 B.n105 163.367
R327 B.n106 B.n87 163.367
R328 B.n110 B.n87 163.367
R329 B.n111 B.n110 163.367
R330 B.n112 B.n111 163.367
R331 B.n112 B.n85 163.367
R332 B.n116 B.n85 163.367
R333 B.n117 B.n116 163.367
R334 B.n118 B.n117 163.367
R335 B.n118 B.n83 163.367
R336 B.n122 B.n83 163.367
R337 B.n123 B.n122 163.367
R338 B.n124 B.n123 163.367
R339 B.n124 B.n81 163.367
R340 B.n128 B.n81 163.367
R341 B.n129 B.n128 163.367
R342 B.n145 B.n75 59.5399
R343 B.n68 B.n67 59.5399
R344 B.n271 B.n29 59.5399
R345 B.n22 B.n21 59.5399
R346 B.n75 B.n74 40.146
R347 B.n67 B.n66 40.146
R348 B.n29 B.n28 40.146
R349 B.n21 B.n20 40.146
R350 B.n301 B.n300 32.6249
R351 B.n257 B.n34 32.6249
R352 B.n175 B.n174 32.6249
R353 B.n131 B.n80 32.6249
R354 B B.n341 18.0485
R355 B.n301 B.n14 10.6151
R356 B.n305 B.n14 10.6151
R357 B.n306 B.n305 10.6151
R358 B.n307 B.n306 10.6151
R359 B.n307 B.n12 10.6151
R360 B.n311 B.n12 10.6151
R361 B.n312 B.n311 10.6151
R362 B.n313 B.n312 10.6151
R363 B.n313 B.n10 10.6151
R364 B.n317 B.n10 10.6151
R365 B.n318 B.n317 10.6151
R366 B.n319 B.n318 10.6151
R367 B.n319 B.n8 10.6151
R368 B.n323 B.n8 10.6151
R369 B.n324 B.n323 10.6151
R370 B.n325 B.n324 10.6151
R371 B.n325 B.n6 10.6151
R372 B.n329 B.n6 10.6151
R373 B.n330 B.n329 10.6151
R374 B.n331 B.n330 10.6151
R375 B.n331 B.n4 10.6151
R376 B.n335 B.n4 10.6151
R377 B.n336 B.n335 10.6151
R378 B.n337 B.n336 10.6151
R379 B.n337 B.n0 10.6151
R380 B.n300 B.n299 10.6151
R381 B.n299 B.n16 10.6151
R382 B.n295 B.n16 10.6151
R383 B.n295 B.n294 10.6151
R384 B.n294 B.n293 10.6151
R385 B.n293 B.n18 10.6151
R386 B.n289 B.n18 10.6151
R387 B.n289 B.n288 10.6151
R388 B.n288 B.n287 10.6151
R389 B.n284 B.n283 10.6151
R390 B.n283 B.n282 10.6151
R391 B.n282 B.n24 10.6151
R392 B.n278 B.n24 10.6151
R393 B.n278 B.n277 10.6151
R394 B.n277 B.n276 10.6151
R395 B.n276 B.n26 10.6151
R396 B.n272 B.n26 10.6151
R397 B.n270 B.n269 10.6151
R398 B.n269 B.n30 10.6151
R399 B.n265 B.n30 10.6151
R400 B.n265 B.n264 10.6151
R401 B.n264 B.n263 10.6151
R402 B.n263 B.n32 10.6151
R403 B.n259 B.n32 10.6151
R404 B.n259 B.n258 10.6151
R405 B.n258 B.n257 10.6151
R406 B.n253 B.n34 10.6151
R407 B.n253 B.n252 10.6151
R408 B.n252 B.n251 10.6151
R409 B.n251 B.n36 10.6151
R410 B.n247 B.n36 10.6151
R411 B.n247 B.n246 10.6151
R412 B.n246 B.n245 10.6151
R413 B.n245 B.n38 10.6151
R414 B.n241 B.n38 10.6151
R415 B.n241 B.n240 10.6151
R416 B.n240 B.n239 10.6151
R417 B.n239 B.n40 10.6151
R418 B.n235 B.n40 10.6151
R419 B.n235 B.n234 10.6151
R420 B.n234 B.n233 10.6151
R421 B.n233 B.n42 10.6151
R422 B.n229 B.n42 10.6151
R423 B.n229 B.n228 10.6151
R424 B.n228 B.n227 10.6151
R425 B.n227 B.n44 10.6151
R426 B.n223 B.n44 10.6151
R427 B.n223 B.n222 10.6151
R428 B.n222 B.n221 10.6151
R429 B.n221 B.n46 10.6151
R430 B.n217 B.n46 10.6151
R431 B.n217 B.n216 10.6151
R432 B.n216 B.n215 10.6151
R433 B.n215 B.n48 10.6151
R434 B.n211 B.n48 10.6151
R435 B.n211 B.n210 10.6151
R436 B.n210 B.n209 10.6151
R437 B.n209 B.n50 10.6151
R438 B.n205 B.n50 10.6151
R439 B.n205 B.n204 10.6151
R440 B.n204 B.n203 10.6151
R441 B.n203 B.n52 10.6151
R442 B.n199 B.n52 10.6151
R443 B.n199 B.n198 10.6151
R444 B.n198 B.n197 10.6151
R445 B.n197 B.n54 10.6151
R446 B.n193 B.n54 10.6151
R447 B.n193 B.n192 10.6151
R448 B.n192 B.n191 10.6151
R449 B.n191 B.n56 10.6151
R450 B.n187 B.n56 10.6151
R451 B.n187 B.n186 10.6151
R452 B.n186 B.n185 10.6151
R453 B.n185 B.n58 10.6151
R454 B.n181 B.n58 10.6151
R455 B.n181 B.n180 10.6151
R456 B.n180 B.n179 10.6151
R457 B.n179 B.n60 10.6151
R458 B.n175 B.n60 10.6151
R459 B.n92 B.n1 10.6151
R460 B.n95 B.n92 10.6151
R461 B.n96 B.n95 10.6151
R462 B.n97 B.n96 10.6151
R463 B.n97 B.n90 10.6151
R464 B.n101 B.n90 10.6151
R465 B.n102 B.n101 10.6151
R466 B.n103 B.n102 10.6151
R467 B.n103 B.n88 10.6151
R468 B.n107 B.n88 10.6151
R469 B.n108 B.n107 10.6151
R470 B.n109 B.n108 10.6151
R471 B.n109 B.n86 10.6151
R472 B.n113 B.n86 10.6151
R473 B.n114 B.n113 10.6151
R474 B.n115 B.n114 10.6151
R475 B.n115 B.n84 10.6151
R476 B.n119 B.n84 10.6151
R477 B.n120 B.n119 10.6151
R478 B.n121 B.n120 10.6151
R479 B.n121 B.n82 10.6151
R480 B.n125 B.n82 10.6151
R481 B.n126 B.n125 10.6151
R482 B.n127 B.n126 10.6151
R483 B.n127 B.n80 10.6151
R484 B.n132 B.n131 10.6151
R485 B.n133 B.n132 10.6151
R486 B.n133 B.n78 10.6151
R487 B.n137 B.n78 10.6151
R488 B.n138 B.n137 10.6151
R489 B.n139 B.n138 10.6151
R490 B.n139 B.n76 10.6151
R491 B.n143 B.n76 10.6151
R492 B.n144 B.n143 10.6151
R493 B.n146 B.n72 10.6151
R494 B.n150 B.n72 10.6151
R495 B.n151 B.n150 10.6151
R496 B.n152 B.n151 10.6151
R497 B.n152 B.n70 10.6151
R498 B.n156 B.n70 10.6151
R499 B.n157 B.n156 10.6151
R500 B.n158 B.n157 10.6151
R501 B.n162 B.n161 10.6151
R502 B.n163 B.n162 10.6151
R503 B.n163 B.n64 10.6151
R504 B.n167 B.n64 10.6151
R505 B.n168 B.n167 10.6151
R506 B.n169 B.n168 10.6151
R507 B.n169 B.n62 10.6151
R508 B.n173 B.n62 10.6151
R509 B.n174 B.n173 10.6151
R510 B.n341 B.n0 8.11757
R511 B.n341 B.n1 8.11757
R512 B.n284 B.n22 6.5566
R513 B.n272 B.n271 6.5566
R514 B.n146 B.n145 6.5566
R515 B.n158 B.n68 6.5566
R516 B.n287 B.n22 4.05904
R517 B.n271 B.n270 4.05904
R518 B.n145 B.n144 4.05904
R519 B.n161 B.n68 4.05904
R520 VN.n0 VN.t0 52.34
R521 VN.n1 VN.t1 52.34
R522 VN.n0 VN.t3 51.9142
R523 VN.n1 VN.t2 51.9142
R524 VN VN.n1 45.183
R525 VN VN.n0 9.44437
R526 VDD2.n2 VDD2.n0 374.993
R527 VDD2.n2 VDD2.n1 344.89
R528 VDD2.n1 VDD2.t3 27.088
R529 VDD2.n1 VDD2.t1 27.088
R530 VDD2.n0 VDD2.t2 27.088
R531 VDD2.n0 VDD2.t0 27.088
R532 VDD2 VDD2.n2 0.0586897
R533 VTAIL.n7 VTAIL.t4 371.149
R534 VTAIL.n0 VTAIL.t7 371.149
R535 VTAIL.n1 VTAIL.t0 371.149
R536 VTAIL.n2 VTAIL.t2 371.149
R537 VTAIL.n6 VTAIL.t1 371.149
R538 VTAIL.n5 VTAIL.t3 371.149
R539 VTAIL.n4 VTAIL.t6 371.149
R540 VTAIL.n3 VTAIL.t5 371.149
R541 VTAIL.n7 VTAIL.n6 15.1858
R542 VTAIL.n3 VTAIL.n2 15.1858
R543 VTAIL.n4 VTAIL.n3 1.78498
R544 VTAIL.n6 VTAIL.n5 1.78498
R545 VTAIL.n2 VTAIL.n1 1.78498
R546 VTAIL VTAIL.n0 0.950931
R547 VTAIL VTAIL.n7 0.834552
R548 VTAIL.n5 VTAIL.n4 0.470328
R549 VTAIL.n1 VTAIL.n0 0.470328
R550 VP.n5 VP.n4 184.171
R551 VP.n14 VP.n13 184.171
R552 VP.n12 VP.n0 161.3
R553 VP.n11 VP.n10 161.3
R554 VP.n9 VP.n1 161.3
R555 VP.n8 VP.n7 161.3
R556 VP.n6 VP.n2 161.3
R557 VP.n3 VP.t2 52.34
R558 VP.n3 VP.t0 51.9142
R559 VP.n4 VP.n3 44.8023
R560 VP.n7 VP.n1 40.577
R561 VP.n11 VP.n1 40.577
R562 VP.n7 VP.n6 24.5923
R563 VP.n12 VP.n11 24.5923
R564 VP.n5 VP.t1 16.6212
R565 VP.n13 VP.t3 16.6212
R566 VP.n6 VP.n5 1.72193
R567 VP.n13 VP.n12 1.72193
R568 VP.n4 VP.n2 0.189894
R569 VP.n8 VP.n2 0.189894
R570 VP.n9 VP.n8 0.189894
R571 VP.n10 VP.n9 0.189894
R572 VP.n10 VP.n0 0.189894
R573 VP.n14 VP.n0 0.189894
R574 VP VP.n14 0.0516364
R575 VDD1 VDD1.n1 375.517
R576 VDD1 VDD1.n0 344.949
R577 VDD1.n0 VDD1.t1 27.088
R578 VDD1.n0 VDD1.t3 27.088
R579 VDD1.n1 VDD1.t2 27.088
R580 VDD1.n1 VDD1.t0 27.088
C0 VDD2 VN 0.72307f
C1 VDD2 w_n2212_n1208# 1.01969f
C2 B VP 1.24607f
C3 B VDD2 0.85695f
C4 VP VTAIL 1.17413f
C5 VDD1 VN 0.1551f
C6 VDD1 w_n2212_n1208# 0.9838f
C7 VN w_n2212_n1208# 3.35298f
C8 VDD2 VTAIL 2.44132f
C9 B VDD1 0.818441f
C10 B VN 0.782926f
C11 VDD2 VP 0.347595f
C12 B w_n2212_n1208# 5.18073f
C13 VDD1 VTAIL 2.39288f
C14 VTAIL VN 1.16002f
C15 VTAIL w_n2212_n1208# 1.38949f
C16 VDD1 VP 0.913807f
C17 VP VN 3.578f
C18 B VTAIL 1.07936f
C19 VP w_n2212_n1208# 3.62808f
C20 VDD1 VDD2 0.817362f
C21 VDD2 VSUBS 0.517623f
C22 VDD1 VSUBS 2.82464f
C23 VTAIL VSUBS 0.338756f
C24 VN VSUBS 4.70754f
C25 VP VSUBS 1.282643f
C26 B VSUBS 2.478726f
C27 w_n2212_n1208# VSUBS 34.3745f
C28 VDD1.t1 VSUBS 0.019671f
C29 VDD1.t3 VSUBS 0.019671f
C30 VDD1.n0 VSUBS 0.064121f
C31 VDD1.t2 VSUBS 0.019671f
C32 VDD1.t0 VSUBS 0.019671f
C33 VDD1.n1 VSUBS 0.126311f
C34 VP.n0 VSUBS 0.057291f
C35 VP.t3 VSUBS 0.24212f
C36 VP.n1 VSUBS 0.046272f
C37 VP.n2 VSUBS 0.057291f
C38 VP.t1 VSUBS 0.24212f
C39 VP.t2 VSUBS 0.537839f
C40 VP.t0 VSUBS 0.534503f
C41 VP.n3 VSUBS 2.05353f
C42 VP.n4 VSUBS 2.26567f
C43 VP.n5 VSUBS 0.282509f
C44 VP.n6 VSUBS 0.057464f
C45 VP.n7 VSUBS 0.113266f
C46 VP.n8 VSUBS 0.057291f
C47 VP.n9 VSUBS 0.057291f
C48 VP.n10 VSUBS 0.057291f
C49 VP.n11 VSUBS 0.113266f
C50 VP.n12 VSUBS 0.057464f
C51 VP.n13 VSUBS 0.282509f
C52 VP.n14 VSUBS 0.061174f
C53 VTAIL.t7 VSUBS 0.092429f
C54 VTAIL.n0 VSUBS 0.247787f
C55 VTAIL.t0 VSUBS 0.092429f
C56 VTAIL.n1 VSUBS 0.300423f
C57 VTAIL.t2 VSUBS 0.092429f
C58 VTAIL.n2 VSUBS 0.714718f
C59 VTAIL.t5 VSUBS 0.092429f
C60 VTAIL.n3 VSUBS 0.714718f
C61 VTAIL.t6 VSUBS 0.092429f
C62 VTAIL.n4 VSUBS 0.300423f
C63 VTAIL.t3 VSUBS 0.092429f
C64 VTAIL.n5 VSUBS 0.300423f
C65 VTAIL.t1 VSUBS 0.092429f
C66 VTAIL.n6 VSUBS 0.714718f
C67 VTAIL.t4 VSUBS 0.092429f
C68 VTAIL.n7 VSUBS 0.654738f
C69 VDD2.t2 VSUBS 0.02032f
C70 VDD2.t0 VSUBS 0.02032f
C71 VDD2.n0 VSUBS 0.12594f
C72 VDD2.t3 VSUBS 0.02032f
C73 VDD2.t1 VSUBS 0.02032f
C74 VDD2.n1 VSUBS 0.066182f
C75 VDD2.n2 VSUBS 1.99877f
C76 VN.t0 VSUBS 0.517114f
C77 VN.t3 VSUBS 0.513908f
C78 VN.n0 VSUBS 0.363767f
C79 VN.t1 VSUBS 0.517114f
C80 VN.t2 VSUBS 0.513908f
C81 VN.n1 VSUBS 2.00698f
C82 B.n0 VSUBS 0.009027f
C83 B.n1 VSUBS 0.009027f
C84 B.n2 VSUBS 0.013351f
C85 B.n3 VSUBS 0.010231f
C86 B.n4 VSUBS 0.010231f
C87 B.n5 VSUBS 0.010231f
C88 B.n6 VSUBS 0.010231f
C89 B.n7 VSUBS 0.010231f
C90 B.n8 VSUBS 0.010231f
C91 B.n9 VSUBS 0.010231f
C92 B.n10 VSUBS 0.010231f
C93 B.n11 VSUBS 0.010231f
C94 B.n12 VSUBS 0.010231f
C95 B.n13 VSUBS 0.010231f
C96 B.n14 VSUBS 0.010231f
C97 B.n15 VSUBS 0.024232f
C98 B.n16 VSUBS 0.010231f
C99 B.n17 VSUBS 0.010231f
C100 B.n18 VSUBS 0.010231f
C101 B.n19 VSUBS 0.010231f
C102 B.t7 VSUBS 0.033083f
C103 B.t8 VSUBS 0.038325f
C104 B.t6 VSUBS 0.152963f
C105 B.n20 VSUBS 0.081013f
C106 B.n21 VSUBS 0.067506f
C107 B.n22 VSUBS 0.023704f
C108 B.n23 VSUBS 0.010231f
C109 B.n24 VSUBS 0.010231f
C110 B.n25 VSUBS 0.010231f
C111 B.n26 VSUBS 0.010231f
C112 B.n27 VSUBS 0.010231f
C113 B.t4 VSUBS 0.033083f
C114 B.t5 VSUBS 0.038325f
C115 B.t3 VSUBS 0.152963f
C116 B.n28 VSUBS 0.081013f
C117 B.n29 VSUBS 0.067506f
C118 B.n30 VSUBS 0.010231f
C119 B.n31 VSUBS 0.010231f
C120 B.n32 VSUBS 0.010231f
C121 B.n33 VSUBS 0.010231f
C122 B.n34 VSUBS 0.023612f
C123 B.n35 VSUBS 0.010231f
C124 B.n36 VSUBS 0.010231f
C125 B.n37 VSUBS 0.010231f
C126 B.n38 VSUBS 0.010231f
C127 B.n39 VSUBS 0.010231f
C128 B.n40 VSUBS 0.010231f
C129 B.n41 VSUBS 0.010231f
C130 B.n42 VSUBS 0.010231f
C131 B.n43 VSUBS 0.010231f
C132 B.n44 VSUBS 0.010231f
C133 B.n45 VSUBS 0.010231f
C134 B.n46 VSUBS 0.010231f
C135 B.n47 VSUBS 0.010231f
C136 B.n48 VSUBS 0.010231f
C137 B.n49 VSUBS 0.010231f
C138 B.n50 VSUBS 0.010231f
C139 B.n51 VSUBS 0.010231f
C140 B.n52 VSUBS 0.010231f
C141 B.n53 VSUBS 0.010231f
C142 B.n54 VSUBS 0.010231f
C143 B.n55 VSUBS 0.010231f
C144 B.n56 VSUBS 0.010231f
C145 B.n57 VSUBS 0.010231f
C146 B.n58 VSUBS 0.010231f
C147 B.n59 VSUBS 0.010231f
C148 B.n60 VSUBS 0.010231f
C149 B.n61 VSUBS 0.024232f
C150 B.n62 VSUBS 0.010231f
C151 B.n63 VSUBS 0.010231f
C152 B.n64 VSUBS 0.010231f
C153 B.n65 VSUBS 0.010231f
C154 B.t2 VSUBS 0.033083f
C155 B.t1 VSUBS 0.038325f
C156 B.t0 VSUBS 0.152963f
C157 B.n66 VSUBS 0.081013f
C158 B.n67 VSUBS 0.067506f
C159 B.n68 VSUBS 0.023704f
C160 B.n69 VSUBS 0.010231f
C161 B.n70 VSUBS 0.010231f
C162 B.n71 VSUBS 0.010231f
C163 B.n72 VSUBS 0.010231f
C164 B.n73 VSUBS 0.010231f
C165 B.t11 VSUBS 0.033083f
C166 B.t10 VSUBS 0.038325f
C167 B.t9 VSUBS 0.152963f
C168 B.n74 VSUBS 0.081013f
C169 B.n75 VSUBS 0.067506f
C170 B.n76 VSUBS 0.010231f
C171 B.n77 VSUBS 0.010231f
C172 B.n78 VSUBS 0.010231f
C173 B.n79 VSUBS 0.010231f
C174 B.n80 VSUBS 0.023612f
C175 B.n81 VSUBS 0.010231f
C176 B.n82 VSUBS 0.010231f
C177 B.n83 VSUBS 0.010231f
C178 B.n84 VSUBS 0.010231f
C179 B.n85 VSUBS 0.010231f
C180 B.n86 VSUBS 0.010231f
C181 B.n87 VSUBS 0.010231f
C182 B.n88 VSUBS 0.010231f
C183 B.n89 VSUBS 0.010231f
C184 B.n90 VSUBS 0.010231f
C185 B.n91 VSUBS 0.010231f
C186 B.n92 VSUBS 0.010231f
C187 B.n93 VSUBS 0.010231f
C188 B.n94 VSUBS 0.010231f
C189 B.n95 VSUBS 0.010231f
C190 B.n96 VSUBS 0.010231f
C191 B.n97 VSUBS 0.010231f
C192 B.n98 VSUBS 0.010231f
C193 B.n99 VSUBS 0.010231f
C194 B.n100 VSUBS 0.010231f
C195 B.n101 VSUBS 0.010231f
C196 B.n102 VSUBS 0.010231f
C197 B.n103 VSUBS 0.010231f
C198 B.n104 VSUBS 0.010231f
C199 B.n105 VSUBS 0.010231f
C200 B.n106 VSUBS 0.010231f
C201 B.n107 VSUBS 0.010231f
C202 B.n108 VSUBS 0.010231f
C203 B.n109 VSUBS 0.010231f
C204 B.n110 VSUBS 0.010231f
C205 B.n111 VSUBS 0.010231f
C206 B.n112 VSUBS 0.010231f
C207 B.n113 VSUBS 0.010231f
C208 B.n114 VSUBS 0.010231f
C209 B.n115 VSUBS 0.010231f
C210 B.n116 VSUBS 0.010231f
C211 B.n117 VSUBS 0.010231f
C212 B.n118 VSUBS 0.010231f
C213 B.n119 VSUBS 0.010231f
C214 B.n120 VSUBS 0.010231f
C215 B.n121 VSUBS 0.010231f
C216 B.n122 VSUBS 0.010231f
C217 B.n123 VSUBS 0.010231f
C218 B.n124 VSUBS 0.010231f
C219 B.n125 VSUBS 0.010231f
C220 B.n126 VSUBS 0.010231f
C221 B.n127 VSUBS 0.010231f
C222 B.n128 VSUBS 0.010231f
C223 B.n129 VSUBS 0.023612f
C224 B.n130 VSUBS 0.024232f
C225 B.n131 VSUBS 0.024232f
C226 B.n132 VSUBS 0.010231f
C227 B.n133 VSUBS 0.010231f
C228 B.n134 VSUBS 0.010231f
C229 B.n135 VSUBS 0.010231f
C230 B.n136 VSUBS 0.010231f
C231 B.n137 VSUBS 0.010231f
C232 B.n138 VSUBS 0.010231f
C233 B.n139 VSUBS 0.010231f
C234 B.n140 VSUBS 0.010231f
C235 B.n141 VSUBS 0.010231f
C236 B.n142 VSUBS 0.010231f
C237 B.n143 VSUBS 0.010231f
C238 B.n144 VSUBS 0.007071f
C239 B.n145 VSUBS 0.023704f
C240 B.n146 VSUBS 0.008275f
C241 B.n147 VSUBS 0.010231f
C242 B.n148 VSUBS 0.010231f
C243 B.n149 VSUBS 0.010231f
C244 B.n150 VSUBS 0.010231f
C245 B.n151 VSUBS 0.010231f
C246 B.n152 VSUBS 0.010231f
C247 B.n153 VSUBS 0.010231f
C248 B.n154 VSUBS 0.010231f
C249 B.n155 VSUBS 0.010231f
C250 B.n156 VSUBS 0.010231f
C251 B.n157 VSUBS 0.010231f
C252 B.n158 VSUBS 0.008275f
C253 B.n159 VSUBS 0.010231f
C254 B.n160 VSUBS 0.010231f
C255 B.n161 VSUBS 0.007071f
C256 B.n162 VSUBS 0.010231f
C257 B.n163 VSUBS 0.010231f
C258 B.n164 VSUBS 0.010231f
C259 B.n165 VSUBS 0.010231f
C260 B.n166 VSUBS 0.010231f
C261 B.n167 VSUBS 0.010231f
C262 B.n168 VSUBS 0.010231f
C263 B.n169 VSUBS 0.010231f
C264 B.n170 VSUBS 0.010231f
C265 B.n171 VSUBS 0.010231f
C266 B.n172 VSUBS 0.010231f
C267 B.n173 VSUBS 0.010231f
C268 B.n174 VSUBS 0.023022f
C269 B.n175 VSUBS 0.024823f
C270 B.n176 VSUBS 0.023612f
C271 B.n177 VSUBS 0.010231f
C272 B.n178 VSUBS 0.010231f
C273 B.n179 VSUBS 0.010231f
C274 B.n180 VSUBS 0.010231f
C275 B.n181 VSUBS 0.010231f
C276 B.n182 VSUBS 0.010231f
C277 B.n183 VSUBS 0.010231f
C278 B.n184 VSUBS 0.010231f
C279 B.n185 VSUBS 0.010231f
C280 B.n186 VSUBS 0.010231f
C281 B.n187 VSUBS 0.010231f
C282 B.n188 VSUBS 0.010231f
C283 B.n189 VSUBS 0.010231f
C284 B.n190 VSUBS 0.010231f
C285 B.n191 VSUBS 0.010231f
C286 B.n192 VSUBS 0.010231f
C287 B.n193 VSUBS 0.010231f
C288 B.n194 VSUBS 0.010231f
C289 B.n195 VSUBS 0.010231f
C290 B.n196 VSUBS 0.010231f
C291 B.n197 VSUBS 0.010231f
C292 B.n198 VSUBS 0.010231f
C293 B.n199 VSUBS 0.010231f
C294 B.n200 VSUBS 0.010231f
C295 B.n201 VSUBS 0.010231f
C296 B.n202 VSUBS 0.010231f
C297 B.n203 VSUBS 0.010231f
C298 B.n204 VSUBS 0.010231f
C299 B.n205 VSUBS 0.010231f
C300 B.n206 VSUBS 0.010231f
C301 B.n207 VSUBS 0.010231f
C302 B.n208 VSUBS 0.010231f
C303 B.n209 VSUBS 0.010231f
C304 B.n210 VSUBS 0.010231f
C305 B.n211 VSUBS 0.010231f
C306 B.n212 VSUBS 0.010231f
C307 B.n213 VSUBS 0.010231f
C308 B.n214 VSUBS 0.010231f
C309 B.n215 VSUBS 0.010231f
C310 B.n216 VSUBS 0.010231f
C311 B.n217 VSUBS 0.010231f
C312 B.n218 VSUBS 0.010231f
C313 B.n219 VSUBS 0.010231f
C314 B.n220 VSUBS 0.010231f
C315 B.n221 VSUBS 0.010231f
C316 B.n222 VSUBS 0.010231f
C317 B.n223 VSUBS 0.010231f
C318 B.n224 VSUBS 0.010231f
C319 B.n225 VSUBS 0.010231f
C320 B.n226 VSUBS 0.010231f
C321 B.n227 VSUBS 0.010231f
C322 B.n228 VSUBS 0.010231f
C323 B.n229 VSUBS 0.010231f
C324 B.n230 VSUBS 0.010231f
C325 B.n231 VSUBS 0.010231f
C326 B.n232 VSUBS 0.010231f
C327 B.n233 VSUBS 0.010231f
C328 B.n234 VSUBS 0.010231f
C329 B.n235 VSUBS 0.010231f
C330 B.n236 VSUBS 0.010231f
C331 B.n237 VSUBS 0.010231f
C332 B.n238 VSUBS 0.010231f
C333 B.n239 VSUBS 0.010231f
C334 B.n240 VSUBS 0.010231f
C335 B.n241 VSUBS 0.010231f
C336 B.n242 VSUBS 0.010231f
C337 B.n243 VSUBS 0.010231f
C338 B.n244 VSUBS 0.010231f
C339 B.n245 VSUBS 0.010231f
C340 B.n246 VSUBS 0.010231f
C341 B.n247 VSUBS 0.010231f
C342 B.n248 VSUBS 0.010231f
C343 B.n249 VSUBS 0.010231f
C344 B.n250 VSUBS 0.010231f
C345 B.n251 VSUBS 0.010231f
C346 B.n252 VSUBS 0.010231f
C347 B.n253 VSUBS 0.010231f
C348 B.n254 VSUBS 0.010231f
C349 B.n255 VSUBS 0.023612f
C350 B.n256 VSUBS 0.024232f
C351 B.n257 VSUBS 0.024232f
C352 B.n258 VSUBS 0.010231f
C353 B.n259 VSUBS 0.010231f
C354 B.n260 VSUBS 0.010231f
C355 B.n261 VSUBS 0.010231f
C356 B.n262 VSUBS 0.010231f
C357 B.n263 VSUBS 0.010231f
C358 B.n264 VSUBS 0.010231f
C359 B.n265 VSUBS 0.010231f
C360 B.n266 VSUBS 0.010231f
C361 B.n267 VSUBS 0.010231f
C362 B.n268 VSUBS 0.010231f
C363 B.n269 VSUBS 0.010231f
C364 B.n270 VSUBS 0.007071f
C365 B.n271 VSUBS 0.023704f
C366 B.n272 VSUBS 0.008275f
C367 B.n273 VSUBS 0.010231f
C368 B.n274 VSUBS 0.010231f
C369 B.n275 VSUBS 0.010231f
C370 B.n276 VSUBS 0.010231f
C371 B.n277 VSUBS 0.010231f
C372 B.n278 VSUBS 0.010231f
C373 B.n279 VSUBS 0.010231f
C374 B.n280 VSUBS 0.010231f
C375 B.n281 VSUBS 0.010231f
C376 B.n282 VSUBS 0.010231f
C377 B.n283 VSUBS 0.010231f
C378 B.n284 VSUBS 0.008275f
C379 B.n285 VSUBS 0.010231f
C380 B.n286 VSUBS 0.010231f
C381 B.n287 VSUBS 0.007071f
C382 B.n288 VSUBS 0.010231f
C383 B.n289 VSUBS 0.010231f
C384 B.n290 VSUBS 0.010231f
C385 B.n291 VSUBS 0.010231f
C386 B.n292 VSUBS 0.010231f
C387 B.n293 VSUBS 0.010231f
C388 B.n294 VSUBS 0.010231f
C389 B.n295 VSUBS 0.010231f
C390 B.n296 VSUBS 0.010231f
C391 B.n297 VSUBS 0.010231f
C392 B.n298 VSUBS 0.010231f
C393 B.n299 VSUBS 0.010231f
C394 B.n300 VSUBS 0.024232f
C395 B.n301 VSUBS 0.023612f
C396 B.n302 VSUBS 0.023612f
C397 B.n303 VSUBS 0.010231f
C398 B.n304 VSUBS 0.010231f
C399 B.n305 VSUBS 0.010231f
C400 B.n306 VSUBS 0.010231f
C401 B.n307 VSUBS 0.010231f
C402 B.n308 VSUBS 0.010231f
C403 B.n309 VSUBS 0.010231f
C404 B.n310 VSUBS 0.010231f
C405 B.n311 VSUBS 0.010231f
C406 B.n312 VSUBS 0.010231f
C407 B.n313 VSUBS 0.010231f
C408 B.n314 VSUBS 0.010231f
C409 B.n315 VSUBS 0.010231f
C410 B.n316 VSUBS 0.010231f
C411 B.n317 VSUBS 0.010231f
C412 B.n318 VSUBS 0.010231f
C413 B.n319 VSUBS 0.010231f
C414 B.n320 VSUBS 0.010231f
C415 B.n321 VSUBS 0.010231f
C416 B.n322 VSUBS 0.010231f
C417 B.n323 VSUBS 0.010231f
C418 B.n324 VSUBS 0.010231f
C419 B.n325 VSUBS 0.010231f
C420 B.n326 VSUBS 0.010231f
C421 B.n327 VSUBS 0.010231f
C422 B.n328 VSUBS 0.010231f
C423 B.n329 VSUBS 0.010231f
C424 B.n330 VSUBS 0.010231f
C425 B.n331 VSUBS 0.010231f
C426 B.n332 VSUBS 0.010231f
C427 B.n333 VSUBS 0.010231f
C428 B.n334 VSUBS 0.010231f
C429 B.n335 VSUBS 0.010231f
C430 B.n336 VSUBS 0.010231f
C431 B.n337 VSUBS 0.010231f
C432 B.n338 VSUBS 0.010231f
C433 B.n339 VSUBS 0.013351f
C434 B.n340 VSUBS 0.014222f
C435 B.n341 VSUBS 0.028282f
.ends

