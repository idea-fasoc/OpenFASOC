* NGSPICE file created from diff_pair_sample_1025.ext - technology: sky130A

.subckt diff_pair_sample_1025 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=3.1515 pd=19.43 as=3.1515 ps=19.43 w=19.1 l=3.87
X1 VDD2.t9 VN.t0 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=7.449 pd=38.98 as=3.1515 ps=19.43 w=19.1 l=3.87
X2 VDD2.t8 VN.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=3.1515 pd=19.43 as=7.449 ps=38.98 w=19.1 l=3.87
X3 VTAIL.t18 VP.t1 VDD1.t4 B.t9 sky130_fd_pr__nfet_01v8 ad=3.1515 pd=19.43 as=3.1515 ps=19.43 w=19.1 l=3.87
X4 VTAIL.t17 VP.t2 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.1515 pd=19.43 as=3.1515 ps=19.43 w=19.1 l=3.87
X5 VDD2.t7 VN.t2 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.1515 pd=19.43 as=3.1515 ps=19.43 w=19.1 l=3.87
X6 VTAIL.t3 VN.t3 VDD2.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=3.1515 pd=19.43 as=3.1515 ps=19.43 w=19.1 l=3.87
X7 VTAIL.t9 VN.t4 VDD2.t5 B.t9 sky130_fd_pr__nfet_01v8 ad=3.1515 pd=19.43 as=3.1515 ps=19.43 w=19.1 l=3.87
X8 VDD1.t2 VP.t3 VTAIL.t16 B.t6 sky130_fd_pr__nfet_01v8 ad=7.449 pd=38.98 as=3.1515 ps=19.43 w=19.1 l=3.87
X9 VDD1.t9 VP.t4 VTAIL.t15 B.t5 sky130_fd_pr__nfet_01v8 ad=3.1515 pd=19.43 as=7.449 ps=38.98 w=19.1 l=3.87
X10 VDD2.t4 VN.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.1515 pd=19.43 as=3.1515 ps=19.43 w=19.1 l=3.87
X11 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=7.449 pd=38.98 as=0 ps=0 w=19.1 l=3.87
X12 VDD1.t8 VP.t5 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=3.1515 pd=19.43 as=3.1515 ps=19.43 w=19.1 l=3.87
X13 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=7.449 pd=38.98 as=0 ps=0 w=19.1 l=3.87
X14 VTAIL.t0 VN.t6 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=3.1515 pd=19.43 as=3.1515 ps=19.43 w=19.1 l=3.87
X15 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=7.449 pd=38.98 as=0 ps=0 w=19.1 l=3.87
X16 VDD1.t7 VP.t6 VTAIL.t13 B.t4 sky130_fd_pr__nfet_01v8 ad=3.1515 pd=19.43 as=3.1515 ps=19.43 w=19.1 l=3.87
X17 VDD1.t6 VP.t7 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=7.449 pd=38.98 as=3.1515 ps=19.43 w=19.1 l=3.87
X18 VDD2.t2 VN.t7 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.1515 pd=19.43 as=7.449 ps=38.98 w=19.1 l=3.87
X19 VTAIL.t11 VP.t8 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=3.1515 pd=19.43 as=3.1515 ps=19.43 w=19.1 l=3.87
X20 VDD1.t0 VP.t9 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=3.1515 pd=19.43 as=7.449 ps=38.98 w=19.1 l=3.87
X21 VTAIL.t8 VN.t8 VDD2.t1 B.t8 sky130_fd_pr__nfet_01v8 ad=3.1515 pd=19.43 as=3.1515 ps=19.43 w=19.1 l=3.87
X22 VDD2.t0 VN.t9 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=7.449 pd=38.98 as=3.1515 ps=19.43 w=19.1 l=3.87
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.449 pd=38.98 as=0 ps=0 w=19.1 l=3.87
R0 VP.n32 VP.n29 161.3
R1 VP.n34 VP.n33 161.3
R2 VP.n35 VP.n28 161.3
R3 VP.n37 VP.n36 161.3
R4 VP.n38 VP.n27 161.3
R5 VP.n40 VP.n39 161.3
R6 VP.n41 VP.n26 161.3
R7 VP.n43 VP.n42 161.3
R8 VP.n44 VP.n25 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n47 VP.n24 161.3
R11 VP.n49 VP.n48 161.3
R12 VP.n50 VP.n23 161.3
R13 VP.n52 VP.n51 161.3
R14 VP.n53 VP.n22 161.3
R15 VP.n55 VP.n54 161.3
R16 VP.n56 VP.n21 161.3
R17 VP.n59 VP.n58 161.3
R18 VP.n60 VP.n20 161.3
R19 VP.n62 VP.n61 161.3
R20 VP.n63 VP.n19 161.3
R21 VP.n65 VP.n64 161.3
R22 VP.n66 VP.n18 161.3
R23 VP.n68 VP.n67 161.3
R24 VP.n69 VP.n17 161.3
R25 VP.n124 VP.n0 161.3
R26 VP.n123 VP.n122 161.3
R27 VP.n121 VP.n1 161.3
R28 VP.n120 VP.n119 161.3
R29 VP.n118 VP.n2 161.3
R30 VP.n117 VP.n116 161.3
R31 VP.n115 VP.n3 161.3
R32 VP.n114 VP.n113 161.3
R33 VP.n111 VP.n4 161.3
R34 VP.n110 VP.n109 161.3
R35 VP.n108 VP.n5 161.3
R36 VP.n107 VP.n106 161.3
R37 VP.n105 VP.n6 161.3
R38 VP.n104 VP.n103 161.3
R39 VP.n102 VP.n7 161.3
R40 VP.n101 VP.n100 161.3
R41 VP.n99 VP.n8 161.3
R42 VP.n98 VP.n97 161.3
R43 VP.n96 VP.n9 161.3
R44 VP.n95 VP.n94 161.3
R45 VP.n93 VP.n10 161.3
R46 VP.n92 VP.n91 161.3
R47 VP.n90 VP.n11 161.3
R48 VP.n89 VP.n88 161.3
R49 VP.n87 VP.n12 161.3
R50 VP.n85 VP.n84 161.3
R51 VP.n83 VP.n13 161.3
R52 VP.n82 VP.n81 161.3
R53 VP.n80 VP.n14 161.3
R54 VP.n79 VP.n78 161.3
R55 VP.n77 VP.n15 161.3
R56 VP.n76 VP.n75 161.3
R57 VP.n74 VP.n16 161.3
R58 VP.n30 VP.t7 151.149
R59 VP.n99 VP.t6 118.944
R60 VP.n73 VP.t3 118.944
R61 VP.n86 VP.t8 118.944
R62 VP.n112 VP.t1 118.944
R63 VP.n125 VP.t9 118.944
R64 VP.n44 VP.t5 118.944
R65 VP.n70 VP.t4 118.944
R66 VP.n57 VP.t0 118.944
R67 VP.n31 VP.t2 118.944
R68 VP.n72 VP.n71 65.602
R69 VP.n31 VP.n30 65.0774
R70 VP.n73 VP.n72 62.5108
R71 VP.n126 VP.n125 62.5108
R72 VP.n71 VP.n70 62.5108
R73 VP.n80 VP.n79 56.4773
R74 VP.n119 VP.n118 56.4773
R75 VP.n64 VP.n63 56.4773
R76 VP.n93 VP.n92 50.148
R77 VP.n106 VP.n105 50.148
R78 VP.n51 VP.n50 50.148
R79 VP.n38 VP.n37 50.148
R80 VP.n94 VP.n93 30.6732
R81 VP.n105 VP.n104 30.6732
R82 VP.n50 VP.n49 30.6732
R83 VP.n39 VP.n38 30.6732
R84 VP.n75 VP.n74 24.3439
R85 VP.n75 VP.n15 24.3439
R86 VP.n79 VP.n15 24.3439
R87 VP.n81 VP.n80 24.3439
R88 VP.n81 VP.n13 24.3439
R89 VP.n85 VP.n13 24.3439
R90 VP.n88 VP.n87 24.3439
R91 VP.n88 VP.n11 24.3439
R92 VP.n92 VP.n11 24.3439
R93 VP.n94 VP.n9 24.3439
R94 VP.n98 VP.n9 24.3439
R95 VP.n99 VP.n98 24.3439
R96 VP.n100 VP.n99 24.3439
R97 VP.n100 VP.n7 24.3439
R98 VP.n104 VP.n7 24.3439
R99 VP.n106 VP.n5 24.3439
R100 VP.n110 VP.n5 24.3439
R101 VP.n111 VP.n110 24.3439
R102 VP.n113 VP.n3 24.3439
R103 VP.n117 VP.n3 24.3439
R104 VP.n118 VP.n117 24.3439
R105 VP.n119 VP.n1 24.3439
R106 VP.n123 VP.n1 24.3439
R107 VP.n124 VP.n123 24.3439
R108 VP.n64 VP.n18 24.3439
R109 VP.n68 VP.n18 24.3439
R110 VP.n69 VP.n68 24.3439
R111 VP.n51 VP.n22 24.3439
R112 VP.n55 VP.n22 24.3439
R113 VP.n56 VP.n55 24.3439
R114 VP.n58 VP.n20 24.3439
R115 VP.n62 VP.n20 24.3439
R116 VP.n63 VP.n62 24.3439
R117 VP.n39 VP.n26 24.3439
R118 VP.n43 VP.n26 24.3439
R119 VP.n44 VP.n43 24.3439
R120 VP.n45 VP.n44 24.3439
R121 VP.n45 VP.n24 24.3439
R122 VP.n49 VP.n24 24.3439
R123 VP.n33 VP.n32 24.3439
R124 VP.n33 VP.n28 24.3439
R125 VP.n37 VP.n28 24.3439
R126 VP.n74 VP.n73 19.4752
R127 VP.n125 VP.n124 19.4752
R128 VP.n70 VP.n69 19.4752
R129 VP.n86 VP.n85 14.6066
R130 VP.n113 VP.n112 14.6066
R131 VP.n58 VP.n57 14.6066
R132 VP.n87 VP.n86 9.73787
R133 VP.n112 VP.n111 9.73787
R134 VP.n57 VP.n56 9.73787
R135 VP.n32 VP.n31 9.73787
R136 VP.n30 VP.n29 2.72002
R137 VP.n71 VP.n17 0.417764
R138 VP.n72 VP.n16 0.417764
R139 VP.n126 VP.n0 0.417764
R140 VP VP.n126 0.394061
R141 VP.n34 VP.n29 0.189894
R142 VP.n35 VP.n34 0.189894
R143 VP.n36 VP.n35 0.189894
R144 VP.n36 VP.n27 0.189894
R145 VP.n40 VP.n27 0.189894
R146 VP.n41 VP.n40 0.189894
R147 VP.n42 VP.n41 0.189894
R148 VP.n42 VP.n25 0.189894
R149 VP.n46 VP.n25 0.189894
R150 VP.n47 VP.n46 0.189894
R151 VP.n48 VP.n47 0.189894
R152 VP.n48 VP.n23 0.189894
R153 VP.n52 VP.n23 0.189894
R154 VP.n53 VP.n52 0.189894
R155 VP.n54 VP.n53 0.189894
R156 VP.n54 VP.n21 0.189894
R157 VP.n59 VP.n21 0.189894
R158 VP.n60 VP.n59 0.189894
R159 VP.n61 VP.n60 0.189894
R160 VP.n61 VP.n19 0.189894
R161 VP.n65 VP.n19 0.189894
R162 VP.n66 VP.n65 0.189894
R163 VP.n67 VP.n66 0.189894
R164 VP.n67 VP.n17 0.189894
R165 VP.n76 VP.n16 0.189894
R166 VP.n77 VP.n76 0.189894
R167 VP.n78 VP.n77 0.189894
R168 VP.n78 VP.n14 0.189894
R169 VP.n82 VP.n14 0.189894
R170 VP.n83 VP.n82 0.189894
R171 VP.n84 VP.n83 0.189894
R172 VP.n84 VP.n12 0.189894
R173 VP.n89 VP.n12 0.189894
R174 VP.n90 VP.n89 0.189894
R175 VP.n91 VP.n90 0.189894
R176 VP.n91 VP.n10 0.189894
R177 VP.n95 VP.n10 0.189894
R178 VP.n96 VP.n95 0.189894
R179 VP.n97 VP.n96 0.189894
R180 VP.n97 VP.n8 0.189894
R181 VP.n101 VP.n8 0.189894
R182 VP.n102 VP.n101 0.189894
R183 VP.n103 VP.n102 0.189894
R184 VP.n103 VP.n6 0.189894
R185 VP.n107 VP.n6 0.189894
R186 VP.n108 VP.n107 0.189894
R187 VP.n109 VP.n108 0.189894
R188 VP.n109 VP.n4 0.189894
R189 VP.n114 VP.n4 0.189894
R190 VP.n115 VP.n114 0.189894
R191 VP.n116 VP.n115 0.189894
R192 VP.n116 VP.n2 0.189894
R193 VP.n120 VP.n2 0.189894
R194 VP.n121 VP.n120 0.189894
R195 VP.n122 VP.n121 0.189894
R196 VP.n122 VP.n0 0.189894
R197 VDD1.n1 VDD1.t6 67.572
R198 VDD1.n3 VDD1.t2 67.5719
R199 VDD1.n5 VDD1.n4 65.5737
R200 VDD1.n1 VDD1.n0 62.9147
R201 VDD1.n7 VDD1.n6 62.9145
R202 VDD1.n3 VDD1.n2 62.9135
R203 VDD1.n7 VDD1.n5 59.7724
R204 VDD1 VDD1.n7 2.65783
R205 VDD1.n6 VDD1.t5 1.03715
R206 VDD1.n6 VDD1.t9 1.03715
R207 VDD1.n0 VDD1.t3 1.03715
R208 VDD1.n0 VDD1.t8 1.03715
R209 VDD1.n4 VDD1.t4 1.03715
R210 VDD1.n4 VDD1.t0 1.03715
R211 VDD1.n2 VDD1.t1 1.03715
R212 VDD1.n2 VDD1.t7 1.03715
R213 VDD1 VDD1.n1 0.963862
R214 VDD1.n5 VDD1.n3 0.850326
R215 VTAIL.n11 VTAIL.t2 47.2725
R216 VTAIL.n17 VTAIL.t5 47.2724
R217 VTAIL.n2 VTAIL.t10 47.2724
R218 VTAIL.n16 VTAIL.t15 47.2724
R219 VTAIL.n15 VTAIL.n14 46.2359
R220 VTAIL.n13 VTAIL.n12 46.2359
R221 VTAIL.n10 VTAIL.n9 46.2359
R222 VTAIL.n8 VTAIL.n7 46.2359
R223 VTAIL.n19 VTAIL.n18 46.2347
R224 VTAIL.n1 VTAIL.n0 46.2347
R225 VTAIL.n4 VTAIL.n3 46.2347
R226 VTAIL.n6 VTAIL.n5 46.2347
R227 VTAIL.n8 VTAIL.n6 36.0738
R228 VTAIL.n17 VTAIL.n16 32.4531
R229 VTAIL.n10 VTAIL.n8 3.62119
R230 VTAIL.n11 VTAIL.n10 3.62119
R231 VTAIL.n15 VTAIL.n13 3.62119
R232 VTAIL.n16 VTAIL.n15 3.62119
R233 VTAIL.n6 VTAIL.n4 3.62119
R234 VTAIL.n4 VTAIL.n2 3.62119
R235 VTAIL.n19 VTAIL.n17 3.62119
R236 VTAIL VTAIL.n1 2.77421
R237 VTAIL.n13 VTAIL.n11 2.28067
R238 VTAIL.n2 VTAIL.n1 2.28067
R239 VTAIL.n18 VTAIL.t1 1.03715
R240 VTAIL.n18 VTAIL.t8 1.03715
R241 VTAIL.n0 VTAIL.t7 1.03715
R242 VTAIL.n0 VTAIL.t3 1.03715
R243 VTAIL.n3 VTAIL.t13 1.03715
R244 VTAIL.n3 VTAIL.t18 1.03715
R245 VTAIL.n5 VTAIL.t16 1.03715
R246 VTAIL.n5 VTAIL.t11 1.03715
R247 VTAIL.n14 VTAIL.t14 1.03715
R248 VTAIL.n14 VTAIL.t19 1.03715
R249 VTAIL.n12 VTAIL.t12 1.03715
R250 VTAIL.n12 VTAIL.t17 1.03715
R251 VTAIL.n9 VTAIL.t4 1.03715
R252 VTAIL.n9 VTAIL.t9 1.03715
R253 VTAIL.n7 VTAIL.t6 1.03715
R254 VTAIL.n7 VTAIL.t0 1.03715
R255 VTAIL VTAIL.n19 0.847483
R256 B.n1076 B.n1075 585
R257 B.n1076 B.n148 585
R258 B.n1079 B.n1078 585
R259 B.n1080 B.n220 585
R260 B.n1082 B.n1081 585
R261 B.n1084 B.n219 585
R262 B.n1087 B.n1086 585
R263 B.n1088 B.n218 585
R264 B.n1090 B.n1089 585
R265 B.n1092 B.n217 585
R266 B.n1095 B.n1094 585
R267 B.n1096 B.n216 585
R268 B.n1098 B.n1097 585
R269 B.n1100 B.n215 585
R270 B.n1103 B.n1102 585
R271 B.n1104 B.n214 585
R272 B.n1106 B.n1105 585
R273 B.n1108 B.n213 585
R274 B.n1111 B.n1110 585
R275 B.n1112 B.n212 585
R276 B.n1114 B.n1113 585
R277 B.n1116 B.n211 585
R278 B.n1119 B.n1118 585
R279 B.n1120 B.n210 585
R280 B.n1122 B.n1121 585
R281 B.n1124 B.n209 585
R282 B.n1127 B.n1126 585
R283 B.n1128 B.n208 585
R284 B.n1130 B.n1129 585
R285 B.n1132 B.n207 585
R286 B.n1135 B.n1134 585
R287 B.n1136 B.n206 585
R288 B.n1138 B.n1137 585
R289 B.n1140 B.n205 585
R290 B.n1143 B.n1142 585
R291 B.n1144 B.n204 585
R292 B.n1146 B.n1145 585
R293 B.n1148 B.n203 585
R294 B.n1151 B.n1150 585
R295 B.n1152 B.n202 585
R296 B.n1154 B.n1153 585
R297 B.n1156 B.n201 585
R298 B.n1159 B.n1158 585
R299 B.n1160 B.n200 585
R300 B.n1162 B.n1161 585
R301 B.n1164 B.n199 585
R302 B.n1167 B.n1166 585
R303 B.n1168 B.n198 585
R304 B.n1170 B.n1169 585
R305 B.n1172 B.n197 585
R306 B.n1175 B.n1174 585
R307 B.n1176 B.n196 585
R308 B.n1178 B.n1177 585
R309 B.n1180 B.n195 585
R310 B.n1183 B.n1182 585
R311 B.n1184 B.n194 585
R312 B.n1186 B.n1185 585
R313 B.n1188 B.n193 585
R314 B.n1191 B.n1190 585
R315 B.n1192 B.n192 585
R316 B.n1194 B.n1193 585
R317 B.n1196 B.n191 585
R318 B.n1199 B.n1198 585
R319 B.n1200 B.n188 585
R320 B.n1203 B.n1202 585
R321 B.n1205 B.n187 585
R322 B.n1208 B.n1207 585
R323 B.n1209 B.n186 585
R324 B.n1211 B.n1210 585
R325 B.n1213 B.n185 585
R326 B.n1216 B.n1215 585
R327 B.n1217 B.n181 585
R328 B.n1219 B.n1218 585
R329 B.n1221 B.n180 585
R330 B.n1224 B.n1223 585
R331 B.n1225 B.n179 585
R332 B.n1227 B.n1226 585
R333 B.n1229 B.n178 585
R334 B.n1232 B.n1231 585
R335 B.n1233 B.n177 585
R336 B.n1235 B.n1234 585
R337 B.n1237 B.n176 585
R338 B.n1240 B.n1239 585
R339 B.n1241 B.n175 585
R340 B.n1243 B.n1242 585
R341 B.n1245 B.n174 585
R342 B.n1248 B.n1247 585
R343 B.n1249 B.n173 585
R344 B.n1251 B.n1250 585
R345 B.n1253 B.n172 585
R346 B.n1256 B.n1255 585
R347 B.n1257 B.n171 585
R348 B.n1259 B.n1258 585
R349 B.n1261 B.n170 585
R350 B.n1264 B.n1263 585
R351 B.n1265 B.n169 585
R352 B.n1267 B.n1266 585
R353 B.n1269 B.n168 585
R354 B.n1272 B.n1271 585
R355 B.n1273 B.n167 585
R356 B.n1275 B.n1274 585
R357 B.n1277 B.n166 585
R358 B.n1280 B.n1279 585
R359 B.n1281 B.n165 585
R360 B.n1283 B.n1282 585
R361 B.n1285 B.n164 585
R362 B.n1288 B.n1287 585
R363 B.n1289 B.n163 585
R364 B.n1291 B.n1290 585
R365 B.n1293 B.n162 585
R366 B.n1296 B.n1295 585
R367 B.n1297 B.n161 585
R368 B.n1299 B.n1298 585
R369 B.n1301 B.n160 585
R370 B.n1304 B.n1303 585
R371 B.n1305 B.n159 585
R372 B.n1307 B.n1306 585
R373 B.n1309 B.n158 585
R374 B.n1312 B.n1311 585
R375 B.n1313 B.n157 585
R376 B.n1315 B.n1314 585
R377 B.n1317 B.n156 585
R378 B.n1320 B.n1319 585
R379 B.n1321 B.n155 585
R380 B.n1323 B.n1322 585
R381 B.n1325 B.n154 585
R382 B.n1328 B.n1327 585
R383 B.n1329 B.n153 585
R384 B.n1331 B.n1330 585
R385 B.n1333 B.n152 585
R386 B.n1336 B.n1335 585
R387 B.n1337 B.n151 585
R388 B.n1339 B.n1338 585
R389 B.n1341 B.n150 585
R390 B.n1344 B.n1343 585
R391 B.n1345 B.n149 585
R392 B.n1074 B.n147 585
R393 B.n1348 B.n147 585
R394 B.n1073 B.n146 585
R395 B.n1349 B.n146 585
R396 B.n1072 B.n145 585
R397 B.n1350 B.n145 585
R398 B.n1071 B.n1070 585
R399 B.n1070 B.n141 585
R400 B.n1069 B.n140 585
R401 B.n1356 B.n140 585
R402 B.n1068 B.n139 585
R403 B.n1357 B.n139 585
R404 B.n1067 B.n138 585
R405 B.n1358 B.n138 585
R406 B.n1066 B.n1065 585
R407 B.n1065 B.n134 585
R408 B.n1064 B.n133 585
R409 B.n1364 B.n133 585
R410 B.n1063 B.n132 585
R411 B.n1365 B.n132 585
R412 B.n1062 B.n131 585
R413 B.n1366 B.n131 585
R414 B.n1061 B.n1060 585
R415 B.n1060 B.n127 585
R416 B.n1059 B.n126 585
R417 B.n1372 B.n126 585
R418 B.n1058 B.n125 585
R419 B.n1373 B.n125 585
R420 B.n1057 B.n124 585
R421 B.n1374 B.n124 585
R422 B.n1056 B.n1055 585
R423 B.n1055 B.n120 585
R424 B.n1054 B.n119 585
R425 B.n1380 B.n119 585
R426 B.n1053 B.n118 585
R427 B.n1381 B.n118 585
R428 B.n1052 B.n117 585
R429 B.n1382 B.n117 585
R430 B.n1051 B.n1050 585
R431 B.n1050 B.n113 585
R432 B.n1049 B.n112 585
R433 B.n1388 B.n112 585
R434 B.n1048 B.n111 585
R435 B.n1389 B.n111 585
R436 B.n1047 B.n110 585
R437 B.n1390 B.n110 585
R438 B.n1046 B.n1045 585
R439 B.n1045 B.n106 585
R440 B.n1044 B.n105 585
R441 B.n1396 B.n105 585
R442 B.n1043 B.n104 585
R443 B.n1397 B.n104 585
R444 B.n1042 B.n103 585
R445 B.n1398 B.n103 585
R446 B.n1041 B.n1040 585
R447 B.n1040 B.n99 585
R448 B.n1039 B.n98 585
R449 B.n1404 B.n98 585
R450 B.n1038 B.n97 585
R451 B.n1405 B.n97 585
R452 B.n1037 B.n96 585
R453 B.n1406 B.n96 585
R454 B.n1036 B.n1035 585
R455 B.n1035 B.n92 585
R456 B.n1034 B.n91 585
R457 B.n1412 B.n91 585
R458 B.n1033 B.n90 585
R459 B.n1413 B.n90 585
R460 B.n1032 B.n89 585
R461 B.n1414 B.n89 585
R462 B.n1031 B.n1030 585
R463 B.n1030 B.n85 585
R464 B.n1029 B.n84 585
R465 B.n1420 B.n84 585
R466 B.n1028 B.n83 585
R467 B.n1421 B.n83 585
R468 B.n1027 B.n82 585
R469 B.n1422 B.n82 585
R470 B.n1026 B.n1025 585
R471 B.n1025 B.n78 585
R472 B.n1024 B.n77 585
R473 B.n1428 B.n77 585
R474 B.n1023 B.n76 585
R475 B.n1429 B.n76 585
R476 B.n1022 B.n75 585
R477 B.n1430 B.n75 585
R478 B.n1021 B.n1020 585
R479 B.n1020 B.n71 585
R480 B.n1019 B.n70 585
R481 B.n1436 B.n70 585
R482 B.n1018 B.n69 585
R483 B.n1437 B.n69 585
R484 B.n1017 B.n68 585
R485 B.n1438 B.n68 585
R486 B.n1016 B.n1015 585
R487 B.n1015 B.n64 585
R488 B.n1014 B.n63 585
R489 B.n1444 B.n63 585
R490 B.n1013 B.n62 585
R491 B.n1445 B.n62 585
R492 B.n1012 B.n61 585
R493 B.n1446 B.n61 585
R494 B.n1011 B.n1010 585
R495 B.n1010 B.n57 585
R496 B.n1009 B.n56 585
R497 B.n1452 B.n56 585
R498 B.n1008 B.n55 585
R499 B.n1453 B.n55 585
R500 B.n1007 B.n54 585
R501 B.n1454 B.n54 585
R502 B.n1006 B.n1005 585
R503 B.n1005 B.n50 585
R504 B.n1004 B.n49 585
R505 B.n1460 B.n49 585
R506 B.n1003 B.n48 585
R507 B.n1461 B.n48 585
R508 B.n1002 B.n47 585
R509 B.n1462 B.n47 585
R510 B.n1001 B.n1000 585
R511 B.n1000 B.n43 585
R512 B.n999 B.n42 585
R513 B.n1468 B.n42 585
R514 B.n998 B.n41 585
R515 B.n1469 B.n41 585
R516 B.n997 B.n40 585
R517 B.n1470 B.n40 585
R518 B.n996 B.n995 585
R519 B.n995 B.n36 585
R520 B.n994 B.n35 585
R521 B.n1476 B.n35 585
R522 B.n993 B.n34 585
R523 B.n1477 B.n34 585
R524 B.n992 B.n33 585
R525 B.n1478 B.n33 585
R526 B.n991 B.n990 585
R527 B.n990 B.n29 585
R528 B.n989 B.n28 585
R529 B.n1484 B.n28 585
R530 B.n988 B.n27 585
R531 B.n1485 B.n27 585
R532 B.n987 B.n26 585
R533 B.n1486 B.n26 585
R534 B.n986 B.n985 585
R535 B.n985 B.n22 585
R536 B.n984 B.n21 585
R537 B.n1492 B.n21 585
R538 B.n983 B.n20 585
R539 B.n1493 B.n20 585
R540 B.n982 B.n19 585
R541 B.n1494 B.n19 585
R542 B.n981 B.n980 585
R543 B.n980 B.n15 585
R544 B.n979 B.n14 585
R545 B.n1500 B.n14 585
R546 B.n978 B.n13 585
R547 B.n1501 B.n13 585
R548 B.n977 B.n12 585
R549 B.n1502 B.n12 585
R550 B.n976 B.n975 585
R551 B.n975 B.n8 585
R552 B.n974 B.n7 585
R553 B.n1508 B.n7 585
R554 B.n973 B.n6 585
R555 B.n1509 B.n6 585
R556 B.n972 B.n5 585
R557 B.n1510 B.n5 585
R558 B.n971 B.n970 585
R559 B.n970 B.n4 585
R560 B.n969 B.n221 585
R561 B.n969 B.n968 585
R562 B.n959 B.n222 585
R563 B.n223 B.n222 585
R564 B.n961 B.n960 585
R565 B.n962 B.n961 585
R566 B.n958 B.n228 585
R567 B.n228 B.n227 585
R568 B.n957 B.n956 585
R569 B.n956 B.n955 585
R570 B.n230 B.n229 585
R571 B.n231 B.n230 585
R572 B.n948 B.n947 585
R573 B.n949 B.n948 585
R574 B.n946 B.n236 585
R575 B.n236 B.n235 585
R576 B.n945 B.n944 585
R577 B.n944 B.n943 585
R578 B.n238 B.n237 585
R579 B.n239 B.n238 585
R580 B.n936 B.n935 585
R581 B.n937 B.n936 585
R582 B.n934 B.n244 585
R583 B.n244 B.n243 585
R584 B.n933 B.n932 585
R585 B.n932 B.n931 585
R586 B.n246 B.n245 585
R587 B.n247 B.n246 585
R588 B.n924 B.n923 585
R589 B.n925 B.n924 585
R590 B.n922 B.n252 585
R591 B.n252 B.n251 585
R592 B.n921 B.n920 585
R593 B.n920 B.n919 585
R594 B.n254 B.n253 585
R595 B.n255 B.n254 585
R596 B.n912 B.n911 585
R597 B.n913 B.n912 585
R598 B.n910 B.n259 585
R599 B.n263 B.n259 585
R600 B.n909 B.n908 585
R601 B.n908 B.n907 585
R602 B.n261 B.n260 585
R603 B.n262 B.n261 585
R604 B.n900 B.n899 585
R605 B.n901 B.n900 585
R606 B.n898 B.n268 585
R607 B.n268 B.n267 585
R608 B.n897 B.n896 585
R609 B.n896 B.n895 585
R610 B.n270 B.n269 585
R611 B.n271 B.n270 585
R612 B.n888 B.n887 585
R613 B.n889 B.n888 585
R614 B.n886 B.n276 585
R615 B.n276 B.n275 585
R616 B.n885 B.n884 585
R617 B.n884 B.n883 585
R618 B.n278 B.n277 585
R619 B.n279 B.n278 585
R620 B.n876 B.n875 585
R621 B.n877 B.n876 585
R622 B.n874 B.n283 585
R623 B.n287 B.n283 585
R624 B.n873 B.n872 585
R625 B.n872 B.n871 585
R626 B.n285 B.n284 585
R627 B.n286 B.n285 585
R628 B.n864 B.n863 585
R629 B.n865 B.n864 585
R630 B.n862 B.n292 585
R631 B.n292 B.n291 585
R632 B.n861 B.n860 585
R633 B.n860 B.n859 585
R634 B.n294 B.n293 585
R635 B.n295 B.n294 585
R636 B.n852 B.n851 585
R637 B.n853 B.n852 585
R638 B.n850 B.n300 585
R639 B.n300 B.n299 585
R640 B.n849 B.n848 585
R641 B.n848 B.n847 585
R642 B.n302 B.n301 585
R643 B.n303 B.n302 585
R644 B.n840 B.n839 585
R645 B.n841 B.n840 585
R646 B.n838 B.n307 585
R647 B.n311 B.n307 585
R648 B.n837 B.n836 585
R649 B.n836 B.n835 585
R650 B.n309 B.n308 585
R651 B.n310 B.n309 585
R652 B.n828 B.n827 585
R653 B.n829 B.n828 585
R654 B.n826 B.n316 585
R655 B.n316 B.n315 585
R656 B.n825 B.n824 585
R657 B.n824 B.n823 585
R658 B.n318 B.n317 585
R659 B.n319 B.n318 585
R660 B.n816 B.n815 585
R661 B.n817 B.n816 585
R662 B.n814 B.n324 585
R663 B.n324 B.n323 585
R664 B.n813 B.n812 585
R665 B.n812 B.n811 585
R666 B.n326 B.n325 585
R667 B.n327 B.n326 585
R668 B.n804 B.n803 585
R669 B.n805 B.n804 585
R670 B.n802 B.n332 585
R671 B.n332 B.n331 585
R672 B.n801 B.n800 585
R673 B.n800 B.n799 585
R674 B.n334 B.n333 585
R675 B.n335 B.n334 585
R676 B.n792 B.n791 585
R677 B.n793 B.n792 585
R678 B.n790 B.n340 585
R679 B.n340 B.n339 585
R680 B.n789 B.n788 585
R681 B.n788 B.n787 585
R682 B.n342 B.n341 585
R683 B.n343 B.n342 585
R684 B.n780 B.n779 585
R685 B.n781 B.n780 585
R686 B.n778 B.n348 585
R687 B.n348 B.n347 585
R688 B.n777 B.n776 585
R689 B.n776 B.n775 585
R690 B.n350 B.n349 585
R691 B.n351 B.n350 585
R692 B.n768 B.n767 585
R693 B.n769 B.n768 585
R694 B.n766 B.n356 585
R695 B.n356 B.n355 585
R696 B.n765 B.n764 585
R697 B.n764 B.n763 585
R698 B.n358 B.n357 585
R699 B.n359 B.n358 585
R700 B.n756 B.n755 585
R701 B.n757 B.n756 585
R702 B.n754 B.n363 585
R703 B.n367 B.n363 585
R704 B.n753 B.n752 585
R705 B.n752 B.n751 585
R706 B.n365 B.n364 585
R707 B.n366 B.n365 585
R708 B.n744 B.n743 585
R709 B.n745 B.n744 585
R710 B.n742 B.n372 585
R711 B.n372 B.n371 585
R712 B.n741 B.n740 585
R713 B.n740 B.n739 585
R714 B.n374 B.n373 585
R715 B.n375 B.n374 585
R716 B.n732 B.n731 585
R717 B.n733 B.n732 585
R718 B.n730 B.n380 585
R719 B.n380 B.n379 585
R720 B.n729 B.n728 585
R721 B.n728 B.n727 585
R722 B.n724 B.n384 585
R723 B.n723 B.n722 585
R724 B.n720 B.n385 585
R725 B.n720 B.n383 585
R726 B.n719 B.n718 585
R727 B.n717 B.n716 585
R728 B.n715 B.n387 585
R729 B.n713 B.n712 585
R730 B.n711 B.n388 585
R731 B.n710 B.n709 585
R732 B.n707 B.n389 585
R733 B.n705 B.n704 585
R734 B.n703 B.n390 585
R735 B.n702 B.n701 585
R736 B.n699 B.n391 585
R737 B.n697 B.n696 585
R738 B.n695 B.n392 585
R739 B.n694 B.n693 585
R740 B.n691 B.n393 585
R741 B.n689 B.n688 585
R742 B.n687 B.n394 585
R743 B.n686 B.n685 585
R744 B.n683 B.n395 585
R745 B.n681 B.n680 585
R746 B.n679 B.n396 585
R747 B.n678 B.n677 585
R748 B.n675 B.n397 585
R749 B.n673 B.n672 585
R750 B.n671 B.n398 585
R751 B.n670 B.n669 585
R752 B.n667 B.n399 585
R753 B.n665 B.n664 585
R754 B.n663 B.n400 585
R755 B.n662 B.n661 585
R756 B.n659 B.n401 585
R757 B.n657 B.n656 585
R758 B.n655 B.n402 585
R759 B.n654 B.n653 585
R760 B.n651 B.n403 585
R761 B.n649 B.n648 585
R762 B.n647 B.n404 585
R763 B.n646 B.n645 585
R764 B.n643 B.n405 585
R765 B.n641 B.n640 585
R766 B.n639 B.n406 585
R767 B.n638 B.n637 585
R768 B.n635 B.n407 585
R769 B.n633 B.n632 585
R770 B.n631 B.n408 585
R771 B.n630 B.n629 585
R772 B.n627 B.n409 585
R773 B.n625 B.n624 585
R774 B.n623 B.n410 585
R775 B.n622 B.n621 585
R776 B.n619 B.n411 585
R777 B.n617 B.n616 585
R778 B.n615 B.n412 585
R779 B.n614 B.n613 585
R780 B.n611 B.n413 585
R781 B.n609 B.n608 585
R782 B.n607 B.n414 585
R783 B.n606 B.n605 585
R784 B.n603 B.n415 585
R785 B.n601 B.n600 585
R786 B.n598 B.n416 585
R787 B.n597 B.n596 585
R788 B.n594 B.n419 585
R789 B.n592 B.n591 585
R790 B.n590 B.n420 585
R791 B.n589 B.n588 585
R792 B.n586 B.n421 585
R793 B.n584 B.n583 585
R794 B.n582 B.n422 585
R795 B.n580 B.n579 585
R796 B.n577 B.n425 585
R797 B.n575 B.n574 585
R798 B.n573 B.n426 585
R799 B.n572 B.n571 585
R800 B.n569 B.n427 585
R801 B.n567 B.n566 585
R802 B.n565 B.n428 585
R803 B.n564 B.n563 585
R804 B.n561 B.n429 585
R805 B.n559 B.n558 585
R806 B.n557 B.n430 585
R807 B.n556 B.n555 585
R808 B.n553 B.n431 585
R809 B.n551 B.n550 585
R810 B.n549 B.n432 585
R811 B.n548 B.n547 585
R812 B.n545 B.n433 585
R813 B.n543 B.n542 585
R814 B.n541 B.n434 585
R815 B.n540 B.n539 585
R816 B.n537 B.n435 585
R817 B.n535 B.n534 585
R818 B.n533 B.n436 585
R819 B.n532 B.n531 585
R820 B.n529 B.n437 585
R821 B.n527 B.n526 585
R822 B.n525 B.n438 585
R823 B.n524 B.n523 585
R824 B.n521 B.n439 585
R825 B.n519 B.n518 585
R826 B.n517 B.n440 585
R827 B.n516 B.n515 585
R828 B.n513 B.n441 585
R829 B.n511 B.n510 585
R830 B.n509 B.n442 585
R831 B.n508 B.n507 585
R832 B.n505 B.n443 585
R833 B.n503 B.n502 585
R834 B.n501 B.n444 585
R835 B.n500 B.n499 585
R836 B.n497 B.n445 585
R837 B.n495 B.n494 585
R838 B.n493 B.n446 585
R839 B.n492 B.n491 585
R840 B.n489 B.n447 585
R841 B.n487 B.n486 585
R842 B.n485 B.n448 585
R843 B.n484 B.n483 585
R844 B.n481 B.n449 585
R845 B.n479 B.n478 585
R846 B.n477 B.n450 585
R847 B.n476 B.n475 585
R848 B.n473 B.n451 585
R849 B.n471 B.n470 585
R850 B.n469 B.n452 585
R851 B.n468 B.n467 585
R852 B.n465 B.n453 585
R853 B.n463 B.n462 585
R854 B.n461 B.n454 585
R855 B.n460 B.n459 585
R856 B.n457 B.n455 585
R857 B.n382 B.n381 585
R858 B.n726 B.n725 585
R859 B.n727 B.n726 585
R860 B.n378 B.n377 585
R861 B.n379 B.n378 585
R862 B.n735 B.n734 585
R863 B.n734 B.n733 585
R864 B.n736 B.n376 585
R865 B.n376 B.n375 585
R866 B.n738 B.n737 585
R867 B.n739 B.n738 585
R868 B.n370 B.n369 585
R869 B.n371 B.n370 585
R870 B.n747 B.n746 585
R871 B.n746 B.n745 585
R872 B.n748 B.n368 585
R873 B.n368 B.n366 585
R874 B.n750 B.n749 585
R875 B.n751 B.n750 585
R876 B.n362 B.n361 585
R877 B.n367 B.n362 585
R878 B.n759 B.n758 585
R879 B.n758 B.n757 585
R880 B.n760 B.n360 585
R881 B.n360 B.n359 585
R882 B.n762 B.n761 585
R883 B.n763 B.n762 585
R884 B.n354 B.n353 585
R885 B.n355 B.n354 585
R886 B.n771 B.n770 585
R887 B.n770 B.n769 585
R888 B.n772 B.n352 585
R889 B.n352 B.n351 585
R890 B.n774 B.n773 585
R891 B.n775 B.n774 585
R892 B.n346 B.n345 585
R893 B.n347 B.n346 585
R894 B.n783 B.n782 585
R895 B.n782 B.n781 585
R896 B.n784 B.n344 585
R897 B.n344 B.n343 585
R898 B.n786 B.n785 585
R899 B.n787 B.n786 585
R900 B.n338 B.n337 585
R901 B.n339 B.n338 585
R902 B.n795 B.n794 585
R903 B.n794 B.n793 585
R904 B.n796 B.n336 585
R905 B.n336 B.n335 585
R906 B.n798 B.n797 585
R907 B.n799 B.n798 585
R908 B.n330 B.n329 585
R909 B.n331 B.n330 585
R910 B.n807 B.n806 585
R911 B.n806 B.n805 585
R912 B.n808 B.n328 585
R913 B.n328 B.n327 585
R914 B.n810 B.n809 585
R915 B.n811 B.n810 585
R916 B.n322 B.n321 585
R917 B.n323 B.n322 585
R918 B.n819 B.n818 585
R919 B.n818 B.n817 585
R920 B.n820 B.n320 585
R921 B.n320 B.n319 585
R922 B.n822 B.n821 585
R923 B.n823 B.n822 585
R924 B.n314 B.n313 585
R925 B.n315 B.n314 585
R926 B.n831 B.n830 585
R927 B.n830 B.n829 585
R928 B.n832 B.n312 585
R929 B.n312 B.n310 585
R930 B.n834 B.n833 585
R931 B.n835 B.n834 585
R932 B.n306 B.n305 585
R933 B.n311 B.n306 585
R934 B.n843 B.n842 585
R935 B.n842 B.n841 585
R936 B.n844 B.n304 585
R937 B.n304 B.n303 585
R938 B.n846 B.n845 585
R939 B.n847 B.n846 585
R940 B.n298 B.n297 585
R941 B.n299 B.n298 585
R942 B.n855 B.n854 585
R943 B.n854 B.n853 585
R944 B.n856 B.n296 585
R945 B.n296 B.n295 585
R946 B.n858 B.n857 585
R947 B.n859 B.n858 585
R948 B.n290 B.n289 585
R949 B.n291 B.n290 585
R950 B.n867 B.n866 585
R951 B.n866 B.n865 585
R952 B.n868 B.n288 585
R953 B.n288 B.n286 585
R954 B.n870 B.n869 585
R955 B.n871 B.n870 585
R956 B.n282 B.n281 585
R957 B.n287 B.n282 585
R958 B.n879 B.n878 585
R959 B.n878 B.n877 585
R960 B.n880 B.n280 585
R961 B.n280 B.n279 585
R962 B.n882 B.n881 585
R963 B.n883 B.n882 585
R964 B.n274 B.n273 585
R965 B.n275 B.n274 585
R966 B.n891 B.n890 585
R967 B.n890 B.n889 585
R968 B.n892 B.n272 585
R969 B.n272 B.n271 585
R970 B.n894 B.n893 585
R971 B.n895 B.n894 585
R972 B.n266 B.n265 585
R973 B.n267 B.n266 585
R974 B.n903 B.n902 585
R975 B.n902 B.n901 585
R976 B.n904 B.n264 585
R977 B.n264 B.n262 585
R978 B.n906 B.n905 585
R979 B.n907 B.n906 585
R980 B.n258 B.n257 585
R981 B.n263 B.n258 585
R982 B.n915 B.n914 585
R983 B.n914 B.n913 585
R984 B.n916 B.n256 585
R985 B.n256 B.n255 585
R986 B.n918 B.n917 585
R987 B.n919 B.n918 585
R988 B.n250 B.n249 585
R989 B.n251 B.n250 585
R990 B.n927 B.n926 585
R991 B.n926 B.n925 585
R992 B.n928 B.n248 585
R993 B.n248 B.n247 585
R994 B.n930 B.n929 585
R995 B.n931 B.n930 585
R996 B.n242 B.n241 585
R997 B.n243 B.n242 585
R998 B.n939 B.n938 585
R999 B.n938 B.n937 585
R1000 B.n940 B.n240 585
R1001 B.n240 B.n239 585
R1002 B.n942 B.n941 585
R1003 B.n943 B.n942 585
R1004 B.n234 B.n233 585
R1005 B.n235 B.n234 585
R1006 B.n951 B.n950 585
R1007 B.n950 B.n949 585
R1008 B.n952 B.n232 585
R1009 B.n232 B.n231 585
R1010 B.n954 B.n953 585
R1011 B.n955 B.n954 585
R1012 B.n226 B.n225 585
R1013 B.n227 B.n226 585
R1014 B.n964 B.n963 585
R1015 B.n963 B.n962 585
R1016 B.n965 B.n224 585
R1017 B.n224 B.n223 585
R1018 B.n967 B.n966 585
R1019 B.n968 B.n967 585
R1020 B.n2 B.n0 585
R1021 B.n4 B.n2 585
R1022 B.n3 B.n1 585
R1023 B.n1509 B.n3 585
R1024 B.n1507 B.n1506 585
R1025 B.n1508 B.n1507 585
R1026 B.n1505 B.n9 585
R1027 B.n9 B.n8 585
R1028 B.n1504 B.n1503 585
R1029 B.n1503 B.n1502 585
R1030 B.n11 B.n10 585
R1031 B.n1501 B.n11 585
R1032 B.n1499 B.n1498 585
R1033 B.n1500 B.n1499 585
R1034 B.n1497 B.n16 585
R1035 B.n16 B.n15 585
R1036 B.n1496 B.n1495 585
R1037 B.n1495 B.n1494 585
R1038 B.n18 B.n17 585
R1039 B.n1493 B.n18 585
R1040 B.n1491 B.n1490 585
R1041 B.n1492 B.n1491 585
R1042 B.n1489 B.n23 585
R1043 B.n23 B.n22 585
R1044 B.n1488 B.n1487 585
R1045 B.n1487 B.n1486 585
R1046 B.n25 B.n24 585
R1047 B.n1485 B.n25 585
R1048 B.n1483 B.n1482 585
R1049 B.n1484 B.n1483 585
R1050 B.n1481 B.n30 585
R1051 B.n30 B.n29 585
R1052 B.n1480 B.n1479 585
R1053 B.n1479 B.n1478 585
R1054 B.n32 B.n31 585
R1055 B.n1477 B.n32 585
R1056 B.n1475 B.n1474 585
R1057 B.n1476 B.n1475 585
R1058 B.n1473 B.n37 585
R1059 B.n37 B.n36 585
R1060 B.n1472 B.n1471 585
R1061 B.n1471 B.n1470 585
R1062 B.n39 B.n38 585
R1063 B.n1469 B.n39 585
R1064 B.n1467 B.n1466 585
R1065 B.n1468 B.n1467 585
R1066 B.n1465 B.n44 585
R1067 B.n44 B.n43 585
R1068 B.n1464 B.n1463 585
R1069 B.n1463 B.n1462 585
R1070 B.n46 B.n45 585
R1071 B.n1461 B.n46 585
R1072 B.n1459 B.n1458 585
R1073 B.n1460 B.n1459 585
R1074 B.n1457 B.n51 585
R1075 B.n51 B.n50 585
R1076 B.n1456 B.n1455 585
R1077 B.n1455 B.n1454 585
R1078 B.n53 B.n52 585
R1079 B.n1453 B.n53 585
R1080 B.n1451 B.n1450 585
R1081 B.n1452 B.n1451 585
R1082 B.n1449 B.n58 585
R1083 B.n58 B.n57 585
R1084 B.n1448 B.n1447 585
R1085 B.n1447 B.n1446 585
R1086 B.n60 B.n59 585
R1087 B.n1445 B.n60 585
R1088 B.n1443 B.n1442 585
R1089 B.n1444 B.n1443 585
R1090 B.n1441 B.n65 585
R1091 B.n65 B.n64 585
R1092 B.n1440 B.n1439 585
R1093 B.n1439 B.n1438 585
R1094 B.n67 B.n66 585
R1095 B.n1437 B.n67 585
R1096 B.n1435 B.n1434 585
R1097 B.n1436 B.n1435 585
R1098 B.n1433 B.n72 585
R1099 B.n72 B.n71 585
R1100 B.n1432 B.n1431 585
R1101 B.n1431 B.n1430 585
R1102 B.n74 B.n73 585
R1103 B.n1429 B.n74 585
R1104 B.n1427 B.n1426 585
R1105 B.n1428 B.n1427 585
R1106 B.n1425 B.n79 585
R1107 B.n79 B.n78 585
R1108 B.n1424 B.n1423 585
R1109 B.n1423 B.n1422 585
R1110 B.n81 B.n80 585
R1111 B.n1421 B.n81 585
R1112 B.n1419 B.n1418 585
R1113 B.n1420 B.n1419 585
R1114 B.n1417 B.n86 585
R1115 B.n86 B.n85 585
R1116 B.n1416 B.n1415 585
R1117 B.n1415 B.n1414 585
R1118 B.n88 B.n87 585
R1119 B.n1413 B.n88 585
R1120 B.n1411 B.n1410 585
R1121 B.n1412 B.n1411 585
R1122 B.n1409 B.n93 585
R1123 B.n93 B.n92 585
R1124 B.n1408 B.n1407 585
R1125 B.n1407 B.n1406 585
R1126 B.n95 B.n94 585
R1127 B.n1405 B.n95 585
R1128 B.n1403 B.n1402 585
R1129 B.n1404 B.n1403 585
R1130 B.n1401 B.n100 585
R1131 B.n100 B.n99 585
R1132 B.n1400 B.n1399 585
R1133 B.n1399 B.n1398 585
R1134 B.n102 B.n101 585
R1135 B.n1397 B.n102 585
R1136 B.n1395 B.n1394 585
R1137 B.n1396 B.n1395 585
R1138 B.n1393 B.n107 585
R1139 B.n107 B.n106 585
R1140 B.n1392 B.n1391 585
R1141 B.n1391 B.n1390 585
R1142 B.n109 B.n108 585
R1143 B.n1389 B.n109 585
R1144 B.n1387 B.n1386 585
R1145 B.n1388 B.n1387 585
R1146 B.n1385 B.n114 585
R1147 B.n114 B.n113 585
R1148 B.n1384 B.n1383 585
R1149 B.n1383 B.n1382 585
R1150 B.n116 B.n115 585
R1151 B.n1381 B.n116 585
R1152 B.n1379 B.n1378 585
R1153 B.n1380 B.n1379 585
R1154 B.n1377 B.n121 585
R1155 B.n121 B.n120 585
R1156 B.n1376 B.n1375 585
R1157 B.n1375 B.n1374 585
R1158 B.n123 B.n122 585
R1159 B.n1373 B.n123 585
R1160 B.n1371 B.n1370 585
R1161 B.n1372 B.n1371 585
R1162 B.n1369 B.n128 585
R1163 B.n128 B.n127 585
R1164 B.n1368 B.n1367 585
R1165 B.n1367 B.n1366 585
R1166 B.n130 B.n129 585
R1167 B.n1365 B.n130 585
R1168 B.n1363 B.n1362 585
R1169 B.n1364 B.n1363 585
R1170 B.n1361 B.n135 585
R1171 B.n135 B.n134 585
R1172 B.n1360 B.n1359 585
R1173 B.n1359 B.n1358 585
R1174 B.n137 B.n136 585
R1175 B.n1357 B.n137 585
R1176 B.n1355 B.n1354 585
R1177 B.n1356 B.n1355 585
R1178 B.n1353 B.n142 585
R1179 B.n142 B.n141 585
R1180 B.n1352 B.n1351 585
R1181 B.n1351 B.n1350 585
R1182 B.n144 B.n143 585
R1183 B.n1349 B.n144 585
R1184 B.n1347 B.n1346 585
R1185 B.n1348 B.n1347 585
R1186 B.n1512 B.n1511 585
R1187 B.n1511 B.n1510 585
R1188 B.n726 B.n384 502.111
R1189 B.n1347 B.n149 502.111
R1190 B.n728 B.n382 502.111
R1191 B.n1076 B.n147 502.111
R1192 B.n423 B.t21 328.341
R1193 B.n417 B.t10 328.341
R1194 B.n182 B.t18 328.341
R1195 B.n189 B.t14 328.341
R1196 B.n1077 B.n148 256.663
R1197 B.n1083 B.n148 256.663
R1198 B.n1085 B.n148 256.663
R1199 B.n1091 B.n148 256.663
R1200 B.n1093 B.n148 256.663
R1201 B.n1099 B.n148 256.663
R1202 B.n1101 B.n148 256.663
R1203 B.n1107 B.n148 256.663
R1204 B.n1109 B.n148 256.663
R1205 B.n1115 B.n148 256.663
R1206 B.n1117 B.n148 256.663
R1207 B.n1123 B.n148 256.663
R1208 B.n1125 B.n148 256.663
R1209 B.n1131 B.n148 256.663
R1210 B.n1133 B.n148 256.663
R1211 B.n1139 B.n148 256.663
R1212 B.n1141 B.n148 256.663
R1213 B.n1147 B.n148 256.663
R1214 B.n1149 B.n148 256.663
R1215 B.n1155 B.n148 256.663
R1216 B.n1157 B.n148 256.663
R1217 B.n1163 B.n148 256.663
R1218 B.n1165 B.n148 256.663
R1219 B.n1171 B.n148 256.663
R1220 B.n1173 B.n148 256.663
R1221 B.n1179 B.n148 256.663
R1222 B.n1181 B.n148 256.663
R1223 B.n1187 B.n148 256.663
R1224 B.n1189 B.n148 256.663
R1225 B.n1195 B.n148 256.663
R1226 B.n1197 B.n148 256.663
R1227 B.n1204 B.n148 256.663
R1228 B.n1206 B.n148 256.663
R1229 B.n1212 B.n148 256.663
R1230 B.n1214 B.n148 256.663
R1231 B.n1220 B.n148 256.663
R1232 B.n1222 B.n148 256.663
R1233 B.n1228 B.n148 256.663
R1234 B.n1230 B.n148 256.663
R1235 B.n1236 B.n148 256.663
R1236 B.n1238 B.n148 256.663
R1237 B.n1244 B.n148 256.663
R1238 B.n1246 B.n148 256.663
R1239 B.n1252 B.n148 256.663
R1240 B.n1254 B.n148 256.663
R1241 B.n1260 B.n148 256.663
R1242 B.n1262 B.n148 256.663
R1243 B.n1268 B.n148 256.663
R1244 B.n1270 B.n148 256.663
R1245 B.n1276 B.n148 256.663
R1246 B.n1278 B.n148 256.663
R1247 B.n1284 B.n148 256.663
R1248 B.n1286 B.n148 256.663
R1249 B.n1292 B.n148 256.663
R1250 B.n1294 B.n148 256.663
R1251 B.n1300 B.n148 256.663
R1252 B.n1302 B.n148 256.663
R1253 B.n1308 B.n148 256.663
R1254 B.n1310 B.n148 256.663
R1255 B.n1316 B.n148 256.663
R1256 B.n1318 B.n148 256.663
R1257 B.n1324 B.n148 256.663
R1258 B.n1326 B.n148 256.663
R1259 B.n1332 B.n148 256.663
R1260 B.n1334 B.n148 256.663
R1261 B.n1340 B.n148 256.663
R1262 B.n1342 B.n148 256.663
R1263 B.n721 B.n383 256.663
R1264 B.n386 B.n383 256.663
R1265 B.n714 B.n383 256.663
R1266 B.n708 B.n383 256.663
R1267 B.n706 B.n383 256.663
R1268 B.n700 B.n383 256.663
R1269 B.n698 B.n383 256.663
R1270 B.n692 B.n383 256.663
R1271 B.n690 B.n383 256.663
R1272 B.n684 B.n383 256.663
R1273 B.n682 B.n383 256.663
R1274 B.n676 B.n383 256.663
R1275 B.n674 B.n383 256.663
R1276 B.n668 B.n383 256.663
R1277 B.n666 B.n383 256.663
R1278 B.n660 B.n383 256.663
R1279 B.n658 B.n383 256.663
R1280 B.n652 B.n383 256.663
R1281 B.n650 B.n383 256.663
R1282 B.n644 B.n383 256.663
R1283 B.n642 B.n383 256.663
R1284 B.n636 B.n383 256.663
R1285 B.n634 B.n383 256.663
R1286 B.n628 B.n383 256.663
R1287 B.n626 B.n383 256.663
R1288 B.n620 B.n383 256.663
R1289 B.n618 B.n383 256.663
R1290 B.n612 B.n383 256.663
R1291 B.n610 B.n383 256.663
R1292 B.n604 B.n383 256.663
R1293 B.n602 B.n383 256.663
R1294 B.n595 B.n383 256.663
R1295 B.n593 B.n383 256.663
R1296 B.n587 B.n383 256.663
R1297 B.n585 B.n383 256.663
R1298 B.n578 B.n383 256.663
R1299 B.n576 B.n383 256.663
R1300 B.n570 B.n383 256.663
R1301 B.n568 B.n383 256.663
R1302 B.n562 B.n383 256.663
R1303 B.n560 B.n383 256.663
R1304 B.n554 B.n383 256.663
R1305 B.n552 B.n383 256.663
R1306 B.n546 B.n383 256.663
R1307 B.n544 B.n383 256.663
R1308 B.n538 B.n383 256.663
R1309 B.n536 B.n383 256.663
R1310 B.n530 B.n383 256.663
R1311 B.n528 B.n383 256.663
R1312 B.n522 B.n383 256.663
R1313 B.n520 B.n383 256.663
R1314 B.n514 B.n383 256.663
R1315 B.n512 B.n383 256.663
R1316 B.n506 B.n383 256.663
R1317 B.n504 B.n383 256.663
R1318 B.n498 B.n383 256.663
R1319 B.n496 B.n383 256.663
R1320 B.n490 B.n383 256.663
R1321 B.n488 B.n383 256.663
R1322 B.n482 B.n383 256.663
R1323 B.n480 B.n383 256.663
R1324 B.n474 B.n383 256.663
R1325 B.n472 B.n383 256.663
R1326 B.n466 B.n383 256.663
R1327 B.n464 B.n383 256.663
R1328 B.n458 B.n383 256.663
R1329 B.n456 B.n383 256.663
R1330 B.n726 B.n378 163.367
R1331 B.n734 B.n378 163.367
R1332 B.n734 B.n376 163.367
R1333 B.n738 B.n376 163.367
R1334 B.n738 B.n370 163.367
R1335 B.n746 B.n370 163.367
R1336 B.n746 B.n368 163.367
R1337 B.n750 B.n368 163.367
R1338 B.n750 B.n362 163.367
R1339 B.n758 B.n362 163.367
R1340 B.n758 B.n360 163.367
R1341 B.n762 B.n360 163.367
R1342 B.n762 B.n354 163.367
R1343 B.n770 B.n354 163.367
R1344 B.n770 B.n352 163.367
R1345 B.n774 B.n352 163.367
R1346 B.n774 B.n346 163.367
R1347 B.n782 B.n346 163.367
R1348 B.n782 B.n344 163.367
R1349 B.n786 B.n344 163.367
R1350 B.n786 B.n338 163.367
R1351 B.n794 B.n338 163.367
R1352 B.n794 B.n336 163.367
R1353 B.n798 B.n336 163.367
R1354 B.n798 B.n330 163.367
R1355 B.n806 B.n330 163.367
R1356 B.n806 B.n328 163.367
R1357 B.n810 B.n328 163.367
R1358 B.n810 B.n322 163.367
R1359 B.n818 B.n322 163.367
R1360 B.n818 B.n320 163.367
R1361 B.n822 B.n320 163.367
R1362 B.n822 B.n314 163.367
R1363 B.n830 B.n314 163.367
R1364 B.n830 B.n312 163.367
R1365 B.n834 B.n312 163.367
R1366 B.n834 B.n306 163.367
R1367 B.n842 B.n306 163.367
R1368 B.n842 B.n304 163.367
R1369 B.n846 B.n304 163.367
R1370 B.n846 B.n298 163.367
R1371 B.n854 B.n298 163.367
R1372 B.n854 B.n296 163.367
R1373 B.n858 B.n296 163.367
R1374 B.n858 B.n290 163.367
R1375 B.n866 B.n290 163.367
R1376 B.n866 B.n288 163.367
R1377 B.n870 B.n288 163.367
R1378 B.n870 B.n282 163.367
R1379 B.n878 B.n282 163.367
R1380 B.n878 B.n280 163.367
R1381 B.n882 B.n280 163.367
R1382 B.n882 B.n274 163.367
R1383 B.n890 B.n274 163.367
R1384 B.n890 B.n272 163.367
R1385 B.n894 B.n272 163.367
R1386 B.n894 B.n266 163.367
R1387 B.n902 B.n266 163.367
R1388 B.n902 B.n264 163.367
R1389 B.n906 B.n264 163.367
R1390 B.n906 B.n258 163.367
R1391 B.n914 B.n258 163.367
R1392 B.n914 B.n256 163.367
R1393 B.n918 B.n256 163.367
R1394 B.n918 B.n250 163.367
R1395 B.n926 B.n250 163.367
R1396 B.n926 B.n248 163.367
R1397 B.n930 B.n248 163.367
R1398 B.n930 B.n242 163.367
R1399 B.n938 B.n242 163.367
R1400 B.n938 B.n240 163.367
R1401 B.n942 B.n240 163.367
R1402 B.n942 B.n234 163.367
R1403 B.n950 B.n234 163.367
R1404 B.n950 B.n232 163.367
R1405 B.n954 B.n232 163.367
R1406 B.n954 B.n226 163.367
R1407 B.n963 B.n226 163.367
R1408 B.n963 B.n224 163.367
R1409 B.n967 B.n224 163.367
R1410 B.n967 B.n2 163.367
R1411 B.n1511 B.n2 163.367
R1412 B.n1511 B.n3 163.367
R1413 B.n1507 B.n3 163.367
R1414 B.n1507 B.n9 163.367
R1415 B.n1503 B.n9 163.367
R1416 B.n1503 B.n11 163.367
R1417 B.n1499 B.n11 163.367
R1418 B.n1499 B.n16 163.367
R1419 B.n1495 B.n16 163.367
R1420 B.n1495 B.n18 163.367
R1421 B.n1491 B.n18 163.367
R1422 B.n1491 B.n23 163.367
R1423 B.n1487 B.n23 163.367
R1424 B.n1487 B.n25 163.367
R1425 B.n1483 B.n25 163.367
R1426 B.n1483 B.n30 163.367
R1427 B.n1479 B.n30 163.367
R1428 B.n1479 B.n32 163.367
R1429 B.n1475 B.n32 163.367
R1430 B.n1475 B.n37 163.367
R1431 B.n1471 B.n37 163.367
R1432 B.n1471 B.n39 163.367
R1433 B.n1467 B.n39 163.367
R1434 B.n1467 B.n44 163.367
R1435 B.n1463 B.n44 163.367
R1436 B.n1463 B.n46 163.367
R1437 B.n1459 B.n46 163.367
R1438 B.n1459 B.n51 163.367
R1439 B.n1455 B.n51 163.367
R1440 B.n1455 B.n53 163.367
R1441 B.n1451 B.n53 163.367
R1442 B.n1451 B.n58 163.367
R1443 B.n1447 B.n58 163.367
R1444 B.n1447 B.n60 163.367
R1445 B.n1443 B.n60 163.367
R1446 B.n1443 B.n65 163.367
R1447 B.n1439 B.n65 163.367
R1448 B.n1439 B.n67 163.367
R1449 B.n1435 B.n67 163.367
R1450 B.n1435 B.n72 163.367
R1451 B.n1431 B.n72 163.367
R1452 B.n1431 B.n74 163.367
R1453 B.n1427 B.n74 163.367
R1454 B.n1427 B.n79 163.367
R1455 B.n1423 B.n79 163.367
R1456 B.n1423 B.n81 163.367
R1457 B.n1419 B.n81 163.367
R1458 B.n1419 B.n86 163.367
R1459 B.n1415 B.n86 163.367
R1460 B.n1415 B.n88 163.367
R1461 B.n1411 B.n88 163.367
R1462 B.n1411 B.n93 163.367
R1463 B.n1407 B.n93 163.367
R1464 B.n1407 B.n95 163.367
R1465 B.n1403 B.n95 163.367
R1466 B.n1403 B.n100 163.367
R1467 B.n1399 B.n100 163.367
R1468 B.n1399 B.n102 163.367
R1469 B.n1395 B.n102 163.367
R1470 B.n1395 B.n107 163.367
R1471 B.n1391 B.n107 163.367
R1472 B.n1391 B.n109 163.367
R1473 B.n1387 B.n109 163.367
R1474 B.n1387 B.n114 163.367
R1475 B.n1383 B.n114 163.367
R1476 B.n1383 B.n116 163.367
R1477 B.n1379 B.n116 163.367
R1478 B.n1379 B.n121 163.367
R1479 B.n1375 B.n121 163.367
R1480 B.n1375 B.n123 163.367
R1481 B.n1371 B.n123 163.367
R1482 B.n1371 B.n128 163.367
R1483 B.n1367 B.n128 163.367
R1484 B.n1367 B.n130 163.367
R1485 B.n1363 B.n130 163.367
R1486 B.n1363 B.n135 163.367
R1487 B.n1359 B.n135 163.367
R1488 B.n1359 B.n137 163.367
R1489 B.n1355 B.n137 163.367
R1490 B.n1355 B.n142 163.367
R1491 B.n1351 B.n142 163.367
R1492 B.n1351 B.n144 163.367
R1493 B.n1347 B.n144 163.367
R1494 B.n722 B.n720 163.367
R1495 B.n720 B.n719 163.367
R1496 B.n716 B.n715 163.367
R1497 B.n713 B.n388 163.367
R1498 B.n709 B.n707 163.367
R1499 B.n705 B.n390 163.367
R1500 B.n701 B.n699 163.367
R1501 B.n697 B.n392 163.367
R1502 B.n693 B.n691 163.367
R1503 B.n689 B.n394 163.367
R1504 B.n685 B.n683 163.367
R1505 B.n681 B.n396 163.367
R1506 B.n677 B.n675 163.367
R1507 B.n673 B.n398 163.367
R1508 B.n669 B.n667 163.367
R1509 B.n665 B.n400 163.367
R1510 B.n661 B.n659 163.367
R1511 B.n657 B.n402 163.367
R1512 B.n653 B.n651 163.367
R1513 B.n649 B.n404 163.367
R1514 B.n645 B.n643 163.367
R1515 B.n641 B.n406 163.367
R1516 B.n637 B.n635 163.367
R1517 B.n633 B.n408 163.367
R1518 B.n629 B.n627 163.367
R1519 B.n625 B.n410 163.367
R1520 B.n621 B.n619 163.367
R1521 B.n617 B.n412 163.367
R1522 B.n613 B.n611 163.367
R1523 B.n609 B.n414 163.367
R1524 B.n605 B.n603 163.367
R1525 B.n601 B.n416 163.367
R1526 B.n596 B.n594 163.367
R1527 B.n592 B.n420 163.367
R1528 B.n588 B.n586 163.367
R1529 B.n584 B.n422 163.367
R1530 B.n579 B.n577 163.367
R1531 B.n575 B.n426 163.367
R1532 B.n571 B.n569 163.367
R1533 B.n567 B.n428 163.367
R1534 B.n563 B.n561 163.367
R1535 B.n559 B.n430 163.367
R1536 B.n555 B.n553 163.367
R1537 B.n551 B.n432 163.367
R1538 B.n547 B.n545 163.367
R1539 B.n543 B.n434 163.367
R1540 B.n539 B.n537 163.367
R1541 B.n535 B.n436 163.367
R1542 B.n531 B.n529 163.367
R1543 B.n527 B.n438 163.367
R1544 B.n523 B.n521 163.367
R1545 B.n519 B.n440 163.367
R1546 B.n515 B.n513 163.367
R1547 B.n511 B.n442 163.367
R1548 B.n507 B.n505 163.367
R1549 B.n503 B.n444 163.367
R1550 B.n499 B.n497 163.367
R1551 B.n495 B.n446 163.367
R1552 B.n491 B.n489 163.367
R1553 B.n487 B.n448 163.367
R1554 B.n483 B.n481 163.367
R1555 B.n479 B.n450 163.367
R1556 B.n475 B.n473 163.367
R1557 B.n471 B.n452 163.367
R1558 B.n467 B.n465 163.367
R1559 B.n463 B.n454 163.367
R1560 B.n459 B.n457 163.367
R1561 B.n728 B.n380 163.367
R1562 B.n732 B.n380 163.367
R1563 B.n732 B.n374 163.367
R1564 B.n740 B.n374 163.367
R1565 B.n740 B.n372 163.367
R1566 B.n744 B.n372 163.367
R1567 B.n744 B.n365 163.367
R1568 B.n752 B.n365 163.367
R1569 B.n752 B.n363 163.367
R1570 B.n756 B.n363 163.367
R1571 B.n756 B.n358 163.367
R1572 B.n764 B.n358 163.367
R1573 B.n764 B.n356 163.367
R1574 B.n768 B.n356 163.367
R1575 B.n768 B.n350 163.367
R1576 B.n776 B.n350 163.367
R1577 B.n776 B.n348 163.367
R1578 B.n780 B.n348 163.367
R1579 B.n780 B.n342 163.367
R1580 B.n788 B.n342 163.367
R1581 B.n788 B.n340 163.367
R1582 B.n792 B.n340 163.367
R1583 B.n792 B.n334 163.367
R1584 B.n800 B.n334 163.367
R1585 B.n800 B.n332 163.367
R1586 B.n804 B.n332 163.367
R1587 B.n804 B.n326 163.367
R1588 B.n812 B.n326 163.367
R1589 B.n812 B.n324 163.367
R1590 B.n816 B.n324 163.367
R1591 B.n816 B.n318 163.367
R1592 B.n824 B.n318 163.367
R1593 B.n824 B.n316 163.367
R1594 B.n828 B.n316 163.367
R1595 B.n828 B.n309 163.367
R1596 B.n836 B.n309 163.367
R1597 B.n836 B.n307 163.367
R1598 B.n840 B.n307 163.367
R1599 B.n840 B.n302 163.367
R1600 B.n848 B.n302 163.367
R1601 B.n848 B.n300 163.367
R1602 B.n852 B.n300 163.367
R1603 B.n852 B.n294 163.367
R1604 B.n860 B.n294 163.367
R1605 B.n860 B.n292 163.367
R1606 B.n864 B.n292 163.367
R1607 B.n864 B.n285 163.367
R1608 B.n872 B.n285 163.367
R1609 B.n872 B.n283 163.367
R1610 B.n876 B.n283 163.367
R1611 B.n876 B.n278 163.367
R1612 B.n884 B.n278 163.367
R1613 B.n884 B.n276 163.367
R1614 B.n888 B.n276 163.367
R1615 B.n888 B.n270 163.367
R1616 B.n896 B.n270 163.367
R1617 B.n896 B.n268 163.367
R1618 B.n900 B.n268 163.367
R1619 B.n900 B.n261 163.367
R1620 B.n908 B.n261 163.367
R1621 B.n908 B.n259 163.367
R1622 B.n912 B.n259 163.367
R1623 B.n912 B.n254 163.367
R1624 B.n920 B.n254 163.367
R1625 B.n920 B.n252 163.367
R1626 B.n924 B.n252 163.367
R1627 B.n924 B.n246 163.367
R1628 B.n932 B.n246 163.367
R1629 B.n932 B.n244 163.367
R1630 B.n936 B.n244 163.367
R1631 B.n936 B.n238 163.367
R1632 B.n944 B.n238 163.367
R1633 B.n944 B.n236 163.367
R1634 B.n948 B.n236 163.367
R1635 B.n948 B.n230 163.367
R1636 B.n956 B.n230 163.367
R1637 B.n956 B.n228 163.367
R1638 B.n961 B.n228 163.367
R1639 B.n961 B.n222 163.367
R1640 B.n969 B.n222 163.367
R1641 B.n970 B.n969 163.367
R1642 B.n970 B.n5 163.367
R1643 B.n6 B.n5 163.367
R1644 B.n7 B.n6 163.367
R1645 B.n975 B.n7 163.367
R1646 B.n975 B.n12 163.367
R1647 B.n13 B.n12 163.367
R1648 B.n14 B.n13 163.367
R1649 B.n980 B.n14 163.367
R1650 B.n980 B.n19 163.367
R1651 B.n20 B.n19 163.367
R1652 B.n21 B.n20 163.367
R1653 B.n985 B.n21 163.367
R1654 B.n985 B.n26 163.367
R1655 B.n27 B.n26 163.367
R1656 B.n28 B.n27 163.367
R1657 B.n990 B.n28 163.367
R1658 B.n990 B.n33 163.367
R1659 B.n34 B.n33 163.367
R1660 B.n35 B.n34 163.367
R1661 B.n995 B.n35 163.367
R1662 B.n995 B.n40 163.367
R1663 B.n41 B.n40 163.367
R1664 B.n42 B.n41 163.367
R1665 B.n1000 B.n42 163.367
R1666 B.n1000 B.n47 163.367
R1667 B.n48 B.n47 163.367
R1668 B.n49 B.n48 163.367
R1669 B.n1005 B.n49 163.367
R1670 B.n1005 B.n54 163.367
R1671 B.n55 B.n54 163.367
R1672 B.n56 B.n55 163.367
R1673 B.n1010 B.n56 163.367
R1674 B.n1010 B.n61 163.367
R1675 B.n62 B.n61 163.367
R1676 B.n63 B.n62 163.367
R1677 B.n1015 B.n63 163.367
R1678 B.n1015 B.n68 163.367
R1679 B.n69 B.n68 163.367
R1680 B.n70 B.n69 163.367
R1681 B.n1020 B.n70 163.367
R1682 B.n1020 B.n75 163.367
R1683 B.n76 B.n75 163.367
R1684 B.n77 B.n76 163.367
R1685 B.n1025 B.n77 163.367
R1686 B.n1025 B.n82 163.367
R1687 B.n83 B.n82 163.367
R1688 B.n84 B.n83 163.367
R1689 B.n1030 B.n84 163.367
R1690 B.n1030 B.n89 163.367
R1691 B.n90 B.n89 163.367
R1692 B.n91 B.n90 163.367
R1693 B.n1035 B.n91 163.367
R1694 B.n1035 B.n96 163.367
R1695 B.n97 B.n96 163.367
R1696 B.n98 B.n97 163.367
R1697 B.n1040 B.n98 163.367
R1698 B.n1040 B.n103 163.367
R1699 B.n104 B.n103 163.367
R1700 B.n105 B.n104 163.367
R1701 B.n1045 B.n105 163.367
R1702 B.n1045 B.n110 163.367
R1703 B.n111 B.n110 163.367
R1704 B.n112 B.n111 163.367
R1705 B.n1050 B.n112 163.367
R1706 B.n1050 B.n117 163.367
R1707 B.n118 B.n117 163.367
R1708 B.n119 B.n118 163.367
R1709 B.n1055 B.n119 163.367
R1710 B.n1055 B.n124 163.367
R1711 B.n125 B.n124 163.367
R1712 B.n126 B.n125 163.367
R1713 B.n1060 B.n126 163.367
R1714 B.n1060 B.n131 163.367
R1715 B.n132 B.n131 163.367
R1716 B.n133 B.n132 163.367
R1717 B.n1065 B.n133 163.367
R1718 B.n1065 B.n138 163.367
R1719 B.n139 B.n138 163.367
R1720 B.n140 B.n139 163.367
R1721 B.n1070 B.n140 163.367
R1722 B.n1070 B.n145 163.367
R1723 B.n146 B.n145 163.367
R1724 B.n147 B.n146 163.367
R1725 B.n1343 B.n1341 163.367
R1726 B.n1339 B.n151 163.367
R1727 B.n1335 B.n1333 163.367
R1728 B.n1331 B.n153 163.367
R1729 B.n1327 B.n1325 163.367
R1730 B.n1323 B.n155 163.367
R1731 B.n1319 B.n1317 163.367
R1732 B.n1315 B.n157 163.367
R1733 B.n1311 B.n1309 163.367
R1734 B.n1307 B.n159 163.367
R1735 B.n1303 B.n1301 163.367
R1736 B.n1299 B.n161 163.367
R1737 B.n1295 B.n1293 163.367
R1738 B.n1291 B.n163 163.367
R1739 B.n1287 B.n1285 163.367
R1740 B.n1283 B.n165 163.367
R1741 B.n1279 B.n1277 163.367
R1742 B.n1275 B.n167 163.367
R1743 B.n1271 B.n1269 163.367
R1744 B.n1267 B.n169 163.367
R1745 B.n1263 B.n1261 163.367
R1746 B.n1259 B.n171 163.367
R1747 B.n1255 B.n1253 163.367
R1748 B.n1251 B.n173 163.367
R1749 B.n1247 B.n1245 163.367
R1750 B.n1243 B.n175 163.367
R1751 B.n1239 B.n1237 163.367
R1752 B.n1235 B.n177 163.367
R1753 B.n1231 B.n1229 163.367
R1754 B.n1227 B.n179 163.367
R1755 B.n1223 B.n1221 163.367
R1756 B.n1219 B.n181 163.367
R1757 B.n1215 B.n1213 163.367
R1758 B.n1211 B.n186 163.367
R1759 B.n1207 B.n1205 163.367
R1760 B.n1203 B.n188 163.367
R1761 B.n1198 B.n1196 163.367
R1762 B.n1194 B.n192 163.367
R1763 B.n1190 B.n1188 163.367
R1764 B.n1186 B.n194 163.367
R1765 B.n1182 B.n1180 163.367
R1766 B.n1178 B.n196 163.367
R1767 B.n1174 B.n1172 163.367
R1768 B.n1170 B.n198 163.367
R1769 B.n1166 B.n1164 163.367
R1770 B.n1162 B.n200 163.367
R1771 B.n1158 B.n1156 163.367
R1772 B.n1154 B.n202 163.367
R1773 B.n1150 B.n1148 163.367
R1774 B.n1146 B.n204 163.367
R1775 B.n1142 B.n1140 163.367
R1776 B.n1138 B.n206 163.367
R1777 B.n1134 B.n1132 163.367
R1778 B.n1130 B.n208 163.367
R1779 B.n1126 B.n1124 163.367
R1780 B.n1122 B.n210 163.367
R1781 B.n1118 B.n1116 163.367
R1782 B.n1114 B.n212 163.367
R1783 B.n1110 B.n1108 163.367
R1784 B.n1106 B.n214 163.367
R1785 B.n1102 B.n1100 163.367
R1786 B.n1098 B.n216 163.367
R1787 B.n1094 B.n1092 163.367
R1788 B.n1090 B.n218 163.367
R1789 B.n1086 B.n1084 163.367
R1790 B.n1082 B.n220 163.367
R1791 B.n1078 B.n1076 163.367
R1792 B.n423 B.t23 149.805
R1793 B.n189 B.t16 149.805
R1794 B.n417 B.t13 149.78
R1795 B.n182 B.t19 149.78
R1796 B.n424 B.n423 81.455
R1797 B.n418 B.n417 81.455
R1798 B.n183 B.n182 81.455
R1799 B.n190 B.n189 81.455
R1800 B.n721 B.n384 71.676
R1801 B.n719 B.n386 71.676
R1802 B.n715 B.n714 71.676
R1803 B.n708 B.n388 71.676
R1804 B.n707 B.n706 71.676
R1805 B.n700 B.n390 71.676
R1806 B.n699 B.n698 71.676
R1807 B.n692 B.n392 71.676
R1808 B.n691 B.n690 71.676
R1809 B.n684 B.n394 71.676
R1810 B.n683 B.n682 71.676
R1811 B.n676 B.n396 71.676
R1812 B.n675 B.n674 71.676
R1813 B.n668 B.n398 71.676
R1814 B.n667 B.n666 71.676
R1815 B.n660 B.n400 71.676
R1816 B.n659 B.n658 71.676
R1817 B.n652 B.n402 71.676
R1818 B.n651 B.n650 71.676
R1819 B.n644 B.n404 71.676
R1820 B.n643 B.n642 71.676
R1821 B.n636 B.n406 71.676
R1822 B.n635 B.n634 71.676
R1823 B.n628 B.n408 71.676
R1824 B.n627 B.n626 71.676
R1825 B.n620 B.n410 71.676
R1826 B.n619 B.n618 71.676
R1827 B.n612 B.n412 71.676
R1828 B.n611 B.n610 71.676
R1829 B.n604 B.n414 71.676
R1830 B.n603 B.n602 71.676
R1831 B.n595 B.n416 71.676
R1832 B.n594 B.n593 71.676
R1833 B.n587 B.n420 71.676
R1834 B.n586 B.n585 71.676
R1835 B.n578 B.n422 71.676
R1836 B.n577 B.n576 71.676
R1837 B.n570 B.n426 71.676
R1838 B.n569 B.n568 71.676
R1839 B.n562 B.n428 71.676
R1840 B.n561 B.n560 71.676
R1841 B.n554 B.n430 71.676
R1842 B.n553 B.n552 71.676
R1843 B.n546 B.n432 71.676
R1844 B.n545 B.n544 71.676
R1845 B.n538 B.n434 71.676
R1846 B.n537 B.n536 71.676
R1847 B.n530 B.n436 71.676
R1848 B.n529 B.n528 71.676
R1849 B.n522 B.n438 71.676
R1850 B.n521 B.n520 71.676
R1851 B.n514 B.n440 71.676
R1852 B.n513 B.n512 71.676
R1853 B.n506 B.n442 71.676
R1854 B.n505 B.n504 71.676
R1855 B.n498 B.n444 71.676
R1856 B.n497 B.n496 71.676
R1857 B.n490 B.n446 71.676
R1858 B.n489 B.n488 71.676
R1859 B.n482 B.n448 71.676
R1860 B.n481 B.n480 71.676
R1861 B.n474 B.n450 71.676
R1862 B.n473 B.n472 71.676
R1863 B.n466 B.n452 71.676
R1864 B.n465 B.n464 71.676
R1865 B.n458 B.n454 71.676
R1866 B.n457 B.n456 71.676
R1867 B.n1342 B.n149 71.676
R1868 B.n1341 B.n1340 71.676
R1869 B.n1334 B.n151 71.676
R1870 B.n1333 B.n1332 71.676
R1871 B.n1326 B.n153 71.676
R1872 B.n1325 B.n1324 71.676
R1873 B.n1318 B.n155 71.676
R1874 B.n1317 B.n1316 71.676
R1875 B.n1310 B.n157 71.676
R1876 B.n1309 B.n1308 71.676
R1877 B.n1302 B.n159 71.676
R1878 B.n1301 B.n1300 71.676
R1879 B.n1294 B.n161 71.676
R1880 B.n1293 B.n1292 71.676
R1881 B.n1286 B.n163 71.676
R1882 B.n1285 B.n1284 71.676
R1883 B.n1278 B.n165 71.676
R1884 B.n1277 B.n1276 71.676
R1885 B.n1270 B.n167 71.676
R1886 B.n1269 B.n1268 71.676
R1887 B.n1262 B.n169 71.676
R1888 B.n1261 B.n1260 71.676
R1889 B.n1254 B.n171 71.676
R1890 B.n1253 B.n1252 71.676
R1891 B.n1246 B.n173 71.676
R1892 B.n1245 B.n1244 71.676
R1893 B.n1238 B.n175 71.676
R1894 B.n1237 B.n1236 71.676
R1895 B.n1230 B.n177 71.676
R1896 B.n1229 B.n1228 71.676
R1897 B.n1222 B.n179 71.676
R1898 B.n1221 B.n1220 71.676
R1899 B.n1214 B.n181 71.676
R1900 B.n1213 B.n1212 71.676
R1901 B.n1206 B.n186 71.676
R1902 B.n1205 B.n1204 71.676
R1903 B.n1197 B.n188 71.676
R1904 B.n1196 B.n1195 71.676
R1905 B.n1189 B.n192 71.676
R1906 B.n1188 B.n1187 71.676
R1907 B.n1181 B.n194 71.676
R1908 B.n1180 B.n1179 71.676
R1909 B.n1173 B.n196 71.676
R1910 B.n1172 B.n1171 71.676
R1911 B.n1165 B.n198 71.676
R1912 B.n1164 B.n1163 71.676
R1913 B.n1157 B.n200 71.676
R1914 B.n1156 B.n1155 71.676
R1915 B.n1149 B.n202 71.676
R1916 B.n1148 B.n1147 71.676
R1917 B.n1141 B.n204 71.676
R1918 B.n1140 B.n1139 71.676
R1919 B.n1133 B.n206 71.676
R1920 B.n1132 B.n1131 71.676
R1921 B.n1125 B.n208 71.676
R1922 B.n1124 B.n1123 71.676
R1923 B.n1117 B.n210 71.676
R1924 B.n1116 B.n1115 71.676
R1925 B.n1109 B.n212 71.676
R1926 B.n1108 B.n1107 71.676
R1927 B.n1101 B.n214 71.676
R1928 B.n1100 B.n1099 71.676
R1929 B.n1093 B.n216 71.676
R1930 B.n1092 B.n1091 71.676
R1931 B.n1085 B.n218 71.676
R1932 B.n1084 B.n1083 71.676
R1933 B.n1077 B.n220 71.676
R1934 B.n1078 B.n1077 71.676
R1935 B.n1083 B.n1082 71.676
R1936 B.n1086 B.n1085 71.676
R1937 B.n1091 B.n1090 71.676
R1938 B.n1094 B.n1093 71.676
R1939 B.n1099 B.n1098 71.676
R1940 B.n1102 B.n1101 71.676
R1941 B.n1107 B.n1106 71.676
R1942 B.n1110 B.n1109 71.676
R1943 B.n1115 B.n1114 71.676
R1944 B.n1118 B.n1117 71.676
R1945 B.n1123 B.n1122 71.676
R1946 B.n1126 B.n1125 71.676
R1947 B.n1131 B.n1130 71.676
R1948 B.n1134 B.n1133 71.676
R1949 B.n1139 B.n1138 71.676
R1950 B.n1142 B.n1141 71.676
R1951 B.n1147 B.n1146 71.676
R1952 B.n1150 B.n1149 71.676
R1953 B.n1155 B.n1154 71.676
R1954 B.n1158 B.n1157 71.676
R1955 B.n1163 B.n1162 71.676
R1956 B.n1166 B.n1165 71.676
R1957 B.n1171 B.n1170 71.676
R1958 B.n1174 B.n1173 71.676
R1959 B.n1179 B.n1178 71.676
R1960 B.n1182 B.n1181 71.676
R1961 B.n1187 B.n1186 71.676
R1962 B.n1190 B.n1189 71.676
R1963 B.n1195 B.n1194 71.676
R1964 B.n1198 B.n1197 71.676
R1965 B.n1204 B.n1203 71.676
R1966 B.n1207 B.n1206 71.676
R1967 B.n1212 B.n1211 71.676
R1968 B.n1215 B.n1214 71.676
R1969 B.n1220 B.n1219 71.676
R1970 B.n1223 B.n1222 71.676
R1971 B.n1228 B.n1227 71.676
R1972 B.n1231 B.n1230 71.676
R1973 B.n1236 B.n1235 71.676
R1974 B.n1239 B.n1238 71.676
R1975 B.n1244 B.n1243 71.676
R1976 B.n1247 B.n1246 71.676
R1977 B.n1252 B.n1251 71.676
R1978 B.n1255 B.n1254 71.676
R1979 B.n1260 B.n1259 71.676
R1980 B.n1263 B.n1262 71.676
R1981 B.n1268 B.n1267 71.676
R1982 B.n1271 B.n1270 71.676
R1983 B.n1276 B.n1275 71.676
R1984 B.n1279 B.n1278 71.676
R1985 B.n1284 B.n1283 71.676
R1986 B.n1287 B.n1286 71.676
R1987 B.n1292 B.n1291 71.676
R1988 B.n1295 B.n1294 71.676
R1989 B.n1300 B.n1299 71.676
R1990 B.n1303 B.n1302 71.676
R1991 B.n1308 B.n1307 71.676
R1992 B.n1311 B.n1310 71.676
R1993 B.n1316 B.n1315 71.676
R1994 B.n1319 B.n1318 71.676
R1995 B.n1324 B.n1323 71.676
R1996 B.n1327 B.n1326 71.676
R1997 B.n1332 B.n1331 71.676
R1998 B.n1335 B.n1334 71.676
R1999 B.n1340 B.n1339 71.676
R2000 B.n1343 B.n1342 71.676
R2001 B.n722 B.n721 71.676
R2002 B.n716 B.n386 71.676
R2003 B.n714 B.n713 71.676
R2004 B.n709 B.n708 71.676
R2005 B.n706 B.n705 71.676
R2006 B.n701 B.n700 71.676
R2007 B.n698 B.n697 71.676
R2008 B.n693 B.n692 71.676
R2009 B.n690 B.n689 71.676
R2010 B.n685 B.n684 71.676
R2011 B.n682 B.n681 71.676
R2012 B.n677 B.n676 71.676
R2013 B.n674 B.n673 71.676
R2014 B.n669 B.n668 71.676
R2015 B.n666 B.n665 71.676
R2016 B.n661 B.n660 71.676
R2017 B.n658 B.n657 71.676
R2018 B.n653 B.n652 71.676
R2019 B.n650 B.n649 71.676
R2020 B.n645 B.n644 71.676
R2021 B.n642 B.n641 71.676
R2022 B.n637 B.n636 71.676
R2023 B.n634 B.n633 71.676
R2024 B.n629 B.n628 71.676
R2025 B.n626 B.n625 71.676
R2026 B.n621 B.n620 71.676
R2027 B.n618 B.n617 71.676
R2028 B.n613 B.n612 71.676
R2029 B.n610 B.n609 71.676
R2030 B.n605 B.n604 71.676
R2031 B.n602 B.n601 71.676
R2032 B.n596 B.n595 71.676
R2033 B.n593 B.n592 71.676
R2034 B.n588 B.n587 71.676
R2035 B.n585 B.n584 71.676
R2036 B.n579 B.n578 71.676
R2037 B.n576 B.n575 71.676
R2038 B.n571 B.n570 71.676
R2039 B.n568 B.n567 71.676
R2040 B.n563 B.n562 71.676
R2041 B.n560 B.n559 71.676
R2042 B.n555 B.n554 71.676
R2043 B.n552 B.n551 71.676
R2044 B.n547 B.n546 71.676
R2045 B.n544 B.n543 71.676
R2046 B.n539 B.n538 71.676
R2047 B.n536 B.n535 71.676
R2048 B.n531 B.n530 71.676
R2049 B.n528 B.n527 71.676
R2050 B.n523 B.n522 71.676
R2051 B.n520 B.n519 71.676
R2052 B.n515 B.n514 71.676
R2053 B.n512 B.n511 71.676
R2054 B.n507 B.n506 71.676
R2055 B.n504 B.n503 71.676
R2056 B.n499 B.n498 71.676
R2057 B.n496 B.n495 71.676
R2058 B.n491 B.n490 71.676
R2059 B.n488 B.n487 71.676
R2060 B.n483 B.n482 71.676
R2061 B.n480 B.n479 71.676
R2062 B.n475 B.n474 71.676
R2063 B.n472 B.n471 71.676
R2064 B.n467 B.n466 71.676
R2065 B.n464 B.n463 71.676
R2066 B.n459 B.n458 71.676
R2067 B.n456 B.n382 71.676
R2068 B.n424 B.t22 68.3507
R2069 B.n190 B.t17 68.3507
R2070 B.n418 B.t12 68.3249
R2071 B.n183 B.t20 68.3249
R2072 B.n727 B.n383 62.7287
R2073 B.n1348 B.n148 62.7287
R2074 B.n581 B.n424 59.5399
R2075 B.n599 B.n418 59.5399
R2076 B.n184 B.n183 59.5399
R2077 B.n1201 B.n190 59.5399
R2078 B.n1346 B.n1345 32.6249
R2079 B.n1075 B.n1074 32.6249
R2080 B.n729 B.n381 32.6249
R2081 B.n725 B.n724 32.6249
R2082 B.n727 B.n379 30.6877
R2083 B.n733 B.n379 30.6877
R2084 B.n733 B.n375 30.6877
R2085 B.n739 B.n375 30.6877
R2086 B.n739 B.n371 30.6877
R2087 B.n745 B.n371 30.6877
R2088 B.n745 B.n366 30.6877
R2089 B.n751 B.n366 30.6877
R2090 B.n751 B.n367 30.6877
R2091 B.n757 B.n359 30.6877
R2092 B.n763 B.n359 30.6877
R2093 B.n763 B.n355 30.6877
R2094 B.n769 B.n355 30.6877
R2095 B.n769 B.n351 30.6877
R2096 B.n775 B.n351 30.6877
R2097 B.n775 B.n347 30.6877
R2098 B.n781 B.n347 30.6877
R2099 B.n781 B.n343 30.6877
R2100 B.n787 B.n343 30.6877
R2101 B.n787 B.n339 30.6877
R2102 B.n793 B.n339 30.6877
R2103 B.n793 B.n335 30.6877
R2104 B.n799 B.n335 30.6877
R2105 B.n805 B.n331 30.6877
R2106 B.n805 B.n327 30.6877
R2107 B.n811 B.n327 30.6877
R2108 B.n811 B.n323 30.6877
R2109 B.n817 B.n323 30.6877
R2110 B.n817 B.n319 30.6877
R2111 B.n823 B.n319 30.6877
R2112 B.n823 B.n315 30.6877
R2113 B.n829 B.n315 30.6877
R2114 B.n829 B.n310 30.6877
R2115 B.n835 B.n310 30.6877
R2116 B.n835 B.n311 30.6877
R2117 B.n841 B.n303 30.6877
R2118 B.n847 B.n303 30.6877
R2119 B.n847 B.n299 30.6877
R2120 B.n853 B.n299 30.6877
R2121 B.n853 B.n295 30.6877
R2122 B.n859 B.n295 30.6877
R2123 B.n859 B.n291 30.6877
R2124 B.n865 B.n291 30.6877
R2125 B.n865 B.n286 30.6877
R2126 B.n871 B.n286 30.6877
R2127 B.n871 B.n287 30.6877
R2128 B.n877 B.n279 30.6877
R2129 B.n883 B.n279 30.6877
R2130 B.n883 B.n275 30.6877
R2131 B.n889 B.n275 30.6877
R2132 B.n889 B.n271 30.6877
R2133 B.n895 B.n271 30.6877
R2134 B.n895 B.n267 30.6877
R2135 B.n901 B.n267 30.6877
R2136 B.n901 B.n262 30.6877
R2137 B.n907 B.n262 30.6877
R2138 B.n907 B.n263 30.6877
R2139 B.n913 B.n255 30.6877
R2140 B.n919 B.n255 30.6877
R2141 B.n919 B.n251 30.6877
R2142 B.n925 B.n251 30.6877
R2143 B.n925 B.n247 30.6877
R2144 B.n931 B.n247 30.6877
R2145 B.n931 B.n243 30.6877
R2146 B.n937 B.n243 30.6877
R2147 B.n937 B.n239 30.6877
R2148 B.n943 B.n239 30.6877
R2149 B.n943 B.n235 30.6877
R2150 B.n949 B.n235 30.6877
R2151 B.n955 B.n231 30.6877
R2152 B.n955 B.n227 30.6877
R2153 B.n962 B.n227 30.6877
R2154 B.n962 B.n223 30.6877
R2155 B.n968 B.n223 30.6877
R2156 B.n968 B.n4 30.6877
R2157 B.n1510 B.n4 30.6877
R2158 B.n1510 B.n1509 30.6877
R2159 B.n1509 B.n1508 30.6877
R2160 B.n1508 B.n8 30.6877
R2161 B.n1502 B.n8 30.6877
R2162 B.n1502 B.n1501 30.6877
R2163 B.n1501 B.n1500 30.6877
R2164 B.n1500 B.n15 30.6877
R2165 B.n1494 B.n1493 30.6877
R2166 B.n1493 B.n1492 30.6877
R2167 B.n1492 B.n22 30.6877
R2168 B.n1486 B.n22 30.6877
R2169 B.n1486 B.n1485 30.6877
R2170 B.n1485 B.n1484 30.6877
R2171 B.n1484 B.n29 30.6877
R2172 B.n1478 B.n29 30.6877
R2173 B.n1478 B.n1477 30.6877
R2174 B.n1477 B.n1476 30.6877
R2175 B.n1476 B.n36 30.6877
R2176 B.n1470 B.n36 30.6877
R2177 B.n1469 B.n1468 30.6877
R2178 B.n1468 B.n43 30.6877
R2179 B.n1462 B.n43 30.6877
R2180 B.n1462 B.n1461 30.6877
R2181 B.n1461 B.n1460 30.6877
R2182 B.n1460 B.n50 30.6877
R2183 B.n1454 B.n50 30.6877
R2184 B.n1454 B.n1453 30.6877
R2185 B.n1453 B.n1452 30.6877
R2186 B.n1452 B.n57 30.6877
R2187 B.n1446 B.n57 30.6877
R2188 B.n1445 B.n1444 30.6877
R2189 B.n1444 B.n64 30.6877
R2190 B.n1438 B.n64 30.6877
R2191 B.n1438 B.n1437 30.6877
R2192 B.n1437 B.n1436 30.6877
R2193 B.n1436 B.n71 30.6877
R2194 B.n1430 B.n71 30.6877
R2195 B.n1430 B.n1429 30.6877
R2196 B.n1429 B.n1428 30.6877
R2197 B.n1428 B.n78 30.6877
R2198 B.n1422 B.n78 30.6877
R2199 B.n1421 B.n1420 30.6877
R2200 B.n1420 B.n85 30.6877
R2201 B.n1414 B.n85 30.6877
R2202 B.n1414 B.n1413 30.6877
R2203 B.n1413 B.n1412 30.6877
R2204 B.n1412 B.n92 30.6877
R2205 B.n1406 B.n92 30.6877
R2206 B.n1406 B.n1405 30.6877
R2207 B.n1405 B.n1404 30.6877
R2208 B.n1404 B.n99 30.6877
R2209 B.n1398 B.n99 30.6877
R2210 B.n1398 B.n1397 30.6877
R2211 B.n1396 B.n106 30.6877
R2212 B.n1390 B.n106 30.6877
R2213 B.n1390 B.n1389 30.6877
R2214 B.n1389 B.n1388 30.6877
R2215 B.n1388 B.n113 30.6877
R2216 B.n1382 B.n113 30.6877
R2217 B.n1382 B.n1381 30.6877
R2218 B.n1381 B.n1380 30.6877
R2219 B.n1380 B.n120 30.6877
R2220 B.n1374 B.n120 30.6877
R2221 B.n1374 B.n1373 30.6877
R2222 B.n1373 B.n1372 30.6877
R2223 B.n1372 B.n127 30.6877
R2224 B.n1366 B.n127 30.6877
R2225 B.n1365 B.n1364 30.6877
R2226 B.n1364 B.n134 30.6877
R2227 B.n1358 B.n134 30.6877
R2228 B.n1358 B.n1357 30.6877
R2229 B.n1357 B.n1356 30.6877
R2230 B.n1356 B.n141 30.6877
R2231 B.n1350 B.n141 30.6877
R2232 B.n1350 B.n1349 30.6877
R2233 B.n1349 B.n1348 30.6877
R2234 B.n263 B.t9 26.6261
R2235 B.t3 B.n1469 26.6261
R2236 B.n841 B.t0 25.7236
R2237 B.n1422 B.t8 25.7236
R2238 B.n799 B.t6 24.821
R2239 B.t5 B.n1396 24.821
R2240 B.t2 B.n231 23.9184
R2241 B.t7 B.n15 23.9184
R2242 B.n757 B.t11 23.0159
R2243 B.n1366 B.t15 23.0159
R2244 B B.n1512 18.0485
R2245 B.n287 B.t4 15.7954
R2246 B.t1 B.n1445 15.7954
R2247 B.n877 B.t4 14.8928
R2248 B.n1446 B.t1 14.8928
R2249 B.n1345 B.n1344 10.6151
R2250 B.n1344 B.n150 10.6151
R2251 B.n1338 B.n150 10.6151
R2252 B.n1338 B.n1337 10.6151
R2253 B.n1337 B.n1336 10.6151
R2254 B.n1336 B.n152 10.6151
R2255 B.n1330 B.n152 10.6151
R2256 B.n1330 B.n1329 10.6151
R2257 B.n1329 B.n1328 10.6151
R2258 B.n1328 B.n154 10.6151
R2259 B.n1322 B.n154 10.6151
R2260 B.n1322 B.n1321 10.6151
R2261 B.n1321 B.n1320 10.6151
R2262 B.n1320 B.n156 10.6151
R2263 B.n1314 B.n156 10.6151
R2264 B.n1314 B.n1313 10.6151
R2265 B.n1313 B.n1312 10.6151
R2266 B.n1312 B.n158 10.6151
R2267 B.n1306 B.n158 10.6151
R2268 B.n1306 B.n1305 10.6151
R2269 B.n1305 B.n1304 10.6151
R2270 B.n1304 B.n160 10.6151
R2271 B.n1298 B.n160 10.6151
R2272 B.n1298 B.n1297 10.6151
R2273 B.n1297 B.n1296 10.6151
R2274 B.n1296 B.n162 10.6151
R2275 B.n1290 B.n162 10.6151
R2276 B.n1290 B.n1289 10.6151
R2277 B.n1289 B.n1288 10.6151
R2278 B.n1288 B.n164 10.6151
R2279 B.n1282 B.n164 10.6151
R2280 B.n1282 B.n1281 10.6151
R2281 B.n1281 B.n1280 10.6151
R2282 B.n1280 B.n166 10.6151
R2283 B.n1274 B.n166 10.6151
R2284 B.n1274 B.n1273 10.6151
R2285 B.n1273 B.n1272 10.6151
R2286 B.n1272 B.n168 10.6151
R2287 B.n1266 B.n168 10.6151
R2288 B.n1266 B.n1265 10.6151
R2289 B.n1265 B.n1264 10.6151
R2290 B.n1264 B.n170 10.6151
R2291 B.n1258 B.n170 10.6151
R2292 B.n1258 B.n1257 10.6151
R2293 B.n1257 B.n1256 10.6151
R2294 B.n1256 B.n172 10.6151
R2295 B.n1250 B.n172 10.6151
R2296 B.n1250 B.n1249 10.6151
R2297 B.n1249 B.n1248 10.6151
R2298 B.n1248 B.n174 10.6151
R2299 B.n1242 B.n174 10.6151
R2300 B.n1242 B.n1241 10.6151
R2301 B.n1241 B.n1240 10.6151
R2302 B.n1240 B.n176 10.6151
R2303 B.n1234 B.n176 10.6151
R2304 B.n1234 B.n1233 10.6151
R2305 B.n1233 B.n1232 10.6151
R2306 B.n1232 B.n178 10.6151
R2307 B.n1226 B.n178 10.6151
R2308 B.n1226 B.n1225 10.6151
R2309 B.n1225 B.n1224 10.6151
R2310 B.n1224 B.n180 10.6151
R2311 B.n1218 B.n1217 10.6151
R2312 B.n1217 B.n1216 10.6151
R2313 B.n1216 B.n185 10.6151
R2314 B.n1210 B.n185 10.6151
R2315 B.n1210 B.n1209 10.6151
R2316 B.n1209 B.n1208 10.6151
R2317 B.n1208 B.n187 10.6151
R2318 B.n1202 B.n187 10.6151
R2319 B.n1200 B.n1199 10.6151
R2320 B.n1199 B.n191 10.6151
R2321 B.n1193 B.n191 10.6151
R2322 B.n1193 B.n1192 10.6151
R2323 B.n1192 B.n1191 10.6151
R2324 B.n1191 B.n193 10.6151
R2325 B.n1185 B.n193 10.6151
R2326 B.n1185 B.n1184 10.6151
R2327 B.n1184 B.n1183 10.6151
R2328 B.n1183 B.n195 10.6151
R2329 B.n1177 B.n195 10.6151
R2330 B.n1177 B.n1176 10.6151
R2331 B.n1176 B.n1175 10.6151
R2332 B.n1175 B.n197 10.6151
R2333 B.n1169 B.n197 10.6151
R2334 B.n1169 B.n1168 10.6151
R2335 B.n1168 B.n1167 10.6151
R2336 B.n1167 B.n199 10.6151
R2337 B.n1161 B.n199 10.6151
R2338 B.n1161 B.n1160 10.6151
R2339 B.n1160 B.n1159 10.6151
R2340 B.n1159 B.n201 10.6151
R2341 B.n1153 B.n201 10.6151
R2342 B.n1153 B.n1152 10.6151
R2343 B.n1152 B.n1151 10.6151
R2344 B.n1151 B.n203 10.6151
R2345 B.n1145 B.n203 10.6151
R2346 B.n1145 B.n1144 10.6151
R2347 B.n1144 B.n1143 10.6151
R2348 B.n1143 B.n205 10.6151
R2349 B.n1137 B.n205 10.6151
R2350 B.n1137 B.n1136 10.6151
R2351 B.n1136 B.n1135 10.6151
R2352 B.n1135 B.n207 10.6151
R2353 B.n1129 B.n207 10.6151
R2354 B.n1129 B.n1128 10.6151
R2355 B.n1128 B.n1127 10.6151
R2356 B.n1127 B.n209 10.6151
R2357 B.n1121 B.n209 10.6151
R2358 B.n1121 B.n1120 10.6151
R2359 B.n1120 B.n1119 10.6151
R2360 B.n1119 B.n211 10.6151
R2361 B.n1113 B.n211 10.6151
R2362 B.n1113 B.n1112 10.6151
R2363 B.n1112 B.n1111 10.6151
R2364 B.n1111 B.n213 10.6151
R2365 B.n1105 B.n213 10.6151
R2366 B.n1105 B.n1104 10.6151
R2367 B.n1104 B.n1103 10.6151
R2368 B.n1103 B.n215 10.6151
R2369 B.n1097 B.n215 10.6151
R2370 B.n1097 B.n1096 10.6151
R2371 B.n1096 B.n1095 10.6151
R2372 B.n1095 B.n217 10.6151
R2373 B.n1089 B.n217 10.6151
R2374 B.n1089 B.n1088 10.6151
R2375 B.n1088 B.n1087 10.6151
R2376 B.n1087 B.n219 10.6151
R2377 B.n1081 B.n219 10.6151
R2378 B.n1081 B.n1080 10.6151
R2379 B.n1080 B.n1079 10.6151
R2380 B.n1079 B.n1075 10.6151
R2381 B.n730 B.n729 10.6151
R2382 B.n731 B.n730 10.6151
R2383 B.n731 B.n373 10.6151
R2384 B.n741 B.n373 10.6151
R2385 B.n742 B.n741 10.6151
R2386 B.n743 B.n742 10.6151
R2387 B.n743 B.n364 10.6151
R2388 B.n753 B.n364 10.6151
R2389 B.n754 B.n753 10.6151
R2390 B.n755 B.n754 10.6151
R2391 B.n755 B.n357 10.6151
R2392 B.n765 B.n357 10.6151
R2393 B.n766 B.n765 10.6151
R2394 B.n767 B.n766 10.6151
R2395 B.n767 B.n349 10.6151
R2396 B.n777 B.n349 10.6151
R2397 B.n778 B.n777 10.6151
R2398 B.n779 B.n778 10.6151
R2399 B.n779 B.n341 10.6151
R2400 B.n789 B.n341 10.6151
R2401 B.n790 B.n789 10.6151
R2402 B.n791 B.n790 10.6151
R2403 B.n791 B.n333 10.6151
R2404 B.n801 B.n333 10.6151
R2405 B.n802 B.n801 10.6151
R2406 B.n803 B.n802 10.6151
R2407 B.n803 B.n325 10.6151
R2408 B.n813 B.n325 10.6151
R2409 B.n814 B.n813 10.6151
R2410 B.n815 B.n814 10.6151
R2411 B.n815 B.n317 10.6151
R2412 B.n825 B.n317 10.6151
R2413 B.n826 B.n825 10.6151
R2414 B.n827 B.n826 10.6151
R2415 B.n827 B.n308 10.6151
R2416 B.n837 B.n308 10.6151
R2417 B.n838 B.n837 10.6151
R2418 B.n839 B.n838 10.6151
R2419 B.n839 B.n301 10.6151
R2420 B.n849 B.n301 10.6151
R2421 B.n850 B.n849 10.6151
R2422 B.n851 B.n850 10.6151
R2423 B.n851 B.n293 10.6151
R2424 B.n861 B.n293 10.6151
R2425 B.n862 B.n861 10.6151
R2426 B.n863 B.n862 10.6151
R2427 B.n863 B.n284 10.6151
R2428 B.n873 B.n284 10.6151
R2429 B.n874 B.n873 10.6151
R2430 B.n875 B.n874 10.6151
R2431 B.n875 B.n277 10.6151
R2432 B.n885 B.n277 10.6151
R2433 B.n886 B.n885 10.6151
R2434 B.n887 B.n886 10.6151
R2435 B.n887 B.n269 10.6151
R2436 B.n897 B.n269 10.6151
R2437 B.n898 B.n897 10.6151
R2438 B.n899 B.n898 10.6151
R2439 B.n899 B.n260 10.6151
R2440 B.n909 B.n260 10.6151
R2441 B.n910 B.n909 10.6151
R2442 B.n911 B.n910 10.6151
R2443 B.n911 B.n253 10.6151
R2444 B.n921 B.n253 10.6151
R2445 B.n922 B.n921 10.6151
R2446 B.n923 B.n922 10.6151
R2447 B.n923 B.n245 10.6151
R2448 B.n933 B.n245 10.6151
R2449 B.n934 B.n933 10.6151
R2450 B.n935 B.n934 10.6151
R2451 B.n935 B.n237 10.6151
R2452 B.n945 B.n237 10.6151
R2453 B.n946 B.n945 10.6151
R2454 B.n947 B.n946 10.6151
R2455 B.n947 B.n229 10.6151
R2456 B.n957 B.n229 10.6151
R2457 B.n958 B.n957 10.6151
R2458 B.n960 B.n958 10.6151
R2459 B.n960 B.n959 10.6151
R2460 B.n959 B.n221 10.6151
R2461 B.n971 B.n221 10.6151
R2462 B.n972 B.n971 10.6151
R2463 B.n973 B.n972 10.6151
R2464 B.n974 B.n973 10.6151
R2465 B.n976 B.n974 10.6151
R2466 B.n977 B.n976 10.6151
R2467 B.n978 B.n977 10.6151
R2468 B.n979 B.n978 10.6151
R2469 B.n981 B.n979 10.6151
R2470 B.n982 B.n981 10.6151
R2471 B.n983 B.n982 10.6151
R2472 B.n984 B.n983 10.6151
R2473 B.n986 B.n984 10.6151
R2474 B.n987 B.n986 10.6151
R2475 B.n988 B.n987 10.6151
R2476 B.n989 B.n988 10.6151
R2477 B.n991 B.n989 10.6151
R2478 B.n992 B.n991 10.6151
R2479 B.n993 B.n992 10.6151
R2480 B.n994 B.n993 10.6151
R2481 B.n996 B.n994 10.6151
R2482 B.n997 B.n996 10.6151
R2483 B.n998 B.n997 10.6151
R2484 B.n999 B.n998 10.6151
R2485 B.n1001 B.n999 10.6151
R2486 B.n1002 B.n1001 10.6151
R2487 B.n1003 B.n1002 10.6151
R2488 B.n1004 B.n1003 10.6151
R2489 B.n1006 B.n1004 10.6151
R2490 B.n1007 B.n1006 10.6151
R2491 B.n1008 B.n1007 10.6151
R2492 B.n1009 B.n1008 10.6151
R2493 B.n1011 B.n1009 10.6151
R2494 B.n1012 B.n1011 10.6151
R2495 B.n1013 B.n1012 10.6151
R2496 B.n1014 B.n1013 10.6151
R2497 B.n1016 B.n1014 10.6151
R2498 B.n1017 B.n1016 10.6151
R2499 B.n1018 B.n1017 10.6151
R2500 B.n1019 B.n1018 10.6151
R2501 B.n1021 B.n1019 10.6151
R2502 B.n1022 B.n1021 10.6151
R2503 B.n1023 B.n1022 10.6151
R2504 B.n1024 B.n1023 10.6151
R2505 B.n1026 B.n1024 10.6151
R2506 B.n1027 B.n1026 10.6151
R2507 B.n1028 B.n1027 10.6151
R2508 B.n1029 B.n1028 10.6151
R2509 B.n1031 B.n1029 10.6151
R2510 B.n1032 B.n1031 10.6151
R2511 B.n1033 B.n1032 10.6151
R2512 B.n1034 B.n1033 10.6151
R2513 B.n1036 B.n1034 10.6151
R2514 B.n1037 B.n1036 10.6151
R2515 B.n1038 B.n1037 10.6151
R2516 B.n1039 B.n1038 10.6151
R2517 B.n1041 B.n1039 10.6151
R2518 B.n1042 B.n1041 10.6151
R2519 B.n1043 B.n1042 10.6151
R2520 B.n1044 B.n1043 10.6151
R2521 B.n1046 B.n1044 10.6151
R2522 B.n1047 B.n1046 10.6151
R2523 B.n1048 B.n1047 10.6151
R2524 B.n1049 B.n1048 10.6151
R2525 B.n1051 B.n1049 10.6151
R2526 B.n1052 B.n1051 10.6151
R2527 B.n1053 B.n1052 10.6151
R2528 B.n1054 B.n1053 10.6151
R2529 B.n1056 B.n1054 10.6151
R2530 B.n1057 B.n1056 10.6151
R2531 B.n1058 B.n1057 10.6151
R2532 B.n1059 B.n1058 10.6151
R2533 B.n1061 B.n1059 10.6151
R2534 B.n1062 B.n1061 10.6151
R2535 B.n1063 B.n1062 10.6151
R2536 B.n1064 B.n1063 10.6151
R2537 B.n1066 B.n1064 10.6151
R2538 B.n1067 B.n1066 10.6151
R2539 B.n1068 B.n1067 10.6151
R2540 B.n1069 B.n1068 10.6151
R2541 B.n1071 B.n1069 10.6151
R2542 B.n1072 B.n1071 10.6151
R2543 B.n1073 B.n1072 10.6151
R2544 B.n1074 B.n1073 10.6151
R2545 B.n724 B.n723 10.6151
R2546 B.n723 B.n385 10.6151
R2547 B.n718 B.n385 10.6151
R2548 B.n718 B.n717 10.6151
R2549 B.n717 B.n387 10.6151
R2550 B.n712 B.n387 10.6151
R2551 B.n712 B.n711 10.6151
R2552 B.n711 B.n710 10.6151
R2553 B.n710 B.n389 10.6151
R2554 B.n704 B.n389 10.6151
R2555 B.n704 B.n703 10.6151
R2556 B.n703 B.n702 10.6151
R2557 B.n702 B.n391 10.6151
R2558 B.n696 B.n391 10.6151
R2559 B.n696 B.n695 10.6151
R2560 B.n695 B.n694 10.6151
R2561 B.n694 B.n393 10.6151
R2562 B.n688 B.n393 10.6151
R2563 B.n688 B.n687 10.6151
R2564 B.n687 B.n686 10.6151
R2565 B.n686 B.n395 10.6151
R2566 B.n680 B.n395 10.6151
R2567 B.n680 B.n679 10.6151
R2568 B.n679 B.n678 10.6151
R2569 B.n678 B.n397 10.6151
R2570 B.n672 B.n397 10.6151
R2571 B.n672 B.n671 10.6151
R2572 B.n671 B.n670 10.6151
R2573 B.n670 B.n399 10.6151
R2574 B.n664 B.n399 10.6151
R2575 B.n664 B.n663 10.6151
R2576 B.n663 B.n662 10.6151
R2577 B.n662 B.n401 10.6151
R2578 B.n656 B.n401 10.6151
R2579 B.n656 B.n655 10.6151
R2580 B.n655 B.n654 10.6151
R2581 B.n654 B.n403 10.6151
R2582 B.n648 B.n403 10.6151
R2583 B.n648 B.n647 10.6151
R2584 B.n647 B.n646 10.6151
R2585 B.n646 B.n405 10.6151
R2586 B.n640 B.n405 10.6151
R2587 B.n640 B.n639 10.6151
R2588 B.n639 B.n638 10.6151
R2589 B.n638 B.n407 10.6151
R2590 B.n632 B.n407 10.6151
R2591 B.n632 B.n631 10.6151
R2592 B.n631 B.n630 10.6151
R2593 B.n630 B.n409 10.6151
R2594 B.n624 B.n409 10.6151
R2595 B.n624 B.n623 10.6151
R2596 B.n623 B.n622 10.6151
R2597 B.n622 B.n411 10.6151
R2598 B.n616 B.n411 10.6151
R2599 B.n616 B.n615 10.6151
R2600 B.n615 B.n614 10.6151
R2601 B.n614 B.n413 10.6151
R2602 B.n608 B.n413 10.6151
R2603 B.n608 B.n607 10.6151
R2604 B.n607 B.n606 10.6151
R2605 B.n606 B.n415 10.6151
R2606 B.n600 B.n415 10.6151
R2607 B.n598 B.n597 10.6151
R2608 B.n597 B.n419 10.6151
R2609 B.n591 B.n419 10.6151
R2610 B.n591 B.n590 10.6151
R2611 B.n590 B.n589 10.6151
R2612 B.n589 B.n421 10.6151
R2613 B.n583 B.n421 10.6151
R2614 B.n583 B.n582 10.6151
R2615 B.n580 B.n425 10.6151
R2616 B.n574 B.n425 10.6151
R2617 B.n574 B.n573 10.6151
R2618 B.n573 B.n572 10.6151
R2619 B.n572 B.n427 10.6151
R2620 B.n566 B.n427 10.6151
R2621 B.n566 B.n565 10.6151
R2622 B.n565 B.n564 10.6151
R2623 B.n564 B.n429 10.6151
R2624 B.n558 B.n429 10.6151
R2625 B.n558 B.n557 10.6151
R2626 B.n557 B.n556 10.6151
R2627 B.n556 B.n431 10.6151
R2628 B.n550 B.n431 10.6151
R2629 B.n550 B.n549 10.6151
R2630 B.n549 B.n548 10.6151
R2631 B.n548 B.n433 10.6151
R2632 B.n542 B.n433 10.6151
R2633 B.n542 B.n541 10.6151
R2634 B.n541 B.n540 10.6151
R2635 B.n540 B.n435 10.6151
R2636 B.n534 B.n435 10.6151
R2637 B.n534 B.n533 10.6151
R2638 B.n533 B.n532 10.6151
R2639 B.n532 B.n437 10.6151
R2640 B.n526 B.n437 10.6151
R2641 B.n526 B.n525 10.6151
R2642 B.n525 B.n524 10.6151
R2643 B.n524 B.n439 10.6151
R2644 B.n518 B.n439 10.6151
R2645 B.n518 B.n517 10.6151
R2646 B.n517 B.n516 10.6151
R2647 B.n516 B.n441 10.6151
R2648 B.n510 B.n441 10.6151
R2649 B.n510 B.n509 10.6151
R2650 B.n509 B.n508 10.6151
R2651 B.n508 B.n443 10.6151
R2652 B.n502 B.n443 10.6151
R2653 B.n502 B.n501 10.6151
R2654 B.n501 B.n500 10.6151
R2655 B.n500 B.n445 10.6151
R2656 B.n494 B.n445 10.6151
R2657 B.n494 B.n493 10.6151
R2658 B.n493 B.n492 10.6151
R2659 B.n492 B.n447 10.6151
R2660 B.n486 B.n447 10.6151
R2661 B.n486 B.n485 10.6151
R2662 B.n485 B.n484 10.6151
R2663 B.n484 B.n449 10.6151
R2664 B.n478 B.n449 10.6151
R2665 B.n478 B.n477 10.6151
R2666 B.n477 B.n476 10.6151
R2667 B.n476 B.n451 10.6151
R2668 B.n470 B.n451 10.6151
R2669 B.n470 B.n469 10.6151
R2670 B.n469 B.n468 10.6151
R2671 B.n468 B.n453 10.6151
R2672 B.n462 B.n453 10.6151
R2673 B.n462 B.n461 10.6151
R2674 B.n461 B.n460 10.6151
R2675 B.n460 B.n455 10.6151
R2676 B.n455 B.n381 10.6151
R2677 B.n725 B.n377 10.6151
R2678 B.n735 B.n377 10.6151
R2679 B.n736 B.n735 10.6151
R2680 B.n737 B.n736 10.6151
R2681 B.n737 B.n369 10.6151
R2682 B.n747 B.n369 10.6151
R2683 B.n748 B.n747 10.6151
R2684 B.n749 B.n748 10.6151
R2685 B.n749 B.n361 10.6151
R2686 B.n759 B.n361 10.6151
R2687 B.n760 B.n759 10.6151
R2688 B.n761 B.n760 10.6151
R2689 B.n761 B.n353 10.6151
R2690 B.n771 B.n353 10.6151
R2691 B.n772 B.n771 10.6151
R2692 B.n773 B.n772 10.6151
R2693 B.n773 B.n345 10.6151
R2694 B.n783 B.n345 10.6151
R2695 B.n784 B.n783 10.6151
R2696 B.n785 B.n784 10.6151
R2697 B.n785 B.n337 10.6151
R2698 B.n795 B.n337 10.6151
R2699 B.n796 B.n795 10.6151
R2700 B.n797 B.n796 10.6151
R2701 B.n797 B.n329 10.6151
R2702 B.n807 B.n329 10.6151
R2703 B.n808 B.n807 10.6151
R2704 B.n809 B.n808 10.6151
R2705 B.n809 B.n321 10.6151
R2706 B.n819 B.n321 10.6151
R2707 B.n820 B.n819 10.6151
R2708 B.n821 B.n820 10.6151
R2709 B.n821 B.n313 10.6151
R2710 B.n831 B.n313 10.6151
R2711 B.n832 B.n831 10.6151
R2712 B.n833 B.n832 10.6151
R2713 B.n833 B.n305 10.6151
R2714 B.n843 B.n305 10.6151
R2715 B.n844 B.n843 10.6151
R2716 B.n845 B.n844 10.6151
R2717 B.n845 B.n297 10.6151
R2718 B.n855 B.n297 10.6151
R2719 B.n856 B.n855 10.6151
R2720 B.n857 B.n856 10.6151
R2721 B.n857 B.n289 10.6151
R2722 B.n867 B.n289 10.6151
R2723 B.n868 B.n867 10.6151
R2724 B.n869 B.n868 10.6151
R2725 B.n869 B.n281 10.6151
R2726 B.n879 B.n281 10.6151
R2727 B.n880 B.n879 10.6151
R2728 B.n881 B.n880 10.6151
R2729 B.n881 B.n273 10.6151
R2730 B.n891 B.n273 10.6151
R2731 B.n892 B.n891 10.6151
R2732 B.n893 B.n892 10.6151
R2733 B.n893 B.n265 10.6151
R2734 B.n903 B.n265 10.6151
R2735 B.n904 B.n903 10.6151
R2736 B.n905 B.n904 10.6151
R2737 B.n905 B.n257 10.6151
R2738 B.n915 B.n257 10.6151
R2739 B.n916 B.n915 10.6151
R2740 B.n917 B.n916 10.6151
R2741 B.n917 B.n249 10.6151
R2742 B.n927 B.n249 10.6151
R2743 B.n928 B.n927 10.6151
R2744 B.n929 B.n928 10.6151
R2745 B.n929 B.n241 10.6151
R2746 B.n939 B.n241 10.6151
R2747 B.n940 B.n939 10.6151
R2748 B.n941 B.n940 10.6151
R2749 B.n941 B.n233 10.6151
R2750 B.n951 B.n233 10.6151
R2751 B.n952 B.n951 10.6151
R2752 B.n953 B.n952 10.6151
R2753 B.n953 B.n225 10.6151
R2754 B.n964 B.n225 10.6151
R2755 B.n965 B.n964 10.6151
R2756 B.n966 B.n965 10.6151
R2757 B.n966 B.n0 10.6151
R2758 B.n1506 B.n1 10.6151
R2759 B.n1506 B.n1505 10.6151
R2760 B.n1505 B.n1504 10.6151
R2761 B.n1504 B.n10 10.6151
R2762 B.n1498 B.n10 10.6151
R2763 B.n1498 B.n1497 10.6151
R2764 B.n1497 B.n1496 10.6151
R2765 B.n1496 B.n17 10.6151
R2766 B.n1490 B.n17 10.6151
R2767 B.n1490 B.n1489 10.6151
R2768 B.n1489 B.n1488 10.6151
R2769 B.n1488 B.n24 10.6151
R2770 B.n1482 B.n24 10.6151
R2771 B.n1482 B.n1481 10.6151
R2772 B.n1481 B.n1480 10.6151
R2773 B.n1480 B.n31 10.6151
R2774 B.n1474 B.n31 10.6151
R2775 B.n1474 B.n1473 10.6151
R2776 B.n1473 B.n1472 10.6151
R2777 B.n1472 B.n38 10.6151
R2778 B.n1466 B.n38 10.6151
R2779 B.n1466 B.n1465 10.6151
R2780 B.n1465 B.n1464 10.6151
R2781 B.n1464 B.n45 10.6151
R2782 B.n1458 B.n45 10.6151
R2783 B.n1458 B.n1457 10.6151
R2784 B.n1457 B.n1456 10.6151
R2785 B.n1456 B.n52 10.6151
R2786 B.n1450 B.n52 10.6151
R2787 B.n1450 B.n1449 10.6151
R2788 B.n1449 B.n1448 10.6151
R2789 B.n1448 B.n59 10.6151
R2790 B.n1442 B.n59 10.6151
R2791 B.n1442 B.n1441 10.6151
R2792 B.n1441 B.n1440 10.6151
R2793 B.n1440 B.n66 10.6151
R2794 B.n1434 B.n66 10.6151
R2795 B.n1434 B.n1433 10.6151
R2796 B.n1433 B.n1432 10.6151
R2797 B.n1432 B.n73 10.6151
R2798 B.n1426 B.n73 10.6151
R2799 B.n1426 B.n1425 10.6151
R2800 B.n1425 B.n1424 10.6151
R2801 B.n1424 B.n80 10.6151
R2802 B.n1418 B.n80 10.6151
R2803 B.n1418 B.n1417 10.6151
R2804 B.n1417 B.n1416 10.6151
R2805 B.n1416 B.n87 10.6151
R2806 B.n1410 B.n87 10.6151
R2807 B.n1410 B.n1409 10.6151
R2808 B.n1409 B.n1408 10.6151
R2809 B.n1408 B.n94 10.6151
R2810 B.n1402 B.n94 10.6151
R2811 B.n1402 B.n1401 10.6151
R2812 B.n1401 B.n1400 10.6151
R2813 B.n1400 B.n101 10.6151
R2814 B.n1394 B.n101 10.6151
R2815 B.n1394 B.n1393 10.6151
R2816 B.n1393 B.n1392 10.6151
R2817 B.n1392 B.n108 10.6151
R2818 B.n1386 B.n108 10.6151
R2819 B.n1386 B.n1385 10.6151
R2820 B.n1385 B.n1384 10.6151
R2821 B.n1384 B.n115 10.6151
R2822 B.n1378 B.n115 10.6151
R2823 B.n1378 B.n1377 10.6151
R2824 B.n1377 B.n1376 10.6151
R2825 B.n1376 B.n122 10.6151
R2826 B.n1370 B.n122 10.6151
R2827 B.n1370 B.n1369 10.6151
R2828 B.n1369 B.n1368 10.6151
R2829 B.n1368 B.n129 10.6151
R2830 B.n1362 B.n129 10.6151
R2831 B.n1362 B.n1361 10.6151
R2832 B.n1361 B.n1360 10.6151
R2833 B.n1360 B.n136 10.6151
R2834 B.n1354 B.n136 10.6151
R2835 B.n1354 B.n1353 10.6151
R2836 B.n1353 B.n1352 10.6151
R2837 B.n1352 B.n143 10.6151
R2838 B.n1346 B.n143 10.6151
R2839 B.n367 B.t11 7.67229
R2840 B.t15 B.n1365 7.67229
R2841 B.n949 B.t2 6.76973
R2842 B.n1494 B.t7 6.76973
R2843 B.n1218 B.n184 6.5566
R2844 B.n1202 B.n1201 6.5566
R2845 B.n599 B.n598 6.5566
R2846 B.n582 B.n581 6.5566
R2847 B.t6 B.n331 5.86717
R2848 B.n1397 B.t5 5.86717
R2849 B.n311 B.t0 4.9646
R2850 B.t8 B.n1421 4.9646
R2851 B.n913 B.t9 4.06204
R2852 B.n1470 B.t3 4.06204
R2853 B.n184 B.n180 4.05904
R2854 B.n1201 B.n1200 4.05904
R2855 B.n600 B.n599 4.05904
R2856 B.n581 B.n580 4.05904
R2857 B.n1512 B.n0 2.81026
R2858 B.n1512 B.n1 2.81026
R2859 VN.n107 VN.n55 161.3
R2860 VN.n106 VN.n105 161.3
R2861 VN.n104 VN.n56 161.3
R2862 VN.n103 VN.n102 161.3
R2863 VN.n101 VN.n57 161.3
R2864 VN.n100 VN.n99 161.3
R2865 VN.n98 VN.n58 161.3
R2866 VN.n97 VN.n96 161.3
R2867 VN.n94 VN.n59 161.3
R2868 VN.n93 VN.n92 161.3
R2869 VN.n91 VN.n60 161.3
R2870 VN.n90 VN.n89 161.3
R2871 VN.n88 VN.n61 161.3
R2872 VN.n87 VN.n86 161.3
R2873 VN.n85 VN.n62 161.3
R2874 VN.n84 VN.n83 161.3
R2875 VN.n82 VN.n63 161.3
R2876 VN.n81 VN.n80 161.3
R2877 VN.n79 VN.n64 161.3
R2878 VN.n78 VN.n77 161.3
R2879 VN.n76 VN.n65 161.3
R2880 VN.n75 VN.n74 161.3
R2881 VN.n73 VN.n66 161.3
R2882 VN.n72 VN.n71 161.3
R2883 VN.n70 VN.n67 161.3
R2884 VN.n52 VN.n0 161.3
R2885 VN.n51 VN.n50 161.3
R2886 VN.n49 VN.n1 161.3
R2887 VN.n48 VN.n47 161.3
R2888 VN.n46 VN.n2 161.3
R2889 VN.n45 VN.n44 161.3
R2890 VN.n43 VN.n3 161.3
R2891 VN.n42 VN.n41 161.3
R2892 VN.n39 VN.n4 161.3
R2893 VN.n38 VN.n37 161.3
R2894 VN.n36 VN.n5 161.3
R2895 VN.n35 VN.n34 161.3
R2896 VN.n33 VN.n6 161.3
R2897 VN.n32 VN.n31 161.3
R2898 VN.n30 VN.n7 161.3
R2899 VN.n29 VN.n28 161.3
R2900 VN.n27 VN.n8 161.3
R2901 VN.n26 VN.n25 161.3
R2902 VN.n24 VN.n9 161.3
R2903 VN.n23 VN.n22 161.3
R2904 VN.n21 VN.n10 161.3
R2905 VN.n20 VN.n19 161.3
R2906 VN.n18 VN.n11 161.3
R2907 VN.n17 VN.n16 161.3
R2908 VN.n15 VN.n12 161.3
R2909 VN.n13 VN.t9 151.149
R2910 VN.n68 VN.t7 151.149
R2911 VN.n27 VN.t5 118.944
R2912 VN.n14 VN.t3 118.944
R2913 VN.n40 VN.t8 118.944
R2914 VN.n53 VN.t1 118.944
R2915 VN.n82 VN.t2 118.944
R2916 VN.n69 VN.t4 118.944
R2917 VN.n95 VN.t6 118.944
R2918 VN.n108 VN.t0 118.944
R2919 VN VN.n109 65.6403
R2920 VN.n14 VN.n13 65.0774
R2921 VN.n69 VN.n68 65.0774
R2922 VN.n54 VN.n53 62.5108
R2923 VN.n109 VN.n108 62.5108
R2924 VN.n47 VN.n46 56.4773
R2925 VN.n102 VN.n101 56.4773
R2926 VN.n21 VN.n20 50.148
R2927 VN.n34 VN.n33 50.148
R2928 VN.n76 VN.n75 50.148
R2929 VN.n89 VN.n88 50.148
R2930 VN.n22 VN.n21 30.6732
R2931 VN.n33 VN.n32 30.6732
R2932 VN.n77 VN.n76 30.6732
R2933 VN.n88 VN.n87 30.6732
R2934 VN.n16 VN.n15 24.3439
R2935 VN.n16 VN.n11 24.3439
R2936 VN.n20 VN.n11 24.3439
R2937 VN.n22 VN.n9 24.3439
R2938 VN.n26 VN.n9 24.3439
R2939 VN.n27 VN.n26 24.3439
R2940 VN.n28 VN.n27 24.3439
R2941 VN.n28 VN.n7 24.3439
R2942 VN.n32 VN.n7 24.3439
R2943 VN.n34 VN.n5 24.3439
R2944 VN.n38 VN.n5 24.3439
R2945 VN.n39 VN.n38 24.3439
R2946 VN.n41 VN.n3 24.3439
R2947 VN.n45 VN.n3 24.3439
R2948 VN.n46 VN.n45 24.3439
R2949 VN.n47 VN.n1 24.3439
R2950 VN.n51 VN.n1 24.3439
R2951 VN.n52 VN.n51 24.3439
R2952 VN.n75 VN.n66 24.3439
R2953 VN.n71 VN.n66 24.3439
R2954 VN.n71 VN.n70 24.3439
R2955 VN.n87 VN.n62 24.3439
R2956 VN.n83 VN.n62 24.3439
R2957 VN.n83 VN.n82 24.3439
R2958 VN.n82 VN.n81 24.3439
R2959 VN.n81 VN.n64 24.3439
R2960 VN.n77 VN.n64 24.3439
R2961 VN.n101 VN.n100 24.3439
R2962 VN.n100 VN.n58 24.3439
R2963 VN.n96 VN.n58 24.3439
R2964 VN.n94 VN.n93 24.3439
R2965 VN.n93 VN.n60 24.3439
R2966 VN.n89 VN.n60 24.3439
R2967 VN.n107 VN.n106 24.3439
R2968 VN.n106 VN.n56 24.3439
R2969 VN.n102 VN.n56 24.3439
R2970 VN.n53 VN.n52 19.4752
R2971 VN.n108 VN.n107 19.4752
R2972 VN.n41 VN.n40 14.6066
R2973 VN.n96 VN.n95 14.6066
R2974 VN.n15 VN.n14 9.73787
R2975 VN.n40 VN.n39 9.73787
R2976 VN.n70 VN.n69 9.73787
R2977 VN.n95 VN.n94 9.73787
R2978 VN.n68 VN.n67 2.72005
R2979 VN.n13 VN.n12 2.72005
R2980 VN.n109 VN.n55 0.417764
R2981 VN.n54 VN.n0 0.417764
R2982 VN VN.n54 0.394061
R2983 VN.n105 VN.n55 0.189894
R2984 VN.n105 VN.n104 0.189894
R2985 VN.n104 VN.n103 0.189894
R2986 VN.n103 VN.n57 0.189894
R2987 VN.n99 VN.n57 0.189894
R2988 VN.n99 VN.n98 0.189894
R2989 VN.n98 VN.n97 0.189894
R2990 VN.n97 VN.n59 0.189894
R2991 VN.n92 VN.n59 0.189894
R2992 VN.n92 VN.n91 0.189894
R2993 VN.n91 VN.n90 0.189894
R2994 VN.n90 VN.n61 0.189894
R2995 VN.n86 VN.n61 0.189894
R2996 VN.n86 VN.n85 0.189894
R2997 VN.n85 VN.n84 0.189894
R2998 VN.n84 VN.n63 0.189894
R2999 VN.n80 VN.n63 0.189894
R3000 VN.n80 VN.n79 0.189894
R3001 VN.n79 VN.n78 0.189894
R3002 VN.n78 VN.n65 0.189894
R3003 VN.n74 VN.n65 0.189894
R3004 VN.n74 VN.n73 0.189894
R3005 VN.n73 VN.n72 0.189894
R3006 VN.n72 VN.n67 0.189894
R3007 VN.n17 VN.n12 0.189894
R3008 VN.n18 VN.n17 0.189894
R3009 VN.n19 VN.n18 0.189894
R3010 VN.n19 VN.n10 0.189894
R3011 VN.n23 VN.n10 0.189894
R3012 VN.n24 VN.n23 0.189894
R3013 VN.n25 VN.n24 0.189894
R3014 VN.n25 VN.n8 0.189894
R3015 VN.n29 VN.n8 0.189894
R3016 VN.n30 VN.n29 0.189894
R3017 VN.n31 VN.n30 0.189894
R3018 VN.n31 VN.n6 0.189894
R3019 VN.n35 VN.n6 0.189894
R3020 VN.n36 VN.n35 0.189894
R3021 VN.n37 VN.n36 0.189894
R3022 VN.n37 VN.n4 0.189894
R3023 VN.n42 VN.n4 0.189894
R3024 VN.n43 VN.n42 0.189894
R3025 VN.n44 VN.n43 0.189894
R3026 VN.n44 VN.n2 0.189894
R3027 VN.n48 VN.n2 0.189894
R3028 VN.n49 VN.n48 0.189894
R3029 VN.n50 VN.n49 0.189894
R3030 VN.n50 VN.n0 0.189894
R3031 VDD2.n1 VDD2.t0 67.5719
R3032 VDD2.n3 VDD2.n2 65.5737
R3033 VDD2 VDD2.n7 65.5719
R3034 VDD2.n4 VDD2.t9 63.9513
R3035 VDD2.n6 VDD2.n5 62.9147
R3036 VDD2.n1 VDD2.n0 62.9135
R3037 VDD2.n4 VDD2.n3 57.3791
R3038 VDD2.n6 VDD2.n4 3.62119
R3039 VDD2.n7 VDD2.t5 1.03715
R3040 VDD2.n7 VDD2.t2 1.03715
R3041 VDD2.n5 VDD2.t3 1.03715
R3042 VDD2.n5 VDD2.t7 1.03715
R3043 VDD2.n2 VDD2.t1 1.03715
R3044 VDD2.n2 VDD2.t8 1.03715
R3045 VDD2.n0 VDD2.t6 1.03715
R3046 VDD2.n0 VDD2.t4 1.03715
R3047 VDD2 VDD2.n6 0.963862
R3048 VDD2.n3 VDD2.n1 0.850326
C0 VN VP 11.6f
C1 VN VDD1 0.155989f
C2 VTAIL VP 18.6803f
C3 VN VDD2 17.821001f
C4 VTAIL VDD1 13.7922f
C5 VTAIL VDD2 13.8516f
C6 VDD1 VP 18.405901f
C7 VN VTAIL 18.664999f
C8 VDD2 VP 0.744755f
C9 VDD1 VDD2 3.00282f
C10 VDD2 B 9.911874f
C11 VDD1 B 9.918755f
C12 VTAIL B 12.054374f
C13 VN B 24.781961f
C14 VP B 23.312342f
C15 VDD2.t0 B 4.21998f
C16 VDD2.t6 B 0.358106f
C17 VDD2.t4 B 0.358106f
C18 VDD2.n0 B 3.27757f
C19 VDD2.n1 B 1.04351f
C20 VDD2.t1 B 0.358106f
C21 VDD2.t8 B 0.358106f
C22 VDD2.n2 B 3.30516f
C23 VDD2.n3 B 3.80482f
C24 VDD2.t9 B 4.19107f
C25 VDD2.n4 B 3.94064f
C26 VDD2.t3 B 0.358106f
C27 VDD2.t7 B 0.358106f
C28 VDD2.n5 B 3.27757f
C29 VDD2.n6 B 0.540689f
C30 VDD2.t5 B 0.358106f
C31 VDD2.t2 B 0.358106f
C32 VDD2.n7 B 3.3051f
C33 VN.n0 B 0.029065f
C34 VN.t1 B 3.14406f
C35 VN.n1 B 0.028934f
C36 VN.n2 B 0.015447f
C37 VN.n3 B 0.028934f
C38 VN.n4 B 0.015447f
C39 VN.t8 B 3.14406f
C40 VN.n5 B 0.028934f
C41 VN.n6 B 0.015447f
C42 VN.n7 B 0.028934f
C43 VN.n8 B 0.015447f
C44 VN.t5 B 3.14406f
C45 VN.n9 B 0.028934f
C46 VN.n10 B 0.015447f
C47 VN.n11 B 0.028934f
C48 VN.n12 B 0.204626f
C49 VN.t3 B 3.14406f
C50 VN.t9 B 3.40007f
C51 VN.n13 B 1.08749f
C52 VN.n14 B 1.13564f
C53 VN.n15 B 0.020363f
C54 VN.n16 B 0.028934f
C55 VN.n17 B 0.015447f
C56 VN.n18 B 0.015447f
C57 VN.n19 B 0.015447f
C58 VN.n20 B 0.028493f
C59 VN.n21 B 0.014622f
C60 VN.n22 B 0.031116f
C61 VN.n23 B 0.015447f
C62 VN.n24 B 0.015447f
C63 VN.n25 B 0.015447f
C64 VN.n26 B 0.028934f
C65 VN.n27 B 1.09557f
C66 VN.n28 B 0.028934f
C67 VN.n29 B 0.015447f
C68 VN.n30 B 0.015447f
C69 VN.n31 B 0.015447f
C70 VN.n32 B 0.031116f
C71 VN.n33 B 0.014622f
C72 VN.n34 B 0.028493f
C73 VN.n35 B 0.015447f
C74 VN.n36 B 0.015447f
C75 VN.n37 B 0.015447f
C76 VN.n38 B 0.028934f
C77 VN.n39 B 0.020363f
C78 VN.n40 B 1.08092f
C79 VN.n41 B 0.02322f
C80 VN.n42 B 0.015447f
C81 VN.n43 B 0.015447f
C82 VN.n44 B 0.015447f
C83 VN.n45 B 0.028934f
C84 VN.n46 B 0.024816f
C85 VN.n47 B 0.020481f
C86 VN.n48 B 0.015447f
C87 VN.n49 B 0.015447f
C88 VN.n50 B 0.015447f
C89 VN.n51 B 0.028934f
C90 VN.n52 B 0.026077f
C91 VN.n53 B 1.14709f
C92 VN.n54 B 0.049112f
C93 VN.n55 B 0.029065f
C94 VN.t0 B 3.14406f
C95 VN.n56 B 0.028934f
C96 VN.n57 B 0.015447f
C97 VN.n58 B 0.028934f
C98 VN.n59 B 0.015447f
C99 VN.t6 B 3.14406f
C100 VN.n60 B 0.028934f
C101 VN.n61 B 0.015447f
C102 VN.n62 B 0.028934f
C103 VN.n63 B 0.015447f
C104 VN.t2 B 3.14406f
C105 VN.n64 B 0.028934f
C106 VN.n65 B 0.015447f
C107 VN.n66 B 0.028934f
C108 VN.n67 B 0.204626f
C109 VN.t4 B 3.14406f
C110 VN.t7 B 3.40007f
C111 VN.n68 B 1.08749f
C112 VN.n69 B 1.13564f
C113 VN.n70 B 0.020363f
C114 VN.n71 B 0.028934f
C115 VN.n72 B 0.015447f
C116 VN.n73 B 0.015447f
C117 VN.n74 B 0.015447f
C118 VN.n75 B 0.028493f
C119 VN.n76 B 0.014622f
C120 VN.n77 B 0.031116f
C121 VN.n78 B 0.015447f
C122 VN.n79 B 0.015447f
C123 VN.n80 B 0.015447f
C124 VN.n81 B 0.028934f
C125 VN.n82 B 1.09557f
C126 VN.n83 B 0.028934f
C127 VN.n84 B 0.015447f
C128 VN.n85 B 0.015447f
C129 VN.n86 B 0.015447f
C130 VN.n87 B 0.031116f
C131 VN.n88 B 0.014622f
C132 VN.n89 B 0.028493f
C133 VN.n90 B 0.015447f
C134 VN.n91 B 0.015447f
C135 VN.n92 B 0.015447f
C136 VN.n93 B 0.028934f
C137 VN.n94 B 0.020363f
C138 VN.n95 B 1.08092f
C139 VN.n96 B 0.02322f
C140 VN.n97 B 0.015447f
C141 VN.n98 B 0.015447f
C142 VN.n99 B 0.015447f
C143 VN.n100 B 0.028934f
C144 VN.n101 B 0.024816f
C145 VN.n102 B 0.020481f
C146 VN.n103 B 0.015447f
C147 VN.n104 B 0.015447f
C148 VN.n105 B 0.015447f
C149 VN.n106 B 0.028934f
C150 VN.n107 B 0.026077f
C151 VN.n108 B 1.14709f
C152 VN.n109 B 1.29526f
C153 VTAIL.t7 B 0.364407f
C154 VTAIL.t3 B 0.364407f
C155 VTAIL.n0 B 3.26706f
C156 VTAIL.n1 B 0.622121f
C157 VTAIL.t10 B 4.17543f
C158 VTAIL.n2 B 0.773477f
C159 VTAIL.t13 B 0.364407f
C160 VTAIL.t18 B 0.364407f
C161 VTAIL.n3 B 3.26706f
C162 VTAIL.n4 B 0.792299f
C163 VTAIL.t16 B 0.364407f
C164 VTAIL.t11 B 0.364407f
C165 VTAIL.n5 B 3.26706f
C166 VTAIL.n6 B 2.68288f
C167 VTAIL.t6 B 0.364407f
C168 VTAIL.t0 B 0.364407f
C169 VTAIL.n7 B 3.26707f
C170 VTAIL.n8 B 2.68287f
C171 VTAIL.t4 B 0.364407f
C172 VTAIL.t9 B 0.364407f
C173 VTAIL.n9 B 3.26707f
C174 VTAIL.n10 B 0.79229f
C175 VTAIL.t2 B 4.17546f
C176 VTAIL.n11 B 0.773446f
C177 VTAIL.t12 B 0.364407f
C178 VTAIL.t17 B 0.364407f
C179 VTAIL.n12 B 3.26707f
C180 VTAIL.n13 B 0.688003f
C181 VTAIL.t14 B 0.364407f
C182 VTAIL.t19 B 0.364407f
C183 VTAIL.n14 B 3.26707f
C184 VTAIL.n15 B 0.79229f
C185 VTAIL.t15 B 4.17543f
C186 VTAIL.n16 B 2.48667f
C187 VTAIL.t5 B 4.17543f
C188 VTAIL.n17 B 2.48667f
C189 VTAIL.t1 B 0.364407f
C190 VTAIL.t8 B 0.364407f
C191 VTAIL.n18 B 3.26706f
C192 VTAIL.n19 B 0.576517f
C193 VDD1.t6 B 4.27002f
C194 VDD1.t3 B 0.362351f
C195 VDD1.t8 B 0.362351f
C196 VDD1.n0 B 3.31643f
C197 VDD1.n1 B 1.06398f
C198 VDD1.t2 B 4.27f
C199 VDD1.t1 B 0.362351f
C200 VDD1.t7 B 0.362351f
C201 VDD1.n2 B 3.31642f
C202 VDD1.n3 B 1.05588f
C203 VDD1.t4 B 0.362351f
C204 VDD1.t0 B 0.362351f
C205 VDD1.n4 B 3.34434f
C206 VDD1.n5 B 4.00851f
C207 VDD1.t5 B 0.362351f
C208 VDD1.t9 B 0.362351f
C209 VDD1.n6 B 3.31641f
C210 VDD1.n7 B 4.05912f
C211 VP.n0 B 0.02944f
C212 VP.t9 B 3.18472f
C213 VP.n1 B 0.029308f
C214 VP.n2 B 0.015647f
C215 VP.n3 B 0.029308f
C216 VP.n4 B 0.015647f
C217 VP.t1 B 3.18472f
C218 VP.n5 B 0.029308f
C219 VP.n6 B 0.015647f
C220 VP.n7 B 0.029308f
C221 VP.n8 B 0.015647f
C222 VP.t6 B 3.18472f
C223 VP.n9 B 0.029308f
C224 VP.n10 B 0.015647f
C225 VP.n11 B 0.029308f
C226 VP.n12 B 0.015647f
C227 VP.t8 B 3.18472f
C228 VP.n13 B 0.029308f
C229 VP.n14 B 0.015647f
C230 VP.n15 B 0.029308f
C231 VP.n16 B 0.02944f
C232 VP.t3 B 3.18472f
C233 VP.n17 B 0.02944f
C234 VP.t4 B 3.18472f
C235 VP.n18 B 0.029308f
C236 VP.n19 B 0.015647f
C237 VP.n20 B 0.029308f
C238 VP.n21 B 0.015647f
C239 VP.t0 B 3.18472f
C240 VP.n22 B 0.029308f
C241 VP.n23 B 0.015647f
C242 VP.n24 B 0.029308f
C243 VP.n25 B 0.015647f
C244 VP.t5 B 3.18472f
C245 VP.n26 B 0.029308f
C246 VP.n27 B 0.015647f
C247 VP.n28 B 0.029308f
C248 VP.n29 B 0.207273f
C249 VP.t2 B 3.18472f
C250 VP.t7 B 3.44404f
C251 VP.n30 B 1.10156f
C252 VP.n31 B 1.15032f
C253 VP.n32 B 0.020626f
C254 VP.n33 B 0.029308f
C255 VP.n34 B 0.015647f
C256 VP.n35 B 0.015647f
C257 VP.n36 B 0.015647f
C258 VP.n37 B 0.028862f
C259 VP.n38 B 0.014811f
C260 VP.n39 B 0.031518f
C261 VP.n40 B 0.015647f
C262 VP.n41 B 0.015647f
C263 VP.n42 B 0.015647f
C264 VP.n43 B 0.029308f
C265 VP.n44 B 1.10974f
C266 VP.n45 B 0.029308f
C267 VP.n46 B 0.015647f
C268 VP.n47 B 0.015647f
C269 VP.n48 B 0.015647f
C270 VP.n49 B 0.031518f
C271 VP.n50 B 0.014811f
C272 VP.n51 B 0.028862f
C273 VP.n52 B 0.015647f
C274 VP.n53 B 0.015647f
C275 VP.n54 B 0.015647f
C276 VP.n55 B 0.029308f
C277 VP.n56 B 0.020626f
C278 VP.n57 B 1.0949f
C279 VP.n58 B 0.02352f
C280 VP.n59 B 0.015647f
C281 VP.n60 B 0.015647f
C282 VP.n61 B 0.015647f
C283 VP.n62 B 0.029308f
C284 VP.n63 B 0.025137f
C285 VP.n64 B 0.020746f
C286 VP.n65 B 0.015647f
C287 VP.n66 B 0.015647f
C288 VP.n67 B 0.015647f
C289 VP.n68 B 0.029308f
C290 VP.n69 B 0.026414f
C291 VP.n70 B 1.16192f
C292 VP.n71 B 1.30864f
C293 VP.n72 B 1.31719f
C294 VP.n73 B 1.16192f
C295 VP.n74 B 0.026414f
C296 VP.n75 B 0.029308f
C297 VP.n76 B 0.015647f
C298 VP.n77 B 0.015647f
C299 VP.n78 B 0.015647f
C300 VP.n79 B 0.020746f
C301 VP.n80 B 0.025137f
C302 VP.n81 B 0.029308f
C303 VP.n82 B 0.015647f
C304 VP.n83 B 0.015647f
C305 VP.n84 B 0.015647f
C306 VP.n85 B 0.02352f
C307 VP.n86 B 1.0949f
C308 VP.n87 B 0.020626f
C309 VP.n88 B 0.029308f
C310 VP.n89 B 0.015647f
C311 VP.n90 B 0.015647f
C312 VP.n91 B 0.015647f
C313 VP.n92 B 0.028862f
C314 VP.n93 B 0.014811f
C315 VP.n94 B 0.031518f
C316 VP.n95 B 0.015647f
C317 VP.n96 B 0.015647f
C318 VP.n97 B 0.015647f
C319 VP.n98 B 0.029308f
C320 VP.n99 B 1.10974f
C321 VP.n100 B 0.029308f
C322 VP.n101 B 0.015647f
C323 VP.n102 B 0.015647f
C324 VP.n103 B 0.015647f
C325 VP.n104 B 0.031518f
C326 VP.n105 B 0.014811f
C327 VP.n106 B 0.028862f
C328 VP.n107 B 0.015647f
C329 VP.n108 B 0.015647f
C330 VP.n109 B 0.015647f
C331 VP.n110 B 0.029308f
C332 VP.n111 B 0.020626f
C333 VP.n112 B 1.0949f
C334 VP.n113 B 0.02352f
C335 VP.n114 B 0.015647f
C336 VP.n115 B 0.015647f
C337 VP.n116 B 0.015647f
C338 VP.n117 B 0.029308f
C339 VP.n118 B 0.025137f
C340 VP.n119 B 0.020746f
C341 VP.n120 B 0.015647f
C342 VP.n121 B 0.015647f
C343 VP.n122 B 0.015647f
C344 VP.n123 B 0.029308f
C345 VP.n124 B 0.026414f
C346 VP.n125 B 1.16192f
C347 VP.n126 B 0.049747f
.ends

