* NGSPICE file created from diff_pair_sample_1111.ext - technology: sky130A

.subckt diff_pair_sample_1111 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 w_n2062_n4022# sky130_fd_pr__pfet_01v8 ad=5.9553 pd=31.32 as=5.9553 ps=31.32 w=15.27 l=2.4
X1 VDD1.t1 VP.t0 VTAIL.t0 w_n2062_n4022# sky130_fd_pr__pfet_01v8 ad=5.9553 pd=31.32 as=5.9553 ps=31.32 w=15.27 l=2.4
X2 B.t11 B.t9 B.t10 w_n2062_n4022# sky130_fd_pr__pfet_01v8 ad=5.9553 pd=31.32 as=0 ps=0 w=15.27 l=2.4
X3 VDD2.t0 VN.t1 VTAIL.t3 w_n2062_n4022# sky130_fd_pr__pfet_01v8 ad=5.9553 pd=31.32 as=5.9553 ps=31.32 w=15.27 l=2.4
X4 B.t8 B.t6 B.t7 w_n2062_n4022# sky130_fd_pr__pfet_01v8 ad=5.9553 pd=31.32 as=0 ps=0 w=15.27 l=2.4
X5 B.t5 B.t3 B.t4 w_n2062_n4022# sky130_fd_pr__pfet_01v8 ad=5.9553 pd=31.32 as=0 ps=0 w=15.27 l=2.4
X6 VDD1.t0 VP.t1 VTAIL.t1 w_n2062_n4022# sky130_fd_pr__pfet_01v8 ad=5.9553 pd=31.32 as=5.9553 ps=31.32 w=15.27 l=2.4
X7 B.t2 B.t0 B.t1 w_n2062_n4022# sky130_fd_pr__pfet_01v8 ad=5.9553 pd=31.32 as=0 ps=0 w=15.27 l=2.4
R0 VN VN.t1 249.207
R1 VN VN.t0 202.844
R2 VTAIL.n2 VTAIL.t0 54.4945
R3 VTAIL.n1 VTAIL.t3 54.4945
R4 VTAIL.n3 VTAIL.t2 54.4944
R5 VTAIL.n0 VTAIL.t1 54.4944
R6 VTAIL.n1 VTAIL.n0 30.2376
R7 VTAIL.n3 VTAIL.n2 27.8841
R8 VTAIL.n2 VTAIL.n1 1.64705
R9 VTAIL VTAIL.n0 1.11688
R10 VTAIL VTAIL.n3 0.530672
R11 VDD2.n0 VDD2.t1 112.704
R12 VDD2.n0 VDD2.t0 71.1733
R13 VDD2 VDD2.n0 0.647052
R14 VP.n0 VP.t0 249.111
R15 VP.n0 VP.t1 202.507
R16 VP VP.n0 0.336784
R17 VDD1 VDD1.t0 113.817
R18 VDD1 VDD1.t1 71.8199
R19 B.n450 B.n449 585
R20 B.n451 B.n74 585
R21 B.n453 B.n452 585
R22 B.n454 B.n73 585
R23 B.n456 B.n455 585
R24 B.n457 B.n72 585
R25 B.n459 B.n458 585
R26 B.n460 B.n71 585
R27 B.n462 B.n461 585
R28 B.n463 B.n70 585
R29 B.n465 B.n464 585
R30 B.n466 B.n69 585
R31 B.n468 B.n467 585
R32 B.n469 B.n68 585
R33 B.n471 B.n470 585
R34 B.n472 B.n67 585
R35 B.n474 B.n473 585
R36 B.n475 B.n66 585
R37 B.n477 B.n476 585
R38 B.n478 B.n65 585
R39 B.n480 B.n479 585
R40 B.n481 B.n64 585
R41 B.n483 B.n482 585
R42 B.n484 B.n63 585
R43 B.n486 B.n485 585
R44 B.n487 B.n62 585
R45 B.n489 B.n488 585
R46 B.n490 B.n61 585
R47 B.n492 B.n491 585
R48 B.n493 B.n60 585
R49 B.n495 B.n494 585
R50 B.n496 B.n59 585
R51 B.n498 B.n497 585
R52 B.n499 B.n58 585
R53 B.n501 B.n500 585
R54 B.n502 B.n57 585
R55 B.n504 B.n503 585
R56 B.n505 B.n56 585
R57 B.n507 B.n506 585
R58 B.n508 B.n55 585
R59 B.n510 B.n509 585
R60 B.n511 B.n54 585
R61 B.n513 B.n512 585
R62 B.n514 B.n53 585
R63 B.n516 B.n515 585
R64 B.n517 B.n52 585
R65 B.n519 B.n518 585
R66 B.n520 B.n51 585
R67 B.n522 B.n521 585
R68 B.n523 B.n47 585
R69 B.n525 B.n524 585
R70 B.n526 B.n46 585
R71 B.n528 B.n527 585
R72 B.n529 B.n45 585
R73 B.n531 B.n530 585
R74 B.n532 B.n44 585
R75 B.n534 B.n533 585
R76 B.n535 B.n43 585
R77 B.n537 B.n536 585
R78 B.n538 B.n42 585
R79 B.n540 B.n539 585
R80 B.n542 B.n39 585
R81 B.n544 B.n543 585
R82 B.n545 B.n38 585
R83 B.n547 B.n546 585
R84 B.n548 B.n37 585
R85 B.n550 B.n549 585
R86 B.n551 B.n36 585
R87 B.n553 B.n552 585
R88 B.n554 B.n35 585
R89 B.n556 B.n555 585
R90 B.n557 B.n34 585
R91 B.n559 B.n558 585
R92 B.n560 B.n33 585
R93 B.n562 B.n561 585
R94 B.n563 B.n32 585
R95 B.n565 B.n564 585
R96 B.n566 B.n31 585
R97 B.n568 B.n567 585
R98 B.n569 B.n30 585
R99 B.n571 B.n570 585
R100 B.n572 B.n29 585
R101 B.n574 B.n573 585
R102 B.n575 B.n28 585
R103 B.n577 B.n576 585
R104 B.n578 B.n27 585
R105 B.n580 B.n579 585
R106 B.n581 B.n26 585
R107 B.n583 B.n582 585
R108 B.n584 B.n25 585
R109 B.n586 B.n585 585
R110 B.n587 B.n24 585
R111 B.n589 B.n588 585
R112 B.n590 B.n23 585
R113 B.n592 B.n591 585
R114 B.n593 B.n22 585
R115 B.n595 B.n594 585
R116 B.n596 B.n21 585
R117 B.n598 B.n597 585
R118 B.n599 B.n20 585
R119 B.n601 B.n600 585
R120 B.n602 B.n19 585
R121 B.n604 B.n603 585
R122 B.n605 B.n18 585
R123 B.n607 B.n606 585
R124 B.n608 B.n17 585
R125 B.n610 B.n609 585
R126 B.n611 B.n16 585
R127 B.n613 B.n612 585
R128 B.n614 B.n15 585
R129 B.n616 B.n615 585
R130 B.n617 B.n14 585
R131 B.n448 B.n75 585
R132 B.n447 B.n446 585
R133 B.n445 B.n76 585
R134 B.n444 B.n443 585
R135 B.n442 B.n77 585
R136 B.n441 B.n440 585
R137 B.n439 B.n78 585
R138 B.n438 B.n437 585
R139 B.n436 B.n79 585
R140 B.n435 B.n434 585
R141 B.n433 B.n80 585
R142 B.n432 B.n431 585
R143 B.n430 B.n81 585
R144 B.n429 B.n428 585
R145 B.n427 B.n82 585
R146 B.n426 B.n425 585
R147 B.n424 B.n83 585
R148 B.n423 B.n422 585
R149 B.n421 B.n84 585
R150 B.n420 B.n419 585
R151 B.n418 B.n85 585
R152 B.n417 B.n416 585
R153 B.n415 B.n86 585
R154 B.n414 B.n413 585
R155 B.n412 B.n87 585
R156 B.n411 B.n410 585
R157 B.n409 B.n88 585
R158 B.n408 B.n407 585
R159 B.n406 B.n89 585
R160 B.n405 B.n404 585
R161 B.n403 B.n90 585
R162 B.n402 B.n401 585
R163 B.n400 B.n91 585
R164 B.n399 B.n398 585
R165 B.n397 B.n92 585
R166 B.n396 B.n395 585
R167 B.n394 B.n93 585
R168 B.n393 B.n392 585
R169 B.n391 B.n94 585
R170 B.n390 B.n389 585
R171 B.n388 B.n95 585
R172 B.n387 B.n386 585
R173 B.n385 B.n96 585
R174 B.n384 B.n383 585
R175 B.n382 B.n97 585
R176 B.n381 B.n380 585
R177 B.n379 B.n98 585
R178 B.n378 B.n377 585
R179 B.n376 B.n99 585
R180 B.n207 B.n206 585
R181 B.n208 B.n159 585
R182 B.n210 B.n209 585
R183 B.n211 B.n158 585
R184 B.n213 B.n212 585
R185 B.n214 B.n157 585
R186 B.n216 B.n215 585
R187 B.n217 B.n156 585
R188 B.n219 B.n218 585
R189 B.n220 B.n155 585
R190 B.n222 B.n221 585
R191 B.n223 B.n154 585
R192 B.n225 B.n224 585
R193 B.n226 B.n153 585
R194 B.n228 B.n227 585
R195 B.n229 B.n152 585
R196 B.n231 B.n230 585
R197 B.n232 B.n151 585
R198 B.n234 B.n233 585
R199 B.n235 B.n150 585
R200 B.n237 B.n236 585
R201 B.n238 B.n149 585
R202 B.n240 B.n239 585
R203 B.n241 B.n148 585
R204 B.n243 B.n242 585
R205 B.n244 B.n147 585
R206 B.n246 B.n245 585
R207 B.n247 B.n146 585
R208 B.n249 B.n248 585
R209 B.n250 B.n145 585
R210 B.n252 B.n251 585
R211 B.n253 B.n144 585
R212 B.n255 B.n254 585
R213 B.n256 B.n143 585
R214 B.n258 B.n257 585
R215 B.n259 B.n142 585
R216 B.n261 B.n260 585
R217 B.n262 B.n141 585
R218 B.n264 B.n263 585
R219 B.n265 B.n140 585
R220 B.n267 B.n266 585
R221 B.n268 B.n139 585
R222 B.n270 B.n269 585
R223 B.n271 B.n138 585
R224 B.n273 B.n272 585
R225 B.n274 B.n137 585
R226 B.n276 B.n275 585
R227 B.n277 B.n136 585
R228 B.n279 B.n278 585
R229 B.n280 B.n135 585
R230 B.n282 B.n281 585
R231 B.n284 B.n132 585
R232 B.n286 B.n285 585
R233 B.n287 B.n131 585
R234 B.n289 B.n288 585
R235 B.n290 B.n130 585
R236 B.n292 B.n291 585
R237 B.n293 B.n129 585
R238 B.n295 B.n294 585
R239 B.n296 B.n128 585
R240 B.n298 B.n297 585
R241 B.n300 B.n299 585
R242 B.n301 B.n124 585
R243 B.n303 B.n302 585
R244 B.n304 B.n123 585
R245 B.n306 B.n305 585
R246 B.n307 B.n122 585
R247 B.n309 B.n308 585
R248 B.n310 B.n121 585
R249 B.n312 B.n311 585
R250 B.n313 B.n120 585
R251 B.n315 B.n314 585
R252 B.n316 B.n119 585
R253 B.n318 B.n317 585
R254 B.n319 B.n118 585
R255 B.n321 B.n320 585
R256 B.n322 B.n117 585
R257 B.n324 B.n323 585
R258 B.n325 B.n116 585
R259 B.n327 B.n326 585
R260 B.n328 B.n115 585
R261 B.n330 B.n329 585
R262 B.n331 B.n114 585
R263 B.n333 B.n332 585
R264 B.n334 B.n113 585
R265 B.n336 B.n335 585
R266 B.n337 B.n112 585
R267 B.n339 B.n338 585
R268 B.n340 B.n111 585
R269 B.n342 B.n341 585
R270 B.n343 B.n110 585
R271 B.n345 B.n344 585
R272 B.n346 B.n109 585
R273 B.n348 B.n347 585
R274 B.n349 B.n108 585
R275 B.n351 B.n350 585
R276 B.n352 B.n107 585
R277 B.n354 B.n353 585
R278 B.n355 B.n106 585
R279 B.n357 B.n356 585
R280 B.n358 B.n105 585
R281 B.n360 B.n359 585
R282 B.n361 B.n104 585
R283 B.n363 B.n362 585
R284 B.n364 B.n103 585
R285 B.n366 B.n365 585
R286 B.n367 B.n102 585
R287 B.n369 B.n368 585
R288 B.n370 B.n101 585
R289 B.n372 B.n371 585
R290 B.n373 B.n100 585
R291 B.n375 B.n374 585
R292 B.n205 B.n160 585
R293 B.n204 B.n203 585
R294 B.n202 B.n161 585
R295 B.n201 B.n200 585
R296 B.n199 B.n162 585
R297 B.n198 B.n197 585
R298 B.n196 B.n163 585
R299 B.n195 B.n194 585
R300 B.n193 B.n164 585
R301 B.n192 B.n191 585
R302 B.n190 B.n165 585
R303 B.n189 B.n188 585
R304 B.n187 B.n166 585
R305 B.n186 B.n185 585
R306 B.n184 B.n167 585
R307 B.n183 B.n182 585
R308 B.n181 B.n168 585
R309 B.n180 B.n179 585
R310 B.n178 B.n169 585
R311 B.n177 B.n176 585
R312 B.n175 B.n170 585
R313 B.n174 B.n173 585
R314 B.n172 B.n171 585
R315 B.n2 B.n0 585
R316 B.n653 B.n1 585
R317 B.n652 B.n651 585
R318 B.n650 B.n3 585
R319 B.n649 B.n648 585
R320 B.n647 B.n4 585
R321 B.n646 B.n645 585
R322 B.n644 B.n5 585
R323 B.n643 B.n642 585
R324 B.n641 B.n6 585
R325 B.n640 B.n639 585
R326 B.n638 B.n7 585
R327 B.n637 B.n636 585
R328 B.n635 B.n8 585
R329 B.n634 B.n633 585
R330 B.n632 B.n9 585
R331 B.n631 B.n630 585
R332 B.n629 B.n10 585
R333 B.n628 B.n627 585
R334 B.n626 B.n11 585
R335 B.n625 B.n624 585
R336 B.n623 B.n12 585
R337 B.n622 B.n621 585
R338 B.n620 B.n13 585
R339 B.n619 B.n618 585
R340 B.n655 B.n654 585
R341 B.n207 B.n160 530.939
R342 B.n618 B.n617 530.939
R343 B.n376 B.n375 530.939
R344 B.n449 B.n448 530.939
R345 B.n125 B.t0 361.06
R346 B.n133 B.t6 361.06
R347 B.n40 B.t9 361.06
R348 B.n48 B.t3 361.06
R349 B.n125 B.t2 165.481
R350 B.n48 B.t4 165.481
R351 B.n133 B.t8 165.462
R352 B.n40 B.t10 165.462
R353 B.n203 B.n160 163.367
R354 B.n203 B.n202 163.367
R355 B.n202 B.n201 163.367
R356 B.n201 B.n162 163.367
R357 B.n197 B.n162 163.367
R358 B.n197 B.n196 163.367
R359 B.n196 B.n195 163.367
R360 B.n195 B.n164 163.367
R361 B.n191 B.n164 163.367
R362 B.n191 B.n190 163.367
R363 B.n190 B.n189 163.367
R364 B.n189 B.n166 163.367
R365 B.n185 B.n166 163.367
R366 B.n185 B.n184 163.367
R367 B.n184 B.n183 163.367
R368 B.n183 B.n168 163.367
R369 B.n179 B.n168 163.367
R370 B.n179 B.n178 163.367
R371 B.n178 B.n177 163.367
R372 B.n177 B.n170 163.367
R373 B.n173 B.n170 163.367
R374 B.n173 B.n172 163.367
R375 B.n172 B.n2 163.367
R376 B.n654 B.n2 163.367
R377 B.n654 B.n653 163.367
R378 B.n653 B.n652 163.367
R379 B.n652 B.n3 163.367
R380 B.n648 B.n3 163.367
R381 B.n648 B.n647 163.367
R382 B.n647 B.n646 163.367
R383 B.n646 B.n5 163.367
R384 B.n642 B.n5 163.367
R385 B.n642 B.n641 163.367
R386 B.n641 B.n640 163.367
R387 B.n640 B.n7 163.367
R388 B.n636 B.n7 163.367
R389 B.n636 B.n635 163.367
R390 B.n635 B.n634 163.367
R391 B.n634 B.n9 163.367
R392 B.n630 B.n9 163.367
R393 B.n630 B.n629 163.367
R394 B.n629 B.n628 163.367
R395 B.n628 B.n11 163.367
R396 B.n624 B.n11 163.367
R397 B.n624 B.n623 163.367
R398 B.n623 B.n622 163.367
R399 B.n622 B.n13 163.367
R400 B.n618 B.n13 163.367
R401 B.n208 B.n207 163.367
R402 B.n209 B.n208 163.367
R403 B.n209 B.n158 163.367
R404 B.n213 B.n158 163.367
R405 B.n214 B.n213 163.367
R406 B.n215 B.n214 163.367
R407 B.n215 B.n156 163.367
R408 B.n219 B.n156 163.367
R409 B.n220 B.n219 163.367
R410 B.n221 B.n220 163.367
R411 B.n221 B.n154 163.367
R412 B.n225 B.n154 163.367
R413 B.n226 B.n225 163.367
R414 B.n227 B.n226 163.367
R415 B.n227 B.n152 163.367
R416 B.n231 B.n152 163.367
R417 B.n232 B.n231 163.367
R418 B.n233 B.n232 163.367
R419 B.n233 B.n150 163.367
R420 B.n237 B.n150 163.367
R421 B.n238 B.n237 163.367
R422 B.n239 B.n238 163.367
R423 B.n239 B.n148 163.367
R424 B.n243 B.n148 163.367
R425 B.n244 B.n243 163.367
R426 B.n245 B.n244 163.367
R427 B.n245 B.n146 163.367
R428 B.n249 B.n146 163.367
R429 B.n250 B.n249 163.367
R430 B.n251 B.n250 163.367
R431 B.n251 B.n144 163.367
R432 B.n255 B.n144 163.367
R433 B.n256 B.n255 163.367
R434 B.n257 B.n256 163.367
R435 B.n257 B.n142 163.367
R436 B.n261 B.n142 163.367
R437 B.n262 B.n261 163.367
R438 B.n263 B.n262 163.367
R439 B.n263 B.n140 163.367
R440 B.n267 B.n140 163.367
R441 B.n268 B.n267 163.367
R442 B.n269 B.n268 163.367
R443 B.n269 B.n138 163.367
R444 B.n273 B.n138 163.367
R445 B.n274 B.n273 163.367
R446 B.n275 B.n274 163.367
R447 B.n275 B.n136 163.367
R448 B.n279 B.n136 163.367
R449 B.n280 B.n279 163.367
R450 B.n281 B.n280 163.367
R451 B.n281 B.n132 163.367
R452 B.n286 B.n132 163.367
R453 B.n287 B.n286 163.367
R454 B.n288 B.n287 163.367
R455 B.n288 B.n130 163.367
R456 B.n292 B.n130 163.367
R457 B.n293 B.n292 163.367
R458 B.n294 B.n293 163.367
R459 B.n294 B.n128 163.367
R460 B.n298 B.n128 163.367
R461 B.n299 B.n298 163.367
R462 B.n299 B.n124 163.367
R463 B.n303 B.n124 163.367
R464 B.n304 B.n303 163.367
R465 B.n305 B.n304 163.367
R466 B.n305 B.n122 163.367
R467 B.n309 B.n122 163.367
R468 B.n310 B.n309 163.367
R469 B.n311 B.n310 163.367
R470 B.n311 B.n120 163.367
R471 B.n315 B.n120 163.367
R472 B.n316 B.n315 163.367
R473 B.n317 B.n316 163.367
R474 B.n317 B.n118 163.367
R475 B.n321 B.n118 163.367
R476 B.n322 B.n321 163.367
R477 B.n323 B.n322 163.367
R478 B.n323 B.n116 163.367
R479 B.n327 B.n116 163.367
R480 B.n328 B.n327 163.367
R481 B.n329 B.n328 163.367
R482 B.n329 B.n114 163.367
R483 B.n333 B.n114 163.367
R484 B.n334 B.n333 163.367
R485 B.n335 B.n334 163.367
R486 B.n335 B.n112 163.367
R487 B.n339 B.n112 163.367
R488 B.n340 B.n339 163.367
R489 B.n341 B.n340 163.367
R490 B.n341 B.n110 163.367
R491 B.n345 B.n110 163.367
R492 B.n346 B.n345 163.367
R493 B.n347 B.n346 163.367
R494 B.n347 B.n108 163.367
R495 B.n351 B.n108 163.367
R496 B.n352 B.n351 163.367
R497 B.n353 B.n352 163.367
R498 B.n353 B.n106 163.367
R499 B.n357 B.n106 163.367
R500 B.n358 B.n357 163.367
R501 B.n359 B.n358 163.367
R502 B.n359 B.n104 163.367
R503 B.n363 B.n104 163.367
R504 B.n364 B.n363 163.367
R505 B.n365 B.n364 163.367
R506 B.n365 B.n102 163.367
R507 B.n369 B.n102 163.367
R508 B.n370 B.n369 163.367
R509 B.n371 B.n370 163.367
R510 B.n371 B.n100 163.367
R511 B.n375 B.n100 163.367
R512 B.n377 B.n376 163.367
R513 B.n377 B.n98 163.367
R514 B.n381 B.n98 163.367
R515 B.n382 B.n381 163.367
R516 B.n383 B.n382 163.367
R517 B.n383 B.n96 163.367
R518 B.n387 B.n96 163.367
R519 B.n388 B.n387 163.367
R520 B.n389 B.n388 163.367
R521 B.n389 B.n94 163.367
R522 B.n393 B.n94 163.367
R523 B.n394 B.n393 163.367
R524 B.n395 B.n394 163.367
R525 B.n395 B.n92 163.367
R526 B.n399 B.n92 163.367
R527 B.n400 B.n399 163.367
R528 B.n401 B.n400 163.367
R529 B.n401 B.n90 163.367
R530 B.n405 B.n90 163.367
R531 B.n406 B.n405 163.367
R532 B.n407 B.n406 163.367
R533 B.n407 B.n88 163.367
R534 B.n411 B.n88 163.367
R535 B.n412 B.n411 163.367
R536 B.n413 B.n412 163.367
R537 B.n413 B.n86 163.367
R538 B.n417 B.n86 163.367
R539 B.n418 B.n417 163.367
R540 B.n419 B.n418 163.367
R541 B.n419 B.n84 163.367
R542 B.n423 B.n84 163.367
R543 B.n424 B.n423 163.367
R544 B.n425 B.n424 163.367
R545 B.n425 B.n82 163.367
R546 B.n429 B.n82 163.367
R547 B.n430 B.n429 163.367
R548 B.n431 B.n430 163.367
R549 B.n431 B.n80 163.367
R550 B.n435 B.n80 163.367
R551 B.n436 B.n435 163.367
R552 B.n437 B.n436 163.367
R553 B.n437 B.n78 163.367
R554 B.n441 B.n78 163.367
R555 B.n442 B.n441 163.367
R556 B.n443 B.n442 163.367
R557 B.n443 B.n76 163.367
R558 B.n447 B.n76 163.367
R559 B.n448 B.n447 163.367
R560 B.n617 B.n616 163.367
R561 B.n616 B.n15 163.367
R562 B.n612 B.n15 163.367
R563 B.n612 B.n611 163.367
R564 B.n611 B.n610 163.367
R565 B.n610 B.n17 163.367
R566 B.n606 B.n17 163.367
R567 B.n606 B.n605 163.367
R568 B.n605 B.n604 163.367
R569 B.n604 B.n19 163.367
R570 B.n600 B.n19 163.367
R571 B.n600 B.n599 163.367
R572 B.n599 B.n598 163.367
R573 B.n598 B.n21 163.367
R574 B.n594 B.n21 163.367
R575 B.n594 B.n593 163.367
R576 B.n593 B.n592 163.367
R577 B.n592 B.n23 163.367
R578 B.n588 B.n23 163.367
R579 B.n588 B.n587 163.367
R580 B.n587 B.n586 163.367
R581 B.n586 B.n25 163.367
R582 B.n582 B.n25 163.367
R583 B.n582 B.n581 163.367
R584 B.n581 B.n580 163.367
R585 B.n580 B.n27 163.367
R586 B.n576 B.n27 163.367
R587 B.n576 B.n575 163.367
R588 B.n575 B.n574 163.367
R589 B.n574 B.n29 163.367
R590 B.n570 B.n29 163.367
R591 B.n570 B.n569 163.367
R592 B.n569 B.n568 163.367
R593 B.n568 B.n31 163.367
R594 B.n564 B.n31 163.367
R595 B.n564 B.n563 163.367
R596 B.n563 B.n562 163.367
R597 B.n562 B.n33 163.367
R598 B.n558 B.n33 163.367
R599 B.n558 B.n557 163.367
R600 B.n557 B.n556 163.367
R601 B.n556 B.n35 163.367
R602 B.n552 B.n35 163.367
R603 B.n552 B.n551 163.367
R604 B.n551 B.n550 163.367
R605 B.n550 B.n37 163.367
R606 B.n546 B.n37 163.367
R607 B.n546 B.n545 163.367
R608 B.n545 B.n544 163.367
R609 B.n544 B.n39 163.367
R610 B.n539 B.n39 163.367
R611 B.n539 B.n538 163.367
R612 B.n538 B.n537 163.367
R613 B.n537 B.n43 163.367
R614 B.n533 B.n43 163.367
R615 B.n533 B.n532 163.367
R616 B.n532 B.n531 163.367
R617 B.n531 B.n45 163.367
R618 B.n527 B.n45 163.367
R619 B.n527 B.n526 163.367
R620 B.n526 B.n525 163.367
R621 B.n525 B.n47 163.367
R622 B.n521 B.n47 163.367
R623 B.n521 B.n520 163.367
R624 B.n520 B.n519 163.367
R625 B.n519 B.n52 163.367
R626 B.n515 B.n52 163.367
R627 B.n515 B.n514 163.367
R628 B.n514 B.n513 163.367
R629 B.n513 B.n54 163.367
R630 B.n509 B.n54 163.367
R631 B.n509 B.n508 163.367
R632 B.n508 B.n507 163.367
R633 B.n507 B.n56 163.367
R634 B.n503 B.n56 163.367
R635 B.n503 B.n502 163.367
R636 B.n502 B.n501 163.367
R637 B.n501 B.n58 163.367
R638 B.n497 B.n58 163.367
R639 B.n497 B.n496 163.367
R640 B.n496 B.n495 163.367
R641 B.n495 B.n60 163.367
R642 B.n491 B.n60 163.367
R643 B.n491 B.n490 163.367
R644 B.n490 B.n489 163.367
R645 B.n489 B.n62 163.367
R646 B.n485 B.n62 163.367
R647 B.n485 B.n484 163.367
R648 B.n484 B.n483 163.367
R649 B.n483 B.n64 163.367
R650 B.n479 B.n64 163.367
R651 B.n479 B.n478 163.367
R652 B.n478 B.n477 163.367
R653 B.n477 B.n66 163.367
R654 B.n473 B.n66 163.367
R655 B.n473 B.n472 163.367
R656 B.n472 B.n471 163.367
R657 B.n471 B.n68 163.367
R658 B.n467 B.n68 163.367
R659 B.n467 B.n466 163.367
R660 B.n466 B.n465 163.367
R661 B.n465 B.n70 163.367
R662 B.n461 B.n70 163.367
R663 B.n461 B.n460 163.367
R664 B.n460 B.n459 163.367
R665 B.n459 B.n72 163.367
R666 B.n455 B.n72 163.367
R667 B.n455 B.n454 163.367
R668 B.n454 B.n453 163.367
R669 B.n453 B.n74 163.367
R670 B.n449 B.n74 163.367
R671 B.n126 B.t1 112.535
R672 B.n49 B.t5 112.535
R673 B.n134 B.t7 112.516
R674 B.n41 B.t11 112.516
R675 B.n127 B.n126 59.5399
R676 B.n283 B.n134 59.5399
R677 B.n541 B.n41 59.5399
R678 B.n50 B.n49 59.5399
R679 B.n126 B.n125 52.946
R680 B.n134 B.n133 52.946
R681 B.n41 B.n40 52.946
R682 B.n49 B.n48 52.946
R683 B.n619 B.n14 34.4981
R684 B.n450 B.n75 34.4981
R685 B.n374 B.n99 34.4981
R686 B.n206 B.n205 34.4981
R687 B B.n655 18.0485
R688 B.n615 B.n14 10.6151
R689 B.n615 B.n614 10.6151
R690 B.n614 B.n613 10.6151
R691 B.n613 B.n16 10.6151
R692 B.n609 B.n16 10.6151
R693 B.n609 B.n608 10.6151
R694 B.n608 B.n607 10.6151
R695 B.n607 B.n18 10.6151
R696 B.n603 B.n18 10.6151
R697 B.n603 B.n602 10.6151
R698 B.n602 B.n601 10.6151
R699 B.n601 B.n20 10.6151
R700 B.n597 B.n20 10.6151
R701 B.n597 B.n596 10.6151
R702 B.n596 B.n595 10.6151
R703 B.n595 B.n22 10.6151
R704 B.n591 B.n22 10.6151
R705 B.n591 B.n590 10.6151
R706 B.n590 B.n589 10.6151
R707 B.n589 B.n24 10.6151
R708 B.n585 B.n24 10.6151
R709 B.n585 B.n584 10.6151
R710 B.n584 B.n583 10.6151
R711 B.n583 B.n26 10.6151
R712 B.n579 B.n26 10.6151
R713 B.n579 B.n578 10.6151
R714 B.n578 B.n577 10.6151
R715 B.n577 B.n28 10.6151
R716 B.n573 B.n28 10.6151
R717 B.n573 B.n572 10.6151
R718 B.n572 B.n571 10.6151
R719 B.n571 B.n30 10.6151
R720 B.n567 B.n30 10.6151
R721 B.n567 B.n566 10.6151
R722 B.n566 B.n565 10.6151
R723 B.n565 B.n32 10.6151
R724 B.n561 B.n32 10.6151
R725 B.n561 B.n560 10.6151
R726 B.n560 B.n559 10.6151
R727 B.n559 B.n34 10.6151
R728 B.n555 B.n34 10.6151
R729 B.n555 B.n554 10.6151
R730 B.n554 B.n553 10.6151
R731 B.n553 B.n36 10.6151
R732 B.n549 B.n36 10.6151
R733 B.n549 B.n548 10.6151
R734 B.n548 B.n547 10.6151
R735 B.n547 B.n38 10.6151
R736 B.n543 B.n38 10.6151
R737 B.n543 B.n542 10.6151
R738 B.n540 B.n42 10.6151
R739 B.n536 B.n42 10.6151
R740 B.n536 B.n535 10.6151
R741 B.n535 B.n534 10.6151
R742 B.n534 B.n44 10.6151
R743 B.n530 B.n44 10.6151
R744 B.n530 B.n529 10.6151
R745 B.n529 B.n528 10.6151
R746 B.n528 B.n46 10.6151
R747 B.n524 B.n523 10.6151
R748 B.n523 B.n522 10.6151
R749 B.n522 B.n51 10.6151
R750 B.n518 B.n51 10.6151
R751 B.n518 B.n517 10.6151
R752 B.n517 B.n516 10.6151
R753 B.n516 B.n53 10.6151
R754 B.n512 B.n53 10.6151
R755 B.n512 B.n511 10.6151
R756 B.n511 B.n510 10.6151
R757 B.n510 B.n55 10.6151
R758 B.n506 B.n55 10.6151
R759 B.n506 B.n505 10.6151
R760 B.n505 B.n504 10.6151
R761 B.n504 B.n57 10.6151
R762 B.n500 B.n57 10.6151
R763 B.n500 B.n499 10.6151
R764 B.n499 B.n498 10.6151
R765 B.n498 B.n59 10.6151
R766 B.n494 B.n59 10.6151
R767 B.n494 B.n493 10.6151
R768 B.n493 B.n492 10.6151
R769 B.n492 B.n61 10.6151
R770 B.n488 B.n61 10.6151
R771 B.n488 B.n487 10.6151
R772 B.n487 B.n486 10.6151
R773 B.n486 B.n63 10.6151
R774 B.n482 B.n63 10.6151
R775 B.n482 B.n481 10.6151
R776 B.n481 B.n480 10.6151
R777 B.n480 B.n65 10.6151
R778 B.n476 B.n65 10.6151
R779 B.n476 B.n475 10.6151
R780 B.n475 B.n474 10.6151
R781 B.n474 B.n67 10.6151
R782 B.n470 B.n67 10.6151
R783 B.n470 B.n469 10.6151
R784 B.n469 B.n468 10.6151
R785 B.n468 B.n69 10.6151
R786 B.n464 B.n69 10.6151
R787 B.n464 B.n463 10.6151
R788 B.n463 B.n462 10.6151
R789 B.n462 B.n71 10.6151
R790 B.n458 B.n71 10.6151
R791 B.n458 B.n457 10.6151
R792 B.n457 B.n456 10.6151
R793 B.n456 B.n73 10.6151
R794 B.n452 B.n73 10.6151
R795 B.n452 B.n451 10.6151
R796 B.n451 B.n450 10.6151
R797 B.n378 B.n99 10.6151
R798 B.n379 B.n378 10.6151
R799 B.n380 B.n379 10.6151
R800 B.n380 B.n97 10.6151
R801 B.n384 B.n97 10.6151
R802 B.n385 B.n384 10.6151
R803 B.n386 B.n385 10.6151
R804 B.n386 B.n95 10.6151
R805 B.n390 B.n95 10.6151
R806 B.n391 B.n390 10.6151
R807 B.n392 B.n391 10.6151
R808 B.n392 B.n93 10.6151
R809 B.n396 B.n93 10.6151
R810 B.n397 B.n396 10.6151
R811 B.n398 B.n397 10.6151
R812 B.n398 B.n91 10.6151
R813 B.n402 B.n91 10.6151
R814 B.n403 B.n402 10.6151
R815 B.n404 B.n403 10.6151
R816 B.n404 B.n89 10.6151
R817 B.n408 B.n89 10.6151
R818 B.n409 B.n408 10.6151
R819 B.n410 B.n409 10.6151
R820 B.n410 B.n87 10.6151
R821 B.n414 B.n87 10.6151
R822 B.n415 B.n414 10.6151
R823 B.n416 B.n415 10.6151
R824 B.n416 B.n85 10.6151
R825 B.n420 B.n85 10.6151
R826 B.n421 B.n420 10.6151
R827 B.n422 B.n421 10.6151
R828 B.n422 B.n83 10.6151
R829 B.n426 B.n83 10.6151
R830 B.n427 B.n426 10.6151
R831 B.n428 B.n427 10.6151
R832 B.n428 B.n81 10.6151
R833 B.n432 B.n81 10.6151
R834 B.n433 B.n432 10.6151
R835 B.n434 B.n433 10.6151
R836 B.n434 B.n79 10.6151
R837 B.n438 B.n79 10.6151
R838 B.n439 B.n438 10.6151
R839 B.n440 B.n439 10.6151
R840 B.n440 B.n77 10.6151
R841 B.n444 B.n77 10.6151
R842 B.n445 B.n444 10.6151
R843 B.n446 B.n445 10.6151
R844 B.n446 B.n75 10.6151
R845 B.n206 B.n159 10.6151
R846 B.n210 B.n159 10.6151
R847 B.n211 B.n210 10.6151
R848 B.n212 B.n211 10.6151
R849 B.n212 B.n157 10.6151
R850 B.n216 B.n157 10.6151
R851 B.n217 B.n216 10.6151
R852 B.n218 B.n217 10.6151
R853 B.n218 B.n155 10.6151
R854 B.n222 B.n155 10.6151
R855 B.n223 B.n222 10.6151
R856 B.n224 B.n223 10.6151
R857 B.n224 B.n153 10.6151
R858 B.n228 B.n153 10.6151
R859 B.n229 B.n228 10.6151
R860 B.n230 B.n229 10.6151
R861 B.n230 B.n151 10.6151
R862 B.n234 B.n151 10.6151
R863 B.n235 B.n234 10.6151
R864 B.n236 B.n235 10.6151
R865 B.n236 B.n149 10.6151
R866 B.n240 B.n149 10.6151
R867 B.n241 B.n240 10.6151
R868 B.n242 B.n241 10.6151
R869 B.n242 B.n147 10.6151
R870 B.n246 B.n147 10.6151
R871 B.n247 B.n246 10.6151
R872 B.n248 B.n247 10.6151
R873 B.n248 B.n145 10.6151
R874 B.n252 B.n145 10.6151
R875 B.n253 B.n252 10.6151
R876 B.n254 B.n253 10.6151
R877 B.n254 B.n143 10.6151
R878 B.n258 B.n143 10.6151
R879 B.n259 B.n258 10.6151
R880 B.n260 B.n259 10.6151
R881 B.n260 B.n141 10.6151
R882 B.n264 B.n141 10.6151
R883 B.n265 B.n264 10.6151
R884 B.n266 B.n265 10.6151
R885 B.n266 B.n139 10.6151
R886 B.n270 B.n139 10.6151
R887 B.n271 B.n270 10.6151
R888 B.n272 B.n271 10.6151
R889 B.n272 B.n137 10.6151
R890 B.n276 B.n137 10.6151
R891 B.n277 B.n276 10.6151
R892 B.n278 B.n277 10.6151
R893 B.n278 B.n135 10.6151
R894 B.n282 B.n135 10.6151
R895 B.n285 B.n284 10.6151
R896 B.n285 B.n131 10.6151
R897 B.n289 B.n131 10.6151
R898 B.n290 B.n289 10.6151
R899 B.n291 B.n290 10.6151
R900 B.n291 B.n129 10.6151
R901 B.n295 B.n129 10.6151
R902 B.n296 B.n295 10.6151
R903 B.n297 B.n296 10.6151
R904 B.n301 B.n300 10.6151
R905 B.n302 B.n301 10.6151
R906 B.n302 B.n123 10.6151
R907 B.n306 B.n123 10.6151
R908 B.n307 B.n306 10.6151
R909 B.n308 B.n307 10.6151
R910 B.n308 B.n121 10.6151
R911 B.n312 B.n121 10.6151
R912 B.n313 B.n312 10.6151
R913 B.n314 B.n313 10.6151
R914 B.n314 B.n119 10.6151
R915 B.n318 B.n119 10.6151
R916 B.n319 B.n318 10.6151
R917 B.n320 B.n319 10.6151
R918 B.n320 B.n117 10.6151
R919 B.n324 B.n117 10.6151
R920 B.n325 B.n324 10.6151
R921 B.n326 B.n325 10.6151
R922 B.n326 B.n115 10.6151
R923 B.n330 B.n115 10.6151
R924 B.n331 B.n330 10.6151
R925 B.n332 B.n331 10.6151
R926 B.n332 B.n113 10.6151
R927 B.n336 B.n113 10.6151
R928 B.n337 B.n336 10.6151
R929 B.n338 B.n337 10.6151
R930 B.n338 B.n111 10.6151
R931 B.n342 B.n111 10.6151
R932 B.n343 B.n342 10.6151
R933 B.n344 B.n343 10.6151
R934 B.n344 B.n109 10.6151
R935 B.n348 B.n109 10.6151
R936 B.n349 B.n348 10.6151
R937 B.n350 B.n349 10.6151
R938 B.n350 B.n107 10.6151
R939 B.n354 B.n107 10.6151
R940 B.n355 B.n354 10.6151
R941 B.n356 B.n355 10.6151
R942 B.n356 B.n105 10.6151
R943 B.n360 B.n105 10.6151
R944 B.n361 B.n360 10.6151
R945 B.n362 B.n361 10.6151
R946 B.n362 B.n103 10.6151
R947 B.n366 B.n103 10.6151
R948 B.n367 B.n366 10.6151
R949 B.n368 B.n367 10.6151
R950 B.n368 B.n101 10.6151
R951 B.n372 B.n101 10.6151
R952 B.n373 B.n372 10.6151
R953 B.n374 B.n373 10.6151
R954 B.n205 B.n204 10.6151
R955 B.n204 B.n161 10.6151
R956 B.n200 B.n161 10.6151
R957 B.n200 B.n199 10.6151
R958 B.n199 B.n198 10.6151
R959 B.n198 B.n163 10.6151
R960 B.n194 B.n163 10.6151
R961 B.n194 B.n193 10.6151
R962 B.n193 B.n192 10.6151
R963 B.n192 B.n165 10.6151
R964 B.n188 B.n165 10.6151
R965 B.n188 B.n187 10.6151
R966 B.n187 B.n186 10.6151
R967 B.n186 B.n167 10.6151
R968 B.n182 B.n167 10.6151
R969 B.n182 B.n181 10.6151
R970 B.n181 B.n180 10.6151
R971 B.n180 B.n169 10.6151
R972 B.n176 B.n169 10.6151
R973 B.n176 B.n175 10.6151
R974 B.n175 B.n174 10.6151
R975 B.n174 B.n171 10.6151
R976 B.n171 B.n0 10.6151
R977 B.n651 B.n1 10.6151
R978 B.n651 B.n650 10.6151
R979 B.n650 B.n649 10.6151
R980 B.n649 B.n4 10.6151
R981 B.n645 B.n4 10.6151
R982 B.n645 B.n644 10.6151
R983 B.n644 B.n643 10.6151
R984 B.n643 B.n6 10.6151
R985 B.n639 B.n6 10.6151
R986 B.n639 B.n638 10.6151
R987 B.n638 B.n637 10.6151
R988 B.n637 B.n8 10.6151
R989 B.n633 B.n8 10.6151
R990 B.n633 B.n632 10.6151
R991 B.n632 B.n631 10.6151
R992 B.n631 B.n10 10.6151
R993 B.n627 B.n10 10.6151
R994 B.n627 B.n626 10.6151
R995 B.n626 B.n625 10.6151
R996 B.n625 B.n12 10.6151
R997 B.n621 B.n12 10.6151
R998 B.n621 B.n620 10.6151
R999 B.n620 B.n619 10.6151
R1000 B.n542 B.n541 9.36635
R1001 B.n524 B.n50 9.36635
R1002 B.n283 B.n282 9.36635
R1003 B.n300 B.n127 9.36635
R1004 B.n655 B.n0 2.81026
R1005 B.n655 B.n1 2.81026
R1006 B.n541 B.n540 1.24928
R1007 B.n50 B.n46 1.24928
R1008 B.n284 B.n283 1.24928
R1009 B.n297 B.n127 1.24928
C0 w_n2062_n4022# VTAIL 3.2369f
C1 VTAIL B 4.29762f
C2 VDD1 VTAIL 5.91836f
C3 VN VDD2 3.42558f
C4 w_n2062_n4022# VP 3.15659f
C5 B VP 1.48486f
C6 VDD1 VP 3.59925f
C7 w_n2062_n4022# B 9.51018f
C8 VTAIL VN 2.92598f
C9 w_n2062_n4022# VDD1 1.98666f
C10 VDD1 B 1.9364f
C11 VN VP 5.9671f
C12 w_n2062_n4022# VN 2.89436f
C13 VN B 1.05455f
C14 VDD1 VN 0.14803f
C15 VTAIL VDD2 5.96659f
C16 VP VDD2 0.324951f
C17 w_n2062_n4022# VDD2 2.01016f
C18 B VDD2 1.9647f
C19 VTAIL VP 2.94034f
C20 VDD1 VDD2 0.651091f
C21 VDD2 VSUBS 0.99778f
C22 VDD1 VSUBS 4.7942f
C23 VTAIL VSUBS 1.112536f
C24 VN VSUBS 8.47045f
C25 VP VSUBS 1.746227f
C26 B VSUBS 4.034677f
C27 w_n2062_n4022# VSUBS 0.101673p
C28 B.n0 VSUBS 0.003635f
C29 B.n1 VSUBS 0.003635f
C30 B.n2 VSUBS 0.005748f
C31 B.n3 VSUBS 0.005748f
C32 B.n4 VSUBS 0.005748f
C33 B.n5 VSUBS 0.005748f
C34 B.n6 VSUBS 0.005748f
C35 B.n7 VSUBS 0.005748f
C36 B.n8 VSUBS 0.005748f
C37 B.n9 VSUBS 0.005748f
C38 B.n10 VSUBS 0.005748f
C39 B.n11 VSUBS 0.005748f
C40 B.n12 VSUBS 0.005748f
C41 B.n13 VSUBS 0.005748f
C42 B.n14 VSUBS 0.014331f
C43 B.n15 VSUBS 0.005748f
C44 B.n16 VSUBS 0.005748f
C45 B.n17 VSUBS 0.005748f
C46 B.n18 VSUBS 0.005748f
C47 B.n19 VSUBS 0.005748f
C48 B.n20 VSUBS 0.005748f
C49 B.n21 VSUBS 0.005748f
C50 B.n22 VSUBS 0.005748f
C51 B.n23 VSUBS 0.005748f
C52 B.n24 VSUBS 0.005748f
C53 B.n25 VSUBS 0.005748f
C54 B.n26 VSUBS 0.005748f
C55 B.n27 VSUBS 0.005748f
C56 B.n28 VSUBS 0.005748f
C57 B.n29 VSUBS 0.005748f
C58 B.n30 VSUBS 0.005748f
C59 B.n31 VSUBS 0.005748f
C60 B.n32 VSUBS 0.005748f
C61 B.n33 VSUBS 0.005748f
C62 B.n34 VSUBS 0.005748f
C63 B.n35 VSUBS 0.005748f
C64 B.n36 VSUBS 0.005748f
C65 B.n37 VSUBS 0.005748f
C66 B.n38 VSUBS 0.005748f
C67 B.n39 VSUBS 0.005748f
C68 B.t11 VSUBS 0.418027f
C69 B.t10 VSUBS 0.434097f
C70 B.t9 VSUBS 1.34175f
C71 B.n40 VSUBS 0.22652f
C72 B.n41 VSUBS 0.058419f
C73 B.n42 VSUBS 0.005748f
C74 B.n43 VSUBS 0.005748f
C75 B.n44 VSUBS 0.005748f
C76 B.n45 VSUBS 0.005748f
C77 B.n46 VSUBS 0.003212f
C78 B.n47 VSUBS 0.005748f
C79 B.t5 VSUBS 0.418016f
C80 B.t4 VSUBS 0.434088f
C81 B.t3 VSUBS 1.34175f
C82 B.n48 VSUBS 0.226529f
C83 B.n49 VSUBS 0.058431f
C84 B.n50 VSUBS 0.013317f
C85 B.n51 VSUBS 0.005748f
C86 B.n52 VSUBS 0.005748f
C87 B.n53 VSUBS 0.005748f
C88 B.n54 VSUBS 0.005748f
C89 B.n55 VSUBS 0.005748f
C90 B.n56 VSUBS 0.005748f
C91 B.n57 VSUBS 0.005748f
C92 B.n58 VSUBS 0.005748f
C93 B.n59 VSUBS 0.005748f
C94 B.n60 VSUBS 0.005748f
C95 B.n61 VSUBS 0.005748f
C96 B.n62 VSUBS 0.005748f
C97 B.n63 VSUBS 0.005748f
C98 B.n64 VSUBS 0.005748f
C99 B.n65 VSUBS 0.005748f
C100 B.n66 VSUBS 0.005748f
C101 B.n67 VSUBS 0.005748f
C102 B.n68 VSUBS 0.005748f
C103 B.n69 VSUBS 0.005748f
C104 B.n70 VSUBS 0.005748f
C105 B.n71 VSUBS 0.005748f
C106 B.n72 VSUBS 0.005748f
C107 B.n73 VSUBS 0.005748f
C108 B.n74 VSUBS 0.005748f
C109 B.n75 VSUBS 0.014205f
C110 B.n76 VSUBS 0.005748f
C111 B.n77 VSUBS 0.005748f
C112 B.n78 VSUBS 0.005748f
C113 B.n79 VSUBS 0.005748f
C114 B.n80 VSUBS 0.005748f
C115 B.n81 VSUBS 0.005748f
C116 B.n82 VSUBS 0.005748f
C117 B.n83 VSUBS 0.005748f
C118 B.n84 VSUBS 0.005748f
C119 B.n85 VSUBS 0.005748f
C120 B.n86 VSUBS 0.005748f
C121 B.n87 VSUBS 0.005748f
C122 B.n88 VSUBS 0.005748f
C123 B.n89 VSUBS 0.005748f
C124 B.n90 VSUBS 0.005748f
C125 B.n91 VSUBS 0.005748f
C126 B.n92 VSUBS 0.005748f
C127 B.n93 VSUBS 0.005748f
C128 B.n94 VSUBS 0.005748f
C129 B.n95 VSUBS 0.005748f
C130 B.n96 VSUBS 0.005748f
C131 B.n97 VSUBS 0.005748f
C132 B.n98 VSUBS 0.005748f
C133 B.n99 VSUBS 0.013562f
C134 B.n100 VSUBS 0.005748f
C135 B.n101 VSUBS 0.005748f
C136 B.n102 VSUBS 0.005748f
C137 B.n103 VSUBS 0.005748f
C138 B.n104 VSUBS 0.005748f
C139 B.n105 VSUBS 0.005748f
C140 B.n106 VSUBS 0.005748f
C141 B.n107 VSUBS 0.005748f
C142 B.n108 VSUBS 0.005748f
C143 B.n109 VSUBS 0.005748f
C144 B.n110 VSUBS 0.005748f
C145 B.n111 VSUBS 0.005748f
C146 B.n112 VSUBS 0.005748f
C147 B.n113 VSUBS 0.005748f
C148 B.n114 VSUBS 0.005748f
C149 B.n115 VSUBS 0.005748f
C150 B.n116 VSUBS 0.005748f
C151 B.n117 VSUBS 0.005748f
C152 B.n118 VSUBS 0.005748f
C153 B.n119 VSUBS 0.005748f
C154 B.n120 VSUBS 0.005748f
C155 B.n121 VSUBS 0.005748f
C156 B.n122 VSUBS 0.005748f
C157 B.n123 VSUBS 0.005748f
C158 B.n124 VSUBS 0.005748f
C159 B.t1 VSUBS 0.418016f
C160 B.t2 VSUBS 0.434088f
C161 B.t0 VSUBS 1.34175f
C162 B.n125 VSUBS 0.226529f
C163 B.n126 VSUBS 0.058431f
C164 B.n127 VSUBS 0.013317f
C165 B.n128 VSUBS 0.005748f
C166 B.n129 VSUBS 0.005748f
C167 B.n130 VSUBS 0.005748f
C168 B.n131 VSUBS 0.005748f
C169 B.n132 VSUBS 0.005748f
C170 B.t7 VSUBS 0.418027f
C171 B.t8 VSUBS 0.434097f
C172 B.t6 VSUBS 1.34175f
C173 B.n133 VSUBS 0.22652f
C174 B.n134 VSUBS 0.058419f
C175 B.n135 VSUBS 0.005748f
C176 B.n136 VSUBS 0.005748f
C177 B.n137 VSUBS 0.005748f
C178 B.n138 VSUBS 0.005748f
C179 B.n139 VSUBS 0.005748f
C180 B.n140 VSUBS 0.005748f
C181 B.n141 VSUBS 0.005748f
C182 B.n142 VSUBS 0.005748f
C183 B.n143 VSUBS 0.005748f
C184 B.n144 VSUBS 0.005748f
C185 B.n145 VSUBS 0.005748f
C186 B.n146 VSUBS 0.005748f
C187 B.n147 VSUBS 0.005748f
C188 B.n148 VSUBS 0.005748f
C189 B.n149 VSUBS 0.005748f
C190 B.n150 VSUBS 0.005748f
C191 B.n151 VSUBS 0.005748f
C192 B.n152 VSUBS 0.005748f
C193 B.n153 VSUBS 0.005748f
C194 B.n154 VSUBS 0.005748f
C195 B.n155 VSUBS 0.005748f
C196 B.n156 VSUBS 0.005748f
C197 B.n157 VSUBS 0.005748f
C198 B.n158 VSUBS 0.005748f
C199 B.n159 VSUBS 0.005748f
C200 B.n160 VSUBS 0.013562f
C201 B.n161 VSUBS 0.005748f
C202 B.n162 VSUBS 0.005748f
C203 B.n163 VSUBS 0.005748f
C204 B.n164 VSUBS 0.005748f
C205 B.n165 VSUBS 0.005748f
C206 B.n166 VSUBS 0.005748f
C207 B.n167 VSUBS 0.005748f
C208 B.n168 VSUBS 0.005748f
C209 B.n169 VSUBS 0.005748f
C210 B.n170 VSUBS 0.005748f
C211 B.n171 VSUBS 0.005748f
C212 B.n172 VSUBS 0.005748f
C213 B.n173 VSUBS 0.005748f
C214 B.n174 VSUBS 0.005748f
C215 B.n175 VSUBS 0.005748f
C216 B.n176 VSUBS 0.005748f
C217 B.n177 VSUBS 0.005748f
C218 B.n178 VSUBS 0.005748f
C219 B.n179 VSUBS 0.005748f
C220 B.n180 VSUBS 0.005748f
C221 B.n181 VSUBS 0.005748f
C222 B.n182 VSUBS 0.005748f
C223 B.n183 VSUBS 0.005748f
C224 B.n184 VSUBS 0.005748f
C225 B.n185 VSUBS 0.005748f
C226 B.n186 VSUBS 0.005748f
C227 B.n187 VSUBS 0.005748f
C228 B.n188 VSUBS 0.005748f
C229 B.n189 VSUBS 0.005748f
C230 B.n190 VSUBS 0.005748f
C231 B.n191 VSUBS 0.005748f
C232 B.n192 VSUBS 0.005748f
C233 B.n193 VSUBS 0.005748f
C234 B.n194 VSUBS 0.005748f
C235 B.n195 VSUBS 0.005748f
C236 B.n196 VSUBS 0.005748f
C237 B.n197 VSUBS 0.005748f
C238 B.n198 VSUBS 0.005748f
C239 B.n199 VSUBS 0.005748f
C240 B.n200 VSUBS 0.005748f
C241 B.n201 VSUBS 0.005748f
C242 B.n202 VSUBS 0.005748f
C243 B.n203 VSUBS 0.005748f
C244 B.n204 VSUBS 0.005748f
C245 B.n205 VSUBS 0.013562f
C246 B.n206 VSUBS 0.014331f
C247 B.n207 VSUBS 0.014331f
C248 B.n208 VSUBS 0.005748f
C249 B.n209 VSUBS 0.005748f
C250 B.n210 VSUBS 0.005748f
C251 B.n211 VSUBS 0.005748f
C252 B.n212 VSUBS 0.005748f
C253 B.n213 VSUBS 0.005748f
C254 B.n214 VSUBS 0.005748f
C255 B.n215 VSUBS 0.005748f
C256 B.n216 VSUBS 0.005748f
C257 B.n217 VSUBS 0.005748f
C258 B.n218 VSUBS 0.005748f
C259 B.n219 VSUBS 0.005748f
C260 B.n220 VSUBS 0.005748f
C261 B.n221 VSUBS 0.005748f
C262 B.n222 VSUBS 0.005748f
C263 B.n223 VSUBS 0.005748f
C264 B.n224 VSUBS 0.005748f
C265 B.n225 VSUBS 0.005748f
C266 B.n226 VSUBS 0.005748f
C267 B.n227 VSUBS 0.005748f
C268 B.n228 VSUBS 0.005748f
C269 B.n229 VSUBS 0.005748f
C270 B.n230 VSUBS 0.005748f
C271 B.n231 VSUBS 0.005748f
C272 B.n232 VSUBS 0.005748f
C273 B.n233 VSUBS 0.005748f
C274 B.n234 VSUBS 0.005748f
C275 B.n235 VSUBS 0.005748f
C276 B.n236 VSUBS 0.005748f
C277 B.n237 VSUBS 0.005748f
C278 B.n238 VSUBS 0.005748f
C279 B.n239 VSUBS 0.005748f
C280 B.n240 VSUBS 0.005748f
C281 B.n241 VSUBS 0.005748f
C282 B.n242 VSUBS 0.005748f
C283 B.n243 VSUBS 0.005748f
C284 B.n244 VSUBS 0.005748f
C285 B.n245 VSUBS 0.005748f
C286 B.n246 VSUBS 0.005748f
C287 B.n247 VSUBS 0.005748f
C288 B.n248 VSUBS 0.005748f
C289 B.n249 VSUBS 0.005748f
C290 B.n250 VSUBS 0.005748f
C291 B.n251 VSUBS 0.005748f
C292 B.n252 VSUBS 0.005748f
C293 B.n253 VSUBS 0.005748f
C294 B.n254 VSUBS 0.005748f
C295 B.n255 VSUBS 0.005748f
C296 B.n256 VSUBS 0.005748f
C297 B.n257 VSUBS 0.005748f
C298 B.n258 VSUBS 0.005748f
C299 B.n259 VSUBS 0.005748f
C300 B.n260 VSUBS 0.005748f
C301 B.n261 VSUBS 0.005748f
C302 B.n262 VSUBS 0.005748f
C303 B.n263 VSUBS 0.005748f
C304 B.n264 VSUBS 0.005748f
C305 B.n265 VSUBS 0.005748f
C306 B.n266 VSUBS 0.005748f
C307 B.n267 VSUBS 0.005748f
C308 B.n268 VSUBS 0.005748f
C309 B.n269 VSUBS 0.005748f
C310 B.n270 VSUBS 0.005748f
C311 B.n271 VSUBS 0.005748f
C312 B.n272 VSUBS 0.005748f
C313 B.n273 VSUBS 0.005748f
C314 B.n274 VSUBS 0.005748f
C315 B.n275 VSUBS 0.005748f
C316 B.n276 VSUBS 0.005748f
C317 B.n277 VSUBS 0.005748f
C318 B.n278 VSUBS 0.005748f
C319 B.n279 VSUBS 0.005748f
C320 B.n280 VSUBS 0.005748f
C321 B.n281 VSUBS 0.005748f
C322 B.n282 VSUBS 0.00541f
C323 B.n283 VSUBS 0.013317f
C324 B.n284 VSUBS 0.003212f
C325 B.n285 VSUBS 0.005748f
C326 B.n286 VSUBS 0.005748f
C327 B.n287 VSUBS 0.005748f
C328 B.n288 VSUBS 0.005748f
C329 B.n289 VSUBS 0.005748f
C330 B.n290 VSUBS 0.005748f
C331 B.n291 VSUBS 0.005748f
C332 B.n292 VSUBS 0.005748f
C333 B.n293 VSUBS 0.005748f
C334 B.n294 VSUBS 0.005748f
C335 B.n295 VSUBS 0.005748f
C336 B.n296 VSUBS 0.005748f
C337 B.n297 VSUBS 0.003212f
C338 B.n298 VSUBS 0.005748f
C339 B.n299 VSUBS 0.005748f
C340 B.n300 VSUBS 0.00541f
C341 B.n301 VSUBS 0.005748f
C342 B.n302 VSUBS 0.005748f
C343 B.n303 VSUBS 0.005748f
C344 B.n304 VSUBS 0.005748f
C345 B.n305 VSUBS 0.005748f
C346 B.n306 VSUBS 0.005748f
C347 B.n307 VSUBS 0.005748f
C348 B.n308 VSUBS 0.005748f
C349 B.n309 VSUBS 0.005748f
C350 B.n310 VSUBS 0.005748f
C351 B.n311 VSUBS 0.005748f
C352 B.n312 VSUBS 0.005748f
C353 B.n313 VSUBS 0.005748f
C354 B.n314 VSUBS 0.005748f
C355 B.n315 VSUBS 0.005748f
C356 B.n316 VSUBS 0.005748f
C357 B.n317 VSUBS 0.005748f
C358 B.n318 VSUBS 0.005748f
C359 B.n319 VSUBS 0.005748f
C360 B.n320 VSUBS 0.005748f
C361 B.n321 VSUBS 0.005748f
C362 B.n322 VSUBS 0.005748f
C363 B.n323 VSUBS 0.005748f
C364 B.n324 VSUBS 0.005748f
C365 B.n325 VSUBS 0.005748f
C366 B.n326 VSUBS 0.005748f
C367 B.n327 VSUBS 0.005748f
C368 B.n328 VSUBS 0.005748f
C369 B.n329 VSUBS 0.005748f
C370 B.n330 VSUBS 0.005748f
C371 B.n331 VSUBS 0.005748f
C372 B.n332 VSUBS 0.005748f
C373 B.n333 VSUBS 0.005748f
C374 B.n334 VSUBS 0.005748f
C375 B.n335 VSUBS 0.005748f
C376 B.n336 VSUBS 0.005748f
C377 B.n337 VSUBS 0.005748f
C378 B.n338 VSUBS 0.005748f
C379 B.n339 VSUBS 0.005748f
C380 B.n340 VSUBS 0.005748f
C381 B.n341 VSUBS 0.005748f
C382 B.n342 VSUBS 0.005748f
C383 B.n343 VSUBS 0.005748f
C384 B.n344 VSUBS 0.005748f
C385 B.n345 VSUBS 0.005748f
C386 B.n346 VSUBS 0.005748f
C387 B.n347 VSUBS 0.005748f
C388 B.n348 VSUBS 0.005748f
C389 B.n349 VSUBS 0.005748f
C390 B.n350 VSUBS 0.005748f
C391 B.n351 VSUBS 0.005748f
C392 B.n352 VSUBS 0.005748f
C393 B.n353 VSUBS 0.005748f
C394 B.n354 VSUBS 0.005748f
C395 B.n355 VSUBS 0.005748f
C396 B.n356 VSUBS 0.005748f
C397 B.n357 VSUBS 0.005748f
C398 B.n358 VSUBS 0.005748f
C399 B.n359 VSUBS 0.005748f
C400 B.n360 VSUBS 0.005748f
C401 B.n361 VSUBS 0.005748f
C402 B.n362 VSUBS 0.005748f
C403 B.n363 VSUBS 0.005748f
C404 B.n364 VSUBS 0.005748f
C405 B.n365 VSUBS 0.005748f
C406 B.n366 VSUBS 0.005748f
C407 B.n367 VSUBS 0.005748f
C408 B.n368 VSUBS 0.005748f
C409 B.n369 VSUBS 0.005748f
C410 B.n370 VSUBS 0.005748f
C411 B.n371 VSUBS 0.005748f
C412 B.n372 VSUBS 0.005748f
C413 B.n373 VSUBS 0.005748f
C414 B.n374 VSUBS 0.014331f
C415 B.n375 VSUBS 0.014331f
C416 B.n376 VSUBS 0.013562f
C417 B.n377 VSUBS 0.005748f
C418 B.n378 VSUBS 0.005748f
C419 B.n379 VSUBS 0.005748f
C420 B.n380 VSUBS 0.005748f
C421 B.n381 VSUBS 0.005748f
C422 B.n382 VSUBS 0.005748f
C423 B.n383 VSUBS 0.005748f
C424 B.n384 VSUBS 0.005748f
C425 B.n385 VSUBS 0.005748f
C426 B.n386 VSUBS 0.005748f
C427 B.n387 VSUBS 0.005748f
C428 B.n388 VSUBS 0.005748f
C429 B.n389 VSUBS 0.005748f
C430 B.n390 VSUBS 0.005748f
C431 B.n391 VSUBS 0.005748f
C432 B.n392 VSUBS 0.005748f
C433 B.n393 VSUBS 0.005748f
C434 B.n394 VSUBS 0.005748f
C435 B.n395 VSUBS 0.005748f
C436 B.n396 VSUBS 0.005748f
C437 B.n397 VSUBS 0.005748f
C438 B.n398 VSUBS 0.005748f
C439 B.n399 VSUBS 0.005748f
C440 B.n400 VSUBS 0.005748f
C441 B.n401 VSUBS 0.005748f
C442 B.n402 VSUBS 0.005748f
C443 B.n403 VSUBS 0.005748f
C444 B.n404 VSUBS 0.005748f
C445 B.n405 VSUBS 0.005748f
C446 B.n406 VSUBS 0.005748f
C447 B.n407 VSUBS 0.005748f
C448 B.n408 VSUBS 0.005748f
C449 B.n409 VSUBS 0.005748f
C450 B.n410 VSUBS 0.005748f
C451 B.n411 VSUBS 0.005748f
C452 B.n412 VSUBS 0.005748f
C453 B.n413 VSUBS 0.005748f
C454 B.n414 VSUBS 0.005748f
C455 B.n415 VSUBS 0.005748f
C456 B.n416 VSUBS 0.005748f
C457 B.n417 VSUBS 0.005748f
C458 B.n418 VSUBS 0.005748f
C459 B.n419 VSUBS 0.005748f
C460 B.n420 VSUBS 0.005748f
C461 B.n421 VSUBS 0.005748f
C462 B.n422 VSUBS 0.005748f
C463 B.n423 VSUBS 0.005748f
C464 B.n424 VSUBS 0.005748f
C465 B.n425 VSUBS 0.005748f
C466 B.n426 VSUBS 0.005748f
C467 B.n427 VSUBS 0.005748f
C468 B.n428 VSUBS 0.005748f
C469 B.n429 VSUBS 0.005748f
C470 B.n430 VSUBS 0.005748f
C471 B.n431 VSUBS 0.005748f
C472 B.n432 VSUBS 0.005748f
C473 B.n433 VSUBS 0.005748f
C474 B.n434 VSUBS 0.005748f
C475 B.n435 VSUBS 0.005748f
C476 B.n436 VSUBS 0.005748f
C477 B.n437 VSUBS 0.005748f
C478 B.n438 VSUBS 0.005748f
C479 B.n439 VSUBS 0.005748f
C480 B.n440 VSUBS 0.005748f
C481 B.n441 VSUBS 0.005748f
C482 B.n442 VSUBS 0.005748f
C483 B.n443 VSUBS 0.005748f
C484 B.n444 VSUBS 0.005748f
C485 B.n445 VSUBS 0.005748f
C486 B.n446 VSUBS 0.005748f
C487 B.n447 VSUBS 0.005748f
C488 B.n448 VSUBS 0.013562f
C489 B.n449 VSUBS 0.014331f
C490 B.n450 VSUBS 0.013688f
C491 B.n451 VSUBS 0.005748f
C492 B.n452 VSUBS 0.005748f
C493 B.n453 VSUBS 0.005748f
C494 B.n454 VSUBS 0.005748f
C495 B.n455 VSUBS 0.005748f
C496 B.n456 VSUBS 0.005748f
C497 B.n457 VSUBS 0.005748f
C498 B.n458 VSUBS 0.005748f
C499 B.n459 VSUBS 0.005748f
C500 B.n460 VSUBS 0.005748f
C501 B.n461 VSUBS 0.005748f
C502 B.n462 VSUBS 0.005748f
C503 B.n463 VSUBS 0.005748f
C504 B.n464 VSUBS 0.005748f
C505 B.n465 VSUBS 0.005748f
C506 B.n466 VSUBS 0.005748f
C507 B.n467 VSUBS 0.005748f
C508 B.n468 VSUBS 0.005748f
C509 B.n469 VSUBS 0.005748f
C510 B.n470 VSUBS 0.005748f
C511 B.n471 VSUBS 0.005748f
C512 B.n472 VSUBS 0.005748f
C513 B.n473 VSUBS 0.005748f
C514 B.n474 VSUBS 0.005748f
C515 B.n475 VSUBS 0.005748f
C516 B.n476 VSUBS 0.005748f
C517 B.n477 VSUBS 0.005748f
C518 B.n478 VSUBS 0.005748f
C519 B.n479 VSUBS 0.005748f
C520 B.n480 VSUBS 0.005748f
C521 B.n481 VSUBS 0.005748f
C522 B.n482 VSUBS 0.005748f
C523 B.n483 VSUBS 0.005748f
C524 B.n484 VSUBS 0.005748f
C525 B.n485 VSUBS 0.005748f
C526 B.n486 VSUBS 0.005748f
C527 B.n487 VSUBS 0.005748f
C528 B.n488 VSUBS 0.005748f
C529 B.n489 VSUBS 0.005748f
C530 B.n490 VSUBS 0.005748f
C531 B.n491 VSUBS 0.005748f
C532 B.n492 VSUBS 0.005748f
C533 B.n493 VSUBS 0.005748f
C534 B.n494 VSUBS 0.005748f
C535 B.n495 VSUBS 0.005748f
C536 B.n496 VSUBS 0.005748f
C537 B.n497 VSUBS 0.005748f
C538 B.n498 VSUBS 0.005748f
C539 B.n499 VSUBS 0.005748f
C540 B.n500 VSUBS 0.005748f
C541 B.n501 VSUBS 0.005748f
C542 B.n502 VSUBS 0.005748f
C543 B.n503 VSUBS 0.005748f
C544 B.n504 VSUBS 0.005748f
C545 B.n505 VSUBS 0.005748f
C546 B.n506 VSUBS 0.005748f
C547 B.n507 VSUBS 0.005748f
C548 B.n508 VSUBS 0.005748f
C549 B.n509 VSUBS 0.005748f
C550 B.n510 VSUBS 0.005748f
C551 B.n511 VSUBS 0.005748f
C552 B.n512 VSUBS 0.005748f
C553 B.n513 VSUBS 0.005748f
C554 B.n514 VSUBS 0.005748f
C555 B.n515 VSUBS 0.005748f
C556 B.n516 VSUBS 0.005748f
C557 B.n517 VSUBS 0.005748f
C558 B.n518 VSUBS 0.005748f
C559 B.n519 VSUBS 0.005748f
C560 B.n520 VSUBS 0.005748f
C561 B.n521 VSUBS 0.005748f
C562 B.n522 VSUBS 0.005748f
C563 B.n523 VSUBS 0.005748f
C564 B.n524 VSUBS 0.00541f
C565 B.n525 VSUBS 0.005748f
C566 B.n526 VSUBS 0.005748f
C567 B.n527 VSUBS 0.005748f
C568 B.n528 VSUBS 0.005748f
C569 B.n529 VSUBS 0.005748f
C570 B.n530 VSUBS 0.005748f
C571 B.n531 VSUBS 0.005748f
C572 B.n532 VSUBS 0.005748f
C573 B.n533 VSUBS 0.005748f
C574 B.n534 VSUBS 0.005748f
C575 B.n535 VSUBS 0.005748f
C576 B.n536 VSUBS 0.005748f
C577 B.n537 VSUBS 0.005748f
C578 B.n538 VSUBS 0.005748f
C579 B.n539 VSUBS 0.005748f
C580 B.n540 VSUBS 0.003212f
C581 B.n541 VSUBS 0.013317f
C582 B.n542 VSUBS 0.00541f
C583 B.n543 VSUBS 0.005748f
C584 B.n544 VSUBS 0.005748f
C585 B.n545 VSUBS 0.005748f
C586 B.n546 VSUBS 0.005748f
C587 B.n547 VSUBS 0.005748f
C588 B.n548 VSUBS 0.005748f
C589 B.n549 VSUBS 0.005748f
C590 B.n550 VSUBS 0.005748f
C591 B.n551 VSUBS 0.005748f
C592 B.n552 VSUBS 0.005748f
C593 B.n553 VSUBS 0.005748f
C594 B.n554 VSUBS 0.005748f
C595 B.n555 VSUBS 0.005748f
C596 B.n556 VSUBS 0.005748f
C597 B.n557 VSUBS 0.005748f
C598 B.n558 VSUBS 0.005748f
C599 B.n559 VSUBS 0.005748f
C600 B.n560 VSUBS 0.005748f
C601 B.n561 VSUBS 0.005748f
C602 B.n562 VSUBS 0.005748f
C603 B.n563 VSUBS 0.005748f
C604 B.n564 VSUBS 0.005748f
C605 B.n565 VSUBS 0.005748f
C606 B.n566 VSUBS 0.005748f
C607 B.n567 VSUBS 0.005748f
C608 B.n568 VSUBS 0.005748f
C609 B.n569 VSUBS 0.005748f
C610 B.n570 VSUBS 0.005748f
C611 B.n571 VSUBS 0.005748f
C612 B.n572 VSUBS 0.005748f
C613 B.n573 VSUBS 0.005748f
C614 B.n574 VSUBS 0.005748f
C615 B.n575 VSUBS 0.005748f
C616 B.n576 VSUBS 0.005748f
C617 B.n577 VSUBS 0.005748f
C618 B.n578 VSUBS 0.005748f
C619 B.n579 VSUBS 0.005748f
C620 B.n580 VSUBS 0.005748f
C621 B.n581 VSUBS 0.005748f
C622 B.n582 VSUBS 0.005748f
C623 B.n583 VSUBS 0.005748f
C624 B.n584 VSUBS 0.005748f
C625 B.n585 VSUBS 0.005748f
C626 B.n586 VSUBS 0.005748f
C627 B.n587 VSUBS 0.005748f
C628 B.n588 VSUBS 0.005748f
C629 B.n589 VSUBS 0.005748f
C630 B.n590 VSUBS 0.005748f
C631 B.n591 VSUBS 0.005748f
C632 B.n592 VSUBS 0.005748f
C633 B.n593 VSUBS 0.005748f
C634 B.n594 VSUBS 0.005748f
C635 B.n595 VSUBS 0.005748f
C636 B.n596 VSUBS 0.005748f
C637 B.n597 VSUBS 0.005748f
C638 B.n598 VSUBS 0.005748f
C639 B.n599 VSUBS 0.005748f
C640 B.n600 VSUBS 0.005748f
C641 B.n601 VSUBS 0.005748f
C642 B.n602 VSUBS 0.005748f
C643 B.n603 VSUBS 0.005748f
C644 B.n604 VSUBS 0.005748f
C645 B.n605 VSUBS 0.005748f
C646 B.n606 VSUBS 0.005748f
C647 B.n607 VSUBS 0.005748f
C648 B.n608 VSUBS 0.005748f
C649 B.n609 VSUBS 0.005748f
C650 B.n610 VSUBS 0.005748f
C651 B.n611 VSUBS 0.005748f
C652 B.n612 VSUBS 0.005748f
C653 B.n613 VSUBS 0.005748f
C654 B.n614 VSUBS 0.005748f
C655 B.n615 VSUBS 0.005748f
C656 B.n616 VSUBS 0.005748f
C657 B.n617 VSUBS 0.014331f
C658 B.n618 VSUBS 0.013562f
C659 B.n619 VSUBS 0.013562f
C660 B.n620 VSUBS 0.005748f
C661 B.n621 VSUBS 0.005748f
C662 B.n622 VSUBS 0.005748f
C663 B.n623 VSUBS 0.005748f
C664 B.n624 VSUBS 0.005748f
C665 B.n625 VSUBS 0.005748f
C666 B.n626 VSUBS 0.005748f
C667 B.n627 VSUBS 0.005748f
C668 B.n628 VSUBS 0.005748f
C669 B.n629 VSUBS 0.005748f
C670 B.n630 VSUBS 0.005748f
C671 B.n631 VSUBS 0.005748f
C672 B.n632 VSUBS 0.005748f
C673 B.n633 VSUBS 0.005748f
C674 B.n634 VSUBS 0.005748f
C675 B.n635 VSUBS 0.005748f
C676 B.n636 VSUBS 0.005748f
C677 B.n637 VSUBS 0.005748f
C678 B.n638 VSUBS 0.005748f
C679 B.n639 VSUBS 0.005748f
C680 B.n640 VSUBS 0.005748f
C681 B.n641 VSUBS 0.005748f
C682 B.n642 VSUBS 0.005748f
C683 B.n643 VSUBS 0.005748f
C684 B.n644 VSUBS 0.005748f
C685 B.n645 VSUBS 0.005748f
C686 B.n646 VSUBS 0.005748f
C687 B.n647 VSUBS 0.005748f
C688 B.n648 VSUBS 0.005748f
C689 B.n649 VSUBS 0.005748f
C690 B.n650 VSUBS 0.005748f
C691 B.n651 VSUBS 0.005748f
C692 B.n652 VSUBS 0.005748f
C693 B.n653 VSUBS 0.005748f
C694 B.n654 VSUBS 0.005748f
C695 B.n655 VSUBS 0.013015f
C696 VDD1.t1 VSUBS 2.55433f
C697 VDD1.t0 VSUBS 3.25483f
C698 VP.t0 VSUBS 5.08099f
C699 VP.t1 VSUBS 4.44731f
C700 VP.n0 VSUBS 6.08271f
C701 VDD2.t1 VSUBS 3.89279f
C702 VDD2.t0 VSUBS 3.08367f
C703 VDD2.n0 VSUBS 4.28f
C704 VTAIL.t1 VSUBS 3.40241f
C705 VTAIL.n0 VSUBS 2.95682f
C706 VTAIL.t3 VSUBS 3.40243f
C707 VTAIL.n1 VSUBS 3.00537f
C708 VTAIL.t0 VSUBS 3.40243f
C709 VTAIL.n2 VSUBS 2.78977f
C710 VTAIL.t2 VSUBS 3.40241f
C711 VTAIL.n3 VSUBS 2.68752f
C712 VN.t0 VSUBS 4.2925f
C713 VN.t1 VSUBS 4.90505f
.ends

