* NGSPICE file created from diff_pair_sample_1113.ext - technology: sky130A

.subckt diff_pair_sample_1113 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.8743 pd=17.75 as=6.7938 ps=35.62 w=17.42 l=0.42
X1 VTAIL.t7 VN.t1 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.8743 pd=17.75 as=2.8743 ps=17.75 w=17.42 l=0.42
X2 VDD2.t3 VN.t2 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.7938 pd=35.62 as=2.8743 ps=17.75 w=17.42 l=0.42
X3 VDD1.t5 VP.t0 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=6.7938 pd=35.62 as=2.8743 ps=17.75 w=17.42 l=0.42
X4 VTAIL.t10 VP.t1 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.8743 pd=17.75 as=2.8743 ps=17.75 w=17.42 l=0.42
X5 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=6.7938 pd=35.62 as=0 ps=0 w=17.42 l=0.42
X6 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=6.7938 pd=35.62 as=0 ps=0 w=17.42 l=0.42
X7 VDD1.t3 VP.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.7938 pd=35.62 as=2.8743 ps=17.75 w=17.42 l=0.42
X8 VDD1.t2 VP.t3 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.8743 pd=17.75 as=6.7938 ps=35.62 w=17.42 l=0.42
X9 VDD2.t2 VN.t3 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.8743 pd=17.75 as=6.7938 ps=35.62 w=17.42 l=0.42
X10 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.7938 pd=35.62 as=0 ps=0 w=17.42 l=0.42
X11 VDD2.t1 VN.t4 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=6.7938 pd=35.62 as=2.8743 ps=17.75 w=17.42 l=0.42
X12 VDD1.t1 VP.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.8743 pd=17.75 as=6.7938 ps=35.62 w=17.42 l=0.42
X13 VTAIL.t8 VP.t5 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.8743 pd=17.75 as=2.8743 ps=17.75 w=17.42 l=0.42
X14 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.7938 pd=35.62 as=0 ps=0 w=17.42 l=0.42
X15 VTAIL.t3 VN.t5 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.8743 pd=17.75 as=2.8743 ps=17.75 w=17.42 l=0.42
R0 VN.n0 VN.t2 1118.83
R1 VN.n4 VN.t3 1118.83
R2 VN.n2 VN.t0 1100.1
R3 VN.n6 VN.t4 1100.1
R4 VN.n1 VN.t5 1094.25
R5 VN.n5 VN.t1 1094.25
R6 VN.n3 VN.n2 161.3
R7 VN.n7 VN.n6 161.3
R8 VN.n7 VN.n4 71.5267
R9 VN.n3 VN.n0 71.5267
R10 VN VN.n7 44.688
R11 VN.n2 VN.n1 42.3581
R12 VN.n6 VN.n5 42.3581
R13 VN.n5 VN.n4 18.712
R14 VN.n1 VN.n0 18.712
R15 VN VN.n3 0.0516364
R16 VTAIL.n394 VTAIL.n302 289.615
R17 VTAIL.n94 VTAIL.n2 289.615
R18 VTAIL.n296 VTAIL.n204 289.615
R19 VTAIL.n196 VTAIL.n104 289.615
R20 VTAIL.n335 VTAIL.n334 185
R21 VTAIL.n337 VTAIL.n336 185
R22 VTAIL.n330 VTAIL.n329 185
R23 VTAIL.n343 VTAIL.n342 185
R24 VTAIL.n345 VTAIL.n344 185
R25 VTAIL.n326 VTAIL.n325 185
R26 VTAIL.n351 VTAIL.n350 185
R27 VTAIL.n353 VTAIL.n352 185
R28 VTAIL.n322 VTAIL.n321 185
R29 VTAIL.n359 VTAIL.n358 185
R30 VTAIL.n361 VTAIL.n360 185
R31 VTAIL.n318 VTAIL.n317 185
R32 VTAIL.n367 VTAIL.n366 185
R33 VTAIL.n369 VTAIL.n368 185
R34 VTAIL.n314 VTAIL.n313 185
R35 VTAIL.n376 VTAIL.n375 185
R36 VTAIL.n377 VTAIL.n312 185
R37 VTAIL.n379 VTAIL.n378 185
R38 VTAIL.n310 VTAIL.n309 185
R39 VTAIL.n385 VTAIL.n384 185
R40 VTAIL.n387 VTAIL.n386 185
R41 VTAIL.n306 VTAIL.n305 185
R42 VTAIL.n393 VTAIL.n392 185
R43 VTAIL.n395 VTAIL.n394 185
R44 VTAIL.n35 VTAIL.n34 185
R45 VTAIL.n37 VTAIL.n36 185
R46 VTAIL.n30 VTAIL.n29 185
R47 VTAIL.n43 VTAIL.n42 185
R48 VTAIL.n45 VTAIL.n44 185
R49 VTAIL.n26 VTAIL.n25 185
R50 VTAIL.n51 VTAIL.n50 185
R51 VTAIL.n53 VTAIL.n52 185
R52 VTAIL.n22 VTAIL.n21 185
R53 VTAIL.n59 VTAIL.n58 185
R54 VTAIL.n61 VTAIL.n60 185
R55 VTAIL.n18 VTAIL.n17 185
R56 VTAIL.n67 VTAIL.n66 185
R57 VTAIL.n69 VTAIL.n68 185
R58 VTAIL.n14 VTAIL.n13 185
R59 VTAIL.n76 VTAIL.n75 185
R60 VTAIL.n77 VTAIL.n12 185
R61 VTAIL.n79 VTAIL.n78 185
R62 VTAIL.n10 VTAIL.n9 185
R63 VTAIL.n85 VTAIL.n84 185
R64 VTAIL.n87 VTAIL.n86 185
R65 VTAIL.n6 VTAIL.n5 185
R66 VTAIL.n93 VTAIL.n92 185
R67 VTAIL.n95 VTAIL.n94 185
R68 VTAIL.n297 VTAIL.n296 185
R69 VTAIL.n295 VTAIL.n294 185
R70 VTAIL.n208 VTAIL.n207 185
R71 VTAIL.n289 VTAIL.n288 185
R72 VTAIL.n287 VTAIL.n286 185
R73 VTAIL.n212 VTAIL.n211 185
R74 VTAIL.n216 VTAIL.n214 185
R75 VTAIL.n281 VTAIL.n280 185
R76 VTAIL.n279 VTAIL.n278 185
R77 VTAIL.n218 VTAIL.n217 185
R78 VTAIL.n273 VTAIL.n272 185
R79 VTAIL.n271 VTAIL.n270 185
R80 VTAIL.n222 VTAIL.n221 185
R81 VTAIL.n265 VTAIL.n264 185
R82 VTAIL.n263 VTAIL.n262 185
R83 VTAIL.n226 VTAIL.n225 185
R84 VTAIL.n257 VTAIL.n256 185
R85 VTAIL.n255 VTAIL.n254 185
R86 VTAIL.n230 VTAIL.n229 185
R87 VTAIL.n249 VTAIL.n248 185
R88 VTAIL.n247 VTAIL.n246 185
R89 VTAIL.n234 VTAIL.n233 185
R90 VTAIL.n241 VTAIL.n240 185
R91 VTAIL.n239 VTAIL.n238 185
R92 VTAIL.n197 VTAIL.n196 185
R93 VTAIL.n195 VTAIL.n194 185
R94 VTAIL.n108 VTAIL.n107 185
R95 VTAIL.n189 VTAIL.n188 185
R96 VTAIL.n187 VTAIL.n186 185
R97 VTAIL.n112 VTAIL.n111 185
R98 VTAIL.n116 VTAIL.n114 185
R99 VTAIL.n181 VTAIL.n180 185
R100 VTAIL.n179 VTAIL.n178 185
R101 VTAIL.n118 VTAIL.n117 185
R102 VTAIL.n173 VTAIL.n172 185
R103 VTAIL.n171 VTAIL.n170 185
R104 VTAIL.n122 VTAIL.n121 185
R105 VTAIL.n165 VTAIL.n164 185
R106 VTAIL.n163 VTAIL.n162 185
R107 VTAIL.n126 VTAIL.n125 185
R108 VTAIL.n157 VTAIL.n156 185
R109 VTAIL.n155 VTAIL.n154 185
R110 VTAIL.n130 VTAIL.n129 185
R111 VTAIL.n149 VTAIL.n148 185
R112 VTAIL.n147 VTAIL.n146 185
R113 VTAIL.n134 VTAIL.n133 185
R114 VTAIL.n141 VTAIL.n140 185
R115 VTAIL.n139 VTAIL.n138 185
R116 VTAIL.n333 VTAIL.t6 147.659
R117 VTAIL.n33 VTAIL.t1 147.659
R118 VTAIL.n237 VTAIL.t9 147.659
R119 VTAIL.n137 VTAIL.t2 147.659
R120 VTAIL.n336 VTAIL.n335 104.615
R121 VTAIL.n336 VTAIL.n329 104.615
R122 VTAIL.n343 VTAIL.n329 104.615
R123 VTAIL.n344 VTAIL.n343 104.615
R124 VTAIL.n344 VTAIL.n325 104.615
R125 VTAIL.n351 VTAIL.n325 104.615
R126 VTAIL.n352 VTAIL.n351 104.615
R127 VTAIL.n352 VTAIL.n321 104.615
R128 VTAIL.n359 VTAIL.n321 104.615
R129 VTAIL.n360 VTAIL.n359 104.615
R130 VTAIL.n360 VTAIL.n317 104.615
R131 VTAIL.n367 VTAIL.n317 104.615
R132 VTAIL.n368 VTAIL.n367 104.615
R133 VTAIL.n368 VTAIL.n313 104.615
R134 VTAIL.n376 VTAIL.n313 104.615
R135 VTAIL.n377 VTAIL.n376 104.615
R136 VTAIL.n378 VTAIL.n377 104.615
R137 VTAIL.n378 VTAIL.n309 104.615
R138 VTAIL.n385 VTAIL.n309 104.615
R139 VTAIL.n386 VTAIL.n385 104.615
R140 VTAIL.n386 VTAIL.n305 104.615
R141 VTAIL.n393 VTAIL.n305 104.615
R142 VTAIL.n394 VTAIL.n393 104.615
R143 VTAIL.n36 VTAIL.n35 104.615
R144 VTAIL.n36 VTAIL.n29 104.615
R145 VTAIL.n43 VTAIL.n29 104.615
R146 VTAIL.n44 VTAIL.n43 104.615
R147 VTAIL.n44 VTAIL.n25 104.615
R148 VTAIL.n51 VTAIL.n25 104.615
R149 VTAIL.n52 VTAIL.n51 104.615
R150 VTAIL.n52 VTAIL.n21 104.615
R151 VTAIL.n59 VTAIL.n21 104.615
R152 VTAIL.n60 VTAIL.n59 104.615
R153 VTAIL.n60 VTAIL.n17 104.615
R154 VTAIL.n67 VTAIL.n17 104.615
R155 VTAIL.n68 VTAIL.n67 104.615
R156 VTAIL.n68 VTAIL.n13 104.615
R157 VTAIL.n76 VTAIL.n13 104.615
R158 VTAIL.n77 VTAIL.n76 104.615
R159 VTAIL.n78 VTAIL.n77 104.615
R160 VTAIL.n78 VTAIL.n9 104.615
R161 VTAIL.n85 VTAIL.n9 104.615
R162 VTAIL.n86 VTAIL.n85 104.615
R163 VTAIL.n86 VTAIL.n5 104.615
R164 VTAIL.n93 VTAIL.n5 104.615
R165 VTAIL.n94 VTAIL.n93 104.615
R166 VTAIL.n296 VTAIL.n295 104.615
R167 VTAIL.n295 VTAIL.n207 104.615
R168 VTAIL.n288 VTAIL.n207 104.615
R169 VTAIL.n288 VTAIL.n287 104.615
R170 VTAIL.n287 VTAIL.n211 104.615
R171 VTAIL.n216 VTAIL.n211 104.615
R172 VTAIL.n280 VTAIL.n216 104.615
R173 VTAIL.n280 VTAIL.n279 104.615
R174 VTAIL.n279 VTAIL.n217 104.615
R175 VTAIL.n272 VTAIL.n217 104.615
R176 VTAIL.n272 VTAIL.n271 104.615
R177 VTAIL.n271 VTAIL.n221 104.615
R178 VTAIL.n264 VTAIL.n221 104.615
R179 VTAIL.n264 VTAIL.n263 104.615
R180 VTAIL.n263 VTAIL.n225 104.615
R181 VTAIL.n256 VTAIL.n225 104.615
R182 VTAIL.n256 VTAIL.n255 104.615
R183 VTAIL.n255 VTAIL.n229 104.615
R184 VTAIL.n248 VTAIL.n229 104.615
R185 VTAIL.n248 VTAIL.n247 104.615
R186 VTAIL.n247 VTAIL.n233 104.615
R187 VTAIL.n240 VTAIL.n233 104.615
R188 VTAIL.n240 VTAIL.n239 104.615
R189 VTAIL.n196 VTAIL.n195 104.615
R190 VTAIL.n195 VTAIL.n107 104.615
R191 VTAIL.n188 VTAIL.n107 104.615
R192 VTAIL.n188 VTAIL.n187 104.615
R193 VTAIL.n187 VTAIL.n111 104.615
R194 VTAIL.n116 VTAIL.n111 104.615
R195 VTAIL.n180 VTAIL.n116 104.615
R196 VTAIL.n180 VTAIL.n179 104.615
R197 VTAIL.n179 VTAIL.n117 104.615
R198 VTAIL.n172 VTAIL.n117 104.615
R199 VTAIL.n172 VTAIL.n171 104.615
R200 VTAIL.n171 VTAIL.n121 104.615
R201 VTAIL.n164 VTAIL.n121 104.615
R202 VTAIL.n164 VTAIL.n163 104.615
R203 VTAIL.n163 VTAIL.n125 104.615
R204 VTAIL.n156 VTAIL.n125 104.615
R205 VTAIL.n156 VTAIL.n155 104.615
R206 VTAIL.n155 VTAIL.n129 104.615
R207 VTAIL.n148 VTAIL.n129 104.615
R208 VTAIL.n148 VTAIL.n147 104.615
R209 VTAIL.n147 VTAIL.n133 104.615
R210 VTAIL.n140 VTAIL.n133 104.615
R211 VTAIL.n140 VTAIL.n139 104.615
R212 VTAIL.n335 VTAIL.t6 52.3082
R213 VTAIL.n35 VTAIL.t1 52.3082
R214 VTAIL.n239 VTAIL.t9 52.3082
R215 VTAIL.n139 VTAIL.t2 52.3082
R216 VTAIL.n203 VTAIL.n202 42.064
R217 VTAIL.n103 VTAIL.n102 42.064
R218 VTAIL.n1 VTAIL.n0 42.0638
R219 VTAIL.n101 VTAIL.n100 42.0638
R220 VTAIL.n399 VTAIL.n398 30.246
R221 VTAIL.n99 VTAIL.n98 30.246
R222 VTAIL.n301 VTAIL.n300 30.246
R223 VTAIL.n201 VTAIL.n200 30.246
R224 VTAIL.n103 VTAIL.n101 28.6772
R225 VTAIL.n399 VTAIL.n301 28.0307
R226 VTAIL.n334 VTAIL.n333 15.6677
R227 VTAIL.n34 VTAIL.n33 15.6677
R228 VTAIL.n238 VTAIL.n237 15.6677
R229 VTAIL.n138 VTAIL.n137 15.6677
R230 VTAIL.n379 VTAIL.n310 13.1884
R231 VTAIL.n79 VTAIL.n10 13.1884
R232 VTAIL.n214 VTAIL.n212 13.1884
R233 VTAIL.n114 VTAIL.n112 13.1884
R234 VTAIL.n337 VTAIL.n332 12.8005
R235 VTAIL.n380 VTAIL.n312 12.8005
R236 VTAIL.n384 VTAIL.n383 12.8005
R237 VTAIL.n37 VTAIL.n32 12.8005
R238 VTAIL.n80 VTAIL.n12 12.8005
R239 VTAIL.n84 VTAIL.n83 12.8005
R240 VTAIL.n286 VTAIL.n285 12.8005
R241 VTAIL.n282 VTAIL.n281 12.8005
R242 VTAIL.n241 VTAIL.n236 12.8005
R243 VTAIL.n186 VTAIL.n185 12.8005
R244 VTAIL.n182 VTAIL.n181 12.8005
R245 VTAIL.n141 VTAIL.n136 12.8005
R246 VTAIL.n338 VTAIL.n330 12.0247
R247 VTAIL.n375 VTAIL.n374 12.0247
R248 VTAIL.n387 VTAIL.n308 12.0247
R249 VTAIL.n38 VTAIL.n30 12.0247
R250 VTAIL.n75 VTAIL.n74 12.0247
R251 VTAIL.n87 VTAIL.n8 12.0247
R252 VTAIL.n289 VTAIL.n210 12.0247
R253 VTAIL.n278 VTAIL.n215 12.0247
R254 VTAIL.n242 VTAIL.n234 12.0247
R255 VTAIL.n189 VTAIL.n110 12.0247
R256 VTAIL.n178 VTAIL.n115 12.0247
R257 VTAIL.n142 VTAIL.n134 12.0247
R258 VTAIL.n342 VTAIL.n341 11.249
R259 VTAIL.n373 VTAIL.n314 11.249
R260 VTAIL.n388 VTAIL.n306 11.249
R261 VTAIL.n42 VTAIL.n41 11.249
R262 VTAIL.n73 VTAIL.n14 11.249
R263 VTAIL.n88 VTAIL.n6 11.249
R264 VTAIL.n290 VTAIL.n208 11.249
R265 VTAIL.n277 VTAIL.n218 11.249
R266 VTAIL.n246 VTAIL.n245 11.249
R267 VTAIL.n190 VTAIL.n108 11.249
R268 VTAIL.n177 VTAIL.n118 11.249
R269 VTAIL.n146 VTAIL.n145 11.249
R270 VTAIL.n345 VTAIL.n328 10.4732
R271 VTAIL.n370 VTAIL.n369 10.4732
R272 VTAIL.n392 VTAIL.n391 10.4732
R273 VTAIL.n45 VTAIL.n28 10.4732
R274 VTAIL.n70 VTAIL.n69 10.4732
R275 VTAIL.n92 VTAIL.n91 10.4732
R276 VTAIL.n294 VTAIL.n293 10.4732
R277 VTAIL.n274 VTAIL.n273 10.4732
R278 VTAIL.n249 VTAIL.n232 10.4732
R279 VTAIL.n194 VTAIL.n193 10.4732
R280 VTAIL.n174 VTAIL.n173 10.4732
R281 VTAIL.n149 VTAIL.n132 10.4732
R282 VTAIL.n346 VTAIL.n326 9.69747
R283 VTAIL.n366 VTAIL.n316 9.69747
R284 VTAIL.n395 VTAIL.n304 9.69747
R285 VTAIL.n46 VTAIL.n26 9.69747
R286 VTAIL.n66 VTAIL.n16 9.69747
R287 VTAIL.n95 VTAIL.n4 9.69747
R288 VTAIL.n297 VTAIL.n206 9.69747
R289 VTAIL.n270 VTAIL.n220 9.69747
R290 VTAIL.n250 VTAIL.n230 9.69747
R291 VTAIL.n197 VTAIL.n106 9.69747
R292 VTAIL.n170 VTAIL.n120 9.69747
R293 VTAIL.n150 VTAIL.n130 9.69747
R294 VTAIL.n398 VTAIL.n397 9.45567
R295 VTAIL.n98 VTAIL.n97 9.45567
R296 VTAIL.n300 VTAIL.n299 9.45567
R297 VTAIL.n200 VTAIL.n199 9.45567
R298 VTAIL.n397 VTAIL.n396 9.3005
R299 VTAIL.n304 VTAIL.n303 9.3005
R300 VTAIL.n391 VTAIL.n390 9.3005
R301 VTAIL.n389 VTAIL.n388 9.3005
R302 VTAIL.n308 VTAIL.n307 9.3005
R303 VTAIL.n383 VTAIL.n382 9.3005
R304 VTAIL.n355 VTAIL.n354 9.3005
R305 VTAIL.n324 VTAIL.n323 9.3005
R306 VTAIL.n349 VTAIL.n348 9.3005
R307 VTAIL.n347 VTAIL.n346 9.3005
R308 VTAIL.n328 VTAIL.n327 9.3005
R309 VTAIL.n341 VTAIL.n340 9.3005
R310 VTAIL.n339 VTAIL.n338 9.3005
R311 VTAIL.n332 VTAIL.n331 9.3005
R312 VTAIL.n357 VTAIL.n356 9.3005
R313 VTAIL.n320 VTAIL.n319 9.3005
R314 VTAIL.n363 VTAIL.n362 9.3005
R315 VTAIL.n365 VTAIL.n364 9.3005
R316 VTAIL.n316 VTAIL.n315 9.3005
R317 VTAIL.n371 VTAIL.n370 9.3005
R318 VTAIL.n373 VTAIL.n372 9.3005
R319 VTAIL.n374 VTAIL.n311 9.3005
R320 VTAIL.n381 VTAIL.n380 9.3005
R321 VTAIL.n97 VTAIL.n96 9.3005
R322 VTAIL.n4 VTAIL.n3 9.3005
R323 VTAIL.n91 VTAIL.n90 9.3005
R324 VTAIL.n89 VTAIL.n88 9.3005
R325 VTAIL.n8 VTAIL.n7 9.3005
R326 VTAIL.n83 VTAIL.n82 9.3005
R327 VTAIL.n55 VTAIL.n54 9.3005
R328 VTAIL.n24 VTAIL.n23 9.3005
R329 VTAIL.n49 VTAIL.n48 9.3005
R330 VTAIL.n47 VTAIL.n46 9.3005
R331 VTAIL.n28 VTAIL.n27 9.3005
R332 VTAIL.n41 VTAIL.n40 9.3005
R333 VTAIL.n39 VTAIL.n38 9.3005
R334 VTAIL.n32 VTAIL.n31 9.3005
R335 VTAIL.n57 VTAIL.n56 9.3005
R336 VTAIL.n20 VTAIL.n19 9.3005
R337 VTAIL.n63 VTAIL.n62 9.3005
R338 VTAIL.n65 VTAIL.n64 9.3005
R339 VTAIL.n16 VTAIL.n15 9.3005
R340 VTAIL.n71 VTAIL.n70 9.3005
R341 VTAIL.n73 VTAIL.n72 9.3005
R342 VTAIL.n74 VTAIL.n11 9.3005
R343 VTAIL.n81 VTAIL.n80 9.3005
R344 VTAIL.n224 VTAIL.n223 9.3005
R345 VTAIL.n267 VTAIL.n266 9.3005
R346 VTAIL.n269 VTAIL.n268 9.3005
R347 VTAIL.n220 VTAIL.n219 9.3005
R348 VTAIL.n275 VTAIL.n274 9.3005
R349 VTAIL.n277 VTAIL.n276 9.3005
R350 VTAIL.n215 VTAIL.n213 9.3005
R351 VTAIL.n283 VTAIL.n282 9.3005
R352 VTAIL.n299 VTAIL.n298 9.3005
R353 VTAIL.n206 VTAIL.n205 9.3005
R354 VTAIL.n293 VTAIL.n292 9.3005
R355 VTAIL.n291 VTAIL.n290 9.3005
R356 VTAIL.n210 VTAIL.n209 9.3005
R357 VTAIL.n285 VTAIL.n284 9.3005
R358 VTAIL.n261 VTAIL.n260 9.3005
R359 VTAIL.n259 VTAIL.n258 9.3005
R360 VTAIL.n228 VTAIL.n227 9.3005
R361 VTAIL.n253 VTAIL.n252 9.3005
R362 VTAIL.n251 VTAIL.n250 9.3005
R363 VTAIL.n232 VTAIL.n231 9.3005
R364 VTAIL.n245 VTAIL.n244 9.3005
R365 VTAIL.n243 VTAIL.n242 9.3005
R366 VTAIL.n236 VTAIL.n235 9.3005
R367 VTAIL.n124 VTAIL.n123 9.3005
R368 VTAIL.n167 VTAIL.n166 9.3005
R369 VTAIL.n169 VTAIL.n168 9.3005
R370 VTAIL.n120 VTAIL.n119 9.3005
R371 VTAIL.n175 VTAIL.n174 9.3005
R372 VTAIL.n177 VTAIL.n176 9.3005
R373 VTAIL.n115 VTAIL.n113 9.3005
R374 VTAIL.n183 VTAIL.n182 9.3005
R375 VTAIL.n199 VTAIL.n198 9.3005
R376 VTAIL.n106 VTAIL.n105 9.3005
R377 VTAIL.n193 VTAIL.n192 9.3005
R378 VTAIL.n191 VTAIL.n190 9.3005
R379 VTAIL.n110 VTAIL.n109 9.3005
R380 VTAIL.n185 VTAIL.n184 9.3005
R381 VTAIL.n161 VTAIL.n160 9.3005
R382 VTAIL.n159 VTAIL.n158 9.3005
R383 VTAIL.n128 VTAIL.n127 9.3005
R384 VTAIL.n153 VTAIL.n152 9.3005
R385 VTAIL.n151 VTAIL.n150 9.3005
R386 VTAIL.n132 VTAIL.n131 9.3005
R387 VTAIL.n145 VTAIL.n144 9.3005
R388 VTAIL.n143 VTAIL.n142 9.3005
R389 VTAIL.n136 VTAIL.n135 9.3005
R390 VTAIL.n350 VTAIL.n349 8.92171
R391 VTAIL.n365 VTAIL.n318 8.92171
R392 VTAIL.n396 VTAIL.n302 8.92171
R393 VTAIL.n50 VTAIL.n49 8.92171
R394 VTAIL.n65 VTAIL.n18 8.92171
R395 VTAIL.n96 VTAIL.n2 8.92171
R396 VTAIL.n298 VTAIL.n204 8.92171
R397 VTAIL.n269 VTAIL.n222 8.92171
R398 VTAIL.n254 VTAIL.n253 8.92171
R399 VTAIL.n198 VTAIL.n104 8.92171
R400 VTAIL.n169 VTAIL.n122 8.92171
R401 VTAIL.n154 VTAIL.n153 8.92171
R402 VTAIL.n353 VTAIL.n324 8.14595
R403 VTAIL.n362 VTAIL.n361 8.14595
R404 VTAIL.n53 VTAIL.n24 8.14595
R405 VTAIL.n62 VTAIL.n61 8.14595
R406 VTAIL.n266 VTAIL.n265 8.14595
R407 VTAIL.n257 VTAIL.n228 8.14595
R408 VTAIL.n166 VTAIL.n165 8.14595
R409 VTAIL.n157 VTAIL.n128 8.14595
R410 VTAIL.n354 VTAIL.n322 7.3702
R411 VTAIL.n358 VTAIL.n320 7.3702
R412 VTAIL.n54 VTAIL.n22 7.3702
R413 VTAIL.n58 VTAIL.n20 7.3702
R414 VTAIL.n262 VTAIL.n224 7.3702
R415 VTAIL.n258 VTAIL.n226 7.3702
R416 VTAIL.n162 VTAIL.n124 7.3702
R417 VTAIL.n158 VTAIL.n126 7.3702
R418 VTAIL.n357 VTAIL.n322 6.59444
R419 VTAIL.n358 VTAIL.n357 6.59444
R420 VTAIL.n57 VTAIL.n22 6.59444
R421 VTAIL.n58 VTAIL.n57 6.59444
R422 VTAIL.n262 VTAIL.n261 6.59444
R423 VTAIL.n261 VTAIL.n226 6.59444
R424 VTAIL.n162 VTAIL.n161 6.59444
R425 VTAIL.n161 VTAIL.n126 6.59444
R426 VTAIL.n354 VTAIL.n353 5.81868
R427 VTAIL.n361 VTAIL.n320 5.81868
R428 VTAIL.n54 VTAIL.n53 5.81868
R429 VTAIL.n61 VTAIL.n20 5.81868
R430 VTAIL.n265 VTAIL.n224 5.81868
R431 VTAIL.n258 VTAIL.n257 5.81868
R432 VTAIL.n165 VTAIL.n124 5.81868
R433 VTAIL.n158 VTAIL.n157 5.81868
R434 VTAIL.n350 VTAIL.n324 5.04292
R435 VTAIL.n362 VTAIL.n318 5.04292
R436 VTAIL.n398 VTAIL.n302 5.04292
R437 VTAIL.n50 VTAIL.n24 5.04292
R438 VTAIL.n62 VTAIL.n18 5.04292
R439 VTAIL.n98 VTAIL.n2 5.04292
R440 VTAIL.n300 VTAIL.n204 5.04292
R441 VTAIL.n266 VTAIL.n222 5.04292
R442 VTAIL.n254 VTAIL.n228 5.04292
R443 VTAIL.n200 VTAIL.n104 5.04292
R444 VTAIL.n166 VTAIL.n122 5.04292
R445 VTAIL.n154 VTAIL.n128 5.04292
R446 VTAIL.n333 VTAIL.n331 4.38563
R447 VTAIL.n33 VTAIL.n31 4.38563
R448 VTAIL.n237 VTAIL.n235 4.38563
R449 VTAIL.n137 VTAIL.n135 4.38563
R450 VTAIL.n349 VTAIL.n326 4.26717
R451 VTAIL.n366 VTAIL.n365 4.26717
R452 VTAIL.n396 VTAIL.n395 4.26717
R453 VTAIL.n49 VTAIL.n26 4.26717
R454 VTAIL.n66 VTAIL.n65 4.26717
R455 VTAIL.n96 VTAIL.n95 4.26717
R456 VTAIL.n298 VTAIL.n297 4.26717
R457 VTAIL.n270 VTAIL.n269 4.26717
R458 VTAIL.n253 VTAIL.n230 4.26717
R459 VTAIL.n198 VTAIL.n197 4.26717
R460 VTAIL.n170 VTAIL.n169 4.26717
R461 VTAIL.n153 VTAIL.n130 4.26717
R462 VTAIL.n346 VTAIL.n345 3.49141
R463 VTAIL.n369 VTAIL.n316 3.49141
R464 VTAIL.n392 VTAIL.n304 3.49141
R465 VTAIL.n46 VTAIL.n45 3.49141
R466 VTAIL.n69 VTAIL.n16 3.49141
R467 VTAIL.n92 VTAIL.n4 3.49141
R468 VTAIL.n294 VTAIL.n206 3.49141
R469 VTAIL.n273 VTAIL.n220 3.49141
R470 VTAIL.n250 VTAIL.n249 3.49141
R471 VTAIL.n194 VTAIL.n106 3.49141
R472 VTAIL.n173 VTAIL.n120 3.49141
R473 VTAIL.n150 VTAIL.n149 3.49141
R474 VTAIL.n342 VTAIL.n328 2.71565
R475 VTAIL.n370 VTAIL.n314 2.71565
R476 VTAIL.n391 VTAIL.n306 2.71565
R477 VTAIL.n42 VTAIL.n28 2.71565
R478 VTAIL.n70 VTAIL.n14 2.71565
R479 VTAIL.n91 VTAIL.n6 2.71565
R480 VTAIL.n293 VTAIL.n208 2.71565
R481 VTAIL.n274 VTAIL.n218 2.71565
R482 VTAIL.n246 VTAIL.n232 2.71565
R483 VTAIL.n193 VTAIL.n108 2.71565
R484 VTAIL.n174 VTAIL.n118 2.71565
R485 VTAIL.n146 VTAIL.n132 2.71565
R486 VTAIL.n341 VTAIL.n330 1.93989
R487 VTAIL.n375 VTAIL.n373 1.93989
R488 VTAIL.n388 VTAIL.n387 1.93989
R489 VTAIL.n41 VTAIL.n30 1.93989
R490 VTAIL.n75 VTAIL.n73 1.93989
R491 VTAIL.n88 VTAIL.n87 1.93989
R492 VTAIL.n290 VTAIL.n289 1.93989
R493 VTAIL.n278 VTAIL.n277 1.93989
R494 VTAIL.n245 VTAIL.n234 1.93989
R495 VTAIL.n190 VTAIL.n189 1.93989
R496 VTAIL.n178 VTAIL.n177 1.93989
R497 VTAIL.n145 VTAIL.n134 1.93989
R498 VTAIL.n338 VTAIL.n337 1.16414
R499 VTAIL.n374 VTAIL.n312 1.16414
R500 VTAIL.n384 VTAIL.n308 1.16414
R501 VTAIL.n38 VTAIL.n37 1.16414
R502 VTAIL.n74 VTAIL.n12 1.16414
R503 VTAIL.n84 VTAIL.n8 1.16414
R504 VTAIL.n286 VTAIL.n210 1.16414
R505 VTAIL.n281 VTAIL.n215 1.16414
R506 VTAIL.n242 VTAIL.n241 1.16414
R507 VTAIL.n186 VTAIL.n110 1.16414
R508 VTAIL.n181 VTAIL.n115 1.16414
R509 VTAIL.n142 VTAIL.n141 1.16414
R510 VTAIL.n0 VTAIL.t4 1.13712
R511 VTAIL.n0 VTAIL.t3 1.13712
R512 VTAIL.n100 VTAIL.t0 1.13712
R513 VTAIL.n100 VTAIL.t10 1.13712
R514 VTAIL.n202 VTAIL.t11 1.13712
R515 VTAIL.n202 VTAIL.t8 1.13712
R516 VTAIL.n102 VTAIL.t5 1.13712
R517 VTAIL.n102 VTAIL.t7 1.13712
R518 VTAIL.n203 VTAIL.n201 0.793603
R519 VTAIL.n99 VTAIL.n1 0.793603
R520 VTAIL.n201 VTAIL.n103 0.647052
R521 VTAIL.n301 VTAIL.n203 0.647052
R522 VTAIL.n101 VTAIL.n99 0.647052
R523 VTAIL VTAIL.n399 0.427224
R524 VTAIL.n334 VTAIL.n332 0.388379
R525 VTAIL.n380 VTAIL.n379 0.388379
R526 VTAIL.n383 VTAIL.n310 0.388379
R527 VTAIL.n34 VTAIL.n32 0.388379
R528 VTAIL.n80 VTAIL.n79 0.388379
R529 VTAIL.n83 VTAIL.n10 0.388379
R530 VTAIL.n285 VTAIL.n212 0.388379
R531 VTAIL.n282 VTAIL.n214 0.388379
R532 VTAIL.n238 VTAIL.n236 0.388379
R533 VTAIL.n185 VTAIL.n112 0.388379
R534 VTAIL.n182 VTAIL.n114 0.388379
R535 VTAIL.n138 VTAIL.n136 0.388379
R536 VTAIL VTAIL.n1 0.220328
R537 VTAIL.n339 VTAIL.n331 0.155672
R538 VTAIL.n340 VTAIL.n339 0.155672
R539 VTAIL.n340 VTAIL.n327 0.155672
R540 VTAIL.n347 VTAIL.n327 0.155672
R541 VTAIL.n348 VTAIL.n347 0.155672
R542 VTAIL.n348 VTAIL.n323 0.155672
R543 VTAIL.n355 VTAIL.n323 0.155672
R544 VTAIL.n356 VTAIL.n355 0.155672
R545 VTAIL.n356 VTAIL.n319 0.155672
R546 VTAIL.n363 VTAIL.n319 0.155672
R547 VTAIL.n364 VTAIL.n363 0.155672
R548 VTAIL.n364 VTAIL.n315 0.155672
R549 VTAIL.n371 VTAIL.n315 0.155672
R550 VTAIL.n372 VTAIL.n371 0.155672
R551 VTAIL.n372 VTAIL.n311 0.155672
R552 VTAIL.n381 VTAIL.n311 0.155672
R553 VTAIL.n382 VTAIL.n381 0.155672
R554 VTAIL.n382 VTAIL.n307 0.155672
R555 VTAIL.n389 VTAIL.n307 0.155672
R556 VTAIL.n390 VTAIL.n389 0.155672
R557 VTAIL.n390 VTAIL.n303 0.155672
R558 VTAIL.n397 VTAIL.n303 0.155672
R559 VTAIL.n39 VTAIL.n31 0.155672
R560 VTAIL.n40 VTAIL.n39 0.155672
R561 VTAIL.n40 VTAIL.n27 0.155672
R562 VTAIL.n47 VTAIL.n27 0.155672
R563 VTAIL.n48 VTAIL.n47 0.155672
R564 VTAIL.n48 VTAIL.n23 0.155672
R565 VTAIL.n55 VTAIL.n23 0.155672
R566 VTAIL.n56 VTAIL.n55 0.155672
R567 VTAIL.n56 VTAIL.n19 0.155672
R568 VTAIL.n63 VTAIL.n19 0.155672
R569 VTAIL.n64 VTAIL.n63 0.155672
R570 VTAIL.n64 VTAIL.n15 0.155672
R571 VTAIL.n71 VTAIL.n15 0.155672
R572 VTAIL.n72 VTAIL.n71 0.155672
R573 VTAIL.n72 VTAIL.n11 0.155672
R574 VTAIL.n81 VTAIL.n11 0.155672
R575 VTAIL.n82 VTAIL.n81 0.155672
R576 VTAIL.n82 VTAIL.n7 0.155672
R577 VTAIL.n89 VTAIL.n7 0.155672
R578 VTAIL.n90 VTAIL.n89 0.155672
R579 VTAIL.n90 VTAIL.n3 0.155672
R580 VTAIL.n97 VTAIL.n3 0.155672
R581 VTAIL.n299 VTAIL.n205 0.155672
R582 VTAIL.n292 VTAIL.n205 0.155672
R583 VTAIL.n292 VTAIL.n291 0.155672
R584 VTAIL.n291 VTAIL.n209 0.155672
R585 VTAIL.n284 VTAIL.n209 0.155672
R586 VTAIL.n284 VTAIL.n283 0.155672
R587 VTAIL.n283 VTAIL.n213 0.155672
R588 VTAIL.n276 VTAIL.n213 0.155672
R589 VTAIL.n276 VTAIL.n275 0.155672
R590 VTAIL.n275 VTAIL.n219 0.155672
R591 VTAIL.n268 VTAIL.n219 0.155672
R592 VTAIL.n268 VTAIL.n267 0.155672
R593 VTAIL.n267 VTAIL.n223 0.155672
R594 VTAIL.n260 VTAIL.n223 0.155672
R595 VTAIL.n260 VTAIL.n259 0.155672
R596 VTAIL.n259 VTAIL.n227 0.155672
R597 VTAIL.n252 VTAIL.n227 0.155672
R598 VTAIL.n252 VTAIL.n251 0.155672
R599 VTAIL.n251 VTAIL.n231 0.155672
R600 VTAIL.n244 VTAIL.n231 0.155672
R601 VTAIL.n244 VTAIL.n243 0.155672
R602 VTAIL.n243 VTAIL.n235 0.155672
R603 VTAIL.n199 VTAIL.n105 0.155672
R604 VTAIL.n192 VTAIL.n105 0.155672
R605 VTAIL.n192 VTAIL.n191 0.155672
R606 VTAIL.n191 VTAIL.n109 0.155672
R607 VTAIL.n184 VTAIL.n109 0.155672
R608 VTAIL.n184 VTAIL.n183 0.155672
R609 VTAIL.n183 VTAIL.n113 0.155672
R610 VTAIL.n176 VTAIL.n113 0.155672
R611 VTAIL.n176 VTAIL.n175 0.155672
R612 VTAIL.n175 VTAIL.n119 0.155672
R613 VTAIL.n168 VTAIL.n119 0.155672
R614 VTAIL.n168 VTAIL.n167 0.155672
R615 VTAIL.n167 VTAIL.n123 0.155672
R616 VTAIL.n160 VTAIL.n123 0.155672
R617 VTAIL.n160 VTAIL.n159 0.155672
R618 VTAIL.n159 VTAIL.n127 0.155672
R619 VTAIL.n152 VTAIL.n127 0.155672
R620 VTAIL.n152 VTAIL.n151 0.155672
R621 VTAIL.n151 VTAIL.n131 0.155672
R622 VTAIL.n144 VTAIL.n131 0.155672
R623 VTAIL.n144 VTAIL.n143 0.155672
R624 VTAIL.n143 VTAIL.n135 0.155672
R625 VDD2.n191 VDD2.n99 289.615
R626 VDD2.n92 VDD2.n0 289.615
R627 VDD2.n192 VDD2.n191 185
R628 VDD2.n190 VDD2.n189 185
R629 VDD2.n103 VDD2.n102 185
R630 VDD2.n184 VDD2.n183 185
R631 VDD2.n182 VDD2.n181 185
R632 VDD2.n107 VDD2.n106 185
R633 VDD2.n111 VDD2.n109 185
R634 VDD2.n176 VDD2.n175 185
R635 VDD2.n174 VDD2.n173 185
R636 VDD2.n113 VDD2.n112 185
R637 VDD2.n168 VDD2.n167 185
R638 VDD2.n166 VDD2.n165 185
R639 VDD2.n117 VDD2.n116 185
R640 VDD2.n160 VDD2.n159 185
R641 VDD2.n158 VDD2.n157 185
R642 VDD2.n121 VDD2.n120 185
R643 VDD2.n152 VDD2.n151 185
R644 VDD2.n150 VDD2.n149 185
R645 VDD2.n125 VDD2.n124 185
R646 VDD2.n144 VDD2.n143 185
R647 VDD2.n142 VDD2.n141 185
R648 VDD2.n129 VDD2.n128 185
R649 VDD2.n136 VDD2.n135 185
R650 VDD2.n134 VDD2.n133 185
R651 VDD2.n33 VDD2.n32 185
R652 VDD2.n35 VDD2.n34 185
R653 VDD2.n28 VDD2.n27 185
R654 VDD2.n41 VDD2.n40 185
R655 VDD2.n43 VDD2.n42 185
R656 VDD2.n24 VDD2.n23 185
R657 VDD2.n49 VDD2.n48 185
R658 VDD2.n51 VDD2.n50 185
R659 VDD2.n20 VDD2.n19 185
R660 VDD2.n57 VDD2.n56 185
R661 VDD2.n59 VDD2.n58 185
R662 VDD2.n16 VDD2.n15 185
R663 VDD2.n65 VDD2.n64 185
R664 VDD2.n67 VDD2.n66 185
R665 VDD2.n12 VDD2.n11 185
R666 VDD2.n74 VDD2.n73 185
R667 VDD2.n75 VDD2.n10 185
R668 VDD2.n77 VDD2.n76 185
R669 VDD2.n8 VDD2.n7 185
R670 VDD2.n83 VDD2.n82 185
R671 VDD2.n85 VDD2.n84 185
R672 VDD2.n4 VDD2.n3 185
R673 VDD2.n91 VDD2.n90 185
R674 VDD2.n93 VDD2.n92 185
R675 VDD2.n132 VDD2.t1 147.659
R676 VDD2.n31 VDD2.t3 147.659
R677 VDD2.n191 VDD2.n190 104.615
R678 VDD2.n190 VDD2.n102 104.615
R679 VDD2.n183 VDD2.n102 104.615
R680 VDD2.n183 VDD2.n182 104.615
R681 VDD2.n182 VDD2.n106 104.615
R682 VDD2.n111 VDD2.n106 104.615
R683 VDD2.n175 VDD2.n111 104.615
R684 VDD2.n175 VDD2.n174 104.615
R685 VDD2.n174 VDD2.n112 104.615
R686 VDD2.n167 VDD2.n112 104.615
R687 VDD2.n167 VDD2.n166 104.615
R688 VDD2.n166 VDD2.n116 104.615
R689 VDD2.n159 VDD2.n116 104.615
R690 VDD2.n159 VDD2.n158 104.615
R691 VDD2.n158 VDD2.n120 104.615
R692 VDD2.n151 VDD2.n120 104.615
R693 VDD2.n151 VDD2.n150 104.615
R694 VDD2.n150 VDD2.n124 104.615
R695 VDD2.n143 VDD2.n124 104.615
R696 VDD2.n143 VDD2.n142 104.615
R697 VDD2.n142 VDD2.n128 104.615
R698 VDD2.n135 VDD2.n128 104.615
R699 VDD2.n135 VDD2.n134 104.615
R700 VDD2.n34 VDD2.n33 104.615
R701 VDD2.n34 VDD2.n27 104.615
R702 VDD2.n41 VDD2.n27 104.615
R703 VDD2.n42 VDD2.n41 104.615
R704 VDD2.n42 VDD2.n23 104.615
R705 VDD2.n49 VDD2.n23 104.615
R706 VDD2.n50 VDD2.n49 104.615
R707 VDD2.n50 VDD2.n19 104.615
R708 VDD2.n57 VDD2.n19 104.615
R709 VDD2.n58 VDD2.n57 104.615
R710 VDD2.n58 VDD2.n15 104.615
R711 VDD2.n65 VDD2.n15 104.615
R712 VDD2.n66 VDD2.n65 104.615
R713 VDD2.n66 VDD2.n11 104.615
R714 VDD2.n74 VDD2.n11 104.615
R715 VDD2.n75 VDD2.n74 104.615
R716 VDD2.n76 VDD2.n75 104.615
R717 VDD2.n76 VDD2.n7 104.615
R718 VDD2.n83 VDD2.n7 104.615
R719 VDD2.n84 VDD2.n83 104.615
R720 VDD2.n84 VDD2.n3 104.615
R721 VDD2.n91 VDD2.n3 104.615
R722 VDD2.n92 VDD2.n91 104.615
R723 VDD2.n98 VDD2.n97 58.8489
R724 VDD2 VDD2.n197 58.846
R725 VDD2.n134 VDD2.t1 52.3082
R726 VDD2.n33 VDD2.t3 52.3082
R727 VDD2.n98 VDD2.n96 47.3543
R728 VDD2.n196 VDD2.n195 46.9247
R729 VDD2.n196 VDD2.n98 40.8338
R730 VDD2.n133 VDD2.n132 15.6677
R731 VDD2.n32 VDD2.n31 15.6677
R732 VDD2.n109 VDD2.n107 13.1884
R733 VDD2.n77 VDD2.n8 13.1884
R734 VDD2.n181 VDD2.n180 12.8005
R735 VDD2.n177 VDD2.n176 12.8005
R736 VDD2.n136 VDD2.n131 12.8005
R737 VDD2.n35 VDD2.n30 12.8005
R738 VDD2.n78 VDD2.n10 12.8005
R739 VDD2.n82 VDD2.n81 12.8005
R740 VDD2.n184 VDD2.n105 12.0247
R741 VDD2.n173 VDD2.n110 12.0247
R742 VDD2.n137 VDD2.n129 12.0247
R743 VDD2.n36 VDD2.n28 12.0247
R744 VDD2.n73 VDD2.n72 12.0247
R745 VDD2.n85 VDD2.n6 12.0247
R746 VDD2.n185 VDD2.n103 11.249
R747 VDD2.n172 VDD2.n113 11.249
R748 VDD2.n141 VDD2.n140 11.249
R749 VDD2.n40 VDD2.n39 11.249
R750 VDD2.n71 VDD2.n12 11.249
R751 VDD2.n86 VDD2.n4 11.249
R752 VDD2.n189 VDD2.n188 10.4732
R753 VDD2.n169 VDD2.n168 10.4732
R754 VDD2.n144 VDD2.n127 10.4732
R755 VDD2.n43 VDD2.n26 10.4732
R756 VDD2.n68 VDD2.n67 10.4732
R757 VDD2.n90 VDD2.n89 10.4732
R758 VDD2.n192 VDD2.n101 9.69747
R759 VDD2.n165 VDD2.n115 9.69747
R760 VDD2.n145 VDD2.n125 9.69747
R761 VDD2.n44 VDD2.n24 9.69747
R762 VDD2.n64 VDD2.n14 9.69747
R763 VDD2.n93 VDD2.n2 9.69747
R764 VDD2.n195 VDD2.n194 9.45567
R765 VDD2.n96 VDD2.n95 9.45567
R766 VDD2.n119 VDD2.n118 9.3005
R767 VDD2.n162 VDD2.n161 9.3005
R768 VDD2.n164 VDD2.n163 9.3005
R769 VDD2.n115 VDD2.n114 9.3005
R770 VDD2.n170 VDD2.n169 9.3005
R771 VDD2.n172 VDD2.n171 9.3005
R772 VDD2.n110 VDD2.n108 9.3005
R773 VDD2.n178 VDD2.n177 9.3005
R774 VDD2.n194 VDD2.n193 9.3005
R775 VDD2.n101 VDD2.n100 9.3005
R776 VDD2.n188 VDD2.n187 9.3005
R777 VDD2.n186 VDD2.n185 9.3005
R778 VDD2.n105 VDD2.n104 9.3005
R779 VDD2.n180 VDD2.n179 9.3005
R780 VDD2.n156 VDD2.n155 9.3005
R781 VDD2.n154 VDD2.n153 9.3005
R782 VDD2.n123 VDD2.n122 9.3005
R783 VDD2.n148 VDD2.n147 9.3005
R784 VDD2.n146 VDD2.n145 9.3005
R785 VDD2.n127 VDD2.n126 9.3005
R786 VDD2.n140 VDD2.n139 9.3005
R787 VDD2.n138 VDD2.n137 9.3005
R788 VDD2.n131 VDD2.n130 9.3005
R789 VDD2.n95 VDD2.n94 9.3005
R790 VDD2.n2 VDD2.n1 9.3005
R791 VDD2.n89 VDD2.n88 9.3005
R792 VDD2.n87 VDD2.n86 9.3005
R793 VDD2.n6 VDD2.n5 9.3005
R794 VDD2.n81 VDD2.n80 9.3005
R795 VDD2.n53 VDD2.n52 9.3005
R796 VDD2.n22 VDD2.n21 9.3005
R797 VDD2.n47 VDD2.n46 9.3005
R798 VDD2.n45 VDD2.n44 9.3005
R799 VDD2.n26 VDD2.n25 9.3005
R800 VDD2.n39 VDD2.n38 9.3005
R801 VDD2.n37 VDD2.n36 9.3005
R802 VDD2.n30 VDD2.n29 9.3005
R803 VDD2.n55 VDD2.n54 9.3005
R804 VDD2.n18 VDD2.n17 9.3005
R805 VDD2.n61 VDD2.n60 9.3005
R806 VDD2.n63 VDD2.n62 9.3005
R807 VDD2.n14 VDD2.n13 9.3005
R808 VDD2.n69 VDD2.n68 9.3005
R809 VDD2.n71 VDD2.n70 9.3005
R810 VDD2.n72 VDD2.n9 9.3005
R811 VDD2.n79 VDD2.n78 9.3005
R812 VDD2.n193 VDD2.n99 8.92171
R813 VDD2.n164 VDD2.n117 8.92171
R814 VDD2.n149 VDD2.n148 8.92171
R815 VDD2.n48 VDD2.n47 8.92171
R816 VDD2.n63 VDD2.n16 8.92171
R817 VDD2.n94 VDD2.n0 8.92171
R818 VDD2.n161 VDD2.n160 8.14595
R819 VDD2.n152 VDD2.n123 8.14595
R820 VDD2.n51 VDD2.n22 8.14595
R821 VDD2.n60 VDD2.n59 8.14595
R822 VDD2.n157 VDD2.n119 7.3702
R823 VDD2.n153 VDD2.n121 7.3702
R824 VDD2.n52 VDD2.n20 7.3702
R825 VDD2.n56 VDD2.n18 7.3702
R826 VDD2.n157 VDD2.n156 6.59444
R827 VDD2.n156 VDD2.n121 6.59444
R828 VDD2.n55 VDD2.n20 6.59444
R829 VDD2.n56 VDD2.n55 6.59444
R830 VDD2.n160 VDD2.n119 5.81868
R831 VDD2.n153 VDD2.n152 5.81868
R832 VDD2.n52 VDD2.n51 5.81868
R833 VDD2.n59 VDD2.n18 5.81868
R834 VDD2.n195 VDD2.n99 5.04292
R835 VDD2.n161 VDD2.n117 5.04292
R836 VDD2.n149 VDD2.n123 5.04292
R837 VDD2.n48 VDD2.n22 5.04292
R838 VDD2.n60 VDD2.n16 5.04292
R839 VDD2.n96 VDD2.n0 5.04292
R840 VDD2.n132 VDD2.n130 4.38563
R841 VDD2.n31 VDD2.n29 4.38563
R842 VDD2.n193 VDD2.n192 4.26717
R843 VDD2.n165 VDD2.n164 4.26717
R844 VDD2.n148 VDD2.n125 4.26717
R845 VDD2.n47 VDD2.n24 4.26717
R846 VDD2.n64 VDD2.n63 4.26717
R847 VDD2.n94 VDD2.n93 4.26717
R848 VDD2.n189 VDD2.n101 3.49141
R849 VDD2.n168 VDD2.n115 3.49141
R850 VDD2.n145 VDD2.n144 3.49141
R851 VDD2.n44 VDD2.n43 3.49141
R852 VDD2.n67 VDD2.n14 3.49141
R853 VDD2.n90 VDD2.n2 3.49141
R854 VDD2.n188 VDD2.n103 2.71565
R855 VDD2.n169 VDD2.n113 2.71565
R856 VDD2.n141 VDD2.n127 2.71565
R857 VDD2.n40 VDD2.n26 2.71565
R858 VDD2.n68 VDD2.n12 2.71565
R859 VDD2.n89 VDD2.n4 2.71565
R860 VDD2.n185 VDD2.n184 1.93989
R861 VDD2.n173 VDD2.n172 1.93989
R862 VDD2.n140 VDD2.n129 1.93989
R863 VDD2.n39 VDD2.n28 1.93989
R864 VDD2.n73 VDD2.n71 1.93989
R865 VDD2.n86 VDD2.n85 1.93989
R866 VDD2.n181 VDD2.n105 1.16414
R867 VDD2.n176 VDD2.n110 1.16414
R868 VDD2.n137 VDD2.n136 1.16414
R869 VDD2.n36 VDD2.n35 1.16414
R870 VDD2.n72 VDD2.n10 1.16414
R871 VDD2.n82 VDD2.n6 1.16414
R872 VDD2.n197 VDD2.t4 1.13712
R873 VDD2.n197 VDD2.t2 1.13712
R874 VDD2.n97 VDD2.t0 1.13712
R875 VDD2.n97 VDD2.t5 1.13712
R876 VDD2 VDD2.n196 0.543603
R877 VDD2.n180 VDD2.n107 0.388379
R878 VDD2.n177 VDD2.n109 0.388379
R879 VDD2.n133 VDD2.n131 0.388379
R880 VDD2.n32 VDD2.n30 0.388379
R881 VDD2.n78 VDD2.n77 0.388379
R882 VDD2.n81 VDD2.n8 0.388379
R883 VDD2.n194 VDD2.n100 0.155672
R884 VDD2.n187 VDD2.n100 0.155672
R885 VDD2.n187 VDD2.n186 0.155672
R886 VDD2.n186 VDD2.n104 0.155672
R887 VDD2.n179 VDD2.n104 0.155672
R888 VDD2.n179 VDD2.n178 0.155672
R889 VDD2.n178 VDD2.n108 0.155672
R890 VDD2.n171 VDD2.n108 0.155672
R891 VDD2.n171 VDD2.n170 0.155672
R892 VDD2.n170 VDD2.n114 0.155672
R893 VDD2.n163 VDD2.n114 0.155672
R894 VDD2.n163 VDD2.n162 0.155672
R895 VDD2.n162 VDD2.n118 0.155672
R896 VDD2.n155 VDD2.n118 0.155672
R897 VDD2.n155 VDD2.n154 0.155672
R898 VDD2.n154 VDD2.n122 0.155672
R899 VDD2.n147 VDD2.n122 0.155672
R900 VDD2.n147 VDD2.n146 0.155672
R901 VDD2.n146 VDD2.n126 0.155672
R902 VDD2.n139 VDD2.n126 0.155672
R903 VDD2.n139 VDD2.n138 0.155672
R904 VDD2.n138 VDD2.n130 0.155672
R905 VDD2.n37 VDD2.n29 0.155672
R906 VDD2.n38 VDD2.n37 0.155672
R907 VDD2.n38 VDD2.n25 0.155672
R908 VDD2.n45 VDD2.n25 0.155672
R909 VDD2.n46 VDD2.n45 0.155672
R910 VDD2.n46 VDD2.n21 0.155672
R911 VDD2.n53 VDD2.n21 0.155672
R912 VDD2.n54 VDD2.n53 0.155672
R913 VDD2.n54 VDD2.n17 0.155672
R914 VDD2.n61 VDD2.n17 0.155672
R915 VDD2.n62 VDD2.n61 0.155672
R916 VDD2.n62 VDD2.n13 0.155672
R917 VDD2.n69 VDD2.n13 0.155672
R918 VDD2.n70 VDD2.n69 0.155672
R919 VDD2.n70 VDD2.n9 0.155672
R920 VDD2.n79 VDD2.n9 0.155672
R921 VDD2.n80 VDD2.n79 0.155672
R922 VDD2.n80 VDD2.n5 0.155672
R923 VDD2.n87 VDD2.n5 0.155672
R924 VDD2.n88 VDD2.n87 0.155672
R925 VDD2.n88 VDD2.n1 0.155672
R926 VDD2.n95 VDD2.n1 0.155672
R927 B.n448 B.t17 1208.28
R928 B.n446 B.t6 1208.28
R929 B.n100 B.t14 1208.28
R930 B.n98 B.t10 1208.28
R931 B.n775 B.n774 585
R932 B.n776 B.n775 585
R933 B.n350 B.n97 585
R934 B.n349 B.n348 585
R935 B.n347 B.n346 585
R936 B.n345 B.n344 585
R937 B.n343 B.n342 585
R938 B.n341 B.n340 585
R939 B.n339 B.n338 585
R940 B.n337 B.n336 585
R941 B.n335 B.n334 585
R942 B.n333 B.n332 585
R943 B.n331 B.n330 585
R944 B.n329 B.n328 585
R945 B.n327 B.n326 585
R946 B.n325 B.n324 585
R947 B.n323 B.n322 585
R948 B.n321 B.n320 585
R949 B.n319 B.n318 585
R950 B.n317 B.n316 585
R951 B.n315 B.n314 585
R952 B.n313 B.n312 585
R953 B.n311 B.n310 585
R954 B.n309 B.n308 585
R955 B.n307 B.n306 585
R956 B.n305 B.n304 585
R957 B.n303 B.n302 585
R958 B.n301 B.n300 585
R959 B.n299 B.n298 585
R960 B.n297 B.n296 585
R961 B.n295 B.n294 585
R962 B.n293 B.n292 585
R963 B.n291 B.n290 585
R964 B.n289 B.n288 585
R965 B.n287 B.n286 585
R966 B.n285 B.n284 585
R967 B.n283 B.n282 585
R968 B.n281 B.n280 585
R969 B.n279 B.n278 585
R970 B.n277 B.n276 585
R971 B.n275 B.n274 585
R972 B.n273 B.n272 585
R973 B.n271 B.n270 585
R974 B.n269 B.n268 585
R975 B.n267 B.n266 585
R976 B.n265 B.n264 585
R977 B.n263 B.n262 585
R978 B.n261 B.n260 585
R979 B.n259 B.n258 585
R980 B.n257 B.n256 585
R981 B.n255 B.n254 585
R982 B.n253 B.n252 585
R983 B.n251 B.n250 585
R984 B.n249 B.n248 585
R985 B.n247 B.n246 585
R986 B.n245 B.n244 585
R987 B.n243 B.n242 585
R988 B.n241 B.n240 585
R989 B.n239 B.n238 585
R990 B.n236 B.n235 585
R991 B.n234 B.n233 585
R992 B.n232 B.n231 585
R993 B.n230 B.n229 585
R994 B.n228 B.n227 585
R995 B.n226 B.n225 585
R996 B.n224 B.n223 585
R997 B.n222 B.n221 585
R998 B.n220 B.n219 585
R999 B.n218 B.n217 585
R1000 B.n216 B.n215 585
R1001 B.n214 B.n213 585
R1002 B.n212 B.n211 585
R1003 B.n210 B.n209 585
R1004 B.n208 B.n207 585
R1005 B.n206 B.n205 585
R1006 B.n204 B.n203 585
R1007 B.n202 B.n201 585
R1008 B.n200 B.n199 585
R1009 B.n198 B.n197 585
R1010 B.n196 B.n195 585
R1011 B.n194 B.n193 585
R1012 B.n192 B.n191 585
R1013 B.n190 B.n189 585
R1014 B.n188 B.n187 585
R1015 B.n186 B.n185 585
R1016 B.n184 B.n183 585
R1017 B.n182 B.n181 585
R1018 B.n180 B.n179 585
R1019 B.n178 B.n177 585
R1020 B.n176 B.n175 585
R1021 B.n174 B.n173 585
R1022 B.n172 B.n171 585
R1023 B.n170 B.n169 585
R1024 B.n168 B.n167 585
R1025 B.n166 B.n165 585
R1026 B.n164 B.n163 585
R1027 B.n162 B.n161 585
R1028 B.n160 B.n159 585
R1029 B.n158 B.n157 585
R1030 B.n156 B.n155 585
R1031 B.n154 B.n153 585
R1032 B.n152 B.n151 585
R1033 B.n150 B.n149 585
R1034 B.n148 B.n147 585
R1035 B.n146 B.n145 585
R1036 B.n144 B.n143 585
R1037 B.n142 B.n141 585
R1038 B.n140 B.n139 585
R1039 B.n138 B.n137 585
R1040 B.n136 B.n135 585
R1041 B.n134 B.n133 585
R1042 B.n132 B.n131 585
R1043 B.n130 B.n129 585
R1044 B.n128 B.n127 585
R1045 B.n126 B.n125 585
R1046 B.n124 B.n123 585
R1047 B.n122 B.n121 585
R1048 B.n120 B.n119 585
R1049 B.n118 B.n117 585
R1050 B.n116 B.n115 585
R1051 B.n114 B.n113 585
R1052 B.n112 B.n111 585
R1053 B.n110 B.n109 585
R1054 B.n108 B.n107 585
R1055 B.n106 B.n105 585
R1056 B.n104 B.n103 585
R1057 B.n773 B.n34 585
R1058 B.n777 B.n34 585
R1059 B.n772 B.n33 585
R1060 B.n778 B.n33 585
R1061 B.n771 B.n770 585
R1062 B.n770 B.n29 585
R1063 B.n769 B.n28 585
R1064 B.n784 B.n28 585
R1065 B.n768 B.n27 585
R1066 B.n785 B.n27 585
R1067 B.n767 B.n26 585
R1068 B.n786 B.n26 585
R1069 B.n766 B.n765 585
R1070 B.n765 B.n22 585
R1071 B.n764 B.n21 585
R1072 B.n792 B.n21 585
R1073 B.n763 B.n20 585
R1074 B.n793 B.n20 585
R1075 B.n762 B.n19 585
R1076 B.n794 B.n19 585
R1077 B.n761 B.n760 585
R1078 B.n760 B.n15 585
R1079 B.n759 B.n14 585
R1080 B.n800 B.n14 585
R1081 B.n758 B.n13 585
R1082 B.n801 B.n13 585
R1083 B.n757 B.n12 585
R1084 B.n802 B.n12 585
R1085 B.n756 B.n755 585
R1086 B.n755 B.n11 585
R1087 B.n754 B.n7 585
R1088 B.n808 B.n7 585
R1089 B.n753 B.n6 585
R1090 B.n809 B.n6 585
R1091 B.n752 B.n5 585
R1092 B.n810 B.n5 585
R1093 B.n751 B.n750 585
R1094 B.n750 B.n4 585
R1095 B.n749 B.n351 585
R1096 B.n749 B.n748 585
R1097 B.n738 B.n352 585
R1098 B.n741 B.n352 585
R1099 B.n740 B.n739 585
R1100 B.n742 B.n740 585
R1101 B.n737 B.n356 585
R1102 B.n360 B.n356 585
R1103 B.n736 B.n735 585
R1104 B.n735 B.n734 585
R1105 B.n358 B.n357 585
R1106 B.n359 B.n358 585
R1107 B.n727 B.n726 585
R1108 B.n728 B.n727 585
R1109 B.n725 B.n365 585
R1110 B.n365 B.n364 585
R1111 B.n724 B.n723 585
R1112 B.n723 B.n722 585
R1113 B.n367 B.n366 585
R1114 B.n368 B.n367 585
R1115 B.n715 B.n714 585
R1116 B.n716 B.n715 585
R1117 B.n713 B.n372 585
R1118 B.n376 B.n372 585
R1119 B.n712 B.n711 585
R1120 B.n711 B.n710 585
R1121 B.n374 B.n373 585
R1122 B.n375 B.n374 585
R1123 B.n703 B.n702 585
R1124 B.n704 B.n703 585
R1125 B.n701 B.n381 585
R1126 B.n381 B.n380 585
R1127 B.n695 B.n694 585
R1128 B.n693 B.n445 585
R1129 B.n692 B.n444 585
R1130 B.n697 B.n444 585
R1131 B.n691 B.n690 585
R1132 B.n689 B.n688 585
R1133 B.n687 B.n686 585
R1134 B.n685 B.n684 585
R1135 B.n683 B.n682 585
R1136 B.n681 B.n680 585
R1137 B.n679 B.n678 585
R1138 B.n677 B.n676 585
R1139 B.n675 B.n674 585
R1140 B.n673 B.n672 585
R1141 B.n671 B.n670 585
R1142 B.n669 B.n668 585
R1143 B.n667 B.n666 585
R1144 B.n665 B.n664 585
R1145 B.n663 B.n662 585
R1146 B.n661 B.n660 585
R1147 B.n659 B.n658 585
R1148 B.n657 B.n656 585
R1149 B.n655 B.n654 585
R1150 B.n653 B.n652 585
R1151 B.n651 B.n650 585
R1152 B.n649 B.n648 585
R1153 B.n647 B.n646 585
R1154 B.n645 B.n644 585
R1155 B.n643 B.n642 585
R1156 B.n641 B.n640 585
R1157 B.n639 B.n638 585
R1158 B.n637 B.n636 585
R1159 B.n635 B.n634 585
R1160 B.n633 B.n632 585
R1161 B.n631 B.n630 585
R1162 B.n629 B.n628 585
R1163 B.n627 B.n626 585
R1164 B.n625 B.n624 585
R1165 B.n623 B.n622 585
R1166 B.n621 B.n620 585
R1167 B.n619 B.n618 585
R1168 B.n617 B.n616 585
R1169 B.n615 B.n614 585
R1170 B.n613 B.n612 585
R1171 B.n611 B.n610 585
R1172 B.n609 B.n608 585
R1173 B.n607 B.n606 585
R1174 B.n605 B.n604 585
R1175 B.n603 B.n602 585
R1176 B.n601 B.n600 585
R1177 B.n599 B.n598 585
R1178 B.n597 B.n596 585
R1179 B.n595 B.n594 585
R1180 B.n593 B.n592 585
R1181 B.n591 B.n590 585
R1182 B.n589 B.n588 585
R1183 B.n587 B.n586 585
R1184 B.n585 B.n584 585
R1185 B.n583 B.n582 585
R1186 B.n580 B.n579 585
R1187 B.n578 B.n577 585
R1188 B.n576 B.n575 585
R1189 B.n574 B.n573 585
R1190 B.n572 B.n571 585
R1191 B.n570 B.n569 585
R1192 B.n568 B.n567 585
R1193 B.n566 B.n565 585
R1194 B.n564 B.n563 585
R1195 B.n562 B.n561 585
R1196 B.n560 B.n559 585
R1197 B.n558 B.n557 585
R1198 B.n556 B.n555 585
R1199 B.n554 B.n553 585
R1200 B.n552 B.n551 585
R1201 B.n550 B.n549 585
R1202 B.n548 B.n547 585
R1203 B.n546 B.n545 585
R1204 B.n544 B.n543 585
R1205 B.n542 B.n541 585
R1206 B.n540 B.n539 585
R1207 B.n538 B.n537 585
R1208 B.n536 B.n535 585
R1209 B.n534 B.n533 585
R1210 B.n532 B.n531 585
R1211 B.n530 B.n529 585
R1212 B.n528 B.n527 585
R1213 B.n526 B.n525 585
R1214 B.n524 B.n523 585
R1215 B.n522 B.n521 585
R1216 B.n520 B.n519 585
R1217 B.n518 B.n517 585
R1218 B.n516 B.n515 585
R1219 B.n514 B.n513 585
R1220 B.n512 B.n511 585
R1221 B.n510 B.n509 585
R1222 B.n508 B.n507 585
R1223 B.n506 B.n505 585
R1224 B.n504 B.n503 585
R1225 B.n502 B.n501 585
R1226 B.n500 B.n499 585
R1227 B.n498 B.n497 585
R1228 B.n496 B.n495 585
R1229 B.n494 B.n493 585
R1230 B.n492 B.n491 585
R1231 B.n490 B.n489 585
R1232 B.n488 B.n487 585
R1233 B.n486 B.n485 585
R1234 B.n484 B.n483 585
R1235 B.n482 B.n481 585
R1236 B.n480 B.n479 585
R1237 B.n478 B.n477 585
R1238 B.n476 B.n475 585
R1239 B.n474 B.n473 585
R1240 B.n472 B.n471 585
R1241 B.n470 B.n469 585
R1242 B.n468 B.n467 585
R1243 B.n466 B.n465 585
R1244 B.n464 B.n463 585
R1245 B.n462 B.n461 585
R1246 B.n460 B.n459 585
R1247 B.n458 B.n457 585
R1248 B.n456 B.n455 585
R1249 B.n454 B.n453 585
R1250 B.n452 B.n451 585
R1251 B.n383 B.n382 585
R1252 B.n700 B.n699 585
R1253 B.n379 B.n378 585
R1254 B.n380 B.n379 585
R1255 B.n706 B.n705 585
R1256 B.n705 B.n704 585
R1257 B.n707 B.n377 585
R1258 B.n377 B.n375 585
R1259 B.n709 B.n708 585
R1260 B.n710 B.n709 585
R1261 B.n371 B.n370 585
R1262 B.n376 B.n371 585
R1263 B.n718 B.n717 585
R1264 B.n717 B.n716 585
R1265 B.n719 B.n369 585
R1266 B.n369 B.n368 585
R1267 B.n721 B.n720 585
R1268 B.n722 B.n721 585
R1269 B.n363 B.n362 585
R1270 B.n364 B.n363 585
R1271 B.n730 B.n729 585
R1272 B.n729 B.n728 585
R1273 B.n731 B.n361 585
R1274 B.n361 B.n359 585
R1275 B.n733 B.n732 585
R1276 B.n734 B.n733 585
R1277 B.n355 B.n354 585
R1278 B.n360 B.n355 585
R1279 B.n744 B.n743 585
R1280 B.n743 B.n742 585
R1281 B.n745 B.n353 585
R1282 B.n741 B.n353 585
R1283 B.n747 B.n746 585
R1284 B.n748 B.n747 585
R1285 B.n2 B.n0 585
R1286 B.n4 B.n2 585
R1287 B.n3 B.n1 585
R1288 B.n809 B.n3 585
R1289 B.n807 B.n806 585
R1290 B.n808 B.n807 585
R1291 B.n805 B.n8 585
R1292 B.n11 B.n8 585
R1293 B.n804 B.n803 585
R1294 B.n803 B.n802 585
R1295 B.n10 B.n9 585
R1296 B.n801 B.n10 585
R1297 B.n799 B.n798 585
R1298 B.n800 B.n799 585
R1299 B.n797 B.n16 585
R1300 B.n16 B.n15 585
R1301 B.n796 B.n795 585
R1302 B.n795 B.n794 585
R1303 B.n18 B.n17 585
R1304 B.n793 B.n18 585
R1305 B.n791 B.n790 585
R1306 B.n792 B.n791 585
R1307 B.n789 B.n23 585
R1308 B.n23 B.n22 585
R1309 B.n788 B.n787 585
R1310 B.n787 B.n786 585
R1311 B.n25 B.n24 585
R1312 B.n785 B.n25 585
R1313 B.n783 B.n782 585
R1314 B.n784 B.n783 585
R1315 B.n781 B.n30 585
R1316 B.n30 B.n29 585
R1317 B.n780 B.n779 585
R1318 B.n779 B.n778 585
R1319 B.n32 B.n31 585
R1320 B.n777 B.n32 585
R1321 B.n812 B.n811 585
R1322 B.n811 B.n810 585
R1323 B.n695 B.n379 463.671
R1324 B.n103 B.n32 463.671
R1325 B.n699 B.n381 463.671
R1326 B.n775 B.n34 463.671
R1327 B.n448 B.t19 389.865
R1328 B.n98 B.t12 389.865
R1329 B.n446 B.t9 389.865
R1330 B.n100 B.t15 389.865
R1331 B.n449 B.t18 375.32
R1332 B.n99 B.t13 375.32
R1333 B.n447 B.t8 375.32
R1334 B.n101 B.t16 375.32
R1335 B.n776 B.n96 256.663
R1336 B.n776 B.n95 256.663
R1337 B.n776 B.n94 256.663
R1338 B.n776 B.n93 256.663
R1339 B.n776 B.n92 256.663
R1340 B.n776 B.n91 256.663
R1341 B.n776 B.n90 256.663
R1342 B.n776 B.n89 256.663
R1343 B.n776 B.n88 256.663
R1344 B.n776 B.n87 256.663
R1345 B.n776 B.n86 256.663
R1346 B.n776 B.n85 256.663
R1347 B.n776 B.n84 256.663
R1348 B.n776 B.n83 256.663
R1349 B.n776 B.n82 256.663
R1350 B.n776 B.n81 256.663
R1351 B.n776 B.n80 256.663
R1352 B.n776 B.n79 256.663
R1353 B.n776 B.n78 256.663
R1354 B.n776 B.n77 256.663
R1355 B.n776 B.n76 256.663
R1356 B.n776 B.n75 256.663
R1357 B.n776 B.n74 256.663
R1358 B.n776 B.n73 256.663
R1359 B.n776 B.n72 256.663
R1360 B.n776 B.n71 256.663
R1361 B.n776 B.n70 256.663
R1362 B.n776 B.n69 256.663
R1363 B.n776 B.n68 256.663
R1364 B.n776 B.n67 256.663
R1365 B.n776 B.n66 256.663
R1366 B.n776 B.n65 256.663
R1367 B.n776 B.n64 256.663
R1368 B.n776 B.n63 256.663
R1369 B.n776 B.n62 256.663
R1370 B.n776 B.n61 256.663
R1371 B.n776 B.n60 256.663
R1372 B.n776 B.n59 256.663
R1373 B.n776 B.n58 256.663
R1374 B.n776 B.n57 256.663
R1375 B.n776 B.n56 256.663
R1376 B.n776 B.n55 256.663
R1377 B.n776 B.n54 256.663
R1378 B.n776 B.n53 256.663
R1379 B.n776 B.n52 256.663
R1380 B.n776 B.n51 256.663
R1381 B.n776 B.n50 256.663
R1382 B.n776 B.n49 256.663
R1383 B.n776 B.n48 256.663
R1384 B.n776 B.n47 256.663
R1385 B.n776 B.n46 256.663
R1386 B.n776 B.n45 256.663
R1387 B.n776 B.n44 256.663
R1388 B.n776 B.n43 256.663
R1389 B.n776 B.n42 256.663
R1390 B.n776 B.n41 256.663
R1391 B.n776 B.n40 256.663
R1392 B.n776 B.n39 256.663
R1393 B.n776 B.n38 256.663
R1394 B.n776 B.n37 256.663
R1395 B.n776 B.n36 256.663
R1396 B.n776 B.n35 256.663
R1397 B.n697 B.n696 256.663
R1398 B.n697 B.n384 256.663
R1399 B.n697 B.n385 256.663
R1400 B.n697 B.n386 256.663
R1401 B.n697 B.n387 256.663
R1402 B.n697 B.n388 256.663
R1403 B.n697 B.n389 256.663
R1404 B.n697 B.n390 256.663
R1405 B.n697 B.n391 256.663
R1406 B.n697 B.n392 256.663
R1407 B.n697 B.n393 256.663
R1408 B.n697 B.n394 256.663
R1409 B.n697 B.n395 256.663
R1410 B.n697 B.n396 256.663
R1411 B.n697 B.n397 256.663
R1412 B.n697 B.n398 256.663
R1413 B.n697 B.n399 256.663
R1414 B.n697 B.n400 256.663
R1415 B.n697 B.n401 256.663
R1416 B.n697 B.n402 256.663
R1417 B.n697 B.n403 256.663
R1418 B.n697 B.n404 256.663
R1419 B.n697 B.n405 256.663
R1420 B.n697 B.n406 256.663
R1421 B.n697 B.n407 256.663
R1422 B.n697 B.n408 256.663
R1423 B.n697 B.n409 256.663
R1424 B.n697 B.n410 256.663
R1425 B.n697 B.n411 256.663
R1426 B.n697 B.n412 256.663
R1427 B.n697 B.n413 256.663
R1428 B.n697 B.n414 256.663
R1429 B.n697 B.n415 256.663
R1430 B.n697 B.n416 256.663
R1431 B.n697 B.n417 256.663
R1432 B.n697 B.n418 256.663
R1433 B.n697 B.n419 256.663
R1434 B.n697 B.n420 256.663
R1435 B.n697 B.n421 256.663
R1436 B.n697 B.n422 256.663
R1437 B.n697 B.n423 256.663
R1438 B.n697 B.n424 256.663
R1439 B.n697 B.n425 256.663
R1440 B.n697 B.n426 256.663
R1441 B.n697 B.n427 256.663
R1442 B.n697 B.n428 256.663
R1443 B.n697 B.n429 256.663
R1444 B.n697 B.n430 256.663
R1445 B.n697 B.n431 256.663
R1446 B.n697 B.n432 256.663
R1447 B.n697 B.n433 256.663
R1448 B.n697 B.n434 256.663
R1449 B.n697 B.n435 256.663
R1450 B.n697 B.n436 256.663
R1451 B.n697 B.n437 256.663
R1452 B.n697 B.n438 256.663
R1453 B.n697 B.n439 256.663
R1454 B.n697 B.n440 256.663
R1455 B.n697 B.n441 256.663
R1456 B.n697 B.n442 256.663
R1457 B.n697 B.n443 256.663
R1458 B.n698 B.n697 256.663
R1459 B.n705 B.n379 163.367
R1460 B.n705 B.n377 163.367
R1461 B.n709 B.n377 163.367
R1462 B.n709 B.n371 163.367
R1463 B.n717 B.n371 163.367
R1464 B.n717 B.n369 163.367
R1465 B.n721 B.n369 163.367
R1466 B.n721 B.n363 163.367
R1467 B.n729 B.n363 163.367
R1468 B.n729 B.n361 163.367
R1469 B.n733 B.n361 163.367
R1470 B.n733 B.n355 163.367
R1471 B.n743 B.n355 163.367
R1472 B.n743 B.n353 163.367
R1473 B.n747 B.n353 163.367
R1474 B.n747 B.n2 163.367
R1475 B.n811 B.n2 163.367
R1476 B.n811 B.n3 163.367
R1477 B.n807 B.n3 163.367
R1478 B.n807 B.n8 163.367
R1479 B.n803 B.n8 163.367
R1480 B.n803 B.n10 163.367
R1481 B.n799 B.n10 163.367
R1482 B.n799 B.n16 163.367
R1483 B.n795 B.n16 163.367
R1484 B.n795 B.n18 163.367
R1485 B.n791 B.n18 163.367
R1486 B.n791 B.n23 163.367
R1487 B.n787 B.n23 163.367
R1488 B.n787 B.n25 163.367
R1489 B.n783 B.n25 163.367
R1490 B.n783 B.n30 163.367
R1491 B.n779 B.n30 163.367
R1492 B.n779 B.n32 163.367
R1493 B.n445 B.n444 163.367
R1494 B.n690 B.n444 163.367
R1495 B.n688 B.n687 163.367
R1496 B.n684 B.n683 163.367
R1497 B.n680 B.n679 163.367
R1498 B.n676 B.n675 163.367
R1499 B.n672 B.n671 163.367
R1500 B.n668 B.n667 163.367
R1501 B.n664 B.n663 163.367
R1502 B.n660 B.n659 163.367
R1503 B.n656 B.n655 163.367
R1504 B.n652 B.n651 163.367
R1505 B.n648 B.n647 163.367
R1506 B.n644 B.n643 163.367
R1507 B.n640 B.n639 163.367
R1508 B.n636 B.n635 163.367
R1509 B.n632 B.n631 163.367
R1510 B.n628 B.n627 163.367
R1511 B.n624 B.n623 163.367
R1512 B.n620 B.n619 163.367
R1513 B.n616 B.n615 163.367
R1514 B.n612 B.n611 163.367
R1515 B.n608 B.n607 163.367
R1516 B.n604 B.n603 163.367
R1517 B.n600 B.n599 163.367
R1518 B.n596 B.n595 163.367
R1519 B.n592 B.n591 163.367
R1520 B.n588 B.n587 163.367
R1521 B.n584 B.n583 163.367
R1522 B.n579 B.n578 163.367
R1523 B.n575 B.n574 163.367
R1524 B.n571 B.n570 163.367
R1525 B.n567 B.n566 163.367
R1526 B.n563 B.n562 163.367
R1527 B.n559 B.n558 163.367
R1528 B.n555 B.n554 163.367
R1529 B.n551 B.n550 163.367
R1530 B.n547 B.n546 163.367
R1531 B.n543 B.n542 163.367
R1532 B.n539 B.n538 163.367
R1533 B.n535 B.n534 163.367
R1534 B.n531 B.n530 163.367
R1535 B.n527 B.n526 163.367
R1536 B.n523 B.n522 163.367
R1537 B.n519 B.n518 163.367
R1538 B.n515 B.n514 163.367
R1539 B.n511 B.n510 163.367
R1540 B.n507 B.n506 163.367
R1541 B.n503 B.n502 163.367
R1542 B.n499 B.n498 163.367
R1543 B.n495 B.n494 163.367
R1544 B.n491 B.n490 163.367
R1545 B.n487 B.n486 163.367
R1546 B.n483 B.n482 163.367
R1547 B.n479 B.n478 163.367
R1548 B.n475 B.n474 163.367
R1549 B.n471 B.n470 163.367
R1550 B.n467 B.n466 163.367
R1551 B.n463 B.n462 163.367
R1552 B.n459 B.n458 163.367
R1553 B.n455 B.n454 163.367
R1554 B.n451 B.n383 163.367
R1555 B.n703 B.n381 163.367
R1556 B.n703 B.n374 163.367
R1557 B.n711 B.n374 163.367
R1558 B.n711 B.n372 163.367
R1559 B.n715 B.n372 163.367
R1560 B.n715 B.n367 163.367
R1561 B.n723 B.n367 163.367
R1562 B.n723 B.n365 163.367
R1563 B.n727 B.n365 163.367
R1564 B.n727 B.n358 163.367
R1565 B.n735 B.n358 163.367
R1566 B.n735 B.n356 163.367
R1567 B.n740 B.n356 163.367
R1568 B.n740 B.n352 163.367
R1569 B.n749 B.n352 163.367
R1570 B.n750 B.n749 163.367
R1571 B.n750 B.n5 163.367
R1572 B.n6 B.n5 163.367
R1573 B.n7 B.n6 163.367
R1574 B.n755 B.n7 163.367
R1575 B.n755 B.n12 163.367
R1576 B.n13 B.n12 163.367
R1577 B.n14 B.n13 163.367
R1578 B.n760 B.n14 163.367
R1579 B.n760 B.n19 163.367
R1580 B.n20 B.n19 163.367
R1581 B.n21 B.n20 163.367
R1582 B.n765 B.n21 163.367
R1583 B.n765 B.n26 163.367
R1584 B.n27 B.n26 163.367
R1585 B.n28 B.n27 163.367
R1586 B.n770 B.n28 163.367
R1587 B.n770 B.n33 163.367
R1588 B.n34 B.n33 163.367
R1589 B.n107 B.n106 163.367
R1590 B.n111 B.n110 163.367
R1591 B.n115 B.n114 163.367
R1592 B.n119 B.n118 163.367
R1593 B.n123 B.n122 163.367
R1594 B.n127 B.n126 163.367
R1595 B.n131 B.n130 163.367
R1596 B.n135 B.n134 163.367
R1597 B.n139 B.n138 163.367
R1598 B.n143 B.n142 163.367
R1599 B.n147 B.n146 163.367
R1600 B.n151 B.n150 163.367
R1601 B.n155 B.n154 163.367
R1602 B.n159 B.n158 163.367
R1603 B.n163 B.n162 163.367
R1604 B.n167 B.n166 163.367
R1605 B.n171 B.n170 163.367
R1606 B.n175 B.n174 163.367
R1607 B.n179 B.n178 163.367
R1608 B.n183 B.n182 163.367
R1609 B.n187 B.n186 163.367
R1610 B.n191 B.n190 163.367
R1611 B.n195 B.n194 163.367
R1612 B.n199 B.n198 163.367
R1613 B.n203 B.n202 163.367
R1614 B.n207 B.n206 163.367
R1615 B.n211 B.n210 163.367
R1616 B.n215 B.n214 163.367
R1617 B.n219 B.n218 163.367
R1618 B.n223 B.n222 163.367
R1619 B.n227 B.n226 163.367
R1620 B.n231 B.n230 163.367
R1621 B.n235 B.n234 163.367
R1622 B.n240 B.n239 163.367
R1623 B.n244 B.n243 163.367
R1624 B.n248 B.n247 163.367
R1625 B.n252 B.n251 163.367
R1626 B.n256 B.n255 163.367
R1627 B.n260 B.n259 163.367
R1628 B.n264 B.n263 163.367
R1629 B.n268 B.n267 163.367
R1630 B.n272 B.n271 163.367
R1631 B.n276 B.n275 163.367
R1632 B.n280 B.n279 163.367
R1633 B.n284 B.n283 163.367
R1634 B.n288 B.n287 163.367
R1635 B.n292 B.n291 163.367
R1636 B.n296 B.n295 163.367
R1637 B.n300 B.n299 163.367
R1638 B.n304 B.n303 163.367
R1639 B.n308 B.n307 163.367
R1640 B.n312 B.n311 163.367
R1641 B.n316 B.n315 163.367
R1642 B.n320 B.n319 163.367
R1643 B.n324 B.n323 163.367
R1644 B.n328 B.n327 163.367
R1645 B.n332 B.n331 163.367
R1646 B.n336 B.n335 163.367
R1647 B.n340 B.n339 163.367
R1648 B.n344 B.n343 163.367
R1649 B.n348 B.n347 163.367
R1650 B.n775 B.n97 163.367
R1651 B.n696 B.n695 71.676
R1652 B.n690 B.n384 71.676
R1653 B.n687 B.n385 71.676
R1654 B.n683 B.n386 71.676
R1655 B.n679 B.n387 71.676
R1656 B.n675 B.n388 71.676
R1657 B.n671 B.n389 71.676
R1658 B.n667 B.n390 71.676
R1659 B.n663 B.n391 71.676
R1660 B.n659 B.n392 71.676
R1661 B.n655 B.n393 71.676
R1662 B.n651 B.n394 71.676
R1663 B.n647 B.n395 71.676
R1664 B.n643 B.n396 71.676
R1665 B.n639 B.n397 71.676
R1666 B.n635 B.n398 71.676
R1667 B.n631 B.n399 71.676
R1668 B.n627 B.n400 71.676
R1669 B.n623 B.n401 71.676
R1670 B.n619 B.n402 71.676
R1671 B.n615 B.n403 71.676
R1672 B.n611 B.n404 71.676
R1673 B.n607 B.n405 71.676
R1674 B.n603 B.n406 71.676
R1675 B.n599 B.n407 71.676
R1676 B.n595 B.n408 71.676
R1677 B.n591 B.n409 71.676
R1678 B.n587 B.n410 71.676
R1679 B.n583 B.n411 71.676
R1680 B.n578 B.n412 71.676
R1681 B.n574 B.n413 71.676
R1682 B.n570 B.n414 71.676
R1683 B.n566 B.n415 71.676
R1684 B.n562 B.n416 71.676
R1685 B.n558 B.n417 71.676
R1686 B.n554 B.n418 71.676
R1687 B.n550 B.n419 71.676
R1688 B.n546 B.n420 71.676
R1689 B.n542 B.n421 71.676
R1690 B.n538 B.n422 71.676
R1691 B.n534 B.n423 71.676
R1692 B.n530 B.n424 71.676
R1693 B.n526 B.n425 71.676
R1694 B.n522 B.n426 71.676
R1695 B.n518 B.n427 71.676
R1696 B.n514 B.n428 71.676
R1697 B.n510 B.n429 71.676
R1698 B.n506 B.n430 71.676
R1699 B.n502 B.n431 71.676
R1700 B.n498 B.n432 71.676
R1701 B.n494 B.n433 71.676
R1702 B.n490 B.n434 71.676
R1703 B.n486 B.n435 71.676
R1704 B.n482 B.n436 71.676
R1705 B.n478 B.n437 71.676
R1706 B.n474 B.n438 71.676
R1707 B.n470 B.n439 71.676
R1708 B.n466 B.n440 71.676
R1709 B.n462 B.n441 71.676
R1710 B.n458 B.n442 71.676
R1711 B.n454 B.n443 71.676
R1712 B.n698 B.n383 71.676
R1713 B.n103 B.n35 71.676
R1714 B.n107 B.n36 71.676
R1715 B.n111 B.n37 71.676
R1716 B.n115 B.n38 71.676
R1717 B.n119 B.n39 71.676
R1718 B.n123 B.n40 71.676
R1719 B.n127 B.n41 71.676
R1720 B.n131 B.n42 71.676
R1721 B.n135 B.n43 71.676
R1722 B.n139 B.n44 71.676
R1723 B.n143 B.n45 71.676
R1724 B.n147 B.n46 71.676
R1725 B.n151 B.n47 71.676
R1726 B.n155 B.n48 71.676
R1727 B.n159 B.n49 71.676
R1728 B.n163 B.n50 71.676
R1729 B.n167 B.n51 71.676
R1730 B.n171 B.n52 71.676
R1731 B.n175 B.n53 71.676
R1732 B.n179 B.n54 71.676
R1733 B.n183 B.n55 71.676
R1734 B.n187 B.n56 71.676
R1735 B.n191 B.n57 71.676
R1736 B.n195 B.n58 71.676
R1737 B.n199 B.n59 71.676
R1738 B.n203 B.n60 71.676
R1739 B.n207 B.n61 71.676
R1740 B.n211 B.n62 71.676
R1741 B.n215 B.n63 71.676
R1742 B.n219 B.n64 71.676
R1743 B.n223 B.n65 71.676
R1744 B.n227 B.n66 71.676
R1745 B.n231 B.n67 71.676
R1746 B.n235 B.n68 71.676
R1747 B.n240 B.n69 71.676
R1748 B.n244 B.n70 71.676
R1749 B.n248 B.n71 71.676
R1750 B.n252 B.n72 71.676
R1751 B.n256 B.n73 71.676
R1752 B.n260 B.n74 71.676
R1753 B.n264 B.n75 71.676
R1754 B.n268 B.n76 71.676
R1755 B.n272 B.n77 71.676
R1756 B.n276 B.n78 71.676
R1757 B.n280 B.n79 71.676
R1758 B.n284 B.n80 71.676
R1759 B.n288 B.n81 71.676
R1760 B.n292 B.n82 71.676
R1761 B.n296 B.n83 71.676
R1762 B.n300 B.n84 71.676
R1763 B.n304 B.n85 71.676
R1764 B.n308 B.n86 71.676
R1765 B.n312 B.n87 71.676
R1766 B.n316 B.n88 71.676
R1767 B.n320 B.n89 71.676
R1768 B.n324 B.n90 71.676
R1769 B.n328 B.n91 71.676
R1770 B.n332 B.n92 71.676
R1771 B.n336 B.n93 71.676
R1772 B.n340 B.n94 71.676
R1773 B.n344 B.n95 71.676
R1774 B.n348 B.n96 71.676
R1775 B.n97 B.n96 71.676
R1776 B.n347 B.n95 71.676
R1777 B.n343 B.n94 71.676
R1778 B.n339 B.n93 71.676
R1779 B.n335 B.n92 71.676
R1780 B.n331 B.n91 71.676
R1781 B.n327 B.n90 71.676
R1782 B.n323 B.n89 71.676
R1783 B.n319 B.n88 71.676
R1784 B.n315 B.n87 71.676
R1785 B.n311 B.n86 71.676
R1786 B.n307 B.n85 71.676
R1787 B.n303 B.n84 71.676
R1788 B.n299 B.n83 71.676
R1789 B.n295 B.n82 71.676
R1790 B.n291 B.n81 71.676
R1791 B.n287 B.n80 71.676
R1792 B.n283 B.n79 71.676
R1793 B.n279 B.n78 71.676
R1794 B.n275 B.n77 71.676
R1795 B.n271 B.n76 71.676
R1796 B.n267 B.n75 71.676
R1797 B.n263 B.n74 71.676
R1798 B.n259 B.n73 71.676
R1799 B.n255 B.n72 71.676
R1800 B.n251 B.n71 71.676
R1801 B.n247 B.n70 71.676
R1802 B.n243 B.n69 71.676
R1803 B.n239 B.n68 71.676
R1804 B.n234 B.n67 71.676
R1805 B.n230 B.n66 71.676
R1806 B.n226 B.n65 71.676
R1807 B.n222 B.n64 71.676
R1808 B.n218 B.n63 71.676
R1809 B.n214 B.n62 71.676
R1810 B.n210 B.n61 71.676
R1811 B.n206 B.n60 71.676
R1812 B.n202 B.n59 71.676
R1813 B.n198 B.n58 71.676
R1814 B.n194 B.n57 71.676
R1815 B.n190 B.n56 71.676
R1816 B.n186 B.n55 71.676
R1817 B.n182 B.n54 71.676
R1818 B.n178 B.n53 71.676
R1819 B.n174 B.n52 71.676
R1820 B.n170 B.n51 71.676
R1821 B.n166 B.n50 71.676
R1822 B.n162 B.n49 71.676
R1823 B.n158 B.n48 71.676
R1824 B.n154 B.n47 71.676
R1825 B.n150 B.n46 71.676
R1826 B.n146 B.n45 71.676
R1827 B.n142 B.n44 71.676
R1828 B.n138 B.n43 71.676
R1829 B.n134 B.n42 71.676
R1830 B.n130 B.n41 71.676
R1831 B.n126 B.n40 71.676
R1832 B.n122 B.n39 71.676
R1833 B.n118 B.n38 71.676
R1834 B.n114 B.n37 71.676
R1835 B.n110 B.n36 71.676
R1836 B.n106 B.n35 71.676
R1837 B.n696 B.n445 71.676
R1838 B.n688 B.n384 71.676
R1839 B.n684 B.n385 71.676
R1840 B.n680 B.n386 71.676
R1841 B.n676 B.n387 71.676
R1842 B.n672 B.n388 71.676
R1843 B.n668 B.n389 71.676
R1844 B.n664 B.n390 71.676
R1845 B.n660 B.n391 71.676
R1846 B.n656 B.n392 71.676
R1847 B.n652 B.n393 71.676
R1848 B.n648 B.n394 71.676
R1849 B.n644 B.n395 71.676
R1850 B.n640 B.n396 71.676
R1851 B.n636 B.n397 71.676
R1852 B.n632 B.n398 71.676
R1853 B.n628 B.n399 71.676
R1854 B.n624 B.n400 71.676
R1855 B.n620 B.n401 71.676
R1856 B.n616 B.n402 71.676
R1857 B.n612 B.n403 71.676
R1858 B.n608 B.n404 71.676
R1859 B.n604 B.n405 71.676
R1860 B.n600 B.n406 71.676
R1861 B.n596 B.n407 71.676
R1862 B.n592 B.n408 71.676
R1863 B.n588 B.n409 71.676
R1864 B.n584 B.n410 71.676
R1865 B.n579 B.n411 71.676
R1866 B.n575 B.n412 71.676
R1867 B.n571 B.n413 71.676
R1868 B.n567 B.n414 71.676
R1869 B.n563 B.n415 71.676
R1870 B.n559 B.n416 71.676
R1871 B.n555 B.n417 71.676
R1872 B.n551 B.n418 71.676
R1873 B.n547 B.n419 71.676
R1874 B.n543 B.n420 71.676
R1875 B.n539 B.n421 71.676
R1876 B.n535 B.n422 71.676
R1877 B.n531 B.n423 71.676
R1878 B.n527 B.n424 71.676
R1879 B.n523 B.n425 71.676
R1880 B.n519 B.n426 71.676
R1881 B.n515 B.n427 71.676
R1882 B.n511 B.n428 71.676
R1883 B.n507 B.n429 71.676
R1884 B.n503 B.n430 71.676
R1885 B.n499 B.n431 71.676
R1886 B.n495 B.n432 71.676
R1887 B.n491 B.n433 71.676
R1888 B.n487 B.n434 71.676
R1889 B.n483 B.n435 71.676
R1890 B.n479 B.n436 71.676
R1891 B.n475 B.n437 71.676
R1892 B.n471 B.n438 71.676
R1893 B.n467 B.n439 71.676
R1894 B.n463 B.n440 71.676
R1895 B.n459 B.n441 71.676
R1896 B.n455 B.n442 71.676
R1897 B.n451 B.n443 71.676
R1898 B.n699 B.n698 71.676
R1899 B.n450 B.n449 59.5399
R1900 B.n581 B.n447 59.5399
R1901 B.n102 B.n101 59.5399
R1902 B.n237 B.n99 59.5399
R1903 B.n697 B.n380 57.6784
R1904 B.n777 B.n776 57.6784
R1905 B.n704 B.n380 32.9593
R1906 B.n704 B.n375 32.9593
R1907 B.n710 B.n375 32.9593
R1908 B.n710 B.n376 32.9593
R1909 B.n716 B.n368 32.9593
R1910 B.n722 B.n368 32.9593
R1911 B.n722 B.n364 32.9593
R1912 B.n728 B.n364 32.9593
R1913 B.n734 B.n359 32.9593
R1914 B.n734 B.n360 32.9593
R1915 B.n742 B.n741 32.9593
R1916 B.n748 B.n4 32.9593
R1917 B.n810 B.n4 32.9593
R1918 B.n810 B.n809 32.9593
R1919 B.n809 B.n808 32.9593
R1920 B.n802 B.n11 32.9593
R1921 B.n801 B.n800 32.9593
R1922 B.n800 B.n15 32.9593
R1923 B.n794 B.n793 32.9593
R1924 B.n793 B.n792 32.9593
R1925 B.n792 B.n22 32.9593
R1926 B.n786 B.n22 32.9593
R1927 B.n785 B.n784 32.9593
R1928 B.n784 B.n29 32.9593
R1929 B.n778 B.n29 32.9593
R1930 B.n778 B.n777 32.9593
R1931 B.n104 B.n31 30.1273
R1932 B.n774 B.n773 30.1273
R1933 B.n701 B.n700 30.1273
R1934 B.n694 B.n378 30.1273
R1935 B.n742 B.t4 30.0512
R1936 B.n802 B.t2 30.0512
R1937 B.n728 B.t0 29.0818
R1938 B.n794 B.t5 29.0818
R1939 B.n748 B.t1 23.2655
R1940 B.n808 B.t3 23.2655
R1941 B B.n812 18.0485
R1942 B.n716 B.t7 17.4493
R1943 B.n786 B.t11 17.4493
R1944 B.n376 B.t7 15.5105
R1945 B.t11 B.n785 15.5105
R1946 B.n449 B.n448 14.546
R1947 B.n447 B.n446 14.546
R1948 B.n101 B.n100 14.546
R1949 B.n99 B.n98 14.546
R1950 B.n105 B.n104 10.6151
R1951 B.n108 B.n105 10.6151
R1952 B.n109 B.n108 10.6151
R1953 B.n112 B.n109 10.6151
R1954 B.n113 B.n112 10.6151
R1955 B.n116 B.n113 10.6151
R1956 B.n117 B.n116 10.6151
R1957 B.n120 B.n117 10.6151
R1958 B.n121 B.n120 10.6151
R1959 B.n124 B.n121 10.6151
R1960 B.n125 B.n124 10.6151
R1961 B.n128 B.n125 10.6151
R1962 B.n129 B.n128 10.6151
R1963 B.n132 B.n129 10.6151
R1964 B.n133 B.n132 10.6151
R1965 B.n136 B.n133 10.6151
R1966 B.n137 B.n136 10.6151
R1967 B.n140 B.n137 10.6151
R1968 B.n141 B.n140 10.6151
R1969 B.n144 B.n141 10.6151
R1970 B.n145 B.n144 10.6151
R1971 B.n148 B.n145 10.6151
R1972 B.n149 B.n148 10.6151
R1973 B.n152 B.n149 10.6151
R1974 B.n153 B.n152 10.6151
R1975 B.n156 B.n153 10.6151
R1976 B.n157 B.n156 10.6151
R1977 B.n160 B.n157 10.6151
R1978 B.n161 B.n160 10.6151
R1979 B.n164 B.n161 10.6151
R1980 B.n165 B.n164 10.6151
R1981 B.n168 B.n165 10.6151
R1982 B.n169 B.n168 10.6151
R1983 B.n172 B.n169 10.6151
R1984 B.n173 B.n172 10.6151
R1985 B.n176 B.n173 10.6151
R1986 B.n177 B.n176 10.6151
R1987 B.n180 B.n177 10.6151
R1988 B.n181 B.n180 10.6151
R1989 B.n184 B.n181 10.6151
R1990 B.n185 B.n184 10.6151
R1991 B.n188 B.n185 10.6151
R1992 B.n189 B.n188 10.6151
R1993 B.n192 B.n189 10.6151
R1994 B.n193 B.n192 10.6151
R1995 B.n196 B.n193 10.6151
R1996 B.n197 B.n196 10.6151
R1997 B.n200 B.n197 10.6151
R1998 B.n201 B.n200 10.6151
R1999 B.n204 B.n201 10.6151
R2000 B.n205 B.n204 10.6151
R2001 B.n208 B.n205 10.6151
R2002 B.n209 B.n208 10.6151
R2003 B.n212 B.n209 10.6151
R2004 B.n213 B.n212 10.6151
R2005 B.n216 B.n213 10.6151
R2006 B.n217 B.n216 10.6151
R2007 B.n221 B.n220 10.6151
R2008 B.n224 B.n221 10.6151
R2009 B.n225 B.n224 10.6151
R2010 B.n228 B.n225 10.6151
R2011 B.n229 B.n228 10.6151
R2012 B.n232 B.n229 10.6151
R2013 B.n233 B.n232 10.6151
R2014 B.n236 B.n233 10.6151
R2015 B.n241 B.n238 10.6151
R2016 B.n242 B.n241 10.6151
R2017 B.n245 B.n242 10.6151
R2018 B.n246 B.n245 10.6151
R2019 B.n249 B.n246 10.6151
R2020 B.n250 B.n249 10.6151
R2021 B.n253 B.n250 10.6151
R2022 B.n254 B.n253 10.6151
R2023 B.n257 B.n254 10.6151
R2024 B.n258 B.n257 10.6151
R2025 B.n261 B.n258 10.6151
R2026 B.n262 B.n261 10.6151
R2027 B.n265 B.n262 10.6151
R2028 B.n266 B.n265 10.6151
R2029 B.n269 B.n266 10.6151
R2030 B.n270 B.n269 10.6151
R2031 B.n273 B.n270 10.6151
R2032 B.n274 B.n273 10.6151
R2033 B.n277 B.n274 10.6151
R2034 B.n278 B.n277 10.6151
R2035 B.n281 B.n278 10.6151
R2036 B.n282 B.n281 10.6151
R2037 B.n285 B.n282 10.6151
R2038 B.n286 B.n285 10.6151
R2039 B.n289 B.n286 10.6151
R2040 B.n290 B.n289 10.6151
R2041 B.n293 B.n290 10.6151
R2042 B.n294 B.n293 10.6151
R2043 B.n297 B.n294 10.6151
R2044 B.n298 B.n297 10.6151
R2045 B.n301 B.n298 10.6151
R2046 B.n302 B.n301 10.6151
R2047 B.n305 B.n302 10.6151
R2048 B.n306 B.n305 10.6151
R2049 B.n309 B.n306 10.6151
R2050 B.n310 B.n309 10.6151
R2051 B.n313 B.n310 10.6151
R2052 B.n314 B.n313 10.6151
R2053 B.n317 B.n314 10.6151
R2054 B.n318 B.n317 10.6151
R2055 B.n321 B.n318 10.6151
R2056 B.n322 B.n321 10.6151
R2057 B.n325 B.n322 10.6151
R2058 B.n326 B.n325 10.6151
R2059 B.n329 B.n326 10.6151
R2060 B.n330 B.n329 10.6151
R2061 B.n333 B.n330 10.6151
R2062 B.n334 B.n333 10.6151
R2063 B.n337 B.n334 10.6151
R2064 B.n338 B.n337 10.6151
R2065 B.n341 B.n338 10.6151
R2066 B.n342 B.n341 10.6151
R2067 B.n345 B.n342 10.6151
R2068 B.n346 B.n345 10.6151
R2069 B.n349 B.n346 10.6151
R2070 B.n350 B.n349 10.6151
R2071 B.n774 B.n350 10.6151
R2072 B.n702 B.n701 10.6151
R2073 B.n702 B.n373 10.6151
R2074 B.n712 B.n373 10.6151
R2075 B.n713 B.n712 10.6151
R2076 B.n714 B.n713 10.6151
R2077 B.n714 B.n366 10.6151
R2078 B.n724 B.n366 10.6151
R2079 B.n725 B.n724 10.6151
R2080 B.n726 B.n725 10.6151
R2081 B.n726 B.n357 10.6151
R2082 B.n736 B.n357 10.6151
R2083 B.n737 B.n736 10.6151
R2084 B.n739 B.n737 10.6151
R2085 B.n739 B.n738 10.6151
R2086 B.n738 B.n351 10.6151
R2087 B.n751 B.n351 10.6151
R2088 B.n752 B.n751 10.6151
R2089 B.n753 B.n752 10.6151
R2090 B.n754 B.n753 10.6151
R2091 B.n756 B.n754 10.6151
R2092 B.n757 B.n756 10.6151
R2093 B.n758 B.n757 10.6151
R2094 B.n759 B.n758 10.6151
R2095 B.n761 B.n759 10.6151
R2096 B.n762 B.n761 10.6151
R2097 B.n763 B.n762 10.6151
R2098 B.n764 B.n763 10.6151
R2099 B.n766 B.n764 10.6151
R2100 B.n767 B.n766 10.6151
R2101 B.n768 B.n767 10.6151
R2102 B.n769 B.n768 10.6151
R2103 B.n771 B.n769 10.6151
R2104 B.n772 B.n771 10.6151
R2105 B.n773 B.n772 10.6151
R2106 B.n694 B.n693 10.6151
R2107 B.n693 B.n692 10.6151
R2108 B.n692 B.n691 10.6151
R2109 B.n691 B.n689 10.6151
R2110 B.n689 B.n686 10.6151
R2111 B.n686 B.n685 10.6151
R2112 B.n685 B.n682 10.6151
R2113 B.n682 B.n681 10.6151
R2114 B.n681 B.n678 10.6151
R2115 B.n678 B.n677 10.6151
R2116 B.n677 B.n674 10.6151
R2117 B.n674 B.n673 10.6151
R2118 B.n673 B.n670 10.6151
R2119 B.n670 B.n669 10.6151
R2120 B.n669 B.n666 10.6151
R2121 B.n666 B.n665 10.6151
R2122 B.n665 B.n662 10.6151
R2123 B.n662 B.n661 10.6151
R2124 B.n661 B.n658 10.6151
R2125 B.n658 B.n657 10.6151
R2126 B.n657 B.n654 10.6151
R2127 B.n654 B.n653 10.6151
R2128 B.n653 B.n650 10.6151
R2129 B.n650 B.n649 10.6151
R2130 B.n649 B.n646 10.6151
R2131 B.n646 B.n645 10.6151
R2132 B.n645 B.n642 10.6151
R2133 B.n642 B.n641 10.6151
R2134 B.n641 B.n638 10.6151
R2135 B.n638 B.n637 10.6151
R2136 B.n637 B.n634 10.6151
R2137 B.n634 B.n633 10.6151
R2138 B.n633 B.n630 10.6151
R2139 B.n630 B.n629 10.6151
R2140 B.n629 B.n626 10.6151
R2141 B.n626 B.n625 10.6151
R2142 B.n625 B.n622 10.6151
R2143 B.n622 B.n621 10.6151
R2144 B.n621 B.n618 10.6151
R2145 B.n618 B.n617 10.6151
R2146 B.n617 B.n614 10.6151
R2147 B.n614 B.n613 10.6151
R2148 B.n613 B.n610 10.6151
R2149 B.n610 B.n609 10.6151
R2150 B.n609 B.n606 10.6151
R2151 B.n606 B.n605 10.6151
R2152 B.n605 B.n602 10.6151
R2153 B.n602 B.n601 10.6151
R2154 B.n601 B.n598 10.6151
R2155 B.n598 B.n597 10.6151
R2156 B.n597 B.n594 10.6151
R2157 B.n594 B.n593 10.6151
R2158 B.n593 B.n590 10.6151
R2159 B.n590 B.n589 10.6151
R2160 B.n589 B.n586 10.6151
R2161 B.n586 B.n585 10.6151
R2162 B.n585 B.n582 10.6151
R2163 B.n580 B.n577 10.6151
R2164 B.n577 B.n576 10.6151
R2165 B.n576 B.n573 10.6151
R2166 B.n573 B.n572 10.6151
R2167 B.n572 B.n569 10.6151
R2168 B.n569 B.n568 10.6151
R2169 B.n568 B.n565 10.6151
R2170 B.n565 B.n564 10.6151
R2171 B.n561 B.n560 10.6151
R2172 B.n560 B.n557 10.6151
R2173 B.n557 B.n556 10.6151
R2174 B.n556 B.n553 10.6151
R2175 B.n553 B.n552 10.6151
R2176 B.n552 B.n549 10.6151
R2177 B.n549 B.n548 10.6151
R2178 B.n548 B.n545 10.6151
R2179 B.n545 B.n544 10.6151
R2180 B.n544 B.n541 10.6151
R2181 B.n541 B.n540 10.6151
R2182 B.n540 B.n537 10.6151
R2183 B.n537 B.n536 10.6151
R2184 B.n536 B.n533 10.6151
R2185 B.n533 B.n532 10.6151
R2186 B.n532 B.n529 10.6151
R2187 B.n529 B.n528 10.6151
R2188 B.n528 B.n525 10.6151
R2189 B.n525 B.n524 10.6151
R2190 B.n524 B.n521 10.6151
R2191 B.n521 B.n520 10.6151
R2192 B.n520 B.n517 10.6151
R2193 B.n517 B.n516 10.6151
R2194 B.n516 B.n513 10.6151
R2195 B.n513 B.n512 10.6151
R2196 B.n512 B.n509 10.6151
R2197 B.n509 B.n508 10.6151
R2198 B.n508 B.n505 10.6151
R2199 B.n505 B.n504 10.6151
R2200 B.n504 B.n501 10.6151
R2201 B.n501 B.n500 10.6151
R2202 B.n500 B.n497 10.6151
R2203 B.n497 B.n496 10.6151
R2204 B.n496 B.n493 10.6151
R2205 B.n493 B.n492 10.6151
R2206 B.n492 B.n489 10.6151
R2207 B.n489 B.n488 10.6151
R2208 B.n488 B.n485 10.6151
R2209 B.n485 B.n484 10.6151
R2210 B.n484 B.n481 10.6151
R2211 B.n481 B.n480 10.6151
R2212 B.n480 B.n477 10.6151
R2213 B.n477 B.n476 10.6151
R2214 B.n476 B.n473 10.6151
R2215 B.n473 B.n472 10.6151
R2216 B.n472 B.n469 10.6151
R2217 B.n469 B.n468 10.6151
R2218 B.n468 B.n465 10.6151
R2219 B.n465 B.n464 10.6151
R2220 B.n464 B.n461 10.6151
R2221 B.n461 B.n460 10.6151
R2222 B.n460 B.n457 10.6151
R2223 B.n457 B.n456 10.6151
R2224 B.n456 B.n453 10.6151
R2225 B.n453 B.n452 10.6151
R2226 B.n452 B.n382 10.6151
R2227 B.n700 B.n382 10.6151
R2228 B.n706 B.n378 10.6151
R2229 B.n707 B.n706 10.6151
R2230 B.n708 B.n707 10.6151
R2231 B.n708 B.n370 10.6151
R2232 B.n718 B.n370 10.6151
R2233 B.n719 B.n718 10.6151
R2234 B.n720 B.n719 10.6151
R2235 B.n720 B.n362 10.6151
R2236 B.n730 B.n362 10.6151
R2237 B.n731 B.n730 10.6151
R2238 B.n732 B.n731 10.6151
R2239 B.n732 B.n354 10.6151
R2240 B.n744 B.n354 10.6151
R2241 B.n745 B.n744 10.6151
R2242 B.n746 B.n745 10.6151
R2243 B.n746 B.n0 10.6151
R2244 B.n806 B.n1 10.6151
R2245 B.n806 B.n805 10.6151
R2246 B.n805 B.n804 10.6151
R2247 B.n804 B.n9 10.6151
R2248 B.n798 B.n9 10.6151
R2249 B.n798 B.n797 10.6151
R2250 B.n797 B.n796 10.6151
R2251 B.n796 B.n17 10.6151
R2252 B.n790 B.n17 10.6151
R2253 B.n790 B.n789 10.6151
R2254 B.n789 B.n788 10.6151
R2255 B.n788 B.n24 10.6151
R2256 B.n782 B.n24 10.6151
R2257 B.n782 B.n781 10.6151
R2258 B.n781 B.n780 10.6151
R2259 B.n780 B.n31 10.6151
R2260 B.n741 B.t1 9.69427
R2261 B.n11 B.t3 9.69427
R2262 B.n220 B.n102 6.5566
R2263 B.n237 B.n236 6.5566
R2264 B.n581 B.n580 6.5566
R2265 B.n564 B.n450 6.5566
R2266 B.n217 B.n102 4.05904
R2267 B.n238 B.n237 4.05904
R2268 B.n582 B.n581 4.05904
R2269 B.n561 B.n450 4.05904
R2270 B.t0 B.n359 3.87801
R2271 B.t5 B.n15 3.87801
R2272 B.n360 B.t4 2.90863
R2273 B.t2 B.n801 2.90863
R2274 B.n812 B.n0 2.81026
R2275 B.n812 B.n1 2.81026
R2276 VP.n1 VP.t0 1118.83
R2277 VP.n8 VP.t4 1100.1
R2278 VP.n6 VP.t2 1100.1
R2279 VP.n3 VP.t3 1100.1
R2280 VP.n7 VP.t1 1094.25
R2281 VP.n2 VP.t5 1094.25
R2282 VP.n9 VP.n8 161.3
R2283 VP.n4 VP.n3 161.3
R2284 VP.n7 VP.n0 161.3
R2285 VP.n6 VP.n5 161.3
R2286 VP.n4 VP.n1 71.5267
R2287 VP.n5 VP.n4 44.3073
R2288 VP.n7 VP.n6 42.3581
R2289 VP.n8 VP.n7 42.3581
R2290 VP.n3 VP.n2 42.3581
R2291 VP.n2 VP.n1 18.712
R2292 VP.n5 VP.n0 0.189894
R2293 VP.n9 VP.n0 0.189894
R2294 VP VP.n9 0.0516364
R2295 VDD1.n92 VDD1.n0 289.615
R2296 VDD1.n189 VDD1.n97 289.615
R2297 VDD1.n93 VDD1.n92 185
R2298 VDD1.n91 VDD1.n90 185
R2299 VDD1.n4 VDD1.n3 185
R2300 VDD1.n85 VDD1.n84 185
R2301 VDD1.n83 VDD1.n82 185
R2302 VDD1.n8 VDD1.n7 185
R2303 VDD1.n12 VDD1.n10 185
R2304 VDD1.n77 VDD1.n76 185
R2305 VDD1.n75 VDD1.n74 185
R2306 VDD1.n14 VDD1.n13 185
R2307 VDD1.n69 VDD1.n68 185
R2308 VDD1.n67 VDD1.n66 185
R2309 VDD1.n18 VDD1.n17 185
R2310 VDD1.n61 VDD1.n60 185
R2311 VDD1.n59 VDD1.n58 185
R2312 VDD1.n22 VDD1.n21 185
R2313 VDD1.n53 VDD1.n52 185
R2314 VDD1.n51 VDD1.n50 185
R2315 VDD1.n26 VDD1.n25 185
R2316 VDD1.n45 VDD1.n44 185
R2317 VDD1.n43 VDD1.n42 185
R2318 VDD1.n30 VDD1.n29 185
R2319 VDD1.n37 VDD1.n36 185
R2320 VDD1.n35 VDD1.n34 185
R2321 VDD1.n130 VDD1.n129 185
R2322 VDD1.n132 VDD1.n131 185
R2323 VDD1.n125 VDD1.n124 185
R2324 VDD1.n138 VDD1.n137 185
R2325 VDD1.n140 VDD1.n139 185
R2326 VDD1.n121 VDD1.n120 185
R2327 VDD1.n146 VDD1.n145 185
R2328 VDD1.n148 VDD1.n147 185
R2329 VDD1.n117 VDD1.n116 185
R2330 VDD1.n154 VDD1.n153 185
R2331 VDD1.n156 VDD1.n155 185
R2332 VDD1.n113 VDD1.n112 185
R2333 VDD1.n162 VDD1.n161 185
R2334 VDD1.n164 VDD1.n163 185
R2335 VDD1.n109 VDD1.n108 185
R2336 VDD1.n171 VDD1.n170 185
R2337 VDD1.n172 VDD1.n107 185
R2338 VDD1.n174 VDD1.n173 185
R2339 VDD1.n105 VDD1.n104 185
R2340 VDD1.n180 VDD1.n179 185
R2341 VDD1.n182 VDD1.n181 185
R2342 VDD1.n101 VDD1.n100 185
R2343 VDD1.n188 VDD1.n187 185
R2344 VDD1.n190 VDD1.n189 185
R2345 VDD1.n33 VDD1.t5 147.659
R2346 VDD1.n128 VDD1.t3 147.659
R2347 VDD1.n92 VDD1.n91 104.615
R2348 VDD1.n91 VDD1.n3 104.615
R2349 VDD1.n84 VDD1.n3 104.615
R2350 VDD1.n84 VDD1.n83 104.615
R2351 VDD1.n83 VDD1.n7 104.615
R2352 VDD1.n12 VDD1.n7 104.615
R2353 VDD1.n76 VDD1.n12 104.615
R2354 VDD1.n76 VDD1.n75 104.615
R2355 VDD1.n75 VDD1.n13 104.615
R2356 VDD1.n68 VDD1.n13 104.615
R2357 VDD1.n68 VDD1.n67 104.615
R2358 VDD1.n67 VDD1.n17 104.615
R2359 VDD1.n60 VDD1.n17 104.615
R2360 VDD1.n60 VDD1.n59 104.615
R2361 VDD1.n59 VDD1.n21 104.615
R2362 VDD1.n52 VDD1.n21 104.615
R2363 VDD1.n52 VDD1.n51 104.615
R2364 VDD1.n51 VDD1.n25 104.615
R2365 VDD1.n44 VDD1.n25 104.615
R2366 VDD1.n44 VDD1.n43 104.615
R2367 VDD1.n43 VDD1.n29 104.615
R2368 VDD1.n36 VDD1.n29 104.615
R2369 VDD1.n36 VDD1.n35 104.615
R2370 VDD1.n131 VDD1.n130 104.615
R2371 VDD1.n131 VDD1.n124 104.615
R2372 VDD1.n138 VDD1.n124 104.615
R2373 VDD1.n139 VDD1.n138 104.615
R2374 VDD1.n139 VDD1.n120 104.615
R2375 VDD1.n146 VDD1.n120 104.615
R2376 VDD1.n147 VDD1.n146 104.615
R2377 VDD1.n147 VDD1.n116 104.615
R2378 VDD1.n154 VDD1.n116 104.615
R2379 VDD1.n155 VDD1.n154 104.615
R2380 VDD1.n155 VDD1.n112 104.615
R2381 VDD1.n162 VDD1.n112 104.615
R2382 VDD1.n163 VDD1.n162 104.615
R2383 VDD1.n163 VDD1.n108 104.615
R2384 VDD1.n171 VDD1.n108 104.615
R2385 VDD1.n172 VDD1.n171 104.615
R2386 VDD1.n173 VDD1.n172 104.615
R2387 VDD1.n173 VDD1.n104 104.615
R2388 VDD1.n180 VDD1.n104 104.615
R2389 VDD1.n181 VDD1.n180 104.615
R2390 VDD1.n181 VDD1.n100 104.615
R2391 VDD1.n188 VDD1.n100 104.615
R2392 VDD1.n189 VDD1.n188 104.615
R2393 VDD1.n195 VDD1.n194 58.8489
R2394 VDD1.n197 VDD1.n196 58.7426
R2395 VDD1.n35 VDD1.t5 52.3082
R2396 VDD1.n130 VDD1.t3 52.3082
R2397 VDD1 VDD1.n96 47.4678
R2398 VDD1.n195 VDD1.n193 47.3543
R2399 VDD1.n197 VDD1.n195 41.7401
R2400 VDD1.n34 VDD1.n33 15.6677
R2401 VDD1.n129 VDD1.n128 15.6677
R2402 VDD1.n10 VDD1.n8 13.1884
R2403 VDD1.n174 VDD1.n105 13.1884
R2404 VDD1.n82 VDD1.n81 12.8005
R2405 VDD1.n78 VDD1.n77 12.8005
R2406 VDD1.n37 VDD1.n32 12.8005
R2407 VDD1.n132 VDD1.n127 12.8005
R2408 VDD1.n175 VDD1.n107 12.8005
R2409 VDD1.n179 VDD1.n178 12.8005
R2410 VDD1.n85 VDD1.n6 12.0247
R2411 VDD1.n74 VDD1.n11 12.0247
R2412 VDD1.n38 VDD1.n30 12.0247
R2413 VDD1.n133 VDD1.n125 12.0247
R2414 VDD1.n170 VDD1.n169 12.0247
R2415 VDD1.n182 VDD1.n103 12.0247
R2416 VDD1.n86 VDD1.n4 11.249
R2417 VDD1.n73 VDD1.n14 11.249
R2418 VDD1.n42 VDD1.n41 11.249
R2419 VDD1.n137 VDD1.n136 11.249
R2420 VDD1.n168 VDD1.n109 11.249
R2421 VDD1.n183 VDD1.n101 11.249
R2422 VDD1.n90 VDD1.n89 10.4732
R2423 VDD1.n70 VDD1.n69 10.4732
R2424 VDD1.n45 VDD1.n28 10.4732
R2425 VDD1.n140 VDD1.n123 10.4732
R2426 VDD1.n165 VDD1.n164 10.4732
R2427 VDD1.n187 VDD1.n186 10.4732
R2428 VDD1.n93 VDD1.n2 9.69747
R2429 VDD1.n66 VDD1.n16 9.69747
R2430 VDD1.n46 VDD1.n26 9.69747
R2431 VDD1.n141 VDD1.n121 9.69747
R2432 VDD1.n161 VDD1.n111 9.69747
R2433 VDD1.n190 VDD1.n99 9.69747
R2434 VDD1.n96 VDD1.n95 9.45567
R2435 VDD1.n193 VDD1.n192 9.45567
R2436 VDD1.n20 VDD1.n19 9.3005
R2437 VDD1.n63 VDD1.n62 9.3005
R2438 VDD1.n65 VDD1.n64 9.3005
R2439 VDD1.n16 VDD1.n15 9.3005
R2440 VDD1.n71 VDD1.n70 9.3005
R2441 VDD1.n73 VDD1.n72 9.3005
R2442 VDD1.n11 VDD1.n9 9.3005
R2443 VDD1.n79 VDD1.n78 9.3005
R2444 VDD1.n95 VDD1.n94 9.3005
R2445 VDD1.n2 VDD1.n1 9.3005
R2446 VDD1.n89 VDD1.n88 9.3005
R2447 VDD1.n87 VDD1.n86 9.3005
R2448 VDD1.n6 VDD1.n5 9.3005
R2449 VDD1.n81 VDD1.n80 9.3005
R2450 VDD1.n57 VDD1.n56 9.3005
R2451 VDD1.n55 VDD1.n54 9.3005
R2452 VDD1.n24 VDD1.n23 9.3005
R2453 VDD1.n49 VDD1.n48 9.3005
R2454 VDD1.n47 VDD1.n46 9.3005
R2455 VDD1.n28 VDD1.n27 9.3005
R2456 VDD1.n41 VDD1.n40 9.3005
R2457 VDD1.n39 VDD1.n38 9.3005
R2458 VDD1.n32 VDD1.n31 9.3005
R2459 VDD1.n192 VDD1.n191 9.3005
R2460 VDD1.n99 VDD1.n98 9.3005
R2461 VDD1.n186 VDD1.n185 9.3005
R2462 VDD1.n184 VDD1.n183 9.3005
R2463 VDD1.n103 VDD1.n102 9.3005
R2464 VDD1.n178 VDD1.n177 9.3005
R2465 VDD1.n150 VDD1.n149 9.3005
R2466 VDD1.n119 VDD1.n118 9.3005
R2467 VDD1.n144 VDD1.n143 9.3005
R2468 VDD1.n142 VDD1.n141 9.3005
R2469 VDD1.n123 VDD1.n122 9.3005
R2470 VDD1.n136 VDD1.n135 9.3005
R2471 VDD1.n134 VDD1.n133 9.3005
R2472 VDD1.n127 VDD1.n126 9.3005
R2473 VDD1.n152 VDD1.n151 9.3005
R2474 VDD1.n115 VDD1.n114 9.3005
R2475 VDD1.n158 VDD1.n157 9.3005
R2476 VDD1.n160 VDD1.n159 9.3005
R2477 VDD1.n111 VDD1.n110 9.3005
R2478 VDD1.n166 VDD1.n165 9.3005
R2479 VDD1.n168 VDD1.n167 9.3005
R2480 VDD1.n169 VDD1.n106 9.3005
R2481 VDD1.n176 VDD1.n175 9.3005
R2482 VDD1.n94 VDD1.n0 8.92171
R2483 VDD1.n65 VDD1.n18 8.92171
R2484 VDD1.n50 VDD1.n49 8.92171
R2485 VDD1.n145 VDD1.n144 8.92171
R2486 VDD1.n160 VDD1.n113 8.92171
R2487 VDD1.n191 VDD1.n97 8.92171
R2488 VDD1.n62 VDD1.n61 8.14595
R2489 VDD1.n53 VDD1.n24 8.14595
R2490 VDD1.n148 VDD1.n119 8.14595
R2491 VDD1.n157 VDD1.n156 8.14595
R2492 VDD1.n58 VDD1.n20 7.3702
R2493 VDD1.n54 VDD1.n22 7.3702
R2494 VDD1.n149 VDD1.n117 7.3702
R2495 VDD1.n153 VDD1.n115 7.3702
R2496 VDD1.n58 VDD1.n57 6.59444
R2497 VDD1.n57 VDD1.n22 6.59444
R2498 VDD1.n152 VDD1.n117 6.59444
R2499 VDD1.n153 VDD1.n152 6.59444
R2500 VDD1.n61 VDD1.n20 5.81868
R2501 VDD1.n54 VDD1.n53 5.81868
R2502 VDD1.n149 VDD1.n148 5.81868
R2503 VDD1.n156 VDD1.n115 5.81868
R2504 VDD1.n96 VDD1.n0 5.04292
R2505 VDD1.n62 VDD1.n18 5.04292
R2506 VDD1.n50 VDD1.n24 5.04292
R2507 VDD1.n145 VDD1.n119 5.04292
R2508 VDD1.n157 VDD1.n113 5.04292
R2509 VDD1.n193 VDD1.n97 5.04292
R2510 VDD1.n33 VDD1.n31 4.38563
R2511 VDD1.n128 VDD1.n126 4.38563
R2512 VDD1.n94 VDD1.n93 4.26717
R2513 VDD1.n66 VDD1.n65 4.26717
R2514 VDD1.n49 VDD1.n26 4.26717
R2515 VDD1.n144 VDD1.n121 4.26717
R2516 VDD1.n161 VDD1.n160 4.26717
R2517 VDD1.n191 VDD1.n190 4.26717
R2518 VDD1.n90 VDD1.n2 3.49141
R2519 VDD1.n69 VDD1.n16 3.49141
R2520 VDD1.n46 VDD1.n45 3.49141
R2521 VDD1.n141 VDD1.n140 3.49141
R2522 VDD1.n164 VDD1.n111 3.49141
R2523 VDD1.n187 VDD1.n99 3.49141
R2524 VDD1.n89 VDD1.n4 2.71565
R2525 VDD1.n70 VDD1.n14 2.71565
R2526 VDD1.n42 VDD1.n28 2.71565
R2527 VDD1.n137 VDD1.n123 2.71565
R2528 VDD1.n165 VDD1.n109 2.71565
R2529 VDD1.n186 VDD1.n101 2.71565
R2530 VDD1.n86 VDD1.n85 1.93989
R2531 VDD1.n74 VDD1.n73 1.93989
R2532 VDD1.n41 VDD1.n30 1.93989
R2533 VDD1.n136 VDD1.n125 1.93989
R2534 VDD1.n170 VDD1.n168 1.93989
R2535 VDD1.n183 VDD1.n182 1.93989
R2536 VDD1.n82 VDD1.n6 1.16414
R2537 VDD1.n77 VDD1.n11 1.16414
R2538 VDD1.n38 VDD1.n37 1.16414
R2539 VDD1.n133 VDD1.n132 1.16414
R2540 VDD1.n169 VDD1.n107 1.16414
R2541 VDD1.n179 VDD1.n103 1.16414
R2542 VDD1.n196 VDD1.t0 1.13712
R2543 VDD1.n196 VDD1.t2 1.13712
R2544 VDD1.n194 VDD1.t4 1.13712
R2545 VDD1.n194 VDD1.t1 1.13712
R2546 VDD1.n81 VDD1.n8 0.388379
R2547 VDD1.n78 VDD1.n10 0.388379
R2548 VDD1.n34 VDD1.n32 0.388379
R2549 VDD1.n129 VDD1.n127 0.388379
R2550 VDD1.n175 VDD1.n174 0.388379
R2551 VDD1.n178 VDD1.n105 0.388379
R2552 VDD1.n95 VDD1.n1 0.155672
R2553 VDD1.n88 VDD1.n1 0.155672
R2554 VDD1.n88 VDD1.n87 0.155672
R2555 VDD1.n87 VDD1.n5 0.155672
R2556 VDD1.n80 VDD1.n5 0.155672
R2557 VDD1.n80 VDD1.n79 0.155672
R2558 VDD1.n79 VDD1.n9 0.155672
R2559 VDD1.n72 VDD1.n9 0.155672
R2560 VDD1.n72 VDD1.n71 0.155672
R2561 VDD1.n71 VDD1.n15 0.155672
R2562 VDD1.n64 VDD1.n15 0.155672
R2563 VDD1.n64 VDD1.n63 0.155672
R2564 VDD1.n63 VDD1.n19 0.155672
R2565 VDD1.n56 VDD1.n19 0.155672
R2566 VDD1.n56 VDD1.n55 0.155672
R2567 VDD1.n55 VDD1.n23 0.155672
R2568 VDD1.n48 VDD1.n23 0.155672
R2569 VDD1.n48 VDD1.n47 0.155672
R2570 VDD1.n47 VDD1.n27 0.155672
R2571 VDD1.n40 VDD1.n27 0.155672
R2572 VDD1.n40 VDD1.n39 0.155672
R2573 VDD1.n39 VDD1.n31 0.155672
R2574 VDD1.n134 VDD1.n126 0.155672
R2575 VDD1.n135 VDD1.n134 0.155672
R2576 VDD1.n135 VDD1.n122 0.155672
R2577 VDD1.n142 VDD1.n122 0.155672
R2578 VDD1.n143 VDD1.n142 0.155672
R2579 VDD1.n143 VDD1.n118 0.155672
R2580 VDD1.n150 VDD1.n118 0.155672
R2581 VDD1.n151 VDD1.n150 0.155672
R2582 VDD1.n151 VDD1.n114 0.155672
R2583 VDD1.n158 VDD1.n114 0.155672
R2584 VDD1.n159 VDD1.n158 0.155672
R2585 VDD1.n159 VDD1.n110 0.155672
R2586 VDD1.n166 VDD1.n110 0.155672
R2587 VDD1.n167 VDD1.n166 0.155672
R2588 VDD1.n167 VDD1.n106 0.155672
R2589 VDD1.n176 VDD1.n106 0.155672
R2590 VDD1.n177 VDD1.n176 0.155672
R2591 VDD1.n177 VDD1.n102 0.155672
R2592 VDD1.n184 VDD1.n102 0.155672
R2593 VDD1.n185 VDD1.n184 0.155672
R2594 VDD1.n185 VDD1.n98 0.155672
R2595 VDD1.n192 VDD1.n98 0.155672
R2596 VDD1 VDD1.n197 0.103948
C0 VTAIL VDD1 16.8916f
C1 VP VTAIL 4.02843f
C2 VTAIL VDD2 16.919f
C3 VN VDD1 0.147401f
C4 VP VN 5.81328f
C5 VN VDD2 4.644259f
C6 VN VTAIL 4.01345f
C7 VP VDD1 4.76439f
C8 VDD1 VDD2 0.613274f
C9 VP VDD2 0.274608f
C10 VDD2 B 5.260126f
C11 VDD1 B 5.225859f
C12 VTAIL B 8.03933f
C13 VN B 7.8097f
C14 VP B 5.284657f
C15 VDD1.n0 B 0.033885f
C16 VDD1.n1 B 0.025844f
C17 VDD1.n2 B 0.013887f
C18 VDD1.n3 B 0.032825f
C19 VDD1.n4 B 0.014704f
C20 VDD1.n5 B 0.025844f
C21 VDD1.n6 B 0.013887f
C22 VDD1.n7 B 0.032825f
C23 VDD1.n8 B 0.014296f
C24 VDD1.n9 B 0.025844f
C25 VDD1.n10 B 0.014296f
C26 VDD1.n11 B 0.013887f
C27 VDD1.n12 B 0.032825f
C28 VDD1.n13 B 0.032825f
C29 VDD1.n14 B 0.014704f
C30 VDD1.n15 B 0.025844f
C31 VDD1.n16 B 0.013887f
C32 VDD1.n17 B 0.032825f
C33 VDD1.n18 B 0.014704f
C34 VDD1.n19 B 0.025844f
C35 VDD1.n20 B 0.013887f
C36 VDD1.n21 B 0.032825f
C37 VDD1.n22 B 0.014704f
C38 VDD1.n23 B 0.025844f
C39 VDD1.n24 B 0.013887f
C40 VDD1.n25 B 0.032825f
C41 VDD1.n26 B 0.014704f
C42 VDD1.n27 B 0.025844f
C43 VDD1.n28 B 0.013887f
C44 VDD1.n29 B 0.032825f
C45 VDD1.n30 B 0.014704f
C46 VDD1.n31 B 1.96808f
C47 VDD1.n32 B 0.013887f
C48 VDD1.t5 B 0.054339f
C49 VDD1.n33 B 0.184241f
C50 VDD1.n34 B 0.019391f
C51 VDD1.n35 B 0.024619f
C52 VDD1.n36 B 0.032825f
C53 VDD1.n37 B 0.014704f
C54 VDD1.n38 B 0.013887f
C55 VDD1.n39 B 0.025844f
C56 VDD1.n40 B 0.025844f
C57 VDD1.n41 B 0.013887f
C58 VDD1.n42 B 0.014704f
C59 VDD1.n43 B 0.032825f
C60 VDD1.n44 B 0.032825f
C61 VDD1.n45 B 0.014704f
C62 VDD1.n46 B 0.013887f
C63 VDD1.n47 B 0.025844f
C64 VDD1.n48 B 0.025844f
C65 VDD1.n49 B 0.013887f
C66 VDD1.n50 B 0.014704f
C67 VDD1.n51 B 0.032825f
C68 VDD1.n52 B 0.032825f
C69 VDD1.n53 B 0.014704f
C70 VDD1.n54 B 0.013887f
C71 VDD1.n55 B 0.025844f
C72 VDD1.n56 B 0.025844f
C73 VDD1.n57 B 0.013887f
C74 VDD1.n58 B 0.014704f
C75 VDD1.n59 B 0.032825f
C76 VDD1.n60 B 0.032825f
C77 VDD1.n61 B 0.014704f
C78 VDD1.n62 B 0.013887f
C79 VDD1.n63 B 0.025844f
C80 VDD1.n64 B 0.025844f
C81 VDD1.n65 B 0.013887f
C82 VDD1.n66 B 0.014704f
C83 VDD1.n67 B 0.032825f
C84 VDD1.n68 B 0.032825f
C85 VDD1.n69 B 0.014704f
C86 VDD1.n70 B 0.013887f
C87 VDD1.n71 B 0.025844f
C88 VDD1.n72 B 0.025844f
C89 VDD1.n73 B 0.013887f
C90 VDD1.n74 B 0.014704f
C91 VDD1.n75 B 0.032825f
C92 VDD1.n76 B 0.032825f
C93 VDD1.n77 B 0.014704f
C94 VDD1.n78 B 0.013887f
C95 VDD1.n79 B 0.025844f
C96 VDD1.n80 B 0.025844f
C97 VDD1.n81 B 0.013887f
C98 VDD1.n82 B 0.014704f
C99 VDD1.n83 B 0.032825f
C100 VDD1.n84 B 0.032825f
C101 VDD1.n85 B 0.014704f
C102 VDD1.n86 B 0.013887f
C103 VDD1.n87 B 0.025844f
C104 VDD1.n88 B 0.025844f
C105 VDD1.n89 B 0.013887f
C106 VDD1.n90 B 0.014704f
C107 VDD1.n91 B 0.032825f
C108 VDD1.n92 B 0.066743f
C109 VDD1.n93 B 0.014704f
C110 VDD1.n94 B 0.013887f
C111 VDD1.n95 B 0.056206f
C112 VDD1.n96 B 0.055729f
C113 VDD1.n97 B 0.033885f
C114 VDD1.n98 B 0.025844f
C115 VDD1.n99 B 0.013887f
C116 VDD1.n100 B 0.032825f
C117 VDD1.n101 B 0.014704f
C118 VDD1.n102 B 0.025844f
C119 VDD1.n103 B 0.013887f
C120 VDD1.n104 B 0.032825f
C121 VDD1.n105 B 0.014296f
C122 VDD1.n106 B 0.025844f
C123 VDD1.n107 B 0.014704f
C124 VDD1.n108 B 0.032825f
C125 VDD1.n109 B 0.014704f
C126 VDD1.n110 B 0.025844f
C127 VDD1.n111 B 0.013887f
C128 VDD1.n112 B 0.032825f
C129 VDD1.n113 B 0.014704f
C130 VDD1.n114 B 0.025844f
C131 VDD1.n115 B 0.013887f
C132 VDD1.n116 B 0.032825f
C133 VDD1.n117 B 0.014704f
C134 VDD1.n118 B 0.025844f
C135 VDD1.n119 B 0.013887f
C136 VDD1.n120 B 0.032825f
C137 VDD1.n121 B 0.014704f
C138 VDD1.n122 B 0.025844f
C139 VDD1.n123 B 0.013887f
C140 VDD1.n124 B 0.032825f
C141 VDD1.n125 B 0.014704f
C142 VDD1.n126 B 1.96808f
C143 VDD1.n127 B 0.013887f
C144 VDD1.t3 B 0.054339f
C145 VDD1.n128 B 0.184241f
C146 VDD1.n129 B 0.019391f
C147 VDD1.n130 B 0.024619f
C148 VDD1.n131 B 0.032825f
C149 VDD1.n132 B 0.014704f
C150 VDD1.n133 B 0.013887f
C151 VDD1.n134 B 0.025844f
C152 VDD1.n135 B 0.025844f
C153 VDD1.n136 B 0.013887f
C154 VDD1.n137 B 0.014704f
C155 VDD1.n138 B 0.032825f
C156 VDD1.n139 B 0.032825f
C157 VDD1.n140 B 0.014704f
C158 VDD1.n141 B 0.013887f
C159 VDD1.n142 B 0.025844f
C160 VDD1.n143 B 0.025844f
C161 VDD1.n144 B 0.013887f
C162 VDD1.n145 B 0.014704f
C163 VDD1.n146 B 0.032825f
C164 VDD1.n147 B 0.032825f
C165 VDD1.n148 B 0.014704f
C166 VDD1.n149 B 0.013887f
C167 VDD1.n150 B 0.025844f
C168 VDD1.n151 B 0.025844f
C169 VDD1.n152 B 0.013887f
C170 VDD1.n153 B 0.014704f
C171 VDD1.n154 B 0.032825f
C172 VDD1.n155 B 0.032825f
C173 VDD1.n156 B 0.014704f
C174 VDD1.n157 B 0.013887f
C175 VDD1.n158 B 0.025844f
C176 VDD1.n159 B 0.025844f
C177 VDD1.n160 B 0.013887f
C178 VDD1.n161 B 0.014704f
C179 VDD1.n162 B 0.032825f
C180 VDD1.n163 B 0.032825f
C181 VDD1.n164 B 0.014704f
C182 VDD1.n165 B 0.013887f
C183 VDD1.n166 B 0.025844f
C184 VDD1.n167 B 0.025844f
C185 VDD1.n168 B 0.013887f
C186 VDD1.n169 B 0.013887f
C187 VDD1.n170 B 0.014704f
C188 VDD1.n171 B 0.032825f
C189 VDD1.n172 B 0.032825f
C190 VDD1.n173 B 0.032825f
C191 VDD1.n174 B 0.014296f
C192 VDD1.n175 B 0.013887f
C193 VDD1.n176 B 0.025844f
C194 VDD1.n177 B 0.025844f
C195 VDD1.n178 B 0.013887f
C196 VDD1.n179 B 0.014704f
C197 VDD1.n180 B 0.032825f
C198 VDD1.n181 B 0.032825f
C199 VDD1.n182 B 0.014704f
C200 VDD1.n183 B 0.013887f
C201 VDD1.n184 B 0.025844f
C202 VDD1.n185 B 0.025844f
C203 VDD1.n186 B 0.013887f
C204 VDD1.n187 B 0.014704f
C205 VDD1.n188 B 0.032825f
C206 VDD1.n189 B 0.066743f
C207 VDD1.n190 B 0.014704f
C208 VDD1.n191 B 0.013887f
C209 VDD1.n192 B 0.056206f
C210 VDD1.n193 B 0.055435f
C211 VDD1.t4 B 0.355763f
C212 VDD1.t1 B 0.355763f
C213 VDD1.n194 B 3.23427f
C214 VDD1.n195 B 2.20997f
C215 VDD1.t0 B 0.355763f
C216 VDD1.t2 B 0.355763f
C217 VDD1.n196 B 3.23374f
C218 VDD1.n197 B 2.68373f
C219 VP.n0 B 0.054436f
C220 VP.t2 B 1.13227f
C221 VP.t0 B 1.13952f
C222 VP.n1 B 0.425992f
C223 VP.t5 B 1.13003f
C224 VP.n2 B 0.442127f
C225 VP.t3 B 1.13227f
C226 VP.n3 B 0.432834f
C227 VP.n4 B 2.57521f
C228 VP.n5 B 2.49668f
C229 VP.n6 B 0.432834f
C230 VP.t1 B 1.13003f
C231 VP.n7 B 0.442127f
C232 VP.t4 B 1.13227f
C233 VP.n8 B 0.432834f
C234 VP.n9 B 0.042186f
C235 VDD2.n0 B 0.033721f
C236 VDD2.n1 B 0.025719f
C237 VDD2.n2 B 0.01382f
C238 VDD2.n3 B 0.032666f
C239 VDD2.n4 B 0.014633f
C240 VDD2.n5 B 0.025719f
C241 VDD2.n6 B 0.01382f
C242 VDD2.n7 B 0.032666f
C243 VDD2.n8 B 0.014227f
C244 VDD2.n9 B 0.025719f
C245 VDD2.n10 B 0.014633f
C246 VDD2.n11 B 0.032666f
C247 VDD2.n12 B 0.014633f
C248 VDD2.n13 B 0.025719f
C249 VDD2.n14 B 0.01382f
C250 VDD2.n15 B 0.032666f
C251 VDD2.n16 B 0.014633f
C252 VDD2.n17 B 0.025719f
C253 VDD2.n18 B 0.01382f
C254 VDD2.n19 B 0.032666f
C255 VDD2.n20 B 0.014633f
C256 VDD2.n21 B 0.025719f
C257 VDD2.n22 B 0.01382f
C258 VDD2.n23 B 0.032666f
C259 VDD2.n24 B 0.014633f
C260 VDD2.n25 B 0.025719f
C261 VDD2.n26 B 0.01382f
C262 VDD2.n27 B 0.032666f
C263 VDD2.n28 B 0.014633f
C264 VDD2.n29 B 1.95855f
C265 VDD2.n30 B 0.01382f
C266 VDD2.t3 B 0.054076f
C267 VDD2.n31 B 0.183349f
C268 VDD2.n32 B 0.019297f
C269 VDD2.n33 B 0.0245f
C270 VDD2.n34 B 0.032666f
C271 VDD2.n35 B 0.014633f
C272 VDD2.n36 B 0.01382f
C273 VDD2.n37 B 0.025719f
C274 VDD2.n38 B 0.025719f
C275 VDD2.n39 B 0.01382f
C276 VDD2.n40 B 0.014633f
C277 VDD2.n41 B 0.032666f
C278 VDD2.n42 B 0.032666f
C279 VDD2.n43 B 0.014633f
C280 VDD2.n44 B 0.01382f
C281 VDD2.n45 B 0.025719f
C282 VDD2.n46 B 0.025719f
C283 VDD2.n47 B 0.01382f
C284 VDD2.n48 B 0.014633f
C285 VDD2.n49 B 0.032666f
C286 VDD2.n50 B 0.032666f
C287 VDD2.n51 B 0.014633f
C288 VDD2.n52 B 0.01382f
C289 VDD2.n53 B 0.025719f
C290 VDD2.n54 B 0.025719f
C291 VDD2.n55 B 0.01382f
C292 VDD2.n56 B 0.014633f
C293 VDD2.n57 B 0.032666f
C294 VDD2.n58 B 0.032666f
C295 VDD2.n59 B 0.014633f
C296 VDD2.n60 B 0.01382f
C297 VDD2.n61 B 0.025719f
C298 VDD2.n62 B 0.025719f
C299 VDD2.n63 B 0.01382f
C300 VDD2.n64 B 0.014633f
C301 VDD2.n65 B 0.032666f
C302 VDD2.n66 B 0.032666f
C303 VDD2.n67 B 0.014633f
C304 VDD2.n68 B 0.01382f
C305 VDD2.n69 B 0.025719f
C306 VDD2.n70 B 0.025719f
C307 VDD2.n71 B 0.01382f
C308 VDD2.n72 B 0.01382f
C309 VDD2.n73 B 0.014633f
C310 VDD2.n74 B 0.032666f
C311 VDD2.n75 B 0.032666f
C312 VDD2.n76 B 0.032666f
C313 VDD2.n77 B 0.014227f
C314 VDD2.n78 B 0.01382f
C315 VDD2.n79 B 0.025719f
C316 VDD2.n80 B 0.025719f
C317 VDD2.n81 B 0.01382f
C318 VDD2.n82 B 0.014633f
C319 VDD2.n83 B 0.032666f
C320 VDD2.n84 B 0.032666f
C321 VDD2.n85 B 0.014633f
C322 VDD2.n86 B 0.01382f
C323 VDD2.n87 B 0.025719f
C324 VDD2.n88 B 0.025719f
C325 VDD2.n89 B 0.01382f
C326 VDD2.n90 B 0.014633f
C327 VDD2.n91 B 0.032666f
C328 VDD2.n92 B 0.06642f
C329 VDD2.n93 B 0.014633f
C330 VDD2.n94 B 0.01382f
C331 VDD2.n95 B 0.055935f
C332 VDD2.n96 B 0.055167f
C333 VDD2.t0 B 0.354041f
C334 VDD2.t5 B 0.354041f
C335 VDD2.n97 B 3.21862f
C336 VDD2.n98 B 2.12552f
C337 VDD2.n99 B 0.033721f
C338 VDD2.n100 B 0.025719f
C339 VDD2.n101 B 0.01382f
C340 VDD2.n102 B 0.032666f
C341 VDD2.n103 B 0.014633f
C342 VDD2.n104 B 0.025719f
C343 VDD2.n105 B 0.01382f
C344 VDD2.n106 B 0.032666f
C345 VDD2.n107 B 0.014227f
C346 VDD2.n108 B 0.025719f
C347 VDD2.n109 B 0.014227f
C348 VDD2.n110 B 0.01382f
C349 VDD2.n111 B 0.032666f
C350 VDD2.n112 B 0.032666f
C351 VDD2.n113 B 0.014633f
C352 VDD2.n114 B 0.025719f
C353 VDD2.n115 B 0.01382f
C354 VDD2.n116 B 0.032666f
C355 VDD2.n117 B 0.014633f
C356 VDD2.n118 B 0.025719f
C357 VDD2.n119 B 0.01382f
C358 VDD2.n120 B 0.032666f
C359 VDD2.n121 B 0.014633f
C360 VDD2.n122 B 0.025719f
C361 VDD2.n123 B 0.01382f
C362 VDD2.n124 B 0.032666f
C363 VDD2.n125 B 0.014633f
C364 VDD2.n126 B 0.025719f
C365 VDD2.n127 B 0.01382f
C366 VDD2.n128 B 0.032666f
C367 VDD2.n129 B 0.014633f
C368 VDD2.n130 B 1.95855f
C369 VDD2.n131 B 0.01382f
C370 VDD2.t1 B 0.054076f
C371 VDD2.n132 B 0.183349f
C372 VDD2.n133 B 0.019297f
C373 VDD2.n134 B 0.0245f
C374 VDD2.n135 B 0.032666f
C375 VDD2.n136 B 0.014633f
C376 VDD2.n137 B 0.01382f
C377 VDD2.n138 B 0.025719f
C378 VDD2.n139 B 0.025719f
C379 VDD2.n140 B 0.01382f
C380 VDD2.n141 B 0.014633f
C381 VDD2.n142 B 0.032666f
C382 VDD2.n143 B 0.032666f
C383 VDD2.n144 B 0.014633f
C384 VDD2.n145 B 0.01382f
C385 VDD2.n146 B 0.025719f
C386 VDD2.n147 B 0.025719f
C387 VDD2.n148 B 0.01382f
C388 VDD2.n149 B 0.014633f
C389 VDD2.n150 B 0.032666f
C390 VDD2.n151 B 0.032666f
C391 VDD2.n152 B 0.014633f
C392 VDD2.n153 B 0.01382f
C393 VDD2.n154 B 0.025719f
C394 VDD2.n155 B 0.025719f
C395 VDD2.n156 B 0.01382f
C396 VDD2.n157 B 0.014633f
C397 VDD2.n158 B 0.032666f
C398 VDD2.n159 B 0.032666f
C399 VDD2.n160 B 0.014633f
C400 VDD2.n161 B 0.01382f
C401 VDD2.n162 B 0.025719f
C402 VDD2.n163 B 0.025719f
C403 VDD2.n164 B 0.01382f
C404 VDD2.n165 B 0.014633f
C405 VDD2.n166 B 0.032666f
C406 VDD2.n167 B 0.032666f
C407 VDD2.n168 B 0.014633f
C408 VDD2.n169 B 0.01382f
C409 VDD2.n170 B 0.025719f
C410 VDD2.n171 B 0.025719f
C411 VDD2.n172 B 0.01382f
C412 VDD2.n173 B 0.014633f
C413 VDD2.n174 B 0.032666f
C414 VDD2.n175 B 0.032666f
C415 VDD2.n176 B 0.014633f
C416 VDD2.n177 B 0.01382f
C417 VDD2.n178 B 0.025719f
C418 VDD2.n179 B 0.025719f
C419 VDD2.n180 B 0.01382f
C420 VDD2.n181 B 0.014633f
C421 VDD2.n182 B 0.032666f
C422 VDD2.n183 B 0.032666f
C423 VDD2.n184 B 0.014633f
C424 VDD2.n185 B 0.01382f
C425 VDD2.n186 B 0.025719f
C426 VDD2.n187 B 0.025719f
C427 VDD2.n188 B 0.01382f
C428 VDD2.n189 B 0.014633f
C429 VDD2.n190 B 0.032666f
C430 VDD2.n191 B 0.06642f
C431 VDD2.n192 B 0.014633f
C432 VDD2.n193 B 0.01382f
C433 VDD2.n194 B 0.055935f
C434 VDD2.n195 B 0.054401f
C435 VDD2.n196 B 2.4534f
C436 VDD2.t4 B 0.354041f
C437 VDD2.t2 B 0.354041f
C438 VDD2.n197 B 3.2186f
C439 VTAIL.t4 B 0.358527f
C440 VTAIL.t3 B 0.358527f
C441 VTAIL.n0 B 3.17405f
C442 VTAIL.n1 B 0.353265f
C443 VTAIL.n2 B 0.034148f
C444 VTAIL.n3 B 0.026045f
C445 VTAIL.n4 B 0.013995f
C446 VTAIL.n5 B 0.03308f
C447 VTAIL.n6 B 0.014819f
C448 VTAIL.n7 B 0.026045f
C449 VTAIL.n8 B 0.013995f
C450 VTAIL.n9 B 0.03308f
C451 VTAIL.n10 B 0.014407f
C452 VTAIL.n11 B 0.026045f
C453 VTAIL.n12 B 0.014819f
C454 VTAIL.n13 B 0.03308f
C455 VTAIL.n14 B 0.014819f
C456 VTAIL.n15 B 0.026045f
C457 VTAIL.n16 B 0.013995f
C458 VTAIL.n17 B 0.03308f
C459 VTAIL.n18 B 0.014819f
C460 VTAIL.n19 B 0.026045f
C461 VTAIL.n20 B 0.013995f
C462 VTAIL.n21 B 0.03308f
C463 VTAIL.n22 B 0.014819f
C464 VTAIL.n23 B 0.026045f
C465 VTAIL.n24 B 0.013995f
C466 VTAIL.n25 B 0.03308f
C467 VTAIL.n26 B 0.014819f
C468 VTAIL.n27 B 0.026045f
C469 VTAIL.n28 B 0.013995f
C470 VTAIL.n29 B 0.03308f
C471 VTAIL.n30 B 0.014819f
C472 VTAIL.n31 B 1.98337f
C473 VTAIL.n32 B 0.013995f
C474 VTAIL.t1 B 0.054761f
C475 VTAIL.n33 B 0.185672f
C476 VTAIL.n34 B 0.019541f
C477 VTAIL.n35 B 0.02481f
C478 VTAIL.n36 B 0.03308f
C479 VTAIL.n37 B 0.014819f
C480 VTAIL.n38 B 0.013995f
C481 VTAIL.n39 B 0.026045f
C482 VTAIL.n40 B 0.026045f
C483 VTAIL.n41 B 0.013995f
C484 VTAIL.n42 B 0.014819f
C485 VTAIL.n43 B 0.03308f
C486 VTAIL.n44 B 0.03308f
C487 VTAIL.n45 B 0.014819f
C488 VTAIL.n46 B 0.013995f
C489 VTAIL.n47 B 0.026045f
C490 VTAIL.n48 B 0.026045f
C491 VTAIL.n49 B 0.013995f
C492 VTAIL.n50 B 0.014819f
C493 VTAIL.n51 B 0.03308f
C494 VTAIL.n52 B 0.03308f
C495 VTAIL.n53 B 0.014819f
C496 VTAIL.n54 B 0.013995f
C497 VTAIL.n55 B 0.026045f
C498 VTAIL.n56 B 0.026045f
C499 VTAIL.n57 B 0.013995f
C500 VTAIL.n58 B 0.014819f
C501 VTAIL.n59 B 0.03308f
C502 VTAIL.n60 B 0.03308f
C503 VTAIL.n61 B 0.014819f
C504 VTAIL.n62 B 0.013995f
C505 VTAIL.n63 B 0.026045f
C506 VTAIL.n64 B 0.026045f
C507 VTAIL.n65 B 0.013995f
C508 VTAIL.n66 B 0.014819f
C509 VTAIL.n67 B 0.03308f
C510 VTAIL.n68 B 0.03308f
C511 VTAIL.n69 B 0.014819f
C512 VTAIL.n70 B 0.013995f
C513 VTAIL.n71 B 0.026045f
C514 VTAIL.n72 B 0.026045f
C515 VTAIL.n73 B 0.013995f
C516 VTAIL.n74 B 0.013995f
C517 VTAIL.n75 B 0.014819f
C518 VTAIL.n76 B 0.03308f
C519 VTAIL.n77 B 0.03308f
C520 VTAIL.n78 B 0.03308f
C521 VTAIL.n79 B 0.014407f
C522 VTAIL.n80 B 0.013995f
C523 VTAIL.n81 B 0.026045f
C524 VTAIL.n82 B 0.026045f
C525 VTAIL.n83 B 0.013995f
C526 VTAIL.n84 B 0.014819f
C527 VTAIL.n85 B 0.03308f
C528 VTAIL.n86 B 0.03308f
C529 VTAIL.n87 B 0.014819f
C530 VTAIL.n88 B 0.013995f
C531 VTAIL.n89 B 0.026045f
C532 VTAIL.n90 B 0.026045f
C533 VTAIL.n91 B 0.013995f
C534 VTAIL.n92 B 0.014819f
C535 VTAIL.n93 B 0.03308f
C536 VTAIL.n94 B 0.067262f
C537 VTAIL.n95 B 0.014819f
C538 VTAIL.n96 B 0.013995f
C539 VTAIL.n97 B 0.056643f
C540 VTAIL.n98 B 0.037076f
C541 VTAIL.n99 B 0.141058f
C542 VTAIL.t0 B 0.358527f
C543 VTAIL.t10 B 0.358527f
C544 VTAIL.n100 B 3.17405f
C545 VTAIL.n101 B 2.0451f
C546 VTAIL.t5 B 0.358527f
C547 VTAIL.t7 B 0.358527f
C548 VTAIL.n102 B 3.17407f
C549 VTAIL.n103 B 2.04508f
C550 VTAIL.n104 B 0.034148f
C551 VTAIL.n105 B 0.026045f
C552 VTAIL.n106 B 0.013995f
C553 VTAIL.n107 B 0.03308f
C554 VTAIL.n108 B 0.014819f
C555 VTAIL.n109 B 0.026045f
C556 VTAIL.n110 B 0.013995f
C557 VTAIL.n111 B 0.03308f
C558 VTAIL.n112 B 0.014407f
C559 VTAIL.n113 B 0.026045f
C560 VTAIL.n114 B 0.014407f
C561 VTAIL.n115 B 0.013995f
C562 VTAIL.n116 B 0.03308f
C563 VTAIL.n117 B 0.03308f
C564 VTAIL.n118 B 0.014819f
C565 VTAIL.n119 B 0.026045f
C566 VTAIL.n120 B 0.013995f
C567 VTAIL.n121 B 0.03308f
C568 VTAIL.n122 B 0.014819f
C569 VTAIL.n123 B 0.026045f
C570 VTAIL.n124 B 0.013995f
C571 VTAIL.n125 B 0.03308f
C572 VTAIL.n126 B 0.014819f
C573 VTAIL.n127 B 0.026045f
C574 VTAIL.n128 B 0.013995f
C575 VTAIL.n129 B 0.03308f
C576 VTAIL.n130 B 0.014819f
C577 VTAIL.n131 B 0.026045f
C578 VTAIL.n132 B 0.013995f
C579 VTAIL.n133 B 0.03308f
C580 VTAIL.n134 B 0.014819f
C581 VTAIL.n135 B 1.98337f
C582 VTAIL.n136 B 0.013995f
C583 VTAIL.t2 B 0.054761f
C584 VTAIL.n137 B 0.185672f
C585 VTAIL.n138 B 0.019541f
C586 VTAIL.n139 B 0.02481f
C587 VTAIL.n140 B 0.03308f
C588 VTAIL.n141 B 0.014819f
C589 VTAIL.n142 B 0.013995f
C590 VTAIL.n143 B 0.026045f
C591 VTAIL.n144 B 0.026045f
C592 VTAIL.n145 B 0.013995f
C593 VTAIL.n146 B 0.014819f
C594 VTAIL.n147 B 0.03308f
C595 VTAIL.n148 B 0.03308f
C596 VTAIL.n149 B 0.014819f
C597 VTAIL.n150 B 0.013995f
C598 VTAIL.n151 B 0.026045f
C599 VTAIL.n152 B 0.026045f
C600 VTAIL.n153 B 0.013995f
C601 VTAIL.n154 B 0.014819f
C602 VTAIL.n155 B 0.03308f
C603 VTAIL.n156 B 0.03308f
C604 VTAIL.n157 B 0.014819f
C605 VTAIL.n158 B 0.013995f
C606 VTAIL.n159 B 0.026045f
C607 VTAIL.n160 B 0.026045f
C608 VTAIL.n161 B 0.013995f
C609 VTAIL.n162 B 0.014819f
C610 VTAIL.n163 B 0.03308f
C611 VTAIL.n164 B 0.03308f
C612 VTAIL.n165 B 0.014819f
C613 VTAIL.n166 B 0.013995f
C614 VTAIL.n167 B 0.026045f
C615 VTAIL.n168 B 0.026045f
C616 VTAIL.n169 B 0.013995f
C617 VTAIL.n170 B 0.014819f
C618 VTAIL.n171 B 0.03308f
C619 VTAIL.n172 B 0.03308f
C620 VTAIL.n173 B 0.014819f
C621 VTAIL.n174 B 0.013995f
C622 VTAIL.n175 B 0.026045f
C623 VTAIL.n176 B 0.026045f
C624 VTAIL.n177 B 0.013995f
C625 VTAIL.n178 B 0.014819f
C626 VTAIL.n179 B 0.03308f
C627 VTAIL.n180 B 0.03308f
C628 VTAIL.n181 B 0.014819f
C629 VTAIL.n182 B 0.013995f
C630 VTAIL.n183 B 0.026045f
C631 VTAIL.n184 B 0.026045f
C632 VTAIL.n185 B 0.013995f
C633 VTAIL.n186 B 0.014819f
C634 VTAIL.n187 B 0.03308f
C635 VTAIL.n188 B 0.03308f
C636 VTAIL.n189 B 0.014819f
C637 VTAIL.n190 B 0.013995f
C638 VTAIL.n191 B 0.026045f
C639 VTAIL.n192 B 0.026045f
C640 VTAIL.n193 B 0.013995f
C641 VTAIL.n194 B 0.014819f
C642 VTAIL.n195 B 0.03308f
C643 VTAIL.n196 B 0.067262f
C644 VTAIL.n197 B 0.014819f
C645 VTAIL.n198 B 0.013995f
C646 VTAIL.n199 B 0.056643f
C647 VTAIL.n200 B 0.037076f
C648 VTAIL.n201 B 0.141058f
C649 VTAIL.t11 B 0.358527f
C650 VTAIL.t8 B 0.358527f
C651 VTAIL.n202 B 3.17407f
C652 VTAIL.n203 B 0.389061f
C653 VTAIL.n204 B 0.034148f
C654 VTAIL.n205 B 0.026045f
C655 VTAIL.n206 B 0.013995f
C656 VTAIL.n207 B 0.03308f
C657 VTAIL.n208 B 0.014819f
C658 VTAIL.n209 B 0.026045f
C659 VTAIL.n210 B 0.013995f
C660 VTAIL.n211 B 0.03308f
C661 VTAIL.n212 B 0.014407f
C662 VTAIL.n213 B 0.026045f
C663 VTAIL.n214 B 0.014407f
C664 VTAIL.n215 B 0.013995f
C665 VTAIL.n216 B 0.03308f
C666 VTAIL.n217 B 0.03308f
C667 VTAIL.n218 B 0.014819f
C668 VTAIL.n219 B 0.026045f
C669 VTAIL.n220 B 0.013995f
C670 VTAIL.n221 B 0.03308f
C671 VTAIL.n222 B 0.014819f
C672 VTAIL.n223 B 0.026045f
C673 VTAIL.n224 B 0.013995f
C674 VTAIL.n225 B 0.03308f
C675 VTAIL.n226 B 0.014819f
C676 VTAIL.n227 B 0.026045f
C677 VTAIL.n228 B 0.013995f
C678 VTAIL.n229 B 0.03308f
C679 VTAIL.n230 B 0.014819f
C680 VTAIL.n231 B 0.026045f
C681 VTAIL.n232 B 0.013995f
C682 VTAIL.n233 B 0.03308f
C683 VTAIL.n234 B 0.014819f
C684 VTAIL.n235 B 1.98337f
C685 VTAIL.n236 B 0.013995f
C686 VTAIL.t9 B 0.054761f
C687 VTAIL.n237 B 0.185672f
C688 VTAIL.n238 B 0.019541f
C689 VTAIL.n239 B 0.02481f
C690 VTAIL.n240 B 0.03308f
C691 VTAIL.n241 B 0.014819f
C692 VTAIL.n242 B 0.013995f
C693 VTAIL.n243 B 0.026045f
C694 VTAIL.n244 B 0.026045f
C695 VTAIL.n245 B 0.013995f
C696 VTAIL.n246 B 0.014819f
C697 VTAIL.n247 B 0.03308f
C698 VTAIL.n248 B 0.03308f
C699 VTAIL.n249 B 0.014819f
C700 VTAIL.n250 B 0.013995f
C701 VTAIL.n251 B 0.026045f
C702 VTAIL.n252 B 0.026045f
C703 VTAIL.n253 B 0.013995f
C704 VTAIL.n254 B 0.014819f
C705 VTAIL.n255 B 0.03308f
C706 VTAIL.n256 B 0.03308f
C707 VTAIL.n257 B 0.014819f
C708 VTAIL.n258 B 0.013995f
C709 VTAIL.n259 B 0.026045f
C710 VTAIL.n260 B 0.026045f
C711 VTAIL.n261 B 0.013995f
C712 VTAIL.n262 B 0.014819f
C713 VTAIL.n263 B 0.03308f
C714 VTAIL.n264 B 0.03308f
C715 VTAIL.n265 B 0.014819f
C716 VTAIL.n266 B 0.013995f
C717 VTAIL.n267 B 0.026045f
C718 VTAIL.n268 B 0.026045f
C719 VTAIL.n269 B 0.013995f
C720 VTAIL.n270 B 0.014819f
C721 VTAIL.n271 B 0.03308f
C722 VTAIL.n272 B 0.03308f
C723 VTAIL.n273 B 0.014819f
C724 VTAIL.n274 B 0.013995f
C725 VTAIL.n275 B 0.026045f
C726 VTAIL.n276 B 0.026045f
C727 VTAIL.n277 B 0.013995f
C728 VTAIL.n278 B 0.014819f
C729 VTAIL.n279 B 0.03308f
C730 VTAIL.n280 B 0.03308f
C731 VTAIL.n281 B 0.014819f
C732 VTAIL.n282 B 0.013995f
C733 VTAIL.n283 B 0.026045f
C734 VTAIL.n284 B 0.026045f
C735 VTAIL.n285 B 0.013995f
C736 VTAIL.n286 B 0.014819f
C737 VTAIL.n287 B 0.03308f
C738 VTAIL.n288 B 0.03308f
C739 VTAIL.n289 B 0.014819f
C740 VTAIL.n290 B 0.013995f
C741 VTAIL.n291 B 0.026045f
C742 VTAIL.n292 B 0.026045f
C743 VTAIL.n293 B 0.013995f
C744 VTAIL.n294 B 0.014819f
C745 VTAIL.n295 B 0.03308f
C746 VTAIL.n296 B 0.067262f
C747 VTAIL.n297 B 0.014819f
C748 VTAIL.n298 B 0.013995f
C749 VTAIL.n299 B 0.056643f
C750 VTAIL.n300 B 0.037076f
C751 VTAIL.n301 B 1.74282f
C752 VTAIL.n302 B 0.034148f
C753 VTAIL.n303 B 0.026045f
C754 VTAIL.n304 B 0.013995f
C755 VTAIL.n305 B 0.03308f
C756 VTAIL.n306 B 0.014819f
C757 VTAIL.n307 B 0.026045f
C758 VTAIL.n308 B 0.013995f
C759 VTAIL.n309 B 0.03308f
C760 VTAIL.n310 B 0.014407f
C761 VTAIL.n311 B 0.026045f
C762 VTAIL.n312 B 0.014819f
C763 VTAIL.n313 B 0.03308f
C764 VTAIL.n314 B 0.014819f
C765 VTAIL.n315 B 0.026045f
C766 VTAIL.n316 B 0.013995f
C767 VTAIL.n317 B 0.03308f
C768 VTAIL.n318 B 0.014819f
C769 VTAIL.n319 B 0.026045f
C770 VTAIL.n320 B 0.013995f
C771 VTAIL.n321 B 0.03308f
C772 VTAIL.n322 B 0.014819f
C773 VTAIL.n323 B 0.026045f
C774 VTAIL.n324 B 0.013995f
C775 VTAIL.n325 B 0.03308f
C776 VTAIL.n326 B 0.014819f
C777 VTAIL.n327 B 0.026045f
C778 VTAIL.n328 B 0.013995f
C779 VTAIL.n329 B 0.03308f
C780 VTAIL.n330 B 0.014819f
C781 VTAIL.n331 B 1.98337f
C782 VTAIL.n332 B 0.013995f
C783 VTAIL.t6 B 0.054761f
C784 VTAIL.n333 B 0.185672f
C785 VTAIL.n334 B 0.019541f
C786 VTAIL.n335 B 0.02481f
C787 VTAIL.n336 B 0.03308f
C788 VTAIL.n337 B 0.014819f
C789 VTAIL.n338 B 0.013995f
C790 VTAIL.n339 B 0.026045f
C791 VTAIL.n340 B 0.026045f
C792 VTAIL.n341 B 0.013995f
C793 VTAIL.n342 B 0.014819f
C794 VTAIL.n343 B 0.03308f
C795 VTAIL.n344 B 0.03308f
C796 VTAIL.n345 B 0.014819f
C797 VTAIL.n346 B 0.013995f
C798 VTAIL.n347 B 0.026045f
C799 VTAIL.n348 B 0.026045f
C800 VTAIL.n349 B 0.013995f
C801 VTAIL.n350 B 0.014819f
C802 VTAIL.n351 B 0.03308f
C803 VTAIL.n352 B 0.03308f
C804 VTAIL.n353 B 0.014819f
C805 VTAIL.n354 B 0.013995f
C806 VTAIL.n355 B 0.026045f
C807 VTAIL.n356 B 0.026045f
C808 VTAIL.n357 B 0.013995f
C809 VTAIL.n358 B 0.014819f
C810 VTAIL.n359 B 0.03308f
C811 VTAIL.n360 B 0.03308f
C812 VTAIL.n361 B 0.014819f
C813 VTAIL.n362 B 0.013995f
C814 VTAIL.n363 B 0.026045f
C815 VTAIL.n364 B 0.026045f
C816 VTAIL.n365 B 0.013995f
C817 VTAIL.n366 B 0.014819f
C818 VTAIL.n367 B 0.03308f
C819 VTAIL.n368 B 0.03308f
C820 VTAIL.n369 B 0.014819f
C821 VTAIL.n370 B 0.013995f
C822 VTAIL.n371 B 0.026045f
C823 VTAIL.n372 B 0.026045f
C824 VTAIL.n373 B 0.013995f
C825 VTAIL.n374 B 0.013995f
C826 VTAIL.n375 B 0.014819f
C827 VTAIL.n376 B 0.03308f
C828 VTAIL.n377 B 0.03308f
C829 VTAIL.n378 B 0.03308f
C830 VTAIL.n379 B 0.014407f
C831 VTAIL.n380 B 0.013995f
C832 VTAIL.n381 B 0.026045f
C833 VTAIL.n382 B 0.026045f
C834 VTAIL.n383 B 0.013995f
C835 VTAIL.n384 B 0.014819f
C836 VTAIL.n385 B 0.03308f
C837 VTAIL.n386 B 0.03308f
C838 VTAIL.n387 B 0.014819f
C839 VTAIL.n388 B 0.013995f
C840 VTAIL.n389 B 0.026045f
C841 VTAIL.n390 B 0.026045f
C842 VTAIL.n391 B 0.013995f
C843 VTAIL.n392 B 0.014819f
C844 VTAIL.n393 B 0.03308f
C845 VTAIL.n394 B 0.067262f
C846 VTAIL.n395 B 0.014819f
C847 VTAIL.n396 B 0.013995f
C848 VTAIL.n397 B 0.056643f
C849 VTAIL.n398 B 0.037076f
C850 VTAIL.n399 B 1.72437f
C851 VN.t2 B 1.11805f
C852 VN.n0 B 0.417965f
C853 VN.t5 B 1.10874f
C854 VN.n1 B 0.433797f
C855 VN.t0 B 1.11094f
C856 VN.n2 B 0.424679f
C857 VN.n3 B 0.161643f
C858 VN.t3 B 1.11805f
C859 VN.n4 B 0.417965f
C860 VN.t4 B 1.11094f
C861 VN.t1 B 1.10874f
C862 VN.n5 B 0.433797f
C863 VN.n6 B 0.424679f
C864 VN.n7 B 2.56164f
.ends

