* NGSPICE file created from diff_pair_sample_1701.ext - technology: sky130A

.subckt diff_pair_sample_1701 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.109 pd=26.98 as=5.109 ps=26.98 w=13.1 l=3.5
X1 VDD1.t1 VP.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=5.109 pd=26.98 as=5.109 ps=26.98 w=13.1 l=3.5
X2 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=5.109 pd=26.98 as=0 ps=0 w=13.1 l=3.5
X3 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.109 pd=26.98 as=5.109 ps=26.98 w=13.1 l=3.5
X4 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=5.109 pd=26.98 as=0 ps=0 w=13.1 l=3.5
X5 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=5.109 pd=26.98 as=5.109 ps=26.98 w=13.1 l=3.5
X6 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=5.109 pd=26.98 as=0 ps=0 w=13.1 l=3.5
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=5.109 pd=26.98 as=0 ps=0 w=13.1 l=3.5
R0 VN VN.t1 176.833
R1 VN VN.t0 129.575
R2 VTAIL.n1 VTAIL.t2 44.5186
R3 VTAIL.n3 VTAIL.t1 44.5183
R4 VTAIL.n0 VTAIL.t0 44.5183
R5 VTAIL.n2 VTAIL.t3 44.5183
R6 VTAIL.n1 VTAIL.n0 30.2634
R7 VTAIL.n3 VTAIL.n2 26.9617
R8 VTAIL.n2 VTAIL.n1 2.12119
R9 VTAIL VTAIL.n0 1.35395
R10 VTAIL VTAIL.n3 0.767741
R11 VDD2.n0 VDD2.t1 102.754
R12 VDD2.n0 VDD2.t0 61.1971
R13 VDD2 VDD2.n0 0.884121
R14 B.n555 B.n113 585
R15 B.n113 B.n58 585
R16 B.n557 B.n556 585
R17 B.n559 B.n112 585
R18 B.n562 B.n561 585
R19 B.n563 B.n111 585
R20 B.n565 B.n564 585
R21 B.n567 B.n110 585
R22 B.n570 B.n569 585
R23 B.n571 B.n109 585
R24 B.n573 B.n572 585
R25 B.n575 B.n108 585
R26 B.n578 B.n577 585
R27 B.n579 B.n107 585
R28 B.n581 B.n580 585
R29 B.n583 B.n106 585
R30 B.n586 B.n585 585
R31 B.n587 B.n105 585
R32 B.n589 B.n588 585
R33 B.n591 B.n104 585
R34 B.n594 B.n593 585
R35 B.n595 B.n103 585
R36 B.n597 B.n596 585
R37 B.n599 B.n102 585
R38 B.n602 B.n601 585
R39 B.n603 B.n101 585
R40 B.n605 B.n604 585
R41 B.n607 B.n100 585
R42 B.n610 B.n609 585
R43 B.n611 B.n99 585
R44 B.n613 B.n612 585
R45 B.n615 B.n98 585
R46 B.n618 B.n617 585
R47 B.n619 B.n97 585
R48 B.n621 B.n620 585
R49 B.n623 B.n96 585
R50 B.n626 B.n625 585
R51 B.n627 B.n95 585
R52 B.n629 B.n628 585
R53 B.n631 B.n94 585
R54 B.n634 B.n633 585
R55 B.n635 B.n93 585
R56 B.n637 B.n636 585
R57 B.n639 B.n92 585
R58 B.n641 B.n640 585
R59 B.n643 B.n642 585
R60 B.n646 B.n645 585
R61 B.n647 B.n87 585
R62 B.n649 B.n648 585
R63 B.n651 B.n86 585
R64 B.n654 B.n653 585
R65 B.n655 B.n85 585
R66 B.n657 B.n656 585
R67 B.n659 B.n84 585
R68 B.n662 B.n661 585
R69 B.n664 B.n81 585
R70 B.n666 B.n665 585
R71 B.n668 B.n80 585
R72 B.n671 B.n670 585
R73 B.n672 B.n79 585
R74 B.n674 B.n673 585
R75 B.n676 B.n78 585
R76 B.n679 B.n678 585
R77 B.n680 B.n77 585
R78 B.n682 B.n681 585
R79 B.n684 B.n76 585
R80 B.n687 B.n686 585
R81 B.n688 B.n75 585
R82 B.n690 B.n689 585
R83 B.n692 B.n74 585
R84 B.n695 B.n694 585
R85 B.n696 B.n73 585
R86 B.n698 B.n697 585
R87 B.n700 B.n72 585
R88 B.n703 B.n702 585
R89 B.n704 B.n71 585
R90 B.n706 B.n705 585
R91 B.n708 B.n70 585
R92 B.n711 B.n710 585
R93 B.n712 B.n69 585
R94 B.n714 B.n713 585
R95 B.n716 B.n68 585
R96 B.n719 B.n718 585
R97 B.n720 B.n67 585
R98 B.n722 B.n721 585
R99 B.n724 B.n66 585
R100 B.n727 B.n726 585
R101 B.n728 B.n65 585
R102 B.n730 B.n729 585
R103 B.n732 B.n64 585
R104 B.n735 B.n734 585
R105 B.n736 B.n63 585
R106 B.n738 B.n737 585
R107 B.n740 B.n62 585
R108 B.n743 B.n742 585
R109 B.n744 B.n61 585
R110 B.n746 B.n745 585
R111 B.n748 B.n60 585
R112 B.n751 B.n750 585
R113 B.n752 B.n59 585
R114 B.n554 B.n57 585
R115 B.n755 B.n57 585
R116 B.n553 B.n56 585
R117 B.n756 B.n56 585
R118 B.n552 B.n55 585
R119 B.n757 B.n55 585
R120 B.n551 B.n550 585
R121 B.n550 B.n51 585
R122 B.n549 B.n50 585
R123 B.n763 B.n50 585
R124 B.n548 B.n49 585
R125 B.n764 B.n49 585
R126 B.n547 B.n48 585
R127 B.n765 B.n48 585
R128 B.n546 B.n545 585
R129 B.n545 B.n44 585
R130 B.n544 B.n43 585
R131 B.n771 B.n43 585
R132 B.n543 B.n42 585
R133 B.n772 B.n42 585
R134 B.n542 B.n41 585
R135 B.n773 B.n41 585
R136 B.n541 B.n540 585
R137 B.n540 B.n37 585
R138 B.n539 B.n36 585
R139 B.n779 B.n36 585
R140 B.n538 B.n35 585
R141 B.n780 B.n35 585
R142 B.n537 B.n34 585
R143 B.n781 B.n34 585
R144 B.n536 B.n535 585
R145 B.n535 B.n30 585
R146 B.n534 B.n29 585
R147 B.n787 B.n29 585
R148 B.n533 B.n28 585
R149 B.n788 B.n28 585
R150 B.n532 B.n27 585
R151 B.n789 B.n27 585
R152 B.n531 B.n530 585
R153 B.n530 B.n23 585
R154 B.n529 B.n22 585
R155 B.n795 B.n22 585
R156 B.n528 B.n21 585
R157 B.n796 B.n21 585
R158 B.n527 B.n20 585
R159 B.n797 B.n20 585
R160 B.n526 B.n525 585
R161 B.n525 B.n19 585
R162 B.n524 B.n15 585
R163 B.n803 B.n15 585
R164 B.n523 B.n14 585
R165 B.n804 B.n14 585
R166 B.n522 B.n13 585
R167 B.n805 B.n13 585
R168 B.n521 B.n520 585
R169 B.n520 B.n12 585
R170 B.n519 B.n518 585
R171 B.n519 B.n8 585
R172 B.n517 B.n7 585
R173 B.n812 B.n7 585
R174 B.n516 B.n6 585
R175 B.n813 B.n6 585
R176 B.n515 B.n5 585
R177 B.n814 B.n5 585
R178 B.n514 B.n513 585
R179 B.n513 B.n4 585
R180 B.n512 B.n114 585
R181 B.n512 B.n511 585
R182 B.n502 B.n115 585
R183 B.n116 B.n115 585
R184 B.n504 B.n503 585
R185 B.n505 B.n504 585
R186 B.n501 B.n121 585
R187 B.n121 B.n120 585
R188 B.n500 B.n499 585
R189 B.n499 B.n498 585
R190 B.n123 B.n122 585
R191 B.n491 B.n123 585
R192 B.n490 B.n489 585
R193 B.n492 B.n490 585
R194 B.n488 B.n128 585
R195 B.n128 B.n127 585
R196 B.n487 B.n486 585
R197 B.n486 B.n485 585
R198 B.n130 B.n129 585
R199 B.n131 B.n130 585
R200 B.n478 B.n477 585
R201 B.n479 B.n478 585
R202 B.n476 B.n136 585
R203 B.n136 B.n135 585
R204 B.n475 B.n474 585
R205 B.n474 B.n473 585
R206 B.n138 B.n137 585
R207 B.n139 B.n138 585
R208 B.n466 B.n465 585
R209 B.n467 B.n466 585
R210 B.n464 B.n144 585
R211 B.n144 B.n143 585
R212 B.n463 B.n462 585
R213 B.n462 B.n461 585
R214 B.n146 B.n145 585
R215 B.n147 B.n146 585
R216 B.n454 B.n453 585
R217 B.n455 B.n454 585
R218 B.n452 B.n152 585
R219 B.n152 B.n151 585
R220 B.n451 B.n450 585
R221 B.n450 B.n449 585
R222 B.n154 B.n153 585
R223 B.n155 B.n154 585
R224 B.n442 B.n441 585
R225 B.n443 B.n442 585
R226 B.n440 B.n160 585
R227 B.n160 B.n159 585
R228 B.n439 B.n438 585
R229 B.n438 B.n437 585
R230 B.n162 B.n161 585
R231 B.n163 B.n162 585
R232 B.n430 B.n429 585
R233 B.n431 B.n430 585
R234 B.n428 B.n168 585
R235 B.n168 B.n167 585
R236 B.n427 B.n426 585
R237 B.n426 B.n425 585
R238 B.n422 B.n172 585
R239 B.n421 B.n420 585
R240 B.n418 B.n173 585
R241 B.n418 B.n171 585
R242 B.n417 B.n416 585
R243 B.n415 B.n414 585
R244 B.n413 B.n175 585
R245 B.n411 B.n410 585
R246 B.n409 B.n176 585
R247 B.n408 B.n407 585
R248 B.n405 B.n177 585
R249 B.n403 B.n402 585
R250 B.n401 B.n178 585
R251 B.n400 B.n399 585
R252 B.n397 B.n179 585
R253 B.n395 B.n394 585
R254 B.n393 B.n180 585
R255 B.n392 B.n391 585
R256 B.n389 B.n181 585
R257 B.n387 B.n386 585
R258 B.n385 B.n182 585
R259 B.n384 B.n383 585
R260 B.n381 B.n183 585
R261 B.n379 B.n378 585
R262 B.n377 B.n184 585
R263 B.n376 B.n375 585
R264 B.n373 B.n185 585
R265 B.n371 B.n370 585
R266 B.n369 B.n186 585
R267 B.n368 B.n367 585
R268 B.n365 B.n187 585
R269 B.n363 B.n362 585
R270 B.n361 B.n188 585
R271 B.n360 B.n359 585
R272 B.n357 B.n189 585
R273 B.n355 B.n354 585
R274 B.n353 B.n190 585
R275 B.n352 B.n351 585
R276 B.n349 B.n191 585
R277 B.n347 B.n346 585
R278 B.n345 B.n192 585
R279 B.n344 B.n343 585
R280 B.n341 B.n193 585
R281 B.n339 B.n338 585
R282 B.n337 B.n194 585
R283 B.n336 B.n335 585
R284 B.n333 B.n332 585
R285 B.n331 B.n330 585
R286 B.n329 B.n199 585
R287 B.n327 B.n326 585
R288 B.n325 B.n200 585
R289 B.n324 B.n323 585
R290 B.n321 B.n201 585
R291 B.n319 B.n318 585
R292 B.n317 B.n202 585
R293 B.n315 B.n314 585
R294 B.n312 B.n205 585
R295 B.n310 B.n309 585
R296 B.n308 B.n206 585
R297 B.n307 B.n306 585
R298 B.n304 B.n207 585
R299 B.n302 B.n301 585
R300 B.n300 B.n208 585
R301 B.n299 B.n298 585
R302 B.n296 B.n209 585
R303 B.n294 B.n293 585
R304 B.n292 B.n210 585
R305 B.n291 B.n290 585
R306 B.n288 B.n211 585
R307 B.n286 B.n285 585
R308 B.n284 B.n212 585
R309 B.n283 B.n282 585
R310 B.n280 B.n213 585
R311 B.n278 B.n277 585
R312 B.n276 B.n214 585
R313 B.n275 B.n274 585
R314 B.n272 B.n215 585
R315 B.n270 B.n269 585
R316 B.n268 B.n216 585
R317 B.n267 B.n266 585
R318 B.n264 B.n217 585
R319 B.n262 B.n261 585
R320 B.n260 B.n218 585
R321 B.n259 B.n258 585
R322 B.n256 B.n219 585
R323 B.n254 B.n253 585
R324 B.n252 B.n220 585
R325 B.n251 B.n250 585
R326 B.n248 B.n221 585
R327 B.n246 B.n245 585
R328 B.n244 B.n222 585
R329 B.n243 B.n242 585
R330 B.n240 B.n223 585
R331 B.n238 B.n237 585
R332 B.n236 B.n224 585
R333 B.n235 B.n234 585
R334 B.n232 B.n225 585
R335 B.n230 B.n229 585
R336 B.n228 B.n227 585
R337 B.n170 B.n169 585
R338 B.n424 B.n423 585
R339 B.n425 B.n424 585
R340 B.n166 B.n165 585
R341 B.n167 B.n166 585
R342 B.n433 B.n432 585
R343 B.n432 B.n431 585
R344 B.n434 B.n164 585
R345 B.n164 B.n163 585
R346 B.n436 B.n435 585
R347 B.n437 B.n436 585
R348 B.n158 B.n157 585
R349 B.n159 B.n158 585
R350 B.n445 B.n444 585
R351 B.n444 B.n443 585
R352 B.n446 B.n156 585
R353 B.n156 B.n155 585
R354 B.n448 B.n447 585
R355 B.n449 B.n448 585
R356 B.n150 B.n149 585
R357 B.n151 B.n150 585
R358 B.n457 B.n456 585
R359 B.n456 B.n455 585
R360 B.n458 B.n148 585
R361 B.n148 B.n147 585
R362 B.n460 B.n459 585
R363 B.n461 B.n460 585
R364 B.n142 B.n141 585
R365 B.n143 B.n142 585
R366 B.n469 B.n468 585
R367 B.n468 B.n467 585
R368 B.n470 B.n140 585
R369 B.n140 B.n139 585
R370 B.n472 B.n471 585
R371 B.n473 B.n472 585
R372 B.n134 B.n133 585
R373 B.n135 B.n134 585
R374 B.n481 B.n480 585
R375 B.n480 B.n479 585
R376 B.n482 B.n132 585
R377 B.n132 B.n131 585
R378 B.n484 B.n483 585
R379 B.n485 B.n484 585
R380 B.n126 B.n125 585
R381 B.n127 B.n126 585
R382 B.n494 B.n493 585
R383 B.n493 B.n492 585
R384 B.n495 B.n124 585
R385 B.n491 B.n124 585
R386 B.n497 B.n496 585
R387 B.n498 B.n497 585
R388 B.n119 B.n118 585
R389 B.n120 B.n119 585
R390 B.n507 B.n506 585
R391 B.n506 B.n505 585
R392 B.n508 B.n117 585
R393 B.n117 B.n116 585
R394 B.n510 B.n509 585
R395 B.n511 B.n510 585
R396 B.n3 B.n0 585
R397 B.n4 B.n3 585
R398 B.n811 B.n1 585
R399 B.n812 B.n811 585
R400 B.n810 B.n809 585
R401 B.n810 B.n8 585
R402 B.n808 B.n9 585
R403 B.n12 B.n9 585
R404 B.n807 B.n806 585
R405 B.n806 B.n805 585
R406 B.n11 B.n10 585
R407 B.n804 B.n11 585
R408 B.n802 B.n801 585
R409 B.n803 B.n802 585
R410 B.n800 B.n16 585
R411 B.n19 B.n16 585
R412 B.n799 B.n798 585
R413 B.n798 B.n797 585
R414 B.n18 B.n17 585
R415 B.n796 B.n18 585
R416 B.n794 B.n793 585
R417 B.n795 B.n794 585
R418 B.n792 B.n24 585
R419 B.n24 B.n23 585
R420 B.n791 B.n790 585
R421 B.n790 B.n789 585
R422 B.n26 B.n25 585
R423 B.n788 B.n26 585
R424 B.n786 B.n785 585
R425 B.n787 B.n786 585
R426 B.n784 B.n31 585
R427 B.n31 B.n30 585
R428 B.n783 B.n782 585
R429 B.n782 B.n781 585
R430 B.n33 B.n32 585
R431 B.n780 B.n33 585
R432 B.n778 B.n777 585
R433 B.n779 B.n778 585
R434 B.n776 B.n38 585
R435 B.n38 B.n37 585
R436 B.n775 B.n774 585
R437 B.n774 B.n773 585
R438 B.n40 B.n39 585
R439 B.n772 B.n40 585
R440 B.n770 B.n769 585
R441 B.n771 B.n770 585
R442 B.n768 B.n45 585
R443 B.n45 B.n44 585
R444 B.n767 B.n766 585
R445 B.n766 B.n765 585
R446 B.n47 B.n46 585
R447 B.n764 B.n47 585
R448 B.n762 B.n761 585
R449 B.n763 B.n762 585
R450 B.n760 B.n52 585
R451 B.n52 B.n51 585
R452 B.n759 B.n758 585
R453 B.n758 B.n757 585
R454 B.n54 B.n53 585
R455 B.n756 B.n54 585
R456 B.n754 B.n753 585
R457 B.n755 B.n754 585
R458 B.n815 B.n814 585
R459 B.n813 B.n2 585
R460 B.n754 B.n59 545.355
R461 B.n113 B.n57 545.355
R462 B.n426 B.n170 545.355
R463 B.n424 B.n172 545.355
R464 B.n82 B.t9 299.296
R465 B.n88 B.t13 299.296
R466 B.n203 B.t6 299.296
R467 B.n195 B.t2 299.296
R468 B.n558 B.n58 256.663
R469 B.n560 B.n58 256.663
R470 B.n566 B.n58 256.663
R471 B.n568 B.n58 256.663
R472 B.n574 B.n58 256.663
R473 B.n576 B.n58 256.663
R474 B.n582 B.n58 256.663
R475 B.n584 B.n58 256.663
R476 B.n590 B.n58 256.663
R477 B.n592 B.n58 256.663
R478 B.n598 B.n58 256.663
R479 B.n600 B.n58 256.663
R480 B.n606 B.n58 256.663
R481 B.n608 B.n58 256.663
R482 B.n614 B.n58 256.663
R483 B.n616 B.n58 256.663
R484 B.n622 B.n58 256.663
R485 B.n624 B.n58 256.663
R486 B.n630 B.n58 256.663
R487 B.n632 B.n58 256.663
R488 B.n638 B.n58 256.663
R489 B.n91 B.n58 256.663
R490 B.n644 B.n58 256.663
R491 B.n650 B.n58 256.663
R492 B.n652 B.n58 256.663
R493 B.n658 B.n58 256.663
R494 B.n660 B.n58 256.663
R495 B.n667 B.n58 256.663
R496 B.n669 B.n58 256.663
R497 B.n675 B.n58 256.663
R498 B.n677 B.n58 256.663
R499 B.n683 B.n58 256.663
R500 B.n685 B.n58 256.663
R501 B.n691 B.n58 256.663
R502 B.n693 B.n58 256.663
R503 B.n699 B.n58 256.663
R504 B.n701 B.n58 256.663
R505 B.n707 B.n58 256.663
R506 B.n709 B.n58 256.663
R507 B.n715 B.n58 256.663
R508 B.n717 B.n58 256.663
R509 B.n723 B.n58 256.663
R510 B.n725 B.n58 256.663
R511 B.n731 B.n58 256.663
R512 B.n733 B.n58 256.663
R513 B.n739 B.n58 256.663
R514 B.n741 B.n58 256.663
R515 B.n747 B.n58 256.663
R516 B.n749 B.n58 256.663
R517 B.n419 B.n171 256.663
R518 B.n174 B.n171 256.663
R519 B.n412 B.n171 256.663
R520 B.n406 B.n171 256.663
R521 B.n404 B.n171 256.663
R522 B.n398 B.n171 256.663
R523 B.n396 B.n171 256.663
R524 B.n390 B.n171 256.663
R525 B.n388 B.n171 256.663
R526 B.n382 B.n171 256.663
R527 B.n380 B.n171 256.663
R528 B.n374 B.n171 256.663
R529 B.n372 B.n171 256.663
R530 B.n366 B.n171 256.663
R531 B.n364 B.n171 256.663
R532 B.n358 B.n171 256.663
R533 B.n356 B.n171 256.663
R534 B.n350 B.n171 256.663
R535 B.n348 B.n171 256.663
R536 B.n342 B.n171 256.663
R537 B.n340 B.n171 256.663
R538 B.n334 B.n171 256.663
R539 B.n198 B.n171 256.663
R540 B.n328 B.n171 256.663
R541 B.n322 B.n171 256.663
R542 B.n320 B.n171 256.663
R543 B.n313 B.n171 256.663
R544 B.n311 B.n171 256.663
R545 B.n305 B.n171 256.663
R546 B.n303 B.n171 256.663
R547 B.n297 B.n171 256.663
R548 B.n295 B.n171 256.663
R549 B.n289 B.n171 256.663
R550 B.n287 B.n171 256.663
R551 B.n281 B.n171 256.663
R552 B.n279 B.n171 256.663
R553 B.n273 B.n171 256.663
R554 B.n271 B.n171 256.663
R555 B.n265 B.n171 256.663
R556 B.n263 B.n171 256.663
R557 B.n257 B.n171 256.663
R558 B.n255 B.n171 256.663
R559 B.n249 B.n171 256.663
R560 B.n247 B.n171 256.663
R561 B.n241 B.n171 256.663
R562 B.n239 B.n171 256.663
R563 B.n233 B.n171 256.663
R564 B.n231 B.n171 256.663
R565 B.n226 B.n171 256.663
R566 B.n817 B.n816 256.663
R567 B.n750 B.n748 163.367
R568 B.n746 B.n61 163.367
R569 B.n742 B.n740 163.367
R570 B.n738 B.n63 163.367
R571 B.n734 B.n732 163.367
R572 B.n730 B.n65 163.367
R573 B.n726 B.n724 163.367
R574 B.n722 B.n67 163.367
R575 B.n718 B.n716 163.367
R576 B.n714 B.n69 163.367
R577 B.n710 B.n708 163.367
R578 B.n706 B.n71 163.367
R579 B.n702 B.n700 163.367
R580 B.n698 B.n73 163.367
R581 B.n694 B.n692 163.367
R582 B.n690 B.n75 163.367
R583 B.n686 B.n684 163.367
R584 B.n682 B.n77 163.367
R585 B.n678 B.n676 163.367
R586 B.n674 B.n79 163.367
R587 B.n670 B.n668 163.367
R588 B.n666 B.n81 163.367
R589 B.n661 B.n659 163.367
R590 B.n657 B.n85 163.367
R591 B.n653 B.n651 163.367
R592 B.n649 B.n87 163.367
R593 B.n645 B.n643 163.367
R594 B.n640 B.n639 163.367
R595 B.n637 B.n93 163.367
R596 B.n633 B.n631 163.367
R597 B.n629 B.n95 163.367
R598 B.n625 B.n623 163.367
R599 B.n621 B.n97 163.367
R600 B.n617 B.n615 163.367
R601 B.n613 B.n99 163.367
R602 B.n609 B.n607 163.367
R603 B.n605 B.n101 163.367
R604 B.n601 B.n599 163.367
R605 B.n597 B.n103 163.367
R606 B.n593 B.n591 163.367
R607 B.n589 B.n105 163.367
R608 B.n585 B.n583 163.367
R609 B.n581 B.n107 163.367
R610 B.n577 B.n575 163.367
R611 B.n573 B.n109 163.367
R612 B.n569 B.n567 163.367
R613 B.n565 B.n111 163.367
R614 B.n561 B.n559 163.367
R615 B.n557 B.n113 163.367
R616 B.n426 B.n168 163.367
R617 B.n430 B.n168 163.367
R618 B.n430 B.n162 163.367
R619 B.n438 B.n162 163.367
R620 B.n438 B.n160 163.367
R621 B.n442 B.n160 163.367
R622 B.n442 B.n154 163.367
R623 B.n450 B.n154 163.367
R624 B.n450 B.n152 163.367
R625 B.n454 B.n152 163.367
R626 B.n454 B.n146 163.367
R627 B.n462 B.n146 163.367
R628 B.n462 B.n144 163.367
R629 B.n466 B.n144 163.367
R630 B.n466 B.n138 163.367
R631 B.n474 B.n138 163.367
R632 B.n474 B.n136 163.367
R633 B.n478 B.n136 163.367
R634 B.n478 B.n130 163.367
R635 B.n486 B.n130 163.367
R636 B.n486 B.n128 163.367
R637 B.n490 B.n128 163.367
R638 B.n490 B.n123 163.367
R639 B.n499 B.n123 163.367
R640 B.n499 B.n121 163.367
R641 B.n504 B.n121 163.367
R642 B.n504 B.n115 163.367
R643 B.n512 B.n115 163.367
R644 B.n513 B.n512 163.367
R645 B.n513 B.n5 163.367
R646 B.n6 B.n5 163.367
R647 B.n7 B.n6 163.367
R648 B.n519 B.n7 163.367
R649 B.n520 B.n519 163.367
R650 B.n520 B.n13 163.367
R651 B.n14 B.n13 163.367
R652 B.n15 B.n14 163.367
R653 B.n525 B.n15 163.367
R654 B.n525 B.n20 163.367
R655 B.n21 B.n20 163.367
R656 B.n22 B.n21 163.367
R657 B.n530 B.n22 163.367
R658 B.n530 B.n27 163.367
R659 B.n28 B.n27 163.367
R660 B.n29 B.n28 163.367
R661 B.n535 B.n29 163.367
R662 B.n535 B.n34 163.367
R663 B.n35 B.n34 163.367
R664 B.n36 B.n35 163.367
R665 B.n540 B.n36 163.367
R666 B.n540 B.n41 163.367
R667 B.n42 B.n41 163.367
R668 B.n43 B.n42 163.367
R669 B.n545 B.n43 163.367
R670 B.n545 B.n48 163.367
R671 B.n49 B.n48 163.367
R672 B.n50 B.n49 163.367
R673 B.n550 B.n50 163.367
R674 B.n550 B.n55 163.367
R675 B.n56 B.n55 163.367
R676 B.n57 B.n56 163.367
R677 B.n420 B.n418 163.367
R678 B.n418 B.n417 163.367
R679 B.n414 B.n413 163.367
R680 B.n411 B.n176 163.367
R681 B.n407 B.n405 163.367
R682 B.n403 B.n178 163.367
R683 B.n399 B.n397 163.367
R684 B.n395 B.n180 163.367
R685 B.n391 B.n389 163.367
R686 B.n387 B.n182 163.367
R687 B.n383 B.n381 163.367
R688 B.n379 B.n184 163.367
R689 B.n375 B.n373 163.367
R690 B.n371 B.n186 163.367
R691 B.n367 B.n365 163.367
R692 B.n363 B.n188 163.367
R693 B.n359 B.n357 163.367
R694 B.n355 B.n190 163.367
R695 B.n351 B.n349 163.367
R696 B.n347 B.n192 163.367
R697 B.n343 B.n341 163.367
R698 B.n339 B.n194 163.367
R699 B.n335 B.n333 163.367
R700 B.n330 B.n329 163.367
R701 B.n327 B.n200 163.367
R702 B.n323 B.n321 163.367
R703 B.n319 B.n202 163.367
R704 B.n314 B.n312 163.367
R705 B.n310 B.n206 163.367
R706 B.n306 B.n304 163.367
R707 B.n302 B.n208 163.367
R708 B.n298 B.n296 163.367
R709 B.n294 B.n210 163.367
R710 B.n290 B.n288 163.367
R711 B.n286 B.n212 163.367
R712 B.n282 B.n280 163.367
R713 B.n278 B.n214 163.367
R714 B.n274 B.n272 163.367
R715 B.n270 B.n216 163.367
R716 B.n266 B.n264 163.367
R717 B.n262 B.n218 163.367
R718 B.n258 B.n256 163.367
R719 B.n254 B.n220 163.367
R720 B.n250 B.n248 163.367
R721 B.n246 B.n222 163.367
R722 B.n242 B.n240 163.367
R723 B.n238 B.n224 163.367
R724 B.n234 B.n232 163.367
R725 B.n230 B.n227 163.367
R726 B.n424 B.n166 163.367
R727 B.n432 B.n166 163.367
R728 B.n432 B.n164 163.367
R729 B.n436 B.n164 163.367
R730 B.n436 B.n158 163.367
R731 B.n444 B.n158 163.367
R732 B.n444 B.n156 163.367
R733 B.n448 B.n156 163.367
R734 B.n448 B.n150 163.367
R735 B.n456 B.n150 163.367
R736 B.n456 B.n148 163.367
R737 B.n460 B.n148 163.367
R738 B.n460 B.n142 163.367
R739 B.n468 B.n142 163.367
R740 B.n468 B.n140 163.367
R741 B.n472 B.n140 163.367
R742 B.n472 B.n134 163.367
R743 B.n480 B.n134 163.367
R744 B.n480 B.n132 163.367
R745 B.n484 B.n132 163.367
R746 B.n484 B.n126 163.367
R747 B.n493 B.n126 163.367
R748 B.n493 B.n124 163.367
R749 B.n497 B.n124 163.367
R750 B.n497 B.n119 163.367
R751 B.n506 B.n119 163.367
R752 B.n506 B.n117 163.367
R753 B.n510 B.n117 163.367
R754 B.n510 B.n3 163.367
R755 B.n815 B.n3 163.367
R756 B.n811 B.n2 163.367
R757 B.n811 B.n810 163.367
R758 B.n810 B.n9 163.367
R759 B.n806 B.n9 163.367
R760 B.n806 B.n11 163.367
R761 B.n802 B.n11 163.367
R762 B.n802 B.n16 163.367
R763 B.n798 B.n16 163.367
R764 B.n798 B.n18 163.367
R765 B.n794 B.n18 163.367
R766 B.n794 B.n24 163.367
R767 B.n790 B.n24 163.367
R768 B.n790 B.n26 163.367
R769 B.n786 B.n26 163.367
R770 B.n786 B.n31 163.367
R771 B.n782 B.n31 163.367
R772 B.n782 B.n33 163.367
R773 B.n778 B.n33 163.367
R774 B.n778 B.n38 163.367
R775 B.n774 B.n38 163.367
R776 B.n774 B.n40 163.367
R777 B.n770 B.n40 163.367
R778 B.n770 B.n45 163.367
R779 B.n766 B.n45 163.367
R780 B.n766 B.n47 163.367
R781 B.n762 B.n47 163.367
R782 B.n762 B.n52 163.367
R783 B.n758 B.n52 163.367
R784 B.n758 B.n54 163.367
R785 B.n754 B.n54 163.367
R786 B.n88 B.t14 145.423
R787 B.n203 B.t8 145.423
R788 B.n82 B.t11 145.405
R789 B.n195 B.t5 145.405
R790 B.n425 B.n171 79.6195
R791 B.n755 B.n58 79.6195
R792 B.n83 B.n82 74.2793
R793 B.n89 B.n88 74.2793
R794 B.n204 B.n203 74.2793
R795 B.n196 B.n195 74.2793
R796 B.n749 B.n59 71.676
R797 B.n748 B.n747 71.676
R798 B.n741 B.n61 71.676
R799 B.n740 B.n739 71.676
R800 B.n733 B.n63 71.676
R801 B.n732 B.n731 71.676
R802 B.n725 B.n65 71.676
R803 B.n724 B.n723 71.676
R804 B.n717 B.n67 71.676
R805 B.n716 B.n715 71.676
R806 B.n709 B.n69 71.676
R807 B.n708 B.n707 71.676
R808 B.n701 B.n71 71.676
R809 B.n700 B.n699 71.676
R810 B.n693 B.n73 71.676
R811 B.n692 B.n691 71.676
R812 B.n685 B.n75 71.676
R813 B.n684 B.n683 71.676
R814 B.n677 B.n77 71.676
R815 B.n676 B.n675 71.676
R816 B.n669 B.n79 71.676
R817 B.n668 B.n667 71.676
R818 B.n660 B.n81 71.676
R819 B.n659 B.n658 71.676
R820 B.n652 B.n85 71.676
R821 B.n651 B.n650 71.676
R822 B.n644 B.n87 71.676
R823 B.n643 B.n91 71.676
R824 B.n639 B.n638 71.676
R825 B.n632 B.n93 71.676
R826 B.n631 B.n630 71.676
R827 B.n624 B.n95 71.676
R828 B.n623 B.n622 71.676
R829 B.n616 B.n97 71.676
R830 B.n615 B.n614 71.676
R831 B.n608 B.n99 71.676
R832 B.n607 B.n606 71.676
R833 B.n600 B.n101 71.676
R834 B.n599 B.n598 71.676
R835 B.n592 B.n103 71.676
R836 B.n591 B.n590 71.676
R837 B.n584 B.n105 71.676
R838 B.n583 B.n582 71.676
R839 B.n576 B.n107 71.676
R840 B.n575 B.n574 71.676
R841 B.n568 B.n109 71.676
R842 B.n567 B.n566 71.676
R843 B.n560 B.n111 71.676
R844 B.n559 B.n558 71.676
R845 B.n558 B.n557 71.676
R846 B.n561 B.n560 71.676
R847 B.n566 B.n565 71.676
R848 B.n569 B.n568 71.676
R849 B.n574 B.n573 71.676
R850 B.n577 B.n576 71.676
R851 B.n582 B.n581 71.676
R852 B.n585 B.n584 71.676
R853 B.n590 B.n589 71.676
R854 B.n593 B.n592 71.676
R855 B.n598 B.n597 71.676
R856 B.n601 B.n600 71.676
R857 B.n606 B.n605 71.676
R858 B.n609 B.n608 71.676
R859 B.n614 B.n613 71.676
R860 B.n617 B.n616 71.676
R861 B.n622 B.n621 71.676
R862 B.n625 B.n624 71.676
R863 B.n630 B.n629 71.676
R864 B.n633 B.n632 71.676
R865 B.n638 B.n637 71.676
R866 B.n640 B.n91 71.676
R867 B.n645 B.n644 71.676
R868 B.n650 B.n649 71.676
R869 B.n653 B.n652 71.676
R870 B.n658 B.n657 71.676
R871 B.n661 B.n660 71.676
R872 B.n667 B.n666 71.676
R873 B.n670 B.n669 71.676
R874 B.n675 B.n674 71.676
R875 B.n678 B.n677 71.676
R876 B.n683 B.n682 71.676
R877 B.n686 B.n685 71.676
R878 B.n691 B.n690 71.676
R879 B.n694 B.n693 71.676
R880 B.n699 B.n698 71.676
R881 B.n702 B.n701 71.676
R882 B.n707 B.n706 71.676
R883 B.n710 B.n709 71.676
R884 B.n715 B.n714 71.676
R885 B.n718 B.n717 71.676
R886 B.n723 B.n722 71.676
R887 B.n726 B.n725 71.676
R888 B.n731 B.n730 71.676
R889 B.n734 B.n733 71.676
R890 B.n739 B.n738 71.676
R891 B.n742 B.n741 71.676
R892 B.n747 B.n746 71.676
R893 B.n750 B.n749 71.676
R894 B.n419 B.n172 71.676
R895 B.n417 B.n174 71.676
R896 B.n413 B.n412 71.676
R897 B.n406 B.n176 71.676
R898 B.n405 B.n404 71.676
R899 B.n398 B.n178 71.676
R900 B.n397 B.n396 71.676
R901 B.n390 B.n180 71.676
R902 B.n389 B.n388 71.676
R903 B.n382 B.n182 71.676
R904 B.n381 B.n380 71.676
R905 B.n374 B.n184 71.676
R906 B.n373 B.n372 71.676
R907 B.n366 B.n186 71.676
R908 B.n365 B.n364 71.676
R909 B.n358 B.n188 71.676
R910 B.n357 B.n356 71.676
R911 B.n350 B.n190 71.676
R912 B.n349 B.n348 71.676
R913 B.n342 B.n192 71.676
R914 B.n341 B.n340 71.676
R915 B.n334 B.n194 71.676
R916 B.n333 B.n198 71.676
R917 B.n329 B.n328 71.676
R918 B.n322 B.n200 71.676
R919 B.n321 B.n320 71.676
R920 B.n313 B.n202 71.676
R921 B.n312 B.n311 71.676
R922 B.n305 B.n206 71.676
R923 B.n304 B.n303 71.676
R924 B.n297 B.n208 71.676
R925 B.n296 B.n295 71.676
R926 B.n289 B.n210 71.676
R927 B.n288 B.n287 71.676
R928 B.n281 B.n212 71.676
R929 B.n280 B.n279 71.676
R930 B.n273 B.n214 71.676
R931 B.n272 B.n271 71.676
R932 B.n265 B.n216 71.676
R933 B.n264 B.n263 71.676
R934 B.n257 B.n218 71.676
R935 B.n256 B.n255 71.676
R936 B.n249 B.n220 71.676
R937 B.n248 B.n247 71.676
R938 B.n241 B.n222 71.676
R939 B.n240 B.n239 71.676
R940 B.n233 B.n224 71.676
R941 B.n232 B.n231 71.676
R942 B.n227 B.n226 71.676
R943 B.n420 B.n419 71.676
R944 B.n414 B.n174 71.676
R945 B.n412 B.n411 71.676
R946 B.n407 B.n406 71.676
R947 B.n404 B.n403 71.676
R948 B.n399 B.n398 71.676
R949 B.n396 B.n395 71.676
R950 B.n391 B.n390 71.676
R951 B.n388 B.n387 71.676
R952 B.n383 B.n382 71.676
R953 B.n380 B.n379 71.676
R954 B.n375 B.n374 71.676
R955 B.n372 B.n371 71.676
R956 B.n367 B.n366 71.676
R957 B.n364 B.n363 71.676
R958 B.n359 B.n358 71.676
R959 B.n356 B.n355 71.676
R960 B.n351 B.n350 71.676
R961 B.n348 B.n347 71.676
R962 B.n343 B.n342 71.676
R963 B.n340 B.n339 71.676
R964 B.n335 B.n334 71.676
R965 B.n330 B.n198 71.676
R966 B.n328 B.n327 71.676
R967 B.n323 B.n322 71.676
R968 B.n320 B.n319 71.676
R969 B.n314 B.n313 71.676
R970 B.n311 B.n310 71.676
R971 B.n306 B.n305 71.676
R972 B.n303 B.n302 71.676
R973 B.n298 B.n297 71.676
R974 B.n295 B.n294 71.676
R975 B.n290 B.n289 71.676
R976 B.n287 B.n286 71.676
R977 B.n282 B.n281 71.676
R978 B.n279 B.n278 71.676
R979 B.n274 B.n273 71.676
R980 B.n271 B.n270 71.676
R981 B.n266 B.n265 71.676
R982 B.n263 B.n262 71.676
R983 B.n258 B.n257 71.676
R984 B.n255 B.n254 71.676
R985 B.n250 B.n249 71.676
R986 B.n247 B.n246 71.676
R987 B.n242 B.n241 71.676
R988 B.n239 B.n238 71.676
R989 B.n234 B.n233 71.676
R990 B.n231 B.n230 71.676
R991 B.n226 B.n170 71.676
R992 B.n816 B.n815 71.676
R993 B.n816 B.n2 71.676
R994 B.n89 B.t15 71.1437
R995 B.n204 B.t7 71.1437
R996 B.n83 B.t12 71.127
R997 B.n196 B.t4 71.127
R998 B.n663 B.n83 59.5399
R999 B.n90 B.n89 59.5399
R1000 B.n316 B.n204 59.5399
R1001 B.n197 B.n196 59.5399
R1002 B.n425 B.n167 40.708
R1003 B.n431 B.n167 40.708
R1004 B.n431 B.n163 40.708
R1005 B.n437 B.n163 40.708
R1006 B.n437 B.n159 40.708
R1007 B.n443 B.n159 40.708
R1008 B.n443 B.n155 40.708
R1009 B.n449 B.n155 40.708
R1010 B.n455 B.n151 40.708
R1011 B.n455 B.n147 40.708
R1012 B.n461 B.n147 40.708
R1013 B.n461 B.n143 40.708
R1014 B.n467 B.n143 40.708
R1015 B.n467 B.n139 40.708
R1016 B.n473 B.n139 40.708
R1017 B.n473 B.n135 40.708
R1018 B.n479 B.n135 40.708
R1019 B.n479 B.n131 40.708
R1020 B.n485 B.n131 40.708
R1021 B.n485 B.n127 40.708
R1022 B.n492 B.n127 40.708
R1023 B.n492 B.n491 40.708
R1024 B.n498 B.n120 40.708
R1025 B.n505 B.n120 40.708
R1026 B.n505 B.n116 40.708
R1027 B.n511 B.n116 40.708
R1028 B.n511 B.n4 40.708
R1029 B.n814 B.n4 40.708
R1030 B.n814 B.n813 40.708
R1031 B.n813 B.n812 40.708
R1032 B.n812 B.n8 40.708
R1033 B.n12 B.n8 40.708
R1034 B.n805 B.n12 40.708
R1035 B.n805 B.n804 40.708
R1036 B.n804 B.n803 40.708
R1037 B.n797 B.n19 40.708
R1038 B.n797 B.n796 40.708
R1039 B.n796 B.n795 40.708
R1040 B.n795 B.n23 40.708
R1041 B.n789 B.n23 40.708
R1042 B.n789 B.n788 40.708
R1043 B.n788 B.n787 40.708
R1044 B.n787 B.n30 40.708
R1045 B.n781 B.n30 40.708
R1046 B.n781 B.n780 40.708
R1047 B.n780 B.n779 40.708
R1048 B.n779 B.n37 40.708
R1049 B.n773 B.n37 40.708
R1050 B.n773 B.n772 40.708
R1051 B.n771 B.n44 40.708
R1052 B.n765 B.n44 40.708
R1053 B.n765 B.n764 40.708
R1054 B.n764 B.n763 40.708
R1055 B.n763 B.n51 40.708
R1056 B.n757 B.n51 40.708
R1057 B.n757 B.n756 40.708
R1058 B.n756 B.n755 40.708
R1059 B.n423 B.n422 35.4346
R1060 B.n427 B.n169 35.4346
R1061 B.n753 B.n752 35.4346
R1062 B.n555 B.n554 35.4346
R1063 B.n449 B.t3 32.327
R1064 B.t10 B.n771 32.327
R1065 B.n498 B.t0 29.9325
R1066 B.n803 B.t1 29.9325
R1067 B B.n817 18.0485
R1068 B.n491 B.t0 10.776
R1069 B.n19 B.t1 10.776
R1070 B.n423 B.n165 10.6151
R1071 B.n433 B.n165 10.6151
R1072 B.n434 B.n433 10.6151
R1073 B.n435 B.n434 10.6151
R1074 B.n435 B.n157 10.6151
R1075 B.n445 B.n157 10.6151
R1076 B.n446 B.n445 10.6151
R1077 B.n447 B.n446 10.6151
R1078 B.n447 B.n149 10.6151
R1079 B.n457 B.n149 10.6151
R1080 B.n458 B.n457 10.6151
R1081 B.n459 B.n458 10.6151
R1082 B.n459 B.n141 10.6151
R1083 B.n469 B.n141 10.6151
R1084 B.n470 B.n469 10.6151
R1085 B.n471 B.n470 10.6151
R1086 B.n471 B.n133 10.6151
R1087 B.n481 B.n133 10.6151
R1088 B.n482 B.n481 10.6151
R1089 B.n483 B.n482 10.6151
R1090 B.n483 B.n125 10.6151
R1091 B.n494 B.n125 10.6151
R1092 B.n495 B.n494 10.6151
R1093 B.n496 B.n495 10.6151
R1094 B.n496 B.n118 10.6151
R1095 B.n507 B.n118 10.6151
R1096 B.n508 B.n507 10.6151
R1097 B.n509 B.n508 10.6151
R1098 B.n509 B.n0 10.6151
R1099 B.n422 B.n421 10.6151
R1100 B.n421 B.n173 10.6151
R1101 B.n416 B.n173 10.6151
R1102 B.n416 B.n415 10.6151
R1103 B.n415 B.n175 10.6151
R1104 B.n410 B.n175 10.6151
R1105 B.n410 B.n409 10.6151
R1106 B.n409 B.n408 10.6151
R1107 B.n408 B.n177 10.6151
R1108 B.n402 B.n177 10.6151
R1109 B.n402 B.n401 10.6151
R1110 B.n401 B.n400 10.6151
R1111 B.n400 B.n179 10.6151
R1112 B.n394 B.n179 10.6151
R1113 B.n394 B.n393 10.6151
R1114 B.n393 B.n392 10.6151
R1115 B.n392 B.n181 10.6151
R1116 B.n386 B.n181 10.6151
R1117 B.n386 B.n385 10.6151
R1118 B.n385 B.n384 10.6151
R1119 B.n384 B.n183 10.6151
R1120 B.n378 B.n183 10.6151
R1121 B.n378 B.n377 10.6151
R1122 B.n377 B.n376 10.6151
R1123 B.n376 B.n185 10.6151
R1124 B.n370 B.n185 10.6151
R1125 B.n370 B.n369 10.6151
R1126 B.n369 B.n368 10.6151
R1127 B.n368 B.n187 10.6151
R1128 B.n362 B.n187 10.6151
R1129 B.n362 B.n361 10.6151
R1130 B.n361 B.n360 10.6151
R1131 B.n360 B.n189 10.6151
R1132 B.n354 B.n189 10.6151
R1133 B.n354 B.n353 10.6151
R1134 B.n353 B.n352 10.6151
R1135 B.n352 B.n191 10.6151
R1136 B.n346 B.n191 10.6151
R1137 B.n346 B.n345 10.6151
R1138 B.n345 B.n344 10.6151
R1139 B.n344 B.n193 10.6151
R1140 B.n338 B.n193 10.6151
R1141 B.n338 B.n337 10.6151
R1142 B.n337 B.n336 10.6151
R1143 B.n332 B.n331 10.6151
R1144 B.n331 B.n199 10.6151
R1145 B.n326 B.n199 10.6151
R1146 B.n326 B.n325 10.6151
R1147 B.n325 B.n324 10.6151
R1148 B.n324 B.n201 10.6151
R1149 B.n318 B.n201 10.6151
R1150 B.n318 B.n317 10.6151
R1151 B.n315 B.n205 10.6151
R1152 B.n309 B.n205 10.6151
R1153 B.n309 B.n308 10.6151
R1154 B.n308 B.n307 10.6151
R1155 B.n307 B.n207 10.6151
R1156 B.n301 B.n207 10.6151
R1157 B.n301 B.n300 10.6151
R1158 B.n300 B.n299 10.6151
R1159 B.n299 B.n209 10.6151
R1160 B.n293 B.n209 10.6151
R1161 B.n293 B.n292 10.6151
R1162 B.n292 B.n291 10.6151
R1163 B.n291 B.n211 10.6151
R1164 B.n285 B.n211 10.6151
R1165 B.n285 B.n284 10.6151
R1166 B.n284 B.n283 10.6151
R1167 B.n283 B.n213 10.6151
R1168 B.n277 B.n213 10.6151
R1169 B.n277 B.n276 10.6151
R1170 B.n276 B.n275 10.6151
R1171 B.n275 B.n215 10.6151
R1172 B.n269 B.n215 10.6151
R1173 B.n269 B.n268 10.6151
R1174 B.n268 B.n267 10.6151
R1175 B.n267 B.n217 10.6151
R1176 B.n261 B.n217 10.6151
R1177 B.n261 B.n260 10.6151
R1178 B.n260 B.n259 10.6151
R1179 B.n259 B.n219 10.6151
R1180 B.n253 B.n219 10.6151
R1181 B.n253 B.n252 10.6151
R1182 B.n252 B.n251 10.6151
R1183 B.n251 B.n221 10.6151
R1184 B.n245 B.n221 10.6151
R1185 B.n245 B.n244 10.6151
R1186 B.n244 B.n243 10.6151
R1187 B.n243 B.n223 10.6151
R1188 B.n237 B.n223 10.6151
R1189 B.n237 B.n236 10.6151
R1190 B.n236 B.n235 10.6151
R1191 B.n235 B.n225 10.6151
R1192 B.n229 B.n225 10.6151
R1193 B.n229 B.n228 10.6151
R1194 B.n228 B.n169 10.6151
R1195 B.n428 B.n427 10.6151
R1196 B.n429 B.n428 10.6151
R1197 B.n429 B.n161 10.6151
R1198 B.n439 B.n161 10.6151
R1199 B.n440 B.n439 10.6151
R1200 B.n441 B.n440 10.6151
R1201 B.n441 B.n153 10.6151
R1202 B.n451 B.n153 10.6151
R1203 B.n452 B.n451 10.6151
R1204 B.n453 B.n452 10.6151
R1205 B.n453 B.n145 10.6151
R1206 B.n463 B.n145 10.6151
R1207 B.n464 B.n463 10.6151
R1208 B.n465 B.n464 10.6151
R1209 B.n465 B.n137 10.6151
R1210 B.n475 B.n137 10.6151
R1211 B.n476 B.n475 10.6151
R1212 B.n477 B.n476 10.6151
R1213 B.n477 B.n129 10.6151
R1214 B.n487 B.n129 10.6151
R1215 B.n488 B.n487 10.6151
R1216 B.n489 B.n488 10.6151
R1217 B.n489 B.n122 10.6151
R1218 B.n500 B.n122 10.6151
R1219 B.n501 B.n500 10.6151
R1220 B.n503 B.n501 10.6151
R1221 B.n503 B.n502 10.6151
R1222 B.n502 B.n114 10.6151
R1223 B.n514 B.n114 10.6151
R1224 B.n515 B.n514 10.6151
R1225 B.n516 B.n515 10.6151
R1226 B.n517 B.n516 10.6151
R1227 B.n518 B.n517 10.6151
R1228 B.n521 B.n518 10.6151
R1229 B.n522 B.n521 10.6151
R1230 B.n523 B.n522 10.6151
R1231 B.n524 B.n523 10.6151
R1232 B.n526 B.n524 10.6151
R1233 B.n527 B.n526 10.6151
R1234 B.n528 B.n527 10.6151
R1235 B.n529 B.n528 10.6151
R1236 B.n531 B.n529 10.6151
R1237 B.n532 B.n531 10.6151
R1238 B.n533 B.n532 10.6151
R1239 B.n534 B.n533 10.6151
R1240 B.n536 B.n534 10.6151
R1241 B.n537 B.n536 10.6151
R1242 B.n538 B.n537 10.6151
R1243 B.n539 B.n538 10.6151
R1244 B.n541 B.n539 10.6151
R1245 B.n542 B.n541 10.6151
R1246 B.n543 B.n542 10.6151
R1247 B.n544 B.n543 10.6151
R1248 B.n546 B.n544 10.6151
R1249 B.n547 B.n546 10.6151
R1250 B.n548 B.n547 10.6151
R1251 B.n549 B.n548 10.6151
R1252 B.n551 B.n549 10.6151
R1253 B.n552 B.n551 10.6151
R1254 B.n553 B.n552 10.6151
R1255 B.n554 B.n553 10.6151
R1256 B.n809 B.n1 10.6151
R1257 B.n809 B.n808 10.6151
R1258 B.n808 B.n807 10.6151
R1259 B.n807 B.n10 10.6151
R1260 B.n801 B.n10 10.6151
R1261 B.n801 B.n800 10.6151
R1262 B.n800 B.n799 10.6151
R1263 B.n799 B.n17 10.6151
R1264 B.n793 B.n17 10.6151
R1265 B.n793 B.n792 10.6151
R1266 B.n792 B.n791 10.6151
R1267 B.n791 B.n25 10.6151
R1268 B.n785 B.n25 10.6151
R1269 B.n785 B.n784 10.6151
R1270 B.n784 B.n783 10.6151
R1271 B.n783 B.n32 10.6151
R1272 B.n777 B.n32 10.6151
R1273 B.n777 B.n776 10.6151
R1274 B.n776 B.n775 10.6151
R1275 B.n775 B.n39 10.6151
R1276 B.n769 B.n39 10.6151
R1277 B.n769 B.n768 10.6151
R1278 B.n768 B.n767 10.6151
R1279 B.n767 B.n46 10.6151
R1280 B.n761 B.n46 10.6151
R1281 B.n761 B.n760 10.6151
R1282 B.n760 B.n759 10.6151
R1283 B.n759 B.n53 10.6151
R1284 B.n753 B.n53 10.6151
R1285 B.n752 B.n751 10.6151
R1286 B.n751 B.n60 10.6151
R1287 B.n745 B.n60 10.6151
R1288 B.n745 B.n744 10.6151
R1289 B.n744 B.n743 10.6151
R1290 B.n743 B.n62 10.6151
R1291 B.n737 B.n62 10.6151
R1292 B.n737 B.n736 10.6151
R1293 B.n736 B.n735 10.6151
R1294 B.n735 B.n64 10.6151
R1295 B.n729 B.n64 10.6151
R1296 B.n729 B.n728 10.6151
R1297 B.n728 B.n727 10.6151
R1298 B.n727 B.n66 10.6151
R1299 B.n721 B.n66 10.6151
R1300 B.n721 B.n720 10.6151
R1301 B.n720 B.n719 10.6151
R1302 B.n719 B.n68 10.6151
R1303 B.n713 B.n68 10.6151
R1304 B.n713 B.n712 10.6151
R1305 B.n712 B.n711 10.6151
R1306 B.n711 B.n70 10.6151
R1307 B.n705 B.n70 10.6151
R1308 B.n705 B.n704 10.6151
R1309 B.n704 B.n703 10.6151
R1310 B.n703 B.n72 10.6151
R1311 B.n697 B.n72 10.6151
R1312 B.n697 B.n696 10.6151
R1313 B.n696 B.n695 10.6151
R1314 B.n695 B.n74 10.6151
R1315 B.n689 B.n74 10.6151
R1316 B.n689 B.n688 10.6151
R1317 B.n688 B.n687 10.6151
R1318 B.n687 B.n76 10.6151
R1319 B.n681 B.n76 10.6151
R1320 B.n681 B.n680 10.6151
R1321 B.n680 B.n679 10.6151
R1322 B.n679 B.n78 10.6151
R1323 B.n673 B.n78 10.6151
R1324 B.n673 B.n672 10.6151
R1325 B.n672 B.n671 10.6151
R1326 B.n671 B.n80 10.6151
R1327 B.n665 B.n80 10.6151
R1328 B.n665 B.n664 10.6151
R1329 B.n662 B.n84 10.6151
R1330 B.n656 B.n84 10.6151
R1331 B.n656 B.n655 10.6151
R1332 B.n655 B.n654 10.6151
R1333 B.n654 B.n86 10.6151
R1334 B.n648 B.n86 10.6151
R1335 B.n648 B.n647 10.6151
R1336 B.n647 B.n646 10.6151
R1337 B.n642 B.n641 10.6151
R1338 B.n641 B.n92 10.6151
R1339 B.n636 B.n92 10.6151
R1340 B.n636 B.n635 10.6151
R1341 B.n635 B.n634 10.6151
R1342 B.n634 B.n94 10.6151
R1343 B.n628 B.n94 10.6151
R1344 B.n628 B.n627 10.6151
R1345 B.n627 B.n626 10.6151
R1346 B.n626 B.n96 10.6151
R1347 B.n620 B.n96 10.6151
R1348 B.n620 B.n619 10.6151
R1349 B.n619 B.n618 10.6151
R1350 B.n618 B.n98 10.6151
R1351 B.n612 B.n98 10.6151
R1352 B.n612 B.n611 10.6151
R1353 B.n611 B.n610 10.6151
R1354 B.n610 B.n100 10.6151
R1355 B.n604 B.n100 10.6151
R1356 B.n604 B.n603 10.6151
R1357 B.n603 B.n602 10.6151
R1358 B.n602 B.n102 10.6151
R1359 B.n596 B.n102 10.6151
R1360 B.n596 B.n595 10.6151
R1361 B.n595 B.n594 10.6151
R1362 B.n594 B.n104 10.6151
R1363 B.n588 B.n104 10.6151
R1364 B.n588 B.n587 10.6151
R1365 B.n587 B.n586 10.6151
R1366 B.n586 B.n106 10.6151
R1367 B.n580 B.n106 10.6151
R1368 B.n580 B.n579 10.6151
R1369 B.n579 B.n578 10.6151
R1370 B.n578 B.n108 10.6151
R1371 B.n572 B.n108 10.6151
R1372 B.n572 B.n571 10.6151
R1373 B.n571 B.n570 10.6151
R1374 B.n570 B.n110 10.6151
R1375 B.n564 B.n110 10.6151
R1376 B.n564 B.n563 10.6151
R1377 B.n563 B.n562 10.6151
R1378 B.n562 B.n112 10.6151
R1379 B.n556 B.n112 10.6151
R1380 B.n556 B.n555 10.6151
R1381 B.t3 B.n151 8.38145
R1382 B.n772 B.t10 8.38145
R1383 B.n817 B.n0 8.11757
R1384 B.n817 B.n1 8.11757
R1385 B.n332 B.n197 6.5566
R1386 B.n317 B.n316 6.5566
R1387 B.n663 B.n662 6.5566
R1388 B.n646 B.n90 6.5566
R1389 B.n336 B.n197 4.05904
R1390 B.n316 B.n315 4.05904
R1391 B.n664 B.n663 4.05904
R1392 B.n642 B.n90 4.05904
R1393 VP.n0 VP.t0 176.925
R1394 VP.n0 VP.t1 129.049
R1395 VP VP.n0 0.526373
R1396 VDD1 VDD1.t0 104.103
R1397 VDD1 VDD1.t1 62.0808
C0 VN VP 6.07698f
C1 VTAIL VP 2.82161f
C2 VDD1 VDD2 0.784661f
C3 VDD1 VN 0.14887f
C4 VDD1 VTAIL 5.51738f
C5 VDD2 VN 3.13541f
C6 VDD1 VP 3.3555f
C7 VDD2 VTAIL 5.57461f
C8 VTAIL VN 2.80737f
C9 VDD2 VP 0.371285f
C10 VDD2 B 4.940294f
C11 VDD1 B 8.343359f
C12 VTAIL B 8.24308f
C13 VN B 11.83073f
C14 VP B 7.586739f
C15 VDD1.t1 B 2.43659f
C16 VDD1.t0 B 3.12247f
C17 VP.t0 B 4.33693f
C18 VP.t1 B 3.66791f
C19 VP.n0 B 4.19791f
C20 VDD2.t1 B 3.03441f
C21 VDD2.t0 B 2.3982f
C22 VDD2.n0 B 3.10101f
C23 VTAIL.t0 B 2.37164f
C24 VTAIL.n0 B 1.86259f
C25 VTAIL.t2 B 2.37165f
C26 VTAIL.n1 B 1.91402f
C27 VTAIL.t3 B 2.37164f
C28 VTAIL.n2 B 1.69269f
C29 VTAIL.t1 B 2.37164f
C30 VTAIL.n3 B 1.60196f
C31 VN.t0 B 3.57226f
C32 VN.t1 B 4.21848f
.ends

