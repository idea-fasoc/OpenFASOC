* NGSPICE file created from diff_pair_sample_0930.ext - technology: sky130A

.subckt diff_pair_sample_0930 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VP.t0 VDD1.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=0.6336 pd=4.17 as=0.6336 ps=4.17 w=3.84 l=1.02
X1 VDD1.t4 VP.t1 VTAIL.t17 B.t2 sky130_fd_pr__nfet_01v8 ad=0.6336 pd=4.17 as=0.6336 ps=4.17 w=3.84 l=1.02
X2 VDD2.t9 VN.t0 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.6336 pd=4.17 as=0.6336 ps=4.17 w=3.84 l=1.02
X3 B.t22 B.t20 B.t21 B.t10 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=8.46 as=0 ps=0 w=3.84 l=1.02
X4 VDD1.t6 VP.t2 VTAIL.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=8.46 as=0.6336 ps=4.17 w=3.84 l=1.02
X5 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=8.46 as=0 ps=0 w=3.84 l=1.02
X6 VDD2.t8 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.6336 pd=4.17 as=1.4976 ps=8.46 w=3.84 l=1.02
X7 VTAIL.t19 VN.t2 VDD2.t7 B.t23 sky130_fd_pr__nfet_01v8 ad=0.6336 pd=4.17 as=0.6336 ps=4.17 w=3.84 l=1.02
X8 VTAIL.t15 VP.t3 VDD1.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=0.6336 pd=4.17 as=0.6336 ps=4.17 w=3.84 l=1.02
X9 VTAIL.t4 VN.t3 VDD2.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=0.6336 pd=4.17 as=0.6336 ps=4.17 w=3.84 l=1.02
X10 VDD2.t5 VN.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.6336 pd=4.17 as=0.6336 ps=4.17 w=3.84 l=1.02
X11 VTAIL.t14 VP.t4 VDD1.t5 B.t23 sky130_fd_pr__nfet_01v8 ad=0.6336 pd=4.17 as=0.6336 ps=4.17 w=3.84 l=1.02
X12 VDD1.t8 VP.t5 VTAIL.t13 B.t7 sky130_fd_pr__nfet_01v8 ad=0.6336 pd=4.17 as=0.6336 ps=4.17 w=3.84 l=1.02
X13 VDD1.t0 VP.t6 VTAIL.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=8.46 as=0.6336 ps=4.17 w=3.84 l=1.02
X14 VDD2.t4 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.6336 pd=4.17 as=1.4976 ps=8.46 w=3.84 l=1.02
X15 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=8.46 as=0 ps=0 w=3.84 l=1.02
X16 VDD1.t3 VP.t7 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=0.6336 pd=4.17 as=1.4976 ps=8.46 w=3.84 l=1.02
X17 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=8.46 as=0 ps=0 w=3.84 l=1.02
X18 VDD2.t3 VN.t6 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=8.46 as=0.6336 ps=4.17 w=3.84 l=1.02
X19 VTAIL.t10 VP.t8 VDD1.t2 B.t6 sky130_fd_pr__nfet_01v8 ad=0.6336 pd=4.17 as=0.6336 ps=4.17 w=3.84 l=1.02
X20 VDD2.t2 VN.t7 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=1.4976 pd=8.46 as=0.6336 ps=4.17 w=3.84 l=1.02
X21 VTAIL.t6 VN.t8 VDD2.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=0.6336 pd=4.17 as=0.6336 ps=4.17 w=3.84 l=1.02
X22 VTAIL.t5 VN.t9 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=0.6336 pd=4.17 as=0.6336 ps=4.17 w=3.84 l=1.02
X23 VDD1.t1 VP.t9 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=0.6336 pd=4.17 as=1.4976 ps=8.46 w=3.84 l=1.02
R0 VP.n10 VP.n7 161.3
R1 VP.n12 VP.n11 161.3
R2 VP.n13 VP.n6 161.3
R3 VP.n16 VP.n15 161.3
R4 VP.n17 VP.n5 161.3
R5 VP.n19 VP.n18 161.3
R6 VP.n21 VP.n4 161.3
R7 VP.n40 VP.n0 161.3
R8 VP.n38 VP.n37 161.3
R9 VP.n36 VP.n1 161.3
R10 VP.n35 VP.n34 161.3
R11 VP.n32 VP.n2 161.3
R12 VP.n31 VP.n30 161.3
R13 VP.n29 VP.n3 161.3
R14 VP.n28 VP.n27 161.3
R15 VP.n9 VP.t6 143.904
R16 VP.n25 VP.t2 129.243
R17 VP.n41 VP.t9 129.243
R18 VP.n22 VP.t7 129.243
R19 VP.n26 VP.t0 90.7299
R20 VP.n33 VP.t5 90.7299
R21 VP.n39 VP.t3 90.7299
R22 VP.n20 VP.t8 90.7299
R23 VP.n14 VP.t1 90.7299
R24 VP.n8 VP.t4 90.7299
R25 VP.n23 VP.n22 80.6037
R26 VP.n42 VP.n41 80.6037
R27 VP.n25 VP.n24 80.6037
R28 VP.n27 VP.n25 53.6107
R29 VP.n41 VP.n40 53.6107
R30 VP.n22 VP.n21 53.6107
R31 VP.n9 VP.n8 48.9084
R32 VP.n32 VP.n31 47.8428
R33 VP.n34 VP.n1 47.8428
R34 VP.n15 VP.n5 47.8428
R35 VP.n13 VP.n12 47.8428
R36 VP.n10 VP.n9 44.2988
R37 VP.n24 VP.n23 38.5279
R38 VP.n31 VP.n3 33.3113
R39 VP.n38 VP.n1 33.3113
R40 VP.n19 VP.n5 33.3113
R41 VP.n12 VP.n7 33.3113
R42 VP.n27 VP.n26 19.674
R43 VP.n40 VP.n39 19.674
R44 VP.n21 VP.n20 19.674
R45 VP.n33 VP.n32 12.2964
R46 VP.n34 VP.n33 12.2964
R47 VP.n14 VP.n13 12.2964
R48 VP.n15 VP.n14 12.2964
R49 VP.n26 VP.n3 4.91887
R50 VP.n39 VP.n38 4.91887
R51 VP.n20 VP.n19 4.91887
R52 VP.n8 VP.n7 4.91887
R53 VP.n23 VP.n4 0.285035
R54 VP.n28 VP.n24 0.285035
R55 VP.n42 VP.n0 0.285035
R56 VP.n11 VP.n10 0.189894
R57 VP.n11 VP.n6 0.189894
R58 VP.n16 VP.n6 0.189894
R59 VP.n17 VP.n16 0.189894
R60 VP.n18 VP.n17 0.189894
R61 VP.n18 VP.n4 0.189894
R62 VP.n29 VP.n28 0.189894
R63 VP.n30 VP.n29 0.189894
R64 VP.n30 VP.n2 0.189894
R65 VP.n35 VP.n2 0.189894
R66 VP.n36 VP.n35 0.189894
R67 VP.n37 VP.n36 0.189894
R68 VP.n37 VP.n0 0.189894
R69 VP VP.n42 0.146778
R70 VDD1.n14 VDD1.n0 289.615
R71 VDD1.n35 VDD1.n21 289.615
R72 VDD1.n15 VDD1.n14 185
R73 VDD1.n13 VDD1.n12 185
R74 VDD1.n4 VDD1.n3 185
R75 VDD1.n7 VDD1.n6 185
R76 VDD1.n28 VDD1.n27 185
R77 VDD1.n25 VDD1.n24 185
R78 VDD1.n34 VDD1.n33 185
R79 VDD1.n36 VDD1.n35 185
R80 VDD1.t0 VDD1.n5 147.888
R81 VDD1.t6 VDD1.n26 147.888
R82 VDD1.n14 VDD1.n13 104.615
R83 VDD1.n13 VDD1.n3 104.615
R84 VDD1.n6 VDD1.n3 104.615
R85 VDD1.n27 VDD1.n24 104.615
R86 VDD1.n34 VDD1.n24 104.615
R87 VDD1.n35 VDD1.n34 104.615
R88 VDD1.n43 VDD1.n42 74.2815
R89 VDD1.n20 VDD1.n19 73.4641
R90 VDD1.n45 VDD1.n44 73.464
R91 VDD1.n41 VDD1.n40 73.464
R92 VDD1.n6 VDD1.t0 52.3082
R93 VDD1.n27 VDD1.t6 52.3082
R94 VDD1.n20 VDD1.n18 50.0279
R95 VDD1.n41 VDD1.n39 50.0279
R96 VDD1.n45 VDD1.n43 33.7186
R97 VDD1.n7 VDD1.n5 15.6496
R98 VDD1.n28 VDD1.n26 15.6496
R99 VDD1.n8 VDD1.n4 12.8005
R100 VDD1.n29 VDD1.n25 12.8005
R101 VDD1.n12 VDD1.n11 12.0247
R102 VDD1.n33 VDD1.n32 12.0247
R103 VDD1.n15 VDD1.n2 11.249
R104 VDD1.n36 VDD1.n23 11.249
R105 VDD1.n16 VDD1.n0 10.4732
R106 VDD1.n37 VDD1.n21 10.4732
R107 VDD1.n18 VDD1.n17 9.45567
R108 VDD1.n39 VDD1.n38 9.45567
R109 VDD1.n17 VDD1.n16 9.3005
R110 VDD1.n2 VDD1.n1 9.3005
R111 VDD1.n11 VDD1.n10 9.3005
R112 VDD1.n9 VDD1.n8 9.3005
R113 VDD1.n38 VDD1.n37 9.3005
R114 VDD1.n23 VDD1.n22 9.3005
R115 VDD1.n32 VDD1.n31 9.3005
R116 VDD1.n30 VDD1.n29 9.3005
R117 VDD1.n44 VDD1.t2 5.15675
R118 VDD1.n44 VDD1.t3 5.15675
R119 VDD1.n19 VDD1.t5 5.15675
R120 VDD1.n19 VDD1.t4 5.15675
R121 VDD1.n42 VDD1.t7 5.15675
R122 VDD1.n42 VDD1.t1 5.15675
R123 VDD1.n40 VDD1.t9 5.15675
R124 VDD1.n40 VDD1.t8 5.15675
R125 VDD1.n9 VDD1.n5 4.40546
R126 VDD1.n30 VDD1.n26 4.40546
R127 VDD1.n18 VDD1.n0 3.49141
R128 VDD1.n39 VDD1.n21 3.49141
R129 VDD1.n16 VDD1.n15 2.71565
R130 VDD1.n37 VDD1.n36 2.71565
R131 VDD1.n12 VDD1.n2 1.93989
R132 VDD1.n33 VDD1.n23 1.93989
R133 VDD1.n11 VDD1.n4 1.16414
R134 VDD1.n32 VDD1.n25 1.16414
R135 VDD1 VDD1.n45 0.815155
R136 VDD1.n8 VDD1.n7 0.388379
R137 VDD1.n29 VDD1.n28 0.388379
R138 VDD1 VDD1.n20 0.349638
R139 VDD1.n43 VDD1.n41 0.236102
R140 VDD1.n17 VDD1.n1 0.155672
R141 VDD1.n10 VDD1.n1 0.155672
R142 VDD1.n10 VDD1.n9 0.155672
R143 VDD1.n31 VDD1.n30 0.155672
R144 VDD1.n31 VDD1.n22 0.155672
R145 VDD1.n38 VDD1.n22 0.155672
R146 VTAIL.n88 VTAIL.n74 289.615
R147 VTAIL.n16 VTAIL.n2 289.615
R148 VTAIL.n68 VTAIL.n54 289.615
R149 VTAIL.n44 VTAIL.n30 289.615
R150 VTAIL.n81 VTAIL.n80 185
R151 VTAIL.n78 VTAIL.n77 185
R152 VTAIL.n87 VTAIL.n86 185
R153 VTAIL.n89 VTAIL.n88 185
R154 VTAIL.n9 VTAIL.n8 185
R155 VTAIL.n6 VTAIL.n5 185
R156 VTAIL.n15 VTAIL.n14 185
R157 VTAIL.n17 VTAIL.n16 185
R158 VTAIL.n69 VTAIL.n68 185
R159 VTAIL.n67 VTAIL.n66 185
R160 VTAIL.n58 VTAIL.n57 185
R161 VTAIL.n61 VTAIL.n60 185
R162 VTAIL.n45 VTAIL.n44 185
R163 VTAIL.n43 VTAIL.n42 185
R164 VTAIL.n34 VTAIL.n33 185
R165 VTAIL.n37 VTAIL.n36 185
R166 VTAIL.t3 VTAIL.n79 147.888
R167 VTAIL.t9 VTAIL.n7 147.888
R168 VTAIL.t11 VTAIL.n59 147.888
R169 VTAIL.t0 VTAIL.n35 147.888
R170 VTAIL.n80 VTAIL.n77 104.615
R171 VTAIL.n87 VTAIL.n77 104.615
R172 VTAIL.n88 VTAIL.n87 104.615
R173 VTAIL.n8 VTAIL.n5 104.615
R174 VTAIL.n15 VTAIL.n5 104.615
R175 VTAIL.n16 VTAIL.n15 104.615
R176 VTAIL.n68 VTAIL.n67 104.615
R177 VTAIL.n67 VTAIL.n57 104.615
R178 VTAIL.n60 VTAIL.n57 104.615
R179 VTAIL.n44 VTAIL.n43 104.615
R180 VTAIL.n43 VTAIL.n33 104.615
R181 VTAIL.n36 VTAIL.n33 104.615
R182 VTAIL.n53 VTAIL.n52 56.7853
R183 VTAIL.n51 VTAIL.n50 56.7853
R184 VTAIL.n29 VTAIL.n28 56.7853
R185 VTAIL.n27 VTAIL.n26 56.7853
R186 VTAIL.n95 VTAIL.n94 56.7852
R187 VTAIL.n1 VTAIL.n0 56.7852
R188 VTAIL.n23 VTAIL.n22 56.7852
R189 VTAIL.n25 VTAIL.n24 56.7852
R190 VTAIL.n80 VTAIL.t3 52.3082
R191 VTAIL.n8 VTAIL.t9 52.3082
R192 VTAIL.n60 VTAIL.t11 52.3082
R193 VTAIL.n36 VTAIL.t0 52.3082
R194 VTAIL.n93 VTAIL.n92 32.1853
R195 VTAIL.n21 VTAIL.n20 32.1853
R196 VTAIL.n73 VTAIL.n72 32.1853
R197 VTAIL.n49 VTAIL.n48 32.1853
R198 VTAIL.n27 VTAIL.n25 18.0048
R199 VTAIL.n93 VTAIL.n73 16.841
R200 VTAIL.n81 VTAIL.n79 15.6496
R201 VTAIL.n9 VTAIL.n7 15.6496
R202 VTAIL.n61 VTAIL.n59 15.6496
R203 VTAIL.n37 VTAIL.n35 15.6496
R204 VTAIL.n82 VTAIL.n78 12.8005
R205 VTAIL.n10 VTAIL.n6 12.8005
R206 VTAIL.n62 VTAIL.n58 12.8005
R207 VTAIL.n38 VTAIL.n34 12.8005
R208 VTAIL.n86 VTAIL.n85 12.0247
R209 VTAIL.n14 VTAIL.n13 12.0247
R210 VTAIL.n66 VTAIL.n65 12.0247
R211 VTAIL.n42 VTAIL.n41 12.0247
R212 VTAIL.n89 VTAIL.n76 11.249
R213 VTAIL.n17 VTAIL.n4 11.249
R214 VTAIL.n69 VTAIL.n56 11.249
R215 VTAIL.n45 VTAIL.n32 11.249
R216 VTAIL.n90 VTAIL.n74 10.4732
R217 VTAIL.n18 VTAIL.n2 10.4732
R218 VTAIL.n70 VTAIL.n54 10.4732
R219 VTAIL.n46 VTAIL.n30 10.4732
R220 VTAIL.n92 VTAIL.n91 9.45567
R221 VTAIL.n20 VTAIL.n19 9.45567
R222 VTAIL.n72 VTAIL.n71 9.45567
R223 VTAIL.n48 VTAIL.n47 9.45567
R224 VTAIL.n91 VTAIL.n90 9.3005
R225 VTAIL.n76 VTAIL.n75 9.3005
R226 VTAIL.n85 VTAIL.n84 9.3005
R227 VTAIL.n83 VTAIL.n82 9.3005
R228 VTAIL.n19 VTAIL.n18 9.3005
R229 VTAIL.n4 VTAIL.n3 9.3005
R230 VTAIL.n13 VTAIL.n12 9.3005
R231 VTAIL.n11 VTAIL.n10 9.3005
R232 VTAIL.n71 VTAIL.n70 9.3005
R233 VTAIL.n56 VTAIL.n55 9.3005
R234 VTAIL.n65 VTAIL.n64 9.3005
R235 VTAIL.n63 VTAIL.n62 9.3005
R236 VTAIL.n47 VTAIL.n46 9.3005
R237 VTAIL.n32 VTAIL.n31 9.3005
R238 VTAIL.n41 VTAIL.n40 9.3005
R239 VTAIL.n39 VTAIL.n38 9.3005
R240 VTAIL.n94 VTAIL.t2 5.15675
R241 VTAIL.n94 VTAIL.t6 5.15675
R242 VTAIL.n0 VTAIL.t1 5.15675
R243 VTAIL.n0 VTAIL.t19 5.15675
R244 VTAIL.n22 VTAIL.t13 5.15675
R245 VTAIL.n22 VTAIL.t15 5.15675
R246 VTAIL.n24 VTAIL.t16 5.15675
R247 VTAIL.n24 VTAIL.t18 5.15675
R248 VTAIL.n52 VTAIL.t17 5.15675
R249 VTAIL.n52 VTAIL.t10 5.15675
R250 VTAIL.n50 VTAIL.t12 5.15675
R251 VTAIL.n50 VTAIL.t14 5.15675
R252 VTAIL.n28 VTAIL.t7 5.15675
R253 VTAIL.n28 VTAIL.t4 5.15675
R254 VTAIL.n26 VTAIL.t8 5.15675
R255 VTAIL.n26 VTAIL.t5 5.15675
R256 VTAIL.n83 VTAIL.n79 4.40546
R257 VTAIL.n11 VTAIL.n7 4.40546
R258 VTAIL.n63 VTAIL.n59 4.40546
R259 VTAIL.n39 VTAIL.n35 4.40546
R260 VTAIL.n92 VTAIL.n74 3.49141
R261 VTAIL.n20 VTAIL.n2 3.49141
R262 VTAIL.n72 VTAIL.n54 3.49141
R263 VTAIL.n48 VTAIL.n30 3.49141
R264 VTAIL.n90 VTAIL.n89 2.71565
R265 VTAIL.n18 VTAIL.n17 2.71565
R266 VTAIL.n70 VTAIL.n69 2.71565
R267 VTAIL.n46 VTAIL.n45 2.71565
R268 VTAIL.n86 VTAIL.n76 1.93989
R269 VTAIL.n14 VTAIL.n4 1.93989
R270 VTAIL.n66 VTAIL.n56 1.93989
R271 VTAIL.n42 VTAIL.n32 1.93989
R272 VTAIL.n29 VTAIL.n27 1.16429
R273 VTAIL.n49 VTAIL.n29 1.16429
R274 VTAIL.n53 VTAIL.n51 1.16429
R275 VTAIL.n73 VTAIL.n53 1.16429
R276 VTAIL.n25 VTAIL.n23 1.16429
R277 VTAIL.n23 VTAIL.n21 1.16429
R278 VTAIL.n95 VTAIL.n93 1.16429
R279 VTAIL.n85 VTAIL.n78 1.16414
R280 VTAIL.n13 VTAIL.n6 1.16414
R281 VTAIL.n65 VTAIL.n58 1.16414
R282 VTAIL.n41 VTAIL.n34 1.16414
R283 VTAIL.n51 VTAIL.n49 1.05222
R284 VTAIL.n21 VTAIL.n1 1.05222
R285 VTAIL VTAIL.n1 0.931535
R286 VTAIL.n82 VTAIL.n81 0.388379
R287 VTAIL.n10 VTAIL.n9 0.388379
R288 VTAIL.n62 VTAIL.n61 0.388379
R289 VTAIL.n38 VTAIL.n37 0.388379
R290 VTAIL VTAIL.n95 0.233259
R291 VTAIL.n84 VTAIL.n83 0.155672
R292 VTAIL.n84 VTAIL.n75 0.155672
R293 VTAIL.n91 VTAIL.n75 0.155672
R294 VTAIL.n12 VTAIL.n11 0.155672
R295 VTAIL.n12 VTAIL.n3 0.155672
R296 VTAIL.n19 VTAIL.n3 0.155672
R297 VTAIL.n71 VTAIL.n55 0.155672
R298 VTAIL.n64 VTAIL.n55 0.155672
R299 VTAIL.n64 VTAIL.n63 0.155672
R300 VTAIL.n47 VTAIL.n31 0.155672
R301 VTAIL.n40 VTAIL.n31 0.155672
R302 VTAIL.n40 VTAIL.n39 0.155672
R303 B.n494 B.n493 585
R304 B.n495 B.n494 585
R305 B.n175 B.n84 585
R306 B.n174 B.n173 585
R307 B.n172 B.n171 585
R308 B.n170 B.n169 585
R309 B.n168 B.n167 585
R310 B.n166 B.n165 585
R311 B.n164 B.n163 585
R312 B.n162 B.n161 585
R313 B.n160 B.n159 585
R314 B.n158 B.n157 585
R315 B.n156 B.n155 585
R316 B.n154 B.n153 585
R317 B.n152 B.n151 585
R318 B.n150 B.n149 585
R319 B.n148 B.n147 585
R320 B.n146 B.n145 585
R321 B.n144 B.n143 585
R322 B.n141 B.n140 585
R323 B.n139 B.n138 585
R324 B.n137 B.n136 585
R325 B.n135 B.n134 585
R326 B.n133 B.n132 585
R327 B.n131 B.n130 585
R328 B.n129 B.n128 585
R329 B.n127 B.n126 585
R330 B.n125 B.n124 585
R331 B.n123 B.n122 585
R332 B.n121 B.n120 585
R333 B.n119 B.n118 585
R334 B.n117 B.n116 585
R335 B.n115 B.n114 585
R336 B.n113 B.n112 585
R337 B.n111 B.n110 585
R338 B.n109 B.n108 585
R339 B.n107 B.n106 585
R340 B.n105 B.n104 585
R341 B.n103 B.n102 585
R342 B.n101 B.n100 585
R343 B.n99 B.n98 585
R344 B.n97 B.n96 585
R345 B.n95 B.n94 585
R346 B.n93 B.n92 585
R347 B.n91 B.n90 585
R348 B.n60 B.n59 585
R349 B.n492 B.n61 585
R350 B.n496 B.n61 585
R351 B.n491 B.n490 585
R352 B.n490 B.n57 585
R353 B.n489 B.n56 585
R354 B.n502 B.n56 585
R355 B.n488 B.n55 585
R356 B.n503 B.n55 585
R357 B.n487 B.n54 585
R358 B.n504 B.n54 585
R359 B.n486 B.n485 585
R360 B.n485 B.n53 585
R361 B.n484 B.n49 585
R362 B.n510 B.n49 585
R363 B.n483 B.n48 585
R364 B.n511 B.n48 585
R365 B.n482 B.n47 585
R366 B.n512 B.n47 585
R367 B.n481 B.n480 585
R368 B.n480 B.n43 585
R369 B.n479 B.n42 585
R370 B.n518 B.n42 585
R371 B.n478 B.n41 585
R372 B.n519 B.n41 585
R373 B.n477 B.n40 585
R374 B.n520 B.n40 585
R375 B.n476 B.n475 585
R376 B.n475 B.n36 585
R377 B.n474 B.n35 585
R378 B.n526 B.n35 585
R379 B.n473 B.n34 585
R380 B.n527 B.n34 585
R381 B.n472 B.n33 585
R382 B.n528 B.n33 585
R383 B.n471 B.n470 585
R384 B.n470 B.n29 585
R385 B.n469 B.n28 585
R386 B.n534 B.n28 585
R387 B.n468 B.n27 585
R388 B.n535 B.n27 585
R389 B.n467 B.n26 585
R390 B.n536 B.n26 585
R391 B.n466 B.n465 585
R392 B.n465 B.n22 585
R393 B.n464 B.n21 585
R394 B.n542 B.n21 585
R395 B.n463 B.n20 585
R396 B.n543 B.n20 585
R397 B.n462 B.n19 585
R398 B.n544 B.n19 585
R399 B.n461 B.n460 585
R400 B.n460 B.n15 585
R401 B.n459 B.n14 585
R402 B.n550 B.n14 585
R403 B.n458 B.n13 585
R404 B.n551 B.n13 585
R405 B.n457 B.n12 585
R406 B.n552 B.n12 585
R407 B.n456 B.n455 585
R408 B.n455 B.n8 585
R409 B.n454 B.n7 585
R410 B.n558 B.n7 585
R411 B.n453 B.n6 585
R412 B.n559 B.n6 585
R413 B.n452 B.n5 585
R414 B.n560 B.n5 585
R415 B.n451 B.n450 585
R416 B.n450 B.n4 585
R417 B.n449 B.n176 585
R418 B.n449 B.n448 585
R419 B.n439 B.n177 585
R420 B.n178 B.n177 585
R421 B.n441 B.n440 585
R422 B.n442 B.n441 585
R423 B.n438 B.n183 585
R424 B.n183 B.n182 585
R425 B.n437 B.n436 585
R426 B.n436 B.n435 585
R427 B.n185 B.n184 585
R428 B.n186 B.n185 585
R429 B.n428 B.n427 585
R430 B.n429 B.n428 585
R431 B.n426 B.n191 585
R432 B.n191 B.n190 585
R433 B.n425 B.n424 585
R434 B.n424 B.n423 585
R435 B.n193 B.n192 585
R436 B.n194 B.n193 585
R437 B.n416 B.n415 585
R438 B.n417 B.n416 585
R439 B.n414 B.n199 585
R440 B.n199 B.n198 585
R441 B.n413 B.n412 585
R442 B.n412 B.n411 585
R443 B.n201 B.n200 585
R444 B.n202 B.n201 585
R445 B.n404 B.n403 585
R446 B.n405 B.n404 585
R447 B.n402 B.n207 585
R448 B.n207 B.n206 585
R449 B.n401 B.n400 585
R450 B.n400 B.n399 585
R451 B.n209 B.n208 585
R452 B.n210 B.n209 585
R453 B.n392 B.n391 585
R454 B.n393 B.n392 585
R455 B.n390 B.n215 585
R456 B.n215 B.n214 585
R457 B.n389 B.n388 585
R458 B.n388 B.n387 585
R459 B.n217 B.n216 585
R460 B.n218 B.n217 585
R461 B.n380 B.n379 585
R462 B.n381 B.n380 585
R463 B.n378 B.n223 585
R464 B.n223 B.n222 585
R465 B.n377 B.n376 585
R466 B.n376 B.n375 585
R467 B.n225 B.n224 585
R468 B.n368 B.n225 585
R469 B.n367 B.n366 585
R470 B.n369 B.n367 585
R471 B.n365 B.n230 585
R472 B.n230 B.n229 585
R473 B.n364 B.n363 585
R474 B.n363 B.n362 585
R475 B.n232 B.n231 585
R476 B.n233 B.n232 585
R477 B.n355 B.n354 585
R478 B.n356 B.n355 585
R479 B.n236 B.n235 585
R480 B.n265 B.n263 585
R481 B.n266 B.n262 585
R482 B.n266 B.n237 585
R483 B.n269 B.n268 585
R484 B.n270 B.n261 585
R485 B.n272 B.n271 585
R486 B.n274 B.n260 585
R487 B.n277 B.n276 585
R488 B.n278 B.n259 585
R489 B.n280 B.n279 585
R490 B.n282 B.n258 585
R491 B.n285 B.n284 585
R492 B.n286 B.n257 585
R493 B.n288 B.n287 585
R494 B.n290 B.n256 585
R495 B.n293 B.n292 585
R496 B.n294 B.n255 585
R497 B.n299 B.n298 585
R498 B.n301 B.n254 585
R499 B.n304 B.n303 585
R500 B.n305 B.n253 585
R501 B.n307 B.n306 585
R502 B.n309 B.n252 585
R503 B.n312 B.n311 585
R504 B.n313 B.n251 585
R505 B.n315 B.n314 585
R506 B.n317 B.n250 585
R507 B.n320 B.n319 585
R508 B.n321 B.n246 585
R509 B.n323 B.n322 585
R510 B.n325 B.n245 585
R511 B.n328 B.n327 585
R512 B.n329 B.n244 585
R513 B.n331 B.n330 585
R514 B.n333 B.n243 585
R515 B.n336 B.n335 585
R516 B.n337 B.n242 585
R517 B.n339 B.n338 585
R518 B.n341 B.n241 585
R519 B.n344 B.n343 585
R520 B.n345 B.n240 585
R521 B.n347 B.n346 585
R522 B.n349 B.n239 585
R523 B.n352 B.n351 585
R524 B.n353 B.n238 585
R525 B.n358 B.n357 585
R526 B.n357 B.n356 585
R527 B.n359 B.n234 585
R528 B.n234 B.n233 585
R529 B.n361 B.n360 585
R530 B.n362 B.n361 585
R531 B.n228 B.n227 585
R532 B.n229 B.n228 585
R533 B.n371 B.n370 585
R534 B.n370 B.n369 585
R535 B.n372 B.n226 585
R536 B.n368 B.n226 585
R537 B.n374 B.n373 585
R538 B.n375 B.n374 585
R539 B.n221 B.n220 585
R540 B.n222 B.n221 585
R541 B.n383 B.n382 585
R542 B.n382 B.n381 585
R543 B.n384 B.n219 585
R544 B.n219 B.n218 585
R545 B.n386 B.n385 585
R546 B.n387 B.n386 585
R547 B.n213 B.n212 585
R548 B.n214 B.n213 585
R549 B.n395 B.n394 585
R550 B.n394 B.n393 585
R551 B.n396 B.n211 585
R552 B.n211 B.n210 585
R553 B.n398 B.n397 585
R554 B.n399 B.n398 585
R555 B.n205 B.n204 585
R556 B.n206 B.n205 585
R557 B.n407 B.n406 585
R558 B.n406 B.n405 585
R559 B.n408 B.n203 585
R560 B.n203 B.n202 585
R561 B.n410 B.n409 585
R562 B.n411 B.n410 585
R563 B.n197 B.n196 585
R564 B.n198 B.n197 585
R565 B.n419 B.n418 585
R566 B.n418 B.n417 585
R567 B.n420 B.n195 585
R568 B.n195 B.n194 585
R569 B.n422 B.n421 585
R570 B.n423 B.n422 585
R571 B.n189 B.n188 585
R572 B.n190 B.n189 585
R573 B.n431 B.n430 585
R574 B.n430 B.n429 585
R575 B.n432 B.n187 585
R576 B.n187 B.n186 585
R577 B.n434 B.n433 585
R578 B.n435 B.n434 585
R579 B.n181 B.n180 585
R580 B.n182 B.n181 585
R581 B.n444 B.n443 585
R582 B.n443 B.n442 585
R583 B.n445 B.n179 585
R584 B.n179 B.n178 585
R585 B.n447 B.n446 585
R586 B.n448 B.n447 585
R587 B.n2 B.n0 585
R588 B.n4 B.n2 585
R589 B.n3 B.n1 585
R590 B.n559 B.n3 585
R591 B.n557 B.n556 585
R592 B.n558 B.n557 585
R593 B.n555 B.n9 585
R594 B.n9 B.n8 585
R595 B.n554 B.n553 585
R596 B.n553 B.n552 585
R597 B.n11 B.n10 585
R598 B.n551 B.n11 585
R599 B.n549 B.n548 585
R600 B.n550 B.n549 585
R601 B.n547 B.n16 585
R602 B.n16 B.n15 585
R603 B.n546 B.n545 585
R604 B.n545 B.n544 585
R605 B.n18 B.n17 585
R606 B.n543 B.n18 585
R607 B.n541 B.n540 585
R608 B.n542 B.n541 585
R609 B.n539 B.n23 585
R610 B.n23 B.n22 585
R611 B.n538 B.n537 585
R612 B.n537 B.n536 585
R613 B.n25 B.n24 585
R614 B.n535 B.n25 585
R615 B.n533 B.n532 585
R616 B.n534 B.n533 585
R617 B.n531 B.n30 585
R618 B.n30 B.n29 585
R619 B.n530 B.n529 585
R620 B.n529 B.n528 585
R621 B.n32 B.n31 585
R622 B.n527 B.n32 585
R623 B.n525 B.n524 585
R624 B.n526 B.n525 585
R625 B.n523 B.n37 585
R626 B.n37 B.n36 585
R627 B.n522 B.n521 585
R628 B.n521 B.n520 585
R629 B.n39 B.n38 585
R630 B.n519 B.n39 585
R631 B.n517 B.n516 585
R632 B.n518 B.n517 585
R633 B.n515 B.n44 585
R634 B.n44 B.n43 585
R635 B.n514 B.n513 585
R636 B.n513 B.n512 585
R637 B.n46 B.n45 585
R638 B.n511 B.n46 585
R639 B.n509 B.n508 585
R640 B.n510 B.n509 585
R641 B.n507 B.n50 585
R642 B.n53 B.n50 585
R643 B.n506 B.n505 585
R644 B.n505 B.n504 585
R645 B.n52 B.n51 585
R646 B.n503 B.n52 585
R647 B.n501 B.n500 585
R648 B.n502 B.n501 585
R649 B.n499 B.n58 585
R650 B.n58 B.n57 585
R651 B.n498 B.n497 585
R652 B.n497 B.n496 585
R653 B.n562 B.n561 585
R654 B.n561 B.n560 585
R655 B.n357 B.n236 473.281
R656 B.n497 B.n60 473.281
R657 B.n355 B.n238 473.281
R658 B.n494 B.n61 473.281
R659 B.n247 B.t13 293.789
R660 B.n295 B.t17 293.789
R661 B.n87 B.t20 293.789
R662 B.n85 B.t9 293.789
R663 B.n495 B.n83 256.663
R664 B.n495 B.n82 256.663
R665 B.n495 B.n81 256.663
R666 B.n495 B.n80 256.663
R667 B.n495 B.n79 256.663
R668 B.n495 B.n78 256.663
R669 B.n495 B.n77 256.663
R670 B.n495 B.n76 256.663
R671 B.n495 B.n75 256.663
R672 B.n495 B.n74 256.663
R673 B.n495 B.n73 256.663
R674 B.n495 B.n72 256.663
R675 B.n495 B.n71 256.663
R676 B.n495 B.n70 256.663
R677 B.n495 B.n69 256.663
R678 B.n495 B.n68 256.663
R679 B.n495 B.n67 256.663
R680 B.n495 B.n66 256.663
R681 B.n495 B.n65 256.663
R682 B.n495 B.n64 256.663
R683 B.n495 B.n63 256.663
R684 B.n495 B.n62 256.663
R685 B.n264 B.n237 256.663
R686 B.n267 B.n237 256.663
R687 B.n273 B.n237 256.663
R688 B.n275 B.n237 256.663
R689 B.n281 B.n237 256.663
R690 B.n283 B.n237 256.663
R691 B.n289 B.n237 256.663
R692 B.n291 B.n237 256.663
R693 B.n300 B.n237 256.663
R694 B.n302 B.n237 256.663
R695 B.n308 B.n237 256.663
R696 B.n310 B.n237 256.663
R697 B.n316 B.n237 256.663
R698 B.n318 B.n237 256.663
R699 B.n324 B.n237 256.663
R700 B.n326 B.n237 256.663
R701 B.n332 B.n237 256.663
R702 B.n334 B.n237 256.663
R703 B.n340 B.n237 256.663
R704 B.n342 B.n237 256.663
R705 B.n348 B.n237 256.663
R706 B.n350 B.n237 256.663
R707 B.n247 B.t16 168.339
R708 B.n85 B.t11 168.339
R709 B.n295 B.t19 168.339
R710 B.n87 B.t21 168.339
R711 B.n357 B.n234 163.367
R712 B.n361 B.n234 163.367
R713 B.n361 B.n228 163.367
R714 B.n370 B.n228 163.367
R715 B.n370 B.n226 163.367
R716 B.n374 B.n226 163.367
R717 B.n374 B.n221 163.367
R718 B.n382 B.n221 163.367
R719 B.n382 B.n219 163.367
R720 B.n386 B.n219 163.367
R721 B.n386 B.n213 163.367
R722 B.n394 B.n213 163.367
R723 B.n394 B.n211 163.367
R724 B.n398 B.n211 163.367
R725 B.n398 B.n205 163.367
R726 B.n406 B.n205 163.367
R727 B.n406 B.n203 163.367
R728 B.n410 B.n203 163.367
R729 B.n410 B.n197 163.367
R730 B.n418 B.n197 163.367
R731 B.n418 B.n195 163.367
R732 B.n422 B.n195 163.367
R733 B.n422 B.n189 163.367
R734 B.n430 B.n189 163.367
R735 B.n430 B.n187 163.367
R736 B.n434 B.n187 163.367
R737 B.n434 B.n181 163.367
R738 B.n443 B.n181 163.367
R739 B.n443 B.n179 163.367
R740 B.n447 B.n179 163.367
R741 B.n447 B.n2 163.367
R742 B.n561 B.n2 163.367
R743 B.n561 B.n3 163.367
R744 B.n557 B.n3 163.367
R745 B.n557 B.n9 163.367
R746 B.n553 B.n9 163.367
R747 B.n553 B.n11 163.367
R748 B.n549 B.n11 163.367
R749 B.n549 B.n16 163.367
R750 B.n545 B.n16 163.367
R751 B.n545 B.n18 163.367
R752 B.n541 B.n18 163.367
R753 B.n541 B.n23 163.367
R754 B.n537 B.n23 163.367
R755 B.n537 B.n25 163.367
R756 B.n533 B.n25 163.367
R757 B.n533 B.n30 163.367
R758 B.n529 B.n30 163.367
R759 B.n529 B.n32 163.367
R760 B.n525 B.n32 163.367
R761 B.n525 B.n37 163.367
R762 B.n521 B.n37 163.367
R763 B.n521 B.n39 163.367
R764 B.n517 B.n39 163.367
R765 B.n517 B.n44 163.367
R766 B.n513 B.n44 163.367
R767 B.n513 B.n46 163.367
R768 B.n509 B.n46 163.367
R769 B.n509 B.n50 163.367
R770 B.n505 B.n50 163.367
R771 B.n505 B.n52 163.367
R772 B.n501 B.n52 163.367
R773 B.n501 B.n58 163.367
R774 B.n497 B.n58 163.367
R775 B.n266 B.n265 163.367
R776 B.n268 B.n266 163.367
R777 B.n272 B.n261 163.367
R778 B.n276 B.n274 163.367
R779 B.n280 B.n259 163.367
R780 B.n284 B.n282 163.367
R781 B.n288 B.n257 163.367
R782 B.n292 B.n290 163.367
R783 B.n299 B.n255 163.367
R784 B.n303 B.n301 163.367
R785 B.n307 B.n253 163.367
R786 B.n311 B.n309 163.367
R787 B.n315 B.n251 163.367
R788 B.n319 B.n317 163.367
R789 B.n323 B.n246 163.367
R790 B.n327 B.n325 163.367
R791 B.n331 B.n244 163.367
R792 B.n335 B.n333 163.367
R793 B.n339 B.n242 163.367
R794 B.n343 B.n341 163.367
R795 B.n347 B.n240 163.367
R796 B.n351 B.n349 163.367
R797 B.n355 B.n232 163.367
R798 B.n363 B.n232 163.367
R799 B.n363 B.n230 163.367
R800 B.n367 B.n230 163.367
R801 B.n367 B.n225 163.367
R802 B.n376 B.n225 163.367
R803 B.n376 B.n223 163.367
R804 B.n380 B.n223 163.367
R805 B.n380 B.n217 163.367
R806 B.n388 B.n217 163.367
R807 B.n388 B.n215 163.367
R808 B.n392 B.n215 163.367
R809 B.n392 B.n209 163.367
R810 B.n400 B.n209 163.367
R811 B.n400 B.n207 163.367
R812 B.n404 B.n207 163.367
R813 B.n404 B.n201 163.367
R814 B.n412 B.n201 163.367
R815 B.n412 B.n199 163.367
R816 B.n416 B.n199 163.367
R817 B.n416 B.n193 163.367
R818 B.n424 B.n193 163.367
R819 B.n424 B.n191 163.367
R820 B.n428 B.n191 163.367
R821 B.n428 B.n185 163.367
R822 B.n436 B.n185 163.367
R823 B.n436 B.n183 163.367
R824 B.n441 B.n183 163.367
R825 B.n441 B.n177 163.367
R826 B.n449 B.n177 163.367
R827 B.n450 B.n449 163.367
R828 B.n450 B.n5 163.367
R829 B.n6 B.n5 163.367
R830 B.n7 B.n6 163.367
R831 B.n455 B.n7 163.367
R832 B.n455 B.n12 163.367
R833 B.n13 B.n12 163.367
R834 B.n14 B.n13 163.367
R835 B.n460 B.n14 163.367
R836 B.n460 B.n19 163.367
R837 B.n20 B.n19 163.367
R838 B.n21 B.n20 163.367
R839 B.n465 B.n21 163.367
R840 B.n465 B.n26 163.367
R841 B.n27 B.n26 163.367
R842 B.n28 B.n27 163.367
R843 B.n470 B.n28 163.367
R844 B.n470 B.n33 163.367
R845 B.n34 B.n33 163.367
R846 B.n35 B.n34 163.367
R847 B.n475 B.n35 163.367
R848 B.n475 B.n40 163.367
R849 B.n41 B.n40 163.367
R850 B.n42 B.n41 163.367
R851 B.n480 B.n42 163.367
R852 B.n480 B.n47 163.367
R853 B.n48 B.n47 163.367
R854 B.n49 B.n48 163.367
R855 B.n485 B.n49 163.367
R856 B.n485 B.n54 163.367
R857 B.n55 B.n54 163.367
R858 B.n56 B.n55 163.367
R859 B.n490 B.n56 163.367
R860 B.n490 B.n61 163.367
R861 B.n92 B.n91 163.367
R862 B.n96 B.n95 163.367
R863 B.n100 B.n99 163.367
R864 B.n104 B.n103 163.367
R865 B.n108 B.n107 163.367
R866 B.n112 B.n111 163.367
R867 B.n116 B.n115 163.367
R868 B.n120 B.n119 163.367
R869 B.n124 B.n123 163.367
R870 B.n128 B.n127 163.367
R871 B.n132 B.n131 163.367
R872 B.n136 B.n135 163.367
R873 B.n140 B.n139 163.367
R874 B.n145 B.n144 163.367
R875 B.n149 B.n148 163.367
R876 B.n153 B.n152 163.367
R877 B.n157 B.n156 163.367
R878 B.n161 B.n160 163.367
R879 B.n165 B.n164 163.367
R880 B.n169 B.n168 163.367
R881 B.n173 B.n172 163.367
R882 B.n494 B.n84 163.367
R883 B.n356 B.n237 143.609
R884 B.n496 B.n495 143.609
R885 B.n248 B.t15 142.157
R886 B.n86 B.t12 142.157
R887 B.n296 B.t18 142.157
R888 B.n88 B.t22 142.157
R889 B.n356 B.n233 82.063
R890 B.n362 B.n233 82.063
R891 B.n362 B.n229 82.063
R892 B.n369 B.n229 82.063
R893 B.n369 B.n368 82.063
R894 B.n375 B.n222 82.063
R895 B.n381 B.n222 82.063
R896 B.n381 B.n218 82.063
R897 B.n387 B.n218 82.063
R898 B.n387 B.n214 82.063
R899 B.n393 B.n214 82.063
R900 B.n399 B.n210 82.063
R901 B.n399 B.n206 82.063
R902 B.n405 B.n206 82.063
R903 B.n411 B.n202 82.063
R904 B.n411 B.n198 82.063
R905 B.n417 B.n198 82.063
R906 B.n423 B.n194 82.063
R907 B.n423 B.n190 82.063
R908 B.n429 B.n190 82.063
R909 B.n435 B.n186 82.063
R910 B.n435 B.n182 82.063
R911 B.n442 B.n182 82.063
R912 B.n448 B.n178 82.063
R913 B.n448 B.n4 82.063
R914 B.n560 B.n4 82.063
R915 B.n560 B.n559 82.063
R916 B.n559 B.n558 82.063
R917 B.n558 B.n8 82.063
R918 B.n552 B.n551 82.063
R919 B.n551 B.n550 82.063
R920 B.n550 B.n15 82.063
R921 B.n544 B.n543 82.063
R922 B.n543 B.n542 82.063
R923 B.n542 B.n22 82.063
R924 B.n536 B.n535 82.063
R925 B.n535 B.n534 82.063
R926 B.n534 B.n29 82.063
R927 B.n528 B.n527 82.063
R928 B.n527 B.n526 82.063
R929 B.n526 B.n36 82.063
R930 B.n520 B.n519 82.063
R931 B.n519 B.n518 82.063
R932 B.n518 B.n43 82.063
R933 B.n512 B.n43 82.063
R934 B.n512 B.n511 82.063
R935 B.n511 B.n510 82.063
R936 B.n504 B.n53 82.063
R937 B.n504 B.n503 82.063
R938 B.n503 B.n502 82.063
R939 B.n502 B.n57 82.063
R940 B.n496 B.n57 82.063
R941 B.n264 B.n236 71.676
R942 B.n268 B.n267 71.676
R943 B.n273 B.n272 71.676
R944 B.n276 B.n275 71.676
R945 B.n281 B.n280 71.676
R946 B.n284 B.n283 71.676
R947 B.n289 B.n288 71.676
R948 B.n292 B.n291 71.676
R949 B.n300 B.n299 71.676
R950 B.n303 B.n302 71.676
R951 B.n308 B.n307 71.676
R952 B.n311 B.n310 71.676
R953 B.n316 B.n315 71.676
R954 B.n319 B.n318 71.676
R955 B.n324 B.n323 71.676
R956 B.n327 B.n326 71.676
R957 B.n332 B.n331 71.676
R958 B.n335 B.n334 71.676
R959 B.n340 B.n339 71.676
R960 B.n343 B.n342 71.676
R961 B.n348 B.n347 71.676
R962 B.n351 B.n350 71.676
R963 B.n62 B.n60 71.676
R964 B.n92 B.n63 71.676
R965 B.n96 B.n64 71.676
R966 B.n100 B.n65 71.676
R967 B.n104 B.n66 71.676
R968 B.n108 B.n67 71.676
R969 B.n112 B.n68 71.676
R970 B.n116 B.n69 71.676
R971 B.n120 B.n70 71.676
R972 B.n124 B.n71 71.676
R973 B.n128 B.n72 71.676
R974 B.n132 B.n73 71.676
R975 B.n136 B.n74 71.676
R976 B.n140 B.n75 71.676
R977 B.n145 B.n76 71.676
R978 B.n149 B.n77 71.676
R979 B.n153 B.n78 71.676
R980 B.n157 B.n79 71.676
R981 B.n161 B.n80 71.676
R982 B.n165 B.n81 71.676
R983 B.n169 B.n82 71.676
R984 B.n173 B.n83 71.676
R985 B.n84 B.n83 71.676
R986 B.n172 B.n82 71.676
R987 B.n168 B.n81 71.676
R988 B.n164 B.n80 71.676
R989 B.n160 B.n79 71.676
R990 B.n156 B.n78 71.676
R991 B.n152 B.n77 71.676
R992 B.n148 B.n76 71.676
R993 B.n144 B.n75 71.676
R994 B.n139 B.n74 71.676
R995 B.n135 B.n73 71.676
R996 B.n131 B.n72 71.676
R997 B.n127 B.n71 71.676
R998 B.n123 B.n70 71.676
R999 B.n119 B.n69 71.676
R1000 B.n115 B.n68 71.676
R1001 B.n111 B.n67 71.676
R1002 B.n107 B.n66 71.676
R1003 B.n103 B.n65 71.676
R1004 B.n99 B.n64 71.676
R1005 B.n95 B.n63 71.676
R1006 B.n91 B.n62 71.676
R1007 B.n265 B.n264 71.676
R1008 B.n267 B.n261 71.676
R1009 B.n274 B.n273 71.676
R1010 B.n275 B.n259 71.676
R1011 B.n282 B.n281 71.676
R1012 B.n283 B.n257 71.676
R1013 B.n290 B.n289 71.676
R1014 B.n291 B.n255 71.676
R1015 B.n301 B.n300 71.676
R1016 B.n302 B.n253 71.676
R1017 B.n309 B.n308 71.676
R1018 B.n310 B.n251 71.676
R1019 B.n317 B.n316 71.676
R1020 B.n318 B.n246 71.676
R1021 B.n325 B.n324 71.676
R1022 B.n326 B.n244 71.676
R1023 B.n333 B.n332 71.676
R1024 B.n334 B.n242 71.676
R1025 B.n341 B.n340 71.676
R1026 B.n342 B.n240 71.676
R1027 B.n349 B.n348 71.676
R1028 B.n350 B.n238 71.676
R1029 B.n249 B.n248 59.5399
R1030 B.n297 B.n296 59.5399
R1031 B.n89 B.n88 59.5399
R1032 B.n142 B.n86 59.5399
R1033 B.n375 B.t14 53.0998
R1034 B.n510 B.t10 53.0998
R1035 B.t0 B.n178 48.2726
R1036 B.t1 B.n8 48.2726
R1037 B.t4 B.n186 45.859
R1038 B.t23 B.n15 45.859
R1039 B.n393 B.t8 43.4454
R1040 B.t7 B.n194 43.4454
R1041 B.t2 B.n22 43.4454
R1042 B.n520 B.t3 43.4454
R1043 B.n405 B.t5 41.0318
R1044 B.t5 B.n202 41.0318
R1045 B.t6 B.n29 41.0318
R1046 B.n528 B.t6 41.0318
R1047 B.t8 B.n210 38.6182
R1048 B.n417 B.t7 38.6182
R1049 B.n536 B.t2 38.6182
R1050 B.t3 B.n36 38.6182
R1051 B.n429 B.t4 36.2046
R1052 B.n544 B.t23 36.2046
R1053 B.n442 B.t0 33.791
R1054 B.n552 B.t1 33.791
R1055 B.n498 B.n59 30.7517
R1056 B.n493 B.n492 30.7517
R1057 B.n354 B.n353 30.7517
R1058 B.n358 B.n235 30.7517
R1059 B.n368 B.t14 28.9637
R1060 B.n53 B.t10 28.9637
R1061 B.n248 B.n247 26.1823
R1062 B.n296 B.n295 26.1823
R1063 B.n88 B.n87 26.1823
R1064 B.n86 B.n85 26.1823
R1065 B B.n562 18.0485
R1066 B.n90 B.n59 10.6151
R1067 B.n93 B.n90 10.6151
R1068 B.n94 B.n93 10.6151
R1069 B.n97 B.n94 10.6151
R1070 B.n98 B.n97 10.6151
R1071 B.n101 B.n98 10.6151
R1072 B.n102 B.n101 10.6151
R1073 B.n105 B.n102 10.6151
R1074 B.n106 B.n105 10.6151
R1075 B.n109 B.n106 10.6151
R1076 B.n110 B.n109 10.6151
R1077 B.n113 B.n110 10.6151
R1078 B.n114 B.n113 10.6151
R1079 B.n117 B.n114 10.6151
R1080 B.n118 B.n117 10.6151
R1081 B.n121 B.n118 10.6151
R1082 B.n122 B.n121 10.6151
R1083 B.n126 B.n125 10.6151
R1084 B.n129 B.n126 10.6151
R1085 B.n130 B.n129 10.6151
R1086 B.n133 B.n130 10.6151
R1087 B.n134 B.n133 10.6151
R1088 B.n137 B.n134 10.6151
R1089 B.n138 B.n137 10.6151
R1090 B.n141 B.n138 10.6151
R1091 B.n146 B.n143 10.6151
R1092 B.n147 B.n146 10.6151
R1093 B.n150 B.n147 10.6151
R1094 B.n151 B.n150 10.6151
R1095 B.n154 B.n151 10.6151
R1096 B.n155 B.n154 10.6151
R1097 B.n158 B.n155 10.6151
R1098 B.n159 B.n158 10.6151
R1099 B.n162 B.n159 10.6151
R1100 B.n163 B.n162 10.6151
R1101 B.n166 B.n163 10.6151
R1102 B.n167 B.n166 10.6151
R1103 B.n170 B.n167 10.6151
R1104 B.n171 B.n170 10.6151
R1105 B.n174 B.n171 10.6151
R1106 B.n175 B.n174 10.6151
R1107 B.n493 B.n175 10.6151
R1108 B.n354 B.n231 10.6151
R1109 B.n364 B.n231 10.6151
R1110 B.n365 B.n364 10.6151
R1111 B.n366 B.n365 10.6151
R1112 B.n366 B.n224 10.6151
R1113 B.n377 B.n224 10.6151
R1114 B.n378 B.n377 10.6151
R1115 B.n379 B.n378 10.6151
R1116 B.n379 B.n216 10.6151
R1117 B.n389 B.n216 10.6151
R1118 B.n390 B.n389 10.6151
R1119 B.n391 B.n390 10.6151
R1120 B.n391 B.n208 10.6151
R1121 B.n401 B.n208 10.6151
R1122 B.n402 B.n401 10.6151
R1123 B.n403 B.n402 10.6151
R1124 B.n403 B.n200 10.6151
R1125 B.n413 B.n200 10.6151
R1126 B.n414 B.n413 10.6151
R1127 B.n415 B.n414 10.6151
R1128 B.n415 B.n192 10.6151
R1129 B.n425 B.n192 10.6151
R1130 B.n426 B.n425 10.6151
R1131 B.n427 B.n426 10.6151
R1132 B.n427 B.n184 10.6151
R1133 B.n437 B.n184 10.6151
R1134 B.n438 B.n437 10.6151
R1135 B.n440 B.n438 10.6151
R1136 B.n440 B.n439 10.6151
R1137 B.n439 B.n176 10.6151
R1138 B.n451 B.n176 10.6151
R1139 B.n452 B.n451 10.6151
R1140 B.n453 B.n452 10.6151
R1141 B.n454 B.n453 10.6151
R1142 B.n456 B.n454 10.6151
R1143 B.n457 B.n456 10.6151
R1144 B.n458 B.n457 10.6151
R1145 B.n459 B.n458 10.6151
R1146 B.n461 B.n459 10.6151
R1147 B.n462 B.n461 10.6151
R1148 B.n463 B.n462 10.6151
R1149 B.n464 B.n463 10.6151
R1150 B.n466 B.n464 10.6151
R1151 B.n467 B.n466 10.6151
R1152 B.n468 B.n467 10.6151
R1153 B.n469 B.n468 10.6151
R1154 B.n471 B.n469 10.6151
R1155 B.n472 B.n471 10.6151
R1156 B.n473 B.n472 10.6151
R1157 B.n474 B.n473 10.6151
R1158 B.n476 B.n474 10.6151
R1159 B.n477 B.n476 10.6151
R1160 B.n478 B.n477 10.6151
R1161 B.n479 B.n478 10.6151
R1162 B.n481 B.n479 10.6151
R1163 B.n482 B.n481 10.6151
R1164 B.n483 B.n482 10.6151
R1165 B.n484 B.n483 10.6151
R1166 B.n486 B.n484 10.6151
R1167 B.n487 B.n486 10.6151
R1168 B.n488 B.n487 10.6151
R1169 B.n489 B.n488 10.6151
R1170 B.n491 B.n489 10.6151
R1171 B.n492 B.n491 10.6151
R1172 B.n263 B.n235 10.6151
R1173 B.n263 B.n262 10.6151
R1174 B.n269 B.n262 10.6151
R1175 B.n270 B.n269 10.6151
R1176 B.n271 B.n270 10.6151
R1177 B.n271 B.n260 10.6151
R1178 B.n277 B.n260 10.6151
R1179 B.n278 B.n277 10.6151
R1180 B.n279 B.n278 10.6151
R1181 B.n279 B.n258 10.6151
R1182 B.n285 B.n258 10.6151
R1183 B.n286 B.n285 10.6151
R1184 B.n287 B.n286 10.6151
R1185 B.n287 B.n256 10.6151
R1186 B.n293 B.n256 10.6151
R1187 B.n294 B.n293 10.6151
R1188 B.n298 B.n294 10.6151
R1189 B.n304 B.n254 10.6151
R1190 B.n305 B.n304 10.6151
R1191 B.n306 B.n305 10.6151
R1192 B.n306 B.n252 10.6151
R1193 B.n312 B.n252 10.6151
R1194 B.n313 B.n312 10.6151
R1195 B.n314 B.n313 10.6151
R1196 B.n314 B.n250 10.6151
R1197 B.n321 B.n320 10.6151
R1198 B.n322 B.n321 10.6151
R1199 B.n322 B.n245 10.6151
R1200 B.n328 B.n245 10.6151
R1201 B.n329 B.n328 10.6151
R1202 B.n330 B.n329 10.6151
R1203 B.n330 B.n243 10.6151
R1204 B.n336 B.n243 10.6151
R1205 B.n337 B.n336 10.6151
R1206 B.n338 B.n337 10.6151
R1207 B.n338 B.n241 10.6151
R1208 B.n344 B.n241 10.6151
R1209 B.n345 B.n344 10.6151
R1210 B.n346 B.n345 10.6151
R1211 B.n346 B.n239 10.6151
R1212 B.n352 B.n239 10.6151
R1213 B.n353 B.n352 10.6151
R1214 B.n359 B.n358 10.6151
R1215 B.n360 B.n359 10.6151
R1216 B.n360 B.n227 10.6151
R1217 B.n371 B.n227 10.6151
R1218 B.n372 B.n371 10.6151
R1219 B.n373 B.n372 10.6151
R1220 B.n373 B.n220 10.6151
R1221 B.n383 B.n220 10.6151
R1222 B.n384 B.n383 10.6151
R1223 B.n385 B.n384 10.6151
R1224 B.n385 B.n212 10.6151
R1225 B.n395 B.n212 10.6151
R1226 B.n396 B.n395 10.6151
R1227 B.n397 B.n396 10.6151
R1228 B.n397 B.n204 10.6151
R1229 B.n407 B.n204 10.6151
R1230 B.n408 B.n407 10.6151
R1231 B.n409 B.n408 10.6151
R1232 B.n409 B.n196 10.6151
R1233 B.n419 B.n196 10.6151
R1234 B.n420 B.n419 10.6151
R1235 B.n421 B.n420 10.6151
R1236 B.n421 B.n188 10.6151
R1237 B.n431 B.n188 10.6151
R1238 B.n432 B.n431 10.6151
R1239 B.n433 B.n432 10.6151
R1240 B.n433 B.n180 10.6151
R1241 B.n444 B.n180 10.6151
R1242 B.n445 B.n444 10.6151
R1243 B.n446 B.n445 10.6151
R1244 B.n446 B.n0 10.6151
R1245 B.n556 B.n1 10.6151
R1246 B.n556 B.n555 10.6151
R1247 B.n555 B.n554 10.6151
R1248 B.n554 B.n10 10.6151
R1249 B.n548 B.n10 10.6151
R1250 B.n548 B.n547 10.6151
R1251 B.n547 B.n546 10.6151
R1252 B.n546 B.n17 10.6151
R1253 B.n540 B.n17 10.6151
R1254 B.n540 B.n539 10.6151
R1255 B.n539 B.n538 10.6151
R1256 B.n538 B.n24 10.6151
R1257 B.n532 B.n24 10.6151
R1258 B.n532 B.n531 10.6151
R1259 B.n531 B.n530 10.6151
R1260 B.n530 B.n31 10.6151
R1261 B.n524 B.n31 10.6151
R1262 B.n524 B.n523 10.6151
R1263 B.n523 B.n522 10.6151
R1264 B.n522 B.n38 10.6151
R1265 B.n516 B.n38 10.6151
R1266 B.n516 B.n515 10.6151
R1267 B.n515 B.n514 10.6151
R1268 B.n514 B.n45 10.6151
R1269 B.n508 B.n45 10.6151
R1270 B.n508 B.n507 10.6151
R1271 B.n507 B.n506 10.6151
R1272 B.n506 B.n51 10.6151
R1273 B.n500 B.n51 10.6151
R1274 B.n500 B.n499 10.6151
R1275 B.n499 B.n498 10.6151
R1276 B.n125 B.n89 6.5566
R1277 B.n142 B.n141 6.5566
R1278 B.n297 B.n254 6.5566
R1279 B.n250 B.n249 6.5566
R1280 B.n122 B.n89 4.05904
R1281 B.n143 B.n142 4.05904
R1282 B.n298 B.n297 4.05904
R1283 B.n320 B.n249 4.05904
R1284 B.n562 B.n0 2.81026
R1285 B.n562 B.n1 2.81026
R1286 VN.n37 VN.n20 161.3
R1287 VN.n35 VN.n34 161.3
R1288 VN.n33 VN.n21 161.3
R1289 VN.n32 VN.n31 161.3
R1290 VN.n29 VN.n22 161.3
R1291 VN.n28 VN.n27 161.3
R1292 VN.n26 VN.n23 161.3
R1293 VN.n17 VN.n0 161.3
R1294 VN.n15 VN.n14 161.3
R1295 VN.n13 VN.n1 161.3
R1296 VN.n12 VN.n11 161.3
R1297 VN.n9 VN.n2 161.3
R1298 VN.n8 VN.n7 161.3
R1299 VN.n6 VN.n3 161.3
R1300 VN.n5 VN.t6 143.904
R1301 VN.n25 VN.t5 143.904
R1302 VN.n18 VN.t1 129.243
R1303 VN.n38 VN.t7 129.243
R1304 VN.n4 VN.t2 90.7299
R1305 VN.n10 VN.t4 90.7299
R1306 VN.n16 VN.t8 90.7299
R1307 VN.n24 VN.t3 90.7299
R1308 VN.n30 VN.t0 90.7299
R1309 VN.n36 VN.t9 90.7299
R1310 VN.n39 VN.n38 80.6037
R1311 VN.n19 VN.n18 80.6037
R1312 VN.n18 VN.n17 53.6107
R1313 VN.n38 VN.n37 53.6107
R1314 VN.n5 VN.n4 48.9084
R1315 VN.n25 VN.n24 48.9084
R1316 VN.n9 VN.n8 47.8428
R1317 VN.n11 VN.n1 47.8428
R1318 VN.n29 VN.n28 47.8428
R1319 VN.n31 VN.n21 47.8428
R1320 VN.n26 VN.n25 44.2988
R1321 VN.n6 VN.n5 44.2988
R1322 VN VN.n39 38.8134
R1323 VN.n8 VN.n3 33.3113
R1324 VN.n15 VN.n1 33.3113
R1325 VN.n28 VN.n23 33.3113
R1326 VN.n35 VN.n21 33.3113
R1327 VN.n17 VN.n16 19.674
R1328 VN.n37 VN.n36 19.674
R1329 VN.n10 VN.n9 12.2964
R1330 VN.n11 VN.n10 12.2964
R1331 VN.n31 VN.n30 12.2964
R1332 VN.n30 VN.n29 12.2964
R1333 VN.n4 VN.n3 4.91887
R1334 VN.n16 VN.n15 4.91887
R1335 VN.n24 VN.n23 4.91887
R1336 VN.n36 VN.n35 4.91887
R1337 VN.n39 VN.n20 0.285035
R1338 VN.n19 VN.n0 0.285035
R1339 VN.n34 VN.n20 0.189894
R1340 VN.n34 VN.n33 0.189894
R1341 VN.n33 VN.n32 0.189894
R1342 VN.n32 VN.n22 0.189894
R1343 VN.n27 VN.n22 0.189894
R1344 VN.n27 VN.n26 0.189894
R1345 VN.n7 VN.n6 0.189894
R1346 VN.n7 VN.n2 0.189894
R1347 VN.n12 VN.n2 0.189894
R1348 VN.n13 VN.n12 0.189894
R1349 VN.n14 VN.n13 0.189894
R1350 VN.n14 VN.n0 0.189894
R1351 VN VN.n19 0.146778
R1352 VDD2.n37 VDD2.n23 289.615
R1353 VDD2.n14 VDD2.n0 289.615
R1354 VDD2.n38 VDD2.n37 185
R1355 VDD2.n36 VDD2.n35 185
R1356 VDD2.n27 VDD2.n26 185
R1357 VDD2.n30 VDD2.n29 185
R1358 VDD2.n7 VDD2.n6 185
R1359 VDD2.n4 VDD2.n3 185
R1360 VDD2.n13 VDD2.n12 185
R1361 VDD2.n15 VDD2.n14 185
R1362 VDD2.t2 VDD2.n28 147.888
R1363 VDD2.t3 VDD2.n5 147.888
R1364 VDD2.n37 VDD2.n36 104.615
R1365 VDD2.n36 VDD2.n26 104.615
R1366 VDD2.n29 VDD2.n26 104.615
R1367 VDD2.n6 VDD2.n3 104.615
R1368 VDD2.n13 VDD2.n3 104.615
R1369 VDD2.n14 VDD2.n13 104.615
R1370 VDD2.n22 VDD2.n21 74.2815
R1371 VDD2 VDD2.n45 74.2786
R1372 VDD2.n44 VDD2.n43 73.4641
R1373 VDD2.n20 VDD2.n19 73.464
R1374 VDD2.n29 VDD2.t2 52.3082
R1375 VDD2.n6 VDD2.t3 52.3082
R1376 VDD2.n20 VDD2.n18 50.0279
R1377 VDD2.n42 VDD2.n41 48.8641
R1378 VDD2.n42 VDD2.n22 32.5537
R1379 VDD2.n30 VDD2.n28 15.6496
R1380 VDD2.n7 VDD2.n5 15.6496
R1381 VDD2.n31 VDD2.n27 12.8005
R1382 VDD2.n8 VDD2.n4 12.8005
R1383 VDD2.n35 VDD2.n34 12.0247
R1384 VDD2.n12 VDD2.n11 12.0247
R1385 VDD2.n38 VDD2.n25 11.249
R1386 VDD2.n15 VDD2.n2 11.249
R1387 VDD2.n39 VDD2.n23 10.4732
R1388 VDD2.n16 VDD2.n0 10.4732
R1389 VDD2.n41 VDD2.n40 9.45567
R1390 VDD2.n18 VDD2.n17 9.45567
R1391 VDD2.n40 VDD2.n39 9.3005
R1392 VDD2.n25 VDD2.n24 9.3005
R1393 VDD2.n34 VDD2.n33 9.3005
R1394 VDD2.n32 VDD2.n31 9.3005
R1395 VDD2.n17 VDD2.n16 9.3005
R1396 VDD2.n2 VDD2.n1 9.3005
R1397 VDD2.n11 VDD2.n10 9.3005
R1398 VDD2.n9 VDD2.n8 9.3005
R1399 VDD2.n45 VDD2.t6 5.15675
R1400 VDD2.n45 VDD2.t4 5.15675
R1401 VDD2.n43 VDD2.t0 5.15675
R1402 VDD2.n43 VDD2.t9 5.15675
R1403 VDD2.n21 VDD2.t1 5.15675
R1404 VDD2.n21 VDD2.t8 5.15675
R1405 VDD2.n19 VDD2.t7 5.15675
R1406 VDD2.n19 VDD2.t5 5.15675
R1407 VDD2.n32 VDD2.n28 4.40546
R1408 VDD2.n9 VDD2.n5 4.40546
R1409 VDD2.n41 VDD2.n23 3.49141
R1410 VDD2.n18 VDD2.n0 3.49141
R1411 VDD2.n39 VDD2.n38 2.71565
R1412 VDD2.n16 VDD2.n15 2.71565
R1413 VDD2.n35 VDD2.n25 1.93989
R1414 VDD2.n12 VDD2.n2 1.93989
R1415 VDD2.n44 VDD2.n42 1.16429
R1416 VDD2.n34 VDD2.n27 1.16414
R1417 VDD2.n11 VDD2.n4 1.16414
R1418 VDD2.n31 VDD2.n30 0.388379
R1419 VDD2.n8 VDD2.n7 0.388379
R1420 VDD2 VDD2.n44 0.349638
R1421 VDD2.n22 VDD2.n20 0.236102
R1422 VDD2.n40 VDD2.n24 0.155672
R1423 VDD2.n33 VDD2.n24 0.155672
R1424 VDD2.n33 VDD2.n32 0.155672
R1425 VDD2.n10 VDD2.n9 0.155672
R1426 VDD2.n10 VDD2.n1 0.155672
R1427 VDD2.n17 VDD2.n1 0.155672
C0 VDD1 VP 3.10375f
C1 VN VTAIL 3.29132f
C2 VDD1 VDD2 1.17185f
C3 VDD1 VN 0.154469f
C4 VP VDD2 0.386358f
C5 VDD1 VTAIL 5.884931f
C6 VP VN 4.55907f
C7 VP VTAIL 3.30556f
C8 VDD2 VN 2.87431f
C9 VDD2 VTAIL 5.92618f
C10 VDD2 B 3.873999f
C11 VDD1 B 3.828153f
C12 VTAIL B 3.57575f
C13 VN B 9.913189f
C14 VP B 8.351677f
C15 VDD2.n0 B 0.031279f
C16 VDD2.n1 B 0.023613f
C17 VDD2.n2 B 0.012689f
C18 VDD2.n3 B 0.029991f
C19 VDD2.n4 B 0.013435f
C20 VDD2.n5 B 0.089609f
C21 VDD2.t3 B 0.049521f
C22 VDD2.n6 B 0.022494f
C23 VDD2.n7 B 0.017652f
C24 VDD2.n8 B 0.012689f
C25 VDD2.n9 B 0.325999f
C26 VDD2.n10 B 0.023613f
C27 VDD2.n11 B 0.012689f
C28 VDD2.n12 B 0.013435f
C29 VDD2.n13 B 0.029991f
C30 VDD2.n14 B 0.061545f
C31 VDD2.n15 B 0.013435f
C32 VDD2.n16 B 0.012689f
C33 VDD2.n17 B 0.054581f
C34 VDD2.n18 B 0.053512f
C35 VDD2.t7 B 0.071654f
C36 VDD2.t5 B 0.071654f
C37 VDD2.n19 B 0.55959f
C38 VDD2.n20 B 0.42199f
C39 VDD2.t1 B 0.071654f
C40 VDD2.t8 B 0.071654f
C41 VDD2.n21 B 0.563367f
C42 VDD2.n22 B 1.49115f
C43 VDD2.n23 B 0.031279f
C44 VDD2.n24 B 0.023613f
C45 VDD2.n25 B 0.012689f
C46 VDD2.n26 B 0.029991f
C47 VDD2.n27 B 0.013435f
C48 VDD2.n28 B 0.089609f
C49 VDD2.t2 B 0.049521f
C50 VDD2.n29 B 0.022494f
C51 VDD2.n30 B 0.017652f
C52 VDD2.n31 B 0.012689f
C53 VDD2.n32 B 0.325999f
C54 VDD2.n33 B 0.023613f
C55 VDD2.n34 B 0.012689f
C56 VDD2.n35 B 0.013435f
C57 VDD2.n36 B 0.029991f
C58 VDD2.n37 B 0.061545f
C59 VDD2.n38 B 0.013435f
C60 VDD2.n39 B 0.012689f
C61 VDD2.n40 B 0.054581f
C62 VDD2.n41 B 0.050394f
C63 VDD2.n42 B 1.53741f
C64 VDD2.t0 B 0.071654f
C65 VDD2.t9 B 0.071654f
C66 VDD2.n43 B 0.559593f
C67 VDD2.n44 B 0.297402f
C68 VDD2.t6 B 0.071654f
C69 VDD2.t4 B 0.071654f
C70 VDD2.n45 B 0.563345f
C71 VN.n0 B 0.05271f
C72 VN.t8 B 0.395956f
C73 VN.n1 B 0.03483f
C74 VN.n2 B 0.039501f
C75 VN.t4 B 0.395956f
C76 VN.n3 B 0.050379f
C77 VN.t6 B 0.482012f
C78 VN.t2 B 0.395956f
C79 VN.n4 B 0.211891f
C80 VN.n5 B 0.239334f
C81 VN.n6 B 0.167417f
C82 VN.n7 B 0.039501f
C83 VN.n8 B 0.03483f
C84 VN.n9 B 0.055873f
C85 VN.n10 B 0.180694f
C86 VN.n11 B 0.055873f
C87 VN.n12 B 0.039501f
C88 VN.n13 B 0.039501f
C89 VN.n14 B 0.039501f
C90 VN.n15 B 0.050379f
C91 VN.n16 B 0.180694f
C92 VN.n17 B 0.052191f
C93 VN.t1 B 0.457307f
C94 VN.n18 B 0.242228f
C95 VN.n19 B 0.036995f
C96 VN.n20 B 0.05271f
C97 VN.t9 B 0.395956f
C98 VN.n21 B 0.03483f
C99 VN.n22 B 0.039501f
C100 VN.t0 B 0.395956f
C101 VN.n23 B 0.050379f
C102 VN.t5 B 0.482012f
C103 VN.t3 B 0.395956f
C104 VN.n24 B 0.211891f
C105 VN.n25 B 0.239334f
C106 VN.n26 B 0.167417f
C107 VN.n27 B 0.039501f
C108 VN.n28 B 0.03483f
C109 VN.n29 B 0.055873f
C110 VN.n30 B 0.180694f
C111 VN.n31 B 0.055873f
C112 VN.n32 B 0.039501f
C113 VN.n33 B 0.039501f
C114 VN.n34 B 0.039501f
C115 VN.n35 B 0.050379f
C116 VN.n36 B 0.180694f
C117 VN.n37 B 0.052191f
C118 VN.t7 B 0.457307f
C119 VN.n38 B 0.242228f
C120 VN.n39 B 1.44225f
C121 VTAIL.t1 B 0.08787f
C122 VTAIL.t19 B 0.08787f
C123 VTAIL.n0 B 0.622195f
C124 VTAIL.n1 B 0.433233f
C125 VTAIL.n2 B 0.038357f
C126 VTAIL.n3 B 0.028957f
C127 VTAIL.n4 B 0.01556f
C128 VTAIL.n5 B 0.036779f
C129 VTAIL.n6 B 0.016476f
C130 VTAIL.n7 B 0.109889f
C131 VTAIL.t9 B 0.060728f
C132 VTAIL.n8 B 0.027584f
C133 VTAIL.n9 B 0.021647f
C134 VTAIL.n10 B 0.01556f
C135 VTAIL.n11 B 0.399778f
C136 VTAIL.n12 B 0.028957f
C137 VTAIL.n13 B 0.01556f
C138 VTAIL.n14 B 0.016476f
C139 VTAIL.n15 B 0.036779f
C140 VTAIL.n16 B 0.075475f
C141 VTAIL.n17 B 0.016476f
C142 VTAIL.n18 B 0.01556f
C143 VTAIL.n19 B 0.066933f
C144 VTAIL.n20 B 0.041805f
C145 VTAIL.n21 B 0.231454f
C146 VTAIL.t13 B 0.08787f
C147 VTAIL.t15 B 0.08787f
C148 VTAIL.n22 B 0.622195f
C149 VTAIL.n23 B 0.465407f
C150 VTAIL.t16 B 0.08787f
C151 VTAIL.t18 B 0.08787f
C152 VTAIL.n24 B 0.622195f
C153 VTAIL.n25 B 1.27622f
C154 VTAIL.t8 B 0.08787f
C155 VTAIL.t5 B 0.08787f
C156 VTAIL.n26 B 0.6222f
C157 VTAIL.n27 B 1.27622f
C158 VTAIL.t7 B 0.08787f
C159 VTAIL.t4 B 0.08787f
C160 VTAIL.n28 B 0.6222f
C161 VTAIL.n29 B 0.465403f
C162 VTAIL.n30 B 0.038357f
C163 VTAIL.n31 B 0.028957f
C164 VTAIL.n32 B 0.01556f
C165 VTAIL.n33 B 0.036779f
C166 VTAIL.n34 B 0.016476f
C167 VTAIL.n35 B 0.109889f
C168 VTAIL.t0 B 0.060728f
C169 VTAIL.n36 B 0.027584f
C170 VTAIL.n37 B 0.021647f
C171 VTAIL.n38 B 0.01556f
C172 VTAIL.n39 B 0.399778f
C173 VTAIL.n40 B 0.028957f
C174 VTAIL.n41 B 0.01556f
C175 VTAIL.n42 B 0.016476f
C176 VTAIL.n43 B 0.036779f
C177 VTAIL.n44 B 0.075475f
C178 VTAIL.n45 B 0.016476f
C179 VTAIL.n46 B 0.01556f
C180 VTAIL.n47 B 0.066933f
C181 VTAIL.n48 B 0.041805f
C182 VTAIL.n49 B 0.231454f
C183 VTAIL.t12 B 0.08787f
C184 VTAIL.t14 B 0.08787f
C185 VTAIL.n50 B 0.6222f
C186 VTAIL.n51 B 0.454946f
C187 VTAIL.t17 B 0.08787f
C188 VTAIL.t10 B 0.08787f
C189 VTAIL.n52 B 0.6222f
C190 VTAIL.n53 B 0.465403f
C191 VTAIL.n54 B 0.038357f
C192 VTAIL.n55 B 0.028957f
C193 VTAIL.n56 B 0.01556f
C194 VTAIL.n57 B 0.036779f
C195 VTAIL.n58 B 0.016476f
C196 VTAIL.n59 B 0.109889f
C197 VTAIL.t11 B 0.060728f
C198 VTAIL.n60 B 0.027584f
C199 VTAIL.n61 B 0.021647f
C200 VTAIL.n62 B 0.01556f
C201 VTAIL.n63 B 0.399778f
C202 VTAIL.n64 B 0.028957f
C203 VTAIL.n65 B 0.01556f
C204 VTAIL.n66 B 0.016476f
C205 VTAIL.n67 B 0.036779f
C206 VTAIL.n68 B 0.075475f
C207 VTAIL.n69 B 0.016476f
C208 VTAIL.n70 B 0.01556f
C209 VTAIL.n71 B 0.066933f
C210 VTAIL.n72 B 0.041805f
C211 VTAIL.n73 B 0.944138f
C212 VTAIL.n74 B 0.038357f
C213 VTAIL.n75 B 0.028957f
C214 VTAIL.n76 B 0.01556f
C215 VTAIL.n77 B 0.036779f
C216 VTAIL.n78 B 0.016476f
C217 VTAIL.n79 B 0.109889f
C218 VTAIL.t3 B 0.060728f
C219 VTAIL.n80 B 0.027584f
C220 VTAIL.n81 B 0.021647f
C221 VTAIL.n82 B 0.01556f
C222 VTAIL.n83 B 0.399778f
C223 VTAIL.n84 B 0.028957f
C224 VTAIL.n85 B 0.01556f
C225 VTAIL.n86 B 0.016476f
C226 VTAIL.n87 B 0.036779f
C227 VTAIL.n88 B 0.075475f
C228 VTAIL.n89 B 0.016476f
C229 VTAIL.n90 B 0.01556f
C230 VTAIL.n91 B 0.066933f
C231 VTAIL.n92 B 0.041805f
C232 VTAIL.n93 B 0.944138f
C233 VTAIL.t2 B 0.08787f
C234 VTAIL.t6 B 0.08787f
C235 VTAIL.n94 B 0.622195f
C236 VTAIL.n95 B 0.378536f
C237 VDD1.n0 B 0.031676f
C238 VDD1.n1 B 0.023913f
C239 VDD1.n2 B 0.01285f
C240 VDD1.n3 B 0.030372f
C241 VDD1.n4 B 0.013606f
C242 VDD1.n5 B 0.090746f
C243 VDD1.t0 B 0.050149f
C244 VDD1.n6 B 0.022779f
C245 VDD1.n7 B 0.017876f
C246 VDD1.n8 B 0.01285f
C247 VDD1.n9 B 0.330136f
C248 VDD1.n10 B 0.023913f
C249 VDD1.n11 B 0.01285f
C250 VDD1.n12 B 0.013606f
C251 VDD1.n13 B 0.030372f
C252 VDD1.n14 B 0.062327f
C253 VDD1.n15 B 0.013606f
C254 VDD1.n16 B 0.01285f
C255 VDD1.n17 B 0.055273f
C256 VDD1.n18 B 0.054191f
C257 VDD1.t5 B 0.072563f
C258 VDD1.t4 B 0.072563f
C259 VDD1.n19 B 0.566694f
C260 VDD1.n20 B 0.433737f
C261 VDD1.n21 B 0.031676f
C262 VDD1.n22 B 0.023913f
C263 VDD1.n23 B 0.01285f
C264 VDD1.n24 B 0.030372f
C265 VDD1.n25 B 0.013606f
C266 VDD1.n26 B 0.090746f
C267 VDD1.t6 B 0.050149f
C268 VDD1.n27 B 0.022779f
C269 VDD1.n28 B 0.017876f
C270 VDD1.n29 B 0.01285f
C271 VDD1.n30 B 0.330136f
C272 VDD1.n31 B 0.023913f
C273 VDD1.n32 B 0.01285f
C274 VDD1.n33 B 0.013606f
C275 VDD1.n34 B 0.030372f
C276 VDD1.n35 B 0.062327f
C277 VDD1.n36 B 0.013606f
C278 VDD1.n37 B 0.01285f
C279 VDD1.n38 B 0.055273f
C280 VDD1.n39 B 0.054191f
C281 VDD1.t9 B 0.072563f
C282 VDD1.t8 B 0.072563f
C283 VDD1.n40 B 0.566692f
C284 VDD1.n41 B 0.427345f
C285 VDD1.t7 B 0.072563f
C286 VDD1.t1 B 0.072563f
C287 VDD1.n42 B 0.570517f
C288 VDD1.n43 B 1.58672f
C289 VDD1.t2 B 0.072563f
C290 VDD1.t3 B 0.072563f
C291 VDD1.n44 B 0.566692f
C292 VDD1.n45 B 1.77955f
C293 VP.n0 B 0.053963f
C294 VP.t3 B 0.405373f
C295 VP.n1 B 0.035659f
C296 VP.n2 B 0.040441f
C297 VP.t5 B 0.405373f
C298 VP.n3 B 0.051578f
C299 VP.n4 B 0.053963f
C300 VP.t7 B 0.468183f
C301 VP.t8 B 0.405373f
C302 VP.n5 B 0.035659f
C303 VP.n6 B 0.040441f
C304 VP.t1 B 0.405373f
C305 VP.n7 B 0.051578f
C306 VP.t4 B 0.405373f
C307 VP.n8 B 0.21693f
C308 VP.t6 B 0.493475f
C309 VP.n9 B 0.245025f
C310 VP.n10 B 0.171399f
C311 VP.n11 B 0.040441f
C312 VP.n12 B 0.035659f
C313 VP.n13 B 0.057202f
C314 VP.n14 B 0.184991f
C315 VP.n15 B 0.057202f
C316 VP.n16 B 0.040441f
C317 VP.n17 B 0.040441f
C318 VP.n18 B 0.040441f
C319 VP.n19 B 0.051578f
C320 VP.n20 B 0.184991f
C321 VP.n21 B 0.053432f
C322 VP.n22 B 0.247989f
C323 VP.n23 B 1.4535f
C324 VP.n24 B 1.49134f
C325 VP.t2 B 0.468183f
C326 VP.n25 B 0.247989f
C327 VP.t0 B 0.405373f
C328 VP.n26 B 0.184991f
C329 VP.n27 B 0.053432f
C330 VP.n28 B 0.053963f
C331 VP.n29 B 0.040441f
C332 VP.n30 B 0.040441f
C333 VP.n31 B 0.035659f
C334 VP.n32 B 0.057202f
C335 VP.n33 B 0.184991f
C336 VP.n34 B 0.057202f
C337 VP.n35 B 0.040441f
C338 VP.n36 B 0.040441f
C339 VP.n37 B 0.040441f
C340 VP.n38 B 0.051578f
C341 VP.n39 B 0.184991f
C342 VP.n40 B 0.053432f
C343 VP.t9 B 0.468183f
C344 VP.n41 B 0.247989f
C345 VP.n42 B 0.037874f
.ends

