* NGSPICE file created from diff_pair_sample_0805.ext - technology: sky130A

.subckt diff_pair_sample_0805 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t7 B.t21 sky130_fd_pr__nfet_01v8 ad=0.13035 pd=1.12 as=0.3081 ps=2.36 w=0.79 l=3.56
X1 VDD2.t7 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.13035 pd=1.12 as=0.13035 ps=1.12 w=0.79 l=3.56
X2 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=0.3081 pd=2.36 as=0 ps=0 w=0.79 l=3.56
X3 VDD1.t6 VP.t1 VTAIL.t4 B.t20 sky130_fd_pr__nfet_01v8 ad=0.13035 pd=1.12 as=0.3081 ps=2.36 w=0.79 l=3.56
X4 VDD1.t5 VP.t2 VTAIL.t6 B.t19 sky130_fd_pr__nfet_01v8 ad=0.13035 pd=1.12 as=0.13035 ps=1.12 w=0.79 l=3.56
X5 VTAIL.t0 VN.t1 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.13035 pd=1.12 as=0.13035 ps=1.12 w=0.79 l=3.56
X6 VTAIL.t3 VP.t3 VDD1.t4 B.t18 sky130_fd_pr__nfet_01v8 ad=0.13035 pd=1.12 as=0.13035 ps=1.12 w=0.79 l=3.56
X7 VTAIL.t13 VN.t2 VDD2.t5 B.t18 sky130_fd_pr__nfet_01v8 ad=0.13035 pd=1.12 as=0.13035 ps=1.12 w=0.79 l=3.56
X8 VDD1.t3 VP.t4 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.13035 pd=1.12 as=0.13035 ps=1.12 w=0.79 l=3.56
X9 VTAIL.t2 VP.t5 VDD1.t2 B.t17 sky130_fd_pr__nfet_01v8 ad=0.3081 pd=2.36 as=0.13035 ps=1.12 w=0.79 l=3.56
X10 VTAIL.t15 VN.t3 VDD2.t4 B.t16 sky130_fd_pr__nfet_01v8 ad=0.3081 pd=2.36 as=0.13035 ps=1.12 w=0.79 l=3.56
X11 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=0.3081 pd=2.36 as=0 ps=0 w=0.79 l=3.56
X12 VDD2.t3 VN.t4 VTAIL.t14 B.t20 sky130_fd_pr__nfet_01v8 ad=0.13035 pd=1.12 as=0.3081 ps=2.36 w=0.79 l=3.56
X13 VTAIL.t12 VN.t5 VDD2.t2 B.t17 sky130_fd_pr__nfet_01v8 ad=0.3081 pd=2.36 as=0.13035 ps=1.12 w=0.79 l=3.56
X14 VTAIL.t9 VP.t6 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.13035 pd=1.12 as=0.13035 ps=1.12 w=0.79 l=3.56
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.3081 pd=2.36 as=0 ps=0 w=0.79 l=3.56
X16 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.3081 pd=2.36 as=0 ps=0 w=0.79 l=3.56
X17 VTAIL.t8 VP.t7 VDD1.t0 B.t16 sky130_fd_pr__nfet_01v8 ad=0.3081 pd=2.36 as=0.13035 ps=1.12 w=0.79 l=3.56
X18 VDD2.t1 VN.t6 VTAIL.t11 B.t21 sky130_fd_pr__nfet_01v8 ad=0.13035 pd=1.12 as=0.3081 ps=2.36 w=0.79 l=3.56
X19 VDD2.t0 VN.t7 VTAIL.t10 B.t19 sky130_fd_pr__nfet_01v8 ad=0.13035 pd=1.12 as=0.13035 ps=1.12 w=0.79 l=3.56
R0 VP.n24 VP.n21 161.3
R1 VP.n26 VP.n25 161.3
R2 VP.n27 VP.n20 161.3
R3 VP.n29 VP.n28 161.3
R4 VP.n30 VP.n19 161.3
R5 VP.n32 VP.n31 161.3
R6 VP.n33 VP.n18 161.3
R7 VP.n36 VP.n35 161.3
R8 VP.n37 VP.n17 161.3
R9 VP.n39 VP.n38 161.3
R10 VP.n40 VP.n16 161.3
R11 VP.n42 VP.n41 161.3
R12 VP.n43 VP.n15 161.3
R13 VP.n45 VP.n44 161.3
R14 VP.n46 VP.n14 161.3
R15 VP.n48 VP.n47 161.3
R16 VP.n89 VP.n88 161.3
R17 VP.n87 VP.n1 161.3
R18 VP.n86 VP.n85 161.3
R19 VP.n84 VP.n2 161.3
R20 VP.n83 VP.n82 161.3
R21 VP.n81 VP.n3 161.3
R22 VP.n80 VP.n79 161.3
R23 VP.n78 VP.n4 161.3
R24 VP.n77 VP.n76 161.3
R25 VP.n74 VP.n5 161.3
R26 VP.n73 VP.n72 161.3
R27 VP.n71 VP.n6 161.3
R28 VP.n70 VP.n69 161.3
R29 VP.n68 VP.n7 161.3
R30 VP.n67 VP.n66 161.3
R31 VP.n65 VP.n8 161.3
R32 VP.n64 VP.n63 161.3
R33 VP.n61 VP.n9 161.3
R34 VP.n60 VP.n59 161.3
R35 VP.n58 VP.n10 161.3
R36 VP.n57 VP.n56 161.3
R37 VP.n55 VP.n11 161.3
R38 VP.n54 VP.n53 161.3
R39 VP.n52 VP.n12 161.3
R40 VP.n51 VP.n50 85.908
R41 VP.n90 VP.n0 85.908
R42 VP.n49 VP.n13 85.908
R43 VP.n23 VP.n22 65.0012
R44 VP.n69 VP.n6 56.5193
R45 VP.n28 VP.n19 56.5193
R46 VP.n56 VP.n10 54.0911
R47 VP.n82 VP.n2 54.0911
R48 VP.n41 VP.n15 54.0911
R49 VP.n51 VP.n49 46.9084
R50 VP.n23 VP.t5 37.5795
R51 VP.n60 VP.n10 26.8957
R52 VP.n82 VP.n81 26.8957
R53 VP.n41 VP.n40 26.8957
R54 VP.n54 VP.n12 24.4675
R55 VP.n55 VP.n54 24.4675
R56 VP.n56 VP.n55 24.4675
R57 VP.n61 VP.n60 24.4675
R58 VP.n63 VP.n61 24.4675
R59 VP.n67 VP.n8 24.4675
R60 VP.n68 VP.n67 24.4675
R61 VP.n69 VP.n68 24.4675
R62 VP.n73 VP.n6 24.4675
R63 VP.n74 VP.n73 24.4675
R64 VP.n76 VP.n74 24.4675
R65 VP.n80 VP.n4 24.4675
R66 VP.n81 VP.n80 24.4675
R67 VP.n86 VP.n2 24.4675
R68 VP.n87 VP.n86 24.4675
R69 VP.n88 VP.n87 24.4675
R70 VP.n45 VP.n15 24.4675
R71 VP.n46 VP.n45 24.4675
R72 VP.n47 VP.n46 24.4675
R73 VP.n32 VP.n19 24.4675
R74 VP.n33 VP.n32 24.4675
R75 VP.n35 VP.n33 24.4675
R76 VP.n39 VP.n17 24.4675
R77 VP.n40 VP.n39 24.4675
R78 VP.n26 VP.n21 24.4675
R79 VP.n27 VP.n26 24.4675
R80 VP.n28 VP.n27 24.4675
R81 VP.n63 VP.n62 14.9254
R82 VP.n75 VP.n4 14.9254
R83 VP.n34 VP.n17 14.9254
R84 VP.n62 VP.n8 9.54263
R85 VP.n76 VP.n75 9.54263
R86 VP.n35 VP.n34 9.54263
R87 VP.n22 VP.n21 9.54263
R88 VP.n50 VP.t7 5.34853
R89 VP.n62 VP.t4 5.34853
R90 VP.n75 VP.t3 5.34853
R91 VP.n0 VP.t1 5.34853
R92 VP.n13 VP.t0 5.34853
R93 VP.n34 VP.t6 5.34853
R94 VP.n22 VP.t2 5.34853
R95 VP.n50 VP.n12 4.15989
R96 VP.n88 VP.n0 4.15989
R97 VP.n47 VP.n13 4.15989
R98 VP.n24 VP.n23 3.34372
R99 VP.n49 VP.n48 0.354971
R100 VP.n52 VP.n51 0.354971
R101 VP.n90 VP.n89 0.354971
R102 VP VP.n90 0.26696
R103 VP.n25 VP.n24 0.189894
R104 VP.n25 VP.n20 0.189894
R105 VP.n29 VP.n20 0.189894
R106 VP.n30 VP.n29 0.189894
R107 VP.n31 VP.n30 0.189894
R108 VP.n31 VP.n18 0.189894
R109 VP.n36 VP.n18 0.189894
R110 VP.n37 VP.n36 0.189894
R111 VP.n38 VP.n37 0.189894
R112 VP.n38 VP.n16 0.189894
R113 VP.n42 VP.n16 0.189894
R114 VP.n43 VP.n42 0.189894
R115 VP.n44 VP.n43 0.189894
R116 VP.n44 VP.n14 0.189894
R117 VP.n48 VP.n14 0.189894
R118 VP.n53 VP.n52 0.189894
R119 VP.n53 VP.n11 0.189894
R120 VP.n57 VP.n11 0.189894
R121 VP.n58 VP.n57 0.189894
R122 VP.n59 VP.n58 0.189894
R123 VP.n59 VP.n9 0.189894
R124 VP.n64 VP.n9 0.189894
R125 VP.n65 VP.n64 0.189894
R126 VP.n66 VP.n65 0.189894
R127 VP.n66 VP.n7 0.189894
R128 VP.n70 VP.n7 0.189894
R129 VP.n71 VP.n70 0.189894
R130 VP.n72 VP.n71 0.189894
R131 VP.n72 VP.n5 0.189894
R132 VP.n77 VP.n5 0.189894
R133 VP.n78 VP.n77 0.189894
R134 VP.n79 VP.n78 0.189894
R135 VP.n79 VP.n3 0.189894
R136 VP.n83 VP.n3 0.189894
R137 VP.n84 VP.n83 0.189894
R138 VP.n85 VP.n84 0.189894
R139 VP.n85 VP.n1 0.189894
R140 VP.n89 VP.n1 0.189894
R141 VTAIL.n15 VTAIL.t11 245.934
R142 VTAIL.n2 VTAIL.t12 245.934
R143 VTAIL.n3 VTAIL.t4 245.934
R144 VTAIL.n6 VTAIL.t8 245.934
R145 VTAIL.n14 VTAIL.t7 245.934
R146 VTAIL.n11 VTAIL.t2 245.934
R147 VTAIL.n10 VTAIL.t14 245.934
R148 VTAIL.n7 VTAIL.t15 245.934
R149 VTAIL.n1 VTAIL.n0 220.87
R150 VTAIL.n5 VTAIL.n4 220.87
R151 VTAIL.n13 VTAIL.n12 220.87
R152 VTAIL.n9 VTAIL.n8 220.87
R153 VTAIL.n0 VTAIL.t10 25.0638
R154 VTAIL.n0 VTAIL.t0 25.0638
R155 VTAIL.n4 VTAIL.t5 25.0638
R156 VTAIL.n4 VTAIL.t3 25.0638
R157 VTAIL.n12 VTAIL.t6 25.0638
R158 VTAIL.n12 VTAIL.t9 25.0638
R159 VTAIL.n8 VTAIL.t1 25.0638
R160 VTAIL.n8 VTAIL.t13 25.0638
R161 VTAIL.n15 VTAIL.n14 16.4014
R162 VTAIL.n7 VTAIL.n6 16.4014
R163 VTAIL.n9 VTAIL.n7 3.35395
R164 VTAIL.n10 VTAIL.n9 3.35395
R165 VTAIL.n13 VTAIL.n11 3.35395
R166 VTAIL.n14 VTAIL.n13 3.35395
R167 VTAIL.n6 VTAIL.n5 3.35395
R168 VTAIL.n5 VTAIL.n3 3.35395
R169 VTAIL.n2 VTAIL.n1 3.35395
R170 VTAIL VTAIL.n15 3.29576
R171 VTAIL.n11 VTAIL.n10 0.470328
R172 VTAIL.n3 VTAIL.n2 0.470328
R173 VTAIL VTAIL.n1 0.0586897
R174 VDD1 VDD1.n0 239.284
R175 VDD1.n3 VDD1.n2 239.171
R176 VDD1.n3 VDD1.n1 239.171
R177 VDD1.n5 VDD1.n4 237.548
R178 VDD1.n5 VDD1.n3 40.0699
R179 VDD1.n4 VDD1.t1 25.0638
R180 VDD1.n4 VDD1.t7 25.0638
R181 VDD1.n0 VDD1.t2 25.0638
R182 VDD1.n0 VDD1.t5 25.0638
R183 VDD1.n2 VDD1.t4 25.0638
R184 VDD1.n2 VDD1.t6 25.0638
R185 VDD1.n1 VDD1.t0 25.0638
R186 VDD1.n1 VDD1.t3 25.0638
R187 VDD1 VDD1.n5 1.61903
R188 B.n672 B.n671 585
R189 B.n673 B.n672 585
R190 B.n190 B.n133 585
R191 B.n189 B.n188 585
R192 B.n187 B.n186 585
R193 B.n185 B.n184 585
R194 B.n183 B.n182 585
R195 B.n181 B.n180 585
R196 B.n179 B.n178 585
R197 B.n177 B.n176 585
R198 B.n175 B.n174 585
R199 B.n173 B.n172 585
R200 B.n171 B.n170 585
R201 B.n169 B.n168 585
R202 B.n167 B.n166 585
R203 B.n165 B.n164 585
R204 B.n163 B.n162 585
R205 B.n161 B.n160 585
R206 B.n159 B.n158 585
R207 B.n156 B.n155 585
R208 B.n154 B.n153 585
R209 B.n152 B.n151 585
R210 B.n150 B.n149 585
R211 B.n148 B.n147 585
R212 B.n146 B.n145 585
R213 B.n144 B.n143 585
R214 B.n142 B.n141 585
R215 B.n140 B.n139 585
R216 B.n670 B.n119 585
R217 B.n674 B.n119 585
R218 B.n669 B.n118 585
R219 B.n675 B.n118 585
R220 B.n668 B.n667 585
R221 B.n667 B.n114 585
R222 B.n666 B.n113 585
R223 B.n681 B.n113 585
R224 B.n665 B.n112 585
R225 B.n682 B.n112 585
R226 B.n664 B.n111 585
R227 B.n683 B.n111 585
R228 B.n663 B.n662 585
R229 B.n662 B.n107 585
R230 B.n661 B.n106 585
R231 B.n689 B.n106 585
R232 B.n660 B.n105 585
R233 B.n690 B.n105 585
R234 B.n659 B.n104 585
R235 B.n691 B.n104 585
R236 B.n658 B.n657 585
R237 B.n657 B.n100 585
R238 B.n656 B.n99 585
R239 B.n697 B.n99 585
R240 B.n655 B.n98 585
R241 B.n698 B.n98 585
R242 B.n654 B.n97 585
R243 B.n699 B.n97 585
R244 B.n653 B.n652 585
R245 B.n652 B.n93 585
R246 B.n651 B.n92 585
R247 B.n705 B.n92 585
R248 B.n650 B.n91 585
R249 B.n706 B.n91 585
R250 B.n649 B.n90 585
R251 B.n707 B.n90 585
R252 B.n648 B.n647 585
R253 B.n647 B.n86 585
R254 B.n646 B.n85 585
R255 B.n713 B.n85 585
R256 B.n645 B.n84 585
R257 B.n714 B.n84 585
R258 B.n644 B.n83 585
R259 B.n715 B.n83 585
R260 B.n643 B.n642 585
R261 B.n642 B.n79 585
R262 B.n641 B.n78 585
R263 B.n721 B.n78 585
R264 B.n640 B.n77 585
R265 B.n722 B.n77 585
R266 B.n639 B.n76 585
R267 B.n723 B.n76 585
R268 B.n638 B.n637 585
R269 B.n637 B.n72 585
R270 B.n636 B.n71 585
R271 B.n729 B.n71 585
R272 B.n635 B.n70 585
R273 B.n730 B.n70 585
R274 B.n634 B.n69 585
R275 B.n731 B.n69 585
R276 B.n633 B.n632 585
R277 B.n632 B.n65 585
R278 B.n631 B.n64 585
R279 B.n737 B.n64 585
R280 B.n630 B.n63 585
R281 B.n738 B.n63 585
R282 B.n629 B.n62 585
R283 B.n739 B.n62 585
R284 B.n628 B.n627 585
R285 B.n627 B.n58 585
R286 B.n626 B.n57 585
R287 B.n745 B.n57 585
R288 B.n625 B.n56 585
R289 B.n746 B.n56 585
R290 B.n624 B.n55 585
R291 B.n747 B.n55 585
R292 B.n623 B.n622 585
R293 B.n622 B.n51 585
R294 B.n621 B.n50 585
R295 B.n753 B.n50 585
R296 B.n620 B.n49 585
R297 B.n754 B.n49 585
R298 B.n619 B.n48 585
R299 B.n755 B.n48 585
R300 B.n618 B.n617 585
R301 B.n617 B.n44 585
R302 B.n616 B.n43 585
R303 B.n761 B.n43 585
R304 B.n615 B.n42 585
R305 B.n762 B.n42 585
R306 B.n614 B.n41 585
R307 B.n763 B.n41 585
R308 B.n613 B.n612 585
R309 B.n612 B.n40 585
R310 B.n611 B.n36 585
R311 B.n769 B.n36 585
R312 B.n610 B.n35 585
R313 B.n770 B.n35 585
R314 B.n609 B.n34 585
R315 B.n771 B.n34 585
R316 B.n608 B.n607 585
R317 B.n607 B.n30 585
R318 B.n606 B.n29 585
R319 B.n777 B.n29 585
R320 B.n605 B.n28 585
R321 B.n778 B.n28 585
R322 B.n604 B.n27 585
R323 B.n779 B.n27 585
R324 B.n603 B.n602 585
R325 B.n602 B.n23 585
R326 B.n601 B.n22 585
R327 B.n785 B.n22 585
R328 B.n600 B.n21 585
R329 B.n786 B.n21 585
R330 B.n599 B.n20 585
R331 B.n787 B.n20 585
R332 B.n598 B.n597 585
R333 B.n597 B.n19 585
R334 B.n596 B.n15 585
R335 B.n793 B.n15 585
R336 B.n595 B.n14 585
R337 B.n794 B.n14 585
R338 B.n594 B.n13 585
R339 B.n795 B.n13 585
R340 B.n593 B.n592 585
R341 B.n592 B.n12 585
R342 B.n591 B.n590 585
R343 B.n591 B.n8 585
R344 B.n589 B.n7 585
R345 B.n802 B.n7 585
R346 B.n588 B.n6 585
R347 B.n803 B.n6 585
R348 B.n587 B.n5 585
R349 B.n804 B.n5 585
R350 B.n586 B.n585 585
R351 B.n585 B.n4 585
R352 B.n584 B.n191 585
R353 B.n584 B.n583 585
R354 B.n574 B.n192 585
R355 B.n193 B.n192 585
R356 B.n576 B.n575 585
R357 B.n577 B.n576 585
R358 B.n573 B.n198 585
R359 B.n198 B.n197 585
R360 B.n572 B.n571 585
R361 B.n571 B.n570 585
R362 B.n200 B.n199 585
R363 B.n563 B.n200 585
R364 B.n562 B.n561 585
R365 B.n564 B.n562 585
R366 B.n560 B.n205 585
R367 B.n205 B.n204 585
R368 B.n559 B.n558 585
R369 B.n558 B.n557 585
R370 B.n207 B.n206 585
R371 B.n208 B.n207 585
R372 B.n550 B.n549 585
R373 B.n551 B.n550 585
R374 B.n548 B.n213 585
R375 B.n213 B.n212 585
R376 B.n547 B.n546 585
R377 B.n546 B.n545 585
R378 B.n215 B.n214 585
R379 B.n216 B.n215 585
R380 B.n538 B.n537 585
R381 B.n539 B.n538 585
R382 B.n536 B.n221 585
R383 B.n221 B.n220 585
R384 B.n535 B.n534 585
R385 B.n534 B.n533 585
R386 B.n223 B.n222 585
R387 B.n526 B.n223 585
R388 B.n525 B.n524 585
R389 B.n527 B.n525 585
R390 B.n523 B.n228 585
R391 B.n228 B.n227 585
R392 B.n522 B.n521 585
R393 B.n521 B.n520 585
R394 B.n230 B.n229 585
R395 B.n231 B.n230 585
R396 B.n513 B.n512 585
R397 B.n514 B.n513 585
R398 B.n511 B.n236 585
R399 B.n236 B.n235 585
R400 B.n510 B.n509 585
R401 B.n509 B.n508 585
R402 B.n238 B.n237 585
R403 B.n239 B.n238 585
R404 B.n501 B.n500 585
R405 B.n502 B.n501 585
R406 B.n499 B.n244 585
R407 B.n244 B.n243 585
R408 B.n498 B.n497 585
R409 B.n497 B.n496 585
R410 B.n246 B.n245 585
R411 B.n247 B.n246 585
R412 B.n489 B.n488 585
R413 B.n490 B.n489 585
R414 B.n487 B.n252 585
R415 B.n252 B.n251 585
R416 B.n486 B.n485 585
R417 B.n485 B.n484 585
R418 B.n254 B.n253 585
R419 B.n255 B.n254 585
R420 B.n477 B.n476 585
R421 B.n478 B.n477 585
R422 B.n475 B.n260 585
R423 B.n260 B.n259 585
R424 B.n474 B.n473 585
R425 B.n473 B.n472 585
R426 B.n262 B.n261 585
R427 B.n263 B.n262 585
R428 B.n465 B.n464 585
R429 B.n466 B.n465 585
R430 B.n463 B.n268 585
R431 B.n268 B.n267 585
R432 B.n462 B.n461 585
R433 B.n461 B.n460 585
R434 B.n270 B.n269 585
R435 B.n271 B.n270 585
R436 B.n453 B.n452 585
R437 B.n454 B.n453 585
R438 B.n451 B.n276 585
R439 B.n276 B.n275 585
R440 B.n450 B.n449 585
R441 B.n449 B.n448 585
R442 B.n278 B.n277 585
R443 B.n279 B.n278 585
R444 B.n441 B.n440 585
R445 B.n442 B.n441 585
R446 B.n439 B.n284 585
R447 B.n284 B.n283 585
R448 B.n438 B.n437 585
R449 B.n437 B.n436 585
R450 B.n286 B.n285 585
R451 B.n287 B.n286 585
R452 B.n429 B.n428 585
R453 B.n430 B.n429 585
R454 B.n427 B.n292 585
R455 B.n292 B.n291 585
R456 B.n426 B.n425 585
R457 B.n425 B.n424 585
R458 B.n294 B.n293 585
R459 B.n295 B.n294 585
R460 B.n417 B.n416 585
R461 B.n418 B.n417 585
R462 B.n415 B.n300 585
R463 B.n300 B.n299 585
R464 B.n414 B.n413 585
R465 B.n413 B.n412 585
R466 B.n302 B.n301 585
R467 B.n303 B.n302 585
R468 B.n405 B.n404 585
R469 B.n406 B.n405 585
R470 B.n403 B.n308 585
R471 B.n308 B.n307 585
R472 B.n402 B.n401 585
R473 B.n401 B.n400 585
R474 B.n310 B.n309 585
R475 B.n311 B.n310 585
R476 B.n393 B.n392 585
R477 B.n394 B.n393 585
R478 B.n391 B.n316 585
R479 B.n316 B.n315 585
R480 B.n385 B.n384 585
R481 B.n383 B.n331 585
R482 B.n382 B.n330 585
R483 B.n387 B.n330 585
R484 B.n381 B.n380 585
R485 B.n379 B.n378 585
R486 B.n377 B.n376 585
R487 B.n375 B.n374 585
R488 B.n373 B.n372 585
R489 B.n371 B.n370 585
R490 B.n369 B.n368 585
R491 B.n367 B.n366 585
R492 B.n365 B.n364 585
R493 B.n363 B.n362 585
R494 B.n361 B.n360 585
R495 B.n359 B.n358 585
R496 B.n357 B.n356 585
R497 B.n355 B.n354 585
R498 B.n353 B.n352 585
R499 B.n350 B.n349 585
R500 B.n348 B.n347 585
R501 B.n346 B.n345 585
R502 B.n344 B.n343 585
R503 B.n342 B.n341 585
R504 B.n340 B.n339 585
R505 B.n338 B.n337 585
R506 B.n318 B.n317 585
R507 B.n390 B.n389 585
R508 B.n314 B.n313 585
R509 B.n315 B.n314 585
R510 B.n396 B.n395 585
R511 B.n395 B.n394 585
R512 B.n397 B.n312 585
R513 B.n312 B.n311 585
R514 B.n399 B.n398 585
R515 B.n400 B.n399 585
R516 B.n306 B.n305 585
R517 B.n307 B.n306 585
R518 B.n408 B.n407 585
R519 B.n407 B.n406 585
R520 B.n409 B.n304 585
R521 B.n304 B.n303 585
R522 B.n411 B.n410 585
R523 B.n412 B.n411 585
R524 B.n298 B.n297 585
R525 B.n299 B.n298 585
R526 B.n420 B.n419 585
R527 B.n419 B.n418 585
R528 B.n421 B.n296 585
R529 B.n296 B.n295 585
R530 B.n423 B.n422 585
R531 B.n424 B.n423 585
R532 B.n290 B.n289 585
R533 B.n291 B.n290 585
R534 B.n432 B.n431 585
R535 B.n431 B.n430 585
R536 B.n433 B.n288 585
R537 B.n288 B.n287 585
R538 B.n435 B.n434 585
R539 B.n436 B.n435 585
R540 B.n282 B.n281 585
R541 B.n283 B.n282 585
R542 B.n444 B.n443 585
R543 B.n443 B.n442 585
R544 B.n445 B.n280 585
R545 B.n280 B.n279 585
R546 B.n447 B.n446 585
R547 B.n448 B.n447 585
R548 B.n274 B.n273 585
R549 B.n275 B.n274 585
R550 B.n456 B.n455 585
R551 B.n455 B.n454 585
R552 B.n457 B.n272 585
R553 B.n272 B.n271 585
R554 B.n459 B.n458 585
R555 B.n460 B.n459 585
R556 B.n266 B.n265 585
R557 B.n267 B.n266 585
R558 B.n468 B.n467 585
R559 B.n467 B.n466 585
R560 B.n469 B.n264 585
R561 B.n264 B.n263 585
R562 B.n471 B.n470 585
R563 B.n472 B.n471 585
R564 B.n258 B.n257 585
R565 B.n259 B.n258 585
R566 B.n480 B.n479 585
R567 B.n479 B.n478 585
R568 B.n481 B.n256 585
R569 B.n256 B.n255 585
R570 B.n483 B.n482 585
R571 B.n484 B.n483 585
R572 B.n250 B.n249 585
R573 B.n251 B.n250 585
R574 B.n492 B.n491 585
R575 B.n491 B.n490 585
R576 B.n493 B.n248 585
R577 B.n248 B.n247 585
R578 B.n495 B.n494 585
R579 B.n496 B.n495 585
R580 B.n242 B.n241 585
R581 B.n243 B.n242 585
R582 B.n504 B.n503 585
R583 B.n503 B.n502 585
R584 B.n505 B.n240 585
R585 B.n240 B.n239 585
R586 B.n507 B.n506 585
R587 B.n508 B.n507 585
R588 B.n234 B.n233 585
R589 B.n235 B.n234 585
R590 B.n516 B.n515 585
R591 B.n515 B.n514 585
R592 B.n517 B.n232 585
R593 B.n232 B.n231 585
R594 B.n519 B.n518 585
R595 B.n520 B.n519 585
R596 B.n226 B.n225 585
R597 B.n227 B.n226 585
R598 B.n529 B.n528 585
R599 B.n528 B.n527 585
R600 B.n530 B.n224 585
R601 B.n526 B.n224 585
R602 B.n532 B.n531 585
R603 B.n533 B.n532 585
R604 B.n219 B.n218 585
R605 B.n220 B.n219 585
R606 B.n541 B.n540 585
R607 B.n540 B.n539 585
R608 B.n542 B.n217 585
R609 B.n217 B.n216 585
R610 B.n544 B.n543 585
R611 B.n545 B.n544 585
R612 B.n211 B.n210 585
R613 B.n212 B.n211 585
R614 B.n553 B.n552 585
R615 B.n552 B.n551 585
R616 B.n554 B.n209 585
R617 B.n209 B.n208 585
R618 B.n556 B.n555 585
R619 B.n557 B.n556 585
R620 B.n203 B.n202 585
R621 B.n204 B.n203 585
R622 B.n566 B.n565 585
R623 B.n565 B.n564 585
R624 B.n567 B.n201 585
R625 B.n563 B.n201 585
R626 B.n569 B.n568 585
R627 B.n570 B.n569 585
R628 B.n196 B.n195 585
R629 B.n197 B.n196 585
R630 B.n579 B.n578 585
R631 B.n578 B.n577 585
R632 B.n580 B.n194 585
R633 B.n194 B.n193 585
R634 B.n582 B.n581 585
R635 B.n583 B.n582 585
R636 B.n3 B.n0 585
R637 B.n4 B.n3 585
R638 B.n801 B.n1 585
R639 B.n802 B.n801 585
R640 B.n800 B.n799 585
R641 B.n800 B.n8 585
R642 B.n798 B.n9 585
R643 B.n12 B.n9 585
R644 B.n797 B.n796 585
R645 B.n796 B.n795 585
R646 B.n11 B.n10 585
R647 B.n794 B.n11 585
R648 B.n792 B.n791 585
R649 B.n793 B.n792 585
R650 B.n790 B.n16 585
R651 B.n19 B.n16 585
R652 B.n789 B.n788 585
R653 B.n788 B.n787 585
R654 B.n18 B.n17 585
R655 B.n786 B.n18 585
R656 B.n784 B.n783 585
R657 B.n785 B.n784 585
R658 B.n782 B.n24 585
R659 B.n24 B.n23 585
R660 B.n781 B.n780 585
R661 B.n780 B.n779 585
R662 B.n26 B.n25 585
R663 B.n778 B.n26 585
R664 B.n776 B.n775 585
R665 B.n777 B.n776 585
R666 B.n774 B.n31 585
R667 B.n31 B.n30 585
R668 B.n773 B.n772 585
R669 B.n772 B.n771 585
R670 B.n33 B.n32 585
R671 B.n770 B.n33 585
R672 B.n768 B.n767 585
R673 B.n769 B.n768 585
R674 B.n766 B.n37 585
R675 B.n40 B.n37 585
R676 B.n765 B.n764 585
R677 B.n764 B.n763 585
R678 B.n39 B.n38 585
R679 B.n762 B.n39 585
R680 B.n760 B.n759 585
R681 B.n761 B.n760 585
R682 B.n758 B.n45 585
R683 B.n45 B.n44 585
R684 B.n757 B.n756 585
R685 B.n756 B.n755 585
R686 B.n47 B.n46 585
R687 B.n754 B.n47 585
R688 B.n752 B.n751 585
R689 B.n753 B.n752 585
R690 B.n750 B.n52 585
R691 B.n52 B.n51 585
R692 B.n749 B.n748 585
R693 B.n748 B.n747 585
R694 B.n54 B.n53 585
R695 B.n746 B.n54 585
R696 B.n744 B.n743 585
R697 B.n745 B.n744 585
R698 B.n742 B.n59 585
R699 B.n59 B.n58 585
R700 B.n741 B.n740 585
R701 B.n740 B.n739 585
R702 B.n61 B.n60 585
R703 B.n738 B.n61 585
R704 B.n736 B.n735 585
R705 B.n737 B.n736 585
R706 B.n734 B.n66 585
R707 B.n66 B.n65 585
R708 B.n733 B.n732 585
R709 B.n732 B.n731 585
R710 B.n68 B.n67 585
R711 B.n730 B.n68 585
R712 B.n728 B.n727 585
R713 B.n729 B.n728 585
R714 B.n726 B.n73 585
R715 B.n73 B.n72 585
R716 B.n725 B.n724 585
R717 B.n724 B.n723 585
R718 B.n75 B.n74 585
R719 B.n722 B.n75 585
R720 B.n720 B.n719 585
R721 B.n721 B.n720 585
R722 B.n718 B.n80 585
R723 B.n80 B.n79 585
R724 B.n717 B.n716 585
R725 B.n716 B.n715 585
R726 B.n82 B.n81 585
R727 B.n714 B.n82 585
R728 B.n712 B.n711 585
R729 B.n713 B.n712 585
R730 B.n710 B.n87 585
R731 B.n87 B.n86 585
R732 B.n709 B.n708 585
R733 B.n708 B.n707 585
R734 B.n89 B.n88 585
R735 B.n706 B.n89 585
R736 B.n704 B.n703 585
R737 B.n705 B.n704 585
R738 B.n702 B.n94 585
R739 B.n94 B.n93 585
R740 B.n701 B.n700 585
R741 B.n700 B.n699 585
R742 B.n96 B.n95 585
R743 B.n698 B.n96 585
R744 B.n696 B.n695 585
R745 B.n697 B.n696 585
R746 B.n694 B.n101 585
R747 B.n101 B.n100 585
R748 B.n693 B.n692 585
R749 B.n692 B.n691 585
R750 B.n103 B.n102 585
R751 B.n690 B.n103 585
R752 B.n688 B.n687 585
R753 B.n689 B.n688 585
R754 B.n686 B.n108 585
R755 B.n108 B.n107 585
R756 B.n685 B.n684 585
R757 B.n684 B.n683 585
R758 B.n110 B.n109 585
R759 B.n682 B.n110 585
R760 B.n680 B.n679 585
R761 B.n681 B.n680 585
R762 B.n678 B.n115 585
R763 B.n115 B.n114 585
R764 B.n677 B.n676 585
R765 B.n676 B.n675 585
R766 B.n117 B.n116 585
R767 B.n674 B.n117 585
R768 B.n805 B.n804 585
R769 B.n803 B.n2 585
R770 B.n139 B.n117 458.866
R771 B.n672 B.n119 458.866
R772 B.n389 B.n316 458.866
R773 B.n385 B.n314 458.866
R774 B.n137 B.t14 310.524
R775 B.n134 B.t4 310.524
R776 B.n335 B.t9 310.524
R777 B.n332 B.t12 310.524
R778 B.n673 B.n132 256.663
R779 B.n673 B.n131 256.663
R780 B.n673 B.n130 256.663
R781 B.n673 B.n129 256.663
R782 B.n673 B.n128 256.663
R783 B.n673 B.n127 256.663
R784 B.n673 B.n126 256.663
R785 B.n673 B.n125 256.663
R786 B.n673 B.n124 256.663
R787 B.n673 B.n123 256.663
R788 B.n673 B.n122 256.663
R789 B.n673 B.n121 256.663
R790 B.n673 B.n120 256.663
R791 B.n387 B.n386 256.663
R792 B.n387 B.n319 256.663
R793 B.n387 B.n320 256.663
R794 B.n387 B.n321 256.663
R795 B.n387 B.n322 256.663
R796 B.n387 B.n323 256.663
R797 B.n387 B.n324 256.663
R798 B.n387 B.n325 256.663
R799 B.n387 B.n326 256.663
R800 B.n387 B.n327 256.663
R801 B.n387 B.n328 256.663
R802 B.n387 B.n329 256.663
R803 B.n388 B.n387 256.663
R804 B.n807 B.n806 256.663
R805 B.n138 B.t15 235.082
R806 B.n135 B.t5 235.082
R807 B.n336 B.t8 235.082
R808 B.n333 B.t11 235.082
R809 B.n137 B.t13 209.965
R810 B.n134 B.t2 209.965
R811 B.n335 B.t6 209.965
R812 B.n332 B.t10 209.965
R813 B.n387 B.n315 201.32
R814 B.n674 B.n673 201.32
R815 B.n143 B.n142 163.367
R816 B.n147 B.n146 163.367
R817 B.n151 B.n150 163.367
R818 B.n155 B.n154 163.367
R819 B.n160 B.n159 163.367
R820 B.n164 B.n163 163.367
R821 B.n168 B.n167 163.367
R822 B.n172 B.n171 163.367
R823 B.n176 B.n175 163.367
R824 B.n180 B.n179 163.367
R825 B.n184 B.n183 163.367
R826 B.n188 B.n187 163.367
R827 B.n672 B.n133 163.367
R828 B.n393 B.n316 163.367
R829 B.n393 B.n310 163.367
R830 B.n401 B.n310 163.367
R831 B.n401 B.n308 163.367
R832 B.n405 B.n308 163.367
R833 B.n405 B.n302 163.367
R834 B.n413 B.n302 163.367
R835 B.n413 B.n300 163.367
R836 B.n417 B.n300 163.367
R837 B.n417 B.n294 163.367
R838 B.n425 B.n294 163.367
R839 B.n425 B.n292 163.367
R840 B.n429 B.n292 163.367
R841 B.n429 B.n286 163.367
R842 B.n437 B.n286 163.367
R843 B.n437 B.n284 163.367
R844 B.n441 B.n284 163.367
R845 B.n441 B.n278 163.367
R846 B.n449 B.n278 163.367
R847 B.n449 B.n276 163.367
R848 B.n453 B.n276 163.367
R849 B.n453 B.n270 163.367
R850 B.n461 B.n270 163.367
R851 B.n461 B.n268 163.367
R852 B.n465 B.n268 163.367
R853 B.n465 B.n262 163.367
R854 B.n473 B.n262 163.367
R855 B.n473 B.n260 163.367
R856 B.n477 B.n260 163.367
R857 B.n477 B.n254 163.367
R858 B.n485 B.n254 163.367
R859 B.n485 B.n252 163.367
R860 B.n489 B.n252 163.367
R861 B.n489 B.n246 163.367
R862 B.n497 B.n246 163.367
R863 B.n497 B.n244 163.367
R864 B.n501 B.n244 163.367
R865 B.n501 B.n238 163.367
R866 B.n509 B.n238 163.367
R867 B.n509 B.n236 163.367
R868 B.n513 B.n236 163.367
R869 B.n513 B.n230 163.367
R870 B.n521 B.n230 163.367
R871 B.n521 B.n228 163.367
R872 B.n525 B.n228 163.367
R873 B.n525 B.n223 163.367
R874 B.n534 B.n223 163.367
R875 B.n534 B.n221 163.367
R876 B.n538 B.n221 163.367
R877 B.n538 B.n215 163.367
R878 B.n546 B.n215 163.367
R879 B.n546 B.n213 163.367
R880 B.n550 B.n213 163.367
R881 B.n550 B.n207 163.367
R882 B.n558 B.n207 163.367
R883 B.n558 B.n205 163.367
R884 B.n562 B.n205 163.367
R885 B.n562 B.n200 163.367
R886 B.n571 B.n200 163.367
R887 B.n571 B.n198 163.367
R888 B.n576 B.n198 163.367
R889 B.n576 B.n192 163.367
R890 B.n584 B.n192 163.367
R891 B.n585 B.n584 163.367
R892 B.n585 B.n5 163.367
R893 B.n6 B.n5 163.367
R894 B.n7 B.n6 163.367
R895 B.n591 B.n7 163.367
R896 B.n592 B.n591 163.367
R897 B.n592 B.n13 163.367
R898 B.n14 B.n13 163.367
R899 B.n15 B.n14 163.367
R900 B.n597 B.n15 163.367
R901 B.n597 B.n20 163.367
R902 B.n21 B.n20 163.367
R903 B.n22 B.n21 163.367
R904 B.n602 B.n22 163.367
R905 B.n602 B.n27 163.367
R906 B.n28 B.n27 163.367
R907 B.n29 B.n28 163.367
R908 B.n607 B.n29 163.367
R909 B.n607 B.n34 163.367
R910 B.n35 B.n34 163.367
R911 B.n36 B.n35 163.367
R912 B.n612 B.n36 163.367
R913 B.n612 B.n41 163.367
R914 B.n42 B.n41 163.367
R915 B.n43 B.n42 163.367
R916 B.n617 B.n43 163.367
R917 B.n617 B.n48 163.367
R918 B.n49 B.n48 163.367
R919 B.n50 B.n49 163.367
R920 B.n622 B.n50 163.367
R921 B.n622 B.n55 163.367
R922 B.n56 B.n55 163.367
R923 B.n57 B.n56 163.367
R924 B.n627 B.n57 163.367
R925 B.n627 B.n62 163.367
R926 B.n63 B.n62 163.367
R927 B.n64 B.n63 163.367
R928 B.n632 B.n64 163.367
R929 B.n632 B.n69 163.367
R930 B.n70 B.n69 163.367
R931 B.n71 B.n70 163.367
R932 B.n637 B.n71 163.367
R933 B.n637 B.n76 163.367
R934 B.n77 B.n76 163.367
R935 B.n78 B.n77 163.367
R936 B.n642 B.n78 163.367
R937 B.n642 B.n83 163.367
R938 B.n84 B.n83 163.367
R939 B.n85 B.n84 163.367
R940 B.n647 B.n85 163.367
R941 B.n647 B.n90 163.367
R942 B.n91 B.n90 163.367
R943 B.n92 B.n91 163.367
R944 B.n652 B.n92 163.367
R945 B.n652 B.n97 163.367
R946 B.n98 B.n97 163.367
R947 B.n99 B.n98 163.367
R948 B.n657 B.n99 163.367
R949 B.n657 B.n104 163.367
R950 B.n105 B.n104 163.367
R951 B.n106 B.n105 163.367
R952 B.n662 B.n106 163.367
R953 B.n662 B.n111 163.367
R954 B.n112 B.n111 163.367
R955 B.n113 B.n112 163.367
R956 B.n667 B.n113 163.367
R957 B.n667 B.n118 163.367
R958 B.n119 B.n118 163.367
R959 B.n331 B.n330 163.367
R960 B.n380 B.n330 163.367
R961 B.n378 B.n377 163.367
R962 B.n374 B.n373 163.367
R963 B.n370 B.n369 163.367
R964 B.n366 B.n365 163.367
R965 B.n362 B.n361 163.367
R966 B.n358 B.n357 163.367
R967 B.n354 B.n353 163.367
R968 B.n349 B.n348 163.367
R969 B.n345 B.n344 163.367
R970 B.n341 B.n340 163.367
R971 B.n337 B.n318 163.367
R972 B.n395 B.n314 163.367
R973 B.n395 B.n312 163.367
R974 B.n399 B.n312 163.367
R975 B.n399 B.n306 163.367
R976 B.n407 B.n306 163.367
R977 B.n407 B.n304 163.367
R978 B.n411 B.n304 163.367
R979 B.n411 B.n298 163.367
R980 B.n419 B.n298 163.367
R981 B.n419 B.n296 163.367
R982 B.n423 B.n296 163.367
R983 B.n423 B.n290 163.367
R984 B.n431 B.n290 163.367
R985 B.n431 B.n288 163.367
R986 B.n435 B.n288 163.367
R987 B.n435 B.n282 163.367
R988 B.n443 B.n282 163.367
R989 B.n443 B.n280 163.367
R990 B.n447 B.n280 163.367
R991 B.n447 B.n274 163.367
R992 B.n455 B.n274 163.367
R993 B.n455 B.n272 163.367
R994 B.n459 B.n272 163.367
R995 B.n459 B.n266 163.367
R996 B.n467 B.n266 163.367
R997 B.n467 B.n264 163.367
R998 B.n471 B.n264 163.367
R999 B.n471 B.n258 163.367
R1000 B.n479 B.n258 163.367
R1001 B.n479 B.n256 163.367
R1002 B.n483 B.n256 163.367
R1003 B.n483 B.n250 163.367
R1004 B.n491 B.n250 163.367
R1005 B.n491 B.n248 163.367
R1006 B.n495 B.n248 163.367
R1007 B.n495 B.n242 163.367
R1008 B.n503 B.n242 163.367
R1009 B.n503 B.n240 163.367
R1010 B.n507 B.n240 163.367
R1011 B.n507 B.n234 163.367
R1012 B.n515 B.n234 163.367
R1013 B.n515 B.n232 163.367
R1014 B.n519 B.n232 163.367
R1015 B.n519 B.n226 163.367
R1016 B.n528 B.n226 163.367
R1017 B.n528 B.n224 163.367
R1018 B.n532 B.n224 163.367
R1019 B.n532 B.n219 163.367
R1020 B.n540 B.n219 163.367
R1021 B.n540 B.n217 163.367
R1022 B.n544 B.n217 163.367
R1023 B.n544 B.n211 163.367
R1024 B.n552 B.n211 163.367
R1025 B.n552 B.n209 163.367
R1026 B.n556 B.n209 163.367
R1027 B.n556 B.n203 163.367
R1028 B.n565 B.n203 163.367
R1029 B.n565 B.n201 163.367
R1030 B.n569 B.n201 163.367
R1031 B.n569 B.n196 163.367
R1032 B.n578 B.n196 163.367
R1033 B.n578 B.n194 163.367
R1034 B.n582 B.n194 163.367
R1035 B.n582 B.n3 163.367
R1036 B.n805 B.n3 163.367
R1037 B.n801 B.n2 163.367
R1038 B.n801 B.n800 163.367
R1039 B.n800 B.n9 163.367
R1040 B.n796 B.n9 163.367
R1041 B.n796 B.n11 163.367
R1042 B.n792 B.n11 163.367
R1043 B.n792 B.n16 163.367
R1044 B.n788 B.n16 163.367
R1045 B.n788 B.n18 163.367
R1046 B.n784 B.n18 163.367
R1047 B.n784 B.n24 163.367
R1048 B.n780 B.n24 163.367
R1049 B.n780 B.n26 163.367
R1050 B.n776 B.n26 163.367
R1051 B.n776 B.n31 163.367
R1052 B.n772 B.n31 163.367
R1053 B.n772 B.n33 163.367
R1054 B.n768 B.n33 163.367
R1055 B.n768 B.n37 163.367
R1056 B.n764 B.n37 163.367
R1057 B.n764 B.n39 163.367
R1058 B.n760 B.n39 163.367
R1059 B.n760 B.n45 163.367
R1060 B.n756 B.n45 163.367
R1061 B.n756 B.n47 163.367
R1062 B.n752 B.n47 163.367
R1063 B.n752 B.n52 163.367
R1064 B.n748 B.n52 163.367
R1065 B.n748 B.n54 163.367
R1066 B.n744 B.n54 163.367
R1067 B.n744 B.n59 163.367
R1068 B.n740 B.n59 163.367
R1069 B.n740 B.n61 163.367
R1070 B.n736 B.n61 163.367
R1071 B.n736 B.n66 163.367
R1072 B.n732 B.n66 163.367
R1073 B.n732 B.n68 163.367
R1074 B.n728 B.n68 163.367
R1075 B.n728 B.n73 163.367
R1076 B.n724 B.n73 163.367
R1077 B.n724 B.n75 163.367
R1078 B.n720 B.n75 163.367
R1079 B.n720 B.n80 163.367
R1080 B.n716 B.n80 163.367
R1081 B.n716 B.n82 163.367
R1082 B.n712 B.n82 163.367
R1083 B.n712 B.n87 163.367
R1084 B.n708 B.n87 163.367
R1085 B.n708 B.n89 163.367
R1086 B.n704 B.n89 163.367
R1087 B.n704 B.n94 163.367
R1088 B.n700 B.n94 163.367
R1089 B.n700 B.n96 163.367
R1090 B.n696 B.n96 163.367
R1091 B.n696 B.n101 163.367
R1092 B.n692 B.n101 163.367
R1093 B.n692 B.n103 163.367
R1094 B.n688 B.n103 163.367
R1095 B.n688 B.n108 163.367
R1096 B.n684 B.n108 163.367
R1097 B.n684 B.n110 163.367
R1098 B.n680 B.n110 163.367
R1099 B.n680 B.n115 163.367
R1100 B.n676 B.n115 163.367
R1101 B.n676 B.n117 163.367
R1102 B.n394 B.n315 123.332
R1103 B.n394 B.n311 123.332
R1104 B.n400 B.n311 123.332
R1105 B.n400 B.n307 123.332
R1106 B.n406 B.n307 123.332
R1107 B.n406 B.n303 123.332
R1108 B.n412 B.n303 123.332
R1109 B.n412 B.n299 123.332
R1110 B.n418 B.n299 123.332
R1111 B.n424 B.n295 123.332
R1112 B.n424 B.n291 123.332
R1113 B.n430 B.n291 123.332
R1114 B.n430 B.n287 123.332
R1115 B.n436 B.n287 123.332
R1116 B.n436 B.n283 123.332
R1117 B.n442 B.n283 123.332
R1118 B.n442 B.n279 123.332
R1119 B.n448 B.n279 123.332
R1120 B.n448 B.n275 123.332
R1121 B.n454 B.n275 123.332
R1122 B.n454 B.n271 123.332
R1123 B.n460 B.n271 123.332
R1124 B.n466 B.n267 123.332
R1125 B.n466 B.n263 123.332
R1126 B.n472 B.n263 123.332
R1127 B.n472 B.n259 123.332
R1128 B.n478 B.n259 123.332
R1129 B.n478 B.n255 123.332
R1130 B.n484 B.n255 123.332
R1131 B.n484 B.n251 123.332
R1132 B.n490 B.n251 123.332
R1133 B.n490 B.n247 123.332
R1134 B.n496 B.n247 123.332
R1135 B.n502 B.n243 123.332
R1136 B.n502 B.n239 123.332
R1137 B.n508 B.n239 123.332
R1138 B.n508 B.n235 123.332
R1139 B.n514 B.n235 123.332
R1140 B.n514 B.n231 123.332
R1141 B.n520 B.n231 123.332
R1142 B.n520 B.n227 123.332
R1143 B.n527 B.n227 123.332
R1144 B.n527 B.n526 123.332
R1145 B.n533 B.n220 123.332
R1146 B.n539 B.n220 123.332
R1147 B.n539 B.n216 123.332
R1148 B.n545 B.n216 123.332
R1149 B.n545 B.n212 123.332
R1150 B.n551 B.n212 123.332
R1151 B.n551 B.n208 123.332
R1152 B.n557 B.n208 123.332
R1153 B.n557 B.n204 123.332
R1154 B.n564 B.n204 123.332
R1155 B.n564 B.n563 123.332
R1156 B.n570 B.n197 123.332
R1157 B.n577 B.n197 123.332
R1158 B.n577 B.n193 123.332
R1159 B.n583 B.n193 123.332
R1160 B.n583 B.n4 123.332
R1161 B.n804 B.n4 123.332
R1162 B.n804 B.n803 123.332
R1163 B.n803 B.n802 123.332
R1164 B.n802 B.n8 123.332
R1165 B.n12 B.n8 123.332
R1166 B.n795 B.n12 123.332
R1167 B.n795 B.n794 123.332
R1168 B.n794 B.n793 123.332
R1169 B.n787 B.n19 123.332
R1170 B.n787 B.n786 123.332
R1171 B.n786 B.n785 123.332
R1172 B.n785 B.n23 123.332
R1173 B.n779 B.n23 123.332
R1174 B.n779 B.n778 123.332
R1175 B.n778 B.n777 123.332
R1176 B.n777 B.n30 123.332
R1177 B.n771 B.n30 123.332
R1178 B.n771 B.n770 123.332
R1179 B.n770 B.n769 123.332
R1180 B.n763 B.n40 123.332
R1181 B.n763 B.n762 123.332
R1182 B.n762 B.n761 123.332
R1183 B.n761 B.n44 123.332
R1184 B.n755 B.n44 123.332
R1185 B.n755 B.n754 123.332
R1186 B.n754 B.n753 123.332
R1187 B.n753 B.n51 123.332
R1188 B.n747 B.n51 123.332
R1189 B.n747 B.n746 123.332
R1190 B.n745 B.n58 123.332
R1191 B.n739 B.n58 123.332
R1192 B.n739 B.n738 123.332
R1193 B.n738 B.n737 123.332
R1194 B.n737 B.n65 123.332
R1195 B.n731 B.n65 123.332
R1196 B.n731 B.n730 123.332
R1197 B.n730 B.n729 123.332
R1198 B.n729 B.n72 123.332
R1199 B.n723 B.n72 123.332
R1200 B.n723 B.n722 123.332
R1201 B.n721 B.n79 123.332
R1202 B.n715 B.n79 123.332
R1203 B.n715 B.n714 123.332
R1204 B.n714 B.n713 123.332
R1205 B.n713 B.n86 123.332
R1206 B.n707 B.n86 123.332
R1207 B.n707 B.n706 123.332
R1208 B.n706 B.n705 123.332
R1209 B.n705 B.n93 123.332
R1210 B.n699 B.n93 123.332
R1211 B.n699 B.n698 123.332
R1212 B.n698 B.n697 123.332
R1213 B.n697 B.n100 123.332
R1214 B.n691 B.n690 123.332
R1215 B.n690 B.n689 123.332
R1216 B.n689 B.n107 123.332
R1217 B.n683 B.n107 123.332
R1218 B.n683 B.n682 123.332
R1219 B.n682 B.n681 123.332
R1220 B.n681 B.n114 123.332
R1221 B.n675 B.n114 123.332
R1222 B.n675 B.n674 123.332
R1223 B.n460 B.t16 105.195
R1224 B.t21 B.n721 105.195
R1225 B.n570 B.t20 101.567
R1226 B.n793 B.t17 101.567
R1227 B.t7 B.n295 97.9395
R1228 B.t3 B.n100 97.9395
R1229 B.n526 B.t18 90.6848
R1230 B.n40 B.t19 90.6848
R1231 B.t1 B.n243 87.0574
R1232 B.n746 B.t0 87.0574
R1233 B.n138 B.n137 75.4429
R1234 B.n135 B.n134 75.4429
R1235 B.n336 B.n335 75.4429
R1236 B.n333 B.n332 75.4429
R1237 B.n139 B.n120 71.676
R1238 B.n143 B.n121 71.676
R1239 B.n147 B.n122 71.676
R1240 B.n151 B.n123 71.676
R1241 B.n155 B.n124 71.676
R1242 B.n160 B.n125 71.676
R1243 B.n164 B.n126 71.676
R1244 B.n168 B.n127 71.676
R1245 B.n172 B.n128 71.676
R1246 B.n176 B.n129 71.676
R1247 B.n180 B.n130 71.676
R1248 B.n184 B.n131 71.676
R1249 B.n188 B.n132 71.676
R1250 B.n133 B.n132 71.676
R1251 B.n187 B.n131 71.676
R1252 B.n183 B.n130 71.676
R1253 B.n179 B.n129 71.676
R1254 B.n175 B.n128 71.676
R1255 B.n171 B.n127 71.676
R1256 B.n167 B.n126 71.676
R1257 B.n163 B.n125 71.676
R1258 B.n159 B.n124 71.676
R1259 B.n154 B.n123 71.676
R1260 B.n150 B.n122 71.676
R1261 B.n146 B.n121 71.676
R1262 B.n142 B.n120 71.676
R1263 B.n386 B.n385 71.676
R1264 B.n380 B.n319 71.676
R1265 B.n377 B.n320 71.676
R1266 B.n373 B.n321 71.676
R1267 B.n369 B.n322 71.676
R1268 B.n365 B.n323 71.676
R1269 B.n361 B.n324 71.676
R1270 B.n357 B.n325 71.676
R1271 B.n353 B.n326 71.676
R1272 B.n348 B.n327 71.676
R1273 B.n344 B.n328 71.676
R1274 B.n340 B.n329 71.676
R1275 B.n388 B.n318 71.676
R1276 B.n386 B.n331 71.676
R1277 B.n378 B.n319 71.676
R1278 B.n374 B.n320 71.676
R1279 B.n370 B.n321 71.676
R1280 B.n366 B.n322 71.676
R1281 B.n362 B.n323 71.676
R1282 B.n358 B.n324 71.676
R1283 B.n354 B.n325 71.676
R1284 B.n349 B.n326 71.676
R1285 B.n345 B.n327 71.676
R1286 B.n341 B.n328 71.676
R1287 B.n337 B.n329 71.676
R1288 B.n389 B.n388 71.676
R1289 B.n806 B.n805 71.676
R1290 B.n806 B.n2 71.676
R1291 B.n157 B.n138 59.5399
R1292 B.n136 B.n135 59.5399
R1293 B.n351 B.n336 59.5399
R1294 B.n334 B.n333 59.5399
R1295 B.n496 B.t1 36.2742
R1296 B.t0 B.n745 36.2742
R1297 B.n533 B.t18 32.6468
R1298 B.n769 B.t19 32.6468
R1299 B.n384 B.n313 29.8151
R1300 B.n391 B.n390 29.8151
R1301 B.n140 B.n116 29.8151
R1302 B.n671 B.n670 29.8151
R1303 B.n418 B.t7 25.3921
R1304 B.n691 B.t3 25.3921
R1305 B.n563 B.t20 21.7647
R1306 B.n19 B.t17 21.7647
R1307 B.t16 B.n267 18.1374
R1308 B.n722 B.t21 18.1374
R1309 B B.n807 18.0485
R1310 B.n396 B.n313 10.6151
R1311 B.n397 B.n396 10.6151
R1312 B.n398 B.n397 10.6151
R1313 B.n398 B.n305 10.6151
R1314 B.n408 B.n305 10.6151
R1315 B.n409 B.n408 10.6151
R1316 B.n410 B.n409 10.6151
R1317 B.n410 B.n297 10.6151
R1318 B.n420 B.n297 10.6151
R1319 B.n421 B.n420 10.6151
R1320 B.n422 B.n421 10.6151
R1321 B.n422 B.n289 10.6151
R1322 B.n432 B.n289 10.6151
R1323 B.n433 B.n432 10.6151
R1324 B.n434 B.n433 10.6151
R1325 B.n434 B.n281 10.6151
R1326 B.n444 B.n281 10.6151
R1327 B.n445 B.n444 10.6151
R1328 B.n446 B.n445 10.6151
R1329 B.n446 B.n273 10.6151
R1330 B.n456 B.n273 10.6151
R1331 B.n457 B.n456 10.6151
R1332 B.n458 B.n457 10.6151
R1333 B.n458 B.n265 10.6151
R1334 B.n468 B.n265 10.6151
R1335 B.n469 B.n468 10.6151
R1336 B.n470 B.n469 10.6151
R1337 B.n470 B.n257 10.6151
R1338 B.n480 B.n257 10.6151
R1339 B.n481 B.n480 10.6151
R1340 B.n482 B.n481 10.6151
R1341 B.n482 B.n249 10.6151
R1342 B.n492 B.n249 10.6151
R1343 B.n493 B.n492 10.6151
R1344 B.n494 B.n493 10.6151
R1345 B.n494 B.n241 10.6151
R1346 B.n504 B.n241 10.6151
R1347 B.n505 B.n504 10.6151
R1348 B.n506 B.n505 10.6151
R1349 B.n506 B.n233 10.6151
R1350 B.n516 B.n233 10.6151
R1351 B.n517 B.n516 10.6151
R1352 B.n518 B.n517 10.6151
R1353 B.n518 B.n225 10.6151
R1354 B.n529 B.n225 10.6151
R1355 B.n530 B.n529 10.6151
R1356 B.n531 B.n530 10.6151
R1357 B.n531 B.n218 10.6151
R1358 B.n541 B.n218 10.6151
R1359 B.n542 B.n541 10.6151
R1360 B.n543 B.n542 10.6151
R1361 B.n543 B.n210 10.6151
R1362 B.n553 B.n210 10.6151
R1363 B.n554 B.n553 10.6151
R1364 B.n555 B.n554 10.6151
R1365 B.n555 B.n202 10.6151
R1366 B.n566 B.n202 10.6151
R1367 B.n567 B.n566 10.6151
R1368 B.n568 B.n567 10.6151
R1369 B.n568 B.n195 10.6151
R1370 B.n579 B.n195 10.6151
R1371 B.n580 B.n579 10.6151
R1372 B.n581 B.n580 10.6151
R1373 B.n581 B.n0 10.6151
R1374 B.n384 B.n383 10.6151
R1375 B.n383 B.n382 10.6151
R1376 B.n382 B.n381 10.6151
R1377 B.n381 B.n379 10.6151
R1378 B.n379 B.n376 10.6151
R1379 B.n376 B.n375 10.6151
R1380 B.n375 B.n372 10.6151
R1381 B.n372 B.n371 10.6151
R1382 B.n368 B.n367 10.6151
R1383 B.n367 B.n364 10.6151
R1384 B.n364 B.n363 10.6151
R1385 B.n363 B.n360 10.6151
R1386 B.n360 B.n359 10.6151
R1387 B.n359 B.n356 10.6151
R1388 B.n356 B.n355 10.6151
R1389 B.n355 B.n352 10.6151
R1390 B.n350 B.n347 10.6151
R1391 B.n347 B.n346 10.6151
R1392 B.n346 B.n343 10.6151
R1393 B.n343 B.n342 10.6151
R1394 B.n342 B.n339 10.6151
R1395 B.n339 B.n338 10.6151
R1396 B.n338 B.n317 10.6151
R1397 B.n390 B.n317 10.6151
R1398 B.n392 B.n391 10.6151
R1399 B.n392 B.n309 10.6151
R1400 B.n402 B.n309 10.6151
R1401 B.n403 B.n402 10.6151
R1402 B.n404 B.n403 10.6151
R1403 B.n404 B.n301 10.6151
R1404 B.n414 B.n301 10.6151
R1405 B.n415 B.n414 10.6151
R1406 B.n416 B.n415 10.6151
R1407 B.n416 B.n293 10.6151
R1408 B.n426 B.n293 10.6151
R1409 B.n427 B.n426 10.6151
R1410 B.n428 B.n427 10.6151
R1411 B.n428 B.n285 10.6151
R1412 B.n438 B.n285 10.6151
R1413 B.n439 B.n438 10.6151
R1414 B.n440 B.n439 10.6151
R1415 B.n440 B.n277 10.6151
R1416 B.n450 B.n277 10.6151
R1417 B.n451 B.n450 10.6151
R1418 B.n452 B.n451 10.6151
R1419 B.n452 B.n269 10.6151
R1420 B.n462 B.n269 10.6151
R1421 B.n463 B.n462 10.6151
R1422 B.n464 B.n463 10.6151
R1423 B.n464 B.n261 10.6151
R1424 B.n474 B.n261 10.6151
R1425 B.n475 B.n474 10.6151
R1426 B.n476 B.n475 10.6151
R1427 B.n476 B.n253 10.6151
R1428 B.n486 B.n253 10.6151
R1429 B.n487 B.n486 10.6151
R1430 B.n488 B.n487 10.6151
R1431 B.n488 B.n245 10.6151
R1432 B.n498 B.n245 10.6151
R1433 B.n499 B.n498 10.6151
R1434 B.n500 B.n499 10.6151
R1435 B.n500 B.n237 10.6151
R1436 B.n510 B.n237 10.6151
R1437 B.n511 B.n510 10.6151
R1438 B.n512 B.n511 10.6151
R1439 B.n512 B.n229 10.6151
R1440 B.n522 B.n229 10.6151
R1441 B.n523 B.n522 10.6151
R1442 B.n524 B.n523 10.6151
R1443 B.n524 B.n222 10.6151
R1444 B.n535 B.n222 10.6151
R1445 B.n536 B.n535 10.6151
R1446 B.n537 B.n536 10.6151
R1447 B.n537 B.n214 10.6151
R1448 B.n547 B.n214 10.6151
R1449 B.n548 B.n547 10.6151
R1450 B.n549 B.n548 10.6151
R1451 B.n549 B.n206 10.6151
R1452 B.n559 B.n206 10.6151
R1453 B.n560 B.n559 10.6151
R1454 B.n561 B.n560 10.6151
R1455 B.n561 B.n199 10.6151
R1456 B.n572 B.n199 10.6151
R1457 B.n573 B.n572 10.6151
R1458 B.n575 B.n573 10.6151
R1459 B.n575 B.n574 10.6151
R1460 B.n574 B.n191 10.6151
R1461 B.n586 B.n191 10.6151
R1462 B.n587 B.n586 10.6151
R1463 B.n588 B.n587 10.6151
R1464 B.n589 B.n588 10.6151
R1465 B.n590 B.n589 10.6151
R1466 B.n593 B.n590 10.6151
R1467 B.n594 B.n593 10.6151
R1468 B.n595 B.n594 10.6151
R1469 B.n596 B.n595 10.6151
R1470 B.n598 B.n596 10.6151
R1471 B.n599 B.n598 10.6151
R1472 B.n600 B.n599 10.6151
R1473 B.n601 B.n600 10.6151
R1474 B.n603 B.n601 10.6151
R1475 B.n604 B.n603 10.6151
R1476 B.n605 B.n604 10.6151
R1477 B.n606 B.n605 10.6151
R1478 B.n608 B.n606 10.6151
R1479 B.n609 B.n608 10.6151
R1480 B.n610 B.n609 10.6151
R1481 B.n611 B.n610 10.6151
R1482 B.n613 B.n611 10.6151
R1483 B.n614 B.n613 10.6151
R1484 B.n615 B.n614 10.6151
R1485 B.n616 B.n615 10.6151
R1486 B.n618 B.n616 10.6151
R1487 B.n619 B.n618 10.6151
R1488 B.n620 B.n619 10.6151
R1489 B.n621 B.n620 10.6151
R1490 B.n623 B.n621 10.6151
R1491 B.n624 B.n623 10.6151
R1492 B.n625 B.n624 10.6151
R1493 B.n626 B.n625 10.6151
R1494 B.n628 B.n626 10.6151
R1495 B.n629 B.n628 10.6151
R1496 B.n630 B.n629 10.6151
R1497 B.n631 B.n630 10.6151
R1498 B.n633 B.n631 10.6151
R1499 B.n634 B.n633 10.6151
R1500 B.n635 B.n634 10.6151
R1501 B.n636 B.n635 10.6151
R1502 B.n638 B.n636 10.6151
R1503 B.n639 B.n638 10.6151
R1504 B.n640 B.n639 10.6151
R1505 B.n641 B.n640 10.6151
R1506 B.n643 B.n641 10.6151
R1507 B.n644 B.n643 10.6151
R1508 B.n645 B.n644 10.6151
R1509 B.n646 B.n645 10.6151
R1510 B.n648 B.n646 10.6151
R1511 B.n649 B.n648 10.6151
R1512 B.n650 B.n649 10.6151
R1513 B.n651 B.n650 10.6151
R1514 B.n653 B.n651 10.6151
R1515 B.n654 B.n653 10.6151
R1516 B.n655 B.n654 10.6151
R1517 B.n656 B.n655 10.6151
R1518 B.n658 B.n656 10.6151
R1519 B.n659 B.n658 10.6151
R1520 B.n660 B.n659 10.6151
R1521 B.n661 B.n660 10.6151
R1522 B.n663 B.n661 10.6151
R1523 B.n664 B.n663 10.6151
R1524 B.n665 B.n664 10.6151
R1525 B.n666 B.n665 10.6151
R1526 B.n668 B.n666 10.6151
R1527 B.n669 B.n668 10.6151
R1528 B.n670 B.n669 10.6151
R1529 B.n799 B.n1 10.6151
R1530 B.n799 B.n798 10.6151
R1531 B.n798 B.n797 10.6151
R1532 B.n797 B.n10 10.6151
R1533 B.n791 B.n10 10.6151
R1534 B.n791 B.n790 10.6151
R1535 B.n790 B.n789 10.6151
R1536 B.n789 B.n17 10.6151
R1537 B.n783 B.n17 10.6151
R1538 B.n783 B.n782 10.6151
R1539 B.n782 B.n781 10.6151
R1540 B.n781 B.n25 10.6151
R1541 B.n775 B.n25 10.6151
R1542 B.n775 B.n774 10.6151
R1543 B.n774 B.n773 10.6151
R1544 B.n773 B.n32 10.6151
R1545 B.n767 B.n32 10.6151
R1546 B.n767 B.n766 10.6151
R1547 B.n766 B.n765 10.6151
R1548 B.n765 B.n38 10.6151
R1549 B.n759 B.n38 10.6151
R1550 B.n759 B.n758 10.6151
R1551 B.n758 B.n757 10.6151
R1552 B.n757 B.n46 10.6151
R1553 B.n751 B.n46 10.6151
R1554 B.n751 B.n750 10.6151
R1555 B.n750 B.n749 10.6151
R1556 B.n749 B.n53 10.6151
R1557 B.n743 B.n53 10.6151
R1558 B.n743 B.n742 10.6151
R1559 B.n742 B.n741 10.6151
R1560 B.n741 B.n60 10.6151
R1561 B.n735 B.n60 10.6151
R1562 B.n735 B.n734 10.6151
R1563 B.n734 B.n733 10.6151
R1564 B.n733 B.n67 10.6151
R1565 B.n727 B.n67 10.6151
R1566 B.n727 B.n726 10.6151
R1567 B.n726 B.n725 10.6151
R1568 B.n725 B.n74 10.6151
R1569 B.n719 B.n74 10.6151
R1570 B.n719 B.n718 10.6151
R1571 B.n718 B.n717 10.6151
R1572 B.n717 B.n81 10.6151
R1573 B.n711 B.n81 10.6151
R1574 B.n711 B.n710 10.6151
R1575 B.n710 B.n709 10.6151
R1576 B.n709 B.n88 10.6151
R1577 B.n703 B.n88 10.6151
R1578 B.n703 B.n702 10.6151
R1579 B.n702 B.n701 10.6151
R1580 B.n701 B.n95 10.6151
R1581 B.n695 B.n95 10.6151
R1582 B.n695 B.n694 10.6151
R1583 B.n694 B.n693 10.6151
R1584 B.n693 B.n102 10.6151
R1585 B.n687 B.n102 10.6151
R1586 B.n687 B.n686 10.6151
R1587 B.n686 B.n685 10.6151
R1588 B.n685 B.n109 10.6151
R1589 B.n679 B.n109 10.6151
R1590 B.n679 B.n678 10.6151
R1591 B.n678 B.n677 10.6151
R1592 B.n677 B.n116 10.6151
R1593 B.n141 B.n140 10.6151
R1594 B.n144 B.n141 10.6151
R1595 B.n145 B.n144 10.6151
R1596 B.n148 B.n145 10.6151
R1597 B.n149 B.n148 10.6151
R1598 B.n152 B.n149 10.6151
R1599 B.n153 B.n152 10.6151
R1600 B.n156 B.n153 10.6151
R1601 B.n161 B.n158 10.6151
R1602 B.n162 B.n161 10.6151
R1603 B.n165 B.n162 10.6151
R1604 B.n166 B.n165 10.6151
R1605 B.n169 B.n166 10.6151
R1606 B.n170 B.n169 10.6151
R1607 B.n173 B.n170 10.6151
R1608 B.n174 B.n173 10.6151
R1609 B.n178 B.n177 10.6151
R1610 B.n181 B.n178 10.6151
R1611 B.n182 B.n181 10.6151
R1612 B.n185 B.n182 10.6151
R1613 B.n186 B.n185 10.6151
R1614 B.n189 B.n186 10.6151
R1615 B.n190 B.n189 10.6151
R1616 B.n671 B.n190 10.6151
R1617 B.n807 B.n0 8.11757
R1618 B.n807 B.n1 8.11757
R1619 B.n368 B.n334 6.5566
R1620 B.n352 B.n351 6.5566
R1621 B.n158 B.n157 6.5566
R1622 B.n174 B.n136 6.5566
R1623 B.n371 B.n334 4.05904
R1624 B.n351 B.n350 4.05904
R1625 B.n157 B.n156 4.05904
R1626 B.n177 B.n136 4.05904
R1627 VN.n72 VN.n71 161.3
R1628 VN.n70 VN.n38 161.3
R1629 VN.n69 VN.n68 161.3
R1630 VN.n67 VN.n39 161.3
R1631 VN.n66 VN.n65 161.3
R1632 VN.n64 VN.n40 161.3
R1633 VN.n63 VN.n62 161.3
R1634 VN.n61 VN.n41 161.3
R1635 VN.n60 VN.n59 161.3
R1636 VN.n58 VN.n42 161.3
R1637 VN.n57 VN.n56 161.3
R1638 VN.n55 VN.n44 161.3
R1639 VN.n54 VN.n53 161.3
R1640 VN.n52 VN.n45 161.3
R1641 VN.n51 VN.n50 161.3
R1642 VN.n49 VN.n46 161.3
R1643 VN.n35 VN.n34 161.3
R1644 VN.n33 VN.n1 161.3
R1645 VN.n32 VN.n31 161.3
R1646 VN.n30 VN.n2 161.3
R1647 VN.n29 VN.n28 161.3
R1648 VN.n27 VN.n3 161.3
R1649 VN.n26 VN.n25 161.3
R1650 VN.n24 VN.n4 161.3
R1651 VN.n23 VN.n22 161.3
R1652 VN.n20 VN.n5 161.3
R1653 VN.n19 VN.n18 161.3
R1654 VN.n17 VN.n6 161.3
R1655 VN.n16 VN.n15 161.3
R1656 VN.n14 VN.n7 161.3
R1657 VN.n13 VN.n12 161.3
R1658 VN.n11 VN.n8 161.3
R1659 VN.n36 VN.n0 85.908
R1660 VN.n73 VN.n37 85.908
R1661 VN.n10 VN.n9 65.0012
R1662 VN.n48 VN.n47 65.0012
R1663 VN.n15 VN.n6 56.5193
R1664 VN.n53 VN.n44 56.5193
R1665 VN.n28 VN.n2 54.0911
R1666 VN.n65 VN.n39 54.0911
R1667 VN VN.n73 47.0738
R1668 VN.n10 VN.t5 37.5796
R1669 VN.n48 VN.t4 37.5796
R1670 VN.n28 VN.n27 26.8957
R1671 VN.n65 VN.n64 26.8957
R1672 VN.n13 VN.n8 24.4675
R1673 VN.n14 VN.n13 24.4675
R1674 VN.n15 VN.n14 24.4675
R1675 VN.n19 VN.n6 24.4675
R1676 VN.n20 VN.n19 24.4675
R1677 VN.n22 VN.n20 24.4675
R1678 VN.n26 VN.n4 24.4675
R1679 VN.n27 VN.n26 24.4675
R1680 VN.n32 VN.n2 24.4675
R1681 VN.n33 VN.n32 24.4675
R1682 VN.n34 VN.n33 24.4675
R1683 VN.n53 VN.n52 24.4675
R1684 VN.n52 VN.n51 24.4675
R1685 VN.n51 VN.n46 24.4675
R1686 VN.n64 VN.n63 24.4675
R1687 VN.n63 VN.n41 24.4675
R1688 VN.n59 VN.n58 24.4675
R1689 VN.n58 VN.n57 24.4675
R1690 VN.n57 VN.n44 24.4675
R1691 VN.n71 VN.n70 24.4675
R1692 VN.n70 VN.n69 24.4675
R1693 VN.n69 VN.n39 24.4675
R1694 VN.n21 VN.n4 14.9254
R1695 VN.n43 VN.n41 14.9254
R1696 VN.n9 VN.n8 9.54263
R1697 VN.n22 VN.n21 9.54263
R1698 VN.n47 VN.n46 9.54263
R1699 VN.n59 VN.n43 9.54263
R1700 VN.n9 VN.t7 5.34853
R1701 VN.n21 VN.t1 5.34853
R1702 VN.n0 VN.t6 5.34853
R1703 VN.n47 VN.t2 5.34853
R1704 VN.n43 VN.t0 5.34853
R1705 VN.n37 VN.t3 5.34853
R1706 VN.n34 VN.n0 4.15989
R1707 VN.n71 VN.n37 4.15989
R1708 VN.n11 VN.n10 3.34374
R1709 VN.n49 VN.n48 3.34374
R1710 VN.n73 VN.n72 0.354971
R1711 VN.n36 VN.n35 0.354971
R1712 VN VN.n36 0.26696
R1713 VN.n72 VN.n38 0.189894
R1714 VN.n68 VN.n38 0.189894
R1715 VN.n68 VN.n67 0.189894
R1716 VN.n67 VN.n66 0.189894
R1717 VN.n66 VN.n40 0.189894
R1718 VN.n62 VN.n40 0.189894
R1719 VN.n62 VN.n61 0.189894
R1720 VN.n61 VN.n60 0.189894
R1721 VN.n60 VN.n42 0.189894
R1722 VN.n56 VN.n42 0.189894
R1723 VN.n56 VN.n55 0.189894
R1724 VN.n55 VN.n54 0.189894
R1725 VN.n54 VN.n45 0.189894
R1726 VN.n50 VN.n45 0.189894
R1727 VN.n50 VN.n49 0.189894
R1728 VN.n12 VN.n11 0.189894
R1729 VN.n12 VN.n7 0.189894
R1730 VN.n16 VN.n7 0.189894
R1731 VN.n17 VN.n16 0.189894
R1732 VN.n18 VN.n17 0.189894
R1733 VN.n18 VN.n5 0.189894
R1734 VN.n23 VN.n5 0.189894
R1735 VN.n24 VN.n23 0.189894
R1736 VN.n25 VN.n24 0.189894
R1737 VN.n25 VN.n3 0.189894
R1738 VN.n29 VN.n3 0.189894
R1739 VN.n30 VN.n29 0.189894
R1740 VN.n31 VN.n30 0.189894
R1741 VN.n31 VN.n1 0.189894
R1742 VN.n35 VN.n1 0.189894
R1743 VDD2.n2 VDD2.n1 239.171
R1744 VDD2.n2 VDD2.n0 239.171
R1745 VDD2 VDD2.n5 239.167
R1746 VDD2.n4 VDD2.n3 237.548
R1747 VDD2.n4 VDD2.n2 39.4868
R1748 VDD2.n5 VDD2.t5 25.0638
R1749 VDD2.n5 VDD2.t3 25.0638
R1750 VDD2.n3 VDD2.t4 25.0638
R1751 VDD2.n3 VDD2.t7 25.0638
R1752 VDD2.n1 VDD2.t6 25.0638
R1753 VDD2.n1 VDD2.t1 25.0638
R1754 VDD2.n0 VDD2.t2 25.0638
R1755 VDD2.n0 VDD2.t0 25.0638
R1756 VDD2 VDD2.n4 1.73541
C0 VDD1 VN 0.160967f
C1 VDD2 VP 0.631884f
C2 VDD1 VTAIL 5.25153f
C3 VDD2 VN 1.05921f
C4 VDD2 VTAIL 5.31238f
C5 VDD2 VDD1 2.27535f
C6 VN VP 6.77436f
C7 VTAIL VP 2.8718f
C8 VDD1 VP 1.52494f
C9 VTAIL VN 2.85769f
C10 VDD2 B 5.451074f
C11 VDD1 B 5.970287f
C12 VTAIL B 3.804905f
C13 VN B 18.49316f
C14 VP B 16.789736f
C15 VDD2.t2 B 0.019167f
C16 VDD2.t0 B 0.019167f
C17 VDD2.n0 B 0.050282f
C18 VDD2.t6 B 0.019167f
C19 VDD2.t1 B 0.019167f
C20 VDD2.n1 B 0.050282f
C21 VDD2.n2 B 3.54469f
C22 VDD2.t4 B 0.019167f
C23 VDD2.t7 B 0.019167f
C24 VDD2.n3 B 0.04632f
C25 VDD2.n4 B 2.79333f
C26 VDD2.t5 B 0.019167f
C27 VDD2.t3 B 0.019167f
C28 VDD2.n5 B 0.05027f
C29 VN.t6 B 0.13648f
C30 VN.n0 B 0.213918f
C31 VN.n1 B 0.029956f
C32 VN.n2 B 0.052506f
C33 VN.n3 B 0.029956f
C34 VN.n4 B 0.045079f
C35 VN.n5 B 0.029956f
C36 VN.n6 B 0.04373f
C37 VN.n7 B 0.029956f
C38 VN.n8 B 0.039015f
C39 VN.t7 B 0.13648f
C40 VN.n9 B 0.206974f
C41 VN.t5 B 0.419484f
C42 VN.n10 B 0.275789f
C43 VN.n11 B 0.374762f
C44 VN.n12 B 0.029956f
C45 VN.n13 B 0.05583f
C46 VN.n14 B 0.05583f
C47 VN.n15 B 0.04373f
C48 VN.n16 B 0.029956f
C49 VN.n17 B 0.029956f
C50 VN.n18 B 0.029956f
C51 VN.n19 B 0.05583f
C52 VN.n20 B 0.05583f
C53 VN.t1 B 0.13648f
C54 VN.n21 B 0.106261f
C55 VN.n22 B 0.039015f
C56 VN.n23 B 0.029956f
C57 VN.n24 B 0.029956f
C58 VN.n25 B 0.029956f
C59 VN.n26 B 0.05583f
C60 VN.n27 B 0.058068f
C61 VN.n28 B 0.032715f
C62 VN.n29 B 0.029956f
C63 VN.n30 B 0.029956f
C64 VN.n31 B 0.029956f
C65 VN.n32 B 0.05583f
C66 VN.n33 B 0.05583f
C67 VN.n34 B 0.032951f
C68 VN.n35 B 0.048348f
C69 VN.n36 B 0.086958f
C70 VN.t3 B 0.13648f
C71 VN.n37 B 0.213918f
C72 VN.n38 B 0.029956f
C73 VN.n39 B 0.052506f
C74 VN.n40 B 0.029956f
C75 VN.n41 B 0.045079f
C76 VN.n42 B 0.029956f
C77 VN.t0 B 0.13648f
C78 VN.n43 B 0.106261f
C79 VN.n44 B 0.04373f
C80 VN.n45 B 0.029956f
C81 VN.n46 B 0.039015f
C82 VN.t4 B 0.419484f
C83 VN.t2 B 0.13648f
C84 VN.n47 B 0.206974f
C85 VN.n48 B 0.275789f
C86 VN.n49 B 0.374762f
C87 VN.n50 B 0.029956f
C88 VN.n51 B 0.05583f
C89 VN.n52 B 0.05583f
C90 VN.n53 B 0.04373f
C91 VN.n54 B 0.029956f
C92 VN.n55 B 0.029956f
C93 VN.n56 B 0.029956f
C94 VN.n57 B 0.05583f
C95 VN.n58 B 0.05583f
C96 VN.n59 B 0.039015f
C97 VN.n60 B 0.029956f
C98 VN.n61 B 0.029956f
C99 VN.n62 B 0.029956f
C100 VN.n63 B 0.05583f
C101 VN.n64 B 0.058068f
C102 VN.n65 B 0.032715f
C103 VN.n66 B 0.029956f
C104 VN.n67 B 0.029956f
C105 VN.n68 B 0.029956f
C106 VN.n69 B 0.05583f
C107 VN.n70 B 0.05583f
C108 VN.n71 B 0.032951f
C109 VN.n72 B 0.048348f
C110 VN.n73 B 1.57803f
C111 VDD1.t2 B 0.018885f
C112 VDD1.t5 B 0.018885f
C113 VDD1.n0 B 0.049891f
C114 VDD1.t0 B 0.018885f
C115 VDD1.t3 B 0.018885f
C116 VDD1.n1 B 0.049543f
C117 VDD1.t4 B 0.018885f
C118 VDD1.t6 B 0.018885f
C119 VDD1.n2 B 0.049543f
C120 VDD1.n3 B 3.55521f
C121 VDD1.t1 B 0.018885f
C122 VDD1.t7 B 0.018885f
C123 VDD1.n4 B 0.045639f
C124 VDD1.n5 B 2.79001f
C125 VTAIL.t10 B 0.030404f
C126 VTAIL.t0 B 0.030404f
C127 VTAIL.n0 B 0.064662f
C128 VTAIL.n1 B 0.604016f
C129 VTAIL.t12 B 0.135641f
C130 VTAIL.n2 B 0.680557f
C131 VTAIL.t4 B 0.135641f
C132 VTAIL.n3 B 0.680557f
C133 VTAIL.t5 B 0.030404f
C134 VTAIL.t3 B 0.030404f
C135 VTAIL.n4 B 0.064662f
C136 VTAIL.n5 B 1.12115f
C137 VTAIL.t8 B 0.135641f
C138 VTAIL.n6 B 1.90154f
C139 VTAIL.t15 B 0.135641f
C140 VTAIL.n7 B 1.90154f
C141 VTAIL.t1 B 0.030404f
C142 VTAIL.t13 B 0.030404f
C143 VTAIL.n8 B 0.064662f
C144 VTAIL.n9 B 1.12115f
C145 VTAIL.t14 B 0.135641f
C146 VTAIL.n10 B 0.680557f
C147 VTAIL.t2 B 0.135641f
C148 VTAIL.n11 B 0.680557f
C149 VTAIL.t6 B 0.030404f
C150 VTAIL.t9 B 0.030404f
C151 VTAIL.n12 B 0.064662f
C152 VTAIL.n13 B 1.12115f
C153 VTAIL.t7 B 0.135641f
C154 VTAIL.n14 B 1.90154f
C155 VTAIL.t11 B 0.135641f
C156 VTAIL.n15 B 1.89241f
C157 VP.t1 B 0.137075f
C158 VP.n0 B 0.214851f
C159 VP.n1 B 0.030086f
C160 VP.n2 B 0.052735f
C161 VP.n3 B 0.030086f
C162 VP.n4 B 0.045275f
C163 VP.n5 B 0.030086f
C164 VP.n6 B 0.043921f
C165 VP.n7 B 0.030086f
C166 VP.n8 B 0.039185f
C167 VP.n9 B 0.030086f
C168 VP.n10 B 0.032858f
C169 VP.n11 B 0.030086f
C170 VP.n12 B 0.033094f
C171 VP.t0 B 0.137075f
C172 VP.n13 B 0.214851f
C173 VP.n14 B 0.030086f
C174 VP.n15 B 0.052735f
C175 VP.n16 B 0.030086f
C176 VP.n17 B 0.045275f
C177 VP.n18 B 0.030086f
C178 VP.n19 B 0.043921f
C179 VP.n20 B 0.030086f
C180 VP.n21 B 0.039185f
C181 VP.t5 B 0.421312f
C182 VP.t2 B 0.137075f
C183 VP.n22 B 0.207877f
C184 VP.n23 B 0.276992f
C185 VP.n24 B 0.376397f
C186 VP.n25 B 0.030086f
C187 VP.n26 B 0.056073f
C188 VP.n27 B 0.056073f
C189 VP.n28 B 0.043921f
C190 VP.n29 B 0.030086f
C191 VP.n30 B 0.030086f
C192 VP.n31 B 0.030086f
C193 VP.n32 B 0.056073f
C194 VP.n33 B 0.056073f
C195 VP.t6 B 0.137075f
C196 VP.n34 B 0.106724f
C197 VP.n35 B 0.039185f
C198 VP.n36 B 0.030086f
C199 VP.n37 B 0.030086f
C200 VP.n38 B 0.030086f
C201 VP.n39 B 0.056073f
C202 VP.n40 B 0.058321f
C203 VP.n41 B 0.032858f
C204 VP.n42 B 0.030086f
C205 VP.n43 B 0.030086f
C206 VP.n44 B 0.030086f
C207 VP.n45 B 0.056073f
C208 VP.n46 B 0.056073f
C209 VP.n47 B 0.033094f
C210 VP.n48 B 0.048559f
C211 VP.n49 B 1.57232f
C212 VP.t7 B 0.137075f
C213 VP.n50 B 0.214851f
C214 VP.n51 B 1.59537f
C215 VP.n52 B 0.048559f
C216 VP.n53 B 0.030086f
C217 VP.n54 B 0.056073f
C218 VP.n55 B 0.056073f
C219 VP.n56 B 0.052735f
C220 VP.n57 B 0.030086f
C221 VP.n58 B 0.030086f
C222 VP.n59 B 0.030086f
C223 VP.n60 B 0.058321f
C224 VP.n61 B 0.056073f
C225 VP.t4 B 0.137075f
C226 VP.n62 B 0.106724f
C227 VP.n63 B 0.045275f
C228 VP.n64 B 0.030086f
C229 VP.n65 B 0.030086f
C230 VP.n66 B 0.030086f
C231 VP.n67 B 0.056073f
C232 VP.n68 B 0.056073f
C233 VP.n69 B 0.043921f
C234 VP.n70 B 0.030086f
C235 VP.n71 B 0.030086f
C236 VP.n72 B 0.030086f
C237 VP.n73 B 0.056073f
C238 VP.n74 B 0.056073f
C239 VP.t3 B 0.137075f
C240 VP.n75 B 0.106724f
C241 VP.n76 B 0.039185f
C242 VP.n77 B 0.030086f
C243 VP.n78 B 0.030086f
C244 VP.n79 B 0.030086f
C245 VP.n80 B 0.056073f
C246 VP.n81 B 0.058321f
C247 VP.n82 B 0.032858f
C248 VP.n83 B 0.030086f
C249 VP.n84 B 0.030086f
C250 VP.n85 B 0.030086f
C251 VP.n86 B 0.056073f
C252 VP.n87 B 0.056073f
C253 VP.n88 B 0.033094f
C254 VP.n89 B 0.048559f
C255 VP.n90 B 0.087338f
.ends

