* NGSPICE file created from diff_pair_sample_1782.ext - technology: sky130A

.subckt diff_pair_sample_1782 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t2 w_n1642_n4174# sky130_fd_pr__pfet_01v8 ad=6.2517 pd=32.84 as=2.64495 ps=16.36 w=16.03 l=0.79
X1 B.t11 B.t9 B.t10 w_n1642_n4174# sky130_fd_pr__pfet_01v8 ad=6.2517 pd=32.84 as=0 ps=0 w=16.03 l=0.79
X2 VTAIL.t2 VP.t0 VDD1.t3 w_n1642_n4174# sky130_fd_pr__pfet_01v8 ad=6.2517 pd=32.84 as=2.64495 ps=16.36 w=16.03 l=0.79
X3 VDD2.t1 VN.t1 VTAIL.t6 w_n1642_n4174# sky130_fd_pr__pfet_01v8 ad=2.64495 pd=16.36 as=6.2517 ps=32.84 w=16.03 l=0.79
X4 B.t8 B.t6 B.t7 w_n1642_n4174# sky130_fd_pr__pfet_01v8 ad=6.2517 pd=32.84 as=0 ps=0 w=16.03 l=0.79
X5 VDD1.t2 VP.t1 VTAIL.t3 w_n1642_n4174# sky130_fd_pr__pfet_01v8 ad=2.64495 pd=16.36 as=6.2517 ps=32.84 w=16.03 l=0.79
X6 VDD2.t0 VN.t2 VTAIL.t5 w_n1642_n4174# sky130_fd_pr__pfet_01v8 ad=2.64495 pd=16.36 as=6.2517 ps=32.84 w=16.03 l=0.79
X7 B.t5 B.t3 B.t4 w_n1642_n4174# sky130_fd_pr__pfet_01v8 ad=6.2517 pd=32.84 as=0 ps=0 w=16.03 l=0.79
X8 VTAIL.t0 VP.t2 VDD1.t1 w_n1642_n4174# sky130_fd_pr__pfet_01v8 ad=6.2517 pd=32.84 as=2.64495 ps=16.36 w=16.03 l=0.79
X9 B.t2 B.t0 B.t1 w_n1642_n4174# sky130_fd_pr__pfet_01v8 ad=6.2517 pd=32.84 as=0 ps=0 w=16.03 l=0.79
X10 VTAIL.t4 VN.t3 VDD2.t3 w_n1642_n4174# sky130_fd_pr__pfet_01v8 ad=6.2517 pd=32.84 as=2.64495 ps=16.36 w=16.03 l=0.79
X11 VDD1.t0 VP.t3 VTAIL.t1 w_n1642_n4174# sky130_fd_pr__pfet_01v8 ad=2.64495 pd=16.36 as=6.2517 ps=32.84 w=16.03 l=0.79
R0 VN.n0 VN.t3 560.043
R1 VN.n1 VN.t2 560.043
R2 VN.n0 VN.t1 559.994
R3 VN.n1 VN.t0 559.994
R4 VN VN.n1 88.8458
R5 VN VN.n0 44.7132
R6 VDD2.n2 VDD2.n0 109.263
R7 VDD2.n2 VDD2.n1 68.8322
R8 VDD2.n1 VDD2.t2 2.02826
R9 VDD2.n1 VDD2.t0 2.02826
R10 VDD2.n0 VDD2.t3 2.02826
R11 VDD2.n0 VDD2.t1 2.02826
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n714 VTAIL.n630 756.745
R14 VTAIL.n84 VTAIL.n0 756.745
R15 VTAIL.n174 VTAIL.n90 756.745
R16 VTAIL.n264 VTAIL.n180 756.745
R17 VTAIL.n624 VTAIL.n540 756.745
R18 VTAIL.n534 VTAIL.n450 756.745
R19 VTAIL.n444 VTAIL.n360 756.745
R20 VTAIL.n354 VTAIL.n270 756.745
R21 VTAIL.n658 VTAIL.n657 585
R22 VTAIL.n663 VTAIL.n662 585
R23 VTAIL.n665 VTAIL.n664 585
R24 VTAIL.n654 VTAIL.n653 585
R25 VTAIL.n671 VTAIL.n670 585
R26 VTAIL.n673 VTAIL.n672 585
R27 VTAIL.n650 VTAIL.n649 585
R28 VTAIL.n679 VTAIL.n678 585
R29 VTAIL.n681 VTAIL.n680 585
R30 VTAIL.n646 VTAIL.n645 585
R31 VTAIL.n687 VTAIL.n686 585
R32 VTAIL.n689 VTAIL.n688 585
R33 VTAIL.n642 VTAIL.n641 585
R34 VTAIL.n695 VTAIL.n694 585
R35 VTAIL.n697 VTAIL.n696 585
R36 VTAIL.n638 VTAIL.n637 585
R37 VTAIL.n704 VTAIL.n703 585
R38 VTAIL.n705 VTAIL.n636 585
R39 VTAIL.n707 VTAIL.n706 585
R40 VTAIL.n634 VTAIL.n633 585
R41 VTAIL.n713 VTAIL.n712 585
R42 VTAIL.n715 VTAIL.n714 585
R43 VTAIL.n28 VTAIL.n27 585
R44 VTAIL.n33 VTAIL.n32 585
R45 VTAIL.n35 VTAIL.n34 585
R46 VTAIL.n24 VTAIL.n23 585
R47 VTAIL.n41 VTAIL.n40 585
R48 VTAIL.n43 VTAIL.n42 585
R49 VTAIL.n20 VTAIL.n19 585
R50 VTAIL.n49 VTAIL.n48 585
R51 VTAIL.n51 VTAIL.n50 585
R52 VTAIL.n16 VTAIL.n15 585
R53 VTAIL.n57 VTAIL.n56 585
R54 VTAIL.n59 VTAIL.n58 585
R55 VTAIL.n12 VTAIL.n11 585
R56 VTAIL.n65 VTAIL.n64 585
R57 VTAIL.n67 VTAIL.n66 585
R58 VTAIL.n8 VTAIL.n7 585
R59 VTAIL.n74 VTAIL.n73 585
R60 VTAIL.n75 VTAIL.n6 585
R61 VTAIL.n77 VTAIL.n76 585
R62 VTAIL.n4 VTAIL.n3 585
R63 VTAIL.n83 VTAIL.n82 585
R64 VTAIL.n85 VTAIL.n84 585
R65 VTAIL.n118 VTAIL.n117 585
R66 VTAIL.n123 VTAIL.n122 585
R67 VTAIL.n125 VTAIL.n124 585
R68 VTAIL.n114 VTAIL.n113 585
R69 VTAIL.n131 VTAIL.n130 585
R70 VTAIL.n133 VTAIL.n132 585
R71 VTAIL.n110 VTAIL.n109 585
R72 VTAIL.n139 VTAIL.n138 585
R73 VTAIL.n141 VTAIL.n140 585
R74 VTAIL.n106 VTAIL.n105 585
R75 VTAIL.n147 VTAIL.n146 585
R76 VTAIL.n149 VTAIL.n148 585
R77 VTAIL.n102 VTAIL.n101 585
R78 VTAIL.n155 VTAIL.n154 585
R79 VTAIL.n157 VTAIL.n156 585
R80 VTAIL.n98 VTAIL.n97 585
R81 VTAIL.n164 VTAIL.n163 585
R82 VTAIL.n165 VTAIL.n96 585
R83 VTAIL.n167 VTAIL.n166 585
R84 VTAIL.n94 VTAIL.n93 585
R85 VTAIL.n173 VTAIL.n172 585
R86 VTAIL.n175 VTAIL.n174 585
R87 VTAIL.n208 VTAIL.n207 585
R88 VTAIL.n213 VTAIL.n212 585
R89 VTAIL.n215 VTAIL.n214 585
R90 VTAIL.n204 VTAIL.n203 585
R91 VTAIL.n221 VTAIL.n220 585
R92 VTAIL.n223 VTAIL.n222 585
R93 VTAIL.n200 VTAIL.n199 585
R94 VTAIL.n229 VTAIL.n228 585
R95 VTAIL.n231 VTAIL.n230 585
R96 VTAIL.n196 VTAIL.n195 585
R97 VTAIL.n237 VTAIL.n236 585
R98 VTAIL.n239 VTAIL.n238 585
R99 VTAIL.n192 VTAIL.n191 585
R100 VTAIL.n245 VTAIL.n244 585
R101 VTAIL.n247 VTAIL.n246 585
R102 VTAIL.n188 VTAIL.n187 585
R103 VTAIL.n254 VTAIL.n253 585
R104 VTAIL.n255 VTAIL.n186 585
R105 VTAIL.n257 VTAIL.n256 585
R106 VTAIL.n184 VTAIL.n183 585
R107 VTAIL.n263 VTAIL.n262 585
R108 VTAIL.n265 VTAIL.n264 585
R109 VTAIL.n625 VTAIL.n624 585
R110 VTAIL.n623 VTAIL.n622 585
R111 VTAIL.n544 VTAIL.n543 585
R112 VTAIL.n617 VTAIL.n616 585
R113 VTAIL.n615 VTAIL.n546 585
R114 VTAIL.n614 VTAIL.n613 585
R115 VTAIL.n549 VTAIL.n547 585
R116 VTAIL.n608 VTAIL.n607 585
R117 VTAIL.n606 VTAIL.n605 585
R118 VTAIL.n553 VTAIL.n552 585
R119 VTAIL.n600 VTAIL.n599 585
R120 VTAIL.n598 VTAIL.n597 585
R121 VTAIL.n557 VTAIL.n556 585
R122 VTAIL.n592 VTAIL.n591 585
R123 VTAIL.n590 VTAIL.n589 585
R124 VTAIL.n561 VTAIL.n560 585
R125 VTAIL.n584 VTAIL.n583 585
R126 VTAIL.n582 VTAIL.n581 585
R127 VTAIL.n565 VTAIL.n564 585
R128 VTAIL.n576 VTAIL.n575 585
R129 VTAIL.n574 VTAIL.n573 585
R130 VTAIL.n569 VTAIL.n568 585
R131 VTAIL.n535 VTAIL.n534 585
R132 VTAIL.n533 VTAIL.n532 585
R133 VTAIL.n454 VTAIL.n453 585
R134 VTAIL.n527 VTAIL.n526 585
R135 VTAIL.n525 VTAIL.n456 585
R136 VTAIL.n524 VTAIL.n523 585
R137 VTAIL.n459 VTAIL.n457 585
R138 VTAIL.n518 VTAIL.n517 585
R139 VTAIL.n516 VTAIL.n515 585
R140 VTAIL.n463 VTAIL.n462 585
R141 VTAIL.n510 VTAIL.n509 585
R142 VTAIL.n508 VTAIL.n507 585
R143 VTAIL.n467 VTAIL.n466 585
R144 VTAIL.n502 VTAIL.n501 585
R145 VTAIL.n500 VTAIL.n499 585
R146 VTAIL.n471 VTAIL.n470 585
R147 VTAIL.n494 VTAIL.n493 585
R148 VTAIL.n492 VTAIL.n491 585
R149 VTAIL.n475 VTAIL.n474 585
R150 VTAIL.n486 VTAIL.n485 585
R151 VTAIL.n484 VTAIL.n483 585
R152 VTAIL.n479 VTAIL.n478 585
R153 VTAIL.n445 VTAIL.n444 585
R154 VTAIL.n443 VTAIL.n442 585
R155 VTAIL.n364 VTAIL.n363 585
R156 VTAIL.n437 VTAIL.n436 585
R157 VTAIL.n435 VTAIL.n366 585
R158 VTAIL.n434 VTAIL.n433 585
R159 VTAIL.n369 VTAIL.n367 585
R160 VTAIL.n428 VTAIL.n427 585
R161 VTAIL.n426 VTAIL.n425 585
R162 VTAIL.n373 VTAIL.n372 585
R163 VTAIL.n420 VTAIL.n419 585
R164 VTAIL.n418 VTAIL.n417 585
R165 VTAIL.n377 VTAIL.n376 585
R166 VTAIL.n412 VTAIL.n411 585
R167 VTAIL.n410 VTAIL.n409 585
R168 VTAIL.n381 VTAIL.n380 585
R169 VTAIL.n404 VTAIL.n403 585
R170 VTAIL.n402 VTAIL.n401 585
R171 VTAIL.n385 VTAIL.n384 585
R172 VTAIL.n396 VTAIL.n395 585
R173 VTAIL.n394 VTAIL.n393 585
R174 VTAIL.n389 VTAIL.n388 585
R175 VTAIL.n355 VTAIL.n354 585
R176 VTAIL.n353 VTAIL.n352 585
R177 VTAIL.n274 VTAIL.n273 585
R178 VTAIL.n347 VTAIL.n346 585
R179 VTAIL.n345 VTAIL.n276 585
R180 VTAIL.n344 VTAIL.n343 585
R181 VTAIL.n279 VTAIL.n277 585
R182 VTAIL.n338 VTAIL.n337 585
R183 VTAIL.n336 VTAIL.n335 585
R184 VTAIL.n283 VTAIL.n282 585
R185 VTAIL.n330 VTAIL.n329 585
R186 VTAIL.n328 VTAIL.n327 585
R187 VTAIL.n287 VTAIL.n286 585
R188 VTAIL.n322 VTAIL.n321 585
R189 VTAIL.n320 VTAIL.n319 585
R190 VTAIL.n291 VTAIL.n290 585
R191 VTAIL.n314 VTAIL.n313 585
R192 VTAIL.n312 VTAIL.n311 585
R193 VTAIL.n295 VTAIL.n294 585
R194 VTAIL.n306 VTAIL.n305 585
R195 VTAIL.n304 VTAIL.n303 585
R196 VTAIL.n299 VTAIL.n298 585
R197 VTAIL.n659 VTAIL.t6 327.466
R198 VTAIL.n29 VTAIL.t4 327.466
R199 VTAIL.n119 VTAIL.t3 327.466
R200 VTAIL.n209 VTAIL.t0 327.466
R201 VTAIL.n570 VTAIL.t1 327.466
R202 VTAIL.n480 VTAIL.t2 327.466
R203 VTAIL.n390 VTAIL.t5 327.466
R204 VTAIL.n300 VTAIL.t7 327.466
R205 VTAIL.n663 VTAIL.n657 171.744
R206 VTAIL.n664 VTAIL.n663 171.744
R207 VTAIL.n664 VTAIL.n653 171.744
R208 VTAIL.n671 VTAIL.n653 171.744
R209 VTAIL.n672 VTAIL.n671 171.744
R210 VTAIL.n672 VTAIL.n649 171.744
R211 VTAIL.n679 VTAIL.n649 171.744
R212 VTAIL.n680 VTAIL.n679 171.744
R213 VTAIL.n680 VTAIL.n645 171.744
R214 VTAIL.n687 VTAIL.n645 171.744
R215 VTAIL.n688 VTAIL.n687 171.744
R216 VTAIL.n688 VTAIL.n641 171.744
R217 VTAIL.n695 VTAIL.n641 171.744
R218 VTAIL.n696 VTAIL.n695 171.744
R219 VTAIL.n696 VTAIL.n637 171.744
R220 VTAIL.n704 VTAIL.n637 171.744
R221 VTAIL.n705 VTAIL.n704 171.744
R222 VTAIL.n706 VTAIL.n705 171.744
R223 VTAIL.n706 VTAIL.n633 171.744
R224 VTAIL.n713 VTAIL.n633 171.744
R225 VTAIL.n714 VTAIL.n713 171.744
R226 VTAIL.n33 VTAIL.n27 171.744
R227 VTAIL.n34 VTAIL.n33 171.744
R228 VTAIL.n34 VTAIL.n23 171.744
R229 VTAIL.n41 VTAIL.n23 171.744
R230 VTAIL.n42 VTAIL.n41 171.744
R231 VTAIL.n42 VTAIL.n19 171.744
R232 VTAIL.n49 VTAIL.n19 171.744
R233 VTAIL.n50 VTAIL.n49 171.744
R234 VTAIL.n50 VTAIL.n15 171.744
R235 VTAIL.n57 VTAIL.n15 171.744
R236 VTAIL.n58 VTAIL.n57 171.744
R237 VTAIL.n58 VTAIL.n11 171.744
R238 VTAIL.n65 VTAIL.n11 171.744
R239 VTAIL.n66 VTAIL.n65 171.744
R240 VTAIL.n66 VTAIL.n7 171.744
R241 VTAIL.n74 VTAIL.n7 171.744
R242 VTAIL.n75 VTAIL.n74 171.744
R243 VTAIL.n76 VTAIL.n75 171.744
R244 VTAIL.n76 VTAIL.n3 171.744
R245 VTAIL.n83 VTAIL.n3 171.744
R246 VTAIL.n84 VTAIL.n83 171.744
R247 VTAIL.n123 VTAIL.n117 171.744
R248 VTAIL.n124 VTAIL.n123 171.744
R249 VTAIL.n124 VTAIL.n113 171.744
R250 VTAIL.n131 VTAIL.n113 171.744
R251 VTAIL.n132 VTAIL.n131 171.744
R252 VTAIL.n132 VTAIL.n109 171.744
R253 VTAIL.n139 VTAIL.n109 171.744
R254 VTAIL.n140 VTAIL.n139 171.744
R255 VTAIL.n140 VTAIL.n105 171.744
R256 VTAIL.n147 VTAIL.n105 171.744
R257 VTAIL.n148 VTAIL.n147 171.744
R258 VTAIL.n148 VTAIL.n101 171.744
R259 VTAIL.n155 VTAIL.n101 171.744
R260 VTAIL.n156 VTAIL.n155 171.744
R261 VTAIL.n156 VTAIL.n97 171.744
R262 VTAIL.n164 VTAIL.n97 171.744
R263 VTAIL.n165 VTAIL.n164 171.744
R264 VTAIL.n166 VTAIL.n165 171.744
R265 VTAIL.n166 VTAIL.n93 171.744
R266 VTAIL.n173 VTAIL.n93 171.744
R267 VTAIL.n174 VTAIL.n173 171.744
R268 VTAIL.n213 VTAIL.n207 171.744
R269 VTAIL.n214 VTAIL.n213 171.744
R270 VTAIL.n214 VTAIL.n203 171.744
R271 VTAIL.n221 VTAIL.n203 171.744
R272 VTAIL.n222 VTAIL.n221 171.744
R273 VTAIL.n222 VTAIL.n199 171.744
R274 VTAIL.n229 VTAIL.n199 171.744
R275 VTAIL.n230 VTAIL.n229 171.744
R276 VTAIL.n230 VTAIL.n195 171.744
R277 VTAIL.n237 VTAIL.n195 171.744
R278 VTAIL.n238 VTAIL.n237 171.744
R279 VTAIL.n238 VTAIL.n191 171.744
R280 VTAIL.n245 VTAIL.n191 171.744
R281 VTAIL.n246 VTAIL.n245 171.744
R282 VTAIL.n246 VTAIL.n187 171.744
R283 VTAIL.n254 VTAIL.n187 171.744
R284 VTAIL.n255 VTAIL.n254 171.744
R285 VTAIL.n256 VTAIL.n255 171.744
R286 VTAIL.n256 VTAIL.n183 171.744
R287 VTAIL.n263 VTAIL.n183 171.744
R288 VTAIL.n264 VTAIL.n263 171.744
R289 VTAIL.n624 VTAIL.n623 171.744
R290 VTAIL.n623 VTAIL.n543 171.744
R291 VTAIL.n616 VTAIL.n543 171.744
R292 VTAIL.n616 VTAIL.n615 171.744
R293 VTAIL.n615 VTAIL.n614 171.744
R294 VTAIL.n614 VTAIL.n547 171.744
R295 VTAIL.n607 VTAIL.n547 171.744
R296 VTAIL.n607 VTAIL.n606 171.744
R297 VTAIL.n606 VTAIL.n552 171.744
R298 VTAIL.n599 VTAIL.n552 171.744
R299 VTAIL.n599 VTAIL.n598 171.744
R300 VTAIL.n598 VTAIL.n556 171.744
R301 VTAIL.n591 VTAIL.n556 171.744
R302 VTAIL.n591 VTAIL.n590 171.744
R303 VTAIL.n590 VTAIL.n560 171.744
R304 VTAIL.n583 VTAIL.n560 171.744
R305 VTAIL.n583 VTAIL.n582 171.744
R306 VTAIL.n582 VTAIL.n564 171.744
R307 VTAIL.n575 VTAIL.n564 171.744
R308 VTAIL.n575 VTAIL.n574 171.744
R309 VTAIL.n574 VTAIL.n568 171.744
R310 VTAIL.n534 VTAIL.n533 171.744
R311 VTAIL.n533 VTAIL.n453 171.744
R312 VTAIL.n526 VTAIL.n453 171.744
R313 VTAIL.n526 VTAIL.n525 171.744
R314 VTAIL.n525 VTAIL.n524 171.744
R315 VTAIL.n524 VTAIL.n457 171.744
R316 VTAIL.n517 VTAIL.n457 171.744
R317 VTAIL.n517 VTAIL.n516 171.744
R318 VTAIL.n516 VTAIL.n462 171.744
R319 VTAIL.n509 VTAIL.n462 171.744
R320 VTAIL.n509 VTAIL.n508 171.744
R321 VTAIL.n508 VTAIL.n466 171.744
R322 VTAIL.n501 VTAIL.n466 171.744
R323 VTAIL.n501 VTAIL.n500 171.744
R324 VTAIL.n500 VTAIL.n470 171.744
R325 VTAIL.n493 VTAIL.n470 171.744
R326 VTAIL.n493 VTAIL.n492 171.744
R327 VTAIL.n492 VTAIL.n474 171.744
R328 VTAIL.n485 VTAIL.n474 171.744
R329 VTAIL.n485 VTAIL.n484 171.744
R330 VTAIL.n484 VTAIL.n478 171.744
R331 VTAIL.n444 VTAIL.n443 171.744
R332 VTAIL.n443 VTAIL.n363 171.744
R333 VTAIL.n436 VTAIL.n363 171.744
R334 VTAIL.n436 VTAIL.n435 171.744
R335 VTAIL.n435 VTAIL.n434 171.744
R336 VTAIL.n434 VTAIL.n367 171.744
R337 VTAIL.n427 VTAIL.n367 171.744
R338 VTAIL.n427 VTAIL.n426 171.744
R339 VTAIL.n426 VTAIL.n372 171.744
R340 VTAIL.n419 VTAIL.n372 171.744
R341 VTAIL.n419 VTAIL.n418 171.744
R342 VTAIL.n418 VTAIL.n376 171.744
R343 VTAIL.n411 VTAIL.n376 171.744
R344 VTAIL.n411 VTAIL.n410 171.744
R345 VTAIL.n410 VTAIL.n380 171.744
R346 VTAIL.n403 VTAIL.n380 171.744
R347 VTAIL.n403 VTAIL.n402 171.744
R348 VTAIL.n402 VTAIL.n384 171.744
R349 VTAIL.n395 VTAIL.n384 171.744
R350 VTAIL.n395 VTAIL.n394 171.744
R351 VTAIL.n394 VTAIL.n388 171.744
R352 VTAIL.n354 VTAIL.n353 171.744
R353 VTAIL.n353 VTAIL.n273 171.744
R354 VTAIL.n346 VTAIL.n273 171.744
R355 VTAIL.n346 VTAIL.n345 171.744
R356 VTAIL.n345 VTAIL.n344 171.744
R357 VTAIL.n344 VTAIL.n277 171.744
R358 VTAIL.n337 VTAIL.n277 171.744
R359 VTAIL.n337 VTAIL.n336 171.744
R360 VTAIL.n336 VTAIL.n282 171.744
R361 VTAIL.n329 VTAIL.n282 171.744
R362 VTAIL.n329 VTAIL.n328 171.744
R363 VTAIL.n328 VTAIL.n286 171.744
R364 VTAIL.n321 VTAIL.n286 171.744
R365 VTAIL.n321 VTAIL.n320 171.744
R366 VTAIL.n320 VTAIL.n290 171.744
R367 VTAIL.n313 VTAIL.n290 171.744
R368 VTAIL.n313 VTAIL.n312 171.744
R369 VTAIL.n312 VTAIL.n294 171.744
R370 VTAIL.n305 VTAIL.n294 171.744
R371 VTAIL.n305 VTAIL.n304 171.744
R372 VTAIL.n304 VTAIL.n298 171.744
R373 VTAIL.t6 VTAIL.n657 85.8723
R374 VTAIL.t4 VTAIL.n27 85.8723
R375 VTAIL.t3 VTAIL.n117 85.8723
R376 VTAIL.t0 VTAIL.n207 85.8723
R377 VTAIL.t1 VTAIL.n568 85.8723
R378 VTAIL.t2 VTAIL.n478 85.8723
R379 VTAIL.t5 VTAIL.n388 85.8723
R380 VTAIL.t7 VTAIL.n298 85.8723
R381 VTAIL.n719 VTAIL.n718 31.2157
R382 VTAIL.n89 VTAIL.n88 31.2157
R383 VTAIL.n179 VTAIL.n178 31.2157
R384 VTAIL.n269 VTAIL.n268 31.2157
R385 VTAIL.n629 VTAIL.n628 31.2157
R386 VTAIL.n539 VTAIL.n538 31.2157
R387 VTAIL.n449 VTAIL.n448 31.2157
R388 VTAIL.n359 VTAIL.n358 31.2157
R389 VTAIL.n719 VTAIL.n629 27.1514
R390 VTAIL.n359 VTAIL.n269 27.1514
R391 VTAIL.n659 VTAIL.n658 16.3895
R392 VTAIL.n29 VTAIL.n28 16.3895
R393 VTAIL.n119 VTAIL.n118 16.3895
R394 VTAIL.n209 VTAIL.n208 16.3895
R395 VTAIL.n570 VTAIL.n569 16.3895
R396 VTAIL.n480 VTAIL.n479 16.3895
R397 VTAIL.n390 VTAIL.n389 16.3895
R398 VTAIL.n300 VTAIL.n299 16.3895
R399 VTAIL.n707 VTAIL.n636 13.1884
R400 VTAIL.n77 VTAIL.n6 13.1884
R401 VTAIL.n167 VTAIL.n96 13.1884
R402 VTAIL.n257 VTAIL.n186 13.1884
R403 VTAIL.n617 VTAIL.n546 13.1884
R404 VTAIL.n527 VTAIL.n456 13.1884
R405 VTAIL.n437 VTAIL.n366 13.1884
R406 VTAIL.n347 VTAIL.n276 13.1884
R407 VTAIL.n662 VTAIL.n661 12.8005
R408 VTAIL.n703 VTAIL.n702 12.8005
R409 VTAIL.n708 VTAIL.n634 12.8005
R410 VTAIL.n32 VTAIL.n31 12.8005
R411 VTAIL.n73 VTAIL.n72 12.8005
R412 VTAIL.n78 VTAIL.n4 12.8005
R413 VTAIL.n122 VTAIL.n121 12.8005
R414 VTAIL.n163 VTAIL.n162 12.8005
R415 VTAIL.n168 VTAIL.n94 12.8005
R416 VTAIL.n212 VTAIL.n211 12.8005
R417 VTAIL.n253 VTAIL.n252 12.8005
R418 VTAIL.n258 VTAIL.n184 12.8005
R419 VTAIL.n618 VTAIL.n544 12.8005
R420 VTAIL.n613 VTAIL.n548 12.8005
R421 VTAIL.n573 VTAIL.n572 12.8005
R422 VTAIL.n528 VTAIL.n454 12.8005
R423 VTAIL.n523 VTAIL.n458 12.8005
R424 VTAIL.n483 VTAIL.n482 12.8005
R425 VTAIL.n438 VTAIL.n364 12.8005
R426 VTAIL.n433 VTAIL.n368 12.8005
R427 VTAIL.n393 VTAIL.n392 12.8005
R428 VTAIL.n348 VTAIL.n274 12.8005
R429 VTAIL.n343 VTAIL.n278 12.8005
R430 VTAIL.n303 VTAIL.n302 12.8005
R431 VTAIL.n665 VTAIL.n656 12.0247
R432 VTAIL.n701 VTAIL.n638 12.0247
R433 VTAIL.n712 VTAIL.n711 12.0247
R434 VTAIL.n35 VTAIL.n26 12.0247
R435 VTAIL.n71 VTAIL.n8 12.0247
R436 VTAIL.n82 VTAIL.n81 12.0247
R437 VTAIL.n125 VTAIL.n116 12.0247
R438 VTAIL.n161 VTAIL.n98 12.0247
R439 VTAIL.n172 VTAIL.n171 12.0247
R440 VTAIL.n215 VTAIL.n206 12.0247
R441 VTAIL.n251 VTAIL.n188 12.0247
R442 VTAIL.n262 VTAIL.n261 12.0247
R443 VTAIL.n622 VTAIL.n621 12.0247
R444 VTAIL.n612 VTAIL.n549 12.0247
R445 VTAIL.n576 VTAIL.n567 12.0247
R446 VTAIL.n532 VTAIL.n531 12.0247
R447 VTAIL.n522 VTAIL.n459 12.0247
R448 VTAIL.n486 VTAIL.n477 12.0247
R449 VTAIL.n442 VTAIL.n441 12.0247
R450 VTAIL.n432 VTAIL.n369 12.0247
R451 VTAIL.n396 VTAIL.n387 12.0247
R452 VTAIL.n352 VTAIL.n351 12.0247
R453 VTAIL.n342 VTAIL.n279 12.0247
R454 VTAIL.n306 VTAIL.n297 12.0247
R455 VTAIL.n666 VTAIL.n654 11.249
R456 VTAIL.n698 VTAIL.n697 11.249
R457 VTAIL.n715 VTAIL.n632 11.249
R458 VTAIL.n36 VTAIL.n24 11.249
R459 VTAIL.n68 VTAIL.n67 11.249
R460 VTAIL.n85 VTAIL.n2 11.249
R461 VTAIL.n126 VTAIL.n114 11.249
R462 VTAIL.n158 VTAIL.n157 11.249
R463 VTAIL.n175 VTAIL.n92 11.249
R464 VTAIL.n216 VTAIL.n204 11.249
R465 VTAIL.n248 VTAIL.n247 11.249
R466 VTAIL.n265 VTAIL.n182 11.249
R467 VTAIL.n625 VTAIL.n542 11.249
R468 VTAIL.n609 VTAIL.n608 11.249
R469 VTAIL.n577 VTAIL.n565 11.249
R470 VTAIL.n535 VTAIL.n452 11.249
R471 VTAIL.n519 VTAIL.n518 11.249
R472 VTAIL.n487 VTAIL.n475 11.249
R473 VTAIL.n445 VTAIL.n362 11.249
R474 VTAIL.n429 VTAIL.n428 11.249
R475 VTAIL.n397 VTAIL.n385 11.249
R476 VTAIL.n355 VTAIL.n272 11.249
R477 VTAIL.n339 VTAIL.n338 11.249
R478 VTAIL.n307 VTAIL.n295 11.249
R479 VTAIL.n670 VTAIL.n669 10.4732
R480 VTAIL.n694 VTAIL.n640 10.4732
R481 VTAIL.n716 VTAIL.n630 10.4732
R482 VTAIL.n40 VTAIL.n39 10.4732
R483 VTAIL.n64 VTAIL.n10 10.4732
R484 VTAIL.n86 VTAIL.n0 10.4732
R485 VTAIL.n130 VTAIL.n129 10.4732
R486 VTAIL.n154 VTAIL.n100 10.4732
R487 VTAIL.n176 VTAIL.n90 10.4732
R488 VTAIL.n220 VTAIL.n219 10.4732
R489 VTAIL.n244 VTAIL.n190 10.4732
R490 VTAIL.n266 VTAIL.n180 10.4732
R491 VTAIL.n626 VTAIL.n540 10.4732
R492 VTAIL.n605 VTAIL.n551 10.4732
R493 VTAIL.n581 VTAIL.n580 10.4732
R494 VTAIL.n536 VTAIL.n450 10.4732
R495 VTAIL.n515 VTAIL.n461 10.4732
R496 VTAIL.n491 VTAIL.n490 10.4732
R497 VTAIL.n446 VTAIL.n360 10.4732
R498 VTAIL.n425 VTAIL.n371 10.4732
R499 VTAIL.n401 VTAIL.n400 10.4732
R500 VTAIL.n356 VTAIL.n270 10.4732
R501 VTAIL.n335 VTAIL.n281 10.4732
R502 VTAIL.n311 VTAIL.n310 10.4732
R503 VTAIL.n673 VTAIL.n652 9.69747
R504 VTAIL.n693 VTAIL.n642 9.69747
R505 VTAIL.n43 VTAIL.n22 9.69747
R506 VTAIL.n63 VTAIL.n12 9.69747
R507 VTAIL.n133 VTAIL.n112 9.69747
R508 VTAIL.n153 VTAIL.n102 9.69747
R509 VTAIL.n223 VTAIL.n202 9.69747
R510 VTAIL.n243 VTAIL.n192 9.69747
R511 VTAIL.n604 VTAIL.n553 9.69747
R512 VTAIL.n584 VTAIL.n563 9.69747
R513 VTAIL.n514 VTAIL.n463 9.69747
R514 VTAIL.n494 VTAIL.n473 9.69747
R515 VTAIL.n424 VTAIL.n373 9.69747
R516 VTAIL.n404 VTAIL.n383 9.69747
R517 VTAIL.n334 VTAIL.n283 9.69747
R518 VTAIL.n314 VTAIL.n293 9.69747
R519 VTAIL.n718 VTAIL.n717 9.45567
R520 VTAIL.n88 VTAIL.n87 9.45567
R521 VTAIL.n178 VTAIL.n177 9.45567
R522 VTAIL.n268 VTAIL.n267 9.45567
R523 VTAIL.n628 VTAIL.n627 9.45567
R524 VTAIL.n538 VTAIL.n537 9.45567
R525 VTAIL.n448 VTAIL.n447 9.45567
R526 VTAIL.n358 VTAIL.n357 9.45567
R527 VTAIL.n717 VTAIL.n716 9.3005
R528 VTAIL.n632 VTAIL.n631 9.3005
R529 VTAIL.n711 VTAIL.n710 9.3005
R530 VTAIL.n709 VTAIL.n708 9.3005
R531 VTAIL.n648 VTAIL.n647 9.3005
R532 VTAIL.n677 VTAIL.n676 9.3005
R533 VTAIL.n675 VTAIL.n674 9.3005
R534 VTAIL.n652 VTAIL.n651 9.3005
R535 VTAIL.n669 VTAIL.n668 9.3005
R536 VTAIL.n667 VTAIL.n666 9.3005
R537 VTAIL.n656 VTAIL.n655 9.3005
R538 VTAIL.n661 VTAIL.n660 9.3005
R539 VTAIL.n683 VTAIL.n682 9.3005
R540 VTAIL.n685 VTAIL.n684 9.3005
R541 VTAIL.n644 VTAIL.n643 9.3005
R542 VTAIL.n691 VTAIL.n690 9.3005
R543 VTAIL.n693 VTAIL.n692 9.3005
R544 VTAIL.n640 VTAIL.n639 9.3005
R545 VTAIL.n699 VTAIL.n698 9.3005
R546 VTAIL.n701 VTAIL.n700 9.3005
R547 VTAIL.n702 VTAIL.n635 9.3005
R548 VTAIL.n87 VTAIL.n86 9.3005
R549 VTAIL.n2 VTAIL.n1 9.3005
R550 VTAIL.n81 VTAIL.n80 9.3005
R551 VTAIL.n79 VTAIL.n78 9.3005
R552 VTAIL.n18 VTAIL.n17 9.3005
R553 VTAIL.n47 VTAIL.n46 9.3005
R554 VTAIL.n45 VTAIL.n44 9.3005
R555 VTAIL.n22 VTAIL.n21 9.3005
R556 VTAIL.n39 VTAIL.n38 9.3005
R557 VTAIL.n37 VTAIL.n36 9.3005
R558 VTAIL.n26 VTAIL.n25 9.3005
R559 VTAIL.n31 VTAIL.n30 9.3005
R560 VTAIL.n53 VTAIL.n52 9.3005
R561 VTAIL.n55 VTAIL.n54 9.3005
R562 VTAIL.n14 VTAIL.n13 9.3005
R563 VTAIL.n61 VTAIL.n60 9.3005
R564 VTAIL.n63 VTAIL.n62 9.3005
R565 VTAIL.n10 VTAIL.n9 9.3005
R566 VTAIL.n69 VTAIL.n68 9.3005
R567 VTAIL.n71 VTAIL.n70 9.3005
R568 VTAIL.n72 VTAIL.n5 9.3005
R569 VTAIL.n177 VTAIL.n176 9.3005
R570 VTAIL.n92 VTAIL.n91 9.3005
R571 VTAIL.n171 VTAIL.n170 9.3005
R572 VTAIL.n169 VTAIL.n168 9.3005
R573 VTAIL.n108 VTAIL.n107 9.3005
R574 VTAIL.n137 VTAIL.n136 9.3005
R575 VTAIL.n135 VTAIL.n134 9.3005
R576 VTAIL.n112 VTAIL.n111 9.3005
R577 VTAIL.n129 VTAIL.n128 9.3005
R578 VTAIL.n127 VTAIL.n126 9.3005
R579 VTAIL.n116 VTAIL.n115 9.3005
R580 VTAIL.n121 VTAIL.n120 9.3005
R581 VTAIL.n143 VTAIL.n142 9.3005
R582 VTAIL.n145 VTAIL.n144 9.3005
R583 VTAIL.n104 VTAIL.n103 9.3005
R584 VTAIL.n151 VTAIL.n150 9.3005
R585 VTAIL.n153 VTAIL.n152 9.3005
R586 VTAIL.n100 VTAIL.n99 9.3005
R587 VTAIL.n159 VTAIL.n158 9.3005
R588 VTAIL.n161 VTAIL.n160 9.3005
R589 VTAIL.n162 VTAIL.n95 9.3005
R590 VTAIL.n267 VTAIL.n266 9.3005
R591 VTAIL.n182 VTAIL.n181 9.3005
R592 VTAIL.n261 VTAIL.n260 9.3005
R593 VTAIL.n259 VTAIL.n258 9.3005
R594 VTAIL.n198 VTAIL.n197 9.3005
R595 VTAIL.n227 VTAIL.n226 9.3005
R596 VTAIL.n225 VTAIL.n224 9.3005
R597 VTAIL.n202 VTAIL.n201 9.3005
R598 VTAIL.n219 VTAIL.n218 9.3005
R599 VTAIL.n217 VTAIL.n216 9.3005
R600 VTAIL.n206 VTAIL.n205 9.3005
R601 VTAIL.n211 VTAIL.n210 9.3005
R602 VTAIL.n233 VTAIL.n232 9.3005
R603 VTAIL.n235 VTAIL.n234 9.3005
R604 VTAIL.n194 VTAIL.n193 9.3005
R605 VTAIL.n241 VTAIL.n240 9.3005
R606 VTAIL.n243 VTAIL.n242 9.3005
R607 VTAIL.n190 VTAIL.n189 9.3005
R608 VTAIL.n249 VTAIL.n248 9.3005
R609 VTAIL.n251 VTAIL.n250 9.3005
R610 VTAIL.n252 VTAIL.n185 9.3005
R611 VTAIL.n596 VTAIL.n595 9.3005
R612 VTAIL.n555 VTAIL.n554 9.3005
R613 VTAIL.n602 VTAIL.n601 9.3005
R614 VTAIL.n604 VTAIL.n603 9.3005
R615 VTAIL.n551 VTAIL.n550 9.3005
R616 VTAIL.n610 VTAIL.n609 9.3005
R617 VTAIL.n612 VTAIL.n611 9.3005
R618 VTAIL.n548 VTAIL.n545 9.3005
R619 VTAIL.n627 VTAIL.n626 9.3005
R620 VTAIL.n542 VTAIL.n541 9.3005
R621 VTAIL.n621 VTAIL.n620 9.3005
R622 VTAIL.n619 VTAIL.n618 9.3005
R623 VTAIL.n594 VTAIL.n593 9.3005
R624 VTAIL.n559 VTAIL.n558 9.3005
R625 VTAIL.n588 VTAIL.n587 9.3005
R626 VTAIL.n586 VTAIL.n585 9.3005
R627 VTAIL.n563 VTAIL.n562 9.3005
R628 VTAIL.n580 VTAIL.n579 9.3005
R629 VTAIL.n578 VTAIL.n577 9.3005
R630 VTAIL.n567 VTAIL.n566 9.3005
R631 VTAIL.n572 VTAIL.n571 9.3005
R632 VTAIL.n506 VTAIL.n505 9.3005
R633 VTAIL.n465 VTAIL.n464 9.3005
R634 VTAIL.n512 VTAIL.n511 9.3005
R635 VTAIL.n514 VTAIL.n513 9.3005
R636 VTAIL.n461 VTAIL.n460 9.3005
R637 VTAIL.n520 VTAIL.n519 9.3005
R638 VTAIL.n522 VTAIL.n521 9.3005
R639 VTAIL.n458 VTAIL.n455 9.3005
R640 VTAIL.n537 VTAIL.n536 9.3005
R641 VTAIL.n452 VTAIL.n451 9.3005
R642 VTAIL.n531 VTAIL.n530 9.3005
R643 VTAIL.n529 VTAIL.n528 9.3005
R644 VTAIL.n504 VTAIL.n503 9.3005
R645 VTAIL.n469 VTAIL.n468 9.3005
R646 VTAIL.n498 VTAIL.n497 9.3005
R647 VTAIL.n496 VTAIL.n495 9.3005
R648 VTAIL.n473 VTAIL.n472 9.3005
R649 VTAIL.n490 VTAIL.n489 9.3005
R650 VTAIL.n488 VTAIL.n487 9.3005
R651 VTAIL.n477 VTAIL.n476 9.3005
R652 VTAIL.n482 VTAIL.n481 9.3005
R653 VTAIL.n416 VTAIL.n415 9.3005
R654 VTAIL.n375 VTAIL.n374 9.3005
R655 VTAIL.n422 VTAIL.n421 9.3005
R656 VTAIL.n424 VTAIL.n423 9.3005
R657 VTAIL.n371 VTAIL.n370 9.3005
R658 VTAIL.n430 VTAIL.n429 9.3005
R659 VTAIL.n432 VTAIL.n431 9.3005
R660 VTAIL.n368 VTAIL.n365 9.3005
R661 VTAIL.n447 VTAIL.n446 9.3005
R662 VTAIL.n362 VTAIL.n361 9.3005
R663 VTAIL.n441 VTAIL.n440 9.3005
R664 VTAIL.n439 VTAIL.n438 9.3005
R665 VTAIL.n414 VTAIL.n413 9.3005
R666 VTAIL.n379 VTAIL.n378 9.3005
R667 VTAIL.n408 VTAIL.n407 9.3005
R668 VTAIL.n406 VTAIL.n405 9.3005
R669 VTAIL.n383 VTAIL.n382 9.3005
R670 VTAIL.n400 VTAIL.n399 9.3005
R671 VTAIL.n398 VTAIL.n397 9.3005
R672 VTAIL.n387 VTAIL.n386 9.3005
R673 VTAIL.n392 VTAIL.n391 9.3005
R674 VTAIL.n326 VTAIL.n325 9.3005
R675 VTAIL.n285 VTAIL.n284 9.3005
R676 VTAIL.n332 VTAIL.n331 9.3005
R677 VTAIL.n334 VTAIL.n333 9.3005
R678 VTAIL.n281 VTAIL.n280 9.3005
R679 VTAIL.n340 VTAIL.n339 9.3005
R680 VTAIL.n342 VTAIL.n341 9.3005
R681 VTAIL.n278 VTAIL.n275 9.3005
R682 VTAIL.n357 VTAIL.n356 9.3005
R683 VTAIL.n272 VTAIL.n271 9.3005
R684 VTAIL.n351 VTAIL.n350 9.3005
R685 VTAIL.n349 VTAIL.n348 9.3005
R686 VTAIL.n324 VTAIL.n323 9.3005
R687 VTAIL.n289 VTAIL.n288 9.3005
R688 VTAIL.n318 VTAIL.n317 9.3005
R689 VTAIL.n316 VTAIL.n315 9.3005
R690 VTAIL.n293 VTAIL.n292 9.3005
R691 VTAIL.n310 VTAIL.n309 9.3005
R692 VTAIL.n308 VTAIL.n307 9.3005
R693 VTAIL.n297 VTAIL.n296 9.3005
R694 VTAIL.n302 VTAIL.n301 9.3005
R695 VTAIL.n674 VTAIL.n650 8.92171
R696 VTAIL.n690 VTAIL.n689 8.92171
R697 VTAIL.n44 VTAIL.n20 8.92171
R698 VTAIL.n60 VTAIL.n59 8.92171
R699 VTAIL.n134 VTAIL.n110 8.92171
R700 VTAIL.n150 VTAIL.n149 8.92171
R701 VTAIL.n224 VTAIL.n200 8.92171
R702 VTAIL.n240 VTAIL.n239 8.92171
R703 VTAIL.n601 VTAIL.n600 8.92171
R704 VTAIL.n585 VTAIL.n561 8.92171
R705 VTAIL.n511 VTAIL.n510 8.92171
R706 VTAIL.n495 VTAIL.n471 8.92171
R707 VTAIL.n421 VTAIL.n420 8.92171
R708 VTAIL.n405 VTAIL.n381 8.92171
R709 VTAIL.n331 VTAIL.n330 8.92171
R710 VTAIL.n315 VTAIL.n291 8.92171
R711 VTAIL.n678 VTAIL.n677 8.14595
R712 VTAIL.n686 VTAIL.n644 8.14595
R713 VTAIL.n48 VTAIL.n47 8.14595
R714 VTAIL.n56 VTAIL.n14 8.14595
R715 VTAIL.n138 VTAIL.n137 8.14595
R716 VTAIL.n146 VTAIL.n104 8.14595
R717 VTAIL.n228 VTAIL.n227 8.14595
R718 VTAIL.n236 VTAIL.n194 8.14595
R719 VTAIL.n597 VTAIL.n555 8.14595
R720 VTAIL.n589 VTAIL.n588 8.14595
R721 VTAIL.n507 VTAIL.n465 8.14595
R722 VTAIL.n499 VTAIL.n498 8.14595
R723 VTAIL.n417 VTAIL.n375 8.14595
R724 VTAIL.n409 VTAIL.n408 8.14595
R725 VTAIL.n327 VTAIL.n285 8.14595
R726 VTAIL.n319 VTAIL.n318 8.14595
R727 VTAIL.n681 VTAIL.n648 7.3702
R728 VTAIL.n685 VTAIL.n646 7.3702
R729 VTAIL.n51 VTAIL.n18 7.3702
R730 VTAIL.n55 VTAIL.n16 7.3702
R731 VTAIL.n141 VTAIL.n108 7.3702
R732 VTAIL.n145 VTAIL.n106 7.3702
R733 VTAIL.n231 VTAIL.n198 7.3702
R734 VTAIL.n235 VTAIL.n196 7.3702
R735 VTAIL.n596 VTAIL.n557 7.3702
R736 VTAIL.n592 VTAIL.n559 7.3702
R737 VTAIL.n506 VTAIL.n467 7.3702
R738 VTAIL.n502 VTAIL.n469 7.3702
R739 VTAIL.n416 VTAIL.n377 7.3702
R740 VTAIL.n412 VTAIL.n379 7.3702
R741 VTAIL.n326 VTAIL.n287 7.3702
R742 VTAIL.n322 VTAIL.n289 7.3702
R743 VTAIL.n682 VTAIL.n681 6.59444
R744 VTAIL.n682 VTAIL.n646 6.59444
R745 VTAIL.n52 VTAIL.n51 6.59444
R746 VTAIL.n52 VTAIL.n16 6.59444
R747 VTAIL.n142 VTAIL.n141 6.59444
R748 VTAIL.n142 VTAIL.n106 6.59444
R749 VTAIL.n232 VTAIL.n231 6.59444
R750 VTAIL.n232 VTAIL.n196 6.59444
R751 VTAIL.n593 VTAIL.n557 6.59444
R752 VTAIL.n593 VTAIL.n592 6.59444
R753 VTAIL.n503 VTAIL.n467 6.59444
R754 VTAIL.n503 VTAIL.n502 6.59444
R755 VTAIL.n413 VTAIL.n377 6.59444
R756 VTAIL.n413 VTAIL.n412 6.59444
R757 VTAIL.n323 VTAIL.n287 6.59444
R758 VTAIL.n323 VTAIL.n322 6.59444
R759 VTAIL.n678 VTAIL.n648 5.81868
R760 VTAIL.n686 VTAIL.n685 5.81868
R761 VTAIL.n48 VTAIL.n18 5.81868
R762 VTAIL.n56 VTAIL.n55 5.81868
R763 VTAIL.n138 VTAIL.n108 5.81868
R764 VTAIL.n146 VTAIL.n145 5.81868
R765 VTAIL.n228 VTAIL.n198 5.81868
R766 VTAIL.n236 VTAIL.n235 5.81868
R767 VTAIL.n597 VTAIL.n596 5.81868
R768 VTAIL.n589 VTAIL.n559 5.81868
R769 VTAIL.n507 VTAIL.n506 5.81868
R770 VTAIL.n499 VTAIL.n469 5.81868
R771 VTAIL.n417 VTAIL.n416 5.81868
R772 VTAIL.n409 VTAIL.n379 5.81868
R773 VTAIL.n327 VTAIL.n326 5.81868
R774 VTAIL.n319 VTAIL.n289 5.81868
R775 VTAIL.n677 VTAIL.n650 5.04292
R776 VTAIL.n689 VTAIL.n644 5.04292
R777 VTAIL.n47 VTAIL.n20 5.04292
R778 VTAIL.n59 VTAIL.n14 5.04292
R779 VTAIL.n137 VTAIL.n110 5.04292
R780 VTAIL.n149 VTAIL.n104 5.04292
R781 VTAIL.n227 VTAIL.n200 5.04292
R782 VTAIL.n239 VTAIL.n194 5.04292
R783 VTAIL.n600 VTAIL.n555 5.04292
R784 VTAIL.n588 VTAIL.n561 5.04292
R785 VTAIL.n510 VTAIL.n465 5.04292
R786 VTAIL.n498 VTAIL.n471 5.04292
R787 VTAIL.n420 VTAIL.n375 5.04292
R788 VTAIL.n408 VTAIL.n381 5.04292
R789 VTAIL.n330 VTAIL.n285 5.04292
R790 VTAIL.n318 VTAIL.n291 5.04292
R791 VTAIL.n674 VTAIL.n673 4.26717
R792 VTAIL.n690 VTAIL.n642 4.26717
R793 VTAIL.n44 VTAIL.n43 4.26717
R794 VTAIL.n60 VTAIL.n12 4.26717
R795 VTAIL.n134 VTAIL.n133 4.26717
R796 VTAIL.n150 VTAIL.n102 4.26717
R797 VTAIL.n224 VTAIL.n223 4.26717
R798 VTAIL.n240 VTAIL.n192 4.26717
R799 VTAIL.n601 VTAIL.n553 4.26717
R800 VTAIL.n585 VTAIL.n584 4.26717
R801 VTAIL.n511 VTAIL.n463 4.26717
R802 VTAIL.n495 VTAIL.n494 4.26717
R803 VTAIL.n421 VTAIL.n373 4.26717
R804 VTAIL.n405 VTAIL.n404 4.26717
R805 VTAIL.n331 VTAIL.n283 4.26717
R806 VTAIL.n315 VTAIL.n314 4.26717
R807 VTAIL.n660 VTAIL.n659 3.70982
R808 VTAIL.n30 VTAIL.n29 3.70982
R809 VTAIL.n120 VTAIL.n119 3.70982
R810 VTAIL.n210 VTAIL.n209 3.70982
R811 VTAIL.n571 VTAIL.n570 3.70982
R812 VTAIL.n481 VTAIL.n480 3.70982
R813 VTAIL.n391 VTAIL.n390 3.70982
R814 VTAIL.n301 VTAIL.n300 3.70982
R815 VTAIL.n670 VTAIL.n652 3.49141
R816 VTAIL.n694 VTAIL.n693 3.49141
R817 VTAIL.n718 VTAIL.n630 3.49141
R818 VTAIL.n40 VTAIL.n22 3.49141
R819 VTAIL.n64 VTAIL.n63 3.49141
R820 VTAIL.n88 VTAIL.n0 3.49141
R821 VTAIL.n130 VTAIL.n112 3.49141
R822 VTAIL.n154 VTAIL.n153 3.49141
R823 VTAIL.n178 VTAIL.n90 3.49141
R824 VTAIL.n220 VTAIL.n202 3.49141
R825 VTAIL.n244 VTAIL.n243 3.49141
R826 VTAIL.n268 VTAIL.n180 3.49141
R827 VTAIL.n628 VTAIL.n540 3.49141
R828 VTAIL.n605 VTAIL.n604 3.49141
R829 VTAIL.n581 VTAIL.n563 3.49141
R830 VTAIL.n538 VTAIL.n450 3.49141
R831 VTAIL.n515 VTAIL.n514 3.49141
R832 VTAIL.n491 VTAIL.n473 3.49141
R833 VTAIL.n448 VTAIL.n360 3.49141
R834 VTAIL.n425 VTAIL.n424 3.49141
R835 VTAIL.n401 VTAIL.n383 3.49141
R836 VTAIL.n358 VTAIL.n270 3.49141
R837 VTAIL.n335 VTAIL.n334 3.49141
R838 VTAIL.n311 VTAIL.n293 3.49141
R839 VTAIL.n669 VTAIL.n654 2.71565
R840 VTAIL.n697 VTAIL.n640 2.71565
R841 VTAIL.n716 VTAIL.n715 2.71565
R842 VTAIL.n39 VTAIL.n24 2.71565
R843 VTAIL.n67 VTAIL.n10 2.71565
R844 VTAIL.n86 VTAIL.n85 2.71565
R845 VTAIL.n129 VTAIL.n114 2.71565
R846 VTAIL.n157 VTAIL.n100 2.71565
R847 VTAIL.n176 VTAIL.n175 2.71565
R848 VTAIL.n219 VTAIL.n204 2.71565
R849 VTAIL.n247 VTAIL.n190 2.71565
R850 VTAIL.n266 VTAIL.n265 2.71565
R851 VTAIL.n626 VTAIL.n625 2.71565
R852 VTAIL.n608 VTAIL.n551 2.71565
R853 VTAIL.n580 VTAIL.n565 2.71565
R854 VTAIL.n536 VTAIL.n535 2.71565
R855 VTAIL.n518 VTAIL.n461 2.71565
R856 VTAIL.n490 VTAIL.n475 2.71565
R857 VTAIL.n446 VTAIL.n445 2.71565
R858 VTAIL.n428 VTAIL.n371 2.71565
R859 VTAIL.n400 VTAIL.n385 2.71565
R860 VTAIL.n356 VTAIL.n355 2.71565
R861 VTAIL.n338 VTAIL.n281 2.71565
R862 VTAIL.n310 VTAIL.n295 2.71565
R863 VTAIL.n666 VTAIL.n665 1.93989
R864 VTAIL.n698 VTAIL.n638 1.93989
R865 VTAIL.n712 VTAIL.n632 1.93989
R866 VTAIL.n36 VTAIL.n35 1.93989
R867 VTAIL.n68 VTAIL.n8 1.93989
R868 VTAIL.n82 VTAIL.n2 1.93989
R869 VTAIL.n126 VTAIL.n125 1.93989
R870 VTAIL.n158 VTAIL.n98 1.93989
R871 VTAIL.n172 VTAIL.n92 1.93989
R872 VTAIL.n216 VTAIL.n215 1.93989
R873 VTAIL.n248 VTAIL.n188 1.93989
R874 VTAIL.n262 VTAIL.n182 1.93989
R875 VTAIL.n622 VTAIL.n542 1.93989
R876 VTAIL.n609 VTAIL.n549 1.93989
R877 VTAIL.n577 VTAIL.n576 1.93989
R878 VTAIL.n532 VTAIL.n452 1.93989
R879 VTAIL.n519 VTAIL.n459 1.93989
R880 VTAIL.n487 VTAIL.n486 1.93989
R881 VTAIL.n442 VTAIL.n362 1.93989
R882 VTAIL.n429 VTAIL.n369 1.93989
R883 VTAIL.n397 VTAIL.n396 1.93989
R884 VTAIL.n352 VTAIL.n272 1.93989
R885 VTAIL.n339 VTAIL.n279 1.93989
R886 VTAIL.n307 VTAIL.n306 1.93989
R887 VTAIL.n662 VTAIL.n656 1.16414
R888 VTAIL.n703 VTAIL.n701 1.16414
R889 VTAIL.n711 VTAIL.n634 1.16414
R890 VTAIL.n32 VTAIL.n26 1.16414
R891 VTAIL.n73 VTAIL.n71 1.16414
R892 VTAIL.n81 VTAIL.n4 1.16414
R893 VTAIL.n122 VTAIL.n116 1.16414
R894 VTAIL.n163 VTAIL.n161 1.16414
R895 VTAIL.n171 VTAIL.n94 1.16414
R896 VTAIL.n212 VTAIL.n206 1.16414
R897 VTAIL.n253 VTAIL.n251 1.16414
R898 VTAIL.n261 VTAIL.n184 1.16414
R899 VTAIL.n621 VTAIL.n544 1.16414
R900 VTAIL.n613 VTAIL.n612 1.16414
R901 VTAIL.n573 VTAIL.n567 1.16414
R902 VTAIL.n531 VTAIL.n454 1.16414
R903 VTAIL.n523 VTAIL.n522 1.16414
R904 VTAIL.n483 VTAIL.n477 1.16414
R905 VTAIL.n441 VTAIL.n364 1.16414
R906 VTAIL.n433 VTAIL.n432 1.16414
R907 VTAIL.n393 VTAIL.n387 1.16414
R908 VTAIL.n351 VTAIL.n274 1.16414
R909 VTAIL.n343 VTAIL.n342 1.16414
R910 VTAIL.n303 VTAIL.n297 1.16414
R911 VTAIL.n449 VTAIL.n359 0.966017
R912 VTAIL.n629 VTAIL.n539 0.966017
R913 VTAIL.n269 VTAIL.n179 0.966017
R914 VTAIL VTAIL.n89 0.541448
R915 VTAIL.n539 VTAIL.n449 0.470328
R916 VTAIL.n179 VTAIL.n89 0.470328
R917 VTAIL VTAIL.n719 0.425069
R918 VTAIL.n661 VTAIL.n658 0.388379
R919 VTAIL.n702 VTAIL.n636 0.388379
R920 VTAIL.n708 VTAIL.n707 0.388379
R921 VTAIL.n31 VTAIL.n28 0.388379
R922 VTAIL.n72 VTAIL.n6 0.388379
R923 VTAIL.n78 VTAIL.n77 0.388379
R924 VTAIL.n121 VTAIL.n118 0.388379
R925 VTAIL.n162 VTAIL.n96 0.388379
R926 VTAIL.n168 VTAIL.n167 0.388379
R927 VTAIL.n211 VTAIL.n208 0.388379
R928 VTAIL.n252 VTAIL.n186 0.388379
R929 VTAIL.n258 VTAIL.n257 0.388379
R930 VTAIL.n618 VTAIL.n617 0.388379
R931 VTAIL.n548 VTAIL.n546 0.388379
R932 VTAIL.n572 VTAIL.n569 0.388379
R933 VTAIL.n528 VTAIL.n527 0.388379
R934 VTAIL.n458 VTAIL.n456 0.388379
R935 VTAIL.n482 VTAIL.n479 0.388379
R936 VTAIL.n438 VTAIL.n437 0.388379
R937 VTAIL.n368 VTAIL.n366 0.388379
R938 VTAIL.n392 VTAIL.n389 0.388379
R939 VTAIL.n348 VTAIL.n347 0.388379
R940 VTAIL.n278 VTAIL.n276 0.388379
R941 VTAIL.n302 VTAIL.n299 0.388379
R942 VTAIL.n660 VTAIL.n655 0.155672
R943 VTAIL.n667 VTAIL.n655 0.155672
R944 VTAIL.n668 VTAIL.n667 0.155672
R945 VTAIL.n668 VTAIL.n651 0.155672
R946 VTAIL.n675 VTAIL.n651 0.155672
R947 VTAIL.n676 VTAIL.n675 0.155672
R948 VTAIL.n676 VTAIL.n647 0.155672
R949 VTAIL.n683 VTAIL.n647 0.155672
R950 VTAIL.n684 VTAIL.n683 0.155672
R951 VTAIL.n684 VTAIL.n643 0.155672
R952 VTAIL.n691 VTAIL.n643 0.155672
R953 VTAIL.n692 VTAIL.n691 0.155672
R954 VTAIL.n692 VTAIL.n639 0.155672
R955 VTAIL.n699 VTAIL.n639 0.155672
R956 VTAIL.n700 VTAIL.n699 0.155672
R957 VTAIL.n700 VTAIL.n635 0.155672
R958 VTAIL.n709 VTAIL.n635 0.155672
R959 VTAIL.n710 VTAIL.n709 0.155672
R960 VTAIL.n710 VTAIL.n631 0.155672
R961 VTAIL.n717 VTAIL.n631 0.155672
R962 VTAIL.n30 VTAIL.n25 0.155672
R963 VTAIL.n37 VTAIL.n25 0.155672
R964 VTAIL.n38 VTAIL.n37 0.155672
R965 VTAIL.n38 VTAIL.n21 0.155672
R966 VTAIL.n45 VTAIL.n21 0.155672
R967 VTAIL.n46 VTAIL.n45 0.155672
R968 VTAIL.n46 VTAIL.n17 0.155672
R969 VTAIL.n53 VTAIL.n17 0.155672
R970 VTAIL.n54 VTAIL.n53 0.155672
R971 VTAIL.n54 VTAIL.n13 0.155672
R972 VTAIL.n61 VTAIL.n13 0.155672
R973 VTAIL.n62 VTAIL.n61 0.155672
R974 VTAIL.n62 VTAIL.n9 0.155672
R975 VTAIL.n69 VTAIL.n9 0.155672
R976 VTAIL.n70 VTAIL.n69 0.155672
R977 VTAIL.n70 VTAIL.n5 0.155672
R978 VTAIL.n79 VTAIL.n5 0.155672
R979 VTAIL.n80 VTAIL.n79 0.155672
R980 VTAIL.n80 VTAIL.n1 0.155672
R981 VTAIL.n87 VTAIL.n1 0.155672
R982 VTAIL.n120 VTAIL.n115 0.155672
R983 VTAIL.n127 VTAIL.n115 0.155672
R984 VTAIL.n128 VTAIL.n127 0.155672
R985 VTAIL.n128 VTAIL.n111 0.155672
R986 VTAIL.n135 VTAIL.n111 0.155672
R987 VTAIL.n136 VTAIL.n135 0.155672
R988 VTAIL.n136 VTAIL.n107 0.155672
R989 VTAIL.n143 VTAIL.n107 0.155672
R990 VTAIL.n144 VTAIL.n143 0.155672
R991 VTAIL.n144 VTAIL.n103 0.155672
R992 VTAIL.n151 VTAIL.n103 0.155672
R993 VTAIL.n152 VTAIL.n151 0.155672
R994 VTAIL.n152 VTAIL.n99 0.155672
R995 VTAIL.n159 VTAIL.n99 0.155672
R996 VTAIL.n160 VTAIL.n159 0.155672
R997 VTAIL.n160 VTAIL.n95 0.155672
R998 VTAIL.n169 VTAIL.n95 0.155672
R999 VTAIL.n170 VTAIL.n169 0.155672
R1000 VTAIL.n170 VTAIL.n91 0.155672
R1001 VTAIL.n177 VTAIL.n91 0.155672
R1002 VTAIL.n210 VTAIL.n205 0.155672
R1003 VTAIL.n217 VTAIL.n205 0.155672
R1004 VTAIL.n218 VTAIL.n217 0.155672
R1005 VTAIL.n218 VTAIL.n201 0.155672
R1006 VTAIL.n225 VTAIL.n201 0.155672
R1007 VTAIL.n226 VTAIL.n225 0.155672
R1008 VTAIL.n226 VTAIL.n197 0.155672
R1009 VTAIL.n233 VTAIL.n197 0.155672
R1010 VTAIL.n234 VTAIL.n233 0.155672
R1011 VTAIL.n234 VTAIL.n193 0.155672
R1012 VTAIL.n241 VTAIL.n193 0.155672
R1013 VTAIL.n242 VTAIL.n241 0.155672
R1014 VTAIL.n242 VTAIL.n189 0.155672
R1015 VTAIL.n249 VTAIL.n189 0.155672
R1016 VTAIL.n250 VTAIL.n249 0.155672
R1017 VTAIL.n250 VTAIL.n185 0.155672
R1018 VTAIL.n259 VTAIL.n185 0.155672
R1019 VTAIL.n260 VTAIL.n259 0.155672
R1020 VTAIL.n260 VTAIL.n181 0.155672
R1021 VTAIL.n267 VTAIL.n181 0.155672
R1022 VTAIL.n627 VTAIL.n541 0.155672
R1023 VTAIL.n620 VTAIL.n541 0.155672
R1024 VTAIL.n620 VTAIL.n619 0.155672
R1025 VTAIL.n619 VTAIL.n545 0.155672
R1026 VTAIL.n611 VTAIL.n545 0.155672
R1027 VTAIL.n611 VTAIL.n610 0.155672
R1028 VTAIL.n610 VTAIL.n550 0.155672
R1029 VTAIL.n603 VTAIL.n550 0.155672
R1030 VTAIL.n603 VTAIL.n602 0.155672
R1031 VTAIL.n602 VTAIL.n554 0.155672
R1032 VTAIL.n595 VTAIL.n554 0.155672
R1033 VTAIL.n595 VTAIL.n594 0.155672
R1034 VTAIL.n594 VTAIL.n558 0.155672
R1035 VTAIL.n587 VTAIL.n558 0.155672
R1036 VTAIL.n587 VTAIL.n586 0.155672
R1037 VTAIL.n586 VTAIL.n562 0.155672
R1038 VTAIL.n579 VTAIL.n562 0.155672
R1039 VTAIL.n579 VTAIL.n578 0.155672
R1040 VTAIL.n578 VTAIL.n566 0.155672
R1041 VTAIL.n571 VTAIL.n566 0.155672
R1042 VTAIL.n537 VTAIL.n451 0.155672
R1043 VTAIL.n530 VTAIL.n451 0.155672
R1044 VTAIL.n530 VTAIL.n529 0.155672
R1045 VTAIL.n529 VTAIL.n455 0.155672
R1046 VTAIL.n521 VTAIL.n455 0.155672
R1047 VTAIL.n521 VTAIL.n520 0.155672
R1048 VTAIL.n520 VTAIL.n460 0.155672
R1049 VTAIL.n513 VTAIL.n460 0.155672
R1050 VTAIL.n513 VTAIL.n512 0.155672
R1051 VTAIL.n512 VTAIL.n464 0.155672
R1052 VTAIL.n505 VTAIL.n464 0.155672
R1053 VTAIL.n505 VTAIL.n504 0.155672
R1054 VTAIL.n504 VTAIL.n468 0.155672
R1055 VTAIL.n497 VTAIL.n468 0.155672
R1056 VTAIL.n497 VTAIL.n496 0.155672
R1057 VTAIL.n496 VTAIL.n472 0.155672
R1058 VTAIL.n489 VTAIL.n472 0.155672
R1059 VTAIL.n489 VTAIL.n488 0.155672
R1060 VTAIL.n488 VTAIL.n476 0.155672
R1061 VTAIL.n481 VTAIL.n476 0.155672
R1062 VTAIL.n447 VTAIL.n361 0.155672
R1063 VTAIL.n440 VTAIL.n361 0.155672
R1064 VTAIL.n440 VTAIL.n439 0.155672
R1065 VTAIL.n439 VTAIL.n365 0.155672
R1066 VTAIL.n431 VTAIL.n365 0.155672
R1067 VTAIL.n431 VTAIL.n430 0.155672
R1068 VTAIL.n430 VTAIL.n370 0.155672
R1069 VTAIL.n423 VTAIL.n370 0.155672
R1070 VTAIL.n423 VTAIL.n422 0.155672
R1071 VTAIL.n422 VTAIL.n374 0.155672
R1072 VTAIL.n415 VTAIL.n374 0.155672
R1073 VTAIL.n415 VTAIL.n414 0.155672
R1074 VTAIL.n414 VTAIL.n378 0.155672
R1075 VTAIL.n407 VTAIL.n378 0.155672
R1076 VTAIL.n407 VTAIL.n406 0.155672
R1077 VTAIL.n406 VTAIL.n382 0.155672
R1078 VTAIL.n399 VTAIL.n382 0.155672
R1079 VTAIL.n399 VTAIL.n398 0.155672
R1080 VTAIL.n398 VTAIL.n386 0.155672
R1081 VTAIL.n391 VTAIL.n386 0.155672
R1082 VTAIL.n357 VTAIL.n271 0.155672
R1083 VTAIL.n350 VTAIL.n271 0.155672
R1084 VTAIL.n350 VTAIL.n349 0.155672
R1085 VTAIL.n349 VTAIL.n275 0.155672
R1086 VTAIL.n341 VTAIL.n275 0.155672
R1087 VTAIL.n341 VTAIL.n340 0.155672
R1088 VTAIL.n340 VTAIL.n280 0.155672
R1089 VTAIL.n333 VTAIL.n280 0.155672
R1090 VTAIL.n333 VTAIL.n332 0.155672
R1091 VTAIL.n332 VTAIL.n284 0.155672
R1092 VTAIL.n325 VTAIL.n284 0.155672
R1093 VTAIL.n325 VTAIL.n324 0.155672
R1094 VTAIL.n324 VTAIL.n288 0.155672
R1095 VTAIL.n317 VTAIL.n288 0.155672
R1096 VTAIL.n317 VTAIL.n316 0.155672
R1097 VTAIL.n316 VTAIL.n292 0.155672
R1098 VTAIL.n309 VTAIL.n292 0.155672
R1099 VTAIL.n309 VTAIL.n308 0.155672
R1100 VTAIL.n308 VTAIL.n296 0.155672
R1101 VTAIL.n301 VTAIL.n296 0.155672
R1102 B.n119 B.t0 691.001
R1103 B.n127 B.t3 691.001
R1104 B.n38 B.t9 691.001
R1105 B.n46 B.t6 691.001
R1106 B.n421 B.n420 585
R1107 B.n422 B.n73 585
R1108 B.n424 B.n423 585
R1109 B.n425 B.n72 585
R1110 B.n427 B.n426 585
R1111 B.n428 B.n71 585
R1112 B.n430 B.n429 585
R1113 B.n431 B.n70 585
R1114 B.n433 B.n432 585
R1115 B.n434 B.n69 585
R1116 B.n436 B.n435 585
R1117 B.n437 B.n68 585
R1118 B.n439 B.n438 585
R1119 B.n440 B.n67 585
R1120 B.n442 B.n441 585
R1121 B.n443 B.n66 585
R1122 B.n445 B.n444 585
R1123 B.n446 B.n65 585
R1124 B.n448 B.n447 585
R1125 B.n449 B.n64 585
R1126 B.n451 B.n450 585
R1127 B.n452 B.n63 585
R1128 B.n454 B.n453 585
R1129 B.n455 B.n62 585
R1130 B.n457 B.n456 585
R1131 B.n458 B.n61 585
R1132 B.n460 B.n459 585
R1133 B.n461 B.n60 585
R1134 B.n463 B.n462 585
R1135 B.n464 B.n59 585
R1136 B.n466 B.n465 585
R1137 B.n467 B.n58 585
R1138 B.n469 B.n468 585
R1139 B.n470 B.n57 585
R1140 B.n472 B.n471 585
R1141 B.n473 B.n56 585
R1142 B.n475 B.n474 585
R1143 B.n476 B.n55 585
R1144 B.n478 B.n477 585
R1145 B.n479 B.n54 585
R1146 B.n481 B.n480 585
R1147 B.n482 B.n53 585
R1148 B.n484 B.n483 585
R1149 B.n485 B.n52 585
R1150 B.n487 B.n486 585
R1151 B.n488 B.n51 585
R1152 B.n490 B.n489 585
R1153 B.n491 B.n50 585
R1154 B.n493 B.n492 585
R1155 B.n494 B.n49 585
R1156 B.n496 B.n495 585
R1157 B.n497 B.n45 585
R1158 B.n499 B.n498 585
R1159 B.n500 B.n44 585
R1160 B.n502 B.n501 585
R1161 B.n503 B.n43 585
R1162 B.n505 B.n504 585
R1163 B.n506 B.n42 585
R1164 B.n508 B.n507 585
R1165 B.n509 B.n41 585
R1166 B.n511 B.n510 585
R1167 B.n512 B.n40 585
R1168 B.n514 B.n513 585
R1169 B.n516 B.n37 585
R1170 B.n518 B.n517 585
R1171 B.n519 B.n36 585
R1172 B.n521 B.n520 585
R1173 B.n522 B.n35 585
R1174 B.n524 B.n523 585
R1175 B.n525 B.n34 585
R1176 B.n527 B.n526 585
R1177 B.n528 B.n33 585
R1178 B.n530 B.n529 585
R1179 B.n531 B.n32 585
R1180 B.n533 B.n532 585
R1181 B.n534 B.n31 585
R1182 B.n536 B.n535 585
R1183 B.n537 B.n30 585
R1184 B.n539 B.n538 585
R1185 B.n540 B.n29 585
R1186 B.n542 B.n541 585
R1187 B.n543 B.n28 585
R1188 B.n545 B.n544 585
R1189 B.n546 B.n27 585
R1190 B.n548 B.n547 585
R1191 B.n549 B.n26 585
R1192 B.n551 B.n550 585
R1193 B.n552 B.n25 585
R1194 B.n554 B.n553 585
R1195 B.n555 B.n24 585
R1196 B.n557 B.n556 585
R1197 B.n558 B.n23 585
R1198 B.n560 B.n559 585
R1199 B.n561 B.n22 585
R1200 B.n563 B.n562 585
R1201 B.n564 B.n21 585
R1202 B.n566 B.n565 585
R1203 B.n567 B.n20 585
R1204 B.n569 B.n568 585
R1205 B.n570 B.n19 585
R1206 B.n572 B.n571 585
R1207 B.n573 B.n18 585
R1208 B.n575 B.n574 585
R1209 B.n576 B.n17 585
R1210 B.n578 B.n577 585
R1211 B.n579 B.n16 585
R1212 B.n581 B.n580 585
R1213 B.n582 B.n15 585
R1214 B.n584 B.n583 585
R1215 B.n585 B.n14 585
R1216 B.n587 B.n586 585
R1217 B.n588 B.n13 585
R1218 B.n590 B.n589 585
R1219 B.n591 B.n12 585
R1220 B.n593 B.n592 585
R1221 B.n594 B.n11 585
R1222 B.n419 B.n74 585
R1223 B.n418 B.n417 585
R1224 B.n416 B.n75 585
R1225 B.n415 B.n414 585
R1226 B.n413 B.n76 585
R1227 B.n412 B.n411 585
R1228 B.n410 B.n77 585
R1229 B.n409 B.n408 585
R1230 B.n407 B.n78 585
R1231 B.n406 B.n405 585
R1232 B.n404 B.n79 585
R1233 B.n403 B.n402 585
R1234 B.n401 B.n80 585
R1235 B.n400 B.n399 585
R1236 B.n398 B.n81 585
R1237 B.n397 B.n396 585
R1238 B.n395 B.n82 585
R1239 B.n394 B.n393 585
R1240 B.n392 B.n83 585
R1241 B.n391 B.n390 585
R1242 B.n389 B.n84 585
R1243 B.n388 B.n387 585
R1244 B.n386 B.n85 585
R1245 B.n385 B.n384 585
R1246 B.n383 B.n86 585
R1247 B.n382 B.n381 585
R1248 B.n380 B.n87 585
R1249 B.n379 B.n378 585
R1250 B.n377 B.n88 585
R1251 B.n376 B.n375 585
R1252 B.n374 B.n89 585
R1253 B.n373 B.n372 585
R1254 B.n371 B.n90 585
R1255 B.n370 B.n369 585
R1256 B.n368 B.n91 585
R1257 B.n367 B.n366 585
R1258 B.n365 B.n92 585
R1259 B.n190 B.n189 585
R1260 B.n191 B.n154 585
R1261 B.n193 B.n192 585
R1262 B.n194 B.n153 585
R1263 B.n196 B.n195 585
R1264 B.n197 B.n152 585
R1265 B.n199 B.n198 585
R1266 B.n200 B.n151 585
R1267 B.n202 B.n201 585
R1268 B.n203 B.n150 585
R1269 B.n205 B.n204 585
R1270 B.n206 B.n149 585
R1271 B.n208 B.n207 585
R1272 B.n209 B.n148 585
R1273 B.n211 B.n210 585
R1274 B.n212 B.n147 585
R1275 B.n214 B.n213 585
R1276 B.n215 B.n146 585
R1277 B.n217 B.n216 585
R1278 B.n218 B.n145 585
R1279 B.n220 B.n219 585
R1280 B.n221 B.n144 585
R1281 B.n223 B.n222 585
R1282 B.n224 B.n143 585
R1283 B.n226 B.n225 585
R1284 B.n227 B.n142 585
R1285 B.n229 B.n228 585
R1286 B.n230 B.n141 585
R1287 B.n232 B.n231 585
R1288 B.n233 B.n140 585
R1289 B.n235 B.n234 585
R1290 B.n236 B.n139 585
R1291 B.n238 B.n237 585
R1292 B.n239 B.n138 585
R1293 B.n241 B.n240 585
R1294 B.n242 B.n137 585
R1295 B.n244 B.n243 585
R1296 B.n245 B.n136 585
R1297 B.n247 B.n246 585
R1298 B.n248 B.n135 585
R1299 B.n250 B.n249 585
R1300 B.n251 B.n134 585
R1301 B.n253 B.n252 585
R1302 B.n254 B.n133 585
R1303 B.n256 B.n255 585
R1304 B.n257 B.n132 585
R1305 B.n259 B.n258 585
R1306 B.n260 B.n131 585
R1307 B.n262 B.n261 585
R1308 B.n263 B.n130 585
R1309 B.n265 B.n264 585
R1310 B.n266 B.n129 585
R1311 B.n268 B.n267 585
R1312 B.n270 B.n126 585
R1313 B.n272 B.n271 585
R1314 B.n273 B.n125 585
R1315 B.n275 B.n274 585
R1316 B.n276 B.n124 585
R1317 B.n278 B.n277 585
R1318 B.n279 B.n123 585
R1319 B.n281 B.n280 585
R1320 B.n282 B.n122 585
R1321 B.n284 B.n283 585
R1322 B.n286 B.n285 585
R1323 B.n287 B.n118 585
R1324 B.n289 B.n288 585
R1325 B.n290 B.n117 585
R1326 B.n292 B.n291 585
R1327 B.n293 B.n116 585
R1328 B.n295 B.n294 585
R1329 B.n296 B.n115 585
R1330 B.n298 B.n297 585
R1331 B.n299 B.n114 585
R1332 B.n301 B.n300 585
R1333 B.n302 B.n113 585
R1334 B.n304 B.n303 585
R1335 B.n305 B.n112 585
R1336 B.n307 B.n306 585
R1337 B.n308 B.n111 585
R1338 B.n310 B.n309 585
R1339 B.n311 B.n110 585
R1340 B.n313 B.n312 585
R1341 B.n314 B.n109 585
R1342 B.n316 B.n315 585
R1343 B.n317 B.n108 585
R1344 B.n319 B.n318 585
R1345 B.n320 B.n107 585
R1346 B.n322 B.n321 585
R1347 B.n323 B.n106 585
R1348 B.n325 B.n324 585
R1349 B.n326 B.n105 585
R1350 B.n328 B.n327 585
R1351 B.n329 B.n104 585
R1352 B.n331 B.n330 585
R1353 B.n332 B.n103 585
R1354 B.n334 B.n333 585
R1355 B.n335 B.n102 585
R1356 B.n337 B.n336 585
R1357 B.n338 B.n101 585
R1358 B.n340 B.n339 585
R1359 B.n341 B.n100 585
R1360 B.n343 B.n342 585
R1361 B.n344 B.n99 585
R1362 B.n346 B.n345 585
R1363 B.n347 B.n98 585
R1364 B.n349 B.n348 585
R1365 B.n350 B.n97 585
R1366 B.n352 B.n351 585
R1367 B.n353 B.n96 585
R1368 B.n355 B.n354 585
R1369 B.n356 B.n95 585
R1370 B.n358 B.n357 585
R1371 B.n359 B.n94 585
R1372 B.n361 B.n360 585
R1373 B.n362 B.n93 585
R1374 B.n364 B.n363 585
R1375 B.n188 B.n155 585
R1376 B.n187 B.n186 585
R1377 B.n185 B.n156 585
R1378 B.n184 B.n183 585
R1379 B.n182 B.n157 585
R1380 B.n181 B.n180 585
R1381 B.n179 B.n158 585
R1382 B.n178 B.n177 585
R1383 B.n176 B.n159 585
R1384 B.n175 B.n174 585
R1385 B.n173 B.n160 585
R1386 B.n172 B.n171 585
R1387 B.n170 B.n161 585
R1388 B.n169 B.n168 585
R1389 B.n167 B.n162 585
R1390 B.n166 B.n165 585
R1391 B.n164 B.n163 585
R1392 B.n2 B.n0 585
R1393 B.n621 B.n1 585
R1394 B.n620 B.n619 585
R1395 B.n618 B.n3 585
R1396 B.n617 B.n616 585
R1397 B.n615 B.n4 585
R1398 B.n614 B.n613 585
R1399 B.n612 B.n5 585
R1400 B.n611 B.n610 585
R1401 B.n609 B.n6 585
R1402 B.n608 B.n607 585
R1403 B.n606 B.n7 585
R1404 B.n605 B.n604 585
R1405 B.n603 B.n8 585
R1406 B.n602 B.n601 585
R1407 B.n600 B.n9 585
R1408 B.n599 B.n598 585
R1409 B.n597 B.n10 585
R1410 B.n596 B.n595 585
R1411 B.n623 B.n622 585
R1412 B.n189 B.n188 540.549
R1413 B.n596 B.n11 540.549
R1414 B.n363 B.n92 540.549
R1415 B.n421 B.n74 540.549
R1416 B.n119 B.t2 469.769
R1417 B.n46 B.t7 469.769
R1418 B.n127 B.t5 469.769
R1419 B.n38 B.t10 469.769
R1420 B.n120 B.t1 448.048
R1421 B.n47 B.t8 448.048
R1422 B.n128 B.t4 448.046
R1423 B.n39 B.t11 448.046
R1424 B.n188 B.n187 163.367
R1425 B.n187 B.n156 163.367
R1426 B.n183 B.n156 163.367
R1427 B.n183 B.n182 163.367
R1428 B.n182 B.n181 163.367
R1429 B.n181 B.n158 163.367
R1430 B.n177 B.n158 163.367
R1431 B.n177 B.n176 163.367
R1432 B.n176 B.n175 163.367
R1433 B.n175 B.n160 163.367
R1434 B.n171 B.n160 163.367
R1435 B.n171 B.n170 163.367
R1436 B.n170 B.n169 163.367
R1437 B.n169 B.n162 163.367
R1438 B.n165 B.n162 163.367
R1439 B.n165 B.n164 163.367
R1440 B.n164 B.n2 163.367
R1441 B.n622 B.n2 163.367
R1442 B.n622 B.n621 163.367
R1443 B.n621 B.n620 163.367
R1444 B.n620 B.n3 163.367
R1445 B.n616 B.n3 163.367
R1446 B.n616 B.n615 163.367
R1447 B.n615 B.n614 163.367
R1448 B.n614 B.n5 163.367
R1449 B.n610 B.n5 163.367
R1450 B.n610 B.n609 163.367
R1451 B.n609 B.n608 163.367
R1452 B.n608 B.n7 163.367
R1453 B.n604 B.n7 163.367
R1454 B.n604 B.n603 163.367
R1455 B.n603 B.n602 163.367
R1456 B.n602 B.n9 163.367
R1457 B.n598 B.n9 163.367
R1458 B.n598 B.n597 163.367
R1459 B.n597 B.n596 163.367
R1460 B.n189 B.n154 163.367
R1461 B.n193 B.n154 163.367
R1462 B.n194 B.n193 163.367
R1463 B.n195 B.n194 163.367
R1464 B.n195 B.n152 163.367
R1465 B.n199 B.n152 163.367
R1466 B.n200 B.n199 163.367
R1467 B.n201 B.n200 163.367
R1468 B.n201 B.n150 163.367
R1469 B.n205 B.n150 163.367
R1470 B.n206 B.n205 163.367
R1471 B.n207 B.n206 163.367
R1472 B.n207 B.n148 163.367
R1473 B.n211 B.n148 163.367
R1474 B.n212 B.n211 163.367
R1475 B.n213 B.n212 163.367
R1476 B.n213 B.n146 163.367
R1477 B.n217 B.n146 163.367
R1478 B.n218 B.n217 163.367
R1479 B.n219 B.n218 163.367
R1480 B.n219 B.n144 163.367
R1481 B.n223 B.n144 163.367
R1482 B.n224 B.n223 163.367
R1483 B.n225 B.n224 163.367
R1484 B.n225 B.n142 163.367
R1485 B.n229 B.n142 163.367
R1486 B.n230 B.n229 163.367
R1487 B.n231 B.n230 163.367
R1488 B.n231 B.n140 163.367
R1489 B.n235 B.n140 163.367
R1490 B.n236 B.n235 163.367
R1491 B.n237 B.n236 163.367
R1492 B.n237 B.n138 163.367
R1493 B.n241 B.n138 163.367
R1494 B.n242 B.n241 163.367
R1495 B.n243 B.n242 163.367
R1496 B.n243 B.n136 163.367
R1497 B.n247 B.n136 163.367
R1498 B.n248 B.n247 163.367
R1499 B.n249 B.n248 163.367
R1500 B.n249 B.n134 163.367
R1501 B.n253 B.n134 163.367
R1502 B.n254 B.n253 163.367
R1503 B.n255 B.n254 163.367
R1504 B.n255 B.n132 163.367
R1505 B.n259 B.n132 163.367
R1506 B.n260 B.n259 163.367
R1507 B.n261 B.n260 163.367
R1508 B.n261 B.n130 163.367
R1509 B.n265 B.n130 163.367
R1510 B.n266 B.n265 163.367
R1511 B.n267 B.n266 163.367
R1512 B.n267 B.n126 163.367
R1513 B.n272 B.n126 163.367
R1514 B.n273 B.n272 163.367
R1515 B.n274 B.n273 163.367
R1516 B.n274 B.n124 163.367
R1517 B.n278 B.n124 163.367
R1518 B.n279 B.n278 163.367
R1519 B.n280 B.n279 163.367
R1520 B.n280 B.n122 163.367
R1521 B.n284 B.n122 163.367
R1522 B.n285 B.n284 163.367
R1523 B.n285 B.n118 163.367
R1524 B.n289 B.n118 163.367
R1525 B.n290 B.n289 163.367
R1526 B.n291 B.n290 163.367
R1527 B.n291 B.n116 163.367
R1528 B.n295 B.n116 163.367
R1529 B.n296 B.n295 163.367
R1530 B.n297 B.n296 163.367
R1531 B.n297 B.n114 163.367
R1532 B.n301 B.n114 163.367
R1533 B.n302 B.n301 163.367
R1534 B.n303 B.n302 163.367
R1535 B.n303 B.n112 163.367
R1536 B.n307 B.n112 163.367
R1537 B.n308 B.n307 163.367
R1538 B.n309 B.n308 163.367
R1539 B.n309 B.n110 163.367
R1540 B.n313 B.n110 163.367
R1541 B.n314 B.n313 163.367
R1542 B.n315 B.n314 163.367
R1543 B.n315 B.n108 163.367
R1544 B.n319 B.n108 163.367
R1545 B.n320 B.n319 163.367
R1546 B.n321 B.n320 163.367
R1547 B.n321 B.n106 163.367
R1548 B.n325 B.n106 163.367
R1549 B.n326 B.n325 163.367
R1550 B.n327 B.n326 163.367
R1551 B.n327 B.n104 163.367
R1552 B.n331 B.n104 163.367
R1553 B.n332 B.n331 163.367
R1554 B.n333 B.n332 163.367
R1555 B.n333 B.n102 163.367
R1556 B.n337 B.n102 163.367
R1557 B.n338 B.n337 163.367
R1558 B.n339 B.n338 163.367
R1559 B.n339 B.n100 163.367
R1560 B.n343 B.n100 163.367
R1561 B.n344 B.n343 163.367
R1562 B.n345 B.n344 163.367
R1563 B.n345 B.n98 163.367
R1564 B.n349 B.n98 163.367
R1565 B.n350 B.n349 163.367
R1566 B.n351 B.n350 163.367
R1567 B.n351 B.n96 163.367
R1568 B.n355 B.n96 163.367
R1569 B.n356 B.n355 163.367
R1570 B.n357 B.n356 163.367
R1571 B.n357 B.n94 163.367
R1572 B.n361 B.n94 163.367
R1573 B.n362 B.n361 163.367
R1574 B.n363 B.n362 163.367
R1575 B.n367 B.n92 163.367
R1576 B.n368 B.n367 163.367
R1577 B.n369 B.n368 163.367
R1578 B.n369 B.n90 163.367
R1579 B.n373 B.n90 163.367
R1580 B.n374 B.n373 163.367
R1581 B.n375 B.n374 163.367
R1582 B.n375 B.n88 163.367
R1583 B.n379 B.n88 163.367
R1584 B.n380 B.n379 163.367
R1585 B.n381 B.n380 163.367
R1586 B.n381 B.n86 163.367
R1587 B.n385 B.n86 163.367
R1588 B.n386 B.n385 163.367
R1589 B.n387 B.n386 163.367
R1590 B.n387 B.n84 163.367
R1591 B.n391 B.n84 163.367
R1592 B.n392 B.n391 163.367
R1593 B.n393 B.n392 163.367
R1594 B.n393 B.n82 163.367
R1595 B.n397 B.n82 163.367
R1596 B.n398 B.n397 163.367
R1597 B.n399 B.n398 163.367
R1598 B.n399 B.n80 163.367
R1599 B.n403 B.n80 163.367
R1600 B.n404 B.n403 163.367
R1601 B.n405 B.n404 163.367
R1602 B.n405 B.n78 163.367
R1603 B.n409 B.n78 163.367
R1604 B.n410 B.n409 163.367
R1605 B.n411 B.n410 163.367
R1606 B.n411 B.n76 163.367
R1607 B.n415 B.n76 163.367
R1608 B.n416 B.n415 163.367
R1609 B.n417 B.n416 163.367
R1610 B.n417 B.n74 163.367
R1611 B.n592 B.n11 163.367
R1612 B.n592 B.n591 163.367
R1613 B.n591 B.n590 163.367
R1614 B.n590 B.n13 163.367
R1615 B.n586 B.n13 163.367
R1616 B.n586 B.n585 163.367
R1617 B.n585 B.n584 163.367
R1618 B.n584 B.n15 163.367
R1619 B.n580 B.n15 163.367
R1620 B.n580 B.n579 163.367
R1621 B.n579 B.n578 163.367
R1622 B.n578 B.n17 163.367
R1623 B.n574 B.n17 163.367
R1624 B.n574 B.n573 163.367
R1625 B.n573 B.n572 163.367
R1626 B.n572 B.n19 163.367
R1627 B.n568 B.n19 163.367
R1628 B.n568 B.n567 163.367
R1629 B.n567 B.n566 163.367
R1630 B.n566 B.n21 163.367
R1631 B.n562 B.n21 163.367
R1632 B.n562 B.n561 163.367
R1633 B.n561 B.n560 163.367
R1634 B.n560 B.n23 163.367
R1635 B.n556 B.n23 163.367
R1636 B.n556 B.n555 163.367
R1637 B.n555 B.n554 163.367
R1638 B.n554 B.n25 163.367
R1639 B.n550 B.n25 163.367
R1640 B.n550 B.n549 163.367
R1641 B.n549 B.n548 163.367
R1642 B.n548 B.n27 163.367
R1643 B.n544 B.n27 163.367
R1644 B.n544 B.n543 163.367
R1645 B.n543 B.n542 163.367
R1646 B.n542 B.n29 163.367
R1647 B.n538 B.n29 163.367
R1648 B.n538 B.n537 163.367
R1649 B.n537 B.n536 163.367
R1650 B.n536 B.n31 163.367
R1651 B.n532 B.n31 163.367
R1652 B.n532 B.n531 163.367
R1653 B.n531 B.n530 163.367
R1654 B.n530 B.n33 163.367
R1655 B.n526 B.n33 163.367
R1656 B.n526 B.n525 163.367
R1657 B.n525 B.n524 163.367
R1658 B.n524 B.n35 163.367
R1659 B.n520 B.n35 163.367
R1660 B.n520 B.n519 163.367
R1661 B.n519 B.n518 163.367
R1662 B.n518 B.n37 163.367
R1663 B.n513 B.n37 163.367
R1664 B.n513 B.n512 163.367
R1665 B.n512 B.n511 163.367
R1666 B.n511 B.n41 163.367
R1667 B.n507 B.n41 163.367
R1668 B.n507 B.n506 163.367
R1669 B.n506 B.n505 163.367
R1670 B.n505 B.n43 163.367
R1671 B.n501 B.n43 163.367
R1672 B.n501 B.n500 163.367
R1673 B.n500 B.n499 163.367
R1674 B.n499 B.n45 163.367
R1675 B.n495 B.n45 163.367
R1676 B.n495 B.n494 163.367
R1677 B.n494 B.n493 163.367
R1678 B.n493 B.n50 163.367
R1679 B.n489 B.n50 163.367
R1680 B.n489 B.n488 163.367
R1681 B.n488 B.n487 163.367
R1682 B.n487 B.n52 163.367
R1683 B.n483 B.n52 163.367
R1684 B.n483 B.n482 163.367
R1685 B.n482 B.n481 163.367
R1686 B.n481 B.n54 163.367
R1687 B.n477 B.n54 163.367
R1688 B.n477 B.n476 163.367
R1689 B.n476 B.n475 163.367
R1690 B.n475 B.n56 163.367
R1691 B.n471 B.n56 163.367
R1692 B.n471 B.n470 163.367
R1693 B.n470 B.n469 163.367
R1694 B.n469 B.n58 163.367
R1695 B.n465 B.n58 163.367
R1696 B.n465 B.n464 163.367
R1697 B.n464 B.n463 163.367
R1698 B.n463 B.n60 163.367
R1699 B.n459 B.n60 163.367
R1700 B.n459 B.n458 163.367
R1701 B.n458 B.n457 163.367
R1702 B.n457 B.n62 163.367
R1703 B.n453 B.n62 163.367
R1704 B.n453 B.n452 163.367
R1705 B.n452 B.n451 163.367
R1706 B.n451 B.n64 163.367
R1707 B.n447 B.n64 163.367
R1708 B.n447 B.n446 163.367
R1709 B.n446 B.n445 163.367
R1710 B.n445 B.n66 163.367
R1711 B.n441 B.n66 163.367
R1712 B.n441 B.n440 163.367
R1713 B.n440 B.n439 163.367
R1714 B.n439 B.n68 163.367
R1715 B.n435 B.n68 163.367
R1716 B.n435 B.n434 163.367
R1717 B.n434 B.n433 163.367
R1718 B.n433 B.n70 163.367
R1719 B.n429 B.n70 163.367
R1720 B.n429 B.n428 163.367
R1721 B.n428 B.n427 163.367
R1722 B.n427 B.n72 163.367
R1723 B.n423 B.n72 163.367
R1724 B.n423 B.n422 163.367
R1725 B.n422 B.n421 163.367
R1726 B.n121 B.n120 59.5399
R1727 B.n269 B.n128 59.5399
R1728 B.n515 B.n39 59.5399
R1729 B.n48 B.n47 59.5399
R1730 B.n595 B.n594 35.1225
R1731 B.n420 B.n419 35.1225
R1732 B.n365 B.n364 35.1225
R1733 B.n190 B.n155 35.1225
R1734 B.n120 B.n119 21.7217
R1735 B.n128 B.n127 21.7217
R1736 B.n39 B.n38 21.7217
R1737 B.n47 B.n46 21.7217
R1738 B B.n623 18.0485
R1739 B.n594 B.n593 10.6151
R1740 B.n593 B.n12 10.6151
R1741 B.n589 B.n12 10.6151
R1742 B.n589 B.n588 10.6151
R1743 B.n588 B.n587 10.6151
R1744 B.n587 B.n14 10.6151
R1745 B.n583 B.n14 10.6151
R1746 B.n583 B.n582 10.6151
R1747 B.n582 B.n581 10.6151
R1748 B.n581 B.n16 10.6151
R1749 B.n577 B.n16 10.6151
R1750 B.n577 B.n576 10.6151
R1751 B.n576 B.n575 10.6151
R1752 B.n575 B.n18 10.6151
R1753 B.n571 B.n18 10.6151
R1754 B.n571 B.n570 10.6151
R1755 B.n570 B.n569 10.6151
R1756 B.n569 B.n20 10.6151
R1757 B.n565 B.n20 10.6151
R1758 B.n565 B.n564 10.6151
R1759 B.n564 B.n563 10.6151
R1760 B.n563 B.n22 10.6151
R1761 B.n559 B.n22 10.6151
R1762 B.n559 B.n558 10.6151
R1763 B.n558 B.n557 10.6151
R1764 B.n557 B.n24 10.6151
R1765 B.n553 B.n24 10.6151
R1766 B.n553 B.n552 10.6151
R1767 B.n552 B.n551 10.6151
R1768 B.n551 B.n26 10.6151
R1769 B.n547 B.n26 10.6151
R1770 B.n547 B.n546 10.6151
R1771 B.n546 B.n545 10.6151
R1772 B.n545 B.n28 10.6151
R1773 B.n541 B.n28 10.6151
R1774 B.n541 B.n540 10.6151
R1775 B.n540 B.n539 10.6151
R1776 B.n539 B.n30 10.6151
R1777 B.n535 B.n30 10.6151
R1778 B.n535 B.n534 10.6151
R1779 B.n534 B.n533 10.6151
R1780 B.n533 B.n32 10.6151
R1781 B.n529 B.n32 10.6151
R1782 B.n529 B.n528 10.6151
R1783 B.n528 B.n527 10.6151
R1784 B.n527 B.n34 10.6151
R1785 B.n523 B.n34 10.6151
R1786 B.n523 B.n522 10.6151
R1787 B.n522 B.n521 10.6151
R1788 B.n521 B.n36 10.6151
R1789 B.n517 B.n36 10.6151
R1790 B.n517 B.n516 10.6151
R1791 B.n514 B.n40 10.6151
R1792 B.n510 B.n40 10.6151
R1793 B.n510 B.n509 10.6151
R1794 B.n509 B.n508 10.6151
R1795 B.n508 B.n42 10.6151
R1796 B.n504 B.n42 10.6151
R1797 B.n504 B.n503 10.6151
R1798 B.n503 B.n502 10.6151
R1799 B.n502 B.n44 10.6151
R1800 B.n498 B.n497 10.6151
R1801 B.n497 B.n496 10.6151
R1802 B.n496 B.n49 10.6151
R1803 B.n492 B.n49 10.6151
R1804 B.n492 B.n491 10.6151
R1805 B.n491 B.n490 10.6151
R1806 B.n490 B.n51 10.6151
R1807 B.n486 B.n51 10.6151
R1808 B.n486 B.n485 10.6151
R1809 B.n485 B.n484 10.6151
R1810 B.n484 B.n53 10.6151
R1811 B.n480 B.n53 10.6151
R1812 B.n480 B.n479 10.6151
R1813 B.n479 B.n478 10.6151
R1814 B.n478 B.n55 10.6151
R1815 B.n474 B.n55 10.6151
R1816 B.n474 B.n473 10.6151
R1817 B.n473 B.n472 10.6151
R1818 B.n472 B.n57 10.6151
R1819 B.n468 B.n57 10.6151
R1820 B.n468 B.n467 10.6151
R1821 B.n467 B.n466 10.6151
R1822 B.n466 B.n59 10.6151
R1823 B.n462 B.n59 10.6151
R1824 B.n462 B.n461 10.6151
R1825 B.n461 B.n460 10.6151
R1826 B.n460 B.n61 10.6151
R1827 B.n456 B.n61 10.6151
R1828 B.n456 B.n455 10.6151
R1829 B.n455 B.n454 10.6151
R1830 B.n454 B.n63 10.6151
R1831 B.n450 B.n63 10.6151
R1832 B.n450 B.n449 10.6151
R1833 B.n449 B.n448 10.6151
R1834 B.n448 B.n65 10.6151
R1835 B.n444 B.n65 10.6151
R1836 B.n444 B.n443 10.6151
R1837 B.n443 B.n442 10.6151
R1838 B.n442 B.n67 10.6151
R1839 B.n438 B.n67 10.6151
R1840 B.n438 B.n437 10.6151
R1841 B.n437 B.n436 10.6151
R1842 B.n436 B.n69 10.6151
R1843 B.n432 B.n69 10.6151
R1844 B.n432 B.n431 10.6151
R1845 B.n431 B.n430 10.6151
R1846 B.n430 B.n71 10.6151
R1847 B.n426 B.n71 10.6151
R1848 B.n426 B.n425 10.6151
R1849 B.n425 B.n424 10.6151
R1850 B.n424 B.n73 10.6151
R1851 B.n420 B.n73 10.6151
R1852 B.n366 B.n365 10.6151
R1853 B.n366 B.n91 10.6151
R1854 B.n370 B.n91 10.6151
R1855 B.n371 B.n370 10.6151
R1856 B.n372 B.n371 10.6151
R1857 B.n372 B.n89 10.6151
R1858 B.n376 B.n89 10.6151
R1859 B.n377 B.n376 10.6151
R1860 B.n378 B.n377 10.6151
R1861 B.n378 B.n87 10.6151
R1862 B.n382 B.n87 10.6151
R1863 B.n383 B.n382 10.6151
R1864 B.n384 B.n383 10.6151
R1865 B.n384 B.n85 10.6151
R1866 B.n388 B.n85 10.6151
R1867 B.n389 B.n388 10.6151
R1868 B.n390 B.n389 10.6151
R1869 B.n390 B.n83 10.6151
R1870 B.n394 B.n83 10.6151
R1871 B.n395 B.n394 10.6151
R1872 B.n396 B.n395 10.6151
R1873 B.n396 B.n81 10.6151
R1874 B.n400 B.n81 10.6151
R1875 B.n401 B.n400 10.6151
R1876 B.n402 B.n401 10.6151
R1877 B.n402 B.n79 10.6151
R1878 B.n406 B.n79 10.6151
R1879 B.n407 B.n406 10.6151
R1880 B.n408 B.n407 10.6151
R1881 B.n408 B.n77 10.6151
R1882 B.n412 B.n77 10.6151
R1883 B.n413 B.n412 10.6151
R1884 B.n414 B.n413 10.6151
R1885 B.n414 B.n75 10.6151
R1886 B.n418 B.n75 10.6151
R1887 B.n419 B.n418 10.6151
R1888 B.n191 B.n190 10.6151
R1889 B.n192 B.n191 10.6151
R1890 B.n192 B.n153 10.6151
R1891 B.n196 B.n153 10.6151
R1892 B.n197 B.n196 10.6151
R1893 B.n198 B.n197 10.6151
R1894 B.n198 B.n151 10.6151
R1895 B.n202 B.n151 10.6151
R1896 B.n203 B.n202 10.6151
R1897 B.n204 B.n203 10.6151
R1898 B.n204 B.n149 10.6151
R1899 B.n208 B.n149 10.6151
R1900 B.n209 B.n208 10.6151
R1901 B.n210 B.n209 10.6151
R1902 B.n210 B.n147 10.6151
R1903 B.n214 B.n147 10.6151
R1904 B.n215 B.n214 10.6151
R1905 B.n216 B.n215 10.6151
R1906 B.n216 B.n145 10.6151
R1907 B.n220 B.n145 10.6151
R1908 B.n221 B.n220 10.6151
R1909 B.n222 B.n221 10.6151
R1910 B.n222 B.n143 10.6151
R1911 B.n226 B.n143 10.6151
R1912 B.n227 B.n226 10.6151
R1913 B.n228 B.n227 10.6151
R1914 B.n228 B.n141 10.6151
R1915 B.n232 B.n141 10.6151
R1916 B.n233 B.n232 10.6151
R1917 B.n234 B.n233 10.6151
R1918 B.n234 B.n139 10.6151
R1919 B.n238 B.n139 10.6151
R1920 B.n239 B.n238 10.6151
R1921 B.n240 B.n239 10.6151
R1922 B.n240 B.n137 10.6151
R1923 B.n244 B.n137 10.6151
R1924 B.n245 B.n244 10.6151
R1925 B.n246 B.n245 10.6151
R1926 B.n246 B.n135 10.6151
R1927 B.n250 B.n135 10.6151
R1928 B.n251 B.n250 10.6151
R1929 B.n252 B.n251 10.6151
R1930 B.n252 B.n133 10.6151
R1931 B.n256 B.n133 10.6151
R1932 B.n257 B.n256 10.6151
R1933 B.n258 B.n257 10.6151
R1934 B.n258 B.n131 10.6151
R1935 B.n262 B.n131 10.6151
R1936 B.n263 B.n262 10.6151
R1937 B.n264 B.n263 10.6151
R1938 B.n264 B.n129 10.6151
R1939 B.n268 B.n129 10.6151
R1940 B.n271 B.n270 10.6151
R1941 B.n271 B.n125 10.6151
R1942 B.n275 B.n125 10.6151
R1943 B.n276 B.n275 10.6151
R1944 B.n277 B.n276 10.6151
R1945 B.n277 B.n123 10.6151
R1946 B.n281 B.n123 10.6151
R1947 B.n282 B.n281 10.6151
R1948 B.n283 B.n282 10.6151
R1949 B.n287 B.n286 10.6151
R1950 B.n288 B.n287 10.6151
R1951 B.n288 B.n117 10.6151
R1952 B.n292 B.n117 10.6151
R1953 B.n293 B.n292 10.6151
R1954 B.n294 B.n293 10.6151
R1955 B.n294 B.n115 10.6151
R1956 B.n298 B.n115 10.6151
R1957 B.n299 B.n298 10.6151
R1958 B.n300 B.n299 10.6151
R1959 B.n300 B.n113 10.6151
R1960 B.n304 B.n113 10.6151
R1961 B.n305 B.n304 10.6151
R1962 B.n306 B.n305 10.6151
R1963 B.n306 B.n111 10.6151
R1964 B.n310 B.n111 10.6151
R1965 B.n311 B.n310 10.6151
R1966 B.n312 B.n311 10.6151
R1967 B.n312 B.n109 10.6151
R1968 B.n316 B.n109 10.6151
R1969 B.n317 B.n316 10.6151
R1970 B.n318 B.n317 10.6151
R1971 B.n318 B.n107 10.6151
R1972 B.n322 B.n107 10.6151
R1973 B.n323 B.n322 10.6151
R1974 B.n324 B.n323 10.6151
R1975 B.n324 B.n105 10.6151
R1976 B.n328 B.n105 10.6151
R1977 B.n329 B.n328 10.6151
R1978 B.n330 B.n329 10.6151
R1979 B.n330 B.n103 10.6151
R1980 B.n334 B.n103 10.6151
R1981 B.n335 B.n334 10.6151
R1982 B.n336 B.n335 10.6151
R1983 B.n336 B.n101 10.6151
R1984 B.n340 B.n101 10.6151
R1985 B.n341 B.n340 10.6151
R1986 B.n342 B.n341 10.6151
R1987 B.n342 B.n99 10.6151
R1988 B.n346 B.n99 10.6151
R1989 B.n347 B.n346 10.6151
R1990 B.n348 B.n347 10.6151
R1991 B.n348 B.n97 10.6151
R1992 B.n352 B.n97 10.6151
R1993 B.n353 B.n352 10.6151
R1994 B.n354 B.n353 10.6151
R1995 B.n354 B.n95 10.6151
R1996 B.n358 B.n95 10.6151
R1997 B.n359 B.n358 10.6151
R1998 B.n360 B.n359 10.6151
R1999 B.n360 B.n93 10.6151
R2000 B.n364 B.n93 10.6151
R2001 B.n186 B.n155 10.6151
R2002 B.n186 B.n185 10.6151
R2003 B.n185 B.n184 10.6151
R2004 B.n184 B.n157 10.6151
R2005 B.n180 B.n157 10.6151
R2006 B.n180 B.n179 10.6151
R2007 B.n179 B.n178 10.6151
R2008 B.n178 B.n159 10.6151
R2009 B.n174 B.n159 10.6151
R2010 B.n174 B.n173 10.6151
R2011 B.n173 B.n172 10.6151
R2012 B.n172 B.n161 10.6151
R2013 B.n168 B.n161 10.6151
R2014 B.n168 B.n167 10.6151
R2015 B.n167 B.n166 10.6151
R2016 B.n166 B.n163 10.6151
R2017 B.n163 B.n0 10.6151
R2018 B.n619 B.n1 10.6151
R2019 B.n619 B.n618 10.6151
R2020 B.n618 B.n617 10.6151
R2021 B.n617 B.n4 10.6151
R2022 B.n613 B.n4 10.6151
R2023 B.n613 B.n612 10.6151
R2024 B.n612 B.n611 10.6151
R2025 B.n611 B.n6 10.6151
R2026 B.n607 B.n6 10.6151
R2027 B.n607 B.n606 10.6151
R2028 B.n606 B.n605 10.6151
R2029 B.n605 B.n8 10.6151
R2030 B.n601 B.n8 10.6151
R2031 B.n601 B.n600 10.6151
R2032 B.n600 B.n599 10.6151
R2033 B.n599 B.n10 10.6151
R2034 B.n595 B.n10 10.6151
R2035 B.n516 B.n515 9.36635
R2036 B.n498 B.n48 9.36635
R2037 B.n269 B.n268 9.36635
R2038 B.n286 B.n121 9.36635
R2039 B.n623 B.n0 2.81026
R2040 B.n623 B.n1 2.81026
R2041 B.n515 B.n514 1.24928
R2042 B.n48 B.n44 1.24928
R2043 B.n270 B.n269 1.24928
R2044 B.n283 B.n121 1.24928
R2045 VP.n1 VP.t0 560.043
R2046 VP.n1 VP.t3 559.994
R2047 VP.n3 VP.t2 539.048
R2048 VP.n5 VP.t1 539.048
R2049 VP.n6 VP.n5 161.3
R2050 VP.n4 VP.n0 161.3
R2051 VP.n3 VP.n2 161.3
R2052 VP.n2 VP.n1 88.4651
R2053 VP.n4 VP.n3 24.1005
R2054 VP.n5 VP.n4 24.1005
R2055 VP.n2 VP.n0 0.189894
R2056 VP.n6 VP.n0 0.189894
R2057 VP VP.n6 0.0516364
R2058 VDD1 VDD1.n1 109.787
R2059 VDD1 VDD1.n0 68.8904
R2060 VDD1.n0 VDD1.t3 2.02826
R2061 VDD1.n0 VDD1.t0 2.02826
R2062 VDD1.n1 VDD1.t1 2.02826
R2063 VDD1.n1 VDD1.t2 2.02826
C0 VTAIL VDD1 8.1878f
C1 VTAIL w_n1642_n4174# 5.11715f
C2 VN VP 5.63223f
C3 VTAIL VDD2 8.229871f
C4 VP VDD1 4.48862f
C5 VP w_n1642_n4174# 2.72842f
C6 VP VDD2 0.278939f
C7 VTAIL B 4.99139f
C8 VN VDD1 0.147171f
C9 VN w_n1642_n4174# 2.52191f
C10 VN VDD2 4.35714f
C11 B VP 1.14544f
C12 w_n1642_n4174# VDD1 1.18938f
C13 VDD2 VDD1 0.587163f
C14 VDD2 w_n1642_n4174# 1.20572f
C15 VTAIL VP 3.83274f
C16 B VN 0.811177f
C17 B VDD1 1.05066f
C18 B w_n1642_n4174# 8.1482f
C19 VTAIL VN 3.81863f
C20 B VDD2 1.07347f
C21 VDD2 VSUBS 0.785947f
C22 VDD1 VSUBS 5.551985f
C23 VTAIL VSUBS 1.077743f
C24 VN VSUBS 6.08383f
C25 VP VSUBS 1.489189f
C26 B VSUBS 3.037818f
C27 w_n1642_n4174# VSUBS 83.9587f
C28 VDD1.t3 VSUBS 0.353741f
C29 VDD1.t0 VSUBS 0.353741f
C30 VDD1.n0 VSUBS 2.89102f
C31 VDD1.t1 VSUBS 0.353741f
C32 VDD1.t2 VSUBS 0.353741f
C33 VDD1.n1 VSUBS 3.73682f
C34 VP.n0 VSUBS 0.056714f
C35 VP.t3 VSUBS 2.06865f
C36 VP.t0 VSUBS 2.06873f
C37 VP.n1 VSUBS 2.80865f
C38 VP.n2 VSUBS 3.8857f
C39 VP.t2 VSUBS 2.03954f
C40 VP.n3 VSUBS 0.774281f
C41 VP.n4 VSUBS 0.01287f
C42 VP.t1 VSUBS 2.03954f
C43 VP.n5 VSUBS 0.774281f
C44 VP.n6 VSUBS 0.043951f
C45 B.n0 VSUBS 0.00488f
C46 B.n1 VSUBS 0.00488f
C47 B.n2 VSUBS 0.007718f
C48 B.n3 VSUBS 0.007718f
C49 B.n4 VSUBS 0.007718f
C50 B.n5 VSUBS 0.007718f
C51 B.n6 VSUBS 0.007718f
C52 B.n7 VSUBS 0.007718f
C53 B.n8 VSUBS 0.007718f
C54 B.n9 VSUBS 0.007718f
C55 B.n10 VSUBS 0.007718f
C56 B.n11 VSUBS 0.019171f
C57 B.n12 VSUBS 0.007718f
C58 B.n13 VSUBS 0.007718f
C59 B.n14 VSUBS 0.007718f
C60 B.n15 VSUBS 0.007718f
C61 B.n16 VSUBS 0.007718f
C62 B.n17 VSUBS 0.007718f
C63 B.n18 VSUBS 0.007718f
C64 B.n19 VSUBS 0.007718f
C65 B.n20 VSUBS 0.007718f
C66 B.n21 VSUBS 0.007718f
C67 B.n22 VSUBS 0.007718f
C68 B.n23 VSUBS 0.007718f
C69 B.n24 VSUBS 0.007718f
C70 B.n25 VSUBS 0.007718f
C71 B.n26 VSUBS 0.007718f
C72 B.n27 VSUBS 0.007718f
C73 B.n28 VSUBS 0.007718f
C74 B.n29 VSUBS 0.007718f
C75 B.n30 VSUBS 0.007718f
C76 B.n31 VSUBS 0.007718f
C77 B.n32 VSUBS 0.007718f
C78 B.n33 VSUBS 0.007718f
C79 B.n34 VSUBS 0.007718f
C80 B.n35 VSUBS 0.007718f
C81 B.n36 VSUBS 0.007718f
C82 B.n37 VSUBS 0.007718f
C83 B.t11 VSUBS 0.334844f
C84 B.t10 VSUBS 0.349495f
C85 B.t9 VSUBS 0.57059f
C86 B.n38 VSUBS 0.448977f
C87 B.n39 VSUBS 0.327851f
C88 B.n40 VSUBS 0.007718f
C89 B.n41 VSUBS 0.007718f
C90 B.n42 VSUBS 0.007718f
C91 B.n43 VSUBS 0.007718f
C92 B.n44 VSUBS 0.004313f
C93 B.n45 VSUBS 0.007718f
C94 B.t8 VSUBS 0.334848f
C95 B.t7 VSUBS 0.349498f
C96 B.t6 VSUBS 0.57059f
C97 B.n46 VSUBS 0.448973f
C98 B.n47 VSUBS 0.327847f
C99 B.n48 VSUBS 0.017881f
C100 B.n49 VSUBS 0.007718f
C101 B.n50 VSUBS 0.007718f
C102 B.n51 VSUBS 0.007718f
C103 B.n52 VSUBS 0.007718f
C104 B.n53 VSUBS 0.007718f
C105 B.n54 VSUBS 0.007718f
C106 B.n55 VSUBS 0.007718f
C107 B.n56 VSUBS 0.007718f
C108 B.n57 VSUBS 0.007718f
C109 B.n58 VSUBS 0.007718f
C110 B.n59 VSUBS 0.007718f
C111 B.n60 VSUBS 0.007718f
C112 B.n61 VSUBS 0.007718f
C113 B.n62 VSUBS 0.007718f
C114 B.n63 VSUBS 0.007718f
C115 B.n64 VSUBS 0.007718f
C116 B.n65 VSUBS 0.007718f
C117 B.n66 VSUBS 0.007718f
C118 B.n67 VSUBS 0.007718f
C119 B.n68 VSUBS 0.007718f
C120 B.n69 VSUBS 0.007718f
C121 B.n70 VSUBS 0.007718f
C122 B.n71 VSUBS 0.007718f
C123 B.n72 VSUBS 0.007718f
C124 B.n73 VSUBS 0.007718f
C125 B.n74 VSUBS 0.018737f
C126 B.n75 VSUBS 0.007718f
C127 B.n76 VSUBS 0.007718f
C128 B.n77 VSUBS 0.007718f
C129 B.n78 VSUBS 0.007718f
C130 B.n79 VSUBS 0.007718f
C131 B.n80 VSUBS 0.007718f
C132 B.n81 VSUBS 0.007718f
C133 B.n82 VSUBS 0.007718f
C134 B.n83 VSUBS 0.007718f
C135 B.n84 VSUBS 0.007718f
C136 B.n85 VSUBS 0.007718f
C137 B.n86 VSUBS 0.007718f
C138 B.n87 VSUBS 0.007718f
C139 B.n88 VSUBS 0.007718f
C140 B.n89 VSUBS 0.007718f
C141 B.n90 VSUBS 0.007718f
C142 B.n91 VSUBS 0.007718f
C143 B.n92 VSUBS 0.018737f
C144 B.n93 VSUBS 0.007718f
C145 B.n94 VSUBS 0.007718f
C146 B.n95 VSUBS 0.007718f
C147 B.n96 VSUBS 0.007718f
C148 B.n97 VSUBS 0.007718f
C149 B.n98 VSUBS 0.007718f
C150 B.n99 VSUBS 0.007718f
C151 B.n100 VSUBS 0.007718f
C152 B.n101 VSUBS 0.007718f
C153 B.n102 VSUBS 0.007718f
C154 B.n103 VSUBS 0.007718f
C155 B.n104 VSUBS 0.007718f
C156 B.n105 VSUBS 0.007718f
C157 B.n106 VSUBS 0.007718f
C158 B.n107 VSUBS 0.007718f
C159 B.n108 VSUBS 0.007718f
C160 B.n109 VSUBS 0.007718f
C161 B.n110 VSUBS 0.007718f
C162 B.n111 VSUBS 0.007718f
C163 B.n112 VSUBS 0.007718f
C164 B.n113 VSUBS 0.007718f
C165 B.n114 VSUBS 0.007718f
C166 B.n115 VSUBS 0.007718f
C167 B.n116 VSUBS 0.007718f
C168 B.n117 VSUBS 0.007718f
C169 B.n118 VSUBS 0.007718f
C170 B.t1 VSUBS 0.334848f
C171 B.t2 VSUBS 0.349498f
C172 B.t0 VSUBS 0.57059f
C173 B.n119 VSUBS 0.448973f
C174 B.n120 VSUBS 0.327847f
C175 B.n121 VSUBS 0.017881f
C176 B.n122 VSUBS 0.007718f
C177 B.n123 VSUBS 0.007718f
C178 B.n124 VSUBS 0.007718f
C179 B.n125 VSUBS 0.007718f
C180 B.n126 VSUBS 0.007718f
C181 B.t4 VSUBS 0.334844f
C182 B.t5 VSUBS 0.349495f
C183 B.t3 VSUBS 0.57059f
C184 B.n127 VSUBS 0.448977f
C185 B.n128 VSUBS 0.327851f
C186 B.n129 VSUBS 0.007718f
C187 B.n130 VSUBS 0.007718f
C188 B.n131 VSUBS 0.007718f
C189 B.n132 VSUBS 0.007718f
C190 B.n133 VSUBS 0.007718f
C191 B.n134 VSUBS 0.007718f
C192 B.n135 VSUBS 0.007718f
C193 B.n136 VSUBS 0.007718f
C194 B.n137 VSUBS 0.007718f
C195 B.n138 VSUBS 0.007718f
C196 B.n139 VSUBS 0.007718f
C197 B.n140 VSUBS 0.007718f
C198 B.n141 VSUBS 0.007718f
C199 B.n142 VSUBS 0.007718f
C200 B.n143 VSUBS 0.007718f
C201 B.n144 VSUBS 0.007718f
C202 B.n145 VSUBS 0.007718f
C203 B.n146 VSUBS 0.007718f
C204 B.n147 VSUBS 0.007718f
C205 B.n148 VSUBS 0.007718f
C206 B.n149 VSUBS 0.007718f
C207 B.n150 VSUBS 0.007718f
C208 B.n151 VSUBS 0.007718f
C209 B.n152 VSUBS 0.007718f
C210 B.n153 VSUBS 0.007718f
C211 B.n154 VSUBS 0.007718f
C212 B.n155 VSUBS 0.018737f
C213 B.n156 VSUBS 0.007718f
C214 B.n157 VSUBS 0.007718f
C215 B.n158 VSUBS 0.007718f
C216 B.n159 VSUBS 0.007718f
C217 B.n160 VSUBS 0.007718f
C218 B.n161 VSUBS 0.007718f
C219 B.n162 VSUBS 0.007718f
C220 B.n163 VSUBS 0.007718f
C221 B.n164 VSUBS 0.007718f
C222 B.n165 VSUBS 0.007718f
C223 B.n166 VSUBS 0.007718f
C224 B.n167 VSUBS 0.007718f
C225 B.n168 VSUBS 0.007718f
C226 B.n169 VSUBS 0.007718f
C227 B.n170 VSUBS 0.007718f
C228 B.n171 VSUBS 0.007718f
C229 B.n172 VSUBS 0.007718f
C230 B.n173 VSUBS 0.007718f
C231 B.n174 VSUBS 0.007718f
C232 B.n175 VSUBS 0.007718f
C233 B.n176 VSUBS 0.007718f
C234 B.n177 VSUBS 0.007718f
C235 B.n178 VSUBS 0.007718f
C236 B.n179 VSUBS 0.007718f
C237 B.n180 VSUBS 0.007718f
C238 B.n181 VSUBS 0.007718f
C239 B.n182 VSUBS 0.007718f
C240 B.n183 VSUBS 0.007718f
C241 B.n184 VSUBS 0.007718f
C242 B.n185 VSUBS 0.007718f
C243 B.n186 VSUBS 0.007718f
C244 B.n187 VSUBS 0.007718f
C245 B.n188 VSUBS 0.018737f
C246 B.n189 VSUBS 0.019171f
C247 B.n190 VSUBS 0.019171f
C248 B.n191 VSUBS 0.007718f
C249 B.n192 VSUBS 0.007718f
C250 B.n193 VSUBS 0.007718f
C251 B.n194 VSUBS 0.007718f
C252 B.n195 VSUBS 0.007718f
C253 B.n196 VSUBS 0.007718f
C254 B.n197 VSUBS 0.007718f
C255 B.n198 VSUBS 0.007718f
C256 B.n199 VSUBS 0.007718f
C257 B.n200 VSUBS 0.007718f
C258 B.n201 VSUBS 0.007718f
C259 B.n202 VSUBS 0.007718f
C260 B.n203 VSUBS 0.007718f
C261 B.n204 VSUBS 0.007718f
C262 B.n205 VSUBS 0.007718f
C263 B.n206 VSUBS 0.007718f
C264 B.n207 VSUBS 0.007718f
C265 B.n208 VSUBS 0.007718f
C266 B.n209 VSUBS 0.007718f
C267 B.n210 VSUBS 0.007718f
C268 B.n211 VSUBS 0.007718f
C269 B.n212 VSUBS 0.007718f
C270 B.n213 VSUBS 0.007718f
C271 B.n214 VSUBS 0.007718f
C272 B.n215 VSUBS 0.007718f
C273 B.n216 VSUBS 0.007718f
C274 B.n217 VSUBS 0.007718f
C275 B.n218 VSUBS 0.007718f
C276 B.n219 VSUBS 0.007718f
C277 B.n220 VSUBS 0.007718f
C278 B.n221 VSUBS 0.007718f
C279 B.n222 VSUBS 0.007718f
C280 B.n223 VSUBS 0.007718f
C281 B.n224 VSUBS 0.007718f
C282 B.n225 VSUBS 0.007718f
C283 B.n226 VSUBS 0.007718f
C284 B.n227 VSUBS 0.007718f
C285 B.n228 VSUBS 0.007718f
C286 B.n229 VSUBS 0.007718f
C287 B.n230 VSUBS 0.007718f
C288 B.n231 VSUBS 0.007718f
C289 B.n232 VSUBS 0.007718f
C290 B.n233 VSUBS 0.007718f
C291 B.n234 VSUBS 0.007718f
C292 B.n235 VSUBS 0.007718f
C293 B.n236 VSUBS 0.007718f
C294 B.n237 VSUBS 0.007718f
C295 B.n238 VSUBS 0.007718f
C296 B.n239 VSUBS 0.007718f
C297 B.n240 VSUBS 0.007718f
C298 B.n241 VSUBS 0.007718f
C299 B.n242 VSUBS 0.007718f
C300 B.n243 VSUBS 0.007718f
C301 B.n244 VSUBS 0.007718f
C302 B.n245 VSUBS 0.007718f
C303 B.n246 VSUBS 0.007718f
C304 B.n247 VSUBS 0.007718f
C305 B.n248 VSUBS 0.007718f
C306 B.n249 VSUBS 0.007718f
C307 B.n250 VSUBS 0.007718f
C308 B.n251 VSUBS 0.007718f
C309 B.n252 VSUBS 0.007718f
C310 B.n253 VSUBS 0.007718f
C311 B.n254 VSUBS 0.007718f
C312 B.n255 VSUBS 0.007718f
C313 B.n256 VSUBS 0.007718f
C314 B.n257 VSUBS 0.007718f
C315 B.n258 VSUBS 0.007718f
C316 B.n259 VSUBS 0.007718f
C317 B.n260 VSUBS 0.007718f
C318 B.n261 VSUBS 0.007718f
C319 B.n262 VSUBS 0.007718f
C320 B.n263 VSUBS 0.007718f
C321 B.n264 VSUBS 0.007718f
C322 B.n265 VSUBS 0.007718f
C323 B.n266 VSUBS 0.007718f
C324 B.n267 VSUBS 0.007718f
C325 B.n268 VSUBS 0.007264f
C326 B.n269 VSUBS 0.017881f
C327 B.n270 VSUBS 0.004313f
C328 B.n271 VSUBS 0.007718f
C329 B.n272 VSUBS 0.007718f
C330 B.n273 VSUBS 0.007718f
C331 B.n274 VSUBS 0.007718f
C332 B.n275 VSUBS 0.007718f
C333 B.n276 VSUBS 0.007718f
C334 B.n277 VSUBS 0.007718f
C335 B.n278 VSUBS 0.007718f
C336 B.n279 VSUBS 0.007718f
C337 B.n280 VSUBS 0.007718f
C338 B.n281 VSUBS 0.007718f
C339 B.n282 VSUBS 0.007718f
C340 B.n283 VSUBS 0.004313f
C341 B.n284 VSUBS 0.007718f
C342 B.n285 VSUBS 0.007718f
C343 B.n286 VSUBS 0.007264f
C344 B.n287 VSUBS 0.007718f
C345 B.n288 VSUBS 0.007718f
C346 B.n289 VSUBS 0.007718f
C347 B.n290 VSUBS 0.007718f
C348 B.n291 VSUBS 0.007718f
C349 B.n292 VSUBS 0.007718f
C350 B.n293 VSUBS 0.007718f
C351 B.n294 VSUBS 0.007718f
C352 B.n295 VSUBS 0.007718f
C353 B.n296 VSUBS 0.007718f
C354 B.n297 VSUBS 0.007718f
C355 B.n298 VSUBS 0.007718f
C356 B.n299 VSUBS 0.007718f
C357 B.n300 VSUBS 0.007718f
C358 B.n301 VSUBS 0.007718f
C359 B.n302 VSUBS 0.007718f
C360 B.n303 VSUBS 0.007718f
C361 B.n304 VSUBS 0.007718f
C362 B.n305 VSUBS 0.007718f
C363 B.n306 VSUBS 0.007718f
C364 B.n307 VSUBS 0.007718f
C365 B.n308 VSUBS 0.007718f
C366 B.n309 VSUBS 0.007718f
C367 B.n310 VSUBS 0.007718f
C368 B.n311 VSUBS 0.007718f
C369 B.n312 VSUBS 0.007718f
C370 B.n313 VSUBS 0.007718f
C371 B.n314 VSUBS 0.007718f
C372 B.n315 VSUBS 0.007718f
C373 B.n316 VSUBS 0.007718f
C374 B.n317 VSUBS 0.007718f
C375 B.n318 VSUBS 0.007718f
C376 B.n319 VSUBS 0.007718f
C377 B.n320 VSUBS 0.007718f
C378 B.n321 VSUBS 0.007718f
C379 B.n322 VSUBS 0.007718f
C380 B.n323 VSUBS 0.007718f
C381 B.n324 VSUBS 0.007718f
C382 B.n325 VSUBS 0.007718f
C383 B.n326 VSUBS 0.007718f
C384 B.n327 VSUBS 0.007718f
C385 B.n328 VSUBS 0.007718f
C386 B.n329 VSUBS 0.007718f
C387 B.n330 VSUBS 0.007718f
C388 B.n331 VSUBS 0.007718f
C389 B.n332 VSUBS 0.007718f
C390 B.n333 VSUBS 0.007718f
C391 B.n334 VSUBS 0.007718f
C392 B.n335 VSUBS 0.007718f
C393 B.n336 VSUBS 0.007718f
C394 B.n337 VSUBS 0.007718f
C395 B.n338 VSUBS 0.007718f
C396 B.n339 VSUBS 0.007718f
C397 B.n340 VSUBS 0.007718f
C398 B.n341 VSUBS 0.007718f
C399 B.n342 VSUBS 0.007718f
C400 B.n343 VSUBS 0.007718f
C401 B.n344 VSUBS 0.007718f
C402 B.n345 VSUBS 0.007718f
C403 B.n346 VSUBS 0.007718f
C404 B.n347 VSUBS 0.007718f
C405 B.n348 VSUBS 0.007718f
C406 B.n349 VSUBS 0.007718f
C407 B.n350 VSUBS 0.007718f
C408 B.n351 VSUBS 0.007718f
C409 B.n352 VSUBS 0.007718f
C410 B.n353 VSUBS 0.007718f
C411 B.n354 VSUBS 0.007718f
C412 B.n355 VSUBS 0.007718f
C413 B.n356 VSUBS 0.007718f
C414 B.n357 VSUBS 0.007718f
C415 B.n358 VSUBS 0.007718f
C416 B.n359 VSUBS 0.007718f
C417 B.n360 VSUBS 0.007718f
C418 B.n361 VSUBS 0.007718f
C419 B.n362 VSUBS 0.007718f
C420 B.n363 VSUBS 0.019171f
C421 B.n364 VSUBS 0.019171f
C422 B.n365 VSUBS 0.018737f
C423 B.n366 VSUBS 0.007718f
C424 B.n367 VSUBS 0.007718f
C425 B.n368 VSUBS 0.007718f
C426 B.n369 VSUBS 0.007718f
C427 B.n370 VSUBS 0.007718f
C428 B.n371 VSUBS 0.007718f
C429 B.n372 VSUBS 0.007718f
C430 B.n373 VSUBS 0.007718f
C431 B.n374 VSUBS 0.007718f
C432 B.n375 VSUBS 0.007718f
C433 B.n376 VSUBS 0.007718f
C434 B.n377 VSUBS 0.007718f
C435 B.n378 VSUBS 0.007718f
C436 B.n379 VSUBS 0.007718f
C437 B.n380 VSUBS 0.007718f
C438 B.n381 VSUBS 0.007718f
C439 B.n382 VSUBS 0.007718f
C440 B.n383 VSUBS 0.007718f
C441 B.n384 VSUBS 0.007718f
C442 B.n385 VSUBS 0.007718f
C443 B.n386 VSUBS 0.007718f
C444 B.n387 VSUBS 0.007718f
C445 B.n388 VSUBS 0.007718f
C446 B.n389 VSUBS 0.007718f
C447 B.n390 VSUBS 0.007718f
C448 B.n391 VSUBS 0.007718f
C449 B.n392 VSUBS 0.007718f
C450 B.n393 VSUBS 0.007718f
C451 B.n394 VSUBS 0.007718f
C452 B.n395 VSUBS 0.007718f
C453 B.n396 VSUBS 0.007718f
C454 B.n397 VSUBS 0.007718f
C455 B.n398 VSUBS 0.007718f
C456 B.n399 VSUBS 0.007718f
C457 B.n400 VSUBS 0.007718f
C458 B.n401 VSUBS 0.007718f
C459 B.n402 VSUBS 0.007718f
C460 B.n403 VSUBS 0.007718f
C461 B.n404 VSUBS 0.007718f
C462 B.n405 VSUBS 0.007718f
C463 B.n406 VSUBS 0.007718f
C464 B.n407 VSUBS 0.007718f
C465 B.n408 VSUBS 0.007718f
C466 B.n409 VSUBS 0.007718f
C467 B.n410 VSUBS 0.007718f
C468 B.n411 VSUBS 0.007718f
C469 B.n412 VSUBS 0.007718f
C470 B.n413 VSUBS 0.007718f
C471 B.n414 VSUBS 0.007718f
C472 B.n415 VSUBS 0.007718f
C473 B.n416 VSUBS 0.007718f
C474 B.n417 VSUBS 0.007718f
C475 B.n418 VSUBS 0.007718f
C476 B.n419 VSUBS 0.019585f
C477 B.n420 VSUBS 0.018323f
C478 B.n421 VSUBS 0.019171f
C479 B.n422 VSUBS 0.007718f
C480 B.n423 VSUBS 0.007718f
C481 B.n424 VSUBS 0.007718f
C482 B.n425 VSUBS 0.007718f
C483 B.n426 VSUBS 0.007718f
C484 B.n427 VSUBS 0.007718f
C485 B.n428 VSUBS 0.007718f
C486 B.n429 VSUBS 0.007718f
C487 B.n430 VSUBS 0.007718f
C488 B.n431 VSUBS 0.007718f
C489 B.n432 VSUBS 0.007718f
C490 B.n433 VSUBS 0.007718f
C491 B.n434 VSUBS 0.007718f
C492 B.n435 VSUBS 0.007718f
C493 B.n436 VSUBS 0.007718f
C494 B.n437 VSUBS 0.007718f
C495 B.n438 VSUBS 0.007718f
C496 B.n439 VSUBS 0.007718f
C497 B.n440 VSUBS 0.007718f
C498 B.n441 VSUBS 0.007718f
C499 B.n442 VSUBS 0.007718f
C500 B.n443 VSUBS 0.007718f
C501 B.n444 VSUBS 0.007718f
C502 B.n445 VSUBS 0.007718f
C503 B.n446 VSUBS 0.007718f
C504 B.n447 VSUBS 0.007718f
C505 B.n448 VSUBS 0.007718f
C506 B.n449 VSUBS 0.007718f
C507 B.n450 VSUBS 0.007718f
C508 B.n451 VSUBS 0.007718f
C509 B.n452 VSUBS 0.007718f
C510 B.n453 VSUBS 0.007718f
C511 B.n454 VSUBS 0.007718f
C512 B.n455 VSUBS 0.007718f
C513 B.n456 VSUBS 0.007718f
C514 B.n457 VSUBS 0.007718f
C515 B.n458 VSUBS 0.007718f
C516 B.n459 VSUBS 0.007718f
C517 B.n460 VSUBS 0.007718f
C518 B.n461 VSUBS 0.007718f
C519 B.n462 VSUBS 0.007718f
C520 B.n463 VSUBS 0.007718f
C521 B.n464 VSUBS 0.007718f
C522 B.n465 VSUBS 0.007718f
C523 B.n466 VSUBS 0.007718f
C524 B.n467 VSUBS 0.007718f
C525 B.n468 VSUBS 0.007718f
C526 B.n469 VSUBS 0.007718f
C527 B.n470 VSUBS 0.007718f
C528 B.n471 VSUBS 0.007718f
C529 B.n472 VSUBS 0.007718f
C530 B.n473 VSUBS 0.007718f
C531 B.n474 VSUBS 0.007718f
C532 B.n475 VSUBS 0.007718f
C533 B.n476 VSUBS 0.007718f
C534 B.n477 VSUBS 0.007718f
C535 B.n478 VSUBS 0.007718f
C536 B.n479 VSUBS 0.007718f
C537 B.n480 VSUBS 0.007718f
C538 B.n481 VSUBS 0.007718f
C539 B.n482 VSUBS 0.007718f
C540 B.n483 VSUBS 0.007718f
C541 B.n484 VSUBS 0.007718f
C542 B.n485 VSUBS 0.007718f
C543 B.n486 VSUBS 0.007718f
C544 B.n487 VSUBS 0.007718f
C545 B.n488 VSUBS 0.007718f
C546 B.n489 VSUBS 0.007718f
C547 B.n490 VSUBS 0.007718f
C548 B.n491 VSUBS 0.007718f
C549 B.n492 VSUBS 0.007718f
C550 B.n493 VSUBS 0.007718f
C551 B.n494 VSUBS 0.007718f
C552 B.n495 VSUBS 0.007718f
C553 B.n496 VSUBS 0.007718f
C554 B.n497 VSUBS 0.007718f
C555 B.n498 VSUBS 0.007264f
C556 B.n499 VSUBS 0.007718f
C557 B.n500 VSUBS 0.007718f
C558 B.n501 VSUBS 0.007718f
C559 B.n502 VSUBS 0.007718f
C560 B.n503 VSUBS 0.007718f
C561 B.n504 VSUBS 0.007718f
C562 B.n505 VSUBS 0.007718f
C563 B.n506 VSUBS 0.007718f
C564 B.n507 VSUBS 0.007718f
C565 B.n508 VSUBS 0.007718f
C566 B.n509 VSUBS 0.007718f
C567 B.n510 VSUBS 0.007718f
C568 B.n511 VSUBS 0.007718f
C569 B.n512 VSUBS 0.007718f
C570 B.n513 VSUBS 0.007718f
C571 B.n514 VSUBS 0.004313f
C572 B.n515 VSUBS 0.017881f
C573 B.n516 VSUBS 0.007264f
C574 B.n517 VSUBS 0.007718f
C575 B.n518 VSUBS 0.007718f
C576 B.n519 VSUBS 0.007718f
C577 B.n520 VSUBS 0.007718f
C578 B.n521 VSUBS 0.007718f
C579 B.n522 VSUBS 0.007718f
C580 B.n523 VSUBS 0.007718f
C581 B.n524 VSUBS 0.007718f
C582 B.n525 VSUBS 0.007718f
C583 B.n526 VSUBS 0.007718f
C584 B.n527 VSUBS 0.007718f
C585 B.n528 VSUBS 0.007718f
C586 B.n529 VSUBS 0.007718f
C587 B.n530 VSUBS 0.007718f
C588 B.n531 VSUBS 0.007718f
C589 B.n532 VSUBS 0.007718f
C590 B.n533 VSUBS 0.007718f
C591 B.n534 VSUBS 0.007718f
C592 B.n535 VSUBS 0.007718f
C593 B.n536 VSUBS 0.007718f
C594 B.n537 VSUBS 0.007718f
C595 B.n538 VSUBS 0.007718f
C596 B.n539 VSUBS 0.007718f
C597 B.n540 VSUBS 0.007718f
C598 B.n541 VSUBS 0.007718f
C599 B.n542 VSUBS 0.007718f
C600 B.n543 VSUBS 0.007718f
C601 B.n544 VSUBS 0.007718f
C602 B.n545 VSUBS 0.007718f
C603 B.n546 VSUBS 0.007718f
C604 B.n547 VSUBS 0.007718f
C605 B.n548 VSUBS 0.007718f
C606 B.n549 VSUBS 0.007718f
C607 B.n550 VSUBS 0.007718f
C608 B.n551 VSUBS 0.007718f
C609 B.n552 VSUBS 0.007718f
C610 B.n553 VSUBS 0.007718f
C611 B.n554 VSUBS 0.007718f
C612 B.n555 VSUBS 0.007718f
C613 B.n556 VSUBS 0.007718f
C614 B.n557 VSUBS 0.007718f
C615 B.n558 VSUBS 0.007718f
C616 B.n559 VSUBS 0.007718f
C617 B.n560 VSUBS 0.007718f
C618 B.n561 VSUBS 0.007718f
C619 B.n562 VSUBS 0.007718f
C620 B.n563 VSUBS 0.007718f
C621 B.n564 VSUBS 0.007718f
C622 B.n565 VSUBS 0.007718f
C623 B.n566 VSUBS 0.007718f
C624 B.n567 VSUBS 0.007718f
C625 B.n568 VSUBS 0.007718f
C626 B.n569 VSUBS 0.007718f
C627 B.n570 VSUBS 0.007718f
C628 B.n571 VSUBS 0.007718f
C629 B.n572 VSUBS 0.007718f
C630 B.n573 VSUBS 0.007718f
C631 B.n574 VSUBS 0.007718f
C632 B.n575 VSUBS 0.007718f
C633 B.n576 VSUBS 0.007718f
C634 B.n577 VSUBS 0.007718f
C635 B.n578 VSUBS 0.007718f
C636 B.n579 VSUBS 0.007718f
C637 B.n580 VSUBS 0.007718f
C638 B.n581 VSUBS 0.007718f
C639 B.n582 VSUBS 0.007718f
C640 B.n583 VSUBS 0.007718f
C641 B.n584 VSUBS 0.007718f
C642 B.n585 VSUBS 0.007718f
C643 B.n586 VSUBS 0.007718f
C644 B.n587 VSUBS 0.007718f
C645 B.n588 VSUBS 0.007718f
C646 B.n589 VSUBS 0.007718f
C647 B.n590 VSUBS 0.007718f
C648 B.n591 VSUBS 0.007718f
C649 B.n592 VSUBS 0.007718f
C650 B.n593 VSUBS 0.007718f
C651 B.n594 VSUBS 0.019171f
C652 B.n595 VSUBS 0.018737f
C653 B.n596 VSUBS 0.018737f
C654 B.n597 VSUBS 0.007718f
C655 B.n598 VSUBS 0.007718f
C656 B.n599 VSUBS 0.007718f
C657 B.n600 VSUBS 0.007718f
C658 B.n601 VSUBS 0.007718f
C659 B.n602 VSUBS 0.007718f
C660 B.n603 VSUBS 0.007718f
C661 B.n604 VSUBS 0.007718f
C662 B.n605 VSUBS 0.007718f
C663 B.n606 VSUBS 0.007718f
C664 B.n607 VSUBS 0.007718f
C665 B.n608 VSUBS 0.007718f
C666 B.n609 VSUBS 0.007718f
C667 B.n610 VSUBS 0.007718f
C668 B.n611 VSUBS 0.007718f
C669 B.n612 VSUBS 0.007718f
C670 B.n613 VSUBS 0.007718f
C671 B.n614 VSUBS 0.007718f
C672 B.n615 VSUBS 0.007718f
C673 B.n616 VSUBS 0.007718f
C674 B.n617 VSUBS 0.007718f
C675 B.n618 VSUBS 0.007718f
C676 B.n619 VSUBS 0.007718f
C677 B.n620 VSUBS 0.007718f
C678 B.n621 VSUBS 0.007718f
C679 B.n622 VSUBS 0.007718f
C680 B.n623 VSUBS 0.017476f
C681 VTAIL.n0 VSUBS 0.02285f
C682 VTAIL.n1 VSUBS 0.022347f
C683 VTAIL.n2 VSUBS 0.012008f
C684 VTAIL.n3 VSUBS 0.028383f
C685 VTAIL.n4 VSUBS 0.012715f
C686 VTAIL.n5 VSUBS 0.022347f
C687 VTAIL.n6 VSUBS 0.012361f
C688 VTAIL.n7 VSUBS 0.028383f
C689 VTAIL.n8 VSUBS 0.012715f
C690 VTAIL.n9 VSUBS 0.022347f
C691 VTAIL.n10 VSUBS 0.012008f
C692 VTAIL.n11 VSUBS 0.028383f
C693 VTAIL.n12 VSUBS 0.012715f
C694 VTAIL.n13 VSUBS 0.022347f
C695 VTAIL.n14 VSUBS 0.012008f
C696 VTAIL.n15 VSUBS 0.028383f
C697 VTAIL.n16 VSUBS 0.012715f
C698 VTAIL.n17 VSUBS 0.022347f
C699 VTAIL.n18 VSUBS 0.012008f
C700 VTAIL.n19 VSUBS 0.028383f
C701 VTAIL.n20 VSUBS 0.012715f
C702 VTAIL.n21 VSUBS 0.022347f
C703 VTAIL.n22 VSUBS 0.012008f
C704 VTAIL.n23 VSUBS 0.028383f
C705 VTAIL.n24 VSUBS 0.012715f
C706 VTAIL.n25 VSUBS 0.022347f
C707 VTAIL.n26 VSUBS 0.012008f
C708 VTAIL.n27 VSUBS 0.021287f
C709 VTAIL.n28 VSUBS 0.018056f
C710 VTAIL.t4 VSUBS 0.060819f
C711 VTAIL.n29 VSUBS 0.164314f
C712 VTAIL.n30 VSUBS 1.53137f
C713 VTAIL.n31 VSUBS 0.012008f
C714 VTAIL.n32 VSUBS 0.012715f
C715 VTAIL.n33 VSUBS 0.028383f
C716 VTAIL.n34 VSUBS 0.028383f
C717 VTAIL.n35 VSUBS 0.012715f
C718 VTAIL.n36 VSUBS 0.012008f
C719 VTAIL.n37 VSUBS 0.022347f
C720 VTAIL.n38 VSUBS 0.022347f
C721 VTAIL.n39 VSUBS 0.012008f
C722 VTAIL.n40 VSUBS 0.012715f
C723 VTAIL.n41 VSUBS 0.028383f
C724 VTAIL.n42 VSUBS 0.028383f
C725 VTAIL.n43 VSUBS 0.012715f
C726 VTAIL.n44 VSUBS 0.012008f
C727 VTAIL.n45 VSUBS 0.022347f
C728 VTAIL.n46 VSUBS 0.022347f
C729 VTAIL.n47 VSUBS 0.012008f
C730 VTAIL.n48 VSUBS 0.012715f
C731 VTAIL.n49 VSUBS 0.028383f
C732 VTAIL.n50 VSUBS 0.028383f
C733 VTAIL.n51 VSUBS 0.012715f
C734 VTAIL.n52 VSUBS 0.012008f
C735 VTAIL.n53 VSUBS 0.022347f
C736 VTAIL.n54 VSUBS 0.022347f
C737 VTAIL.n55 VSUBS 0.012008f
C738 VTAIL.n56 VSUBS 0.012715f
C739 VTAIL.n57 VSUBS 0.028383f
C740 VTAIL.n58 VSUBS 0.028383f
C741 VTAIL.n59 VSUBS 0.012715f
C742 VTAIL.n60 VSUBS 0.012008f
C743 VTAIL.n61 VSUBS 0.022347f
C744 VTAIL.n62 VSUBS 0.022347f
C745 VTAIL.n63 VSUBS 0.012008f
C746 VTAIL.n64 VSUBS 0.012715f
C747 VTAIL.n65 VSUBS 0.028383f
C748 VTAIL.n66 VSUBS 0.028383f
C749 VTAIL.n67 VSUBS 0.012715f
C750 VTAIL.n68 VSUBS 0.012008f
C751 VTAIL.n69 VSUBS 0.022347f
C752 VTAIL.n70 VSUBS 0.022347f
C753 VTAIL.n71 VSUBS 0.012008f
C754 VTAIL.n72 VSUBS 0.012008f
C755 VTAIL.n73 VSUBS 0.012715f
C756 VTAIL.n74 VSUBS 0.028383f
C757 VTAIL.n75 VSUBS 0.028383f
C758 VTAIL.n76 VSUBS 0.028383f
C759 VTAIL.n77 VSUBS 0.012361f
C760 VTAIL.n78 VSUBS 0.012008f
C761 VTAIL.n79 VSUBS 0.022347f
C762 VTAIL.n80 VSUBS 0.022347f
C763 VTAIL.n81 VSUBS 0.012008f
C764 VTAIL.n82 VSUBS 0.012715f
C765 VTAIL.n83 VSUBS 0.028383f
C766 VTAIL.n84 VSUBS 0.062908f
C767 VTAIL.n85 VSUBS 0.012715f
C768 VTAIL.n86 VSUBS 0.012008f
C769 VTAIL.n87 VSUBS 0.050127f
C770 VTAIL.n88 VSUBS 0.031331f
C771 VTAIL.n89 VSUBS 0.091007f
C772 VTAIL.n90 VSUBS 0.02285f
C773 VTAIL.n91 VSUBS 0.022347f
C774 VTAIL.n92 VSUBS 0.012008f
C775 VTAIL.n93 VSUBS 0.028383f
C776 VTAIL.n94 VSUBS 0.012715f
C777 VTAIL.n95 VSUBS 0.022347f
C778 VTAIL.n96 VSUBS 0.012361f
C779 VTAIL.n97 VSUBS 0.028383f
C780 VTAIL.n98 VSUBS 0.012715f
C781 VTAIL.n99 VSUBS 0.022347f
C782 VTAIL.n100 VSUBS 0.012008f
C783 VTAIL.n101 VSUBS 0.028383f
C784 VTAIL.n102 VSUBS 0.012715f
C785 VTAIL.n103 VSUBS 0.022347f
C786 VTAIL.n104 VSUBS 0.012008f
C787 VTAIL.n105 VSUBS 0.028383f
C788 VTAIL.n106 VSUBS 0.012715f
C789 VTAIL.n107 VSUBS 0.022347f
C790 VTAIL.n108 VSUBS 0.012008f
C791 VTAIL.n109 VSUBS 0.028383f
C792 VTAIL.n110 VSUBS 0.012715f
C793 VTAIL.n111 VSUBS 0.022347f
C794 VTAIL.n112 VSUBS 0.012008f
C795 VTAIL.n113 VSUBS 0.028383f
C796 VTAIL.n114 VSUBS 0.012715f
C797 VTAIL.n115 VSUBS 0.022347f
C798 VTAIL.n116 VSUBS 0.012008f
C799 VTAIL.n117 VSUBS 0.021287f
C800 VTAIL.n118 VSUBS 0.018056f
C801 VTAIL.t3 VSUBS 0.060819f
C802 VTAIL.n119 VSUBS 0.164314f
C803 VTAIL.n120 VSUBS 1.53137f
C804 VTAIL.n121 VSUBS 0.012008f
C805 VTAIL.n122 VSUBS 0.012715f
C806 VTAIL.n123 VSUBS 0.028383f
C807 VTAIL.n124 VSUBS 0.028383f
C808 VTAIL.n125 VSUBS 0.012715f
C809 VTAIL.n126 VSUBS 0.012008f
C810 VTAIL.n127 VSUBS 0.022347f
C811 VTAIL.n128 VSUBS 0.022347f
C812 VTAIL.n129 VSUBS 0.012008f
C813 VTAIL.n130 VSUBS 0.012715f
C814 VTAIL.n131 VSUBS 0.028383f
C815 VTAIL.n132 VSUBS 0.028383f
C816 VTAIL.n133 VSUBS 0.012715f
C817 VTAIL.n134 VSUBS 0.012008f
C818 VTAIL.n135 VSUBS 0.022347f
C819 VTAIL.n136 VSUBS 0.022347f
C820 VTAIL.n137 VSUBS 0.012008f
C821 VTAIL.n138 VSUBS 0.012715f
C822 VTAIL.n139 VSUBS 0.028383f
C823 VTAIL.n140 VSUBS 0.028383f
C824 VTAIL.n141 VSUBS 0.012715f
C825 VTAIL.n142 VSUBS 0.012008f
C826 VTAIL.n143 VSUBS 0.022347f
C827 VTAIL.n144 VSUBS 0.022347f
C828 VTAIL.n145 VSUBS 0.012008f
C829 VTAIL.n146 VSUBS 0.012715f
C830 VTAIL.n147 VSUBS 0.028383f
C831 VTAIL.n148 VSUBS 0.028383f
C832 VTAIL.n149 VSUBS 0.012715f
C833 VTAIL.n150 VSUBS 0.012008f
C834 VTAIL.n151 VSUBS 0.022347f
C835 VTAIL.n152 VSUBS 0.022347f
C836 VTAIL.n153 VSUBS 0.012008f
C837 VTAIL.n154 VSUBS 0.012715f
C838 VTAIL.n155 VSUBS 0.028383f
C839 VTAIL.n156 VSUBS 0.028383f
C840 VTAIL.n157 VSUBS 0.012715f
C841 VTAIL.n158 VSUBS 0.012008f
C842 VTAIL.n159 VSUBS 0.022347f
C843 VTAIL.n160 VSUBS 0.022347f
C844 VTAIL.n161 VSUBS 0.012008f
C845 VTAIL.n162 VSUBS 0.012008f
C846 VTAIL.n163 VSUBS 0.012715f
C847 VTAIL.n164 VSUBS 0.028383f
C848 VTAIL.n165 VSUBS 0.028383f
C849 VTAIL.n166 VSUBS 0.028383f
C850 VTAIL.n167 VSUBS 0.012361f
C851 VTAIL.n168 VSUBS 0.012008f
C852 VTAIL.n169 VSUBS 0.022347f
C853 VTAIL.n170 VSUBS 0.022347f
C854 VTAIL.n171 VSUBS 0.012008f
C855 VTAIL.n172 VSUBS 0.012715f
C856 VTAIL.n173 VSUBS 0.028383f
C857 VTAIL.n174 VSUBS 0.062908f
C858 VTAIL.n175 VSUBS 0.012715f
C859 VTAIL.n176 VSUBS 0.012008f
C860 VTAIL.n177 VSUBS 0.050127f
C861 VTAIL.n178 VSUBS 0.031331f
C862 VTAIL.n179 VSUBS 0.121578f
C863 VTAIL.n180 VSUBS 0.02285f
C864 VTAIL.n181 VSUBS 0.022347f
C865 VTAIL.n182 VSUBS 0.012008f
C866 VTAIL.n183 VSUBS 0.028383f
C867 VTAIL.n184 VSUBS 0.012715f
C868 VTAIL.n185 VSUBS 0.022347f
C869 VTAIL.n186 VSUBS 0.012361f
C870 VTAIL.n187 VSUBS 0.028383f
C871 VTAIL.n188 VSUBS 0.012715f
C872 VTAIL.n189 VSUBS 0.022347f
C873 VTAIL.n190 VSUBS 0.012008f
C874 VTAIL.n191 VSUBS 0.028383f
C875 VTAIL.n192 VSUBS 0.012715f
C876 VTAIL.n193 VSUBS 0.022347f
C877 VTAIL.n194 VSUBS 0.012008f
C878 VTAIL.n195 VSUBS 0.028383f
C879 VTAIL.n196 VSUBS 0.012715f
C880 VTAIL.n197 VSUBS 0.022347f
C881 VTAIL.n198 VSUBS 0.012008f
C882 VTAIL.n199 VSUBS 0.028383f
C883 VTAIL.n200 VSUBS 0.012715f
C884 VTAIL.n201 VSUBS 0.022347f
C885 VTAIL.n202 VSUBS 0.012008f
C886 VTAIL.n203 VSUBS 0.028383f
C887 VTAIL.n204 VSUBS 0.012715f
C888 VTAIL.n205 VSUBS 0.022347f
C889 VTAIL.n206 VSUBS 0.012008f
C890 VTAIL.n207 VSUBS 0.021287f
C891 VTAIL.n208 VSUBS 0.018056f
C892 VTAIL.t0 VSUBS 0.060819f
C893 VTAIL.n209 VSUBS 0.164314f
C894 VTAIL.n210 VSUBS 1.53137f
C895 VTAIL.n211 VSUBS 0.012008f
C896 VTAIL.n212 VSUBS 0.012715f
C897 VTAIL.n213 VSUBS 0.028383f
C898 VTAIL.n214 VSUBS 0.028383f
C899 VTAIL.n215 VSUBS 0.012715f
C900 VTAIL.n216 VSUBS 0.012008f
C901 VTAIL.n217 VSUBS 0.022347f
C902 VTAIL.n218 VSUBS 0.022347f
C903 VTAIL.n219 VSUBS 0.012008f
C904 VTAIL.n220 VSUBS 0.012715f
C905 VTAIL.n221 VSUBS 0.028383f
C906 VTAIL.n222 VSUBS 0.028383f
C907 VTAIL.n223 VSUBS 0.012715f
C908 VTAIL.n224 VSUBS 0.012008f
C909 VTAIL.n225 VSUBS 0.022347f
C910 VTAIL.n226 VSUBS 0.022347f
C911 VTAIL.n227 VSUBS 0.012008f
C912 VTAIL.n228 VSUBS 0.012715f
C913 VTAIL.n229 VSUBS 0.028383f
C914 VTAIL.n230 VSUBS 0.028383f
C915 VTAIL.n231 VSUBS 0.012715f
C916 VTAIL.n232 VSUBS 0.012008f
C917 VTAIL.n233 VSUBS 0.022347f
C918 VTAIL.n234 VSUBS 0.022347f
C919 VTAIL.n235 VSUBS 0.012008f
C920 VTAIL.n236 VSUBS 0.012715f
C921 VTAIL.n237 VSUBS 0.028383f
C922 VTAIL.n238 VSUBS 0.028383f
C923 VTAIL.n239 VSUBS 0.012715f
C924 VTAIL.n240 VSUBS 0.012008f
C925 VTAIL.n241 VSUBS 0.022347f
C926 VTAIL.n242 VSUBS 0.022347f
C927 VTAIL.n243 VSUBS 0.012008f
C928 VTAIL.n244 VSUBS 0.012715f
C929 VTAIL.n245 VSUBS 0.028383f
C930 VTAIL.n246 VSUBS 0.028383f
C931 VTAIL.n247 VSUBS 0.012715f
C932 VTAIL.n248 VSUBS 0.012008f
C933 VTAIL.n249 VSUBS 0.022347f
C934 VTAIL.n250 VSUBS 0.022347f
C935 VTAIL.n251 VSUBS 0.012008f
C936 VTAIL.n252 VSUBS 0.012008f
C937 VTAIL.n253 VSUBS 0.012715f
C938 VTAIL.n254 VSUBS 0.028383f
C939 VTAIL.n255 VSUBS 0.028383f
C940 VTAIL.n256 VSUBS 0.028383f
C941 VTAIL.n257 VSUBS 0.012361f
C942 VTAIL.n258 VSUBS 0.012008f
C943 VTAIL.n259 VSUBS 0.022347f
C944 VTAIL.n260 VSUBS 0.022347f
C945 VTAIL.n261 VSUBS 0.012008f
C946 VTAIL.n262 VSUBS 0.012715f
C947 VTAIL.n263 VSUBS 0.028383f
C948 VTAIL.n264 VSUBS 0.062908f
C949 VTAIL.n265 VSUBS 0.012715f
C950 VTAIL.n266 VSUBS 0.012008f
C951 VTAIL.n267 VSUBS 0.050127f
C952 VTAIL.n268 VSUBS 0.031331f
C953 VTAIL.n269 VSUBS 1.45587f
C954 VTAIL.n270 VSUBS 0.02285f
C955 VTAIL.n271 VSUBS 0.022347f
C956 VTAIL.n272 VSUBS 0.012008f
C957 VTAIL.n273 VSUBS 0.028383f
C958 VTAIL.n274 VSUBS 0.012715f
C959 VTAIL.n275 VSUBS 0.022347f
C960 VTAIL.n276 VSUBS 0.012361f
C961 VTAIL.n277 VSUBS 0.028383f
C962 VTAIL.n278 VSUBS 0.012008f
C963 VTAIL.n279 VSUBS 0.012715f
C964 VTAIL.n280 VSUBS 0.022347f
C965 VTAIL.n281 VSUBS 0.012008f
C966 VTAIL.n282 VSUBS 0.028383f
C967 VTAIL.n283 VSUBS 0.012715f
C968 VTAIL.n284 VSUBS 0.022347f
C969 VTAIL.n285 VSUBS 0.012008f
C970 VTAIL.n286 VSUBS 0.028383f
C971 VTAIL.n287 VSUBS 0.012715f
C972 VTAIL.n288 VSUBS 0.022347f
C973 VTAIL.n289 VSUBS 0.012008f
C974 VTAIL.n290 VSUBS 0.028383f
C975 VTAIL.n291 VSUBS 0.012715f
C976 VTAIL.n292 VSUBS 0.022347f
C977 VTAIL.n293 VSUBS 0.012008f
C978 VTAIL.n294 VSUBS 0.028383f
C979 VTAIL.n295 VSUBS 0.012715f
C980 VTAIL.n296 VSUBS 0.022347f
C981 VTAIL.n297 VSUBS 0.012008f
C982 VTAIL.n298 VSUBS 0.021287f
C983 VTAIL.n299 VSUBS 0.018056f
C984 VTAIL.t7 VSUBS 0.060819f
C985 VTAIL.n300 VSUBS 0.164314f
C986 VTAIL.n301 VSUBS 1.53137f
C987 VTAIL.n302 VSUBS 0.012008f
C988 VTAIL.n303 VSUBS 0.012715f
C989 VTAIL.n304 VSUBS 0.028383f
C990 VTAIL.n305 VSUBS 0.028383f
C991 VTAIL.n306 VSUBS 0.012715f
C992 VTAIL.n307 VSUBS 0.012008f
C993 VTAIL.n308 VSUBS 0.022347f
C994 VTAIL.n309 VSUBS 0.022347f
C995 VTAIL.n310 VSUBS 0.012008f
C996 VTAIL.n311 VSUBS 0.012715f
C997 VTAIL.n312 VSUBS 0.028383f
C998 VTAIL.n313 VSUBS 0.028383f
C999 VTAIL.n314 VSUBS 0.012715f
C1000 VTAIL.n315 VSUBS 0.012008f
C1001 VTAIL.n316 VSUBS 0.022347f
C1002 VTAIL.n317 VSUBS 0.022347f
C1003 VTAIL.n318 VSUBS 0.012008f
C1004 VTAIL.n319 VSUBS 0.012715f
C1005 VTAIL.n320 VSUBS 0.028383f
C1006 VTAIL.n321 VSUBS 0.028383f
C1007 VTAIL.n322 VSUBS 0.012715f
C1008 VTAIL.n323 VSUBS 0.012008f
C1009 VTAIL.n324 VSUBS 0.022347f
C1010 VTAIL.n325 VSUBS 0.022347f
C1011 VTAIL.n326 VSUBS 0.012008f
C1012 VTAIL.n327 VSUBS 0.012715f
C1013 VTAIL.n328 VSUBS 0.028383f
C1014 VTAIL.n329 VSUBS 0.028383f
C1015 VTAIL.n330 VSUBS 0.012715f
C1016 VTAIL.n331 VSUBS 0.012008f
C1017 VTAIL.n332 VSUBS 0.022347f
C1018 VTAIL.n333 VSUBS 0.022347f
C1019 VTAIL.n334 VSUBS 0.012008f
C1020 VTAIL.n335 VSUBS 0.012715f
C1021 VTAIL.n336 VSUBS 0.028383f
C1022 VTAIL.n337 VSUBS 0.028383f
C1023 VTAIL.n338 VSUBS 0.012715f
C1024 VTAIL.n339 VSUBS 0.012008f
C1025 VTAIL.n340 VSUBS 0.022347f
C1026 VTAIL.n341 VSUBS 0.022347f
C1027 VTAIL.n342 VSUBS 0.012008f
C1028 VTAIL.n343 VSUBS 0.012715f
C1029 VTAIL.n344 VSUBS 0.028383f
C1030 VTAIL.n345 VSUBS 0.028383f
C1031 VTAIL.n346 VSUBS 0.028383f
C1032 VTAIL.n347 VSUBS 0.012361f
C1033 VTAIL.n348 VSUBS 0.012008f
C1034 VTAIL.n349 VSUBS 0.022347f
C1035 VTAIL.n350 VSUBS 0.022347f
C1036 VTAIL.n351 VSUBS 0.012008f
C1037 VTAIL.n352 VSUBS 0.012715f
C1038 VTAIL.n353 VSUBS 0.028383f
C1039 VTAIL.n354 VSUBS 0.062908f
C1040 VTAIL.n355 VSUBS 0.012715f
C1041 VTAIL.n356 VSUBS 0.012008f
C1042 VTAIL.n357 VSUBS 0.050127f
C1043 VTAIL.n358 VSUBS 0.031331f
C1044 VTAIL.n359 VSUBS 1.45587f
C1045 VTAIL.n360 VSUBS 0.02285f
C1046 VTAIL.n361 VSUBS 0.022347f
C1047 VTAIL.n362 VSUBS 0.012008f
C1048 VTAIL.n363 VSUBS 0.028383f
C1049 VTAIL.n364 VSUBS 0.012715f
C1050 VTAIL.n365 VSUBS 0.022347f
C1051 VTAIL.n366 VSUBS 0.012361f
C1052 VTAIL.n367 VSUBS 0.028383f
C1053 VTAIL.n368 VSUBS 0.012008f
C1054 VTAIL.n369 VSUBS 0.012715f
C1055 VTAIL.n370 VSUBS 0.022347f
C1056 VTAIL.n371 VSUBS 0.012008f
C1057 VTAIL.n372 VSUBS 0.028383f
C1058 VTAIL.n373 VSUBS 0.012715f
C1059 VTAIL.n374 VSUBS 0.022347f
C1060 VTAIL.n375 VSUBS 0.012008f
C1061 VTAIL.n376 VSUBS 0.028383f
C1062 VTAIL.n377 VSUBS 0.012715f
C1063 VTAIL.n378 VSUBS 0.022347f
C1064 VTAIL.n379 VSUBS 0.012008f
C1065 VTAIL.n380 VSUBS 0.028383f
C1066 VTAIL.n381 VSUBS 0.012715f
C1067 VTAIL.n382 VSUBS 0.022347f
C1068 VTAIL.n383 VSUBS 0.012008f
C1069 VTAIL.n384 VSUBS 0.028383f
C1070 VTAIL.n385 VSUBS 0.012715f
C1071 VTAIL.n386 VSUBS 0.022347f
C1072 VTAIL.n387 VSUBS 0.012008f
C1073 VTAIL.n388 VSUBS 0.021287f
C1074 VTAIL.n389 VSUBS 0.018056f
C1075 VTAIL.t5 VSUBS 0.060819f
C1076 VTAIL.n390 VSUBS 0.164314f
C1077 VTAIL.n391 VSUBS 1.53137f
C1078 VTAIL.n392 VSUBS 0.012008f
C1079 VTAIL.n393 VSUBS 0.012715f
C1080 VTAIL.n394 VSUBS 0.028383f
C1081 VTAIL.n395 VSUBS 0.028383f
C1082 VTAIL.n396 VSUBS 0.012715f
C1083 VTAIL.n397 VSUBS 0.012008f
C1084 VTAIL.n398 VSUBS 0.022347f
C1085 VTAIL.n399 VSUBS 0.022347f
C1086 VTAIL.n400 VSUBS 0.012008f
C1087 VTAIL.n401 VSUBS 0.012715f
C1088 VTAIL.n402 VSUBS 0.028383f
C1089 VTAIL.n403 VSUBS 0.028383f
C1090 VTAIL.n404 VSUBS 0.012715f
C1091 VTAIL.n405 VSUBS 0.012008f
C1092 VTAIL.n406 VSUBS 0.022347f
C1093 VTAIL.n407 VSUBS 0.022347f
C1094 VTAIL.n408 VSUBS 0.012008f
C1095 VTAIL.n409 VSUBS 0.012715f
C1096 VTAIL.n410 VSUBS 0.028383f
C1097 VTAIL.n411 VSUBS 0.028383f
C1098 VTAIL.n412 VSUBS 0.012715f
C1099 VTAIL.n413 VSUBS 0.012008f
C1100 VTAIL.n414 VSUBS 0.022347f
C1101 VTAIL.n415 VSUBS 0.022347f
C1102 VTAIL.n416 VSUBS 0.012008f
C1103 VTAIL.n417 VSUBS 0.012715f
C1104 VTAIL.n418 VSUBS 0.028383f
C1105 VTAIL.n419 VSUBS 0.028383f
C1106 VTAIL.n420 VSUBS 0.012715f
C1107 VTAIL.n421 VSUBS 0.012008f
C1108 VTAIL.n422 VSUBS 0.022347f
C1109 VTAIL.n423 VSUBS 0.022347f
C1110 VTAIL.n424 VSUBS 0.012008f
C1111 VTAIL.n425 VSUBS 0.012715f
C1112 VTAIL.n426 VSUBS 0.028383f
C1113 VTAIL.n427 VSUBS 0.028383f
C1114 VTAIL.n428 VSUBS 0.012715f
C1115 VTAIL.n429 VSUBS 0.012008f
C1116 VTAIL.n430 VSUBS 0.022347f
C1117 VTAIL.n431 VSUBS 0.022347f
C1118 VTAIL.n432 VSUBS 0.012008f
C1119 VTAIL.n433 VSUBS 0.012715f
C1120 VTAIL.n434 VSUBS 0.028383f
C1121 VTAIL.n435 VSUBS 0.028383f
C1122 VTAIL.n436 VSUBS 0.028383f
C1123 VTAIL.n437 VSUBS 0.012361f
C1124 VTAIL.n438 VSUBS 0.012008f
C1125 VTAIL.n439 VSUBS 0.022347f
C1126 VTAIL.n440 VSUBS 0.022347f
C1127 VTAIL.n441 VSUBS 0.012008f
C1128 VTAIL.n442 VSUBS 0.012715f
C1129 VTAIL.n443 VSUBS 0.028383f
C1130 VTAIL.n444 VSUBS 0.062908f
C1131 VTAIL.n445 VSUBS 0.012715f
C1132 VTAIL.n446 VSUBS 0.012008f
C1133 VTAIL.n447 VSUBS 0.050127f
C1134 VTAIL.n448 VSUBS 0.031331f
C1135 VTAIL.n449 VSUBS 0.121578f
C1136 VTAIL.n450 VSUBS 0.02285f
C1137 VTAIL.n451 VSUBS 0.022347f
C1138 VTAIL.n452 VSUBS 0.012008f
C1139 VTAIL.n453 VSUBS 0.028383f
C1140 VTAIL.n454 VSUBS 0.012715f
C1141 VTAIL.n455 VSUBS 0.022347f
C1142 VTAIL.n456 VSUBS 0.012361f
C1143 VTAIL.n457 VSUBS 0.028383f
C1144 VTAIL.n458 VSUBS 0.012008f
C1145 VTAIL.n459 VSUBS 0.012715f
C1146 VTAIL.n460 VSUBS 0.022347f
C1147 VTAIL.n461 VSUBS 0.012008f
C1148 VTAIL.n462 VSUBS 0.028383f
C1149 VTAIL.n463 VSUBS 0.012715f
C1150 VTAIL.n464 VSUBS 0.022347f
C1151 VTAIL.n465 VSUBS 0.012008f
C1152 VTAIL.n466 VSUBS 0.028383f
C1153 VTAIL.n467 VSUBS 0.012715f
C1154 VTAIL.n468 VSUBS 0.022347f
C1155 VTAIL.n469 VSUBS 0.012008f
C1156 VTAIL.n470 VSUBS 0.028383f
C1157 VTAIL.n471 VSUBS 0.012715f
C1158 VTAIL.n472 VSUBS 0.022347f
C1159 VTAIL.n473 VSUBS 0.012008f
C1160 VTAIL.n474 VSUBS 0.028383f
C1161 VTAIL.n475 VSUBS 0.012715f
C1162 VTAIL.n476 VSUBS 0.022347f
C1163 VTAIL.n477 VSUBS 0.012008f
C1164 VTAIL.n478 VSUBS 0.021287f
C1165 VTAIL.n479 VSUBS 0.018056f
C1166 VTAIL.t2 VSUBS 0.060819f
C1167 VTAIL.n480 VSUBS 0.164314f
C1168 VTAIL.n481 VSUBS 1.53137f
C1169 VTAIL.n482 VSUBS 0.012008f
C1170 VTAIL.n483 VSUBS 0.012715f
C1171 VTAIL.n484 VSUBS 0.028383f
C1172 VTAIL.n485 VSUBS 0.028383f
C1173 VTAIL.n486 VSUBS 0.012715f
C1174 VTAIL.n487 VSUBS 0.012008f
C1175 VTAIL.n488 VSUBS 0.022347f
C1176 VTAIL.n489 VSUBS 0.022347f
C1177 VTAIL.n490 VSUBS 0.012008f
C1178 VTAIL.n491 VSUBS 0.012715f
C1179 VTAIL.n492 VSUBS 0.028383f
C1180 VTAIL.n493 VSUBS 0.028383f
C1181 VTAIL.n494 VSUBS 0.012715f
C1182 VTAIL.n495 VSUBS 0.012008f
C1183 VTAIL.n496 VSUBS 0.022347f
C1184 VTAIL.n497 VSUBS 0.022347f
C1185 VTAIL.n498 VSUBS 0.012008f
C1186 VTAIL.n499 VSUBS 0.012715f
C1187 VTAIL.n500 VSUBS 0.028383f
C1188 VTAIL.n501 VSUBS 0.028383f
C1189 VTAIL.n502 VSUBS 0.012715f
C1190 VTAIL.n503 VSUBS 0.012008f
C1191 VTAIL.n504 VSUBS 0.022347f
C1192 VTAIL.n505 VSUBS 0.022347f
C1193 VTAIL.n506 VSUBS 0.012008f
C1194 VTAIL.n507 VSUBS 0.012715f
C1195 VTAIL.n508 VSUBS 0.028383f
C1196 VTAIL.n509 VSUBS 0.028383f
C1197 VTAIL.n510 VSUBS 0.012715f
C1198 VTAIL.n511 VSUBS 0.012008f
C1199 VTAIL.n512 VSUBS 0.022347f
C1200 VTAIL.n513 VSUBS 0.022347f
C1201 VTAIL.n514 VSUBS 0.012008f
C1202 VTAIL.n515 VSUBS 0.012715f
C1203 VTAIL.n516 VSUBS 0.028383f
C1204 VTAIL.n517 VSUBS 0.028383f
C1205 VTAIL.n518 VSUBS 0.012715f
C1206 VTAIL.n519 VSUBS 0.012008f
C1207 VTAIL.n520 VSUBS 0.022347f
C1208 VTAIL.n521 VSUBS 0.022347f
C1209 VTAIL.n522 VSUBS 0.012008f
C1210 VTAIL.n523 VSUBS 0.012715f
C1211 VTAIL.n524 VSUBS 0.028383f
C1212 VTAIL.n525 VSUBS 0.028383f
C1213 VTAIL.n526 VSUBS 0.028383f
C1214 VTAIL.n527 VSUBS 0.012361f
C1215 VTAIL.n528 VSUBS 0.012008f
C1216 VTAIL.n529 VSUBS 0.022347f
C1217 VTAIL.n530 VSUBS 0.022347f
C1218 VTAIL.n531 VSUBS 0.012008f
C1219 VTAIL.n532 VSUBS 0.012715f
C1220 VTAIL.n533 VSUBS 0.028383f
C1221 VTAIL.n534 VSUBS 0.062908f
C1222 VTAIL.n535 VSUBS 0.012715f
C1223 VTAIL.n536 VSUBS 0.012008f
C1224 VTAIL.n537 VSUBS 0.050127f
C1225 VTAIL.n538 VSUBS 0.031331f
C1226 VTAIL.n539 VSUBS 0.121578f
C1227 VTAIL.n540 VSUBS 0.02285f
C1228 VTAIL.n541 VSUBS 0.022347f
C1229 VTAIL.n542 VSUBS 0.012008f
C1230 VTAIL.n543 VSUBS 0.028383f
C1231 VTAIL.n544 VSUBS 0.012715f
C1232 VTAIL.n545 VSUBS 0.022347f
C1233 VTAIL.n546 VSUBS 0.012361f
C1234 VTAIL.n547 VSUBS 0.028383f
C1235 VTAIL.n548 VSUBS 0.012008f
C1236 VTAIL.n549 VSUBS 0.012715f
C1237 VTAIL.n550 VSUBS 0.022347f
C1238 VTAIL.n551 VSUBS 0.012008f
C1239 VTAIL.n552 VSUBS 0.028383f
C1240 VTAIL.n553 VSUBS 0.012715f
C1241 VTAIL.n554 VSUBS 0.022347f
C1242 VTAIL.n555 VSUBS 0.012008f
C1243 VTAIL.n556 VSUBS 0.028383f
C1244 VTAIL.n557 VSUBS 0.012715f
C1245 VTAIL.n558 VSUBS 0.022347f
C1246 VTAIL.n559 VSUBS 0.012008f
C1247 VTAIL.n560 VSUBS 0.028383f
C1248 VTAIL.n561 VSUBS 0.012715f
C1249 VTAIL.n562 VSUBS 0.022347f
C1250 VTAIL.n563 VSUBS 0.012008f
C1251 VTAIL.n564 VSUBS 0.028383f
C1252 VTAIL.n565 VSUBS 0.012715f
C1253 VTAIL.n566 VSUBS 0.022347f
C1254 VTAIL.n567 VSUBS 0.012008f
C1255 VTAIL.n568 VSUBS 0.021287f
C1256 VTAIL.n569 VSUBS 0.018056f
C1257 VTAIL.t1 VSUBS 0.060819f
C1258 VTAIL.n570 VSUBS 0.164314f
C1259 VTAIL.n571 VSUBS 1.53137f
C1260 VTAIL.n572 VSUBS 0.012008f
C1261 VTAIL.n573 VSUBS 0.012715f
C1262 VTAIL.n574 VSUBS 0.028383f
C1263 VTAIL.n575 VSUBS 0.028383f
C1264 VTAIL.n576 VSUBS 0.012715f
C1265 VTAIL.n577 VSUBS 0.012008f
C1266 VTAIL.n578 VSUBS 0.022347f
C1267 VTAIL.n579 VSUBS 0.022347f
C1268 VTAIL.n580 VSUBS 0.012008f
C1269 VTAIL.n581 VSUBS 0.012715f
C1270 VTAIL.n582 VSUBS 0.028383f
C1271 VTAIL.n583 VSUBS 0.028383f
C1272 VTAIL.n584 VSUBS 0.012715f
C1273 VTAIL.n585 VSUBS 0.012008f
C1274 VTAIL.n586 VSUBS 0.022347f
C1275 VTAIL.n587 VSUBS 0.022347f
C1276 VTAIL.n588 VSUBS 0.012008f
C1277 VTAIL.n589 VSUBS 0.012715f
C1278 VTAIL.n590 VSUBS 0.028383f
C1279 VTAIL.n591 VSUBS 0.028383f
C1280 VTAIL.n592 VSUBS 0.012715f
C1281 VTAIL.n593 VSUBS 0.012008f
C1282 VTAIL.n594 VSUBS 0.022347f
C1283 VTAIL.n595 VSUBS 0.022347f
C1284 VTAIL.n596 VSUBS 0.012008f
C1285 VTAIL.n597 VSUBS 0.012715f
C1286 VTAIL.n598 VSUBS 0.028383f
C1287 VTAIL.n599 VSUBS 0.028383f
C1288 VTAIL.n600 VSUBS 0.012715f
C1289 VTAIL.n601 VSUBS 0.012008f
C1290 VTAIL.n602 VSUBS 0.022347f
C1291 VTAIL.n603 VSUBS 0.022347f
C1292 VTAIL.n604 VSUBS 0.012008f
C1293 VTAIL.n605 VSUBS 0.012715f
C1294 VTAIL.n606 VSUBS 0.028383f
C1295 VTAIL.n607 VSUBS 0.028383f
C1296 VTAIL.n608 VSUBS 0.012715f
C1297 VTAIL.n609 VSUBS 0.012008f
C1298 VTAIL.n610 VSUBS 0.022347f
C1299 VTAIL.n611 VSUBS 0.022347f
C1300 VTAIL.n612 VSUBS 0.012008f
C1301 VTAIL.n613 VSUBS 0.012715f
C1302 VTAIL.n614 VSUBS 0.028383f
C1303 VTAIL.n615 VSUBS 0.028383f
C1304 VTAIL.n616 VSUBS 0.028383f
C1305 VTAIL.n617 VSUBS 0.012361f
C1306 VTAIL.n618 VSUBS 0.012008f
C1307 VTAIL.n619 VSUBS 0.022347f
C1308 VTAIL.n620 VSUBS 0.022347f
C1309 VTAIL.n621 VSUBS 0.012008f
C1310 VTAIL.n622 VSUBS 0.012715f
C1311 VTAIL.n623 VSUBS 0.028383f
C1312 VTAIL.n624 VSUBS 0.062908f
C1313 VTAIL.n625 VSUBS 0.012715f
C1314 VTAIL.n626 VSUBS 0.012008f
C1315 VTAIL.n627 VSUBS 0.050127f
C1316 VTAIL.n628 VSUBS 0.031331f
C1317 VTAIL.n629 VSUBS 1.45587f
C1318 VTAIL.n630 VSUBS 0.02285f
C1319 VTAIL.n631 VSUBS 0.022347f
C1320 VTAIL.n632 VSUBS 0.012008f
C1321 VTAIL.n633 VSUBS 0.028383f
C1322 VTAIL.n634 VSUBS 0.012715f
C1323 VTAIL.n635 VSUBS 0.022347f
C1324 VTAIL.n636 VSUBS 0.012361f
C1325 VTAIL.n637 VSUBS 0.028383f
C1326 VTAIL.n638 VSUBS 0.012715f
C1327 VTAIL.n639 VSUBS 0.022347f
C1328 VTAIL.n640 VSUBS 0.012008f
C1329 VTAIL.n641 VSUBS 0.028383f
C1330 VTAIL.n642 VSUBS 0.012715f
C1331 VTAIL.n643 VSUBS 0.022347f
C1332 VTAIL.n644 VSUBS 0.012008f
C1333 VTAIL.n645 VSUBS 0.028383f
C1334 VTAIL.n646 VSUBS 0.012715f
C1335 VTAIL.n647 VSUBS 0.022347f
C1336 VTAIL.n648 VSUBS 0.012008f
C1337 VTAIL.n649 VSUBS 0.028383f
C1338 VTAIL.n650 VSUBS 0.012715f
C1339 VTAIL.n651 VSUBS 0.022347f
C1340 VTAIL.n652 VSUBS 0.012008f
C1341 VTAIL.n653 VSUBS 0.028383f
C1342 VTAIL.n654 VSUBS 0.012715f
C1343 VTAIL.n655 VSUBS 0.022347f
C1344 VTAIL.n656 VSUBS 0.012008f
C1345 VTAIL.n657 VSUBS 0.021287f
C1346 VTAIL.n658 VSUBS 0.018056f
C1347 VTAIL.t6 VSUBS 0.060819f
C1348 VTAIL.n659 VSUBS 0.164314f
C1349 VTAIL.n660 VSUBS 1.53137f
C1350 VTAIL.n661 VSUBS 0.012008f
C1351 VTAIL.n662 VSUBS 0.012715f
C1352 VTAIL.n663 VSUBS 0.028383f
C1353 VTAIL.n664 VSUBS 0.028383f
C1354 VTAIL.n665 VSUBS 0.012715f
C1355 VTAIL.n666 VSUBS 0.012008f
C1356 VTAIL.n667 VSUBS 0.022347f
C1357 VTAIL.n668 VSUBS 0.022347f
C1358 VTAIL.n669 VSUBS 0.012008f
C1359 VTAIL.n670 VSUBS 0.012715f
C1360 VTAIL.n671 VSUBS 0.028383f
C1361 VTAIL.n672 VSUBS 0.028383f
C1362 VTAIL.n673 VSUBS 0.012715f
C1363 VTAIL.n674 VSUBS 0.012008f
C1364 VTAIL.n675 VSUBS 0.022347f
C1365 VTAIL.n676 VSUBS 0.022347f
C1366 VTAIL.n677 VSUBS 0.012008f
C1367 VTAIL.n678 VSUBS 0.012715f
C1368 VTAIL.n679 VSUBS 0.028383f
C1369 VTAIL.n680 VSUBS 0.028383f
C1370 VTAIL.n681 VSUBS 0.012715f
C1371 VTAIL.n682 VSUBS 0.012008f
C1372 VTAIL.n683 VSUBS 0.022347f
C1373 VTAIL.n684 VSUBS 0.022347f
C1374 VTAIL.n685 VSUBS 0.012008f
C1375 VTAIL.n686 VSUBS 0.012715f
C1376 VTAIL.n687 VSUBS 0.028383f
C1377 VTAIL.n688 VSUBS 0.028383f
C1378 VTAIL.n689 VSUBS 0.012715f
C1379 VTAIL.n690 VSUBS 0.012008f
C1380 VTAIL.n691 VSUBS 0.022347f
C1381 VTAIL.n692 VSUBS 0.022347f
C1382 VTAIL.n693 VSUBS 0.012008f
C1383 VTAIL.n694 VSUBS 0.012715f
C1384 VTAIL.n695 VSUBS 0.028383f
C1385 VTAIL.n696 VSUBS 0.028383f
C1386 VTAIL.n697 VSUBS 0.012715f
C1387 VTAIL.n698 VSUBS 0.012008f
C1388 VTAIL.n699 VSUBS 0.022347f
C1389 VTAIL.n700 VSUBS 0.022347f
C1390 VTAIL.n701 VSUBS 0.012008f
C1391 VTAIL.n702 VSUBS 0.012008f
C1392 VTAIL.n703 VSUBS 0.012715f
C1393 VTAIL.n704 VSUBS 0.028383f
C1394 VTAIL.n705 VSUBS 0.028383f
C1395 VTAIL.n706 VSUBS 0.028383f
C1396 VTAIL.n707 VSUBS 0.012361f
C1397 VTAIL.n708 VSUBS 0.012008f
C1398 VTAIL.n709 VSUBS 0.022347f
C1399 VTAIL.n710 VSUBS 0.022347f
C1400 VTAIL.n711 VSUBS 0.012008f
C1401 VTAIL.n712 VSUBS 0.012715f
C1402 VTAIL.n713 VSUBS 0.028383f
C1403 VTAIL.n714 VSUBS 0.062908f
C1404 VTAIL.n715 VSUBS 0.012715f
C1405 VTAIL.n716 VSUBS 0.012008f
C1406 VTAIL.n717 VSUBS 0.050127f
C1407 VTAIL.n718 VSUBS 0.031331f
C1408 VTAIL.n719 VSUBS 1.41692f
C1409 VDD2.t3 VSUBS 0.353829f
C1410 VDD2.t1 VSUBS 0.353829f
C1411 VDD2.n0 VSUBS 3.71017f
C1412 VDD2.t2 VSUBS 0.353829f
C1413 VDD2.t0 VSUBS 0.353829f
C1414 VDD2.n1 VSUBS 2.89119f
C1415 VDD2.n2 VSUBS 4.49041f
C1416 VN.t3 VSUBS 2.02163f
C1417 VN.t1 VSUBS 2.02156f
C1418 VN.n0 VSUBS 1.46949f
C1419 VN.t2 VSUBS 2.02163f
C1420 VN.t0 VSUBS 2.02156f
C1421 VN.n1 VSUBS 2.76833f
.ends

