* NGSPICE file created from diff_pair_sample_0069.ext - technology: sky130A

.subckt diff_pair_sample_0069 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t9 w_n2594_n1740# sky130_fd_pr__pfet_01v8 ad=0.6369 pd=4.19 as=1.5054 ps=8.5 w=3.86 l=1.7
X1 VTAIL.t3 VN.t0 VDD2.t5 w_n2594_n1740# sky130_fd_pr__pfet_01v8 ad=0.6369 pd=4.19 as=0.6369 ps=4.19 w=3.86 l=1.7
X2 VDD2.t4 VN.t1 VTAIL.t0 w_n2594_n1740# sky130_fd_pr__pfet_01v8 ad=1.5054 pd=8.5 as=0.6369 ps=4.19 w=3.86 l=1.7
X3 VDD1.t4 VP.t1 VTAIL.t7 w_n2594_n1740# sky130_fd_pr__pfet_01v8 ad=0.6369 pd=4.19 as=1.5054 ps=8.5 w=3.86 l=1.7
X4 B.t11 B.t9 B.t10 w_n2594_n1740# sky130_fd_pr__pfet_01v8 ad=1.5054 pd=8.5 as=0 ps=0 w=3.86 l=1.7
X5 VDD2.t3 VN.t2 VTAIL.t1 w_n2594_n1740# sky130_fd_pr__pfet_01v8 ad=1.5054 pd=8.5 as=0.6369 ps=4.19 w=3.86 l=1.7
X6 VTAIL.t8 VP.t2 VDD1.t3 w_n2594_n1740# sky130_fd_pr__pfet_01v8 ad=0.6369 pd=4.19 as=0.6369 ps=4.19 w=3.86 l=1.7
X7 VTAIL.t4 VN.t3 VDD2.t2 w_n2594_n1740# sky130_fd_pr__pfet_01v8 ad=0.6369 pd=4.19 as=0.6369 ps=4.19 w=3.86 l=1.7
X8 VDD1.t2 VP.t3 VTAIL.t10 w_n2594_n1740# sky130_fd_pr__pfet_01v8 ad=1.5054 pd=8.5 as=0.6369 ps=4.19 w=3.86 l=1.7
X9 VDD2.t1 VN.t4 VTAIL.t5 w_n2594_n1740# sky130_fd_pr__pfet_01v8 ad=0.6369 pd=4.19 as=1.5054 ps=8.5 w=3.86 l=1.7
X10 VDD1.t1 VP.t4 VTAIL.t6 w_n2594_n1740# sky130_fd_pr__pfet_01v8 ad=1.5054 pd=8.5 as=0.6369 ps=4.19 w=3.86 l=1.7
X11 VDD2.t0 VN.t5 VTAIL.t2 w_n2594_n1740# sky130_fd_pr__pfet_01v8 ad=0.6369 pd=4.19 as=1.5054 ps=8.5 w=3.86 l=1.7
X12 B.t8 B.t6 B.t7 w_n2594_n1740# sky130_fd_pr__pfet_01v8 ad=1.5054 pd=8.5 as=0 ps=0 w=3.86 l=1.7
X13 B.t5 B.t3 B.t4 w_n2594_n1740# sky130_fd_pr__pfet_01v8 ad=1.5054 pd=8.5 as=0 ps=0 w=3.86 l=1.7
X14 B.t2 B.t0 B.t1 w_n2594_n1740# sky130_fd_pr__pfet_01v8 ad=1.5054 pd=8.5 as=0 ps=0 w=3.86 l=1.7
X15 VTAIL.t11 VP.t5 VDD1.t0 w_n2594_n1740# sky130_fd_pr__pfet_01v8 ad=0.6369 pd=4.19 as=0.6369 ps=4.19 w=3.86 l=1.7
R0 VP.n18 VP.n17 184.417
R1 VP.n33 VP.n32 184.417
R2 VP.n16 VP.n15 184.417
R3 VP.n10 VP.n9 161.3
R4 VP.n11 VP.n6 161.3
R5 VP.n13 VP.n12 161.3
R6 VP.n14 VP.n5 161.3
R7 VP.n31 VP.n0 161.3
R8 VP.n30 VP.n29 161.3
R9 VP.n28 VP.n1 161.3
R10 VP.n27 VP.n26 161.3
R11 VP.n25 VP.n2 161.3
R12 VP.n24 VP.n23 161.3
R13 VP.n22 VP.n3 161.3
R14 VP.n21 VP.n20 161.3
R15 VP.n19 VP.n4 161.3
R16 VP.n7 VP.t3 88.0093
R17 VP.n25 VP.t5 54.7217
R18 VP.n18 VP.t4 54.7217
R19 VP.n32 VP.t1 54.7217
R20 VP.n8 VP.t2 54.7217
R21 VP.n15 VP.t0 54.7217
R22 VP.n8 VP.n7 44.7248
R23 VP.n20 VP.n3 42.0302
R24 VP.n30 VP.n1 42.0302
R25 VP.n13 VP.n6 42.0302
R26 VP.n24 VP.n3 39.1239
R27 VP.n26 VP.n1 39.1239
R28 VP.n9 VP.n6 39.1239
R29 VP.n17 VP.n16 38.8225
R30 VP.n20 VP.n19 24.5923
R31 VP.n25 VP.n24 24.5923
R32 VP.n26 VP.n25 24.5923
R33 VP.n31 VP.n30 24.5923
R34 VP.n14 VP.n13 24.5923
R35 VP.n9 VP.n8 24.5923
R36 VP.n10 VP.n7 12.4115
R37 VP.n19 VP.n18 1.47601
R38 VP.n32 VP.n31 1.47601
R39 VP.n15 VP.n14 1.47601
R40 VP.n11 VP.n10 0.189894
R41 VP.n12 VP.n11 0.189894
R42 VP.n12 VP.n5 0.189894
R43 VP.n16 VP.n5 0.189894
R44 VP.n17 VP.n4 0.189894
R45 VP.n21 VP.n4 0.189894
R46 VP.n22 VP.n21 0.189894
R47 VP.n23 VP.n22 0.189894
R48 VP.n23 VP.n2 0.189894
R49 VP.n27 VP.n2 0.189894
R50 VP.n28 VP.n27 0.189894
R51 VP.n29 VP.n28 0.189894
R52 VP.n29 VP.n0 0.189894
R53 VP.n33 VP.n0 0.189894
R54 VP VP.n33 0.0516364
R55 VTAIL.n82 VTAIL.n68 756.745
R56 VTAIL.n16 VTAIL.n2 756.745
R57 VTAIL.n62 VTAIL.n48 756.745
R58 VTAIL.n40 VTAIL.n26 756.745
R59 VTAIL.n75 VTAIL.n74 585
R60 VTAIL.n72 VTAIL.n71 585
R61 VTAIL.n81 VTAIL.n80 585
R62 VTAIL.n83 VTAIL.n82 585
R63 VTAIL.n9 VTAIL.n8 585
R64 VTAIL.n6 VTAIL.n5 585
R65 VTAIL.n15 VTAIL.n14 585
R66 VTAIL.n17 VTAIL.n16 585
R67 VTAIL.n63 VTAIL.n62 585
R68 VTAIL.n61 VTAIL.n60 585
R69 VTAIL.n52 VTAIL.n51 585
R70 VTAIL.n55 VTAIL.n54 585
R71 VTAIL.n41 VTAIL.n40 585
R72 VTAIL.n39 VTAIL.n38 585
R73 VTAIL.n30 VTAIL.n29 585
R74 VTAIL.n33 VTAIL.n32 585
R75 VTAIL.t2 VTAIL.n73 330.707
R76 VTAIL.t7 VTAIL.n7 330.707
R77 VTAIL.t9 VTAIL.n53 330.707
R78 VTAIL.t5 VTAIL.n31 330.707
R79 VTAIL.n74 VTAIL.n71 171.744
R80 VTAIL.n81 VTAIL.n71 171.744
R81 VTAIL.n82 VTAIL.n81 171.744
R82 VTAIL.n8 VTAIL.n5 171.744
R83 VTAIL.n15 VTAIL.n5 171.744
R84 VTAIL.n16 VTAIL.n15 171.744
R85 VTAIL.n62 VTAIL.n61 171.744
R86 VTAIL.n61 VTAIL.n51 171.744
R87 VTAIL.n54 VTAIL.n51 171.744
R88 VTAIL.n40 VTAIL.n39 171.744
R89 VTAIL.n39 VTAIL.n29 171.744
R90 VTAIL.n32 VTAIL.n29 171.744
R91 VTAIL.n47 VTAIL.n46 97.2774
R92 VTAIL.n25 VTAIL.n24 97.2774
R93 VTAIL.n1 VTAIL.n0 97.2773
R94 VTAIL.n23 VTAIL.n22 97.2773
R95 VTAIL.n74 VTAIL.t2 85.8723
R96 VTAIL.n8 VTAIL.t7 85.8723
R97 VTAIL.n54 VTAIL.t9 85.8723
R98 VTAIL.n32 VTAIL.t5 85.8723
R99 VTAIL.n87 VTAIL.n86 32.5732
R100 VTAIL.n21 VTAIL.n20 32.5732
R101 VTAIL.n67 VTAIL.n66 32.5732
R102 VTAIL.n45 VTAIL.n44 32.5732
R103 VTAIL.n25 VTAIL.n23 19.1945
R104 VTAIL.n87 VTAIL.n67 17.4445
R105 VTAIL.n75 VTAIL.n73 16.3201
R106 VTAIL.n9 VTAIL.n7 16.3201
R107 VTAIL.n55 VTAIL.n53 16.3201
R108 VTAIL.n33 VTAIL.n31 16.3201
R109 VTAIL.n76 VTAIL.n72 12.8005
R110 VTAIL.n10 VTAIL.n6 12.8005
R111 VTAIL.n56 VTAIL.n52 12.8005
R112 VTAIL.n34 VTAIL.n30 12.8005
R113 VTAIL.n80 VTAIL.n79 12.0247
R114 VTAIL.n14 VTAIL.n13 12.0247
R115 VTAIL.n60 VTAIL.n59 12.0247
R116 VTAIL.n38 VTAIL.n37 12.0247
R117 VTAIL.n83 VTAIL.n70 11.249
R118 VTAIL.n17 VTAIL.n4 11.249
R119 VTAIL.n63 VTAIL.n50 11.249
R120 VTAIL.n41 VTAIL.n28 11.249
R121 VTAIL.n84 VTAIL.n68 10.4732
R122 VTAIL.n18 VTAIL.n2 10.4732
R123 VTAIL.n64 VTAIL.n48 10.4732
R124 VTAIL.n42 VTAIL.n26 10.4732
R125 VTAIL.n86 VTAIL.n85 9.45567
R126 VTAIL.n20 VTAIL.n19 9.45567
R127 VTAIL.n66 VTAIL.n65 9.45567
R128 VTAIL.n44 VTAIL.n43 9.45567
R129 VTAIL.n85 VTAIL.n84 9.3005
R130 VTAIL.n70 VTAIL.n69 9.3005
R131 VTAIL.n79 VTAIL.n78 9.3005
R132 VTAIL.n77 VTAIL.n76 9.3005
R133 VTAIL.n19 VTAIL.n18 9.3005
R134 VTAIL.n4 VTAIL.n3 9.3005
R135 VTAIL.n13 VTAIL.n12 9.3005
R136 VTAIL.n11 VTAIL.n10 9.3005
R137 VTAIL.n65 VTAIL.n64 9.3005
R138 VTAIL.n50 VTAIL.n49 9.3005
R139 VTAIL.n59 VTAIL.n58 9.3005
R140 VTAIL.n57 VTAIL.n56 9.3005
R141 VTAIL.n43 VTAIL.n42 9.3005
R142 VTAIL.n28 VTAIL.n27 9.3005
R143 VTAIL.n37 VTAIL.n36 9.3005
R144 VTAIL.n35 VTAIL.n34 9.3005
R145 VTAIL.n0 VTAIL.t1 8.42148
R146 VTAIL.n0 VTAIL.t3 8.42148
R147 VTAIL.n22 VTAIL.t6 8.42148
R148 VTAIL.n22 VTAIL.t11 8.42148
R149 VTAIL.n46 VTAIL.t10 8.42148
R150 VTAIL.n46 VTAIL.t8 8.42148
R151 VTAIL.n24 VTAIL.t0 8.42148
R152 VTAIL.n24 VTAIL.t4 8.42148
R153 VTAIL.n77 VTAIL.n73 3.78097
R154 VTAIL.n11 VTAIL.n7 3.78097
R155 VTAIL.n57 VTAIL.n53 3.78097
R156 VTAIL.n35 VTAIL.n31 3.78097
R157 VTAIL.n86 VTAIL.n68 3.49141
R158 VTAIL.n20 VTAIL.n2 3.49141
R159 VTAIL.n66 VTAIL.n48 3.49141
R160 VTAIL.n44 VTAIL.n26 3.49141
R161 VTAIL.n84 VTAIL.n83 2.71565
R162 VTAIL.n18 VTAIL.n17 2.71565
R163 VTAIL.n64 VTAIL.n63 2.71565
R164 VTAIL.n42 VTAIL.n41 2.71565
R165 VTAIL.n80 VTAIL.n70 1.93989
R166 VTAIL.n14 VTAIL.n4 1.93989
R167 VTAIL.n60 VTAIL.n50 1.93989
R168 VTAIL.n38 VTAIL.n28 1.93989
R169 VTAIL.n45 VTAIL.n25 1.7505
R170 VTAIL.n67 VTAIL.n47 1.7505
R171 VTAIL.n23 VTAIL.n21 1.7505
R172 VTAIL.n47 VTAIL.n45 1.34533
R173 VTAIL.n21 VTAIL.n1 1.34533
R174 VTAIL VTAIL.n87 1.25481
R175 VTAIL.n79 VTAIL.n72 1.16414
R176 VTAIL.n13 VTAIL.n6 1.16414
R177 VTAIL.n59 VTAIL.n52 1.16414
R178 VTAIL.n37 VTAIL.n30 1.16414
R179 VTAIL VTAIL.n1 0.49619
R180 VTAIL.n76 VTAIL.n75 0.388379
R181 VTAIL.n10 VTAIL.n9 0.388379
R182 VTAIL.n56 VTAIL.n55 0.388379
R183 VTAIL.n34 VTAIL.n33 0.388379
R184 VTAIL.n78 VTAIL.n77 0.155672
R185 VTAIL.n78 VTAIL.n69 0.155672
R186 VTAIL.n85 VTAIL.n69 0.155672
R187 VTAIL.n12 VTAIL.n11 0.155672
R188 VTAIL.n12 VTAIL.n3 0.155672
R189 VTAIL.n19 VTAIL.n3 0.155672
R190 VTAIL.n65 VTAIL.n49 0.155672
R191 VTAIL.n58 VTAIL.n49 0.155672
R192 VTAIL.n58 VTAIL.n57 0.155672
R193 VTAIL.n43 VTAIL.n27 0.155672
R194 VTAIL.n36 VTAIL.n27 0.155672
R195 VTAIL.n36 VTAIL.n35 0.155672
R196 VDD1.n14 VDD1.n0 756.745
R197 VDD1.n33 VDD1.n19 756.745
R198 VDD1.n15 VDD1.n14 585
R199 VDD1.n13 VDD1.n12 585
R200 VDD1.n4 VDD1.n3 585
R201 VDD1.n7 VDD1.n6 585
R202 VDD1.n26 VDD1.n25 585
R203 VDD1.n23 VDD1.n22 585
R204 VDD1.n32 VDD1.n31 585
R205 VDD1.n34 VDD1.n33 585
R206 VDD1.t2 VDD1.n5 330.707
R207 VDD1.t1 VDD1.n24 330.707
R208 VDD1.n14 VDD1.n13 171.744
R209 VDD1.n13 VDD1.n3 171.744
R210 VDD1.n6 VDD1.n3 171.744
R211 VDD1.n25 VDD1.n22 171.744
R212 VDD1.n32 VDD1.n22 171.744
R213 VDD1.n33 VDD1.n32 171.744
R214 VDD1.n39 VDD1.n38 114.338
R215 VDD1.n41 VDD1.n40 113.957
R216 VDD1.n6 VDD1.t2 85.8723
R217 VDD1.n25 VDD1.t1 85.8723
R218 VDD1 VDD1.n18 50.6227
R219 VDD1.n39 VDD1.n37 50.5092
R220 VDD1.n41 VDD1.n39 34.1884
R221 VDD1.n7 VDD1.n5 16.3201
R222 VDD1.n26 VDD1.n24 16.3201
R223 VDD1.n8 VDD1.n4 12.8005
R224 VDD1.n27 VDD1.n23 12.8005
R225 VDD1.n12 VDD1.n11 12.0247
R226 VDD1.n31 VDD1.n30 12.0247
R227 VDD1.n15 VDD1.n2 11.249
R228 VDD1.n34 VDD1.n21 11.249
R229 VDD1.n16 VDD1.n0 10.4732
R230 VDD1.n35 VDD1.n19 10.4732
R231 VDD1.n18 VDD1.n17 9.45567
R232 VDD1.n37 VDD1.n36 9.45567
R233 VDD1.n17 VDD1.n16 9.3005
R234 VDD1.n2 VDD1.n1 9.3005
R235 VDD1.n11 VDD1.n10 9.3005
R236 VDD1.n9 VDD1.n8 9.3005
R237 VDD1.n36 VDD1.n35 9.3005
R238 VDD1.n21 VDD1.n20 9.3005
R239 VDD1.n30 VDD1.n29 9.3005
R240 VDD1.n28 VDD1.n27 9.3005
R241 VDD1.n40 VDD1.t3 8.42148
R242 VDD1.n40 VDD1.t5 8.42148
R243 VDD1.n38 VDD1.t0 8.42148
R244 VDD1.n38 VDD1.t4 8.42148
R245 VDD1.n9 VDD1.n5 3.78097
R246 VDD1.n28 VDD1.n24 3.78097
R247 VDD1.n18 VDD1.n0 3.49141
R248 VDD1.n37 VDD1.n19 3.49141
R249 VDD1.n16 VDD1.n15 2.71565
R250 VDD1.n35 VDD1.n34 2.71565
R251 VDD1.n12 VDD1.n2 1.93989
R252 VDD1.n31 VDD1.n21 1.93989
R253 VDD1.n11 VDD1.n4 1.16414
R254 VDD1.n30 VDD1.n23 1.16414
R255 VDD1.n8 VDD1.n7 0.388379
R256 VDD1.n27 VDD1.n26 0.388379
R257 VDD1 VDD1.n41 0.37981
R258 VDD1.n17 VDD1.n1 0.155672
R259 VDD1.n10 VDD1.n1 0.155672
R260 VDD1.n10 VDD1.n9 0.155672
R261 VDD1.n29 VDD1.n28 0.155672
R262 VDD1.n29 VDD1.n20 0.155672
R263 VDD1.n36 VDD1.n20 0.155672
R264 VN.n11 VN.n10 184.417
R265 VN.n23 VN.n22 184.417
R266 VN.n21 VN.n12 161.3
R267 VN.n20 VN.n19 161.3
R268 VN.n18 VN.n13 161.3
R269 VN.n17 VN.n16 161.3
R270 VN.n9 VN.n0 161.3
R271 VN.n8 VN.n7 161.3
R272 VN.n6 VN.n1 161.3
R273 VN.n5 VN.n4 161.3
R274 VN.n2 VN.t2 88.0093
R275 VN.n14 VN.t4 88.0093
R276 VN.n3 VN.t0 54.7217
R277 VN.n10 VN.t5 54.7217
R278 VN.n15 VN.t3 54.7217
R279 VN.n22 VN.t1 54.7217
R280 VN.n15 VN.n14 44.7248
R281 VN.n3 VN.n2 44.7248
R282 VN.n8 VN.n1 42.0302
R283 VN.n20 VN.n13 42.0302
R284 VN VN.n23 39.2032
R285 VN.n4 VN.n1 39.1239
R286 VN.n16 VN.n13 39.1239
R287 VN.n4 VN.n3 24.5923
R288 VN.n9 VN.n8 24.5923
R289 VN.n16 VN.n15 24.5923
R290 VN.n21 VN.n20 24.5923
R291 VN.n17 VN.n14 12.4115
R292 VN.n5 VN.n2 12.4115
R293 VN.n10 VN.n9 1.47601
R294 VN.n22 VN.n21 1.47601
R295 VN.n23 VN.n12 0.189894
R296 VN.n19 VN.n12 0.189894
R297 VN.n19 VN.n18 0.189894
R298 VN.n18 VN.n17 0.189894
R299 VN.n6 VN.n5 0.189894
R300 VN.n7 VN.n6 0.189894
R301 VN.n7 VN.n0 0.189894
R302 VN.n11 VN.n0 0.189894
R303 VN VN.n11 0.0516364
R304 VDD2.n35 VDD2.n21 756.745
R305 VDD2.n14 VDD2.n0 756.745
R306 VDD2.n36 VDD2.n35 585
R307 VDD2.n34 VDD2.n33 585
R308 VDD2.n25 VDD2.n24 585
R309 VDD2.n28 VDD2.n27 585
R310 VDD2.n7 VDD2.n6 585
R311 VDD2.n4 VDD2.n3 585
R312 VDD2.n13 VDD2.n12 585
R313 VDD2.n15 VDD2.n14 585
R314 VDD2.t4 VDD2.n26 330.707
R315 VDD2.t3 VDD2.n5 330.707
R316 VDD2.n35 VDD2.n34 171.744
R317 VDD2.n34 VDD2.n24 171.744
R318 VDD2.n27 VDD2.n24 171.744
R319 VDD2.n6 VDD2.n3 171.744
R320 VDD2.n13 VDD2.n3 171.744
R321 VDD2.n14 VDD2.n13 171.744
R322 VDD2.n20 VDD2.n19 114.338
R323 VDD2 VDD2.n41 114.335
R324 VDD2.n27 VDD2.t4 85.8723
R325 VDD2.n6 VDD2.t3 85.8723
R326 VDD2.n20 VDD2.n18 50.5092
R327 VDD2.n40 VDD2.n39 49.252
R328 VDD2.n40 VDD2.n20 32.7304
R329 VDD2.n28 VDD2.n26 16.3201
R330 VDD2.n7 VDD2.n5 16.3201
R331 VDD2.n29 VDD2.n25 12.8005
R332 VDD2.n8 VDD2.n4 12.8005
R333 VDD2.n33 VDD2.n32 12.0247
R334 VDD2.n12 VDD2.n11 12.0247
R335 VDD2.n36 VDD2.n23 11.249
R336 VDD2.n15 VDD2.n2 11.249
R337 VDD2.n37 VDD2.n21 10.4732
R338 VDD2.n16 VDD2.n0 10.4732
R339 VDD2.n39 VDD2.n38 9.45567
R340 VDD2.n18 VDD2.n17 9.45567
R341 VDD2.n38 VDD2.n37 9.3005
R342 VDD2.n23 VDD2.n22 9.3005
R343 VDD2.n32 VDD2.n31 9.3005
R344 VDD2.n30 VDD2.n29 9.3005
R345 VDD2.n17 VDD2.n16 9.3005
R346 VDD2.n2 VDD2.n1 9.3005
R347 VDD2.n11 VDD2.n10 9.3005
R348 VDD2.n9 VDD2.n8 9.3005
R349 VDD2.n41 VDD2.t2 8.42148
R350 VDD2.n41 VDD2.t1 8.42148
R351 VDD2.n19 VDD2.t5 8.42148
R352 VDD2.n19 VDD2.t0 8.42148
R353 VDD2.n30 VDD2.n26 3.78097
R354 VDD2.n9 VDD2.n5 3.78097
R355 VDD2.n39 VDD2.n21 3.49141
R356 VDD2.n18 VDD2.n0 3.49141
R357 VDD2.n37 VDD2.n36 2.71565
R358 VDD2.n16 VDD2.n15 2.71565
R359 VDD2.n33 VDD2.n23 1.93989
R360 VDD2.n12 VDD2.n2 1.93989
R361 VDD2 VDD2.n40 1.37119
R362 VDD2.n32 VDD2.n25 1.16414
R363 VDD2.n11 VDD2.n4 1.16414
R364 VDD2.n29 VDD2.n28 0.388379
R365 VDD2.n8 VDD2.n7 0.388379
R366 VDD2.n38 VDD2.n22 0.155672
R367 VDD2.n31 VDD2.n22 0.155672
R368 VDD2.n31 VDD2.n30 0.155672
R369 VDD2.n10 VDD2.n9 0.155672
R370 VDD2.n10 VDD2.n1 0.155672
R371 VDD2.n17 VDD2.n1 0.155672
R372 B.n333 B.n44 585
R373 B.n335 B.n334 585
R374 B.n336 B.n43 585
R375 B.n338 B.n337 585
R376 B.n339 B.n42 585
R377 B.n341 B.n340 585
R378 B.n342 B.n41 585
R379 B.n344 B.n343 585
R380 B.n345 B.n40 585
R381 B.n347 B.n346 585
R382 B.n348 B.n39 585
R383 B.n350 B.n349 585
R384 B.n351 B.n38 585
R385 B.n353 B.n352 585
R386 B.n354 B.n37 585
R387 B.n356 B.n355 585
R388 B.n357 B.n36 585
R389 B.n359 B.n358 585
R390 B.n361 B.n33 585
R391 B.n363 B.n362 585
R392 B.n364 B.n32 585
R393 B.n366 B.n365 585
R394 B.n367 B.n31 585
R395 B.n369 B.n368 585
R396 B.n370 B.n30 585
R397 B.n372 B.n371 585
R398 B.n373 B.n27 585
R399 B.n376 B.n375 585
R400 B.n377 B.n26 585
R401 B.n379 B.n378 585
R402 B.n380 B.n25 585
R403 B.n382 B.n381 585
R404 B.n383 B.n24 585
R405 B.n385 B.n384 585
R406 B.n386 B.n23 585
R407 B.n388 B.n387 585
R408 B.n389 B.n22 585
R409 B.n391 B.n390 585
R410 B.n392 B.n21 585
R411 B.n394 B.n393 585
R412 B.n395 B.n20 585
R413 B.n397 B.n396 585
R414 B.n398 B.n19 585
R415 B.n400 B.n399 585
R416 B.n401 B.n18 585
R417 B.n332 B.n331 585
R418 B.n330 B.n45 585
R419 B.n329 B.n328 585
R420 B.n327 B.n46 585
R421 B.n326 B.n325 585
R422 B.n324 B.n47 585
R423 B.n323 B.n322 585
R424 B.n321 B.n48 585
R425 B.n320 B.n319 585
R426 B.n318 B.n49 585
R427 B.n317 B.n316 585
R428 B.n315 B.n50 585
R429 B.n314 B.n313 585
R430 B.n312 B.n51 585
R431 B.n311 B.n310 585
R432 B.n309 B.n52 585
R433 B.n308 B.n307 585
R434 B.n306 B.n53 585
R435 B.n305 B.n304 585
R436 B.n303 B.n54 585
R437 B.n302 B.n301 585
R438 B.n300 B.n55 585
R439 B.n299 B.n298 585
R440 B.n297 B.n56 585
R441 B.n296 B.n295 585
R442 B.n294 B.n57 585
R443 B.n293 B.n292 585
R444 B.n291 B.n58 585
R445 B.n290 B.n289 585
R446 B.n288 B.n59 585
R447 B.n287 B.n286 585
R448 B.n285 B.n60 585
R449 B.n284 B.n283 585
R450 B.n282 B.n61 585
R451 B.n281 B.n280 585
R452 B.n279 B.n62 585
R453 B.n278 B.n277 585
R454 B.n276 B.n63 585
R455 B.n275 B.n274 585
R456 B.n273 B.n64 585
R457 B.n272 B.n271 585
R458 B.n270 B.n65 585
R459 B.n269 B.n268 585
R460 B.n267 B.n66 585
R461 B.n266 B.n265 585
R462 B.n264 B.n67 585
R463 B.n263 B.n262 585
R464 B.n261 B.n68 585
R465 B.n260 B.n259 585
R466 B.n258 B.n69 585
R467 B.n257 B.n256 585
R468 B.n255 B.n70 585
R469 B.n254 B.n253 585
R470 B.n252 B.n71 585
R471 B.n251 B.n250 585
R472 B.n249 B.n72 585
R473 B.n248 B.n247 585
R474 B.n246 B.n73 585
R475 B.n245 B.n244 585
R476 B.n243 B.n74 585
R477 B.n242 B.n241 585
R478 B.n240 B.n75 585
R479 B.n239 B.n238 585
R480 B.n237 B.n76 585
R481 B.n236 B.n235 585
R482 B.n167 B.n166 585
R483 B.n168 B.n103 585
R484 B.n170 B.n169 585
R485 B.n171 B.n102 585
R486 B.n173 B.n172 585
R487 B.n174 B.n101 585
R488 B.n176 B.n175 585
R489 B.n177 B.n100 585
R490 B.n179 B.n178 585
R491 B.n180 B.n99 585
R492 B.n182 B.n181 585
R493 B.n183 B.n98 585
R494 B.n185 B.n184 585
R495 B.n186 B.n97 585
R496 B.n188 B.n187 585
R497 B.n189 B.n96 585
R498 B.n191 B.n190 585
R499 B.n192 B.n93 585
R500 B.n195 B.n194 585
R501 B.n196 B.n92 585
R502 B.n198 B.n197 585
R503 B.n199 B.n91 585
R504 B.n201 B.n200 585
R505 B.n202 B.n90 585
R506 B.n204 B.n203 585
R507 B.n205 B.n89 585
R508 B.n207 B.n206 585
R509 B.n209 B.n208 585
R510 B.n210 B.n85 585
R511 B.n212 B.n211 585
R512 B.n213 B.n84 585
R513 B.n215 B.n214 585
R514 B.n216 B.n83 585
R515 B.n218 B.n217 585
R516 B.n219 B.n82 585
R517 B.n221 B.n220 585
R518 B.n222 B.n81 585
R519 B.n224 B.n223 585
R520 B.n225 B.n80 585
R521 B.n227 B.n226 585
R522 B.n228 B.n79 585
R523 B.n230 B.n229 585
R524 B.n231 B.n78 585
R525 B.n233 B.n232 585
R526 B.n234 B.n77 585
R527 B.n165 B.n104 585
R528 B.n164 B.n163 585
R529 B.n162 B.n105 585
R530 B.n161 B.n160 585
R531 B.n159 B.n106 585
R532 B.n158 B.n157 585
R533 B.n156 B.n107 585
R534 B.n155 B.n154 585
R535 B.n153 B.n108 585
R536 B.n152 B.n151 585
R537 B.n150 B.n109 585
R538 B.n149 B.n148 585
R539 B.n147 B.n110 585
R540 B.n146 B.n145 585
R541 B.n144 B.n111 585
R542 B.n143 B.n142 585
R543 B.n141 B.n112 585
R544 B.n140 B.n139 585
R545 B.n138 B.n113 585
R546 B.n137 B.n136 585
R547 B.n135 B.n114 585
R548 B.n134 B.n133 585
R549 B.n132 B.n115 585
R550 B.n131 B.n130 585
R551 B.n129 B.n116 585
R552 B.n128 B.n127 585
R553 B.n126 B.n117 585
R554 B.n125 B.n124 585
R555 B.n123 B.n118 585
R556 B.n122 B.n121 585
R557 B.n120 B.n119 585
R558 B.n2 B.n0 585
R559 B.n449 B.n1 585
R560 B.n448 B.n447 585
R561 B.n446 B.n3 585
R562 B.n445 B.n444 585
R563 B.n443 B.n4 585
R564 B.n442 B.n441 585
R565 B.n440 B.n5 585
R566 B.n439 B.n438 585
R567 B.n437 B.n6 585
R568 B.n436 B.n435 585
R569 B.n434 B.n7 585
R570 B.n433 B.n432 585
R571 B.n431 B.n8 585
R572 B.n430 B.n429 585
R573 B.n428 B.n9 585
R574 B.n427 B.n426 585
R575 B.n425 B.n10 585
R576 B.n424 B.n423 585
R577 B.n422 B.n11 585
R578 B.n421 B.n420 585
R579 B.n419 B.n12 585
R580 B.n418 B.n417 585
R581 B.n416 B.n13 585
R582 B.n415 B.n414 585
R583 B.n413 B.n14 585
R584 B.n412 B.n411 585
R585 B.n410 B.n15 585
R586 B.n409 B.n408 585
R587 B.n407 B.n16 585
R588 B.n406 B.n405 585
R589 B.n404 B.n17 585
R590 B.n403 B.n402 585
R591 B.n451 B.n450 585
R592 B.n166 B.n165 492.5
R593 B.n402 B.n401 492.5
R594 B.n236 B.n77 492.5
R595 B.n333 B.n332 492.5
R596 B.n86 B.t11 272.284
R597 B.n34 B.t1 272.284
R598 B.n94 B.t8 272.284
R599 B.n28 B.t4 272.284
R600 B.n86 B.t9 260.836
R601 B.n94 B.t6 260.836
R602 B.n28 B.t3 260.836
R603 B.n34 B.t0 260.836
R604 B.n87 B.t10 232.915
R605 B.n35 B.t2 232.915
R606 B.n95 B.t7 232.915
R607 B.n29 B.t5 232.915
R608 B.n165 B.n164 163.367
R609 B.n164 B.n105 163.367
R610 B.n160 B.n105 163.367
R611 B.n160 B.n159 163.367
R612 B.n159 B.n158 163.367
R613 B.n158 B.n107 163.367
R614 B.n154 B.n107 163.367
R615 B.n154 B.n153 163.367
R616 B.n153 B.n152 163.367
R617 B.n152 B.n109 163.367
R618 B.n148 B.n109 163.367
R619 B.n148 B.n147 163.367
R620 B.n147 B.n146 163.367
R621 B.n146 B.n111 163.367
R622 B.n142 B.n111 163.367
R623 B.n142 B.n141 163.367
R624 B.n141 B.n140 163.367
R625 B.n140 B.n113 163.367
R626 B.n136 B.n113 163.367
R627 B.n136 B.n135 163.367
R628 B.n135 B.n134 163.367
R629 B.n134 B.n115 163.367
R630 B.n130 B.n115 163.367
R631 B.n130 B.n129 163.367
R632 B.n129 B.n128 163.367
R633 B.n128 B.n117 163.367
R634 B.n124 B.n117 163.367
R635 B.n124 B.n123 163.367
R636 B.n123 B.n122 163.367
R637 B.n122 B.n119 163.367
R638 B.n119 B.n2 163.367
R639 B.n450 B.n2 163.367
R640 B.n450 B.n449 163.367
R641 B.n449 B.n448 163.367
R642 B.n448 B.n3 163.367
R643 B.n444 B.n3 163.367
R644 B.n444 B.n443 163.367
R645 B.n443 B.n442 163.367
R646 B.n442 B.n5 163.367
R647 B.n438 B.n5 163.367
R648 B.n438 B.n437 163.367
R649 B.n437 B.n436 163.367
R650 B.n436 B.n7 163.367
R651 B.n432 B.n7 163.367
R652 B.n432 B.n431 163.367
R653 B.n431 B.n430 163.367
R654 B.n430 B.n9 163.367
R655 B.n426 B.n9 163.367
R656 B.n426 B.n425 163.367
R657 B.n425 B.n424 163.367
R658 B.n424 B.n11 163.367
R659 B.n420 B.n11 163.367
R660 B.n420 B.n419 163.367
R661 B.n419 B.n418 163.367
R662 B.n418 B.n13 163.367
R663 B.n414 B.n13 163.367
R664 B.n414 B.n413 163.367
R665 B.n413 B.n412 163.367
R666 B.n412 B.n15 163.367
R667 B.n408 B.n15 163.367
R668 B.n408 B.n407 163.367
R669 B.n407 B.n406 163.367
R670 B.n406 B.n17 163.367
R671 B.n402 B.n17 163.367
R672 B.n166 B.n103 163.367
R673 B.n170 B.n103 163.367
R674 B.n171 B.n170 163.367
R675 B.n172 B.n171 163.367
R676 B.n172 B.n101 163.367
R677 B.n176 B.n101 163.367
R678 B.n177 B.n176 163.367
R679 B.n178 B.n177 163.367
R680 B.n178 B.n99 163.367
R681 B.n182 B.n99 163.367
R682 B.n183 B.n182 163.367
R683 B.n184 B.n183 163.367
R684 B.n184 B.n97 163.367
R685 B.n188 B.n97 163.367
R686 B.n189 B.n188 163.367
R687 B.n190 B.n189 163.367
R688 B.n190 B.n93 163.367
R689 B.n195 B.n93 163.367
R690 B.n196 B.n195 163.367
R691 B.n197 B.n196 163.367
R692 B.n197 B.n91 163.367
R693 B.n201 B.n91 163.367
R694 B.n202 B.n201 163.367
R695 B.n203 B.n202 163.367
R696 B.n203 B.n89 163.367
R697 B.n207 B.n89 163.367
R698 B.n208 B.n207 163.367
R699 B.n208 B.n85 163.367
R700 B.n212 B.n85 163.367
R701 B.n213 B.n212 163.367
R702 B.n214 B.n213 163.367
R703 B.n214 B.n83 163.367
R704 B.n218 B.n83 163.367
R705 B.n219 B.n218 163.367
R706 B.n220 B.n219 163.367
R707 B.n220 B.n81 163.367
R708 B.n224 B.n81 163.367
R709 B.n225 B.n224 163.367
R710 B.n226 B.n225 163.367
R711 B.n226 B.n79 163.367
R712 B.n230 B.n79 163.367
R713 B.n231 B.n230 163.367
R714 B.n232 B.n231 163.367
R715 B.n232 B.n77 163.367
R716 B.n237 B.n236 163.367
R717 B.n238 B.n237 163.367
R718 B.n238 B.n75 163.367
R719 B.n242 B.n75 163.367
R720 B.n243 B.n242 163.367
R721 B.n244 B.n243 163.367
R722 B.n244 B.n73 163.367
R723 B.n248 B.n73 163.367
R724 B.n249 B.n248 163.367
R725 B.n250 B.n249 163.367
R726 B.n250 B.n71 163.367
R727 B.n254 B.n71 163.367
R728 B.n255 B.n254 163.367
R729 B.n256 B.n255 163.367
R730 B.n256 B.n69 163.367
R731 B.n260 B.n69 163.367
R732 B.n261 B.n260 163.367
R733 B.n262 B.n261 163.367
R734 B.n262 B.n67 163.367
R735 B.n266 B.n67 163.367
R736 B.n267 B.n266 163.367
R737 B.n268 B.n267 163.367
R738 B.n268 B.n65 163.367
R739 B.n272 B.n65 163.367
R740 B.n273 B.n272 163.367
R741 B.n274 B.n273 163.367
R742 B.n274 B.n63 163.367
R743 B.n278 B.n63 163.367
R744 B.n279 B.n278 163.367
R745 B.n280 B.n279 163.367
R746 B.n280 B.n61 163.367
R747 B.n284 B.n61 163.367
R748 B.n285 B.n284 163.367
R749 B.n286 B.n285 163.367
R750 B.n286 B.n59 163.367
R751 B.n290 B.n59 163.367
R752 B.n291 B.n290 163.367
R753 B.n292 B.n291 163.367
R754 B.n292 B.n57 163.367
R755 B.n296 B.n57 163.367
R756 B.n297 B.n296 163.367
R757 B.n298 B.n297 163.367
R758 B.n298 B.n55 163.367
R759 B.n302 B.n55 163.367
R760 B.n303 B.n302 163.367
R761 B.n304 B.n303 163.367
R762 B.n304 B.n53 163.367
R763 B.n308 B.n53 163.367
R764 B.n309 B.n308 163.367
R765 B.n310 B.n309 163.367
R766 B.n310 B.n51 163.367
R767 B.n314 B.n51 163.367
R768 B.n315 B.n314 163.367
R769 B.n316 B.n315 163.367
R770 B.n316 B.n49 163.367
R771 B.n320 B.n49 163.367
R772 B.n321 B.n320 163.367
R773 B.n322 B.n321 163.367
R774 B.n322 B.n47 163.367
R775 B.n326 B.n47 163.367
R776 B.n327 B.n326 163.367
R777 B.n328 B.n327 163.367
R778 B.n328 B.n45 163.367
R779 B.n332 B.n45 163.367
R780 B.n401 B.n400 163.367
R781 B.n400 B.n19 163.367
R782 B.n396 B.n19 163.367
R783 B.n396 B.n395 163.367
R784 B.n395 B.n394 163.367
R785 B.n394 B.n21 163.367
R786 B.n390 B.n21 163.367
R787 B.n390 B.n389 163.367
R788 B.n389 B.n388 163.367
R789 B.n388 B.n23 163.367
R790 B.n384 B.n23 163.367
R791 B.n384 B.n383 163.367
R792 B.n383 B.n382 163.367
R793 B.n382 B.n25 163.367
R794 B.n378 B.n25 163.367
R795 B.n378 B.n377 163.367
R796 B.n377 B.n376 163.367
R797 B.n376 B.n27 163.367
R798 B.n371 B.n27 163.367
R799 B.n371 B.n370 163.367
R800 B.n370 B.n369 163.367
R801 B.n369 B.n31 163.367
R802 B.n365 B.n31 163.367
R803 B.n365 B.n364 163.367
R804 B.n364 B.n363 163.367
R805 B.n363 B.n33 163.367
R806 B.n358 B.n33 163.367
R807 B.n358 B.n357 163.367
R808 B.n357 B.n356 163.367
R809 B.n356 B.n37 163.367
R810 B.n352 B.n37 163.367
R811 B.n352 B.n351 163.367
R812 B.n351 B.n350 163.367
R813 B.n350 B.n39 163.367
R814 B.n346 B.n39 163.367
R815 B.n346 B.n345 163.367
R816 B.n345 B.n344 163.367
R817 B.n344 B.n41 163.367
R818 B.n340 B.n41 163.367
R819 B.n340 B.n339 163.367
R820 B.n339 B.n338 163.367
R821 B.n338 B.n43 163.367
R822 B.n334 B.n43 163.367
R823 B.n334 B.n333 163.367
R824 B.n88 B.n87 59.5399
R825 B.n193 B.n95 59.5399
R826 B.n374 B.n29 59.5399
R827 B.n360 B.n35 59.5399
R828 B.n87 B.n86 39.3702
R829 B.n95 B.n94 39.3702
R830 B.n29 B.n28 39.3702
R831 B.n35 B.n34 39.3702
R832 B.n403 B.n18 32.0005
R833 B.n331 B.n44 32.0005
R834 B.n235 B.n234 32.0005
R835 B.n167 B.n104 32.0005
R836 B B.n451 18.0485
R837 B.n399 B.n18 10.6151
R838 B.n399 B.n398 10.6151
R839 B.n398 B.n397 10.6151
R840 B.n397 B.n20 10.6151
R841 B.n393 B.n20 10.6151
R842 B.n393 B.n392 10.6151
R843 B.n392 B.n391 10.6151
R844 B.n391 B.n22 10.6151
R845 B.n387 B.n22 10.6151
R846 B.n387 B.n386 10.6151
R847 B.n386 B.n385 10.6151
R848 B.n385 B.n24 10.6151
R849 B.n381 B.n24 10.6151
R850 B.n381 B.n380 10.6151
R851 B.n380 B.n379 10.6151
R852 B.n379 B.n26 10.6151
R853 B.n375 B.n26 10.6151
R854 B.n373 B.n372 10.6151
R855 B.n372 B.n30 10.6151
R856 B.n368 B.n30 10.6151
R857 B.n368 B.n367 10.6151
R858 B.n367 B.n366 10.6151
R859 B.n366 B.n32 10.6151
R860 B.n362 B.n32 10.6151
R861 B.n362 B.n361 10.6151
R862 B.n359 B.n36 10.6151
R863 B.n355 B.n36 10.6151
R864 B.n355 B.n354 10.6151
R865 B.n354 B.n353 10.6151
R866 B.n353 B.n38 10.6151
R867 B.n349 B.n38 10.6151
R868 B.n349 B.n348 10.6151
R869 B.n348 B.n347 10.6151
R870 B.n347 B.n40 10.6151
R871 B.n343 B.n40 10.6151
R872 B.n343 B.n342 10.6151
R873 B.n342 B.n341 10.6151
R874 B.n341 B.n42 10.6151
R875 B.n337 B.n42 10.6151
R876 B.n337 B.n336 10.6151
R877 B.n336 B.n335 10.6151
R878 B.n335 B.n44 10.6151
R879 B.n235 B.n76 10.6151
R880 B.n239 B.n76 10.6151
R881 B.n240 B.n239 10.6151
R882 B.n241 B.n240 10.6151
R883 B.n241 B.n74 10.6151
R884 B.n245 B.n74 10.6151
R885 B.n246 B.n245 10.6151
R886 B.n247 B.n246 10.6151
R887 B.n247 B.n72 10.6151
R888 B.n251 B.n72 10.6151
R889 B.n252 B.n251 10.6151
R890 B.n253 B.n252 10.6151
R891 B.n253 B.n70 10.6151
R892 B.n257 B.n70 10.6151
R893 B.n258 B.n257 10.6151
R894 B.n259 B.n258 10.6151
R895 B.n259 B.n68 10.6151
R896 B.n263 B.n68 10.6151
R897 B.n264 B.n263 10.6151
R898 B.n265 B.n264 10.6151
R899 B.n265 B.n66 10.6151
R900 B.n269 B.n66 10.6151
R901 B.n270 B.n269 10.6151
R902 B.n271 B.n270 10.6151
R903 B.n271 B.n64 10.6151
R904 B.n275 B.n64 10.6151
R905 B.n276 B.n275 10.6151
R906 B.n277 B.n276 10.6151
R907 B.n277 B.n62 10.6151
R908 B.n281 B.n62 10.6151
R909 B.n282 B.n281 10.6151
R910 B.n283 B.n282 10.6151
R911 B.n283 B.n60 10.6151
R912 B.n287 B.n60 10.6151
R913 B.n288 B.n287 10.6151
R914 B.n289 B.n288 10.6151
R915 B.n289 B.n58 10.6151
R916 B.n293 B.n58 10.6151
R917 B.n294 B.n293 10.6151
R918 B.n295 B.n294 10.6151
R919 B.n295 B.n56 10.6151
R920 B.n299 B.n56 10.6151
R921 B.n300 B.n299 10.6151
R922 B.n301 B.n300 10.6151
R923 B.n301 B.n54 10.6151
R924 B.n305 B.n54 10.6151
R925 B.n306 B.n305 10.6151
R926 B.n307 B.n306 10.6151
R927 B.n307 B.n52 10.6151
R928 B.n311 B.n52 10.6151
R929 B.n312 B.n311 10.6151
R930 B.n313 B.n312 10.6151
R931 B.n313 B.n50 10.6151
R932 B.n317 B.n50 10.6151
R933 B.n318 B.n317 10.6151
R934 B.n319 B.n318 10.6151
R935 B.n319 B.n48 10.6151
R936 B.n323 B.n48 10.6151
R937 B.n324 B.n323 10.6151
R938 B.n325 B.n324 10.6151
R939 B.n325 B.n46 10.6151
R940 B.n329 B.n46 10.6151
R941 B.n330 B.n329 10.6151
R942 B.n331 B.n330 10.6151
R943 B.n168 B.n167 10.6151
R944 B.n169 B.n168 10.6151
R945 B.n169 B.n102 10.6151
R946 B.n173 B.n102 10.6151
R947 B.n174 B.n173 10.6151
R948 B.n175 B.n174 10.6151
R949 B.n175 B.n100 10.6151
R950 B.n179 B.n100 10.6151
R951 B.n180 B.n179 10.6151
R952 B.n181 B.n180 10.6151
R953 B.n181 B.n98 10.6151
R954 B.n185 B.n98 10.6151
R955 B.n186 B.n185 10.6151
R956 B.n187 B.n186 10.6151
R957 B.n187 B.n96 10.6151
R958 B.n191 B.n96 10.6151
R959 B.n192 B.n191 10.6151
R960 B.n194 B.n92 10.6151
R961 B.n198 B.n92 10.6151
R962 B.n199 B.n198 10.6151
R963 B.n200 B.n199 10.6151
R964 B.n200 B.n90 10.6151
R965 B.n204 B.n90 10.6151
R966 B.n205 B.n204 10.6151
R967 B.n206 B.n205 10.6151
R968 B.n210 B.n209 10.6151
R969 B.n211 B.n210 10.6151
R970 B.n211 B.n84 10.6151
R971 B.n215 B.n84 10.6151
R972 B.n216 B.n215 10.6151
R973 B.n217 B.n216 10.6151
R974 B.n217 B.n82 10.6151
R975 B.n221 B.n82 10.6151
R976 B.n222 B.n221 10.6151
R977 B.n223 B.n222 10.6151
R978 B.n223 B.n80 10.6151
R979 B.n227 B.n80 10.6151
R980 B.n228 B.n227 10.6151
R981 B.n229 B.n228 10.6151
R982 B.n229 B.n78 10.6151
R983 B.n233 B.n78 10.6151
R984 B.n234 B.n233 10.6151
R985 B.n163 B.n104 10.6151
R986 B.n163 B.n162 10.6151
R987 B.n162 B.n161 10.6151
R988 B.n161 B.n106 10.6151
R989 B.n157 B.n106 10.6151
R990 B.n157 B.n156 10.6151
R991 B.n156 B.n155 10.6151
R992 B.n155 B.n108 10.6151
R993 B.n151 B.n108 10.6151
R994 B.n151 B.n150 10.6151
R995 B.n150 B.n149 10.6151
R996 B.n149 B.n110 10.6151
R997 B.n145 B.n110 10.6151
R998 B.n145 B.n144 10.6151
R999 B.n144 B.n143 10.6151
R1000 B.n143 B.n112 10.6151
R1001 B.n139 B.n112 10.6151
R1002 B.n139 B.n138 10.6151
R1003 B.n138 B.n137 10.6151
R1004 B.n137 B.n114 10.6151
R1005 B.n133 B.n114 10.6151
R1006 B.n133 B.n132 10.6151
R1007 B.n132 B.n131 10.6151
R1008 B.n131 B.n116 10.6151
R1009 B.n127 B.n116 10.6151
R1010 B.n127 B.n126 10.6151
R1011 B.n126 B.n125 10.6151
R1012 B.n125 B.n118 10.6151
R1013 B.n121 B.n118 10.6151
R1014 B.n121 B.n120 10.6151
R1015 B.n120 B.n0 10.6151
R1016 B.n447 B.n1 10.6151
R1017 B.n447 B.n446 10.6151
R1018 B.n446 B.n445 10.6151
R1019 B.n445 B.n4 10.6151
R1020 B.n441 B.n4 10.6151
R1021 B.n441 B.n440 10.6151
R1022 B.n440 B.n439 10.6151
R1023 B.n439 B.n6 10.6151
R1024 B.n435 B.n6 10.6151
R1025 B.n435 B.n434 10.6151
R1026 B.n434 B.n433 10.6151
R1027 B.n433 B.n8 10.6151
R1028 B.n429 B.n8 10.6151
R1029 B.n429 B.n428 10.6151
R1030 B.n428 B.n427 10.6151
R1031 B.n427 B.n10 10.6151
R1032 B.n423 B.n10 10.6151
R1033 B.n423 B.n422 10.6151
R1034 B.n422 B.n421 10.6151
R1035 B.n421 B.n12 10.6151
R1036 B.n417 B.n12 10.6151
R1037 B.n417 B.n416 10.6151
R1038 B.n416 B.n415 10.6151
R1039 B.n415 B.n14 10.6151
R1040 B.n411 B.n14 10.6151
R1041 B.n411 B.n410 10.6151
R1042 B.n410 B.n409 10.6151
R1043 B.n409 B.n16 10.6151
R1044 B.n405 B.n16 10.6151
R1045 B.n405 B.n404 10.6151
R1046 B.n404 B.n403 10.6151
R1047 B.n374 B.n373 6.5566
R1048 B.n361 B.n360 6.5566
R1049 B.n194 B.n193 6.5566
R1050 B.n206 B.n88 6.5566
R1051 B.n375 B.n374 4.05904
R1052 B.n360 B.n359 4.05904
R1053 B.n193 B.n192 4.05904
R1054 B.n209 B.n88 4.05904
R1055 B.n451 B.n0 2.81026
R1056 B.n451 B.n1 2.81026
C0 VDD2 VDD1 1.07994f
C1 VN VP 4.54882f
C2 VDD2 w_n2594_n1740# 1.54341f
C3 B VN 0.890188f
C4 VTAIL VP 2.64301f
C5 w_n2594_n1740# VDD1 1.48758f
C6 VTAIL B 1.57398f
C7 VDD2 VN 2.21548f
C8 VTAIL VDD2 4.37184f
C9 VDD1 VN 0.154008f
C10 w_n2594_n1740# VN 4.54589f
C11 B VP 1.44117f
C12 VTAIL VDD1 4.32559f
C13 VTAIL w_n2594_n1740# 1.70852f
C14 VDD2 VP 0.386203f
C15 B VDD2 1.27726f
C16 VDD1 VP 2.44551f
C17 VTAIL VN 2.62881f
C18 B VDD1 1.22458f
C19 w_n2594_n1740# VP 4.87767f
C20 B w_n2594_n1740# 6.16026f
C21 VDD2 VSUBS 1.118838f
C22 VDD1 VSUBS 1.172147f
C23 VTAIL VSUBS 0.480949f
C24 VN VSUBS 4.64369f
C25 VP VSUBS 1.756335f
C26 B VSUBS 2.899783f
C27 w_n2594_n1740# VSUBS 56.870895f
C28 B.n0 VSUBS 0.004592f
C29 B.n1 VSUBS 0.004592f
C30 B.n2 VSUBS 0.007262f
C31 B.n3 VSUBS 0.007262f
C32 B.n4 VSUBS 0.007262f
C33 B.n5 VSUBS 0.007262f
C34 B.n6 VSUBS 0.007262f
C35 B.n7 VSUBS 0.007262f
C36 B.n8 VSUBS 0.007262f
C37 B.n9 VSUBS 0.007262f
C38 B.n10 VSUBS 0.007262f
C39 B.n11 VSUBS 0.007262f
C40 B.n12 VSUBS 0.007262f
C41 B.n13 VSUBS 0.007262f
C42 B.n14 VSUBS 0.007262f
C43 B.n15 VSUBS 0.007262f
C44 B.n16 VSUBS 0.007262f
C45 B.n17 VSUBS 0.007262f
C46 B.n18 VSUBS 0.017206f
C47 B.n19 VSUBS 0.007262f
C48 B.n20 VSUBS 0.007262f
C49 B.n21 VSUBS 0.007262f
C50 B.n22 VSUBS 0.007262f
C51 B.n23 VSUBS 0.007262f
C52 B.n24 VSUBS 0.007262f
C53 B.n25 VSUBS 0.007262f
C54 B.n26 VSUBS 0.007262f
C55 B.n27 VSUBS 0.007262f
C56 B.t5 VSUBS 0.057748f
C57 B.t4 VSUBS 0.072627f
C58 B.t3 VSUBS 0.322309f
C59 B.n28 VSUBS 0.130708f
C60 B.n29 VSUBS 0.113262f
C61 B.n30 VSUBS 0.007262f
C62 B.n31 VSUBS 0.007262f
C63 B.n32 VSUBS 0.007262f
C64 B.n33 VSUBS 0.007262f
C65 B.t2 VSUBS 0.057749f
C66 B.t1 VSUBS 0.072627f
C67 B.t0 VSUBS 0.322309f
C68 B.n34 VSUBS 0.130708f
C69 B.n35 VSUBS 0.113261f
C70 B.n36 VSUBS 0.007262f
C71 B.n37 VSUBS 0.007262f
C72 B.n38 VSUBS 0.007262f
C73 B.n39 VSUBS 0.007262f
C74 B.n40 VSUBS 0.007262f
C75 B.n41 VSUBS 0.007262f
C76 B.n42 VSUBS 0.007262f
C77 B.n43 VSUBS 0.007262f
C78 B.n44 VSUBS 0.01633f
C79 B.n45 VSUBS 0.007262f
C80 B.n46 VSUBS 0.007262f
C81 B.n47 VSUBS 0.007262f
C82 B.n48 VSUBS 0.007262f
C83 B.n49 VSUBS 0.007262f
C84 B.n50 VSUBS 0.007262f
C85 B.n51 VSUBS 0.007262f
C86 B.n52 VSUBS 0.007262f
C87 B.n53 VSUBS 0.007262f
C88 B.n54 VSUBS 0.007262f
C89 B.n55 VSUBS 0.007262f
C90 B.n56 VSUBS 0.007262f
C91 B.n57 VSUBS 0.007262f
C92 B.n58 VSUBS 0.007262f
C93 B.n59 VSUBS 0.007262f
C94 B.n60 VSUBS 0.007262f
C95 B.n61 VSUBS 0.007262f
C96 B.n62 VSUBS 0.007262f
C97 B.n63 VSUBS 0.007262f
C98 B.n64 VSUBS 0.007262f
C99 B.n65 VSUBS 0.007262f
C100 B.n66 VSUBS 0.007262f
C101 B.n67 VSUBS 0.007262f
C102 B.n68 VSUBS 0.007262f
C103 B.n69 VSUBS 0.007262f
C104 B.n70 VSUBS 0.007262f
C105 B.n71 VSUBS 0.007262f
C106 B.n72 VSUBS 0.007262f
C107 B.n73 VSUBS 0.007262f
C108 B.n74 VSUBS 0.007262f
C109 B.n75 VSUBS 0.007262f
C110 B.n76 VSUBS 0.007262f
C111 B.n77 VSUBS 0.017206f
C112 B.n78 VSUBS 0.007262f
C113 B.n79 VSUBS 0.007262f
C114 B.n80 VSUBS 0.007262f
C115 B.n81 VSUBS 0.007262f
C116 B.n82 VSUBS 0.007262f
C117 B.n83 VSUBS 0.007262f
C118 B.n84 VSUBS 0.007262f
C119 B.n85 VSUBS 0.007262f
C120 B.t10 VSUBS 0.057749f
C121 B.t11 VSUBS 0.072627f
C122 B.t9 VSUBS 0.322309f
C123 B.n86 VSUBS 0.130708f
C124 B.n87 VSUBS 0.113261f
C125 B.n88 VSUBS 0.016826f
C126 B.n89 VSUBS 0.007262f
C127 B.n90 VSUBS 0.007262f
C128 B.n91 VSUBS 0.007262f
C129 B.n92 VSUBS 0.007262f
C130 B.n93 VSUBS 0.007262f
C131 B.t7 VSUBS 0.057748f
C132 B.t8 VSUBS 0.072627f
C133 B.t6 VSUBS 0.322309f
C134 B.n94 VSUBS 0.130708f
C135 B.n95 VSUBS 0.113262f
C136 B.n96 VSUBS 0.007262f
C137 B.n97 VSUBS 0.007262f
C138 B.n98 VSUBS 0.007262f
C139 B.n99 VSUBS 0.007262f
C140 B.n100 VSUBS 0.007262f
C141 B.n101 VSUBS 0.007262f
C142 B.n102 VSUBS 0.007262f
C143 B.n103 VSUBS 0.007262f
C144 B.n104 VSUBS 0.01633f
C145 B.n105 VSUBS 0.007262f
C146 B.n106 VSUBS 0.007262f
C147 B.n107 VSUBS 0.007262f
C148 B.n108 VSUBS 0.007262f
C149 B.n109 VSUBS 0.007262f
C150 B.n110 VSUBS 0.007262f
C151 B.n111 VSUBS 0.007262f
C152 B.n112 VSUBS 0.007262f
C153 B.n113 VSUBS 0.007262f
C154 B.n114 VSUBS 0.007262f
C155 B.n115 VSUBS 0.007262f
C156 B.n116 VSUBS 0.007262f
C157 B.n117 VSUBS 0.007262f
C158 B.n118 VSUBS 0.007262f
C159 B.n119 VSUBS 0.007262f
C160 B.n120 VSUBS 0.007262f
C161 B.n121 VSUBS 0.007262f
C162 B.n122 VSUBS 0.007262f
C163 B.n123 VSUBS 0.007262f
C164 B.n124 VSUBS 0.007262f
C165 B.n125 VSUBS 0.007262f
C166 B.n126 VSUBS 0.007262f
C167 B.n127 VSUBS 0.007262f
C168 B.n128 VSUBS 0.007262f
C169 B.n129 VSUBS 0.007262f
C170 B.n130 VSUBS 0.007262f
C171 B.n131 VSUBS 0.007262f
C172 B.n132 VSUBS 0.007262f
C173 B.n133 VSUBS 0.007262f
C174 B.n134 VSUBS 0.007262f
C175 B.n135 VSUBS 0.007262f
C176 B.n136 VSUBS 0.007262f
C177 B.n137 VSUBS 0.007262f
C178 B.n138 VSUBS 0.007262f
C179 B.n139 VSUBS 0.007262f
C180 B.n140 VSUBS 0.007262f
C181 B.n141 VSUBS 0.007262f
C182 B.n142 VSUBS 0.007262f
C183 B.n143 VSUBS 0.007262f
C184 B.n144 VSUBS 0.007262f
C185 B.n145 VSUBS 0.007262f
C186 B.n146 VSUBS 0.007262f
C187 B.n147 VSUBS 0.007262f
C188 B.n148 VSUBS 0.007262f
C189 B.n149 VSUBS 0.007262f
C190 B.n150 VSUBS 0.007262f
C191 B.n151 VSUBS 0.007262f
C192 B.n152 VSUBS 0.007262f
C193 B.n153 VSUBS 0.007262f
C194 B.n154 VSUBS 0.007262f
C195 B.n155 VSUBS 0.007262f
C196 B.n156 VSUBS 0.007262f
C197 B.n157 VSUBS 0.007262f
C198 B.n158 VSUBS 0.007262f
C199 B.n159 VSUBS 0.007262f
C200 B.n160 VSUBS 0.007262f
C201 B.n161 VSUBS 0.007262f
C202 B.n162 VSUBS 0.007262f
C203 B.n163 VSUBS 0.007262f
C204 B.n164 VSUBS 0.007262f
C205 B.n165 VSUBS 0.01633f
C206 B.n166 VSUBS 0.017206f
C207 B.n167 VSUBS 0.017206f
C208 B.n168 VSUBS 0.007262f
C209 B.n169 VSUBS 0.007262f
C210 B.n170 VSUBS 0.007262f
C211 B.n171 VSUBS 0.007262f
C212 B.n172 VSUBS 0.007262f
C213 B.n173 VSUBS 0.007262f
C214 B.n174 VSUBS 0.007262f
C215 B.n175 VSUBS 0.007262f
C216 B.n176 VSUBS 0.007262f
C217 B.n177 VSUBS 0.007262f
C218 B.n178 VSUBS 0.007262f
C219 B.n179 VSUBS 0.007262f
C220 B.n180 VSUBS 0.007262f
C221 B.n181 VSUBS 0.007262f
C222 B.n182 VSUBS 0.007262f
C223 B.n183 VSUBS 0.007262f
C224 B.n184 VSUBS 0.007262f
C225 B.n185 VSUBS 0.007262f
C226 B.n186 VSUBS 0.007262f
C227 B.n187 VSUBS 0.007262f
C228 B.n188 VSUBS 0.007262f
C229 B.n189 VSUBS 0.007262f
C230 B.n190 VSUBS 0.007262f
C231 B.n191 VSUBS 0.007262f
C232 B.n192 VSUBS 0.00502f
C233 B.n193 VSUBS 0.016826f
C234 B.n194 VSUBS 0.005874f
C235 B.n195 VSUBS 0.007262f
C236 B.n196 VSUBS 0.007262f
C237 B.n197 VSUBS 0.007262f
C238 B.n198 VSUBS 0.007262f
C239 B.n199 VSUBS 0.007262f
C240 B.n200 VSUBS 0.007262f
C241 B.n201 VSUBS 0.007262f
C242 B.n202 VSUBS 0.007262f
C243 B.n203 VSUBS 0.007262f
C244 B.n204 VSUBS 0.007262f
C245 B.n205 VSUBS 0.007262f
C246 B.n206 VSUBS 0.005874f
C247 B.n207 VSUBS 0.007262f
C248 B.n208 VSUBS 0.007262f
C249 B.n209 VSUBS 0.00502f
C250 B.n210 VSUBS 0.007262f
C251 B.n211 VSUBS 0.007262f
C252 B.n212 VSUBS 0.007262f
C253 B.n213 VSUBS 0.007262f
C254 B.n214 VSUBS 0.007262f
C255 B.n215 VSUBS 0.007262f
C256 B.n216 VSUBS 0.007262f
C257 B.n217 VSUBS 0.007262f
C258 B.n218 VSUBS 0.007262f
C259 B.n219 VSUBS 0.007262f
C260 B.n220 VSUBS 0.007262f
C261 B.n221 VSUBS 0.007262f
C262 B.n222 VSUBS 0.007262f
C263 B.n223 VSUBS 0.007262f
C264 B.n224 VSUBS 0.007262f
C265 B.n225 VSUBS 0.007262f
C266 B.n226 VSUBS 0.007262f
C267 B.n227 VSUBS 0.007262f
C268 B.n228 VSUBS 0.007262f
C269 B.n229 VSUBS 0.007262f
C270 B.n230 VSUBS 0.007262f
C271 B.n231 VSUBS 0.007262f
C272 B.n232 VSUBS 0.007262f
C273 B.n233 VSUBS 0.007262f
C274 B.n234 VSUBS 0.017206f
C275 B.n235 VSUBS 0.01633f
C276 B.n236 VSUBS 0.01633f
C277 B.n237 VSUBS 0.007262f
C278 B.n238 VSUBS 0.007262f
C279 B.n239 VSUBS 0.007262f
C280 B.n240 VSUBS 0.007262f
C281 B.n241 VSUBS 0.007262f
C282 B.n242 VSUBS 0.007262f
C283 B.n243 VSUBS 0.007262f
C284 B.n244 VSUBS 0.007262f
C285 B.n245 VSUBS 0.007262f
C286 B.n246 VSUBS 0.007262f
C287 B.n247 VSUBS 0.007262f
C288 B.n248 VSUBS 0.007262f
C289 B.n249 VSUBS 0.007262f
C290 B.n250 VSUBS 0.007262f
C291 B.n251 VSUBS 0.007262f
C292 B.n252 VSUBS 0.007262f
C293 B.n253 VSUBS 0.007262f
C294 B.n254 VSUBS 0.007262f
C295 B.n255 VSUBS 0.007262f
C296 B.n256 VSUBS 0.007262f
C297 B.n257 VSUBS 0.007262f
C298 B.n258 VSUBS 0.007262f
C299 B.n259 VSUBS 0.007262f
C300 B.n260 VSUBS 0.007262f
C301 B.n261 VSUBS 0.007262f
C302 B.n262 VSUBS 0.007262f
C303 B.n263 VSUBS 0.007262f
C304 B.n264 VSUBS 0.007262f
C305 B.n265 VSUBS 0.007262f
C306 B.n266 VSUBS 0.007262f
C307 B.n267 VSUBS 0.007262f
C308 B.n268 VSUBS 0.007262f
C309 B.n269 VSUBS 0.007262f
C310 B.n270 VSUBS 0.007262f
C311 B.n271 VSUBS 0.007262f
C312 B.n272 VSUBS 0.007262f
C313 B.n273 VSUBS 0.007262f
C314 B.n274 VSUBS 0.007262f
C315 B.n275 VSUBS 0.007262f
C316 B.n276 VSUBS 0.007262f
C317 B.n277 VSUBS 0.007262f
C318 B.n278 VSUBS 0.007262f
C319 B.n279 VSUBS 0.007262f
C320 B.n280 VSUBS 0.007262f
C321 B.n281 VSUBS 0.007262f
C322 B.n282 VSUBS 0.007262f
C323 B.n283 VSUBS 0.007262f
C324 B.n284 VSUBS 0.007262f
C325 B.n285 VSUBS 0.007262f
C326 B.n286 VSUBS 0.007262f
C327 B.n287 VSUBS 0.007262f
C328 B.n288 VSUBS 0.007262f
C329 B.n289 VSUBS 0.007262f
C330 B.n290 VSUBS 0.007262f
C331 B.n291 VSUBS 0.007262f
C332 B.n292 VSUBS 0.007262f
C333 B.n293 VSUBS 0.007262f
C334 B.n294 VSUBS 0.007262f
C335 B.n295 VSUBS 0.007262f
C336 B.n296 VSUBS 0.007262f
C337 B.n297 VSUBS 0.007262f
C338 B.n298 VSUBS 0.007262f
C339 B.n299 VSUBS 0.007262f
C340 B.n300 VSUBS 0.007262f
C341 B.n301 VSUBS 0.007262f
C342 B.n302 VSUBS 0.007262f
C343 B.n303 VSUBS 0.007262f
C344 B.n304 VSUBS 0.007262f
C345 B.n305 VSUBS 0.007262f
C346 B.n306 VSUBS 0.007262f
C347 B.n307 VSUBS 0.007262f
C348 B.n308 VSUBS 0.007262f
C349 B.n309 VSUBS 0.007262f
C350 B.n310 VSUBS 0.007262f
C351 B.n311 VSUBS 0.007262f
C352 B.n312 VSUBS 0.007262f
C353 B.n313 VSUBS 0.007262f
C354 B.n314 VSUBS 0.007262f
C355 B.n315 VSUBS 0.007262f
C356 B.n316 VSUBS 0.007262f
C357 B.n317 VSUBS 0.007262f
C358 B.n318 VSUBS 0.007262f
C359 B.n319 VSUBS 0.007262f
C360 B.n320 VSUBS 0.007262f
C361 B.n321 VSUBS 0.007262f
C362 B.n322 VSUBS 0.007262f
C363 B.n323 VSUBS 0.007262f
C364 B.n324 VSUBS 0.007262f
C365 B.n325 VSUBS 0.007262f
C366 B.n326 VSUBS 0.007262f
C367 B.n327 VSUBS 0.007262f
C368 B.n328 VSUBS 0.007262f
C369 B.n329 VSUBS 0.007262f
C370 B.n330 VSUBS 0.007262f
C371 B.n331 VSUBS 0.017206f
C372 B.n332 VSUBS 0.01633f
C373 B.n333 VSUBS 0.017206f
C374 B.n334 VSUBS 0.007262f
C375 B.n335 VSUBS 0.007262f
C376 B.n336 VSUBS 0.007262f
C377 B.n337 VSUBS 0.007262f
C378 B.n338 VSUBS 0.007262f
C379 B.n339 VSUBS 0.007262f
C380 B.n340 VSUBS 0.007262f
C381 B.n341 VSUBS 0.007262f
C382 B.n342 VSUBS 0.007262f
C383 B.n343 VSUBS 0.007262f
C384 B.n344 VSUBS 0.007262f
C385 B.n345 VSUBS 0.007262f
C386 B.n346 VSUBS 0.007262f
C387 B.n347 VSUBS 0.007262f
C388 B.n348 VSUBS 0.007262f
C389 B.n349 VSUBS 0.007262f
C390 B.n350 VSUBS 0.007262f
C391 B.n351 VSUBS 0.007262f
C392 B.n352 VSUBS 0.007262f
C393 B.n353 VSUBS 0.007262f
C394 B.n354 VSUBS 0.007262f
C395 B.n355 VSUBS 0.007262f
C396 B.n356 VSUBS 0.007262f
C397 B.n357 VSUBS 0.007262f
C398 B.n358 VSUBS 0.007262f
C399 B.n359 VSUBS 0.00502f
C400 B.n360 VSUBS 0.016826f
C401 B.n361 VSUBS 0.005874f
C402 B.n362 VSUBS 0.007262f
C403 B.n363 VSUBS 0.007262f
C404 B.n364 VSUBS 0.007262f
C405 B.n365 VSUBS 0.007262f
C406 B.n366 VSUBS 0.007262f
C407 B.n367 VSUBS 0.007262f
C408 B.n368 VSUBS 0.007262f
C409 B.n369 VSUBS 0.007262f
C410 B.n370 VSUBS 0.007262f
C411 B.n371 VSUBS 0.007262f
C412 B.n372 VSUBS 0.007262f
C413 B.n373 VSUBS 0.005874f
C414 B.n374 VSUBS 0.016826f
C415 B.n375 VSUBS 0.00502f
C416 B.n376 VSUBS 0.007262f
C417 B.n377 VSUBS 0.007262f
C418 B.n378 VSUBS 0.007262f
C419 B.n379 VSUBS 0.007262f
C420 B.n380 VSUBS 0.007262f
C421 B.n381 VSUBS 0.007262f
C422 B.n382 VSUBS 0.007262f
C423 B.n383 VSUBS 0.007262f
C424 B.n384 VSUBS 0.007262f
C425 B.n385 VSUBS 0.007262f
C426 B.n386 VSUBS 0.007262f
C427 B.n387 VSUBS 0.007262f
C428 B.n388 VSUBS 0.007262f
C429 B.n389 VSUBS 0.007262f
C430 B.n390 VSUBS 0.007262f
C431 B.n391 VSUBS 0.007262f
C432 B.n392 VSUBS 0.007262f
C433 B.n393 VSUBS 0.007262f
C434 B.n394 VSUBS 0.007262f
C435 B.n395 VSUBS 0.007262f
C436 B.n396 VSUBS 0.007262f
C437 B.n397 VSUBS 0.007262f
C438 B.n398 VSUBS 0.007262f
C439 B.n399 VSUBS 0.007262f
C440 B.n400 VSUBS 0.007262f
C441 B.n401 VSUBS 0.017206f
C442 B.n402 VSUBS 0.01633f
C443 B.n403 VSUBS 0.01633f
C444 B.n404 VSUBS 0.007262f
C445 B.n405 VSUBS 0.007262f
C446 B.n406 VSUBS 0.007262f
C447 B.n407 VSUBS 0.007262f
C448 B.n408 VSUBS 0.007262f
C449 B.n409 VSUBS 0.007262f
C450 B.n410 VSUBS 0.007262f
C451 B.n411 VSUBS 0.007262f
C452 B.n412 VSUBS 0.007262f
C453 B.n413 VSUBS 0.007262f
C454 B.n414 VSUBS 0.007262f
C455 B.n415 VSUBS 0.007262f
C456 B.n416 VSUBS 0.007262f
C457 B.n417 VSUBS 0.007262f
C458 B.n418 VSUBS 0.007262f
C459 B.n419 VSUBS 0.007262f
C460 B.n420 VSUBS 0.007262f
C461 B.n421 VSUBS 0.007262f
C462 B.n422 VSUBS 0.007262f
C463 B.n423 VSUBS 0.007262f
C464 B.n424 VSUBS 0.007262f
C465 B.n425 VSUBS 0.007262f
C466 B.n426 VSUBS 0.007262f
C467 B.n427 VSUBS 0.007262f
C468 B.n428 VSUBS 0.007262f
C469 B.n429 VSUBS 0.007262f
C470 B.n430 VSUBS 0.007262f
C471 B.n431 VSUBS 0.007262f
C472 B.n432 VSUBS 0.007262f
C473 B.n433 VSUBS 0.007262f
C474 B.n434 VSUBS 0.007262f
C475 B.n435 VSUBS 0.007262f
C476 B.n436 VSUBS 0.007262f
C477 B.n437 VSUBS 0.007262f
C478 B.n438 VSUBS 0.007262f
C479 B.n439 VSUBS 0.007262f
C480 B.n440 VSUBS 0.007262f
C481 B.n441 VSUBS 0.007262f
C482 B.n442 VSUBS 0.007262f
C483 B.n443 VSUBS 0.007262f
C484 B.n444 VSUBS 0.007262f
C485 B.n445 VSUBS 0.007262f
C486 B.n446 VSUBS 0.007262f
C487 B.n447 VSUBS 0.007262f
C488 B.n448 VSUBS 0.007262f
C489 B.n449 VSUBS 0.007262f
C490 B.n450 VSUBS 0.007262f
C491 B.n451 VSUBS 0.016445f
C492 VDD2.n0 VSUBS 0.023468f
C493 VDD2.n1 VSUBS 0.022303f
C494 VDD2.n2 VSUBS 0.011985f
C495 VDD2.n3 VSUBS 0.028327f
C496 VDD2.n4 VSUBS 0.01269f
C497 VDD2.n5 VSUBS 0.08538f
C498 VDD2.t3 VSUBS 0.062148f
C499 VDD2.n6 VSUBS 0.021246f
C500 VDD2.n7 VSUBS 0.017818f
C501 VDD2.n8 VSUBS 0.011985f
C502 VDD2.n9 VSUBS 0.292808f
C503 VDD2.n10 VSUBS 0.022303f
C504 VDD2.n11 VSUBS 0.011985f
C505 VDD2.n12 VSUBS 0.01269f
C506 VDD2.n13 VSUBS 0.028327f
C507 VDD2.n14 VSUBS 0.06504f
C508 VDD2.n15 VSUBS 0.01269f
C509 VDD2.n16 VSUBS 0.011985f
C510 VDD2.n17 VSUBS 0.052162f
C511 VDD2.n18 VSUBS 0.051301f
C512 VDD2.t5 VSUBS 0.068031f
C513 VDD2.t0 VSUBS 0.068031f
C514 VDD2.n19 VSUBS 0.394489f
C515 VDD2.n20 VSUBS 1.73767f
C516 VDD2.n21 VSUBS 0.023468f
C517 VDD2.n22 VSUBS 0.022303f
C518 VDD2.n23 VSUBS 0.011985f
C519 VDD2.n24 VSUBS 0.028327f
C520 VDD2.n25 VSUBS 0.01269f
C521 VDD2.n26 VSUBS 0.08538f
C522 VDD2.t4 VSUBS 0.062148f
C523 VDD2.n27 VSUBS 0.021246f
C524 VDD2.n28 VSUBS 0.017818f
C525 VDD2.n29 VSUBS 0.011985f
C526 VDD2.n30 VSUBS 0.292808f
C527 VDD2.n31 VSUBS 0.022303f
C528 VDD2.n32 VSUBS 0.011985f
C529 VDD2.n33 VSUBS 0.01269f
C530 VDD2.n34 VSUBS 0.028327f
C531 VDD2.n35 VSUBS 0.06504f
C532 VDD2.n36 VSUBS 0.01269f
C533 VDD2.n37 VSUBS 0.011985f
C534 VDD2.n38 VSUBS 0.052162f
C535 VDD2.n39 VSUBS 0.047965f
C536 VDD2.n40 VSUBS 1.48993f
C537 VDD2.t2 VSUBS 0.068031f
C538 VDD2.t1 VSUBS 0.068031f
C539 VDD2.n41 VSUBS 0.394472f
C540 VN.n0 VSUBS 0.050758f
C541 VN.t5 VSUBS 0.852826f
C542 VN.n1 VSUBS 0.041141f
C543 VN.t2 VSUBS 1.07429f
C544 VN.n2 VSUBS 0.453961f
C545 VN.t0 VSUBS 0.852826f
C546 VN.n3 VSUBS 0.490662f
C547 VN.n4 VSUBS 0.10103f
C548 VN.n5 VSUBS 0.367881f
C549 VN.n6 VSUBS 0.050758f
C550 VN.n7 VSUBS 0.050758f
C551 VN.n8 VSUBS 0.099525f
C552 VN.n9 VSUBS 0.050447f
C553 VN.n10 VSUBS 0.458636f
C554 VN.n11 VSUBS 0.053814f
C555 VN.n12 VSUBS 0.050758f
C556 VN.t1 VSUBS 0.852826f
C557 VN.n13 VSUBS 0.041141f
C558 VN.t4 VSUBS 1.07429f
C559 VN.n14 VSUBS 0.453961f
C560 VN.t3 VSUBS 0.852826f
C561 VN.n15 VSUBS 0.490662f
C562 VN.n16 VSUBS 0.10103f
C563 VN.n17 VSUBS 0.367881f
C564 VN.n18 VSUBS 0.050758f
C565 VN.n19 VSUBS 0.050758f
C566 VN.n20 VSUBS 0.099525f
C567 VN.n21 VSUBS 0.050447f
C568 VN.n22 VSUBS 0.458636f
C569 VN.n23 VSUBS 1.87874f
C570 VDD1.n0 VSUBS 0.023529f
C571 VDD1.n1 VSUBS 0.022362f
C572 VDD1.n2 VSUBS 0.012016f
C573 VDD1.n3 VSUBS 0.028402f
C574 VDD1.n4 VSUBS 0.012723f
C575 VDD1.n5 VSUBS 0.085605f
C576 VDD1.t2 VSUBS 0.062312f
C577 VDD1.n6 VSUBS 0.021302f
C578 VDD1.n7 VSUBS 0.017865f
C579 VDD1.n8 VSUBS 0.012016f
C580 VDD1.n9 VSUBS 0.293581f
C581 VDD1.n10 VSUBS 0.022362f
C582 VDD1.n11 VSUBS 0.012016f
C583 VDD1.n12 VSUBS 0.012723f
C584 VDD1.n13 VSUBS 0.028402f
C585 VDD1.n14 VSUBS 0.065211f
C586 VDD1.n15 VSUBS 0.012723f
C587 VDD1.n16 VSUBS 0.012016f
C588 VDD1.n17 VSUBS 0.052299f
C589 VDD1.n18 VSUBS 0.051941f
C590 VDD1.n19 VSUBS 0.023529f
C591 VDD1.n20 VSUBS 0.022362f
C592 VDD1.n21 VSUBS 0.012016f
C593 VDD1.n22 VSUBS 0.028402f
C594 VDD1.n23 VSUBS 0.012723f
C595 VDD1.n24 VSUBS 0.085605f
C596 VDD1.t1 VSUBS 0.062312f
C597 VDD1.n25 VSUBS 0.021302f
C598 VDD1.n26 VSUBS 0.017865f
C599 VDD1.n27 VSUBS 0.012016f
C600 VDD1.n28 VSUBS 0.293581f
C601 VDD1.n29 VSUBS 0.022362f
C602 VDD1.n30 VSUBS 0.012016f
C603 VDD1.n31 VSUBS 0.012723f
C604 VDD1.n32 VSUBS 0.028402f
C605 VDD1.n33 VSUBS 0.065211f
C606 VDD1.n34 VSUBS 0.012723f
C607 VDD1.n35 VSUBS 0.012016f
C608 VDD1.n36 VSUBS 0.052299f
C609 VDD1.n37 VSUBS 0.051436f
C610 VDD1.t0 VSUBS 0.06821f
C611 VDD1.t4 VSUBS 0.06821f
C612 VDD1.n38 VSUBS 0.395529f
C613 VDD1.n39 VSUBS 1.82698f
C614 VDD1.t3 VSUBS 0.06821f
C615 VDD1.t5 VSUBS 0.06821f
C616 VDD1.n40 VSUBS 0.393938f
C617 VDD1.n41 VSUBS 1.82398f
C618 VTAIL.t1 VSUBS 0.086027f
C619 VTAIL.t3 VSUBS 0.086027f
C620 VTAIL.n0 VSUBS 0.430292f
C621 VTAIL.n1 VSUBS 0.588962f
C622 VTAIL.n2 VSUBS 0.029676f
C623 VTAIL.n3 VSUBS 0.028203f
C624 VTAIL.n4 VSUBS 0.015155f
C625 VTAIL.n5 VSUBS 0.035821f
C626 VTAIL.n6 VSUBS 0.016047f
C627 VTAIL.n7 VSUBS 0.107966f
C628 VTAIL.t7 VSUBS 0.078588f
C629 VTAIL.n8 VSUBS 0.026866f
C630 VTAIL.n9 VSUBS 0.022531f
C631 VTAIL.n10 VSUBS 0.015155f
C632 VTAIL.n11 VSUBS 0.370267f
C633 VTAIL.n12 VSUBS 0.028203f
C634 VTAIL.n13 VSUBS 0.015155f
C635 VTAIL.n14 VSUBS 0.016047f
C636 VTAIL.n15 VSUBS 0.035821f
C637 VTAIL.n16 VSUBS 0.082245f
C638 VTAIL.n17 VSUBS 0.016047f
C639 VTAIL.n18 VSUBS 0.015155f
C640 VTAIL.n19 VSUBS 0.065961f
C641 VTAIL.n20 VSUBS 0.041185f
C642 VTAIL.n21 VSUBS 0.30577f
C643 VTAIL.t6 VSUBS 0.086027f
C644 VTAIL.t11 VSUBS 0.086027f
C645 VTAIL.n22 VSUBS 0.430292f
C646 VTAIL.n23 VSUBS 1.58431f
C647 VTAIL.t0 VSUBS 0.086027f
C648 VTAIL.t4 VSUBS 0.086027f
C649 VTAIL.n24 VSUBS 0.430295f
C650 VTAIL.n25 VSUBS 1.58431f
C651 VTAIL.n26 VSUBS 0.029676f
C652 VTAIL.n27 VSUBS 0.028203f
C653 VTAIL.n28 VSUBS 0.015155f
C654 VTAIL.n29 VSUBS 0.035821f
C655 VTAIL.n30 VSUBS 0.016047f
C656 VTAIL.n31 VSUBS 0.107966f
C657 VTAIL.t5 VSUBS 0.078588f
C658 VTAIL.n32 VSUBS 0.026866f
C659 VTAIL.n33 VSUBS 0.022531f
C660 VTAIL.n34 VSUBS 0.015155f
C661 VTAIL.n35 VSUBS 0.370267f
C662 VTAIL.n36 VSUBS 0.028203f
C663 VTAIL.n37 VSUBS 0.015155f
C664 VTAIL.n38 VSUBS 0.016047f
C665 VTAIL.n39 VSUBS 0.035821f
C666 VTAIL.n40 VSUBS 0.082245f
C667 VTAIL.n41 VSUBS 0.016047f
C668 VTAIL.n42 VSUBS 0.015155f
C669 VTAIL.n43 VSUBS 0.065961f
C670 VTAIL.n44 VSUBS 0.041185f
C671 VTAIL.n45 VSUBS 0.30577f
C672 VTAIL.t10 VSUBS 0.086027f
C673 VTAIL.t8 VSUBS 0.086027f
C674 VTAIL.n46 VSUBS 0.430295f
C675 VTAIL.n47 VSUBS 0.702946f
C676 VTAIL.n48 VSUBS 0.029676f
C677 VTAIL.n49 VSUBS 0.028203f
C678 VTAIL.n50 VSUBS 0.015155f
C679 VTAIL.n51 VSUBS 0.035821f
C680 VTAIL.n52 VSUBS 0.016047f
C681 VTAIL.n53 VSUBS 0.107966f
C682 VTAIL.t9 VSUBS 0.078588f
C683 VTAIL.n54 VSUBS 0.026866f
C684 VTAIL.n55 VSUBS 0.022531f
C685 VTAIL.n56 VSUBS 0.015155f
C686 VTAIL.n57 VSUBS 0.370267f
C687 VTAIL.n58 VSUBS 0.028203f
C688 VTAIL.n59 VSUBS 0.015155f
C689 VTAIL.n60 VSUBS 0.016047f
C690 VTAIL.n61 VSUBS 0.035821f
C691 VTAIL.n62 VSUBS 0.082245f
C692 VTAIL.n63 VSUBS 0.016047f
C693 VTAIL.n64 VSUBS 0.015155f
C694 VTAIL.n65 VSUBS 0.065961f
C695 VTAIL.n66 VSUBS 0.041185f
C696 VTAIL.n67 VSUBS 1.02809f
C697 VTAIL.n68 VSUBS 0.029676f
C698 VTAIL.n69 VSUBS 0.028203f
C699 VTAIL.n70 VSUBS 0.015155f
C700 VTAIL.n71 VSUBS 0.035821f
C701 VTAIL.n72 VSUBS 0.016047f
C702 VTAIL.n73 VSUBS 0.107966f
C703 VTAIL.t2 VSUBS 0.078588f
C704 VTAIL.n74 VSUBS 0.026866f
C705 VTAIL.n75 VSUBS 0.022531f
C706 VTAIL.n76 VSUBS 0.015155f
C707 VTAIL.n77 VSUBS 0.370267f
C708 VTAIL.n78 VSUBS 0.028203f
C709 VTAIL.n79 VSUBS 0.015155f
C710 VTAIL.n80 VSUBS 0.016047f
C711 VTAIL.n81 VSUBS 0.035821f
C712 VTAIL.n82 VSUBS 0.082245f
C713 VTAIL.n83 VSUBS 0.016047f
C714 VTAIL.n84 VSUBS 0.015155f
C715 VTAIL.n85 VSUBS 0.065961f
C716 VTAIL.n86 VSUBS 0.041185f
C717 VTAIL.n87 VSUBS 0.983048f
C718 VP.n0 VSUBS 0.05324f
C719 VP.t1 VSUBS 0.89453f
C720 VP.n1 VSUBS 0.043153f
C721 VP.n2 VSUBS 0.05324f
C722 VP.t5 VSUBS 0.89453f
C723 VP.n3 VSUBS 0.043153f
C724 VP.n4 VSUBS 0.05324f
C725 VP.t4 VSUBS 0.89453f
C726 VP.n5 VSUBS 0.05324f
C727 VP.t0 VSUBS 0.89453f
C728 VP.n6 VSUBS 0.043153f
C729 VP.t3 VSUBS 1.12683f
C730 VP.n7 VSUBS 0.476161f
C731 VP.t2 VSUBS 0.89453f
C732 VP.n8 VSUBS 0.514657f
C733 VP.n9 VSUBS 0.105971f
C734 VP.n10 VSUBS 0.385871f
C735 VP.n11 VSUBS 0.05324f
C736 VP.n12 VSUBS 0.05324f
C737 VP.n13 VSUBS 0.104392f
C738 VP.n14 VSUBS 0.052914f
C739 VP.n15 VSUBS 0.481064f
C740 VP.n16 VSUBS 1.93549f
C741 VP.n17 VSUBS 1.98493f
C742 VP.n18 VSUBS 0.481064f
C743 VP.n19 VSUBS 0.052914f
C744 VP.n20 VSUBS 0.104392f
C745 VP.n21 VSUBS 0.05324f
C746 VP.n22 VSUBS 0.05324f
C747 VP.n23 VSUBS 0.05324f
C748 VP.n24 VSUBS 0.105971f
C749 VP.n25 VSUBS 0.425089f
C750 VP.n26 VSUBS 0.105971f
C751 VP.n27 VSUBS 0.05324f
C752 VP.n28 VSUBS 0.05324f
C753 VP.n29 VSUBS 0.05324f
C754 VP.n30 VSUBS 0.104392f
C755 VP.n31 VSUBS 0.052914f
C756 VP.n32 VSUBS 0.481064f
C757 VP.n33 VSUBS 0.056445f
.ends

