* NGSPICE file created from diff_pair_sample_0889.ext - technology: sky130A

.subckt diff_pair_sample_0889 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=2.8509 pd=15.4 as=0 ps=0 w=7.31 l=3.53
X1 VDD1.t3 VP.t0 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.20615 pd=7.64 as=2.8509 ps=15.4 w=7.31 l=3.53
X2 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=2.8509 pd=15.4 as=0 ps=0 w=7.31 l=3.53
X3 VTAIL.t3 VN.t0 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.8509 pd=15.4 as=1.20615 ps=7.64 w=7.31 l=3.53
X4 VTAIL.t0 VN.t1 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.8509 pd=15.4 as=1.20615 ps=7.64 w=7.31 l=3.53
X5 VTAIL.t7 VP.t1 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.8509 pd=15.4 as=1.20615 ps=7.64 w=7.31 l=3.53
X6 VDD1.t1 VP.t2 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=1.20615 pd=7.64 as=2.8509 ps=15.4 w=7.31 l=3.53
X7 VDD2.t1 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.20615 pd=7.64 as=2.8509 ps=15.4 w=7.31 l=3.53
X8 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.8509 pd=15.4 as=0 ps=0 w=7.31 l=3.53
X9 VDD2.t0 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.20615 pd=7.64 as=2.8509 ps=15.4 w=7.31 l=3.53
X10 VTAIL.t4 VP.t3 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=2.8509 pd=15.4 as=1.20615 ps=7.64 w=7.31 l=3.53
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.8509 pd=15.4 as=0 ps=0 w=7.31 l=3.53
R0 B.n545 B.n115 585
R1 B.n115 B.n78 585
R2 B.n547 B.n546 585
R3 B.n549 B.n114 585
R4 B.n552 B.n551 585
R5 B.n553 B.n113 585
R6 B.n555 B.n554 585
R7 B.n557 B.n112 585
R8 B.n560 B.n559 585
R9 B.n561 B.n111 585
R10 B.n563 B.n562 585
R11 B.n565 B.n110 585
R12 B.n568 B.n567 585
R13 B.n569 B.n109 585
R14 B.n571 B.n570 585
R15 B.n573 B.n108 585
R16 B.n576 B.n575 585
R17 B.n577 B.n107 585
R18 B.n579 B.n578 585
R19 B.n581 B.n106 585
R20 B.n584 B.n583 585
R21 B.n585 B.n105 585
R22 B.n587 B.n586 585
R23 B.n589 B.n104 585
R24 B.n592 B.n591 585
R25 B.n593 B.n103 585
R26 B.n595 B.n594 585
R27 B.n597 B.n102 585
R28 B.n600 B.n599 585
R29 B.n602 B.n99 585
R30 B.n604 B.n603 585
R31 B.n606 B.n98 585
R32 B.n609 B.n608 585
R33 B.n610 B.n97 585
R34 B.n612 B.n611 585
R35 B.n614 B.n96 585
R36 B.n617 B.n616 585
R37 B.n618 B.n93 585
R38 B.n621 B.n620 585
R39 B.n623 B.n92 585
R40 B.n626 B.n625 585
R41 B.n627 B.n91 585
R42 B.n629 B.n628 585
R43 B.n631 B.n90 585
R44 B.n634 B.n633 585
R45 B.n635 B.n89 585
R46 B.n637 B.n636 585
R47 B.n639 B.n88 585
R48 B.n642 B.n641 585
R49 B.n643 B.n87 585
R50 B.n645 B.n644 585
R51 B.n647 B.n86 585
R52 B.n650 B.n649 585
R53 B.n651 B.n85 585
R54 B.n653 B.n652 585
R55 B.n655 B.n84 585
R56 B.n658 B.n657 585
R57 B.n659 B.n83 585
R58 B.n661 B.n660 585
R59 B.n663 B.n82 585
R60 B.n666 B.n665 585
R61 B.n667 B.n81 585
R62 B.n669 B.n668 585
R63 B.n671 B.n80 585
R64 B.n674 B.n673 585
R65 B.n675 B.n79 585
R66 B.n544 B.n77 585
R67 B.n678 B.n77 585
R68 B.n543 B.n76 585
R69 B.n679 B.n76 585
R70 B.n542 B.n75 585
R71 B.n680 B.n75 585
R72 B.n541 B.n540 585
R73 B.n540 B.n71 585
R74 B.n539 B.n70 585
R75 B.n686 B.n70 585
R76 B.n538 B.n69 585
R77 B.n687 B.n69 585
R78 B.n537 B.n68 585
R79 B.n688 B.n68 585
R80 B.n536 B.n535 585
R81 B.n535 B.n64 585
R82 B.n534 B.n63 585
R83 B.n694 B.n63 585
R84 B.n533 B.n62 585
R85 B.n695 B.n62 585
R86 B.n532 B.n61 585
R87 B.n696 B.n61 585
R88 B.n531 B.n530 585
R89 B.n530 B.n57 585
R90 B.n529 B.n56 585
R91 B.n702 B.n56 585
R92 B.n528 B.n55 585
R93 B.n703 B.n55 585
R94 B.n527 B.n54 585
R95 B.n704 B.n54 585
R96 B.n526 B.n525 585
R97 B.n525 B.n50 585
R98 B.n524 B.n49 585
R99 B.n710 B.n49 585
R100 B.n523 B.n48 585
R101 B.n711 B.n48 585
R102 B.n522 B.n47 585
R103 B.n712 B.n47 585
R104 B.n521 B.n520 585
R105 B.n520 B.n43 585
R106 B.n519 B.n42 585
R107 B.n718 B.n42 585
R108 B.n518 B.n41 585
R109 B.n719 B.n41 585
R110 B.n517 B.n40 585
R111 B.n720 B.n40 585
R112 B.n516 B.n515 585
R113 B.n515 B.n39 585
R114 B.n514 B.n35 585
R115 B.n726 B.n35 585
R116 B.n513 B.n34 585
R117 B.n727 B.n34 585
R118 B.n512 B.n33 585
R119 B.n728 B.n33 585
R120 B.n511 B.n510 585
R121 B.n510 B.n29 585
R122 B.n509 B.n28 585
R123 B.n734 B.n28 585
R124 B.n508 B.n27 585
R125 B.n735 B.n27 585
R126 B.n507 B.n26 585
R127 B.n736 B.n26 585
R128 B.n506 B.n505 585
R129 B.n505 B.n22 585
R130 B.n504 B.n21 585
R131 B.n742 B.n21 585
R132 B.n503 B.n20 585
R133 B.n743 B.n20 585
R134 B.n502 B.n19 585
R135 B.n744 B.n19 585
R136 B.n501 B.n500 585
R137 B.n500 B.n15 585
R138 B.n499 B.n14 585
R139 B.n750 B.n14 585
R140 B.n498 B.n13 585
R141 B.n751 B.n13 585
R142 B.n497 B.n12 585
R143 B.n752 B.n12 585
R144 B.n496 B.n495 585
R145 B.n495 B.n8 585
R146 B.n494 B.n7 585
R147 B.n758 B.n7 585
R148 B.n493 B.n6 585
R149 B.n759 B.n6 585
R150 B.n492 B.n5 585
R151 B.n760 B.n5 585
R152 B.n491 B.n490 585
R153 B.n490 B.n4 585
R154 B.n489 B.n116 585
R155 B.n489 B.n488 585
R156 B.n479 B.n117 585
R157 B.n118 B.n117 585
R158 B.n481 B.n480 585
R159 B.n482 B.n481 585
R160 B.n478 B.n123 585
R161 B.n123 B.n122 585
R162 B.n477 B.n476 585
R163 B.n476 B.n475 585
R164 B.n125 B.n124 585
R165 B.n126 B.n125 585
R166 B.n468 B.n467 585
R167 B.n469 B.n468 585
R168 B.n466 B.n131 585
R169 B.n131 B.n130 585
R170 B.n465 B.n464 585
R171 B.n464 B.n463 585
R172 B.n133 B.n132 585
R173 B.n134 B.n133 585
R174 B.n456 B.n455 585
R175 B.n457 B.n456 585
R176 B.n454 B.n139 585
R177 B.n139 B.n138 585
R178 B.n453 B.n452 585
R179 B.n452 B.n451 585
R180 B.n141 B.n140 585
R181 B.n142 B.n141 585
R182 B.n444 B.n443 585
R183 B.n445 B.n444 585
R184 B.n442 B.n147 585
R185 B.n147 B.n146 585
R186 B.n441 B.n440 585
R187 B.n440 B.n439 585
R188 B.n149 B.n148 585
R189 B.n432 B.n149 585
R190 B.n431 B.n430 585
R191 B.n433 B.n431 585
R192 B.n429 B.n154 585
R193 B.n154 B.n153 585
R194 B.n428 B.n427 585
R195 B.n427 B.n426 585
R196 B.n156 B.n155 585
R197 B.n157 B.n156 585
R198 B.n419 B.n418 585
R199 B.n420 B.n419 585
R200 B.n417 B.n162 585
R201 B.n162 B.n161 585
R202 B.n416 B.n415 585
R203 B.n415 B.n414 585
R204 B.n164 B.n163 585
R205 B.n165 B.n164 585
R206 B.n407 B.n406 585
R207 B.n408 B.n407 585
R208 B.n405 B.n170 585
R209 B.n170 B.n169 585
R210 B.n404 B.n403 585
R211 B.n403 B.n402 585
R212 B.n172 B.n171 585
R213 B.n173 B.n172 585
R214 B.n395 B.n394 585
R215 B.n396 B.n395 585
R216 B.n393 B.n178 585
R217 B.n178 B.n177 585
R218 B.n392 B.n391 585
R219 B.n391 B.n390 585
R220 B.n180 B.n179 585
R221 B.n181 B.n180 585
R222 B.n383 B.n382 585
R223 B.n384 B.n383 585
R224 B.n381 B.n186 585
R225 B.n186 B.n185 585
R226 B.n380 B.n379 585
R227 B.n379 B.n378 585
R228 B.n188 B.n187 585
R229 B.n189 B.n188 585
R230 B.n371 B.n370 585
R231 B.n372 B.n371 585
R232 B.n369 B.n194 585
R233 B.n194 B.n193 585
R234 B.n368 B.n367 585
R235 B.n367 B.n366 585
R236 B.n363 B.n198 585
R237 B.n362 B.n361 585
R238 B.n359 B.n199 585
R239 B.n359 B.n197 585
R240 B.n358 B.n357 585
R241 B.n356 B.n355 585
R242 B.n354 B.n201 585
R243 B.n352 B.n351 585
R244 B.n350 B.n202 585
R245 B.n349 B.n348 585
R246 B.n346 B.n203 585
R247 B.n344 B.n343 585
R248 B.n342 B.n204 585
R249 B.n341 B.n340 585
R250 B.n338 B.n205 585
R251 B.n336 B.n335 585
R252 B.n334 B.n206 585
R253 B.n333 B.n332 585
R254 B.n330 B.n207 585
R255 B.n328 B.n327 585
R256 B.n326 B.n208 585
R257 B.n325 B.n324 585
R258 B.n322 B.n209 585
R259 B.n320 B.n319 585
R260 B.n318 B.n210 585
R261 B.n317 B.n316 585
R262 B.n314 B.n211 585
R263 B.n312 B.n311 585
R264 B.n310 B.n212 585
R265 B.n308 B.n307 585
R266 B.n305 B.n215 585
R267 B.n303 B.n302 585
R268 B.n301 B.n216 585
R269 B.n300 B.n299 585
R270 B.n297 B.n217 585
R271 B.n295 B.n294 585
R272 B.n293 B.n218 585
R273 B.n292 B.n291 585
R274 B.n289 B.n288 585
R275 B.n287 B.n286 585
R276 B.n285 B.n223 585
R277 B.n283 B.n282 585
R278 B.n281 B.n224 585
R279 B.n280 B.n279 585
R280 B.n277 B.n225 585
R281 B.n275 B.n274 585
R282 B.n273 B.n226 585
R283 B.n272 B.n271 585
R284 B.n269 B.n227 585
R285 B.n267 B.n266 585
R286 B.n265 B.n228 585
R287 B.n264 B.n263 585
R288 B.n261 B.n229 585
R289 B.n259 B.n258 585
R290 B.n257 B.n230 585
R291 B.n256 B.n255 585
R292 B.n253 B.n231 585
R293 B.n251 B.n250 585
R294 B.n249 B.n232 585
R295 B.n248 B.n247 585
R296 B.n245 B.n233 585
R297 B.n243 B.n242 585
R298 B.n241 B.n234 585
R299 B.n240 B.n239 585
R300 B.n237 B.n235 585
R301 B.n196 B.n195 585
R302 B.n365 B.n364 585
R303 B.n366 B.n365 585
R304 B.n192 B.n191 585
R305 B.n193 B.n192 585
R306 B.n374 B.n373 585
R307 B.n373 B.n372 585
R308 B.n375 B.n190 585
R309 B.n190 B.n189 585
R310 B.n377 B.n376 585
R311 B.n378 B.n377 585
R312 B.n184 B.n183 585
R313 B.n185 B.n184 585
R314 B.n386 B.n385 585
R315 B.n385 B.n384 585
R316 B.n387 B.n182 585
R317 B.n182 B.n181 585
R318 B.n389 B.n388 585
R319 B.n390 B.n389 585
R320 B.n176 B.n175 585
R321 B.n177 B.n176 585
R322 B.n398 B.n397 585
R323 B.n397 B.n396 585
R324 B.n399 B.n174 585
R325 B.n174 B.n173 585
R326 B.n401 B.n400 585
R327 B.n402 B.n401 585
R328 B.n168 B.n167 585
R329 B.n169 B.n168 585
R330 B.n410 B.n409 585
R331 B.n409 B.n408 585
R332 B.n411 B.n166 585
R333 B.n166 B.n165 585
R334 B.n413 B.n412 585
R335 B.n414 B.n413 585
R336 B.n160 B.n159 585
R337 B.n161 B.n160 585
R338 B.n422 B.n421 585
R339 B.n421 B.n420 585
R340 B.n423 B.n158 585
R341 B.n158 B.n157 585
R342 B.n425 B.n424 585
R343 B.n426 B.n425 585
R344 B.n152 B.n151 585
R345 B.n153 B.n152 585
R346 B.n435 B.n434 585
R347 B.n434 B.n433 585
R348 B.n436 B.n150 585
R349 B.n432 B.n150 585
R350 B.n438 B.n437 585
R351 B.n439 B.n438 585
R352 B.n145 B.n144 585
R353 B.n146 B.n145 585
R354 B.n447 B.n446 585
R355 B.n446 B.n445 585
R356 B.n448 B.n143 585
R357 B.n143 B.n142 585
R358 B.n450 B.n449 585
R359 B.n451 B.n450 585
R360 B.n137 B.n136 585
R361 B.n138 B.n137 585
R362 B.n459 B.n458 585
R363 B.n458 B.n457 585
R364 B.n460 B.n135 585
R365 B.n135 B.n134 585
R366 B.n462 B.n461 585
R367 B.n463 B.n462 585
R368 B.n129 B.n128 585
R369 B.n130 B.n129 585
R370 B.n471 B.n470 585
R371 B.n470 B.n469 585
R372 B.n472 B.n127 585
R373 B.n127 B.n126 585
R374 B.n474 B.n473 585
R375 B.n475 B.n474 585
R376 B.n121 B.n120 585
R377 B.n122 B.n121 585
R378 B.n484 B.n483 585
R379 B.n483 B.n482 585
R380 B.n485 B.n119 585
R381 B.n119 B.n118 585
R382 B.n487 B.n486 585
R383 B.n488 B.n487 585
R384 B.n2 B.n0 585
R385 B.n4 B.n2 585
R386 B.n3 B.n1 585
R387 B.n759 B.n3 585
R388 B.n757 B.n756 585
R389 B.n758 B.n757 585
R390 B.n755 B.n9 585
R391 B.n9 B.n8 585
R392 B.n754 B.n753 585
R393 B.n753 B.n752 585
R394 B.n11 B.n10 585
R395 B.n751 B.n11 585
R396 B.n749 B.n748 585
R397 B.n750 B.n749 585
R398 B.n747 B.n16 585
R399 B.n16 B.n15 585
R400 B.n746 B.n745 585
R401 B.n745 B.n744 585
R402 B.n18 B.n17 585
R403 B.n743 B.n18 585
R404 B.n741 B.n740 585
R405 B.n742 B.n741 585
R406 B.n739 B.n23 585
R407 B.n23 B.n22 585
R408 B.n738 B.n737 585
R409 B.n737 B.n736 585
R410 B.n25 B.n24 585
R411 B.n735 B.n25 585
R412 B.n733 B.n732 585
R413 B.n734 B.n733 585
R414 B.n731 B.n30 585
R415 B.n30 B.n29 585
R416 B.n730 B.n729 585
R417 B.n729 B.n728 585
R418 B.n32 B.n31 585
R419 B.n727 B.n32 585
R420 B.n725 B.n724 585
R421 B.n726 B.n725 585
R422 B.n723 B.n36 585
R423 B.n39 B.n36 585
R424 B.n722 B.n721 585
R425 B.n721 B.n720 585
R426 B.n38 B.n37 585
R427 B.n719 B.n38 585
R428 B.n717 B.n716 585
R429 B.n718 B.n717 585
R430 B.n715 B.n44 585
R431 B.n44 B.n43 585
R432 B.n714 B.n713 585
R433 B.n713 B.n712 585
R434 B.n46 B.n45 585
R435 B.n711 B.n46 585
R436 B.n709 B.n708 585
R437 B.n710 B.n709 585
R438 B.n707 B.n51 585
R439 B.n51 B.n50 585
R440 B.n706 B.n705 585
R441 B.n705 B.n704 585
R442 B.n53 B.n52 585
R443 B.n703 B.n53 585
R444 B.n701 B.n700 585
R445 B.n702 B.n701 585
R446 B.n699 B.n58 585
R447 B.n58 B.n57 585
R448 B.n698 B.n697 585
R449 B.n697 B.n696 585
R450 B.n60 B.n59 585
R451 B.n695 B.n60 585
R452 B.n693 B.n692 585
R453 B.n694 B.n693 585
R454 B.n691 B.n65 585
R455 B.n65 B.n64 585
R456 B.n690 B.n689 585
R457 B.n689 B.n688 585
R458 B.n67 B.n66 585
R459 B.n687 B.n67 585
R460 B.n685 B.n684 585
R461 B.n686 B.n685 585
R462 B.n683 B.n72 585
R463 B.n72 B.n71 585
R464 B.n682 B.n681 585
R465 B.n681 B.n680 585
R466 B.n74 B.n73 585
R467 B.n679 B.n74 585
R468 B.n677 B.n676 585
R469 B.n678 B.n677 585
R470 B.n762 B.n761 585
R471 B.n761 B.n760 585
R472 B.n365 B.n198 545.355
R473 B.n677 B.n79 545.355
R474 B.n367 B.n196 545.355
R475 B.n115 B.n77 545.355
R476 B.n219 B.t17 276.252
R477 B.n100 B.t6 276.252
R478 B.n213 B.t11 276.252
R479 B.n94 B.t13 276.252
R480 B.n219 B.t15 259.027
R481 B.n213 B.t8 259.027
R482 B.n94 B.t12 259.027
R483 B.n100 B.t4 259.027
R484 B.n548 B.n78 256.663
R485 B.n550 B.n78 256.663
R486 B.n556 B.n78 256.663
R487 B.n558 B.n78 256.663
R488 B.n564 B.n78 256.663
R489 B.n566 B.n78 256.663
R490 B.n572 B.n78 256.663
R491 B.n574 B.n78 256.663
R492 B.n580 B.n78 256.663
R493 B.n582 B.n78 256.663
R494 B.n588 B.n78 256.663
R495 B.n590 B.n78 256.663
R496 B.n596 B.n78 256.663
R497 B.n598 B.n78 256.663
R498 B.n605 B.n78 256.663
R499 B.n607 B.n78 256.663
R500 B.n613 B.n78 256.663
R501 B.n615 B.n78 256.663
R502 B.n622 B.n78 256.663
R503 B.n624 B.n78 256.663
R504 B.n630 B.n78 256.663
R505 B.n632 B.n78 256.663
R506 B.n638 B.n78 256.663
R507 B.n640 B.n78 256.663
R508 B.n646 B.n78 256.663
R509 B.n648 B.n78 256.663
R510 B.n654 B.n78 256.663
R511 B.n656 B.n78 256.663
R512 B.n662 B.n78 256.663
R513 B.n664 B.n78 256.663
R514 B.n670 B.n78 256.663
R515 B.n672 B.n78 256.663
R516 B.n360 B.n197 256.663
R517 B.n200 B.n197 256.663
R518 B.n353 B.n197 256.663
R519 B.n347 B.n197 256.663
R520 B.n345 B.n197 256.663
R521 B.n339 B.n197 256.663
R522 B.n337 B.n197 256.663
R523 B.n331 B.n197 256.663
R524 B.n329 B.n197 256.663
R525 B.n323 B.n197 256.663
R526 B.n321 B.n197 256.663
R527 B.n315 B.n197 256.663
R528 B.n313 B.n197 256.663
R529 B.n306 B.n197 256.663
R530 B.n304 B.n197 256.663
R531 B.n298 B.n197 256.663
R532 B.n296 B.n197 256.663
R533 B.n290 B.n197 256.663
R534 B.n222 B.n197 256.663
R535 B.n284 B.n197 256.663
R536 B.n278 B.n197 256.663
R537 B.n276 B.n197 256.663
R538 B.n270 B.n197 256.663
R539 B.n268 B.n197 256.663
R540 B.n262 B.n197 256.663
R541 B.n260 B.n197 256.663
R542 B.n254 B.n197 256.663
R543 B.n252 B.n197 256.663
R544 B.n246 B.n197 256.663
R545 B.n244 B.n197 256.663
R546 B.n238 B.n197 256.663
R547 B.n236 B.n197 256.663
R548 B.n220 B.t16 201.392
R549 B.n101 B.t7 201.392
R550 B.n214 B.t10 201.392
R551 B.n95 B.t14 201.392
R552 B.n365 B.n192 163.367
R553 B.n373 B.n192 163.367
R554 B.n373 B.n190 163.367
R555 B.n377 B.n190 163.367
R556 B.n377 B.n184 163.367
R557 B.n385 B.n184 163.367
R558 B.n385 B.n182 163.367
R559 B.n389 B.n182 163.367
R560 B.n389 B.n176 163.367
R561 B.n397 B.n176 163.367
R562 B.n397 B.n174 163.367
R563 B.n401 B.n174 163.367
R564 B.n401 B.n168 163.367
R565 B.n409 B.n168 163.367
R566 B.n409 B.n166 163.367
R567 B.n413 B.n166 163.367
R568 B.n413 B.n160 163.367
R569 B.n421 B.n160 163.367
R570 B.n421 B.n158 163.367
R571 B.n425 B.n158 163.367
R572 B.n425 B.n152 163.367
R573 B.n434 B.n152 163.367
R574 B.n434 B.n150 163.367
R575 B.n438 B.n150 163.367
R576 B.n438 B.n145 163.367
R577 B.n446 B.n145 163.367
R578 B.n446 B.n143 163.367
R579 B.n450 B.n143 163.367
R580 B.n450 B.n137 163.367
R581 B.n458 B.n137 163.367
R582 B.n458 B.n135 163.367
R583 B.n462 B.n135 163.367
R584 B.n462 B.n129 163.367
R585 B.n470 B.n129 163.367
R586 B.n470 B.n127 163.367
R587 B.n474 B.n127 163.367
R588 B.n474 B.n121 163.367
R589 B.n483 B.n121 163.367
R590 B.n483 B.n119 163.367
R591 B.n487 B.n119 163.367
R592 B.n487 B.n2 163.367
R593 B.n761 B.n2 163.367
R594 B.n761 B.n3 163.367
R595 B.n757 B.n3 163.367
R596 B.n757 B.n9 163.367
R597 B.n753 B.n9 163.367
R598 B.n753 B.n11 163.367
R599 B.n749 B.n11 163.367
R600 B.n749 B.n16 163.367
R601 B.n745 B.n16 163.367
R602 B.n745 B.n18 163.367
R603 B.n741 B.n18 163.367
R604 B.n741 B.n23 163.367
R605 B.n737 B.n23 163.367
R606 B.n737 B.n25 163.367
R607 B.n733 B.n25 163.367
R608 B.n733 B.n30 163.367
R609 B.n729 B.n30 163.367
R610 B.n729 B.n32 163.367
R611 B.n725 B.n32 163.367
R612 B.n725 B.n36 163.367
R613 B.n721 B.n36 163.367
R614 B.n721 B.n38 163.367
R615 B.n717 B.n38 163.367
R616 B.n717 B.n44 163.367
R617 B.n713 B.n44 163.367
R618 B.n713 B.n46 163.367
R619 B.n709 B.n46 163.367
R620 B.n709 B.n51 163.367
R621 B.n705 B.n51 163.367
R622 B.n705 B.n53 163.367
R623 B.n701 B.n53 163.367
R624 B.n701 B.n58 163.367
R625 B.n697 B.n58 163.367
R626 B.n697 B.n60 163.367
R627 B.n693 B.n60 163.367
R628 B.n693 B.n65 163.367
R629 B.n689 B.n65 163.367
R630 B.n689 B.n67 163.367
R631 B.n685 B.n67 163.367
R632 B.n685 B.n72 163.367
R633 B.n681 B.n72 163.367
R634 B.n681 B.n74 163.367
R635 B.n677 B.n74 163.367
R636 B.n361 B.n359 163.367
R637 B.n359 B.n358 163.367
R638 B.n355 B.n354 163.367
R639 B.n352 B.n202 163.367
R640 B.n348 B.n346 163.367
R641 B.n344 B.n204 163.367
R642 B.n340 B.n338 163.367
R643 B.n336 B.n206 163.367
R644 B.n332 B.n330 163.367
R645 B.n328 B.n208 163.367
R646 B.n324 B.n322 163.367
R647 B.n320 B.n210 163.367
R648 B.n316 B.n314 163.367
R649 B.n312 B.n212 163.367
R650 B.n307 B.n305 163.367
R651 B.n303 B.n216 163.367
R652 B.n299 B.n297 163.367
R653 B.n295 B.n218 163.367
R654 B.n291 B.n289 163.367
R655 B.n286 B.n285 163.367
R656 B.n283 B.n224 163.367
R657 B.n279 B.n277 163.367
R658 B.n275 B.n226 163.367
R659 B.n271 B.n269 163.367
R660 B.n267 B.n228 163.367
R661 B.n263 B.n261 163.367
R662 B.n259 B.n230 163.367
R663 B.n255 B.n253 163.367
R664 B.n251 B.n232 163.367
R665 B.n247 B.n245 163.367
R666 B.n243 B.n234 163.367
R667 B.n239 B.n237 163.367
R668 B.n367 B.n194 163.367
R669 B.n371 B.n194 163.367
R670 B.n371 B.n188 163.367
R671 B.n379 B.n188 163.367
R672 B.n379 B.n186 163.367
R673 B.n383 B.n186 163.367
R674 B.n383 B.n180 163.367
R675 B.n391 B.n180 163.367
R676 B.n391 B.n178 163.367
R677 B.n395 B.n178 163.367
R678 B.n395 B.n172 163.367
R679 B.n403 B.n172 163.367
R680 B.n403 B.n170 163.367
R681 B.n407 B.n170 163.367
R682 B.n407 B.n164 163.367
R683 B.n415 B.n164 163.367
R684 B.n415 B.n162 163.367
R685 B.n419 B.n162 163.367
R686 B.n419 B.n156 163.367
R687 B.n427 B.n156 163.367
R688 B.n427 B.n154 163.367
R689 B.n431 B.n154 163.367
R690 B.n431 B.n149 163.367
R691 B.n440 B.n149 163.367
R692 B.n440 B.n147 163.367
R693 B.n444 B.n147 163.367
R694 B.n444 B.n141 163.367
R695 B.n452 B.n141 163.367
R696 B.n452 B.n139 163.367
R697 B.n456 B.n139 163.367
R698 B.n456 B.n133 163.367
R699 B.n464 B.n133 163.367
R700 B.n464 B.n131 163.367
R701 B.n468 B.n131 163.367
R702 B.n468 B.n125 163.367
R703 B.n476 B.n125 163.367
R704 B.n476 B.n123 163.367
R705 B.n481 B.n123 163.367
R706 B.n481 B.n117 163.367
R707 B.n489 B.n117 163.367
R708 B.n490 B.n489 163.367
R709 B.n490 B.n5 163.367
R710 B.n6 B.n5 163.367
R711 B.n7 B.n6 163.367
R712 B.n495 B.n7 163.367
R713 B.n495 B.n12 163.367
R714 B.n13 B.n12 163.367
R715 B.n14 B.n13 163.367
R716 B.n500 B.n14 163.367
R717 B.n500 B.n19 163.367
R718 B.n20 B.n19 163.367
R719 B.n21 B.n20 163.367
R720 B.n505 B.n21 163.367
R721 B.n505 B.n26 163.367
R722 B.n27 B.n26 163.367
R723 B.n28 B.n27 163.367
R724 B.n510 B.n28 163.367
R725 B.n510 B.n33 163.367
R726 B.n34 B.n33 163.367
R727 B.n35 B.n34 163.367
R728 B.n515 B.n35 163.367
R729 B.n515 B.n40 163.367
R730 B.n41 B.n40 163.367
R731 B.n42 B.n41 163.367
R732 B.n520 B.n42 163.367
R733 B.n520 B.n47 163.367
R734 B.n48 B.n47 163.367
R735 B.n49 B.n48 163.367
R736 B.n525 B.n49 163.367
R737 B.n525 B.n54 163.367
R738 B.n55 B.n54 163.367
R739 B.n56 B.n55 163.367
R740 B.n530 B.n56 163.367
R741 B.n530 B.n61 163.367
R742 B.n62 B.n61 163.367
R743 B.n63 B.n62 163.367
R744 B.n535 B.n63 163.367
R745 B.n535 B.n68 163.367
R746 B.n69 B.n68 163.367
R747 B.n70 B.n69 163.367
R748 B.n540 B.n70 163.367
R749 B.n540 B.n75 163.367
R750 B.n76 B.n75 163.367
R751 B.n77 B.n76 163.367
R752 B.n673 B.n671 163.367
R753 B.n669 B.n81 163.367
R754 B.n665 B.n663 163.367
R755 B.n661 B.n83 163.367
R756 B.n657 B.n655 163.367
R757 B.n653 B.n85 163.367
R758 B.n649 B.n647 163.367
R759 B.n645 B.n87 163.367
R760 B.n641 B.n639 163.367
R761 B.n637 B.n89 163.367
R762 B.n633 B.n631 163.367
R763 B.n629 B.n91 163.367
R764 B.n625 B.n623 163.367
R765 B.n621 B.n93 163.367
R766 B.n616 B.n614 163.367
R767 B.n612 B.n97 163.367
R768 B.n608 B.n606 163.367
R769 B.n604 B.n99 163.367
R770 B.n599 B.n597 163.367
R771 B.n595 B.n103 163.367
R772 B.n591 B.n589 163.367
R773 B.n587 B.n105 163.367
R774 B.n583 B.n581 163.367
R775 B.n579 B.n107 163.367
R776 B.n575 B.n573 163.367
R777 B.n571 B.n109 163.367
R778 B.n567 B.n565 163.367
R779 B.n563 B.n111 163.367
R780 B.n559 B.n557 163.367
R781 B.n555 B.n113 163.367
R782 B.n551 B.n549 163.367
R783 B.n547 B.n115 163.367
R784 B.n366 B.n197 117.999
R785 B.n678 B.n78 117.999
R786 B.n220 B.n219 74.8611
R787 B.n214 B.n213 74.8611
R788 B.n95 B.n94 74.8611
R789 B.n101 B.n100 74.8611
R790 B.n360 B.n198 71.676
R791 B.n358 B.n200 71.676
R792 B.n354 B.n353 71.676
R793 B.n347 B.n202 71.676
R794 B.n346 B.n345 71.676
R795 B.n339 B.n204 71.676
R796 B.n338 B.n337 71.676
R797 B.n331 B.n206 71.676
R798 B.n330 B.n329 71.676
R799 B.n323 B.n208 71.676
R800 B.n322 B.n321 71.676
R801 B.n315 B.n210 71.676
R802 B.n314 B.n313 71.676
R803 B.n306 B.n212 71.676
R804 B.n305 B.n304 71.676
R805 B.n298 B.n216 71.676
R806 B.n297 B.n296 71.676
R807 B.n290 B.n218 71.676
R808 B.n289 B.n222 71.676
R809 B.n285 B.n284 71.676
R810 B.n278 B.n224 71.676
R811 B.n277 B.n276 71.676
R812 B.n270 B.n226 71.676
R813 B.n269 B.n268 71.676
R814 B.n262 B.n228 71.676
R815 B.n261 B.n260 71.676
R816 B.n254 B.n230 71.676
R817 B.n253 B.n252 71.676
R818 B.n246 B.n232 71.676
R819 B.n245 B.n244 71.676
R820 B.n238 B.n234 71.676
R821 B.n237 B.n236 71.676
R822 B.n672 B.n79 71.676
R823 B.n671 B.n670 71.676
R824 B.n664 B.n81 71.676
R825 B.n663 B.n662 71.676
R826 B.n656 B.n83 71.676
R827 B.n655 B.n654 71.676
R828 B.n648 B.n85 71.676
R829 B.n647 B.n646 71.676
R830 B.n640 B.n87 71.676
R831 B.n639 B.n638 71.676
R832 B.n632 B.n89 71.676
R833 B.n631 B.n630 71.676
R834 B.n624 B.n91 71.676
R835 B.n623 B.n622 71.676
R836 B.n615 B.n93 71.676
R837 B.n614 B.n613 71.676
R838 B.n607 B.n97 71.676
R839 B.n606 B.n605 71.676
R840 B.n598 B.n99 71.676
R841 B.n597 B.n596 71.676
R842 B.n590 B.n103 71.676
R843 B.n589 B.n588 71.676
R844 B.n582 B.n105 71.676
R845 B.n581 B.n580 71.676
R846 B.n574 B.n107 71.676
R847 B.n573 B.n572 71.676
R848 B.n566 B.n109 71.676
R849 B.n565 B.n564 71.676
R850 B.n558 B.n111 71.676
R851 B.n557 B.n556 71.676
R852 B.n550 B.n113 71.676
R853 B.n549 B.n548 71.676
R854 B.n548 B.n547 71.676
R855 B.n551 B.n550 71.676
R856 B.n556 B.n555 71.676
R857 B.n559 B.n558 71.676
R858 B.n564 B.n563 71.676
R859 B.n567 B.n566 71.676
R860 B.n572 B.n571 71.676
R861 B.n575 B.n574 71.676
R862 B.n580 B.n579 71.676
R863 B.n583 B.n582 71.676
R864 B.n588 B.n587 71.676
R865 B.n591 B.n590 71.676
R866 B.n596 B.n595 71.676
R867 B.n599 B.n598 71.676
R868 B.n605 B.n604 71.676
R869 B.n608 B.n607 71.676
R870 B.n613 B.n612 71.676
R871 B.n616 B.n615 71.676
R872 B.n622 B.n621 71.676
R873 B.n625 B.n624 71.676
R874 B.n630 B.n629 71.676
R875 B.n633 B.n632 71.676
R876 B.n638 B.n637 71.676
R877 B.n641 B.n640 71.676
R878 B.n646 B.n645 71.676
R879 B.n649 B.n648 71.676
R880 B.n654 B.n653 71.676
R881 B.n657 B.n656 71.676
R882 B.n662 B.n661 71.676
R883 B.n665 B.n664 71.676
R884 B.n670 B.n669 71.676
R885 B.n673 B.n672 71.676
R886 B.n361 B.n360 71.676
R887 B.n355 B.n200 71.676
R888 B.n353 B.n352 71.676
R889 B.n348 B.n347 71.676
R890 B.n345 B.n344 71.676
R891 B.n340 B.n339 71.676
R892 B.n337 B.n336 71.676
R893 B.n332 B.n331 71.676
R894 B.n329 B.n328 71.676
R895 B.n324 B.n323 71.676
R896 B.n321 B.n320 71.676
R897 B.n316 B.n315 71.676
R898 B.n313 B.n312 71.676
R899 B.n307 B.n306 71.676
R900 B.n304 B.n303 71.676
R901 B.n299 B.n298 71.676
R902 B.n296 B.n295 71.676
R903 B.n291 B.n290 71.676
R904 B.n286 B.n222 71.676
R905 B.n284 B.n283 71.676
R906 B.n279 B.n278 71.676
R907 B.n276 B.n275 71.676
R908 B.n271 B.n270 71.676
R909 B.n268 B.n267 71.676
R910 B.n263 B.n262 71.676
R911 B.n260 B.n259 71.676
R912 B.n255 B.n254 71.676
R913 B.n252 B.n251 71.676
R914 B.n247 B.n246 71.676
R915 B.n244 B.n243 71.676
R916 B.n239 B.n238 71.676
R917 B.n236 B.n196 71.676
R918 B.n221 B.n220 59.5399
R919 B.n309 B.n214 59.5399
R920 B.n619 B.n95 59.5399
R921 B.n601 B.n101 59.5399
R922 B.n366 B.n193 59.4363
R923 B.n372 B.n193 59.4363
R924 B.n372 B.n189 59.4363
R925 B.n378 B.n189 59.4363
R926 B.n378 B.n185 59.4363
R927 B.n384 B.n185 59.4363
R928 B.n384 B.n181 59.4363
R929 B.n390 B.n181 59.4363
R930 B.n396 B.n177 59.4363
R931 B.n396 B.n173 59.4363
R932 B.n402 B.n173 59.4363
R933 B.n402 B.n169 59.4363
R934 B.n408 B.n169 59.4363
R935 B.n408 B.n165 59.4363
R936 B.n414 B.n165 59.4363
R937 B.n414 B.n161 59.4363
R938 B.n420 B.n161 59.4363
R939 B.n420 B.n157 59.4363
R940 B.n426 B.n157 59.4363
R941 B.n426 B.n153 59.4363
R942 B.n433 B.n153 59.4363
R943 B.n433 B.n432 59.4363
R944 B.n439 B.n146 59.4363
R945 B.n445 B.n146 59.4363
R946 B.n445 B.n142 59.4363
R947 B.n451 B.n142 59.4363
R948 B.n451 B.n138 59.4363
R949 B.n457 B.n138 59.4363
R950 B.n457 B.n134 59.4363
R951 B.n463 B.n134 59.4363
R952 B.n463 B.n130 59.4363
R953 B.n469 B.n130 59.4363
R954 B.n475 B.n126 59.4363
R955 B.n475 B.n122 59.4363
R956 B.n482 B.n122 59.4363
R957 B.n482 B.n118 59.4363
R958 B.n488 B.n118 59.4363
R959 B.n488 B.n4 59.4363
R960 B.n760 B.n4 59.4363
R961 B.n760 B.n759 59.4363
R962 B.n759 B.n758 59.4363
R963 B.n758 B.n8 59.4363
R964 B.n752 B.n8 59.4363
R965 B.n752 B.n751 59.4363
R966 B.n751 B.n750 59.4363
R967 B.n750 B.n15 59.4363
R968 B.n744 B.n743 59.4363
R969 B.n743 B.n742 59.4363
R970 B.n742 B.n22 59.4363
R971 B.n736 B.n22 59.4363
R972 B.n736 B.n735 59.4363
R973 B.n735 B.n734 59.4363
R974 B.n734 B.n29 59.4363
R975 B.n728 B.n29 59.4363
R976 B.n728 B.n727 59.4363
R977 B.n727 B.n726 59.4363
R978 B.n720 B.n39 59.4363
R979 B.n720 B.n719 59.4363
R980 B.n719 B.n718 59.4363
R981 B.n718 B.n43 59.4363
R982 B.n712 B.n43 59.4363
R983 B.n712 B.n711 59.4363
R984 B.n711 B.n710 59.4363
R985 B.n710 B.n50 59.4363
R986 B.n704 B.n50 59.4363
R987 B.n704 B.n703 59.4363
R988 B.n703 B.n702 59.4363
R989 B.n702 B.n57 59.4363
R990 B.n696 B.n57 59.4363
R991 B.n696 B.n695 59.4363
R992 B.n694 B.n64 59.4363
R993 B.n688 B.n64 59.4363
R994 B.n688 B.n687 59.4363
R995 B.n687 B.n686 59.4363
R996 B.n686 B.n71 59.4363
R997 B.n680 B.n71 59.4363
R998 B.n680 B.n679 59.4363
R999 B.n679 B.n678 59.4363
R1000 B.n390 B.t9 48.0736
R1001 B.t5 B.n694 48.0736
R1002 B.n469 B.t1 42.8293
R1003 B.n744 B.t0 42.8293
R1004 B.n439 B.t3 37.5849
R1005 B.n726 B.t2 37.5849
R1006 B.n545 B.n544 35.4346
R1007 B.n676 B.n675 35.4346
R1008 B.n368 B.n195 35.4346
R1009 B.n364 B.n363 35.4346
R1010 B.n432 B.t3 21.8519
R1011 B.n39 B.t2 21.8519
R1012 B B.n762 18.0485
R1013 B.t1 B.n126 16.6076
R1014 B.t0 B.n15 16.6076
R1015 B.t9 B.n177 11.3632
R1016 B.n695 B.t5 11.3632
R1017 B.n675 B.n674 10.6151
R1018 B.n674 B.n80 10.6151
R1019 B.n668 B.n80 10.6151
R1020 B.n668 B.n667 10.6151
R1021 B.n667 B.n666 10.6151
R1022 B.n666 B.n82 10.6151
R1023 B.n660 B.n82 10.6151
R1024 B.n660 B.n659 10.6151
R1025 B.n659 B.n658 10.6151
R1026 B.n658 B.n84 10.6151
R1027 B.n652 B.n84 10.6151
R1028 B.n652 B.n651 10.6151
R1029 B.n651 B.n650 10.6151
R1030 B.n650 B.n86 10.6151
R1031 B.n644 B.n86 10.6151
R1032 B.n644 B.n643 10.6151
R1033 B.n643 B.n642 10.6151
R1034 B.n642 B.n88 10.6151
R1035 B.n636 B.n88 10.6151
R1036 B.n636 B.n635 10.6151
R1037 B.n635 B.n634 10.6151
R1038 B.n634 B.n90 10.6151
R1039 B.n628 B.n90 10.6151
R1040 B.n628 B.n627 10.6151
R1041 B.n627 B.n626 10.6151
R1042 B.n626 B.n92 10.6151
R1043 B.n620 B.n92 10.6151
R1044 B.n618 B.n617 10.6151
R1045 B.n617 B.n96 10.6151
R1046 B.n611 B.n96 10.6151
R1047 B.n611 B.n610 10.6151
R1048 B.n610 B.n609 10.6151
R1049 B.n609 B.n98 10.6151
R1050 B.n603 B.n98 10.6151
R1051 B.n603 B.n602 10.6151
R1052 B.n600 B.n102 10.6151
R1053 B.n594 B.n102 10.6151
R1054 B.n594 B.n593 10.6151
R1055 B.n593 B.n592 10.6151
R1056 B.n592 B.n104 10.6151
R1057 B.n586 B.n104 10.6151
R1058 B.n586 B.n585 10.6151
R1059 B.n585 B.n584 10.6151
R1060 B.n584 B.n106 10.6151
R1061 B.n578 B.n106 10.6151
R1062 B.n578 B.n577 10.6151
R1063 B.n577 B.n576 10.6151
R1064 B.n576 B.n108 10.6151
R1065 B.n570 B.n108 10.6151
R1066 B.n570 B.n569 10.6151
R1067 B.n569 B.n568 10.6151
R1068 B.n568 B.n110 10.6151
R1069 B.n562 B.n110 10.6151
R1070 B.n562 B.n561 10.6151
R1071 B.n561 B.n560 10.6151
R1072 B.n560 B.n112 10.6151
R1073 B.n554 B.n112 10.6151
R1074 B.n554 B.n553 10.6151
R1075 B.n553 B.n552 10.6151
R1076 B.n552 B.n114 10.6151
R1077 B.n546 B.n114 10.6151
R1078 B.n546 B.n545 10.6151
R1079 B.n369 B.n368 10.6151
R1080 B.n370 B.n369 10.6151
R1081 B.n370 B.n187 10.6151
R1082 B.n380 B.n187 10.6151
R1083 B.n381 B.n380 10.6151
R1084 B.n382 B.n381 10.6151
R1085 B.n382 B.n179 10.6151
R1086 B.n392 B.n179 10.6151
R1087 B.n393 B.n392 10.6151
R1088 B.n394 B.n393 10.6151
R1089 B.n394 B.n171 10.6151
R1090 B.n404 B.n171 10.6151
R1091 B.n405 B.n404 10.6151
R1092 B.n406 B.n405 10.6151
R1093 B.n406 B.n163 10.6151
R1094 B.n416 B.n163 10.6151
R1095 B.n417 B.n416 10.6151
R1096 B.n418 B.n417 10.6151
R1097 B.n418 B.n155 10.6151
R1098 B.n428 B.n155 10.6151
R1099 B.n429 B.n428 10.6151
R1100 B.n430 B.n429 10.6151
R1101 B.n430 B.n148 10.6151
R1102 B.n441 B.n148 10.6151
R1103 B.n442 B.n441 10.6151
R1104 B.n443 B.n442 10.6151
R1105 B.n443 B.n140 10.6151
R1106 B.n453 B.n140 10.6151
R1107 B.n454 B.n453 10.6151
R1108 B.n455 B.n454 10.6151
R1109 B.n455 B.n132 10.6151
R1110 B.n465 B.n132 10.6151
R1111 B.n466 B.n465 10.6151
R1112 B.n467 B.n466 10.6151
R1113 B.n467 B.n124 10.6151
R1114 B.n477 B.n124 10.6151
R1115 B.n478 B.n477 10.6151
R1116 B.n480 B.n478 10.6151
R1117 B.n480 B.n479 10.6151
R1118 B.n479 B.n116 10.6151
R1119 B.n491 B.n116 10.6151
R1120 B.n492 B.n491 10.6151
R1121 B.n493 B.n492 10.6151
R1122 B.n494 B.n493 10.6151
R1123 B.n496 B.n494 10.6151
R1124 B.n497 B.n496 10.6151
R1125 B.n498 B.n497 10.6151
R1126 B.n499 B.n498 10.6151
R1127 B.n501 B.n499 10.6151
R1128 B.n502 B.n501 10.6151
R1129 B.n503 B.n502 10.6151
R1130 B.n504 B.n503 10.6151
R1131 B.n506 B.n504 10.6151
R1132 B.n507 B.n506 10.6151
R1133 B.n508 B.n507 10.6151
R1134 B.n509 B.n508 10.6151
R1135 B.n511 B.n509 10.6151
R1136 B.n512 B.n511 10.6151
R1137 B.n513 B.n512 10.6151
R1138 B.n514 B.n513 10.6151
R1139 B.n516 B.n514 10.6151
R1140 B.n517 B.n516 10.6151
R1141 B.n518 B.n517 10.6151
R1142 B.n519 B.n518 10.6151
R1143 B.n521 B.n519 10.6151
R1144 B.n522 B.n521 10.6151
R1145 B.n523 B.n522 10.6151
R1146 B.n524 B.n523 10.6151
R1147 B.n526 B.n524 10.6151
R1148 B.n527 B.n526 10.6151
R1149 B.n528 B.n527 10.6151
R1150 B.n529 B.n528 10.6151
R1151 B.n531 B.n529 10.6151
R1152 B.n532 B.n531 10.6151
R1153 B.n533 B.n532 10.6151
R1154 B.n534 B.n533 10.6151
R1155 B.n536 B.n534 10.6151
R1156 B.n537 B.n536 10.6151
R1157 B.n538 B.n537 10.6151
R1158 B.n539 B.n538 10.6151
R1159 B.n541 B.n539 10.6151
R1160 B.n542 B.n541 10.6151
R1161 B.n543 B.n542 10.6151
R1162 B.n544 B.n543 10.6151
R1163 B.n363 B.n362 10.6151
R1164 B.n362 B.n199 10.6151
R1165 B.n357 B.n199 10.6151
R1166 B.n357 B.n356 10.6151
R1167 B.n356 B.n201 10.6151
R1168 B.n351 B.n201 10.6151
R1169 B.n351 B.n350 10.6151
R1170 B.n350 B.n349 10.6151
R1171 B.n349 B.n203 10.6151
R1172 B.n343 B.n203 10.6151
R1173 B.n343 B.n342 10.6151
R1174 B.n342 B.n341 10.6151
R1175 B.n341 B.n205 10.6151
R1176 B.n335 B.n205 10.6151
R1177 B.n335 B.n334 10.6151
R1178 B.n334 B.n333 10.6151
R1179 B.n333 B.n207 10.6151
R1180 B.n327 B.n207 10.6151
R1181 B.n327 B.n326 10.6151
R1182 B.n326 B.n325 10.6151
R1183 B.n325 B.n209 10.6151
R1184 B.n319 B.n209 10.6151
R1185 B.n319 B.n318 10.6151
R1186 B.n318 B.n317 10.6151
R1187 B.n317 B.n211 10.6151
R1188 B.n311 B.n211 10.6151
R1189 B.n311 B.n310 10.6151
R1190 B.n308 B.n215 10.6151
R1191 B.n302 B.n215 10.6151
R1192 B.n302 B.n301 10.6151
R1193 B.n301 B.n300 10.6151
R1194 B.n300 B.n217 10.6151
R1195 B.n294 B.n217 10.6151
R1196 B.n294 B.n293 10.6151
R1197 B.n293 B.n292 10.6151
R1198 B.n288 B.n287 10.6151
R1199 B.n287 B.n223 10.6151
R1200 B.n282 B.n223 10.6151
R1201 B.n282 B.n281 10.6151
R1202 B.n281 B.n280 10.6151
R1203 B.n280 B.n225 10.6151
R1204 B.n274 B.n225 10.6151
R1205 B.n274 B.n273 10.6151
R1206 B.n273 B.n272 10.6151
R1207 B.n272 B.n227 10.6151
R1208 B.n266 B.n227 10.6151
R1209 B.n266 B.n265 10.6151
R1210 B.n265 B.n264 10.6151
R1211 B.n264 B.n229 10.6151
R1212 B.n258 B.n229 10.6151
R1213 B.n258 B.n257 10.6151
R1214 B.n257 B.n256 10.6151
R1215 B.n256 B.n231 10.6151
R1216 B.n250 B.n231 10.6151
R1217 B.n250 B.n249 10.6151
R1218 B.n249 B.n248 10.6151
R1219 B.n248 B.n233 10.6151
R1220 B.n242 B.n233 10.6151
R1221 B.n242 B.n241 10.6151
R1222 B.n241 B.n240 10.6151
R1223 B.n240 B.n235 10.6151
R1224 B.n235 B.n195 10.6151
R1225 B.n364 B.n191 10.6151
R1226 B.n374 B.n191 10.6151
R1227 B.n375 B.n374 10.6151
R1228 B.n376 B.n375 10.6151
R1229 B.n376 B.n183 10.6151
R1230 B.n386 B.n183 10.6151
R1231 B.n387 B.n386 10.6151
R1232 B.n388 B.n387 10.6151
R1233 B.n388 B.n175 10.6151
R1234 B.n398 B.n175 10.6151
R1235 B.n399 B.n398 10.6151
R1236 B.n400 B.n399 10.6151
R1237 B.n400 B.n167 10.6151
R1238 B.n410 B.n167 10.6151
R1239 B.n411 B.n410 10.6151
R1240 B.n412 B.n411 10.6151
R1241 B.n412 B.n159 10.6151
R1242 B.n422 B.n159 10.6151
R1243 B.n423 B.n422 10.6151
R1244 B.n424 B.n423 10.6151
R1245 B.n424 B.n151 10.6151
R1246 B.n435 B.n151 10.6151
R1247 B.n436 B.n435 10.6151
R1248 B.n437 B.n436 10.6151
R1249 B.n437 B.n144 10.6151
R1250 B.n447 B.n144 10.6151
R1251 B.n448 B.n447 10.6151
R1252 B.n449 B.n448 10.6151
R1253 B.n449 B.n136 10.6151
R1254 B.n459 B.n136 10.6151
R1255 B.n460 B.n459 10.6151
R1256 B.n461 B.n460 10.6151
R1257 B.n461 B.n128 10.6151
R1258 B.n471 B.n128 10.6151
R1259 B.n472 B.n471 10.6151
R1260 B.n473 B.n472 10.6151
R1261 B.n473 B.n120 10.6151
R1262 B.n484 B.n120 10.6151
R1263 B.n485 B.n484 10.6151
R1264 B.n486 B.n485 10.6151
R1265 B.n486 B.n0 10.6151
R1266 B.n756 B.n1 10.6151
R1267 B.n756 B.n755 10.6151
R1268 B.n755 B.n754 10.6151
R1269 B.n754 B.n10 10.6151
R1270 B.n748 B.n10 10.6151
R1271 B.n748 B.n747 10.6151
R1272 B.n747 B.n746 10.6151
R1273 B.n746 B.n17 10.6151
R1274 B.n740 B.n17 10.6151
R1275 B.n740 B.n739 10.6151
R1276 B.n739 B.n738 10.6151
R1277 B.n738 B.n24 10.6151
R1278 B.n732 B.n24 10.6151
R1279 B.n732 B.n731 10.6151
R1280 B.n731 B.n730 10.6151
R1281 B.n730 B.n31 10.6151
R1282 B.n724 B.n31 10.6151
R1283 B.n724 B.n723 10.6151
R1284 B.n723 B.n722 10.6151
R1285 B.n722 B.n37 10.6151
R1286 B.n716 B.n37 10.6151
R1287 B.n716 B.n715 10.6151
R1288 B.n715 B.n714 10.6151
R1289 B.n714 B.n45 10.6151
R1290 B.n708 B.n45 10.6151
R1291 B.n708 B.n707 10.6151
R1292 B.n707 B.n706 10.6151
R1293 B.n706 B.n52 10.6151
R1294 B.n700 B.n52 10.6151
R1295 B.n700 B.n699 10.6151
R1296 B.n699 B.n698 10.6151
R1297 B.n698 B.n59 10.6151
R1298 B.n692 B.n59 10.6151
R1299 B.n692 B.n691 10.6151
R1300 B.n691 B.n690 10.6151
R1301 B.n690 B.n66 10.6151
R1302 B.n684 B.n66 10.6151
R1303 B.n684 B.n683 10.6151
R1304 B.n683 B.n682 10.6151
R1305 B.n682 B.n73 10.6151
R1306 B.n676 B.n73 10.6151
R1307 B.n619 B.n618 6.5566
R1308 B.n602 B.n601 6.5566
R1309 B.n309 B.n308 6.5566
R1310 B.n292 B.n221 6.5566
R1311 B.n620 B.n619 4.05904
R1312 B.n601 B.n600 4.05904
R1313 B.n310 B.n309 4.05904
R1314 B.n288 B.n221 4.05904
R1315 B.n762 B.n0 2.81026
R1316 B.n762 B.n1 2.81026
R1317 VP.n19 VP.n18 161.3
R1318 VP.n17 VP.n1 161.3
R1319 VP.n16 VP.n15 161.3
R1320 VP.n14 VP.n2 161.3
R1321 VP.n13 VP.n12 161.3
R1322 VP.n11 VP.n3 161.3
R1323 VP.n10 VP.n9 161.3
R1324 VP.n8 VP.n4 161.3
R1325 VP.n5 VP.t1 84.4852
R1326 VP.n5 VP.t0 83.2584
R1327 VP.n7 VP.n6 81.2593
R1328 VP.n20 VP.n0 81.2593
R1329 VP.n12 VP.n2 56.5193
R1330 VP.n6 VP.t3 49.9073
R1331 VP.n0 VP.t2 49.9073
R1332 VP.n7 VP.n5 47.8266
R1333 VP.n10 VP.n4 24.4675
R1334 VP.n11 VP.n10 24.4675
R1335 VP.n12 VP.n11 24.4675
R1336 VP.n16 VP.n2 24.4675
R1337 VP.n17 VP.n16 24.4675
R1338 VP.n18 VP.n17 24.4675
R1339 VP.n6 VP.n4 8.80862
R1340 VP.n18 VP.n0 8.80862
R1341 VP.n8 VP.n7 0.354971
R1342 VP.n20 VP.n19 0.354971
R1343 VP VP.n20 0.26696
R1344 VP.n9 VP.n8 0.189894
R1345 VP.n9 VP.n3 0.189894
R1346 VP.n13 VP.n3 0.189894
R1347 VP.n14 VP.n13 0.189894
R1348 VP.n15 VP.n14 0.189894
R1349 VP.n15 VP.n1 0.189894
R1350 VP.n19 VP.n1 0.189894
R1351 VTAIL.n282 VTAIL.n252 214.453
R1352 VTAIL.n30 VTAIL.n0 214.453
R1353 VTAIL.n66 VTAIL.n36 214.453
R1354 VTAIL.n102 VTAIL.n72 214.453
R1355 VTAIL.n246 VTAIL.n216 214.453
R1356 VTAIL.n210 VTAIL.n180 214.453
R1357 VTAIL.n174 VTAIL.n144 214.453
R1358 VTAIL.n138 VTAIL.n108 214.453
R1359 VTAIL.n265 VTAIL.n264 185
R1360 VTAIL.n267 VTAIL.n266 185
R1361 VTAIL.n260 VTAIL.n259 185
R1362 VTAIL.n273 VTAIL.n272 185
R1363 VTAIL.n275 VTAIL.n274 185
R1364 VTAIL.n256 VTAIL.n255 185
R1365 VTAIL.n281 VTAIL.n280 185
R1366 VTAIL.n283 VTAIL.n282 185
R1367 VTAIL.n13 VTAIL.n12 185
R1368 VTAIL.n15 VTAIL.n14 185
R1369 VTAIL.n8 VTAIL.n7 185
R1370 VTAIL.n21 VTAIL.n20 185
R1371 VTAIL.n23 VTAIL.n22 185
R1372 VTAIL.n4 VTAIL.n3 185
R1373 VTAIL.n29 VTAIL.n28 185
R1374 VTAIL.n31 VTAIL.n30 185
R1375 VTAIL.n49 VTAIL.n48 185
R1376 VTAIL.n51 VTAIL.n50 185
R1377 VTAIL.n44 VTAIL.n43 185
R1378 VTAIL.n57 VTAIL.n56 185
R1379 VTAIL.n59 VTAIL.n58 185
R1380 VTAIL.n40 VTAIL.n39 185
R1381 VTAIL.n65 VTAIL.n64 185
R1382 VTAIL.n67 VTAIL.n66 185
R1383 VTAIL.n85 VTAIL.n84 185
R1384 VTAIL.n87 VTAIL.n86 185
R1385 VTAIL.n80 VTAIL.n79 185
R1386 VTAIL.n93 VTAIL.n92 185
R1387 VTAIL.n95 VTAIL.n94 185
R1388 VTAIL.n76 VTAIL.n75 185
R1389 VTAIL.n101 VTAIL.n100 185
R1390 VTAIL.n103 VTAIL.n102 185
R1391 VTAIL.n247 VTAIL.n246 185
R1392 VTAIL.n245 VTAIL.n244 185
R1393 VTAIL.n220 VTAIL.n219 185
R1394 VTAIL.n239 VTAIL.n238 185
R1395 VTAIL.n237 VTAIL.n236 185
R1396 VTAIL.n224 VTAIL.n223 185
R1397 VTAIL.n231 VTAIL.n230 185
R1398 VTAIL.n229 VTAIL.n228 185
R1399 VTAIL.n211 VTAIL.n210 185
R1400 VTAIL.n209 VTAIL.n208 185
R1401 VTAIL.n184 VTAIL.n183 185
R1402 VTAIL.n203 VTAIL.n202 185
R1403 VTAIL.n201 VTAIL.n200 185
R1404 VTAIL.n188 VTAIL.n187 185
R1405 VTAIL.n195 VTAIL.n194 185
R1406 VTAIL.n193 VTAIL.n192 185
R1407 VTAIL.n175 VTAIL.n174 185
R1408 VTAIL.n173 VTAIL.n172 185
R1409 VTAIL.n148 VTAIL.n147 185
R1410 VTAIL.n167 VTAIL.n166 185
R1411 VTAIL.n165 VTAIL.n164 185
R1412 VTAIL.n152 VTAIL.n151 185
R1413 VTAIL.n159 VTAIL.n158 185
R1414 VTAIL.n157 VTAIL.n156 185
R1415 VTAIL.n139 VTAIL.n138 185
R1416 VTAIL.n137 VTAIL.n136 185
R1417 VTAIL.n112 VTAIL.n111 185
R1418 VTAIL.n131 VTAIL.n130 185
R1419 VTAIL.n129 VTAIL.n128 185
R1420 VTAIL.n116 VTAIL.n115 185
R1421 VTAIL.n123 VTAIL.n122 185
R1422 VTAIL.n121 VTAIL.n120 185
R1423 VTAIL.n263 VTAIL.t2 149.524
R1424 VTAIL.n11 VTAIL.t0 149.524
R1425 VTAIL.n47 VTAIL.t5 149.524
R1426 VTAIL.n83 VTAIL.t4 149.524
R1427 VTAIL.n227 VTAIL.t6 149.524
R1428 VTAIL.n191 VTAIL.t7 149.524
R1429 VTAIL.n155 VTAIL.t1 149.524
R1430 VTAIL.n119 VTAIL.t3 149.524
R1431 VTAIL.n266 VTAIL.n265 104.615
R1432 VTAIL.n266 VTAIL.n259 104.615
R1433 VTAIL.n273 VTAIL.n259 104.615
R1434 VTAIL.n274 VTAIL.n273 104.615
R1435 VTAIL.n274 VTAIL.n255 104.615
R1436 VTAIL.n281 VTAIL.n255 104.615
R1437 VTAIL.n282 VTAIL.n281 104.615
R1438 VTAIL.n14 VTAIL.n13 104.615
R1439 VTAIL.n14 VTAIL.n7 104.615
R1440 VTAIL.n21 VTAIL.n7 104.615
R1441 VTAIL.n22 VTAIL.n21 104.615
R1442 VTAIL.n22 VTAIL.n3 104.615
R1443 VTAIL.n29 VTAIL.n3 104.615
R1444 VTAIL.n30 VTAIL.n29 104.615
R1445 VTAIL.n50 VTAIL.n49 104.615
R1446 VTAIL.n50 VTAIL.n43 104.615
R1447 VTAIL.n57 VTAIL.n43 104.615
R1448 VTAIL.n58 VTAIL.n57 104.615
R1449 VTAIL.n58 VTAIL.n39 104.615
R1450 VTAIL.n65 VTAIL.n39 104.615
R1451 VTAIL.n66 VTAIL.n65 104.615
R1452 VTAIL.n86 VTAIL.n85 104.615
R1453 VTAIL.n86 VTAIL.n79 104.615
R1454 VTAIL.n93 VTAIL.n79 104.615
R1455 VTAIL.n94 VTAIL.n93 104.615
R1456 VTAIL.n94 VTAIL.n75 104.615
R1457 VTAIL.n101 VTAIL.n75 104.615
R1458 VTAIL.n102 VTAIL.n101 104.615
R1459 VTAIL.n246 VTAIL.n245 104.615
R1460 VTAIL.n245 VTAIL.n219 104.615
R1461 VTAIL.n238 VTAIL.n219 104.615
R1462 VTAIL.n238 VTAIL.n237 104.615
R1463 VTAIL.n237 VTAIL.n223 104.615
R1464 VTAIL.n230 VTAIL.n223 104.615
R1465 VTAIL.n230 VTAIL.n229 104.615
R1466 VTAIL.n210 VTAIL.n209 104.615
R1467 VTAIL.n209 VTAIL.n183 104.615
R1468 VTAIL.n202 VTAIL.n183 104.615
R1469 VTAIL.n202 VTAIL.n201 104.615
R1470 VTAIL.n201 VTAIL.n187 104.615
R1471 VTAIL.n194 VTAIL.n187 104.615
R1472 VTAIL.n194 VTAIL.n193 104.615
R1473 VTAIL.n174 VTAIL.n173 104.615
R1474 VTAIL.n173 VTAIL.n147 104.615
R1475 VTAIL.n166 VTAIL.n147 104.615
R1476 VTAIL.n166 VTAIL.n165 104.615
R1477 VTAIL.n165 VTAIL.n151 104.615
R1478 VTAIL.n158 VTAIL.n151 104.615
R1479 VTAIL.n158 VTAIL.n157 104.615
R1480 VTAIL.n138 VTAIL.n137 104.615
R1481 VTAIL.n137 VTAIL.n111 104.615
R1482 VTAIL.n130 VTAIL.n111 104.615
R1483 VTAIL.n130 VTAIL.n129 104.615
R1484 VTAIL.n129 VTAIL.n115 104.615
R1485 VTAIL.n122 VTAIL.n115 104.615
R1486 VTAIL.n122 VTAIL.n121 104.615
R1487 VTAIL.n265 VTAIL.t2 52.3082
R1488 VTAIL.n13 VTAIL.t0 52.3082
R1489 VTAIL.n49 VTAIL.t5 52.3082
R1490 VTAIL.n85 VTAIL.t4 52.3082
R1491 VTAIL.n229 VTAIL.t6 52.3082
R1492 VTAIL.n193 VTAIL.t7 52.3082
R1493 VTAIL.n157 VTAIL.t1 52.3082
R1494 VTAIL.n121 VTAIL.t3 52.3082
R1495 VTAIL.n287 VTAIL.n286 36.646
R1496 VTAIL.n35 VTAIL.n34 36.646
R1497 VTAIL.n71 VTAIL.n70 36.646
R1498 VTAIL.n107 VTAIL.n106 36.646
R1499 VTAIL.n251 VTAIL.n250 36.646
R1500 VTAIL.n215 VTAIL.n214 36.646
R1501 VTAIL.n179 VTAIL.n178 36.646
R1502 VTAIL.n143 VTAIL.n142 36.646
R1503 VTAIL.n287 VTAIL.n251 21.9962
R1504 VTAIL.n143 VTAIL.n107 21.9962
R1505 VTAIL.n284 VTAIL.n283 12.8005
R1506 VTAIL.n32 VTAIL.n31 12.8005
R1507 VTAIL.n68 VTAIL.n67 12.8005
R1508 VTAIL.n104 VTAIL.n103 12.8005
R1509 VTAIL.n248 VTAIL.n247 12.8005
R1510 VTAIL.n212 VTAIL.n211 12.8005
R1511 VTAIL.n176 VTAIL.n175 12.8005
R1512 VTAIL.n140 VTAIL.n139 12.8005
R1513 VTAIL.n280 VTAIL.n254 12.0247
R1514 VTAIL.n28 VTAIL.n2 12.0247
R1515 VTAIL.n64 VTAIL.n38 12.0247
R1516 VTAIL.n100 VTAIL.n74 12.0247
R1517 VTAIL.n244 VTAIL.n218 12.0247
R1518 VTAIL.n208 VTAIL.n182 12.0247
R1519 VTAIL.n172 VTAIL.n146 12.0247
R1520 VTAIL.n136 VTAIL.n110 12.0247
R1521 VTAIL.n279 VTAIL.n256 11.249
R1522 VTAIL.n27 VTAIL.n4 11.249
R1523 VTAIL.n63 VTAIL.n40 11.249
R1524 VTAIL.n99 VTAIL.n76 11.249
R1525 VTAIL.n243 VTAIL.n220 11.249
R1526 VTAIL.n207 VTAIL.n184 11.249
R1527 VTAIL.n171 VTAIL.n148 11.249
R1528 VTAIL.n135 VTAIL.n112 11.249
R1529 VTAIL.n276 VTAIL.n275 10.4732
R1530 VTAIL.n24 VTAIL.n23 10.4732
R1531 VTAIL.n60 VTAIL.n59 10.4732
R1532 VTAIL.n96 VTAIL.n95 10.4732
R1533 VTAIL.n240 VTAIL.n239 10.4732
R1534 VTAIL.n204 VTAIL.n203 10.4732
R1535 VTAIL.n168 VTAIL.n167 10.4732
R1536 VTAIL.n132 VTAIL.n131 10.4732
R1537 VTAIL.n264 VTAIL.n263 10.2747
R1538 VTAIL.n12 VTAIL.n11 10.2747
R1539 VTAIL.n48 VTAIL.n47 10.2747
R1540 VTAIL.n84 VTAIL.n83 10.2747
R1541 VTAIL.n228 VTAIL.n227 10.2747
R1542 VTAIL.n192 VTAIL.n191 10.2747
R1543 VTAIL.n156 VTAIL.n155 10.2747
R1544 VTAIL.n120 VTAIL.n119 10.2747
R1545 VTAIL.n272 VTAIL.n258 9.69747
R1546 VTAIL.n20 VTAIL.n6 9.69747
R1547 VTAIL.n56 VTAIL.n42 9.69747
R1548 VTAIL.n92 VTAIL.n78 9.69747
R1549 VTAIL.n236 VTAIL.n222 9.69747
R1550 VTAIL.n200 VTAIL.n186 9.69747
R1551 VTAIL.n164 VTAIL.n150 9.69747
R1552 VTAIL.n128 VTAIL.n114 9.69747
R1553 VTAIL.n286 VTAIL.n285 9.45567
R1554 VTAIL.n34 VTAIL.n33 9.45567
R1555 VTAIL.n70 VTAIL.n69 9.45567
R1556 VTAIL.n106 VTAIL.n105 9.45567
R1557 VTAIL.n250 VTAIL.n249 9.45567
R1558 VTAIL.n214 VTAIL.n213 9.45567
R1559 VTAIL.n178 VTAIL.n177 9.45567
R1560 VTAIL.n142 VTAIL.n141 9.45567
R1561 VTAIL.n262 VTAIL.n261 9.3005
R1562 VTAIL.n269 VTAIL.n268 9.3005
R1563 VTAIL.n271 VTAIL.n270 9.3005
R1564 VTAIL.n258 VTAIL.n257 9.3005
R1565 VTAIL.n277 VTAIL.n276 9.3005
R1566 VTAIL.n279 VTAIL.n278 9.3005
R1567 VTAIL.n254 VTAIL.n253 9.3005
R1568 VTAIL.n285 VTAIL.n284 9.3005
R1569 VTAIL.n10 VTAIL.n9 9.3005
R1570 VTAIL.n17 VTAIL.n16 9.3005
R1571 VTAIL.n19 VTAIL.n18 9.3005
R1572 VTAIL.n6 VTAIL.n5 9.3005
R1573 VTAIL.n25 VTAIL.n24 9.3005
R1574 VTAIL.n27 VTAIL.n26 9.3005
R1575 VTAIL.n2 VTAIL.n1 9.3005
R1576 VTAIL.n33 VTAIL.n32 9.3005
R1577 VTAIL.n46 VTAIL.n45 9.3005
R1578 VTAIL.n53 VTAIL.n52 9.3005
R1579 VTAIL.n55 VTAIL.n54 9.3005
R1580 VTAIL.n42 VTAIL.n41 9.3005
R1581 VTAIL.n61 VTAIL.n60 9.3005
R1582 VTAIL.n63 VTAIL.n62 9.3005
R1583 VTAIL.n38 VTAIL.n37 9.3005
R1584 VTAIL.n69 VTAIL.n68 9.3005
R1585 VTAIL.n82 VTAIL.n81 9.3005
R1586 VTAIL.n89 VTAIL.n88 9.3005
R1587 VTAIL.n91 VTAIL.n90 9.3005
R1588 VTAIL.n78 VTAIL.n77 9.3005
R1589 VTAIL.n97 VTAIL.n96 9.3005
R1590 VTAIL.n99 VTAIL.n98 9.3005
R1591 VTAIL.n74 VTAIL.n73 9.3005
R1592 VTAIL.n105 VTAIL.n104 9.3005
R1593 VTAIL.n226 VTAIL.n225 9.3005
R1594 VTAIL.n233 VTAIL.n232 9.3005
R1595 VTAIL.n235 VTAIL.n234 9.3005
R1596 VTAIL.n222 VTAIL.n221 9.3005
R1597 VTAIL.n241 VTAIL.n240 9.3005
R1598 VTAIL.n243 VTAIL.n242 9.3005
R1599 VTAIL.n218 VTAIL.n217 9.3005
R1600 VTAIL.n249 VTAIL.n248 9.3005
R1601 VTAIL.n190 VTAIL.n189 9.3005
R1602 VTAIL.n197 VTAIL.n196 9.3005
R1603 VTAIL.n199 VTAIL.n198 9.3005
R1604 VTAIL.n186 VTAIL.n185 9.3005
R1605 VTAIL.n205 VTAIL.n204 9.3005
R1606 VTAIL.n207 VTAIL.n206 9.3005
R1607 VTAIL.n182 VTAIL.n181 9.3005
R1608 VTAIL.n213 VTAIL.n212 9.3005
R1609 VTAIL.n154 VTAIL.n153 9.3005
R1610 VTAIL.n161 VTAIL.n160 9.3005
R1611 VTAIL.n163 VTAIL.n162 9.3005
R1612 VTAIL.n150 VTAIL.n149 9.3005
R1613 VTAIL.n169 VTAIL.n168 9.3005
R1614 VTAIL.n171 VTAIL.n170 9.3005
R1615 VTAIL.n146 VTAIL.n145 9.3005
R1616 VTAIL.n177 VTAIL.n176 9.3005
R1617 VTAIL.n118 VTAIL.n117 9.3005
R1618 VTAIL.n125 VTAIL.n124 9.3005
R1619 VTAIL.n127 VTAIL.n126 9.3005
R1620 VTAIL.n114 VTAIL.n113 9.3005
R1621 VTAIL.n133 VTAIL.n132 9.3005
R1622 VTAIL.n135 VTAIL.n134 9.3005
R1623 VTAIL.n110 VTAIL.n109 9.3005
R1624 VTAIL.n141 VTAIL.n140 9.3005
R1625 VTAIL.n271 VTAIL.n260 8.92171
R1626 VTAIL.n19 VTAIL.n8 8.92171
R1627 VTAIL.n55 VTAIL.n44 8.92171
R1628 VTAIL.n91 VTAIL.n80 8.92171
R1629 VTAIL.n235 VTAIL.n224 8.92171
R1630 VTAIL.n199 VTAIL.n188 8.92171
R1631 VTAIL.n163 VTAIL.n152 8.92171
R1632 VTAIL.n127 VTAIL.n116 8.92171
R1633 VTAIL.n286 VTAIL.n252 8.2187
R1634 VTAIL.n34 VTAIL.n0 8.2187
R1635 VTAIL.n70 VTAIL.n36 8.2187
R1636 VTAIL.n106 VTAIL.n72 8.2187
R1637 VTAIL.n250 VTAIL.n216 8.2187
R1638 VTAIL.n214 VTAIL.n180 8.2187
R1639 VTAIL.n178 VTAIL.n144 8.2187
R1640 VTAIL.n142 VTAIL.n108 8.2187
R1641 VTAIL.n268 VTAIL.n267 8.14595
R1642 VTAIL.n16 VTAIL.n15 8.14595
R1643 VTAIL.n52 VTAIL.n51 8.14595
R1644 VTAIL.n88 VTAIL.n87 8.14595
R1645 VTAIL.n232 VTAIL.n231 8.14595
R1646 VTAIL.n196 VTAIL.n195 8.14595
R1647 VTAIL.n160 VTAIL.n159 8.14595
R1648 VTAIL.n124 VTAIL.n123 8.14595
R1649 VTAIL.n264 VTAIL.n262 7.3702
R1650 VTAIL.n12 VTAIL.n10 7.3702
R1651 VTAIL.n48 VTAIL.n46 7.3702
R1652 VTAIL.n84 VTAIL.n82 7.3702
R1653 VTAIL.n228 VTAIL.n226 7.3702
R1654 VTAIL.n192 VTAIL.n190 7.3702
R1655 VTAIL.n156 VTAIL.n154 7.3702
R1656 VTAIL.n120 VTAIL.n118 7.3702
R1657 VTAIL.n267 VTAIL.n262 5.81868
R1658 VTAIL.n15 VTAIL.n10 5.81868
R1659 VTAIL.n51 VTAIL.n46 5.81868
R1660 VTAIL.n87 VTAIL.n82 5.81868
R1661 VTAIL.n231 VTAIL.n226 5.81868
R1662 VTAIL.n195 VTAIL.n190 5.81868
R1663 VTAIL.n159 VTAIL.n154 5.81868
R1664 VTAIL.n123 VTAIL.n118 5.81868
R1665 VTAIL.n284 VTAIL.n252 5.3904
R1666 VTAIL.n32 VTAIL.n0 5.3904
R1667 VTAIL.n68 VTAIL.n36 5.3904
R1668 VTAIL.n104 VTAIL.n72 5.3904
R1669 VTAIL.n248 VTAIL.n216 5.3904
R1670 VTAIL.n212 VTAIL.n180 5.3904
R1671 VTAIL.n176 VTAIL.n144 5.3904
R1672 VTAIL.n140 VTAIL.n108 5.3904
R1673 VTAIL.n268 VTAIL.n260 5.04292
R1674 VTAIL.n16 VTAIL.n8 5.04292
R1675 VTAIL.n52 VTAIL.n44 5.04292
R1676 VTAIL.n88 VTAIL.n80 5.04292
R1677 VTAIL.n232 VTAIL.n224 5.04292
R1678 VTAIL.n196 VTAIL.n188 5.04292
R1679 VTAIL.n160 VTAIL.n152 5.04292
R1680 VTAIL.n124 VTAIL.n116 5.04292
R1681 VTAIL.n272 VTAIL.n271 4.26717
R1682 VTAIL.n20 VTAIL.n19 4.26717
R1683 VTAIL.n56 VTAIL.n55 4.26717
R1684 VTAIL.n92 VTAIL.n91 4.26717
R1685 VTAIL.n236 VTAIL.n235 4.26717
R1686 VTAIL.n200 VTAIL.n199 4.26717
R1687 VTAIL.n164 VTAIL.n163 4.26717
R1688 VTAIL.n128 VTAIL.n127 4.26717
R1689 VTAIL.n275 VTAIL.n258 3.49141
R1690 VTAIL.n23 VTAIL.n6 3.49141
R1691 VTAIL.n59 VTAIL.n42 3.49141
R1692 VTAIL.n95 VTAIL.n78 3.49141
R1693 VTAIL.n239 VTAIL.n222 3.49141
R1694 VTAIL.n203 VTAIL.n186 3.49141
R1695 VTAIL.n167 VTAIL.n150 3.49141
R1696 VTAIL.n131 VTAIL.n114 3.49141
R1697 VTAIL.n179 VTAIL.n143 3.32809
R1698 VTAIL.n251 VTAIL.n215 3.32809
R1699 VTAIL.n107 VTAIL.n71 3.32809
R1700 VTAIL.n263 VTAIL.n261 2.84305
R1701 VTAIL.n11 VTAIL.n9 2.84305
R1702 VTAIL.n47 VTAIL.n45 2.84305
R1703 VTAIL.n83 VTAIL.n81 2.84305
R1704 VTAIL.n227 VTAIL.n225 2.84305
R1705 VTAIL.n191 VTAIL.n189 2.84305
R1706 VTAIL.n155 VTAIL.n153 2.84305
R1707 VTAIL.n119 VTAIL.n117 2.84305
R1708 VTAIL.n276 VTAIL.n256 2.71565
R1709 VTAIL.n24 VTAIL.n4 2.71565
R1710 VTAIL.n60 VTAIL.n40 2.71565
R1711 VTAIL.n96 VTAIL.n76 2.71565
R1712 VTAIL.n240 VTAIL.n220 2.71565
R1713 VTAIL.n204 VTAIL.n184 2.71565
R1714 VTAIL.n168 VTAIL.n148 2.71565
R1715 VTAIL.n132 VTAIL.n112 2.71565
R1716 VTAIL.n280 VTAIL.n279 1.93989
R1717 VTAIL.n28 VTAIL.n27 1.93989
R1718 VTAIL.n64 VTAIL.n63 1.93989
R1719 VTAIL.n100 VTAIL.n99 1.93989
R1720 VTAIL.n244 VTAIL.n243 1.93989
R1721 VTAIL.n208 VTAIL.n207 1.93989
R1722 VTAIL.n172 VTAIL.n171 1.93989
R1723 VTAIL.n136 VTAIL.n135 1.93989
R1724 VTAIL VTAIL.n35 1.72248
R1725 VTAIL VTAIL.n287 1.6061
R1726 VTAIL.n283 VTAIL.n254 1.16414
R1727 VTAIL.n31 VTAIL.n2 1.16414
R1728 VTAIL.n67 VTAIL.n38 1.16414
R1729 VTAIL.n103 VTAIL.n74 1.16414
R1730 VTAIL.n247 VTAIL.n218 1.16414
R1731 VTAIL.n211 VTAIL.n182 1.16414
R1732 VTAIL.n175 VTAIL.n146 1.16414
R1733 VTAIL.n139 VTAIL.n110 1.16414
R1734 VTAIL.n215 VTAIL.n179 0.470328
R1735 VTAIL.n71 VTAIL.n35 0.470328
R1736 VTAIL.n269 VTAIL.n261 0.155672
R1737 VTAIL.n270 VTAIL.n269 0.155672
R1738 VTAIL.n270 VTAIL.n257 0.155672
R1739 VTAIL.n277 VTAIL.n257 0.155672
R1740 VTAIL.n278 VTAIL.n277 0.155672
R1741 VTAIL.n278 VTAIL.n253 0.155672
R1742 VTAIL.n285 VTAIL.n253 0.155672
R1743 VTAIL.n17 VTAIL.n9 0.155672
R1744 VTAIL.n18 VTAIL.n17 0.155672
R1745 VTAIL.n18 VTAIL.n5 0.155672
R1746 VTAIL.n25 VTAIL.n5 0.155672
R1747 VTAIL.n26 VTAIL.n25 0.155672
R1748 VTAIL.n26 VTAIL.n1 0.155672
R1749 VTAIL.n33 VTAIL.n1 0.155672
R1750 VTAIL.n53 VTAIL.n45 0.155672
R1751 VTAIL.n54 VTAIL.n53 0.155672
R1752 VTAIL.n54 VTAIL.n41 0.155672
R1753 VTAIL.n61 VTAIL.n41 0.155672
R1754 VTAIL.n62 VTAIL.n61 0.155672
R1755 VTAIL.n62 VTAIL.n37 0.155672
R1756 VTAIL.n69 VTAIL.n37 0.155672
R1757 VTAIL.n89 VTAIL.n81 0.155672
R1758 VTAIL.n90 VTAIL.n89 0.155672
R1759 VTAIL.n90 VTAIL.n77 0.155672
R1760 VTAIL.n97 VTAIL.n77 0.155672
R1761 VTAIL.n98 VTAIL.n97 0.155672
R1762 VTAIL.n98 VTAIL.n73 0.155672
R1763 VTAIL.n105 VTAIL.n73 0.155672
R1764 VTAIL.n249 VTAIL.n217 0.155672
R1765 VTAIL.n242 VTAIL.n217 0.155672
R1766 VTAIL.n242 VTAIL.n241 0.155672
R1767 VTAIL.n241 VTAIL.n221 0.155672
R1768 VTAIL.n234 VTAIL.n221 0.155672
R1769 VTAIL.n234 VTAIL.n233 0.155672
R1770 VTAIL.n233 VTAIL.n225 0.155672
R1771 VTAIL.n213 VTAIL.n181 0.155672
R1772 VTAIL.n206 VTAIL.n181 0.155672
R1773 VTAIL.n206 VTAIL.n205 0.155672
R1774 VTAIL.n205 VTAIL.n185 0.155672
R1775 VTAIL.n198 VTAIL.n185 0.155672
R1776 VTAIL.n198 VTAIL.n197 0.155672
R1777 VTAIL.n197 VTAIL.n189 0.155672
R1778 VTAIL.n177 VTAIL.n145 0.155672
R1779 VTAIL.n170 VTAIL.n145 0.155672
R1780 VTAIL.n170 VTAIL.n169 0.155672
R1781 VTAIL.n169 VTAIL.n149 0.155672
R1782 VTAIL.n162 VTAIL.n149 0.155672
R1783 VTAIL.n162 VTAIL.n161 0.155672
R1784 VTAIL.n161 VTAIL.n153 0.155672
R1785 VTAIL.n141 VTAIL.n109 0.155672
R1786 VTAIL.n134 VTAIL.n109 0.155672
R1787 VTAIL.n134 VTAIL.n133 0.155672
R1788 VTAIL.n133 VTAIL.n113 0.155672
R1789 VTAIL.n126 VTAIL.n113 0.155672
R1790 VTAIL.n126 VTAIL.n125 0.155672
R1791 VTAIL.n125 VTAIL.n117 0.155672
R1792 VDD1 VDD1.n1 109.62
R1793 VDD1 VDD1.n0 69.1536
R1794 VDD1.n0 VDD1.t2 2.70912
R1795 VDD1.n0 VDD1.t3 2.70912
R1796 VDD1.n1 VDD1.t0 2.70912
R1797 VDD1.n1 VDD1.t1 2.70912
R1798 VN.n1 VN.t2 84.4854
R1799 VN.n0 VN.t1 84.4854
R1800 VN.n0 VN.t3 83.2583
R1801 VN.n1 VN.t0 83.2583
R1802 VN VN.n1 47.992
R1803 VN VN.n0 2.17003
R1804 VDD2.n2 VDD2.n0 109.094
R1805 VDD2.n2 VDD2.n1 69.0954
R1806 VDD2.n1 VDD2.t3 2.70912
R1807 VDD2.n1 VDD2.t1 2.70912
R1808 VDD2.n0 VDD2.t2 2.70912
R1809 VDD2.n0 VDD2.t0 2.70912
R1810 VDD2 VDD2.n2 0.0586897
C0 VTAIL VN 3.43646f
C1 VDD2 VN 3.15947f
C2 VP VN 5.99373f
C3 VDD1 VN 0.149991f
C4 VDD2 VTAIL 4.71186f
C5 VTAIL VP 3.45057f
C6 VDD1 VTAIL 4.65142f
C7 VDD2 VP 0.453634f
C8 VDD2 VDD1 1.24939f
C9 VDD1 VP 3.46214f
C10 VDD2 B 3.94455f
C11 VDD1 B 8.06793f
C12 VTAIL B 7.739665f
C13 VN B 12.18721f
C14 VP B 10.59844f
C15 VDD2.t2 B 0.161823f
C16 VDD2.t0 B 0.161823f
C17 VDD2.n0 B 1.93172f
C18 VDD2.t3 B 0.161823f
C19 VDD2.t1 B 0.161823f
C20 VDD2.n1 B 1.39169f
C21 VDD2.n2 B 3.6229f
C22 VN.t3 B 1.8835f
C23 VN.t1 B 1.89407f
C24 VN.n0 B 1.11447f
C25 VN.t2 B 1.89407f
C26 VN.t0 B 1.8835f
C27 VN.n1 B 2.45018f
C28 VDD1.t2 B 0.165797f
C29 VDD1.t3 B 0.165797f
C30 VDD1.n0 B 1.42633f
C31 VDD1.t0 B 0.165797f
C32 VDD1.t1 B 0.165797f
C33 VDD1.n1 B 2.00485f
C34 VTAIL.n0 B 0.027298f
C35 VTAIL.n1 B 0.019278f
C36 VTAIL.n2 B 0.010359f
C37 VTAIL.n3 B 0.024485f
C38 VTAIL.n4 B 0.010969f
C39 VTAIL.n5 B 0.019278f
C40 VTAIL.n6 B 0.010359f
C41 VTAIL.n7 B 0.024485f
C42 VTAIL.n8 B 0.010969f
C43 VTAIL.n9 B 0.570311f
C44 VTAIL.n10 B 0.010359f
C45 VTAIL.t0 B 0.040898f
C46 VTAIL.n11 B 0.104336f
C47 VTAIL.n12 B 0.017309f
C48 VTAIL.n13 B 0.018364f
C49 VTAIL.n14 B 0.024485f
C50 VTAIL.n15 B 0.010969f
C51 VTAIL.n16 B 0.010359f
C52 VTAIL.n17 B 0.019278f
C53 VTAIL.n18 B 0.019278f
C54 VTAIL.n19 B 0.010359f
C55 VTAIL.n20 B 0.010969f
C56 VTAIL.n21 B 0.024485f
C57 VTAIL.n22 B 0.024485f
C58 VTAIL.n23 B 0.010969f
C59 VTAIL.n24 B 0.010359f
C60 VTAIL.n25 B 0.019278f
C61 VTAIL.n26 B 0.019278f
C62 VTAIL.n27 B 0.010359f
C63 VTAIL.n28 B 0.010969f
C64 VTAIL.n29 B 0.024485f
C65 VTAIL.n30 B 0.051045f
C66 VTAIL.n31 B 0.010969f
C67 VTAIL.n32 B 0.020256f
C68 VTAIL.n33 B 0.050618f
C69 VTAIL.n34 B 0.053982f
C70 VTAIL.n35 B 0.156046f
C71 VTAIL.n36 B 0.027298f
C72 VTAIL.n37 B 0.019278f
C73 VTAIL.n38 B 0.010359f
C74 VTAIL.n39 B 0.024485f
C75 VTAIL.n40 B 0.010969f
C76 VTAIL.n41 B 0.019278f
C77 VTAIL.n42 B 0.010359f
C78 VTAIL.n43 B 0.024485f
C79 VTAIL.n44 B 0.010969f
C80 VTAIL.n45 B 0.570311f
C81 VTAIL.n46 B 0.010359f
C82 VTAIL.t5 B 0.040898f
C83 VTAIL.n47 B 0.104336f
C84 VTAIL.n48 B 0.017309f
C85 VTAIL.n49 B 0.018364f
C86 VTAIL.n50 B 0.024485f
C87 VTAIL.n51 B 0.010969f
C88 VTAIL.n52 B 0.010359f
C89 VTAIL.n53 B 0.019278f
C90 VTAIL.n54 B 0.019278f
C91 VTAIL.n55 B 0.010359f
C92 VTAIL.n56 B 0.010969f
C93 VTAIL.n57 B 0.024485f
C94 VTAIL.n58 B 0.024485f
C95 VTAIL.n59 B 0.010969f
C96 VTAIL.n60 B 0.010359f
C97 VTAIL.n61 B 0.019278f
C98 VTAIL.n62 B 0.019278f
C99 VTAIL.n63 B 0.010359f
C100 VTAIL.n64 B 0.010969f
C101 VTAIL.n65 B 0.024485f
C102 VTAIL.n66 B 0.051045f
C103 VTAIL.n67 B 0.010969f
C104 VTAIL.n68 B 0.020256f
C105 VTAIL.n69 B 0.050618f
C106 VTAIL.n70 B 0.053982f
C107 VTAIL.n71 B 0.255783f
C108 VTAIL.n72 B 0.027298f
C109 VTAIL.n73 B 0.019278f
C110 VTAIL.n74 B 0.010359f
C111 VTAIL.n75 B 0.024485f
C112 VTAIL.n76 B 0.010969f
C113 VTAIL.n77 B 0.019278f
C114 VTAIL.n78 B 0.010359f
C115 VTAIL.n79 B 0.024485f
C116 VTAIL.n80 B 0.010969f
C117 VTAIL.n81 B 0.570311f
C118 VTAIL.n82 B 0.010359f
C119 VTAIL.t4 B 0.040898f
C120 VTAIL.n83 B 0.104336f
C121 VTAIL.n84 B 0.017309f
C122 VTAIL.n85 B 0.018364f
C123 VTAIL.n86 B 0.024485f
C124 VTAIL.n87 B 0.010969f
C125 VTAIL.n88 B 0.010359f
C126 VTAIL.n89 B 0.019278f
C127 VTAIL.n90 B 0.019278f
C128 VTAIL.n91 B 0.010359f
C129 VTAIL.n92 B 0.010969f
C130 VTAIL.n93 B 0.024485f
C131 VTAIL.n94 B 0.024485f
C132 VTAIL.n95 B 0.010969f
C133 VTAIL.n96 B 0.010359f
C134 VTAIL.n97 B 0.019278f
C135 VTAIL.n98 B 0.019278f
C136 VTAIL.n99 B 0.010359f
C137 VTAIL.n100 B 0.010969f
C138 VTAIL.n101 B 0.024485f
C139 VTAIL.n102 B 0.051045f
C140 VTAIL.n103 B 0.010969f
C141 VTAIL.n104 B 0.020256f
C142 VTAIL.n105 B 0.050618f
C143 VTAIL.n106 B 0.053982f
C144 VTAIL.n107 B 1.08663f
C145 VTAIL.n108 B 0.027298f
C146 VTAIL.n109 B 0.019278f
C147 VTAIL.n110 B 0.010359f
C148 VTAIL.n111 B 0.024485f
C149 VTAIL.n112 B 0.010969f
C150 VTAIL.n113 B 0.019278f
C151 VTAIL.n114 B 0.010359f
C152 VTAIL.n115 B 0.024485f
C153 VTAIL.n116 B 0.010969f
C154 VTAIL.n117 B 0.570311f
C155 VTAIL.n118 B 0.010359f
C156 VTAIL.t3 B 0.040899f
C157 VTAIL.n119 B 0.104336f
C158 VTAIL.n120 B 0.017309f
C159 VTAIL.n121 B 0.018364f
C160 VTAIL.n122 B 0.024485f
C161 VTAIL.n123 B 0.010969f
C162 VTAIL.n124 B 0.010359f
C163 VTAIL.n125 B 0.019278f
C164 VTAIL.n126 B 0.019278f
C165 VTAIL.n127 B 0.010359f
C166 VTAIL.n128 B 0.010969f
C167 VTAIL.n129 B 0.024485f
C168 VTAIL.n130 B 0.024485f
C169 VTAIL.n131 B 0.010969f
C170 VTAIL.n132 B 0.010359f
C171 VTAIL.n133 B 0.019278f
C172 VTAIL.n134 B 0.019278f
C173 VTAIL.n135 B 0.010359f
C174 VTAIL.n136 B 0.010969f
C175 VTAIL.n137 B 0.024485f
C176 VTAIL.n138 B 0.051045f
C177 VTAIL.n139 B 0.010969f
C178 VTAIL.n140 B 0.020256f
C179 VTAIL.n141 B 0.050618f
C180 VTAIL.n142 B 0.053982f
C181 VTAIL.n143 B 1.08663f
C182 VTAIL.n144 B 0.027298f
C183 VTAIL.n145 B 0.019278f
C184 VTAIL.n146 B 0.010359f
C185 VTAIL.n147 B 0.024485f
C186 VTAIL.n148 B 0.010969f
C187 VTAIL.n149 B 0.019278f
C188 VTAIL.n150 B 0.010359f
C189 VTAIL.n151 B 0.024485f
C190 VTAIL.n152 B 0.010969f
C191 VTAIL.n153 B 0.570311f
C192 VTAIL.n154 B 0.010359f
C193 VTAIL.t1 B 0.040899f
C194 VTAIL.n155 B 0.104336f
C195 VTAIL.n156 B 0.017309f
C196 VTAIL.n157 B 0.018364f
C197 VTAIL.n158 B 0.024485f
C198 VTAIL.n159 B 0.010969f
C199 VTAIL.n160 B 0.010359f
C200 VTAIL.n161 B 0.019278f
C201 VTAIL.n162 B 0.019278f
C202 VTAIL.n163 B 0.010359f
C203 VTAIL.n164 B 0.010969f
C204 VTAIL.n165 B 0.024485f
C205 VTAIL.n166 B 0.024485f
C206 VTAIL.n167 B 0.010969f
C207 VTAIL.n168 B 0.010359f
C208 VTAIL.n169 B 0.019278f
C209 VTAIL.n170 B 0.019278f
C210 VTAIL.n171 B 0.010359f
C211 VTAIL.n172 B 0.010969f
C212 VTAIL.n173 B 0.024485f
C213 VTAIL.n174 B 0.051045f
C214 VTAIL.n175 B 0.010969f
C215 VTAIL.n176 B 0.020256f
C216 VTAIL.n177 B 0.050618f
C217 VTAIL.n178 B 0.053982f
C218 VTAIL.n179 B 0.255783f
C219 VTAIL.n180 B 0.027298f
C220 VTAIL.n181 B 0.019278f
C221 VTAIL.n182 B 0.010359f
C222 VTAIL.n183 B 0.024485f
C223 VTAIL.n184 B 0.010969f
C224 VTAIL.n185 B 0.019278f
C225 VTAIL.n186 B 0.010359f
C226 VTAIL.n187 B 0.024485f
C227 VTAIL.n188 B 0.010969f
C228 VTAIL.n189 B 0.570311f
C229 VTAIL.n190 B 0.010359f
C230 VTAIL.t7 B 0.040899f
C231 VTAIL.n191 B 0.104336f
C232 VTAIL.n192 B 0.017309f
C233 VTAIL.n193 B 0.018364f
C234 VTAIL.n194 B 0.024485f
C235 VTAIL.n195 B 0.010969f
C236 VTAIL.n196 B 0.010359f
C237 VTAIL.n197 B 0.019278f
C238 VTAIL.n198 B 0.019278f
C239 VTAIL.n199 B 0.010359f
C240 VTAIL.n200 B 0.010969f
C241 VTAIL.n201 B 0.024485f
C242 VTAIL.n202 B 0.024485f
C243 VTAIL.n203 B 0.010969f
C244 VTAIL.n204 B 0.010359f
C245 VTAIL.n205 B 0.019278f
C246 VTAIL.n206 B 0.019278f
C247 VTAIL.n207 B 0.010359f
C248 VTAIL.n208 B 0.010969f
C249 VTAIL.n209 B 0.024485f
C250 VTAIL.n210 B 0.051045f
C251 VTAIL.n211 B 0.010969f
C252 VTAIL.n212 B 0.020256f
C253 VTAIL.n213 B 0.050618f
C254 VTAIL.n214 B 0.053982f
C255 VTAIL.n215 B 0.255783f
C256 VTAIL.n216 B 0.027298f
C257 VTAIL.n217 B 0.019278f
C258 VTAIL.n218 B 0.010359f
C259 VTAIL.n219 B 0.024485f
C260 VTAIL.n220 B 0.010969f
C261 VTAIL.n221 B 0.019278f
C262 VTAIL.n222 B 0.010359f
C263 VTAIL.n223 B 0.024485f
C264 VTAIL.n224 B 0.010969f
C265 VTAIL.n225 B 0.570311f
C266 VTAIL.n226 B 0.010359f
C267 VTAIL.t6 B 0.040899f
C268 VTAIL.n227 B 0.104336f
C269 VTAIL.n228 B 0.017309f
C270 VTAIL.n229 B 0.018364f
C271 VTAIL.n230 B 0.024485f
C272 VTAIL.n231 B 0.010969f
C273 VTAIL.n232 B 0.010359f
C274 VTAIL.n233 B 0.019278f
C275 VTAIL.n234 B 0.019278f
C276 VTAIL.n235 B 0.010359f
C277 VTAIL.n236 B 0.010969f
C278 VTAIL.n237 B 0.024485f
C279 VTAIL.n238 B 0.024485f
C280 VTAIL.n239 B 0.010969f
C281 VTAIL.n240 B 0.010359f
C282 VTAIL.n241 B 0.019278f
C283 VTAIL.n242 B 0.019278f
C284 VTAIL.n243 B 0.010359f
C285 VTAIL.n244 B 0.010969f
C286 VTAIL.n245 B 0.024485f
C287 VTAIL.n246 B 0.051045f
C288 VTAIL.n247 B 0.010969f
C289 VTAIL.n248 B 0.020256f
C290 VTAIL.n249 B 0.050618f
C291 VTAIL.n250 B 0.053982f
C292 VTAIL.n251 B 1.08663f
C293 VTAIL.n252 B 0.027298f
C294 VTAIL.n253 B 0.019278f
C295 VTAIL.n254 B 0.010359f
C296 VTAIL.n255 B 0.024485f
C297 VTAIL.n256 B 0.010969f
C298 VTAIL.n257 B 0.019278f
C299 VTAIL.n258 B 0.010359f
C300 VTAIL.n259 B 0.024485f
C301 VTAIL.n260 B 0.010969f
C302 VTAIL.n261 B 0.570311f
C303 VTAIL.n262 B 0.010359f
C304 VTAIL.t2 B 0.040898f
C305 VTAIL.n263 B 0.104336f
C306 VTAIL.n264 B 0.017309f
C307 VTAIL.n265 B 0.018364f
C308 VTAIL.n266 B 0.024485f
C309 VTAIL.n267 B 0.010969f
C310 VTAIL.n268 B 0.010359f
C311 VTAIL.n269 B 0.019278f
C312 VTAIL.n270 B 0.019278f
C313 VTAIL.n271 B 0.010359f
C314 VTAIL.n272 B 0.010969f
C315 VTAIL.n273 B 0.024485f
C316 VTAIL.n274 B 0.024485f
C317 VTAIL.n275 B 0.010969f
C318 VTAIL.n276 B 0.010359f
C319 VTAIL.n277 B 0.019278f
C320 VTAIL.n278 B 0.019278f
C321 VTAIL.n279 B 0.010359f
C322 VTAIL.n280 B 0.010969f
C323 VTAIL.n281 B 0.024485f
C324 VTAIL.n282 B 0.051045f
C325 VTAIL.n283 B 0.010969f
C326 VTAIL.n284 B 0.020256f
C327 VTAIL.n285 B 0.050618f
C328 VTAIL.n286 B 0.053982f
C329 VTAIL.n287 B 0.97966f
C330 VP.t2 B 1.6397f
C331 VP.n0 B 0.685276f
C332 VP.n1 B 0.023757f
C333 VP.n2 B 0.034682f
C334 VP.n3 B 0.023757f
C335 VP.n4 B 0.030287f
C336 VP.t1 B 1.95921f
C337 VP.t0 B 1.94829f
C338 VP.n5 B 2.52464f
C339 VP.t3 B 1.6397f
C340 VP.n6 B 0.685276f
C341 VP.n7 B 1.27794f
C342 VP.n8 B 0.038344f
C343 VP.n9 B 0.023757f
C344 VP.n10 B 0.044278f
C345 VP.n11 B 0.044278f
C346 VP.n12 B 0.034682f
C347 VP.n13 B 0.023757f
C348 VP.n14 B 0.023757f
C349 VP.n15 B 0.023757f
C350 VP.n16 B 0.044278f
C351 VP.n17 B 0.044278f
C352 VP.n18 B 0.030287f
C353 VP.n19 B 0.038344f
C354 VP.n20 B 0.06514f
.ends

