* NGSPICE file created from diff_pair_sample_1163.ext - technology: sky130A

.subckt diff_pair_sample_1163 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.0771 pd=16.56 as=3.0771 ps=16.56 w=7.89 l=2.64
X1 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.0771 pd=16.56 as=3.0771 ps=16.56 w=7.89 l=2.64
X2 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=3.0771 pd=16.56 as=0 ps=0 w=7.89 l=2.64
X3 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=3.0771 pd=16.56 as=0 ps=0 w=7.89 l=2.64
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.0771 pd=16.56 as=0 ps=0 w=7.89 l=2.64
X5 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=3.0771 pd=16.56 as=3.0771 ps=16.56 w=7.89 l=2.64
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.0771 pd=16.56 as=0 ps=0 w=7.89 l=2.64
X7 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.0771 pd=16.56 as=3.0771 ps=16.56 w=7.89 l=2.64
R0 VN VN.t1 154.774
R1 VN VN.t0 113.553
R2 VTAIL.n162 VTAIL.n126 289.615
R3 VTAIL.n36 VTAIL.n0 289.615
R4 VTAIL.n120 VTAIL.n84 289.615
R5 VTAIL.n78 VTAIL.n42 289.615
R6 VTAIL.n138 VTAIL.n137 185
R7 VTAIL.n143 VTAIL.n142 185
R8 VTAIL.n145 VTAIL.n144 185
R9 VTAIL.n134 VTAIL.n133 185
R10 VTAIL.n151 VTAIL.n150 185
R11 VTAIL.n153 VTAIL.n152 185
R12 VTAIL.n130 VTAIL.n129 185
R13 VTAIL.n160 VTAIL.n159 185
R14 VTAIL.n161 VTAIL.n128 185
R15 VTAIL.n163 VTAIL.n162 185
R16 VTAIL.n12 VTAIL.n11 185
R17 VTAIL.n17 VTAIL.n16 185
R18 VTAIL.n19 VTAIL.n18 185
R19 VTAIL.n8 VTAIL.n7 185
R20 VTAIL.n25 VTAIL.n24 185
R21 VTAIL.n27 VTAIL.n26 185
R22 VTAIL.n4 VTAIL.n3 185
R23 VTAIL.n34 VTAIL.n33 185
R24 VTAIL.n35 VTAIL.n2 185
R25 VTAIL.n37 VTAIL.n36 185
R26 VTAIL.n121 VTAIL.n120 185
R27 VTAIL.n119 VTAIL.n86 185
R28 VTAIL.n118 VTAIL.n117 185
R29 VTAIL.n89 VTAIL.n87 185
R30 VTAIL.n112 VTAIL.n111 185
R31 VTAIL.n110 VTAIL.n109 185
R32 VTAIL.n93 VTAIL.n92 185
R33 VTAIL.n104 VTAIL.n103 185
R34 VTAIL.n102 VTAIL.n101 185
R35 VTAIL.n97 VTAIL.n96 185
R36 VTAIL.n79 VTAIL.n78 185
R37 VTAIL.n77 VTAIL.n44 185
R38 VTAIL.n76 VTAIL.n75 185
R39 VTAIL.n47 VTAIL.n45 185
R40 VTAIL.n70 VTAIL.n69 185
R41 VTAIL.n68 VTAIL.n67 185
R42 VTAIL.n51 VTAIL.n50 185
R43 VTAIL.n62 VTAIL.n61 185
R44 VTAIL.n60 VTAIL.n59 185
R45 VTAIL.n55 VTAIL.n54 185
R46 VTAIL.n139 VTAIL.t3 149.524
R47 VTAIL.n13 VTAIL.t0 149.524
R48 VTAIL.n98 VTAIL.t1 149.524
R49 VTAIL.n56 VTAIL.t2 149.524
R50 VTAIL.n143 VTAIL.n137 104.615
R51 VTAIL.n144 VTAIL.n143 104.615
R52 VTAIL.n144 VTAIL.n133 104.615
R53 VTAIL.n151 VTAIL.n133 104.615
R54 VTAIL.n152 VTAIL.n151 104.615
R55 VTAIL.n152 VTAIL.n129 104.615
R56 VTAIL.n160 VTAIL.n129 104.615
R57 VTAIL.n161 VTAIL.n160 104.615
R58 VTAIL.n162 VTAIL.n161 104.615
R59 VTAIL.n17 VTAIL.n11 104.615
R60 VTAIL.n18 VTAIL.n17 104.615
R61 VTAIL.n18 VTAIL.n7 104.615
R62 VTAIL.n25 VTAIL.n7 104.615
R63 VTAIL.n26 VTAIL.n25 104.615
R64 VTAIL.n26 VTAIL.n3 104.615
R65 VTAIL.n34 VTAIL.n3 104.615
R66 VTAIL.n35 VTAIL.n34 104.615
R67 VTAIL.n36 VTAIL.n35 104.615
R68 VTAIL.n120 VTAIL.n119 104.615
R69 VTAIL.n119 VTAIL.n118 104.615
R70 VTAIL.n118 VTAIL.n87 104.615
R71 VTAIL.n111 VTAIL.n87 104.615
R72 VTAIL.n111 VTAIL.n110 104.615
R73 VTAIL.n110 VTAIL.n92 104.615
R74 VTAIL.n103 VTAIL.n92 104.615
R75 VTAIL.n103 VTAIL.n102 104.615
R76 VTAIL.n102 VTAIL.n96 104.615
R77 VTAIL.n78 VTAIL.n77 104.615
R78 VTAIL.n77 VTAIL.n76 104.615
R79 VTAIL.n76 VTAIL.n45 104.615
R80 VTAIL.n69 VTAIL.n45 104.615
R81 VTAIL.n69 VTAIL.n68 104.615
R82 VTAIL.n68 VTAIL.n50 104.615
R83 VTAIL.n61 VTAIL.n50 104.615
R84 VTAIL.n61 VTAIL.n60 104.615
R85 VTAIL.n60 VTAIL.n54 104.615
R86 VTAIL.t3 VTAIL.n137 52.3082
R87 VTAIL.t0 VTAIL.n11 52.3082
R88 VTAIL.t1 VTAIL.n96 52.3082
R89 VTAIL.t2 VTAIL.n54 52.3082
R90 VTAIL.n167 VTAIL.n166 33.9308
R91 VTAIL.n41 VTAIL.n40 33.9308
R92 VTAIL.n125 VTAIL.n124 33.9308
R93 VTAIL.n83 VTAIL.n82 33.9308
R94 VTAIL.n83 VTAIL.n41 24.2893
R95 VTAIL.n167 VTAIL.n125 21.7289
R96 VTAIL.n163 VTAIL.n128 13.1884
R97 VTAIL.n37 VTAIL.n2 13.1884
R98 VTAIL.n121 VTAIL.n86 13.1884
R99 VTAIL.n79 VTAIL.n44 13.1884
R100 VTAIL.n159 VTAIL.n158 12.8005
R101 VTAIL.n164 VTAIL.n126 12.8005
R102 VTAIL.n33 VTAIL.n32 12.8005
R103 VTAIL.n38 VTAIL.n0 12.8005
R104 VTAIL.n122 VTAIL.n84 12.8005
R105 VTAIL.n117 VTAIL.n88 12.8005
R106 VTAIL.n80 VTAIL.n42 12.8005
R107 VTAIL.n75 VTAIL.n46 12.8005
R108 VTAIL.n157 VTAIL.n130 12.0247
R109 VTAIL.n31 VTAIL.n4 12.0247
R110 VTAIL.n116 VTAIL.n89 12.0247
R111 VTAIL.n74 VTAIL.n47 12.0247
R112 VTAIL.n154 VTAIL.n153 11.249
R113 VTAIL.n28 VTAIL.n27 11.249
R114 VTAIL.n113 VTAIL.n112 11.249
R115 VTAIL.n71 VTAIL.n70 11.249
R116 VTAIL.n150 VTAIL.n132 10.4732
R117 VTAIL.n24 VTAIL.n6 10.4732
R118 VTAIL.n109 VTAIL.n91 10.4732
R119 VTAIL.n67 VTAIL.n49 10.4732
R120 VTAIL.n139 VTAIL.n138 10.2747
R121 VTAIL.n13 VTAIL.n12 10.2747
R122 VTAIL.n98 VTAIL.n97 10.2747
R123 VTAIL.n56 VTAIL.n55 10.2747
R124 VTAIL.n149 VTAIL.n134 9.69747
R125 VTAIL.n23 VTAIL.n8 9.69747
R126 VTAIL.n108 VTAIL.n93 9.69747
R127 VTAIL.n66 VTAIL.n51 9.69747
R128 VTAIL.n166 VTAIL.n165 9.45567
R129 VTAIL.n40 VTAIL.n39 9.45567
R130 VTAIL.n124 VTAIL.n123 9.45567
R131 VTAIL.n82 VTAIL.n81 9.45567
R132 VTAIL.n165 VTAIL.n164 9.3005
R133 VTAIL.n141 VTAIL.n140 9.3005
R134 VTAIL.n136 VTAIL.n135 9.3005
R135 VTAIL.n147 VTAIL.n146 9.3005
R136 VTAIL.n149 VTAIL.n148 9.3005
R137 VTAIL.n132 VTAIL.n131 9.3005
R138 VTAIL.n155 VTAIL.n154 9.3005
R139 VTAIL.n157 VTAIL.n156 9.3005
R140 VTAIL.n158 VTAIL.n127 9.3005
R141 VTAIL.n39 VTAIL.n38 9.3005
R142 VTAIL.n15 VTAIL.n14 9.3005
R143 VTAIL.n10 VTAIL.n9 9.3005
R144 VTAIL.n21 VTAIL.n20 9.3005
R145 VTAIL.n23 VTAIL.n22 9.3005
R146 VTAIL.n6 VTAIL.n5 9.3005
R147 VTAIL.n29 VTAIL.n28 9.3005
R148 VTAIL.n31 VTAIL.n30 9.3005
R149 VTAIL.n32 VTAIL.n1 9.3005
R150 VTAIL.n100 VTAIL.n99 9.3005
R151 VTAIL.n95 VTAIL.n94 9.3005
R152 VTAIL.n106 VTAIL.n105 9.3005
R153 VTAIL.n108 VTAIL.n107 9.3005
R154 VTAIL.n91 VTAIL.n90 9.3005
R155 VTAIL.n114 VTAIL.n113 9.3005
R156 VTAIL.n116 VTAIL.n115 9.3005
R157 VTAIL.n88 VTAIL.n85 9.3005
R158 VTAIL.n123 VTAIL.n122 9.3005
R159 VTAIL.n58 VTAIL.n57 9.3005
R160 VTAIL.n53 VTAIL.n52 9.3005
R161 VTAIL.n64 VTAIL.n63 9.3005
R162 VTAIL.n66 VTAIL.n65 9.3005
R163 VTAIL.n49 VTAIL.n48 9.3005
R164 VTAIL.n72 VTAIL.n71 9.3005
R165 VTAIL.n74 VTAIL.n73 9.3005
R166 VTAIL.n46 VTAIL.n43 9.3005
R167 VTAIL.n81 VTAIL.n80 9.3005
R168 VTAIL.n146 VTAIL.n145 8.92171
R169 VTAIL.n20 VTAIL.n19 8.92171
R170 VTAIL.n105 VTAIL.n104 8.92171
R171 VTAIL.n63 VTAIL.n62 8.92171
R172 VTAIL.n142 VTAIL.n136 8.14595
R173 VTAIL.n16 VTAIL.n10 8.14595
R174 VTAIL.n101 VTAIL.n95 8.14595
R175 VTAIL.n59 VTAIL.n53 8.14595
R176 VTAIL.n141 VTAIL.n138 7.3702
R177 VTAIL.n15 VTAIL.n12 7.3702
R178 VTAIL.n100 VTAIL.n97 7.3702
R179 VTAIL.n58 VTAIL.n55 7.3702
R180 VTAIL.n142 VTAIL.n141 5.81868
R181 VTAIL.n16 VTAIL.n15 5.81868
R182 VTAIL.n101 VTAIL.n100 5.81868
R183 VTAIL.n59 VTAIL.n58 5.81868
R184 VTAIL.n145 VTAIL.n136 5.04292
R185 VTAIL.n19 VTAIL.n10 5.04292
R186 VTAIL.n104 VTAIL.n95 5.04292
R187 VTAIL.n62 VTAIL.n53 5.04292
R188 VTAIL.n146 VTAIL.n134 4.26717
R189 VTAIL.n20 VTAIL.n8 4.26717
R190 VTAIL.n105 VTAIL.n93 4.26717
R191 VTAIL.n63 VTAIL.n51 4.26717
R192 VTAIL.n150 VTAIL.n149 3.49141
R193 VTAIL.n24 VTAIL.n23 3.49141
R194 VTAIL.n109 VTAIL.n108 3.49141
R195 VTAIL.n67 VTAIL.n66 3.49141
R196 VTAIL.n140 VTAIL.n139 2.84304
R197 VTAIL.n14 VTAIL.n13 2.84304
R198 VTAIL.n99 VTAIL.n98 2.84304
R199 VTAIL.n57 VTAIL.n56 2.84304
R200 VTAIL.n153 VTAIL.n132 2.71565
R201 VTAIL.n27 VTAIL.n6 2.71565
R202 VTAIL.n112 VTAIL.n91 2.71565
R203 VTAIL.n70 VTAIL.n49 2.71565
R204 VTAIL.n154 VTAIL.n130 1.93989
R205 VTAIL.n28 VTAIL.n4 1.93989
R206 VTAIL.n113 VTAIL.n89 1.93989
R207 VTAIL.n71 VTAIL.n47 1.93989
R208 VTAIL.n125 VTAIL.n83 1.7505
R209 VTAIL VTAIL.n41 1.1686
R210 VTAIL.n159 VTAIL.n157 1.16414
R211 VTAIL.n166 VTAIL.n126 1.16414
R212 VTAIL.n33 VTAIL.n31 1.16414
R213 VTAIL.n40 VTAIL.n0 1.16414
R214 VTAIL.n124 VTAIL.n84 1.16414
R215 VTAIL.n117 VTAIL.n116 1.16414
R216 VTAIL.n82 VTAIL.n42 1.16414
R217 VTAIL.n75 VTAIL.n74 1.16414
R218 VTAIL VTAIL.n167 0.582397
R219 VTAIL.n158 VTAIL.n128 0.388379
R220 VTAIL.n164 VTAIL.n163 0.388379
R221 VTAIL.n32 VTAIL.n2 0.388379
R222 VTAIL.n38 VTAIL.n37 0.388379
R223 VTAIL.n122 VTAIL.n121 0.388379
R224 VTAIL.n88 VTAIL.n86 0.388379
R225 VTAIL.n80 VTAIL.n79 0.388379
R226 VTAIL.n46 VTAIL.n44 0.388379
R227 VTAIL.n140 VTAIL.n135 0.155672
R228 VTAIL.n147 VTAIL.n135 0.155672
R229 VTAIL.n148 VTAIL.n147 0.155672
R230 VTAIL.n148 VTAIL.n131 0.155672
R231 VTAIL.n155 VTAIL.n131 0.155672
R232 VTAIL.n156 VTAIL.n155 0.155672
R233 VTAIL.n156 VTAIL.n127 0.155672
R234 VTAIL.n165 VTAIL.n127 0.155672
R235 VTAIL.n14 VTAIL.n9 0.155672
R236 VTAIL.n21 VTAIL.n9 0.155672
R237 VTAIL.n22 VTAIL.n21 0.155672
R238 VTAIL.n22 VTAIL.n5 0.155672
R239 VTAIL.n29 VTAIL.n5 0.155672
R240 VTAIL.n30 VTAIL.n29 0.155672
R241 VTAIL.n30 VTAIL.n1 0.155672
R242 VTAIL.n39 VTAIL.n1 0.155672
R243 VTAIL.n123 VTAIL.n85 0.155672
R244 VTAIL.n115 VTAIL.n85 0.155672
R245 VTAIL.n115 VTAIL.n114 0.155672
R246 VTAIL.n114 VTAIL.n90 0.155672
R247 VTAIL.n107 VTAIL.n90 0.155672
R248 VTAIL.n107 VTAIL.n106 0.155672
R249 VTAIL.n106 VTAIL.n94 0.155672
R250 VTAIL.n99 VTAIL.n94 0.155672
R251 VTAIL.n81 VTAIL.n43 0.155672
R252 VTAIL.n73 VTAIL.n43 0.155672
R253 VTAIL.n73 VTAIL.n72 0.155672
R254 VTAIL.n72 VTAIL.n48 0.155672
R255 VTAIL.n65 VTAIL.n48 0.155672
R256 VTAIL.n65 VTAIL.n64 0.155672
R257 VTAIL.n64 VTAIL.n52 0.155672
R258 VTAIL.n57 VTAIL.n52 0.155672
R259 VDD2.n77 VDD2.n41 289.615
R260 VDD2.n36 VDD2.n0 289.615
R261 VDD2.n78 VDD2.n77 185
R262 VDD2.n76 VDD2.n43 185
R263 VDD2.n75 VDD2.n74 185
R264 VDD2.n46 VDD2.n44 185
R265 VDD2.n69 VDD2.n68 185
R266 VDD2.n67 VDD2.n66 185
R267 VDD2.n50 VDD2.n49 185
R268 VDD2.n61 VDD2.n60 185
R269 VDD2.n59 VDD2.n58 185
R270 VDD2.n54 VDD2.n53 185
R271 VDD2.n12 VDD2.n11 185
R272 VDD2.n17 VDD2.n16 185
R273 VDD2.n19 VDD2.n18 185
R274 VDD2.n8 VDD2.n7 185
R275 VDD2.n25 VDD2.n24 185
R276 VDD2.n27 VDD2.n26 185
R277 VDD2.n4 VDD2.n3 185
R278 VDD2.n34 VDD2.n33 185
R279 VDD2.n35 VDD2.n2 185
R280 VDD2.n37 VDD2.n36 185
R281 VDD2.n55 VDD2.t0 149.524
R282 VDD2.n13 VDD2.t1 149.524
R283 VDD2.n77 VDD2.n76 104.615
R284 VDD2.n76 VDD2.n75 104.615
R285 VDD2.n75 VDD2.n44 104.615
R286 VDD2.n68 VDD2.n44 104.615
R287 VDD2.n68 VDD2.n67 104.615
R288 VDD2.n67 VDD2.n49 104.615
R289 VDD2.n60 VDD2.n49 104.615
R290 VDD2.n60 VDD2.n59 104.615
R291 VDD2.n59 VDD2.n53 104.615
R292 VDD2.n17 VDD2.n11 104.615
R293 VDD2.n18 VDD2.n17 104.615
R294 VDD2.n18 VDD2.n7 104.615
R295 VDD2.n25 VDD2.n7 104.615
R296 VDD2.n26 VDD2.n25 104.615
R297 VDD2.n26 VDD2.n3 104.615
R298 VDD2.n34 VDD2.n3 104.615
R299 VDD2.n35 VDD2.n34 104.615
R300 VDD2.n36 VDD2.n35 104.615
R301 VDD2.n82 VDD2.n40 86.1915
R302 VDD2.t0 VDD2.n53 52.3082
R303 VDD2.t1 VDD2.n11 52.3082
R304 VDD2.n82 VDD2.n81 50.6096
R305 VDD2.n78 VDD2.n43 13.1884
R306 VDD2.n37 VDD2.n2 13.1884
R307 VDD2.n79 VDD2.n41 12.8005
R308 VDD2.n74 VDD2.n45 12.8005
R309 VDD2.n33 VDD2.n32 12.8005
R310 VDD2.n38 VDD2.n0 12.8005
R311 VDD2.n73 VDD2.n46 12.0247
R312 VDD2.n31 VDD2.n4 12.0247
R313 VDD2.n70 VDD2.n69 11.249
R314 VDD2.n28 VDD2.n27 11.249
R315 VDD2.n66 VDD2.n48 10.4732
R316 VDD2.n24 VDD2.n6 10.4732
R317 VDD2.n55 VDD2.n54 10.2747
R318 VDD2.n13 VDD2.n12 10.2747
R319 VDD2.n65 VDD2.n50 9.69747
R320 VDD2.n23 VDD2.n8 9.69747
R321 VDD2.n81 VDD2.n80 9.45567
R322 VDD2.n40 VDD2.n39 9.45567
R323 VDD2.n57 VDD2.n56 9.3005
R324 VDD2.n52 VDD2.n51 9.3005
R325 VDD2.n63 VDD2.n62 9.3005
R326 VDD2.n65 VDD2.n64 9.3005
R327 VDD2.n48 VDD2.n47 9.3005
R328 VDD2.n71 VDD2.n70 9.3005
R329 VDD2.n73 VDD2.n72 9.3005
R330 VDD2.n45 VDD2.n42 9.3005
R331 VDD2.n80 VDD2.n79 9.3005
R332 VDD2.n39 VDD2.n38 9.3005
R333 VDD2.n15 VDD2.n14 9.3005
R334 VDD2.n10 VDD2.n9 9.3005
R335 VDD2.n21 VDD2.n20 9.3005
R336 VDD2.n23 VDD2.n22 9.3005
R337 VDD2.n6 VDD2.n5 9.3005
R338 VDD2.n29 VDD2.n28 9.3005
R339 VDD2.n31 VDD2.n30 9.3005
R340 VDD2.n32 VDD2.n1 9.3005
R341 VDD2.n62 VDD2.n61 8.92171
R342 VDD2.n20 VDD2.n19 8.92171
R343 VDD2.n58 VDD2.n52 8.14595
R344 VDD2.n16 VDD2.n10 8.14595
R345 VDD2.n57 VDD2.n54 7.3702
R346 VDD2.n15 VDD2.n12 7.3702
R347 VDD2.n58 VDD2.n57 5.81868
R348 VDD2.n16 VDD2.n15 5.81868
R349 VDD2.n61 VDD2.n52 5.04292
R350 VDD2.n19 VDD2.n10 5.04292
R351 VDD2.n62 VDD2.n50 4.26717
R352 VDD2.n20 VDD2.n8 4.26717
R353 VDD2.n66 VDD2.n65 3.49141
R354 VDD2.n24 VDD2.n23 3.49141
R355 VDD2.n56 VDD2.n55 2.84304
R356 VDD2.n14 VDD2.n13 2.84304
R357 VDD2.n69 VDD2.n48 2.71565
R358 VDD2.n27 VDD2.n6 2.71565
R359 VDD2.n70 VDD2.n46 1.93989
R360 VDD2.n28 VDD2.n4 1.93989
R361 VDD2.n81 VDD2.n41 1.16414
R362 VDD2.n74 VDD2.n73 1.16414
R363 VDD2.n33 VDD2.n31 1.16414
R364 VDD2.n40 VDD2.n0 1.16414
R365 VDD2 VDD2.n82 0.698776
R366 VDD2.n79 VDD2.n78 0.388379
R367 VDD2.n45 VDD2.n43 0.388379
R368 VDD2.n32 VDD2.n2 0.388379
R369 VDD2.n38 VDD2.n37 0.388379
R370 VDD2.n80 VDD2.n42 0.155672
R371 VDD2.n72 VDD2.n42 0.155672
R372 VDD2.n72 VDD2.n71 0.155672
R373 VDD2.n71 VDD2.n47 0.155672
R374 VDD2.n64 VDD2.n47 0.155672
R375 VDD2.n64 VDD2.n63 0.155672
R376 VDD2.n63 VDD2.n51 0.155672
R377 VDD2.n56 VDD2.n51 0.155672
R378 VDD2.n14 VDD2.n9 0.155672
R379 VDD2.n21 VDD2.n9 0.155672
R380 VDD2.n22 VDD2.n21 0.155672
R381 VDD2.n22 VDD2.n5 0.155672
R382 VDD2.n29 VDD2.n5 0.155672
R383 VDD2.n30 VDD2.n29 0.155672
R384 VDD2.n30 VDD2.n1 0.155672
R385 VDD2.n39 VDD2.n1 0.155672
R386 B.n562 B.n561 585
R387 B.n563 B.n562 585
R388 B.n225 B.n84 585
R389 B.n224 B.n223 585
R390 B.n222 B.n221 585
R391 B.n220 B.n219 585
R392 B.n218 B.n217 585
R393 B.n216 B.n215 585
R394 B.n214 B.n213 585
R395 B.n212 B.n211 585
R396 B.n210 B.n209 585
R397 B.n208 B.n207 585
R398 B.n206 B.n205 585
R399 B.n204 B.n203 585
R400 B.n202 B.n201 585
R401 B.n200 B.n199 585
R402 B.n198 B.n197 585
R403 B.n196 B.n195 585
R404 B.n194 B.n193 585
R405 B.n192 B.n191 585
R406 B.n190 B.n189 585
R407 B.n188 B.n187 585
R408 B.n186 B.n185 585
R409 B.n184 B.n183 585
R410 B.n182 B.n181 585
R411 B.n180 B.n179 585
R412 B.n178 B.n177 585
R413 B.n176 B.n175 585
R414 B.n174 B.n173 585
R415 B.n172 B.n171 585
R416 B.n170 B.n169 585
R417 B.n167 B.n166 585
R418 B.n165 B.n164 585
R419 B.n163 B.n162 585
R420 B.n161 B.n160 585
R421 B.n159 B.n158 585
R422 B.n157 B.n156 585
R423 B.n155 B.n154 585
R424 B.n153 B.n152 585
R425 B.n151 B.n150 585
R426 B.n149 B.n148 585
R427 B.n147 B.n146 585
R428 B.n145 B.n144 585
R429 B.n143 B.n142 585
R430 B.n141 B.n140 585
R431 B.n139 B.n138 585
R432 B.n137 B.n136 585
R433 B.n135 B.n134 585
R434 B.n133 B.n132 585
R435 B.n131 B.n130 585
R436 B.n129 B.n128 585
R437 B.n127 B.n126 585
R438 B.n125 B.n124 585
R439 B.n123 B.n122 585
R440 B.n121 B.n120 585
R441 B.n119 B.n118 585
R442 B.n117 B.n116 585
R443 B.n115 B.n114 585
R444 B.n113 B.n112 585
R445 B.n111 B.n110 585
R446 B.n109 B.n108 585
R447 B.n107 B.n106 585
R448 B.n105 B.n104 585
R449 B.n103 B.n102 585
R450 B.n101 B.n100 585
R451 B.n99 B.n98 585
R452 B.n97 B.n96 585
R453 B.n95 B.n94 585
R454 B.n93 B.n92 585
R455 B.n91 B.n90 585
R456 B.n560 B.n49 585
R457 B.n564 B.n49 585
R458 B.n559 B.n48 585
R459 B.n565 B.n48 585
R460 B.n558 B.n557 585
R461 B.n557 B.n44 585
R462 B.n556 B.n43 585
R463 B.n571 B.n43 585
R464 B.n555 B.n42 585
R465 B.n572 B.n42 585
R466 B.n554 B.n41 585
R467 B.n573 B.n41 585
R468 B.n553 B.n552 585
R469 B.n552 B.n37 585
R470 B.n551 B.n36 585
R471 B.n579 B.n36 585
R472 B.n550 B.n35 585
R473 B.n580 B.n35 585
R474 B.n549 B.n34 585
R475 B.n581 B.n34 585
R476 B.n548 B.n547 585
R477 B.n547 B.n30 585
R478 B.n546 B.n29 585
R479 B.n587 B.n29 585
R480 B.n545 B.n28 585
R481 B.n588 B.n28 585
R482 B.n544 B.n27 585
R483 B.n589 B.n27 585
R484 B.n543 B.n542 585
R485 B.n542 B.n23 585
R486 B.n541 B.n22 585
R487 B.n595 B.n22 585
R488 B.n540 B.n21 585
R489 B.n596 B.n21 585
R490 B.n539 B.n20 585
R491 B.n597 B.n20 585
R492 B.n538 B.n537 585
R493 B.n537 B.n16 585
R494 B.n536 B.n15 585
R495 B.n603 B.n15 585
R496 B.n535 B.n14 585
R497 B.n604 B.n14 585
R498 B.n534 B.n13 585
R499 B.n605 B.n13 585
R500 B.n533 B.n532 585
R501 B.n532 B.n12 585
R502 B.n531 B.n530 585
R503 B.n531 B.n8 585
R504 B.n529 B.n7 585
R505 B.n612 B.n7 585
R506 B.n528 B.n6 585
R507 B.n613 B.n6 585
R508 B.n527 B.n5 585
R509 B.n614 B.n5 585
R510 B.n526 B.n525 585
R511 B.n525 B.n4 585
R512 B.n524 B.n226 585
R513 B.n524 B.n523 585
R514 B.n514 B.n227 585
R515 B.n228 B.n227 585
R516 B.n516 B.n515 585
R517 B.n517 B.n516 585
R518 B.n513 B.n233 585
R519 B.n233 B.n232 585
R520 B.n512 B.n511 585
R521 B.n511 B.n510 585
R522 B.n235 B.n234 585
R523 B.n236 B.n235 585
R524 B.n503 B.n502 585
R525 B.n504 B.n503 585
R526 B.n501 B.n241 585
R527 B.n241 B.n240 585
R528 B.n500 B.n499 585
R529 B.n499 B.n498 585
R530 B.n243 B.n242 585
R531 B.n244 B.n243 585
R532 B.n491 B.n490 585
R533 B.n492 B.n491 585
R534 B.n489 B.n249 585
R535 B.n249 B.n248 585
R536 B.n488 B.n487 585
R537 B.n487 B.n486 585
R538 B.n251 B.n250 585
R539 B.n252 B.n251 585
R540 B.n479 B.n478 585
R541 B.n480 B.n479 585
R542 B.n477 B.n257 585
R543 B.n257 B.n256 585
R544 B.n476 B.n475 585
R545 B.n475 B.n474 585
R546 B.n259 B.n258 585
R547 B.n260 B.n259 585
R548 B.n467 B.n466 585
R549 B.n468 B.n467 585
R550 B.n465 B.n265 585
R551 B.n265 B.n264 585
R552 B.n464 B.n463 585
R553 B.n463 B.n462 585
R554 B.n267 B.n266 585
R555 B.n268 B.n267 585
R556 B.n455 B.n454 585
R557 B.n456 B.n455 585
R558 B.n453 B.n273 585
R559 B.n273 B.n272 585
R560 B.n447 B.n446 585
R561 B.n445 B.n309 585
R562 B.n444 B.n308 585
R563 B.n449 B.n308 585
R564 B.n443 B.n442 585
R565 B.n441 B.n440 585
R566 B.n439 B.n438 585
R567 B.n437 B.n436 585
R568 B.n435 B.n434 585
R569 B.n433 B.n432 585
R570 B.n431 B.n430 585
R571 B.n429 B.n428 585
R572 B.n427 B.n426 585
R573 B.n425 B.n424 585
R574 B.n423 B.n422 585
R575 B.n421 B.n420 585
R576 B.n419 B.n418 585
R577 B.n417 B.n416 585
R578 B.n415 B.n414 585
R579 B.n413 B.n412 585
R580 B.n411 B.n410 585
R581 B.n409 B.n408 585
R582 B.n407 B.n406 585
R583 B.n405 B.n404 585
R584 B.n403 B.n402 585
R585 B.n401 B.n400 585
R586 B.n399 B.n398 585
R587 B.n397 B.n396 585
R588 B.n395 B.n394 585
R589 B.n393 B.n392 585
R590 B.n391 B.n390 585
R591 B.n388 B.n387 585
R592 B.n386 B.n385 585
R593 B.n384 B.n383 585
R594 B.n382 B.n381 585
R595 B.n380 B.n379 585
R596 B.n378 B.n377 585
R597 B.n376 B.n375 585
R598 B.n374 B.n373 585
R599 B.n372 B.n371 585
R600 B.n370 B.n369 585
R601 B.n368 B.n367 585
R602 B.n366 B.n365 585
R603 B.n364 B.n363 585
R604 B.n362 B.n361 585
R605 B.n360 B.n359 585
R606 B.n358 B.n357 585
R607 B.n356 B.n355 585
R608 B.n354 B.n353 585
R609 B.n352 B.n351 585
R610 B.n350 B.n349 585
R611 B.n348 B.n347 585
R612 B.n346 B.n345 585
R613 B.n344 B.n343 585
R614 B.n342 B.n341 585
R615 B.n340 B.n339 585
R616 B.n338 B.n337 585
R617 B.n336 B.n335 585
R618 B.n334 B.n333 585
R619 B.n332 B.n331 585
R620 B.n330 B.n329 585
R621 B.n328 B.n327 585
R622 B.n326 B.n325 585
R623 B.n324 B.n323 585
R624 B.n322 B.n321 585
R625 B.n320 B.n319 585
R626 B.n318 B.n317 585
R627 B.n316 B.n315 585
R628 B.n275 B.n274 585
R629 B.n452 B.n451 585
R630 B.n271 B.n270 585
R631 B.n272 B.n271 585
R632 B.n458 B.n457 585
R633 B.n457 B.n456 585
R634 B.n459 B.n269 585
R635 B.n269 B.n268 585
R636 B.n461 B.n460 585
R637 B.n462 B.n461 585
R638 B.n263 B.n262 585
R639 B.n264 B.n263 585
R640 B.n470 B.n469 585
R641 B.n469 B.n468 585
R642 B.n471 B.n261 585
R643 B.n261 B.n260 585
R644 B.n473 B.n472 585
R645 B.n474 B.n473 585
R646 B.n255 B.n254 585
R647 B.n256 B.n255 585
R648 B.n482 B.n481 585
R649 B.n481 B.n480 585
R650 B.n483 B.n253 585
R651 B.n253 B.n252 585
R652 B.n485 B.n484 585
R653 B.n486 B.n485 585
R654 B.n247 B.n246 585
R655 B.n248 B.n247 585
R656 B.n494 B.n493 585
R657 B.n493 B.n492 585
R658 B.n495 B.n245 585
R659 B.n245 B.n244 585
R660 B.n497 B.n496 585
R661 B.n498 B.n497 585
R662 B.n239 B.n238 585
R663 B.n240 B.n239 585
R664 B.n506 B.n505 585
R665 B.n505 B.n504 585
R666 B.n507 B.n237 585
R667 B.n237 B.n236 585
R668 B.n509 B.n508 585
R669 B.n510 B.n509 585
R670 B.n231 B.n230 585
R671 B.n232 B.n231 585
R672 B.n519 B.n518 585
R673 B.n518 B.n517 585
R674 B.n520 B.n229 585
R675 B.n229 B.n228 585
R676 B.n522 B.n521 585
R677 B.n523 B.n522 585
R678 B.n3 B.n0 585
R679 B.n4 B.n3 585
R680 B.n611 B.n1 585
R681 B.n612 B.n611 585
R682 B.n610 B.n609 585
R683 B.n610 B.n8 585
R684 B.n608 B.n9 585
R685 B.n12 B.n9 585
R686 B.n607 B.n606 585
R687 B.n606 B.n605 585
R688 B.n11 B.n10 585
R689 B.n604 B.n11 585
R690 B.n602 B.n601 585
R691 B.n603 B.n602 585
R692 B.n600 B.n17 585
R693 B.n17 B.n16 585
R694 B.n599 B.n598 585
R695 B.n598 B.n597 585
R696 B.n19 B.n18 585
R697 B.n596 B.n19 585
R698 B.n594 B.n593 585
R699 B.n595 B.n594 585
R700 B.n592 B.n24 585
R701 B.n24 B.n23 585
R702 B.n591 B.n590 585
R703 B.n590 B.n589 585
R704 B.n26 B.n25 585
R705 B.n588 B.n26 585
R706 B.n586 B.n585 585
R707 B.n587 B.n586 585
R708 B.n584 B.n31 585
R709 B.n31 B.n30 585
R710 B.n583 B.n582 585
R711 B.n582 B.n581 585
R712 B.n33 B.n32 585
R713 B.n580 B.n33 585
R714 B.n578 B.n577 585
R715 B.n579 B.n578 585
R716 B.n576 B.n38 585
R717 B.n38 B.n37 585
R718 B.n575 B.n574 585
R719 B.n574 B.n573 585
R720 B.n40 B.n39 585
R721 B.n572 B.n40 585
R722 B.n570 B.n569 585
R723 B.n571 B.n570 585
R724 B.n568 B.n45 585
R725 B.n45 B.n44 585
R726 B.n567 B.n566 585
R727 B.n566 B.n565 585
R728 B.n47 B.n46 585
R729 B.n564 B.n47 585
R730 B.n615 B.n614 585
R731 B.n613 B.n2 585
R732 B.n90 B.n47 482.89
R733 B.n562 B.n49 482.89
R734 B.n451 B.n273 482.89
R735 B.n447 B.n271 482.89
R736 B.n87 B.t6 280.132
R737 B.n85 B.t10 280.132
R738 B.n312 B.t2 280.132
R739 B.n310 B.t13 280.132
R740 B.n85 B.t11 268.757
R741 B.n312 B.t5 268.757
R742 B.n87 B.t8 268.757
R743 B.n310 B.t15 268.757
R744 B.n563 B.n83 256.663
R745 B.n563 B.n82 256.663
R746 B.n563 B.n81 256.663
R747 B.n563 B.n80 256.663
R748 B.n563 B.n79 256.663
R749 B.n563 B.n78 256.663
R750 B.n563 B.n77 256.663
R751 B.n563 B.n76 256.663
R752 B.n563 B.n75 256.663
R753 B.n563 B.n74 256.663
R754 B.n563 B.n73 256.663
R755 B.n563 B.n72 256.663
R756 B.n563 B.n71 256.663
R757 B.n563 B.n70 256.663
R758 B.n563 B.n69 256.663
R759 B.n563 B.n68 256.663
R760 B.n563 B.n67 256.663
R761 B.n563 B.n66 256.663
R762 B.n563 B.n65 256.663
R763 B.n563 B.n64 256.663
R764 B.n563 B.n63 256.663
R765 B.n563 B.n62 256.663
R766 B.n563 B.n61 256.663
R767 B.n563 B.n60 256.663
R768 B.n563 B.n59 256.663
R769 B.n563 B.n58 256.663
R770 B.n563 B.n57 256.663
R771 B.n563 B.n56 256.663
R772 B.n563 B.n55 256.663
R773 B.n563 B.n54 256.663
R774 B.n563 B.n53 256.663
R775 B.n563 B.n52 256.663
R776 B.n563 B.n51 256.663
R777 B.n563 B.n50 256.663
R778 B.n449 B.n448 256.663
R779 B.n449 B.n276 256.663
R780 B.n449 B.n277 256.663
R781 B.n449 B.n278 256.663
R782 B.n449 B.n279 256.663
R783 B.n449 B.n280 256.663
R784 B.n449 B.n281 256.663
R785 B.n449 B.n282 256.663
R786 B.n449 B.n283 256.663
R787 B.n449 B.n284 256.663
R788 B.n449 B.n285 256.663
R789 B.n449 B.n286 256.663
R790 B.n449 B.n287 256.663
R791 B.n449 B.n288 256.663
R792 B.n449 B.n289 256.663
R793 B.n449 B.n290 256.663
R794 B.n449 B.n291 256.663
R795 B.n449 B.n292 256.663
R796 B.n449 B.n293 256.663
R797 B.n449 B.n294 256.663
R798 B.n449 B.n295 256.663
R799 B.n449 B.n296 256.663
R800 B.n449 B.n297 256.663
R801 B.n449 B.n298 256.663
R802 B.n449 B.n299 256.663
R803 B.n449 B.n300 256.663
R804 B.n449 B.n301 256.663
R805 B.n449 B.n302 256.663
R806 B.n449 B.n303 256.663
R807 B.n449 B.n304 256.663
R808 B.n449 B.n305 256.663
R809 B.n449 B.n306 256.663
R810 B.n449 B.n307 256.663
R811 B.n450 B.n449 256.663
R812 B.n617 B.n616 256.663
R813 B.n86 B.t12 211.157
R814 B.n313 B.t4 211.157
R815 B.n88 B.t9 211.157
R816 B.n311 B.t14 211.157
R817 B.n94 B.n93 163.367
R818 B.n98 B.n97 163.367
R819 B.n102 B.n101 163.367
R820 B.n106 B.n105 163.367
R821 B.n110 B.n109 163.367
R822 B.n114 B.n113 163.367
R823 B.n118 B.n117 163.367
R824 B.n122 B.n121 163.367
R825 B.n126 B.n125 163.367
R826 B.n130 B.n129 163.367
R827 B.n134 B.n133 163.367
R828 B.n138 B.n137 163.367
R829 B.n142 B.n141 163.367
R830 B.n146 B.n145 163.367
R831 B.n150 B.n149 163.367
R832 B.n154 B.n153 163.367
R833 B.n158 B.n157 163.367
R834 B.n162 B.n161 163.367
R835 B.n166 B.n165 163.367
R836 B.n171 B.n170 163.367
R837 B.n175 B.n174 163.367
R838 B.n179 B.n178 163.367
R839 B.n183 B.n182 163.367
R840 B.n187 B.n186 163.367
R841 B.n191 B.n190 163.367
R842 B.n195 B.n194 163.367
R843 B.n199 B.n198 163.367
R844 B.n203 B.n202 163.367
R845 B.n207 B.n206 163.367
R846 B.n211 B.n210 163.367
R847 B.n215 B.n214 163.367
R848 B.n219 B.n218 163.367
R849 B.n223 B.n222 163.367
R850 B.n562 B.n84 163.367
R851 B.n455 B.n273 163.367
R852 B.n455 B.n267 163.367
R853 B.n463 B.n267 163.367
R854 B.n463 B.n265 163.367
R855 B.n467 B.n265 163.367
R856 B.n467 B.n259 163.367
R857 B.n475 B.n259 163.367
R858 B.n475 B.n257 163.367
R859 B.n479 B.n257 163.367
R860 B.n479 B.n251 163.367
R861 B.n487 B.n251 163.367
R862 B.n487 B.n249 163.367
R863 B.n491 B.n249 163.367
R864 B.n491 B.n243 163.367
R865 B.n499 B.n243 163.367
R866 B.n499 B.n241 163.367
R867 B.n503 B.n241 163.367
R868 B.n503 B.n235 163.367
R869 B.n511 B.n235 163.367
R870 B.n511 B.n233 163.367
R871 B.n516 B.n233 163.367
R872 B.n516 B.n227 163.367
R873 B.n524 B.n227 163.367
R874 B.n525 B.n524 163.367
R875 B.n525 B.n5 163.367
R876 B.n6 B.n5 163.367
R877 B.n7 B.n6 163.367
R878 B.n531 B.n7 163.367
R879 B.n532 B.n531 163.367
R880 B.n532 B.n13 163.367
R881 B.n14 B.n13 163.367
R882 B.n15 B.n14 163.367
R883 B.n537 B.n15 163.367
R884 B.n537 B.n20 163.367
R885 B.n21 B.n20 163.367
R886 B.n22 B.n21 163.367
R887 B.n542 B.n22 163.367
R888 B.n542 B.n27 163.367
R889 B.n28 B.n27 163.367
R890 B.n29 B.n28 163.367
R891 B.n547 B.n29 163.367
R892 B.n547 B.n34 163.367
R893 B.n35 B.n34 163.367
R894 B.n36 B.n35 163.367
R895 B.n552 B.n36 163.367
R896 B.n552 B.n41 163.367
R897 B.n42 B.n41 163.367
R898 B.n43 B.n42 163.367
R899 B.n557 B.n43 163.367
R900 B.n557 B.n48 163.367
R901 B.n49 B.n48 163.367
R902 B.n309 B.n308 163.367
R903 B.n442 B.n308 163.367
R904 B.n440 B.n439 163.367
R905 B.n436 B.n435 163.367
R906 B.n432 B.n431 163.367
R907 B.n428 B.n427 163.367
R908 B.n424 B.n423 163.367
R909 B.n420 B.n419 163.367
R910 B.n416 B.n415 163.367
R911 B.n412 B.n411 163.367
R912 B.n408 B.n407 163.367
R913 B.n404 B.n403 163.367
R914 B.n400 B.n399 163.367
R915 B.n396 B.n395 163.367
R916 B.n392 B.n391 163.367
R917 B.n387 B.n386 163.367
R918 B.n383 B.n382 163.367
R919 B.n379 B.n378 163.367
R920 B.n375 B.n374 163.367
R921 B.n371 B.n370 163.367
R922 B.n367 B.n366 163.367
R923 B.n363 B.n362 163.367
R924 B.n359 B.n358 163.367
R925 B.n355 B.n354 163.367
R926 B.n351 B.n350 163.367
R927 B.n347 B.n346 163.367
R928 B.n343 B.n342 163.367
R929 B.n339 B.n338 163.367
R930 B.n335 B.n334 163.367
R931 B.n331 B.n330 163.367
R932 B.n327 B.n326 163.367
R933 B.n323 B.n322 163.367
R934 B.n319 B.n318 163.367
R935 B.n315 B.n275 163.367
R936 B.n457 B.n271 163.367
R937 B.n457 B.n269 163.367
R938 B.n461 B.n269 163.367
R939 B.n461 B.n263 163.367
R940 B.n469 B.n263 163.367
R941 B.n469 B.n261 163.367
R942 B.n473 B.n261 163.367
R943 B.n473 B.n255 163.367
R944 B.n481 B.n255 163.367
R945 B.n481 B.n253 163.367
R946 B.n485 B.n253 163.367
R947 B.n485 B.n247 163.367
R948 B.n493 B.n247 163.367
R949 B.n493 B.n245 163.367
R950 B.n497 B.n245 163.367
R951 B.n497 B.n239 163.367
R952 B.n505 B.n239 163.367
R953 B.n505 B.n237 163.367
R954 B.n509 B.n237 163.367
R955 B.n509 B.n231 163.367
R956 B.n518 B.n231 163.367
R957 B.n518 B.n229 163.367
R958 B.n522 B.n229 163.367
R959 B.n522 B.n3 163.367
R960 B.n615 B.n3 163.367
R961 B.n611 B.n2 163.367
R962 B.n611 B.n610 163.367
R963 B.n610 B.n9 163.367
R964 B.n606 B.n9 163.367
R965 B.n606 B.n11 163.367
R966 B.n602 B.n11 163.367
R967 B.n602 B.n17 163.367
R968 B.n598 B.n17 163.367
R969 B.n598 B.n19 163.367
R970 B.n594 B.n19 163.367
R971 B.n594 B.n24 163.367
R972 B.n590 B.n24 163.367
R973 B.n590 B.n26 163.367
R974 B.n586 B.n26 163.367
R975 B.n586 B.n31 163.367
R976 B.n582 B.n31 163.367
R977 B.n582 B.n33 163.367
R978 B.n578 B.n33 163.367
R979 B.n578 B.n38 163.367
R980 B.n574 B.n38 163.367
R981 B.n574 B.n40 163.367
R982 B.n570 B.n40 163.367
R983 B.n570 B.n45 163.367
R984 B.n566 B.n45 163.367
R985 B.n566 B.n47 163.367
R986 B.n449 B.n272 107.787
R987 B.n564 B.n563 107.787
R988 B.n90 B.n50 71.676
R989 B.n94 B.n51 71.676
R990 B.n98 B.n52 71.676
R991 B.n102 B.n53 71.676
R992 B.n106 B.n54 71.676
R993 B.n110 B.n55 71.676
R994 B.n114 B.n56 71.676
R995 B.n118 B.n57 71.676
R996 B.n122 B.n58 71.676
R997 B.n126 B.n59 71.676
R998 B.n130 B.n60 71.676
R999 B.n134 B.n61 71.676
R1000 B.n138 B.n62 71.676
R1001 B.n142 B.n63 71.676
R1002 B.n146 B.n64 71.676
R1003 B.n150 B.n65 71.676
R1004 B.n154 B.n66 71.676
R1005 B.n158 B.n67 71.676
R1006 B.n162 B.n68 71.676
R1007 B.n166 B.n69 71.676
R1008 B.n171 B.n70 71.676
R1009 B.n175 B.n71 71.676
R1010 B.n179 B.n72 71.676
R1011 B.n183 B.n73 71.676
R1012 B.n187 B.n74 71.676
R1013 B.n191 B.n75 71.676
R1014 B.n195 B.n76 71.676
R1015 B.n199 B.n77 71.676
R1016 B.n203 B.n78 71.676
R1017 B.n207 B.n79 71.676
R1018 B.n211 B.n80 71.676
R1019 B.n215 B.n81 71.676
R1020 B.n219 B.n82 71.676
R1021 B.n223 B.n83 71.676
R1022 B.n84 B.n83 71.676
R1023 B.n222 B.n82 71.676
R1024 B.n218 B.n81 71.676
R1025 B.n214 B.n80 71.676
R1026 B.n210 B.n79 71.676
R1027 B.n206 B.n78 71.676
R1028 B.n202 B.n77 71.676
R1029 B.n198 B.n76 71.676
R1030 B.n194 B.n75 71.676
R1031 B.n190 B.n74 71.676
R1032 B.n186 B.n73 71.676
R1033 B.n182 B.n72 71.676
R1034 B.n178 B.n71 71.676
R1035 B.n174 B.n70 71.676
R1036 B.n170 B.n69 71.676
R1037 B.n165 B.n68 71.676
R1038 B.n161 B.n67 71.676
R1039 B.n157 B.n66 71.676
R1040 B.n153 B.n65 71.676
R1041 B.n149 B.n64 71.676
R1042 B.n145 B.n63 71.676
R1043 B.n141 B.n62 71.676
R1044 B.n137 B.n61 71.676
R1045 B.n133 B.n60 71.676
R1046 B.n129 B.n59 71.676
R1047 B.n125 B.n58 71.676
R1048 B.n121 B.n57 71.676
R1049 B.n117 B.n56 71.676
R1050 B.n113 B.n55 71.676
R1051 B.n109 B.n54 71.676
R1052 B.n105 B.n53 71.676
R1053 B.n101 B.n52 71.676
R1054 B.n97 B.n51 71.676
R1055 B.n93 B.n50 71.676
R1056 B.n448 B.n447 71.676
R1057 B.n442 B.n276 71.676
R1058 B.n439 B.n277 71.676
R1059 B.n435 B.n278 71.676
R1060 B.n431 B.n279 71.676
R1061 B.n427 B.n280 71.676
R1062 B.n423 B.n281 71.676
R1063 B.n419 B.n282 71.676
R1064 B.n415 B.n283 71.676
R1065 B.n411 B.n284 71.676
R1066 B.n407 B.n285 71.676
R1067 B.n403 B.n286 71.676
R1068 B.n399 B.n287 71.676
R1069 B.n395 B.n288 71.676
R1070 B.n391 B.n289 71.676
R1071 B.n386 B.n290 71.676
R1072 B.n382 B.n291 71.676
R1073 B.n378 B.n292 71.676
R1074 B.n374 B.n293 71.676
R1075 B.n370 B.n294 71.676
R1076 B.n366 B.n295 71.676
R1077 B.n362 B.n296 71.676
R1078 B.n358 B.n297 71.676
R1079 B.n354 B.n298 71.676
R1080 B.n350 B.n299 71.676
R1081 B.n346 B.n300 71.676
R1082 B.n342 B.n301 71.676
R1083 B.n338 B.n302 71.676
R1084 B.n334 B.n303 71.676
R1085 B.n330 B.n304 71.676
R1086 B.n326 B.n305 71.676
R1087 B.n322 B.n306 71.676
R1088 B.n318 B.n307 71.676
R1089 B.n450 B.n275 71.676
R1090 B.n448 B.n309 71.676
R1091 B.n440 B.n276 71.676
R1092 B.n436 B.n277 71.676
R1093 B.n432 B.n278 71.676
R1094 B.n428 B.n279 71.676
R1095 B.n424 B.n280 71.676
R1096 B.n420 B.n281 71.676
R1097 B.n416 B.n282 71.676
R1098 B.n412 B.n283 71.676
R1099 B.n408 B.n284 71.676
R1100 B.n404 B.n285 71.676
R1101 B.n400 B.n286 71.676
R1102 B.n396 B.n287 71.676
R1103 B.n392 B.n288 71.676
R1104 B.n387 B.n289 71.676
R1105 B.n383 B.n290 71.676
R1106 B.n379 B.n291 71.676
R1107 B.n375 B.n292 71.676
R1108 B.n371 B.n293 71.676
R1109 B.n367 B.n294 71.676
R1110 B.n363 B.n295 71.676
R1111 B.n359 B.n296 71.676
R1112 B.n355 B.n297 71.676
R1113 B.n351 B.n298 71.676
R1114 B.n347 B.n299 71.676
R1115 B.n343 B.n300 71.676
R1116 B.n339 B.n301 71.676
R1117 B.n335 B.n302 71.676
R1118 B.n331 B.n303 71.676
R1119 B.n327 B.n304 71.676
R1120 B.n323 B.n305 71.676
R1121 B.n319 B.n306 71.676
R1122 B.n315 B.n307 71.676
R1123 B.n451 B.n450 71.676
R1124 B.n616 B.n615 71.676
R1125 B.n616 B.n2 71.676
R1126 B.n89 B.n88 59.5399
R1127 B.n168 B.n86 59.5399
R1128 B.n314 B.n313 59.5399
R1129 B.n389 B.n311 59.5399
R1130 B.n88 B.n87 57.6005
R1131 B.n86 B.n85 57.6005
R1132 B.n313 B.n312 57.6005
R1133 B.n311 B.n310 57.6005
R1134 B.n456 B.n272 56.8178
R1135 B.n456 B.n268 56.8178
R1136 B.n462 B.n268 56.8178
R1137 B.n462 B.n264 56.8178
R1138 B.n468 B.n264 56.8178
R1139 B.n468 B.n260 56.8178
R1140 B.n474 B.n260 56.8178
R1141 B.n480 B.n256 56.8178
R1142 B.n480 B.n252 56.8178
R1143 B.n486 B.n252 56.8178
R1144 B.n486 B.n248 56.8178
R1145 B.n492 B.n248 56.8178
R1146 B.n492 B.n244 56.8178
R1147 B.n498 B.n244 56.8178
R1148 B.n498 B.n240 56.8178
R1149 B.n504 B.n240 56.8178
R1150 B.n504 B.n236 56.8178
R1151 B.n510 B.n236 56.8178
R1152 B.n517 B.n232 56.8178
R1153 B.n517 B.n228 56.8178
R1154 B.n523 B.n228 56.8178
R1155 B.n523 B.n4 56.8178
R1156 B.n614 B.n4 56.8178
R1157 B.n614 B.n613 56.8178
R1158 B.n613 B.n612 56.8178
R1159 B.n612 B.n8 56.8178
R1160 B.n12 B.n8 56.8178
R1161 B.n605 B.n12 56.8178
R1162 B.n605 B.n604 56.8178
R1163 B.n603 B.n16 56.8178
R1164 B.n597 B.n16 56.8178
R1165 B.n597 B.n596 56.8178
R1166 B.n596 B.n595 56.8178
R1167 B.n595 B.n23 56.8178
R1168 B.n589 B.n23 56.8178
R1169 B.n589 B.n588 56.8178
R1170 B.n588 B.n587 56.8178
R1171 B.n587 B.n30 56.8178
R1172 B.n581 B.n30 56.8178
R1173 B.n581 B.n580 56.8178
R1174 B.n579 B.n37 56.8178
R1175 B.n573 B.n37 56.8178
R1176 B.n573 B.n572 56.8178
R1177 B.n572 B.n571 56.8178
R1178 B.n571 B.n44 56.8178
R1179 B.n565 B.n44 56.8178
R1180 B.n565 B.n564 56.8178
R1181 B.n474 B.t3 33.4225
R1182 B.t7 B.n579 33.4225
R1183 B.n446 B.n270 31.3761
R1184 B.n453 B.n452 31.3761
R1185 B.n561 B.n560 31.3761
R1186 B.n91 B.n46 31.3761
R1187 B.n510 B.t0 30.0803
R1188 B.t1 B.n603 30.0803
R1189 B.t0 B.n232 26.7381
R1190 B.n604 B.t1 26.7381
R1191 B.t3 B.n256 23.3959
R1192 B.n580 B.t7 23.3959
R1193 B B.n617 18.0485
R1194 B.n458 B.n270 10.6151
R1195 B.n459 B.n458 10.6151
R1196 B.n460 B.n459 10.6151
R1197 B.n460 B.n262 10.6151
R1198 B.n470 B.n262 10.6151
R1199 B.n471 B.n470 10.6151
R1200 B.n472 B.n471 10.6151
R1201 B.n472 B.n254 10.6151
R1202 B.n482 B.n254 10.6151
R1203 B.n483 B.n482 10.6151
R1204 B.n484 B.n483 10.6151
R1205 B.n484 B.n246 10.6151
R1206 B.n494 B.n246 10.6151
R1207 B.n495 B.n494 10.6151
R1208 B.n496 B.n495 10.6151
R1209 B.n496 B.n238 10.6151
R1210 B.n506 B.n238 10.6151
R1211 B.n507 B.n506 10.6151
R1212 B.n508 B.n507 10.6151
R1213 B.n508 B.n230 10.6151
R1214 B.n519 B.n230 10.6151
R1215 B.n520 B.n519 10.6151
R1216 B.n521 B.n520 10.6151
R1217 B.n521 B.n0 10.6151
R1218 B.n446 B.n445 10.6151
R1219 B.n445 B.n444 10.6151
R1220 B.n444 B.n443 10.6151
R1221 B.n443 B.n441 10.6151
R1222 B.n441 B.n438 10.6151
R1223 B.n438 B.n437 10.6151
R1224 B.n437 B.n434 10.6151
R1225 B.n434 B.n433 10.6151
R1226 B.n433 B.n430 10.6151
R1227 B.n430 B.n429 10.6151
R1228 B.n429 B.n426 10.6151
R1229 B.n426 B.n425 10.6151
R1230 B.n425 B.n422 10.6151
R1231 B.n422 B.n421 10.6151
R1232 B.n421 B.n418 10.6151
R1233 B.n418 B.n417 10.6151
R1234 B.n417 B.n414 10.6151
R1235 B.n414 B.n413 10.6151
R1236 B.n413 B.n410 10.6151
R1237 B.n410 B.n409 10.6151
R1238 B.n409 B.n406 10.6151
R1239 B.n406 B.n405 10.6151
R1240 B.n405 B.n402 10.6151
R1241 B.n402 B.n401 10.6151
R1242 B.n401 B.n398 10.6151
R1243 B.n398 B.n397 10.6151
R1244 B.n397 B.n394 10.6151
R1245 B.n394 B.n393 10.6151
R1246 B.n393 B.n390 10.6151
R1247 B.n388 B.n385 10.6151
R1248 B.n385 B.n384 10.6151
R1249 B.n384 B.n381 10.6151
R1250 B.n381 B.n380 10.6151
R1251 B.n380 B.n377 10.6151
R1252 B.n377 B.n376 10.6151
R1253 B.n376 B.n373 10.6151
R1254 B.n373 B.n372 10.6151
R1255 B.n369 B.n368 10.6151
R1256 B.n368 B.n365 10.6151
R1257 B.n365 B.n364 10.6151
R1258 B.n364 B.n361 10.6151
R1259 B.n361 B.n360 10.6151
R1260 B.n360 B.n357 10.6151
R1261 B.n357 B.n356 10.6151
R1262 B.n356 B.n353 10.6151
R1263 B.n353 B.n352 10.6151
R1264 B.n352 B.n349 10.6151
R1265 B.n349 B.n348 10.6151
R1266 B.n348 B.n345 10.6151
R1267 B.n345 B.n344 10.6151
R1268 B.n344 B.n341 10.6151
R1269 B.n341 B.n340 10.6151
R1270 B.n340 B.n337 10.6151
R1271 B.n337 B.n336 10.6151
R1272 B.n336 B.n333 10.6151
R1273 B.n333 B.n332 10.6151
R1274 B.n332 B.n329 10.6151
R1275 B.n329 B.n328 10.6151
R1276 B.n328 B.n325 10.6151
R1277 B.n325 B.n324 10.6151
R1278 B.n324 B.n321 10.6151
R1279 B.n321 B.n320 10.6151
R1280 B.n320 B.n317 10.6151
R1281 B.n317 B.n316 10.6151
R1282 B.n316 B.n274 10.6151
R1283 B.n452 B.n274 10.6151
R1284 B.n454 B.n453 10.6151
R1285 B.n454 B.n266 10.6151
R1286 B.n464 B.n266 10.6151
R1287 B.n465 B.n464 10.6151
R1288 B.n466 B.n465 10.6151
R1289 B.n466 B.n258 10.6151
R1290 B.n476 B.n258 10.6151
R1291 B.n477 B.n476 10.6151
R1292 B.n478 B.n477 10.6151
R1293 B.n478 B.n250 10.6151
R1294 B.n488 B.n250 10.6151
R1295 B.n489 B.n488 10.6151
R1296 B.n490 B.n489 10.6151
R1297 B.n490 B.n242 10.6151
R1298 B.n500 B.n242 10.6151
R1299 B.n501 B.n500 10.6151
R1300 B.n502 B.n501 10.6151
R1301 B.n502 B.n234 10.6151
R1302 B.n512 B.n234 10.6151
R1303 B.n513 B.n512 10.6151
R1304 B.n515 B.n513 10.6151
R1305 B.n515 B.n514 10.6151
R1306 B.n514 B.n226 10.6151
R1307 B.n526 B.n226 10.6151
R1308 B.n527 B.n526 10.6151
R1309 B.n528 B.n527 10.6151
R1310 B.n529 B.n528 10.6151
R1311 B.n530 B.n529 10.6151
R1312 B.n533 B.n530 10.6151
R1313 B.n534 B.n533 10.6151
R1314 B.n535 B.n534 10.6151
R1315 B.n536 B.n535 10.6151
R1316 B.n538 B.n536 10.6151
R1317 B.n539 B.n538 10.6151
R1318 B.n540 B.n539 10.6151
R1319 B.n541 B.n540 10.6151
R1320 B.n543 B.n541 10.6151
R1321 B.n544 B.n543 10.6151
R1322 B.n545 B.n544 10.6151
R1323 B.n546 B.n545 10.6151
R1324 B.n548 B.n546 10.6151
R1325 B.n549 B.n548 10.6151
R1326 B.n550 B.n549 10.6151
R1327 B.n551 B.n550 10.6151
R1328 B.n553 B.n551 10.6151
R1329 B.n554 B.n553 10.6151
R1330 B.n555 B.n554 10.6151
R1331 B.n556 B.n555 10.6151
R1332 B.n558 B.n556 10.6151
R1333 B.n559 B.n558 10.6151
R1334 B.n560 B.n559 10.6151
R1335 B.n609 B.n1 10.6151
R1336 B.n609 B.n608 10.6151
R1337 B.n608 B.n607 10.6151
R1338 B.n607 B.n10 10.6151
R1339 B.n601 B.n10 10.6151
R1340 B.n601 B.n600 10.6151
R1341 B.n600 B.n599 10.6151
R1342 B.n599 B.n18 10.6151
R1343 B.n593 B.n18 10.6151
R1344 B.n593 B.n592 10.6151
R1345 B.n592 B.n591 10.6151
R1346 B.n591 B.n25 10.6151
R1347 B.n585 B.n25 10.6151
R1348 B.n585 B.n584 10.6151
R1349 B.n584 B.n583 10.6151
R1350 B.n583 B.n32 10.6151
R1351 B.n577 B.n32 10.6151
R1352 B.n577 B.n576 10.6151
R1353 B.n576 B.n575 10.6151
R1354 B.n575 B.n39 10.6151
R1355 B.n569 B.n39 10.6151
R1356 B.n569 B.n568 10.6151
R1357 B.n568 B.n567 10.6151
R1358 B.n567 B.n46 10.6151
R1359 B.n92 B.n91 10.6151
R1360 B.n95 B.n92 10.6151
R1361 B.n96 B.n95 10.6151
R1362 B.n99 B.n96 10.6151
R1363 B.n100 B.n99 10.6151
R1364 B.n103 B.n100 10.6151
R1365 B.n104 B.n103 10.6151
R1366 B.n107 B.n104 10.6151
R1367 B.n108 B.n107 10.6151
R1368 B.n111 B.n108 10.6151
R1369 B.n112 B.n111 10.6151
R1370 B.n115 B.n112 10.6151
R1371 B.n116 B.n115 10.6151
R1372 B.n119 B.n116 10.6151
R1373 B.n120 B.n119 10.6151
R1374 B.n123 B.n120 10.6151
R1375 B.n124 B.n123 10.6151
R1376 B.n127 B.n124 10.6151
R1377 B.n128 B.n127 10.6151
R1378 B.n131 B.n128 10.6151
R1379 B.n132 B.n131 10.6151
R1380 B.n135 B.n132 10.6151
R1381 B.n136 B.n135 10.6151
R1382 B.n139 B.n136 10.6151
R1383 B.n140 B.n139 10.6151
R1384 B.n143 B.n140 10.6151
R1385 B.n144 B.n143 10.6151
R1386 B.n147 B.n144 10.6151
R1387 B.n148 B.n147 10.6151
R1388 B.n152 B.n151 10.6151
R1389 B.n155 B.n152 10.6151
R1390 B.n156 B.n155 10.6151
R1391 B.n159 B.n156 10.6151
R1392 B.n160 B.n159 10.6151
R1393 B.n163 B.n160 10.6151
R1394 B.n164 B.n163 10.6151
R1395 B.n167 B.n164 10.6151
R1396 B.n172 B.n169 10.6151
R1397 B.n173 B.n172 10.6151
R1398 B.n176 B.n173 10.6151
R1399 B.n177 B.n176 10.6151
R1400 B.n180 B.n177 10.6151
R1401 B.n181 B.n180 10.6151
R1402 B.n184 B.n181 10.6151
R1403 B.n185 B.n184 10.6151
R1404 B.n188 B.n185 10.6151
R1405 B.n189 B.n188 10.6151
R1406 B.n192 B.n189 10.6151
R1407 B.n193 B.n192 10.6151
R1408 B.n196 B.n193 10.6151
R1409 B.n197 B.n196 10.6151
R1410 B.n200 B.n197 10.6151
R1411 B.n201 B.n200 10.6151
R1412 B.n204 B.n201 10.6151
R1413 B.n205 B.n204 10.6151
R1414 B.n208 B.n205 10.6151
R1415 B.n209 B.n208 10.6151
R1416 B.n212 B.n209 10.6151
R1417 B.n213 B.n212 10.6151
R1418 B.n216 B.n213 10.6151
R1419 B.n217 B.n216 10.6151
R1420 B.n220 B.n217 10.6151
R1421 B.n221 B.n220 10.6151
R1422 B.n224 B.n221 10.6151
R1423 B.n225 B.n224 10.6151
R1424 B.n561 B.n225 10.6151
R1425 B.n617 B.n0 8.11757
R1426 B.n617 B.n1 8.11757
R1427 B.n389 B.n388 6.5566
R1428 B.n372 B.n314 6.5566
R1429 B.n151 B.n89 6.5566
R1430 B.n168 B.n167 6.5566
R1431 B.n390 B.n389 4.05904
R1432 B.n369 B.n314 4.05904
R1433 B.n148 B.n89 4.05904
R1434 B.n169 B.n168 4.05904
R1435 VP.n0 VP.t1 154.772
R1436 VP.n0 VP.t0 113.123
R1437 VP VP.n0 0.431811
R1438 VDD1.n36 VDD1.n0 289.615
R1439 VDD1.n77 VDD1.n41 289.615
R1440 VDD1.n37 VDD1.n36 185
R1441 VDD1.n35 VDD1.n2 185
R1442 VDD1.n34 VDD1.n33 185
R1443 VDD1.n5 VDD1.n3 185
R1444 VDD1.n28 VDD1.n27 185
R1445 VDD1.n26 VDD1.n25 185
R1446 VDD1.n9 VDD1.n8 185
R1447 VDD1.n20 VDD1.n19 185
R1448 VDD1.n18 VDD1.n17 185
R1449 VDD1.n13 VDD1.n12 185
R1450 VDD1.n53 VDD1.n52 185
R1451 VDD1.n58 VDD1.n57 185
R1452 VDD1.n60 VDD1.n59 185
R1453 VDD1.n49 VDD1.n48 185
R1454 VDD1.n66 VDD1.n65 185
R1455 VDD1.n68 VDD1.n67 185
R1456 VDD1.n45 VDD1.n44 185
R1457 VDD1.n75 VDD1.n74 185
R1458 VDD1.n76 VDD1.n43 185
R1459 VDD1.n78 VDD1.n77 185
R1460 VDD1.n14 VDD1.t0 149.524
R1461 VDD1.n54 VDD1.t1 149.524
R1462 VDD1.n36 VDD1.n35 104.615
R1463 VDD1.n35 VDD1.n34 104.615
R1464 VDD1.n34 VDD1.n3 104.615
R1465 VDD1.n27 VDD1.n3 104.615
R1466 VDD1.n27 VDD1.n26 104.615
R1467 VDD1.n26 VDD1.n8 104.615
R1468 VDD1.n19 VDD1.n8 104.615
R1469 VDD1.n19 VDD1.n18 104.615
R1470 VDD1.n18 VDD1.n12 104.615
R1471 VDD1.n58 VDD1.n52 104.615
R1472 VDD1.n59 VDD1.n58 104.615
R1473 VDD1.n59 VDD1.n48 104.615
R1474 VDD1.n66 VDD1.n48 104.615
R1475 VDD1.n67 VDD1.n66 104.615
R1476 VDD1.n67 VDD1.n44 104.615
R1477 VDD1.n75 VDD1.n44 104.615
R1478 VDD1.n76 VDD1.n75 104.615
R1479 VDD1.n77 VDD1.n76 104.615
R1480 VDD1 VDD1.n81 87.3564
R1481 VDD1.t0 VDD1.n12 52.3082
R1482 VDD1.t1 VDD1.n52 52.3082
R1483 VDD1 VDD1.n40 51.3079
R1484 VDD1.n37 VDD1.n2 13.1884
R1485 VDD1.n78 VDD1.n43 13.1884
R1486 VDD1.n38 VDD1.n0 12.8005
R1487 VDD1.n33 VDD1.n4 12.8005
R1488 VDD1.n74 VDD1.n73 12.8005
R1489 VDD1.n79 VDD1.n41 12.8005
R1490 VDD1.n32 VDD1.n5 12.0247
R1491 VDD1.n72 VDD1.n45 12.0247
R1492 VDD1.n29 VDD1.n28 11.249
R1493 VDD1.n69 VDD1.n68 11.249
R1494 VDD1.n25 VDD1.n7 10.4732
R1495 VDD1.n65 VDD1.n47 10.4732
R1496 VDD1.n14 VDD1.n13 10.2747
R1497 VDD1.n54 VDD1.n53 10.2747
R1498 VDD1.n24 VDD1.n9 9.69747
R1499 VDD1.n64 VDD1.n49 9.69747
R1500 VDD1.n40 VDD1.n39 9.45567
R1501 VDD1.n81 VDD1.n80 9.45567
R1502 VDD1.n16 VDD1.n15 9.3005
R1503 VDD1.n11 VDD1.n10 9.3005
R1504 VDD1.n22 VDD1.n21 9.3005
R1505 VDD1.n24 VDD1.n23 9.3005
R1506 VDD1.n7 VDD1.n6 9.3005
R1507 VDD1.n30 VDD1.n29 9.3005
R1508 VDD1.n32 VDD1.n31 9.3005
R1509 VDD1.n4 VDD1.n1 9.3005
R1510 VDD1.n39 VDD1.n38 9.3005
R1511 VDD1.n80 VDD1.n79 9.3005
R1512 VDD1.n56 VDD1.n55 9.3005
R1513 VDD1.n51 VDD1.n50 9.3005
R1514 VDD1.n62 VDD1.n61 9.3005
R1515 VDD1.n64 VDD1.n63 9.3005
R1516 VDD1.n47 VDD1.n46 9.3005
R1517 VDD1.n70 VDD1.n69 9.3005
R1518 VDD1.n72 VDD1.n71 9.3005
R1519 VDD1.n73 VDD1.n42 9.3005
R1520 VDD1.n21 VDD1.n20 8.92171
R1521 VDD1.n61 VDD1.n60 8.92171
R1522 VDD1.n17 VDD1.n11 8.14595
R1523 VDD1.n57 VDD1.n51 8.14595
R1524 VDD1.n16 VDD1.n13 7.3702
R1525 VDD1.n56 VDD1.n53 7.3702
R1526 VDD1.n17 VDD1.n16 5.81868
R1527 VDD1.n57 VDD1.n56 5.81868
R1528 VDD1.n20 VDD1.n11 5.04292
R1529 VDD1.n60 VDD1.n51 5.04292
R1530 VDD1.n21 VDD1.n9 4.26717
R1531 VDD1.n61 VDD1.n49 4.26717
R1532 VDD1.n25 VDD1.n24 3.49141
R1533 VDD1.n65 VDD1.n64 3.49141
R1534 VDD1.n15 VDD1.n14 2.84304
R1535 VDD1.n55 VDD1.n54 2.84304
R1536 VDD1.n28 VDD1.n7 2.71565
R1537 VDD1.n68 VDD1.n47 2.71565
R1538 VDD1.n29 VDD1.n5 1.93989
R1539 VDD1.n69 VDD1.n45 1.93989
R1540 VDD1.n40 VDD1.n0 1.16414
R1541 VDD1.n33 VDD1.n32 1.16414
R1542 VDD1.n74 VDD1.n72 1.16414
R1543 VDD1.n81 VDD1.n41 1.16414
R1544 VDD1.n38 VDD1.n37 0.388379
R1545 VDD1.n4 VDD1.n2 0.388379
R1546 VDD1.n73 VDD1.n43 0.388379
R1547 VDD1.n79 VDD1.n78 0.388379
R1548 VDD1.n39 VDD1.n1 0.155672
R1549 VDD1.n31 VDD1.n1 0.155672
R1550 VDD1.n31 VDD1.n30 0.155672
R1551 VDD1.n30 VDD1.n6 0.155672
R1552 VDD1.n23 VDD1.n6 0.155672
R1553 VDD1.n23 VDD1.n22 0.155672
R1554 VDD1.n22 VDD1.n10 0.155672
R1555 VDD1.n15 VDD1.n10 0.155672
R1556 VDD1.n55 VDD1.n50 0.155672
R1557 VDD1.n62 VDD1.n50 0.155672
R1558 VDD1.n63 VDD1.n62 0.155672
R1559 VDD1.n63 VDD1.n46 0.155672
R1560 VDD1.n70 VDD1.n46 0.155672
R1561 VDD1.n71 VDD1.n70 0.155672
R1562 VDD1.n71 VDD1.n42 0.155672
R1563 VDD1.n80 VDD1.n42 0.155672
C0 VP VN 4.71747f
C1 VTAIL VDD1 3.98979f
C2 VP VDD2 0.334421f
C3 VN VDD1 0.14814f
C4 VDD2 VDD1 0.678958f
C5 VN VTAIL 1.77182f
C6 VDD2 VTAIL 4.04165f
C7 VP VDD1 2.10153f
C8 VN VDD2 1.91705f
C9 VP VTAIL 1.78604f
C10 VDD2 B 3.665515f
C11 VDD1 B 6.16475f
C12 VTAIL B 5.68337f
C13 VN B 8.23652f
C14 VP B 6.172545f
C15 VDD1.n0 B 0.02728f
C16 VDD1.n1 B 0.020914f
C17 VDD1.n2 B 0.011569f
C18 VDD1.n3 B 0.026563f
C19 VDD1.n4 B 0.011238f
C20 VDD1.n5 B 0.011899f
C21 VDD1.n6 B 0.020914f
C22 VDD1.n7 B 0.011238f
C23 VDD1.n8 B 0.026563f
C24 VDD1.n9 B 0.011899f
C25 VDD1.n10 B 0.020914f
C26 VDD1.n11 B 0.011238f
C27 VDD1.n12 B 0.019922f
C28 VDD1.n13 B 0.018778f
C29 VDD1.t0 B 0.044414f
C30 VDD1.n14 B 0.11781f
C31 VDD1.n15 B 0.672718f
C32 VDD1.n16 B 0.011238f
C33 VDD1.n17 B 0.011899f
C34 VDD1.n18 B 0.026563f
C35 VDD1.n19 B 0.026563f
C36 VDD1.n20 B 0.011899f
C37 VDD1.n21 B 0.011238f
C38 VDD1.n22 B 0.020914f
C39 VDD1.n23 B 0.020914f
C40 VDD1.n24 B 0.011238f
C41 VDD1.n25 B 0.011899f
C42 VDD1.n26 B 0.026563f
C43 VDD1.n27 B 0.026563f
C44 VDD1.n28 B 0.011899f
C45 VDD1.n29 B 0.011238f
C46 VDD1.n30 B 0.020914f
C47 VDD1.n31 B 0.020914f
C48 VDD1.n32 B 0.011238f
C49 VDD1.n33 B 0.011899f
C50 VDD1.n34 B 0.026563f
C51 VDD1.n35 B 0.026563f
C52 VDD1.n36 B 0.053762f
C53 VDD1.n37 B 0.011569f
C54 VDD1.n38 B 0.011238f
C55 VDD1.n39 B 0.050913f
C56 VDD1.n40 B 0.045404f
C57 VDD1.n41 B 0.02728f
C58 VDD1.n42 B 0.020914f
C59 VDD1.n43 B 0.011569f
C60 VDD1.n44 B 0.026563f
C61 VDD1.n45 B 0.011899f
C62 VDD1.n46 B 0.020914f
C63 VDD1.n47 B 0.011238f
C64 VDD1.n48 B 0.026563f
C65 VDD1.n49 B 0.011899f
C66 VDD1.n50 B 0.020914f
C67 VDD1.n51 B 0.011238f
C68 VDD1.n52 B 0.019922f
C69 VDD1.n53 B 0.018778f
C70 VDD1.t1 B 0.044414f
C71 VDD1.n54 B 0.11781f
C72 VDD1.n55 B 0.672718f
C73 VDD1.n56 B 0.011238f
C74 VDD1.n57 B 0.011899f
C75 VDD1.n58 B 0.026563f
C76 VDD1.n59 B 0.026563f
C77 VDD1.n60 B 0.011899f
C78 VDD1.n61 B 0.011238f
C79 VDD1.n62 B 0.020914f
C80 VDD1.n63 B 0.020914f
C81 VDD1.n64 B 0.011238f
C82 VDD1.n65 B 0.011899f
C83 VDD1.n66 B 0.026563f
C84 VDD1.n67 B 0.026563f
C85 VDD1.n68 B 0.011899f
C86 VDD1.n69 B 0.011238f
C87 VDD1.n70 B 0.020914f
C88 VDD1.n71 B 0.020914f
C89 VDD1.n72 B 0.011238f
C90 VDD1.n73 B 0.011238f
C91 VDD1.n74 B 0.011899f
C92 VDD1.n75 B 0.026563f
C93 VDD1.n76 B 0.026563f
C94 VDD1.n77 B 0.053762f
C95 VDD1.n78 B 0.011569f
C96 VDD1.n79 B 0.011238f
C97 VDD1.n80 B 0.050913f
C98 VDD1.n81 B 0.526537f
C99 VP.t0 B 1.7305f
C100 VP.t1 B 2.17671f
C101 VP.n0 B 2.82432f
C102 VDD2.n0 B 0.018118f
C103 VDD2.n1 B 0.01389f
C104 VDD2.n2 B 0.007683f
C105 VDD2.n3 B 0.017642f
C106 VDD2.n4 B 0.007903f
C107 VDD2.n5 B 0.01389f
C108 VDD2.n6 B 0.007464f
C109 VDD2.n7 B 0.017642f
C110 VDD2.n8 B 0.007903f
C111 VDD2.n9 B 0.01389f
C112 VDD2.n10 B 0.007464f
C113 VDD2.n11 B 0.013231f
C114 VDD2.n12 B 0.012472f
C115 VDD2.t1 B 0.029497f
C116 VDD2.n13 B 0.078243f
C117 VDD2.n14 B 0.446784f
C118 VDD2.n15 B 0.007464f
C119 VDD2.n16 B 0.007903f
C120 VDD2.n17 B 0.017642f
C121 VDD2.n18 B 0.017642f
C122 VDD2.n19 B 0.007903f
C123 VDD2.n20 B 0.007464f
C124 VDD2.n21 B 0.01389f
C125 VDD2.n22 B 0.01389f
C126 VDD2.n23 B 0.007464f
C127 VDD2.n24 B 0.007903f
C128 VDD2.n25 B 0.017642f
C129 VDD2.n26 B 0.017642f
C130 VDD2.n27 B 0.007903f
C131 VDD2.n28 B 0.007464f
C132 VDD2.n29 B 0.01389f
C133 VDD2.n30 B 0.01389f
C134 VDD2.n31 B 0.007464f
C135 VDD2.n32 B 0.007464f
C136 VDD2.n33 B 0.007903f
C137 VDD2.n34 B 0.017642f
C138 VDD2.n35 B 0.017642f
C139 VDD2.n36 B 0.035706f
C140 VDD2.n37 B 0.007683f
C141 VDD2.n38 B 0.007464f
C142 VDD2.n39 B 0.033814f
C143 VDD2.n40 B 0.324747f
C144 VDD2.n41 B 0.018118f
C145 VDD2.n42 B 0.01389f
C146 VDD2.n43 B 0.007683f
C147 VDD2.n44 B 0.017642f
C148 VDD2.n45 B 0.007464f
C149 VDD2.n46 B 0.007903f
C150 VDD2.n47 B 0.01389f
C151 VDD2.n48 B 0.007464f
C152 VDD2.n49 B 0.017642f
C153 VDD2.n50 B 0.007903f
C154 VDD2.n51 B 0.01389f
C155 VDD2.n52 B 0.007464f
C156 VDD2.n53 B 0.013231f
C157 VDD2.n54 B 0.012472f
C158 VDD2.t0 B 0.029497f
C159 VDD2.n55 B 0.078243f
C160 VDD2.n56 B 0.446784f
C161 VDD2.n57 B 0.007464f
C162 VDD2.n58 B 0.007903f
C163 VDD2.n59 B 0.017642f
C164 VDD2.n60 B 0.017642f
C165 VDD2.n61 B 0.007903f
C166 VDD2.n62 B 0.007464f
C167 VDD2.n63 B 0.01389f
C168 VDD2.n64 B 0.01389f
C169 VDD2.n65 B 0.007464f
C170 VDD2.n66 B 0.007903f
C171 VDD2.n67 B 0.017642f
C172 VDD2.n68 B 0.017642f
C173 VDD2.n69 B 0.007903f
C174 VDD2.n70 B 0.007464f
C175 VDD2.n71 B 0.01389f
C176 VDD2.n72 B 0.01389f
C177 VDD2.n73 B 0.007464f
C178 VDD2.n74 B 0.007903f
C179 VDD2.n75 B 0.017642f
C180 VDD2.n76 B 0.017642f
C181 VDD2.n77 B 0.035706f
C182 VDD2.n78 B 0.007683f
C183 VDD2.n79 B 0.007464f
C184 VDD2.n80 B 0.033814f
C185 VDD2.n81 B 0.029353f
C186 VDD2.n82 B 1.46878f
C187 VTAIL.n0 B 0.01991f
C188 VTAIL.n1 B 0.015264f
C189 VTAIL.n2 B 0.008443f
C190 VTAIL.n3 B 0.019387f
C191 VTAIL.n4 B 0.008685f
C192 VTAIL.n5 B 0.015264f
C193 VTAIL.n6 B 0.008202f
C194 VTAIL.n7 B 0.019387f
C195 VTAIL.n8 B 0.008685f
C196 VTAIL.n9 B 0.015264f
C197 VTAIL.n10 B 0.008202f
C198 VTAIL.n11 B 0.01454f
C199 VTAIL.n12 B 0.013705f
C200 VTAIL.t0 B 0.032414f
C201 VTAIL.n13 B 0.085981f
C202 VTAIL.n14 B 0.490969f
C203 VTAIL.n15 B 0.008202f
C204 VTAIL.n16 B 0.008685f
C205 VTAIL.n17 B 0.019387f
C206 VTAIL.n18 B 0.019387f
C207 VTAIL.n19 B 0.008685f
C208 VTAIL.n20 B 0.008202f
C209 VTAIL.n21 B 0.015264f
C210 VTAIL.n22 B 0.015264f
C211 VTAIL.n23 B 0.008202f
C212 VTAIL.n24 B 0.008685f
C213 VTAIL.n25 B 0.019387f
C214 VTAIL.n26 B 0.019387f
C215 VTAIL.n27 B 0.008685f
C216 VTAIL.n28 B 0.008202f
C217 VTAIL.n29 B 0.015264f
C218 VTAIL.n30 B 0.015264f
C219 VTAIL.n31 B 0.008202f
C220 VTAIL.n32 B 0.008202f
C221 VTAIL.n33 B 0.008685f
C222 VTAIL.n34 B 0.019387f
C223 VTAIL.n35 B 0.019387f
C224 VTAIL.n36 B 0.039237f
C225 VTAIL.n37 B 0.008443f
C226 VTAIL.n38 B 0.008202f
C227 VTAIL.n39 B 0.037158f
C228 VTAIL.n40 B 0.02173f
C229 VTAIL.n41 B 0.865265f
C230 VTAIL.n42 B 0.01991f
C231 VTAIL.n43 B 0.015264f
C232 VTAIL.n44 B 0.008443f
C233 VTAIL.n45 B 0.019387f
C234 VTAIL.n46 B 0.008202f
C235 VTAIL.n47 B 0.008685f
C236 VTAIL.n48 B 0.015264f
C237 VTAIL.n49 B 0.008202f
C238 VTAIL.n50 B 0.019387f
C239 VTAIL.n51 B 0.008685f
C240 VTAIL.n52 B 0.015264f
C241 VTAIL.n53 B 0.008202f
C242 VTAIL.n54 B 0.01454f
C243 VTAIL.n55 B 0.013705f
C244 VTAIL.t2 B 0.032414f
C245 VTAIL.n56 B 0.085981f
C246 VTAIL.n57 B 0.490969f
C247 VTAIL.n58 B 0.008202f
C248 VTAIL.n59 B 0.008685f
C249 VTAIL.n60 B 0.019387f
C250 VTAIL.n61 B 0.019387f
C251 VTAIL.n62 B 0.008685f
C252 VTAIL.n63 B 0.008202f
C253 VTAIL.n64 B 0.015264f
C254 VTAIL.n65 B 0.015264f
C255 VTAIL.n66 B 0.008202f
C256 VTAIL.n67 B 0.008685f
C257 VTAIL.n68 B 0.019387f
C258 VTAIL.n69 B 0.019387f
C259 VTAIL.n70 B 0.008685f
C260 VTAIL.n71 B 0.008202f
C261 VTAIL.n72 B 0.015264f
C262 VTAIL.n73 B 0.015264f
C263 VTAIL.n74 B 0.008202f
C264 VTAIL.n75 B 0.008685f
C265 VTAIL.n76 B 0.019387f
C266 VTAIL.n77 B 0.019387f
C267 VTAIL.n78 B 0.039237f
C268 VTAIL.n79 B 0.008443f
C269 VTAIL.n80 B 0.008202f
C270 VTAIL.n81 B 0.037158f
C271 VTAIL.n82 B 0.02173f
C272 VTAIL.n83 B 0.893885f
C273 VTAIL.n84 B 0.01991f
C274 VTAIL.n85 B 0.015264f
C275 VTAIL.n86 B 0.008443f
C276 VTAIL.n87 B 0.019387f
C277 VTAIL.n88 B 0.008202f
C278 VTAIL.n89 B 0.008685f
C279 VTAIL.n90 B 0.015264f
C280 VTAIL.n91 B 0.008202f
C281 VTAIL.n92 B 0.019387f
C282 VTAIL.n93 B 0.008685f
C283 VTAIL.n94 B 0.015264f
C284 VTAIL.n95 B 0.008202f
C285 VTAIL.n96 B 0.01454f
C286 VTAIL.n97 B 0.013705f
C287 VTAIL.t1 B 0.032414f
C288 VTAIL.n98 B 0.085981f
C289 VTAIL.n99 B 0.490969f
C290 VTAIL.n100 B 0.008202f
C291 VTAIL.n101 B 0.008685f
C292 VTAIL.n102 B 0.019387f
C293 VTAIL.n103 B 0.019387f
C294 VTAIL.n104 B 0.008685f
C295 VTAIL.n105 B 0.008202f
C296 VTAIL.n106 B 0.015264f
C297 VTAIL.n107 B 0.015264f
C298 VTAIL.n108 B 0.008202f
C299 VTAIL.n109 B 0.008685f
C300 VTAIL.n110 B 0.019387f
C301 VTAIL.n111 B 0.019387f
C302 VTAIL.n112 B 0.008685f
C303 VTAIL.n113 B 0.008202f
C304 VTAIL.n114 B 0.015264f
C305 VTAIL.n115 B 0.015264f
C306 VTAIL.n116 B 0.008202f
C307 VTAIL.n117 B 0.008685f
C308 VTAIL.n118 B 0.019387f
C309 VTAIL.n119 B 0.019387f
C310 VTAIL.n120 B 0.039237f
C311 VTAIL.n121 B 0.008443f
C312 VTAIL.n122 B 0.008202f
C313 VTAIL.n123 B 0.037158f
C314 VTAIL.n124 B 0.02173f
C315 VTAIL.n125 B 0.767959f
C316 VTAIL.n126 B 0.01991f
C317 VTAIL.n127 B 0.015264f
C318 VTAIL.n128 B 0.008443f
C319 VTAIL.n129 B 0.019387f
C320 VTAIL.n130 B 0.008685f
C321 VTAIL.n131 B 0.015264f
C322 VTAIL.n132 B 0.008202f
C323 VTAIL.n133 B 0.019387f
C324 VTAIL.n134 B 0.008685f
C325 VTAIL.n135 B 0.015264f
C326 VTAIL.n136 B 0.008202f
C327 VTAIL.n137 B 0.01454f
C328 VTAIL.n138 B 0.013705f
C329 VTAIL.t3 B 0.032414f
C330 VTAIL.n139 B 0.085981f
C331 VTAIL.n140 B 0.490969f
C332 VTAIL.n141 B 0.008202f
C333 VTAIL.n142 B 0.008685f
C334 VTAIL.n143 B 0.019387f
C335 VTAIL.n144 B 0.019387f
C336 VTAIL.n145 B 0.008685f
C337 VTAIL.n146 B 0.008202f
C338 VTAIL.n147 B 0.015264f
C339 VTAIL.n148 B 0.015264f
C340 VTAIL.n149 B 0.008202f
C341 VTAIL.n150 B 0.008685f
C342 VTAIL.n151 B 0.019387f
C343 VTAIL.n152 B 0.019387f
C344 VTAIL.n153 B 0.008685f
C345 VTAIL.n154 B 0.008202f
C346 VTAIL.n155 B 0.015264f
C347 VTAIL.n156 B 0.015264f
C348 VTAIL.n157 B 0.008202f
C349 VTAIL.n158 B 0.008202f
C350 VTAIL.n159 B 0.008685f
C351 VTAIL.n160 B 0.019387f
C352 VTAIL.n161 B 0.019387f
C353 VTAIL.n162 B 0.039237f
C354 VTAIL.n163 B 0.008443f
C355 VTAIL.n164 B 0.008202f
C356 VTAIL.n165 B 0.037158f
C357 VTAIL.n166 B 0.02173f
C358 VTAIL.n167 B 0.710509f
C359 VN.t0 B 1.19112f
C360 VN.t1 B 1.49766f
.ends

