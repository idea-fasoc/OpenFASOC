* NGSPICE file created from diff_pair_sample_1213.ext - technology: sky130A

.subckt diff_pair_sample_1213 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.65835 pd=4.32 as=1.5561 ps=8.76 w=3.99 l=3.68
X1 VDD2.t5 VN.t0 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=0.65835 pd=4.32 as=1.5561 ps=8.76 w=3.99 l=3.68
X2 VDD2.t4 VN.t1 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=1.5561 pd=8.76 as=0.65835 ps=4.32 w=3.99 l=3.68
X3 VDD1.t4 VP.t1 VTAIL.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.5561 pd=8.76 as=0.65835 ps=4.32 w=3.99 l=3.68
X4 VDD1.t3 VP.t2 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=0.65835 pd=4.32 as=1.5561 ps=8.76 w=3.99 l=3.68
X5 VTAIL.t10 VN.t2 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.65835 pd=4.32 as=0.65835 ps=4.32 w=3.99 l=3.68
X6 VTAIL.t0 VP.t3 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.65835 pd=4.32 as=0.65835 ps=4.32 w=3.99 l=3.68
X7 VDD2.t2 VN.t3 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=0.65835 pd=4.32 as=1.5561 ps=8.76 w=3.99 l=3.68
X8 VDD2.t1 VN.t4 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=1.5561 pd=8.76 as=0.65835 ps=4.32 w=3.99 l=3.68
X9 VDD1.t1 VP.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.5561 pd=8.76 as=0.65835 ps=4.32 w=3.99 l=3.68
X10 VTAIL.t4 VP.t5 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.65835 pd=4.32 as=0.65835 ps=4.32 w=3.99 l=3.68
X11 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.68
X12 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.68
X13 VTAIL.t7 VN.t5 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.65835 pd=4.32 as=0.65835 ps=4.32 w=3.99 l=3.68
X14 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.68
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.68
R0 VP.n16 VP.n13 161.3
R1 VP.n18 VP.n17 161.3
R2 VP.n19 VP.n12 161.3
R3 VP.n21 VP.n20 161.3
R4 VP.n22 VP.n11 161.3
R5 VP.n24 VP.n23 161.3
R6 VP.n25 VP.n10 161.3
R7 VP.n27 VP.n26 161.3
R8 VP.n56 VP.n55 161.3
R9 VP.n54 VP.n1 161.3
R10 VP.n53 VP.n52 161.3
R11 VP.n51 VP.n2 161.3
R12 VP.n50 VP.n49 161.3
R13 VP.n48 VP.n3 161.3
R14 VP.n47 VP.n46 161.3
R15 VP.n45 VP.n4 161.3
R16 VP.n44 VP.n43 161.3
R17 VP.n42 VP.n5 161.3
R18 VP.n41 VP.n40 161.3
R19 VP.n39 VP.n6 161.3
R20 VP.n38 VP.n37 161.3
R21 VP.n36 VP.n7 161.3
R22 VP.n35 VP.n34 161.3
R23 VP.n33 VP.n8 161.3
R24 VP.n32 VP.n31 161.3
R25 VP.n30 VP.n29 89.5781
R26 VP.n57 VP.n0 89.5781
R27 VP.n28 VP.n9 89.5781
R28 VP.n15 VP.t4 58.3843
R29 VP.n15 VP.n14 50.4792
R30 VP.n29 VP.n28 46.8289
R31 VP.n37 VP.n36 40.979
R32 VP.n49 VP.n2 40.979
R33 VP.n20 VP.n11 40.979
R34 VP.n37 VP.n6 40.0078
R35 VP.n49 VP.n48 40.0078
R36 VP.n20 VP.n19 40.0078
R37 VP.n43 VP.t5 26.1307
R38 VP.n30 VP.t1 26.1307
R39 VP.n0 VP.t0 26.1307
R40 VP.n14 VP.t3 26.1307
R41 VP.n9 VP.t2 26.1307
R42 VP.n31 VP.n8 24.4675
R43 VP.n35 VP.n8 24.4675
R44 VP.n36 VP.n35 24.4675
R45 VP.n41 VP.n6 24.4675
R46 VP.n42 VP.n41 24.4675
R47 VP.n43 VP.n42 24.4675
R48 VP.n43 VP.n4 24.4675
R49 VP.n47 VP.n4 24.4675
R50 VP.n48 VP.n47 24.4675
R51 VP.n53 VP.n2 24.4675
R52 VP.n54 VP.n53 24.4675
R53 VP.n55 VP.n54 24.4675
R54 VP.n24 VP.n11 24.4675
R55 VP.n25 VP.n24 24.4675
R56 VP.n26 VP.n25 24.4675
R57 VP.n14 VP.n13 24.4675
R58 VP.n18 VP.n13 24.4675
R59 VP.n19 VP.n18 24.4675
R60 VP.n16 VP.n15 2.51577
R61 VP.n31 VP.n30 0.48984
R62 VP.n55 VP.n0 0.48984
R63 VP.n26 VP.n9 0.48984
R64 VP.n28 VP.n27 0.354971
R65 VP.n32 VP.n29 0.354971
R66 VP.n57 VP.n56 0.354971
R67 VP VP.n57 0.26696
R68 VP.n17 VP.n16 0.189894
R69 VP.n17 VP.n12 0.189894
R70 VP.n21 VP.n12 0.189894
R71 VP.n22 VP.n21 0.189894
R72 VP.n23 VP.n22 0.189894
R73 VP.n23 VP.n10 0.189894
R74 VP.n27 VP.n10 0.189894
R75 VP.n33 VP.n32 0.189894
R76 VP.n34 VP.n33 0.189894
R77 VP.n34 VP.n7 0.189894
R78 VP.n38 VP.n7 0.189894
R79 VP.n39 VP.n38 0.189894
R80 VP.n40 VP.n39 0.189894
R81 VP.n40 VP.n5 0.189894
R82 VP.n44 VP.n5 0.189894
R83 VP.n45 VP.n44 0.189894
R84 VP.n46 VP.n45 0.189894
R85 VP.n46 VP.n3 0.189894
R86 VP.n50 VP.n3 0.189894
R87 VP.n51 VP.n50 0.189894
R88 VP.n52 VP.n51 0.189894
R89 VP.n52 VP.n1 0.189894
R90 VP.n56 VP.n1 0.189894
R91 VTAIL.n82 VTAIL.n68 289.615
R92 VTAIL.n16 VTAIL.n2 289.615
R93 VTAIL.n62 VTAIL.n48 289.615
R94 VTAIL.n40 VTAIL.n26 289.615
R95 VTAIL.n75 VTAIL.n74 185
R96 VTAIL.n72 VTAIL.n71 185
R97 VTAIL.n81 VTAIL.n80 185
R98 VTAIL.n83 VTAIL.n82 185
R99 VTAIL.n9 VTAIL.n8 185
R100 VTAIL.n6 VTAIL.n5 185
R101 VTAIL.n15 VTAIL.n14 185
R102 VTAIL.n17 VTAIL.n16 185
R103 VTAIL.n63 VTAIL.n62 185
R104 VTAIL.n61 VTAIL.n60 185
R105 VTAIL.n52 VTAIL.n51 185
R106 VTAIL.n55 VTAIL.n54 185
R107 VTAIL.n41 VTAIL.n40 185
R108 VTAIL.n39 VTAIL.n38 185
R109 VTAIL.n30 VTAIL.n29 185
R110 VTAIL.n33 VTAIL.n32 185
R111 VTAIL.t9 VTAIL.n73 147.888
R112 VTAIL.t5 VTAIL.n7 147.888
R113 VTAIL.t2 VTAIL.n53 147.888
R114 VTAIL.t8 VTAIL.n31 147.888
R115 VTAIL.n74 VTAIL.n71 104.615
R116 VTAIL.n81 VTAIL.n71 104.615
R117 VTAIL.n82 VTAIL.n81 104.615
R118 VTAIL.n8 VTAIL.n5 104.615
R119 VTAIL.n15 VTAIL.n5 104.615
R120 VTAIL.n16 VTAIL.n15 104.615
R121 VTAIL.n62 VTAIL.n61 104.615
R122 VTAIL.n61 VTAIL.n51 104.615
R123 VTAIL.n54 VTAIL.n51 104.615
R124 VTAIL.n40 VTAIL.n39 104.615
R125 VTAIL.n39 VTAIL.n29 104.615
R126 VTAIL.n32 VTAIL.n29 104.615
R127 VTAIL.n47 VTAIL.n46 59.6944
R128 VTAIL.n25 VTAIL.n24 59.6944
R129 VTAIL.n1 VTAIL.n0 59.6943
R130 VTAIL.n23 VTAIL.n22 59.6943
R131 VTAIL.n74 VTAIL.t9 52.3082
R132 VTAIL.n8 VTAIL.t5 52.3082
R133 VTAIL.n54 VTAIL.t2 52.3082
R134 VTAIL.n32 VTAIL.t8 52.3082
R135 VTAIL.n87 VTAIL.n86 35.0944
R136 VTAIL.n21 VTAIL.n20 35.0944
R137 VTAIL.n67 VTAIL.n66 35.0944
R138 VTAIL.n45 VTAIL.n44 35.0944
R139 VTAIL.n25 VTAIL.n23 22.7203
R140 VTAIL.n87 VTAIL.n67 19.2634
R141 VTAIL.n75 VTAIL.n73 15.6496
R142 VTAIL.n9 VTAIL.n7 15.6496
R143 VTAIL.n55 VTAIL.n53 15.6496
R144 VTAIL.n33 VTAIL.n31 15.6496
R145 VTAIL.n76 VTAIL.n72 12.8005
R146 VTAIL.n10 VTAIL.n6 12.8005
R147 VTAIL.n56 VTAIL.n52 12.8005
R148 VTAIL.n34 VTAIL.n30 12.8005
R149 VTAIL.n80 VTAIL.n79 12.0247
R150 VTAIL.n14 VTAIL.n13 12.0247
R151 VTAIL.n60 VTAIL.n59 12.0247
R152 VTAIL.n38 VTAIL.n37 12.0247
R153 VTAIL.n83 VTAIL.n70 11.249
R154 VTAIL.n17 VTAIL.n4 11.249
R155 VTAIL.n63 VTAIL.n50 11.249
R156 VTAIL.n41 VTAIL.n28 11.249
R157 VTAIL.n84 VTAIL.n68 10.4732
R158 VTAIL.n18 VTAIL.n2 10.4732
R159 VTAIL.n64 VTAIL.n48 10.4732
R160 VTAIL.n42 VTAIL.n26 10.4732
R161 VTAIL.n86 VTAIL.n85 9.45567
R162 VTAIL.n20 VTAIL.n19 9.45567
R163 VTAIL.n66 VTAIL.n65 9.45567
R164 VTAIL.n44 VTAIL.n43 9.45567
R165 VTAIL.n85 VTAIL.n84 9.3005
R166 VTAIL.n70 VTAIL.n69 9.3005
R167 VTAIL.n79 VTAIL.n78 9.3005
R168 VTAIL.n77 VTAIL.n76 9.3005
R169 VTAIL.n19 VTAIL.n18 9.3005
R170 VTAIL.n4 VTAIL.n3 9.3005
R171 VTAIL.n13 VTAIL.n12 9.3005
R172 VTAIL.n11 VTAIL.n10 9.3005
R173 VTAIL.n65 VTAIL.n64 9.3005
R174 VTAIL.n50 VTAIL.n49 9.3005
R175 VTAIL.n59 VTAIL.n58 9.3005
R176 VTAIL.n57 VTAIL.n56 9.3005
R177 VTAIL.n43 VTAIL.n42 9.3005
R178 VTAIL.n28 VTAIL.n27 9.3005
R179 VTAIL.n37 VTAIL.n36 9.3005
R180 VTAIL.n35 VTAIL.n34 9.3005
R181 VTAIL.n0 VTAIL.t11 4.96291
R182 VTAIL.n0 VTAIL.t7 4.96291
R183 VTAIL.n22 VTAIL.t3 4.96291
R184 VTAIL.n22 VTAIL.t4 4.96291
R185 VTAIL.n46 VTAIL.t1 4.96291
R186 VTAIL.n46 VTAIL.t0 4.96291
R187 VTAIL.n24 VTAIL.t6 4.96291
R188 VTAIL.n24 VTAIL.t10 4.96291
R189 VTAIL.n77 VTAIL.n73 4.40546
R190 VTAIL.n11 VTAIL.n7 4.40546
R191 VTAIL.n57 VTAIL.n53 4.40546
R192 VTAIL.n35 VTAIL.n31 4.40546
R193 VTAIL.n86 VTAIL.n68 3.49141
R194 VTAIL.n20 VTAIL.n2 3.49141
R195 VTAIL.n66 VTAIL.n48 3.49141
R196 VTAIL.n44 VTAIL.n26 3.49141
R197 VTAIL.n45 VTAIL.n25 3.4574
R198 VTAIL.n67 VTAIL.n47 3.4574
R199 VTAIL.n23 VTAIL.n21 3.4574
R200 VTAIL.n84 VTAIL.n83 2.71565
R201 VTAIL.n18 VTAIL.n17 2.71565
R202 VTAIL.n64 VTAIL.n63 2.71565
R203 VTAIL.n42 VTAIL.n41 2.71565
R204 VTAIL VTAIL.n87 2.53498
R205 VTAIL.n47 VTAIL.n45 2.19878
R206 VTAIL.n21 VTAIL.n1 2.19878
R207 VTAIL.n80 VTAIL.n70 1.93989
R208 VTAIL.n14 VTAIL.n4 1.93989
R209 VTAIL.n60 VTAIL.n50 1.93989
R210 VTAIL.n38 VTAIL.n28 1.93989
R211 VTAIL.n79 VTAIL.n72 1.16414
R212 VTAIL.n13 VTAIL.n6 1.16414
R213 VTAIL.n59 VTAIL.n52 1.16414
R214 VTAIL.n37 VTAIL.n30 1.16414
R215 VTAIL VTAIL.n1 0.922914
R216 VTAIL.n76 VTAIL.n75 0.388379
R217 VTAIL.n10 VTAIL.n9 0.388379
R218 VTAIL.n56 VTAIL.n55 0.388379
R219 VTAIL.n34 VTAIL.n33 0.388379
R220 VTAIL.n78 VTAIL.n77 0.155672
R221 VTAIL.n78 VTAIL.n69 0.155672
R222 VTAIL.n85 VTAIL.n69 0.155672
R223 VTAIL.n12 VTAIL.n11 0.155672
R224 VTAIL.n12 VTAIL.n3 0.155672
R225 VTAIL.n19 VTAIL.n3 0.155672
R226 VTAIL.n65 VTAIL.n49 0.155672
R227 VTAIL.n58 VTAIL.n49 0.155672
R228 VTAIL.n58 VTAIL.n57 0.155672
R229 VTAIL.n43 VTAIL.n27 0.155672
R230 VTAIL.n36 VTAIL.n27 0.155672
R231 VTAIL.n36 VTAIL.n35 0.155672
R232 VDD1.n14 VDD1.n0 289.615
R233 VDD1.n33 VDD1.n19 289.615
R234 VDD1.n15 VDD1.n14 185
R235 VDD1.n13 VDD1.n12 185
R236 VDD1.n4 VDD1.n3 185
R237 VDD1.n7 VDD1.n6 185
R238 VDD1.n26 VDD1.n25 185
R239 VDD1.n23 VDD1.n22 185
R240 VDD1.n32 VDD1.n31 185
R241 VDD1.n34 VDD1.n33 185
R242 VDD1.t1 VDD1.n5 147.888
R243 VDD1.t4 VDD1.n24 147.888
R244 VDD1.n14 VDD1.n13 104.615
R245 VDD1.n13 VDD1.n3 104.615
R246 VDD1.n6 VDD1.n3 104.615
R247 VDD1.n25 VDD1.n22 104.615
R248 VDD1.n32 VDD1.n22 104.615
R249 VDD1.n33 VDD1.n32 104.615
R250 VDD1.n39 VDD1.n38 77.1819
R251 VDD1.n41 VDD1.n40 76.3731
R252 VDD1 VDD1.n18 54.4241
R253 VDD1.n39 VDD1.n37 54.3106
R254 VDD1.n6 VDD1.t1 52.3082
R255 VDD1.n25 VDD1.t4 52.3082
R256 VDD1.n41 VDD1.n39 40.7013
R257 VDD1.n7 VDD1.n5 15.6496
R258 VDD1.n26 VDD1.n24 15.6496
R259 VDD1.n8 VDD1.n4 12.8005
R260 VDD1.n27 VDD1.n23 12.8005
R261 VDD1.n12 VDD1.n11 12.0247
R262 VDD1.n31 VDD1.n30 12.0247
R263 VDD1.n15 VDD1.n2 11.249
R264 VDD1.n34 VDD1.n21 11.249
R265 VDD1.n16 VDD1.n0 10.4732
R266 VDD1.n35 VDD1.n19 10.4732
R267 VDD1.n18 VDD1.n17 9.45567
R268 VDD1.n37 VDD1.n36 9.45567
R269 VDD1.n17 VDD1.n16 9.3005
R270 VDD1.n2 VDD1.n1 9.3005
R271 VDD1.n11 VDD1.n10 9.3005
R272 VDD1.n9 VDD1.n8 9.3005
R273 VDD1.n36 VDD1.n35 9.3005
R274 VDD1.n21 VDD1.n20 9.3005
R275 VDD1.n30 VDD1.n29 9.3005
R276 VDD1.n28 VDD1.n27 9.3005
R277 VDD1.n40 VDD1.t2 4.96291
R278 VDD1.n40 VDD1.t3 4.96291
R279 VDD1.n38 VDD1.t0 4.96291
R280 VDD1.n38 VDD1.t5 4.96291
R281 VDD1.n9 VDD1.n5 4.40546
R282 VDD1.n28 VDD1.n24 4.40546
R283 VDD1.n18 VDD1.n0 3.49141
R284 VDD1.n37 VDD1.n19 3.49141
R285 VDD1.n16 VDD1.n15 2.71565
R286 VDD1.n35 VDD1.n34 2.71565
R287 VDD1.n12 VDD1.n2 1.93989
R288 VDD1.n31 VDD1.n21 1.93989
R289 VDD1.n11 VDD1.n4 1.16414
R290 VDD1.n30 VDD1.n23 1.16414
R291 VDD1 VDD1.n41 0.806535
R292 VDD1.n8 VDD1.n7 0.388379
R293 VDD1.n27 VDD1.n26 0.388379
R294 VDD1.n17 VDD1.n1 0.155672
R295 VDD1.n10 VDD1.n1 0.155672
R296 VDD1.n10 VDD1.n9 0.155672
R297 VDD1.n29 VDD1.n28 0.155672
R298 VDD1.n29 VDD1.n20 0.155672
R299 VDD1.n36 VDD1.n20 0.155672
R300 B.n681 B.n680 585
R301 B.n216 B.n124 585
R302 B.n215 B.n214 585
R303 B.n213 B.n212 585
R304 B.n211 B.n210 585
R305 B.n209 B.n208 585
R306 B.n207 B.n206 585
R307 B.n205 B.n204 585
R308 B.n203 B.n202 585
R309 B.n201 B.n200 585
R310 B.n199 B.n198 585
R311 B.n197 B.n196 585
R312 B.n195 B.n194 585
R313 B.n193 B.n192 585
R314 B.n191 B.n190 585
R315 B.n189 B.n188 585
R316 B.n187 B.n186 585
R317 B.n185 B.n184 585
R318 B.n183 B.n182 585
R319 B.n181 B.n180 585
R320 B.n179 B.n178 585
R321 B.n177 B.n176 585
R322 B.n175 B.n174 585
R323 B.n173 B.n172 585
R324 B.n171 B.n170 585
R325 B.n169 B.n168 585
R326 B.n167 B.n166 585
R327 B.n165 B.n164 585
R328 B.n163 B.n162 585
R329 B.n161 B.n160 585
R330 B.n159 B.n158 585
R331 B.n157 B.n156 585
R332 B.n155 B.n154 585
R333 B.n153 B.n152 585
R334 B.n151 B.n150 585
R335 B.n149 B.n148 585
R336 B.n147 B.n146 585
R337 B.n145 B.n144 585
R338 B.n143 B.n142 585
R339 B.n141 B.n140 585
R340 B.n139 B.n138 585
R341 B.n137 B.n136 585
R342 B.n135 B.n134 585
R343 B.n133 B.n132 585
R344 B.n102 B.n101 585
R345 B.n686 B.n685 585
R346 B.n679 B.n125 585
R347 B.n125 B.n99 585
R348 B.n678 B.n98 585
R349 B.n690 B.n98 585
R350 B.n677 B.n97 585
R351 B.n691 B.n97 585
R352 B.n676 B.n96 585
R353 B.n692 B.n96 585
R354 B.n675 B.n674 585
R355 B.n674 B.n92 585
R356 B.n673 B.n91 585
R357 B.n698 B.n91 585
R358 B.n672 B.n90 585
R359 B.n699 B.n90 585
R360 B.n671 B.n89 585
R361 B.n700 B.n89 585
R362 B.n670 B.n669 585
R363 B.n669 B.n85 585
R364 B.n668 B.n84 585
R365 B.n706 B.n84 585
R366 B.n667 B.n83 585
R367 B.n707 B.n83 585
R368 B.n666 B.n82 585
R369 B.n708 B.n82 585
R370 B.n665 B.n664 585
R371 B.n664 B.n78 585
R372 B.n663 B.n77 585
R373 B.n714 B.n77 585
R374 B.n662 B.n76 585
R375 B.n715 B.n76 585
R376 B.n661 B.n75 585
R377 B.n716 B.n75 585
R378 B.n660 B.n659 585
R379 B.n659 B.n71 585
R380 B.n658 B.n70 585
R381 B.n722 B.n70 585
R382 B.n657 B.n69 585
R383 B.n723 B.n69 585
R384 B.n656 B.n68 585
R385 B.n724 B.n68 585
R386 B.n655 B.n654 585
R387 B.n654 B.n64 585
R388 B.n653 B.n63 585
R389 B.n730 B.n63 585
R390 B.n652 B.n62 585
R391 B.n731 B.n62 585
R392 B.n651 B.n61 585
R393 B.n732 B.n61 585
R394 B.n650 B.n649 585
R395 B.n649 B.n60 585
R396 B.n648 B.n56 585
R397 B.n738 B.n56 585
R398 B.n647 B.n55 585
R399 B.n739 B.n55 585
R400 B.n646 B.n54 585
R401 B.n740 B.n54 585
R402 B.n645 B.n644 585
R403 B.n644 B.n50 585
R404 B.n643 B.n49 585
R405 B.n746 B.n49 585
R406 B.n642 B.n48 585
R407 B.n747 B.n48 585
R408 B.n641 B.n47 585
R409 B.n748 B.n47 585
R410 B.n640 B.n639 585
R411 B.n639 B.n43 585
R412 B.n638 B.n42 585
R413 B.n754 B.n42 585
R414 B.n637 B.n41 585
R415 B.n755 B.n41 585
R416 B.n636 B.n40 585
R417 B.n756 B.n40 585
R418 B.n635 B.n634 585
R419 B.n634 B.n39 585
R420 B.n633 B.n35 585
R421 B.n762 B.n35 585
R422 B.n632 B.n34 585
R423 B.n763 B.n34 585
R424 B.n631 B.n33 585
R425 B.n764 B.n33 585
R426 B.n630 B.n629 585
R427 B.n629 B.n29 585
R428 B.n628 B.n28 585
R429 B.n770 B.n28 585
R430 B.n627 B.n27 585
R431 B.n771 B.n27 585
R432 B.n626 B.n26 585
R433 B.n772 B.n26 585
R434 B.n625 B.n624 585
R435 B.n624 B.n22 585
R436 B.n623 B.n21 585
R437 B.n778 B.n21 585
R438 B.n622 B.n20 585
R439 B.n779 B.n20 585
R440 B.n621 B.n19 585
R441 B.n780 B.n19 585
R442 B.n620 B.n619 585
R443 B.n619 B.t1 585
R444 B.n618 B.n15 585
R445 B.n786 B.n15 585
R446 B.n617 B.n14 585
R447 B.n787 B.n14 585
R448 B.n616 B.n13 585
R449 B.n788 B.n13 585
R450 B.n615 B.n614 585
R451 B.n614 B.n12 585
R452 B.n613 B.n612 585
R453 B.n613 B.n8 585
R454 B.n611 B.n7 585
R455 B.n795 B.n7 585
R456 B.n610 B.n6 585
R457 B.n796 B.n6 585
R458 B.n609 B.n5 585
R459 B.n797 B.n5 585
R460 B.n608 B.n607 585
R461 B.n607 B.n4 585
R462 B.n606 B.n217 585
R463 B.n606 B.n605 585
R464 B.n596 B.n218 585
R465 B.n219 B.n218 585
R466 B.n598 B.n597 585
R467 B.n599 B.n598 585
R468 B.n595 B.n224 585
R469 B.n224 B.n223 585
R470 B.n594 B.n593 585
R471 B.n593 B.n592 585
R472 B.n226 B.n225 585
R473 B.t5 B.n226 585
R474 B.n585 B.n584 585
R475 B.n586 B.n585 585
R476 B.n583 B.n231 585
R477 B.n231 B.n230 585
R478 B.n582 B.n581 585
R479 B.n581 B.n580 585
R480 B.n233 B.n232 585
R481 B.n234 B.n233 585
R482 B.n573 B.n572 585
R483 B.n574 B.n573 585
R484 B.n571 B.n239 585
R485 B.n239 B.n238 585
R486 B.n570 B.n569 585
R487 B.n569 B.n568 585
R488 B.n241 B.n240 585
R489 B.n242 B.n241 585
R490 B.n561 B.n560 585
R491 B.n562 B.n561 585
R492 B.n559 B.n247 585
R493 B.n247 B.n246 585
R494 B.n558 B.n557 585
R495 B.n557 B.n556 585
R496 B.n249 B.n248 585
R497 B.n549 B.n249 585
R498 B.n548 B.n547 585
R499 B.n550 B.n548 585
R500 B.n546 B.n254 585
R501 B.n254 B.n253 585
R502 B.n545 B.n544 585
R503 B.n544 B.n543 585
R504 B.n256 B.n255 585
R505 B.n257 B.n256 585
R506 B.n536 B.n535 585
R507 B.n537 B.n536 585
R508 B.n534 B.n262 585
R509 B.n262 B.n261 585
R510 B.n533 B.n532 585
R511 B.n532 B.n531 585
R512 B.n264 B.n263 585
R513 B.n265 B.n264 585
R514 B.n524 B.n523 585
R515 B.n525 B.n524 585
R516 B.n522 B.n270 585
R517 B.n270 B.n269 585
R518 B.n521 B.n520 585
R519 B.n520 B.n519 585
R520 B.n272 B.n271 585
R521 B.n512 B.n272 585
R522 B.n511 B.n510 585
R523 B.n513 B.n511 585
R524 B.n509 B.n277 585
R525 B.n277 B.n276 585
R526 B.n508 B.n507 585
R527 B.n507 B.n506 585
R528 B.n279 B.n278 585
R529 B.n280 B.n279 585
R530 B.n499 B.n498 585
R531 B.n500 B.n499 585
R532 B.n497 B.n285 585
R533 B.n285 B.n284 585
R534 B.n496 B.n495 585
R535 B.n495 B.n494 585
R536 B.n287 B.n286 585
R537 B.n288 B.n287 585
R538 B.n487 B.n486 585
R539 B.n488 B.n487 585
R540 B.n485 B.n293 585
R541 B.n293 B.n292 585
R542 B.n484 B.n483 585
R543 B.n483 B.n482 585
R544 B.n295 B.n294 585
R545 B.n296 B.n295 585
R546 B.n475 B.n474 585
R547 B.n476 B.n475 585
R548 B.n473 B.n301 585
R549 B.n301 B.n300 585
R550 B.n472 B.n471 585
R551 B.n471 B.n470 585
R552 B.n303 B.n302 585
R553 B.n304 B.n303 585
R554 B.n463 B.n462 585
R555 B.n464 B.n463 585
R556 B.n461 B.n309 585
R557 B.n309 B.n308 585
R558 B.n460 B.n459 585
R559 B.n459 B.n458 585
R560 B.n311 B.n310 585
R561 B.n312 B.n311 585
R562 B.n451 B.n450 585
R563 B.n452 B.n451 585
R564 B.n449 B.n317 585
R565 B.n317 B.n316 585
R566 B.n448 B.n447 585
R567 B.n447 B.n446 585
R568 B.n319 B.n318 585
R569 B.n320 B.n319 585
R570 B.n442 B.n441 585
R571 B.n323 B.n322 585
R572 B.n438 B.n437 585
R573 B.n439 B.n438 585
R574 B.n436 B.n346 585
R575 B.n435 B.n434 585
R576 B.n433 B.n432 585
R577 B.n431 B.n430 585
R578 B.n429 B.n428 585
R579 B.n427 B.n426 585
R580 B.n425 B.n424 585
R581 B.n423 B.n422 585
R582 B.n421 B.n420 585
R583 B.n419 B.n418 585
R584 B.n417 B.n416 585
R585 B.n415 B.n414 585
R586 B.n413 B.n412 585
R587 B.n411 B.n410 585
R588 B.n409 B.n408 585
R589 B.n406 B.n405 585
R590 B.n404 B.n403 585
R591 B.n402 B.n401 585
R592 B.n400 B.n399 585
R593 B.n398 B.n397 585
R594 B.n396 B.n395 585
R595 B.n394 B.n393 585
R596 B.n392 B.n391 585
R597 B.n390 B.n389 585
R598 B.n388 B.n387 585
R599 B.n385 B.n384 585
R600 B.n383 B.n382 585
R601 B.n381 B.n380 585
R602 B.n379 B.n378 585
R603 B.n377 B.n376 585
R604 B.n375 B.n374 585
R605 B.n373 B.n372 585
R606 B.n371 B.n370 585
R607 B.n369 B.n368 585
R608 B.n367 B.n366 585
R609 B.n365 B.n364 585
R610 B.n363 B.n362 585
R611 B.n361 B.n360 585
R612 B.n359 B.n358 585
R613 B.n357 B.n356 585
R614 B.n355 B.n354 585
R615 B.n353 B.n352 585
R616 B.n351 B.n345 585
R617 B.n439 B.n345 585
R618 B.n443 B.n321 585
R619 B.n321 B.n320 585
R620 B.n445 B.n444 585
R621 B.n446 B.n445 585
R622 B.n315 B.n314 585
R623 B.n316 B.n315 585
R624 B.n454 B.n453 585
R625 B.n453 B.n452 585
R626 B.n455 B.n313 585
R627 B.n313 B.n312 585
R628 B.n457 B.n456 585
R629 B.n458 B.n457 585
R630 B.n307 B.n306 585
R631 B.n308 B.n307 585
R632 B.n466 B.n465 585
R633 B.n465 B.n464 585
R634 B.n467 B.n305 585
R635 B.n305 B.n304 585
R636 B.n469 B.n468 585
R637 B.n470 B.n469 585
R638 B.n299 B.n298 585
R639 B.n300 B.n299 585
R640 B.n478 B.n477 585
R641 B.n477 B.n476 585
R642 B.n479 B.n297 585
R643 B.n297 B.n296 585
R644 B.n481 B.n480 585
R645 B.n482 B.n481 585
R646 B.n291 B.n290 585
R647 B.n292 B.n291 585
R648 B.n490 B.n489 585
R649 B.n489 B.n488 585
R650 B.n491 B.n289 585
R651 B.n289 B.n288 585
R652 B.n493 B.n492 585
R653 B.n494 B.n493 585
R654 B.n283 B.n282 585
R655 B.n284 B.n283 585
R656 B.n502 B.n501 585
R657 B.n501 B.n500 585
R658 B.n503 B.n281 585
R659 B.n281 B.n280 585
R660 B.n505 B.n504 585
R661 B.n506 B.n505 585
R662 B.n275 B.n274 585
R663 B.n276 B.n275 585
R664 B.n515 B.n514 585
R665 B.n514 B.n513 585
R666 B.n516 B.n273 585
R667 B.n512 B.n273 585
R668 B.n518 B.n517 585
R669 B.n519 B.n518 585
R670 B.n268 B.n267 585
R671 B.n269 B.n268 585
R672 B.n527 B.n526 585
R673 B.n526 B.n525 585
R674 B.n528 B.n266 585
R675 B.n266 B.n265 585
R676 B.n530 B.n529 585
R677 B.n531 B.n530 585
R678 B.n260 B.n259 585
R679 B.n261 B.n260 585
R680 B.n539 B.n538 585
R681 B.n538 B.n537 585
R682 B.n540 B.n258 585
R683 B.n258 B.n257 585
R684 B.n542 B.n541 585
R685 B.n543 B.n542 585
R686 B.n252 B.n251 585
R687 B.n253 B.n252 585
R688 B.n552 B.n551 585
R689 B.n551 B.n550 585
R690 B.n553 B.n250 585
R691 B.n549 B.n250 585
R692 B.n555 B.n554 585
R693 B.n556 B.n555 585
R694 B.n245 B.n244 585
R695 B.n246 B.n245 585
R696 B.n564 B.n563 585
R697 B.n563 B.n562 585
R698 B.n565 B.n243 585
R699 B.n243 B.n242 585
R700 B.n567 B.n566 585
R701 B.n568 B.n567 585
R702 B.n237 B.n236 585
R703 B.n238 B.n237 585
R704 B.n576 B.n575 585
R705 B.n575 B.n574 585
R706 B.n577 B.n235 585
R707 B.n235 B.n234 585
R708 B.n579 B.n578 585
R709 B.n580 B.n579 585
R710 B.n229 B.n228 585
R711 B.n230 B.n229 585
R712 B.n588 B.n587 585
R713 B.n587 B.n586 585
R714 B.n589 B.n227 585
R715 B.n227 B.t5 585
R716 B.n591 B.n590 585
R717 B.n592 B.n591 585
R718 B.n222 B.n221 585
R719 B.n223 B.n222 585
R720 B.n601 B.n600 585
R721 B.n600 B.n599 585
R722 B.n602 B.n220 585
R723 B.n220 B.n219 585
R724 B.n604 B.n603 585
R725 B.n605 B.n604 585
R726 B.n3 B.n0 585
R727 B.n4 B.n3 585
R728 B.n794 B.n1 585
R729 B.n795 B.n794 585
R730 B.n793 B.n792 585
R731 B.n793 B.n8 585
R732 B.n791 B.n9 585
R733 B.n12 B.n9 585
R734 B.n790 B.n789 585
R735 B.n789 B.n788 585
R736 B.n11 B.n10 585
R737 B.n787 B.n11 585
R738 B.n785 B.n784 585
R739 B.n786 B.n785 585
R740 B.n783 B.n16 585
R741 B.n16 B.t1 585
R742 B.n782 B.n781 585
R743 B.n781 B.n780 585
R744 B.n18 B.n17 585
R745 B.n779 B.n18 585
R746 B.n777 B.n776 585
R747 B.n778 B.n777 585
R748 B.n775 B.n23 585
R749 B.n23 B.n22 585
R750 B.n774 B.n773 585
R751 B.n773 B.n772 585
R752 B.n25 B.n24 585
R753 B.n771 B.n25 585
R754 B.n769 B.n768 585
R755 B.n770 B.n769 585
R756 B.n767 B.n30 585
R757 B.n30 B.n29 585
R758 B.n766 B.n765 585
R759 B.n765 B.n764 585
R760 B.n32 B.n31 585
R761 B.n763 B.n32 585
R762 B.n761 B.n760 585
R763 B.n762 B.n761 585
R764 B.n759 B.n36 585
R765 B.n39 B.n36 585
R766 B.n758 B.n757 585
R767 B.n757 B.n756 585
R768 B.n38 B.n37 585
R769 B.n755 B.n38 585
R770 B.n753 B.n752 585
R771 B.n754 B.n753 585
R772 B.n751 B.n44 585
R773 B.n44 B.n43 585
R774 B.n750 B.n749 585
R775 B.n749 B.n748 585
R776 B.n46 B.n45 585
R777 B.n747 B.n46 585
R778 B.n745 B.n744 585
R779 B.n746 B.n745 585
R780 B.n743 B.n51 585
R781 B.n51 B.n50 585
R782 B.n742 B.n741 585
R783 B.n741 B.n740 585
R784 B.n53 B.n52 585
R785 B.n739 B.n53 585
R786 B.n737 B.n736 585
R787 B.n738 B.n737 585
R788 B.n735 B.n57 585
R789 B.n60 B.n57 585
R790 B.n734 B.n733 585
R791 B.n733 B.n732 585
R792 B.n59 B.n58 585
R793 B.n731 B.n59 585
R794 B.n729 B.n728 585
R795 B.n730 B.n729 585
R796 B.n727 B.n65 585
R797 B.n65 B.n64 585
R798 B.n726 B.n725 585
R799 B.n725 B.n724 585
R800 B.n67 B.n66 585
R801 B.n723 B.n67 585
R802 B.n721 B.n720 585
R803 B.n722 B.n721 585
R804 B.n719 B.n72 585
R805 B.n72 B.n71 585
R806 B.n718 B.n717 585
R807 B.n717 B.n716 585
R808 B.n74 B.n73 585
R809 B.n715 B.n74 585
R810 B.n713 B.n712 585
R811 B.n714 B.n713 585
R812 B.n711 B.n79 585
R813 B.n79 B.n78 585
R814 B.n710 B.n709 585
R815 B.n709 B.n708 585
R816 B.n81 B.n80 585
R817 B.n707 B.n81 585
R818 B.n705 B.n704 585
R819 B.n706 B.n705 585
R820 B.n703 B.n86 585
R821 B.n86 B.n85 585
R822 B.n702 B.n701 585
R823 B.n701 B.n700 585
R824 B.n88 B.n87 585
R825 B.n699 B.n88 585
R826 B.n697 B.n696 585
R827 B.n698 B.n697 585
R828 B.n695 B.n93 585
R829 B.n93 B.n92 585
R830 B.n694 B.n693 585
R831 B.n693 B.n692 585
R832 B.n95 B.n94 585
R833 B.n691 B.n95 585
R834 B.n689 B.n688 585
R835 B.n690 B.n689 585
R836 B.n687 B.n100 585
R837 B.n100 B.n99 585
R838 B.n798 B.n797 585
R839 B.n796 B.n2 585
R840 B.n685 B.n100 439.647
R841 B.n681 B.n125 439.647
R842 B.n345 B.n319 439.647
R843 B.n441 B.n321 439.647
R844 B.n683 B.n682 256.663
R845 B.n683 B.n123 256.663
R846 B.n683 B.n122 256.663
R847 B.n683 B.n121 256.663
R848 B.n683 B.n120 256.663
R849 B.n683 B.n119 256.663
R850 B.n683 B.n118 256.663
R851 B.n683 B.n117 256.663
R852 B.n683 B.n116 256.663
R853 B.n683 B.n115 256.663
R854 B.n683 B.n114 256.663
R855 B.n683 B.n113 256.663
R856 B.n683 B.n112 256.663
R857 B.n683 B.n111 256.663
R858 B.n683 B.n110 256.663
R859 B.n683 B.n109 256.663
R860 B.n683 B.n108 256.663
R861 B.n683 B.n107 256.663
R862 B.n683 B.n106 256.663
R863 B.n683 B.n105 256.663
R864 B.n683 B.n104 256.663
R865 B.n683 B.n103 256.663
R866 B.n684 B.n683 256.663
R867 B.n440 B.n439 256.663
R868 B.n439 B.n324 256.663
R869 B.n439 B.n325 256.663
R870 B.n439 B.n326 256.663
R871 B.n439 B.n327 256.663
R872 B.n439 B.n328 256.663
R873 B.n439 B.n329 256.663
R874 B.n439 B.n330 256.663
R875 B.n439 B.n331 256.663
R876 B.n439 B.n332 256.663
R877 B.n439 B.n333 256.663
R878 B.n439 B.n334 256.663
R879 B.n439 B.n335 256.663
R880 B.n439 B.n336 256.663
R881 B.n439 B.n337 256.663
R882 B.n439 B.n338 256.663
R883 B.n439 B.n339 256.663
R884 B.n439 B.n340 256.663
R885 B.n439 B.n341 256.663
R886 B.n439 B.n342 256.663
R887 B.n439 B.n343 256.663
R888 B.n439 B.n344 256.663
R889 B.n800 B.n799 256.663
R890 B.n129 B.t14 235.379
R891 B.n126 B.t6 235.379
R892 B.n349 B.t17 235.379
R893 B.n347 B.t10 235.379
R894 B.n126 B.t8 222.835
R895 B.n349 B.t19 222.835
R896 B.n129 B.t15 222.835
R897 B.n347 B.t13 222.835
R898 B.n132 B.n102 163.367
R899 B.n136 B.n135 163.367
R900 B.n140 B.n139 163.367
R901 B.n144 B.n143 163.367
R902 B.n148 B.n147 163.367
R903 B.n152 B.n151 163.367
R904 B.n156 B.n155 163.367
R905 B.n160 B.n159 163.367
R906 B.n164 B.n163 163.367
R907 B.n168 B.n167 163.367
R908 B.n172 B.n171 163.367
R909 B.n176 B.n175 163.367
R910 B.n180 B.n179 163.367
R911 B.n184 B.n183 163.367
R912 B.n188 B.n187 163.367
R913 B.n192 B.n191 163.367
R914 B.n196 B.n195 163.367
R915 B.n200 B.n199 163.367
R916 B.n204 B.n203 163.367
R917 B.n208 B.n207 163.367
R918 B.n212 B.n211 163.367
R919 B.n214 B.n124 163.367
R920 B.n447 B.n319 163.367
R921 B.n447 B.n317 163.367
R922 B.n451 B.n317 163.367
R923 B.n451 B.n311 163.367
R924 B.n459 B.n311 163.367
R925 B.n459 B.n309 163.367
R926 B.n463 B.n309 163.367
R927 B.n463 B.n303 163.367
R928 B.n471 B.n303 163.367
R929 B.n471 B.n301 163.367
R930 B.n475 B.n301 163.367
R931 B.n475 B.n295 163.367
R932 B.n483 B.n295 163.367
R933 B.n483 B.n293 163.367
R934 B.n487 B.n293 163.367
R935 B.n487 B.n287 163.367
R936 B.n495 B.n287 163.367
R937 B.n495 B.n285 163.367
R938 B.n499 B.n285 163.367
R939 B.n499 B.n279 163.367
R940 B.n507 B.n279 163.367
R941 B.n507 B.n277 163.367
R942 B.n511 B.n277 163.367
R943 B.n511 B.n272 163.367
R944 B.n520 B.n272 163.367
R945 B.n520 B.n270 163.367
R946 B.n524 B.n270 163.367
R947 B.n524 B.n264 163.367
R948 B.n532 B.n264 163.367
R949 B.n532 B.n262 163.367
R950 B.n536 B.n262 163.367
R951 B.n536 B.n256 163.367
R952 B.n544 B.n256 163.367
R953 B.n544 B.n254 163.367
R954 B.n548 B.n254 163.367
R955 B.n548 B.n249 163.367
R956 B.n557 B.n249 163.367
R957 B.n557 B.n247 163.367
R958 B.n561 B.n247 163.367
R959 B.n561 B.n241 163.367
R960 B.n569 B.n241 163.367
R961 B.n569 B.n239 163.367
R962 B.n573 B.n239 163.367
R963 B.n573 B.n233 163.367
R964 B.n581 B.n233 163.367
R965 B.n581 B.n231 163.367
R966 B.n585 B.n231 163.367
R967 B.n585 B.n226 163.367
R968 B.n593 B.n226 163.367
R969 B.n593 B.n224 163.367
R970 B.n598 B.n224 163.367
R971 B.n598 B.n218 163.367
R972 B.n606 B.n218 163.367
R973 B.n607 B.n606 163.367
R974 B.n607 B.n5 163.367
R975 B.n6 B.n5 163.367
R976 B.n7 B.n6 163.367
R977 B.n613 B.n7 163.367
R978 B.n614 B.n613 163.367
R979 B.n614 B.n13 163.367
R980 B.n14 B.n13 163.367
R981 B.n15 B.n14 163.367
R982 B.n619 B.n15 163.367
R983 B.n619 B.n19 163.367
R984 B.n20 B.n19 163.367
R985 B.n21 B.n20 163.367
R986 B.n624 B.n21 163.367
R987 B.n624 B.n26 163.367
R988 B.n27 B.n26 163.367
R989 B.n28 B.n27 163.367
R990 B.n629 B.n28 163.367
R991 B.n629 B.n33 163.367
R992 B.n34 B.n33 163.367
R993 B.n35 B.n34 163.367
R994 B.n634 B.n35 163.367
R995 B.n634 B.n40 163.367
R996 B.n41 B.n40 163.367
R997 B.n42 B.n41 163.367
R998 B.n639 B.n42 163.367
R999 B.n639 B.n47 163.367
R1000 B.n48 B.n47 163.367
R1001 B.n49 B.n48 163.367
R1002 B.n644 B.n49 163.367
R1003 B.n644 B.n54 163.367
R1004 B.n55 B.n54 163.367
R1005 B.n56 B.n55 163.367
R1006 B.n649 B.n56 163.367
R1007 B.n649 B.n61 163.367
R1008 B.n62 B.n61 163.367
R1009 B.n63 B.n62 163.367
R1010 B.n654 B.n63 163.367
R1011 B.n654 B.n68 163.367
R1012 B.n69 B.n68 163.367
R1013 B.n70 B.n69 163.367
R1014 B.n659 B.n70 163.367
R1015 B.n659 B.n75 163.367
R1016 B.n76 B.n75 163.367
R1017 B.n77 B.n76 163.367
R1018 B.n664 B.n77 163.367
R1019 B.n664 B.n82 163.367
R1020 B.n83 B.n82 163.367
R1021 B.n84 B.n83 163.367
R1022 B.n669 B.n84 163.367
R1023 B.n669 B.n89 163.367
R1024 B.n90 B.n89 163.367
R1025 B.n91 B.n90 163.367
R1026 B.n674 B.n91 163.367
R1027 B.n674 B.n96 163.367
R1028 B.n97 B.n96 163.367
R1029 B.n98 B.n97 163.367
R1030 B.n125 B.n98 163.367
R1031 B.n438 B.n323 163.367
R1032 B.n438 B.n346 163.367
R1033 B.n434 B.n433 163.367
R1034 B.n430 B.n429 163.367
R1035 B.n426 B.n425 163.367
R1036 B.n422 B.n421 163.367
R1037 B.n418 B.n417 163.367
R1038 B.n414 B.n413 163.367
R1039 B.n410 B.n409 163.367
R1040 B.n405 B.n404 163.367
R1041 B.n401 B.n400 163.367
R1042 B.n397 B.n396 163.367
R1043 B.n393 B.n392 163.367
R1044 B.n389 B.n388 163.367
R1045 B.n384 B.n383 163.367
R1046 B.n380 B.n379 163.367
R1047 B.n376 B.n375 163.367
R1048 B.n372 B.n371 163.367
R1049 B.n368 B.n367 163.367
R1050 B.n364 B.n363 163.367
R1051 B.n360 B.n359 163.367
R1052 B.n356 B.n355 163.367
R1053 B.n352 B.n345 163.367
R1054 B.n445 B.n321 163.367
R1055 B.n445 B.n315 163.367
R1056 B.n453 B.n315 163.367
R1057 B.n453 B.n313 163.367
R1058 B.n457 B.n313 163.367
R1059 B.n457 B.n307 163.367
R1060 B.n465 B.n307 163.367
R1061 B.n465 B.n305 163.367
R1062 B.n469 B.n305 163.367
R1063 B.n469 B.n299 163.367
R1064 B.n477 B.n299 163.367
R1065 B.n477 B.n297 163.367
R1066 B.n481 B.n297 163.367
R1067 B.n481 B.n291 163.367
R1068 B.n489 B.n291 163.367
R1069 B.n489 B.n289 163.367
R1070 B.n493 B.n289 163.367
R1071 B.n493 B.n283 163.367
R1072 B.n501 B.n283 163.367
R1073 B.n501 B.n281 163.367
R1074 B.n505 B.n281 163.367
R1075 B.n505 B.n275 163.367
R1076 B.n514 B.n275 163.367
R1077 B.n514 B.n273 163.367
R1078 B.n518 B.n273 163.367
R1079 B.n518 B.n268 163.367
R1080 B.n526 B.n268 163.367
R1081 B.n526 B.n266 163.367
R1082 B.n530 B.n266 163.367
R1083 B.n530 B.n260 163.367
R1084 B.n538 B.n260 163.367
R1085 B.n538 B.n258 163.367
R1086 B.n542 B.n258 163.367
R1087 B.n542 B.n252 163.367
R1088 B.n551 B.n252 163.367
R1089 B.n551 B.n250 163.367
R1090 B.n555 B.n250 163.367
R1091 B.n555 B.n245 163.367
R1092 B.n563 B.n245 163.367
R1093 B.n563 B.n243 163.367
R1094 B.n567 B.n243 163.367
R1095 B.n567 B.n237 163.367
R1096 B.n575 B.n237 163.367
R1097 B.n575 B.n235 163.367
R1098 B.n579 B.n235 163.367
R1099 B.n579 B.n229 163.367
R1100 B.n587 B.n229 163.367
R1101 B.n587 B.n227 163.367
R1102 B.n591 B.n227 163.367
R1103 B.n591 B.n222 163.367
R1104 B.n600 B.n222 163.367
R1105 B.n600 B.n220 163.367
R1106 B.n604 B.n220 163.367
R1107 B.n604 B.n3 163.367
R1108 B.n798 B.n3 163.367
R1109 B.n794 B.n2 163.367
R1110 B.n794 B.n793 163.367
R1111 B.n793 B.n9 163.367
R1112 B.n789 B.n9 163.367
R1113 B.n789 B.n11 163.367
R1114 B.n785 B.n11 163.367
R1115 B.n785 B.n16 163.367
R1116 B.n781 B.n16 163.367
R1117 B.n781 B.n18 163.367
R1118 B.n777 B.n18 163.367
R1119 B.n777 B.n23 163.367
R1120 B.n773 B.n23 163.367
R1121 B.n773 B.n25 163.367
R1122 B.n769 B.n25 163.367
R1123 B.n769 B.n30 163.367
R1124 B.n765 B.n30 163.367
R1125 B.n765 B.n32 163.367
R1126 B.n761 B.n32 163.367
R1127 B.n761 B.n36 163.367
R1128 B.n757 B.n36 163.367
R1129 B.n757 B.n38 163.367
R1130 B.n753 B.n38 163.367
R1131 B.n753 B.n44 163.367
R1132 B.n749 B.n44 163.367
R1133 B.n749 B.n46 163.367
R1134 B.n745 B.n46 163.367
R1135 B.n745 B.n51 163.367
R1136 B.n741 B.n51 163.367
R1137 B.n741 B.n53 163.367
R1138 B.n737 B.n53 163.367
R1139 B.n737 B.n57 163.367
R1140 B.n733 B.n57 163.367
R1141 B.n733 B.n59 163.367
R1142 B.n729 B.n59 163.367
R1143 B.n729 B.n65 163.367
R1144 B.n725 B.n65 163.367
R1145 B.n725 B.n67 163.367
R1146 B.n721 B.n67 163.367
R1147 B.n721 B.n72 163.367
R1148 B.n717 B.n72 163.367
R1149 B.n717 B.n74 163.367
R1150 B.n713 B.n74 163.367
R1151 B.n713 B.n79 163.367
R1152 B.n709 B.n79 163.367
R1153 B.n709 B.n81 163.367
R1154 B.n705 B.n81 163.367
R1155 B.n705 B.n86 163.367
R1156 B.n701 B.n86 163.367
R1157 B.n701 B.n88 163.367
R1158 B.n697 B.n88 163.367
R1159 B.n697 B.n93 163.367
R1160 B.n693 B.n93 163.367
R1161 B.n693 B.n95 163.367
R1162 B.n689 B.n95 163.367
R1163 B.n689 B.n100 163.367
R1164 B.n127 B.t9 145.066
R1165 B.n350 B.t18 145.066
R1166 B.n130 B.t16 145.066
R1167 B.n348 B.t12 145.066
R1168 B.n439 B.n320 129.412
R1169 B.n683 B.n99 129.412
R1170 B.n446 B.n320 80.7344
R1171 B.n446 B.n316 80.7344
R1172 B.n452 B.n316 80.7344
R1173 B.n452 B.n312 80.7344
R1174 B.n458 B.n312 80.7344
R1175 B.n458 B.n308 80.7344
R1176 B.n464 B.n308 80.7344
R1177 B.n464 B.n304 80.7344
R1178 B.n470 B.n304 80.7344
R1179 B.n476 B.n300 80.7344
R1180 B.n476 B.n296 80.7344
R1181 B.n482 B.n296 80.7344
R1182 B.n482 B.n292 80.7344
R1183 B.n488 B.n292 80.7344
R1184 B.n488 B.n288 80.7344
R1185 B.n494 B.n288 80.7344
R1186 B.n494 B.n284 80.7344
R1187 B.n500 B.n284 80.7344
R1188 B.n500 B.n280 80.7344
R1189 B.n506 B.n280 80.7344
R1190 B.n506 B.n276 80.7344
R1191 B.n513 B.n276 80.7344
R1192 B.n513 B.n512 80.7344
R1193 B.n519 B.n269 80.7344
R1194 B.n525 B.n269 80.7344
R1195 B.n525 B.n265 80.7344
R1196 B.n531 B.n265 80.7344
R1197 B.n531 B.n261 80.7344
R1198 B.n537 B.n261 80.7344
R1199 B.n537 B.n257 80.7344
R1200 B.n543 B.n257 80.7344
R1201 B.n543 B.n253 80.7344
R1202 B.n550 B.n253 80.7344
R1203 B.n550 B.n549 80.7344
R1204 B.n556 B.n246 80.7344
R1205 B.n562 B.n246 80.7344
R1206 B.n562 B.n242 80.7344
R1207 B.n568 B.n242 80.7344
R1208 B.n568 B.n238 80.7344
R1209 B.n574 B.n238 80.7344
R1210 B.n574 B.n234 80.7344
R1211 B.n580 B.n234 80.7344
R1212 B.n580 B.n230 80.7344
R1213 B.n586 B.n230 80.7344
R1214 B.n586 B.t5 80.7344
R1215 B.n592 B.t5 80.7344
R1216 B.n592 B.n223 80.7344
R1217 B.n599 B.n223 80.7344
R1218 B.n599 B.n219 80.7344
R1219 B.n605 B.n219 80.7344
R1220 B.n605 B.n4 80.7344
R1221 B.n797 B.n4 80.7344
R1222 B.n797 B.n796 80.7344
R1223 B.n796 B.n795 80.7344
R1224 B.n795 B.n8 80.7344
R1225 B.n12 B.n8 80.7344
R1226 B.n788 B.n12 80.7344
R1227 B.n788 B.n787 80.7344
R1228 B.n787 B.n786 80.7344
R1229 B.n786 B.t1 80.7344
R1230 B.n780 B.t1 80.7344
R1231 B.n780 B.n779 80.7344
R1232 B.n779 B.n778 80.7344
R1233 B.n778 B.n22 80.7344
R1234 B.n772 B.n22 80.7344
R1235 B.n772 B.n771 80.7344
R1236 B.n771 B.n770 80.7344
R1237 B.n770 B.n29 80.7344
R1238 B.n764 B.n29 80.7344
R1239 B.n764 B.n763 80.7344
R1240 B.n763 B.n762 80.7344
R1241 B.n756 B.n39 80.7344
R1242 B.n756 B.n755 80.7344
R1243 B.n755 B.n754 80.7344
R1244 B.n754 B.n43 80.7344
R1245 B.n748 B.n43 80.7344
R1246 B.n748 B.n747 80.7344
R1247 B.n747 B.n746 80.7344
R1248 B.n746 B.n50 80.7344
R1249 B.n740 B.n50 80.7344
R1250 B.n740 B.n739 80.7344
R1251 B.n739 B.n738 80.7344
R1252 B.n732 B.n60 80.7344
R1253 B.n732 B.n731 80.7344
R1254 B.n731 B.n730 80.7344
R1255 B.n730 B.n64 80.7344
R1256 B.n724 B.n64 80.7344
R1257 B.n724 B.n723 80.7344
R1258 B.n723 B.n722 80.7344
R1259 B.n722 B.n71 80.7344
R1260 B.n716 B.n71 80.7344
R1261 B.n716 B.n715 80.7344
R1262 B.n715 B.n714 80.7344
R1263 B.n714 B.n78 80.7344
R1264 B.n708 B.n78 80.7344
R1265 B.n708 B.n707 80.7344
R1266 B.n706 B.n85 80.7344
R1267 B.n700 B.n85 80.7344
R1268 B.n700 B.n699 80.7344
R1269 B.n699 B.n698 80.7344
R1270 B.n698 B.n92 80.7344
R1271 B.n692 B.n92 80.7344
R1272 B.n692 B.n691 80.7344
R1273 B.n691 B.n690 80.7344
R1274 B.n690 B.n99 80.7344
R1275 B.n130 B.n129 77.7702
R1276 B.n127 B.n126 77.7702
R1277 B.n350 B.n349 77.7702
R1278 B.n348 B.n347 77.7702
R1279 B.n685 B.n684 71.676
R1280 B.n132 B.n103 71.676
R1281 B.n136 B.n104 71.676
R1282 B.n140 B.n105 71.676
R1283 B.n144 B.n106 71.676
R1284 B.n148 B.n107 71.676
R1285 B.n152 B.n108 71.676
R1286 B.n156 B.n109 71.676
R1287 B.n160 B.n110 71.676
R1288 B.n164 B.n111 71.676
R1289 B.n168 B.n112 71.676
R1290 B.n172 B.n113 71.676
R1291 B.n176 B.n114 71.676
R1292 B.n180 B.n115 71.676
R1293 B.n184 B.n116 71.676
R1294 B.n188 B.n117 71.676
R1295 B.n192 B.n118 71.676
R1296 B.n196 B.n119 71.676
R1297 B.n200 B.n120 71.676
R1298 B.n204 B.n121 71.676
R1299 B.n208 B.n122 71.676
R1300 B.n212 B.n123 71.676
R1301 B.n682 B.n124 71.676
R1302 B.n682 B.n681 71.676
R1303 B.n214 B.n123 71.676
R1304 B.n211 B.n122 71.676
R1305 B.n207 B.n121 71.676
R1306 B.n203 B.n120 71.676
R1307 B.n199 B.n119 71.676
R1308 B.n195 B.n118 71.676
R1309 B.n191 B.n117 71.676
R1310 B.n187 B.n116 71.676
R1311 B.n183 B.n115 71.676
R1312 B.n179 B.n114 71.676
R1313 B.n175 B.n113 71.676
R1314 B.n171 B.n112 71.676
R1315 B.n167 B.n111 71.676
R1316 B.n163 B.n110 71.676
R1317 B.n159 B.n109 71.676
R1318 B.n155 B.n108 71.676
R1319 B.n151 B.n107 71.676
R1320 B.n147 B.n106 71.676
R1321 B.n143 B.n105 71.676
R1322 B.n139 B.n104 71.676
R1323 B.n135 B.n103 71.676
R1324 B.n684 B.n102 71.676
R1325 B.n441 B.n440 71.676
R1326 B.n346 B.n324 71.676
R1327 B.n433 B.n325 71.676
R1328 B.n429 B.n326 71.676
R1329 B.n425 B.n327 71.676
R1330 B.n421 B.n328 71.676
R1331 B.n417 B.n329 71.676
R1332 B.n413 B.n330 71.676
R1333 B.n409 B.n331 71.676
R1334 B.n404 B.n332 71.676
R1335 B.n400 B.n333 71.676
R1336 B.n396 B.n334 71.676
R1337 B.n392 B.n335 71.676
R1338 B.n388 B.n336 71.676
R1339 B.n383 B.n337 71.676
R1340 B.n379 B.n338 71.676
R1341 B.n375 B.n339 71.676
R1342 B.n371 B.n340 71.676
R1343 B.n367 B.n341 71.676
R1344 B.n363 B.n342 71.676
R1345 B.n359 B.n343 71.676
R1346 B.n355 B.n344 71.676
R1347 B.n440 B.n323 71.676
R1348 B.n434 B.n324 71.676
R1349 B.n430 B.n325 71.676
R1350 B.n426 B.n326 71.676
R1351 B.n422 B.n327 71.676
R1352 B.n418 B.n328 71.676
R1353 B.n414 B.n329 71.676
R1354 B.n410 B.n330 71.676
R1355 B.n405 B.n331 71.676
R1356 B.n401 B.n332 71.676
R1357 B.n397 B.n333 71.676
R1358 B.n393 B.n334 71.676
R1359 B.n389 B.n335 71.676
R1360 B.n384 B.n336 71.676
R1361 B.n380 B.n337 71.676
R1362 B.n376 B.n338 71.676
R1363 B.n372 B.n339 71.676
R1364 B.n368 B.n340 71.676
R1365 B.n364 B.n341 71.676
R1366 B.n360 B.n342 71.676
R1367 B.n356 B.n343 71.676
R1368 B.n352 B.n344 71.676
R1369 B.n799 B.n798 71.676
R1370 B.n799 B.n2 71.676
R1371 B.n556 B.t0 64.1128
R1372 B.n762 B.t2 64.1128
R1373 B.n131 B.n130 59.5399
R1374 B.n128 B.n127 59.5399
R1375 B.n386 B.n350 59.5399
R1376 B.n407 B.n348 59.5399
R1377 B.t11 B.n300 47.4911
R1378 B.n519 B.t4 47.4911
R1379 B.n738 B.t3 47.4911
R1380 B.n707 B.t7 47.4911
R1381 B.n470 B.t11 33.2439
R1382 B.n512 B.t4 33.2439
R1383 B.n60 B.t3 33.2439
R1384 B.t7 B.n706 33.2439
R1385 B.n443 B.n442 28.5664
R1386 B.n351 B.n318 28.5664
R1387 B.n687 B.n686 28.5664
R1388 B.n680 B.n679 28.5664
R1389 B B.n800 18.0485
R1390 B.n549 B.t0 16.6222
R1391 B.n39 B.t2 16.6222
R1392 B.n444 B.n443 10.6151
R1393 B.n444 B.n314 10.6151
R1394 B.n454 B.n314 10.6151
R1395 B.n455 B.n454 10.6151
R1396 B.n456 B.n455 10.6151
R1397 B.n456 B.n306 10.6151
R1398 B.n466 B.n306 10.6151
R1399 B.n467 B.n466 10.6151
R1400 B.n468 B.n467 10.6151
R1401 B.n468 B.n298 10.6151
R1402 B.n478 B.n298 10.6151
R1403 B.n479 B.n478 10.6151
R1404 B.n480 B.n479 10.6151
R1405 B.n480 B.n290 10.6151
R1406 B.n490 B.n290 10.6151
R1407 B.n491 B.n490 10.6151
R1408 B.n492 B.n491 10.6151
R1409 B.n492 B.n282 10.6151
R1410 B.n502 B.n282 10.6151
R1411 B.n503 B.n502 10.6151
R1412 B.n504 B.n503 10.6151
R1413 B.n504 B.n274 10.6151
R1414 B.n515 B.n274 10.6151
R1415 B.n516 B.n515 10.6151
R1416 B.n517 B.n516 10.6151
R1417 B.n517 B.n267 10.6151
R1418 B.n527 B.n267 10.6151
R1419 B.n528 B.n527 10.6151
R1420 B.n529 B.n528 10.6151
R1421 B.n529 B.n259 10.6151
R1422 B.n539 B.n259 10.6151
R1423 B.n540 B.n539 10.6151
R1424 B.n541 B.n540 10.6151
R1425 B.n541 B.n251 10.6151
R1426 B.n552 B.n251 10.6151
R1427 B.n553 B.n552 10.6151
R1428 B.n554 B.n553 10.6151
R1429 B.n554 B.n244 10.6151
R1430 B.n564 B.n244 10.6151
R1431 B.n565 B.n564 10.6151
R1432 B.n566 B.n565 10.6151
R1433 B.n566 B.n236 10.6151
R1434 B.n576 B.n236 10.6151
R1435 B.n577 B.n576 10.6151
R1436 B.n578 B.n577 10.6151
R1437 B.n578 B.n228 10.6151
R1438 B.n588 B.n228 10.6151
R1439 B.n589 B.n588 10.6151
R1440 B.n590 B.n589 10.6151
R1441 B.n590 B.n221 10.6151
R1442 B.n601 B.n221 10.6151
R1443 B.n602 B.n601 10.6151
R1444 B.n603 B.n602 10.6151
R1445 B.n603 B.n0 10.6151
R1446 B.n442 B.n322 10.6151
R1447 B.n437 B.n322 10.6151
R1448 B.n437 B.n436 10.6151
R1449 B.n436 B.n435 10.6151
R1450 B.n435 B.n432 10.6151
R1451 B.n432 B.n431 10.6151
R1452 B.n431 B.n428 10.6151
R1453 B.n428 B.n427 10.6151
R1454 B.n427 B.n424 10.6151
R1455 B.n424 B.n423 10.6151
R1456 B.n423 B.n420 10.6151
R1457 B.n420 B.n419 10.6151
R1458 B.n419 B.n416 10.6151
R1459 B.n416 B.n415 10.6151
R1460 B.n415 B.n412 10.6151
R1461 B.n412 B.n411 10.6151
R1462 B.n411 B.n408 10.6151
R1463 B.n406 B.n403 10.6151
R1464 B.n403 B.n402 10.6151
R1465 B.n402 B.n399 10.6151
R1466 B.n399 B.n398 10.6151
R1467 B.n398 B.n395 10.6151
R1468 B.n395 B.n394 10.6151
R1469 B.n394 B.n391 10.6151
R1470 B.n391 B.n390 10.6151
R1471 B.n390 B.n387 10.6151
R1472 B.n385 B.n382 10.6151
R1473 B.n382 B.n381 10.6151
R1474 B.n381 B.n378 10.6151
R1475 B.n378 B.n377 10.6151
R1476 B.n377 B.n374 10.6151
R1477 B.n374 B.n373 10.6151
R1478 B.n373 B.n370 10.6151
R1479 B.n370 B.n369 10.6151
R1480 B.n369 B.n366 10.6151
R1481 B.n366 B.n365 10.6151
R1482 B.n365 B.n362 10.6151
R1483 B.n362 B.n361 10.6151
R1484 B.n361 B.n358 10.6151
R1485 B.n358 B.n357 10.6151
R1486 B.n357 B.n354 10.6151
R1487 B.n354 B.n353 10.6151
R1488 B.n353 B.n351 10.6151
R1489 B.n448 B.n318 10.6151
R1490 B.n449 B.n448 10.6151
R1491 B.n450 B.n449 10.6151
R1492 B.n450 B.n310 10.6151
R1493 B.n460 B.n310 10.6151
R1494 B.n461 B.n460 10.6151
R1495 B.n462 B.n461 10.6151
R1496 B.n462 B.n302 10.6151
R1497 B.n472 B.n302 10.6151
R1498 B.n473 B.n472 10.6151
R1499 B.n474 B.n473 10.6151
R1500 B.n474 B.n294 10.6151
R1501 B.n484 B.n294 10.6151
R1502 B.n485 B.n484 10.6151
R1503 B.n486 B.n485 10.6151
R1504 B.n486 B.n286 10.6151
R1505 B.n496 B.n286 10.6151
R1506 B.n497 B.n496 10.6151
R1507 B.n498 B.n497 10.6151
R1508 B.n498 B.n278 10.6151
R1509 B.n508 B.n278 10.6151
R1510 B.n509 B.n508 10.6151
R1511 B.n510 B.n509 10.6151
R1512 B.n510 B.n271 10.6151
R1513 B.n521 B.n271 10.6151
R1514 B.n522 B.n521 10.6151
R1515 B.n523 B.n522 10.6151
R1516 B.n523 B.n263 10.6151
R1517 B.n533 B.n263 10.6151
R1518 B.n534 B.n533 10.6151
R1519 B.n535 B.n534 10.6151
R1520 B.n535 B.n255 10.6151
R1521 B.n545 B.n255 10.6151
R1522 B.n546 B.n545 10.6151
R1523 B.n547 B.n546 10.6151
R1524 B.n547 B.n248 10.6151
R1525 B.n558 B.n248 10.6151
R1526 B.n559 B.n558 10.6151
R1527 B.n560 B.n559 10.6151
R1528 B.n560 B.n240 10.6151
R1529 B.n570 B.n240 10.6151
R1530 B.n571 B.n570 10.6151
R1531 B.n572 B.n571 10.6151
R1532 B.n572 B.n232 10.6151
R1533 B.n582 B.n232 10.6151
R1534 B.n583 B.n582 10.6151
R1535 B.n584 B.n583 10.6151
R1536 B.n584 B.n225 10.6151
R1537 B.n594 B.n225 10.6151
R1538 B.n595 B.n594 10.6151
R1539 B.n597 B.n595 10.6151
R1540 B.n597 B.n596 10.6151
R1541 B.n596 B.n217 10.6151
R1542 B.n608 B.n217 10.6151
R1543 B.n609 B.n608 10.6151
R1544 B.n610 B.n609 10.6151
R1545 B.n611 B.n610 10.6151
R1546 B.n612 B.n611 10.6151
R1547 B.n615 B.n612 10.6151
R1548 B.n616 B.n615 10.6151
R1549 B.n617 B.n616 10.6151
R1550 B.n618 B.n617 10.6151
R1551 B.n620 B.n618 10.6151
R1552 B.n621 B.n620 10.6151
R1553 B.n622 B.n621 10.6151
R1554 B.n623 B.n622 10.6151
R1555 B.n625 B.n623 10.6151
R1556 B.n626 B.n625 10.6151
R1557 B.n627 B.n626 10.6151
R1558 B.n628 B.n627 10.6151
R1559 B.n630 B.n628 10.6151
R1560 B.n631 B.n630 10.6151
R1561 B.n632 B.n631 10.6151
R1562 B.n633 B.n632 10.6151
R1563 B.n635 B.n633 10.6151
R1564 B.n636 B.n635 10.6151
R1565 B.n637 B.n636 10.6151
R1566 B.n638 B.n637 10.6151
R1567 B.n640 B.n638 10.6151
R1568 B.n641 B.n640 10.6151
R1569 B.n642 B.n641 10.6151
R1570 B.n643 B.n642 10.6151
R1571 B.n645 B.n643 10.6151
R1572 B.n646 B.n645 10.6151
R1573 B.n647 B.n646 10.6151
R1574 B.n648 B.n647 10.6151
R1575 B.n650 B.n648 10.6151
R1576 B.n651 B.n650 10.6151
R1577 B.n652 B.n651 10.6151
R1578 B.n653 B.n652 10.6151
R1579 B.n655 B.n653 10.6151
R1580 B.n656 B.n655 10.6151
R1581 B.n657 B.n656 10.6151
R1582 B.n658 B.n657 10.6151
R1583 B.n660 B.n658 10.6151
R1584 B.n661 B.n660 10.6151
R1585 B.n662 B.n661 10.6151
R1586 B.n663 B.n662 10.6151
R1587 B.n665 B.n663 10.6151
R1588 B.n666 B.n665 10.6151
R1589 B.n667 B.n666 10.6151
R1590 B.n668 B.n667 10.6151
R1591 B.n670 B.n668 10.6151
R1592 B.n671 B.n670 10.6151
R1593 B.n672 B.n671 10.6151
R1594 B.n673 B.n672 10.6151
R1595 B.n675 B.n673 10.6151
R1596 B.n676 B.n675 10.6151
R1597 B.n677 B.n676 10.6151
R1598 B.n678 B.n677 10.6151
R1599 B.n679 B.n678 10.6151
R1600 B.n792 B.n1 10.6151
R1601 B.n792 B.n791 10.6151
R1602 B.n791 B.n790 10.6151
R1603 B.n790 B.n10 10.6151
R1604 B.n784 B.n10 10.6151
R1605 B.n784 B.n783 10.6151
R1606 B.n783 B.n782 10.6151
R1607 B.n782 B.n17 10.6151
R1608 B.n776 B.n17 10.6151
R1609 B.n776 B.n775 10.6151
R1610 B.n775 B.n774 10.6151
R1611 B.n774 B.n24 10.6151
R1612 B.n768 B.n24 10.6151
R1613 B.n768 B.n767 10.6151
R1614 B.n767 B.n766 10.6151
R1615 B.n766 B.n31 10.6151
R1616 B.n760 B.n31 10.6151
R1617 B.n760 B.n759 10.6151
R1618 B.n759 B.n758 10.6151
R1619 B.n758 B.n37 10.6151
R1620 B.n752 B.n37 10.6151
R1621 B.n752 B.n751 10.6151
R1622 B.n751 B.n750 10.6151
R1623 B.n750 B.n45 10.6151
R1624 B.n744 B.n45 10.6151
R1625 B.n744 B.n743 10.6151
R1626 B.n743 B.n742 10.6151
R1627 B.n742 B.n52 10.6151
R1628 B.n736 B.n52 10.6151
R1629 B.n736 B.n735 10.6151
R1630 B.n735 B.n734 10.6151
R1631 B.n734 B.n58 10.6151
R1632 B.n728 B.n58 10.6151
R1633 B.n728 B.n727 10.6151
R1634 B.n727 B.n726 10.6151
R1635 B.n726 B.n66 10.6151
R1636 B.n720 B.n66 10.6151
R1637 B.n720 B.n719 10.6151
R1638 B.n719 B.n718 10.6151
R1639 B.n718 B.n73 10.6151
R1640 B.n712 B.n73 10.6151
R1641 B.n712 B.n711 10.6151
R1642 B.n711 B.n710 10.6151
R1643 B.n710 B.n80 10.6151
R1644 B.n704 B.n80 10.6151
R1645 B.n704 B.n703 10.6151
R1646 B.n703 B.n702 10.6151
R1647 B.n702 B.n87 10.6151
R1648 B.n696 B.n87 10.6151
R1649 B.n696 B.n695 10.6151
R1650 B.n695 B.n694 10.6151
R1651 B.n694 B.n94 10.6151
R1652 B.n688 B.n94 10.6151
R1653 B.n688 B.n687 10.6151
R1654 B.n686 B.n101 10.6151
R1655 B.n133 B.n101 10.6151
R1656 B.n134 B.n133 10.6151
R1657 B.n137 B.n134 10.6151
R1658 B.n138 B.n137 10.6151
R1659 B.n141 B.n138 10.6151
R1660 B.n142 B.n141 10.6151
R1661 B.n145 B.n142 10.6151
R1662 B.n146 B.n145 10.6151
R1663 B.n149 B.n146 10.6151
R1664 B.n150 B.n149 10.6151
R1665 B.n153 B.n150 10.6151
R1666 B.n154 B.n153 10.6151
R1667 B.n157 B.n154 10.6151
R1668 B.n158 B.n157 10.6151
R1669 B.n161 B.n158 10.6151
R1670 B.n162 B.n161 10.6151
R1671 B.n166 B.n165 10.6151
R1672 B.n169 B.n166 10.6151
R1673 B.n170 B.n169 10.6151
R1674 B.n173 B.n170 10.6151
R1675 B.n174 B.n173 10.6151
R1676 B.n177 B.n174 10.6151
R1677 B.n178 B.n177 10.6151
R1678 B.n181 B.n178 10.6151
R1679 B.n182 B.n181 10.6151
R1680 B.n186 B.n185 10.6151
R1681 B.n189 B.n186 10.6151
R1682 B.n190 B.n189 10.6151
R1683 B.n193 B.n190 10.6151
R1684 B.n194 B.n193 10.6151
R1685 B.n197 B.n194 10.6151
R1686 B.n198 B.n197 10.6151
R1687 B.n201 B.n198 10.6151
R1688 B.n202 B.n201 10.6151
R1689 B.n205 B.n202 10.6151
R1690 B.n206 B.n205 10.6151
R1691 B.n209 B.n206 10.6151
R1692 B.n210 B.n209 10.6151
R1693 B.n213 B.n210 10.6151
R1694 B.n215 B.n213 10.6151
R1695 B.n216 B.n215 10.6151
R1696 B.n680 B.n216 10.6151
R1697 B.n408 B.n407 9.36635
R1698 B.n386 B.n385 9.36635
R1699 B.n162 B.n131 9.36635
R1700 B.n185 B.n128 9.36635
R1701 B.n800 B.n0 8.11757
R1702 B.n800 B.n1 8.11757
R1703 B.n407 B.n406 1.24928
R1704 B.n387 B.n386 1.24928
R1705 B.n165 B.n131 1.24928
R1706 B.n182 B.n128 1.24928
R1707 VN.n38 VN.n37 161.3
R1708 VN.n36 VN.n21 161.3
R1709 VN.n35 VN.n34 161.3
R1710 VN.n33 VN.n22 161.3
R1711 VN.n32 VN.n31 161.3
R1712 VN.n30 VN.n23 161.3
R1713 VN.n29 VN.n28 161.3
R1714 VN.n27 VN.n24 161.3
R1715 VN.n18 VN.n17 161.3
R1716 VN.n16 VN.n1 161.3
R1717 VN.n15 VN.n14 161.3
R1718 VN.n13 VN.n2 161.3
R1719 VN.n12 VN.n11 161.3
R1720 VN.n10 VN.n3 161.3
R1721 VN.n9 VN.n8 161.3
R1722 VN.n7 VN.n4 161.3
R1723 VN.n19 VN.n0 89.5781
R1724 VN.n39 VN.n20 89.5781
R1725 VN.n26 VN.t3 58.3844
R1726 VN.n6 VN.t1 58.3844
R1727 VN.n26 VN.n25 50.4792
R1728 VN.n6 VN.n5 50.4792
R1729 VN VN.n39 46.9942
R1730 VN.n11 VN.n2 40.979
R1731 VN.n31 VN.n22 40.979
R1732 VN.n11 VN.n10 40.0078
R1733 VN.n31 VN.n30 40.0078
R1734 VN.n5 VN.t5 26.1307
R1735 VN.n0 VN.t0 26.1307
R1736 VN.n25 VN.t2 26.1307
R1737 VN.n20 VN.t4 26.1307
R1738 VN.n5 VN.n4 24.4675
R1739 VN.n9 VN.n4 24.4675
R1740 VN.n10 VN.n9 24.4675
R1741 VN.n15 VN.n2 24.4675
R1742 VN.n16 VN.n15 24.4675
R1743 VN.n17 VN.n16 24.4675
R1744 VN.n30 VN.n29 24.4675
R1745 VN.n29 VN.n24 24.4675
R1746 VN.n25 VN.n24 24.4675
R1747 VN.n37 VN.n36 24.4675
R1748 VN.n36 VN.n35 24.4675
R1749 VN.n35 VN.n22 24.4675
R1750 VN.n27 VN.n26 2.51578
R1751 VN.n7 VN.n6 2.51578
R1752 VN.n17 VN.n0 0.48984
R1753 VN.n37 VN.n20 0.48984
R1754 VN.n39 VN.n38 0.354971
R1755 VN.n19 VN.n18 0.354971
R1756 VN VN.n19 0.26696
R1757 VN.n38 VN.n21 0.189894
R1758 VN.n34 VN.n21 0.189894
R1759 VN.n34 VN.n33 0.189894
R1760 VN.n33 VN.n32 0.189894
R1761 VN.n32 VN.n23 0.189894
R1762 VN.n28 VN.n23 0.189894
R1763 VN.n28 VN.n27 0.189894
R1764 VN.n8 VN.n7 0.189894
R1765 VN.n8 VN.n3 0.189894
R1766 VN.n12 VN.n3 0.189894
R1767 VN.n13 VN.n12 0.189894
R1768 VN.n14 VN.n13 0.189894
R1769 VN.n14 VN.n1 0.189894
R1770 VN.n18 VN.n1 0.189894
R1771 VDD2.n35 VDD2.n21 289.615
R1772 VDD2.n14 VDD2.n0 289.615
R1773 VDD2.n36 VDD2.n35 185
R1774 VDD2.n34 VDD2.n33 185
R1775 VDD2.n25 VDD2.n24 185
R1776 VDD2.n28 VDD2.n27 185
R1777 VDD2.n7 VDD2.n6 185
R1778 VDD2.n4 VDD2.n3 185
R1779 VDD2.n13 VDD2.n12 185
R1780 VDD2.n15 VDD2.n14 185
R1781 VDD2.t1 VDD2.n26 147.888
R1782 VDD2.t4 VDD2.n5 147.888
R1783 VDD2.n35 VDD2.n34 104.615
R1784 VDD2.n34 VDD2.n24 104.615
R1785 VDD2.n27 VDD2.n24 104.615
R1786 VDD2.n6 VDD2.n3 104.615
R1787 VDD2.n13 VDD2.n3 104.615
R1788 VDD2.n14 VDD2.n13 104.615
R1789 VDD2.n20 VDD2.n19 77.1819
R1790 VDD2 VDD2.n41 77.1791
R1791 VDD2.n20 VDD2.n18 54.3106
R1792 VDD2.n27 VDD2.t1 52.3082
R1793 VDD2.n6 VDD2.t4 52.3082
R1794 VDD2.n40 VDD2.n39 51.7732
R1795 VDD2.n40 VDD2.n20 38.3899
R1796 VDD2.n28 VDD2.n26 15.6496
R1797 VDD2.n7 VDD2.n5 15.6496
R1798 VDD2.n29 VDD2.n25 12.8005
R1799 VDD2.n8 VDD2.n4 12.8005
R1800 VDD2.n33 VDD2.n32 12.0247
R1801 VDD2.n12 VDD2.n11 12.0247
R1802 VDD2.n36 VDD2.n23 11.249
R1803 VDD2.n15 VDD2.n2 11.249
R1804 VDD2.n37 VDD2.n21 10.4732
R1805 VDD2.n16 VDD2.n0 10.4732
R1806 VDD2.n39 VDD2.n38 9.45567
R1807 VDD2.n18 VDD2.n17 9.45567
R1808 VDD2.n38 VDD2.n37 9.3005
R1809 VDD2.n23 VDD2.n22 9.3005
R1810 VDD2.n32 VDD2.n31 9.3005
R1811 VDD2.n30 VDD2.n29 9.3005
R1812 VDD2.n17 VDD2.n16 9.3005
R1813 VDD2.n2 VDD2.n1 9.3005
R1814 VDD2.n11 VDD2.n10 9.3005
R1815 VDD2.n9 VDD2.n8 9.3005
R1816 VDD2.n41 VDD2.t3 4.96291
R1817 VDD2.n41 VDD2.t2 4.96291
R1818 VDD2.n19 VDD2.t0 4.96291
R1819 VDD2.n19 VDD2.t5 4.96291
R1820 VDD2.n30 VDD2.n26 4.40546
R1821 VDD2.n9 VDD2.n5 4.40546
R1822 VDD2.n39 VDD2.n21 3.49141
R1823 VDD2.n18 VDD2.n0 3.49141
R1824 VDD2.n37 VDD2.n36 2.71565
R1825 VDD2.n16 VDD2.n15 2.71565
R1826 VDD2 VDD2.n40 2.65136
R1827 VDD2.n33 VDD2.n23 1.93989
R1828 VDD2.n12 VDD2.n2 1.93989
R1829 VDD2.n32 VDD2.n25 1.16414
R1830 VDD2.n11 VDD2.n4 1.16414
R1831 VDD2.n29 VDD2.n28 0.388379
R1832 VDD2.n8 VDD2.n7 0.388379
R1833 VDD2.n38 VDD2.n22 0.155672
R1834 VDD2.n31 VDD2.n22 0.155672
R1835 VDD2.n31 VDD2.n30 0.155672
R1836 VDD2.n10 VDD2.n9 0.155672
R1837 VDD2.n10 VDD2.n1 0.155672
R1838 VDD2.n17 VDD2.n1 0.155672
C0 VTAIL VP 3.69133f
C1 VTAIL VN 3.6771f
C2 VDD1 VTAIL 5.52924f
C3 VDD2 VP 0.554053f
C4 VDD2 VN 2.64293f
C5 VN VP 6.50306f
C6 VDD1 VDD2 1.8264f
C7 VDD1 VP 3.038f
C8 VDD1 VN 0.156308f
C9 VDD2 VTAIL 5.58949f
C10 VDD2 B 5.382374f
C11 VDD1 B 5.569437f
C12 VTAIL B 4.787744f
C13 VN B 15.3645f
C14 VP B 13.994438f
C15 VDD2.n0 B 0.031576f
C16 VDD2.n1 B 0.022146f
C17 VDD2.n2 B 0.0119f
C18 VDD2.n3 B 0.028127f
C19 VDD2.n4 B 0.0126f
C20 VDD2.n5 B 0.085583f
C21 VDD2.t4 B 0.046804f
C22 VDD2.n6 B 0.021096f
C23 VDD2.n7 B 0.016555f
C24 VDD2.n8 B 0.0119f
C25 VDD2.n9 B 0.319902f
C26 VDD2.n10 B 0.022146f
C27 VDD2.n11 B 0.0119f
C28 VDD2.n12 B 0.0126f
C29 VDD2.n13 B 0.028127f
C30 VDD2.n14 B 0.061684f
C31 VDD2.n15 B 0.0126f
C32 VDD2.n16 B 0.0119f
C33 VDD2.n17 B 0.055727f
C34 VDD2.n18 B 0.060571f
C35 VDD2.t0 B 0.069826f
C36 VDD2.t5 B 0.069826f
C37 VDD2.n19 B 0.553155f
C38 VDD2.n20 B 2.3481f
C39 VDD2.n21 B 0.031576f
C40 VDD2.n22 B 0.022146f
C41 VDD2.n23 B 0.0119f
C42 VDD2.n24 B 0.028127f
C43 VDD2.n25 B 0.0126f
C44 VDD2.n26 B 0.085583f
C45 VDD2.t1 B 0.046804f
C46 VDD2.n27 B 0.021096f
C47 VDD2.n28 B 0.016555f
C48 VDD2.n29 B 0.0119f
C49 VDD2.n30 B 0.319902f
C50 VDD2.n31 B 0.022146f
C51 VDD2.n32 B 0.0119f
C52 VDD2.n33 B 0.0126f
C53 VDD2.n34 B 0.028127f
C54 VDD2.n35 B 0.061684f
C55 VDD2.n36 B 0.0126f
C56 VDD2.n37 B 0.0119f
C57 VDD2.n38 B 0.055727f
C58 VDD2.n39 B 0.049989f
C59 VDD2.n40 B 1.97859f
C60 VDD2.t3 B 0.069826f
C61 VDD2.t2 B 0.069826f
C62 VDD2.n41 B 0.553129f
C63 VN.t0 B 0.900706f
C64 VN.n0 B 0.433662f
C65 VN.n1 B 0.023884f
C66 VN.n2 B 0.047348f
C67 VN.n3 B 0.023884f
C68 VN.n4 B 0.044514f
C69 VN.t5 B 0.900706f
C70 VN.n5 B 0.44714f
C71 VN.t1 B 1.19715f
C72 VN.n6 B 0.444248f
C73 VN.n7 B 0.304484f
C74 VN.n8 B 0.023884f
C75 VN.n9 B 0.044514f
C76 VN.n10 B 0.047587f
C77 VN.n11 B 0.019317f
C78 VN.n12 B 0.023884f
C79 VN.n13 B 0.023884f
C80 VN.n14 B 0.023884f
C81 VN.n15 B 0.044514f
C82 VN.n16 B 0.044514f
C83 VN.n17 B 0.022977f
C84 VN.n18 B 0.038548f
C85 VN.n19 B 0.073315f
C86 VN.t4 B 0.900706f
C87 VN.n20 B 0.433662f
C88 VN.n21 B 0.023884f
C89 VN.n22 B 0.047348f
C90 VN.n23 B 0.023884f
C91 VN.n24 B 0.044514f
C92 VN.t3 B 1.19715f
C93 VN.t2 B 0.900706f
C94 VN.n25 B 0.44714f
C95 VN.n26 B 0.444248f
C96 VN.n27 B 0.304484f
C97 VN.n28 B 0.023884f
C98 VN.n29 B 0.044514f
C99 VN.n30 B 0.047587f
C100 VN.n31 B 0.019317f
C101 VN.n32 B 0.023884f
C102 VN.n33 B 0.023884f
C103 VN.n34 B 0.023884f
C104 VN.n35 B 0.044514f
C105 VN.n36 B 0.044514f
C106 VN.n37 B 0.022977f
C107 VN.n38 B 0.038548f
C108 VN.n39 B 1.25882f
C109 VDD1.n0 B 0.032408f
C110 VDD1.n1 B 0.022729f
C111 VDD1.n2 B 0.012214f
C112 VDD1.n3 B 0.028869f
C113 VDD1.n4 B 0.012932f
C114 VDD1.n5 B 0.087838f
C115 VDD1.t1 B 0.048037f
C116 VDD1.n6 B 0.021651f
C117 VDD1.n7 B 0.016991f
C118 VDD1.n8 B 0.012214f
C119 VDD1.n9 B 0.328331f
C120 VDD1.n10 B 0.022729f
C121 VDD1.n11 B 0.012214f
C122 VDD1.n12 B 0.012932f
C123 VDD1.n13 B 0.028869f
C124 VDD1.n14 B 0.063309f
C125 VDD1.n15 B 0.012932f
C126 VDD1.n16 B 0.012214f
C127 VDD1.n17 B 0.057195f
C128 VDD1.n18 B 0.063024f
C129 VDD1.n19 B 0.032408f
C130 VDD1.n20 B 0.022729f
C131 VDD1.n21 B 0.012214f
C132 VDD1.n22 B 0.028869f
C133 VDD1.n23 B 0.012932f
C134 VDD1.n24 B 0.087838f
C135 VDD1.t4 B 0.048037f
C136 VDD1.n25 B 0.021651f
C137 VDD1.n26 B 0.016991f
C138 VDD1.n27 B 0.012214f
C139 VDD1.n28 B 0.328331f
C140 VDD1.n29 B 0.022729f
C141 VDD1.n30 B 0.012214f
C142 VDD1.n31 B 0.012932f
C143 VDD1.n32 B 0.028869f
C144 VDD1.n33 B 0.063309f
C145 VDD1.n34 B 0.012932f
C146 VDD1.n35 B 0.012214f
C147 VDD1.n36 B 0.057195f
C148 VDD1.n37 B 0.062167f
C149 VDD1.t0 B 0.071665f
C150 VDD1.t5 B 0.071665f
C151 VDD1.n38 B 0.567729f
C152 VDD1.n39 B 2.54051f
C153 VDD1.t2 B 0.071665f
C154 VDD1.t3 B 0.071665f
C155 VDD1.n40 B 0.562495f
C156 VDD1.n41 B 2.24216f
C157 VTAIL.t11 B 0.098522f
C158 VTAIL.t7 B 0.098522f
C159 VTAIL.n0 B 0.706868f
C160 VTAIL.n1 B 0.581822f
C161 VTAIL.n2 B 0.044553f
C162 VTAIL.n3 B 0.031247f
C163 VTAIL.n4 B 0.016791f
C164 VTAIL.n5 B 0.039687f
C165 VTAIL.n6 B 0.017778f
C166 VTAIL.n7 B 0.120755f
C167 VTAIL.t5 B 0.066039f
C168 VTAIL.n8 B 0.029765f
C169 VTAIL.n9 B 0.023358f
C170 VTAIL.n10 B 0.016791f
C171 VTAIL.n11 B 0.451372f
C172 VTAIL.n12 B 0.031247f
C173 VTAIL.n13 B 0.016791f
C174 VTAIL.n14 B 0.017778f
C175 VTAIL.n15 B 0.039687f
C176 VTAIL.n16 B 0.087034f
C177 VTAIL.n17 B 0.017778f
C178 VTAIL.n18 B 0.016791f
C179 VTAIL.n19 B 0.078628f
C180 VTAIL.n20 B 0.049003f
C181 VTAIL.n21 B 0.599694f
C182 VTAIL.t3 B 0.098522f
C183 VTAIL.t4 B 0.098522f
C184 VTAIL.n22 B 0.706868f
C185 VTAIL.n23 B 2.08255f
C186 VTAIL.t6 B 0.098522f
C187 VTAIL.t10 B 0.098522f
C188 VTAIL.n24 B 0.706872f
C189 VTAIL.n25 B 2.08254f
C190 VTAIL.n26 B 0.044553f
C191 VTAIL.n27 B 0.031247f
C192 VTAIL.n28 B 0.016791f
C193 VTAIL.n29 B 0.039687f
C194 VTAIL.n30 B 0.017778f
C195 VTAIL.n31 B 0.120755f
C196 VTAIL.t8 B 0.066039f
C197 VTAIL.n32 B 0.029765f
C198 VTAIL.n33 B 0.023358f
C199 VTAIL.n34 B 0.016791f
C200 VTAIL.n35 B 0.451372f
C201 VTAIL.n36 B 0.031247f
C202 VTAIL.n37 B 0.016791f
C203 VTAIL.n38 B 0.017778f
C204 VTAIL.n39 B 0.039687f
C205 VTAIL.n40 B 0.087034f
C206 VTAIL.n41 B 0.017778f
C207 VTAIL.n42 B 0.016791f
C208 VTAIL.n43 B 0.078628f
C209 VTAIL.n44 B 0.049003f
C210 VTAIL.n45 B 0.599694f
C211 VTAIL.t1 B 0.098522f
C212 VTAIL.t0 B 0.098522f
C213 VTAIL.n46 B 0.706872f
C214 VTAIL.n47 B 0.836999f
C215 VTAIL.n48 B 0.044553f
C216 VTAIL.n49 B 0.031247f
C217 VTAIL.n50 B 0.016791f
C218 VTAIL.n51 B 0.039687f
C219 VTAIL.n52 B 0.017778f
C220 VTAIL.n53 B 0.120755f
C221 VTAIL.t2 B 0.066039f
C222 VTAIL.n54 B 0.029765f
C223 VTAIL.n55 B 0.023358f
C224 VTAIL.n56 B 0.016791f
C225 VTAIL.n57 B 0.451372f
C226 VTAIL.n58 B 0.031247f
C227 VTAIL.n59 B 0.016791f
C228 VTAIL.n60 B 0.017778f
C229 VTAIL.n61 B 0.039687f
C230 VTAIL.n62 B 0.087034f
C231 VTAIL.n63 B 0.017778f
C232 VTAIL.n64 B 0.016791f
C233 VTAIL.n65 B 0.078628f
C234 VTAIL.n66 B 0.049003f
C235 VTAIL.n67 B 1.49718f
C236 VTAIL.n68 B 0.044553f
C237 VTAIL.n69 B 0.031247f
C238 VTAIL.n70 B 0.016791f
C239 VTAIL.n71 B 0.039687f
C240 VTAIL.n72 B 0.017778f
C241 VTAIL.n73 B 0.120755f
C242 VTAIL.t9 B 0.066039f
C243 VTAIL.n74 B 0.029765f
C244 VTAIL.n75 B 0.023358f
C245 VTAIL.n76 B 0.016791f
C246 VTAIL.n77 B 0.451372f
C247 VTAIL.n78 B 0.031247f
C248 VTAIL.n79 B 0.016791f
C249 VTAIL.n80 B 0.017778f
C250 VTAIL.n81 B 0.039687f
C251 VTAIL.n82 B 0.087034f
C252 VTAIL.n83 B 0.017778f
C253 VTAIL.n84 B 0.016791f
C254 VTAIL.n85 B 0.078628f
C255 VTAIL.n86 B 0.049003f
C256 VTAIL.n87 B 1.40431f
C257 VP.t0 B 0.931296f
C258 VP.n0 B 0.44839f
C259 VP.n1 B 0.024695f
C260 VP.n2 B 0.048956f
C261 VP.n3 B 0.024695f
C262 VP.n4 B 0.046026f
C263 VP.n5 B 0.024695f
C264 VP.t5 B 0.931296f
C265 VP.n6 B 0.049203f
C266 VP.n7 B 0.024695f
C267 VP.n8 B 0.046026f
C268 VP.t2 B 0.931296f
C269 VP.n9 B 0.44839f
C270 VP.n10 B 0.024695f
C271 VP.n11 B 0.048956f
C272 VP.n12 B 0.024695f
C273 VP.n13 B 0.046026f
C274 VP.t4 B 1.2378f
C275 VP.t3 B 0.931296f
C276 VP.n14 B 0.462325f
C277 VP.n15 B 0.459337f
C278 VP.n16 B 0.314826f
C279 VP.n17 B 0.024695f
C280 VP.n18 B 0.046026f
C281 VP.n19 B 0.049203f
C282 VP.n20 B 0.019973f
C283 VP.n21 B 0.024695f
C284 VP.n22 B 0.024695f
C285 VP.n23 B 0.024695f
C286 VP.n24 B 0.046026f
C287 VP.n25 B 0.046026f
C288 VP.n26 B 0.023757f
C289 VP.n27 B 0.039858f
C290 VP.n28 B 1.29123f
C291 VP.n29 B 1.31018f
C292 VP.t1 B 0.931296f
C293 VP.n30 B 0.44839f
C294 VP.n31 B 0.023757f
C295 VP.n32 B 0.039858f
C296 VP.n33 B 0.024695f
C297 VP.n34 B 0.024695f
C298 VP.n35 B 0.046026f
C299 VP.n36 B 0.048956f
C300 VP.n37 B 0.019973f
C301 VP.n38 B 0.024695f
C302 VP.n39 B 0.024695f
C303 VP.n40 B 0.024695f
C304 VP.n41 B 0.046026f
C305 VP.n42 B 0.046026f
C306 VP.n43 B 0.384756f
C307 VP.n44 B 0.024695f
C308 VP.n45 B 0.024695f
C309 VP.n46 B 0.024695f
C310 VP.n47 B 0.046026f
C311 VP.n48 B 0.049203f
C312 VP.n49 B 0.019973f
C313 VP.n50 B 0.024695f
C314 VP.n51 B 0.024695f
C315 VP.n52 B 0.024695f
C316 VP.n53 B 0.046026f
C317 VP.n54 B 0.046026f
C318 VP.n55 B 0.023757f
C319 VP.n56 B 0.039858f
C320 VP.n57 B 0.075805f
.ends

