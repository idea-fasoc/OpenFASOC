* NGSPICE file created from diff_pair_sample_0316.ext - technology: sky130A

.subckt diff_pair_sample_0316 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t15 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=1.31175 pd=8.28 as=1.31175 ps=8.28 w=7.95 l=3.84
X1 VTAIL.t1 VN.t0 VDD2.t9 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=1.31175 pd=8.28 as=1.31175 ps=8.28 w=7.95 l=3.84
X2 VTAIL.t5 VN.t1 VDD2.t8 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=1.31175 pd=8.28 as=1.31175 ps=8.28 w=7.95 l=3.84
X3 VTAIL.t16 VP.t1 VDD1.t8 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=1.31175 pd=8.28 as=1.31175 ps=8.28 w=7.95 l=3.84
X4 VDD1.t7 VP.t2 VTAIL.t10 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=3.1005 pd=16.68 as=1.31175 ps=8.28 w=7.95 l=3.84
X5 VDD2.t7 VN.t2 VTAIL.t2 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=1.31175 pd=8.28 as=3.1005 ps=16.68 w=7.95 l=3.84
X6 VDD1.t6 VP.t3 VTAIL.t11 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=1.31175 pd=8.28 as=3.1005 ps=16.68 w=7.95 l=3.84
X7 VDD2.t6 VN.t3 VTAIL.t0 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=1.31175 pd=8.28 as=3.1005 ps=16.68 w=7.95 l=3.84
X8 VDD2.t5 VN.t4 VTAIL.t7 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=3.1005 pd=16.68 as=1.31175 ps=8.28 w=7.95 l=3.84
X9 VDD1.t5 VP.t4 VTAIL.t9 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=3.1005 pd=16.68 as=1.31175 ps=8.28 w=7.95 l=3.84
X10 B.t11 B.t9 B.t10 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=3.1005 pd=16.68 as=0 ps=0 w=7.95 l=3.84
X11 VDD2.t4 VN.t5 VTAIL.t4 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=3.1005 pd=16.68 as=1.31175 ps=8.28 w=7.95 l=3.84
X12 B.t8 B.t6 B.t7 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=3.1005 pd=16.68 as=0 ps=0 w=7.95 l=3.84
X13 VTAIL.t19 VN.t6 VDD2.t3 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=1.31175 pd=8.28 as=1.31175 ps=8.28 w=7.95 l=3.84
X14 VTAIL.t17 VP.t5 VDD1.t4 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=1.31175 pd=8.28 as=1.31175 ps=8.28 w=7.95 l=3.84
X15 B.t5 B.t3 B.t4 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=3.1005 pd=16.68 as=0 ps=0 w=7.95 l=3.84
X16 VTAIL.t13 VP.t6 VDD1.t3 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=1.31175 pd=8.28 as=1.31175 ps=8.28 w=7.95 l=3.84
X17 B.t2 B.t0 B.t1 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=3.1005 pd=16.68 as=0 ps=0 w=7.95 l=3.84
X18 VTAIL.t12 VP.t7 VDD1.t2 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=1.31175 pd=8.28 as=1.31175 ps=8.28 w=7.95 l=3.84
X19 VDD2.t2 VN.t7 VTAIL.t3 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=1.31175 pd=8.28 as=1.31175 ps=8.28 w=7.95 l=3.84
X20 VDD2.t1 VN.t8 VTAIL.t8 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=1.31175 pd=8.28 as=1.31175 ps=8.28 w=7.95 l=3.84
X21 VDD1.t1 VP.t8 VTAIL.t18 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=1.31175 pd=8.28 as=3.1005 ps=16.68 w=7.95 l=3.84
X22 VTAIL.t6 VN.t9 VDD2.t0 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=1.31175 pd=8.28 as=1.31175 ps=8.28 w=7.95 l=3.84
X23 VDD1.t0 VP.t9 VTAIL.t14 w_n5974_n2558# sky130_fd_pr__pfet_01v8 ad=1.31175 pd=8.28 as=1.31175 ps=8.28 w=7.95 l=3.84
R0 VP.n34 VP.n33 161.3
R1 VP.n35 VP.n30 161.3
R2 VP.n37 VP.n36 161.3
R3 VP.n38 VP.n29 161.3
R4 VP.n40 VP.n39 161.3
R5 VP.n41 VP.n28 161.3
R6 VP.n43 VP.n42 161.3
R7 VP.n44 VP.n27 161.3
R8 VP.n47 VP.n46 161.3
R9 VP.n48 VP.n26 161.3
R10 VP.n50 VP.n49 161.3
R11 VP.n51 VP.n25 161.3
R12 VP.n53 VP.n52 161.3
R13 VP.n54 VP.n24 161.3
R14 VP.n56 VP.n55 161.3
R15 VP.n57 VP.n23 161.3
R16 VP.n60 VP.n59 161.3
R17 VP.n61 VP.n22 161.3
R18 VP.n63 VP.n62 161.3
R19 VP.n64 VP.n21 161.3
R20 VP.n66 VP.n65 161.3
R21 VP.n67 VP.n20 161.3
R22 VP.n69 VP.n68 161.3
R23 VP.n70 VP.n19 161.3
R24 VP.n72 VP.n71 161.3
R25 VP.n129 VP.n128 161.3
R26 VP.n127 VP.n1 161.3
R27 VP.n126 VP.n125 161.3
R28 VP.n124 VP.n2 161.3
R29 VP.n123 VP.n122 161.3
R30 VP.n121 VP.n3 161.3
R31 VP.n120 VP.n119 161.3
R32 VP.n118 VP.n4 161.3
R33 VP.n117 VP.n116 161.3
R34 VP.n114 VP.n5 161.3
R35 VP.n113 VP.n112 161.3
R36 VP.n111 VP.n6 161.3
R37 VP.n110 VP.n109 161.3
R38 VP.n108 VP.n7 161.3
R39 VP.n107 VP.n106 161.3
R40 VP.n105 VP.n8 161.3
R41 VP.n104 VP.n103 161.3
R42 VP.n101 VP.n9 161.3
R43 VP.n100 VP.n99 161.3
R44 VP.n98 VP.n10 161.3
R45 VP.n97 VP.n96 161.3
R46 VP.n95 VP.n11 161.3
R47 VP.n94 VP.n93 161.3
R48 VP.n92 VP.n12 161.3
R49 VP.n91 VP.n90 161.3
R50 VP.n88 VP.n13 161.3
R51 VP.n87 VP.n86 161.3
R52 VP.n85 VP.n14 161.3
R53 VP.n84 VP.n83 161.3
R54 VP.n82 VP.n15 161.3
R55 VP.n81 VP.n80 161.3
R56 VP.n79 VP.n16 161.3
R57 VP.n78 VP.n77 161.3
R58 VP.n76 VP.n17 161.3
R59 VP.n75 VP.n74 85.6633
R60 VP.n130 VP.n0 85.6633
R61 VP.n73 VP.n18 85.6633
R62 VP.n31 VP.t2 83.1449
R63 VP.n74 VP.n73 56.8743
R64 VP.n96 VP.n95 56.5193
R65 VP.n109 VP.n108 56.5193
R66 VP.n52 VP.n51 56.5193
R67 VP.n39 VP.n38 56.5193
R68 VP.n32 VP.n31 54.4796
R69 VP.n75 VP.t4 49.895
R70 VP.n89 VP.t1 49.895
R71 VP.n102 VP.t9 49.895
R72 VP.n115 VP.t6 49.895
R73 VP.n0 VP.t3 49.895
R74 VP.n18 VP.t8 49.895
R75 VP.n58 VP.t5 49.895
R76 VP.n45 VP.t0 49.895
R77 VP.n32 VP.t7 49.895
R78 VP.n82 VP.n81 40.979
R79 VP.n122 VP.n2 40.979
R80 VP.n65 VP.n20 40.979
R81 VP.n83 VP.n82 40.0078
R82 VP.n122 VP.n121 40.0078
R83 VP.n65 VP.n64 40.0078
R84 VP.n77 VP.n76 24.4675
R85 VP.n77 VP.n16 24.4675
R86 VP.n81 VP.n16 24.4675
R87 VP.n83 VP.n14 24.4675
R88 VP.n87 VP.n14 24.4675
R89 VP.n88 VP.n87 24.4675
R90 VP.n90 VP.n12 24.4675
R91 VP.n94 VP.n12 24.4675
R92 VP.n95 VP.n94 24.4675
R93 VP.n96 VP.n10 24.4675
R94 VP.n100 VP.n10 24.4675
R95 VP.n101 VP.n100 24.4675
R96 VP.n103 VP.n8 24.4675
R97 VP.n107 VP.n8 24.4675
R98 VP.n108 VP.n107 24.4675
R99 VP.n109 VP.n6 24.4675
R100 VP.n113 VP.n6 24.4675
R101 VP.n114 VP.n113 24.4675
R102 VP.n116 VP.n4 24.4675
R103 VP.n120 VP.n4 24.4675
R104 VP.n121 VP.n120 24.4675
R105 VP.n126 VP.n2 24.4675
R106 VP.n127 VP.n126 24.4675
R107 VP.n128 VP.n127 24.4675
R108 VP.n69 VP.n20 24.4675
R109 VP.n70 VP.n69 24.4675
R110 VP.n71 VP.n70 24.4675
R111 VP.n52 VP.n24 24.4675
R112 VP.n56 VP.n24 24.4675
R113 VP.n57 VP.n56 24.4675
R114 VP.n59 VP.n22 24.4675
R115 VP.n63 VP.n22 24.4675
R116 VP.n64 VP.n63 24.4675
R117 VP.n39 VP.n28 24.4675
R118 VP.n43 VP.n28 24.4675
R119 VP.n44 VP.n43 24.4675
R120 VP.n46 VP.n26 24.4675
R121 VP.n50 VP.n26 24.4675
R122 VP.n51 VP.n50 24.4675
R123 VP.n33 VP.n30 24.4675
R124 VP.n37 VP.n30 24.4675
R125 VP.n38 VP.n37 24.4675
R126 VP.n90 VP.n89 20.5528
R127 VP.n115 VP.n114 20.5528
R128 VP.n58 VP.n57 20.5528
R129 VP.n33 VP.n32 20.5528
R130 VP.n102 VP.n101 12.234
R131 VP.n103 VP.n102 12.234
R132 VP.n45 VP.n44 12.234
R133 VP.n46 VP.n45 12.234
R134 VP.n76 VP.n75 4.40456
R135 VP.n128 VP.n0 4.40456
R136 VP.n71 VP.n18 4.40456
R137 VP.n89 VP.n88 3.91522
R138 VP.n116 VP.n115 3.91522
R139 VP.n59 VP.n58 3.91522
R140 VP.n34 VP.n31 2.43001
R141 VP.n73 VP.n72 0.354971
R142 VP.n74 VP.n17 0.354971
R143 VP.n130 VP.n129 0.354971
R144 VP VP.n130 0.26696
R145 VP.n35 VP.n34 0.189894
R146 VP.n36 VP.n35 0.189894
R147 VP.n36 VP.n29 0.189894
R148 VP.n40 VP.n29 0.189894
R149 VP.n41 VP.n40 0.189894
R150 VP.n42 VP.n41 0.189894
R151 VP.n42 VP.n27 0.189894
R152 VP.n47 VP.n27 0.189894
R153 VP.n48 VP.n47 0.189894
R154 VP.n49 VP.n48 0.189894
R155 VP.n49 VP.n25 0.189894
R156 VP.n53 VP.n25 0.189894
R157 VP.n54 VP.n53 0.189894
R158 VP.n55 VP.n54 0.189894
R159 VP.n55 VP.n23 0.189894
R160 VP.n60 VP.n23 0.189894
R161 VP.n61 VP.n60 0.189894
R162 VP.n62 VP.n61 0.189894
R163 VP.n62 VP.n21 0.189894
R164 VP.n66 VP.n21 0.189894
R165 VP.n67 VP.n66 0.189894
R166 VP.n68 VP.n67 0.189894
R167 VP.n68 VP.n19 0.189894
R168 VP.n72 VP.n19 0.189894
R169 VP.n78 VP.n17 0.189894
R170 VP.n79 VP.n78 0.189894
R171 VP.n80 VP.n79 0.189894
R172 VP.n80 VP.n15 0.189894
R173 VP.n84 VP.n15 0.189894
R174 VP.n85 VP.n84 0.189894
R175 VP.n86 VP.n85 0.189894
R176 VP.n86 VP.n13 0.189894
R177 VP.n91 VP.n13 0.189894
R178 VP.n92 VP.n91 0.189894
R179 VP.n93 VP.n92 0.189894
R180 VP.n93 VP.n11 0.189894
R181 VP.n97 VP.n11 0.189894
R182 VP.n98 VP.n97 0.189894
R183 VP.n99 VP.n98 0.189894
R184 VP.n99 VP.n9 0.189894
R185 VP.n104 VP.n9 0.189894
R186 VP.n105 VP.n104 0.189894
R187 VP.n106 VP.n105 0.189894
R188 VP.n106 VP.n7 0.189894
R189 VP.n110 VP.n7 0.189894
R190 VP.n111 VP.n110 0.189894
R191 VP.n112 VP.n111 0.189894
R192 VP.n112 VP.n5 0.189894
R193 VP.n117 VP.n5 0.189894
R194 VP.n118 VP.n117 0.189894
R195 VP.n119 VP.n118 0.189894
R196 VP.n119 VP.n3 0.189894
R197 VP.n123 VP.n3 0.189894
R198 VP.n124 VP.n123 0.189894
R199 VP.n125 VP.n124 0.189894
R200 VP.n125 VP.n1 0.189894
R201 VP.n129 VP.n1 0.189894
R202 VTAIL.n176 VTAIL.n140 756.745
R203 VTAIL.n38 VTAIL.n2 756.745
R204 VTAIL.n134 VTAIL.n98 756.745
R205 VTAIL.n88 VTAIL.n52 756.745
R206 VTAIL.n152 VTAIL.n151 585
R207 VTAIL.n157 VTAIL.n156 585
R208 VTAIL.n159 VTAIL.n158 585
R209 VTAIL.n148 VTAIL.n147 585
R210 VTAIL.n165 VTAIL.n164 585
R211 VTAIL.n167 VTAIL.n166 585
R212 VTAIL.n144 VTAIL.n143 585
R213 VTAIL.n174 VTAIL.n173 585
R214 VTAIL.n175 VTAIL.n142 585
R215 VTAIL.n177 VTAIL.n176 585
R216 VTAIL.n14 VTAIL.n13 585
R217 VTAIL.n19 VTAIL.n18 585
R218 VTAIL.n21 VTAIL.n20 585
R219 VTAIL.n10 VTAIL.n9 585
R220 VTAIL.n27 VTAIL.n26 585
R221 VTAIL.n29 VTAIL.n28 585
R222 VTAIL.n6 VTAIL.n5 585
R223 VTAIL.n36 VTAIL.n35 585
R224 VTAIL.n37 VTAIL.n4 585
R225 VTAIL.n39 VTAIL.n38 585
R226 VTAIL.n135 VTAIL.n134 585
R227 VTAIL.n133 VTAIL.n100 585
R228 VTAIL.n132 VTAIL.n131 585
R229 VTAIL.n103 VTAIL.n101 585
R230 VTAIL.n126 VTAIL.n125 585
R231 VTAIL.n124 VTAIL.n123 585
R232 VTAIL.n107 VTAIL.n106 585
R233 VTAIL.n118 VTAIL.n117 585
R234 VTAIL.n116 VTAIL.n115 585
R235 VTAIL.n111 VTAIL.n110 585
R236 VTAIL.n89 VTAIL.n88 585
R237 VTAIL.n87 VTAIL.n54 585
R238 VTAIL.n86 VTAIL.n85 585
R239 VTAIL.n57 VTAIL.n55 585
R240 VTAIL.n80 VTAIL.n79 585
R241 VTAIL.n78 VTAIL.n77 585
R242 VTAIL.n61 VTAIL.n60 585
R243 VTAIL.n72 VTAIL.n71 585
R244 VTAIL.n70 VTAIL.n69 585
R245 VTAIL.n65 VTAIL.n64 585
R246 VTAIL.n153 VTAIL.t2 329.043
R247 VTAIL.n15 VTAIL.t11 329.043
R248 VTAIL.n112 VTAIL.t18 329.043
R249 VTAIL.n66 VTAIL.t0 329.043
R250 VTAIL.n157 VTAIL.n151 171.744
R251 VTAIL.n158 VTAIL.n157 171.744
R252 VTAIL.n158 VTAIL.n147 171.744
R253 VTAIL.n165 VTAIL.n147 171.744
R254 VTAIL.n166 VTAIL.n165 171.744
R255 VTAIL.n166 VTAIL.n143 171.744
R256 VTAIL.n174 VTAIL.n143 171.744
R257 VTAIL.n175 VTAIL.n174 171.744
R258 VTAIL.n176 VTAIL.n175 171.744
R259 VTAIL.n19 VTAIL.n13 171.744
R260 VTAIL.n20 VTAIL.n19 171.744
R261 VTAIL.n20 VTAIL.n9 171.744
R262 VTAIL.n27 VTAIL.n9 171.744
R263 VTAIL.n28 VTAIL.n27 171.744
R264 VTAIL.n28 VTAIL.n5 171.744
R265 VTAIL.n36 VTAIL.n5 171.744
R266 VTAIL.n37 VTAIL.n36 171.744
R267 VTAIL.n38 VTAIL.n37 171.744
R268 VTAIL.n134 VTAIL.n133 171.744
R269 VTAIL.n133 VTAIL.n132 171.744
R270 VTAIL.n132 VTAIL.n101 171.744
R271 VTAIL.n125 VTAIL.n101 171.744
R272 VTAIL.n125 VTAIL.n124 171.744
R273 VTAIL.n124 VTAIL.n106 171.744
R274 VTAIL.n117 VTAIL.n106 171.744
R275 VTAIL.n117 VTAIL.n116 171.744
R276 VTAIL.n116 VTAIL.n110 171.744
R277 VTAIL.n88 VTAIL.n87 171.744
R278 VTAIL.n87 VTAIL.n86 171.744
R279 VTAIL.n86 VTAIL.n55 171.744
R280 VTAIL.n79 VTAIL.n55 171.744
R281 VTAIL.n79 VTAIL.n78 171.744
R282 VTAIL.n78 VTAIL.n60 171.744
R283 VTAIL.n71 VTAIL.n60 171.744
R284 VTAIL.n71 VTAIL.n70 171.744
R285 VTAIL.n70 VTAIL.n64 171.744
R286 VTAIL.t2 VTAIL.n151 85.8723
R287 VTAIL.t11 VTAIL.n13 85.8723
R288 VTAIL.t18 VTAIL.n110 85.8723
R289 VTAIL.t0 VTAIL.n64 85.8723
R290 VTAIL.n97 VTAIL.n96 68.5895
R291 VTAIL.n95 VTAIL.n94 68.5895
R292 VTAIL.n51 VTAIL.n50 68.5895
R293 VTAIL.n49 VTAIL.n48 68.5895
R294 VTAIL.n183 VTAIL.n182 68.5894
R295 VTAIL.n1 VTAIL.n0 68.5894
R296 VTAIL.n45 VTAIL.n44 68.5894
R297 VTAIL.n47 VTAIL.n46 68.5894
R298 VTAIL.n181 VTAIL.n180 35.0944
R299 VTAIL.n43 VTAIL.n42 35.0944
R300 VTAIL.n139 VTAIL.n138 35.0944
R301 VTAIL.n93 VTAIL.n92 35.0944
R302 VTAIL.n49 VTAIL.n47 26.41
R303 VTAIL.n181 VTAIL.n139 22.8152
R304 VTAIL.n177 VTAIL.n142 13.1884
R305 VTAIL.n39 VTAIL.n4 13.1884
R306 VTAIL.n135 VTAIL.n100 13.1884
R307 VTAIL.n89 VTAIL.n54 13.1884
R308 VTAIL.n173 VTAIL.n172 12.8005
R309 VTAIL.n178 VTAIL.n140 12.8005
R310 VTAIL.n35 VTAIL.n34 12.8005
R311 VTAIL.n40 VTAIL.n2 12.8005
R312 VTAIL.n136 VTAIL.n98 12.8005
R313 VTAIL.n131 VTAIL.n102 12.8005
R314 VTAIL.n90 VTAIL.n52 12.8005
R315 VTAIL.n85 VTAIL.n56 12.8005
R316 VTAIL.n171 VTAIL.n144 12.0247
R317 VTAIL.n33 VTAIL.n6 12.0247
R318 VTAIL.n130 VTAIL.n103 12.0247
R319 VTAIL.n84 VTAIL.n57 12.0247
R320 VTAIL.n168 VTAIL.n167 11.249
R321 VTAIL.n30 VTAIL.n29 11.249
R322 VTAIL.n127 VTAIL.n126 11.249
R323 VTAIL.n81 VTAIL.n80 11.249
R324 VTAIL.n153 VTAIL.n152 10.7238
R325 VTAIL.n15 VTAIL.n14 10.7238
R326 VTAIL.n112 VTAIL.n111 10.7238
R327 VTAIL.n66 VTAIL.n65 10.7238
R328 VTAIL.n164 VTAIL.n146 10.4732
R329 VTAIL.n26 VTAIL.n8 10.4732
R330 VTAIL.n123 VTAIL.n105 10.4732
R331 VTAIL.n77 VTAIL.n59 10.4732
R332 VTAIL.n163 VTAIL.n148 9.69747
R333 VTAIL.n25 VTAIL.n10 9.69747
R334 VTAIL.n122 VTAIL.n107 9.69747
R335 VTAIL.n76 VTAIL.n61 9.69747
R336 VTAIL.n180 VTAIL.n179 9.45567
R337 VTAIL.n42 VTAIL.n41 9.45567
R338 VTAIL.n138 VTAIL.n137 9.45567
R339 VTAIL.n92 VTAIL.n91 9.45567
R340 VTAIL.n179 VTAIL.n178 9.3005
R341 VTAIL.n155 VTAIL.n154 9.3005
R342 VTAIL.n150 VTAIL.n149 9.3005
R343 VTAIL.n161 VTAIL.n160 9.3005
R344 VTAIL.n163 VTAIL.n162 9.3005
R345 VTAIL.n146 VTAIL.n145 9.3005
R346 VTAIL.n169 VTAIL.n168 9.3005
R347 VTAIL.n171 VTAIL.n170 9.3005
R348 VTAIL.n172 VTAIL.n141 9.3005
R349 VTAIL.n41 VTAIL.n40 9.3005
R350 VTAIL.n17 VTAIL.n16 9.3005
R351 VTAIL.n12 VTAIL.n11 9.3005
R352 VTAIL.n23 VTAIL.n22 9.3005
R353 VTAIL.n25 VTAIL.n24 9.3005
R354 VTAIL.n8 VTAIL.n7 9.3005
R355 VTAIL.n31 VTAIL.n30 9.3005
R356 VTAIL.n33 VTAIL.n32 9.3005
R357 VTAIL.n34 VTAIL.n3 9.3005
R358 VTAIL.n114 VTAIL.n113 9.3005
R359 VTAIL.n109 VTAIL.n108 9.3005
R360 VTAIL.n120 VTAIL.n119 9.3005
R361 VTAIL.n122 VTAIL.n121 9.3005
R362 VTAIL.n105 VTAIL.n104 9.3005
R363 VTAIL.n128 VTAIL.n127 9.3005
R364 VTAIL.n130 VTAIL.n129 9.3005
R365 VTAIL.n102 VTAIL.n99 9.3005
R366 VTAIL.n137 VTAIL.n136 9.3005
R367 VTAIL.n68 VTAIL.n67 9.3005
R368 VTAIL.n63 VTAIL.n62 9.3005
R369 VTAIL.n74 VTAIL.n73 9.3005
R370 VTAIL.n76 VTAIL.n75 9.3005
R371 VTAIL.n59 VTAIL.n58 9.3005
R372 VTAIL.n82 VTAIL.n81 9.3005
R373 VTAIL.n84 VTAIL.n83 9.3005
R374 VTAIL.n56 VTAIL.n53 9.3005
R375 VTAIL.n91 VTAIL.n90 9.3005
R376 VTAIL.n160 VTAIL.n159 8.92171
R377 VTAIL.n22 VTAIL.n21 8.92171
R378 VTAIL.n119 VTAIL.n118 8.92171
R379 VTAIL.n73 VTAIL.n72 8.92171
R380 VTAIL.n156 VTAIL.n150 8.14595
R381 VTAIL.n18 VTAIL.n12 8.14595
R382 VTAIL.n115 VTAIL.n109 8.14595
R383 VTAIL.n69 VTAIL.n63 8.14595
R384 VTAIL.n155 VTAIL.n152 7.3702
R385 VTAIL.n17 VTAIL.n14 7.3702
R386 VTAIL.n114 VTAIL.n111 7.3702
R387 VTAIL.n68 VTAIL.n65 7.3702
R388 VTAIL.n156 VTAIL.n155 5.81868
R389 VTAIL.n18 VTAIL.n17 5.81868
R390 VTAIL.n115 VTAIL.n114 5.81868
R391 VTAIL.n69 VTAIL.n68 5.81868
R392 VTAIL.n159 VTAIL.n150 5.04292
R393 VTAIL.n21 VTAIL.n12 5.04292
R394 VTAIL.n118 VTAIL.n109 5.04292
R395 VTAIL.n72 VTAIL.n63 5.04292
R396 VTAIL.n160 VTAIL.n148 4.26717
R397 VTAIL.n22 VTAIL.n10 4.26717
R398 VTAIL.n119 VTAIL.n107 4.26717
R399 VTAIL.n73 VTAIL.n61 4.26717
R400 VTAIL.n182 VTAIL.t8 4.08918
R401 VTAIL.n182 VTAIL.t5 4.08918
R402 VTAIL.n0 VTAIL.t4 4.08918
R403 VTAIL.n0 VTAIL.t19 4.08918
R404 VTAIL.n44 VTAIL.t14 4.08918
R405 VTAIL.n44 VTAIL.t13 4.08918
R406 VTAIL.n46 VTAIL.t9 4.08918
R407 VTAIL.n46 VTAIL.t16 4.08918
R408 VTAIL.n96 VTAIL.t15 4.08918
R409 VTAIL.n96 VTAIL.t17 4.08918
R410 VTAIL.n94 VTAIL.t10 4.08918
R411 VTAIL.n94 VTAIL.t12 4.08918
R412 VTAIL.n50 VTAIL.t3 4.08918
R413 VTAIL.n50 VTAIL.t6 4.08918
R414 VTAIL.n48 VTAIL.t7 4.08918
R415 VTAIL.n48 VTAIL.t1 4.08918
R416 VTAIL.n51 VTAIL.n49 3.59533
R417 VTAIL.n93 VTAIL.n51 3.59533
R418 VTAIL.n97 VTAIL.n95 3.59533
R419 VTAIL.n139 VTAIL.n97 3.59533
R420 VTAIL.n47 VTAIL.n45 3.59533
R421 VTAIL.n45 VTAIL.n43 3.59533
R422 VTAIL.n183 VTAIL.n181 3.59533
R423 VTAIL.n164 VTAIL.n163 3.49141
R424 VTAIL.n26 VTAIL.n25 3.49141
R425 VTAIL.n123 VTAIL.n122 3.49141
R426 VTAIL.n77 VTAIL.n76 3.49141
R427 VTAIL VTAIL.n1 2.75481
R428 VTAIL.n167 VTAIL.n146 2.71565
R429 VTAIL.n29 VTAIL.n8 2.71565
R430 VTAIL.n126 VTAIL.n105 2.71565
R431 VTAIL.n80 VTAIL.n59 2.71565
R432 VTAIL.n154 VTAIL.n153 2.4129
R433 VTAIL.n16 VTAIL.n15 2.4129
R434 VTAIL.n113 VTAIL.n112 2.4129
R435 VTAIL.n67 VTAIL.n66 2.4129
R436 VTAIL.n95 VTAIL.n93 2.26774
R437 VTAIL.n43 VTAIL.n1 2.26774
R438 VTAIL.n168 VTAIL.n144 1.93989
R439 VTAIL.n30 VTAIL.n6 1.93989
R440 VTAIL.n127 VTAIL.n103 1.93989
R441 VTAIL.n81 VTAIL.n57 1.93989
R442 VTAIL.n173 VTAIL.n171 1.16414
R443 VTAIL.n180 VTAIL.n140 1.16414
R444 VTAIL.n35 VTAIL.n33 1.16414
R445 VTAIL.n42 VTAIL.n2 1.16414
R446 VTAIL.n138 VTAIL.n98 1.16414
R447 VTAIL.n131 VTAIL.n130 1.16414
R448 VTAIL.n92 VTAIL.n52 1.16414
R449 VTAIL.n85 VTAIL.n84 1.16414
R450 VTAIL VTAIL.n183 0.841017
R451 VTAIL.n172 VTAIL.n142 0.388379
R452 VTAIL.n178 VTAIL.n177 0.388379
R453 VTAIL.n34 VTAIL.n4 0.388379
R454 VTAIL.n40 VTAIL.n39 0.388379
R455 VTAIL.n136 VTAIL.n135 0.388379
R456 VTAIL.n102 VTAIL.n100 0.388379
R457 VTAIL.n90 VTAIL.n89 0.388379
R458 VTAIL.n56 VTAIL.n54 0.388379
R459 VTAIL.n154 VTAIL.n149 0.155672
R460 VTAIL.n161 VTAIL.n149 0.155672
R461 VTAIL.n162 VTAIL.n161 0.155672
R462 VTAIL.n162 VTAIL.n145 0.155672
R463 VTAIL.n169 VTAIL.n145 0.155672
R464 VTAIL.n170 VTAIL.n169 0.155672
R465 VTAIL.n170 VTAIL.n141 0.155672
R466 VTAIL.n179 VTAIL.n141 0.155672
R467 VTAIL.n16 VTAIL.n11 0.155672
R468 VTAIL.n23 VTAIL.n11 0.155672
R469 VTAIL.n24 VTAIL.n23 0.155672
R470 VTAIL.n24 VTAIL.n7 0.155672
R471 VTAIL.n31 VTAIL.n7 0.155672
R472 VTAIL.n32 VTAIL.n31 0.155672
R473 VTAIL.n32 VTAIL.n3 0.155672
R474 VTAIL.n41 VTAIL.n3 0.155672
R475 VTAIL.n137 VTAIL.n99 0.155672
R476 VTAIL.n129 VTAIL.n99 0.155672
R477 VTAIL.n129 VTAIL.n128 0.155672
R478 VTAIL.n128 VTAIL.n104 0.155672
R479 VTAIL.n121 VTAIL.n104 0.155672
R480 VTAIL.n121 VTAIL.n120 0.155672
R481 VTAIL.n120 VTAIL.n108 0.155672
R482 VTAIL.n113 VTAIL.n108 0.155672
R483 VTAIL.n91 VTAIL.n53 0.155672
R484 VTAIL.n83 VTAIL.n53 0.155672
R485 VTAIL.n83 VTAIL.n82 0.155672
R486 VTAIL.n82 VTAIL.n58 0.155672
R487 VTAIL.n75 VTAIL.n58 0.155672
R488 VTAIL.n75 VTAIL.n74 0.155672
R489 VTAIL.n74 VTAIL.n62 0.155672
R490 VTAIL.n67 VTAIL.n62 0.155672
R491 VDD1.n36 VDD1.n0 756.745
R492 VDD1.n79 VDD1.n43 756.745
R493 VDD1.n37 VDD1.n36 585
R494 VDD1.n35 VDD1.n2 585
R495 VDD1.n34 VDD1.n33 585
R496 VDD1.n5 VDD1.n3 585
R497 VDD1.n28 VDD1.n27 585
R498 VDD1.n26 VDD1.n25 585
R499 VDD1.n9 VDD1.n8 585
R500 VDD1.n20 VDD1.n19 585
R501 VDD1.n18 VDD1.n17 585
R502 VDD1.n13 VDD1.n12 585
R503 VDD1.n55 VDD1.n54 585
R504 VDD1.n60 VDD1.n59 585
R505 VDD1.n62 VDD1.n61 585
R506 VDD1.n51 VDD1.n50 585
R507 VDD1.n68 VDD1.n67 585
R508 VDD1.n70 VDD1.n69 585
R509 VDD1.n47 VDD1.n46 585
R510 VDD1.n77 VDD1.n76 585
R511 VDD1.n78 VDD1.n45 585
R512 VDD1.n80 VDD1.n79 585
R513 VDD1.n14 VDD1.t7 329.043
R514 VDD1.n56 VDD1.t5 329.043
R515 VDD1.n36 VDD1.n35 171.744
R516 VDD1.n35 VDD1.n34 171.744
R517 VDD1.n34 VDD1.n3 171.744
R518 VDD1.n27 VDD1.n3 171.744
R519 VDD1.n27 VDD1.n26 171.744
R520 VDD1.n26 VDD1.n8 171.744
R521 VDD1.n19 VDD1.n8 171.744
R522 VDD1.n19 VDD1.n18 171.744
R523 VDD1.n18 VDD1.n12 171.744
R524 VDD1.n60 VDD1.n54 171.744
R525 VDD1.n61 VDD1.n60 171.744
R526 VDD1.n61 VDD1.n50 171.744
R527 VDD1.n68 VDD1.n50 171.744
R528 VDD1.n69 VDD1.n68 171.744
R529 VDD1.n69 VDD1.n46 171.744
R530 VDD1.n77 VDD1.n46 171.744
R531 VDD1.n78 VDD1.n77 171.744
R532 VDD1.n79 VDD1.n78 171.744
R533 VDD1.n87 VDD1.n86 87.9089
R534 VDD1.t7 VDD1.n12 85.8723
R535 VDD1.t5 VDD1.n54 85.8723
R536 VDD1.n42 VDD1.n41 85.2683
R537 VDD1.n89 VDD1.n88 85.2682
R538 VDD1.n85 VDD1.n84 85.2682
R539 VDD1.n42 VDD1.n40 55.3681
R540 VDD1.n85 VDD1.n83 55.3681
R541 VDD1.n89 VDD1.n87 50.0246
R542 VDD1.n37 VDD1.n2 13.1884
R543 VDD1.n80 VDD1.n45 13.1884
R544 VDD1.n38 VDD1.n0 12.8005
R545 VDD1.n33 VDD1.n4 12.8005
R546 VDD1.n76 VDD1.n75 12.8005
R547 VDD1.n81 VDD1.n43 12.8005
R548 VDD1.n32 VDD1.n5 12.0247
R549 VDD1.n74 VDD1.n47 12.0247
R550 VDD1.n29 VDD1.n28 11.249
R551 VDD1.n71 VDD1.n70 11.249
R552 VDD1.n14 VDD1.n13 10.7238
R553 VDD1.n56 VDD1.n55 10.7238
R554 VDD1.n25 VDD1.n7 10.4732
R555 VDD1.n67 VDD1.n49 10.4732
R556 VDD1.n24 VDD1.n9 9.69747
R557 VDD1.n66 VDD1.n51 9.69747
R558 VDD1.n40 VDD1.n39 9.45567
R559 VDD1.n83 VDD1.n82 9.45567
R560 VDD1.n16 VDD1.n15 9.3005
R561 VDD1.n11 VDD1.n10 9.3005
R562 VDD1.n22 VDD1.n21 9.3005
R563 VDD1.n24 VDD1.n23 9.3005
R564 VDD1.n7 VDD1.n6 9.3005
R565 VDD1.n30 VDD1.n29 9.3005
R566 VDD1.n32 VDD1.n31 9.3005
R567 VDD1.n4 VDD1.n1 9.3005
R568 VDD1.n39 VDD1.n38 9.3005
R569 VDD1.n82 VDD1.n81 9.3005
R570 VDD1.n58 VDD1.n57 9.3005
R571 VDD1.n53 VDD1.n52 9.3005
R572 VDD1.n64 VDD1.n63 9.3005
R573 VDD1.n66 VDD1.n65 9.3005
R574 VDD1.n49 VDD1.n48 9.3005
R575 VDD1.n72 VDD1.n71 9.3005
R576 VDD1.n74 VDD1.n73 9.3005
R577 VDD1.n75 VDD1.n44 9.3005
R578 VDD1.n21 VDD1.n20 8.92171
R579 VDD1.n63 VDD1.n62 8.92171
R580 VDD1.n17 VDD1.n11 8.14595
R581 VDD1.n59 VDD1.n53 8.14595
R582 VDD1.n16 VDD1.n13 7.3702
R583 VDD1.n58 VDD1.n55 7.3702
R584 VDD1.n17 VDD1.n16 5.81868
R585 VDD1.n59 VDD1.n58 5.81868
R586 VDD1.n20 VDD1.n11 5.04292
R587 VDD1.n62 VDD1.n53 5.04292
R588 VDD1.n21 VDD1.n9 4.26717
R589 VDD1.n63 VDD1.n51 4.26717
R590 VDD1.n88 VDD1.t4 4.08918
R591 VDD1.n88 VDD1.t1 4.08918
R592 VDD1.n41 VDD1.t2 4.08918
R593 VDD1.n41 VDD1.t9 4.08918
R594 VDD1.n86 VDD1.t3 4.08918
R595 VDD1.n86 VDD1.t6 4.08918
R596 VDD1.n84 VDD1.t8 4.08918
R597 VDD1.n84 VDD1.t0 4.08918
R598 VDD1.n25 VDD1.n24 3.49141
R599 VDD1.n67 VDD1.n66 3.49141
R600 VDD1.n28 VDD1.n7 2.71565
R601 VDD1.n70 VDD1.n49 2.71565
R602 VDD1 VDD1.n89 2.63843
R603 VDD1.n15 VDD1.n14 2.4129
R604 VDD1.n57 VDD1.n56 2.4129
R605 VDD1.n29 VDD1.n5 1.93989
R606 VDD1.n71 VDD1.n47 1.93989
R607 VDD1.n40 VDD1.n0 1.16414
R608 VDD1.n33 VDD1.n32 1.16414
R609 VDD1.n76 VDD1.n74 1.16414
R610 VDD1.n83 VDD1.n43 1.16414
R611 VDD1 VDD1.n42 0.957397
R612 VDD1.n87 VDD1.n85 0.843861
R613 VDD1.n38 VDD1.n37 0.388379
R614 VDD1.n4 VDD1.n2 0.388379
R615 VDD1.n75 VDD1.n45 0.388379
R616 VDD1.n81 VDD1.n80 0.388379
R617 VDD1.n39 VDD1.n1 0.155672
R618 VDD1.n31 VDD1.n1 0.155672
R619 VDD1.n31 VDD1.n30 0.155672
R620 VDD1.n30 VDD1.n6 0.155672
R621 VDD1.n23 VDD1.n6 0.155672
R622 VDD1.n23 VDD1.n22 0.155672
R623 VDD1.n22 VDD1.n10 0.155672
R624 VDD1.n15 VDD1.n10 0.155672
R625 VDD1.n57 VDD1.n52 0.155672
R626 VDD1.n64 VDD1.n52 0.155672
R627 VDD1.n65 VDD1.n64 0.155672
R628 VDD1.n65 VDD1.n48 0.155672
R629 VDD1.n72 VDD1.n48 0.155672
R630 VDD1.n73 VDD1.n72 0.155672
R631 VDD1.n73 VDD1.n44 0.155672
R632 VDD1.n82 VDD1.n44 0.155672
R633 VN.n110 VN.n109 161.3
R634 VN.n108 VN.n57 161.3
R635 VN.n107 VN.n106 161.3
R636 VN.n105 VN.n58 161.3
R637 VN.n104 VN.n103 161.3
R638 VN.n102 VN.n59 161.3
R639 VN.n101 VN.n100 161.3
R640 VN.n99 VN.n60 161.3
R641 VN.n98 VN.n97 161.3
R642 VN.n95 VN.n61 161.3
R643 VN.n94 VN.n93 161.3
R644 VN.n92 VN.n62 161.3
R645 VN.n91 VN.n90 161.3
R646 VN.n89 VN.n63 161.3
R647 VN.n88 VN.n87 161.3
R648 VN.n86 VN.n64 161.3
R649 VN.n85 VN.n84 161.3
R650 VN.n82 VN.n65 161.3
R651 VN.n81 VN.n80 161.3
R652 VN.n79 VN.n66 161.3
R653 VN.n78 VN.n77 161.3
R654 VN.n76 VN.n67 161.3
R655 VN.n75 VN.n74 161.3
R656 VN.n73 VN.n68 161.3
R657 VN.n72 VN.n71 161.3
R658 VN.n54 VN.n53 161.3
R659 VN.n52 VN.n1 161.3
R660 VN.n51 VN.n50 161.3
R661 VN.n49 VN.n2 161.3
R662 VN.n48 VN.n47 161.3
R663 VN.n46 VN.n3 161.3
R664 VN.n45 VN.n44 161.3
R665 VN.n43 VN.n4 161.3
R666 VN.n42 VN.n41 161.3
R667 VN.n39 VN.n5 161.3
R668 VN.n38 VN.n37 161.3
R669 VN.n36 VN.n6 161.3
R670 VN.n35 VN.n34 161.3
R671 VN.n33 VN.n7 161.3
R672 VN.n32 VN.n31 161.3
R673 VN.n30 VN.n8 161.3
R674 VN.n29 VN.n28 161.3
R675 VN.n26 VN.n9 161.3
R676 VN.n25 VN.n24 161.3
R677 VN.n23 VN.n10 161.3
R678 VN.n22 VN.n21 161.3
R679 VN.n20 VN.n11 161.3
R680 VN.n19 VN.n18 161.3
R681 VN.n17 VN.n12 161.3
R682 VN.n16 VN.n15 161.3
R683 VN.n55 VN.n0 85.6633
R684 VN.n111 VN.n56 85.6633
R685 VN.n69 VN.t3 83.145
R686 VN.n13 VN.t5 83.145
R687 VN VN.n111 57.0397
R688 VN.n21 VN.n20 56.5193
R689 VN.n34 VN.n33 56.5193
R690 VN.n77 VN.n76 56.5193
R691 VN.n90 VN.n89 56.5193
R692 VN.n14 VN.n13 54.4796
R693 VN.n70 VN.n69 54.4796
R694 VN.n14 VN.t6 49.895
R695 VN.n27 VN.t8 49.895
R696 VN.n40 VN.t1 49.895
R697 VN.n0 VN.t2 49.895
R698 VN.n70 VN.t9 49.895
R699 VN.n83 VN.t7 49.895
R700 VN.n96 VN.t0 49.895
R701 VN.n56 VN.t4 49.895
R702 VN.n47 VN.n2 40.979
R703 VN.n103 VN.n58 40.979
R704 VN.n47 VN.n46 40.0078
R705 VN.n103 VN.n102 40.0078
R706 VN.n15 VN.n12 24.4675
R707 VN.n19 VN.n12 24.4675
R708 VN.n20 VN.n19 24.4675
R709 VN.n21 VN.n10 24.4675
R710 VN.n25 VN.n10 24.4675
R711 VN.n26 VN.n25 24.4675
R712 VN.n28 VN.n8 24.4675
R713 VN.n32 VN.n8 24.4675
R714 VN.n33 VN.n32 24.4675
R715 VN.n34 VN.n6 24.4675
R716 VN.n38 VN.n6 24.4675
R717 VN.n39 VN.n38 24.4675
R718 VN.n41 VN.n4 24.4675
R719 VN.n45 VN.n4 24.4675
R720 VN.n46 VN.n45 24.4675
R721 VN.n51 VN.n2 24.4675
R722 VN.n52 VN.n51 24.4675
R723 VN.n53 VN.n52 24.4675
R724 VN.n76 VN.n75 24.4675
R725 VN.n75 VN.n68 24.4675
R726 VN.n71 VN.n68 24.4675
R727 VN.n89 VN.n88 24.4675
R728 VN.n88 VN.n64 24.4675
R729 VN.n84 VN.n64 24.4675
R730 VN.n82 VN.n81 24.4675
R731 VN.n81 VN.n66 24.4675
R732 VN.n77 VN.n66 24.4675
R733 VN.n102 VN.n101 24.4675
R734 VN.n101 VN.n60 24.4675
R735 VN.n97 VN.n60 24.4675
R736 VN.n95 VN.n94 24.4675
R737 VN.n94 VN.n62 24.4675
R738 VN.n90 VN.n62 24.4675
R739 VN.n109 VN.n108 24.4675
R740 VN.n108 VN.n107 24.4675
R741 VN.n107 VN.n58 24.4675
R742 VN.n15 VN.n14 20.5528
R743 VN.n40 VN.n39 20.5528
R744 VN.n71 VN.n70 20.5528
R745 VN.n96 VN.n95 20.5528
R746 VN.n27 VN.n26 12.234
R747 VN.n28 VN.n27 12.234
R748 VN.n84 VN.n83 12.234
R749 VN.n83 VN.n82 12.234
R750 VN.n53 VN.n0 4.40456
R751 VN.n109 VN.n56 4.40456
R752 VN.n41 VN.n40 3.91522
R753 VN.n97 VN.n96 3.91522
R754 VN.n72 VN.n69 2.43002
R755 VN.n16 VN.n13 2.43002
R756 VN.n111 VN.n110 0.354971
R757 VN.n55 VN.n54 0.354971
R758 VN VN.n55 0.26696
R759 VN.n110 VN.n57 0.189894
R760 VN.n106 VN.n57 0.189894
R761 VN.n106 VN.n105 0.189894
R762 VN.n105 VN.n104 0.189894
R763 VN.n104 VN.n59 0.189894
R764 VN.n100 VN.n59 0.189894
R765 VN.n100 VN.n99 0.189894
R766 VN.n99 VN.n98 0.189894
R767 VN.n98 VN.n61 0.189894
R768 VN.n93 VN.n61 0.189894
R769 VN.n93 VN.n92 0.189894
R770 VN.n92 VN.n91 0.189894
R771 VN.n91 VN.n63 0.189894
R772 VN.n87 VN.n63 0.189894
R773 VN.n87 VN.n86 0.189894
R774 VN.n86 VN.n85 0.189894
R775 VN.n85 VN.n65 0.189894
R776 VN.n80 VN.n65 0.189894
R777 VN.n80 VN.n79 0.189894
R778 VN.n79 VN.n78 0.189894
R779 VN.n78 VN.n67 0.189894
R780 VN.n74 VN.n67 0.189894
R781 VN.n74 VN.n73 0.189894
R782 VN.n73 VN.n72 0.189894
R783 VN.n17 VN.n16 0.189894
R784 VN.n18 VN.n17 0.189894
R785 VN.n18 VN.n11 0.189894
R786 VN.n22 VN.n11 0.189894
R787 VN.n23 VN.n22 0.189894
R788 VN.n24 VN.n23 0.189894
R789 VN.n24 VN.n9 0.189894
R790 VN.n29 VN.n9 0.189894
R791 VN.n30 VN.n29 0.189894
R792 VN.n31 VN.n30 0.189894
R793 VN.n31 VN.n7 0.189894
R794 VN.n35 VN.n7 0.189894
R795 VN.n36 VN.n35 0.189894
R796 VN.n37 VN.n36 0.189894
R797 VN.n37 VN.n5 0.189894
R798 VN.n42 VN.n5 0.189894
R799 VN.n43 VN.n42 0.189894
R800 VN.n44 VN.n43 0.189894
R801 VN.n44 VN.n3 0.189894
R802 VN.n48 VN.n3 0.189894
R803 VN.n49 VN.n48 0.189894
R804 VN.n50 VN.n49 0.189894
R805 VN.n50 VN.n1 0.189894
R806 VN.n54 VN.n1 0.189894
R807 VDD2.n81 VDD2.n45 756.745
R808 VDD2.n36 VDD2.n0 756.745
R809 VDD2.n82 VDD2.n81 585
R810 VDD2.n80 VDD2.n47 585
R811 VDD2.n79 VDD2.n78 585
R812 VDD2.n50 VDD2.n48 585
R813 VDD2.n73 VDD2.n72 585
R814 VDD2.n71 VDD2.n70 585
R815 VDD2.n54 VDD2.n53 585
R816 VDD2.n65 VDD2.n64 585
R817 VDD2.n63 VDD2.n62 585
R818 VDD2.n58 VDD2.n57 585
R819 VDD2.n12 VDD2.n11 585
R820 VDD2.n17 VDD2.n16 585
R821 VDD2.n19 VDD2.n18 585
R822 VDD2.n8 VDD2.n7 585
R823 VDD2.n25 VDD2.n24 585
R824 VDD2.n27 VDD2.n26 585
R825 VDD2.n4 VDD2.n3 585
R826 VDD2.n34 VDD2.n33 585
R827 VDD2.n35 VDD2.n2 585
R828 VDD2.n37 VDD2.n36 585
R829 VDD2.n59 VDD2.t5 329.043
R830 VDD2.n13 VDD2.t4 329.043
R831 VDD2.n81 VDD2.n80 171.744
R832 VDD2.n80 VDD2.n79 171.744
R833 VDD2.n79 VDD2.n48 171.744
R834 VDD2.n72 VDD2.n48 171.744
R835 VDD2.n72 VDD2.n71 171.744
R836 VDD2.n71 VDD2.n53 171.744
R837 VDD2.n64 VDD2.n53 171.744
R838 VDD2.n64 VDD2.n63 171.744
R839 VDD2.n63 VDD2.n57 171.744
R840 VDD2.n17 VDD2.n11 171.744
R841 VDD2.n18 VDD2.n17 171.744
R842 VDD2.n18 VDD2.n7 171.744
R843 VDD2.n25 VDD2.n7 171.744
R844 VDD2.n26 VDD2.n25 171.744
R845 VDD2.n26 VDD2.n3 171.744
R846 VDD2.n34 VDD2.n3 171.744
R847 VDD2.n35 VDD2.n34 171.744
R848 VDD2.n36 VDD2.n35 171.744
R849 VDD2.n44 VDD2.n43 87.9089
R850 VDD2 VDD2.n89 87.9061
R851 VDD2.t5 VDD2.n57 85.8723
R852 VDD2.t4 VDD2.n11 85.8723
R853 VDD2.n88 VDD2.n87 85.2683
R854 VDD2.n42 VDD2.n41 85.2682
R855 VDD2.n42 VDD2.n40 55.3681
R856 VDD2.n86 VDD2.n85 51.7732
R857 VDD2.n86 VDD2.n44 47.6442
R858 VDD2.n82 VDD2.n47 13.1884
R859 VDD2.n37 VDD2.n2 13.1884
R860 VDD2.n83 VDD2.n45 12.8005
R861 VDD2.n78 VDD2.n49 12.8005
R862 VDD2.n33 VDD2.n32 12.8005
R863 VDD2.n38 VDD2.n0 12.8005
R864 VDD2.n77 VDD2.n50 12.0247
R865 VDD2.n31 VDD2.n4 12.0247
R866 VDD2.n74 VDD2.n73 11.249
R867 VDD2.n28 VDD2.n27 11.249
R868 VDD2.n59 VDD2.n58 10.7238
R869 VDD2.n13 VDD2.n12 10.7238
R870 VDD2.n70 VDD2.n52 10.4732
R871 VDD2.n24 VDD2.n6 10.4732
R872 VDD2.n69 VDD2.n54 9.69747
R873 VDD2.n23 VDD2.n8 9.69747
R874 VDD2.n85 VDD2.n84 9.45567
R875 VDD2.n40 VDD2.n39 9.45567
R876 VDD2.n61 VDD2.n60 9.3005
R877 VDD2.n56 VDD2.n55 9.3005
R878 VDD2.n67 VDD2.n66 9.3005
R879 VDD2.n69 VDD2.n68 9.3005
R880 VDD2.n52 VDD2.n51 9.3005
R881 VDD2.n75 VDD2.n74 9.3005
R882 VDD2.n77 VDD2.n76 9.3005
R883 VDD2.n49 VDD2.n46 9.3005
R884 VDD2.n84 VDD2.n83 9.3005
R885 VDD2.n39 VDD2.n38 9.3005
R886 VDD2.n15 VDD2.n14 9.3005
R887 VDD2.n10 VDD2.n9 9.3005
R888 VDD2.n21 VDD2.n20 9.3005
R889 VDD2.n23 VDD2.n22 9.3005
R890 VDD2.n6 VDD2.n5 9.3005
R891 VDD2.n29 VDD2.n28 9.3005
R892 VDD2.n31 VDD2.n30 9.3005
R893 VDD2.n32 VDD2.n1 9.3005
R894 VDD2.n66 VDD2.n65 8.92171
R895 VDD2.n20 VDD2.n19 8.92171
R896 VDD2.n62 VDD2.n56 8.14595
R897 VDD2.n16 VDD2.n10 8.14595
R898 VDD2.n61 VDD2.n58 7.3702
R899 VDD2.n15 VDD2.n12 7.3702
R900 VDD2.n62 VDD2.n61 5.81868
R901 VDD2.n16 VDD2.n15 5.81868
R902 VDD2.n65 VDD2.n56 5.04292
R903 VDD2.n19 VDD2.n10 5.04292
R904 VDD2.n66 VDD2.n54 4.26717
R905 VDD2.n20 VDD2.n8 4.26717
R906 VDD2.n89 VDD2.t0 4.08918
R907 VDD2.n89 VDD2.t6 4.08918
R908 VDD2.n87 VDD2.t9 4.08918
R909 VDD2.n87 VDD2.t2 4.08918
R910 VDD2.n43 VDD2.t8 4.08918
R911 VDD2.n43 VDD2.t7 4.08918
R912 VDD2.n41 VDD2.t3 4.08918
R913 VDD2.n41 VDD2.t1 4.08918
R914 VDD2.n88 VDD2.n86 3.59533
R915 VDD2.n70 VDD2.n69 3.49141
R916 VDD2.n24 VDD2.n23 3.49141
R917 VDD2.n73 VDD2.n52 2.71565
R918 VDD2.n27 VDD2.n6 2.71565
R919 VDD2.n60 VDD2.n59 2.4129
R920 VDD2.n14 VDD2.n13 2.4129
R921 VDD2.n74 VDD2.n50 1.93989
R922 VDD2.n28 VDD2.n4 1.93989
R923 VDD2.n85 VDD2.n45 1.16414
R924 VDD2.n78 VDD2.n77 1.16414
R925 VDD2.n33 VDD2.n31 1.16414
R926 VDD2.n40 VDD2.n0 1.16414
R927 VDD2 VDD2.n88 0.957397
R928 VDD2.n44 VDD2.n42 0.843861
R929 VDD2.n83 VDD2.n82 0.388379
R930 VDD2.n49 VDD2.n47 0.388379
R931 VDD2.n32 VDD2.n2 0.388379
R932 VDD2.n38 VDD2.n37 0.388379
R933 VDD2.n84 VDD2.n46 0.155672
R934 VDD2.n76 VDD2.n46 0.155672
R935 VDD2.n76 VDD2.n75 0.155672
R936 VDD2.n75 VDD2.n51 0.155672
R937 VDD2.n68 VDD2.n51 0.155672
R938 VDD2.n68 VDD2.n67 0.155672
R939 VDD2.n67 VDD2.n55 0.155672
R940 VDD2.n60 VDD2.n55 0.155672
R941 VDD2.n14 VDD2.n9 0.155672
R942 VDD2.n21 VDD2.n9 0.155672
R943 VDD2.n22 VDD2.n21 0.155672
R944 VDD2.n22 VDD2.n5 0.155672
R945 VDD2.n29 VDD2.n5 0.155672
R946 VDD2.n30 VDD2.n29 0.155672
R947 VDD2.n30 VDD2.n1 0.155672
R948 VDD2.n39 VDD2.n1 0.155672
R949 B.n467 B.n466 585
R950 B.n465 B.n164 585
R951 B.n464 B.n463 585
R952 B.n462 B.n165 585
R953 B.n461 B.n460 585
R954 B.n459 B.n166 585
R955 B.n458 B.n457 585
R956 B.n456 B.n167 585
R957 B.n455 B.n454 585
R958 B.n453 B.n168 585
R959 B.n452 B.n451 585
R960 B.n450 B.n169 585
R961 B.n449 B.n448 585
R962 B.n447 B.n170 585
R963 B.n446 B.n445 585
R964 B.n444 B.n171 585
R965 B.n443 B.n442 585
R966 B.n441 B.n172 585
R967 B.n440 B.n439 585
R968 B.n438 B.n173 585
R969 B.n437 B.n436 585
R970 B.n435 B.n174 585
R971 B.n434 B.n433 585
R972 B.n432 B.n175 585
R973 B.n431 B.n430 585
R974 B.n429 B.n176 585
R975 B.n428 B.n427 585
R976 B.n426 B.n177 585
R977 B.n425 B.n424 585
R978 B.n423 B.n178 585
R979 B.n422 B.n421 585
R980 B.n417 B.n179 585
R981 B.n416 B.n415 585
R982 B.n414 B.n180 585
R983 B.n413 B.n412 585
R984 B.n411 B.n181 585
R985 B.n410 B.n409 585
R986 B.n408 B.n182 585
R987 B.n407 B.n406 585
R988 B.n404 B.n183 585
R989 B.n403 B.n402 585
R990 B.n401 B.n186 585
R991 B.n400 B.n399 585
R992 B.n398 B.n187 585
R993 B.n397 B.n396 585
R994 B.n395 B.n188 585
R995 B.n394 B.n393 585
R996 B.n392 B.n189 585
R997 B.n391 B.n390 585
R998 B.n389 B.n190 585
R999 B.n388 B.n387 585
R1000 B.n386 B.n191 585
R1001 B.n385 B.n384 585
R1002 B.n383 B.n192 585
R1003 B.n382 B.n381 585
R1004 B.n380 B.n193 585
R1005 B.n379 B.n378 585
R1006 B.n377 B.n194 585
R1007 B.n376 B.n375 585
R1008 B.n374 B.n195 585
R1009 B.n373 B.n372 585
R1010 B.n371 B.n196 585
R1011 B.n370 B.n369 585
R1012 B.n368 B.n197 585
R1013 B.n367 B.n366 585
R1014 B.n365 B.n198 585
R1015 B.n364 B.n363 585
R1016 B.n362 B.n199 585
R1017 B.n361 B.n360 585
R1018 B.n468 B.n163 585
R1019 B.n470 B.n469 585
R1020 B.n471 B.n162 585
R1021 B.n473 B.n472 585
R1022 B.n474 B.n161 585
R1023 B.n476 B.n475 585
R1024 B.n477 B.n160 585
R1025 B.n479 B.n478 585
R1026 B.n480 B.n159 585
R1027 B.n482 B.n481 585
R1028 B.n483 B.n158 585
R1029 B.n485 B.n484 585
R1030 B.n486 B.n157 585
R1031 B.n488 B.n487 585
R1032 B.n489 B.n156 585
R1033 B.n491 B.n490 585
R1034 B.n492 B.n155 585
R1035 B.n494 B.n493 585
R1036 B.n495 B.n154 585
R1037 B.n497 B.n496 585
R1038 B.n498 B.n153 585
R1039 B.n500 B.n499 585
R1040 B.n501 B.n152 585
R1041 B.n503 B.n502 585
R1042 B.n504 B.n151 585
R1043 B.n506 B.n505 585
R1044 B.n507 B.n150 585
R1045 B.n509 B.n508 585
R1046 B.n510 B.n149 585
R1047 B.n512 B.n511 585
R1048 B.n513 B.n148 585
R1049 B.n515 B.n514 585
R1050 B.n516 B.n147 585
R1051 B.n518 B.n517 585
R1052 B.n519 B.n146 585
R1053 B.n521 B.n520 585
R1054 B.n522 B.n145 585
R1055 B.n524 B.n523 585
R1056 B.n525 B.n144 585
R1057 B.n527 B.n526 585
R1058 B.n528 B.n143 585
R1059 B.n530 B.n529 585
R1060 B.n531 B.n142 585
R1061 B.n533 B.n532 585
R1062 B.n534 B.n141 585
R1063 B.n536 B.n535 585
R1064 B.n537 B.n140 585
R1065 B.n539 B.n538 585
R1066 B.n540 B.n139 585
R1067 B.n542 B.n541 585
R1068 B.n543 B.n138 585
R1069 B.n545 B.n544 585
R1070 B.n546 B.n137 585
R1071 B.n548 B.n547 585
R1072 B.n549 B.n136 585
R1073 B.n551 B.n550 585
R1074 B.n552 B.n135 585
R1075 B.n554 B.n553 585
R1076 B.n555 B.n134 585
R1077 B.n557 B.n556 585
R1078 B.n558 B.n133 585
R1079 B.n560 B.n559 585
R1080 B.n561 B.n132 585
R1081 B.n563 B.n562 585
R1082 B.n564 B.n131 585
R1083 B.n566 B.n565 585
R1084 B.n567 B.n130 585
R1085 B.n569 B.n568 585
R1086 B.n570 B.n129 585
R1087 B.n572 B.n571 585
R1088 B.n573 B.n128 585
R1089 B.n575 B.n574 585
R1090 B.n576 B.n127 585
R1091 B.n578 B.n577 585
R1092 B.n579 B.n126 585
R1093 B.n581 B.n580 585
R1094 B.n582 B.n125 585
R1095 B.n584 B.n583 585
R1096 B.n585 B.n124 585
R1097 B.n587 B.n586 585
R1098 B.n588 B.n123 585
R1099 B.n590 B.n589 585
R1100 B.n591 B.n122 585
R1101 B.n593 B.n592 585
R1102 B.n594 B.n121 585
R1103 B.n596 B.n595 585
R1104 B.n597 B.n120 585
R1105 B.n599 B.n598 585
R1106 B.n600 B.n119 585
R1107 B.n602 B.n601 585
R1108 B.n603 B.n118 585
R1109 B.n605 B.n604 585
R1110 B.n606 B.n117 585
R1111 B.n608 B.n607 585
R1112 B.n609 B.n116 585
R1113 B.n611 B.n610 585
R1114 B.n612 B.n115 585
R1115 B.n614 B.n613 585
R1116 B.n615 B.n114 585
R1117 B.n617 B.n616 585
R1118 B.n618 B.n113 585
R1119 B.n620 B.n619 585
R1120 B.n621 B.n112 585
R1121 B.n623 B.n622 585
R1122 B.n624 B.n111 585
R1123 B.n626 B.n625 585
R1124 B.n627 B.n110 585
R1125 B.n629 B.n628 585
R1126 B.n630 B.n109 585
R1127 B.n632 B.n631 585
R1128 B.n633 B.n108 585
R1129 B.n635 B.n634 585
R1130 B.n636 B.n107 585
R1131 B.n638 B.n637 585
R1132 B.n639 B.n106 585
R1133 B.n641 B.n640 585
R1134 B.n642 B.n105 585
R1135 B.n644 B.n643 585
R1136 B.n645 B.n104 585
R1137 B.n647 B.n646 585
R1138 B.n648 B.n103 585
R1139 B.n650 B.n649 585
R1140 B.n651 B.n102 585
R1141 B.n653 B.n652 585
R1142 B.n654 B.n101 585
R1143 B.n656 B.n655 585
R1144 B.n657 B.n100 585
R1145 B.n659 B.n658 585
R1146 B.n660 B.n99 585
R1147 B.n662 B.n661 585
R1148 B.n663 B.n98 585
R1149 B.n665 B.n664 585
R1150 B.n666 B.n97 585
R1151 B.n668 B.n667 585
R1152 B.n669 B.n96 585
R1153 B.n671 B.n670 585
R1154 B.n672 B.n95 585
R1155 B.n674 B.n673 585
R1156 B.n675 B.n94 585
R1157 B.n677 B.n676 585
R1158 B.n678 B.n93 585
R1159 B.n680 B.n679 585
R1160 B.n681 B.n92 585
R1161 B.n683 B.n682 585
R1162 B.n684 B.n91 585
R1163 B.n686 B.n685 585
R1164 B.n687 B.n90 585
R1165 B.n689 B.n688 585
R1166 B.n690 B.n89 585
R1167 B.n692 B.n691 585
R1168 B.n693 B.n88 585
R1169 B.n695 B.n694 585
R1170 B.n696 B.n87 585
R1171 B.n698 B.n697 585
R1172 B.n699 B.n86 585
R1173 B.n701 B.n700 585
R1174 B.n702 B.n85 585
R1175 B.n704 B.n703 585
R1176 B.n705 B.n84 585
R1177 B.n707 B.n706 585
R1178 B.n708 B.n83 585
R1179 B.n710 B.n709 585
R1180 B.n711 B.n82 585
R1181 B.n713 B.n712 585
R1182 B.n818 B.n817 585
R1183 B.n816 B.n43 585
R1184 B.n815 B.n814 585
R1185 B.n813 B.n44 585
R1186 B.n812 B.n811 585
R1187 B.n810 B.n45 585
R1188 B.n809 B.n808 585
R1189 B.n807 B.n46 585
R1190 B.n806 B.n805 585
R1191 B.n804 B.n47 585
R1192 B.n803 B.n802 585
R1193 B.n801 B.n48 585
R1194 B.n800 B.n799 585
R1195 B.n798 B.n49 585
R1196 B.n797 B.n796 585
R1197 B.n795 B.n50 585
R1198 B.n794 B.n793 585
R1199 B.n792 B.n51 585
R1200 B.n791 B.n790 585
R1201 B.n789 B.n52 585
R1202 B.n788 B.n787 585
R1203 B.n786 B.n53 585
R1204 B.n785 B.n784 585
R1205 B.n783 B.n54 585
R1206 B.n782 B.n781 585
R1207 B.n780 B.n55 585
R1208 B.n779 B.n778 585
R1209 B.n777 B.n56 585
R1210 B.n776 B.n775 585
R1211 B.n774 B.n57 585
R1212 B.n772 B.n771 585
R1213 B.n770 B.n60 585
R1214 B.n769 B.n768 585
R1215 B.n767 B.n61 585
R1216 B.n766 B.n765 585
R1217 B.n764 B.n62 585
R1218 B.n763 B.n762 585
R1219 B.n761 B.n63 585
R1220 B.n760 B.n759 585
R1221 B.n758 B.n757 585
R1222 B.n756 B.n67 585
R1223 B.n755 B.n754 585
R1224 B.n753 B.n68 585
R1225 B.n752 B.n751 585
R1226 B.n750 B.n69 585
R1227 B.n749 B.n748 585
R1228 B.n747 B.n70 585
R1229 B.n746 B.n745 585
R1230 B.n744 B.n71 585
R1231 B.n743 B.n742 585
R1232 B.n741 B.n72 585
R1233 B.n740 B.n739 585
R1234 B.n738 B.n73 585
R1235 B.n737 B.n736 585
R1236 B.n735 B.n74 585
R1237 B.n734 B.n733 585
R1238 B.n732 B.n75 585
R1239 B.n731 B.n730 585
R1240 B.n729 B.n76 585
R1241 B.n728 B.n727 585
R1242 B.n726 B.n77 585
R1243 B.n725 B.n724 585
R1244 B.n723 B.n78 585
R1245 B.n722 B.n721 585
R1246 B.n720 B.n79 585
R1247 B.n719 B.n718 585
R1248 B.n717 B.n80 585
R1249 B.n716 B.n715 585
R1250 B.n714 B.n81 585
R1251 B.n819 B.n42 585
R1252 B.n821 B.n820 585
R1253 B.n822 B.n41 585
R1254 B.n824 B.n823 585
R1255 B.n825 B.n40 585
R1256 B.n827 B.n826 585
R1257 B.n828 B.n39 585
R1258 B.n830 B.n829 585
R1259 B.n831 B.n38 585
R1260 B.n833 B.n832 585
R1261 B.n834 B.n37 585
R1262 B.n836 B.n835 585
R1263 B.n837 B.n36 585
R1264 B.n839 B.n838 585
R1265 B.n840 B.n35 585
R1266 B.n842 B.n841 585
R1267 B.n843 B.n34 585
R1268 B.n845 B.n844 585
R1269 B.n846 B.n33 585
R1270 B.n848 B.n847 585
R1271 B.n849 B.n32 585
R1272 B.n851 B.n850 585
R1273 B.n852 B.n31 585
R1274 B.n854 B.n853 585
R1275 B.n855 B.n30 585
R1276 B.n857 B.n856 585
R1277 B.n858 B.n29 585
R1278 B.n860 B.n859 585
R1279 B.n861 B.n28 585
R1280 B.n863 B.n862 585
R1281 B.n864 B.n27 585
R1282 B.n866 B.n865 585
R1283 B.n867 B.n26 585
R1284 B.n869 B.n868 585
R1285 B.n870 B.n25 585
R1286 B.n872 B.n871 585
R1287 B.n873 B.n24 585
R1288 B.n875 B.n874 585
R1289 B.n876 B.n23 585
R1290 B.n878 B.n877 585
R1291 B.n879 B.n22 585
R1292 B.n881 B.n880 585
R1293 B.n882 B.n21 585
R1294 B.n884 B.n883 585
R1295 B.n885 B.n20 585
R1296 B.n887 B.n886 585
R1297 B.n888 B.n19 585
R1298 B.n890 B.n889 585
R1299 B.n891 B.n18 585
R1300 B.n893 B.n892 585
R1301 B.n894 B.n17 585
R1302 B.n896 B.n895 585
R1303 B.n897 B.n16 585
R1304 B.n899 B.n898 585
R1305 B.n900 B.n15 585
R1306 B.n902 B.n901 585
R1307 B.n903 B.n14 585
R1308 B.n905 B.n904 585
R1309 B.n906 B.n13 585
R1310 B.n908 B.n907 585
R1311 B.n909 B.n12 585
R1312 B.n911 B.n910 585
R1313 B.n912 B.n11 585
R1314 B.n914 B.n913 585
R1315 B.n915 B.n10 585
R1316 B.n917 B.n916 585
R1317 B.n918 B.n9 585
R1318 B.n920 B.n919 585
R1319 B.n921 B.n8 585
R1320 B.n923 B.n922 585
R1321 B.n924 B.n7 585
R1322 B.n926 B.n925 585
R1323 B.n927 B.n6 585
R1324 B.n929 B.n928 585
R1325 B.n930 B.n5 585
R1326 B.n932 B.n931 585
R1327 B.n933 B.n4 585
R1328 B.n935 B.n934 585
R1329 B.n936 B.n3 585
R1330 B.n938 B.n937 585
R1331 B.n939 B.n0 585
R1332 B.n2 B.n1 585
R1333 B.n241 B.n240 585
R1334 B.n242 B.n239 585
R1335 B.n244 B.n243 585
R1336 B.n245 B.n238 585
R1337 B.n247 B.n246 585
R1338 B.n248 B.n237 585
R1339 B.n250 B.n249 585
R1340 B.n251 B.n236 585
R1341 B.n253 B.n252 585
R1342 B.n254 B.n235 585
R1343 B.n256 B.n255 585
R1344 B.n257 B.n234 585
R1345 B.n259 B.n258 585
R1346 B.n260 B.n233 585
R1347 B.n262 B.n261 585
R1348 B.n263 B.n232 585
R1349 B.n265 B.n264 585
R1350 B.n266 B.n231 585
R1351 B.n268 B.n267 585
R1352 B.n269 B.n230 585
R1353 B.n271 B.n270 585
R1354 B.n272 B.n229 585
R1355 B.n274 B.n273 585
R1356 B.n275 B.n228 585
R1357 B.n277 B.n276 585
R1358 B.n278 B.n227 585
R1359 B.n280 B.n279 585
R1360 B.n281 B.n226 585
R1361 B.n283 B.n282 585
R1362 B.n284 B.n225 585
R1363 B.n286 B.n285 585
R1364 B.n287 B.n224 585
R1365 B.n289 B.n288 585
R1366 B.n290 B.n223 585
R1367 B.n292 B.n291 585
R1368 B.n293 B.n222 585
R1369 B.n295 B.n294 585
R1370 B.n296 B.n221 585
R1371 B.n298 B.n297 585
R1372 B.n299 B.n220 585
R1373 B.n301 B.n300 585
R1374 B.n302 B.n219 585
R1375 B.n304 B.n303 585
R1376 B.n305 B.n218 585
R1377 B.n307 B.n306 585
R1378 B.n308 B.n217 585
R1379 B.n310 B.n309 585
R1380 B.n311 B.n216 585
R1381 B.n313 B.n312 585
R1382 B.n314 B.n215 585
R1383 B.n316 B.n315 585
R1384 B.n317 B.n214 585
R1385 B.n319 B.n318 585
R1386 B.n320 B.n213 585
R1387 B.n322 B.n321 585
R1388 B.n323 B.n212 585
R1389 B.n325 B.n324 585
R1390 B.n326 B.n211 585
R1391 B.n328 B.n327 585
R1392 B.n329 B.n210 585
R1393 B.n331 B.n330 585
R1394 B.n332 B.n209 585
R1395 B.n334 B.n333 585
R1396 B.n335 B.n208 585
R1397 B.n337 B.n336 585
R1398 B.n338 B.n207 585
R1399 B.n340 B.n339 585
R1400 B.n341 B.n206 585
R1401 B.n343 B.n342 585
R1402 B.n344 B.n205 585
R1403 B.n346 B.n345 585
R1404 B.n347 B.n204 585
R1405 B.n349 B.n348 585
R1406 B.n350 B.n203 585
R1407 B.n352 B.n351 585
R1408 B.n353 B.n202 585
R1409 B.n355 B.n354 585
R1410 B.n356 B.n201 585
R1411 B.n358 B.n357 585
R1412 B.n359 B.n200 585
R1413 B.n360 B.n359 530.939
R1414 B.n466 B.n163 530.939
R1415 B.n712 B.n81 530.939
R1416 B.n819 B.n818 530.939
R1417 B.n418 B.t7 383.594
R1418 B.n64 B.t5 383.594
R1419 B.n184 B.t1 383.594
R1420 B.n58 B.t11 383.594
R1421 B.n419 B.t8 302.721
R1422 B.n65 B.t4 302.721
R1423 B.n185 B.t2 302.721
R1424 B.n59 B.t10 302.721
R1425 B.n184 B.t0 259.269
R1426 B.n418 B.t6 259.269
R1427 B.n64 B.t3 259.269
R1428 B.n58 B.t9 259.269
R1429 B.n941 B.n940 256.663
R1430 B.n940 B.n939 235.042
R1431 B.n940 B.n2 235.042
R1432 B.n360 B.n199 163.367
R1433 B.n364 B.n199 163.367
R1434 B.n365 B.n364 163.367
R1435 B.n366 B.n365 163.367
R1436 B.n366 B.n197 163.367
R1437 B.n370 B.n197 163.367
R1438 B.n371 B.n370 163.367
R1439 B.n372 B.n371 163.367
R1440 B.n372 B.n195 163.367
R1441 B.n376 B.n195 163.367
R1442 B.n377 B.n376 163.367
R1443 B.n378 B.n377 163.367
R1444 B.n378 B.n193 163.367
R1445 B.n382 B.n193 163.367
R1446 B.n383 B.n382 163.367
R1447 B.n384 B.n383 163.367
R1448 B.n384 B.n191 163.367
R1449 B.n388 B.n191 163.367
R1450 B.n389 B.n388 163.367
R1451 B.n390 B.n389 163.367
R1452 B.n390 B.n189 163.367
R1453 B.n394 B.n189 163.367
R1454 B.n395 B.n394 163.367
R1455 B.n396 B.n395 163.367
R1456 B.n396 B.n187 163.367
R1457 B.n400 B.n187 163.367
R1458 B.n401 B.n400 163.367
R1459 B.n402 B.n401 163.367
R1460 B.n402 B.n183 163.367
R1461 B.n407 B.n183 163.367
R1462 B.n408 B.n407 163.367
R1463 B.n409 B.n408 163.367
R1464 B.n409 B.n181 163.367
R1465 B.n413 B.n181 163.367
R1466 B.n414 B.n413 163.367
R1467 B.n415 B.n414 163.367
R1468 B.n415 B.n179 163.367
R1469 B.n422 B.n179 163.367
R1470 B.n423 B.n422 163.367
R1471 B.n424 B.n423 163.367
R1472 B.n424 B.n177 163.367
R1473 B.n428 B.n177 163.367
R1474 B.n429 B.n428 163.367
R1475 B.n430 B.n429 163.367
R1476 B.n430 B.n175 163.367
R1477 B.n434 B.n175 163.367
R1478 B.n435 B.n434 163.367
R1479 B.n436 B.n435 163.367
R1480 B.n436 B.n173 163.367
R1481 B.n440 B.n173 163.367
R1482 B.n441 B.n440 163.367
R1483 B.n442 B.n441 163.367
R1484 B.n442 B.n171 163.367
R1485 B.n446 B.n171 163.367
R1486 B.n447 B.n446 163.367
R1487 B.n448 B.n447 163.367
R1488 B.n448 B.n169 163.367
R1489 B.n452 B.n169 163.367
R1490 B.n453 B.n452 163.367
R1491 B.n454 B.n453 163.367
R1492 B.n454 B.n167 163.367
R1493 B.n458 B.n167 163.367
R1494 B.n459 B.n458 163.367
R1495 B.n460 B.n459 163.367
R1496 B.n460 B.n165 163.367
R1497 B.n464 B.n165 163.367
R1498 B.n465 B.n464 163.367
R1499 B.n466 B.n465 163.367
R1500 B.n712 B.n711 163.367
R1501 B.n711 B.n710 163.367
R1502 B.n710 B.n83 163.367
R1503 B.n706 B.n83 163.367
R1504 B.n706 B.n705 163.367
R1505 B.n705 B.n704 163.367
R1506 B.n704 B.n85 163.367
R1507 B.n700 B.n85 163.367
R1508 B.n700 B.n699 163.367
R1509 B.n699 B.n698 163.367
R1510 B.n698 B.n87 163.367
R1511 B.n694 B.n87 163.367
R1512 B.n694 B.n693 163.367
R1513 B.n693 B.n692 163.367
R1514 B.n692 B.n89 163.367
R1515 B.n688 B.n89 163.367
R1516 B.n688 B.n687 163.367
R1517 B.n687 B.n686 163.367
R1518 B.n686 B.n91 163.367
R1519 B.n682 B.n91 163.367
R1520 B.n682 B.n681 163.367
R1521 B.n681 B.n680 163.367
R1522 B.n680 B.n93 163.367
R1523 B.n676 B.n93 163.367
R1524 B.n676 B.n675 163.367
R1525 B.n675 B.n674 163.367
R1526 B.n674 B.n95 163.367
R1527 B.n670 B.n95 163.367
R1528 B.n670 B.n669 163.367
R1529 B.n669 B.n668 163.367
R1530 B.n668 B.n97 163.367
R1531 B.n664 B.n97 163.367
R1532 B.n664 B.n663 163.367
R1533 B.n663 B.n662 163.367
R1534 B.n662 B.n99 163.367
R1535 B.n658 B.n99 163.367
R1536 B.n658 B.n657 163.367
R1537 B.n657 B.n656 163.367
R1538 B.n656 B.n101 163.367
R1539 B.n652 B.n101 163.367
R1540 B.n652 B.n651 163.367
R1541 B.n651 B.n650 163.367
R1542 B.n650 B.n103 163.367
R1543 B.n646 B.n103 163.367
R1544 B.n646 B.n645 163.367
R1545 B.n645 B.n644 163.367
R1546 B.n644 B.n105 163.367
R1547 B.n640 B.n105 163.367
R1548 B.n640 B.n639 163.367
R1549 B.n639 B.n638 163.367
R1550 B.n638 B.n107 163.367
R1551 B.n634 B.n107 163.367
R1552 B.n634 B.n633 163.367
R1553 B.n633 B.n632 163.367
R1554 B.n632 B.n109 163.367
R1555 B.n628 B.n109 163.367
R1556 B.n628 B.n627 163.367
R1557 B.n627 B.n626 163.367
R1558 B.n626 B.n111 163.367
R1559 B.n622 B.n111 163.367
R1560 B.n622 B.n621 163.367
R1561 B.n621 B.n620 163.367
R1562 B.n620 B.n113 163.367
R1563 B.n616 B.n113 163.367
R1564 B.n616 B.n615 163.367
R1565 B.n615 B.n614 163.367
R1566 B.n614 B.n115 163.367
R1567 B.n610 B.n115 163.367
R1568 B.n610 B.n609 163.367
R1569 B.n609 B.n608 163.367
R1570 B.n608 B.n117 163.367
R1571 B.n604 B.n117 163.367
R1572 B.n604 B.n603 163.367
R1573 B.n603 B.n602 163.367
R1574 B.n602 B.n119 163.367
R1575 B.n598 B.n119 163.367
R1576 B.n598 B.n597 163.367
R1577 B.n597 B.n596 163.367
R1578 B.n596 B.n121 163.367
R1579 B.n592 B.n121 163.367
R1580 B.n592 B.n591 163.367
R1581 B.n591 B.n590 163.367
R1582 B.n590 B.n123 163.367
R1583 B.n586 B.n123 163.367
R1584 B.n586 B.n585 163.367
R1585 B.n585 B.n584 163.367
R1586 B.n584 B.n125 163.367
R1587 B.n580 B.n125 163.367
R1588 B.n580 B.n579 163.367
R1589 B.n579 B.n578 163.367
R1590 B.n578 B.n127 163.367
R1591 B.n574 B.n127 163.367
R1592 B.n574 B.n573 163.367
R1593 B.n573 B.n572 163.367
R1594 B.n572 B.n129 163.367
R1595 B.n568 B.n129 163.367
R1596 B.n568 B.n567 163.367
R1597 B.n567 B.n566 163.367
R1598 B.n566 B.n131 163.367
R1599 B.n562 B.n131 163.367
R1600 B.n562 B.n561 163.367
R1601 B.n561 B.n560 163.367
R1602 B.n560 B.n133 163.367
R1603 B.n556 B.n133 163.367
R1604 B.n556 B.n555 163.367
R1605 B.n555 B.n554 163.367
R1606 B.n554 B.n135 163.367
R1607 B.n550 B.n135 163.367
R1608 B.n550 B.n549 163.367
R1609 B.n549 B.n548 163.367
R1610 B.n548 B.n137 163.367
R1611 B.n544 B.n137 163.367
R1612 B.n544 B.n543 163.367
R1613 B.n543 B.n542 163.367
R1614 B.n542 B.n139 163.367
R1615 B.n538 B.n139 163.367
R1616 B.n538 B.n537 163.367
R1617 B.n537 B.n536 163.367
R1618 B.n536 B.n141 163.367
R1619 B.n532 B.n141 163.367
R1620 B.n532 B.n531 163.367
R1621 B.n531 B.n530 163.367
R1622 B.n530 B.n143 163.367
R1623 B.n526 B.n143 163.367
R1624 B.n526 B.n525 163.367
R1625 B.n525 B.n524 163.367
R1626 B.n524 B.n145 163.367
R1627 B.n520 B.n145 163.367
R1628 B.n520 B.n519 163.367
R1629 B.n519 B.n518 163.367
R1630 B.n518 B.n147 163.367
R1631 B.n514 B.n147 163.367
R1632 B.n514 B.n513 163.367
R1633 B.n513 B.n512 163.367
R1634 B.n512 B.n149 163.367
R1635 B.n508 B.n149 163.367
R1636 B.n508 B.n507 163.367
R1637 B.n507 B.n506 163.367
R1638 B.n506 B.n151 163.367
R1639 B.n502 B.n151 163.367
R1640 B.n502 B.n501 163.367
R1641 B.n501 B.n500 163.367
R1642 B.n500 B.n153 163.367
R1643 B.n496 B.n153 163.367
R1644 B.n496 B.n495 163.367
R1645 B.n495 B.n494 163.367
R1646 B.n494 B.n155 163.367
R1647 B.n490 B.n155 163.367
R1648 B.n490 B.n489 163.367
R1649 B.n489 B.n488 163.367
R1650 B.n488 B.n157 163.367
R1651 B.n484 B.n157 163.367
R1652 B.n484 B.n483 163.367
R1653 B.n483 B.n482 163.367
R1654 B.n482 B.n159 163.367
R1655 B.n478 B.n159 163.367
R1656 B.n478 B.n477 163.367
R1657 B.n477 B.n476 163.367
R1658 B.n476 B.n161 163.367
R1659 B.n472 B.n161 163.367
R1660 B.n472 B.n471 163.367
R1661 B.n471 B.n470 163.367
R1662 B.n470 B.n163 163.367
R1663 B.n818 B.n43 163.367
R1664 B.n814 B.n43 163.367
R1665 B.n814 B.n813 163.367
R1666 B.n813 B.n812 163.367
R1667 B.n812 B.n45 163.367
R1668 B.n808 B.n45 163.367
R1669 B.n808 B.n807 163.367
R1670 B.n807 B.n806 163.367
R1671 B.n806 B.n47 163.367
R1672 B.n802 B.n47 163.367
R1673 B.n802 B.n801 163.367
R1674 B.n801 B.n800 163.367
R1675 B.n800 B.n49 163.367
R1676 B.n796 B.n49 163.367
R1677 B.n796 B.n795 163.367
R1678 B.n795 B.n794 163.367
R1679 B.n794 B.n51 163.367
R1680 B.n790 B.n51 163.367
R1681 B.n790 B.n789 163.367
R1682 B.n789 B.n788 163.367
R1683 B.n788 B.n53 163.367
R1684 B.n784 B.n53 163.367
R1685 B.n784 B.n783 163.367
R1686 B.n783 B.n782 163.367
R1687 B.n782 B.n55 163.367
R1688 B.n778 B.n55 163.367
R1689 B.n778 B.n777 163.367
R1690 B.n777 B.n776 163.367
R1691 B.n776 B.n57 163.367
R1692 B.n771 B.n57 163.367
R1693 B.n771 B.n770 163.367
R1694 B.n770 B.n769 163.367
R1695 B.n769 B.n61 163.367
R1696 B.n765 B.n61 163.367
R1697 B.n765 B.n764 163.367
R1698 B.n764 B.n763 163.367
R1699 B.n763 B.n63 163.367
R1700 B.n759 B.n63 163.367
R1701 B.n759 B.n758 163.367
R1702 B.n758 B.n67 163.367
R1703 B.n754 B.n67 163.367
R1704 B.n754 B.n753 163.367
R1705 B.n753 B.n752 163.367
R1706 B.n752 B.n69 163.367
R1707 B.n748 B.n69 163.367
R1708 B.n748 B.n747 163.367
R1709 B.n747 B.n746 163.367
R1710 B.n746 B.n71 163.367
R1711 B.n742 B.n71 163.367
R1712 B.n742 B.n741 163.367
R1713 B.n741 B.n740 163.367
R1714 B.n740 B.n73 163.367
R1715 B.n736 B.n73 163.367
R1716 B.n736 B.n735 163.367
R1717 B.n735 B.n734 163.367
R1718 B.n734 B.n75 163.367
R1719 B.n730 B.n75 163.367
R1720 B.n730 B.n729 163.367
R1721 B.n729 B.n728 163.367
R1722 B.n728 B.n77 163.367
R1723 B.n724 B.n77 163.367
R1724 B.n724 B.n723 163.367
R1725 B.n723 B.n722 163.367
R1726 B.n722 B.n79 163.367
R1727 B.n718 B.n79 163.367
R1728 B.n718 B.n717 163.367
R1729 B.n717 B.n716 163.367
R1730 B.n716 B.n81 163.367
R1731 B.n820 B.n819 163.367
R1732 B.n820 B.n41 163.367
R1733 B.n824 B.n41 163.367
R1734 B.n825 B.n824 163.367
R1735 B.n826 B.n825 163.367
R1736 B.n826 B.n39 163.367
R1737 B.n830 B.n39 163.367
R1738 B.n831 B.n830 163.367
R1739 B.n832 B.n831 163.367
R1740 B.n832 B.n37 163.367
R1741 B.n836 B.n37 163.367
R1742 B.n837 B.n836 163.367
R1743 B.n838 B.n837 163.367
R1744 B.n838 B.n35 163.367
R1745 B.n842 B.n35 163.367
R1746 B.n843 B.n842 163.367
R1747 B.n844 B.n843 163.367
R1748 B.n844 B.n33 163.367
R1749 B.n848 B.n33 163.367
R1750 B.n849 B.n848 163.367
R1751 B.n850 B.n849 163.367
R1752 B.n850 B.n31 163.367
R1753 B.n854 B.n31 163.367
R1754 B.n855 B.n854 163.367
R1755 B.n856 B.n855 163.367
R1756 B.n856 B.n29 163.367
R1757 B.n860 B.n29 163.367
R1758 B.n861 B.n860 163.367
R1759 B.n862 B.n861 163.367
R1760 B.n862 B.n27 163.367
R1761 B.n866 B.n27 163.367
R1762 B.n867 B.n866 163.367
R1763 B.n868 B.n867 163.367
R1764 B.n868 B.n25 163.367
R1765 B.n872 B.n25 163.367
R1766 B.n873 B.n872 163.367
R1767 B.n874 B.n873 163.367
R1768 B.n874 B.n23 163.367
R1769 B.n878 B.n23 163.367
R1770 B.n879 B.n878 163.367
R1771 B.n880 B.n879 163.367
R1772 B.n880 B.n21 163.367
R1773 B.n884 B.n21 163.367
R1774 B.n885 B.n884 163.367
R1775 B.n886 B.n885 163.367
R1776 B.n886 B.n19 163.367
R1777 B.n890 B.n19 163.367
R1778 B.n891 B.n890 163.367
R1779 B.n892 B.n891 163.367
R1780 B.n892 B.n17 163.367
R1781 B.n896 B.n17 163.367
R1782 B.n897 B.n896 163.367
R1783 B.n898 B.n897 163.367
R1784 B.n898 B.n15 163.367
R1785 B.n902 B.n15 163.367
R1786 B.n903 B.n902 163.367
R1787 B.n904 B.n903 163.367
R1788 B.n904 B.n13 163.367
R1789 B.n908 B.n13 163.367
R1790 B.n909 B.n908 163.367
R1791 B.n910 B.n909 163.367
R1792 B.n910 B.n11 163.367
R1793 B.n914 B.n11 163.367
R1794 B.n915 B.n914 163.367
R1795 B.n916 B.n915 163.367
R1796 B.n916 B.n9 163.367
R1797 B.n920 B.n9 163.367
R1798 B.n921 B.n920 163.367
R1799 B.n922 B.n921 163.367
R1800 B.n922 B.n7 163.367
R1801 B.n926 B.n7 163.367
R1802 B.n927 B.n926 163.367
R1803 B.n928 B.n927 163.367
R1804 B.n928 B.n5 163.367
R1805 B.n932 B.n5 163.367
R1806 B.n933 B.n932 163.367
R1807 B.n934 B.n933 163.367
R1808 B.n934 B.n3 163.367
R1809 B.n938 B.n3 163.367
R1810 B.n939 B.n938 163.367
R1811 B.n240 B.n2 163.367
R1812 B.n240 B.n239 163.367
R1813 B.n244 B.n239 163.367
R1814 B.n245 B.n244 163.367
R1815 B.n246 B.n245 163.367
R1816 B.n246 B.n237 163.367
R1817 B.n250 B.n237 163.367
R1818 B.n251 B.n250 163.367
R1819 B.n252 B.n251 163.367
R1820 B.n252 B.n235 163.367
R1821 B.n256 B.n235 163.367
R1822 B.n257 B.n256 163.367
R1823 B.n258 B.n257 163.367
R1824 B.n258 B.n233 163.367
R1825 B.n262 B.n233 163.367
R1826 B.n263 B.n262 163.367
R1827 B.n264 B.n263 163.367
R1828 B.n264 B.n231 163.367
R1829 B.n268 B.n231 163.367
R1830 B.n269 B.n268 163.367
R1831 B.n270 B.n269 163.367
R1832 B.n270 B.n229 163.367
R1833 B.n274 B.n229 163.367
R1834 B.n275 B.n274 163.367
R1835 B.n276 B.n275 163.367
R1836 B.n276 B.n227 163.367
R1837 B.n280 B.n227 163.367
R1838 B.n281 B.n280 163.367
R1839 B.n282 B.n281 163.367
R1840 B.n282 B.n225 163.367
R1841 B.n286 B.n225 163.367
R1842 B.n287 B.n286 163.367
R1843 B.n288 B.n287 163.367
R1844 B.n288 B.n223 163.367
R1845 B.n292 B.n223 163.367
R1846 B.n293 B.n292 163.367
R1847 B.n294 B.n293 163.367
R1848 B.n294 B.n221 163.367
R1849 B.n298 B.n221 163.367
R1850 B.n299 B.n298 163.367
R1851 B.n300 B.n299 163.367
R1852 B.n300 B.n219 163.367
R1853 B.n304 B.n219 163.367
R1854 B.n305 B.n304 163.367
R1855 B.n306 B.n305 163.367
R1856 B.n306 B.n217 163.367
R1857 B.n310 B.n217 163.367
R1858 B.n311 B.n310 163.367
R1859 B.n312 B.n311 163.367
R1860 B.n312 B.n215 163.367
R1861 B.n316 B.n215 163.367
R1862 B.n317 B.n316 163.367
R1863 B.n318 B.n317 163.367
R1864 B.n318 B.n213 163.367
R1865 B.n322 B.n213 163.367
R1866 B.n323 B.n322 163.367
R1867 B.n324 B.n323 163.367
R1868 B.n324 B.n211 163.367
R1869 B.n328 B.n211 163.367
R1870 B.n329 B.n328 163.367
R1871 B.n330 B.n329 163.367
R1872 B.n330 B.n209 163.367
R1873 B.n334 B.n209 163.367
R1874 B.n335 B.n334 163.367
R1875 B.n336 B.n335 163.367
R1876 B.n336 B.n207 163.367
R1877 B.n340 B.n207 163.367
R1878 B.n341 B.n340 163.367
R1879 B.n342 B.n341 163.367
R1880 B.n342 B.n205 163.367
R1881 B.n346 B.n205 163.367
R1882 B.n347 B.n346 163.367
R1883 B.n348 B.n347 163.367
R1884 B.n348 B.n203 163.367
R1885 B.n352 B.n203 163.367
R1886 B.n353 B.n352 163.367
R1887 B.n354 B.n353 163.367
R1888 B.n354 B.n201 163.367
R1889 B.n358 B.n201 163.367
R1890 B.n359 B.n358 163.367
R1891 B.n185 B.n184 80.8732
R1892 B.n419 B.n418 80.8732
R1893 B.n65 B.n64 80.8732
R1894 B.n59 B.n58 80.8732
R1895 B.n405 B.n185 59.5399
R1896 B.n420 B.n419 59.5399
R1897 B.n66 B.n65 59.5399
R1898 B.n773 B.n59 59.5399
R1899 B.n817 B.n42 34.4981
R1900 B.n714 B.n713 34.4981
R1901 B.n468 B.n467 34.4981
R1902 B.n361 B.n200 34.4981
R1903 B B.n941 18.0485
R1904 B.n821 B.n42 10.6151
R1905 B.n822 B.n821 10.6151
R1906 B.n823 B.n822 10.6151
R1907 B.n823 B.n40 10.6151
R1908 B.n827 B.n40 10.6151
R1909 B.n828 B.n827 10.6151
R1910 B.n829 B.n828 10.6151
R1911 B.n829 B.n38 10.6151
R1912 B.n833 B.n38 10.6151
R1913 B.n834 B.n833 10.6151
R1914 B.n835 B.n834 10.6151
R1915 B.n835 B.n36 10.6151
R1916 B.n839 B.n36 10.6151
R1917 B.n840 B.n839 10.6151
R1918 B.n841 B.n840 10.6151
R1919 B.n841 B.n34 10.6151
R1920 B.n845 B.n34 10.6151
R1921 B.n846 B.n845 10.6151
R1922 B.n847 B.n846 10.6151
R1923 B.n847 B.n32 10.6151
R1924 B.n851 B.n32 10.6151
R1925 B.n852 B.n851 10.6151
R1926 B.n853 B.n852 10.6151
R1927 B.n853 B.n30 10.6151
R1928 B.n857 B.n30 10.6151
R1929 B.n858 B.n857 10.6151
R1930 B.n859 B.n858 10.6151
R1931 B.n859 B.n28 10.6151
R1932 B.n863 B.n28 10.6151
R1933 B.n864 B.n863 10.6151
R1934 B.n865 B.n864 10.6151
R1935 B.n865 B.n26 10.6151
R1936 B.n869 B.n26 10.6151
R1937 B.n870 B.n869 10.6151
R1938 B.n871 B.n870 10.6151
R1939 B.n871 B.n24 10.6151
R1940 B.n875 B.n24 10.6151
R1941 B.n876 B.n875 10.6151
R1942 B.n877 B.n876 10.6151
R1943 B.n877 B.n22 10.6151
R1944 B.n881 B.n22 10.6151
R1945 B.n882 B.n881 10.6151
R1946 B.n883 B.n882 10.6151
R1947 B.n883 B.n20 10.6151
R1948 B.n887 B.n20 10.6151
R1949 B.n888 B.n887 10.6151
R1950 B.n889 B.n888 10.6151
R1951 B.n889 B.n18 10.6151
R1952 B.n893 B.n18 10.6151
R1953 B.n894 B.n893 10.6151
R1954 B.n895 B.n894 10.6151
R1955 B.n895 B.n16 10.6151
R1956 B.n899 B.n16 10.6151
R1957 B.n900 B.n899 10.6151
R1958 B.n901 B.n900 10.6151
R1959 B.n901 B.n14 10.6151
R1960 B.n905 B.n14 10.6151
R1961 B.n906 B.n905 10.6151
R1962 B.n907 B.n906 10.6151
R1963 B.n907 B.n12 10.6151
R1964 B.n911 B.n12 10.6151
R1965 B.n912 B.n911 10.6151
R1966 B.n913 B.n912 10.6151
R1967 B.n913 B.n10 10.6151
R1968 B.n917 B.n10 10.6151
R1969 B.n918 B.n917 10.6151
R1970 B.n919 B.n918 10.6151
R1971 B.n919 B.n8 10.6151
R1972 B.n923 B.n8 10.6151
R1973 B.n924 B.n923 10.6151
R1974 B.n925 B.n924 10.6151
R1975 B.n925 B.n6 10.6151
R1976 B.n929 B.n6 10.6151
R1977 B.n930 B.n929 10.6151
R1978 B.n931 B.n930 10.6151
R1979 B.n931 B.n4 10.6151
R1980 B.n935 B.n4 10.6151
R1981 B.n936 B.n935 10.6151
R1982 B.n937 B.n936 10.6151
R1983 B.n937 B.n0 10.6151
R1984 B.n817 B.n816 10.6151
R1985 B.n816 B.n815 10.6151
R1986 B.n815 B.n44 10.6151
R1987 B.n811 B.n44 10.6151
R1988 B.n811 B.n810 10.6151
R1989 B.n810 B.n809 10.6151
R1990 B.n809 B.n46 10.6151
R1991 B.n805 B.n46 10.6151
R1992 B.n805 B.n804 10.6151
R1993 B.n804 B.n803 10.6151
R1994 B.n803 B.n48 10.6151
R1995 B.n799 B.n48 10.6151
R1996 B.n799 B.n798 10.6151
R1997 B.n798 B.n797 10.6151
R1998 B.n797 B.n50 10.6151
R1999 B.n793 B.n50 10.6151
R2000 B.n793 B.n792 10.6151
R2001 B.n792 B.n791 10.6151
R2002 B.n791 B.n52 10.6151
R2003 B.n787 B.n52 10.6151
R2004 B.n787 B.n786 10.6151
R2005 B.n786 B.n785 10.6151
R2006 B.n785 B.n54 10.6151
R2007 B.n781 B.n54 10.6151
R2008 B.n781 B.n780 10.6151
R2009 B.n780 B.n779 10.6151
R2010 B.n779 B.n56 10.6151
R2011 B.n775 B.n56 10.6151
R2012 B.n775 B.n774 10.6151
R2013 B.n772 B.n60 10.6151
R2014 B.n768 B.n60 10.6151
R2015 B.n768 B.n767 10.6151
R2016 B.n767 B.n766 10.6151
R2017 B.n766 B.n62 10.6151
R2018 B.n762 B.n62 10.6151
R2019 B.n762 B.n761 10.6151
R2020 B.n761 B.n760 10.6151
R2021 B.n757 B.n756 10.6151
R2022 B.n756 B.n755 10.6151
R2023 B.n755 B.n68 10.6151
R2024 B.n751 B.n68 10.6151
R2025 B.n751 B.n750 10.6151
R2026 B.n750 B.n749 10.6151
R2027 B.n749 B.n70 10.6151
R2028 B.n745 B.n70 10.6151
R2029 B.n745 B.n744 10.6151
R2030 B.n744 B.n743 10.6151
R2031 B.n743 B.n72 10.6151
R2032 B.n739 B.n72 10.6151
R2033 B.n739 B.n738 10.6151
R2034 B.n738 B.n737 10.6151
R2035 B.n737 B.n74 10.6151
R2036 B.n733 B.n74 10.6151
R2037 B.n733 B.n732 10.6151
R2038 B.n732 B.n731 10.6151
R2039 B.n731 B.n76 10.6151
R2040 B.n727 B.n76 10.6151
R2041 B.n727 B.n726 10.6151
R2042 B.n726 B.n725 10.6151
R2043 B.n725 B.n78 10.6151
R2044 B.n721 B.n78 10.6151
R2045 B.n721 B.n720 10.6151
R2046 B.n720 B.n719 10.6151
R2047 B.n719 B.n80 10.6151
R2048 B.n715 B.n80 10.6151
R2049 B.n715 B.n714 10.6151
R2050 B.n713 B.n82 10.6151
R2051 B.n709 B.n82 10.6151
R2052 B.n709 B.n708 10.6151
R2053 B.n708 B.n707 10.6151
R2054 B.n707 B.n84 10.6151
R2055 B.n703 B.n84 10.6151
R2056 B.n703 B.n702 10.6151
R2057 B.n702 B.n701 10.6151
R2058 B.n701 B.n86 10.6151
R2059 B.n697 B.n86 10.6151
R2060 B.n697 B.n696 10.6151
R2061 B.n696 B.n695 10.6151
R2062 B.n695 B.n88 10.6151
R2063 B.n691 B.n88 10.6151
R2064 B.n691 B.n690 10.6151
R2065 B.n690 B.n689 10.6151
R2066 B.n689 B.n90 10.6151
R2067 B.n685 B.n90 10.6151
R2068 B.n685 B.n684 10.6151
R2069 B.n684 B.n683 10.6151
R2070 B.n683 B.n92 10.6151
R2071 B.n679 B.n92 10.6151
R2072 B.n679 B.n678 10.6151
R2073 B.n678 B.n677 10.6151
R2074 B.n677 B.n94 10.6151
R2075 B.n673 B.n94 10.6151
R2076 B.n673 B.n672 10.6151
R2077 B.n672 B.n671 10.6151
R2078 B.n671 B.n96 10.6151
R2079 B.n667 B.n96 10.6151
R2080 B.n667 B.n666 10.6151
R2081 B.n666 B.n665 10.6151
R2082 B.n665 B.n98 10.6151
R2083 B.n661 B.n98 10.6151
R2084 B.n661 B.n660 10.6151
R2085 B.n660 B.n659 10.6151
R2086 B.n659 B.n100 10.6151
R2087 B.n655 B.n100 10.6151
R2088 B.n655 B.n654 10.6151
R2089 B.n654 B.n653 10.6151
R2090 B.n653 B.n102 10.6151
R2091 B.n649 B.n102 10.6151
R2092 B.n649 B.n648 10.6151
R2093 B.n648 B.n647 10.6151
R2094 B.n647 B.n104 10.6151
R2095 B.n643 B.n104 10.6151
R2096 B.n643 B.n642 10.6151
R2097 B.n642 B.n641 10.6151
R2098 B.n641 B.n106 10.6151
R2099 B.n637 B.n106 10.6151
R2100 B.n637 B.n636 10.6151
R2101 B.n636 B.n635 10.6151
R2102 B.n635 B.n108 10.6151
R2103 B.n631 B.n108 10.6151
R2104 B.n631 B.n630 10.6151
R2105 B.n630 B.n629 10.6151
R2106 B.n629 B.n110 10.6151
R2107 B.n625 B.n110 10.6151
R2108 B.n625 B.n624 10.6151
R2109 B.n624 B.n623 10.6151
R2110 B.n623 B.n112 10.6151
R2111 B.n619 B.n112 10.6151
R2112 B.n619 B.n618 10.6151
R2113 B.n618 B.n617 10.6151
R2114 B.n617 B.n114 10.6151
R2115 B.n613 B.n114 10.6151
R2116 B.n613 B.n612 10.6151
R2117 B.n612 B.n611 10.6151
R2118 B.n611 B.n116 10.6151
R2119 B.n607 B.n116 10.6151
R2120 B.n607 B.n606 10.6151
R2121 B.n606 B.n605 10.6151
R2122 B.n605 B.n118 10.6151
R2123 B.n601 B.n118 10.6151
R2124 B.n601 B.n600 10.6151
R2125 B.n600 B.n599 10.6151
R2126 B.n599 B.n120 10.6151
R2127 B.n595 B.n120 10.6151
R2128 B.n595 B.n594 10.6151
R2129 B.n594 B.n593 10.6151
R2130 B.n593 B.n122 10.6151
R2131 B.n589 B.n122 10.6151
R2132 B.n589 B.n588 10.6151
R2133 B.n588 B.n587 10.6151
R2134 B.n587 B.n124 10.6151
R2135 B.n583 B.n124 10.6151
R2136 B.n583 B.n582 10.6151
R2137 B.n582 B.n581 10.6151
R2138 B.n581 B.n126 10.6151
R2139 B.n577 B.n126 10.6151
R2140 B.n577 B.n576 10.6151
R2141 B.n576 B.n575 10.6151
R2142 B.n575 B.n128 10.6151
R2143 B.n571 B.n128 10.6151
R2144 B.n571 B.n570 10.6151
R2145 B.n570 B.n569 10.6151
R2146 B.n569 B.n130 10.6151
R2147 B.n565 B.n130 10.6151
R2148 B.n565 B.n564 10.6151
R2149 B.n564 B.n563 10.6151
R2150 B.n563 B.n132 10.6151
R2151 B.n559 B.n132 10.6151
R2152 B.n559 B.n558 10.6151
R2153 B.n558 B.n557 10.6151
R2154 B.n557 B.n134 10.6151
R2155 B.n553 B.n134 10.6151
R2156 B.n553 B.n552 10.6151
R2157 B.n552 B.n551 10.6151
R2158 B.n551 B.n136 10.6151
R2159 B.n547 B.n136 10.6151
R2160 B.n547 B.n546 10.6151
R2161 B.n546 B.n545 10.6151
R2162 B.n545 B.n138 10.6151
R2163 B.n541 B.n138 10.6151
R2164 B.n541 B.n540 10.6151
R2165 B.n540 B.n539 10.6151
R2166 B.n539 B.n140 10.6151
R2167 B.n535 B.n140 10.6151
R2168 B.n535 B.n534 10.6151
R2169 B.n534 B.n533 10.6151
R2170 B.n533 B.n142 10.6151
R2171 B.n529 B.n142 10.6151
R2172 B.n529 B.n528 10.6151
R2173 B.n528 B.n527 10.6151
R2174 B.n527 B.n144 10.6151
R2175 B.n523 B.n144 10.6151
R2176 B.n523 B.n522 10.6151
R2177 B.n522 B.n521 10.6151
R2178 B.n521 B.n146 10.6151
R2179 B.n517 B.n146 10.6151
R2180 B.n517 B.n516 10.6151
R2181 B.n516 B.n515 10.6151
R2182 B.n515 B.n148 10.6151
R2183 B.n511 B.n148 10.6151
R2184 B.n511 B.n510 10.6151
R2185 B.n510 B.n509 10.6151
R2186 B.n509 B.n150 10.6151
R2187 B.n505 B.n150 10.6151
R2188 B.n505 B.n504 10.6151
R2189 B.n504 B.n503 10.6151
R2190 B.n503 B.n152 10.6151
R2191 B.n499 B.n152 10.6151
R2192 B.n499 B.n498 10.6151
R2193 B.n498 B.n497 10.6151
R2194 B.n497 B.n154 10.6151
R2195 B.n493 B.n154 10.6151
R2196 B.n493 B.n492 10.6151
R2197 B.n492 B.n491 10.6151
R2198 B.n491 B.n156 10.6151
R2199 B.n487 B.n156 10.6151
R2200 B.n487 B.n486 10.6151
R2201 B.n486 B.n485 10.6151
R2202 B.n485 B.n158 10.6151
R2203 B.n481 B.n158 10.6151
R2204 B.n481 B.n480 10.6151
R2205 B.n480 B.n479 10.6151
R2206 B.n479 B.n160 10.6151
R2207 B.n475 B.n160 10.6151
R2208 B.n475 B.n474 10.6151
R2209 B.n474 B.n473 10.6151
R2210 B.n473 B.n162 10.6151
R2211 B.n469 B.n162 10.6151
R2212 B.n469 B.n468 10.6151
R2213 B.n241 B.n1 10.6151
R2214 B.n242 B.n241 10.6151
R2215 B.n243 B.n242 10.6151
R2216 B.n243 B.n238 10.6151
R2217 B.n247 B.n238 10.6151
R2218 B.n248 B.n247 10.6151
R2219 B.n249 B.n248 10.6151
R2220 B.n249 B.n236 10.6151
R2221 B.n253 B.n236 10.6151
R2222 B.n254 B.n253 10.6151
R2223 B.n255 B.n254 10.6151
R2224 B.n255 B.n234 10.6151
R2225 B.n259 B.n234 10.6151
R2226 B.n260 B.n259 10.6151
R2227 B.n261 B.n260 10.6151
R2228 B.n261 B.n232 10.6151
R2229 B.n265 B.n232 10.6151
R2230 B.n266 B.n265 10.6151
R2231 B.n267 B.n266 10.6151
R2232 B.n267 B.n230 10.6151
R2233 B.n271 B.n230 10.6151
R2234 B.n272 B.n271 10.6151
R2235 B.n273 B.n272 10.6151
R2236 B.n273 B.n228 10.6151
R2237 B.n277 B.n228 10.6151
R2238 B.n278 B.n277 10.6151
R2239 B.n279 B.n278 10.6151
R2240 B.n279 B.n226 10.6151
R2241 B.n283 B.n226 10.6151
R2242 B.n284 B.n283 10.6151
R2243 B.n285 B.n284 10.6151
R2244 B.n285 B.n224 10.6151
R2245 B.n289 B.n224 10.6151
R2246 B.n290 B.n289 10.6151
R2247 B.n291 B.n290 10.6151
R2248 B.n291 B.n222 10.6151
R2249 B.n295 B.n222 10.6151
R2250 B.n296 B.n295 10.6151
R2251 B.n297 B.n296 10.6151
R2252 B.n297 B.n220 10.6151
R2253 B.n301 B.n220 10.6151
R2254 B.n302 B.n301 10.6151
R2255 B.n303 B.n302 10.6151
R2256 B.n303 B.n218 10.6151
R2257 B.n307 B.n218 10.6151
R2258 B.n308 B.n307 10.6151
R2259 B.n309 B.n308 10.6151
R2260 B.n309 B.n216 10.6151
R2261 B.n313 B.n216 10.6151
R2262 B.n314 B.n313 10.6151
R2263 B.n315 B.n314 10.6151
R2264 B.n315 B.n214 10.6151
R2265 B.n319 B.n214 10.6151
R2266 B.n320 B.n319 10.6151
R2267 B.n321 B.n320 10.6151
R2268 B.n321 B.n212 10.6151
R2269 B.n325 B.n212 10.6151
R2270 B.n326 B.n325 10.6151
R2271 B.n327 B.n326 10.6151
R2272 B.n327 B.n210 10.6151
R2273 B.n331 B.n210 10.6151
R2274 B.n332 B.n331 10.6151
R2275 B.n333 B.n332 10.6151
R2276 B.n333 B.n208 10.6151
R2277 B.n337 B.n208 10.6151
R2278 B.n338 B.n337 10.6151
R2279 B.n339 B.n338 10.6151
R2280 B.n339 B.n206 10.6151
R2281 B.n343 B.n206 10.6151
R2282 B.n344 B.n343 10.6151
R2283 B.n345 B.n344 10.6151
R2284 B.n345 B.n204 10.6151
R2285 B.n349 B.n204 10.6151
R2286 B.n350 B.n349 10.6151
R2287 B.n351 B.n350 10.6151
R2288 B.n351 B.n202 10.6151
R2289 B.n355 B.n202 10.6151
R2290 B.n356 B.n355 10.6151
R2291 B.n357 B.n356 10.6151
R2292 B.n357 B.n200 10.6151
R2293 B.n362 B.n361 10.6151
R2294 B.n363 B.n362 10.6151
R2295 B.n363 B.n198 10.6151
R2296 B.n367 B.n198 10.6151
R2297 B.n368 B.n367 10.6151
R2298 B.n369 B.n368 10.6151
R2299 B.n369 B.n196 10.6151
R2300 B.n373 B.n196 10.6151
R2301 B.n374 B.n373 10.6151
R2302 B.n375 B.n374 10.6151
R2303 B.n375 B.n194 10.6151
R2304 B.n379 B.n194 10.6151
R2305 B.n380 B.n379 10.6151
R2306 B.n381 B.n380 10.6151
R2307 B.n381 B.n192 10.6151
R2308 B.n385 B.n192 10.6151
R2309 B.n386 B.n385 10.6151
R2310 B.n387 B.n386 10.6151
R2311 B.n387 B.n190 10.6151
R2312 B.n391 B.n190 10.6151
R2313 B.n392 B.n391 10.6151
R2314 B.n393 B.n392 10.6151
R2315 B.n393 B.n188 10.6151
R2316 B.n397 B.n188 10.6151
R2317 B.n398 B.n397 10.6151
R2318 B.n399 B.n398 10.6151
R2319 B.n399 B.n186 10.6151
R2320 B.n403 B.n186 10.6151
R2321 B.n404 B.n403 10.6151
R2322 B.n406 B.n182 10.6151
R2323 B.n410 B.n182 10.6151
R2324 B.n411 B.n410 10.6151
R2325 B.n412 B.n411 10.6151
R2326 B.n412 B.n180 10.6151
R2327 B.n416 B.n180 10.6151
R2328 B.n417 B.n416 10.6151
R2329 B.n421 B.n417 10.6151
R2330 B.n425 B.n178 10.6151
R2331 B.n426 B.n425 10.6151
R2332 B.n427 B.n426 10.6151
R2333 B.n427 B.n176 10.6151
R2334 B.n431 B.n176 10.6151
R2335 B.n432 B.n431 10.6151
R2336 B.n433 B.n432 10.6151
R2337 B.n433 B.n174 10.6151
R2338 B.n437 B.n174 10.6151
R2339 B.n438 B.n437 10.6151
R2340 B.n439 B.n438 10.6151
R2341 B.n439 B.n172 10.6151
R2342 B.n443 B.n172 10.6151
R2343 B.n444 B.n443 10.6151
R2344 B.n445 B.n444 10.6151
R2345 B.n445 B.n170 10.6151
R2346 B.n449 B.n170 10.6151
R2347 B.n450 B.n449 10.6151
R2348 B.n451 B.n450 10.6151
R2349 B.n451 B.n168 10.6151
R2350 B.n455 B.n168 10.6151
R2351 B.n456 B.n455 10.6151
R2352 B.n457 B.n456 10.6151
R2353 B.n457 B.n166 10.6151
R2354 B.n461 B.n166 10.6151
R2355 B.n462 B.n461 10.6151
R2356 B.n463 B.n462 10.6151
R2357 B.n463 B.n164 10.6151
R2358 B.n467 B.n164 10.6151
R2359 B.n941 B.n0 8.11757
R2360 B.n941 B.n1 8.11757
R2361 B.n773 B.n772 6.5566
R2362 B.n760 B.n66 6.5566
R2363 B.n406 B.n405 6.5566
R2364 B.n421 B.n420 6.5566
R2365 B.n774 B.n773 4.05904
R2366 B.n757 B.n66 4.05904
R2367 B.n405 B.n404 4.05904
R2368 B.n420 B.n178 4.05904
C0 w_n5974_n2558# VP 13.8597f
C1 w_n5974_n2558# VDD1 2.97927f
C2 w_n5974_n2558# VN 13.0781f
C3 w_n5974_n2558# VTAIL 2.84104f
C4 VP VDD1 8.31531f
C5 VDD2 w_n5974_n2558# 3.18726f
C6 VP VN 9.47596f
C7 VN VDD1 0.156075f
C8 VP VTAIL 9.11629f
C9 VTAIL VDD1 9.47981f
C10 w_n5974_n2558# B 11.495901f
C11 VDD2 VP 0.741078f
C12 VN VTAIL 9.10173f
C13 VDD2 VDD1 2.98117f
C14 VDD2 VN 7.733439f
C15 VDD2 VTAIL 9.54067f
C16 B VP 2.8724f
C17 B VDD1 2.63399f
C18 B VN 1.55123f
C19 B VTAIL 3.22623f
C20 VDD2 B 2.8002f
C21 VDD2 VSUBS 2.59836f
C22 VDD1 VSUBS 2.405853f
C23 VTAIL VSUBS 1.480338f
C24 VN VSUBS 9.771741f
C25 VP VSUBS 5.674374f
C26 B VSUBS 6.562293f
C27 w_n5974_n2558# VSUBS 0.189615p
C28 B.n0 VSUBS 0.009123f
C29 B.n1 VSUBS 0.009123f
C30 B.n2 VSUBS 0.013492f
C31 B.n3 VSUBS 0.010339f
C32 B.n4 VSUBS 0.010339f
C33 B.n5 VSUBS 0.010339f
C34 B.n6 VSUBS 0.010339f
C35 B.n7 VSUBS 0.010339f
C36 B.n8 VSUBS 0.010339f
C37 B.n9 VSUBS 0.010339f
C38 B.n10 VSUBS 0.010339f
C39 B.n11 VSUBS 0.010339f
C40 B.n12 VSUBS 0.010339f
C41 B.n13 VSUBS 0.010339f
C42 B.n14 VSUBS 0.010339f
C43 B.n15 VSUBS 0.010339f
C44 B.n16 VSUBS 0.010339f
C45 B.n17 VSUBS 0.010339f
C46 B.n18 VSUBS 0.010339f
C47 B.n19 VSUBS 0.010339f
C48 B.n20 VSUBS 0.010339f
C49 B.n21 VSUBS 0.010339f
C50 B.n22 VSUBS 0.010339f
C51 B.n23 VSUBS 0.010339f
C52 B.n24 VSUBS 0.010339f
C53 B.n25 VSUBS 0.010339f
C54 B.n26 VSUBS 0.010339f
C55 B.n27 VSUBS 0.010339f
C56 B.n28 VSUBS 0.010339f
C57 B.n29 VSUBS 0.010339f
C58 B.n30 VSUBS 0.010339f
C59 B.n31 VSUBS 0.010339f
C60 B.n32 VSUBS 0.010339f
C61 B.n33 VSUBS 0.010339f
C62 B.n34 VSUBS 0.010339f
C63 B.n35 VSUBS 0.010339f
C64 B.n36 VSUBS 0.010339f
C65 B.n37 VSUBS 0.010339f
C66 B.n38 VSUBS 0.010339f
C67 B.n39 VSUBS 0.010339f
C68 B.n40 VSUBS 0.010339f
C69 B.n41 VSUBS 0.010339f
C70 B.n42 VSUBS 0.02434f
C71 B.n43 VSUBS 0.010339f
C72 B.n44 VSUBS 0.010339f
C73 B.n45 VSUBS 0.010339f
C74 B.n46 VSUBS 0.010339f
C75 B.n47 VSUBS 0.010339f
C76 B.n48 VSUBS 0.010339f
C77 B.n49 VSUBS 0.010339f
C78 B.n50 VSUBS 0.010339f
C79 B.n51 VSUBS 0.010339f
C80 B.n52 VSUBS 0.010339f
C81 B.n53 VSUBS 0.010339f
C82 B.n54 VSUBS 0.010339f
C83 B.n55 VSUBS 0.010339f
C84 B.n56 VSUBS 0.010339f
C85 B.n57 VSUBS 0.010339f
C86 B.t10 VSUBS 0.185479f
C87 B.t11 VSUBS 0.243402f
C88 B.t9 VSUBS 2.14522f
C89 B.n58 VSUBS 0.394957f
C90 B.n59 VSUBS 0.289488f
C91 B.n60 VSUBS 0.010339f
C92 B.n61 VSUBS 0.010339f
C93 B.n62 VSUBS 0.010339f
C94 B.n63 VSUBS 0.010339f
C95 B.t4 VSUBS 0.185482f
C96 B.t5 VSUBS 0.243405f
C97 B.t3 VSUBS 2.14522f
C98 B.n64 VSUBS 0.394955f
C99 B.n65 VSUBS 0.289485f
C100 B.n66 VSUBS 0.023955f
C101 B.n67 VSUBS 0.010339f
C102 B.n68 VSUBS 0.010339f
C103 B.n69 VSUBS 0.010339f
C104 B.n70 VSUBS 0.010339f
C105 B.n71 VSUBS 0.010339f
C106 B.n72 VSUBS 0.010339f
C107 B.n73 VSUBS 0.010339f
C108 B.n74 VSUBS 0.010339f
C109 B.n75 VSUBS 0.010339f
C110 B.n76 VSUBS 0.010339f
C111 B.n77 VSUBS 0.010339f
C112 B.n78 VSUBS 0.010339f
C113 B.n79 VSUBS 0.010339f
C114 B.n80 VSUBS 0.010339f
C115 B.n81 VSUBS 0.025835f
C116 B.n82 VSUBS 0.010339f
C117 B.n83 VSUBS 0.010339f
C118 B.n84 VSUBS 0.010339f
C119 B.n85 VSUBS 0.010339f
C120 B.n86 VSUBS 0.010339f
C121 B.n87 VSUBS 0.010339f
C122 B.n88 VSUBS 0.010339f
C123 B.n89 VSUBS 0.010339f
C124 B.n90 VSUBS 0.010339f
C125 B.n91 VSUBS 0.010339f
C126 B.n92 VSUBS 0.010339f
C127 B.n93 VSUBS 0.010339f
C128 B.n94 VSUBS 0.010339f
C129 B.n95 VSUBS 0.010339f
C130 B.n96 VSUBS 0.010339f
C131 B.n97 VSUBS 0.010339f
C132 B.n98 VSUBS 0.010339f
C133 B.n99 VSUBS 0.010339f
C134 B.n100 VSUBS 0.010339f
C135 B.n101 VSUBS 0.010339f
C136 B.n102 VSUBS 0.010339f
C137 B.n103 VSUBS 0.010339f
C138 B.n104 VSUBS 0.010339f
C139 B.n105 VSUBS 0.010339f
C140 B.n106 VSUBS 0.010339f
C141 B.n107 VSUBS 0.010339f
C142 B.n108 VSUBS 0.010339f
C143 B.n109 VSUBS 0.010339f
C144 B.n110 VSUBS 0.010339f
C145 B.n111 VSUBS 0.010339f
C146 B.n112 VSUBS 0.010339f
C147 B.n113 VSUBS 0.010339f
C148 B.n114 VSUBS 0.010339f
C149 B.n115 VSUBS 0.010339f
C150 B.n116 VSUBS 0.010339f
C151 B.n117 VSUBS 0.010339f
C152 B.n118 VSUBS 0.010339f
C153 B.n119 VSUBS 0.010339f
C154 B.n120 VSUBS 0.010339f
C155 B.n121 VSUBS 0.010339f
C156 B.n122 VSUBS 0.010339f
C157 B.n123 VSUBS 0.010339f
C158 B.n124 VSUBS 0.010339f
C159 B.n125 VSUBS 0.010339f
C160 B.n126 VSUBS 0.010339f
C161 B.n127 VSUBS 0.010339f
C162 B.n128 VSUBS 0.010339f
C163 B.n129 VSUBS 0.010339f
C164 B.n130 VSUBS 0.010339f
C165 B.n131 VSUBS 0.010339f
C166 B.n132 VSUBS 0.010339f
C167 B.n133 VSUBS 0.010339f
C168 B.n134 VSUBS 0.010339f
C169 B.n135 VSUBS 0.010339f
C170 B.n136 VSUBS 0.010339f
C171 B.n137 VSUBS 0.010339f
C172 B.n138 VSUBS 0.010339f
C173 B.n139 VSUBS 0.010339f
C174 B.n140 VSUBS 0.010339f
C175 B.n141 VSUBS 0.010339f
C176 B.n142 VSUBS 0.010339f
C177 B.n143 VSUBS 0.010339f
C178 B.n144 VSUBS 0.010339f
C179 B.n145 VSUBS 0.010339f
C180 B.n146 VSUBS 0.010339f
C181 B.n147 VSUBS 0.010339f
C182 B.n148 VSUBS 0.010339f
C183 B.n149 VSUBS 0.010339f
C184 B.n150 VSUBS 0.010339f
C185 B.n151 VSUBS 0.010339f
C186 B.n152 VSUBS 0.010339f
C187 B.n153 VSUBS 0.010339f
C188 B.n154 VSUBS 0.010339f
C189 B.n155 VSUBS 0.010339f
C190 B.n156 VSUBS 0.010339f
C191 B.n157 VSUBS 0.010339f
C192 B.n158 VSUBS 0.010339f
C193 B.n159 VSUBS 0.010339f
C194 B.n160 VSUBS 0.010339f
C195 B.n161 VSUBS 0.010339f
C196 B.n162 VSUBS 0.010339f
C197 B.n163 VSUBS 0.02434f
C198 B.n164 VSUBS 0.010339f
C199 B.n165 VSUBS 0.010339f
C200 B.n166 VSUBS 0.010339f
C201 B.n167 VSUBS 0.010339f
C202 B.n168 VSUBS 0.010339f
C203 B.n169 VSUBS 0.010339f
C204 B.n170 VSUBS 0.010339f
C205 B.n171 VSUBS 0.010339f
C206 B.n172 VSUBS 0.010339f
C207 B.n173 VSUBS 0.010339f
C208 B.n174 VSUBS 0.010339f
C209 B.n175 VSUBS 0.010339f
C210 B.n176 VSUBS 0.010339f
C211 B.n177 VSUBS 0.010339f
C212 B.n178 VSUBS 0.007146f
C213 B.n179 VSUBS 0.010339f
C214 B.n180 VSUBS 0.010339f
C215 B.n181 VSUBS 0.010339f
C216 B.n182 VSUBS 0.010339f
C217 B.n183 VSUBS 0.010339f
C218 B.t2 VSUBS 0.185479f
C219 B.t1 VSUBS 0.243402f
C220 B.t0 VSUBS 2.14522f
C221 B.n184 VSUBS 0.394957f
C222 B.n185 VSUBS 0.289488f
C223 B.n186 VSUBS 0.010339f
C224 B.n187 VSUBS 0.010339f
C225 B.n188 VSUBS 0.010339f
C226 B.n189 VSUBS 0.010339f
C227 B.n190 VSUBS 0.010339f
C228 B.n191 VSUBS 0.010339f
C229 B.n192 VSUBS 0.010339f
C230 B.n193 VSUBS 0.010339f
C231 B.n194 VSUBS 0.010339f
C232 B.n195 VSUBS 0.010339f
C233 B.n196 VSUBS 0.010339f
C234 B.n197 VSUBS 0.010339f
C235 B.n198 VSUBS 0.010339f
C236 B.n199 VSUBS 0.010339f
C237 B.n200 VSUBS 0.02434f
C238 B.n201 VSUBS 0.010339f
C239 B.n202 VSUBS 0.010339f
C240 B.n203 VSUBS 0.010339f
C241 B.n204 VSUBS 0.010339f
C242 B.n205 VSUBS 0.010339f
C243 B.n206 VSUBS 0.010339f
C244 B.n207 VSUBS 0.010339f
C245 B.n208 VSUBS 0.010339f
C246 B.n209 VSUBS 0.010339f
C247 B.n210 VSUBS 0.010339f
C248 B.n211 VSUBS 0.010339f
C249 B.n212 VSUBS 0.010339f
C250 B.n213 VSUBS 0.010339f
C251 B.n214 VSUBS 0.010339f
C252 B.n215 VSUBS 0.010339f
C253 B.n216 VSUBS 0.010339f
C254 B.n217 VSUBS 0.010339f
C255 B.n218 VSUBS 0.010339f
C256 B.n219 VSUBS 0.010339f
C257 B.n220 VSUBS 0.010339f
C258 B.n221 VSUBS 0.010339f
C259 B.n222 VSUBS 0.010339f
C260 B.n223 VSUBS 0.010339f
C261 B.n224 VSUBS 0.010339f
C262 B.n225 VSUBS 0.010339f
C263 B.n226 VSUBS 0.010339f
C264 B.n227 VSUBS 0.010339f
C265 B.n228 VSUBS 0.010339f
C266 B.n229 VSUBS 0.010339f
C267 B.n230 VSUBS 0.010339f
C268 B.n231 VSUBS 0.010339f
C269 B.n232 VSUBS 0.010339f
C270 B.n233 VSUBS 0.010339f
C271 B.n234 VSUBS 0.010339f
C272 B.n235 VSUBS 0.010339f
C273 B.n236 VSUBS 0.010339f
C274 B.n237 VSUBS 0.010339f
C275 B.n238 VSUBS 0.010339f
C276 B.n239 VSUBS 0.010339f
C277 B.n240 VSUBS 0.010339f
C278 B.n241 VSUBS 0.010339f
C279 B.n242 VSUBS 0.010339f
C280 B.n243 VSUBS 0.010339f
C281 B.n244 VSUBS 0.010339f
C282 B.n245 VSUBS 0.010339f
C283 B.n246 VSUBS 0.010339f
C284 B.n247 VSUBS 0.010339f
C285 B.n248 VSUBS 0.010339f
C286 B.n249 VSUBS 0.010339f
C287 B.n250 VSUBS 0.010339f
C288 B.n251 VSUBS 0.010339f
C289 B.n252 VSUBS 0.010339f
C290 B.n253 VSUBS 0.010339f
C291 B.n254 VSUBS 0.010339f
C292 B.n255 VSUBS 0.010339f
C293 B.n256 VSUBS 0.010339f
C294 B.n257 VSUBS 0.010339f
C295 B.n258 VSUBS 0.010339f
C296 B.n259 VSUBS 0.010339f
C297 B.n260 VSUBS 0.010339f
C298 B.n261 VSUBS 0.010339f
C299 B.n262 VSUBS 0.010339f
C300 B.n263 VSUBS 0.010339f
C301 B.n264 VSUBS 0.010339f
C302 B.n265 VSUBS 0.010339f
C303 B.n266 VSUBS 0.010339f
C304 B.n267 VSUBS 0.010339f
C305 B.n268 VSUBS 0.010339f
C306 B.n269 VSUBS 0.010339f
C307 B.n270 VSUBS 0.010339f
C308 B.n271 VSUBS 0.010339f
C309 B.n272 VSUBS 0.010339f
C310 B.n273 VSUBS 0.010339f
C311 B.n274 VSUBS 0.010339f
C312 B.n275 VSUBS 0.010339f
C313 B.n276 VSUBS 0.010339f
C314 B.n277 VSUBS 0.010339f
C315 B.n278 VSUBS 0.010339f
C316 B.n279 VSUBS 0.010339f
C317 B.n280 VSUBS 0.010339f
C318 B.n281 VSUBS 0.010339f
C319 B.n282 VSUBS 0.010339f
C320 B.n283 VSUBS 0.010339f
C321 B.n284 VSUBS 0.010339f
C322 B.n285 VSUBS 0.010339f
C323 B.n286 VSUBS 0.010339f
C324 B.n287 VSUBS 0.010339f
C325 B.n288 VSUBS 0.010339f
C326 B.n289 VSUBS 0.010339f
C327 B.n290 VSUBS 0.010339f
C328 B.n291 VSUBS 0.010339f
C329 B.n292 VSUBS 0.010339f
C330 B.n293 VSUBS 0.010339f
C331 B.n294 VSUBS 0.010339f
C332 B.n295 VSUBS 0.010339f
C333 B.n296 VSUBS 0.010339f
C334 B.n297 VSUBS 0.010339f
C335 B.n298 VSUBS 0.010339f
C336 B.n299 VSUBS 0.010339f
C337 B.n300 VSUBS 0.010339f
C338 B.n301 VSUBS 0.010339f
C339 B.n302 VSUBS 0.010339f
C340 B.n303 VSUBS 0.010339f
C341 B.n304 VSUBS 0.010339f
C342 B.n305 VSUBS 0.010339f
C343 B.n306 VSUBS 0.010339f
C344 B.n307 VSUBS 0.010339f
C345 B.n308 VSUBS 0.010339f
C346 B.n309 VSUBS 0.010339f
C347 B.n310 VSUBS 0.010339f
C348 B.n311 VSUBS 0.010339f
C349 B.n312 VSUBS 0.010339f
C350 B.n313 VSUBS 0.010339f
C351 B.n314 VSUBS 0.010339f
C352 B.n315 VSUBS 0.010339f
C353 B.n316 VSUBS 0.010339f
C354 B.n317 VSUBS 0.010339f
C355 B.n318 VSUBS 0.010339f
C356 B.n319 VSUBS 0.010339f
C357 B.n320 VSUBS 0.010339f
C358 B.n321 VSUBS 0.010339f
C359 B.n322 VSUBS 0.010339f
C360 B.n323 VSUBS 0.010339f
C361 B.n324 VSUBS 0.010339f
C362 B.n325 VSUBS 0.010339f
C363 B.n326 VSUBS 0.010339f
C364 B.n327 VSUBS 0.010339f
C365 B.n328 VSUBS 0.010339f
C366 B.n329 VSUBS 0.010339f
C367 B.n330 VSUBS 0.010339f
C368 B.n331 VSUBS 0.010339f
C369 B.n332 VSUBS 0.010339f
C370 B.n333 VSUBS 0.010339f
C371 B.n334 VSUBS 0.010339f
C372 B.n335 VSUBS 0.010339f
C373 B.n336 VSUBS 0.010339f
C374 B.n337 VSUBS 0.010339f
C375 B.n338 VSUBS 0.010339f
C376 B.n339 VSUBS 0.010339f
C377 B.n340 VSUBS 0.010339f
C378 B.n341 VSUBS 0.010339f
C379 B.n342 VSUBS 0.010339f
C380 B.n343 VSUBS 0.010339f
C381 B.n344 VSUBS 0.010339f
C382 B.n345 VSUBS 0.010339f
C383 B.n346 VSUBS 0.010339f
C384 B.n347 VSUBS 0.010339f
C385 B.n348 VSUBS 0.010339f
C386 B.n349 VSUBS 0.010339f
C387 B.n350 VSUBS 0.010339f
C388 B.n351 VSUBS 0.010339f
C389 B.n352 VSUBS 0.010339f
C390 B.n353 VSUBS 0.010339f
C391 B.n354 VSUBS 0.010339f
C392 B.n355 VSUBS 0.010339f
C393 B.n356 VSUBS 0.010339f
C394 B.n357 VSUBS 0.010339f
C395 B.n358 VSUBS 0.010339f
C396 B.n359 VSUBS 0.02434f
C397 B.n360 VSUBS 0.025835f
C398 B.n361 VSUBS 0.025835f
C399 B.n362 VSUBS 0.010339f
C400 B.n363 VSUBS 0.010339f
C401 B.n364 VSUBS 0.010339f
C402 B.n365 VSUBS 0.010339f
C403 B.n366 VSUBS 0.010339f
C404 B.n367 VSUBS 0.010339f
C405 B.n368 VSUBS 0.010339f
C406 B.n369 VSUBS 0.010339f
C407 B.n370 VSUBS 0.010339f
C408 B.n371 VSUBS 0.010339f
C409 B.n372 VSUBS 0.010339f
C410 B.n373 VSUBS 0.010339f
C411 B.n374 VSUBS 0.010339f
C412 B.n375 VSUBS 0.010339f
C413 B.n376 VSUBS 0.010339f
C414 B.n377 VSUBS 0.010339f
C415 B.n378 VSUBS 0.010339f
C416 B.n379 VSUBS 0.010339f
C417 B.n380 VSUBS 0.010339f
C418 B.n381 VSUBS 0.010339f
C419 B.n382 VSUBS 0.010339f
C420 B.n383 VSUBS 0.010339f
C421 B.n384 VSUBS 0.010339f
C422 B.n385 VSUBS 0.010339f
C423 B.n386 VSUBS 0.010339f
C424 B.n387 VSUBS 0.010339f
C425 B.n388 VSUBS 0.010339f
C426 B.n389 VSUBS 0.010339f
C427 B.n390 VSUBS 0.010339f
C428 B.n391 VSUBS 0.010339f
C429 B.n392 VSUBS 0.010339f
C430 B.n393 VSUBS 0.010339f
C431 B.n394 VSUBS 0.010339f
C432 B.n395 VSUBS 0.010339f
C433 B.n396 VSUBS 0.010339f
C434 B.n397 VSUBS 0.010339f
C435 B.n398 VSUBS 0.010339f
C436 B.n399 VSUBS 0.010339f
C437 B.n400 VSUBS 0.010339f
C438 B.n401 VSUBS 0.010339f
C439 B.n402 VSUBS 0.010339f
C440 B.n403 VSUBS 0.010339f
C441 B.n404 VSUBS 0.007146f
C442 B.n405 VSUBS 0.023955f
C443 B.n406 VSUBS 0.008363f
C444 B.n407 VSUBS 0.010339f
C445 B.n408 VSUBS 0.010339f
C446 B.n409 VSUBS 0.010339f
C447 B.n410 VSUBS 0.010339f
C448 B.n411 VSUBS 0.010339f
C449 B.n412 VSUBS 0.010339f
C450 B.n413 VSUBS 0.010339f
C451 B.n414 VSUBS 0.010339f
C452 B.n415 VSUBS 0.010339f
C453 B.n416 VSUBS 0.010339f
C454 B.n417 VSUBS 0.010339f
C455 B.t8 VSUBS 0.185482f
C456 B.t7 VSUBS 0.243405f
C457 B.t6 VSUBS 2.14522f
C458 B.n418 VSUBS 0.394955f
C459 B.n419 VSUBS 0.289485f
C460 B.n420 VSUBS 0.023955f
C461 B.n421 VSUBS 0.008363f
C462 B.n422 VSUBS 0.010339f
C463 B.n423 VSUBS 0.010339f
C464 B.n424 VSUBS 0.010339f
C465 B.n425 VSUBS 0.010339f
C466 B.n426 VSUBS 0.010339f
C467 B.n427 VSUBS 0.010339f
C468 B.n428 VSUBS 0.010339f
C469 B.n429 VSUBS 0.010339f
C470 B.n430 VSUBS 0.010339f
C471 B.n431 VSUBS 0.010339f
C472 B.n432 VSUBS 0.010339f
C473 B.n433 VSUBS 0.010339f
C474 B.n434 VSUBS 0.010339f
C475 B.n435 VSUBS 0.010339f
C476 B.n436 VSUBS 0.010339f
C477 B.n437 VSUBS 0.010339f
C478 B.n438 VSUBS 0.010339f
C479 B.n439 VSUBS 0.010339f
C480 B.n440 VSUBS 0.010339f
C481 B.n441 VSUBS 0.010339f
C482 B.n442 VSUBS 0.010339f
C483 B.n443 VSUBS 0.010339f
C484 B.n444 VSUBS 0.010339f
C485 B.n445 VSUBS 0.010339f
C486 B.n446 VSUBS 0.010339f
C487 B.n447 VSUBS 0.010339f
C488 B.n448 VSUBS 0.010339f
C489 B.n449 VSUBS 0.010339f
C490 B.n450 VSUBS 0.010339f
C491 B.n451 VSUBS 0.010339f
C492 B.n452 VSUBS 0.010339f
C493 B.n453 VSUBS 0.010339f
C494 B.n454 VSUBS 0.010339f
C495 B.n455 VSUBS 0.010339f
C496 B.n456 VSUBS 0.010339f
C497 B.n457 VSUBS 0.010339f
C498 B.n458 VSUBS 0.010339f
C499 B.n459 VSUBS 0.010339f
C500 B.n460 VSUBS 0.010339f
C501 B.n461 VSUBS 0.010339f
C502 B.n462 VSUBS 0.010339f
C503 B.n463 VSUBS 0.010339f
C504 B.n464 VSUBS 0.010339f
C505 B.n465 VSUBS 0.010339f
C506 B.n466 VSUBS 0.025835f
C507 B.n467 VSUBS 0.024679f
C508 B.n468 VSUBS 0.025497f
C509 B.n469 VSUBS 0.010339f
C510 B.n470 VSUBS 0.010339f
C511 B.n471 VSUBS 0.010339f
C512 B.n472 VSUBS 0.010339f
C513 B.n473 VSUBS 0.010339f
C514 B.n474 VSUBS 0.010339f
C515 B.n475 VSUBS 0.010339f
C516 B.n476 VSUBS 0.010339f
C517 B.n477 VSUBS 0.010339f
C518 B.n478 VSUBS 0.010339f
C519 B.n479 VSUBS 0.010339f
C520 B.n480 VSUBS 0.010339f
C521 B.n481 VSUBS 0.010339f
C522 B.n482 VSUBS 0.010339f
C523 B.n483 VSUBS 0.010339f
C524 B.n484 VSUBS 0.010339f
C525 B.n485 VSUBS 0.010339f
C526 B.n486 VSUBS 0.010339f
C527 B.n487 VSUBS 0.010339f
C528 B.n488 VSUBS 0.010339f
C529 B.n489 VSUBS 0.010339f
C530 B.n490 VSUBS 0.010339f
C531 B.n491 VSUBS 0.010339f
C532 B.n492 VSUBS 0.010339f
C533 B.n493 VSUBS 0.010339f
C534 B.n494 VSUBS 0.010339f
C535 B.n495 VSUBS 0.010339f
C536 B.n496 VSUBS 0.010339f
C537 B.n497 VSUBS 0.010339f
C538 B.n498 VSUBS 0.010339f
C539 B.n499 VSUBS 0.010339f
C540 B.n500 VSUBS 0.010339f
C541 B.n501 VSUBS 0.010339f
C542 B.n502 VSUBS 0.010339f
C543 B.n503 VSUBS 0.010339f
C544 B.n504 VSUBS 0.010339f
C545 B.n505 VSUBS 0.010339f
C546 B.n506 VSUBS 0.010339f
C547 B.n507 VSUBS 0.010339f
C548 B.n508 VSUBS 0.010339f
C549 B.n509 VSUBS 0.010339f
C550 B.n510 VSUBS 0.010339f
C551 B.n511 VSUBS 0.010339f
C552 B.n512 VSUBS 0.010339f
C553 B.n513 VSUBS 0.010339f
C554 B.n514 VSUBS 0.010339f
C555 B.n515 VSUBS 0.010339f
C556 B.n516 VSUBS 0.010339f
C557 B.n517 VSUBS 0.010339f
C558 B.n518 VSUBS 0.010339f
C559 B.n519 VSUBS 0.010339f
C560 B.n520 VSUBS 0.010339f
C561 B.n521 VSUBS 0.010339f
C562 B.n522 VSUBS 0.010339f
C563 B.n523 VSUBS 0.010339f
C564 B.n524 VSUBS 0.010339f
C565 B.n525 VSUBS 0.010339f
C566 B.n526 VSUBS 0.010339f
C567 B.n527 VSUBS 0.010339f
C568 B.n528 VSUBS 0.010339f
C569 B.n529 VSUBS 0.010339f
C570 B.n530 VSUBS 0.010339f
C571 B.n531 VSUBS 0.010339f
C572 B.n532 VSUBS 0.010339f
C573 B.n533 VSUBS 0.010339f
C574 B.n534 VSUBS 0.010339f
C575 B.n535 VSUBS 0.010339f
C576 B.n536 VSUBS 0.010339f
C577 B.n537 VSUBS 0.010339f
C578 B.n538 VSUBS 0.010339f
C579 B.n539 VSUBS 0.010339f
C580 B.n540 VSUBS 0.010339f
C581 B.n541 VSUBS 0.010339f
C582 B.n542 VSUBS 0.010339f
C583 B.n543 VSUBS 0.010339f
C584 B.n544 VSUBS 0.010339f
C585 B.n545 VSUBS 0.010339f
C586 B.n546 VSUBS 0.010339f
C587 B.n547 VSUBS 0.010339f
C588 B.n548 VSUBS 0.010339f
C589 B.n549 VSUBS 0.010339f
C590 B.n550 VSUBS 0.010339f
C591 B.n551 VSUBS 0.010339f
C592 B.n552 VSUBS 0.010339f
C593 B.n553 VSUBS 0.010339f
C594 B.n554 VSUBS 0.010339f
C595 B.n555 VSUBS 0.010339f
C596 B.n556 VSUBS 0.010339f
C597 B.n557 VSUBS 0.010339f
C598 B.n558 VSUBS 0.010339f
C599 B.n559 VSUBS 0.010339f
C600 B.n560 VSUBS 0.010339f
C601 B.n561 VSUBS 0.010339f
C602 B.n562 VSUBS 0.010339f
C603 B.n563 VSUBS 0.010339f
C604 B.n564 VSUBS 0.010339f
C605 B.n565 VSUBS 0.010339f
C606 B.n566 VSUBS 0.010339f
C607 B.n567 VSUBS 0.010339f
C608 B.n568 VSUBS 0.010339f
C609 B.n569 VSUBS 0.010339f
C610 B.n570 VSUBS 0.010339f
C611 B.n571 VSUBS 0.010339f
C612 B.n572 VSUBS 0.010339f
C613 B.n573 VSUBS 0.010339f
C614 B.n574 VSUBS 0.010339f
C615 B.n575 VSUBS 0.010339f
C616 B.n576 VSUBS 0.010339f
C617 B.n577 VSUBS 0.010339f
C618 B.n578 VSUBS 0.010339f
C619 B.n579 VSUBS 0.010339f
C620 B.n580 VSUBS 0.010339f
C621 B.n581 VSUBS 0.010339f
C622 B.n582 VSUBS 0.010339f
C623 B.n583 VSUBS 0.010339f
C624 B.n584 VSUBS 0.010339f
C625 B.n585 VSUBS 0.010339f
C626 B.n586 VSUBS 0.010339f
C627 B.n587 VSUBS 0.010339f
C628 B.n588 VSUBS 0.010339f
C629 B.n589 VSUBS 0.010339f
C630 B.n590 VSUBS 0.010339f
C631 B.n591 VSUBS 0.010339f
C632 B.n592 VSUBS 0.010339f
C633 B.n593 VSUBS 0.010339f
C634 B.n594 VSUBS 0.010339f
C635 B.n595 VSUBS 0.010339f
C636 B.n596 VSUBS 0.010339f
C637 B.n597 VSUBS 0.010339f
C638 B.n598 VSUBS 0.010339f
C639 B.n599 VSUBS 0.010339f
C640 B.n600 VSUBS 0.010339f
C641 B.n601 VSUBS 0.010339f
C642 B.n602 VSUBS 0.010339f
C643 B.n603 VSUBS 0.010339f
C644 B.n604 VSUBS 0.010339f
C645 B.n605 VSUBS 0.010339f
C646 B.n606 VSUBS 0.010339f
C647 B.n607 VSUBS 0.010339f
C648 B.n608 VSUBS 0.010339f
C649 B.n609 VSUBS 0.010339f
C650 B.n610 VSUBS 0.010339f
C651 B.n611 VSUBS 0.010339f
C652 B.n612 VSUBS 0.010339f
C653 B.n613 VSUBS 0.010339f
C654 B.n614 VSUBS 0.010339f
C655 B.n615 VSUBS 0.010339f
C656 B.n616 VSUBS 0.010339f
C657 B.n617 VSUBS 0.010339f
C658 B.n618 VSUBS 0.010339f
C659 B.n619 VSUBS 0.010339f
C660 B.n620 VSUBS 0.010339f
C661 B.n621 VSUBS 0.010339f
C662 B.n622 VSUBS 0.010339f
C663 B.n623 VSUBS 0.010339f
C664 B.n624 VSUBS 0.010339f
C665 B.n625 VSUBS 0.010339f
C666 B.n626 VSUBS 0.010339f
C667 B.n627 VSUBS 0.010339f
C668 B.n628 VSUBS 0.010339f
C669 B.n629 VSUBS 0.010339f
C670 B.n630 VSUBS 0.010339f
C671 B.n631 VSUBS 0.010339f
C672 B.n632 VSUBS 0.010339f
C673 B.n633 VSUBS 0.010339f
C674 B.n634 VSUBS 0.010339f
C675 B.n635 VSUBS 0.010339f
C676 B.n636 VSUBS 0.010339f
C677 B.n637 VSUBS 0.010339f
C678 B.n638 VSUBS 0.010339f
C679 B.n639 VSUBS 0.010339f
C680 B.n640 VSUBS 0.010339f
C681 B.n641 VSUBS 0.010339f
C682 B.n642 VSUBS 0.010339f
C683 B.n643 VSUBS 0.010339f
C684 B.n644 VSUBS 0.010339f
C685 B.n645 VSUBS 0.010339f
C686 B.n646 VSUBS 0.010339f
C687 B.n647 VSUBS 0.010339f
C688 B.n648 VSUBS 0.010339f
C689 B.n649 VSUBS 0.010339f
C690 B.n650 VSUBS 0.010339f
C691 B.n651 VSUBS 0.010339f
C692 B.n652 VSUBS 0.010339f
C693 B.n653 VSUBS 0.010339f
C694 B.n654 VSUBS 0.010339f
C695 B.n655 VSUBS 0.010339f
C696 B.n656 VSUBS 0.010339f
C697 B.n657 VSUBS 0.010339f
C698 B.n658 VSUBS 0.010339f
C699 B.n659 VSUBS 0.010339f
C700 B.n660 VSUBS 0.010339f
C701 B.n661 VSUBS 0.010339f
C702 B.n662 VSUBS 0.010339f
C703 B.n663 VSUBS 0.010339f
C704 B.n664 VSUBS 0.010339f
C705 B.n665 VSUBS 0.010339f
C706 B.n666 VSUBS 0.010339f
C707 B.n667 VSUBS 0.010339f
C708 B.n668 VSUBS 0.010339f
C709 B.n669 VSUBS 0.010339f
C710 B.n670 VSUBS 0.010339f
C711 B.n671 VSUBS 0.010339f
C712 B.n672 VSUBS 0.010339f
C713 B.n673 VSUBS 0.010339f
C714 B.n674 VSUBS 0.010339f
C715 B.n675 VSUBS 0.010339f
C716 B.n676 VSUBS 0.010339f
C717 B.n677 VSUBS 0.010339f
C718 B.n678 VSUBS 0.010339f
C719 B.n679 VSUBS 0.010339f
C720 B.n680 VSUBS 0.010339f
C721 B.n681 VSUBS 0.010339f
C722 B.n682 VSUBS 0.010339f
C723 B.n683 VSUBS 0.010339f
C724 B.n684 VSUBS 0.010339f
C725 B.n685 VSUBS 0.010339f
C726 B.n686 VSUBS 0.010339f
C727 B.n687 VSUBS 0.010339f
C728 B.n688 VSUBS 0.010339f
C729 B.n689 VSUBS 0.010339f
C730 B.n690 VSUBS 0.010339f
C731 B.n691 VSUBS 0.010339f
C732 B.n692 VSUBS 0.010339f
C733 B.n693 VSUBS 0.010339f
C734 B.n694 VSUBS 0.010339f
C735 B.n695 VSUBS 0.010339f
C736 B.n696 VSUBS 0.010339f
C737 B.n697 VSUBS 0.010339f
C738 B.n698 VSUBS 0.010339f
C739 B.n699 VSUBS 0.010339f
C740 B.n700 VSUBS 0.010339f
C741 B.n701 VSUBS 0.010339f
C742 B.n702 VSUBS 0.010339f
C743 B.n703 VSUBS 0.010339f
C744 B.n704 VSUBS 0.010339f
C745 B.n705 VSUBS 0.010339f
C746 B.n706 VSUBS 0.010339f
C747 B.n707 VSUBS 0.010339f
C748 B.n708 VSUBS 0.010339f
C749 B.n709 VSUBS 0.010339f
C750 B.n710 VSUBS 0.010339f
C751 B.n711 VSUBS 0.010339f
C752 B.n712 VSUBS 0.02434f
C753 B.n713 VSUBS 0.02434f
C754 B.n714 VSUBS 0.025835f
C755 B.n715 VSUBS 0.010339f
C756 B.n716 VSUBS 0.010339f
C757 B.n717 VSUBS 0.010339f
C758 B.n718 VSUBS 0.010339f
C759 B.n719 VSUBS 0.010339f
C760 B.n720 VSUBS 0.010339f
C761 B.n721 VSUBS 0.010339f
C762 B.n722 VSUBS 0.010339f
C763 B.n723 VSUBS 0.010339f
C764 B.n724 VSUBS 0.010339f
C765 B.n725 VSUBS 0.010339f
C766 B.n726 VSUBS 0.010339f
C767 B.n727 VSUBS 0.010339f
C768 B.n728 VSUBS 0.010339f
C769 B.n729 VSUBS 0.010339f
C770 B.n730 VSUBS 0.010339f
C771 B.n731 VSUBS 0.010339f
C772 B.n732 VSUBS 0.010339f
C773 B.n733 VSUBS 0.010339f
C774 B.n734 VSUBS 0.010339f
C775 B.n735 VSUBS 0.010339f
C776 B.n736 VSUBS 0.010339f
C777 B.n737 VSUBS 0.010339f
C778 B.n738 VSUBS 0.010339f
C779 B.n739 VSUBS 0.010339f
C780 B.n740 VSUBS 0.010339f
C781 B.n741 VSUBS 0.010339f
C782 B.n742 VSUBS 0.010339f
C783 B.n743 VSUBS 0.010339f
C784 B.n744 VSUBS 0.010339f
C785 B.n745 VSUBS 0.010339f
C786 B.n746 VSUBS 0.010339f
C787 B.n747 VSUBS 0.010339f
C788 B.n748 VSUBS 0.010339f
C789 B.n749 VSUBS 0.010339f
C790 B.n750 VSUBS 0.010339f
C791 B.n751 VSUBS 0.010339f
C792 B.n752 VSUBS 0.010339f
C793 B.n753 VSUBS 0.010339f
C794 B.n754 VSUBS 0.010339f
C795 B.n755 VSUBS 0.010339f
C796 B.n756 VSUBS 0.010339f
C797 B.n757 VSUBS 0.007146f
C798 B.n758 VSUBS 0.010339f
C799 B.n759 VSUBS 0.010339f
C800 B.n760 VSUBS 0.008363f
C801 B.n761 VSUBS 0.010339f
C802 B.n762 VSUBS 0.010339f
C803 B.n763 VSUBS 0.010339f
C804 B.n764 VSUBS 0.010339f
C805 B.n765 VSUBS 0.010339f
C806 B.n766 VSUBS 0.010339f
C807 B.n767 VSUBS 0.010339f
C808 B.n768 VSUBS 0.010339f
C809 B.n769 VSUBS 0.010339f
C810 B.n770 VSUBS 0.010339f
C811 B.n771 VSUBS 0.010339f
C812 B.n772 VSUBS 0.008363f
C813 B.n773 VSUBS 0.023955f
C814 B.n774 VSUBS 0.007146f
C815 B.n775 VSUBS 0.010339f
C816 B.n776 VSUBS 0.010339f
C817 B.n777 VSUBS 0.010339f
C818 B.n778 VSUBS 0.010339f
C819 B.n779 VSUBS 0.010339f
C820 B.n780 VSUBS 0.010339f
C821 B.n781 VSUBS 0.010339f
C822 B.n782 VSUBS 0.010339f
C823 B.n783 VSUBS 0.010339f
C824 B.n784 VSUBS 0.010339f
C825 B.n785 VSUBS 0.010339f
C826 B.n786 VSUBS 0.010339f
C827 B.n787 VSUBS 0.010339f
C828 B.n788 VSUBS 0.010339f
C829 B.n789 VSUBS 0.010339f
C830 B.n790 VSUBS 0.010339f
C831 B.n791 VSUBS 0.010339f
C832 B.n792 VSUBS 0.010339f
C833 B.n793 VSUBS 0.010339f
C834 B.n794 VSUBS 0.010339f
C835 B.n795 VSUBS 0.010339f
C836 B.n796 VSUBS 0.010339f
C837 B.n797 VSUBS 0.010339f
C838 B.n798 VSUBS 0.010339f
C839 B.n799 VSUBS 0.010339f
C840 B.n800 VSUBS 0.010339f
C841 B.n801 VSUBS 0.010339f
C842 B.n802 VSUBS 0.010339f
C843 B.n803 VSUBS 0.010339f
C844 B.n804 VSUBS 0.010339f
C845 B.n805 VSUBS 0.010339f
C846 B.n806 VSUBS 0.010339f
C847 B.n807 VSUBS 0.010339f
C848 B.n808 VSUBS 0.010339f
C849 B.n809 VSUBS 0.010339f
C850 B.n810 VSUBS 0.010339f
C851 B.n811 VSUBS 0.010339f
C852 B.n812 VSUBS 0.010339f
C853 B.n813 VSUBS 0.010339f
C854 B.n814 VSUBS 0.010339f
C855 B.n815 VSUBS 0.010339f
C856 B.n816 VSUBS 0.010339f
C857 B.n817 VSUBS 0.025835f
C858 B.n818 VSUBS 0.025835f
C859 B.n819 VSUBS 0.02434f
C860 B.n820 VSUBS 0.010339f
C861 B.n821 VSUBS 0.010339f
C862 B.n822 VSUBS 0.010339f
C863 B.n823 VSUBS 0.010339f
C864 B.n824 VSUBS 0.010339f
C865 B.n825 VSUBS 0.010339f
C866 B.n826 VSUBS 0.010339f
C867 B.n827 VSUBS 0.010339f
C868 B.n828 VSUBS 0.010339f
C869 B.n829 VSUBS 0.010339f
C870 B.n830 VSUBS 0.010339f
C871 B.n831 VSUBS 0.010339f
C872 B.n832 VSUBS 0.010339f
C873 B.n833 VSUBS 0.010339f
C874 B.n834 VSUBS 0.010339f
C875 B.n835 VSUBS 0.010339f
C876 B.n836 VSUBS 0.010339f
C877 B.n837 VSUBS 0.010339f
C878 B.n838 VSUBS 0.010339f
C879 B.n839 VSUBS 0.010339f
C880 B.n840 VSUBS 0.010339f
C881 B.n841 VSUBS 0.010339f
C882 B.n842 VSUBS 0.010339f
C883 B.n843 VSUBS 0.010339f
C884 B.n844 VSUBS 0.010339f
C885 B.n845 VSUBS 0.010339f
C886 B.n846 VSUBS 0.010339f
C887 B.n847 VSUBS 0.010339f
C888 B.n848 VSUBS 0.010339f
C889 B.n849 VSUBS 0.010339f
C890 B.n850 VSUBS 0.010339f
C891 B.n851 VSUBS 0.010339f
C892 B.n852 VSUBS 0.010339f
C893 B.n853 VSUBS 0.010339f
C894 B.n854 VSUBS 0.010339f
C895 B.n855 VSUBS 0.010339f
C896 B.n856 VSUBS 0.010339f
C897 B.n857 VSUBS 0.010339f
C898 B.n858 VSUBS 0.010339f
C899 B.n859 VSUBS 0.010339f
C900 B.n860 VSUBS 0.010339f
C901 B.n861 VSUBS 0.010339f
C902 B.n862 VSUBS 0.010339f
C903 B.n863 VSUBS 0.010339f
C904 B.n864 VSUBS 0.010339f
C905 B.n865 VSUBS 0.010339f
C906 B.n866 VSUBS 0.010339f
C907 B.n867 VSUBS 0.010339f
C908 B.n868 VSUBS 0.010339f
C909 B.n869 VSUBS 0.010339f
C910 B.n870 VSUBS 0.010339f
C911 B.n871 VSUBS 0.010339f
C912 B.n872 VSUBS 0.010339f
C913 B.n873 VSUBS 0.010339f
C914 B.n874 VSUBS 0.010339f
C915 B.n875 VSUBS 0.010339f
C916 B.n876 VSUBS 0.010339f
C917 B.n877 VSUBS 0.010339f
C918 B.n878 VSUBS 0.010339f
C919 B.n879 VSUBS 0.010339f
C920 B.n880 VSUBS 0.010339f
C921 B.n881 VSUBS 0.010339f
C922 B.n882 VSUBS 0.010339f
C923 B.n883 VSUBS 0.010339f
C924 B.n884 VSUBS 0.010339f
C925 B.n885 VSUBS 0.010339f
C926 B.n886 VSUBS 0.010339f
C927 B.n887 VSUBS 0.010339f
C928 B.n888 VSUBS 0.010339f
C929 B.n889 VSUBS 0.010339f
C930 B.n890 VSUBS 0.010339f
C931 B.n891 VSUBS 0.010339f
C932 B.n892 VSUBS 0.010339f
C933 B.n893 VSUBS 0.010339f
C934 B.n894 VSUBS 0.010339f
C935 B.n895 VSUBS 0.010339f
C936 B.n896 VSUBS 0.010339f
C937 B.n897 VSUBS 0.010339f
C938 B.n898 VSUBS 0.010339f
C939 B.n899 VSUBS 0.010339f
C940 B.n900 VSUBS 0.010339f
C941 B.n901 VSUBS 0.010339f
C942 B.n902 VSUBS 0.010339f
C943 B.n903 VSUBS 0.010339f
C944 B.n904 VSUBS 0.010339f
C945 B.n905 VSUBS 0.010339f
C946 B.n906 VSUBS 0.010339f
C947 B.n907 VSUBS 0.010339f
C948 B.n908 VSUBS 0.010339f
C949 B.n909 VSUBS 0.010339f
C950 B.n910 VSUBS 0.010339f
C951 B.n911 VSUBS 0.010339f
C952 B.n912 VSUBS 0.010339f
C953 B.n913 VSUBS 0.010339f
C954 B.n914 VSUBS 0.010339f
C955 B.n915 VSUBS 0.010339f
C956 B.n916 VSUBS 0.010339f
C957 B.n917 VSUBS 0.010339f
C958 B.n918 VSUBS 0.010339f
C959 B.n919 VSUBS 0.010339f
C960 B.n920 VSUBS 0.010339f
C961 B.n921 VSUBS 0.010339f
C962 B.n922 VSUBS 0.010339f
C963 B.n923 VSUBS 0.010339f
C964 B.n924 VSUBS 0.010339f
C965 B.n925 VSUBS 0.010339f
C966 B.n926 VSUBS 0.010339f
C967 B.n927 VSUBS 0.010339f
C968 B.n928 VSUBS 0.010339f
C969 B.n929 VSUBS 0.010339f
C970 B.n930 VSUBS 0.010339f
C971 B.n931 VSUBS 0.010339f
C972 B.n932 VSUBS 0.010339f
C973 B.n933 VSUBS 0.010339f
C974 B.n934 VSUBS 0.010339f
C975 B.n935 VSUBS 0.010339f
C976 B.n936 VSUBS 0.010339f
C977 B.n937 VSUBS 0.010339f
C978 B.n938 VSUBS 0.010339f
C979 B.n939 VSUBS 0.013492f
C980 B.n940 VSUBS 0.014373f
C981 B.n941 VSUBS 0.028581f
C982 VDD2.n0 VSUBS 0.035606f
C983 VDD2.n1 VSUBS 0.033703f
C984 VDD2.n2 VSUBS 0.018643f
C985 VDD2.n3 VSUBS 0.042807f
C986 VDD2.n4 VSUBS 0.019176f
C987 VDD2.n5 VSUBS 0.033703f
C988 VDD2.n6 VSUBS 0.018111f
C989 VDD2.n7 VSUBS 0.042807f
C990 VDD2.n8 VSUBS 0.019176f
C991 VDD2.n9 VSUBS 0.033703f
C992 VDD2.n10 VSUBS 0.018111f
C993 VDD2.n11 VSUBS 0.032105f
C994 VDD2.n12 VSUBS 0.032201f
C995 VDD2.t4 VSUBS 0.091942f
C996 VDD2.n13 VSUBS 0.203846f
C997 VDD2.n14 VSUBS 1.05756f
C998 VDD2.n15 VSUBS 0.018111f
C999 VDD2.n16 VSUBS 0.019176f
C1000 VDD2.n17 VSUBS 0.042807f
C1001 VDD2.n18 VSUBS 0.042807f
C1002 VDD2.n19 VSUBS 0.019176f
C1003 VDD2.n20 VSUBS 0.018111f
C1004 VDD2.n21 VSUBS 0.033703f
C1005 VDD2.n22 VSUBS 0.033703f
C1006 VDD2.n23 VSUBS 0.018111f
C1007 VDD2.n24 VSUBS 0.019176f
C1008 VDD2.n25 VSUBS 0.042807f
C1009 VDD2.n26 VSUBS 0.042807f
C1010 VDD2.n27 VSUBS 0.019176f
C1011 VDD2.n28 VSUBS 0.018111f
C1012 VDD2.n29 VSUBS 0.033703f
C1013 VDD2.n30 VSUBS 0.033703f
C1014 VDD2.n31 VSUBS 0.018111f
C1015 VDD2.n32 VSUBS 0.018111f
C1016 VDD2.n33 VSUBS 0.019176f
C1017 VDD2.n34 VSUBS 0.042807f
C1018 VDD2.n35 VSUBS 0.042807f
C1019 VDD2.n36 VSUBS 0.098771f
C1020 VDD2.n37 VSUBS 0.018643f
C1021 VDD2.n38 VSUBS 0.018111f
C1022 VDD2.n39 VSUBS 0.084809f
C1023 VDD2.n40 VSUBS 0.102699f
C1024 VDD2.t3 VSUBS 0.211734f
C1025 VDD2.t1 VSUBS 0.211734f
C1026 VDD2.n41 VSUBS 1.53333f
C1027 VDD2.n42 VSUBS 1.47944f
C1028 VDD2.t8 VSUBS 0.211734f
C1029 VDD2.t7 VSUBS 0.211734f
C1030 VDD2.n43 VSUBS 1.57112f
C1031 VDD2.n44 VSUBS 4.73879f
C1032 VDD2.n45 VSUBS 0.035606f
C1033 VDD2.n46 VSUBS 0.033703f
C1034 VDD2.n47 VSUBS 0.018643f
C1035 VDD2.n48 VSUBS 0.042807f
C1036 VDD2.n49 VSUBS 0.018111f
C1037 VDD2.n50 VSUBS 0.019176f
C1038 VDD2.n51 VSUBS 0.033703f
C1039 VDD2.n52 VSUBS 0.018111f
C1040 VDD2.n53 VSUBS 0.042807f
C1041 VDD2.n54 VSUBS 0.019176f
C1042 VDD2.n55 VSUBS 0.033703f
C1043 VDD2.n56 VSUBS 0.018111f
C1044 VDD2.n57 VSUBS 0.032105f
C1045 VDD2.n58 VSUBS 0.032201f
C1046 VDD2.t5 VSUBS 0.091942f
C1047 VDD2.n59 VSUBS 0.203846f
C1048 VDD2.n60 VSUBS 1.05756f
C1049 VDD2.n61 VSUBS 0.018111f
C1050 VDD2.n62 VSUBS 0.019176f
C1051 VDD2.n63 VSUBS 0.042807f
C1052 VDD2.n64 VSUBS 0.042807f
C1053 VDD2.n65 VSUBS 0.019176f
C1054 VDD2.n66 VSUBS 0.018111f
C1055 VDD2.n67 VSUBS 0.033703f
C1056 VDD2.n68 VSUBS 0.033703f
C1057 VDD2.n69 VSUBS 0.018111f
C1058 VDD2.n70 VSUBS 0.019176f
C1059 VDD2.n71 VSUBS 0.042807f
C1060 VDD2.n72 VSUBS 0.042807f
C1061 VDD2.n73 VSUBS 0.019176f
C1062 VDD2.n74 VSUBS 0.018111f
C1063 VDD2.n75 VSUBS 0.033703f
C1064 VDD2.n76 VSUBS 0.033703f
C1065 VDD2.n77 VSUBS 0.018111f
C1066 VDD2.n78 VSUBS 0.019176f
C1067 VDD2.n79 VSUBS 0.042807f
C1068 VDD2.n80 VSUBS 0.042807f
C1069 VDD2.n81 VSUBS 0.098771f
C1070 VDD2.n82 VSUBS 0.018643f
C1071 VDD2.n83 VSUBS 0.018111f
C1072 VDD2.n84 VSUBS 0.084809f
C1073 VDD2.n85 VSUBS 0.072881f
C1074 VDD2.n86 VSUBS 4.13238f
C1075 VDD2.t9 VSUBS 0.211734f
C1076 VDD2.t2 VSUBS 0.211734f
C1077 VDD2.n87 VSUBS 1.53334f
C1078 VDD2.n88 VSUBS 1.06141f
C1079 VDD2.t0 VSUBS 0.211734f
C1080 VDD2.t6 VSUBS 0.211734f
C1081 VDD2.n89 VSUBS 1.57107f
C1082 VN.t2 VSUBS 2.20927f
C1083 VN.n0 VSUBS 0.897859f
C1084 VN.n1 VSUBS 0.026953f
C1085 VN.n2 VSUBS 0.053432f
C1086 VN.n3 VSUBS 0.026953f
C1087 VN.n4 VSUBS 0.050234f
C1088 VN.n5 VSUBS 0.026953f
C1089 VN.t1 VSUBS 2.20927f
C1090 VN.n6 VSUBS 0.050234f
C1091 VN.n7 VSUBS 0.026953f
C1092 VN.n8 VSUBS 0.050234f
C1093 VN.n9 VSUBS 0.026953f
C1094 VN.t8 VSUBS 2.20927f
C1095 VN.n10 VSUBS 0.050234f
C1096 VN.n11 VSUBS 0.026953f
C1097 VN.n12 VSUBS 0.050234f
C1098 VN.t5 VSUBS 2.61326f
C1099 VN.n13 VSUBS 0.856492f
C1100 VN.t6 VSUBS 2.20927f
C1101 VN.n14 VSUBS 0.899754f
C1102 VN.n15 VSUBS 0.046266f
C1103 VN.n16 VSUBS 0.346905f
C1104 VN.n17 VSUBS 0.026953f
C1105 VN.n18 VSUBS 0.026953f
C1106 VN.n19 VSUBS 0.050234f
C1107 VN.n20 VSUBS 0.032965f
C1108 VN.n21 VSUBS 0.045734f
C1109 VN.n22 VSUBS 0.026953f
C1110 VN.n23 VSUBS 0.026953f
C1111 VN.n24 VSUBS 0.026953f
C1112 VN.n25 VSUBS 0.050234f
C1113 VN.n26 VSUBS 0.037834f
C1114 VN.n27 VSUBS 0.793453f
C1115 VN.n28 VSUBS 0.037834f
C1116 VN.n29 VSUBS 0.026953f
C1117 VN.n30 VSUBS 0.026953f
C1118 VN.n31 VSUBS 0.026953f
C1119 VN.n32 VSUBS 0.050234f
C1120 VN.n33 VSUBS 0.045734f
C1121 VN.n34 VSUBS 0.032965f
C1122 VN.n35 VSUBS 0.026953f
C1123 VN.n36 VSUBS 0.026953f
C1124 VN.n37 VSUBS 0.026953f
C1125 VN.n38 VSUBS 0.050234f
C1126 VN.n39 VSUBS 0.046266f
C1127 VN.n40 VSUBS 0.793453f
C1128 VN.n41 VSUBS 0.029401f
C1129 VN.n42 VSUBS 0.026953f
C1130 VN.n43 VSUBS 0.026953f
C1131 VN.n44 VSUBS 0.026953f
C1132 VN.n45 VSUBS 0.050234f
C1133 VN.n46 VSUBS 0.053702f
C1134 VN.n47 VSUBS 0.021799f
C1135 VN.n48 VSUBS 0.026953f
C1136 VN.n49 VSUBS 0.026953f
C1137 VN.n50 VSUBS 0.026953f
C1138 VN.n51 VSUBS 0.050234f
C1139 VN.n52 VSUBS 0.050234f
C1140 VN.n53 VSUBS 0.029897f
C1141 VN.n54 VSUBS 0.043502f
C1142 VN.n55 VSUBS 0.082135f
C1143 VN.t4 VSUBS 2.20927f
C1144 VN.n56 VSUBS 0.897859f
C1145 VN.n57 VSUBS 0.026953f
C1146 VN.n58 VSUBS 0.053432f
C1147 VN.n59 VSUBS 0.026953f
C1148 VN.n60 VSUBS 0.050234f
C1149 VN.n61 VSUBS 0.026953f
C1150 VN.t0 VSUBS 2.20927f
C1151 VN.n62 VSUBS 0.050234f
C1152 VN.n63 VSUBS 0.026953f
C1153 VN.n64 VSUBS 0.050234f
C1154 VN.n65 VSUBS 0.026953f
C1155 VN.t7 VSUBS 2.20927f
C1156 VN.n66 VSUBS 0.050234f
C1157 VN.n67 VSUBS 0.026953f
C1158 VN.n68 VSUBS 0.050234f
C1159 VN.t3 VSUBS 2.61326f
C1160 VN.n69 VSUBS 0.856492f
C1161 VN.t9 VSUBS 2.20927f
C1162 VN.n70 VSUBS 0.899754f
C1163 VN.n71 VSUBS 0.046266f
C1164 VN.n72 VSUBS 0.346905f
C1165 VN.n73 VSUBS 0.026953f
C1166 VN.n74 VSUBS 0.026953f
C1167 VN.n75 VSUBS 0.050234f
C1168 VN.n76 VSUBS 0.032965f
C1169 VN.n77 VSUBS 0.045734f
C1170 VN.n78 VSUBS 0.026953f
C1171 VN.n79 VSUBS 0.026953f
C1172 VN.n80 VSUBS 0.026953f
C1173 VN.n81 VSUBS 0.050234f
C1174 VN.n82 VSUBS 0.037834f
C1175 VN.n83 VSUBS 0.793453f
C1176 VN.n84 VSUBS 0.037834f
C1177 VN.n85 VSUBS 0.026953f
C1178 VN.n86 VSUBS 0.026953f
C1179 VN.n87 VSUBS 0.026953f
C1180 VN.n88 VSUBS 0.050234f
C1181 VN.n89 VSUBS 0.045734f
C1182 VN.n90 VSUBS 0.032965f
C1183 VN.n91 VSUBS 0.026953f
C1184 VN.n92 VSUBS 0.026953f
C1185 VN.n93 VSUBS 0.026953f
C1186 VN.n94 VSUBS 0.050234f
C1187 VN.n95 VSUBS 0.046266f
C1188 VN.n96 VSUBS 0.793453f
C1189 VN.n97 VSUBS 0.029401f
C1190 VN.n98 VSUBS 0.026953f
C1191 VN.n99 VSUBS 0.026953f
C1192 VN.n100 VSUBS 0.026953f
C1193 VN.n101 VSUBS 0.050234f
C1194 VN.n102 VSUBS 0.053702f
C1195 VN.n103 VSUBS 0.021799f
C1196 VN.n104 VSUBS 0.026953f
C1197 VN.n105 VSUBS 0.026953f
C1198 VN.n106 VSUBS 0.026953f
C1199 VN.n107 VSUBS 0.050234f
C1200 VN.n108 VSUBS 0.050234f
C1201 VN.n109 VSUBS 0.029897f
C1202 VN.n110 VSUBS 0.043502f
C1203 VN.n111 VSUBS 1.86477f
C1204 VDD1.n0 VSUBS 0.035708f
C1205 VDD1.n1 VSUBS 0.0338f
C1206 VDD1.n2 VSUBS 0.018697f
C1207 VDD1.n3 VSUBS 0.04293f
C1208 VDD1.n4 VSUBS 0.018163f
C1209 VDD1.n5 VSUBS 0.019231f
C1210 VDD1.n6 VSUBS 0.0338f
C1211 VDD1.n7 VSUBS 0.018163f
C1212 VDD1.n8 VSUBS 0.04293f
C1213 VDD1.n9 VSUBS 0.019231f
C1214 VDD1.n10 VSUBS 0.0338f
C1215 VDD1.n11 VSUBS 0.018163f
C1216 VDD1.n12 VSUBS 0.032197f
C1217 VDD1.n13 VSUBS 0.032293f
C1218 VDD1.t7 VSUBS 0.092206f
C1219 VDD1.n14 VSUBS 0.204431f
C1220 VDD1.n15 VSUBS 1.0606f
C1221 VDD1.n16 VSUBS 0.018163f
C1222 VDD1.n17 VSUBS 0.019231f
C1223 VDD1.n18 VSUBS 0.04293f
C1224 VDD1.n19 VSUBS 0.04293f
C1225 VDD1.n20 VSUBS 0.019231f
C1226 VDD1.n21 VSUBS 0.018163f
C1227 VDD1.n22 VSUBS 0.0338f
C1228 VDD1.n23 VSUBS 0.0338f
C1229 VDD1.n24 VSUBS 0.018163f
C1230 VDD1.n25 VSUBS 0.019231f
C1231 VDD1.n26 VSUBS 0.04293f
C1232 VDD1.n27 VSUBS 0.04293f
C1233 VDD1.n28 VSUBS 0.019231f
C1234 VDD1.n29 VSUBS 0.018163f
C1235 VDD1.n30 VSUBS 0.0338f
C1236 VDD1.n31 VSUBS 0.0338f
C1237 VDD1.n32 VSUBS 0.018163f
C1238 VDD1.n33 VSUBS 0.019231f
C1239 VDD1.n34 VSUBS 0.04293f
C1240 VDD1.n35 VSUBS 0.04293f
C1241 VDD1.n36 VSUBS 0.099054f
C1242 VDD1.n37 VSUBS 0.018697f
C1243 VDD1.n38 VSUBS 0.018163f
C1244 VDD1.n39 VSUBS 0.085052f
C1245 VDD1.n40 VSUBS 0.102993f
C1246 VDD1.t2 VSUBS 0.212341f
C1247 VDD1.t9 VSUBS 0.212341f
C1248 VDD1.n41 VSUBS 1.53774f
C1249 VDD1.n42 VSUBS 1.49512f
C1250 VDD1.n43 VSUBS 0.035708f
C1251 VDD1.n44 VSUBS 0.0338f
C1252 VDD1.n45 VSUBS 0.018697f
C1253 VDD1.n46 VSUBS 0.04293f
C1254 VDD1.n47 VSUBS 0.019231f
C1255 VDD1.n48 VSUBS 0.0338f
C1256 VDD1.n49 VSUBS 0.018163f
C1257 VDD1.n50 VSUBS 0.04293f
C1258 VDD1.n51 VSUBS 0.019231f
C1259 VDD1.n52 VSUBS 0.0338f
C1260 VDD1.n53 VSUBS 0.018163f
C1261 VDD1.n54 VSUBS 0.032197f
C1262 VDD1.n55 VSUBS 0.032293f
C1263 VDD1.t5 VSUBS 0.092206f
C1264 VDD1.n56 VSUBS 0.204431f
C1265 VDD1.n57 VSUBS 1.0606f
C1266 VDD1.n58 VSUBS 0.018163f
C1267 VDD1.n59 VSUBS 0.019231f
C1268 VDD1.n60 VSUBS 0.04293f
C1269 VDD1.n61 VSUBS 0.04293f
C1270 VDD1.n62 VSUBS 0.019231f
C1271 VDD1.n63 VSUBS 0.018163f
C1272 VDD1.n64 VSUBS 0.0338f
C1273 VDD1.n65 VSUBS 0.0338f
C1274 VDD1.n66 VSUBS 0.018163f
C1275 VDD1.n67 VSUBS 0.019231f
C1276 VDD1.n68 VSUBS 0.04293f
C1277 VDD1.n69 VSUBS 0.04293f
C1278 VDD1.n70 VSUBS 0.019231f
C1279 VDD1.n71 VSUBS 0.018163f
C1280 VDD1.n72 VSUBS 0.0338f
C1281 VDD1.n73 VSUBS 0.0338f
C1282 VDD1.n74 VSUBS 0.018163f
C1283 VDD1.n75 VSUBS 0.018163f
C1284 VDD1.n76 VSUBS 0.019231f
C1285 VDD1.n77 VSUBS 0.04293f
C1286 VDD1.n78 VSUBS 0.04293f
C1287 VDD1.n79 VSUBS 0.099054f
C1288 VDD1.n80 VSUBS 0.018697f
C1289 VDD1.n81 VSUBS 0.018163f
C1290 VDD1.n82 VSUBS 0.085052f
C1291 VDD1.n83 VSUBS 0.102993f
C1292 VDD1.t8 VSUBS 0.212341f
C1293 VDD1.t0 VSUBS 0.212341f
C1294 VDD1.n84 VSUBS 1.53773f
C1295 VDD1.n85 VSUBS 1.48369f
C1296 VDD1.t3 VSUBS 0.212341f
C1297 VDD1.t6 VSUBS 0.212341f
C1298 VDD1.n86 VSUBS 1.57563f
C1299 VDD1.n87 VSUBS 4.96293f
C1300 VDD1.t4 VSUBS 0.212341f
C1301 VDD1.t1 VSUBS 0.212341f
C1302 VDD1.n88 VSUBS 1.53773f
C1303 VDD1.n89 VSUBS 4.85912f
C1304 VTAIL.t4 VSUBS 0.204468f
C1305 VTAIL.t19 VSUBS 0.204468f
C1306 VTAIL.n0 VSUBS 1.34905f
C1307 VTAIL.n1 VSUBS 1.1617f
C1308 VTAIL.n2 VSUBS 0.034384f
C1309 VTAIL.n3 VSUBS 0.032547f
C1310 VTAIL.n4 VSUBS 0.018003f
C1311 VTAIL.n5 VSUBS 0.041338f
C1312 VTAIL.n6 VSUBS 0.018518f
C1313 VTAIL.n7 VSUBS 0.032547f
C1314 VTAIL.n8 VSUBS 0.017489f
C1315 VTAIL.n9 VSUBS 0.041338f
C1316 VTAIL.n10 VSUBS 0.018518f
C1317 VTAIL.n11 VSUBS 0.032547f
C1318 VTAIL.n12 VSUBS 0.017489f
C1319 VTAIL.n13 VSUBS 0.031003f
C1320 VTAIL.n14 VSUBS 0.031096f
C1321 VTAIL.t11 VSUBS 0.088787f
C1322 VTAIL.n15 VSUBS 0.196852f
C1323 VTAIL.n16 VSUBS 1.02128f
C1324 VTAIL.n17 VSUBS 0.017489f
C1325 VTAIL.n18 VSUBS 0.018518f
C1326 VTAIL.n19 VSUBS 0.041338f
C1327 VTAIL.n20 VSUBS 0.041338f
C1328 VTAIL.n21 VSUBS 0.018518f
C1329 VTAIL.n22 VSUBS 0.017489f
C1330 VTAIL.n23 VSUBS 0.032547f
C1331 VTAIL.n24 VSUBS 0.032547f
C1332 VTAIL.n25 VSUBS 0.017489f
C1333 VTAIL.n26 VSUBS 0.018518f
C1334 VTAIL.n27 VSUBS 0.041338f
C1335 VTAIL.n28 VSUBS 0.041338f
C1336 VTAIL.n29 VSUBS 0.018518f
C1337 VTAIL.n30 VSUBS 0.017489f
C1338 VTAIL.n31 VSUBS 0.032547f
C1339 VTAIL.n32 VSUBS 0.032547f
C1340 VTAIL.n33 VSUBS 0.017489f
C1341 VTAIL.n34 VSUBS 0.017489f
C1342 VTAIL.n35 VSUBS 0.018518f
C1343 VTAIL.n36 VSUBS 0.041338f
C1344 VTAIL.n37 VSUBS 0.041338f
C1345 VTAIL.n38 VSUBS 0.095382f
C1346 VTAIL.n39 VSUBS 0.018003f
C1347 VTAIL.n40 VSUBS 0.017489f
C1348 VTAIL.n41 VSUBS 0.081899f
C1349 VTAIL.n42 VSUBS 0.047956f
C1350 VTAIL.n43 VSUBS 0.646338f
C1351 VTAIL.t14 VSUBS 0.204468f
C1352 VTAIL.t13 VSUBS 0.204468f
C1353 VTAIL.n44 VSUBS 1.34905f
C1354 VTAIL.n45 VSUBS 1.38907f
C1355 VTAIL.t9 VSUBS 0.204468f
C1356 VTAIL.t16 VSUBS 0.204468f
C1357 VTAIL.n46 VSUBS 1.34905f
C1358 VTAIL.n47 VSUBS 2.92691f
C1359 VTAIL.t7 VSUBS 0.204468f
C1360 VTAIL.t1 VSUBS 0.204468f
C1361 VTAIL.n48 VSUBS 1.34906f
C1362 VTAIL.n49 VSUBS 2.9269f
C1363 VTAIL.t3 VSUBS 0.204468f
C1364 VTAIL.t6 VSUBS 0.204468f
C1365 VTAIL.n50 VSUBS 1.34906f
C1366 VTAIL.n51 VSUBS 1.38906f
C1367 VTAIL.n52 VSUBS 0.034384f
C1368 VTAIL.n53 VSUBS 0.032547f
C1369 VTAIL.n54 VSUBS 0.018003f
C1370 VTAIL.n55 VSUBS 0.041338f
C1371 VTAIL.n56 VSUBS 0.017489f
C1372 VTAIL.n57 VSUBS 0.018518f
C1373 VTAIL.n58 VSUBS 0.032547f
C1374 VTAIL.n59 VSUBS 0.017489f
C1375 VTAIL.n60 VSUBS 0.041338f
C1376 VTAIL.n61 VSUBS 0.018518f
C1377 VTAIL.n62 VSUBS 0.032547f
C1378 VTAIL.n63 VSUBS 0.017489f
C1379 VTAIL.n64 VSUBS 0.031003f
C1380 VTAIL.n65 VSUBS 0.031096f
C1381 VTAIL.t0 VSUBS 0.088787f
C1382 VTAIL.n66 VSUBS 0.196852f
C1383 VTAIL.n67 VSUBS 1.02128f
C1384 VTAIL.n68 VSUBS 0.017489f
C1385 VTAIL.n69 VSUBS 0.018518f
C1386 VTAIL.n70 VSUBS 0.041338f
C1387 VTAIL.n71 VSUBS 0.041338f
C1388 VTAIL.n72 VSUBS 0.018518f
C1389 VTAIL.n73 VSUBS 0.017489f
C1390 VTAIL.n74 VSUBS 0.032547f
C1391 VTAIL.n75 VSUBS 0.032547f
C1392 VTAIL.n76 VSUBS 0.017489f
C1393 VTAIL.n77 VSUBS 0.018518f
C1394 VTAIL.n78 VSUBS 0.041338f
C1395 VTAIL.n79 VSUBS 0.041338f
C1396 VTAIL.n80 VSUBS 0.018518f
C1397 VTAIL.n81 VSUBS 0.017489f
C1398 VTAIL.n82 VSUBS 0.032547f
C1399 VTAIL.n83 VSUBS 0.032547f
C1400 VTAIL.n84 VSUBS 0.017489f
C1401 VTAIL.n85 VSUBS 0.018518f
C1402 VTAIL.n86 VSUBS 0.041338f
C1403 VTAIL.n87 VSUBS 0.041338f
C1404 VTAIL.n88 VSUBS 0.095382f
C1405 VTAIL.n89 VSUBS 0.018003f
C1406 VTAIL.n90 VSUBS 0.017489f
C1407 VTAIL.n91 VSUBS 0.081899f
C1408 VTAIL.n92 VSUBS 0.047956f
C1409 VTAIL.n93 VSUBS 0.646338f
C1410 VTAIL.t10 VSUBS 0.204468f
C1411 VTAIL.t12 VSUBS 0.204468f
C1412 VTAIL.n94 VSUBS 1.34906f
C1413 VTAIL.n95 VSUBS 1.24983f
C1414 VTAIL.t15 VSUBS 0.204468f
C1415 VTAIL.t17 VSUBS 0.204468f
C1416 VTAIL.n96 VSUBS 1.34906f
C1417 VTAIL.n97 VSUBS 1.38906f
C1418 VTAIL.n98 VSUBS 0.034384f
C1419 VTAIL.n99 VSUBS 0.032547f
C1420 VTAIL.n100 VSUBS 0.018003f
C1421 VTAIL.n101 VSUBS 0.041338f
C1422 VTAIL.n102 VSUBS 0.017489f
C1423 VTAIL.n103 VSUBS 0.018518f
C1424 VTAIL.n104 VSUBS 0.032547f
C1425 VTAIL.n105 VSUBS 0.017489f
C1426 VTAIL.n106 VSUBS 0.041338f
C1427 VTAIL.n107 VSUBS 0.018518f
C1428 VTAIL.n108 VSUBS 0.032547f
C1429 VTAIL.n109 VSUBS 0.017489f
C1430 VTAIL.n110 VSUBS 0.031003f
C1431 VTAIL.n111 VSUBS 0.031096f
C1432 VTAIL.t18 VSUBS 0.088787f
C1433 VTAIL.n112 VSUBS 0.196852f
C1434 VTAIL.n113 VSUBS 1.02128f
C1435 VTAIL.n114 VSUBS 0.017489f
C1436 VTAIL.n115 VSUBS 0.018518f
C1437 VTAIL.n116 VSUBS 0.041338f
C1438 VTAIL.n117 VSUBS 0.041338f
C1439 VTAIL.n118 VSUBS 0.018518f
C1440 VTAIL.n119 VSUBS 0.017489f
C1441 VTAIL.n120 VSUBS 0.032547f
C1442 VTAIL.n121 VSUBS 0.032547f
C1443 VTAIL.n122 VSUBS 0.017489f
C1444 VTAIL.n123 VSUBS 0.018518f
C1445 VTAIL.n124 VSUBS 0.041338f
C1446 VTAIL.n125 VSUBS 0.041338f
C1447 VTAIL.n126 VSUBS 0.018518f
C1448 VTAIL.n127 VSUBS 0.017489f
C1449 VTAIL.n128 VSUBS 0.032547f
C1450 VTAIL.n129 VSUBS 0.032547f
C1451 VTAIL.n130 VSUBS 0.017489f
C1452 VTAIL.n131 VSUBS 0.018518f
C1453 VTAIL.n132 VSUBS 0.041338f
C1454 VTAIL.n133 VSUBS 0.041338f
C1455 VTAIL.n134 VSUBS 0.095382f
C1456 VTAIL.n135 VSUBS 0.018003f
C1457 VTAIL.n136 VSUBS 0.017489f
C1458 VTAIL.n137 VSUBS 0.081899f
C1459 VTAIL.n138 VSUBS 0.047956f
C1460 VTAIL.n139 VSUBS 1.94641f
C1461 VTAIL.n140 VSUBS 0.034384f
C1462 VTAIL.n141 VSUBS 0.032547f
C1463 VTAIL.n142 VSUBS 0.018003f
C1464 VTAIL.n143 VSUBS 0.041338f
C1465 VTAIL.n144 VSUBS 0.018518f
C1466 VTAIL.n145 VSUBS 0.032547f
C1467 VTAIL.n146 VSUBS 0.017489f
C1468 VTAIL.n147 VSUBS 0.041338f
C1469 VTAIL.n148 VSUBS 0.018518f
C1470 VTAIL.n149 VSUBS 0.032547f
C1471 VTAIL.n150 VSUBS 0.017489f
C1472 VTAIL.n151 VSUBS 0.031003f
C1473 VTAIL.n152 VSUBS 0.031096f
C1474 VTAIL.t2 VSUBS 0.088787f
C1475 VTAIL.n153 VSUBS 0.196852f
C1476 VTAIL.n154 VSUBS 1.02128f
C1477 VTAIL.n155 VSUBS 0.017489f
C1478 VTAIL.n156 VSUBS 0.018518f
C1479 VTAIL.n157 VSUBS 0.041338f
C1480 VTAIL.n158 VSUBS 0.041338f
C1481 VTAIL.n159 VSUBS 0.018518f
C1482 VTAIL.n160 VSUBS 0.017489f
C1483 VTAIL.n161 VSUBS 0.032547f
C1484 VTAIL.n162 VSUBS 0.032547f
C1485 VTAIL.n163 VSUBS 0.017489f
C1486 VTAIL.n164 VSUBS 0.018518f
C1487 VTAIL.n165 VSUBS 0.041338f
C1488 VTAIL.n166 VSUBS 0.041338f
C1489 VTAIL.n167 VSUBS 0.018518f
C1490 VTAIL.n168 VSUBS 0.017489f
C1491 VTAIL.n169 VSUBS 0.032547f
C1492 VTAIL.n170 VSUBS 0.032547f
C1493 VTAIL.n171 VSUBS 0.017489f
C1494 VTAIL.n172 VSUBS 0.017489f
C1495 VTAIL.n173 VSUBS 0.018518f
C1496 VTAIL.n174 VSUBS 0.041338f
C1497 VTAIL.n175 VSUBS 0.041338f
C1498 VTAIL.n176 VSUBS 0.095382f
C1499 VTAIL.n177 VSUBS 0.018003f
C1500 VTAIL.n178 VSUBS 0.017489f
C1501 VTAIL.n179 VSUBS 0.081899f
C1502 VTAIL.n180 VSUBS 0.047956f
C1503 VTAIL.n181 VSUBS 1.94641f
C1504 VTAIL.t8 VSUBS 0.204468f
C1505 VTAIL.t5 VSUBS 0.204468f
C1506 VTAIL.n182 VSUBS 1.34905f
C1507 VTAIL.n183 VSUBS 1.10022f
C1508 VP.t3 VSUBS 2.45274f
C1509 VP.n0 VSUBS 0.996807f
C1510 VP.n1 VSUBS 0.029924f
C1511 VP.n2 VSUBS 0.05932f
C1512 VP.n3 VSUBS 0.029924f
C1513 VP.n4 VSUBS 0.05577f
C1514 VP.n5 VSUBS 0.029924f
C1515 VP.t6 VSUBS 2.45274f
C1516 VP.n6 VSUBS 0.05577f
C1517 VP.n7 VSUBS 0.029924f
C1518 VP.n8 VSUBS 0.05577f
C1519 VP.n9 VSUBS 0.029924f
C1520 VP.t9 VSUBS 2.45274f
C1521 VP.n10 VSUBS 0.05577f
C1522 VP.n11 VSUBS 0.029924f
C1523 VP.n12 VSUBS 0.05577f
C1524 VP.n13 VSUBS 0.029924f
C1525 VP.t1 VSUBS 2.45274f
C1526 VP.n14 VSUBS 0.05577f
C1527 VP.n15 VSUBS 0.029924f
C1528 VP.n16 VSUBS 0.05577f
C1529 VP.n17 VSUBS 0.048296f
C1530 VP.t4 VSUBS 2.45274f
C1531 VP.t8 VSUBS 2.45274f
C1532 VP.n18 VSUBS 0.996807f
C1533 VP.n19 VSUBS 0.029924f
C1534 VP.n20 VSUBS 0.05932f
C1535 VP.n21 VSUBS 0.029924f
C1536 VP.n22 VSUBS 0.05577f
C1537 VP.n23 VSUBS 0.029924f
C1538 VP.t5 VSUBS 2.45274f
C1539 VP.n24 VSUBS 0.05577f
C1540 VP.n25 VSUBS 0.029924f
C1541 VP.n26 VSUBS 0.05577f
C1542 VP.n27 VSUBS 0.029924f
C1543 VP.t0 VSUBS 2.45274f
C1544 VP.n28 VSUBS 0.05577f
C1545 VP.n29 VSUBS 0.029924f
C1546 VP.n30 VSUBS 0.05577f
C1547 VP.t2 VSUBS 2.90125f
C1548 VP.n31 VSUBS 0.950882f
C1549 VP.t7 VSUBS 2.45274f
C1550 VP.n32 VSUBS 0.998911f
C1551 VP.n33 VSUBS 0.051365f
C1552 VP.n34 VSUBS 0.385136f
C1553 VP.n35 VSUBS 0.029924f
C1554 VP.n36 VSUBS 0.029924f
C1555 VP.n37 VSUBS 0.05577f
C1556 VP.n38 VSUBS 0.036598f
C1557 VP.n39 VSUBS 0.050774f
C1558 VP.n40 VSUBS 0.029924f
C1559 VP.n41 VSUBS 0.029924f
C1560 VP.n42 VSUBS 0.029924f
C1561 VP.n43 VSUBS 0.05577f
C1562 VP.n44 VSUBS 0.042003f
C1563 VP.n45 VSUBS 0.880895f
C1564 VP.n46 VSUBS 0.042003f
C1565 VP.n47 VSUBS 0.029924f
C1566 VP.n48 VSUBS 0.029924f
C1567 VP.n49 VSUBS 0.029924f
C1568 VP.n50 VSUBS 0.05577f
C1569 VP.n51 VSUBS 0.050774f
C1570 VP.n52 VSUBS 0.036598f
C1571 VP.n53 VSUBS 0.029924f
C1572 VP.n54 VSUBS 0.029924f
C1573 VP.n55 VSUBS 0.029924f
C1574 VP.n56 VSUBS 0.05577f
C1575 VP.n57 VSUBS 0.051365f
C1576 VP.n58 VSUBS 0.880895f
C1577 VP.n59 VSUBS 0.032642f
C1578 VP.n60 VSUBS 0.029924f
C1579 VP.n61 VSUBS 0.029924f
C1580 VP.n62 VSUBS 0.029924f
C1581 VP.n63 VSUBS 0.05577f
C1582 VP.n64 VSUBS 0.05962f
C1583 VP.n65 VSUBS 0.024201f
C1584 VP.n66 VSUBS 0.029924f
C1585 VP.n67 VSUBS 0.029924f
C1586 VP.n68 VSUBS 0.029924f
C1587 VP.n69 VSUBS 0.05577f
C1588 VP.n70 VSUBS 0.05577f
C1589 VP.n71 VSUBS 0.033192f
C1590 VP.n72 VSUBS 0.048296f
C1591 VP.n73 VSUBS 2.05855f
C1592 VP.n74 VSUBS 2.07746f
C1593 VP.n75 VSUBS 0.996807f
C1594 VP.n76 VSUBS 0.033192f
C1595 VP.n77 VSUBS 0.05577f
C1596 VP.n78 VSUBS 0.029924f
C1597 VP.n79 VSUBS 0.029924f
C1598 VP.n80 VSUBS 0.029924f
C1599 VP.n81 VSUBS 0.05932f
C1600 VP.n82 VSUBS 0.024201f
C1601 VP.n83 VSUBS 0.05962f
C1602 VP.n84 VSUBS 0.029924f
C1603 VP.n85 VSUBS 0.029924f
C1604 VP.n86 VSUBS 0.029924f
C1605 VP.n87 VSUBS 0.05577f
C1606 VP.n88 VSUBS 0.032642f
C1607 VP.n89 VSUBS 0.880895f
C1608 VP.n90 VSUBS 0.051365f
C1609 VP.n91 VSUBS 0.029924f
C1610 VP.n92 VSUBS 0.029924f
C1611 VP.n93 VSUBS 0.029924f
C1612 VP.n94 VSUBS 0.05577f
C1613 VP.n95 VSUBS 0.036598f
C1614 VP.n96 VSUBS 0.050774f
C1615 VP.n97 VSUBS 0.029924f
C1616 VP.n98 VSUBS 0.029924f
C1617 VP.n99 VSUBS 0.029924f
C1618 VP.n100 VSUBS 0.05577f
C1619 VP.n101 VSUBS 0.042003f
C1620 VP.n102 VSUBS 0.880895f
C1621 VP.n103 VSUBS 0.042003f
C1622 VP.n104 VSUBS 0.029924f
C1623 VP.n105 VSUBS 0.029924f
C1624 VP.n106 VSUBS 0.029924f
C1625 VP.n107 VSUBS 0.05577f
C1626 VP.n108 VSUBS 0.050774f
C1627 VP.n109 VSUBS 0.036598f
C1628 VP.n110 VSUBS 0.029924f
C1629 VP.n111 VSUBS 0.029924f
C1630 VP.n112 VSUBS 0.029924f
C1631 VP.n113 VSUBS 0.05577f
C1632 VP.n114 VSUBS 0.051365f
C1633 VP.n115 VSUBS 0.880895f
C1634 VP.n116 VSUBS 0.032642f
C1635 VP.n117 VSUBS 0.029924f
C1636 VP.n118 VSUBS 0.029924f
C1637 VP.n119 VSUBS 0.029924f
C1638 VP.n120 VSUBS 0.05577f
C1639 VP.n121 VSUBS 0.05962f
C1640 VP.n122 VSUBS 0.024201f
C1641 VP.n123 VSUBS 0.029924f
C1642 VP.n124 VSUBS 0.029924f
C1643 VP.n125 VSUBS 0.029924f
C1644 VP.n126 VSUBS 0.05577f
C1645 VP.n127 VSUBS 0.05577f
C1646 VP.n128 VSUBS 0.033192f
C1647 VP.n129 VSUBS 0.048296f
C1648 VP.n130 VSUBS 0.091186f
.ends

