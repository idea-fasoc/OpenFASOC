* NGSPICE file created from diff_pair_sample_1274.ext - technology: sky130A

.subckt diff_pair_sample_1274 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t10 w_n4700_n3898# sky130_fd_pr__pfet_01v8 ad=2.41725 pd=14.98 as=5.7135 ps=30.08 w=14.65 l=3.4
X1 VDD1.t6 VP.t1 VTAIL.t9 w_n4700_n3898# sky130_fd_pr__pfet_01v8 ad=2.41725 pd=14.98 as=2.41725 ps=14.98 w=14.65 l=3.4
X2 B.t11 B.t9 B.t10 w_n4700_n3898# sky130_fd_pr__pfet_01v8 ad=5.7135 pd=30.08 as=0 ps=0 w=14.65 l=3.4
X3 VTAIL.t1 VN.t0 VDD2.t7 w_n4700_n3898# sky130_fd_pr__pfet_01v8 ad=5.7135 pd=30.08 as=2.41725 ps=14.98 w=14.65 l=3.4
X4 VDD1.t5 VP.t2 VTAIL.t15 w_n4700_n3898# sky130_fd_pr__pfet_01v8 ad=2.41725 pd=14.98 as=5.7135 ps=30.08 w=14.65 l=3.4
X5 VTAIL.t3 VN.t1 VDD2.t6 w_n4700_n3898# sky130_fd_pr__pfet_01v8 ad=5.7135 pd=30.08 as=2.41725 ps=14.98 w=14.65 l=3.4
X6 B.t8 B.t6 B.t7 w_n4700_n3898# sky130_fd_pr__pfet_01v8 ad=5.7135 pd=30.08 as=0 ps=0 w=14.65 l=3.4
X7 VTAIL.t7 VN.t2 VDD2.t5 w_n4700_n3898# sky130_fd_pr__pfet_01v8 ad=2.41725 pd=14.98 as=2.41725 ps=14.98 w=14.65 l=3.4
X8 VTAIL.t14 VP.t3 VDD1.t4 w_n4700_n3898# sky130_fd_pr__pfet_01v8 ad=5.7135 pd=30.08 as=2.41725 ps=14.98 w=14.65 l=3.4
X9 VTAIL.t0 VN.t3 VDD2.t4 w_n4700_n3898# sky130_fd_pr__pfet_01v8 ad=2.41725 pd=14.98 as=2.41725 ps=14.98 w=14.65 l=3.4
X10 VDD2.t3 VN.t4 VTAIL.t5 w_n4700_n3898# sky130_fd_pr__pfet_01v8 ad=2.41725 pd=14.98 as=5.7135 ps=30.08 w=14.65 l=3.4
X11 VTAIL.t13 VP.t4 VDD1.t3 w_n4700_n3898# sky130_fd_pr__pfet_01v8 ad=2.41725 pd=14.98 as=2.41725 ps=14.98 w=14.65 l=3.4
X12 VDD1.t2 VP.t5 VTAIL.t8 w_n4700_n3898# sky130_fd_pr__pfet_01v8 ad=2.41725 pd=14.98 as=2.41725 ps=14.98 w=14.65 l=3.4
X13 VTAIL.t11 VP.t6 VDD1.t1 w_n4700_n3898# sky130_fd_pr__pfet_01v8 ad=2.41725 pd=14.98 as=2.41725 ps=14.98 w=14.65 l=3.4
X14 VDD2.t2 VN.t5 VTAIL.t6 w_n4700_n3898# sky130_fd_pr__pfet_01v8 ad=2.41725 pd=14.98 as=2.41725 ps=14.98 w=14.65 l=3.4
X15 B.t5 B.t3 B.t4 w_n4700_n3898# sky130_fd_pr__pfet_01v8 ad=5.7135 pd=30.08 as=0 ps=0 w=14.65 l=3.4
X16 VTAIL.t12 VP.t7 VDD1.t0 w_n4700_n3898# sky130_fd_pr__pfet_01v8 ad=5.7135 pd=30.08 as=2.41725 ps=14.98 w=14.65 l=3.4
X17 VDD2.t1 VN.t6 VTAIL.t4 w_n4700_n3898# sky130_fd_pr__pfet_01v8 ad=2.41725 pd=14.98 as=2.41725 ps=14.98 w=14.65 l=3.4
X18 B.t2 B.t0 B.t1 w_n4700_n3898# sky130_fd_pr__pfet_01v8 ad=5.7135 pd=30.08 as=0 ps=0 w=14.65 l=3.4
X19 VDD2.t0 VN.t7 VTAIL.t2 w_n4700_n3898# sky130_fd_pr__pfet_01v8 ad=2.41725 pd=14.98 as=5.7135 ps=30.08 w=14.65 l=3.4
R0 VP.n24 VP.n21 161.3
R1 VP.n26 VP.n25 161.3
R2 VP.n27 VP.n20 161.3
R3 VP.n29 VP.n28 161.3
R4 VP.n30 VP.n19 161.3
R5 VP.n32 VP.n31 161.3
R6 VP.n33 VP.n18 161.3
R7 VP.n35 VP.n34 161.3
R8 VP.n37 VP.n36 161.3
R9 VP.n38 VP.n16 161.3
R10 VP.n40 VP.n39 161.3
R11 VP.n41 VP.n15 161.3
R12 VP.n43 VP.n42 161.3
R13 VP.n44 VP.n14 161.3
R14 VP.n46 VP.n45 161.3
R15 VP.n83 VP.n82 161.3
R16 VP.n81 VP.n1 161.3
R17 VP.n80 VP.n79 161.3
R18 VP.n78 VP.n2 161.3
R19 VP.n77 VP.n76 161.3
R20 VP.n75 VP.n3 161.3
R21 VP.n74 VP.n73 161.3
R22 VP.n72 VP.n71 161.3
R23 VP.n70 VP.n5 161.3
R24 VP.n69 VP.n68 161.3
R25 VP.n67 VP.n6 161.3
R26 VP.n66 VP.n65 161.3
R27 VP.n64 VP.n7 161.3
R28 VP.n63 VP.n62 161.3
R29 VP.n61 VP.n8 161.3
R30 VP.n60 VP.n59 161.3
R31 VP.n57 VP.n9 161.3
R32 VP.n56 VP.n55 161.3
R33 VP.n54 VP.n10 161.3
R34 VP.n53 VP.n52 161.3
R35 VP.n51 VP.n11 161.3
R36 VP.n50 VP.n49 161.3
R37 VP.n23 VP.t7 136.925
R38 VP.n12 VP.t3 103.844
R39 VP.n58 VP.t1 103.844
R40 VP.n4 VP.t6 103.844
R41 VP.n0 VP.t0 103.844
R42 VP.n13 VP.t2 103.844
R43 VP.n17 VP.t4 103.844
R44 VP.n22 VP.t5 103.844
R45 VP.n48 VP.n12 73.1852
R46 VP.n84 VP.n0 73.1852
R47 VP.n47 VP.n13 73.1852
R48 VP.n23 VP.n22 68.9427
R49 VP.n48 VP.n47 56.8175
R50 VP.n65 VP.n6 56.5193
R51 VP.n28 VP.n19 56.5193
R52 VP.n56 VP.n10 42.4359
R53 VP.n76 VP.n2 42.4359
R54 VP.n39 VP.n15 42.4359
R55 VP.n52 VP.n10 38.5509
R56 VP.n80 VP.n2 38.5509
R57 VP.n43 VP.n15 38.5509
R58 VP.n51 VP.n50 24.4675
R59 VP.n52 VP.n51 24.4675
R60 VP.n57 VP.n56 24.4675
R61 VP.n59 VP.n57 24.4675
R62 VP.n63 VP.n8 24.4675
R63 VP.n64 VP.n63 24.4675
R64 VP.n65 VP.n64 24.4675
R65 VP.n69 VP.n6 24.4675
R66 VP.n70 VP.n69 24.4675
R67 VP.n71 VP.n70 24.4675
R68 VP.n75 VP.n74 24.4675
R69 VP.n76 VP.n75 24.4675
R70 VP.n81 VP.n80 24.4675
R71 VP.n82 VP.n81 24.4675
R72 VP.n44 VP.n43 24.4675
R73 VP.n45 VP.n44 24.4675
R74 VP.n32 VP.n19 24.4675
R75 VP.n33 VP.n32 24.4675
R76 VP.n34 VP.n33 24.4675
R77 VP.n38 VP.n37 24.4675
R78 VP.n39 VP.n38 24.4675
R79 VP.n26 VP.n21 24.4675
R80 VP.n27 VP.n26 24.4675
R81 VP.n28 VP.n27 24.4675
R82 VP.n59 VP.n58 18.8401
R83 VP.n74 VP.n4 18.8401
R84 VP.n37 VP.n17 18.8401
R85 VP.n50 VP.n12 16.8827
R86 VP.n82 VP.n0 16.8827
R87 VP.n45 VP.n13 16.8827
R88 VP.n58 VP.n8 5.62791
R89 VP.n71 VP.n4 5.62791
R90 VP.n34 VP.n17 5.62791
R91 VP.n22 VP.n21 5.62791
R92 VP.n24 VP.n23 4.05577
R93 VP.n47 VP.n46 0.354971
R94 VP.n49 VP.n48 0.354971
R95 VP.n84 VP.n83 0.354971
R96 VP VP.n84 0.26696
R97 VP.n25 VP.n24 0.189894
R98 VP.n25 VP.n20 0.189894
R99 VP.n29 VP.n20 0.189894
R100 VP.n30 VP.n29 0.189894
R101 VP.n31 VP.n30 0.189894
R102 VP.n31 VP.n18 0.189894
R103 VP.n35 VP.n18 0.189894
R104 VP.n36 VP.n35 0.189894
R105 VP.n36 VP.n16 0.189894
R106 VP.n40 VP.n16 0.189894
R107 VP.n41 VP.n40 0.189894
R108 VP.n42 VP.n41 0.189894
R109 VP.n42 VP.n14 0.189894
R110 VP.n46 VP.n14 0.189894
R111 VP.n49 VP.n11 0.189894
R112 VP.n53 VP.n11 0.189894
R113 VP.n54 VP.n53 0.189894
R114 VP.n55 VP.n54 0.189894
R115 VP.n55 VP.n9 0.189894
R116 VP.n60 VP.n9 0.189894
R117 VP.n61 VP.n60 0.189894
R118 VP.n62 VP.n61 0.189894
R119 VP.n62 VP.n7 0.189894
R120 VP.n66 VP.n7 0.189894
R121 VP.n67 VP.n66 0.189894
R122 VP.n68 VP.n67 0.189894
R123 VP.n68 VP.n5 0.189894
R124 VP.n72 VP.n5 0.189894
R125 VP.n73 VP.n72 0.189894
R126 VP.n73 VP.n3 0.189894
R127 VP.n77 VP.n3 0.189894
R128 VP.n78 VP.n77 0.189894
R129 VP.n79 VP.n78 0.189894
R130 VP.n79 VP.n1 0.189894
R131 VP.n83 VP.n1 0.189894
R132 VTAIL.n658 VTAIL.n582 756.745
R133 VTAIL.n78 VTAIL.n2 756.745
R134 VTAIL.n160 VTAIL.n84 756.745
R135 VTAIL.n244 VTAIL.n168 756.745
R136 VTAIL.n576 VTAIL.n500 756.745
R137 VTAIL.n492 VTAIL.n416 756.745
R138 VTAIL.n410 VTAIL.n334 756.745
R139 VTAIL.n326 VTAIL.n250 756.745
R140 VTAIL.n609 VTAIL.n608 585
R141 VTAIL.n606 VTAIL.n605 585
R142 VTAIL.n615 VTAIL.n614 585
R143 VTAIL.n617 VTAIL.n616 585
R144 VTAIL.n602 VTAIL.n601 585
R145 VTAIL.n623 VTAIL.n622 585
R146 VTAIL.n625 VTAIL.n624 585
R147 VTAIL.n598 VTAIL.n597 585
R148 VTAIL.n631 VTAIL.n630 585
R149 VTAIL.n633 VTAIL.n632 585
R150 VTAIL.n594 VTAIL.n593 585
R151 VTAIL.n639 VTAIL.n638 585
R152 VTAIL.n641 VTAIL.n640 585
R153 VTAIL.n590 VTAIL.n589 585
R154 VTAIL.n647 VTAIL.n646 585
R155 VTAIL.n650 VTAIL.n649 585
R156 VTAIL.n648 VTAIL.n586 585
R157 VTAIL.n655 VTAIL.n585 585
R158 VTAIL.n657 VTAIL.n656 585
R159 VTAIL.n659 VTAIL.n658 585
R160 VTAIL.n29 VTAIL.n28 585
R161 VTAIL.n26 VTAIL.n25 585
R162 VTAIL.n35 VTAIL.n34 585
R163 VTAIL.n37 VTAIL.n36 585
R164 VTAIL.n22 VTAIL.n21 585
R165 VTAIL.n43 VTAIL.n42 585
R166 VTAIL.n45 VTAIL.n44 585
R167 VTAIL.n18 VTAIL.n17 585
R168 VTAIL.n51 VTAIL.n50 585
R169 VTAIL.n53 VTAIL.n52 585
R170 VTAIL.n14 VTAIL.n13 585
R171 VTAIL.n59 VTAIL.n58 585
R172 VTAIL.n61 VTAIL.n60 585
R173 VTAIL.n10 VTAIL.n9 585
R174 VTAIL.n67 VTAIL.n66 585
R175 VTAIL.n70 VTAIL.n69 585
R176 VTAIL.n68 VTAIL.n6 585
R177 VTAIL.n75 VTAIL.n5 585
R178 VTAIL.n77 VTAIL.n76 585
R179 VTAIL.n79 VTAIL.n78 585
R180 VTAIL.n111 VTAIL.n110 585
R181 VTAIL.n108 VTAIL.n107 585
R182 VTAIL.n117 VTAIL.n116 585
R183 VTAIL.n119 VTAIL.n118 585
R184 VTAIL.n104 VTAIL.n103 585
R185 VTAIL.n125 VTAIL.n124 585
R186 VTAIL.n127 VTAIL.n126 585
R187 VTAIL.n100 VTAIL.n99 585
R188 VTAIL.n133 VTAIL.n132 585
R189 VTAIL.n135 VTAIL.n134 585
R190 VTAIL.n96 VTAIL.n95 585
R191 VTAIL.n141 VTAIL.n140 585
R192 VTAIL.n143 VTAIL.n142 585
R193 VTAIL.n92 VTAIL.n91 585
R194 VTAIL.n149 VTAIL.n148 585
R195 VTAIL.n152 VTAIL.n151 585
R196 VTAIL.n150 VTAIL.n88 585
R197 VTAIL.n157 VTAIL.n87 585
R198 VTAIL.n159 VTAIL.n158 585
R199 VTAIL.n161 VTAIL.n160 585
R200 VTAIL.n195 VTAIL.n194 585
R201 VTAIL.n192 VTAIL.n191 585
R202 VTAIL.n201 VTAIL.n200 585
R203 VTAIL.n203 VTAIL.n202 585
R204 VTAIL.n188 VTAIL.n187 585
R205 VTAIL.n209 VTAIL.n208 585
R206 VTAIL.n211 VTAIL.n210 585
R207 VTAIL.n184 VTAIL.n183 585
R208 VTAIL.n217 VTAIL.n216 585
R209 VTAIL.n219 VTAIL.n218 585
R210 VTAIL.n180 VTAIL.n179 585
R211 VTAIL.n225 VTAIL.n224 585
R212 VTAIL.n227 VTAIL.n226 585
R213 VTAIL.n176 VTAIL.n175 585
R214 VTAIL.n233 VTAIL.n232 585
R215 VTAIL.n236 VTAIL.n235 585
R216 VTAIL.n234 VTAIL.n172 585
R217 VTAIL.n241 VTAIL.n171 585
R218 VTAIL.n243 VTAIL.n242 585
R219 VTAIL.n245 VTAIL.n244 585
R220 VTAIL.n577 VTAIL.n576 585
R221 VTAIL.n575 VTAIL.n574 585
R222 VTAIL.n573 VTAIL.n503 585
R223 VTAIL.n507 VTAIL.n504 585
R224 VTAIL.n568 VTAIL.n567 585
R225 VTAIL.n566 VTAIL.n565 585
R226 VTAIL.n509 VTAIL.n508 585
R227 VTAIL.n560 VTAIL.n559 585
R228 VTAIL.n558 VTAIL.n557 585
R229 VTAIL.n513 VTAIL.n512 585
R230 VTAIL.n552 VTAIL.n551 585
R231 VTAIL.n550 VTAIL.n549 585
R232 VTAIL.n517 VTAIL.n516 585
R233 VTAIL.n544 VTAIL.n543 585
R234 VTAIL.n542 VTAIL.n541 585
R235 VTAIL.n521 VTAIL.n520 585
R236 VTAIL.n536 VTAIL.n535 585
R237 VTAIL.n534 VTAIL.n533 585
R238 VTAIL.n525 VTAIL.n524 585
R239 VTAIL.n528 VTAIL.n527 585
R240 VTAIL.n493 VTAIL.n492 585
R241 VTAIL.n491 VTAIL.n490 585
R242 VTAIL.n489 VTAIL.n419 585
R243 VTAIL.n423 VTAIL.n420 585
R244 VTAIL.n484 VTAIL.n483 585
R245 VTAIL.n482 VTAIL.n481 585
R246 VTAIL.n425 VTAIL.n424 585
R247 VTAIL.n476 VTAIL.n475 585
R248 VTAIL.n474 VTAIL.n473 585
R249 VTAIL.n429 VTAIL.n428 585
R250 VTAIL.n468 VTAIL.n467 585
R251 VTAIL.n466 VTAIL.n465 585
R252 VTAIL.n433 VTAIL.n432 585
R253 VTAIL.n460 VTAIL.n459 585
R254 VTAIL.n458 VTAIL.n457 585
R255 VTAIL.n437 VTAIL.n436 585
R256 VTAIL.n452 VTAIL.n451 585
R257 VTAIL.n450 VTAIL.n449 585
R258 VTAIL.n441 VTAIL.n440 585
R259 VTAIL.n444 VTAIL.n443 585
R260 VTAIL.n411 VTAIL.n410 585
R261 VTAIL.n409 VTAIL.n408 585
R262 VTAIL.n407 VTAIL.n337 585
R263 VTAIL.n341 VTAIL.n338 585
R264 VTAIL.n402 VTAIL.n401 585
R265 VTAIL.n400 VTAIL.n399 585
R266 VTAIL.n343 VTAIL.n342 585
R267 VTAIL.n394 VTAIL.n393 585
R268 VTAIL.n392 VTAIL.n391 585
R269 VTAIL.n347 VTAIL.n346 585
R270 VTAIL.n386 VTAIL.n385 585
R271 VTAIL.n384 VTAIL.n383 585
R272 VTAIL.n351 VTAIL.n350 585
R273 VTAIL.n378 VTAIL.n377 585
R274 VTAIL.n376 VTAIL.n375 585
R275 VTAIL.n355 VTAIL.n354 585
R276 VTAIL.n370 VTAIL.n369 585
R277 VTAIL.n368 VTAIL.n367 585
R278 VTAIL.n359 VTAIL.n358 585
R279 VTAIL.n362 VTAIL.n361 585
R280 VTAIL.n327 VTAIL.n326 585
R281 VTAIL.n325 VTAIL.n324 585
R282 VTAIL.n323 VTAIL.n253 585
R283 VTAIL.n257 VTAIL.n254 585
R284 VTAIL.n318 VTAIL.n317 585
R285 VTAIL.n316 VTAIL.n315 585
R286 VTAIL.n259 VTAIL.n258 585
R287 VTAIL.n310 VTAIL.n309 585
R288 VTAIL.n308 VTAIL.n307 585
R289 VTAIL.n263 VTAIL.n262 585
R290 VTAIL.n302 VTAIL.n301 585
R291 VTAIL.n300 VTAIL.n299 585
R292 VTAIL.n267 VTAIL.n266 585
R293 VTAIL.n294 VTAIL.n293 585
R294 VTAIL.n292 VTAIL.n291 585
R295 VTAIL.n271 VTAIL.n270 585
R296 VTAIL.n286 VTAIL.n285 585
R297 VTAIL.n284 VTAIL.n283 585
R298 VTAIL.n275 VTAIL.n274 585
R299 VTAIL.n278 VTAIL.n277 585
R300 VTAIL.t15 VTAIL.n526 327.466
R301 VTAIL.t12 VTAIL.n442 327.466
R302 VTAIL.t5 VTAIL.n360 327.466
R303 VTAIL.t3 VTAIL.n276 327.466
R304 VTAIL.t2 VTAIL.n607 327.466
R305 VTAIL.t1 VTAIL.n27 327.466
R306 VTAIL.t10 VTAIL.n109 327.466
R307 VTAIL.t14 VTAIL.n193 327.466
R308 VTAIL.n608 VTAIL.n605 171.744
R309 VTAIL.n615 VTAIL.n605 171.744
R310 VTAIL.n616 VTAIL.n615 171.744
R311 VTAIL.n616 VTAIL.n601 171.744
R312 VTAIL.n623 VTAIL.n601 171.744
R313 VTAIL.n624 VTAIL.n623 171.744
R314 VTAIL.n624 VTAIL.n597 171.744
R315 VTAIL.n631 VTAIL.n597 171.744
R316 VTAIL.n632 VTAIL.n631 171.744
R317 VTAIL.n632 VTAIL.n593 171.744
R318 VTAIL.n639 VTAIL.n593 171.744
R319 VTAIL.n640 VTAIL.n639 171.744
R320 VTAIL.n640 VTAIL.n589 171.744
R321 VTAIL.n647 VTAIL.n589 171.744
R322 VTAIL.n649 VTAIL.n647 171.744
R323 VTAIL.n649 VTAIL.n648 171.744
R324 VTAIL.n648 VTAIL.n585 171.744
R325 VTAIL.n657 VTAIL.n585 171.744
R326 VTAIL.n658 VTAIL.n657 171.744
R327 VTAIL.n28 VTAIL.n25 171.744
R328 VTAIL.n35 VTAIL.n25 171.744
R329 VTAIL.n36 VTAIL.n35 171.744
R330 VTAIL.n36 VTAIL.n21 171.744
R331 VTAIL.n43 VTAIL.n21 171.744
R332 VTAIL.n44 VTAIL.n43 171.744
R333 VTAIL.n44 VTAIL.n17 171.744
R334 VTAIL.n51 VTAIL.n17 171.744
R335 VTAIL.n52 VTAIL.n51 171.744
R336 VTAIL.n52 VTAIL.n13 171.744
R337 VTAIL.n59 VTAIL.n13 171.744
R338 VTAIL.n60 VTAIL.n59 171.744
R339 VTAIL.n60 VTAIL.n9 171.744
R340 VTAIL.n67 VTAIL.n9 171.744
R341 VTAIL.n69 VTAIL.n67 171.744
R342 VTAIL.n69 VTAIL.n68 171.744
R343 VTAIL.n68 VTAIL.n5 171.744
R344 VTAIL.n77 VTAIL.n5 171.744
R345 VTAIL.n78 VTAIL.n77 171.744
R346 VTAIL.n110 VTAIL.n107 171.744
R347 VTAIL.n117 VTAIL.n107 171.744
R348 VTAIL.n118 VTAIL.n117 171.744
R349 VTAIL.n118 VTAIL.n103 171.744
R350 VTAIL.n125 VTAIL.n103 171.744
R351 VTAIL.n126 VTAIL.n125 171.744
R352 VTAIL.n126 VTAIL.n99 171.744
R353 VTAIL.n133 VTAIL.n99 171.744
R354 VTAIL.n134 VTAIL.n133 171.744
R355 VTAIL.n134 VTAIL.n95 171.744
R356 VTAIL.n141 VTAIL.n95 171.744
R357 VTAIL.n142 VTAIL.n141 171.744
R358 VTAIL.n142 VTAIL.n91 171.744
R359 VTAIL.n149 VTAIL.n91 171.744
R360 VTAIL.n151 VTAIL.n149 171.744
R361 VTAIL.n151 VTAIL.n150 171.744
R362 VTAIL.n150 VTAIL.n87 171.744
R363 VTAIL.n159 VTAIL.n87 171.744
R364 VTAIL.n160 VTAIL.n159 171.744
R365 VTAIL.n194 VTAIL.n191 171.744
R366 VTAIL.n201 VTAIL.n191 171.744
R367 VTAIL.n202 VTAIL.n201 171.744
R368 VTAIL.n202 VTAIL.n187 171.744
R369 VTAIL.n209 VTAIL.n187 171.744
R370 VTAIL.n210 VTAIL.n209 171.744
R371 VTAIL.n210 VTAIL.n183 171.744
R372 VTAIL.n217 VTAIL.n183 171.744
R373 VTAIL.n218 VTAIL.n217 171.744
R374 VTAIL.n218 VTAIL.n179 171.744
R375 VTAIL.n225 VTAIL.n179 171.744
R376 VTAIL.n226 VTAIL.n225 171.744
R377 VTAIL.n226 VTAIL.n175 171.744
R378 VTAIL.n233 VTAIL.n175 171.744
R379 VTAIL.n235 VTAIL.n233 171.744
R380 VTAIL.n235 VTAIL.n234 171.744
R381 VTAIL.n234 VTAIL.n171 171.744
R382 VTAIL.n243 VTAIL.n171 171.744
R383 VTAIL.n244 VTAIL.n243 171.744
R384 VTAIL.n576 VTAIL.n575 171.744
R385 VTAIL.n575 VTAIL.n503 171.744
R386 VTAIL.n507 VTAIL.n503 171.744
R387 VTAIL.n567 VTAIL.n507 171.744
R388 VTAIL.n567 VTAIL.n566 171.744
R389 VTAIL.n566 VTAIL.n508 171.744
R390 VTAIL.n559 VTAIL.n508 171.744
R391 VTAIL.n559 VTAIL.n558 171.744
R392 VTAIL.n558 VTAIL.n512 171.744
R393 VTAIL.n551 VTAIL.n512 171.744
R394 VTAIL.n551 VTAIL.n550 171.744
R395 VTAIL.n550 VTAIL.n516 171.744
R396 VTAIL.n543 VTAIL.n516 171.744
R397 VTAIL.n543 VTAIL.n542 171.744
R398 VTAIL.n542 VTAIL.n520 171.744
R399 VTAIL.n535 VTAIL.n520 171.744
R400 VTAIL.n535 VTAIL.n534 171.744
R401 VTAIL.n534 VTAIL.n524 171.744
R402 VTAIL.n527 VTAIL.n524 171.744
R403 VTAIL.n492 VTAIL.n491 171.744
R404 VTAIL.n491 VTAIL.n419 171.744
R405 VTAIL.n423 VTAIL.n419 171.744
R406 VTAIL.n483 VTAIL.n423 171.744
R407 VTAIL.n483 VTAIL.n482 171.744
R408 VTAIL.n482 VTAIL.n424 171.744
R409 VTAIL.n475 VTAIL.n424 171.744
R410 VTAIL.n475 VTAIL.n474 171.744
R411 VTAIL.n474 VTAIL.n428 171.744
R412 VTAIL.n467 VTAIL.n428 171.744
R413 VTAIL.n467 VTAIL.n466 171.744
R414 VTAIL.n466 VTAIL.n432 171.744
R415 VTAIL.n459 VTAIL.n432 171.744
R416 VTAIL.n459 VTAIL.n458 171.744
R417 VTAIL.n458 VTAIL.n436 171.744
R418 VTAIL.n451 VTAIL.n436 171.744
R419 VTAIL.n451 VTAIL.n450 171.744
R420 VTAIL.n450 VTAIL.n440 171.744
R421 VTAIL.n443 VTAIL.n440 171.744
R422 VTAIL.n410 VTAIL.n409 171.744
R423 VTAIL.n409 VTAIL.n337 171.744
R424 VTAIL.n341 VTAIL.n337 171.744
R425 VTAIL.n401 VTAIL.n341 171.744
R426 VTAIL.n401 VTAIL.n400 171.744
R427 VTAIL.n400 VTAIL.n342 171.744
R428 VTAIL.n393 VTAIL.n342 171.744
R429 VTAIL.n393 VTAIL.n392 171.744
R430 VTAIL.n392 VTAIL.n346 171.744
R431 VTAIL.n385 VTAIL.n346 171.744
R432 VTAIL.n385 VTAIL.n384 171.744
R433 VTAIL.n384 VTAIL.n350 171.744
R434 VTAIL.n377 VTAIL.n350 171.744
R435 VTAIL.n377 VTAIL.n376 171.744
R436 VTAIL.n376 VTAIL.n354 171.744
R437 VTAIL.n369 VTAIL.n354 171.744
R438 VTAIL.n369 VTAIL.n368 171.744
R439 VTAIL.n368 VTAIL.n358 171.744
R440 VTAIL.n361 VTAIL.n358 171.744
R441 VTAIL.n326 VTAIL.n325 171.744
R442 VTAIL.n325 VTAIL.n253 171.744
R443 VTAIL.n257 VTAIL.n253 171.744
R444 VTAIL.n317 VTAIL.n257 171.744
R445 VTAIL.n317 VTAIL.n316 171.744
R446 VTAIL.n316 VTAIL.n258 171.744
R447 VTAIL.n309 VTAIL.n258 171.744
R448 VTAIL.n309 VTAIL.n308 171.744
R449 VTAIL.n308 VTAIL.n262 171.744
R450 VTAIL.n301 VTAIL.n262 171.744
R451 VTAIL.n301 VTAIL.n300 171.744
R452 VTAIL.n300 VTAIL.n266 171.744
R453 VTAIL.n293 VTAIL.n266 171.744
R454 VTAIL.n293 VTAIL.n292 171.744
R455 VTAIL.n292 VTAIL.n270 171.744
R456 VTAIL.n285 VTAIL.n270 171.744
R457 VTAIL.n285 VTAIL.n284 171.744
R458 VTAIL.n284 VTAIL.n274 171.744
R459 VTAIL.n277 VTAIL.n274 171.744
R460 VTAIL.n608 VTAIL.t2 85.8723
R461 VTAIL.n28 VTAIL.t1 85.8723
R462 VTAIL.n110 VTAIL.t10 85.8723
R463 VTAIL.n194 VTAIL.t14 85.8723
R464 VTAIL.n527 VTAIL.t15 85.8723
R465 VTAIL.n443 VTAIL.t12 85.8723
R466 VTAIL.n361 VTAIL.t5 85.8723
R467 VTAIL.n277 VTAIL.t3 85.8723
R468 VTAIL.n499 VTAIL.n498 54.2817
R469 VTAIL.n333 VTAIL.n332 54.2817
R470 VTAIL.n1 VTAIL.n0 54.2815
R471 VTAIL.n167 VTAIL.n166 54.2815
R472 VTAIL.n663 VTAIL.n662 32.3793
R473 VTAIL.n83 VTAIL.n82 32.3793
R474 VTAIL.n165 VTAIL.n164 32.3793
R475 VTAIL.n249 VTAIL.n248 32.3793
R476 VTAIL.n581 VTAIL.n580 32.3793
R477 VTAIL.n497 VTAIL.n496 32.3793
R478 VTAIL.n415 VTAIL.n414 32.3793
R479 VTAIL.n331 VTAIL.n330 32.3793
R480 VTAIL.n663 VTAIL.n581 28.2117
R481 VTAIL.n331 VTAIL.n249 28.2117
R482 VTAIL.n609 VTAIL.n607 16.3895
R483 VTAIL.n29 VTAIL.n27 16.3895
R484 VTAIL.n111 VTAIL.n109 16.3895
R485 VTAIL.n195 VTAIL.n193 16.3895
R486 VTAIL.n528 VTAIL.n526 16.3895
R487 VTAIL.n444 VTAIL.n442 16.3895
R488 VTAIL.n362 VTAIL.n360 16.3895
R489 VTAIL.n278 VTAIL.n276 16.3895
R490 VTAIL.n656 VTAIL.n655 13.1884
R491 VTAIL.n76 VTAIL.n75 13.1884
R492 VTAIL.n158 VTAIL.n157 13.1884
R493 VTAIL.n242 VTAIL.n241 13.1884
R494 VTAIL.n574 VTAIL.n573 13.1884
R495 VTAIL.n490 VTAIL.n489 13.1884
R496 VTAIL.n408 VTAIL.n407 13.1884
R497 VTAIL.n324 VTAIL.n323 13.1884
R498 VTAIL.n610 VTAIL.n606 12.8005
R499 VTAIL.n654 VTAIL.n586 12.8005
R500 VTAIL.n659 VTAIL.n584 12.8005
R501 VTAIL.n30 VTAIL.n26 12.8005
R502 VTAIL.n74 VTAIL.n6 12.8005
R503 VTAIL.n79 VTAIL.n4 12.8005
R504 VTAIL.n112 VTAIL.n108 12.8005
R505 VTAIL.n156 VTAIL.n88 12.8005
R506 VTAIL.n161 VTAIL.n86 12.8005
R507 VTAIL.n196 VTAIL.n192 12.8005
R508 VTAIL.n240 VTAIL.n172 12.8005
R509 VTAIL.n245 VTAIL.n170 12.8005
R510 VTAIL.n577 VTAIL.n502 12.8005
R511 VTAIL.n572 VTAIL.n504 12.8005
R512 VTAIL.n529 VTAIL.n525 12.8005
R513 VTAIL.n493 VTAIL.n418 12.8005
R514 VTAIL.n488 VTAIL.n420 12.8005
R515 VTAIL.n445 VTAIL.n441 12.8005
R516 VTAIL.n411 VTAIL.n336 12.8005
R517 VTAIL.n406 VTAIL.n338 12.8005
R518 VTAIL.n363 VTAIL.n359 12.8005
R519 VTAIL.n327 VTAIL.n252 12.8005
R520 VTAIL.n322 VTAIL.n254 12.8005
R521 VTAIL.n279 VTAIL.n275 12.8005
R522 VTAIL.n614 VTAIL.n613 12.0247
R523 VTAIL.n651 VTAIL.n650 12.0247
R524 VTAIL.n660 VTAIL.n582 12.0247
R525 VTAIL.n34 VTAIL.n33 12.0247
R526 VTAIL.n71 VTAIL.n70 12.0247
R527 VTAIL.n80 VTAIL.n2 12.0247
R528 VTAIL.n116 VTAIL.n115 12.0247
R529 VTAIL.n153 VTAIL.n152 12.0247
R530 VTAIL.n162 VTAIL.n84 12.0247
R531 VTAIL.n200 VTAIL.n199 12.0247
R532 VTAIL.n237 VTAIL.n236 12.0247
R533 VTAIL.n246 VTAIL.n168 12.0247
R534 VTAIL.n578 VTAIL.n500 12.0247
R535 VTAIL.n569 VTAIL.n568 12.0247
R536 VTAIL.n533 VTAIL.n532 12.0247
R537 VTAIL.n494 VTAIL.n416 12.0247
R538 VTAIL.n485 VTAIL.n484 12.0247
R539 VTAIL.n449 VTAIL.n448 12.0247
R540 VTAIL.n412 VTAIL.n334 12.0247
R541 VTAIL.n403 VTAIL.n402 12.0247
R542 VTAIL.n367 VTAIL.n366 12.0247
R543 VTAIL.n328 VTAIL.n250 12.0247
R544 VTAIL.n319 VTAIL.n318 12.0247
R545 VTAIL.n283 VTAIL.n282 12.0247
R546 VTAIL.n617 VTAIL.n604 11.249
R547 VTAIL.n646 VTAIL.n588 11.249
R548 VTAIL.n37 VTAIL.n24 11.249
R549 VTAIL.n66 VTAIL.n8 11.249
R550 VTAIL.n119 VTAIL.n106 11.249
R551 VTAIL.n148 VTAIL.n90 11.249
R552 VTAIL.n203 VTAIL.n190 11.249
R553 VTAIL.n232 VTAIL.n174 11.249
R554 VTAIL.n565 VTAIL.n506 11.249
R555 VTAIL.n536 VTAIL.n523 11.249
R556 VTAIL.n481 VTAIL.n422 11.249
R557 VTAIL.n452 VTAIL.n439 11.249
R558 VTAIL.n399 VTAIL.n340 11.249
R559 VTAIL.n370 VTAIL.n357 11.249
R560 VTAIL.n315 VTAIL.n256 11.249
R561 VTAIL.n286 VTAIL.n273 11.249
R562 VTAIL.n618 VTAIL.n602 10.4732
R563 VTAIL.n645 VTAIL.n590 10.4732
R564 VTAIL.n38 VTAIL.n22 10.4732
R565 VTAIL.n65 VTAIL.n10 10.4732
R566 VTAIL.n120 VTAIL.n104 10.4732
R567 VTAIL.n147 VTAIL.n92 10.4732
R568 VTAIL.n204 VTAIL.n188 10.4732
R569 VTAIL.n231 VTAIL.n176 10.4732
R570 VTAIL.n564 VTAIL.n509 10.4732
R571 VTAIL.n537 VTAIL.n521 10.4732
R572 VTAIL.n480 VTAIL.n425 10.4732
R573 VTAIL.n453 VTAIL.n437 10.4732
R574 VTAIL.n398 VTAIL.n343 10.4732
R575 VTAIL.n371 VTAIL.n355 10.4732
R576 VTAIL.n314 VTAIL.n259 10.4732
R577 VTAIL.n287 VTAIL.n271 10.4732
R578 VTAIL.n622 VTAIL.n621 9.69747
R579 VTAIL.n642 VTAIL.n641 9.69747
R580 VTAIL.n42 VTAIL.n41 9.69747
R581 VTAIL.n62 VTAIL.n61 9.69747
R582 VTAIL.n124 VTAIL.n123 9.69747
R583 VTAIL.n144 VTAIL.n143 9.69747
R584 VTAIL.n208 VTAIL.n207 9.69747
R585 VTAIL.n228 VTAIL.n227 9.69747
R586 VTAIL.n561 VTAIL.n560 9.69747
R587 VTAIL.n541 VTAIL.n540 9.69747
R588 VTAIL.n477 VTAIL.n476 9.69747
R589 VTAIL.n457 VTAIL.n456 9.69747
R590 VTAIL.n395 VTAIL.n394 9.69747
R591 VTAIL.n375 VTAIL.n374 9.69747
R592 VTAIL.n311 VTAIL.n310 9.69747
R593 VTAIL.n291 VTAIL.n290 9.69747
R594 VTAIL.n662 VTAIL.n661 9.45567
R595 VTAIL.n82 VTAIL.n81 9.45567
R596 VTAIL.n164 VTAIL.n163 9.45567
R597 VTAIL.n248 VTAIL.n247 9.45567
R598 VTAIL.n580 VTAIL.n579 9.45567
R599 VTAIL.n496 VTAIL.n495 9.45567
R600 VTAIL.n414 VTAIL.n413 9.45567
R601 VTAIL.n330 VTAIL.n329 9.45567
R602 VTAIL.n661 VTAIL.n660 9.3005
R603 VTAIL.n584 VTAIL.n583 9.3005
R604 VTAIL.n629 VTAIL.n628 9.3005
R605 VTAIL.n627 VTAIL.n626 9.3005
R606 VTAIL.n600 VTAIL.n599 9.3005
R607 VTAIL.n621 VTAIL.n620 9.3005
R608 VTAIL.n619 VTAIL.n618 9.3005
R609 VTAIL.n604 VTAIL.n603 9.3005
R610 VTAIL.n613 VTAIL.n612 9.3005
R611 VTAIL.n611 VTAIL.n610 9.3005
R612 VTAIL.n596 VTAIL.n595 9.3005
R613 VTAIL.n635 VTAIL.n634 9.3005
R614 VTAIL.n637 VTAIL.n636 9.3005
R615 VTAIL.n592 VTAIL.n591 9.3005
R616 VTAIL.n643 VTAIL.n642 9.3005
R617 VTAIL.n645 VTAIL.n644 9.3005
R618 VTAIL.n588 VTAIL.n587 9.3005
R619 VTAIL.n652 VTAIL.n651 9.3005
R620 VTAIL.n654 VTAIL.n653 9.3005
R621 VTAIL.n81 VTAIL.n80 9.3005
R622 VTAIL.n4 VTAIL.n3 9.3005
R623 VTAIL.n49 VTAIL.n48 9.3005
R624 VTAIL.n47 VTAIL.n46 9.3005
R625 VTAIL.n20 VTAIL.n19 9.3005
R626 VTAIL.n41 VTAIL.n40 9.3005
R627 VTAIL.n39 VTAIL.n38 9.3005
R628 VTAIL.n24 VTAIL.n23 9.3005
R629 VTAIL.n33 VTAIL.n32 9.3005
R630 VTAIL.n31 VTAIL.n30 9.3005
R631 VTAIL.n16 VTAIL.n15 9.3005
R632 VTAIL.n55 VTAIL.n54 9.3005
R633 VTAIL.n57 VTAIL.n56 9.3005
R634 VTAIL.n12 VTAIL.n11 9.3005
R635 VTAIL.n63 VTAIL.n62 9.3005
R636 VTAIL.n65 VTAIL.n64 9.3005
R637 VTAIL.n8 VTAIL.n7 9.3005
R638 VTAIL.n72 VTAIL.n71 9.3005
R639 VTAIL.n74 VTAIL.n73 9.3005
R640 VTAIL.n163 VTAIL.n162 9.3005
R641 VTAIL.n86 VTAIL.n85 9.3005
R642 VTAIL.n131 VTAIL.n130 9.3005
R643 VTAIL.n129 VTAIL.n128 9.3005
R644 VTAIL.n102 VTAIL.n101 9.3005
R645 VTAIL.n123 VTAIL.n122 9.3005
R646 VTAIL.n121 VTAIL.n120 9.3005
R647 VTAIL.n106 VTAIL.n105 9.3005
R648 VTAIL.n115 VTAIL.n114 9.3005
R649 VTAIL.n113 VTAIL.n112 9.3005
R650 VTAIL.n98 VTAIL.n97 9.3005
R651 VTAIL.n137 VTAIL.n136 9.3005
R652 VTAIL.n139 VTAIL.n138 9.3005
R653 VTAIL.n94 VTAIL.n93 9.3005
R654 VTAIL.n145 VTAIL.n144 9.3005
R655 VTAIL.n147 VTAIL.n146 9.3005
R656 VTAIL.n90 VTAIL.n89 9.3005
R657 VTAIL.n154 VTAIL.n153 9.3005
R658 VTAIL.n156 VTAIL.n155 9.3005
R659 VTAIL.n247 VTAIL.n246 9.3005
R660 VTAIL.n170 VTAIL.n169 9.3005
R661 VTAIL.n215 VTAIL.n214 9.3005
R662 VTAIL.n213 VTAIL.n212 9.3005
R663 VTAIL.n186 VTAIL.n185 9.3005
R664 VTAIL.n207 VTAIL.n206 9.3005
R665 VTAIL.n205 VTAIL.n204 9.3005
R666 VTAIL.n190 VTAIL.n189 9.3005
R667 VTAIL.n199 VTAIL.n198 9.3005
R668 VTAIL.n197 VTAIL.n196 9.3005
R669 VTAIL.n182 VTAIL.n181 9.3005
R670 VTAIL.n221 VTAIL.n220 9.3005
R671 VTAIL.n223 VTAIL.n222 9.3005
R672 VTAIL.n178 VTAIL.n177 9.3005
R673 VTAIL.n229 VTAIL.n228 9.3005
R674 VTAIL.n231 VTAIL.n230 9.3005
R675 VTAIL.n174 VTAIL.n173 9.3005
R676 VTAIL.n238 VTAIL.n237 9.3005
R677 VTAIL.n240 VTAIL.n239 9.3005
R678 VTAIL.n554 VTAIL.n553 9.3005
R679 VTAIL.n556 VTAIL.n555 9.3005
R680 VTAIL.n511 VTAIL.n510 9.3005
R681 VTAIL.n562 VTAIL.n561 9.3005
R682 VTAIL.n564 VTAIL.n563 9.3005
R683 VTAIL.n506 VTAIL.n505 9.3005
R684 VTAIL.n570 VTAIL.n569 9.3005
R685 VTAIL.n572 VTAIL.n571 9.3005
R686 VTAIL.n579 VTAIL.n578 9.3005
R687 VTAIL.n502 VTAIL.n501 9.3005
R688 VTAIL.n515 VTAIL.n514 9.3005
R689 VTAIL.n548 VTAIL.n547 9.3005
R690 VTAIL.n546 VTAIL.n545 9.3005
R691 VTAIL.n519 VTAIL.n518 9.3005
R692 VTAIL.n540 VTAIL.n539 9.3005
R693 VTAIL.n538 VTAIL.n537 9.3005
R694 VTAIL.n523 VTAIL.n522 9.3005
R695 VTAIL.n532 VTAIL.n531 9.3005
R696 VTAIL.n530 VTAIL.n529 9.3005
R697 VTAIL.n470 VTAIL.n469 9.3005
R698 VTAIL.n472 VTAIL.n471 9.3005
R699 VTAIL.n427 VTAIL.n426 9.3005
R700 VTAIL.n478 VTAIL.n477 9.3005
R701 VTAIL.n480 VTAIL.n479 9.3005
R702 VTAIL.n422 VTAIL.n421 9.3005
R703 VTAIL.n486 VTAIL.n485 9.3005
R704 VTAIL.n488 VTAIL.n487 9.3005
R705 VTAIL.n495 VTAIL.n494 9.3005
R706 VTAIL.n418 VTAIL.n417 9.3005
R707 VTAIL.n431 VTAIL.n430 9.3005
R708 VTAIL.n464 VTAIL.n463 9.3005
R709 VTAIL.n462 VTAIL.n461 9.3005
R710 VTAIL.n435 VTAIL.n434 9.3005
R711 VTAIL.n456 VTAIL.n455 9.3005
R712 VTAIL.n454 VTAIL.n453 9.3005
R713 VTAIL.n439 VTAIL.n438 9.3005
R714 VTAIL.n448 VTAIL.n447 9.3005
R715 VTAIL.n446 VTAIL.n445 9.3005
R716 VTAIL.n388 VTAIL.n387 9.3005
R717 VTAIL.n390 VTAIL.n389 9.3005
R718 VTAIL.n345 VTAIL.n344 9.3005
R719 VTAIL.n396 VTAIL.n395 9.3005
R720 VTAIL.n398 VTAIL.n397 9.3005
R721 VTAIL.n340 VTAIL.n339 9.3005
R722 VTAIL.n404 VTAIL.n403 9.3005
R723 VTAIL.n406 VTAIL.n405 9.3005
R724 VTAIL.n413 VTAIL.n412 9.3005
R725 VTAIL.n336 VTAIL.n335 9.3005
R726 VTAIL.n349 VTAIL.n348 9.3005
R727 VTAIL.n382 VTAIL.n381 9.3005
R728 VTAIL.n380 VTAIL.n379 9.3005
R729 VTAIL.n353 VTAIL.n352 9.3005
R730 VTAIL.n374 VTAIL.n373 9.3005
R731 VTAIL.n372 VTAIL.n371 9.3005
R732 VTAIL.n357 VTAIL.n356 9.3005
R733 VTAIL.n366 VTAIL.n365 9.3005
R734 VTAIL.n364 VTAIL.n363 9.3005
R735 VTAIL.n304 VTAIL.n303 9.3005
R736 VTAIL.n306 VTAIL.n305 9.3005
R737 VTAIL.n261 VTAIL.n260 9.3005
R738 VTAIL.n312 VTAIL.n311 9.3005
R739 VTAIL.n314 VTAIL.n313 9.3005
R740 VTAIL.n256 VTAIL.n255 9.3005
R741 VTAIL.n320 VTAIL.n319 9.3005
R742 VTAIL.n322 VTAIL.n321 9.3005
R743 VTAIL.n329 VTAIL.n328 9.3005
R744 VTAIL.n252 VTAIL.n251 9.3005
R745 VTAIL.n265 VTAIL.n264 9.3005
R746 VTAIL.n298 VTAIL.n297 9.3005
R747 VTAIL.n296 VTAIL.n295 9.3005
R748 VTAIL.n269 VTAIL.n268 9.3005
R749 VTAIL.n290 VTAIL.n289 9.3005
R750 VTAIL.n288 VTAIL.n287 9.3005
R751 VTAIL.n273 VTAIL.n272 9.3005
R752 VTAIL.n282 VTAIL.n281 9.3005
R753 VTAIL.n280 VTAIL.n279 9.3005
R754 VTAIL.n625 VTAIL.n600 8.92171
R755 VTAIL.n638 VTAIL.n592 8.92171
R756 VTAIL.n45 VTAIL.n20 8.92171
R757 VTAIL.n58 VTAIL.n12 8.92171
R758 VTAIL.n127 VTAIL.n102 8.92171
R759 VTAIL.n140 VTAIL.n94 8.92171
R760 VTAIL.n211 VTAIL.n186 8.92171
R761 VTAIL.n224 VTAIL.n178 8.92171
R762 VTAIL.n557 VTAIL.n511 8.92171
R763 VTAIL.n544 VTAIL.n519 8.92171
R764 VTAIL.n473 VTAIL.n427 8.92171
R765 VTAIL.n460 VTAIL.n435 8.92171
R766 VTAIL.n391 VTAIL.n345 8.92171
R767 VTAIL.n378 VTAIL.n353 8.92171
R768 VTAIL.n307 VTAIL.n261 8.92171
R769 VTAIL.n294 VTAIL.n269 8.92171
R770 VTAIL.n626 VTAIL.n598 8.14595
R771 VTAIL.n637 VTAIL.n594 8.14595
R772 VTAIL.n46 VTAIL.n18 8.14595
R773 VTAIL.n57 VTAIL.n14 8.14595
R774 VTAIL.n128 VTAIL.n100 8.14595
R775 VTAIL.n139 VTAIL.n96 8.14595
R776 VTAIL.n212 VTAIL.n184 8.14595
R777 VTAIL.n223 VTAIL.n180 8.14595
R778 VTAIL.n556 VTAIL.n513 8.14595
R779 VTAIL.n545 VTAIL.n517 8.14595
R780 VTAIL.n472 VTAIL.n429 8.14595
R781 VTAIL.n461 VTAIL.n433 8.14595
R782 VTAIL.n390 VTAIL.n347 8.14595
R783 VTAIL.n379 VTAIL.n351 8.14595
R784 VTAIL.n306 VTAIL.n263 8.14595
R785 VTAIL.n295 VTAIL.n267 8.14595
R786 VTAIL.n630 VTAIL.n629 7.3702
R787 VTAIL.n634 VTAIL.n633 7.3702
R788 VTAIL.n50 VTAIL.n49 7.3702
R789 VTAIL.n54 VTAIL.n53 7.3702
R790 VTAIL.n132 VTAIL.n131 7.3702
R791 VTAIL.n136 VTAIL.n135 7.3702
R792 VTAIL.n216 VTAIL.n215 7.3702
R793 VTAIL.n220 VTAIL.n219 7.3702
R794 VTAIL.n553 VTAIL.n552 7.3702
R795 VTAIL.n549 VTAIL.n548 7.3702
R796 VTAIL.n469 VTAIL.n468 7.3702
R797 VTAIL.n465 VTAIL.n464 7.3702
R798 VTAIL.n387 VTAIL.n386 7.3702
R799 VTAIL.n383 VTAIL.n382 7.3702
R800 VTAIL.n303 VTAIL.n302 7.3702
R801 VTAIL.n299 VTAIL.n298 7.3702
R802 VTAIL.n630 VTAIL.n596 6.59444
R803 VTAIL.n633 VTAIL.n596 6.59444
R804 VTAIL.n50 VTAIL.n16 6.59444
R805 VTAIL.n53 VTAIL.n16 6.59444
R806 VTAIL.n132 VTAIL.n98 6.59444
R807 VTAIL.n135 VTAIL.n98 6.59444
R808 VTAIL.n216 VTAIL.n182 6.59444
R809 VTAIL.n219 VTAIL.n182 6.59444
R810 VTAIL.n552 VTAIL.n515 6.59444
R811 VTAIL.n549 VTAIL.n515 6.59444
R812 VTAIL.n468 VTAIL.n431 6.59444
R813 VTAIL.n465 VTAIL.n431 6.59444
R814 VTAIL.n386 VTAIL.n349 6.59444
R815 VTAIL.n383 VTAIL.n349 6.59444
R816 VTAIL.n302 VTAIL.n265 6.59444
R817 VTAIL.n299 VTAIL.n265 6.59444
R818 VTAIL.n629 VTAIL.n598 5.81868
R819 VTAIL.n634 VTAIL.n594 5.81868
R820 VTAIL.n49 VTAIL.n18 5.81868
R821 VTAIL.n54 VTAIL.n14 5.81868
R822 VTAIL.n131 VTAIL.n100 5.81868
R823 VTAIL.n136 VTAIL.n96 5.81868
R824 VTAIL.n215 VTAIL.n184 5.81868
R825 VTAIL.n220 VTAIL.n180 5.81868
R826 VTAIL.n553 VTAIL.n513 5.81868
R827 VTAIL.n548 VTAIL.n517 5.81868
R828 VTAIL.n469 VTAIL.n429 5.81868
R829 VTAIL.n464 VTAIL.n433 5.81868
R830 VTAIL.n387 VTAIL.n347 5.81868
R831 VTAIL.n382 VTAIL.n351 5.81868
R832 VTAIL.n303 VTAIL.n263 5.81868
R833 VTAIL.n298 VTAIL.n267 5.81868
R834 VTAIL.n626 VTAIL.n625 5.04292
R835 VTAIL.n638 VTAIL.n637 5.04292
R836 VTAIL.n46 VTAIL.n45 5.04292
R837 VTAIL.n58 VTAIL.n57 5.04292
R838 VTAIL.n128 VTAIL.n127 5.04292
R839 VTAIL.n140 VTAIL.n139 5.04292
R840 VTAIL.n212 VTAIL.n211 5.04292
R841 VTAIL.n224 VTAIL.n223 5.04292
R842 VTAIL.n557 VTAIL.n556 5.04292
R843 VTAIL.n545 VTAIL.n544 5.04292
R844 VTAIL.n473 VTAIL.n472 5.04292
R845 VTAIL.n461 VTAIL.n460 5.04292
R846 VTAIL.n391 VTAIL.n390 5.04292
R847 VTAIL.n379 VTAIL.n378 5.04292
R848 VTAIL.n307 VTAIL.n306 5.04292
R849 VTAIL.n295 VTAIL.n294 5.04292
R850 VTAIL.n622 VTAIL.n600 4.26717
R851 VTAIL.n641 VTAIL.n592 4.26717
R852 VTAIL.n42 VTAIL.n20 4.26717
R853 VTAIL.n61 VTAIL.n12 4.26717
R854 VTAIL.n124 VTAIL.n102 4.26717
R855 VTAIL.n143 VTAIL.n94 4.26717
R856 VTAIL.n208 VTAIL.n186 4.26717
R857 VTAIL.n227 VTAIL.n178 4.26717
R858 VTAIL.n560 VTAIL.n511 4.26717
R859 VTAIL.n541 VTAIL.n519 4.26717
R860 VTAIL.n476 VTAIL.n427 4.26717
R861 VTAIL.n457 VTAIL.n435 4.26717
R862 VTAIL.n394 VTAIL.n345 4.26717
R863 VTAIL.n375 VTAIL.n353 4.26717
R864 VTAIL.n310 VTAIL.n261 4.26717
R865 VTAIL.n291 VTAIL.n269 4.26717
R866 VTAIL.n611 VTAIL.n607 3.70982
R867 VTAIL.n31 VTAIL.n27 3.70982
R868 VTAIL.n113 VTAIL.n109 3.70982
R869 VTAIL.n197 VTAIL.n193 3.70982
R870 VTAIL.n530 VTAIL.n526 3.70982
R871 VTAIL.n446 VTAIL.n442 3.70982
R872 VTAIL.n364 VTAIL.n360 3.70982
R873 VTAIL.n280 VTAIL.n276 3.70982
R874 VTAIL.n621 VTAIL.n602 3.49141
R875 VTAIL.n642 VTAIL.n590 3.49141
R876 VTAIL.n41 VTAIL.n22 3.49141
R877 VTAIL.n62 VTAIL.n10 3.49141
R878 VTAIL.n123 VTAIL.n104 3.49141
R879 VTAIL.n144 VTAIL.n92 3.49141
R880 VTAIL.n207 VTAIL.n188 3.49141
R881 VTAIL.n228 VTAIL.n176 3.49141
R882 VTAIL.n561 VTAIL.n509 3.49141
R883 VTAIL.n540 VTAIL.n521 3.49141
R884 VTAIL.n477 VTAIL.n425 3.49141
R885 VTAIL.n456 VTAIL.n437 3.49141
R886 VTAIL.n395 VTAIL.n343 3.49141
R887 VTAIL.n374 VTAIL.n355 3.49141
R888 VTAIL.n311 VTAIL.n259 3.49141
R889 VTAIL.n290 VTAIL.n271 3.49141
R890 VTAIL.n333 VTAIL.n331 3.21602
R891 VTAIL.n415 VTAIL.n333 3.21602
R892 VTAIL.n499 VTAIL.n497 3.21602
R893 VTAIL.n581 VTAIL.n499 3.21602
R894 VTAIL.n249 VTAIL.n167 3.21602
R895 VTAIL.n167 VTAIL.n165 3.21602
R896 VTAIL.n83 VTAIL.n1 3.21602
R897 VTAIL VTAIL.n663 3.15783
R898 VTAIL.n618 VTAIL.n617 2.71565
R899 VTAIL.n646 VTAIL.n645 2.71565
R900 VTAIL.n38 VTAIL.n37 2.71565
R901 VTAIL.n66 VTAIL.n65 2.71565
R902 VTAIL.n120 VTAIL.n119 2.71565
R903 VTAIL.n148 VTAIL.n147 2.71565
R904 VTAIL.n204 VTAIL.n203 2.71565
R905 VTAIL.n232 VTAIL.n231 2.71565
R906 VTAIL.n565 VTAIL.n564 2.71565
R907 VTAIL.n537 VTAIL.n536 2.71565
R908 VTAIL.n481 VTAIL.n480 2.71565
R909 VTAIL.n453 VTAIL.n452 2.71565
R910 VTAIL.n399 VTAIL.n398 2.71565
R911 VTAIL.n371 VTAIL.n370 2.71565
R912 VTAIL.n315 VTAIL.n314 2.71565
R913 VTAIL.n287 VTAIL.n286 2.71565
R914 VTAIL.n0 VTAIL.t4 2.21927
R915 VTAIL.n0 VTAIL.t7 2.21927
R916 VTAIL.n166 VTAIL.t9 2.21927
R917 VTAIL.n166 VTAIL.t11 2.21927
R918 VTAIL.n498 VTAIL.t8 2.21927
R919 VTAIL.n498 VTAIL.t13 2.21927
R920 VTAIL.n332 VTAIL.t6 2.21927
R921 VTAIL.n332 VTAIL.t0 2.21927
R922 VTAIL.n614 VTAIL.n604 1.93989
R923 VTAIL.n650 VTAIL.n588 1.93989
R924 VTAIL.n662 VTAIL.n582 1.93989
R925 VTAIL.n34 VTAIL.n24 1.93989
R926 VTAIL.n70 VTAIL.n8 1.93989
R927 VTAIL.n82 VTAIL.n2 1.93989
R928 VTAIL.n116 VTAIL.n106 1.93989
R929 VTAIL.n152 VTAIL.n90 1.93989
R930 VTAIL.n164 VTAIL.n84 1.93989
R931 VTAIL.n200 VTAIL.n190 1.93989
R932 VTAIL.n236 VTAIL.n174 1.93989
R933 VTAIL.n248 VTAIL.n168 1.93989
R934 VTAIL.n580 VTAIL.n500 1.93989
R935 VTAIL.n568 VTAIL.n506 1.93989
R936 VTAIL.n533 VTAIL.n523 1.93989
R937 VTAIL.n496 VTAIL.n416 1.93989
R938 VTAIL.n484 VTAIL.n422 1.93989
R939 VTAIL.n449 VTAIL.n439 1.93989
R940 VTAIL.n414 VTAIL.n334 1.93989
R941 VTAIL.n402 VTAIL.n340 1.93989
R942 VTAIL.n367 VTAIL.n357 1.93989
R943 VTAIL.n330 VTAIL.n250 1.93989
R944 VTAIL.n318 VTAIL.n256 1.93989
R945 VTAIL.n283 VTAIL.n273 1.93989
R946 VTAIL.n613 VTAIL.n606 1.16414
R947 VTAIL.n651 VTAIL.n586 1.16414
R948 VTAIL.n660 VTAIL.n659 1.16414
R949 VTAIL.n33 VTAIL.n26 1.16414
R950 VTAIL.n71 VTAIL.n6 1.16414
R951 VTAIL.n80 VTAIL.n79 1.16414
R952 VTAIL.n115 VTAIL.n108 1.16414
R953 VTAIL.n153 VTAIL.n88 1.16414
R954 VTAIL.n162 VTAIL.n161 1.16414
R955 VTAIL.n199 VTAIL.n192 1.16414
R956 VTAIL.n237 VTAIL.n172 1.16414
R957 VTAIL.n246 VTAIL.n245 1.16414
R958 VTAIL.n578 VTAIL.n577 1.16414
R959 VTAIL.n569 VTAIL.n504 1.16414
R960 VTAIL.n532 VTAIL.n525 1.16414
R961 VTAIL.n494 VTAIL.n493 1.16414
R962 VTAIL.n485 VTAIL.n420 1.16414
R963 VTAIL.n448 VTAIL.n441 1.16414
R964 VTAIL.n412 VTAIL.n411 1.16414
R965 VTAIL.n403 VTAIL.n338 1.16414
R966 VTAIL.n366 VTAIL.n359 1.16414
R967 VTAIL.n328 VTAIL.n327 1.16414
R968 VTAIL.n319 VTAIL.n254 1.16414
R969 VTAIL.n282 VTAIL.n275 1.16414
R970 VTAIL.n497 VTAIL.n415 0.470328
R971 VTAIL.n165 VTAIL.n83 0.470328
R972 VTAIL.n610 VTAIL.n609 0.388379
R973 VTAIL.n655 VTAIL.n654 0.388379
R974 VTAIL.n656 VTAIL.n584 0.388379
R975 VTAIL.n30 VTAIL.n29 0.388379
R976 VTAIL.n75 VTAIL.n74 0.388379
R977 VTAIL.n76 VTAIL.n4 0.388379
R978 VTAIL.n112 VTAIL.n111 0.388379
R979 VTAIL.n157 VTAIL.n156 0.388379
R980 VTAIL.n158 VTAIL.n86 0.388379
R981 VTAIL.n196 VTAIL.n195 0.388379
R982 VTAIL.n241 VTAIL.n240 0.388379
R983 VTAIL.n242 VTAIL.n170 0.388379
R984 VTAIL.n574 VTAIL.n502 0.388379
R985 VTAIL.n573 VTAIL.n572 0.388379
R986 VTAIL.n529 VTAIL.n528 0.388379
R987 VTAIL.n490 VTAIL.n418 0.388379
R988 VTAIL.n489 VTAIL.n488 0.388379
R989 VTAIL.n445 VTAIL.n444 0.388379
R990 VTAIL.n408 VTAIL.n336 0.388379
R991 VTAIL.n407 VTAIL.n406 0.388379
R992 VTAIL.n363 VTAIL.n362 0.388379
R993 VTAIL.n324 VTAIL.n252 0.388379
R994 VTAIL.n323 VTAIL.n322 0.388379
R995 VTAIL.n279 VTAIL.n278 0.388379
R996 VTAIL.n612 VTAIL.n611 0.155672
R997 VTAIL.n612 VTAIL.n603 0.155672
R998 VTAIL.n619 VTAIL.n603 0.155672
R999 VTAIL.n620 VTAIL.n619 0.155672
R1000 VTAIL.n620 VTAIL.n599 0.155672
R1001 VTAIL.n627 VTAIL.n599 0.155672
R1002 VTAIL.n628 VTAIL.n627 0.155672
R1003 VTAIL.n628 VTAIL.n595 0.155672
R1004 VTAIL.n635 VTAIL.n595 0.155672
R1005 VTAIL.n636 VTAIL.n635 0.155672
R1006 VTAIL.n636 VTAIL.n591 0.155672
R1007 VTAIL.n643 VTAIL.n591 0.155672
R1008 VTAIL.n644 VTAIL.n643 0.155672
R1009 VTAIL.n644 VTAIL.n587 0.155672
R1010 VTAIL.n652 VTAIL.n587 0.155672
R1011 VTAIL.n653 VTAIL.n652 0.155672
R1012 VTAIL.n653 VTAIL.n583 0.155672
R1013 VTAIL.n661 VTAIL.n583 0.155672
R1014 VTAIL.n32 VTAIL.n31 0.155672
R1015 VTAIL.n32 VTAIL.n23 0.155672
R1016 VTAIL.n39 VTAIL.n23 0.155672
R1017 VTAIL.n40 VTAIL.n39 0.155672
R1018 VTAIL.n40 VTAIL.n19 0.155672
R1019 VTAIL.n47 VTAIL.n19 0.155672
R1020 VTAIL.n48 VTAIL.n47 0.155672
R1021 VTAIL.n48 VTAIL.n15 0.155672
R1022 VTAIL.n55 VTAIL.n15 0.155672
R1023 VTAIL.n56 VTAIL.n55 0.155672
R1024 VTAIL.n56 VTAIL.n11 0.155672
R1025 VTAIL.n63 VTAIL.n11 0.155672
R1026 VTAIL.n64 VTAIL.n63 0.155672
R1027 VTAIL.n64 VTAIL.n7 0.155672
R1028 VTAIL.n72 VTAIL.n7 0.155672
R1029 VTAIL.n73 VTAIL.n72 0.155672
R1030 VTAIL.n73 VTAIL.n3 0.155672
R1031 VTAIL.n81 VTAIL.n3 0.155672
R1032 VTAIL.n114 VTAIL.n113 0.155672
R1033 VTAIL.n114 VTAIL.n105 0.155672
R1034 VTAIL.n121 VTAIL.n105 0.155672
R1035 VTAIL.n122 VTAIL.n121 0.155672
R1036 VTAIL.n122 VTAIL.n101 0.155672
R1037 VTAIL.n129 VTAIL.n101 0.155672
R1038 VTAIL.n130 VTAIL.n129 0.155672
R1039 VTAIL.n130 VTAIL.n97 0.155672
R1040 VTAIL.n137 VTAIL.n97 0.155672
R1041 VTAIL.n138 VTAIL.n137 0.155672
R1042 VTAIL.n138 VTAIL.n93 0.155672
R1043 VTAIL.n145 VTAIL.n93 0.155672
R1044 VTAIL.n146 VTAIL.n145 0.155672
R1045 VTAIL.n146 VTAIL.n89 0.155672
R1046 VTAIL.n154 VTAIL.n89 0.155672
R1047 VTAIL.n155 VTAIL.n154 0.155672
R1048 VTAIL.n155 VTAIL.n85 0.155672
R1049 VTAIL.n163 VTAIL.n85 0.155672
R1050 VTAIL.n198 VTAIL.n197 0.155672
R1051 VTAIL.n198 VTAIL.n189 0.155672
R1052 VTAIL.n205 VTAIL.n189 0.155672
R1053 VTAIL.n206 VTAIL.n205 0.155672
R1054 VTAIL.n206 VTAIL.n185 0.155672
R1055 VTAIL.n213 VTAIL.n185 0.155672
R1056 VTAIL.n214 VTAIL.n213 0.155672
R1057 VTAIL.n214 VTAIL.n181 0.155672
R1058 VTAIL.n221 VTAIL.n181 0.155672
R1059 VTAIL.n222 VTAIL.n221 0.155672
R1060 VTAIL.n222 VTAIL.n177 0.155672
R1061 VTAIL.n229 VTAIL.n177 0.155672
R1062 VTAIL.n230 VTAIL.n229 0.155672
R1063 VTAIL.n230 VTAIL.n173 0.155672
R1064 VTAIL.n238 VTAIL.n173 0.155672
R1065 VTAIL.n239 VTAIL.n238 0.155672
R1066 VTAIL.n239 VTAIL.n169 0.155672
R1067 VTAIL.n247 VTAIL.n169 0.155672
R1068 VTAIL.n579 VTAIL.n501 0.155672
R1069 VTAIL.n571 VTAIL.n501 0.155672
R1070 VTAIL.n571 VTAIL.n570 0.155672
R1071 VTAIL.n570 VTAIL.n505 0.155672
R1072 VTAIL.n563 VTAIL.n505 0.155672
R1073 VTAIL.n563 VTAIL.n562 0.155672
R1074 VTAIL.n562 VTAIL.n510 0.155672
R1075 VTAIL.n555 VTAIL.n510 0.155672
R1076 VTAIL.n555 VTAIL.n554 0.155672
R1077 VTAIL.n554 VTAIL.n514 0.155672
R1078 VTAIL.n547 VTAIL.n514 0.155672
R1079 VTAIL.n547 VTAIL.n546 0.155672
R1080 VTAIL.n546 VTAIL.n518 0.155672
R1081 VTAIL.n539 VTAIL.n518 0.155672
R1082 VTAIL.n539 VTAIL.n538 0.155672
R1083 VTAIL.n538 VTAIL.n522 0.155672
R1084 VTAIL.n531 VTAIL.n522 0.155672
R1085 VTAIL.n531 VTAIL.n530 0.155672
R1086 VTAIL.n495 VTAIL.n417 0.155672
R1087 VTAIL.n487 VTAIL.n417 0.155672
R1088 VTAIL.n487 VTAIL.n486 0.155672
R1089 VTAIL.n486 VTAIL.n421 0.155672
R1090 VTAIL.n479 VTAIL.n421 0.155672
R1091 VTAIL.n479 VTAIL.n478 0.155672
R1092 VTAIL.n478 VTAIL.n426 0.155672
R1093 VTAIL.n471 VTAIL.n426 0.155672
R1094 VTAIL.n471 VTAIL.n470 0.155672
R1095 VTAIL.n470 VTAIL.n430 0.155672
R1096 VTAIL.n463 VTAIL.n430 0.155672
R1097 VTAIL.n463 VTAIL.n462 0.155672
R1098 VTAIL.n462 VTAIL.n434 0.155672
R1099 VTAIL.n455 VTAIL.n434 0.155672
R1100 VTAIL.n455 VTAIL.n454 0.155672
R1101 VTAIL.n454 VTAIL.n438 0.155672
R1102 VTAIL.n447 VTAIL.n438 0.155672
R1103 VTAIL.n447 VTAIL.n446 0.155672
R1104 VTAIL.n413 VTAIL.n335 0.155672
R1105 VTAIL.n405 VTAIL.n335 0.155672
R1106 VTAIL.n405 VTAIL.n404 0.155672
R1107 VTAIL.n404 VTAIL.n339 0.155672
R1108 VTAIL.n397 VTAIL.n339 0.155672
R1109 VTAIL.n397 VTAIL.n396 0.155672
R1110 VTAIL.n396 VTAIL.n344 0.155672
R1111 VTAIL.n389 VTAIL.n344 0.155672
R1112 VTAIL.n389 VTAIL.n388 0.155672
R1113 VTAIL.n388 VTAIL.n348 0.155672
R1114 VTAIL.n381 VTAIL.n348 0.155672
R1115 VTAIL.n381 VTAIL.n380 0.155672
R1116 VTAIL.n380 VTAIL.n352 0.155672
R1117 VTAIL.n373 VTAIL.n352 0.155672
R1118 VTAIL.n373 VTAIL.n372 0.155672
R1119 VTAIL.n372 VTAIL.n356 0.155672
R1120 VTAIL.n365 VTAIL.n356 0.155672
R1121 VTAIL.n365 VTAIL.n364 0.155672
R1122 VTAIL.n329 VTAIL.n251 0.155672
R1123 VTAIL.n321 VTAIL.n251 0.155672
R1124 VTAIL.n321 VTAIL.n320 0.155672
R1125 VTAIL.n320 VTAIL.n255 0.155672
R1126 VTAIL.n313 VTAIL.n255 0.155672
R1127 VTAIL.n313 VTAIL.n312 0.155672
R1128 VTAIL.n312 VTAIL.n260 0.155672
R1129 VTAIL.n305 VTAIL.n260 0.155672
R1130 VTAIL.n305 VTAIL.n304 0.155672
R1131 VTAIL.n304 VTAIL.n264 0.155672
R1132 VTAIL.n297 VTAIL.n264 0.155672
R1133 VTAIL.n297 VTAIL.n296 0.155672
R1134 VTAIL.n296 VTAIL.n268 0.155672
R1135 VTAIL.n289 VTAIL.n268 0.155672
R1136 VTAIL.n289 VTAIL.n288 0.155672
R1137 VTAIL.n288 VTAIL.n272 0.155672
R1138 VTAIL.n281 VTAIL.n272 0.155672
R1139 VTAIL.n281 VTAIL.n280 0.155672
R1140 VTAIL VTAIL.n1 0.0586897
R1141 VDD1 VDD1.n0 72.6265
R1142 VDD1.n3 VDD1.n2 72.5127
R1143 VDD1.n3 VDD1.n1 72.5127
R1144 VDD1.n5 VDD1.n4 70.9603
R1145 VDD1.n5 VDD1.n3 51.3974
R1146 VDD1.n4 VDD1.t3 2.21927
R1147 VDD1.n4 VDD1.t5 2.21927
R1148 VDD1.n0 VDD1.t0 2.21927
R1149 VDD1.n0 VDD1.t2 2.21927
R1150 VDD1.n2 VDD1.t1 2.21927
R1151 VDD1.n2 VDD1.t7 2.21927
R1152 VDD1.n1 VDD1.t4 2.21927
R1153 VDD1.n1 VDD1.t6 2.21927
R1154 VDD1 VDD1.n5 1.55007
R1155 B.n693 B.n692 585
R1156 B.n694 B.n91 585
R1157 B.n696 B.n695 585
R1158 B.n697 B.n90 585
R1159 B.n699 B.n698 585
R1160 B.n700 B.n89 585
R1161 B.n702 B.n701 585
R1162 B.n703 B.n88 585
R1163 B.n705 B.n704 585
R1164 B.n706 B.n87 585
R1165 B.n708 B.n707 585
R1166 B.n709 B.n86 585
R1167 B.n711 B.n710 585
R1168 B.n712 B.n85 585
R1169 B.n714 B.n713 585
R1170 B.n715 B.n84 585
R1171 B.n717 B.n716 585
R1172 B.n718 B.n83 585
R1173 B.n720 B.n719 585
R1174 B.n721 B.n82 585
R1175 B.n723 B.n722 585
R1176 B.n724 B.n81 585
R1177 B.n726 B.n725 585
R1178 B.n727 B.n80 585
R1179 B.n729 B.n728 585
R1180 B.n730 B.n79 585
R1181 B.n732 B.n731 585
R1182 B.n733 B.n78 585
R1183 B.n735 B.n734 585
R1184 B.n736 B.n77 585
R1185 B.n738 B.n737 585
R1186 B.n739 B.n76 585
R1187 B.n741 B.n740 585
R1188 B.n742 B.n75 585
R1189 B.n744 B.n743 585
R1190 B.n745 B.n74 585
R1191 B.n747 B.n746 585
R1192 B.n748 B.n73 585
R1193 B.n750 B.n749 585
R1194 B.n751 B.n72 585
R1195 B.n753 B.n752 585
R1196 B.n754 B.n71 585
R1197 B.n756 B.n755 585
R1198 B.n757 B.n70 585
R1199 B.n759 B.n758 585
R1200 B.n760 B.n69 585
R1201 B.n762 B.n761 585
R1202 B.n763 B.n68 585
R1203 B.n765 B.n764 585
R1204 B.n767 B.n65 585
R1205 B.n769 B.n768 585
R1206 B.n770 B.n64 585
R1207 B.n772 B.n771 585
R1208 B.n773 B.n63 585
R1209 B.n775 B.n774 585
R1210 B.n776 B.n62 585
R1211 B.n778 B.n777 585
R1212 B.n779 B.n61 585
R1213 B.n781 B.n780 585
R1214 B.n783 B.n782 585
R1215 B.n784 B.n57 585
R1216 B.n786 B.n785 585
R1217 B.n787 B.n56 585
R1218 B.n789 B.n788 585
R1219 B.n790 B.n55 585
R1220 B.n792 B.n791 585
R1221 B.n793 B.n54 585
R1222 B.n795 B.n794 585
R1223 B.n796 B.n53 585
R1224 B.n798 B.n797 585
R1225 B.n799 B.n52 585
R1226 B.n801 B.n800 585
R1227 B.n802 B.n51 585
R1228 B.n804 B.n803 585
R1229 B.n805 B.n50 585
R1230 B.n807 B.n806 585
R1231 B.n808 B.n49 585
R1232 B.n810 B.n809 585
R1233 B.n811 B.n48 585
R1234 B.n813 B.n812 585
R1235 B.n814 B.n47 585
R1236 B.n816 B.n815 585
R1237 B.n817 B.n46 585
R1238 B.n819 B.n818 585
R1239 B.n820 B.n45 585
R1240 B.n822 B.n821 585
R1241 B.n823 B.n44 585
R1242 B.n825 B.n824 585
R1243 B.n826 B.n43 585
R1244 B.n828 B.n827 585
R1245 B.n829 B.n42 585
R1246 B.n831 B.n830 585
R1247 B.n832 B.n41 585
R1248 B.n834 B.n833 585
R1249 B.n835 B.n40 585
R1250 B.n837 B.n836 585
R1251 B.n838 B.n39 585
R1252 B.n840 B.n839 585
R1253 B.n841 B.n38 585
R1254 B.n843 B.n842 585
R1255 B.n844 B.n37 585
R1256 B.n846 B.n845 585
R1257 B.n847 B.n36 585
R1258 B.n849 B.n848 585
R1259 B.n850 B.n35 585
R1260 B.n852 B.n851 585
R1261 B.n853 B.n34 585
R1262 B.n855 B.n854 585
R1263 B.n691 B.n92 585
R1264 B.n690 B.n689 585
R1265 B.n688 B.n93 585
R1266 B.n687 B.n686 585
R1267 B.n685 B.n94 585
R1268 B.n684 B.n683 585
R1269 B.n682 B.n95 585
R1270 B.n681 B.n680 585
R1271 B.n679 B.n96 585
R1272 B.n678 B.n677 585
R1273 B.n676 B.n97 585
R1274 B.n675 B.n674 585
R1275 B.n673 B.n98 585
R1276 B.n672 B.n671 585
R1277 B.n670 B.n99 585
R1278 B.n669 B.n668 585
R1279 B.n667 B.n100 585
R1280 B.n666 B.n665 585
R1281 B.n664 B.n101 585
R1282 B.n663 B.n662 585
R1283 B.n661 B.n102 585
R1284 B.n660 B.n659 585
R1285 B.n658 B.n103 585
R1286 B.n657 B.n656 585
R1287 B.n655 B.n104 585
R1288 B.n654 B.n653 585
R1289 B.n652 B.n105 585
R1290 B.n651 B.n650 585
R1291 B.n649 B.n106 585
R1292 B.n648 B.n647 585
R1293 B.n646 B.n107 585
R1294 B.n645 B.n644 585
R1295 B.n643 B.n108 585
R1296 B.n642 B.n641 585
R1297 B.n640 B.n109 585
R1298 B.n639 B.n638 585
R1299 B.n637 B.n110 585
R1300 B.n636 B.n635 585
R1301 B.n634 B.n111 585
R1302 B.n633 B.n632 585
R1303 B.n631 B.n112 585
R1304 B.n630 B.n629 585
R1305 B.n628 B.n113 585
R1306 B.n627 B.n626 585
R1307 B.n625 B.n114 585
R1308 B.n624 B.n623 585
R1309 B.n622 B.n115 585
R1310 B.n621 B.n620 585
R1311 B.n619 B.n116 585
R1312 B.n618 B.n617 585
R1313 B.n616 B.n117 585
R1314 B.n615 B.n614 585
R1315 B.n613 B.n118 585
R1316 B.n612 B.n611 585
R1317 B.n610 B.n119 585
R1318 B.n609 B.n608 585
R1319 B.n607 B.n120 585
R1320 B.n606 B.n605 585
R1321 B.n604 B.n121 585
R1322 B.n603 B.n602 585
R1323 B.n601 B.n122 585
R1324 B.n600 B.n599 585
R1325 B.n598 B.n123 585
R1326 B.n597 B.n596 585
R1327 B.n595 B.n124 585
R1328 B.n594 B.n593 585
R1329 B.n592 B.n125 585
R1330 B.n591 B.n590 585
R1331 B.n589 B.n126 585
R1332 B.n588 B.n587 585
R1333 B.n586 B.n127 585
R1334 B.n585 B.n584 585
R1335 B.n583 B.n128 585
R1336 B.n582 B.n581 585
R1337 B.n580 B.n129 585
R1338 B.n579 B.n578 585
R1339 B.n577 B.n130 585
R1340 B.n576 B.n575 585
R1341 B.n574 B.n131 585
R1342 B.n573 B.n572 585
R1343 B.n571 B.n132 585
R1344 B.n570 B.n569 585
R1345 B.n568 B.n133 585
R1346 B.n567 B.n566 585
R1347 B.n565 B.n134 585
R1348 B.n564 B.n563 585
R1349 B.n562 B.n135 585
R1350 B.n561 B.n560 585
R1351 B.n559 B.n136 585
R1352 B.n558 B.n557 585
R1353 B.n556 B.n137 585
R1354 B.n555 B.n554 585
R1355 B.n553 B.n138 585
R1356 B.n552 B.n551 585
R1357 B.n550 B.n139 585
R1358 B.n549 B.n548 585
R1359 B.n547 B.n140 585
R1360 B.n546 B.n545 585
R1361 B.n544 B.n141 585
R1362 B.n543 B.n542 585
R1363 B.n541 B.n142 585
R1364 B.n540 B.n539 585
R1365 B.n538 B.n143 585
R1366 B.n537 B.n536 585
R1367 B.n535 B.n144 585
R1368 B.n534 B.n533 585
R1369 B.n532 B.n145 585
R1370 B.n531 B.n530 585
R1371 B.n529 B.n146 585
R1372 B.n528 B.n527 585
R1373 B.n526 B.n147 585
R1374 B.n525 B.n524 585
R1375 B.n523 B.n148 585
R1376 B.n522 B.n521 585
R1377 B.n520 B.n149 585
R1378 B.n519 B.n518 585
R1379 B.n517 B.n150 585
R1380 B.n516 B.n515 585
R1381 B.n514 B.n151 585
R1382 B.n513 B.n512 585
R1383 B.n511 B.n152 585
R1384 B.n510 B.n509 585
R1385 B.n508 B.n153 585
R1386 B.n507 B.n506 585
R1387 B.n505 B.n154 585
R1388 B.n504 B.n503 585
R1389 B.n502 B.n155 585
R1390 B.n339 B.n338 585
R1391 B.n340 B.n213 585
R1392 B.n342 B.n341 585
R1393 B.n343 B.n212 585
R1394 B.n345 B.n344 585
R1395 B.n346 B.n211 585
R1396 B.n348 B.n347 585
R1397 B.n349 B.n210 585
R1398 B.n351 B.n350 585
R1399 B.n352 B.n209 585
R1400 B.n354 B.n353 585
R1401 B.n355 B.n208 585
R1402 B.n357 B.n356 585
R1403 B.n358 B.n207 585
R1404 B.n360 B.n359 585
R1405 B.n361 B.n206 585
R1406 B.n363 B.n362 585
R1407 B.n364 B.n205 585
R1408 B.n366 B.n365 585
R1409 B.n367 B.n204 585
R1410 B.n369 B.n368 585
R1411 B.n370 B.n203 585
R1412 B.n372 B.n371 585
R1413 B.n373 B.n202 585
R1414 B.n375 B.n374 585
R1415 B.n376 B.n201 585
R1416 B.n378 B.n377 585
R1417 B.n379 B.n200 585
R1418 B.n381 B.n380 585
R1419 B.n382 B.n199 585
R1420 B.n384 B.n383 585
R1421 B.n385 B.n198 585
R1422 B.n387 B.n386 585
R1423 B.n388 B.n197 585
R1424 B.n390 B.n389 585
R1425 B.n391 B.n196 585
R1426 B.n393 B.n392 585
R1427 B.n394 B.n195 585
R1428 B.n396 B.n395 585
R1429 B.n397 B.n194 585
R1430 B.n399 B.n398 585
R1431 B.n400 B.n193 585
R1432 B.n402 B.n401 585
R1433 B.n403 B.n192 585
R1434 B.n405 B.n404 585
R1435 B.n406 B.n191 585
R1436 B.n408 B.n407 585
R1437 B.n409 B.n190 585
R1438 B.n411 B.n410 585
R1439 B.n413 B.n187 585
R1440 B.n415 B.n414 585
R1441 B.n416 B.n186 585
R1442 B.n418 B.n417 585
R1443 B.n419 B.n185 585
R1444 B.n421 B.n420 585
R1445 B.n422 B.n184 585
R1446 B.n424 B.n423 585
R1447 B.n425 B.n183 585
R1448 B.n427 B.n426 585
R1449 B.n429 B.n428 585
R1450 B.n430 B.n179 585
R1451 B.n432 B.n431 585
R1452 B.n433 B.n178 585
R1453 B.n435 B.n434 585
R1454 B.n436 B.n177 585
R1455 B.n438 B.n437 585
R1456 B.n439 B.n176 585
R1457 B.n441 B.n440 585
R1458 B.n442 B.n175 585
R1459 B.n444 B.n443 585
R1460 B.n445 B.n174 585
R1461 B.n447 B.n446 585
R1462 B.n448 B.n173 585
R1463 B.n450 B.n449 585
R1464 B.n451 B.n172 585
R1465 B.n453 B.n452 585
R1466 B.n454 B.n171 585
R1467 B.n456 B.n455 585
R1468 B.n457 B.n170 585
R1469 B.n459 B.n458 585
R1470 B.n460 B.n169 585
R1471 B.n462 B.n461 585
R1472 B.n463 B.n168 585
R1473 B.n465 B.n464 585
R1474 B.n466 B.n167 585
R1475 B.n468 B.n467 585
R1476 B.n469 B.n166 585
R1477 B.n471 B.n470 585
R1478 B.n472 B.n165 585
R1479 B.n474 B.n473 585
R1480 B.n475 B.n164 585
R1481 B.n477 B.n476 585
R1482 B.n478 B.n163 585
R1483 B.n480 B.n479 585
R1484 B.n481 B.n162 585
R1485 B.n483 B.n482 585
R1486 B.n484 B.n161 585
R1487 B.n486 B.n485 585
R1488 B.n487 B.n160 585
R1489 B.n489 B.n488 585
R1490 B.n490 B.n159 585
R1491 B.n492 B.n491 585
R1492 B.n493 B.n158 585
R1493 B.n495 B.n494 585
R1494 B.n496 B.n157 585
R1495 B.n498 B.n497 585
R1496 B.n499 B.n156 585
R1497 B.n501 B.n500 585
R1498 B.n337 B.n214 585
R1499 B.n336 B.n335 585
R1500 B.n334 B.n215 585
R1501 B.n333 B.n332 585
R1502 B.n331 B.n216 585
R1503 B.n330 B.n329 585
R1504 B.n328 B.n217 585
R1505 B.n327 B.n326 585
R1506 B.n325 B.n218 585
R1507 B.n324 B.n323 585
R1508 B.n322 B.n219 585
R1509 B.n321 B.n320 585
R1510 B.n319 B.n220 585
R1511 B.n318 B.n317 585
R1512 B.n316 B.n221 585
R1513 B.n315 B.n314 585
R1514 B.n313 B.n222 585
R1515 B.n312 B.n311 585
R1516 B.n310 B.n223 585
R1517 B.n309 B.n308 585
R1518 B.n307 B.n224 585
R1519 B.n306 B.n305 585
R1520 B.n304 B.n225 585
R1521 B.n303 B.n302 585
R1522 B.n301 B.n226 585
R1523 B.n300 B.n299 585
R1524 B.n298 B.n227 585
R1525 B.n297 B.n296 585
R1526 B.n295 B.n228 585
R1527 B.n294 B.n293 585
R1528 B.n292 B.n229 585
R1529 B.n291 B.n290 585
R1530 B.n289 B.n230 585
R1531 B.n288 B.n287 585
R1532 B.n286 B.n231 585
R1533 B.n285 B.n284 585
R1534 B.n283 B.n232 585
R1535 B.n282 B.n281 585
R1536 B.n280 B.n233 585
R1537 B.n279 B.n278 585
R1538 B.n277 B.n234 585
R1539 B.n276 B.n275 585
R1540 B.n274 B.n235 585
R1541 B.n273 B.n272 585
R1542 B.n271 B.n236 585
R1543 B.n270 B.n269 585
R1544 B.n268 B.n237 585
R1545 B.n267 B.n266 585
R1546 B.n265 B.n238 585
R1547 B.n264 B.n263 585
R1548 B.n262 B.n239 585
R1549 B.n261 B.n260 585
R1550 B.n259 B.n240 585
R1551 B.n258 B.n257 585
R1552 B.n256 B.n241 585
R1553 B.n255 B.n254 585
R1554 B.n253 B.n242 585
R1555 B.n252 B.n251 585
R1556 B.n250 B.n243 585
R1557 B.n249 B.n248 585
R1558 B.n247 B.n244 585
R1559 B.n246 B.n245 585
R1560 B.n2 B.n0 585
R1561 B.n949 B.n1 585
R1562 B.n948 B.n947 585
R1563 B.n946 B.n3 585
R1564 B.n945 B.n944 585
R1565 B.n943 B.n4 585
R1566 B.n942 B.n941 585
R1567 B.n940 B.n5 585
R1568 B.n939 B.n938 585
R1569 B.n937 B.n6 585
R1570 B.n936 B.n935 585
R1571 B.n934 B.n7 585
R1572 B.n933 B.n932 585
R1573 B.n931 B.n8 585
R1574 B.n930 B.n929 585
R1575 B.n928 B.n9 585
R1576 B.n927 B.n926 585
R1577 B.n925 B.n10 585
R1578 B.n924 B.n923 585
R1579 B.n922 B.n11 585
R1580 B.n921 B.n920 585
R1581 B.n919 B.n12 585
R1582 B.n918 B.n917 585
R1583 B.n916 B.n13 585
R1584 B.n915 B.n914 585
R1585 B.n913 B.n14 585
R1586 B.n912 B.n911 585
R1587 B.n910 B.n15 585
R1588 B.n909 B.n908 585
R1589 B.n907 B.n16 585
R1590 B.n906 B.n905 585
R1591 B.n904 B.n17 585
R1592 B.n903 B.n902 585
R1593 B.n901 B.n18 585
R1594 B.n900 B.n899 585
R1595 B.n898 B.n19 585
R1596 B.n897 B.n896 585
R1597 B.n895 B.n20 585
R1598 B.n894 B.n893 585
R1599 B.n892 B.n21 585
R1600 B.n891 B.n890 585
R1601 B.n889 B.n22 585
R1602 B.n888 B.n887 585
R1603 B.n886 B.n23 585
R1604 B.n885 B.n884 585
R1605 B.n883 B.n24 585
R1606 B.n882 B.n881 585
R1607 B.n880 B.n25 585
R1608 B.n879 B.n878 585
R1609 B.n877 B.n26 585
R1610 B.n876 B.n875 585
R1611 B.n874 B.n27 585
R1612 B.n873 B.n872 585
R1613 B.n871 B.n28 585
R1614 B.n870 B.n869 585
R1615 B.n868 B.n29 585
R1616 B.n867 B.n866 585
R1617 B.n865 B.n30 585
R1618 B.n864 B.n863 585
R1619 B.n862 B.n31 585
R1620 B.n861 B.n860 585
R1621 B.n859 B.n32 585
R1622 B.n858 B.n857 585
R1623 B.n856 B.n33 585
R1624 B.n951 B.n950 585
R1625 B.n338 B.n337 526.135
R1626 B.n854 B.n33 526.135
R1627 B.n500 B.n155 526.135
R1628 B.n692 B.n691 526.135
R1629 B.n180 B.t11 495.502
R1630 B.n66 B.t7 495.502
R1631 B.n188 B.t2 495.502
R1632 B.n58 B.t4 495.502
R1633 B.n181 B.t10 423.163
R1634 B.n67 B.t8 423.163
R1635 B.n189 B.t1 423.163
R1636 B.n59 B.t5 423.163
R1637 B.n180 B.t9 312.844
R1638 B.n188 B.t0 312.844
R1639 B.n58 B.t3 312.844
R1640 B.n66 B.t6 312.844
R1641 B.n337 B.n336 163.367
R1642 B.n336 B.n215 163.367
R1643 B.n332 B.n215 163.367
R1644 B.n332 B.n331 163.367
R1645 B.n331 B.n330 163.367
R1646 B.n330 B.n217 163.367
R1647 B.n326 B.n217 163.367
R1648 B.n326 B.n325 163.367
R1649 B.n325 B.n324 163.367
R1650 B.n324 B.n219 163.367
R1651 B.n320 B.n219 163.367
R1652 B.n320 B.n319 163.367
R1653 B.n319 B.n318 163.367
R1654 B.n318 B.n221 163.367
R1655 B.n314 B.n221 163.367
R1656 B.n314 B.n313 163.367
R1657 B.n313 B.n312 163.367
R1658 B.n312 B.n223 163.367
R1659 B.n308 B.n223 163.367
R1660 B.n308 B.n307 163.367
R1661 B.n307 B.n306 163.367
R1662 B.n306 B.n225 163.367
R1663 B.n302 B.n225 163.367
R1664 B.n302 B.n301 163.367
R1665 B.n301 B.n300 163.367
R1666 B.n300 B.n227 163.367
R1667 B.n296 B.n227 163.367
R1668 B.n296 B.n295 163.367
R1669 B.n295 B.n294 163.367
R1670 B.n294 B.n229 163.367
R1671 B.n290 B.n229 163.367
R1672 B.n290 B.n289 163.367
R1673 B.n289 B.n288 163.367
R1674 B.n288 B.n231 163.367
R1675 B.n284 B.n231 163.367
R1676 B.n284 B.n283 163.367
R1677 B.n283 B.n282 163.367
R1678 B.n282 B.n233 163.367
R1679 B.n278 B.n233 163.367
R1680 B.n278 B.n277 163.367
R1681 B.n277 B.n276 163.367
R1682 B.n276 B.n235 163.367
R1683 B.n272 B.n235 163.367
R1684 B.n272 B.n271 163.367
R1685 B.n271 B.n270 163.367
R1686 B.n270 B.n237 163.367
R1687 B.n266 B.n237 163.367
R1688 B.n266 B.n265 163.367
R1689 B.n265 B.n264 163.367
R1690 B.n264 B.n239 163.367
R1691 B.n260 B.n239 163.367
R1692 B.n260 B.n259 163.367
R1693 B.n259 B.n258 163.367
R1694 B.n258 B.n241 163.367
R1695 B.n254 B.n241 163.367
R1696 B.n254 B.n253 163.367
R1697 B.n253 B.n252 163.367
R1698 B.n252 B.n243 163.367
R1699 B.n248 B.n243 163.367
R1700 B.n248 B.n247 163.367
R1701 B.n247 B.n246 163.367
R1702 B.n246 B.n2 163.367
R1703 B.n950 B.n2 163.367
R1704 B.n950 B.n949 163.367
R1705 B.n949 B.n948 163.367
R1706 B.n948 B.n3 163.367
R1707 B.n944 B.n3 163.367
R1708 B.n944 B.n943 163.367
R1709 B.n943 B.n942 163.367
R1710 B.n942 B.n5 163.367
R1711 B.n938 B.n5 163.367
R1712 B.n938 B.n937 163.367
R1713 B.n937 B.n936 163.367
R1714 B.n936 B.n7 163.367
R1715 B.n932 B.n7 163.367
R1716 B.n932 B.n931 163.367
R1717 B.n931 B.n930 163.367
R1718 B.n930 B.n9 163.367
R1719 B.n926 B.n9 163.367
R1720 B.n926 B.n925 163.367
R1721 B.n925 B.n924 163.367
R1722 B.n924 B.n11 163.367
R1723 B.n920 B.n11 163.367
R1724 B.n920 B.n919 163.367
R1725 B.n919 B.n918 163.367
R1726 B.n918 B.n13 163.367
R1727 B.n914 B.n13 163.367
R1728 B.n914 B.n913 163.367
R1729 B.n913 B.n912 163.367
R1730 B.n912 B.n15 163.367
R1731 B.n908 B.n15 163.367
R1732 B.n908 B.n907 163.367
R1733 B.n907 B.n906 163.367
R1734 B.n906 B.n17 163.367
R1735 B.n902 B.n17 163.367
R1736 B.n902 B.n901 163.367
R1737 B.n901 B.n900 163.367
R1738 B.n900 B.n19 163.367
R1739 B.n896 B.n19 163.367
R1740 B.n896 B.n895 163.367
R1741 B.n895 B.n894 163.367
R1742 B.n894 B.n21 163.367
R1743 B.n890 B.n21 163.367
R1744 B.n890 B.n889 163.367
R1745 B.n889 B.n888 163.367
R1746 B.n888 B.n23 163.367
R1747 B.n884 B.n23 163.367
R1748 B.n884 B.n883 163.367
R1749 B.n883 B.n882 163.367
R1750 B.n882 B.n25 163.367
R1751 B.n878 B.n25 163.367
R1752 B.n878 B.n877 163.367
R1753 B.n877 B.n876 163.367
R1754 B.n876 B.n27 163.367
R1755 B.n872 B.n27 163.367
R1756 B.n872 B.n871 163.367
R1757 B.n871 B.n870 163.367
R1758 B.n870 B.n29 163.367
R1759 B.n866 B.n29 163.367
R1760 B.n866 B.n865 163.367
R1761 B.n865 B.n864 163.367
R1762 B.n864 B.n31 163.367
R1763 B.n860 B.n31 163.367
R1764 B.n860 B.n859 163.367
R1765 B.n859 B.n858 163.367
R1766 B.n858 B.n33 163.367
R1767 B.n338 B.n213 163.367
R1768 B.n342 B.n213 163.367
R1769 B.n343 B.n342 163.367
R1770 B.n344 B.n343 163.367
R1771 B.n344 B.n211 163.367
R1772 B.n348 B.n211 163.367
R1773 B.n349 B.n348 163.367
R1774 B.n350 B.n349 163.367
R1775 B.n350 B.n209 163.367
R1776 B.n354 B.n209 163.367
R1777 B.n355 B.n354 163.367
R1778 B.n356 B.n355 163.367
R1779 B.n356 B.n207 163.367
R1780 B.n360 B.n207 163.367
R1781 B.n361 B.n360 163.367
R1782 B.n362 B.n361 163.367
R1783 B.n362 B.n205 163.367
R1784 B.n366 B.n205 163.367
R1785 B.n367 B.n366 163.367
R1786 B.n368 B.n367 163.367
R1787 B.n368 B.n203 163.367
R1788 B.n372 B.n203 163.367
R1789 B.n373 B.n372 163.367
R1790 B.n374 B.n373 163.367
R1791 B.n374 B.n201 163.367
R1792 B.n378 B.n201 163.367
R1793 B.n379 B.n378 163.367
R1794 B.n380 B.n379 163.367
R1795 B.n380 B.n199 163.367
R1796 B.n384 B.n199 163.367
R1797 B.n385 B.n384 163.367
R1798 B.n386 B.n385 163.367
R1799 B.n386 B.n197 163.367
R1800 B.n390 B.n197 163.367
R1801 B.n391 B.n390 163.367
R1802 B.n392 B.n391 163.367
R1803 B.n392 B.n195 163.367
R1804 B.n396 B.n195 163.367
R1805 B.n397 B.n396 163.367
R1806 B.n398 B.n397 163.367
R1807 B.n398 B.n193 163.367
R1808 B.n402 B.n193 163.367
R1809 B.n403 B.n402 163.367
R1810 B.n404 B.n403 163.367
R1811 B.n404 B.n191 163.367
R1812 B.n408 B.n191 163.367
R1813 B.n409 B.n408 163.367
R1814 B.n410 B.n409 163.367
R1815 B.n410 B.n187 163.367
R1816 B.n415 B.n187 163.367
R1817 B.n416 B.n415 163.367
R1818 B.n417 B.n416 163.367
R1819 B.n417 B.n185 163.367
R1820 B.n421 B.n185 163.367
R1821 B.n422 B.n421 163.367
R1822 B.n423 B.n422 163.367
R1823 B.n423 B.n183 163.367
R1824 B.n427 B.n183 163.367
R1825 B.n428 B.n427 163.367
R1826 B.n428 B.n179 163.367
R1827 B.n432 B.n179 163.367
R1828 B.n433 B.n432 163.367
R1829 B.n434 B.n433 163.367
R1830 B.n434 B.n177 163.367
R1831 B.n438 B.n177 163.367
R1832 B.n439 B.n438 163.367
R1833 B.n440 B.n439 163.367
R1834 B.n440 B.n175 163.367
R1835 B.n444 B.n175 163.367
R1836 B.n445 B.n444 163.367
R1837 B.n446 B.n445 163.367
R1838 B.n446 B.n173 163.367
R1839 B.n450 B.n173 163.367
R1840 B.n451 B.n450 163.367
R1841 B.n452 B.n451 163.367
R1842 B.n452 B.n171 163.367
R1843 B.n456 B.n171 163.367
R1844 B.n457 B.n456 163.367
R1845 B.n458 B.n457 163.367
R1846 B.n458 B.n169 163.367
R1847 B.n462 B.n169 163.367
R1848 B.n463 B.n462 163.367
R1849 B.n464 B.n463 163.367
R1850 B.n464 B.n167 163.367
R1851 B.n468 B.n167 163.367
R1852 B.n469 B.n468 163.367
R1853 B.n470 B.n469 163.367
R1854 B.n470 B.n165 163.367
R1855 B.n474 B.n165 163.367
R1856 B.n475 B.n474 163.367
R1857 B.n476 B.n475 163.367
R1858 B.n476 B.n163 163.367
R1859 B.n480 B.n163 163.367
R1860 B.n481 B.n480 163.367
R1861 B.n482 B.n481 163.367
R1862 B.n482 B.n161 163.367
R1863 B.n486 B.n161 163.367
R1864 B.n487 B.n486 163.367
R1865 B.n488 B.n487 163.367
R1866 B.n488 B.n159 163.367
R1867 B.n492 B.n159 163.367
R1868 B.n493 B.n492 163.367
R1869 B.n494 B.n493 163.367
R1870 B.n494 B.n157 163.367
R1871 B.n498 B.n157 163.367
R1872 B.n499 B.n498 163.367
R1873 B.n500 B.n499 163.367
R1874 B.n504 B.n155 163.367
R1875 B.n505 B.n504 163.367
R1876 B.n506 B.n505 163.367
R1877 B.n506 B.n153 163.367
R1878 B.n510 B.n153 163.367
R1879 B.n511 B.n510 163.367
R1880 B.n512 B.n511 163.367
R1881 B.n512 B.n151 163.367
R1882 B.n516 B.n151 163.367
R1883 B.n517 B.n516 163.367
R1884 B.n518 B.n517 163.367
R1885 B.n518 B.n149 163.367
R1886 B.n522 B.n149 163.367
R1887 B.n523 B.n522 163.367
R1888 B.n524 B.n523 163.367
R1889 B.n524 B.n147 163.367
R1890 B.n528 B.n147 163.367
R1891 B.n529 B.n528 163.367
R1892 B.n530 B.n529 163.367
R1893 B.n530 B.n145 163.367
R1894 B.n534 B.n145 163.367
R1895 B.n535 B.n534 163.367
R1896 B.n536 B.n535 163.367
R1897 B.n536 B.n143 163.367
R1898 B.n540 B.n143 163.367
R1899 B.n541 B.n540 163.367
R1900 B.n542 B.n541 163.367
R1901 B.n542 B.n141 163.367
R1902 B.n546 B.n141 163.367
R1903 B.n547 B.n546 163.367
R1904 B.n548 B.n547 163.367
R1905 B.n548 B.n139 163.367
R1906 B.n552 B.n139 163.367
R1907 B.n553 B.n552 163.367
R1908 B.n554 B.n553 163.367
R1909 B.n554 B.n137 163.367
R1910 B.n558 B.n137 163.367
R1911 B.n559 B.n558 163.367
R1912 B.n560 B.n559 163.367
R1913 B.n560 B.n135 163.367
R1914 B.n564 B.n135 163.367
R1915 B.n565 B.n564 163.367
R1916 B.n566 B.n565 163.367
R1917 B.n566 B.n133 163.367
R1918 B.n570 B.n133 163.367
R1919 B.n571 B.n570 163.367
R1920 B.n572 B.n571 163.367
R1921 B.n572 B.n131 163.367
R1922 B.n576 B.n131 163.367
R1923 B.n577 B.n576 163.367
R1924 B.n578 B.n577 163.367
R1925 B.n578 B.n129 163.367
R1926 B.n582 B.n129 163.367
R1927 B.n583 B.n582 163.367
R1928 B.n584 B.n583 163.367
R1929 B.n584 B.n127 163.367
R1930 B.n588 B.n127 163.367
R1931 B.n589 B.n588 163.367
R1932 B.n590 B.n589 163.367
R1933 B.n590 B.n125 163.367
R1934 B.n594 B.n125 163.367
R1935 B.n595 B.n594 163.367
R1936 B.n596 B.n595 163.367
R1937 B.n596 B.n123 163.367
R1938 B.n600 B.n123 163.367
R1939 B.n601 B.n600 163.367
R1940 B.n602 B.n601 163.367
R1941 B.n602 B.n121 163.367
R1942 B.n606 B.n121 163.367
R1943 B.n607 B.n606 163.367
R1944 B.n608 B.n607 163.367
R1945 B.n608 B.n119 163.367
R1946 B.n612 B.n119 163.367
R1947 B.n613 B.n612 163.367
R1948 B.n614 B.n613 163.367
R1949 B.n614 B.n117 163.367
R1950 B.n618 B.n117 163.367
R1951 B.n619 B.n618 163.367
R1952 B.n620 B.n619 163.367
R1953 B.n620 B.n115 163.367
R1954 B.n624 B.n115 163.367
R1955 B.n625 B.n624 163.367
R1956 B.n626 B.n625 163.367
R1957 B.n626 B.n113 163.367
R1958 B.n630 B.n113 163.367
R1959 B.n631 B.n630 163.367
R1960 B.n632 B.n631 163.367
R1961 B.n632 B.n111 163.367
R1962 B.n636 B.n111 163.367
R1963 B.n637 B.n636 163.367
R1964 B.n638 B.n637 163.367
R1965 B.n638 B.n109 163.367
R1966 B.n642 B.n109 163.367
R1967 B.n643 B.n642 163.367
R1968 B.n644 B.n643 163.367
R1969 B.n644 B.n107 163.367
R1970 B.n648 B.n107 163.367
R1971 B.n649 B.n648 163.367
R1972 B.n650 B.n649 163.367
R1973 B.n650 B.n105 163.367
R1974 B.n654 B.n105 163.367
R1975 B.n655 B.n654 163.367
R1976 B.n656 B.n655 163.367
R1977 B.n656 B.n103 163.367
R1978 B.n660 B.n103 163.367
R1979 B.n661 B.n660 163.367
R1980 B.n662 B.n661 163.367
R1981 B.n662 B.n101 163.367
R1982 B.n666 B.n101 163.367
R1983 B.n667 B.n666 163.367
R1984 B.n668 B.n667 163.367
R1985 B.n668 B.n99 163.367
R1986 B.n672 B.n99 163.367
R1987 B.n673 B.n672 163.367
R1988 B.n674 B.n673 163.367
R1989 B.n674 B.n97 163.367
R1990 B.n678 B.n97 163.367
R1991 B.n679 B.n678 163.367
R1992 B.n680 B.n679 163.367
R1993 B.n680 B.n95 163.367
R1994 B.n684 B.n95 163.367
R1995 B.n685 B.n684 163.367
R1996 B.n686 B.n685 163.367
R1997 B.n686 B.n93 163.367
R1998 B.n690 B.n93 163.367
R1999 B.n691 B.n690 163.367
R2000 B.n854 B.n853 163.367
R2001 B.n853 B.n852 163.367
R2002 B.n852 B.n35 163.367
R2003 B.n848 B.n35 163.367
R2004 B.n848 B.n847 163.367
R2005 B.n847 B.n846 163.367
R2006 B.n846 B.n37 163.367
R2007 B.n842 B.n37 163.367
R2008 B.n842 B.n841 163.367
R2009 B.n841 B.n840 163.367
R2010 B.n840 B.n39 163.367
R2011 B.n836 B.n39 163.367
R2012 B.n836 B.n835 163.367
R2013 B.n835 B.n834 163.367
R2014 B.n834 B.n41 163.367
R2015 B.n830 B.n41 163.367
R2016 B.n830 B.n829 163.367
R2017 B.n829 B.n828 163.367
R2018 B.n828 B.n43 163.367
R2019 B.n824 B.n43 163.367
R2020 B.n824 B.n823 163.367
R2021 B.n823 B.n822 163.367
R2022 B.n822 B.n45 163.367
R2023 B.n818 B.n45 163.367
R2024 B.n818 B.n817 163.367
R2025 B.n817 B.n816 163.367
R2026 B.n816 B.n47 163.367
R2027 B.n812 B.n47 163.367
R2028 B.n812 B.n811 163.367
R2029 B.n811 B.n810 163.367
R2030 B.n810 B.n49 163.367
R2031 B.n806 B.n49 163.367
R2032 B.n806 B.n805 163.367
R2033 B.n805 B.n804 163.367
R2034 B.n804 B.n51 163.367
R2035 B.n800 B.n51 163.367
R2036 B.n800 B.n799 163.367
R2037 B.n799 B.n798 163.367
R2038 B.n798 B.n53 163.367
R2039 B.n794 B.n53 163.367
R2040 B.n794 B.n793 163.367
R2041 B.n793 B.n792 163.367
R2042 B.n792 B.n55 163.367
R2043 B.n788 B.n55 163.367
R2044 B.n788 B.n787 163.367
R2045 B.n787 B.n786 163.367
R2046 B.n786 B.n57 163.367
R2047 B.n782 B.n57 163.367
R2048 B.n782 B.n781 163.367
R2049 B.n781 B.n61 163.367
R2050 B.n777 B.n61 163.367
R2051 B.n777 B.n776 163.367
R2052 B.n776 B.n775 163.367
R2053 B.n775 B.n63 163.367
R2054 B.n771 B.n63 163.367
R2055 B.n771 B.n770 163.367
R2056 B.n770 B.n769 163.367
R2057 B.n769 B.n65 163.367
R2058 B.n764 B.n65 163.367
R2059 B.n764 B.n763 163.367
R2060 B.n763 B.n762 163.367
R2061 B.n762 B.n69 163.367
R2062 B.n758 B.n69 163.367
R2063 B.n758 B.n757 163.367
R2064 B.n757 B.n756 163.367
R2065 B.n756 B.n71 163.367
R2066 B.n752 B.n71 163.367
R2067 B.n752 B.n751 163.367
R2068 B.n751 B.n750 163.367
R2069 B.n750 B.n73 163.367
R2070 B.n746 B.n73 163.367
R2071 B.n746 B.n745 163.367
R2072 B.n745 B.n744 163.367
R2073 B.n744 B.n75 163.367
R2074 B.n740 B.n75 163.367
R2075 B.n740 B.n739 163.367
R2076 B.n739 B.n738 163.367
R2077 B.n738 B.n77 163.367
R2078 B.n734 B.n77 163.367
R2079 B.n734 B.n733 163.367
R2080 B.n733 B.n732 163.367
R2081 B.n732 B.n79 163.367
R2082 B.n728 B.n79 163.367
R2083 B.n728 B.n727 163.367
R2084 B.n727 B.n726 163.367
R2085 B.n726 B.n81 163.367
R2086 B.n722 B.n81 163.367
R2087 B.n722 B.n721 163.367
R2088 B.n721 B.n720 163.367
R2089 B.n720 B.n83 163.367
R2090 B.n716 B.n83 163.367
R2091 B.n716 B.n715 163.367
R2092 B.n715 B.n714 163.367
R2093 B.n714 B.n85 163.367
R2094 B.n710 B.n85 163.367
R2095 B.n710 B.n709 163.367
R2096 B.n709 B.n708 163.367
R2097 B.n708 B.n87 163.367
R2098 B.n704 B.n87 163.367
R2099 B.n704 B.n703 163.367
R2100 B.n703 B.n702 163.367
R2101 B.n702 B.n89 163.367
R2102 B.n698 B.n89 163.367
R2103 B.n698 B.n697 163.367
R2104 B.n697 B.n696 163.367
R2105 B.n696 B.n91 163.367
R2106 B.n692 B.n91 163.367
R2107 B.n181 B.n180 72.3399
R2108 B.n189 B.n188 72.3399
R2109 B.n59 B.n58 72.3399
R2110 B.n67 B.n66 72.3399
R2111 B.n182 B.n181 59.5399
R2112 B.n412 B.n189 59.5399
R2113 B.n60 B.n59 59.5399
R2114 B.n766 B.n67 59.5399
R2115 B.n856 B.n855 34.1859
R2116 B.n693 B.n92 34.1859
R2117 B.n502 B.n501 34.1859
R2118 B.n339 B.n214 34.1859
R2119 B B.n951 18.0485
R2120 B.n855 B.n34 10.6151
R2121 B.n851 B.n34 10.6151
R2122 B.n851 B.n850 10.6151
R2123 B.n850 B.n849 10.6151
R2124 B.n849 B.n36 10.6151
R2125 B.n845 B.n36 10.6151
R2126 B.n845 B.n844 10.6151
R2127 B.n844 B.n843 10.6151
R2128 B.n843 B.n38 10.6151
R2129 B.n839 B.n38 10.6151
R2130 B.n839 B.n838 10.6151
R2131 B.n838 B.n837 10.6151
R2132 B.n837 B.n40 10.6151
R2133 B.n833 B.n40 10.6151
R2134 B.n833 B.n832 10.6151
R2135 B.n832 B.n831 10.6151
R2136 B.n831 B.n42 10.6151
R2137 B.n827 B.n42 10.6151
R2138 B.n827 B.n826 10.6151
R2139 B.n826 B.n825 10.6151
R2140 B.n825 B.n44 10.6151
R2141 B.n821 B.n44 10.6151
R2142 B.n821 B.n820 10.6151
R2143 B.n820 B.n819 10.6151
R2144 B.n819 B.n46 10.6151
R2145 B.n815 B.n46 10.6151
R2146 B.n815 B.n814 10.6151
R2147 B.n814 B.n813 10.6151
R2148 B.n813 B.n48 10.6151
R2149 B.n809 B.n48 10.6151
R2150 B.n809 B.n808 10.6151
R2151 B.n808 B.n807 10.6151
R2152 B.n807 B.n50 10.6151
R2153 B.n803 B.n50 10.6151
R2154 B.n803 B.n802 10.6151
R2155 B.n802 B.n801 10.6151
R2156 B.n801 B.n52 10.6151
R2157 B.n797 B.n52 10.6151
R2158 B.n797 B.n796 10.6151
R2159 B.n796 B.n795 10.6151
R2160 B.n795 B.n54 10.6151
R2161 B.n791 B.n54 10.6151
R2162 B.n791 B.n790 10.6151
R2163 B.n790 B.n789 10.6151
R2164 B.n789 B.n56 10.6151
R2165 B.n785 B.n56 10.6151
R2166 B.n785 B.n784 10.6151
R2167 B.n784 B.n783 10.6151
R2168 B.n780 B.n779 10.6151
R2169 B.n779 B.n778 10.6151
R2170 B.n778 B.n62 10.6151
R2171 B.n774 B.n62 10.6151
R2172 B.n774 B.n773 10.6151
R2173 B.n773 B.n772 10.6151
R2174 B.n772 B.n64 10.6151
R2175 B.n768 B.n64 10.6151
R2176 B.n768 B.n767 10.6151
R2177 B.n765 B.n68 10.6151
R2178 B.n761 B.n68 10.6151
R2179 B.n761 B.n760 10.6151
R2180 B.n760 B.n759 10.6151
R2181 B.n759 B.n70 10.6151
R2182 B.n755 B.n70 10.6151
R2183 B.n755 B.n754 10.6151
R2184 B.n754 B.n753 10.6151
R2185 B.n753 B.n72 10.6151
R2186 B.n749 B.n72 10.6151
R2187 B.n749 B.n748 10.6151
R2188 B.n748 B.n747 10.6151
R2189 B.n747 B.n74 10.6151
R2190 B.n743 B.n74 10.6151
R2191 B.n743 B.n742 10.6151
R2192 B.n742 B.n741 10.6151
R2193 B.n741 B.n76 10.6151
R2194 B.n737 B.n76 10.6151
R2195 B.n737 B.n736 10.6151
R2196 B.n736 B.n735 10.6151
R2197 B.n735 B.n78 10.6151
R2198 B.n731 B.n78 10.6151
R2199 B.n731 B.n730 10.6151
R2200 B.n730 B.n729 10.6151
R2201 B.n729 B.n80 10.6151
R2202 B.n725 B.n80 10.6151
R2203 B.n725 B.n724 10.6151
R2204 B.n724 B.n723 10.6151
R2205 B.n723 B.n82 10.6151
R2206 B.n719 B.n82 10.6151
R2207 B.n719 B.n718 10.6151
R2208 B.n718 B.n717 10.6151
R2209 B.n717 B.n84 10.6151
R2210 B.n713 B.n84 10.6151
R2211 B.n713 B.n712 10.6151
R2212 B.n712 B.n711 10.6151
R2213 B.n711 B.n86 10.6151
R2214 B.n707 B.n86 10.6151
R2215 B.n707 B.n706 10.6151
R2216 B.n706 B.n705 10.6151
R2217 B.n705 B.n88 10.6151
R2218 B.n701 B.n88 10.6151
R2219 B.n701 B.n700 10.6151
R2220 B.n700 B.n699 10.6151
R2221 B.n699 B.n90 10.6151
R2222 B.n695 B.n90 10.6151
R2223 B.n695 B.n694 10.6151
R2224 B.n694 B.n693 10.6151
R2225 B.n503 B.n502 10.6151
R2226 B.n503 B.n154 10.6151
R2227 B.n507 B.n154 10.6151
R2228 B.n508 B.n507 10.6151
R2229 B.n509 B.n508 10.6151
R2230 B.n509 B.n152 10.6151
R2231 B.n513 B.n152 10.6151
R2232 B.n514 B.n513 10.6151
R2233 B.n515 B.n514 10.6151
R2234 B.n515 B.n150 10.6151
R2235 B.n519 B.n150 10.6151
R2236 B.n520 B.n519 10.6151
R2237 B.n521 B.n520 10.6151
R2238 B.n521 B.n148 10.6151
R2239 B.n525 B.n148 10.6151
R2240 B.n526 B.n525 10.6151
R2241 B.n527 B.n526 10.6151
R2242 B.n527 B.n146 10.6151
R2243 B.n531 B.n146 10.6151
R2244 B.n532 B.n531 10.6151
R2245 B.n533 B.n532 10.6151
R2246 B.n533 B.n144 10.6151
R2247 B.n537 B.n144 10.6151
R2248 B.n538 B.n537 10.6151
R2249 B.n539 B.n538 10.6151
R2250 B.n539 B.n142 10.6151
R2251 B.n543 B.n142 10.6151
R2252 B.n544 B.n543 10.6151
R2253 B.n545 B.n544 10.6151
R2254 B.n545 B.n140 10.6151
R2255 B.n549 B.n140 10.6151
R2256 B.n550 B.n549 10.6151
R2257 B.n551 B.n550 10.6151
R2258 B.n551 B.n138 10.6151
R2259 B.n555 B.n138 10.6151
R2260 B.n556 B.n555 10.6151
R2261 B.n557 B.n556 10.6151
R2262 B.n557 B.n136 10.6151
R2263 B.n561 B.n136 10.6151
R2264 B.n562 B.n561 10.6151
R2265 B.n563 B.n562 10.6151
R2266 B.n563 B.n134 10.6151
R2267 B.n567 B.n134 10.6151
R2268 B.n568 B.n567 10.6151
R2269 B.n569 B.n568 10.6151
R2270 B.n569 B.n132 10.6151
R2271 B.n573 B.n132 10.6151
R2272 B.n574 B.n573 10.6151
R2273 B.n575 B.n574 10.6151
R2274 B.n575 B.n130 10.6151
R2275 B.n579 B.n130 10.6151
R2276 B.n580 B.n579 10.6151
R2277 B.n581 B.n580 10.6151
R2278 B.n581 B.n128 10.6151
R2279 B.n585 B.n128 10.6151
R2280 B.n586 B.n585 10.6151
R2281 B.n587 B.n586 10.6151
R2282 B.n587 B.n126 10.6151
R2283 B.n591 B.n126 10.6151
R2284 B.n592 B.n591 10.6151
R2285 B.n593 B.n592 10.6151
R2286 B.n593 B.n124 10.6151
R2287 B.n597 B.n124 10.6151
R2288 B.n598 B.n597 10.6151
R2289 B.n599 B.n598 10.6151
R2290 B.n599 B.n122 10.6151
R2291 B.n603 B.n122 10.6151
R2292 B.n604 B.n603 10.6151
R2293 B.n605 B.n604 10.6151
R2294 B.n605 B.n120 10.6151
R2295 B.n609 B.n120 10.6151
R2296 B.n610 B.n609 10.6151
R2297 B.n611 B.n610 10.6151
R2298 B.n611 B.n118 10.6151
R2299 B.n615 B.n118 10.6151
R2300 B.n616 B.n615 10.6151
R2301 B.n617 B.n616 10.6151
R2302 B.n617 B.n116 10.6151
R2303 B.n621 B.n116 10.6151
R2304 B.n622 B.n621 10.6151
R2305 B.n623 B.n622 10.6151
R2306 B.n623 B.n114 10.6151
R2307 B.n627 B.n114 10.6151
R2308 B.n628 B.n627 10.6151
R2309 B.n629 B.n628 10.6151
R2310 B.n629 B.n112 10.6151
R2311 B.n633 B.n112 10.6151
R2312 B.n634 B.n633 10.6151
R2313 B.n635 B.n634 10.6151
R2314 B.n635 B.n110 10.6151
R2315 B.n639 B.n110 10.6151
R2316 B.n640 B.n639 10.6151
R2317 B.n641 B.n640 10.6151
R2318 B.n641 B.n108 10.6151
R2319 B.n645 B.n108 10.6151
R2320 B.n646 B.n645 10.6151
R2321 B.n647 B.n646 10.6151
R2322 B.n647 B.n106 10.6151
R2323 B.n651 B.n106 10.6151
R2324 B.n652 B.n651 10.6151
R2325 B.n653 B.n652 10.6151
R2326 B.n653 B.n104 10.6151
R2327 B.n657 B.n104 10.6151
R2328 B.n658 B.n657 10.6151
R2329 B.n659 B.n658 10.6151
R2330 B.n659 B.n102 10.6151
R2331 B.n663 B.n102 10.6151
R2332 B.n664 B.n663 10.6151
R2333 B.n665 B.n664 10.6151
R2334 B.n665 B.n100 10.6151
R2335 B.n669 B.n100 10.6151
R2336 B.n670 B.n669 10.6151
R2337 B.n671 B.n670 10.6151
R2338 B.n671 B.n98 10.6151
R2339 B.n675 B.n98 10.6151
R2340 B.n676 B.n675 10.6151
R2341 B.n677 B.n676 10.6151
R2342 B.n677 B.n96 10.6151
R2343 B.n681 B.n96 10.6151
R2344 B.n682 B.n681 10.6151
R2345 B.n683 B.n682 10.6151
R2346 B.n683 B.n94 10.6151
R2347 B.n687 B.n94 10.6151
R2348 B.n688 B.n687 10.6151
R2349 B.n689 B.n688 10.6151
R2350 B.n689 B.n92 10.6151
R2351 B.n340 B.n339 10.6151
R2352 B.n341 B.n340 10.6151
R2353 B.n341 B.n212 10.6151
R2354 B.n345 B.n212 10.6151
R2355 B.n346 B.n345 10.6151
R2356 B.n347 B.n346 10.6151
R2357 B.n347 B.n210 10.6151
R2358 B.n351 B.n210 10.6151
R2359 B.n352 B.n351 10.6151
R2360 B.n353 B.n352 10.6151
R2361 B.n353 B.n208 10.6151
R2362 B.n357 B.n208 10.6151
R2363 B.n358 B.n357 10.6151
R2364 B.n359 B.n358 10.6151
R2365 B.n359 B.n206 10.6151
R2366 B.n363 B.n206 10.6151
R2367 B.n364 B.n363 10.6151
R2368 B.n365 B.n364 10.6151
R2369 B.n365 B.n204 10.6151
R2370 B.n369 B.n204 10.6151
R2371 B.n370 B.n369 10.6151
R2372 B.n371 B.n370 10.6151
R2373 B.n371 B.n202 10.6151
R2374 B.n375 B.n202 10.6151
R2375 B.n376 B.n375 10.6151
R2376 B.n377 B.n376 10.6151
R2377 B.n377 B.n200 10.6151
R2378 B.n381 B.n200 10.6151
R2379 B.n382 B.n381 10.6151
R2380 B.n383 B.n382 10.6151
R2381 B.n383 B.n198 10.6151
R2382 B.n387 B.n198 10.6151
R2383 B.n388 B.n387 10.6151
R2384 B.n389 B.n388 10.6151
R2385 B.n389 B.n196 10.6151
R2386 B.n393 B.n196 10.6151
R2387 B.n394 B.n393 10.6151
R2388 B.n395 B.n394 10.6151
R2389 B.n395 B.n194 10.6151
R2390 B.n399 B.n194 10.6151
R2391 B.n400 B.n399 10.6151
R2392 B.n401 B.n400 10.6151
R2393 B.n401 B.n192 10.6151
R2394 B.n405 B.n192 10.6151
R2395 B.n406 B.n405 10.6151
R2396 B.n407 B.n406 10.6151
R2397 B.n407 B.n190 10.6151
R2398 B.n411 B.n190 10.6151
R2399 B.n414 B.n413 10.6151
R2400 B.n414 B.n186 10.6151
R2401 B.n418 B.n186 10.6151
R2402 B.n419 B.n418 10.6151
R2403 B.n420 B.n419 10.6151
R2404 B.n420 B.n184 10.6151
R2405 B.n424 B.n184 10.6151
R2406 B.n425 B.n424 10.6151
R2407 B.n426 B.n425 10.6151
R2408 B.n430 B.n429 10.6151
R2409 B.n431 B.n430 10.6151
R2410 B.n431 B.n178 10.6151
R2411 B.n435 B.n178 10.6151
R2412 B.n436 B.n435 10.6151
R2413 B.n437 B.n436 10.6151
R2414 B.n437 B.n176 10.6151
R2415 B.n441 B.n176 10.6151
R2416 B.n442 B.n441 10.6151
R2417 B.n443 B.n442 10.6151
R2418 B.n443 B.n174 10.6151
R2419 B.n447 B.n174 10.6151
R2420 B.n448 B.n447 10.6151
R2421 B.n449 B.n448 10.6151
R2422 B.n449 B.n172 10.6151
R2423 B.n453 B.n172 10.6151
R2424 B.n454 B.n453 10.6151
R2425 B.n455 B.n454 10.6151
R2426 B.n455 B.n170 10.6151
R2427 B.n459 B.n170 10.6151
R2428 B.n460 B.n459 10.6151
R2429 B.n461 B.n460 10.6151
R2430 B.n461 B.n168 10.6151
R2431 B.n465 B.n168 10.6151
R2432 B.n466 B.n465 10.6151
R2433 B.n467 B.n466 10.6151
R2434 B.n467 B.n166 10.6151
R2435 B.n471 B.n166 10.6151
R2436 B.n472 B.n471 10.6151
R2437 B.n473 B.n472 10.6151
R2438 B.n473 B.n164 10.6151
R2439 B.n477 B.n164 10.6151
R2440 B.n478 B.n477 10.6151
R2441 B.n479 B.n478 10.6151
R2442 B.n479 B.n162 10.6151
R2443 B.n483 B.n162 10.6151
R2444 B.n484 B.n483 10.6151
R2445 B.n485 B.n484 10.6151
R2446 B.n485 B.n160 10.6151
R2447 B.n489 B.n160 10.6151
R2448 B.n490 B.n489 10.6151
R2449 B.n491 B.n490 10.6151
R2450 B.n491 B.n158 10.6151
R2451 B.n495 B.n158 10.6151
R2452 B.n496 B.n495 10.6151
R2453 B.n497 B.n496 10.6151
R2454 B.n497 B.n156 10.6151
R2455 B.n501 B.n156 10.6151
R2456 B.n335 B.n214 10.6151
R2457 B.n335 B.n334 10.6151
R2458 B.n334 B.n333 10.6151
R2459 B.n333 B.n216 10.6151
R2460 B.n329 B.n216 10.6151
R2461 B.n329 B.n328 10.6151
R2462 B.n328 B.n327 10.6151
R2463 B.n327 B.n218 10.6151
R2464 B.n323 B.n218 10.6151
R2465 B.n323 B.n322 10.6151
R2466 B.n322 B.n321 10.6151
R2467 B.n321 B.n220 10.6151
R2468 B.n317 B.n220 10.6151
R2469 B.n317 B.n316 10.6151
R2470 B.n316 B.n315 10.6151
R2471 B.n315 B.n222 10.6151
R2472 B.n311 B.n222 10.6151
R2473 B.n311 B.n310 10.6151
R2474 B.n310 B.n309 10.6151
R2475 B.n309 B.n224 10.6151
R2476 B.n305 B.n224 10.6151
R2477 B.n305 B.n304 10.6151
R2478 B.n304 B.n303 10.6151
R2479 B.n303 B.n226 10.6151
R2480 B.n299 B.n226 10.6151
R2481 B.n299 B.n298 10.6151
R2482 B.n298 B.n297 10.6151
R2483 B.n297 B.n228 10.6151
R2484 B.n293 B.n228 10.6151
R2485 B.n293 B.n292 10.6151
R2486 B.n292 B.n291 10.6151
R2487 B.n291 B.n230 10.6151
R2488 B.n287 B.n230 10.6151
R2489 B.n287 B.n286 10.6151
R2490 B.n286 B.n285 10.6151
R2491 B.n285 B.n232 10.6151
R2492 B.n281 B.n232 10.6151
R2493 B.n281 B.n280 10.6151
R2494 B.n280 B.n279 10.6151
R2495 B.n279 B.n234 10.6151
R2496 B.n275 B.n234 10.6151
R2497 B.n275 B.n274 10.6151
R2498 B.n274 B.n273 10.6151
R2499 B.n273 B.n236 10.6151
R2500 B.n269 B.n236 10.6151
R2501 B.n269 B.n268 10.6151
R2502 B.n268 B.n267 10.6151
R2503 B.n267 B.n238 10.6151
R2504 B.n263 B.n238 10.6151
R2505 B.n263 B.n262 10.6151
R2506 B.n262 B.n261 10.6151
R2507 B.n261 B.n240 10.6151
R2508 B.n257 B.n240 10.6151
R2509 B.n257 B.n256 10.6151
R2510 B.n256 B.n255 10.6151
R2511 B.n255 B.n242 10.6151
R2512 B.n251 B.n242 10.6151
R2513 B.n251 B.n250 10.6151
R2514 B.n250 B.n249 10.6151
R2515 B.n249 B.n244 10.6151
R2516 B.n245 B.n244 10.6151
R2517 B.n245 B.n0 10.6151
R2518 B.n947 B.n1 10.6151
R2519 B.n947 B.n946 10.6151
R2520 B.n946 B.n945 10.6151
R2521 B.n945 B.n4 10.6151
R2522 B.n941 B.n4 10.6151
R2523 B.n941 B.n940 10.6151
R2524 B.n940 B.n939 10.6151
R2525 B.n939 B.n6 10.6151
R2526 B.n935 B.n6 10.6151
R2527 B.n935 B.n934 10.6151
R2528 B.n934 B.n933 10.6151
R2529 B.n933 B.n8 10.6151
R2530 B.n929 B.n8 10.6151
R2531 B.n929 B.n928 10.6151
R2532 B.n928 B.n927 10.6151
R2533 B.n927 B.n10 10.6151
R2534 B.n923 B.n10 10.6151
R2535 B.n923 B.n922 10.6151
R2536 B.n922 B.n921 10.6151
R2537 B.n921 B.n12 10.6151
R2538 B.n917 B.n12 10.6151
R2539 B.n917 B.n916 10.6151
R2540 B.n916 B.n915 10.6151
R2541 B.n915 B.n14 10.6151
R2542 B.n911 B.n14 10.6151
R2543 B.n911 B.n910 10.6151
R2544 B.n910 B.n909 10.6151
R2545 B.n909 B.n16 10.6151
R2546 B.n905 B.n16 10.6151
R2547 B.n905 B.n904 10.6151
R2548 B.n904 B.n903 10.6151
R2549 B.n903 B.n18 10.6151
R2550 B.n899 B.n18 10.6151
R2551 B.n899 B.n898 10.6151
R2552 B.n898 B.n897 10.6151
R2553 B.n897 B.n20 10.6151
R2554 B.n893 B.n20 10.6151
R2555 B.n893 B.n892 10.6151
R2556 B.n892 B.n891 10.6151
R2557 B.n891 B.n22 10.6151
R2558 B.n887 B.n22 10.6151
R2559 B.n887 B.n886 10.6151
R2560 B.n886 B.n885 10.6151
R2561 B.n885 B.n24 10.6151
R2562 B.n881 B.n24 10.6151
R2563 B.n881 B.n880 10.6151
R2564 B.n880 B.n879 10.6151
R2565 B.n879 B.n26 10.6151
R2566 B.n875 B.n26 10.6151
R2567 B.n875 B.n874 10.6151
R2568 B.n874 B.n873 10.6151
R2569 B.n873 B.n28 10.6151
R2570 B.n869 B.n28 10.6151
R2571 B.n869 B.n868 10.6151
R2572 B.n868 B.n867 10.6151
R2573 B.n867 B.n30 10.6151
R2574 B.n863 B.n30 10.6151
R2575 B.n863 B.n862 10.6151
R2576 B.n862 B.n861 10.6151
R2577 B.n861 B.n32 10.6151
R2578 B.n857 B.n32 10.6151
R2579 B.n857 B.n856 10.6151
R2580 B.n783 B.n60 9.36635
R2581 B.n766 B.n765 9.36635
R2582 B.n412 B.n411 9.36635
R2583 B.n429 B.n182 9.36635
R2584 B.n951 B.n0 2.81026
R2585 B.n951 B.n1 2.81026
R2586 B.n780 B.n60 1.24928
R2587 B.n767 B.n766 1.24928
R2588 B.n413 B.n412 1.24928
R2589 B.n426 B.n182 1.24928
R2590 VN.n68 VN.n67 161.3
R2591 VN.n66 VN.n36 161.3
R2592 VN.n65 VN.n64 161.3
R2593 VN.n63 VN.n37 161.3
R2594 VN.n62 VN.n61 161.3
R2595 VN.n60 VN.n38 161.3
R2596 VN.n59 VN.n58 161.3
R2597 VN.n57 VN.n56 161.3
R2598 VN.n55 VN.n40 161.3
R2599 VN.n54 VN.n53 161.3
R2600 VN.n52 VN.n41 161.3
R2601 VN.n51 VN.n50 161.3
R2602 VN.n49 VN.n42 161.3
R2603 VN.n48 VN.n47 161.3
R2604 VN.n46 VN.n43 161.3
R2605 VN.n33 VN.n32 161.3
R2606 VN.n31 VN.n1 161.3
R2607 VN.n30 VN.n29 161.3
R2608 VN.n28 VN.n2 161.3
R2609 VN.n27 VN.n26 161.3
R2610 VN.n25 VN.n3 161.3
R2611 VN.n24 VN.n23 161.3
R2612 VN.n22 VN.n21 161.3
R2613 VN.n20 VN.n5 161.3
R2614 VN.n19 VN.n18 161.3
R2615 VN.n17 VN.n6 161.3
R2616 VN.n16 VN.n15 161.3
R2617 VN.n14 VN.n7 161.3
R2618 VN.n13 VN.n12 161.3
R2619 VN.n11 VN.n8 161.3
R2620 VN.n45 VN.t4 136.927
R2621 VN.n10 VN.t0 136.927
R2622 VN.n9 VN.t6 103.844
R2623 VN.n4 VN.t2 103.844
R2624 VN.n0 VN.t7 103.844
R2625 VN.n44 VN.t3 103.844
R2626 VN.n39 VN.t5 103.844
R2627 VN.n35 VN.t1 103.844
R2628 VN.n34 VN.n0 73.1852
R2629 VN.n69 VN.n35 73.1852
R2630 VN.n10 VN.n9 68.9426
R2631 VN.n45 VN.n44 68.9426
R2632 VN VN.n69 56.9829
R2633 VN.n15 VN.n6 56.5193
R2634 VN.n50 VN.n41 56.5193
R2635 VN.n26 VN.n2 42.4359
R2636 VN.n61 VN.n37 42.4359
R2637 VN.n30 VN.n2 38.5509
R2638 VN.n65 VN.n37 38.5509
R2639 VN.n13 VN.n8 24.4675
R2640 VN.n14 VN.n13 24.4675
R2641 VN.n15 VN.n14 24.4675
R2642 VN.n19 VN.n6 24.4675
R2643 VN.n20 VN.n19 24.4675
R2644 VN.n21 VN.n20 24.4675
R2645 VN.n25 VN.n24 24.4675
R2646 VN.n26 VN.n25 24.4675
R2647 VN.n31 VN.n30 24.4675
R2648 VN.n32 VN.n31 24.4675
R2649 VN.n50 VN.n49 24.4675
R2650 VN.n49 VN.n48 24.4675
R2651 VN.n48 VN.n43 24.4675
R2652 VN.n61 VN.n60 24.4675
R2653 VN.n60 VN.n59 24.4675
R2654 VN.n56 VN.n55 24.4675
R2655 VN.n55 VN.n54 24.4675
R2656 VN.n54 VN.n41 24.4675
R2657 VN.n67 VN.n66 24.4675
R2658 VN.n66 VN.n65 24.4675
R2659 VN.n24 VN.n4 18.8401
R2660 VN.n59 VN.n39 18.8401
R2661 VN.n32 VN.n0 16.8827
R2662 VN.n67 VN.n35 16.8827
R2663 VN.n9 VN.n8 5.62791
R2664 VN.n21 VN.n4 5.62791
R2665 VN.n44 VN.n43 5.62791
R2666 VN.n56 VN.n39 5.62791
R2667 VN.n11 VN.n10 4.0558
R2668 VN.n46 VN.n45 4.05579
R2669 VN.n69 VN.n68 0.354971
R2670 VN.n34 VN.n33 0.354971
R2671 VN VN.n34 0.26696
R2672 VN.n68 VN.n36 0.189894
R2673 VN.n64 VN.n36 0.189894
R2674 VN.n64 VN.n63 0.189894
R2675 VN.n63 VN.n62 0.189894
R2676 VN.n62 VN.n38 0.189894
R2677 VN.n58 VN.n38 0.189894
R2678 VN.n58 VN.n57 0.189894
R2679 VN.n57 VN.n40 0.189894
R2680 VN.n53 VN.n40 0.189894
R2681 VN.n53 VN.n52 0.189894
R2682 VN.n52 VN.n51 0.189894
R2683 VN.n51 VN.n42 0.189894
R2684 VN.n47 VN.n42 0.189894
R2685 VN.n47 VN.n46 0.189894
R2686 VN.n12 VN.n11 0.189894
R2687 VN.n12 VN.n7 0.189894
R2688 VN.n16 VN.n7 0.189894
R2689 VN.n17 VN.n16 0.189894
R2690 VN.n18 VN.n17 0.189894
R2691 VN.n18 VN.n5 0.189894
R2692 VN.n22 VN.n5 0.189894
R2693 VN.n23 VN.n22 0.189894
R2694 VN.n23 VN.n3 0.189894
R2695 VN.n27 VN.n3 0.189894
R2696 VN.n28 VN.n27 0.189894
R2697 VN.n29 VN.n28 0.189894
R2698 VN.n29 VN.n1 0.189894
R2699 VN.n33 VN.n1 0.189894
R2700 VDD2.n2 VDD2.n1 72.5127
R2701 VDD2.n2 VDD2.n0 72.5127
R2702 VDD2 VDD2.n5 72.5099
R2703 VDD2.n4 VDD2.n3 70.9605
R2704 VDD2.n4 VDD2.n2 50.8144
R2705 VDD2.n5 VDD2.t4 2.21927
R2706 VDD2.n5 VDD2.t3 2.21927
R2707 VDD2.n3 VDD2.t6 2.21927
R2708 VDD2.n3 VDD2.t2 2.21927
R2709 VDD2.n1 VDD2.t5 2.21927
R2710 VDD2.n1 VDD2.t0 2.21927
R2711 VDD2.n0 VDD2.t7 2.21927
R2712 VDD2.n0 VDD2.t1 2.21927
R2713 VDD2 VDD2.n4 1.66645
C0 VP B 2.47362f
C1 VTAIL VDD1 9.151f
C2 VP VN 9.12969f
C3 VP VDD2 0.604402f
C4 VDD1 w_n4700_n3898# 2.27708f
C5 VTAIL B 6.22558f
C6 VN VTAIL 11.5553f
C7 VTAIL VDD2 9.21078f
C8 w_n4700_n3898# B 12.0829f
C9 VN w_n4700_n3898# 9.833691f
C10 VDD1 B 1.9648f
C11 VDD2 w_n4700_n3898# 2.42535f
C12 VN VDD1 0.152777f
C13 VDD1 VDD2 2.1888f
C14 VP VTAIL 11.5694f
C15 VP w_n4700_n3898# 10.446199f
C16 VP VDD1 11.476f
C17 VN B 1.44257f
C18 VDD2 B 2.086f
C19 VN VDD2 11.0262f
C20 VTAIL w_n4700_n3898# 4.86745f
C21 VDD2 VSUBS 2.406486f
C22 VDD1 VSUBS 3.09197f
C23 VTAIL VSUBS 1.593666f
C24 VN VSUBS 7.89006f
C25 VP VSUBS 4.508628f
C26 B VSUBS 6.119827f
C27 w_n4700_n3898# VSUBS 0.224754p
C28 VDD2.t7 VSUBS 0.370973f
C29 VDD2.t1 VSUBS 0.370973f
C30 VDD2.n0 VSUBS 3.02424f
C31 VDD2.t5 VSUBS 0.370973f
C32 VDD2.t0 VSUBS 0.370973f
C33 VDD2.n1 VSUBS 3.02424f
C34 VDD2.n2 VSUBS 5.69353f
C35 VDD2.t6 VSUBS 0.370973f
C36 VDD2.t2 VSUBS 0.370973f
C37 VDD2.n3 VSUBS 3.00034f
C38 VDD2.n4 VSUBS 4.74153f
C39 VDD2.t4 VSUBS 0.370973f
C40 VDD2.t3 VSUBS 0.370973f
C41 VDD2.n5 VSUBS 3.02418f
C42 VN.t7 VSUBS 3.22797f
C43 VN.n0 VSUBS 1.22199f
C44 VN.n1 VSUBS 0.023663f
C45 VN.n2 VSUBS 0.019251f
C46 VN.n3 VSUBS 0.023663f
C47 VN.t2 VSUBS 3.22797f
C48 VN.n4 VSUBS 1.12281f
C49 VN.n5 VSUBS 0.023663f
C50 VN.n6 VSUBS 0.034543f
C51 VN.n7 VSUBS 0.023663f
C52 VN.n8 VSUBS 0.027335f
C53 VN.t6 VSUBS 3.22797f
C54 VN.n9 VSUBS 1.19774f
C55 VN.t0 VSUBS 3.54139f
C56 VN.n10 VSUBS 1.14423f
C57 VN.n11 VSUBS 0.279934f
C58 VN.n12 VSUBS 0.023663f
C59 VN.n13 VSUBS 0.044102f
C60 VN.n14 VSUBS 0.044102f
C61 VN.n15 VSUBS 0.034543f
C62 VN.n16 VSUBS 0.023663f
C63 VN.n17 VSUBS 0.023663f
C64 VN.n18 VSUBS 0.023663f
C65 VN.n19 VSUBS 0.044102f
C66 VN.n20 VSUBS 0.044102f
C67 VN.n21 VSUBS 0.027335f
C68 VN.n22 VSUBS 0.023663f
C69 VN.n23 VSUBS 0.023663f
C70 VN.n24 VSUBS 0.039093f
C71 VN.n25 VSUBS 0.044102f
C72 VN.n26 VSUBS 0.046497f
C73 VN.n27 VSUBS 0.023663f
C74 VN.n28 VSUBS 0.023663f
C75 VN.n29 VSUBS 0.023663f
C76 VN.n30 VSUBS 0.047441f
C77 VN.n31 VSUBS 0.044102f
C78 VN.n32 VSUBS 0.037351f
C79 VN.n33 VSUBS 0.038191f
C80 VN.n34 VSUBS 0.055955f
C81 VN.t1 VSUBS 3.22797f
C82 VN.n35 VSUBS 1.22199f
C83 VN.n36 VSUBS 0.023663f
C84 VN.n37 VSUBS 0.019251f
C85 VN.n38 VSUBS 0.023663f
C86 VN.t5 VSUBS 3.22797f
C87 VN.n39 VSUBS 1.12281f
C88 VN.n40 VSUBS 0.023663f
C89 VN.n41 VSUBS 0.034543f
C90 VN.n42 VSUBS 0.023663f
C91 VN.n43 VSUBS 0.027335f
C92 VN.t4 VSUBS 3.54139f
C93 VN.t3 VSUBS 3.22797f
C94 VN.n44 VSUBS 1.19774f
C95 VN.n45 VSUBS 1.14423f
C96 VN.n46 VSUBS 0.279934f
C97 VN.n47 VSUBS 0.023663f
C98 VN.n48 VSUBS 0.044102f
C99 VN.n49 VSUBS 0.044102f
C100 VN.n50 VSUBS 0.034543f
C101 VN.n51 VSUBS 0.023663f
C102 VN.n52 VSUBS 0.023663f
C103 VN.n53 VSUBS 0.023663f
C104 VN.n54 VSUBS 0.044102f
C105 VN.n55 VSUBS 0.044102f
C106 VN.n56 VSUBS 0.027335f
C107 VN.n57 VSUBS 0.023663f
C108 VN.n58 VSUBS 0.023663f
C109 VN.n59 VSUBS 0.039093f
C110 VN.n60 VSUBS 0.044102f
C111 VN.n61 VSUBS 0.046497f
C112 VN.n62 VSUBS 0.023663f
C113 VN.n63 VSUBS 0.023663f
C114 VN.n64 VSUBS 0.023663f
C115 VN.n65 VSUBS 0.047441f
C116 VN.n66 VSUBS 0.044102f
C117 VN.n67 VSUBS 0.037351f
C118 VN.n68 VSUBS 0.038191f
C119 VN.n69 VSUBS 1.61935f
C120 B.n0 VSUBS 0.004735f
C121 B.n1 VSUBS 0.004735f
C122 B.n2 VSUBS 0.007488f
C123 B.n3 VSUBS 0.007488f
C124 B.n4 VSUBS 0.007488f
C125 B.n5 VSUBS 0.007488f
C126 B.n6 VSUBS 0.007488f
C127 B.n7 VSUBS 0.007488f
C128 B.n8 VSUBS 0.007488f
C129 B.n9 VSUBS 0.007488f
C130 B.n10 VSUBS 0.007488f
C131 B.n11 VSUBS 0.007488f
C132 B.n12 VSUBS 0.007488f
C133 B.n13 VSUBS 0.007488f
C134 B.n14 VSUBS 0.007488f
C135 B.n15 VSUBS 0.007488f
C136 B.n16 VSUBS 0.007488f
C137 B.n17 VSUBS 0.007488f
C138 B.n18 VSUBS 0.007488f
C139 B.n19 VSUBS 0.007488f
C140 B.n20 VSUBS 0.007488f
C141 B.n21 VSUBS 0.007488f
C142 B.n22 VSUBS 0.007488f
C143 B.n23 VSUBS 0.007488f
C144 B.n24 VSUBS 0.007488f
C145 B.n25 VSUBS 0.007488f
C146 B.n26 VSUBS 0.007488f
C147 B.n27 VSUBS 0.007488f
C148 B.n28 VSUBS 0.007488f
C149 B.n29 VSUBS 0.007488f
C150 B.n30 VSUBS 0.007488f
C151 B.n31 VSUBS 0.007488f
C152 B.n32 VSUBS 0.007488f
C153 B.n33 VSUBS 0.017822f
C154 B.n34 VSUBS 0.007488f
C155 B.n35 VSUBS 0.007488f
C156 B.n36 VSUBS 0.007488f
C157 B.n37 VSUBS 0.007488f
C158 B.n38 VSUBS 0.007488f
C159 B.n39 VSUBS 0.007488f
C160 B.n40 VSUBS 0.007488f
C161 B.n41 VSUBS 0.007488f
C162 B.n42 VSUBS 0.007488f
C163 B.n43 VSUBS 0.007488f
C164 B.n44 VSUBS 0.007488f
C165 B.n45 VSUBS 0.007488f
C166 B.n46 VSUBS 0.007488f
C167 B.n47 VSUBS 0.007488f
C168 B.n48 VSUBS 0.007488f
C169 B.n49 VSUBS 0.007488f
C170 B.n50 VSUBS 0.007488f
C171 B.n51 VSUBS 0.007488f
C172 B.n52 VSUBS 0.007488f
C173 B.n53 VSUBS 0.007488f
C174 B.n54 VSUBS 0.007488f
C175 B.n55 VSUBS 0.007488f
C176 B.n56 VSUBS 0.007488f
C177 B.n57 VSUBS 0.007488f
C178 B.t5 VSUBS 0.290142f
C179 B.t4 VSUBS 0.333988f
C180 B.t3 VSUBS 2.44063f
C181 B.n58 VSUBS 0.530323f
C182 B.n59 VSUBS 0.311012f
C183 B.n60 VSUBS 0.017349f
C184 B.n61 VSUBS 0.007488f
C185 B.n62 VSUBS 0.007488f
C186 B.n63 VSUBS 0.007488f
C187 B.n64 VSUBS 0.007488f
C188 B.n65 VSUBS 0.007488f
C189 B.t8 VSUBS 0.290146f
C190 B.t7 VSUBS 0.333991f
C191 B.t6 VSUBS 2.44063f
C192 B.n66 VSUBS 0.53032f
C193 B.n67 VSUBS 0.311009f
C194 B.n68 VSUBS 0.007488f
C195 B.n69 VSUBS 0.007488f
C196 B.n70 VSUBS 0.007488f
C197 B.n71 VSUBS 0.007488f
C198 B.n72 VSUBS 0.007488f
C199 B.n73 VSUBS 0.007488f
C200 B.n74 VSUBS 0.007488f
C201 B.n75 VSUBS 0.007488f
C202 B.n76 VSUBS 0.007488f
C203 B.n77 VSUBS 0.007488f
C204 B.n78 VSUBS 0.007488f
C205 B.n79 VSUBS 0.007488f
C206 B.n80 VSUBS 0.007488f
C207 B.n81 VSUBS 0.007488f
C208 B.n82 VSUBS 0.007488f
C209 B.n83 VSUBS 0.007488f
C210 B.n84 VSUBS 0.007488f
C211 B.n85 VSUBS 0.007488f
C212 B.n86 VSUBS 0.007488f
C213 B.n87 VSUBS 0.007488f
C214 B.n88 VSUBS 0.007488f
C215 B.n89 VSUBS 0.007488f
C216 B.n90 VSUBS 0.007488f
C217 B.n91 VSUBS 0.007488f
C218 B.n92 VSUBS 0.018667f
C219 B.n93 VSUBS 0.007488f
C220 B.n94 VSUBS 0.007488f
C221 B.n95 VSUBS 0.007488f
C222 B.n96 VSUBS 0.007488f
C223 B.n97 VSUBS 0.007488f
C224 B.n98 VSUBS 0.007488f
C225 B.n99 VSUBS 0.007488f
C226 B.n100 VSUBS 0.007488f
C227 B.n101 VSUBS 0.007488f
C228 B.n102 VSUBS 0.007488f
C229 B.n103 VSUBS 0.007488f
C230 B.n104 VSUBS 0.007488f
C231 B.n105 VSUBS 0.007488f
C232 B.n106 VSUBS 0.007488f
C233 B.n107 VSUBS 0.007488f
C234 B.n108 VSUBS 0.007488f
C235 B.n109 VSUBS 0.007488f
C236 B.n110 VSUBS 0.007488f
C237 B.n111 VSUBS 0.007488f
C238 B.n112 VSUBS 0.007488f
C239 B.n113 VSUBS 0.007488f
C240 B.n114 VSUBS 0.007488f
C241 B.n115 VSUBS 0.007488f
C242 B.n116 VSUBS 0.007488f
C243 B.n117 VSUBS 0.007488f
C244 B.n118 VSUBS 0.007488f
C245 B.n119 VSUBS 0.007488f
C246 B.n120 VSUBS 0.007488f
C247 B.n121 VSUBS 0.007488f
C248 B.n122 VSUBS 0.007488f
C249 B.n123 VSUBS 0.007488f
C250 B.n124 VSUBS 0.007488f
C251 B.n125 VSUBS 0.007488f
C252 B.n126 VSUBS 0.007488f
C253 B.n127 VSUBS 0.007488f
C254 B.n128 VSUBS 0.007488f
C255 B.n129 VSUBS 0.007488f
C256 B.n130 VSUBS 0.007488f
C257 B.n131 VSUBS 0.007488f
C258 B.n132 VSUBS 0.007488f
C259 B.n133 VSUBS 0.007488f
C260 B.n134 VSUBS 0.007488f
C261 B.n135 VSUBS 0.007488f
C262 B.n136 VSUBS 0.007488f
C263 B.n137 VSUBS 0.007488f
C264 B.n138 VSUBS 0.007488f
C265 B.n139 VSUBS 0.007488f
C266 B.n140 VSUBS 0.007488f
C267 B.n141 VSUBS 0.007488f
C268 B.n142 VSUBS 0.007488f
C269 B.n143 VSUBS 0.007488f
C270 B.n144 VSUBS 0.007488f
C271 B.n145 VSUBS 0.007488f
C272 B.n146 VSUBS 0.007488f
C273 B.n147 VSUBS 0.007488f
C274 B.n148 VSUBS 0.007488f
C275 B.n149 VSUBS 0.007488f
C276 B.n150 VSUBS 0.007488f
C277 B.n151 VSUBS 0.007488f
C278 B.n152 VSUBS 0.007488f
C279 B.n153 VSUBS 0.007488f
C280 B.n154 VSUBS 0.007488f
C281 B.n155 VSUBS 0.017822f
C282 B.n156 VSUBS 0.007488f
C283 B.n157 VSUBS 0.007488f
C284 B.n158 VSUBS 0.007488f
C285 B.n159 VSUBS 0.007488f
C286 B.n160 VSUBS 0.007488f
C287 B.n161 VSUBS 0.007488f
C288 B.n162 VSUBS 0.007488f
C289 B.n163 VSUBS 0.007488f
C290 B.n164 VSUBS 0.007488f
C291 B.n165 VSUBS 0.007488f
C292 B.n166 VSUBS 0.007488f
C293 B.n167 VSUBS 0.007488f
C294 B.n168 VSUBS 0.007488f
C295 B.n169 VSUBS 0.007488f
C296 B.n170 VSUBS 0.007488f
C297 B.n171 VSUBS 0.007488f
C298 B.n172 VSUBS 0.007488f
C299 B.n173 VSUBS 0.007488f
C300 B.n174 VSUBS 0.007488f
C301 B.n175 VSUBS 0.007488f
C302 B.n176 VSUBS 0.007488f
C303 B.n177 VSUBS 0.007488f
C304 B.n178 VSUBS 0.007488f
C305 B.n179 VSUBS 0.007488f
C306 B.t10 VSUBS 0.290146f
C307 B.t11 VSUBS 0.333991f
C308 B.t9 VSUBS 2.44063f
C309 B.n180 VSUBS 0.53032f
C310 B.n181 VSUBS 0.311009f
C311 B.n182 VSUBS 0.017349f
C312 B.n183 VSUBS 0.007488f
C313 B.n184 VSUBS 0.007488f
C314 B.n185 VSUBS 0.007488f
C315 B.n186 VSUBS 0.007488f
C316 B.n187 VSUBS 0.007488f
C317 B.t1 VSUBS 0.290142f
C318 B.t2 VSUBS 0.333988f
C319 B.t0 VSUBS 2.44063f
C320 B.n188 VSUBS 0.530323f
C321 B.n189 VSUBS 0.311012f
C322 B.n190 VSUBS 0.007488f
C323 B.n191 VSUBS 0.007488f
C324 B.n192 VSUBS 0.007488f
C325 B.n193 VSUBS 0.007488f
C326 B.n194 VSUBS 0.007488f
C327 B.n195 VSUBS 0.007488f
C328 B.n196 VSUBS 0.007488f
C329 B.n197 VSUBS 0.007488f
C330 B.n198 VSUBS 0.007488f
C331 B.n199 VSUBS 0.007488f
C332 B.n200 VSUBS 0.007488f
C333 B.n201 VSUBS 0.007488f
C334 B.n202 VSUBS 0.007488f
C335 B.n203 VSUBS 0.007488f
C336 B.n204 VSUBS 0.007488f
C337 B.n205 VSUBS 0.007488f
C338 B.n206 VSUBS 0.007488f
C339 B.n207 VSUBS 0.007488f
C340 B.n208 VSUBS 0.007488f
C341 B.n209 VSUBS 0.007488f
C342 B.n210 VSUBS 0.007488f
C343 B.n211 VSUBS 0.007488f
C344 B.n212 VSUBS 0.007488f
C345 B.n213 VSUBS 0.007488f
C346 B.n214 VSUBS 0.017822f
C347 B.n215 VSUBS 0.007488f
C348 B.n216 VSUBS 0.007488f
C349 B.n217 VSUBS 0.007488f
C350 B.n218 VSUBS 0.007488f
C351 B.n219 VSUBS 0.007488f
C352 B.n220 VSUBS 0.007488f
C353 B.n221 VSUBS 0.007488f
C354 B.n222 VSUBS 0.007488f
C355 B.n223 VSUBS 0.007488f
C356 B.n224 VSUBS 0.007488f
C357 B.n225 VSUBS 0.007488f
C358 B.n226 VSUBS 0.007488f
C359 B.n227 VSUBS 0.007488f
C360 B.n228 VSUBS 0.007488f
C361 B.n229 VSUBS 0.007488f
C362 B.n230 VSUBS 0.007488f
C363 B.n231 VSUBS 0.007488f
C364 B.n232 VSUBS 0.007488f
C365 B.n233 VSUBS 0.007488f
C366 B.n234 VSUBS 0.007488f
C367 B.n235 VSUBS 0.007488f
C368 B.n236 VSUBS 0.007488f
C369 B.n237 VSUBS 0.007488f
C370 B.n238 VSUBS 0.007488f
C371 B.n239 VSUBS 0.007488f
C372 B.n240 VSUBS 0.007488f
C373 B.n241 VSUBS 0.007488f
C374 B.n242 VSUBS 0.007488f
C375 B.n243 VSUBS 0.007488f
C376 B.n244 VSUBS 0.007488f
C377 B.n245 VSUBS 0.007488f
C378 B.n246 VSUBS 0.007488f
C379 B.n247 VSUBS 0.007488f
C380 B.n248 VSUBS 0.007488f
C381 B.n249 VSUBS 0.007488f
C382 B.n250 VSUBS 0.007488f
C383 B.n251 VSUBS 0.007488f
C384 B.n252 VSUBS 0.007488f
C385 B.n253 VSUBS 0.007488f
C386 B.n254 VSUBS 0.007488f
C387 B.n255 VSUBS 0.007488f
C388 B.n256 VSUBS 0.007488f
C389 B.n257 VSUBS 0.007488f
C390 B.n258 VSUBS 0.007488f
C391 B.n259 VSUBS 0.007488f
C392 B.n260 VSUBS 0.007488f
C393 B.n261 VSUBS 0.007488f
C394 B.n262 VSUBS 0.007488f
C395 B.n263 VSUBS 0.007488f
C396 B.n264 VSUBS 0.007488f
C397 B.n265 VSUBS 0.007488f
C398 B.n266 VSUBS 0.007488f
C399 B.n267 VSUBS 0.007488f
C400 B.n268 VSUBS 0.007488f
C401 B.n269 VSUBS 0.007488f
C402 B.n270 VSUBS 0.007488f
C403 B.n271 VSUBS 0.007488f
C404 B.n272 VSUBS 0.007488f
C405 B.n273 VSUBS 0.007488f
C406 B.n274 VSUBS 0.007488f
C407 B.n275 VSUBS 0.007488f
C408 B.n276 VSUBS 0.007488f
C409 B.n277 VSUBS 0.007488f
C410 B.n278 VSUBS 0.007488f
C411 B.n279 VSUBS 0.007488f
C412 B.n280 VSUBS 0.007488f
C413 B.n281 VSUBS 0.007488f
C414 B.n282 VSUBS 0.007488f
C415 B.n283 VSUBS 0.007488f
C416 B.n284 VSUBS 0.007488f
C417 B.n285 VSUBS 0.007488f
C418 B.n286 VSUBS 0.007488f
C419 B.n287 VSUBS 0.007488f
C420 B.n288 VSUBS 0.007488f
C421 B.n289 VSUBS 0.007488f
C422 B.n290 VSUBS 0.007488f
C423 B.n291 VSUBS 0.007488f
C424 B.n292 VSUBS 0.007488f
C425 B.n293 VSUBS 0.007488f
C426 B.n294 VSUBS 0.007488f
C427 B.n295 VSUBS 0.007488f
C428 B.n296 VSUBS 0.007488f
C429 B.n297 VSUBS 0.007488f
C430 B.n298 VSUBS 0.007488f
C431 B.n299 VSUBS 0.007488f
C432 B.n300 VSUBS 0.007488f
C433 B.n301 VSUBS 0.007488f
C434 B.n302 VSUBS 0.007488f
C435 B.n303 VSUBS 0.007488f
C436 B.n304 VSUBS 0.007488f
C437 B.n305 VSUBS 0.007488f
C438 B.n306 VSUBS 0.007488f
C439 B.n307 VSUBS 0.007488f
C440 B.n308 VSUBS 0.007488f
C441 B.n309 VSUBS 0.007488f
C442 B.n310 VSUBS 0.007488f
C443 B.n311 VSUBS 0.007488f
C444 B.n312 VSUBS 0.007488f
C445 B.n313 VSUBS 0.007488f
C446 B.n314 VSUBS 0.007488f
C447 B.n315 VSUBS 0.007488f
C448 B.n316 VSUBS 0.007488f
C449 B.n317 VSUBS 0.007488f
C450 B.n318 VSUBS 0.007488f
C451 B.n319 VSUBS 0.007488f
C452 B.n320 VSUBS 0.007488f
C453 B.n321 VSUBS 0.007488f
C454 B.n322 VSUBS 0.007488f
C455 B.n323 VSUBS 0.007488f
C456 B.n324 VSUBS 0.007488f
C457 B.n325 VSUBS 0.007488f
C458 B.n326 VSUBS 0.007488f
C459 B.n327 VSUBS 0.007488f
C460 B.n328 VSUBS 0.007488f
C461 B.n329 VSUBS 0.007488f
C462 B.n330 VSUBS 0.007488f
C463 B.n331 VSUBS 0.007488f
C464 B.n332 VSUBS 0.007488f
C465 B.n333 VSUBS 0.007488f
C466 B.n334 VSUBS 0.007488f
C467 B.n335 VSUBS 0.007488f
C468 B.n336 VSUBS 0.007488f
C469 B.n337 VSUBS 0.017822f
C470 B.n338 VSUBS 0.018296f
C471 B.n339 VSUBS 0.018296f
C472 B.n340 VSUBS 0.007488f
C473 B.n341 VSUBS 0.007488f
C474 B.n342 VSUBS 0.007488f
C475 B.n343 VSUBS 0.007488f
C476 B.n344 VSUBS 0.007488f
C477 B.n345 VSUBS 0.007488f
C478 B.n346 VSUBS 0.007488f
C479 B.n347 VSUBS 0.007488f
C480 B.n348 VSUBS 0.007488f
C481 B.n349 VSUBS 0.007488f
C482 B.n350 VSUBS 0.007488f
C483 B.n351 VSUBS 0.007488f
C484 B.n352 VSUBS 0.007488f
C485 B.n353 VSUBS 0.007488f
C486 B.n354 VSUBS 0.007488f
C487 B.n355 VSUBS 0.007488f
C488 B.n356 VSUBS 0.007488f
C489 B.n357 VSUBS 0.007488f
C490 B.n358 VSUBS 0.007488f
C491 B.n359 VSUBS 0.007488f
C492 B.n360 VSUBS 0.007488f
C493 B.n361 VSUBS 0.007488f
C494 B.n362 VSUBS 0.007488f
C495 B.n363 VSUBS 0.007488f
C496 B.n364 VSUBS 0.007488f
C497 B.n365 VSUBS 0.007488f
C498 B.n366 VSUBS 0.007488f
C499 B.n367 VSUBS 0.007488f
C500 B.n368 VSUBS 0.007488f
C501 B.n369 VSUBS 0.007488f
C502 B.n370 VSUBS 0.007488f
C503 B.n371 VSUBS 0.007488f
C504 B.n372 VSUBS 0.007488f
C505 B.n373 VSUBS 0.007488f
C506 B.n374 VSUBS 0.007488f
C507 B.n375 VSUBS 0.007488f
C508 B.n376 VSUBS 0.007488f
C509 B.n377 VSUBS 0.007488f
C510 B.n378 VSUBS 0.007488f
C511 B.n379 VSUBS 0.007488f
C512 B.n380 VSUBS 0.007488f
C513 B.n381 VSUBS 0.007488f
C514 B.n382 VSUBS 0.007488f
C515 B.n383 VSUBS 0.007488f
C516 B.n384 VSUBS 0.007488f
C517 B.n385 VSUBS 0.007488f
C518 B.n386 VSUBS 0.007488f
C519 B.n387 VSUBS 0.007488f
C520 B.n388 VSUBS 0.007488f
C521 B.n389 VSUBS 0.007488f
C522 B.n390 VSUBS 0.007488f
C523 B.n391 VSUBS 0.007488f
C524 B.n392 VSUBS 0.007488f
C525 B.n393 VSUBS 0.007488f
C526 B.n394 VSUBS 0.007488f
C527 B.n395 VSUBS 0.007488f
C528 B.n396 VSUBS 0.007488f
C529 B.n397 VSUBS 0.007488f
C530 B.n398 VSUBS 0.007488f
C531 B.n399 VSUBS 0.007488f
C532 B.n400 VSUBS 0.007488f
C533 B.n401 VSUBS 0.007488f
C534 B.n402 VSUBS 0.007488f
C535 B.n403 VSUBS 0.007488f
C536 B.n404 VSUBS 0.007488f
C537 B.n405 VSUBS 0.007488f
C538 B.n406 VSUBS 0.007488f
C539 B.n407 VSUBS 0.007488f
C540 B.n408 VSUBS 0.007488f
C541 B.n409 VSUBS 0.007488f
C542 B.n410 VSUBS 0.007488f
C543 B.n411 VSUBS 0.007047f
C544 B.n412 VSUBS 0.017349f
C545 B.n413 VSUBS 0.004184f
C546 B.n414 VSUBS 0.007488f
C547 B.n415 VSUBS 0.007488f
C548 B.n416 VSUBS 0.007488f
C549 B.n417 VSUBS 0.007488f
C550 B.n418 VSUBS 0.007488f
C551 B.n419 VSUBS 0.007488f
C552 B.n420 VSUBS 0.007488f
C553 B.n421 VSUBS 0.007488f
C554 B.n422 VSUBS 0.007488f
C555 B.n423 VSUBS 0.007488f
C556 B.n424 VSUBS 0.007488f
C557 B.n425 VSUBS 0.007488f
C558 B.n426 VSUBS 0.004184f
C559 B.n427 VSUBS 0.007488f
C560 B.n428 VSUBS 0.007488f
C561 B.n429 VSUBS 0.007047f
C562 B.n430 VSUBS 0.007488f
C563 B.n431 VSUBS 0.007488f
C564 B.n432 VSUBS 0.007488f
C565 B.n433 VSUBS 0.007488f
C566 B.n434 VSUBS 0.007488f
C567 B.n435 VSUBS 0.007488f
C568 B.n436 VSUBS 0.007488f
C569 B.n437 VSUBS 0.007488f
C570 B.n438 VSUBS 0.007488f
C571 B.n439 VSUBS 0.007488f
C572 B.n440 VSUBS 0.007488f
C573 B.n441 VSUBS 0.007488f
C574 B.n442 VSUBS 0.007488f
C575 B.n443 VSUBS 0.007488f
C576 B.n444 VSUBS 0.007488f
C577 B.n445 VSUBS 0.007488f
C578 B.n446 VSUBS 0.007488f
C579 B.n447 VSUBS 0.007488f
C580 B.n448 VSUBS 0.007488f
C581 B.n449 VSUBS 0.007488f
C582 B.n450 VSUBS 0.007488f
C583 B.n451 VSUBS 0.007488f
C584 B.n452 VSUBS 0.007488f
C585 B.n453 VSUBS 0.007488f
C586 B.n454 VSUBS 0.007488f
C587 B.n455 VSUBS 0.007488f
C588 B.n456 VSUBS 0.007488f
C589 B.n457 VSUBS 0.007488f
C590 B.n458 VSUBS 0.007488f
C591 B.n459 VSUBS 0.007488f
C592 B.n460 VSUBS 0.007488f
C593 B.n461 VSUBS 0.007488f
C594 B.n462 VSUBS 0.007488f
C595 B.n463 VSUBS 0.007488f
C596 B.n464 VSUBS 0.007488f
C597 B.n465 VSUBS 0.007488f
C598 B.n466 VSUBS 0.007488f
C599 B.n467 VSUBS 0.007488f
C600 B.n468 VSUBS 0.007488f
C601 B.n469 VSUBS 0.007488f
C602 B.n470 VSUBS 0.007488f
C603 B.n471 VSUBS 0.007488f
C604 B.n472 VSUBS 0.007488f
C605 B.n473 VSUBS 0.007488f
C606 B.n474 VSUBS 0.007488f
C607 B.n475 VSUBS 0.007488f
C608 B.n476 VSUBS 0.007488f
C609 B.n477 VSUBS 0.007488f
C610 B.n478 VSUBS 0.007488f
C611 B.n479 VSUBS 0.007488f
C612 B.n480 VSUBS 0.007488f
C613 B.n481 VSUBS 0.007488f
C614 B.n482 VSUBS 0.007488f
C615 B.n483 VSUBS 0.007488f
C616 B.n484 VSUBS 0.007488f
C617 B.n485 VSUBS 0.007488f
C618 B.n486 VSUBS 0.007488f
C619 B.n487 VSUBS 0.007488f
C620 B.n488 VSUBS 0.007488f
C621 B.n489 VSUBS 0.007488f
C622 B.n490 VSUBS 0.007488f
C623 B.n491 VSUBS 0.007488f
C624 B.n492 VSUBS 0.007488f
C625 B.n493 VSUBS 0.007488f
C626 B.n494 VSUBS 0.007488f
C627 B.n495 VSUBS 0.007488f
C628 B.n496 VSUBS 0.007488f
C629 B.n497 VSUBS 0.007488f
C630 B.n498 VSUBS 0.007488f
C631 B.n499 VSUBS 0.007488f
C632 B.n500 VSUBS 0.018296f
C633 B.n501 VSUBS 0.018296f
C634 B.n502 VSUBS 0.017822f
C635 B.n503 VSUBS 0.007488f
C636 B.n504 VSUBS 0.007488f
C637 B.n505 VSUBS 0.007488f
C638 B.n506 VSUBS 0.007488f
C639 B.n507 VSUBS 0.007488f
C640 B.n508 VSUBS 0.007488f
C641 B.n509 VSUBS 0.007488f
C642 B.n510 VSUBS 0.007488f
C643 B.n511 VSUBS 0.007488f
C644 B.n512 VSUBS 0.007488f
C645 B.n513 VSUBS 0.007488f
C646 B.n514 VSUBS 0.007488f
C647 B.n515 VSUBS 0.007488f
C648 B.n516 VSUBS 0.007488f
C649 B.n517 VSUBS 0.007488f
C650 B.n518 VSUBS 0.007488f
C651 B.n519 VSUBS 0.007488f
C652 B.n520 VSUBS 0.007488f
C653 B.n521 VSUBS 0.007488f
C654 B.n522 VSUBS 0.007488f
C655 B.n523 VSUBS 0.007488f
C656 B.n524 VSUBS 0.007488f
C657 B.n525 VSUBS 0.007488f
C658 B.n526 VSUBS 0.007488f
C659 B.n527 VSUBS 0.007488f
C660 B.n528 VSUBS 0.007488f
C661 B.n529 VSUBS 0.007488f
C662 B.n530 VSUBS 0.007488f
C663 B.n531 VSUBS 0.007488f
C664 B.n532 VSUBS 0.007488f
C665 B.n533 VSUBS 0.007488f
C666 B.n534 VSUBS 0.007488f
C667 B.n535 VSUBS 0.007488f
C668 B.n536 VSUBS 0.007488f
C669 B.n537 VSUBS 0.007488f
C670 B.n538 VSUBS 0.007488f
C671 B.n539 VSUBS 0.007488f
C672 B.n540 VSUBS 0.007488f
C673 B.n541 VSUBS 0.007488f
C674 B.n542 VSUBS 0.007488f
C675 B.n543 VSUBS 0.007488f
C676 B.n544 VSUBS 0.007488f
C677 B.n545 VSUBS 0.007488f
C678 B.n546 VSUBS 0.007488f
C679 B.n547 VSUBS 0.007488f
C680 B.n548 VSUBS 0.007488f
C681 B.n549 VSUBS 0.007488f
C682 B.n550 VSUBS 0.007488f
C683 B.n551 VSUBS 0.007488f
C684 B.n552 VSUBS 0.007488f
C685 B.n553 VSUBS 0.007488f
C686 B.n554 VSUBS 0.007488f
C687 B.n555 VSUBS 0.007488f
C688 B.n556 VSUBS 0.007488f
C689 B.n557 VSUBS 0.007488f
C690 B.n558 VSUBS 0.007488f
C691 B.n559 VSUBS 0.007488f
C692 B.n560 VSUBS 0.007488f
C693 B.n561 VSUBS 0.007488f
C694 B.n562 VSUBS 0.007488f
C695 B.n563 VSUBS 0.007488f
C696 B.n564 VSUBS 0.007488f
C697 B.n565 VSUBS 0.007488f
C698 B.n566 VSUBS 0.007488f
C699 B.n567 VSUBS 0.007488f
C700 B.n568 VSUBS 0.007488f
C701 B.n569 VSUBS 0.007488f
C702 B.n570 VSUBS 0.007488f
C703 B.n571 VSUBS 0.007488f
C704 B.n572 VSUBS 0.007488f
C705 B.n573 VSUBS 0.007488f
C706 B.n574 VSUBS 0.007488f
C707 B.n575 VSUBS 0.007488f
C708 B.n576 VSUBS 0.007488f
C709 B.n577 VSUBS 0.007488f
C710 B.n578 VSUBS 0.007488f
C711 B.n579 VSUBS 0.007488f
C712 B.n580 VSUBS 0.007488f
C713 B.n581 VSUBS 0.007488f
C714 B.n582 VSUBS 0.007488f
C715 B.n583 VSUBS 0.007488f
C716 B.n584 VSUBS 0.007488f
C717 B.n585 VSUBS 0.007488f
C718 B.n586 VSUBS 0.007488f
C719 B.n587 VSUBS 0.007488f
C720 B.n588 VSUBS 0.007488f
C721 B.n589 VSUBS 0.007488f
C722 B.n590 VSUBS 0.007488f
C723 B.n591 VSUBS 0.007488f
C724 B.n592 VSUBS 0.007488f
C725 B.n593 VSUBS 0.007488f
C726 B.n594 VSUBS 0.007488f
C727 B.n595 VSUBS 0.007488f
C728 B.n596 VSUBS 0.007488f
C729 B.n597 VSUBS 0.007488f
C730 B.n598 VSUBS 0.007488f
C731 B.n599 VSUBS 0.007488f
C732 B.n600 VSUBS 0.007488f
C733 B.n601 VSUBS 0.007488f
C734 B.n602 VSUBS 0.007488f
C735 B.n603 VSUBS 0.007488f
C736 B.n604 VSUBS 0.007488f
C737 B.n605 VSUBS 0.007488f
C738 B.n606 VSUBS 0.007488f
C739 B.n607 VSUBS 0.007488f
C740 B.n608 VSUBS 0.007488f
C741 B.n609 VSUBS 0.007488f
C742 B.n610 VSUBS 0.007488f
C743 B.n611 VSUBS 0.007488f
C744 B.n612 VSUBS 0.007488f
C745 B.n613 VSUBS 0.007488f
C746 B.n614 VSUBS 0.007488f
C747 B.n615 VSUBS 0.007488f
C748 B.n616 VSUBS 0.007488f
C749 B.n617 VSUBS 0.007488f
C750 B.n618 VSUBS 0.007488f
C751 B.n619 VSUBS 0.007488f
C752 B.n620 VSUBS 0.007488f
C753 B.n621 VSUBS 0.007488f
C754 B.n622 VSUBS 0.007488f
C755 B.n623 VSUBS 0.007488f
C756 B.n624 VSUBS 0.007488f
C757 B.n625 VSUBS 0.007488f
C758 B.n626 VSUBS 0.007488f
C759 B.n627 VSUBS 0.007488f
C760 B.n628 VSUBS 0.007488f
C761 B.n629 VSUBS 0.007488f
C762 B.n630 VSUBS 0.007488f
C763 B.n631 VSUBS 0.007488f
C764 B.n632 VSUBS 0.007488f
C765 B.n633 VSUBS 0.007488f
C766 B.n634 VSUBS 0.007488f
C767 B.n635 VSUBS 0.007488f
C768 B.n636 VSUBS 0.007488f
C769 B.n637 VSUBS 0.007488f
C770 B.n638 VSUBS 0.007488f
C771 B.n639 VSUBS 0.007488f
C772 B.n640 VSUBS 0.007488f
C773 B.n641 VSUBS 0.007488f
C774 B.n642 VSUBS 0.007488f
C775 B.n643 VSUBS 0.007488f
C776 B.n644 VSUBS 0.007488f
C777 B.n645 VSUBS 0.007488f
C778 B.n646 VSUBS 0.007488f
C779 B.n647 VSUBS 0.007488f
C780 B.n648 VSUBS 0.007488f
C781 B.n649 VSUBS 0.007488f
C782 B.n650 VSUBS 0.007488f
C783 B.n651 VSUBS 0.007488f
C784 B.n652 VSUBS 0.007488f
C785 B.n653 VSUBS 0.007488f
C786 B.n654 VSUBS 0.007488f
C787 B.n655 VSUBS 0.007488f
C788 B.n656 VSUBS 0.007488f
C789 B.n657 VSUBS 0.007488f
C790 B.n658 VSUBS 0.007488f
C791 B.n659 VSUBS 0.007488f
C792 B.n660 VSUBS 0.007488f
C793 B.n661 VSUBS 0.007488f
C794 B.n662 VSUBS 0.007488f
C795 B.n663 VSUBS 0.007488f
C796 B.n664 VSUBS 0.007488f
C797 B.n665 VSUBS 0.007488f
C798 B.n666 VSUBS 0.007488f
C799 B.n667 VSUBS 0.007488f
C800 B.n668 VSUBS 0.007488f
C801 B.n669 VSUBS 0.007488f
C802 B.n670 VSUBS 0.007488f
C803 B.n671 VSUBS 0.007488f
C804 B.n672 VSUBS 0.007488f
C805 B.n673 VSUBS 0.007488f
C806 B.n674 VSUBS 0.007488f
C807 B.n675 VSUBS 0.007488f
C808 B.n676 VSUBS 0.007488f
C809 B.n677 VSUBS 0.007488f
C810 B.n678 VSUBS 0.007488f
C811 B.n679 VSUBS 0.007488f
C812 B.n680 VSUBS 0.007488f
C813 B.n681 VSUBS 0.007488f
C814 B.n682 VSUBS 0.007488f
C815 B.n683 VSUBS 0.007488f
C816 B.n684 VSUBS 0.007488f
C817 B.n685 VSUBS 0.007488f
C818 B.n686 VSUBS 0.007488f
C819 B.n687 VSUBS 0.007488f
C820 B.n688 VSUBS 0.007488f
C821 B.n689 VSUBS 0.007488f
C822 B.n690 VSUBS 0.007488f
C823 B.n691 VSUBS 0.017822f
C824 B.n692 VSUBS 0.018296f
C825 B.n693 VSUBS 0.017451f
C826 B.n694 VSUBS 0.007488f
C827 B.n695 VSUBS 0.007488f
C828 B.n696 VSUBS 0.007488f
C829 B.n697 VSUBS 0.007488f
C830 B.n698 VSUBS 0.007488f
C831 B.n699 VSUBS 0.007488f
C832 B.n700 VSUBS 0.007488f
C833 B.n701 VSUBS 0.007488f
C834 B.n702 VSUBS 0.007488f
C835 B.n703 VSUBS 0.007488f
C836 B.n704 VSUBS 0.007488f
C837 B.n705 VSUBS 0.007488f
C838 B.n706 VSUBS 0.007488f
C839 B.n707 VSUBS 0.007488f
C840 B.n708 VSUBS 0.007488f
C841 B.n709 VSUBS 0.007488f
C842 B.n710 VSUBS 0.007488f
C843 B.n711 VSUBS 0.007488f
C844 B.n712 VSUBS 0.007488f
C845 B.n713 VSUBS 0.007488f
C846 B.n714 VSUBS 0.007488f
C847 B.n715 VSUBS 0.007488f
C848 B.n716 VSUBS 0.007488f
C849 B.n717 VSUBS 0.007488f
C850 B.n718 VSUBS 0.007488f
C851 B.n719 VSUBS 0.007488f
C852 B.n720 VSUBS 0.007488f
C853 B.n721 VSUBS 0.007488f
C854 B.n722 VSUBS 0.007488f
C855 B.n723 VSUBS 0.007488f
C856 B.n724 VSUBS 0.007488f
C857 B.n725 VSUBS 0.007488f
C858 B.n726 VSUBS 0.007488f
C859 B.n727 VSUBS 0.007488f
C860 B.n728 VSUBS 0.007488f
C861 B.n729 VSUBS 0.007488f
C862 B.n730 VSUBS 0.007488f
C863 B.n731 VSUBS 0.007488f
C864 B.n732 VSUBS 0.007488f
C865 B.n733 VSUBS 0.007488f
C866 B.n734 VSUBS 0.007488f
C867 B.n735 VSUBS 0.007488f
C868 B.n736 VSUBS 0.007488f
C869 B.n737 VSUBS 0.007488f
C870 B.n738 VSUBS 0.007488f
C871 B.n739 VSUBS 0.007488f
C872 B.n740 VSUBS 0.007488f
C873 B.n741 VSUBS 0.007488f
C874 B.n742 VSUBS 0.007488f
C875 B.n743 VSUBS 0.007488f
C876 B.n744 VSUBS 0.007488f
C877 B.n745 VSUBS 0.007488f
C878 B.n746 VSUBS 0.007488f
C879 B.n747 VSUBS 0.007488f
C880 B.n748 VSUBS 0.007488f
C881 B.n749 VSUBS 0.007488f
C882 B.n750 VSUBS 0.007488f
C883 B.n751 VSUBS 0.007488f
C884 B.n752 VSUBS 0.007488f
C885 B.n753 VSUBS 0.007488f
C886 B.n754 VSUBS 0.007488f
C887 B.n755 VSUBS 0.007488f
C888 B.n756 VSUBS 0.007488f
C889 B.n757 VSUBS 0.007488f
C890 B.n758 VSUBS 0.007488f
C891 B.n759 VSUBS 0.007488f
C892 B.n760 VSUBS 0.007488f
C893 B.n761 VSUBS 0.007488f
C894 B.n762 VSUBS 0.007488f
C895 B.n763 VSUBS 0.007488f
C896 B.n764 VSUBS 0.007488f
C897 B.n765 VSUBS 0.007047f
C898 B.n766 VSUBS 0.017349f
C899 B.n767 VSUBS 0.004184f
C900 B.n768 VSUBS 0.007488f
C901 B.n769 VSUBS 0.007488f
C902 B.n770 VSUBS 0.007488f
C903 B.n771 VSUBS 0.007488f
C904 B.n772 VSUBS 0.007488f
C905 B.n773 VSUBS 0.007488f
C906 B.n774 VSUBS 0.007488f
C907 B.n775 VSUBS 0.007488f
C908 B.n776 VSUBS 0.007488f
C909 B.n777 VSUBS 0.007488f
C910 B.n778 VSUBS 0.007488f
C911 B.n779 VSUBS 0.007488f
C912 B.n780 VSUBS 0.004184f
C913 B.n781 VSUBS 0.007488f
C914 B.n782 VSUBS 0.007488f
C915 B.n783 VSUBS 0.007047f
C916 B.n784 VSUBS 0.007488f
C917 B.n785 VSUBS 0.007488f
C918 B.n786 VSUBS 0.007488f
C919 B.n787 VSUBS 0.007488f
C920 B.n788 VSUBS 0.007488f
C921 B.n789 VSUBS 0.007488f
C922 B.n790 VSUBS 0.007488f
C923 B.n791 VSUBS 0.007488f
C924 B.n792 VSUBS 0.007488f
C925 B.n793 VSUBS 0.007488f
C926 B.n794 VSUBS 0.007488f
C927 B.n795 VSUBS 0.007488f
C928 B.n796 VSUBS 0.007488f
C929 B.n797 VSUBS 0.007488f
C930 B.n798 VSUBS 0.007488f
C931 B.n799 VSUBS 0.007488f
C932 B.n800 VSUBS 0.007488f
C933 B.n801 VSUBS 0.007488f
C934 B.n802 VSUBS 0.007488f
C935 B.n803 VSUBS 0.007488f
C936 B.n804 VSUBS 0.007488f
C937 B.n805 VSUBS 0.007488f
C938 B.n806 VSUBS 0.007488f
C939 B.n807 VSUBS 0.007488f
C940 B.n808 VSUBS 0.007488f
C941 B.n809 VSUBS 0.007488f
C942 B.n810 VSUBS 0.007488f
C943 B.n811 VSUBS 0.007488f
C944 B.n812 VSUBS 0.007488f
C945 B.n813 VSUBS 0.007488f
C946 B.n814 VSUBS 0.007488f
C947 B.n815 VSUBS 0.007488f
C948 B.n816 VSUBS 0.007488f
C949 B.n817 VSUBS 0.007488f
C950 B.n818 VSUBS 0.007488f
C951 B.n819 VSUBS 0.007488f
C952 B.n820 VSUBS 0.007488f
C953 B.n821 VSUBS 0.007488f
C954 B.n822 VSUBS 0.007488f
C955 B.n823 VSUBS 0.007488f
C956 B.n824 VSUBS 0.007488f
C957 B.n825 VSUBS 0.007488f
C958 B.n826 VSUBS 0.007488f
C959 B.n827 VSUBS 0.007488f
C960 B.n828 VSUBS 0.007488f
C961 B.n829 VSUBS 0.007488f
C962 B.n830 VSUBS 0.007488f
C963 B.n831 VSUBS 0.007488f
C964 B.n832 VSUBS 0.007488f
C965 B.n833 VSUBS 0.007488f
C966 B.n834 VSUBS 0.007488f
C967 B.n835 VSUBS 0.007488f
C968 B.n836 VSUBS 0.007488f
C969 B.n837 VSUBS 0.007488f
C970 B.n838 VSUBS 0.007488f
C971 B.n839 VSUBS 0.007488f
C972 B.n840 VSUBS 0.007488f
C973 B.n841 VSUBS 0.007488f
C974 B.n842 VSUBS 0.007488f
C975 B.n843 VSUBS 0.007488f
C976 B.n844 VSUBS 0.007488f
C977 B.n845 VSUBS 0.007488f
C978 B.n846 VSUBS 0.007488f
C979 B.n847 VSUBS 0.007488f
C980 B.n848 VSUBS 0.007488f
C981 B.n849 VSUBS 0.007488f
C982 B.n850 VSUBS 0.007488f
C983 B.n851 VSUBS 0.007488f
C984 B.n852 VSUBS 0.007488f
C985 B.n853 VSUBS 0.007488f
C986 B.n854 VSUBS 0.018296f
C987 B.n855 VSUBS 0.018296f
C988 B.n856 VSUBS 0.017822f
C989 B.n857 VSUBS 0.007488f
C990 B.n858 VSUBS 0.007488f
C991 B.n859 VSUBS 0.007488f
C992 B.n860 VSUBS 0.007488f
C993 B.n861 VSUBS 0.007488f
C994 B.n862 VSUBS 0.007488f
C995 B.n863 VSUBS 0.007488f
C996 B.n864 VSUBS 0.007488f
C997 B.n865 VSUBS 0.007488f
C998 B.n866 VSUBS 0.007488f
C999 B.n867 VSUBS 0.007488f
C1000 B.n868 VSUBS 0.007488f
C1001 B.n869 VSUBS 0.007488f
C1002 B.n870 VSUBS 0.007488f
C1003 B.n871 VSUBS 0.007488f
C1004 B.n872 VSUBS 0.007488f
C1005 B.n873 VSUBS 0.007488f
C1006 B.n874 VSUBS 0.007488f
C1007 B.n875 VSUBS 0.007488f
C1008 B.n876 VSUBS 0.007488f
C1009 B.n877 VSUBS 0.007488f
C1010 B.n878 VSUBS 0.007488f
C1011 B.n879 VSUBS 0.007488f
C1012 B.n880 VSUBS 0.007488f
C1013 B.n881 VSUBS 0.007488f
C1014 B.n882 VSUBS 0.007488f
C1015 B.n883 VSUBS 0.007488f
C1016 B.n884 VSUBS 0.007488f
C1017 B.n885 VSUBS 0.007488f
C1018 B.n886 VSUBS 0.007488f
C1019 B.n887 VSUBS 0.007488f
C1020 B.n888 VSUBS 0.007488f
C1021 B.n889 VSUBS 0.007488f
C1022 B.n890 VSUBS 0.007488f
C1023 B.n891 VSUBS 0.007488f
C1024 B.n892 VSUBS 0.007488f
C1025 B.n893 VSUBS 0.007488f
C1026 B.n894 VSUBS 0.007488f
C1027 B.n895 VSUBS 0.007488f
C1028 B.n896 VSUBS 0.007488f
C1029 B.n897 VSUBS 0.007488f
C1030 B.n898 VSUBS 0.007488f
C1031 B.n899 VSUBS 0.007488f
C1032 B.n900 VSUBS 0.007488f
C1033 B.n901 VSUBS 0.007488f
C1034 B.n902 VSUBS 0.007488f
C1035 B.n903 VSUBS 0.007488f
C1036 B.n904 VSUBS 0.007488f
C1037 B.n905 VSUBS 0.007488f
C1038 B.n906 VSUBS 0.007488f
C1039 B.n907 VSUBS 0.007488f
C1040 B.n908 VSUBS 0.007488f
C1041 B.n909 VSUBS 0.007488f
C1042 B.n910 VSUBS 0.007488f
C1043 B.n911 VSUBS 0.007488f
C1044 B.n912 VSUBS 0.007488f
C1045 B.n913 VSUBS 0.007488f
C1046 B.n914 VSUBS 0.007488f
C1047 B.n915 VSUBS 0.007488f
C1048 B.n916 VSUBS 0.007488f
C1049 B.n917 VSUBS 0.007488f
C1050 B.n918 VSUBS 0.007488f
C1051 B.n919 VSUBS 0.007488f
C1052 B.n920 VSUBS 0.007488f
C1053 B.n921 VSUBS 0.007488f
C1054 B.n922 VSUBS 0.007488f
C1055 B.n923 VSUBS 0.007488f
C1056 B.n924 VSUBS 0.007488f
C1057 B.n925 VSUBS 0.007488f
C1058 B.n926 VSUBS 0.007488f
C1059 B.n927 VSUBS 0.007488f
C1060 B.n928 VSUBS 0.007488f
C1061 B.n929 VSUBS 0.007488f
C1062 B.n930 VSUBS 0.007488f
C1063 B.n931 VSUBS 0.007488f
C1064 B.n932 VSUBS 0.007488f
C1065 B.n933 VSUBS 0.007488f
C1066 B.n934 VSUBS 0.007488f
C1067 B.n935 VSUBS 0.007488f
C1068 B.n936 VSUBS 0.007488f
C1069 B.n937 VSUBS 0.007488f
C1070 B.n938 VSUBS 0.007488f
C1071 B.n939 VSUBS 0.007488f
C1072 B.n940 VSUBS 0.007488f
C1073 B.n941 VSUBS 0.007488f
C1074 B.n942 VSUBS 0.007488f
C1075 B.n943 VSUBS 0.007488f
C1076 B.n944 VSUBS 0.007488f
C1077 B.n945 VSUBS 0.007488f
C1078 B.n946 VSUBS 0.007488f
C1079 B.n947 VSUBS 0.007488f
C1080 B.n948 VSUBS 0.007488f
C1081 B.n949 VSUBS 0.007488f
C1082 B.n950 VSUBS 0.007488f
C1083 B.n951 VSUBS 0.016955f
C1084 VDD1.t0 VSUBS 0.346006f
C1085 VDD1.t2 VSUBS 0.346006f
C1086 VDD1.n0 VSUBS 2.82255f
C1087 VDD1.t4 VSUBS 0.346006f
C1088 VDD1.t6 VSUBS 0.346006f
C1089 VDD1.n1 VSUBS 2.8207f
C1090 VDD1.t1 VSUBS 0.346006f
C1091 VDD1.t7 VSUBS 0.346006f
C1092 VDD1.n2 VSUBS 2.8207f
C1093 VDD1.n3 VSUBS 5.37198f
C1094 VDD1.t3 VSUBS 0.346006f
C1095 VDD1.t5 VSUBS 0.346006f
C1096 VDD1.n4 VSUBS 2.7984f
C1097 VDD1.n5 VSUBS 4.45999f
C1098 VTAIL.t4 VSUBS 0.288917f
C1099 VTAIL.t7 VSUBS 0.288917f
C1100 VTAIL.n0 VSUBS 2.19191f
C1101 VTAIL.n1 VSUBS 0.850017f
C1102 VTAIL.n2 VSUBS 0.025307f
C1103 VTAIL.n3 VSUBS 0.024956f
C1104 VTAIL.n4 VSUBS 0.01341f
C1105 VTAIL.n5 VSUBS 0.031698f
C1106 VTAIL.n6 VSUBS 0.014199f
C1107 VTAIL.n7 VSUBS 0.024956f
C1108 VTAIL.n8 VSUBS 0.01341f
C1109 VTAIL.n9 VSUBS 0.031698f
C1110 VTAIL.n10 VSUBS 0.014199f
C1111 VTAIL.n11 VSUBS 0.024956f
C1112 VTAIL.n12 VSUBS 0.01341f
C1113 VTAIL.n13 VSUBS 0.031698f
C1114 VTAIL.n14 VSUBS 0.014199f
C1115 VTAIL.n15 VSUBS 0.024956f
C1116 VTAIL.n16 VSUBS 0.01341f
C1117 VTAIL.n17 VSUBS 0.031698f
C1118 VTAIL.n18 VSUBS 0.014199f
C1119 VTAIL.n19 VSUBS 0.024956f
C1120 VTAIL.n20 VSUBS 0.01341f
C1121 VTAIL.n21 VSUBS 0.031698f
C1122 VTAIL.n22 VSUBS 0.014199f
C1123 VTAIL.n23 VSUBS 0.024956f
C1124 VTAIL.n24 VSUBS 0.01341f
C1125 VTAIL.n25 VSUBS 0.031698f
C1126 VTAIL.n26 VSUBS 0.014199f
C1127 VTAIL.n27 VSUBS 0.173345f
C1128 VTAIL.t1 VSUBS 0.067836f
C1129 VTAIL.n28 VSUBS 0.023773f
C1130 VTAIL.n29 VSUBS 0.020164f
C1131 VTAIL.n30 VSUBS 0.01341f
C1132 VTAIL.n31 VSUBS 1.55386f
C1133 VTAIL.n32 VSUBS 0.024956f
C1134 VTAIL.n33 VSUBS 0.01341f
C1135 VTAIL.n34 VSUBS 0.014199f
C1136 VTAIL.n35 VSUBS 0.031698f
C1137 VTAIL.n36 VSUBS 0.031698f
C1138 VTAIL.n37 VSUBS 0.014199f
C1139 VTAIL.n38 VSUBS 0.01341f
C1140 VTAIL.n39 VSUBS 0.024956f
C1141 VTAIL.n40 VSUBS 0.024956f
C1142 VTAIL.n41 VSUBS 0.01341f
C1143 VTAIL.n42 VSUBS 0.014199f
C1144 VTAIL.n43 VSUBS 0.031698f
C1145 VTAIL.n44 VSUBS 0.031698f
C1146 VTAIL.n45 VSUBS 0.014199f
C1147 VTAIL.n46 VSUBS 0.01341f
C1148 VTAIL.n47 VSUBS 0.024956f
C1149 VTAIL.n48 VSUBS 0.024956f
C1150 VTAIL.n49 VSUBS 0.01341f
C1151 VTAIL.n50 VSUBS 0.014199f
C1152 VTAIL.n51 VSUBS 0.031698f
C1153 VTAIL.n52 VSUBS 0.031698f
C1154 VTAIL.n53 VSUBS 0.014199f
C1155 VTAIL.n54 VSUBS 0.01341f
C1156 VTAIL.n55 VSUBS 0.024956f
C1157 VTAIL.n56 VSUBS 0.024956f
C1158 VTAIL.n57 VSUBS 0.01341f
C1159 VTAIL.n58 VSUBS 0.014199f
C1160 VTAIL.n59 VSUBS 0.031698f
C1161 VTAIL.n60 VSUBS 0.031698f
C1162 VTAIL.n61 VSUBS 0.014199f
C1163 VTAIL.n62 VSUBS 0.01341f
C1164 VTAIL.n63 VSUBS 0.024956f
C1165 VTAIL.n64 VSUBS 0.024956f
C1166 VTAIL.n65 VSUBS 0.01341f
C1167 VTAIL.n66 VSUBS 0.014199f
C1168 VTAIL.n67 VSUBS 0.031698f
C1169 VTAIL.n68 VSUBS 0.031698f
C1170 VTAIL.n69 VSUBS 0.031698f
C1171 VTAIL.n70 VSUBS 0.014199f
C1172 VTAIL.n71 VSUBS 0.01341f
C1173 VTAIL.n72 VSUBS 0.024956f
C1174 VTAIL.n73 VSUBS 0.024956f
C1175 VTAIL.n74 VSUBS 0.01341f
C1176 VTAIL.n75 VSUBS 0.013805f
C1177 VTAIL.n76 VSUBS 0.013805f
C1178 VTAIL.n77 VSUBS 0.031698f
C1179 VTAIL.n78 VSUBS 0.069534f
C1180 VTAIL.n79 VSUBS 0.014199f
C1181 VTAIL.n80 VSUBS 0.01341f
C1182 VTAIL.n81 VSUBS 0.058026f
C1183 VTAIL.n82 VSUBS 0.034659f
C1184 VTAIL.n83 VSUBS 0.317864f
C1185 VTAIL.n84 VSUBS 0.025307f
C1186 VTAIL.n85 VSUBS 0.024956f
C1187 VTAIL.n86 VSUBS 0.01341f
C1188 VTAIL.n87 VSUBS 0.031698f
C1189 VTAIL.n88 VSUBS 0.014199f
C1190 VTAIL.n89 VSUBS 0.024956f
C1191 VTAIL.n90 VSUBS 0.01341f
C1192 VTAIL.n91 VSUBS 0.031698f
C1193 VTAIL.n92 VSUBS 0.014199f
C1194 VTAIL.n93 VSUBS 0.024956f
C1195 VTAIL.n94 VSUBS 0.01341f
C1196 VTAIL.n95 VSUBS 0.031698f
C1197 VTAIL.n96 VSUBS 0.014199f
C1198 VTAIL.n97 VSUBS 0.024956f
C1199 VTAIL.n98 VSUBS 0.01341f
C1200 VTAIL.n99 VSUBS 0.031698f
C1201 VTAIL.n100 VSUBS 0.014199f
C1202 VTAIL.n101 VSUBS 0.024956f
C1203 VTAIL.n102 VSUBS 0.01341f
C1204 VTAIL.n103 VSUBS 0.031698f
C1205 VTAIL.n104 VSUBS 0.014199f
C1206 VTAIL.n105 VSUBS 0.024956f
C1207 VTAIL.n106 VSUBS 0.01341f
C1208 VTAIL.n107 VSUBS 0.031698f
C1209 VTAIL.n108 VSUBS 0.014199f
C1210 VTAIL.n109 VSUBS 0.173345f
C1211 VTAIL.t10 VSUBS 0.067836f
C1212 VTAIL.n110 VSUBS 0.023773f
C1213 VTAIL.n111 VSUBS 0.020164f
C1214 VTAIL.n112 VSUBS 0.01341f
C1215 VTAIL.n113 VSUBS 1.55386f
C1216 VTAIL.n114 VSUBS 0.024956f
C1217 VTAIL.n115 VSUBS 0.01341f
C1218 VTAIL.n116 VSUBS 0.014199f
C1219 VTAIL.n117 VSUBS 0.031698f
C1220 VTAIL.n118 VSUBS 0.031698f
C1221 VTAIL.n119 VSUBS 0.014199f
C1222 VTAIL.n120 VSUBS 0.01341f
C1223 VTAIL.n121 VSUBS 0.024956f
C1224 VTAIL.n122 VSUBS 0.024956f
C1225 VTAIL.n123 VSUBS 0.01341f
C1226 VTAIL.n124 VSUBS 0.014199f
C1227 VTAIL.n125 VSUBS 0.031698f
C1228 VTAIL.n126 VSUBS 0.031698f
C1229 VTAIL.n127 VSUBS 0.014199f
C1230 VTAIL.n128 VSUBS 0.01341f
C1231 VTAIL.n129 VSUBS 0.024956f
C1232 VTAIL.n130 VSUBS 0.024956f
C1233 VTAIL.n131 VSUBS 0.01341f
C1234 VTAIL.n132 VSUBS 0.014199f
C1235 VTAIL.n133 VSUBS 0.031698f
C1236 VTAIL.n134 VSUBS 0.031698f
C1237 VTAIL.n135 VSUBS 0.014199f
C1238 VTAIL.n136 VSUBS 0.01341f
C1239 VTAIL.n137 VSUBS 0.024956f
C1240 VTAIL.n138 VSUBS 0.024956f
C1241 VTAIL.n139 VSUBS 0.01341f
C1242 VTAIL.n140 VSUBS 0.014199f
C1243 VTAIL.n141 VSUBS 0.031698f
C1244 VTAIL.n142 VSUBS 0.031698f
C1245 VTAIL.n143 VSUBS 0.014199f
C1246 VTAIL.n144 VSUBS 0.01341f
C1247 VTAIL.n145 VSUBS 0.024956f
C1248 VTAIL.n146 VSUBS 0.024956f
C1249 VTAIL.n147 VSUBS 0.01341f
C1250 VTAIL.n148 VSUBS 0.014199f
C1251 VTAIL.n149 VSUBS 0.031698f
C1252 VTAIL.n150 VSUBS 0.031698f
C1253 VTAIL.n151 VSUBS 0.031698f
C1254 VTAIL.n152 VSUBS 0.014199f
C1255 VTAIL.n153 VSUBS 0.01341f
C1256 VTAIL.n154 VSUBS 0.024956f
C1257 VTAIL.n155 VSUBS 0.024956f
C1258 VTAIL.n156 VSUBS 0.01341f
C1259 VTAIL.n157 VSUBS 0.013805f
C1260 VTAIL.n158 VSUBS 0.013805f
C1261 VTAIL.n159 VSUBS 0.031698f
C1262 VTAIL.n160 VSUBS 0.069534f
C1263 VTAIL.n161 VSUBS 0.014199f
C1264 VTAIL.n162 VSUBS 0.01341f
C1265 VTAIL.n163 VSUBS 0.058026f
C1266 VTAIL.n164 VSUBS 0.034659f
C1267 VTAIL.n165 VSUBS 0.317864f
C1268 VTAIL.t9 VSUBS 0.288917f
C1269 VTAIL.t11 VSUBS 0.288917f
C1270 VTAIL.n166 VSUBS 2.19191f
C1271 VTAIL.n167 VSUBS 1.10391f
C1272 VTAIL.n168 VSUBS 0.025307f
C1273 VTAIL.n169 VSUBS 0.024956f
C1274 VTAIL.n170 VSUBS 0.01341f
C1275 VTAIL.n171 VSUBS 0.031698f
C1276 VTAIL.n172 VSUBS 0.014199f
C1277 VTAIL.n173 VSUBS 0.024956f
C1278 VTAIL.n174 VSUBS 0.01341f
C1279 VTAIL.n175 VSUBS 0.031698f
C1280 VTAIL.n176 VSUBS 0.014199f
C1281 VTAIL.n177 VSUBS 0.024956f
C1282 VTAIL.n178 VSUBS 0.01341f
C1283 VTAIL.n179 VSUBS 0.031698f
C1284 VTAIL.n180 VSUBS 0.014199f
C1285 VTAIL.n181 VSUBS 0.024956f
C1286 VTAIL.n182 VSUBS 0.01341f
C1287 VTAIL.n183 VSUBS 0.031698f
C1288 VTAIL.n184 VSUBS 0.014199f
C1289 VTAIL.n185 VSUBS 0.024956f
C1290 VTAIL.n186 VSUBS 0.01341f
C1291 VTAIL.n187 VSUBS 0.031698f
C1292 VTAIL.n188 VSUBS 0.014199f
C1293 VTAIL.n189 VSUBS 0.024956f
C1294 VTAIL.n190 VSUBS 0.01341f
C1295 VTAIL.n191 VSUBS 0.031698f
C1296 VTAIL.n192 VSUBS 0.014199f
C1297 VTAIL.n193 VSUBS 0.173345f
C1298 VTAIL.t14 VSUBS 0.067836f
C1299 VTAIL.n194 VSUBS 0.023773f
C1300 VTAIL.n195 VSUBS 0.020164f
C1301 VTAIL.n196 VSUBS 0.01341f
C1302 VTAIL.n197 VSUBS 1.55386f
C1303 VTAIL.n198 VSUBS 0.024956f
C1304 VTAIL.n199 VSUBS 0.01341f
C1305 VTAIL.n200 VSUBS 0.014199f
C1306 VTAIL.n201 VSUBS 0.031698f
C1307 VTAIL.n202 VSUBS 0.031698f
C1308 VTAIL.n203 VSUBS 0.014199f
C1309 VTAIL.n204 VSUBS 0.01341f
C1310 VTAIL.n205 VSUBS 0.024956f
C1311 VTAIL.n206 VSUBS 0.024956f
C1312 VTAIL.n207 VSUBS 0.01341f
C1313 VTAIL.n208 VSUBS 0.014199f
C1314 VTAIL.n209 VSUBS 0.031698f
C1315 VTAIL.n210 VSUBS 0.031698f
C1316 VTAIL.n211 VSUBS 0.014199f
C1317 VTAIL.n212 VSUBS 0.01341f
C1318 VTAIL.n213 VSUBS 0.024956f
C1319 VTAIL.n214 VSUBS 0.024956f
C1320 VTAIL.n215 VSUBS 0.01341f
C1321 VTAIL.n216 VSUBS 0.014199f
C1322 VTAIL.n217 VSUBS 0.031698f
C1323 VTAIL.n218 VSUBS 0.031698f
C1324 VTAIL.n219 VSUBS 0.014199f
C1325 VTAIL.n220 VSUBS 0.01341f
C1326 VTAIL.n221 VSUBS 0.024956f
C1327 VTAIL.n222 VSUBS 0.024956f
C1328 VTAIL.n223 VSUBS 0.01341f
C1329 VTAIL.n224 VSUBS 0.014199f
C1330 VTAIL.n225 VSUBS 0.031698f
C1331 VTAIL.n226 VSUBS 0.031698f
C1332 VTAIL.n227 VSUBS 0.014199f
C1333 VTAIL.n228 VSUBS 0.01341f
C1334 VTAIL.n229 VSUBS 0.024956f
C1335 VTAIL.n230 VSUBS 0.024956f
C1336 VTAIL.n231 VSUBS 0.01341f
C1337 VTAIL.n232 VSUBS 0.014199f
C1338 VTAIL.n233 VSUBS 0.031698f
C1339 VTAIL.n234 VSUBS 0.031698f
C1340 VTAIL.n235 VSUBS 0.031698f
C1341 VTAIL.n236 VSUBS 0.014199f
C1342 VTAIL.n237 VSUBS 0.01341f
C1343 VTAIL.n238 VSUBS 0.024956f
C1344 VTAIL.n239 VSUBS 0.024956f
C1345 VTAIL.n240 VSUBS 0.01341f
C1346 VTAIL.n241 VSUBS 0.013805f
C1347 VTAIL.n242 VSUBS 0.013805f
C1348 VTAIL.n243 VSUBS 0.031698f
C1349 VTAIL.n244 VSUBS 0.069534f
C1350 VTAIL.n245 VSUBS 0.014199f
C1351 VTAIL.n246 VSUBS 0.01341f
C1352 VTAIL.n247 VSUBS 0.058026f
C1353 VTAIL.n248 VSUBS 0.034659f
C1354 VTAIL.n249 VSUBS 1.89325f
C1355 VTAIL.n250 VSUBS 0.025307f
C1356 VTAIL.n251 VSUBS 0.024956f
C1357 VTAIL.n252 VSUBS 0.01341f
C1358 VTAIL.n253 VSUBS 0.031698f
C1359 VTAIL.n254 VSUBS 0.014199f
C1360 VTAIL.n255 VSUBS 0.024956f
C1361 VTAIL.n256 VSUBS 0.01341f
C1362 VTAIL.n257 VSUBS 0.031698f
C1363 VTAIL.n258 VSUBS 0.031698f
C1364 VTAIL.n259 VSUBS 0.014199f
C1365 VTAIL.n260 VSUBS 0.024956f
C1366 VTAIL.n261 VSUBS 0.01341f
C1367 VTAIL.n262 VSUBS 0.031698f
C1368 VTAIL.n263 VSUBS 0.014199f
C1369 VTAIL.n264 VSUBS 0.024956f
C1370 VTAIL.n265 VSUBS 0.01341f
C1371 VTAIL.n266 VSUBS 0.031698f
C1372 VTAIL.n267 VSUBS 0.014199f
C1373 VTAIL.n268 VSUBS 0.024956f
C1374 VTAIL.n269 VSUBS 0.01341f
C1375 VTAIL.n270 VSUBS 0.031698f
C1376 VTAIL.n271 VSUBS 0.014199f
C1377 VTAIL.n272 VSUBS 0.024956f
C1378 VTAIL.n273 VSUBS 0.01341f
C1379 VTAIL.n274 VSUBS 0.031698f
C1380 VTAIL.n275 VSUBS 0.014199f
C1381 VTAIL.n276 VSUBS 0.173345f
C1382 VTAIL.t3 VSUBS 0.067836f
C1383 VTAIL.n277 VSUBS 0.023773f
C1384 VTAIL.n278 VSUBS 0.020164f
C1385 VTAIL.n279 VSUBS 0.01341f
C1386 VTAIL.n280 VSUBS 1.55386f
C1387 VTAIL.n281 VSUBS 0.024956f
C1388 VTAIL.n282 VSUBS 0.01341f
C1389 VTAIL.n283 VSUBS 0.014199f
C1390 VTAIL.n284 VSUBS 0.031698f
C1391 VTAIL.n285 VSUBS 0.031698f
C1392 VTAIL.n286 VSUBS 0.014199f
C1393 VTAIL.n287 VSUBS 0.01341f
C1394 VTAIL.n288 VSUBS 0.024956f
C1395 VTAIL.n289 VSUBS 0.024956f
C1396 VTAIL.n290 VSUBS 0.01341f
C1397 VTAIL.n291 VSUBS 0.014199f
C1398 VTAIL.n292 VSUBS 0.031698f
C1399 VTAIL.n293 VSUBS 0.031698f
C1400 VTAIL.n294 VSUBS 0.014199f
C1401 VTAIL.n295 VSUBS 0.01341f
C1402 VTAIL.n296 VSUBS 0.024956f
C1403 VTAIL.n297 VSUBS 0.024956f
C1404 VTAIL.n298 VSUBS 0.01341f
C1405 VTAIL.n299 VSUBS 0.014199f
C1406 VTAIL.n300 VSUBS 0.031698f
C1407 VTAIL.n301 VSUBS 0.031698f
C1408 VTAIL.n302 VSUBS 0.014199f
C1409 VTAIL.n303 VSUBS 0.01341f
C1410 VTAIL.n304 VSUBS 0.024956f
C1411 VTAIL.n305 VSUBS 0.024956f
C1412 VTAIL.n306 VSUBS 0.01341f
C1413 VTAIL.n307 VSUBS 0.014199f
C1414 VTAIL.n308 VSUBS 0.031698f
C1415 VTAIL.n309 VSUBS 0.031698f
C1416 VTAIL.n310 VSUBS 0.014199f
C1417 VTAIL.n311 VSUBS 0.01341f
C1418 VTAIL.n312 VSUBS 0.024956f
C1419 VTAIL.n313 VSUBS 0.024956f
C1420 VTAIL.n314 VSUBS 0.01341f
C1421 VTAIL.n315 VSUBS 0.014199f
C1422 VTAIL.n316 VSUBS 0.031698f
C1423 VTAIL.n317 VSUBS 0.031698f
C1424 VTAIL.n318 VSUBS 0.014199f
C1425 VTAIL.n319 VSUBS 0.01341f
C1426 VTAIL.n320 VSUBS 0.024956f
C1427 VTAIL.n321 VSUBS 0.024956f
C1428 VTAIL.n322 VSUBS 0.01341f
C1429 VTAIL.n323 VSUBS 0.013805f
C1430 VTAIL.n324 VSUBS 0.013805f
C1431 VTAIL.n325 VSUBS 0.031698f
C1432 VTAIL.n326 VSUBS 0.069534f
C1433 VTAIL.n327 VSUBS 0.014199f
C1434 VTAIL.n328 VSUBS 0.01341f
C1435 VTAIL.n329 VSUBS 0.058026f
C1436 VTAIL.n330 VSUBS 0.034659f
C1437 VTAIL.n331 VSUBS 1.89325f
C1438 VTAIL.t6 VSUBS 0.288917f
C1439 VTAIL.t0 VSUBS 0.288917f
C1440 VTAIL.n332 VSUBS 2.19192f
C1441 VTAIL.n333 VSUBS 1.1039f
C1442 VTAIL.n334 VSUBS 0.025307f
C1443 VTAIL.n335 VSUBS 0.024956f
C1444 VTAIL.n336 VSUBS 0.01341f
C1445 VTAIL.n337 VSUBS 0.031698f
C1446 VTAIL.n338 VSUBS 0.014199f
C1447 VTAIL.n339 VSUBS 0.024956f
C1448 VTAIL.n340 VSUBS 0.01341f
C1449 VTAIL.n341 VSUBS 0.031698f
C1450 VTAIL.n342 VSUBS 0.031698f
C1451 VTAIL.n343 VSUBS 0.014199f
C1452 VTAIL.n344 VSUBS 0.024956f
C1453 VTAIL.n345 VSUBS 0.01341f
C1454 VTAIL.n346 VSUBS 0.031698f
C1455 VTAIL.n347 VSUBS 0.014199f
C1456 VTAIL.n348 VSUBS 0.024956f
C1457 VTAIL.n349 VSUBS 0.01341f
C1458 VTAIL.n350 VSUBS 0.031698f
C1459 VTAIL.n351 VSUBS 0.014199f
C1460 VTAIL.n352 VSUBS 0.024956f
C1461 VTAIL.n353 VSUBS 0.01341f
C1462 VTAIL.n354 VSUBS 0.031698f
C1463 VTAIL.n355 VSUBS 0.014199f
C1464 VTAIL.n356 VSUBS 0.024956f
C1465 VTAIL.n357 VSUBS 0.01341f
C1466 VTAIL.n358 VSUBS 0.031698f
C1467 VTAIL.n359 VSUBS 0.014199f
C1468 VTAIL.n360 VSUBS 0.173345f
C1469 VTAIL.t5 VSUBS 0.067836f
C1470 VTAIL.n361 VSUBS 0.023773f
C1471 VTAIL.n362 VSUBS 0.020164f
C1472 VTAIL.n363 VSUBS 0.01341f
C1473 VTAIL.n364 VSUBS 1.55386f
C1474 VTAIL.n365 VSUBS 0.024956f
C1475 VTAIL.n366 VSUBS 0.01341f
C1476 VTAIL.n367 VSUBS 0.014199f
C1477 VTAIL.n368 VSUBS 0.031698f
C1478 VTAIL.n369 VSUBS 0.031698f
C1479 VTAIL.n370 VSUBS 0.014199f
C1480 VTAIL.n371 VSUBS 0.01341f
C1481 VTAIL.n372 VSUBS 0.024956f
C1482 VTAIL.n373 VSUBS 0.024956f
C1483 VTAIL.n374 VSUBS 0.01341f
C1484 VTAIL.n375 VSUBS 0.014199f
C1485 VTAIL.n376 VSUBS 0.031698f
C1486 VTAIL.n377 VSUBS 0.031698f
C1487 VTAIL.n378 VSUBS 0.014199f
C1488 VTAIL.n379 VSUBS 0.01341f
C1489 VTAIL.n380 VSUBS 0.024956f
C1490 VTAIL.n381 VSUBS 0.024956f
C1491 VTAIL.n382 VSUBS 0.01341f
C1492 VTAIL.n383 VSUBS 0.014199f
C1493 VTAIL.n384 VSUBS 0.031698f
C1494 VTAIL.n385 VSUBS 0.031698f
C1495 VTAIL.n386 VSUBS 0.014199f
C1496 VTAIL.n387 VSUBS 0.01341f
C1497 VTAIL.n388 VSUBS 0.024956f
C1498 VTAIL.n389 VSUBS 0.024956f
C1499 VTAIL.n390 VSUBS 0.01341f
C1500 VTAIL.n391 VSUBS 0.014199f
C1501 VTAIL.n392 VSUBS 0.031698f
C1502 VTAIL.n393 VSUBS 0.031698f
C1503 VTAIL.n394 VSUBS 0.014199f
C1504 VTAIL.n395 VSUBS 0.01341f
C1505 VTAIL.n396 VSUBS 0.024956f
C1506 VTAIL.n397 VSUBS 0.024956f
C1507 VTAIL.n398 VSUBS 0.01341f
C1508 VTAIL.n399 VSUBS 0.014199f
C1509 VTAIL.n400 VSUBS 0.031698f
C1510 VTAIL.n401 VSUBS 0.031698f
C1511 VTAIL.n402 VSUBS 0.014199f
C1512 VTAIL.n403 VSUBS 0.01341f
C1513 VTAIL.n404 VSUBS 0.024956f
C1514 VTAIL.n405 VSUBS 0.024956f
C1515 VTAIL.n406 VSUBS 0.01341f
C1516 VTAIL.n407 VSUBS 0.013805f
C1517 VTAIL.n408 VSUBS 0.013805f
C1518 VTAIL.n409 VSUBS 0.031698f
C1519 VTAIL.n410 VSUBS 0.069534f
C1520 VTAIL.n411 VSUBS 0.014199f
C1521 VTAIL.n412 VSUBS 0.01341f
C1522 VTAIL.n413 VSUBS 0.058026f
C1523 VTAIL.n414 VSUBS 0.034659f
C1524 VTAIL.n415 VSUBS 0.317864f
C1525 VTAIL.n416 VSUBS 0.025307f
C1526 VTAIL.n417 VSUBS 0.024956f
C1527 VTAIL.n418 VSUBS 0.01341f
C1528 VTAIL.n419 VSUBS 0.031698f
C1529 VTAIL.n420 VSUBS 0.014199f
C1530 VTAIL.n421 VSUBS 0.024956f
C1531 VTAIL.n422 VSUBS 0.01341f
C1532 VTAIL.n423 VSUBS 0.031698f
C1533 VTAIL.n424 VSUBS 0.031698f
C1534 VTAIL.n425 VSUBS 0.014199f
C1535 VTAIL.n426 VSUBS 0.024956f
C1536 VTAIL.n427 VSUBS 0.01341f
C1537 VTAIL.n428 VSUBS 0.031698f
C1538 VTAIL.n429 VSUBS 0.014199f
C1539 VTAIL.n430 VSUBS 0.024956f
C1540 VTAIL.n431 VSUBS 0.01341f
C1541 VTAIL.n432 VSUBS 0.031698f
C1542 VTAIL.n433 VSUBS 0.014199f
C1543 VTAIL.n434 VSUBS 0.024956f
C1544 VTAIL.n435 VSUBS 0.01341f
C1545 VTAIL.n436 VSUBS 0.031698f
C1546 VTAIL.n437 VSUBS 0.014199f
C1547 VTAIL.n438 VSUBS 0.024956f
C1548 VTAIL.n439 VSUBS 0.01341f
C1549 VTAIL.n440 VSUBS 0.031698f
C1550 VTAIL.n441 VSUBS 0.014199f
C1551 VTAIL.n442 VSUBS 0.173345f
C1552 VTAIL.t12 VSUBS 0.067836f
C1553 VTAIL.n443 VSUBS 0.023773f
C1554 VTAIL.n444 VSUBS 0.020164f
C1555 VTAIL.n445 VSUBS 0.01341f
C1556 VTAIL.n446 VSUBS 1.55386f
C1557 VTAIL.n447 VSUBS 0.024956f
C1558 VTAIL.n448 VSUBS 0.01341f
C1559 VTAIL.n449 VSUBS 0.014199f
C1560 VTAIL.n450 VSUBS 0.031698f
C1561 VTAIL.n451 VSUBS 0.031698f
C1562 VTAIL.n452 VSUBS 0.014199f
C1563 VTAIL.n453 VSUBS 0.01341f
C1564 VTAIL.n454 VSUBS 0.024956f
C1565 VTAIL.n455 VSUBS 0.024956f
C1566 VTAIL.n456 VSUBS 0.01341f
C1567 VTAIL.n457 VSUBS 0.014199f
C1568 VTAIL.n458 VSUBS 0.031698f
C1569 VTAIL.n459 VSUBS 0.031698f
C1570 VTAIL.n460 VSUBS 0.014199f
C1571 VTAIL.n461 VSUBS 0.01341f
C1572 VTAIL.n462 VSUBS 0.024956f
C1573 VTAIL.n463 VSUBS 0.024956f
C1574 VTAIL.n464 VSUBS 0.01341f
C1575 VTAIL.n465 VSUBS 0.014199f
C1576 VTAIL.n466 VSUBS 0.031698f
C1577 VTAIL.n467 VSUBS 0.031698f
C1578 VTAIL.n468 VSUBS 0.014199f
C1579 VTAIL.n469 VSUBS 0.01341f
C1580 VTAIL.n470 VSUBS 0.024956f
C1581 VTAIL.n471 VSUBS 0.024956f
C1582 VTAIL.n472 VSUBS 0.01341f
C1583 VTAIL.n473 VSUBS 0.014199f
C1584 VTAIL.n474 VSUBS 0.031698f
C1585 VTAIL.n475 VSUBS 0.031698f
C1586 VTAIL.n476 VSUBS 0.014199f
C1587 VTAIL.n477 VSUBS 0.01341f
C1588 VTAIL.n478 VSUBS 0.024956f
C1589 VTAIL.n479 VSUBS 0.024956f
C1590 VTAIL.n480 VSUBS 0.01341f
C1591 VTAIL.n481 VSUBS 0.014199f
C1592 VTAIL.n482 VSUBS 0.031698f
C1593 VTAIL.n483 VSUBS 0.031698f
C1594 VTAIL.n484 VSUBS 0.014199f
C1595 VTAIL.n485 VSUBS 0.01341f
C1596 VTAIL.n486 VSUBS 0.024956f
C1597 VTAIL.n487 VSUBS 0.024956f
C1598 VTAIL.n488 VSUBS 0.01341f
C1599 VTAIL.n489 VSUBS 0.013805f
C1600 VTAIL.n490 VSUBS 0.013805f
C1601 VTAIL.n491 VSUBS 0.031698f
C1602 VTAIL.n492 VSUBS 0.069534f
C1603 VTAIL.n493 VSUBS 0.014199f
C1604 VTAIL.n494 VSUBS 0.01341f
C1605 VTAIL.n495 VSUBS 0.058026f
C1606 VTAIL.n496 VSUBS 0.034659f
C1607 VTAIL.n497 VSUBS 0.317864f
C1608 VTAIL.t8 VSUBS 0.288917f
C1609 VTAIL.t13 VSUBS 0.288917f
C1610 VTAIL.n498 VSUBS 2.19192f
C1611 VTAIL.n499 VSUBS 1.1039f
C1612 VTAIL.n500 VSUBS 0.025307f
C1613 VTAIL.n501 VSUBS 0.024956f
C1614 VTAIL.n502 VSUBS 0.01341f
C1615 VTAIL.n503 VSUBS 0.031698f
C1616 VTAIL.n504 VSUBS 0.014199f
C1617 VTAIL.n505 VSUBS 0.024956f
C1618 VTAIL.n506 VSUBS 0.01341f
C1619 VTAIL.n507 VSUBS 0.031698f
C1620 VTAIL.n508 VSUBS 0.031698f
C1621 VTAIL.n509 VSUBS 0.014199f
C1622 VTAIL.n510 VSUBS 0.024956f
C1623 VTAIL.n511 VSUBS 0.01341f
C1624 VTAIL.n512 VSUBS 0.031698f
C1625 VTAIL.n513 VSUBS 0.014199f
C1626 VTAIL.n514 VSUBS 0.024956f
C1627 VTAIL.n515 VSUBS 0.01341f
C1628 VTAIL.n516 VSUBS 0.031698f
C1629 VTAIL.n517 VSUBS 0.014199f
C1630 VTAIL.n518 VSUBS 0.024956f
C1631 VTAIL.n519 VSUBS 0.01341f
C1632 VTAIL.n520 VSUBS 0.031698f
C1633 VTAIL.n521 VSUBS 0.014199f
C1634 VTAIL.n522 VSUBS 0.024956f
C1635 VTAIL.n523 VSUBS 0.01341f
C1636 VTAIL.n524 VSUBS 0.031698f
C1637 VTAIL.n525 VSUBS 0.014199f
C1638 VTAIL.n526 VSUBS 0.173345f
C1639 VTAIL.t15 VSUBS 0.067836f
C1640 VTAIL.n527 VSUBS 0.023773f
C1641 VTAIL.n528 VSUBS 0.020164f
C1642 VTAIL.n529 VSUBS 0.01341f
C1643 VTAIL.n530 VSUBS 1.55386f
C1644 VTAIL.n531 VSUBS 0.024956f
C1645 VTAIL.n532 VSUBS 0.01341f
C1646 VTAIL.n533 VSUBS 0.014199f
C1647 VTAIL.n534 VSUBS 0.031698f
C1648 VTAIL.n535 VSUBS 0.031698f
C1649 VTAIL.n536 VSUBS 0.014199f
C1650 VTAIL.n537 VSUBS 0.01341f
C1651 VTAIL.n538 VSUBS 0.024956f
C1652 VTAIL.n539 VSUBS 0.024956f
C1653 VTAIL.n540 VSUBS 0.01341f
C1654 VTAIL.n541 VSUBS 0.014199f
C1655 VTAIL.n542 VSUBS 0.031698f
C1656 VTAIL.n543 VSUBS 0.031698f
C1657 VTAIL.n544 VSUBS 0.014199f
C1658 VTAIL.n545 VSUBS 0.01341f
C1659 VTAIL.n546 VSUBS 0.024956f
C1660 VTAIL.n547 VSUBS 0.024956f
C1661 VTAIL.n548 VSUBS 0.01341f
C1662 VTAIL.n549 VSUBS 0.014199f
C1663 VTAIL.n550 VSUBS 0.031698f
C1664 VTAIL.n551 VSUBS 0.031698f
C1665 VTAIL.n552 VSUBS 0.014199f
C1666 VTAIL.n553 VSUBS 0.01341f
C1667 VTAIL.n554 VSUBS 0.024956f
C1668 VTAIL.n555 VSUBS 0.024956f
C1669 VTAIL.n556 VSUBS 0.01341f
C1670 VTAIL.n557 VSUBS 0.014199f
C1671 VTAIL.n558 VSUBS 0.031698f
C1672 VTAIL.n559 VSUBS 0.031698f
C1673 VTAIL.n560 VSUBS 0.014199f
C1674 VTAIL.n561 VSUBS 0.01341f
C1675 VTAIL.n562 VSUBS 0.024956f
C1676 VTAIL.n563 VSUBS 0.024956f
C1677 VTAIL.n564 VSUBS 0.01341f
C1678 VTAIL.n565 VSUBS 0.014199f
C1679 VTAIL.n566 VSUBS 0.031698f
C1680 VTAIL.n567 VSUBS 0.031698f
C1681 VTAIL.n568 VSUBS 0.014199f
C1682 VTAIL.n569 VSUBS 0.01341f
C1683 VTAIL.n570 VSUBS 0.024956f
C1684 VTAIL.n571 VSUBS 0.024956f
C1685 VTAIL.n572 VSUBS 0.01341f
C1686 VTAIL.n573 VSUBS 0.013805f
C1687 VTAIL.n574 VSUBS 0.013805f
C1688 VTAIL.n575 VSUBS 0.031698f
C1689 VTAIL.n576 VSUBS 0.069534f
C1690 VTAIL.n577 VSUBS 0.014199f
C1691 VTAIL.n578 VSUBS 0.01341f
C1692 VTAIL.n579 VSUBS 0.058026f
C1693 VTAIL.n580 VSUBS 0.034659f
C1694 VTAIL.n581 VSUBS 1.89325f
C1695 VTAIL.n582 VSUBS 0.025307f
C1696 VTAIL.n583 VSUBS 0.024956f
C1697 VTAIL.n584 VSUBS 0.01341f
C1698 VTAIL.n585 VSUBS 0.031698f
C1699 VTAIL.n586 VSUBS 0.014199f
C1700 VTAIL.n587 VSUBS 0.024956f
C1701 VTAIL.n588 VSUBS 0.01341f
C1702 VTAIL.n589 VSUBS 0.031698f
C1703 VTAIL.n590 VSUBS 0.014199f
C1704 VTAIL.n591 VSUBS 0.024956f
C1705 VTAIL.n592 VSUBS 0.01341f
C1706 VTAIL.n593 VSUBS 0.031698f
C1707 VTAIL.n594 VSUBS 0.014199f
C1708 VTAIL.n595 VSUBS 0.024956f
C1709 VTAIL.n596 VSUBS 0.01341f
C1710 VTAIL.n597 VSUBS 0.031698f
C1711 VTAIL.n598 VSUBS 0.014199f
C1712 VTAIL.n599 VSUBS 0.024956f
C1713 VTAIL.n600 VSUBS 0.01341f
C1714 VTAIL.n601 VSUBS 0.031698f
C1715 VTAIL.n602 VSUBS 0.014199f
C1716 VTAIL.n603 VSUBS 0.024956f
C1717 VTAIL.n604 VSUBS 0.01341f
C1718 VTAIL.n605 VSUBS 0.031698f
C1719 VTAIL.n606 VSUBS 0.014199f
C1720 VTAIL.n607 VSUBS 0.173345f
C1721 VTAIL.t2 VSUBS 0.067836f
C1722 VTAIL.n608 VSUBS 0.023773f
C1723 VTAIL.n609 VSUBS 0.020164f
C1724 VTAIL.n610 VSUBS 0.01341f
C1725 VTAIL.n611 VSUBS 1.55386f
C1726 VTAIL.n612 VSUBS 0.024956f
C1727 VTAIL.n613 VSUBS 0.01341f
C1728 VTAIL.n614 VSUBS 0.014199f
C1729 VTAIL.n615 VSUBS 0.031698f
C1730 VTAIL.n616 VSUBS 0.031698f
C1731 VTAIL.n617 VSUBS 0.014199f
C1732 VTAIL.n618 VSUBS 0.01341f
C1733 VTAIL.n619 VSUBS 0.024956f
C1734 VTAIL.n620 VSUBS 0.024956f
C1735 VTAIL.n621 VSUBS 0.01341f
C1736 VTAIL.n622 VSUBS 0.014199f
C1737 VTAIL.n623 VSUBS 0.031698f
C1738 VTAIL.n624 VSUBS 0.031698f
C1739 VTAIL.n625 VSUBS 0.014199f
C1740 VTAIL.n626 VSUBS 0.01341f
C1741 VTAIL.n627 VSUBS 0.024956f
C1742 VTAIL.n628 VSUBS 0.024956f
C1743 VTAIL.n629 VSUBS 0.01341f
C1744 VTAIL.n630 VSUBS 0.014199f
C1745 VTAIL.n631 VSUBS 0.031698f
C1746 VTAIL.n632 VSUBS 0.031698f
C1747 VTAIL.n633 VSUBS 0.014199f
C1748 VTAIL.n634 VSUBS 0.01341f
C1749 VTAIL.n635 VSUBS 0.024956f
C1750 VTAIL.n636 VSUBS 0.024956f
C1751 VTAIL.n637 VSUBS 0.01341f
C1752 VTAIL.n638 VSUBS 0.014199f
C1753 VTAIL.n639 VSUBS 0.031698f
C1754 VTAIL.n640 VSUBS 0.031698f
C1755 VTAIL.n641 VSUBS 0.014199f
C1756 VTAIL.n642 VSUBS 0.01341f
C1757 VTAIL.n643 VSUBS 0.024956f
C1758 VTAIL.n644 VSUBS 0.024956f
C1759 VTAIL.n645 VSUBS 0.01341f
C1760 VTAIL.n646 VSUBS 0.014199f
C1761 VTAIL.n647 VSUBS 0.031698f
C1762 VTAIL.n648 VSUBS 0.031698f
C1763 VTAIL.n649 VSUBS 0.031698f
C1764 VTAIL.n650 VSUBS 0.014199f
C1765 VTAIL.n651 VSUBS 0.01341f
C1766 VTAIL.n652 VSUBS 0.024956f
C1767 VTAIL.n653 VSUBS 0.024956f
C1768 VTAIL.n654 VSUBS 0.01341f
C1769 VTAIL.n655 VSUBS 0.013805f
C1770 VTAIL.n656 VSUBS 0.013805f
C1771 VTAIL.n657 VSUBS 0.031698f
C1772 VTAIL.n658 VSUBS 0.069534f
C1773 VTAIL.n659 VSUBS 0.014199f
C1774 VTAIL.n660 VSUBS 0.01341f
C1775 VTAIL.n661 VSUBS 0.058026f
C1776 VTAIL.n662 VSUBS 0.034659f
C1777 VTAIL.n663 VSUBS 1.88857f
C1778 VP.t0 VSUBS 3.5108f
C1779 VP.n0 VSUBS 1.32906f
C1780 VP.n1 VSUBS 0.025736f
C1781 VP.n2 VSUBS 0.020938f
C1782 VP.n3 VSUBS 0.025736f
C1783 VP.t6 VSUBS 3.5108f
C1784 VP.n4 VSUBS 1.22119f
C1785 VP.n5 VSUBS 0.025736f
C1786 VP.n6 VSUBS 0.03757f
C1787 VP.n7 VSUBS 0.025736f
C1788 VP.n8 VSUBS 0.02973f
C1789 VP.n9 VSUBS 0.025736f
C1790 VP.n10 VSUBS 0.020938f
C1791 VP.n11 VSUBS 0.025736f
C1792 VP.t3 VSUBS 3.5108f
C1793 VP.n12 VSUBS 1.32906f
C1794 VP.t2 VSUBS 3.5108f
C1795 VP.n13 VSUBS 1.32906f
C1796 VP.n14 VSUBS 0.025736f
C1797 VP.n15 VSUBS 0.020938f
C1798 VP.n16 VSUBS 0.025736f
C1799 VP.t4 VSUBS 3.5108f
C1800 VP.n17 VSUBS 1.22119f
C1801 VP.n18 VSUBS 0.025736f
C1802 VP.n19 VSUBS 0.03757f
C1803 VP.n20 VSUBS 0.025736f
C1804 VP.n21 VSUBS 0.02973f
C1805 VP.t7 VSUBS 3.85168f
C1806 VP.t5 VSUBS 3.5108f
C1807 VP.n22 VSUBS 1.30268f
C1808 VP.n23 VSUBS 1.24449f
C1809 VP.n24 VSUBS 0.304462f
C1810 VP.n25 VSUBS 0.025736f
C1811 VP.n26 VSUBS 0.047966f
C1812 VP.n27 VSUBS 0.047966f
C1813 VP.n28 VSUBS 0.03757f
C1814 VP.n29 VSUBS 0.025736f
C1815 VP.n30 VSUBS 0.025736f
C1816 VP.n31 VSUBS 0.025736f
C1817 VP.n32 VSUBS 0.047966f
C1818 VP.n33 VSUBS 0.047966f
C1819 VP.n34 VSUBS 0.02973f
C1820 VP.n35 VSUBS 0.025736f
C1821 VP.n36 VSUBS 0.025736f
C1822 VP.n37 VSUBS 0.042518f
C1823 VP.n38 VSUBS 0.047966f
C1824 VP.n39 VSUBS 0.050571f
C1825 VP.n40 VSUBS 0.025736f
C1826 VP.n41 VSUBS 0.025736f
C1827 VP.n42 VSUBS 0.025736f
C1828 VP.n43 VSUBS 0.051597f
C1829 VP.n44 VSUBS 0.047966f
C1830 VP.n45 VSUBS 0.040624f
C1831 VP.n46 VSUBS 0.041538f
C1832 VP.n47 VSUBS 1.75115f
C1833 VP.n48 VSUBS 1.76743f
C1834 VP.n49 VSUBS 0.041538f
C1835 VP.n50 VSUBS 0.040624f
C1836 VP.n51 VSUBS 0.047966f
C1837 VP.n52 VSUBS 0.051597f
C1838 VP.n53 VSUBS 0.025736f
C1839 VP.n54 VSUBS 0.025736f
C1840 VP.n55 VSUBS 0.025736f
C1841 VP.n56 VSUBS 0.050571f
C1842 VP.n57 VSUBS 0.047966f
C1843 VP.t1 VSUBS 3.5108f
C1844 VP.n58 VSUBS 1.22119f
C1845 VP.n59 VSUBS 0.042518f
C1846 VP.n60 VSUBS 0.025736f
C1847 VP.n61 VSUBS 0.025736f
C1848 VP.n62 VSUBS 0.025736f
C1849 VP.n63 VSUBS 0.047966f
C1850 VP.n64 VSUBS 0.047966f
C1851 VP.n65 VSUBS 0.03757f
C1852 VP.n66 VSUBS 0.025736f
C1853 VP.n67 VSUBS 0.025736f
C1854 VP.n68 VSUBS 0.025736f
C1855 VP.n69 VSUBS 0.047966f
C1856 VP.n70 VSUBS 0.047966f
C1857 VP.n71 VSUBS 0.02973f
C1858 VP.n72 VSUBS 0.025736f
C1859 VP.n73 VSUBS 0.025736f
C1860 VP.n74 VSUBS 0.042518f
C1861 VP.n75 VSUBS 0.047966f
C1862 VP.n76 VSUBS 0.050571f
C1863 VP.n77 VSUBS 0.025736f
C1864 VP.n78 VSUBS 0.025736f
C1865 VP.n79 VSUBS 0.025736f
C1866 VP.n80 VSUBS 0.051597f
C1867 VP.n81 VSUBS 0.047966f
C1868 VP.n82 VSUBS 0.040624f
C1869 VP.n83 VSUBS 0.041538f
C1870 VP.n84 VSUBS 0.060857f
.ends

