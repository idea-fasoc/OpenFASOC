* NGSPICE file created from diff_pair_sample_0845.ext - technology: sky130A

.subckt diff_pair_sample_0845 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t14 VP.t0 VDD1.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.1582 pd=13.41 as=2.1582 ps=13.41 w=13.08 l=3.31
X1 VDD1.t3 VP.t1 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=2.1582 pd=13.41 as=5.1012 ps=26.94 w=13.08 l=3.31
X2 VTAIL.t12 VP.t2 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=5.1012 pd=26.94 as=2.1582 ps=13.41 w=13.08 l=3.31
X3 VTAIL.t1 VN.t0 VDD2.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=5.1012 pd=26.94 as=2.1582 ps=13.41 w=13.08 l=3.31
X4 VTAIL.t0 VN.t1 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=5.1012 pd=26.94 as=2.1582 ps=13.41 w=13.08 l=3.31
X5 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=5.1012 pd=26.94 as=0 ps=0 w=13.08 l=3.31
X6 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=5.1012 pd=26.94 as=0 ps=0 w=13.08 l=3.31
X7 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=5.1012 pd=26.94 as=0 ps=0 w=13.08 l=3.31
X8 VDD2.t5 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1582 pd=13.41 as=2.1582 ps=13.41 w=13.08 l=3.31
X9 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.1012 pd=26.94 as=0 ps=0 w=13.08 l=3.31
X10 VDD2.t4 VN.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.1582 pd=13.41 as=2.1582 ps=13.41 w=13.08 l=3.31
X11 VTAIL.t11 VP.t3 VDD1.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=2.1582 pd=13.41 as=2.1582 ps=13.41 w=13.08 l=3.31
X12 VTAIL.t15 VN.t4 VDD2.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=2.1582 pd=13.41 as=2.1582 ps=13.41 w=13.08 l=3.31
X13 VDD1.t4 VP.t4 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=2.1582 pd=13.41 as=2.1582 ps=13.41 w=13.08 l=3.31
X14 VDD1.t1 VP.t5 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1582 pd=13.41 as=2.1582 ps=13.41 w=13.08 l=3.31
X15 VDD2.t2 VN.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.1582 pd=13.41 as=5.1012 ps=26.94 w=13.08 l=3.31
X16 VTAIL.t5 VN.t6 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=2.1582 pd=13.41 as=2.1582 ps=13.41 w=13.08 l=3.31
X17 VTAIL.t8 VP.t6 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.1012 pd=26.94 as=2.1582 ps=13.41 w=13.08 l=3.31
X18 VDD1.t7 VP.t7 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=2.1582 pd=13.41 as=5.1012 ps=26.94 w=13.08 l=3.31
X19 VDD2.t0 VN.t7 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.1582 pd=13.41 as=5.1012 ps=26.94 w=13.08 l=3.31
R0 VP.n24 VP.n21 161.3
R1 VP.n26 VP.n25 161.3
R2 VP.n27 VP.n20 161.3
R3 VP.n29 VP.n28 161.3
R4 VP.n30 VP.n19 161.3
R5 VP.n32 VP.n31 161.3
R6 VP.n33 VP.n18 161.3
R7 VP.n35 VP.n34 161.3
R8 VP.n37 VP.n36 161.3
R9 VP.n38 VP.n16 161.3
R10 VP.n40 VP.n39 161.3
R11 VP.n41 VP.n15 161.3
R12 VP.n43 VP.n42 161.3
R13 VP.n44 VP.n14 161.3
R14 VP.n46 VP.n45 161.3
R15 VP.n83 VP.n82 161.3
R16 VP.n81 VP.n1 161.3
R17 VP.n80 VP.n79 161.3
R18 VP.n78 VP.n2 161.3
R19 VP.n77 VP.n76 161.3
R20 VP.n75 VP.n3 161.3
R21 VP.n74 VP.n73 161.3
R22 VP.n72 VP.n71 161.3
R23 VP.n70 VP.n5 161.3
R24 VP.n69 VP.n68 161.3
R25 VP.n67 VP.n6 161.3
R26 VP.n66 VP.n65 161.3
R27 VP.n64 VP.n7 161.3
R28 VP.n63 VP.n62 161.3
R29 VP.n61 VP.n8 161.3
R30 VP.n60 VP.n59 161.3
R31 VP.n57 VP.n9 161.3
R32 VP.n56 VP.n55 161.3
R33 VP.n54 VP.n10 161.3
R34 VP.n53 VP.n52 161.3
R35 VP.n51 VP.n11 161.3
R36 VP.n50 VP.n49 161.3
R37 VP.n23 VP.t6 127.492
R38 VP.n12 VP.t2 95.2355
R39 VP.n58 VP.t5 95.2355
R40 VP.n4 VP.t3 95.2355
R41 VP.n0 VP.t1 95.2355
R42 VP.n13 VP.t7 95.2355
R43 VP.n17 VP.t0 95.2355
R44 VP.n22 VP.t4 95.2355
R45 VP.n48 VP.n12 79.917
R46 VP.n84 VP.n0 79.917
R47 VP.n47 VP.n13 79.917
R48 VP.n23 VP.n22 71.3663
R49 VP.n65 VP.n6 56.5617
R50 VP.n28 VP.n19 56.5617
R51 VP.n48 VP.n47 55.0829
R52 VP.n56 VP.n10 51.2335
R53 VP.n76 VP.n2 51.2335
R54 VP.n39 VP.n15 51.2335
R55 VP.n52 VP.n10 29.9206
R56 VP.n80 VP.n2 29.9206
R57 VP.n43 VP.n15 29.9206
R58 VP.n51 VP.n50 24.5923
R59 VP.n52 VP.n51 24.5923
R60 VP.n57 VP.n56 24.5923
R61 VP.n59 VP.n57 24.5923
R62 VP.n63 VP.n8 24.5923
R63 VP.n64 VP.n63 24.5923
R64 VP.n65 VP.n64 24.5923
R65 VP.n69 VP.n6 24.5923
R66 VP.n70 VP.n69 24.5923
R67 VP.n71 VP.n70 24.5923
R68 VP.n75 VP.n74 24.5923
R69 VP.n76 VP.n75 24.5923
R70 VP.n81 VP.n80 24.5923
R71 VP.n82 VP.n81 24.5923
R72 VP.n44 VP.n43 24.5923
R73 VP.n45 VP.n44 24.5923
R74 VP.n32 VP.n19 24.5923
R75 VP.n33 VP.n32 24.5923
R76 VP.n34 VP.n33 24.5923
R77 VP.n38 VP.n37 24.5923
R78 VP.n39 VP.n38 24.5923
R79 VP.n26 VP.n21 24.5923
R80 VP.n27 VP.n26 24.5923
R81 VP.n28 VP.n27 24.5923
R82 VP.n59 VP.n58 21.1495
R83 VP.n74 VP.n4 21.1495
R84 VP.n37 VP.n17 21.1495
R85 VP.n50 VP.n12 10.3291
R86 VP.n82 VP.n0 10.3291
R87 VP.n45 VP.n13 10.3291
R88 VP.n24 VP.n23 4.37639
R89 VP.n58 VP.n8 3.44336
R90 VP.n71 VP.n4 3.44336
R91 VP.n34 VP.n17 3.44336
R92 VP.n22 VP.n21 3.44336
R93 VP.n47 VP.n46 0.354861
R94 VP.n49 VP.n48 0.354861
R95 VP.n84 VP.n83 0.354861
R96 VP VP.n84 0.267071
R97 VP.n25 VP.n24 0.189894
R98 VP.n25 VP.n20 0.189894
R99 VP.n29 VP.n20 0.189894
R100 VP.n30 VP.n29 0.189894
R101 VP.n31 VP.n30 0.189894
R102 VP.n31 VP.n18 0.189894
R103 VP.n35 VP.n18 0.189894
R104 VP.n36 VP.n35 0.189894
R105 VP.n36 VP.n16 0.189894
R106 VP.n40 VP.n16 0.189894
R107 VP.n41 VP.n40 0.189894
R108 VP.n42 VP.n41 0.189894
R109 VP.n42 VP.n14 0.189894
R110 VP.n46 VP.n14 0.189894
R111 VP.n49 VP.n11 0.189894
R112 VP.n53 VP.n11 0.189894
R113 VP.n54 VP.n53 0.189894
R114 VP.n55 VP.n54 0.189894
R115 VP.n55 VP.n9 0.189894
R116 VP.n60 VP.n9 0.189894
R117 VP.n61 VP.n60 0.189894
R118 VP.n62 VP.n61 0.189894
R119 VP.n62 VP.n7 0.189894
R120 VP.n66 VP.n7 0.189894
R121 VP.n67 VP.n66 0.189894
R122 VP.n68 VP.n67 0.189894
R123 VP.n68 VP.n5 0.189894
R124 VP.n72 VP.n5 0.189894
R125 VP.n73 VP.n72 0.189894
R126 VP.n73 VP.n3 0.189894
R127 VP.n77 VP.n3 0.189894
R128 VP.n78 VP.n77 0.189894
R129 VP.n79 VP.n78 0.189894
R130 VP.n79 VP.n1 0.189894
R131 VP.n83 VP.n1 0.189894
R132 VDD1 VDD1.n0 60.9252
R133 VDD1.n3 VDD1.n2 60.8116
R134 VDD1.n3 VDD1.n1 60.8116
R135 VDD1.n5 VDD1.n4 59.2979
R136 VDD1.n5 VDD1.n3 49.6949
R137 VDD1.n4 VDD1.t6 1.51426
R138 VDD1.n4 VDD1.t7 1.51426
R139 VDD1.n0 VDD1.t0 1.51426
R140 VDD1.n0 VDD1.t4 1.51426
R141 VDD1.n2 VDD1.t5 1.51426
R142 VDD1.n2 VDD1.t3 1.51426
R143 VDD1.n1 VDD1.t2 1.51426
R144 VDD1.n1 VDD1.t1 1.51426
R145 VDD1 VDD1.n5 1.51128
R146 VTAIL.n11 VTAIL.t8 44.133
R147 VTAIL.n10 VTAIL.t3 44.133
R148 VTAIL.n7 VTAIL.t1 44.133
R149 VTAIL.n15 VTAIL.t4 44.1328
R150 VTAIL.n2 VTAIL.t0 44.1328
R151 VTAIL.n3 VTAIL.t13 44.1328
R152 VTAIL.n6 VTAIL.t12 44.1328
R153 VTAIL.n14 VTAIL.t7 44.1328
R154 VTAIL.n13 VTAIL.n12 42.6192
R155 VTAIL.n9 VTAIL.n8 42.6192
R156 VTAIL.n1 VTAIL.n0 42.6192
R157 VTAIL.n5 VTAIL.n4 42.6192
R158 VTAIL.n15 VTAIL.n14 26.7807
R159 VTAIL.n7 VTAIL.n6 26.7807
R160 VTAIL.n9 VTAIL.n7 3.13843
R161 VTAIL.n10 VTAIL.n9 3.13843
R162 VTAIL.n13 VTAIL.n11 3.13843
R163 VTAIL.n14 VTAIL.n13 3.13843
R164 VTAIL.n6 VTAIL.n5 3.13843
R165 VTAIL.n5 VTAIL.n3 3.13843
R166 VTAIL.n2 VTAIL.n1 3.13843
R167 VTAIL VTAIL.n15 3.08024
R168 VTAIL.n0 VTAIL.t6 1.51426
R169 VTAIL.n0 VTAIL.t5 1.51426
R170 VTAIL.n4 VTAIL.t9 1.51426
R171 VTAIL.n4 VTAIL.t11 1.51426
R172 VTAIL.n12 VTAIL.t10 1.51426
R173 VTAIL.n12 VTAIL.t14 1.51426
R174 VTAIL.n8 VTAIL.t2 1.51426
R175 VTAIL.n8 VTAIL.t15 1.51426
R176 VTAIL.n11 VTAIL.n10 0.470328
R177 VTAIL.n3 VTAIL.n2 0.470328
R178 VTAIL VTAIL.n1 0.0586897
R179 B.n1000 B.n999 585
R180 B.n1001 B.n1000 585
R181 B.n363 B.n162 585
R182 B.n362 B.n361 585
R183 B.n360 B.n359 585
R184 B.n358 B.n357 585
R185 B.n356 B.n355 585
R186 B.n354 B.n353 585
R187 B.n352 B.n351 585
R188 B.n350 B.n349 585
R189 B.n348 B.n347 585
R190 B.n346 B.n345 585
R191 B.n344 B.n343 585
R192 B.n342 B.n341 585
R193 B.n340 B.n339 585
R194 B.n338 B.n337 585
R195 B.n336 B.n335 585
R196 B.n334 B.n333 585
R197 B.n332 B.n331 585
R198 B.n330 B.n329 585
R199 B.n328 B.n327 585
R200 B.n326 B.n325 585
R201 B.n324 B.n323 585
R202 B.n322 B.n321 585
R203 B.n320 B.n319 585
R204 B.n318 B.n317 585
R205 B.n316 B.n315 585
R206 B.n314 B.n313 585
R207 B.n312 B.n311 585
R208 B.n310 B.n309 585
R209 B.n308 B.n307 585
R210 B.n306 B.n305 585
R211 B.n304 B.n303 585
R212 B.n302 B.n301 585
R213 B.n300 B.n299 585
R214 B.n298 B.n297 585
R215 B.n296 B.n295 585
R216 B.n294 B.n293 585
R217 B.n292 B.n291 585
R218 B.n290 B.n289 585
R219 B.n288 B.n287 585
R220 B.n286 B.n285 585
R221 B.n284 B.n283 585
R222 B.n282 B.n281 585
R223 B.n280 B.n279 585
R224 B.n278 B.n277 585
R225 B.n276 B.n275 585
R226 B.n274 B.n273 585
R227 B.n272 B.n271 585
R228 B.n270 B.n269 585
R229 B.n268 B.n267 585
R230 B.n266 B.n265 585
R231 B.n264 B.n263 585
R232 B.n262 B.n261 585
R233 B.n260 B.n259 585
R234 B.n257 B.n256 585
R235 B.n255 B.n254 585
R236 B.n253 B.n252 585
R237 B.n251 B.n250 585
R238 B.n249 B.n248 585
R239 B.n247 B.n246 585
R240 B.n245 B.n244 585
R241 B.n243 B.n242 585
R242 B.n241 B.n240 585
R243 B.n239 B.n238 585
R244 B.n237 B.n236 585
R245 B.n235 B.n234 585
R246 B.n233 B.n232 585
R247 B.n231 B.n230 585
R248 B.n229 B.n228 585
R249 B.n227 B.n226 585
R250 B.n225 B.n224 585
R251 B.n223 B.n222 585
R252 B.n221 B.n220 585
R253 B.n219 B.n218 585
R254 B.n217 B.n216 585
R255 B.n215 B.n214 585
R256 B.n213 B.n212 585
R257 B.n211 B.n210 585
R258 B.n209 B.n208 585
R259 B.n207 B.n206 585
R260 B.n205 B.n204 585
R261 B.n203 B.n202 585
R262 B.n201 B.n200 585
R263 B.n199 B.n198 585
R264 B.n197 B.n196 585
R265 B.n195 B.n194 585
R266 B.n193 B.n192 585
R267 B.n191 B.n190 585
R268 B.n189 B.n188 585
R269 B.n187 B.n186 585
R270 B.n185 B.n184 585
R271 B.n183 B.n182 585
R272 B.n181 B.n180 585
R273 B.n179 B.n178 585
R274 B.n177 B.n176 585
R275 B.n175 B.n174 585
R276 B.n173 B.n172 585
R277 B.n171 B.n170 585
R278 B.n169 B.n168 585
R279 B.n998 B.n112 585
R280 B.n1002 B.n112 585
R281 B.n997 B.n111 585
R282 B.n1003 B.n111 585
R283 B.n996 B.n995 585
R284 B.n995 B.n107 585
R285 B.n994 B.n106 585
R286 B.n1009 B.n106 585
R287 B.n993 B.n105 585
R288 B.n1010 B.n105 585
R289 B.n992 B.n104 585
R290 B.n1011 B.n104 585
R291 B.n991 B.n990 585
R292 B.n990 B.n100 585
R293 B.n989 B.n99 585
R294 B.n1017 B.n99 585
R295 B.n988 B.n98 585
R296 B.n1018 B.n98 585
R297 B.n987 B.n97 585
R298 B.n1019 B.n97 585
R299 B.n986 B.n985 585
R300 B.n985 B.n93 585
R301 B.n984 B.n92 585
R302 B.n1025 B.n92 585
R303 B.n983 B.n91 585
R304 B.n1026 B.n91 585
R305 B.n982 B.n90 585
R306 B.n1027 B.n90 585
R307 B.n981 B.n980 585
R308 B.n980 B.n86 585
R309 B.n979 B.n85 585
R310 B.n1033 B.n85 585
R311 B.n978 B.n84 585
R312 B.n1034 B.n84 585
R313 B.n977 B.n83 585
R314 B.n1035 B.n83 585
R315 B.n976 B.n975 585
R316 B.n975 B.n79 585
R317 B.n974 B.n78 585
R318 B.n1041 B.n78 585
R319 B.n973 B.n77 585
R320 B.n1042 B.n77 585
R321 B.n972 B.n76 585
R322 B.n1043 B.n76 585
R323 B.n971 B.n970 585
R324 B.n970 B.n75 585
R325 B.n969 B.n71 585
R326 B.n1049 B.n71 585
R327 B.n968 B.n70 585
R328 B.n1050 B.n70 585
R329 B.n967 B.n69 585
R330 B.n1051 B.n69 585
R331 B.n966 B.n965 585
R332 B.n965 B.n65 585
R333 B.n964 B.n64 585
R334 B.n1057 B.n64 585
R335 B.n963 B.n63 585
R336 B.n1058 B.n63 585
R337 B.n962 B.n62 585
R338 B.n1059 B.n62 585
R339 B.n961 B.n960 585
R340 B.n960 B.n58 585
R341 B.n959 B.n57 585
R342 B.n1065 B.n57 585
R343 B.n958 B.n56 585
R344 B.n1066 B.n56 585
R345 B.n957 B.n55 585
R346 B.n1067 B.n55 585
R347 B.n956 B.n955 585
R348 B.n955 B.n51 585
R349 B.n954 B.n50 585
R350 B.n1073 B.n50 585
R351 B.n953 B.n49 585
R352 B.n1074 B.n49 585
R353 B.n952 B.n48 585
R354 B.n1075 B.n48 585
R355 B.n951 B.n950 585
R356 B.n950 B.n44 585
R357 B.n949 B.n43 585
R358 B.n1081 B.n43 585
R359 B.n948 B.n42 585
R360 B.n1082 B.n42 585
R361 B.n947 B.n41 585
R362 B.n1083 B.n41 585
R363 B.n946 B.n945 585
R364 B.n945 B.n37 585
R365 B.n944 B.n36 585
R366 B.n1089 B.n36 585
R367 B.n943 B.n35 585
R368 B.n1090 B.n35 585
R369 B.n942 B.n34 585
R370 B.n1091 B.n34 585
R371 B.n941 B.n940 585
R372 B.n940 B.n30 585
R373 B.n939 B.n29 585
R374 B.n1097 B.n29 585
R375 B.n938 B.n28 585
R376 B.n1098 B.n28 585
R377 B.n937 B.n27 585
R378 B.n1099 B.n27 585
R379 B.n936 B.n935 585
R380 B.n935 B.n23 585
R381 B.n934 B.n22 585
R382 B.n1105 B.n22 585
R383 B.n933 B.n21 585
R384 B.n1106 B.n21 585
R385 B.n932 B.n20 585
R386 B.n1107 B.n20 585
R387 B.n931 B.n930 585
R388 B.n930 B.n19 585
R389 B.n929 B.n15 585
R390 B.n1113 B.n15 585
R391 B.n928 B.n14 585
R392 B.n1114 B.n14 585
R393 B.n927 B.n13 585
R394 B.n1115 B.n13 585
R395 B.n926 B.n925 585
R396 B.n925 B.n12 585
R397 B.n924 B.n923 585
R398 B.n924 B.n8 585
R399 B.n922 B.n7 585
R400 B.n1122 B.n7 585
R401 B.n921 B.n6 585
R402 B.n1123 B.n6 585
R403 B.n920 B.n5 585
R404 B.n1124 B.n5 585
R405 B.n919 B.n918 585
R406 B.n918 B.n4 585
R407 B.n917 B.n364 585
R408 B.n917 B.n916 585
R409 B.n907 B.n365 585
R410 B.n366 B.n365 585
R411 B.n909 B.n908 585
R412 B.n910 B.n909 585
R413 B.n906 B.n371 585
R414 B.n371 B.n370 585
R415 B.n905 B.n904 585
R416 B.n904 B.n903 585
R417 B.n373 B.n372 585
R418 B.n896 B.n373 585
R419 B.n895 B.n894 585
R420 B.n897 B.n895 585
R421 B.n893 B.n378 585
R422 B.n378 B.n377 585
R423 B.n892 B.n891 585
R424 B.n891 B.n890 585
R425 B.n380 B.n379 585
R426 B.n381 B.n380 585
R427 B.n883 B.n882 585
R428 B.n884 B.n883 585
R429 B.n881 B.n386 585
R430 B.n386 B.n385 585
R431 B.n880 B.n879 585
R432 B.n879 B.n878 585
R433 B.n388 B.n387 585
R434 B.n389 B.n388 585
R435 B.n871 B.n870 585
R436 B.n872 B.n871 585
R437 B.n869 B.n394 585
R438 B.n394 B.n393 585
R439 B.n868 B.n867 585
R440 B.n867 B.n866 585
R441 B.n396 B.n395 585
R442 B.n397 B.n396 585
R443 B.n859 B.n858 585
R444 B.n860 B.n859 585
R445 B.n857 B.n402 585
R446 B.n402 B.n401 585
R447 B.n856 B.n855 585
R448 B.n855 B.n854 585
R449 B.n404 B.n403 585
R450 B.n405 B.n404 585
R451 B.n847 B.n846 585
R452 B.n848 B.n847 585
R453 B.n845 B.n410 585
R454 B.n410 B.n409 585
R455 B.n844 B.n843 585
R456 B.n843 B.n842 585
R457 B.n412 B.n411 585
R458 B.n413 B.n412 585
R459 B.n835 B.n834 585
R460 B.n836 B.n835 585
R461 B.n833 B.n418 585
R462 B.n418 B.n417 585
R463 B.n832 B.n831 585
R464 B.n831 B.n830 585
R465 B.n420 B.n419 585
R466 B.n421 B.n420 585
R467 B.n823 B.n822 585
R468 B.n824 B.n823 585
R469 B.n821 B.n426 585
R470 B.n426 B.n425 585
R471 B.n820 B.n819 585
R472 B.n819 B.n818 585
R473 B.n428 B.n427 585
R474 B.n429 B.n428 585
R475 B.n811 B.n810 585
R476 B.n812 B.n811 585
R477 B.n809 B.n434 585
R478 B.n434 B.n433 585
R479 B.n808 B.n807 585
R480 B.n807 B.n806 585
R481 B.n436 B.n435 585
R482 B.n799 B.n436 585
R483 B.n798 B.n797 585
R484 B.n800 B.n798 585
R485 B.n796 B.n441 585
R486 B.n441 B.n440 585
R487 B.n795 B.n794 585
R488 B.n794 B.n793 585
R489 B.n443 B.n442 585
R490 B.n444 B.n443 585
R491 B.n786 B.n785 585
R492 B.n787 B.n786 585
R493 B.n784 B.n449 585
R494 B.n449 B.n448 585
R495 B.n783 B.n782 585
R496 B.n782 B.n781 585
R497 B.n451 B.n450 585
R498 B.n452 B.n451 585
R499 B.n774 B.n773 585
R500 B.n775 B.n774 585
R501 B.n772 B.n457 585
R502 B.n457 B.n456 585
R503 B.n771 B.n770 585
R504 B.n770 B.n769 585
R505 B.n459 B.n458 585
R506 B.n460 B.n459 585
R507 B.n762 B.n761 585
R508 B.n763 B.n762 585
R509 B.n760 B.n464 585
R510 B.n468 B.n464 585
R511 B.n759 B.n758 585
R512 B.n758 B.n757 585
R513 B.n466 B.n465 585
R514 B.n467 B.n466 585
R515 B.n750 B.n749 585
R516 B.n751 B.n750 585
R517 B.n748 B.n473 585
R518 B.n473 B.n472 585
R519 B.n747 B.n746 585
R520 B.n746 B.n745 585
R521 B.n475 B.n474 585
R522 B.n476 B.n475 585
R523 B.n738 B.n737 585
R524 B.n739 B.n738 585
R525 B.n736 B.n481 585
R526 B.n481 B.n480 585
R527 B.n730 B.n729 585
R528 B.n728 B.n532 585
R529 B.n727 B.n531 585
R530 B.n732 B.n531 585
R531 B.n726 B.n725 585
R532 B.n724 B.n723 585
R533 B.n722 B.n721 585
R534 B.n720 B.n719 585
R535 B.n718 B.n717 585
R536 B.n716 B.n715 585
R537 B.n714 B.n713 585
R538 B.n712 B.n711 585
R539 B.n710 B.n709 585
R540 B.n708 B.n707 585
R541 B.n706 B.n705 585
R542 B.n704 B.n703 585
R543 B.n702 B.n701 585
R544 B.n700 B.n699 585
R545 B.n698 B.n697 585
R546 B.n696 B.n695 585
R547 B.n694 B.n693 585
R548 B.n692 B.n691 585
R549 B.n690 B.n689 585
R550 B.n688 B.n687 585
R551 B.n686 B.n685 585
R552 B.n684 B.n683 585
R553 B.n682 B.n681 585
R554 B.n680 B.n679 585
R555 B.n678 B.n677 585
R556 B.n676 B.n675 585
R557 B.n674 B.n673 585
R558 B.n672 B.n671 585
R559 B.n670 B.n669 585
R560 B.n668 B.n667 585
R561 B.n666 B.n665 585
R562 B.n664 B.n663 585
R563 B.n662 B.n661 585
R564 B.n660 B.n659 585
R565 B.n658 B.n657 585
R566 B.n656 B.n655 585
R567 B.n654 B.n653 585
R568 B.n652 B.n651 585
R569 B.n650 B.n649 585
R570 B.n648 B.n647 585
R571 B.n646 B.n645 585
R572 B.n644 B.n643 585
R573 B.n642 B.n641 585
R574 B.n640 B.n639 585
R575 B.n638 B.n637 585
R576 B.n636 B.n635 585
R577 B.n634 B.n633 585
R578 B.n632 B.n631 585
R579 B.n630 B.n629 585
R580 B.n628 B.n627 585
R581 B.n626 B.n625 585
R582 B.n623 B.n622 585
R583 B.n621 B.n620 585
R584 B.n619 B.n618 585
R585 B.n617 B.n616 585
R586 B.n615 B.n614 585
R587 B.n613 B.n612 585
R588 B.n611 B.n610 585
R589 B.n609 B.n608 585
R590 B.n607 B.n606 585
R591 B.n605 B.n604 585
R592 B.n603 B.n602 585
R593 B.n601 B.n600 585
R594 B.n599 B.n598 585
R595 B.n597 B.n596 585
R596 B.n595 B.n594 585
R597 B.n593 B.n592 585
R598 B.n591 B.n590 585
R599 B.n589 B.n588 585
R600 B.n587 B.n586 585
R601 B.n585 B.n584 585
R602 B.n583 B.n582 585
R603 B.n581 B.n580 585
R604 B.n579 B.n578 585
R605 B.n577 B.n576 585
R606 B.n575 B.n574 585
R607 B.n573 B.n572 585
R608 B.n571 B.n570 585
R609 B.n569 B.n568 585
R610 B.n567 B.n566 585
R611 B.n565 B.n564 585
R612 B.n563 B.n562 585
R613 B.n561 B.n560 585
R614 B.n559 B.n558 585
R615 B.n557 B.n556 585
R616 B.n555 B.n554 585
R617 B.n553 B.n552 585
R618 B.n551 B.n550 585
R619 B.n549 B.n548 585
R620 B.n547 B.n546 585
R621 B.n545 B.n544 585
R622 B.n543 B.n542 585
R623 B.n541 B.n540 585
R624 B.n539 B.n538 585
R625 B.n483 B.n482 585
R626 B.n735 B.n734 585
R627 B.n479 B.n478 585
R628 B.n480 B.n479 585
R629 B.n741 B.n740 585
R630 B.n740 B.n739 585
R631 B.n742 B.n477 585
R632 B.n477 B.n476 585
R633 B.n744 B.n743 585
R634 B.n745 B.n744 585
R635 B.n471 B.n470 585
R636 B.n472 B.n471 585
R637 B.n753 B.n752 585
R638 B.n752 B.n751 585
R639 B.n754 B.n469 585
R640 B.n469 B.n467 585
R641 B.n756 B.n755 585
R642 B.n757 B.n756 585
R643 B.n463 B.n462 585
R644 B.n468 B.n463 585
R645 B.n765 B.n764 585
R646 B.n764 B.n763 585
R647 B.n766 B.n461 585
R648 B.n461 B.n460 585
R649 B.n768 B.n767 585
R650 B.n769 B.n768 585
R651 B.n455 B.n454 585
R652 B.n456 B.n455 585
R653 B.n777 B.n776 585
R654 B.n776 B.n775 585
R655 B.n778 B.n453 585
R656 B.n453 B.n452 585
R657 B.n780 B.n779 585
R658 B.n781 B.n780 585
R659 B.n447 B.n446 585
R660 B.n448 B.n447 585
R661 B.n789 B.n788 585
R662 B.n788 B.n787 585
R663 B.n790 B.n445 585
R664 B.n445 B.n444 585
R665 B.n792 B.n791 585
R666 B.n793 B.n792 585
R667 B.n439 B.n438 585
R668 B.n440 B.n439 585
R669 B.n802 B.n801 585
R670 B.n801 B.n800 585
R671 B.n803 B.n437 585
R672 B.n799 B.n437 585
R673 B.n805 B.n804 585
R674 B.n806 B.n805 585
R675 B.n432 B.n431 585
R676 B.n433 B.n432 585
R677 B.n814 B.n813 585
R678 B.n813 B.n812 585
R679 B.n815 B.n430 585
R680 B.n430 B.n429 585
R681 B.n817 B.n816 585
R682 B.n818 B.n817 585
R683 B.n424 B.n423 585
R684 B.n425 B.n424 585
R685 B.n826 B.n825 585
R686 B.n825 B.n824 585
R687 B.n827 B.n422 585
R688 B.n422 B.n421 585
R689 B.n829 B.n828 585
R690 B.n830 B.n829 585
R691 B.n416 B.n415 585
R692 B.n417 B.n416 585
R693 B.n838 B.n837 585
R694 B.n837 B.n836 585
R695 B.n839 B.n414 585
R696 B.n414 B.n413 585
R697 B.n841 B.n840 585
R698 B.n842 B.n841 585
R699 B.n408 B.n407 585
R700 B.n409 B.n408 585
R701 B.n850 B.n849 585
R702 B.n849 B.n848 585
R703 B.n851 B.n406 585
R704 B.n406 B.n405 585
R705 B.n853 B.n852 585
R706 B.n854 B.n853 585
R707 B.n400 B.n399 585
R708 B.n401 B.n400 585
R709 B.n862 B.n861 585
R710 B.n861 B.n860 585
R711 B.n863 B.n398 585
R712 B.n398 B.n397 585
R713 B.n865 B.n864 585
R714 B.n866 B.n865 585
R715 B.n392 B.n391 585
R716 B.n393 B.n392 585
R717 B.n874 B.n873 585
R718 B.n873 B.n872 585
R719 B.n875 B.n390 585
R720 B.n390 B.n389 585
R721 B.n877 B.n876 585
R722 B.n878 B.n877 585
R723 B.n384 B.n383 585
R724 B.n385 B.n384 585
R725 B.n886 B.n885 585
R726 B.n885 B.n884 585
R727 B.n887 B.n382 585
R728 B.n382 B.n381 585
R729 B.n889 B.n888 585
R730 B.n890 B.n889 585
R731 B.n376 B.n375 585
R732 B.n377 B.n376 585
R733 B.n899 B.n898 585
R734 B.n898 B.n897 585
R735 B.n900 B.n374 585
R736 B.n896 B.n374 585
R737 B.n902 B.n901 585
R738 B.n903 B.n902 585
R739 B.n369 B.n368 585
R740 B.n370 B.n369 585
R741 B.n912 B.n911 585
R742 B.n911 B.n910 585
R743 B.n913 B.n367 585
R744 B.n367 B.n366 585
R745 B.n915 B.n914 585
R746 B.n916 B.n915 585
R747 B.n3 B.n0 585
R748 B.n4 B.n3 585
R749 B.n1121 B.n1 585
R750 B.n1122 B.n1121 585
R751 B.n1120 B.n1119 585
R752 B.n1120 B.n8 585
R753 B.n1118 B.n9 585
R754 B.n12 B.n9 585
R755 B.n1117 B.n1116 585
R756 B.n1116 B.n1115 585
R757 B.n11 B.n10 585
R758 B.n1114 B.n11 585
R759 B.n1112 B.n1111 585
R760 B.n1113 B.n1112 585
R761 B.n1110 B.n16 585
R762 B.n19 B.n16 585
R763 B.n1109 B.n1108 585
R764 B.n1108 B.n1107 585
R765 B.n18 B.n17 585
R766 B.n1106 B.n18 585
R767 B.n1104 B.n1103 585
R768 B.n1105 B.n1104 585
R769 B.n1102 B.n24 585
R770 B.n24 B.n23 585
R771 B.n1101 B.n1100 585
R772 B.n1100 B.n1099 585
R773 B.n26 B.n25 585
R774 B.n1098 B.n26 585
R775 B.n1096 B.n1095 585
R776 B.n1097 B.n1096 585
R777 B.n1094 B.n31 585
R778 B.n31 B.n30 585
R779 B.n1093 B.n1092 585
R780 B.n1092 B.n1091 585
R781 B.n33 B.n32 585
R782 B.n1090 B.n33 585
R783 B.n1088 B.n1087 585
R784 B.n1089 B.n1088 585
R785 B.n1086 B.n38 585
R786 B.n38 B.n37 585
R787 B.n1085 B.n1084 585
R788 B.n1084 B.n1083 585
R789 B.n40 B.n39 585
R790 B.n1082 B.n40 585
R791 B.n1080 B.n1079 585
R792 B.n1081 B.n1080 585
R793 B.n1078 B.n45 585
R794 B.n45 B.n44 585
R795 B.n1077 B.n1076 585
R796 B.n1076 B.n1075 585
R797 B.n47 B.n46 585
R798 B.n1074 B.n47 585
R799 B.n1072 B.n1071 585
R800 B.n1073 B.n1072 585
R801 B.n1070 B.n52 585
R802 B.n52 B.n51 585
R803 B.n1069 B.n1068 585
R804 B.n1068 B.n1067 585
R805 B.n54 B.n53 585
R806 B.n1066 B.n54 585
R807 B.n1064 B.n1063 585
R808 B.n1065 B.n1064 585
R809 B.n1062 B.n59 585
R810 B.n59 B.n58 585
R811 B.n1061 B.n1060 585
R812 B.n1060 B.n1059 585
R813 B.n61 B.n60 585
R814 B.n1058 B.n61 585
R815 B.n1056 B.n1055 585
R816 B.n1057 B.n1056 585
R817 B.n1054 B.n66 585
R818 B.n66 B.n65 585
R819 B.n1053 B.n1052 585
R820 B.n1052 B.n1051 585
R821 B.n68 B.n67 585
R822 B.n1050 B.n68 585
R823 B.n1048 B.n1047 585
R824 B.n1049 B.n1048 585
R825 B.n1046 B.n72 585
R826 B.n75 B.n72 585
R827 B.n1045 B.n1044 585
R828 B.n1044 B.n1043 585
R829 B.n74 B.n73 585
R830 B.n1042 B.n74 585
R831 B.n1040 B.n1039 585
R832 B.n1041 B.n1040 585
R833 B.n1038 B.n80 585
R834 B.n80 B.n79 585
R835 B.n1037 B.n1036 585
R836 B.n1036 B.n1035 585
R837 B.n82 B.n81 585
R838 B.n1034 B.n82 585
R839 B.n1032 B.n1031 585
R840 B.n1033 B.n1032 585
R841 B.n1030 B.n87 585
R842 B.n87 B.n86 585
R843 B.n1029 B.n1028 585
R844 B.n1028 B.n1027 585
R845 B.n89 B.n88 585
R846 B.n1026 B.n89 585
R847 B.n1024 B.n1023 585
R848 B.n1025 B.n1024 585
R849 B.n1022 B.n94 585
R850 B.n94 B.n93 585
R851 B.n1021 B.n1020 585
R852 B.n1020 B.n1019 585
R853 B.n96 B.n95 585
R854 B.n1018 B.n96 585
R855 B.n1016 B.n1015 585
R856 B.n1017 B.n1016 585
R857 B.n1014 B.n101 585
R858 B.n101 B.n100 585
R859 B.n1013 B.n1012 585
R860 B.n1012 B.n1011 585
R861 B.n103 B.n102 585
R862 B.n1010 B.n103 585
R863 B.n1008 B.n1007 585
R864 B.n1009 B.n1008 585
R865 B.n1006 B.n108 585
R866 B.n108 B.n107 585
R867 B.n1005 B.n1004 585
R868 B.n1004 B.n1003 585
R869 B.n110 B.n109 585
R870 B.n1002 B.n110 585
R871 B.n1125 B.n1124 585
R872 B.n1123 B.n2 585
R873 B.n168 B.n110 535.745
R874 B.n1000 B.n112 535.745
R875 B.n734 B.n481 535.745
R876 B.n730 B.n479 535.745
R877 B.n166 B.t16 304.151
R878 B.n163 B.t8 304.151
R879 B.n536 B.t19 304.151
R880 B.n533 B.t12 304.151
R881 B.n1001 B.n161 256.663
R882 B.n1001 B.n160 256.663
R883 B.n1001 B.n159 256.663
R884 B.n1001 B.n158 256.663
R885 B.n1001 B.n157 256.663
R886 B.n1001 B.n156 256.663
R887 B.n1001 B.n155 256.663
R888 B.n1001 B.n154 256.663
R889 B.n1001 B.n153 256.663
R890 B.n1001 B.n152 256.663
R891 B.n1001 B.n151 256.663
R892 B.n1001 B.n150 256.663
R893 B.n1001 B.n149 256.663
R894 B.n1001 B.n148 256.663
R895 B.n1001 B.n147 256.663
R896 B.n1001 B.n146 256.663
R897 B.n1001 B.n145 256.663
R898 B.n1001 B.n144 256.663
R899 B.n1001 B.n143 256.663
R900 B.n1001 B.n142 256.663
R901 B.n1001 B.n141 256.663
R902 B.n1001 B.n140 256.663
R903 B.n1001 B.n139 256.663
R904 B.n1001 B.n138 256.663
R905 B.n1001 B.n137 256.663
R906 B.n1001 B.n136 256.663
R907 B.n1001 B.n135 256.663
R908 B.n1001 B.n134 256.663
R909 B.n1001 B.n133 256.663
R910 B.n1001 B.n132 256.663
R911 B.n1001 B.n131 256.663
R912 B.n1001 B.n130 256.663
R913 B.n1001 B.n129 256.663
R914 B.n1001 B.n128 256.663
R915 B.n1001 B.n127 256.663
R916 B.n1001 B.n126 256.663
R917 B.n1001 B.n125 256.663
R918 B.n1001 B.n124 256.663
R919 B.n1001 B.n123 256.663
R920 B.n1001 B.n122 256.663
R921 B.n1001 B.n121 256.663
R922 B.n1001 B.n120 256.663
R923 B.n1001 B.n119 256.663
R924 B.n1001 B.n118 256.663
R925 B.n1001 B.n117 256.663
R926 B.n1001 B.n116 256.663
R927 B.n1001 B.n115 256.663
R928 B.n1001 B.n114 256.663
R929 B.n1001 B.n113 256.663
R930 B.n732 B.n731 256.663
R931 B.n732 B.n484 256.663
R932 B.n732 B.n485 256.663
R933 B.n732 B.n486 256.663
R934 B.n732 B.n487 256.663
R935 B.n732 B.n488 256.663
R936 B.n732 B.n489 256.663
R937 B.n732 B.n490 256.663
R938 B.n732 B.n491 256.663
R939 B.n732 B.n492 256.663
R940 B.n732 B.n493 256.663
R941 B.n732 B.n494 256.663
R942 B.n732 B.n495 256.663
R943 B.n732 B.n496 256.663
R944 B.n732 B.n497 256.663
R945 B.n732 B.n498 256.663
R946 B.n732 B.n499 256.663
R947 B.n732 B.n500 256.663
R948 B.n732 B.n501 256.663
R949 B.n732 B.n502 256.663
R950 B.n732 B.n503 256.663
R951 B.n732 B.n504 256.663
R952 B.n732 B.n505 256.663
R953 B.n732 B.n506 256.663
R954 B.n732 B.n507 256.663
R955 B.n732 B.n508 256.663
R956 B.n732 B.n509 256.663
R957 B.n732 B.n510 256.663
R958 B.n732 B.n511 256.663
R959 B.n732 B.n512 256.663
R960 B.n732 B.n513 256.663
R961 B.n732 B.n514 256.663
R962 B.n732 B.n515 256.663
R963 B.n732 B.n516 256.663
R964 B.n732 B.n517 256.663
R965 B.n732 B.n518 256.663
R966 B.n732 B.n519 256.663
R967 B.n732 B.n520 256.663
R968 B.n732 B.n521 256.663
R969 B.n732 B.n522 256.663
R970 B.n732 B.n523 256.663
R971 B.n732 B.n524 256.663
R972 B.n732 B.n525 256.663
R973 B.n732 B.n526 256.663
R974 B.n732 B.n527 256.663
R975 B.n732 B.n528 256.663
R976 B.n732 B.n529 256.663
R977 B.n732 B.n530 256.663
R978 B.n733 B.n732 256.663
R979 B.n1127 B.n1126 256.663
R980 B.n172 B.n171 163.367
R981 B.n176 B.n175 163.367
R982 B.n180 B.n179 163.367
R983 B.n184 B.n183 163.367
R984 B.n188 B.n187 163.367
R985 B.n192 B.n191 163.367
R986 B.n196 B.n195 163.367
R987 B.n200 B.n199 163.367
R988 B.n204 B.n203 163.367
R989 B.n208 B.n207 163.367
R990 B.n212 B.n211 163.367
R991 B.n216 B.n215 163.367
R992 B.n220 B.n219 163.367
R993 B.n224 B.n223 163.367
R994 B.n228 B.n227 163.367
R995 B.n232 B.n231 163.367
R996 B.n236 B.n235 163.367
R997 B.n240 B.n239 163.367
R998 B.n244 B.n243 163.367
R999 B.n248 B.n247 163.367
R1000 B.n252 B.n251 163.367
R1001 B.n256 B.n255 163.367
R1002 B.n261 B.n260 163.367
R1003 B.n265 B.n264 163.367
R1004 B.n269 B.n268 163.367
R1005 B.n273 B.n272 163.367
R1006 B.n277 B.n276 163.367
R1007 B.n281 B.n280 163.367
R1008 B.n285 B.n284 163.367
R1009 B.n289 B.n288 163.367
R1010 B.n293 B.n292 163.367
R1011 B.n297 B.n296 163.367
R1012 B.n301 B.n300 163.367
R1013 B.n305 B.n304 163.367
R1014 B.n309 B.n308 163.367
R1015 B.n313 B.n312 163.367
R1016 B.n317 B.n316 163.367
R1017 B.n321 B.n320 163.367
R1018 B.n325 B.n324 163.367
R1019 B.n329 B.n328 163.367
R1020 B.n333 B.n332 163.367
R1021 B.n337 B.n336 163.367
R1022 B.n341 B.n340 163.367
R1023 B.n345 B.n344 163.367
R1024 B.n349 B.n348 163.367
R1025 B.n353 B.n352 163.367
R1026 B.n357 B.n356 163.367
R1027 B.n361 B.n360 163.367
R1028 B.n1000 B.n162 163.367
R1029 B.n738 B.n481 163.367
R1030 B.n738 B.n475 163.367
R1031 B.n746 B.n475 163.367
R1032 B.n746 B.n473 163.367
R1033 B.n750 B.n473 163.367
R1034 B.n750 B.n466 163.367
R1035 B.n758 B.n466 163.367
R1036 B.n758 B.n464 163.367
R1037 B.n762 B.n464 163.367
R1038 B.n762 B.n459 163.367
R1039 B.n770 B.n459 163.367
R1040 B.n770 B.n457 163.367
R1041 B.n774 B.n457 163.367
R1042 B.n774 B.n451 163.367
R1043 B.n782 B.n451 163.367
R1044 B.n782 B.n449 163.367
R1045 B.n786 B.n449 163.367
R1046 B.n786 B.n443 163.367
R1047 B.n794 B.n443 163.367
R1048 B.n794 B.n441 163.367
R1049 B.n798 B.n441 163.367
R1050 B.n798 B.n436 163.367
R1051 B.n807 B.n436 163.367
R1052 B.n807 B.n434 163.367
R1053 B.n811 B.n434 163.367
R1054 B.n811 B.n428 163.367
R1055 B.n819 B.n428 163.367
R1056 B.n819 B.n426 163.367
R1057 B.n823 B.n426 163.367
R1058 B.n823 B.n420 163.367
R1059 B.n831 B.n420 163.367
R1060 B.n831 B.n418 163.367
R1061 B.n835 B.n418 163.367
R1062 B.n835 B.n412 163.367
R1063 B.n843 B.n412 163.367
R1064 B.n843 B.n410 163.367
R1065 B.n847 B.n410 163.367
R1066 B.n847 B.n404 163.367
R1067 B.n855 B.n404 163.367
R1068 B.n855 B.n402 163.367
R1069 B.n859 B.n402 163.367
R1070 B.n859 B.n396 163.367
R1071 B.n867 B.n396 163.367
R1072 B.n867 B.n394 163.367
R1073 B.n871 B.n394 163.367
R1074 B.n871 B.n388 163.367
R1075 B.n879 B.n388 163.367
R1076 B.n879 B.n386 163.367
R1077 B.n883 B.n386 163.367
R1078 B.n883 B.n380 163.367
R1079 B.n891 B.n380 163.367
R1080 B.n891 B.n378 163.367
R1081 B.n895 B.n378 163.367
R1082 B.n895 B.n373 163.367
R1083 B.n904 B.n373 163.367
R1084 B.n904 B.n371 163.367
R1085 B.n909 B.n371 163.367
R1086 B.n909 B.n365 163.367
R1087 B.n917 B.n365 163.367
R1088 B.n918 B.n917 163.367
R1089 B.n918 B.n5 163.367
R1090 B.n6 B.n5 163.367
R1091 B.n7 B.n6 163.367
R1092 B.n924 B.n7 163.367
R1093 B.n925 B.n924 163.367
R1094 B.n925 B.n13 163.367
R1095 B.n14 B.n13 163.367
R1096 B.n15 B.n14 163.367
R1097 B.n930 B.n15 163.367
R1098 B.n930 B.n20 163.367
R1099 B.n21 B.n20 163.367
R1100 B.n22 B.n21 163.367
R1101 B.n935 B.n22 163.367
R1102 B.n935 B.n27 163.367
R1103 B.n28 B.n27 163.367
R1104 B.n29 B.n28 163.367
R1105 B.n940 B.n29 163.367
R1106 B.n940 B.n34 163.367
R1107 B.n35 B.n34 163.367
R1108 B.n36 B.n35 163.367
R1109 B.n945 B.n36 163.367
R1110 B.n945 B.n41 163.367
R1111 B.n42 B.n41 163.367
R1112 B.n43 B.n42 163.367
R1113 B.n950 B.n43 163.367
R1114 B.n950 B.n48 163.367
R1115 B.n49 B.n48 163.367
R1116 B.n50 B.n49 163.367
R1117 B.n955 B.n50 163.367
R1118 B.n955 B.n55 163.367
R1119 B.n56 B.n55 163.367
R1120 B.n57 B.n56 163.367
R1121 B.n960 B.n57 163.367
R1122 B.n960 B.n62 163.367
R1123 B.n63 B.n62 163.367
R1124 B.n64 B.n63 163.367
R1125 B.n965 B.n64 163.367
R1126 B.n965 B.n69 163.367
R1127 B.n70 B.n69 163.367
R1128 B.n71 B.n70 163.367
R1129 B.n970 B.n71 163.367
R1130 B.n970 B.n76 163.367
R1131 B.n77 B.n76 163.367
R1132 B.n78 B.n77 163.367
R1133 B.n975 B.n78 163.367
R1134 B.n975 B.n83 163.367
R1135 B.n84 B.n83 163.367
R1136 B.n85 B.n84 163.367
R1137 B.n980 B.n85 163.367
R1138 B.n980 B.n90 163.367
R1139 B.n91 B.n90 163.367
R1140 B.n92 B.n91 163.367
R1141 B.n985 B.n92 163.367
R1142 B.n985 B.n97 163.367
R1143 B.n98 B.n97 163.367
R1144 B.n99 B.n98 163.367
R1145 B.n990 B.n99 163.367
R1146 B.n990 B.n104 163.367
R1147 B.n105 B.n104 163.367
R1148 B.n106 B.n105 163.367
R1149 B.n995 B.n106 163.367
R1150 B.n995 B.n111 163.367
R1151 B.n112 B.n111 163.367
R1152 B.n532 B.n531 163.367
R1153 B.n725 B.n531 163.367
R1154 B.n723 B.n722 163.367
R1155 B.n719 B.n718 163.367
R1156 B.n715 B.n714 163.367
R1157 B.n711 B.n710 163.367
R1158 B.n707 B.n706 163.367
R1159 B.n703 B.n702 163.367
R1160 B.n699 B.n698 163.367
R1161 B.n695 B.n694 163.367
R1162 B.n691 B.n690 163.367
R1163 B.n687 B.n686 163.367
R1164 B.n683 B.n682 163.367
R1165 B.n679 B.n678 163.367
R1166 B.n675 B.n674 163.367
R1167 B.n671 B.n670 163.367
R1168 B.n667 B.n666 163.367
R1169 B.n663 B.n662 163.367
R1170 B.n659 B.n658 163.367
R1171 B.n655 B.n654 163.367
R1172 B.n651 B.n650 163.367
R1173 B.n647 B.n646 163.367
R1174 B.n643 B.n642 163.367
R1175 B.n639 B.n638 163.367
R1176 B.n635 B.n634 163.367
R1177 B.n631 B.n630 163.367
R1178 B.n627 B.n626 163.367
R1179 B.n622 B.n621 163.367
R1180 B.n618 B.n617 163.367
R1181 B.n614 B.n613 163.367
R1182 B.n610 B.n609 163.367
R1183 B.n606 B.n605 163.367
R1184 B.n602 B.n601 163.367
R1185 B.n598 B.n597 163.367
R1186 B.n594 B.n593 163.367
R1187 B.n590 B.n589 163.367
R1188 B.n586 B.n585 163.367
R1189 B.n582 B.n581 163.367
R1190 B.n578 B.n577 163.367
R1191 B.n574 B.n573 163.367
R1192 B.n570 B.n569 163.367
R1193 B.n566 B.n565 163.367
R1194 B.n562 B.n561 163.367
R1195 B.n558 B.n557 163.367
R1196 B.n554 B.n553 163.367
R1197 B.n550 B.n549 163.367
R1198 B.n546 B.n545 163.367
R1199 B.n542 B.n541 163.367
R1200 B.n538 B.n483 163.367
R1201 B.n740 B.n479 163.367
R1202 B.n740 B.n477 163.367
R1203 B.n744 B.n477 163.367
R1204 B.n744 B.n471 163.367
R1205 B.n752 B.n471 163.367
R1206 B.n752 B.n469 163.367
R1207 B.n756 B.n469 163.367
R1208 B.n756 B.n463 163.367
R1209 B.n764 B.n463 163.367
R1210 B.n764 B.n461 163.367
R1211 B.n768 B.n461 163.367
R1212 B.n768 B.n455 163.367
R1213 B.n776 B.n455 163.367
R1214 B.n776 B.n453 163.367
R1215 B.n780 B.n453 163.367
R1216 B.n780 B.n447 163.367
R1217 B.n788 B.n447 163.367
R1218 B.n788 B.n445 163.367
R1219 B.n792 B.n445 163.367
R1220 B.n792 B.n439 163.367
R1221 B.n801 B.n439 163.367
R1222 B.n801 B.n437 163.367
R1223 B.n805 B.n437 163.367
R1224 B.n805 B.n432 163.367
R1225 B.n813 B.n432 163.367
R1226 B.n813 B.n430 163.367
R1227 B.n817 B.n430 163.367
R1228 B.n817 B.n424 163.367
R1229 B.n825 B.n424 163.367
R1230 B.n825 B.n422 163.367
R1231 B.n829 B.n422 163.367
R1232 B.n829 B.n416 163.367
R1233 B.n837 B.n416 163.367
R1234 B.n837 B.n414 163.367
R1235 B.n841 B.n414 163.367
R1236 B.n841 B.n408 163.367
R1237 B.n849 B.n408 163.367
R1238 B.n849 B.n406 163.367
R1239 B.n853 B.n406 163.367
R1240 B.n853 B.n400 163.367
R1241 B.n861 B.n400 163.367
R1242 B.n861 B.n398 163.367
R1243 B.n865 B.n398 163.367
R1244 B.n865 B.n392 163.367
R1245 B.n873 B.n392 163.367
R1246 B.n873 B.n390 163.367
R1247 B.n877 B.n390 163.367
R1248 B.n877 B.n384 163.367
R1249 B.n885 B.n384 163.367
R1250 B.n885 B.n382 163.367
R1251 B.n889 B.n382 163.367
R1252 B.n889 B.n376 163.367
R1253 B.n898 B.n376 163.367
R1254 B.n898 B.n374 163.367
R1255 B.n902 B.n374 163.367
R1256 B.n902 B.n369 163.367
R1257 B.n911 B.n369 163.367
R1258 B.n911 B.n367 163.367
R1259 B.n915 B.n367 163.367
R1260 B.n915 B.n3 163.367
R1261 B.n1125 B.n3 163.367
R1262 B.n1121 B.n2 163.367
R1263 B.n1121 B.n1120 163.367
R1264 B.n1120 B.n9 163.367
R1265 B.n1116 B.n9 163.367
R1266 B.n1116 B.n11 163.367
R1267 B.n1112 B.n11 163.367
R1268 B.n1112 B.n16 163.367
R1269 B.n1108 B.n16 163.367
R1270 B.n1108 B.n18 163.367
R1271 B.n1104 B.n18 163.367
R1272 B.n1104 B.n24 163.367
R1273 B.n1100 B.n24 163.367
R1274 B.n1100 B.n26 163.367
R1275 B.n1096 B.n26 163.367
R1276 B.n1096 B.n31 163.367
R1277 B.n1092 B.n31 163.367
R1278 B.n1092 B.n33 163.367
R1279 B.n1088 B.n33 163.367
R1280 B.n1088 B.n38 163.367
R1281 B.n1084 B.n38 163.367
R1282 B.n1084 B.n40 163.367
R1283 B.n1080 B.n40 163.367
R1284 B.n1080 B.n45 163.367
R1285 B.n1076 B.n45 163.367
R1286 B.n1076 B.n47 163.367
R1287 B.n1072 B.n47 163.367
R1288 B.n1072 B.n52 163.367
R1289 B.n1068 B.n52 163.367
R1290 B.n1068 B.n54 163.367
R1291 B.n1064 B.n54 163.367
R1292 B.n1064 B.n59 163.367
R1293 B.n1060 B.n59 163.367
R1294 B.n1060 B.n61 163.367
R1295 B.n1056 B.n61 163.367
R1296 B.n1056 B.n66 163.367
R1297 B.n1052 B.n66 163.367
R1298 B.n1052 B.n68 163.367
R1299 B.n1048 B.n68 163.367
R1300 B.n1048 B.n72 163.367
R1301 B.n1044 B.n72 163.367
R1302 B.n1044 B.n74 163.367
R1303 B.n1040 B.n74 163.367
R1304 B.n1040 B.n80 163.367
R1305 B.n1036 B.n80 163.367
R1306 B.n1036 B.n82 163.367
R1307 B.n1032 B.n82 163.367
R1308 B.n1032 B.n87 163.367
R1309 B.n1028 B.n87 163.367
R1310 B.n1028 B.n89 163.367
R1311 B.n1024 B.n89 163.367
R1312 B.n1024 B.n94 163.367
R1313 B.n1020 B.n94 163.367
R1314 B.n1020 B.n96 163.367
R1315 B.n1016 B.n96 163.367
R1316 B.n1016 B.n101 163.367
R1317 B.n1012 B.n101 163.367
R1318 B.n1012 B.n103 163.367
R1319 B.n1008 B.n103 163.367
R1320 B.n1008 B.n108 163.367
R1321 B.n1004 B.n108 163.367
R1322 B.n1004 B.n110 163.367
R1323 B.n163 B.t10 141.352
R1324 B.n536 B.t21 141.352
R1325 B.n166 B.t17 141.335
R1326 B.n533 B.t15 141.335
R1327 B.n732 B.n480 79.7063
R1328 B.n1002 B.n1001 79.7063
R1329 B.n168 B.n113 71.676
R1330 B.n172 B.n114 71.676
R1331 B.n176 B.n115 71.676
R1332 B.n180 B.n116 71.676
R1333 B.n184 B.n117 71.676
R1334 B.n188 B.n118 71.676
R1335 B.n192 B.n119 71.676
R1336 B.n196 B.n120 71.676
R1337 B.n200 B.n121 71.676
R1338 B.n204 B.n122 71.676
R1339 B.n208 B.n123 71.676
R1340 B.n212 B.n124 71.676
R1341 B.n216 B.n125 71.676
R1342 B.n220 B.n126 71.676
R1343 B.n224 B.n127 71.676
R1344 B.n228 B.n128 71.676
R1345 B.n232 B.n129 71.676
R1346 B.n236 B.n130 71.676
R1347 B.n240 B.n131 71.676
R1348 B.n244 B.n132 71.676
R1349 B.n248 B.n133 71.676
R1350 B.n252 B.n134 71.676
R1351 B.n256 B.n135 71.676
R1352 B.n261 B.n136 71.676
R1353 B.n265 B.n137 71.676
R1354 B.n269 B.n138 71.676
R1355 B.n273 B.n139 71.676
R1356 B.n277 B.n140 71.676
R1357 B.n281 B.n141 71.676
R1358 B.n285 B.n142 71.676
R1359 B.n289 B.n143 71.676
R1360 B.n293 B.n144 71.676
R1361 B.n297 B.n145 71.676
R1362 B.n301 B.n146 71.676
R1363 B.n305 B.n147 71.676
R1364 B.n309 B.n148 71.676
R1365 B.n313 B.n149 71.676
R1366 B.n317 B.n150 71.676
R1367 B.n321 B.n151 71.676
R1368 B.n325 B.n152 71.676
R1369 B.n329 B.n153 71.676
R1370 B.n333 B.n154 71.676
R1371 B.n337 B.n155 71.676
R1372 B.n341 B.n156 71.676
R1373 B.n345 B.n157 71.676
R1374 B.n349 B.n158 71.676
R1375 B.n353 B.n159 71.676
R1376 B.n357 B.n160 71.676
R1377 B.n361 B.n161 71.676
R1378 B.n162 B.n161 71.676
R1379 B.n360 B.n160 71.676
R1380 B.n356 B.n159 71.676
R1381 B.n352 B.n158 71.676
R1382 B.n348 B.n157 71.676
R1383 B.n344 B.n156 71.676
R1384 B.n340 B.n155 71.676
R1385 B.n336 B.n154 71.676
R1386 B.n332 B.n153 71.676
R1387 B.n328 B.n152 71.676
R1388 B.n324 B.n151 71.676
R1389 B.n320 B.n150 71.676
R1390 B.n316 B.n149 71.676
R1391 B.n312 B.n148 71.676
R1392 B.n308 B.n147 71.676
R1393 B.n304 B.n146 71.676
R1394 B.n300 B.n145 71.676
R1395 B.n296 B.n144 71.676
R1396 B.n292 B.n143 71.676
R1397 B.n288 B.n142 71.676
R1398 B.n284 B.n141 71.676
R1399 B.n280 B.n140 71.676
R1400 B.n276 B.n139 71.676
R1401 B.n272 B.n138 71.676
R1402 B.n268 B.n137 71.676
R1403 B.n264 B.n136 71.676
R1404 B.n260 B.n135 71.676
R1405 B.n255 B.n134 71.676
R1406 B.n251 B.n133 71.676
R1407 B.n247 B.n132 71.676
R1408 B.n243 B.n131 71.676
R1409 B.n239 B.n130 71.676
R1410 B.n235 B.n129 71.676
R1411 B.n231 B.n128 71.676
R1412 B.n227 B.n127 71.676
R1413 B.n223 B.n126 71.676
R1414 B.n219 B.n125 71.676
R1415 B.n215 B.n124 71.676
R1416 B.n211 B.n123 71.676
R1417 B.n207 B.n122 71.676
R1418 B.n203 B.n121 71.676
R1419 B.n199 B.n120 71.676
R1420 B.n195 B.n119 71.676
R1421 B.n191 B.n118 71.676
R1422 B.n187 B.n117 71.676
R1423 B.n183 B.n116 71.676
R1424 B.n179 B.n115 71.676
R1425 B.n175 B.n114 71.676
R1426 B.n171 B.n113 71.676
R1427 B.n731 B.n730 71.676
R1428 B.n725 B.n484 71.676
R1429 B.n722 B.n485 71.676
R1430 B.n718 B.n486 71.676
R1431 B.n714 B.n487 71.676
R1432 B.n710 B.n488 71.676
R1433 B.n706 B.n489 71.676
R1434 B.n702 B.n490 71.676
R1435 B.n698 B.n491 71.676
R1436 B.n694 B.n492 71.676
R1437 B.n690 B.n493 71.676
R1438 B.n686 B.n494 71.676
R1439 B.n682 B.n495 71.676
R1440 B.n678 B.n496 71.676
R1441 B.n674 B.n497 71.676
R1442 B.n670 B.n498 71.676
R1443 B.n666 B.n499 71.676
R1444 B.n662 B.n500 71.676
R1445 B.n658 B.n501 71.676
R1446 B.n654 B.n502 71.676
R1447 B.n650 B.n503 71.676
R1448 B.n646 B.n504 71.676
R1449 B.n642 B.n505 71.676
R1450 B.n638 B.n506 71.676
R1451 B.n634 B.n507 71.676
R1452 B.n630 B.n508 71.676
R1453 B.n626 B.n509 71.676
R1454 B.n621 B.n510 71.676
R1455 B.n617 B.n511 71.676
R1456 B.n613 B.n512 71.676
R1457 B.n609 B.n513 71.676
R1458 B.n605 B.n514 71.676
R1459 B.n601 B.n515 71.676
R1460 B.n597 B.n516 71.676
R1461 B.n593 B.n517 71.676
R1462 B.n589 B.n518 71.676
R1463 B.n585 B.n519 71.676
R1464 B.n581 B.n520 71.676
R1465 B.n577 B.n521 71.676
R1466 B.n573 B.n522 71.676
R1467 B.n569 B.n523 71.676
R1468 B.n565 B.n524 71.676
R1469 B.n561 B.n525 71.676
R1470 B.n557 B.n526 71.676
R1471 B.n553 B.n527 71.676
R1472 B.n549 B.n528 71.676
R1473 B.n545 B.n529 71.676
R1474 B.n541 B.n530 71.676
R1475 B.n733 B.n483 71.676
R1476 B.n731 B.n532 71.676
R1477 B.n723 B.n484 71.676
R1478 B.n719 B.n485 71.676
R1479 B.n715 B.n486 71.676
R1480 B.n711 B.n487 71.676
R1481 B.n707 B.n488 71.676
R1482 B.n703 B.n489 71.676
R1483 B.n699 B.n490 71.676
R1484 B.n695 B.n491 71.676
R1485 B.n691 B.n492 71.676
R1486 B.n687 B.n493 71.676
R1487 B.n683 B.n494 71.676
R1488 B.n679 B.n495 71.676
R1489 B.n675 B.n496 71.676
R1490 B.n671 B.n497 71.676
R1491 B.n667 B.n498 71.676
R1492 B.n663 B.n499 71.676
R1493 B.n659 B.n500 71.676
R1494 B.n655 B.n501 71.676
R1495 B.n651 B.n502 71.676
R1496 B.n647 B.n503 71.676
R1497 B.n643 B.n504 71.676
R1498 B.n639 B.n505 71.676
R1499 B.n635 B.n506 71.676
R1500 B.n631 B.n507 71.676
R1501 B.n627 B.n508 71.676
R1502 B.n622 B.n509 71.676
R1503 B.n618 B.n510 71.676
R1504 B.n614 B.n511 71.676
R1505 B.n610 B.n512 71.676
R1506 B.n606 B.n513 71.676
R1507 B.n602 B.n514 71.676
R1508 B.n598 B.n515 71.676
R1509 B.n594 B.n516 71.676
R1510 B.n590 B.n517 71.676
R1511 B.n586 B.n518 71.676
R1512 B.n582 B.n519 71.676
R1513 B.n578 B.n520 71.676
R1514 B.n574 B.n521 71.676
R1515 B.n570 B.n522 71.676
R1516 B.n566 B.n523 71.676
R1517 B.n562 B.n524 71.676
R1518 B.n558 B.n525 71.676
R1519 B.n554 B.n526 71.676
R1520 B.n550 B.n527 71.676
R1521 B.n546 B.n528 71.676
R1522 B.n542 B.n529 71.676
R1523 B.n538 B.n530 71.676
R1524 B.n734 B.n733 71.676
R1525 B.n1126 B.n1125 71.676
R1526 B.n1126 B.n2 71.676
R1527 B.n164 B.t11 70.7582
R1528 B.n537 B.t20 70.7582
R1529 B.n167 B.t18 70.7415
R1530 B.n534 B.t14 70.7415
R1531 B.n167 B.n166 70.5944
R1532 B.n164 B.n163 70.5944
R1533 B.n537 B.n536 70.5944
R1534 B.n534 B.n533 70.5944
R1535 B.n258 B.n167 59.5399
R1536 B.n165 B.n164 59.5399
R1537 B.n624 B.n537 59.5399
R1538 B.n535 B.n534 59.5399
R1539 B.n739 B.n480 40.7523
R1540 B.n739 B.n476 40.7523
R1541 B.n745 B.n476 40.7523
R1542 B.n745 B.n472 40.7523
R1543 B.n751 B.n472 40.7523
R1544 B.n751 B.n467 40.7523
R1545 B.n757 B.n467 40.7523
R1546 B.n757 B.n468 40.7523
R1547 B.n763 B.n460 40.7523
R1548 B.n769 B.n460 40.7523
R1549 B.n769 B.n456 40.7523
R1550 B.n775 B.n456 40.7523
R1551 B.n775 B.n452 40.7523
R1552 B.n781 B.n452 40.7523
R1553 B.n781 B.n448 40.7523
R1554 B.n787 B.n448 40.7523
R1555 B.n787 B.n444 40.7523
R1556 B.n793 B.n444 40.7523
R1557 B.n793 B.n440 40.7523
R1558 B.n800 B.n440 40.7523
R1559 B.n800 B.n799 40.7523
R1560 B.n806 B.n433 40.7523
R1561 B.n812 B.n433 40.7523
R1562 B.n812 B.n429 40.7523
R1563 B.n818 B.n429 40.7523
R1564 B.n818 B.n425 40.7523
R1565 B.n824 B.n425 40.7523
R1566 B.n824 B.n421 40.7523
R1567 B.n830 B.n421 40.7523
R1568 B.n830 B.n417 40.7523
R1569 B.n836 B.n417 40.7523
R1570 B.n842 B.n413 40.7523
R1571 B.n842 B.n409 40.7523
R1572 B.n848 B.n409 40.7523
R1573 B.n848 B.n405 40.7523
R1574 B.n854 B.n405 40.7523
R1575 B.n854 B.n401 40.7523
R1576 B.n860 B.n401 40.7523
R1577 B.n860 B.n397 40.7523
R1578 B.n866 B.n397 40.7523
R1579 B.n872 B.n393 40.7523
R1580 B.n872 B.n389 40.7523
R1581 B.n878 B.n389 40.7523
R1582 B.n878 B.n385 40.7523
R1583 B.n884 B.n385 40.7523
R1584 B.n884 B.n381 40.7523
R1585 B.n890 B.n381 40.7523
R1586 B.n890 B.n377 40.7523
R1587 B.n897 B.n377 40.7523
R1588 B.n897 B.n896 40.7523
R1589 B.n903 B.n370 40.7523
R1590 B.n910 B.n370 40.7523
R1591 B.n910 B.n366 40.7523
R1592 B.n916 B.n366 40.7523
R1593 B.n916 B.n4 40.7523
R1594 B.n1124 B.n4 40.7523
R1595 B.n1124 B.n1123 40.7523
R1596 B.n1123 B.n1122 40.7523
R1597 B.n1122 B.n8 40.7523
R1598 B.n12 B.n8 40.7523
R1599 B.n1115 B.n12 40.7523
R1600 B.n1115 B.n1114 40.7523
R1601 B.n1114 B.n1113 40.7523
R1602 B.n1107 B.n19 40.7523
R1603 B.n1107 B.n1106 40.7523
R1604 B.n1106 B.n1105 40.7523
R1605 B.n1105 B.n23 40.7523
R1606 B.n1099 B.n23 40.7523
R1607 B.n1099 B.n1098 40.7523
R1608 B.n1098 B.n1097 40.7523
R1609 B.n1097 B.n30 40.7523
R1610 B.n1091 B.n30 40.7523
R1611 B.n1091 B.n1090 40.7523
R1612 B.n1089 B.n37 40.7523
R1613 B.n1083 B.n37 40.7523
R1614 B.n1083 B.n1082 40.7523
R1615 B.n1082 B.n1081 40.7523
R1616 B.n1081 B.n44 40.7523
R1617 B.n1075 B.n44 40.7523
R1618 B.n1075 B.n1074 40.7523
R1619 B.n1074 B.n1073 40.7523
R1620 B.n1073 B.n51 40.7523
R1621 B.n1067 B.n1066 40.7523
R1622 B.n1066 B.n1065 40.7523
R1623 B.n1065 B.n58 40.7523
R1624 B.n1059 B.n58 40.7523
R1625 B.n1059 B.n1058 40.7523
R1626 B.n1058 B.n1057 40.7523
R1627 B.n1057 B.n65 40.7523
R1628 B.n1051 B.n65 40.7523
R1629 B.n1051 B.n1050 40.7523
R1630 B.n1050 B.n1049 40.7523
R1631 B.n1043 B.n75 40.7523
R1632 B.n1043 B.n1042 40.7523
R1633 B.n1042 B.n1041 40.7523
R1634 B.n1041 B.n79 40.7523
R1635 B.n1035 B.n79 40.7523
R1636 B.n1035 B.n1034 40.7523
R1637 B.n1034 B.n1033 40.7523
R1638 B.n1033 B.n86 40.7523
R1639 B.n1027 B.n86 40.7523
R1640 B.n1027 B.n1026 40.7523
R1641 B.n1026 B.n1025 40.7523
R1642 B.n1025 B.n93 40.7523
R1643 B.n1019 B.n93 40.7523
R1644 B.n1018 B.n1017 40.7523
R1645 B.n1017 B.n100 40.7523
R1646 B.n1011 B.n100 40.7523
R1647 B.n1011 B.n1010 40.7523
R1648 B.n1010 B.n1009 40.7523
R1649 B.n1009 B.n107 40.7523
R1650 B.n1003 B.n107 40.7523
R1651 B.n1003 B.n1002 40.7523
R1652 B.t2 B.n413 35.3587
R1653 B.t5 B.n51 35.3587
R1654 B.n729 B.n478 34.8103
R1655 B.n736 B.n735 34.8103
R1656 B.n999 B.n998 34.8103
R1657 B.n169 B.n109 34.8103
R1658 B.n866 B.t7 34.1601
R1659 B.t6 B.n1089 34.1601
R1660 B.n806 B.t1 23.3729
R1661 B.n1049 B.t4 23.3729
R1662 B.n896 B.t3 22.1743
R1663 B.n19 B.t0 22.1743
R1664 B.n468 B.t13 20.9757
R1665 B.t9 B.n1018 20.9757
R1666 B.n763 B.t13 19.7771
R1667 B.n1019 B.t9 19.7771
R1668 B.n903 B.t3 18.5785
R1669 B.n1113 B.t0 18.5785
R1670 B B.n1127 18.0485
R1671 B.n799 B.t1 17.38
R1672 B.n75 B.t4 17.38
R1673 B.n741 B.n478 10.6151
R1674 B.n742 B.n741 10.6151
R1675 B.n743 B.n742 10.6151
R1676 B.n743 B.n470 10.6151
R1677 B.n753 B.n470 10.6151
R1678 B.n754 B.n753 10.6151
R1679 B.n755 B.n754 10.6151
R1680 B.n755 B.n462 10.6151
R1681 B.n765 B.n462 10.6151
R1682 B.n766 B.n765 10.6151
R1683 B.n767 B.n766 10.6151
R1684 B.n767 B.n454 10.6151
R1685 B.n777 B.n454 10.6151
R1686 B.n778 B.n777 10.6151
R1687 B.n779 B.n778 10.6151
R1688 B.n779 B.n446 10.6151
R1689 B.n789 B.n446 10.6151
R1690 B.n790 B.n789 10.6151
R1691 B.n791 B.n790 10.6151
R1692 B.n791 B.n438 10.6151
R1693 B.n802 B.n438 10.6151
R1694 B.n803 B.n802 10.6151
R1695 B.n804 B.n803 10.6151
R1696 B.n804 B.n431 10.6151
R1697 B.n814 B.n431 10.6151
R1698 B.n815 B.n814 10.6151
R1699 B.n816 B.n815 10.6151
R1700 B.n816 B.n423 10.6151
R1701 B.n826 B.n423 10.6151
R1702 B.n827 B.n826 10.6151
R1703 B.n828 B.n827 10.6151
R1704 B.n828 B.n415 10.6151
R1705 B.n838 B.n415 10.6151
R1706 B.n839 B.n838 10.6151
R1707 B.n840 B.n839 10.6151
R1708 B.n840 B.n407 10.6151
R1709 B.n850 B.n407 10.6151
R1710 B.n851 B.n850 10.6151
R1711 B.n852 B.n851 10.6151
R1712 B.n852 B.n399 10.6151
R1713 B.n862 B.n399 10.6151
R1714 B.n863 B.n862 10.6151
R1715 B.n864 B.n863 10.6151
R1716 B.n864 B.n391 10.6151
R1717 B.n874 B.n391 10.6151
R1718 B.n875 B.n874 10.6151
R1719 B.n876 B.n875 10.6151
R1720 B.n876 B.n383 10.6151
R1721 B.n886 B.n383 10.6151
R1722 B.n887 B.n886 10.6151
R1723 B.n888 B.n887 10.6151
R1724 B.n888 B.n375 10.6151
R1725 B.n899 B.n375 10.6151
R1726 B.n900 B.n899 10.6151
R1727 B.n901 B.n900 10.6151
R1728 B.n901 B.n368 10.6151
R1729 B.n912 B.n368 10.6151
R1730 B.n913 B.n912 10.6151
R1731 B.n914 B.n913 10.6151
R1732 B.n914 B.n0 10.6151
R1733 B.n729 B.n728 10.6151
R1734 B.n728 B.n727 10.6151
R1735 B.n727 B.n726 10.6151
R1736 B.n726 B.n724 10.6151
R1737 B.n724 B.n721 10.6151
R1738 B.n721 B.n720 10.6151
R1739 B.n720 B.n717 10.6151
R1740 B.n717 B.n716 10.6151
R1741 B.n716 B.n713 10.6151
R1742 B.n713 B.n712 10.6151
R1743 B.n712 B.n709 10.6151
R1744 B.n709 B.n708 10.6151
R1745 B.n708 B.n705 10.6151
R1746 B.n705 B.n704 10.6151
R1747 B.n704 B.n701 10.6151
R1748 B.n701 B.n700 10.6151
R1749 B.n700 B.n697 10.6151
R1750 B.n697 B.n696 10.6151
R1751 B.n696 B.n693 10.6151
R1752 B.n693 B.n692 10.6151
R1753 B.n692 B.n689 10.6151
R1754 B.n689 B.n688 10.6151
R1755 B.n688 B.n685 10.6151
R1756 B.n685 B.n684 10.6151
R1757 B.n684 B.n681 10.6151
R1758 B.n681 B.n680 10.6151
R1759 B.n680 B.n677 10.6151
R1760 B.n677 B.n676 10.6151
R1761 B.n676 B.n673 10.6151
R1762 B.n673 B.n672 10.6151
R1763 B.n672 B.n669 10.6151
R1764 B.n669 B.n668 10.6151
R1765 B.n668 B.n665 10.6151
R1766 B.n665 B.n664 10.6151
R1767 B.n664 B.n661 10.6151
R1768 B.n661 B.n660 10.6151
R1769 B.n660 B.n657 10.6151
R1770 B.n657 B.n656 10.6151
R1771 B.n656 B.n653 10.6151
R1772 B.n653 B.n652 10.6151
R1773 B.n652 B.n649 10.6151
R1774 B.n649 B.n648 10.6151
R1775 B.n648 B.n645 10.6151
R1776 B.n645 B.n644 10.6151
R1777 B.n641 B.n640 10.6151
R1778 B.n640 B.n637 10.6151
R1779 B.n637 B.n636 10.6151
R1780 B.n636 B.n633 10.6151
R1781 B.n633 B.n632 10.6151
R1782 B.n632 B.n629 10.6151
R1783 B.n629 B.n628 10.6151
R1784 B.n628 B.n625 10.6151
R1785 B.n623 B.n620 10.6151
R1786 B.n620 B.n619 10.6151
R1787 B.n619 B.n616 10.6151
R1788 B.n616 B.n615 10.6151
R1789 B.n615 B.n612 10.6151
R1790 B.n612 B.n611 10.6151
R1791 B.n611 B.n608 10.6151
R1792 B.n608 B.n607 10.6151
R1793 B.n607 B.n604 10.6151
R1794 B.n604 B.n603 10.6151
R1795 B.n603 B.n600 10.6151
R1796 B.n600 B.n599 10.6151
R1797 B.n599 B.n596 10.6151
R1798 B.n596 B.n595 10.6151
R1799 B.n595 B.n592 10.6151
R1800 B.n592 B.n591 10.6151
R1801 B.n591 B.n588 10.6151
R1802 B.n588 B.n587 10.6151
R1803 B.n587 B.n584 10.6151
R1804 B.n584 B.n583 10.6151
R1805 B.n583 B.n580 10.6151
R1806 B.n580 B.n579 10.6151
R1807 B.n579 B.n576 10.6151
R1808 B.n576 B.n575 10.6151
R1809 B.n575 B.n572 10.6151
R1810 B.n572 B.n571 10.6151
R1811 B.n571 B.n568 10.6151
R1812 B.n568 B.n567 10.6151
R1813 B.n567 B.n564 10.6151
R1814 B.n564 B.n563 10.6151
R1815 B.n563 B.n560 10.6151
R1816 B.n560 B.n559 10.6151
R1817 B.n559 B.n556 10.6151
R1818 B.n556 B.n555 10.6151
R1819 B.n555 B.n552 10.6151
R1820 B.n552 B.n551 10.6151
R1821 B.n551 B.n548 10.6151
R1822 B.n548 B.n547 10.6151
R1823 B.n547 B.n544 10.6151
R1824 B.n544 B.n543 10.6151
R1825 B.n543 B.n540 10.6151
R1826 B.n540 B.n539 10.6151
R1827 B.n539 B.n482 10.6151
R1828 B.n735 B.n482 10.6151
R1829 B.n737 B.n736 10.6151
R1830 B.n737 B.n474 10.6151
R1831 B.n747 B.n474 10.6151
R1832 B.n748 B.n747 10.6151
R1833 B.n749 B.n748 10.6151
R1834 B.n749 B.n465 10.6151
R1835 B.n759 B.n465 10.6151
R1836 B.n760 B.n759 10.6151
R1837 B.n761 B.n760 10.6151
R1838 B.n761 B.n458 10.6151
R1839 B.n771 B.n458 10.6151
R1840 B.n772 B.n771 10.6151
R1841 B.n773 B.n772 10.6151
R1842 B.n773 B.n450 10.6151
R1843 B.n783 B.n450 10.6151
R1844 B.n784 B.n783 10.6151
R1845 B.n785 B.n784 10.6151
R1846 B.n785 B.n442 10.6151
R1847 B.n795 B.n442 10.6151
R1848 B.n796 B.n795 10.6151
R1849 B.n797 B.n796 10.6151
R1850 B.n797 B.n435 10.6151
R1851 B.n808 B.n435 10.6151
R1852 B.n809 B.n808 10.6151
R1853 B.n810 B.n809 10.6151
R1854 B.n810 B.n427 10.6151
R1855 B.n820 B.n427 10.6151
R1856 B.n821 B.n820 10.6151
R1857 B.n822 B.n821 10.6151
R1858 B.n822 B.n419 10.6151
R1859 B.n832 B.n419 10.6151
R1860 B.n833 B.n832 10.6151
R1861 B.n834 B.n833 10.6151
R1862 B.n834 B.n411 10.6151
R1863 B.n844 B.n411 10.6151
R1864 B.n845 B.n844 10.6151
R1865 B.n846 B.n845 10.6151
R1866 B.n846 B.n403 10.6151
R1867 B.n856 B.n403 10.6151
R1868 B.n857 B.n856 10.6151
R1869 B.n858 B.n857 10.6151
R1870 B.n858 B.n395 10.6151
R1871 B.n868 B.n395 10.6151
R1872 B.n869 B.n868 10.6151
R1873 B.n870 B.n869 10.6151
R1874 B.n870 B.n387 10.6151
R1875 B.n880 B.n387 10.6151
R1876 B.n881 B.n880 10.6151
R1877 B.n882 B.n881 10.6151
R1878 B.n882 B.n379 10.6151
R1879 B.n892 B.n379 10.6151
R1880 B.n893 B.n892 10.6151
R1881 B.n894 B.n893 10.6151
R1882 B.n894 B.n372 10.6151
R1883 B.n905 B.n372 10.6151
R1884 B.n906 B.n905 10.6151
R1885 B.n908 B.n906 10.6151
R1886 B.n908 B.n907 10.6151
R1887 B.n907 B.n364 10.6151
R1888 B.n919 B.n364 10.6151
R1889 B.n920 B.n919 10.6151
R1890 B.n921 B.n920 10.6151
R1891 B.n922 B.n921 10.6151
R1892 B.n923 B.n922 10.6151
R1893 B.n926 B.n923 10.6151
R1894 B.n927 B.n926 10.6151
R1895 B.n928 B.n927 10.6151
R1896 B.n929 B.n928 10.6151
R1897 B.n931 B.n929 10.6151
R1898 B.n932 B.n931 10.6151
R1899 B.n933 B.n932 10.6151
R1900 B.n934 B.n933 10.6151
R1901 B.n936 B.n934 10.6151
R1902 B.n937 B.n936 10.6151
R1903 B.n938 B.n937 10.6151
R1904 B.n939 B.n938 10.6151
R1905 B.n941 B.n939 10.6151
R1906 B.n942 B.n941 10.6151
R1907 B.n943 B.n942 10.6151
R1908 B.n944 B.n943 10.6151
R1909 B.n946 B.n944 10.6151
R1910 B.n947 B.n946 10.6151
R1911 B.n948 B.n947 10.6151
R1912 B.n949 B.n948 10.6151
R1913 B.n951 B.n949 10.6151
R1914 B.n952 B.n951 10.6151
R1915 B.n953 B.n952 10.6151
R1916 B.n954 B.n953 10.6151
R1917 B.n956 B.n954 10.6151
R1918 B.n957 B.n956 10.6151
R1919 B.n958 B.n957 10.6151
R1920 B.n959 B.n958 10.6151
R1921 B.n961 B.n959 10.6151
R1922 B.n962 B.n961 10.6151
R1923 B.n963 B.n962 10.6151
R1924 B.n964 B.n963 10.6151
R1925 B.n966 B.n964 10.6151
R1926 B.n967 B.n966 10.6151
R1927 B.n968 B.n967 10.6151
R1928 B.n969 B.n968 10.6151
R1929 B.n971 B.n969 10.6151
R1930 B.n972 B.n971 10.6151
R1931 B.n973 B.n972 10.6151
R1932 B.n974 B.n973 10.6151
R1933 B.n976 B.n974 10.6151
R1934 B.n977 B.n976 10.6151
R1935 B.n978 B.n977 10.6151
R1936 B.n979 B.n978 10.6151
R1937 B.n981 B.n979 10.6151
R1938 B.n982 B.n981 10.6151
R1939 B.n983 B.n982 10.6151
R1940 B.n984 B.n983 10.6151
R1941 B.n986 B.n984 10.6151
R1942 B.n987 B.n986 10.6151
R1943 B.n988 B.n987 10.6151
R1944 B.n989 B.n988 10.6151
R1945 B.n991 B.n989 10.6151
R1946 B.n992 B.n991 10.6151
R1947 B.n993 B.n992 10.6151
R1948 B.n994 B.n993 10.6151
R1949 B.n996 B.n994 10.6151
R1950 B.n997 B.n996 10.6151
R1951 B.n998 B.n997 10.6151
R1952 B.n1119 B.n1 10.6151
R1953 B.n1119 B.n1118 10.6151
R1954 B.n1118 B.n1117 10.6151
R1955 B.n1117 B.n10 10.6151
R1956 B.n1111 B.n10 10.6151
R1957 B.n1111 B.n1110 10.6151
R1958 B.n1110 B.n1109 10.6151
R1959 B.n1109 B.n17 10.6151
R1960 B.n1103 B.n17 10.6151
R1961 B.n1103 B.n1102 10.6151
R1962 B.n1102 B.n1101 10.6151
R1963 B.n1101 B.n25 10.6151
R1964 B.n1095 B.n25 10.6151
R1965 B.n1095 B.n1094 10.6151
R1966 B.n1094 B.n1093 10.6151
R1967 B.n1093 B.n32 10.6151
R1968 B.n1087 B.n32 10.6151
R1969 B.n1087 B.n1086 10.6151
R1970 B.n1086 B.n1085 10.6151
R1971 B.n1085 B.n39 10.6151
R1972 B.n1079 B.n39 10.6151
R1973 B.n1079 B.n1078 10.6151
R1974 B.n1078 B.n1077 10.6151
R1975 B.n1077 B.n46 10.6151
R1976 B.n1071 B.n46 10.6151
R1977 B.n1071 B.n1070 10.6151
R1978 B.n1070 B.n1069 10.6151
R1979 B.n1069 B.n53 10.6151
R1980 B.n1063 B.n53 10.6151
R1981 B.n1063 B.n1062 10.6151
R1982 B.n1062 B.n1061 10.6151
R1983 B.n1061 B.n60 10.6151
R1984 B.n1055 B.n60 10.6151
R1985 B.n1055 B.n1054 10.6151
R1986 B.n1054 B.n1053 10.6151
R1987 B.n1053 B.n67 10.6151
R1988 B.n1047 B.n67 10.6151
R1989 B.n1047 B.n1046 10.6151
R1990 B.n1046 B.n1045 10.6151
R1991 B.n1045 B.n73 10.6151
R1992 B.n1039 B.n73 10.6151
R1993 B.n1039 B.n1038 10.6151
R1994 B.n1038 B.n1037 10.6151
R1995 B.n1037 B.n81 10.6151
R1996 B.n1031 B.n81 10.6151
R1997 B.n1031 B.n1030 10.6151
R1998 B.n1030 B.n1029 10.6151
R1999 B.n1029 B.n88 10.6151
R2000 B.n1023 B.n88 10.6151
R2001 B.n1023 B.n1022 10.6151
R2002 B.n1022 B.n1021 10.6151
R2003 B.n1021 B.n95 10.6151
R2004 B.n1015 B.n95 10.6151
R2005 B.n1015 B.n1014 10.6151
R2006 B.n1014 B.n1013 10.6151
R2007 B.n1013 B.n102 10.6151
R2008 B.n1007 B.n102 10.6151
R2009 B.n1007 B.n1006 10.6151
R2010 B.n1006 B.n1005 10.6151
R2011 B.n1005 B.n109 10.6151
R2012 B.n170 B.n169 10.6151
R2013 B.n173 B.n170 10.6151
R2014 B.n174 B.n173 10.6151
R2015 B.n177 B.n174 10.6151
R2016 B.n178 B.n177 10.6151
R2017 B.n181 B.n178 10.6151
R2018 B.n182 B.n181 10.6151
R2019 B.n185 B.n182 10.6151
R2020 B.n186 B.n185 10.6151
R2021 B.n189 B.n186 10.6151
R2022 B.n190 B.n189 10.6151
R2023 B.n193 B.n190 10.6151
R2024 B.n194 B.n193 10.6151
R2025 B.n197 B.n194 10.6151
R2026 B.n198 B.n197 10.6151
R2027 B.n201 B.n198 10.6151
R2028 B.n202 B.n201 10.6151
R2029 B.n205 B.n202 10.6151
R2030 B.n206 B.n205 10.6151
R2031 B.n209 B.n206 10.6151
R2032 B.n210 B.n209 10.6151
R2033 B.n213 B.n210 10.6151
R2034 B.n214 B.n213 10.6151
R2035 B.n217 B.n214 10.6151
R2036 B.n218 B.n217 10.6151
R2037 B.n221 B.n218 10.6151
R2038 B.n222 B.n221 10.6151
R2039 B.n225 B.n222 10.6151
R2040 B.n226 B.n225 10.6151
R2041 B.n229 B.n226 10.6151
R2042 B.n230 B.n229 10.6151
R2043 B.n233 B.n230 10.6151
R2044 B.n234 B.n233 10.6151
R2045 B.n237 B.n234 10.6151
R2046 B.n238 B.n237 10.6151
R2047 B.n241 B.n238 10.6151
R2048 B.n242 B.n241 10.6151
R2049 B.n245 B.n242 10.6151
R2050 B.n246 B.n245 10.6151
R2051 B.n249 B.n246 10.6151
R2052 B.n250 B.n249 10.6151
R2053 B.n253 B.n250 10.6151
R2054 B.n254 B.n253 10.6151
R2055 B.n257 B.n254 10.6151
R2056 B.n262 B.n259 10.6151
R2057 B.n263 B.n262 10.6151
R2058 B.n266 B.n263 10.6151
R2059 B.n267 B.n266 10.6151
R2060 B.n270 B.n267 10.6151
R2061 B.n271 B.n270 10.6151
R2062 B.n274 B.n271 10.6151
R2063 B.n275 B.n274 10.6151
R2064 B.n279 B.n278 10.6151
R2065 B.n282 B.n279 10.6151
R2066 B.n283 B.n282 10.6151
R2067 B.n286 B.n283 10.6151
R2068 B.n287 B.n286 10.6151
R2069 B.n290 B.n287 10.6151
R2070 B.n291 B.n290 10.6151
R2071 B.n294 B.n291 10.6151
R2072 B.n295 B.n294 10.6151
R2073 B.n298 B.n295 10.6151
R2074 B.n299 B.n298 10.6151
R2075 B.n302 B.n299 10.6151
R2076 B.n303 B.n302 10.6151
R2077 B.n306 B.n303 10.6151
R2078 B.n307 B.n306 10.6151
R2079 B.n310 B.n307 10.6151
R2080 B.n311 B.n310 10.6151
R2081 B.n314 B.n311 10.6151
R2082 B.n315 B.n314 10.6151
R2083 B.n318 B.n315 10.6151
R2084 B.n319 B.n318 10.6151
R2085 B.n322 B.n319 10.6151
R2086 B.n323 B.n322 10.6151
R2087 B.n326 B.n323 10.6151
R2088 B.n327 B.n326 10.6151
R2089 B.n330 B.n327 10.6151
R2090 B.n331 B.n330 10.6151
R2091 B.n334 B.n331 10.6151
R2092 B.n335 B.n334 10.6151
R2093 B.n338 B.n335 10.6151
R2094 B.n339 B.n338 10.6151
R2095 B.n342 B.n339 10.6151
R2096 B.n343 B.n342 10.6151
R2097 B.n346 B.n343 10.6151
R2098 B.n347 B.n346 10.6151
R2099 B.n350 B.n347 10.6151
R2100 B.n351 B.n350 10.6151
R2101 B.n354 B.n351 10.6151
R2102 B.n355 B.n354 10.6151
R2103 B.n358 B.n355 10.6151
R2104 B.n359 B.n358 10.6151
R2105 B.n362 B.n359 10.6151
R2106 B.n363 B.n362 10.6151
R2107 B.n999 B.n363 10.6151
R2108 B.n1127 B.n0 8.11757
R2109 B.n1127 B.n1 8.11757
R2110 B.t7 B.n393 6.59271
R2111 B.n1090 B.t6 6.59271
R2112 B.n641 B.n535 6.5566
R2113 B.n625 B.n624 6.5566
R2114 B.n259 B.n258 6.5566
R2115 B.n275 B.n165 6.5566
R2116 B.n836 B.t2 5.39413
R2117 B.n1067 B.t5 5.39413
R2118 B.n644 B.n535 4.05904
R2119 B.n624 B.n623 4.05904
R2120 B.n258 B.n257 4.05904
R2121 B.n278 B.n165 4.05904
R2122 VN.n68 VN.n67 161.3
R2123 VN.n66 VN.n36 161.3
R2124 VN.n65 VN.n64 161.3
R2125 VN.n63 VN.n37 161.3
R2126 VN.n62 VN.n61 161.3
R2127 VN.n60 VN.n38 161.3
R2128 VN.n59 VN.n58 161.3
R2129 VN.n57 VN.n56 161.3
R2130 VN.n55 VN.n40 161.3
R2131 VN.n54 VN.n53 161.3
R2132 VN.n52 VN.n41 161.3
R2133 VN.n51 VN.n50 161.3
R2134 VN.n49 VN.n42 161.3
R2135 VN.n48 VN.n47 161.3
R2136 VN.n46 VN.n43 161.3
R2137 VN.n33 VN.n32 161.3
R2138 VN.n31 VN.n1 161.3
R2139 VN.n30 VN.n29 161.3
R2140 VN.n28 VN.n2 161.3
R2141 VN.n27 VN.n26 161.3
R2142 VN.n25 VN.n3 161.3
R2143 VN.n24 VN.n23 161.3
R2144 VN.n22 VN.n21 161.3
R2145 VN.n20 VN.n5 161.3
R2146 VN.n19 VN.n18 161.3
R2147 VN.n17 VN.n6 161.3
R2148 VN.n16 VN.n15 161.3
R2149 VN.n14 VN.n7 161.3
R2150 VN.n13 VN.n12 161.3
R2151 VN.n11 VN.n8 161.3
R2152 VN.n45 VN.t5 127.492
R2153 VN.n10 VN.t1 127.492
R2154 VN.n9 VN.t3 95.2355
R2155 VN.n4 VN.t6 95.2355
R2156 VN.n0 VN.t7 95.2355
R2157 VN.n44 VN.t4 95.2355
R2158 VN.n39 VN.t2 95.2355
R2159 VN.n35 VN.t0 95.2355
R2160 VN.n34 VN.n0 79.917
R2161 VN.n69 VN.n35 79.917
R2162 VN.n10 VN.n9 71.3663
R2163 VN.n45 VN.n44 71.3663
R2164 VN.n15 VN.n6 56.5617
R2165 VN.n50 VN.n41 56.5617
R2166 VN VN.n69 55.2481
R2167 VN.n26 VN.n2 51.2335
R2168 VN.n61 VN.n37 51.2335
R2169 VN.n30 VN.n2 29.9206
R2170 VN.n65 VN.n37 29.9206
R2171 VN.n13 VN.n8 24.5923
R2172 VN.n14 VN.n13 24.5923
R2173 VN.n15 VN.n14 24.5923
R2174 VN.n19 VN.n6 24.5923
R2175 VN.n20 VN.n19 24.5923
R2176 VN.n21 VN.n20 24.5923
R2177 VN.n25 VN.n24 24.5923
R2178 VN.n26 VN.n25 24.5923
R2179 VN.n31 VN.n30 24.5923
R2180 VN.n32 VN.n31 24.5923
R2181 VN.n50 VN.n49 24.5923
R2182 VN.n49 VN.n48 24.5923
R2183 VN.n48 VN.n43 24.5923
R2184 VN.n61 VN.n60 24.5923
R2185 VN.n60 VN.n59 24.5923
R2186 VN.n56 VN.n55 24.5923
R2187 VN.n55 VN.n54 24.5923
R2188 VN.n54 VN.n41 24.5923
R2189 VN.n67 VN.n66 24.5923
R2190 VN.n66 VN.n65 24.5923
R2191 VN.n24 VN.n4 21.1495
R2192 VN.n59 VN.n39 21.1495
R2193 VN.n32 VN.n0 10.3291
R2194 VN.n67 VN.n35 10.3291
R2195 VN.n46 VN.n45 4.37641
R2196 VN.n11 VN.n10 4.37641
R2197 VN.n9 VN.n8 3.44336
R2198 VN.n21 VN.n4 3.44336
R2199 VN.n44 VN.n43 3.44336
R2200 VN.n56 VN.n39 3.44336
R2201 VN.n69 VN.n68 0.354861
R2202 VN.n34 VN.n33 0.354861
R2203 VN VN.n34 0.267071
R2204 VN.n68 VN.n36 0.189894
R2205 VN.n64 VN.n36 0.189894
R2206 VN.n64 VN.n63 0.189894
R2207 VN.n63 VN.n62 0.189894
R2208 VN.n62 VN.n38 0.189894
R2209 VN.n58 VN.n38 0.189894
R2210 VN.n58 VN.n57 0.189894
R2211 VN.n57 VN.n40 0.189894
R2212 VN.n53 VN.n40 0.189894
R2213 VN.n53 VN.n52 0.189894
R2214 VN.n52 VN.n51 0.189894
R2215 VN.n51 VN.n42 0.189894
R2216 VN.n47 VN.n42 0.189894
R2217 VN.n47 VN.n46 0.189894
R2218 VN.n12 VN.n11 0.189894
R2219 VN.n12 VN.n7 0.189894
R2220 VN.n16 VN.n7 0.189894
R2221 VN.n17 VN.n16 0.189894
R2222 VN.n18 VN.n17 0.189894
R2223 VN.n18 VN.n5 0.189894
R2224 VN.n22 VN.n5 0.189894
R2225 VN.n23 VN.n22 0.189894
R2226 VN.n23 VN.n3 0.189894
R2227 VN.n27 VN.n3 0.189894
R2228 VN.n28 VN.n27 0.189894
R2229 VN.n29 VN.n28 0.189894
R2230 VN.n29 VN.n1 0.189894
R2231 VN.n33 VN.n1 0.189894
R2232 VDD2.n2 VDD2.n1 60.8116
R2233 VDD2.n2 VDD2.n0 60.8116
R2234 VDD2 VDD2.n5 60.8086
R2235 VDD2.n4 VDD2.n3 59.298
R2236 VDD2.n4 VDD2.n2 49.1118
R2237 VDD2 VDD2.n4 1.62766
R2238 VDD2.n5 VDD2.t3 1.51426
R2239 VDD2.n5 VDD2.t2 1.51426
R2240 VDD2.n3 VDD2.t7 1.51426
R2241 VDD2.n3 VDD2.t5 1.51426
R2242 VDD2.n1 VDD2.t1 1.51426
R2243 VDD2.n1 VDD2.t0 1.51426
R2244 VDD2.n0 VDD2.t6 1.51426
R2245 VDD2.n0 VDD2.t4 1.51426
C0 VDD2 VTAIL 8.709411f
C1 VDD1 VTAIL 8.65023f
C2 VP VN 8.72782f
C3 VP VDD2 0.595474f
C4 VP VDD1 10.286901f
C5 VN VDD2 9.84647f
C6 VN VDD1 0.153263f
C7 VP VTAIL 10.441401f
C8 VDD1 VDD2 2.14406f
C9 VN VTAIL 10.4273f
C10 VDD2 B 6.199242f
C11 VDD1 B 6.718574f
C12 VTAIL B 11.62276f
C13 VN B 18.318329f
C14 VP B 16.954744f
C15 VDD2.t6 B 0.276673f
C16 VDD2.t4 B 0.276673f
C17 VDD2.n0 B 2.49024f
C18 VDD2.t1 B 0.276673f
C19 VDD2.t0 B 0.276673f
C20 VDD2.n1 B 2.49024f
C21 VDD2.n2 B 4.03243f
C22 VDD2.t7 B 0.276673f
C23 VDD2.t5 B 0.276673f
C24 VDD2.n3 B 2.47434f
C25 VDD2.n4 B 3.51628f
C26 VDD2.t3 B 0.276673f
C27 VDD2.t2 B 0.276673f
C28 VDD2.n5 B 2.49019f
C29 VN.t7 B 2.20392f
C30 VN.n0 B 0.839054f
C31 VN.n1 B 0.018639f
C32 VN.n2 B 0.018142f
C33 VN.n3 B 0.018639f
C34 VN.t6 B 2.20392f
C35 VN.n4 B 0.770916f
C36 VN.n5 B 0.018639f
C37 VN.n6 B 0.027095f
C38 VN.n7 B 0.018639f
C39 VN.n8 B 0.01989f
C40 VN.t3 B 2.20392f
C41 VN.n9 B 0.827599f
C42 VN.t1 B 2.43179f
C43 VN.n10 B 0.792726f
C44 VN.n11 B 0.22042f
C45 VN.n12 B 0.018639f
C46 VN.n13 B 0.034565f
C47 VN.n14 B 0.034565f
C48 VN.n15 B 0.027095f
C49 VN.n16 B 0.018639f
C50 VN.n17 B 0.018639f
C51 VN.n18 B 0.018639f
C52 VN.n19 B 0.034565f
C53 VN.n20 B 0.034565f
C54 VN.n21 B 0.01989f
C55 VN.n22 B 0.018639f
C56 VN.n23 B 0.018639f
C57 VN.n24 B 0.032176f
C58 VN.n25 B 0.034565f
C59 VN.n26 B 0.033678f
C60 VN.n27 B 0.018639f
C61 VN.n28 B 0.018639f
C62 VN.n29 B 0.018639f
C63 VN.n30 B 0.036935f
C64 VN.n31 B 0.034565f
C65 VN.n32 B 0.024668f
C66 VN.n33 B 0.030079f
C67 VN.n34 B 0.048158f
C68 VN.t0 B 2.20392f
C69 VN.n35 B 0.839054f
C70 VN.n36 B 0.018639f
C71 VN.n37 B 0.018142f
C72 VN.n38 B 0.018639f
C73 VN.t2 B 2.20392f
C74 VN.n39 B 0.770916f
C75 VN.n40 B 0.018639f
C76 VN.n41 B 0.027095f
C77 VN.n42 B 0.018639f
C78 VN.n43 B 0.01989f
C79 VN.t5 B 2.43179f
C80 VN.t4 B 2.20392f
C81 VN.n44 B 0.827599f
C82 VN.n45 B 0.792726f
C83 VN.n46 B 0.22042f
C84 VN.n47 B 0.018639f
C85 VN.n48 B 0.034565f
C86 VN.n49 B 0.034565f
C87 VN.n50 B 0.027095f
C88 VN.n51 B 0.018639f
C89 VN.n52 B 0.018639f
C90 VN.n53 B 0.018639f
C91 VN.n54 B 0.034565f
C92 VN.n55 B 0.034565f
C93 VN.n56 B 0.01989f
C94 VN.n57 B 0.018639f
C95 VN.n58 B 0.018639f
C96 VN.n59 B 0.032176f
C97 VN.n60 B 0.034565f
C98 VN.n61 B 0.033678f
C99 VN.n62 B 0.018639f
C100 VN.n63 B 0.018639f
C101 VN.n64 B 0.018639f
C102 VN.n65 B 0.036935f
C103 VN.n66 B 0.034565f
C104 VN.n67 B 0.024668f
C105 VN.n68 B 0.030079f
C106 VN.n69 B 1.22456f
C107 VTAIL.t6 B 0.206661f
C108 VTAIL.t5 B 0.206661f
C109 VTAIL.n0 B 1.78353f
C110 VTAIL.n1 B 0.412485f
C111 VTAIL.t0 B 2.27373f
C112 VTAIL.n2 B 0.512432f
C113 VTAIL.t13 B 2.27373f
C114 VTAIL.n3 B 0.512432f
C115 VTAIL.t9 B 0.206661f
C116 VTAIL.t11 B 0.206661f
C117 VTAIL.n4 B 1.78353f
C118 VTAIL.n5 B 0.610896f
C119 VTAIL.t12 B 2.27373f
C120 VTAIL.n6 B 1.68236f
C121 VTAIL.t1 B 2.27373f
C122 VTAIL.n7 B 1.68235f
C123 VTAIL.t2 B 0.206661f
C124 VTAIL.t15 B 0.206661f
C125 VTAIL.n8 B 1.78353f
C126 VTAIL.n9 B 0.610898f
C127 VTAIL.t3 B 2.27373f
C128 VTAIL.n10 B 0.512426f
C129 VTAIL.t8 B 2.27373f
C130 VTAIL.n11 B 0.512426f
C131 VTAIL.t10 B 0.206661f
C132 VTAIL.t14 B 0.206661f
C133 VTAIL.n12 B 1.78353f
C134 VTAIL.n13 B 0.610898f
C135 VTAIL.t7 B 2.27373f
C136 VTAIL.n14 B 1.68236f
C137 VTAIL.t4 B 2.27373f
C138 VTAIL.n15 B 1.67861f
C139 VDD1.t0 B 0.282035f
C140 VDD1.t4 B 0.282035f
C141 VDD1.n0 B 2.53994f
C142 VDD1.t2 B 0.282035f
C143 VDD1.t1 B 0.282035f
C144 VDD1.n1 B 2.5385f
C145 VDD1.t5 B 0.282035f
C146 VDD1.t3 B 0.282035f
C147 VDD1.n2 B 2.5385f
C148 VDD1.n3 B 4.16696f
C149 VDD1.t6 B 0.282035f
C150 VDD1.t7 B 0.282035f
C151 VDD1.n4 B 2.52228f
C152 VDD1.n5 B 3.6186f
C153 VP.t1 B 2.24409f
C154 VP.n0 B 0.854345f
C155 VP.n1 B 0.018979f
C156 VP.n2 B 0.018473f
C157 VP.n3 B 0.018979f
C158 VP.t3 B 2.24409f
C159 VP.n4 B 0.784965f
C160 VP.n5 B 0.018979f
C161 VP.n6 B 0.027589f
C162 VP.n7 B 0.018979f
C163 VP.n8 B 0.020253f
C164 VP.n9 B 0.018979f
C165 VP.n10 B 0.018473f
C166 VP.n11 B 0.018979f
C167 VP.t2 B 2.24409f
C168 VP.n12 B 0.854345f
C169 VP.t7 B 2.24409f
C170 VP.n13 B 0.854345f
C171 VP.n14 B 0.018979f
C172 VP.n15 B 0.018473f
C173 VP.n16 B 0.018979f
C174 VP.t0 B 2.24409f
C175 VP.n17 B 0.784965f
C176 VP.n18 B 0.018979f
C177 VP.n19 B 0.027589f
C178 VP.n20 B 0.018979f
C179 VP.n21 B 0.020253f
C180 VP.t6 B 2.47611f
C181 VP.t4 B 2.24409f
C182 VP.n22 B 0.842682f
C183 VP.n23 B 0.807174f
C184 VP.n24 B 0.224438f
C185 VP.n25 B 0.018979f
C186 VP.n26 B 0.035195f
C187 VP.n27 B 0.035195f
C188 VP.n28 B 0.027589f
C189 VP.n29 B 0.018979f
C190 VP.n30 B 0.018979f
C191 VP.n31 B 0.018979f
C192 VP.n32 B 0.035195f
C193 VP.n33 B 0.035195f
C194 VP.n34 B 0.020253f
C195 VP.n35 B 0.018979f
C196 VP.n36 B 0.018979f
C197 VP.n37 B 0.032762f
C198 VP.n38 B 0.035195f
C199 VP.n39 B 0.034291f
C200 VP.n40 B 0.018979f
C201 VP.n41 B 0.018979f
C202 VP.n42 B 0.018979f
C203 VP.n43 B 0.037608f
C204 VP.n44 B 0.035195f
C205 VP.n45 B 0.025117f
C206 VP.n46 B 0.030627f
C207 VP.n47 B 1.23936f
C208 VP.n48 B 1.25178f
C209 VP.n49 B 0.030627f
C210 VP.n50 B 0.025117f
C211 VP.n51 B 0.035195f
C212 VP.n52 B 0.037608f
C213 VP.n53 B 0.018979f
C214 VP.n54 B 0.018979f
C215 VP.n55 B 0.018979f
C216 VP.n56 B 0.034291f
C217 VP.n57 B 0.035195f
C218 VP.t5 B 2.24409f
C219 VP.n58 B 0.784965f
C220 VP.n59 B 0.032762f
C221 VP.n60 B 0.018979f
C222 VP.n61 B 0.018979f
C223 VP.n62 B 0.018979f
C224 VP.n63 B 0.035195f
C225 VP.n64 B 0.035195f
C226 VP.n65 B 0.027589f
C227 VP.n66 B 0.018979f
C228 VP.n67 B 0.018979f
C229 VP.n68 B 0.018979f
C230 VP.n69 B 0.035195f
C231 VP.n70 B 0.035195f
C232 VP.n71 B 0.020253f
C233 VP.n72 B 0.018979f
C234 VP.n73 B 0.018979f
C235 VP.n74 B 0.032762f
C236 VP.n75 B 0.035195f
C237 VP.n76 B 0.034291f
C238 VP.n77 B 0.018979f
C239 VP.n78 B 0.018979f
C240 VP.n79 B 0.018979f
C241 VP.n80 B 0.037608f
C242 VP.n81 B 0.035195f
C243 VP.n82 B 0.025117f
C244 VP.n83 B 0.030627f
C245 VP.n84 B 0.049035f
.ends

