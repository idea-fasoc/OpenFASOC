* NGSPICE file created from diff_pair_sample_1097.ext - technology: sky130A

.subckt diff_pair_sample_1097 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t14 VP.t0 VDD1.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=2.25555 pd=14 as=2.25555 ps=14 w=13.67 l=1.31
X1 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=5.3313 pd=28.12 as=0 ps=0 w=13.67 l=1.31
X2 VTAIL.t6 VN.t0 VDD2.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=2.25555 pd=14 as=2.25555 ps=14 w=13.67 l=1.31
X3 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=5.3313 pd=28.12 as=0 ps=0 w=13.67 l=1.31
X4 VDD2.t6 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.25555 pd=14 as=2.25555 ps=14 w=13.67 l=1.31
X5 VDD1.t7 VP.t1 VTAIL.t13 B.t4 sky130_fd_pr__nfet_01v8 ad=2.25555 pd=14 as=5.3313 ps=28.12 w=13.67 l=1.31
X6 VTAIL.t15 VN.t2 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=2.25555 pd=14 as=2.25555 ps=14 w=13.67 l=1.31
X7 VDD2.t4 VN.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.25555 pd=14 as=5.3313 ps=28.12 w=13.67 l=1.31
X8 VDD2.t3 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.25555 pd=14 as=2.25555 ps=14 w=13.67 l=1.31
X9 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=5.3313 pd=28.12 as=0 ps=0 w=13.67 l=1.31
X10 VTAIL.t12 VP.t2 VDD1.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.3313 pd=28.12 as=2.25555 ps=14 w=13.67 l=1.31
X11 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.3313 pd=28.12 as=0 ps=0 w=13.67 l=1.31
X12 VDD1.t2 VP.t3 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=2.25555 pd=14 as=5.3313 ps=28.12 w=13.67 l=1.31
X13 VDD2.t2 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.25555 pd=14 as=5.3313 ps=28.12 w=13.67 l=1.31
X14 VTAIL.t2 VN.t6 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=5.3313 pd=28.12 as=2.25555 ps=14 w=13.67 l=1.31
X15 VTAIL.t10 VP.t4 VDD1.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=2.25555 pd=14 as=2.25555 ps=14 w=13.67 l=1.31
X16 VDD1.t5 VP.t5 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=2.25555 pd=14 as=2.25555 ps=14 w=13.67 l=1.31
X17 VTAIL.t5 VN.t7 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=5.3313 pd=28.12 as=2.25555 ps=14 w=13.67 l=1.31
X18 VDD1.t4 VP.t6 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=2.25555 pd=14 as=2.25555 ps=14 w=13.67 l=1.31
X19 VTAIL.t7 VP.t7 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=5.3313 pd=28.12 as=2.25555 ps=14 w=13.67 l=1.31
R0 VP.n11 VP.t7 279.003
R1 VP.n5 VP.t2 251.487
R2 VP.n29 VP.t5 251.487
R3 VP.n36 VP.t0 251.487
R4 VP.n43 VP.t1 251.487
R5 VP.n23 VP.t3 251.487
R6 VP.n16 VP.t4 251.487
R7 VP.n10 VP.t6 251.487
R8 VP.n25 VP.n5 175.492
R9 VP.n44 VP.n43 175.492
R10 VP.n24 VP.n23 175.492
R11 VP.n12 VP.n9 161.3
R12 VP.n14 VP.n13 161.3
R13 VP.n15 VP.n8 161.3
R14 VP.n18 VP.n17 161.3
R15 VP.n19 VP.n7 161.3
R16 VP.n21 VP.n20 161.3
R17 VP.n22 VP.n6 161.3
R18 VP.n42 VP.n0 161.3
R19 VP.n41 VP.n40 161.3
R20 VP.n39 VP.n1 161.3
R21 VP.n38 VP.n37 161.3
R22 VP.n35 VP.n2 161.3
R23 VP.n34 VP.n33 161.3
R24 VP.n32 VP.n3 161.3
R25 VP.n31 VP.n30 161.3
R26 VP.n28 VP.n4 161.3
R27 VP.n27 VP.n26 161.3
R28 VP.n11 VP.n10 62.0576
R29 VP.n35 VP.n34 56.5193
R30 VP.n15 VP.n14 56.5193
R31 VP.n30 VP.n28 51.1773
R32 VP.n41 VP.n1 51.1773
R33 VP.n21 VP.n7 51.1773
R34 VP.n25 VP.n24 46.0081
R35 VP.n28 VP.n27 29.8095
R36 VP.n42 VP.n41 29.8095
R37 VP.n22 VP.n21 29.8095
R38 VP.n12 VP.n11 27.6443
R39 VP.n34 VP.n3 24.4675
R40 VP.n37 VP.n35 24.4675
R41 VP.n17 VP.n15 24.4675
R42 VP.n14 VP.n9 24.4675
R43 VP.n30 VP.n29 21.0421
R44 VP.n36 VP.n1 21.0421
R45 VP.n16 VP.n7 21.0421
R46 VP.n27 VP.n5 10.2766
R47 VP.n43 VP.n42 10.2766
R48 VP.n23 VP.n22 10.2766
R49 VP.n29 VP.n3 3.42588
R50 VP.n37 VP.n36 3.42588
R51 VP.n17 VP.n16 3.42588
R52 VP.n10 VP.n9 3.42588
R53 VP.n13 VP.n12 0.189894
R54 VP.n13 VP.n8 0.189894
R55 VP.n18 VP.n8 0.189894
R56 VP.n19 VP.n18 0.189894
R57 VP.n20 VP.n19 0.189894
R58 VP.n20 VP.n6 0.189894
R59 VP.n24 VP.n6 0.189894
R60 VP.n26 VP.n25 0.189894
R61 VP.n26 VP.n4 0.189894
R62 VP.n31 VP.n4 0.189894
R63 VP.n32 VP.n31 0.189894
R64 VP.n33 VP.n32 0.189894
R65 VP.n33 VP.n2 0.189894
R66 VP.n38 VP.n2 0.189894
R67 VP.n39 VP.n38 0.189894
R68 VP.n40 VP.n39 0.189894
R69 VP.n40 VP.n0 0.189894
R70 VP.n44 VP.n0 0.189894
R71 VP VP.n44 0.0516364
R72 VDD1 VDD1.n0 63.9655
R73 VDD1.n3 VDD1.n2 63.8518
R74 VDD1.n3 VDD1.n1 63.8518
R75 VDD1.n5 VDD1.n4 63.2003
R76 VDD1.n5 VDD1.n3 42.4449
R77 VDD1.n4 VDD1.t1 1.44893
R78 VDD1.n4 VDD1.t2 1.44893
R79 VDD1.n0 VDD1.t3 1.44893
R80 VDD1.n0 VDD1.t4 1.44893
R81 VDD1.n2 VDD1.t0 1.44893
R82 VDD1.n2 VDD1.t7 1.44893
R83 VDD1.n1 VDD1.t6 1.44893
R84 VDD1.n1 VDD1.t5 1.44893
R85 VDD1 VDD1.n5 0.649207
R86 VTAIL.n11 VTAIL.t7 47.9701
R87 VTAIL.n10 VTAIL.t4 47.9701
R88 VTAIL.n7 VTAIL.t5 47.9701
R89 VTAIL.n15 VTAIL.t0 47.9699
R90 VTAIL.n2 VTAIL.t2 47.9699
R91 VTAIL.n3 VTAIL.t13 47.9699
R92 VTAIL.n6 VTAIL.t12 47.9699
R93 VTAIL.n14 VTAIL.t11 47.9699
R94 VTAIL.n13 VTAIL.n12 46.5217
R95 VTAIL.n9 VTAIL.n8 46.5217
R96 VTAIL.n1 VTAIL.n0 46.5215
R97 VTAIL.n5 VTAIL.n4 46.5215
R98 VTAIL.n15 VTAIL.n14 25.5652
R99 VTAIL.n7 VTAIL.n6 25.5652
R100 VTAIL.n0 VTAIL.t1 1.44893
R101 VTAIL.n0 VTAIL.t6 1.44893
R102 VTAIL.n4 VTAIL.t9 1.44893
R103 VTAIL.n4 VTAIL.t14 1.44893
R104 VTAIL.n12 VTAIL.t8 1.44893
R105 VTAIL.n12 VTAIL.t10 1.44893
R106 VTAIL.n8 VTAIL.t3 1.44893
R107 VTAIL.n8 VTAIL.t15 1.44893
R108 VTAIL.n9 VTAIL.n7 1.41429
R109 VTAIL.n10 VTAIL.n9 1.41429
R110 VTAIL.n13 VTAIL.n11 1.41429
R111 VTAIL.n14 VTAIL.n13 1.41429
R112 VTAIL.n6 VTAIL.n5 1.41429
R113 VTAIL.n5 VTAIL.n3 1.41429
R114 VTAIL.n2 VTAIL.n1 1.41429
R115 VTAIL VTAIL.n15 1.3561
R116 VTAIL.n11 VTAIL.n10 0.470328
R117 VTAIL.n3 VTAIL.n2 0.470328
R118 VTAIL VTAIL.n1 0.0586897
R119 B.n784 B.n783 585
R120 B.n785 B.n784 585
R121 B.n320 B.n113 585
R122 B.n319 B.n318 585
R123 B.n317 B.n316 585
R124 B.n315 B.n314 585
R125 B.n313 B.n312 585
R126 B.n311 B.n310 585
R127 B.n309 B.n308 585
R128 B.n307 B.n306 585
R129 B.n305 B.n304 585
R130 B.n303 B.n302 585
R131 B.n301 B.n300 585
R132 B.n299 B.n298 585
R133 B.n297 B.n296 585
R134 B.n295 B.n294 585
R135 B.n293 B.n292 585
R136 B.n291 B.n290 585
R137 B.n289 B.n288 585
R138 B.n287 B.n286 585
R139 B.n285 B.n284 585
R140 B.n283 B.n282 585
R141 B.n281 B.n280 585
R142 B.n279 B.n278 585
R143 B.n277 B.n276 585
R144 B.n275 B.n274 585
R145 B.n273 B.n272 585
R146 B.n271 B.n270 585
R147 B.n269 B.n268 585
R148 B.n267 B.n266 585
R149 B.n265 B.n264 585
R150 B.n263 B.n262 585
R151 B.n261 B.n260 585
R152 B.n259 B.n258 585
R153 B.n257 B.n256 585
R154 B.n255 B.n254 585
R155 B.n253 B.n252 585
R156 B.n251 B.n250 585
R157 B.n249 B.n248 585
R158 B.n247 B.n246 585
R159 B.n245 B.n244 585
R160 B.n243 B.n242 585
R161 B.n241 B.n240 585
R162 B.n239 B.n238 585
R163 B.n237 B.n236 585
R164 B.n235 B.n234 585
R165 B.n233 B.n232 585
R166 B.n231 B.n230 585
R167 B.n229 B.n228 585
R168 B.n227 B.n226 585
R169 B.n225 B.n224 585
R170 B.n223 B.n222 585
R171 B.n221 B.n220 585
R172 B.n219 B.n218 585
R173 B.n217 B.n216 585
R174 B.n215 B.n214 585
R175 B.n213 B.n212 585
R176 B.n210 B.n209 585
R177 B.n208 B.n207 585
R178 B.n206 B.n205 585
R179 B.n204 B.n203 585
R180 B.n202 B.n201 585
R181 B.n200 B.n199 585
R182 B.n198 B.n197 585
R183 B.n196 B.n195 585
R184 B.n194 B.n193 585
R185 B.n192 B.n191 585
R186 B.n190 B.n189 585
R187 B.n188 B.n187 585
R188 B.n186 B.n185 585
R189 B.n184 B.n183 585
R190 B.n182 B.n181 585
R191 B.n180 B.n179 585
R192 B.n178 B.n177 585
R193 B.n176 B.n175 585
R194 B.n174 B.n173 585
R195 B.n172 B.n171 585
R196 B.n170 B.n169 585
R197 B.n168 B.n167 585
R198 B.n166 B.n165 585
R199 B.n164 B.n163 585
R200 B.n162 B.n161 585
R201 B.n160 B.n159 585
R202 B.n158 B.n157 585
R203 B.n156 B.n155 585
R204 B.n154 B.n153 585
R205 B.n152 B.n151 585
R206 B.n150 B.n149 585
R207 B.n148 B.n147 585
R208 B.n146 B.n145 585
R209 B.n144 B.n143 585
R210 B.n142 B.n141 585
R211 B.n140 B.n139 585
R212 B.n138 B.n137 585
R213 B.n136 B.n135 585
R214 B.n134 B.n133 585
R215 B.n132 B.n131 585
R216 B.n130 B.n129 585
R217 B.n128 B.n127 585
R218 B.n126 B.n125 585
R219 B.n124 B.n123 585
R220 B.n122 B.n121 585
R221 B.n120 B.n119 585
R222 B.n60 B.n59 585
R223 B.n782 B.n61 585
R224 B.n786 B.n61 585
R225 B.n781 B.n780 585
R226 B.n780 B.n57 585
R227 B.n779 B.n56 585
R228 B.n792 B.n56 585
R229 B.n778 B.n55 585
R230 B.n793 B.n55 585
R231 B.n777 B.n54 585
R232 B.n794 B.n54 585
R233 B.n776 B.n775 585
R234 B.n775 B.n53 585
R235 B.n774 B.n49 585
R236 B.n800 B.n49 585
R237 B.n773 B.n48 585
R238 B.n801 B.n48 585
R239 B.n772 B.n47 585
R240 B.n802 B.n47 585
R241 B.n771 B.n770 585
R242 B.n770 B.n43 585
R243 B.n769 B.n42 585
R244 B.n808 B.n42 585
R245 B.n768 B.n41 585
R246 B.n809 B.n41 585
R247 B.n767 B.n40 585
R248 B.n810 B.n40 585
R249 B.n766 B.n765 585
R250 B.n765 B.n39 585
R251 B.n764 B.n35 585
R252 B.n816 B.n35 585
R253 B.n763 B.n34 585
R254 B.n817 B.n34 585
R255 B.n762 B.n33 585
R256 B.n818 B.n33 585
R257 B.n761 B.n760 585
R258 B.n760 B.n29 585
R259 B.n759 B.n28 585
R260 B.n824 B.n28 585
R261 B.n758 B.n27 585
R262 B.n825 B.n27 585
R263 B.n757 B.n26 585
R264 B.n826 B.n26 585
R265 B.n756 B.n755 585
R266 B.n755 B.n22 585
R267 B.n754 B.n21 585
R268 B.n832 B.n21 585
R269 B.n753 B.n20 585
R270 B.n833 B.n20 585
R271 B.n752 B.n19 585
R272 B.n834 B.n19 585
R273 B.n751 B.n750 585
R274 B.n750 B.n15 585
R275 B.n749 B.n14 585
R276 B.n840 B.n14 585
R277 B.n748 B.n13 585
R278 B.n841 B.n13 585
R279 B.n747 B.n12 585
R280 B.n842 B.n12 585
R281 B.n746 B.n745 585
R282 B.n745 B.n8 585
R283 B.n744 B.n7 585
R284 B.n848 B.n7 585
R285 B.n743 B.n6 585
R286 B.n849 B.n6 585
R287 B.n742 B.n5 585
R288 B.n850 B.n5 585
R289 B.n741 B.n740 585
R290 B.n740 B.n4 585
R291 B.n739 B.n321 585
R292 B.n739 B.n738 585
R293 B.n729 B.n322 585
R294 B.n323 B.n322 585
R295 B.n731 B.n730 585
R296 B.n732 B.n731 585
R297 B.n728 B.n327 585
R298 B.n331 B.n327 585
R299 B.n727 B.n726 585
R300 B.n726 B.n725 585
R301 B.n329 B.n328 585
R302 B.n330 B.n329 585
R303 B.n718 B.n717 585
R304 B.n719 B.n718 585
R305 B.n716 B.n335 585
R306 B.n339 B.n335 585
R307 B.n715 B.n714 585
R308 B.n714 B.n713 585
R309 B.n337 B.n336 585
R310 B.n338 B.n337 585
R311 B.n706 B.n705 585
R312 B.n707 B.n706 585
R313 B.n704 B.n344 585
R314 B.n344 B.n343 585
R315 B.n703 B.n702 585
R316 B.n702 B.n701 585
R317 B.n346 B.n345 585
R318 B.n347 B.n346 585
R319 B.n694 B.n693 585
R320 B.n695 B.n694 585
R321 B.n692 B.n352 585
R322 B.n352 B.n351 585
R323 B.n691 B.n690 585
R324 B.n690 B.n689 585
R325 B.n354 B.n353 585
R326 B.n682 B.n354 585
R327 B.n681 B.n680 585
R328 B.n683 B.n681 585
R329 B.n679 B.n359 585
R330 B.n359 B.n358 585
R331 B.n678 B.n677 585
R332 B.n677 B.n676 585
R333 B.n361 B.n360 585
R334 B.n362 B.n361 585
R335 B.n669 B.n668 585
R336 B.n670 B.n669 585
R337 B.n667 B.n367 585
R338 B.n367 B.n366 585
R339 B.n666 B.n665 585
R340 B.n665 B.n664 585
R341 B.n369 B.n368 585
R342 B.n657 B.n369 585
R343 B.n656 B.n655 585
R344 B.n658 B.n656 585
R345 B.n654 B.n374 585
R346 B.n374 B.n373 585
R347 B.n653 B.n652 585
R348 B.n652 B.n651 585
R349 B.n376 B.n375 585
R350 B.n377 B.n376 585
R351 B.n644 B.n643 585
R352 B.n645 B.n644 585
R353 B.n380 B.n379 585
R354 B.n437 B.n436 585
R355 B.n438 B.n434 585
R356 B.n434 B.n381 585
R357 B.n440 B.n439 585
R358 B.n442 B.n433 585
R359 B.n445 B.n444 585
R360 B.n446 B.n432 585
R361 B.n448 B.n447 585
R362 B.n450 B.n431 585
R363 B.n453 B.n452 585
R364 B.n454 B.n430 585
R365 B.n456 B.n455 585
R366 B.n458 B.n429 585
R367 B.n461 B.n460 585
R368 B.n462 B.n428 585
R369 B.n464 B.n463 585
R370 B.n466 B.n427 585
R371 B.n469 B.n468 585
R372 B.n470 B.n426 585
R373 B.n472 B.n471 585
R374 B.n474 B.n425 585
R375 B.n477 B.n476 585
R376 B.n478 B.n424 585
R377 B.n480 B.n479 585
R378 B.n482 B.n423 585
R379 B.n485 B.n484 585
R380 B.n486 B.n422 585
R381 B.n488 B.n487 585
R382 B.n490 B.n421 585
R383 B.n493 B.n492 585
R384 B.n494 B.n420 585
R385 B.n496 B.n495 585
R386 B.n498 B.n419 585
R387 B.n501 B.n500 585
R388 B.n502 B.n418 585
R389 B.n504 B.n503 585
R390 B.n506 B.n417 585
R391 B.n509 B.n508 585
R392 B.n510 B.n416 585
R393 B.n512 B.n511 585
R394 B.n514 B.n415 585
R395 B.n517 B.n516 585
R396 B.n518 B.n414 585
R397 B.n520 B.n519 585
R398 B.n522 B.n413 585
R399 B.n525 B.n524 585
R400 B.n526 B.n410 585
R401 B.n529 B.n528 585
R402 B.n531 B.n409 585
R403 B.n534 B.n533 585
R404 B.n535 B.n408 585
R405 B.n537 B.n536 585
R406 B.n539 B.n407 585
R407 B.n542 B.n541 585
R408 B.n543 B.n406 585
R409 B.n548 B.n547 585
R410 B.n550 B.n405 585
R411 B.n553 B.n552 585
R412 B.n554 B.n404 585
R413 B.n556 B.n555 585
R414 B.n558 B.n403 585
R415 B.n561 B.n560 585
R416 B.n562 B.n402 585
R417 B.n564 B.n563 585
R418 B.n566 B.n401 585
R419 B.n569 B.n568 585
R420 B.n570 B.n400 585
R421 B.n572 B.n571 585
R422 B.n574 B.n399 585
R423 B.n577 B.n576 585
R424 B.n578 B.n398 585
R425 B.n580 B.n579 585
R426 B.n582 B.n397 585
R427 B.n585 B.n584 585
R428 B.n586 B.n396 585
R429 B.n588 B.n587 585
R430 B.n590 B.n395 585
R431 B.n593 B.n592 585
R432 B.n594 B.n394 585
R433 B.n596 B.n595 585
R434 B.n598 B.n393 585
R435 B.n601 B.n600 585
R436 B.n602 B.n392 585
R437 B.n604 B.n603 585
R438 B.n606 B.n391 585
R439 B.n609 B.n608 585
R440 B.n610 B.n390 585
R441 B.n612 B.n611 585
R442 B.n614 B.n389 585
R443 B.n617 B.n616 585
R444 B.n618 B.n388 585
R445 B.n620 B.n619 585
R446 B.n622 B.n387 585
R447 B.n625 B.n624 585
R448 B.n626 B.n386 585
R449 B.n628 B.n627 585
R450 B.n630 B.n385 585
R451 B.n633 B.n632 585
R452 B.n634 B.n384 585
R453 B.n636 B.n635 585
R454 B.n638 B.n383 585
R455 B.n641 B.n640 585
R456 B.n642 B.n382 585
R457 B.n647 B.n646 585
R458 B.n646 B.n645 585
R459 B.n648 B.n378 585
R460 B.n378 B.n377 585
R461 B.n650 B.n649 585
R462 B.n651 B.n650 585
R463 B.n372 B.n371 585
R464 B.n373 B.n372 585
R465 B.n660 B.n659 585
R466 B.n659 B.n658 585
R467 B.n661 B.n370 585
R468 B.n657 B.n370 585
R469 B.n663 B.n662 585
R470 B.n664 B.n663 585
R471 B.n365 B.n364 585
R472 B.n366 B.n365 585
R473 B.n672 B.n671 585
R474 B.n671 B.n670 585
R475 B.n673 B.n363 585
R476 B.n363 B.n362 585
R477 B.n675 B.n674 585
R478 B.n676 B.n675 585
R479 B.n357 B.n356 585
R480 B.n358 B.n357 585
R481 B.n685 B.n684 585
R482 B.n684 B.n683 585
R483 B.n686 B.n355 585
R484 B.n682 B.n355 585
R485 B.n688 B.n687 585
R486 B.n689 B.n688 585
R487 B.n350 B.n349 585
R488 B.n351 B.n350 585
R489 B.n697 B.n696 585
R490 B.n696 B.n695 585
R491 B.n698 B.n348 585
R492 B.n348 B.n347 585
R493 B.n700 B.n699 585
R494 B.n701 B.n700 585
R495 B.n342 B.n341 585
R496 B.n343 B.n342 585
R497 B.n709 B.n708 585
R498 B.n708 B.n707 585
R499 B.n710 B.n340 585
R500 B.n340 B.n338 585
R501 B.n712 B.n711 585
R502 B.n713 B.n712 585
R503 B.n334 B.n333 585
R504 B.n339 B.n334 585
R505 B.n721 B.n720 585
R506 B.n720 B.n719 585
R507 B.n722 B.n332 585
R508 B.n332 B.n330 585
R509 B.n724 B.n723 585
R510 B.n725 B.n724 585
R511 B.n326 B.n325 585
R512 B.n331 B.n326 585
R513 B.n734 B.n733 585
R514 B.n733 B.n732 585
R515 B.n735 B.n324 585
R516 B.n324 B.n323 585
R517 B.n737 B.n736 585
R518 B.n738 B.n737 585
R519 B.n2 B.n0 585
R520 B.n4 B.n2 585
R521 B.n3 B.n1 585
R522 B.n849 B.n3 585
R523 B.n847 B.n846 585
R524 B.n848 B.n847 585
R525 B.n845 B.n9 585
R526 B.n9 B.n8 585
R527 B.n844 B.n843 585
R528 B.n843 B.n842 585
R529 B.n11 B.n10 585
R530 B.n841 B.n11 585
R531 B.n839 B.n838 585
R532 B.n840 B.n839 585
R533 B.n837 B.n16 585
R534 B.n16 B.n15 585
R535 B.n836 B.n835 585
R536 B.n835 B.n834 585
R537 B.n18 B.n17 585
R538 B.n833 B.n18 585
R539 B.n831 B.n830 585
R540 B.n832 B.n831 585
R541 B.n829 B.n23 585
R542 B.n23 B.n22 585
R543 B.n828 B.n827 585
R544 B.n827 B.n826 585
R545 B.n25 B.n24 585
R546 B.n825 B.n25 585
R547 B.n823 B.n822 585
R548 B.n824 B.n823 585
R549 B.n821 B.n30 585
R550 B.n30 B.n29 585
R551 B.n820 B.n819 585
R552 B.n819 B.n818 585
R553 B.n32 B.n31 585
R554 B.n817 B.n32 585
R555 B.n815 B.n814 585
R556 B.n816 B.n815 585
R557 B.n813 B.n36 585
R558 B.n39 B.n36 585
R559 B.n812 B.n811 585
R560 B.n811 B.n810 585
R561 B.n38 B.n37 585
R562 B.n809 B.n38 585
R563 B.n807 B.n806 585
R564 B.n808 B.n807 585
R565 B.n805 B.n44 585
R566 B.n44 B.n43 585
R567 B.n804 B.n803 585
R568 B.n803 B.n802 585
R569 B.n46 B.n45 585
R570 B.n801 B.n46 585
R571 B.n799 B.n798 585
R572 B.n800 B.n799 585
R573 B.n797 B.n50 585
R574 B.n53 B.n50 585
R575 B.n796 B.n795 585
R576 B.n795 B.n794 585
R577 B.n52 B.n51 585
R578 B.n793 B.n52 585
R579 B.n791 B.n790 585
R580 B.n792 B.n791 585
R581 B.n789 B.n58 585
R582 B.n58 B.n57 585
R583 B.n788 B.n787 585
R584 B.n787 B.n786 585
R585 B.n852 B.n851 585
R586 B.n851 B.n850 585
R587 B.n646 B.n380 506.916
R588 B.n787 B.n60 506.916
R589 B.n644 B.n382 506.916
R590 B.n784 B.n61 506.916
R591 B.n544 B.t19 456.142
R592 B.n411 B.t15 456.142
R593 B.n117 B.t12 456.142
R594 B.n114 B.t8 456.142
R595 B.n785 B.n112 256.663
R596 B.n785 B.n111 256.663
R597 B.n785 B.n110 256.663
R598 B.n785 B.n109 256.663
R599 B.n785 B.n108 256.663
R600 B.n785 B.n107 256.663
R601 B.n785 B.n106 256.663
R602 B.n785 B.n105 256.663
R603 B.n785 B.n104 256.663
R604 B.n785 B.n103 256.663
R605 B.n785 B.n102 256.663
R606 B.n785 B.n101 256.663
R607 B.n785 B.n100 256.663
R608 B.n785 B.n99 256.663
R609 B.n785 B.n98 256.663
R610 B.n785 B.n97 256.663
R611 B.n785 B.n96 256.663
R612 B.n785 B.n95 256.663
R613 B.n785 B.n94 256.663
R614 B.n785 B.n93 256.663
R615 B.n785 B.n92 256.663
R616 B.n785 B.n91 256.663
R617 B.n785 B.n90 256.663
R618 B.n785 B.n89 256.663
R619 B.n785 B.n88 256.663
R620 B.n785 B.n87 256.663
R621 B.n785 B.n86 256.663
R622 B.n785 B.n85 256.663
R623 B.n785 B.n84 256.663
R624 B.n785 B.n83 256.663
R625 B.n785 B.n82 256.663
R626 B.n785 B.n81 256.663
R627 B.n785 B.n80 256.663
R628 B.n785 B.n79 256.663
R629 B.n785 B.n78 256.663
R630 B.n785 B.n77 256.663
R631 B.n785 B.n76 256.663
R632 B.n785 B.n75 256.663
R633 B.n785 B.n74 256.663
R634 B.n785 B.n73 256.663
R635 B.n785 B.n72 256.663
R636 B.n785 B.n71 256.663
R637 B.n785 B.n70 256.663
R638 B.n785 B.n69 256.663
R639 B.n785 B.n68 256.663
R640 B.n785 B.n67 256.663
R641 B.n785 B.n66 256.663
R642 B.n785 B.n65 256.663
R643 B.n785 B.n64 256.663
R644 B.n785 B.n63 256.663
R645 B.n785 B.n62 256.663
R646 B.n435 B.n381 256.663
R647 B.n441 B.n381 256.663
R648 B.n443 B.n381 256.663
R649 B.n449 B.n381 256.663
R650 B.n451 B.n381 256.663
R651 B.n457 B.n381 256.663
R652 B.n459 B.n381 256.663
R653 B.n465 B.n381 256.663
R654 B.n467 B.n381 256.663
R655 B.n473 B.n381 256.663
R656 B.n475 B.n381 256.663
R657 B.n481 B.n381 256.663
R658 B.n483 B.n381 256.663
R659 B.n489 B.n381 256.663
R660 B.n491 B.n381 256.663
R661 B.n497 B.n381 256.663
R662 B.n499 B.n381 256.663
R663 B.n505 B.n381 256.663
R664 B.n507 B.n381 256.663
R665 B.n513 B.n381 256.663
R666 B.n515 B.n381 256.663
R667 B.n521 B.n381 256.663
R668 B.n523 B.n381 256.663
R669 B.n530 B.n381 256.663
R670 B.n532 B.n381 256.663
R671 B.n538 B.n381 256.663
R672 B.n540 B.n381 256.663
R673 B.n549 B.n381 256.663
R674 B.n551 B.n381 256.663
R675 B.n557 B.n381 256.663
R676 B.n559 B.n381 256.663
R677 B.n565 B.n381 256.663
R678 B.n567 B.n381 256.663
R679 B.n573 B.n381 256.663
R680 B.n575 B.n381 256.663
R681 B.n581 B.n381 256.663
R682 B.n583 B.n381 256.663
R683 B.n589 B.n381 256.663
R684 B.n591 B.n381 256.663
R685 B.n597 B.n381 256.663
R686 B.n599 B.n381 256.663
R687 B.n605 B.n381 256.663
R688 B.n607 B.n381 256.663
R689 B.n613 B.n381 256.663
R690 B.n615 B.n381 256.663
R691 B.n621 B.n381 256.663
R692 B.n623 B.n381 256.663
R693 B.n629 B.n381 256.663
R694 B.n631 B.n381 256.663
R695 B.n637 B.n381 256.663
R696 B.n639 B.n381 256.663
R697 B.n646 B.n378 163.367
R698 B.n650 B.n378 163.367
R699 B.n650 B.n372 163.367
R700 B.n659 B.n372 163.367
R701 B.n659 B.n370 163.367
R702 B.n663 B.n370 163.367
R703 B.n663 B.n365 163.367
R704 B.n671 B.n365 163.367
R705 B.n671 B.n363 163.367
R706 B.n675 B.n363 163.367
R707 B.n675 B.n357 163.367
R708 B.n684 B.n357 163.367
R709 B.n684 B.n355 163.367
R710 B.n688 B.n355 163.367
R711 B.n688 B.n350 163.367
R712 B.n696 B.n350 163.367
R713 B.n696 B.n348 163.367
R714 B.n700 B.n348 163.367
R715 B.n700 B.n342 163.367
R716 B.n708 B.n342 163.367
R717 B.n708 B.n340 163.367
R718 B.n712 B.n340 163.367
R719 B.n712 B.n334 163.367
R720 B.n720 B.n334 163.367
R721 B.n720 B.n332 163.367
R722 B.n724 B.n332 163.367
R723 B.n724 B.n326 163.367
R724 B.n733 B.n326 163.367
R725 B.n733 B.n324 163.367
R726 B.n737 B.n324 163.367
R727 B.n737 B.n2 163.367
R728 B.n851 B.n2 163.367
R729 B.n851 B.n3 163.367
R730 B.n847 B.n3 163.367
R731 B.n847 B.n9 163.367
R732 B.n843 B.n9 163.367
R733 B.n843 B.n11 163.367
R734 B.n839 B.n11 163.367
R735 B.n839 B.n16 163.367
R736 B.n835 B.n16 163.367
R737 B.n835 B.n18 163.367
R738 B.n831 B.n18 163.367
R739 B.n831 B.n23 163.367
R740 B.n827 B.n23 163.367
R741 B.n827 B.n25 163.367
R742 B.n823 B.n25 163.367
R743 B.n823 B.n30 163.367
R744 B.n819 B.n30 163.367
R745 B.n819 B.n32 163.367
R746 B.n815 B.n32 163.367
R747 B.n815 B.n36 163.367
R748 B.n811 B.n36 163.367
R749 B.n811 B.n38 163.367
R750 B.n807 B.n38 163.367
R751 B.n807 B.n44 163.367
R752 B.n803 B.n44 163.367
R753 B.n803 B.n46 163.367
R754 B.n799 B.n46 163.367
R755 B.n799 B.n50 163.367
R756 B.n795 B.n50 163.367
R757 B.n795 B.n52 163.367
R758 B.n791 B.n52 163.367
R759 B.n791 B.n58 163.367
R760 B.n787 B.n58 163.367
R761 B.n436 B.n434 163.367
R762 B.n440 B.n434 163.367
R763 B.n444 B.n442 163.367
R764 B.n448 B.n432 163.367
R765 B.n452 B.n450 163.367
R766 B.n456 B.n430 163.367
R767 B.n460 B.n458 163.367
R768 B.n464 B.n428 163.367
R769 B.n468 B.n466 163.367
R770 B.n472 B.n426 163.367
R771 B.n476 B.n474 163.367
R772 B.n480 B.n424 163.367
R773 B.n484 B.n482 163.367
R774 B.n488 B.n422 163.367
R775 B.n492 B.n490 163.367
R776 B.n496 B.n420 163.367
R777 B.n500 B.n498 163.367
R778 B.n504 B.n418 163.367
R779 B.n508 B.n506 163.367
R780 B.n512 B.n416 163.367
R781 B.n516 B.n514 163.367
R782 B.n520 B.n414 163.367
R783 B.n524 B.n522 163.367
R784 B.n529 B.n410 163.367
R785 B.n533 B.n531 163.367
R786 B.n537 B.n408 163.367
R787 B.n541 B.n539 163.367
R788 B.n548 B.n406 163.367
R789 B.n552 B.n550 163.367
R790 B.n556 B.n404 163.367
R791 B.n560 B.n558 163.367
R792 B.n564 B.n402 163.367
R793 B.n568 B.n566 163.367
R794 B.n572 B.n400 163.367
R795 B.n576 B.n574 163.367
R796 B.n580 B.n398 163.367
R797 B.n584 B.n582 163.367
R798 B.n588 B.n396 163.367
R799 B.n592 B.n590 163.367
R800 B.n596 B.n394 163.367
R801 B.n600 B.n598 163.367
R802 B.n604 B.n392 163.367
R803 B.n608 B.n606 163.367
R804 B.n612 B.n390 163.367
R805 B.n616 B.n614 163.367
R806 B.n620 B.n388 163.367
R807 B.n624 B.n622 163.367
R808 B.n628 B.n386 163.367
R809 B.n632 B.n630 163.367
R810 B.n636 B.n384 163.367
R811 B.n640 B.n638 163.367
R812 B.n644 B.n376 163.367
R813 B.n652 B.n376 163.367
R814 B.n652 B.n374 163.367
R815 B.n656 B.n374 163.367
R816 B.n656 B.n369 163.367
R817 B.n665 B.n369 163.367
R818 B.n665 B.n367 163.367
R819 B.n669 B.n367 163.367
R820 B.n669 B.n361 163.367
R821 B.n677 B.n361 163.367
R822 B.n677 B.n359 163.367
R823 B.n681 B.n359 163.367
R824 B.n681 B.n354 163.367
R825 B.n690 B.n354 163.367
R826 B.n690 B.n352 163.367
R827 B.n694 B.n352 163.367
R828 B.n694 B.n346 163.367
R829 B.n702 B.n346 163.367
R830 B.n702 B.n344 163.367
R831 B.n706 B.n344 163.367
R832 B.n706 B.n337 163.367
R833 B.n714 B.n337 163.367
R834 B.n714 B.n335 163.367
R835 B.n718 B.n335 163.367
R836 B.n718 B.n329 163.367
R837 B.n726 B.n329 163.367
R838 B.n726 B.n327 163.367
R839 B.n731 B.n327 163.367
R840 B.n731 B.n322 163.367
R841 B.n739 B.n322 163.367
R842 B.n740 B.n739 163.367
R843 B.n740 B.n5 163.367
R844 B.n6 B.n5 163.367
R845 B.n7 B.n6 163.367
R846 B.n745 B.n7 163.367
R847 B.n745 B.n12 163.367
R848 B.n13 B.n12 163.367
R849 B.n14 B.n13 163.367
R850 B.n750 B.n14 163.367
R851 B.n750 B.n19 163.367
R852 B.n20 B.n19 163.367
R853 B.n21 B.n20 163.367
R854 B.n755 B.n21 163.367
R855 B.n755 B.n26 163.367
R856 B.n27 B.n26 163.367
R857 B.n28 B.n27 163.367
R858 B.n760 B.n28 163.367
R859 B.n760 B.n33 163.367
R860 B.n34 B.n33 163.367
R861 B.n35 B.n34 163.367
R862 B.n765 B.n35 163.367
R863 B.n765 B.n40 163.367
R864 B.n41 B.n40 163.367
R865 B.n42 B.n41 163.367
R866 B.n770 B.n42 163.367
R867 B.n770 B.n47 163.367
R868 B.n48 B.n47 163.367
R869 B.n49 B.n48 163.367
R870 B.n775 B.n49 163.367
R871 B.n775 B.n54 163.367
R872 B.n55 B.n54 163.367
R873 B.n56 B.n55 163.367
R874 B.n780 B.n56 163.367
R875 B.n780 B.n61 163.367
R876 B.n121 B.n120 163.367
R877 B.n125 B.n124 163.367
R878 B.n129 B.n128 163.367
R879 B.n133 B.n132 163.367
R880 B.n137 B.n136 163.367
R881 B.n141 B.n140 163.367
R882 B.n145 B.n144 163.367
R883 B.n149 B.n148 163.367
R884 B.n153 B.n152 163.367
R885 B.n157 B.n156 163.367
R886 B.n161 B.n160 163.367
R887 B.n165 B.n164 163.367
R888 B.n169 B.n168 163.367
R889 B.n173 B.n172 163.367
R890 B.n177 B.n176 163.367
R891 B.n181 B.n180 163.367
R892 B.n185 B.n184 163.367
R893 B.n189 B.n188 163.367
R894 B.n193 B.n192 163.367
R895 B.n197 B.n196 163.367
R896 B.n201 B.n200 163.367
R897 B.n205 B.n204 163.367
R898 B.n209 B.n208 163.367
R899 B.n214 B.n213 163.367
R900 B.n218 B.n217 163.367
R901 B.n222 B.n221 163.367
R902 B.n226 B.n225 163.367
R903 B.n230 B.n229 163.367
R904 B.n234 B.n233 163.367
R905 B.n238 B.n237 163.367
R906 B.n242 B.n241 163.367
R907 B.n246 B.n245 163.367
R908 B.n250 B.n249 163.367
R909 B.n254 B.n253 163.367
R910 B.n258 B.n257 163.367
R911 B.n262 B.n261 163.367
R912 B.n266 B.n265 163.367
R913 B.n270 B.n269 163.367
R914 B.n274 B.n273 163.367
R915 B.n278 B.n277 163.367
R916 B.n282 B.n281 163.367
R917 B.n286 B.n285 163.367
R918 B.n290 B.n289 163.367
R919 B.n294 B.n293 163.367
R920 B.n298 B.n297 163.367
R921 B.n302 B.n301 163.367
R922 B.n306 B.n305 163.367
R923 B.n310 B.n309 163.367
R924 B.n314 B.n313 163.367
R925 B.n318 B.n317 163.367
R926 B.n784 B.n113 163.367
R927 B.n544 B.t21 100.754
R928 B.n114 B.t10 100.754
R929 B.n411 B.t18 100.737
R930 B.n117 B.t13 100.737
R931 B.n645 B.n381 80.7078
R932 B.n786 B.n785 80.7078
R933 B.n435 B.n380 71.676
R934 B.n441 B.n440 71.676
R935 B.n444 B.n443 71.676
R936 B.n449 B.n448 71.676
R937 B.n452 B.n451 71.676
R938 B.n457 B.n456 71.676
R939 B.n460 B.n459 71.676
R940 B.n465 B.n464 71.676
R941 B.n468 B.n467 71.676
R942 B.n473 B.n472 71.676
R943 B.n476 B.n475 71.676
R944 B.n481 B.n480 71.676
R945 B.n484 B.n483 71.676
R946 B.n489 B.n488 71.676
R947 B.n492 B.n491 71.676
R948 B.n497 B.n496 71.676
R949 B.n500 B.n499 71.676
R950 B.n505 B.n504 71.676
R951 B.n508 B.n507 71.676
R952 B.n513 B.n512 71.676
R953 B.n516 B.n515 71.676
R954 B.n521 B.n520 71.676
R955 B.n524 B.n523 71.676
R956 B.n530 B.n529 71.676
R957 B.n533 B.n532 71.676
R958 B.n538 B.n537 71.676
R959 B.n541 B.n540 71.676
R960 B.n549 B.n548 71.676
R961 B.n552 B.n551 71.676
R962 B.n557 B.n556 71.676
R963 B.n560 B.n559 71.676
R964 B.n565 B.n564 71.676
R965 B.n568 B.n567 71.676
R966 B.n573 B.n572 71.676
R967 B.n576 B.n575 71.676
R968 B.n581 B.n580 71.676
R969 B.n584 B.n583 71.676
R970 B.n589 B.n588 71.676
R971 B.n592 B.n591 71.676
R972 B.n597 B.n596 71.676
R973 B.n600 B.n599 71.676
R974 B.n605 B.n604 71.676
R975 B.n608 B.n607 71.676
R976 B.n613 B.n612 71.676
R977 B.n616 B.n615 71.676
R978 B.n621 B.n620 71.676
R979 B.n624 B.n623 71.676
R980 B.n629 B.n628 71.676
R981 B.n632 B.n631 71.676
R982 B.n637 B.n636 71.676
R983 B.n640 B.n639 71.676
R984 B.n62 B.n60 71.676
R985 B.n121 B.n63 71.676
R986 B.n125 B.n64 71.676
R987 B.n129 B.n65 71.676
R988 B.n133 B.n66 71.676
R989 B.n137 B.n67 71.676
R990 B.n141 B.n68 71.676
R991 B.n145 B.n69 71.676
R992 B.n149 B.n70 71.676
R993 B.n153 B.n71 71.676
R994 B.n157 B.n72 71.676
R995 B.n161 B.n73 71.676
R996 B.n165 B.n74 71.676
R997 B.n169 B.n75 71.676
R998 B.n173 B.n76 71.676
R999 B.n177 B.n77 71.676
R1000 B.n181 B.n78 71.676
R1001 B.n185 B.n79 71.676
R1002 B.n189 B.n80 71.676
R1003 B.n193 B.n81 71.676
R1004 B.n197 B.n82 71.676
R1005 B.n201 B.n83 71.676
R1006 B.n205 B.n84 71.676
R1007 B.n209 B.n85 71.676
R1008 B.n214 B.n86 71.676
R1009 B.n218 B.n87 71.676
R1010 B.n222 B.n88 71.676
R1011 B.n226 B.n89 71.676
R1012 B.n230 B.n90 71.676
R1013 B.n234 B.n91 71.676
R1014 B.n238 B.n92 71.676
R1015 B.n242 B.n93 71.676
R1016 B.n246 B.n94 71.676
R1017 B.n250 B.n95 71.676
R1018 B.n254 B.n96 71.676
R1019 B.n258 B.n97 71.676
R1020 B.n262 B.n98 71.676
R1021 B.n266 B.n99 71.676
R1022 B.n270 B.n100 71.676
R1023 B.n274 B.n101 71.676
R1024 B.n278 B.n102 71.676
R1025 B.n282 B.n103 71.676
R1026 B.n286 B.n104 71.676
R1027 B.n290 B.n105 71.676
R1028 B.n294 B.n106 71.676
R1029 B.n298 B.n107 71.676
R1030 B.n302 B.n108 71.676
R1031 B.n306 B.n109 71.676
R1032 B.n310 B.n110 71.676
R1033 B.n314 B.n111 71.676
R1034 B.n318 B.n112 71.676
R1035 B.n113 B.n112 71.676
R1036 B.n317 B.n111 71.676
R1037 B.n313 B.n110 71.676
R1038 B.n309 B.n109 71.676
R1039 B.n305 B.n108 71.676
R1040 B.n301 B.n107 71.676
R1041 B.n297 B.n106 71.676
R1042 B.n293 B.n105 71.676
R1043 B.n289 B.n104 71.676
R1044 B.n285 B.n103 71.676
R1045 B.n281 B.n102 71.676
R1046 B.n277 B.n101 71.676
R1047 B.n273 B.n100 71.676
R1048 B.n269 B.n99 71.676
R1049 B.n265 B.n98 71.676
R1050 B.n261 B.n97 71.676
R1051 B.n257 B.n96 71.676
R1052 B.n253 B.n95 71.676
R1053 B.n249 B.n94 71.676
R1054 B.n245 B.n93 71.676
R1055 B.n241 B.n92 71.676
R1056 B.n237 B.n91 71.676
R1057 B.n233 B.n90 71.676
R1058 B.n229 B.n89 71.676
R1059 B.n225 B.n88 71.676
R1060 B.n221 B.n87 71.676
R1061 B.n217 B.n86 71.676
R1062 B.n213 B.n85 71.676
R1063 B.n208 B.n84 71.676
R1064 B.n204 B.n83 71.676
R1065 B.n200 B.n82 71.676
R1066 B.n196 B.n81 71.676
R1067 B.n192 B.n80 71.676
R1068 B.n188 B.n79 71.676
R1069 B.n184 B.n78 71.676
R1070 B.n180 B.n77 71.676
R1071 B.n176 B.n76 71.676
R1072 B.n172 B.n75 71.676
R1073 B.n168 B.n74 71.676
R1074 B.n164 B.n73 71.676
R1075 B.n160 B.n72 71.676
R1076 B.n156 B.n71 71.676
R1077 B.n152 B.n70 71.676
R1078 B.n148 B.n69 71.676
R1079 B.n144 B.n68 71.676
R1080 B.n140 B.n67 71.676
R1081 B.n136 B.n66 71.676
R1082 B.n132 B.n65 71.676
R1083 B.n128 B.n64 71.676
R1084 B.n124 B.n63 71.676
R1085 B.n120 B.n62 71.676
R1086 B.n436 B.n435 71.676
R1087 B.n442 B.n441 71.676
R1088 B.n443 B.n432 71.676
R1089 B.n450 B.n449 71.676
R1090 B.n451 B.n430 71.676
R1091 B.n458 B.n457 71.676
R1092 B.n459 B.n428 71.676
R1093 B.n466 B.n465 71.676
R1094 B.n467 B.n426 71.676
R1095 B.n474 B.n473 71.676
R1096 B.n475 B.n424 71.676
R1097 B.n482 B.n481 71.676
R1098 B.n483 B.n422 71.676
R1099 B.n490 B.n489 71.676
R1100 B.n491 B.n420 71.676
R1101 B.n498 B.n497 71.676
R1102 B.n499 B.n418 71.676
R1103 B.n506 B.n505 71.676
R1104 B.n507 B.n416 71.676
R1105 B.n514 B.n513 71.676
R1106 B.n515 B.n414 71.676
R1107 B.n522 B.n521 71.676
R1108 B.n523 B.n410 71.676
R1109 B.n531 B.n530 71.676
R1110 B.n532 B.n408 71.676
R1111 B.n539 B.n538 71.676
R1112 B.n540 B.n406 71.676
R1113 B.n550 B.n549 71.676
R1114 B.n551 B.n404 71.676
R1115 B.n558 B.n557 71.676
R1116 B.n559 B.n402 71.676
R1117 B.n566 B.n565 71.676
R1118 B.n567 B.n400 71.676
R1119 B.n574 B.n573 71.676
R1120 B.n575 B.n398 71.676
R1121 B.n582 B.n581 71.676
R1122 B.n583 B.n396 71.676
R1123 B.n590 B.n589 71.676
R1124 B.n591 B.n394 71.676
R1125 B.n598 B.n597 71.676
R1126 B.n599 B.n392 71.676
R1127 B.n606 B.n605 71.676
R1128 B.n607 B.n390 71.676
R1129 B.n614 B.n613 71.676
R1130 B.n615 B.n388 71.676
R1131 B.n622 B.n621 71.676
R1132 B.n623 B.n386 71.676
R1133 B.n630 B.n629 71.676
R1134 B.n631 B.n384 71.676
R1135 B.n638 B.n637 71.676
R1136 B.n639 B.n382 71.676
R1137 B.n545 B.t20 68.9484
R1138 B.n115 B.t11 68.9484
R1139 B.n412 B.t17 68.9307
R1140 B.n118 B.t14 68.9307
R1141 B.n546 B.n545 59.5399
R1142 B.n527 B.n412 59.5399
R1143 B.n211 B.n118 59.5399
R1144 B.n116 B.n115 59.5399
R1145 B.n645 B.n377 39.4832
R1146 B.n651 B.n377 39.4832
R1147 B.n651 B.n373 39.4832
R1148 B.n658 B.n373 39.4832
R1149 B.n658 B.n657 39.4832
R1150 B.n664 B.n366 39.4832
R1151 B.n670 B.n366 39.4832
R1152 B.n670 B.n362 39.4832
R1153 B.n676 B.n362 39.4832
R1154 B.n676 B.n358 39.4832
R1155 B.n683 B.n358 39.4832
R1156 B.n683 B.n682 39.4832
R1157 B.n689 B.n351 39.4832
R1158 B.n695 B.n351 39.4832
R1159 B.n695 B.n347 39.4832
R1160 B.n701 B.n347 39.4832
R1161 B.n707 B.n343 39.4832
R1162 B.n707 B.n338 39.4832
R1163 B.n713 B.n338 39.4832
R1164 B.n713 B.n339 39.4832
R1165 B.n719 B.n330 39.4832
R1166 B.n725 B.n330 39.4832
R1167 B.n725 B.n331 39.4832
R1168 B.n732 B.n323 39.4832
R1169 B.n738 B.n323 39.4832
R1170 B.n738 B.n4 39.4832
R1171 B.n850 B.n4 39.4832
R1172 B.n850 B.n849 39.4832
R1173 B.n849 B.n848 39.4832
R1174 B.n848 B.n8 39.4832
R1175 B.n842 B.n8 39.4832
R1176 B.n841 B.n840 39.4832
R1177 B.n840 B.n15 39.4832
R1178 B.n834 B.n15 39.4832
R1179 B.n833 B.n832 39.4832
R1180 B.n832 B.n22 39.4832
R1181 B.n826 B.n22 39.4832
R1182 B.n826 B.n825 39.4832
R1183 B.n824 B.n29 39.4832
R1184 B.n818 B.n29 39.4832
R1185 B.n818 B.n817 39.4832
R1186 B.n817 B.n816 39.4832
R1187 B.n810 B.n39 39.4832
R1188 B.n810 B.n809 39.4832
R1189 B.n809 B.n808 39.4832
R1190 B.n808 B.n43 39.4832
R1191 B.n802 B.n43 39.4832
R1192 B.n802 B.n801 39.4832
R1193 B.n801 B.n800 39.4832
R1194 B.n794 B.n53 39.4832
R1195 B.n794 B.n793 39.4832
R1196 B.n793 B.n792 39.4832
R1197 B.n792 B.n57 39.4832
R1198 B.n786 B.n57 39.4832
R1199 B.n331 B.t4 38.9026
R1200 B.t2 B.n841 38.9026
R1201 B.n719 B.t7 33.0963
R1202 B.n834 B.t1 33.0963
R1203 B.n788 B.n59 32.9371
R1204 B.n783 B.n782 32.9371
R1205 B.n643 B.n642 32.9371
R1206 B.n647 B.n379 32.9371
R1207 B.n545 B.n544 31.8066
R1208 B.n412 B.n411 31.8066
R1209 B.n118 B.n117 31.8066
R1210 B.n115 B.n114 31.8066
R1211 B.t3 B.n343 26.1288
R1212 B.n825 B.t6 26.1288
R1213 B.n664 B.t16 20.3225
R1214 B.n682 B.t5 20.3225
R1215 B.n39 B.t0 20.3225
R1216 B.n800 B.t9 20.3225
R1217 B.n657 B.t16 19.1612
R1218 B.n689 B.t5 19.1612
R1219 B.n816 B.t0 19.1612
R1220 B.n53 B.t9 19.1612
R1221 B B.n852 18.0485
R1222 B.n701 B.t3 13.3549
R1223 B.t6 B.n824 13.3549
R1224 B.n119 B.n59 10.6151
R1225 B.n122 B.n119 10.6151
R1226 B.n123 B.n122 10.6151
R1227 B.n126 B.n123 10.6151
R1228 B.n127 B.n126 10.6151
R1229 B.n130 B.n127 10.6151
R1230 B.n131 B.n130 10.6151
R1231 B.n134 B.n131 10.6151
R1232 B.n135 B.n134 10.6151
R1233 B.n138 B.n135 10.6151
R1234 B.n139 B.n138 10.6151
R1235 B.n142 B.n139 10.6151
R1236 B.n143 B.n142 10.6151
R1237 B.n146 B.n143 10.6151
R1238 B.n147 B.n146 10.6151
R1239 B.n150 B.n147 10.6151
R1240 B.n151 B.n150 10.6151
R1241 B.n154 B.n151 10.6151
R1242 B.n155 B.n154 10.6151
R1243 B.n158 B.n155 10.6151
R1244 B.n159 B.n158 10.6151
R1245 B.n162 B.n159 10.6151
R1246 B.n163 B.n162 10.6151
R1247 B.n166 B.n163 10.6151
R1248 B.n167 B.n166 10.6151
R1249 B.n170 B.n167 10.6151
R1250 B.n171 B.n170 10.6151
R1251 B.n174 B.n171 10.6151
R1252 B.n175 B.n174 10.6151
R1253 B.n178 B.n175 10.6151
R1254 B.n179 B.n178 10.6151
R1255 B.n182 B.n179 10.6151
R1256 B.n183 B.n182 10.6151
R1257 B.n186 B.n183 10.6151
R1258 B.n187 B.n186 10.6151
R1259 B.n190 B.n187 10.6151
R1260 B.n191 B.n190 10.6151
R1261 B.n194 B.n191 10.6151
R1262 B.n195 B.n194 10.6151
R1263 B.n198 B.n195 10.6151
R1264 B.n199 B.n198 10.6151
R1265 B.n202 B.n199 10.6151
R1266 B.n203 B.n202 10.6151
R1267 B.n206 B.n203 10.6151
R1268 B.n207 B.n206 10.6151
R1269 B.n210 B.n207 10.6151
R1270 B.n215 B.n212 10.6151
R1271 B.n216 B.n215 10.6151
R1272 B.n219 B.n216 10.6151
R1273 B.n220 B.n219 10.6151
R1274 B.n223 B.n220 10.6151
R1275 B.n224 B.n223 10.6151
R1276 B.n227 B.n224 10.6151
R1277 B.n228 B.n227 10.6151
R1278 B.n232 B.n231 10.6151
R1279 B.n235 B.n232 10.6151
R1280 B.n236 B.n235 10.6151
R1281 B.n239 B.n236 10.6151
R1282 B.n240 B.n239 10.6151
R1283 B.n243 B.n240 10.6151
R1284 B.n244 B.n243 10.6151
R1285 B.n247 B.n244 10.6151
R1286 B.n248 B.n247 10.6151
R1287 B.n251 B.n248 10.6151
R1288 B.n252 B.n251 10.6151
R1289 B.n255 B.n252 10.6151
R1290 B.n256 B.n255 10.6151
R1291 B.n259 B.n256 10.6151
R1292 B.n260 B.n259 10.6151
R1293 B.n263 B.n260 10.6151
R1294 B.n264 B.n263 10.6151
R1295 B.n267 B.n264 10.6151
R1296 B.n268 B.n267 10.6151
R1297 B.n271 B.n268 10.6151
R1298 B.n272 B.n271 10.6151
R1299 B.n275 B.n272 10.6151
R1300 B.n276 B.n275 10.6151
R1301 B.n279 B.n276 10.6151
R1302 B.n280 B.n279 10.6151
R1303 B.n283 B.n280 10.6151
R1304 B.n284 B.n283 10.6151
R1305 B.n287 B.n284 10.6151
R1306 B.n288 B.n287 10.6151
R1307 B.n291 B.n288 10.6151
R1308 B.n292 B.n291 10.6151
R1309 B.n295 B.n292 10.6151
R1310 B.n296 B.n295 10.6151
R1311 B.n299 B.n296 10.6151
R1312 B.n300 B.n299 10.6151
R1313 B.n303 B.n300 10.6151
R1314 B.n304 B.n303 10.6151
R1315 B.n307 B.n304 10.6151
R1316 B.n308 B.n307 10.6151
R1317 B.n311 B.n308 10.6151
R1318 B.n312 B.n311 10.6151
R1319 B.n315 B.n312 10.6151
R1320 B.n316 B.n315 10.6151
R1321 B.n319 B.n316 10.6151
R1322 B.n320 B.n319 10.6151
R1323 B.n783 B.n320 10.6151
R1324 B.n643 B.n375 10.6151
R1325 B.n653 B.n375 10.6151
R1326 B.n654 B.n653 10.6151
R1327 B.n655 B.n654 10.6151
R1328 B.n655 B.n368 10.6151
R1329 B.n666 B.n368 10.6151
R1330 B.n667 B.n666 10.6151
R1331 B.n668 B.n667 10.6151
R1332 B.n668 B.n360 10.6151
R1333 B.n678 B.n360 10.6151
R1334 B.n679 B.n678 10.6151
R1335 B.n680 B.n679 10.6151
R1336 B.n680 B.n353 10.6151
R1337 B.n691 B.n353 10.6151
R1338 B.n692 B.n691 10.6151
R1339 B.n693 B.n692 10.6151
R1340 B.n693 B.n345 10.6151
R1341 B.n703 B.n345 10.6151
R1342 B.n704 B.n703 10.6151
R1343 B.n705 B.n704 10.6151
R1344 B.n705 B.n336 10.6151
R1345 B.n715 B.n336 10.6151
R1346 B.n716 B.n715 10.6151
R1347 B.n717 B.n716 10.6151
R1348 B.n717 B.n328 10.6151
R1349 B.n727 B.n328 10.6151
R1350 B.n728 B.n727 10.6151
R1351 B.n730 B.n728 10.6151
R1352 B.n730 B.n729 10.6151
R1353 B.n729 B.n321 10.6151
R1354 B.n741 B.n321 10.6151
R1355 B.n742 B.n741 10.6151
R1356 B.n743 B.n742 10.6151
R1357 B.n744 B.n743 10.6151
R1358 B.n746 B.n744 10.6151
R1359 B.n747 B.n746 10.6151
R1360 B.n748 B.n747 10.6151
R1361 B.n749 B.n748 10.6151
R1362 B.n751 B.n749 10.6151
R1363 B.n752 B.n751 10.6151
R1364 B.n753 B.n752 10.6151
R1365 B.n754 B.n753 10.6151
R1366 B.n756 B.n754 10.6151
R1367 B.n757 B.n756 10.6151
R1368 B.n758 B.n757 10.6151
R1369 B.n759 B.n758 10.6151
R1370 B.n761 B.n759 10.6151
R1371 B.n762 B.n761 10.6151
R1372 B.n763 B.n762 10.6151
R1373 B.n764 B.n763 10.6151
R1374 B.n766 B.n764 10.6151
R1375 B.n767 B.n766 10.6151
R1376 B.n768 B.n767 10.6151
R1377 B.n769 B.n768 10.6151
R1378 B.n771 B.n769 10.6151
R1379 B.n772 B.n771 10.6151
R1380 B.n773 B.n772 10.6151
R1381 B.n774 B.n773 10.6151
R1382 B.n776 B.n774 10.6151
R1383 B.n777 B.n776 10.6151
R1384 B.n778 B.n777 10.6151
R1385 B.n779 B.n778 10.6151
R1386 B.n781 B.n779 10.6151
R1387 B.n782 B.n781 10.6151
R1388 B.n437 B.n379 10.6151
R1389 B.n438 B.n437 10.6151
R1390 B.n439 B.n438 10.6151
R1391 B.n439 B.n433 10.6151
R1392 B.n445 B.n433 10.6151
R1393 B.n446 B.n445 10.6151
R1394 B.n447 B.n446 10.6151
R1395 B.n447 B.n431 10.6151
R1396 B.n453 B.n431 10.6151
R1397 B.n454 B.n453 10.6151
R1398 B.n455 B.n454 10.6151
R1399 B.n455 B.n429 10.6151
R1400 B.n461 B.n429 10.6151
R1401 B.n462 B.n461 10.6151
R1402 B.n463 B.n462 10.6151
R1403 B.n463 B.n427 10.6151
R1404 B.n469 B.n427 10.6151
R1405 B.n470 B.n469 10.6151
R1406 B.n471 B.n470 10.6151
R1407 B.n471 B.n425 10.6151
R1408 B.n477 B.n425 10.6151
R1409 B.n478 B.n477 10.6151
R1410 B.n479 B.n478 10.6151
R1411 B.n479 B.n423 10.6151
R1412 B.n485 B.n423 10.6151
R1413 B.n486 B.n485 10.6151
R1414 B.n487 B.n486 10.6151
R1415 B.n487 B.n421 10.6151
R1416 B.n493 B.n421 10.6151
R1417 B.n494 B.n493 10.6151
R1418 B.n495 B.n494 10.6151
R1419 B.n495 B.n419 10.6151
R1420 B.n501 B.n419 10.6151
R1421 B.n502 B.n501 10.6151
R1422 B.n503 B.n502 10.6151
R1423 B.n503 B.n417 10.6151
R1424 B.n509 B.n417 10.6151
R1425 B.n510 B.n509 10.6151
R1426 B.n511 B.n510 10.6151
R1427 B.n511 B.n415 10.6151
R1428 B.n517 B.n415 10.6151
R1429 B.n518 B.n517 10.6151
R1430 B.n519 B.n518 10.6151
R1431 B.n519 B.n413 10.6151
R1432 B.n525 B.n413 10.6151
R1433 B.n526 B.n525 10.6151
R1434 B.n528 B.n409 10.6151
R1435 B.n534 B.n409 10.6151
R1436 B.n535 B.n534 10.6151
R1437 B.n536 B.n535 10.6151
R1438 B.n536 B.n407 10.6151
R1439 B.n542 B.n407 10.6151
R1440 B.n543 B.n542 10.6151
R1441 B.n547 B.n543 10.6151
R1442 B.n553 B.n405 10.6151
R1443 B.n554 B.n553 10.6151
R1444 B.n555 B.n554 10.6151
R1445 B.n555 B.n403 10.6151
R1446 B.n561 B.n403 10.6151
R1447 B.n562 B.n561 10.6151
R1448 B.n563 B.n562 10.6151
R1449 B.n563 B.n401 10.6151
R1450 B.n569 B.n401 10.6151
R1451 B.n570 B.n569 10.6151
R1452 B.n571 B.n570 10.6151
R1453 B.n571 B.n399 10.6151
R1454 B.n577 B.n399 10.6151
R1455 B.n578 B.n577 10.6151
R1456 B.n579 B.n578 10.6151
R1457 B.n579 B.n397 10.6151
R1458 B.n585 B.n397 10.6151
R1459 B.n586 B.n585 10.6151
R1460 B.n587 B.n586 10.6151
R1461 B.n587 B.n395 10.6151
R1462 B.n593 B.n395 10.6151
R1463 B.n594 B.n593 10.6151
R1464 B.n595 B.n594 10.6151
R1465 B.n595 B.n393 10.6151
R1466 B.n601 B.n393 10.6151
R1467 B.n602 B.n601 10.6151
R1468 B.n603 B.n602 10.6151
R1469 B.n603 B.n391 10.6151
R1470 B.n609 B.n391 10.6151
R1471 B.n610 B.n609 10.6151
R1472 B.n611 B.n610 10.6151
R1473 B.n611 B.n389 10.6151
R1474 B.n617 B.n389 10.6151
R1475 B.n618 B.n617 10.6151
R1476 B.n619 B.n618 10.6151
R1477 B.n619 B.n387 10.6151
R1478 B.n625 B.n387 10.6151
R1479 B.n626 B.n625 10.6151
R1480 B.n627 B.n626 10.6151
R1481 B.n627 B.n385 10.6151
R1482 B.n633 B.n385 10.6151
R1483 B.n634 B.n633 10.6151
R1484 B.n635 B.n634 10.6151
R1485 B.n635 B.n383 10.6151
R1486 B.n641 B.n383 10.6151
R1487 B.n642 B.n641 10.6151
R1488 B.n648 B.n647 10.6151
R1489 B.n649 B.n648 10.6151
R1490 B.n649 B.n371 10.6151
R1491 B.n660 B.n371 10.6151
R1492 B.n661 B.n660 10.6151
R1493 B.n662 B.n661 10.6151
R1494 B.n662 B.n364 10.6151
R1495 B.n672 B.n364 10.6151
R1496 B.n673 B.n672 10.6151
R1497 B.n674 B.n673 10.6151
R1498 B.n674 B.n356 10.6151
R1499 B.n685 B.n356 10.6151
R1500 B.n686 B.n685 10.6151
R1501 B.n687 B.n686 10.6151
R1502 B.n687 B.n349 10.6151
R1503 B.n697 B.n349 10.6151
R1504 B.n698 B.n697 10.6151
R1505 B.n699 B.n698 10.6151
R1506 B.n699 B.n341 10.6151
R1507 B.n709 B.n341 10.6151
R1508 B.n710 B.n709 10.6151
R1509 B.n711 B.n710 10.6151
R1510 B.n711 B.n333 10.6151
R1511 B.n721 B.n333 10.6151
R1512 B.n722 B.n721 10.6151
R1513 B.n723 B.n722 10.6151
R1514 B.n723 B.n325 10.6151
R1515 B.n734 B.n325 10.6151
R1516 B.n735 B.n734 10.6151
R1517 B.n736 B.n735 10.6151
R1518 B.n736 B.n0 10.6151
R1519 B.n846 B.n1 10.6151
R1520 B.n846 B.n845 10.6151
R1521 B.n845 B.n844 10.6151
R1522 B.n844 B.n10 10.6151
R1523 B.n838 B.n10 10.6151
R1524 B.n838 B.n837 10.6151
R1525 B.n837 B.n836 10.6151
R1526 B.n836 B.n17 10.6151
R1527 B.n830 B.n17 10.6151
R1528 B.n830 B.n829 10.6151
R1529 B.n829 B.n828 10.6151
R1530 B.n828 B.n24 10.6151
R1531 B.n822 B.n24 10.6151
R1532 B.n822 B.n821 10.6151
R1533 B.n821 B.n820 10.6151
R1534 B.n820 B.n31 10.6151
R1535 B.n814 B.n31 10.6151
R1536 B.n814 B.n813 10.6151
R1537 B.n813 B.n812 10.6151
R1538 B.n812 B.n37 10.6151
R1539 B.n806 B.n37 10.6151
R1540 B.n806 B.n805 10.6151
R1541 B.n805 B.n804 10.6151
R1542 B.n804 B.n45 10.6151
R1543 B.n798 B.n45 10.6151
R1544 B.n798 B.n797 10.6151
R1545 B.n797 B.n796 10.6151
R1546 B.n796 B.n51 10.6151
R1547 B.n790 B.n51 10.6151
R1548 B.n790 B.n789 10.6151
R1549 B.n789 B.n788 10.6151
R1550 B.n212 B.n211 6.5566
R1551 B.n228 B.n116 6.5566
R1552 B.n528 B.n527 6.5566
R1553 B.n547 B.n546 6.5566
R1554 B.n339 B.t7 6.38741
R1555 B.t1 B.n833 6.38741
R1556 B.n211 B.n210 4.05904
R1557 B.n231 B.n116 4.05904
R1558 B.n527 B.n526 4.05904
R1559 B.n546 B.n405 4.05904
R1560 B.n852 B.n0 2.81026
R1561 B.n852 B.n1 2.81026
R1562 B.n732 B.t4 0.581128
R1563 B.n842 B.t2 0.581128
R1564 VN.n5 VN.t6 279.003
R1565 VN.n25 VN.t3 279.003
R1566 VN.n4 VN.t1 251.487
R1567 VN.n10 VN.t0 251.487
R1568 VN.n17 VN.t5 251.487
R1569 VN.n24 VN.t2 251.487
R1570 VN.n22 VN.t4 251.487
R1571 VN.n36 VN.t7 251.487
R1572 VN.n18 VN.n17 175.492
R1573 VN.n37 VN.n36 175.492
R1574 VN.n35 VN.n19 161.3
R1575 VN.n34 VN.n33 161.3
R1576 VN.n32 VN.n20 161.3
R1577 VN.n31 VN.n30 161.3
R1578 VN.n29 VN.n21 161.3
R1579 VN.n28 VN.n27 161.3
R1580 VN.n26 VN.n23 161.3
R1581 VN.n16 VN.n0 161.3
R1582 VN.n15 VN.n14 161.3
R1583 VN.n13 VN.n1 161.3
R1584 VN.n12 VN.n11 161.3
R1585 VN.n9 VN.n2 161.3
R1586 VN.n8 VN.n7 161.3
R1587 VN.n6 VN.n3 161.3
R1588 VN.n5 VN.n4 62.0576
R1589 VN.n25 VN.n24 62.0576
R1590 VN.n9 VN.n8 56.5193
R1591 VN.n29 VN.n28 56.5193
R1592 VN.n15 VN.n1 51.1773
R1593 VN.n34 VN.n20 51.1773
R1594 VN VN.n37 46.3888
R1595 VN.n16 VN.n15 29.8095
R1596 VN.n35 VN.n34 29.8095
R1597 VN.n26 VN.n25 27.6443
R1598 VN.n6 VN.n5 27.6443
R1599 VN.n8 VN.n3 24.4675
R1600 VN.n11 VN.n9 24.4675
R1601 VN.n28 VN.n23 24.4675
R1602 VN.n30 VN.n29 24.4675
R1603 VN.n10 VN.n1 21.0421
R1604 VN.n22 VN.n20 21.0421
R1605 VN.n17 VN.n16 10.2766
R1606 VN.n36 VN.n35 10.2766
R1607 VN.n4 VN.n3 3.42588
R1608 VN.n11 VN.n10 3.42588
R1609 VN.n24 VN.n23 3.42588
R1610 VN.n30 VN.n22 3.42588
R1611 VN.n37 VN.n19 0.189894
R1612 VN.n33 VN.n19 0.189894
R1613 VN.n33 VN.n32 0.189894
R1614 VN.n32 VN.n31 0.189894
R1615 VN.n31 VN.n21 0.189894
R1616 VN.n27 VN.n21 0.189894
R1617 VN.n27 VN.n26 0.189894
R1618 VN.n7 VN.n6 0.189894
R1619 VN.n7 VN.n2 0.189894
R1620 VN.n12 VN.n2 0.189894
R1621 VN.n13 VN.n12 0.189894
R1622 VN.n14 VN.n13 0.189894
R1623 VN.n14 VN.n0 0.189894
R1624 VN.n18 VN.n0 0.189894
R1625 VN VN.n18 0.0516364
R1626 VDD2.n2 VDD2.n1 63.8518
R1627 VDD2.n2 VDD2.n0 63.8518
R1628 VDD2 VDD2.n5 63.849
R1629 VDD2.n4 VDD2.n3 63.2005
R1630 VDD2.n4 VDD2.n2 41.8618
R1631 VDD2.n5 VDD2.t5 1.44893
R1632 VDD2.n5 VDD2.t4 1.44893
R1633 VDD2.n3 VDD2.t0 1.44893
R1634 VDD2.n3 VDD2.t3 1.44893
R1635 VDD2.n1 VDD2.t7 1.44893
R1636 VDD2.n1 VDD2.t2 1.44893
R1637 VDD2.n0 VDD2.t1 1.44893
R1638 VDD2.n0 VDD2.t6 1.44893
R1639 VDD2 VDD2.n4 0.765586
C0 VDD1 VP 8.4123f
C1 VDD1 VN 0.149246f
C2 VP VN 6.39672f
C3 VDD2 VDD1 1.13131f
C4 VDD2 VP 0.382251f
C5 VDD2 VN 8.18004f
C6 VDD1 VTAIL 9.60307f
C7 VP VTAIL 8.1076f
C8 VN VTAIL 8.093491f
C9 VDD2 VTAIL 9.648839f
C10 VDD2 B 4.201219f
C11 VDD1 B 4.500046f
C12 VTAIL B 10.462293f
C13 VN B 10.865089f
C14 VP B 9.136149f
C15 VDD2.t1 B 0.272565f
C16 VDD2.t6 B 0.272565f
C17 VDD2.n0 B 2.45889f
C18 VDD2.t7 B 0.272565f
C19 VDD2.t2 B 0.272565f
C20 VDD2.n1 B 2.45889f
C21 VDD2.n2 B 2.64617f
C22 VDD2.t0 B 0.272565f
C23 VDD2.t3 B 0.272565f
C24 VDD2.n3 B 2.455f
C25 VDD2.n4 B 2.65003f
C26 VDD2.t5 B 0.272565f
C27 VDD2.t4 B 0.272565f
C28 VDD2.n5 B 2.45886f
C29 VN.n0 B 0.03303f
C30 VN.t5 B 1.61723f
C31 VN.n1 B 0.055716f
C32 VN.n2 B 0.03303f
C33 VN.n3 B 0.035423f
C34 VN.t6 B 1.68499f
C35 VN.t1 B 1.61723f
C36 VN.n4 B 0.62701f
C37 VN.n5 B 0.666554f
C38 VN.n6 B 0.173291f
C39 VN.n7 B 0.03303f
C40 VN.n8 B 0.048218f
C41 VN.n9 B 0.048218f
C42 VN.t0 B 1.61723f
C43 VN.n10 B 0.582943f
C44 VN.n11 B 0.035423f
C45 VN.n12 B 0.03303f
C46 VN.n13 B 0.03303f
C47 VN.n14 B 0.03303f
C48 VN.n15 B 0.032219f
C49 VN.n16 B 0.048179f
C50 VN.n17 B 0.640643f
C51 VN.n18 B 0.030674f
C52 VN.n19 B 0.03303f
C53 VN.t7 B 1.61723f
C54 VN.n20 B 0.055716f
C55 VN.n21 B 0.03303f
C56 VN.t4 B 1.61723f
C57 VN.n22 B 0.582943f
C58 VN.n23 B 0.035423f
C59 VN.t3 B 1.68499f
C60 VN.t2 B 1.61723f
C61 VN.n24 B 0.62701f
C62 VN.n25 B 0.666554f
C63 VN.n26 B 0.173291f
C64 VN.n27 B 0.03303f
C65 VN.n28 B 0.048218f
C66 VN.n29 B 0.048218f
C67 VN.n30 B 0.035423f
C68 VN.n31 B 0.03303f
C69 VN.n32 B 0.03303f
C70 VN.n33 B 0.03303f
C71 VN.n34 B 0.032219f
C72 VN.n35 B 0.048179f
C73 VN.n36 B 0.640643f
C74 VN.n37 B 1.60675f
C75 VTAIL.t1 B 0.20415f
C76 VTAIL.t6 B 0.20415f
C77 VTAIL.n0 B 1.78563f
C78 VTAIL.n1 B 0.268922f
C79 VTAIL.t2 B 2.27784f
C80 VTAIL.n2 B 0.358553f
C81 VTAIL.t13 B 2.27784f
C82 VTAIL.n3 B 0.358553f
C83 VTAIL.t9 B 0.20415f
C84 VTAIL.t14 B 0.20415f
C85 VTAIL.n4 B 1.78563f
C86 VTAIL.n5 B 0.351471f
C87 VTAIL.t12 B 2.27784f
C88 VTAIL.n6 B 1.39037f
C89 VTAIL.t5 B 2.27784f
C90 VTAIL.n7 B 1.39036f
C91 VTAIL.t3 B 0.20415f
C92 VTAIL.t15 B 0.20415f
C93 VTAIL.n8 B 1.78563f
C94 VTAIL.n9 B 0.351469f
C95 VTAIL.t4 B 2.27784f
C96 VTAIL.n10 B 0.35855f
C97 VTAIL.t7 B 2.27784f
C98 VTAIL.n11 B 0.35855f
C99 VTAIL.t8 B 0.20415f
C100 VTAIL.t10 B 0.20415f
C101 VTAIL.n12 B 1.78563f
C102 VTAIL.n13 B 0.351469f
C103 VTAIL.t11 B 2.27784f
C104 VTAIL.n14 B 1.39037f
C105 VTAIL.t0 B 2.27784f
C106 VTAIL.n15 B 1.38682f
C107 VDD1.t3 B 0.274192f
C108 VDD1.t4 B 0.274192f
C109 VDD1.n0 B 2.47434f
C110 VDD1.t6 B 0.274192f
C111 VDD1.t5 B 0.274192f
C112 VDD1.n1 B 2.47357f
C113 VDD1.t0 B 0.274192f
C114 VDD1.t7 B 0.274192f
C115 VDD1.n2 B 2.47357f
C116 VDD1.n3 B 2.71558f
C117 VDD1.t1 B 0.274192f
C118 VDD1.t2 B 0.274192f
C119 VDD1.n4 B 2.46965f
C120 VDD1.n5 B 2.69647f
C121 VP.n0 B 0.03339f
C122 VP.t1 B 1.63482f
C123 VP.n1 B 0.056322f
C124 VP.n2 B 0.03339f
C125 VP.n3 B 0.035808f
C126 VP.n4 B 0.03339f
C127 VP.t2 B 1.63482f
C128 VP.n5 B 0.647612f
C129 VP.n6 B 0.03339f
C130 VP.t3 B 1.63482f
C131 VP.n7 B 0.056322f
C132 VP.n8 B 0.03339f
C133 VP.n9 B 0.035808f
C134 VP.t7 B 1.70332f
C135 VP.t6 B 1.63482f
C136 VP.n10 B 0.63383f
C137 VP.n11 B 0.673805f
C138 VP.n12 B 0.175176f
C139 VP.n13 B 0.03339f
C140 VP.n14 B 0.048743f
C141 VP.n15 B 0.048743f
C142 VP.t4 B 1.63482f
C143 VP.n16 B 0.589284f
C144 VP.n17 B 0.035808f
C145 VP.n18 B 0.03339f
C146 VP.n19 B 0.03339f
C147 VP.n20 B 0.03339f
C148 VP.n21 B 0.032569f
C149 VP.n22 B 0.048703f
C150 VP.n23 B 0.647612f
C151 VP.n24 B 1.60243f
C152 VP.n25 B 1.62851f
C153 VP.n26 B 0.03339f
C154 VP.n27 B 0.048703f
C155 VP.n28 B 0.032569f
C156 VP.t5 B 1.63482f
C157 VP.n29 B 0.589284f
C158 VP.n30 B 0.056322f
C159 VP.n31 B 0.03339f
C160 VP.n32 B 0.03339f
C161 VP.n33 B 0.03339f
C162 VP.n34 B 0.048743f
C163 VP.n35 B 0.048743f
C164 VP.t0 B 1.63482f
C165 VP.n36 B 0.589284f
C166 VP.n37 B 0.035808f
C167 VP.n38 B 0.03339f
C168 VP.n39 B 0.03339f
C169 VP.n40 B 0.03339f
C170 VP.n41 B 0.032569f
C171 VP.n42 B 0.048703f
C172 VP.n43 B 0.647612f
C173 VP.n44 B 0.031007f
.ends

