* NGSPICE file created from diff_pair_sample_0781.ext - technology: sky130A

.subckt diff_pair_sample_0781 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t17 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=1.0803 pd=6.32 as=0.45705 ps=3.1 w=2.77 l=0.67
X1 B.t11 B.t9 B.t10 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=1.0803 pd=6.32 as=0 ps=0 w=2.77 l=0.67
X2 VTAIL.t5 VP.t0 VDD1.t9 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=0.45705 pd=3.1 as=0.45705 ps=3.1 w=2.77 l=0.67
X3 VDD2.t8 VN.t1 VTAIL.t13 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=0.45705 pd=3.1 as=0.45705 ps=3.1 w=2.77 l=0.67
X4 B.t8 B.t6 B.t7 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=1.0803 pd=6.32 as=0 ps=0 w=2.77 l=0.67
X5 VDD2.t7 VN.t2 VTAIL.t10 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=1.0803 pd=6.32 as=0.45705 ps=3.1 w=2.77 l=0.67
X6 VDD1.t8 VP.t1 VTAIL.t0 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=0.45705 pd=3.1 as=1.0803 ps=6.32 w=2.77 l=0.67
X7 VDD2.t6 VN.t3 VTAIL.t12 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=0.45705 pd=3.1 as=0.45705 ps=3.1 w=2.77 l=0.67
X8 VDD1.t7 VP.t2 VTAIL.t19 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=0.45705 pd=3.1 as=0.45705 ps=3.1 w=2.77 l=0.67
X9 VTAIL.t2 VP.t3 VDD1.t6 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=0.45705 pd=3.1 as=0.45705 ps=3.1 w=2.77 l=0.67
X10 B.t5 B.t3 B.t4 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=1.0803 pd=6.32 as=0 ps=0 w=2.77 l=0.67
X11 VDD1.t5 VP.t4 VTAIL.t1 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=1.0803 pd=6.32 as=0.45705 ps=3.1 w=2.77 l=0.67
X12 VDD2.t5 VN.t4 VTAIL.t15 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=0.45705 pd=3.1 as=1.0803 ps=6.32 w=2.77 l=0.67
X13 VDD2.t4 VN.t5 VTAIL.t16 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=0.45705 pd=3.1 as=1.0803 ps=6.32 w=2.77 l=0.67
X14 B.t2 B.t0 B.t1 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=1.0803 pd=6.32 as=0 ps=0 w=2.77 l=0.67
X15 VDD1.t4 VP.t5 VTAIL.t18 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=0.45705 pd=3.1 as=1.0803 ps=6.32 w=2.77 l=0.67
X16 VTAIL.t14 VN.t6 VDD2.t3 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=0.45705 pd=3.1 as=0.45705 ps=3.1 w=2.77 l=0.67
X17 VDD1.t3 VP.t6 VTAIL.t3 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=0.45705 pd=3.1 as=0.45705 ps=3.1 w=2.77 l=0.67
X18 VTAIL.t8 VN.t7 VDD2.t2 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=0.45705 pd=3.1 as=0.45705 ps=3.1 w=2.77 l=0.67
X19 VTAIL.t9 VN.t8 VDD2.t1 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=0.45705 pd=3.1 as=0.45705 ps=3.1 w=2.77 l=0.67
X20 VTAIL.t11 VN.t9 VDD2.t0 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=0.45705 pd=3.1 as=0.45705 ps=3.1 w=2.77 l=0.67
X21 VTAIL.t7 VP.t7 VDD1.t2 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=0.45705 pd=3.1 as=0.45705 ps=3.1 w=2.77 l=0.67
X22 VTAIL.t6 VP.t8 VDD1.t1 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=0.45705 pd=3.1 as=0.45705 ps=3.1 w=2.77 l=0.67
X23 VDD1.t0 VP.t9 VTAIL.t4 w_n2170_n1522# sky130_fd_pr__pfet_01v8 ad=1.0803 pd=6.32 as=0.45705 ps=3.1 w=2.77 l=0.67
R0 VN.n3 VN.t2 179.625
R1 VN.n17 VN.t4 179.625
R2 VN.n13 VN.n12 161.3
R3 VN.n27 VN.n26 161.3
R4 VN.n25 VN.n14 161.3
R5 VN.n24 VN.n23 161.3
R6 VN.n22 VN.n15 161.3
R7 VN.n21 VN.n20 161.3
R8 VN.n19 VN.n16 161.3
R9 VN.n11 VN.n0 161.3
R10 VN.n10 VN.n9 161.3
R11 VN.n8 VN.n1 161.3
R12 VN.n7 VN.n6 161.3
R13 VN.n5 VN.n2 161.3
R14 VN.n4 VN.t7 158.629
R15 VN.n6 VN.t3 158.629
R16 VN.n10 VN.t9 158.629
R17 VN.n12 VN.t5 158.629
R18 VN.n18 VN.t8 158.629
R19 VN.n20 VN.t1 158.629
R20 VN.n24 VN.t6 158.629
R21 VN.n26 VN.t0 158.629
R22 VN.n17 VN.n16 44.8515
R23 VN.n3 VN.n2 44.8515
R24 VN VN.n27 35.9569
R25 VN.n5 VN.n4 24.1005
R26 VN.n6 VN.n5 24.1005
R27 VN.n6 VN.n1 24.1005
R28 VN.n10 VN.n1 24.1005
R29 VN.n11 VN.n10 24.1005
R30 VN.n12 VN.n11 24.1005
R31 VN.n20 VN.n19 24.1005
R32 VN.n19 VN.n18 24.1005
R33 VN.n24 VN.n15 24.1005
R34 VN.n20 VN.n15 24.1005
R35 VN.n26 VN.n25 24.1005
R36 VN.n25 VN.n24 24.1005
R37 VN.n4 VN.n3 20.9471
R38 VN.n18 VN.n17 20.9471
R39 VN.n27 VN.n14 0.189894
R40 VN.n23 VN.n14 0.189894
R41 VN.n23 VN.n22 0.189894
R42 VN.n22 VN.n21 0.189894
R43 VN.n21 VN.n16 0.189894
R44 VN.n7 VN.n2 0.189894
R45 VN.n8 VN.n7 0.189894
R46 VN.n9 VN.n8 0.189894
R47 VN.n9 VN.n0 0.189894
R48 VN.n13 VN.n0 0.189894
R49 VN VN.n13 0.0516364
R50 VTAIL.n11 VTAIL.t15 133.321
R51 VTAIL.n17 VTAIL.t16 133.32
R52 VTAIL.n2 VTAIL.t0 133.32
R53 VTAIL.n16 VTAIL.t18 133.32
R54 VTAIL.n15 VTAIL.n14 121.585
R55 VTAIL.n13 VTAIL.n12 121.585
R56 VTAIL.n10 VTAIL.n9 121.585
R57 VTAIL.n8 VTAIL.n7 121.585
R58 VTAIL.n19 VTAIL.n18 121.585
R59 VTAIL.n1 VTAIL.n0 121.585
R60 VTAIL.n4 VTAIL.n3 121.585
R61 VTAIL.n6 VTAIL.n5 121.585
R62 VTAIL.n8 VTAIL.n6 16.4789
R63 VTAIL.n17 VTAIL.n16 15.6169
R64 VTAIL.n18 VTAIL.t12 11.7352
R65 VTAIL.n18 VTAIL.t11 11.7352
R66 VTAIL.n0 VTAIL.t10 11.7352
R67 VTAIL.n0 VTAIL.t8 11.7352
R68 VTAIL.n3 VTAIL.t19 11.7352
R69 VTAIL.n3 VTAIL.t7 11.7352
R70 VTAIL.n5 VTAIL.t1 11.7352
R71 VTAIL.n5 VTAIL.t6 11.7352
R72 VTAIL.n14 VTAIL.t3 11.7352
R73 VTAIL.n14 VTAIL.t5 11.7352
R74 VTAIL.n12 VTAIL.t4 11.7352
R75 VTAIL.n12 VTAIL.t2 11.7352
R76 VTAIL.n9 VTAIL.t13 11.7352
R77 VTAIL.n9 VTAIL.t9 11.7352
R78 VTAIL.n7 VTAIL.t17 11.7352
R79 VTAIL.n7 VTAIL.t14 11.7352
R80 VTAIL.n13 VTAIL.n11 0.901362
R81 VTAIL.n2 VTAIL.n1 0.901362
R82 VTAIL.n10 VTAIL.n8 0.862569
R83 VTAIL.n11 VTAIL.n10 0.862569
R84 VTAIL.n15 VTAIL.n13 0.862569
R85 VTAIL.n16 VTAIL.n15 0.862569
R86 VTAIL.n6 VTAIL.n4 0.862569
R87 VTAIL.n4 VTAIL.n2 0.862569
R88 VTAIL.n19 VTAIL.n17 0.862569
R89 VTAIL VTAIL.n1 0.705241
R90 VTAIL VTAIL.n19 0.157828
R91 VDD2.n1 VDD2.t7 150.861
R92 VDD2.n4 VDD2.t9 149.999
R93 VDD2.n3 VDD2.n2 138.856
R94 VDD2 VDD2.n7 138.852
R95 VDD2.n6 VDD2.n5 138.264
R96 VDD2.n1 VDD2.n0 138.263
R97 VDD2.n4 VDD2.n3 30.1981
R98 VDD2.n7 VDD2.t1 11.7352
R99 VDD2.n7 VDD2.t5 11.7352
R100 VDD2.n5 VDD2.t3 11.7352
R101 VDD2.n5 VDD2.t8 11.7352
R102 VDD2.n2 VDD2.t0 11.7352
R103 VDD2.n2 VDD2.t4 11.7352
R104 VDD2.n0 VDD2.t2 11.7352
R105 VDD2.n0 VDD2.t6 11.7352
R106 VDD2.n6 VDD2.n4 0.862569
R107 VDD2 VDD2.n6 0.274207
R108 VDD2.n3 VDD2.n1 0.160671
R109 B.n194 B.n193 585
R110 B.n192 B.n65 585
R111 B.n191 B.n190 585
R112 B.n189 B.n66 585
R113 B.n188 B.n187 585
R114 B.n186 B.n67 585
R115 B.n185 B.n184 585
R116 B.n183 B.n68 585
R117 B.n182 B.n181 585
R118 B.n180 B.n69 585
R119 B.n179 B.n178 585
R120 B.n177 B.n70 585
R121 B.n176 B.n175 585
R122 B.n174 B.n71 585
R123 B.n173 B.n172 585
R124 B.n168 B.n72 585
R125 B.n167 B.n166 585
R126 B.n165 B.n73 585
R127 B.n164 B.n163 585
R128 B.n162 B.n74 585
R129 B.n161 B.n160 585
R130 B.n159 B.n75 585
R131 B.n158 B.n157 585
R132 B.n156 B.n76 585
R133 B.n154 B.n153 585
R134 B.n152 B.n79 585
R135 B.n151 B.n150 585
R136 B.n149 B.n80 585
R137 B.n148 B.n147 585
R138 B.n146 B.n81 585
R139 B.n145 B.n144 585
R140 B.n143 B.n82 585
R141 B.n142 B.n141 585
R142 B.n140 B.n83 585
R143 B.n139 B.n138 585
R144 B.n137 B.n84 585
R145 B.n136 B.n135 585
R146 B.n134 B.n85 585
R147 B.n195 B.n64 585
R148 B.n197 B.n196 585
R149 B.n198 B.n63 585
R150 B.n200 B.n199 585
R151 B.n201 B.n62 585
R152 B.n203 B.n202 585
R153 B.n204 B.n61 585
R154 B.n206 B.n205 585
R155 B.n207 B.n60 585
R156 B.n209 B.n208 585
R157 B.n210 B.n59 585
R158 B.n212 B.n211 585
R159 B.n213 B.n58 585
R160 B.n215 B.n214 585
R161 B.n216 B.n57 585
R162 B.n218 B.n217 585
R163 B.n219 B.n56 585
R164 B.n221 B.n220 585
R165 B.n222 B.n55 585
R166 B.n224 B.n223 585
R167 B.n225 B.n54 585
R168 B.n227 B.n226 585
R169 B.n228 B.n53 585
R170 B.n230 B.n229 585
R171 B.n231 B.n52 585
R172 B.n233 B.n232 585
R173 B.n234 B.n51 585
R174 B.n236 B.n235 585
R175 B.n237 B.n50 585
R176 B.n239 B.n238 585
R177 B.n240 B.n49 585
R178 B.n242 B.n241 585
R179 B.n243 B.n48 585
R180 B.n245 B.n244 585
R181 B.n246 B.n47 585
R182 B.n248 B.n247 585
R183 B.n249 B.n46 585
R184 B.n251 B.n250 585
R185 B.n252 B.n45 585
R186 B.n254 B.n253 585
R187 B.n255 B.n44 585
R188 B.n257 B.n256 585
R189 B.n258 B.n43 585
R190 B.n260 B.n259 585
R191 B.n261 B.n42 585
R192 B.n263 B.n262 585
R193 B.n264 B.n41 585
R194 B.n266 B.n265 585
R195 B.n267 B.n40 585
R196 B.n269 B.n268 585
R197 B.n270 B.n39 585
R198 B.n272 B.n271 585
R199 B.n330 B.n329 585
R200 B.n328 B.n15 585
R201 B.n327 B.n326 585
R202 B.n325 B.n16 585
R203 B.n324 B.n323 585
R204 B.n322 B.n17 585
R205 B.n321 B.n320 585
R206 B.n319 B.n18 585
R207 B.n318 B.n317 585
R208 B.n316 B.n19 585
R209 B.n315 B.n314 585
R210 B.n313 B.n20 585
R211 B.n312 B.n311 585
R212 B.n310 B.n21 585
R213 B.n308 B.n307 585
R214 B.n306 B.n24 585
R215 B.n305 B.n304 585
R216 B.n303 B.n25 585
R217 B.n302 B.n301 585
R218 B.n300 B.n26 585
R219 B.n299 B.n298 585
R220 B.n297 B.n27 585
R221 B.n296 B.n295 585
R222 B.n294 B.n28 585
R223 B.n293 B.n292 585
R224 B.n291 B.n29 585
R225 B.n290 B.n289 585
R226 B.n288 B.n33 585
R227 B.n287 B.n286 585
R228 B.n285 B.n34 585
R229 B.n284 B.n283 585
R230 B.n282 B.n35 585
R231 B.n281 B.n280 585
R232 B.n279 B.n36 585
R233 B.n278 B.n277 585
R234 B.n276 B.n37 585
R235 B.n275 B.n274 585
R236 B.n273 B.n38 585
R237 B.n331 B.n14 585
R238 B.n333 B.n332 585
R239 B.n334 B.n13 585
R240 B.n336 B.n335 585
R241 B.n337 B.n12 585
R242 B.n339 B.n338 585
R243 B.n340 B.n11 585
R244 B.n342 B.n341 585
R245 B.n343 B.n10 585
R246 B.n345 B.n344 585
R247 B.n346 B.n9 585
R248 B.n348 B.n347 585
R249 B.n349 B.n8 585
R250 B.n351 B.n350 585
R251 B.n352 B.n7 585
R252 B.n354 B.n353 585
R253 B.n355 B.n6 585
R254 B.n357 B.n356 585
R255 B.n358 B.n5 585
R256 B.n360 B.n359 585
R257 B.n361 B.n4 585
R258 B.n363 B.n362 585
R259 B.n364 B.n3 585
R260 B.n366 B.n365 585
R261 B.n367 B.n0 585
R262 B.n2 B.n1 585
R263 B.n98 B.n97 585
R264 B.n100 B.n99 585
R265 B.n101 B.n96 585
R266 B.n103 B.n102 585
R267 B.n104 B.n95 585
R268 B.n106 B.n105 585
R269 B.n107 B.n94 585
R270 B.n109 B.n108 585
R271 B.n110 B.n93 585
R272 B.n112 B.n111 585
R273 B.n113 B.n92 585
R274 B.n115 B.n114 585
R275 B.n116 B.n91 585
R276 B.n118 B.n117 585
R277 B.n119 B.n90 585
R278 B.n121 B.n120 585
R279 B.n122 B.n89 585
R280 B.n124 B.n123 585
R281 B.n125 B.n88 585
R282 B.n127 B.n126 585
R283 B.n128 B.n87 585
R284 B.n130 B.n129 585
R285 B.n131 B.n86 585
R286 B.n133 B.n132 585
R287 B.n134 B.n133 583.793
R288 B.n193 B.n64 583.793
R289 B.n271 B.n38 583.793
R290 B.n331 B.n330 583.793
R291 B.n77 B.t0 302.988
R292 B.n169 B.t3 302.988
R293 B.n30 B.t6 302.988
R294 B.n22 B.t9 302.988
R295 B.n369 B.n368 256.663
R296 B.n368 B.n367 235.042
R297 B.n368 B.n2 235.042
R298 B.n135 B.n134 163.367
R299 B.n135 B.n84 163.367
R300 B.n139 B.n84 163.367
R301 B.n140 B.n139 163.367
R302 B.n141 B.n140 163.367
R303 B.n141 B.n82 163.367
R304 B.n145 B.n82 163.367
R305 B.n146 B.n145 163.367
R306 B.n147 B.n146 163.367
R307 B.n147 B.n80 163.367
R308 B.n151 B.n80 163.367
R309 B.n152 B.n151 163.367
R310 B.n153 B.n152 163.367
R311 B.n153 B.n76 163.367
R312 B.n158 B.n76 163.367
R313 B.n159 B.n158 163.367
R314 B.n160 B.n159 163.367
R315 B.n160 B.n74 163.367
R316 B.n164 B.n74 163.367
R317 B.n165 B.n164 163.367
R318 B.n166 B.n165 163.367
R319 B.n166 B.n72 163.367
R320 B.n173 B.n72 163.367
R321 B.n174 B.n173 163.367
R322 B.n175 B.n174 163.367
R323 B.n175 B.n70 163.367
R324 B.n179 B.n70 163.367
R325 B.n180 B.n179 163.367
R326 B.n181 B.n180 163.367
R327 B.n181 B.n68 163.367
R328 B.n185 B.n68 163.367
R329 B.n186 B.n185 163.367
R330 B.n187 B.n186 163.367
R331 B.n187 B.n66 163.367
R332 B.n191 B.n66 163.367
R333 B.n192 B.n191 163.367
R334 B.n193 B.n192 163.367
R335 B.n271 B.n270 163.367
R336 B.n270 B.n269 163.367
R337 B.n269 B.n40 163.367
R338 B.n265 B.n40 163.367
R339 B.n265 B.n264 163.367
R340 B.n264 B.n263 163.367
R341 B.n263 B.n42 163.367
R342 B.n259 B.n42 163.367
R343 B.n259 B.n258 163.367
R344 B.n258 B.n257 163.367
R345 B.n257 B.n44 163.367
R346 B.n253 B.n44 163.367
R347 B.n253 B.n252 163.367
R348 B.n252 B.n251 163.367
R349 B.n251 B.n46 163.367
R350 B.n247 B.n46 163.367
R351 B.n247 B.n246 163.367
R352 B.n246 B.n245 163.367
R353 B.n245 B.n48 163.367
R354 B.n241 B.n48 163.367
R355 B.n241 B.n240 163.367
R356 B.n240 B.n239 163.367
R357 B.n239 B.n50 163.367
R358 B.n235 B.n50 163.367
R359 B.n235 B.n234 163.367
R360 B.n234 B.n233 163.367
R361 B.n233 B.n52 163.367
R362 B.n229 B.n52 163.367
R363 B.n229 B.n228 163.367
R364 B.n228 B.n227 163.367
R365 B.n227 B.n54 163.367
R366 B.n223 B.n54 163.367
R367 B.n223 B.n222 163.367
R368 B.n222 B.n221 163.367
R369 B.n221 B.n56 163.367
R370 B.n217 B.n56 163.367
R371 B.n217 B.n216 163.367
R372 B.n216 B.n215 163.367
R373 B.n215 B.n58 163.367
R374 B.n211 B.n58 163.367
R375 B.n211 B.n210 163.367
R376 B.n210 B.n209 163.367
R377 B.n209 B.n60 163.367
R378 B.n205 B.n60 163.367
R379 B.n205 B.n204 163.367
R380 B.n204 B.n203 163.367
R381 B.n203 B.n62 163.367
R382 B.n199 B.n62 163.367
R383 B.n199 B.n198 163.367
R384 B.n198 B.n197 163.367
R385 B.n197 B.n64 163.367
R386 B.n330 B.n15 163.367
R387 B.n326 B.n15 163.367
R388 B.n326 B.n325 163.367
R389 B.n325 B.n324 163.367
R390 B.n324 B.n17 163.367
R391 B.n320 B.n17 163.367
R392 B.n320 B.n319 163.367
R393 B.n319 B.n318 163.367
R394 B.n318 B.n19 163.367
R395 B.n314 B.n19 163.367
R396 B.n314 B.n313 163.367
R397 B.n313 B.n312 163.367
R398 B.n312 B.n21 163.367
R399 B.n307 B.n21 163.367
R400 B.n307 B.n306 163.367
R401 B.n306 B.n305 163.367
R402 B.n305 B.n25 163.367
R403 B.n301 B.n25 163.367
R404 B.n301 B.n300 163.367
R405 B.n300 B.n299 163.367
R406 B.n299 B.n27 163.367
R407 B.n295 B.n27 163.367
R408 B.n295 B.n294 163.367
R409 B.n294 B.n293 163.367
R410 B.n293 B.n29 163.367
R411 B.n289 B.n29 163.367
R412 B.n289 B.n288 163.367
R413 B.n288 B.n287 163.367
R414 B.n287 B.n34 163.367
R415 B.n283 B.n34 163.367
R416 B.n283 B.n282 163.367
R417 B.n282 B.n281 163.367
R418 B.n281 B.n36 163.367
R419 B.n277 B.n36 163.367
R420 B.n277 B.n276 163.367
R421 B.n276 B.n275 163.367
R422 B.n275 B.n38 163.367
R423 B.n332 B.n331 163.367
R424 B.n332 B.n13 163.367
R425 B.n336 B.n13 163.367
R426 B.n337 B.n336 163.367
R427 B.n338 B.n337 163.367
R428 B.n338 B.n11 163.367
R429 B.n342 B.n11 163.367
R430 B.n343 B.n342 163.367
R431 B.n344 B.n343 163.367
R432 B.n344 B.n9 163.367
R433 B.n348 B.n9 163.367
R434 B.n349 B.n348 163.367
R435 B.n350 B.n349 163.367
R436 B.n350 B.n7 163.367
R437 B.n354 B.n7 163.367
R438 B.n355 B.n354 163.367
R439 B.n356 B.n355 163.367
R440 B.n356 B.n5 163.367
R441 B.n360 B.n5 163.367
R442 B.n361 B.n360 163.367
R443 B.n362 B.n361 163.367
R444 B.n362 B.n3 163.367
R445 B.n366 B.n3 163.367
R446 B.n367 B.n366 163.367
R447 B.n98 B.n2 163.367
R448 B.n99 B.n98 163.367
R449 B.n99 B.n96 163.367
R450 B.n103 B.n96 163.367
R451 B.n104 B.n103 163.367
R452 B.n105 B.n104 163.367
R453 B.n105 B.n94 163.367
R454 B.n109 B.n94 163.367
R455 B.n110 B.n109 163.367
R456 B.n111 B.n110 163.367
R457 B.n111 B.n92 163.367
R458 B.n115 B.n92 163.367
R459 B.n116 B.n115 163.367
R460 B.n117 B.n116 163.367
R461 B.n117 B.n90 163.367
R462 B.n121 B.n90 163.367
R463 B.n122 B.n121 163.367
R464 B.n123 B.n122 163.367
R465 B.n123 B.n88 163.367
R466 B.n127 B.n88 163.367
R467 B.n128 B.n127 163.367
R468 B.n129 B.n128 163.367
R469 B.n129 B.n86 163.367
R470 B.n133 B.n86 163.367
R471 B.n169 B.t4 161.055
R472 B.n30 B.t8 161.055
R473 B.n77 B.t1 161.054
R474 B.n22 B.t11 161.054
R475 B.n170 B.t5 141.661
R476 B.n31 B.t7 141.661
R477 B.n78 B.t2 141.661
R478 B.n23 B.t10 141.661
R479 B.n155 B.n78 59.5399
R480 B.n171 B.n170 59.5399
R481 B.n32 B.n31 59.5399
R482 B.n309 B.n23 59.5399
R483 B.n329 B.n14 37.9322
R484 B.n273 B.n272 37.9322
R485 B.n195 B.n194 37.9322
R486 B.n132 B.n85 37.9322
R487 B.n78 B.n77 19.3944
R488 B.n170 B.n169 19.3944
R489 B.n31 B.n30 19.3944
R490 B.n23 B.n22 19.3944
R491 B B.n369 18.0485
R492 B.n333 B.n14 10.6151
R493 B.n334 B.n333 10.6151
R494 B.n335 B.n334 10.6151
R495 B.n335 B.n12 10.6151
R496 B.n339 B.n12 10.6151
R497 B.n340 B.n339 10.6151
R498 B.n341 B.n340 10.6151
R499 B.n341 B.n10 10.6151
R500 B.n345 B.n10 10.6151
R501 B.n346 B.n345 10.6151
R502 B.n347 B.n346 10.6151
R503 B.n347 B.n8 10.6151
R504 B.n351 B.n8 10.6151
R505 B.n352 B.n351 10.6151
R506 B.n353 B.n352 10.6151
R507 B.n353 B.n6 10.6151
R508 B.n357 B.n6 10.6151
R509 B.n358 B.n357 10.6151
R510 B.n359 B.n358 10.6151
R511 B.n359 B.n4 10.6151
R512 B.n363 B.n4 10.6151
R513 B.n364 B.n363 10.6151
R514 B.n365 B.n364 10.6151
R515 B.n365 B.n0 10.6151
R516 B.n329 B.n328 10.6151
R517 B.n328 B.n327 10.6151
R518 B.n327 B.n16 10.6151
R519 B.n323 B.n16 10.6151
R520 B.n323 B.n322 10.6151
R521 B.n322 B.n321 10.6151
R522 B.n321 B.n18 10.6151
R523 B.n317 B.n18 10.6151
R524 B.n317 B.n316 10.6151
R525 B.n316 B.n315 10.6151
R526 B.n315 B.n20 10.6151
R527 B.n311 B.n20 10.6151
R528 B.n311 B.n310 10.6151
R529 B.n308 B.n24 10.6151
R530 B.n304 B.n24 10.6151
R531 B.n304 B.n303 10.6151
R532 B.n303 B.n302 10.6151
R533 B.n302 B.n26 10.6151
R534 B.n298 B.n26 10.6151
R535 B.n298 B.n297 10.6151
R536 B.n297 B.n296 10.6151
R537 B.n296 B.n28 10.6151
R538 B.n292 B.n291 10.6151
R539 B.n291 B.n290 10.6151
R540 B.n290 B.n33 10.6151
R541 B.n286 B.n33 10.6151
R542 B.n286 B.n285 10.6151
R543 B.n285 B.n284 10.6151
R544 B.n284 B.n35 10.6151
R545 B.n280 B.n35 10.6151
R546 B.n280 B.n279 10.6151
R547 B.n279 B.n278 10.6151
R548 B.n278 B.n37 10.6151
R549 B.n274 B.n37 10.6151
R550 B.n274 B.n273 10.6151
R551 B.n272 B.n39 10.6151
R552 B.n268 B.n39 10.6151
R553 B.n268 B.n267 10.6151
R554 B.n267 B.n266 10.6151
R555 B.n266 B.n41 10.6151
R556 B.n262 B.n41 10.6151
R557 B.n262 B.n261 10.6151
R558 B.n261 B.n260 10.6151
R559 B.n260 B.n43 10.6151
R560 B.n256 B.n43 10.6151
R561 B.n256 B.n255 10.6151
R562 B.n255 B.n254 10.6151
R563 B.n254 B.n45 10.6151
R564 B.n250 B.n45 10.6151
R565 B.n250 B.n249 10.6151
R566 B.n249 B.n248 10.6151
R567 B.n248 B.n47 10.6151
R568 B.n244 B.n47 10.6151
R569 B.n244 B.n243 10.6151
R570 B.n243 B.n242 10.6151
R571 B.n242 B.n49 10.6151
R572 B.n238 B.n49 10.6151
R573 B.n238 B.n237 10.6151
R574 B.n237 B.n236 10.6151
R575 B.n236 B.n51 10.6151
R576 B.n232 B.n51 10.6151
R577 B.n232 B.n231 10.6151
R578 B.n231 B.n230 10.6151
R579 B.n230 B.n53 10.6151
R580 B.n226 B.n53 10.6151
R581 B.n226 B.n225 10.6151
R582 B.n225 B.n224 10.6151
R583 B.n224 B.n55 10.6151
R584 B.n220 B.n55 10.6151
R585 B.n220 B.n219 10.6151
R586 B.n219 B.n218 10.6151
R587 B.n218 B.n57 10.6151
R588 B.n214 B.n57 10.6151
R589 B.n214 B.n213 10.6151
R590 B.n213 B.n212 10.6151
R591 B.n212 B.n59 10.6151
R592 B.n208 B.n59 10.6151
R593 B.n208 B.n207 10.6151
R594 B.n207 B.n206 10.6151
R595 B.n206 B.n61 10.6151
R596 B.n202 B.n61 10.6151
R597 B.n202 B.n201 10.6151
R598 B.n201 B.n200 10.6151
R599 B.n200 B.n63 10.6151
R600 B.n196 B.n63 10.6151
R601 B.n196 B.n195 10.6151
R602 B.n97 B.n1 10.6151
R603 B.n100 B.n97 10.6151
R604 B.n101 B.n100 10.6151
R605 B.n102 B.n101 10.6151
R606 B.n102 B.n95 10.6151
R607 B.n106 B.n95 10.6151
R608 B.n107 B.n106 10.6151
R609 B.n108 B.n107 10.6151
R610 B.n108 B.n93 10.6151
R611 B.n112 B.n93 10.6151
R612 B.n113 B.n112 10.6151
R613 B.n114 B.n113 10.6151
R614 B.n114 B.n91 10.6151
R615 B.n118 B.n91 10.6151
R616 B.n119 B.n118 10.6151
R617 B.n120 B.n119 10.6151
R618 B.n120 B.n89 10.6151
R619 B.n124 B.n89 10.6151
R620 B.n125 B.n124 10.6151
R621 B.n126 B.n125 10.6151
R622 B.n126 B.n87 10.6151
R623 B.n130 B.n87 10.6151
R624 B.n131 B.n130 10.6151
R625 B.n132 B.n131 10.6151
R626 B.n136 B.n85 10.6151
R627 B.n137 B.n136 10.6151
R628 B.n138 B.n137 10.6151
R629 B.n138 B.n83 10.6151
R630 B.n142 B.n83 10.6151
R631 B.n143 B.n142 10.6151
R632 B.n144 B.n143 10.6151
R633 B.n144 B.n81 10.6151
R634 B.n148 B.n81 10.6151
R635 B.n149 B.n148 10.6151
R636 B.n150 B.n149 10.6151
R637 B.n150 B.n79 10.6151
R638 B.n154 B.n79 10.6151
R639 B.n157 B.n156 10.6151
R640 B.n157 B.n75 10.6151
R641 B.n161 B.n75 10.6151
R642 B.n162 B.n161 10.6151
R643 B.n163 B.n162 10.6151
R644 B.n163 B.n73 10.6151
R645 B.n167 B.n73 10.6151
R646 B.n168 B.n167 10.6151
R647 B.n172 B.n168 10.6151
R648 B.n176 B.n71 10.6151
R649 B.n177 B.n176 10.6151
R650 B.n178 B.n177 10.6151
R651 B.n178 B.n69 10.6151
R652 B.n182 B.n69 10.6151
R653 B.n183 B.n182 10.6151
R654 B.n184 B.n183 10.6151
R655 B.n184 B.n67 10.6151
R656 B.n188 B.n67 10.6151
R657 B.n189 B.n188 10.6151
R658 B.n190 B.n189 10.6151
R659 B.n190 B.n65 10.6151
R660 B.n194 B.n65 10.6151
R661 B.n310 B.n309 9.36635
R662 B.n292 B.n32 9.36635
R663 B.n155 B.n154 9.36635
R664 B.n171 B.n71 9.36635
R665 B.n369 B.n0 8.11757
R666 B.n369 B.n1 8.11757
R667 B.n309 B.n308 1.24928
R668 B.n32 B.n28 1.24928
R669 B.n156 B.n155 1.24928
R670 B.n172 B.n171 1.24928
R671 VP.n7 VP.t9 179.625
R672 VP.n31 VP.n30 161.3
R673 VP.n10 VP.n9 161.3
R674 VP.n11 VP.n6 161.3
R675 VP.n13 VP.n12 161.3
R676 VP.n14 VP.n5 161.3
R677 VP.n15 VP.n4 161.3
R678 VP.n17 VP.n16 161.3
R679 VP.n29 VP.n0 161.3
R680 VP.n28 VP.n27 161.3
R681 VP.n26 VP.n1 161.3
R682 VP.n25 VP.n24 161.3
R683 VP.n23 VP.n2 161.3
R684 VP.n22 VP.n21 161.3
R685 VP.n20 VP.n3 161.3
R686 VP.n19 VP.n18 161.3
R687 VP.n18 VP.t4 158.629
R688 VP.n22 VP.t8 158.629
R689 VP.n24 VP.t2 158.629
R690 VP.n28 VP.t7 158.629
R691 VP.n30 VP.t1 158.629
R692 VP.n16 VP.t5 158.629
R693 VP.n14 VP.t0 158.629
R694 VP.n6 VP.t6 158.629
R695 VP.n8 VP.t3 158.629
R696 VP.n10 VP.n7 44.8515
R697 VP.n19 VP.n17 35.5763
R698 VP.n18 VP.n3 24.1005
R699 VP.n22 VP.n3 24.1005
R700 VP.n23 VP.n22 24.1005
R701 VP.n24 VP.n23 24.1005
R702 VP.n24 VP.n1 24.1005
R703 VP.n28 VP.n1 24.1005
R704 VP.n29 VP.n28 24.1005
R705 VP.n30 VP.n29 24.1005
R706 VP.n15 VP.n14 24.1005
R707 VP.n16 VP.n15 24.1005
R708 VP.n13 VP.n6 24.1005
R709 VP.n14 VP.n13 24.1005
R710 VP.n9 VP.n8 24.1005
R711 VP.n9 VP.n6 24.1005
R712 VP.n8 VP.n7 20.9471
R713 VP.n11 VP.n10 0.189894
R714 VP.n12 VP.n11 0.189894
R715 VP.n12 VP.n5 0.189894
R716 VP.n5 VP.n4 0.189894
R717 VP.n17 VP.n4 0.189894
R718 VP.n20 VP.n19 0.189894
R719 VP.n21 VP.n20 0.189894
R720 VP.n21 VP.n2 0.189894
R721 VP.n25 VP.n2 0.189894
R722 VP.n26 VP.n25 0.189894
R723 VP.n27 VP.n26 0.189894
R724 VP.n27 VP.n0 0.189894
R725 VP.n31 VP.n0 0.189894
R726 VP VP.n31 0.0516364
R727 VDD1.n1 VDD1.t0 150.861
R728 VDD1.n3 VDD1.t5 150.861
R729 VDD1.n5 VDD1.n4 138.856
R730 VDD1.n1 VDD1.n0 138.264
R731 VDD1.n7 VDD1.n6 138.264
R732 VDD1.n3 VDD1.n2 138.263
R733 VDD1.n7 VDD1.n5 31.2121
R734 VDD1.n6 VDD1.t9 11.7352
R735 VDD1.n6 VDD1.t4 11.7352
R736 VDD1.n0 VDD1.t6 11.7352
R737 VDD1.n0 VDD1.t3 11.7352
R738 VDD1.n4 VDD1.t2 11.7352
R739 VDD1.n4 VDD1.t8 11.7352
R740 VDD1.n2 VDD1.t1 11.7352
R741 VDD1.n2 VDD1.t7 11.7352
R742 VDD1 VDD1.n7 0.588862
R743 VDD1 VDD1.n1 0.274207
R744 VDD1.n5 VDD1.n3 0.160671
C0 VDD1 VN 0.153921f
C1 w_n2170_n1522# B 4.7132f
C2 VDD1 VP 2.03619f
C3 VDD1 VDD2 0.947807f
C4 VTAIL VN 2.13554f
C5 VTAIL VP 2.14976f
C6 VTAIL VDD2 5.2945f
C7 VN B 0.679935f
C8 VN w_n2170_n1522# 3.88148f
C9 VP B 1.13386f
C10 VDD2 B 1.06222f
C11 VTAIL VDD1 5.2554f
C12 VP w_n2170_n1522# 4.15533f
C13 VDD2 w_n2170_n1522# 1.37668f
C14 VDD1 B 1.019f
C15 VDD1 w_n2170_n1522# 1.33418f
C16 VP VN 3.85378f
C17 VDD2 VN 1.85034f
C18 VTAIL B 1.04922f
C19 VDD2 VP 0.341882f
C20 VTAIL w_n2170_n1522# 1.53023f
C21 VDD2 VSUBS 0.811569f
C22 VDD1 VSUBS 0.847012f
C23 VTAIL VSUBS 0.349668f
C24 VN VSUBS 3.99088f
C25 VP VSUBS 1.318763f
C26 B VSUBS 2.093441f
C27 w_n2170_n1522# VSUBS 41.8984f
C28 VDD1.t0 VSUBS 0.402593f
C29 VDD1.t6 VSUBS 0.054758f
C30 VDD1.t3 VSUBS 0.054758f
C31 VDD1.n0 VSUBS 0.280212f
C32 VDD1.n1 VSUBS 0.807021f
C33 VDD1.t5 VSUBS 0.402592f
C34 VDD1.t1 VSUBS 0.054758f
C35 VDD1.t7 VSUBS 0.054758f
C36 VDD1.n2 VSUBS 0.280211f
C37 VDD1.n3 VSUBS 0.801492f
C38 VDD1.t2 VSUBS 0.054758f
C39 VDD1.t8 VSUBS 0.054758f
C40 VDD1.n4 VSUBS 0.282053f
C41 VDD1.n5 VSUBS 1.51949f
C42 VDD1.t9 VSUBS 0.054758f
C43 VDD1.t4 VSUBS 0.054758f
C44 VDD1.n6 VSUBS 0.280211f
C45 VDD1.n7 VSUBS 1.73657f
C46 VP.n0 VSUBS 0.071708f
C47 VP.n1 VSUBS 0.016272f
C48 VP.n2 VSUBS 0.071708f
C49 VP.n3 VSUBS 0.016272f
C50 VP.n4 VSUBS 0.071708f
C51 VP.t5 VSUBS 0.401684f
C52 VP.t0 VSUBS 0.401684f
C53 VP.n5 VSUBS 0.071708f
C54 VP.t6 VSUBS 0.401684f
C55 VP.n6 VSUBS 0.243818f
C56 VP.t9 VSUBS 0.429967f
C57 VP.n7 VSUBS 0.220758f
C58 VP.t3 VSUBS 0.401684f
C59 VP.n8 VSUBS 0.248983f
C60 VP.n9 VSUBS 0.016272f
C61 VP.n10 VSUBS 0.292937f
C62 VP.n11 VSUBS 0.071708f
C63 VP.n12 VSUBS 0.071708f
C64 VP.n13 VSUBS 0.016272f
C65 VP.n14 VSUBS 0.243818f
C66 VP.n15 VSUBS 0.016272f
C67 VP.n16 VSUBS 0.236523f
C68 VP.n17 VSUBS 2.20458f
C69 VP.t4 VSUBS 0.401684f
C70 VP.n18 VSUBS 0.236523f
C71 VP.n19 VSUBS 2.27704f
C72 VP.n20 VSUBS 0.071708f
C73 VP.n21 VSUBS 0.071708f
C74 VP.t8 VSUBS 0.401684f
C75 VP.n22 VSUBS 0.243818f
C76 VP.n23 VSUBS 0.016272f
C77 VP.t2 VSUBS 0.401684f
C78 VP.n24 VSUBS 0.243818f
C79 VP.n25 VSUBS 0.071708f
C80 VP.n26 VSUBS 0.071708f
C81 VP.n27 VSUBS 0.071708f
C82 VP.t7 VSUBS 0.401684f
C83 VP.n28 VSUBS 0.243818f
C84 VP.n29 VSUBS 0.016272f
C85 VP.t1 VSUBS 0.401684f
C86 VP.n30 VSUBS 0.236523f
C87 VP.n31 VSUBS 0.055571f
C88 B.n0 VSUBS 0.007049f
C89 B.n1 VSUBS 0.007049f
C90 B.n2 VSUBS 0.010425f
C91 B.n3 VSUBS 0.007989f
C92 B.n4 VSUBS 0.007989f
C93 B.n5 VSUBS 0.007989f
C94 B.n6 VSUBS 0.007989f
C95 B.n7 VSUBS 0.007989f
C96 B.n8 VSUBS 0.007989f
C97 B.n9 VSUBS 0.007989f
C98 B.n10 VSUBS 0.007989f
C99 B.n11 VSUBS 0.007989f
C100 B.n12 VSUBS 0.007989f
C101 B.n13 VSUBS 0.007989f
C102 B.n14 VSUBS 0.02029f
C103 B.n15 VSUBS 0.007989f
C104 B.n16 VSUBS 0.007989f
C105 B.n17 VSUBS 0.007989f
C106 B.n18 VSUBS 0.007989f
C107 B.n19 VSUBS 0.007989f
C108 B.n20 VSUBS 0.007989f
C109 B.n21 VSUBS 0.007989f
C110 B.t10 VSUBS 0.074584f
C111 B.t11 VSUBS 0.08088f
C112 B.t9 VSUBS 0.097425f
C113 B.n22 VSUBS 0.070615f
C114 B.n23 VSUBS 0.063679f
C115 B.n24 VSUBS 0.007989f
C116 B.n25 VSUBS 0.007989f
C117 B.n26 VSUBS 0.007989f
C118 B.n27 VSUBS 0.007989f
C119 B.n28 VSUBS 0.004464f
C120 B.n29 VSUBS 0.007989f
C121 B.t7 VSUBS 0.074584f
C122 B.t8 VSUBS 0.08088f
C123 B.t6 VSUBS 0.097425f
C124 B.n30 VSUBS 0.070615f
C125 B.n31 VSUBS 0.063679f
C126 B.n32 VSUBS 0.018509f
C127 B.n33 VSUBS 0.007989f
C128 B.n34 VSUBS 0.007989f
C129 B.n35 VSUBS 0.007989f
C130 B.n36 VSUBS 0.007989f
C131 B.n37 VSUBS 0.007989f
C132 B.n38 VSUBS 0.021063f
C133 B.n39 VSUBS 0.007989f
C134 B.n40 VSUBS 0.007989f
C135 B.n41 VSUBS 0.007989f
C136 B.n42 VSUBS 0.007989f
C137 B.n43 VSUBS 0.007989f
C138 B.n44 VSUBS 0.007989f
C139 B.n45 VSUBS 0.007989f
C140 B.n46 VSUBS 0.007989f
C141 B.n47 VSUBS 0.007989f
C142 B.n48 VSUBS 0.007989f
C143 B.n49 VSUBS 0.007989f
C144 B.n50 VSUBS 0.007989f
C145 B.n51 VSUBS 0.007989f
C146 B.n52 VSUBS 0.007989f
C147 B.n53 VSUBS 0.007989f
C148 B.n54 VSUBS 0.007989f
C149 B.n55 VSUBS 0.007989f
C150 B.n56 VSUBS 0.007989f
C151 B.n57 VSUBS 0.007989f
C152 B.n58 VSUBS 0.007989f
C153 B.n59 VSUBS 0.007989f
C154 B.n60 VSUBS 0.007989f
C155 B.n61 VSUBS 0.007989f
C156 B.n62 VSUBS 0.007989f
C157 B.n63 VSUBS 0.007989f
C158 B.n64 VSUBS 0.02029f
C159 B.n65 VSUBS 0.007989f
C160 B.n66 VSUBS 0.007989f
C161 B.n67 VSUBS 0.007989f
C162 B.n68 VSUBS 0.007989f
C163 B.n69 VSUBS 0.007989f
C164 B.n70 VSUBS 0.007989f
C165 B.n71 VSUBS 0.007519f
C166 B.n72 VSUBS 0.007989f
C167 B.n73 VSUBS 0.007989f
C168 B.n74 VSUBS 0.007989f
C169 B.n75 VSUBS 0.007989f
C170 B.n76 VSUBS 0.007989f
C171 B.t2 VSUBS 0.074584f
C172 B.t1 VSUBS 0.08088f
C173 B.t0 VSUBS 0.097425f
C174 B.n77 VSUBS 0.070615f
C175 B.n78 VSUBS 0.063679f
C176 B.n79 VSUBS 0.007989f
C177 B.n80 VSUBS 0.007989f
C178 B.n81 VSUBS 0.007989f
C179 B.n82 VSUBS 0.007989f
C180 B.n83 VSUBS 0.007989f
C181 B.n84 VSUBS 0.007989f
C182 B.n85 VSUBS 0.021063f
C183 B.n86 VSUBS 0.007989f
C184 B.n87 VSUBS 0.007989f
C185 B.n88 VSUBS 0.007989f
C186 B.n89 VSUBS 0.007989f
C187 B.n90 VSUBS 0.007989f
C188 B.n91 VSUBS 0.007989f
C189 B.n92 VSUBS 0.007989f
C190 B.n93 VSUBS 0.007989f
C191 B.n94 VSUBS 0.007989f
C192 B.n95 VSUBS 0.007989f
C193 B.n96 VSUBS 0.007989f
C194 B.n97 VSUBS 0.007989f
C195 B.n98 VSUBS 0.007989f
C196 B.n99 VSUBS 0.007989f
C197 B.n100 VSUBS 0.007989f
C198 B.n101 VSUBS 0.007989f
C199 B.n102 VSUBS 0.007989f
C200 B.n103 VSUBS 0.007989f
C201 B.n104 VSUBS 0.007989f
C202 B.n105 VSUBS 0.007989f
C203 B.n106 VSUBS 0.007989f
C204 B.n107 VSUBS 0.007989f
C205 B.n108 VSUBS 0.007989f
C206 B.n109 VSUBS 0.007989f
C207 B.n110 VSUBS 0.007989f
C208 B.n111 VSUBS 0.007989f
C209 B.n112 VSUBS 0.007989f
C210 B.n113 VSUBS 0.007989f
C211 B.n114 VSUBS 0.007989f
C212 B.n115 VSUBS 0.007989f
C213 B.n116 VSUBS 0.007989f
C214 B.n117 VSUBS 0.007989f
C215 B.n118 VSUBS 0.007989f
C216 B.n119 VSUBS 0.007989f
C217 B.n120 VSUBS 0.007989f
C218 B.n121 VSUBS 0.007989f
C219 B.n122 VSUBS 0.007989f
C220 B.n123 VSUBS 0.007989f
C221 B.n124 VSUBS 0.007989f
C222 B.n125 VSUBS 0.007989f
C223 B.n126 VSUBS 0.007989f
C224 B.n127 VSUBS 0.007989f
C225 B.n128 VSUBS 0.007989f
C226 B.n129 VSUBS 0.007989f
C227 B.n130 VSUBS 0.007989f
C228 B.n131 VSUBS 0.007989f
C229 B.n132 VSUBS 0.02029f
C230 B.n133 VSUBS 0.02029f
C231 B.n134 VSUBS 0.021063f
C232 B.n135 VSUBS 0.007989f
C233 B.n136 VSUBS 0.007989f
C234 B.n137 VSUBS 0.007989f
C235 B.n138 VSUBS 0.007989f
C236 B.n139 VSUBS 0.007989f
C237 B.n140 VSUBS 0.007989f
C238 B.n141 VSUBS 0.007989f
C239 B.n142 VSUBS 0.007989f
C240 B.n143 VSUBS 0.007989f
C241 B.n144 VSUBS 0.007989f
C242 B.n145 VSUBS 0.007989f
C243 B.n146 VSUBS 0.007989f
C244 B.n147 VSUBS 0.007989f
C245 B.n148 VSUBS 0.007989f
C246 B.n149 VSUBS 0.007989f
C247 B.n150 VSUBS 0.007989f
C248 B.n151 VSUBS 0.007989f
C249 B.n152 VSUBS 0.007989f
C250 B.n153 VSUBS 0.007989f
C251 B.n154 VSUBS 0.007519f
C252 B.n155 VSUBS 0.018509f
C253 B.n156 VSUBS 0.004464f
C254 B.n157 VSUBS 0.007989f
C255 B.n158 VSUBS 0.007989f
C256 B.n159 VSUBS 0.007989f
C257 B.n160 VSUBS 0.007989f
C258 B.n161 VSUBS 0.007989f
C259 B.n162 VSUBS 0.007989f
C260 B.n163 VSUBS 0.007989f
C261 B.n164 VSUBS 0.007989f
C262 B.n165 VSUBS 0.007989f
C263 B.n166 VSUBS 0.007989f
C264 B.n167 VSUBS 0.007989f
C265 B.n168 VSUBS 0.007989f
C266 B.t5 VSUBS 0.074584f
C267 B.t4 VSUBS 0.08088f
C268 B.t3 VSUBS 0.097425f
C269 B.n169 VSUBS 0.070615f
C270 B.n170 VSUBS 0.063679f
C271 B.n171 VSUBS 0.018509f
C272 B.n172 VSUBS 0.004464f
C273 B.n173 VSUBS 0.007989f
C274 B.n174 VSUBS 0.007989f
C275 B.n175 VSUBS 0.007989f
C276 B.n176 VSUBS 0.007989f
C277 B.n177 VSUBS 0.007989f
C278 B.n178 VSUBS 0.007989f
C279 B.n179 VSUBS 0.007989f
C280 B.n180 VSUBS 0.007989f
C281 B.n181 VSUBS 0.007989f
C282 B.n182 VSUBS 0.007989f
C283 B.n183 VSUBS 0.007989f
C284 B.n184 VSUBS 0.007989f
C285 B.n185 VSUBS 0.007989f
C286 B.n186 VSUBS 0.007989f
C287 B.n187 VSUBS 0.007989f
C288 B.n188 VSUBS 0.007989f
C289 B.n189 VSUBS 0.007989f
C290 B.n190 VSUBS 0.007989f
C291 B.n191 VSUBS 0.007989f
C292 B.n192 VSUBS 0.007989f
C293 B.n193 VSUBS 0.021063f
C294 B.n194 VSUBS 0.02025f
C295 B.n195 VSUBS 0.021102f
C296 B.n196 VSUBS 0.007989f
C297 B.n197 VSUBS 0.007989f
C298 B.n198 VSUBS 0.007989f
C299 B.n199 VSUBS 0.007989f
C300 B.n200 VSUBS 0.007989f
C301 B.n201 VSUBS 0.007989f
C302 B.n202 VSUBS 0.007989f
C303 B.n203 VSUBS 0.007989f
C304 B.n204 VSUBS 0.007989f
C305 B.n205 VSUBS 0.007989f
C306 B.n206 VSUBS 0.007989f
C307 B.n207 VSUBS 0.007989f
C308 B.n208 VSUBS 0.007989f
C309 B.n209 VSUBS 0.007989f
C310 B.n210 VSUBS 0.007989f
C311 B.n211 VSUBS 0.007989f
C312 B.n212 VSUBS 0.007989f
C313 B.n213 VSUBS 0.007989f
C314 B.n214 VSUBS 0.007989f
C315 B.n215 VSUBS 0.007989f
C316 B.n216 VSUBS 0.007989f
C317 B.n217 VSUBS 0.007989f
C318 B.n218 VSUBS 0.007989f
C319 B.n219 VSUBS 0.007989f
C320 B.n220 VSUBS 0.007989f
C321 B.n221 VSUBS 0.007989f
C322 B.n222 VSUBS 0.007989f
C323 B.n223 VSUBS 0.007989f
C324 B.n224 VSUBS 0.007989f
C325 B.n225 VSUBS 0.007989f
C326 B.n226 VSUBS 0.007989f
C327 B.n227 VSUBS 0.007989f
C328 B.n228 VSUBS 0.007989f
C329 B.n229 VSUBS 0.007989f
C330 B.n230 VSUBS 0.007989f
C331 B.n231 VSUBS 0.007989f
C332 B.n232 VSUBS 0.007989f
C333 B.n233 VSUBS 0.007989f
C334 B.n234 VSUBS 0.007989f
C335 B.n235 VSUBS 0.007989f
C336 B.n236 VSUBS 0.007989f
C337 B.n237 VSUBS 0.007989f
C338 B.n238 VSUBS 0.007989f
C339 B.n239 VSUBS 0.007989f
C340 B.n240 VSUBS 0.007989f
C341 B.n241 VSUBS 0.007989f
C342 B.n242 VSUBS 0.007989f
C343 B.n243 VSUBS 0.007989f
C344 B.n244 VSUBS 0.007989f
C345 B.n245 VSUBS 0.007989f
C346 B.n246 VSUBS 0.007989f
C347 B.n247 VSUBS 0.007989f
C348 B.n248 VSUBS 0.007989f
C349 B.n249 VSUBS 0.007989f
C350 B.n250 VSUBS 0.007989f
C351 B.n251 VSUBS 0.007989f
C352 B.n252 VSUBS 0.007989f
C353 B.n253 VSUBS 0.007989f
C354 B.n254 VSUBS 0.007989f
C355 B.n255 VSUBS 0.007989f
C356 B.n256 VSUBS 0.007989f
C357 B.n257 VSUBS 0.007989f
C358 B.n258 VSUBS 0.007989f
C359 B.n259 VSUBS 0.007989f
C360 B.n260 VSUBS 0.007989f
C361 B.n261 VSUBS 0.007989f
C362 B.n262 VSUBS 0.007989f
C363 B.n263 VSUBS 0.007989f
C364 B.n264 VSUBS 0.007989f
C365 B.n265 VSUBS 0.007989f
C366 B.n266 VSUBS 0.007989f
C367 B.n267 VSUBS 0.007989f
C368 B.n268 VSUBS 0.007989f
C369 B.n269 VSUBS 0.007989f
C370 B.n270 VSUBS 0.007989f
C371 B.n271 VSUBS 0.02029f
C372 B.n272 VSUBS 0.02029f
C373 B.n273 VSUBS 0.021063f
C374 B.n274 VSUBS 0.007989f
C375 B.n275 VSUBS 0.007989f
C376 B.n276 VSUBS 0.007989f
C377 B.n277 VSUBS 0.007989f
C378 B.n278 VSUBS 0.007989f
C379 B.n279 VSUBS 0.007989f
C380 B.n280 VSUBS 0.007989f
C381 B.n281 VSUBS 0.007989f
C382 B.n282 VSUBS 0.007989f
C383 B.n283 VSUBS 0.007989f
C384 B.n284 VSUBS 0.007989f
C385 B.n285 VSUBS 0.007989f
C386 B.n286 VSUBS 0.007989f
C387 B.n287 VSUBS 0.007989f
C388 B.n288 VSUBS 0.007989f
C389 B.n289 VSUBS 0.007989f
C390 B.n290 VSUBS 0.007989f
C391 B.n291 VSUBS 0.007989f
C392 B.n292 VSUBS 0.007519f
C393 B.n293 VSUBS 0.007989f
C394 B.n294 VSUBS 0.007989f
C395 B.n295 VSUBS 0.007989f
C396 B.n296 VSUBS 0.007989f
C397 B.n297 VSUBS 0.007989f
C398 B.n298 VSUBS 0.007989f
C399 B.n299 VSUBS 0.007989f
C400 B.n300 VSUBS 0.007989f
C401 B.n301 VSUBS 0.007989f
C402 B.n302 VSUBS 0.007989f
C403 B.n303 VSUBS 0.007989f
C404 B.n304 VSUBS 0.007989f
C405 B.n305 VSUBS 0.007989f
C406 B.n306 VSUBS 0.007989f
C407 B.n307 VSUBS 0.007989f
C408 B.n308 VSUBS 0.004464f
C409 B.n309 VSUBS 0.018509f
C410 B.n310 VSUBS 0.007519f
C411 B.n311 VSUBS 0.007989f
C412 B.n312 VSUBS 0.007989f
C413 B.n313 VSUBS 0.007989f
C414 B.n314 VSUBS 0.007989f
C415 B.n315 VSUBS 0.007989f
C416 B.n316 VSUBS 0.007989f
C417 B.n317 VSUBS 0.007989f
C418 B.n318 VSUBS 0.007989f
C419 B.n319 VSUBS 0.007989f
C420 B.n320 VSUBS 0.007989f
C421 B.n321 VSUBS 0.007989f
C422 B.n322 VSUBS 0.007989f
C423 B.n323 VSUBS 0.007989f
C424 B.n324 VSUBS 0.007989f
C425 B.n325 VSUBS 0.007989f
C426 B.n326 VSUBS 0.007989f
C427 B.n327 VSUBS 0.007989f
C428 B.n328 VSUBS 0.007989f
C429 B.n329 VSUBS 0.021063f
C430 B.n330 VSUBS 0.021063f
C431 B.n331 VSUBS 0.02029f
C432 B.n332 VSUBS 0.007989f
C433 B.n333 VSUBS 0.007989f
C434 B.n334 VSUBS 0.007989f
C435 B.n335 VSUBS 0.007989f
C436 B.n336 VSUBS 0.007989f
C437 B.n337 VSUBS 0.007989f
C438 B.n338 VSUBS 0.007989f
C439 B.n339 VSUBS 0.007989f
C440 B.n340 VSUBS 0.007989f
C441 B.n341 VSUBS 0.007989f
C442 B.n342 VSUBS 0.007989f
C443 B.n343 VSUBS 0.007989f
C444 B.n344 VSUBS 0.007989f
C445 B.n345 VSUBS 0.007989f
C446 B.n346 VSUBS 0.007989f
C447 B.n347 VSUBS 0.007989f
C448 B.n348 VSUBS 0.007989f
C449 B.n349 VSUBS 0.007989f
C450 B.n350 VSUBS 0.007989f
C451 B.n351 VSUBS 0.007989f
C452 B.n352 VSUBS 0.007989f
C453 B.n353 VSUBS 0.007989f
C454 B.n354 VSUBS 0.007989f
C455 B.n355 VSUBS 0.007989f
C456 B.n356 VSUBS 0.007989f
C457 B.n357 VSUBS 0.007989f
C458 B.n358 VSUBS 0.007989f
C459 B.n359 VSUBS 0.007989f
C460 B.n360 VSUBS 0.007989f
C461 B.n361 VSUBS 0.007989f
C462 B.n362 VSUBS 0.007989f
C463 B.n363 VSUBS 0.007989f
C464 B.n364 VSUBS 0.007989f
C465 B.n365 VSUBS 0.007989f
C466 B.n366 VSUBS 0.007989f
C467 B.n367 VSUBS 0.010425f
C468 B.n368 VSUBS 0.011105f
C469 B.n369 VSUBS 0.022083f
C470 VDD2.t7 VSUBS 0.29604f
C471 VDD2.t2 VSUBS 0.040265f
C472 VDD2.t6 VSUBS 0.040265f
C473 VDD2.n0 VSUBS 0.206049f
C474 VDD2.n1 VSUBS 0.589365f
C475 VDD2.t0 VSUBS 0.040265f
C476 VDD2.t4 VSUBS 0.040265f
C477 VDD2.n2 VSUBS 0.207403f
C478 VDD2.n3 VSUBS 1.06431f
C479 VDD2.t9 VSUBS 0.294304f
C480 VDD2.n4 VSUBS 1.24873f
C481 VDD2.t3 VSUBS 0.040265f
C482 VDD2.t8 VSUBS 0.040265f
C483 VDD2.n5 VSUBS 0.206049f
C484 VDD2.n6 VSUBS 0.29121f
C485 VDD2.t1 VSUBS 0.040265f
C486 VDD2.t5 VSUBS 0.040265f
C487 VDD2.n7 VSUBS 0.207393f
C488 VTAIL.t10 VSUBS 0.067366f
C489 VTAIL.t8 VSUBS 0.067366f
C490 VTAIL.n0 VSUBS 0.294149f
C491 VTAIL.n1 VSUBS 0.542551f
C492 VTAIL.t0 VSUBS 0.441742f
C493 VTAIL.n2 VSUBS 0.594286f
C494 VTAIL.t19 VSUBS 0.067366f
C495 VTAIL.t7 VSUBS 0.067366f
C496 VTAIL.n3 VSUBS 0.294149f
C497 VTAIL.n4 VSUBS 0.554306f
C498 VTAIL.t1 VSUBS 0.067366f
C499 VTAIL.t6 VSUBS 0.067366f
C500 VTAIL.n5 VSUBS 0.294149f
C501 VTAIL.n6 VSUBS 1.29465f
C502 VTAIL.t17 VSUBS 0.067366f
C503 VTAIL.t14 VSUBS 0.067366f
C504 VTAIL.n7 VSUBS 0.29415f
C505 VTAIL.n8 VSUBS 1.29465f
C506 VTAIL.t13 VSUBS 0.067366f
C507 VTAIL.t9 VSUBS 0.067366f
C508 VTAIL.n9 VSUBS 0.29415f
C509 VTAIL.n10 VSUBS 0.554305f
C510 VTAIL.t15 VSUBS 0.441743f
C511 VTAIL.n11 VSUBS 0.594284f
C512 VTAIL.t4 VSUBS 0.067366f
C513 VTAIL.t2 VSUBS 0.067366f
C514 VTAIL.n12 VSUBS 0.29415f
C515 VTAIL.n13 VSUBS 0.558152f
C516 VTAIL.t3 VSUBS 0.067366f
C517 VTAIL.t5 VSUBS 0.067366f
C518 VTAIL.n14 VSUBS 0.29415f
C519 VTAIL.n15 VSUBS 0.554305f
C520 VTAIL.t18 VSUBS 0.441742f
C521 VTAIL.n16 VSUBS 1.24529f
C522 VTAIL.t16 VSUBS 0.441742f
C523 VTAIL.n17 VSUBS 1.24529f
C524 VTAIL.t12 VSUBS 0.067366f
C525 VTAIL.t11 VSUBS 0.067366f
C526 VTAIL.n18 VSUBS 0.294149f
C527 VTAIL.n19 VSUBS 0.484419f
C528 VN.n0 VSUBS 0.057712f
C529 VN.n1 VSUBS 0.013096f
C530 VN.n2 VSUBS 0.235763f
C531 VN.t2 VSUBS 0.346049f
C532 VN.n3 VSUBS 0.177672f
C533 VN.t7 VSUBS 0.323286f
C534 VN.n4 VSUBS 0.200388f
C535 VN.n5 VSUBS 0.013096f
C536 VN.t3 VSUBS 0.323286f
C537 VN.n6 VSUBS 0.196231f
C538 VN.n7 VSUBS 0.057712f
C539 VN.n8 VSUBS 0.057712f
C540 VN.n9 VSUBS 0.057712f
C541 VN.t9 VSUBS 0.323286f
C542 VN.n10 VSUBS 0.196231f
C543 VN.n11 VSUBS 0.013096f
C544 VN.t5 VSUBS 0.323286f
C545 VN.n12 VSUBS 0.19036f
C546 VN.n13 VSUBS 0.044725f
C547 VN.n14 VSUBS 0.057712f
C548 VN.n15 VSUBS 0.013096f
C549 VN.t6 VSUBS 0.323286f
C550 VN.n16 VSUBS 0.235763f
C551 VN.t4 VSUBS 0.346049f
C552 VN.n17 VSUBS 0.177672f
C553 VN.t8 VSUBS 0.323286f
C554 VN.n18 VSUBS 0.200388f
C555 VN.n19 VSUBS 0.013096f
C556 VN.t1 VSUBS 0.323286f
C557 VN.n20 VSUBS 0.196231f
C558 VN.n21 VSUBS 0.057712f
C559 VN.n22 VSUBS 0.057712f
C560 VN.n23 VSUBS 0.057712f
C561 VN.n24 VSUBS 0.196231f
C562 VN.n25 VSUBS 0.013096f
C563 VN.t0 VSUBS 0.323286f
C564 VN.n26 VSUBS 0.19036f
C565 VN.n27 VSUBS 1.81262f
.ends

