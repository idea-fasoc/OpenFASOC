* NGSPICE file created from diff_pair_sample_0540.ext - technology: sky130A

.subckt diff_pair_sample_0540 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.15 as=0.3003 ps=2.15 w=1.82 l=0.58
X1 VTAIL.t12 VP.t1 VDD1.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.7098 pd=4.42 as=0.3003 ps=2.15 w=1.82 l=0.58
X2 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=0.7098 pd=4.42 as=0 ps=0 w=1.82 l=0.58
X3 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=0.7098 pd=4.42 as=0 ps=0 w=1.82 l=0.58
X4 VDD2.t7 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.15 as=0.3003 ps=2.15 w=1.82 l=0.58
X5 VTAIL.t3 VN.t1 VDD2.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7098 pd=4.42 as=0.3003 ps=2.15 w=1.82 l=0.58
X6 VDD1.t5 VP.t2 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.15 as=0.3003 ps=2.15 w=1.82 l=0.58
X7 VTAIL.t4 VN.t2 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.15 as=0.3003 ps=2.15 w=1.82 l=0.58
X8 VTAIL.t8 VP.t3 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.15 as=0.3003 ps=2.15 w=1.82 l=0.58
X9 VDD2.t4 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.15 as=0.3003 ps=2.15 w=1.82 l=0.58
X10 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=0.7098 pd=4.42 as=0 ps=0 w=1.82 l=0.58
X11 VTAIL.t9 VP.t4 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.15 as=0.3003 ps=2.15 w=1.82 l=0.58
X12 VDD2.t3 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.15 as=0.7098 ps=4.42 w=1.82 l=0.58
X13 VDD1.t2 VP.t5 VTAIL.t15 B.t5 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.15 as=0.7098 ps=4.42 w=1.82 l=0.58
X14 VDD1.t1 VP.t6 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.15 as=0.7098 ps=4.42 w=1.82 l=0.58
X15 VTAIL.t14 VP.t7 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7098 pd=4.42 as=0.3003 ps=2.15 w=1.82 l=0.58
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.7098 pd=4.42 as=0 ps=0 w=1.82 l=0.58
X17 VTAIL.t7 VN.t5 VDD2.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.15 as=0.3003 ps=2.15 w=1.82 l=0.58
X18 VTAIL.t6 VN.t6 VDD2.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=0.7098 pd=4.42 as=0.3003 ps=2.15 w=1.82 l=0.58
X19 VDD2.t0 VN.t7 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.15 as=0.7098 ps=4.42 w=1.82 l=0.58
R0 VP.n4 VP.t1 170.853
R1 VP.n19 VP.n18 161.3
R2 VP.n6 VP.n3 161.3
R3 VP.n7 VP.n2 161.3
R4 VP.n9 VP.n8 161.3
R5 VP.n17 VP.n0 161.3
R6 VP.n16 VP.n15 161.3
R7 VP.n14 VP.n1 161.3
R8 VP.n13 VP.n12 161.3
R9 VP.n11 VP.n10 161.3
R10 VP.n11 VP.t7 144.185
R11 VP.n1 VP.t0 144.185
R12 VP.n16 VP.t3 144.185
R13 VP.n18 VP.t6 144.185
R14 VP.n8 VP.t5 144.185
R15 VP.n6 VP.t4 144.185
R16 VP.n5 VP.t2 144.185
R17 VP.n16 VP.n1 48.2005
R18 VP.n6 VP.n5 48.2005
R19 VP.n12 VP.n11 47.4702
R20 VP.n18 VP.n17 47.4702
R21 VP.n8 VP.n7 47.4702
R22 VP.n4 VP.n3 45.1192
R23 VP.n10 VP.n9 33.7429
R24 VP.n5 VP.n4 13.6377
R25 VP.n12 VP.n1 0.730803
R26 VP.n17 VP.n16 0.730803
R27 VP.n7 VP.n6 0.730803
R28 VP.n3 VP.n2 0.189894
R29 VP.n9 VP.n2 0.189894
R30 VP.n13 VP.n10 0.189894
R31 VP.n14 VP.n13 0.189894
R32 VP.n15 VP.n14 0.189894
R33 VP.n15 VP.n0 0.189894
R34 VP.n19 VP.n0 0.189894
R35 VP VP.n19 0.0516364
R36 VTAIL.n66 VTAIL.n64 289.615
R37 VTAIL.n4 VTAIL.n2 289.615
R38 VTAIL.n12 VTAIL.n10 289.615
R39 VTAIL.n22 VTAIL.n20 289.615
R40 VTAIL.n58 VTAIL.n56 289.615
R41 VTAIL.n48 VTAIL.n46 289.615
R42 VTAIL.n40 VTAIL.n38 289.615
R43 VTAIL.n30 VTAIL.n28 289.615
R44 VTAIL.n67 VTAIL.n66 185
R45 VTAIL.n5 VTAIL.n4 185
R46 VTAIL.n13 VTAIL.n12 185
R47 VTAIL.n23 VTAIL.n22 185
R48 VTAIL.n59 VTAIL.n58 185
R49 VTAIL.n49 VTAIL.n48 185
R50 VTAIL.n41 VTAIL.n40 185
R51 VTAIL.n31 VTAIL.n30 185
R52 VTAIL.t5 VTAIL.n65 164.876
R53 VTAIL.t6 VTAIL.n3 164.876
R54 VTAIL.t13 VTAIL.n11 164.876
R55 VTAIL.t14 VTAIL.n21 164.876
R56 VTAIL.t15 VTAIL.n57 164.876
R57 VTAIL.t12 VTAIL.n47 164.876
R58 VTAIL.t0 VTAIL.n39 164.876
R59 VTAIL.t3 VTAIL.n29 164.876
R60 VTAIL.n55 VTAIL.n54 85.5201
R61 VTAIL.n37 VTAIL.n36 85.5201
R62 VTAIL.n1 VTAIL.n0 85.52
R63 VTAIL.n19 VTAIL.n18 85.52
R64 VTAIL.n66 VTAIL.t5 52.3082
R65 VTAIL.n4 VTAIL.t6 52.3082
R66 VTAIL.n12 VTAIL.t13 52.3082
R67 VTAIL.n22 VTAIL.t14 52.3082
R68 VTAIL.n58 VTAIL.t15 52.3082
R69 VTAIL.n48 VTAIL.t12 52.3082
R70 VTAIL.n40 VTAIL.t0 52.3082
R71 VTAIL.n30 VTAIL.t3 52.3082
R72 VTAIL.n71 VTAIL.n70 34.9005
R73 VTAIL.n9 VTAIL.n8 34.9005
R74 VTAIL.n17 VTAIL.n16 34.9005
R75 VTAIL.n27 VTAIL.n26 34.9005
R76 VTAIL.n63 VTAIL.n62 34.9005
R77 VTAIL.n53 VTAIL.n52 34.9005
R78 VTAIL.n45 VTAIL.n44 34.9005
R79 VTAIL.n35 VTAIL.n34 34.9005
R80 VTAIL.n67 VTAIL.n65 14.7318
R81 VTAIL.n5 VTAIL.n3 14.7318
R82 VTAIL.n13 VTAIL.n11 14.7318
R83 VTAIL.n23 VTAIL.n21 14.7318
R84 VTAIL.n59 VTAIL.n57 14.7318
R85 VTAIL.n49 VTAIL.n47 14.7318
R86 VTAIL.n41 VTAIL.n39 14.7318
R87 VTAIL.n31 VTAIL.n29 14.7318
R88 VTAIL.n71 VTAIL.n63 14.7203
R89 VTAIL.n35 VTAIL.n27 14.7203
R90 VTAIL.n68 VTAIL.n64 12.8005
R91 VTAIL.n6 VTAIL.n2 12.8005
R92 VTAIL.n14 VTAIL.n10 12.8005
R93 VTAIL.n24 VTAIL.n20 12.8005
R94 VTAIL.n60 VTAIL.n56 12.8005
R95 VTAIL.n50 VTAIL.n46 12.8005
R96 VTAIL.n42 VTAIL.n38 12.8005
R97 VTAIL.n32 VTAIL.n28 12.8005
R98 VTAIL.n0 VTAIL.t1 10.8796
R99 VTAIL.n0 VTAIL.t4 10.8796
R100 VTAIL.n18 VTAIL.t11 10.8796
R101 VTAIL.n18 VTAIL.t8 10.8796
R102 VTAIL.n54 VTAIL.t10 10.8796
R103 VTAIL.n54 VTAIL.t9 10.8796
R104 VTAIL.n36 VTAIL.t2 10.8796
R105 VTAIL.n36 VTAIL.t7 10.8796
R106 VTAIL.n70 VTAIL.n69 9.45567
R107 VTAIL.n8 VTAIL.n7 9.45567
R108 VTAIL.n16 VTAIL.n15 9.45567
R109 VTAIL.n26 VTAIL.n25 9.45567
R110 VTAIL.n62 VTAIL.n61 9.45567
R111 VTAIL.n52 VTAIL.n51 9.45567
R112 VTAIL.n44 VTAIL.n43 9.45567
R113 VTAIL.n34 VTAIL.n33 9.45567
R114 VTAIL.n69 VTAIL.n68 9.3005
R115 VTAIL.n7 VTAIL.n6 9.3005
R116 VTAIL.n15 VTAIL.n14 9.3005
R117 VTAIL.n25 VTAIL.n24 9.3005
R118 VTAIL.n61 VTAIL.n60 9.3005
R119 VTAIL.n51 VTAIL.n50 9.3005
R120 VTAIL.n43 VTAIL.n42 9.3005
R121 VTAIL.n33 VTAIL.n32 9.3005
R122 VTAIL.n69 VTAIL.n65 5.62509
R123 VTAIL.n7 VTAIL.n3 5.62509
R124 VTAIL.n15 VTAIL.n11 5.62509
R125 VTAIL.n25 VTAIL.n21 5.62509
R126 VTAIL.n61 VTAIL.n57 5.62509
R127 VTAIL.n51 VTAIL.n47 5.62509
R128 VTAIL.n43 VTAIL.n39 5.62509
R129 VTAIL.n33 VTAIL.n29 5.62509
R130 VTAIL.n70 VTAIL.n64 1.16414
R131 VTAIL.n8 VTAIL.n2 1.16414
R132 VTAIL.n16 VTAIL.n10 1.16414
R133 VTAIL.n26 VTAIL.n20 1.16414
R134 VTAIL.n62 VTAIL.n56 1.16414
R135 VTAIL.n52 VTAIL.n46 1.16414
R136 VTAIL.n44 VTAIL.n38 1.16414
R137 VTAIL.n34 VTAIL.n28 1.16414
R138 VTAIL.n37 VTAIL.n35 0.784983
R139 VTAIL.n45 VTAIL.n37 0.784983
R140 VTAIL.n55 VTAIL.n53 0.784983
R141 VTAIL.n63 VTAIL.n55 0.784983
R142 VTAIL.n27 VTAIL.n19 0.784983
R143 VTAIL.n19 VTAIL.n17 0.784983
R144 VTAIL.n9 VTAIL.n1 0.784983
R145 VTAIL VTAIL.n71 0.726793
R146 VTAIL.n53 VTAIL.n45 0.470328
R147 VTAIL.n17 VTAIL.n9 0.470328
R148 VTAIL.n68 VTAIL.n67 0.388379
R149 VTAIL.n6 VTAIL.n5 0.388379
R150 VTAIL.n14 VTAIL.n13 0.388379
R151 VTAIL.n24 VTAIL.n23 0.388379
R152 VTAIL.n60 VTAIL.n59 0.388379
R153 VTAIL.n50 VTAIL.n49 0.388379
R154 VTAIL.n42 VTAIL.n41 0.388379
R155 VTAIL.n32 VTAIL.n31 0.388379
R156 VTAIL VTAIL.n1 0.0586897
R157 VDD1 VDD1.n0 102.65
R158 VDD1.n3 VDD1.n2 102.535
R159 VDD1.n3 VDD1.n1 102.535
R160 VDD1.n5 VDD1.n4 102.198
R161 VDD1.n5 VDD1.n3 29.3974
R162 VDD1.n4 VDD1.t3 10.8796
R163 VDD1.n4 VDD1.t2 10.8796
R164 VDD1.n0 VDD1.t6 10.8796
R165 VDD1.n0 VDD1.t5 10.8796
R166 VDD1.n2 VDD1.t4 10.8796
R167 VDD1.n2 VDD1.t1 10.8796
R168 VDD1.n1 VDD1.t0 10.8796
R169 VDD1.n1 VDD1.t7 10.8796
R170 VDD1 VDD1.n5 0.334552
R171 B.n350 B.n349 585
R172 B.n351 B.n350 585
R173 B.n128 B.n59 585
R174 B.n127 B.n126 585
R175 B.n125 B.n124 585
R176 B.n123 B.n122 585
R177 B.n121 B.n120 585
R178 B.n119 B.n118 585
R179 B.n117 B.n116 585
R180 B.n115 B.n114 585
R181 B.n113 B.n112 585
R182 B.n111 B.n110 585
R183 B.n109 B.n108 585
R184 B.n106 B.n105 585
R185 B.n104 B.n103 585
R186 B.n102 B.n101 585
R187 B.n100 B.n99 585
R188 B.n98 B.n97 585
R189 B.n96 B.n95 585
R190 B.n94 B.n93 585
R191 B.n92 B.n91 585
R192 B.n90 B.n89 585
R193 B.n88 B.n87 585
R194 B.n86 B.n85 585
R195 B.n84 B.n83 585
R196 B.n82 B.n81 585
R197 B.n80 B.n79 585
R198 B.n78 B.n77 585
R199 B.n76 B.n75 585
R200 B.n74 B.n73 585
R201 B.n72 B.n71 585
R202 B.n70 B.n69 585
R203 B.n68 B.n67 585
R204 B.n66 B.n65 585
R205 B.n348 B.n42 585
R206 B.n352 B.n42 585
R207 B.n347 B.n41 585
R208 B.n353 B.n41 585
R209 B.n346 B.n345 585
R210 B.n345 B.n37 585
R211 B.n344 B.n36 585
R212 B.n359 B.n36 585
R213 B.n343 B.n35 585
R214 B.n360 B.n35 585
R215 B.n342 B.n34 585
R216 B.n361 B.n34 585
R217 B.n341 B.n340 585
R218 B.n340 B.n30 585
R219 B.n339 B.n29 585
R220 B.n367 B.n29 585
R221 B.n338 B.n28 585
R222 B.n368 B.n28 585
R223 B.n337 B.n27 585
R224 B.n369 B.n27 585
R225 B.n336 B.n335 585
R226 B.n335 B.n26 585
R227 B.n334 B.n22 585
R228 B.n375 B.n22 585
R229 B.n333 B.n21 585
R230 B.n376 B.n21 585
R231 B.n332 B.n20 585
R232 B.n377 B.n20 585
R233 B.n331 B.n330 585
R234 B.n330 B.n16 585
R235 B.n329 B.n15 585
R236 B.n383 B.n15 585
R237 B.n328 B.n14 585
R238 B.n384 B.n14 585
R239 B.n327 B.n13 585
R240 B.n385 B.n13 585
R241 B.n326 B.n325 585
R242 B.n325 B.n12 585
R243 B.n324 B.n323 585
R244 B.n324 B.n8 585
R245 B.n322 B.n7 585
R246 B.n392 B.n7 585
R247 B.n321 B.n6 585
R248 B.n393 B.n6 585
R249 B.n320 B.n5 585
R250 B.n394 B.n5 585
R251 B.n319 B.n318 585
R252 B.n318 B.n4 585
R253 B.n317 B.n129 585
R254 B.n317 B.n316 585
R255 B.n306 B.n130 585
R256 B.n309 B.n130 585
R257 B.n308 B.n307 585
R258 B.n310 B.n308 585
R259 B.n305 B.n135 585
R260 B.n135 B.n134 585
R261 B.n304 B.n303 585
R262 B.n303 B.n302 585
R263 B.n137 B.n136 585
R264 B.n138 B.n137 585
R265 B.n295 B.n294 585
R266 B.n296 B.n295 585
R267 B.n293 B.n143 585
R268 B.n143 B.n142 585
R269 B.n292 B.n291 585
R270 B.n291 B.n290 585
R271 B.n145 B.n144 585
R272 B.n283 B.n145 585
R273 B.n282 B.n281 585
R274 B.n284 B.n282 585
R275 B.n280 B.n150 585
R276 B.n150 B.n149 585
R277 B.n279 B.n278 585
R278 B.n278 B.n277 585
R279 B.n152 B.n151 585
R280 B.n153 B.n152 585
R281 B.n270 B.n269 585
R282 B.n271 B.n270 585
R283 B.n268 B.n157 585
R284 B.n161 B.n157 585
R285 B.n267 B.n266 585
R286 B.n266 B.n265 585
R287 B.n159 B.n158 585
R288 B.n160 B.n159 585
R289 B.n258 B.n257 585
R290 B.n259 B.n258 585
R291 B.n256 B.n166 585
R292 B.n166 B.n165 585
R293 B.n250 B.n249 585
R294 B.n248 B.n184 585
R295 B.n247 B.n183 585
R296 B.n252 B.n183 585
R297 B.n246 B.n245 585
R298 B.n244 B.n243 585
R299 B.n242 B.n241 585
R300 B.n240 B.n239 585
R301 B.n238 B.n237 585
R302 B.n236 B.n235 585
R303 B.n234 B.n233 585
R304 B.n232 B.n231 585
R305 B.n230 B.n229 585
R306 B.n227 B.n226 585
R307 B.n225 B.n224 585
R308 B.n223 B.n222 585
R309 B.n221 B.n220 585
R310 B.n219 B.n218 585
R311 B.n217 B.n216 585
R312 B.n215 B.n214 585
R313 B.n213 B.n212 585
R314 B.n211 B.n210 585
R315 B.n209 B.n208 585
R316 B.n207 B.n206 585
R317 B.n205 B.n204 585
R318 B.n203 B.n202 585
R319 B.n201 B.n200 585
R320 B.n199 B.n198 585
R321 B.n197 B.n196 585
R322 B.n195 B.n194 585
R323 B.n193 B.n192 585
R324 B.n191 B.n190 585
R325 B.n168 B.n167 585
R326 B.n255 B.n254 585
R327 B.n164 B.n163 585
R328 B.n165 B.n164 585
R329 B.n261 B.n260 585
R330 B.n260 B.n259 585
R331 B.n262 B.n162 585
R332 B.n162 B.n160 585
R333 B.n264 B.n263 585
R334 B.n265 B.n264 585
R335 B.n156 B.n155 585
R336 B.n161 B.n156 585
R337 B.n273 B.n272 585
R338 B.n272 B.n271 585
R339 B.n274 B.n154 585
R340 B.n154 B.n153 585
R341 B.n276 B.n275 585
R342 B.n277 B.n276 585
R343 B.n148 B.n147 585
R344 B.n149 B.n148 585
R345 B.n286 B.n285 585
R346 B.n285 B.n284 585
R347 B.n287 B.n146 585
R348 B.n283 B.n146 585
R349 B.n289 B.n288 585
R350 B.n290 B.n289 585
R351 B.n141 B.n140 585
R352 B.n142 B.n141 585
R353 B.n298 B.n297 585
R354 B.n297 B.n296 585
R355 B.n299 B.n139 585
R356 B.n139 B.n138 585
R357 B.n301 B.n300 585
R358 B.n302 B.n301 585
R359 B.n133 B.n132 585
R360 B.n134 B.n133 585
R361 B.n312 B.n311 585
R362 B.n311 B.n310 585
R363 B.n313 B.n131 585
R364 B.n309 B.n131 585
R365 B.n315 B.n314 585
R366 B.n316 B.n315 585
R367 B.n3 B.n0 585
R368 B.n4 B.n3 585
R369 B.n391 B.n1 585
R370 B.n392 B.n391 585
R371 B.n390 B.n389 585
R372 B.n390 B.n8 585
R373 B.n388 B.n9 585
R374 B.n12 B.n9 585
R375 B.n387 B.n386 585
R376 B.n386 B.n385 585
R377 B.n11 B.n10 585
R378 B.n384 B.n11 585
R379 B.n382 B.n381 585
R380 B.n383 B.n382 585
R381 B.n380 B.n17 585
R382 B.n17 B.n16 585
R383 B.n379 B.n378 585
R384 B.n378 B.n377 585
R385 B.n19 B.n18 585
R386 B.n376 B.n19 585
R387 B.n374 B.n373 585
R388 B.n375 B.n374 585
R389 B.n372 B.n23 585
R390 B.n26 B.n23 585
R391 B.n371 B.n370 585
R392 B.n370 B.n369 585
R393 B.n25 B.n24 585
R394 B.n368 B.n25 585
R395 B.n366 B.n365 585
R396 B.n367 B.n366 585
R397 B.n364 B.n31 585
R398 B.n31 B.n30 585
R399 B.n363 B.n362 585
R400 B.n362 B.n361 585
R401 B.n33 B.n32 585
R402 B.n360 B.n33 585
R403 B.n358 B.n357 585
R404 B.n359 B.n358 585
R405 B.n356 B.n38 585
R406 B.n38 B.n37 585
R407 B.n355 B.n354 585
R408 B.n354 B.n353 585
R409 B.n40 B.n39 585
R410 B.n352 B.n40 585
R411 B.n395 B.n394 585
R412 B.n393 B.n2 585
R413 B.n65 B.n40 492.5
R414 B.n350 B.n42 492.5
R415 B.n254 B.n166 492.5
R416 B.n250 B.n164 492.5
R417 B.n60 B.t19 281.101
R418 B.n187 B.t8 281.101
R419 B.n62 B.t12 280.786
R420 B.n185 B.t16 280.786
R421 B.n351 B.n58 256.663
R422 B.n351 B.n57 256.663
R423 B.n351 B.n56 256.663
R424 B.n351 B.n55 256.663
R425 B.n351 B.n54 256.663
R426 B.n351 B.n53 256.663
R427 B.n351 B.n52 256.663
R428 B.n351 B.n51 256.663
R429 B.n351 B.n50 256.663
R430 B.n351 B.n49 256.663
R431 B.n351 B.n48 256.663
R432 B.n351 B.n47 256.663
R433 B.n351 B.n46 256.663
R434 B.n351 B.n45 256.663
R435 B.n351 B.n44 256.663
R436 B.n351 B.n43 256.663
R437 B.n252 B.n251 256.663
R438 B.n252 B.n169 256.663
R439 B.n252 B.n170 256.663
R440 B.n252 B.n171 256.663
R441 B.n252 B.n172 256.663
R442 B.n252 B.n173 256.663
R443 B.n252 B.n174 256.663
R444 B.n252 B.n175 256.663
R445 B.n252 B.n176 256.663
R446 B.n252 B.n177 256.663
R447 B.n252 B.n178 256.663
R448 B.n252 B.n179 256.663
R449 B.n252 B.n180 256.663
R450 B.n252 B.n181 256.663
R451 B.n252 B.n182 256.663
R452 B.n253 B.n252 256.663
R453 B.n397 B.n396 256.663
R454 B.n252 B.n165 190.698
R455 B.n352 B.n351 190.698
R456 B.n69 B.n68 163.367
R457 B.n73 B.n72 163.367
R458 B.n77 B.n76 163.367
R459 B.n81 B.n80 163.367
R460 B.n85 B.n84 163.367
R461 B.n89 B.n88 163.367
R462 B.n93 B.n92 163.367
R463 B.n97 B.n96 163.367
R464 B.n101 B.n100 163.367
R465 B.n105 B.n104 163.367
R466 B.n110 B.n109 163.367
R467 B.n114 B.n113 163.367
R468 B.n118 B.n117 163.367
R469 B.n122 B.n121 163.367
R470 B.n126 B.n125 163.367
R471 B.n350 B.n59 163.367
R472 B.n258 B.n166 163.367
R473 B.n258 B.n159 163.367
R474 B.n266 B.n159 163.367
R475 B.n266 B.n157 163.367
R476 B.n270 B.n157 163.367
R477 B.n270 B.n152 163.367
R478 B.n278 B.n152 163.367
R479 B.n278 B.n150 163.367
R480 B.n282 B.n150 163.367
R481 B.n282 B.n145 163.367
R482 B.n291 B.n145 163.367
R483 B.n291 B.n143 163.367
R484 B.n295 B.n143 163.367
R485 B.n295 B.n137 163.367
R486 B.n303 B.n137 163.367
R487 B.n303 B.n135 163.367
R488 B.n308 B.n135 163.367
R489 B.n308 B.n130 163.367
R490 B.n317 B.n130 163.367
R491 B.n318 B.n317 163.367
R492 B.n318 B.n5 163.367
R493 B.n6 B.n5 163.367
R494 B.n7 B.n6 163.367
R495 B.n324 B.n7 163.367
R496 B.n325 B.n324 163.367
R497 B.n325 B.n13 163.367
R498 B.n14 B.n13 163.367
R499 B.n15 B.n14 163.367
R500 B.n330 B.n15 163.367
R501 B.n330 B.n20 163.367
R502 B.n21 B.n20 163.367
R503 B.n22 B.n21 163.367
R504 B.n335 B.n22 163.367
R505 B.n335 B.n27 163.367
R506 B.n28 B.n27 163.367
R507 B.n29 B.n28 163.367
R508 B.n340 B.n29 163.367
R509 B.n340 B.n34 163.367
R510 B.n35 B.n34 163.367
R511 B.n36 B.n35 163.367
R512 B.n345 B.n36 163.367
R513 B.n345 B.n41 163.367
R514 B.n42 B.n41 163.367
R515 B.n184 B.n183 163.367
R516 B.n245 B.n183 163.367
R517 B.n243 B.n242 163.367
R518 B.n239 B.n238 163.367
R519 B.n235 B.n234 163.367
R520 B.n231 B.n230 163.367
R521 B.n226 B.n225 163.367
R522 B.n222 B.n221 163.367
R523 B.n218 B.n217 163.367
R524 B.n214 B.n213 163.367
R525 B.n210 B.n209 163.367
R526 B.n206 B.n205 163.367
R527 B.n202 B.n201 163.367
R528 B.n198 B.n197 163.367
R529 B.n194 B.n193 163.367
R530 B.n190 B.n168 163.367
R531 B.n260 B.n164 163.367
R532 B.n260 B.n162 163.367
R533 B.n264 B.n162 163.367
R534 B.n264 B.n156 163.367
R535 B.n272 B.n156 163.367
R536 B.n272 B.n154 163.367
R537 B.n276 B.n154 163.367
R538 B.n276 B.n148 163.367
R539 B.n285 B.n148 163.367
R540 B.n285 B.n146 163.367
R541 B.n289 B.n146 163.367
R542 B.n289 B.n141 163.367
R543 B.n297 B.n141 163.367
R544 B.n297 B.n139 163.367
R545 B.n301 B.n139 163.367
R546 B.n301 B.n133 163.367
R547 B.n311 B.n133 163.367
R548 B.n311 B.n131 163.367
R549 B.n315 B.n131 163.367
R550 B.n315 B.n3 163.367
R551 B.n395 B.n3 163.367
R552 B.n391 B.n2 163.367
R553 B.n391 B.n390 163.367
R554 B.n390 B.n9 163.367
R555 B.n386 B.n9 163.367
R556 B.n386 B.n11 163.367
R557 B.n382 B.n11 163.367
R558 B.n382 B.n17 163.367
R559 B.n378 B.n17 163.367
R560 B.n378 B.n19 163.367
R561 B.n374 B.n19 163.367
R562 B.n374 B.n23 163.367
R563 B.n370 B.n23 163.367
R564 B.n370 B.n25 163.367
R565 B.n366 B.n25 163.367
R566 B.n366 B.n31 163.367
R567 B.n362 B.n31 163.367
R568 B.n362 B.n33 163.367
R569 B.n358 B.n33 163.367
R570 B.n358 B.n38 163.367
R571 B.n354 B.n38 163.367
R572 B.n354 B.n40 163.367
R573 B.n60 B.t20 137.369
R574 B.n187 B.t11 137.369
R575 B.n62 B.t14 137.369
R576 B.n185 B.t18 137.369
R577 B.n61 B.t21 119.722
R578 B.n188 B.t10 119.722
R579 B.n63 B.t15 119.722
R580 B.n186 B.t17 119.722
R581 B.n259 B.n165 105.427
R582 B.n259 B.n160 105.427
R583 B.n265 B.n160 105.427
R584 B.n265 B.n161 105.427
R585 B.n271 B.n153 105.427
R586 B.n277 B.n153 105.427
R587 B.n277 B.n149 105.427
R588 B.n284 B.n149 105.427
R589 B.n284 B.n283 105.427
R590 B.n290 B.n142 105.427
R591 B.n296 B.n142 105.427
R592 B.n302 B.n138 105.427
R593 B.n310 B.n134 105.427
R594 B.n310 B.n309 105.427
R595 B.n316 B.n4 105.427
R596 B.n394 B.n4 105.427
R597 B.n394 B.n393 105.427
R598 B.n393 B.n392 105.427
R599 B.n392 B.n8 105.427
R600 B.n385 B.n12 105.427
R601 B.n385 B.n384 105.427
R602 B.n383 B.n16 105.427
R603 B.n377 B.n376 105.427
R604 B.n376 B.n375 105.427
R605 B.n369 B.n26 105.427
R606 B.n369 B.n368 105.427
R607 B.n368 B.n367 105.427
R608 B.n367 B.n30 105.427
R609 B.n361 B.n30 105.427
R610 B.n360 B.n359 105.427
R611 B.n359 B.n37 105.427
R612 B.n353 B.n37 105.427
R613 B.n353 B.n352 105.427
R614 B.n302 B.t7 93.0238
R615 B.t1 B.n383 93.0238
R616 B.t2 B.n138 83.7214
R617 B.t4 B.n16 83.7214
R618 B.n65 B.n43 71.676
R619 B.n69 B.n44 71.676
R620 B.n73 B.n45 71.676
R621 B.n77 B.n46 71.676
R622 B.n81 B.n47 71.676
R623 B.n85 B.n48 71.676
R624 B.n89 B.n49 71.676
R625 B.n93 B.n50 71.676
R626 B.n97 B.n51 71.676
R627 B.n101 B.n52 71.676
R628 B.n105 B.n53 71.676
R629 B.n110 B.n54 71.676
R630 B.n114 B.n55 71.676
R631 B.n118 B.n56 71.676
R632 B.n122 B.n57 71.676
R633 B.n126 B.n58 71.676
R634 B.n59 B.n58 71.676
R635 B.n125 B.n57 71.676
R636 B.n121 B.n56 71.676
R637 B.n117 B.n55 71.676
R638 B.n113 B.n54 71.676
R639 B.n109 B.n53 71.676
R640 B.n104 B.n52 71.676
R641 B.n100 B.n51 71.676
R642 B.n96 B.n50 71.676
R643 B.n92 B.n49 71.676
R644 B.n88 B.n48 71.676
R645 B.n84 B.n47 71.676
R646 B.n80 B.n46 71.676
R647 B.n76 B.n45 71.676
R648 B.n72 B.n44 71.676
R649 B.n68 B.n43 71.676
R650 B.n251 B.n250 71.676
R651 B.n245 B.n169 71.676
R652 B.n242 B.n170 71.676
R653 B.n238 B.n171 71.676
R654 B.n234 B.n172 71.676
R655 B.n230 B.n173 71.676
R656 B.n225 B.n174 71.676
R657 B.n221 B.n175 71.676
R658 B.n217 B.n176 71.676
R659 B.n213 B.n177 71.676
R660 B.n209 B.n178 71.676
R661 B.n205 B.n179 71.676
R662 B.n201 B.n180 71.676
R663 B.n197 B.n181 71.676
R664 B.n193 B.n182 71.676
R665 B.n253 B.n168 71.676
R666 B.n251 B.n184 71.676
R667 B.n243 B.n169 71.676
R668 B.n239 B.n170 71.676
R669 B.n235 B.n171 71.676
R670 B.n231 B.n172 71.676
R671 B.n226 B.n173 71.676
R672 B.n222 B.n174 71.676
R673 B.n218 B.n175 71.676
R674 B.n214 B.n176 71.676
R675 B.n210 B.n177 71.676
R676 B.n206 B.n178 71.676
R677 B.n202 B.n179 71.676
R678 B.n198 B.n180 71.676
R679 B.n194 B.n181 71.676
R680 B.n190 B.n182 71.676
R681 B.n254 B.n253 71.676
R682 B.n396 B.n395 71.676
R683 B.n396 B.n2 71.676
R684 B.n161 B.t9 68.2176
R685 B.t13 B.n360 68.2176
R686 B.n64 B.n63 59.5399
R687 B.n107 B.n61 59.5399
R688 B.n189 B.n188 59.5399
R689 B.n228 B.n186 59.5399
R690 B.n309 B.t0 58.9152
R691 B.n12 B.t6 58.9152
R692 B.n283 B.t3 55.8145
R693 B.n26 B.t5 55.8145
R694 B.n290 B.t3 49.6129
R695 B.n375 B.t5 49.6129
R696 B.n316 B.t0 46.5121
R697 B.t6 B.n8 46.5121
R698 B.n271 B.t9 37.2098
R699 B.n361 B.t13 37.2098
R700 B.n249 B.n163 32.0005
R701 B.n256 B.n255 32.0005
R702 B.n349 B.n348 32.0005
R703 B.n66 B.n39 32.0005
R704 B.n296 B.t2 21.7059
R705 B.n377 B.t4 21.7059
R706 B B.n397 18.0485
R707 B.n63 B.n62 17.649
R708 B.n61 B.n60 17.649
R709 B.n188 B.n187 17.649
R710 B.n186 B.n185 17.649
R711 B.t7 B.n134 12.4036
R712 B.n384 B.t1 12.4036
R713 B.n261 B.n163 10.6151
R714 B.n262 B.n261 10.6151
R715 B.n263 B.n262 10.6151
R716 B.n263 B.n155 10.6151
R717 B.n273 B.n155 10.6151
R718 B.n274 B.n273 10.6151
R719 B.n275 B.n274 10.6151
R720 B.n275 B.n147 10.6151
R721 B.n286 B.n147 10.6151
R722 B.n287 B.n286 10.6151
R723 B.n288 B.n287 10.6151
R724 B.n288 B.n140 10.6151
R725 B.n298 B.n140 10.6151
R726 B.n299 B.n298 10.6151
R727 B.n300 B.n299 10.6151
R728 B.n300 B.n132 10.6151
R729 B.n312 B.n132 10.6151
R730 B.n313 B.n312 10.6151
R731 B.n314 B.n313 10.6151
R732 B.n314 B.n0 10.6151
R733 B.n249 B.n248 10.6151
R734 B.n248 B.n247 10.6151
R735 B.n247 B.n246 10.6151
R736 B.n246 B.n244 10.6151
R737 B.n244 B.n241 10.6151
R738 B.n241 B.n240 10.6151
R739 B.n240 B.n237 10.6151
R740 B.n237 B.n236 10.6151
R741 B.n236 B.n233 10.6151
R742 B.n233 B.n232 10.6151
R743 B.n232 B.n229 10.6151
R744 B.n227 B.n224 10.6151
R745 B.n224 B.n223 10.6151
R746 B.n223 B.n220 10.6151
R747 B.n220 B.n219 10.6151
R748 B.n219 B.n216 10.6151
R749 B.n216 B.n215 10.6151
R750 B.n215 B.n212 10.6151
R751 B.n212 B.n211 10.6151
R752 B.n208 B.n207 10.6151
R753 B.n207 B.n204 10.6151
R754 B.n204 B.n203 10.6151
R755 B.n203 B.n200 10.6151
R756 B.n200 B.n199 10.6151
R757 B.n199 B.n196 10.6151
R758 B.n196 B.n195 10.6151
R759 B.n195 B.n192 10.6151
R760 B.n192 B.n191 10.6151
R761 B.n191 B.n167 10.6151
R762 B.n255 B.n167 10.6151
R763 B.n257 B.n256 10.6151
R764 B.n257 B.n158 10.6151
R765 B.n267 B.n158 10.6151
R766 B.n268 B.n267 10.6151
R767 B.n269 B.n268 10.6151
R768 B.n269 B.n151 10.6151
R769 B.n279 B.n151 10.6151
R770 B.n280 B.n279 10.6151
R771 B.n281 B.n280 10.6151
R772 B.n281 B.n144 10.6151
R773 B.n292 B.n144 10.6151
R774 B.n293 B.n292 10.6151
R775 B.n294 B.n293 10.6151
R776 B.n294 B.n136 10.6151
R777 B.n304 B.n136 10.6151
R778 B.n305 B.n304 10.6151
R779 B.n307 B.n305 10.6151
R780 B.n307 B.n306 10.6151
R781 B.n306 B.n129 10.6151
R782 B.n319 B.n129 10.6151
R783 B.n320 B.n319 10.6151
R784 B.n321 B.n320 10.6151
R785 B.n322 B.n321 10.6151
R786 B.n323 B.n322 10.6151
R787 B.n326 B.n323 10.6151
R788 B.n327 B.n326 10.6151
R789 B.n328 B.n327 10.6151
R790 B.n329 B.n328 10.6151
R791 B.n331 B.n329 10.6151
R792 B.n332 B.n331 10.6151
R793 B.n333 B.n332 10.6151
R794 B.n334 B.n333 10.6151
R795 B.n336 B.n334 10.6151
R796 B.n337 B.n336 10.6151
R797 B.n338 B.n337 10.6151
R798 B.n339 B.n338 10.6151
R799 B.n341 B.n339 10.6151
R800 B.n342 B.n341 10.6151
R801 B.n343 B.n342 10.6151
R802 B.n344 B.n343 10.6151
R803 B.n346 B.n344 10.6151
R804 B.n347 B.n346 10.6151
R805 B.n348 B.n347 10.6151
R806 B.n389 B.n1 10.6151
R807 B.n389 B.n388 10.6151
R808 B.n388 B.n387 10.6151
R809 B.n387 B.n10 10.6151
R810 B.n381 B.n10 10.6151
R811 B.n381 B.n380 10.6151
R812 B.n380 B.n379 10.6151
R813 B.n379 B.n18 10.6151
R814 B.n373 B.n18 10.6151
R815 B.n373 B.n372 10.6151
R816 B.n372 B.n371 10.6151
R817 B.n371 B.n24 10.6151
R818 B.n365 B.n24 10.6151
R819 B.n365 B.n364 10.6151
R820 B.n364 B.n363 10.6151
R821 B.n363 B.n32 10.6151
R822 B.n357 B.n32 10.6151
R823 B.n357 B.n356 10.6151
R824 B.n356 B.n355 10.6151
R825 B.n355 B.n39 10.6151
R826 B.n67 B.n66 10.6151
R827 B.n70 B.n67 10.6151
R828 B.n71 B.n70 10.6151
R829 B.n74 B.n71 10.6151
R830 B.n75 B.n74 10.6151
R831 B.n78 B.n75 10.6151
R832 B.n79 B.n78 10.6151
R833 B.n82 B.n79 10.6151
R834 B.n83 B.n82 10.6151
R835 B.n86 B.n83 10.6151
R836 B.n87 B.n86 10.6151
R837 B.n91 B.n90 10.6151
R838 B.n94 B.n91 10.6151
R839 B.n95 B.n94 10.6151
R840 B.n98 B.n95 10.6151
R841 B.n99 B.n98 10.6151
R842 B.n102 B.n99 10.6151
R843 B.n103 B.n102 10.6151
R844 B.n106 B.n103 10.6151
R845 B.n111 B.n108 10.6151
R846 B.n112 B.n111 10.6151
R847 B.n115 B.n112 10.6151
R848 B.n116 B.n115 10.6151
R849 B.n119 B.n116 10.6151
R850 B.n120 B.n119 10.6151
R851 B.n123 B.n120 10.6151
R852 B.n124 B.n123 10.6151
R853 B.n127 B.n124 10.6151
R854 B.n128 B.n127 10.6151
R855 B.n349 B.n128 10.6151
R856 B.n397 B.n0 8.11757
R857 B.n397 B.n1 8.11757
R858 B.n228 B.n227 6.4005
R859 B.n211 B.n189 6.4005
R860 B.n90 B.n64 6.4005
R861 B.n107 B.n106 6.4005
R862 B.n229 B.n228 4.21513
R863 B.n208 B.n189 4.21513
R864 B.n87 B.n64 4.21513
R865 B.n108 B.n107 4.21513
R866 VN.n2 VN.t6 170.853
R867 VN.n10 VN.t4 170.853
R868 VN.n7 VN.n6 161.3
R869 VN.n15 VN.n14 161.3
R870 VN.n13 VN.n8 161.3
R871 VN.n12 VN.n11 161.3
R872 VN.n5 VN.n0 161.3
R873 VN.n4 VN.n3 161.3
R874 VN.n1 VN.t3 144.185
R875 VN.n4 VN.t2 144.185
R876 VN.n6 VN.t7 144.185
R877 VN.n9 VN.t5 144.185
R878 VN.n12 VN.t0 144.185
R879 VN.n14 VN.t1 144.185
R880 VN.n4 VN.n1 48.2005
R881 VN.n12 VN.n9 48.2005
R882 VN.n6 VN.n5 47.4702
R883 VN.n14 VN.n13 47.4702
R884 VN.n11 VN.n10 45.1192
R885 VN.n3 VN.n2 45.1192
R886 VN VN.n15 34.1236
R887 VN.n2 VN.n1 13.6377
R888 VN.n10 VN.n9 13.6377
R889 VN.n5 VN.n4 0.730803
R890 VN.n13 VN.n12 0.730803
R891 VN.n15 VN.n8 0.189894
R892 VN.n11 VN.n8 0.189894
R893 VN.n3 VN.n0 0.189894
R894 VN.n7 VN.n0 0.189894
R895 VN VN.n7 0.0516364
R896 VDD2.n2 VDD2.n1 102.535
R897 VDD2.n2 VDD2.n0 102.535
R898 VDD2 VDD2.n5 102.532
R899 VDD2.n4 VDD2.n3 102.198
R900 VDD2.n4 VDD2.n2 28.8144
R901 VDD2.n5 VDD2.t2 10.8796
R902 VDD2.n5 VDD2.t3 10.8796
R903 VDD2.n3 VDD2.t6 10.8796
R904 VDD2.n3 VDD2.t7 10.8796
R905 VDD2.n1 VDD2.t5 10.8796
R906 VDD2.n1 VDD2.t0 10.8796
R907 VDD2.n0 VDD2.t1 10.8796
R908 VDD2.n0 VDD2.t4 10.8796
R909 VDD2 VDD2.n4 0.450931
C0 VDD1 VP 1.2298f
C1 VDD2 VP 0.311216f
C2 VTAIL VP 1.31266f
C3 VN VDD1 0.153766f
C4 VDD2 VN 1.0736f
C5 VN VTAIL 1.29855f
C6 VN VP 3.31859f
C7 VDD2 VDD1 0.767187f
C8 VDD1 VTAIL 3.53261f
C9 VDD2 VTAIL 3.57348f
C10 VDD2 B 2.442323f
C11 VDD1 B 2.648872f
C12 VTAIL B 2.894035f
C13 VN B 6.268318f
C14 VP B 5.318074f
C15 VDD2.t1 B 0.029442f
C16 VDD2.t4 B 0.029442f
C17 VDD2.n0 B 0.189413f
C18 VDD2.t5 B 0.029442f
C19 VDD2.t0 B 0.029442f
C20 VDD2.n1 B 0.189413f
C21 VDD2.n2 B 1.18454f
C22 VDD2.t6 B 0.029442f
C23 VDD2.t7 B 0.029442f
C24 VDD2.n3 B 0.188668f
C25 VDD2.n4 B 1.14643f
C26 VDD2.t2 B 0.029442f
C27 VDD2.t3 B 0.029442f
C28 VDD2.n5 B 0.189403f
C29 VN.n0 B 0.028611f
C30 VN.t3 B 0.094406f
C31 VN.n1 B 0.076874f
C32 VN.t6 B 0.105419f
C33 VN.n2 B 0.060226f
C34 VN.n3 B 0.119323f
C35 VN.t2 B 0.094406f
C36 VN.n4 B 0.070603f
C37 VN.n5 B 0.006492f
C38 VN.t7 B 0.094406f
C39 VN.n6 B 0.070427f
C40 VN.n7 B 0.022173f
C41 VN.n8 B 0.028611f
C42 VN.t5 B 0.094406f
C43 VN.n9 B 0.076874f
C44 VN.t0 B 0.094406f
C45 VN.t4 B 0.105419f
C46 VN.n10 B 0.060226f
C47 VN.n11 B 0.119323f
C48 VN.n12 B 0.070603f
C49 VN.n13 B 0.006492f
C50 VN.t1 B 0.094406f
C51 VN.n14 B 0.070427f
C52 VN.n15 B 0.81257f
C53 VDD1.t6 B 0.028035f
C54 VDD1.t5 B 0.028035f
C55 VDD1.n0 B 0.180628f
C56 VDD1.t0 B 0.028035f
C57 VDD1.t7 B 0.028035f
C58 VDD1.n1 B 0.180364f
C59 VDD1.t4 B 0.028035f
C60 VDD1.t1 B 0.028035f
C61 VDD1.n2 B 0.180364f
C62 VDD1.n3 B 1.16978f
C63 VDD1.t3 B 0.028035f
C64 VDD1.t2 B 0.028035f
C65 VDD1.n4 B 0.179654f
C66 VDD1.n5 B 1.11451f
C67 VTAIL.t1 B 0.028969f
C68 VTAIL.t4 B 0.028969f
C69 VTAIL.n0 B 0.158833f
C70 VTAIL.n1 B 0.195375f
C71 VTAIL.n2 B 0.026952f
C72 VTAIL.n3 B 0.063171f
C73 VTAIL.t6 B 0.045071f
C74 VTAIL.n4 B 0.046583f
C75 VTAIL.n5 B 0.013334f
C76 VTAIL.n6 B 0.010823f
C77 VTAIL.n7 B 0.123694f
C78 VTAIL.n8 B 0.029511f
C79 VTAIL.n9 B 0.100789f
C80 VTAIL.n10 B 0.026952f
C81 VTAIL.n11 B 0.063171f
C82 VTAIL.t13 B 0.045071f
C83 VTAIL.n12 B 0.046583f
C84 VTAIL.n13 B 0.013334f
C85 VTAIL.n14 B 0.010823f
C86 VTAIL.n15 B 0.123694f
C87 VTAIL.n16 B 0.029511f
C88 VTAIL.n17 B 0.100789f
C89 VTAIL.t11 B 0.028969f
C90 VTAIL.t8 B 0.028969f
C91 VTAIL.n18 B 0.158833f
C92 VTAIL.n19 B 0.242513f
C93 VTAIL.n20 B 0.026952f
C94 VTAIL.n21 B 0.063171f
C95 VTAIL.t14 B 0.045071f
C96 VTAIL.n22 B 0.046583f
C97 VTAIL.n23 B 0.013334f
C98 VTAIL.n24 B 0.010823f
C99 VTAIL.n25 B 0.123694f
C100 VTAIL.n26 B 0.029511f
C101 VTAIL.n27 B 0.496646f
C102 VTAIL.n28 B 0.026952f
C103 VTAIL.n29 B 0.063171f
C104 VTAIL.t3 B 0.045071f
C105 VTAIL.n30 B 0.046583f
C106 VTAIL.n31 B 0.013334f
C107 VTAIL.n32 B 0.010823f
C108 VTAIL.n33 B 0.123694f
C109 VTAIL.n34 B 0.029511f
C110 VTAIL.n35 B 0.496646f
C111 VTAIL.t2 B 0.028969f
C112 VTAIL.t7 B 0.028969f
C113 VTAIL.n36 B 0.158834f
C114 VTAIL.n37 B 0.242512f
C115 VTAIL.n38 B 0.026952f
C116 VTAIL.n39 B 0.063171f
C117 VTAIL.t0 B 0.045071f
C118 VTAIL.n40 B 0.046583f
C119 VTAIL.n41 B 0.013334f
C120 VTAIL.n42 B 0.010823f
C121 VTAIL.n43 B 0.123694f
C122 VTAIL.n44 B 0.029511f
C123 VTAIL.n45 B 0.100789f
C124 VTAIL.n46 B 0.026952f
C125 VTAIL.n47 B 0.063171f
C126 VTAIL.t12 B 0.045071f
C127 VTAIL.n48 B 0.046583f
C128 VTAIL.n49 B 0.013334f
C129 VTAIL.n50 B 0.010823f
C130 VTAIL.n51 B 0.123694f
C131 VTAIL.n52 B 0.029511f
C132 VTAIL.n53 B 0.100789f
C133 VTAIL.t10 B 0.028969f
C134 VTAIL.t9 B 0.028969f
C135 VTAIL.n54 B 0.158834f
C136 VTAIL.n55 B 0.242512f
C137 VTAIL.n56 B 0.026952f
C138 VTAIL.n57 B 0.063171f
C139 VTAIL.t15 B 0.045071f
C140 VTAIL.n58 B 0.046583f
C141 VTAIL.n59 B 0.013334f
C142 VTAIL.n60 B 0.010823f
C143 VTAIL.n61 B 0.123694f
C144 VTAIL.n62 B 0.029511f
C145 VTAIL.n63 B 0.496646f
C146 VTAIL.n64 B 0.026952f
C147 VTAIL.n65 B 0.063171f
C148 VTAIL.t5 B 0.045071f
C149 VTAIL.n66 B 0.046583f
C150 VTAIL.n67 B 0.013334f
C151 VTAIL.n68 B 0.010823f
C152 VTAIL.n69 B 0.123694f
C153 VTAIL.n70 B 0.029511f
C154 VTAIL.n71 B 0.492869f
C155 VP.n0 B 0.028964f
C156 VP.t0 B 0.095571f
C157 VP.n1 B 0.071474f
C158 VP.n2 B 0.028964f
C159 VP.t5 B 0.095571f
C160 VP.t4 B 0.095571f
C161 VP.n3 B 0.120795f
C162 VP.t2 B 0.095571f
C163 VP.t1 B 0.10672f
C164 VP.n4 B 0.060969f
C165 VP.n5 B 0.077823f
C166 VP.n6 B 0.071474f
C167 VP.n7 B 0.006573f
C168 VP.n8 B 0.071296f
C169 VP.n9 B 0.80329f
C170 VP.n10 B 0.834057f
C171 VP.t7 B 0.095571f
C172 VP.n11 B 0.071296f
C173 VP.n12 B 0.006573f
C174 VP.n13 B 0.028964f
C175 VP.n14 B 0.028964f
C176 VP.n15 B 0.028964f
C177 VP.t3 B 0.095571f
C178 VP.n16 B 0.071474f
C179 VP.n17 B 0.006573f
C180 VP.t6 B 0.095571f
C181 VP.n18 B 0.071296f
C182 VP.n19 B 0.022446f
.ends

