* NGSPICE file created from diff_pair_sample_1259.ext - technology: sky130A

.subckt diff_pair_sample_1259 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=0.2223 pd=1.92 as=0 ps=0 w=0.57 l=1.5
X1 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=0.2223 pd=1.92 as=0 ps=0 w=0.57 l=1.5
X2 VDD2.t1 VN.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.2223 pd=1.92 as=0.2223 ps=1.92 w=0.57 l=1.5
X3 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2223 pd=1.92 as=0 ps=0 w=0.57 l=1.5
X4 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.2223 pd=1.92 as=0.2223 ps=1.92 w=0.57 l=1.5
X5 VDD2.t0 VN.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2223 pd=1.92 as=0.2223 ps=1.92 w=0.57 l=1.5
X6 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2223 pd=1.92 as=0.2223 ps=1.92 w=0.57 l=1.5
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2223 pd=1.92 as=0 ps=0 w=0.57 l=1.5
R0 B.n292 B.n291 585
R1 B.n103 B.n51 585
R2 B.n102 B.n101 585
R3 B.n100 B.n99 585
R4 B.n98 B.n97 585
R5 B.n96 B.n95 585
R6 B.n94 B.n93 585
R7 B.n92 B.n91 585
R8 B.n90 B.n89 585
R9 B.n88 B.n87 585
R10 B.n86 B.n85 585
R11 B.n84 B.n83 585
R12 B.n82 B.n81 585
R13 B.n80 B.n79 585
R14 B.n78 B.n77 585
R15 B.n76 B.n75 585
R16 B.n74 B.n73 585
R17 B.n72 B.n71 585
R18 B.n70 B.n69 585
R19 B.n68 B.n67 585
R20 B.n66 B.n65 585
R21 B.n64 B.n63 585
R22 B.n62 B.n61 585
R23 B.n60 B.n59 585
R24 B.n39 B.n38 585
R25 B.n297 B.n296 585
R26 B.n290 B.n52 585
R27 B.n52 B.n36 585
R28 B.n289 B.n35 585
R29 B.n301 B.n35 585
R30 B.n288 B.n34 585
R31 B.n302 B.n34 585
R32 B.n287 B.n33 585
R33 B.n303 B.n33 585
R34 B.n286 B.n285 585
R35 B.n285 B.n29 585
R36 B.n284 B.n28 585
R37 B.n309 B.n28 585
R38 B.n283 B.n27 585
R39 B.n310 B.n27 585
R40 B.n282 B.n26 585
R41 B.n311 B.n26 585
R42 B.n281 B.n280 585
R43 B.n280 B.n22 585
R44 B.n279 B.n21 585
R45 B.n317 B.n21 585
R46 B.n278 B.n20 585
R47 B.n318 B.n20 585
R48 B.n277 B.n19 585
R49 B.n319 B.n19 585
R50 B.n276 B.n275 585
R51 B.n275 B.n15 585
R52 B.n274 B.n14 585
R53 B.n325 B.n14 585
R54 B.n273 B.n13 585
R55 B.n326 B.n13 585
R56 B.n272 B.n12 585
R57 B.n327 B.n12 585
R58 B.n271 B.n270 585
R59 B.n270 B.n8 585
R60 B.n269 B.n7 585
R61 B.n333 B.n7 585
R62 B.n268 B.n6 585
R63 B.n334 B.n6 585
R64 B.n267 B.n5 585
R65 B.n335 B.n5 585
R66 B.n266 B.n265 585
R67 B.n265 B.n4 585
R68 B.n264 B.n104 585
R69 B.n264 B.n263 585
R70 B.n254 B.n105 585
R71 B.n106 B.n105 585
R72 B.n256 B.n255 585
R73 B.n257 B.n256 585
R74 B.n253 B.n110 585
R75 B.n114 B.n110 585
R76 B.n252 B.n251 585
R77 B.n251 B.n250 585
R78 B.n112 B.n111 585
R79 B.n113 B.n112 585
R80 B.n243 B.n242 585
R81 B.n244 B.n243 585
R82 B.n241 B.n119 585
R83 B.n119 B.n118 585
R84 B.n240 B.n239 585
R85 B.n239 B.n238 585
R86 B.n121 B.n120 585
R87 B.n122 B.n121 585
R88 B.n231 B.n230 585
R89 B.n232 B.n231 585
R90 B.n229 B.n126 585
R91 B.n130 B.n126 585
R92 B.n228 B.n227 585
R93 B.n227 B.n226 585
R94 B.n128 B.n127 585
R95 B.n129 B.n128 585
R96 B.n219 B.n218 585
R97 B.n220 B.n219 585
R98 B.n217 B.n135 585
R99 B.n135 B.n134 585
R100 B.n216 B.n215 585
R101 B.n215 B.n214 585
R102 B.n137 B.n136 585
R103 B.n138 B.n137 585
R104 B.n210 B.n209 585
R105 B.n141 B.n140 585
R106 B.n206 B.n205 585
R107 B.n207 B.n206 585
R108 B.n204 B.n154 585
R109 B.n203 B.n202 585
R110 B.n201 B.n200 585
R111 B.n199 B.n198 585
R112 B.n197 B.n196 585
R113 B.n194 B.n193 585
R114 B.n192 B.n191 585
R115 B.n190 B.n189 585
R116 B.n188 B.n187 585
R117 B.n186 B.n185 585
R118 B.n184 B.n183 585
R119 B.n182 B.n181 585
R120 B.n180 B.n179 585
R121 B.n178 B.n177 585
R122 B.n176 B.n175 585
R123 B.n173 B.n172 585
R124 B.n171 B.n170 585
R125 B.n169 B.n168 585
R126 B.n167 B.n166 585
R127 B.n165 B.n164 585
R128 B.n163 B.n162 585
R129 B.n161 B.n160 585
R130 B.n159 B.n153 585
R131 B.n207 B.n153 585
R132 B.n211 B.n139 585
R133 B.n139 B.n138 585
R134 B.n213 B.n212 585
R135 B.n214 B.n213 585
R136 B.n133 B.n132 585
R137 B.n134 B.n133 585
R138 B.n222 B.n221 585
R139 B.n221 B.n220 585
R140 B.n223 B.n131 585
R141 B.n131 B.n129 585
R142 B.n225 B.n224 585
R143 B.n226 B.n225 585
R144 B.n125 B.n124 585
R145 B.n130 B.n125 585
R146 B.n234 B.n233 585
R147 B.n233 B.n232 585
R148 B.n235 B.n123 585
R149 B.n123 B.n122 585
R150 B.n237 B.n236 585
R151 B.n238 B.n237 585
R152 B.n117 B.n116 585
R153 B.n118 B.n117 585
R154 B.n246 B.n245 585
R155 B.n245 B.n244 585
R156 B.n247 B.n115 585
R157 B.n115 B.n113 585
R158 B.n249 B.n248 585
R159 B.n250 B.n249 585
R160 B.n109 B.n108 585
R161 B.n114 B.n109 585
R162 B.n259 B.n258 585
R163 B.n258 B.n257 585
R164 B.n260 B.n107 585
R165 B.n107 B.n106 585
R166 B.n262 B.n261 585
R167 B.n263 B.n262 585
R168 B.n2 B.n0 585
R169 B.n4 B.n2 585
R170 B.n3 B.n1 585
R171 B.n334 B.n3 585
R172 B.n332 B.n331 585
R173 B.n333 B.n332 585
R174 B.n330 B.n9 585
R175 B.n9 B.n8 585
R176 B.n329 B.n328 585
R177 B.n328 B.n327 585
R178 B.n11 B.n10 585
R179 B.n326 B.n11 585
R180 B.n324 B.n323 585
R181 B.n325 B.n324 585
R182 B.n322 B.n16 585
R183 B.n16 B.n15 585
R184 B.n321 B.n320 585
R185 B.n320 B.n319 585
R186 B.n18 B.n17 585
R187 B.n318 B.n18 585
R188 B.n316 B.n315 585
R189 B.n317 B.n316 585
R190 B.n314 B.n23 585
R191 B.n23 B.n22 585
R192 B.n313 B.n312 585
R193 B.n312 B.n311 585
R194 B.n25 B.n24 585
R195 B.n310 B.n25 585
R196 B.n308 B.n307 585
R197 B.n309 B.n308 585
R198 B.n306 B.n30 585
R199 B.n30 B.n29 585
R200 B.n305 B.n304 585
R201 B.n304 B.n303 585
R202 B.n32 B.n31 585
R203 B.n302 B.n32 585
R204 B.n300 B.n299 585
R205 B.n301 B.n300 585
R206 B.n298 B.n37 585
R207 B.n37 B.n36 585
R208 B.n337 B.n336 585
R209 B.n336 B.n335 585
R210 B.n209 B.n139 444.452
R211 B.n296 B.n37 444.452
R212 B.n153 B.n137 444.452
R213 B.n292 B.n52 444.452
R214 B.n157 B.t12 275.979
R215 B.n155 B.t15 275.979
R216 B.n56 B.t4 275.979
R217 B.n53 B.t7 275.979
R218 B.n294 B.n293 256.663
R219 B.n294 B.n50 256.663
R220 B.n294 B.n49 256.663
R221 B.n294 B.n48 256.663
R222 B.n294 B.n47 256.663
R223 B.n294 B.n46 256.663
R224 B.n294 B.n45 256.663
R225 B.n294 B.n44 256.663
R226 B.n294 B.n43 256.663
R227 B.n294 B.n42 256.663
R228 B.n294 B.n41 256.663
R229 B.n294 B.n40 256.663
R230 B.n295 B.n294 256.663
R231 B.n208 B.n207 256.663
R232 B.n207 B.n142 256.663
R233 B.n207 B.n143 256.663
R234 B.n207 B.n144 256.663
R235 B.n207 B.n145 256.663
R236 B.n207 B.n146 256.663
R237 B.n207 B.n147 256.663
R238 B.n207 B.n148 256.663
R239 B.n207 B.n149 256.663
R240 B.n207 B.n150 256.663
R241 B.n207 B.n151 256.663
R242 B.n207 B.n152 256.663
R243 B.n158 B.t11 240.488
R244 B.n156 B.t14 240.488
R245 B.n57 B.t5 240.488
R246 B.n54 B.t8 240.488
R247 B.n207 B.n138 216.424
R248 B.n294 B.n36 216.424
R249 B.n157 B.t9 207.549
R250 B.n155 B.t13 207.549
R251 B.n56 B.t2 207.549
R252 B.n53 B.t6 207.549
R253 B.n213 B.n139 163.367
R254 B.n213 B.n133 163.367
R255 B.n221 B.n133 163.367
R256 B.n221 B.n131 163.367
R257 B.n225 B.n131 163.367
R258 B.n225 B.n125 163.367
R259 B.n233 B.n125 163.367
R260 B.n233 B.n123 163.367
R261 B.n237 B.n123 163.367
R262 B.n237 B.n117 163.367
R263 B.n245 B.n117 163.367
R264 B.n245 B.n115 163.367
R265 B.n249 B.n115 163.367
R266 B.n249 B.n109 163.367
R267 B.n258 B.n109 163.367
R268 B.n258 B.n107 163.367
R269 B.n262 B.n107 163.367
R270 B.n262 B.n2 163.367
R271 B.n336 B.n2 163.367
R272 B.n336 B.n3 163.367
R273 B.n332 B.n3 163.367
R274 B.n332 B.n9 163.367
R275 B.n328 B.n9 163.367
R276 B.n328 B.n11 163.367
R277 B.n324 B.n11 163.367
R278 B.n324 B.n16 163.367
R279 B.n320 B.n16 163.367
R280 B.n320 B.n18 163.367
R281 B.n316 B.n18 163.367
R282 B.n316 B.n23 163.367
R283 B.n312 B.n23 163.367
R284 B.n312 B.n25 163.367
R285 B.n308 B.n25 163.367
R286 B.n308 B.n30 163.367
R287 B.n304 B.n30 163.367
R288 B.n304 B.n32 163.367
R289 B.n300 B.n32 163.367
R290 B.n300 B.n37 163.367
R291 B.n206 B.n141 163.367
R292 B.n206 B.n154 163.367
R293 B.n202 B.n201 163.367
R294 B.n198 B.n197 163.367
R295 B.n193 B.n192 163.367
R296 B.n189 B.n188 163.367
R297 B.n185 B.n184 163.367
R298 B.n181 B.n180 163.367
R299 B.n177 B.n176 163.367
R300 B.n172 B.n171 163.367
R301 B.n168 B.n167 163.367
R302 B.n164 B.n163 163.367
R303 B.n160 B.n153 163.367
R304 B.n215 B.n137 163.367
R305 B.n215 B.n135 163.367
R306 B.n219 B.n135 163.367
R307 B.n219 B.n128 163.367
R308 B.n227 B.n128 163.367
R309 B.n227 B.n126 163.367
R310 B.n231 B.n126 163.367
R311 B.n231 B.n121 163.367
R312 B.n239 B.n121 163.367
R313 B.n239 B.n119 163.367
R314 B.n243 B.n119 163.367
R315 B.n243 B.n112 163.367
R316 B.n251 B.n112 163.367
R317 B.n251 B.n110 163.367
R318 B.n256 B.n110 163.367
R319 B.n256 B.n105 163.367
R320 B.n264 B.n105 163.367
R321 B.n265 B.n264 163.367
R322 B.n265 B.n5 163.367
R323 B.n6 B.n5 163.367
R324 B.n7 B.n6 163.367
R325 B.n270 B.n7 163.367
R326 B.n270 B.n12 163.367
R327 B.n13 B.n12 163.367
R328 B.n14 B.n13 163.367
R329 B.n275 B.n14 163.367
R330 B.n275 B.n19 163.367
R331 B.n20 B.n19 163.367
R332 B.n21 B.n20 163.367
R333 B.n280 B.n21 163.367
R334 B.n280 B.n26 163.367
R335 B.n27 B.n26 163.367
R336 B.n28 B.n27 163.367
R337 B.n285 B.n28 163.367
R338 B.n285 B.n33 163.367
R339 B.n34 B.n33 163.367
R340 B.n35 B.n34 163.367
R341 B.n52 B.n35 163.367
R342 B.n59 B.n39 163.367
R343 B.n63 B.n62 163.367
R344 B.n67 B.n66 163.367
R345 B.n71 B.n70 163.367
R346 B.n75 B.n74 163.367
R347 B.n79 B.n78 163.367
R348 B.n83 B.n82 163.367
R349 B.n87 B.n86 163.367
R350 B.n91 B.n90 163.367
R351 B.n95 B.n94 163.367
R352 B.n99 B.n98 163.367
R353 B.n101 B.n51 163.367
R354 B.n214 B.n138 127.974
R355 B.n214 B.n134 127.974
R356 B.n220 B.n134 127.974
R357 B.n220 B.n129 127.974
R358 B.n226 B.n129 127.974
R359 B.n226 B.n130 127.974
R360 B.n232 B.n122 127.974
R361 B.n238 B.n122 127.974
R362 B.n238 B.n118 127.974
R363 B.n244 B.n118 127.974
R364 B.n244 B.n113 127.974
R365 B.n250 B.n113 127.974
R366 B.n250 B.n114 127.974
R367 B.n257 B.n106 127.974
R368 B.n263 B.n106 127.974
R369 B.n263 B.n4 127.974
R370 B.n335 B.n4 127.974
R371 B.n335 B.n334 127.974
R372 B.n334 B.n333 127.974
R373 B.n333 B.n8 127.974
R374 B.n327 B.n8 127.974
R375 B.n326 B.n325 127.974
R376 B.n325 B.n15 127.974
R377 B.n319 B.n15 127.974
R378 B.n319 B.n318 127.974
R379 B.n318 B.n317 127.974
R380 B.n317 B.n22 127.974
R381 B.n311 B.n22 127.974
R382 B.n310 B.n309 127.974
R383 B.n309 B.n29 127.974
R384 B.n303 B.n29 127.974
R385 B.n303 B.n302 127.974
R386 B.n302 B.n301 127.974
R387 B.n301 B.n36 127.974
R388 B.n232 B.t10 112.918
R389 B.n311 B.t3 112.918
R390 B.n114 B.t0 90.3341
R391 B.t1 B.n326 90.3341
R392 B.n209 B.n208 71.676
R393 B.n154 B.n142 71.676
R394 B.n201 B.n143 71.676
R395 B.n197 B.n144 71.676
R396 B.n192 B.n145 71.676
R397 B.n188 B.n146 71.676
R398 B.n184 B.n147 71.676
R399 B.n180 B.n148 71.676
R400 B.n176 B.n149 71.676
R401 B.n171 B.n150 71.676
R402 B.n167 B.n151 71.676
R403 B.n163 B.n152 71.676
R404 B.n296 B.n295 71.676
R405 B.n59 B.n40 71.676
R406 B.n63 B.n41 71.676
R407 B.n67 B.n42 71.676
R408 B.n71 B.n43 71.676
R409 B.n75 B.n44 71.676
R410 B.n79 B.n45 71.676
R411 B.n83 B.n46 71.676
R412 B.n87 B.n47 71.676
R413 B.n91 B.n48 71.676
R414 B.n95 B.n49 71.676
R415 B.n99 B.n50 71.676
R416 B.n293 B.n51 71.676
R417 B.n293 B.n292 71.676
R418 B.n101 B.n50 71.676
R419 B.n98 B.n49 71.676
R420 B.n94 B.n48 71.676
R421 B.n90 B.n47 71.676
R422 B.n86 B.n46 71.676
R423 B.n82 B.n45 71.676
R424 B.n78 B.n44 71.676
R425 B.n74 B.n43 71.676
R426 B.n70 B.n42 71.676
R427 B.n66 B.n41 71.676
R428 B.n62 B.n40 71.676
R429 B.n295 B.n39 71.676
R430 B.n208 B.n141 71.676
R431 B.n202 B.n142 71.676
R432 B.n198 B.n143 71.676
R433 B.n193 B.n144 71.676
R434 B.n189 B.n145 71.676
R435 B.n185 B.n146 71.676
R436 B.n181 B.n147 71.676
R437 B.n177 B.n148 71.676
R438 B.n172 B.n149 71.676
R439 B.n168 B.n150 71.676
R440 B.n164 B.n151 71.676
R441 B.n160 B.n152 71.676
R442 B.n174 B.n158 59.5399
R443 B.n195 B.n156 59.5399
R444 B.n58 B.n57 59.5399
R445 B.n55 B.n54 59.5399
R446 B.n257 B.t0 37.6395
R447 B.n327 B.t1 37.6395
R448 B.n158 B.n157 35.4914
R449 B.n156 B.n155 35.4914
R450 B.n57 B.n56 35.4914
R451 B.n54 B.n53 35.4914
R452 B.n291 B.n290 28.8785
R453 B.n298 B.n297 28.8785
R454 B.n159 B.n136 28.8785
R455 B.n211 B.n210 28.8785
R456 B B.n337 18.0485
R457 B.n130 B.t10 15.0561
R458 B.t3 B.n310 15.0561
R459 B.n297 B.n38 10.6151
R460 B.n60 B.n38 10.6151
R461 B.n61 B.n60 10.6151
R462 B.n64 B.n61 10.6151
R463 B.n65 B.n64 10.6151
R464 B.n68 B.n65 10.6151
R465 B.n69 B.n68 10.6151
R466 B.n73 B.n72 10.6151
R467 B.n76 B.n73 10.6151
R468 B.n77 B.n76 10.6151
R469 B.n80 B.n77 10.6151
R470 B.n81 B.n80 10.6151
R471 B.n84 B.n81 10.6151
R472 B.n85 B.n84 10.6151
R473 B.n88 B.n85 10.6151
R474 B.n89 B.n88 10.6151
R475 B.n93 B.n92 10.6151
R476 B.n96 B.n93 10.6151
R477 B.n97 B.n96 10.6151
R478 B.n100 B.n97 10.6151
R479 B.n102 B.n100 10.6151
R480 B.n103 B.n102 10.6151
R481 B.n291 B.n103 10.6151
R482 B.n216 B.n136 10.6151
R483 B.n217 B.n216 10.6151
R484 B.n218 B.n217 10.6151
R485 B.n218 B.n127 10.6151
R486 B.n228 B.n127 10.6151
R487 B.n229 B.n228 10.6151
R488 B.n230 B.n229 10.6151
R489 B.n230 B.n120 10.6151
R490 B.n240 B.n120 10.6151
R491 B.n241 B.n240 10.6151
R492 B.n242 B.n241 10.6151
R493 B.n242 B.n111 10.6151
R494 B.n252 B.n111 10.6151
R495 B.n253 B.n252 10.6151
R496 B.n255 B.n253 10.6151
R497 B.n255 B.n254 10.6151
R498 B.n254 B.n104 10.6151
R499 B.n266 B.n104 10.6151
R500 B.n267 B.n266 10.6151
R501 B.n268 B.n267 10.6151
R502 B.n269 B.n268 10.6151
R503 B.n271 B.n269 10.6151
R504 B.n272 B.n271 10.6151
R505 B.n273 B.n272 10.6151
R506 B.n274 B.n273 10.6151
R507 B.n276 B.n274 10.6151
R508 B.n277 B.n276 10.6151
R509 B.n278 B.n277 10.6151
R510 B.n279 B.n278 10.6151
R511 B.n281 B.n279 10.6151
R512 B.n282 B.n281 10.6151
R513 B.n283 B.n282 10.6151
R514 B.n284 B.n283 10.6151
R515 B.n286 B.n284 10.6151
R516 B.n287 B.n286 10.6151
R517 B.n288 B.n287 10.6151
R518 B.n289 B.n288 10.6151
R519 B.n290 B.n289 10.6151
R520 B.n210 B.n140 10.6151
R521 B.n205 B.n140 10.6151
R522 B.n205 B.n204 10.6151
R523 B.n204 B.n203 10.6151
R524 B.n203 B.n200 10.6151
R525 B.n200 B.n199 10.6151
R526 B.n199 B.n196 10.6151
R527 B.n194 B.n191 10.6151
R528 B.n191 B.n190 10.6151
R529 B.n190 B.n187 10.6151
R530 B.n187 B.n186 10.6151
R531 B.n186 B.n183 10.6151
R532 B.n183 B.n182 10.6151
R533 B.n182 B.n179 10.6151
R534 B.n179 B.n178 10.6151
R535 B.n178 B.n175 10.6151
R536 B.n173 B.n170 10.6151
R537 B.n170 B.n169 10.6151
R538 B.n169 B.n166 10.6151
R539 B.n166 B.n165 10.6151
R540 B.n165 B.n162 10.6151
R541 B.n162 B.n161 10.6151
R542 B.n161 B.n159 10.6151
R543 B.n212 B.n211 10.6151
R544 B.n212 B.n132 10.6151
R545 B.n222 B.n132 10.6151
R546 B.n223 B.n222 10.6151
R547 B.n224 B.n223 10.6151
R548 B.n224 B.n124 10.6151
R549 B.n234 B.n124 10.6151
R550 B.n235 B.n234 10.6151
R551 B.n236 B.n235 10.6151
R552 B.n236 B.n116 10.6151
R553 B.n246 B.n116 10.6151
R554 B.n247 B.n246 10.6151
R555 B.n248 B.n247 10.6151
R556 B.n248 B.n108 10.6151
R557 B.n259 B.n108 10.6151
R558 B.n260 B.n259 10.6151
R559 B.n261 B.n260 10.6151
R560 B.n261 B.n0 10.6151
R561 B.n331 B.n1 10.6151
R562 B.n331 B.n330 10.6151
R563 B.n330 B.n329 10.6151
R564 B.n329 B.n10 10.6151
R565 B.n323 B.n10 10.6151
R566 B.n323 B.n322 10.6151
R567 B.n322 B.n321 10.6151
R568 B.n321 B.n17 10.6151
R569 B.n315 B.n17 10.6151
R570 B.n315 B.n314 10.6151
R571 B.n314 B.n313 10.6151
R572 B.n313 B.n24 10.6151
R573 B.n307 B.n24 10.6151
R574 B.n307 B.n306 10.6151
R575 B.n306 B.n305 10.6151
R576 B.n305 B.n31 10.6151
R577 B.n299 B.n31 10.6151
R578 B.n299 B.n298 10.6151
R579 B.n69 B.n58 9.36635
R580 B.n92 B.n55 9.36635
R581 B.n196 B.n195 9.36635
R582 B.n174 B.n173 9.36635
R583 B.n337 B.n0 2.81026
R584 B.n337 B.n1 2.81026
R585 B.n72 B.n58 1.24928
R586 B.n89 B.n55 1.24928
R587 B.n195 B.n194 1.24928
R588 B.n175 B.n174 1.24928
R589 VN VN.t1 149.477
R590 VN VN.t0 116.257
R591 VTAIL.n3 VTAIL.t2 251.34
R592 VTAIL.n0 VTAIL.t0 251.34
R593 VTAIL.n2 VTAIL.t1 251.34
R594 VTAIL.n1 VTAIL.t3 251.34
R595 VTAIL.n1 VTAIL.n0 16.0134
R596 VTAIL.n3 VTAIL.n2 14.4358
R597 VTAIL.n2 VTAIL.n1 1.25912
R598 VTAIL VTAIL.n0 0.922914
R599 VTAIL VTAIL.n3 0.336707
R600 VDD2.n0 VDD2.t1 295.325
R601 VDD2.n0 VDD2.t0 268.019
R602 VDD2 VDD2.n0 0.453086
R603 VP.n0 VP.t0 149.191
R604 VP.n0 VP.t1 116.112
R605 VP VP.n0 0.146778
R606 VDD1 VDD1.t0 296.245
R607 VDD1 VDD1.t1 268.471
C0 VTAIL VDD2 1.71647f
C1 VTAIL VN 0.665334f
C2 VP VTAIL 0.679455f
C3 VDD1 VDD2 0.54415f
C4 VDD1 VN 0.156021f
C5 VP VDD1 0.494804f
C6 VN VDD2 0.357251f
C7 VP VDD2 0.295445f
C8 VP VN 2.82999f
C9 VDD1 VTAIL 1.6707f
C10 VDD2 B 1.87838f
C11 VDD1 B 2.0377f
C12 VTAIL B 1.86327f
C13 VN B 6.16166f
C14 VP B 3.999485f
C15 VP.t0 B 0.49318f
C16 VP.t1 B 0.24092f
C17 VP.n0 B 2.02504f
C18 VN.t0 B 0.236386f
C19 VN.t1 B 0.490344f
.ends

