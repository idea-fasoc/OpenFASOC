* NGSPICE file created from diff_pair_sample_0010.ext - technology: sky130A

.subckt diff_pair_sample_0010 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=2.0319 pd=11.2 as=0 ps=0 w=5.21 l=1.84
X1 VTAIL.t16 VP.t0 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=0.85965 pd=5.54 as=0.85965 ps=5.54 w=5.21 l=1.84
X2 VDD1.t2 VP.t1 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=2.0319 pd=11.2 as=0.85965 ps=5.54 w=5.21 l=1.84
X3 VTAIL.t14 VP.t2 VDD1.t3 B.t8 sky130_fd_pr__nfet_01v8 ad=0.85965 pd=5.54 as=0.85965 ps=5.54 w=5.21 l=1.84
X4 VDD1.t4 VP.t3 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=0.85965 pd=5.54 as=0.85965 ps=5.54 w=5.21 l=1.84
X5 VTAIL.t6 VN.t0 VDD2.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=0.85965 pd=5.54 as=0.85965 ps=5.54 w=5.21 l=1.84
X6 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=2.0319 pd=11.2 as=0 ps=0 w=5.21 l=1.84
X7 VTAIL.t2 VN.t1 VDD2.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=0.85965 pd=5.54 as=0.85965 ps=5.54 w=5.21 l=1.84
X8 VDD1.t5 VP.t4 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=0.85965 pd=5.54 as=2.0319 ps=11.2 w=5.21 l=1.84
X9 VTAIL.t3 VN.t2 VDD2.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=0.85965 pd=5.54 as=0.85965 ps=5.54 w=5.21 l=1.84
X10 VDD2.t6 VN.t3 VTAIL.t18 B.t1 sky130_fd_pr__nfet_01v8 ad=0.85965 pd=5.54 as=2.0319 ps=11.2 w=5.21 l=1.84
X11 VTAIL.t11 VP.t5 VDD1.t1 B.t9 sky130_fd_pr__nfet_01v8 ad=0.85965 pd=5.54 as=0.85965 ps=5.54 w=5.21 l=1.84
X12 VDD2.t5 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.85965 pd=5.54 as=0.85965 ps=5.54 w=5.21 l=1.84
X13 VTAIL.t10 VP.t6 VDD1.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=0.85965 pd=5.54 as=0.85965 ps=5.54 w=5.21 l=1.84
X14 VDD1.t7 VP.t7 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=0.85965 pd=5.54 as=2.0319 ps=11.2 w=5.21 l=1.84
X15 VDD2.t4 VN.t5 VTAIL.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=0.85965 pd=5.54 as=2.0319 ps=11.2 w=5.21 l=1.84
X16 VDD1.t8 VP.t8 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=0.85965 pd=5.54 as=0.85965 ps=5.54 w=5.21 l=1.84
X17 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=2.0319 pd=11.2 as=0 ps=0 w=5.21 l=1.84
X18 VDD1.t6 VP.t9 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=2.0319 pd=11.2 as=0.85965 ps=5.54 w=5.21 l=1.84
X19 VTAIL.t19 VN.t6 VDD2.t3 B.t8 sky130_fd_pr__nfet_01v8 ad=0.85965 pd=5.54 as=0.85965 ps=5.54 w=5.21 l=1.84
X20 VDD2.t2 VN.t7 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.0319 pd=11.2 as=0.85965 ps=5.54 w=5.21 l=1.84
X21 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.0319 pd=11.2 as=0 ps=0 w=5.21 l=1.84
X22 VDD2.t1 VN.t8 VTAIL.t17 B.t7 sky130_fd_pr__nfet_01v8 ad=2.0319 pd=11.2 as=0.85965 ps=5.54 w=5.21 l=1.84
X23 VDD2.t0 VN.t9 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.85965 pd=5.54 as=0.85965 ps=5.54 w=5.21 l=1.84
R0 B.n545 B.n544 585
R1 B.n545 B.n86 585
R2 B.n548 B.n547 585
R3 B.n549 B.n117 585
R4 B.n551 B.n550 585
R5 B.n553 B.n116 585
R6 B.n556 B.n555 585
R7 B.n557 B.n115 585
R8 B.n559 B.n558 585
R9 B.n561 B.n114 585
R10 B.n564 B.n563 585
R11 B.n565 B.n113 585
R12 B.n567 B.n566 585
R13 B.n569 B.n112 585
R14 B.n572 B.n571 585
R15 B.n573 B.n111 585
R16 B.n575 B.n574 585
R17 B.n577 B.n110 585
R18 B.n580 B.n579 585
R19 B.n581 B.n109 585
R20 B.n583 B.n582 585
R21 B.n585 B.n108 585
R22 B.n588 B.n587 585
R23 B.n590 B.n105 585
R24 B.n592 B.n591 585
R25 B.n594 B.n104 585
R26 B.n597 B.n596 585
R27 B.n598 B.n103 585
R28 B.n600 B.n599 585
R29 B.n602 B.n102 585
R30 B.n604 B.n603 585
R31 B.n606 B.n605 585
R32 B.n609 B.n608 585
R33 B.n610 B.n97 585
R34 B.n612 B.n611 585
R35 B.n614 B.n96 585
R36 B.n617 B.n616 585
R37 B.n618 B.n95 585
R38 B.n620 B.n619 585
R39 B.n622 B.n94 585
R40 B.n625 B.n624 585
R41 B.n626 B.n93 585
R42 B.n628 B.n627 585
R43 B.n630 B.n92 585
R44 B.n633 B.n632 585
R45 B.n634 B.n91 585
R46 B.n636 B.n635 585
R47 B.n638 B.n90 585
R48 B.n641 B.n640 585
R49 B.n642 B.n89 585
R50 B.n644 B.n643 585
R51 B.n646 B.n88 585
R52 B.n649 B.n648 585
R53 B.n650 B.n87 585
R54 B.n543 B.n85 585
R55 B.n653 B.n85 585
R56 B.n542 B.n84 585
R57 B.n654 B.n84 585
R58 B.n541 B.n83 585
R59 B.n655 B.n83 585
R60 B.n540 B.n539 585
R61 B.n539 B.n79 585
R62 B.n538 B.n78 585
R63 B.n661 B.n78 585
R64 B.n537 B.n77 585
R65 B.n662 B.n77 585
R66 B.n536 B.n76 585
R67 B.n663 B.n76 585
R68 B.n535 B.n534 585
R69 B.n534 B.n72 585
R70 B.n533 B.n71 585
R71 B.n669 B.n71 585
R72 B.n532 B.n70 585
R73 B.n670 B.n70 585
R74 B.n531 B.n69 585
R75 B.n671 B.n69 585
R76 B.n530 B.n529 585
R77 B.n529 B.n65 585
R78 B.n528 B.n64 585
R79 B.n677 B.n64 585
R80 B.n527 B.n63 585
R81 B.n678 B.n63 585
R82 B.n526 B.n62 585
R83 B.n679 B.n62 585
R84 B.n525 B.n524 585
R85 B.n524 B.n58 585
R86 B.n523 B.n57 585
R87 B.n685 B.n57 585
R88 B.n522 B.n56 585
R89 B.n686 B.n56 585
R90 B.n521 B.n55 585
R91 B.n687 B.n55 585
R92 B.n520 B.n519 585
R93 B.n519 B.n51 585
R94 B.n518 B.n50 585
R95 B.n693 B.n50 585
R96 B.n517 B.n49 585
R97 B.n694 B.n49 585
R98 B.n516 B.n48 585
R99 B.n695 B.n48 585
R100 B.n515 B.n514 585
R101 B.n514 B.n44 585
R102 B.n513 B.n43 585
R103 B.n701 B.n43 585
R104 B.n512 B.n42 585
R105 B.n702 B.n42 585
R106 B.n511 B.n41 585
R107 B.n703 B.n41 585
R108 B.n510 B.n509 585
R109 B.n509 B.n37 585
R110 B.n508 B.n36 585
R111 B.n709 B.n36 585
R112 B.n507 B.n35 585
R113 B.n710 B.n35 585
R114 B.n506 B.n34 585
R115 B.n711 B.n34 585
R116 B.n505 B.n504 585
R117 B.n504 B.n30 585
R118 B.n503 B.n29 585
R119 B.n717 B.n29 585
R120 B.n502 B.n28 585
R121 B.n718 B.n28 585
R122 B.n501 B.n27 585
R123 B.n719 B.n27 585
R124 B.n500 B.n499 585
R125 B.n499 B.n26 585
R126 B.n498 B.n22 585
R127 B.n725 B.n22 585
R128 B.n497 B.n21 585
R129 B.n726 B.n21 585
R130 B.n496 B.n20 585
R131 B.n727 B.n20 585
R132 B.n495 B.n494 585
R133 B.n494 B.n16 585
R134 B.n493 B.n15 585
R135 B.n733 B.n15 585
R136 B.n492 B.n14 585
R137 B.n734 B.n14 585
R138 B.n491 B.n13 585
R139 B.n735 B.n13 585
R140 B.n490 B.n489 585
R141 B.n489 B.n12 585
R142 B.n488 B.n487 585
R143 B.n488 B.n8 585
R144 B.n486 B.n7 585
R145 B.n742 B.n7 585
R146 B.n485 B.n6 585
R147 B.n743 B.n6 585
R148 B.n484 B.n5 585
R149 B.n744 B.n5 585
R150 B.n483 B.n482 585
R151 B.n482 B.n4 585
R152 B.n481 B.n118 585
R153 B.n481 B.n480 585
R154 B.n471 B.n119 585
R155 B.n120 B.n119 585
R156 B.n473 B.n472 585
R157 B.n474 B.n473 585
R158 B.n470 B.n124 585
R159 B.n128 B.n124 585
R160 B.n469 B.n468 585
R161 B.n468 B.n467 585
R162 B.n126 B.n125 585
R163 B.n127 B.n126 585
R164 B.n460 B.n459 585
R165 B.n461 B.n460 585
R166 B.n458 B.n133 585
R167 B.n133 B.n132 585
R168 B.n457 B.n456 585
R169 B.n456 B.n455 585
R170 B.n135 B.n134 585
R171 B.n448 B.n135 585
R172 B.n447 B.n446 585
R173 B.n449 B.n447 585
R174 B.n445 B.n140 585
R175 B.n140 B.n139 585
R176 B.n444 B.n443 585
R177 B.n443 B.n442 585
R178 B.n142 B.n141 585
R179 B.n143 B.n142 585
R180 B.n435 B.n434 585
R181 B.n436 B.n435 585
R182 B.n433 B.n148 585
R183 B.n148 B.n147 585
R184 B.n432 B.n431 585
R185 B.n431 B.n430 585
R186 B.n150 B.n149 585
R187 B.n151 B.n150 585
R188 B.n423 B.n422 585
R189 B.n424 B.n423 585
R190 B.n421 B.n156 585
R191 B.n156 B.n155 585
R192 B.n420 B.n419 585
R193 B.n419 B.n418 585
R194 B.n158 B.n157 585
R195 B.n159 B.n158 585
R196 B.n411 B.n410 585
R197 B.n412 B.n411 585
R198 B.n409 B.n164 585
R199 B.n164 B.n163 585
R200 B.n408 B.n407 585
R201 B.n407 B.n406 585
R202 B.n166 B.n165 585
R203 B.n167 B.n166 585
R204 B.n399 B.n398 585
R205 B.n400 B.n399 585
R206 B.n397 B.n172 585
R207 B.n172 B.n171 585
R208 B.n396 B.n395 585
R209 B.n395 B.n394 585
R210 B.n174 B.n173 585
R211 B.n175 B.n174 585
R212 B.n387 B.n386 585
R213 B.n388 B.n387 585
R214 B.n385 B.n180 585
R215 B.n180 B.n179 585
R216 B.n384 B.n383 585
R217 B.n383 B.n382 585
R218 B.n182 B.n181 585
R219 B.n183 B.n182 585
R220 B.n375 B.n374 585
R221 B.n376 B.n375 585
R222 B.n373 B.n188 585
R223 B.n188 B.n187 585
R224 B.n372 B.n371 585
R225 B.n371 B.n370 585
R226 B.n190 B.n189 585
R227 B.n191 B.n190 585
R228 B.n363 B.n362 585
R229 B.n364 B.n363 585
R230 B.n361 B.n196 585
R231 B.n196 B.n195 585
R232 B.n360 B.n359 585
R233 B.n359 B.n358 585
R234 B.n198 B.n197 585
R235 B.n199 B.n198 585
R236 B.n351 B.n350 585
R237 B.n352 B.n351 585
R238 B.n349 B.n204 585
R239 B.n204 B.n203 585
R240 B.n348 B.n347 585
R241 B.n347 B.n346 585
R242 B.n343 B.n208 585
R243 B.n342 B.n341 585
R244 B.n339 B.n209 585
R245 B.n339 B.n207 585
R246 B.n338 B.n337 585
R247 B.n336 B.n335 585
R248 B.n334 B.n211 585
R249 B.n332 B.n331 585
R250 B.n330 B.n212 585
R251 B.n329 B.n328 585
R252 B.n326 B.n213 585
R253 B.n324 B.n323 585
R254 B.n322 B.n214 585
R255 B.n321 B.n320 585
R256 B.n318 B.n215 585
R257 B.n316 B.n315 585
R258 B.n314 B.n216 585
R259 B.n313 B.n312 585
R260 B.n310 B.n217 585
R261 B.n308 B.n307 585
R262 B.n306 B.n218 585
R263 B.n305 B.n304 585
R264 B.n302 B.n219 585
R265 B.n300 B.n299 585
R266 B.n298 B.n220 585
R267 B.n297 B.n296 585
R268 B.n294 B.n224 585
R269 B.n292 B.n291 585
R270 B.n290 B.n225 585
R271 B.n289 B.n288 585
R272 B.n286 B.n226 585
R273 B.n284 B.n283 585
R274 B.n281 B.n227 585
R275 B.n280 B.n279 585
R276 B.n277 B.n230 585
R277 B.n275 B.n274 585
R278 B.n273 B.n231 585
R279 B.n272 B.n271 585
R280 B.n269 B.n232 585
R281 B.n267 B.n266 585
R282 B.n265 B.n233 585
R283 B.n264 B.n263 585
R284 B.n261 B.n234 585
R285 B.n259 B.n258 585
R286 B.n257 B.n235 585
R287 B.n256 B.n255 585
R288 B.n253 B.n236 585
R289 B.n251 B.n250 585
R290 B.n249 B.n237 585
R291 B.n248 B.n247 585
R292 B.n245 B.n238 585
R293 B.n243 B.n242 585
R294 B.n241 B.n240 585
R295 B.n206 B.n205 585
R296 B.n345 B.n344 585
R297 B.n346 B.n345 585
R298 B.n202 B.n201 585
R299 B.n203 B.n202 585
R300 B.n354 B.n353 585
R301 B.n353 B.n352 585
R302 B.n355 B.n200 585
R303 B.n200 B.n199 585
R304 B.n357 B.n356 585
R305 B.n358 B.n357 585
R306 B.n194 B.n193 585
R307 B.n195 B.n194 585
R308 B.n366 B.n365 585
R309 B.n365 B.n364 585
R310 B.n367 B.n192 585
R311 B.n192 B.n191 585
R312 B.n369 B.n368 585
R313 B.n370 B.n369 585
R314 B.n186 B.n185 585
R315 B.n187 B.n186 585
R316 B.n378 B.n377 585
R317 B.n377 B.n376 585
R318 B.n379 B.n184 585
R319 B.n184 B.n183 585
R320 B.n381 B.n380 585
R321 B.n382 B.n381 585
R322 B.n178 B.n177 585
R323 B.n179 B.n178 585
R324 B.n390 B.n389 585
R325 B.n389 B.n388 585
R326 B.n391 B.n176 585
R327 B.n176 B.n175 585
R328 B.n393 B.n392 585
R329 B.n394 B.n393 585
R330 B.n170 B.n169 585
R331 B.n171 B.n170 585
R332 B.n402 B.n401 585
R333 B.n401 B.n400 585
R334 B.n403 B.n168 585
R335 B.n168 B.n167 585
R336 B.n405 B.n404 585
R337 B.n406 B.n405 585
R338 B.n162 B.n161 585
R339 B.n163 B.n162 585
R340 B.n414 B.n413 585
R341 B.n413 B.n412 585
R342 B.n415 B.n160 585
R343 B.n160 B.n159 585
R344 B.n417 B.n416 585
R345 B.n418 B.n417 585
R346 B.n154 B.n153 585
R347 B.n155 B.n154 585
R348 B.n426 B.n425 585
R349 B.n425 B.n424 585
R350 B.n427 B.n152 585
R351 B.n152 B.n151 585
R352 B.n429 B.n428 585
R353 B.n430 B.n429 585
R354 B.n146 B.n145 585
R355 B.n147 B.n146 585
R356 B.n438 B.n437 585
R357 B.n437 B.n436 585
R358 B.n439 B.n144 585
R359 B.n144 B.n143 585
R360 B.n441 B.n440 585
R361 B.n442 B.n441 585
R362 B.n138 B.n137 585
R363 B.n139 B.n138 585
R364 B.n451 B.n450 585
R365 B.n450 B.n449 585
R366 B.n452 B.n136 585
R367 B.n448 B.n136 585
R368 B.n454 B.n453 585
R369 B.n455 B.n454 585
R370 B.n131 B.n130 585
R371 B.n132 B.n131 585
R372 B.n463 B.n462 585
R373 B.n462 B.n461 585
R374 B.n464 B.n129 585
R375 B.n129 B.n127 585
R376 B.n466 B.n465 585
R377 B.n467 B.n466 585
R378 B.n123 B.n122 585
R379 B.n128 B.n123 585
R380 B.n476 B.n475 585
R381 B.n475 B.n474 585
R382 B.n477 B.n121 585
R383 B.n121 B.n120 585
R384 B.n479 B.n478 585
R385 B.n480 B.n479 585
R386 B.n3 B.n0 585
R387 B.n4 B.n3 585
R388 B.n741 B.n1 585
R389 B.n742 B.n741 585
R390 B.n740 B.n739 585
R391 B.n740 B.n8 585
R392 B.n738 B.n9 585
R393 B.n12 B.n9 585
R394 B.n737 B.n736 585
R395 B.n736 B.n735 585
R396 B.n11 B.n10 585
R397 B.n734 B.n11 585
R398 B.n732 B.n731 585
R399 B.n733 B.n732 585
R400 B.n730 B.n17 585
R401 B.n17 B.n16 585
R402 B.n729 B.n728 585
R403 B.n728 B.n727 585
R404 B.n19 B.n18 585
R405 B.n726 B.n19 585
R406 B.n724 B.n723 585
R407 B.n725 B.n724 585
R408 B.n722 B.n23 585
R409 B.n26 B.n23 585
R410 B.n721 B.n720 585
R411 B.n720 B.n719 585
R412 B.n25 B.n24 585
R413 B.n718 B.n25 585
R414 B.n716 B.n715 585
R415 B.n717 B.n716 585
R416 B.n714 B.n31 585
R417 B.n31 B.n30 585
R418 B.n713 B.n712 585
R419 B.n712 B.n711 585
R420 B.n33 B.n32 585
R421 B.n710 B.n33 585
R422 B.n708 B.n707 585
R423 B.n709 B.n708 585
R424 B.n706 B.n38 585
R425 B.n38 B.n37 585
R426 B.n705 B.n704 585
R427 B.n704 B.n703 585
R428 B.n40 B.n39 585
R429 B.n702 B.n40 585
R430 B.n700 B.n699 585
R431 B.n701 B.n700 585
R432 B.n698 B.n45 585
R433 B.n45 B.n44 585
R434 B.n697 B.n696 585
R435 B.n696 B.n695 585
R436 B.n47 B.n46 585
R437 B.n694 B.n47 585
R438 B.n692 B.n691 585
R439 B.n693 B.n692 585
R440 B.n690 B.n52 585
R441 B.n52 B.n51 585
R442 B.n689 B.n688 585
R443 B.n688 B.n687 585
R444 B.n54 B.n53 585
R445 B.n686 B.n54 585
R446 B.n684 B.n683 585
R447 B.n685 B.n684 585
R448 B.n682 B.n59 585
R449 B.n59 B.n58 585
R450 B.n681 B.n680 585
R451 B.n680 B.n679 585
R452 B.n61 B.n60 585
R453 B.n678 B.n61 585
R454 B.n676 B.n675 585
R455 B.n677 B.n676 585
R456 B.n674 B.n66 585
R457 B.n66 B.n65 585
R458 B.n673 B.n672 585
R459 B.n672 B.n671 585
R460 B.n68 B.n67 585
R461 B.n670 B.n68 585
R462 B.n668 B.n667 585
R463 B.n669 B.n668 585
R464 B.n666 B.n73 585
R465 B.n73 B.n72 585
R466 B.n665 B.n664 585
R467 B.n664 B.n663 585
R468 B.n75 B.n74 585
R469 B.n662 B.n75 585
R470 B.n660 B.n659 585
R471 B.n661 B.n660 585
R472 B.n658 B.n80 585
R473 B.n80 B.n79 585
R474 B.n657 B.n656 585
R475 B.n656 B.n655 585
R476 B.n82 B.n81 585
R477 B.n654 B.n82 585
R478 B.n652 B.n651 585
R479 B.n653 B.n652 585
R480 B.n745 B.n744 585
R481 B.n743 B.n2 585
R482 B.n652 B.n87 473.281
R483 B.n545 B.n85 473.281
R484 B.n347 B.n206 473.281
R485 B.n345 B.n208 473.281
R486 B.n98 B.t10 274.755
R487 B.n106 B.t21 274.755
R488 B.n228 B.t14 274.755
R489 B.n221 B.t18 274.755
R490 B.n546 B.n86 256.663
R491 B.n552 B.n86 256.663
R492 B.n554 B.n86 256.663
R493 B.n560 B.n86 256.663
R494 B.n562 B.n86 256.663
R495 B.n568 B.n86 256.663
R496 B.n570 B.n86 256.663
R497 B.n576 B.n86 256.663
R498 B.n578 B.n86 256.663
R499 B.n584 B.n86 256.663
R500 B.n586 B.n86 256.663
R501 B.n593 B.n86 256.663
R502 B.n595 B.n86 256.663
R503 B.n601 B.n86 256.663
R504 B.n101 B.n86 256.663
R505 B.n607 B.n86 256.663
R506 B.n613 B.n86 256.663
R507 B.n615 B.n86 256.663
R508 B.n621 B.n86 256.663
R509 B.n623 B.n86 256.663
R510 B.n629 B.n86 256.663
R511 B.n631 B.n86 256.663
R512 B.n637 B.n86 256.663
R513 B.n639 B.n86 256.663
R514 B.n645 B.n86 256.663
R515 B.n647 B.n86 256.663
R516 B.n340 B.n207 256.663
R517 B.n210 B.n207 256.663
R518 B.n333 B.n207 256.663
R519 B.n327 B.n207 256.663
R520 B.n325 B.n207 256.663
R521 B.n319 B.n207 256.663
R522 B.n317 B.n207 256.663
R523 B.n311 B.n207 256.663
R524 B.n309 B.n207 256.663
R525 B.n303 B.n207 256.663
R526 B.n301 B.n207 256.663
R527 B.n295 B.n207 256.663
R528 B.n293 B.n207 256.663
R529 B.n287 B.n207 256.663
R530 B.n285 B.n207 256.663
R531 B.n278 B.n207 256.663
R532 B.n276 B.n207 256.663
R533 B.n270 B.n207 256.663
R534 B.n268 B.n207 256.663
R535 B.n262 B.n207 256.663
R536 B.n260 B.n207 256.663
R537 B.n254 B.n207 256.663
R538 B.n252 B.n207 256.663
R539 B.n246 B.n207 256.663
R540 B.n244 B.n207 256.663
R541 B.n239 B.n207 256.663
R542 B.n747 B.n746 256.663
R543 B.n106 B.t22 207.302
R544 B.n228 B.t17 207.302
R545 B.n98 B.t12 207.302
R546 B.n221 B.t20 207.302
R547 B.n107 B.t23 165.216
R548 B.n229 B.t16 165.216
R549 B.n99 B.t13 165.216
R550 B.n222 B.t19 165.216
R551 B.n648 B.n646 163.367
R552 B.n644 B.n89 163.367
R553 B.n640 B.n638 163.367
R554 B.n636 B.n91 163.367
R555 B.n632 B.n630 163.367
R556 B.n628 B.n93 163.367
R557 B.n624 B.n622 163.367
R558 B.n620 B.n95 163.367
R559 B.n616 B.n614 163.367
R560 B.n612 B.n97 163.367
R561 B.n608 B.n606 163.367
R562 B.n603 B.n602 163.367
R563 B.n600 B.n103 163.367
R564 B.n596 B.n594 163.367
R565 B.n592 B.n105 163.367
R566 B.n587 B.n585 163.367
R567 B.n583 B.n109 163.367
R568 B.n579 B.n577 163.367
R569 B.n575 B.n111 163.367
R570 B.n571 B.n569 163.367
R571 B.n567 B.n113 163.367
R572 B.n563 B.n561 163.367
R573 B.n559 B.n115 163.367
R574 B.n555 B.n553 163.367
R575 B.n551 B.n117 163.367
R576 B.n547 B.n545 163.367
R577 B.n347 B.n204 163.367
R578 B.n351 B.n204 163.367
R579 B.n351 B.n198 163.367
R580 B.n359 B.n198 163.367
R581 B.n359 B.n196 163.367
R582 B.n363 B.n196 163.367
R583 B.n363 B.n190 163.367
R584 B.n371 B.n190 163.367
R585 B.n371 B.n188 163.367
R586 B.n375 B.n188 163.367
R587 B.n375 B.n182 163.367
R588 B.n383 B.n182 163.367
R589 B.n383 B.n180 163.367
R590 B.n387 B.n180 163.367
R591 B.n387 B.n174 163.367
R592 B.n395 B.n174 163.367
R593 B.n395 B.n172 163.367
R594 B.n399 B.n172 163.367
R595 B.n399 B.n166 163.367
R596 B.n407 B.n166 163.367
R597 B.n407 B.n164 163.367
R598 B.n411 B.n164 163.367
R599 B.n411 B.n158 163.367
R600 B.n419 B.n158 163.367
R601 B.n419 B.n156 163.367
R602 B.n423 B.n156 163.367
R603 B.n423 B.n150 163.367
R604 B.n431 B.n150 163.367
R605 B.n431 B.n148 163.367
R606 B.n435 B.n148 163.367
R607 B.n435 B.n142 163.367
R608 B.n443 B.n142 163.367
R609 B.n443 B.n140 163.367
R610 B.n447 B.n140 163.367
R611 B.n447 B.n135 163.367
R612 B.n456 B.n135 163.367
R613 B.n456 B.n133 163.367
R614 B.n460 B.n133 163.367
R615 B.n460 B.n126 163.367
R616 B.n468 B.n126 163.367
R617 B.n468 B.n124 163.367
R618 B.n473 B.n124 163.367
R619 B.n473 B.n119 163.367
R620 B.n481 B.n119 163.367
R621 B.n482 B.n481 163.367
R622 B.n482 B.n5 163.367
R623 B.n6 B.n5 163.367
R624 B.n7 B.n6 163.367
R625 B.n488 B.n7 163.367
R626 B.n489 B.n488 163.367
R627 B.n489 B.n13 163.367
R628 B.n14 B.n13 163.367
R629 B.n15 B.n14 163.367
R630 B.n494 B.n15 163.367
R631 B.n494 B.n20 163.367
R632 B.n21 B.n20 163.367
R633 B.n22 B.n21 163.367
R634 B.n499 B.n22 163.367
R635 B.n499 B.n27 163.367
R636 B.n28 B.n27 163.367
R637 B.n29 B.n28 163.367
R638 B.n504 B.n29 163.367
R639 B.n504 B.n34 163.367
R640 B.n35 B.n34 163.367
R641 B.n36 B.n35 163.367
R642 B.n509 B.n36 163.367
R643 B.n509 B.n41 163.367
R644 B.n42 B.n41 163.367
R645 B.n43 B.n42 163.367
R646 B.n514 B.n43 163.367
R647 B.n514 B.n48 163.367
R648 B.n49 B.n48 163.367
R649 B.n50 B.n49 163.367
R650 B.n519 B.n50 163.367
R651 B.n519 B.n55 163.367
R652 B.n56 B.n55 163.367
R653 B.n57 B.n56 163.367
R654 B.n524 B.n57 163.367
R655 B.n524 B.n62 163.367
R656 B.n63 B.n62 163.367
R657 B.n64 B.n63 163.367
R658 B.n529 B.n64 163.367
R659 B.n529 B.n69 163.367
R660 B.n70 B.n69 163.367
R661 B.n71 B.n70 163.367
R662 B.n534 B.n71 163.367
R663 B.n534 B.n76 163.367
R664 B.n77 B.n76 163.367
R665 B.n78 B.n77 163.367
R666 B.n539 B.n78 163.367
R667 B.n539 B.n83 163.367
R668 B.n84 B.n83 163.367
R669 B.n85 B.n84 163.367
R670 B.n341 B.n339 163.367
R671 B.n339 B.n338 163.367
R672 B.n335 B.n334 163.367
R673 B.n332 B.n212 163.367
R674 B.n328 B.n326 163.367
R675 B.n324 B.n214 163.367
R676 B.n320 B.n318 163.367
R677 B.n316 B.n216 163.367
R678 B.n312 B.n310 163.367
R679 B.n308 B.n218 163.367
R680 B.n304 B.n302 163.367
R681 B.n300 B.n220 163.367
R682 B.n296 B.n294 163.367
R683 B.n292 B.n225 163.367
R684 B.n288 B.n286 163.367
R685 B.n284 B.n227 163.367
R686 B.n279 B.n277 163.367
R687 B.n275 B.n231 163.367
R688 B.n271 B.n269 163.367
R689 B.n267 B.n233 163.367
R690 B.n263 B.n261 163.367
R691 B.n259 B.n235 163.367
R692 B.n255 B.n253 163.367
R693 B.n251 B.n237 163.367
R694 B.n247 B.n245 163.367
R695 B.n243 B.n240 163.367
R696 B.n345 B.n202 163.367
R697 B.n353 B.n202 163.367
R698 B.n353 B.n200 163.367
R699 B.n357 B.n200 163.367
R700 B.n357 B.n194 163.367
R701 B.n365 B.n194 163.367
R702 B.n365 B.n192 163.367
R703 B.n369 B.n192 163.367
R704 B.n369 B.n186 163.367
R705 B.n377 B.n186 163.367
R706 B.n377 B.n184 163.367
R707 B.n381 B.n184 163.367
R708 B.n381 B.n178 163.367
R709 B.n389 B.n178 163.367
R710 B.n389 B.n176 163.367
R711 B.n393 B.n176 163.367
R712 B.n393 B.n170 163.367
R713 B.n401 B.n170 163.367
R714 B.n401 B.n168 163.367
R715 B.n405 B.n168 163.367
R716 B.n405 B.n162 163.367
R717 B.n413 B.n162 163.367
R718 B.n413 B.n160 163.367
R719 B.n417 B.n160 163.367
R720 B.n417 B.n154 163.367
R721 B.n425 B.n154 163.367
R722 B.n425 B.n152 163.367
R723 B.n429 B.n152 163.367
R724 B.n429 B.n146 163.367
R725 B.n437 B.n146 163.367
R726 B.n437 B.n144 163.367
R727 B.n441 B.n144 163.367
R728 B.n441 B.n138 163.367
R729 B.n450 B.n138 163.367
R730 B.n450 B.n136 163.367
R731 B.n454 B.n136 163.367
R732 B.n454 B.n131 163.367
R733 B.n462 B.n131 163.367
R734 B.n462 B.n129 163.367
R735 B.n466 B.n129 163.367
R736 B.n466 B.n123 163.367
R737 B.n475 B.n123 163.367
R738 B.n475 B.n121 163.367
R739 B.n479 B.n121 163.367
R740 B.n479 B.n3 163.367
R741 B.n745 B.n3 163.367
R742 B.n741 B.n2 163.367
R743 B.n741 B.n740 163.367
R744 B.n740 B.n9 163.367
R745 B.n736 B.n9 163.367
R746 B.n736 B.n11 163.367
R747 B.n732 B.n11 163.367
R748 B.n732 B.n17 163.367
R749 B.n728 B.n17 163.367
R750 B.n728 B.n19 163.367
R751 B.n724 B.n19 163.367
R752 B.n724 B.n23 163.367
R753 B.n720 B.n23 163.367
R754 B.n720 B.n25 163.367
R755 B.n716 B.n25 163.367
R756 B.n716 B.n31 163.367
R757 B.n712 B.n31 163.367
R758 B.n712 B.n33 163.367
R759 B.n708 B.n33 163.367
R760 B.n708 B.n38 163.367
R761 B.n704 B.n38 163.367
R762 B.n704 B.n40 163.367
R763 B.n700 B.n40 163.367
R764 B.n700 B.n45 163.367
R765 B.n696 B.n45 163.367
R766 B.n696 B.n47 163.367
R767 B.n692 B.n47 163.367
R768 B.n692 B.n52 163.367
R769 B.n688 B.n52 163.367
R770 B.n688 B.n54 163.367
R771 B.n684 B.n54 163.367
R772 B.n684 B.n59 163.367
R773 B.n680 B.n59 163.367
R774 B.n680 B.n61 163.367
R775 B.n676 B.n61 163.367
R776 B.n676 B.n66 163.367
R777 B.n672 B.n66 163.367
R778 B.n672 B.n68 163.367
R779 B.n668 B.n68 163.367
R780 B.n668 B.n73 163.367
R781 B.n664 B.n73 163.367
R782 B.n664 B.n75 163.367
R783 B.n660 B.n75 163.367
R784 B.n660 B.n80 163.367
R785 B.n656 B.n80 163.367
R786 B.n656 B.n82 163.367
R787 B.n652 B.n82 163.367
R788 B.n346 B.n207 122.748
R789 B.n653 B.n86 122.748
R790 B.n647 B.n87 71.676
R791 B.n646 B.n645 71.676
R792 B.n639 B.n89 71.676
R793 B.n638 B.n637 71.676
R794 B.n631 B.n91 71.676
R795 B.n630 B.n629 71.676
R796 B.n623 B.n93 71.676
R797 B.n622 B.n621 71.676
R798 B.n615 B.n95 71.676
R799 B.n614 B.n613 71.676
R800 B.n607 B.n97 71.676
R801 B.n606 B.n101 71.676
R802 B.n602 B.n601 71.676
R803 B.n595 B.n103 71.676
R804 B.n594 B.n593 71.676
R805 B.n586 B.n105 71.676
R806 B.n585 B.n584 71.676
R807 B.n578 B.n109 71.676
R808 B.n577 B.n576 71.676
R809 B.n570 B.n111 71.676
R810 B.n569 B.n568 71.676
R811 B.n562 B.n113 71.676
R812 B.n561 B.n560 71.676
R813 B.n554 B.n115 71.676
R814 B.n553 B.n552 71.676
R815 B.n546 B.n117 71.676
R816 B.n547 B.n546 71.676
R817 B.n552 B.n551 71.676
R818 B.n555 B.n554 71.676
R819 B.n560 B.n559 71.676
R820 B.n563 B.n562 71.676
R821 B.n568 B.n567 71.676
R822 B.n571 B.n570 71.676
R823 B.n576 B.n575 71.676
R824 B.n579 B.n578 71.676
R825 B.n584 B.n583 71.676
R826 B.n587 B.n586 71.676
R827 B.n593 B.n592 71.676
R828 B.n596 B.n595 71.676
R829 B.n601 B.n600 71.676
R830 B.n603 B.n101 71.676
R831 B.n608 B.n607 71.676
R832 B.n613 B.n612 71.676
R833 B.n616 B.n615 71.676
R834 B.n621 B.n620 71.676
R835 B.n624 B.n623 71.676
R836 B.n629 B.n628 71.676
R837 B.n632 B.n631 71.676
R838 B.n637 B.n636 71.676
R839 B.n640 B.n639 71.676
R840 B.n645 B.n644 71.676
R841 B.n648 B.n647 71.676
R842 B.n340 B.n208 71.676
R843 B.n338 B.n210 71.676
R844 B.n334 B.n333 71.676
R845 B.n327 B.n212 71.676
R846 B.n326 B.n325 71.676
R847 B.n319 B.n214 71.676
R848 B.n318 B.n317 71.676
R849 B.n311 B.n216 71.676
R850 B.n310 B.n309 71.676
R851 B.n303 B.n218 71.676
R852 B.n302 B.n301 71.676
R853 B.n295 B.n220 71.676
R854 B.n294 B.n293 71.676
R855 B.n287 B.n225 71.676
R856 B.n286 B.n285 71.676
R857 B.n278 B.n227 71.676
R858 B.n277 B.n276 71.676
R859 B.n270 B.n231 71.676
R860 B.n269 B.n268 71.676
R861 B.n262 B.n233 71.676
R862 B.n261 B.n260 71.676
R863 B.n254 B.n235 71.676
R864 B.n253 B.n252 71.676
R865 B.n246 B.n237 71.676
R866 B.n245 B.n244 71.676
R867 B.n240 B.n239 71.676
R868 B.n341 B.n340 71.676
R869 B.n335 B.n210 71.676
R870 B.n333 B.n332 71.676
R871 B.n328 B.n327 71.676
R872 B.n325 B.n324 71.676
R873 B.n320 B.n319 71.676
R874 B.n317 B.n316 71.676
R875 B.n312 B.n311 71.676
R876 B.n309 B.n308 71.676
R877 B.n304 B.n303 71.676
R878 B.n301 B.n300 71.676
R879 B.n296 B.n295 71.676
R880 B.n293 B.n292 71.676
R881 B.n288 B.n287 71.676
R882 B.n285 B.n284 71.676
R883 B.n279 B.n278 71.676
R884 B.n276 B.n275 71.676
R885 B.n271 B.n270 71.676
R886 B.n268 B.n267 71.676
R887 B.n263 B.n262 71.676
R888 B.n260 B.n259 71.676
R889 B.n255 B.n254 71.676
R890 B.n252 B.n251 71.676
R891 B.n247 B.n246 71.676
R892 B.n244 B.n243 71.676
R893 B.n239 B.n206 71.676
R894 B.n746 B.n745 71.676
R895 B.n746 B.n2 71.676
R896 B.n346 B.n203 71.3405
R897 B.n352 B.n203 71.3405
R898 B.n352 B.n199 71.3405
R899 B.n358 B.n199 71.3405
R900 B.n358 B.n195 71.3405
R901 B.n364 B.n195 71.3405
R902 B.n370 B.n191 71.3405
R903 B.n370 B.n187 71.3405
R904 B.n376 B.n187 71.3405
R905 B.n376 B.n183 71.3405
R906 B.n382 B.n183 71.3405
R907 B.n382 B.n179 71.3405
R908 B.n388 B.n179 71.3405
R909 B.n388 B.n175 71.3405
R910 B.n394 B.n175 71.3405
R911 B.n400 B.n171 71.3405
R912 B.n400 B.n167 71.3405
R913 B.n406 B.n167 71.3405
R914 B.n406 B.n163 71.3405
R915 B.n412 B.n163 71.3405
R916 B.n418 B.n159 71.3405
R917 B.n418 B.n155 71.3405
R918 B.n424 B.n155 71.3405
R919 B.n424 B.n151 71.3405
R920 B.n430 B.n151 71.3405
R921 B.n436 B.n147 71.3405
R922 B.n436 B.n143 71.3405
R923 B.n442 B.n143 71.3405
R924 B.n442 B.n139 71.3405
R925 B.n449 B.n139 71.3405
R926 B.n449 B.n448 71.3405
R927 B.n455 B.n132 71.3405
R928 B.n461 B.n132 71.3405
R929 B.n461 B.n127 71.3405
R930 B.n467 B.n127 71.3405
R931 B.n467 B.n128 71.3405
R932 B.n474 B.n120 71.3405
R933 B.n480 B.n120 71.3405
R934 B.n480 B.n4 71.3405
R935 B.n744 B.n4 71.3405
R936 B.n744 B.n743 71.3405
R937 B.n743 B.n742 71.3405
R938 B.n742 B.n8 71.3405
R939 B.n12 B.n8 71.3405
R940 B.n735 B.n12 71.3405
R941 B.n734 B.n733 71.3405
R942 B.n733 B.n16 71.3405
R943 B.n727 B.n16 71.3405
R944 B.n727 B.n726 71.3405
R945 B.n726 B.n725 71.3405
R946 B.n719 B.n26 71.3405
R947 B.n719 B.n718 71.3405
R948 B.n718 B.n717 71.3405
R949 B.n717 B.n30 71.3405
R950 B.n711 B.n30 71.3405
R951 B.n711 B.n710 71.3405
R952 B.n709 B.n37 71.3405
R953 B.n703 B.n37 71.3405
R954 B.n703 B.n702 71.3405
R955 B.n702 B.n701 71.3405
R956 B.n701 B.n44 71.3405
R957 B.n695 B.n694 71.3405
R958 B.n694 B.n693 71.3405
R959 B.n693 B.n51 71.3405
R960 B.n687 B.n51 71.3405
R961 B.n687 B.n686 71.3405
R962 B.n685 B.n58 71.3405
R963 B.n679 B.n58 71.3405
R964 B.n679 B.n678 71.3405
R965 B.n678 B.n677 71.3405
R966 B.n677 B.n65 71.3405
R967 B.n671 B.n65 71.3405
R968 B.n671 B.n670 71.3405
R969 B.n670 B.n669 71.3405
R970 B.n669 B.n72 71.3405
R971 B.n663 B.n662 71.3405
R972 B.n662 B.n661 71.3405
R973 B.n661 B.n79 71.3405
R974 B.n655 B.n79 71.3405
R975 B.n655 B.n654 71.3405
R976 B.n654 B.n653 71.3405
R977 B.n430 B.t0 67.144
R978 B.t3 B.n709 67.144
R979 B.n100 B.n99 59.5399
R980 B.n589 B.n107 59.5399
R981 B.n282 B.n229 59.5399
R982 B.n223 B.n222 59.5399
R983 B.t7 B.n171 58.7511
R984 B.n686 B.t1 58.7511
R985 B.n128 B.t6 50.3582
R986 B.t5 B.n734 50.3582
R987 B.n455 B.t4 48.2599
R988 B.n725 B.t2 48.2599
R989 B.n99 B.n98 42.0853
R990 B.n107 B.n106 42.0853
R991 B.n229 B.n228 42.0853
R992 B.n222 B.n221 42.0853
R993 B.n364 B.t15 41.9652
R994 B.n663 B.t11 41.9652
R995 B.n412 B.t9 39.867
R996 B.n695 B.t8 39.867
R997 B.t9 B.n159 31.474
R998 B.t8 B.n44 31.474
R999 B.n344 B.n343 30.7517
R1000 B.n348 B.n205 30.7517
R1001 B.n544 B.n543 30.7517
R1002 B.n651 B.n650 30.7517
R1003 B.t15 B.n191 29.3758
R1004 B.t11 B.n72 29.3758
R1005 B.n448 B.t4 23.0811
R1006 B.n26 B.t2 23.0811
R1007 B.n474 B.t6 20.9829
R1008 B.n735 B.t5 20.9829
R1009 B B.n747 18.0485
R1010 B.n394 B.t7 12.5899
R1011 B.t1 B.n685 12.5899
R1012 B.n344 B.n201 10.6151
R1013 B.n354 B.n201 10.6151
R1014 B.n355 B.n354 10.6151
R1015 B.n356 B.n355 10.6151
R1016 B.n356 B.n193 10.6151
R1017 B.n366 B.n193 10.6151
R1018 B.n367 B.n366 10.6151
R1019 B.n368 B.n367 10.6151
R1020 B.n368 B.n185 10.6151
R1021 B.n378 B.n185 10.6151
R1022 B.n379 B.n378 10.6151
R1023 B.n380 B.n379 10.6151
R1024 B.n380 B.n177 10.6151
R1025 B.n390 B.n177 10.6151
R1026 B.n391 B.n390 10.6151
R1027 B.n392 B.n391 10.6151
R1028 B.n392 B.n169 10.6151
R1029 B.n402 B.n169 10.6151
R1030 B.n403 B.n402 10.6151
R1031 B.n404 B.n403 10.6151
R1032 B.n404 B.n161 10.6151
R1033 B.n414 B.n161 10.6151
R1034 B.n415 B.n414 10.6151
R1035 B.n416 B.n415 10.6151
R1036 B.n416 B.n153 10.6151
R1037 B.n426 B.n153 10.6151
R1038 B.n427 B.n426 10.6151
R1039 B.n428 B.n427 10.6151
R1040 B.n428 B.n145 10.6151
R1041 B.n438 B.n145 10.6151
R1042 B.n439 B.n438 10.6151
R1043 B.n440 B.n439 10.6151
R1044 B.n440 B.n137 10.6151
R1045 B.n451 B.n137 10.6151
R1046 B.n452 B.n451 10.6151
R1047 B.n453 B.n452 10.6151
R1048 B.n453 B.n130 10.6151
R1049 B.n463 B.n130 10.6151
R1050 B.n464 B.n463 10.6151
R1051 B.n465 B.n464 10.6151
R1052 B.n465 B.n122 10.6151
R1053 B.n476 B.n122 10.6151
R1054 B.n477 B.n476 10.6151
R1055 B.n478 B.n477 10.6151
R1056 B.n478 B.n0 10.6151
R1057 B.n343 B.n342 10.6151
R1058 B.n342 B.n209 10.6151
R1059 B.n337 B.n209 10.6151
R1060 B.n337 B.n336 10.6151
R1061 B.n336 B.n211 10.6151
R1062 B.n331 B.n211 10.6151
R1063 B.n331 B.n330 10.6151
R1064 B.n330 B.n329 10.6151
R1065 B.n329 B.n213 10.6151
R1066 B.n323 B.n213 10.6151
R1067 B.n323 B.n322 10.6151
R1068 B.n322 B.n321 10.6151
R1069 B.n321 B.n215 10.6151
R1070 B.n315 B.n215 10.6151
R1071 B.n315 B.n314 10.6151
R1072 B.n314 B.n313 10.6151
R1073 B.n313 B.n217 10.6151
R1074 B.n307 B.n217 10.6151
R1075 B.n307 B.n306 10.6151
R1076 B.n306 B.n305 10.6151
R1077 B.n305 B.n219 10.6151
R1078 B.n299 B.n298 10.6151
R1079 B.n298 B.n297 10.6151
R1080 B.n297 B.n224 10.6151
R1081 B.n291 B.n224 10.6151
R1082 B.n291 B.n290 10.6151
R1083 B.n290 B.n289 10.6151
R1084 B.n289 B.n226 10.6151
R1085 B.n283 B.n226 10.6151
R1086 B.n281 B.n280 10.6151
R1087 B.n280 B.n230 10.6151
R1088 B.n274 B.n230 10.6151
R1089 B.n274 B.n273 10.6151
R1090 B.n273 B.n272 10.6151
R1091 B.n272 B.n232 10.6151
R1092 B.n266 B.n232 10.6151
R1093 B.n266 B.n265 10.6151
R1094 B.n265 B.n264 10.6151
R1095 B.n264 B.n234 10.6151
R1096 B.n258 B.n234 10.6151
R1097 B.n258 B.n257 10.6151
R1098 B.n257 B.n256 10.6151
R1099 B.n256 B.n236 10.6151
R1100 B.n250 B.n236 10.6151
R1101 B.n250 B.n249 10.6151
R1102 B.n249 B.n248 10.6151
R1103 B.n248 B.n238 10.6151
R1104 B.n242 B.n238 10.6151
R1105 B.n242 B.n241 10.6151
R1106 B.n241 B.n205 10.6151
R1107 B.n349 B.n348 10.6151
R1108 B.n350 B.n349 10.6151
R1109 B.n350 B.n197 10.6151
R1110 B.n360 B.n197 10.6151
R1111 B.n361 B.n360 10.6151
R1112 B.n362 B.n361 10.6151
R1113 B.n362 B.n189 10.6151
R1114 B.n372 B.n189 10.6151
R1115 B.n373 B.n372 10.6151
R1116 B.n374 B.n373 10.6151
R1117 B.n374 B.n181 10.6151
R1118 B.n384 B.n181 10.6151
R1119 B.n385 B.n384 10.6151
R1120 B.n386 B.n385 10.6151
R1121 B.n386 B.n173 10.6151
R1122 B.n396 B.n173 10.6151
R1123 B.n397 B.n396 10.6151
R1124 B.n398 B.n397 10.6151
R1125 B.n398 B.n165 10.6151
R1126 B.n408 B.n165 10.6151
R1127 B.n409 B.n408 10.6151
R1128 B.n410 B.n409 10.6151
R1129 B.n410 B.n157 10.6151
R1130 B.n420 B.n157 10.6151
R1131 B.n421 B.n420 10.6151
R1132 B.n422 B.n421 10.6151
R1133 B.n422 B.n149 10.6151
R1134 B.n432 B.n149 10.6151
R1135 B.n433 B.n432 10.6151
R1136 B.n434 B.n433 10.6151
R1137 B.n434 B.n141 10.6151
R1138 B.n444 B.n141 10.6151
R1139 B.n445 B.n444 10.6151
R1140 B.n446 B.n445 10.6151
R1141 B.n446 B.n134 10.6151
R1142 B.n457 B.n134 10.6151
R1143 B.n458 B.n457 10.6151
R1144 B.n459 B.n458 10.6151
R1145 B.n459 B.n125 10.6151
R1146 B.n469 B.n125 10.6151
R1147 B.n470 B.n469 10.6151
R1148 B.n472 B.n470 10.6151
R1149 B.n472 B.n471 10.6151
R1150 B.n471 B.n118 10.6151
R1151 B.n483 B.n118 10.6151
R1152 B.n484 B.n483 10.6151
R1153 B.n485 B.n484 10.6151
R1154 B.n486 B.n485 10.6151
R1155 B.n487 B.n486 10.6151
R1156 B.n490 B.n487 10.6151
R1157 B.n491 B.n490 10.6151
R1158 B.n492 B.n491 10.6151
R1159 B.n493 B.n492 10.6151
R1160 B.n495 B.n493 10.6151
R1161 B.n496 B.n495 10.6151
R1162 B.n497 B.n496 10.6151
R1163 B.n498 B.n497 10.6151
R1164 B.n500 B.n498 10.6151
R1165 B.n501 B.n500 10.6151
R1166 B.n502 B.n501 10.6151
R1167 B.n503 B.n502 10.6151
R1168 B.n505 B.n503 10.6151
R1169 B.n506 B.n505 10.6151
R1170 B.n507 B.n506 10.6151
R1171 B.n508 B.n507 10.6151
R1172 B.n510 B.n508 10.6151
R1173 B.n511 B.n510 10.6151
R1174 B.n512 B.n511 10.6151
R1175 B.n513 B.n512 10.6151
R1176 B.n515 B.n513 10.6151
R1177 B.n516 B.n515 10.6151
R1178 B.n517 B.n516 10.6151
R1179 B.n518 B.n517 10.6151
R1180 B.n520 B.n518 10.6151
R1181 B.n521 B.n520 10.6151
R1182 B.n522 B.n521 10.6151
R1183 B.n523 B.n522 10.6151
R1184 B.n525 B.n523 10.6151
R1185 B.n526 B.n525 10.6151
R1186 B.n527 B.n526 10.6151
R1187 B.n528 B.n527 10.6151
R1188 B.n530 B.n528 10.6151
R1189 B.n531 B.n530 10.6151
R1190 B.n532 B.n531 10.6151
R1191 B.n533 B.n532 10.6151
R1192 B.n535 B.n533 10.6151
R1193 B.n536 B.n535 10.6151
R1194 B.n537 B.n536 10.6151
R1195 B.n538 B.n537 10.6151
R1196 B.n540 B.n538 10.6151
R1197 B.n541 B.n540 10.6151
R1198 B.n542 B.n541 10.6151
R1199 B.n543 B.n542 10.6151
R1200 B.n739 B.n1 10.6151
R1201 B.n739 B.n738 10.6151
R1202 B.n738 B.n737 10.6151
R1203 B.n737 B.n10 10.6151
R1204 B.n731 B.n10 10.6151
R1205 B.n731 B.n730 10.6151
R1206 B.n730 B.n729 10.6151
R1207 B.n729 B.n18 10.6151
R1208 B.n723 B.n18 10.6151
R1209 B.n723 B.n722 10.6151
R1210 B.n722 B.n721 10.6151
R1211 B.n721 B.n24 10.6151
R1212 B.n715 B.n24 10.6151
R1213 B.n715 B.n714 10.6151
R1214 B.n714 B.n713 10.6151
R1215 B.n713 B.n32 10.6151
R1216 B.n707 B.n32 10.6151
R1217 B.n707 B.n706 10.6151
R1218 B.n706 B.n705 10.6151
R1219 B.n705 B.n39 10.6151
R1220 B.n699 B.n39 10.6151
R1221 B.n699 B.n698 10.6151
R1222 B.n698 B.n697 10.6151
R1223 B.n697 B.n46 10.6151
R1224 B.n691 B.n46 10.6151
R1225 B.n691 B.n690 10.6151
R1226 B.n690 B.n689 10.6151
R1227 B.n689 B.n53 10.6151
R1228 B.n683 B.n53 10.6151
R1229 B.n683 B.n682 10.6151
R1230 B.n682 B.n681 10.6151
R1231 B.n681 B.n60 10.6151
R1232 B.n675 B.n60 10.6151
R1233 B.n675 B.n674 10.6151
R1234 B.n674 B.n673 10.6151
R1235 B.n673 B.n67 10.6151
R1236 B.n667 B.n67 10.6151
R1237 B.n667 B.n666 10.6151
R1238 B.n666 B.n665 10.6151
R1239 B.n665 B.n74 10.6151
R1240 B.n659 B.n74 10.6151
R1241 B.n659 B.n658 10.6151
R1242 B.n658 B.n657 10.6151
R1243 B.n657 B.n81 10.6151
R1244 B.n651 B.n81 10.6151
R1245 B.n650 B.n649 10.6151
R1246 B.n649 B.n88 10.6151
R1247 B.n643 B.n88 10.6151
R1248 B.n643 B.n642 10.6151
R1249 B.n642 B.n641 10.6151
R1250 B.n641 B.n90 10.6151
R1251 B.n635 B.n90 10.6151
R1252 B.n635 B.n634 10.6151
R1253 B.n634 B.n633 10.6151
R1254 B.n633 B.n92 10.6151
R1255 B.n627 B.n92 10.6151
R1256 B.n627 B.n626 10.6151
R1257 B.n626 B.n625 10.6151
R1258 B.n625 B.n94 10.6151
R1259 B.n619 B.n94 10.6151
R1260 B.n619 B.n618 10.6151
R1261 B.n618 B.n617 10.6151
R1262 B.n617 B.n96 10.6151
R1263 B.n611 B.n96 10.6151
R1264 B.n611 B.n610 10.6151
R1265 B.n610 B.n609 10.6151
R1266 B.n605 B.n604 10.6151
R1267 B.n604 B.n102 10.6151
R1268 B.n599 B.n102 10.6151
R1269 B.n599 B.n598 10.6151
R1270 B.n598 B.n597 10.6151
R1271 B.n597 B.n104 10.6151
R1272 B.n591 B.n104 10.6151
R1273 B.n591 B.n590 10.6151
R1274 B.n588 B.n108 10.6151
R1275 B.n582 B.n108 10.6151
R1276 B.n582 B.n581 10.6151
R1277 B.n581 B.n580 10.6151
R1278 B.n580 B.n110 10.6151
R1279 B.n574 B.n110 10.6151
R1280 B.n574 B.n573 10.6151
R1281 B.n573 B.n572 10.6151
R1282 B.n572 B.n112 10.6151
R1283 B.n566 B.n112 10.6151
R1284 B.n566 B.n565 10.6151
R1285 B.n565 B.n564 10.6151
R1286 B.n564 B.n114 10.6151
R1287 B.n558 B.n114 10.6151
R1288 B.n558 B.n557 10.6151
R1289 B.n557 B.n556 10.6151
R1290 B.n556 B.n116 10.6151
R1291 B.n550 B.n116 10.6151
R1292 B.n550 B.n549 10.6151
R1293 B.n549 B.n548 10.6151
R1294 B.n548 B.n544 10.6151
R1295 B.n747 B.n0 8.11757
R1296 B.n747 B.n1 8.11757
R1297 B.n299 B.n223 6.5566
R1298 B.n283 B.n282 6.5566
R1299 B.n605 B.n100 6.5566
R1300 B.n590 B.n589 6.5566
R1301 B.t0 B.n147 4.19697
R1302 B.n710 B.t3 4.19697
R1303 B.n223 B.n219 4.05904
R1304 B.n282 B.n281 4.05904
R1305 B.n609 B.n100 4.05904
R1306 B.n589 B.n588 4.05904
R1307 VP.n42 VP.n9 181.363
R1308 VP.n74 VP.n73 181.363
R1309 VP.n41 VP.n40 181.363
R1310 VP.n19 VP.n16 161.3
R1311 VP.n21 VP.n20 161.3
R1312 VP.n22 VP.n15 161.3
R1313 VP.n24 VP.n23 161.3
R1314 VP.n26 VP.n14 161.3
R1315 VP.n28 VP.n27 161.3
R1316 VP.n29 VP.n13 161.3
R1317 VP.n31 VP.n30 161.3
R1318 VP.n33 VP.n12 161.3
R1319 VP.n35 VP.n34 161.3
R1320 VP.n36 VP.n11 161.3
R1321 VP.n38 VP.n37 161.3
R1322 VP.n39 VP.n10 161.3
R1323 VP.n72 VP.n0 161.3
R1324 VP.n71 VP.n70 161.3
R1325 VP.n69 VP.n1 161.3
R1326 VP.n68 VP.n67 161.3
R1327 VP.n66 VP.n2 161.3
R1328 VP.n64 VP.n63 161.3
R1329 VP.n62 VP.n3 161.3
R1330 VP.n61 VP.n60 161.3
R1331 VP.n59 VP.n4 161.3
R1332 VP.n57 VP.n56 161.3
R1333 VP.n55 VP.n5 161.3
R1334 VP.n54 VP.n53 161.3
R1335 VP.n52 VP.n6 161.3
R1336 VP.n50 VP.n49 161.3
R1337 VP.n48 VP.n7 161.3
R1338 VP.n47 VP.n46 161.3
R1339 VP.n45 VP.n8 161.3
R1340 VP.n44 VP.n43 161.3
R1341 VP.n17 VP.t9 103.059
R1342 VP.n9 VP.t1 68.2402
R1343 VP.n51 VP.t5 68.2402
R1344 VP.n58 VP.t8 68.2402
R1345 VP.n65 VP.t0 68.2402
R1346 VP.n73 VP.t4 68.2402
R1347 VP.n40 VP.t7 68.2402
R1348 VP.n32 VP.t2 68.2402
R1349 VP.n25 VP.t3 68.2402
R1350 VP.n18 VP.t6 68.2402
R1351 VP.n53 VP.n5 56.5193
R1352 VP.n60 VP.n3 56.5193
R1353 VP.n27 VP.n13 56.5193
R1354 VP.n20 VP.n15 56.5193
R1355 VP.n18 VP.n17 48.825
R1356 VP.n42 VP.n41 43.7619
R1357 VP.n46 VP.n45 40.979
R1358 VP.n71 VP.n1 40.979
R1359 VP.n38 VP.n11 40.979
R1360 VP.n46 VP.n7 40.0078
R1361 VP.n67 VP.n1 40.0078
R1362 VP.n34 VP.n11 40.0078
R1363 VP.n45 VP.n44 24.4675
R1364 VP.n50 VP.n7 24.4675
R1365 VP.n53 VP.n52 24.4675
R1366 VP.n57 VP.n5 24.4675
R1367 VP.n60 VP.n59 24.4675
R1368 VP.n64 VP.n3 24.4675
R1369 VP.n67 VP.n66 24.4675
R1370 VP.n72 VP.n71 24.4675
R1371 VP.n39 VP.n38 24.4675
R1372 VP.n31 VP.n13 24.4675
R1373 VP.n34 VP.n33 24.4675
R1374 VP.n24 VP.n15 24.4675
R1375 VP.n27 VP.n26 24.4675
R1376 VP.n20 VP.n19 24.4675
R1377 VP.n52 VP.n51 20.5528
R1378 VP.n65 VP.n64 20.5528
R1379 VP.n32 VP.n31 20.5528
R1380 VP.n19 VP.n18 20.5528
R1381 VP.n17 VP.n16 12.2488
R1382 VP.n58 VP.n57 12.234
R1383 VP.n59 VP.n58 12.234
R1384 VP.n25 VP.n24 12.234
R1385 VP.n26 VP.n25 12.234
R1386 VP.n44 VP.n9 4.40456
R1387 VP.n73 VP.n72 4.40456
R1388 VP.n40 VP.n39 4.40456
R1389 VP.n51 VP.n50 3.91522
R1390 VP.n66 VP.n65 3.91522
R1391 VP.n33 VP.n32 3.91522
R1392 VP.n21 VP.n16 0.189894
R1393 VP.n22 VP.n21 0.189894
R1394 VP.n23 VP.n22 0.189894
R1395 VP.n23 VP.n14 0.189894
R1396 VP.n28 VP.n14 0.189894
R1397 VP.n29 VP.n28 0.189894
R1398 VP.n30 VP.n29 0.189894
R1399 VP.n30 VP.n12 0.189894
R1400 VP.n35 VP.n12 0.189894
R1401 VP.n36 VP.n35 0.189894
R1402 VP.n37 VP.n36 0.189894
R1403 VP.n37 VP.n10 0.189894
R1404 VP.n41 VP.n10 0.189894
R1405 VP.n43 VP.n42 0.189894
R1406 VP.n43 VP.n8 0.189894
R1407 VP.n47 VP.n8 0.189894
R1408 VP.n48 VP.n47 0.189894
R1409 VP.n49 VP.n48 0.189894
R1410 VP.n49 VP.n6 0.189894
R1411 VP.n54 VP.n6 0.189894
R1412 VP.n55 VP.n54 0.189894
R1413 VP.n56 VP.n55 0.189894
R1414 VP.n56 VP.n4 0.189894
R1415 VP.n61 VP.n4 0.189894
R1416 VP.n62 VP.n61 0.189894
R1417 VP.n63 VP.n62 0.189894
R1418 VP.n63 VP.n2 0.189894
R1419 VP.n68 VP.n2 0.189894
R1420 VP.n69 VP.n68 0.189894
R1421 VP.n70 VP.n69 0.189894
R1422 VP.n70 VP.n0 0.189894
R1423 VP.n74 VP.n0 0.189894
R1424 VP VP.n74 0.0516364
R1425 VDD1.n22 VDD1.n0 289.615
R1426 VDD1.n51 VDD1.n29 289.615
R1427 VDD1.n23 VDD1.n22 185
R1428 VDD1.n21 VDD1.n20 185
R1429 VDD1.n4 VDD1.n3 185
R1430 VDD1.n15 VDD1.n14 185
R1431 VDD1.n13 VDD1.n12 185
R1432 VDD1.n8 VDD1.n7 185
R1433 VDD1.n37 VDD1.n36 185
R1434 VDD1.n42 VDD1.n41 185
R1435 VDD1.n44 VDD1.n43 185
R1436 VDD1.n33 VDD1.n32 185
R1437 VDD1.n50 VDD1.n49 185
R1438 VDD1.n52 VDD1.n51 185
R1439 VDD1.n9 VDD1.t6 147.672
R1440 VDD1.n38 VDD1.t2 147.672
R1441 VDD1.n22 VDD1.n21 104.615
R1442 VDD1.n21 VDD1.n3 104.615
R1443 VDD1.n14 VDD1.n3 104.615
R1444 VDD1.n14 VDD1.n13 104.615
R1445 VDD1.n13 VDD1.n7 104.615
R1446 VDD1.n42 VDD1.n36 104.615
R1447 VDD1.n43 VDD1.n42 104.615
R1448 VDD1.n43 VDD1.n32 104.615
R1449 VDD1.n50 VDD1.n32 104.615
R1450 VDD1.n51 VDD1.n50 104.615
R1451 VDD1.n59 VDD1.n58 68.6452
R1452 VDD1.n28 VDD1.n27 67.2977
R1453 VDD1.n61 VDD1.n60 67.2975
R1454 VDD1.n57 VDD1.n56 67.2975
R1455 VDD1.t6 VDD1.n7 52.3082
R1456 VDD1.t2 VDD1.n36 52.3082
R1457 VDD1.n28 VDD1.n26 49.3773
R1458 VDD1.n57 VDD1.n55 49.3773
R1459 VDD1.n61 VDD1.n59 38.6108
R1460 VDD1.n9 VDD1.n8 15.6666
R1461 VDD1.n38 VDD1.n37 15.6666
R1462 VDD1.n12 VDD1.n11 12.8005
R1463 VDD1.n41 VDD1.n40 12.8005
R1464 VDD1.n15 VDD1.n6 12.0247
R1465 VDD1.n44 VDD1.n35 12.0247
R1466 VDD1.n16 VDD1.n4 11.249
R1467 VDD1.n45 VDD1.n33 11.249
R1468 VDD1.n20 VDD1.n19 10.4732
R1469 VDD1.n49 VDD1.n48 10.4732
R1470 VDD1.n23 VDD1.n2 9.69747
R1471 VDD1.n52 VDD1.n31 9.69747
R1472 VDD1.n26 VDD1.n25 9.45567
R1473 VDD1.n55 VDD1.n54 9.45567
R1474 VDD1.n25 VDD1.n24 9.3005
R1475 VDD1.n2 VDD1.n1 9.3005
R1476 VDD1.n19 VDD1.n18 9.3005
R1477 VDD1.n17 VDD1.n16 9.3005
R1478 VDD1.n6 VDD1.n5 9.3005
R1479 VDD1.n11 VDD1.n10 9.3005
R1480 VDD1.n54 VDD1.n53 9.3005
R1481 VDD1.n31 VDD1.n30 9.3005
R1482 VDD1.n48 VDD1.n47 9.3005
R1483 VDD1.n46 VDD1.n45 9.3005
R1484 VDD1.n35 VDD1.n34 9.3005
R1485 VDD1.n40 VDD1.n39 9.3005
R1486 VDD1.n24 VDD1.n0 8.92171
R1487 VDD1.n53 VDD1.n29 8.92171
R1488 VDD1.n26 VDD1.n0 5.04292
R1489 VDD1.n55 VDD1.n29 5.04292
R1490 VDD1.n10 VDD1.n9 4.38687
R1491 VDD1.n39 VDD1.n38 4.38687
R1492 VDD1.n24 VDD1.n23 4.26717
R1493 VDD1.n53 VDD1.n52 4.26717
R1494 VDD1.n60 VDD1.t3 3.80088
R1495 VDD1.n60 VDD1.t7 3.80088
R1496 VDD1.n27 VDD1.t9 3.80088
R1497 VDD1.n27 VDD1.t4 3.80088
R1498 VDD1.n58 VDD1.t0 3.80088
R1499 VDD1.n58 VDD1.t5 3.80088
R1500 VDD1.n56 VDD1.t1 3.80088
R1501 VDD1.n56 VDD1.t8 3.80088
R1502 VDD1.n20 VDD1.n2 3.49141
R1503 VDD1.n49 VDD1.n31 3.49141
R1504 VDD1.n19 VDD1.n4 2.71565
R1505 VDD1.n48 VDD1.n33 2.71565
R1506 VDD1.n16 VDD1.n15 1.93989
R1507 VDD1.n45 VDD1.n44 1.93989
R1508 VDD1 VDD1.n61 1.34533
R1509 VDD1.n12 VDD1.n6 1.16414
R1510 VDD1.n41 VDD1.n35 1.16414
R1511 VDD1 VDD1.n28 0.526362
R1512 VDD1.n59 VDD1.n57 0.412826
R1513 VDD1.n11 VDD1.n8 0.388379
R1514 VDD1.n40 VDD1.n37 0.388379
R1515 VDD1.n25 VDD1.n1 0.155672
R1516 VDD1.n18 VDD1.n1 0.155672
R1517 VDD1.n18 VDD1.n17 0.155672
R1518 VDD1.n17 VDD1.n5 0.155672
R1519 VDD1.n10 VDD1.n5 0.155672
R1520 VDD1.n39 VDD1.n34 0.155672
R1521 VDD1.n46 VDD1.n34 0.155672
R1522 VDD1.n47 VDD1.n46 0.155672
R1523 VDD1.n47 VDD1.n30 0.155672
R1524 VDD1.n54 VDD1.n30 0.155672
R1525 VTAIL.n120 VTAIL.n98 289.615
R1526 VTAIL.n24 VTAIL.n2 289.615
R1527 VTAIL.n92 VTAIL.n70 289.615
R1528 VTAIL.n60 VTAIL.n38 289.615
R1529 VTAIL.n106 VTAIL.n105 185
R1530 VTAIL.n111 VTAIL.n110 185
R1531 VTAIL.n113 VTAIL.n112 185
R1532 VTAIL.n102 VTAIL.n101 185
R1533 VTAIL.n119 VTAIL.n118 185
R1534 VTAIL.n121 VTAIL.n120 185
R1535 VTAIL.n10 VTAIL.n9 185
R1536 VTAIL.n15 VTAIL.n14 185
R1537 VTAIL.n17 VTAIL.n16 185
R1538 VTAIL.n6 VTAIL.n5 185
R1539 VTAIL.n23 VTAIL.n22 185
R1540 VTAIL.n25 VTAIL.n24 185
R1541 VTAIL.n93 VTAIL.n92 185
R1542 VTAIL.n91 VTAIL.n90 185
R1543 VTAIL.n74 VTAIL.n73 185
R1544 VTAIL.n85 VTAIL.n84 185
R1545 VTAIL.n83 VTAIL.n82 185
R1546 VTAIL.n78 VTAIL.n77 185
R1547 VTAIL.n61 VTAIL.n60 185
R1548 VTAIL.n59 VTAIL.n58 185
R1549 VTAIL.n42 VTAIL.n41 185
R1550 VTAIL.n53 VTAIL.n52 185
R1551 VTAIL.n51 VTAIL.n50 185
R1552 VTAIL.n46 VTAIL.n45 185
R1553 VTAIL.n107 VTAIL.t18 147.672
R1554 VTAIL.n11 VTAIL.t12 147.672
R1555 VTAIL.n79 VTAIL.t9 147.672
R1556 VTAIL.n47 VTAIL.t1 147.672
R1557 VTAIL.n111 VTAIL.n105 104.615
R1558 VTAIL.n112 VTAIL.n111 104.615
R1559 VTAIL.n112 VTAIL.n101 104.615
R1560 VTAIL.n119 VTAIL.n101 104.615
R1561 VTAIL.n120 VTAIL.n119 104.615
R1562 VTAIL.n15 VTAIL.n9 104.615
R1563 VTAIL.n16 VTAIL.n15 104.615
R1564 VTAIL.n16 VTAIL.n5 104.615
R1565 VTAIL.n23 VTAIL.n5 104.615
R1566 VTAIL.n24 VTAIL.n23 104.615
R1567 VTAIL.n92 VTAIL.n91 104.615
R1568 VTAIL.n91 VTAIL.n73 104.615
R1569 VTAIL.n84 VTAIL.n73 104.615
R1570 VTAIL.n84 VTAIL.n83 104.615
R1571 VTAIL.n83 VTAIL.n77 104.615
R1572 VTAIL.n60 VTAIL.n59 104.615
R1573 VTAIL.n59 VTAIL.n41 104.615
R1574 VTAIL.n52 VTAIL.n41 104.615
R1575 VTAIL.n52 VTAIL.n51 104.615
R1576 VTAIL.n51 VTAIL.n45 104.615
R1577 VTAIL.t18 VTAIL.n105 52.3082
R1578 VTAIL.t12 VTAIL.n9 52.3082
R1579 VTAIL.t9 VTAIL.n77 52.3082
R1580 VTAIL.t1 VTAIL.n45 52.3082
R1581 VTAIL.n69 VTAIL.n68 50.6189
R1582 VTAIL.n67 VTAIL.n66 50.6189
R1583 VTAIL.n37 VTAIL.n36 50.6189
R1584 VTAIL.n35 VTAIL.n34 50.6189
R1585 VTAIL.n127 VTAIL.n126 50.6187
R1586 VTAIL.n1 VTAIL.n0 50.6187
R1587 VTAIL.n31 VTAIL.n30 50.6187
R1588 VTAIL.n33 VTAIL.n32 50.6187
R1589 VTAIL.n125 VTAIL.n124 30.8278
R1590 VTAIL.n29 VTAIL.n28 30.8278
R1591 VTAIL.n97 VTAIL.n96 30.8278
R1592 VTAIL.n65 VTAIL.n64 30.8278
R1593 VTAIL.n35 VTAIL.n33 20.5996
R1594 VTAIL.n125 VTAIL.n97 18.7289
R1595 VTAIL.n107 VTAIL.n106 15.6666
R1596 VTAIL.n11 VTAIL.n10 15.6666
R1597 VTAIL.n79 VTAIL.n78 15.6666
R1598 VTAIL.n47 VTAIL.n46 15.6666
R1599 VTAIL.n110 VTAIL.n109 12.8005
R1600 VTAIL.n14 VTAIL.n13 12.8005
R1601 VTAIL.n82 VTAIL.n81 12.8005
R1602 VTAIL.n50 VTAIL.n49 12.8005
R1603 VTAIL.n113 VTAIL.n104 12.0247
R1604 VTAIL.n17 VTAIL.n8 12.0247
R1605 VTAIL.n85 VTAIL.n76 12.0247
R1606 VTAIL.n53 VTAIL.n44 12.0247
R1607 VTAIL.n114 VTAIL.n102 11.249
R1608 VTAIL.n18 VTAIL.n6 11.249
R1609 VTAIL.n86 VTAIL.n74 11.249
R1610 VTAIL.n54 VTAIL.n42 11.249
R1611 VTAIL.n118 VTAIL.n117 10.4732
R1612 VTAIL.n22 VTAIL.n21 10.4732
R1613 VTAIL.n90 VTAIL.n89 10.4732
R1614 VTAIL.n58 VTAIL.n57 10.4732
R1615 VTAIL.n121 VTAIL.n100 9.69747
R1616 VTAIL.n25 VTAIL.n4 9.69747
R1617 VTAIL.n93 VTAIL.n72 9.69747
R1618 VTAIL.n61 VTAIL.n40 9.69747
R1619 VTAIL.n124 VTAIL.n123 9.45567
R1620 VTAIL.n28 VTAIL.n27 9.45567
R1621 VTAIL.n96 VTAIL.n95 9.45567
R1622 VTAIL.n64 VTAIL.n63 9.45567
R1623 VTAIL.n123 VTAIL.n122 9.3005
R1624 VTAIL.n100 VTAIL.n99 9.3005
R1625 VTAIL.n117 VTAIL.n116 9.3005
R1626 VTAIL.n115 VTAIL.n114 9.3005
R1627 VTAIL.n104 VTAIL.n103 9.3005
R1628 VTAIL.n109 VTAIL.n108 9.3005
R1629 VTAIL.n27 VTAIL.n26 9.3005
R1630 VTAIL.n4 VTAIL.n3 9.3005
R1631 VTAIL.n21 VTAIL.n20 9.3005
R1632 VTAIL.n19 VTAIL.n18 9.3005
R1633 VTAIL.n8 VTAIL.n7 9.3005
R1634 VTAIL.n13 VTAIL.n12 9.3005
R1635 VTAIL.n95 VTAIL.n94 9.3005
R1636 VTAIL.n72 VTAIL.n71 9.3005
R1637 VTAIL.n89 VTAIL.n88 9.3005
R1638 VTAIL.n87 VTAIL.n86 9.3005
R1639 VTAIL.n76 VTAIL.n75 9.3005
R1640 VTAIL.n81 VTAIL.n80 9.3005
R1641 VTAIL.n63 VTAIL.n62 9.3005
R1642 VTAIL.n40 VTAIL.n39 9.3005
R1643 VTAIL.n57 VTAIL.n56 9.3005
R1644 VTAIL.n55 VTAIL.n54 9.3005
R1645 VTAIL.n44 VTAIL.n43 9.3005
R1646 VTAIL.n49 VTAIL.n48 9.3005
R1647 VTAIL.n122 VTAIL.n98 8.92171
R1648 VTAIL.n26 VTAIL.n2 8.92171
R1649 VTAIL.n94 VTAIL.n70 8.92171
R1650 VTAIL.n62 VTAIL.n38 8.92171
R1651 VTAIL.n124 VTAIL.n98 5.04292
R1652 VTAIL.n28 VTAIL.n2 5.04292
R1653 VTAIL.n96 VTAIL.n70 5.04292
R1654 VTAIL.n64 VTAIL.n38 5.04292
R1655 VTAIL.n108 VTAIL.n107 4.38687
R1656 VTAIL.n12 VTAIL.n11 4.38687
R1657 VTAIL.n80 VTAIL.n79 4.38687
R1658 VTAIL.n48 VTAIL.n47 4.38687
R1659 VTAIL.n122 VTAIL.n121 4.26717
R1660 VTAIL.n26 VTAIL.n25 4.26717
R1661 VTAIL.n94 VTAIL.n93 4.26717
R1662 VTAIL.n62 VTAIL.n61 4.26717
R1663 VTAIL.n126 VTAIL.t4 3.80088
R1664 VTAIL.n126 VTAIL.t19 3.80088
R1665 VTAIL.n0 VTAIL.t5 3.80088
R1666 VTAIL.n0 VTAIL.t2 3.80088
R1667 VTAIL.n30 VTAIL.t8 3.80088
R1668 VTAIL.n30 VTAIL.t16 3.80088
R1669 VTAIL.n32 VTAIL.t15 3.80088
R1670 VTAIL.n32 VTAIL.t11 3.80088
R1671 VTAIL.n68 VTAIL.t13 3.80088
R1672 VTAIL.n68 VTAIL.t14 3.80088
R1673 VTAIL.n66 VTAIL.t7 3.80088
R1674 VTAIL.n66 VTAIL.t10 3.80088
R1675 VTAIL.n36 VTAIL.t0 3.80088
R1676 VTAIL.n36 VTAIL.t3 3.80088
R1677 VTAIL.n34 VTAIL.t17 3.80088
R1678 VTAIL.n34 VTAIL.t6 3.80088
R1679 VTAIL.n118 VTAIL.n100 3.49141
R1680 VTAIL.n22 VTAIL.n4 3.49141
R1681 VTAIL.n90 VTAIL.n72 3.49141
R1682 VTAIL.n58 VTAIL.n40 3.49141
R1683 VTAIL.n117 VTAIL.n102 2.71565
R1684 VTAIL.n21 VTAIL.n6 2.71565
R1685 VTAIL.n89 VTAIL.n74 2.71565
R1686 VTAIL.n57 VTAIL.n42 2.71565
R1687 VTAIL.n114 VTAIL.n113 1.93989
R1688 VTAIL.n18 VTAIL.n17 1.93989
R1689 VTAIL.n86 VTAIL.n85 1.93989
R1690 VTAIL.n54 VTAIL.n53 1.93989
R1691 VTAIL.n37 VTAIL.n35 1.87119
R1692 VTAIL.n65 VTAIL.n37 1.87119
R1693 VTAIL.n69 VTAIL.n67 1.87119
R1694 VTAIL.n97 VTAIL.n69 1.87119
R1695 VTAIL.n33 VTAIL.n31 1.87119
R1696 VTAIL.n31 VTAIL.n29 1.87119
R1697 VTAIL.n127 VTAIL.n125 1.87119
R1698 VTAIL VTAIL.n1 1.46171
R1699 VTAIL.n67 VTAIL.n65 1.40567
R1700 VTAIL.n29 VTAIL.n1 1.40567
R1701 VTAIL.n110 VTAIL.n104 1.16414
R1702 VTAIL.n14 VTAIL.n8 1.16414
R1703 VTAIL.n82 VTAIL.n76 1.16414
R1704 VTAIL.n50 VTAIL.n44 1.16414
R1705 VTAIL VTAIL.n127 0.409983
R1706 VTAIL.n109 VTAIL.n106 0.388379
R1707 VTAIL.n13 VTAIL.n10 0.388379
R1708 VTAIL.n81 VTAIL.n78 0.388379
R1709 VTAIL.n49 VTAIL.n46 0.388379
R1710 VTAIL.n108 VTAIL.n103 0.155672
R1711 VTAIL.n115 VTAIL.n103 0.155672
R1712 VTAIL.n116 VTAIL.n115 0.155672
R1713 VTAIL.n116 VTAIL.n99 0.155672
R1714 VTAIL.n123 VTAIL.n99 0.155672
R1715 VTAIL.n12 VTAIL.n7 0.155672
R1716 VTAIL.n19 VTAIL.n7 0.155672
R1717 VTAIL.n20 VTAIL.n19 0.155672
R1718 VTAIL.n20 VTAIL.n3 0.155672
R1719 VTAIL.n27 VTAIL.n3 0.155672
R1720 VTAIL.n95 VTAIL.n71 0.155672
R1721 VTAIL.n88 VTAIL.n71 0.155672
R1722 VTAIL.n88 VTAIL.n87 0.155672
R1723 VTAIL.n87 VTAIL.n75 0.155672
R1724 VTAIL.n80 VTAIL.n75 0.155672
R1725 VTAIL.n63 VTAIL.n39 0.155672
R1726 VTAIL.n56 VTAIL.n39 0.155672
R1727 VTAIL.n56 VTAIL.n55 0.155672
R1728 VTAIL.n55 VTAIL.n43 0.155672
R1729 VTAIL.n48 VTAIL.n43 0.155672
R1730 VN.n31 VN.n30 181.363
R1731 VN.n63 VN.n62 181.363
R1732 VN.n61 VN.n32 161.3
R1733 VN.n60 VN.n59 161.3
R1734 VN.n58 VN.n33 161.3
R1735 VN.n57 VN.n56 161.3
R1736 VN.n55 VN.n34 161.3
R1737 VN.n53 VN.n52 161.3
R1738 VN.n51 VN.n35 161.3
R1739 VN.n50 VN.n49 161.3
R1740 VN.n48 VN.n36 161.3
R1741 VN.n46 VN.n45 161.3
R1742 VN.n44 VN.n37 161.3
R1743 VN.n43 VN.n42 161.3
R1744 VN.n41 VN.n38 161.3
R1745 VN.n29 VN.n0 161.3
R1746 VN.n28 VN.n27 161.3
R1747 VN.n26 VN.n1 161.3
R1748 VN.n25 VN.n24 161.3
R1749 VN.n23 VN.n2 161.3
R1750 VN.n21 VN.n20 161.3
R1751 VN.n19 VN.n3 161.3
R1752 VN.n18 VN.n17 161.3
R1753 VN.n16 VN.n4 161.3
R1754 VN.n14 VN.n13 161.3
R1755 VN.n12 VN.n5 161.3
R1756 VN.n11 VN.n10 161.3
R1757 VN.n9 VN.n6 161.3
R1758 VN.n7 VN.t7 103.059
R1759 VN.n39 VN.t5 103.059
R1760 VN.n8 VN.t1 68.2402
R1761 VN.n15 VN.t9 68.2402
R1762 VN.n22 VN.t6 68.2402
R1763 VN.n30 VN.t3 68.2402
R1764 VN.n40 VN.t2 68.2402
R1765 VN.n47 VN.t4 68.2402
R1766 VN.n54 VN.t0 68.2402
R1767 VN.n62 VN.t8 68.2402
R1768 VN.n10 VN.n5 56.5193
R1769 VN.n17 VN.n3 56.5193
R1770 VN.n42 VN.n37 56.5193
R1771 VN.n49 VN.n35 56.5193
R1772 VN.n8 VN.n7 48.825
R1773 VN.n40 VN.n39 48.825
R1774 VN VN.n63 44.1425
R1775 VN.n28 VN.n1 40.979
R1776 VN.n60 VN.n33 40.979
R1777 VN.n24 VN.n1 40.0078
R1778 VN.n56 VN.n33 40.0078
R1779 VN.n10 VN.n9 24.4675
R1780 VN.n14 VN.n5 24.4675
R1781 VN.n17 VN.n16 24.4675
R1782 VN.n21 VN.n3 24.4675
R1783 VN.n24 VN.n23 24.4675
R1784 VN.n29 VN.n28 24.4675
R1785 VN.n42 VN.n41 24.4675
R1786 VN.n49 VN.n48 24.4675
R1787 VN.n46 VN.n37 24.4675
R1788 VN.n56 VN.n55 24.4675
R1789 VN.n53 VN.n35 24.4675
R1790 VN.n61 VN.n60 24.4675
R1791 VN.n9 VN.n8 20.5528
R1792 VN.n22 VN.n21 20.5528
R1793 VN.n41 VN.n40 20.5528
R1794 VN.n54 VN.n53 20.5528
R1795 VN.n39 VN.n38 12.2488
R1796 VN.n7 VN.n6 12.2488
R1797 VN.n15 VN.n14 12.234
R1798 VN.n16 VN.n15 12.234
R1799 VN.n48 VN.n47 12.234
R1800 VN.n47 VN.n46 12.234
R1801 VN.n30 VN.n29 4.40456
R1802 VN.n62 VN.n61 4.40456
R1803 VN.n23 VN.n22 3.91522
R1804 VN.n55 VN.n54 3.91522
R1805 VN.n63 VN.n32 0.189894
R1806 VN.n59 VN.n32 0.189894
R1807 VN.n59 VN.n58 0.189894
R1808 VN.n58 VN.n57 0.189894
R1809 VN.n57 VN.n34 0.189894
R1810 VN.n52 VN.n34 0.189894
R1811 VN.n52 VN.n51 0.189894
R1812 VN.n51 VN.n50 0.189894
R1813 VN.n50 VN.n36 0.189894
R1814 VN.n45 VN.n36 0.189894
R1815 VN.n45 VN.n44 0.189894
R1816 VN.n44 VN.n43 0.189894
R1817 VN.n43 VN.n38 0.189894
R1818 VN.n11 VN.n6 0.189894
R1819 VN.n12 VN.n11 0.189894
R1820 VN.n13 VN.n12 0.189894
R1821 VN.n13 VN.n4 0.189894
R1822 VN.n18 VN.n4 0.189894
R1823 VN.n19 VN.n18 0.189894
R1824 VN.n20 VN.n19 0.189894
R1825 VN.n20 VN.n2 0.189894
R1826 VN.n25 VN.n2 0.189894
R1827 VN.n26 VN.n25 0.189894
R1828 VN.n27 VN.n26 0.189894
R1829 VN.n27 VN.n0 0.189894
R1830 VN.n31 VN.n0 0.189894
R1831 VN VN.n31 0.0516364
R1832 VDD2.n53 VDD2.n31 289.615
R1833 VDD2.n22 VDD2.n0 289.615
R1834 VDD2.n54 VDD2.n53 185
R1835 VDD2.n52 VDD2.n51 185
R1836 VDD2.n35 VDD2.n34 185
R1837 VDD2.n46 VDD2.n45 185
R1838 VDD2.n44 VDD2.n43 185
R1839 VDD2.n39 VDD2.n38 185
R1840 VDD2.n8 VDD2.n7 185
R1841 VDD2.n13 VDD2.n12 185
R1842 VDD2.n15 VDD2.n14 185
R1843 VDD2.n4 VDD2.n3 185
R1844 VDD2.n21 VDD2.n20 185
R1845 VDD2.n23 VDD2.n22 185
R1846 VDD2.n40 VDD2.t1 147.672
R1847 VDD2.n9 VDD2.t2 147.672
R1848 VDD2.n53 VDD2.n52 104.615
R1849 VDD2.n52 VDD2.n34 104.615
R1850 VDD2.n45 VDD2.n34 104.615
R1851 VDD2.n45 VDD2.n44 104.615
R1852 VDD2.n44 VDD2.n38 104.615
R1853 VDD2.n13 VDD2.n7 104.615
R1854 VDD2.n14 VDD2.n13 104.615
R1855 VDD2.n14 VDD2.n3 104.615
R1856 VDD2.n21 VDD2.n3 104.615
R1857 VDD2.n22 VDD2.n21 104.615
R1858 VDD2.n30 VDD2.n29 68.6452
R1859 VDD2 VDD2.n61 68.6424
R1860 VDD2.n60 VDD2.n59 67.2977
R1861 VDD2.n28 VDD2.n27 67.2975
R1862 VDD2.t1 VDD2.n38 52.3082
R1863 VDD2.t2 VDD2.n7 52.3082
R1864 VDD2.n28 VDD2.n26 49.3773
R1865 VDD2.n58 VDD2.n57 47.5066
R1866 VDD2.n58 VDD2.n30 37.0924
R1867 VDD2.n40 VDD2.n39 15.6666
R1868 VDD2.n9 VDD2.n8 15.6666
R1869 VDD2.n43 VDD2.n42 12.8005
R1870 VDD2.n12 VDD2.n11 12.8005
R1871 VDD2.n46 VDD2.n37 12.0247
R1872 VDD2.n15 VDD2.n6 12.0247
R1873 VDD2.n47 VDD2.n35 11.249
R1874 VDD2.n16 VDD2.n4 11.249
R1875 VDD2.n51 VDD2.n50 10.4732
R1876 VDD2.n20 VDD2.n19 10.4732
R1877 VDD2.n54 VDD2.n33 9.69747
R1878 VDD2.n23 VDD2.n2 9.69747
R1879 VDD2.n57 VDD2.n56 9.45567
R1880 VDD2.n26 VDD2.n25 9.45567
R1881 VDD2.n56 VDD2.n55 9.3005
R1882 VDD2.n33 VDD2.n32 9.3005
R1883 VDD2.n50 VDD2.n49 9.3005
R1884 VDD2.n48 VDD2.n47 9.3005
R1885 VDD2.n37 VDD2.n36 9.3005
R1886 VDD2.n42 VDD2.n41 9.3005
R1887 VDD2.n25 VDD2.n24 9.3005
R1888 VDD2.n2 VDD2.n1 9.3005
R1889 VDD2.n19 VDD2.n18 9.3005
R1890 VDD2.n17 VDD2.n16 9.3005
R1891 VDD2.n6 VDD2.n5 9.3005
R1892 VDD2.n11 VDD2.n10 9.3005
R1893 VDD2.n55 VDD2.n31 8.92171
R1894 VDD2.n24 VDD2.n0 8.92171
R1895 VDD2.n57 VDD2.n31 5.04292
R1896 VDD2.n26 VDD2.n0 5.04292
R1897 VDD2.n41 VDD2.n40 4.38687
R1898 VDD2.n10 VDD2.n9 4.38687
R1899 VDD2.n55 VDD2.n54 4.26717
R1900 VDD2.n24 VDD2.n23 4.26717
R1901 VDD2.n61 VDD2.t7 3.80088
R1902 VDD2.n61 VDD2.t4 3.80088
R1903 VDD2.n59 VDD2.t9 3.80088
R1904 VDD2.n59 VDD2.t5 3.80088
R1905 VDD2.n29 VDD2.t3 3.80088
R1906 VDD2.n29 VDD2.t6 3.80088
R1907 VDD2.n27 VDD2.t8 3.80088
R1908 VDD2.n27 VDD2.t0 3.80088
R1909 VDD2.n51 VDD2.n33 3.49141
R1910 VDD2.n20 VDD2.n2 3.49141
R1911 VDD2.n50 VDD2.n35 2.71565
R1912 VDD2.n19 VDD2.n4 2.71565
R1913 VDD2.n47 VDD2.n46 1.93989
R1914 VDD2.n16 VDD2.n15 1.93989
R1915 VDD2.n60 VDD2.n58 1.87119
R1916 VDD2.n43 VDD2.n37 1.16414
R1917 VDD2.n12 VDD2.n6 1.16414
R1918 VDD2 VDD2.n60 0.526362
R1919 VDD2.n30 VDD2.n28 0.412826
R1920 VDD2.n42 VDD2.n39 0.388379
R1921 VDD2.n11 VDD2.n8 0.388379
R1922 VDD2.n56 VDD2.n32 0.155672
R1923 VDD2.n49 VDD2.n32 0.155672
R1924 VDD2.n49 VDD2.n48 0.155672
R1925 VDD2.n48 VDD2.n36 0.155672
R1926 VDD2.n41 VDD2.n36 0.155672
R1927 VDD2.n10 VDD2.n5 0.155672
R1928 VDD2.n17 VDD2.n5 0.155672
R1929 VDD2.n18 VDD2.n17 0.155672
R1930 VDD2.n18 VDD2.n1 0.155672
R1931 VDD2.n25 VDD2.n1 0.155672
C0 VDD2 VP 0.489976f
C1 VTAIL VDD1 6.78849f
C2 VP VDD1 4.88539f
C3 VDD2 VN 4.55356f
C4 VP VTAIL 5.33702f
C5 VN VDD1 0.151468f
C6 VN VTAIL 5.3228f
C7 VDD2 VDD1 1.67791f
C8 VN VP 6.01874f
C9 VDD2 VTAIL 6.83545f
C10 VDD2 B 5.091876f
C11 VDD1 B 5.076347f
C12 VTAIL B 4.615823f
C13 VN B 13.8172f
C14 VP B 12.343748f
C15 VDD2.n0 B 0.03029f
C16 VDD2.n1 B 0.022751f
C17 VDD2.n2 B 0.012225f
C18 VDD2.n3 B 0.028896f
C19 VDD2.n4 B 0.012945f
C20 VDD2.n5 B 0.022751f
C21 VDD2.n6 B 0.012225f
C22 VDD2.n7 B 0.021672f
C23 VDD2.n8 B 0.017066f
C24 VDD2.t2 B 0.047127f
C25 VDD2.n9 B 0.093017f
C26 VDD2.n10 B 0.458715f
C27 VDD2.n11 B 0.012225f
C28 VDD2.n12 B 0.012945f
C29 VDD2.n13 B 0.028896f
C30 VDD2.n14 B 0.028896f
C31 VDD2.n15 B 0.012945f
C32 VDD2.n16 B 0.012225f
C33 VDD2.n17 B 0.022751f
C34 VDD2.n18 B 0.022751f
C35 VDD2.n19 B 0.012225f
C36 VDD2.n20 B 0.012945f
C37 VDD2.n21 B 0.028896f
C38 VDD2.n22 B 0.05957f
C39 VDD2.n23 B 0.012945f
C40 VDD2.n24 B 0.012225f
C41 VDD2.n25 B 0.050412f
C42 VDD2.n26 B 0.055492f
C43 VDD2.t8 B 0.093668f
C44 VDD2.t0 B 0.093668f
C45 VDD2.n27 B 0.766874f
C46 VDD2.n28 B 0.523825f
C47 VDD2.t3 B 0.093668f
C48 VDD2.t6 B 0.093668f
C49 VDD2.n29 B 0.775272f
C50 VDD2.n30 B 1.90519f
C51 VDD2.n31 B 0.03029f
C52 VDD2.n32 B 0.022751f
C53 VDD2.n33 B 0.012225f
C54 VDD2.n34 B 0.028896f
C55 VDD2.n35 B 0.012945f
C56 VDD2.n36 B 0.022751f
C57 VDD2.n37 B 0.012225f
C58 VDD2.n38 B 0.021672f
C59 VDD2.n39 B 0.017066f
C60 VDD2.t1 B 0.047127f
C61 VDD2.n40 B 0.093017f
C62 VDD2.n41 B 0.458715f
C63 VDD2.n42 B 0.012225f
C64 VDD2.n43 B 0.012945f
C65 VDD2.n44 B 0.028896f
C66 VDD2.n45 B 0.028896f
C67 VDD2.n46 B 0.012945f
C68 VDD2.n47 B 0.012225f
C69 VDD2.n48 B 0.022751f
C70 VDD2.n49 B 0.022751f
C71 VDD2.n50 B 0.012225f
C72 VDD2.n51 B 0.012945f
C73 VDD2.n52 B 0.028896f
C74 VDD2.n53 B 0.05957f
C75 VDD2.n54 B 0.012945f
C76 VDD2.n55 B 0.012225f
C77 VDD2.n56 B 0.050412f
C78 VDD2.n57 B 0.048684f
C79 VDD2.n58 B 1.87421f
C80 VDD2.t9 B 0.093668f
C81 VDD2.t5 B 0.093668f
C82 VDD2.n59 B 0.766878f
C83 VDD2.n60 B 0.357972f
C84 VDD2.t7 B 0.093668f
C85 VDD2.t4 B 0.093668f
C86 VDD2.n61 B 0.775243f
C87 VN.n0 B 0.029329f
C88 VN.t3 B 0.737526f
C89 VN.n1 B 0.02372f
C90 VN.n2 B 0.029329f
C91 VN.t6 B 0.737526f
C92 VN.n3 B 0.035871f
C93 VN.n4 B 0.029329f
C94 VN.t9 B 0.737526f
C95 VN.n5 B 0.049764f
C96 VN.n6 B 0.217251f
C97 VN.t1 B 0.737526f
C98 VN.t7 B 0.883214f
C99 VN.n7 B 0.348749f
C100 VN.n8 B 0.364974f
C101 VN.n9 B 0.050344f
C102 VN.n10 B 0.035871f
C103 VN.n11 B 0.029329f
C104 VN.n12 B 0.029329f
C105 VN.n13 B 0.029329f
C106 VN.n14 B 0.041168f
C107 VN.n15 B 0.289633f
C108 VN.n16 B 0.041168f
C109 VN.n17 B 0.049764f
C110 VN.n18 B 0.029329f
C111 VN.n19 B 0.029329f
C112 VN.n20 B 0.029329f
C113 VN.n21 B 0.050344f
C114 VN.n22 B 0.289633f
C115 VN.n23 B 0.031993f
C116 VN.n24 B 0.058435f
C117 VN.n25 B 0.029329f
C118 VN.n26 B 0.029329f
C119 VN.n27 B 0.029329f
C120 VN.n28 B 0.058141f
C121 VN.n29 B 0.032533f
C122 VN.n30 B 0.358889f
C123 VN.n31 B 0.031343f
C124 VN.n32 B 0.029329f
C125 VN.t8 B 0.737526f
C126 VN.n33 B 0.02372f
C127 VN.n34 B 0.029329f
C128 VN.t0 B 0.737526f
C129 VN.n35 B 0.035871f
C130 VN.n36 B 0.029329f
C131 VN.t4 B 0.737526f
C132 VN.n37 B 0.049764f
C133 VN.n38 B 0.217251f
C134 VN.t2 B 0.737526f
C135 VN.t5 B 0.883214f
C136 VN.n39 B 0.348749f
C137 VN.n40 B 0.364974f
C138 VN.n41 B 0.050344f
C139 VN.n42 B 0.035871f
C140 VN.n43 B 0.029329f
C141 VN.n44 B 0.029329f
C142 VN.n45 B 0.029329f
C143 VN.n46 B 0.041168f
C144 VN.n47 B 0.289633f
C145 VN.n48 B 0.041168f
C146 VN.n49 B 0.049764f
C147 VN.n50 B 0.029329f
C148 VN.n51 B 0.029329f
C149 VN.n52 B 0.029329f
C150 VN.n53 B 0.050344f
C151 VN.n54 B 0.289633f
C152 VN.n55 B 0.031993f
C153 VN.n56 B 0.058435f
C154 VN.n57 B 0.029329f
C155 VN.n58 B 0.029329f
C156 VN.n59 B 0.029329f
C157 VN.n60 B 0.058141f
C158 VN.n61 B 0.032533f
C159 VN.n62 B 0.358889f
C160 VN.n63 B 1.32304f
C161 VTAIL.t5 B 0.116116f
C162 VTAIL.t2 B 0.116116f
C163 VTAIL.n0 B 0.877964f
C164 VTAIL.n1 B 0.520814f
C165 VTAIL.n2 B 0.037549f
C166 VTAIL.n3 B 0.028203f
C167 VTAIL.n4 B 0.015155f
C168 VTAIL.n5 B 0.035821f
C169 VTAIL.n6 B 0.016047f
C170 VTAIL.n7 B 0.028203f
C171 VTAIL.n8 B 0.015155f
C172 VTAIL.n9 B 0.026866f
C173 VTAIL.n10 B 0.021155f
C174 VTAIL.t12 B 0.058421f
C175 VTAIL.n11 B 0.115308f
C176 VTAIL.n12 B 0.568645f
C177 VTAIL.n13 B 0.015155f
C178 VTAIL.n14 B 0.016047f
C179 VTAIL.n15 B 0.035821f
C180 VTAIL.n16 B 0.035821f
C181 VTAIL.n17 B 0.016047f
C182 VTAIL.n18 B 0.015155f
C183 VTAIL.n19 B 0.028203f
C184 VTAIL.n20 B 0.028203f
C185 VTAIL.n21 B 0.015155f
C186 VTAIL.n22 B 0.016047f
C187 VTAIL.n23 B 0.035821f
C188 VTAIL.n24 B 0.073846f
C189 VTAIL.n25 B 0.016047f
C190 VTAIL.n26 B 0.015155f
C191 VTAIL.n27 B 0.062494f
C192 VTAIL.n28 B 0.040855f
C193 VTAIL.n29 B 0.320269f
C194 VTAIL.t8 B 0.116116f
C195 VTAIL.t16 B 0.116116f
C196 VTAIL.n30 B 0.877964f
C197 VTAIL.n31 B 0.600332f
C198 VTAIL.t15 B 0.116116f
C199 VTAIL.t11 B 0.116116f
C200 VTAIL.n32 B 0.877964f
C201 VTAIL.n33 B 1.56161f
C202 VTAIL.t17 B 0.116116f
C203 VTAIL.t6 B 0.116116f
C204 VTAIL.n34 B 0.877971f
C205 VTAIL.n35 B 1.5616f
C206 VTAIL.t0 B 0.116116f
C207 VTAIL.t3 B 0.116116f
C208 VTAIL.n36 B 0.877971f
C209 VTAIL.n37 B 0.600326f
C210 VTAIL.n38 B 0.037549f
C211 VTAIL.n39 B 0.028203f
C212 VTAIL.n40 B 0.015155f
C213 VTAIL.n41 B 0.035821f
C214 VTAIL.n42 B 0.016047f
C215 VTAIL.n43 B 0.028203f
C216 VTAIL.n44 B 0.015155f
C217 VTAIL.n45 B 0.026866f
C218 VTAIL.n46 B 0.021155f
C219 VTAIL.t1 B 0.058421f
C220 VTAIL.n47 B 0.115308f
C221 VTAIL.n48 B 0.568645f
C222 VTAIL.n49 B 0.015155f
C223 VTAIL.n50 B 0.016047f
C224 VTAIL.n51 B 0.035821f
C225 VTAIL.n52 B 0.035821f
C226 VTAIL.n53 B 0.016047f
C227 VTAIL.n54 B 0.015155f
C228 VTAIL.n55 B 0.028203f
C229 VTAIL.n56 B 0.028203f
C230 VTAIL.n57 B 0.015155f
C231 VTAIL.n58 B 0.016047f
C232 VTAIL.n59 B 0.035821f
C233 VTAIL.n60 B 0.073846f
C234 VTAIL.n61 B 0.016047f
C235 VTAIL.n62 B 0.015155f
C236 VTAIL.n63 B 0.062494f
C237 VTAIL.n64 B 0.040855f
C238 VTAIL.n65 B 0.320269f
C239 VTAIL.t7 B 0.116116f
C240 VTAIL.t10 B 0.116116f
C241 VTAIL.n66 B 0.877971f
C242 VTAIL.n67 B 0.558021f
C243 VTAIL.t13 B 0.116116f
C244 VTAIL.t14 B 0.116116f
C245 VTAIL.n68 B 0.877971f
C246 VTAIL.n69 B 0.600326f
C247 VTAIL.n70 B 0.037549f
C248 VTAIL.n71 B 0.028203f
C249 VTAIL.n72 B 0.015155f
C250 VTAIL.n73 B 0.035821f
C251 VTAIL.n74 B 0.016047f
C252 VTAIL.n75 B 0.028203f
C253 VTAIL.n76 B 0.015155f
C254 VTAIL.n77 B 0.026866f
C255 VTAIL.n78 B 0.021155f
C256 VTAIL.t9 B 0.058421f
C257 VTAIL.n79 B 0.115308f
C258 VTAIL.n80 B 0.568645f
C259 VTAIL.n81 B 0.015155f
C260 VTAIL.n82 B 0.016047f
C261 VTAIL.n83 B 0.035821f
C262 VTAIL.n84 B 0.035821f
C263 VTAIL.n85 B 0.016047f
C264 VTAIL.n86 B 0.015155f
C265 VTAIL.n87 B 0.028203f
C266 VTAIL.n88 B 0.028203f
C267 VTAIL.n89 B 0.015155f
C268 VTAIL.n90 B 0.016047f
C269 VTAIL.n91 B 0.035821f
C270 VTAIL.n92 B 0.073846f
C271 VTAIL.n93 B 0.016047f
C272 VTAIL.n94 B 0.015155f
C273 VTAIL.n95 B 0.062494f
C274 VTAIL.n96 B 0.040855f
C275 VTAIL.n97 B 1.15385f
C276 VTAIL.n98 B 0.037549f
C277 VTAIL.n99 B 0.028203f
C278 VTAIL.n100 B 0.015155f
C279 VTAIL.n101 B 0.035821f
C280 VTAIL.n102 B 0.016047f
C281 VTAIL.n103 B 0.028203f
C282 VTAIL.n104 B 0.015155f
C283 VTAIL.n105 B 0.026866f
C284 VTAIL.n106 B 0.021155f
C285 VTAIL.t18 B 0.058421f
C286 VTAIL.n107 B 0.115308f
C287 VTAIL.n108 B 0.568645f
C288 VTAIL.n109 B 0.015155f
C289 VTAIL.n110 B 0.016047f
C290 VTAIL.n111 B 0.035821f
C291 VTAIL.n112 B 0.035821f
C292 VTAIL.n113 B 0.016047f
C293 VTAIL.n114 B 0.015155f
C294 VTAIL.n115 B 0.028203f
C295 VTAIL.n116 B 0.028203f
C296 VTAIL.n117 B 0.015155f
C297 VTAIL.n118 B 0.016047f
C298 VTAIL.n119 B 0.035821f
C299 VTAIL.n120 B 0.073846f
C300 VTAIL.n121 B 0.016047f
C301 VTAIL.n122 B 0.015155f
C302 VTAIL.n123 B 0.062494f
C303 VTAIL.n124 B 0.040855f
C304 VTAIL.n125 B 1.15385f
C305 VTAIL.t4 B 0.116116f
C306 VTAIL.t19 B 0.116116f
C307 VTAIL.n126 B 0.877964f
C308 VTAIL.n127 B 0.467541f
C309 VDD1.n0 B 0.03086f
C310 VDD1.n1 B 0.023179f
C311 VDD1.n2 B 0.012455f
C312 VDD1.n3 B 0.02944f
C313 VDD1.n4 B 0.013188f
C314 VDD1.n5 B 0.023179f
C315 VDD1.n6 B 0.012455f
C316 VDD1.n7 B 0.02208f
C317 VDD1.n8 B 0.017386f
C318 VDD1.t6 B 0.048013f
C319 VDD1.n9 B 0.094766f
C320 VDD1.n10 B 0.467342f
C321 VDD1.n11 B 0.012455f
C322 VDD1.n12 B 0.013188f
C323 VDD1.n13 B 0.02944f
C324 VDD1.n14 B 0.02944f
C325 VDD1.n15 B 0.013188f
C326 VDD1.n16 B 0.012455f
C327 VDD1.n17 B 0.023179f
C328 VDD1.n18 B 0.023179f
C329 VDD1.n19 B 0.012455f
C330 VDD1.n20 B 0.013188f
C331 VDD1.n21 B 0.02944f
C332 VDD1.n22 B 0.06069f
C333 VDD1.n23 B 0.013188f
C334 VDD1.n24 B 0.012455f
C335 VDD1.n25 B 0.051361f
C336 VDD1.n26 B 0.056536f
C337 VDD1.t9 B 0.09543f
C338 VDD1.t4 B 0.09543f
C339 VDD1.n27 B 0.7813f
C340 VDD1.n28 B 0.540849f
C341 VDD1.n29 B 0.03086f
C342 VDD1.n30 B 0.023179f
C343 VDD1.n31 B 0.012455f
C344 VDD1.n32 B 0.02944f
C345 VDD1.n33 B 0.013188f
C346 VDD1.n34 B 0.023179f
C347 VDD1.n35 B 0.012455f
C348 VDD1.n36 B 0.02208f
C349 VDD1.n37 B 0.017386f
C350 VDD1.t2 B 0.048013f
C351 VDD1.n38 B 0.094766f
C352 VDD1.n39 B 0.467342f
C353 VDD1.n40 B 0.012455f
C354 VDD1.n41 B 0.013188f
C355 VDD1.n42 B 0.02944f
C356 VDD1.n43 B 0.02944f
C357 VDD1.n44 B 0.013188f
C358 VDD1.n45 B 0.012455f
C359 VDD1.n46 B 0.023179f
C360 VDD1.n47 B 0.023179f
C361 VDD1.n48 B 0.012455f
C362 VDD1.n49 B 0.013188f
C363 VDD1.n50 B 0.02944f
C364 VDD1.n51 B 0.06069f
C365 VDD1.n52 B 0.013188f
C366 VDD1.n53 B 0.012455f
C367 VDD1.n54 B 0.051361f
C368 VDD1.n55 B 0.056536f
C369 VDD1.t1 B 0.09543f
C370 VDD1.t8 B 0.09543f
C371 VDD1.n56 B 0.781296f
C372 VDD1.n57 B 0.533677f
C373 VDD1.t0 B 0.09543f
C374 VDD1.t5 B 0.09543f
C375 VDD1.n58 B 0.789852f
C376 VDD1.n59 B 2.03396f
C377 VDD1.t3 B 0.09543f
C378 VDD1.t7 B 0.09543f
C379 VDD1.n60 B 0.781296f
C380 VDD1.n61 B 2.15426f
C381 VP.n0 B 0.02996f
C382 VP.t4 B 0.753395f
C383 VP.n1 B 0.024231f
C384 VP.n2 B 0.02996f
C385 VP.t0 B 0.753395f
C386 VP.n3 B 0.036643f
C387 VP.n4 B 0.02996f
C388 VP.t8 B 0.753395f
C389 VP.n5 B 0.050835f
C390 VP.n6 B 0.02996f
C391 VP.t5 B 0.753395f
C392 VP.n7 B 0.059693f
C393 VP.n8 B 0.02996f
C394 VP.t1 B 0.753395f
C395 VP.n9 B 0.366611f
C396 VP.n10 B 0.02996f
C397 VP.t7 B 0.753395f
C398 VP.n11 B 0.024231f
C399 VP.n12 B 0.02996f
C400 VP.t2 B 0.753395f
C401 VP.n13 B 0.036643f
C402 VP.n14 B 0.02996f
C403 VP.t3 B 0.753395f
C404 VP.n15 B 0.050835f
C405 VP.n16 B 0.221926f
C406 VP.t6 B 0.753395f
C407 VP.t9 B 0.902218f
C408 VP.n17 B 0.356253f
C409 VP.n18 B 0.372827f
C410 VP.n19 B 0.051427f
C411 VP.n20 B 0.036643f
C412 VP.n21 B 0.02996f
C413 VP.n22 B 0.02996f
C414 VP.n23 B 0.02996f
C415 VP.n24 B 0.042054f
C416 VP.n25 B 0.295865f
C417 VP.n26 B 0.042054f
C418 VP.n27 B 0.050835f
C419 VP.n28 B 0.02996f
C420 VP.n29 B 0.02996f
C421 VP.n30 B 0.02996f
C422 VP.n31 B 0.051427f
C423 VP.n32 B 0.295865f
C424 VP.n33 B 0.032681f
C425 VP.n34 B 0.059693f
C426 VP.n35 B 0.02996f
C427 VP.n36 B 0.02996f
C428 VP.n37 B 0.02996f
C429 VP.n38 B 0.059392f
C430 VP.n39 B 0.033232f
C431 VP.n40 B 0.366611f
C432 VP.n41 B 1.33189f
C433 VP.n42 B 1.3565f
C434 VP.n43 B 0.02996f
C435 VP.n44 B 0.033232f
C436 VP.n45 B 0.059392f
C437 VP.n46 B 0.024231f
C438 VP.n47 B 0.02996f
C439 VP.n48 B 0.02996f
C440 VP.n49 B 0.02996f
C441 VP.n50 B 0.032681f
C442 VP.n51 B 0.295865f
C443 VP.n52 B 0.051427f
C444 VP.n53 B 0.036643f
C445 VP.n54 B 0.02996f
C446 VP.n55 B 0.02996f
C447 VP.n56 B 0.02996f
C448 VP.n57 B 0.042054f
C449 VP.n58 B 0.295865f
C450 VP.n59 B 0.042054f
C451 VP.n60 B 0.050835f
C452 VP.n61 B 0.02996f
C453 VP.n62 B 0.02996f
C454 VP.n63 B 0.02996f
C455 VP.n64 B 0.051427f
C456 VP.n65 B 0.295865f
C457 VP.n66 B 0.032681f
C458 VP.n67 B 0.059693f
C459 VP.n68 B 0.02996f
C460 VP.n69 B 0.02996f
C461 VP.n70 B 0.02996f
C462 VP.n71 B 0.059392f
C463 VP.n72 B 0.033232f
C464 VP.n73 B 0.366611f
C465 VP.n74 B 0.032017f
.ends

