* NGSPICE file created from diff_pair_sample_1086.ext - technology: sky130A

.subckt diff_pair_sample_1086 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t3 w_n3514_n2012# sky130_fd_pr__pfet_01v8 ad=0.8613 pd=5.55 as=0.8613 ps=5.55 w=5.22 l=2.85
X1 VDD1.t1 VP.t1 VTAIL.t10 w_n3514_n2012# sky130_fd_pr__pfet_01v8 ad=0.8613 pd=5.55 as=2.0358 ps=11.22 w=5.22 l=2.85
X2 VDD1.t2 VP.t2 VTAIL.t9 w_n3514_n2012# sky130_fd_pr__pfet_01v8 ad=0.8613 pd=5.55 as=2.0358 ps=11.22 w=5.22 l=2.85
X3 VDD2.t5 VN.t0 VTAIL.t0 w_n3514_n2012# sky130_fd_pr__pfet_01v8 ad=0.8613 pd=5.55 as=2.0358 ps=11.22 w=5.22 l=2.85
X4 B.t11 B.t9 B.t10 w_n3514_n2012# sky130_fd_pr__pfet_01v8 ad=2.0358 pd=11.22 as=0 ps=0 w=5.22 l=2.85
X5 B.t8 B.t6 B.t7 w_n3514_n2012# sky130_fd_pr__pfet_01v8 ad=2.0358 pd=11.22 as=0 ps=0 w=5.22 l=2.85
X6 VDD1.t0 VP.t3 VTAIL.t8 w_n3514_n2012# sky130_fd_pr__pfet_01v8 ad=2.0358 pd=11.22 as=0.8613 ps=5.55 w=5.22 l=2.85
X7 VDD2.t4 VN.t1 VTAIL.t5 w_n3514_n2012# sky130_fd_pr__pfet_01v8 ad=0.8613 pd=5.55 as=2.0358 ps=11.22 w=5.22 l=2.85
X8 VTAIL.t1 VN.t2 VDD2.t3 w_n3514_n2012# sky130_fd_pr__pfet_01v8 ad=0.8613 pd=5.55 as=0.8613 ps=5.55 w=5.22 l=2.85
X9 B.t5 B.t3 B.t4 w_n3514_n2012# sky130_fd_pr__pfet_01v8 ad=2.0358 pd=11.22 as=0 ps=0 w=5.22 l=2.85
X10 VDD2.t2 VN.t3 VTAIL.t4 w_n3514_n2012# sky130_fd_pr__pfet_01v8 ad=2.0358 pd=11.22 as=0.8613 ps=5.55 w=5.22 l=2.85
X11 B.t2 B.t0 B.t1 w_n3514_n2012# sky130_fd_pr__pfet_01v8 ad=2.0358 pd=11.22 as=0 ps=0 w=5.22 l=2.85
X12 VTAIL.t7 VP.t4 VDD1.t4 w_n3514_n2012# sky130_fd_pr__pfet_01v8 ad=0.8613 pd=5.55 as=0.8613 ps=5.55 w=5.22 l=2.85
X13 VDD2.t1 VN.t4 VTAIL.t3 w_n3514_n2012# sky130_fd_pr__pfet_01v8 ad=2.0358 pd=11.22 as=0.8613 ps=5.55 w=5.22 l=2.85
X14 VDD1.t5 VP.t5 VTAIL.t6 w_n3514_n2012# sky130_fd_pr__pfet_01v8 ad=2.0358 pd=11.22 as=0.8613 ps=5.55 w=5.22 l=2.85
X15 VTAIL.t2 VN.t5 VDD2.t0 w_n3514_n2012# sky130_fd_pr__pfet_01v8 ad=0.8613 pd=5.55 as=0.8613 ps=5.55 w=5.22 l=2.85
R0 VP.n13 VP.n10 161.3
R1 VP.n15 VP.n14 161.3
R2 VP.n16 VP.n9 161.3
R3 VP.n18 VP.n17 161.3
R4 VP.n19 VP.n8 161.3
R5 VP.n21 VP.n20 161.3
R6 VP.n43 VP.n42 161.3
R7 VP.n41 VP.n1 161.3
R8 VP.n40 VP.n39 161.3
R9 VP.n38 VP.n2 161.3
R10 VP.n37 VP.n36 161.3
R11 VP.n35 VP.n3 161.3
R12 VP.n33 VP.n32 161.3
R13 VP.n31 VP.n4 161.3
R14 VP.n30 VP.n29 161.3
R15 VP.n28 VP.n5 161.3
R16 VP.n27 VP.n26 161.3
R17 VP.n25 VP.n6 161.3
R18 VP.n11 VP.t3 75.972
R19 VP.n24 VP.n23 69.0966
R20 VP.n44 VP.n0 69.0966
R21 VP.n22 VP.n7 69.0966
R22 VP.n12 VP.n11 61.6484
R23 VP.n29 VP.n28 56.0773
R24 VP.n40 VP.n2 56.0773
R25 VP.n18 VP.n9 56.0773
R26 VP.n24 VP.n22 44.6208
R27 VP.n23 VP.t5 44.1416
R28 VP.n34 VP.t0 44.1416
R29 VP.n0 VP.t1 44.1416
R30 VP.n7 VP.t2 44.1416
R31 VP.n12 VP.t4 44.1416
R32 VP.n28 VP.n27 25.0767
R33 VP.n41 VP.n40 25.0767
R34 VP.n19 VP.n18 25.0767
R35 VP.n27 VP.n6 24.5923
R36 VP.n29 VP.n4 24.5923
R37 VP.n33 VP.n4 24.5923
R38 VP.n36 VP.n35 24.5923
R39 VP.n36 VP.n2 24.5923
R40 VP.n42 VP.n41 24.5923
R41 VP.n20 VP.n19 24.5923
R42 VP.n14 VP.n13 24.5923
R43 VP.n14 VP.n9 24.5923
R44 VP.n23 VP.n6 21.1495
R45 VP.n42 VP.n0 21.1495
R46 VP.n20 VP.n7 21.1495
R47 VP.n34 VP.n33 12.2964
R48 VP.n35 VP.n34 12.2964
R49 VP.n13 VP.n12 12.2964
R50 VP.n11 VP.n10 5.45928
R51 VP.n22 VP.n21 0.354861
R52 VP.n25 VP.n24 0.354861
R53 VP.n44 VP.n43 0.354861
R54 VP VP.n44 0.267071
R55 VP.n15 VP.n10 0.189894
R56 VP.n16 VP.n15 0.189894
R57 VP.n17 VP.n16 0.189894
R58 VP.n17 VP.n8 0.189894
R59 VP.n21 VP.n8 0.189894
R60 VP.n26 VP.n25 0.189894
R61 VP.n26 VP.n5 0.189894
R62 VP.n30 VP.n5 0.189894
R63 VP.n31 VP.n30 0.189894
R64 VP.n32 VP.n31 0.189894
R65 VP.n32 VP.n3 0.189894
R66 VP.n37 VP.n3 0.189894
R67 VP.n38 VP.n37 0.189894
R68 VP.n39 VP.n38 0.189894
R69 VP.n39 VP.n1 0.189894
R70 VP.n43 VP.n1 0.189894
R71 VDD1.n22 VDD1.n0 756.745
R72 VDD1.n49 VDD1.n27 756.745
R73 VDD1.n23 VDD1.n22 585
R74 VDD1.n21 VDD1.n20 585
R75 VDD1.n4 VDD1.n3 585
R76 VDD1.n15 VDD1.n14 585
R77 VDD1.n13 VDD1.n12 585
R78 VDD1.n8 VDD1.n7 585
R79 VDD1.n35 VDD1.n34 585
R80 VDD1.n40 VDD1.n39 585
R81 VDD1.n42 VDD1.n41 585
R82 VDD1.n31 VDD1.n30 585
R83 VDD1.n48 VDD1.n47 585
R84 VDD1.n50 VDD1.n49 585
R85 VDD1.n9 VDD1.t0 327.856
R86 VDD1.n36 VDD1.t5 327.856
R87 VDD1.n22 VDD1.n21 171.744
R88 VDD1.n21 VDD1.n3 171.744
R89 VDD1.n14 VDD1.n3 171.744
R90 VDD1.n14 VDD1.n13 171.744
R91 VDD1.n13 VDD1.n7 171.744
R92 VDD1.n40 VDD1.n34 171.744
R93 VDD1.n41 VDD1.n40 171.744
R94 VDD1.n41 VDD1.n30 171.744
R95 VDD1.n48 VDD1.n30 171.744
R96 VDD1.n49 VDD1.n48 171.744
R97 VDD1.n55 VDD1.n54 96.7971
R98 VDD1.n57 VDD1.n56 96.1671
R99 VDD1.t0 VDD1.n7 85.8723
R100 VDD1.t5 VDD1.n34 85.8723
R101 VDD1 VDD1.n26 49.8147
R102 VDD1.n55 VDD1.n53 49.7012
R103 VDD1.n57 VDD1.n55 39.0785
R104 VDD1.n9 VDD1.n8 16.381
R105 VDD1.n36 VDD1.n35 16.381
R106 VDD1.n12 VDD1.n11 12.8005
R107 VDD1.n39 VDD1.n38 12.8005
R108 VDD1.n15 VDD1.n6 12.0247
R109 VDD1.n42 VDD1.n33 12.0247
R110 VDD1.n16 VDD1.n4 11.249
R111 VDD1.n43 VDD1.n31 11.249
R112 VDD1.n20 VDD1.n19 10.4732
R113 VDD1.n47 VDD1.n46 10.4732
R114 VDD1.n23 VDD1.n2 9.69747
R115 VDD1.n50 VDD1.n29 9.69747
R116 VDD1.n26 VDD1.n25 9.45567
R117 VDD1.n53 VDD1.n52 9.45567
R118 VDD1.n25 VDD1.n24 9.3005
R119 VDD1.n2 VDD1.n1 9.3005
R120 VDD1.n19 VDD1.n18 9.3005
R121 VDD1.n17 VDD1.n16 9.3005
R122 VDD1.n6 VDD1.n5 9.3005
R123 VDD1.n11 VDD1.n10 9.3005
R124 VDD1.n52 VDD1.n51 9.3005
R125 VDD1.n29 VDD1.n28 9.3005
R126 VDD1.n46 VDD1.n45 9.3005
R127 VDD1.n44 VDD1.n43 9.3005
R128 VDD1.n33 VDD1.n32 9.3005
R129 VDD1.n38 VDD1.n37 9.3005
R130 VDD1.n24 VDD1.n0 8.92171
R131 VDD1.n51 VDD1.n27 8.92171
R132 VDD1.n56 VDD1.t4 6.22751
R133 VDD1.n56 VDD1.t2 6.22751
R134 VDD1.n54 VDD1.t3 6.22751
R135 VDD1.n54 VDD1.t1 6.22751
R136 VDD1.n26 VDD1.n0 5.04292
R137 VDD1.n53 VDD1.n27 5.04292
R138 VDD1.n24 VDD1.n23 4.26717
R139 VDD1.n51 VDD1.n50 4.26717
R140 VDD1.n10 VDD1.n9 3.71853
R141 VDD1.n37 VDD1.n36 3.71853
R142 VDD1.n20 VDD1.n2 3.49141
R143 VDD1.n47 VDD1.n29 3.49141
R144 VDD1.n19 VDD1.n4 2.71565
R145 VDD1.n46 VDD1.n31 2.71565
R146 VDD1.n16 VDD1.n15 1.93989
R147 VDD1.n43 VDD1.n42 1.93989
R148 VDD1.n12 VDD1.n6 1.16414
R149 VDD1.n39 VDD1.n33 1.16414
R150 VDD1 VDD1.n57 0.627655
R151 VDD1.n11 VDD1.n8 0.388379
R152 VDD1.n38 VDD1.n35 0.388379
R153 VDD1.n25 VDD1.n1 0.155672
R154 VDD1.n18 VDD1.n1 0.155672
R155 VDD1.n18 VDD1.n17 0.155672
R156 VDD1.n17 VDD1.n5 0.155672
R157 VDD1.n10 VDD1.n5 0.155672
R158 VDD1.n37 VDD1.n32 0.155672
R159 VDD1.n44 VDD1.n32 0.155672
R160 VDD1.n45 VDD1.n44 0.155672
R161 VDD1.n45 VDD1.n28 0.155672
R162 VDD1.n52 VDD1.n28 0.155672
R163 VTAIL.n114 VTAIL.n92 756.745
R164 VTAIL.n24 VTAIL.n2 756.745
R165 VTAIL.n86 VTAIL.n64 756.745
R166 VTAIL.n56 VTAIL.n34 756.745
R167 VTAIL.n100 VTAIL.n99 585
R168 VTAIL.n105 VTAIL.n104 585
R169 VTAIL.n107 VTAIL.n106 585
R170 VTAIL.n96 VTAIL.n95 585
R171 VTAIL.n113 VTAIL.n112 585
R172 VTAIL.n115 VTAIL.n114 585
R173 VTAIL.n10 VTAIL.n9 585
R174 VTAIL.n15 VTAIL.n14 585
R175 VTAIL.n17 VTAIL.n16 585
R176 VTAIL.n6 VTAIL.n5 585
R177 VTAIL.n23 VTAIL.n22 585
R178 VTAIL.n25 VTAIL.n24 585
R179 VTAIL.n87 VTAIL.n86 585
R180 VTAIL.n85 VTAIL.n84 585
R181 VTAIL.n68 VTAIL.n67 585
R182 VTAIL.n79 VTAIL.n78 585
R183 VTAIL.n77 VTAIL.n76 585
R184 VTAIL.n72 VTAIL.n71 585
R185 VTAIL.n57 VTAIL.n56 585
R186 VTAIL.n55 VTAIL.n54 585
R187 VTAIL.n38 VTAIL.n37 585
R188 VTAIL.n49 VTAIL.n48 585
R189 VTAIL.n47 VTAIL.n46 585
R190 VTAIL.n42 VTAIL.n41 585
R191 VTAIL.n101 VTAIL.t0 327.856
R192 VTAIL.n11 VTAIL.t10 327.856
R193 VTAIL.n73 VTAIL.t9 327.856
R194 VTAIL.n43 VTAIL.t5 327.856
R195 VTAIL.n105 VTAIL.n99 171.744
R196 VTAIL.n106 VTAIL.n105 171.744
R197 VTAIL.n106 VTAIL.n95 171.744
R198 VTAIL.n113 VTAIL.n95 171.744
R199 VTAIL.n114 VTAIL.n113 171.744
R200 VTAIL.n15 VTAIL.n9 171.744
R201 VTAIL.n16 VTAIL.n15 171.744
R202 VTAIL.n16 VTAIL.n5 171.744
R203 VTAIL.n23 VTAIL.n5 171.744
R204 VTAIL.n24 VTAIL.n23 171.744
R205 VTAIL.n86 VTAIL.n85 171.744
R206 VTAIL.n85 VTAIL.n67 171.744
R207 VTAIL.n78 VTAIL.n67 171.744
R208 VTAIL.n78 VTAIL.n77 171.744
R209 VTAIL.n77 VTAIL.n71 171.744
R210 VTAIL.n56 VTAIL.n55 171.744
R211 VTAIL.n55 VTAIL.n37 171.744
R212 VTAIL.n48 VTAIL.n37 171.744
R213 VTAIL.n48 VTAIL.n47 171.744
R214 VTAIL.n47 VTAIL.n41 171.744
R215 VTAIL.t0 VTAIL.n99 85.8723
R216 VTAIL.t10 VTAIL.n9 85.8723
R217 VTAIL.t9 VTAIL.n71 85.8723
R218 VTAIL.t5 VTAIL.n41 85.8723
R219 VTAIL.n63 VTAIL.n62 79.4885
R220 VTAIL.n33 VTAIL.n32 79.4885
R221 VTAIL.n1 VTAIL.n0 79.4883
R222 VTAIL.n31 VTAIL.n30 79.4883
R223 VTAIL.n119 VTAIL.n118 31.0217
R224 VTAIL.n29 VTAIL.n28 31.0217
R225 VTAIL.n91 VTAIL.n90 31.0217
R226 VTAIL.n61 VTAIL.n60 31.0217
R227 VTAIL.n33 VTAIL.n31 22.3496
R228 VTAIL.n119 VTAIL.n91 19.6083
R229 VTAIL.n101 VTAIL.n100 16.381
R230 VTAIL.n11 VTAIL.n10 16.381
R231 VTAIL.n73 VTAIL.n72 16.381
R232 VTAIL.n43 VTAIL.n42 16.381
R233 VTAIL.n104 VTAIL.n103 12.8005
R234 VTAIL.n14 VTAIL.n13 12.8005
R235 VTAIL.n76 VTAIL.n75 12.8005
R236 VTAIL.n46 VTAIL.n45 12.8005
R237 VTAIL.n107 VTAIL.n98 12.0247
R238 VTAIL.n17 VTAIL.n8 12.0247
R239 VTAIL.n79 VTAIL.n70 12.0247
R240 VTAIL.n49 VTAIL.n40 12.0247
R241 VTAIL.n108 VTAIL.n96 11.249
R242 VTAIL.n18 VTAIL.n6 11.249
R243 VTAIL.n80 VTAIL.n68 11.249
R244 VTAIL.n50 VTAIL.n38 11.249
R245 VTAIL.n112 VTAIL.n111 10.4732
R246 VTAIL.n22 VTAIL.n21 10.4732
R247 VTAIL.n84 VTAIL.n83 10.4732
R248 VTAIL.n54 VTAIL.n53 10.4732
R249 VTAIL.n115 VTAIL.n94 9.69747
R250 VTAIL.n25 VTAIL.n4 9.69747
R251 VTAIL.n87 VTAIL.n66 9.69747
R252 VTAIL.n57 VTAIL.n36 9.69747
R253 VTAIL.n118 VTAIL.n117 9.45567
R254 VTAIL.n28 VTAIL.n27 9.45567
R255 VTAIL.n90 VTAIL.n89 9.45567
R256 VTAIL.n60 VTAIL.n59 9.45567
R257 VTAIL.n117 VTAIL.n116 9.3005
R258 VTAIL.n94 VTAIL.n93 9.3005
R259 VTAIL.n111 VTAIL.n110 9.3005
R260 VTAIL.n109 VTAIL.n108 9.3005
R261 VTAIL.n98 VTAIL.n97 9.3005
R262 VTAIL.n103 VTAIL.n102 9.3005
R263 VTAIL.n27 VTAIL.n26 9.3005
R264 VTAIL.n4 VTAIL.n3 9.3005
R265 VTAIL.n21 VTAIL.n20 9.3005
R266 VTAIL.n19 VTAIL.n18 9.3005
R267 VTAIL.n8 VTAIL.n7 9.3005
R268 VTAIL.n13 VTAIL.n12 9.3005
R269 VTAIL.n89 VTAIL.n88 9.3005
R270 VTAIL.n66 VTAIL.n65 9.3005
R271 VTAIL.n83 VTAIL.n82 9.3005
R272 VTAIL.n81 VTAIL.n80 9.3005
R273 VTAIL.n70 VTAIL.n69 9.3005
R274 VTAIL.n75 VTAIL.n74 9.3005
R275 VTAIL.n59 VTAIL.n58 9.3005
R276 VTAIL.n36 VTAIL.n35 9.3005
R277 VTAIL.n53 VTAIL.n52 9.3005
R278 VTAIL.n51 VTAIL.n50 9.3005
R279 VTAIL.n40 VTAIL.n39 9.3005
R280 VTAIL.n45 VTAIL.n44 9.3005
R281 VTAIL.n116 VTAIL.n92 8.92171
R282 VTAIL.n26 VTAIL.n2 8.92171
R283 VTAIL.n88 VTAIL.n64 8.92171
R284 VTAIL.n58 VTAIL.n34 8.92171
R285 VTAIL.n0 VTAIL.t4 6.22751
R286 VTAIL.n0 VTAIL.t1 6.22751
R287 VTAIL.n30 VTAIL.t6 6.22751
R288 VTAIL.n30 VTAIL.t11 6.22751
R289 VTAIL.n62 VTAIL.t8 6.22751
R290 VTAIL.n62 VTAIL.t7 6.22751
R291 VTAIL.n32 VTAIL.t3 6.22751
R292 VTAIL.n32 VTAIL.t2 6.22751
R293 VTAIL.n118 VTAIL.n92 5.04292
R294 VTAIL.n28 VTAIL.n2 5.04292
R295 VTAIL.n90 VTAIL.n64 5.04292
R296 VTAIL.n60 VTAIL.n34 5.04292
R297 VTAIL.n116 VTAIL.n115 4.26717
R298 VTAIL.n26 VTAIL.n25 4.26717
R299 VTAIL.n88 VTAIL.n87 4.26717
R300 VTAIL.n58 VTAIL.n57 4.26717
R301 VTAIL.n74 VTAIL.n73 3.71853
R302 VTAIL.n44 VTAIL.n43 3.71853
R303 VTAIL.n102 VTAIL.n101 3.71853
R304 VTAIL.n12 VTAIL.n11 3.71853
R305 VTAIL.n112 VTAIL.n94 3.49141
R306 VTAIL.n22 VTAIL.n4 3.49141
R307 VTAIL.n84 VTAIL.n66 3.49141
R308 VTAIL.n54 VTAIL.n36 3.49141
R309 VTAIL.n61 VTAIL.n33 2.74188
R310 VTAIL.n91 VTAIL.n63 2.74188
R311 VTAIL.n31 VTAIL.n29 2.74188
R312 VTAIL.n111 VTAIL.n96 2.71565
R313 VTAIL.n21 VTAIL.n6 2.71565
R314 VTAIL.n83 VTAIL.n68 2.71565
R315 VTAIL.n53 VTAIL.n38 2.71565
R316 VTAIL VTAIL.n119 1.99834
R317 VTAIL.n108 VTAIL.n107 1.93989
R318 VTAIL.n18 VTAIL.n17 1.93989
R319 VTAIL.n80 VTAIL.n79 1.93989
R320 VTAIL.n50 VTAIL.n49 1.93989
R321 VTAIL.n63 VTAIL.n61 1.84102
R322 VTAIL.n29 VTAIL.n1 1.84102
R323 VTAIL.n104 VTAIL.n98 1.16414
R324 VTAIL.n14 VTAIL.n8 1.16414
R325 VTAIL.n76 VTAIL.n70 1.16414
R326 VTAIL.n46 VTAIL.n40 1.16414
R327 VTAIL VTAIL.n1 0.744035
R328 VTAIL.n103 VTAIL.n100 0.388379
R329 VTAIL.n13 VTAIL.n10 0.388379
R330 VTAIL.n75 VTAIL.n72 0.388379
R331 VTAIL.n45 VTAIL.n42 0.388379
R332 VTAIL.n102 VTAIL.n97 0.155672
R333 VTAIL.n109 VTAIL.n97 0.155672
R334 VTAIL.n110 VTAIL.n109 0.155672
R335 VTAIL.n110 VTAIL.n93 0.155672
R336 VTAIL.n117 VTAIL.n93 0.155672
R337 VTAIL.n12 VTAIL.n7 0.155672
R338 VTAIL.n19 VTAIL.n7 0.155672
R339 VTAIL.n20 VTAIL.n19 0.155672
R340 VTAIL.n20 VTAIL.n3 0.155672
R341 VTAIL.n27 VTAIL.n3 0.155672
R342 VTAIL.n89 VTAIL.n65 0.155672
R343 VTAIL.n82 VTAIL.n65 0.155672
R344 VTAIL.n82 VTAIL.n81 0.155672
R345 VTAIL.n81 VTAIL.n69 0.155672
R346 VTAIL.n74 VTAIL.n69 0.155672
R347 VTAIL.n59 VTAIL.n35 0.155672
R348 VTAIL.n52 VTAIL.n35 0.155672
R349 VTAIL.n52 VTAIL.n51 0.155672
R350 VTAIL.n51 VTAIL.n39 0.155672
R351 VTAIL.n44 VTAIL.n39 0.155672
R352 VN.n30 VN.n29 161.3
R353 VN.n28 VN.n17 161.3
R354 VN.n27 VN.n26 161.3
R355 VN.n25 VN.n18 161.3
R356 VN.n24 VN.n23 161.3
R357 VN.n22 VN.n19 161.3
R358 VN.n14 VN.n13 161.3
R359 VN.n12 VN.n1 161.3
R360 VN.n11 VN.n10 161.3
R361 VN.n9 VN.n2 161.3
R362 VN.n8 VN.n7 161.3
R363 VN.n6 VN.n3 161.3
R364 VN.n20 VN.t1 75.9722
R365 VN.n4 VN.t3 75.9722
R366 VN.n15 VN.n0 69.0966
R367 VN.n31 VN.n16 69.0966
R368 VN.n5 VN.n4 61.6484
R369 VN.n21 VN.n20 61.6484
R370 VN.n11 VN.n2 56.0773
R371 VN.n27 VN.n18 56.0773
R372 VN VN.n31 44.786
R373 VN.n5 VN.t2 44.1416
R374 VN.n0 VN.t0 44.1416
R375 VN.n21 VN.t5 44.1416
R376 VN.n16 VN.t4 44.1416
R377 VN.n12 VN.n11 25.0767
R378 VN.n28 VN.n27 25.0767
R379 VN.n7 VN.n6 24.5923
R380 VN.n7 VN.n2 24.5923
R381 VN.n13 VN.n12 24.5923
R382 VN.n23 VN.n18 24.5923
R383 VN.n23 VN.n22 24.5923
R384 VN.n29 VN.n28 24.5923
R385 VN.n13 VN.n0 21.1495
R386 VN.n29 VN.n16 21.1495
R387 VN.n6 VN.n5 12.2964
R388 VN.n22 VN.n21 12.2964
R389 VN.n20 VN.n19 5.45931
R390 VN.n4 VN.n3 5.45931
R391 VN.n31 VN.n30 0.354861
R392 VN.n15 VN.n14 0.354861
R393 VN VN.n15 0.267071
R394 VN.n30 VN.n17 0.189894
R395 VN.n26 VN.n17 0.189894
R396 VN.n26 VN.n25 0.189894
R397 VN.n25 VN.n24 0.189894
R398 VN.n24 VN.n19 0.189894
R399 VN.n8 VN.n3 0.189894
R400 VN.n9 VN.n8 0.189894
R401 VN.n10 VN.n9 0.189894
R402 VN.n10 VN.n1 0.189894
R403 VN.n14 VN.n1 0.189894
R404 VDD2.n51 VDD2.n29 756.745
R405 VDD2.n22 VDD2.n0 756.745
R406 VDD2.n52 VDD2.n51 585
R407 VDD2.n50 VDD2.n49 585
R408 VDD2.n33 VDD2.n32 585
R409 VDD2.n44 VDD2.n43 585
R410 VDD2.n42 VDD2.n41 585
R411 VDD2.n37 VDD2.n36 585
R412 VDD2.n8 VDD2.n7 585
R413 VDD2.n13 VDD2.n12 585
R414 VDD2.n15 VDD2.n14 585
R415 VDD2.n4 VDD2.n3 585
R416 VDD2.n21 VDD2.n20 585
R417 VDD2.n23 VDD2.n22 585
R418 VDD2.n38 VDD2.t1 327.856
R419 VDD2.n9 VDD2.t2 327.856
R420 VDD2.n51 VDD2.n50 171.744
R421 VDD2.n50 VDD2.n32 171.744
R422 VDD2.n43 VDD2.n32 171.744
R423 VDD2.n43 VDD2.n42 171.744
R424 VDD2.n42 VDD2.n36 171.744
R425 VDD2.n13 VDD2.n7 171.744
R426 VDD2.n14 VDD2.n13 171.744
R427 VDD2.n14 VDD2.n3 171.744
R428 VDD2.n21 VDD2.n3 171.744
R429 VDD2.n22 VDD2.n21 171.744
R430 VDD2.n28 VDD2.n27 96.7971
R431 VDD2 VDD2.n57 96.7943
R432 VDD2.t1 VDD2.n36 85.8723
R433 VDD2.t2 VDD2.n7 85.8723
R434 VDD2.n28 VDD2.n26 49.7012
R435 VDD2.n56 VDD2.n55 47.7005
R436 VDD2.n56 VDD2.n28 37.1248
R437 VDD2.n38 VDD2.n37 16.381
R438 VDD2.n9 VDD2.n8 16.381
R439 VDD2.n41 VDD2.n40 12.8005
R440 VDD2.n12 VDD2.n11 12.8005
R441 VDD2.n44 VDD2.n35 12.0247
R442 VDD2.n15 VDD2.n6 12.0247
R443 VDD2.n45 VDD2.n33 11.249
R444 VDD2.n16 VDD2.n4 11.249
R445 VDD2.n49 VDD2.n48 10.4732
R446 VDD2.n20 VDD2.n19 10.4732
R447 VDD2.n52 VDD2.n31 9.69747
R448 VDD2.n23 VDD2.n2 9.69747
R449 VDD2.n55 VDD2.n54 9.45567
R450 VDD2.n26 VDD2.n25 9.45567
R451 VDD2.n54 VDD2.n53 9.3005
R452 VDD2.n31 VDD2.n30 9.3005
R453 VDD2.n48 VDD2.n47 9.3005
R454 VDD2.n46 VDD2.n45 9.3005
R455 VDD2.n35 VDD2.n34 9.3005
R456 VDD2.n40 VDD2.n39 9.3005
R457 VDD2.n25 VDD2.n24 9.3005
R458 VDD2.n2 VDD2.n1 9.3005
R459 VDD2.n19 VDD2.n18 9.3005
R460 VDD2.n17 VDD2.n16 9.3005
R461 VDD2.n6 VDD2.n5 9.3005
R462 VDD2.n11 VDD2.n10 9.3005
R463 VDD2.n53 VDD2.n29 8.92171
R464 VDD2.n24 VDD2.n0 8.92171
R465 VDD2.n57 VDD2.t0 6.22751
R466 VDD2.n57 VDD2.t4 6.22751
R467 VDD2.n27 VDD2.t3 6.22751
R468 VDD2.n27 VDD2.t5 6.22751
R469 VDD2.n55 VDD2.n29 5.04292
R470 VDD2.n26 VDD2.n0 5.04292
R471 VDD2.n53 VDD2.n52 4.26717
R472 VDD2.n24 VDD2.n23 4.26717
R473 VDD2.n39 VDD2.n38 3.71853
R474 VDD2.n10 VDD2.n9 3.71853
R475 VDD2.n49 VDD2.n31 3.49141
R476 VDD2.n20 VDD2.n2 3.49141
R477 VDD2.n48 VDD2.n33 2.71565
R478 VDD2.n19 VDD2.n4 2.71565
R479 VDD2 VDD2.n56 2.11472
R480 VDD2.n45 VDD2.n44 1.93989
R481 VDD2.n16 VDD2.n15 1.93989
R482 VDD2.n41 VDD2.n35 1.16414
R483 VDD2.n12 VDD2.n6 1.16414
R484 VDD2.n40 VDD2.n37 0.388379
R485 VDD2.n11 VDD2.n8 0.388379
R486 VDD2.n54 VDD2.n30 0.155672
R487 VDD2.n47 VDD2.n30 0.155672
R488 VDD2.n47 VDD2.n46 0.155672
R489 VDD2.n46 VDD2.n34 0.155672
R490 VDD2.n39 VDD2.n34 0.155672
R491 VDD2.n10 VDD2.n5 0.155672
R492 VDD2.n17 VDD2.n5 0.155672
R493 VDD2.n18 VDD2.n17 0.155672
R494 VDD2.n18 VDD2.n1 0.155672
R495 VDD2.n25 VDD2.n1 0.155672
R496 B.n301 B.n300 585
R497 B.n299 B.n102 585
R498 B.n298 B.n297 585
R499 B.n296 B.n103 585
R500 B.n295 B.n294 585
R501 B.n293 B.n104 585
R502 B.n292 B.n291 585
R503 B.n290 B.n105 585
R504 B.n289 B.n288 585
R505 B.n287 B.n106 585
R506 B.n286 B.n285 585
R507 B.n284 B.n107 585
R508 B.n283 B.n282 585
R509 B.n281 B.n108 585
R510 B.n280 B.n279 585
R511 B.n278 B.n109 585
R512 B.n277 B.n276 585
R513 B.n275 B.n110 585
R514 B.n274 B.n273 585
R515 B.n272 B.n111 585
R516 B.n271 B.n270 585
R517 B.n269 B.n112 585
R518 B.n268 B.n267 585
R519 B.n263 B.n113 585
R520 B.n262 B.n261 585
R521 B.n260 B.n114 585
R522 B.n259 B.n258 585
R523 B.n257 B.n115 585
R524 B.n256 B.n255 585
R525 B.n254 B.n116 585
R526 B.n253 B.n252 585
R527 B.n250 B.n117 585
R528 B.n249 B.n248 585
R529 B.n247 B.n120 585
R530 B.n246 B.n245 585
R531 B.n244 B.n121 585
R532 B.n243 B.n242 585
R533 B.n241 B.n122 585
R534 B.n240 B.n239 585
R535 B.n238 B.n123 585
R536 B.n237 B.n236 585
R537 B.n235 B.n124 585
R538 B.n234 B.n233 585
R539 B.n232 B.n125 585
R540 B.n231 B.n230 585
R541 B.n229 B.n126 585
R542 B.n228 B.n227 585
R543 B.n226 B.n127 585
R544 B.n225 B.n224 585
R545 B.n223 B.n128 585
R546 B.n222 B.n221 585
R547 B.n220 B.n129 585
R548 B.n219 B.n218 585
R549 B.n302 B.n101 585
R550 B.n304 B.n303 585
R551 B.n305 B.n100 585
R552 B.n307 B.n306 585
R553 B.n308 B.n99 585
R554 B.n310 B.n309 585
R555 B.n311 B.n98 585
R556 B.n313 B.n312 585
R557 B.n314 B.n97 585
R558 B.n316 B.n315 585
R559 B.n317 B.n96 585
R560 B.n319 B.n318 585
R561 B.n320 B.n95 585
R562 B.n322 B.n321 585
R563 B.n323 B.n94 585
R564 B.n325 B.n324 585
R565 B.n326 B.n93 585
R566 B.n328 B.n327 585
R567 B.n329 B.n92 585
R568 B.n331 B.n330 585
R569 B.n332 B.n91 585
R570 B.n334 B.n333 585
R571 B.n335 B.n90 585
R572 B.n337 B.n336 585
R573 B.n338 B.n89 585
R574 B.n340 B.n339 585
R575 B.n341 B.n88 585
R576 B.n343 B.n342 585
R577 B.n344 B.n87 585
R578 B.n346 B.n345 585
R579 B.n347 B.n86 585
R580 B.n349 B.n348 585
R581 B.n350 B.n85 585
R582 B.n352 B.n351 585
R583 B.n353 B.n84 585
R584 B.n355 B.n354 585
R585 B.n356 B.n83 585
R586 B.n358 B.n357 585
R587 B.n359 B.n82 585
R588 B.n361 B.n360 585
R589 B.n362 B.n81 585
R590 B.n364 B.n363 585
R591 B.n365 B.n80 585
R592 B.n367 B.n366 585
R593 B.n368 B.n79 585
R594 B.n370 B.n369 585
R595 B.n371 B.n78 585
R596 B.n373 B.n372 585
R597 B.n374 B.n77 585
R598 B.n376 B.n375 585
R599 B.n377 B.n76 585
R600 B.n379 B.n378 585
R601 B.n380 B.n75 585
R602 B.n382 B.n381 585
R603 B.n383 B.n74 585
R604 B.n385 B.n384 585
R605 B.n386 B.n73 585
R606 B.n388 B.n387 585
R607 B.n389 B.n72 585
R608 B.n391 B.n390 585
R609 B.n392 B.n71 585
R610 B.n394 B.n393 585
R611 B.n395 B.n70 585
R612 B.n397 B.n396 585
R613 B.n398 B.n69 585
R614 B.n400 B.n399 585
R615 B.n401 B.n68 585
R616 B.n403 B.n402 585
R617 B.n404 B.n67 585
R618 B.n406 B.n405 585
R619 B.n407 B.n66 585
R620 B.n409 B.n408 585
R621 B.n410 B.n65 585
R622 B.n412 B.n411 585
R623 B.n413 B.n64 585
R624 B.n415 B.n414 585
R625 B.n416 B.n63 585
R626 B.n418 B.n417 585
R627 B.n419 B.n62 585
R628 B.n421 B.n420 585
R629 B.n422 B.n61 585
R630 B.n424 B.n423 585
R631 B.n425 B.n60 585
R632 B.n427 B.n426 585
R633 B.n428 B.n59 585
R634 B.n430 B.n429 585
R635 B.n431 B.n58 585
R636 B.n433 B.n432 585
R637 B.n434 B.n57 585
R638 B.n436 B.n435 585
R639 B.n437 B.n56 585
R640 B.n439 B.n438 585
R641 B.n520 B.n519 585
R642 B.n518 B.n25 585
R643 B.n517 B.n516 585
R644 B.n515 B.n26 585
R645 B.n514 B.n513 585
R646 B.n512 B.n27 585
R647 B.n511 B.n510 585
R648 B.n509 B.n28 585
R649 B.n508 B.n507 585
R650 B.n506 B.n29 585
R651 B.n505 B.n504 585
R652 B.n503 B.n30 585
R653 B.n502 B.n501 585
R654 B.n500 B.n31 585
R655 B.n499 B.n498 585
R656 B.n497 B.n32 585
R657 B.n496 B.n495 585
R658 B.n494 B.n33 585
R659 B.n493 B.n492 585
R660 B.n491 B.n34 585
R661 B.n490 B.n489 585
R662 B.n488 B.n35 585
R663 B.n486 B.n485 585
R664 B.n484 B.n38 585
R665 B.n483 B.n482 585
R666 B.n481 B.n39 585
R667 B.n480 B.n479 585
R668 B.n478 B.n40 585
R669 B.n477 B.n476 585
R670 B.n475 B.n41 585
R671 B.n474 B.n473 585
R672 B.n472 B.n471 585
R673 B.n470 B.n45 585
R674 B.n469 B.n468 585
R675 B.n467 B.n46 585
R676 B.n466 B.n465 585
R677 B.n464 B.n47 585
R678 B.n463 B.n462 585
R679 B.n461 B.n48 585
R680 B.n460 B.n459 585
R681 B.n458 B.n49 585
R682 B.n457 B.n456 585
R683 B.n455 B.n50 585
R684 B.n454 B.n453 585
R685 B.n452 B.n51 585
R686 B.n451 B.n450 585
R687 B.n449 B.n52 585
R688 B.n448 B.n447 585
R689 B.n446 B.n53 585
R690 B.n445 B.n444 585
R691 B.n443 B.n54 585
R692 B.n442 B.n441 585
R693 B.n440 B.n55 585
R694 B.n521 B.n24 585
R695 B.n523 B.n522 585
R696 B.n524 B.n23 585
R697 B.n526 B.n525 585
R698 B.n527 B.n22 585
R699 B.n529 B.n528 585
R700 B.n530 B.n21 585
R701 B.n532 B.n531 585
R702 B.n533 B.n20 585
R703 B.n535 B.n534 585
R704 B.n536 B.n19 585
R705 B.n538 B.n537 585
R706 B.n539 B.n18 585
R707 B.n541 B.n540 585
R708 B.n542 B.n17 585
R709 B.n544 B.n543 585
R710 B.n545 B.n16 585
R711 B.n547 B.n546 585
R712 B.n548 B.n15 585
R713 B.n550 B.n549 585
R714 B.n551 B.n14 585
R715 B.n553 B.n552 585
R716 B.n554 B.n13 585
R717 B.n556 B.n555 585
R718 B.n557 B.n12 585
R719 B.n559 B.n558 585
R720 B.n560 B.n11 585
R721 B.n562 B.n561 585
R722 B.n563 B.n10 585
R723 B.n565 B.n564 585
R724 B.n566 B.n9 585
R725 B.n568 B.n567 585
R726 B.n569 B.n8 585
R727 B.n571 B.n570 585
R728 B.n572 B.n7 585
R729 B.n574 B.n573 585
R730 B.n575 B.n6 585
R731 B.n577 B.n576 585
R732 B.n578 B.n5 585
R733 B.n580 B.n579 585
R734 B.n581 B.n4 585
R735 B.n583 B.n582 585
R736 B.n584 B.n3 585
R737 B.n586 B.n585 585
R738 B.n587 B.n0 585
R739 B.n2 B.n1 585
R740 B.n153 B.n152 585
R741 B.n154 B.n151 585
R742 B.n156 B.n155 585
R743 B.n157 B.n150 585
R744 B.n159 B.n158 585
R745 B.n160 B.n149 585
R746 B.n162 B.n161 585
R747 B.n163 B.n148 585
R748 B.n165 B.n164 585
R749 B.n166 B.n147 585
R750 B.n168 B.n167 585
R751 B.n169 B.n146 585
R752 B.n171 B.n170 585
R753 B.n172 B.n145 585
R754 B.n174 B.n173 585
R755 B.n175 B.n144 585
R756 B.n177 B.n176 585
R757 B.n178 B.n143 585
R758 B.n180 B.n179 585
R759 B.n181 B.n142 585
R760 B.n183 B.n182 585
R761 B.n184 B.n141 585
R762 B.n186 B.n185 585
R763 B.n187 B.n140 585
R764 B.n189 B.n188 585
R765 B.n190 B.n139 585
R766 B.n192 B.n191 585
R767 B.n193 B.n138 585
R768 B.n195 B.n194 585
R769 B.n196 B.n137 585
R770 B.n198 B.n197 585
R771 B.n199 B.n136 585
R772 B.n201 B.n200 585
R773 B.n202 B.n135 585
R774 B.n204 B.n203 585
R775 B.n205 B.n134 585
R776 B.n207 B.n206 585
R777 B.n208 B.n133 585
R778 B.n210 B.n209 585
R779 B.n211 B.n132 585
R780 B.n213 B.n212 585
R781 B.n214 B.n131 585
R782 B.n216 B.n215 585
R783 B.n217 B.n130 585
R784 B.n218 B.n217 497.305
R785 B.n300 B.n101 497.305
R786 B.n438 B.n55 497.305
R787 B.n521 B.n520 497.305
R788 B.n264 B.t7 316.158
R789 B.n42 B.t2 316.158
R790 B.n118 B.t10 316.158
R791 B.n36 B.t5 316.158
R792 B.n589 B.n588 256.663
R793 B.n265 B.t8 254.484
R794 B.n43 B.t1 254.484
R795 B.n119 B.t11 254.484
R796 B.n37 B.t4 254.484
R797 B.n118 B.t9 252.536
R798 B.n264 B.t6 252.536
R799 B.n42 B.t0 252.536
R800 B.n36 B.t3 252.536
R801 B.n588 B.n587 235.042
R802 B.n588 B.n2 235.042
R803 B.n218 B.n129 163.367
R804 B.n222 B.n129 163.367
R805 B.n223 B.n222 163.367
R806 B.n224 B.n223 163.367
R807 B.n224 B.n127 163.367
R808 B.n228 B.n127 163.367
R809 B.n229 B.n228 163.367
R810 B.n230 B.n229 163.367
R811 B.n230 B.n125 163.367
R812 B.n234 B.n125 163.367
R813 B.n235 B.n234 163.367
R814 B.n236 B.n235 163.367
R815 B.n236 B.n123 163.367
R816 B.n240 B.n123 163.367
R817 B.n241 B.n240 163.367
R818 B.n242 B.n241 163.367
R819 B.n242 B.n121 163.367
R820 B.n246 B.n121 163.367
R821 B.n247 B.n246 163.367
R822 B.n248 B.n247 163.367
R823 B.n248 B.n117 163.367
R824 B.n253 B.n117 163.367
R825 B.n254 B.n253 163.367
R826 B.n255 B.n254 163.367
R827 B.n255 B.n115 163.367
R828 B.n259 B.n115 163.367
R829 B.n260 B.n259 163.367
R830 B.n261 B.n260 163.367
R831 B.n261 B.n113 163.367
R832 B.n268 B.n113 163.367
R833 B.n269 B.n268 163.367
R834 B.n270 B.n269 163.367
R835 B.n270 B.n111 163.367
R836 B.n274 B.n111 163.367
R837 B.n275 B.n274 163.367
R838 B.n276 B.n275 163.367
R839 B.n276 B.n109 163.367
R840 B.n280 B.n109 163.367
R841 B.n281 B.n280 163.367
R842 B.n282 B.n281 163.367
R843 B.n282 B.n107 163.367
R844 B.n286 B.n107 163.367
R845 B.n287 B.n286 163.367
R846 B.n288 B.n287 163.367
R847 B.n288 B.n105 163.367
R848 B.n292 B.n105 163.367
R849 B.n293 B.n292 163.367
R850 B.n294 B.n293 163.367
R851 B.n294 B.n103 163.367
R852 B.n298 B.n103 163.367
R853 B.n299 B.n298 163.367
R854 B.n300 B.n299 163.367
R855 B.n438 B.n437 163.367
R856 B.n437 B.n436 163.367
R857 B.n436 B.n57 163.367
R858 B.n432 B.n57 163.367
R859 B.n432 B.n431 163.367
R860 B.n431 B.n430 163.367
R861 B.n430 B.n59 163.367
R862 B.n426 B.n59 163.367
R863 B.n426 B.n425 163.367
R864 B.n425 B.n424 163.367
R865 B.n424 B.n61 163.367
R866 B.n420 B.n61 163.367
R867 B.n420 B.n419 163.367
R868 B.n419 B.n418 163.367
R869 B.n418 B.n63 163.367
R870 B.n414 B.n63 163.367
R871 B.n414 B.n413 163.367
R872 B.n413 B.n412 163.367
R873 B.n412 B.n65 163.367
R874 B.n408 B.n65 163.367
R875 B.n408 B.n407 163.367
R876 B.n407 B.n406 163.367
R877 B.n406 B.n67 163.367
R878 B.n402 B.n67 163.367
R879 B.n402 B.n401 163.367
R880 B.n401 B.n400 163.367
R881 B.n400 B.n69 163.367
R882 B.n396 B.n69 163.367
R883 B.n396 B.n395 163.367
R884 B.n395 B.n394 163.367
R885 B.n394 B.n71 163.367
R886 B.n390 B.n71 163.367
R887 B.n390 B.n389 163.367
R888 B.n389 B.n388 163.367
R889 B.n388 B.n73 163.367
R890 B.n384 B.n73 163.367
R891 B.n384 B.n383 163.367
R892 B.n383 B.n382 163.367
R893 B.n382 B.n75 163.367
R894 B.n378 B.n75 163.367
R895 B.n378 B.n377 163.367
R896 B.n377 B.n376 163.367
R897 B.n376 B.n77 163.367
R898 B.n372 B.n77 163.367
R899 B.n372 B.n371 163.367
R900 B.n371 B.n370 163.367
R901 B.n370 B.n79 163.367
R902 B.n366 B.n79 163.367
R903 B.n366 B.n365 163.367
R904 B.n365 B.n364 163.367
R905 B.n364 B.n81 163.367
R906 B.n360 B.n81 163.367
R907 B.n360 B.n359 163.367
R908 B.n359 B.n358 163.367
R909 B.n358 B.n83 163.367
R910 B.n354 B.n83 163.367
R911 B.n354 B.n353 163.367
R912 B.n353 B.n352 163.367
R913 B.n352 B.n85 163.367
R914 B.n348 B.n85 163.367
R915 B.n348 B.n347 163.367
R916 B.n347 B.n346 163.367
R917 B.n346 B.n87 163.367
R918 B.n342 B.n87 163.367
R919 B.n342 B.n341 163.367
R920 B.n341 B.n340 163.367
R921 B.n340 B.n89 163.367
R922 B.n336 B.n89 163.367
R923 B.n336 B.n335 163.367
R924 B.n335 B.n334 163.367
R925 B.n334 B.n91 163.367
R926 B.n330 B.n91 163.367
R927 B.n330 B.n329 163.367
R928 B.n329 B.n328 163.367
R929 B.n328 B.n93 163.367
R930 B.n324 B.n93 163.367
R931 B.n324 B.n323 163.367
R932 B.n323 B.n322 163.367
R933 B.n322 B.n95 163.367
R934 B.n318 B.n95 163.367
R935 B.n318 B.n317 163.367
R936 B.n317 B.n316 163.367
R937 B.n316 B.n97 163.367
R938 B.n312 B.n97 163.367
R939 B.n312 B.n311 163.367
R940 B.n311 B.n310 163.367
R941 B.n310 B.n99 163.367
R942 B.n306 B.n99 163.367
R943 B.n306 B.n305 163.367
R944 B.n305 B.n304 163.367
R945 B.n304 B.n101 163.367
R946 B.n520 B.n25 163.367
R947 B.n516 B.n25 163.367
R948 B.n516 B.n515 163.367
R949 B.n515 B.n514 163.367
R950 B.n514 B.n27 163.367
R951 B.n510 B.n27 163.367
R952 B.n510 B.n509 163.367
R953 B.n509 B.n508 163.367
R954 B.n508 B.n29 163.367
R955 B.n504 B.n29 163.367
R956 B.n504 B.n503 163.367
R957 B.n503 B.n502 163.367
R958 B.n502 B.n31 163.367
R959 B.n498 B.n31 163.367
R960 B.n498 B.n497 163.367
R961 B.n497 B.n496 163.367
R962 B.n496 B.n33 163.367
R963 B.n492 B.n33 163.367
R964 B.n492 B.n491 163.367
R965 B.n491 B.n490 163.367
R966 B.n490 B.n35 163.367
R967 B.n485 B.n35 163.367
R968 B.n485 B.n484 163.367
R969 B.n484 B.n483 163.367
R970 B.n483 B.n39 163.367
R971 B.n479 B.n39 163.367
R972 B.n479 B.n478 163.367
R973 B.n478 B.n477 163.367
R974 B.n477 B.n41 163.367
R975 B.n473 B.n41 163.367
R976 B.n473 B.n472 163.367
R977 B.n472 B.n45 163.367
R978 B.n468 B.n45 163.367
R979 B.n468 B.n467 163.367
R980 B.n467 B.n466 163.367
R981 B.n466 B.n47 163.367
R982 B.n462 B.n47 163.367
R983 B.n462 B.n461 163.367
R984 B.n461 B.n460 163.367
R985 B.n460 B.n49 163.367
R986 B.n456 B.n49 163.367
R987 B.n456 B.n455 163.367
R988 B.n455 B.n454 163.367
R989 B.n454 B.n51 163.367
R990 B.n450 B.n51 163.367
R991 B.n450 B.n449 163.367
R992 B.n449 B.n448 163.367
R993 B.n448 B.n53 163.367
R994 B.n444 B.n53 163.367
R995 B.n444 B.n443 163.367
R996 B.n443 B.n442 163.367
R997 B.n442 B.n55 163.367
R998 B.n522 B.n521 163.367
R999 B.n522 B.n23 163.367
R1000 B.n526 B.n23 163.367
R1001 B.n527 B.n526 163.367
R1002 B.n528 B.n527 163.367
R1003 B.n528 B.n21 163.367
R1004 B.n532 B.n21 163.367
R1005 B.n533 B.n532 163.367
R1006 B.n534 B.n533 163.367
R1007 B.n534 B.n19 163.367
R1008 B.n538 B.n19 163.367
R1009 B.n539 B.n538 163.367
R1010 B.n540 B.n539 163.367
R1011 B.n540 B.n17 163.367
R1012 B.n544 B.n17 163.367
R1013 B.n545 B.n544 163.367
R1014 B.n546 B.n545 163.367
R1015 B.n546 B.n15 163.367
R1016 B.n550 B.n15 163.367
R1017 B.n551 B.n550 163.367
R1018 B.n552 B.n551 163.367
R1019 B.n552 B.n13 163.367
R1020 B.n556 B.n13 163.367
R1021 B.n557 B.n556 163.367
R1022 B.n558 B.n557 163.367
R1023 B.n558 B.n11 163.367
R1024 B.n562 B.n11 163.367
R1025 B.n563 B.n562 163.367
R1026 B.n564 B.n563 163.367
R1027 B.n564 B.n9 163.367
R1028 B.n568 B.n9 163.367
R1029 B.n569 B.n568 163.367
R1030 B.n570 B.n569 163.367
R1031 B.n570 B.n7 163.367
R1032 B.n574 B.n7 163.367
R1033 B.n575 B.n574 163.367
R1034 B.n576 B.n575 163.367
R1035 B.n576 B.n5 163.367
R1036 B.n580 B.n5 163.367
R1037 B.n581 B.n580 163.367
R1038 B.n582 B.n581 163.367
R1039 B.n582 B.n3 163.367
R1040 B.n586 B.n3 163.367
R1041 B.n587 B.n586 163.367
R1042 B.n152 B.n2 163.367
R1043 B.n152 B.n151 163.367
R1044 B.n156 B.n151 163.367
R1045 B.n157 B.n156 163.367
R1046 B.n158 B.n157 163.367
R1047 B.n158 B.n149 163.367
R1048 B.n162 B.n149 163.367
R1049 B.n163 B.n162 163.367
R1050 B.n164 B.n163 163.367
R1051 B.n164 B.n147 163.367
R1052 B.n168 B.n147 163.367
R1053 B.n169 B.n168 163.367
R1054 B.n170 B.n169 163.367
R1055 B.n170 B.n145 163.367
R1056 B.n174 B.n145 163.367
R1057 B.n175 B.n174 163.367
R1058 B.n176 B.n175 163.367
R1059 B.n176 B.n143 163.367
R1060 B.n180 B.n143 163.367
R1061 B.n181 B.n180 163.367
R1062 B.n182 B.n181 163.367
R1063 B.n182 B.n141 163.367
R1064 B.n186 B.n141 163.367
R1065 B.n187 B.n186 163.367
R1066 B.n188 B.n187 163.367
R1067 B.n188 B.n139 163.367
R1068 B.n192 B.n139 163.367
R1069 B.n193 B.n192 163.367
R1070 B.n194 B.n193 163.367
R1071 B.n194 B.n137 163.367
R1072 B.n198 B.n137 163.367
R1073 B.n199 B.n198 163.367
R1074 B.n200 B.n199 163.367
R1075 B.n200 B.n135 163.367
R1076 B.n204 B.n135 163.367
R1077 B.n205 B.n204 163.367
R1078 B.n206 B.n205 163.367
R1079 B.n206 B.n133 163.367
R1080 B.n210 B.n133 163.367
R1081 B.n211 B.n210 163.367
R1082 B.n212 B.n211 163.367
R1083 B.n212 B.n131 163.367
R1084 B.n216 B.n131 163.367
R1085 B.n217 B.n216 163.367
R1086 B.n119 B.n118 61.6732
R1087 B.n265 B.n264 61.6732
R1088 B.n43 B.n42 61.6732
R1089 B.n37 B.n36 61.6732
R1090 B.n251 B.n119 59.5399
R1091 B.n266 B.n265 59.5399
R1092 B.n44 B.n43 59.5399
R1093 B.n487 B.n37 59.5399
R1094 B.n519 B.n24 32.3127
R1095 B.n440 B.n439 32.3127
R1096 B.n302 B.n301 32.3127
R1097 B.n219 B.n130 32.3127
R1098 B B.n589 18.0485
R1099 B.n523 B.n24 10.6151
R1100 B.n524 B.n523 10.6151
R1101 B.n525 B.n524 10.6151
R1102 B.n525 B.n22 10.6151
R1103 B.n529 B.n22 10.6151
R1104 B.n530 B.n529 10.6151
R1105 B.n531 B.n530 10.6151
R1106 B.n531 B.n20 10.6151
R1107 B.n535 B.n20 10.6151
R1108 B.n536 B.n535 10.6151
R1109 B.n537 B.n536 10.6151
R1110 B.n537 B.n18 10.6151
R1111 B.n541 B.n18 10.6151
R1112 B.n542 B.n541 10.6151
R1113 B.n543 B.n542 10.6151
R1114 B.n543 B.n16 10.6151
R1115 B.n547 B.n16 10.6151
R1116 B.n548 B.n547 10.6151
R1117 B.n549 B.n548 10.6151
R1118 B.n549 B.n14 10.6151
R1119 B.n553 B.n14 10.6151
R1120 B.n554 B.n553 10.6151
R1121 B.n555 B.n554 10.6151
R1122 B.n555 B.n12 10.6151
R1123 B.n559 B.n12 10.6151
R1124 B.n560 B.n559 10.6151
R1125 B.n561 B.n560 10.6151
R1126 B.n561 B.n10 10.6151
R1127 B.n565 B.n10 10.6151
R1128 B.n566 B.n565 10.6151
R1129 B.n567 B.n566 10.6151
R1130 B.n567 B.n8 10.6151
R1131 B.n571 B.n8 10.6151
R1132 B.n572 B.n571 10.6151
R1133 B.n573 B.n572 10.6151
R1134 B.n573 B.n6 10.6151
R1135 B.n577 B.n6 10.6151
R1136 B.n578 B.n577 10.6151
R1137 B.n579 B.n578 10.6151
R1138 B.n579 B.n4 10.6151
R1139 B.n583 B.n4 10.6151
R1140 B.n584 B.n583 10.6151
R1141 B.n585 B.n584 10.6151
R1142 B.n585 B.n0 10.6151
R1143 B.n519 B.n518 10.6151
R1144 B.n518 B.n517 10.6151
R1145 B.n517 B.n26 10.6151
R1146 B.n513 B.n26 10.6151
R1147 B.n513 B.n512 10.6151
R1148 B.n512 B.n511 10.6151
R1149 B.n511 B.n28 10.6151
R1150 B.n507 B.n28 10.6151
R1151 B.n507 B.n506 10.6151
R1152 B.n506 B.n505 10.6151
R1153 B.n505 B.n30 10.6151
R1154 B.n501 B.n30 10.6151
R1155 B.n501 B.n500 10.6151
R1156 B.n500 B.n499 10.6151
R1157 B.n499 B.n32 10.6151
R1158 B.n495 B.n32 10.6151
R1159 B.n495 B.n494 10.6151
R1160 B.n494 B.n493 10.6151
R1161 B.n493 B.n34 10.6151
R1162 B.n489 B.n34 10.6151
R1163 B.n489 B.n488 10.6151
R1164 B.n486 B.n38 10.6151
R1165 B.n482 B.n38 10.6151
R1166 B.n482 B.n481 10.6151
R1167 B.n481 B.n480 10.6151
R1168 B.n480 B.n40 10.6151
R1169 B.n476 B.n40 10.6151
R1170 B.n476 B.n475 10.6151
R1171 B.n475 B.n474 10.6151
R1172 B.n471 B.n470 10.6151
R1173 B.n470 B.n469 10.6151
R1174 B.n469 B.n46 10.6151
R1175 B.n465 B.n46 10.6151
R1176 B.n465 B.n464 10.6151
R1177 B.n464 B.n463 10.6151
R1178 B.n463 B.n48 10.6151
R1179 B.n459 B.n48 10.6151
R1180 B.n459 B.n458 10.6151
R1181 B.n458 B.n457 10.6151
R1182 B.n457 B.n50 10.6151
R1183 B.n453 B.n50 10.6151
R1184 B.n453 B.n452 10.6151
R1185 B.n452 B.n451 10.6151
R1186 B.n451 B.n52 10.6151
R1187 B.n447 B.n52 10.6151
R1188 B.n447 B.n446 10.6151
R1189 B.n446 B.n445 10.6151
R1190 B.n445 B.n54 10.6151
R1191 B.n441 B.n54 10.6151
R1192 B.n441 B.n440 10.6151
R1193 B.n439 B.n56 10.6151
R1194 B.n435 B.n56 10.6151
R1195 B.n435 B.n434 10.6151
R1196 B.n434 B.n433 10.6151
R1197 B.n433 B.n58 10.6151
R1198 B.n429 B.n58 10.6151
R1199 B.n429 B.n428 10.6151
R1200 B.n428 B.n427 10.6151
R1201 B.n427 B.n60 10.6151
R1202 B.n423 B.n60 10.6151
R1203 B.n423 B.n422 10.6151
R1204 B.n422 B.n421 10.6151
R1205 B.n421 B.n62 10.6151
R1206 B.n417 B.n62 10.6151
R1207 B.n417 B.n416 10.6151
R1208 B.n416 B.n415 10.6151
R1209 B.n415 B.n64 10.6151
R1210 B.n411 B.n64 10.6151
R1211 B.n411 B.n410 10.6151
R1212 B.n410 B.n409 10.6151
R1213 B.n409 B.n66 10.6151
R1214 B.n405 B.n66 10.6151
R1215 B.n405 B.n404 10.6151
R1216 B.n404 B.n403 10.6151
R1217 B.n403 B.n68 10.6151
R1218 B.n399 B.n68 10.6151
R1219 B.n399 B.n398 10.6151
R1220 B.n398 B.n397 10.6151
R1221 B.n397 B.n70 10.6151
R1222 B.n393 B.n70 10.6151
R1223 B.n393 B.n392 10.6151
R1224 B.n392 B.n391 10.6151
R1225 B.n391 B.n72 10.6151
R1226 B.n387 B.n72 10.6151
R1227 B.n387 B.n386 10.6151
R1228 B.n386 B.n385 10.6151
R1229 B.n385 B.n74 10.6151
R1230 B.n381 B.n74 10.6151
R1231 B.n381 B.n380 10.6151
R1232 B.n380 B.n379 10.6151
R1233 B.n379 B.n76 10.6151
R1234 B.n375 B.n76 10.6151
R1235 B.n375 B.n374 10.6151
R1236 B.n374 B.n373 10.6151
R1237 B.n373 B.n78 10.6151
R1238 B.n369 B.n78 10.6151
R1239 B.n369 B.n368 10.6151
R1240 B.n368 B.n367 10.6151
R1241 B.n367 B.n80 10.6151
R1242 B.n363 B.n80 10.6151
R1243 B.n363 B.n362 10.6151
R1244 B.n362 B.n361 10.6151
R1245 B.n361 B.n82 10.6151
R1246 B.n357 B.n82 10.6151
R1247 B.n357 B.n356 10.6151
R1248 B.n356 B.n355 10.6151
R1249 B.n355 B.n84 10.6151
R1250 B.n351 B.n84 10.6151
R1251 B.n351 B.n350 10.6151
R1252 B.n350 B.n349 10.6151
R1253 B.n349 B.n86 10.6151
R1254 B.n345 B.n86 10.6151
R1255 B.n345 B.n344 10.6151
R1256 B.n344 B.n343 10.6151
R1257 B.n343 B.n88 10.6151
R1258 B.n339 B.n88 10.6151
R1259 B.n339 B.n338 10.6151
R1260 B.n338 B.n337 10.6151
R1261 B.n337 B.n90 10.6151
R1262 B.n333 B.n90 10.6151
R1263 B.n333 B.n332 10.6151
R1264 B.n332 B.n331 10.6151
R1265 B.n331 B.n92 10.6151
R1266 B.n327 B.n92 10.6151
R1267 B.n327 B.n326 10.6151
R1268 B.n326 B.n325 10.6151
R1269 B.n325 B.n94 10.6151
R1270 B.n321 B.n94 10.6151
R1271 B.n321 B.n320 10.6151
R1272 B.n320 B.n319 10.6151
R1273 B.n319 B.n96 10.6151
R1274 B.n315 B.n96 10.6151
R1275 B.n315 B.n314 10.6151
R1276 B.n314 B.n313 10.6151
R1277 B.n313 B.n98 10.6151
R1278 B.n309 B.n98 10.6151
R1279 B.n309 B.n308 10.6151
R1280 B.n308 B.n307 10.6151
R1281 B.n307 B.n100 10.6151
R1282 B.n303 B.n100 10.6151
R1283 B.n303 B.n302 10.6151
R1284 B.n153 B.n1 10.6151
R1285 B.n154 B.n153 10.6151
R1286 B.n155 B.n154 10.6151
R1287 B.n155 B.n150 10.6151
R1288 B.n159 B.n150 10.6151
R1289 B.n160 B.n159 10.6151
R1290 B.n161 B.n160 10.6151
R1291 B.n161 B.n148 10.6151
R1292 B.n165 B.n148 10.6151
R1293 B.n166 B.n165 10.6151
R1294 B.n167 B.n166 10.6151
R1295 B.n167 B.n146 10.6151
R1296 B.n171 B.n146 10.6151
R1297 B.n172 B.n171 10.6151
R1298 B.n173 B.n172 10.6151
R1299 B.n173 B.n144 10.6151
R1300 B.n177 B.n144 10.6151
R1301 B.n178 B.n177 10.6151
R1302 B.n179 B.n178 10.6151
R1303 B.n179 B.n142 10.6151
R1304 B.n183 B.n142 10.6151
R1305 B.n184 B.n183 10.6151
R1306 B.n185 B.n184 10.6151
R1307 B.n185 B.n140 10.6151
R1308 B.n189 B.n140 10.6151
R1309 B.n190 B.n189 10.6151
R1310 B.n191 B.n190 10.6151
R1311 B.n191 B.n138 10.6151
R1312 B.n195 B.n138 10.6151
R1313 B.n196 B.n195 10.6151
R1314 B.n197 B.n196 10.6151
R1315 B.n197 B.n136 10.6151
R1316 B.n201 B.n136 10.6151
R1317 B.n202 B.n201 10.6151
R1318 B.n203 B.n202 10.6151
R1319 B.n203 B.n134 10.6151
R1320 B.n207 B.n134 10.6151
R1321 B.n208 B.n207 10.6151
R1322 B.n209 B.n208 10.6151
R1323 B.n209 B.n132 10.6151
R1324 B.n213 B.n132 10.6151
R1325 B.n214 B.n213 10.6151
R1326 B.n215 B.n214 10.6151
R1327 B.n215 B.n130 10.6151
R1328 B.n220 B.n219 10.6151
R1329 B.n221 B.n220 10.6151
R1330 B.n221 B.n128 10.6151
R1331 B.n225 B.n128 10.6151
R1332 B.n226 B.n225 10.6151
R1333 B.n227 B.n226 10.6151
R1334 B.n227 B.n126 10.6151
R1335 B.n231 B.n126 10.6151
R1336 B.n232 B.n231 10.6151
R1337 B.n233 B.n232 10.6151
R1338 B.n233 B.n124 10.6151
R1339 B.n237 B.n124 10.6151
R1340 B.n238 B.n237 10.6151
R1341 B.n239 B.n238 10.6151
R1342 B.n239 B.n122 10.6151
R1343 B.n243 B.n122 10.6151
R1344 B.n244 B.n243 10.6151
R1345 B.n245 B.n244 10.6151
R1346 B.n245 B.n120 10.6151
R1347 B.n249 B.n120 10.6151
R1348 B.n250 B.n249 10.6151
R1349 B.n252 B.n116 10.6151
R1350 B.n256 B.n116 10.6151
R1351 B.n257 B.n256 10.6151
R1352 B.n258 B.n257 10.6151
R1353 B.n258 B.n114 10.6151
R1354 B.n262 B.n114 10.6151
R1355 B.n263 B.n262 10.6151
R1356 B.n267 B.n263 10.6151
R1357 B.n271 B.n112 10.6151
R1358 B.n272 B.n271 10.6151
R1359 B.n273 B.n272 10.6151
R1360 B.n273 B.n110 10.6151
R1361 B.n277 B.n110 10.6151
R1362 B.n278 B.n277 10.6151
R1363 B.n279 B.n278 10.6151
R1364 B.n279 B.n108 10.6151
R1365 B.n283 B.n108 10.6151
R1366 B.n284 B.n283 10.6151
R1367 B.n285 B.n284 10.6151
R1368 B.n285 B.n106 10.6151
R1369 B.n289 B.n106 10.6151
R1370 B.n290 B.n289 10.6151
R1371 B.n291 B.n290 10.6151
R1372 B.n291 B.n104 10.6151
R1373 B.n295 B.n104 10.6151
R1374 B.n296 B.n295 10.6151
R1375 B.n297 B.n296 10.6151
R1376 B.n297 B.n102 10.6151
R1377 B.n301 B.n102 10.6151
R1378 B.n589 B.n0 8.11757
R1379 B.n589 B.n1 8.11757
R1380 B.n487 B.n486 6.5566
R1381 B.n474 B.n44 6.5566
R1382 B.n252 B.n251 6.5566
R1383 B.n267 B.n266 6.5566
R1384 B.n488 B.n487 4.05904
R1385 B.n471 B.n44 4.05904
R1386 B.n251 B.n250 4.05904
R1387 B.n266 B.n112 4.05904
C0 w_n3514_n2012# VDD2 1.97634f
C1 VDD1 VP 3.5205f
C2 VTAIL w_n3514_n2012# 2.05059f
C3 VN B 1.17048f
C4 B VDD2 1.70012f
C5 VN VP 5.91272f
C6 VN VDD1 0.151481f
C7 VDD2 VP 0.483514f
C8 VDD1 VDD2 1.5042f
C9 VTAIL B 2.22987f
C10 B w_n3514_n2012# 8.134601f
C11 VTAIL VP 3.90037f
C12 VTAIL VDD1 5.40802f
C13 w_n3514_n2012# VP 7.05278f
C14 VN VDD2 3.1947f
C15 VDD1 w_n3514_n2012# 1.88357f
C16 VTAIL VN 3.88619f
C17 VN w_n3514_n2012# 6.59786f
C18 B VP 1.9314f
C19 VTAIL VDD2 5.46222f
C20 VDD1 B 1.61988f
C21 VDD2 VSUBS 1.464097f
C22 VDD1 VSUBS 1.609359f
C23 VTAIL VSUBS 0.688722f
C24 VN VSUBS 5.8157f
C25 VP VSUBS 2.680531f
C26 B VSUBS 4.06793f
C27 w_n3514_n2012# VSUBS 88.5106f
C28 B.n0 VSUBS 0.006993f
C29 B.n1 VSUBS 0.006993f
C30 B.n2 VSUBS 0.010342f
C31 B.n3 VSUBS 0.007925f
C32 B.n4 VSUBS 0.007925f
C33 B.n5 VSUBS 0.007925f
C34 B.n6 VSUBS 0.007925f
C35 B.n7 VSUBS 0.007925f
C36 B.n8 VSUBS 0.007925f
C37 B.n9 VSUBS 0.007925f
C38 B.n10 VSUBS 0.007925f
C39 B.n11 VSUBS 0.007925f
C40 B.n12 VSUBS 0.007925f
C41 B.n13 VSUBS 0.007925f
C42 B.n14 VSUBS 0.007925f
C43 B.n15 VSUBS 0.007925f
C44 B.n16 VSUBS 0.007925f
C45 B.n17 VSUBS 0.007925f
C46 B.n18 VSUBS 0.007925f
C47 B.n19 VSUBS 0.007925f
C48 B.n20 VSUBS 0.007925f
C49 B.n21 VSUBS 0.007925f
C50 B.n22 VSUBS 0.007925f
C51 B.n23 VSUBS 0.007925f
C52 B.n24 VSUBS 0.017919f
C53 B.n25 VSUBS 0.007925f
C54 B.n26 VSUBS 0.007925f
C55 B.n27 VSUBS 0.007925f
C56 B.n28 VSUBS 0.007925f
C57 B.n29 VSUBS 0.007925f
C58 B.n30 VSUBS 0.007925f
C59 B.n31 VSUBS 0.007925f
C60 B.n32 VSUBS 0.007925f
C61 B.n33 VSUBS 0.007925f
C62 B.n34 VSUBS 0.007925f
C63 B.n35 VSUBS 0.007925f
C64 B.t4 VSUBS 0.086195f
C65 B.t5 VSUBS 0.115492f
C66 B.t3 VSUBS 0.80487f
C67 B.n36 VSUBS 0.197856f
C68 B.n37 VSUBS 0.16149f
C69 B.n38 VSUBS 0.007925f
C70 B.n39 VSUBS 0.007925f
C71 B.n40 VSUBS 0.007925f
C72 B.n41 VSUBS 0.007925f
C73 B.t1 VSUBS 0.086197f
C74 B.t2 VSUBS 0.115493f
C75 B.t0 VSUBS 0.80487f
C76 B.n42 VSUBS 0.197855f
C77 B.n43 VSUBS 0.161488f
C78 B.n44 VSUBS 0.018362f
C79 B.n45 VSUBS 0.007925f
C80 B.n46 VSUBS 0.007925f
C81 B.n47 VSUBS 0.007925f
C82 B.n48 VSUBS 0.007925f
C83 B.n49 VSUBS 0.007925f
C84 B.n50 VSUBS 0.007925f
C85 B.n51 VSUBS 0.007925f
C86 B.n52 VSUBS 0.007925f
C87 B.n53 VSUBS 0.007925f
C88 B.n54 VSUBS 0.007925f
C89 B.n55 VSUBS 0.018911f
C90 B.n56 VSUBS 0.007925f
C91 B.n57 VSUBS 0.007925f
C92 B.n58 VSUBS 0.007925f
C93 B.n59 VSUBS 0.007925f
C94 B.n60 VSUBS 0.007925f
C95 B.n61 VSUBS 0.007925f
C96 B.n62 VSUBS 0.007925f
C97 B.n63 VSUBS 0.007925f
C98 B.n64 VSUBS 0.007925f
C99 B.n65 VSUBS 0.007925f
C100 B.n66 VSUBS 0.007925f
C101 B.n67 VSUBS 0.007925f
C102 B.n68 VSUBS 0.007925f
C103 B.n69 VSUBS 0.007925f
C104 B.n70 VSUBS 0.007925f
C105 B.n71 VSUBS 0.007925f
C106 B.n72 VSUBS 0.007925f
C107 B.n73 VSUBS 0.007925f
C108 B.n74 VSUBS 0.007925f
C109 B.n75 VSUBS 0.007925f
C110 B.n76 VSUBS 0.007925f
C111 B.n77 VSUBS 0.007925f
C112 B.n78 VSUBS 0.007925f
C113 B.n79 VSUBS 0.007925f
C114 B.n80 VSUBS 0.007925f
C115 B.n81 VSUBS 0.007925f
C116 B.n82 VSUBS 0.007925f
C117 B.n83 VSUBS 0.007925f
C118 B.n84 VSUBS 0.007925f
C119 B.n85 VSUBS 0.007925f
C120 B.n86 VSUBS 0.007925f
C121 B.n87 VSUBS 0.007925f
C122 B.n88 VSUBS 0.007925f
C123 B.n89 VSUBS 0.007925f
C124 B.n90 VSUBS 0.007925f
C125 B.n91 VSUBS 0.007925f
C126 B.n92 VSUBS 0.007925f
C127 B.n93 VSUBS 0.007925f
C128 B.n94 VSUBS 0.007925f
C129 B.n95 VSUBS 0.007925f
C130 B.n96 VSUBS 0.007925f
C131 B.n97 VSUBS 0.007925f
C132 B.n98 VSUBS 0.007925f
C133 B.n99 VSUBS 0.007925f
C134 B.n100 VSUBS 0.007925f
C135 B.n101 VSUBS 0.017919f
C136 B.n102 VSUBS 0.007925f
C137 B.n103 VSUBS 0.007925f
C138 B.n104 VSUBS 0.007925f
C139 B.n105 VSUBS 0.007925f
C140 B.n106 VSUBS 0.007925f
C141 B.n107 VSUBS 0.007925f
C142 B.n108 VSUBS 0.007925f
C143 B.n109 VSUBS 0.007925f
C144 B.n110 VSUBS 0.007925f
C145 B.n111 VSUBS 0.007925f
C146 B.n112 VSUBS 0.005478f
C147 B.n113 VSUBS 0.007925f
C148 B.n114 VSUBS 0.007925f
C149 B.n115 VSUBS 0.007925f
C150 B.n116 VSUBS 0.007925f
C151 B.n117 VSUBS 0.007925f
C152 B.t11 VSUBS 0.086195f
C153 B.t10 VSUBS 0.115492f
C154 B.t9 VSUBS 0.80487f
C155 B.n118 VSUBS 0.197856f
C156 B.n119 VSUBS 0.16149f
C157 B.n120 VSUBS 0.007925f
C158 B.n121 VSUBS 0.007925f
C159 B.n122 VSUBS 0.007925f
C160 B.n123 VSUBS 0.007925f
C161 B.n124 VSUBS 0.007925f
C162 B.n125 VSUBS 0.007925f
C163 B.n126 VSUBS 0.007925f
C164 B.n127 VSUBS 0.007925f
C165 B.n128 VSUBS 0.007925f
C166 B.n129 VSUBS 0.007925f
C167 B.n130 VSUBS 0.017919f
C168 B.n131 VSUBS 0.007925f
C169 B.n132 VSUBS 0.007925f
C170 B.n133 VSUBS 0.007925f
C171 B.n134 VSUBS 0.007925f
C172 B.n135 VSUBS 0.007925f
C173 B.n136 VSUBS 0.007925f
C174 B.n137 VSUBS 0.007925f
C175 B.n138 VSUBS 0.007925f
C176 B.n139 VSUBS 0.007925f
C177 B.n140 VSUBS 0.007925f
C178 B.n141 VSUBS 0.007925f
C179 B.n142 VSUBS 0.007925f
C180 B.n143 VSUBS 0.007925f
C181 B.n144 VSUBS 0.007925f
C182 B.n145 VSUBS 0.007925f
C183 B.n146 VSUBS 0.007925f
C184 B.n147 VSUBS 0.007925f
C185 B.n148 VSUBS 0.007925f
C186 B.n149 VSUBS 0.007925f
C187 B.n150 VSUBS 0.007925f
C188 B.n151 VSUBS 0.007925f
C189 B.n152 VSUBS 0.007925f
C190 B.n153 VSUBS 0.007925f
C191 B.n154 VSUBS 0.007925f
C192 B.n155 VSUBS 0.007925f
C193 B.n156 VSUBS 0.007925f
C194 B.n157 VSUBS 0.007925f
C195 B.n158 VSUBS 0.007925f
C196 B.n159 VSUBS 0.007925f
C197 B.n160 VSUBS 0.007925f
C198 B.n161 VSUBS 0.007925f
C199 B.n162 VSUBS 0.007925f
C200 B.n163 VSUBS 0.007925f
C201 B.n164 VSUBS 0.007925f
C202 B.n165 VSUBS 0.007925f
C203 B.n166 VSUBS 0.007925f
C204 B.n167 VSUBS 0.007925f
C205 B.n168 VSUBS 0.007925f
C206 B.n169 VSUBS 0.007925f
C207 B.n170 VSUBS 0.007925f
C208 B.n171 VSUBS 0.007925f
C209 B.n172 VSUBS 0.007925f
C210 B.n173 VSUBS 0.007925f
C211 B.n174 VSUBS 0.007925f
C212 B.n175 VSUBS 0.007925f
C213 B.n176 VSUBS 0.007925f
C214 B.n177 VSUBS 0.007925f
C215 B.n178 VSUBS 0.007925f
C216 B.n179 VSUBS 0.007925f
C217 B.n180 VSUBS 0.007925f
C218 B.n181 VSUBS 0.007925f
C219 B.n182 VSUBS 0.007925f
C220 B.n183 VSUBS 0.007925f
C221 B.n184 VSUBS 0.007925f
C222 B.n185 VSUBS 0.007925f
C223 B.n186 VSUBS 0.007925f
C224 B.n187 VSUBS 0.007925f
C225 B.n188 VSUBS 0.007925f
C226 B.n189 VSUBS 0.007925f
C227 B.n190 VSUBS 0.007925f
C228 B.n191 VSUBS 0.007925f
C229 B.n192 VSUBS 0.007925f
C230 B.n193 VSUBS 0.007925f
C231 B.n194 VSUBS 0.007925f
C232 B.n195 VSUBS 0.007925f
C233 B.n196 VSUBS 0.007925f
C234 B.n197 VSUBS 0.007925f
C235 B.n198 VSUBS 0.007925f
C236 B.n199 VSUBS 0.007925f
C237 B.n200 VSUBS 0.007925f
C238 B.n201 VSUBS 0.007925f
C239 B.n202 VSUBS 0.007925f
C240 B.n203 VSUBS 0.007925f
C241 B.n204 VSUBS 0.007925f
C242 B.n205 VSUBS 0.007925f
C243 B.n206 VSUBS 0.007925f
C244 B.n207 VSUBS 0.007925f
C245 B.n208 VSUBS 0.007925f
C246 B.n209 VSUBS 0.007925f
C247 B.n210 VSUBS 0.007925f
C248 B.n211 VSUBS 0.007925f
C249 B.n212 VSUBS 0.007925f
C250 B.n213 VSUBS 0.007925f
C251 B.n214 VSUBS 0.007925f
C252 B.n215 VSUBS 0.007925f
C253 B.n216 VSUBS 0.007925f
C254 B.n217 VSUBS 0.017919f
C255 B.n218 VSUBS 0.018911f
C256 B.n219 VSUBS 0.018911f
C257 B.n220 VSUBS 0.007925f
C258 B.n221 VSUBS 0.007925f
C259 B.n222 VSUBS 0.007925f
C260 B.n223 VSUBS 0.007925f
C261 B.n224 VSUBS 0.007925f
C262 B.n225 VSUBS 0.007925f
C263 B.n226 VSUBS 0.007925f
C264 B.n227 VSUBS 0.007925f
C265 B.n228 VSUBS 0.007925f
C266 B.n229 VSUBS 0.007925f
C267 B.n230 VSUBS 0.007925f
C268 B.n231 VSUBS 0.007925f
C269 B.n232 VSUBS 0.007925f
C270 B.n233 VSUBS 0.007925f
C271 B.n234 VSUBS 0.007925f
C272 B.n235 VSUBS 0.007925f
C273 B.n236 VSUBS 0.007925f
C274 B.n237 VSUBS 0.007925f
C275 B.n238 VSUBS 0.007925f
C276 B.n239 VSUBS 0.007925f
C277 B.n240 VSUBS 0.007925f
C278 B.n241 VSUBS 0.007925f
C279 B.n242 VSUBS 0.007925f
C280 B.n243 VSUBS 0.007925f
C281 B.n244 VSUBS 0.007925f
C282 B.n245 VSUBS 0.007925f
C283 B.n246 VSUBS 0.007925f
C284 B.n247 VSUBS 0.007925f
C285 B.n248 VSUBS 0.007925f
C286 B.n249 VSUBS 0.007925f
C287 B.n250 VSUBS 0.005478f
C288 B.n251 VSUBS 0.018362f
C289 B.n252 VSUBS 0.00641f
C290 B.n253 VSUBS 0.007925f
C291 B.n254 VSUBS 0.007925f
C292 B.n255 VSUBS 0.007925f
C293 B.n256 VSUBS 0.007925f
C294 B.n257 VSUBS 0.007925f
C295 B.n258 VSUBS 0.007925f
C296 B.n259 VSUBS 0.007925f
C297 B.n260 VSUBS 0.007925f
C298 B.n261 VSUBS 0.007925f
C299 B.n262 VSUBS 0.007925f
C300 B.n263 VSUBS 0.007925f
C301 B.t8 VSUBS 0.086197f
C302 B.t7 VSUBS 0.115493f
C303 B.t6 VSUBS 0.80487f
C304 B.n264 VSUBS 0.197855f
C305 B.n265 VSUBS 0.161488f
C306 B.n266 VSUBS 0.018362f
C307 B.n267 VSUBS 0.00641f
C308 B.n268 VSUBS 0.007925f
C309 B.n269 VSUBS 0.007925f
C310 B.n270 VSUBS 0.007925f
C311 B.n271 VSUBS 0.007925f
C312 B.n272 VSUBS 0.007925f
C313 B.n273 VSUBS 0.007925f
C314 B.n274 VSUBS 0.007925f
C315 B.n275 VSUBS 0.007925f
C316 B.n276 VSUBS 0.007925f
C317 B.n277 VSUBS 0.007925f
C318 B.n278 VSUBS 0.007925f
C319 B.n279 VSUBS 0.007925f
C320 B.n280 VSUBS 0.007925f
C321 B.n281 VSUBS 0.007925f
C322 B.n282 VSUBS 0.007925f
C323 B.n283 VSUBS 0.007925f
C324 B.n284 VSUBS 0.007925f
C325 B.n285 VSUBS 0.007925f
C326 B.n286 VSUBS 0.007925f
C327 B.n287 VSUBS 0.007925f
C328 B.n288 VSUBS 0.007925f
C329 B.n289 VSUBS 0.007925f
C330 B.n290 VSUBS 0.007925f
C331 B.n291 VSUBS 0.007925f
C332 B.n292 VSUBS 0.007925f
C333 B.n293 VSUBS 0.007925f
C334 B.n294 VSUBS 0.007925f
C335 B.n295 VSUBS 0.007925f
C336 B.n296 VSUBS 0.007925f
C337 B.n297 VSUBS 0.007925f
C338 B.n298 VSUBS 0.007925f
C339 B.n299 VSUBS 0.007925f
C340 B.n300 VSUBS 0.018911f
C341 B.n301 VSUBS 0.017965f
C342 B.n302 VSUBS 0.018865f
C343 B.n303 VSUBS 0.007925f
C344 B.n304 VSUBS 0.007925f
C345 B.n305 VSUBS 0.007925f
C346 B.n306 VSUBS 0.007925f
C347 B.n307 VSUBS 0.007925f
C348 B.n308 VSUBS 0.007925f
C349 B.n309 VSUBS 0.007925f
C350 B.n310 VSUBS 0.007925f
C351 B.n311 VSUBS 0.007925f
C352 B.n312 VSUBS 0.007925f
C353 B.n313 VSUBS 0.007925f
C354 B.n314 VSUBS 0.007925f
C355 B.n315 VSUBS 0.007925f
C356 B.n316 VSUBS 0.007925f
C357 B.n317 VSUBS 0.007925f
C358 B.n318 VSUBS 0.007925f
C359 B.n319 VSUBS 0.007925f
C360 B.n320 VSUBS 0.007925f
C361 B.n321 VSUBS 0.007925f
C362 B.n322 VSUBS 0.007925f
C363 B.n323 VSUBS 0.007925f
C364 B.n324 VSUBS 0.007925f
C365 B.n325 VSUBS 0.007925f
C366 B.n326 VSUBS 0.007925f
C367 B.n327 VSUBS 0.007925f
C368 B.n328 VSUBS 0.007925f
C369 B.n329 VSUBS 0.007925f
C370 B.n330 VSUBS 0.007925f
C371 B.n331 VSUBS 0.007925f
C372 B.n332 VSUBS 0.007925f
C373 B.n333 VSUBS 0.007925f
C374 B.n334 VSUBS 0.007925f
C375 B.n335 VSUBS 0.007925f
C376 B.n336 VSUBS 0.007925f
C377 B.n337 VSUBS 0.007925f
C378 B.n338 VSUBS 0.007925f
C379 B.n339 VSUBS 0.007925f
C380 B.n340 VSUBS 0.007925f
C381 B.n341 VSUBS 0.007925f
C382 B.n342 VSUBS 0.007925f
C383 B.n343 VSUBS 0.007925f
C384 B.n344 VSUBS 0.007925f
C385 B.n345 VSUBS 0.007925f
C386 B.n346 VSUBS 0.007925f
C387 B.n347 VSUBS 0.007925f
C388 B.n348 VSUBS 0.007925f
C389 B.n349 VSUBS 0.007925f
C390 B.n350 VSUBS 0.007925f
C391 B.n351 VSUBS 0.007925f
C392 B.n352 VSUBS 0.007925f
C393 B.n353 VSUBS 0.007925f
C394 B.n354 VSUBS 0.007925f
C395 B.n355 VSUBS 0.007925f
C396 B.n356 VSUBS 0.007925f
C397 B.n357 VSUBS 0.007925f
C398 B.n358 VSUBS 0.007925f
C399 B.n359 VSUBS 0.007925f
C400 B.n360 VSUBS 0.007925f
C401 B.n361 VSUBS 0.007925f
C402 B.n362 VSUBS 0.007925f
C403 B.n363 VSUBS 0.007925f
C404 B.n364 VSUBS 0.007925f
C405 B.n365 VSUBS 0.007925f
C406 B.n366 VSUBS 0.007925f
C407 B.n367 VSUBS 0.007925f
C408 B.n368 VSUBS 0.007925f
C409 B.n369 VSUBS 0.007925f
C410 B.n370 VSUBS 0.007925f
C411 B.n371 VSUBS 0.007925f
C412 B.n372 VSUBS 0.007925f
C413 B.n373 VSUBS 0.007925f
C414 B.n374 VSUBS 0.007925f
C415 B.n375 VSUBS 0.007925f
C416 B.n376 VSUBS 0.007925f
C417 B.n377 VSUBS 0.007925f
C418 B.n378 VSUBS 0.007925f
C419 B.n379 VSUBS 0.007925f
C420 B.n380 VSUBS 0.007925f
C421 B.n381 VSUBS 0.007925f
C422 B.n382 VSUBS 0.007925f
C423 B.n383 VSUBS 0.007925f
C424 B.n384 VSUBS 0.007925f
C425 B.n385 VSUBS 0.007925f
C426 B.n386 VSUBS 0.007925f
C427 B.n387 VSUBS 0.007925f
C428 B.n388 VSUBS 0.007925f
C429 B.n389 VSUBS 0.007925f
C430 B.n390 VSUBS 0.007925f
C431 B.n391 VSUBS 0.007925f
C432 B.n392 VSUBS 0.007925f
C433 B.n393 VSUBS 0.007925f
C434 B.n394 VSUBS 0.007925f
C435 B.n395 VSUBS 0.007925f
C436 B.n396 VSUBS 0.007925f
C437 B.n397 VSUBS 0.007925f
C438 B.n398 VSUBS 0.007925f
C439 B.n399 VSUBS 0.007925f
C440 B.n400 VSUBS 0.007925f
C441 B.n401 VSUBS 0.007925f
C442 B.n402 VSUBS 0.007925f
C443 B.n403 VSUBS 0.007925f
C444 B.n404 VSUBS 0.007925f
C445 B.n405 VSUBS 0.007925f
C446 B.n406 VSUBS 0.007925f
C447 B.n407 VSUBS 0.007925f
C448 B.n408 VSUBS 0.007925f
C449 B.n409 VSUBS 0.007925f
C450 B.n410 VSUBS 0.007925f
C451 B.n411 VSUBS 0.007925f
C452 B.n412 VSUBS 0.007925f
C453 B.n413 VSUBS 0.007925f
C454 B.n414 VSUBS 0.007925f
C455 B.n415 VSUBS 0.007925f
C456 B.n416 VSUBS 0.007925f
C457 B.n417 VSUBS 0.007925f
C458 B.n418 VSUBS 0.007925f
C459 B.n419 VSUBS 0.007925f
C460 B.n420 VSUBS 0.007925f
C461 B.n421 VSUBS 0.007925f
C462 B.n422 VSUBS 0.007925f
C463 B.n423 VSUBS 0.007925f
C464 B.n424 VSUBS 0.007925f
C465 B.n425 VSUBS 0.007925f
C466 B.n426 VSUBS 0.007925f
C467 B.n427 VSUBS 0.007925f
C468 B.n428 VSUBS 0.007925f
C469 B.n429 VSUBS 0.007925f
C470 B.n430 VSUBS 0.007925f
C471 B.n431 VSUBS 0.007925f
C472 B.n432 VSUBS 0.007925f
C473 B.n433 VSUBS 0.007925f
C474 B.n434 VSUBS 0.007925f
C475 B.n435 VSUBS 0.007925f
C476 B.n436 VSUBS 0.007925f
C477 B.n437 VSUBS 0.007925f
C478 B.n438 VSUBS 0.017919f
C479 B.n439 VSUBS 0.017919f
C480 B.n440 VSUBS 0.018911f
C481 B.n441 VSUBS 0.007925f
C482 B.n442 VSUBS 0.007925f
C483 B.n443 VSUBS 0.007925f
C484 B.n444 VSUBS 0.007925f
C485 B.n445 VSUBS 0.007925f
C486 B.n446 VSUBS 0.007925f
C487 B.n447 VSUBS 0.007925f
C488 B.n448 VSUBS 0.007925f
C489 B.n449 VSUBS 0.007925f
C490 B.n450 VSUBS 0.007925f
C491 B.n451 VSUBS 0.007925f
C492 B.n452 VSUBS 0.007925f
C493 B.n453 VSUBS 0.007925f
C494 B.n454 VSUBS 0.007925f
C495 B.n455 VSUBS 0.007925f
C496 B.n456 VSUBS 0.007925f
C497 B.n457 VSUBS 0.007925f
C498 B.n458 VSUBS 0.007925f
C499 B.n459 VSUBS 0.007925f
C500 B.n460 VSUBS 0.007925f
C501 B.n461 VSUBS 0.007925f
C502 B.n462 VSUBS 0.007925f
C503 B.n463 VSUBS 0.007925f
C504 B.n464 VSUBS 0.007925f
C505 B.n465 VSUBS 0.007925f
C506 B.n466 VSUBS 0.007925f
C507 B.n467 VSUBS 0.007925f
C508 B.n468 VSUBS 0.007925f
C509 B.n469 VSUBS 0.007925f
C510 B.n470 VSUBS 0.007925f
C511 B.n471 VSUBS 0.005478f
C512 B.n472 VSUBS 0.007925f
C513 B.n473 VSUBS 0.007925f
C514 B.n474 VSUBS 0.00641f
C515 B.n475 VSUBS 0.007925f
C516 B.n476 VSUBS 0.007925f
C517 B.n477 VSUBS 0.007925f
C518 B.n478 VSUBS 0.007925f
C519 B.n479 VSUBS 0.007925f
C520 B.n480 VSUBS 0.007925f
C521 B.n481 VSUBS 0.007925f
C522 B.n482 VSUBS 0.007925f
C523 B.n483 VSUBS 0.007925f
C524 B.n484 VSUBS 0.007925f
C525 B.n485 VSUBS 0.007925f
C526 B.n486 VSUBS 0.00641f
C527 B.n487 VSUBS 0.018362f
C528 B.n488 VSUBS 0.005478f
C529 B.n489 VSUBS 0.007925f
C530 B.n490 VSUBS 0.007925f
C531 B.n491 VSUBS 0.007925f
C532 B.n492 VSUBS 0.007925f
C533 B.n493 VSUBS 0.007925f
C534 B.n494 VSUBS 0.007925f
C535 B.n495 VSUBS 0.007925f
C536 B.n496 VSUBS 0.007925f
C537 B.n497 VSUBS 0.007925f
C538 B.n498 VSUBS 0.007925f
C539 B.n499 VSUBS 0.007925f
C540 B.n500 VSUBS 0.007925f
C541 B.n501 VSUBS 0.007925f
C542 B.n502 VSUBS 0.007925f
C543 B.n503 VSUBS 0.007925f
C544 B.n504 VSUBS 0.007925f
C545 B.n505 VSUBS 0.007925f
C546 B.n506 VSUBS 0.007925f
C547 B.n507 VSUBS 0.007925f
C548 B.n508 VSUBS 0.007925f
C549 B.n509 VSUBS 0.007925f
C550 B.n510 VSUBS 0.007925f
C551 B.n511 VSUBS 0.007925f
C552 B.n512 VSUBS 0.007925f
C553 B.n513 VSUBS 0.007925f
C554 B.n514 VSUBS 0.007925f
C555 B.n515 VSUBS 0.007925f
C556 B.n516 VSUBS 0.007925f
C557 B.n517 VSUBS 0.007925f
C558 B.n518 VSUBS 0.007925f
C559 B.n519 VSUBS 0.018911f
C560 B.n520 VSUBS 0.018911f
C561 B.n521 VSUBS 0.017919f
C562 B.n522 VSUBS 0.007925f
C563 B.n523 VSUBS 0.007925f
C564 B.n524 VSUBS 0.007925f
C565 B.n525 VSUBS 0.007925f
C566 B.n526 VSUBS 0.007925f
C567 B.n527 VSUBS 0.007925f
C568 B.n528 VSUBS 0.007925f
C569 B.n529 VSUBS 0.007925f
C570 B.n530 VSUBS 0.007925f
C571 B.n531 VSUBS 0.007925f
C572 B.n532 VSUBS 0.007925f
C573 B.n533 VSUBS 0.007925f
C574 B.n534 VSUBS 0.007925f
C575 B.n535 VSUBS 0.007925f
C576 B.n536 VSUBS 0.007925f
C577 B.n537 VSUBS 0.007925f
C578 B.n538 VSUBS 0.007925f
C579 B.n539 VSUBS 0.007925f
C580 B.n540 VSUBS 0.007925f
C581 B.n541 VSUBS 0.007925f
C582 B.n542 VSUBS 0.007925f
C583 B.n543 VSUBS 0.007925f
C584 B.n544 VSUBS 0.007925f
C585 B.n545 VSUBS 0.007925f
C586 B.n546 VSUBS 0.007925f
C587 B.n547 VSUBS 0.007925f
C588 B.n548 VSUBS 0.007925f
C589 B.n549 VSUBS 0.007925f
C590 B.n550 VSUBS 0.007925f
C591 B.n551 VSUBS 0.007925f
C592 B.n552 VSUBS 0.007925f
C593 B.n553 VSUBS 0.007925f
C594 B.n554 VSUBS 0.007925f
C595 B.n555 VSUBS 0.007925f
C596 B.n556 VSUBS 0.007925f
C597 B.n557 VSUBS 0.007925f
C598 B.n558 VSUBS 0.007925f
C599 B.n559 VSUBS 0.007925f
C600 B.n560 VSUBS 0.007925f
C601 B.n561 VSUBS 0.007925f
C602 B.n562 VSUBS 0.007925f
C603 B.n563 VSUBS 0.007925f
C604 B.n564 VSUBS 0.007925f
C605 B.n565 VSUBS 0.007925f
C606 B.n566 VSUBS 0.007925f
C607 B.n567 VSUBS 0.007925f
C608 B.n568 VSUBS 0.007925f
C609 B.n569 VSUBS 0.007925f
C610 B.n570 VSUBS 0.007925f
C611 B.n571 VSUBS 0.007925f
C612 B.n572 VSUBS 0.007925f
C613 B.n573 VSUBS 0.007925f
C614 B.n574 VSUBS 0.007925f
C615 B.n575 VSUBS 0.007925f
C616 B.n576 VSUBS 0.007925f
C617 B.n577 VSUBS 0.007925f
C618 B.n578 VSUBS 0.007925f
C619 B.n579 VSUBS 0.007925f
C620 B.n580 VSUBS 0.007925f
C621 B.n581 VSUBS 0.007925f
C622 B.n582 VSUBS 0.007925f
C623 B.n583 VSUBS 0.007925f
C624 B.n584 VSUBS 0.007925f
C625 B.n585 VSUBS 0.007925f
C626 B.n586 VSUBS 0.007925f
C627 B.n587 VSUBS 0.010342f
C628 B.n588 VSUBS 0.011017f
C629 B.n589 VSUBS 0.021909f
C630 VDD2.n0 VSUBS 0.023206f
C631 VDD2.n1 VSUBS 0.022055f
C632 VDD2.n2 VSUBS 0.011851f
C633 VDD2.n3 VSUBS 0.028012f
C634 VDD2.n4 VSUBS 0.012548f
C635 VDD2.n5 VSUBS 0.022055f
C636 VDD2.n6 VSUBS 0.011851f
C637 VDD2.n7 VSUBS 0.021009f
C638 VDD2.n8 VSUBS 0.017793f
C639 VDD2.t2 VSUBS 0.060278f
C640 VDD2.n9 VSUBS 0.092593f
C641 VDD2.n10 VSUBS 0.427474f
C642 VDD2.n11 VSUBS 0.011851f
C643 VDD2.n12 VSUBS 0.012548f
C644 VDD2.n13 VSUBS 0.028012f
C645 VDD2.n14 VSUBS 0.028012f
C646 VDD2.n15 VSUBS 0.012548f
C647 VDD2.n16 VSUBS 0.011851f
C648 VDD2.n17 VSUBS 0.022055f
C649 VDD2.n18 VSUBS 0.022055f
C650 VDD2.n19 VSUBS 0.011851f
C651 VDD2.n20 VSUBS 0.012548f
C652 VDD2.n21 VSUBS 0.028012f
C653 VDD2.n22 VSUBS 0.064315f
C654 VDD2.n23 VSUBS 0.012548f
C655 VDD2.n24 VSUBS 0.011851f
C656 VDD2.n25 VSUBS 0.049171f
C657 VDD2.n26 VSUBS 0.054777f
C658 VDD2.t3 VSUBS 0.090976f
C659 VDD2.t5 VSUBS 0.090976f
C660 VDD2.n27 VSUBS 0.581736f
C661 VDD2.n28 VSUBS 2.25726f
C662 VDD2.n29 VSUBS 0.023206f
C663 VDD2.n30 VSUBS 0.022055f
C664 VDD2.n31 VSUBS 0.011851f
C665 VDD2.n32 VSUBS 0.028012f
C666 VDD2.n33 VSUBS 0.012548f
C667 VDD2.n34 VSUBS 0.022055f
C668 VDD2.n35 VSUBS 0.011851f
C669 VDD2.n36 VSUBS 0.021009f
C670 VDD2.n37 VSUBS 0.017793f
C671 VDD2.t1 VSUBS 0.060278f
C672 VDD2.n38 VSUBS 0.092593f
C673 VDD2.n39 VSUBS 0.427474f
C674 VDD2.n40 VSUBS 0.011851f
C675 VDD2.n41 VSUBS 0.012548f
C676 VDD2.n42 VSUBS 0.028012f
C677 VDD2.n43 VSUBS 0.028012f
C678 VDD2.n44 VSUBS 0.012548f
C679 VDD2.n45 VSUBS 0.011851f
C680 VDD2.n46 VSUBS 0.022055f
C681 VDD2.n47 VSUBS 0.022055f
C682 VDD2.n48 VSUBS 0.011851f
C683 VDD2.n49 VSUBS 0.012548f
C684 VDD2.n50 VSUBS 0.028012f
C685 VDD2.n51 VSUBS 0.064315f
C686 VDD2.n52 VSUBS 0.012548f
C687 VDD2.n53 VSUBS 0.011851f
C688 VDD2.n54 VSUBS 0.049171f
C689 VDD2.n55 VSUBS 0.047375f
C690 VDD2.n56 VSUBS 1.85019f
C691 VDD2.t0 VSUBS 0.090976f
C692 VDD2.t4 VSUBS 0.090976f
C693 VDD2.n57 VSUBS 0.581712f
C694 VN.t0 VSUBS 1.50334f
C695 VN.n0 VSUBS 0.717767f
C696 VN.n1 VSUBS 0.038518f
C697 VN.n2 VSUBS 0.065488f
C698 VN.n3 VSUBS 0.409075f
C699 VN.t2 VSUBS 1.50334f
C700 VN.t3 VSUBS 1.84682f
C701 VN.n4 VSUBS 0.663672f
C702 VN.n5 VSUBS 0.688939f
C703 VN.n6 VSUBS 0.053796f
C704 VN.n7 VSUBS 0.071427f
C705 VN.n8 VSUBS 0.038518f
C706 VN.n9 VSUBS 0.038518f
C707 VN.n10 VSUBS 0.038518f
C708 VN.n11 VSUBS 0.045827f
C709 VN.n12 VSUBS 0.072095f
C710 VN.n13 VSUBS 0.066491f
C711 VN.n14 VSUBS 0.062157f
C712 VN.n15 VSUBS 0.076454f
C713 VN.t4 VSUBS 1.50334f
C714 VN.n16 VSUBS 0.717767f
C715 VN.n17 VSUBS 0.038518f
C716 VN.n18 VSUBS 0.065488f
C717 VN.n19 VSUBS 0.409075f
C718 VN.t5 VSUBS 1.50334f
C719 VN.t1 VSUBS 1.84682f
C720 VN.n20 VSUBS 0.663672f
C721 VN.n21 VSUBS 0.688939f
C722 VN.n22 VSUBS 0.053796f
C723 VN.n23 VSUBS 0.071427f
C724 VN.n24 VSUBS 0.038518f
C725 VN.n25 VSUBS 0.038518f
C726 VN.n26 VSUBS 0.038518f
C727 VN.n27 VSUBS 0.045827f
C728 VN.n28 VSUBS 0.072095f
C729 VN.n29 VSUBS 0.066491f
C730 VN.n30 VSUBS 0.062157f
C731 VN.n31 VSUBS 1.84948f
C732 VTAIL.t4 VSUBS 0.143488f
C733 VTAIL.t1 VSUBS 0.143488f
C734 VTAIL.n0 VSUBS 0.799013f
C735 VTAIL.n1 VSUBS 0.897158f
C736 VTAIL.n2 VSUBS 0.036601f
C737 VTAIL.n3 VSUBS 0.034785f
C738 VTAIL.n4 VSUBS 0.018692f
C739 VTAIL.n5 VSUBS 0.044181f
C740 VTAIL.n6 VSUBS 0.019791f
C741 VTAIL.n7 VSUBS 0.034785f
C742 VTAIL.n8 VSUBS 0.018692f
C743 VTAIL.n9 VSUBS 0.033136f
C744 VTAIL.n10 VSUBS 0.028064f
C745 VTAIL.t10 VSUBS 0.095071f
C746 VTAIL.n11 VSUBS 0.146038f
C747 VTAIL.n12 VSUBS 0.674217f
C748 VTAIL.n13 VSUBS 0.018692f
C749 VTAIL.n14 VSUBS 0.019791f
C750 VTAIL.n15 VSUBS 0.044181f
C751 VTAIL.n16 VSUBS 0.044181f
C752 VTAIL.n17 VSUBS 0.019791f
C753 VTAIL.n18 VSUBS 0.018692f
C754 VTAIL.n19 VSUBS 0.034785f
C755 VTAIL.n20 VSUBS 0.034785f
C756 VTAIL.n21 VSUBS 0.018692f
C757 VTAIL.n22 VSUBS 0.019791f
C758 VTAIL.n23 VSUBS 0.044181f
C759 VTAIL.n24 VSUBS 0.101439f
C760 VTAIL.n25 VSUBS 0.019791f
C761 VTAIL.n26 VSUBS 0.018692f
C762 VTAIL.n27 VSUBS 0.077552f
C763 VTAIL.n28 VSUBS 0.050679f
C764 VTAIL.n29 VSUBS 0.541661f
C765 VTAIL.t6 VSUBS 0.143488f
C766 VTAIL.t11 VSUBS 0.143488f
C767 VTAIL.n30 VSUBS 0.799013f
C768 VTAIL.n31 VSUBS 2.50622f
C769 VTAIL.t3 VSUBS 0.143488f
C770 VTAIL.t2 VSUBS 0.143488f
C771 VTAIL.n32 VSUBS 0.799019f
C772 VTAIL.n33 VSUBS 2.50621f
C773 VTAIL.n34 VSUBS 0.036601f
C774 VTAIL.n35 VSUBS 0.034785f
C775 VTAIL.n36 VSUBS 0.018692f
C776 VTAIL.n37 VSUBS 0.044181f
C777 VTAIL.n38 VSUBS 0.019791f
C778 VTAIL.n39 VSUBS 0.034785f
C779 VTAIL.n40 VSUBS 0.018692f
C780 VTAIL.n41 VSUBS 0.033136f
C781 VTAIL.n42 VSUBS 0.028064f
C782 VTAIL.t5 VSUBS 0.095071f
C783 VTAIL.n43 VSUBS 0.146038f
C784 VTAIL.n44 VSUBS 0.674217f
C785 VTAIL.n45 VSUBS 0.018692f
C786 VTAIL.n46 VSUBS 0.019791f
C787 VTAIL.n47 VSUBS 0.044181f
C788 VTAIL.n48 VSUBS 0.044181f
C789 VTAIL.n49 VSUBS 0.019791f
C790 VTAIL.n50 VSUBS 0.018692f
C791 VTAIL.n51 VSUBS 0.034785f
C792 VTAIL.n52 VSUBS 0.034785f
C793 VTAIL.n53 VSUBS 0.018692f
C794 VTAIL.n54 VSUBS 0.019791f
C795 VTAIL.n55 VSUBS 0.044181f
C796 VTAIL.n56 VSUBS 0.101439f
C797 VTAIL.n57 VSUBS 0.019791f
C798 VTAIL.n58 VSUBS 0.018692f
C799 VTAIL.n59 VSUBS 0.077552f
C800 VTAIL.n60 VSUBS 0.050679f
C801 VTAIL.n61 VSUBS 0.541661f
C802 VTAIL.t8 VSUBS 0.143488f
C803 VTAIL.t7 VSUBS 0.143488f
C804 VTAIL.n62 VSUBS 0.799019f
C805 VTAIL.n63 VSUBS 1.12108f
C806 VTAIL.n64 VSUBS 0.036601f
C807 VTAIL.n65 VSUBS 0.034785f
C808 VTAIL.n66 VSUBS 0.018692f
C809 VTAIL.n67 VSUBS 0.044181f
C810 VTAIL.n68 VSUBS 0.019791f
C811 VTAIL.n69 VSUBS 0.034785f
C812 VTAIL.n70 VSUBS 0.018692f
C813 VTAIL.n71 VSUBS 0.033136f
C814 VTAIL.n72 VSUBS 0.028064f
C815 VTAIL.t9 VSUBS 0.095071f
C816 VTAIL.n73 VSUBS 0.146038f
C817 VTAIL.n74 VSUBS 0.674217f
C818 VTAIL.n75 VSUBS 0.018692f
C819 VTAIL.n76 VSUBS 0.019791f
C820 VTAIL.n77 VSUBS 0.044181f
C821 VTAIL.n78 VSUBS 0.044181f
C822 VTAIL.n79 VSUBS 0.019791f
C823 VTAIL.n80 VSUBS 0.018692f
C824 VTAIL.n81 VSUBS 0.034785f
C825 VTAIL.n82 VSUBS 0.034785f
C826 VTAIL.n83 VSUBS 0.018692f
C827 VTAIL.n84 VSUBS 0.019791f
C828 VTAIL.n85 VSUBS 0.044181f
C829 VTAIL.n86 VSUBS 0.101439f
C830 VTAIL.n87 VSUBS 0.019791f
C831 VTAIL.n88 VSUBS 0.018692f
C832 VTAIL.n89 VSUBS 0.077552f
C833 VTAIL.n90 VSUBS 0.050679f
C834 VTAIL.n91 VSUBS 1.61953f
C835 VTAIL.n92 VSUBS 0.036601f
C836 VTAIL.n93 VSUBS 0.034785f
C837 VTAIL.n94 VSUBS 0.018692f
C838 VTAIL.n95 VSUBS 0.044181f
C839 VTAIL.n96 VSUBS 0.019791f
C840 VTAIL.n97 VSUBS 0.034785f
C841 VTAIL.n98 VSUBS 0.018692f
C842 VTAIL.n99 VSUBS 0.033136f
C843 VTAIL.n100 VSUBS 0.028064f
C844 VTAIL.t0 VSUBS 0.095071f
C845 VTAIL.n101 VSUBS 0.146038f
C846 VTAIL.n102 VSUBS 0.674217f
C847 VTAIL.n103 VSUBS 0.018692f
C848 VTAIL.n104 VSUBS 0.019791f
C849 VTAIL.n105 VSUBS 0.044181f
C850 VTAIL.n106 VSUBS 0.044181f
C851 VTAIL.n107 VSUBS 0.019791f
C852 VTAIL.n108 VSUBS 0.018692f
C853 VTAIL.n109 VSUBS 0.034785f
C854 VTAIL.n110 VSUBS 0.034785f
C855 VTAIL.n111 VSUBS 0.018692f
C856 VTAIL.n112 VSUBS 0.019791f
C857 VTAIL.n113 VSUBS 0.044181f
C858 VTAIL.n114 VSUBS 0.101439f
C859 VTAIL.n115 VSUBS 0.019791f
C860 VTAIL.n116 VSUBS 0.018692f
C861 VTAIL.n117 VSUBS 0.077552f
C862 VTAIL.n118 VSUBS 0.050679f
C863 VTAIL.n119 VSUBS 1.53619f
C864 VDD1.n0 VSUBS 0.02352f
C865 VDD1.n1 VSUBS 0.022352f
C866 VDD1.n2 VSUBS 0.012011f
C867 VDD1.n3 VSUBS 0.02839f
C868 VDD1.n4 VSUBS 0.012718f
C869 VDD1.n5 VSUBS 0.022352f
C870 VDD1.n6 VSUBS 0.012011f
C871 VDD1.n7 VSUBS 0.021293f
C872 VDD1.n8 VSUBS 0.018034f
C873 VDD1.t0 VSUBS 0.061092f
C874 VDD1.n9 VSUBS 0.093842f
C875 VDD1.n10 VSUBS 0.433244f
C876 VDD1.n11 VSUBS 0.012011f
C877 VDD1.n12 VSUBS 0.012718f
C878 VDD1.n13 VSUBS 0.02839f
C879 VDD1.n14 VSUBS 0.02839f
C880 VDD1.n15 VSUBS 0.012718f
C881 VDD1.n16 VSUBS 0.012011f
C882 VDD1.n17 VSUBS 0.022352f
C883 VDD1.n18 VSUBS 0.022352f
C884 VDD1.n19 VSUBS 0.012011f
C885 VDD1.n20 VSUBS 0.012718f
C886 VDD1.n21 VSUBS 0.02839f
C887 VDD1.n22 VSUBS 0.065183f
C888 VDD1.n23 VSUBS 0.012718f
C889 VDD1.n24 VSUBS 0.012011f
C890 VDD1.n25 VSUBS 0.049834f
C891 VDD1.n26 VSUBS 0.05626f
C892 VDD1.n27 VSUBS 0.02352f
C893 VDD1.n28 VSUBS 0.022352f
C894 VDD1.n29 VSUBS 0.012011f
C895 VDD1.n30 VSUBS 0.02839f
C896 VDD1.n31 VSUBS 0.012718f
C897 VDD1.n32 VSUBS 0.022352f
C898 VDD1.n33 VSUBS 0.012011f
C899 VDD1.n34 VSUBS 0.021293f
C900 VDD1.n35 VSUBS 0.018034f
C901 VDD1.t5 VSUBS 0.061092f
C902 VDD1.n36 VSUBS 0.093842f
C903 VDD1.n37 VSUBS 0.433245f
C904 VDD1.n38 VSUBS 0.012011f
C905 VDD1.n39 VSUBS 0.012718f
C906 VDD1.n40 VSUBS 0.02839f
C907 VDD1.n41 VSUBS 0.02839f
C908 VDD1.n42 VSUBS 0.012718f
C909 VDD1.n43 VSUBS 0.012011f
C910 VDD1.n44 VSUBS 0.022352f
C911 VDD1.n45 VSUBS 0.022352f
C912 VDD1.n46 VSUBS 0.012011f
C913 VDD1.n47 VSUBS 0.012718f
C914 VDD1.n48 VSUBS 0.02839f
C915 VDD1.n49 VSUBS 0.065183f
C916 VDD1.n50 VSUBS 0.012718f
C917 VDD1.n51 VSUBS 0.012011f
C918 VDD1.n52 VSUBS 0.049834f
C919 VDD1.n53 VSUBS 0.055516f
C920 VDD1.t3 VSUBS 0.092204f
C921 VDD1.t1 VSUBS 0.092204f
C922 VDD1.n54 VSUBS 0.589589f
C923 VDD1.n55 VSUBS 2.39851f
C924 VDD1.t4 VSUBS 0.092204f
C925 VDD1.t2 VSUBS 0.092204f
C926 VDD1.n56 VSUBS 0.585676f
C927 VDD1.n57 VSUBS 2.25283f
C928 VP.t1 VSUBS 1.56904f
C929 VP.n0 VSUBS 0.749133f
C930 VP.n1 VSUBS 0.040201f
C931 VP.n2 VSUBS 0.06835f
C932 VP.n3 VSUBS 0.040201f
C933 VP.t0 VSUBS 1.56904f
C934 VP.n4 VSUBS 0.074549f
C935 VP.n5 VSUBS 0.040201f
C936 VP.n6 VSUBS 0.069396f
C937 VP.t2 VSUBS 1.56904f
C938 VP.n7 VSUBS 0.749133f
C939 VP.n8 VSUBS 0.040201f
C940 VP.n9 VSUBS 0.06835f
C941 VP.n10 VSUBS 0.426952f
C942 VP.t4 VSUBS 1.56904f
C943 VP.t3 VSUBS 1.92753f
C944 VP.n11 VSUBS 0.692675f
C945 VP.n12 VSUBS 0.719045f
C946 VP.n13 VSUBS 0.056147f
C947 VP.n14 VSUBS 0.074549f
C948 VP.n15 VSUBS 0.040201f
C949 VP.n16 VSUBS 0.040201f
C950 VP.n17 VSUBS 0.040201f
C951 VP.n18 VSUBS 0.04783f
C952 VP.n19 VSUBS 0.075245f
C953 VP.n20 VSUBS 0.069396f
C954 VP.n21 VSUBS 0.064873f
C955 VP.n22 VSUBS 1.91316f
C956 VP.t5 VSUBS 1.56904f
C957 VP.n23 VSUBS 0.749133f
C958 VP.n24 VSUBS 1.94564f
C959 VP.n25 VSUBS 0.064873f
C960 VP.n26 VSUBS 0.040201f
C961 VP.n27 VSUBS 0.075245f
C962 VP.n28 VSUBS 0.04783f
C963 VP.n29 VSUBS 0.06835f
C964 VP.n30 VSUBS 0.040201f
C965 VP.n31 VSUBS 0.040201f
C966 VP.n32 VSUBS 0.040201f
C967 VP.n33 VSUBS 0.056147f
C968 VP.n34 VSUBS 0.595491f
C969 VP.n35 VSUBS 0.056147f
C970 VP.n36 VSUBS 0.074549f
C971 VP.n37 VSUBS 0.040201f
C972 VP.n38 VSUBS 0.040201f
C973 VP.n39 VSUBS 0.040201f
C974 VP.n40 VSUBS 0.04783f
C975 VP.n41 VSUBS 0.075245f
C976 VP.n42 VSUBS 0.069396f
C977 VP.n43 VSUBS 0.064873f
C978 VP.n44 VSUBS 0.079795f
.ends

