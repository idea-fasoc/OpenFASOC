* NGSPICE file created from diff_pair_sample_1583.ext - technology: sky130A

.subckt diff_pair_sample_1583 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=2.0982 pd=11.54 as=0 ps=0 w=5.38 l=2.43
X1 VDD1.t9 VP.t0 VTAIL.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=2.0982 ps=11.54 w=5.38 l=2.43
X2 VDD1.t8 VP.t1 VTAIL.t19 B.t2 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=2.0982 ps=11.54 w=5.38 l=2.43
X3 VTAIL.t17 VP.t2 VDD1.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=0.8877 ps=5.71 w=5.38 l=2.43
X4 VDD2.t9 VN.t0 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=0.8877 ps=5.71 w=5.38 l=2.43
X5 VDD2.t8 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=0.8877 ps=5.71 w=5.38 l=2.43
X6 VDD1.t6 VP.t3 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=2.0982 pd=11.54 as=0.8877 ps=5.71 w=5.38 l=2.43
X7 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=2.0982 pd=11.54 as=0 ps=0 w=5.38 l=2.43
X8 VTAIL.t5 VN.t2 VDD2.t7 B.t8 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=0.8877 ps=5.71 w=5.38 l=2.43
X9 VTAIL.t18 VP.t4 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=0.8877 ps=5.71 w=5.38 l=2.43
X10 VDD2.t6 VN.t3 VTAIL.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=2.0982 pd=11.54 as=0.8877 ps=5.71 w=5.38 l=2.43
X11 VTAIL.t9 VN.t4 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=0.8877 ps=5.71 w=5.38 l=2.43
X12 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=2.0982 pd=11.54 as=0 ps=0 w=5.38 l=2.43
X13 VTAIL.t12 VP.t5 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=0.8877 ps=5.71 w=5.38 l=2.43
X14 VDD1.t3 VP.t6 VTAIL.t15 B.t6 sky130_fd_pr__nfet_01v8 ad=2.0982 pd=11.54 as=0.8877 ps=5.71 w=5.38 l=2.43
X15 VDD2.t4 VN.t5 VTAIL.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=2.0982 pd=11.54 as=0.8877 ps=5.71 w=5.38 l=2.43
X16 VDD2.t3 VN.t6 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=2.0982 ps=11.54 w=5.38 l=2.43
X17 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.0982 pd=11.54 as=0 ps=0 w=5.38 l=2.43
X18 VDD1.t2 VP.t7 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=0.8877 ps=5.71 w=5.38 l=2.43
X19 VTAIL.t1 VN.t7 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=0.8877 ps=5.71 w=5.38 l=2.43
X20 VTAIL.t7 VN.t8 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=0.8877 ps=5.71 w=5.38 l=2.43
X21 VDD2.t0 VN.t9 VTAIL.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=2.0982 ps=11.54 w=5.38 l=2.43
X22 VTAIL.t16 VP.t8 VDD1.t1 B.t8 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=0.8877 ps=5.71 w=5.38 l=2.43
X23 VDD1.t0 VP.t9 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=0.8877 pd=5.71 as=0.8877 ps=5.71 w=5.38 l=2.43
R0 B.n739 B.n738 585
R1 B.n242 B.n131 585
R2 B.n241 B.n240 585
R3 B.n239 B.n238 585
R4 B.n237 B.n236 585
R5 B.n235 B.n234 585
R6 B.n233 B.n232 585
R7 B.n231 B.n230 585
R8 B.n229 B.n228 585
R9 B.n227 B.n226 585
R10 B.n225 B.n224 585
R11 B.n223 B.n222 585
R12 B.n221 B.n220 585
R13 B.n219 B.n218 585
R14 B.n217 B.n216 585
R15 B.n215 B.n214 585
R16 B.n213 B.n212 585
R17 B.n211 B.n210 585
R18 B.n209 B.n208 585
R19 B.n207 B.n206 585
R20 B.n205 B.n204 585
R21 B.n203 B.n202 585
R22 B.n201 B.n200 585
R23 B.n199 B.n198 585
R24 B.n197 B.n196 585
R25 B.n195 B.n194 585
R26 B.n193 B.n192 585
R27 B.n191 B.n190 585
R28 B.n189 B.n188 585
R29 B.n187 B.n186 585
R30 B.n185 B.n184 585
R31 B.n183 B.n182 585
R32 B.n181 B.n180 585
R33 B.n179 B.n178 585
R34 B.n177 B.n176 585
R35 B.n175 B.n174 585
R36 B.n173 B.n172 585
R37 B.n171 B.n170 585
R38 B.n169 B.n168 585
R39 B.n167 B.n166 585
R40 B.n165 B.n164 585
R41 B.n163 B.n162 585
R42 B.n161 B.n160 585
R43 B.n159 B.n158 585
R44 B.n157 B.n156 585
R45 B.n155 B.n154 585
R46 B.n153 B.n152 585
R47 B.n151 B.n150 585
R48 B.n149 B.n148 585
R49 B.n147 B.n146 585
R50 B.n145 B.n144 585
R51 B.n143 B.n142 585
R52 B.n141 B.n140 585
R53 B.n139 B.n138 585
R54 B.n737 B.n104 585
R55 B.n742 B.n104 585
R56 B.n736 B.n103 585
R57 B.n743 B.n103 585
R58 B.n735 B.n734 585
R59 B.n734 B.n99 585
R60 B.n733 B.n98 585
R61 B.n749 B.n98 585
R62 B.n732 B.n97 585
R63 B.n750 B.n97 585
R64 B.n731 B.n96 585
R65 B.n751 B.n96 585
R66 B.n730 B.n729 585
R67 B.n729 B.n92 585
R68 B.n728 B.n91 585
R69 B.n757 B.n91 585
R70 B.n727 B.n90 585
R71 B.n758 B.n90 585
R72 B.n726 B.n89 585
R73 B.n759 B.n89 585
R74 B.n725 B.n724 585
R75 B.n724 B.n85 585
R76 B.n723 B.n84 585
R77 B.n765 B.n84 585
R78 B.n722 B.n83 585
R79 B.n766 B.n83 585
R80 B.n721 B.n82 585
R81 B.n767 B.n82 585
R82 B.n720 B.n719 585
R83 B.n719 B.n78 585
R84 B.n718 B.n77 585
R85 B.n773 B.n77 585
R86 B.n717 B.n76 585
R87 B.n774 B.n76 585
R88 B.n716 B.n75 585
R89 B.n775 B.n75 585
R90 B.n715 B.n714 585
R91 B.n714 B.n74 585
R92 B.n713 B.n70 585
R93 B.n781 B.n70 585
R94 B.n712 B.n69 585
R95 B.n782 B.n69 585
R96 B.n711 B.n68 585
R97 B.n783 B.n68 585
R98 B.n710 B.n709 585
R99 B.n709 B.n64 585
R100 B.n708 B.n63 585
R101 B.n789 B.n63 585
R102 B.n707 B.n62 585
R103 B.n790 B.n62 585
R104 B.n706 B.n61 585
R105 B.n791 B.n61 585
R106 B.n705 B.n704 585
R107 B.n704 B.n60 585
R108 B.n703 B.n56 585
R109 B.n797 B.n56 585
R110 B.n702 B.n55 585
R111 B.n798 B.n55 585
R112 B.n701 B.n54 585
R113 B.n799 B.n54 585
R114 B.n700 B.n699 585
R115 B.n699 B.n50 585
R116 B.n698 B.n49 585
R117 B.n805 B.n49 585
R118 B.n697 B.n48 585
R119 B.n806 B.n48 585
R120 B.n696 B.n47 585
R121 B.n807 B.n47 585
R122 B.n695 B.n694 585
R123 B.n694 B.n43 585
R124 B.n693 B.n42 585
R125 B.n813 B.n42 585
R126 B.n692 B.n41 585
R127 B.n814 B.n41 585
R128 B.n691 B.n40 585
R129 B.n815 B.n40 585
R130 B.n690 B.n689 585
R131 B.n689 B.n36 585
R132 B.n688 B.n35 585
R133 B.n821 B.n35 585
R134 B.n687 B.n34 585
R135 B.n822 B.n34 585
R136 B.n686 B.n33 585
R137 B.n823 B.n33 585
R138 B.n685 B.n684 585
R139 B.n684 B.n29 585
R140 B.n683 B.n28 585
R141 B.n829 B.n28 585
R142 B.n682 B.n27 585
R143 B.n830 B.n27 585
R144 B.n681 B.n26 585
R145 B.n831 B.n26 585
R146 B.n680 B.n679 585
R147 B.n679 B.n22 585
R148 B.n678 B.n21 585
R149 B.n837 B.n21 585
R150 B.n677 B.n20 585
R151 B.n838 B.n20 585
R152 B.n676 B.n19 585
R153 B.n839 B.n19 585
R154 B.n675 B.n674 585
R155 B.n674 B.n15 585
R156 B.n673 B.n14 585
R157 B.n845 B.n14 585
R158 B.n672 B.n13 585
R159 B.n846 B.n13 585
R160 B.n671 B.n12 585
R161 B.n847 B.n12 585
R162 B.n670 B.n669 585
R163 B.n669 B.n8 585
R164 B.n668 B.n7 585
R165 B.n853 B.n7 585
R166 B.n667 B.n6 585
R167 B.n854 B.n6 585
R168 B.n666 B.n5 585
R169 B.n855 B.n5 585
R170 B.n665 B.n664 585
R171 B.n664 B.n4 585
R172 B.n663 B.n243 585
R173 B.n663 B.n662 585
R174 B.n653 B.n244 585
R175 B.n245 B.n244 585
R176 B.n655 B.n654 585
R177 B.n656 B.n655 585
R178 B.n652 B.n250 585
R179 B.n250 B.n249 585
R180 B.n651 B.n650 585
R181 B.n650 B.n649 585
R182 B.n252 B.n251 585
R183 B.n253 B.n252 585
R184 B.n642 B.n641 585
R185 B.n643 B.n642 585
R186 B.n640 B.n258 585
R187 B.n258 B.n257 585
R188 B.n639 B.n638 585
R189 B.n638 B.n637 585
R190 B.n260 B.n259 585
R191 B.n261 B.n260 585
R192 B.n630 B.n629 585
R193 B.n631 B.n630 585
R194 B.n628 B.n266 585
R195 B.n266 B.n265 585
R196 B.n627 B.n626 585
R197 B.n626 B.n625 585
R198 B.n268 B.n267 585
R199 B.n269 B.n268 585
R200 B.n618 B.n617 585
R201 B.n619 B.n618 585
R202 B.n616 B.n274 585
R203 B.n274 B.n273 585
R204 B.n615 B.n614 585
R205 B.n614 B.n613 585
R206 B.n276 B.n275 585
R207 B.n277 B.n276 585
R208 B.n606 B.n605 585
R209 B.n607 B.n606 585
R210 B.n604 B.n282 585
R211 B.n282 B.n281 585
R212 B.n603 B.n602 585
R213 B.n602 B.n601 585
R214 B.n284 B.n283 585
R215 B.n285 B.n284 585
R216 B.n594 B.n593 585
R217 B.n595 B.n594 585
R218 B.n592 B.n290 585
R219 B.n290 B.n289 585
R220 B.n591 B.n590 585
R221 B.n590 B.n589 585
R222 B.n292 B.n291 585
R223 B.n293 B.n292 585
R224 B.n582 B.n581 585
R225 B.n583 B.n582 585
R226 B.n580 B.n298 585
R227 B.n298 B.n297 585
R228 B.n579 B.n578 585
R229 B.n578 B.n577 585
R230 B.n300 B.n299 585
R231 B.n570 B.n300 585
R232 B.n569 B.n568 585
R233 B.n571 B.n569 585
R234 B.n567 B.n305 585
R235 B.n305 B.n304 585
R236 B.n566 B.n565 585
R237 B.n565 B.n564 585
R238 B.n307 B.n306 585
R239 B.n308 B.n307 585
R240 B.n557 B.n556 585
R241 B.n558 B.n557 585
R242 B.n555 B.n313 585
R243 B.n313 B.n312 585
R244 B.n554 B.n553 585
R245 B.n553 B.n552 585
R246 B.n315 B.n314 585
R247 B.n545 B.n315 585
R248 B.n544 B.n543 585
R249 B.n546 B.n544 585
R250 B.n542 B.n320 585
R251 B.n320 B.n319 585
R252 B.n541 B.n540 585
R253 B.n540 B.n539 585
R254 B.n322 B.n321 585
R255 B.n323 B.n322 585
R256 B.n532 B.n531 585
R257 B.n533 B.n532 585
R258 B.n530 B.n328 585
R259 B.n328 B.n327 585
R260 B.n529 B.n528 585
R261 B.n528 B.n527 585
R262 B.n330 B.n329 585
R263 B.n331 B.n330 585
R264 B.n520 B.n519 585
R265 B.n521 B.n520 585
R266 B.n518 B.n336 585
R267 B.n336 B.n335 585
R268 B.n517 B.n516 585
R269 B.n516 B.n515 585
R270 B.n338 B.n337 585
R271 B.n339 B.n338 585
R272 B.n508 B.n507 585
R273 B.n509 B.n508 585
R274 B.n506 B.n344 585
R275 B.n344 B.n343 585
R276 B.n505 B.n504 585
R277 B.n504 B.n503 585
R278 B.n346 B.n345 585
R279 B.n347 B.n346 585
R280 B.n496 B.n495 585
R281 B.n497 B.n496 585
R282 B.n494 B.n352 585
R283 B.n352 B.n351 585
R284 B.n489 B.n488 585
R285 B.n487 B.n381 585
R286 B.n486 B.n380 585
R287 B.n491 B.n380 585
R288 B.n485 B.n484 585
R289 B.n483 B.n482 585
R290 B.n481 B.n480 585
R291 B.n479 B.n478 585
R292 B.n477 B.n476 585
R293 B.n475 B.n474 585
R294 B.n473 B.n472 585
R295 B.n471 B.n470 585
R296 B.n469 B.n468 585
R297 B.n467 B.n466 585
R298 B.n465 B.n464 585
R299 B.n463 B.n462 585
R300 B.n461 B.n460 585
R301 B.n459 B.n458 585
R302 B.n457 B.n456 585
R303 B.n455 B.n454 585
R304 B.n453 B.n452 585
R305 B.n451 B.n450 585
R306 B.n449 B.n448 585
R307 B.n446 B.n445 585
R308 B.n444 B.n443 585
R309 B.n442 B.n441 585
R310 B.n440 B.n439 585
R311 B.n438 B.n437 585
R312 B.n436 B.n435 585
R313 B.n434 B.n433 585
R314 B.n432 B.n431 585
R315 B.n430 B.n429 585
R316 B.n428 B.n427 585
R317 B.n425 B.n424 585
R318 B.n423 B.n422 585
R319 B.n421 B.n420 585
R320 B.n419 B.n418 585
R321 B.n417 B.n416 585
R322 B.n415 B.n414 585
R323 B.n413 B.n412 585
R324 B.n411 B.n410 585
R325 B.n409 B.n408 585
R326 B.n407 B.n406 585
R327 B.n405 B.n404 585
R328 B.n403 B.n402 585
R329 B.n401 B.n400 585
R330 B.n399 B.n398 585
R331 B.n397 B.n396 585
R332 B.n395 B.n394 585
R333 B.n393 B.n392 585
R334 B.n391 B.n390 585
R335 B.n389 B.n388 585
R336 B.n387 B.n386 585
R337 B.n354 B.n353 585
R338 B.n493 B.n492 585
R339 B.n492 B.n491 585
R340 B.n350 B.n349 585
R341 B.n351 B.n350 585
R342 B.n499 B.n498 585
R343 B.n498 B.n497 585
R344 B.n500 B.n348 585
R345 B.n348 B.n347 585
R346 B.n502 B.n501 585
R347 B.n503 B.n502 585
R348 B.n342 B.n341 585
R349 B.n343 B.n342 585
R350 B.n511 B.n510 585
R351 B.n510 B.n509 585
R352 B.n512 B.n340 585
R353 B.n340 B.n339 585
R354 B.n514 B.n513 585
R355 B.n515 B.n514 585
R356 B.n334 B.n333 585
R357 B.n335 B.n334 585
R358 B.n523 B.n522 585
R359 B.n522 B.n521 585
R360 B.n524 B.n332 585
R361 B.n332 B.n331 585
R362 B.n526 B.n525 585
R363 B.n527 B.n526 585
R364 B.n326 B.n325 585
R365 B.n327 B.n326 585
R366 B.n535 B.n534 585
R367 B.n534 B.n533 585
R368 B.n536 B.n324 585
R369 B.n324 B.n323 585
R370 B.n538 B.n537 585
R371 B.n539 B.n538 585
R372 B.n318 B.n317 585
R373 B.n319 B.n318 585
R374 B.n548 B.n547 585
R375 B.n547 B.n546 585
R376 B.n549 B.n316 585
R377 B.n545 B.n316 585
R378 B.n551 B.n550 585
R379 B.n552 B.n551 585
R380 B.n311 B.n310 585
R381 B.n312 B.n311 585
R382 B.n560 B.n559 585
R383 B.n559 B.n558 585
R384 B.n561 B.n309 585
R385 B.n309 B.n308 585
R386 B.n563 B.n562 585
R387 B.n564 B.n563 585
R388 B.n303 B.n302 585
R389 B.n304 B.n303 585
R390 B.n573 B.n572 585
R391 B.n572 B.n571 585
R392 B.n574 B.n301 585
R393 B.n570 B.n301 585
R394 B.n576 B.n575 585
R395 B.n577 B.n576 585
R396 B.n296 B.n295 585
R397 B.n297 B.n296 585
R398 B.n585 B.n584 585
R399 B.n584 B.n583 585
R400 B.n586 B.n294 585
R401 B.n294 B.n293 585
R402 B.n588 B.n587 585
R403 B.n589 B.n588 585
R404 B.n288 B.n287 585
R405 B.n289 B.n288 585
R406 B.n597 B.n596 585
R407 B.n596 B.n595 585
R408 B.n598 B.n286 585
R409 B.n286 B.n285 585
R410 B.n600 B.n599 585
R411 B.n601 B.n600 585
R412 B.n280 B.n279 585
R413 B.n281 B.n280 585
R414 B.n609 B.n608 585
R415 B.n608 B.n607 585
R416 B.n610 B.n278 585
R417 B.n278 B.n277 585
R418 B.n612 B.n611 585
R419 B.n613 B.n612 585
R420 B.n272 B.n271 585
R421 B.n273 B.n272 585
R422 B.n621 B.n620 585
R423 B.n620 B.n619 585
R424 B.n622 B.n270 585
R425 B.n270 B.n269 585
R426 B.n624 B.n623 585
R427 B.n625 B.n624 585
R428 B.n264 B.n263 585
R429 B.n265 B.n264 585
R430 B.n633 B.n632 585
R431 B.n632 B.n631 585
R432 B.n634 B.n262 585
R433 B.n262 B.n261 585
R434 B.n636 B.n635 585
R435 B.n637 B.n636 585
R436 B.n256 B.n255 585
R437 B.n257 B.n256 585
R438 B.n645 B.n644 585
R439 B.n644 B.n643 585
R440 B.n646 B.n254 585
R441 B.n254 B.n253 585
R442 B.n648 B.n647 585
R443 B.n649 B.n648 585
R444 B.n248 B.n247 585
R445 B.n249 B.n248 585
R446 B.n658 B.n657 585
R447 B.n657 B.n656 585
R448 B.n659 B.n246 585
R449 B.n246 B.n245 585
R450 B.n661 B.n660 585
R451 B.n662 B.n661 585
R452 B.n2 B.n0 585
R453 B.n4 B.n2 585
R454 B.n3 B.n1 585
R455 B.n854 B.n3 585
R456 B.n852 B.n851 585
R457 B.n853 B.n852 585
R458 B.n850 B.n9 585
R459 B.n9 B.n8 585
R460 B.n849 B.n848 585
R461 B.n848 B.n847 585
R462 B.n11 B.n10 585
R463 B.n846 B.n11 585
R464 B.n844 B.n843 585
R465 B.n845 B.n844 585
R466 B.n842 B.n16 585
R467 B.n16 B.n15 585
R468 B.n841 B.n840 585
R469 B.n840 B.n839 585
R470 B.n18 B.n17 585
R471 B.n838 B.n18 585
R472 B.n836 B.n835 585
R473 B.n837 B.n836 585
R474 B.n834 B.n23 585
R475 B.n23 B.n22 585
R476 B.n833 B.n832 585
R477 B.n832 B.n831 585
R478 B.n25 B.n24 585
R479 B.n830 B.n25 585
R480 B.n828 B.n827 585
R481 B.n829 B.n828 585
R482 B.n826 B.n30 585
R483 B.n30 B.n29 585
R484 B.n825 B.n824 585
R485 B.n824 B.n823 585
R486 B.n32 B.n31 585
R487 B.n822 B.n32 585
R488 B.n820 B.n819 585
R489 B.n821 B.n820 585
R490 B.n818 B.n37 585
R491 B.n37 B.n36 585
R492 B.n817 B.n816 585
R493 B.n816 B.n815 585
R494 B.n39 B.n38 585
R495 B.n814 B.n39 585
R496 B.n812 B.n811 585
R497 B.n813 B.n812 585
R498 B.n810 B.n44 585
R499 B.n44 B.n43 585
R500 B.n809 B.n808 585
R501 B.n808 B.n807 585
R502 B.n46 B.n45 585
R503 B.n806 B.n46 585
R504 B.n804 B.n803 585
R505 B.n805 B.n804 585
R506 B.n802 B.n51 585
R507 B.n51 B.n50 585
R508 B.n801 B.n800 585
R509 B.n800 B.n799 585
R510 B.n53 B.n52 585
R511 B.n798 B.n53 585
R512 B.n796 B.n795 585
R513 B.n797 B.n796 585
R514 B.n794 B.n57 585
R515 B.n60 B.n57 585
R516 B.n793 B.n792 585
R517 B.n792 B.n791 585
R518 B.n59 B.n58 585
R519 B.n790 B.n59 585
R520 B.n788 B.n787 585
R521 B.n789 B.n788 585
R522 B.n786 B.n65 585
R523 B.n65 B.n64 585
R524 B.n785 B.n784 585
R525 B.n784 B.n783 585
R526 B.n67 B.n66 585
R527 B.n782 B.n67 585
R528 B.n780 B.n779 585
R529 B.n781 B.n780 585
R530 B.n778 B.n71 585
R531 B.n74 B.n71 585
R532 B.n777 B.n776 585
R533 B.n776 B.n775 585
R534 B.n73 B.n72 585
R535 B.n774 B.n73 585
R536 B.n772 B.n771 585
R537 B.n773 B.n772 585
R538 B.n770 B.n79 585
R539 B.n79 B.n78 585
R540 B.n769 B.n768 585
R541 B.n768 B.n767 585
R542 B.n81 B.n80 585
R543 B.n766 B.n81 585
R544 B.n764 B.n763 585
R545 B.n765 B.n764 585
R546 B.n762 B.n86 585
R547 B.n86 B.n85 585
R548 B.n761 B.n760 585
R549 B.n760 B.n759 585
R550 B.n88 B.n87 585
R551 B.n758 B.n88 585
R552 B.n756 B.n755 585
R553 B.n757 B.n756 585
R554 B.n754 B.n93 585
R555 B.n93 B.n92 585
R556 B.n753 B.n752 585
R557 B.n752 B.n751 585
R558 B.n95 B.n94 585
R559 B.n750 B.n95 585
R560 B.n748 B.n747 585
R561 B.n749 B.n748 585
R562 B.n746 B.n100 585
R563 B.n100 B.n99 585
R564 B.n745 B.n744 585
R565 B.n744 B.n743 585
R566 B.n102 B.n101 585
R567 B.n742 B.n102 585
R568 B.n857 B.n856 585
R569 B.n856 B.n855 585
R570 B.n489 B.n350 458.866
R571 B.n138 B.n102 458.866
R572 B.n492 B.n352 458.866
R573 B.n739 B.n104 458.866
R574 B.n384 B.t21 261.132
R575 B.n382 B.t14 261.132
R576 B.n135 B.t18 261.132
R577 B.n132 B.t10 261.132
R578 B.n741 B.n740 256.663
R579 B.n741 B.n130 256.663
R580 B.n741 B.n129 256.663
R581 B.n741 B.n128 256.663
R582 B.n741 B.n127 256.663
R583 B.n741 B.n126 256.663
R584 B.n741 B.n125 256.663
R585 B.n741 B.n124 256.663
R586 B.n741 B.n123 256.663
R587 B.n741 B.n122 256.663
R588 B.n741 B.n121 256.663
R589 B.n741 B.n120 256.663
R590 B.n741 B.n119 256.663
R591 B.n741 B.n118 256.663
R592 B.n741 B.n117 256.663
R593 B.n741 B.n116 256.663
R594 B.n741 B.n115 256.663
R595 B.n741 B.n114 256.663
R596 B.n741 B.n113 256.663
R597 B.n741 B.n112 256.663
R598 B.n741 B.n111 256.663
R599 B.n741 B.n110 256.663
R600 B.n741 B.n109 256.663
R601 B.n741 B.n108 256.663
R602 B.n741 B.n107 256.663
R603 B.n741 B.n106 256.663
R604 B.n741 B.n105 256.663
R605 B.n491 B.n490 256.663
R606 B.n491 B.n355 256.663
R607 B.n491 B.n356 256.663
R608 B.n491 B.n357 256.663
R609 B.n491 B.n358 256.663
R610 B.n491 B.n359 256.663
R611 B.n491 B.n360 256.663
R612 B.n491 B.n361 256.663
R613 B.n491 B.n362 256.663
R614 B.n491 B.n363 256.663
R615 B.n491 B.n364 256.663
R616 B.n491 B.n365 256.663
R617 B.n491 B.n366 256.663
R618 B.n491 B.n367 256.663
R619 B.n491 B.n368 256.663
R620 B.n491 B.n369 256.663
R621 B.n491 B.n370 256.663
R622 B.n491 B.n371 256.663
R623 B.n491 B.n372 256.663
R624 B.n491 B.n373 256.663
R625 B.n491 B.n374 256.663
R626 B.n491 B.n375 256.663
R627 B.n491 B.n376 256.663
R628 B.n491 B.n377 256.663
R629 B.n491 B.n378 256.663
R630 B.n491 B.n379 256.663
R631 B.n384 B.t23 222.041
R632 B.n132 B.t12 222.041
R633 B.n382 B.t17 222.041
R634 B.n135 B.t19 222.041
R635 B.n385 B.t22 168.513
R636 B.n133 B.t13 168.513
R637 B.n383 B.t16 168.513
R638 B.n136 B.t20 168.513
R639 B.n498 B.n350 163.367
R640 B.n498 B.n348 163.367
R641 B.n502 B.n348 163.367
R642 B.n502 B.n342 163.367
R643 B.n510 B.n342 163.367
R644 B.n510 B.n340 163.367
R645 B.n514 B.n340 163.367
R646 B.n514 B.n334 163.367
R647 B.n522 B.n334 163.367
R648 B.n522 B.n332 163.367
R649 B.n526 B.n332 163.367
R650 B.n526 B.n326 163.367
R651 B.n534 B.n326 163.367
R652 B.n534 B.n324 163.367
R653 B.n538 B.n324 163.367
R654 B.n538 B.n318 163.367
R655 B.n547 B.n318 163.367
R656 B.n547 B.n316 163.367
R657 B.n551 B.n316 163.367
R658 B.n551 B.n311 163.367
R659 B.n559 B.n311 163.367
R660 B.n559 B.n309 163.367
R661 B.n563 B.n309 163.367
R662 B.n563 B.n303 163.367
R663 B.n572 B.n303 163.367
R664 B.n572 B.n301 163.367
R665 B.n576 B.n301 163.367
R666 B.n576 B.n296 163.367
R667 B.n584 B.n296 163.367
R668 B.n584 B.n294 163.367
R669 B.n588 B.n294 163.367
R670 B.n588 B.n288 163.367
R671 B.n596 B.n288 163.367
R672 B.n596 B.n286 163.367
R673 B.n600 B.n286 163.367
R674 B.n600 B.n280 163.367
R675 B.n608 B.n280 163.367
R676 B.n608 B.n278 163.367
R677 B.n612 B.n278 163.367
R678 B.n612 B.n272 163.367
R679 B.n620 B.n272 163.367
R680 B.n620 B.n270 163.367
R681 B.n624 B.n270 163.367
R682 B.n624 B.n264 163.367
R683 B.n632 B.n264 163.367
R684 B.n632 B.n262 163.367
R685 B.n636 B.n262 163.367
R686 B.n636 B.n256 163.367
R687 B.n644 B.n256 163.367
R688 B.n644 B.n254 163.367
R689 B.n648 B.n254 163.367
R690 B.n648 B.n248 163.367
R691 B.n657 B.n248 163.367
R692 B.n657 B.n246 163.367
R693 B.n661 B.n246 163.367
R694 B.n661 B.n2 163.367
R695 B.n856 B.n2 163.367
R696 B.n856 B.n3 163.367
R697 B.n852 B.n3 163.367
R698 B.n852 B.n9 163.367
R699 B.n848 B.n9 163.367
R700 B.n848 B.n11 163.367
R701 B.n844 B.n11 163.367
R702 B.n844 B.n16 163.367
R703 B.n840 B.n16 163.367
R704 B.n840 B.n18 163.367
R705 B.n836 B.n18 163.367
R706 B.n836 B.n23 163.367
R707 B.n832 B.n23 163.367
R708 B.n832 B.n25 163.367
R709 B.n828 B.n25 163.367
R710 B.n828 B.n30 163.367
R711 B.n824 B.n30 163.367
R712 B.n824 B.n32 163.367
R713 B.n820 B.n32 163.367
R714 B.n820 B.n37 163.367
R715 B.n816 B.n37 163.367
R716 B.n816 B.n39 163.367
R717 B.n812 B.n39 163.367
R718 B.n812 B.n44 163.367
R719 B.n808 B.n44 163.367
R720 B.n808 B.n46 163.367
R721 B.n804 B.n46 163.367
R722 B.n804 B.n51 163.367
R723 B.n800 B.n51 163.367
R724 B.n800 B.n53 163.367
R725 B.n796 B.n53 163.367
R726 B.n796 B.n57 163.367
R727 B.n792 B.n57 163.367
R728 B.n792 B.n59 163.367
R729 B.n788 B.n59 163.367
R730 B.n788 B.n65 163.367
R731 B.n784 B.n65 163.367
R732 B.n784 B.n67 163.367
R733 B.n780 B.n67 163.367
R734 B.n780 B.n71 163.367
R735 B.n776 B.n71 163.367
R736 B.n776 B.n73 163.367
R737 B.n772 B.n73 163.367
R738 B.n772 B.n79 163.367
R739 B.n768 B.n79 163.367
R740 B.n768 B.n81 163.367
R741 B.n764 B.n81 163.367
R742 B.n764 B.n86 163.367
R743 B.n760 B.n86 163.367
R744 B.n760 B.n88 163.367
R745 B.n756 B.n88 163.367
R746 B.n756 B.n93 163.367
R747 B.n752 B.n93 163.367
R748 B.n752 B.n95 163.367
R749 B.n748 B.n95 163.367
R750 B.n748 B.n100 163.367
R751 B.n744 B.n100 163.367
R752 B.n744 B.n102 163.367
R753 B.n381 B.n380 163.367
R754 B.n484 B.n380 163.367
R755 B.n482 B.n481 163.367
R756 B.n478 B.n477 163.367
R757 B.n474 B.n473 163.367
R758 B.n470 B.n469 163.367
R759 B.n466 B.n465 163.367
R760 B.n462 B.n461 163.367
R761 B.n458 B.n457 163.367
R762 B.n454 B.n453 163.367
R763 B.n450 B.n449 163.367
R764 B.n445 B.n444 163.367
R765 B.n441 B.n440 163.367
R766 B.n437 B.n436 163.367
R767 B.n433 B.n432 163.367
R768 B.n429 B.n428 163.367
R769 B.n424 B.n423 163.367
R770 B.n420 B.n419 163.367
R771 B.n416 B.n415 163.367
R772 B.n412 B.n411 163.367
R773 B.n408 B.n407 163.367
R774 B.n404 B.n403 163.367
R775 B.n400 B.n399 163.367
R776 B.n396 B.n395 163.367
R777 B.n392 B.n391 163.367
R778 B.n388 B.n387 163.367
R779 B.n492 B.n354 163.367
R780 B.n496 B.n352 163.367
R781 B.n496 B.n346 163.367
R782 B.n504 B.n346 163.367
R783 B.n504 B.n344 163.367
R784 B.n508 B.n344 163.367
R785 B.n508 B.n338 163.367
R786 B.n516 B.n338 163.367
R787 B.n516 B.n336 163.367
R788 B.n520 B.n336 163.367
R789 B.n520 B.n330 163.367
R790 B.n528 B.n330 163.367
R791 B.n528 B.n328 163.367
R792 B.n532 B.n328 163.367
R793 B.n532 B.n322 163.367
R794 B.n540 B.n322 163.367
R795 B.n540 B.n320 163.367
R796 B.n544 B.n320 163.367
R797 B.n544 B.n315 163.367
R798 B.n553 B.n315 163.367
R799 B.n553 B.n313 163.367
R800 B.n557 B.n313 163.367
R801 B.n557 B.n307 163.367
R802 B.n565 B.n307 163.367
R803 B.n565 B.n305 163.367
R804 B.n569 B.n305 163.367
R805 B.n569 B.n300 163.367
R806 B.n578 B.n300 163.367
R807 B.n578 B.n298 163.367
R808 B.n582 B.n298 163.367
R809 B.n582 B.n292 163.367
R810 B.n590 B.n292 163.367
R811 B.n590 B.n290 163.367
R812 B.n594 B.n290 163.367
R813 B.n594 B.n284 163.367
R814 B.n602 B.n284 163.367
R815 B.n602 B.n282 163.367
R816 B.n606 B.n282 163.367
R817 B.n606 B.n276 163.367
R818 B.n614 B.n276 163.367
R819 B.n614 B.n274 163.367
R820 B.n618 B.n274 163.367
R821 B.n618 B.n268 163.367
R822 B.n626 B.n268 163.367
R823 B.n626 B.n266 163.367
R824 B.n630 B.n266 163.367
R825 B.n630 B.n260 163.367
R826 B.n638 B.n260 163.367
R827 B.n638 B.n258 163.367
R828 B.n642 B.n258 163.367
R829 B.n642 B.n252 163.367
R830 B.n650 B.n252 163.367
R831 B.n650 B.n250 163.367
R832 B.n655 B.n250 163.367
R833 B.n655 B.n244 163.367
R834 B.n663 B.n244 163.367
R835 B.n664 B.n663 163.367
R836 B.n664 B.n5 163.367
R837 B.n6 B.n5 163.367
R838 B.n7 B.n6 163.367
R839 B.n669 B.n7 163.367
R840 B.n669 B.n12 163.367
R841 B.n13 B.n12 163.367
R842 B.n14 B.n13 163.367
R843 B.n674 B.n14 163.367
R844 B.n674 B.n19 163.367
R845 B.n20 B.n19 163.367
R846 B.n21 B.n20 163.367
R847 B.n679 B.n21 163.367
R848 B.n679 B.n26 163.367
R849 B.n27 B.n26 163.367
R850 B.n28 B.n27 163.367
R851 B.n684 B.n28 163.367
R852 B.n684 B.n33 163.367
R853 B.n34 B.n33 163.367
R854 B.n35 B.n34 163.367
R855 B.n689 B.n35 163.367
R856 B.n689 B.n40 163.367
R857 B.n41 B.n40 163.367
R858 B.n42 B.n41 163.367
R859 B.n694 B.n42 163.367
R860 B.n694 B.n47 163.367
R861 B.n48 B.n47 163.367
R862 B.n49 B.n48 163.367
R863 B.n699 B.n49 163.367
R864 B.n699 B.n54 163.367
R865 B.n55 B.n54 163.367
R866 B.n56 B.n55 163.367
R867 B.n704 B.n56 163.367
R868 B.n704 B.n61 163.367
R869 B.n62 B.n61 163.367
R870 B.n63 B.n62 163.367
R871 B.n709 B.n63 163.367
R872 B.n709 B.n68 163.367
R873 B.n69 B.n68 163.367
R874 B.n70 B.n69 163.367
R875 B.n714 B.n70 163.367
R876 B.n714 B.n75 163.367
R877 B.n76 B.n75 163.367
R878 B.n77 B.n76 163.367
R879 B.n719 B.n77 163.367
R880 B.n719 B.n82 163.367
R881 B.n83 B.n82 163.367
R882 B.n84 B.n83 163.367
R883 B.n724 B.n84 163.367
R884 B.n724 B.n89 163.367
R885 B.n90 B.n89 163.367
R886 B.n91 B.n90 163.367
R887 B.n729 B.n91 163.367
R888 B.n729 B.n96 163.367
R889 B.n97 B.n96 163.367
R890 B.n98 B.n97 163.367
R891 B.n734 B.n98 163.367
R892 B.n734 B.n103 163.367
R893 B.n104 B.n103 163.367
R894 B.n142 B.n141 163.367
R895 B.n146 B.n145 163.367
R896 B.n150 B.n149 163.367
R897 B.n154 B.n153 163.367
R898 B.n158 B.n157 163.367
R899 B.n162 B.n161 163.367
R900 B.n166 B.n165 163.367
R901 B.n170 B.n169 163.367
R902 B.n174 B.n173 163.367
R903 B.n178 B.n177 163.367
R904 B.n182 B.n181 163.367
R905 B.n186 B.n185 163.367
R906 B.n190 B.n189 163.367
R907 B.n194 B.n193 163.367
R908 B.n198 B.n197 163.367
R909 B.n202 B.n201 163.367
R910 B.n206 B.n205 163.367
R911 B.n210 B.n209 163.367
R912 B.n214 B.n213 163.367
R913 B.n218 B.n217 163.367
R914 B.n222 B.n221 163.367
R915 B.n226 B.n225 163.367
R916 B.n230 B.n229 163.367
R917 B.n234 B.n233 163.367
R918 B.n238 B.n237 163.367
R919 B.n240 B.n131 163.367
R920 B.n491 B.n351 114.594
R921 B.n742 B.n741 114.594
R922 B.n490 B.n489 71.676
R923 B.n484 B.n355 71.676
R924 B.n481 B.n356 71.676
R925 B.n477 B.n357 71.676
R926 B.n473 B.n358 71.676
R927 B.n469 B.n359 71.676
R928 B.n465 B.n360 71.676
R929 B.n461 B.n361 71.676
R930 B.n457 B.n362 71.676
R931 B.n453 B.n363 71.676
R932 B.n449 B.n364 71.676
R933 B.n444 B.n365 71.676
R934 B.n440 B.n366 71.676
R935 B.n436 B.n367 71.676
R936 B.n432 B.n368 71.676
R937 B.n428 B.n369 71.676
R938 B.n423 B.n370 71.676
R939 B.n419 B.n371 71.676
R940 B.n415 B.n372 71.676
R941 B.n411 B.n373 71.676
R942 B.n407 B.n374 71.676
R943 B.n403 B.n375 71.676
R944 B.n399 B.n376 71.676
R945 B.n395 B.n377 71.676
R946 B.n391 B.n378 71.676
R947 B.n387 B.n379 71.676
R948 B.n138 B.n105 71.676
R949 B.n142 B.n106 71.676
R950 B.n146 B.n107 71.676
R951 B.n150 B.n108 71.676
R952 B.n154 B.n109 71.676
R953 B.n158 B.n110 71.676
R954 B.n162 B.n111 71.676
R955 B.n166 B.n112 71.676
R956 B.n170 B.n113 71.676
R957 B.n174 B.n114 71.676
R958 B.n178 B.n115 71.676
R959 B.n182 B.n116 71.676
R960 B.n186 B.n117 71.676
R961 B.n190 B.n118 71.676
R962 B.n194 B.n119 71.676
R963 B.n198 B.n120 71.676
R964 B.n202 B.n121 71.676
R965 B.n206 B.n122 71.676
R966 B.n210 B.n123 71.676
R967 B.n214 B.n124 71.676
R968 B.n218 B.n125 71.676
R969 B.n222 B.n126 71.676
R970 B.n226 B.n127 71.676
R971 B.n230 B.n128 71.676
R972 B.n234 B.n129 71.676
R973 B.n238 B.n130 71.676
R974 B.n740 B.n131 71.676
R975 B.n740 B.n739 71.676
R976 B.n240 B.n130 71.676
R977 B.n237 B.n129 71.676
R978 B.n233 B.n128 71.676
R979 B.n229 B.n127 71.676
R980 B.n225 B.n126 71.676
R981 B.n221 B.n125 71.676
R982 B.n217 B.n124 71.676
R983 B.n213 B.n123 71.676
R984 B.n209 B.n122 71.676
R985 B.n205 B.n121 71.676
R986 B.n201 B.n120 71.676
R987 B.n197 B.n119 71.676
R988 B.n193 B.n118 71.676
R989 B.n189 B.n117 71.676
R990 B.n185 B.n116 71.676
R991 B.n181 B.n115 71.676
R992 B.n177 B.n114 71.676
R993 B.n173 B.n113 71.676
R994 B.n169 B.n112 71.676
R995 B.n165 B.n111 71.676
R996 B.n161 B.n110 71.676
R997 B.n157 B.n109 71.676
R998 B.n153 B.n108 71.676
R999 B.n149 B.n107 71.676
R1000 B.n145 B.n106 71.676
R1001 B.n141 B.n105 71.676
R1002 B.n490 B.n381 71.676
R1003 B.n482 B.n355 71.676
R1004 B.n478 B.n356 71.676
R1005 B.n474 B.n357 71.676
R1006 B.n470 B.n358 71.676
R1007 B.n466 B.n359 71.676
R1008 B.n462 B.n360 71.676
R1009 B.n458 B.n361 71.676
R1010 B.n454 B.n362 71.676
R1011 B.n450 B.n363 71.676
R1012 B.n445 B.n364 71.676
R1013 B.n441 B.n365 71.676
R1014 B.n437 B.n366 71.676
R1015 B.n433 B.n367 71.676
R1016 B.n429 B.n368 71.676
R1017 B.n424 B.n369 71.676
R1018 B.n420 B.n370 71.676
R1019 B.n416 B.n371 71.676
R1020 B.n412 B.n372 71.676
R1021 B.n408 B.n373 71.676
R1022 B.n404 B.n374 71.676
R1023 B.n400 B.n375 71.676
R1024 B.n396 B.n376 71.676
R1025 B.n392 B.n377 71.676
R1026 B.n388 B.n378 71.676
R1027 B.n379 B.n354 71.676
R1028 B.n497 B.n351 70.2023
R1029 B.n497 B.n347 70.2023
R1030 B.n503 B.n347 70.2023
R1031 B.n503 B.n343 70.2023
R1032 B.n509 B.n343 70.2023
R1033 B.n509 B.n339 70.2023
R1034 B.n515 B.n339 70.2023
R1035 B.n521 B.n335 70.2023
R1036 B.n521 B.n331 70.2023
R1037 B.n527 B.n331 70.2023
R1038 B.n527 B.n327 70.2023
R1039 B.n533 B.n327 70.2023
R1040 B.n533 B.n323 70.2023
R1041 B.n539 B.n323 70.2023
R1042 B.n539 B.n319 70.2023
R1043 B.n546 B.n319 70.2023
R1044 B.n546 B.n545 70.2023
R1045 B.n552 B.n312 70.2023
R1046 B.n558 B.n312 70.2023
R1047 B.n558 B.n308 70.2023
R1048 B.n564 B.n308 70.2023
R1049 B.n564 B.n304 70.2023
R1050 B.n571 B.n304 70.2023
R1051 B.n571 B.n570 70.2023
R1052 B.n577 B.n297 70.2023
R1053 B.n583 B.n297 70.2023
R1054 B.n583 B.n293 70.2023
R1055 B.n589 B.n293 70.2023
R1056 B.n589 B.n289 70.2023
R1057 B.n595 B.n289 70.2023
R1058 B.n595 B.n285 70.2023
R1059 B.n601 B.n285 70.2023
R1060 B.n607 B.n281 70.2023
R1061 B.n607 B.n277 70.2023
R1062 B.n613 B.n277 70.2023
R1063 B.n613 B.n273 70.2023
R1064 B.n619 B.n273 70.2023
R1065 B.n619 B.n269 70.2023
R1066 B.n625 B.n269 70.2023
R1067 B.n631 B.n265 70.2023
R1068 B.n631 B.n261 70.2023
R1069 B.n637 B.n261 70.2023
R1070 B.n637 B.n257 70.2023
R1071 B.n643 B.n257 70.2023
R1072 B.n643 B.n253 70.2023
R1073 B.n649 B.n253 70.2023
R1074 B.n656 B.n249 70.2023
R1075 B.n656 B.n245 70.2023
R1076 B.n662 B.n245 70.2023
R1077 B.n662 B.n4 70.2023
R1078 B.n855 B.n4 70.2023
R1079 B.n855 B.n854 70.2023
R1080 B.n854 B.n853 70.2023
R1081 B.n853 B.n8 70.2023
R1082 B.n847 B.n8 70.2023
R1083 B.n847 B.n846 70.2023
R1084 B.n845 B.n15 70.2023
R1085 B.n839 B.n15 70.2023
R1086 B.n839 B.n838 70.2023
R1087 B.n838 B.n837 70.2023
R1088 B.n837 B.n22 70.2023
R1089 B.n831 B.n22 70.2023
R1090 B.n831 B.n830 70.2023
R1091 B.n829 B.n29 70.2023
R1092 B.n823 B.n29 70.2023
R1093 B.n823 B.n822 70.2023
R1094 B.n822 B.n821 70.2023
R1095 B.n821 B.n36 70.2023
R1096 B.n815 B.n36 70.2023
R1097 B.n815 B.n814 70.2023
R1098 B.n813 B.n43 70.2023
R1099 B.n807 B.n43 70.2023
R1100 B.n807 B.n806 70.2023
R1101 B.n806 B.n805 70.2023
R1102 B.n805 B.n50 70.2023
R1103 B.n799 B.n50 70.2023
R1104 B.n799 B.n798 70.2023
R1105 B.n798 B.n797 70.2023
R1106 B.n791 B.n60 70.2023
R1107 B.n791 B.n790 70.2023
R1108 B.n790 B.n789 70.2023
R1109 B.n789 B.n64 70.2023
R1110 B.n783 B.n64 70.2023
R1111 B.n783 B.n782 70.2023
R1112 B.n782 B.n781 70.2023
R1113 B.n775 B.n74 70.2023
R1114 B.n775 B.n774 70.2023
R1115 B.n774 B.n773 70.2023
R1116 B.n773 B.n78 70.2023
R1117 B.n767 B.n78 70.2023
R1118 B.n767 B.n766 70.2023
R1119 B.n766 B.n765 70.2023
R1120 B.n765 B.n85 70.2023
R1121 B.n759 B.n85 70.2023
R1122 B.n759 B.n758 70.2023
R1123 B.n757 B.n92 70.2023
R1124 B.n751 B.n92 70.2023
R1125 B.n751 B.n750 70.2023
R1126 B.n750 B.n749 70.2023
R1127 B.n749 B.n99 70.2023
R1128 B.n743 B.n99 70.2023
R1129 B.n743 B.n742 70.2023
R1130 B.n570 B.t4 69.1699
R1131 B.n60 B.t1 69.1699
R1132 B.t3 B.n281 62.9756
R1133 B.n814 B.t0 62.9756
R1134 B.n545 B.t7 60.9109
R1135 B.n74 B.t9 60.9109
R1136 B.n426 B.n385 59.5399
R1137 B.n447 B.n383 59.5399
R1138 B.n137 B.n136 59.5399
R1139 B.n134 B.n133 59.5399
R1140 B.t8 B.n265 54.7166
R1141 B.n830 B.t5 54.7166
R1142 B.n385 B.n384 53.5278
R1143 B.n383 B.n382 53.5278
R1144 B.n136 B.n135 53.5278
R1145 B.n133 B.n132 53.5278
R1146 B.t2 B.n249 46.4576
R1147 B.n846 B.t6 46.4576
R1148 B.n515 B.t15 38.1985
R1149 B.t11 B.n757 38.1985
R1150 B.t15 B.n335 32.0043
R1151 B.n758 B.t11 32.0043
R1152 B.n139 B.n101 29.8151
R1153 B.n494 B.n493 29.8151
R1154 B.n488 B.n349 29.8151
R1155 B.n738 B.n737 29.8151
R1156 B.n649 B.t2 23.7452
R1157 B.t6 B.n845 23.7452
R1158 B B.n857 18.0485
R1159 B.n625 B.t8 15.4862
R1160 B.t5 B.n829 15.4862
R1161 B.n140 B.n139 10.6151
R1162 B.n143 B.n140 10.6151
R1163 B.n144 B.n143 10.6151
R1164 B.n147 B.n144 10.6151
R1165 B.n148 B.n147 10.6151
R1166 B.n151 B.n148 10.6151
R1167 B.n152 B.n151 10.6151
R1168 B.n155 B.n152 10.6151
R1169 B.n156 B.n155 10.6151
R1170 B.n159 B.n156 10.6151
R1171 B.n160 B.n159 10.6151
R1172 B.n163 B.n160 10.6151
R1173 B.n164 B.n163 10.6151
R1174 B.n167 B.n164 10.6151
R1175 B.n168 B.n167 10.6151
R1176 B.n171 B.n168 10.6151
R1177 B.n172 B.n171 10.6151
R1178 B.n175 B.n172 10.6151
R1179 B.n176 B.n175 10.6151
R1180 B.n179 B.n176 10.6151
R1181 B.n180 B.n179 10.6151
R1182 B.n184 B.n183 10.6151
R1183 B.n187 B.n184 10.6151
R1184 B.n188 B.n187 10.6151
R1185 B.n191 B.n188 10.6151
R1186 B.n192 B.n191 10.6151
R1187 B.n195 B.n192 10.6151
R1188 B.n196 B.n195 10.6151
R1189 B.n199 B.n196 10.6151
R1190 B.n200 B.n199 10.6151
R1191 B.n204 B.n203 10.6151
R1192 B.n207 B.n204 10.6151
R1193 B.n208 B.n207 10.6151
R1194 B.n211 B.n208 10.6151
R1195 B.n212 B.n211 10.6151
R1196 B.n215 B.n212 10.6151
R1197 B.n216 B.n215 10.6151
R1198 B.n219 B.n216 10.6151
R1199 B.n220 B.n219 10.6151
R1200 B.n223 B.n220 10.6151
R1201 B.n224 B.n223 10.6151
R1202 B.n227 B.n224 10.6151
R1203 B.n228 B.n227 10.6151
R1204 B.n231 B.n228 10.6151
R1205 B.n232 B.n231 10.6151
R1206 B.n235 B.n232 10.6151
R1207 B.n236 B.n235 10.6151
R1208 B.n239 B.n236 10.6151
R1209 B.n241 B.n239 10.6151
R1210 B.n242 B.n241 10.6151
R1211 B.n738 B.n242 10.6151
R1212 B.n495 B.n494 10.6151
R1213 B.n495 B.n345 10.6151
R1214 B.n505 B.n345 10.6151
R1215 B.n506 B.n505 10.6151
R1216 B.n507 B.n506 10.6151
R1217 B.n507 B.n337 10.6151
R1218 B.n517 B.n337 10.6151
R1219 B.n518 B.n517 10.6151
R1220 B.n519 B.n518 10.6151
R1221 B.n519 B.n329 10.6151
R1222 B.n529 B.n329 10.6151
R1223 B.n530 B.n529 10.6151
R1224 B.n531 B.n530 10.6151
R1225 B.n531 B.n321 10.6151
R1226 B.n541 B.n321 10.6151
R1227 B.n542 B.n541 10.6151
R1228 B.n543 B.n542 10.6151
R1229 B.n543 B.n314 10.6151
R1230 B.n554 B.n314 10.6151
R1231 B.n555 B.n554 10.6151
R1232 B.n556 B.n555 10.6151
R1233 B.n556 B.n306 10.6151
R1234 B.n566 B.n306 10.6151
R1235 B.n567 B.n566 10.6151
R1236 B.n568 B.n567 10.6151
R1237 B.n568 B.n299 10.6151
R1238 B.n579 B.n299 10.6151
R1239 B.n580 B.n579 10.6151
R1240 B.n581 B.n580 10.6151
R1241 B.n581 B.n291 10.6151
R1242 B.n591 B.n291 10.6151
R1243 B.n592 B.n591 10.6151
R1244 B.n593 B.n592 10.6151
R1245 B.n593 B.n283 10.6151
R1246 B.n603 B.n283 10.6151
R1247 B.n604 B.n603 10.6151
R1248 B.n605 B.n604 10.6151
R1249 B.n605 B.n275 10.6151
R1250 B.n615 B.n275 10.6151
R1251 B.n616 B.n615 10.6151
R1252 B.n617 B.n616 10.6151
R1253 B.n617 B.n267 10.6151
R1254 B.n627 B.n267 10.6151
R1255 B.n628 B.n627 10.6151
R1256 B.n629 B.n628 10.6151
R1257 B.n629 B.n259 10.6151
R1258 B.n639 B.n259 10.6151
R1259 B.n640 B.n639 10.6151
R1260 B.n641 B.n640 10.6151
R1261 B.n641 B.n251 10.6151
R1262 B.n651 B.n251 10.6151
R1263 B.n652 B.n651 10.6151
R1264 B.n654 B.n652 10.6151
R1265 B.n654 B.n653 10.6151
R1266 B.n653 B.n243 10.6151
R1267 B.n665 B.n243 10.6151
R1268 B.n666 B.n665 10.6151
R1269 B.n667 B.n666 10.6151
R1270 B.n668 B.n667 10.6151
R1271 B.n670 B.n668 10.6151
R1272 B.n671 B.n670 10.6151
R1273 B.n672 B.n671 10.6151
R1274 B.n673 B.n672 10.6151
R1275 B.n675 B.n673 10.6151
R1276 B.n676 B.n675 10.6151
R1277 B.n677 B.n676 10.6151
R1278 B.n678 B.n677 10.6151
R1279 B.n680 B.n678 10.6151
R1280 B.n681 B.n680 10.6151
R1281 B.n682 B.n681 10.6151
R1282 B.n683 B.n682 10.6151
R1283 B.n685 B.n683 10.6151
R1284 B.n686 B.n685 10.6151
R1285 B.n687 B.n686 10.6151
R1286 B.n688 B.n687 10.6151
R1287 B.n690 B.n688 10.6151
R1288 B.n691 B.n690 10.6151
R1289 B.n692 B.n691 10.6151
R1290 B.n693 B.n692 10.6151
R1291 B.n695 B.n693 10.6151
R1292 B.n696 B.n695 10.6151
R1293 B.n697 B.n696 10.6151
R1294 B.n698 B.n697 10.6151
R1295 B.n700 B.n698 10.6151
R1296 B.n701 B.n700 10.6151
R1297 B.n702 B.n701 10.6151
R1298 B.n703 B.n702 10.6151
R1299 B.n705 B.n703 10.6151
R1300 B.n706 B.n705 10.6151
R1301 B.n707 B.n706 10.6151
R1302 B.n708 B.n707 10.6151
R1303 B.n710 B.n708 10.6151
R1304 B.n711 B.n710 10.6151
R1305 B.n712 B.n711 10.6151
R1306 B.n713 B.n712 10.6151
R1307 B.n715 B.n713 10.6151
R1308 B.n716 B.n715 10.6151
R1309 B.n717 B.n716 10.6151
R1310 B.n718 B.n717 10.6151
R1311 B.n720 B.n718 10.6151
R1312 B.n721 B.n720 10.6151
R1313 B.n722 B.n721 10.6151
R1314 B.n723 B.n722 10.6151
R1315 B.n725 B.n723 10.6151
R1316 B.n726 B.n725 10.6151
R1317 B.n727 B.n726 10.6151
R1318 B.n728 B.n727 10.6151
R1319 B.n730 B.n728 10.6151
R1320 B.n731 B.n730 10.6151
R1321 B.n732 B.n731 10.6151
R1322 B.n733 B.n732 10.6151
R1323 B.n735 B.n733 10.6151
R1324 B.n736 B.n735 10.6151
R1325 B.n737 B.n736 10.6151
R1326 B.n488 B.n487 10.6151
R1327 B.n487 B.n486 10.6151
R1328 B.n486 B.n485 10.6151
R1329 B.n485 B.n483 10.6151
R1330 B.n483 B.n480 10.6151
R1331 B.n480 B.n479 10.6151
R1332 B.n479 B.n476 10.6151
R1333 B.n476 B.n475 10.6151
R1334 B.n475 B.n472 10.6151
R1335 B.n472 B.n471 10.6151
R1336 B.n471 B.n468 10.6151
R1337 B.n468 B.n467 10.6151
R1338 B.n467 B.n464 10.6151
R1339 B.n464 B.n463 10.6151
R1340 B.n463 B.n460 10.6151
R1341 B.n460 B.n459 10.6151
R1342 B.n459 B.n456 10.6151
R1343 B.n456 B.n455 10.6151
R1344 B.n455 B.n452 10.6151
R1345 B.n452 B.n451 10.6151
R1346 B.n451 B.n448 10.6151
R1347 B.n446 B.n443 10.6151
R1348 B.n443 B.n442 10.6151
R1349 B.n442 B.n439 10.6151
R1350 B.n439 B.n438 10.6151
R1351 B.n438 B.n435 10.6151
R1352 B.n435 B.n434 10.6151
R1353 B.n434 B.n431 10.6151
R1354 B.n431 B.n430 10.6151
R1355 B.n430 B.n427 10.6151
R1356 B.n425 B.n422 10.6151
R1357 B.n422 B.n421 10.6151
R1358 B.n421 B.n418 10.6151
R1359 B.n418 B.n417 10.6151
R1360 B.n417 B.n414 10.6151
R1361 B.n414 B.n413 10.6151
R1362 B.n413 B.n410 10.6151
R1363 B.n410 B.n409 10.6151
R1364 B.n409 B.n406 10.6151
R1365 B.n406 B.n405 10.6151
R1366 B.n405 B.n402 10.6151
R1367 B.n402 B.n401 10.6151
R1368 B.n401 B.n398 10.6151
R1369 B.n398 B.n397 10.6151
R1370 B.n397 B.n394 10.6151
R1371 B.n394 B.n393 10.6151
R1372 B.n393 B.n390 10.6151
R1373 B.n390 B.n389 10.6151
R1374 B.n389 B.n386 10.6151
R1375 B.n386 B.n353 10.6151
R1376 B.n493 B.n353 10.6151
R1377 B.n499 B.n349 10.6151
R1378 B.n500 B.n499 10.6151
R1379 B.n501 B.n500 10.6151
R1380 B.n501 B.n341 10.6151
R1381 B.n511 B.n341 10.6151
R1382 B.n512 B.n511 10.6151
R1383 B.n513 B.n512 10.6151
R1384 B.n513 B.n333 10.6151
R1385 B.n523 B.n333 10.6151
R1386 B.n524 B.n523 10.6151
R1387 B.n525 B.n524 10.6151
R1388 B.n525 B.n325 10.6151
R1389 B.n535 B.n325 10.6151
R1390 B.n536 B.n535 10.6151
R1391 B.n537 B.n536 10.6151
R1392 B.n537 B.n317 10.6151
R1393 B.n548 B.n317 10.6151
R1394 B.n549 B.n548 10.6151
R1395 B.n550 B.n549 10.6151
R1396 B.n550 B.n310 10.6151
R1397 B.n560 B.n310 10.6151
R1398 B.n561 B.n560 10.6151
R1399 B.n562 B.n561 10.6151
R1400 B.n562 B.n302 10.6151
R1401 B.n573 B.n302 10.6151
R1402 B.n574 B.n573 10.6151
R1403 B.n575 B.n574 10.6151
R1404 B.n575 B.n295 10.6151
R1405 B.n585 B.n295 10.6151
R1406 B.n586 B.n585 10.6151
R1407 B.n587 B.n586 10.6151
R1408 B.n587 B.n287 10.6151
R1409 B.n597 B.n287 10.6151
R1410 B.n598 B.n597 10.6151
R1411 B.n599 B.n598 10.6151
R1412 B.n599 B.n279 10.6151
R1413 B.n609 B.n279 10.6151
R1414 B.n610 B.n609 10.6151
R1415 B.n611 B.n610 10.6151
R1416 B.n611 B.n271 10.6151
R1417 B.n621 B.n271 10.6151
R1418 B.n622 B.n621 10.6151
R1419 B.n623 B.n622 10.6151
R1420 B.n623 B.n263 10.6151
R1421 B.n633 B.n263 10.6151
R1422 B.n634 B.n633 10.6151
R1423 B.n635 B.n634 10.6151
R1424 B.n635 B.n255 10.6151
R1425 B.n645 B.n255 10.6151
R1426 B.n646 B.n645 10.6151
R1427 B.n647 B.n646 10.6151
R1428 B.n647 B.n247 10.6151
R1429 B.n658 B.n247 10.6151
R1430 B.n659 B.n658 10.6151
R1431 B.n660 B.n659 10.6151
R1432 B.n660 B.n0 10.6151
R1433 B.n851 B.n1 10.6151
R1434 B.n851 B.n850 10.6151
R1435 B.n850 B.n849 10.6151
R1436 B.n849 B.n10 10.6151
R1437 B.n843 B.n10 10.6151
R1438 B.n843 B.n842 10.6151
R1439 B.n842 B.n841 10.6151
R1440 B.n841 B.n17 10.6151
R1441 B.n835 B.n17 10.6151
R1442 B.n835 B.n834 10.6151
R1443 B.n834 B.n833 10.6151
R1444 B.n833 B.n24 10.6151
R1445 B.n827 B.n24 10.6151
R1446 B.n827 B.n826 10.6151
R1447 B.n826 B.n825 10.6151
R1448 B.n825 B.n31 10.6151
R1449 B.n819 B.n31 10.6151
R1450 B.n819 B.n818 10.6151
R1451 B.n818 B.n817 10.6151
R1452 B.n817 B.n38 10.6151
R1453 B.n811 B.n38 10.6151
R1454 B.n811 B.n810 10.6151
R1455 B.n810 B.n809 10.6151
R1456 B.n809 B.n45 10.6151
R1457 B.n803 B.n45 10.6151
R1458 B.n803 B.n802 10.6151
R1459 B.n802 B.n801 10.6151
R1460 B.n801 B.n52 10.6151
R1461 B.n795 B.n52 10.6151
R1462 B.n795 B.n794 10.6151
R1463 B.n794 B.n793 10.6151
R1464 B.n793 B.n58 10.6151
R1465 B.n787 B.n58 10.6151
R1466 B.n787 B.n786 10.6151
R1467 B.n786 B.n785 10.6151
R1468 B.n785 B.n66 10.6151
R1469 B.n779 B.n66 10.6151
R1470 B.n779 B.n778 10.6151
R1471 B.n778 B.n777 10.6151
R1472 B.n777 B.n72 10.6151
R1473 B.n771 B.n72 10.6151
R1474 B.n771 B.n770 10.6151
R1475 B.n770 B.n769 10.6151
R1476 B.n769 B.n80 10.6151
R1477 B.n763 B.n80 10.6151
R1478 B.n763 B.n762 10.6151
R1479 B.n762 B.n761 10.6151
R1480 B.n761 B.n87 10.6151
R1481 B.n755 B.n87 10.6151
R1482 B.n755 B.n754 10.6151
R1483 B.n754 B.n753 10.6151
R1484 B.n753 B.n94 10.6151
R1485 B.n747 B.n94 10.6151
R1486 B.n747 B.n746 10.6151
R1487 B.n746 B.n745 10.6151
R1488 B.n745 B.n101 10.6151
R1489 B.n180 B.n137 9.36635
R1490 B.n203 B.n134 9.36635
R1491 B.n448 B.n447 9.36635
R1492 B.n426 B.n425 9.36635
R1493 B.n552 B.t7 9.29191
R1494 B.n781 B.t9 9.29191
R1495 B.n601 B.t3 7.22715
R1496 B.t0 B.n813 7.22715
R1497 B.n857 B.n0 2.81026
R1498 B.n857 B.n1 2.81026
R1499 B.n183 B.n137 1.24928
R1500 B.n200 B.n134 1.24928
R1501 B.n447 B.n446 1.24928
R1502 B.n427 B.n426 1.24928
R1503 B.n577 B.t4 1.03288
R1504 B.n797 B.t1 1.03288
R1505 VP.n23 VP.n20 161.3
R1506 VP.n25 VP.n24 161.3
R1507 VP.n26 VP.n19 161.3
R1508 VP.n28 VP.n27 161.3
R1509 VP.n29 VP.n18 161.3
R1510 VP.n32 VP.n31 161.3
R1511 VP.n33 VP.n17 161.3
R1512 VP.n35 VP.n34 161.3
R1513 VP.n36 VP.n16 161.3
R1514 VP.n38 VP.n37 161.3
R1515 VP.n39 VP.n15 161.3
R1516 VP.n41 VP.n40 161.3
R1517 VP.n43 VP.n14 161.3
R1518 VP.n45 VP.n44 161.3
R1519 VP.n46 VP.n13 161.3
R1520 VP.n48 VP.n47 161.3
R1521 VP.n49 VP.n12 161.3
R1522 VP.n88 VP.n0 161.3
R1523 VP.n87 VP.n86 161.3
R1524 VP.n85 VP.n1 161.3
R1525 VP.n84 VP.n83 161.3
R1526 VP.n82 VP.n2 161.3
R1527 VP.n80 VP.n79 161.3
R1528 VP.n78 VP.n3 161.3
R1529 VP.n77 VP.n76 161.3
R1530 VP.n75 VP.n4 161.3
R1531 VP.n74 VP.n73 161.3
R1532 VP.n72 VP.n5 161.3
R1533 VP.n71 VP.n70 161.3
R1534 VP.n68 VP.n6 161.3
R1535 VP.n67 VP.n66 161.3
R1536 VP.n65 VP.n7 161.3
R1537 VP.n64 VP.n63 161.3
R1538 VP.n62 VP.n8 161.3
R1539 VP.n60 VP.n59 161.3
R1540 VP.n58 VP.n9 161.3
R1541 VP.n57 VP.n56 161.3
R1542 VP.n55 VP.n10 161.3
R1543 VP.n54 VP.n53 161.3
R1544 VP.n52 VP.n11 97.6287
R1545 VP.n90 VP.n89 97.6287
R1546 VP.n51 VP.n50 97.6287
R1547 VP.n21 VP.t6 85.2357
R1548 VP.n22 VP.n21 72.2118
R1549 VP.n11 VP.t3 53.3577
R1550 VP.n61 VP.t5 53.3577
R1551 VP.n69 VP.t7 53.3577
R1552 VP.n81 VP.t8 53.3577
R1553 VP.n89 VP.t1 53.3577
R1554 VP.n50 VP.t0 53.3577
R1555 VP.n42 VP.t4 53.3577
R1556 VP.n30 VP.t9 53.3577
R1557 VP.n22 VP.t2 53.3577
R1558 VP.n67 VP.n7 53.171
R1559 VP.n76 VP.n75 53.171
R1560 VP.n37 VP.n36 53.171
R1561 VP.n28 VP.n19 53.171
R1562 VP.n56 VP.n9 51.2335
R1563 VP.n83 VP.n1 51.2335
R1564 VP.n44 VP.n13 51.2335
R1565 VP.n52 VP.n51 47.2042
R1566 VP.n56 VP.n55 29.9206
R1567 VP.n87 VP.n1 29.9206
R1568 VP.n48 VP.n13 29.9206
R1569 VP.n68 VP.n67 27.983
R1570 VP.n75 VP.n74 27.983
R1571 VP.n36 VP.n35 27.983
R1572 VP.n29 VP.n28 27.983
R1573 VP.n55 VP.n54 24.5923
R1574 VP.n60 VP.n9 24.5923
R1575 VP.n63 VP.n62 24.5923
R1576 VP.n63 VP.n7 24.5923
R1577 VP.n70 VP.n68 24.5923
R1578 VP.n74 VP.n5 24.5923
R1579 VP.n76 VP.n3 24.5923
R1580 VP.n80 VP.n3 24.5923
R1581 VP.n83 VP.n82 24.5923
R1582 VP.n88 VP.n87 24.5923
R1583 VP.n49 VP.n48 24.5923
R1584 VP.n37 VP.n15 24.5923
R1585 VP.n41 VP.n15 24.5923
R1586 VP.n44 VP.n43 24.5923
R1587 VP.n31 VP.n29 24.5923
R1588 VP.n35 VP.n17 24.5923
R1589 VP.n24 VP.n23 24.5923
R1590 VP.n24 VP.n19 24.5923
R1591 VP.n61 VP.n60 24.1005
R1592 VP.n82 VP.n81 24.1005
R1593 VP.n43 VP.n42 24.1005
R1594 VP.n54 VP.n11 13.2801
R1595 VP.n89 VP.n88 13.2801
R1596 VP.n50 VP.n49 13.2801
R1597 VP.n70 VP.n69 12.2964
R1598 VP.n69 VP.n5 12.2964
R1599 VP.n31 VP.n30 12.2964
R1600 VP.n30 VP.n17 12.2964
R1601 VP.n21 VP.n20 9.68946
R1602 VP.n62 VP.n61 0.492337
R1603 VP.n81 VP.n80 0.492337
R1604 VP.n42 VP.n41 0.492337
R1605 VP.n23 VP.n22 0.492337
R1606 VP.n51 VP.n12 0.278335
R1607 VP.n53 VP.n52 0.278335
R1608 VP.n90 VP.n0 0.278335
R1609 VP.n25 VP.n20 0.189894
R1610 VP.n26 VP.n25 0.189894
R1611 VP.n27 VP.n26 0.189894
R1612 VP.n27 VP.n18 0.189894
R1613 VP.n32 VP.n18 0.189894
R1614 VP.n33 VP.n32 0.189894
R1615 VP.n34 VP.n33 0.189894
R1616 VP.n34 VP.n16 0.189894
R1617 VP.n38 VP.n16 0.189894
R1618 VP.n39 VP.n38 0.189894
R1619 VP.n40 VP.n39 0.189894
R1620 VP.n40 VP.n14 0.189894
R1621 VP.n45 VP.n14 0.189894
R1622 VP.n46 VP.n45 0.189894
R1623 VP.n47 VP.n46 0.189894
R1624 VP.n47 VP.n12 0.189894
R1625 VP.n53 VP.n10 0.189894
R1626 VP.n57 VP.n10 0.189894
R1627 VP.n58 VP.n57 0.189894
R1628 VP.n59 VP.n58 0.189894
R1629 VP.n59 VP.n8 0.189894
R1630 VP.n64 VP.n8 0.189894
R1631 VP.n65 VP.n64 0.189894
R1632 VP.n66 VP.n65 0.189894
R1633 VP.n66 VP.n6 0.189894
R1634 VP.n71 VP.n6 0.189894
R1635 VP.n72 VP.n71 0.189894
R1636 VP.n73 VP.n72 0.189894
R1637 VP.n73 VP.n4 0.189894
R1638 VP.n77 VP.n4 0.189894
R1639 VP.n78 VP.n77 0.189894
R1640 VP.n79 VP.n78 0.189894
R1641 VP.n79 VP.n2 0.189894
R1642 VP.n84 VP.n2 0.189894
R1643 VP.n85 VP.n84 0.189894
R1644 VP.n86 VP.n85 0.189894
R1645 VP.n86 VP.n0 0.189894
R1646 VP VP.n90 0.153485
R1647 VTAIL.n120 VTAIL.n98 289.615
R1648 VTAIL.n24 VTAIL.n2 289.615
R1649 VTAIL.n92 VTAIL.n70 289.615
R1650 VTAIL.n60 VTAIL.n38 289.615
R1651 VTAIL.n106 VTAIL.n105 185
R1652 VTAIL.n111 VTAIL.n110 185
R1653 VTAIL.n113 VTAIL.n112 185
R1654 VTAIL.n102 VTAIL.n101 185
R1655 VTAIL.n119 VTAIL.n118 185
R1656 VTAIL.n121 VTAIL.n120 185
R1657 VTAIL.n10 VTAIL.n9 185
R1658 VTAIL.n15 VTAIL.n14 185
R1659 VTAIL.n17 VTAIL.n16 185
R1660 VTAIL.n6 VTAIL.n5 185
R1661 VTAIL.n23 VTAIL.n22 185
R1662 VTAIL.n25 VTAIL.n24 185
R1663 VTAIL.n93 VTAIL.n92 185
R1664 VTAIL.n91 VTAIL.n90 185
R1665 VTAIL.n74 VTAIL.n73 185
R1666 VTAIL.n85 VTAIL.n84 185
R1667 VTAIL.n83 VTAIL.n82 185
R1668 VTAIL.n78 VTAIL.n77 185
R1669 VTAIL.n61 VTAIL.n60 185
R1670 VTAIL.n59 VTAIL.n58 185
R1671 VTAIL.n42 VTAIL.n41 185
R1672 VTAIL.n53 VTAIL.n52 185
R1673 VTAIL.n51 VTAIL.n50 185
R1674 VTAIL.n46 VTAIL.n45 185
R1675 VTAIL.n107 VTAIL.t6 147.672
R1676 VTAIL.n11 VTAIL.t19 147.672
R1677 VTAIL.n79 VTAIL.t10 147.672
R1678 VTAIL.n47 VTAIL.t2 147.672
R1679 VTAIL.n111 VTAIL.n105 104.615
R1680 VTAIL.n112 VTAIL.n111 104.615
R1681 VTAIL.n112 VTAIL.n101 104.615
R1682 VTAIL.n119 VTAIL.n101 104.615
R1683 VTAIL.n120 VTAIL.n119 104.615
R1684 VTAIL.n15 VTAIL.n9 104.615
R1685 VTAIL.n16 VTAIL.n15 104.615
R1686 VTAIL.n16 VTAIL.n5 104.615
R1687 VTAIL.n23 VTAIL.n5 104.615
R1688 VTAIL.n24 VTAIL.n23 104.615
R1689 VTAIL.n92 VTAIL.n91 104.615
R1690 VTAIL.n91 VTAIL.n73 104.615
R1691 VTAIL.n84 VTAIL.n73 104.615
R1692 VTAIL.n84 VTAIL.n83 104.615
R1693 VTAIL.n83 VTAIL.n77 104.615
R1694 VTAIL.n60 VTAIL.n59 104.615
R1695 VTAIL.n59 VTAIL.n41 104.615
R1696 VTAIL.n52 VTAIL.n41 104.615
R1697 VTAIL.n52 VTAIL.n51 104.615
R1698 VTAIL.n51 VTAIL.n45 104.615
R1699 VTAIL.n69 VTAIL.n68 53.9159
R1700 VTAIL.n67 VTAIL.n66 53.9159
R1701 VTAIL.n37 VTAIL.n36 53.9159
R1702 VTAIL.n35 VTAIL.n34 53.9159
R1703 VTAIL.n127 VTAIL.n126 53.9157
R1704 VTAIL.n1 VTAIL.n0 53.9157
R1705 VTAIL.n31 VTAIL.n30 53.9157
R1706 VTAIL.n33 VTAIL.n32 53.9157
R1707 VTAIL.t6 VTAIL.n105 52.3082
R1708 VTAIL.t19 VTAIL.n9 52.3082
R1709 VTAIL.t10 VTAIL.n77 52.3082
R1710 VTAIL.t2 VTAIL.n45 52.3082
R1711 VTAIL.n125 VTAIL.n124 34.1247
R1712 VTAIL.n29 VTAIL.n28 34.1247
R1713 VTAIL.n97 VTAIL.n96 34.1247
R1714 VTAIL.n65 VTAIL.n64 34.1247
R1715 VTAIL.n35 VTAIL.n33 21.7634
R1716 VTAIL.n125 VTAIL.n97 19.3841
R1717 VTAIL.n107 VTAIL.n106 15.6666
R1718 VTAIL.n11 VTAIL.n10 15.6666
R1719 VTAIL.n79 VTAIL.n78 15.6666
R1720 VTAIL.n47 VTAIL.n46 15.6666
R1721 VTAIL.n110 VTAIL.n109 12.8005
R1722 VTAIL.n14 VTAIL.n13 12.8005
R1723 VTAIL.n82 VTAIL.n81 12.8005
R1724 VTAIL.n50 VTAIL.n49 12.8005
R1725 VTAIL.n113 VTAIL.n104 12.0247
R1726 VTAIL.n17 VTAIL.n8 12.0247
R1727 VTAIL.n85 VTAIL.n76 12.0247
R1728 VTAIL.n53 VTAIL.n44 12.0247
R1729 VTAIL.n114 VTAIL.n102 11.249
R1730 VTAIL.n18 VTAIL.n6 11.249
R1731 VTAIL.n86 VTAIL.n74 11.249
R1732 VTAIL.n54 VTAIL.n42 11.249
R1733 VTAIL.n118 VTAIL.n117 10.4732
R1734 VTAIL.n22 VTAIL.n21 10.4732
R1735 VTAIL.n90 VTAIL.n89 10.4732
R1736 VTAIL.n58 VTAIL.n57 10.4732
R1737 VTAIL.n121 VTAIL.n100 9.69747
R1738 VTAIL.n25 VTAIL.n4 9.69747
R1739 VTAIL.n93 VTAIL.n72 9.69747
R1740 VTAIL.n61 VTAIL.n40 9.69747
R1741 VTAIL.n124 VTAIL.n123 9.45567
R1742 VTAIL.n28 VTAIL.n27 9.45567
R1743 VTAIL.n96 VTAIL.n95 9.45567
R1744 VTAIL.n64 VTAIL.n63 9.45567
R1745 VTAIL.n123 VTAIL.n122 9.3005
R1746 VTAIL.n100 VTAIL.n99 9.3005
R1747 VTAIL.n117 VTAIL.n116 9.3005
R1748 VTAIL.n115 VTAIL.n114 9.3005
R1749 VTAIL.n104 VTAIL.n103 9.3005
R1750 VTAIL.n109 VTAIL.n108 9.3005
R1751 VTAIL.n27 VTAIL.n26 9.3005
R1752 VTAIL.n4 VTAIL.n3 9.3005
R1753 VTAIL.n21 VTAIL.n20 9.3005
R1754 VTAIL.n19 VTAIL.n18 9.3005
R1755 VTAIL.n8 VTAIL.n7 9.3005
R1756 VTAIL.n13 VTAIL.n12 9.3005
R1757 VTAIL.n95 VTAIL.n94 9.3005
R1758 VTAIL.n72 VTAIL.n71 9.3005
R1759 VTAIL.n89 VTAIL.n88 9.3005
R1760 VTAIL.n87 VTAIL.n86 9.3005
R1761 VTAIL.n76 VTAIL.n75 9.3005
R1762 VTAIL.n81 VTAIL.n80 9.3005
R1763 VTAIL.n63 VTAIL.n62 9.3005
R1764 VTAIL.n40 VTAIL.n39 9.3005
R1765 VTAIL.n57 VTAIL.n56 9.3005
R1766 VTAIL.n55 VTAIL.n54 9.3005
R1767 VTAIL.n44 VTAIL.n43 9.3005
R1768 VTAIL.n49 VTAIL.n48 9.3005
R1769 VTAIL.n122 VTAIL.n98 8.92171
R1770 VTAIL.n26 VTAIL.n2 8.92171
R1771 VTAIL.n94 VTAIL.n70 8.92171
R1772 VTAIL.n62 VTAIL.n38 8.92171
R1773 VTAIL.n124 VTAIL.n98 5.04292
R1774 VTAIL.n28 VTAIL.n2 5.04292
R1775 VTAIL.n96 VTAIL.n70 5.04292
R1776 VTAIL.n64 VTAIL.n38 5.04292
R1777 VTAIL.n108 VTAIL.n107 4.38687
R1778 VTAIL.n12 VTAIL.n11 4.38687
R1779 VTAIL.n80 VTAIL.n79 4.38687
R1780 VTAIL.n48 VTAIL.n47 4.38687
R1781 VTAIL.n122 VTAIL.n121 4.26717
R1782 VTAIL.n26 VTAIL.n25 4.26717
R1783 VTAIL.n94 VTAIL.n93 4.26717
R1784 VTAIL.n62 VTAIL.n61 4.26717
R1785 VTAIL.n126 VTAIL.t0 3.6808
R1786 VTAIL.n126 VTAIL.t7 3.6808
R1787 VTAIL.n0 VTAIL.t3 3.6808
R1788 VTAIL.n0 VTAIL.t9 3.6808
R1789 VTAIL.n30 VTAIL.t13 3.6808
R1790 VTAIL.n30 VTAIL.t16 3.6808
R1791 VTAIL.n32 VTAIL.t11 3.6808
R1792 VTAIL.n32 VTAIL.t12 3.6808
R1793 VTAIL.n68 VTAIL.t14 3.6808
R1794 VTAIL.n68 VTAIL.t18 3.6808
R1795 VTAIL.n66 VTAIL.t15 3.6808
R1796 VTAIL.n66 VTAIL.t17 3.6808
R1797 VTAIL.n36 VTAIL.t8 3.6808
R1798 VTAIL.n36 VTAIL.t5 3.6808
R1799 VTAIL.n34 VTAIL.t4 3.6808
R1800 VTAIL.n34 VTAIL.t1 3.6808
R1801 VTAIL.n118 VTAIL.n100 3.49141
R1802 VTAIL.n22 VTAIL.n4 3.49141
R1803 VTAIL.n90 VTAIL.n72 3.49141
R1804 VTAIL.n58 VTAIL.n40 3.49141
R1805 VTAIL.n117 VTAIL.n102 2.71565
R1806 VTAIL.n21 VTAIL.n6 2.71565
R1807 VTAIL.n89 VTAIL.n74 2.71565
R1808 VTAIL.n57 VTAIL.n42 2.71565
R1809 VTAIL.n37 VTAIL.n35 2.37981
R1810 VTAIL.n65 VTAIL.n37 2.37981
R1811 VTAIL.n69 VTAIL.n67 2.37981
R1812 VTAIL.n97 VTAIL.n69 2.37981
R1813 VTAIL.n33 VTAIL.n31 2.37981
R1814 VTAIL.n31 VTAIL.n29 2.37981
R1815 VTAIL.n127 VTAIL.n125 2.37981
R1816 VTAIL.n114 VTAIL.n113 1.93989
R1817 VTAIL.n18 VTAIL.n17 1.93989
R1818 VTAIL.n86 VTAIL.n85 1.93989
R1819 VTAIL.n54 VTAIL.n53 1.93989
R1820 VTAIL VTAIL.n1 1.84317
R1821 VTAIL.n67 VTAIL.n65 1.65998
R1822 VTAIL.n29 VTAIL.n1 1.65998
R1823 VTAIL.n110 VTAIL.n104 1.16414
R1824 VTAIL.n14 VTAIL.n8 1.16414
R1825 VTAIL.n82 VTAIL.n76 1.16414
R1826 VTAIL.n50 VTAIL.n44 1.16414
R1827 VTAIL VTAIL.n127 0.537138
R1828 VTAIL.n109 VTAIL.n106 0.388379
R1829 VTAIL.n13 VTAIL.n10 0.388379
R1830 VTAIL.n81 VTAIL.n78 0.388379
R1831 VTAIL.n49 VTAIL.n46 0.388379
R1832 VTAIL.n108 VTAIL.n103 0.155672
R1833 VTAIL.n115 VTAIL.n103 0.155672
R1834 VTAIL.n116 VTAIL.n115 0.155672
R1835 VTAIL.n116 VTAIL.n99 0.155672
R1836 VTAIL.n123 VTAIL.n99 0.155672
R1837 VTAIL.n12 VTAIL.n7 0.155672
R1838 VTAIL.n19 VTAIL.n7 0.155672
R1839 VTAIL.n20 VTAIL.n19 0.155672
R1840 VTAIL.n20 VTAIL.n3 0.155672
R1841 VTAIL.n27 VTAIL.n3 0.155672
R1842 VTAIL.n95 VTAIL.n71 0.155672
R1843 VTAIL.n88 VTAIL.n71 0.155672
R1844 VTAIL.n88 VTAIL.n87 0.155672
R1845 VTAIL.n87 VTAIL.n75 0.155672
R1846 VTAIL.n80 VTAIL.n75 0.155672
R1847 VTAIL.n63 VTAIL.n39 0.155672
R1848 VTAIL.n56 VTAIL.n39 0.155672
R1849 VTAIL.n56 VTAIL.n55 0.155672
R1850 VTAIL.n55 VTAIL.n43 0.155672
R1851 VTAIL.n48 VTAIL.n43 0.155672
R1852 VDD1.n22 VDD1.n0 289.615
R1853 VDD1.n51 VDD1.n29 289.615
R1854 VDD1.n23 VDD1.n22 185
R1855 VDD1.n21 VDD1.n20 185
R1856 VDD1.n4 VDD1.n3 185
R1857 VDD1.n15 VDD1.n14 185
R1858 VDD1.n13 VDD1.n12 185
R1859 VDD1.n8 VDD1.n7 185
R1860 VDD1.n37 VDD1.n36 185
R1861 VDD1.n42 VDD1.n41 185
R1862 VDD1.n44 VDD1.n43 185
R1863 VDD1.n33 VDD1.n32 185
R1864 VDD1.n50 VDD1.n49 185
R1865 VDD1.n52 VDD1.n51 185
R1866 VDD1.n9 VDD1.t3 147.672
R1867 VDD1.n38 VDD1.t6 147.672
R1868 VDD1.n22 VDD1.n21 104.615
R1869 VDD1.n21 VDD1.n3 104.615
R1870 VDD1.n14 VDD1.n3 104.615
R1871 VDD1.n14 VDD1.n13 104.615
R1872 VDD1.n13 VDD1.n7 104.615
R1873 VDD1.n42 VDD1.n36 104.615
R1874 VDD1.n43 VDD1.n42 104.615
R1875 VDD1.n43 VDD1.n32 104.615
R1876 VDD1.n50 VDD1.n32 104.615
R1877 VDD1.n51 VDD1.n50 104.615
R1878 VDD1.n59 VDD1.n58 72.3236
R1879 VDD1.n28 VDD1.n27 70.5946
R1880 VDD1.n61 VDD1.n60 70.5945
R1881 VDD1.n57 VDD1.n56 70.5945
R1882 VDD1.n28 VDD1.n26 53.1828
R1883 VDD1.n57 VDD1.n55 53.1828
R1884 VDD1.t3 VDD1.n7 52.3082
R1885 VDD1.t6 VDD1.n36 52.3082
R1886 VDD1.n61 VDD1.n59 41.4276
R1887 VDD1.n9 VDD1.n8 15.6666
R1888 VDD1.n38 VDD1.n37 15.6666
R1889 VDD1.n12 VDD1.n11 12.8005
R1890 VDD1.n41 VDD1.n40 12.8005
R1891 VDD1.n15 VDD1.n6 12.0247
R1892 VDD1.n44 VDD1.n35 12.0247
R1893 VDD1.n16 VDD1.n4 11.249
R1894 VDD1.n45 VDD1.n33 11.249
R1895 VDD1.n20 VDD1.n19 10.4732
R1896 VDD1.n49 VDD1.n48 10.4732
R1897 VDD1.n23 VDD1.n2 9.69747
R1898 VDD1.n52 VDD1.n31 9.69747
R1899 VDD1.n26 VDD1.n25 9.45567
R1900 VDD1.n55 VDD1.n54 9.45567
R1901 VDD1.n25 VDD1.n24 9.3005
R1902 VDD1.n2 VDD1.n1 9.3005
R1903 VDD1.n19 VDD1.n18 9.3005
R1904 VDD1.n17 VDD1.n16 9.3005
R1905 VDD1.n6 VDD1.n5 9.3005
R1906 VDD1.n11 VDD1.n10 9.3005
R1907 VDD1.n54 VDD1.n53 9.3005
R1908 VDD1.n31 VDD1.n30 9.3005
R1909 VDD1.n48 VDD1.n47 9.3005
R1910 VDD1.n46 VDD1.n45 9.3005
R1911 VDD1.n35 VDD1.n34 9.3005
R1912 VDD1.n40 VDD1.n39 9.3005
R1913 VDD1.n24 VDD1.n0 8.92171
R1914 VDD1.n53 VDD1.n29 8.92171
R1915 VDD1.n26 VDD1.n0 5.04292
R1916 VDD1.n55 VDD1.n29 5.04292
R1917 VDD1.n10 VDD1.n9 4.38687
R1918 VDD1.n39 VDD1.n38 4.38687
R1919 VDD1.n24 VDD1.n23 4.26717
R1920 VDD1.n53 VDD1.n52 4.26717
R1921 VDD1.n60 VDD1.t5 3.6808
R1922 VDD1.n60 VDD1.t9 3.6808
R1923 VDD1.n27 VDD1.t7 3.6808
R1924 VDD1.n27 VDD1.t0 3.6808
R1925 VDD1.n58 VDD1.t1 3.6808
R1926 VDD1.n58 VDD1.t8 3.6808
R1927 VDD1.n56 VDD1.t4 3.6808
R1928 VDD1.n56 VDD1.t2 3.6808
R1929 VDD1.n20 VDD1.n2 3.49141
R1930 VDD1.n49 VDD1.n31 3.49141
R1931 VDD1.n19 VDD1.n4 2.71565
R1932 VDD1.n48 VDD1.n33 2.71565
R1933 VDD1.n16 VDD1.n15 1.93989
R1934 VDD1.n45 VDD1.n44 1.93989
R1935 VDD1 VDD1.n61 1.72679
R1936 VDD1.n12 VDD1.n6 1.16414
R1937 VDD1.n41 VDD1.n35 1.16414
R1938 VDD1 VDD1.n28 0.653517
R1939 VDD1.n59 VDD1.n57 0.539982
R1940 VDD1.n11 VDD1.n8 0.388379
R1941 VDD1.n40 VDD1.n37 0.388379
R1942 VDD1.n25 VDD1.n1 0.155672
R1943 VDD1.n18 VDD1.n1 0.155672
R1944 VDD1.n18 VDD1.n17 0.155672
R1945 VDD1.n17 VDD1.n5 0.155672
R1946 VDD1.n10 VDD1.n5 0.155672
R1947 VDD1.n39 VDD1.n34 0.155672
R1948 VDD1.n46 VDD1.n34 0.155672
R1949 VDD1.n47 VDD1.n46 0.155672
R1950 VDD1.n47 VDD1.n30 0.155672
R1951 VDD1.n54 VDD1.n30 0.155672
R1952 VN.n77 VN.n40 161.3
R1953 VN.n76 VN.n75 161.3
R1954 VN.n74 VN.n41 161.3
R1955 VN.n73 VN.n72 161.3
R1956 VN.n71 VN.n42 161.3
R1957 VN.n69 VN.n68 161.3
R1958 VN.n67 VN.n43 161.3
R1959 VN.n66 VN.n65 161.3
R1960 VN.n64 VN.n44 161.3
R1961 VN.n63 VN.n62 161.3
R1962 VN.n61 VN.n45 161.3
R1963 VN.n60 VN.n59 161.3
R1964 VN.n58 VN.n46 161.3
R1965 VN.n57 VN.n56 161.3
R1966 VN.n55 VN.n48 161.3
R1967 VN.n54 VN.n53 161.3
R1968 VN.n52 VN.n49 161.3
R1969 VN.n37 VN.n0 161.3
R1970 VN.n36 VN.n35 161.3
R1971 VN.n34 VN.n1 161.3
R1972 VN.n33 VN.n32 161.3
R1973 VN.n31 VN.n2 161.3
R1974 VN.n29 VN.n28 161.3
R1975 VN.n27 VN.n3 161.3
R1976 VN.n26 VN.n25 161.3
R1977 VN.n24 VN.n4 161.3
R1978 VN.n23 VN.n22 161.3
R1979 VN.n21 VN.n5 161.3
R1980 VN.n20 VN.n19 161.3
R1981 VN.n17 VN.n6 161.3
R1982 VN.n16 VN.n15 161.3
R1983 VN.n14 VN.n7 161.3
R1984 VN.n13 VN.n12 161.3
R1985 VN.n11 VN.n8 161.3
R1986 VN.n39 VN.n38 97.6287
R1987 VN.n79 VN.n78 97.6287
R1988 VN.n9 VN.t5 85.2357
R1989 VN.n50 VN.t6 85.2357
R1990 VN.n10 VN.n9 72.2118
R1991 VN.n51 VN.n50 72.2118
R1992 VN.n10 VN.t4 53.3577
R1993 VN.n18 VN.t1 53.3577
R1994 VN.n30 VN.t8 53.3577
R1995 VN.n38 VN.t9 53.3577
R1996 VN.n51 VN.t2 53.3577
R1997 VN.n47 VN.t0 53.3577
R1998 VN.n70 VN.t7 53.3577
R1999 VN.n78 VN.t3 53.3577
R2000 VN.n16 VN.n7 53.171
R2001 VN.n25 VN.n24 53.171
R2002 VN.n57 VN.n48 53.171
R2003 VN.n65 VN.n64 53.171
R2004 VN.n32 VN.n1 51.2335
R2005 VN.n72 VN.n41 51.2335
R2006 VN VN.n79 47.483
R2007 VN.n36 VN.n1 29.9206
R2008 VN.n76 VN.n41 29.9206
R2009 VN.n17 VN.n16 27.983
R2010 VN.n24 VN.n23 27.983
R2011 VN.n58 VN.n57 27.983
R2012 VN.n64 VN.n63 27.983
R2013 VN.n12 VN.n11 24.5923
R2014 VN.n12 VN.n7 24.5923
R2015 VN.n19 VN.n17 24.5923
R2016 VN.n23 VN.n5 24.5923
R2017 VN.n25 VN.n3 24.5923
R2018 VN.n29 VN.n3 24.5923
R2019 VN.n32 VN.n31 24.5923
R2020 VN.n37 VN.n36 24.5923
R2021 VN.n53 VN.n48 24.5923
R2022 VN.n53 VN.n52 24.5923
R2023 VN.n63 VN.n45 24.5923
R2024 VN.n59 VN.n58 24.5923
R2025 VN.n72 VN.n71 24.5923
R2026 VN.n69 VN.n43 24.5923
R2027 VN.n65 VN.n43 24.5923
R2028 VN.n77 VN.n76 24.5923
R2029 VN.n31 VN.n30 24.1005
R2030 VN.n71 VN.n70 24.1005
R2031 VN.n38 VN.n37 13.2801
R2032 VN.n78 VN.n77 13.2801
R2033 VN.n19 VN.n18 12.2964
R2034 VN.n18 VN.n5 12.2964
R2035 VN.n47 VN.n45 12.2964
R2036 VN.n59 VN.n47 12.2964
R2037 VN.n50 VN.n49 9.68946
R2038 VN.n9 VN.n8 9.68946
R2039 VN.n11 VN.n10 0.492337
R2040 VN.n30 VN.n29 0.492337
R2041 VN.n52 VN.n51 0.492337
R2042 VN.n70 VN.n69 0.492337
R2043 VN.n79 VN.n40 0.278335
R2044 VN.n39 VN.n0 0.278335
R2045 VN.n75 VN.n40 0.189894
R2046 VN.n75 VN.n74 0.189894
R2047 VN.n74 VN.n73 0.189894
R2048 VN.n73 VN.n42 0.189894
R2049 VN.n68 VN.n42 0.189894
R2050 VN.n68 VN.n67 0.189894
R2051 VN.n67 VN.n66 0.189894
R2052 VN.n66 VN.n44 0.189894
R2053 VN.n62 VN.n44 0.189894
R2054 VN.n62 VN.n61 0.189894
R2055 VN.n61 VN.n60 0.189894
R2056 VN.n60 VN.n46 0.189894
R2057 VN.n56 VN.n46 0.189894
R2058 VN.n56 VN.n55 0.189894
R2059 VN.n55 VN.n54 0.189894
R2060 VN.n54 VN.n49 0.189894
R2061 VN.n13 VN.n8 0.189894
R2062 VN.n14 VN.n13 0.189894
R2063 VN.n15 VN.n14 0.189894
R2064 VN.n15 VN.n6 0.189894
R2065 VN.n20 VN.n6 0.189894
R2066 VN.n21 VN.n20 0.189894
R2067 VN.n22 VN.n21 0.189894
R2068 VN.n22 VN.n4 0.189894
R2069 VN.n26 VN.n4 0.189894
R2070 VN.n27 VN.n26 0.189894
R2071 VN.n28 VN.n27 0.189894
R2072 VN.n28 VN.n2 0.189894
R2073 VN.n33 VN.n2 0.189894
R2074 VN.n34 VN.n33 0.189894
R2075 VN.n35 VN.n34 0.189894
R2076 VN.n35 VN.n0 0.189894
R2077 VN VN.n39 0.153485
R2078 VDD2.n53 VDD2.n31 289.615
R2079 VDD2.n22 VDD2.n0 289.615
R2080 VDD2.n54 VDD2.n53 185
R2081 VDD2.n52 VDD2.n51 185
R2082 VDD2.n35 VDD2.n34 185
R2083 VDD2.n46 VDD2.n45 185
R2084 VDD2.n44 VDD2.n43 185
R2085 VDD2.n39 VDD2.n38 185
R2086 VDD2.n8 VDD2.n7 185
R2087 VDD2.n13 VDD2.n12 185
R2088 VDD2.n15 VDD2.n14 185
R2089 VDD2.n4 VDD2.n3 185
R2090 VDD2.n21 VDD2.n20 185
R2091 VDD2.n23 VDD2.n22 185
R2092 VDD2.n40 VDD2.t6 147.672
R2093 VDD2.n9 VDD2.t4 147.672
R2094 VDD2.n53 VDD2.n52 104.615
R2095 VDD2.n52 VDD2.n34 104.615
R2096 VDD2.n45 VDD2.n34 104.615
R2097 VDD2.n45 VDD2.n44 104.615
R2098 VDD2.n44 VDD2.n38 104.615
R2099 VDD2.n13 VDD2.n7 104.615
R2100 VDD2.n14 VDD2.n13 104.615
R2101 VDD2.n14 VDD2.n3 104.615
R2102 VDD2.n21 VDD2.n3 104.615
R2103 VDD2.n22 VDD2.n21 104.615
R2104 VDD2.n30 VDD2.n29 72.3236
R2105 VDD2 VDD2.n61 72.3208
R2106 VDD2.n60 VDD2.n59 70.5946
R2107 VDD2.n28 VDD2.n27 70.5945
R2108 VDD2.n28 VDD2.n26 53.1828
R2109 VDD2.t6 VDD2.n38 52.3082
R2110 VDD2.t4 VDD2.n7 52.3082
R2111 VDD2.n58 VDD2.n57 50.8035
R2112 VDD2.n58 VDD2.n30 39.6549
R2113 VDD2.n40 VDD2.n39 15.6666
R2114 VDD2.n9 VDD2.n8 15.6666
R2115 VDD2.n43 VDD2.n42 12.8005
R2116 VDD2.n12 VDD2.n11 12.8005
R2117 VDD2.n46 VDD2.n37 12.0247
R2118 VDD2.n15 VDD2.n6 12.0247
R2119 VDD2.n47 VDD2.n35 11.249
R2120 VDD2.n16 VDD2.n4 11.249
R2121 VDD2.n51 VDD2.n50 10.4732
R2122 VDD2.n20 VDD2.n19 10.4732
R2123 VDD2.n54 VDD2.n33 9.69747
R2124 VDD2.n23 VDD2.n2 9.69747
R2125 VDD2.n57 VDD2.n56 9.45567
R2126 VDD2.n26 VDD2.n25 9.45567
R2127 VDD2.n56 VDD2.n55 9.3005
R2128 VDD2.n33 VDD2.n32 9.3005
R2129 VDD2.n50 VDD2.n49 9.3005
R2130 VDD2.n48 VDD2.n47 9.3005
R2131 VDD2.n37 VDD2.n36 9.3005
R2132 VDD2.n42 VDD2.n41 9.3005
R2133 VDD2.n25 VDD2.n24 9.3005
R2134 VDD2.n2 VDD2.n1 9.3005
R2135 VDD2.n19 VDD2.n18 9.3005
R2136 VDD2.n17 VDD2.n16 9.3005
R2137 VDD2.n6 VDD2.n5 9.3005
R2138 VDD2.n11 VDD2.n10 9.3005
R2139 VDD2.n55 VDD2.n31 8.92171
R2140 VDD2.n24 VDD2.n0 8.92171
R2141 VDD2.n57 VDD2.n31 5.04292
R2142 VDD2.n26 VDD2.n0 5.04292
R2143 VDD2.n41 VDD2.n40 4.38687
R2144 VDD2.n10 VDD2.n9 4.38687
R2145 VDD2.n55 VDD2.n54 4.26717
R2146 VDD2.n24 VDD2.n23 4.26717
R2147 VDD2.n61 VDD2.t7 3.6808
R2148 VDD2.n61 VDD2.t3 3.6808
R2149 VDD2.n59 VDD2.t2 3.6808
R2150 VDD2.n59 VDD2.t9 3.6808
R2151 VDD2.n29 VDD2.t1 3.6808
R2152 VDD2.n29 VDD2.t0 3.6808
R2153 VDD2.n27 VDD2.t5 3.6808
R2154 VDD2.n27 VDD2.t8 3.6808
R2155 VDD2.n51 VDD2.n33 3.49141
R2156 VDD2.n20 VDD2.n2 3.49141
R2157 VDD2.n50 VDD2.n35 2.71565
R2158 VDD2.n19 VDD2.n4 2.71565
R2159 VDD2.n60 VDD2.n58 2.37981
R2160 VDD2.n47 VDD2.n46 1.93989
R2161 VDD2.n16 VDD2.n15 1.93989
R2162 VDD2.n43 VDD2.n37 1.16414
R2163 VDD2.n12 VDD2.n6 1.16414
R2164 VDD2 VDD2.n60 0.653517
R2165 VDD2.n30 VDD2.n28 0.539982
R2166 VDD2.n42 VDD2.n39 0.388379
R2167 VDD2.n11 VDD2.n8 0.388379
R2168 VDD2.n56 VDD2.n32 0.155672
R2169 VDD2.n49 VDD2.n32 0.155672
R2170 VDD2.n49 VDD2.n48 0.155672
R2171 VDD2.n48 VDD2.n36 0.155672
R2172 VDD2.n41 VDD2.n36 0.155672
R2173 VDD2.n10 VDD2.n5 0.155672
R2174 VDD2.n17 VDD2.n5 0.155672
R2175 VDD2.n18 VDD2.n17 0.155672
R2176 VDD2.n18 VDD2.n1 0.155672
R2177 VDD2.n25 VDD2.n1 0.155672
C0 VTAIL VDD1 7.21256f
C1 VDD2 VDD1 2.06282f
C2 VN VTAIL 6.06196f
C3 VDD2 VN 5.00119f
C4 VDD2 VTAIL 7.26381f
C5 VP VDD1 5.40684f
C6 VN VP 6.9147f
C7 VN VDD1 0.153283f
C8 VP VTAIL 6.07616f
C9 VDD2 VP 0.565657f
C10 VDD2 B 5.904286f
C11 VDD1 B 5.823256f
C12 VTAIL B 5.032638f
C13 VN B 16.63641f
C14 VP B 15.18273f
C15 VDD2.n0 B 0.038317f
C16 VDD2.n1 B 0.026497f
C17 VDD2.n2 B 0.014238f
C18 VDD2.n3 B 0.033654f
C19 VDD2.n4 B 0.015076f
C20 VDD2.n5 B 0.026497f
C21 VDD2.n6 B 0.014238f
C22 VDD2.n7 B 0.025241f
C23 VDD2.n8 B 0.019875f
C24 VDD2.t4 B 0.055018f
C25 VDD2.n9 B 0.109703f
C26 VDD2.n10 B 0.554531f
C27 VDD2.n11 B 0.014238f
C28 VDD2.n12 B 0.015076f
C29 VDD2.n13 B 0.033654f
C30 VDD2.n14 B 0.033654f
C31 VDD2.n15 B 0.015076f
C32 VDD2.n16 B 0.014238f
C33 VDD2.n17 B 0.026497f
C34 VDD2.n18 B 0.026497f
C35 VDD2.n19 B 0.014238f
C36 VDD2.n20 B 0.015076f
C37 VDD2.n21 B 0.033654f
C38 VDD2.n22 B 0.074753f
C39 VDD2.n23 B 0.015076f
C40 VDD2.n24 B 0.014238f
C41 VDD2.n25 B 0.064867f
C42 VDD2.n26 B 0.071863f
C43 VDD2.t5 B 0.112651f
C44 VDD2.t8 B 0.112651f
C45 VDD2.n27 B 0.926876f
C46 VDD2.n28 B 0.707557f
C47 VDD2.t1 B 0.112651f
C48 VDD2.t0 B 0.112651f
C49 VDD2.n29 B 0.940605f
C50 VDD2.n30 B 2.55564f
C51 VDD2.n31 B 0.038317f
C52 VDD2.n32 B 0.026497f
C53 VDD2.n33 B 0.014238f
C54 VDD2.n34 B 0.033654f
C55 VDD2.n35 B 0.015076f
C56 VDD2.n36 B 0.026497f
C57 VDD2.n37 B 0.014238f
C58 VDD2.n38 B 0.025241f
C59 VDD2.n39 B 0.019875f
C60 VDD2.t6 B 0.055018f
C61 VDD2.n40 B 0.109703f
C62 VDD2.n41 B 0.554531f
C63 VDD2.n42 B 0.014238f
C64 VDD2.n43 B 0.015076f
C65 VDD2.n44 B 0.033654f
C66 VDD2.n45 B 0.033654f
C67 VDD2.n46 B 0.015076f
C68 VDD2.n47 B 0.014238f
C69 VDD2.n48 B 0.026497f
C70 VDD2.n49 B 0.026497f
C71 VDD2.n50 B 0.014238f
C72 VDD2.n51 B 0.015076f
C73 VDD2.n52 B 0.033654f
C74 VDD2.n53 B 0.074753f
C75 VDD2.n54 B 0.015076f
C76 VDD2.n55 B 0.014238f
C77 VDD2.n56 B 0.064867f
C78 VDD2.n57 B 0.060399f
C79 VDD2.n58 B 2.44653f
C80 VDD2.t2 B 0.112651f
C81 VDD2.t9 B 0.112651f
C82 VDD2.n59 B 0.926881f
C83 VDD2.n60 B 0.471332f
C84 VDD2.t7 B 0.112651f
C85 VDD2.t3 B 0.112651f
C86 VDD2.n61 B 0.940569f
C87 VN.n0 B 0.033378f
C88 VN.t9 B 0.870148f
C89 VN.n1 B 0.024644f
C90 VN.n2 B 0.025319f
C91 VN.t8 B 0.870148f
C92 VN.n3 B 0.046951f
C93 VN.n4 B 0.025319f
C94 VN.n5 B 0.035362f
C95 VN.n6 B 0.025319f
C96 VN.n7 B 0.044709f
C97 VN.n8 B 0.221338f
C98 VN.t4 B 0.870148f
C99 VN.t5 B 1.04823f
C100 VN.n9 B 0.389407f
C101 VN.n10 B 0.392343f
C102 VN.n11 B 0.024236f
C103 VN.n12 B 0.046951f
C104 VN.n13 B 0.025319f
C105 VN.n14 B 0.025319f
C106 VN.n15 B 0.025319f
C107 VN.n16 B 0.026485f
C108 VN.n17 B 0.049367f
C109 VN.t1 B 0.870148f
C110 VN.n18 B 0.332386f
C111 VN.n19 B 0.035362f
C112 VN.n20 B 0.025319f
C113 VN.n21 B 0.025319f
C114 VN.n22 B 0.025319f
C115 VN.n23 B 0.049367f
C116 VN.n24 B 0.026485f
C117 VN.n25 B 0.044709f
C118 VN.n26 B 0.025319f
C119 VN.n27 B 0.025319f
C120 VN.n28 B 0.025319f
C121 VN.n29 B 0.024236f
C122 VN.n30 B 0.332386f
C123 VN.n31 B 0.046488f
C124 VN.n32 B 0.045746f
C125 VN.n33 B 0.025319f
C126 VN.n34 B 0.025319f
C127 VN.n35 B 0.025319f
C128 VN.n36 B 0.050171f
C129 VN.n37 B 0.036289f
C130 VN.n38 B 0.415565f
C131 VN.n39 B 0.037758f
C132 VN.n40 B 0.033378f
C133 VN.t3 B 0.870148f
C134 VN.n41 B 0.024644f
C135 VN.n42 B 0.025319f
C136 VN.t7 B 0.870148f
C137 VN.n43 B 0.046951f
C138 VN.n44 B 0.025319f
C139 VN.n45 B 0.035362f
C140 VN.n46 B 0.025319f
C141 VN.t0 B 0.870148f
C142 VN.n47 B 0.332386f
C143 VN.n48 B 0.044709f
C144 VN.n49 B 0.221338f
C145 VN.t2 B 0.870148f
C146 VN.t6 B 1.04823f
C147 VN.n50 B 0.389407f
C148 VN.n51 B 0.392343f
C149 VN.n52 B 0.024236f
C150 VN.n53 B 0.046951f
C151 VN.n54 B 0.025319f
C152 VN.n55 B 0.025319f
C153 VN.n56 B 0.025319f
C154 VN.n57 B 0.026485f
C155 VN.n58 B 0.049367f
C156 VN.n59 B 0.035362f
C157 VN.n60 B 0.025319f
C158 VN.n61 B 0.025319f
C159 VN.n62 B 0.025319f
C160 VN.n63 B 0.049367f
C161 VN.n64 B 0.026485f
C162 VN.n65 B 0.044709f
C163 VN.n66 B 0.025319f
C164 VN.n67 B 0.025319f
C165 VN.n68 B 0.025319f
C166 VN.n69 B 0.024236f
C167 VN.n70 B 0.332386f
C168 VN.n71 B 0.046488f
C169 VN.n72 B 0.045746f
C170 VN.n73 B 0.025319f
C171 VN.n74 B 0.025319f
C172 VN.n75 B 0.025319f
C173 VN.n76 B 0.050171f
C174 VN.n77 B 0.036289f
C175 VN.n78 B 0.415565f
C176 VN.n79 B 1.3033f
C177 VDD1.n0 B 0.038851f
C178 VDD1.n1 B 0.026867f
C179 VDD1.n2 B 0.014437f
C180 VDD1.n3 B 0.034124f
C181 VDD1.n4 B 0.015286f
C182 VDD1.n5 B 0.026867f
C183 VDD1.n6 B 0.014437f
C184 VDD1.n7 B 0.025593f
C185 VDD1.n8 B 0.020153f
C186 VDD1.t3 B 0.055785f
C187 VDD1.n9 B 0.111233f
C188 VDD1.n10 B 0.562263f
C189 VDD1.n11 B 0.014437f
C190 VDD1.n12 B 0.015286f
C191 VDD1.n13 B 0.034124f
C192 VDD1.n14 B 0.034124f
C193 VDD1.n15 B 0.015286f
C194 VDD1.n16 B 0.014437f
C195 VDD1.n17 B 0.026867f
C196 VDD1.n18 B 0.026867f
C197 VDD1.n19 B 0.014437f
C198 VDD1.n20 B 0.015286f
C199 VDD1.n21 B 0.034124f
C200 VDD1.n22 B 0.075795f
C201 VDD1.n23 B 0.015286f
C202 VDD1.n24 B 0.014437f
C203 VDD1.n25 B 0.065771f
C204 VDD1.n26 B 0.072865f
C205 VDD1.t7 B 0.114222f
C206 VDD1.t0 B 0.114222f
C207 VDD1.n27 B 0.939803f
C208 VDD1.n28 B 0.726092f
C209 VDD1.n29 B 0.038851f
C210 VDD1.n30 B 0.026867f
C211 VDD1.n31 B 0.014437f
C212 VDD1.n32 B 0.034124f
C213 VDD1.n33 B 0.015286f
C214 VDD1.n34 B 0.026867f
C215 VDD1.n35 B 0.014437f
C216 VDD1.n36 B 0.025593f
C217 VDD1.n37 B 0.020153f
C218 VDD1.t6 B 0.055785f
C219 VDD1.n38 B 0.111233f
C220 VDD1.n39 B 0.562263f
C221 VDD1.n40 B 0.014437f
C222 VDD1.n41 B 0.015286f
C223 VDD1.n42 B 0.034124f
C224 VDD1.n43 B 0.034124f
C225 VDD1.n44 B 0.015286f
C226 VDD1.n45 B 0.014437f
C227 VDD1.n46 B 0.026867f
C228 VDD1.n47 B 0.026867f
C229 VDD1.n48 B 0.014437f
C230 VDD1.n49 B 0.015286f
C231 VDD1.n50 B 0.034124f
C232 VDD1.n51 B 0.075795f
C233 VDD1.n52 B 0.015286f
C234 VDD1.n53 B 0.014437f
C235 VDD1.n54 B 0.065771f
C236 VDD1.n55 B 0.072865f
C237 VDD1.t4 B 0.114222f
C238 VDD1.t2 B 0.114222f
C239 VDD1.n56 B 0.939799f
C240 VDD1.n57 B 0.717422f
C241 VDD1.t1 B 0.114222f
C242 VDD1.t8 B 0.114222f
C243 VDD1.n58 B 0.95372f
C244 VDD1.n59 B 2.71507f
C245 VDD1.t5 B 0.114222f
C246 VDD1.t9 B 0.114222f
C247 VDD1.n60 B 0.939799f
C248 VDD1.n61 B 2.77791f
C249 VTAIL.t3 B 0.123622f
C250 VTAIL.t9 B 0.123622f
C251 VTAIL.n0 B 0.946737f
C252 VTAIL.n1 B 0.592142f
C253 VTAIL.n2 B 0.042048f
C254 VTAIL.n3 B 0.029078f
C255 VTAIL.n4 B 0.015625f
C256 VTAIL.n5 B 0.036932f
C257 VTAIL.n6 B 0.016544f
C258 VTAIL.n7 B 0.029078f
C259 VTAIL.n8 B 0.015625f
C260 VTAIL.n9 B 0.027699f
C261 VTAIL.n10 B 0.021811f
C262 VTAIL.t19 B 0.060376f
C263 VTAIL.n11 B 0.120387f
C264 VTAIL.n12 B 0.608536f
C265 VTAIL.n13 B 0.015625f
C266 VTAIL.n14 B 0.016544f
C267 VTAIL.n15 B 0.036932f
C268 VTAIL.n16 B 0.036932f
C269 VTAIL.n17 B 0.016544f
C270 VTAIL.n18 B 0.015625f
C271 VTAIL.n19 B 0.029078f
C272 VTAIL.n20 B 0.029078f
C273 VTAIL.n21 B 0.015625f
C274 VTAIL.n22 B 0.016544f
C275 VTAIL.n23 B 0.036932f
C276 VTAIL.n24 B 0.082033f
C277 VTAIL.n25 B 0.016544f
C278 VTAIL.n26 B 0.015625f
C279 VTAIL.n27 B 0.071184f
C280 VTAIL.n28 B 0.046234f
C281 VTAIL.n29 B 0.405492f
C282 VTAIL.t13 B 0.123622f
C283 VTAIL.t16 B 0.123622f
C284 VTAIL.n30 B 0.946737f
C285 VTAIL.n31 B 0.709866f
C286 VTAIL.t11 B 0.123622f
C287 VTAIL.t12 B 0.123622f
C288 VTAIL.n32 B 0.946737f
C289 VTAIL.n33 B 1.76233f
C290 VTAIL.t4 B 0.123622f
C291 VTAIL.t1 B 0.123622f
C292 VTAIL.n34 B 0.946743f
C293 VTAIL.n35 B 1.76232f
C294 VTAIL.t8 B 0.123622f
C295 VTAIL.t5 B 0.123622f
C296 VTAIL.n36 B 0.946743f
C297 VTAIL.n37 B 0.70986f
C298 VTAIL.n38 B 0.042048f
C299 VTAIL.n39 B 0.029078f
C300 VTAIL.n40 B 0.015625f
C301 VTAIL.n41 B 0.036932f
C302 VTAIL.n42 B 0.016544f
C303 VTAIL.n43 B 0.029078f
C304 VTAIL.n44 B 0.015625f
C305 VTAIL.n45 B 0.027699f
C306 VTAIL.n46 B 0.021811f
C307 VTAIL.t2 B 0.060376f
C308 VTAIL.n47 B 0.120387f
C309 VTAIL.n48 B 0.608536f
C310 VTAIL.n49 B 0.015625f
C311 VTAIL.n50 B 0.016544f
C312 VTAIL.n51 B 0.036932f
C313 VTAIL.n52 B 0.036932f
C314 VTAIL.n53 B 0.016544f
C315 VTAIL.n54 B 0.015625f
C316 VTAIL.n55 B 0.029078f
C317 VTAIL.n56 B 0.029078f
C318 VTAIL.n57 B 0.015625f
C319 VTAIL.n58 B 0.016544f
C320 VTAIL.n59 B 0.036932f
C321 VTAIL.n60 B 0.082033f
C322 VTAIL.n61 B 0.016544f
C323 VTAIL.n62 B 0.015625f
C324 VTAIL.n63 B 0.071184f
C325 VTAIL.n64 B 0.046234f
C326 VTAIL.n65 B 0.405492f
C327 VTAIL.t15 B 0.123622f
C328 VTAIL.t17 B 0.123622f
C329 VTAIL.n66 B 0.946743f
C330 VTAIL.n67 B 0.642416f
C331 VTAIL.t14 B 0.123622f
C332 VTAIL.t18 B 0.123622f
C333 VTAIL.n68 B 0.946743f
C334 VTAIL.n69 B 0.70986f
C335 VTAIL.n70 B 0.042048f
C336 VTAIL.n71 B 0.029078f
C337 VTAIL.n72 B 0.015625f
C338 VTAIL.n73 B 0.036932f
C339 VTAIL.n74 B 0.016544f
C340 VTAIL.n75 B 0.029078f
C341 VTAIL.n76 B 0.015625f
C342 VTAIL.n77 B 0.027699f
C343 VTAIL.n78 B 0.021811f
C344 VTAIL.t10 B 0.060376f
C345 VTAIL.n79 B 0.120387f
C346 VTAIL.n80 B 0.608536f
C347 VTAIL.n81 B 0.015625f
C348 VTAIL.n82 B 0.016544f
C349 VTAIL.n83 B 0.036932f
C350 VTAIL.n84 B 0.036932f
C351 VTAIL.n85 B 0.016544f
C352 VTAIL.n86 B 0.015625f
C353 VTAIL.n87 B 0.029078f
C354 VTAIL.n88 B 0.029078f
C355 VTAIL.n89 B 0.015625f
C356 VTAIL.n90 B 0.016544f
C357 VTAIL.n91 B 0.036932f
C358 VTAIL.n92 B 0.082033f
C359 VTAIL.n93 B 0.016544f
C360 VTAIL.n94 B 0.015625f
C361 VTAIL.n95 B 0.071184f
C362 VTAIL.n96 B 0.046234f
C363 VTAIL.n97 B 1.30247f
C364 VTAIL.n98 B 0.042048f
C365 VTAIL.n99 B 0.029078f
C366 VTAIL.n100 B 0.015625f
C367 VTAIL.n101 B 0.036932f
C368 VTAIL.n102 B 0.016544f
C369 VTAIL.n103 B 0.029078f
C370 VTAIL.n104 B 0.015625f
C371 VTAIL.n105 B 0.027699f
C372 VTAIL.n106 B 0.021811f
C373 VTAIL.t6 B 0.060376f
C374 VTAIL.n107 B 0.120387f
C375 VTAIL.n108 B 0.608536f
C376 VTAIL.n109 B 0.015625f
C377 VTAIL.n110 B 0.016544f
C378 VTAIL.n111 B 0.036932f
C379 VTAIL.n112 B 0.036932f
C380 VTAIL.n113 B 0.016544f
C381 VTAIL.n114 B 0.015625f
C382 VTAIL.n115 B 0.029078f
C383 VTAIL.n116 B 0.029078f
C384 VTAIL.n117 B 0.015625f
C385 VTAIL.n118 B 0.016544f
C386 VTAIL.n119 B 0.036932f
C387 VTAIL.n120 B 0.082033f
C388 VTAIL.n121 B 0.016544f
C389 VTAIL.n122 B 0.015625f
C390 VTAIL.n123 B 0.071184f
C391 VTAIL.n124 B 0.046234f
C392 VTAIL.n125 B 1.30247f
C393 VTAIL.t0 B 0.123622f
C394 VTAIL.t7 B 0.123622f
C395 VTAIL.n126 B 0.946737f
C396 VTAIL.n127 B 0.537217f
C397 VP.n0 B 0.034188f
C398 VP.t1 B 0.891247f
C399 VP.n1 B 0.025241f
C400 VP.n2 B 0.025933f
C401 VP.t8 B 0.891247f
C402 VP.n3 B 0.04809f
C403 VP.n4 B 0.025933f
C404 VP.n5 B 0.036219f
C405 VP.n6 B 0.025933f
C406 VP.n7 B 0.045793f
C407 VP.n8 B 0.025933f
C408 VP.t5 B 0.891247f
C409 VP.n9 B 0.046855f
C410 VP.n10 B 0.025933f
C411 VP.t3 B 0.891247f
C412 VP.n11 B 0.425642f
C413 VP.n12 B 0.034188f
C414 VP.t0 B 0.891247f
C415 VP.n13 B 0.025241f
C416 VP.n14 B 0.025933f
C417 VP.t4 B 0.891247f
C418 VP.n15 B 0.04809f
C419 VP.n16 B 0.025933f
C420 VP.n17 B 0.036219f
C421 VP.n18 B 0.025933f
C422 VP.n19 B 0.045793f
C423 VP.n20 B 0.226705f
C424 VP.t2 B 0.891247f
C425 VP.t6 B 1.07365f
C426 VP.n21 B 0.398849f
C427 VP.n22 B 0.401856f
C428 VP.n23 B 0.024824f
C429 VP.n24 B 0.04809f
C430 VP.n25 B 0.025933f
C431 VP.n26 B 0.025933f
C432 VP.n27 B 0.025933f
C433 VP.n28 B 0.027127f
C434 VP.n29 B 0.050564f
C435 VP.t9 B 0.891247f
C436 VP.n30 B 0.340445f
C437 VP.n31 B 0.036219f
C438 VP.n32 B 0.025933f
C439 VP.n33 B 0.025933f
C440 VP.n34 B 0.025933f
C441 VP.n35 B 0.050564f
C442 VP.n36 B 0.027127f
C443 VP.n37 B 0.045793f
C444 VP.n38 B 0.025933f
C445 VP.n39 B 0.025933f
C446 VP.n40 B 0.025933f
C447 VP.n41 B 0.024824f
C448 VP.n42 B 0.340445f
C449 VP.n43 B 0.047615f
C450 VP.n44 B 0.046855f
C451 VP.n45 B 0.025933f
C452 VP.n46 B 0.025933f
C453 VP.n47 B 0.025933f
C454 VP.n48 B 0.051387f
C455 VP.n49 B 0.037169f
C456 VP.n50 B 0.425642f
C457 VP.n51 B 1.32084f
C458 VP.n52 B 1.34065f
C459 VP.n53 B 0.034188f
C460 VP.n54 B 0.037169f
C461 VP.n55 B 0.051387f
C462 VP.n56 B 0.025241f
C463 VP.n57 B 0.025933f
C464 VP.n58 B 0.025933f
C465 VP.n59 B 0.025933f
C466 VP.n60 B 0.047615f
C467 VP.n61 B 0.340445f
C468 VP.n62 B 0.024824f
C469 VP.n63 B 0.04809f
C470 VP.n64 B 0.025933f
C471 VP.n65 B 0.025933f
C472 VP.n66 B 0.025933f
C473 VP.n67 B 0.027127f
C474 VP.n68 B 0.050564f
C475 VP.t7 B 0.891247f
C476 VP.n69 B 0.340445f
C477 VP.n70 B 0.036219f
C478 VP.n71 B 0.025933f
C479 VP.n72 B 0.025933f
C480 VP.n73 B 0.025933f
C481 VP.n74 B 0.050564f
C482 VP.n75 B 0.027127f
C483 VP.n76 B 0.045793f
C484 VP.n77 B 0.025933f
C485 VP.n78 B 0.025933f
C486 VP.n79 B 0.025933f
C487 VP.n80 B 0.024824f
C488 VP.n81 B 0.340445f
C489 VP.n82 B 0.047615f
C490 VP.n83 B 0.046855f
C491 VP.n84 B 0.025933f
C492 VP.n85 B 0.025933f
C493 VP.n86 B 0.025933f
C494 VP.n87 B 0.051387f
C495 VP.n88 B 0.037169f
C496 VP.n89 B 0.425642f
C497 VP.n90 B 0.038674f
.ends

