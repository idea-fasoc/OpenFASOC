* NGSPICE file created from diff_pair_sample_1005.ext - technology: sky130A

.subckt diff_pair_sample_1005 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5155 pd=13.68 as=0 ps=0 w=6.45 l=1.79
X1 VTAIL.t7 VP.t0 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.5155 pd=13.68 as=1.06425 ps=6.78 w=6.45 l=1.79
X2 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=2.5155 pd=13.68 as=0 ps=0 w=6.45 l=1.79
X3 VDD1.t0 VP.t1 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.06425 pd=6.78 as=2.5155 ps=13.68 w=6.45 l=1.79
X4 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.5155 pd=13.68 as=0 ps=0 w=6.45 l=1.79
X5 VDD2.t3 VN.t0 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.06425 pd=6.78 as=2.5155 ps=13.68 w=6.45 l=1.79
X6 VTAIL.t0 VN.t1 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.5155 pd=13.68 as=1.06425 ps=6.78 w=6.45 l=1.79
X7 VTAIL.t5 VP.t2 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5155 pd=13.68 as=1.06425 ps=6.78 w=6.45 l=1.79
X8 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5155 pd=13.68 as=0 ps=0 w=6.45 l=1.79
X9 VTAIL.t1 VN.t2 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5155 pd=13.68 as=1.06425 ps=6.78 w=6.45 l=1.79
X10 VDD2.t0 VN.t3 VTAIL.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=1.06425 pd=6.78 as=2.5155 ps=13.68 w=6.45 l=1.79
X11 VDD1.t3 VP.t3 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=1.06425 pd=6.78 as=2.5155 ps=13.68 w=6.45 l=1.79
R0 B.n526 B.n525 585
R1 B.n202 B.n82 585
R2 B.n201 B.n200 585
R3 B.n199 B.n198 585
R4 B.n197 B.n196 585
R5 B.n195 B.n194 585
R6 B.n193 B.n192 585
R7 B.n191 B.n190 585
R8 B.n189 B.n188 585
R9 B.n187 B.n186 585
R10 B.n185 B.n184 585
R11 B.n183 B.n182 585
R12 B.n181 B.n180 585
R13 B.n179 B.n178 585
R14 B.n177 B.n176 585
R15 B.n175 B.n174 585
R16 B.n173 B.n172 585
R17 B.n171 B.n170 585
R18 B.n169 B.n168 585
R19 B.n167 B.n166 585
R20 B.n165 B.n164 585
R21 B.n163 B.n162 585
R22 B.n161 B.n160 585
R23 B.n159 B.n158 585
R24 B.n157 B.n156 585
R25 B.n154 B.n153 585
R26 B.n152 B.n151 585
R27 B.n150 B.n149 585
R28 B.n148 B.n147 585
R29 B.n146 B.n145 585
R30 B.n144 B.n143 585
R31 B.n142 B.n141 585
R32 B.n140 B.n139 585
R33 B.n138 B.n137 585
R34 B.n136 B.n135 585
R35 B.n133 B.n132 585
R36 B.n131 B.n130 585
R37 B.n129 B.n128 585
R38 B.n127 B.n126 585
R39 B.n125 B.n124 585
R40 B.n123 B.n122 585
R41 B.n121 B.n120 585
R42 B.n119 B.n118 585
R43 B.n117 B.n116 585
R44 B.n115 B.n114 585
R45 B.n113 B.n112 585
R46 B.n111 B.n110 585
R47 B.n109 B.n108 585
R48 B.n107 B.n106 585
R49 B.n105 B.n104 585
R50 B.n103 B.n102 585
R51 B.n101 B.n100 585
R52 B.n99 B.n98 585
R53 B.n97 B.n96 585
R54 B.n95 B.n94 585
R55 B.n93 B.n92 585
R56 B.n91 B.n90 585
R57 B.n89 B.n88 585
R58 B.n53 B.n52 585
R59 B.n531 B.n530 585
R60 B.n524 B.n83 585
R61 B.n83 B.n50 585
R62 B.n523 B.n49 585
R63 B.n535 B.n49 585
R64 B.n522 B.n48 585
R65 B.n536 B.n48 585
R66 B.n521 B.n47 585
R67 B.n537 B.n47 585
R68 B.n520 B.n519 585
R69 B.n519 B.n43 585
R70 B.n518 B.n42 585
R71 B.n543 B.n42 585
R72 B.n517 B.n41 585
R73 B.n544 B.n41 585
R74 B.n516 B.n40 585
R75 B.n545 B.n40 585
R76 B.n515 B.n514 585
R77 B.n514 B.n36 585
R78 B.n513 B.n35 585
R79 B.n551 B.n35 585
R80 B.n512 B.n34 585
R81 B.n552 B.n34 585
R82 B.n511 B.n33 585
R83 B.n553 B.n33 585
R84 B.n510 B.n509 585
R85 B.n509 B.n29 585
R86 B.n508 B.n28 585
R87 B.n559 B.n28 585
R88 B.n507 B.n27 585
R89 B.n560 B.n27 585
R90 B.n506 B.n26 585
R91 B.n561 B.n26 585
R92 B.n505 B.n504 585
R93 B.n504 B.n25 585
R94 B.n503 B.n21 585
R95 B.n567 B.n21 585
R96 B.n502 B.n20 585
R97 B.n568 B.n20 585
R98 B.n501 B.n19 585
R99 B.n569 B.n19 585
R100 B.n500 B.n499 585
R101 B.n499 B.n15 585
R102 B.n498 B.n14 585
R103 B.n575 B.n14 585
R104 B.n497 B.n13 585
R105 B.n576 B.n13 585
R106 B.n496 B.n12 585
R107 B.n577 B.n12 585
R108 B.n495 B.n494 585
R109 B.n494 B.n8 585
R110 B.n493 B.n7 585
R111 B.n583 B.n7 585
R112 B.n492 B.n6 585
R113 B.n584 B.n6 585
R114 B.n491 B.n5 585
R115 B.n585 B.n5 585
R116 B.n490 B.n489 585
R117 B.n489 B.n4 585
R118 B.n488 B.n203 585
R119 B.n488 B.n487 585
R120 B.n478 B.n204 585
R121 B.n205 B.n204 585
R122 B.n480 B.n479 585
R123 B.n481 B.n480 585
R124 B.n477 B.n209 585
R125 B.n213 B.n209 585
R126 B.n476 B.n475 585
R127 B.n475 B.n474 585
R128 B.n211 B.n210 585
R129 B.n212 B.n211 585
R130 B.n467 B.n466 585
R131 B.n468 B.n467 585
R132 B.n465 B.n218 585
R133 B.n218 B.n217 585
R134 B.n464 B.n463 585
R135 B.n463 B.n462 585
R136 B.n220 B.n219 585
R137 B.n455 B.n220 585
R138 B.n454 B.n453 585
R139 B.n456 B.n454 585
R140 B.n452 B.n225 585
R141 B.n225 B.n224 585
R142 B.n451 B.n450 585
R143 B.n450 B.n449 585
R144 B.n227 B.n226 585
R145 B.n228 B.n227 585
R146 B.n442 B.n441 585
R147 B.n443 B.n442 585
R148 B.n440 B.n233 585
R149 B.n233 B.n232 585
R150 B.n439 B.n438 585
R151 B.n438 B.n437 585
R152 B.n235 B.n234 585
R153 B.n236 B.n235 585
R154 B.n430 B.n429 585
R155 B.n431 B.n430 585
R156 B.n428 B.n240 585
R157 B.n244 B.n240 585
R158 B.n427 B.n426 585
R159 B.n426 B.n425 585
R160 B.n242 B.n241 585
R161 B.n243 B.n242 585
R162 B.n418 B.n417 585
R163 B.n419 B.n418 585
R164 B.n416 B.n249 585
R165 B.n249 B.n248 585
R166 B.n415 B.n414 585
R167 B.n414 B.n413 585
R168 B.n251 B.n250 585
R169 B.n252 B.n251 585
R170 B.n409 B.n408 585
R171 B.n255 B.n254 585
R172 B.n405 B.n404 585
R173 B.n406 B.n405 585
R174 B.n403 B.n285 585
R175 B.n402 B.n401 585
R176 B.n400 B.n399 585
R177 B.n398 B.n397 585
R178 B.n396 B.n395 585
R179 B.n394 B.n393 585
R180 B.n392 B.n391 585
R181 B.n390 B.n389 585
R182 B.n388 B.n387 585
R183 B.n386 B.n385 585
R184 B.n384 B.n383 585
R185 B.n382 B.n381 585
R186 B.n380 B.n379 585
R187 B.n378 B.n377 585
R188 B.n376 B.n375 585
R189 B.n374 B.n373 585
R190 B.n372 B.n371 585
R191 B.n370 B.n369 585
R192 B.n368 B.n367 585
R193 B.n366 B.n365 585
R194 B.n364 B.n363 585
R195 B.n362 B.n361 585
R196 B.n360 B.n359 585
R197 B.n358 B.n357 585
R198 B.n356 B.n355 585
R199 B.n354 B.n353 585
R200 B.n352 B.n351 585
R201 B.n350 B.n349 585
R202 B.n348 B.n347 585
R203 B.n346 B.n345 585
R204 B.n344 B.n343 585
R205 B.n342 B.n341 585
R206 B.n340 B.n339 585
R207 B.n338 B.n337 585
R208 B.n336 B.n335 585
R209 B.n334 B.n333 585
R210 B.n332 B.n331 585
R211 B.n330 B.n329 585
R212 B.n328 B.n327 585
R213 B.n326 B.n325 585
R214 B.n324 B.n323 585
R215 B.n322 B.n321 585
R216 B.n320 B.n319 585
R217 B.n318 B.n317 585
R218 B.n316 B.n315 585
R219 B.n314 B.n313 585
R220 B.n312 B.n311 585
R221 B.n310 B.n309 585
R222 B.n308 B.n307 585
R223 B.n306 B.n305 585
R224 B.n304 B.n303 585
R225 B.n302 B.n301 585
R226 B.n300 B.n299 585
R227 B.n298 B.n297 585
R228 B.n296 B.n295 585
R229 B.n294 B.n293 585
R230 B.n292 B.n284 585
R231 B.n406 B.n284 585
R232 B.n410 B.n253 585
R233 B.n253 B.n252 585
R234 B.n412 B.n411 585
R235 B.n413 B.n412 585
R236 B.n247 B.n246 585
R237 B.n248 B.n247 585
R238 B.n421 B.n420 585
R239 B.n420 B.n419 585
R240 B.n422 B.n245 585
R241 B.n245 B.n243 585
R242 B.n424 B.n423 585
R243 B.n425 B.n424 585
R244 B.n239 B.n238 585
R245 B.n244 B.n239 585
R246 B.n433 B.n432 585
R247 B.n432 B.n431 585
R248 B.n434 B.n237 585
R249 B.n237 B.n236 585
R250 B.n436 B.n435 585
R251 B.n437 B.n436 585
R252 B.n231 B.n230 585
R253 B.n232 B.n231 585
R254 B.n445 B.n444 585
R255 B.n444 B.n443 585
R256 B.n446 B.n229 585
R257 B.n229 B.n228 585
R258 B.n448 B.n447 585
R259 B.n449 B.n448 585
R260 B.n223 B.n222 585
R261 B.n224 B.n223 585
R262 B.n458 B.n457 585
R263 B.n457 B.n456 585
R264 B.n459 B.n221 585
R265 B.n455 B.n221 585
R266 B.n461 B.n460 585
R267 B.n462 B.n461 585
R268 B.n216 B.n215 585
R269 B.n217 B.n216 585
R270 B.n470 B.n469 585
R271 B.n469 B.n468 585
R272 B.n471 B.n214 585
R273 B.n214 B.n212 585
R274 B.n473 B.n472 585
R275 B.n474 B.n473 585
R276 B.n208 B.n207 585
R277 B.n213 B.n208 585
R278 B.n483 B.n482 585
R279 B.n482 B.n481 585
R280 B.n484 B.n206 585
R281 B.n206 B.n205 585
R282 B.n486 B.n485 585
R283 B.n487 B.n486 585
R284 B.n2 B.n0 585
R285 B.n4 B.n2 585
R286 B.n3 B.n1 585
R287 B.n584 B.n3 585
R288 B.n582 B.n581 585
R289 B.n583 B.n582 585
R290 B.n580 B.n9 585
R291 B.n9 B.n8 585
R292 B.n579 B.n578 585
R293 B.n578 B.n577 585
R294 B.n11 B.n10 585
R295 B.n576 B.n11 585
R296 B.n574 B.n573 585
R297 B.n575 B.n574 585
R298 B.n572 B.n16 585
R299 B.n16 B.n15 585
R300 B.n571 B.n570 585
R301 B.n570 B.n569 585
R302 B.n18 B.n17 585
R303 B.n568 B.n18 585
R304 B.n566 B.n565 585
R305 B.n567 B.n566 585
R306 B.n564 B.n22 585
R307 B.n25 B.n22 585
R308 B.n563 B.n562 585
R309 B.n562 B.n561 585
R310 B.n24 B.n23 585
R311 B.n560 B.n24 585
R312 B.n558 B.n557 585
R313 B.n559 B.n558 585
R314 B.n556 B.n30 585
R315 B.n30 B.n29 585
R316 B.n555 B.n554 585
R317 B.n554 B.n553 585
R318 B.n32 B.n31 585
R319 B.n552 B.n32 585
R320 B.n550 B.n549 585
R321 B.n551 B.n550 585
R322 B.n548 B.n37 585
R323 B.n37 B.n36 585
R324 B.n547 B.n546 585
R325 B.n546 B.n545 585
R326 B.n39 B.n38 585
R327 B.n544 B.n39 585
R328 B.n542 B.n541 585
R329 B.n543 B.n542 585
R330 B.n540 B.n44 585
R331 B.n44 B.n43 585
R332 B.n539 B.n538 585
R333 B.n538 B.n537 585
R334 B.n46 B.n45 585
R335 B.n536 B.n46 585
R336 B.n534 B.n533 585
R337 B.n535 B.n534 585
R338 B.n532 B.n51 585
R339 B.n51 B.n50 585
R340 B.n587 B.n586 585
R341 B.n586 B.n585 585
R342 B.n408 B.n253 482.89
R343 B.n530 B.n51 482.89
R344 B.n284 B.n251 482.89
R345 B.n526 B.n83 482.89
R346 B.n289 B.t8 293.219
R347 B.n286 B.t12 293.219
R348 B.n86 B.t15 293.219
R349 B.n84 B.t4 293.219
R350 B.n528 B.n527 256.663
R351 B.n528 B.n81 256.663
R352 B.n528 B.n80 256.663
R353 B.n528 B.n79 256.663
R354 B.n528 B.n78 256.663
R355 B.n528 B.n77 256.663
R356 B.n528 B.n76 256.663
R357 B.n528 B.n75 256.663
R358 B.n528 B.n74 256.663
R359 B.n528 B.n73 256.663
R360 B.n528 B.n72 256.663
R361 B.n528 B.n71 256.663
R362 B.n528 B.n70 256.663
R363 B.n528 B.n69 256.663
R364 B.n528 B.n68 256.663
R365 B.n528 B.n67 256.663
R366 B.n528 B.n66 256.663
R367 B.n528 B.n65 256.663
R368 B.n528 B.n64 256.663
R369 B.n528 B.n63 256.663
R370 B.n528 B.n62 256.663
R371 B.n528 B.n61 256.663
R372 B.n528 B.n60 256.663
R373 B.n528 B.n59 256.663
R374 B.n528 B.n58 256.663
R375 B.n528 B.n57 256.663
R376 B.n528 B.n56 256.663
R377 B.n528 B.n55 256.663
R378 B.n528 B.n54 256.663
R379 B.n529 B.n528 256.663
R380 B.n407 B.n406 256.663
R381 B.n406 B.n256 256.663
R382 B.n406 B.n257 256.663
R383 B.n406 B.n258 256.663
R384 B.n406 B.n259 256.663
R385 B.n406 B.n260 256.663
R386 B.n406 B.n261 256.663
R387 B.n406 B.n262 256.663
R388 B.n406 B.n263 256.663
R389 B.n406 B.n264 256.663
R390 B.n406 B.n265 256.663
R391 B.n406 B.n266 256.663
R392 B.n406 B.n267 256.663
R393 B.n406 B.n268 256.663
R394 B.n406 B.n269 256.663
R395 B.n406 B.n270 256.663
R396 B.n406 B.n271 256.663
R397 B.n406 B.n272 256.663
R398 B.n406 B.n273 256.663
R399 B.n406 B.n274 256.663
R400 B.n406 B.n275 256.663
R401 B.n406 B.n276 256.663
R402 B.n406 B.n277 256.663
R403 B.n406 B.n278 256.663
R404 B.n406 B.n279 256.663
R405 B.n406 B.n280 256.663
R406 B.n406 B.n281 256.663
R407 B.n406 B.n282 256.663
R408 B.n406 B.n283 256.663
R409 B.n412 B.n253 163.367
R410 B.n412 B.n247 163.367
R411 B.n420 B.n247 163.367
R412 B.n420 B.n245 163.367
R413 B.n424 B.n245 163.367
R414 B.n424 B.n239 163.367
R415 B.n432 B.n239 163.367
R416 B.n432 B.n237 163.367
R417 B.n436 B.n237 163.367
R418 B.n436 B.n231 163.367
R419 B.n444 B.n231 163.367
R420 B.n444 B.n229 163.367
R421 B.n448 B.n229 163.367
R422 B.n448 B.n223 163.367
R423 B.n457 B.n223 163.367
R424 B.n457 B.n221 163.367
R425 B.n461 B.n221 163.367
R426 B.n461 B.n216 163.367
R427 B.n469 B.n216 163.367
R428 B.n469 B.n214 163.367
R429 B.n473 B.n214 163.367
R430 B.n473 B.n208 163.367
R431 B.n482 B.n208 163.367
R432 B.n482 B.n206 163.367
R433 B.n486 B.n206 163.367
R434 B.n486 B.n2 163.367
R435 B.n586 B.n2 163.367
R436 B.n586 B.n3 163.367
R437 B.n582 B.n3 163.367
R438 B.n582 B.n9 163.367
R439 B.n578 B.n9 163.367
R440 B.n578 B.n11 163.367
R441 B.n574 B.n11 163.367
R442 B.n574 B.n16 163.367
R443 B.n570 B.n16 163.367
R444 B.n570 B.n18 163.367
R445 B.n566 B.n18 163.367
R446 B.n566 B.n22 163.367
R447 B.n562 B.n22 163.367
R448 B.n562 B.n24 163.367
R449 B.n558 B.n24 163.367
R450 B.n558 B.n30 163.367
R451 B.n554 B.n30 163.367
R452 B.n554 B.n32 163.367
R453 B.n550 B.n32 163.367
R454 B.n550 B.n37 163.367
R455 B.n546 B.n37 163.367
R456 B.n546 B.n39 163.367
R457 B.n542 B.n39 163.367
R458 B.n542 B.n44 163.367
R459 B.n538 B.n44 163.367
R460 B.n538 B.n46 163.367
R461 B.n534 B.n46 163.367
R462 B.n534 B.n51 163.367
R463 B.n405 B.n255 163.367
R464 B.n405 B.n285 163.367
R465 B.n401 B.n400 163.367
R466 B.n397 B.n396 163.367
R467 B.n393 B.n392 163.367
R468 B.n389 B.n388 163.367
R469 B.n385 B.n384 163.367
R470 B.n381 B.n380 163.367
R471 B.n377 B.n376 163.367
R472 B.n373 B.n372 163.367
R473 B.n369 B.n368 163.367
R474 B.n365 B.n364 163.367
R475 B.n361 B.n360 163.367
R476 B.n357 B.n356 163.367
R477 B.n353 B.n352 163.367
R478 B.n349 B.n348 163.367
R479 B.n345 B.n344 163.367
R480 B.n341 B.n340 163.367
R481 B.n337 B.n336 163.367
R482 B.n333 B.n332 163.367
R483 B.n329 B.n328 163.367
R484 B.n325 B.n324 163.367
R485 B.n321 B.n320 163.367
R486 B.n317 B.n316 163.367
R487 B.n313 B.n312 163.367
R488 B.n309 B.n308 163.367
R489 B.n305 B.n304 163.367
R490 B.n301 B.n300 163.367
R491 B.n297 B.n296 163.367
R492 B.n293 B.n284 163.367
R493 B.n414 B.n251 163.367
R494 B.n414 B.n249 163.367
R495 B.n418 B.n249 163.367
R496 B.n418 B.n242 163.367
R497 B.n426 B.n242 163.367
R498 B.n426 B.n240 163.367
R499 B.n430 B.n240 163.367
R500 B.n430 B.n235 163.367
R501 B.n438 B.n235 163.367
R502 B.n438 B.n233 163.367
R503 B.n442 B.n233 163.367
R504 B.n442 B.n227 163.367
R505 B.n450 B.n227 163.367
R506 B.n450 B.n225 163.367
R507 B.n454 B.n225 163.367
R508 B.n454 B.n220 163.367
R509 B.n463 B.n220 163.367
R510 B.n463 B.n218 163.367
R511 B.n467 B.n218 163.367
R512 B.n467 B.n211 163.367
R513 B.n475 B.n211 163.367
R514 B.n475 B.n209 163.367
R515 B.n480 B.n209 163.367
R516 B.n480 B.n204 163.367
R517 B.n488 B.n204 163.367
R518 B.n489 B.n488 163.367
R519 B.n489 B.n5 163.367
R520 B.n6 B.n5 163.367
R521 B.n7 B.n6 163.367
R522 B.n494 B.n7 163.367
R523 B.n494 B.n12 163.367
R524 B.n13 B.n12 163.367
R525 B.n14 B.n13 163.367
R526 B.n499 B.n14 163.367
R527 B.n499 B.n19 163.367
R528 B.n20 B.n19 163.367
R529 B.n21 B.n20 163.367
R530 B.n504 B.n21 163.367
R531 B.n504 B.n26 163.367
R532 B.n27 B.n26 163.367
R533 B.n28 B.n27 163.367
R534 B.n509 B.n28 163.367
R535 B.n509 B.n33 163.367
R536 B.n34 B.n33 163.367
R537 B.n35 B.n34 163.367
R538 B.n514 B.n35 163.367
R539 B.n514 B.n40 163.367
R540 B.n41 B.n40 163.367
R541 B.n42 B.n41 163.367
R542 B.n519 B.n42 163.367
R543 B.n519 B.n47 163.367
R544 B.n48 B.n47 163.367
R545 B.n49 B.n48 163.367
R546 B.n83 B.n49 163.367
R547 B.n88 B.n53 163.367
R548 B.n92 B.n91 163.367
R549 B.n96 B.n95 163.367
R550 B.n100 B.n99 163.367
R551 B.n104 B.n103 163.367
R552 B.n108 B.n107 163.367
R553 B.n112 B.n111 163.367
R554 B.n116 B.n115 163.367
R555 B.n120 B.n119 163.367
R556 B.n124 B.n123 163.367
R557 B.n128 B.n127 163.367
R558 B.n132 B.n131 163.367
R559 B.n137 B.n136 163.367
R560 B.n141 B.n140 163.367
R561 B.n145 B.n144 163.367
R562 B.n149 B.n148 163.367
R563 B.n153 B.n152 163.367
R564 B.n158 B.n157 163.367
R565 B.n162 B.n161 163.367
R566 B.n166 B.n165 163.367
R567 B.n170 B.n169 163.367
R568 B.n174 B.n173 163.367
R569 B.n178 B.n177 163.367
R570 B.n182 B.n181 163.367
R571 B.n186 B.n185 163.367
R572 B.n190 B.n189 163.367
R573 B.n194 B.n193 163.367
R574 B.n198 B.n197 163.367
R575 B.n200 B.n82 163.367
R576 B.n289 B.t11 116.728
R577 B.n84 B.t6 116.728
R578 B.n286 B.t14 116.722
R579 B.n86 B.t16 116.722
R580 B.n406 B.n252 104.136
R581 B.n528 B.n50 104.136
R582 B.n290 B.t10 75.6129
R583 B.n85 B.t7 75.6129
R584 B.n287 B.t13 75.6061
R585 B.n87 B.t17 75.6061
R586 B.n408 B.n407 71.676
R587 B.n285 B.n256 71.676
R588 B.n400 B.n257 71.676
R589 B.n396 B.n258 71.676
R590 B.n392 B.n259 71.676
R591 B.n388 B.n260 71.676
R592 B.n384 B.n261 71.676
R593 B.n380 B.n262 71.676
R594 B.n376 B.n263 71.676
R595 B.n372 B.n264 71.676
R596 B.n368 B.n265 71.676
R597 B.n364 B.n266 71.676
R598 B.n360 B.n267 71.676
R599 B.n356 B.n268 71.676
R600 B.n352 B.n269 71.676
R601 B.n348 B.n270 71.676
R602 B.n344 B.n271 71.676
R603 B.n340 B.n272 71.676
R604 B.n336 B.n273 71.676
R605 B.n332 B.n274 71.676
R606 B.n328 B.n275 71.676
R607 B.n324 B.n276 71.676
R608 B.n320 B.n277 71.676
R609 B.n316 B.n278 71.676
R610 B.n312 B.n279 71.676
R611 B.n308 B.n280 71.676
R612 B.n304 B.n281 71.676
R613 B.n300 B.n282 71.676
R614 B.n296 B.n283 71.676
R615 B.n530 B.n529 71.676
R616 B.n88 B.n54 71.676
R617 B.n92 B.n55 71.676
R618 B.n96 B.n56 71.676
R619 B.n100 B.n57 71.676
R620 B.n104 B.n58 71.676
R621 B.n108 B.n59 71.676
R622 B.n112 B.n60 71.676
R623 B.n116 B.n61 71.676
R624 B.n120 B.n62 71.676
R625 B.n124 B.n63 71.676
R626 B.n128 B.n64 71.676
R627 B.n132 B.n65 71.676
R628 B.n137 B.n66 71.676
R629 B.n141 B.n67 71.676
R630 B.n145 B.n68 71.676
R631 B.n149 B.n69 71.676
R632 B.n153 B.n70 71.676
R633 B.n158 B.n71 71.676
R634 B.n162 B.n72 71.676
R635 B.n166 B.n73 71.676
R636 B.n170 B.n74 71.676
R637 B.n174 B.n75 71.676
R638 B.n178 B.n76 71.676
R639 B.n182 B.n77 71.676
R640 B.n186 B.n78 71.676
R641 B.n190 B.n79 71.676
R642 B.n194 B.n80 71.676
R643 B.n198 B.n81 71.676
R644 B.n527 B.n82 71.676
R645 B.n527 B.n526 71.676
R646 B.n200 B.n81 71.676
R647 B.n197 B.n80 71.676
R648 B.n193 B.n79 71.676
R649 B.n189 B.n78 71.676
R650 B.n185 B.n77 71.676
R651 B.n181 B.n76 71.676
R652 B.n177 B.n75 71.676
R653 B.n173 B.n74 71.676
R654 B.n169 B.n73 71.676
R655 B.n165 B.n72 71.676
R656 B.n161 B.n71 71.676
R657 B.n157 B.n70 71.676
R658 B.n152 B.n69 71.676
R659 B.n148 B.n68 71.676
R660 B.n144 B.n67 71.676
R661 B.n140 B.n66 71.676
R662 B.n136 B.n65 71.676
R663 B.n131 B.n64 71.676
R664 B.n127 B.n63 71.676
R665 B.n123 B.n62 71.676
R666 B.n119 B.n61 71.676
R667 B.n115 B.n60 71.676
R668 B.n111 B.n59 71.676
R669 B.n107 B.n58 71.676
R670 B.n103 B.n57 71.676
R671 B.n99 B.n56 71.676
R672 B.n95 B.n55 71.676
R673 B.n91 B.n54 71.676
R674 B.n529 B.n53 71.676
R675 B.n407 B.n255 71.676
R676 B.n401 B.n256 71.676
R677 B.n397 B.n257 71.676
R678 B.n393 B.n258 71.676
R679 B.n389 B.n259 71.676
R680 B.n385 B.n260 71.676
R681 B.n381 B.n261 71.676
R682 B.n377 B.n262 71.676
R683 B.n373 B.n263 71.676
R684 B.n369 B.n264 71.676
R685 B.n365 B.n265 71.676
R686 B.n361 B.n266 71.676
R687 B.n357 B.n267 71.676
R688 B.n353 B.n268 71.676
R689 B.n349 B.n269 71.676
R690 B.n345 B.n270 71.676
R691 B.n341 B.n271 71.676
R692 B.n337 B.n272 71.676
R693 B.n333 B.n273 71.676
R694 B.n329 B.n274 71.676
R695 B.n325 B.n275 71.676
R696 B.n321 B.n276 71.676
R697 B.n317 B.n277 71.676
R698 B.n313 B.n278 71.676
R699 B.n309 B.n279 71.676
R700 B.n305 B.n280 71.676
R701 B.n301 B.n281 71.676
R702 B.n297 B.n282 71.676
R703 B.n293 B.n283 71.676
R704 B.n413 B.n252 63.7958
R705 B.n413 B.n248 63.7958
R706 B.n419 B.n248 63.7958
R707 B.n419 B.n243 63.7958
R708 B.n425 B.n243 63.7958
R709 B.n425 B.n244 63.7958
R710 B.n431 B.n236 63.7958
R711 B.n437 B.n236 63.7958
R712 B.n437 B.n232 63.7958
R713 B.n443 B.n232 63.7958
R714 B.n443 B.n228 63.7958
R715 B.n449 B.n228 63.7958
R716 B.n449 B.n224 63.7958
R717 B.n456 B.n224 63.7958
R718 B.n456 B.n455 63.7958
R719 B.n462 B.n217 63.7958
R720 B.n468 B.n217 63.7958
R721 B.n468 B.n212 63.7958
R722 B.n474 B.n212 63.7958
R723 B.n474 B.n213 63.7958
R724 B.n481 B.n205 63.7958
R725 B.n487 B.n205 63.7958
R726 B.n487 B.n4 63.7958
R727 B.n585 B.n4 63.7958
R728 B.n585 B.n584 63.7958
R729 B.n584 B.n583 63.7958
R730 B.n583 B.n8 63.7958
R731 B.n577 B.n8 63.7958
R732 B.n576 B.n575 63.7958
R733 B.n575 B.n15 63.7958
R734 B.n569 B.n15 63.7958
R735 B.n569 B.n568 63.7958
R736 B.n568 B.n567 63.7958
R737 B.n561 B.n25 63.7958
R738 B.n561 B.n560 63.7958
R739 B.n560 B.n559 63.7958
R740 B.n559 B.n29 63.7958
R741 B.n553 B.n29 63.7958
R742 B.n553 B.n552 63.7958
R743 B.n552 B.n551 63.7958
R744 B.n551 B.n36 63.7958
R745 B.n545 B.n36 63.7958
R746 B.n544 B.n543 63.7958
R747 B.n543 B.n43 63.7958
R748 B.n537 B.n43 63.7958
R749 B.n537 B.n536 63.7958
R750 B.n536 B.n535 63.7958
R751 B.n535 B.n50 63.7958
R752 B.n462 B.t0 60.9813
R753 B.n567 B.t2 60.9813
R754 B.n291 B.n290 59.5399
R755 B.n288 B.n287 59.5399
R756 B.n134 B.n87 59.5399
R757 B.n155 B.n85 59.5399
R758 B.n481 B.t3 45.9706
R759 B.n577 B.t1 45.9706
R760 B.n290 B.n289 41.1157
R761 B.n287 B.n286 41.1157
R762 B.n87 B.n86 41.1157
R763 B.n85 B.n84 41.1157
R764 B.n244 B.t9 38.4653
R765 B.t5 B.n544 38.4653
R766 B.n532 B.n531 31.3761
R767 B.n525 B.n524 31.3761
R768 B.n292 B.n250 31.3761
R769 B.n410 B.n409 31.3761
R770 B.n431 B.t9 25.331
R771 B.n545 B.t5 25.331
R772 B B.n587 18.0485
R773 B.n213 B.t3 17.8257
R774 B.t1 B.n576 17.8257
R775 B.n531 B.n52 10.6151
R776 B.n89 B.n52 10.6151
R777 B.n90 B.n89 10.6151
R778 B.n93 B.n90 10.6151
R779 B.n94 B.n93 10.6151
R780 B.n97 B.n94 10.6151
R781 B.n98 B.n97 10.6151
R782 B.n101 B.n98 10.6151
R783 B.n102 B.n101 10.6151
R784 B.n105 B.n102 10.6151
R785 B.n106 B.n105 10.6151
R786 B.n109 B.n106 10.6151
R787 B.n110 B.n109 10.6151
R788 B.n113 B.n110 10.6151
R789 B.n114 B.n113 10.6151
R790 B.n117 B.n114 10.6151
R791 B.n118 B.n117 10.6151
R792 B.n121 B.n118 10.6151
R793 B.n122 B.n121 10.6151
R794 B.n125 B.n122 10.6151
R795 B.n126 B.n125 10.6151
R796 B.n129 B.n126 10.6151
R797 B.n130 B.n129 10.6151
R798 B.n133 B.n130 10.6151
R799 B.n138 B.n135 10.6151
R800 B.n139 B.n138 10.6151
R801 B.n142 B.n139 10.6151
R802 B.n143 B.n142 10.6151
R803 B.n146 B.n143 10.6151
R804 B.n147 B.n146 10.6151
R805 B.n150 B.n147 10.6151
R806 B.n151 B.n150 10.6151
R807 B.n154 B.n151 10.6151
R808 B.n159 B.n156 10.6151
R809 B.n160 B.n159 10.6151
R810 B.n163 B.n160 10.6151
R811 B.n164 B.n163 10.6151
R812 B.n167 B.n164 10.6151
R813 B.n168 B.n167 10.6151
R814 B.n171 B.n168 10.6151
R815 B.n172 B.n171 10.6151
R816 B.n175 B.n172 10.6151
R817 B.n176 B.n175 10.6151
R818 B.n179 B.n176 10.6151
R819 B.n180 B.n179 10.6151
R820 B.n183 B.n180 10.6151
R821 B.n184 B.n183 10.6151
R822 B.n187 B.n184 10.6151
R823 B.n188 B.n187 10.6151
R824 B.n191 B.n188 10.6151
R825 B.n192 B.n191 10.6151
R826 B.n195 B.n192 10.6151
R827 B.n196 B.n195 10.6151
R828 B.n199 B.n196 10.6151
R829 B.n201 B.n199 10.6151
R830 B.n202 B.n201 10.6151
R831 B.n525 B.n202 10.6151
R832 B.n415 B.n250 10.6151
R833 B.n416 B.n415 10.6151
R834 B.n417 B.n416 10.6151
R835 B.n417 B.n241 10.6151
R836 B.n427 B.n241 10.6151
R837 B.n428 B.n427 10.6151
R838 B.n429 B.n428 10.6151
R839 B.n429 B.n234 10.6151
R840 B.n439 B.n234 10.6151
R841 B.n440 B.n439 10.6151
R842 B.n441 B.n440 10.6151
R843 B.n441 B.n226 10.6151
R844 B.n451 B.n226 10.6151
R845 B.n452 B.n451 10.6151
R846 B.n453 B.n452 10.6151
R847 B.n453 B.n219 10.6151
R848 B.n464 B.n219 10.6151
R849 B.n465 B.n464 10.6151
R850 B.n466 B.n465 10.6151
R851 B.n466 B.n210 10.6151
R852 B.n476 B.n210 10.6151
R853 B.n477 B.n476 10.6151
R854 B.n479 B.n477 10.6151
R855 B.n479 B.n478 10.6151
R856 B.n478 B.n203 10.6151
R857 B.n490 B.n203 10.6151
R858 B.n491 B.n490 10.6151
R859 B.n492 B.n491 10.6151
R860 B.n493 B.n492 10.6151
R861 B.n495 B.n493 10.6151
R862 B.n496 B.n495 10.6151
R863 B.n497 B.n496 10.6151
R864 B.n498 B.n497 10.6151
R865 B.n500 B.n498 10.6151
R866 B.n501 B.n500 10.6151
R867 B.n502 B.n501 10.6151
R868 B.n503 B.n502 10.6151
R869 B.n505 B.n503 10.6151
R870 B.n506 B.n505 10.6151
R871 B.n507 B.n506 10.6151
R872 B.n508 B.n507 10.6151
R873 B.n510 B.n508 10.6151
R874 B.n511 B.n510 10.6151
R875 B.n512 B.n511 10.6151
R876 B.n513 B.n512 10.6151
R877 B.n515 B.n513 10.6151
R878 B.n516 B.n515 10.6151
R879 B.n517 B.n516 10.6151
R880 B.n518 B.n517 10.6151
R881 B.n520 B.n518 10.6151
R882 B.n521 B.n520 10.6151
R883 B.n522 B.n521 10.6151
R884 B.n523 B.n522 10.6151
R885 B.n524 B.n523 10.6151
R886 B.n409 B.n254 10.6151
R887 B.n404 B.n254 10.6151
R888 B.n404 B.n403 10.6151
R889 B.n403 B.n402 10.6151
R890 B.n402 B.n399 10.6151
R891 B.n399 B.n398 10.6151
R892 B.n398 B.n395 10.6151
R893 B.n395 B.n394 10.6151
R894 B.n394 B.n391 10.6151
R895 B.n391 B.n390 10.6151
R896 B.n390 B.n387 10.6151
R897 B.n387 B.n386 10.6151
R898 B.n386 B.n383 10.6151
R899 B.n383 B.n382 10.6151
R900 B.n382 B.n379 10.6151
R901 B.n379 B.n378 10.6151
R902 B.n378 B.n375 10.6151
R903 B.n375 B.n374 10.6151
R904 B.n374 B.n371 10.6151
R905 B.n371 B.n370 10.6151
R906 B.n370 B.n367 10.6151
R907 B.n367 B.n366 10.6151
R908 B.n366 B.n363 10.6151
R909 B.n363 B.n362 10.6151
R910 B.n359 B.n358 10.6151
R911 B.n358 B.n355 10.6151
R912 B.n355 B.n354 10.6151
R913 B.n354 B.n351 10.6151
R914 B.n351 B.n350 10.6151
R915 B.n350 B.n347 10.6151
R916 B.n347 B.n346 10.6151
R917 B.n346 B.n343 10.6151
R918 B.n343 B.n342 10.6151
R919 B.n339 B.n338 10.6151
R920 B.n338 B.n335 10.6151
R921 B.n335 B.n334 10.6151
R922 B.n334 B.n331 10.6151
R923 B.n331 B.n330 10.6151
R924 B.n330 B.n327 10.6151
R925 B.n327 B.n326 10.6151
R926 B.n326 B.n323 10.6151
R927 B.n323 B.n322 10.6151
R928 B.n322 B.n319 10.6151
R929 B.n319 B.n318 10.6151
R930 B.n318 B.n315 10.6151
R931 B.n315 B.n314 10.6151
R932 B.n314 B.n311 10.6151
R933 B.n311 B.n310 10.6151
R934 B.n310 B.n307 10.6151
R935 B.n307 B.n306 10.6151
R936 B.n306 B.n303 10.6151
R937 B.n303 B.n302 10.6151
R938 B.n302 B.n299 10.6151
R939 B.n299 B.n298 10.6151
R940 B.n298 B.n295 10.6151
R941 B.n295 B.n294 10.6151
R942 B.n294 B.n292 10.6151
R943 B.n411 B.n410 10.6151
R944 B.n411 B.n246 10.6151
R945 B.n421 B.n246 10.6151
R946 B.n422 B.n421 10.6151
R947 B.n423 B.n422 10.6151
R948 B.n423 B.n238 10.6151
R949 B.n433 B.n238 10.6151
R950 B.n434 B.n433 10.6151
R951 B.n435 B.n434 10.6151
R952 B.n435 B.n230 10.6151
R953 B.n445 B.n230 10.6151
R954 B.n446 B.n445 10.6151
R955 B.n447 B.n446 10.6151
R956 B.n447 B.n222 10.6151
R957 B.n458 B.n222 10.6151
R958 B.n459 B.n458 10.6151
R959 B.n460 B.n459 10.6151
R960 B.n460 B.n215 10.6151
R961 B.n470 B.n215 10.6151
R962 B.n471 B.n470 10.6151
R963 B.n472 B.n471 10.6151
R964 B.n472 B.n207 10.6151
R965 B.n483 B.n207 10.6151
R966 B.n484 B.n483 10.6151
R967 B.n485 B.n484 10.6151
R968 B.n485 B.n0 10.6151
R969 B.n581 B.n1 10.6151
R970 B.n581 B.n580 10.6151
R971 B.n580 B.n579 10.6151
R972 B.n579 B.n10 10.6151
R973 B.n573 B.n10 10.6151
R974 B.n573 B.n572 10.6151
R975 B.n572 B.n571 10.6151
R976 B.n571 B.n17 10.6151
R977 B.n565 B.n17 10.6151
R978 B.n565 B.n564 10.6151
R979 B.n564 B.n563 10.6151
R980 B.n563 B.n23 10.6151
R981 B.n557 B.n23 10.6151
R982 B.n557 B.n556 10.6151
R983 B.n556 B.n555 10.6151
R984 B.n555 B.n31 10.6151
R985 B.n549 B.n31 10.6151
R986 B.n549 B.n548 10.6151
R987 B.n548 B.n547 10.6151
R988 B.n547 B.n38 10.6151
R989 B.n541 B.n38 10.6151
R990 B.n541 B.n540 10.6151
R991 B.n540 B.n539 10.6151
R992 B.n539 B.n45 10.6151
R993 B.n533 B.n45 10.6151
R994 B.n533 B.n532 10.6151
R995 B.n134 B.n133 9.36635
R996 B.n156 B.n155 9.36635
R997 B.n362 B.n288 9.36635
R998 B.n339 B.n291 9.36635
R999 B.n455 B.t0 2.815
R1000 B.n25 B.t2 2.815
R1001 B.n587 B.n0 2.81026
R1002 B.n587 B.n1 2.81026
R1003 B.n135 B.n134 1.24928
R1004 B.n155 B.n154 1.24928
R1005 B.n359 B.n288 1.24928
R1006 B.n342 B.n291 1.24928
R1007 VP.n5 VP.n4 182.832
R1008 VP.n14 VP.n13 182.832
R1009 VP.n12 VP.n0 161.3
R1010 VP.n11 VP.n10 161.3
R1011 VP.n9 VP.n1 161.3
R1012 VP.n8 VP.n7 161.3
R1013 VP.n6 VP.n2 161.3
R1014 VP.n3 VP.t2 123.237
R1015 VP.n3 VP.t3 122.808
R1016 VP.n5 VP.t0 86.8413
R1017 VP.n13 VP.t1 86.8413
R1018 VP.n4 VP.n3 48.8667
R1019 VP.n7 VP.n1 40.4934
R1020 VP.n11 VP.n1 40.4934
R1021 VP.n7 VP.n6 24.4675
R1022 VP.n12 VP.n11 24.4675
R1023 VP.n6 VP.n5 2.93654
R1024 VP.n13 VP.n12 2.93654
R1025 VP.n4 VP.n2 0.189894
R1026 VP.n8 VP.n2 0.189894
R1027 VP.n9 VP.n8 0.189894
R1028 VP.n10 VP.n9 0.189894
R1029 VP.n10 VP.n0 0.189894
R1030 VP.n14 VP.n0 0.189894
R1031 VP VP.n14 0.0516364
R1032 VDD1 VDD1.n1 103.624
R1033 VDD1 VDD1.n0 68.3995
R1034 VDD1.n0 VDD1.t2 3.07027
R1035 VDD1.n0 VDD1.t3 3.07027
R1036 VDD1.n1 VDD1.t1 3.07027
R1037 VDD1.n1 VDD1.t0 3.07027
R1038 VTAIL.n5 VTAIL.t5 54.7324
R1039 VTAIL.n4 VTAIL.t2 54.7324
R1040 VTAIL.n3 VTAIL.t0 54.7324
R1041 VTAIL.n6 VTAIL.t4 54.7323
R1042 VTAIL.n7 VTAIL.t3 54.7323
R1043 VTAIL.n0 VTAIL.t1 54.7323
R1044 VTAIL.n1 VTAIL.t6 54.7323
R1045 VTAIL.n2 VTAIL.t7 54.7323
R1046 VTAIL.n7 VTAIL.n6 19.7548
R1047 VTAIL.n3 VTAIL.n2 19.7548
R1048 VTAIL.n4 VTAIL.n3 1.82809
R1049 VTAIL.n6 VTAIL.n5 1.82809
R1050 VTAIL.n2 VTAIL.n1 1.82809
R1051 VTAIL VTAIL.n0 0.972483
R1052 VTAIL VTAIL.n7 0.856103
R1053 VTAIL.n5 VTAIL.n4 0.470328
R1054 VTAIL.n1 VTAIL.n0 0.470328
R1055 VN.n0 VN.t2 123.237
R1056 VN.n1 VN.t0 123.237
R1057 VN.n0 VN.t3 122.808
R1058 VN.n1 VN.t1 122.808
R1059 VN VN.n1 49.2473
R1060 VN VN.n0 9.34203
R1061 VDD2.n2 VDD2.n0 103.1
R1062 VDD2.n2 VDD2.n1 68.3413
R1063 VDD2.n1 VDD2.t2 3.07027
R1064 VDD2.n1 VDD2.t3 3.07027
R1065 VDD2.n0 VDD2.t1 3.07027
R1066 VDD2.n0 VDD2.t0 3.07027
R1067 VDD2 VDD2.n2 0.0586897
C0 VDD1 VN 0.14809f
C1 VDD2 VN 2.50668f
C2 VP VTAIL 2.62831f
C3 VTAIL VN 2.6142f
C4 VDD2 VDD1 0.8293f
C5 VTAIL VDD1 3.87649f
C6 VDD2 VTAIL 3.92527f
C7 VP VN 4.57933f
C8 VP VDD1 2.70064f
C9 VP VDD2 0.342585f
C10 VDD2 B 2.871164f
C11 VDD1 B 6.1766f
C12 VTAIL B 6.115292f
C13 VN B 8.684099f
C14 VP B 6.725471f
C15 VDD2.t1 B 0.137403f
C16 VDD2.t0 B 0.137403f
C17 VDD2.n0 B 1.58125f
C18 VDD2.t2 B 0.137403f
C19 VDD2.t3 B 0.137403f
C20 VDD2.n1 B 1.15647f
C21 VDD2.n2 B 2.94812f
C22 VN.t2 B 1.22009f
C23 VN.t3 B 1.21811f
C24 VN.n0 B 0.866169f
C25 VN.t0 B 1.22009f
C26 VN.t1 B 1.21811f
C27 VN.n1 B 2.1061f
C28 VTAIL.t1 B 0.940676f
C29 VTAIL.n0 B 0.306154f
C30 VTAIL.t6 B 0.940676f
C31 VTAIL.n1 B 0.356534f
C32 VTAIL.t7 B 0.940676f
C33 VTAIL.n2 B 1.01211f
C34 VTAIL.t0 B 0.940681f
C35 VTAIL.n3 B 1.01211f
C36 VTAIL.t2 B 0.940681f
C37 VTAIL.n4 B 0.356529f
C38 VTAIL.t5 B 0.940681f
C39 VTAIL.n5 B 0.356529f
C40 VTAIL.t4 B 0.940676f
C41 VTAIL.n6 B 1.01211f
C42 VTAIL.t3 B 0.940676f
C43 VTAIL.n7 B 0.954882f
C44 VDD1.t2 B 0.139526f
C45 VDD1.t3 B 0.139526f
C46 VDD1.n0 B 1.17468f
C47 VDD1.t1 B 0.139526f
C48 VDD1.t0 B 0.139526f
C49 VDD1.n1 B 1.62888f
C50 VP.n0 B 0.035182f
C51 VP.t1 B 1.07951f
C52 VP.n1 B 0.028441f
C53 VP.n2 B 0.035182f
C54 VP.t0 B 1.07951f
C55 VP.t2 B 1.25146f
C56 VP.t3 B 1.24943f
C57 VP.n3 B 2.13918f
C58 VP.n4 B 1.64877f
C59 VP.n5 B 0.489658f
C60 VP.n6 B 0.037082f
C61 VP.n7 B 0.069923f
C62 VP.n8 B 0.035182f
C63 VP.n9 B 0.035182f
C64 VP.n10 B 0.035182f
C65 VP.n11 B 0.069923f
C66 VP.n12 B 0.037082f
C67 VP.n13 B 0.489658f
C68 VP.n14 B 0.037655f
.ends

