* NGSPICE file created from diff_pair_sample_1323.ext - technology: sky130A

.subckt diff_pair_sample_1323 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=0.7761 pd=4.76 as=0 ps=0 w=1.99 l=1.97
X1 VDD1.t1 VP.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7761 pd=4.76 as=0.7761 ps=4.76 w=1.99 l=1.97
X2 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=0.7761 pd=4.76 as=0 ps=0 w=1.99 l=1.97
X3 VDD1.t0 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7761 pd=4.76 as=0.7761 ps=4.76 w=1.99 l=1.97
X4 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7761 pd=4.76 as=0.7761 ps=4.76 w=1.99 l=1.97
X5 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7761 pd=4.76 as=0 ps=0 w=1.99 l=1.97
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7761 pd=4.76 as=0 ps=0 w=1.99 l=1.97
X7 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7761 pd=4.76 as=0.7761 ps=4.76 w=1.99 l=1.97
R0 B.n354 B.n353 585
R1 B.n130 B.n59 585
R2 B.n129 B.n128 585
R3 B.n127 B.n126 585
R4 B.n125 B.n124 585
R5 B.n123 B.n122 585
R6 B.n121 B.n120 585
R7 B.n119 B.n118 585
R8 B.n117 B.n116 585
R9 B.n115 B.n114 585
R10 B.n113 B.n112 585
R11 B.n111 B.n110 585
R12 B.n109 B.n108 585
R13 B.n107 B.n106 585
R14 B.n105 B.n104 585
R15 B.n103 B.n102 585
R16 B.n101 B.n100 585
R17 B.n99 B.n98 585
R18 B.n97 B.n96 585
R19 B.n95 B.n94 585
R20 B.n93 B.n92 585
R21 B.n91 B.n90 585
R22 B.n89 B.n88 585
R23 B.n87 B.n86 585
R24 B.n85 B.n84 585
R25 B.n83 B.n82 585
R26 B.n81 B.n80 585
R27 B.n79 B.n78 585
R28 B.n77 B.n76 585
R29 B.n75 B.n74 585
R30 B.n73 B.n72 585
R31 B.n71 B.n70 585
R32 B.n69 B.n68 585
R33 B.n67 B.n66 585
R34 B.n352 B.n42 585
R35 B.n357 B.n42 585
R36 B.n351 B.n41 585
R37 B.n358 B.n41 585
R38 B.n350 B.n349 585
R39 B.n349 B.n37 585
R40 B.n348 B.n36 585
R41 B.n364 B.n36 585
R42 B.n347 B.n35 585
R43 B.n365 B.n35 585
R44 B.n346 B.n34 585
R45 B.n366 B.n34 585
R46 B.n345 B.n344 585
R47 B.n344 B.n33 585
R48 B.n343 B.n29 585
R49 B.n372 B.n29 585
R50 B.n342 B.n28 585
R51 B.n373 B.n28 585
R52 B.n341 B.n27 585
R53 B.n374 B.n27 585
R54 B.n340 B.n339 585
R55 B.n339 B.n23 585
R56 B.n338 B.n22 585
R57 B.n380 B.n22 585
R58 B.n337 B.n21 585
R59 B.n381 B.n21 585
R60 B.n336 B.n20 585
R61 B.n382 B.n20 585
R62 B.n335 B.n334 585
R63 B.n334 B.n16 585
R64 B.n333 B.n15 585
R65 B.n388 B.n15 585
R66 B.n332 B.n14 585
R67 B.n389 B.n14 585
R68 B.n331 B.n13 585
R69 B.n390 B.n13 585
R70 B.n330 B.n329 585
R71 B.n329 B.n12 585
R72 B.n328 B.n327 585
R73 B.n328 B.n8 585
R74 B.n326 B.n7 585
R75 B.n397 B.n7 585
R76 B.n325 B.n6 585
R77 B.n398 B.n6 585
R78 B.n324 B.n5 585
R79 B.n399 B.n5 585
R80 B.n323 B.n322 585
R81 B.n322 B.n4 585
R82 B.n321 B.n131 585
R83 B.n321 B.n320 585
R84 B.n311 B.n132 585
R85 B.n133 B.n132 585
R86 B.n313 B.n312 585
R87 B.n314 B.n313 585
R88 B.n310 B.n137 585
R89 B.n141 B.n137 585
R90 B.n309 B.n308 585
R91 B.n308 B.n307 585
R92 B.n139 B.n138 585
R93 B.n140 B.n139 585
R94 B.n300 B.n299 585
R95 B.n301 B.n300 585
R96 B.n298 B.n146 585
R97 B.n146 B.n145 585
R98 B.n297 B.n296 585
R99 B.n296 B.n295 585
R100 B.n148 B.n147 585
R101 B.n149 B.n148 585
R102 B.n288 B.n287 585
R103 B.n289 B.n288 585
R104 B.n286 B.n154 585
R105 B.n154 B.n153 585
R106 B.n285 B.n284 585
R107 B.n284 B.n283 585
R108 B.n156 B.n155 585
R109 B.n276 B.n156 585
R110 B.n275 B.n274 585
R111 B.n277 B.n275 585
R112 B.n273 B.n161 585
R113 B.n161 B.n160 585
R114 B.n272 B.n271 585
R115 B.n271 B.n270 585
R116 B.n163 B.n162 585
R117 B.n164 B.n163 585
R118 B.n263 B.n262 585
R119 B.n264 B.n263 585
R120 B.n261 B.n169 585
R121 B.n169 B.n168 585
R122 B.n256 B.n255 585
R123 B.n254 B.n188 585
R124 B.n253 B.n187 585
R125 B.n258 B.n187 585
R126 B.n252 B.n251 585
R127 B.n250 B.n249 585
R128 B.n248 B.n247 585
R129 B.n246 B.n245 585
R130 B.n244 B.n243 585
R131 B.n242 B.n241 585
R132 B.n240 B.n239 585
R133 B.n238 B.n237 585
R134 B.n236 B.n235 585
R135 B.n233 B.n232 585
R136 B.n231 B.n230 585
R137 B.n229 B.n228 585
R138 B.n227 B.n226 585
R139 B.n225 B.n224 585
R140 B.n223 B.n222 585
R141 B.n221 B.n220 585
R142 B.n219 B.n218 585
R143 B.n217 B.n216 585
R144 B.n215 B.n214 585
R145 B.n212 B.n211 585
R146 B.n210 B.n209 585
R147 B.n208 B.n207 585
R148 B.n206 B.n205 585
R149 B.n204 B.n203 585
R150 B.n202 B.n201 585
R151 B.n200 B.n199 585
R152 B.n198 B.n197 585
R153 B.n196 B.n195 585
R154 B.n194 B.n193 585
R155 B.n171 B.n170 585
R156 B.n260 B.n259 585
R157 B.n259 B.n258 585
R158 B.n167 B.n166 585
R159 B.n168 B.n167 585
R160 B.n266 B.n265 585
R161 B.n265 B.n264 585
R162 B.n267 B.n165 585
R163 B.n165 B.n164 585
R164 B.n269 B.n268 585
R165 B.n270 B.n269 585
R166 B.n159 B.n158 585
R167 B.n160 B.n159 585
R168 B.n279 B.n278 585
R169 B.n278 B.n277 585
R170 B.n280 B.n157 585
R171 B.n276 B.n157 585
R172 B.n282 B.n281 585
R173 B.n283 B.n282 585
R174 B.n152 B.n151 585
R175 B.n153 B.n152 585
R176 B.n291 B.n290 585
R177 B.n290 B.n289 585
R178 B.n292 B.n150 585
R179 B.n150 B.n149 585
R180 B.n294 B.n293 585
R181 B.n295 B.n294 585
R182 B.n144 B.n143 585
R183 B.n145 B.n144 585
R184 B.n303 B.n302 585
R185 B.n302 B.n301 585
R186 B.n304 B.n142 585
R187 B.n142 B.n140 585
R188 B.n306 B.n305 585
R189 B.n307 B.n306 585
R190 B.n136 B.n135 585
R191 B.n141 B.n136 585
R192 B.n316 B.n315 585
R193 B.n315 B.n314 585
R194 B.n317 B.n134 585
R195 B.n134 B.n133 585
R196 B.n319 B.n318 585
R197 B.n320 B.n319 585
R198 B.n3 B.n0 585
R199 B.n4 B.n3 585
R200 B.n396 B.n1 585
R201 B.n397 B.n396 585
R202 B.n395 B.n394 585
R203 B.n395 B.n8 585
R204 B.n393 B.n9 585
R205 B.n12 B.n9 585
R206 B.n392 B.n391 585
R207 B.n391 B.n390 585
R208 B.n11 B.n10 585
R209 B.n389 B.n11 585
R210 B.n387 B.n386 585
R211 B.n388 B.n387 585
R212 B.n385 B.n17 585
R213 B.n17 B.n16 585
R214 B.n384 B.n383 585
R215 B.n383 B.n382 585
R216 B.n19 B.n18 585
R217 B.n381 B.n19 585
R218 B.n379 B.n378 585
R219 B.n380 B.n379 585
R220 B.n377 B.n24 585
R221 B.n24 B.n23 585
R222 B.n376 B.n375 585
R223 B.n375 B.n374 585
R224 B.n26 B.n25 585
R225 B.n373 B.n26 585
R226 B.n371 B.n370 585
R227 B.n372 B.n371 585
R228 B.n369 B.n30 585
R229 B.n33 B.n30 585
R230 B.n368 B.n367 585
R231 B.n367 B.n366 585
R232 B.n32 B.n31 585
R233 B.n365 B.n32 585
R234 B.n363 B.n362 585
R235 B.n364 B.n363 585
R236 B.n361 B.n38 585
R237 B.n38 B.n37 585
R238 B.n360 B.n359 585
R239 B.n359 B.n358 585
R240 B.n40 B.n39 585
R241 B.n357 B.n40 585
R242 B.n400 B.n399 585
R243 B.n398 B.n2 585
R244 B.n66 B.n40 516.524
R245 B.n354 B.n42 516.524
R246 B.n259 B.n169 516.524
R247 B.n256 B.n167 516.524
R248 B.n356 B.n355 256.663
R249 B.n356 B.n58 256.663
R250 B.n356 B.n57 256.663
R251 B.n356 B.n56 256.663
R252 B.n356 B.n55 256.663
R253 B.n356 B.n54 256.663
R254 B.n356 B.n53 256.663
R255 B.n356 B.n52 256.663
R256 B.n356 B.n51 256.663
R257 B.n356 B.n50 256.663
R258 B.n356 B.n49 256.663
R259 B.n356 B.n48 256.663
R260 B.n356 B.n47 256.663
R261 B.n356 B.n46 256.663
R262 B.n356 B.n45 256.663
R263 B.n356 B.n44 256.663
R264 B.n356 B.n43 256.663
R265 B.n258 B.n257 256.663
R266 B.n258 B.n172 256.663
R267 B.n258 B.n173 256.663
R268 B.n258 B.n174 256.663
R269 B.n258 B.n175 256.663
R270 B.n258 B.n176 256.663
R271 B.n258 B.n177 256.663
R272 B.n258 B.n178 256.663
R273 B.n258 B.n179 256.663
R274 B.n258 B.n180 256.663
R275 B.n258 B.n181 256.663
R276 B.n258 B.n182 256.663
R277 B.n258 B.n183 256.663
R278 B.n258 B.n184 256.663
R279 B.n258 B.n185 256.663
R280 B.n258 B.n186 256.663
R281 B.n402 B.n401 256.663
R282 B.n63 B.t9 231.191
R283 B.n60 B.t13 231.191
R284 B.n191 B.t6 231.191
R285 B.n189 B.t2 231.191
R286 B.n258 B.n168 201.376
R287 B.n357 B.n356 201.376
R288 B.n60 B.t14 167.43
R289 B.n191 B.t8 167.43
R290 B.n63 B.t11 167.43
R291 B.n189 B.t5 167.43
R292 B.n70 B.n69 163.367
R293 B.n74 B.n73 163.367
R294 B.n78 B.n77 163.367
R295 B.n82 B.n81 163.367
R296 B.n86 B.n85 163.367
R297 B.n90 B.n89 163.367
R298 B.n94 B.n93 163.367
R299 B.n98 B.n97 163.367
R300 B.n102 B.n101 163.367
R301 B.n106 B.n105 163.367
R302 B.n110 B.n109 163.367
R303 B.n114 B.n113 163.367
R304 B.n118 B.n117 163.367
R305 B.n122 B.n121 163.367
R306 B.n126 B.n125 163.367
R307 B.n128 B.n59 163.367
R308 B.n263 B.n169 163.367
R309 B.n263 B.n163 163.367
R310 B.n271 B.n163 163.367
R311 B.n271 B.n161 163.367
R312 B.n275 B.n161 163.367
R313 B.n275 B.n156 163.367
R314 B.n284 B.n156 163.367
R315 B.n284 B.n154 163.367
R316 B.n288 B.n154 163.367
R317 B.n288 B.n148 163.367
R318 B.n296 B.n148 163.367
R319 B.n296 B.n146 163.367
R320 B.n300 B.n146 163.367
R321 B.n300 B.n139 163.367
R322 B.n308 B.n139 163.367
R323 B.n308 B.n137 163.367
R324 B.n313 B.n137 163.367
R325 B.n313 B.n132 163.367
R326 B.n321 B.n132 163.367
R327 B.n322 B.n321 163.367
R328 B.n322 B.n5 163.367
R329 B.n6 B.n5 163.367
R330 B.n7 B.n6 163.367
R331 B.n328 B.n7 163.367
R332 B.n329 B.n328 163.367
R333 B.n329 B.n13 163.367
R334 B.n14 B.n13 163.367
R335 B.n15 B.n14 163.367
R336 B.n334 B.n15 163.367
R337 B.n334 B.n20 163.367
R338 B.n21 B.n20 163.367
R339 B.n22 B.n21 163.367
R340 B.n339 B.n22 163.367
R341 B.n339 B.n27 163.367
R342 B.n28 B.n27 163.367
R343 B.n29 B.n28 163.367
R344 B.n344 B.n29 163.367
R345 B.n344 B.n34 163.367
R346 B.n35 B.n34 163.367
R347 B.n36 B.n35 163.367
R348 B.n349 B.n36 163.367
R349 B.n349 B.n41 163.367
R350 B.n42 B.n41 163.367
R351 B.n188 B.n187 163.367
R352 B.n251 B.n187 163.367
R353 B.n249 B.n248 163.367
R354 B.n245 B.n244 163.367
R355 B.n241 B.n240 163.367
R356 B.n237 B.n236 163.367
R357 B.n232 B.n231 163.367
R358 B.n228 B.n227 163.367
R359 B.n224 B.n223 163.367
R360 B.n220 B.n219 163.367
R361 B.n216 B.n215 163.367
R362 B.n211 B.n210 163.367
R363 B.n207 B.n206 163.367
R364 B.n203 B.n202 163.367
R365 B.n199 B.n198 163.367
R366 B.n195 B.n194 163.367
R367 B.n259 B.n171 163.367
R368 B.n265 B.n167 163.367
R369 B.n265 B.n165 163.367
R370 B.n269 B.n165 163.367
R371 B.n269 B.n159 163.367
R372 B.n278 B.n159 163.367
R373 B.n278 B.n157 163.367
R374 B.n282 B.n157 163.367
R375 B.n282 B.n152 163.367
R376 B.n290 B.n152 163.367
R377 B.n290 B.n150 163.367
R378 B.n294 B.n150 163.367
R379 B.n294 B.n144 163.367
R380 B.n302 B.n144 163.367
R381 B.n302 B.n142 163.367
R382 B.n306 B.n142 163.367
R383 B.n306 B.n136 163.367
R384 B.n315 B.n136 163.367
R385 B.n315 B.n134 163.367
R386 B.n319 B.n134 163.367
R387 B.n319 B.n3 163.367
R388 B.n400 B.n3 163.367
R389 B.n396 B.n2 163.367
R390 B.n396 B.n395 163.367
R391 B.n395 B.n9 163.367
R392 B.n391 B.n9 163.367
R393 B.n391 B.n11 163.367
R394 B.n387 B.n11 163.367
R395 B.n387 B.n17 163.367
R396 B.n383 B.n17 163.367
R397 B.n383 B.n19 163.367
R398 B.n379 B.n19 163.367
R399 B.n379 B.n24 163.367
R400 B.n375 B.n24 163.367
R401 B.n375 B.n26 163.367
R402 B.n371 B.n26 163.367
R403 B.n371 B.n30 163.367
R404 B.n367 B.n30 163.367
R405 B.n367 B.n32 163.367
R406 B.n363 B.n32 163.367
R407 B.n363 B.n38 163.367
R408 B.n359 B.n38 163.367
R409 B.n359 B.n40 163.367
R410 B.n61 B.t15 122.825
R411 B.n192 B.t7 122.825
R412 B.n64 B.t12 122.825
R413 B.n190 B.t4 122.825
R414 B.n264 B.n168 102.96
R415 B.n264 B.n164 102.96
R416 B.n270 B.n164 102.96
R417 B.n270 B.n160 102.96
R418 B.n277 B.n160 102.96
R419 B.n277 B.n276 102.96
R420 B.n283 B.n153 102.96
R421 B.n289 B.n153 102.96
R422 B.n289 B.n149 102.96
R423 B.n295 B.n149 102.96
R424 B.n295 B.n145 102.96
R425 B.n301 B.n145 102.96
R426 B.n301 B.n140 102.96
R427 B.n307 B.n140 102.96
R428 B.n307 B.n141 102.96
R429 B.n314 B.n133 102.96
R430 B.n320 B.n133 102.96
R431 B.n320 B.n4 102.96
R432 B.n399 B.n4 102.96
R433 B.n399 B.n398 102.96
R434 B.n398 B.n397 102.96
R435 B.n397 B.n8 102.96
R436 B.n12 B.n8 102.96
R437 B.n390 B.n12 102.96
R438 B.n389 B.n388 102.96
R439 B.n388 B.n16 102.96
R440 B.n382 B.n16 102.96
R441 B.n382 B.n381 102.96
R442 B.n381 B.n380 102.96
R443 B.n380 B.n23 102.96
R444 B.n374 B.n23 102.96
R445 B.n374 B.n373 102.96
R446 B.n373 B.n372 102.96
R447 B.n366 B.n33 102.96
R448 B.n366 B.n365 102.96
R449 B.n365 B.n364 102.96
R450 B.n364 B.n37 102.96
R451 B.n358 B.n37 102.96
R452 B.n358 B.n357 102.96
R453 B.n66 B.n43 71.676
R454 B.n70 B.n44 71.676
R455 B.n74 B.n45 71.676
R456 B.n78 B.n46 71.676
R457 B.n82 B.n47 71.676
R458 B.n86 B.n48 71.676
R459 B.n90 B.n49 71.676
R460 B.n94 B.n50 71.676
R461 B.n98 B.n51 71.676
R462 B.n102 B.n52 71.676
R463 B.n106 B.n53 71.676
R464 B.n110 B.n54 71.676
R465 B.n114 B.n55 71.676
R466 B.n118 B.n56 71.676
R467 B.n122 B.n57 71.676
R468 B.n126 B.n58 71.676
R469 B.n355 B.n59 71.676
R470 B.n355 B.n354 71.676
R471 B.n128 B.n58 71.676
R472 B.n125 B.n57 71.676
R473 B.n121 B.n56 71.676
R474 B.n117 B.n55 71.676
R475 B.n113 B.n54 71.676
R476 B.n109 B.n53 71.676
R477 B.n105 B.n52 71.676
R478 B.n101 B.n51 71.676
R479 B.n97 B.n50 71.676
R480 B.n93 B.n49 71.676
R481 B.n89 B.n48 71.676
R482 B.n85 B.n47 71.676
R483 B.n81 B.n46 71.676
R484 B.n77 B.n45 71.676
R485 B.n73 B.n44 71.676
R486 B.n69 B.n43 71.676
R487 B.n257 B.n256 71.676
R488 B.n251 B.n172 71.676
R489 B.n248 B.n173 71.676
R490 B.n244 B.n174 71.676
R491 B.n240 B.n175 71.676
R492 B.n236 B.n176 71.676
R493 B.n231 B.n177 71.676
R494 B.n227 B.n178 71.676
R495 B.n223 B.n179 71.676
R496 B.n219 B.n180 71.676
R497 B.n215 B.n181 71.676
R498 B.n210 B.n182 71.676
R499 B.n206 B.n183 71.676
R500 B.n202 B.n184 71.676
R501 B.n198 B.n185 71.676
R502 B.n194 B.n186 71.676
R503 B.n257 B.n188 71.676
R504 B.n249 B.n172 71.676
R505 B.n245 B.n173 71.676
R506 B.n241 B.n174 71.676
R507 B.n237 B.n175 71.676
R508 B.n232 B.n176 71.676
R509 B.n228 B.n177 71.676
R510 B.n224 B.n178 71.676
R511 B.n220 B.n179 71.676
R512 B.n216 B.n180 71.676
R513 B.n211 B.n181 71.676
R514 B.n207 B.n182 71.676
R515 B.n203 B.n183 71.676
R516 B.n199 B.n184 71.676
R517 B.n195 B.n185 71.676
R518 B.n186 B.n171 71.676
R519 B.n401 B.n400 71.676
R520 B.n401 B.n2 71.676
R521 B.n65 B.n64 59.5399
R522 B.n62 B.n61 59.5399
R523 B.n213 B.n192 59.5399
R524 B.n234 B.n190 59.5399
R525 B.n276 B.t3 56.0225
R526 B.n33 B.t10 56.0225
R527 B.n141 B.t0 52.9943
R528 B.t1 B.n389 52.9943
R529 B.n314 B.t0 49.9661
R530 B.n390 B.t1 49.9661
R531 B.n283 B.t3 46.9379
R532 B.n372 B.t10 46.9379
R533 B.n64 B.n63 44.6066
R534 B.n61 B.n60 44.6066
R535 B.n192 B.n191 44.6066
R536 B.n190 B.n189 44.6066
R537 B.n255 B.n166 33.5615
R538 B.n261 B.n260 33.5615
R539 B.n353 B.n352 33.5615
R540 B.n67 B.n39 33.5615
R541 B B.n402 18.0485
R542 B.n266 B.n166 10.6151
R543 B.n267 B.n266 10.6151
R544 B.n268 B.n267 10.6151
R545 B.n268 B.n158 10.6151
R546 B.n279 B.n158 10.6151
R547 B.n280 B.n279 10.6151
R548 B.n281 B.n280 10.6151
R549 B.n281 B.n151 10.6151
R550 B.n291 B.n151 10.6151
R551 B.n292 B.n291 10.6151
R552 B.n293 B.n292 10.6151
R553 B.n293 B.n143 10.6151
R554 B.n303 B.n143 10.6151
R555 B.n304 B.n303 10.6151
R556 B.n305 B.n304 10.6151
R557 B.n305 B.n135 10.6151
R558 B.n316 B.n135 10.6151
R559 B.n317 B.n316 10.6151
R560 B.n318 B.n317 10.6151
R561 B.n318 B.n0 10.6151
R562 B.n255 B.n254 10.6151
R563 B.n254 B.n253 10.6151
R564 B.n253 B.n252 10.6151
R565 B.n252 B.n250 10.6151
R566 B.n250 B.n247 10.6151
R567 B.n247 B.n246 10.6151
R568 B.n246 B.n243 10.6151
R569 B.n243 B.n242 10.6151
R570 B.n242 B.n239 10.6151
R571 B.n239 B.n238 10.6151
R572 B.n238 B.n235 10.6151
R573 B.n233 B.n230 10.6151
R574 B.n230 B.n229 10.6151
R575 B.n229 B.n226 10.6151
R576 B.n226 B.n225 10.6151
R577 B.n225 B.n222 10.6151
R578 B.n222 B.n221 10.6151
R579 B.n221 B.n218 10.6151
R580 B.n218 B.n217 10.6151
R581 B.n217 B.n214 10.6151
R582 B.n212 B.n209 10.6151
R583 B.n209 B.n208 10.6151
R584 B.n208 B.n205 10.6151
R585 B.n205 B.n204 10.6151
R586 B.n204 B.n201 10.6151
R587 B.n201 B.n200 10.6151
R588 B.n200 B.n197 10.6151
R589 B.n197 B.n196 10.6151
R590 B.n196 B.n193 10.6151
R591 B.n193 B.n170 10.6151
R592 B.n260 B.n170 10.6151
R593 B.n262 B.n261 10.6151
R594 B.n262 B.n162 10.6151
R595 B.n272 B.n162 10.6151
R596 B.n273 B.n272 10.6151
R597 B.n274 B.n273 10.6151
R598 B.n274 B.n155 10.6151
R599 B.n285 B.n155 10.6151
R600 B.n286 B.n285 10.6151
R601 B.n287 B.n286 10.6151
R602 B.n287 B.n147 10.6151
R603 B.n297 B.n147 10.6151
R604 B.n298 B.n297 10.6151
R605 B.n299 B.n298 10.6151
R606 B.n299 B.n138 10.6151
R607 B.n309 B.n138 10.6151
R608 B.n310 B.n309 10.6151
R609 B.n312 B.n310 10.6151
R610 B.n312 B.n311 10.6151
R611 B.n311 B.n131 10.6151
R612 B.n323 B.n131 10.6151
R613 B.n324 B.n323 10.6151
R614 B.n325 B.n324 10.6151
R615 B.n326 B.n325 10.6151
R616 B.n327 B.n326 10.6151
R617 B.n330 B.n327 10.6151
R618 B.n331 B.n330 10.6151
R619 B.n332 B.n331 10.6151
R620 B.n333 B.n332 10.6151
R621 B.n335 B.n333 10.6151
R622 B.n336 B.n335 10.6151
R623 B.n337 B.n336 10.6151
R624 B.n338 B.n337 10.6151
R625 B.n340 B.n338 10.6151
R626 B.n341 B.n340 10.6151
R627 B.n342 B.n341 10.6151
R628 B.n343 B.n342 10.6151
R629 B.n345 B.n343 10.6151
R630 B.n346 B.n345 10.6151
R631 B.n347 B.n346 10.6151
R632 B.n348 B.n347 10.6151
R633 B.n350 B.n348 10.6151
R634 B.n351 B.n350 10.6151
R635 B.n352 B.n351 10.6151
R636 B.n394 B.n1 10.6151
R637 B.n394 B.n393 10.6151
R638 B.n393 B.n392 10.6151
R639 B.n392 B.n10 10.6151
R640 B.n386 B.n10 10.6151
R641 B.n386 B.n385 10.6151
R642 B.n385 B.n384 10.6151
R643 B.n384 B.n18 10.6151
R644 B.n378 B.n18 10.6151
R645 B.n378 B.n377 10.6151
R646 B.n377 B.n376 10.6151
R647 B.n376 B.n25 10.6151
R648 B.n370 B.n25 10.6151
R649 B.n370 B.n369 10.6151
R650 B.n369 B.n368 10.6151
R651 B.n368 B.n31 10.6151
R652 B.n362 B.n31 10.6151
R653 B.n362 B.n361 10.6151
R654 B.n361 B.n360 10.6151
R655 B.n360 B.n39 10.6151
R656 B.n68 B.n67 10.6151
R657 B.n71 B.n68 10.6151
R658 B.n72 B.n71 10.6151
R659 B.n75 B.n72 10.6151
R660 B.n76 B.n75 10.6151
R661 B.n79 B.n76 10.6151
R662 B.n80 B.n79 10.6151
R663 B.n83 B.n80 10.6151
R664 B.n84 B.n83 10.6151
R665 B.n87 B.n84 10.6151
R666 B.n88 B.n87 10.6151
R667 B.n92 B.n91 10.6151
R668 B.n95 B.n92 10.6151
R669 B.n96 B.n95 10.6151
R670 B.n99 B.n96 10.6151
R671 B.n100 B.n99 10.6151
R672 B.n103 B.n100 10.6151
R673 B.n104 B.n103 10.6151
R674 B.n107 B.n104 10.6151
R675 B.n108 B.n107 10.6151
R676 B.n112 B.n111 10.6151
R677 B.n115 B.n112 10.6151
R678 B.n116 B.n115 10.6151
R679 B.n119 B.n116 10.6151
R680 B.n120 B.n119 10.6151
R681 B.n123 B.n120 10.6151
R682 B.n124 B.n123 10.6151
R683 B.n127 B.n124 10.6151
R684 B.n129 B.n127 10.6151
R685 B.n130 B.n129 10.6151
R686 B.n353 B.n130 10.6151
R687 B.n235 B.n234 9.36635
R688 B.n213 B.n212 9.36635
R689 B.n88 B.n65 9.36635
R690 B.n111 B.n62 9.36635
R691 B.n402 B.n0 8.11757
R692 B.n402 B.n1 8.11757
R693 B.n234 B.n233 1.24928
R694 B.n214 B.n213 1.24928
R695 B.n91 B.n65 1.24928
R696 B.n108 B.n62 1.24928
R697 VP.n0 VP.t1 118.609
R698 VP.n0 VP.t0 83.2059
R699 VP VP.n0 0.241678
R700 VTAIL.n26 VTAIL.n24 289.615
R701 VTAIL.n2 VTAIL.n0 289.615
R702 VTAIL.n18 VTAIL.n16 289.615
R703 VTAIL.n10 VTAIL.n8 289.615
R704 VTAIL.n27 VTAIL.n26 185
R705 VTAIL.n3 VTAIL.n2 185
R706 VTAIL.n19 VTAIL.n18 185
R707 VTAIL.n11 VTAIL.n10 185
R708 VTAIL.t1 VTAIL.n25 167.117
R709 VTAIL.t2 VTAIL.n1 167.117
R710 VTAIL.t3 VTAIL.n17 167.117
R711 VTAIL.t0 VTAIL.n9 167.117
R712 VTAIL.n26 VTAIL.t1 52.3082
R713 VTAIL.n2 VTAIL.t2 52.3082
R714 VTAIL.n18 VTAIL.t3 52.3082
R715 VTAIL.n10 VTAIL.t0 52.3082
R716 VTAIL.n31 VTAIL.n30 31.2157
R717 VTAIL.n7 VTAIL.n6 31.2157
R718 VTAIL.n23 VTAIL.n22 31.2157
R719 VTAIL.n15 VTAIL.n14 31.2157
R720 VTAIL.n15 VTAIL.n7 18.0479
R721 VTAIL.n31 VTAIL.n23 16.0652
R722 VTAIL.n27 VTAIL.n25 9.71174
R723 VTAIL.n3 VTAIL.n1 9.71174
R724 VTAIL.n19 VTAIL.n17 9.71174
R725 VTAIL.n11 VTAIL.n9 9.71174
R726 VTAIL.n30 VTAIL.n29 9.45567
R727 VTAIL.n6 VTAIL.n5 9.45567
R728 VTAIL.n22 VTAIL.n21 9.45567
R729 VTAIL.n14 VTAIL.n13 9.45567
R730 VTAIL.n29 VTAIL.n28 9.3005
R731 VTAIL.n5 VTAIL.n4 9.3005
R732 VTAIL.n21 VTAIL.n20 9.3005
R733 VTAIL.n13 VTAIL.n12 9.3005
R734 VTAIL.n30 VTAIL.n24 8.14595
R735 VTAIL.n6 VTAIL.n0 8.14595
R736 VTAIL.n22 VTAIL.n16 8.14595
R737 VTAIL.n14 VTAIL.n8 8.14595
R738 VTAIL.n28 VTAIL.n27 7.3702
R739 VTAIL.n4 VTAIL.n3 7.3702
R740 VTAIL.n20 VTAIL.n19 7.3702
R741 VTAIL.n12 VTAIL.n11 7.3702
R742 VTAIL.n28 VTAIL.n24 5.81868
R743 VTAIL.n4 VTAIL.n0 5.81868
R744 VTAIL.n20 VTAIL.n16 5.81868
R745 VTAIL.n12 VTAIL.n8 5.81868
R746 VTAIL.n29 VTAIL.n25 3.44771
R747 VTAIL.n5 VTAIL.n1 3.44771
R748 VTAIL.n21 VTAIL.n17 3.44771
R749 VTAIL.n13 VTAIL.n9 3.44771
R750 VTAIL.n23 VTAIL.n15 1.46171
R751 VTAIL VTAIL.n7 1.02421
R752 VTAIL VTAIL.n31 0.438
R753 VDD1.n2 VDD1.n0 289.615
R754 VDD1.n9 VDD1.n7 289.615
R755 VDD1.n3 VDD1.n2 185
R756 VDD1.n10 VDD1.n9 185
R757 VDD1.t0 VDD1.n1 167.117
R758 VDD1.t1 VDD1.n8 167.117
R759 VDD1 VDD1.n13 78.2554
R760 VDD1.n2 VDD1.t0 52.3082
R761 VDD1.n9 VDD1.t1 52.3082
R762 VDD1 VDD1.n6 48.4483
R763 VDD1.n3 VDD1.n1 9.71174
R764 VDD1.n10 VDD1.n8 9.71174
R765 VDD1.n6 VDD1.n5 9.45567
R766 VDD1.n13 VDD1.n12 9.45567
R767 VDD1.n5 VDD1.n4 9.3005
R768 VDD1.n12 VDD1.n11 9.3005
R769 VDD1.n6 VDD1.n0 8.14595
R770 VDD1.n13 VDD1.n7 8.14595
R771 VDD1.n4 VDD1.n3 7.3702
R772 VDD1.n11 VDD1.n10 7.3702
R773 VDD1.n4 VDD1.n0 5.81868
R774 VDD1.n11 VDD1.n7 5.81868
R775 VDD1.n5 VDD1.n1 3.44771
R776 VDD1.n12 VDD1.n8 3.44771
R777 VN VN.t0 118.799
R778 VN VN.t1 83.4471
R779 VDD2.n9 VDD2.n7 289.615
R780 VDD2.n2 VDD2.n0 289.615
R781 VDD2.n10 VDD2.n9 185
R782 VDD2.n3 VDD2.n2 185
R783 VDD2.t1 VDD2.n8 167.117
R784 VDD2.t0 VDD2.n1 167.117
R785 VDD2.n14 VDD2.n6 77.2349
R786 VDD2.n9 VDD2.t1 52.3082
R787 VDD2.n2 VDD2.t0 52.3082
R788 VDD2.n14 VDD2.n13 47.8944
R789 VDD2.n10 VDD2.n8 9.71174
R790 VDD2.n3 VDD2.n1 9.71174
R791 VDD2.n13 VDD2.n12 9.45567
R792 VDD2.n6 VDD2.n5 9.45567
R793 VDD2.n12 VDD2.n11 9.3005
R794 VDD2.n5 VDD2.n4 9.3005
R795 VDD2.n13 VDD2.n7 8.14595
R796 VDD2.n6 VDD2.n0 8.14595
R797 VDD2.n11 VDD2.n10 7.3702
R798 VDD2.n4 VDD2.n3 7.3702
R799 VDD2.n11 VDD2.n7 5.81868
R800 VDD2.n4 VDD2.n0 5.81868
R801 VDD2.n12 VDD2.n8 3.44771
R802 VDD2.n5 VDD2.n1 3.44771
R803 VDD2 VDD2.n14 0.554379
C0 VN VDD1 0.154145f
C1 VDD2 VN 0.649116f
C2 VTAIL VDD1 2.22574f
C3 VDD2 VTAIL 2.2743f
C4 VN VP 3.31199f
C5 VDD2 VDD1 0.598364f
C6 VTAIL VP 0.867925f
C7 VN VTAIL 0.853777f
C8 VP VDD1 0.806161f
C9 VDD2 VP 0.31271f
C10 VDD2 B 2.377634f
C11 VDD1 B 3.78336f
C12 VTAIL B 2.780811f
C13 VN B 6.77614f
C14 VP B 4.738392f
C15 VDD2.n0 B 0.025187f
C16 VDD2.n1 B 0.055769f
C17 VDD2.t0 B 0.041869f
C18 VDD2.n2 B 0.043612f
C19 VDD2.n3 B 0.014125f
C20 VDD2.n4 B 0.009316f
C21 VDD2.n5 B 0.122702f
C22 VDD2.n6 B 0.269957f
C23 VDD2.n7 B 0.025187f
C24 VDD2.n8 B 0.055769f
C25 VDD2.t1 B 0.041869f
C26 VDD2.n9 B 0.043612f
C27 VDD2.n10 B 0.014125f
C28 VDD2.n11 B 0.009316f
C29 VDD2.n12 B 0.122702f
C30 VDD2.n13 B 0.039575f
C31 VDD2.n14 B 1.2785f
C32 VN.t1 B 0.506802f
C33 VN.t0 B 0.842328f
C34 VDD1.n0 B 0.023439f
C35 VDD1.n1 B 0.0519f
C36 VDD1.t0 B 0.038964f
C37 VDD1.n2 B 0.040586f
C38 VDD1.n3 B 0.013145f
C39 VDD1.n4 B 0.00867f
C40 VDD1.n5 B 0.114188f
C41 VDD1.n6 B 0.037506f
C42 VDD1.n7 B 0.023439f
C43 VDD1.n8 B 0.0519f
C44 VDD1.t1 B 0.038964f
C45 VDD1.n9 B 0.040586f
C46 VDD1.n10 B 0.013145f
C47 VDD1.n11 B 0.00867f
C48 VDD1.n12 B 0.114188f
C49 VDD1.n13 B 0.273806f
C50 VTAIL.n0 B 0.030357f
C51 VTAIL.n1 B 0.067216f
C52 VTAIL.t2 B 0.050463f
C53 VTAIL.n2 B 0.052563f
C54 VTAIL.n3 B 0.017025f
C55 VTAIL.n4 B 0.011228f
C56 VTAIL.n5 B 0.147887f
C57 VTAIL.n6 B 0.033258f
C58 VTAIL.n7 B 0.752295f
C59 VTAIL.n8 B 0.030357f
C60 VTAIL.n9 B 0.067216f
C61 VTAIL.t0 B 0.050463f
C62 VTAIL.n10 B 0.052563f
C63 VTAIL.n11 B 0.017025f
C64 VTAIL.n12 B 0.011228f
C65 VTAIL.n13 B 0.147887f
C66 VTAIL.n14 B 0.033258f
C67 VTAIL.n15 B 0.781752f
C68 VTAIL.n16 B 0.030357f
C69 VTAIL.n17 B 0.067216f
C70 VTAIL.t3 B 0.050463f
C71 VTAIL.n18 B 0.052563f
C72 VTAIL.n19 B 0.017025f
C73 VTAIL.n20 B 0.011228f
C74 VTAIL.n21 B 0.147887f
C75 VTAIL.n22 B 0.033258f
C76 VTAIL.n23 B 0.648255f
C77 VTAIL.n24 B 0.030357f
C78 VTAIL.n25 B 0.067216f
C79 VTAIL.t1 B 0.050463f
C80 VTAIL.n26 B 0.052563f
C81 VTAIL.n27 B 0.017025f
C82 VTAIL.n28 B 0.011228f
C83 VTAIL.n29 B 0.147887f
C84 VTAIL.n30 B 0.033258f
C85 VTAIL.n31 B 0.579331f
C86 VP.t1 B 0.847676f
C87 VP.t0 B 0.513043f
C88 VP.n0 B 1.88739f
.ends

