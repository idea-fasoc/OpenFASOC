* NGSPICE file created from diff_pair_sample_1562.ext - technology: sky130A

.subckt diff_pair_sample_1562 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=0.234 pd=1.98 as=0 ps=0 w=0.6 l=0.68
X1 VDD2.t9 VN.t0 VTAIL.t19 B.t3 sky130_fd_pr__nfet_01v8 ad=0.099 pd=0.93 as=0.099 ps=0.93 w=0.6 l=0.68
X2 VTAIL.t5 VP.t0 VDD1.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=0.099 pd=0.93 as=0.099 ps=0.93 w=0.6 l=0.68
X3 VDD1.t8 VP.t1 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=0.234 pd=1.98 as=0.099 ps=0.93 w=0.6 l=0.68
X4 VTAIL.t18 VN.t1 VDD2.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=0.099 pd=0.93 as=0.099 ps=0.93 w=0.6 l=0.68
X5 VDD1.t7 VP.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.099 pd=0.93 as=0.234 ps=1.98 w=0.6 l=0.68
X6 VTAIL.t13 VN.t2 VDD2.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=0.099 pd=0.93 as=0.099 ps=0.93 w=0.6 l=0.68
X7 VDD2.t6 VN.t3 VTAIL.t11 B.t9 sky130_fd_pr__nfet_01v8 ad=0.234 pd=1.98 as=0.099 ps=0.93 w=0.6 l=0.68
X8 VDD1.t6 VP.t3 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=0.234 pd=1.98 as=0.099 ps=0.93 w=0.6 l=0.68
X9 VDD2.t5 VN.t4 VTAIL.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=0.234 pd=1.98 as=0.099 ps=0.93 w=0.6 l=0.68
X10 VDD2.t4 VN.t5 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=0.099 pd=0.93 as=0.234 ps=1.98 w=0.6 l=0.68
X11 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=0.234 pd=1.98 as=0 ps=0 w=0.6 l=0.68
X12 VTAIL.t14 VN.t6 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.099 pd=0.93 as=0.099 ps=0.93 w=0.6 l=0.68
X13 VDD2.t2 VN.t7 VTAIL.t17 B.t4 sky130_fd_pr__nfet_01v8 ad=0.099 pd=0.93 as=0.099 ps=0.93 w=0.6 l=0.68
X14 VTAIL.t1 VP.t4 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.099 pd=0.93 as=0.099 ps=0.93 w=0.6 l=0.68
X15 VDD2.t1 VN.t8 VTAIL.t12 B.t0 sky130_fd_pr__nfet_01v8 ad=0.099 pd=0.93 as=0.234 ps=1.98 w=0.6 l=0.68
X16 VTAIL.t15 VN.t9 VDD2.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=0.099 pd=0.93 as=0.099 ps=0.93 w=0.6 l=0.68
X17 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=0.234 pd=1.98 as=0 ps=0 w=0.6 l=0.68
X18 VDD1.t4 VP.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.099 pd=0.93 as=0.099 ps=0.93 w=0.6 l=0.68
X19 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.234 pd=1.98 as=0 ps=0 w=0.6 l=0.68
X20 VDD1.t3 VP.t6 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.099 pd=0.93 as=0.234 ps=1.98 w=0.6 l=0.68
X21 VTAIL.t2 VP.t7 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.099 pd=0.93 as=0.099 ps=0.93 w=0.6 l=0.68
X22 VDD1.t1 VP.t8 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.099 pd=0.93 as=0.099 ps=0.93 w=0.6 l=0.68
X23 VTAIL.t6 VP.t9 VDD1.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=0.099 pd=0.93 as=0.099 ps=0.93 w=0.6 l=0.68
R0 B.n300 B.n299 585
R1 B.n302 B.n68 585
R2 B.n305 B.n304 585
R3 B.n306 B.n67 585
R4 B.n308 B.n307 585
R5 B.n310 B.n66 585
R6 B.n312 B.n311 585
R7 B.n314 B.n313 585
R8 B.n317 B.n316 585
R9 B.n318 B.n61 585
R10 B.n320 B.n319 585
R11 B.n322 B.n60 585
R12 B.n325 B.n324 585
R13 B.n326 B.n59 585
R14 B.n328 B.n327 585
R15 B.n330 B.n58 585
R16 B.n333 B.n332 585
R17 B.n334 B.n55 585
R18 B.n337 B.n336 585
R19 B.n339 B.n54 585
R20 B.n342 B.n341 585
R21 B.n343 B.n53 585
R22 B.n345 B.n344 585
R23 B.n347 B.n52 585
R24 B.n350 B.n349 585
R25 B.n351 B.n51 585
R26 B.n298 B.n49 585
R27 B.n354 B.n49 585
R28 B.n297 B.n48 585
R29 B.n355 B.n48 585
R30 B.n296 B.n47 585
R31 B.n356 B.n47 585
R32 B.n295 B.n294 585
R33 B.n294 B.n43 585
R34 B.n293 B.n42 585
R35 B.n362 B.n42 585
R36 B.n292 B.n41 585
R37 B.n363 B.n41 585
R38 B.n291 B.n40 585
R39 B.n364 B.n40 585
R40 B.n290 B.n289 585
R41 B.n289 B.n36 585
R42 B.n288 B.n35 585
R43 B.n370 B.n35 585
R44 B.n287 B.n34 585
R45 B.n371 B.n34 585
R46 B.n286 B.n33 585
R47 B.n372 B.n33 585
R48 B.n285 B.n284 585
R49 B.n284 B.n32 585
R50 B.n283 B.n28 585
R51 B.n378 B.n28 585
R52 B.n282 B.n27 585
R53 B.n379 B.n27 585
R54 B.n281 B.n26 585
R55 B.t1 B.n26 585
R56 B.n280 B.n279 585
R57 B.n279 B.n22 585
R58 B.n278 B.n21 585
R59 B.n385 B.n21 585
R60 B.n277 B.n20 585
R61 B.n386 B.n20 585
R62 B.n276 B.n19 585
R63 B.n387 B.n19 585
R64 B.n275 B.n274 585
R65 B.n274 B.n18 585
R66 B.n273 B.n14 585
R67 B.n393 B.n14 585
R68 B.n272 B.n13 585
R69 B.n394 B.n13 585
R70 B.n271 B.n12 585
R71 B.n395 B.n12 585
R72 B.n270 B.n269 585
R73 B.n269 B.n8 585
R74 B.n268 B.n7 585
R75 B.n401 B.n7 585
R76 B.n267 B.n6 585
R77 B.n402 B.n6 585
R78 B.n266 B.n5 585
R79 B.n403 B.n5 585
R80 B.n265 B.n264 585
R81 B.n264 B.n4 585
R82 B.n263 B.n69 585
R83 B.n263 B.n262 585
R84 B.n253 B.n70 585
R85 B.n71 B.n70 585
R86 B.n255 B.n254 585
R87 B.n256 B.n255 585
R88 B.n252 B.n76 585
R89 B.n76 B.n75 585
R90 B.n251 B.n250 585
R91 B.n250 B.n249 585
R92 B.n78 B.n77 585
R93 B.n242 B.n78 585
R94 B.n241 B.n240 585
R95 B.n243 B.n241 585
R96 B.n239 B.n83 585
R97 B.n83 B.n82 585
R98 B.n238 B.n237 585
R99 B.n237 B.n236 585
R100 B.n85 B.n84 585
R101 B.n86 B.n85 585
R102 B.n230 B.n229 585
R103 B.t6 B.n230 585
R104 B.n228 B.n91 585
R105 B.n91 B.n90 585
R106 B.n227 B.n226 585
R107 B.n226 B.n225 585
R108 B.n93 B.n92 585
R109 B.n218 B.n93 585
R110 B.n217 B.n216 585
R111 B.n219 B.n217 585
R112 B.n215 B.n98 585
R113 B.n98 B.n97 585
R114 B.n214 B.n213 585
R115 B.n213 B.n212 585
R116 B.n100 B.n99 585
R117 B.n101 B.n100 585
R118 B.n205 B.n204 585
R119 B.n206 B.n205 585
R120 B.n203 B.n106 585
R121 B.n106 B.n105 585
R122 B.n202 B.n201 585
R123 B.n201 B.n200 585
R124 B.n108 B.n107 585
R125 B.n109 B.n108 585
R126 B.n193 B.n192 585
R127 B.n194 B.n193 585
R128 B.n191 B.n114 585
R129 B.n114 B.n113 585
R130 B.n190 B.n189 585
R131 B.n189 B.n188 585
R132 B.n185 B.n118 585
R133 B.n184 B.n183 585
R134 B.n181 B.n119 585
R135 B.n181 B.n117 585
R136 B.n180 B.n179 585
R137 B.n178 B.n177 585
R138 B.n176 B.n121 585
R139 B.n174 B.n173 585
R140 B.n172 B.n122 585
R141 B.n170 B.n169 585
R142 B.n167 B.n125 585
R143 B.n165 B.n164 585
R144 B.n163 B.n126 585
R145 B.n162 B.n161 585
R146 B.n159 B.n127 585
R147 B.n157 B.n156 585
R148 B.n155 B.n128 585
R149 B.n154 B.n153 585
R150 B.n151 B.n129 585
R151 B.n149 B.n148 585
R152 B.n147 B.n130 585
R153 B.n146 B.n145 585
R154 B.n143 B.n134 585
R155 B.n141 B.n140 585
R156 B.n139 B.n135 585
R157 B.n138 B.n137 585
R158 B.n116 B.n115 585
R159 B.n117 B.n116 585
R160 B.n187 B.n186 585
R161 B.n188 B.n187 585
R162 B.n112 B.n111 585
R163 B.n113 B.n112 585
R164 B.n196 B.n195 585
R165 B.n195 B.n194 585
R166 B.n197 B.n110 585
R167 B.n110 B.n109 585
R168 B.n199 B.n198 585
R169 B.n200 B.n199 585
R170 B.n104 B.n103 585
R171 B.n105 B.n104 585
R172 B.n208 B.n207 585
R173 B.n207 B.n206 585
R174 B.n209 B.n102 585
R175 B.n102 B.n101 585
R176 B.n211 B.n210 585
R177 B.n212 B.n211 585
R178 B.n96 B.n95 585
R179 B.n97 B.n96 585
R180 B.n221 B.n220 585
R181 B.n220 B.n219 585
R182 B.n222 B.n94 585
R183 B.n218 B.n94 585
R184 B.n224 B.n223 585
R185 B.n225 B.n224 585
R186 B.n89 B.n88 585
R187 B.n90 B.n89 585
R188 B.n232 B.n231 585
R189 B.n231 B.t6 585
R190 B.n233 B.n87 585
R191 B.n87 B.n86 585
R192 B.n235 B.n234 585
R193 B.n236 B.n235 585
R194 B.n81 B.n80 585
R195 B.n82 B.n81 585
R196 B.n245 B.n244 585
R197 B.n244 B.n243 585
R198 B.n246 B.n79 585
R199 B.n242 B.n79 585
R200 B.n248 B.n247 585
R201 B.n249 B.n248 585
R202 B.n74 B.n73 585
R203 B.n75 B.n74 585
R204 B.n258 B.n257 585
R205 B.n257 B.n256 585
R206 B.n259 B.n72 585
R207 B.n72 B.n71 585
R208 B.n261 B.n260 585
R209 B.n262 B.n261 585
R210 B.n2 B.n0 585
R211 B.n4 B.n2 585
R212 B.n3 B.n1 585
R213 B.n402 B.n3 585
R214 B.n400 B.n399 585
R215 B.n401 B.n400 585
R216 B.n398 B.n9 585
R217 B.n9 B.n8 585
R218 B.n397 B.n396 585
R219 B.n396 B.n395 585
R220 B.n11 B.n10 585
R221 B.n394 B.n11 585
R222 B.n392 B.n391 585
R223 B.n393 B.n392 585
R224 B.n390 B.n15 585
R225 B.n18 B.n15 585
R226 B.n389 B.n388 585
R227 B.n388 B.n387 585
R228 B.n17 B.n16 585
R229 B.n386 B.n17 585
R230 B.n384 B.n383 585
R231 B.n385 B.n384 585
R232 B.n382 B.n23 585
R233 B.n23 B.n22 585
R234 B.n381 B.n380 585
R235 B.n380 B.t1 585
R236 B.n25 B.n24 585
R237 B.n379 B.n25 585
R238 B.n377 B.n376 585
R239 B.n378 B.n377 585
R240 B.n375 B.n29 585
R241 B.n32 B.n29 585
R242 B.n374 B.n373 585
R243 B.n373 B.n372 585
R244 B.n31 B.n30 585
R245 B.n371 B.n31 585
R246 B.n369 B.n368 585
R247 B.n370 B.n369 585
R248 B.n367 B.n37 585
R249 B.n37 B.n36 585
R250 B.n366 B.n365 585
R251 B.n365 B.n364 585
R252 B.n39 B.n38 585
R253 B.n363 B.n39 585
R254 B.n361 B.n360 585
R255 B.n362 B.n361 585
R256 B.n359 B.n44 585
R257 B.n44 B.n43 585
R258 B.n358 B.n357 585
R259 B.n357 B.n356 585
R260 B.n46 B.n45 585
R261 B.n355 B.n46 585
R262 B.n353 B.n352 585
R263 B.n354 B.n353 585
R264 B.n405 B.n404 585
R265 B.n404 B.n403 585
R266 B.n187 B.n118 468.476
R267 B.n353 B.n51 468.476
R268 B.n189 B.n116 468.476
R269 B.n300 B.n49 468.476
R270 B.n131 B.t20 258.921
R271 B.n123 B.t23 258.921
R272 B.n56 B.t15 258.921
R273 B.n62 B.t12 258.921
R274 B.n301 B.n50 256.663
R275 B.n303 B.n50 256.663
R276 B.n309 B.n50 256.663
R277 B.n65 B.n50 256.663
R278 B.n315 B.n50 256.663
R279 B.n321 B.n50 256.663
R280 B.n323 B.n50 256.663
R281 B.n329 B.n50 256.663
R282 B.n331 B.n50 256.663
R283 B.n338 B.n50 256.663
R284 B.n340 B.n50 256.663
R285 B.n346 B.n50 256.663
R286 B.n348 B.n50 256.663
R287 B.n182 B.n117 256.663
R288 B.n120 B.n117 256.663
R289 B.n175 B.n117 256.663
R290 B.n168 B.n117 256.663
R291 B.n166 B.n117 256.663
R292 B.n160 B.n117 256.663
R293 B.n158 B.n117 256.663
R294 B.n152 B.n117 256.663
R295 B.n150 B.n117 256.663
R296 B.n144 B.n117 256.663
R297 B.n142 B.n117 256.663
R298 B.n136 B.n117 256.663
R299 B.n132 B.t19 239.333
R300 B.n124 B.t22 239.333
R301 B.n57 B.t16 239.333
R302 B.n63 B.t13 239.333
R303 B.n131 B.t17 224.483
R304 B.n123 B.t21 224.483
R305 B.n56 B.t14 224.483
R306 B.n62 B.t10 224.483
R307 B.n188 B.n117 222.81
R308 B.n354 B.n50 222.81
R309 B.n187 B.n112 163.367
R310 B.n195 B.n112 163.367
R311 B.n195 B.n110 163.367
R312 B.n199 B.n110 163.367
R313 B.n199 B.n104 163.367
R314 B.n207 B.n104 163.367
R315 B.n207 B.n102 163.367
R316 B.n211 B.n102 163.367
R317 B.n211 B.n96 163.367
R318 B.n220 B.n96 163.367
R319 B.n220 B.n94 163.367
R320 B.n224 B.n94 163.367
R321 B.n224 B.n89 163.367
R322 B.n231 B.n89 163.367
R323 B.n231 B.n87 163.367
R324 B.n235 B.n87 163.367
R325 B.n235 B.n81 163.367
R326 B.n244 B.n81 163.367
R327 B.n244 B.n79 163.367
R328 B.n248 B.n79 163.367
R329 B.n248 B.n74 163.367
R330 B.n257 B.n74 163.367
R331 B.n257 B.n72 163.367
R332 B.n261 B.n72 163.367
R333 B.n261 B.n2 163.367
R334 B.n404 B.n2 163.367
R335 B.n404 B.n3 163.367
R336 B.n400 B.n3 163.367
R337 B.n400 B.n9 163.367
R338 B.n396 B.n9 163.367
R339 B.n396 B.n11 163.367
R340 B.n392 B.n11 163.367
R341 B.n392 B.n15 163.367
R342 B.n388 B.n15 163.367
R343 B.n388 B.n17 163.367
R344 B.n384 B.n17 163.367
R345 B.n384 B.n23 163.367
R346 B.n380 B.n23 163.367
R347 B.n380 B.n25 163.367
R348 B.n377 B.n25 163.367
R349 B.n377 B.n29 163.367
R350 B.n373 B.n29 163.367
R351 B.n373 B.n31 163.367
R352 B.n369 B.n31 163.367
R353 B.n369 B.n37 163.367
R354 B.n365 B.n37 163.367
R355 B.n365 B.n39 163.367
R356 B.n361 B.n39 163.367
R357 B.n361 B.n44 163.367
R358 B.n357 B.n44 163.367
R359 B.n357 B.n46 163.367
R360 B.n353 B.n46 163.367
R361 B.n183 B.n181 163.367
R362 B.n181 B.n180 163.367
R363 B.n177 B.n176 163.367
R364 B.n174 B.n122 163.367
R365 B.n169 B.n167 163.367
R366 B.n165 B.n126 163.367
R367 B.n161 B.n159 163.367
R368 B.n157 B.n128 163.367
R369 B.n153 B.n151 163.367
R370 B.n149 B.n130 163.367
R371 B.n145 B.n143 163.367
R372 B.n141 B.n135 163.367
R373 B.n137 B.n116 163.367
R374 B.n189 B.n114 163.367
R375 B.n193 B.n114 163.367
R376 B.n193 B.n108 163.367
R377 B.n201 B.n108 163.367
R378 B.n201 B.n106 163.367
R379 B.n205 B.n106 163.367
R380 B.n205 B.n100 163.367
R381 B.n213 B.n100 163.367
R382 B.n213 B.n98 163.367
R383 B.n217 B.n98 163.367
R384 B.n217 B.n93 163.367
R385 B.n226 B.n93 163.367
R386 B.n226 B.n91 163.367
R387 B.n230 B.n91 163.367
R388 B.n230 B.n85 163.367
R389 B.n237 B.n85 163.367
R390 B.n237 B.n83 163.367
R391 B.n241 B.n83 163.367
R392 B.n241 B.n78 163.367
R393 B.n250 B.n78 163.367
R394 B.n250 B.n76 163.367
R395 B.n255 B.n76 163.367
R396 B.n255 B.n70 163.367
R397 B.n263 B.n70 163.367
R398 B.n264 B.n263 163.367
R399 B.n264 B.n5 163.367
R400 B.n6 B.n5 163.367
R401 B.n7 B.n6 163.367
R402 B.n269 B.n7 163.367
R403 B.n269 B.n12 163.367
R404 B.n13 B.n12 163.367
R405 B.n14 B.n13 163.367
R406 B.n274 B.n14 163.367
R407 B.n274 B.n19 163.367
R408 B.n20 B.n19 163.367
R409 B.n21 B.n20 163.367
R410 B.n279 B.n21 163.367
R411 B.n279 B.n26 163.367
R412 B.n27 B.n26 163.367
R413 B.n28 B.n27 163.367
R414 B.n284 B.n28 163.367
R415 B.n284 B.n33 163.367
R416 B.n34 B.n33 163.367
R417 B.n35 B.n34 163.367
R418 B.n289 B.n35 163.367
R419 B.n289 B.n40 163.367
R420 B.n41 B.n40 163.367
R421 B.n42 B.n41 163.367
R422 B.n294 B.n42 163.367
R423 B.n294 B.n47 163.367
R424 B.n48 B.n47 163.367
R425 B.n49 B.n48 163.367
R426 B.n349 B.n347 163.367
R427 B.n345 B.n53 163.367
R428 B.n341 B.n339 163.367
R429 B.n337 B.n55 163.367
R430 B.n332 B.n330 163.367
R431 B.n328 B.n59 163.367
R432 B.n324 B.n322 163.367
R433 B.n320 B.n61 163.367
R434 B.n316 B.n314 163.367
R435 B.n311 B.n310 163.367
R436 B.n308 B.n67 163.367
R437 B.n304 B.n302 163.367
R438 B.n188 B.n113 127.32
R439 B.n194 B.n113 127.32
R440 B.n194 B.n109 127.32
R441 B.n200 B.n109 127.32
R442 B.n206 B.n105 127.32
R443 B.n206 B.n101 127.32
R444 B.n212 B.n101 127.32
R445 B.n212 B.n97 127.32
R446 B.n219 B.n97 127.32
R447 B.n219 B.n218 127.32
R448 B.n225 B.n90 127.32
R449 B.t6 B.n90 127.32
R450 B.t6 B.n86 127.32
R451 B.n236 B.n86 127.32
R452 B.n243 B.n82 127.32
R453 B.n243 B.n242 127.32
R454 B.n249 B.n75 127.32
R455 B.n256 B.n75 127.32
R456 B.n262 B.n71 127.32
R457 B.n262 B.n4 127.32
R458 B.n403 B.n4 127.32
R459 B.n403 B.n402 127.32
R460 B.n402 B.n401 127.32
R461 B.n401 B.n8 127.32
R462 B.n395 B.n394 127.32
R463 B.n394 B.n393 127.32
R464 B.n387 B.n18 127.32
R465 B.n387 B.n386 127.32
R466 B.n385 B.n22 127.32
R467 B.t1 B.n22 127.32
R468 B.t1 B.n379 127.32
R469 B.n379 B.n378 127.32
R470 B.n372 B.n32 127.32
R471 B.n372 B.n371 127.32
R472 B.n371 B.n370 127.32
R473 B.n370 B.n36 127.32
R474 B.n364 B.n36 127.32
R475 B.n364 B.n363 127.32
R476 B.n362 B.n43 127.32
R477 B.n356 B.n43 127.32
R478 B.n356 B.n355 127.32
R479 B.n355 B.n354 127.32
R480 B.n225 B.t8 123.575
R481 B.n236 B.t3 123.575
R482 B.t4 B.n385 123.575
R483 B.n378 B.t0 123.575
R484 B.n242 B.t2 119.831
R485 B.n18 B.t5 119.831
R486 B.n256 B.t7 116.085
R487 B.n395 B.t9 116.085
R488 B.n200 B.t18 108.597
R489 B.t11 B.n362 108.597
R490 B.n182 B.n118 71.676
R491 B.n180 B.n120 71.676
R492 B.n176 B.n175 71.676
R493 B.n168 B.n122 71.676
R494 B.n167 B.n166 71.676
R495 B.n160 B.n126 71.676
R496 B.n159 B.n158 71.676
R497 B.n152 B.n128 71.676
R498 B.n151 B.n150 71.676
R499 B.n144 B.n130 71.676
R500 B.n143 B.n142 71.676
R501 B.n136 B.n135 71.676
R502 B.n348 B.n51 71.676
R503 B.n347 B.n346 71.676
R504 B.n340 B.n53 71.676
R505 B.n339 B.n338 71.676
R506 B.n331 B.n55 71.676
R507 B.n330 B.n329 71.676
R508 B.n323 B.n59 71.676
R509 B.n322 B.n321 71.676
R510 B.n315 B.n61 71.676
R511 B.n314 B.n65 71.676
R512 B.n310 B.n309 71.676
R513 B.n303 B.n67 71.676
R514 B.n302 B.n301 71.676
R515 B.n301 B.n300 71.676
R516 B.n304 B.n303 71.676
R517 B.n309 B.n308 71.676
R518 B.n311 B.n65 71.676
R519 B.n316 B.n315 71.676
R520 B.n321 B.n320 71.676
R521 B.n324 B.n323 71.676
R522 B.n329 B.n328 71.676
R523 B.n332 B.n331 71.676
R524 B.n338 B.n337 71.676
R525 B.n341 B.n340 71.676
R526 B.n346 B.n345 71.676
R527 B.n349 B.n348 71.676
R528 B.n183 B.n182 71.676
R529 B.n177 B.n120 71.676
R530 B.n175 B.n174 71.676
R531 B.n169 B.n168 71.676
R532 B.n166 B.n165 71.676
R533 B.n161 B.n160 71.676
R534 B.n158 B.n157 71.676
R535 B.n153 B.n152 71.676
R536 B.n150 B.n149 71.676
R537 B.n145 B.n144 71.676
R538 B.n142 B.n141 71.676
R539 B.n137 B.n136 71.676
R540 B.n133 B.n132 59.5399
R541 B.n171 B.n124 59.5399
R542 B.n335 B.n57 59.5399
R543 B.n64 B.n63 59.5399
R544 B.n352 B.n351 30.4395
R545 B.n299 B.n298 30.4395
R546 B.n190 B.n115 30.4395
R547 B.n186 B.n185 30.4395
R548 B.n132 B.n131 19.5884
R549 B.n124 B.n123 19.5884
R550 B.n57 B.n56 19.5884
R551 B.n63 B.n62 19.5884
R552 B.t18 B.n105 18.7239
R553 B.n363 B.t11 18.7239
R554 B B.n405 18.0485
R555 B.t7 B.n71 11.2345
R556 B.t9 B.n8 11.2345
R557 B.n351 B.n350 10.6151
R558 B.n350 B.n52 10.6151
R559 B.n344 B.n52 10.6151
R560 B.n344 B.n343 10.6151
R561 B.n343 B.n342 10.6151
R562 B.n342 B.n54 10.6151
R563 B.n336 B.n54 10.6151
R564 B.n334 B.n333 10.6151
R565 B.n333 B.n58 10.6151
R566 B.n327 B.n58 10.6151
R567 B.n327 B.n326 10.6151
R568 B.n326 B.n325 10.6151
R569 B.n325 B.n60 10.6151
R570 B.n319 B.n60 10.6151
R571 B.n319 B.n318 10.6151
R572 B.n318 B.n317 10.6151
R573 B.n313 B.n312 10.6151
R574 B.n312 B.n66 10.6151
R575 B.n307 B.n66 10.6151
R576 B.n307 B.n306 10.6151
R577 B.n306 B.n305 10.6151
R578 B.n305 B.n68 10.6151
R579 B.n299 B.n68 10.6151
R580 B.n191 B.n190 10.6151
R581 B.n192 B.n191 10.6151
R582 B.n192 B.n107 10.6151
R583 B.n202 B.n107 10.6151
R584 B.n203 B.n202 10.6151
R585 B.n204 B.n203 10.6151
R586 B.n204 B.n99 10.6151
R587 B.n214 B.n99 10.6151
R588 B.n215 B.n214 10.6151
R589 B.n216 B.n215 10.6151
R590 B.n216 B.n92 10.6151
R591 B.n227 B.n92 10.6151
R592 B.n228 B.n227 10.6151
R593 B.n229 B.n228 10.6151
R594 B.n229 B.n84 10.6151
R595 B.n238 B.n84 10.6151
R596 B.n239 B.n238 10.6151
R597 B.n240 B.n239 10.6151
R598 B.n240 B.n77 10.6151
R599 B.n251 B.n77 10.6151
R600 B.n252 B.n251 10.6151
R601 B.n254 B.n252 10.6151
R602 B.n254 B.n253 10.6151
R603 B.n253 B.n69 10.6151
R604 B.n265 B.n69 10.6151
R605 B.n266 B.n265 10.6151
R606 B.n267 B.n266 10.6151
R607 B.n268 B.n267 10.6151
R608 B.n270 B.n268 10.6151
R609 B.n271 B.n270 10.6151
R610 B.n272 B.n271 10.6151
R611 B.n273 B.n272 10.6151
R612 B.n275 B.n273 10.6151
R613 B.n276 B.n275 10.6151
R614 B.n277 B.n276 10.6151
R615 B.n278 B.n277 10.6151
R616 B.n280 B.n278 10.6151
R617 B.n281 B.n280 10.6151
R618 B.n282 B.n281 10.6151
R619 B.n283 B.n282 10.6151
R620 B.n285 B.n283 10.6151
R621 B.n286 B.n285 10.6151
R622 B.n287 B.n286 10.6151
R623 B.n288 B.n287 10.6151
R624 B.n290 B.n288 10.6151
R625 B.n291 B.n290 10.6151
R626 B.n292 B.n291 10.6151
R627 B.n293 B.n292 10.6151
R628 B.n295 B.n293 10.6151
R629 B.n296 B.n295 10.6151
R630 B.n297 B.n296 10.6151
R631 B.n298 B.n297 10.6151
R632 B.n185 B.n184 10.6151
R633 B.n184 B.n119 10.6151
R634 B.n179 B.n119 10.6151
R635 B.n179 B.n178 10.6151
R636 B.n178 B.n121 10.6151
R637 B.n173 B.n121 10.6151
R638 B.n173 B.n172 10.6151
R639 B.n170 B.n125 10.6151
R640 B.n164 B.n125 10.6151
R641 B.n164 B.n163 10.6151
R642 B.n163 B.n162 10.6151
R643 B.n162 B.n127 10.6151
R644 B.n156 B.n127 10.6151
R645 B.n156 B.n155 10.6151
R646 B.n155 B.n154 10.6151
R647 B.n154 B.n129 10.6151
R648 B.n148 B.n147 10.6151
R649 B.n147 B.n146 10.6151
R650 B.n146 B.n134 10.6151
R651 B.n140 B.n134 10.6151
R652 B.n140 B.n139 10.6151
R653 B.n139 B.n138 10.6151
R654 B.n138 B.n115 10.6151
R655 B.n186 B.n111 10.6151
R656 B.n196 B.n111 10.6151
R657 B.n197 B.n196 10.6151
R658 B.n198 B.n197 10.6151
R659 B.n198 B.n103 10.6151
R660 B.n208 B.n103 10.6151
R661 B.n209 B.n208 10.6151
R662 B.n210 B.n209 10.6151
R663 B.n210 B.n95 10.6151
R664 B.n221 B.n95 10.6151
R665 B.n222 B.n221 10.6151
R666 B.n223 B.n222 10.6151
R667 B.n223 B.n88 10.6151
R668 B.n232 B.n88 10.6151
R669 B.n233 B.n232 10.6151
R670 B.n234 B.n233 10.6151
R671 B.n234 B.n80 10.6151
R672 B.n245 B.n80 10.6151
R673 B.n246 B.n245 10.6151
R674 B.n247 B.n246 10.6151
R675 B.n247 B.n73 10.6151
R676 B.n258 B.n73 10.6151
R677 B.n259 B.n258 10.6151
R678 B.n260 B.n259 10.6151
R679 B.n260 B.n0 10.6151
R680 B.n399 B.n1 10.6151
R681 B.n399 B.n398 10.6151
R682 B.n398 B.n397 10.6151
R683 B.n397 B.n10 10.6151
R684 B.n391 B.n10 10.6151
R685 B.n391 B.n390 10.6151
R686 B.n390 B.n389 10.6151
R687 B.n389 B.n16 10.6151
R688 B.n383 B.n16 10.6151
R689 B.n383 B.n382 10.6151
R690 B.n382 B.n381 10.6151
R691 B.n381 B.n24 10.6151
R692 B.n376 B.n24 10.6151
R693 B.n376 B.n375 10.6151
R694 B.n375 B.n374 10.6151
R695 B.n374 B.n30 10.6151
R696 B.n368 B.n30 10.6151
R697 B.n368 B.n367 10.6151
R698 B.n367 B.n366 10.6151
R699 B.n366 B.n38 10.6151
R700 B.n360 B.n38 10.6151
R701 B.n360 B.n359 10.6151
R702 B.n359 B.n358 10.6151
R703 B.n358 B.n45 10.6151
R704 B.n352 B.n45 10.6151
R705 B.n336 B.n335 9.36635
R706 B.n313 B.n64 9.36635
R707 B.n172 B.n171 9.36635
R708 B.n148 B.n133 9.36635
R709 B.n249 B.t2 7.48986
R710 B.n393 B.t5 7.48986
R711 B.n218 B.t8 3.74518
R712 B.t3 B.n82 3.74518
R713 B.n386 B.t4 3.74518
R714 B.n32 B.t0 3.74518
R715 B.n405 B.n0 2.81026
R716 B.n405 B.n1 2.81026
R717 B.n335 B.n334 1.24928
R718 B.n317 B.n64 1.24928
R719 B.n171 B.n170 1.24928
R720 B.n133 B.n129 1.24928
R721 VN.n13 VN.n12 161.3
R722 VN.n27 VN.n26 161.3
R723 VN.n25 VN.n14 161.3
R724 VN.n24 VN.n23 161.3
R725 VN.n22 VN.n15 161.3
R726 VN.n21 VN.n20 161.3
R727 VN.n19 VN.n16 161.3
R728 VN.n11 VN.n0 161.3
R729 VN.n10 VN.n9 161.3
R730 VN.n8 VN.n1 161.3
R731 VN.n7 VN.n6 161.3
R732 VN.n5 VN.n2 161.3
R733 VN.n3 VN.t3 101.338
R734 VN.n17 VN.t5 101.338
R735 VN.n4 VN.t2 79.7431
R736 VN.n6 VN.t7 79.7431
R737 VN.n10 VN.t6 79.7431
R738 VN.n12 VN.t8 79.7431
R739 VN.n18 VN.t1 79.7431
R740 VN.n20 VN.t0 79.7431
R741 VN.n24 VN.t9 79.7431
R742 VN.n26 VN.t4 79.7431
R743 VN.n17 VN.n16 44.8545
R744 VN.n3 VN.n2 44.8545
R745 VN VN.n27 34.385
R746 VN.n12 VN.n11 26.2914
R747 VN.n26 VN.n25 26.2914
R748 VN.n5 VN.n4 24.8308
R749 VN.n10 VN.n1 24.8308
R750 VN.n19 VN.n18 24.8308
R751 VN.n24 VN.n15 24.8308
R752 VN.n6 VN.n5 23.3702
R753 VN.n6 VN.n1 23.3702
R754 VN.n20 VN.n19 23.3702
R755 VN.n20 VN.n15 23.3702
R756 VN.n11 VN.n10 21.9096
R757 VN.n25 VN.n24 21.9096
R758 VN.n4 VN.n3 20.3348
R759 VN.n18 VN.n17 20.3348
R760 VN.n27 VN.n14 0.189894
R761 VN.n23 VN.n14 0.189894
R762 VN.n23 VN.n22 0.189894
R763 VN.n22 VN.n21 0.189894
R764 VN.n21 VN.n16 0.189894
R765 VN.n7 VN.n2 0.189894
R766 VN.n8 VN.n7 0.189894
R767 VN.n9 VN.n8 0.189894
R768 VN.n9 VN.n0 0.189894
R769 VN.n13 VN.n0 0.189894
R770 VN VN.n13 0.0516364
R771 VTAIL.n17 VTAIL.t12 250.185
R772 VTAIL.n2 VTAIL.t7 250.185
R773 VTAIL.n16 VTAIL.t0 250.185
R774 VTAIL.n11 VTAIL.t10 250.185
R775 VTAIL.n19 VTAIL.n18 217.185
R776 VTAIL.n1 VTAIL.n0 217.185
R777 VTAIL.n4 VTAIL.n3 217.185
R778 VTAIL.n6 VTAIL.n5 217.185
R779 VTAIL.n15 VTAIL.n14 217.185
R780 VTAIL.n13 VTAIL.n12 217.185
R781 VTAIL.n10 VTAIL.n9 217.185
R782 VTAIL.n8 VTAIL.n7 217.185
R783 VTAIL.n18 VTAIL.t17 33.0005
R784 VTAIL.n18 VTAIL.t14 33.0005
R785 VTAIL.n0 VTAIL.t11 33.0005
R786 VTAIL.n0 VTAIL.t13 33.0005
R787 VTAIL.n3 VTAIL.t3 33.0005
R788 VTAIL.n3 VTAIL.t2 33.0005
R789 VTAIL.n5 VTAIL.t8 33.0005
R790 VTAIL.n5 VTAIL.t6 33.0005
R791 VTAIL.n14 VTAIL.t4 33.0005
R792 VTAIL.n14 VTAIL.t1 33.0005
R793 VTAIL.n12 VTAIL.t9 33.0005
R794 VTAIL.n12 VTAIL.t5 33.0005
R795 VTAIL.n9 VTAIL.t19 33.0005
R796 VTAIL.n9 VTAIL.t18 33.0005
R797 VTAIL.n7 VTAIL.t16 33.0005
R798 VTAIL.n7 VTAIL.t15 33.0005
R799 VTAIL.n8 VTAIL.n6 14.6255
R800 VTAIL.n17 VTAIL.n16 13.7548
R801 VTAIL.n13 VTAIL.n11 0.905672
R802 VTAIL.n2 VTAIL.n1 0.905672
R803 VTAIL.n10 VTAIL.n8 0.87119
R804 VTAIL.n11 VTAIL.n10 0.87119
R805 VTAIL.n15 VTAIL.n13 0.87119
R806 VTAIL.n16 VTAIL.n15 0.87119
R807 VTAIL.n6 VTAIL.n4 0.87119
R808 VTAIL.n4 VTAIL.n2 0.87119
R809 VTAIL.n19 VTAIL.n17 0.87119
R810 VTAIL VTAIL.n1 0.711707
R811 VTAIL VTAIL.n19 0.159983
R812 VDD2.n1 VDD2.t6 267.735
R813 VDD2.n4 VDD2.t5 266.865
R814 VDD2.n3 VDD2.n2 234.462
R815 VDD2 VDD2.n7 234.458
R816 VDD2.n6 VDD2.n5 233.864
R817 VDD2.n1 VDD2.n0 233.864
R818 VDD2.n7 VDD2.t8 33.0005
R819 VDD2.n7 VDD2.t4 33.0005
R820 VDD2.n5 VDD2.t0 33.0005
R821 VDD2.n5 VDD2.t9 33.0005
R822 VDD2.n2 VDD2.t3 33.0005
R823 VDD2.n2 VDD2.t1 33.0005
R824 VDD2.n0 VDD2.t7 33.0005
R825 VDD2.n0 VDD2.t2 33.0005
R826 VDD2.n4 VDD2.n3 28.3683
R827 VDD2.n6 VDD2.n4 0.87119
R828 VDD2 VDD2.n6 0.276362
R829 VDD2.n3 VDD2.n1 0.162826
R830 VP.n31 VP.n30 161.3
R831 VP.n10 VP.n9 161.3
R832 VP.n11 VP.n6 161.3
R833 VP.n13 VP.n12 161.3
R834 VP.n14 VP.n5 161.3
R835 VP.n15 VP.n4 161.3
R836 VP.n17 VP.n16 161.3
R837 VP.n29 VP.n0 161.3
R838 VP.n28 VP.n27 161.3
R839 VP.n26 VP.n1 161.3
R840 VP.n25 VP.n24 161.3
R841 VP.n23 VP.n2 161.3
R842 VP.n22 VP.n21 161.3
R843 VP.n20 VP.n3 161.3
R844 VP.n19 VP.n18 161.3
R845 VP.n7 VP.t3 101.338
R846 VP.n18 VP.t1 79.7431
R847 VP.n22 VP.t9 79.7431
R848 VP.n24 VP.t8 79.7431
R849 VP.n28 VP.t7 79.7431
R850 VP.n30 VP.t6 79.7431
R851 VP.n16 VP.t2 79.7431
R852 VP.n14 VP.t4 79.7431
R853 VP.n6 VP.t5 79.7431
R854 VP.n8 VP.t0 79.7431
R855 VP.n10 VP.n7 44.8545
R856 VP.n19 VP.n17 34.0043
R857 VP.n18 VP.n3 26.2914
R858 VP.n30 VP.n29 26.2914
R859 VP.n16 VP.n15 26.2914
R860 VP.n23 VP.n22 24.8308
R861 VP.n28 VP.n1 24.8308
R862 VP.n14 VP.n13 24.8308
R863 VP.n9 VP.n8 24.8308
R864 VP.n24 VP.n23 23.3702
R865 VP.n24 VP.n1 23.3702
R866 VP.n13 VP.n6 23.3702
R867 VP.n9 VP.n6 23.3702
R868 VP.n22 VP.n3 21.9096
R869 VP.n29 VP.n28 21.9096
R870 VP.n15 VP.n14 21.9096
R871 VP.n8 VP.n7 20.3348
R872 VP.n11 VP.n10 0.189894
R873 VP.n12 VP.n11 0.189894
R874 VP.n12 VP.n5 0.189894
R875 VP.n5 VP.n4 0.189894
R876 VP.n17 VP.n4 0.189894
R877 VP.n20 VP.n19 0.189894
R878 VP.n21 VP.n20 0.189894
R879 VP.n21 VP.n2 0.189894
R880 VP.n25 VP.n2 0.189894
R881 VP.n26 VP.n25 0.189894
R882 VP.n27 VP.n26 0.189894
R883 VP.n27 VP.n0 0.189894
R884 VP.n31 VP.n0 0.189894
R885 VP VP.n31 0.0516364
R886 VDD1.n1 VDD1.t6 267.735
R887 VDD1.n3 VDD1.t8 267.735
R888 VDD1.n5 VDD1.n4 234.462
R889 VDD1.n7 VDD1.n6 233.864
R890 VDD1.n1 VDD1.n0 233.864
R891 VDD1.n3 VDD1.n2 233.864
R892 VDD1.n6 VDD1.t5 33.0005
R893 VDD1.n6 VDD1.t7 33.0005
R894 VDD1.n0 VDD1.t9 33.0005
R895 VDD1.n0 VDD1.t4 33.0005
R896 VDD1.n4 VDD1.t2 33.0005
R897 VDD1.n4 VDD1.t3 33.0005
R898 VDD1.n2 VDD1.t0 33.0005
R899 VDD1.n2 VDD1.t1 33.0005
R900 VDD1.n7 VDD1.n5 29.3867
R901 VDD1 VDD1.n7 0.595328
R902 VDD1 VDD1.n1 0.276362
R903 VDD1.n5 VDD1.n3 0.162826
C0 VDD2 VDD1 0.953768f
C1 VDD2 VN 0.750587f
C2 VDD1 VN 0.156801f
C3 VP VTAIL 1.25434f
C4 VDD2 VP 0.346617f
C5 VDD1 VP 0.938035f
C6 VN VP 3.47268f
C7 VDD2 VTAIL 3.12619f
C8 VDD1 VTAIL 3.0858f
C9 VN VTAIL 1.2402f
C10 VDD2 B 2.735265f
C11 VDD1 B 2.810792f
C12 VTAIL B 2.047037f
C13 VN B 7.467394f
C14 VP B 6.427934f
C15 VDD1.t6 B 0.050538f
C16 VDD1.t9 B 0.010549f
C17 VDD1.t4 B 0.010549f
C18 VDD1.n0 B 0.026917f
C19 VDD1.n1 B 0.270553f
C20 VDD1.t8 B 0.050538f
C21 VDD1.t0 B 0.010549f
C22 VDD1.t1 B 0.010549f
C23 VDD1.n2 B 0.026917f
C24 VDD1.n3 B 0.265591f
C25 VDD1.t2 B 0.010549f
C26 VDD1.t3 B 0.010549f
C27 VDD1.n4 B 0.027353f
C28 VDD1.n5 B 1.03539f
C29 VDD1.t5 B 0.010549f
C30 VDD1.t7 B 0.010549f
C31 VDD1.n6 B 0.026917f
C32 VDD1.n7 B 1.17247f
C33 VP.n0 B 0.031425f
C34 VP.n1 B 0.007131f
C35 VP.n2 B 0.031425f
C36 VP.n3 B 0.007131f
C37 VP.n4 B 0.031425f
C38 VP.t2 B 0.048906f
C39 VP.t4 B 0.048906f
C40 VP.n5 B 0.031425f
C41 VP.t5 B 0.048906f
C42 VP.n6 B 0.065026f
C43 VP.t3 B 0.062636f
C44 VP.n7 B 0.053797f
C45 VP.t0 B 0.048906f
C46 VP.n8 B 0.067569f
C47 VP.n9 B 0.007131f
C48 VP.n10 B 0.129334f
C49 VP.n11 B 0.031425f
C50 VP.n12 B 0.031425f
C51 VP.n13 B 0.007131f
C52 VP.n14 B 0.065026f
C53 VP.n15 B 0.007131f
C54 VP.n16 B 0.062313f
C55 VP.n17 B 0.885022f
C56 VP.t1 B 0.048906f
C57 VP.n18 B 0.062313f
C58 VP.n19 B 0.918146f
C59 VP.n20 B 0.031425f
C60 VP.n21 B 0.031425f
C61 VP.t9 B 0.048906f
C62 VP.n22 B 0.065026f
C63 VP.n23 B 0.007131f
C64 VP.t8 B 0.048906f
C65 VP.n24 B 0.065026f
C66 VP.n25 B 0.031425f
C67 VP.n26 B 0.031425f
C68 VP.n27 B 0.031425f
C69 VP.t7 B 0.048906f
C70 VP.n28 B 0.065026f
C71 VP.n29 B 0.007131f
C72 VP.t6 B 0.048906f
C73 VP.n30 B 0.062313f
C74 VP.n31 B 0.024353f
C75 VDD2.t6 B 0.051914f
C76 VDD2.t7 B 0.010837f
C77 VDD2.t2 B 0.010837f
C78 VDD2.n0 B 0.02765f
C79 VDD2.n1 B 0.272823f
C80 VDD2.t3 B 0.010837f
C81 VDD2.t1 B 0.010837f
C82 VDD2.n2 B 0.028098f
C83 VDD2.n3 B 0.999003f
C84 VDD2.t5 B 0.05147f
C85 VDD2.n4 B 1.14649f
C86 VDD2.t0 B 0.010837f
C87 VDD2.t9 B 0.010837f
C88 VDD2.n5 B 0.02765f
C89 VDD2.n6 B 0.14187f
C90 VDD2.t8 B 0.010837f
C91 VDD2.t4 B 0.010837f
C92 VDD2.n7 B 0.028093f
C93 VTAIL.t11 B 0.016749f
C94 VTAIL.t13 B 0.016749f
C95 VTAIL.n0 B 0.036436f
C96 VTAIL.n1 B 0.231042f
C97 VTAIL.t7 B 0.073493f
C98 VTAIL.n2 B 0.257817f
C99 VTAIL.t3 B 0.016749f
C100 VTAIL.t2 B 0.016749f
C101 VTAIL.n3 B 0.036436f
C102 VTAIL.n4 B 0.24527f
C103 VTAIL.t8 B 0.016749f
C104 VTAIL.t6 B 0.016749f
C105 VTAIL.n5 B 0.036436f
C106 VTAIL.n6 B 0.883105f
C107 VTAIL.t16 B 0.016749f
C108 VTAIL.t15 B 0.016749f
C109 VTAIL.n7 B 0.036436f
C110 VTAIL.n8 B 0.883105f
C111 VTAIL.t19 B 0.016749f
C112 VTAIL.t18 B 0.016749f
C113 VTAIL.n9 B 0.036436f
C114 VTAIL.n10 B 0.24527f
C115 VTAIL.t10 B 0.073493f
C116 VTAIL.n11 B 0.257817f
C117 VTAIL.t9 B 0.016749f
C118 VTAIL.t5 B 0.016749f
C119 VTAIL.n12 B 0.036436f
C120 VTAIL.n13 B 0.249195f
C121 VTAIL.t4 B 0.016749f
C122 VTAIL.t1 B 0.016749f
C123 VTAIL.n14 B 0.036436f
C124 VTAIL.n15 B 0.24527f
C125 VTAIL.t0 B 0.073493f
C126 VTAIL.n16 B 0.79262f
C127 VTAIL.t12 B 0.073493f
C128 VTAIL.n17 B 0.79262f
C129 VTAIL.t17 B 0.016749f
C130 VTAIL.t14 B 0.016749f
C131 VTAIL.n18 B 0.036436f
C132 VTAIL.n19 B 0.164316f
C133 VN.n0 B 0.031033f
C134 VN.n1 B 0.007042f
C135 VN.n2 B 0.127722f
C136 VN.t3 B 0.061856f
C137 VN.n3 B 0.053127f
C138 VN.t2 B 0.048297f
C139 VN.n4 B 0.066727f
C140 VN.n5 B 0.007042f
C141 VN.t7 B 0.048297f
C142 VN.n6 B 0.064215f
C143 VN.n7 B 0.031033f
C144 VN.n8 B 0.031033f
C145 VN.n9 B 0.031033f
C146 VN.t6 B 0.048297f
C147 VN.n10 B 0.064215f
C148 VN.n11 B 0.007042f
C149 VN.t8 B 0.048297f
C150 VN.n12 B 0.061537f
C151 VN.n13 B 0.024049f
C152 VN.n14 B 0.031033f
C153 VN.n15 B 0.007042f
C154 VN.t9 B 0.048297f
C155 VN.n16 B 0.127722f
C156 VN.t5 B 0.061856f
C157 VN.n17 B 0.053127f
C158 VN.t1 B 0.048297f
C159 VN.n18 B 0.066727f
C160 VN.n19 B 0.007042f
C161 VN.t0 B 0.048297f
C162 VN.n20 B 0.064215f
C163 VN.n21 B 0.031033f
C164 VN.n22 B 0.031033f
C165 VN.n23 B 0.031033f
C166 VN.n24 B 0.064215f
C167 VN.n25 B 0.007042f
C168 VN.t4 B 0.048297f
C169 VN.n26 B 0.061537f
C170 VN.n27 B 0.894663f
.ends

