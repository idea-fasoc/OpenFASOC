* NGSPICE file created from diff_pair_sample_0764.ext - technology: sky130A

.subckt diff_pair_sample_0764 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=1.48335 pd=9.32 as=3.5061 ps=18.76 w=8.99 l=2.54
X1 VTAIL.t6 VP.t1 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=3.5061 pd=18.76 as=1.48335 ps=9.32 w=8.99 l=2.54
X2 VDD1.t1 VP.t2 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=1.48335 pd=9.32 as=3.5061 ps=18.76 w=8.99 l=2.54
X3 VDD2.t3 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.48335 pd=9.32 as=3.5061 ps=18.76 w=8.99 l=2.54
X4 VTAIL.t3 VN.t1 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=3.5061 pd=18.76 as=1.48335 ps=9.32 w=8.99 l=2.54
X5 VTAIL.t7 VP.t3 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.5061 pd=18.76 as=1.48335 ps=9.32 w=8.99 l=2.54
X6 VTAIL.t0 VN.t2 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=3.5061 pd=18.76 as=1.48335 ps=9.32 w=8.99 l=2.54
X7 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=3.5061 pd=18.76 as=0 ps=0 w=8.99 l=2.54
X8 VDD2.t0 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.48335 pd=9.32 as=3.5061 ps=18.76 w=8.99 l=2.54
X9 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=3.5061 pd=18.76 as=0 ps=0 w=8.99 l=2.54
X10 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=3.5061 pd=18.76 as=0 ps=0 w=8.99 l=2.54
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.5061 pd=18.76 as=0 ps=0 w=8.99 l=2.54
R0 VP.n14 VP.n0 161.3
R1 VP.n13 VP.n12 161.3
R2 VP.n11 VP.n1 161.3
R3 VP.n10 VP.n9 161.3
R4 VP.n8 VP.n2 161.3
R5 VP.n7 VP.n6 161.3
R6 VP.n4 VP.t3 121.041
R7 VP.n4 VP.t0 120.276
R8 VP.n5 VP.n3 101.704
R9 VP.n16 VP.n15 101.704
R10 VP.n3 VP.t1 85.2993
R11 VP.n15 VP.t2 85.2993
R12 VP.n9 VP.n1 56.5193
R13 VP.n5 VP.n4 48.2728
R14 VP.n8 VP.n7 24.4675
R15 VP.n9 VP.n8 24.4675
R16 VP.n13 VP.n1 24.4675
R17 VP.n14 VP.n13 24.4675
R18 VP.n7 VP.n3 9.05329
R19 VP.n15 VP.n14 9.05329
R20 VP.n6 VP.n5 0.278367
R21 VP.n16 VP.n0 0.278367
R22 VP.n6 VP.n2 0.189894
R23 VP.n10 VP.n2 0.189894
R24 VP.n11 VP.n10 0.189894
R25 VP.n12 VP.n11 0.189894
R26 VP.n12 VP.n0 0.189894
R27 VP VP.n16 0.153454
R28 VTAIL.n5 VTAIL.t7 50.8673
R29 VTAIL.n4 VTAIL.t2 50.8673
R30 VTAIL.n3 VTAIL.t3 50.8673
R31 VTAIL.n7 VTAIL.t1 50.8671
R32 VTAIL.n0 VTAIL.t0 50.8671
R33 VTAIL.n1 VTAIL.t4 50.8671
R34 VTAIL.n2 VTAIL.t6 50.8671
R35 VTAIL.n6 VTAIL.t5 50.8671
R36 VTAIL.n7 VTAIL.n6 22.591
R37 VTAIL.n3 VTAIL.n2 22.591
R38 VTAIL.n4 VTAIL.n3 2.47464
R39 VTAIL.n6 VTAIL.n5 2.47464
R40 VTAIL.n2 VTAIL.n1 2.47464
R41 VTAIL VTAIL.n0 1.29576
R42 VTAIL VTAIL.n7 1.17938
R43 VTAIL.n5 VTAIL.n4 0.470328
R44 VTAIL.n1 VTAIL.n0 0.470328
R45 VDD1 VDD1.n1 104.755
R46 VDD1 VDD1.n0 65.4017
R47 VDD1.n0 VDD1.t0 2.20295
R48 VDD1.n0 VDD1.t3 2.20295
R49 VDD1.n1 VDD1.t2 2.20295
R50 VDD1.n1 VDD1.t1 2.20295
R51 B.n656 B.n655 585
R52 B.n657 B.n656 585
R53 B.n254 B.n101 585
R54 B.n253 B.n252 585
R55 B.n251 B.n250 585
R56 B.n249 B.n248 585
R57 B.n247 B.n246 585
R58 B.n245 B.n244 585
R59 B.n243 B.n242 585
R60 B.n241 B.n240 585
R61 B.n239 B.n238 585
R62 B.n237 B.n236 585
R63 B.n235 B.n234 585
R64 B.n233 B.n232 585
R65 B.n231 B.n230 585
R66 B.n229 B.n228 585
R67 B.n227 B.n226 585
R68 B.n225 B.n224 585
R69 B.n223 B.n222 585
R70 B.n221 B.n220 585
R71 B.n219 B.n218 585
R72 B.n217 B.n216 585
R73 B.n215 B.n214 585
R74 B.n213 B.n212 585
R75 B.n211 B.n210 585
R76 B.n209 B.n208 585
R77 B.n207 B.n206 585
R78 B.n205 B.n204 585
R79 B.n203 B.n202 585
R80 B.n201 B.n200 585
R81 B.n199 B.n198 585
R82 B.n197 B.n196 585
R83 B.n195 B.n194 585
R84 B.n193 B.n192 585
R85 B.n191 B.n190 585
R86 B.n189 B.n188 585
R87 B.n187 B.n186 585
R88 B.n185 B.n184 585
R89 B.n183 B.n182 585
R90 B.n181 B.n180 585
R91 B.n179 B.n178 585
R92 B.n177 B.n176 585
R93 B.n175 B.n174 585
R94 B.n172 B.n171 585
R95 B.n170 B.n169 585
R96 B.n168 B.n167 585
R97 B.n166 B.n165 585
R98 B.n164 B.n163 585
R99 B.n162 B.n161 585
R100 B.n160 B.n159 585
R101 B.n158 B.n157 585
R102 B.n156 B.n155 585
R103 B.n154 B.n153 585
R104 B.n152 B.n151 585
R105 B.n150 B.n149 585
R106 B.n148 B.n147 585
R107 B.n146 B.n145 585
R108 B.n144 B.n143 585
R109 B.n142 B.n141 585
R110 B.n140 B.n139 585
R111 B.n138 B.n137 585
R112 B.n136 B.n135 585
R113 B.n134 B.n133 585
R114 B.n132 B.n131 585
R115 B.n130 B.n129 585
R116 B.n128 B.n127 585
R117 B.n126 B.n125 585
R118 B.n124 B.n123 585
R119 B.n122 B.n121 585
R120 B.n120 B.n119 585
R121 B.n118 B.n117 585
R122 B.n116 B.n115 585
R123 B.n114 B.n113 585
R124 B.n112 B.n111 585
R125 B.n110 B.n109 585
R126 B.n108 B.n107 585
R127 B.n654 B.n63 585
R128 B.n658 B.n63 585
R129 B.n653 B.n62 585
R130 B.n659 B.n62 585
R131 B.n652 B.n651 585
R132 B.n651 B.n58 585
R133 B.n650 B.n57 585
R134 B.n665 B.n57 585
R135 B.n649 B.n56 585
R136 B.n666 B.n56 585
R137 B.n648 B.n55 585
R138 B.n667 B.n55 585
R139 B.n647 B.n646 585
R140 B.n646 B.n51 585
R141 B.n645 B.n50 585
R142 B.n673 B.n50 585
R143 B.n644 B.n49 585
R144 B.n674 B.n49 585
R145 B.n643 B.n48 585
R146 B.n675 B.n48 585
R147 B.n642 B.n641 585
R148 B.n641 B.n44 585
R149 B.n640 B.n43 585
R150 B.n681 B.n43 585
R151 B.n639 B.n42 585
R152 B.n682 B.n42 585
R153 B.n638 B.n41 585
R154 B.n683 B.n41 585
R155 B.n637 B.n636 585
R156 B.n636 B.n37 585
R157 B.n635 B.n36 585
R158 B.n689 B.n36 585
R159 B.n634 B.n35 585
R160 B.n690 B.n35 585
R161 B.n633 B.n34 585
R162 B.n691 B.n34 585
R163 B.n632 B.n631 585
R164 B.n631 B.n30 585
R165 B.n630 B.n29 585
R166 B.n697 B.n29 585
R167 B.n629 B.n28 585
R168 B.n698 B.n28 585
R169 B.n628 B.n27 585
R170 B.n699 B.n27 585
R171 B.n627 B.n626 585
R172 B.n626 B.n23 585
R173 B.n625 B.n22 585
R174 B.n705 B.n22 585
R175 B.n624 B.n21 585
R176 B.n706 B.n21 585
R177 B.n623 B.n20 585
R178 B.n707 B.n20 585
R179 B.n622 B.n621 585
R180 B.n621 B.n16 585
R181 B.n620 B.n15 585
R182 B.n713 B.n15 585
R183 B.n619 B.n14 585
R184 B.n714 B.n14 585
R185 B.n618 B.n13 585
R186 B.n715 B.n13 585
R187 B.n617 B.n616 585
R188 B.n616 B.n12 585
R189 B.n615 B.n614 585
R190 B.n615 B.n8 585
R191 B.n613 B.n7 585
R192 B.n722 B.n7 585
R193 B.n612 B.n6 585
R194 B.n723 B.n6 585
R195 B.n611 B.n5 585
R196 B.n724 B.n5 585
R197 B.n610 B.n609 585
R198 B.n609 B.n4 585
R199 B.n608 B.n255 585
R200 B.n608 B.n607 585
R201 B.n598 B.n256 585
R202 B.n257 B.n256 585
R203 B.n600 B.n599 585
R204 B.n601 B.n600 585
R205 B.n597 B.n262 585
R206 B.n262 B.n261 585
R207 B.n596 B.n595 585
R208 B.n595 B.n594 585
R209 B.n264 B.n263 585
R210 B.n265 B.n264 585
R211 B.n587 B.n586 585
R212 B.n588 B.n587 585
R213 B.n585 B.n270 585
R214 B.n270 B.n269 585
R215 B.n584 B.n583 585
R216 B.n583 B.n582 585
R217 B.n272 B.n271 585
R218 B.n273 B.n272 585
R219 B.n575 B.n574 585
R220 B.n576 B.n575 585
R221 B.n573 B.n278 585
R222 B.n278 B.n277 585
R223 B.n572 B.n571 585
R224 B.n571 B.n570 585
R225 B.n280 B.n279 585
R226 B.n281 B.n280 585
R227 B.n563 B.n562 585
R228 B.n564 B.n563 585
R229 B.n561 B.n286 585
R230 B.n286 B.n285 585
R231 B.n560 B.n559 585
R232 B.n559 B.n558 585
R233 B.n288 B.n287 585
R234 B.n289 B.n288 585
R235 B.n551 B.n550 585
R236 B.n552 B.n551 585
R237 B.n549 B.n294 585
R238 B.n294 B.n293 585
R239 B.n548 B.n547 585
R240 B.n547 B.n546 585
R241 B.n296 B.n295 585
R242 B.n297 B.n296 585
R243 B.n539 B.n538 585
R244 B.n540 B.n539 585
R245 B.n537 B.n302 585
R246 B.n302 B.n301 585
R247 B.n536 B.n535 585
R248 B.n535 B.n534 585
R249 B.n304 B.n303 585
R250 B.n305 B.n304 585
R251 B.n527 B.n526 585
R252 B.n528 B.n527 585
R253 B.n525 B.n310 585
R254 B.n310 B.n309 585
R255 B.n524 B.n523 585
R256 B.n523 B.n522 585
R257 B.n312 B.n311 585
R258 B.n313 B.n312 585
R259 B.n515 B.n514 585
R260 B.n516 B.n515 585
R261 B.n513 B.n318 585
R262 B.n318 B.n317 585
R263 B.n507 B.n506 585
R264 B.n505 B.n357 585
R265 B.n504 B.n356 585
R266 B.n509 B.n356 585
R267 B.n503 B.n502 585
R268 B.n501 B.n500 585
R269 B.n499 B.n498 585
R270 B.n497 B.n496 585
R271 B.n495 B.n494 585
R272 B.n493 B.n492 585
R273 B.n491 B.n490 585
R274 B.n489 B.n488 585
R275 B.n487 B.n486 585
R276 B.n485 B.n484 585
R277 B.n483 B.n482 585
R278 B.n481 B.n480 585
R279 B.n479 B.n478 585
R280 B.n477 B.n476 585
R281 B.n475 B.n474 585
R282 B.n473 B.n472 585
R283 B.n471 B.n470 585
R284 B.n469 B.n468 585
R285 B.n467 B.n466 585
R286 B.n465 B.n464 585
R287 B.n463 B.n462 585
R288 B.n461 B.n460 585
R289 B.n459 B.n458 585
R290 B.n457 B.n456 585
R291 B.n455 B.n454 585
R292 B.n453 B.n452 585
R293 B.n451 B.n450 585
R294 B.n449 B.n448 585
R295 B.n447 B.n446 585
R296 B.n445 B.n444 585
R297 B.n443 B.n442 585
R298 B.n441 B.n440 585
R299 B.n439 B.n438 585
R300 B.n437 B.n436 585
R301 B.n435 B.n434 585
R302 B.n433 B.n432 585
R303 B.n431 B.n430 585
R304 B.n429 B.n428 585
R305 B.n427 B.n426 585
R306 B.n424 B.n423 585
R307 B.n422 B.n421 585
R308 B.n420 B.n419 585
R309 B.n418 B.n417 585
R310 B.n416 B.n415 585
R311 B.n414 B.n413 585
R312 B.n412 B.n411 585
R313 B.n410 B.n409 585
R314 B.n408 B.n407 585
R315 B.n406 B.n405 585
R316 B.n404 B.n403 585
R317 B.n402 B.n401 585
R318 B.n400 B.n399 585
R319 B.n398 B.n397 585
R320 B.n396 B.n395 585
R321 B.n394 B.n393 585
R322 B.n392 B.n391 585
R323 B.n390 B.n389 585
R324 B.n388 B.n387 585
R325 B.n386 B.n385 585
R326 B.n384 B.n383 585
R327 B.n382 B.n381 585
R328 B.n380 B.n379 585
R329 B.n378 B.n377 585
R330 B.n376 B.n375 585
R331 B.n374 B.n373 585
R332 B.n372 B.n371 585
R333 B.n370 B.n369 585
R334 B.n368 B.n367 585
R335 B.n366 B.n365 585
R336 B.n364 B.n363 585
R337 B.n320 B.n319 585
R338 B.n512 B.n511 585
R339 B.n316 B.n315 585
R340 B.n317 B.n316 585
R341 B.n518 B.n517 585
R342 B.n517 B.n516 585
R343 B.n519 B.n314 585
R344 B.n314 B.n313 585
R345 B.n521 B.n520 585
R346 B.n522 B.n521 585
R347 B.n308 B.n307 585
R348 B.n309 B.n308 585
R349 B.n530 B.n529 585
R350 B.n529 B.n528 585
R351 B.n531 B.n306 585
R352 B.n306 B.n305 585
R353 B.n533 B.n532 585
R354 B.n534 B.n533 585
R355 B.n300 B.n299 585
R356 B.n301 B.n300 585
R357 B.n542 B.n541 585
R358 B.n541 B.n540 585
R359 B.n543 B.n298 585
R360 B.n298 B.n297 585
R361 B.n545 B.n544 585
R362 B.n546 B.n545 585
R363 B.n292 B.n291 585
R364 B.n293 B.n292 585
R365 B.n554 B.n553 585
R366 B.n553 B.n552 585
R367 B.n555 B.n290 585
R368 B.n290 B.n289 585
R369 B.n557 B.n556 585
R370 B.n558 B.n557 585
R371 B.n284 B.n283 585
R372 B.n285 B.n284 585
R373 B.n566 B.n565 585
R374 B.n565 B.n564 585
R375 B.n567 B.n282 585
R376 B.n282 B.n281 585
R377 B.n569 B.n568 585
R378 B.n570 B.n569 585
R379 B.n276 B.n275 585
R380 B.n277 B.n276 585
R381 B.n578 B.n577 585
R382 B.n577 B.n576 585
R383 B.n579 B.n274 585
R384 B.n274 B.n273 585
R385 B.n581 B.n580 585
R386 B.n582 B.n581 585
R387 B.n268 B.n267 585
R388 B.n269 B.n268 585
R389 B.n590 B.n589 585
R390 B.n589 B.n588 585
R391 B.n591 B.n266 585
R392 B.n266 B.n265 585
R393 B.n593 B.n592 585
R394 B.n594 B.n593 585
R395 B.n260 B.n259 585
R396 B.n261 B.n260 585
R397 B.n603 B.n602 585
R398 B.n602 B.n601 585
R399 B.n604 B.n258 585
R400 B.n258 B.n257 585
R401 B.n606 B.n605 585
R402 B.n607 B.n606 585
R403 B.n3 B.n0 585
R404 B.n4 B.n3 585
R405 B.n721 B.n1 585
R406 B.n722 B.n721 585
R407 B.n720 B.n719 585
R408 B.n720 B.n8 585
R409 B.n718 B.n9 585
R410 B.n12 B.n9 585
R411 B.n717 B.n716 585
R412 B.n716 B.n715 585
R413 B.n11 B.n10 585
R414 B.n714 B.n11 585
R415 B.n712 B.n711 585
R416 B.n713 B.n712 585
R417 B.n710 B.n17 585
R418 B.n17 B.n16 585
R419 B.n709 B.n708 585
R420 B.n708 B.n707 585
R421 B.n19 B.n18 585
R422 B.n706 B.n19 585
R423 B.n704 B.n703 585
R424 B.n705 B.n704 585
R425 B.n702 B.n24 585
R426 B.n24 B.n23 585
R427 B.n701 B.n700 585
R428 B.n700 B.n699 585
R429 B.n26 B.n25 585
R430 B.n698 B.n26 585
R431 B.n696 B.n695 585
R432 B.n697 B.n696 585
R433 B.n694 B.n31 585
R434 B.n31 B.n30 585
R435 B.n693 B.n692 585
R436 B.n692 B.n691 585
R437 B.n33 B.n32 585
R438 B.n690 B.n33 585
R439 B.n688 B.n687 585
R440 B.n689 B.n688 585
R441 B.n686 B.n38 585
R442 B.n38 B.n37 585
R443 B.n685 B.n684 585
R444 B.n684 B.n683 585
R445 B.n40 B.n39 585
R446 B.n682 B.n40 585
R447 B.n680 B.n679 585
R448 B.n681 B.n680 585
R449 B.n678 B.n45 585
R450 B.n45 B.n44 585
R451 B.n677 B.n676 585
R452 B.n676 B.n675 585
R453 B.n47 B.n46 585
R454 B.n674 B.n47 585
R455 B.n672 B.n671 585
R456 B.n673 B.n672 585
R457 B.n670 B.n52 585
R458 B.n52 B.n51 585
R459 B.n669 B.n668 585
R460 B.n668 B.n667 585
R461 B.n54 B.n53 585
R462 B.n666 B.n54 585
R463 B.n664 B.n663 585
R464 B.n665 B.n664 585
R465 B.n662 B.n59 585
R466 B.n59 B.n58 585
R467 B.n661 B.n660 585
R468 B.n660 B.n659 585
R469 B.n61 B.n60 585
R470 B.n658 B.n61 585
R471 B.n725 B.n724 585
R472 B.n723 B.n2 585
R473 B.n107 B.n61 497.305
R474 B.n656 B.n63 497.305
R475 B.n511 B.n318 497.305
R476 B.n507 B.n316 497.305
R477 B.n105 B.t8 293.253
R478 B.n102 B.t4 293.253
R479 B.n361 B.t11 293.253
R480 B.n358 B.t15 293.253
R481 B.n657 B.n100 256.663
R482 B.n657 B.n99 256.663
R483 B.n657 B.n98 256.663
R484 B.n657 B.n97 256.663
R485 B.n657 B.n96 256.663
R486 B.n657 B.n95 256.663
R487 B.n657 B.n94 256.663
R488 B.n657 B.n93 256.663
R489 B.n657 B.n92 256.663
R490 B.n657 B.n91 256.663
R491 B.n657 B.n90 256.663
R492 B.n657 B.n89 256.663
R493 B.n657 B.n88 256.663
R494 B.n657 B.n87 256.663
R495 B.n657 B.n86 256.663
R496 B.n657 B.n85 256.663
R497 B.n657 B.n84 256.663
R498 B.n657 B.n83 256.663
R499 B.n657 B.n82 256.663
R500 B.n657 B.n81 256.663
R501 B.n657 B.n80 256.663
R502 B.n657 B.n79 256.663
R503 B.n657 B.n78 256.663
R504 B.n657 B.n77 256.663
R505 B.n657 B.n76 256.663
R506 B.n657 B.n75 256.663
R507 B.n657 B.n74 256.663
R508 B.n657 B.n73 256.663
R509 B.n657 B.n72 256.663
R510 B.n657 B.n71 256.663
R511 B.n657 B.n70 256.663
R512 B.n657 B.n69 256.663
R513 B.n657 B.n68 256.663
R514 B.n657 B.n67 256.663
R515 B.n657 B.n66 256.663
R516 B.n657 B.n65 256.663
R517 B.n657 B.n64 256.663
R518 B.n509 B.n508 256.663
R519 B.n509 B.n321 256.663
R520 B.n509 B.n322 256.663
R521 B.n509 B.n323 256.663
R522 B.n509 B.n324 256.663
R523 B.n509 B.n325 256.663
R524 B.n509 B.n326 256.663
R525 B.n509 B.n327 256.663
R526 B.n509 B.n328 256.663
R527 B.n509 B.n329 256.663
R528 B.n509 B.n330 256.663
R529 B.n509 B.n331 256.663
R530 B.n509 B.n332 256.663
R531 B.n509 B.n333 256.663
R532 B.n509 B.n334 256.663
R533 B.n509 B.n335 256.663
R534 B.n509 B.n336 256.663
R535 B.n509 B.n337 256.663
R536 B.n509 B.n338 256.663
R537 B.n509 B.n339 256.663
R538 B.n509 B.n340 256.663
R539 B.n509 B.n341 256.663
R540 B.n509 B.n342 256.663
R541 B.n509 B.n343 256.663
R542 B.n509 B.n344 256.663
R543 B.n509 B.n345 256.663
R544 B.n509 B.n346 256.663
R545 B.n509 B.n347 256.663
R546 B.n509 B.n348 256.663
R547 B.n509 B.n349 256.663
R548 B.n509 B.n350 256.663
R549 B.n509 B.n351 256.663
R550 B.n509 B.n352 256.663
R551 B.n509 B.n353 256.663
R552 B.n509 B.n354 256.663
R553 B.n509 B.n355 256.663
R554 B.n510 B.n509 256.663
R555 B.n727 B.n726 256.663
R556 B.n111 B.n110 163.367
R557 B.n115 B.n114 163.367
R558 B.n119 B.n118 163.367
R559 B.n123 B.n122 163.367
R560 B.n127 B.n126 163.367
R561 B.n131 B.n130 163.367
R562 B.n135 B.n134 163.367
R563 B.n139 B.n138 163.367
R564 B.n143 B.n142 163.367
R565 B.n147 B.n146 163.367
R566 B.n151 B.n150 163.367
R567 B.n155 B.n154 163.367
R568 B.n159 B.n158 163.367
R569 B.n163 B.n162 163.367
R570 B.n167 B.n166 163.367
R571 B.n171 B.n170 163.367
R572 B.n176 B.n175 163.367
R573 B.n180 B.n179 163.367
R574 B.n184 B.n183 163.367
R575 B.n188 B.n187 163.367
R576 B.n192 B.n191 163.367
R577 B.n196 B.n195 163.367
R578 B.n200 B.n199 163.367
R579 B.n204 B.n203 163.367
R580 B.n208 B.n207 163.367
R581 B.n212 B.n211 163.367
R582 B.n216 B.n215 163.367
R583 B.n220 B.n219 163.367
R584 B.n224 B.n223 163.367
R585 B.n228 B.n227 163.367
R586 B.n232 B.n231 163.367
R587 B.n236 B.n235 163.367
R588 B.n240 B.n239 163.367
R589 B.n244 B.n243 163.367
R590 B.n248 B.n247 163.367
R591 B.n252 B.n251 163.367
R592 B.n656 B.n101 163.367
R593 B.n515 B.n318 163.367
R594 B.n515 B.n312 163.367
R595 B.n523 B.n312 163.367
R596 B.n523 B.n310 163.367
R597 B.n527 B.n310 163.367
R598 B.n527 B.n304 163.367
R599 B.n535 B.n304 163.367
R600 B.n535 B.n302 163.367
R601 B.n539 B.n302 163.367
R602 B.n539 B.n296 163.367
R603 B.n547 B.n296 163.367
R604 B.n547 B.n294 163.367
R605 B.n551 B.n294 163.367
R606 B.n551 B.n288 163.367
R607 B.n559 B.n288 163.367
R608 B.n559 B.n286 163.367
R609 B.n563 B.n286 163.367
R610 B.n563 B.n280 163.367
R611 B.n571 B.n280 163.367
R612 B.n571 B.n278 163.367
R613 B.n575 B.n278 163.367
R614 B.n575 B.n272 163.367
R615 B.n583 B.n272 163.367
R616 B.n583 B.n270 163.367
R617 B.n587 B.n270 163.367
R618 B.n587 B.n264 163.367
R619 B.n595 B.n264 163.367
R620 B.n595 B.n262 163.367
R621 B.n600 B.n262 163.367
R622 B.n600 B.n256 163.367
R623 B.n608 B.n256 163.367
R624 B.n609 B.n608 163.367
R625 B.n609 B.n5 163.367
R626 B.n6 B.n5 163.367
R627 B.n7 B.n6 163.367
R628 B.n615 B.n7 163.367
R629 B.n616 B.n615 163.367
R630 B.n616 B.n13 163.367
R631 B.n14 B.n13 163.367
R632 B.n15 B.n14 163.367
R633 B.n621 B.n15 163.367
R634 B.n621 B.n20 163.367
R635 B.n21 B.n20 163.367
R636 B.n22 B.n21 163.367
R637 B.n626 B.n22 163.367
R638 B.n626 B.n27 163.367
R639 B.n28 B.n27 163.367
R640 B.n29 B.n28 163.367
R641 B.n631 B.n29 163.367
R642 B.n631 B.n34 163.367
R643 B.n35 B.n34 163.367
R644 B.n36 B.n35 163.367
R645 B.n636 B.n36 163.367
R646 B.n636 B.n41 163.367
R647 B.n42 B.n41 163.367
R648 B.n43 B.n42 163.367
R649 B.n641 B.n43 163.367
R650 B.n641 B.n48 163.367
R651 B.n49 B.n48 163.367
R652 B.n50 B.n49 163.367
R653 B.n646 B.n50 163.367
R654 B.n646 B.n55 163.367
R655 B.n56 B.n55 163.367
R656 B.n57 B.n56 163.367
R657 B.n651 B.n57 163.367
R658 B.n651 B.n62 163.367
R659 B.n63 B.n62 163.367
R660 B.n357 B.n356 163.367
R661 B.n502 B.n356 163.367
R662 B.n500 B.n499 163.367
R663 B.n496 B.n495 163.367
R664 B.n492 B.n491 163.367
R665 B.n488 B.n487 163.367
R666 B.n484 B.n483 163.367
R667 B.n480 B.n479 163.367
R668 B.n476 B.n475 163.367
R669 B.n472 B.n471 163.367
R670 B.n468 B.n467 163.367
R671 B.n464 B.n463 163.367
R672 B.n460 B.n459 163.367
R673 B.n456 B.n455 163.367
R674 B.n452 B.n451 163.367
R675 B.n448 B.n447 163.367
R676 B.n444 B.n443 163.367
R677 B.n440 B.n439 163.367
R678 B.n436 B.n435 163.367
R679 B.n432 B.n431 163.367
R680 B.n428 B.n427 163.367
R681 B.n423 B.n422 163.367
R682 B.n419 B.n418 163.367
R683 B.n415 B.n414 163.367
R684 B.n411 B.n410 163.367
R685 B.n407 B.n406 163.367
R686 B.n403 B.n402 163.367
R687 B.n399 B.n398 163.367
R688 B.n395 B.n394 163.367
R689 B.n391 B.n390 163.367
R690 B.n387 B.n386 163.367
R691 B.n383 B.n382 163.367
R692 B.n379 B.n378 163.367
R693 B.n375 B.n374 163.367
R694 B.n371 B.n370 163.367
R695 B.n367 B.n366 163.367
R696 B.n363 B.n320 163.367
R697 B.n517 B.n316 163.367
R698 B.n517 B.n314 163.367
R699 B.n521 B.n314 163.367
R700 B.n521 B.n308 163.367
R701 B.n529 B.n308 163.367
R702 B.n529 B.n306 163.367
R703 B.n533 B.n306 163.367
R704 B.n533 B.n300 163.367
R705 B.n541 B.n300 163.367
R706 B.n541 B.n298 163.367
R707 B.n545 B.n298 163.367
R708 B.n545 B.n292 163.367
R709 B.n553 B.n292 163.367
R710 B.n553 B.n290 163.367
R711 B.n557 B.n290 163.367
R712 B.n557 B.n284 163.367
R713 B.n565 B.n284 163.367
R714 B.n565 B.n282 163.367
R715 B.n569 B.n282 163.367
R716 B.n569 B.n276 163.367
R717 B.n577 B.n276 163.367
R718 B.n577 B.n274 163.367
R719 B.n581 B.n274 163.367
R720 B.n581 B.n268 163.367
R721 B.n589 B.n268 163.367
R722 B.n589 B.n266 163.367
R723 B.n593 B.n266 163.367
R724 B.n593 B.n260 163.367
R725 B.n602 B.n260 163.367
R726 B.n602 B.n258 163.367
R727 B.n606 B.n258 163.367
R728 B.n606 B.n3 163.367
R729 B.n725 B.n3 163.367
R730 B.n721 B.n2 163.367
R731 B.n721 B.n720 163.367
R732 B.n720 B.n9 163.367
R733 B.n716 B.n9 163.367
R734 B.n716 B.n11 163.367
R735 B.n712 B.n11 163.367
R736 B.n712 B.n17 163.367
R737 B.n708 B.n17 163.367
R738 B.n708 B.n19 163.367
R739 B.n704 B.n19 163.367
R740 B.n704 B.n24 163.367
R741 B.n700 B.n24 163.367
R742 B.n700 B.n26 163.367
R743 B.n696 B.n26 163.367
R744 B.n696 B.n31 163.367
R745 B.n692 B.n31 163.367
R746 B.n692 B.n33 163.367
R747 B.n688 B.n33 163.367
R748 B.n688 B.n38 163.367
R749 B.n684 B.n38 163.367
R750 B.n684 B.n40 163.367
R751 B.n680 B.n40 163.367
R752 B.n680 B.n45 163.367
R753 B.n676 B.n45 163.367
R754 B.n676 B.n47 163.367
R755 B.n672 B.n47 163.367
R756 B.n672 B.n52 163.367
R757 B.n668 B.n52 163.367
R758 B.n668 B.n54 163.367
R759 B.n664 B.n54 163.367
R760 B.n664 B.n59 163.367
R761 B.n660 B.n59 163.367
R762 B.n660 B.n61 163.367
R763 B.n102 B.t6 126.907
R764 B.n361 B.t14 126.907
R765 B.n105 B.t9 126.897
R766 B.n358 B.t17 126.897
R767 B.n509 B.n317 91.7636
R768 B.n658 B.n657 91.7636
R769 B.n107 B.n64 71.676
R770 B.n111 B.n65 71.676
R771 B.n115 B.n66 71.676
R772 B.n119 B.n67 71.676
R773 B.n123 B.n68 71.676
R774 B.n127 B.n69 71.676
R775 B.n131 B.n70 71.676
R776 B.n135 B.n71 71.676
R777 B.n139 B.n72 71.676
R778 B.n143 B.n73 71.676
R779 B.n147 B.n74 71.676
R780 B.n151 B.n75 71.676
R781 B.n155 B.n76 71.676
R782 B.n159 B.n77 71.676
R783 B.n163 B.n78 71.676
R784 B.n167 B.n79 71.676
R785 B.n171 B.n80 71.676
R786 B.n176 B.n81 71.676
R787 B.n180 B.n82 71.676
R788 B.n184 B.n83 71.676
R789 B.n188 B.n84 71.676
R790 B.n192 B.n85 71.676
R791 B.n196 B.n86 71.676
R792 B.n200 B.n87 71.676
R793 B.n204 B.n88 71.676
R794 B.n208 B.n89 71.676
R795 B.n212 B.n90 71.676
R796 B.n216 B.n91 71.676
R797 B.n220 B.n92 71.676
R798 B.n224 B.n93 71.676
R799 B.n228 B.n94 71.676
R800 B.n232 B.n95 71.676
R801 B.n236 B.n96 71.676
R802 B.n240 B.n97 71.676
R803 B.n244 B.n98 71.676
R804 B.n248 B.n99 71.676
R805 B.n252 B.n100 71.676
R806 B.n101 B.n100 71.676
R807 B.n251 B.n99 71.676
R808 B.n247 B.n98 71.676
R809 B.n243 B.n97 71.676
R810 B.n239 B.n96 71.676
R811 B.n235 B.n95 71.676
R812 B.n231 B.n94 71.676
R813 B.n227 B.n93 71.676
R814 B.n223 B.n92 71.676
R815 B.n219 B.n91 71.676
R816 B.n215 B.n90 71.676
R817 B.n211 B.n89 71.676
R818 B.n207 B.n88 71.676
R819 B.n203 B.n87 71.676
R820 B.n199 B.n86 71.676
R821 B.n195 B.n85 71.676
R822 B.n191 B.n84 71.676
R823 B.n187 B.n83 71.676
R824 B.n183 B.n82 71.676
R825 B.n179 B.n81 71.676
R826 B.n175 B.n80 71.676
R827 B.n170 B.n79 71.676
R828 B.n166 B.n78 71.676
R829 B.n162 B.n77 71.676
R830 B.n158 B.n76 71.676
R831 B.n154 B.n75 71.676
R832 B.n150 B.n74 71.676
R833 B.n146 B.n73 71.676
R834 B.n142 B.n72 71.676
R835 B.n138 B.n71 71.676
R836 B.n134 B.n70 71.676
R837 B.n130 B.n69 71.676
R838 B.n126 B.n68 71.676
R839 B.n122 B.n67 71.676
R840 B.n118 B.n66 71.676
R841 B.n114 B.n65 71.676
R842 B.n110 B.n64 71.676
R843 B.n508 B.n507 71.676
R844 B.n502 B.n321 71.676
R845 B.n499 B.n322 71.676
R846 B.n495 B.n323 71.676
R847 B.n491 B.n324 71.676
R848 B.n487 B.n325 71.676
R849 B.n483 B.n326 71.676
R850 B.n479 B.n327 71.676
R851 B.n475 B.n328 71.676
R852 B.n471 B.n329 71.676
R853 B.n467 B.n330 71.676
R854 B.n463 B.n331 71.676
R855 B.n459 B.n332 71.676
R856 B.n455 B.n333 71.676
R857 B.n451 B.n334 71.676
R858 B.n447 B.n335 71.676
R859 B.n443 B.n336 71.676
R860 B.n439 B.n337 71.676
R861 B.n435 B.n338 71.676
R862 B.n431 B.n339 71.676
R863 B.n427 B.n340 71.676
R864 B.n422 B.n341 71.676
R865 B.n418 B.n342 71.676
R866 B.n414 B.n343 71.676
R867 B.n410 B.n344 71.676
R868 B.n406 B.n345 71.676
R869 B.n402 B.n346 71.676
R870 B.n398 B.n347 71.676
R871 B.n394 B.n348 71.676
R872 B.n390 B.n349 71.676
R873 B.n386 B.n350 71.676
R874 B.n382 B.n351 71.676
R875 B.n378 B.n352 71.676
R876 B.n374 B.n353 71.676
R877 B.n370 B.n354 71.676
R878 B.n366 B.n355 71.676
R879 B.n510 B.n320 71.676
R880 B.n508 B.n357 71.676
R881 B.n500 B.n321 71.676
R882 B.n496 B.n322 71.676
R883 B.n492 B.n323 71.676
R884 B.n488 B.n324 71.676
R885 B.n484 B.n325 71.676
R886 B.n480 B.n326 71.676
R887 B.n476 B.n327 71.676
R888 B.n472 B.n328 71.676
R889 B.n468 B.n329 71.676
R890 B.n464 B.n330 71.676
R891 B.n460 B.n331 71.676
R892 B.n456 B.n332 71.676
R893 B.n452 B.n333 71.676
R894 B.n448 B.n334 71.676
R895 B.n444 B.n335 71.676
R896 B.n440 B.n336 71.676
R897 B.n436 B.n337 71.676
R898 B.n432 B.n338 71.676
R899 B.n428 B.n339 71.676
R900 B.n423 B.n340 71.676
R901 B.n419 B.n341 71.676
R902 B.n415 B.n342 71.676
R903 B.n411 B.n343 71.676
R904 B.n407 B.n344 71.676
R905 B.n403 B.n345 71.676
R906 B.n399 B.n346 71.676
R907 B.n395 B.n347 71.676
R908 B.n391 B.n348 71.676
R909 B.n387 B.n349 71.676
R910 B.n383 B.n350 71.676
R911 B.n379 B.n351 71.676
R912 B.n375 B.n352 71.676
R913 B.n371 B.n353 71.676
R914 B.n367 B.n354 71.676
R915 B.n363 B.n355 71.676
R916 B.n511 B.n510 71.676
R917 B.n726 B.n725 71.676
R918 B.n726 B.n2 71.676
R919 B.n103 B.t7 71.2471
R920 B.n362 B.t13 71.2471
R921 B.n106 B.t10 71.2364
R922 B.n359 B.t16 71.2364
R923 B.n173 B.n106 59.5399
R924 B.n104 B.n103 59.5399
R925 B.n425 B.n362 59.5399
R926 B.n360 B.n359 59.5399
R927 B.n106 B.n105 55.6611
R928 B.n103 B.n102 55.6611
R929 B.n362 B.n361 55.6611
R930 B.n359 B.n358 55.6611
R931 B.n516 B.n317 52.4365
R932 B.n516 B.n313 52.4365
R933 B.n522 B.n313 52.4365
R934 B.n522 B.n309 52.4365
R935 B.n528 B.n309 52.4365
R936 B.n528 B.n305 52.4365
R937 B.n534 B.n305 52.4365
R938 B.n540 B.n301 52.4365
R939 B.n540 B.n297 52.4365
R940 B.n546 B.n297 52.4365
R941 B.n546 B.n293 52.4365
R942 B.n552 B.n293 52.4365
R943 B.n552 B.n289 52.4365
R944 B.n558 B.n289 52.4365
R945 B.n558 B.n285 52.4365
R946 B.n564 B.n285 52.4365
R947 B.n564 B.n281 52.4365
R948 B.n570 B.n281 52.4365
R949 B.n576 B.n277 52.4365
R950 B.n576 B.n273 52.4365
R951 B.n582 B.n273 52.4365
R952 B.n582 B.n269 52.4365
R953 B.n588 B.n269 52.4365
R954 B.n588 B.n265 52.4365
R955 B.n594 B.n265 52.4365
R956 B.n601 B.n261 52.4365
R957 B.n601 B.n257 52.4365
R958 B.n607 B.n257 52.4365
R959 B.n607 B.n4 52.4365
R960 B.n724 B.n4 52.4365
R961 B.n724 B.n723 52.4365
R962 B.n723 B.n722 52.4365
R963 B.n722 B.n8 52.4365
R964 B.n12 B.n8 52.4365
R965 B.n715 B.n12 52.4365
R966 B.n715 B.n714 52.4365
R967 B.n713 B.n16 52.4365
R968 B.n707 B.n16 52.4365
R969 B.n707 B.n706 52.4365
R970 B.n706 B.n705 52.4365
R971 B.n705 B.n23 52.4365
R972 B.n699 B.n23 52.4365
R973 B.n699 B.n698 52.4365
R974 B.n697 B.n30 52.4365
R975 B.n691 B.n30 52.4365
R976 B.n691 B.n690 52.4365
R977 B.n690 B.n689 52.4365
R978 B.n689 B.n37 52.4365
R979 B.n683 B.n37 52.4365
R980 B.n683 B.n682 52.4365
R981 B.n682 B.n681 52.4365
R982 B.n681 B.n44 52.4365
R983 B.n675 B.n44 52.4365
R984 B.n675 B.n674 52.4365
R985 B.n673 B.n51 52.4365
R986 B.n667 B.n51 52.4365
R987 B.n667 B.n666 52.4365
R988 B.n666 B.n665 52.4365
R989 B.n665 B.n58 52.4365
R990 B.n659 B.n58 52.4365
R991 B.n659 B.n658 52.4365
R992 B.t3 B.n277 40.0986
R993 B.n698 B.t1 40.0986
R994 B.n594 B.t2 35.4719
R995 B.t0 B.n713 35.4719
R996 B.n506 B.n315 32.3127
R997 B.n513 B.n512 32.3127
R998 B.n655 B.n654 32.3127
R999 B.n108 B.n60 32.3127
R1000 B.n534 B.t12 30.8452
R1001 B.t5 B.n673 30.8452
R1002 B.t12 B.n301 21.5918
R1003 B.n674 B.t5 21.5918
R1004 B B.n727 18.0485
R1005 B.t2 B.n261 16.9651
R1006 B.n714 B.t0 16.9651
R1007 B.n570 B.t3 12.3384
R1008 B.t1 B.n697 12.3384
R1009 B.n518 B.n315 10.6151
R1010 B.n519 B.n518 10.6151
R1011 B.n520 B.n519 10.6151
R1012 B.n520 B.n307 10.6151
R1013 B.n530 B.n307 10.6151
R1014 B.n531 B.n530 10.6151
R1015 B.n532 B.n531 10.6151
R1016 B.n532 B.n299 10.6151
R1017 B.n542 B.n299 10.6151
R1018 B.n543 B.n542 10.6151
R1019 B.n544 B.n543 10.6151
R1020 B.n544 B.n291 10.6151
R1021 B.n554 B.n291 10.6151
R1022 B.n555 B.n554 10.6151
R1023 B.n556 B.n555 10.6151
R1024 B.n556 B.n283 10.6151
R1025 B.n566 B.n283 10.6151
R1026 B.n567 B.n566 10.6151
R1027 B.n568 B.n567 10.6151
R1028 B.n568 B.n275 10.6151
R1029 B.n578 B.n275 10.6151
R1030 B.n579 B.n578 10.6151
R1031 B.n580 B.n579 10.6151
R1032 B.n580 B.n267 10.6151
R1033 B.n590 B.n267 10.6151
R1034 B.n591 B.n590 10.6151
R1035 B.n592 B.n591 10.6151
R1036 B.n592 B.n259 10.6151
R1037 B.n603 B.n259 10.6151
R1038 B.n604 B.n603 10.6151
R1039 B.n605 B.n604 10.6151
R1040 B.n605 B.n0 10.6151
R1041 B.n506 B.n505 10.6151
R1042 B.n505 B.n504 10.6151
R1043 B.n504 B.n503 10.6151
R1044 B.n503 B.n501 10.6151
R1045 B.n501 B.n498 10.6151
R1046 B.n498 B.n497 10.6151
R1047 B.n497 B.n494 10.6151
R1048 B.n494 B.n493 10.6151
R1049 B.n493 B.n490 10.6151
R1050 B.n490 B.n489 10.6151
R1051 B.n489 B.n486 10.6151
R1052 B.n486 B.n485 10.6151
R1053 B.n485 B.n482 10.6151
R1054 B.n482 B.n481 10.6151
R1055 B.n481 B.n478 10.6151
R1056 B.n478 B.n477 10.6151
R1057 B.n477 B.n474 10.6151
R1058 B.n474 B.n473 10.6151
R1059 B.n473 B.n470 10.6151
R1060 B.n470 B.n469 10.6151
R1061 B.n469 B.n466 10.6151
R1062 B.n466 B.n465 10.6151
R1063 B.n465 B.n462 10.6151
R1064 B.n462 B.n461 10.6151
R1065 B.n461 B.n458 10.6151
R1066 B.n458 B.n457 10.6151
R1067 B.n457 B.n454 10.6151
R1068 B.n454 B.n453 10.6151
R1069 B.n453 B.n450 10.6151
R1070 B.n450 B.n449 10.6151
R1071 B.n449 B.n446 10.6151
R1072 B.n446 B.n445 10.6151
R1073 B.n442 B.n441 10.6151
R1074 B.n441 B.n438 10.6151
R1075 B.n438 B.n437 10.6151
R1076 B.n437 B.n434 10.6151
R1077 B.n434 B.n433 10.6151
R1078 B.n433 B.n430 10.6151
R1079 B.n430 B.n429 10.6151
R1080 B.n429 B.n426 10.6151
R1081 B.n424 B.n421 10.6151
R1082 B.n421 B.n420 10.6151
R1083 B.n420 B.n417 10.6151
R1084 B.n417 B.n416 10.6151
R1085 B.n416 B.n413 10.6151
R1086 B.n413 B.n412 10.6151
R1087 B.n412 B.n409 10.6151
R1088 B.n409 B.n408 10.6151
R1089 B.n408 B.n405 10.6151
R1090 B.n405 B.n404 10.6151
R1091 B.n404 B.n401 10.6151
R1092 B.n401 B.n400 10.6151
R1093 B.n400 B.n397 10.6151
R1094 B.n397 B.n396 10.6151
R1095 B.n396 B.n393 10.6151
R1096 B.n393 B.n392 10.6151
R1097 B.n392 B.n389 10.6151
R1098 B.n389 B.n388 10.6151
R1099 B.n388 B.n385 10.6151
R1100 B.n385 B.n384 10.6151
R1101 B.n384 B.n381 10.6151
R1102 B.n381 B.n380 10.6151
R1103 B.n380 B.n377 10.6151
R1104 B.n377 B.n376 10.6151
R1105 B.n376 B.n373 10.6151
R1106 B.n373 B.n372 10.6151
R1107 B.n372 B.n369 10.6151
R1108 B.n369 B.n368 10.6151
R1109 B.n368 B.n365 10.6151
R1110 B.n365 B.n364 10.6151
R1111 B.n364 B.n319 10.6151
R1112 B.n512 B.n319 10.6151
R1113 B.n514 B.n513 10.6151
R1114 B.n514 B.n311 10.6151
R1115 B.n524 B.n311 10.6151
R1116 B.n525 B.n524 10.6151
R1117 B.n526 B.n525 10.6151
R1118 B.n526 B.n303 10.6151
R1119 B.n536 B.n303 10.6151
R1120 B.n537 B.n536 10.6151
R1121 B.n538 B.n537 10.6151
R1122 B.n538 B.n295 10.6151
R1123 B.n548 B.n295 10.6151
R1124 B.n549 B.n548 10.6151
R1125 B.n550 B.n549 10.6151
R1126 B.n550 B.n287 10.6151
R1127 B.n560 B.n287 10.6151
R1128 B.n561 B.n560 10.6151
R1129 B.n562 B.n561 10.6151
R1130 B.n562 B.n279 10.6151
R1131 B.n572 B.n279 10.6151
R1132 B.n573 B.n572 10.6151
R1133 B.n574 B.n573 10.6151
R1134 B.n574 B.n271 10.6151
R1135 B.n584 B.n271 10.6151
R1136 B.n585 B.n584 10.6151
R1137 B.n586 B.n585 10.6151
R1138 B.n586 B.n263 10.6151
R1139 B.n596 B.n263 10.6151
R1140 B.n597 B.n596 10.6151
R1141 B.n599 B.n597 10.6151
R1142 B.n599 B.n598 10.6151
R1143 B.n598 B.n255 10.6151
R1144 B.n610 B.n255 10.6151
R1145 B.n611 B.n610 10.6151
R1146 B.n612 B.n611 10.6151
R1147 B.n613 B.n612 10.6151
R1148 B.n614 B.n613 10.6151
R1149 B.n617 B.n614 10.6151
R1150 B.n618 B.n617 10.6151
R1151 B.n619 B.n618 10.6151
R1152 B.n620 B.n619 10.6151
R1153 B.n622 B.n620 10.6151
R1154 B.n623 B.n622 10.6151
R1155 B.n624 B.n623 10.6151
R1156 B.n625 B.n624 10.6151
R1157 B.n627 B.n625 10.6151
R1158 B.n628 B.n627 10.6151
R1159 B.n629 B.n628 10.6151
R1160 B.n630 B.n629 10.6151
R1161 B.n632 B.n630 10.6151
R1162 B.n633 B.n632 10.6151
R1163 B.n634 B.n633 10.6151
R1164 B.n635 B.n634 10.6151
R1165 B.n637 B.n635 10.6151
R1166 B.n638 B.n637 10.6151
R1167 B.n639 B.n638 10.6151
R1168 B.n640 B.n639 10.6151
R1169 B.n642 B.n640 10.6151
R1170 B.n643 B.n642 10.6151
R1171 B.n644 B.n643 10.6151
R1172 B.n645 B.n644 10.6151
R1173 B.n647 B.n645 10.6151
R1174 B.n648 B.n647 10.6151
R1175 B.n649 B.n648 10.6151
R1176 B.n650 B.n649 10.6151
R1177 B.n652 B.n650 10.6151
R1178 B.n653 B.n652 10.6151
R1179 B.n654 B.n653 10.6151
R1180 B.n719 B.n1 10.6151
R1181 B.n719 B.n718 10.6151
R1182 B.n718 B.n717 10.6151
R1183 B.n717 B.n10 10.6151
R1184 B.n711 B.n10 10.6151
R1185 B.n711 B.n710 10.6151
R1186 B.n710 B.n709 10.6151
R1187 B.n709 B.n18 10.6151
R1188 B.n703 B.n18 10.6151
R1189 B.n703 B.n702 10.6151
R1190 B.n702 B.n701 10.6151
R1191 B.n701 B.n25 10.6151
R1192 B.n695 B.n25 10.6151
R1193 B.n695 B.n694 10.6151
R1194 B.n694 B.n693 10.6151
R1195 B.n693 B.n32 10.6151
R1196 B.n687 B.n32 10.6151
R1197 B.n687 B.n686 10.6151
R1198 B.n686 B.n685 10.6151
R1199 B.n685 B.n39 10.6151
R1200 B.n679 B.n39 10.6151
R1201 B.n679 B.n678 10.6151
R1202 B.n678 B.n677 10.6151
R1203 B.n677 B.n46 10.6151
R1204 B.n671 B.n46 10.6151
R1205 B.n671 B.n670 10.6151
R1206 B.n670 B.n669 10.6151
R1207 B.n669 B.n53 10.6151
R1208 B.n663 B.n53 10.6151
R1209 B.n663 B.n662 10.6151
R1210 B.n662 B.n661 10.6151
R1211 B.n661 B.n60 10.6151
R1212 B.n109 B.n108 10.6151
R1213 B.n112 B.n109 10.6151
R1214 B.n113 B.n112 10.6151
R1215 B.n116 B.n113 10.6151
R1216 B.n117 B.n116 10.6151
R1217 B.n120 B.n117 10.6151
R1218 B.n121 B.n120 10.6151
R1219 B.n124 B.n121 10.6151
R1220 B.n125 B.n124 10.6151
R1221 B.n128 B.n125 10.6151
R1222 B.n129 B.n128 10.6151
R1223 B.n132 B.n129 10.6151
R1224 B.n133 B.n132 10.6151
R1225 B.n136 B.n133 10.6151
R1226 B.n137 B.n136 10.6151
R1227 B.n140 B.n137 10.6151
R1228 B.n141 B.n140 10.6151
R1229 B.n144 B.n141 10.6151
R1230 B.n145 B.n144 10.6151
R1231 B.n148 B.n145 10.6151
R1232 B.n149 B.n148 10.6151
R1233 B.n152 B.n149 10.6151
R1234 B.n153 B.n152 10.6151
R1235 B.n156 B.n153 10.6151
R1236 B.n157 B.n156 10.6151
R1237 B.n160 B.n157 10.6151
R1238 B.n161 B.n160 10.6151
R1239 B.n164 B.n161 10.6151
R1240 B.n165 B.n164 10.6151
R1241 B.n168 B.n165 10.6151
R1242 B.n169 B.n168 10.6151
R1243 B.n172 B.n169 10.6151
R1244 B.n177 B.n174 10.6151
R1245 B.n178 B.n177 10.6151
R1246 B.n181 B.n178 10.6151
R1247 B.n182 B.n181 10.6151
R1248 B.n185 B.n182 10.6151
R1249 B.n186 B.n185 10.6151
R1250 B.n189 B.n186 10.6151
R1251 B.n190 B.n189 10.6151
R1252 B.n194 B.n193 10.6151
R1253 B.n197 B.n194 10.6151
R1254 B.n198 B.n197 10.6151
R1255 B.n201 B.n198 10.6151
R1256 B.n202 B.n201 10.6151
R1257 B.n205 B.n202 10.6151
R1258 B.n206 B.n205 10.6151
R1259 B.n209 B.n206 10.6151
R1260 B.n210 B.n209 10.6151
R1261 B.n213 B.n210 10.6151
R1262 B.n214 B.n213 10.6151
R1263 B.n217 B.n214 10.6151
R1264 B.n218 B.n217 10.6151
R1265 B.n221 B.n218 10.6151
R1266 B.n222 B.n221 10.6151
R1267 B.n225 B.n222 10.6151
R1268 B.n226 B.n225 10.6151
R1269 B.n229 B.n226 10.6151
R1270 B.n230 B.n229 10.6151
R1271 B.n233 B.n230 10.6151
R1272 B.n234 B.n233 10.6151
R1273 B.n237 B.n234 10.6151
R1274 B.n238 B.n237 10.6151
R1275 B.n241 B.n238 10.6151
R1276 B.n242 B.n241 10.6151
R1277 B.n245 B.n242 10.6151
R1278 B.n246 B.n245 10.6151
R1279 B.n249 B.n246 10.6151
R1280 B.n250 B.n249 10.6151
R1281 B.n253 B.n250 10.6151
R1282 B.n254 B.n253 10.6151
R1283 B.n655 B.n254 10.6151
R1284 B.n727 B.n0 8.11757
R1285 B.n727 B.n1 8.11757
R1286 B.n442 B.n360 6.5566
R1287 B.n426 B.n425 6.5566
R1288 B.n174 B.n173 6.5566
R1289 B.n190 B.n104 6.5566
R1290 B.n445 B.n360 4.05904
R1291 B.n425 B.n424 4.05904
R1292 B.n173 B.n172 4.05904
R1293 B.n193 B.n104 4.05904
R1294 VN.n0 VN.t2 121.041
R1295 VN.n1 VN.t3 121.041
R1296 VN.n0 VN.t0 120.276
R1297 VN.n1 VN.t1 120.276
R1298 VN VN.n1 48.5517
R1299 VN VN.n0 4.44942
R1300 VDD2.n2 VDD2.n0 104.231
R1301 VDD2.n2 VDD2.n1 65.3435
R1302 VDD2.n1 VDD2.t2 2.20295
R1303 VDD2.n1 VDD2.t0 2.20295
R1304 VDD2.n0 VDD2.t1 2.20295
R1305 VDD2.n0 VDD2.t3 2.20295
R1306 VDD2 VDD2.n2 0.0586897
C0 VTAIL VDD2 4.72982f
C1 VDD1 VP 3.8596f
C2 VDD1 VDD2 1.01961f
C3 VN VTAIL 3.65574f
C4 VDD2 VP 0.390622f
C5 VN VDD1 0.14908f
C6 VDD1 VTAIL 4.67602f
C7 VN VP 5.59058f
C8 VN VDD2 3.61879f
C9 VTAIL VP 3.66985f
C10 VDD2 B 3.492941f
C11 VDD1 B 7.34688f
C12 VTAIL B 8.238849f
C13 VN B 10.3425f
C14 VP B 8.603067f
C15 VDD2.t1 B 0.191342f
C16 VDD2.t3 B 0.191342f
C17 VDD2.n0 B 2.22117f
C18 VDD2.t2 B 0.191342f
C19 VDD2.t0 B 0.191342f
C20 VDD2.n1 B 1.67332f
C21 VDD2.n2 B 3.41962f
C22 VN.t2 B 1.88473f
C23 VN.t0 B 1.87998f
C24 VN.n0 B 1.19674f
C25 VN.t3 B 1.88473f
C26 VN.t1 B 1.87998f
C27 VN.n1 B 2.53893f
C28 VDD1.t0 B 0.19591f
C29 VDD1.t3 B 0.19591f
C30 VDD1.n0 B 1.71367f
C31 VDD1.t2 B 0.19591f
C32 VDD1.t1 B 0.19591f
C33 VDD1.n1 B 2.2997f
C34 VTAIL.t0 B 1.32336f
C35 VTAIL.n0 B 0.316871f
C36 VTAIL.t4 B 1.32336f
C37 VTAIL.n1 B 0.383264f
C38 VTAIL.t6 B 1.32336f
C39 VTAIL.n2 B 1.17003f
C40 VTAIL.t3 B 1.32336f
C41 VTAIL.n3 B 1.17002f
C42 VTAIL.t2 B 1.32336f
C43 VTAIL.n4 B 0.38326f
C44 VTAIL.t7 B 1.32336f
C45 VTAIL.n5 B 0.38326f
C46 VTAIL.t5 B 1.32336f
C47 VTAIL.n6 B 1.17003f
C48 VTAIL.t1 B 1.32336f
C49 VTAIL.n7 B 1.09708f
C50 VP.n0 B 0.036395f
C51 VP.t2 B 1.70105f
C52 VP.n1 B 0.040299f
C53 VP.n2 B 0.027605f
C54 VP.t1 B 1.70105f
C55 VP.n3 B 0.70317f
C56 VP.t0 B 1.92936f
C57 VP.t3 B 1.93423f
C58 VP.n4 B 2.59102f
C59 VP.n5 B 1.42055f
C60 VP.n6 B 0.036395f
C61 VP.n7 B 0.035445f
C62 VP.n8 B 0.051449f
C63 VP.n9 B 0.040299f
C64 VP.n10 B 0.027605f
C65 VP.n11 B 0.027605f
C66 VP.n12 B 0.027605f
C67 VP.n13 B 0.051449f
C68 VP.n14 B 0.035445f
C69 VP.n15 B 0.70317f
C70 VP.n16 B 0.045035f
.ends

