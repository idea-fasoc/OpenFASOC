* NGSPICE file created from diff_pair_sample_0665.ext - technology: sky130A

.subckt diff_pair_sample_0665 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=6.24 pd=32.78 as=0 ps=0 w=16 l=3.56
X1 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=6.24 pd=32.78 as=0 ps=0 w=16 l=3.56
X2 VDD1.t3 VP.t0 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.64 pd=16.33 as=6.24 ps=32.78 w=16 l=3.56
X3 VTAIL.t0 VN.t0 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=6.24 pd=32.78 as=2.64 ps=16.33 w=16 l=3.56
X4 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.24 pd=32.78 as=0 ps=0 w=16 l=3.56
X5 VTAIL.t1 VN.t1 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=6.24 pd=32.78 as=2.64 ps=16.33 w=16 l=3.56
X6 VDD1.t2 VP.t1 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.64 pd=16.33 as=6.24 ps=32.78 w=16 l=3.56
X7 VTAIL.t7 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=6.24 pd=32.78 as=2.64 ps=16.33 w=16 l=3.56
X8 VDD2.t1 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.64 pd=16.33 as=6.24 ps=32.78 w=16 l=3.56
X9 VDD2.t0 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.64 pd=16.33 as=6.24 ps=32.78 w=16 l=3.56
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.24 pd=32.78 as=0 ps=0 w=16 l=3.56
X11 VTAIL.t6 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=6.24 pd=32.78 as=2.64 ps=16.33 w=16 l=3.56
R0 B.n702 B.n701 585
R1 B.n704 B.n142 585
R2 B.n707 B.n706 585
R3 B.n708 B.n141 585
R4 B.n710 B.n709 585
R5 B.n712 B.n140 585
R6 B.n715 B.n714 585
R7 B.n716 B.n139 585
R8 B.n718 B.n717 585
R9 B.n720 B.n138 585
R10 B.n723 B.n722 585
R11 B.n724 B.n137 585
R12 B.n726 B.n725 585
R13 B.n728 B.n136 585
R14 B.n731 B.n730 585
R15 B.n732 B.n135 585
R16 B.n734 B.n733 585
R17 B.n736 B.n134 585
R18 B.n739 B.n738 585
R19 B.n740 B.n133 585
R20 B.n742 B.n741 585
R21 B.n744 B.n132 585
R22 B.n747 B.n746 585
R23 B.n748 B.n131 585
R24 B.n750 B.n749 585
R25 B.n752 B.n130 585
R26 B.n755 B.n754 585
R27 B.n756 B.n129 585
R28 B.n758 B.n757 585
R29 B.n760 B.n128 585
R30 B.n763 B.n762 585
R31 B.n764 B.n127 585
R32 B.n766 B.n765 585
R33 B.n768 B.n126 585
R34 B.n771 B.n770 585
R35 B.n772 B.n125 585
R36 B.n774 B.n773 585
R37 B.n776 B.n124 585
R38 B.n779 B.n778 585
R39 B.n780 B.n123 585
R40 B.n782 B.n781 585
R41 B.n784 B.n122 585
R42 B.n787 B.n786 585
R43 B.n788 B.n121 585
R44 B.n790 B.n789 585
R45 B.n792 B.n120 585
R46 B.n795 B.n794 585
R47 B.n796 B.n119 585
R48 B.n798 B.n797 585
R49 B.n800 B.n118 585
R50 B.n803 B.n802 585
R51 B.n804 B.n114 585
R52 B.n806 B.n805 585
R53 B.n808 B.n113 585
R54 B.n811 B.n810 585
R55 B.n812 B.n112 585
R56 B.n814 B.n813 585
R57 B.n816 B.n111 585
R58 B.n819 B.n818 585
R59 B.n820 B.n110 585
R60 B.n822 B.n821 585
R61 B.n824 B.n109 585
R62 B.n827 B.n826 585
R63 B.n829 B.n106 585
R64 B.n831 B.n830 585
R65 B.n833 B.n105 585
R66 B.n836 B.n835 585
R67 B.n837 B.n104 585
R68 B.n839 B.n838 585
R69 B.n841 B.n103 585
R70 B.n844 B.n843 585
R71 B.n845 B.n102 585
R72 B.n847 B.n846 585
R73 B.n849 B.n101 585
R74 B.n852 B.n851 585
R75 B.n853 B.n100 585
R76 B.n855 B.n854 585
R77 B.n857 B.n99 585
R78 B.n860 B.n859 585
R79 B.n861 B.n98 585
R80 B.n863 B.n862 585
R81 B.n865 B.n97 585
R82 B.n868 B.n867 585
R83 B.n869 B.n96 585
R84 B.n871 B.n870 585
R85 B.n873 B.n95 585
R86 B.n876 B.n875 585
R87 B.n877 B.n94 585
R88 B.n879 B.n878 585
R89 B.n881 B.n93 585
R90 B.n884 B.n883 585
R91 B.n885 B.n92 585
R92 B.n887 B.n886 585
R93 B.n889 B.n91 585
R94 B.n892 B.n891 585
R95 B.n893 B.n90 585
R96 B.n895 B.n894 585
R97 B.n897 B.n89 585
R98 B.n900 B.n899 585
R99 B.n901 B.n88 585
R100 B.n903 B.n902 585
R101 B.n905 B.n87 585
R102 B.n908 B.n907 585
R103 B.n909 B.n86 585
R104 B.n911 B.n910 585
R105 B.n913 B.n85 585
R106 B.n916 B.n915 585
R107 B.n917 B.n84 585
R108 B.n919 B.n918 585
R109 B.n921 B.n83 585
R110 B.n924 B.n923 585
R111 B.n925 B.n82 585
R112 B.n927 B.n926 585
R113 B.n929 B.n81 585
R114 B.n932 B.n931 585
R115 B.n933 B.n80 585
R116 B.n700 B.n78 585
R117 B.n936 B.n78 585
R118 B.n699 B.n77 585
R119 B.n937 B.n77 585
R120 B.n698 B.n76 585
R121 B.n938 B.n76 585
R122 B.n697 B.n696 585
R123 B.n696 B.n72 585
R124 B.n695 B.n71 585
R125 B.n944 B.n71 585
R126 B.n694 B.n70 585
R127 B.n945 B.n70 585
R128 B.n693 B.n69 585
R129 B.n946 B.n69 585
R130 B.n692 B.n691 585
R131 B.n691 B.n65 585
R132 B.n690 B.n64 585
R133 B.n952 B.n64 585
R134 B.n689 B.n63 585
R135 B.n953 B.n63 585
R136 B.n688 B.n62 585
R137 B.n954 B.n62 585
R138 B.n687 B.n686 585
R139 B.n686 B.n58 585
R140 B.n685 B.n57 585
R141 B.n960 B.n57 585
R142 B.n684 B.n56 585
R143 B.n961 B.n56 585
R144 B.n683 B.n55 585
R145 B.n962 B.n55 585
R146 B.n682 B.n681 585
R147 B.n681 B.n51 585
R148 B.n680 B.n50 585
R149 B.n968 B.n50 585
R150 B.n679 B.n49 585
R151 B.n969 B.n49 585
R152 B.n678 B.n48 585
R153 B.n970 B.n48 585
R154 B.n677 B.n676 585
R155 B.n676 B.n44 585
R156 B.n675 B.n43 585
R157 B.n976 B.n43 585
R158 B.n674 B.n42 585
R159 B.n977 B.n42 585
R160 B.n673 B.n41 585
R161 B.n978 B.n41 585
R162 B.n672 B.n671 585
R163 B.n671 B.n40 585
R164 B.n670 B.n36 585
R165 B.n984 B.n36 585
R166 B.n669 B.n35 585
R167 B.n985 B.n35 585
R168 B.n668 B.n34 585
R169 B.n986 B.n34 585
R170 B.n667 B.n666 585
R171 B.n666 B.n30 585
R172 B.n665 B.n29 585
R173 B.n992 B.n29 585
R174 B.n664 B.n28 585
R175 B.n993 B.n28 585
R176 B.n663 B.n27 585
R177 B.n994 B.n27 585
R178 B.n662 B.n661 585
R179 B.n661 B.n23 585
R180 B.n660 B.n22 585
R181 B.n1000 B.n22 585
R182 B.n659 B.n21 585
R183 B.n1001 B.n21 585
R184 B.n658 B.n20 585
R185 B.n1002 B.n20 585
R186 B.n657 B.n656 585
R187 B.n656 B.n19 585
R188 B.n655 B.n15 585
R189 B.n1008 B.n15 585
R190 B.n654 B.n14 585
R191 B.n1009 B.n14 585
R192 B.n653 B.n13 585
R193 B.n1010 B.n13 585
R194 B.n652 B.n651 585
R195 B.n651 B.n12 585
R196 B.n650 B.n649 585
R197 B.n650 B.n8 585
R198 B.n648 B.n7 585
R199 B.n1017 B.n7 585
R200 B.n647 B.n6 585
R201 B.n1018 B.n6 585
R202 B.n646 B.n5 585
R203 B.n1019 B.n5 585
R204 B.n645 B.n644 585
R205 B.n644 B.n4 585
R206 B.n643 B.n143 585
R207 B.n643 B.n642 585
R208 B.n633 B.n144 585
R209 B.n145 B.n144 585
R210 B.n635 B.n634 585
R211 B.n636 B.n635 585
R212 B.n632 B.n150 585
R213 B.n150 B.n149 585
R214 B.n631 B.n630 585
R215 B.n630 B.n629 585
R216 B.n152 B.n151 585
R217 B.n622 B.n152 585
R218 B.n621 B.n620 585
R219 B.n623 B.n621 585
R220 B.n619 B.n157 585
R221 B.n157 B.n156 585
R222 B.n618 B.n617 585
R223 B.n617 B.n616 585
R224 B.n159 B.n158 585
R225 B.n160 B.n159 585
R226 B.n609 B.n608 585
R227 B.n610 B.n609 585
R228 B.n607 B.n165 585
R229 B.n165 B.n164 585
R230 B.n606 B.n605 585
R231 B.n605 B.n604 585
R232 B.n167 B.n166 585
R233 B.n168 B.n167 585
R234 B.n597 B.n596 585
R235 B.n598 B.n597 585
R236 B.n595 B.n173 585
R237 B.n173 B.n172 585
R238 B.n594 B.n593 585
R239 B.n593 B.n592 585
R240 B.n175 B.n174 585
R241 B.n585 B.n175 585
R242 B.n584 B.n583 585
R243 B.n586 B.n584 585
R244 B.n582 B.n180 585
R245 B.n180 B.n179 585
R246 B.n581 B.n580 585
R247 B.n580 B.n579 585
R248 B.n182 B.n181 585
R249 B.n183 B.n182 585
R250 B.n572 B.n571 585
R251 B.n573 B.n572 585
R252 B.n570 B.n188 585
R253 B.n188 B.n187 585
R254 B.n569 B.n568 585
R255 B.n568 B.n567 585
R256 B.n190 B.n189 585
R257 B.n191 B.n190 585
R258 B.n560 B.n559 585
R259 B.n561 B.n560 585
R260 B.n558 B.n196 585
R261 B.n196 B.n195 585
R262 B.n557 B.n556 585
R263 B.n556 B.n555 585
R264 B.n198 B.n197 585
R265 B.n199 B.n198 585
R266 B.n548 B.n547 585
R267 B.n549 B.n548 585
R268 B.n546 B.n203 585
R269 B.n207 B.n203 585
R270 B.n545 B.n544 585
R271 B.n544 B.n543 585
R272 B.n205 B.n204 585
R273 B.n206 B.n205 585
R274 B.n536 B.n535 585
R275 B.n537 B.n536 585
R276 B.n534 B.n212 585
R277 B.n212 B.n211 585
R278 B.n533 B.n532 585
R279 B.n532 B.n531 585
R280 B.n214 B.n213 585
R281 B.n215 B.n214 585
R282 B.n524 B.n523 585
R283 B.n525 B.n524 585
R284 B.n522 B.n220 585
R285 B.n220 B.n219 585
R286 B.n521 B.n520 585
R287 B.n520 B.n519 585
R288 B.n516 B.n224 585
R289 B.n515 B.n514 585
R290 B.n512 B.n225 585
R291 B.n512 B.n223 585
R292 B.n511 B.n510 585
R293 B.n509 B.n508 585
R294 B.n507 B.n227 585
R295 B.n505 B.n504 585
R296 B.n503 B.n228 585
R297 B.n502 B.n501 585
R298 B.n499 B.n229 585
R299 B.n497 B.n496 585
R300 B.n495 B.n230 585
R301 B.n494 B.n493 585
R302 B.n491 B.n231 585
R303 B.n489 B.n488 585
R304 B.n487 B.n232 585
R305 B.n486 B.n485 585
R306 B.n483 B.n233 585
R307 B.n481 B.n480 585
R308 B.n479 B.n234 585
R309 B.n478 B.n477 585
R310 B.n475 B.n235 585
R311 B.n473 B.n472 585
R312 B.n471 B.n236 585
R313 B.n470 B.n469 585
R314 B.n467 B.n237 585
R315 B.n465 B.n464 585
R316 B.n463 B.n238 585
R317 B.n462 B.n461 585
R318 B.n459 B.n239 585
R319 B.n457 B.n456 585
R320 B.n455 B.n240 585
R321 B.n454 B.n453 585
R322 B.n451 B.n241 585
R323 B.n449 B.n448 585
R324 B.n447 B.n242 585
R325 B.n446 B.n445 585
R326 B.n443 B.n243 585
R327 B.n441 B.n440 585
R328 B.n439 B.n244 585
R329 B.n438 B.n437 585
R330 B.n435 B.n245 585
R331 B.n433 B.n432 585
R332 B.n431 B.n246 585
R333 B.n430 B.n429 585
R334 B.n427 B.n247 585
R335 B.n425 B.n424 585
R336 B.n423 B.n248 585
R337 B.n422 B.n421 585
R338 B.n419 B.n249 585
R339 B.n417 B.n416 585
R340 B.n415 B.n250 585
R341 B.n414 B.n413 585
R342 B.n411 B.n410 585
R343 B.n409 B.n408 585
R344 B.n407 B.n255 585
R345 B.n405 B.n404 585
R346 B.n403 B.n256 585
R347 B.n402 B.n401 585
R348 B.n399 B.n257 585
R349 B.n397 B.n396 585
R350 B.n395 B.n258 585
R351 B.n394 B.n393 585
R352 B.n391 B.n390 585
R353 B.n389 B.n388 585
R354 B.n387 B.n263 585
R355 B.n385 B.n384 585
R356 B.n383 B.n264 585
R357 B.n382 B.n381 585
R358 B.n379 B.n265 585
R359 B.n377 B.n376 585
R360 B.n375 B.n266 585
R361 B.n374 B.n373 585
R362 B.n371 B.n267 585
R363 B.n369 B.n368 585
R364 B.n367 B.n268 585
R365 B.n366 B.n365 585
R366 B.n363 B.n269 585
R367 B.n361 B.n360 585
R368 B.n359 B.n270 585
R369 B.n358 B.n357 585
R370 B.n355 B.n271 585
R371 B.n353 B.n352 585
R372 B.n351 B.n272 585
R373 B.n350 B.n349 585
R374 B.n347 B.n273 585
R375 B.n345 B.n344 585
R376 B.n343 B.n274 585
R377 B.n342 B.n341 585
R378 B.n339 B.n275 585
R379 B.n337 B.n336 585
R380 B.n335 B.n276 585
R381 B.n334 B.n333 585
R382 B.n331 B.n277 585
R383 B.n329 B.n328 585
R384 B.n327 B.n278 585
R385 B.n326 B.n325 585
R386 B.n323 B.n279 585
R387 B.n321 B.n320 585
R388 B.n319 B.n280 585
R389 B.n318 B.n317 585
R390 B.n315 B.n281 585
R391 B.n313 B.n312 585
R392 B.n311 B.n282 585
R393 B.n310 B.n309 585
R394 B.n307 B.n283 585
R395 B.n305 B.n304 585
R396 B.n303 B.n284 585
R397 B.n302 B.n301 585
R398 B.n299 B.n285 585
R399 B.n297 B.n296 585
R400 B.n295 B.n286 585
R401 B.n294 B.n293 585
R402 B.n291 B.n287 585
R403 B.n289 B.n288 585
R404 B.n222 B.n221 585
R405 B.n223 B.n222 585
R406 B.n518 B.n517 585
R407 B.n519 B.n518 585
R408 B.n218 B.n217 585
R409 B.n219 B.n218 585
R410 B.n527 B.n526 585
R411 B.n526 B.n525 585
R412 B.n528 B.n216 585
R413 B.n216 B.n215 585
R414 B.n530 B.n529 585
R415 B.n531 B.n530 585
R416 B.n210 B.n209 585
R417 B.n211 B.n210 585
R418 B.n539 B.n538 585
R419 B.n538 B.n537 585
R420 B.n540 B.n208 585
R421 B.n208 B.n206 585
R422 B.n542 B.n541 585
R423 B.n543 B.n542 585
R424 B.n202 B.n201 585
R425 B.n207 B.n202 585
R426 B.n551 B.n550 585
R427 B.n550 B.n549 585
R428 B.n552 B.n200 585
R429 B.n200 B.n199 585
R430 B.n554 B.n553 585
R431 B.n555 B.n554 585
R432 B.n194 B.n193 585
R433 B.n195 B.n194 585
R434 B.n563 B.n562 585
R435 B.n562 B.n561 585
R436 B.n564 B.n192 585
R437 B.n192 B.n191 585
R438 B.n566 B.n565 585
R439 B.n567 B.n566 585
R440 B.n186 B.n185 585
R441 B.n187 B.n186 585
R442 B.n575 B.n574 585
R443 B.n574 B.n573 585
R444 B.n576 B.n184 585
R445 B.n184 B.n183 585
R446 B.n578 B.n577 585
R447 B.n579 B.n578 585
R448 B.n178 B.n177 585
R449 B.n179 B.n178 585
R450 B.n588 B.n587 585
R451 B.n587 B.n586 585
R452 B.n589 B.n176 585
R453 B.n585 B.n176 585
R454 B.n591 B.n590 585
R455 B.n592 B.n591 585
R456 B.n171 B.n170 585
R457 B.n172 B.n171 585
R458 B.n600 B.n599 585
R459 B.n599 B.n598 585
R460 B.n601 B.n169 585
R461 B.n169 B.n168 585
R462 B.n603 B.n602 585
R463 B.n604 B.n603 585
R464 B.n163 B.n162 585
R465 B.n164 B.n163 585
R466 B.n612 B.n611 585
R467 B.n611 B.n610 585
R468 B.n613 B.n161 585
R469 B.n161 B.n160 585
R470 B.n615 B.n614 585
R471 B.n616 B.n615 585
R472 B.n155 B.n154 585
R473 B.n156 B.n155 585
R474 B.n625 B.n624 585
R475 B.n624 B.n623 585
R476 B.n626 B.n153 585
R477 B.n622 B.n153 585
R478 B.n628 B.n627 585
R479 B.n629 B.n628 585
R480 B.n148 B.n147 585
R481 B.n149 B.n148 585
R482 B.n638 B.n637 585
R483 B.n637 B.n636 585
R484 B.n639 B.n146 585
R485 B.n146 B.n145 585
R486 B.n641 B.n640 585
R487 B.n642 B.n641 585
R488 B.n3 B.n0 585
R489 B.n4 B.n3 585
R490 B.n1016 B.n1 585
R491 B.n1017 B.n1016 585
R492 B.n1015 B.n1014 585
R493 B.n1015 B.n8 585
R494 B.n1013 B.n9 585
R495 B.n12 B.n9 585
R496 B.n1012 B.n1011 585
R497 B.n1011 B.n1010 585
R498 B.n11 B.n10 585
R499 B.n1009 B.n11 585
R500 B.n1007 B.n1006 585
R501 B.n1008 B.n1007 585
R502 B.n1005 B.n16 585
R503 B.n19 B.n16 585
R504 B.n1004 B.n1003 585
R505 B.n1003 B.n1002 585
R506 B.n18 B.n17 585
R507 B.n1001 B.n18 585
R508 B.n999 B.n998 585
R509 B.n1000 B.n999 585
R510 B.n997 B.n24 585
R511 B.n24 B.n23 585
R512 B.n996 B.n995 585
R513 B.n995 B.n994 585
R514 B.n26 B.n25 585
R515 B.n993 B.n26 585
R516 B.n991 B.n990 585
R517 B.n992 B.n991 585
R518 B.n989 B.n31 585
R519 B.n31 B.n30 585
R520 B.n988 B.n987 585
R521 B.n987 B.n986 585
R522 B.n33 B.n32 585
R523 B.n985 B.n33 585
R524 B.n983 B.n982 585
R525 B.n984 B.n983 585
R526 B.n981 B.n37 585
R527 B.n40 B.n37 585
R528 B.n980 B.n979 585
R529 B.n979 B.n978 585
R530 B.n39 B.n38 585
R531 B.n977 B.n39 585
R532 B.n975 B.n974 585
R533 B.n976 B.n975 585
R534 B.n973 B.n45 585
R535 B.n45 B.n44 585
R536 B.n972 B.n971 585
R537 B.n971 B.n970 585
R538 B.n47 B.n46 585
R539 B.n969 B.n47 585
R540 B.n967 B.n966 585
R541 B.n968 B.n967 585
R542 B.n965 B.n52 585
R543 B.n52 B.n51 585
R544 B.n964 B.n963 585
R545 B.n963 B.n962 585
R546 B.n54 B.n53 585
R547 B.n961 B.n54 585
R548 B.n959 B.n958 585
R549 B.n960 B.n959 585
R550 B.n957 B.n59 585
R551 B.n59 B.n58 585
R552 B.n956 B.n955 585
R553 B.n955 B.n954 585
R554 B.n61 B.n60 585
R555 B.n953 B.n61 585
R556 B.n951 B.n950 585
R557 B.n952 B.n951 585
R558 B.n949 B.n66 585
R559 B.n66 B.n65 585
R560 B.n948 B.n947 585
R561 B.n947 B.n946 585
R562 B.n68 B.n67 585
R563 B.n945 B.n68 585
R564 B.n943 B.n942 585
R565 B.n944 B.n943 585
R566 B.n941 B.n73 585
R567 B.n73 B.n72 585
R568 B.n940 B.n939 585
R569 B.n939 B.n938 585
R570 B.n75 B.n74 585
R571 B.n937 B.n75 585
R572 B.n935 B.n934 585
R573 B.n936 B.n935 585
R574 B.n1020 B.n1019 585
R575 B.n1018 B.n2 585
R576 B.n935 B.n80 516.524
R577 B.n702 B.n78 516.524
R578 B.n520 B.n222 516.524
R579 B.n518 B.n224 516.524
R580 B.n107 B.t10 426.173
R581 B.n115 B.t16 426.173
R582 B.n259 B.t14 426.173
R583 B.n251 B.t7 426.173
R584 B.n116 B.t17 350.731
R585 B.n260 B.t13 350.731
R586 B.n108 B.t11 350.731
R587 B.n252 B.t6 350.731
R588 B.n107 B.t8 317.462
R589 B.n115 B.t15 317.462
R590 B.n259 B.t12 317.462
R591 B.n251 B.t4 317.462
R592 B.n703 B.n79 256.663
R593 B.n705 B.n79 256.663
R594 B.n711 B.n79 256.663
R595 B.n713 B.n79 256.663
R596 B.n719 B.n79 256.663
R597 B.n721 B.n79 256.663
R598 B.n727 B.n79 256.663
R599 B.n729 B.n79 256.663
R600 B.n735 B.n79 256.663
R601 B.n737 B.n79 256.663
R602 B.n743 B.n79 256.663
R603 B.n745 B.n79 256.663
R604 B.n751 B.n79 256.663
R605 B.n753 B.n79 256.663
R606 B.n759 B.n79 256.663
R607 B.n761 B.n79 256.663
R608 B.n767 B.n79 256.663
R609 B.n769 B.n79 256.663
R610 B.n775 B.n79 256.663
R611 B.n777 B.n79 256.663
R612 B.n783 B.n79 256.663
R613 B.n785 B.n79 256.663
R614 B.n791 B.n79 256.663
R615 B.n793 B.n79 256.663
R616 B.n799 B.n79 256.663
R617 B.n801 B.n79 256.663
R618 B.n807 B.n79 256.663
R619 B.n809 B.n79 256.663
R620 B.n815 B.n79 256.663
R621 B.n817 B.n79 256.663
R622 B.n823 B.n79 256.663
R623 B.n825 B.n79 256.663
R624 B.n832 B.n79 256.663
R625 B.n834 B.n79 256.663
R626 B.n840 B.n79 256.663
R627 B.n842 B.n79 256.663
R628 B.n848 B.n79 256.663
R629 B.n850 B.n79 256.663
R630 B.n856 B.n79 256.663
R631 B.n858 B.n79 256.663
R632 B.n864 B.n79 256.663
R633 B.n866 B.n79 256.663
R634 B.n872 B.n79 256.663
R635 B.n874 B.n79 256.663
R636 B.n880 B.n79 256.663
R637 B.n882 B.n79 256.663
R638 B.n888 B.n79 256.663
R639 B.n890 B.n79 256.663
R640 B.n896 B.n79 256.663
R641 B.n898 B.n79 256.663
R642 B.n904 B.n79 256.663
R643 B.n906 B.n79 256.663
R644 B.n912 B.n79 256.663
R645 B.n914 B.n79 256.663
R646 B.n920 B.n79 256.663
R647 B.n922 B.n79 256.663
R648 B.n928 B.n79 256.663
R649 B.n930 B.n79 256.663
R650 B.n513 B.n223 256.663
R651 B.n226 B.n223 256.663
R652 B.n506 B.n223 256.663
R653 B.n500 B.n223 256.663
R654 B.n498 B.n223 256.663
R655 B.n492 B.n223 256.663
R656 B.n490 B.n223 256.663
R657 B.n484 B.n223 256.663
R658 B.n482 B.n223 256.663
R659 B.n476 B.n223 256.663
R660 B.n474 B.n223 256.663
R661 B.n468 B.n223 256.663
R662 B.n466 B.n223 256.663
R663 B.n460 B.n223 256.663
R664 B.n458 B.n223 256.663
R665 B.n452 B.n223 256.663
R666 B.n450 B.n223 256.663
R667 B.n444 B.n223 256.663
R668 B.n442 B.n223 256.663
R669 B.n436 B.n223 256.663
R670 B.n434 B.n223 256.663
R671 B.n428 B.n223 256.663
R672 B.n426 B.n223 256.663
R673 B.n420 B.n223 256.663
R674 B.n418 B.n223 256.663
R675 B.n412 B.n223 256.663
R676 B.n254 B.n223 256.663
R677 B.n406 B.n223 256.663
R678 B.n400 B.n223 256.663
R679 B.n398 B.n223 256.663
R680 B.n392 B.n223 256.663
R681 B.n262 B.n223 256.663
R682 B.n386 B.n223 256.663
R683 B.n380 B.n223 256.663
R684 B.n378 B.n223 256.663
R685 B.n372 B.n223 256.663
R686 B.n370 B.n223 256.663
R687 B.n364 B.n223 256.663
R688 B.n362 B.n223 256.663
R689 B.n356 B.n223 256.663
R690 B.n354 B.n223 256.663
R691 B.n348 B.n223 256.663
R692 B.n346 B.n223 256.663
R693 B.n340 B.n223 256.663
R694 B.n338 B.n223 256.663
R695 B.n332 B.n223 256.663
R696 B.n330 B.n223 256.663
R697 B.n324 B.n223 256.663
R698 B.n322 B.n223 256.663
R699 B.n316 B.n223 256.663
R700 B.n314 B.n223 256.663
R701 B.n308 B.n223 256.663
R702 B.n306 B.n223 256.663
R703 B.n300 B.n223 256.663
R704 B.n298 B.n223 256.663
R705 B.n292 B.n223 256.663
R706 B.n290 B.n223 256.663
R707 B.n1022 B.n1021 256.663
R708 B.n931 B.n929 163.367
R709 B.n927 B.n82 163.367
R710 B.n923 B.n921 163.367
R711 B.n919 B.n84 163.367
R712 B.n915 B.n913 163.367
R713 B.n911 B.n86 163.367
R714 B.n907 B.n905 163.367
R715 B.n903 B.n88 163.367
R716 B.n899 B.n897 163.367
R717 B.n895 B.n90 163.367
R718 B.n891 B.n889 163.367
R719 B.n887 B.n92 163.367
R720 B.n883 B.n881 163.367
R721 B.n879 B.n94 163.367
R722 B.n875 B.n873 163.367
R723 B.n871 B.n96 163.367
R724 B.n867 B.n865 163.367
R725 B.n863 B.n98 163.367
R726 B.n859 B.n857 163.367
R727 B.n855 B.n100 163.367
R728 B.n851 B.n849 163.367
R729 B.n847 B.n102 163.367
R730 B.n843 B.n841 163.367
R731 B.n839 B.n104 163.367
R732 B.n835 B.n833 163.367
R733 B.n831 B.n106 163.367
R734 B.n826 B.n824 163.367
R735 B.n822 B.n110 163.367
R736 B.n818 B.n816 163.367
R737 B.n814 B.n112 163.367
R738 B.n810 B.n808 163.367
R739 B.n806 B.n114 163.367
R740 B.n802 B.n800 163.367
R741 B.n798 B.n119 163.367
R742 B.n794 B.n792 163.367
R743 B.n790 B.n121 163.367
R744 B.n786 B.n784 163.367
R745 B.n782 B.n123 163.367
R746 B.n778 B.n776 163.367
R747 B.n774 B.n125 163.367
R748 B.n770 B.n768 163.367
R749 B.n766 B.n127 163.367
R750 B.n762 B.n760 163.367
R751 B.n758 B.n129 163.367
R752 B.n754 B.n752 163.367
R753 B.n750 B.n131 163.367
R754 B.n746 B.n744 163.367
R755 B.n742 B.n133 163.367
R756 B.n738 B.n736 163.367
R757 B.n734 B.n135 163.367
R758 B.n730 B.n728 163.367
R759 B.n726 B.n137 163.367
R760 B.n722 B.n720 163.367
R761 B.n718 B.n139 163.367
R762 B.n714 B.n712 163.367
R763 B.n710 B.n141 163.367
R764 B.n706 B.n704 163.367
R765 B.n520 B.n220 163.367
R766 B.n524 B.n220 163.367
R767 B.n524 B.n214 163.367
R768 B.n532 B.n214 163.367
R769 B.n532 B.n212 163.367
R770 B.n536 B.n212 163.367
R771 B.n536 B.n205 163.367
R772 B.n544 B.n205 163.367
R773 B.n544 B.n203 163.367
R774 B.n548 B.n203 163.367
R775 B.n548 B.n198 163.367
R776 B.n556 B.n198 163.367
R777 B.n556 B.n196 163.367
R778 B.n560 B.n196 163.367
R779 B.n560 B.n190 163.367
R780 B.n568 B.n190 163.367
R781 B.n568 B.n188 163.367
R782 B.n572 B.n188 163.367
R783 B.n572 B.n182 163.367
R784 B.n580 B.n182 163.367
R785 B.n580 B.n180 163.367
R786 B.n584 B.n180 163.367
R787 B.n584 B.n175 163.367
R788 B.n593 B.n175 163.367
R789 B.n593 B.n173 163.367
R790 B.n597 B.n173 163.367
R791 B.n597 B.n167 163.367
R792 B.n605 B.n167 163.367
R793 B.n605 B.n165 163.367
R794 B.n609 B.n165 163.367
R795 B.n609 B.n159 163.367
R796 B.n617 B.n159 163.367
R797 B.n617 B.n157 163.367
R798 B.n621 B.n157 163.367
R799 B.n621 B.n152 163.367
R800 B.n630 B.n152 163.367
R801 B.n630 B.n150 163.367
R802 B.n635 B.n150 163.367
R803 B.n635 B.n144 163.367
R804 B.n643 B.n144 163.367
R805 B.n644 B.n643 163.367
R806 B.n644 B.n5 163.367
R807 B.n6 B.n5 163.367
R808 B.n7 B.n6 163.367
R809 B.n650 B.n7 163.367
R810 B.n651 B.n650 163.367
R811 B.n651 B.n13 163.367
R812 B.n14 B.n13 163.367
R813 B.n15 B.n14 163.367
R814 B.n656 B.n15 163.367
R815 B.n656 B.n20 163.367
R816 B.n21 B.n20 163.367
R817 B.n22 B.n21 163.367
R818 B.n661 B.n22 163.367
R819 B.n661 B.n27 163.367
R820 B.n28 B.n27 163.367
R821 B.n29 B.n28 163.367
R822 B.n666 B.n29 163.367
R823 B.n666 B.n34 163.367
R824 B.n35 B.n34 163.367
R825 B.n36 B.n35 163.367
R826 B.n671 B.n36 163.367
R827 B.n671 B.n41 163.367
R828 B.n42 B.n41 163.367
R829 B.n43 B.n42 163.367
R830 B.n676 B.n43 163.367
R831 B.n676 B.n48 163.367
R832 B.n49 B.n48 163.367
R833 B.n50 B.n49 163.367
R834 B.n681 B.n50 163.367
R835 B.n681 B.n55 163.367
R836 B.n56 B.n55 163.367
R837 B.n57 B.n56 163.367
R838 B.n686 B.n57 163.367
R839 B.n686 B.n62 163.367
R840 B.n63 B.n62 163.367
R841 B.n64 B.n63 163.367
R842 B.n691 B.n64 163.367
R843 B.n691 B.n69 163.367
R844 B.n70 B.n69 163.367
R845 B.n71 B.n70 163.367
R846 B.n696 B.n71 163.367
R847 B.n696 B.n76 163.367
R848 B.n77 B.n76 163.367
R849 B.n78 B.n77 163.367
R850 B.n514 B.n512 163.367
R851 B.n512 B.n511 163.367
R852 B.n508 B.n507 163.367
R853 B.n505 B.n228 163.367
R854 B.n501 B.n499 163.367
R855 B.n497 B.n230 163.367
R856 B.n493 B.n491 163.367
R857 B.n489 B.n232 163.367
R858 B.n485 B.n483 163.367
R859 B.n481 B.n234 163.367
R860 B.n477 B.n475 163.367
R861 B.n473 B.n236 163.367
R862 B.n469 B.n467 163.367
R863 B.n465 B.n238 163.367
R864 B.n461 B.n459 163.367
R865 B.n457 B.n240 163.367
R866 B.n453 B.n451 163.367
R867 B.n449 B.n242 163.367
R868 B.n445 B.n443 163.367
R869 B.n441 B.n244 163.367
R870 B.n437 B.n435 163.367
R871 B.n433 B.n246 163.367
R872 B.n429 B.n427 163.367
R873 B.n425 B.n248 163.367
R874 B.n421 B.n419 163.367
R875 B.n417 B.n250 163.367
R876 B.n413 B.n411 163.367
R877 B.n408 B.n407 163.367
R878 B.n405 B.n256 163.367
R879 B.n401 B.n399 163.367
R880 B.n397 B.n258 163.367
R881 B.n393 B.n391 163.367
R882 B.n388 B.n387 163.367
R883 B.n385 B.n264 163.367
R884 B.n381 B.n379 163.367
R885 B.n377 B.n266 163.367
R886 B.n373 B.n371 163.367
R887 B.n369 B.n268 163.367
R888 B.n365 B.n363 163.367
R889 B.n361 B.n270 163.367
R890 B.n357 B.n355 163.367
R891 B.n353 B.n272 163.367
R892 B.n349 B.n347 163.367
R893 B.n345 B.n274 163.367
R894 B.n341 B.n339 163.367
R895 B.n337 B.n276 163.367
R896 B.n333 B.n331 163.367
R897 B.n329 B.n278 163.367
R898 B.n325 B.n323 163.367
R899 B.n321 B.n280 163.367
R900 B.n317 B.n315 163.367
R901 B.n313 B.n282 163.367
R902 B.n309 B.n307 163.367
R903 B.n305 B.n284 163.367
R904 B.n301 B.n299 163.367
R905 B.n297 B.n286 163.367
R906 B.n293 B.n291 163.367
R907 B.n289 B.n222 163.367
R908 B.n518 B.n218 163.367
R909 B.n526 B.n218 163.367
R910 B.n526 B.n216 163.367
R911 B.n530 B.n216 163.367
R912 B.n530 B.n210 163.367
R913 B.n538 B.n210 163.367
R914 B.n538 B.n208 163.367
R915 B.n542 B.n208 163.367
R916 B.n542 B.n202 163.367
R917 B.n550 B.n202 163.367
R918 B.n550 B.n200 163.367
R919 B.n554 B.n200 163.367
R920 B.n554 B.n194 163.367
R921 B.n562 B.n194 163.367
R922 B.n562 B.n192 163.367
R923 B.n566 B.n192 163.367
R924 B.n566 B.n186 163.367
R925 B.n574 B.n186 163.367
R926 B.n574 B.n184 163.367
R927 B.n578 B.n184 163.367
R928 B.n578 B.n178 163.367
R929 B.n587 B.n178 163.367
R930 B.n587 B.n176 163.367
R931 B.n591 B.n176 163.367
R932 B.n591 B.n171 163.367
R933 B.n599 B.n171 163.367
R934 B.n599 B.n169 163.367
R935 B.n603 B.n169 163.367
R936 B.n603 B.n163 163.367
R937 B.n611 B.n163 163.367
R938 B.n611 B.n161 163.367
R939 B.n615 B.n161 163.367
R940 B.n615 B.n155 163.367
R941 B.n624 B.n155 163.367
R942 B.n624 B.n153 163.367
R943 B.n628 B.n153 163.367
R944 B.n628 B.n148 163.367
R945 B.n637 B.n148 163.367
R946 B.n637 B.n146 163.367
R947 B.n641 B.n146 163.367
R948 B.n641 B.n3 163.367
R949 B.n1020 B.n3 163.367
R950 B.n1016 B.n2 163.367
R951 B.n1016 B.n1015 163.367
R952 B.n1015 B.n9 163.367
R953 B.n1011 B.n9 163.367
R954 B.n1011 B.n11 163.367
R955 B.n1007 B.n11 163.367
R956 B.n1007 B.n16 163.367
R957 B.n1003 B.n16 163.367
R958 B.n1003 B.n18 163.367
R959 B.n999 B.n18 163.367
R960 B.n999 B.n24 163.367
R961 B.n995 B.n24 163.367
R962 B.n995 B.n26 163.367
R963 B.n991 B.n26 163.367
R964 B.n991 B.n31 163.367
R965 B.n987 B.n31 163.367
R966 B.n987 B.n33 163.367
R967 B.n983 B.n33 163.367
R968 B.n983 B.n37 163.367
R969 B.n979 B.n37 163.367
R970 B.n979 B.n39 163.367
R971 B.n975 B.n39 163.367
R972 B.n975 B.n45 163.367
R973 B.n971 B.n45 163.367
R974 B.n971 B.n47 163.367
R975 B.n967 B.n47 163.367
R976 B.n967 B.n52 163.367
R977 B.n963 B.n52 163.367
R978 B.n963 B.n54 163.367
R979 B.n959 B.n54 163.367
R980 B.n959 B.n59 163.367
R981 B.n955 B.n59 163.367
R982 B.n955 B.n61 163.367
R983 B.n951 B.n61 163.367
R984 B.n951 B.n66 163.367
R985 B.n947 B.n66 163.367
R986 B.n947 B.n68 163.367
R987 B.n943 B.n68 163.367
R988 B.n943 B.n73 163.367
R989 B.n939 B.n73 163.367
R990 B.n939 B.n75 163.367
R991 B.n935 B.n75 163.367
R992 B.n108 B.n107 75.4429
R993 B.n116 B.n115 75.4429
R994 B.n260 B.n259 75.4429
R995 B.n252 B.n251 75.4429
R996 B.n930 B.n80 71.676
R997 B.n929 B.n928 71.676
R998 B.n922 B.n82 71.676
R999 B.n921 B.n920 71.676
R1000 B.n914 B.n84 71.676
R1001 B.n913 B.n912 71.676
R1002 B.n906 B.n86 71.676
R1003 B.n905 B.n904 71.676
R1004 B.n898 B.n88 71.676
R1005 B.n897 B.n896 71.676
R1006 B.n890 B.n90 71.676
R1007 B.n889 B.n888 71.676
R1008 B.n882 B.n92 71.676
R1009 B.n881 B.n880 71.676
R1010 B.n874 B.n94 71.676
R1011 B.n873 B.n872 71.676
R1012 B.n866 B.n96 71.676
R1013 B.n865 B.n864 71.676
R1014 B.n858 B.n98 71.676
R1015 B.n857 B.n856 71.676
R1016 B.n850 B.n100 71.676
R1017 B.n849 B.n848 71.676
R1018 B.n842 B.n102 71.676
R1019 B.n841 B.n840 71.676
R1020 B.n834 B.n104 71.676
R1021 B.n833 B.n832 71.676
R1022 B.n825 B.n106 71.676
R1023 B.n824 B.n823 71.676
R1024 B.n817 B.n110 71.676
R1025 B.n816 B.n815 71.676
R1026 B.n809 B.n112 71.676
R1027 B.n808 B.n807 71.676
R1028 B.n801 B.n114 71.676
R1029 B.n800 B.n799 71.676
R1030 B.n793 B.n119 71.676
R1031 B.n792 B.n791 71.676
R1032 B.n785 B.n121 71.676
R1033 B.n784 B.n783 71.676
R1034 B.n777 B.n123 71.676
R1035 B.n776 B.n775 71.676
R1036 B.n769 B.n125 71.676
R1037 B.n768 B.n767 71.676
R1038 B.n761 B.n127 71.676
R1039 B.n760 B.n759 71.676
R1040 B.n753 B.n129 71.676
R1041 B.n752 B.n751 71.676
R1042 B.n745 B.n131 71.676
R1043 B.n744 B.n743 71.676
R1044 B.n737 B.n133 71.676
R1045 B.n736 B.n735 71.676
R1046 B.n729 B.n135 71.676
R1047 B.n728 B.n727 71.676
R1048 B.n721 B.n137 71.676
R1049 B.n720 B.n719 71.676
R1050 B.n713 B.n139 71.676
R1051 B.n712 B.n711 71.676
R1052 B.n705 B.n141 71.676
R1053 B.n704 B.n703 71.676
R1054 B.n703 B.n702 71.676
R1055 B.n706 B.n705 71.676
R1056 B.n711 B.n710 71.676
R1057 B.n714 B.n713 71.676
R1058 B.n719 B.n718 71.676
R1059 B.n722 B.n721 71.676
R1060 B.n727 B.n726 71.676
R1061 B.n730 B.n729 71.676
R1062 B.n735 B.n734 71.676
R1063 B.n738 B.n737 71.676
R1064 B.n743 B.n742 71.676
R1065 B.n746 B.n745 71.676
R1066 B.n751 B.n750 71.676
R1067 B.n754 B.n753 71.676
R1068 B.n759 B.n758 71.676
R1069 B.n762 B.n761 71.676
R1070 B.n767 B.n766 71.676
R1071 B.n770 B.n769 71.676
R1072 B.n775 B.n774 71.676
R1073 B.n778 B.n777 71.676
R1074 B.n783 B.n782 71.676
R1075 B.n786 B.n785 71.676
R1076 B.n791 B.n790 71.676
R1077 B.n794 B.n793 71.676
R1078 B.n799 B.n798 71.676
R1079 B.n802 B.n801 71.676
R1080 B.n807 B.n806 71.676
R1081 B.n810 B.n809 71.676
R1082 B.n815 B.n814 71.676
R1083 B.n818 B.n817 71.676
R1084 B.n823 B.n822 71.676
R1085 B.n826 B.n825 71.676
R1086 B.n832 B.n831 71.676
R1087 B.n835 B.n834 71.676
R1088 B.n840 B.n839 71.676
R1089 B.n843 B.n842 71.676
R1090 B.n848 B.n847 71.676
R1091 B.n851 B.n850 71.676
R1092 B.n856 B.n855 71.676
R1093 B.n859 B.n858 71.676
R1094 B.n864 B.n863 71.676
R1095 B.n867 B.n866 71.676
R1096 B.n872 B.n871 71.676
R1097 B.n875 B.n874 71.676
R1098 B.n880 B.n879 71.676
R1099 B.n883 B.n882 71.676
R1100 B.n888 B.n887 71.676
R1101 B.n891 B.n890 71.676
R1102 B.n896 B.n895 71.676
R1103 B.n899 B.n898 71.676
R1104 B.n904 B.n903 71.676
R1105 B.n907 B.n906 71.676
R1106 B.n912 B.n911 71.676
R1107 B.n915 B.n914 71.676
R1108 B.n920 B.n919 71.676
R1109 B.n923 B.n922 71.676
R1110 B.n928 B.n927 71.676
R1111 B.n931 B.n930 71.676
R1112 B.n513 B.n224 71.676
R1113 B.n511 B.n226 71.676
R1114 B.n507 B.n506 71.676
R1115 B.n500 B.n228 71.676
R1116 B.n499 B.n498 71.676
R1117 B.n492 B.n230 71.676
R1118 B.n491 B.n490 71.676
R1119 B.n484 B.n232 71.676
R1120 B.n483 B.n482 71.676
R1121 B.n476 B.n234 71.676
R1122 B.n475 B.n474 71.676
R1123 B.n468 B.n236 71.676
R1124 B.n467 B.n466 71.676
R1125 B.n460 B.n238 71.676
R1126 B.n459 B.n458 71.676
R1127 B.n452 B.n240 71.676
R1128 B.n451 B.n450 71.676
R1129 B.n444 B.n242 71.676
R1130 B.n443 B.n442 71.676
R1131 B.n436 B.n244 71.676
R1132 B.n435 B.n434 71.676
R1133 B.n428 B.n246 71.676
R1134 B.n427 B.n426 71.676
R1135 B.n420 B.n248 71.676
R1136 B.n419 B.n418 71.676
R1137 B.n412 B.n250 71.676
R1138 B.n411 B.n254 71.676
R1139 B.n407 B.n406 71.676
R1140 B.n400 B.n256 71.676
R1141 B.n399 B.n398 71.676
R1142 B.n392 B.n258 71.676
R1143 B.n391 B.n262 71.676
R1144 B.n387 B.n386 71.676
R1145 B.n380 B.n264 71.676
R1146 B.n379 B.n378 71.676
R1147 B.n372 B.n266 71.676
R1148 B.n371 B.n370 71.676
R1149 B.n364 B.n268 71.676
R1150 B.n363 B.n362 71.676
R1151 B.n356 B.n270 71.676
R1152 B.n355 B.n354 71.676
R1153 B.n348 B.n272 71.676
R1154 B.n347 B.n346 71.676
R1155 B.n340 B.n274 71.676
R1156 B.n339 B.n338 71.676
R1157 B.n332 B.n276 71.676
R1158 B.n331 B.n330 71.676
R1159 B.n324 B.n278 71.676
R1160 B.n323 B.n322 71.676
R1161 B.n316 B.n280 71.676
R1162 B.n315 B.n314 71.676
R1163 B.n308 B.n282 71.676
R1164 B.n307 B.n306 71.676
R1165 B.n300 B.n284 71.676
R1166 B.n299 B.n298 71.676
R1167 B.n292 B.n286 71.676
R1168 B.n291 B.n290 71.676
R1169 B.n514 B.n513 71.676
R1170 B.n508 B.n226 71.676
R1171 B.n506 B.n505 71.676
R1172 B.n501 B.n500 71.676
R1173 B.n498 B.n497 71.676
R1174 B.n493 B.n492 71.676
R1175 B.n490 B.n489 71.676
R1176 B.n485 B.n484 71.676
R1177 B.n482 B.n481 71.676
R1178 B.n477 B.n476 71.676
R1179 B.n474 B.n473 71.676
R1180 B.n469 B.n468 71.676
R1181 B.n466 B.n465 71.676
R1182 B.n461 B.n460 71.676
R1183 B.n458 B.n457 71.676
R1184 B.n453 B.n452 71.676
R1185 B.n450 B.n449 71.676
R1186 B.n445 B.n444 71.676
R1187 B.n442 B.n441 71.676
R1188 B.n437 B.n436 71.676
R1189 B.n434 B.n433 71.676
R1190 B.n429 B.n428 71.676
R1191 B.n426 B.n425 71.676
R1192 B.n421 B.n420 71.676
R1193 B.n418 B.n417 71.676
R1194 B.n413 B.n412 71.676
R1195 B.n408 B.n254 71.676
R1196 B.n406 B.n405 71.676
R1197 B.n401 B.n400 71.676
R1198 B.n398 B.n397 71.676
R1199 B.n393 B.n392 71.676
R1200 B.n388 B.n262 71.676
R1201 B.n386 B.n385 71.676
R1202 B.n381 B.n380 71.676
R1203 B.n378 B.n377 71.676
R1204 B.n373 B.n372 71.676
R1205 B.n370 B.n369 71.676
R1206 B.n365 B.n364 71.676
R1207 B.n362 B.n361 71.676
R1208 B.n357 B.n356 71.676
R1209 B.n354 B.n353 71.676
R1210 B.n349 B.n348 71.676
R1211 B.n346 B.n345 71.676
R1212 B.n341 B.n340 71.676
R1213 B.n338 B.n337 71.676
R1214 B.n333 B.n332 71.676
R1215 B.n330 B.n329 71.676
R1216 B.n325 B.n324 71.676
R1217 B.n322 B.n321 71.676
R1218 B.n317 B.n316 71.676
R1219 B.n314 B.n313 71.676
R1220 B.n309 B.n308 71.676
R1221 B.n306 B.n305 71.676
R1222 B.n301 B.n300 71.676
R1223 B.n298 B.n297 71.676
R1224 B.n293 B.n292 71.676
R1225 B.n290 B.n289 71.676
R1226 B.n1021 B.n1020 71.676
R1227 B.n1021 B.n2 71.676
R1228 B.n519 B.n223 61.5281
R1229 B.n936 B.n79 61.5281
R1230 B.n828 B.n108 59.5399
R1231 B.n117 B.n116 59.5399
R1232 B.n261 B.n260 59.5399
R1233 B.n253 B.n252 59.5399
R1234 B.n519 B.n219 35.1591
R1235 B.n525 B.n219 35.1591
R1236 B.n525 B.n215 35.1591
R1237 B.n531 B.n215 35.1591
R1238 B.n531 B.n211 35.1591
R1239 B.n537 B.n211 35.1591
R1240 B.n537 B.n206 35.1591
R1241 B.n543 B.n206 35.1591
R1242 B.n543 B.n207 35.1591
R1243 B.n549 B.n199 35.1591
R1244 B.n555 B.n199 35.1591
R1245 B.n555 B.n195 35.1591
R1246 B.n561 B.n195 35.1591
R1247 B.n561 B.n191 35.1591
R1248 B.n567 B.n191 35.1591
R1249 B.n567 B.n187 35.1591
R1250 B.n573 B.n187 35.1591
R1251 B.n573 B.n183 35.1591
R1252 B.n579 B.n183 35.1591
R1253 B.n579 B.n179 35.1591
R1254 B.n586 B.n179 35.1591
R1255 B.n586 B.n585 35.1591
R1256 B.n592 B.n172 35.1591
R1257 B.n598 B.n172 35.1591
R1258 B.n598 B.n168 35.1591
R1259 B.n604 B.n168 35.1591
R1260 B.n604 B.n164 35.1591
R1261 B.n610 B.n164 35.1591
R1262 B.n610 B.n160 35.1591
R1263 B.n616 B.n160 35.1591
R1264 B.n616 B.n156 35.1591
R1265 B.n623 B.n156 35.1591
R1266 B.n623 B.n622 35.1591
R1267 B.n629 B.n149 35.1591
R1268 B.n636 B.n149 35.1591
R1269 B.n636 B.n145 35.1591
R1270 B.n642 B.n145 35.1591
R1271 B.n642 B.n4 35.1591
R1272 B.n1019 B.n4 35.1591
R1273 B.n1019 B.n1018 35.1591
R1274 B.n1018 B.n1017 35.1591
R1275 B.n1017 B.n8 35.1591
R1276 B.n12 B.n8 35.1591
R1277 B.n1010 B.n12 35.1591
R1278 B.n1010 B.n1009 35.1591
R1279 B.n1009 B.n1008 35.1591
R1280 B.n1002 B.n19 35.1591
R1281 B.n1002 B.n1001 35.1591
R1282 B.n1001 B.n1000 35.1591
R1283 B.n1000 B.n23 35.1591
R1284 B.n994 B.n23 35.1591
R1285 B.n994 B.n993 35.1591
R1286 B.n993 B.n992 35.1591
R1287 B.n992 B.n30 35.1591
R1288 B.n986 B.n30 35.1591
R1289 B.n986 B.n985 35.1591
R1290 B.n985 B.n984 35.1591
R1291 B.n978 B.n40 35.1591
R1292 B.n978 B.n977 35.1591
R1293 B.n977 B.n976 35.1591
R1294 B.n976 B.n44 35.1591
R1295 B.n970 B.n44 35.1591
R1296 B.n970 B.n969 35.1591
R1297 B.n969 B.n968 35.1591
R1298 B.n968 B.n51 35.1591
R1299 B.n962 B.n51 35.1591
R1300 B.n962 B.n961 35.1591
R1301 B.n961 B.n960 35.1591
R1302 B.n960 B.n58 35.1591
R1303 B.n954 B.n58 35.1591
R1304 B.n953 B.n952 35.1591
R1305 B.n952 B.n65 35.1591
R1306 B.n946 B.n65 35.1591
R1307 B.n946 B.n945 35.1591
R1308 B.n945 B.n944 35.1591
R1309 B.n944 B.n72 35.1591
R1310 B.n938 B.n72 35.1591
R1311 B.n938 B.n937 35.1591
R1312 B.n937 B.n936 35.1591
R1313 B.n517 B.n516 33.5615
R1314 B.n521 B.n221 33.5615
R1315 B.n701 B.n700 33.5615
R1316 B.n934 B.n933 33.5615
R1317 B.n549 B.t5 32.0569
R1318 B.n954 B.t9 32.0569
R1319 B.n629 B.t3 28.9547
R1320 B.n1008 B.t0 28.9547
R1321 B.n585 B.t1 25.8524
R1322 B.n40 B.t2 25.8524
R1323 B B.n1022 18.0485
R1324 B.n517 B.n217 10.6151
R1325 B.n527 B.n217 10.6151
R1326 B.n528 B.n527 10.6151
R1327 B.n529 B.n528 10.6151
R1328 B.n529 B.n209 10.6151
R1329 B.n539 B.n209 10.6151
R1330 B.n540 B.n539 10.6151
R1331 B.n541 B.n540 10.6151
R1332 B.n541 B.n201 10.6151
R1333 B.n551 B.n201 10.6151
R1334 B.n552 B.n551 10.6151
R1335 B.n553 B.n552 10.6151
R1336 B.n553 B.n193 10.6151
R1337 B.n563 B.n193 10.6151
R1338 B.n564 B.n563 10.6151
R1339 B.n565 B.n564 10.6151
R1340 B.n565 B.n185 10.6151
R1341 B.n575 B.n185 10.6151
R1342 B.n576 B.n575 10.6151
R1343 B.n577 B.n576 10.6151
R1344 B.n577 B.n177 10.6151
R1345 B.n588 B.n177 10.6151
R1346 B.n589 B.n588 10.6151
R1347 B.n590 B.n589 10.6151
R1348 B.n590 B.n170 10.6151
R1349 B.n600 B.n170 10.6151
R1350 B.n601 B.n600 10.6151
R1351 B.n602 B.n601 10.6151
R1352 B.n602 B.n162 10.6151
R1353 B.n612 B.n162 10.6151
R1354 B.n613 B.n612 10.6151
R1355 B.n614 B.n613 10.6151
R1356 B.n614 B.n154 10.6151
R1357 B.n625 B.n154 10.6151
R1358 B.n626 B.n625 10.6151
R1359 B.n627 B.n626 10.6151
R1360 B.n627 B.n147 10.6151
R1361 B.n638 B.n147 10.6151
R1362 B.n639 B.n638 10.6151
R1363 B.n640 B.n639 10.6151
R1364 B.n640 B.n0 10.6151
R1365 B.n516 B.n515 10.6151
R1366 B.n515 B.n225 10.6151
R1367 B.n510 B.n225 10.6151
R1368 B.n510 B.n509 10.6151
R1369 B.n509 B.n227 10.6151
R1370 B.n504 B.n227 10.6151
R1371 B.n504 B.n503 10.6151
R1372 B.n503 B.n502 10.6151
R1373 B.n502 B.n229 10.6151
R1374 B.n496 B.n229 10.6151
R1375 B.n496 B.n495 10.6151
R1376 B.n495 B.n494 10.6151
R1377 B.n494 B.n231 10.6151
R1378 B.n488 B.n231 10.6151
R1379 B.n488 B.n487 10.6151
R1380 B.n487 B.n486 10.6151
R1381 B.n486 B.n233 10.6151
R1382 B.n480 B.n233 10.6151
R1383 B.n480 B.n479 10.6151
R1384 B.n479 B.n478 10.6151
R1385 B.n478 B.n235 10.6151
R1386 B.n472 B.n235 10.6151
R1387 B.n472 B.n471 10.6151
R1388 B.n471 B.n470 10.6151
R1389 B.n470 B.n237 10.6151
R1390 B.n464 B.n237 10.6151
R1391 B.n464 B.n463 10.6151
R1392 B.n463 B.n462 10.6151
R1393 B.n462 B.n239 10.6151
R1394 B.n456 B.n239 10.6151
R1395 B.n456 B.n455 10.6151
R1396 B.n455 B.n454 10.6151
R1397 B.n454 B.n241 10.6151
R1398 B.n448 B.n241 10.6151
R1399 B.n448 B.n447 10.6151
R1400 B.n447 B.n446 10.6151
R1401 B.n446 B.n243 10.6151
R1402 B.n440 B.n243 10.6151
R1403 B.n440 B.n439 10.6151
R1404 B.n439 B.n438 10.6151
R1405 B.n438 B.n245 10.6151
R1406 B.n432 B.n245 10.6151
R1407 B.n432 B.n431 10.6151
R1408 B.n431 B.n430 10.6151
R1409 B.n430 B.n247 10.6151
R1410 B.n424 B.n247 10.6151
R1411 B.n424 B.n423 10.6151
R1412 B.n423 B.n422 10.6151
R1413 B.n422 B.n249 10.6151
R1414 B.n416 B.n249 10.6151
R1415 B.n416 B.n415 10.6151
R1416 B.n415 B.n414 10.6151
R1417 B.n410 B.n409 10.6151
R1418 B.n409 B.n255 10.6151
R1419 B.n404 B.n255 10.6151
R1420 B.n404 B.n403 10.6151
R1421 B.n403 B.n402 10.6151
R1422 B.n402 B.n257 10.6151
R1423 B.n396 B.n257 10.6151
R1424 B.n396 B.n395 10.6151
R1425 B.n395 B.n394 10.6151
R1426 B.n390 B.n389 10.6151
R1427 B.n389 B.n263 10.6151
R1428 B.n384 B.n263 10.6151
R1429 B.n384 B.n383 10.6151
R1430 B.n383 B.n382 10.6151
R1431 B.n382 B.n265 10.6151
R1432 B.n376 B.n265 10.6151
R1433 B.n376 B.n375 10.6151
R1434 B.n375 B.n374 10.6151
R1435 B.n374 B.n267 10.6151
R1436 B.n368 B.n267 10.6151
R1437 B.n368 B.n367 10.6151
R1438 B.n367 B.n366 10.6151
R1439 B.n366 B.n269 10.6151
R1440 B.n360 B.n269 10.6151
R1441 B.n360 B.n359 10.6151
R1442 B.n359 B.n358 10.6151
R1443 B.n358 B.n271 10.6151
R1444 B.n352 B.n271 10.6151
R1445 B.n352 B.n351 10.6151
R1446 B.n351 B.n350 10.6151
R1447 B.n350 B.n273 10.6151
R1448 B.n344 B.n273 10.6151
R1449 B.n344 B.n343 10.6151
R1450 B.n343 B.n342 10.6151
R1451 B.n342 B.n275 10.6151
R1452 B.n336 B.n275 10.6151
R1453 B.n336 B.n335 10.6151
R1454 B.n335 B.n334 10.6151
R1455 B.n334 B.n277 10.6151
R1456 B.n328 B.n277 10.6151
R1457 B.n328 B.n327 10.6151
R1458 B.n327 B.n326 10.6151
R1459 B.n326 B.n279 10.6151
R1460 B.n320 B.n279 10.6151
R1461 B.n320 B.n319 10.6151
R1462 B.n319 B.n318 10.6151
R1463 B.n318 B.n281 10.6151
R1464 B.n312 B.n281 10.6151
R1465 B.n312 B.n311 10.6151
R1466 B.n311 B.n310 10.6151
R1467 B.n310 B.n283 10.6151
R1468 B.n304 B.n283 10.6151
R1469 B.n304 B.n303 10.6151
R1470 B.n303 B.n302 10.6151
R1471 B.n302 B.n285 10.6151
R1472 B.n296 B.n285 10.6151
R1473 B.n296 B.n295 10.6151
R1474 B.n295 B.n294 10.6151
R1475 B.n294 B.n287 10.6151
R1476 B.n288 B.n287 10.6151
R1477 B.n288 B.n221 10.6151
R1478 B.n522 B.n521 10.6151
R1479 B.n523 B.n522 10.6151
R1480 B.n523 B.n213 10.6151
R1481 B.n533 B.n213 10.6151
R1482 B.n534 B.n533 10.6151
R1483 B.n535 B.n534 10.6151
R1484 B.n535 B.n204 10.6151
R1485 B.n545 B.n204 10.6151
R1486 B.n546 B.n545 10.6151
R1487 B.n547 B.n546 10.6151
R1488 B.n547 B.n197 10.6151
R1489 B.n557 B.n197 10.6151
R1490 B.n558 B.n557 10.6151
R1491 B.n559 B.n558 10.6151
R1492 B.n559 B.n189 10.6151
R1493 B.n569 B.n189 10.6151
R1494 B.n570 B.n569 10.6151
R1495 B.n571 B.n570 10.6151
R1496 B.n571 B.n181 10.6151
R1497 B.n581 B.n181 10.6151
R1498 B.n582 B.n581 10.6151
R1499 B.n583 B.n582 10.6151
R1500 B.n583 B.n174 10.6151
R1501 B.n594 B.n174 10.6151
R1502 B.n595 B.n594 10.6151
R1503 B.n596 B.n595 10.6151
R1504 B.n596 B.n166 10.6151
R1505 B.n606 B.n166 10.6151
R1506 B.n607 B.n606 10.6151
R1507 B.n608 B.n607 10.6151
R1508 B.n608 B.n158 10.6151
R1509 B.n618 B.n158 10.6151
R1510 B.n619 B.n618 10.6151
R1511 B.n620 B.n619 10.6151
R1512 B.n620 B.n151 10.6151
R1513 B.n631 B.n151 10.6151
R1514 B.n632 B.n631 10.6151
R1515 B.n634 B.n632 10.6151
R1516 B.n634 B.n633 10.6151
R1517 B.n633 B.n143 10.6151
R1518 B.n645 B.n143 10.6151
R1519 B.n646 B.n645 10.6151
R1520 B.n647 B.n646 10.6151
R1521 B.n648 B.n647 10.6151
R1522 B.n649 B.n648 10.6151
R1523 B.n652 B.n649 10.6151
R1524 B.n653 B.n652 10.6151
R1525 B.n654 B.n653 10.6151
R1526 B.n655 B.n654 10.6151
R1527 B.n657 B.n655 10.6151
R1528 B.n658 B.n657 10.6151
R1529 B.n659 B.n658 10.6151
R1530 B.n660 B.n659 10.6151
R1531 B.n662 B.n660 10.6151
R1532 B.n663 B.n662 10.6151
R1533 B.n664 B.n663 10.6151
R1534 B.n665 B.n664 10.6151
R1535 B.n667 B.n665 10.6151
R1536 B.n668 B.n667 10.6151
R1537 B.n669 B.n668 10.6151
R1538 B.n670 B.n669 10.6151
R1539 B.n672 B.n670 10.6151
R1540 B.n673 B.n672 10.6151
R1541 B.n674 B.n673 10.6151
R1542 B.n675 B.n674 10.6151
R1543 B.n677 B.n675 10.6151
R1544 B.n678 B.n677 10.6151
R1545 B.n679 B.n678 10.6151
R1546 B.n680 B.n679 10.6151
R1547 B.n682 B.n680 10.6151
R1548 B.n683 B.n682 10.6151
R1549 B.n684 B.n683 10.6151
R1550 B.n685 B.n684 10.6151
R1551 B.n687 B.n685 10.6151
R1552 B.n688 B.n687 10.6151
R1553 B.n689 B.n688 10.6151
R1554 B.n690 B.n689 10.6151
R1555 B.n692 B.n690 10.6151
R1556 B.n693 B.n692 10.6151
R1557 B.n694 B.n693 10.6151
R1558 B.n695 B.n694 10.6151
R1559 B.n697 B.n695 10.6151
R1560 B.n698 B.n697 10.6151
R1561 B.n699 B.n698 10.6151
R1562 B.n700 B.n699 10.6151
R1563 B.n1014 B.n1 10.6151
R1564 B.n1014 B.n1013 10.6151
R1565 B.n1013 B.n1012 10.6151
R1566 B.n1012 B.n10 10.6151
R1567 B.n1006 B.n10 10.6151
R1568 B.n1006 B.n1005 10.6151
R1569 B.n1005 B.n1004 10.6151
R1570 B.n1004 B.n17 10.6151
R1571 B.n998 B.n17 10.6151
R1572 B.n998 B.n997 10.6151
R1573 B.n997 B.n996 10.6151
R1574 B.n996 B.n25 10.6151
R1575 B.n990 B.n25 10.6151
R1576 B.n990 B.n989 10.6151
R1577 B.n989 B.n988 10.6151
R1578 B.n988 B.n32 10.6151
R1579 B.n982 B.n32 10.6151
R1580 B.n982 B.n981 10.6151
R1581 B.n981 B.n980 10.6151
R1582 B.n980 B.n38 10.6151
R1583 B.n974 B.n38 10.6151
R1584 B.n974 B.n973 10.6151
R1585 B.n973 B.n972 10.6151
R1586 B.n972 B.n46 10.6151
R1587 B.n966 B.n46 10.6151
R1588 B.n966 B.n965 10.6151
R1589 B.n965 B.n964 10.6151
R1590 B.n964 B.n53 10.6151
R1591 B.n958 B.n53 10.6151
R1592 B.n958 B.n957 10.6151
R1593 B.n957 B.n956 10.6151
R1594 B.n956 B.n60 10.6151
R1595 B.n950 B.n60 10.6151
R1596 B.n950 B.n949 10.6151
R1597 B.n949 B.n948 10.6151
R1598 B.n948 B.n67 10.6151
R1599 B.n942 B.n67 10.6151
R1600 B.n942 B.n941 10.6151
R1601 B.n941 B.n940 10.6151
R1602 B.n940 B.n74 10.6151
R1603 B.n934 B.n74 10.6151
R1604 B.n933 B.n932 10.6151
R1605 B.n932 B.n81 10.6151
R1606 B.n926 B.n81 10.6151
R1607 B.n926 B.n925 10.6151
R1608 B.n925 B.n924 10.6151
R1609 B.n924 B.n83 10.6151
R1610 B.n918 B.n83 10.6151
R1611 B.n918 B.n917 10.6151
R1612 B.n917 B.n916 10.6151
R1613 B.n916 B.n85 10.6151
R1614 B.n910 B.n85 10.6151
R1615 B.n910 B.n909 10.6151
R1616 B.n909 B.n908 10.6151
R1617 B.n908 B.n87 10.6151
R1618 B.n902 B.n87 10.6151
R1619 B.n902 B.n901 10.6151
R1620 B.n901 B.n900 10.6151
R1621 B.n900 B.n89 10.6151
R1622 B.n894 B.n89 10.6151
R1623 B.n894 B.n893 10.6151
R1624 B.n893 B.n892 10.6151
R1625 B.n892 B.n91 10.6151
R1626 B.n886 B.n91 10.6151
R1627 B.n886 B.n885 10.6151
R1628 B.n885 B.n884 10.6151
R1629 B.n884 B.n93 10.6151
R1630 B.n878 B.n93 10.6151
R1631 B.n878 B.n877 10.6151
R1632 B.n877 B.n876 10.6151
R1633 B.n876 B.n95 10.6151
R1634 B.n870 B.n95 10.6151
R1635 B.n870 B.n869 10.6151
R1636 B.n869 B.n868 10.6151
R1637 B.n868 B.n97 10.6151
R1638 B.n862 B.n97 10.6151
R1639 B.n862 B.n861 10.6151
R1640 B.n861 B.n860 10.6151
R1641 B.n860 B.n99 10.6151
R1642 B.n854 B.n99 10.6151
R1643 B.n854 B.n853 10.6151
R1644 B.n853 B.n852 10.6151
R1645 B.n852 B.n101 10.6151
R1646 B.n846 B.n101 10.6151
R1647 B.n846 B.n845 10.6151
R1648 B.n845 B.n844 10.6151
R1649 B.n844 B.n103 10.6151
R1650 B.n838 B.n103 10.6151
R1651 B.n838 B.n837 10.6151
R1652 B.n837 B.n836 10.6151
R1653 B.n836 B.n105 10.6151
R1654 B.n830 B.n105 10.6151
R1655 B.n830 B.n829 10.6151
R1656 B.n827 B.n109 10.6151
R1657 B.n821 B.n109 10.6151
R1658 B.n821 B.n820 10.6151
R1659 B.n820 B.n819 10.6151
R1660 B.n819 B.n111 10.6151
R1661 B.n813 B.n111 10.6151
R1662 B.n813 B.n812 10.6151
R1663 B.n812 B.n811 10.6151
R1664 B.n811 B.n113 10.6151
R1665 B.n805 B.n804 10.6151
R1666 B.n804 B.n803 10.6151
R1667 B.n803 B.n118 10.6151
R1668 B.n797 B.n118 10.6151
R1669 B.n797 B.n796 10.6151
R1670 B.n796 B.n795 10.6151
R1671 B.n795 B.n120 10.6151
R1672 B.n789 B.n120 10.6151
R1673 B.n789 B.n788 10.6151
R1674 B.n788 B.n787 10.6151
R1675 B.n787 B.n122 10.6151
R1676 B.n781 B.n122 10.6151
R1677 B.n781 B.n780 10.6151
R1678 B.n780 B.n779 10.6151
R1679 B.n779 B.n124 10.6151
R1680 B.n773 B.n124 10.6151
R1681 B.n773 B.n772 10.6151
R1682 B.n772 B.n771 10.6151
R1683 B.n771 B.n126 10.6151
R1684 B.n765 B.n126 10.6151
R1685 B.n765 B.n764 10.6151
R1686 B.n764 B.n763 10.6151
R1687 B.n763 B.n128 10.6151
R1688 B.n757 B.n128 10.6151
R1689 B.n757 B.n756 10.6151
R1690 B.n756 B.n755 10.6151
R1691 B.n755 B.n130 10.6151
R1692 B.n749 B.n130 10.6151
R1693 B.n749 B.n748 10.6151
R1694 B.n748 B.n747 10.6151
R1695 B.n747 B.n132 10.6151
R1696 B.n741 B.n132 10.6151
R1697 B.n741 B.n740 10.6151
R1698 B.n740 B.n739 10.6151
R1699 B.n739 B.n134 10.6151
R1700 B.n733 B.n134 10.6151
R1701 B.n733 B.n732 10.6151
R1702 B.n732 B.n731 10.6151
R1703 B.n731 B.n136 10.6151
R1704 B.n725 B.n136 10.6151
R1705 B.n725 B.n724 10.6151
R1706 B.n724 B.n723 10.6151
R1707 B.n723 B.n138 10.6151
R1708 B.n717 B.n138 10.6151
R1709 B.n717 B.n716 10.6151
R1710 B.n716 B.n715 10.6151
R1711 B.n715 B.n140 10.6151
R1712 B.n709 B.n140 10.6151
R1713 B.n709 B.n708 10.6151
R1714 B.n708 B.n707 10.6151
R1715 B.n707 B.n142 10.6151
R1716 B.n701 B.n142 10.6151
R1717 B.n414 B.n253 9.36635
R1718 B.n390 B.n261 9.36635
R1719 B.n829 B.n828 9.36635
R1720 B.n805 B.n117 9.36635
R1721 B.n592 B.t1 9.3072
R1722 B.n984 B.t2 9.3072
R1723 B.n1022 B.n0 8.11757
R1724 B.n1022 B.n1 8.11757
R1725 B.n622 B.t3 6.20497
R1726 B.n19 B.t0 6.20497
R1727 B.n207 B.t5 3.10273
R1728 B.t9 B.n953 3.10273
R1729 B.n410 B.n253 1.24928
R1730 B.n394 B.n261 1.24928
R1731 B.n828 B.n827 1.24928
R1732 B.n117 B.n113 1.24928
R1733 VP.n19 VP.n18 161.3
R1734 VP.n17 VP.n1 161.3
R1735 VP.n16 VP.n15 161.3
R1736 VP.n14 VP.n2 161.3
R1737 VP.n13 VP.n12 161.3
R1738 VP.n11 VP.n3 161.3
R1739 VP.n10 VP.n9 161.3
R1740 VP.n8 VP.n4 161.3
R1741 VP.n5 VP.t2 143.103
R1742 VP.n5 VP.t0 141.869
R1743 VP.n6 VP.t3 108.316
R1744 VP.n0 VP.t1 108.316
R1745 VP.n7 VP.n6 80.6547
R1746 VP.n20 VP.n0 80.6547
R1747 VP.n12 VP.n2 56.5617
R1748 VP.n7 VP.n5 54.4854
R1749 VP.n10 VP.n4 24.5923
R1750 VP.n11 VP.n10 24.5923
R1751 VP.n12 VP.n11 24.5923
R1752 VP.n16 VP.n2 24.5923
R1753 VP.n17 VP.n16 24.5923
R1754 VP.n18 VP.n17 24.5923
R1755 VP.n6 VP.n4 9.59132
R1756 VP.n18 VP.n0 9.59132
R1757 VP.n8 VP.n7 0.354861
R1758 VP.n20 VP.n19 0.354861
R1759 VP VP.n20 0.267071
R1760 VP.n9 VP.n8 0.189894
R1761 VP.n9 VP.n3 0.189894
R1762 VP.n13 VP.n3 0.189894
R1763 VP.n14 VP.n13 0.189894
R1764 VP.n15 VP.n14 0.189894
R1765 VP.n15 VP.n1 0.189894
R1766 VP.n19 VP.n1 0.189894
R1767 VTAIL.n714 VTAIL.n630 289.615
R1768 VTAIL.n84 VTAIL.n0 289.615
R1769 VTAIL.n174 VTAIL.n90 289.615
R1770 VTAIL.n264 VTAIL.n180 289.615
R1771 VTAIL.n624 VTAIL.n540 289.615
R1772 VTAIL.n534 VTAIL.n450 289.615
R1773 VTAIL.n444 VTAIL.n360 289.615
R1774 VTAIL.n354 VTAIL.n270 289.615
R1775 VTAIL.n658 VTAIL.n657 185
R1776 VTAIL.n663 VTAIL.n662 185
R1777 VTAIL.n665 VTAIL.n664 185
R1778 VTAIL.n654 VTAIL.n653 185
R1779 VTAIL.n671 VTAIL.n670 185
R1780 VTAIL.n673 VTAIL.n672 185
R1781 VTAIL.n650 VTAIL.n649 185
R1782 VTAIL.n679 VTAIL.n678 185
R1783 VTAIL.n681 VTAIL.n680 185
R1784 VTAIL.n646 VTAIL.n645 185
R1785 VTAIL.n687 VTAIL.n686 185
R1786 VTAIL.n689 VTAIL.n688 185
R1787 VTAIL.n642 VTAIL.n641 185
R1788 VTAIL.n695 VTAIL.n694 185
R1789 VTAIL.n697 VTAIL.n696 185
R1790 VTAIL.n638 VTAIL.n637 185
R1791 VTAIL.n704 VTAIL.n703 185
R1792 VTAIL.n705 VTAIL.n636 185
R1793 VTAIL.n707 VTAIL.n706 185
R1794 VTAIL.n634 VTAIL.n633 185
R1795 VTAIL.n713 VTAIL.n712 185
R1796 VTAIL.n715 VTAIL.n714 185
R1797 VTAIL.n28 VTAIL.n27 185
R1798 VTAIL.n33 VTAIL.n32 185
R1799 VTAIL.n35 VTAIL.n34 185
R1800 VTAIL.n24 VTAIL.n23 185
R1801 VTAIL.n41 VTAIL.n40 185
R1802 VTAIL.n43 VTAIL.n42 185
R1803 VTAIL.n20 VTAIL.n19 185
R1804 VTAIL.n49 VTAIL.n48 185
R1805 VTAIL.n51 VTAIL.n50 185
R1806 VTAIL.n16 VTAIL.n15 185
R1807 VTAIL.n57 VTAIL.n56 185
R1808 VTAIL.n59 VTAIL.n58 185
R1809 VTAIL.n12 VTAIL.n11 185
R1810 VTAIL.n65 VTAIL.n64 185
R1811 VTAIL.n67 VTAIL.n66 185
R1812 VTAIL.n8 VTAIL.n7 185
R1813 VTAIL.n74 VTAIL.n73 185
R1814 VTAIL.n75 VTAIL.n6 185
R1815 VTAIL.n77 VTAIL.n76 185
R1816 VTAIL.n4 VTAIL.n3 185
R1817 VTAIL.n83 VTAIL.n82 185
R1818 VTAIL.n85 VTAIL.n84 185
R1819 VTAIL.n118 VTAIL.n117 185
R1820 VTAIL.n123 VTAIL.n122 185
R1821 VTAIL.n125 VTAIL.n124 185
R1822 VTAIL.n114 VTAIL.n113 185
R1823 VTAIL.n131 VTAIL.n130 185
R1824 VTAIL.n133 VTAIL.n132 185
R1825 VTAIL.n110 VTAIL.n109 185
R1826 VTAIL.n139 VTAIL.n138 185
R1827 VTAIL.n141 VTAIL.n140 185
R1828 VTAIL.n106 VTAIL.n105 185
R1829 VTAIL.n147 VTAIL.n146 185
R1830 VTAIL.n149 VTAIL.n148 185
R1831 VTAIL.n102 VTAIL.n101 185
R1832 VTAIL.n155 VTAIL.n154 185
R1833 VTAIL.n157 VTAIL.n156 185
R1834 VTAIL.n98 VTAIL.n97 185
R1835 VTAIL.n164 VTAIL.n163 185
R1836 VTAIL.n165 VTAIL.n96 185
R1837 VTAIL.n167 VTAIL.n166 185
R1838 VTAIL.n94 VTAIL.n93 185
R1839 VTAIL.n173 VTAIL.n172 185
R1840 VTAIL.n175 VTAIL.n174 185
R1841 VTAIL.n208 VTAIL.n207 185
R1842 VTAIL.n213 VTAIL.n212 185
R1843 VTAIL.n215 VTAIL.n214 185
R1844 VTAIL.n204 VTAIL.n203 185
R1845 VTAIL.n221 VTAIL.n220 185
R1846 VTAIL.n223 VTAIL.n222 185
R1847 VTAIL.n200 VTAIL.n199 185
R1848 VTAIL.n229 VTAIL.n228 185
R1849 VTAIL.n231 VTAIL.n230 185
R1850 VTAIL.n196 VTAIL.n195 185
R1851 VTAIL.n237 VTAIL.n236 185
R1852 VTAIL.n239 VTAIL.n238 185
R1853 VTAIL.n192 VTAIL.n191 185
R1854 VTAIL.n245 VTAIL.n244 185
R1855 VTAIL.n247 VTAIL.n246 185
R1856 VTAIL.n188 VTAIL.n187 185
R1857 VTAIL.n254 VTAIL.n253 185
R1858 VTAIL.n255 VTAIL.n186 185
R1859 VTAIL.n257 VTAIL.n256 185
R1860 VTAIL.n184 VTAIL.n183 185
R1861 VTAIL.n263 VTAIL.n262 185
R1862 VTAIL.n265 VTAIL.n264 185
R1863 VTAIL.n625 VTAIL.n624 185
R1864 VTAIL.n623 VTAIL.n622 185
R1865 VTAIL.n544 VTAIL.n543 185
R1866 VTAIL.n617 VTAIL.n616 185
R1867 VTAIL.n615 VTAIL.n546 185
R1868 VTAIL.n614 VTAIL.n613 185
R1869 VTAIL.n549 VTAIL.n547 185
R1870 VTAIL.n608 VTAIL.n607 185
R1871 VTAIL.n606 VTAIL.n605 185
R1872 VTAIL.n553 VTAIL.n552 185
R1873 VTAIL.n600 VTAIL.n599 185
R1874 VTAIL.n598 VTAIL.n597 185
R1875 VTAIL.n557 VTAIL.n556 185
R1876 VTAIL.n592 VTAIL.n591 185
R1877 VTAIL.n590 VTAIL.n589 185
R1878 VTAIL.n561 VTAIL.n560 185
R1879 VTAIL.n584 VTAIL.n583 185
R1880 VTAIL.n582 VTAIL.n581 185
R1881 VTAIL.n565 VTAIL.n564 185
R1882 VTAIL.n576 VTAIL.n575 185
R1883 VTAIL.n574 VTAIL.n573 185
R1884 VTAIL.n569 VTAIL.n568 185
R1885 VTAIL.n535 VTAIL.n534 185
R1886 VTAIL.n533 VTAIL.n532 185
R1887 VTAIL.n454 VTAIL.n453 185
R1888 VTAIL.n527 VTAIL.n526 185
R1889 VTAIL.n525 VTAIL.n456 185
R1890 VTAIL.n524 VTAIL.n523 185
R1891 VTAIL.n459 VTAIL.n457 185
R1892 VTAIL.n518 VTAIL.n517 185
R1893 VTAIL.n516 VTAIL.n515 185
R1894 VTAIL.n463 VTAIL.n462 185
R1895 VTAIL.n510 VTAIL.n509 185
R1896 VTAIL.n508 VTAIL.n507 185
R1897 VTAIL.n467 VTAIL.n466 185
R1898 VTAIL.n502 VTAIL.n501 185
R1899 VTAIL.n500 VTAIL.n499 185
R1900 VTAIL.n471 VTAIL.n470 185
R1901 VTAIL.n494 VTAIL.n493 185
R1902 VTAIL.n492 VTAIL.n491 185
R1903 VTAIL.n475 VTAIL.n474 185
R1904 VTAIL.n486 VTAIL.n485 185
R1905 VTAIL.n484 VTAIL.n483 185
R1906 VTAIL.n479 VTAIL.n478 185
R1907 VTAIL.n445 VTAIL.n444 185
R1908 VTAIL.n443 VTAIL.n442 185
R1909 VTAIL.n364 VTAIL.n363 185
R1910 VTAIL.n437 VTAIL.n436 185
R1911 VTAIL.n435 VTAIL.n366 185
R1912 VTAIL.n434 VTAIL.n433 185
R1913 VTAIL.n369 VTAIL.n367 185
R1914 VTAIL.n428 VTAIL.n427 185
R1915 VTAIL.n426 VTAIL.n425 185
R1916 VTAIL.n373 VTAIL.n372 185
R1917 VTAIL.n420 VTAIL.n419 185
R1918 VTAIL.n418 VTAIL.n417 185
R1919 VTAIL.n377 VTAIL.n376 185
R1920 VTAIL.n412 VTAIL.n411 185
R1921 VTAIL.n410 VTAIL.n409 185
R1922 VTAIL.n381 VTAIL.n380 185
R1923 VTAIL.n404 VTAIL.n403 185
R1924 VTAIL.n402 VTAIL.n401 185
R1925 VTAIL.n385 VTAIL.n384 185
R1926 VTAIL.n396 VTAIL.n395 185
R1927 VTAIL.n394 VTAIL.n393 185
R1928 VTAIL.n389 VTAIL.n388 185
R1929 VTAIL.n355 VTAIL.n354 185
R1930 VTAIL.n353 VTAIL.n352 185
R1931 VTAIL.n274 VTAIL.n273 185
R1932 VTAIL.n347 VTAIL.n346 185
R1933 VTAIL.n345 VTAIL.n276 185
R1934 VTAIL.n344 VTAIL.n343 185
R1935 VTAIL.n279 VTAIL.n277 185
R1936 VTAIL.n338 VTAIL.n337 185
R1937 VTAIL.n336 VTAIL.n335 185
R1938 VTAIL.n283 VTAIL.n282 185
R1939 VTAIL.n330 VTAIL.n329 185
R1940 VTAIL.n328 VTAIL.n327 185
R1941 VTAIL.n287 VTAIL.n286 185
R1942 VTAIL.n322 VTAIL.n321 185
R1943 VTAIL.n320 VTAIL.n319 185
R1944 VTAIL.n291 VTAIL.n290 185
R1945 VTAIL.n314 VTAIL.n313 185
R1946 VTAIL.n312 VTAIL.n311 185
R1947 VTAIL.n295 VTAIL.n294 185
R1948 VTAIL.n306 VTAIL.n305 185
R1949 VTAIL.n304 VTAIL.n303 185
R1950 VTAIL.n299 VTAIL.n298 185
R1951 VTAIL.n659 VTAIL.t2 147.659
R1952 VTAIL.n29 VTAIL.t0 147.659
R1953 VTAIL.n119 VTAIL.t4 147.659
R1954 VTAIL.n209 VTAIL.t6 147.659
R1955 VTAIL.n570 VTAIL.t5 147.659
R1956 VTAIL.n480 VTAIL.t7 147.659
R1957 VTAIL.n390 VTAIL.t3 147.659
R1958 VTAIL.n300 VTAIL.t1 147.659
R1959 VTAIL.n663 VTAIL.n657 104.615
R1960 VTAIL.n664 VTAIL.n663 104.615
R1961 VTAIL.n664 VTAIL.n653 104.615
R1962 VTAIL.n671 VTAIL.n653 104.615
R1963 VTAIL.n672 VTAIL.n671 104.615
R1964 VTAIL.n672 VTAIL.n649 104.615
R1965 VTAIL.n679 VTAIL.n649 104.615
R1966 VTAIL.n680 VTAIL.n679 104.615
R1967 VTAIL.n680 VTAIL.n645 104.615
R1968 VTAIL.n687 VTAIL.n645 104.615
R1969 VTAIL.n688 VTAIL.n687 104.615
R1970 VTAIL.n688 VTAIL.n641 104.615
R1971 VTAIL.n695 VTAIL.n641 104.615
R1972 VTAIL.n696 VTAIL.n695 104.615
R1973 VTAIL.n696 VTAIL.n637 104.615
R1974 VTAIL.n704 VTAIL.n637 104.615
R1975 VTAIL.n705 VTAIL.n704 104.615
R1976 VTAIL.n706 VTAIL.n705 104.615
R1977 VTAIL.n706 VTAIL.n633 104.615
R1978 VTAIL.n713 VTAIL.n633 104.615
R1979 VTAIL.n714 VTAIL.n713 104.615
R1980 VTAIL.n33 VTAIL.n27 104.615
R1981 VTAIL.n34 VTAIL.n33 104.615
R1982 VTAIL.n34 VTAIL.n23 104.615
R1983 VTAIL.n41 VTAIL.n23 104.615
R1984 VTAIL.n42 VTAIL.n41 104.615
R1985 VTAIL.n42 VTAIL.n19 104.615
R1986 VTAIL.n49 VTAIL.n19 104.615
R1987 VTAIL.n50 VTAIL.n49 104.615
R1988 VTAIL.n50 VTAIL.n15 104.615
R1989 VTAIL.n57 VTAIL.n15 104.615
R1990 VTAIL.n58 VTAIL.n57 104.615
R1991 VTAIL.n58 VTAIL.n11 104.615
R1992 VTAIL.n65 VTAIL.n11 104.615
R1993 VTAIL.n66 VTAIL.n65 104.615
R1994 VTAIL.n66 VTAIL.n7 104.615
R1995 VTAIL.n74 VTAIL.n7 104.615
R1996 VTAIL.n75 VTAIL.n74 104.615
R1997 VTAIL.n76 VTAIL.n75 104.615
R1998 VTAIL.n76 VTAIL.n3 104.615
R1999 VTAIL.n83 VTAIL.n3 104.615
R2000 VTAIL.n84 VTAIL.n83 104.615
R2001 VTAIL.n123 VTAIL.n117 104.615
R2002 VTAIL.n124 VTAIL.n123 104.615
R2003 VTAIL.n124 VTAIL.n113 104.615
R2004 VTAIL.n131 VTAIL.n113 104.615
R2005 VTAIL.n132 VTAIL.n131 104.615
R2006 VTAIL.n132 VTAIL.n109 104.615
R2007 VTAIL.n139 VTAIL.n109 104.615
R2008 VTAIL.n140 VTAIL.n139 104.615
R2009 VTAIL.n140 VTAIL.n105 104.615
R2010 VTAIL.n147 VTAIL.n105 104.615
R2011 VTAIL.n148 VTAIL.n147 104.615
R2012 VTAIL.n148 VTAIL.n101 104.615
R2013 VTAIL.n155 VTAIL.n101 104.615
R2014 VTAIL.n156 VTAIL.n155 104.615
R2015 VTAIL.n156 VTAIL.n97 104.615
R2016 VTAIL.n164 VTAIL.n97 104.615
R2017 VTAIL.n165 VTAIL.n164 104.615
R2018 VTAIL.n166 VTAIL.n165 104.615
R2019 VTAIL.n166 VTAIL.n93 104.615
R2020 VTAIL.n173 VTAIL.n93 104.615
R2021 VTAIL.n174 VTAIL.n173 104.615
R2022 VTAIL.n213 VTAIL.n207 104.615
R2023 VTAIL.n214 VTAIL.n213 104.615
R2024 VTAIL.n214 VTAIL.n203 104.615
R2025 VTAIL.n221 VTAIL.n203 104.615
R2026 VTAIL.n222 VTAIL.n221 104.615
R2027 VTAIL.n222 VTAIL.n199 104.615
R2028 VTAIL.n229 VTAIL.n199 104.615
R2029 VTAIL.n230 VTAIL.n229 104.615
R2030 VTAIL.n230 VTAIL.n195 104.615
R2031 VTAIL.n237 VTAIL.n195 104.615
R2032 VTAIL.n238 VTAIL.n237 104.615
R2033 VTAIL.n238 VTAIL.n191 104.615
R2034 VTAIL.n245 VTAIL.n191 104.615
R2035 VTAIL.n246 VTAIL.n245 104.615
R2036 VTAIL.n246 VTAIL.n187 104.615
R2037 VTAIL.n254 VTAIL.n187 104.615
R2038 VTAIL.n255 VTAIL.n254 104.615
R2039 VTAIL.n256 VTAIL.n255 104.615
R2040 VTAIL.n256 VTAIL.n183 104.615
R2041 VTAIL.n263 VTAIL.n183 104.615
R2042 VTAIL.n264 VTAIL.n263 104.615
R2043 VTAIL.n624 VTAIL.n623 104.615
R2044 VTAIL.n623 VTAIL.n543 104.615
R2045 VTAIL.n616 VTAIL.n543 104.615
R2046 VTAIL.n616 VTAIL.n615 104.615
R2047 VTAIL.n615 VTAIL.n614 104.615
R2048 VTAIL.n614 VTAIL.n547 104.615
R2049 VTAIL.n607 VTAIL.n547 104.615
R2050 VTAIL.n607 VTAIL.n606 104.615
R2051 VTAIL.n606 VTAIL.n552 104.615
R2052 VTAIL.n599 VTAIL.n552 104.615
R2053 VTAIL.n599 VTAIL.n598 104.615
R2054 VTAIL.n598 VTAIL.n556 104.615
R2055 VTAIL.n591 VTAIL.n556 104.615
R2056 VTAIL.n591 VTAIL.n590 104.615
R2057 VTAIL.n590 VTAIL.n560 104.615
R2058 VTAIL.n583 VTAIL.n560 104.615
R2059 VTAIL.n583 VTAIL.n582 104.615
R2060 VTAIL.n582 VTAIL.n564 104.615
R2061 VTAIL.n575 VTAIL.n564 104.615
R2062 VTAIL.n575 VTAIL.n574 104.615
R2063 VTAIL.n574 VTAIL.n568 104.615
R2064 VTAIL.n534 VTAIL.n533 104.615
R2065 VTAIL.n533 VTAIL.n453 104.615
R2066 VTAIL.n526 VTAIL.n453 104.615
R2067 VTAIL.n526 VTAIL.n525 104.615
R2068 VTAIL.n525 VTAIL.n524 104.615
R2069 VTAIL.n524 VTAIL.n457 104.615
R2070 VTAIL.n517 VTAIL.n457 104.615
R2071 VTAIL.n517 VTAIL.n516 104.615
R2072 VTAIL.n516 VTAIL.n462 104.615
R2073 VTAIL.n509 VTAIL.n462 104.615
R2074 VTAIL.n509 VTAIL.n508 104.615
R2075 VTAIL.n508 VTAIL.n466 104.615
R2076 VTAIL.n501 VTAIL.n466 104.615
R2077 VTAIL.n501 VTAIL.n500 104.615
R2078 VTAIL.n500 VTAIL.n470 104.615
R2079 VTAIL.n493 VTAIL.n470 104.615
R2080 VTAIL.n493 VTAIL.n492 104.615
R2081 VTAIL.n492 VTAIL.n474 104.615
R2082 VTAIL.n485 VTAIL.n474 104.615
R2083 VTAIL.n485 VTAIL.n484 104.615
R2084 VTAIL.n484 VTAIL.n478 104.615
R2085 VTAIL.n444 VTAIL.n443 104.615
R2086 VTAIL.n443 VTAIL.n363 104.615
R2087 VTAIL.n436 VTAIL.n363 104.615
R2088 VTAIL.n436 VTAIL.n435 104.615
R2089 VTAIL.n435 VTAIL.n434 104.615
R2090 VTAIL.n434 VTAIL.n367 104.615
R2091 VTAIL.n427 VTAIL.n367 104.615
R2092 VTAIL.n427 VTAIL.n426 104.615
R2093 VTAIL.n426 VTAIL.n372 104.615
R2094 VTAIL.n419 VTAIL.n372 104.615
R2095 VTAIL.n419 VTAIL.n418 104.615
R2096 VTAIL.n418 VTAIL.n376 104.615
R2097 VTAIL.n411 VTAIL.n376 104.615
R2098 VTAIL.n411 VTAIL.n410 104.615
R2099 VTAIL.n410 VTAIL.n380 104.615
R2100 VTAIL.n403 VTAIL.n380 104.615
R2101 VTAIL.n403 VTAIL.n402 104.615
R2102 VTAIL.n402 VTAIL.n384 104.615
R2103 VTAIL.n395 VTAIL.n384 104.615
R2104 VTAIL.n395 VTAIL.n394 104.615
R2105 VTAIL.n394 VTAIL.n388 104.615
R2106 VTAIL.n354 VTAIL.n353 104.615
R2107 VTAIL.n353 VTAIL.n273 104.615
R2108 VTAIL.n346 VTAIL.n273 104.615
R2109 VTAIL.n346 VTAIL.n345 104.615
R2110 VTAIL.n345 VTAIL.n344 104.615
R2111 VTAIL.n344 VTAIL.n277 104.615
R2112 VTAIL.n337 VTAIL.n277 104.615
R2113 VTAIL.n337 VTAIL.n336 104.615
R2114 VTAIL.n336 VTAIL.n282 104.615
R2115 VTAIL.n329 VTAIL.n282 104.615
R2116 VTAIL.n329 VTAIL.n328 104.615
R2117 VTAIL.n328 VTAIL.n286 104.615
R2118 VTAIL.n321 VTAIL.n286 104.615
R2119 VTAIL.n321 VTAIL.n320 104.615
R2120 VTAIL.n320 VTAIL.n290 104.615
R2121 VTAIL.n313 VTAIL.n290 104.615
R2122 VTAIL.n313 VTAIL.n312 104.615
R2123 VTAIL.n312 VTAIL.n294 104.615
R2124 VTAIL.n305 VTAIL.n294 104.615
R2125 VTAIL.n305 VTAIL.n304 104.615
R2126 VTAIL.n304 VTAIL.n298 104.615
R2127 VTAIL.t2 VTAIL.n657 52.3082
R2128 VTAIL.t0 VTAIL.n27 52.3082
R2129 VTAIL.t4 VTAIL.n117 52.3082
R2130 VTAIL.t6 VTAIL.n207 52.3082
R2131 VTAIL.t5 VTAIL.n568 52.3082
R2132 VTAIL.t7 VTAIL.n478 52.3082
R2133 VTAIL.t3 VTAIL.n388 52.3082
R2134 VTAIL.t1 VTAIL.n298 52.3082
R2135 VTAIL.n719 VTAIL.n718 30.6338
R2136 VTAIL.n89 VTAIL.n88 30.6338
R2137 VTAIL.n179 VTAIL.n178 30.6338
R2138 VTAIL.n269 VTAIL.n268 30.6338
R2139 VTAIL.n629 VTAIL.n628 30.6338
R2140 VTAIL.n539 VTAIL.n538 30.6338
R2141 VTAIL.n449 VTAIL.n448 30.6338
R2142 VTAIL.n359 VTAIL.n358 30.6338
R2143 VTAIL.n719 VTAIL.n629 29.5134
R2144 VTAIL.n359 VTAIL.n269 29.5134
R2145 VTAIL.n659 VTAIL.n658 15.6677
R2146 VTAIL.n29 VTAIL.n28 15.6677
R2147 VTAIL.n119 VTAIL.n118 15.6677
R2148 VTAIL.n209 VTAIL.n208 15.6677
R2149 VTAIL.n570 VTAIL.n569 15.6677
R2150 VTAIL.n480 VTAIL.n479 15.6677
R2151 VTAIL.n390 VTAIL.n389 15.6677
R2152 VTAIL.n300 VTAIL.n299 15.6677
R2153 VTAIL.n707 VTAIL.n636 13.1884
R2154 VTAIL.n77 VTAIL.n6 13.1884
R2155 VTAIL.n167 VTAIL.n96 13.1884
R2156 VTAIL.n257 VTAIL.n186 13.1884
R2157 VTAIL.n617 VTAIL.n546 13.1884
R2158 VTAIL.n527 VTAIL.n456 13.1884
R2159 VTAIL.n437 VTAIL.n366 13.1884
R2160 VTAIL.n347 VTAIL.n276 13.1884
R2161 VTAIL.n662 VTAIL.n661 12.8005
R2162 VTAIL.n703 VTAIL.n702 12.8005
R2163 VTAIL.n708 VTAIL.n634 12.8005
R2164 VTAIL.n32 VTAIL.n31 12.8005
R2165 VTAIL.n73 VTAIL.n72 12.8005
R2166 VTAIL.n78 VTAIL.n4 12.8005
R2167 VTAIL.n122 VTAIL.n121 12.8005
R2168 VTAIL.n163 VTAIL.n162 12.8005
R2169 VTAIL.n168 VTAIL.n94 12.8005
R2170 VTAIL.n212 VTAIL.n211 12.8005
R2171 VTAIL.n253 VTAIL.n252 12.8005
R2172 VTAIL.n258 VTAIL.n184 12.8005
R2173 VTAIL.n618 VTAIL.n544 12.8005
R2174 VTAIL.n613 VTAIL.n548 12.8005
R2175 VTAIL.n573 VTAIL.n572 12.8005
R2176 VTAIL.n528 VTAIL.n454 12.8005
R2177 VTAIL.n523 VTAIL.n458 12.8005
R2178 VTAIL.n483 VTAIL.n482 12.8005
R2179 VTAIL.n438 VTAIL.n364 12.8005
R2180 VTAIL.n433 VTAIL.n368 12.8005
R2181 VTAIL.n393 VTAIL.n392 12.8005
R2182 VTAIL.n348 VTAIL.n274 12.8005
R2183 VTAIL.n343 VTAIL.n278 12.8005
R2184 VTAIL.n303 VTAIL.n302 12.8005
R2185 VTAIL.n665 VTAIL.n656 12.0247
R2186 VTAIL.n701 VTAIL.n638 12.0247
R2187 VTAIL.n712 VTAIL.n711 12.0247
R2188 VTAIL.n35 VTAIL.n26 12.0247
R2189 VTAIL.n71 VTAIL.n8 12.0247
R2190 VTAIL.n82 VTAIL.n81 12.0247
R2191 VTAIL.n125 VTAIL.n116 12.0247
R2192 VTAIL.n161 VTAIL.n98 12.0247
R2193 VTAIL.n172 VTAIL.n171 12.0247
R2194 VTAIL.n215 VTAIL.n206 12.0247
R2195 VTAIL.n251 VTAIL.n188 12.0247
R2196 VTAIL.n262 VTAIL.n261 12.0247
R2197 VTAIL.n622 VTAIL.n621 12.0247
R2198 VTAIL.n612 VTAIL.n549 12.0247
R2199 VTAIL.n576 VTAIL.n567 12.0247
R2200 VTAIL.n532 VTAIL.n531 12.0247
R2201 VTAIL.n522 VTAIL.n459 12.0247
R2202 VTAIL.n486 VTAIL.n477 12.0247
R2203 VTAIL.n442 VTAIL.n441 12.0247
R2204 VTAIL.n432 VTAIL.n369 12.0247
R2205 VTAIL.n396 VTAIL.n387 12.0247
R2206 VTAIL.n352 VTAIL.n351 12.0247
R2207 VTAIL.n342 VTAIL.n279 12.0247
R2208 VTAIL.n306 VTAIL.n297 12.0247
R2209 VTAIL.n666 VTAIL.n654 11.249
R2210 VTAIL.n698 VTAIL.n697 11.249
R2211 VTAIL.n715 VTAIL.n632 11.249
R2212 VTAIL.n36 VTAIL.n24 11.249
R2213 VTAIL.n68 VTAIL.n67 11.249
R2214 VTAIL.n85 VTAIL.n2 11.249
R2215 VTAIL.n126 VTAIL.n114 11.249
R2216 VTAIL.n158 VTAIL.n157 11.249
R2217 VTAIL.n175 VTAIL.n92 11.249
R2218 VTAIL.n216 VTAIL.n204 11.249
R2219 VTAIL.n248 VTAIL.n247 11.249
R2220 VTAIL.n265 VTAIL.n182 11.249
R2221 VTAIL.n625 VTAIL.n542 11.249
R2222 VTAIL.n609 VTAIL.n608 11.249
R2223 VTAIL.n577 VTAIL.n565 11.249
R2224 VTAIL.n535 VTAIL.n452 11.249
R2225 VTAIL.n519 VTAIL.n518 11.249
R2226 VTAIL.n487 VTAIL.n475 11.249
R2227 VTAIL.n445 VTAIL.n362 11.249
R2228 VTAIL.n429 VTAIL.n428 11.249
R2229 VTAIL.n397 VTAIL.n385 11.249
R2230 VTAIL.n355 VTAIL.n272 11.249
R2231 VTAIL.n339 VTAIL.n338 11.249
R2232 VTAIL.n307 VTAIL.n295 11.249
R2233 VTAIL.n670 VTAIL.n669 10.4732
R2234 VTAIL.n694 VTAIL.n640 10.4732
R2235 VTAIL.n716 VTAIL.n630 10.4732
R2236 VTAIL.n40 VTAIL.n39 10.4732
R2237 VTAIL.n64 VTAIL.n10 10.4732
R2238 VTAIL.n86 VTAIL.n0 10.4732
R2239 VTAIL.n130 VTAIL.n129 10.4732
R2240 VTAIL.n154 VTAIL.n100 10.4732
R2241 VTAIL.n176 VTAIL.n90 10.4732
R2242 VTAIL.n220 VTAIL.n219 10.4732
R2243 VTAIL.n244 VTAIL.n190 10.4732
R2244 VTAIL.n266 VTAIL.n180 10.4732
R2245 VTAIL.n626 VTAIL.n540 10.4732
R2246 VTAIL.n605 VTAIL.n551 10.4732
R2247 VTAIL.n581 VTAIL.n580 10.4732
R2248 VTAIL.n536 VTAIL.n450 10.4732
R2249 VTAIL.n515 VTAIL.n461 10.4732
R2250 VTAIL.n491 VTAIL.n490 10.4732
R2251 VTAIL.n446 VTAIL.n360 10.4732
R2252 VTAIL.n425 VTAIL.n371 10.4732
R2253 VTAIL.n401 VTAIL.n400 10.4732
R2254 VTAIL.n356 VTAIL.n270 10.4732
R2255 VTAIL.n335 VTAIL.n281 10.4732
R2256 VTAIL.n311 VTAIL.n310 10.4732
R2257 VTAIL.n673 VTAIL.n652 9.69747
R2258 VTAIL.n693 VTAIL.n642 9.69747
R2259 VTAIL.n43 VTAIL.n22 9.69747
R2260 VTAIL.n63 VTAIL.n12 9.69747
R2261 VTAIL.n133 VTAIL.n112 9.69747
R2262 VTAIL.n153 VTAIL.n102 9.69747
R2263 VTAIL.n223 VTAIL.n202 9.69747
R2264 VTAIL.n243 VTAIL.n192 9.69747
R2265 VTAIL.n604 VTAIL.n553 9.69747
R2266 VTAIL.n584 VTAIL.n563 9.69747
R2267 VTAIL.n514 VTAIL.n463 9.69747
R2268 VTAIL.n494 VTAIL.n473 9.69747
R2269 VTAIL.n424 VTAIL.n373 9.69747
R2270 VTAIL.n404 VTAIL.n383 9.69747
R2271 VTAIL.n334 VTAIL.n283 9.69747
R2272 VTAIL.n314 VTAIL.n293 9.69747
R2273 VTAIL.n718 VTAIL.n717 9.45567
R2274 VTAIL.n88 VTAIL.n87 9.45567
R2275 VTAIL.n178 VTAIL.n177 9.45567
R2276 VTAIL.n268 VTAIL.n267 9.45567
R2277 VTAIL.n628 VTAIL.n627 9.45567
R2278 VTAIL.n538 VTAIL.n537 9.45567
R2279 VTAIL.n448 VTAIL.n447 9.45567
R2280 VTAIL.n358 VTAIL.n357 9.45567
R2281 VTAIL.n717 VTAIL.n716 9.3005
R2282 VTAIL.n632 VTAIL.n631 9.3005
R2283 VTAIL.n711 VTAIL.n710 9.3005
R2284 VTAIL.n709 VTAIL.n708 9.3005
R2285 VTAIL.n648 VTAIL.n647 9.3005
R2286 VTAIL.n677 VTAIL.n676 9.3005
R2287 VTAIL.n675 VTAIL.n674 9.3005
R2288 VTAIL.n652 VTAIL.n651 9.3005
R2289 VTAIL.n669 VTAIL.n668 9.3005
R2290 VTAIL.n667 VTAIL.n666 9.3005
R2291 VTAIL.n656 VTAIL.n655 9.3005
R2292 VTAIL.n661 VTAIL.n660 9.3005
R2293 VTAIL.n683 VTAIL.n682 9.3005
R2294 VTAIL.n685 VTAIL.n684 9.3005
R2295 VTAIL.n644 VTAIL.n643 9.3005
R2296 VTAIL.n691 VTAIL.n690 9.3005
R2297 VTAIL.n693 VTAIL.n692 9.3005
R2298 VTAIL.n640 VTAIL.n639 9.3005
R2299 VTAIL.n699 VTAIL.n698 9.3005
R2300 VTAIL.n701 VTAIL.n700 9.3005
R2301 VTAIL.n702 VTAIL.n635 9.3005
R2302 VTAIL.n87 VTAIL.n86 9.3005
R2303 VTAIL.n2 VTAIL.n1 9.3005
R2304 VTAIL.n81 VTAIL.n80 9.3005
R2305 VTAIL.n79 VTAIL.n78 9.3005
R2306 VTAIL.n18 VTAIL.n17 9.3005
R2307 VTAIL.n47 VTAIL.n46 9.3005
R2308 VTAIL.n45 VTAIL.n44 9.3005
R2309 VTAIL.n22 VTAIL.n21 9.3005
R2310 VTAIL.n39 VTAIL.n38 9.3005
R2311 VTAIL.n37 VTAIL.n36 9.3005
R2312 VTAIL.n26 VTAIL.n25 9.3005
R2313 VTAIL.n31 VTAIL.n30 9.3005
R2314 VTAIL.n53 VTAIL.n52 9.3005
R2315 VTAIL.n55 VTAIL.n54 9.3005
R2316 VTAIL.n14 VTAIL.n13 9.3005
R2317 VTAIL.n61 VTAIL.n60 9.3005
R2318 VTAIL.n63 VTAIL.n62 9.3005
R2319 VTAIL.n10 VTAIL.n9 9.3005
R2320 VTAIL.n69 VTAIL.n68 9.3005
R2321 VTAIL.n71 VTAIL.n70 9.3005
R2322 VTAIL.n72 VTAIL.n5 9.3005
R2323 VTAIL.n177 VTAIL.n176 9.3005
R2324 VTAIL.n92 VTAIL.n91 9.3005
R2325 VTAIL.n171 VTAIL.n170 9.3005
R2326 VTAIL.n169 VTAIL.n168 9.3005
R2327 VTAIL.n108 VTAIL.n107 9.3005
R2328 VTAIL.n137 VTAIL.n136 9.3005
R2329 VTAIL.n135 VTAIL.n134 9.3005
R2330 VTAIL.n112 VTAIL.n111 9.3005
R2331 VTAIL.n129 VTAIL.n128 9.3005
R2332 VTAIL.n127 VTAIL.n126 9.3005
R2333 VTAIL.n116 VTAIL.n115 9.3005
R2334 VTAIL.n121 VTAIL.n120 9.3005
R2335 VTAIL.n143 VTAIL.n142 9.3005
R2336 VTAIL.n145 VTAIL.n144 9.3005
R2337 VTAIL.n104 VTAIL.n103 9.3005
R2338 VTAIL.n151 VTAIL.n150 9.3005
R2339 VTAIL.n153 VTAIL.n152 9.3005
R2340 VTAIL.n100 VTAIL.n99 9.3005
R2341 VTAIL.n159 VTAIL.n158 9.3005
R2342 VTAIL.n161 VTAIL.n160 9.3005
R2343 VTAIL.n162 VTAIL.n95 9.3005
R2344 VTAIL.n267 VTAIL.n266 9.3005
R2345 VTAIL.n182 VTAIL.n181 9.3005
R2346 VTAIL.n261 VTAIL.n260 9.3005
R2347 VTAIL.n259 VTAIL.n258 9.3005
R2348 VTAIL.n198 VTAIL.n197 9.3005
R2349 VTAIL.n227 VTAIL.n226 9.3005
R2350 VTAIL.n225 VTAIL.n224 9.3005
R2351 VTAIL.n202 VTAIL.n201 9.3005
R2352 VTAIL.n219 VTAIL.n218 9.3005
R2353 VTAIL.n217 VTAIL.n216 9.3005
R2354 VTAIL.n206 VTAIL.n205 9.3005
R2355 VTAIL.n211 VTAIL.n210 9.3005
R2356 VTAIL.n233 VTAIL.n232 9.3005
R2357 VTAIL.n235 VTAIL.n234 9.3005
R2358 VTAIL.n194 VTAIL.n193 9.3005
R2359 VTAIL.n241 VTAIL.n240 9.3005
R2360 VTAIL.n243 VTAIL.n242 9.3005
R2361 VTAIL.n190 VTAIL.n189 9.3005
R2362 VTAIL.n249 VTAIL.n248 9.3005
R2363 VTAIL.n251 VTAIL.n250 9.3005
R2364 VTAIL.n252 VTAIL.n185 9.3005
R2365 VTAIL.n596 VTAIL.n595 9.3005
R2366 VTAIL.n555 VTAIL.n554 9.3005
R2367 VTAIL.n602 VTAIL.n601 9.3005
R2368 VTAIL.n604 VTAIL.n603 9.3005
R2369 VTAIL.n551 VTAIL.n550 9.3005
R2370 VTAIL.n610 VTAIL.n609 9.3005
R2371 VTAIL.n612 VTAIL.n611 9.3005
R2372 VTAIL.n548 VTAIL.n545 9.3005
R2373 VTAIL.n627 VTAIL.n626 9.3005
R2374 VTAIL.n542 VTAIL.n541 9.3005
R2375 VTAIL.n621 VTAIL.n620 9.3005
R2376 VTAIL.n619 VTAIL.n618 9.3005
R2377 VTAIL.n594 VTAIL.n593 9.3005
R2378 VTAIL.n559 VTAIL.n558 9.3005
R2379 VTAIL.n588 VTAIL.n587 9.3005
R2380 VTAIL.n586 VTAIL.n585 9.3005
R2381 VTAIL.n563 VTAIL.n562 9.3005
R2382 VTAIL.n580 VTAIL.n579 9.3005
R2383 VTAIL.n578 VTAIL.n577 9.3005
R2384 VTAIL.n567 VTAIL.n566 9.3005
R2385 VTAIL.n572 VTAIL.n571 9.3005
R2386 VTAIL.n506 VTAIL.n505 9.3005
R2387 VTAIL.n465 VTAIL.n464 9.3005
R2388 VTAIL.n512 VTAIL.n511 9.3005
R2389 VTAIL.n514 VTAIL.n513 9.3005
R2390 VTAIL.n461 VTAIL.n460 9.3005
R2391 VTAIL.n520 VTAIL.n519 9.3005
R2392 VTAIL.n522 VTAIL.n521 9.3005
R2393 VTAIL.n458 VTAIL.n455 9.3005
R2394 VTAIL.n537 VTAIL.n536 9.3005
R2395 VTAIL.n452 VTAIL.n451 9.3005
R2396 VTAIL.n531 VTAIL.n530 9.3005
R2397 VTAIL.n529 VTAIL.n528 9.3005
R2398 VTAIL.n504 VTAIL.n503 9.3005
R2399 VTAIL.n469 VTAIL.n468 9.3005
R2400 VTAIL.n498 VTAIL.n497 9.3005
R2401 VTAIL.n496 VTAIL.n495 9.3005
R2402 VTAIL.n473 VTAIL.n472 9.3005
R2403 VTAIL.n490 VTAIL.n489 9.3005
R2404 VTAIL.n488 VTAIL.n487 9.3005
R2405 VTAIL.n477 VTAIL.n476 9.3005
R2406 VTAIL.n482 VTAIL.n481 9.3005
R2407 VTAIL.n416 VTAIL.n415 9.3005
R2408 VTAIL.n375 VTAIL.n374 9.3005
R2409 VTAIL.n422 VTAIL.n421 9.3005
R2410 VTAIL.n424 VTAIL.n423 9.3005
R2411 VTAIL.n371 VTAIL.n370 9.3005
R2412 VTAIL.n430 VTAIL.n429 9.3005
R2413 VTAIL.n432 VTAIL.n431 9.3005
R2414 VTAIL.n368 VTAIL.n365 9.3005
R2415 VTAIL.n447 VTAIL.n446 9.3005
R2416 VTAIL.n362 VTAIL.n361 9.3005
R2417 VTAIL.n441 VTAIL.n440 9.3005
R2418 VTAIL.n439 VTAIL.n438 9.3005
R2419 VTAIL.n414 VTAIL.n413 9.3005
R2420 VTAIL.n379 VTAIL.n378 9.3005
R2421 VTAIL.n408 VTAIL.n407 9.3005
R2422 VTAIL.n406 VTAIL.n405 9.3005
R2423 VTAIL.n383 VTAIL.n382 9.3005
R2424 VTAIL.n400 VTAIL.n399 9.3005
R2425 VTAIL.n398 VTAIL.n397 9.3005
R2426 VTAIL.n387 VTAIL.n386 9.3005
R2427 VTAIL.n392 VTAIL.n391 9.3005
R2428 VTAIL.n326 VTAIL.n325 9.3005
R2429 VTAIL.n285 VTAIL.n284 9.3005
R2430 VTAIL.n332 VTAIL.n331 9.3005
R2431 VTAIL.n334 VTAIL.n333 9.3005
R2432 VTAIL.n281 VTAIL.n280 9.3005
R2433 VTAIL.n340 VTAIL.n339 9.3005
R2434 VTAIL.n342 VTAIL.n341 9.3005
R2435 VTAIL.n278 VTAIL.n275 9.3005
R2436 VTAIL.n357 VTAIL.n356 9.3005
R2437 VTAIL.n272 VTAIL.n271 9.3005
R2438 VTAIL.n351 VTAIL.n350 9.3005
R2439 VTAIL.n349 VTAIL.n348 9.3005
R2440 VTAIL.n324 VTAIL.n323 9.3005
R2441 VTAIL.n289 VTAIL.n288 9.3005
R2442 VTAIL.n318 VTAIL.n317 9.3005
R2443 VTAIL.n316 VTAIL.n315 9.3005
R2444 VTAIL.n293 VTAIL.n292 9.3005
R2445 VTAIL.n310 VTAIL.n309 9.3005
R2446 VTAIL.n308 VTAIL.n307 9.3005
R2447 VTAIL.n297 VTAIL.n296 9.3005
R2448 VTAIL.n302 VTAIL.n301 9.3005
R2449 VTAIL.n674 VTAIL.n650 8.92171
R2450 VTAIL.n690 VTAIL.n689 8.92171
R2451 VTAIL.n44 VTAIL.n20 8.92171
R2452 VTAIL.n60 VTAIL.n59 8.92171
R2453 VTAIL.n134 VTAIL.n110 8.92171
R2454 VTAIL.n150 VTAIL.n149 8.92171
R2455 VTAIL.n224 VTAIL.n200 8.92171
R2456 VTAIL.n240 VTAIL.n239 8.92171
R2457 VTAIL.n601 VTAIL.n600 8.92171
R2458 VTAIL.n585 VTAIL.n561 8.92171
R2459 VTAIL.n511 VTAIL.n510 8.92171
R2460 VTAIL.n495 VTAIL.n471 8.92171
R2461 VTAIL.n421 VTAIL.n420 8.92171
R2462 VTAIL.n405 VTAIL.n381 8.92171
R2463 VTAIL.n331 VTAIL.n330 8.92171
R2464 VTAIL.n315 VTAIL.n291 8.92171
R2465 VTAIL.n678 VTAIL.n677 8.14595
R2466 VTAIL.n686 VTAIL.n644 8.14595
R2467 VTAIL.n48 VTAIL.n47 8.14595
R2468 VTAIL.n56 VTAIL.n14 8.14595
R2469 VTAIL.n138 VTAIL.n137 8.14595
R2470 VTAIL.n146 VTAIL.n104 8.14595
R2471 VTAIL.n228 VTAIL.n227 8.14595
R2472 VTAIL.n236 VTAIL.n194 8.14595
R2473 VTAIL.n597 VTAIL.n555 8.14595
R2474 VTAIL.n589 VTAIL.n588 8.14595
R2475 VTAIL.n507 VTAIL.n465 8.14595
R2476 VTAIL.n499 VTAIL.n498 8.14595
R2477 VTAIL.n417 VTAIL.n375 8.14595
R2478 VTAIL.n409 VTAIL.n408 8.14595
R2479 VTAIL.n327 VTAIL.n285 8.14595
R2480 VTAIL.n319 VTAIL.n318 8.14595
R2481 VTAIL.n681 VTAIL.n648 7.3702
R2482 VTAIL.n685 VTAIL.n646 7.3702
R2483 VTAIL.n51 VTAIL.n18 7.3702
R2484 VTAIL.n55 VTAIL.n16 7.3702
R2485 VTAIL.n141 VTAIL.n108 7.3702
R2486 VTAIL.n145 VTAIL.n106 7.3702
R2487 VTAIL.n231 VTAIL.n198 7.3702
R2488 VTAIL.n235 VTAIL.n196 7.3702
R2489 VTAIL.n596 VTAIL.n557 7.3702
R2490 VTAIL.n592 VTAIL.n559 7.3702
R2491 VTAIL.n506 VTAIL.n467 7.3702
R2492 VTAIL.n502 VTAIL.n469 7.3702
R2493 VTAIL.n416 VTAIL.n377 7.3702
R2494 VTAIL.n412 VTAIL.n379 7.3702
R2495 VTAIL.n326 VTAIL.n287 7.3702
R2496 VTAIL.n322 VTAIL.n289 7.3702
R2497 VTAIL.n682 VTAIL.n681 6.59444
R2498 VTAIL.n682 VTAIL.n646 6.59444
R2499 VTAIL.n52 VTAIL.n51 6.59444
R2500 VTAIL.n52 VTAIL.n16 6.59444
R2501 VTAIL.n142 VTAIL.n141 6.59444
R2502 VTAIL.n142 VTAIL.n106 6.59444
R2503 VTAIL.n232 VTAIL.n231 6.59444
R2504 VTAIL.n232 VTAIL.n196 6.59444
R2505 VTAIL.n593 VTAIL.n557 6.59444
R2506 VTAIL.n593 VTAIL.n592 6.59444
R2507 VTAIL.n503 VTAIL.n467 6.59444
R2508 VTAIL.n503 VTAIL.n502 6.59444
R2509 VTAIL.n413 VTAIL.n377 6.59444
R2510 VTAIL.n413 VTAIL.n412 6.59444
R2511 VTAIL.n323 VTAIL.n287 6.59444
R2512 VTAIL.n323 VTAIL.n322 6.59444
R2513 VTAIL.n678 VTAIL.n648 5.81868
R2514 VTAIL.n686 VTAIL.n685 5.81868
R2515 VTAIL.n48 VTAIL.n18 5.81868
R2516 VTAIL.n56 VTAIL.n55 5.81868
R2517 VTAIL.n138 VTAIL.n108 5.81868
R2518 VTAIL.n146 VTAIL.n145 5.81868
R2519 VTAIL.n228 VTAIL.n198 5.81868
R2520 VTAIL.n236 VTAIL.n235 5.81868
R2521 VTAIL.n597 VTAIL.n596 5.81868
R2522 VTAIL.n589 VTAIL.n559 5.81868
R2523 VTAIL.n507 VTAIL.n506 5.81868
R2524 VTAIL.n499 VTAIL.n469 5.81868
R2525 VTAIL.n417 VTAIL.n416 5.81868
R2526 VTAIL.n409 VTAIL.n379 5.81868
R2527 VTAIL.n327 VTAIL.n326 5.81868
R2528 VTAIL.n319 VTAIL.n289 5.81868
R2529 VTAIL.n677 VTAIL.n650 5.04292
R2530 VTAIL.n689 VTAIL.n644 5.04292
R2531 VTAIL.n47 VTAIL.n20 5.04292
R2532 VTAIL.n59 VTAIL.n14 5.04292
R2533 VTAIL.n137 VTAIL.n110 5.04292
R2534 VTAIL.n149 VTAIL.n104 5.04292
R2535 VTAIL.n227 VTAIL.n200 5.04292
R2536 VTAIL.n239 VTAIL.n194 5.04292
R2537 VTAIL.n600 VTAIL.n555 5.04292
R2538 VTAIL.n588 VTAIL.n561 5.04292
R2539 VTAIL.n510 VTAIL.n465 5.04292
R2540 VTAIL.n498 VTAIL.n471 5.04292
R2541 VTAIL.n420 VTAIL.n375 5.04292
R2542 VTAIL.n408 VTAIL.n381 5.04292
R2543 VTAIL.n330 VTAIL.n285 5.04292
R2544 VTAIL.n318 VTAIL.n291 5.04292
R2545 VTAIL.n660 VTAIL.n659 4.38563
R2546 VTAIL.n30 VTAIL.n29 4.38563
R2547 VTAIL.n120 VTAIL.n119 4.38563
R2548 VTAIL.n210 VTAIL.n209 4.38563
R2549 VTAIL.n571 VTAIL.n570 4.38563
R2550 VTAIL.n481 VTAIL.n480 4.38563
R2551 VTAIL.n391 VTAIL.n390 4.38563
R2552 VTAIL.n301 VTAIL.n300 4.38563
R2553 VTAIL.n674 VTAIL.n673 4.26717
R2554 VTAIL.n690 VTAIL.n642 4.26717
R2555 VTAIL.n44 VTAIL.n43 4.26717
R2556 VTAIL.n60 VTAIL.n12 4.26717
R2557 VTAIL.n134 VTAIL.n133 4.26717
R2558 VTAIL.n150 VTAIL.n102 4.26717
R2559 VTAIL.n224 VTAIL.n223 4.26717
R2560 VTAIL.n240 VTAIL.n192 4.26717
R2561 VTAIL.n601 VTAIL.n553 4.26717
R2562 VTAIL.n585 VTAIL.n584 4.26717
R2563 VTAIL.n511 VTAIL.n463 4.26717
R2564 VTAIL.n495 VTAIL.n494 4.26717
R2565 VTAIL.n421 VTAIL.n373 4.26717
R2566 VTAIL.n405 VTAIL.n404 4.26717
R2567 VTAIL.n331 VTAIL.n283 4.26717
R2568 VTAIL.n315 VTAIL.n314 4.26717
R2569 VTAIL.n670 VTAIL.n652 3.49141
R2570 VTAIL.n694 VTAIL.n693 3.49141
R2571 VTAIL.n718 VTAIL.n630 3.49141
R2572 VTAIL.n40 VTAIL.n22 3.49141
R2573 VTAIL.n64 VTAIL.n63 3.49141
R2574 VTAIL.n88 VTAIL.n0 3.49141
R2575 VTAIL.n130 VTAIL.n112 3.49141
R2576 VTAIL.n154 VTAIL.n153 3.49141
R2577 VTAIL.n178 VTAIL.n90 3.49141
R2578 VTAIL.n220 VTAIL.n202 3.49141
R2579 VTAIL.n244 VTAIL.n243 3.49141
R2580 VTAIL.n268 VTAIL.n180 3.49141
R2581 VTAIL.n628 VTAIL.n540 3.49141
R2582 VTAIL.n605 VTAIL.n604 3.49141
R2583 VTAIL.n581 VTAIL.n563 3.49141
R2584 VTAIL.n538 VTAIL.n450 3.49141
R2585 VTAIL.n515 VTAIL.n514 3.49141
R2586 VTAIL.n491 VTAIL.n473 3.49141
R2587 VTAIL.n448 VTAIL.n360 3.49141
R2588 VTAIL.n425 VTAIL.n424 3.49141
R2589 VTAIL.n401 VTAIL.n383 3.49141
R2590 VTAIL.n358 VTAIL.n270 3.49141
R2591 VTAIL.n335 VTAIL.n334 3.49141
R2592 VTAIL.n311 VTAIL.n293 3.49141
R2593 VTAIL.n449 VTAIL.n359 3.35395
R2594 VTAIL.n629 VTAIL.n539 3.35395
R2595 VTAIL.n269 VTAIL.n179 3.35395
R2596 VTAIL.n669 VTAIL.n654 2.71565
R2597 VTAIL.n697 VTAIL.n640 2.71565
R2598 VTAIL.n716 VTAIL.n715 2.71565
R2599 VTAIL.n39 VTAIL.n24 2.71565
R2600 VTAIL.n67 VTAIL.n10 2.71565
R2601 VTAIL.n86 VTAIL.n85 2.71565
R2602 VTAIL.n129 VTAIL.n114 2.71565
R2603 VTAIL.n157 VTAIL.n100 2.71565
R2604 VTAIL.n176 VTAIL.n175 2.71565
R2605 VTAIL.n219 VTAIL.n204 2.71565
R2606 VTAIL.n247 VTAIL.n190 2.71565
R2607 VTAIL.n266 VTAIL.n265 2.71565
R2608 VTAIL.n626 VTAIL.n625 2.71565
R2609 VTAIL.n608 VTAIL.n551 2.71565
R2610 VTAIL.n580 VTAIL.n565 2.71565
R2611 VTAIL.n536 VTAIL.n535 2.71565
R2612 VTAIL.n518 VTAIL.n461 2.71565
R2613 VTAIL.n490 VTAIL.n475 2.71565
R2614 VTAIL.n446 VTAIL.n445 2.71565
R2615 VTAIL.n428 VTAIL.n371 2.71565
R2616 VTAIL.n400 VTAIL.n385 2.71565
R2617 VTAIL.n356 VTAIL.n355 2.71565
R2618 VTAIL.n338 VTAIL.n281 2.71565
R2619 VTAIL.n310 VTAIL.n295 2.71565
R2620 VTAIL.n666 VTAIL.n665 1.93989
R2621 VTAIL.n698 VTAIL.n638 1.93989
R2622 VTAIL.n712 VTAIL.n632 1.93989
R2623 VTAIL.n36 VTAIL.n35 1.93989
R2624 VTAIL.n68 VTAIL.n8 1.93989
R2625 VTAIL.n82 VTAIL.n2 1.93989
R2626 VTAIL.n126 VTAIL.n125 1.93989
R2627 VTAIL.n158 VTAIL.n98 1.93989
R2628 VTAIL.n172 VTAIL.n92 1.93989
R2629 VTAIL.n216 VTAIL.n215 1.93989
R2630 VTAIL.n248 VTAIL.n188 1.93989
R2631 VTAIL.n262 VTAIL.n182 1.93989
R2632 VTAIL.n622 VTAIL.n542 1.93989
R2633 VTAIL.n609 VTAIL.n549 1.93989
R2634 VTAIL.n577 VTAIL.n576 1.93989
R2635 VTAIL.n532 VTAIL.n452 1.93989
R2636 VTAIL.n519 VTAIL.n459 1.93989
R2637 VTAIL.n487 VTAIL.n486 1.93989
R2638 VTAIL.n442 VTAIL.n362 1.93989
R2639 VTAIL.n429 VTAIL.n369 1.93989
R2640 VTAIL.n397 VTAIL.n396 1.93989
R2641 VTAIL.n352 VTAIL.n272 1.93989
R2642 VTAIL.n339 VTAIL.n279 1.93989
R2643 VTAIL.n307 VTAIL.n306 1.93989
R2644 VTAIL VTAIL.n89 1.73541
R2645 VTAIL VTAIL.n719 1.61903
R2646 VTAIL.n662 VTAIL.n656 1.16414
R2647 VTAIL.n703 VTAIL.n701 1.16414
R2648 VTAIL.n711 VTAIL.n634 1.16414
R2649 VTAIL.n32 VTAIL.n26 1.16414
R2650 VTAIL.n73 VTAIL.n71 1.16414
R2651 VTAIL.n81 VTAIL.n4 1.16414
R2652 VTAIL.n122 VTAIL.n116 1.16414
R2653 VTAIL.n163 VTAIL.n161 1.16414
R2654 VTAIL.n171 VTAIL.n94 1.16414
R2655 VTAIL.n212 VTAIL.n206 1.16414
R2656 VTAIL.n253 VTAIL.n251 1.16414
R2657 VTAIL.n261 VTAIL.n184 1.16414
R2658 VTAIL.n621 VTAIL.n544 1.16414
R2659 VTAIL.n613 VTAIL.n612 1.16414
R2660 VTAIL.n573 VTAIL.n567 1.16414
R2661 VTAIL.n531 VTAIL.n454 1.16414
R2662 VTAIL.n523 VTAIL.n522 1.16414
R2663 VTAIL.n483 VTAIL.n477 1.16414
R2664 VTAIL.n441 VTAIL.n364 1.16414
R2665 VTAIL.n433 VTAIL.n432 1.16414
R2666 VTAIL.n393 VTAIL.n387 1.16414
R2667 VTAIL.n351 VTAIL.n274 1.16414
R2668 VTAIL.n343 VTAIL.n342 1.16414
R2669 VTAIL.n303 VTAIL.n297 1.16414
R2670 VTAIL.n539 VTAIL.n449 0.470328
R2671 VTAIL.n179 VTAIL.n89 0.470328
R2672 VTAIL.n661 VTAIL.n658 0.388379
R2673 VTAIL.n702 VTAIL.n636 0.388379
R2674 VTAIL.n708 VTAIL.n707 0.388379
R2675 VTAIL.n31 VTAIL.n28 0.388379
R2676 VTAIL.n72 VTAIL.n6 0.388379
R2677 VTAIL.n78 VTAIL.n77 0.388379
R2678 VTAIL.n121 VTAIL.n118 0.388379
R2679 VTAIL.n162 VTAIL.n96 0.388379
R2680 VTAIL.n168 VTAIL.n167 0.388379
R2681 VTAIL.n211 VTAIL.n208 0.388379
R2682 VTAIL.n252 VTAIL.n186 0.388379
R2683 VTAIL.n258 VTAIL.n257 0.388379
R2684 VTAIL.n618 VTAIL.n617 0.388379
R2685 VTAIL.n548 VTAIL.n546 0.388379
R2686 VTAIL.n572 VTAIL.n569 0.388379
R2687 VTAIL.n528 VTAIL.n527 0.388379
R2688 VTAIL.n458 VTAIL.n456 0.388379
R2689 VTAIL.n482 VTAIL.n479 0.388379
R2690 VTAIL.n438 VTAIL.n437 0.388379
R2691 VTAIL.n368 VTAIL.n366 0.388379
R2692 VTAIL.n392 VTAIL.n389 0.388379
R2693 VTAIL.n348 VTAIL.n347 0.388379
R2694 VTAIL.n278 VTAIL.n276 0.388379
R2695 VTAIL.n302 VTAIL.n299 0.388379
R2696 VTAIL.n660 VTAIL.n655 0.155672
R2697 VTAIL.n667 VTAIL.n655 0.155672
R2698 VTAIL.n668 VTAIL.n667 0.155672
R2699 VTAIL.n668 VTAIL.n651 0.155672
R2700 VTAIL.n675 VTAIL.n651 0.155672
R2701 VTAIL.n676 VTAIL.n675 0.155672
R2702 VTAIL.n676 VTAIL.n647 0.155672
R2703 VTAIL.n683 VTAIL.n647 0.155672
R2704 VTAIL.n684 VTAIL.n683 0.155672
R2705 VTAIL.n684 VTAIL.n643 0.155672
R2706 VTAIL.n691 VTAIL.n643 0.155672
R2707 VTAIL.n692 VTAIL.n691 0.155672
R2708 VTAIL.n692 VTAIL.n639 0.155672
R2709 VTAIL.n699 VTAIL.n639 0.155672
R2710 VTAIL.n700 VTAIL.n699 0.155672
R2711 VTAIL.n700 VTAIL.n635 0.155672
R2712 VTAIL.n709 VTAIL.n635 0.155672
R2713 VTAIL.n710 VTAIL.n709 0.155672
R2714 VTAIL.n710 VTAIL.n631 0.155672
R2715 VTAIL.n717 VTAIL.n631 0.155672
R2716 VTAIL.n30 VTAIL.n25 0.155672
R2717 VTAIL.n37 VTAIL.n25 0.155672
R2718 VTAIL.n38 VTAIL.n37 0.155672
R2719 VTAIL.n38 VTAIL.n21 0.155672
R2720 VTAIL.n45 VTAIL.n21 0.155672
R2721 VTAIL.n46 VTAIL.n45 0.155672
R2722 VTAIL.n46 VTAIL.n17 0.155672
R2723 VTAIL.n53 VTAIL.n17 0.155672
R2724 VTAIL.n54 VTAIL.n53 0.155672
R2725 VTAIL.n54 VTAIL.n13 0.155672
R2726 VTAIL.n61 VTAIL.n13 0.155672
R2727 VTAIL.n62 VTAIL.n61 0.155672
R2728 VTAIL.n62 VTAIL.n9 0.155672
R2729 VTAIL.n69 VTAIL.n9 0.155672
R2730 VTAIL.n70 VTAIL.n69 0.155672
R2731 VTAIL.n70 VTAIL.n5 0.155672
R2732 VTAIL.n79 VTAIL.n5 0.155672
R2733 VTAIL.n80 VTAIL.n79 0.155672
R2734 VTAIL.n80 VTAIL.n1 0.155672
R2735 VTAIL.n87 VTAIL.n1 0.155672
R2736 VTAIL.n120 VTAIL.n115 0.155672
R2737 VTAIL.n127 VTAIL.n115 0.155672
R2738 VTAIL.n128 VTAIL.n127 0.155672
R2739 VTAIL.n128 VTAIL.n111 0.155672
R2740 VTAIL.n135 VTAIL.n111 0.155672
R2741 VTAIL.n136 VTAIL.n135 0.155672
R2742 VTAIL.n136 VTAIL.n107 0.155672
R2743 VTAIL.n143 VTAIL.n107 0.155672
R2744 VTAIL.n144 VTAIL.n143 0.155672
R2745 VTAIL.n144 VTAIL.n103 0.155672
R2746 VTAIL.n151 VTAIL.n103 0.155672
R2747 VTAIL.n152 VTAIL.n151 0.155672
R2748 VTAIL.n152 VTAIL.n99 0.155672
R2749 VTAIL.n159 VTAIL.n99 0.155672
R2750 VTAIL.n160 VTAIL.n159 0.155672
R2751 VTAIL.n160 VTAIL.n95 0.155672
R2752 VTAIL.n169 VTAIL.n95 0.155672
R2753 VTAIL.n170 VTAIL.n169 0.155672
R2754 VTAIL.n170 VTAIL.n91 0.155672
R2755 VTAIL.n177 VTAIL.n91 0.155672
R2756 VTAIL.n210 VTAIL.n205 0.155672
R2757 VTAIL.n217 VTAIL.n205 0.155672
R2758 VTAIL.n218 VTAIL.n217 0.155672
R2759 VTAIL.n218 VTAIL.n201 0.155672
R2760 VTAIL.n225 VTAIL.n201 0.155672
R2761 VTAIL.n226 VTAIL.n225 0.155672
R2762 VTAIL.n226 VTAIL.n197 0.155672
R2763 VTAIL.n233 VTAIL.n197 0.155672
R2764 VTAIL.n234 VTAIL.n233 0.155672
R2765 VTAIL.n234 VTAIL.n193 0.155672
R2766 VTAIL.n241 VTAIL.n193 0.155672
R2767 VTAIL.n242 VTAIL.n241 0.155672
R2768 VTAIL.n242 VTAIL.n189 0.155672
R2769 VTAIL.n249 VTAIL.n189 0.155672
R2770 VTAIL.n250 VTAIL.n249 0.155672
R2771 VTAIL.n250 VTAIL.n185 0.155672
R2772 VTAIL.n259 VTAIL.n185 0.155672
R2773 VTAIL.n260 VTAIL.n259 0.155672
R2774 VTAIL.n260 VTAIL.n181 0.155672
R2775 VTAIL.n267 VTAIL.n181 0.155672
R2776 VTAIL.n627 VTAIL.n541 0.155672
R2777 VTAIL.n620 VTAIL.n541 0.155672
R2778 VTAIL.n620 VTAIL.n619 0.155672
R2779 VTAIL.n619 VTAIL.n545 0.155672
R2780 VTAIL.n611 VTAIL.n545 0.155672
R2781 VTAIL.n611 VTAIL.n610 0.155672
R2782 VTAIL.n610 VTAIL.n550 0.155672
R2783 VTAIL.n603 VTAIL.n550 0.155672
R2784 VTAIL.n603 VTAIL.n602 0.155672
R2785 VTAIL.n602 VTAIL.n554 0.155672
R2786 VTAIL.n595 VTAIL.n554 0.155672
R2787 VTAIL.n595 VTAIL.n594 0.155672
R2788 VTAIL.n594 VTAIL.n558 0.155672
R2789 VTAIL.n587 VTAIL.n558 0.155672
R2790 VTAIL.n587 VTAIL.n586 0.155672
R2791 VTAIL.n586 VTAIL.n562 0.155672
R2792 VTAIL.n579 VTAIL.n562 0.155672
R2793 VTAIL.n579 VTAIL.n578 0.155672
R2794 VTAIL.n578 VTAIL.n566 0.155672
R2795 VTAIL.n571 VTAIL.n566 0.155672
R2796 VTAIL.n537 VTAIL.n451 0.155672
R2797 VTAIL.n530 VTAIL.n451 0.155672
R2798 VTAIL.n530 VTAIL.n529 0.155672
R2799 VTAIL.n529 VTAIL.n455 0.155672
R2800 VTAIL.n521 VTAIL.n455 0.155672
R2801 VTAIL.n521 VTAIL.n520 0.155672
R2802 VTAIL.n520 VTAIL.n460 0.155672
R2803 VTAIL.n513 VTAIL.n460 0.155672
R2804 VTAIL.n513 VTAIL.n512 0.155672
R2805 VTAIL.n512 VTAIL.n464 0.155672
R2806 VTAIL.n505 VTAIL.n464 0.155672
R2807 VTAIL.n505 VTAIL.n504 0.155672
R2808 VTAIL.n504 VTAIL.n468 0.155672
R2809 VTAIL.n497 VTAIL.n468 0.155672
R2810 VTAIL.n497 VTAIL.n496 0.155672
R2811 VTAIL.n496 VTAIL.n472 0.155672
R2812 VTAIL.n489 VTAIL.n472 0.155672
R2813 VTAIL.n489 VTAIL.n488 0.155672
R2814 VTAIL.n488 VTAIL.n476 0.155672
R2815 VTAIL.n481 VTAIL.n476 0.155672
R2816 VTAIL.n447 VTAIL.n361 0.155672
R2817 VTAIL.n440 VTAIL.n361 0.155672
R2818 VTAIL.n440 VTAIL.n439 0.155672
R2819 VTAIL.n439 VTAIL.n365 0.155672
R2820 VTAIL.n431 VTAIL.n365 0.155672
R2821 VTAIL.n431 VTAIL.n430 0.155672
R2822 VTAIL.n430 VTAIL.n370 0.155672
R2823 VTAIL.n423 VTAIL.n370 0.155672
R2824 VTAIL.n423 VTAIL.n422 0.155672
R2825 VTAIL.n422 VTAIL.n374 0.155672
R2826 VTAIL.n415 VTAIL.n374 0.155672
R2827 VTAIL.n415 VTAIL.n414 0.155672
R2828 VTAIL.n414 VTAIL.n378 0.155672
R2829 VTAIL.n407 VTAIL.n378 0.155672
R2830 VTAIL.n407 VTAIL.n406 0.155672
R2831 VTAIL.n406 VTAIL.n382 0.155672
R2832 VTAIL.n399 VTAIL.n382 0.155672
R2833 VTAIL.n399 VTAIL.n398 0.155672
R2834 VTAIL.n398 VTAIL.n386 0.155672
R2835 VTAIL.n391 VTAIL.n386 0.155672
R2836 VTAIL.n357 VTAIL.n271 0.155672
R2837 VTAIL.n350 VTAIL.n271 0.155672
R2838 VTAIL.n350 VTAIL.n349 0.155672
R2839 VTAIL.n349 VTAIL.n275 0.155672
R2840 VTAIL.n341 VTAIL.n275 0.155672
R2841 VTAIL.n341 VTAIL.n340 0.155672
R2842 VTAIL.n340 VTAIL.n280 0.155672
R2843 VTAIL.n333 VTAIL.n280 0.155672
R2844 VTAIL.n333 VTAIL.n332 0.155672
R2845 VTAIL.n332 VTAIL.n284 0.155672
R2846 VTAIL.n325 VTAIL.n284 0.155672
R2847 VTAIL.n325 VTAIL.n324 0.155672
R2848 VTAIL.n324 VTAIL.n288 0.155672
R2849 VTAIL.n317 VTAIL.n288 0.155672
R2850 VTAIL.n317 VTAIL.n316 0.155672
R2851 VTAIL.n316 VTAIL.n292 0.155672
R2852 VTAIL.n309 VTAIL.n292 0.155672
R2853 VTAIL.n309 VTAIL.n308 0.155672
R2854 VTAIL.n308 VTAIL.n296 0.155672
R2855 VTAIL.n301 VTAIL.n296 0.155672
R2856 VDD1 VDD1.n1 107.32
R2857 VDD1 VDD1.n0 59.2842
R2858 VDD1.n0 VDD1.t1 1.238
R2859 VDD1.n0 VDD1.t3 1.238
R2860 VDD1.n1 VDD1.t0 1.238
R2861 VDD1.n1 VDD1.t2 1.238
R2862 VN.n1 VN.t3 143.103
R2863 VN.n0 VN.t0 143.103
R2864 VN.n0 VN.t2 141.869
R2865 VN.n1 VN.t1 141.869
R2866 VN VN.n1 54.6506
R2867 VN VN.n0 2.1317
R2868 VDD2.n2 VDD2.n0 106.794
R2869 VDD2.n2 VDD2.n1 59.226
R2870 VDD2.n1 VDD2.t2 1.238
R2871 VDD2.n1 VDD2.t0 1.238
R2872 VDD2.n0 VDD2.t3 1.238
R2873 VDD2.n0 VDD2.t1 1.238
R2874 VDD2 VDD2.n2 0.0586897
C0 VDD1 VN 0.150352f
C1 VDD2 VP 0.455877f
C2 VDD1 VTAIL 6.511549f
C3 VDD2 VN 6.54116f
C4 VDD2 VTAIL 6.57219f
C5 VDD1 VDD2 1.25721f
C6 VN VP 7.61882f
C7 VTAIL VP 6.42284f
C8 VN VTAIL 6.40874f
C9 VDD1 VP 6.8457f
C10 VDD2 B 4.626031f
C11 VDD1 B 9.47387f
C12 VTAIL B 13.033222f
C13 VN B 12.85069f
C14 VP B 11.245019f
C15 VDD2.t3 B 0.33882f
C16 VDD2.t1 B 0.33882f
C17 VDD2.n0 B 3.96414f
C18 VDD2.t2 B 0.33882f
C19 VDD2.t0 B 0.33882f
C20 VDD2.n1 B 3.06923f
C21 VDD2.n2 B 4.416009f
C22 VN.t2 B 3.38016f
C23 VN.t0 B 3.39028f
C24 VN.n0 B 2.05149f
C25 VN.t3 B 3.39028f
C26 VN.t1 B 3.38016f
C27 VN.n1 B 3.41735f
C28 VDD1.t1 B 0.341413f
C29 VDD1.t3 B 0.341413f
C30 VDD1.n0 B 3.09325f
C31 VDD1.t0 B 0.341413f
C32 VDD1.t2 B 0.341413f
C33 VDD1.n1 B 4.02367f
C34 VTAIL.n0 B 0.02037f
C35 VTAIL.n1 B 0.016031f
C36 VTAIL.n2 B 0.008614f
C37 VTAIL.n3 B 0.020361f
C38 VTAIL.n4 B 0.009121f
C39 VTAIL.n5 B 0.016031f
C40 VTAIL.n6 B 0.008868f
C41 VTAIL.n7 B 0.020361f
C42 VTAIL.n8 B 0.009121f
C43 VTAIL.n9 B 0.016031f
C44 VTAIL.n10 B 0.008614f
C45 VTAIL.n11 B 0.020361f
C46 VTAIL.n12 B 0.009121f
C47 VTAIL.n13 B 0.016031f
C48 VTAIL.n14 B 0.008614f
C49 VTAIL.n15 B 0.020361f
C50 VTAIL.n16 B 0.009121f
C51 VTAIL.n17 B 0.016031f
C52 VTAIL.n18 B 0.008614f
C53 VTAIL.n19 B 0.020361f
C54 VTAIL.n20 B 0.009121f
C55 VTAIL.n21 B 0.016031f
C56 VTAIL.n22 B 0.008614f
C57 VTAIL.n23 B 0.020361f
C58 VTAIL.n24 B 0.009121f
C59 VTAIL.n25 B 0.016031f
C60 VTAIL.n26 B 0.008614f
C61 VTAIL.n27 B 0.015271f
C62 VTAIL.n28 B 0.012028f
C63 VTAIL.t0 B 0.033628f
C64 VTAIL.n29 B 0.108576f
C65 VTAIL.n30 B 1.11646f
C66 VTAIL.n31 B 0.008614f
C67 VTAIL.n32 B 0.009121f
C68 VTAIL.n33 B 0.020361f
C69 VTAIL.n34 B 0.020361f
C70 VTAIL.n35 B 0.009121f
C71 VTAIL.n36 B 0.008614f
C72 VTAIL.n37 B 0.016031f
C73 VTAIL.n38 B 0.016031f
C74 VTAIL.n39 B 0.008614f
C75 VTAIL.n40 B 0.009121f
C76 VTAIL.n41 B 0.020361f
C77 VTAIL.n42 B 0.020361f
C78 VTAIL.n43 B 0.009121f
C79 VTAIL.n44 B 0.008614f
C80 VTAIL.n45 B 0.016031f
C81 VTAIL.n46 B 0.016031f
C82 VTAIL.n47 B 0.008614f
C83 VTAIL.n48 B 0.009121f
C84 VTAIL.n49 B 0.020361f
C85 VTAIL.n50 B 0.020361f
C86 VTAIL.n51 B 0.009121f
C87 VTAIL.n52 B 0.008614f
C88 VTAIL.n53 B 0.016031f
C89 VTAIL.n54 B 0.016031f
C90 VTAIL.n55 B 0.008614f
C91 VTAIL.n56 B 0.009121f
C92 VTAIL.n57 B 0.020361f
C93 VTAIL.n58 B 0.020361f
C94 VTAIL.n59 B 0.009121f
C95 VTAIL.n60 B 0.008614f
C96 VTAIL.n61 B 0.016031f
C97 VTAIL.n62 B 0.016031f
C98 VTAIL.n63 B 0.008614f
C99 VTAIL.n64 B 0.009121f
C100 VTAIL.n65 B 0.020361f
C101 VTAIL.n66 B 0.020361f
C102 VTAIL.n67 B 0.009121f
C103 VTAIL.n68 B 0.008614f
C104 VTAIL.n69 B 0.016031f
C105 VTAIL.n70 B 0.016031f
C106 VTAIL.n71 B 0.008614f
C107 VTAIL.n72 B 0.008614f
C108 VTAIL.n73 B 0.009121f
C109 VTAIL.n74 B 0.020361f
C110 VTAIL.n75 B 0.020361f
C111 VTAIL.n76 B 0.020361f
C112 VTAIL.n77 B 0.008868f
C113 VTAIL.n78 B 0.008614f
C114 VTAIL.n79 B 0.016031f
C115 VTAIL.n80 B 0.016031f
C116 VTAIL.n81 B 0.008614f
C117 VTAIL.n82 B 0.009121f
C118 VTAIL.n83 B 0.020361f
C119 VTAIL.n84 B 0.040253f
C120 VTAIL.n85 B 0.009121f
C121 VTAIL.n86 B 0.008614f
C122 VTAIL.n87 B 0.035303f
C123 VTAIL.n88 B 0.022075f
C124 VTAIL.n89 B 0.12659f
C125 VTAIL.n90 B 0.02037f
C126 VTAIL.n91 B 0.016031f
C127 VTAIL.n92 B 0.008614f
C128 VTAIL.n93 B 0.020361f
C129 VTAIL.n94 B 0.009121f
C130 VTAIL.n95 B 0.016031f
C131 VTAIL.n96 B 0.008868f
C132 VTAIL.n97 B 0.020361f
C133 VTAIL.n98 B 0.009121f
C134 VTAIL.n99 B 0.016031f
C135 VTAIL.n100 B 0.008614f
C136 VTAIL.n101 B 0.020361f
C137 VTAIL.n102 B 0.009121f
C138 VTAIL.n103 B 0.016031f
C139 VTAIL.n104 B 0.008614f
C140 VTAIL.n105 B 0.020361f
C141 VTAIL.n106 B 0.009121f
C142 VTAIL.n107 B 0.016031f
C143 VTAIL.n108 B 0.008614f
C144 VTAIL.n109 B 0.020361f
C145 VTAIL.n110 B 0.009121f
C146 VTAIL.n111 B 0.016031f
C147 VTAIL.n112 B 0.008614f
C148 VTAIL.n113 B 0.020361f
C149 VTAIL.n114 B 0.009121f
C150 VTAIL.n115 B 0.016031f
C151 VTAIL.n116 B 0.008614f
C152 VTAIL.n117 B 0.015271f
C153 VTAIL.n118 B 0.012028f
C154 VTAIL.t4 B 0.033628f
C155 VTAIL.n119 B 0.108576f
C156 VTAIL.n120 B 1.11646f
C157 VTAIL.n121 B 0.008614f
C158 VTAIL.n122 B 0.009121f
C159 VTAIL.n123 B 0.020361f
C160 VTAIL.n124 B 0.020361f
C161 VTAIL.n125 B 0.009121f
C162 VTAIL.n126 B 0.008614f
C163 VTAIL.n127 B 0.016031f
C164 VTAIL.n128 B 0.016031f
C165 VTAIL.n129 B 0.008614f
C166 VTAIL.n130 B 0.009121f
C167 VTAIL.n131 B 0.020361f
C168 VTAIL.n132 B 0.020361f
C169 VTAIL.n133 B 0.009121f
C170 VTAIL.n134 B 0.008614f
C171 VTAIL.n135 B 0.016031f
C172 VTAIL.n136 B 0.016031f
C173 VTAIL.n137 B 0.008614f
C174 VTAIL.n138 B 0.009121f
C175 VTAIL.n139 B 0.020361f
C176 VTAIL.n140 B 0.020361f
C177 VTAIL.n141 B 0.009121f
C178 VTAIL.n142 B 0.008614f
C179 VTAIL.n143 B 0.016031f
C180 VTAIL.n144 B 0.016031f
C181 VTAIL.n145 B 0.008614f
C182 VTAIL.n146 B 0.009121f
C183 VTAIL.n147 B 0.020361f
C184 VTAIL.n148 B 0.020361f
C185 VTAIL.n149 B 0.009121f
C186 VTAIL.n150 B 0.008614f
C187 VTAIL.n151 B 0.016031f
C188 VTAIL.n152 B 0.016031f
C189 VTAIL.n153 B 0.008614f
C190 VTAIL.n154 B 0.009121f
C191 VTAIL.n155 B 0.020361f
C192 VTAIL.n156 B 0.020361f
C193 VTAIL.n157 B 0.009121f
C194 VTAIL.n158 B 0.008614f
C195 VTAIL.n159 B 0.016031f
C196 VTAIL.n160 B 0.016031f
C197 VTAIL.n161 B 0.008614f
C198 VTAIL.n162 B 0.008614f
C199 VTAIL.n163 B 0.009121f
C200 VTAIL.n164 B 0.020361f
C201 VTAIL.n165 B 0.020361f
C202 VTAIL.n166 B 0.020361f
C203 VTAIL.n167 B 0.008868f
C204 VTAIL.n168 B 0.008614f
C205 VTAIL.n169 B 0.016031f
C206 VTAIL.n170 B 0.016031f
C207 VTAIL.n171 B 0.008614f
C208 VTAIL.n172 B 0.009121f
C209 VTAIL.n173 B 0.020361f
C210 VTAIL.n174 B 0.040253f
C211 VTAIL.n175 B 0.009121f
C212 VTAIL.n176 B 0.008614f
C213 VTAIL.n177 B 0.035303f
C214 VTAIL.n178 B 0.022075f
C215 VTAIL.n179 B 0.210195f
C216 VTAIL.n180 B 0.02037f
C217 VTAIL.n181 B 0.016031f
C218 VTAIL.n182 B 0.008614f
C219 VTAIL.n183 B 0.020361f
C220 VTAIL.n184 B 0.009121f
C221 VTAIL.n185 B 0.016031f
C222 VTAIL.n186 B 0.008868f
C223 VTAIL.n187 B 0.020361f
C224 VTAIL.n188 B 0.009121f
C225 VTAIL.n189 B 0.016031f
C226 VTAIL.n190 B 0.008614f
C227 VTAIL.n191 B 0.020361f
C228 VTAIL.n192 B 0.009121f
C229 VTAIL.n193 B 0.016031f
C230 VTAIL.n194 B 0.008614f
C231 VTAIL.n195 B 0.020361f
C232 VTAIL.n196 B 0.009121f
C233 VTAIL.n197 B 0.016031f
C234 VTAIL.n198 B 0.008614f
C235 VTAIL.n199 B 0.020361f
C236 VTAIL.n200 B 0.009121f
C237 VTAIL.n201 B 0.016031f
C238 VTAIL.n202 B 0.008614f
C239 VTAIL.n203 B 0.020361f
C240 VTAIL.n204 B 0.009121f
C241 VTAIL.n205 B 0.016031f
C242 VTAIL.n206 B 0.008614f
C243 VTAIL.n207 B 0.015271f
C244 VTAIL.n208 B 0.012028f
C245 VTAIL.t6 B 0.033628f
C246 VTAIL.n209 B 0.108576f
C247 VTAIL.n210 B 1.11646f
C248 VTAIL.n211 B 0.008614f
C249 VTAIL.n212 B 0.009121f
C250 VTAIL.n213 B 0.020361f
C251 VTAIL.n214 B 0.020361f
C252 VTAIL.n215 B 0.009121f
C253 VTAIL.n216 B 0.008614f
C254 VTAIL.n217 B 0.016031f
C255 VTAIL.n218 B 0.016031f
C256 VTAIL.n219 B 0.008614f
C257 VTAIL.n220 B 0.009121f
C258 VTAIL.n221 B 0.020361f
C259 VTAIL.n222 B 0.020361f
C260 VTAIL.n223 B 0.009121f
C261 VTAIL.n224 B 0.008614f
C262 VTAIL.n225 B 0.016031f
C263 VTAIL.n226 B 0.016031f
C264 VTAIL.n227 B 0.008614f
C265 VTAIL.n228 B 0.009121f
C266 VTAIL.n229 B 0.020361f
C267 VTAIL.n230 B 0.020361f
C268 VTAIL.n231 B 0.009121f
C269 VTAIL.n232 B 0.008614f
C270 VTAIL.n233 B 0.016031f
C271 VTAIL.n234 B 0.016031f
C272 VTAIL.n235 B 0.008614f
C273 VTAIL.n236 B 0.009121f
C274 VTAIL.n237 B 0.020361f
C275 VTAIL.n238 B 0.020361f
C276 VTAIL.n239 B 0.009121f
C277 VTAIL.n240 B 0.008614f
C278 VTAIL.n241 B 0.016031f
C279 VTAIL.n242 B 0.016031f
C280 VTAIL.n243 B 0.008614f
C281 VTAIL.n244 B 0.009121f
C282 VTAIL.n245 B 0.020361f
C283 VTAIL.n246 B 0.020361f
C284 VTAIL.n247 B 0.009121f
C285 VTAIL.n248 B 0.008614f
C286 VTAIL.n249 B 0.016031f
C287 VTAIL.n250 B 0.016031f
C288 VTAIL.n251 B 0.008614f
C289 VTAIL.n252 B 0.008614f
C290 VTAIL.n253 B 0.009121f
C291 VTAIL.n254 B 0.020361f
C292 VTAIL.n255 B 0.020361f
C293 VTAIL.n256 B 0.020361f
C294 VTAIL.n257 B 0.008868f
C295 VTAIL.n258 B 0.008614f
C296 VTAIL.n259 B 0.016031f
C297 VTAIL.n260 B 0.016031f
C298 VTAIL.n261 B 0.008614f
C299 VTAIL.n262 B 0.009121f
C300 VTAIL.n263 B 0.020361f
C301 VTAIL.n264 B 0.040253f
C302 VTAIL.n265 B 0.009121f
C303 VTAIL.n266 B 0.008614f
C304 VTAIL.n267 B 0.035303f
C305 VTAIL.n268 B 0.022075f
C306 VTAIL.n269 B 1.28939f
C307 VTAIL.n270 B 0.02037f
C308 VTAIL.n271 B 0.016031f
C309 VTAIL.n272 B 0.008614f
C310 VTAIL.n273 B 0.020361f
C311 VTAIL.n274 B 0.009121f
C312 VTAIL.n275 B 0.016031f
C313 VTAIL.n276 B 0.008868f
C314 VTAIL.n277 B 0.020361f
C315 VTAIL.n278 B 0.008614f
C316 VTAIL.n279 B 0.009121f
C317 VTAIL.n280 B 0.016031f
C318 VTAIL.n281 B 0.008614f
C319 VTAIL.n282 B 0.020361f
C320 VTAIL.n283 B 0.009121f
C321 VTAIL.n284 B 0.016031f
C322 VTAIL.n285 B 0.008614f
C323 VTAIL.n286 B 0.020361f
C324 VTAIL.n287 B 0.009121f
C325 VTAIL.n288 B 0.016031f
C326 VTAIL.n289 B 0.008614f
C327 VTAIL.n290 B 0.020361f
C328 VTAIL.n291 B 0.009121f
C329 VTAIL.n292 B 0.016031f
C330 VTAIL.n293 B 0.008614f
C331 VTAIL.n294 B 0.020361f
C332 VTAIL.n295 B 0.009121f
C333 VTAIL.n296 B 0.016031f
C334 VTAIL.n297 B 0.008614f
C335 VTAIL.n298 B 0.015271f
C336 VTAIL.n299 B 0.012028f
C337 VTAIL.t1 B 0.033628f
C338 VTAIL.n300 B 0.108576f
C339 VTAIL.n301 B 1.11646f
C340 VTAIL.n302 B 0.008614f
C341 VTAIL.n303 B 0.009121f
C342 VTAIL.n304 B 0.020361f
C343 VTAIL.n305 B 0.020361f
C344 VTAIL.n306 B 0.009121f
C345 VTAIL.n307 B 0.008614f
C346 VTAIL.n308 B 0.016031f
C347 VTAIL.n309 B 0.016031f
C348 VTAIL.n310 B 0.008614f
C349 VTAIL.n311 B 0.009121f
C350 VTAIL.n312 B 0.020361f
C351 VTAIL.n313 B 0.020361f
C352 VTAIL.n314 B 0.009121f
C353 VTAIL.n315 B 0.008614f
C354 VTAIL.n316 B 0.016031f
C355 VTAIL.n317 B 0.016031f
C356 VTAIL.n318 B 0.008614f
C357 VTAIL.n319 B 0.009121f
C358 VTAIL.n320 B 0.020361f
C359 VTAIL.n321 B 0.020361f
C360 VTAIL.n322 B 0.009121f
C361 VTAIL.n323 B 0.008614f
C362 VTAIL.n324 B 0.016031f
C363 VTAIL.n325 B 0.016031f
C364 VTAIL.n326 B 0.008614f
C365 VTAIL.n327 B 0.009121f
C366 VTAIL.n328 B 0.020361f
C367 VTAIL.n329 B 0.020361f
C368 VTAIL.n330 B 0.009121f
C369 VTAIL.n331 B 0.008614f
C370 VTAIL.n332 B 0.016031f
C371 VTAIL.n333 B 0.016031f
C372 VTAIL.n334 B 0.008614f
C373 VTAIL.n335 B 0.009121f
C374 VTAIL.n336 B 0.020361f
C375 VTAIL.n337 B 0.020361f
C376 VTAIL.n338 B 0.009121f
C377 VTAIL.n339 B 0.008614f
C378 VTAIL.n340 B 0.016031f
C379 VTAIL.n341 B 0.016031f
C380 VTAIL.n342 B 0.008614f
C381 VTAIL.n343 B 0.009121f
C382 VTAIL.n344 B 0.020361f
C383 VTAIL.n345 B 0.020361f
C384 VTAIL.n346 B 0.020361f
C385 VTAIL.n347 B 0.008868f
C386 VTAIL.n348 B 0.008614f
C387 VTAIL.n349 B 0.016031f
C388 VTAIL.n350 B 0.016031f
C389 VTAIL.n351 B 0.008614f
C390 VTAIL.n352 B 0.009121f
C391 VTAIL.n353 B 0.020361f
C392 VTAIL.n354 B 0.040253f
C393 VTAIL.n355 B 0.009121f
C394 VTAIL.n356 B 0.008614f
C395 VTAIL.n357 B 0.035303f
C396 VTAIL.n358 B 0.022075f
C397 VTAIL.n359 B 1.28939f
C398 VTAIL.n360 B 0.02037f
C399 VTAIL.n361 B 0.016031f
C400 VTAIL.n362 B 0.008614f
C401 VTAIL.n363 B 0.020361f
C402 VTAIL.n364 B 0.009121f
C403 VTAIL.n365 B 0.016031f
C404 VTAIL.n366 B 0.008868f
C405 VTAIL.n367 B 0.020361f
C406 VTAIL.n368 B 0.008614f
C407 VTAIL.n369 B 0.009121f
C408 VTAIL.n370 B 0.016031f
C409 VTAIL.n371 B 0.008614f
C410 VTAIL.n372 B 0.020361f
C411 VTAIL.n373 B 0.009121f
C412 VTAIL.n374 B 0.016031f
C413 VTAIL.n375 B 0.008614f
C414 VTAIL.n376 B 0.020361f
C415 VTAIL.n377 B 0.009121f
C416 VTAIL.n378 B 0.016031f
C417 VTAIL.n379 B 0.008614f
C418 VTAIL.n380 B 0.020361f
C419 VTAIL.n381 B 0.009121f
C420 VTAIL.n382 B 0.016031f
C421 VTAIL.n383 B 0.008614f
C422 VTAIL.n384 B 0.020361f
C423 VTAIL.n385 B 0.009121f
C424 VTAIL.n386 B 0.016031f
C425 VTAIL.n387 B 0.008614f
C426 VTAIL.n388 B 0.015271f
C427 VTAIL.n389 B 0.012028f
C428 VTAIL.t3 B 0.033628f
C429 VTAIL.n390 B 0.108576f
C430 VTAIL.n391 B 1.11646f
C431 VTAIL.n392 B 0.008614f
C432 VTAIL.n393 B 0.009121f
C433 VTAIL.n394 B 0.020361f
C434 VTAIL.n395 B 0.020361f
C435 VTAIL.n396 B 0.009121f
C436 VTAIL.n397 B 0.008614f
C437 VTAIL.n398 B 0.016031f
C438 VTAIL.n399 B 0.016031f
C439 VTAIL.n400 B 0.008614f
C440 VTAIL.n401 B 0.009121f
C441 VTAIL.n402 B 0.020361f
C442 VTAIL.n403 B 0.020361f
C443 VTAIL.n404 B 0.009121f
C444 VTAIL.n405 B 0.008614f
C445 VTAIL.n406 B 0.016031f
C446 VTAIL.n407 B 0.016031f
C447 VTAIL.n408 B 0.008614f
C448 VTAIL.n409 B 0.009121f
C449 VTAIL.n410 B 0.020361f
C450 VTAIL.n411 B 0.020361f
C451 VTAIL.n412 B 0.009121f
C452 VTAIL.n413 B 0.008614f
C453 VTAIL.n414 B 0.016031f
C454 VTAIL.n415 B 0.016031f
C455 VTAIL.n416 B 0.008614f
C456 VTAIL.n417 B 0.009121f
C457 VTAIL.n418 B 0.020361f
C458 VTAIL.n419 B 0.020361f
C459 VTAIL.n420 B 0.009121f
C460 VTAIL.n421 B 0.008614f
C461 VTAIL.n422 B 0.016031f
C462 VTAIL.n423 B 0.016031f
C463 VTAIL.n424 B 0.008614f
C464 VTAIL.n425 B 0.009121f
C465 VTAIL.n426 B 0.020361f
C466 VTAIL.n427 B 0.020361f
C467 VTAIL.n428 B 0.009121f
C468 VTAIL.n429 B 0.008614f
C469 VTAIL.n430 B 0.016031f
C470 VTAIL.n431 B 0.016031f
C471 VTAIL.n432 B 0.008614f
C472 VTAIL.n433 B 0.009121f
C473 VTAIL.n434 B 0.020361f
C474 VTAIL.n435 B 0.020361f
C475 VTAIL.n436 B 0.020361f
C476 VTAIL.n437 B 0.008868f
C477 VTAIL.n438 B 0.008614f
C478 VTAIL.n439 B 0.016031f
C479 VTAIL.n440 B 0.016031f
C480 VTAIL.n441 B 0.008614f
C481 VTAIL.n442 B 0.009121f
C482 VTAIL.n443 B 0.020361f
C483 VTAIL.n444 B 0.040253f
C484 VTAIL.n445 B 0.009121f
C485 VTAIL.n446 B 0.008614f
C486 VTAIL.n447 B 0.035303f
C487 VTAIL.n448 B 0.022075f
C488 VTAIL.n449 B 0.210195f
C489 VTAIL.n450 B 0.02037f
C490 VTAIL.n451 B 0.016031f
C491 VTAIL.n452 B 0.008614f
C492 VTAIL.n453 B 0.020361f
C493 VTAIL.n454 B 0.009121f
C494 VTAIL.n455 B 0.016031f
C495 VTAIL.n456 B 0.008868f
C496 VTAIL.n457 B 0.020361f
C497 VTAIL.n458 B 0.008614f
C498 VTAIL.n459 B 0.009121f
C499 VTAIL.n460 B 0.016031f
C500 VTAIL.n461 B 0.008614f
C501 VTAIL.n462 B 0.020361f
C502 VTAIL.n463 B 0.009121f
C503 VTAIL.n464 B 0.016031f
C504 VTAIL.n465 B 0.008614f
C505 VTAIL.n466 B 0.020361f
C506 VTAIL.n467 B 0.009121f
C507 VTAIL.n468 B 0.016031f
C508 VTAIL.n469 B 0.008614f
C509 VTAIL.n470 B 0.020361f
C510 VTAIL.n471 B 0.009121f
C511 VTAIL.n472 B 0.016031f
C512 VTAIL.n473 B 0.008614f
C513 VTAIL.n474 B 0.020361f
C514 VTAIL.n475 B 0.009121f
C515 VTAIL.n476 B 0.016031f
C516 VTAIL.n477 B 0.008614f
C517 VTAIL.n478 B 0.015271f
C518 VTAIL.n479 B 0.012028f
C519 VTAIL.t7 B 0.033628f
C520 VTAIL.n480 B 0.108576f
C521 VTAIL.n481 B 1.11646f
C522 VTAIL.n482 B 0.008614f
C523 VTAIL.n483 B 0.009121f
C524 VTAIL.n484 B 0.020361f
C525 VTAIL.n485 B 0.020361f
C526 VTAIL.n486 B 0.009121f
C527 VTAIL.n487 B 0.008614f
C528 VTAIL.n488 B 0.016031f
C529 VTAIL.n489 B 0.016031f
C530 VTAIL.n490 B 0.008614f
C531 VTAIL.n491 B 0.009121f
C532 VTAIL.n492 B 0.020361f
C533 VTAIL.n493 B 0.020361f
C534 VTAIL.n494 B 0.009121f
C535 VTAIL.n495 B 0.008614f
C536 VTAIL.n496 B 0.016031f
C537 VTAIL.n497 B 0.016031f
C538 VTAIL.n498 B 0.008614f
C539 VTAIL.n499 B 0.009121f
C540 VTAIL.n500 B 0.020361f
C541 VTAIL.n501 B 0.020361f
C542 VTAIL.n502 B 0.009121f
C543 VTAIL.n503 B 0.008614f
C544 VTAIL.n504 B 0.016031f
C545 VTAIL.n505 B 0.016031f
C546 VTAIL.n506 B 0.008614f
C547 VTAIL.n507 B 0.009121f
C548 VTAIL.n508 B 0.020361f
C549 VTAIL.n509 B 0.020361f
C550 VTAIL.n510 B 0.009121f
C551 VTAIL.n511 B 0.008614f
C552 VTAIL.n512 B 0.016031f
C553 VTAIL.n513 B 0.016031f
C554 VTAIL.n514 B 0.008614f
C555 VTAIL.n515 B 0.009121f
C556 VTAIL.n516 B 0.020361f
C557 VTAIL.n517 B 0.020361f
C558 VTAIL.n518 B 0.009121f
C559 VTAIL.n519 B 0.008614f
C560 VTAIL.n520 B 0.016031f
C561 VTAIL.n521 B 0.016031f
C562 VTAIL.n522 B 0.008614f
C563 VTAIL.n523 B 0.009121f
C564 VTAIL.n524 B 0.020361f
C565 VTAIL.n525 B 0.020361f
C566 VTAIL.n526 B 0.020361f
C567 VTAIL.n527 B 0.008868f
C568 VTAIL.n528 B 0.008614f
C569 VTAIL.n529 B 0.016031f
C570 VTAIL.n530 B 0.016031f
C571 VTAIL.n531 B 0.008614f
C572 VTAIL.n532 B 0.009121f
C573 VTAIL.n533 B 0.020361f
C574 VTAIL.n534 B 0.040253f
C575 VTAIL.n535 B 0.009121f
C576 VTAIL.n536 B 0.008614f
C577 VTAIL.n537 B 0.035303f
C578 VTAIL.n538 B 0.022075f
C579 VTAIL.n539 B 0.210195f
C580 VTAIL.n540 B 0.02037f
C581 VTAIL.n541 B 0.016031f
C582 VTAIL.n542 B 0.008614f
C583 VTAIL.n543 B 0.020361f
C584 VTAIL.n544 B 0.009121f
C585 VTAIL.n545 B 0.016031f
C586 VTAIL.n546 B 0.008868f
C587 VTAIL.n547 B 0.020361f
C588 VTAIL.n548 B 0.008614f
C589 VTAIL.n549 B 0.009121f
C590 VTAIL.n550 B 0.016031f
C591 VTAIL.n551 B 0.008614f
C592 VTAIL.n552 B 0.020361f
C593 VTAIL.n553 B 0.009121f
C594 VTAIL.n554 B 0.016031f
C595 VTAIL.n555 B 0.008614f
C596 VTAIL.n556 B 0.020361f
C597 VTAIL.n557 B 0.009121f
C598 VTAIL.n558 B 0.016031f
C599 VTAIL.n559 B 0.008614f
C600 VTAIL.n560 B 0.020361f
C601 VTAIL.n561 B 0.009121f
C602 VTAIL.n562 B 0.016031f
C603 VTAIL.n563 B 0.008614f
C604 VTAIL.n564 B 0.020361f
C605 VTAIL.n565 B 0.009121f
C606 VTAIL.n566 B 0.016031f
C607 VTAIL.n567 B 0.008614f
C608 VTAIL.n568 B 0.015271f
C609 VTAIL.n569 B 0.012028f
C610 VTAIL.t5 B 0.033628f
C611 VTAIL.n570 B 0.108576f
C612 VTAIL.n571 B 1.11646f
C613 VTAIL.n572 B 0.008614f
C614 VTAIL.n573 B 0.009121f
C615 VTAIL.n574 B 0.020361f
C616 VTAIL.n575 B 0.020361f
C617 VTAIL.n576 B 0.009121f
C618 VTAIL.n577 B 0.008614f
C619 VTAIL.n578 B 0.016031f
C620 VTAIL.n579 B 0.016031f
C621 VTAIL.n580 B 0.008614f
C622 VTAIL.n581 B 0.009121f
C623 VTAIL.n582 B 0.020361f
C624 VTAIL.n583 B 0.020361f
C625 VTAIL.n584 B 0.009121f
C626 VTAIL.n585 B 0.008614f
C627 VTAIL.n586 B 0.016031f
C628 VTAIL.n587 B 0.016031f
C629 VTAIL.n588 B 0.008614f
C630 VTAIL.n589 B 0.009121f
C631 VTAIL.n590 B 0.020361f
C632 VTAIL.n591 B 0.020361f
C633 VTAIL.n592 B 0.009121f
C634 VTAIL.n593 B 0.008614f
C635 VTAIL.n594 B 0.016031f
C636 VTAIL.n595 B 0.016031f
C637 VTAIL.n596 B 0.008614f
C638 VTAIL.n597 B 0.009121f
C639 VTAIL.n598 B 0.020361f
C640 VTAIL.n599 B 0.020361f
C641 VTAIL.n600 B 0.009121f
C642 VTAIL.n601 B 0.008614f
C643 VTAIL.n602 B 0.016031f
C644 VTAIL.n603 B 0.016031f
C645 VTAIL.n604 B 0.008614f
C646 VTAIL.n605 B 0.009121f
C647 VTAIL.n606 B 0.020361f
C648 VTAIL.n607 B 0.020361f
C649 VTAIL.n608 B 0.009121f
C650 VTAIL.n609 B 0.008614f
C651 VTAIL.n610 B 0.016031f
C652 VTAIL.n611 B 0.016031f
C653 VTAIL.n612 B 0.008614f
C654 VTAIL.n613 B 0.009121f
C655 VTAIL.n614 B 0.020361f
C656 VTAIL.n615 B 0.020361f
C657 VTAIL.n616 B 0.020361f
C658 VTAIL.n617 B 0.008868f
C659 VTAIL.n618 B 0.008614f
C660 VTAIL.n619 B 0.016031f
C661 VTAIL.n620 B 0.016031f
C662 VTAIL.n621 B 0.008614f
C663 VTAIL.n622 B 0.009121f
C664 VTAIL.n623 B 0.020361f
C665 VTAIL.n624 B 0.040253f
C666 VTAIL.n625 B 0.009121f
C667 VTAIL.n626 B 0.008614f
C668 VTAIL.n627 B 0.035303f
C669 VTAIL.n628 B 0.022075f
C670 VTAIL.n629 B 1.28939f
C671 VTAIL.n630 B 0.02037f
C672 VTAIL.n631 B 0.016031f
C673 VTAIL.n632 B 0.008614f
C674 VTAIL.n633 B 0.020361f
C675 VTAIL.n634 B 0.009121f
C676 VTAIL.n635 B 0.016031f
C677 VTAIL.n636 B 0.008868f
C678 VTAIL.n637 B 0.020361f
C679 VTAIL.n638 B 0.009121f
C680 VTAIL.n639 B 0.016031f
C681 VTAIL.n640 B 0.008614f
C682 VTAIL.n641 B 0.020361f
C683 VTAIL.n642 B 0.009121f
C684 VTAIL.n643 B 0.016031f
C685 VTAIL.n644 B 0.008614f
C686 VTAIL.n645 B 0.020361f
C687 VTAIL.n646 B 0.009121f
C688 VTAIL.n647 B 0.016031f
C689 VTAIL.n648 B 0.008614f
C690 VTAIL.n649 B 0.020361f
C691 VTAIL.n650 B 0.009121f
C692 VTAIL.n651 B 0.016031f
C693 VTAIL.n652 B 0.008614f
C694 VTAIL.n653 B 0.020361f
C695 VTAIL.n654 B 0.009121f
C696 VTAIL.n655 B 0.016031f
C697 VTAIL.n656 B 0.008614f
C698 VTAIL.n657 B 0.015271f
C699 VTAIL.n658 B 0.012028f
C700 VTAIL.t2 B 0.033628f
C701 VTAIL.n659 B 0.108576f
C702 VTAIL.n660 B 1.11646f
C703 VTAIL.n661 B 0.008614f
C704 VTAIL.n662 B 0.009121f
C705 VTAIL.n663 B 0.020361f
C706 VTAIL.n664 B 0.020361f
C707 VTAIL.n665 B 0.009121f
C708 VTAIL.n666 B 0.008614f
C709 VTAIL.n667 B 0.016031f
C710 VTAIL.n668 B 0.016031f
C711 VTAIL.n669 B 0.008614f
C712 VTAIL.n670 B 0.009121f
C713 VTAIL.n671 B 0.020361f
C714 VTAIL.n672 B 0.020361f
C715 VTAIL.n673 B 0.009121f
C716 VTAIL.n674 B 0.008614f
C717 VTAIL.n675 B 0.016031f
C718 VTAIL.n676 B 0.016031f
C719 VTAIL.n677 B 0.008614f
C720 VTAIL.n678 B 0.009121f
C721 VTAIL.n679 B 0.020361f
C722 VTAIL.n680 B 0.020361f
C723 VTAIL.n681 B 0.009121f
C724 VTAIL.n682 B 0.008614f
C725 VTAIL.n683 B 0.016031f
C726 VTAIL.n684 B 0.016031f
C727 VTAIL.n685 B 0.008614f
C728 VTAIL.n686 B 0.009121f
C729 VTAIL.n687 B 0.020361f
C730 VTAIL.n688 B 0.020361f
C731 VTAIL.n689 B 0.009121f
C732 VTAIL.n690 B 0.008614f
C733 VTAIL.n691 B 0.016031f
C734 VTAIL.n692 B 0.016031f
C735 VTAIL.n693 B 0.008614f
C736 VTAIL.n694 B 0.009121f
C737 VTAIL.n695 B 0.020361f
C738 VTAIL.n696 B 0.020361f
C739 VTAIL.n697 B 0.009121f
C740 VTAIL.n698 B 0.008614f
C741 VTAIL.n699 B 0.016031f
C742 VTAIL.n700 B 0.016031f
C743 VTAIL.n701 B 0.008614f
C744 VTAIL.n702 B 0.008614f
C745 VTAIL.n703 B 0.009121f
C746 VTAIL.n704 B 0.020361f
C747 VTAIL.n705 B 0.020361f
C748 VTAIL.n706 B 0.020361f
C749 VTAIL.n707 B 0.008868f
C750 VTAIL.n708 B 0.008614f
C751 VTAIL.n709 B 0.016031f
C752 VTAIL.n710 B 0.016031f
C753 VTAIL.n711 B 0.008614f
C754 VTAIL.n712 B 0.009121f
C755 VTAIL.n713 B 0.020361f
C756 VTAIL.n714 B 0.040253f
C757 VTAIL.n715 B 0.009121f
C758 VTAIL.n716 B 0.008614f
C759 VTAIL.n717 B 0.035303f
C760 VTAIL.n718 B 0.022075f
C761 VTAIL.n719 B 1.19978f
C762 VP.t1 B 3.14176f
C763 VP.n0 B 1.16565f
C764 VP.n1 B 0.020101f
C765 VP.n2 B 0.029219f
C766 VP.n3 B 0.020101f
C767 VP.n4 B 0.02605f
C768 VP.t2 B 3.44457f
C769 VP.t0 B 3.43428f
C770 VP.n5 B 3.46411f
C771 VP.t3 B 3.14176f
C772 VP.n6 B 1.16565f
C773 VP.n7 B 1.30007f
C774 VP.n8 B 0.032437f
C775 VP.n9 B 0.020101f
C776 VP.n10 B 0.037274f
C777 VP.n11 B 0.037274f
C778 VP.n12 B 0.029219f
C779 VP.n13 B 0.020101f
C780 VP.n14 B 0.020101f
C781 VP.n15 B 0.020101f
C782 VP.n16 B 0.037274f
C783 VP.n17 B 0.037274f
C784 VP.n18 B 0.02605f
C785 VP.n19 B 0.032437f
C786 VP.n20 B 0.054824f
.ends

