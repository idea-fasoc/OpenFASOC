* NGSPICE file created from diff_pair_sample_0434.ext - technology: sky130A

.subckt diff_pair_sample_0434 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=3.19605 pd=19.7 as=3.19605 ps=19.7 w=19.37 l=1.58
X1 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=7.5543 pd=39.52 as=0 ps=0 w=19.37 l=1.58
X2 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=7.5543 pd=39.52 as=0 ps=0 w=19.37 l=1.58
X3 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.5543 pd=39.52 as=0 ps=0 w=19.37 l=1.58
X4 VTAIL.t1 VN.t0 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=3.19605 pd=19.7 as=3.19605 ps=19.7 w=19.37 l=1.58
X5 VDD1.t5 VP.t1 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=7.5543 pd=39.52 as=3.19605 ps=19.7 w=19.37 l=1.58
X6 VTAIL.t5 VN.t1 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=3.19605 pd=19.7 as=3.19605 ps=19.7 w=19.37 l=1.58
X7 VTAIL.t9 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.19605 pd=19.7 as=3.19605 ps=19.7 w=19.37 l=1.58
X8 VDD2.t3 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.19605 pd=19.7 as=7.5543 ps=39.52 w=19.37 l=1.58
X9 VDD1.t0 VP.t3 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=3.19605 pd=19.7 as=7.5543 ps=39.52 w=19.37 l=1.58
X10 VDD2.t2 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.19605 pd=19.7 as=7.5543 ps=39.52 w=19.37 l=1.58
X11 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.5543 pd=39.52 as=0 ps=0 w=19.37 l=1.58
X12 VDD2.t1 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=7.5543 pd=39.52 as=3.19605 ps=19.7 w=19.37 l=1.58
X13 VDD1.t2 VP.t4 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=3.19605 pd=19.7 as=7.5543 ps=39.52 w=19.37 l=1.58
X14 VDD1.t4 VP.t5 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=7.5543 pd=39.52 as=3.19605 ps=19.7 w=19.37 l=1.58
X15 VDD2.t0 VN.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=7.5543 pd=39.52 as=3.19605 ps=19.7 w=19.37 l=1.58
R0 VP.n6 VP.t1 328.036
R1 VP.n17 VP.t5 295.454
R2 VP.n24 VP.t2 295.454
R3 VP.n31 VP.t4 295.454
R4 VP.n14 VP.t3 295.454
R5 VP.n7 VP.t0 295.454
R6 VP.n17 VP.n16 177.939
R7 VP.n32 VP.n31 177.939
R8 VP.n15 VP.n14 177.939
R9 VP.n9 VP.n8 161.3
R10 VP.n10 VP.n5 161.3
R11 VP.n12 VP.n11 161.3
R12 VP.n13 VP.n4 161.3
R13 VP.n30 VP.n0 161.3
R14 VP.n29 VP.n28 161.3
R15 VP.n27 VP.n1 161.3
R16 VP.n26 VP.n25 161.3
R17 VP.n23 VP.n2 161.3
R18 VP.n22 VP.n21 161.3
R19 VP.n20 VP.n3 161.3
R20 VP.n19 VP.n18 161.3
R21 VP.n22 VP.n3 56.5193
R22 VP.n29 VP.n1 56.5193
R23 VP.n12 VP.n5 56.5193
R24 VP.n7 VP.n6 53.9242
R25 VP.n16 VP.n15 50.171
R26 VP.n18 VP.n3 24.4675
R27 VP.n23 VP.n22 24.4675
R28 VP.n25 VP.n1 24.4675
R29 VP.n30 VP.n29 24.4675
R30 VP.n13 VP.n12 24.4675
R31 VP.n8 VP.n5 24.4675
R32 VP.n9 VP.n6 17.9991
R33 VP.n24 VP.n23 12.234
R34 VP.n25 VP.n24 12.234
R35 VP.n8 VP.n7 12.234
R36 VP.n18 VP.n17 7.82994
R37 VP.n31 VP.n30 7.82994
R38 VP.n14 VP.n13 7.82994
R39 VP.n10 VP.n9 0.189894
R40 VP.n11 VP.n10 0.189894
R41 VP.n11 VP.n4 0.189894
R42 VP.n15 VP.n4 0.189894
R43 VP.n19 VP.n16 0.189894
R44 VP.n20 VP.n19 0.189894
R45 VP.n21 VP.n20 0.189894
R46 VP.n21 VP.n2 0.189894
R47 VP.n26 VP.n2 0.189894
R48 VP.n27 VP.n26 0.189894
R49 VP.n28 VP.n27 0.189894
R50 VP.n28 VP.n0 0.189894
R51 VP.n32 VP.n0 0.189894
R52 VP VP.n32 0.0516364
R53 VDD1 VDD1.t5 63.8961
R54 VDD1.n1 VDD1.t4 63.7824
R55 VDD1.n1 VDD1.n0 61.9371
R56 VDD1.n3 VDD1.n2 61.5807
R57 VDD1.n3 VDD1.n1 47.1711
R58 VDD1.n2 VDD1.t3 1.0227
R59 VDD1.n2 VDD1.t0 1.0227
R60 VDD1.n0 VDD1.t1 1.0227
R61 VDD1.n0 VDD1.t2 1.0227
R62 VDD1 VDD1.n3 0.353948
R63 VTAIL.n7 VTAIL.t2 45.9243
R64 VTAIL.n10 VTAIL.t8 45.924
R65 VTAIL.n11 VTAIL.t0 45.924
R66 VTAIL.n2 VTAIL.t7 45.924
R67 VTAIL.n9 VTAIL.n8 44.9021
R68 VTAIL.n6 VTAIL.n5 44.9021
R69 VTAIL.n1 VTAIL.n0 44.902
R70 VTAIL.n4 VTAIL.n3 44.902
R71 VTAIL.n6 VTAIL.n4 32.3583
R72 VTAIL.n11 VTAIL.n10 30.7117
R73 VTAIL.n7 VTAIL.n6 1.64705
R74 VTAIL.n10 VTAIL.n9 1.64705
R75 VTAIL.n4 VTAIL.n2 1.64705
R76 VTAIL.n9 VTAIL.n7 1.2936
R77 VTAIL.n2 VTAIL.n1 1.2936
R78 VTAIL VTAIL.n11 1.17722
R79 VTAIL.n0 VTAIL.t3 1.0227
R80 VTAIL.n0 VTAIL.t5 1.0227
R81 VTAIL.n3 VTAIL.t6 1.0227
R82 VTAIL.n3 VTAIL.t9 1.0227
R83 VTAIL.n8 VTAIL.t10 1.0227
R84 VTAIL.n8 VTAIL.t11 1.0227
R85 VTAIL.n5 VTAIL.t4 1.0227
R86 VTAIL.n5 VTAIL.t1 1.0227
R87 VTAIL VTAIL.n1 0.470328
R88 B.n666 B.n665 585
R89 B.n668 B.n130 585
R90 B.n671 B.n670 585
R91 B.n672 B.n129 585
R92 B.n674 B.n673 585
R93 B.n676 B.n128 585
R94 B.n679 B.n678 585
R95 B.n680 B.n127 585
R96 B.n682 B.n681 585
R97 B.n684 B.n126 585
R98 B.n687 B.n686 585
R99 B.n688 B.n125 585
R100 B.n690 B.n689 585
R101 B.n692 B.n124 585
R102 B.n695 B.n694 585
R103 B.n696 B.n123 585
R104 B.n698 B.n697 585
R105 B.n700 B.n122 585
R106 B.n703 B.n702 585
R107 B.n704 B.n121 585
R108 B.n706 B.n705 585
R109 B.n708 B.n120 585
R110 B.n711 B.n710 585
R111 B.n712 B.n119 585
R112 B.n714 B.n713 585
R113 B.n716 B.n118 585
R114 B.n719 B.n718 585
R115 B.n720 B.n117 585
R116 B.n722 B.n721 585
R117 B.n724 B.n116 585
R118 B.n727 B.n726 585
R119 B.n728 B.n115 585
R120 B.n730 B.n729 585
R121 B.n732 B.n114 585
R122 B.n735 B.n734 585
R123 B.n736 B.n113 585
R124 B.n738 B.n737 585
R125 B.n740 B.n112 585
R126 B.n743 B.n742 585
R127 B.n744 B.n111 585
R128 B.n746 B.n745 585
R129 B.n748 B.n110 585
R130 B.n751 B.n750 585
R131 B.n752 B.n109 585
R132 B.n754 B.n753 585
R133 B.n756 B.n108 585
R134 B.n759 B.n758 585
R135 B.n760 B.n107 585
R136 B.n762 B.n761 585
R137 B.n764 B.n106 585
R138 B.n767 B.n766 585
R139 B.n768 B.n105 585
R140 B.n770 B.n769 585
R141 B.n772 B.n104 585
R142 B.n775 B.n774 585
R143 B.n776 B.n103 585
R144 B.n778 B.n777 585
R145 B.n780 B.n102 585
R146 B.n783 B.n782 585
R147 B.n784 B.n101 585
R148 B.n786 B.n785 585
R149 B.n788 B.n100 585
R150 B.n791 B.n790 585
R151 B.n793 B.n97 585
R152 B.n795 B.n794 585
R153 B.n797 B.n96 585
R154 B.n800 B.n799 585
R155 B.n801 B.n95 585
R156 B.n803 B.n802 585
R157 B.n805 B.n94 585
R158 B.n808 B.n807 585
R159 B.n809 B.n90 585
R160 B.n811 B.n810 585
R161 B.n813 B.n89 585
R162 B.n816 B.n815 585
R163 B.n817 B.n88 585
R164 B.n819 B.n818 585
R165 B.n821 B.n87 585
R166 B.n824 B.n823 585
R167 B.n825 B.n86 585
R168 B.n827 B.n826 585
R169 B.n829 B.n85 585
R170 B.n832 B.n831 585
R171 B.n833 B.n84 585
R172 B.n835 B.n834 585
R173 B.n837 B.n83 585
R174 B.n840 B.n839 585
R175 B.n841 B.n82 585
R176 B.n843 B.n842 585
R177 B.n845 B.n81 585
R178 B.n848 B.n847 585
R179 B.n849 B.n80 585
R180 B.n851 B.n850 585
R181 B.n853 B.n79 585
R182 B.n856 B.n855 585
R183 B.n857 B.n78 585
R184 B.n859 B.n858 585
R185 B.n861 B.n77 585
R186 B.n864 B.n863 585
R187 B.n865 B.n76 585
R188 B.n867 B.n866 585
R189 B.n869 B.n75 585
R190 B.n872 B.n871 585
R191 B.n873 B.n74 585
R192 B.n875 B.n874 585
R193 B.n877 B.n73 585
R194 B.n880 B.n879 585
R195 B.n881 B.n72 585
R196 B.n883 B.n882 585
R197 B.n885 B.n71 585
R198 B.n888 B.n887 585
R199 B.n889 B.n70 585
R200 B.n891 B.n890 585
R201 B.n893 B.n69 585
R202 B.n896 B.n895 585
R203 B.n897 B.n68 585
R204 B.n899 B.n898 585
R205 B.n901 B.n67 585
R206 B.n904 B.n903 585
R207 B.n905 B.n66 585
R208 B.n907 B.n906 585
R209 B.n909 B.n65 585
R210 B.n912 B.n911 585
R211 B.n913 B.n64 585
R212 B.n915 B.n914 585
R213 B.n917 B.n63 585
R214 B.n920 B.n919 585
R215 B.n921 B.n62 585
R216 B.n923 B.n922 585
R217 B.n925 B.n61 585
R218 B.n928 B.n927 585
R219 B.n929 B.n60 585
R220 B.n931 B.n930 585
R221 B.n933 B.n59 585
R222 B.n936 B.n935 585
R223 B.n937 B.n58 585
R224 B.n664 B.n56 585
R225 B.n940 B.n56 585
R226 B.n663 B.n55 585
R227 B.n941 B.n55 585
R228 B.n662 B.n54 585
R229 B.n942 B.n54 585
R230 B.n661 B.n660 585
R231 B.n660 B.n50 585
R232 B.n659 B.n49 585
R233 B.n948 B.n49 585
R234 B.n658 B.n48 585
R235 B.n949 B.n48 585
R236 B.n657 B.n47 585
R237 B.n950 B.n47 585
R238 B.n656 B.n655 585
R239 B.n655 B.n43 585
R240 B.n654 B.n42 585
R241 B.n956 B.n42 585
R242 B.n653 B.n41 585
R243 B.n957 B.n41 585
R244 B.n652 B.n40 585
R245 B.n958 B.n40 585
R246 B.n651 B.n650 585
R247 B.n650 B.n36 585
R248 B.n649 B.n35 585
R249 B.n964 B.n35 585
R250 B.n648 B.n34 585
R251 B.n965 B.n34 585
R252 B.n647 B.n33 585
R253 B.n966 B.n33 585
R254 B.n646 B.n645 585
R255 B.n645 B.n29 585
R256 B.n644 B.n28 585
R257 B.n972 B.n28 585
R258 B.n643 B.n27 585
R259 B.n973 B.n27 585
R260 B.n642 B.n26 585
R261 B.n974 B.n26 585
R262 B.n641 B.n640 585
R263 B.n640 B.n22 585
R264 B.n639 B.n21 585
R265 B.n980 B.n21 585
R266 B.n638 B.n20 585
R267 B.n981 B.n20 585
R268 B.n637 B.n19 585
R269 B.n982 B.n19 585
R270 B.n636 B.n635 585
R271 B.n635 B.n15 585
R272 B.n634 B.n14 585
R273 B.n988 B.n14 585
R274 B.n633 B.n13 585
R275 B.n989 B.n13 585
R276 B.n632 B.n12 585
R277 B.n990 B.n12 585
R278 B.n631 B.n630 585
R279 B.n630 B.n629 585
R280 B.n628 B.n627 585
R281 B.n628 B.n8 585
R282 B.n626 B.n7 585
R283 B.n997 B.n7 585
R284 B.n625 B.n6 585
R285 B.n998 B.n6 585
R286 B.n624 B.n5 585
R287 B.n999 B.n5 585
R288 B.n623 B.n622 585
R289 B.n622 B.n4 585
R290 B.n621 B.n131 585
R291 B.n621 B.n620 585
R292 B.n611 B.n132 585
R293 B.n133 B.n132 585
R294 B.n613 B.n612 585
R295 B.n614 B.n613 585
R296 B.n610 B.n138 585
R297 B.n138 B.n137 585
R298 B.n609 B.n608 585
R299 B.n608 B.n607 585
R300 B.n140 B.n139 585
R301 B.n141 B.n140 585
R302 B.n600 B.n599 585
R303 B.n601 B.n600 585
R304 B.n598 B.n146 585
R305 B.n146 B.n145 585
R306 B.n597 B.n596 585
R307 B.n596 B.n595 585
R308 B.n148 B.n147 585
R309 B.n149 B.n148 585
R310 B.n588 B.n587 585
R311 B.n589 B.n588 585
R312 B.n586 B.n154 585
R313 B.n154 B.n153 585
R314 B.n585 B.n584 585
R315 B.n584 B.n583 585
R316 B.n156 B.n155 585
R317 B.n157 B.n156 585
R318 B.n576 B.n575 585
R319 B.n577 B.n576 585
R320 B.n574 B.n162 585
R321 B.n162 B.n161 585
R322 B.n573 B.n572 585
R323 B.n572 B.n571 585
R324 B.n164 B.n163 585
R325 B.n165 B.n164 585
R326 B.n564 B.n563 585
R327 B.n565 B.n564 585
R328 B.n562 B.n170 585
R329 B.n170 B.n169 585
R330 B.n561 B.n560 585
R331 B.n560 B.n559 585
R332 B.n172 B.n171 585
R333 B.n173 B.n172 585
R334 B.n552 B.n551 585
R335 B.n553 B.n552 585
R336 B.n550 B.n178 585
R337 B.n178 B.n177 585
R338 B.n549 B.n548 585
R339 B.n548 B.n547 585
R340 B.n180 B.n179 585
R341 B.n181 B.n180 585
R342 B.n540 B.n539 585
R343 B.n541 B.n540 585
R344 B.n538 B.n186 585
R345 B.n186 B.n185 585
R346 B.n537 B.n536 585
R347 B.n536 B.n535 585
R348 B.n532 B.n190 585
R349 B.n531 B.n530 585
R350 B.n528 B.n191 585
R351 B.n528 B.n189 585
R352 B.n527 B.n526 585
R353 B.n525 B.n524 585
R354 B.n523 B.n193 585
R355 B.n521 B.n520 585
R356 B.n519 B.n194 585
R357 B.n518 B.n517 585
R358 B.n515 B.n195 585
R359 B.n513 B.n512 585
R360 B.n511 B.n196 585
R361 B.n510 B.n509 585
R362 B.n507 B.n197 585
R363 B.n505 B.n504 585
R364 B.n503 B.n198 585
R365 B.n502 B.n501 585
R366 B.n499 B.n199 585
R367 B.n497 B.n496 585
R368 B.n495 B.n200 585
R369 B.n494 B.n493 585
R370 B.n491 B.n201 585
R371 B.n489 B.n488 585
R372 B.n487 B.n202 585
R373 B.n486 B.n485 585
R374 B.n483 B.n203 585
R375 B.n481 B.n480 585
R376 B.n479 B.n204 585
R377 B.n478 B.n477 585
R378 B.n475 B.n205 585
R379 B.n473 B.n472 585
R380 B.n471 B.n206 585
R381 B.n470 B.n469 585
R382 B.n467 B.n207 585
R383 B.n465 B.n464 585
R384 B.n463 B.n208 585
R385 B.n462 B.n461 585
R386 B.n459 B.n209 585
R387 B.n457 B.n456 585
R388 B.n455 B.n210 585
R389 B.n454 B.n453 585
R390 B.n451 B.n211 585
R391 B.n449 B.n448 585
R392 B.n447 B.n212 585
R393 B.n446 B.n445 585
R394 B.n443 B.n213 585
R395 B.n441 B.n440 585
R396 B.n439 B.n214 585
R397 B.n438 B.n437 585
R398 B.n435 B.n215 585
R399 B.n433 B.n432 585
R400 B.n431 B.n216 585
R401 B.n430 B.n429 585
R402 B.n427 B.n217 585
R403 B.n425 B.n424 585
R404 B.n423 B.n218 585
R405 B.n422 B.n421 585
R406 B.n419 B.n219 585
R407 B.n417 B.n416 585
R408 B.n415 B.n220 585
R409 B.n414 B.n413 585
R410 B.n411 B.n221 585
R411 B.n409 B.n408 585
R412 B.n406 B.n222 585
R413 B.n405 B.n404 585
R414 B.n402 B.n225 585
R415 B.n400 B.n399 585
R416 B.n398 B.n226 585
R417 B.n397 B.n396 585
R418 B.n394 B.n227 585
R419 B.n392 B.n391 585
R420 B.n390 B.n228 585
R421 B.n389 B.n388 585
R422 B.n386 B.n385 585
R423 B.n384 B.n383 585
R424 B.n382 B.n233 585
R425 B.n380 B.n379 585
R426 B.n378 B.n234 585
R427 B.n377 B.n376 585
R428 B.n374 B.n235 585
R429 B.n372 B.n371 585
R430 B.n370 B.n236 585
R431 B.n369 B.n368 585
R432 B.n366 B.n237 585
R433 B.n364 B.n363 585
R434 B.n362 B.n238 585
R435 B.n361 B.n360 585
R436 B.n358 B.n239 585
R437 B.n356 B.n355 585
R438 B.n354 B.n240 585
R439 B.n353 B.n352 585
R440 B.n350 B.n241 585
R441 B.n348 B.n347 585
R442 B.n346 B.n242 585
R443 B.n345 B.n344 585
R444 B.n342 B.n243 585
R445 B.n340 B.n339 585
R446 B.n338 B.n244 585
R447 B.n337 B.n336 585
R448 B.n334 B.n245 585
R449 B.n332 B.n331 585
R450 B.n330 B.n246 585
R451 B.n329 B.n328 585
R452 B.n326 B.n247 585
R453 B.n324 B.n323 585
R454 B.n322 B.n248 585
R455 B.n321 B.n320 585
R456 B.n318 B.n249 585
R457 B.n316 B.n315 585
R458 B.n314 B.n250 585
R459 B.n313 B.n312 585
R460 B.n310 B.n251 585
R461 B.n308 B.n307 585
R462 B.n306 B.n252 585
R463 B.n305 B.n304 585
R464 B.n302 B.n253 585
R465 B.n300 B.n299 585
R466 B.n298 B.n254 585
R467 B.n297 B.n296 585
R468 B.n294 B.n255 585
R469 B.n292 B.n291 585
R470 B.n290 B.n256 585
R471 B.n289 B.n288 585
R472 B.n286 B.n257 585
R473 B.n284 B.n283 585
R474 B.n282 B.n258 585
R475 B.n281 B.n280 585
R476 B.n278 B.n259 585
R477 B.n276 B.n275 585
R478 B.n274 B.n260 585
R479 B.n273 B.n272 585
R480 B.n270 B.n261 585
R481 B.n268 B.n267 585
R482 B.n266 B.n262 585
R483 B.n265 B.n264 585
R484 B.n188 B.n187 585
R485 B.n189 B.n188 585
R486 B.n534 B.n533 585
R487 B.n535 B.n534 585
R488 B.n184 B.n183 585
R489 B.n185 B.n184 585
R490 B.n543 B.n542 585
R491 B.n542 B.n541 585
R492 B.n544 B.n182 585
R493 B.n182 B.n181 585
R494 B.n546 B.n545 585
R495 B.n547 B.n546 585
R496 B.n176 B.n175 585
R497 B.n177 B.n176 585
R498 B.n555 B.n554 585
R499 B.n554 B.n553 585
R500 B.n556 B.n174 585
R501 B.n174 B.n173 585
R502 B.n558 B.n557 585
R503 B.n559 B.n558 585
R504 B.n168 B.n167 585
R505 B.n169 B.n168 585
R506 B.n567 B.n566 585
R507 B.n566 B.n565 585
R508 B.n568 B.n166 585
R509 B.n166 B.n165 585
R510 B.n570 B.n569 585
R511 B.n571 B.n570 585
R512 B.n160 B.n159 585
R513 B.n161 B.n160 585
R514 B.n579 B.n578 585
R515 B.n578 B.n577 585
R516 B.n580 B.n158 585
R517 B.n158 B.n157 585
R518 B.n582 B.n581 585
R519 B.n583 B.n582 585
R520 B.n152 B.n151 585
R521 B.n153 B.n152 585
R522 B.n591 B.n590 585
R523 B.n590 B.n589 585
R524 B.n592 B.n150 585
R525 B.n150 B.n149 585
R526 B.n594 B.n593 585
R527 B.n595 B.n594 585
R528 B.n144 B.n143 585
R529 B.n145 B.n144 585
R530 B.n603 B.n602 585
R531 B.n602 B.n601 585
R532 B.n604 B.n142 585
R533 B.n142 B.n141 585
R534 B.n606 B.n605 585
R535 B.n607 B.n606 585
R536 B.n136 B.n135 585
R537 B.n137 B.n136 585
R538 B.n616 B.n615 585
R539 B.n615 B.n614 585
R540 B.n617 B.n134 585
R541 B.n134 B.n133 585
R542 B.n619 B.n618 585
R543 B.n620 B.n619 585
R544 B.n3 B.n0 585
R545 B.n4 B.n3 585
R546 B.n996 B.n1 585
R547 B.n997 B.n996 585
R548 B.n995 B.n994 585
R549 B.n995 B.n8 585
R550 B.n993 B.n9 585
R551 B.n629 B.n9 585
R552 B.n992 B.n991 585
R553 B.n991 B.n990 585
R554 B.n11 B.n10 585
R555 B.n989 B.n11 585
R556 B.n987 B.n986 585
R557 B.n988 B.n987 585
R558 B.n985 B.n16 585
R559 B.n16 B.n15 585
R560 B.n984 B.n983 585
R561 B.n983 B.n982 585
R562 B.n18 B.n17 585
R563 B.n981 B.n18 585
R564 B.n979 B.n978 585
R565 B.n980 B.n979 585
R566 B.n977 B.n23 585
R567 B.n23 B.n22 585
R568 B.n976 B.n975 585
R569 B.n975 B.n974 585
R570 B.n25 B.n24 585
R571 B.n973 B.n25 585
R572 B.n971 B.n970 585
R573 B.n972 B.n971 585
R574 B.n969 B.n30 585
R575 B.n30 B.n29 585
R576 B.n968 B.n967 585
R577 B.n967 B.n966 585
R578 B.n32 B.n31 585
R579 B.n965 B.n32 585
R580 B.n963 B.n962 585
R581 B.n964 B.n963 585
R582 B.n961 B.n37 585
R583 B.n37 B.n36 585
R584 B.n960 B.n959 585
R585 B.n959 B.n958 585
R586 B.n39 B.n38 585
R587 B.n957 B.n39 585
R588 B.n955 B.n954 585
R589 B.n956 B.n955 585
R590 B.n953 B.n44 585
R591 B.n44 B.n43 585
R592 B.n952 B.n951 585
R593 B.n951 B.n950 585
R594 B.n46 B.n45 585
R595 B.n949 B.n46 585
R596 B.n947 B.n946 585
R597 B.n948 B.n947 585
R598 B.n945 B.n51 585
R599 B.n51 B.n50 585
R600 B.n944 B.n943 585
R601 B.n943 B.n942 585
R602 B.n53 B.n52 585
R603 B.n941 B.n53 585
R604 B.n939 B.n938 585
R605 B.n940 B.n939 585
R606 B.n1000 B.n999 585
R607 B.n998 B.n2 585
R608 B.n939 B.n58 526.135
R609 B.n666 B.n56 526.135
R610 B.n536 B.n188 526.135
R611 B.n534 B.n190 526.135
R612 B.n91 B.t6 501.18
R613 B.n98 B.t17 501.18
R614 B.n229 B.t14 501.18
R615 B.n223 B.t10 501.18
R616 B.n667 B.n57 256.663
R617 B.n669 B.n57 256.663
R618 B.n675 B.n57 256.663
R619 B.n677 B.n57 256.663
R620 B.n683 B.n57 256.663
R621 B.n685 B.n57 256.663
R622 B.n691 B.n57 256.663
R623 B.n693 B.n57 256.663
R624 B.n699 B.n57 256.663
R625 B.n701 B.n57 256.663
R626 B.n707 B.n57 256.663
R627 B.n709 B.n57 256.663
R628 B.n715 B.n57 256.663
R629 B.n717 B.n57 256.663
R630 B.n723 B.n57 256.663
R631 B.n725 B.n57 256.663
R632 B.n731 B.n57 256.663
R633 B.n733 B.n57 256.663
R634 B.n739 B.n57 256.663
R635 B.n741 B.n57 256.663
R636 B.n747 B.n57 256.663
R637 B.n749 B.n57 256.663
R638 B.n755 B.n57 256.663
R639 B.n757 B.n57 256.663
R640 B.n763 B.n57 256.663
R641 B.n765 B.n57 256.663
R642 B.n771 B.n57 256.663
R643 B.n773 B.n57 256.663
R644 B.n779 B.n57 256.663
R645 B.n781 B.n57 256.663
R646 B.n787 B.n57 256.663
R647 B.n789 B.n57 256.663
R648 B.n796 B.n57 256.663
R649 B.n798 B.n57 256.663
R650 B.n804 B.n57 256.663
R651 B.n806 B.n57 256.663
R652 B.n812 B.n57 256.663
R653 B.n814 B.n57 256.663
R654 B.n820 B.n57 256.663
R655 B.n822 B.n57 256.663
R656 B.n828 B.n57 256.663
R657 B.n830 B.n57 256.663
R658 B.n836 B.n57 256.663
R659 B.n838 B.n57 256.663
R660 B.n844 B.n57 256.663
R661 B.n846 B.n57 256.663
R662 B.n852 B.n57 256.663
R663 B.n854 B.n57 256.663
R664 B.n860 B.n57 256.663
R665 B.n862 B.n57 256.663
R666 B.n868 B.n57 256.663
R667 B.n870 B.n57 256.663
R668 B.n876 B.n57 256.663
R669 B.n878 B.n57 256.663
R670 B.n884 B.n57 256.663
R671 B.n886 B.n57 256.663
R672 B.n892 B.n57 256.663
R673 B.n894 B.n57 256.663
R674 B.n900 B.n57 256.663
R675 B.n902 B.n57 256.663
R676 B.n908 B.n57 256.663
R677 B.n910 B.n57 256.663
R678 B.n916 B.n57 256.663
R679 B.n918 B.n57 256.663
R680 B.n924 B.n57 256.663
R681 B.n926 B.n57 256.663
R682 B.n932 B.n57 256.663
R683 B.n934 B.n57 256.663
R684 B.n529 B.n189 256.663
R685 B.n192 B.n189 256.663
R686 B.n522 B.n189 256.663
R687 B.n516 B.n189 256.663
R688 B.n514 B.n189 256.663
R689 B.n508 B.n189 256.663
R690 B.n506 B.n189 256.663
R691 B.n500 B.n189 256.663
R692 B.n498 B.n189 256.663
R693 B.n492 B.n189 256.663
R694 B.n490 B.n189 256.663
R695 B.n484 B.n189 256.663
R696 B.n482 B.n189 256.663
R697 B.n476 B.n189 256.663
R698 B.n474 B.n189 256.663
R699 B.n468 B.n189 256.663
R700 B.n466 B.n189 256.663
R701 B.n460 B.n189 256.663
R702 B.n458 B.n189 256.663
R703 B.n452 B.n189 256.663
R704 B.n450 B.n189 256.663
R705 B.n444 B.n189 256.663
R706 B.n442 B.n189 256.663
R707 B.n436 B.n189 256.663
R708 B.n434 B.n189 256.663
R709 B.n428 B.n189 256.663
R710 B.n426 B.n189 256.663
R711 B.n420 B.n189 256.663
R712 B.n418 B.n189 256.663
R713 B.n412 B.n189 256.663
R714 B.n410 B.n189 256.663
R715 B.n403 B.n189 256.663
R716 B.n401 B.n189 256.663
R717 B.n395 B.n189 256.663
R718 B.n393 B.n189 256.663
R719 B.n387 B.n189 256.663
R720 B.n232 B.n189 256.663
R721 B.n381 B.n189 256.663
R722 B.n375 B.n189 256.663
R723 B.n373 B.n189 256.663
R724 B.n367 B.n189 256.663
R725 B.n365 B.n189 256.663
R726 B.n359 B.n189 256.663
R727 B.n357 B.n189 256.663
R728 B.n351 B.n189 256.663
R729 B.n349 B.n189 256.663
R730 B.n343 B.n189 256.663
R731 B.n341 B.n189 256.663
R732 B.n335 B.n189 256.663
R733 B.n333 B.n189 256.663
R734 B.n327 B.n189 256.663
R735 B.n325 B.n189 256.663
R736 B.n319 B.n189 256.663
R737 B.n317 B.n189 256.663
R738 B.n311 B.n189 256.663
R739 B.n309 B.n189 256.663
R740 B.n303 B.n189 256.663
R741 B.n301 B.n189 256.663
R742 B.n295 B.n189 256.663
R743 B.n293 B.n189 256.663
R744 B.n287 B.n189 256.663
R745 B.n285 B.n189 256.663
R746 B.n279 B.n189 256.663
R747 B.n277 B.n189 256.663
R748 B.n271 B.n189 256.663
R749 B.n269 B.n189 256.663
R750 B.n263 B.n189 256.663
R751 B.n1002 B.n1001 256.663
R752 B.n935 B.n933 163.367
R753 B.n931 B.n60 163.367
R754 B.n927 B.n925 163.367
R755 B.n923 B.n62 163.367
R756 B.n919 B.n917 163.367
R757 B.n915 B.n64 163.367
R758 B.n911 B.n909 163.367
R759 B.n907 B.n66 163.367
R760 B.n903 B.n901 163.367
R761 B.n899 B.n68 163.367
R762 B.n895 B.n893 163.367
R763 B.n891 B.n70 163.367
R764 B.n887 B.n885 163.367
R765 B.n883 B.n72 163.367
R766 B.n879 B.n877 163.367
R767 B.n875 B.n74 163.367
R768 B.n871 B.n869 163.367
R769 B.n867 B.n76 163.367
R770 B.n863 B.n861 163.367
R771 B.n859 B.n78 163.367
R772 B.n855 B.n853 163.367
R773 B.n851 B.n80 163.367
R774 B.n847 B.n845 163.367
R775 B.n843 B.n82 163.367
R776 B.n839 B.n837 163.367
R777 B.n835 B.n84 163.367
R778 B.n831 B.n829 163.367
R779 B.n827 B.n86 163.367
R780 B.n823 B.n821 163.367
R781 B.n819 B.n88 163.367
R782 B.n815 B.n813 163.367
R783 B.n811 B.n90 163.367
R784 B.n807 B.n805 163.367
R785 B.n803 B.n95 163.367
R786 B.n799 B.n797 163.367
R787 B.n795 B.n97 163.367
R788 B.n790 B.n788 163.367
R789 B.n786 B.n101 163.367
R790 B.n782 B.n780 163.367
R791 B.n778 B.n103 163.367
R792 B.n774 B.n772 163.367
R793 B.n770 B.n105 163.367
R794 B.n766 B.n764 163.367
R795 B.n762 B.n107 163.367
R796 B.n758 B.n756 163.367
R797 B.n754 B.n109 163.367
R798 B.n750 B.n748 163.367
R799 B.n746 B.n111 163.367
R800 B.n742 B.n740 163.367
R801 B.n738 B.n113 163.367
R802 B.n734 B.n732 163.367
R803 B.n730 B.n115 163.367
R804 B.n726 B.n724 163.367
R805 B.n722 B.n117 163.367
R806 B.n718 B.n716 163.367
R807 B.n714 B.n119 163.367
R808 B.n710 B.n708 163.367
R809 B.n706 B.n121 163.367
R810 B.n702 B.n700 163.367
R811 B.n698 B.n123 163.367
R812 B.n694 B.n692 163.367
R813 B.n690 B.n125 163.367
R814 B.n686 B.n684 163.367
R815 B.n682 B.n127 163.367
R816 B.n678 B.n676 163.367
R817 B.n674 B.n129 163.367
R818 B.n670 B.n668 163.367
R819 B.n536 B.n186 163.367
R820 B.n540 B.n186 163.367
R821 B.n540 B.n180 163.367
R822 B.n548 B.n180 163.367
R823 B.n548 B.n178 163.367
R824 B.n552 B.n178 163.367
R825 B.n552 B.n172 163.367
R826 B.n560 B.n172 163.367
R827 B.n560 B.n170 163.367
R828 B.n564 B.n170 163.367
R829 B.n564 B.n164 163.367
R830 B.n572 B.n164 163.367
R831 B.n572 B.n162 163.367
R832 B.n576 B.n162 163.367
R833 B.n576 B.n156 163.367
R834 B.n584 B.n156 163.367
R835 B.n584 B.n154 163.367
R836 B.n588 B.n154 163.367
R837 B.n588 B.n148 163.367
R838 B.n596 B.n148 163.367
R839 B.n596 B.n146 163.367
R840 B.n600 B.n146 163.367
R841 B.n600 B.n140 163.367
R842 B.n608 B.n140 163.367
R843 B.n608 B.n138 163.367
R844 B.n613 B.n138 163.367
R845 B.n613 B.n132 163.367
R846 B.n621 B.n132 163.367
R847 B.n622 B.n621 163.367
R848 B.n622 B.n5 163.367
R849 B.n6 B.n5 163.367
R850 B.n7 B.n6 163.367
R851 B.n628 B.n7 163.367
R852 B.n630 B.n628 163.367
R853 B.n630 B.n12 163.367
R854 B.n13 B.n12 163.367
R855 B.n14 B.n13 163.367
R856 B.n635 B.n14 163.367
R857 B.n635 B.n19 163.367
R858 B.n20 B.n19 163.367
R859 B.n21 B.n20 163.367
R860 B.n640 B.n21 163.367
R861 B.n640 B.n26 163.367
R862 B.n27 B.n26 163.367
R863 B.n28 B.n27 163.367
R864 B.n645 B.n28 163.367
R865 B.n645 B.n33 163.367
R866 B.n34 B.n33 163.367
R867 B.n35 B.n34 163.367
R868 B.n650 B.n35 163.367
R869 B.n650 B.n40 163.367
R870 B.n41 B.n40 163.367
R871 B.n42 B.n41 163.367
R872 B.n655 B.n42 163.367
R873 B.n655 B.n47 163.367
R874 B.n48 B.n47 163.367
R875 B.n49 B.n48 163.367
R876 B.n660 B.n49 163.367
R877 B.n660 B.n54 163.367
R878 B.n55 B.n54 163.367
R879 B.n56 B.n55 163.367
R880 B.n530 B.n528 163.367
R881 B.n528 B.n527 163.367
R882 B.n524 B.n523 163.367
R883 B.n521 B.n194 163.367
R884 B.n517 B.n515 163.367
R885 B.n513 B.n196 163.367
R886 B.n509 B.n507 163.367
R887 B.n505 B.n198 163.367
R888 B.n501 B.n499 163.367
R889 B.n497 B.n200 163.367
R890 B.n493 B.n491 163.367
R891 B.n489 B.n202 163.367
R892 B.n485 B.n483 163.367
R893 B.n481 B.n204 163.367
R894 B.n477 B.n475 163.367
R895 B.n473 B.n206 163.367
R896 B.n469 B.n467 163.367
R897 B.n465 B.n208 163.367
R898 B.n461 B.n459 163.367
R899 B.n457 B.n210 163.367
R900 B.n453 B.n451 163.367
R901 B.n449 B.n212 163.367
R902 B.n445 B.n443 163.367
R903 B.n441 B.n214 163.367
R904 B.n437 B.n435 163.367
R905 B.n433 B.n216 163.367
R906 B.n429 B.n427 163.367
R907 B.n425 B.n218 163.367
R908 B.n421 B.n419 163.367
R909 B.n417 B.n220 163.367
R910 B.n413 B.n411 163.367
R911 B.n409 B.n222 163.367
R912 B.n404 B.n402 163.367
R913 B.n400 B.n226 163.367
R914 B.n396 B.n394 163.367
R915 B.n392 B.n228 163.367
R916 B.n388 B.n386 163.367
R917 B.n383 B.n382 163.367
R918 B.n380 B.n234 163.367
R919 B.n376 B.n374 163.367
R920 B.n372 B.n236 163.367
R921 B.n368 B.n366 163.367
R922 B.n364 B.n238 163.367
R923 B.n360 B.n358 163.367
R924 B.n356 B.n240 163.367
R925 B.n352 B.n350 163.367
R926 B.n348 B.n242 163.367
R927 B.n344 B.n342 163.367
R928 B.n340 B.n244 163.367
R929 B.n336 B.n334 163.367
R930 B.n332 B.n246 163.367
R931 B.n328 B.n326 163.367
R932 B.n324 B.n248 163.367
R933 B.n320 B.n318 163.367
R934 B.n316 B.n250 163.367
R935 B.n312 B.n310 163.367
R936 B.n308 B.n252 163.367
R937 B.n304 B.n302 163.367
R938 B.n300 B.n254 163.367
R939 B.n296 B.n294 163.367
R940 B.n292 B.n256 163.367
R941 B.n288 B.n286 163.367
R942 B.n284 B.n258 163.367
R943 B.n280 B.n278 163.367
R944 B.n276 B.n260 163.367
R945 B.n272 B.n270 163.367
R946 B.n268 B.n262 163.367
R947 B.n264 B.n188 163.367
R948 B.n534 B.n184 163.367
R949 B.n542 B.n184 163.367
R950 B.n542 B.n182 163.367
R951 B.n546 B.n182 163.367
R952 B.n546 B.n176 163.367
R953 B.n554 B.n176 163.367
R954 B.n554 B.n174 163.367
R955 B.n558 B.n174 163.367
R956 B.n558 B.n168 163.367
R957 B.n566 B.n168 163.367
R958 B.n566 B.n166 163.367
R959 B.n570 B.n166 163.367
R960 B.n570 B.n160 163.367
R961 B.n578 B.n160 163.367
R962 B.n578 B.n158 163.367
R963 B.n582 B.n158 163.367
R964 B.n582 B.n152 163.367
R965 B.n590 B.n152 163.367
R966 B.n590 B.n150 163.367
R967 B.n594 B.n150 163.367
R968 B.n594 B.n144 163.367
R969 B.n602 B.n144 163.367
R970 B.n602 B.n142 163.367
R971 B.n606 B.n142 163.367
R972 B.n606 B.n136 163.367
R973 B.n615 B.n136 163.367
R974 B.n615 B.n134 163.367
R975 B.n619 B.n134 163.367
R976 B.n619 B.n3 163.367
R977 B.n1000 B.n3 163.367
R978 B.n996 B.n2 163.367
R979 B.n996 B.n995 163.367
R980 B.n995 B.n9 163.367
R981 B.n991 B.n9 163.367
R982 B.n991 B.n11 163.367
R983 B.n987 B.n11 163.367
R984 B.n987 B.n16 163.367
R985 B.n983 B.n16 163.367
R986 B.n983 B.n18 163.367
R987 B.n979 B.n18 163.367
R988 B.n979 B.n23 163.367
R989 B.n975 B.n23 163.367
R990 B.n975 B.n25 163.367
R991 B.n971 B.n25 163.367
R992 B.n971 B.n30 163.367
R993 B.n967 B.n30 163.367
R994 B.n967 B.n32 163.367
R995 B.n963 B.n32 163.367
R996 B.n963 B.n37 163.367
R997 B.n959 B.n37 163.367
R998 B.n959 B.n39 163.367
R999 B.n955 B.n39 163.367
R1000 B.n955 B.n44 163.367
R1001 B.n951 B.n44 163.367
R1002 B.n951 B.n46 163.367
R1003 B.n947 B.n46 163.367
R1004 B.n947 B.n51 163.367
R1005 B.n943 B.n51 163.367
R1006 B.n943 B.n53 163.367
R1007 B.n939 B.n53 163.367
R1008 B.n98 B.t18 110.615
R1009 B.n229 B.t16 110.615
R1010 B.n91 B.t8 110.59
R1011 B.n223 B.t13 110.59
R1012 B.n99 B.t19 73.5726
R1013 B.n230 B.t15 73.5726
R1014 B.n92 B.t9 73.5469
R1015 B.n224 B.t12 73.5469
R1016 B.n934 B.n58 71.676
R1017 B.n933 B.n932 71.676
R1018 B.n926 B.n60 71.676
R1019 B.n925 B.n924 71.676
R1020 B.n918 B.n62 71.676
R1021 B.n917 B.n916 71.676
R1022 B.n910 B.n64 71.676
R1023 B.n909 B.n908 71.676
R1024 B.n902 B.n66 71.676
R1025 B.n901 B.n900 71.676
R1026 B.n894 B.n68 71.676
R1027 B.n893 B.n892 71.676
R1028 B.n886 B.n70 71.676
R1029 B.n885 B.n884 71.676
R1030 B.n878 B.n72 71.676
R1031 B.n877 B.n876 71.676
R1032 B.n870 B.n74 71.676
R1033 B.n869 B.n868 71.676
R1034 B.n862 B.n76 71.676
R1035 B.n861 B.n860 71.676
R1036 B.n854 B.n78 71.676
R1037 B.n853 B.n852 71.676
R1038 B.n846 B.n80 71.676
R1039 B.n845 B.n844 71.676
R1040 B.n838 B.n82 71.676
R1041 B.n837 B.n836 71.676
R1042 B.n830 B.n84 71.676
R1043 B.n829 B.n828 71.676
R1044 B.n822 B.n86 71.676
R1045 B.n821 B.n820 71.676
R1046 B.n814 B.n88 71.676
R1047 B.n813 B.n812 71.676
R1048 B.n806 B.n90 71.676
R1049 B.n805 B.n804 71.676
R1050 B.n798 B.n95 71.676
R1051 B.n797 B.n796 71.676
R1052 B.n789 B.n97 71.676
R1053 B.n788 B.n787 71.676
R1054 B.n781 B.n101 71.676
R1055 B.n780 B.n779 71.676
R1056 B.n773 B.n103 71.676
R1057 B.n772 B.n771 71.676
R1058 B.n765 B.n105 71.676
R1059 B.n764 B.n763 71.676
R1060 B.n757 B.n107 71.676
R1061 B.n756 B.n755 71.676
R1062 B.n749 B.n109 71.676
R1063 B.n748 B.n747 71.676
R1064 B.n741 B.n111 71.676
R1065 B.n740 B.n739 71.676
R1066 B.n733 B.n113 71.676
R1067 B.n732 B.n731 71.676
R1068 B.n725 B.n115 71.676
R1069 B.n724 B.n723 71.676
R1070 B.n717 B.n117 71.676
R1071 B.n716 B.n715 71.676
R1072 B.n709 B.n119 71.676
R1073 B.n708 B.n707 71.676
R1074 B.n701 B.n121 71.676
R1075 B.n700 B.n699 71.676
R1076 B.n693 B.n123 71.676
R1077 B.n692 B.n691 71.676
R1078 B.n685 B.n125 71.676
R1079 B.n684 B.n683 71.676
R1080 B.n677 B.n127 71.676
R1081 B.n676 B.n675 71.676
R1082 B.n669 B.n129 71.676
R1083 B.n668 B.n667 71.676
R1084 B.n667 B.n666 71.676
R1085 B.n670 B.n669 71.676
R1086 B.n675 B.n674 71.676
R1087 B.n678 B.n677 71.676
R1088 B.n683 B.n682 71.676
R1089 B.n686 B.n685 71.676
R1090 B.n691 B.n690 71.676
R1091 B.n694 B.n693 71.676
R1092 B.n699 B.n698 71.676
R1093 B.n702 B.n701 71.676
R1094 B.n707 B.n706 71.676
R1095 B.n710 B.n709 71.676
R1096 B.n715 B.n714 71.676
R1097 B.n718 B.n717 71.676
R1098 B.n723 B.n722 71.676
R1099 B.n726 B.n725 71.676
R1100 B.n731 B.n730 71.676
R1101 B.n734 B.n733 71.676
R1102 B.n739 B.n738 71.676
R1103 B.n742 B.n741 71.676
R1104 B.n747 B.n746 71.676
R1105 B.n750 B.n749 71.676
R1106 B.n755 B.n754 71.676
R1107 B.n758 B.n757 71.676
R1108 B.n763 B.n762 71.676
R1109 B.n766 B.n765 71.676
R1110 B.n771 B.n770 71.676
R1111 B.n774 B.n773 71.676
R1112 B.n779 B.n778 71.676
R1113 B.n782 B.n781 71.676
R1114 B.n787 B.n786 71.676
R1115 B.n790 B.n789 71.676
R1116 B.n796 B.n795 71.676
R1117 B.n799 B.n798 71.676
R1118 B.n804 B.n803 71.676
R1119 B.n807 B.n806 71.676
R1120 B.n812 B.n811 71.676
R1121 B.n815 B.n814 71.676
R1122 B.n820 B.n819 71.676
R1123 B.n823 B.n822 71.676
R1124 B.n828 B.n827 71.676
R1125 B.n831 B.n830 71.676
R1126 B.n836 B.n835 71.676
R1127 B.n839 B.n838 71.676
R1128 B.n844 B.n843 71.676
R1129 B.n847 B.n846 71.676
R1130 B.n852 B.n851 71.676
R1131 B.n855 B.n854 71.676
R1132 B.n860 B.n859 71.676
R1133 B.n863 B.n862 71.676
R1134 B.n868 B.n867 71.676
R1135 B.n871 B.n870 71.676
R1136 B.n876 B.n875 71.676
R1137 B.n879 B.n878 71.676
R1138 B.n884 B.n883 71.676
R1139 B.n887 B.n886 71.676
R1140 B.n892 B.n891 71.676
R1141 B.n895 B.n894 71.676
R1142 B.n900 B.n899 71.676
R1143 B.n903 B.n902 71.676
R1144 B.n908 B.n907 71.676
R1145 B.n911 B.n910 71.676
R1146 B.n916 B.n915 71.676
R1147 B.n919 B.n918 71.676
R1148 B.n924 B.n923 71.676
R1149 B.n927 B.n926 71.676
R1150 B.n932 B.n931 71.676
R1151 B.n935 B.n934 71.676
R1152 B.n529 B.n190 71.676
R1153 B.n527 B.n192 71.676
R1154 B.n523 B.n522 71.676
R1155 B.n516 B.n194 71.676
R1156 B.n515 B.n514 71.676
R1157 B.n508 B.n196 71.676
R1158 B.n507 B.n506 71.676
R1159 B.n500 B.n198 71.676
R1160 B.n499 B.n498 71.676
R1161 B.n492 B.n200 71.676
R1162 B.n491 B.n490 71.676
R1163 B.n484 B.n202 71.676
R1164 B.n483 B.n482 71.676
R1165 B.n476 B.n204 71.676
R1166 B.n475 B.n474 71.676
R1167 B.n468 B.n206 71.676
R1168 B.n467 B.n466 71.676
R1169 B.n460 B.n208 71.676
R1170 B.n459 B.n458 71.676
R1171 B.n452 B.n210 71.676
R1172 B.n451 B.n450 71.676
R1173 B.n444 B.n212 71.676
R1174 B.n443 B.n442 71.676
R1175 B.n436 B.n214 71.676
R1176 B.n435 B.n434 71.676
R1177 B.n428 B.n216 71.676
R1178 B.n427 B.n426 71.676
R1179 B.n420 B.n218 71.676
R1180 B.n419 B.n418 71.676
R1181 B.n412 B.n220 71.676
R1182 B.n411 B.n410 71.676
R1183 B.n403 B.n222 71.676
R1184 B.n402 B.n401 71.676
R1185 B.n395 B.n226 71.676
R1186 B.n394 B.n393 71.676
R1187 B.n387 B.n228 71.676
R1188 B.n386 B.n232 71.676
R1189 B.n382 B.n381 71.676
R1190 B.n375 B.n234 71.676
R1191 B.n374 B.n373 71.676
R1192 B.n367 B.n236 71.676
R1193 B.n366 B.n365 71.676
R1194 B.n359 B.n238 71.676
R1195 B.n358 B.n357 71.676
R1196 B.n351 B.n240 71.676
R1197 B.n350 B.n349 71.676
R1198 B.n343 B.n242 71.676
R1199 B.n342 B.n341 71.676
R1200 B.n335 B.n244 71.676
R1201 B.n334 B.n333 71.676
R1202 B.n327 B.n246 71.676
R1203 B.n326 B.n325 71.676
R1204 B.n319 B.n248 71.676
R1205 B.n318 B.n317 71.676
R1206 B.n311 B.n250 71.676
R1207 B.n310 B.n309 71.676
R1208 B.n303 B.n252 71.676
R1209 B.n302 B.n301 71.676
R1210 B.n295 B.n254 71.676
R1211 B.n294 B.n293 71.676
R1212 B.n287 B.n256 71.676
R1213 B.n286 B.n285 71.676
R1214 B.n279 B.n258 71.676
R1215 B.n278 B.n277 71.676
R1216 B.n271 B.n260 71.676
R1217 B.n270 B.n269 71.676
R1218 B.n263 B.n262 71.676
R1219 B.n530 B.n529 71.676
R1220 B.n524 B.n192 71.676
R1221 B.n522 B.n521 71.676
R1222 B.n517 B.n516 71.676
R1223 B.n514 B.n513 71.676
R1224 B.n509 B.n508 71.676
R1225 B.n506 B.n505 71.676
R1226 B.n501 B.n500 71.676
R1227 B.n498 B.n497 71.676
R1228 B.n493 B.n492 71.676
R1229 B.n490 B.n489 71.676
R1230 B.n485 B.n484 71.676
R1231 B.n482 B.n481 71.676
R1232 B.n477 B.n476 71.676
R1233 B.n474 B.n473 71.676
R1234 B.n469 B.n468 71.676
R1235 B.n466 B.n465 71.676
R1236 B.n461 B.n460 71.676
R1237 B.n458 B.n457 71.676
R1238 B.n453 B.n452 71.676
R1239 B.n450 B.n449 71.676
R1240 B.n445 B.n444 71.676
R1241 B.n442 B.n441 71.676
R1242 B.n437 B.n436 71.676
R1243 B.n434 B.n433 71.676
R1244 B.n429 B.n428 71.676
R1245 B.n426 B.n425 71.676
R1246 B.n421 B.n420 71.676
R1247 B.n418 B.n417 71.676
R1248 B.n413 B.n412 71.676
R1249 B.n410 B.n409 71.676
R1250 B.n404 B.n403 71.676
R1251 B.n401 B.n400 71.676
R1252 B.n396 B.n395 71.676
R1253 B.n393 B.n392 71.676
R1254 B.n388 B.n387 71.676
R1255 B.n383 B.n232 71.676
R1256 B.n381 B.n380 71.676
R1257 B.n376 B.n375 71.676
R1258 B.n373 B.n372 71.676
R1259 B.n368 B.n367 71.676
R1260 B.n365 B.n364 71.676
R1261 B.n360 B.n359 71.676
R1262 B.n357 B.n356 71.676
R1263 B.n352 B.n351 71.676
R1264 B.n349 B.n348 71.676
R1265 B.n344 B.n343 71.676
R1266 B.n341 B.n340 71.676
R1267 B.n336 B.n335 71.676
R1268 B.n333 B.n332 71.676
R1269 B.n328 B.n327 71.676
R1270 B.n325 B.n324 71.676
R1271 B.n320 B.n319 71.676
R1272 B.n317 B.n316 71.676
R1273 B.n312 B.n311 71.676
R1274 B.n309 B.n308 71.676
R1275 B.n304 B.n303 71.676
R1276 B.n301 B.n300 71.676
R1277 B.n296 B.n295 71.676
R1278 B.n293 B.n292 71.676
R1279 B.n288 B.n287 71.676
R1280 B.n285 B.n284 71.676
R1281 B.n280 B.n279 71.676
R1282 B.n277 B.n276 71.676
R1283 B.n272 B.n271 71.676
R1284 B.n269 B.n268 71.676
R1285 B.n264 B.n263 71.676
R1286 B.n1001 B.n1000 71.676
R1287 B.n1001 B.n2 71.676
R1288 B.n93 B.n92 59.5399
R1289 B.n792 B.n99 59.5399
R1290 B.n231 B.n230 59.5399
R1291 B.n407 B.n224 59.5399
R1292 B.n535 B.n189 57.5781
R1293 B.n940 B.n57 57.5781
R1294 B.n92 B.n91 37.0429
R1295 B.n99 B.n98 37.0429
R1296 B.n230 B.n229 37.0429
R1297 B.n224 B.n223 37.0429
R1298 B.n533 B.n532 34.1859
R1299 B.n537 B.n187 34.1859
R1300 B.n665 B.n664 34.1859
R1301 B.n938 B.n937 34.1859
R1302 B.n535 B.n185 30.3515
R1303 B.n541 B.n185 30.3515
R1304 B.n541 B.n181 30.3515
R1305 B.n547 B.n181 30.3515
R1306 B.n547 B.n177 30.3515
R1307 B.n553 B.n177 30.3515
R1308 B.n559 B.n173 30.3515
R1309 B.n559 B.n169 30.3515
R1310 B.n565 B.n169 30.3515
R1311 B.n565 B.n165 30.3515
R1312 B.n571 B.n165 30.3515
R1313 B.n571 B.n161 30.3515
R1314 B.n577 B.n161 30.3515
R1315 B.n583 B.n157 30.3515
R1316 B.n583 B.n153 30.3515
R1317 B.n589 B.n153 30.3515
R1318 B.n589 B.n149 30.3515
R1319 B.n595 B.n149 30.3515
R1320 B.n601 B.n145 30.3515
R1321 B.n601 B.n141 30.3515
R1322 B.n607 B.n141 30.3515
R1323 B.n607 B.n137 30.3515
R1324 B.n614 B.n137 30.3515
R1325 B.n620 B.n133 30.3515
R1326 B.n620 B.n4 30.3515
R1327 B.n999 B.n4 30.3515
R1328 B.n999 B.n998 30.3515
R1329 B.n998 B.n997 30.3515
R1330 B.n997 B.n8 30.3515
R1331 B.n629 B.n8 30.3515
R1332 B.n990 B.n989 30.3515
R1333 B.n989 B.n988 30.3515
R1334 B.n988 B.n15 30.3515
R1335 B.n982 B.n15 30.3515
R1336 B.n982 B.n981 30.3515
R1337 B.n980 B.n22 30.3515
R1338 B.n974 B.n22 30.3515
R1339 B.n974 B.n973 30.3515
R1340 B.n973 B.n972 30.3515
R1341 B.n972 B.n29 30.3515
R1342 B.n966 B.n965 30.3515
R1343 B.n965 B.n964 30.3515
R1344 B.n964 B.n36 30.3515
R1345 B.n958 B.n36 30.3515
R1346 B.n958 B.n957 30.3515
R1347 B.n957 B.n956 30.3515
R1348 B.n956 B.n43 30.3515
R1349 B.n950 B.n949 30.3515
R1350 B.n949 B.n948 30.3515
R1351 B.n948 B.n50 30.3515
R1352 B.n942 B.n50 30.3515
R1353 B.n942 B.n941 30.3515
R1354 B.n941 B.n940 30.3515
R1355 B.t11 B.n173 29.4588
R1356 B.t7 B.n43 29.4588
R1357 B.t2 B.n133 27.6735
R1358 B.n629 B.t3 27.6735
R1359 B.n577 B.t4 25.8881
R1360 B.n966 B.t0 25.8881
R1361 B B.n1002 18.0485
R1362 B.t1 B.n145 16.0687
R1363 B.n981 B.t5 16.0687
R1364 B.n595 B.t1 14.2833
R1365 B.t5 B.n980 14.2833
R1366 B.n533 B.n183 10.6151
R1367 B.n543 B.n183 10.6151
R1368 B.n544 B.n543 10.6151
R1369 B.n545 B.n544 10.6151
R1370 B.n545 B.n175 10.6151
R1371 B.n555 B.n175 10.6151
R1372 B.n556 B.n555 10.6151
R1373 B.n557 B.n556 10.6151
R1374 B.n557 B.n167 10.6151
R1375 B.n567 B.n167 10.6151
R1376 B.n568 B.n567 10.6151
R1377 B.n569 B.n568 10.6151
R1378 B.n569 B.n159 10.6151
R1379 B.n579 B.n159 10.6151
R1380 B.n580 B.n579 10.6151
R1381 B.n581 B.n580 10.6151
R1382 B.n581 B.n151 10.6151
R1383 B.n591 B.n151 10.6151
R1384 B.n592 B.n591 10.6151
R1385 B.n593 B.n592 10.6151
R1386 B.n593 B.n143 10.6151
R1387 B.n603 B.n143 10.6151
R1388 B.n604 B.n603 10.6151
R1389 B.n605 B.n604 10.6151
R1390 B.n605 B.n135 10.6151
R1391 B.n616 B.n135 10.6151
R1392 B.n617 B.n616 10.6151
R1393 B.n618 B.n617 10.6151
R1394 B.n618 B.n0 10.6151
R1395 B.n532 B.n531 10.6151
R1396 B.n531 B.n191 10.6151
R1397 B.n526 B.n191 10.6151
R1398 B.n526 B.n525 10.6151
R1399 B.n525 B.n193 10.6151
R1400 B.n520 B.n193 10.6151
R1401 B.n520 B.n519 10.6151
R1402 B.n519 B.n518 10.6151
R1403 B.n518 B.n195 10.6151
R1404 B.n512 B.n195 10.6151
R1405 B.n512 B.n511 10.6151
R1406 B.n511 B.n510 10.6151
R1407 B.n510 B.n197 10.6151
R1408 B.n504 B.n197 10.6151
R1409 B.n504 B.n503 10.6151
R1410 B.n503 B.n502 10.6151
R1411 B.n502 B.n199 10.6151
R1412 B.n496 B.n199 10.6151
R1413 B.n496 B.n495 10.6151
R1414 B.n495 B.n494 10.6151
R1415 B.n494 B.n201 10.6151
R1416 B.n488 B.n201 10.6151
R1417 B.n488 B.n487 10.6151
R1418 B.n487 B.n486 10.6151
R1419 B.n486 B.n203 10.6151
R1420 B.n480 B.n203 10.6151
R1421 B.n480 B.n479 10.6151
R1422 B.n479 B.n478 10.6151
R1423 B.n478 B.n205 10.6151
R1424 B.n472 B.n205 10.6151
R1425 B.n472 B.n471 10.6151
R1426 B.n471 B.n470 10.6151
R1427 B.n470 B.n207 10.6151
R1428 B.n464 B.n207 10.6151
R1429 B.n464 B.n463 10.6151
R1430 B.n463 B.n462 10.6151
R1431 B.n462 B.n209 10.6151
R1432 B.n456 B.n209 10.6151
R1433 B.n456 B.n455 10.6151
R1434 B.n455 B.n454 10.6151
R1435 B.n454 B.n211 10.6151
R1436 B.n448 B.n211 10.6151
R1437 B.n448 B.n447 10.6151
R1438 B.n447 B.n446 10.6151
R1439 B.n446 B.n213 10.6151
R1440 B.n440 B.n213 10.6151
R1441 B.n440 B.n439 10.6151
R1442 B.n439 B.n438 10.6151
R1443 B.n438 B.n215 10.6151
R1444 B.n432 B.n215 10.6151
R1445 B.n432 B.n431 10.6151
R1446 B.n431 B.n430 10.6151
R1447 B.n430 B.n217 10.6151
R1448 B.n424 B.n217 10.6151
R1449 B.n424 B.n423 10.6151
R1450 B.n423 B.n422 10.6151
R1451 B.n422 B.n219 10.6151
R1452 B.n416 B.n219 10.6151
R1453 B.n416 B.n415 10.6151
R1454 B.n415 B.n414 10.6151
R1455 B.n414 B.n221 10.6151
R1456 B.n408 B.n221 10.6151
R1457 B.n406 B.n405 10.6151
R1458 B.n405 B.n225 10.6151
R1459 B.n399 B.n225 10.6151
R1460 B.n399 B.n398 10.6151
R1461 B.n398 B.n397 10.6151
R1462 B.n397 B.n227 10.6151
R1463 B.n391 B.n227 10.6151
R1464 B.n391 B.n390 10.6151
R1465 B.n390 B.n389 10.6151
R1466 B.n385 B.n384 10.6151
R1467 B.n384 B.n233 10.6151
R1468 B.n379 B.n233 10.6151
R1469 B.n379 B.n378 10.6151
R1470 B.n378 B.n377 10.6151
R1471 B.n377 B.n235 10.6151
R1472 B.n371 B.n235 10.6151
R1473 B.n371 B.n370 10.6151
R1474 B.n370 B.n369 10.6151
R1475 B.n369 B.n237 10.6151
R1476 B.n363 B.n237 10.6151
R1477 B.n363 B.n362 10.6151
R1478 B.n362 B.n361 10.6151
R1479 B.n361 B.n239 10.6151
R1480 B.n355 B.n239 10.6151
R1481 B.n355 B.n354 10.6151
R1482 B.n354 B.n353 10.6151
R1483 B.n353 B.n241 10.6151
R1484 B.n347 B.n241 10.6151
R1485 B.n347 B.n346 10.6151
R1486 B.n346 B.n345 10.6151
R1487 B.n345 B.n243 10.6151
R1488 B.n339 B.n243 10.6151
R1489 B.n339 B.n338 10.6151
R1490 B.n338 B.n337 10.6151
R1491 B.n337 B.n245 10.6151
R1492 B.n331 B.n245 10.6151
R1493 B.n331 B.n330 10.6151
R1494 B.n330 B.n329 10.6151
R1495 B.n329 B.n247 10.6151
R1496 B.n323 B.n247 10.6151
R1497 B.n323 B.n322 10.6151
R1498 B.n322 B.n321 10.6151
R1499 B.n321 B.n249 10.6151
R1500 B.n315 B.n249 10.6151
R1501 B.n315 B.n314 10.6151
R1502 B.n314 B.n313 10.6151
R1503 B.n313 B.n251 10.6151
R1504 B.n307 B.n251 10.6151
R1505 B.n307 B.n306 10.6151
R1506 B.n306 B.n305 10.6151
R1507 B.n305 B.n253 10.6151
R1508 B.n299 B.n253 10.6151
R1509 B.n299 B.n298 10.6151
R1510 B.n298 B.n297 10.6151
R1511 B.n297 B.n255 10.6151
R1512 B.n291 B.n255 10.6151
R1513 B.n291 B.n290 10.6151
R1514 B.n290 B.n289 10.6151
R1515 B.n289 B.n257 10.6151
R1516 B.n283 B.n257 10.6151
R1517 B.n283 B.n282 10.6151
R1518 B.n282 B.n281 10.6151
R1519 B.n281 B.n259 10.6151
R1520 B.n275 B.n259 10.6151
R1521 B.n275 B.n274 10.6151
R1522 B.n274 B.n273 10.6151
R1523 B.n273 B.n261 10.6151
R1524 B.n267 B.n261 10.6151
R1525 B.n267 B.n266 10.6151
R1526 B.n266 B.n265 10.6151
R1527 B.n265 B.n187 10.6151
R1528 B.n538 B.n537 10.6151
R1529 B.n539 B.n538 10.6151
R1530 B.n539 B.n179 10.6151
R1531 B.n549 B.n179 10.6151
R1532 B.n550 B.n549 10.6151
R1533 B.n551 B.n550 10.6151
R1534 B.n551 B.n171 10.6151
R1535 B.n561 B.n171 10.6151
R1536 B.n562 B.n561 10.6151
R1537 B.n563 B.n562 10.6151
R1538 B.n563 B.n163 10.6151
R1539 B.n573 B.n163 10.6151
R1540 B.n574 B.n573 10.6151
R1541 B.n575 B.n574 10.6151
R1542 B.n575 B.n155 10.6151
R1543 B.n585 B.n155 10.6151
R1544 B.n586 B.n585 10.6151
R1545 B.n587 B.n586 10.6151
R1546 B.n587 B.n147 10.6151
R1547 B.n597 B.n147 10.6151
R1548 B.n598 B.n597 10.6151
R1549 B.n599 B.n598 10.6151
R1550 B.n599 B.n139 10.6151
R1551 B.n609 B.n139 10.6151
R1552 B.n610 B.n609 10.6151
R1553 B.n612 B.n610 10.6151
R1554 B.n612 B.n611 10.6151
R1555 B.n611 B.n131 10.6151
R1556 B.n623 B.n131 10.6151
R1557 B.n624 B.n623 10.6151
R1558 B.n625 B.n624 10.6151
R1559 B.n626 B.n625 10.6151
R1560 B.n627 B.n626 10.6151
R1561 B.n631 B.n627 10.6151
R1562 B.n632 B.n631 10.6151
R1563 B.n633 B.n632 10.6151
R1564 B.n634 B.n633 10.6151
R1565 B.n636 B.n634 10.6151
R1566 B.n637 B.n636 10.6151
R1567 B.n638 B.n637 10.6151
R1568 B.n639 B.n638 10.6151
R1569 B.n641 B.n639 10.6151
R1570 B.n642 B.n641 10.6151
R1571 B.n643 B.n642 10.6151
R1572 B.n644 B.n643 10.6151
R1573 B.n646 B.n644 10.6151
R1574 B.n647 B.n646 10.6151
R1575 B.n648 B.n647 10.6151
R1576 B.n649 B.n648 10.6151
R1577 B.n651 B.n649 10.6151
R1578 B.n652 B.n651 10.6151
R1579 B.n653 B.n652 10.6151
R1580 B.n654 B.n653 10.6151
R1581 B.n656 B.n654 10.6151
R1582 B.n657 B.n656 10.6151
R1583 B.n658 B.n657 10.6151
R1584 B.n659 B.n658 10.6151
R1585 B.n661 B.n659 10.6151
R1586 B.n662 B.n661 10.6151
R1587 B.n663 B.n662 10.6151
R1588 B.n664 B.n663 10.6151
R1589 B.n994 B.n1 10.6151
R1590 B.n994 B.n993 10.6151
R1591 B.n993 B.n992 10.6151
R1592 B.n992 B.n10 10.6151
R1593 B.n986 B.n10 10.6151
R1594 B.n986 B.n985 10.6151
R1595 B.n985 B.n984 10.6151
R1596 B.n984 B.n17 10.6151
R1597 B.n978 B.n17 10.6151
R1598 B.n978 B.n977 10.6151
R1599 B.n977 B.n976 10.6151
R1600 B.n976 B.n24 10.6151
R1601 B.n970 B.n24 10.6151
R1602 B.n970 B.n969 10.6151
R1603 B.n969 B.n968 10.6151
R1604 B.n968 B.n31 10.6151
R1605 B.n962 B.n31 10.6151
R1606 B.n962 B.n961 10.6151
R1607 B.n961 B.n960 10.6151
R1608 B.n960 B.n38 10.6151
R1609 B.n954 B.n38 10.6151
R1610 B.n954 B.n953 10.6151
R1611 B.n953 B.n952 10.6151
R1612 B.n952 B.n45 10.6151
R1613 B.n946 B.n45 10.6151
R1614 B.n946 B.n945 10.6151
R1615 B.n945 B.n944 10.6151
R1616 B.n944 B.n52 10.6151
R1617 B.n938 B.n52 10.6151
R1618 B.n937 B.n936 10.6151
R1619 B.n936 B.n59 10.6151
R1620 B.n930 B.n59 10.6151
R1621 B.n930 B.n929 10.6151
R1622 B.n929 B.n928 10.6151
R1623 B.n928 B.n61 10.6151
R1624 B.n922 B.n61 10.6151
R1625 B.n922 B.n921 10.6151
R1626 B.n921 B.n920 10.6151
R1627 B.n920 B.n63 10.6151
R1628 B.n914 B.n63 10.6151
R1629 B.n914 B.n913 10.6151
R1630 B.n913 B.n912 10.6151
R1631 B.n912 B.n65 10.6151
R1632 B.n906 B.n65 10.6151
R1633 B.n906 B.n905 10.6151
R1634 B.n905 B.n904 10.6151
R1635 B.n904 B.n67 10.6151
R1636 B.n898 B.n67 10.6151
R1637 B.n898 B.n897 10.6151
R1638 B.n897 B.n896 10.6151
R1639 B.n896 B.n69 10.6151
R1640 B.n890 B.n69 10.6151
R1641 B.n890 B.n889 10.6151
R1642 B.n889 B.n888 10.6151
R1643 B.n888 B.n71 10.6151
R1644 B.n882 B.n71 10.6151
R1645 B.n882 B.n881 10.6151
R1646 B.n881 B.n880 10.6151
R1647 B.n880 B.n73 10.6151
R1648 B.n874 B.n73 10.6151
R1649 B.n874 B.n873 10.6151
R1650 B.n873 B.n872 10.6151
R1651 B.n872 B.n75 10.6151
R1652 B.n866 B.n75 10.6151
R1653 B.n866 B.n865 10.6151
R1654 B.n865 B.n864 10.6151
R1655 B.n864 B.n77 10.6151
R1656 B.n858 B.n77 10.6151
R1657 B.n858 B.n857 10.6151
R1658 B.n857 B.n856 10.6151
R1659 B.n856 B.n79 10.6151
R1660 B.n850 B.n79 10.6151
R1661 B.n850 B.n849 10.6151
R1662 B.n849 B.n848 10.6151
R1663 B.n848 B.n81 10.6151
R1664 B.n842 B.n81 10.6151
R1665 B.n842 B.n841 10.6151
R1666 B.n841 B.n840 10.6151
R1667 B.n840 B.n83 10.6151
R1668 B.n834 B.n83 10.6151
R1669 B.n834 B.n833 10.6151
R1670 B.n833 B.n832 10.6151
R1671 B.n832 B.n85 10.6151
R1672 B.n826 B.n85 10.6151
R1673 B.n826 B.n825 10.6151
R1674 B.n825 B.n824 10.6151
R1675 B.n824 B.n87 10.6151
R1676 B.n818 B.n87 10.6151
R1677 B.n818 B.n817 10.6151
R1678 B.n817 B.n816 10.6151
R1679 B.n816 B.n89 10.6151
R1680 B.n810 B.n809 10.6151
R1681 B.n809 B.n808 10.6151
R1682 B.n808 B.n94 10.6151
R1683 B.n802 B.n94 10.6151
R1684 B.n802 B.n801 10.6151
R1685 B.n801 B.n800 10.6151
R1686 B.n800 B.n96 10.6151
R1687 B.n794 B.n96 10.6151
R1688 B.n794 B.n793 10.6151
R1689 B.n791 B.n100 10.6151
R1690 B.n785 B.n100 10.6151
R1691 B.n785 B.n784 10.6151
R1692 B.n784 B.n783 10.6151
R1693 B.n783 B.n102 10.6151
R1694 B.n777 B.n102 10.6151
R1695 B.n777 B.n776 10.6151
R1696 B.n776 B.n775 10.6151
R1697 B.n775 B.n104 10.6151
R1698 B.n769 B.n104 10.6151
R1699 B.n769 B.n768 10.6151
R1700 B.n768 B.n767 10.6151
R1701 B.n767 B.n106 10.6151
R1702 B.n761 B.n106 10.6151
R1703 B.n761 B.n760 10.6151
R1704 B.n760 B.n759 10.6151
R1705 B.n759 B.n108 10.6151
R1706 B.n753 B.n108 10.6151
R1707 B.n753 B.n752 10.6151
R1708 B.n752 B.n751 10.6151
R1709 B.n751 B.n110 10.6151
R1710 B.n745 B.n110 10.6151
R1711 B.n745 B.n744 10.6151
R1712 B.n744 B.n743 10.6151
R1713 B.n743 B.n112 10.6151
R1714 B.n737 B.n112 10.6151
R1715 B.n737 B.n736 10.6151
R1716 B.n736 B.n735 10.6151
R1717 B.n735 B.n114 10.6151
R1718 B.n729 B.n114 10.6151
R1719 B.n729 B.n728 10.6151
R1720 B.n728 B.n727 10.6151
R1721 B.n727 B.n116 10.6151
R1722 B.n721 B.n116 10.6151
R1723 B.n721 B.n720 10.6151
R1724 B.n720 B.n719 10.6151
R1725 B.n719 B.n118 10.6151
R1726 B.n713 B.n118 10.6151
R1727 B.n713 B.n712 10.6151
R1728 B.n712 B.n711 10.6151
R1729 B.n711 B.n120 10.6151
R1730 B.n705 B.n120 10.6151
R1731 B.n705 B.n704 10.6151
R1732 B.n704 B.n703 10.6151
R1733 B.n703 B.n122 10.6151
R1734 B.n697 B.n122 10.6151
R1735 B.n697 B.n696 10.6151
R1736 B.n696 B.n695 10.6151
R1737 B.n695 B.n124 10.6151
R1738 B.n689 B.n124 10.6151
R1739 B.n689 B.n688 10.6151
R1740 B.n688 B.n687 10.6151
R1741 B.n687 B.n126 10.6151
R1742 B.n681 B.n126 10.6151
R1743 B.n681 B.n680 10.6151
R1744 B.n680 B.n679 10.6151
R1745 B.n679 B.n128 10.6151
R1746 B.n673 B.n128 10.6151
R1747 B.n673 B.n672 10.6151
R1748 B.n672 B.n671 10.6151
R1749 B.n671 B.n130 10.6151
R1750 B.n665 B.n130 10.6151
R1751 B.n408 B.n407 9.36635
R1752 B.n385 B.n231 9.36635
R1753 B.n93 B.n89 9.36635
R1754 B.n792 B.n791 9.36635
R1755 B.n1002 B.n0 8.11757
R1756 B.n1002 B.n1 8.11757
R1757 B.t4 B.n157 4.46388
R1758 B.t0 B.n29 4.46388
R1759 B.n614 B.t2 2.67853
R1760 B.n990 B.t3 2.67853
R1761 B.n407 B.n406 1.24928
R1762 B.n389 B.n231 1.24928
R1763 B.n810 B.n93 1.24928
R1764 B.n793 B.n792 1.24928
R1765 B.n553 B.t11 0.893176
R1766 B.n950 B.t7 0.893176
R1767 VN.n2 VN.t4 328.036
R1768 VN.n14 VN.t2 328.036
R1769 VN.n3 VN.t1 295.454
R1770 VN.n10 VN.t3 295.454
R1771 VN.n15 VN.t0 295.454
R1772 VN.n22 VN.t5 295.454
R1773 VN.n11 VN.n10 177.939
R1774 VN.n23 VN.n22 177.939
R1775 VN.n21 VN.n12 161.3
R1776 VN.n20 VN.n19 161.3
R1777 VN.n18 VN.n13 161.3
R1778 VN.n17 VN.n16 161.3
R1779 VN.n9 VN.n0 161.3
R1780 VN.n8 VN.n7 161.3
R1781 VN.n6 VN.n1 161.3
R1782 VN.n5 VN.n4 161.3
R1783 VN.n8 VN.n1 56.5193
R1784 VN.n20 VN.n13 56.5193
R1785 VN.n3 VN.n2 53.9242
R1786 VN.n15 VN.n14 53.9242
R1787 VN VN.n23 50.5516
R1788 VN.n4 VN.n1 24.4675
R1789 VN.n9 VN.n8 24.4675
R1790 VN.n16 VN.n13 24.4675
R1791 VN.n21 VN.n20 24.4675
R1792 VN.n17 VN.n14 17.9992
R1793 VN.n5 VN.n2 17.9992
R1794 VN.n4 VN.n3 12.234
R1795 VN.n16 VN.n15 12.234
R1796 VN.n10 VN.n9 7.82994
R1797 VN.n22 VN.n21 7.82994
R1798 VN.n23 VN.n12 0.189894
R1799 VN.n19 VN.n12 0.189894
R1800 VN.n19 VN.n18 0.189894
R1801 VN.n18 VN.n17 0.189894
R1802 VN.n6 VN.n5 0.189894
R1803 VN.n7 VN.n6 0.189894
R1804 VN.n7 VN.n0 0.189894
R1805 VN.n11 VN.n0 0.189894
R1806 VN VN.n11 0.0516364
R1807 VDD2.n1 VDD2.t1 63.7824
R1808 VDD2.n2 VDD2.t0 62.603
R1809 VDD2.n1 VDD2.n0 61.9371
R1810 VDD2 VDD2.n3 61.9341
R1811 VDD2.n2 VDD2.n1 45.7649
R1812 VDD2 VDD2.n2 1.2936
R1813 VDD2.n3 VDD2.t5 1.0227
R1814 VDD2.n3 VDD2.t3 1.0227
R1815 VDD2.n0 VDD2.t4 1.0227
R1816 VDD2.n0 VDD2.t2 1.0227
C0 VDD2 VDD1 1.0391f
C1 VN VTAIL 9.033191f
C2 VN VDD2 9.41275f
C3 VTAIL VP 9.047781f
C4 VDD2 VP 0.372827f
C5 VN VDD1 0.149412f
C6 VTAIL VDD2 11.2619f
C7 VP VDD1 9.63072f
C8 VN VP 7.30025f
C9 VTAIL VDD1 11.222f
C10 VDD2 B 6.495961f
C11 VDD1 B 6.769022f
C12 VTAIL B 9.946615f
C13 VN B 10.71558f
C14 VP B 8.912826f
C15 VDD2.t1 B 3.86242f
C16 VDD2.t4 B 0.329952f
C17 VDD2.t2 B 0.329952f
C18 VDD2.n0 B 3.0169f
C19 VDD2.n1 B 2.52788f
C20 VDD2.t0 B 3.85634f
C21 VDD2.n2 B 2.66028f
C22 VDD2.t5 B 0.329952f
C23 VDD2.t3 B 0.329952f
C24 VDD2.n3 B 3.01687f
C25 VN.n0 B 0.030443f
C26 VN.t3 B 2.56615f
C27 VN.n1 B 0.040627f
C28 VN.t4 B 2.66756f
C29 VN.n2 B 0.974464f
C30 VN.t1 B 2.56615f
C31 VN.n3 B 0.957073f
C32 VN.n4 B 0.042733f
C33 VN.n5 B 0.193467f
C34 VN.n6 B 0.030443f
C35 VN.n7 B 0.030443f
C36 VN.n8 B 0.048262f
C37 VN.n9 B 0.03769f
C38 VN.n10 B 0.961997f
C39 VN.n11 B 0.030155f
C40 VN.n12 B 0.030443f
C41 VN.t5 B 2.56615f
C42 VN.n13 B 0.040627f
C43 VN.t2 B 2.66756f
C44 VN.n14 B 0.974464f
C45 VN.t0 B 2.56615f
C46 VN.n15 B 0.957073f
C47 VN.n16 B 0.042733f
C48 VN.n17 B 0.193467f
C49 VN.n18 B 0.030443f
C50 VN.n19 B 0.030443f
C51 VN.n20 B 0.048262f
C52 VN.n21 B 0.03769f
C53 VN.n22 B 0.961997f
C54 VN.n23 B 1.68997f
C55 VTAIL.t3 B 0.33976f
C56 VTAIL.t5 B 0.33976f
C57 VTAIL.n0 B 3.0376f
C58 VTAIL.n1 B 0.347673f
C59 VTAIL.t7 B 3.88353f
C60 VTAIL.n2 B 0.512522f
C61 VTAIL.t6 B 0.33976f
C62 VTAIL.t9 B 0.33976f
C63 VTAIL.n3 B 3.0376f
C64 VTAIL.n4 B 2.07071f
C65 VTAIL.t4 B 0.33976f
C66 VTAIL.t1 B 0.33976f
C67 VTAIL.n5 B 3.03759f
C68 VTAIL.n6 B 2.07071f
C69 VTAIL.t2 B 3.88354f
C70 VTAIL.n7 B 0.512518f
C71 VTAIL.t10 B 0.33976f
C72 VTAIL.t11 B 0.33976f
C73 VTAIL.n8 B 3.03759f
C74 VTAIL.n9 B 0.431843f
C75 VTAIL.t8 B 3.88353f
C76 VTAIL.n10 B 2.03363f
C77 VTAIL.t0 B 3.88353f
C78 VTAIL.n11 B 2.00002f
C79 VDD1.t5 B 3.86694f
C80 VDD1.t4 B 3.86621f
C81 VDD1.t1 B 0.330276f
C82 VDD1.t2 B 0.330276f
C83 VDD1.n0 B 3.01986f
C84 VDD1.n1 B 2.61805f
C85 VDD1.t3 B 0.330276f
C86 VDD1.t0 B 0.330276f
C87 VDD1.n2 B 3.01796f
C88 VDD1.n3 B 2.64547f
C89 VP.n0 B 0.030732f
C90 VP.t4 B 2.59044f
C91 VP.n1 B 0.041012f
C92 VP.n2 B 0.030732f
C93 VP.t2 B 2.59044f
C94 VP.n3 B 0.048719f
C95 VP.n4 B 0.030732f
C96 VP.t3 B 2.59044f
C97 VP.n5 B 0.041012f
C98 VP.t1 B 2.69281f
C99 VP.n6 B 0.983685f
C100 VP.t0 B 2.59044f
C101 VP.n7 B 0.96613f
C102 VP.n8 B 0.043137f
C103 VP.n9 B 0.195298f
C104 VP.n10 B 0.030732f
C105 VP.n11 B 0.030732f
C106 VP.n12 B 0.048719f
C107 VP.n13 B 0.038047f
C108 VP.n14 B 0.9711f
C109 VP.n15 B 1.68599f
C110 VP.n16 B 1.70801f
C111 VP.t5 B 2.59044f
C112 VP.n17 B 0.9711f
C113 VP.n18 B 0.038047f
C114 VP.n19 B 0.030732f
C115 VP.n20 B 0.030732f
C116 VP.n21 B 0.030732f
C117 VP.n22 B 0.041012f
C118 VP.n23 B 0.043137f
C119 VP.n24 B 0.906876f
C120 VP.n25 B 0.043137f
C121 VP.n26 B 0.030732f
C122 VP.n27 B 0.030732f
C123 VP.n28 B 0.030732f
C124 VP.n29 B 0.048719f
C125 VP.n30 B 0.038047f
C126 VP.n31 B 0.9711f
C127 VP.n32 B 0.03044f
.ends

