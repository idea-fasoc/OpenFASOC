* NGSPICE file created from diff_pair_sample_0071.ext - technology: sky130A

.subckt diff_pair_sample_0071 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6224 pd=9.1 as=0 ps=0 w=4.16 l=1.38
X1 VTAIL.t7 VN.t0 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6224 pd=9.1 as=0.6864 ps=4.49 w=4.16 l=1.38
X2 VTAIL.t6 VN.t1 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6224 pd=9.1 as=0.6864 ps=4.49 w=4.16 l=1.38
X3 VDD1.t3 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=4.49 as=1.6224 ps=9.1 w=4.16 l=1.38
X4 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=1.6224 pd=9.1 as=0 ps=0 w=4.16 l=1.38
X5 VDD2.t3 VN.t2 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=4.49 as=1.6224 ps=9.1 w=4.16 l=1.38
X6 VTAIL.t3 VP.t1 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6224 pd=9.1 as=0.6864 ps=4.49 w=4.16 l=1.38
X7 VTAIL.t0 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6224 pd=9.1 as=0.6864 ps=4.49 w=4.16 l=1.38
X8 VDD2.t2 VN.t3 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=4.49 as=1.6224 ps=9.1 w=4.16 l=1.38
X9 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.6224 pd=9.1 as=0 ps=0 w=4.16 l=1.38
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6224 pd=9.1 as=0 ps=0 w=4.16 l=1.38
X11 VDD1.t0 VP.t3 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.6864 pd=4.49 as=1.6224 ps=9.1 w=4.16 l=1.38
R0 B.n430 B.n429 585
R1 B.n431 B.n430 585
R2 B.n163 B.n69 585
R3 B.n162 B.n161 585
R4 B.n160 B.n159 585
R5 B.n158 B.n157 585
R6 B.n156 B.n155 585
R7 B.n154 B.n153 585
R8 B.n152 B.n151 585
R9 B.n150 B.n149 585
R10 B.n148 B.n147 585
R11 B.n146 B.n145 585
R12 B.n144 B.n143 585
R13 B.n142 B.n141 585
R14 B.n140 B.n139 585
R15 B.n138 B.n137 585
R16 B.n136 B.n135 585
R17 B.n134 B.n133 585
R18 B.n132 B.n131 585
R19 B.n130 B.n129 585
R20 B.n128 B.n127 585
R21 B.n126 B.n125 585
R22 B.n124 B.n123 585
R23 B.n122 B.n121 585
R24 B.n120 B.n119 585
R25 B.n118 B.n117 585
R26 B.n116 B.n115 585
R27 B.n114 B.n113 585
R28 B.n112 B.n111 585
R29 B.n109 B.n108 585
R30 B.n107 B.n106 585
R31 B.n105 B.n104 585
R32 B.n103 B.n102 585
R33 B.n101 B.n100 585
R34 B.n99 B.n98 585
R35 B.n97 B.n96 585
R36 B.n95 B.n94 585
R37 B.n93 B.n92 585
R38 B.n91 B.n90 585
R39 B.n89 B.n88 585
R40 B.n87 B.n86 585
R41 B.n85 B.n84 585
R42 B.n83 B.n82 585
R43 B.n81 B.n80 585
R44 B.n79 B.n78 585
R45 B.n77 B.n76 585
R46 B.n46 B.n45 585
R47 B.n434 B.n433 585
R48 B.n428 B.n70 585
R49 B.n70 B.n43 585
R50 B.n427 B.n42 585
R51 B.n438 B.n42 585
R52 B.n426 B.n41 585
R53 B.n439 B.n41 585
R54 B.n425 B.n40 585
R55 B.n440 B.n40 585
R56 B.n424 B.n423 585
R57 B.n423 B.n36 585
R58 B.n422 B.n35 585
R59 B.n446 B.n35 585
R60 B.n421 B.n34 585
R61 B.n447 B.n34 585
R62 B.n420 B.n33 585
R63 B.n448 B.n33 585
R64 B.n419 B.n418 585
R65 B.n418 B.n29 585
R66 B.n417 B.n28 585
R67 B.n454 B.n28 585
R68 B.n416 B.n27 585
R69 B.n455 B.n27 585
R70 B.n415 B.n26 585
R71 B.n456 B.n26 585
R72 B.n414 B.n413 585
R73 B.n413 B.n22 585
R74 B.n412 B.n21 585
R75 B.n462 B.n21 585
R76 B.n411 B.n20 585
R77 B.n463 B.n20 585
R78 B.n410 B.n19 585
R79 B.n464 B.n19 585
R80 B.n409 B.n408 585
R81 B.n408 B.n15 585
R82 B.n407 B.n14 585
R83 B.n470 B.n14 585
R84 B.n406 B.n13 585
R85 B.n471 B.n13 585
R86 B.n405 B.n12 585
R87 B.n472 B.n12 585
R88 B.n404 B.n403 585
R89 B.n403 B.n8 585
R90 B.n402 B.n7 585
R91 B.n478 B.n7 585
R92 B.n401 B.n6 585
R93 B.n479 B.n6 585
R94 B.n400 B.n5 585
R95 B.n480 B.n5 585
R96 B.n399 B.n398 585
R97 B.n398 B.n4 585
R98 B.n397 B.n164 585
R99 B.n397 B.n396 585
R100 B.n387 B.n165 585
R101 B.n166 B.n165 585
R102 B.n389 B.n388 585
R103 B.n390 B.n389 585
R104 B.n386 B.n170 585
R105 B.n174 B.n170 585
R106 B.n385 B.n384 585
R107 B.n384 B.n383 585
R108 B.n172 B.n171 585
R109 B.n173 B.n172 585
R110 B.n376 B.n375 585
R111 B.n377 B.n376 585
R112 B.n374 B.n179 585
R113 B.n179 B.n178 585
R114 B.n373 B.n372 585
R115 B.n372 B.n371 585
R116 B.n181 B.n180 585
R117 B.n182 B.n181 585
R118 B.n364 B.n363 585
R119 B.n365 B.n364 585
R120 B.n362 B.n187 585
R121 B.n187 B.n186 585
R122 B.n361 B.n360 585
R123 B.n360 B.n359 585
R124 B.n189 B.n188 585
R125 B.n190 B.n189 585
R126 B.n352 B.n351 585
R127 B.n353 B.n352 585
R128 B.n350 B.n195 585
R129 B.n195 B.n194 585
R130 B.n349 B.n348 585
R131 B.n348 B.n347 585
R132 B.n197 B.n196 585
R133 B.n198 B.n197 585
R134 B.n340 B.n339 585
R135 B.n341 B.n340 585
R136 B.n338 B.n203 585
R137 B.n203 B.n202 585
R138 B.n337 B.n336 585
R139 B.n336 B.n335 585
R140 B.n205 B.n204 585
R141 B.n206 B.n205 585
R142 B.n331 B.n330 585
R143 B.n209 B.n208 585
R144 B.n327 B.n326 585
R145 B.n328 B.n327 585
R146 B.n325 B.n232 585
R147 B.n324 B.n323 585
R148 B.n322 B.n321 585
R149 B.n320 B.n319 585
R150 B.n318 B.n317 585
R151 B.n316 B.n315 585
R152 B.n314 B.n313 585
R153 B.n312 B.n311 585
R154 B.n310 B.n309 585
R155 B.n308 B.n307 585
R156 B.n306 B.n305 585
R157 B.n304 B.n303 585
R158 B.n302 B.n301 585
R159 B.n300 B.n299 585
R160 B.n298 B.n297 585
R161 B.n296 B.n295 585
R162 B.n294 B.n293 585
R163 B.n292 B.n291 585
R164 B.n290 B.n289 585
R165 B.n288 B.n287 585
R166 B.n286 B.n285 585
R167 B.n284 B.n283 585
R168 B.n282 B.n281 585
R169 B.n280 B.n279 585
R170 B.n278 B.n277 585
R171 B.n275 B.n274 585
R172 B.n273 B.n272 585
R173 B.n271 B.n270 585
R174 B.n269 B.n268 585
R175 B.n267 B.n266 585
R176 B.n265 B.n264 585
R177 B.n263 B.n262 585
R178 B.n261 B.n260 585
R179 B.n259 B.n258 585
R180 B.n257 B.n256 585
R181 B.n255 B.n254 585
R182 B.n253 B.n252 585
R183 B.n251 B.n250 585
R184 B.n249 B.n248 585
R185 B.n247 B.n246 585
R186 B.n245 B.n244 585
R187 B.n243 B.n242 585
R188 B.n241 B.n240 585
R189 B.n239 B.n238 585
R190 B.n332 B.n207 585
R191 B.n207 B.n206 585
R192 B.n334 B.n333 585
R193 B.n335 B.n334 585
R194 B.n201 B.n200 585
R195 B.n202 B.n201 585
R196 B.n343 B.n342 585
R197 B.n342 B.n341 585
R198 B.n344 B.n199 585
R199 B.n199 B.n198 585
R200 B.n346 B.n345 585
R201 B.n347 B.n346 585
R202 B.n193 B.n192 585
R203 B.n194 B.n193 585
R204 B.n355 B.n354 585
R205 B.n354 B.n353 585
R206 B.n356 B.n191 585
R207 B.n191 B.n190 585
R208 B.n358 B.n357 585
R209 B.n359 B.n358 585
R210 B.n185 B.n184 585
R211 B.n186 B.n185 585
R212 B.n367 B.n366 585
R213 B.n366 B.n365 585
R214 B.n368 B.n183 585
R215 B.n183 B.n182 585
R216 B.n370 B.n369 585
R217 B.n371 B.n370 585
R218 B.n177 B.n176 585
R219 B.n178 B.n177 585
R220 B.n379 B.n378 585
R221 B.n378 B.n377 585
R222 B.n380 B.n175 585
R223 B.n175 B.n173 585
R224 B.n382 B.n381 585
R225 B.n383 B.n382 585
R226 B.n169 B.n168 585
R227 B.n174 B.n169 585
R228 B.n392 B.n391 585
R229 B.n391 B.n390 585
R230 B.n393 B.n167 585
R231 B.n167 B.n166 585
R232 B.n395 B.n394 585
R233 B.n396 B.n395 585
R234 B.n2 B.n0 585
R235 B.n4 B.n2 585
R236 B.n3 B.n1 585
R237 B.n479 B.n3 585
R238 B.n477 B.n476 585
R239 B.n478 B.n477 585
R240 B.n475 B.n9 585
R241 B.n9 B.n8 585
R242 B.n474 B.n473 585
R243 B.n473 B.n472 585
R244 B.n11 B.n10 585
R245 B.n471 B.n11 585
R246 B.n469 B.n468 585
R247 B.n470 B.n469 585
R248 B.n467 B.n16 585
R249 B.n16 B.n15 585
R250 B.n466 B.n465 585
R251 B.n465 B.n464 585
R252 B.n18 B.n17 585
R253 B.n463 B.n18 585
R254 B.n461 B.n460 585
R255 B.n462 B.n461 585
R256 B.n459 B.n23 585
R257 B.n23 B.n22 585
R258 B.n458 B.n457 585
R259 B.n457 B.n456 585
R260 B.n25 B.n24 585
R261 B.n455 B.n25 585
R262 B.n453 B.n452 585
R263 B.n454 B.n453 585
R264 B.n451 B.n30 585
R265 B.n30 B.n29 585
R266 B.n450 B.n449 585
R267 B.n449 B.n448 585
R268 B.n32 B.n31 585
R269 B.n447 B.n32 585
R270 B.n445 B.n444 585
R271 B.n446 B.n445 585
R272 B.n443 B.n37 585
R273 B.n37 B.n36 585
R274 B.n442 B.n441 585
R275 B.n441 B.n440 585
R276 B.n39 B.n38 585
R277 B.n439 B.n39 585
R278 B.n437 B.n436 585
R279 B.n438 B.n437 585
R280 B.n435 B.n44 585
R281 B.n44 B.n43 585
R282 B.n482 B.n481 585
R283 B.n481 B.n480 585
R284 B.n330 B.n207 506.916
R285 B.n433 B.n44 506.916
R286 B.n238 B.n205 506.916
R287 B.n430 B.n70 506.916
R288 B.n236 B.t8 277.613
R289 B.n233 B.t12 277.613
R290 B.n74 B.t15 277.613
R291 B.n71 B.t4 277.613
R292 B.n431 B.n68 256.663
R293 B.n431 B.n67 256.663
R294 B.n431 B.n66 256.663
R295 B.n431 B.n65 256.663
R296 B.n431 B.n64 256.663
R297 B.n431 B.n63 256.663
R298 B.n431 B.n62 256.663
R299 B.n431 B.n61 256.663
R300 B.n431 B.n60 256.663
R301 B.n431 B.n59 256.663
R302 B.n431 B.n58 256.663
R303 B.n431 B.n57 256.663
R304 B.n431 B.n56 256.663
R305 B.n431 B.n55 256.663
R306 B.n431 B.n54 256.663
R307 B.n431 B.n53 256.663
R308 B.n431 B.n52 256.663
R309 B.n431 B.n51 256.663
R310 B.n431 B.n50 256.663
R311 B.n431 B.n49 256.663
R312 B.n431 B.n48 256.663
R313 B.n431 B.n47 256.663
R314 B.n432 B.n431 256.663
R315 B.n329 B.n328 256.663
R316 B.n328 B.n210 256.663
R317 B.n328 B.n211 256.663
R318 B.n328 B.n212 256.663
R319 B.n328 B.n213 256.663
R320 B.n328 B.n214 256.663
R321 B.n328 B.n215 256.663
R322 B.n328 B.n216 256.663
R323 B.n328 B.n217 256.663
R324 B.n328 B.n218 256.663
R325 B.n328 B.n219 256.663
R326 B.n328 B.n220 256.663
R327 B.n328 B.n221 256.663
R328 B.n328 B.n222 256.663
R329 B.n328 B.n223 256.663
R330 B.n328 B.n224 256.663
R331 B.n328 B.n225 256.663
R332 B.n328 B.n226 256.663
R333 B.n328 B.n227 256.663
R334 B.n328 B.n228 256.663
R335 B.n328 B.n229 256.663
R336 B.n328 B.n230 256.663
R337 B.n328 B.n231 256.663
R338 B.n334 B.n207 163.367
R339 B.n334 B.n201 163.367
R340 B.n342 B.n201 163.367
R341 B.n342 B.n199 163.367
R342 B.n346 B.n199 163.367
R343 B.n346 B.n193 163.367
R344 B.n354 B.n193 163.367
R345 B.n354 B.n191 163.367
R346 B.n358 B.n191 163.367
R347 B.n358 B.n185 163.367
R348 B.n366 B.n185 163.367
R349 B.n366 B.n183 163.367
R350 B.n370 B.n183 163.367
R351 B.n370 B.n177 163.367
R352 B.n378 B.n177 163.367
R353 B.n378 B.n175 163.367
R354 B.n382 B.n175 163.367
R355 B.n382 B.n169 163.367
R356 B.n391 B.n169 163.367
R357 B.n391 B.n167 163.367
R358 B.n395 B.n167 163.367
R359 B.n395 B.n2 163.367
R360 B.n481 B.n2 163.367
R361 B.n481 B.n3 163.367
R362 B.n477 B.n3 163.367
R363 B.n477 B.n9 163.367
R364 B.n473 B.n9 163.367
R365 B.n473 B.n11 163.367
R366 B.n469 B.n11 163.367
R367 B.n469 B.n16 163.367
R368 B.n465 B.n16 163.367
R369 B.n465 B.n18 163.367
R370 B.n461 B.n18 163.367
R371 B.n461 B.n23 163.367
R372 B.n457 B.n23 163.367
R373 B.n457 B.n25 163.367
R374 B.n453 B.n25 163.367
R375 B.n453 B.n30 163.367
R376 B.n449 B.n30 163.367
R377 B.n449 B.n32 163.367
R378 B.n445 B.n32 163.367
R379 B.n445 B.n37 163.367
R380 B.n441 B.n37 163.367
R381 B.n441 B.n39 163.367
R382 B.n437 B.n39 163.367
R383 B.n437 B.n44 163.367
R384 B.n327 B.n209 163.367
R385 B.n327 B.n232 163.367
R386 B.n323 B.n322 163.367
R387 B.n319 B.n318 163.367
R388 B.n315 B.n314 163.367
R389 B.n311 B.n310 163.367
R390 B.n307 B.n306 163.367
R391 B.n303 B.n302 163.367
R392 B.n299 B.n298 163.367
R393 B.n295 B.n294 163.367
R394 B.n291 B.n290 163.367
R395 B.n287 B.n286 163.367
R396 B.n283 B.n282 163.367
R397 B.n279 B.n278 163.367
R398 B.n274 B.n273 163.367
R399 B.n270 B.n269 163.367
R400 B.n266 B.n265 163.367
R401 B.n262 B.n261 163.367
R402 B.n258 B.n257 163.367
R403 B.n254 B.n253 163.367
R404 B.n250 B.n249 163.367
R405 B.n246 B.n245 163.367
R406 B.n242 B.n241 163.367
R407 B.n336 B.n205 163.367
R408 B.n336 B.n203 163.367
R409 B.n340 B.n203 163.367
R410 B.n340 B.n197 163.367
R411 B.n348 B.n197 163.367
R412 B.n348 B.n195 163.367
R413 B.n352 B.n195 163.367
R414 B.n352 B.n189 163.367
R415 B.n360 B.n189 163.367
R416 B.n360 B.n187 163.367
R417 B.n364 B.n187 163.367
R418 B.n364 B.n181 163.367
R419 B.n372 B.n181 163.367
R420 B.n372 B.n179 163.367
R421 B.n376 B.n179 163.367
R422 B.n376 B.n172 163.367
R423 B.n384 B.n172 163.367
R424 B.n384 B.n170 163.367
R425 B.n389 B.n170 163.367
R426 B.n389 B.n165 163.367
R427 B.n397 B.n165 163.367
R428 B.n398 B.n397 163.367
R429 B.n398 B.n5 163.367
R430 B.n6 B.n5 163.367
R431 B.n7 B.n6 163.367
R432 B.n403 B.n7 163.367
R433 B.n403 B.n12 163.367
R434 B.n13 B.n12 163.367
R435 B.n14 B.n13 163.367
R436 B.n408 B.n14 163.367
R437 B.n408 B.n19 163.367
R438 B.n20 B.n19 163.367
R439 B.n21 B.n20 163.367
R440 B.n413 B.n21 163.367
R441 B.n413 B.n26 163.367
R442 B.n27 B.n26 163.367
R443 B.n28 B.n27 163.367
R444 B.n418 B.n28 163.367
R445 B.n418 B.n33 163.367
R446 B.n34 B.n33 163.367
R447 B.n35 B.n34 163.367
R448 B.n423 B.n35 163.367
R449 B.n423 B.n40 163.367
R450 B.n41 B.n40 163.367
R451 B.n42 B.n41 163.367
R452 B.n70 B.n42 163.367
R453 B.n76 B.n46 163.367
R454 B.n80 B.n79 163.367
R455 B.n84 B.n83 163.367
R456 B.n88 B.n87 163.367
R457 B.n92 B.n91 163.367
R458 B.n96 B.n95 163.367
R459 B.n100 B.n99 163.367
R460 B.n104 B.n103 163.367
R461 B.n108 B.n107 163.367
R462 B.n113 B.n112 163.367
R463 B.n117 B.n116 163.367
R464 B.n121 B.n120 163.367
R465 B.n125 B.n124 163.367
R466 B.n129 B.n128 163.367
R467 B.n133 B.n132 163.367
R468 B.n137 B.n136 163.367
R469 B.n141 B.n140 163.367
R470 B.n145 B.n144 163.367
R471 B.n149 B.n148 163.367
R472 B.n153 B.n152 163.367
R473 B.n157 B.n156 163.367
R474 B.n161 B.n160 163.367
R475 B.n430 B.n69 163.367
R476 B.n328 B.n206 159.725
R477 B.n431 B.n43 159.725
R478 B.n236 B.t11 105.889
R479 B.n71 B.t6 105.889
R480 B.n233 B.t14 105.885
R481 B.n74 B.t16 105.885
R482 B.n335 B.n206 79.2798
R483 B.n335 B.n202 79.2798
R484 B.n341 B.n202 79.2798
R485 B.n341 B.n198 79.2798
R486 B.n347 B.n198 79.2798
R487 B.n353 B.n194 79.2798
R488 B.n353 B.n190 79.2798
R489 B.n359 B.n190 79.2798
R490 B.n359 B.n186 79.2798
R491 B.n365 B.n186 79.2798
R492 B.n365 B.n182 79.2798
R493 B.n371 B.n182 79.2798
R494 B.n377 B.n178 79.2798
R495 B.n377 B.n173 79.2798
R496 B.n383 B.n173 79.2798
R497 B.n383 B.n174 79.2798
R498 B.n390 B.n166 79.2798
R499 B.n396 B.n166 79.2798
R500 B.n396 B.n4 79.2798
R501 B.n480 B.n4 79.2798
R502 B.n480 B.n479 79.2798
R503 B.n479 B.n478 79.2798
R504 B.n478 B.n8 79.2798
R505 B.n472 B.n8 79.2798
R506 B.n471 B.n470 79.2798
R507 B.n470 B.n15 79.2798
R508 B.n464 B.n15 79.2798
R509 B.n464 B.n463 79.2798
R510 B.n462 B.n22 79.2798
R511 B.n456 B.n22 79.2798
R512 B.n456 B.n455 79.2798
R513 B.n455 B.n454 79.2798
R514 B.n454 B.n29 79.2798
R515 B.n448 B.n29 79.2798
R516 B.n448 B.n447 79.2798
R517 B.n446 B.n36 79.2798
R518 B.n440 B.n36 79.2798
R519 B.n440 B.n439 79.2798
R520 B.n439 B.n438 79.2798
R521 B.n438 B.n43 79.2798
R522 B.n237 B.t10 72.7256
R523 B.n72 B.t7 72.7256
R524 B.n234 B.t13 72.7218
R525 B.n75 B.t17 72.7218
R526 B.n330 B.n329 71.676
R527 B.n232 B.n210 71.676
R528 B.n322 B.n211 71.676
R529 B.n318 B.n212 71.676
R530 B.n314 B.n213 71.676
R531 B.n310 B.n214 71.676
R532 B.n306 B.n215 71.676
R533 B.n302 B.n216 71.676
R534 B.n298 B.n217 71.676
R535 B.n294 B.n218 71.676
R536 B.n290 B.n219 71.676
R537 B.n286 B.n220 71.676
R538 B.n282 B.n221 71.676
R539 B.n278 B.n222 71.676
R540 B.n273 B.n223 71.676
R541 B.n269 B.n224 71.676
R542 B.n265 B.n225 71.676
R543 B.n261 B.n226 71.676
R544 B.n257 B.n227 71.676
R545 B.n253 B.n228 71.676
R546 B.n249 B.n229 71.676
R547 B.n245 B.n230 71.676
R548 B.n241 B.n231 71.676
R549 B.n433 B.n432 71.676
R550 B.n76 B.n47 71.676
R551 B.n80 B.n48 71.676
R552 B.n84 B.n49 71.676
R553 B.n88 B.n50 71.676
R554 B.n92 B.n51 71.676
R555 B.n96 B.n52 71.676
R556 B.n100 B.n53 71.676
R557 B.n104 B.n54 71.676
R558 B.n108 B.n55 71.676
R559 B.n113 B.n56 71.676
R560 B.n117 B.n57 71.676
R561 B.n121 B.n58 71.676
R562 B.n125 B.n59 71.676
R563 B.n129 B.n60 71.676
R564 B.n133 B.n61 71.676
R565 B.n137 B.n62 71.676
R566 B.n141 B.n63 71.676
R567 B.n145 B.n64 71.676
R568 B.n149 B.n65 71.676
R569 B.n153 B.n66 71.676
R570 B.n157 B.n67 71.676
R571 B.n161 B.n68 71.676
R572 B.n69 B.n68 71.676
R573 B.n160 B.n67 71.676
R574 B.n156 B.n66 71.676
R575 B.n152 B.n65 71.676
R576 B.n148 B.n64 71.676
R577 B.n144 B.n63 71.676
R578 B.n140 B.n62 71.676
R579 B.n136 B.n61 71.676
R580 B.n132 B.n60 71.676
R581 B.n128 B.n59 71.676
R582 B.n124 B.n58 71.676
R583 B.n120 B.n57 71.676
R584 B.n116 B.n56 71.676
R585 B.n112 B.n55 71.676
R586 B.n107 B.n54 71.676
R587 B.n103 B.n53 71.676
R588 B.n99 B.n52 71.676
R589 B.n95 B.n51 71.676
R590 B.n91 B.n50 71.676
R591 B.n87 B.n49 71.676
R592 B.n83 B.n48 71.676
R593 B.n79 B.n47 71.676
R594 B.n432 B.n46 71.676
R595 B.n329 B.n209 71.676
R596 B.n323 B.n210 71.676
R597 B.n319 B.n211 71.676
R598 B.n315 B.n212 71.676
R599 B.n311 B.n213 71.676
R600 B.n307 B.n214 71.676
R601 B.n303 B.n215 71.676
R602 B.n299 B.n216 71.676
R603 B.n295 B.n217 71.676
R604 B.n291 B.n218 71.676
R605 B.n287 B.n219 71.676
R606 B.n283 B.n220 71.676
R607 B.n279 B.n221 71.676
R608 B.n274 B.n222 71.676
R609 B.n270 B.n223 71.676
R610 B.n266 B.n224 71.676
R611 B.n262 B.n225 71.676
R612 B.n258 B.n226 71.676
R613 B.n254 B.n227 71.676
R614 B.n250 B.n228 71.676
R615 B.n246 B.n229 71.676
R616 B.n242 B.n230 71.676
R617 B.n238 B.n231 71.676
R618 B.n174 B.t2 69.9528
R619 B.t1 B.n471 69.9528
R620 B.n371 B.t3 67.6211
R621 B.t0 B.n462 67.6211
R622 B.n276 B.n237 59.5399
R623 B.n235 B.n234 59.5399
R624 B.n110 B.n75 59.5399
R625 B.n73 B.n72 59.5399
R626 B.n347 B.t9 48.9671
R627 B.t5 B.n446 48.9671
R628 B.n237 B.n236 33.1641
R629 B.n234 B.n233 33.1641
R630 B.n75 B.n74 33.1641
R631 B.n72 B.n71 33.1641
R632 B.n435 B.n434 32.9371
R633 B.n429 B.n428 32.9371
R634 B.n239 B.n204 32.9371
R635 B.n332 B.n331 32.9371
R636 B.t9 B.n194 30.3132
R637 B.n447 B.t5 30.3132
R638 B B.n482 18.0485
R639 B.t3 B.n178 11.6592
R640 B.n463 B.t0 11.6592
R641 B.n434 B.n45 10.6151
R642 B.n77 B.n45 10.6151
R643 B.n78 B.n77 10.6151
R644 B.n81 B.n78 10.6151
R645 B.n82 B.n81 10.6151
R646 B.n85 B.n82 10.6151
R647 B.n86 B.n85 10.6151
R648 B.n89 B.n86 10.6151
R649 B.n90 B.n89 10.6151
R650 B.n93 B.n90 10.6151
R651 B.n94 B.n93 10.6151
R652 B.n97 B.n94 10.6151
R653 B.n98 B.n97 10.6151
R654 B.n101 B.n98 10.6151
R655 B.n102 B.n101 10.6151
R656 B.n105 B.n102 10.6151
R657 B.n106 B.n105 10.6151
R658 B.n109 B.n106 10.6151
R659 B.n114 B.n111 10.6151
R660 B.n115 B.n114 10.6151
R661 B.n118 B.n115 10.6151
R662 B.n119 B.n118 10.6151
R663 B.n122 B.n119 10.6151
R664 B.n123 B.n122 10.6151
R665 B.n126 B.n123 10.6151
R666 B.n127 B.n126 10.6151
R667 B.n131 B.n130 10.6151
R668 B.n134 B.n131 10.6151
R669 B.n135 B.n134 10.6151
R670 B.n138 B.n135 10.6151
R671 B.n139 B.n138 10.6151
R672 B.n142 B.n139 10.6151
R673 B.n143 B.n142 10.6151
R674 B.n146 B.n143 10.6151
R675 B.n147 B.n146 10.6151
R676 B.n150 B.n147 10.6151
R677 B.n151 B.n150 10.6151
R678 B.n154 B.n151 10.6151
R679 B.n155 B.n154 10.6151
R680 B.n158 B.n155 10.6151
R681 B.n159 B.n158 10.6151
R682 B.n162 B.n159 10.6151
R683 B.n163 B.n162 10.6151
R684 B.n429 B.n163 10.6151
R685 B.n337 B.n204 10.6151
R686 B.n338 B.n337 10.6151
R687 B.n339 B.n338 10.6151
R688 B.n339 B.n196 10.6151
R689 B.n349 B.n196 10.6151
R690 B.n350 B.n349 10.6151
R691 B.n351 B.n350 10.6151
R692 B.n351 B.n188 10.6151
R693 B.n361 B.n188 10.6151
R694 B.n362 B.n361 10.6151
R695 B.n363 B.n362 10.6151
R696 B.n363 B.n180 10.6151
R697 B.n373 B.n180 10.6151
R698 B.n374 B.n373 10.6151
R699 B.n375 B.n374 10.6151
R700 B.n375 B.n171 10.6151
R701 B.n385 B.n171 10.6151
R702 B.n386 B.n385 10.6151
R703 B.n388 B.n386 10.6151
R704 B.n388 B.n387 10.6151
R705 B.n387 B.n164 10.6151
R706 B.n399 B.n164 10.6151
R707 B.n400 B.n399 10.6151
R708 B.n401 B.n400 10.6151
R709 B.n402 B.n401 10.6151
R710 B.n404 B.n402 10.6151
R711 B.n405 B.n404 10.6151
R712 B.n406 B.n405 10.6151
R713 B.n407 B.n406 10.6151
R714 B.n409 B.n407 10.6151
R715 B.n410 B.n409 10.6151
R716 B.n411 B.n410 10.6151
R717 B.n412 B.n411 10.6151
R718 B.n414 B.n412 10.6151
R719 B.n415 B.n414 10.6151
R720 B.n416 B.n415 10.6151
R721 B.n417 B.n416 10.6151
R722 B.n419 B.n417 10.6151
R723 B.n420 B.n419 10.6151
R724 B.n421 B.n420 10.6151
R725 B.n422 B.n421 10.6151
R726 B.n424 B.n422 10.6151
R727 B.n425 B.n424 10.6151
R728 B.n426 B.n425 10.6151
R729 B.n427 B.n426 10.6151
R730 B.n428 B.n427 10.6151
R731 B.n331 B.n208 10.6151
R732 B.n326 B.n208 10.6151
R733 B.n326 B.n325 10.6151
R734 B.n325 B.n324 10.6151
R735 B.n324 B.n321 10.6151
R736 B.n321 B.n320 10.6151
R737 B.n320 B.n317 10.6151
R738 B.n317 B.n316 10.6151
R739 B.n316 B.n313 10.6151
R740 B.n313 B.n312 10.6151
R741 B.n312 B.n309 10.6151
R742 B.n309 B.n308 10.6151
R743 B.n308 B.n305 10.6151
R744 B.n305 B.n304 10.6151
R745 B.n304 B.n301 10.6151
R746 B.n301 B.n300 10.6151
R747 B.n300 B.n297 10.6151
R748 B.n297 B.n296 10.6151
R749 B.n293 B.n292 10.6151
R750 B.n292 B.n289 10.6151
R751 B.n289 B.n288 10.6151
R752 B.n288 B.n285 10.6151
R753 B.n285 B.n284 10.6151
R754 B.n284 B.n281 10.6151
R755 B.n281 B.n280 10.6151
R756 B.n280 B.n277 10.6151
R757 B.n275 B.n272 10.6151
R758 B.n272 B.n271 10.6151
R759 B.n271 B.n268 10.6151
R760 B.n268 B.n267 10.6151
R761 B.n267 B.n264 10.6151
R762 B.n264 B.n263 10.6151
R763 B.n263 B.n260 10.6151
R764 B.n260 B.n259 10.6151
R765 B.n259 B.n256 10.6151
R766 B.n256 B.n255 10.6151
R767 B.n255 B.n252 10.6151
R768 B.n252 B.n251 10.6151
R769 B.n251 B.n248 10.6151
R770 B.n248 B.n247 10.6151
R771 B.n247 B.n244 10.6151
R772 B.n244 B.n243 10.6151
R773 B.n243 B.n240 10.6151
R774 B.n240 B.n239 10.6151
R775 B.n333 B.n332 10.6151
R776 B.n333 B.n200 10.6151
R777 B.n343 B.n200 10.6151
R778 B.n344 B.n343 10.6151
R779 B.n345 B.n344 10.6151
R780 B.n345 B.n192 10.6151
R781 B.n355 B.n192 10.6151
R782 B.n356 B.n355 10.6151
R783 B.n357 B.n356 10.6151
R784 B.n357 B.n184 10.6151
R785 B.n367 B.n184 10.6151
R786 B.n368 B.n367 10.6151
R787 B.n369 B.n368 10.6151
R788 B.n369 B.n176 10.6151
R789 B.n379 B.n176 10.6151
R790 B.n380 B.n379 10.6151
R791 B.n381 B.n380 10.6151
R792 B.n381 B.n168 10.6151
R793 B.n392 B.n168 10.6151
R794 B.n393 B.n392 10.6151
R795 B.n394 B.n393 10.6151
R796 B.n394 B.n0 10.6151
R797 B.n476 B.n1 10.6151
R798 B.n476 B.n475 10.6151
R799 B.n475 B.n474 10.6151
R800 B.n474 B.n10 10.6151
R801 B.n468 B.n10 10.6151
R802 B.n468 B.n467 10.6151
R803 B.n467 B.n466 10.6151
R804 B.n466 B.n17 10.6151
R805 B.n460 B.n17 10.6151
R806 B.n460 B.n459 10.6151
R807 B.n459 B.n458 10.6151
R808 B.n458 B.n24 10.6151
R809 B.n452 B.n24 10.6151
R810 B.n452 B.n451 10.6151
R811 B.n451 B.n450 10.6151
R812 B.n450 B.n31 10.6151
R813 B.n444 B.n31 10.6151
R814 B.n444 B.n443 10.6151
R815 B.n443 B.n442 10.6151
R816 B.n442 B.n38 10.6151
R817 B.n436 B.n38 10.6151
R818 B.n436 B.n435 10.6151
R819 B.n390 B.t2 9.32747
R820 B.n472 B.t1 9.32747
R821 B.n111 B.n110 6.5566
R822 B.n127 B.n73 6.5566
R823 B.n293 B.n235 6.5566
R824 B.n277 B.n276 6.5566
R825 B.n110 B.n109 4.05904
R826 B.n130 B.n73 4.05904
R827 B.n296 B.n235 4.05904
R828 B.n276 B.n275 4.05904
R829 B.n482 B.n0 2.81026
R830 B.n482 B.n1 2.81026
R831 VN.n0 VN.t1 111.29
R832 VN.n1 VN.t3 111.29
R833 VN.n0 VN.t2 111.056
R834 VN.n1 VN.t0 111.056
R835 VN VN.n1 54.5602
R836 VN VN.n0 17.564
R837 VDD2.n2 VDD2.n0 102.865
R838 VDD2.n2 VDD2.n1 71.1425
R839 VDD2.n1 VDD2.t0 4.76012
R840 VDD2.n1 VDD2.t2 4.76012
R841 VDD2.n0 VDD2.t1 4.76012
R842 VDD2.n0 VDD2.t3 4.76012
R843 VDD2 VDD2.n2 0.0586897
R844 VTAIL.n5 VTAIL.t0 59.2235
R845 VTAIL.n4 VTAIL.t4 59.2235
R846 VTAIL.n3 VTAIL.t7 59.2235
R847 VTAIL.n6 VTAIL.t1 59.2233
R848 VTAIL.n7 VTAIL.t5 59.2233
R849 VTAIL.n0 VTAIL.t6 59.2233
R850 VTAIL.n1 VTAIL.t2 59.2233
R851 VTAIL.n2 VTAIL.t3 59.2233
R852 VTAIL.n7 VTAIL.n6 17.4272
R853 VTAIL.n3 VTAIL.n2 17.4272
R854 VTAIL.n4 VTAIL.n3 1.47464
R855 VTAIL.n6 VTAIL.n5 1.47464
R856 VTAIL.n2 VTAIL.n1 1.47464
R857 VTAIL VTAIL.n0 0.795759
R858 VTAIL VTAIL.n7 0.679379
R859 VTAIL.n5 VTAIL.n4 0.470328
R860 VTAIL.n1 VTAIL.n0 0.470328
R861 VP.n4 VP.n3 168.433
R862 VP.n10 VP.n9 168.433
R863 VP.n8 VP.n0 161.3
R864 VP.n7 VP.n6 161.3
R865 VP.n5 VP.n1 161.3
R866 VP.n2 VP.t2 111.29
R867 VP.n2 VP.t3 111.056
R868 VP.n3 VP.t1 72.6498
R869 VP.n9 VP.t0 72.6498
R870 VP.n4 VP.n2 54.1795
R871 VP.n7 VP.n1 40.577
R872 VP.n8 VP.n7 40.577
R873 VP.n3 VP.n1 17.4607
R874 VP.n9 VP.n8 17.4607
R875 VP.n5 VP.n4 0.189894
R876 VP.n6 VP.n5 0.189894
R877 VP.n6 VP.n0 0.189894
R878 VP.n10 VP.n0 0.189894
R879 VP VP.n10 0.0516364
R880 VDD1 VDD1.n1 103.391
R881 VDD1 VDD1.n0 71.2007
R882 VDD1.n0 VDD1.t1 4.76012
R883 VDD1.n0 VDD1.t0 4.76012
R884 VDD1.n1 VDD1.t2 4.76012
R885 VDD1.n1 VDD1.t3 4.76012
C0 VN VP 3.85905f
C1 VTAIL VN 1.74967f
C2 VDD1 VN 0.152218f
C3 VDD2 VP 0.321353f
C4 VDD2 VTAIL 3.19934f
C5 VDD2 VDD1 0.728177f
C6 VTAIL VP 1.76378f
C7 VDD1 VP 1.78722f
C8 VDD1 VTAIL 3.15332f
C9 VDD2 VN 1.61888f
C10 VDD2 B 2.415358f
C11 VDD1 B 4.35045f
C12 VTAIL B 4.516457f
C13 VN B 6.89174f
C14 VP B 5.660497f
C15 VDD1.t1 B 0.058116f
C16 VDD1.t0 B 0.058116f
C17 VDD1.n0 B 0.460389f
C18 VDD1.t2 B 0.058116f
C19 VDD1.t3 B 0.058116f
C20 VDD1.n1 B 0.692572f
C21 VP.n0 B 0.022073f
C22 VP.t0 B 0.326663f
C23 VP.n1 B 0.037779f
C24 VP.t2 B 0.403185f
C25 VP.t3 B 0.402719f
C26 VP.n2 B 0.869008f
C27 VP.t1 B 0.326663f
C28 VP.n3 B 0.186874f
C29 VP.n4 B 1.00618f
C30 VP.n5 B 0.022073f
C31 VP.n6 B 0.022073f
C32 VP.n7 B 0.017827f
C33 VP.n8 B 0.037779f
C34 VP.n9 B 0.186874f
C35 VP.n10 B 0.019241f
C36 VTAIL.t6 B 0.391808f
C37 VTAIL.n0 B 0.196496f
C38 VTAIL.t2 B 0.391808f
C39 VTAIL.n1 B 0.224776f
C40 VTAIL.t3 B 0.391808f
C41 VTAIL.n2 B 0.591608f
C42 VTAIL.t7 B 0.39181f
C43 VTAIL.n3 B 0.591606f
C44 VTAIL.t4 B 0.39181f
C45 VTAIL.n4 B 0.224774f
C46 VTAIL.t0 B 0.39181f
C47 VTAIL.n5 B 0.224774f
C48 VTAIL.t1 B 0.391808f
C49 VTAIL.n6 B 0.591608f
C50 VTAIL.t5 B 0.391808f
C51 VTAIL.n7 B 0.55848f
C52 VDD2.t1 B 0.059326f
C53 VDD2.t3 B 0.059326f
C54 VDD2.n0 B 0.692941f
C55 VDD2.t0 B 0.059326f
C56 VDD2.t2 B 0.059326f
C57 VDD2.n1 B 0.469785f
C58 VDD2.n2 B 1.71036f
C59 VN.t1 B 0.400002f
C60 VN.t2 B 0.39954f
C61 VN.n0 B 0.313601f
C62 VN.t3 B 0.400002f
C63 VN.t0 B 0.39954f
C64 VN.n1 B 0.873828f
.ends

