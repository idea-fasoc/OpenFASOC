* NGSPICE file created from diff_pair_sample_0854.ext - technology: sky130A

.subckt diff_pair_sample_0854 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t5 w_n2800_n4698# sky130_fd_pr__pfet_01v8 ad=7.2735 pd=38.08 as=3.07725 ps=18.98 w=18.65 l=1.5
X1 B.t11 B.t9 B.t10 w_n2800_n4698# sky130_fd_pr__pfet_01v8 ad=7.2735 pd=38.08 as=0 ps=0 w=18.65 l=1.5
X2 VDD1.t4 VP.t1 VTAIL.t14 w_n2800_n4698# sky130_fd_pr__pfet_01v8 ad=3.07725 pd=18.98 as=3.07725 ps=18.98 w=18.65 l=1.5
X3 VTAIL.t4 VN.t0 VDD2.t7 w_n2800_n4698# sky130_fd_pr__pfet_01v8 ad=3.07725 pd=18.98 as=3.07725 ps=18.98 w=18.65 l=1.5
X4 VTAIL.t13 VP.t2 VDD1.t3 w_n2800_n4698# sky130_fd_pr__pfet_01v8 ad=7.2735 pd=38.08 as=3.07725 ps=18.98 w=18.65 l=1.5
X5 VDD2.t6 VN.t1 VTAIL.t3 w_n2800_n4698# sky130_fd_pr__pfet_01v8 ad=3.07725 pd=18.98 as=7.2735 ps=38.08 w=18.65 l=1.5
X6 VDD2.t5 VN.t2 VTAIL.t6 w_n2800_n4698# sky130_fd_pr__pfet_01v8 ad=3.07725 pd=18.98 as=3.07725 ps=18.98 w=18.65 l=1.5
X7 VTAIL.t12 VP.t3 VDD1.t2 w_n2800_n4698# sky130_fd_pr__pfet_01v8 ad=3.07725 pd=18.98 as=3.07725 ps=18.98 w=18.65 l=1.5
X8 VDD2.t4 VN.t3 VTAIL.t7 w_n2800_n4698# sky130_fd_pr__pfet_01v8 ad=3.07725 pd=18.98 as=7.2735 ps=38.08 w=18.65 l=1.5
X9 VTAIL.t2 VN.t4 VDD2.t3 w_n2800_n4698# sky130_fd_pr__pfet_01v8 ad=7.2735 pd=38.08 as=3.07725 ps=18.98 w=18.65 l=1.5
X10 VDD1.t7 VP.t4 VTAIL.t11 w_n2800_n4698# sky130_fd_pr__pfet_01v8 ad=3.07725 pd=18.98 as=7.2735 ps=38.08 w=18.65 l=1.5
X11 VTAIL.t1 VN.t5 VDD2.t2 w_n2800_n4698# sky130_fd_pr__pfet_01v8 ad=3.07725 pd=18.98 as=3.07725 ps=18.98 w=18.65 l=1.5
X12 VDD1.t6 VP.t5 VTAIL.t10 w_n2800_n4698# sky130_fd_pr__pfet_01v8 ad=3.07725 pd=18.98 as=3.07725 ps=18.98 w=18.65 l=1.5
X13 VDD1.t1 VP.t6 VTAIL.t9 w_n2800_n4698# sky130_fd_pr__pfet_01v8 ad=3.07725 pd=18.98 as=7.2735 ps=38.08 w=18.65 l=1.5
X14 B.t8 B.t6 B.t7 w_n2800_n4698# sky130_fd_pr__pfet_01v8 ad=7.2735 pd=38.08 as=0 ps=0 w=18.65 l=1.5
X15 B.t5 B.t3 B.t4 w_n2800_n4698# sky130_fd_pr__pfet_01v8 ad=7.2735 pd=38.08 as=0 ps=0 w=18.65 l=1.5
X16 VTAIL.t8 VP.t7 VDD1.t0 w_n2800_n4698# sky130_fd_pr__pfet_01v8 ad=3.07725 pd=18.98 as=3.07725 ps=18.98 w=18.65 l=1.5
X17 VTAIL.t5 VN.t6 VDD2.t1 w_n2800_n4698# sky130_fd_pr__pfet_01v8 ad=7.2735 pd=38.08 as=3.07725 ps=18.98 w=18.65 l=1.5
X18 B.t2 B.t0 B.t1 w_n2800_n4698# sky130_fd_pr__pfet_01v8 ad=7.2735 pd=38.08 as=0 ps=0 w=18.65 l=1.5
X19 VDD2.t0 VN.t7 VTAIL.t0 w_n2800_n4698# sky130_fd_pr__pfet_01v8 ad=3.07725 pd=18.98 as=3.07725 ps=18.98 w=18.65 l=1.5
R0 VP.n11 VP.t2 334.392
R1 VP.n25 VP.t0 299.644
R2 VP.n31 VP.t5 299.644
R3 VP.n38 VP.t3 299.644
R4 VP.n45 VP.t4 299.644
R5 VP.n23 VP.t6 299.644
R6 VP.n16 VP.t7 299.644
R7 VP.n10 VP.t1 299.644
R8 VP.n26 VP.n25 173.779
R9 VP.n46 VP.n45 173.779
R10 VP.n24 VP.n23 173.779
R11 VP.n12 VP.n9 161.3
R12 VP.n14 VP.n13 161.3
R13 VP.n15 VP.n8 161.3
R14 VP.n18 VP.n17 161.3
R15 VP.n19 VP.n7 161.3
R16 VP.n21 VP.n20 161.3
R17 VP.n22 VP.n6 161.3
R18 VP.n44 VP.n0 161.3
R19 VP.n43 VP.n42 161.3
R20 VP.n41 VP.n1 161.3
R21 VP.n40 VP.n39 161.3
R22 VP.n37 VP.n2 161.3
R23 VP.n36 VP.n35 161.3
R24 VP.n34 VP.n3 161.3
R25 VP.n33 VP.n32 161.3
R26 VP.n30 VP.n4 161.3
R27 VP.n29 VP.n28 161.3
R28 VP.n27 VP.n5 161.3
R29 VP.n30 VP.n29 56.5193
R30 VP.n43 VP.n1 56.5193
R31 VP.n21 VP.n7 56.5193
R32 VP.n26 VP.n24 50.7429
R33 VP.n11 VP.n10 46.2606
R34 VP.n36 VP.n3 40.4934
R35 VP.n37 VP.n36 40.4934
R36 VP.n15 VP.n14 40.4934
R37 VP.n14 VP.n9 40.4934
R38 VP.n29 VP.n5 24.4675
R39 VP.n32 VP.n30 24.4675
R40 VP.n39 VP.n1 24.4675
R41 VP.n44 VP.n43 24.4675
R42 VP.n22 VP.n21 24.4675
R43 VP.n17 VP.n7 24.4675
R44 VP.n31 VP.n3 20.3081
R45 VP.n38 VP.n37 20.3081
R46 VP.n16 VP.n15 20.3081
R47 VP.n10 VP.n9 20.3081
R48 VP.n12 VP.n11 17.5886
R49 VP.n25 VP.n5 11.9893
R50 VP.n45 VP.n44 11.9893
R51 VP.n23 VP.n22 11.9893
R52 VP.n32 VP.n31 4.15989
R53 VP.n39 VP.n38 4.15989
R54 VP.n17 VP.n16 4.15989
R55 VP.n13 VP.n12 0.189894
R56 VP.n13 VP.n8 0.189894
R57 VP.n18 VP.n8 0.189894
R58 VP.n19 VP.n18 0.189894
R59 VP.n20 VP.n19 0.189894
R60 VP.n20 VP.n6 0.189894
R61 VP.n24 VP.n6 0.189894
R62 VP.n27 VP.n26 0.189894
R63 VP.n28 VP.n27 0.189894
R64 VP.n28 VP.n4 0.189894
R65 VP.n33 VP.n4 0.189894
R66 VP.n34 VP.n33 0.189894
R67 VP.n35 VP.n34 0.189894
R68 VP.n35 VP.n2 0.189894
R69 VP.n40 VP.n2 0.189894
R70 VP.n41 VP.n40 0.189894
R71 VP.n42 VP.n41 0.189894
R72 VP.n42 VP.n0 0.189894
R73 VP.n46 VP.n0 0.189894
R74 VP VP.n46 0.0516364
R75 VDD1 VDD1.n0 70.3492
R76 VDD1.n3 VDD1.n2 70.2354
R77 VDD1.n3 VDD1.n1 70.2354
R78 VDD1.n5 VDD1.n4 69.502
R79 VDD1.n5 VDD1.n3 47.475
R80 VDD1.n4 VDD1.t0 1.7434
R81 VDD1.n4 VDD1.t1 1.7434
R82 VDD1.n0 VDD1.t3 1.7434
R83 VDD1.n0 VDD1.t4 1.7434
R84 VDD1.n2 VDD1.t2 1.7434
R85 VDD1.n2 VDD1.t7 1.7434
R86 VDD1.n1 VDD1.t5 1.7434
R87 VDD1.n1 VDD1.t6 1.7434
R88 VDD1 VDD1.n5 0.731103
R89 VTAIL.n11 VTAIL.t13 54.5663
R90 VTAIL.n10 VTAIL.t3 54.5663
R91 VTAIL.n7 VTAIL.t5 54.5663
R92 VTAIL.n14 VTAIL.t9 54.5661
R93 VTAIL.n15 VTAIL.t7 54.5661
R94 VTAIL.n2 VTAIL.t2 54.5661
R95 VTAIL.n3 VTAIL.t11 54.5661
R96 VTAIL.n6 VTAIL.t15 54.5661
R97 VTAIL.n13 VTAIL.n12 52.8234
R98 VTAIL.n9 VTAIL.n8 52.8234
R99 VTAIL.n1 VTAIL.n0 52.8232
R100 VTAIL.n5 VTAIL.n4 52.8232
R101 VTAIL.n15 VTAIL.n14 30.0221
R102 VTAIL.n7 VTAIL.n6 30.0221
R103 VTAIL.n0 VTAIL.t6 1.7434
R104 VTAIL.n0 VTAIL.t1 1.7434
R105 VTAIL.n4 VTAIL.t10 1.7434
R106 VTAIL.n4 VTAIL.t12 1.7434
R107 VTAIL.n12 VTAIL.t14 1.7434
R108 VTAIL.n12 VTAIL.t8 1.7434
R109 VTAIL.n8 VTAIL.t0 1.7434
R110 VTAIL.n8 VTAIL.t4 1.7434
R111 VTAIL.n9 VTAIL.n7 1.57809
R112 VTAIL.n10 VTAIL.n9 1.57809
R113 VTAIL.n13 VTAIL.n11 1.57809
R114 VTAIL.n14 VTAIL.n13 1.57809
R115 VTAIL.n6 VTAIL.n5 1.57809
R116 VTAIL.n5 VTAIL.n3 1.57809
R117 VTAIL.n2 VTAIL.n1 1.57809
R118 VTAIL VTAIL.n15 1.5199
R119 VTAIL.n11 VTAIL.n10 0.470328
R120 VTAIL.n3 VTAIL.n2 0.470328
R121 VTAIL VTAIL.n1 0.0586897
R122 B.n571 B.n570 585
R123 B.n572 B.n89 585
R124 B.n574 B.n573 585
R125 B.n575 B.n88 585
R126 B.n577 B.n576 585
R127 B.n578 B.n87 585
R128 B.n580 B.n579 585
R129 B.n581 B.n86 585
R130 B.n583 B.n582 585
R131 B.n584 B.n85 585
R132 B.n586 B.n585 585
R133 B.n587 B.n84 585
R134 B.n589 B.n588 585
R135 B.n590 B.n83 585
R136 B.n592 B.n591 585
R137 B.n593 B.n82 585
R138 B.n595 B.n594 585
R139 B.n596 B.n81 585
R140 B.n598 B.n597 585
R141 B.n599 B.n80 585
R142 B.n601 B.n600 585
R143 B.n602 B.n79 585
R144 B.n604 B.n603 585
R145 B.n605 B.n78 585
R146 B.n607 B.n606 585
R147 B.n608 B.n77 585
R148 B.n610 B.n609 585
R149 B.n611 B.n76 585
R150 B.n613 B.n612 585
R151 B.n614 B.n75 585
R152 B.n616 B.n615 585
R153 B.n617 B.n74 585
R154 B.n619 B.n618 585
R155 B.n620 B.n73 585
R156 B.n622 B.n621 585
R157 B.n623 B.n72 585
R158 B.n625 B.n624 585
R159 B.n626 B.n71 585
R160 B.n628 B.n627 585
R161 B.n629 B.n70 585
R162 B.n631 B.n630 585
R163 B.n632 B.n69 585
R164 B.n634 B.n633 585
R165 B.n635 B.n68 585
R166 B.n637 B.n636 585
R167 B.n638 B.n67 585
R168 B.n640 B.n639 585
R169 B.n641 B.n66 585
R170 B.n643 B.n642 585
R171 B.n644 B.n65 585
R172 B.n646 B.n645 585
R173 B.n647 B.n64 585
R174 B.n649 B.n648 585
R175 B.n650 B.n63 585
R176 B.n652 B.n651 585
R177 B.n653 B.n62 585
R178 B.n655 B.n654 585
R179 B.n656 B.n61 585
R180 B.n658 B.n657 585
R181 B.n659 B.n60 585
R182 B.n661 B.n660 585
R183 B.n663 B.n57 585
R184 B.n665 B.n664 585
R185 B.n666 B.n56 585
R186 B.n668 B.n667 585
R187 B.n669 B.n55 585
R188 B.n671 B.n670 585
R189 B.n672 B.n54 585
R190 B.n674 B.n673 585
R191 B.n675 B.n53 585
R192 B.n677 B.n676 585
R193 B.n679 B.n678 585
R194 B.n680 B.n49 585
R195 B.n682 B.n681 585
R196 B.n683 B.n48 585
R197 B.n685 B.n684 585
R198 B.n686 B.n47 585
R199 B.n688 B.n687 585
R200 B.n689 B.n46 585
R201 B.n691 B.n690 585
R202 B.n692 B.n45 585
R203 B.n694 B.n693 585
R204 B.n695 B.n44 585
R205 B.n697 B.n696 585
R206 B.n698 B.n43 585
R207 B.n700 B.n699 585
R208 B.n701 B.n42 585
R209 B.n703 B.n702 585
R210 B.n704 B.n41 585
R211 B.n706 B.n705 585
R212 B.n707 B.n40 585
R213 B.n709 B.n708 585
R214 B.n710 B.n39 585
R215 B.n712 B.n711 585
R216 B.n713 B.n38 585
R217 B.n715 B.n714 585
R218 B.n716 B.n37 585
R219 B.n718 B.n717 585
R220 B.n719 B.n36 585
R221 B.n721 B.n720 585
R222 B.n722 B.n35 585
R223 B.n724 B.n723 585
R224 B.n725 B.n34 585
R225 B.n727 B.n726 585
R226 B.n728 B.n33 585
R227 B.n730 B.n729 585
R228 B.n731 B.n32 585
R229 B.n733 B.n732 585
R230 B.n734 B.n31 585
R231 B.n736 B.n735 585
R232 B.n737 B.n30 585
R233 B.n739 B.n738 585
R234 B.n740 B.n29 585
R235 B.n742 B.n741 585
R236 B.n743 B.n28 585
R237 B.n745 B.n744 585
R238 B.n746 B.n27 585
R239 B.n748 B.n747 585
R240 B.n749 B.n26 585
R241 B.n751 B.n750 585
R242 B.n752 B.n25 585
R243 B.n754 B.n753 585
R244 B.n755 B.n24 585
R245 B.n757 B.n756 585
R246 B.n758 B.n23 585
R247 B.n760 B.n759 585
R248 B.n761 B.n22 585
R249 B.n763 B.n762 585
R250 B.n764 B.n21 585
R251 B.n766 B.n765 585
R252 B.n767 B.n20 585
R253 B.n769 B.n768 585
R254 B.n569 B.n90 585
R255 B.n568 B.n567 585
R256 B.n566 B.n91 585
R257 B.n565 B.n564 585
R258 B.n563 B.n92 585
R259 B.n562 B.n561 585
R260 B.n560 B.n93 585
R261 B.n559 B.n558 585
R262 B.n557 B.n94 585
R263 B.n556 B.n555 585
R264 B.n554 B.n95 585
R265 B.n553 B.n552 585
R266 B.n551 B.n96 585
R267 B.n550 B.n549 585
R268 B.n548 B.n97 585
R269 B.n547 B.n546 585
R270 B.n545 B.n98 585
R271 B.n544 B.n543 585
R272 B.n542 B.n99 585
R273 B.n541 B.n540 585
R274 B.n539 B.n100 585
R275 B.n538 B.n537 585
R276 B.n536 B.n101 585
R277 B.n535 B.n534 585
R278 B.n533 B.n102 585
R279 B.n532 B.n531 585
R280 B.n530 B.n103 585
R281 B.n529 B.n528 585
R282 B.n527 B.n104 585
R283 B.n526 B.n525 585
R284 B.n524 B.n105 585
R285 B.n523 B.n522 585
R286 B.n521 B.n106 585
R287 B.n520 B.n519 585
R288 B.n518 B.n107 585
R289 B.n517 B.n516 585
R290 B.n515 B.n108 585
R291 B.n514 B.n513 585
R292 B.n512 B.n109 585
R293 B.n511 B.n510 585
R294 B.n509 B.n110 585
R295 B.n508 B.n507 585
R296 B.n506 B.n111 585
R297 B.n505 B.n504 585
R298 B.n503 B.n112 585
R299 B.n502 B.n501 585
R300 B.n500 B.n113 585
R301 B.n499 B.n498 585
R302 B.n497 B.n114 585
R303 B.n496 B.n495 585
R304 B.n494 B.n115 585
R305 B.n493 B.n492 585
R306 B.n491 B.n116 585
R307 B.n490 B.n489 585
R308 B.n488 B.n117 585
R309 B.n487 B.n486 585
R310 B.n485 B.n118 585
R311 B.n484 B.n483 585
R312 B.n482 B.n119 585
R313 B.n481 B.n480 585
R314 B.n479 B.n120 585
R315 B.n478 B.n477 585
R316 B.n476 B.n121 585
R317 B.n475 B.n474 585
R318 B.n473 B.n122 585
R319 B.n472 B.n471 585
R320 B.n470 B.n123 585
R321 B.n469 B.n468 585
R322 B.n467 B.n124 585
R323 B.n466 B.n465 585
R324 B.n464 B.n125 585
R325 B.n265 B.n264 585
R326 B.n266 B.n195 585
R327 B.n268 B.n267 585
R328 B.n269 B.n194 585
R329 B.n271 B.n270 585
R330 B.n272 B.n193 585
R331 B.n274 B.n273 585
R332 B.n275 B.n192 585
R333 B.n277 B.n276 585
R334 B.n278 B.n191 585
R335 B.n280 B.n279 585
R336 B.n281 B.n190 585
R337 B.n283 B.n282 585
R338 B.n284 B.n189 585
R339 B.n286 B.n285 585
R340 B.n287 B.n188 585
R341 B.n289 B.n288 585
R342 B.n290 B.n187 585
R343 B.n292 B.n291 585
R344 B.n293 B.n186 585
R345 B.n295 B.n294 585
R346 B.n296 B.n185 585
R347 B.n298 B.n297 585
R348 B.n299 B.n184 585
R349 B.n301 B.n300 585
R350 B.n302 B.n183 585
R351 B.n304 B.n303 585
R352 B.n305 B.n182 585
R353 B.n307 B.n306 585
R354 B.n308 B.n181 585
R355 B.n310 B.n309 585
R356 B.n311 B.n180 585
R357 B.n313 B.n312 585
R358 B.n314 B.n179 585
R359 B.n316 B.n315 585
R360 B.n317 B.n178 585
R361 B.n319 B.n318 585
R362 B.n320 B.n177 585
R363 B.n322 B.n321 585
R364 B.n323 B.n176 585
R365 B.n325 B.n324 585
R366 B.n326 B.n175 585
R367 B.n328 B.n327 585
R368 B.n329 B.n174 585
R369 B.n331 B.n330 585
R370 B.n332 B.n173 585
R371 B.n334 B.n333 585
R372 B.n335 B.n172 585
R373 B.n337 B.n336 585
R374 B.n338 B.n171 585
R375 B.n340 B.n339 585
R376 B.n341 B.n170 585
R377 B.n343 B.n342 585
R378 B.n344 B.n169 585
R379 B.n346 B.n345 585
R380 B.n347 B.n168 585
R381 B.n349 B.n348 585
R382 B.n350 B.n167 585
R383 B.n352 B.n351 585
R384 B.n353 B.n166 585
R385 B.n355 B.n354 585
R386 B.n357 B.n163 585
R387 B.n359 B.n358 585
R388 B.n360 B.n162 585
R389 B.n362 B.n361 585
R390 B.n363 B.n161 585
R391 B.n365 B.n364 585
R392 B.n366 B.n160 585
R393 B.n368 B.n367 585
R394 B.n369 B.n159 585
R395 B.n371 B.n370 585
R396 B.n373 B.n372 585
R397 B.n374 B.n155 585
R398 B.n376 B.n375 585
R399 B.n377 B.n154 585
R400 B.n379 B.n378 585
R401 B.n380 B.n153 585
R402 B.n382 B.n381 585
R403 B.n383 B.n152 585
R404 B.n385 B.n384 585
R405 B.n386 B.n151 585
R406 B.n388 B.n387 585
R407 B.n389 B.n150 585
R408 B.n391 B.n390 585
R409 B.n392 B.n149 585
R410 B.n394 B.n393 585
R411 B.n395 B.n148 585
R412 B.n397 B.n396 585
R413 B.n398 B.n147 585
R414 B.n400 B.n399 585
R415 B.n401 B.n146 585
R416 B.n403 B.n402 585
R417 B.n404 B.n145 585
R418 B.n406 B.n405 585
R419 B.n407 B.n144 585
R420 B.n409 B.n408 585
R421 B.n410 B.n143 585
R422 B.n412 B.n411 585
R423 B.n413 B.n142 585
R424 B.n415 B.n414 585
R425 B.n416 B.n141 585
R426 B.n418 B.n417 585
R427 B.n419 B.n140 585
R428 B.n421 B.n420 585
R429 B.n422 B.n139 585
R430 B.n424 B.n423 585
R431 B.n425 B.n138 585
R432 B.n427 B.n426 585
R433 B.n428 B.n137 585
R434 B.n430 B.n429 585
R435 B.n431 B.n136 585
R436 B.n433 B.n432 585
R437 B.n434 B.n135 585
R438 B.n436 B.n435 585
R439 B.n437 B.n134 585
R440 B.n439 B.n438 585
R441 B.n440 B.n133 585
R442 B.n442 B.n441 585
R443 B.n443 B.n132 585
R444 B.n445 B.n444 585
R445 B.n446 B.n131 585
R446 B.n448 B.n447 585
R447 B.n449 B.n130 585
R448 B.n451 B.n450 585
R449 B.n452 B.n129 585
R450 B.n454 B.n453 585
R451 B.n455 B.n128 585
R452 B.n457 B.n456 585
R453 B.n458 B.n127 585
R454 B.n460 B.n459 585
R455 B.n461 B.n126 585
R456 B.n463 B.n462 585
R457 B.n263 B.n196 585
R458 B.n262 B.n261 585
R459 B.n260 B.n197 585
R460 B.n259 B.n258 585
R461 B.n257 B.n198 585
R462 B.n256 B.n255 585
R463 B.n254 B.n199 585
R464 B.n253 B.n252 585
R465 B.n251 B.n200 585
R466 B.n250 B.n249 585
R467 B.n248 B.n201 585
R468 B.n247 B.n246 585
R469 B.n245 B.n202 585
R470 B.n244 B.n243 585
R471 B.n242 B.n203 585
R472 B.n241 B.n240 585
R473 B.n239 B.n204 585
R474 B.n238 B.n237 585
R475 B.n236 B.n205 585
R476 B.n235 B.n234 585
R477 B.n233 B.n206 585
R478 B.n232 B.n231 585
R479 B.n230 B.n207 585
R480 B.n229 B.n228 585
R481 B.n227 B.n208 585
R482 B.n226 B.n225 585
R483 B.n224 B.n209 585
R484 B.n223 B.n222 585
R485 B.n221 B.n210 585
R486 B.n220 B.n219 585
R487 B.n218 B.n211 585
R488 B.n217 B.n216 585
R489 B.n215 B.n212 585
R490 B.n214 B.n213 585
R491 B.n2 B.n0 585
R492 B.n821 B.n1 585
R493 B.n820 B.n819 585
R494 B.n818 B.n3 585
R495 B.n817 B.n816 585
R496 B.n815 B.n4 585
R497 B.n814 B.n813 585
R498 B.n812 B.n5 585
R499 B.n811 B.n810 585
R500 B.n809 B.n6 585
R501 B.n808 B.n807 585
R502 B.n806 B.n7 585
R503 B.n805 B.n804 585
R504 B.n803 B.n8 585
R505 B.n802 B.n801 585
R506 B.n800 B.n9 585
R507 B.n799 B.n798 585
R508 B.n797 B.n10 585
R509 B.n796 B.n795 585
R510 B.n794 B.n11 585
R511 B.n793 B.n792 585
R512 B.n791 B.n12 585
R513 B.n790 B.n789 585
R514 B.n788 B.n13 585
R515 B.n787 B.n786 585
R516 B.n785 B.n14 585
R517 B.n784 B.n783 585
R518 B.n782 B.n15 585
R519 B.n781 B.n780 585
R520 B.n779 B.n16 585
R521 B.n778 B.n777 585
R522 B.n776 B.n17 585
R523 B.n775 B.n774 585
R524 B.n773 B.n18 585
R525 B.n772 B.n771 585
R526 B.n770 B.n19 585
R527 B.n823 B.n822 585
R528 B.n156 B.t6 505.084
R529 B.n164 B.t9 505.084
R530 B.n50 B.t0 505.084
R531 B.n58 B.t3 505.084
R532 B.n264 B.n263 497.305
R533 B.n768 B.n19 497.305
R534 B.n462 B.n125 497.305
R535 B.n570 B.n569 497.305
R536 B.n263 B.n262 163.367
R537 B.n262 B.n197 163.367
R538 B.n258 B.n197 163.367
R539 B.n258 B.n257 163.367
R540 B.n257 B.n256 163.367
R541 B.n256 B.n199 163.367
R542 B.n252 B.n199 163.367
R543 B.n252 B.n251 163.367
R544 B.n251 B.n250 163.367
R545 B.n250 B.n201 163.367
R546 B.n246 B.n201 163.367
R547 B.n246 B.n245 163.367
R548 B.n245 B.n244 163.367
R549 B.n244 B.n203 163.367
R550 B.n240 B.n203 163.367
R551 B.n240 B.n239 163.367
R552 B.n239 B.n238 163.367
R553 B.n238 B.n205 163.367
R554 B.n234 B.n205 163.367
R555 B.n234 B.n233 163.367
R556 B.n233 B.n232 163.367
R557 B.n232 B.n207 163.367
R558 B.n228 B.n207 163.367
R559 B.n228 B.n227 163.367
R560 B.n227 B.n226 163.367
R561 B.n226 B.n209 163.367
R562 B.n222 B.n209 163.367
R563 B.n222 B.n221 163.367
R564 B.n221 B.n220 163.367
R565 B.n220 B.n211 163.367
R566 B.n216 B.n211 163.367
R567 B.n216 B.n215 163.367
R568 B.n215 B.n214 163.367
R569 B.n214 B.n2 163.367
R570 B.n822 B.n2 163.367
R571 B.n822 B.n821 163.367
R572 B.n821 B.n820 163.367
R573 B.n820 B.n3 163.367
R574 B.n816 B.n3 163.367
R575 B.n816 B.n815 163.367
R576 B.n815 B.n814 163.367
R577 B.n814 B.n5 163.367
R578 B.n810 B.n5 163.367
R579 B.n810 B.n809 163.367
R580 B.n809 B.n808 163.367
R581 B.n808 B.n7 163.367
R582 B.n804 B.n7 163.367
R583 B.n804 B.n803 163.367
R584 B.n803 B.n802 163.367
R585 B.n802 B.n9 163.367
R586 B.n798 B.n9 163.367
R587 B.n798 B.n797 163.367
R588 B.n797 B.n796 163.367
R589 B.n796 B.n11 163.367
R590 B.n792 B.n11 163.367
R591 B.n792 B.n791 163.367
R592 B.n791 B.n790 163.367
R593 B.n790 B.n13 163.367
R594 B.n786 B.n13 163.367
R595 B.n786 B.n785 163.367
R596 B.n785 B.n784 163.367
R597 B.n784 B.n15 163.367
R598 B.n780 B.n15 163.367
R599 B.n780 B.n779 163.367
R600 B.n779 B.n778 163.367
R601 B.n778 B.n17 163.367
R602 B.n774 B.n17 163.367
R603 B.n774 B.n773 163.367
R604 B.n773 B.n772 163.367
R605 B.n772 B.n19 163.367
R606 B.n264 B.n195 163.367
R607 B.n268 B.n195 163.367
R608 B.n269 B.n268 163.367
R609 B.n270 B.n269 163.367
R610 B.n270 B.n193 163.367
R611 B.n274 B.n193 163.367
R612 B.n275 B.n274 163.367
R613 B.n276 B.n275 163.367
R614 B.n276 B.n191 163.367
R615 B.n280 B.n191 163.367
R616 B.n281 B.n280 163.367
R617 B.n282 B.n281 163.367
R618 B.n282 B.n189 163.367
R619 B.n286 B.n189 163.367
R620 B.n287 B.n286 163.367
R621 B.n288 B.n287 163.367
R622 B.n288 B.n187 163.367
R623 B.n292 B.n187 163.367
R624 B.n293 B.n292 163.367
R625 B.n294 B.n293 163.367
R626 B.n294 B.n185 163.367
R627 B.n298 B.n185 163.367
R628 B.n299 B.n298 163.367
R629 B.n300 B.n299 163.367
R630 B.n300 B.n183 163.367
R631 B.n304 B.n183 163.367
R632 B.n305 B.n304 163.367
R633 B.n306 B.n305 163.367
R634 B.n306 B.n181 163.367
R635 B.n310 B.n181 163.367
R636 B.n311 B.n310 163.367
R637 B.n312 B.n311 163.367
R638 B.n312 B.n179 163.367
R639 B.n316 B.n179 163.367
R640 B.n317 B.n316 163.367
R641 B.n318 B.n317 163.367
R642 B.n318 B.n177 163.367
R643 B.n322 B.n177 163.367
R644 B.n323 B.n322 163.367
R645 B.n324 B.n323 163.367
R646 B.n324 B.n175 163.367
R647 B.n328 B.n175 163.367
R648 B.n329 B.n328 163.367
R649 B.n330 B.n329 163.367
R650 B.n330 B.n173 163.367
R651 B.n334 B.n173 163.367
R652 B.n335 B.n334 163.367
R653 B.n336 B.n335 163.367
R654 B.n336 B.n171 163.367
R655 B.n340 B.n171 163.367
R656 B.n341 B.n340 163.367
R657 B.n342 B.n341 163.367
R658 B.n342 B.n169 163.367
R659 B.n346 B.n169 163.367
R660 B.n347 B.n346 163.367
R661 B.n348 B.n347 163.367
R662 B.n348 B.n167 163.367
R663 B.n352 B.n167 163.367
R664 B.n353 B.n352 163.367
R665 B.n354 B.n353 163.367
R666 B.n354 B.n163 163.367
R667 B.n359 B.n163 163.367
R668 B.n360 B.n359 163.367
R669 B.n361 B.n360 163.367
R670 B.n361 B.n161 163.367
R671 B.n365 B.n161 163.367
R672 B.n366 B.n365 163.367
R673 B.n367 B.n366 163.367
R674 B.n367 B.n159 163.367
R675 B.n371 B.n159 163.367
R676 B.n372 B.n371 163.367
R677 B.n372 B.n155 163.367
R678 B.n376 B.n155 163.367
R679 B.n377 B.n376 163.367
R680 B.n378 B.n377 163.367
R681 B.n378 B.n153 163.367
R682 B.n382 B.n153 163.367
R683 B.n383 B.n382 163.367
R684 B.n384 B.n383 163.367
R685 B.n384 B.n151 163.367
R686 B.n388 B.n151 163.367
R687 B.n389 B.n388 163.367
R688 B.n390 B.n389 163.367
R689 B.n390 B.n149 163.367
R690 B.n394 B.n149 163.367
R691 B.n395 B.n394 163.367
R692 B.n396 B.n395 163.367
R693 B.n396 B.n147 163.367
R694 B.n400 B.n147 163.367
R695 B.n401 B.n400 163.367
R696 B.n402 B.n401 163.367
R697 B.n402 B.n145 163.367
R698 B.n406 B.n145 163.367
R699 B.n407 B.n406 163.367
R700 B.n408 B.n407 163.367
R701 B.n408 B.n143 163.367
R702 B.n412 B.n143 163.367
R703 B.n413 B.n412 163.367
R704 B.n414 B.n413 163.367
R705 B.n414 B.n141 163.367
R706 B.n418 B.n141 163.367
R707 B.n419 B.n418 163.367
R708 B.n420 B.n419 163.367
R709 B.n420 B.n139 163.367
R710 B.n424 B.n139 163.367
R711 B.n425 B.n424 163.367
R712 B.n426 B.n425 163.367
R713 B.n426 B.n137 163.367
R714 B.n430 B.n137 163.367
R715 B.n431 B.n430 163.367
R716 B.n432 B.n431 163.367
R717 B.n432 B.n135 163.367
R718 B.n436 B.n135 163.367
R719 B.n437 B.n436 163.367
R720 B.n438 B.n437 163.367
R721 B.n438 B.n133 163.367
R722 B.n442 B.n133 163.367
R723 B.n443 B.n442 163.367
R724 B.n444 B.n443 163.367
R725 B.n444 B.n131 163.367
R726 B.n448 B.n131 163.367
R727 B.n449 B.n448 163.367
R728 B.n450 B.n449 163.367
R729 B.n450 B.n129 163.367
R730 B.n454 B.n129 163.367
R731 B.n455 B.n454 163.367
R732 B.n456 B.n455 163.367
R733 B.n456 B.n127 163.367
R734 B.n460 B.n127 163.367
R735 B.n461 B.n460 163.367
R736 B.n462 B.n461 163.367
R737 B.n466 B.n125 163.367
R738 B.n467 B.n466 163.367
R739 B.n468 B.n467 163.367
R740 B.n468 B.n123 163.367
R741 B.n472 B.n123 163.367
R742 B.n473 B.n472 163.367
R743 B.n474 B.n473 163.367
R744 B.n474 B.n121 163.367
R745 B.n478 B.n121 163.367
R746 B.n479 B.n478 163.367
R747 B.n480 B.n479 163.367
R748 B.n480 B.n119 163.367
R749 B.n484 B.n119 163.367
R750 B.n485 B.n484 163.367
R751 B.n486 B.n485 163.367
R752 B.n486 B.n117 163.367
R753 B.n490 B.n117 163.367
R754 B.n491 B.n490 163.367
R755 B.n492 B.n491 163.367
R756 B.n492 B.n115 163.367
R757 B.n496 B.n115 163.367
R758 B.n497 B.n496 163.367
R759 B.n498 B.n497 163.367
R760 B.n498 B.n113 163.367
R761 B.n502 B.n113 163.367
R762 B.n503 B.n502 163.367
R763 B.n504 B.n503 163.367
R764 B.n504 B.n111 163.367
R765 B.n508 B.n111 163.367
R766 B.n509 B.n508 163.367
R767 B.n510 B.n509 163.367
R768 B.n510 B.n109 163.367
R769 B.n514 B.n109 163.367
R770 B.n515 B.n514 163.367
R771 B.n516 B.n515 163.367
R772 B.n516 B.n107 163.367
R773 B.n520 B.n107 163.367
R774 B.n521 B.n520 163.367
R775 B.n522 B.n521 163.367
R776 B.n522 B.n105 163.367
R777 B.n526 B.n105 163.367
R778 B.n527 B.n526 163.367
R779 B.n528 B.n527 163.367
R780 B.n528 B.n103 163.367
R781 B.n532 B.n103 163.367
R782 B.n533 B.n532 163.367
R783 B.n534 B.n533 163.367
R784 B.n534 B.n101 163.367
R785 B.n538 B.n101 163.367
R786 B.n539 B.n538 163.367
R787 B.n540 B.n539 163.367
R788 B.n540 B.n99 163.367
R789 B.n544 B.n99 163.367
R790 B.n545 B.n544 163.367
R791 B.n546 B.n545 163.367
R792 B.n546 B.n97 163.367
R793 B.n550 B.n97 163.367
R794 B.n551 B.n550 163.367
R795 B.n552 B.n551 163.367
R796 B.n552 B.n95 163.367
R797 B.n556 B.n95 163.367
R798 B.n557 B.n556 163.367
R799 B.n558 B.n557 163.367
R800 B.n558 B.n93 163.367
R801 B.n562 B.n93 163.367
R802 B.n563 B.n562 163.367
R803 B.n564 B.n563 163.367
R804 B.n564 B.n91 163.367
R805 B.n568 B.n91 163.367
R806 B.n569 B.n568 163.367
R807 B.n768 B.n767 163.367
R808 B.n767 B.n766 163.367
R809 B.n766 B.n21 163.367
R810 B.n762 B.n21 163.367
R811 B.n762 B.n761 163.367
R812 B.n761 B.n760 163.367
R813 B.n760 B.n23 163.367
R814 B.n756 B.n23 163.367
R815 B.n756 B.n755 163.367
R816 B.n755 B.n754 163.367
R817 B.n754 B.n25 163.367
R818 B.n750 B.n25 163.367
R819 B.n750 B.n749 163.367
R820 B.n749 B.n748 163.367
R821 B.n748 B.n27 163.367
R822 B.n744 B.n27 163.367
R823 B.n744 B.n743 163.367
R824 B.n743 B.n742 163.367
R825 B.n742 B.n29 163.367
R826 B.n738 B.n29 163.367
R827 B.n738 B.n737 163.367
R828 B.n737 B.n736 163.367
R829 B.n736 B.n31 163.367
R830 B.n732 B.n31 163.367
R831 B.n732 B.n731 163.367
R832 B.n731 B.n730 163.367
R833 B.n730 B.n33 163.367
R834 B.n726 B.n33 163.367
R835 B.n726 B.n725 163.367
R836 B.n725 B.n724 163.367
R837 B.n724 B.n35 163.367
R838 B.n720 B.n35 163.367
R839 B.n720 B.n719 163.367
R840 B.n719 B.n718 163.367
R841 B.n718 B.n37 163.367
R842 B.n714 B.n37 163.367
R843 B.n714 B.n713 163.367
R844 B.n713 B.n712 163.367
R845 B.n712 B.n39 163.367
R846 B.n708 B.n39 163.367
R847 B.n708 B.n707 163.367
R848 B.n707 B.n706 163.367
R849 B.n706 B.n41 163.367
R850 B.n702 B.n41 163.367
R851 B.n702 B.n701 163.367
R852 B.n701 B.n700 163.367
R853 B.n700 B.n43 163.367
R854 B.n696 B.n43 163.367
R855 B.n696 B.n695 163.367
R856 B.n695 B.n694 163.367
R857 B.n694 B.n45 163.367
R858 B.n690 B.n45 163.367
R859 B.n690 B.n689 163.367
R860 B.n689 B.n688 163.367
R861 B.n688 B.n47 163.367
R862 B.n684 B.n47 163.367
R863 B.n684 B.n683 163.367
R864 B.n683 B.n682 163.367
R865 B.n682 B.n49 163.367
R866 B.n678 B.n49 163.367
R867 B.n678 B.n677 163.367
R868 B.n677 B.n53 163.367
R869 B.n673 B.n53 163.367
R870 B.n673 B.n672 163.367
R871 B.n672 B.n671 163.367
R872 B.n671 B.n55 163.367
R873 B.n667 B.n55 163.367
R874 B.n667 B.n666 163.367
R875 B.n666 B.n665 163.367
R876 B.n665 B.n57 163.367
R877 B.n660 B.n57 163.367
R878 B.n660 B.n659 163.367
R879 B.n659 B.n658 163.367
R880 B.n658 B.n61 163.367
R881 B.n654 B.n61 163.367
R882 B.n654 B.n653 163.367
R883 B.n653 B.n652 163.367
R884 B.n652 B.n63 163.367
R885 B.n648 B.n63 163.367
R886 B.n648 B.n647 163.367
R887 B.n647 B.n646 163.367
R888 B.n646 B.n65 163.367
R889 B.n642 B.n65 163.367
R890 B.n642 B.n641 163.367
R891 B.n641 B.n640 163.367
R892 B.n640 B.n67 163.367
R893 B.n636 B.n67 163.367
R894 B.n636 B.n635 163.367
R895 B.n635 B.n634 163.367
R896 B.n634 B.n69 163.367
R897 B.n630 B.n69 163.367
R898 B.n630 B.n629 163.367
R899 B.n629 B.n628 163.367
R900 B.n628 B.n71 163.367
R901 B.n624 B.n71 163.367
R902 B.n624 B.n623 163.367
R903 B.n623 B.n622 163.367
R904 B.n622 B.n73 163.367
R905 B.n618 B.n73 163.367
R906 B.n618 B.n617 163.367
R907 B.n617 B.n616 163.367
R908 B.n616 B.n75 163.367
R909 B.n612 B.n75 163.367
R910 B.n612 B.n611 163.367
R911 B.n611 B.n610 163.367
R912 B.n610 B.n77 163.367
R913 B.n606 B.n77 163.367
R914 B.n606 B.n605 163.367
R915 B.n605 B.n604 163.367
R916 B.n604 B.n79 163.367
R917 B.n600 B.n79 163.367
R918 B.n600 B.n599 163.367
R919 B.n599 B.n598 163.367
R920 B.n598 B.n81 163.367
R921 B.n594 B.n81 163.367
R922 B.n594 B.n593 163.367
R923 B.n593 B.n592 163.367
R924 B.n592 B.n83 163.367
R925 B.n588 B.n83 163.367
R926 B.n588 B.n587 163.367
R927 B.n587 B.n586 163.367
R928 B.n586 B.n85 163.367
R929 B.n582 B.n85 163.367
R930 B.n582 B.n581 163.367
R931 B.n581 B.n580 163.367
R932 B.n580 B.n87 163.367
R933 B.n576 B.n87 163.367
R934 B.n576 B.n575 163.367
R935 B.n575 B.n574 163.367
R936 B.n574 B.n89 163.367
R937 B.n570 B.n89 163.367
R938 B.n156 B.t8 147.256
R939 B.n58 B.t4 147.256
R940 B.n164 B.t11 147.232
R941 B.n50 B.t1 147.232
R942 B.n157 B.t7 111.766
R943 B.n59 B.t5 111.766
R944 B.n165 B.t10 111.743
R945 B.n51 B.t2 111.743
R946 B.n158 B.n157 59.5399
R947 B.n356 B.n165 59.5399
R948 B.n52 B.n51 59.5399
R949 B.n662 B.n59 59.5399
R950 B.n157 B.n156 35.4914
R951 B.n165 B.n164 35.4914
R952 B.n51 B.n50 35.4914
R953 B.n59 B.n58 35.4914
R954 B.n770 B.n769 32.3127
R955 B.n571 B.n90 32.3127
R956 B.n464 B.n463 32.3127
R957 B.n265 B.n196 32.3127
R958 B B.n823 18.0485
R959 B.n769 B.n20 10.6151
R960 B.n765 B.n20 10.6151
R961 B.n765 B.n764 10.6151
R962 B.n764 B.n763 10.6151
R963 B.n763 B.n22 10.6151
R964 B.n759 B.n22 10.6151
R965 B.n759 B.n758 10.6151
R966 B.n758 B.n757 10.6151
R967 B.n757 B.n24 10.6151
R968 B.n753 B.n24 10.6151
R969 B.n753 B.n752 10.6151
R970 B.n752 B.n751 10.6151
R971 B.n751 B.n26 10.6151
R972 B.n747 B.n26 10.6151
R973 B.n747 B.n746 10.6151
R974 B.n746 B.n745 10.6151
R975 B.n745 B.n28 10.6151
R976 B.n741 B.n28 10.6151
R977 B.n741 B.n740 10.6151
R978 B.n740 B.n739 10.6151
R979 B.n739 B.n30 10.6151
R980 B.n735 B.n30 10.6151
R981 B.n735 B.n734 10.6151
R982 B.n734 B.n733 10.6151
R983 B.n733 B.n32 10.6151
R984 B.n729 B.n32 10.6151
R985 B.n729 B.n728 10.6151
R986 B.n728 B.n727 10.6151
R987 B.n727 B.n34 10.6151
R988 B.n723 B.n34 10.6151
R989 B.n723 B.n722 10.6151
R990 B.n722 B.n721 10.6151
R991 B.n721 B.n36 10.6151
R992 B.n717 B.n36 10.6151
R993 B.n717 B.n716 10.6151
R994 B.n716 B.n715 10.6151
R995 B.n715 B.n38 10.6151
R996 B.n711 B.n38 10.6151
R997 B.n711 B.n710 10.6151
R998 B.n710 B.n709 10.6151
R999 B.n709 B.n40 10.6151
R1000 B.n705 B.n40 10.6151
R1001 B.n705 B.n704 10.6151
R1002 B.n704 B.n703 10.6151
R1003 B.n703 B.n42 10.6151
R1004 B.n699 B.n42 10.6151
R1005 B.n699 B.n698 10.6151
R1006 B.n698 B.n697 10.6151
R1007 B.n697 B.n44 10.6151
R1008 B.n693 B.n44 10.6151
R1009 B.n693 B.n692 10.6151
R1010 B.n692 B.n691 10.6151
R1011 B.n691 B.n46 10.6151
R1012 B.n687 B.n46 10.6151
R1013 B.n687 B.n686 10.6151
R1014 B.n686 B.n685 10.6151
R1015 B.n685 B.n48 10.6151
R1016 B.n681 B.n48 10.6151
R1017 B.n681 B.n680 10.6151
R1018 B.n680 B.n679 10.6151
R1019 B.n676 B.n675 10.6151
R1020 B.n675 B.n674 10.6151
R1021 B.n674 B.n54 10.6151
R1022 B.n670 B.n54 10.6151
R1023 B.n670 B.n669 10.6151
R1024 B.n669 B.n668 10.6151
R1025 B.n668 B.n56 10.6151
R1026 B.n664 B.n56 10.6151
R1027 B.n664 B.n663 10.6151
R1028 B.n661 B.n60 10.6151
R1029 B.n657 B.n60 10.6151
R1030 B.n657 B.n656 10.6151
R1031 B.n656 B.n655 10.6151
R1032 B.n655 B.n62 10.6151
R1033 B.n651 B.n62 10.6151
R1034 B.n651 B.n650 10.6151
R1035 B.n650 B.n649 10.6151
R1036 B.n649 B.n64 10.6151
R1037 B.n645 B.n64 10.6151
R1038 B.n645 B.n644 10.6151
R1039 B.n644 B.n643 10.6151
R1040 B.n643 B.n66 10.6151
R1041 B.n639 B.n66 10.6151
R1042 B.n639 B.n638 10.6151
R1043 B.n638 B.n637 10.6151
R1044 B.n637 B.n68 10.6151
R1045 B.n633 B.n68 10.6151
R1046 B.n633 B.n632 10.6151
R1047 B.n632 B.n631 10.6151
R1048 B.n631 B.n70 10.6151
R1049 B.n627 B.n70 10.6151
R1050 B.n627 B.n626 10.6151
R1051 B.n626 B.n625 10.6151
R1052 B.n625 B.n72 10.6151
R1053 B.n621 B.n72 10.6151
R1054 B.n621 B.n620 10.6151
R1055 B.n620 B.n619 10.6151
R1056 B.n619 B.n74 10.6151
R1057 B.n615 B.n74 10.6151
R1058 B.n615 B.n614 10.6151
R1059 B.n614 B.n613 10.6151
R1060 B.n613 B.n76 10.6151
R1061 B.n609 B.n76 10.6151
R1062 B.n609 B.n608 10.6151
R1063 B.n608 B.n607 10.6151
R1064 B.n607 B.n78 10.6151
R1065 B.n603 B.n78 10.6151
R1066 B.n603 B.n602 10.6151
R1067 B.n602 B.n601 10.6151
R1068 B.n601 B.n80 10.6151
R1069 B.n597 B.n80 10.6151
R1070 B.n597 B.n596 10.6151
R1071 B.n596 B.n595 10.6151
R1072 B.n595 B.n82 10.6151
R1073 B.n591 B.n82 10.6151
R1074 B.n591 B.n590 10.6151
R1075 B.n590 B.n589 10.6151
R1076 B.n589 B.n84 10.6151
R1077 B.n585 B.n84 10.6151
R1078 B.n585 B.n584 10.6151
R1079 B.n584 B.n583 10.6151
R1080 B.n583 B.n86 10.6151
R1081 B.n579 B.n86 10.6151
R1082 B.n579 B.n578 10.6151
R1083 B.n578 B.n577 10.6151
R1084 B.n577 B.n88 10.6151
R1085 B.n573 B.n88 10.6151
R1086 B.n573 B.n572 10.6151
R1087 B.n572 B.n571 10.6151
R1088 B.n465 B.n464 10.6151
R1089 B.n465 B.n124 10.6151
R1090 B.n469 B.n124 10.6151
R1091 B.n470 B.n469 10.6151
R1092 B.n471 B.n470 10.6151
R1093 B.n471 B.n122 10.6151
R1094 B.n475 B.n122 10.6151
R1095 B.n476 B.n475 10.6151
R1096 B.n477 B.n476 10.6151
R1097 B.n477 B.n120 10.6151
R1098 B.n481 B.n120 10.6151
R1099 B.n482 B.n481 10.6151
R1100 B.n483 B.n482 10.6151
R1101 B.n483 B.n118 10.6151
R1102 B.n487 B.n118 10.6151
R1103 B.n488 B.n487 10.6151
R1104 B.n489 B.n488 10.6151
R1105 B.n489 B.n116 10.6151
R1106 B.n493 B.n116 10.6151
R1107 B.n494 B.n493 10.6151
R1108 B.n495 B.n494 10.6151
R1109 B.n495 B.n114 10.6151
R1110 B.n499 B.n114 10.6151
R1111 B.n500 B.n499 10.6151
R1112 B.n501 B.n500 10.6151
R1113 B.n501 B.n112 10.6151
R1114 B.n505 B.n112 10.6151
R1115 B.n506 B.n505 10.6151
R1116 B.n507 B.n506 10.6151
R1117 B.n507 B.n110 10.6151
R1118 B.n511 B.n110 10.6151
R1119 B.n512 B.n511 10.6151
R1120 B.n513 B.n512 10.6151
R1121 B.n513 B.n108 10.6151
R1122 B.n517 B.n108 10.6151
R1123 B.n518 B.n517 10.6151
R1124 B.n519 B.n518 10.6151
R1125 B.n519 B.n106 10.6151
R1126 B.n523 B.n106 10.6151
R1127 B.n524 B.n523 10.6151
R1128 B.n525 B.n524 10.6151
R1129 B.n525 B.n104 10.6151
R1130 B.n529 B.n104 10.6151
R1131 B.n530 B.n529 10.6151
R1132 B.n531 B.n530 10.6151
R1133 B.n531 B.n102 10.6151
R1134 B.n535 B.n102 10.6151
R1135 B.n536 B.n535 10.6151
R1136 B.n537 B.n536 10.6151
R1137 B.n537 B.n100 10.6151
R1138 B.n541 B.n100 10.6151
R1139 B.n542 B.n541 10.6151
R1140 B.n543 B.n542 10.6151
R1141 B.n543 B.n98 10.6151
R1142 B.n547 B.n98 10.6151
R1143 B.n548 B.n547 10.6151
R1144 B.n549 B.n548 10.6151
R1145 B.n549 B.n96 10.6151
R1146 B.n553 B.n96 10.6151
R1147 B.n554 B.n553 10.6151
R1148 B.n555 B.n554 10.6151
R1149 B.n555 B.n94 10.6151
R1150 B.n559 B.n94 10.6151
R1151 B.n560 B.n559 10.6151
R1152 B.n561 B.n560 10.6151
R1153 B.n561 B.n92 10.6151
R1154 B.n565 B.n92 10.6151
R1155 B.n566 B.n565 10.6151
R1156 B.n567 B.n566 10.6151
R1157 B.n567 B.n90 10.6151
R1158 B.n266 B.n265 10.6151
R1159 B.n267 B.n266 10.6151
R1160 B.n267 B.n194 10.6151
R1161 B.n271 B.n194 10.6151
R1162 B.n272 B.n271 10.6151
R1163 B.n273 B.n272 10.6151
R1164 B.n273 B.n192 10.6151
R1165 B.n277 B.n192 10.6151
R1166 B.n278 B.n277 10.6151
R1167 B.n279 B.n278 10.6151
R1168 B.n279 B.n190 10.6151
R1169 B.n283 B.n190 10.6151
R1170 B.n284 B.n283 10.6151
R1171 B.n285 B.n284 10.6151
R1172 B.n285 B.n188 10.6151
R1173 B.n289 B.n188 10.6151
R1174 B.n290 B.n289 10.6151
R1175 B.n291 B.n290 10.6151
R1176 B.n291 B.n186 10.6151
R1177 B.n295 B.n186 10.6151
R1178 B.n296 B.n295 10.6151
R1179 B.n297 B.n296 10.6151
R1180 B.n297 B.n184 10.6151
R1181 B.n301 B.n184 10.6151
R1182 B.n302 B.n301 10.6151
R1183 B.n303 B.n302 10.6151
R1184 B.n303 B.n182 10.6151
R1185 B.n307 B.n182 10.6151
R1186 B.n308 B.n307 10.6151
R1187 B.n309 B.n308 10.6151
R1188 B.n309 B.n180 10.6151
R1189 B.n313 B.n180 10.6151
R1190 B.n314 B.n313 10.6151
R1191 B.n315 B.n314 10.6151
R1192 B.n315 B.n178 10.6151
R1193 B.n319 B.n178 10.6151
R1194 B.n320 B.n319 10.6151
R1195 B.n321 B.n320 10.6151
R1196 B.n321 B.n176 10.6151
R1197 B.n325 B.n176 10.6151
R1198 B.n326 B.n325 10.6151
R1199 B.n327 B.n326 10.6151
R1200 B.n327 B.n174 10.6151
R1201 B.n331 B.n174 10.6151
R1202 B.n332 B.n331 10.6151
R1203 B.n333 B.n332 10.6151
R1204 B.n333 B.n172 10.6151
R1205 B.n337 B.n172 10.6151
R1206 B.n338 B.n337 10.6151
R1207 B.n339 B.n338 10.6151
R1208 B.n339 B.n170 10.6151
R1209 B.n343 B.n170 10.6151
R1210 B.n344 B.n343 10.6151
R1211 B.n345 B.n344 10.6151
R1212 B.n345 B.n168 10.6151
R1213 B.n349 B.n168 10.6151
R1214 B.n350 B.n349 10.6151
R1215 B.n351 B.n350 10.6151
R1216 B.n351 B.n166 10.6151
R1217 B.n355 B.n166 10.6151
R1218 B.n358 B.n357 10.6151
R1219 B.n358 B.n162 10.6151
R1220 B.n362 B.n162 10.6151
R1221 B.n363 B.n362 10.6151
R1222 B.n364 B.n363 10.6151
R1223 B.n364 B.n160 10.6151
R1224 B.n368 B.n160 10.6151
R1225 B.n369 B.n368 10.6151
R1226 B.n370 B.n369 10.6151
R1227 B.n374 B.n373 10.6151
R1228 B.n375 B.n374 10.6151
R1229 B.n375 B.n154 10.6151
R1230 B.n379 B.n154 10.6151
R1231 B.n380 B.n379 10.6151
R1232 B.n381 B.n380 10.6151
R1233 B.n381 B.n152 10.6151
R1234 B.n385 B.n152 10.6151
R1235 B.n386 B.n385 10.6151
R1236 B.n387 B.n386 10.6151
R1237 B.n387 B.n150 10.6151
R1238 B.n391 B.n150 10.6151
R1239 B.n392 B.n391 10.6151
R1240 B.n393 B.n392 10.6151
R1241 B.n393 B.n148 10.6151
R1242 B.n397 B.n148 10.6151
R1243 B.n398 B.n397 10.6151
R1244 B.n399 B.n398 10.6151
R1245 B.n399 B.n146 10.6151
R1246 B.n403 B.n146 10.6151
R1247 B.n404 B.n403 10.6151
R1248 B.n405 B.n404 10.6151
R1249 B.n405 B.n144 10.6151
R1250 B.n409 B.n144 10.6151
R1251 B.n410 B.n409 10.6151
R1252 B.n411 B.n410 10.6151
R1253 B.n411 B.n142 10.6151
R1254 B.n415 B.n142 10.6151
R1255 B.n416 B.n415 10.6151
R1256 B.n417 B.n416 10.6151
R1257 B.n417 B.n140 10.6151
R1258 B.n421 B.n140 10.6151
R1259 B.n422 B.n421 10.6151
R1260 B.n423 B.n422 10.6151
R1261 B.n423 B.n138 10.6151
R1262 B.n427 B.n138 10.6151
R1263 B.n428 B.n427 10.6151
R1264 B.n429 B.n428 10.6151
R1265 B.n429 B.n136 10.6151
R1266 B.n433 B.n136 10.6151
R1267 B.n434 B.n433 10.6151
R1268 B.n435 B.n434 10.6151
R1269 B.n435 B.n134 10.6151
R1270 B.n439 B.n134 10.6151
R1271 B.n440 B.n439 10.6151
R1272 B.n441 B.n440 10.6151
R1273 B.n441 B.n132 10.6151
R1274 B.n445 B.n132 10.6151
R1275 B.n446 B.n445 10.6151
R1276 B.n447 B.n446 10.6151
R1277 B.n447 B.n130 10.6151
R1278 B.n451 B.n130 10.6151
R1279 B.n452 B.n451 10.6151
R1280 B.n453 B.n452 10.6151
R1281 B.n453 B.n128 10.6151
R1282 B.n457 B.n128 10.6151
R1283 B.n458 B.n457 10.6151
R1284 B.n459 B.n458 10.6151
R1285 B.n459 B.n126 10.6151
R1286 B.n463 B.n126 10.6151
R1287 B.n261 B.n196 10.6151
R1288 B.n261 B.n260 10.6151
R1289 B.n260 B.n259 10.6151
R1290 B.n259 B.n198 10.6151
R1291 B.n255 B.n198 10.6151
R1292 B.n255 B.n254 10.6151
R1293 B.n254 B.n253 10.6151
R1294 B.n253 B.n200 10.6151
R1295 B.n249 B.n200 10.6151
R1296 B.n249 B.n248 10.6151
R1297 B.n248 B.n247 10.6151
R1298 B.n247 B.n202 10.6151
R1299 B.n243 B.n202 10.6151
R1300 B.n243 B.n242 10.6151
R1301 B.n242 B.n241 10.6151
R1302 B.n241 B.n204 10.6151
R1303 B.n237 B.n204 10.6151
R1304 B.n237 B.n236 10.6151
R1305 B.n236 B.n235 10.6151
R1306 B.n235 B.n206 10.6151
R1307 B.n231 B.n206 10.6151
R1308 B.n231 B.n230 10.6151
R1309 B.n230 B.n229 10.6151
R1310 B.n229 B.n208 10.6151
R1311 B.n225 B.n208 10.6151
R1312 B.n225 B.n224 10.6151
R1313 B.n224 B.n223 10.6151
R1314 B.n223 B.n210 10.6151
R1315 B.n219 B.n210 10.6151
R1316 B.n219 B.n218 10.6151
R1317 B.n218 B.n217 10.6151
R1318 B.n217 B.n212 10.6151
R1319 B.n213 B.n212 10.6151
R1320 B.n213 B.n0 10.6151
R1321 B.n819 B.n1 10.6151
R1322 B.n819 B.n818 10.6151
R1323 B.n818 B.n817 10.6151
R1324 B.n817 B.n4 10.6151
R1325 B.n813 B.n4 10.6151
R1326 B.n813 B.n812 10.6151
R1327 B.n812 B.n811 10.6151
R1328 B.n811 B.n6 10.6151
R1329 B.n807 B.n6 10.6151
R1330 B.n807 B.n806 10.6151
R1331 B.n806 B.n805 10.6151
R1332 B.n805 B.n8 10.6151
R1333 B.n801 B.n8 10.6151
R1334 B.n801 B.n800 10.6151
R1335 B.n800 B.n799 10.6151
R1336 B.n799 B.n10 10.6151
R1337 B.n795 B.n10 10.6151
R1338 B.n795 B.n794 10.6151
R1339 B.n794 B.n793 10.6151
R1340 B.n793 B.n12 10.6151
R1341 B.n789 B.n12 10.6151
R1342 B.n789 B.n788 10.6151
R1343 B.n788 B.n787 10.6151
R1344 B.n787 B.n14 10.6151
R1345 B.n783 B.n14 10.6151
R1346 B.n783 B.n782 10.6151
R1347 B.n782 B.n781 10.6151
R1348 B.n781 B.n16 10.6151
R1349 B.n777 B.n16 10.6151
R1350 B.n777 B.n776 10.6151
R1351 B.n776 B.n775 10.6151
R1352 B.n775 B.n18 10.6151
R1353 B.n771 B.n18 10.6151
R1354 B.n771 B.n770 10.6151
R1355 B.n679 B.n52 9.36635
R1356 B.n662 B.n661 9.36635
R1357 B.n356 B.n355 9.36635
R1358 B.n373 B.n158 9.36635
R1359 B.n823 B.n0 2.81026
R1360 B.n823 B.n1 2.81026
R1361 B.n676 B.n52 1.24928
R1362 B.n663 B.n662 1.24928
R1363 B.n357 B.n356 1.24928
R1364 B.n370 B.n158 1.24928
R1365 VN.n5 VN.t4 334.392
R1366 VN.n24 VN.t1 334.392
R1367 VN.n4 VN.t2 299.644
R1368 VN.n10 VN.t5 299.644
R1369 VN.n17 VN.t3 299.644
R1370 VN.n23 VN.t0 299.644
R1371 VN.n29 VN.t7 299.644
R1372 VN.n36 VN.t6 299.644
R1373 VN.n18 VN.n17 173.779
R1374 VN.n37 VN.n36 173.779
R1375 VN.n35 VN.n19 161.3
R1376 VN.n34 VN.n33 161.3
R1377 VN.n32 VN.n20 161.3
R1378 VN.n31 VN.n30 161.3
R1379 VN.n28 VN.n21 161.3
R1380 VN.n27 VN.n26 161.3
R1381 VN.n25 VN.n22 161.3
R1382 VN.n16 VN.n0 161.3
R1383 VN.n15 VN.n14 161.3
R1384 VN.n13 VN.n1 161.3
R1385 VN.n12 VN.n11 161.3
R1386 VN.n9 VN.n2 161.3
R1387 VN.n8 VN.n7 161.3
R1388 VN.n6 VN.n3 161.3
R1389 VN.n15 VN.n1 56.5193
R1390 VN.n34 VN.n20 56.5193
R1391 VN VN.n37 51.1236
R1392 VN.n5 VN.n4 46.2606
R1393 VN.n24 VN.n23 46.2606
R1394 VN.n8 VN.n3 40.4934
R1395 VN.n9 VN.n8 40.4934
R1396 VN.n27 VN.n22 40.4934
R1397 VN.n28 VN.n27 40.4934
R1398 VN.n11 VN.n1 24.4675
R1399 VN.n16 VN.n15 24.4675
R1400 VN.n30 VN.n20 24.4675
R1401 VN.n35 VN.n34 24.4675
R1402 VN.n4 VN.n3 20.3081
R1403 VN.n10 VN.n9 20.3081
R1404 VN.n23 VN.n22 20.3081
R1405 VN.n29 VN.n28 20.3081
R1406 VN.n25 VN.n24 17.5886
R1407 VN.n6 VN.n5 17.5886
R1408 VN.n17 VN.n16 11.9893
R1409 VN.n36 VN.n35 11.9893
R1410 VN.n11 VN.n10 4.15989
R1411 VN.n30 VN.n29 4.15989
R1412 VN.n37 VN.n19 0.189894
R1413 VN.n33 VN.n19 0.189894
R1414 VN.n33 VN.n32 0.189894
R1415 VN.n32 VN.n31 0.189894
R1416 VN.n31 VN.n21 0.189894
R1417 VN.n26 VN.n21 0.189894
R1418 VN.n26 VN.n25 0.189894
R1419 VN.n7 VN.n6 0.189894
R1420 VN.n7 VN.n2 0.189894
R1421 VN.n12 VN.n2 0.189894
R1422 VN.n13 VN.n12 0.189894
R1423 VN.n14 VN.n13 0.189894
R1424 VN.n14 VN.n0 0.189894
R1425 VN.n18 VN.n0 0.189894
R1426 VN VN.n18 0.0516364
R1427 VDD2.n2 VDD2.n1 70.2354
R1428 VDD2.n2 VDD2.n0 70.2354
R1429 VDD2 VDD2.n5 70.2326
R1430 VDD2.n4 VDD2.n3 69.5022
R1431 VDD2.n4 VDD2.n2 46.892
R1432 VDD2.n5 VDD2.t7 1.7434
R1433 VDD2.n5 VDD2.t6 1.7434
R1434 VDD2.n3 VDD2.t1 1.7434
R1435 VDD2.n3 VDD2.t0 1.7434
R1436 VDD2.n1 VDD2.t2 1.7434
R1437 VDD2.n1 VDD2.t4 1.7434
R1438 VDD2.n0 VDD2.t3 1.7434
R1439 VDD2.n0 VDD2.t5 1.7434
R1440 VDD2 VDD2.n4 0.847483
C0 VN VTAIL 11.3044f
C1 VP VDD2 0.402688f
C2 VP w_n2800_n4698# 5.87141f
C3 B VDD2 1.55511f
C4 VP VDD1 11.773499f
C5 B w_n2800_n4698# 10.2949f
C6 B VDD1 1.49366f
C7 VN VDD2 11.5215f
C8 VP B 1.64531f
C9 VN w_n2800_n4698# 5.51115f
C10 VN VDD1 0.149808f
C11 VTAIL VDD2 11.595901f
C12 w_n2800_n4698# VTAIL 5.71847f
C13 VN VP 7.54714f
C14 VTAIL VDD1 11.5488f
C15 VN B 1.04726f
C16 VP VTAIL 11.3185f
C17 B VTAIL 6.40422f
C18 w_n2800_n4698# VDD2 1.84067f
C19 VDD1 VDD2 1.22323f
C20 w_n2800_n4698# VDD1 1.77209f
C21 VDD2 VSUBS 1.675347f
C22 VDD1 VSUBS 2.12405f
C23 VTAIL VSUBS 1.418197f
C24 VN VSUBS 5.77284f
C25 VP VSUBS 2.697304f
C26 B VSUBS 4.33756f
C27 w_n2800_n4698# VSUBS 0.160776p
C28 VDD2.t3 VSUBS 0.36891f
C29 VDD2.t5 VSUBS 0.36891f
C30 VDD2.n0 VSUBS 3.08849f
C31 VDD2.t2 VSUBS 0.36891f
C32 VDD2.t4 VSUBS 0.36891f
C33 VDD2.n1 VSUBS 3.08849f
C34 VDD2.n2 VSUBS 3.62804f
C35 VDD2.t1 VSUBS 0.36891f
C36 VDD2.t0 VSUBS 0.36891f
C37 VDD2.n3 VSUBS 3.08129f
C38 VDD2.n4 VSUBS 3.36498f
C39 VDD2.t7 VSUBS 0.36891f
C40 VDD2.t6 VSUBS 0.36891f
C41 VDD2.n5 VSUBS 3.08844f
C42 VN.n0 VSUBS 0.03544f
C43 VN.t3 VSUBS 2.72884f
C44 VN.n1 VSUBS 0.059637f
C45 VN.n2 VSUBS 0.03544f
C46 VN.t5 VSUBS 2.72884f
C47 VN.n3 VSUBS 0.064892f
C48 VN.t4 VSUBS 2.84288f
C49 VN.t2 VSUBS 2.72884f
C50 VN.n4 VSUBS 1.03593f
C51 VN.n5 VSUBS 1.03949f
C52 VN.n6 VSUBS 0.225346f
C53 VN.n7 VSUBS 0.03544f
C54 VN.n8 VSUBS 0.02865f
C55 VN.n9 VSUBS 0.064892f
C56 VN.n10 VSUBS 0.958775f
C57 VN.n11 VSUBS 0.038984f
C58 VN.n12 VSUBS 0.03544f
C59 VN.n13 VSUBS 0.03544f
C60 VN.n14 VSUBS 0.03544f
C61 VN.n15 VSUBS 0.043836f
C62 VN.n16 VSUBS 0.049419f
C63 VN.n17 VSUBS 1.03491f
C64 VN.n18 VSUBS 0.033355f
C65 VN.n19 VSUBS 0.03544f
C66 VN.t6 VSUBS 2.72884f
C67 VN.n20 VSUBS 0.059637f
C68 VN.n21 VSUBS 0.03544f
C69 VN.t7 VSUBS 2.72884f
C70 VN.n22 VSUBS 0.064892f
C71 VN.t1 VSUBS 2.84288f
C72 VN.t0 VSUBS 2.72884f
C73 VN.n23 VSUBS 1.03593f
C74 VN.n24 VSUBS 1.03949f
C75 VN.n25 VSUBS 0.225346f
C76 VN.n26 VSUBS 0.03544f
C77 VN.n27 VSUBS 0.02865f
C78 VN.n28 VSUBS 0.064892f
C79 VN.n29 VSUBS 0.958775f
C80 VN.n30 VSUBS 0.038984f
C81 VN.n31 VSUBS 0.03544f
C82 VN.n32 VSUBS 0.03544f
C83 VN.n33 VSUBS 0.03544f
C84 VN.n34 VSUBS 0.043836f
C85 VN.n35 VSUBS 0.049419f
C86 VN.n36 VSUBS 1.03491f
C87 VN.n37 VSUBS 1.99874f
C88 B.n0 VSUBS 0.004311f
C89 B.n1 VSUBS 0.004311f
C90 B.n2 VSUBS 0.006817f
C91 B.n3 VSUBS 0.006817f
C92 B.n4 VSUBS 0.006817f
C93 B.n5 VSUBS 0.006817f
C94 B.n6 VSUBS 0.006817f
C95 B.n7 VSUBS 0.006817f
C96 B.n8 VSUBS 0.006817f
C97 B.n9 VSUBS 0.006817f
C98 B.n10 VSUBS 0.006817f
C99 B.n11 VSUBS 0.006817f
C100 B.n12 VSUBS 0.006817f
C101 B.n13 VSUBS 0.006817f
C102 B.n14 VSUBS 0.006817f
C103 B.n15 VSUBS 0.006817f
C104 B.n16 VSUBS 0.006817f
C105 B.n17 VSUBS 0.006817f
C106 B.n18 VSUBS 0.006817f
C107 B.n19 VSUBS 0.015414f
C108 B.n20 VSUBS 0.006817f
C109 B.n21 VSUBS 0.006817f
C110 B.n22 VSUBS 0.006817f
C111 B.n23 VSUBS 0.006817f
C112 B.n24 VSUBS 0.006817f
C113 B.n25 VSUBS 0.006817f
C114 B.n26 VSUBS 0.006817f
C115 B.n27 VSUBS 0.006817f
C116 B.n28 VSUBS 0.006817f
C117 B.n29 VSUBS 0.006817f
C118 B.n30 VSUBS 0.006817f
C119 B.n31 VSUBS 0.006817f
C120 B.n32 VSUBS 0.006817f
C121 B.n33 VSUBS 0.006817f
C122 B.n34 VSUBS 0.006817f
C123 B.n35 VSUBS 0.006817f
C124 B.n36 VSUBS 0.006817f
C125 B.n37 VSUBS 0.006817f
C126 B.n38 VSUBS 0.006817f
C127 B.n39 VSUBS 0.006817f
C128 B.n40 VSUBS 0.006817f
C129 B.n41 VSUBS 0.006817f
C130 B.n42 VSUBS 0.006817f
C131 B.n43 VSUBS 0.006817f
C132 B.n44 VSUBS 0.006817f
C133 B.n45 VSUBS 0.006817f
C134 B.n46 VSUBS 0.006817f
C135 B.n47 VSUBS 0.006817f
C136 B.n48 VSUBS 0.006817f
C137 B.n49 VSUBS 0.006817f
C138 B.t2 VSUBS 0.614714f
C139 B.t1 VSUBS 0.62823f
C140 B.t0 VSUBS 1.15583f
C141 B.n50 VSUBS 0.274957f
C142 B.n51 VSUBS 0.065795f
C143 B.n52 VSUBS 0.015795f
C144 B.n53 VSUBS 0.006817f
C145 B.n54 VSUBS 0.006817f
C146 B.n55 VSUBS 0.006817f
C147 B.n56 VSUBS 0.006817f
C148 B.n57 VSUBS 0.006817f
C149 B.t5 VSUBS 0.614691f
C150 B.t4 VSUBS 0.628211f
C151 B.t3 VSUBS 1.15583f
C152 B.n58 VSUBS 0.274977f
C153 B.n59 VSUBS 0.065819f
C154 B.n60 VSUBS 0.006817f
C155 B.n61 VSUBS 0.006817f
C156 B.n62 VSUBS 0.006817f
C157 B.n63 VSUBS 0.006817f
C158 B.n64 VSUBS 0.006817f
C159 B.n65 VSUBS 0.006817f
C160 B.n66 VSUBS 0.006817f
C161 B.n67 VSUBS 0.006817f
C162 B.n68 VSUBS 0.006817f
C163 B.n69 VSUBS 0.006817f
C164 B.n70 VSUBS 0.006817f
C165 B.n71 VSUBS 0.006817f
C166 B.n72 VSUBS 0.006817f
C167 B.n73 VSUBS 0.006817f
C168 B.n74 VSUBS 0.006817f
C169 B.n75 VSUBS 0.006817f
C170 B.n76 VSUBS 0.006817f
C171 B.n77 VSUBS 0.006817f
C172 B.n78 VSUBS 0.006817f
C173 B.n79 VSUBS 0.006817f
C174 B.n80 VSUBS 0.006817f
C175 B.n81 VSUBS 0.006817f
C176 B.n82 VSUBS 0.006817f
C177 B.n83 VSUBS 0.006817f
C178 B.n84 VSUBS 0.006817f
C179 B.n85 VSUBS 0.006817f
C180 B.n86 VSUBS 0.006817f
C181 B.n87 VSUBS 0.006817f
C182 B.n88 VSUBS 0.006817f
C183 B.n89 VSUBS 0.006817f
C184 B.n90 VSUBS 0.016228f
C185 B.n91 VSUBS 0.006817f
C186 B.n92 VSUBS 0.006817f
C187 B.n93 VSUBS 0.006817f
C188 B.n94 VSUBS 0.006817f
C189 B.n95 VSUBS 0.006817f
C190 B.n96 VSUBS 0.006817f
C191 B.n97 VSUBS 0.006817f
C192 B.n98 VSUBS 0.006817f
C193 B.n99 VSUBS 0.006817f
C194 B.n100 VSUBS 0.006817f
C195 B.n101 VSUBS 0.006817f
C196 B.n102 VSUBS 0.006817f
C197 B.n103 VSUBS 0.006817f
C198 B.n104 VSUBS 0.006817f
C199 B.n105 VSUBS 0.006817f
C200 B.n106 VSUBS 0.006817f
C201 B.n107 VSUBS 0.006817f
C202 B.n108 VSUBS 0.006817f
C203 B.n109 VSUBS 0.006817f
C204 B.n110 VSUBS 0.006817f
C205 B.n111 VSUBS 0.006817f
C206 B.n112 VSUBS 0.006817f
C207 B.n113 VSUBS 0.006817f
C208 B.n114 VSUBS 0.006817f
C209 B.n115 VSUBS 0.006817f
C210 B.n116 VSUBS 0.006817f
C211 B.n117 VSUBS 0.006817f
C212 B.n118 VSUBS 0.006817f
C213 B.n119 VSUBS 0.006817f
C214 B.n120 VSUBS 0.006817f
C215 B.n121 VSUBS 0.006817f
C216 B.n122 VSUBS 0.006817f
C217 B.n123 VSUBS 0.006817f
C218 B.n124 VSUBS 0.006817f
C219 B.n125 VSUBS 0.015414f
C220 B.n126 VSUBS 0.006817f
C221 B.n127 VSUBS 0.006817f
C222 B.n128 VSUBS 0.006817f
C223 B.n129 VSUBS 0.006817f
C224 B.n130 VSUBS 0.006817f
C225 B.n131 VSUBS 0.006817f
C226 B.n132 VSUBS 0.006817f
C227 B.n133 VSUBS 0.006817f
C228 B.n134 VSUBS 0.006817f
C229 B.n135 VSUBS 0.006817f
C230 B.n136 VSUBS 0.006817f
C231 B.n137 VSUBS 0.006817f
C232 B.n138 VSUBS 0.006817f
C233 B.n139 VSUBS 0.006817f
C234 B.n140 VSUBS 0.006817f
C235 B.n141 VSUBS 0.006817f
C236 B.n142 VSUBS 0.006817f
C237 B.n143 VSUBS 0.006817f
C238 B.n144 VSUBS 0.006817f
C239 B.n145 VSUBS 0.006817f
C240 B.n146 VSUBS 0.006817f
C241 B.n147 VSUBS 0.006817f
C242 B.n148 VSUBS 0.006817f
C243 B.n149 VSUBS 0.006817f
C244 B.n150 VSUBS 0.006817f
C245 B.n151 VSUBS 0.006817f
C246 B.n152 VSUBS 0.006817f
C247 B.n153 VSUBS 0.006817f
C248 B.n154 VSUBS 0.006817f
C249 B.n155 VSUBS 0.006817f
C250 B.t7 VSUBS 0.614691f
C251 B.t8 VSUBS 0.628211f
C252 B.t6 VSUBS 1.15583f
C253 B.n156 VSUBS 0.274977f
C254 B.n157 VSUBS 0.065819f
C255 B.n158 VSUBS 0.015795f
C256 B.n159 VSUBS 0.006817f
C257 B.n160 VSUBS 0.006817f
C258 B.n161 VSUBS 0.006817f
C259 B.n162 VSUBS 0.006817f
C260 B.n163 VSUBS 0.006817f
C261 B.t10 VSUBS 0.614714f
C262 B.t11 VSUBS 0.62823f
C263 B.t9 VSUBS 1.15583f
C264 B.n164 VSUBS 0.274957f
C265 B.n165 VSUBS 0.065795f
C266 B.n166 VSUBS 0.006817f
C267 B.n167 VSUBS 0.006817f
C268 B.n168 VSUBS 0.006817f
C269 B.n169 VSUBS 0.006817f
C270 B.n170 VSUBS 0.006817f
C271 B.n171 VSUBS 0.006817f
C272 B.n172 VSUBS 0.006817f
C273 B.n173 VSUBS 0.006817f
C274 B.n174 VSUBS 0.006817f
C275 B.n175 VSUBS 0.006817f
C276 B.n176 VSUBS 0.006817f
C277 B.n177 VSUBS 0.006817f
C278 B.n178 VSUBS 0.006817f
C279 B.n179 VSUBS 0.006817f
C280 B.n180 VSUBS 0.006817f
C281 B.n181 VSUBS 0.006817f
C282 B.n182 VSUBS 0.006817f
C283 B.n183 VSUBS 0.006817f
C284 B.n184 VSUBS 0.006817f
C285 B.n185 VSUBS 0.006817f
C286 B.n186 VSUBS 0.006817f
C287 B.n187 VSUBS 0.006817f
C288 B.n188 VSUBS 0.006817f
C289 B.n189 VSUBS 0.006817f
C290 B.n190 VSUBS 0.006817f
C291 B.n191 VSUBS 0.006817f
C292 B.n192 VSUBS 0.006817f
C293 B.n193 VSUBS 0.006817f
C294 B.n194 VSUBS 0.006817f
C295 B.n195 VSUBS 0.006817f
C296 B.n196 VSUBS 0.015414f
C297 B.n197 VSUBS 0.006817f
C298 B.n198 VSUBS 0.006817f
C299 B.n199 VSUBS 0.006817f
C300 B.n200 VSUBS 0.006817f
C301 B.n201 VSUBS 0.006817f
C302 B.n202 VSUBS 0.006817f
C303 B.n203 VSUBS 0.006817f
C304 B.n204 VSUBS 0.006817f
C305 B.n205 VSUBS 0.006817f
C306 B.n206 VSUBS 0.006817f
C307 B.n207 VSUBS 0.006817f
C308 B.n208 VSUBS 0.006817f
C309 B.n209 VSUBS 0.006817f
C310 B.n210 VSUBS 0.006817f
C311 B.n211 VSUBS 0.006817f
C312 B.n212 VSUBS 0.006817f
C313 B.n213 VSUBS 0.006817f
C314 B.n214 VSUBS 0.006817f
C315 B.n215 VSUBS 0.006817f
C316 B.n216 VSUBS 0.006817f
C317 B.n217 VSUBS 0.006817f
C318 B.n218 VSUBS 0.006817f
C319 B.n219 VSUBS 0.006817f
C320 B.n220 VSUBS 0.006817f
C321 B.n221 VSUBS 0.006817f
C322 B.n222 VSUBS 0.006817f
C323 B.n223 VSUBS 0.006817f
C324 B.n224 VSUBS 0.006817f
C325 B.n225 VSUBS 0.006817f
C326 B.n226 VSUBS 0.006817f
C327 B.n227 VSUBS 0.006817f
C328 B.n228 VSUBS 0.006817f
C329 B.n229 VSUBS 0.006817f
C330 B.n230 VSUBS 0.006817f
C331 B.n231 VSUBS 0.006817f
C332 B.n232 VSUBS 0.006817f
C333 B.n233 VSUBS 0.006817f
C334 B.n234 VSUBS 0.006817f
C335 B.n235 VSUBS 0.006817f
C336 B.n236 VSUBS 0.006817f
C337 B.n237 VSUBS 0.006817f
C338 B.n238 VSUBS 0.006817f
C339 B.n239 VSUBS 0.006817f
C340 B.n240 VSUBS 0.006817f
C341 B.n241 VSUBS 0.006817f
C342 B.n242 VSUBS 0.006817f
C343 B.n243 VSUBS 0.006817f
C344 B.n244 VSUBS 0.006817f
C345 B.n245 VSUBS 0.006817f
C346 B.n246 VSUBS 0.006817f
C347 B.n247 VSUBS 0.006817f
C348 B.n248 VSUBS 0.006817f
C349 B.n249 VSUBS 0.006817f
C350 B.n250 VSUBS 0.006817f
C351 B.n251 VSUBS 0.006817f
C352 B.n252 VSUBS 0.006817f
C353 B.n253 VSUBS 0.006817f
C354 B.n254 VSUBS 0.006817f
C355 B.n255 VSUBS 0.006817f
C356 B.n256 VSUBS 0.006817f
C357 B.n257 VSUBS 0.006817f
C358 B.n258 VSUBS 0.006817f
C359 B.n259 VSUBS 0.006817f
C360 B.n260 VSUBS 0.006817f
C361 B.n261 VSUBS 0.006817f
C362 B.n262 VSUBS 0.006817f
C363 B.n263 VSUBS 0.015414f
C364 B.n264 VSUBS 0.016267f
C365 B.n265 VSUBS 0.016267f
C366 B.n266 VSUBS 0.006817f
C367 B.n267 VSUBS 0.006817f
C368 B.n268 VSUBS 0.006817f
C369 B.n269 VSUBS 0.006817f
C370 B.n270 VSUBS 0.006817f
C371 B.n271 VSUBS 0.006817f
C372 B.n272 VSUBS 0.006817f
C373 B.n273 VSUBS 0.006817f
C374 B.n274 VSUBS 0.006817f
C375 B.n275 VSUBS 0.006817f
C376 B.n276 VSUBS 0.006817f
C377 B.n277 VSUBS 0.006817f
C378 B.n278 VSUBS 0.006817f
C379 B.n279 VSUBS 0.006817f
C380 B.n280 VSUBS 0.006817f
C381 B.n281 VSUBS 0.006817f
C382 B.n282 VSUBS 0.006817f
C383 B.n283 VSUBS 0.006817f
C384 B.n284 VSUBS 0.006817f
C385 B.n285 VSUBS 0.006817f
C386 B.n286 VSUBS 0.006817f
C387 B.n287 VSUBS 0.006817f
C388 B.n288 VSUBS 0.006817f
C389 B.n289 VSUBS 0.006817f
C390 B.n290 VSUBS 0.006817f
C391 B.n291 VSUBS 0.006817f
C392 B.n292 VSUBS 0.006817f
C393 B.n293 VSUBS 0.006817f
C394 B.n294 VSUBS 0.006817f
C395 B.n295 VSUBS 0.006817f
C396 B.n296 VSUBS 0.006817f
C397 B.n297 VSUBS 0.006817f
C398 B.n298 VSUBS 0.006817f
C399 B.n299 VSUBS 0.006817f
C400 B.n300 VSUBS 0.006817f
C401 B.n301 VSUBS 0.006817f
C402 B.n302 VSUBS 0.006817f
C403 B.n303 VSUBS 0.006817f
C404 B.n304 VSUBS 0.006817f
C405 B.n305 VSUBS 0.006817f
C406 B.n306 VSUBS 0.006817f
C407 B.n307 VSUBS 0.006817f
C408 B.n308 VSUBS 0.006817f
C409 B.n309 VSUBS 0.006817f
C410 B.n310 VSUBS 0.006817f
C411 B.n311 VSUBS 0.006817f
C412 B.n312 VSUBS 0.006817f
C413 B.n313 VSUBS 0.006817f
C414 B.n314 VSUBS 0.006817f
C415 B.n315 VSUBS 0.006817f
C416 B.n316 VSUBS 0.006817f
C417 B.n317 VSUBS 0.006817f
C418 B.n318 VSUBS 0.006817f
C419 B.n319 VSUBS 0.006817f
C420 B.n320 VSUBS 0.006817f
C421 B.n321 VSUBS 0.006817f
C422 B.n322 VSUBS 0.006817f
C423 B.n323 VSUBS 0.006817f
C424 B.n324 VSUBS 0.006817f
C425 B.n325 VSUBS 0.006817f
C426 B.n326 VSUBS 0.006817f
C427 B.n327 VSUBS 0.006817f
C428 B.n328 VSUBS 0.006817f
C429 B.n329 VSUBS 0.006817f
C430 B.n330 VSUBS 0.006817f
C431 B.n331 VSUBS 0.006817f
C432 B.n332 VSUBS 0.006817f
C433 B.n333 VSUBS 0.006817f
C434 B.n334 VSUBS 0.006817f
C435 B.n335 VSUBS 0.006817f
C436 B.n336 VSUBS 0.006817f
C437 B.n337 VSUBS 0.006817f
C438 B.n338 VSUBS 0.006817f
C439 B.n339 VSUBS 0.006817f
C440 B.n340 VSUBS 0.006817f
C441 B.n341 VSUBS 0.006817f
C442 B.n342 VSUBS 0.006817f
C443 B.n343 VSUBS 0.006817f
C444 B.n344 VSUBS 0.006817f
C445 B.n345 VSUBS 0.006817f
C446 B.n346 VSUBS 0.006817f
C447 B.n347 VSUBS 0.006817f
C448 B.n348 VSUBS 0.006817f
C449 B.n349 VSUBS 0.006817f
C450 B.n350 VSUBS 0.006817f
C451 B.n351 VSUBS 0.006817f
C452 B.n352 VSUBS 0.006817f
C453 B.n353 VSUBS 0.006817f
C454 B.n354 VSUBS 0.006817f
C455 B.n355 VSUBS 0.006416f
C456 B.n356 VSUBS 0.015795f
C457 B.n357 VSUBS 0.00381f
C458 B.n358 VSUBS 0.006817f
C459 B.n359 VSUBS 0.006817f
C460 B.n360 VSUBS 0.006817f
C461 B.n361 VSUBS 0.006817f
C462 B.n362 VSUBS 0.006817f
C463 B.n363 VSUBS 0.006817f
C464 B.n364 VSUBS 0.006817f
C465 B.n365 VSUBS 0.006817f
C466 B.n366 VSUBS 0.006817f
C467 B.n367 VSUBS 0.006817f
C468 B.n368 VSUBS 0.006817f
C469 B.n369 VSUBS 0.006817f
C470 B.n370 VSUBS 0.00381f
C471 B.n371 VSUBS 0.006817f
C472 B.n372 VSUBS 0.006817f
C473 B.n373 VSUBS 0.006416f
C474 B.n374 VSUBS 0.006817f
C475 B.n375 VSUBS 0.006817f
C476 B.n376 VSUBS 0.006817f
C477 B.n377 VSUBS 0.006817f
C478 B.n378 VSUBS 0.006817f
C479 B.n379 VSUBS 0.006817f
C480 B.n380 VSUBS 0.006817f
C481 B.n381 VSUBS 0.006817f
C482 B.n382 VSUBS 0.006817f
C483 B.n383 VSUBS 0.006817f
C484 B.n384 VSUBS 0.006817f
C485 B.n385 VSUBS 0.006817f
C486 B.n386 VSUBS 0.006817f
C487 B.n387 VSUBS 0.006817f
C488 B.n388 VSUBS 0.006817f
C489 B.n389 VSUBS 0.006817f
C490 B.n390 VSUBS 0.006817f
C491 B.n391 VSUBS 0.006817f
C492 B.n392 VSUBS 0.006817f
C493 B.n393 VSUBS 0.006817f
C494 B.n394 VSUBS 0.006817f
C495 B.n395 VSUBS 0.006817f
C496 B.n396 VSUBS 0.006817f
C497 B.n397 VSUBS 0.006817f
C498 B.n398 VSUBS 0.006817f
C499 B.n399 VSUBS 0.006817f
C500 B.n400 VSUBS 0.006817f
C501 B.n401 VSUBS 0.006817f
C502 B.n402 VSUBS 0.006817f
C503 B.n403 VSUBS 0.006817f
C504 B.n404 VSUBS 0.006817f
C505 B.n405 VSUBS 0.006817f
C506 B.n406 VSUBS 0.006817f
C507 B.n407 VSUBS 0.006817f
C508 B.n408 VSUBS 0.006817f
C509 B.n409 VSUBS 0.006817f
C510 B.n410 VSUBS 0.006817f
C511 B.n411 VSUBS 0.006817f
C512 B.n412 VSUBS 0.006817f
C513 B.n413 VSUBS 0.006817f
C514 B.n414 VSUBS 0.006817f
C515 B.n415 VSUBS 0.006817f
C516 B.n416 VSUBS 0.006817f
C517 B.n417 VSUBS 0.006817f
C518 B.n418 VSUBS 0.006817f
C519 B.n419 VSUBS 0.006817f
C520 B.n420 VSUBS 0.006817f
C521 B.n421 VSUBS 0.006817f
C522 B.n422 VSUBS 0.006817f
C523 B.n423 VSUBS 0.006817f
C524 B.n424 VSUBS 0.006817f
C525 B.n425 VSUBS 0.006817f
C526 B.n426 VSUBS 0.006817f
C527 B.n427 VSUBS 0.006817f
C528 B.n428 VSUBS 0.006817f
C529 B.n429 VSUBS 0.006817f
C530 B.n430 VSUBS 0.006817f
C531 B.n431 VSUBS 0.006817f
C532 B.n432 VSUBS 0.006817f
C533 B.n433 VSUBS 0.006817f
C534 B.n434 VSUBS 0.006817f
C535 B.n435 VSUBS 0.006817f
C536 B.n436 VSUBS 0.006817f
C537 B.n437 VSUBS 0.006817f
C538 B.n438 VSUBS 0.006817f
C539 B.n439 VSUBS 0.006817f
C540 B.n440 VSUBS 0.006817f
C541 B.n441 VSUBS 0.006817f
C542 B.n442 VSUBS 0.006817f
C543 B.n443 VSUBS 0.006817f
C544 B.n444 VSUBS 0.006817f
C545 B.n445 VSUBS 0.006817f
C546 B.n446 VSUBS 0.006817f
C547 B.n447 VSUBS 0.006817f
C548 B.n448 VSUBS 0.006817f
C549 B.n449 VSUBS 0.006817f
C550 B.n450 VSUBS 0.006817f
C551 B.n451 VSUBS 0.006817f
C552 B.n452 VSUBS 0.006817f
C553 B.n453 VSUBS 0.006817f
C554 B.n454 VSUBS 0.006817f
C555 B.n455 VSUBS 0.006817f
C556 B.n456 VSUBS 0.006817f
C557 B.n457 VSUBS 0.006817f
C558 B.n458 VSUBS 0.006817f
C559 B.n459 VSUBS 0.006817f
C560 B.n460 VSUBS 0.006817f
C561 B.n461 VSUBS 0.006817f
C562 B.n462 VSUBS 0.016267f
C563 B.n463 VSUBS 0.016267f
C564 B.n464 VSUBS 0.015414f
C565 B.n465 VSUBS 0.006817f
C566 B.n466 VSUBS 0.006817f
C567 B.n467 VSUBS 0.006817f
C568 B.n468 VSUBS 0.006817f
C569 B.n469 VSUBS 0.006817f
C570 B.n470 VSUBS 0.006817f
C571 B.n471 VSUBS 0.006817f
C572 B.n472 VSUBS 0.006817f
C573 B.n473 VSUBS 0.006817f
C574 B.n474 VSUBS 0.006817f
C575 B.n475 VSUBS 0.006817f
C576 B.n476 VSUBS 0.006817f
C577 B.n477 VSUBS 0.006817f
C578 B.n478 VSUBS 0.006817f
C579 B.n479 VSUBS 0.006817f
C580 B.n480 VSUBS 0.006817f
C581 B.n481 VSUBS 0.006817f
C582 B.n482 VSUBS 0.006817f
C583 B.n483 VSUBS 0.006817f
C584 B.n484 VSUBS 0.006817f
C585 B.n485 VSUBS 0.006817f
C586 B.n486 VSUBS 0.006817f
C587 B.n487 VSUBS 0.006817f
C588 B.n488 VSUBS 0.006817f
C589 B.n489 VSUBS 0.006817f
C590 B.n490 VSUBS 0.006817f
C591 B.n491 VSUBS 0.006817f
C592 B.n492 VSUBS 0.006817f
C593 B.n493 VSUBS 0.006817f
C594 B.n494 VSUBS 0.006817f
C595 B.n495 VSUBS 0.006817f
C596 B.n496 VSUBS 0.006817f
C597 B.n497 VSUBS 0.006817f
C598 B.n498 VSUBS 0.006817f
C599 B.n499 VSUBS 0.006817f
C600 B.n500 VSUBS 0.006817f
C601 B.n501 VSUBS 0.006817f
C602 B.n502 VSUBS 0.006817f
C603 B.n503 VSUBS 0.006817f
C604 B.n504 VSUBS 0.006817f
C605 B.n505 VSUBS 0.006817f
C606 B.n506 VSUBS 0.006817f
C607 B.n507 VSUBS 0.006817f
C608 B.n508 VSUBS 0.006817f
C609 B.n509 VSUBS 0.006817f
C610 B.n510 VSUBS 0.006817f
C611 B.n511 VSUBS 0.006817f
C612 B.n512 VSUBS 0.006817f
C613 B.n513 VSUBS 0.006817f
C614 B.n514 VSUBS 0.006817f
C615 B.n515 VSUBS 0.006817f
C616 B.n516 VSUBS 0.006817f
C617 B.n517 VSUBS 0.006817f
C618 B.n518 VSUBS 0.006817f
C619 B.n519 VSUBS 0.006817f
C620 B.n520 VSUBS 0.006817f
C621 B.n521 VSUBS 0.006817f
C622 B.n522 VSUBS 0.006817f
C623 B.n523 VSUBS 0.006817f
C624 B.n524 VSUBS 0.006817f
C625 B.n525 VSUBS 0.006817f
C626 B.n526 VSUBS 0.006817f
C627 B.n527 VSUBS 0.006817f
C628 B.n528 VSUBS 0.006817f
C629 B.n529 VSUBS 0.006817f
C630 B.n530 VSUBS 0.006817f
C631 B.n531 VSUBS 0.006817f
C632 B.n532 VSUBS 0.006817f
C633 B.n533 VSUBS 0.006817f
C634 B.n534 VSUBS 0.006817f
C635 B.n535 VSUBS 0.006817f
C636 B.n536 VSUBS 0.006817f
C637 B.n537 VSUBS 0.006817f
C638 B.n538 VSUBS 0.006817f
C639 B.n539 VSUBS 0.006817f
C640 B.n540 VSUBS 0.006817f
C641 B.n541 VSUBS 0.006817f
C642 B.n542 VSUBS 0.006817f
C643 B.n543 VSUBS 0.006817f
C644 B.n544 VSUBS 0.006817f
C645 B.n545 VSUBS 0.006817f
C646 B.n546 VSUBS 0.006817f
C647 B.n547 VSUBS 0.006817f
C648 B.n548 VSUBS 0.006817f
C649 B.n549 VSUBS 0.006817f
C650 B.n550 VSUBS 0.006817f
C651 B.n551 VSUBS 0.006817f
C652 B.n552 VSUBS 0.006817f
C653 B.n553 VSUBS 0.006817f
C654 B.n554 VSUBS 0.006817f
C655 B.n555 VSUBS 0.006817f
C656 B.n556 VSUBS 0.006817f
C657 B.n557 VSUBS 0.006817f
C658 B.n558 VSUBS 0.006817f
C659 B.n559 VSUBS 0.006817f
C660 B.n560 VSUBS 0.006817f
C661 B.n561 VSUBS 0.006817f
C662 B.n562 VSUBS 0.006817f
C663 B.n563 VSUBS 0.006817f
C664 B.n564 VSUBS 0.006817f
C665 B.n565 VSUBS 0.006817f
C666 B.n566 VSUBS 0.006817f
C667 B.n567 VSUBS 0.006817f
C668 B.n568 VSUBS 0.006817f
C669 B.n569 VSUBS 0.015414f
C670 B.n570 VSUBS 0.016267f
C671 B.n571 VSUBS 0.015453f
C672 B.n572 VSUBS 0.006817f
C673 B.n573 VSUBS 0.006817f
C674 B.n574 VSUBS 0.006817f
C675 B.n575 VSUBS 0.006817f
C676 B.n576 VSUBS 0.006817f
C677 B.n577 VSUBS 0.006817f
C678 B.n578 VSUBS 0.006817f
C679 B.n579 VSUBS 0.006817f
C680 B.n580 VSUBS 0.006817f
C681 B.n581 VSUBS 0.006817f
C682 B.n582 VSUBS 0.006817f
C683 B.n583 VSUBS 0.006817f
C684 B.n584 VSUBS 0.006817f
C685 B.n585 VSUBS 0.006817f
C686 B.n586 VSUBS 0.006817f
C687 B.n587 VSUBS 0.006817f
C688 B.n588 VSUBS 0.006817f
C689 B.n589 VSUBS 0.006817f
C690 B.n590 VSUBS 0.006817f
C691 B.n591 VSUBS 0.006817f
C692 B.n592 VSUBS 0.006817f
C693 B.n593 VSUBS 0.006817f
C694 B.n594 VSUBS 0.006817f
C695 B.n595 VSUBS 0.006817f
C696 B.n596 VSUBS 0.006817f
C697 B.n597 VSUBS 0.006817f
C698 B.n598 VSUBS 0.006817f
C699 B.n599 VSUBS 0.006817f
C700 B.n600 VSUBS 0.006817f
C701 B.n601 VSUBS 0.006817f
C702 B.n602 VSUBS 0.006817f
C703 B.n603 VSUBS 0.006817f
C704 B.n604 VSUBS 0.006817f
C705 B.n605 VSUBS 0.006817f
C706 B.n606 VSUBS 0.006817f
C707 B.n607 VSUBS 0.006817f
C708 B.n608 VSUBS 0.006817f
C709 B.n609 VSUBS 0.006817f
C710 B.n610 VSUBS 0.006817f
C711 B.n611 VSUBS 0.006817f
C712 B.n612 VSUBS 0.006817f
C713 B.n613 VSUBS 0.006817f
C714 B.n614 VSUBS 0.006817f
C715 B.n615 VSUBS 0.006817f
C716 B.n616 VSUBS 0.006817f
C717 B.n617 VSUBS 0.006817f
C718 B.n618 VSUBS 0.006817f
C719 B.n619 VSUBS 0.006817f
C720 B.n620 VSUBS 0.006817f
C721 B.n621 VSUBS 0.006817f
C722 B.n622 VSUBS 0.006817f
C723 B.n623 VSUBS 0.006817f
C724 B.n624 VSUBS 0.006817f
C725 B.n625 VSUBS 0.006817f
C726 B.n626 VSUBS 0.006817f
C727 B.n627 VSUBS 0.006817f
C728 B.n628 VSUBS 0.006817f
C729 B.n629 VSUBS 0.006817f
C730 B.n630 VSUBS 0.006817f
C731 B.n631 VSUBS 0.006817f
C732 B.n632 VSUBS 0.006817f
C733 B.n633 VSUBS 0.006817f
C734 B.n634 VSUBS 0.006817f
C735 B.n635 VSUBS 0.006817f
C736 B.n636 VSUBS 0.006817f
C737 B.n637 VSUBS 0.006817f
C738 B.n638 VSUBS 0.006817f
C739 B.n639 VSUBS 0.006817f
C740 B.n640 VSUBS 0.006817f
C741 B.n641 VSUBS 0.006817f
C742 B.n642 VSUBS 0.006817f
C743 B.n643 VSUBS 0.006817f
C744 B.n644 VSUBS 0.006817f
C745 B.n645 VSUBS 0.006817f
C746 B.n646 VSUBS 0.006817f
C747 B.n647 VSUBS 0.006817f
C748 B.n648 VSUBS 0.006817f
C749 B.n649 VSUBS 0.006817f
C750 B.n650 VSUBS 0.006817f
C751 B.n651 VSUBS 0.006817f
C752 B.n652 VSUBS 0.006817f
C753 B.n653 VSUBS 0.006817f
C754 B.n654 VSUBS 0.006817f
C755 B.n655 VSUBS 0.006817f
C756 B.n656 VSUBS 0.006817f
C757 B.n657 VSUBS 0.006817f
C758 B.n658 VSUBS 0.006817f
C759 B.n659 VSUBS 0.006817f
C760 B.n660 VSUBS 0.006817f
C761 B.n661 VSUBS 0.006416f
C762 B.n662 VSUBS 0.015795f
C763 B.n663 VSUBS 0.00381f
C764 B.n664 VSUBS 0.006817f
C765 B.n665 VSUBS 0.006817f
C766 B.n666 VSUBS 0.006817f
C767 B.n667 VSUBS 0.006817f
C768 B.n668 VSUBS 0.006817f
C769 B.n669 VSUBS 0.006817f
C770 B.n670 VSUBS 0.006817f
C771 B.n671 VSUBS 0.006817f
C772 B.n672 VSUBS 0.006817f
C773 B.n673 VSUBS 0.006817f
C774 B.n674 VSUBS 0.006817f
C775 B.n675 VSUBS 0.006817f
C776 B.n676 VSUBS 0.00381f
C777 B.n677 VSUBS 0.006817f
C778 B.n678 VSUBS 0.006817f
C779 B.n679 VSUBS 0.006416f
C780 B.n680 VSUBS 0.006817f
C781 B.n681 VSUBS 0.006817f
C782 B.n682 VSUBS 0.006817f
C783 B.n683 VSUBS 0.006817f
C784 B.n684 VSUBS 0.006817f
C785 B.n685 VSUBS 0.006817f
C786 B.n686 VSUBS 0.006817f
C787 B.n687 VSUBS 0.006817f
C788 B.n688 VSUBS 0.006817f
C789 B.n689 VSUBS 0.006817f
C790 B.n690 VSUBS 0.006817f
C791 B.n691 VSUBS 0.006817f
C792 B.n692 VSUBS 0.006817f
C793 B.n693 VSUBS 0.006817f
C794 B.n694 VSUBS 0.006817f
C795 B.n695 VSUBS 0.006817f
C796 B.n696 VSUBS 0.006817f
C797 B.n697 VSUBS 0.006817f
C798 B.n698 VSUBS 0.006817f
C799 B.n699 VSUBS 0.006817f
C800 B.n700 VSUBS 0.006817f
C801 B.n701 VSUBS 0.006817f
C802 B.n702 VSUBS 0.006817f
C803 B.n703 VSUBS 0.006817f
C804 B.n704 VSUBS 0.006817f
C805 B.n705 VSUBS 0.006817f
C806 B.n706 VSUBS 0.006817f
C807 B.n707 VSUBS 0.006817f
C808 B.n708 VSUBS 0.006817f
C809 B.n709 VSUBS 0.006817f
C810 B.n710 VSUBS 0.006817f
C811 B.n711 VSUBS 0.006817f
C812 B.n712 VSUBS 0.006817f
C813 B.n713 VSUBS 0.006817f
C814 B.n714 VSUBS 0.006817f
C815 B.n715 VSUBS 0.006817f
C816 B.n716 VSUBS 0.006817f
C817 B.n717 VSUBS 0.006817f
C818 B.n718 VSUBS 0.006817f
C819 B.n719 VSUBS 0.006817f
C820 B.n720 VSUBS 0.006817f
C821 B.n721 VSUBS 0.006817f
C822 B.n722 VSUBS 0.006817f
C823 B.n723 VSUBS 0.006817f
C824 B.n724 VSUBS 0.006817f
C825 B.n725 VSUBS 0.006817f
C826 B.n726 VSUBS 0.006817f
C827 B.n727 VSUBS 0.006817f
C828 B.n728 VSUBS 0.006817f
C829 B.n729 VSUBS 0.006817f
C830 B.n730 VSUBS 0.006817f
C831 B.n731 VSUBS 0.006817f
C832 B.n732 VSUBS 0.006817f
C833 B.n733 VSUBS 0.006817f
C834 B.n734 VSUBS 0.006817f
C835 B.n735 VSUBS 0.006817f
C836 B.n736 VSUBS 0.006817f
C837 B.n737 VSUBS 0.006817f
C838 B.n738 VSUBS 0.006817f
C839 B.n739 VSUBS 0.006817f
C840 B.n740 VSUBS 0.006817f
C841 B.n741 VSUBS 0.006817f
C842 B.n742 VSUBS 0.006817f
C843 B.n743 VSUBS 0.006817f
C844 B.n744 VSUBS 0.006817f
C845 B.n745 VSUBS 0.006817f
C846 B.n746 VSUBS 0.006817f
C847 B.n747 VSUBS 0.006817f
C848 B.n748 VSUBS 0.006817f
C849 B.n749 VSUBS 0.006817f
C850 B.n750 VSUBS 0.006817f
C851 B.n751 VSUBS 0.006817f
C852 B.n752 VSUBS 0.006817f
C853 B.n753 VSUBS 0.006817f
C854 B.n754 VSUBS 0.006817f
C855 B.n755 VSUBS 0.006817f
C856 B.n756 VSUBS 0.006817f
C857 B.n757 VSUBS 0.006817f
C858 B.n758 VSUBS 0.006817f
C859 B.n759 VSUBS 0.006817f
C860 B.n760 VSUBS 0.006817f
C861 B.n761 VSUBS 0.006817f
C862 B.n762 VSUBS 0.006817f
C863 B.n763 VSUBS 0.006817f
C864 B.n764 VSUBS 0.006817f
C865 B.n765 VSUBS 0.006817f
C866 B.n766 VSUBS 0.006817f
C867 B.n767 VSUBS 0.006817f
C868 B.n768 VSUBS 0.016267f
C869 B.n769 VSUBS 0.016267f
C870 B.n770 VSUBS 0.015414f
C871 B.n771 VSUBS 0.006817f
C872 B.n772 VSUBS 0.006817f
C873 B.n773 VSUBS 0.006817f
C874 B.n774 VSUBS 0.006817f
C875 B.n775 VSUBS 0.006817f
C876 B.n776 VSUBS 0.006817f
C877 B.n777 VSUBS 0.006817f
C878 B.n778 VSUBS 0.006817f
C879 B.n779 VSUBS 0.006817f
C880 B.n780 VSUBS 0.006817f
C881 B.n781 VSUBS 0.006817f
C882 B.n782 VSUBS 0.006817f
C883 B.n783 VSUBS 0.006817f
C884 B.n784 VSUBS 0.006817f
C885 B.n785 VSUBS 0.006817f
C886 B.n786 VSUBS 0.006817f
C887 B.n787 VSUBS 0.006817f
C888 B.n788 VSUBS 0.006817f
C889 B.n789 VSUBS 0.006817f
C890 B.n790 VSUBS 0.006817f
C891 B.n791 VSUBS 0.006817f
C892 B.n792 VSUBS 0.006817f
C893 B.n793 VSUBS 0.006817f
C894 B.n794 VSUBS 0.006817f
C895 B.n795 VSUBS 0.006817f
C896 B.n796 VSUBS 0.006817f
C897 B.n797 VSUBS 0.006817f
C898 B.n798 VSUBS 0.006817f
C899 B.n799 VSUBS 0.006817f
C900 B.n800 VSUBS 0.006817f
C901 B.n801 VSUBS 0.006817f
C902 B.n802 VSUBS 0.006817f
C903 B.n803 VSUBS 0.006817f
C904 B.n804 VSUBS 0.006817f
C905 B.n805 VSUBS 0.006817f
C906 B.n806 VSUBS 0.006817f
C907 B.n807 VSUBS 0.006817f
C908 B.n808 VSUBS 0.006817f
C909 B.n809 VSUBS 0.006817f
C910 B.n810 VSUBS 0.006817f
C911 B.n811 VSUBS 0.006817f
C912 B.n812 VSUBS 0.006817f
C913 B.n813 VSUBS 0.006817f
C914 B.n814 VSUBS 0.006817f
C915 B.n815 VSUBS 0.006817f
C916 B.n816 VSUBS 0.006817f
C917 B.n817 VSUBS 0.006817f
C918 B.n818 VSUBS 0.006817f
C919 B.n819 VSUBS 0.006817f
C920 B.n820 VSUBS 0.006817f
C921 B.n821 VSUBS 0.006817f
C922 B.n822 VSUBS 0.006817f
C923 B.n823 VSUBS 0.015437f
C924 VTAIL.t6 VSUBS 0.339956f
C925 VTAIL.t1 VSUBS 0.339956f
C926 VTAIL.n0 VSUBS 2.69749f
C927 VTAIL.n1 VSUBS 0.686169f
C928 VTAIL.t2 VSUBS 3.51972f
C929 VTAIL.n2 VSUBS 0.821692f
C930 VTAIL.t11 VSUBS 3.51972f
C931 VTAIL.n3 VSUBS 0.821692f
C932 VTAIL.t10 VSUBS 0.339956f
C933 VTAIL.t12 VSUBS 0.339956f
C934 VTAIL.n4 VSUBS 2.69749f
C935 VTAIL.n5 VSUBS 0.799101f
C936 VTAIL.t15 VSUBS 3.51972f
C937 VTAIL.n6 VSUBS 2.41236f
C938 VTAIL.t5 VSUBS 3.51975f
C939 VTAIL.n7 VSUBS 2.41234f
C940 VTAIL.t0 VSUBS 0.339956f
C941 VTAIL.t4 VSUBS 0.339956f
C942 VTAIL.n8 VSUBS 2.6975f
C943 VTAIL.n9 VSUBS 0.799096f
C944 VTAIL.t3 VSUBS 3.51975f
C945 VTAIL.n10 VSUBS 0.821666f
C946 VTAIL.t13 VSUBS 3.51975f
C947 VTAIL.n11 VSUBS 0.821666f
C948 VTAIL.t14 VSUBS 0.339956f
C949 VTAIL.t8 VSUBS 0.339956f
C950 VTAIL.n12 VSUBS 2.6975f
C951 VTAIL.n13 VSUBS 0.799096f
C952 VTAIL.t9 VSUBS 3.51972f
C953 VTAIL.n14 VSUBS 2.41236f
C954 VTAIL.t7 VSUBS 3.51972f
C955 VTAIL.n15 VSUBS 2.40804f
C956 VDD1.t3 VSUBS 0.370621f
C957 VDD1.t4 VSUBS 0.370621f
C958 VDD1.n0 VSUBS 3.10403f
C959 VDD1.t5 VSUBS 0.370621f
C960 VDD1.t6 VSUBS 0.370621f
C961 VDD1.n1 VSUBS 3.10281f
C962 VDD1.t2 VSUBS 0.370621f
C963 VDD1.t7 VSUBS 0.370621f
C964 VDD1.n2 VSUBS 3.10281f
C965 VDD1.n3 VSUBS 3.69758f
C966 VDD1.t0 VSUBS 0.370621f
C967 VDD1.t1 VSUBS 0.370621f
C968 VDD1.n4 VSUBS 3.09557f
C969 VDD1.n5 VSUBS 3.41132f
C970 VP.n0 VSUBS 0.036184f
C971 VP.t4 VSUBS 2.78608f
C972 VP.n1 VSUBS 0.060888f
C973 VP.n2 VSUBS 0.036184f
C974 VP.t3 VSUBS 2.78608f
C975 VP.n3 VSUBS 0.066253f
C976 VP.n4 VSUBS 0.036184f
C977 VP.n5 VSUBS 0.050456f
C978 VP.n6 VSUBS 0.036184f
C979 VP.t6 VSUBS 2.78608f
C980 VP.n7 VSUBS 0.060888f
C981 VP.n8 VSUBS 0.036184f
C982 VP.t7 VSUBS 2.78608f
C983 VP.n9 VSUBS 0.066253f
C984 VP.t2 VSUBS 2.90251f
C985 VP.t1 VSUBS 2.78608f
C986 VP.n10 VSUBS 1.05766f
C987 VP.n11 VSUBS 1.06129f
C988 VP.n12 VSUBS 0.230073f
C989 VP.n13 VSUBS 0.036184f
C990 VP.n14 VSUBS 0.029251f
C991 VP.n15 VSUBS 0.066253f
C992 VP.n16 VSUBS 0.978884f
C993 VP.n17 VSUBS 0.039802f
C994 VP.n18 VSUBS 0.036184f
C995 VP.n19 VSUBS 0.036184f
C996 VP.n20 VSUBS 0.036184f
C997 VP.n21 VSUBS 0.044755f
C998 VP.n22 VSUBS 0.050456f
C999 VP.n23 VSUBS 1.05662f
C1000 VP.n24 VSUBS 2.01716f
C1001 VP.t0 VSUBS 2.78608f
C1002 VP.n25 VSUBS 1.05662f
C1003 VP.n26 VSUBS 2.04279f
C1004 VP.n27 VSUBS 0.036184f
C1005 VP.n28 VSUBS 0.036184f
C1006 VP.n29 VSUBS 0.044755f
C1007 VP.n30 VSUBS 0.060888f
C1008 VP.t5 VSUBS 2.78608f
C1009 VP.n31 VSUBS 0.978884f
C1010 VP.n32 VSUBS 0.039802f
C1011 VP.n33 VSUBS 0.036184f
C1012 VP.n34 VSUBS 0.036184f
C1013 VP.n35 VSUBS 0.036184f
C1014 VP.n36 VSUBS 0.029251f
C1015 VP.n37 VSUBS 0.066253f
C1016 VP.n38 VSUBS 0.978884f
C1017 VP.n39 VSUBS 0.039802f
C1018 VP.n40 VSUBS 0.036184f
C1019 VP.n41 VSUBS 0.036184f
C1020 VP.n42 VSUBS 0.036184f
C1021 VP.n43 VSUBS 0.044755f
C1022 VP.n44 VSUBS 0.050456f
C1023 VP.n45 VSUBS 1.05662f
C1024 VP.n46 VSUBS 0.034055f
.ends

