* NGSPICE file created from diff_pair_sample_0023.ext - technology: sky130A

.subckt diff_pair_sample_0023 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VN.t0 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=1.46
X1 VDD2.t4 VN.t1 VTAIL.t17 B.t8 sky130_fd_pr__nfet_01v8 ad=3.4281 pd=18.36 as=1.45035 ps=9.12 w=8.79 l=1.46
X2 VDD1.t9 VP.t0 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=3.4281 pd=18.36 as=1.45035 ps=9.12 w=8.79 l=1.46
X3 VDD2.t2 VN.t2 VTAIL.t16 B.t3 sky130_fd_pr__nfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=1.46
X4 VDD1.t8 VP.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.45035 pd=9.12 as=3.4281 ps=18.36 w=8.79 l=1.46
X5 B.t22 B.t20 B.t21 B.t17 sky130_fd_pr__nfet_01v8 ad=3.4281 pd=18.36 as=0 ps=0 w=8.79 l=1.46
X6 VDD2.t1 VN.t3 VTAIL.t15 B.t4 sky130_fd_pr__nfet_01v8 ad=1.45035 pd=9.12 as=3.4281 ps=18.36 w=8.79 l=1.46
X7 B.t19 B.t16 B.t18 B.t17 sky130_fd_pr__nfet_01v8 ad=3.4281 pd=18.36 as=0 ps=0 w=8.79 l=1.46
X8 VTAIL.t6 VP.t2 VDD1.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=1.46
X9 VDD2.t6 VN.t4 VTAIL.t14 B.t2 sky130_fd_pr__nfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=1.46
X10 VTAIL.t13 VN.t5 VDD2.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=1.46
X11 VTAIL.t1 VP.t3 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=1.46
X12 VTAIL.t0 VP.t4 VDD1.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=1.46
X13 VDD1.t4 VP.t5 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=3.4281 pd=18.36 as=1.45035 ps=9.12 w=8.79 l=1.46
X14 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=3.4281 pd=18.36 as=0 ps=0 w=8.79 l=1.46
X15 VDD1.t3 VP.t6 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.45035 pd=9.12 as=3.4281 ps=18.36 w=8.79 l=1.46
X16 VDD1.t2 VP.t7 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=1.46
X17 VTAIL.t19 VP.t8 VDD1.t1 B.t23 sky130_fd_pr__nfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=1.46
X18 VDD2.t9 VN.t6 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=1.45035 pd=9.12 as=3.4281 ps=18.36 w=8.79 l=1.46
X19 VTAIL.t11 VN.t7 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=1.46
X20 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=3.4281 pd=18.36 as=0 ps=0 w=8.79 l=1.46
X21 VDD1.t0 VP.t9 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=1.46
X22 VTAIL.t10 VN.t8 VDD2.t8 B.t23 sky130_fd_pr__nfet_01v8 ad=1.45035 pd=9.12 as=1.45035 ps=9.12 w=8.79 l=1.46
X23 VDD2.t7 VN.t9 VTAIL.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=3.4281 pd=18.36 as=1.45035 ps=9.12 w=8.79 l=1.46
R0 VN.n26 VN.n25 181.852
R1 VN.n53 VN.n52 181.852
R2 VN.n7 VN.t9 175.512
R3 VN.n34 VN.t6 175.512
R4 VN.n51 VN.n27 161.3
R5 VN.n50 VN.n49 161.3
R6 VN.n48 VN.n28 161.3
R7 VN.n47 VN.n46 161.3
R8 VN.n44 VN.n29 161.3
R9 VN.n43 VN.n42 161.3
R10 VN.n41 VN.n30 161.3
R11 VN.n40 VN.n39 161.3
R12 VN.n38 VN.n31 161.3
R13 VN.n37 VN.n36 161.3
R14 VN.n35 VN.n32 161.3
R15 VN.n24 VN.n0 161.3
R16 VN.n23 VN.n22 161.3
R17 VN.n21 VN.n1 161.3
R18 VN.n20 VN.n19 161.3
R19 VN.n17 VN.n2 161.3
R20 VN.n16 VN.n15 161.3
R21 VN.n14 VN.n3 161.3
R22 VN.n13 VN.n12 161.3
R23 VN.n11 VN.n4 161.3
R24 VN.n10 VN.n9 161.3
R25 VN.n8 VN.n5 161.3
R26 VN.n12 VN.t2 145.095
R27 VN.n6 VN.t7 145.095
R28 VN.n18 VN.t5 145.095
R29 VN.n25 VN.t3 145.095
R30 VN.n39 VN.t4 145.095
R31 VN.n33 VN.t0 145.095
R32 VN.n45 VN.t8 145.095
R33 VN.n52 VN.t1 145.095
R34 VN.n23 VN.n1 56.5193
R35 VN.n50 VN.n28 56.5193
R36 VN.n7 VN.n6 51.5804
R37 VN.n34 VN.n33 51.5804
R38 VN.n11 VN.n10 50.6917
R39 VN.n16 VN.n3 50.6917
R40 VN.n38 VN.n37 50.6917
R41 VN.n43 VN.n30 50.6917
R42 VN VN.n53 44.688
R43 VN.n10 VN.n5 30.2951
R44 VN.n17 VN.n16 30.2951
R45 VN.n37 VN.n32 30.2951
R46 VN.n44 VN.n43 30.2951
R47 VN.n12 VN.n11 24.4675
R48 VN.n12 VN.n3 24.4675
R49 VN.n19 VN.n1 24.4675
R50 VN.n24 VN.n23 24.4675
R51 VN.n39 VN.n30 24.4675
R52 VN.n39 VN.n38 24.4675
R53 VN.n46 VN.n28 24.4675
R54 VN.n51 VN.n50 24.4675
R55 VN.n35 VN.n34 18.3855
R56 VN.n8 VN.n7 18.3855
R57 VN.n6 VN.n5 14.1914
R58 VN.n18 VN.n17 14.1914
R59 VN.n33 VN.n32 14.1914
R60 VN.n45 VN.n44 14.1914
R61 VN.n19 VN.n18 10.2766
R62 VN.n46 VN.n45 10.2766
R63 VN.n25 VN.n24 3.91522
R64 VN.n52 VN.n51 3.91522
R65 VN.n53 VN.n27 0.189894
R66 VN.n49 VN.n27 0.189894
R67 VN.n49 VN.n48 0.189894
R68 VN.n48 VN.n47 0.189894
R69 VN.n47 VN.n29 0.189894
R70 VN.n42 VN.n29 0.189894
R71 VN.n42 VN.n41 0.189894
R72 VN.n41 VN.n40 0.189894
R73 VN.n40 VN.n31 0.189894
R74 VN.n36 VN.n31 0.189894
R75 VN.n36 VN.n35 0.189894
R76 VN.n9 VN.n8 0.189894
R77 VN.n9 VN.n4 0.189894
R78 VN.n13 VN.n4 0.189894
R79 VN.n14 VN.n13 0.189894
R80 VN.n15 VN.n14 0.189894
R81 VN.n15 VN.n2 0.189894
R82 VN.n20 VN.n2 0.189894
R83 VN.n21 VN.n20 0.189894
R84 VN.n22 VN.n21 0.189894
R85 VN.n22 VN.n0 0.189894
R86 VN.n26 VN.n0 0.189894
R87 VN VN.n26 0.0516364
R88 VDD2.n93 VDD2.n51 289.615
R89 VDD2.n42 VDD2.n0 289.615
R90 VDD2.n94 VDD2.n93 185
R91 VDD2.n92 VDD2.n91 185
R92 VDD2.n55 VDD2.n54 185
R93 VDD2.n86 VDD2.n85 185
R94 VDD2.n84 VDD2.n83 185
R95 VDD2.n59 VDD2.n58 185
R96 VDD2.n78 VDD2.n77 185
R97 VDD2.n76 VDD2.n75 185
R98 VDD2.n63 VDD2.n62 185
R99 VDD2.n70 VDD2.n69 185
R100 VDD2.n68 VDD2.n67 185
R101 VDD2.n17 VDD2.n16 185
R102 VDD2.n19 VDD2.n18 185
R103 VDD2.n12 VDD2.n11 185
R104 VDD2.n25 VDD2.n24 185
R105 VDD2.n27 VDD2.n26 185
R106 VDD2.n8 VDD2.n7 185
R107 VDD2.n33 VDD2.n32 185
R108 VDD2.n35 VDD2.n34 185
R109 VDD2.n4 VDD2.n3 185
R110 VDD2.n41 VDD2.n40 185
R111 VDD2.n43 VDD2.n42 185
R112 VDD2.n66 VDD2.t4 147.659
R113 VDD2.n15 VDD2.t7 147.659
R114 VDD2.n93 VDD2.n92 104.615
R115 VDD2.n92 VDD2.n54 104.615
R116 VDD2.n85 VDD2.n54 104.615
R117 VDD2.n85 VDD2.n84 104.615
R118 VDD2.n84 VDD2.n58 104.615
R119 VDD2.n77 VDD2.n58 104.615
R120 VDD2.n77 VDD2.n76 104.615
R121 VDD2.n76 VDD2.n62 104.615
R122 VDD2.n69 VDD2.n62 104.615
R123 VDD2.n69 VDD2.n68 104.615
R124 VDD2.n18 VDD2.n17 104.615
R125 VDD2.n18 VDD2.n11 104.615
R126 VDD2.n25 VDD2.n11 104.615
R127 VDD2.n26 VDD2.n25 104.615
R128 VDD2.n26 VDD2.n7 104.615
R129 VDD2.n33 VDD2.n7 104.615
R130 VDD2.n34 VDD2.n33 104.615
R131 VDD2.n34 VDD2.n3 104.615
R132 VDD2.n41 VDD2.n3 104.615
R133 VDD2.n42 VDD2.n41 104.615
R134 VDD2.n50 VDD2.n49 63.2945
R135 VDD2 VDD2.n101 63.2918
R136 VDD2.n100 VDD2.n99 62.1927
R137 VDD2.n48 VDD2.n47 62.1925
R138 VDD2.n68 VDD2.t4 52.3082
R139 VDD2.n17 VDD2.t7 52.3082
R140 VDD2.n48 VDD2.n46 48.6618
R141 VDD2.n98 VDD2.n97 47.1187
R142 VDD2.n98 VDD2.n50 38.6226
R143 VDD2.n67 VDD2.n66 15.6677
R144 VDD2.n16 VDD2.n15 15.6677
R145 VDD2.n70 VDD2.n65 12.8005
R146 VDD2.n19 VDD2.n14 12.8005
R147 VDD2.n71 VDD2.n63 12.0247
R148 VDD2.n20 VDD2.n12 12.0247
R149 VDD2.n75 VDD2.n74 11.249
R150 VDD2.n24 VDD2.n23 11.249
R151 VDD2.n78 VDD2.n61 10.4732
R152 VDD2.n27 VDD2.n10 10.4732
R153 VDD2.n79 VDD2.n59 9.69747
R154 VDD2.n28 VDD2.n8 9.69747
R155 VDD2.n97 VDD2.n96 9.45567
R156 VDD2.n46 VDD2.n45 9.45567
R157 VDD2.n53 VDD2.n52 9.3005
R158 VDD2.n96 VDD2.n95 9.3005
R159 VDD2.n90 VDD2.n89 9.3005
R160 VDD2.n88 VDD2.n87 9.3005
R161 VDD2.n57 VDD2.n56 9.3005
R162 VDD2.n82 VDD2.n81 9.3005
R163 VDD2.n80 VDD2.n79 9.3005
R164 VDD2.n61 VDD2.n60 9.3005
R165 VDD2.n74 VDD2.n73 9.3005
R166 VDD2.n72 VDD2.n71 9.3005
R167 VDD2.n65 VDD2.n64 9.3005
R168 VDD2.n39 VDD2.n38 9.3005
R169 VDD2.n2 VDD2.n1 9.3005
R170 VDD2.n45 VDD2.n44 9.3005
R171 VDD2.n6 VDD2.n5 9.3005
R172 VDD2.n31 VDD2.n30 9.3005
R173 VDD2.n29 VDD2.n28 9.3005
R174 VDD2.n10 VDD2.n9 9.3005
R175 VDD2.n23 VDD2.n22 9.3005
R176 VDD2.n21 VDD2.n20 9.3005
R177 VDD2.n14 VDD2.n13 9.3005
R178 VDD2.n37 VDD2.n36 9.3005
R179 VDD2.n97 VDD2.n51 8.92171
R180 VDD2.n83 VDD2.n82 8.92171
R181 VDD2.n32 VDD2.n31 8.92171
R182 VDD2.n46 VDD2.n0 8.92171
R183 VDD2.n95 VDD2.n94 8.14595
R184 VDD2.n86 VDD2.n57 8.14595
R185 VDD2.n35 VDD2.n6 8.14595
R186 VDD2.n44 VDD2.n43 8.14595
R187 VDD2.n91 VDD2.n53 7.3702
R188 VDD2.n87 VDD2.n55 7.3702
R189 VDD2.n36 VDD2.n4 7.3702
R190 VDD2.n40 VDD2.n2 7.3702
R191 VDD2.n91 VDD2.n90 6.59444
R192 VDD2.n90 VDD2.n55 6.59444
R193 VDD2.n39 VDD2.n4 6.59444
R194 VDD2.n40 VDD2.n39 6.59444
R195 VDD2.n94 VDD2.n53 5.81868
R196 VDD2.n87 VDD2.n86 5.81868
R197 VDD2.n36 VDD2.n35 5.81868
R198 VDD2.n43 VDD2.n2 5.81868
R199 VDD2.n95 VDD2.n51 5.04292
R200 VDD2.n83 VDD2.n57 5.04292
R201 VDD2.n32 VDD2.n6 5.04292
R202 VDD2.n44 VDD2.n0 5.04292
R203 VDD2.n66 VDD2.n64 4.38563
R204 VDD2.n15 VDD2.n13 4.38563
R205 VDD2.n82 VDD2.n59 4.26717
R206 VDD2.n31 VDD2.n8 4.26717
R207 VDD2.n79 VDD2.n78 3.49141
R208 VDD2.n28 VDD2.n27 3.49141
R209 VDD2.n75 VDD2.n61 2.71565
R210 VDD2.n24 VDD2.n10 2.71565
R211 VDD2.n101 VDD2.t3 2.25306
R212 VDD2.n101 VDD2.t9 2.25306
R213 VDD2.n99 VDD2.t8 2.25306
R214 VDD2.n99 VDD2.t6 2.25306
R215 VDD2.n49 VDD2.t0 2.25306
R216 VDD2.n49 VDD2.t1 2.25306
R217 VDD2.n47 VDD2.t5 2.25306
R218 VDD2.n47 VDD2.t2 2.25306
R219 VDD2.n74 VDD2.n63 1.93989
R220 VDD2.n23 VDD2.n12 1.93989
R221 VDD2.n100 VDD2.n98 1.5436
R222 VDD2.n71 VDD2.n70 1.16414
R223 VDD2.n20 VDD2.n19 1.16414
R224 VDD2 VDD2.n100 0.444466
R225 VDD2.n67 VDD2.n65 0.388379
R226 VDD2.n16 VDD2.n14 0.388379
R227 VDD2.n50 VDD2.n48 0.33093
R228 VDD2.n96 VDD2.n52 0.155672
R229 VDD2.n89 VDD2.n52 0.155672
R230 VDD2.n89 VDD2.n88 0.155672
R231 VDD2.n88 VDD2.n56 0.155672
R232 VDD2.n81 VDD2.n56 0.155672
R233 VDD2.n81 VDD2.n80 0.155672
R234 VDD2.n80 VDD2.n60 0.155672
R235 VDD2.n73 VDD2.n60 0.155672
R236 VDD2.n73 VDD2.n72 0.155672
R237 VDD2.n72 VDD2.n64 0.155672
R238 VDD2.n21 VDD2.n13 0.155672
R239 VDD2.n22 VDD2.n21 0.155672
R240 VDD2.n22 VDD2.n9 0.155672
R241 VDD2.n29 VDD2.n9 0.155672
R242 VDD2.n30 VDD2.n29 0.155672
R243 VDD2.n30 VDD2.n5 0.155672
R244 VDD2.n37 VDD2.n5 0.155672
R245 VDD2.n38 VDD2.n37 0.155672
R246 VDD2.n38 VDD2.n1 0.155672
R247 VDD2.n45 VDD2.n1 0.155672
R248 VTAIL.n200 VTAIL.n158 289.615
R249 VTAIL.n44 VTAIL.n2 289.615
R250 VTAIL.n152 VTAIL.n110 289.615
R251 VTAIL.n100 VTAIL.n58 289.615
R252 VTAIL.n175 VTAIL.n174 185
R253 VTAIL.n177 VTAIL.n176 185
R254 VTAIL.n170 VTAIL.n169 185
R255 VTAIL.n183 VTAIL.n182 185
R256 VTAIL.n185 VTAIL.n184 185
R257 VTAIL.n166 VTAIL.n165 185
R258 VTAIL.n191 VTAIL.n190 185
R259 VTAIL.n193 VTAIL.n192 185
R260 VTAIL.n162 VTAIL.n161 185
R261 VTAIL.n199 VTAIL.n198 185
R262 VTAIL.n201 VTAIL.n200 185
R263 VTAIL.n19 VTAIL.n18 185
R264 VTAIL.n21 VTAIL.n20 185
R265 VTAIL.n14 VTAIL.n13 185
R266 VTAIL.n27 VTAIL.n26 185
R267 VTAIL.n29 VTAIL.n28 185
R268 VTAIL.n10 VTAIL.n9 185
R269 VTAIL.n35 VTAIL.n34 185
R270 VTAIL.n37 VTAIL.n36 185
R271 VTAIL.n6 VTAIL.n5 185
R272 VTAIL.n43 VTAIL.n42 185
R273 VTAIL.n45 VTAIL.n44 185
R274 VTAIL.n153 VTAIL.n152 185
R275 VTAIL.n151 VTAIL.n150 185
R276 VTAIL.n114 VTAIL.n113 185
R277 VTAIL.n145 VTAIL.n144 185
R278 VTAIL.n143 VTAIL.n142 185
R279 VTAIL.n118 VTAIL.n117 185
R280 VTAIL.n137 VTAIL.n136 185
R281 VTAIL.n135 VTAIL.n134 185
R282 VTAIL.n122 VTAIL.n121 185
R283 VTAIL.n129 VTAIL.n128 185
R284 VTAIL.n127 VTAIL.n126 185
R285 VTAIL.n101 VTAIL.n100 185
R286 VTAIL.n99 VTAIL.n98 185
R287 VTAIL.n62 VTAIL.n61 185
R288 VTAIL.n93 VTAIL.n92 185
R289 VTAIL.n91 VTAIL.n90 185
R290 VTAIL.n66 VTAIL.n65 185
R291 VTAIL.n85 VTAIL.n84 185
R292 VTAIL.n83 VTAIL.n82 185
R293 VTAIL.n70 VTAIL.n69 185
R294 VTAIL.n77 VTAIL.n76 185
R295 VTAIL.n75 VTAIL.n74 185
R296 VTAIL.n73 VTAIL.t12 147.659
R297 VTAIL.n173 VTAIL.t15 147.659
R298 VTAIL.n17 VTAIL.t5 147.659
R299 VTAIL.n125 VTAIL.t4 147.659
R300 VTAIL.n176 VTAIL.n175 104.615
R301 VTAIL.n176 VTAIL.n169 104.615
R302 VTAIL.n183 VTAIL.n169 104.615
R303 VTAIL.n184 VTAIL.n183 104.615
R304 VTAIL.n184 VTAIL.n165 104.615
R305 VTAIL.n191 VTAIL.n165 104.615
R306 VTAIL.n192 VTAIL.n191 104.615
R307 VTAIL.n192 VTAIL.n161 104.615
R308 VTAIL.n199 VTAIL.n161 104.615
R309 VTAIL.n200 VTAIL.n199 104.615
R310 VTAIL.n20 VTAIL.n19 104.615
R311 VTAIL.n20 VTAIL.n13 104.615
R312 VTAIL.n27 VTAIL.n13 104.615
R313 VTAIL.n28 VTAIL.n27 104.615
R314 VTAIL.n28 VTAIL.n9 104.615
R315 VTAIL.n35 VTAIL.n9 104.615
R316 VTAIL.n36 VTAIL.n35 104.615
R317 VTAIL.n36 VTAIL.n5 104.615
R318 VTAIL.n43 VTAIL.n5 104.615
R319 VTAIL.n44 VTAIL.n43 104.615
R320 VTAIL.n152 VTAIL.n151 104.615
R321 VTAIL.n151 VTAIL.n113 104.615
R322 VTAIL.n144 VTAIL.n113 104.615
R323 VTAIL.n144 VTAIL.n143 104.615
R324 VTAIL.n143 VTAIL.n117 104.615
R325 VTAIL.n136 VTAIL.n117 104.615
R326 VTAIL.n136 VTAIL.n135 104.615
R327 VTAIL.n135 VTAIL.n121 104.615
R328 VTAIL.n128 VTAIL.n121 104.615
R329 VTAIL.n128 VTAIL.n127 104.615
R330 VTAIL.n100 VTAIL.n99 104.615
R331 VTAIL.n99 VTAIL.n61 104.615
R332 VTAIL.n92 VTAIL.n61 104.615
R333 VTAIL.n92 VTAIL.n91 104.615
R334 VTAIL.n91 VTAIL.n65 104.615
R335 VTAIL.n84 VTAIL.n65 104.615
R336 VTAIL.n84 VTAIL.n83 104.615
R337 VTAIL.n83 VTAIL.n69 104.615
R338 VTAIL.n76 VTAIL.n69 104.615
R339 VTAIL.n76 VTAIL.n75 104.615
R340 VTAIL.n175 VTAIL.t15 52.3082
R341 VTAIL.n19 VTAIL.t5 52.3082
R342 VTAIL.n127 VTAIL.t4 52.3082
R343 VTAIL.n75 VTAIL.t12 52.3082
R344 VTAIL.n109 VTAIL.n108 45.5139
R345 VTAIL.n107 VTAIL.n106 45.5139
R346 VTAIL.n57 VTAIL.n56 45.5139
R347 VTAIL.n55 VTAIL.n54 45.5139
R348 VTAIL.n207 VTAIL.n206 45.5137
R349 VTAIL.n1 VTAIL.n0 45.5137
R350 VTAIL.n51 VTAIL.n50 45.5137
R351 VTAIL.n53 VTAIL.n52 45.5137
R352 VTAIL.n205 VTAIL.n204 30.4399
R353 VTAIL.n49 VTAIL.n48 30.4399
R354 VTAIL.n157 VTAIL.n156 30.4399
R355 VTAIL.n105 VTAIL.n104 30.4399
R356 VTAIL.n55 VTAIL.n53 23.0307
R357 VTAIL.n205 VTAIL.n157 21.4876
R358 VTAIL.n174 VTAIL.n173 15.6677
R359 VTAIL.n18 VTAIL.n17 15.6677
R360 VTAIL.n126 VTAIL.n125 15.6677
R361 VTAIL.n74 VTAIL.n73 15.6677
R362 VTAIL.n177 VTAIL.n172 12.8005
R363 VTAIL.n21 VTAIL.n16 12.8005
R364 VTAIL.n129 VTAIL.n124 12.8005
R365 VTAIL.n77 VTAIL.n72 12.8005
R366 VTAIL.n178 VTAIL.n170 12.0247
R367 VTAIL.n22 VTAIL.n14 12.0247
R368 VTAIL.n130 VTAIL.n122 12.0247
R369 VTAIL.n78 VTAIL.n70 12.0247
R370 VTAIL.n182 VTAIL.n181 11.249
R371 VTAIL.n26 VTAIL.n25 11.249
R372 VTAIL.n134 VTAIL.n133 11.249
R373 VTAIL.n82 VTAIL.n81 11.249
R374 VTAIL.n185 VTAIL.n168 10.4732
R375 VTAIL.n29 VTAIL.n12 10.4732
R376 VTAIL.n137 VTAIL.n120 10.4732
R377 VTAIL.n85 VTAIL.n68 10.4732
R378 VTAIL.n186 VTAIL.n166 9.69747
R379 VTAIL.n30 VTAIL.n10 9.69747
R380 VTAIL.n138 VTAIL.n118 9.69747
R381 VTAIL.n86 VTAIL.n66 9.69747
R382 VTAIL.n204 VTAIL.n203 9.45567
R383 VTAIL.n48 VTAIL.n47 9.45567
R384 VTAIL.n156 VTAIL.n155 9.45567
R385 VTAIL.n104 VTAIL.n103 9.45567
R386 VTAIL.n197 VTAIL.n196 9.3005
R387 VTAIL.n160 VTAIL.n159 9.3005
R388 VTAIL.n203 VTAIL.n202 9.3005
R389 VTAIL.n164 VTAIL.n163 9.3005
R390 VTAIL.n189 VTAIL.n188 9.3005
R391 VTAIL.n187 VTAIL.n186 9.3005
R392 VTAIL.n168 VTAIL.n167 9.3005
R393 VTAIL.n181 VTAIL.n180 9.3005
R394 VTAIL.n179 VTAIL.n178 9.3005
R395 VTAIL.n172 VTAIL.n171 9.3005
R396 VTAIL.n195 VTAIL.n194 9.3005
R397 VTAIL.n41 VTAIL.n40 9.3005
R398 VTAIL.n4 VTAIL.n3 9.3005
R399 VTAIL.n47 VTAIL.n46 9.3005
R400 VTAIL.n8 VTAIL.n7 9.3005
R401 VTAIL.n33 VTAIL.n32 9.3005
R402 VTAIL.n31 VTAIL.n30 9.3005
R403 VTAIL.n12 VTAIL.n11 9.3005
R404 VTAIL.n25 VTAIL.n24 9.3005
R405 VTAIL.n23 VTAIL.n22 9.3005
R406 VTAIL.n16 VTAIL.n15 9.3005
R407 VTAIL.n39 VTAIL.n38 9.3005
R408 VTAIL.n112 VTAIL.n111 9.3005
R409 VTAIL.n149 VTAIL.n148 9.3005
R410 VTAIL.n147 VTAIL.n146 9.3005
R411 VTAIL.n116 VTAIL.n115 9.3005
R412 VTAIL.n141 VTAIL.n140 9.3005
R413 VTAIL.n139 VTAIL.n138 9.3005
R414 VTAIL.n120 VTAIL.n119 9.3005
R415 VTAIL.n133 VTAIL.n132 9.3005
R416 VTAIL.n131 VTAIL.n130 9.3005
R417 VTAIL.n124 VTAIL.n123 9.3005
R418 VTAIL.n155 VTAIL.n154 9.3005
R419 VTAIL.n60 VTAIL.n59 9.3005
R420 VTAIL.n103 VTAIL.n102 9.3005
R421 VTAIL.n97 VTAIL.n96 9.3005
R422 VTAIL.n95 VTAIL.n94 9.3005
R423 VTAIL.n64 VTAIL.n63 9.3005
R424 VTAIL.n89 VTAIL.n88 9.3005
R425 VTAIL.n87 VTAIL.n86 9.3005
R426 VTAIL.n68 VTAIL.n67 9.3005
R427 VTAIL.n81 VTAIL.n80 9.3005
R428 VTAIL.n79 VTAIL.n78 9.3005
R429 VTAIL.n72 VTAIL.n71 9.3005
R430 VTAIL.n190 VTAIL.n189 8.92171
R431 VTAIL.n204 VTAIL.n158 8.92171
R432 VTAIL.n34 VTAIL.n33 8.92171
R433 VTAIL.n48 VTAIL.n2 8.92171
R434 VTAIL.n156 VTAIL.n110 8.92171
R435 VTAIL.n142 VTAIL.n141 8.92171
R436 VTAIL.n104 VTAIL.n58 8.92171
R437 VTAIL.n90 VTAIL.n89 8.92171
R438 VTAIL.n193 VTAIL.n164 8.14595
R439 VTAIL.n202 VTAIL.n201 8.14595
R440 VTAIL.n37 VTAIL.n8 8.14595
R441 VTAIL.n46 VTAIL.n45 8.14595
R442 VTAIL.n154 VTAIL.n153 8.14595
R443 VTAIL.n145 VTAIL.n116 8.14595
R444 VTAIL.n102 VTAIL.n101 8.14595
R445 VTAIL.n93 VTAIL.n64 8.14595
R446 VTAIL.n194 VTAIL.n162 7.3702
R447 VTAIL.n198 VTAIL.n160 7.3702
R448 VTAIL.n38 VTAIL.n6 7.3702
R449 VTAIL.n42 VTAIL.n4 7.3702
R450 VTAIL.n150 VTAIL.n112 7.3702
R451 VTAIL.n146 VTAIL.n114 7.3702
R452 VTAIL.n98 VTAIL.n60 7.3702
R453 VTAIL.n94 VTAIL.n62 7.3702
R454 VTAIL.n197 VTAIL.n162 6.59444
R455 VTAIL.n198 VTAIL.n197 6.59444
R456 VTAIL.n41 VTAIL.n6 6.59444
R457 VTAIL.n42 VTAIL.n41 6.59444
R458 VTAIL.n150 VTAIL.n149 6.59444
R459 VTAIL.n149 VTAIL.n114 6.59444
R460 VTAIL.n98 VTAIL.n97 6.59444
R461 VTAIL.n97 VTAIL.n62 6.59444
R462 VTAIL.n194 VTAIL.n193 5.81868
R463 VTAIL.n201 VTAIL.n160 5.81868
R464 VTAIL.n38 VTAIL.n37 5.81868
R465 VTAIL.n45 VTAIL.n4 5.81868
R466 VTAIL.n153 VTAIL.n112 5.81868
R467 VTAIL.n146 VTAIL.n145 5.81868
R468 VTAIL.n101 VTAIL.n60 5.81868
R469 VTAIL.n94 VTAIL.n93 5.81868
R470 VTAIL.n190 VTAIL.n164 5.04292
R471 VTAIL.n202 VTAIL.n158 5.04292
R472 VTAIL.n34 VTAIL.n8 5.04292
R473 VTAIL.n46 VTAIL.n2 5.04292
R474 VTAIL.n154 VTAIL.n110 5.04292
R475 VTAIL.n142 VTAIL.n116 5.04292
R476 VTAIL.n102 VTAIL.n58 5.04292
R477 VTAIL.n90 VTAIL.n64 5.04292
R478 VTAIL.n173 VTAIL.n171 4.38563
R479 VTAIL.n17 VTAIL.n15 4.38563
R480 VTAIL.n125 VTAIL.n123 4.38563
R481 VTAIL.n73 VTAIL.n71 4.38563
R482 VTAIL.n189 VTAIL.n166 4.26717
R483 VTAIL.n33 VTAIL.n10 4.26717
R484 VTAIL.n141 VTAIL.n118 4.26717
R485 VTAIL.n89 VTAIL.n66 4.26717
R486 VTAIL.n186 VTAIL.n185 3.49141
R487 VTAIL.n30 VTAIL.n29 3.49141
R488 VTAIL.n138 VTAIL.n137 3.49141
R489 VTAIL.n86 VTAIL.n85 3.49141
R490 VTAIL.n182 VTAIL.n168 2.71565
R491 VTAIL.n26 VTAIL.n12 2.71565
R492 VTAIL.n134 VTAIL.n120 2.71565
R493 VTAIL.n82 VTAIL.n68 2.71565
R494 VTAIL.n206 VTAIL.t16 2.25306
R495 VTAIL.n206 VTAIL.t13 2.25306
R496 VTAIL.n0 VTAIL.t9 2.25306
R497 VTAIL.n0 VTAIL.t11 2.25306
R498 VTAIL.n50 VTAIL.t2 2.25306
R499 VTAIL.n50 VTAIL.t0 2.25306
R500 VTAIL.n52 VTAIL.t8 2.25306
R501 VTAIL.n52 VTAIL.t19 2.25306
R502 VTAIL.n108 VTAIL.t3 2.25306
R503 VTAIL.n108 VTAIL.t6 2.25306
R504 VTAIL.n106 VTAIL.t7 2.25306
R505 VTAIL.n106 VTAIL.t1 2.25306
R506 VTAIL.n56 VTAIL.t14 2.25306
R507 VTAIL.n56 VTAIL.t18 2.25306
R508 VTAIL.n54 VTAIL.t17 2.25306
R509 VTAIL.n54 VTAIL.t10 2.25306
R510 VTAIL.n181 VTAIL.n170 1.93989
R511 VTAIL.n25 VTAIL.n14 1.93989
R512 VTAIL.n133 VTAIL.n122 1.93989
R513 VTAIL.n81 VTAIL.n70 1.93989
R514 VTAIL.n57 VTAIL.n55 1.5436
R515 VTAIL.n105 VTAIL.n57 1.5436
R516 VTAIL.n109 VTAIL.n107 1.5436
R517 VTAIL.n157 VTAIL.n109 1.5436
R518 VTAIL.n53 VTAIL.n51 1.5436
R519 VTAIL.n51 VTAIL.n49 1.5436
R520 VTAIL.n207 VTAIL.n205 1.5436
R521 VTAIL.n107 VTAIL.n105 1.24188
R522 VTAIL.n49 VTAIL.n1 1.24188
R523 VTAIL VTAIL.n1 1.21602
R524 VTAIL.n178 VTAIL.n177 1.16414
R525 VTAIL.n22 VTAIL.n21 1.16414
R526 VTAIL.n130 VTAIL.n129 1.16414
R527 VTAIL.n78 VTAIL.n77 1.16414
R528 VTAIL.n174 VTAIL.n172 0.388379
R529 VTAIL.n18 VTAIL.n16 0.388379
R530 VTAIL.n126 VTAIL.n124 0.388379
R531 VTAIL.n74 VTAIL.n72 0.388379
R532 VTAIL VTAIL.n207 0.328086
R533 VTAIL.n179 VTAIL.n171 0.155672
R534 VTAIL.n180 VTAIL.n179 0.155672
R535 VTAIL.n180 VTAIL.n167 0.155672
R536 VTAIL.n187 VTAIL.n167 0.155672
R537 VTAIL.n188 VTAIL.n187 0.155672
R538 VTAIL.n188 VTAIL.n163 0.155672
R539 VTAIL.n195 VTAIL.n163 0.155672
R540 VTAIL.n196 VTAIL.n195 0.155672
R541 VTAIL.n196 VTAIL.n159 0.155672
R542 VTAIL.n203 VTAIL.n159 0.155672
R543 VTAIL.n23 VTAIL.n15 0.155672
R544 VTAIL.n24 VTAIL.n23 0.155672
R545 VTAIL.n24 VTAIL.n11 0.155672
R546 VTAIL.n31 VTAIL.n11 0.155672
R547 VTAIL.n32 VTAIL.n31 0.155672
R548 VTAIL.n32 VTAIL.n7 0.155672
R549 VTAIL.n39 VTAIL.n7 0.155672
R550 VTAIL.n40 VTAIL.n39 0.155672
R551 VTAIL.n40 VTAIL.n3 0.155672
R552 VTAIL.n47 VTAIL.n3 0.155672
R553 VTAIL.n155 VTAIL.n111 0.155672
R554 VTAIL.n148 VTAIL.n111 0.155672
R555 VTAIL.n148 VTAIL.n147 0.155672
R556 VTAIL.n147 VTAIL.n115 0.155672
R557 VTAIL.n140 VTAIL.n115 0.155672
R558 VTAIL.n140 VTAIL.n139 0.155672
R559 VTAIL.n139 VTAIL.n119 0.155672
R560 VTAIL.n132 VTAIL.n119 0.155672
R561 VTAIL.n132 VTAIL.n131 0.155672
R562 VTAIL.n131 VTAIL.n123 0.155672
R563 VTAIL.n103 VTAIL.n59 0.155672
R564 VTAIL.n96 VTAIL.n59 0.155672
R565 VTAIL.n96 VTAIL.n95 0.155672
R566 VTAIL.n95 VTAIL.n63 0.155672
R567 VTAIL.n88 VTAIL.n63 0.155672
R568 VTAIL.n88 VTAIL.n87 0.155672
R569 VTAIL.n87 VTAIL.n67 0.155672
R570 VTAIL.n80 VTAIL.n67 0.155672
R571 VTAIL.n80 VTAIL.n79 0.155672
R572 VTAIL.n79 VTAIL.n71 0.155672
R573 B.n694 B.n693 585
R574 B.n258 B.n110 585
R575 B.n257 B.n256 585
R576 B.n255 B.n254 585
R577 B.n253 B.n252 585
R578 B.n251 B.n250 585
R579 B.n249 B.n248 585
R580 B.n247 B.n246 585
R581 B.n245 B.n244 585
R582 B.n243 B.n242 585
R583 B.n241 B.n240 585
R584 B.n239 B.n238 585
R585 B.n237 B.n236 585
R586 B.n235 B.n234 585
R587 B.n233 B.n232 585
R588 B.n231 B.n230 585
R589 B.n229 B.n228 585
R590 B.n227 B.n226 585
R591 B.n225 B.n224 585
R592 B.n223 B.n222 585
R593 B.n221 B.n220 585
R594 B.n219 B.n218 585
R595 B.n217 B.n216 585
R596 B.n215 B.n214 585
R597 B.n213 B.n212 585
R598 B.n211 B.n210 585
R599 B.n209 B.n208 585
R600 B.n207 B.n206 585
R601 B.n205 B.n204 585
R602 B.n203 B.n202 585
R603 B.n201 B.n200 585
R604 B.n199 B.n198 585
R605 B.n197 B.n196 585
R606 B.n195 B.n194 585
R607 B.n193 B.n192 585
R608 B.n191 B.n190 585
R609 B.n189 B.n188 585
R610 B.n187 B.n186 585
R611 B.n185 B.n184 585
R612 B.n183 B.n182 585
R613 B.n181 B.n180 585
R614 B.n179 B.n178 585
R615 B.n177 B.n176 585
R616 B.n175 B.n174 585
R617 B.n173 B.n172 585
R618 B.n171 B.n170 585
R619 B.n169 B.n168 585
R620 B.n167 B.n166 585
R621 B.n165 B.n164 585
R622 B.n163 B.n162 585
R623 B.n161 B.n160 585
R624 B.n159 B.n158 585
R625 B.n157 B.n156 585
R626 B.n155 B.n154 585
R627 B.n153 B.n152 585
R628 B.n151 B.n150 585
R629 B.n149 B.n148 585
R630 B.n147 B.n146 585
R631 B.n145 B.n144 585
R632 B.n143 B.n142 585
R633 B.n141 B.n140 585
R634 B.n139 B.n138 585
R635 B.n137 B.n136 585
R636 B.n135 B.n134 585
R637 B.n133 B.n132 585
R638 B.n131 B.n130 585
R639 B.n129 B.n128 585
R640 B.n127 B.n126 585
R641 B.n125 B.n124 585
R642 B.n123 B.n122 585
R643 B.n121 B.n120 585
R644 B.n119 B.n118 585
R645 B.n74 B.n73 585
R646 B.n699 B.n698 585
R647 B.n692 B.n111 585
R648 B.n111 B.n71 585
R649 B.n691 B.n70 585
R650 B.n703 B.n70 585
R651 B.n690 B.n69 585
R652 B.n704 B.n69 585
R653 B.n689 B.n68 585
R654 B.n705 B.n68 585
R655 B.n688 B.n687 585
R656 B.n687 B.n64 585
R657 B.n686 B.n63 585
R658 B.n711 B.n63 585
R659 B.n685 B.n62 585
R660 B.n712 B.n62 585
R661 B.n684 B.n61 585
R662 B.n713 B.n61 585
R663 B.n683 B.n682 585
R664 B.n682 B.n57 585
R665 B.n681 B.n56 585
R666 B.n719 B.n56 585
R667 B.n680 B.n55 585
R668 B.n720 B.n55 585
R669 B.n679 B.n54 585
R670 B.n721 B.n54 585
R671 B.n678 B.n677 585
R672 B.n677 B.n50 585
R673 B.n676 B.n49 585
R674 B.n727 B.n49 585
R675 B.n675 B.n48 585
R676 B.n728 B.n48 585
R677 B.n674 B.n47 585
R678 B.n729 B.n47 585
R679 B.n673 B.n672 585
R680 B.n672 B.n43 585
R681 B.n671 B.n42 585
R682 B.n735 B.n42 585
R683 B.n670 B.n41 585
R684 B.n736 B.n41 585
R685 B.n669 B.n40 585
R686 B.n737 B.n40 585
R687 B.n668 B.n667 585
R688 B.n667 B.n36 585
R689 B.n666 B.n35 585
R690 B.n743 B.n35 585
R691 B.n665 B.n34 585
R692 B.n744 B.n34 585
R693 B.n664 B.n33 585
R694 B.n745 B.n33 585
R695 B.n663 B.n662 585
R696 B.n662 B.n32 585
R697 B.n661 B.n28 585
R698 B.n751 B.n28 585
R699 B.n660 B.n27 585
R700 B.n752 B.n27 585
R701 B.n659 B.n26 585
R702 B.n753 B.n26 585
R703 B.n658 B.n657 585
R704 B.n657 B.n22 585
R705 B.n656 B.n21 585
R706 B.n759 B.n21 585
R707 B.n655 B.n20 585
R708 B.t1 B.n20 585
R709 B.n654 B.n19 585
R710 B.n760 B.n19 585
R711 B.n653 B.n652 585
R712 B.n652 B.n15 585
R713 B.n651 B.n14 585
R714 B.n766 B.n14 585
R715 B.n650 B.n13 585
R716 B.n767 B.n13 585
R717 B.n649 B.n12 585
R718 B.n768 B.n12 585
R719 B.n648 B.n647 585
R720 B.n647 B.n646 585
R721 B.n645 B.n644 585
R722 B.n645 B.n8 585
R723 B.n643 B.n7 585
R724 B.n775 B.n7 585
R725 B.n642 B.n6 585
R726 B.n776 B.n6 585
R727 B.n641 B.n5 585
R728 B.n777 B.n5 585
R729 B.n640 B.n639 585
R730 B.n639 B.n4 585
R731 B.n638 B.n259 585
R732 B.n638 B.n637 585
R733 B.n628 B.n260 585
R734 B.n261 B.n260 585
R735 B.n630 B.n629 585
R736 B.n631 B.n630 585
R737 B.n627 B.n266 585
R738 B.n266 B.n265 585
R739 B.n626 B.n625 585
R740 B.n625 B.n624 585
R741 B.n268 B.n267 585
R742 B.n269 B.n268 585
R743 B.n617 B.n616 585
R744 B.n618 B.n617 585
R745 B.n615 B.n273 585
R746 B.n273 B.t0 585
R747 B.n614 B.n613 585
R748 B.n613 B.n612 585
R749 B.n275 B.n274 585
R750 B.n276 B.n275 585
R751 B.n605 B.n604 585
R752 B.n606 B.n605 585
R753 B.n603 B.n281 585
R754 B.n281 B.n280 585
R755 B.n602 B.n601 585
R756 B.n601 B.n600 585
R757 B.n283 B.n282 585
R758 B.n593 B.n283 585
R759 B.n592 B.n591 585
R760 B.n594 B.n592 585
R761 B.n590 B.n288 585
R762 B.n288 B.n287 585
R763 B.n589 B.n588 585
R764 B.n588 B.n587 585
R765 B.n290 B.n289 585
R766 B.n291 B.n290 585
R767 B.n580 B.n579 585
R768 B.n581 B.n580 585
R769 B.n578 B.n296 585
R770 B.n296 B.n295 585
R771 B.n577 B.n576 585
R772 B.n576 B.n575 585
R773 B.n298 B.n297 585
R774 B.n299 B.n298 585
R775 B.n568 B.n567 585
R776 B.n569 B.n568 585
R777 B.n566 B.n303 585
R778 B.n307 B.n303 585
R779 B.n565 B.n564 585
R780 B.n564 B.n563 585
R781 B.n305 B.n304 585
R782 B.n306 B.n305 585
R783 B.n556 B.n555 585
R784 B.n557 B.n556 585
R785 B.n554 B.n312 585
R786 B.n312 B.n311 585
R787 B.n553 B.n552 585
R788 B.n552 B.n551 585
R789 B.n314 B.n313 585
R790 B.n315 B.n314 585
R791 B.n544 B.n543 585
R792 B.n545 B.n544 585
R793 B.n542 B.n320 585
R794 B.n320 B.n319 585
R795 B.n541 B.n540 585
R796 B.n540 B.n539 585
R797 B.n322 B.n321 585
R798 B.n323 B.n322 585
R799 B.n532 B.n531 585
R800 B.n533 B.n532 585
R801 B.n530 B.n328 585
R802 B.n328 B.n327 585
R803 B.n529 B.n528 585
R804 B.n528 B.n527 585
R805 B.n330 B.n329 585
R806 B.n331 B.n330 585
R807 B.n523 B.n522 585
R808 B.n334 B.n333 585
R809 B.n519 B.n518 585
R810 B.n520 B.n519 585
R811 B.n517 B.n371 585
R812 B.n516 B.n515 585
R813 B.n514 B.n513 585
R814 B.n512 B.n511 585
R815 B.n510 B.n509 585
R816 B.n508 B.n507 585
R817 B.n506 B.n505 585
R818 B.n504 B.n503 585
R819 B.n502 B.n501 585
R820 B.n500 B.n499 585
R821 B.n498 B.n497 585
R822 B.n496 B.n495 585
R823 B.n494 B.n493 585
R824 B.n492 B.n491 585
R825 B.n490 B.n489 585
R826 B.n488 B.n487 585
R827 B.n486 B.n485 585
R828 B.n484 B.n483 585
R829 B.n482 B.n481 585
R830 B.n480 B.n479 585
R831 B.n478 B.n477 585
R832 B.n476 B.n475 585
R833 B.n474 B.n473 585
R834 B.n472 B.n471 585
R835 B.n470 B.n469 585
R836 B.n468 B.n467 585
R837 B.n466 B.n465 585
R838 B.n464 B.n463 585
R839 B.n462 B.n461 585
R840 B.n459 B.n458 585
R841 B.n457 B.n456 585
R842 B.n455 B.n454 585
R843 B.n453 B.n452 585
R844 B.n451 B.n450 585
R845 B.n449 B.n448 585
R846 B.n447 B.n446 585
R847 B.n445 B.n444 585
R848 B.n443 B.n442 585
R849 B.n441 B.n440 585
R850 B.n438 B.n437 585
R851 B.n436 B.n435 585
R852 B.n434 B.n433 585
R853 B.n432 B.n431 585
R854 B.n430 B.n429 585
R855 B.n428 B.n427 585
R856 B.n426 B.n425 585
R857 B.n424 B.n423 585
R858 B.n422 B.n421 585
R859 B.n420 B.n419 585
R860 B.n418 B.n417 585
R861 B.n416 B.n415 585
R862 B.n414 B.n413 585
R863 B.n412 B.n411 585
R864 B.n410 B.n409 585
R865 B.n408 B.n407 585
R866 B.n406 B.n405 585
R867 B.n404 B.n403 585
R868 B.n402 B.n401 585
R869 B.n400 B.n399 585
R870 B.n398 B.n397 585
R871 B.n396 B.n395 585
R872 B.n394 B.n393 585
R873 B.n392 B.n391 585
R874 B.n390 B.n389 585
R875 B.n388 B.n387 585
R876 B.n386 B.n385 585
R877 B.n384 B.n383 585
R878 B.n382 B.n381 585
R879 B.n380 B.n379 585
R880 B.n378 B.n377 585
R881 B.n376 B.n370 585
R882 B.n520 B.n370 585
R883 B.n524 B.n332 585
R884 B.n332 B.n331 585
R885 B.n526 B.n525 585
R886 B.n527 B.n526 585
R887 B.n326 B.n325 585
R888 B.n327 B.n326 585
R889 B.n535 B.n534 585
R890 B.n534 B.n533 585
R891 B.n536 B.n324 585
R892 B.n324 B.n323 585
R893 B.n538 B.n537 585
R894 B.n539 B.n538 585
R895 B.n318 B.n317 585
R896 B.n319 B.n318 585
R897 B.n547 B.n546 585
R898 B.n546 B.n545 585
R899 B.n548 B.n316 585
R900 B.n316 B.n315 585
R901 B.n550 B.n549 585
R902 B.n551 B.n550 585
R903 B.n310 B.n309 585
R904 B.n311 B.n310 585
R905 B.n559 B.n558 585
R906 B.n558 B.n557 585
R907 B.n560 B.n308 585
R908 B.n308 B.n306 585
R909 B.n562 B.n561 585
R910 B.n563 B.n562 585
R911 B.n302 B.n301 585
R912 B.n307 B.n302 585
R913 B.n571 B.n570 585
R914 B.n570 B.n569 585
R915 B.n572 B.n300 585
R916 B.n300 B.n299 585
R917 B.n574 B.n573 585
R918 B.n575 B.n574 585
R919 B.n294 B.n293 585
R920 B.n295 B.n294 585
R921 B.n583 B.n582 585
R922 B.n582 B.n581 585
R923 B.n584 B.n292 585
R924 B.n292 B.n291 585
R925 B.n586 B.n585 585
R926 B.n587 B.n586 585
R927 B.n286 B.n285 585
R928 B.n287 B.n286 585
R929 B.n596 B.n595 585
R930 B.n595 B.n594 585
R931 B.n597 B.n284 585
R932 B.n593 B.n284 585
R933 B.n599 B.n598 585
R934 B.n600 B.n599 585
R935 B.n279 B.n278 585
R936 B.n280 B.n279 585
R937 B.n608 B.n607 585
R938 B.n607 B.n606 585
R939 B.n609 B.n277 585
R940 B.n277 B.n276 585
R941 B.n611 B.n610 585
R942 B.n612 B.n611 585
R943 B.n272 B.n271 585
R944 B.t0 B.n272 585
R945 B.n620 B.n619 585
R946 B.n619 B.n618 585
R947 B.n621 B.n270 585
R948 B.n270 B.n269 585
R949 B.n623 B.n622 585
R950 B.n624 B.n623 585
R951 B.n264 B.n263 585
R952 B.n265 B.n264 585
R953 B.n633 B.n632 585
R954 B.n632 B.n631 585
R955 B.n634 B.n262 585
R956 B.n262 B.n261 585
R957 B.n636 B.n635 585
R958 B.n637 B.n636 585
R959 B.n3 B.n0 585
R960 B.n4 B.n3 585
R961 B.n774 B.n1 585
R962 B.n775 B.n774 585
R963 B.n773 B.n772 585
R964 B.n773 B.n8 585
R965 B.n771 B.n9 585
R966 B.n646 B.n9 585
R967 B.n770 B.n769 585
R968 B.n769 B.n768 585
R969 B.n11 B.n10 585
R970 B.n767 B.n11 585
R971 B.n765 B.n764 585
R972 B.n766 B.n765 585
R973 B.n763 B.n16 585
R974 B.n16 B.n15 585
R975 B.n762 B.n761 585
R976 B.n761 B.n760 585
R977 B.n18 B.n17 585
R978 B.t1 B.n18 585
R979 B.n758 B.n757 585
R980 B.n759 B.n758 585
R981 B.n756 B.n23 585
R982 B.n23 B.n22 585
R983 B.n755 B.n754 585
R984 B.n754 B.n753 585
R985 B.n25 B.n24 585
R986 B.n752 B.n25 585
R987 B.n750 B.n749 585
R988 B.n751 B.n750 585
R989 B.n748 B.n29 585
R990 B.n32 B.n29 585
R991 B.n747 B.n746 585
R992 B.n746 B.n745 585
R993 B.n31 B.n30 585
R994 B.n744 B.n31 585
R995 B.n742 B.n741 585
R996 B.n743 B.n742 585
R997 B.n740 B.n37 585
R998 B.n37 B.n36 585
R999 B.n739 B.n738 585
R1000 B.n738 B.n737 585
R1001 B.n39 B.n38 585
R1002 B.n736 B.n39 585
R1003 B.n734 B.n733 585
R1004 B.n735 B.n734 585
R1005 B.n732 B.n44 585
R1006 B.n44 B.n43 585
R1007 B.n731 B.n730 585
R1008 B.n730 B.n729 585
R1009 B.n46 B.n45 585
R1010 B.n728 B.n46 585
R1011 B.n726 B.n725 585
R1012 B.n727 B.n726 585
R1013 B.n724 B.n51 585
R1014 B.n51 B.n50 585
R1015 B.n723 B.n722 585
R1016 B.n722 B.n721 585
R1017 B.n53 B.n52 585
R1018 B.n720 B.n53 585
R1019 B.n718 B.n717 585
R1020 B.n719 B.n718 585
R1021 B.n716 B.n58 585
R1022 B.n58 B.n57 585
R1023 B.n715 B.n714 585
R1024 B.n714 B.n713 585
R1025 B.n60 B.n59 585
R1026 B.n712 B.n60 585
R1027 B.n710 B.n709 585
R1028 B.n711 B.n710 585
R1029 B.n708 B.n65 585
R1030 B.n65 B.n64 585
R1031 B.n707 B.n706 585
R1032 B.n706 B.n705 585
R1033 B.n67 B.n66 585
R1034 B.n704 B.n67 585
R1035 B.n702 B.n701 585
R1036 B.n703 B.n702 585
R1037 B.n700 B.n72 585
R1038 B.n72 B.n71 585
R1039 B.n778 B.n777 585
R1040 B.n776 B.n2 585
R1041 B.n698 B.n72 526.135
R1042 B.n694 B.n111 526.135
R1043 B.n370 B.n330 526.135
R1044 B.n522 B.n332 526.135
R1045 B.n115 B.t20 350.382
R1046 B.n112 B.t16 350.382
R1047 B.n374 B.t13 350.382
R1048 B.n372 B.t9 350.382
R1049 B.n112 B.t18 261.849
R1050 B.n374 B.t15 261.849
R1051 B.n115 B.t21 261.849
R1052 B.n372 B.t12 261.849
R1053 B.n696 B.n695 256.663
R1054 B.n696 B.n109 256.663
R1055 B.n696 B.n108 256.663
R1056 B.n696 B.n107 256.663
R1057 B.n696 B.n106 256.663
R1058 B.n696 B.n105 256.663
R1059 B.n696 B.n104 256.663
R1060 B.n696 B.n103 256.663
R1061 B.n696 B.n102 256.663
R1062 B.n696 B.n101 256.663
R1063 B.n696 B.n100 256.663
R1064 B.n696 B.n99 256.663
R1065 B.n696 B.n98 256.663
R1066 B.n696 B.n97 256.663
R1067 B.n696 B.n96 256.663
R1068 B.n696 B.n95 256.663
R1069 B.n696 B.n94 256.663
R1070 B.n696 B.n93 256.663
R1071 B.n696 B.n92 256.663
R1072 B.n696 B.n91 256.663
R1073 B.n696 B.n90 256.663
R1074 B.n696 B.n89 256.663
R1075 B.n696 B.n88 256.663
R1076 B.n696 B.n87 256.663
R1077 B.n696 B.n86 256.663
R1078 B.n696 B.n85 256.663
R1079 B.n696 B.n84 256.663
R1080 B.n696 B.n83 256.663
R1081 B.n696 B.n82 256.663
R1082 B.n696 B.n81 256.663
R1083 B.n696 B.n80 256.663
R1084 B.n696 B.n79 256.663
R1085 B.n696 B.n78 256.663
R1086 B.n696 B.n77 256.663
R1087 B.n696 B.n76 256.663
R1088 B.n696 B.n75 256.663
R1089 B.n697 B.n696 256.663
R1090 B.n521 B.n520 256.663
R1091 B.n520 B.n335 256.663
R1092 B.n520 B.n336 256.663
R1093 B.n520 B.n337 256.663
R1094 B.n520 B.n338 256.663
R1095 B.n520 B.n339 256.663
R1096 B.n520 B.n340 256.663
R1097 B.n520 B.n341 256.663
R1098 B.n520 B.n342 256.663
R1099 B.n520 B.n343 256.663
R1100 B.n520 B.n344 256.663
R1101 B.n520 B.n345 256.663
R1102 B.n520 B.n346 256.663
R1103 B.n520 B.n347 256.663
R1104 B.n520 B.n348 256.663
R1105 B.n520 B.n349 256.663
R1106 B.n520 B.n350 256.663
R1107 B.n520 B.n351 256.663
R1108 B.n520 B.n352 256.663
R1109 B.n520 B.n353 256.663
R1110 B.n520 B.n354 256.663
R1111 B.n520 B.n355 256.663
R1112 B.n520 B.n356 256.663
R1113 B.n520 B.n357 256.663
R1114 B.n520 B.n358 256.663
R1115 B.n520 B.n359 256.663
R1116 B.n520 B.n360 256.663
R1117 B.n520 B.n361 256.663
R1118 B.n520 B.n362 256.663
R1119 B.n520 B.n363 256.663
R1120 B.n520 B.n364 256.663
R1121 B.n520 B.n365 256.663
R1122 B.n520 B.n366 256.663
R1123 B.n520 B.n367 256.663
R1124 B.n520 B.n368 256.663
R1125 B.n520 B.n369 256.663
R1126 B.n780 B.n779 256.663
R1127 B.n113 B.t19 227.133
R1128 B.n375 B.t14 227.133
R1129 B.n116 B.t22 227.133
R1130 B.n373 B.t11 227.133
R1131 B.n118 B.n74 163.367
R1132 B.n122 B.n121 163.367
R1133 B.n126 B.n125 163.367
R1134 B.n130 B.n129 163.367
R1135 B.n134 B.n133 163.367
R1136 B.n138 B.n137 163.367
R1137 B.n142 B.n141 163.367
R1138 B.n146 B.n145 163.367
R1139 B.n150 B.n149 163.367
R1140 B.n154 B.n153 163.367
R1141 B.n158 B.n157 163.367
R1142 B.n162 B.n161 163.367
R1143 B.n166 B.n165 163.367
R1144 B.n170 B.n169 163.367
R1145 B.n174 B.n173 163.367
R1146 B.n178 B.n177 163.367
R1147 B.n182 B.n181 163.367
R1148 B.n186 B.n185 163.367
R1149 B.n190 B.n189 163.367
R1150 B.n194 B.n193 163.367
R1151 B.n198 B.n197 163.367
R1152 B.n202 B.n201 163.367
R1153 B.n206 B.n205 163.367
R1154 B.n210 B.n209 163.367
R1155 B.n214 B.n213 163.367
R1156 B.n218 B.n217 163.367
R1157 B.n222 B.n221 163.367
R1158 B.n226 B.n225 163.367
R1159 B.n230 B.n229 163.367
R1160 B.n234 B.n233 163.367
R1161 B.n238 B.n237 163.367
R1162 B.n242 B.n241 163.367
R1163 B.n246 B.n245 163.367
R1164 B.n250 B.n249 163.367
R1165 B.n254 B.n253 163.367
R1166 B.n256 B.n110 163.367
R1167 B.n528 B.n330 163.367
R1168 B.n528 B.n328 163.367
R1169 B.n532 B.n328 163.367
R1170 B.n532 B.n322 163.367
R1171 B.n540 B.n322 163.367
R1172 B.n540 B.n320 163.367
R1173 B.n544 B.n320 163.367
R1174 B.n544 B.n314 163.367
R1175 B.n552 B.n314 163.367
R1176 B.n552 B.n312 163.367
R1177 B.n556 B.n312 163.367
R1178 B.n556 B.n305 163.367
R1179 B.n564 B.n305 163.367
R1180 B.n564 B.n303 163.367
R1181 B.n568 B.n303 163.367
R1182 B.n568 B.n298 163.367
R1183 B.n576 B.n298 163.367
R1184 B.n576 B.n296 163.367
R1185 B.n580 B.n296 163.367
R1186 B.n580 B.n290 163.367
R1187 B.n588 B.n290 163.367
R1188 B.n588 B.n288 163.367
R1189 B.n592 B.n288 163.367
R1190 B.n592 B.n283 163.367
R1191 B.n601 B.n283 163.367
R1192 B.n601 B.n281 163.367
R1193 B.n605 B.n281 163.367
R1194 B.n605 B.n275 163.367
R1195 B.n613 B.n275 163.367
R1196 B.n613 B.n273 163.367
R1197 B.n617 B.n273 163.367
R1198 B.n617 B.n268 163.367
R1199 B.n625 B.n268 163.367
R1200 B.n625 B.n266 163.367
R1201 B.n630 B.n266 163.367
R1202 B.n630 B.n260 163.367
R1203 B.n638 B.n260 163.367
R1204 B.n639 B.n638 163.367
R1205 B.n639 B.n5 163.367
R1206 B.n6 B.n5 163.367
R1207 B.n7 B.n6 163.367
R1208 B.n645 B.n7 163.367
R1209 B.n647 B.n645 163.367
R1210 B.n647 B.n12 163.367
R1211 B.n13 B.n12 163.367
R1212 B.n14 B.n13 163.367
R1213 B.n652 B.n14 163.367
R1214 B.n652 B.n19 163.367
R1215 B.n20 B.n19 163.367
R1216 B.n21 B.n20 163.367
R1217 B.n657 B.n21 163.367
R1218 B.n657 B.n26 163.367
R1219 B.n27 B.n26 163.367
R1220 B.n28 B.n27 163.367
R1221 B.n662 B.n28 163.367
R1222 B.n662 B.n33 163.367
R1223 B.n34 B.n33 163.367
R1224 B.n35 B.n34 163.367
R1225 B.n667 B.n35 163.367
R1226 B.n667 B.n40 163.367
R1227 B.n41 B.n40 163.367
R1228 B.n42 B.n41 163.367
R1229 B.n672 B.n42 163.367
R1230 B.n672 B.n47 163.367
R1231 B.n48 B.n47 163.367
R1232 B.n49 B.n48 163.367
R1233 B.n677 B.n49 163.367
R1234 B.n677 B.n54 163.367
R1235 B.n55 B.n54 163.367
R1236 B.n56 B.n55 163.367
R1237 B.n682 B.n56 163.367
R1238 B.n682 B.n61 163.367
R1239 B.n62 B.n61 163.367
R1240 B.n63 B.n62 163.367
R1241 B.n687 B.n63 163.367
R1242 B.n687 B.n68 163.367
R1243 B.n69 B.n68 163.367
R1244 B.n70 B.n69 163.367
R1245 B.n111 B.n70 163.367
R1246 B.n519 B.n334 163.367
R1247 B.n519 B.n371 163.367
R1248 B.n515 B.n514 163.367
R1249 B.n511 B.n510 163.367
R1250 B.n507 B.n506 163.367
R1251 B.n503 B.n502 163.367
R1252 B.n499 B.n498 163.367
R1253 B.n495 B.n494 163.367
R1254 B.n491 B.n490 163.367
R1255 B.n487 B.n486 163.367
R1256 B.n483 B.n482 163.367
R1257 B.n479 B.n478 163.367
R1258 B.n475 B.n474 163.367
R1259 B.n471 B.n470 163.367
R1260 B.n467 B.n466 163.367
R1261 B.n463 B.n462 163.367
R1262 B.n458 B.n457 163.367
R1263 B.n454 B.n453 163.367
R1264 B.n450 B.n449 163.367
R1265 B.n446 B.n445 163.367
R1266 B.n442 B.n441 163.367
R1267 B.n437 B.n436 163.367
R1268 B.n433 B.n432 163.367
R1269 B.n429 B.n428 163.367
R1270 B.n425 B.n424 163.367
R1271 B.n421 B.n420 163.367
R1272 B.n417 B.n416 163.367
R1273 B.n413 B.n412 163.367
R1274 B.n409 B.n408 163.367
R1275 B.n405 B.n404 163.367
R1276 B.n401 B.n400 163.367
R1277 B.n397 B.n396 163.367
R1278 B.n393 B.n392 163.367
R1279 B.n389 B.n388 163.367
R1280 B.n385 B.n384 163.367
R1281 B.n381 B.n380 163.367
R1282 B.n377 B.n370 163.367
R1283 B.n526 B.n332 163.367
R1284 B.n526 B.n326 163.367
R1285 B.n534 B.n326 163.367
R1286 B.n534 B.n324 163.367
R1287 B.n538 B.n324 163.367
R1288 B.n538 B.n318 163.367
R1289 B.n546 B.n318 163.367
R1290 B.n546 B.n316 163.367
R1291 B.n550 B.n316 163.367
R1292 B.n550 B.n310 163.367
R1293 B.n558 B.n310 163.367
R1294 B.n558 B.n308 163.367
R1295 B.n562 B.n308 163.367
R1296 B.n562 B.n302 163.367
R1297 B.n570 B.n302 163.367
R1298 B.n570 B.n300 163.367
R1299 B.n574 B.n300 163.367
R1300 B.n574 B.n294 163.367
R1301 B.n582 B.n294 163.367
R1302 B.n582 B.n292 163.367
R1303 B.n586 B.n292 163.367
R1304 B.n586 B.n286 163.367
R1305 B.n595 B.n286 163.367
R1306 B.n595 B.n284 163.367
R1307 B.n599 B.n284 163.367
R1308 B.n599 B.n279 163.367
R1309 B.n607 B.n279 163.367
R1310 B.n607 B.n277 163.367
R1311 B.n611 B.n277 163.367
R1312 B.n611 B.n272 163.367
R1313 B.n619 B.n272 163.367
R1314 B.n619 B.n270 163.367
R1315 B.n623 B.n270 163.367
R1316 B.n623 B.n264 163.367
R1317 B.n632 B.n264 163.367
R1318 B.n632 B.n262 163.367
R1319 B.n636 B.n262 163.367
R1320 B.n636 B.n3 163.367
R1321 B.n778 B.n3 163.367
R1322 B.n774 B.n2 163.367
R1323 B.n774 B.n773 163.367
R1324 B.n773 B.n9 163.367
R1325 B.n769 B.n9 163.367
R1326 B.n769 B.n11 163.367
R1327 B.n765 B.n11 163.367
R1328 B.n765 B.n16 163.367
R1329 B.n761 B.n16 163.367
R1330 B.n761 B.n18 163.367
R1331 B.n758 B.n18 163.367
R1332 B.n758 B.n23 163.367
R1333 B.n754 B.n23 163.367
R1334 B.n754 B.n25 163.367
R1335 B.n750 B.n25 163.367
R1336 B.n750 B.n29 163.367
R1337 B.n746 B.n29 163.367
R1338 B.n746 B.n31 163.367
R1339 B.n742 B.n31 163.367
R1340 B.n742 B.n37 163.367
R1341 B.n738 B.n37 163.367
R1342 B.n738 B.n39 163.367
R1343 B.n734 B.n39 163.367
R1344 B.n734 B.n44 163.367
R1345 B.n730 B.n44 163.367
R1346 B.n730 B.n46 163.367
R1347 B.n726 B.n46 163.367
R1348 B.n726 B.n51 163.367
R1349 B.n722 B.n51 163.367
R1350 B.n722 B.n53 163.367
R1351 B.n718 B.n53 163.367
R1352 B.n718 B.n58 163.367
R1353 B.n714 B.n58 163.367
R1354 B.n714 B.n60 163.367
R1355 B.n710 B.n60 163.367
R1356 B.n710 B.n65 163.367
R1357 B.n706 B.n65 163.367
R1358 B.n706 B.n67 163.367
R1359 B.n702 B.n67 163.367
R1360 B.n702 B.n72 163.367
R1361 B.n520 B.n331 107.145
R1362 B.n696 B.n71 107.145
R1363 B.n698 B.n697 71.676
R1364 B.n118 B.n75 71.676
R1365 B.n122 B.n76 71.676
R1366 B.n126 B.n77 71.676
R1367 B.n130 B.n78 71.676
R1368 B.n134 B.n79 71.676
R1369 B.n138 B.n80 71.676
R1370 B.n142 B.n81 71.676
R1371 B.n146 B.n82 71.676
R1372 B.n150 B.n83 71.676
R1373 B.n154 B.n84 71.676
R1374 B.n158 B.n85 71.676
R1375 B.n162 B.n86 71.676
R1376 B.n166 B.n87 71.676
R1377 B.n170 B.n88 71.676
R1378 B.n174 B.n89 71.676
R1379 B.n178 B.n90 71.676
R1380 B.n182 B.n91 71.676
R1381 B.n186 B.n92 71.676
R1382 B.n190 B.n93 71.676
R1383 B.n194 B.n94 71.676
R1384 B.n198 B.n95 71.676
R1385 B.n202 B.n96 71.676
R1386 B.n206 B.n97 71.676
R1387 B.n210 B.n98 71.676
R1388 B.n214 B.n99 71.676
R1389 B.n218 B.n100 71.676
R1390 B.n222 B.n101 71.676
R1391 B.n226 B.n102 71.676
R1392 B.n230 B.n103 71.676
R1393 B.n234 B.n104 71.676
R1394 B.n238 B.n105 71.676
R1395 B.n242 B.n106 71.676
R1396 B.n246 B.n107 71.676
R1397 B.n250 B.n108 71.676
R1398 B.n254 B.n109 71.676
R1399 B.n695 B.n110 71.676
R1400 B.n695 B.n694 71.676
R1401 B.n256 B.n109 71.676
R1402 B.n253 B.n108 71.676
R1403 B.n249 B.n107 71.676
R1404 B.n245 B.n106 71.676
R1405 B.n241 B.n105 71.676
R1406 B.n237 B.n104 71.676
R1407 B.n233 B.n103 71.676
R1408 B.n229 B.n102 71.676
R1409 B.n225 B.n101 71.676
R1410 B.n221 B.n100 71.676
R1411 B.n217 B.n99 71.676
R1412 B.n213 B.n98 71.676
R1413 B.n209 B.n97 71.676
R1414 B.n205 B.n96 71.676
R1415 B.n201 B.n95 71.676
R1416 B.n197 B.n94 71.676
R1417 B.n193 B.n93 71.676
R1418 B.n189 B.n92 71.676
R1419 B.n185 B.n91 71.676
R1420 B.n181 B.n90 71.676
R1421 B.n177 B.n89 71.676
R1422 B.n173 B.n88 71.676
R1423 B.n169 B.n87 71.676
R1424 B.n165 B.n86 71.676
R1425 B.n161 B.n85 71.676
R1426 B.n157 B.n84 71.676
R1427 B.n153 B.n83 71.676
R1428 B.n149 B.n82 71.676
R1429 B.n145 B.n81 71.676
R1430 B.n141 B.n80 71.676
R1431 B.n137 B.n79 71.676
R1432 B.n133 B.n78 71.676
R1433 B.n129 B.n77 71.676
R1434 B.n125 B.n76 71.676
R1435 B.n121 B.n75 71.676
R1436 B.n697 B.n74 71.676
R1437 B.n522 B.n521 71.676
R1438 B.n371 B.n335 71.676
R1439 B.n514 B.n336 71.676
R1440 B.n510 B.n337 71.676
R1441 B.n506 B.n338 71.676
R1442 B.n502 B.n339 71.676
R1443 B.n498 B.n340 71.676
R1444 B.n494 B.n341 71.676
R1445 B.n490 B.n342 71.676
R1446 B.n486 B.n343 71.676
R1447 B.n482 B.n344 71.676
R1448 B.n478 B.n345 71.676
R1449 B.n474 B.n346 71.676
R1450 B.n470 B.n347 71.676
R1451 B.n466 B.n348 71.676
R1452 B.n462 B.n349 71.676
R1453 B.n457 B.n350 71.676
R1454 B.n453 B.n351 71.676
R1455 B.n449 B.n352 71.676
R1456 B.n445 B.n353 71.676
R1457 B.n441 B.n354 71.676
R1458 B.n436 B.n355 71.676
R1459 B.n432 B.n356 71.676
R1460 B.n428 B.n357 71.676
R1461 B.n424 B.n358 71.676
R1462 B.n420 B.n359 71.676
R1463 B.n416 B.n360 71.676
R1464 B.n412 B.n361 71.676
R1465 B.n408 B.n362 71.676
R1466 B.n404 B.n363 71.676
R1467 B.n400 B.n364 71.676
R1468 B.n396 B.n365 71.676
R1469 B.n392 B.n366 71.676
R1470 B.n388 B.n367 71.676
R1471 B.n384 B.n368 71.676
R1472 B.n380 B.n369 71.676
R1473 B.n521 B.n334 71.676
R1474 B.n515 B.n335 71.676
R1475 B.n511 B.n336 71.676
R1476 B.n507 B.n337 71.676
R1477 B.n503 B.n338 71.676
R1478 B.n499 B.n339 71.676
R1479 B.n495 B.n340 71.676
R1480 B.n491 B.n341 71.676
R1481 B.n487 B.n342 71.676
R1482 B.n483 B.n343 71.676
R1483 B.n479 B.n344 71.676
R1484 B.n475 B.n345 71.676
R1485 B.n471 B.n346 71.676
R1486 B.n467 B.n347 71.676
R1487 B.n463 B.n348 71.676
R1488 B.n458 B.n349 71.676
R1489 B.n454 B.n350 71.676
R1490 B.n450 B.n351 71.676
R1491 B.n446 B.n352 71.676
R1492 B.n442 B.n353 71.676
R1493 B.n437 B.n354 71.676
R1494 B.n433 B.n355 71.676
R1495 B.n429 B.n356 71.676
R1496 B.n425 B.n357 71.676
R1497 B.n421 B.n358 71.676
R1498 B.n417 B.n359 71.676
R1499 B.n413 B.n360 71.676
R1500 B.n409 B.n361 71.676
R1501 B.n405 B.n362 71.676
R1502 B.n401 B.n363 71.676
R1503 B.n397 B.n364 71.676
R1504 B.n393 B.n365 71.676
R1505 B.n389 B.n366 71.676
R1506 B.n385 B.n367 71.676
R1507 B.n381 B.n368 71.676
R1508 B.n377 B.n369 71.676
R1509 B.n779 B.n778 71.676
R1510 B.n779 B.n2 71.676
R1511 B.n117 B.n116 59.5399
R1512 B.n114 B.n113 59.5399
R1513 B.n439 B.n375 59.5399
R1514 B.n460 B.n373 59.5399
R1515 B.n527 B.n331 53.1822
R1516 B.n527 B.n327 53.1822
R1517 B.n533 B.n327 53.1822
R1518 B.n533 B.n323 53.1822
R1519 B.n539 B.n323 53.1822
R1520 B.n545 B.n319 53.1822
R1521 B.n545 B.n315 53.1822
R1522 B.n551 B.n315 53.1822
R1523 B.n551 B.n311 53.1822
R1524 B.n557 B.n311 53.1822
R1525 B.n557 B.n306 53.1822
R1526 B.n563 B.n306 53.1822
R1527 B.n563 B.n307 53.1822
R1528 B.n569 B.n299 53.1822
R1529 B.n575 B.n299 53.1822
R1530 B.n575 B.n295 53.1822
R1531 B.n581 B.n295 53.1822
R1532 B.n587 B.n291 53.1822
R1533 B.n587 B.n287 53.1822
R1534 B.n594 B.n287 53.1822
R1535 B.n594 B.n593 53.1822
R1536 B.n600 B.n280 53.1822
R1537 B.n606 B.n280 53.1822
R1538 B.n606 B.n276 53.1822
R1539 B.n612 B.n276 53.1822
R1540 B.n612 B.t0 53.1822
R1541 B.n618 B.t0 53.1822
R1542 B.n618 B.n269 53.1822
R1543 B.n624 B.n269 53.1822
R1544 B.n624 B.n265 53.1822
R1545 B.n631 B.n265 53.1822
R1546 B.n637 B.n261 53.1822
R1547 B.n637 B.n4 53.1822
R1548 B.n777 B.n4 53.1822
R1549 B.n777 B.n776 53.1822
R1550 B.n776 B.n775 53.1822
R1551 B.n775 B.n8 53.1822
R1552 B.n646 B.n8 53.1822
R1553 B.n768 B.n767 53.1822
R1554 B.n767 B.n766 53.1822
R1555 B.n766 B.n15 53.1822
R1556 B.n760 B.n15 53.1822
R1557 B.n760 B.t1 53.1822
R1558 B.t1 B.n759 53.1822
R1559 B.n759 B.n22 53.1822
R1560 B.n753 B.n22 53.1822
R1561 B.n753 B.n752 53.1822
R1562 B.n752 B.n751 53.1822
R1563 B.n745 B.n32 53.1822
R1564 B.n745 B.n744 53.1822
R1565 B.n744 B.n743 53.1822
R1566 B.n743 B.n36 53.1822
R1567 B.n737 B.n736 53.1822
R1568 B.n736 B.n735 53.1822
R1569 B.n735 B.n43 53.1822
R1570 B.n729 B.n43 53.1822
R1571 B.n728 B.n727 53.1822
R1572 B.n727 B.n50 53.1822
R1573 B.n721 B.n50 53.1822
R1574 B.n721 B.n720 53.1822
R1575 B.n720 B.n719 53.1822
R1576 B.n719 B.n57 53.1822
R1577 B.n713 B.n57 53.1822
R1578 B.n713 B.n712 53.1822
R1579 B.n711 B.n64 53.1822
R1580 B.n705 B.n64 53.1822
R1581 B.n705 B.n704 53.1822
R1582 B.n704 B.n703 53.1822
R1583 B.n703 B.n71 53.1822
R1584 B.n569 B.t8 42.233
R1585 B.n729 B.t4 42.233
R1586 B.n539 B.t10 39.1047
R1587 B.n593 B.t2 39.1047
R1588 B.t5 B.n261 39.1047
R1589 B.n646 B.t7 39.1047
R1590 B.n32 B.t3 39.1047
R1591 B.t17 B.n711 39.1047
R1592 B.n116 B.n115 34.7157
R1593 B.n113 B.n112 34.7157
R1594 B.n375 B.n374 34.7157
R1595 B.n373 B.n372 34.7157
R1596 B.n524 B.n523 34.1859
R1597 B.n376 B.n329 34.1859
R1598 B.n693 B.n692 34.1859
R1599 B.n700 B.n699 34.1859
R1600 B.t23 B.n291 28.1555
R1601 B.t6 B.n36 28.1555
R1602 B.n581 B.t23 25.0272
R1603 B.n737 B.t6 25.0272
R1604 B B.n780 18.0485
R1605 B.t10 B.n319 14.078
R1606 B.n600 B.t2 14.078
R1607 B.n631 B.t5 14.078
R1608 B.n768 B.t7 14.078
R1609 B.n751 B.t3 14.078
R1610 B.n712 B.t17 14.078
R1611 B.n307 B.t8 10.9497
R1612 B.t4 B.n728 10.9497
R1613 B.n525 B.n524 10.6151
R1614 B.n525 B.n325 10.6151
R1615 B.n535 B.n325 10.6151
R1616 B.n536 B.n535 10.6151
R1617 B.n537 B.n536 10.6151
R1618 B.n537 B.n317 10.6151
R1619 B.n547 B.n317 10.6151
R1620 B.n548 B.n547 10.6151
R1621 B.n549 B.n548 10.6151
R1622 B.n549 B.n309 10.6151
R1623 B.n559 B.n309 10.6151
R1624 B.n560 B.n559 10.6151
R1625 B.n561 B.n560 10.6151
R1626 B.n561 B.n301 10.6151
R1627 B.n571 B.n301 10.6151
R1628 B.n572 B.n571 10.6151
R1629 B.n573 B.n572 10.6151
R1630 B.n573 B.n293 10.6151
R1631 B.n583 B.n293 10.6151
R1632 B.n584 B.n583 10.6151
R1633 B.n585 B.n584 10.6151
R1634 B.n585 B.n285 10.6151
R1635 B.n596 B.n285 10.6151
R1636 B.n597 B.n596 10.6151
R1637 B.n598 B.n597 10.6151
R1638 B.n598 B.n278 10.6151
R1639 B.n608 B.n278 10.6151
R1640 B.n609 B.n608 10.6151
R1641 B.n610 B.n609 10.6151
R1642 B.n610 B.n271 10.6151
R1643 B.n620 B.n271 10.6151
R1644 B.n621 B.n620 10.6151
R1645 B.n622 B.n621 10.6151
R1646 B.n622 B.n263 10.6151
R1647 B.n633 B.n263 10.6151
R1648 B.n634 B.n633 10.6151
R1649 B.n635 B.n634 10.6151
R1650 B.n635 B.n0 10.6151
R1651 B.n523 B.n333 10.6151
R1652 B.n518 B.n333 10.6151
R1653 B.n518 B.n517 10.6151
R1654 B.n517 B.n516 10.6151
R1655 B.n516 B.n513 10.6151
R1656 B.n513 B.n512 10.6151
R1657 B.n512 B.n509 10.6151
R1658 B.n509 B.n508 10.6151
R1659 B.n508 B.n505 10.6151
R1660 B.n505 B.n504 10.6151
R1661 B.n504 B.n501 10.6151
R1662 B.n501 B.n500 10.6151
R1663 B.n500 B.n497 10.6151
R1664 B.n497 B.n496 10.6151
R1665 B.n496 B.n493 10.6151
R1666 B.n493 B.n492 10.6151
R1667 B.n492 B.n489 10.6151
R1668 B.n489 B.n488 10.6151
R1669 B.n488 B.n485 10.6151
R1670 B.n485 B.n484 10.6151
R1671 B.n484 B.n481 10.6151
R1672 B.n481 B.n480 10.6151
R1673 B.n480 B.n477 10.6151
R1674 B.n477 B.n476 10.6151
R1675 B.n476 B.n473 10.6151
R1676 B.n473 B.n472 10.6151
R1677 B.n472 B.n469 10.6151
R1678 B.n469 B.n468 10.6151
R1679 B.n468 B.n465 10.6151
R1680 B.n465 B.n464 10.6151
R1681 B.n464 B.n461 10.6151
R1682 B.n459 B.n456 10.6151
R1683 B.n456 B.n455 10.6151
R1684 B.n455 B.n452 10.6151
R1685 B.n452 B.n451 10.6151
R1686 B.n451 B.n448 10.6151
R1687 B.n448 B.n447 10.6151
R1688 B.n447 B.n444 10.6151
R1689 B.n444 B.n443 10.6151
R1690 B.n443 B.n440 10.6151
R1691 B.n438 B.n435 10.6151
R1692 B.n435 B.n434 10.6151
R1693 B.n434 B.n431 10.6151
R1694 B.n431 B.n430 10.6151
R1695 B.n430 B.n427 10.6151
R1696 B.n427 B.n426 10.6151
R1697 B.n426 B.n423 10.6151
R1698 B.n423 B.n422 10.6151
R1699 B.n422 B.n419 10.6151
R1700 B.n419 B.n418 10.6151
R1701 B.n418 B.n415 10.6151
R1702 B.n415 B.n414 10.6151
R1703 B.n414 B.n411 10.6151
R1704 B.n411 B.n410 10.6151
R1705 B.n410 B.n407 10.6151
R1706 B.n407 B.n406 10.6151
R1707 B.n406 B.n403 10.6151
R1708 B.n403 B.n402 10.6151
R1709 B.n402 B.n399 10.6151
R1710 B.n399 B.n398 10.6151
R1711 B.n398 B.n395 10.6151
R1712 B.n395 B.n394 10.6151
R1713 B.n394 B.n391 10.6151
R1714 B.n391 B.n390 10.6151
R1715 B.n390 B.n387 10.6151
R1716 B.n387 B.n386 10.6151
R1717 B.n386 B.n383 10.6151
R1718 B.n383 B.n382 10.6151
R1719 B.n382 B.n379 10.6151
R1720 B.n379 B.n378 10.6151
R1721 B.n378 B.n376 10.6151
R1722 B.n529 B.n329 10.6151
R1723 B.n530 B.n529 10.6151
R1724 B.n531 B.n530 10.6151
R1725 B.n531 B.n321 10.6151
R1726 B.n541 B.n321 10.6151
R1727 B.n542 B.n541 10.6151
R1728 B.n543 B.n542 10.6151
R1729 B.n543 B.n313 10.6151
R1730 B.n553 B.n313 10.6151
R1731 B.n554 B.n553 10.6151
R1732 B.n555 B.n554 10.6151
R1733 B.n555 B.n304 10.6151
R1734 B.n565 B.n304 10.6151
R1735 B.n566 B.n565 10.6151
R1736 B.n567 B.n566 10.6151
R1737 B.n567 B.n297 10.6151
R1738 B.n577 B.n297 10.6151
R1739 B.n578 B.n577 10.6151
R1740 B.n579 B.n578 10.6151
R1741 B.n579 B.n289 10.6151
R1742 B.n589 B.n289 10.6151
R1743 B.n590 B.n589 10.6151
R1744 B.n591 B.n590 10.6151
R1745 B.n591 B.n282 10.6151
R1746 B.n602 B.n282 10.6151
R1747 B.n603 B.n602 10.6151
R1748 B.n604 B.n603 10.6151
R1749 B.n604 B.n274 10.6151
R1750 B.n614 B.n274 10.6151
R1751 B.n615 B.n614 10.6151
R1752 B.n616 B.n615 10.6151
R1753 B.n616 B.n267 10.6151
R1754 B.n626 B.n267 10.6151
R1755 B.n627 B.n626 10.6151
R1756 B.n629 B.n627 10.6151
R1757 B.n629 B.n628 10.6151
R1758 B.n628 B.n259 10.6151
R1759 B.n640 B.n259 10.6151
R1760 B.n641 B.n640 10.6151
R1761 B.n642 B.n641 10.6151
R1762 B.n643 B.n642 10.6151
R1763 B.n644 B.n643 10.6151
R1764 B.n648 B.n644 10.6151
R1765 B.n649 B.n648 10.6151
R1766 B.n650 B.n649 10.6151
R1767 B.n651 B.n650 10.6151
R1768 B.n653 B.n651 10.6151
R1769 B.n654 B.n653 10.6151
R1770 B.n655 B.n654 10.6151
R1771 B.n656 B.n655 10.6151
R1772 B.n658 B.n656 10.6151
R1773 B.n659 B.n658 10.6151
R1774 B.n660 B.n659 10.6151
R1775 B.n661 B.n660 10.6151
R1776 B.n663 B.n661 10.6151
R1777 B.n664 B.n663 10.6151
R1778 B.n665 B.n664 10.6151
R1779 B.n666 B.n665 10.6151
R1780 B.n668 B.n666 10.6151
R1781 B.n669 B.n668 10.6151
R1782 B.n670 B.n669 10.6151
R1783 B.n671 B.n670 10.6151
R1784 B.n673 B.n671 10.6151
R1785 B.n674 B.n673 10.6151
R1786 B.n675 B.n674 10.6151
R1787 B.n676 B.n675 10.6151
R1788 B.n678 B.n676 10.6151
R1789 B.n679 B.n678 10.6151
R1790 B.n680 B.n679 10.6151
R1791 B.n681 B.n680 10.6151
R1792 B.n683 B.n681 10.6151
R1793 B.n684 B.n683 10.6151
R1794 B.n685 B.n684 10.6151
R1795 B.n686 B.n685 10.6151
R1796 B.n688 B.n686 10.6151
R1797 B.n689 B.n688 10.6151
R1798 B.n690 B.n689 10.6151
R1799 B.n691 B.n690 10.6151
R1800 B.n692 B.n691 10.6151
R1801 B.n772 B.n1 10.6151
R1802 B.n772 B.n771 10.6151
R1803 B.n771 B.n770 10.6151
R1804 B.n770 B.n10 10.6151
R1805 B.n764 B.n10 10.6151
R1806 B.n764 B.n763 10.6151
R1807 B.n763 B.n762 10.6151
R1808 B.n762 B.n17 10.6151
R1809 B.n757 B.n17 10.6151
R1810 B.n757 B.n756 10.6151
R1811 B.n756 B.n755 10.6151
R1812 B.n755 B.n24 10.6151
R1813 B.n749 B.n24 10.6151
R1814 B.n749 B.n748 10.6151
R1815 B.n748 B.n747 10.6151
R1816 B.n747 B.n30 10.6151
R1817 B.n741 B.n30 10.6151
R1818 B.n741 B.n740 10.6151
R1819 B.n740 B.n739 10.6151
R1820 B.n739 B.n38 10.6151
R1821 B.n733 B.n38 10.6151
R1822 B.n733 B.n732 10.6151
R1823 B.n732 B.n731 10.6151
R1824 B.n731 B.n45 10.6151
R1825 B.n725 B.n45 10.6151
R1826 B.n725 B.n724 10.6151
R1827 B.n724 B.n723 10.6151
R1828 B.n723 B.n52 10.6151
R1829 B.n717 B.n52 10.6151
R1830 B.n717 B.n716 10.6151
R1831 B.n716 B.n715 10.6151
R1832 B.n715 B.n59 10.6151
R1833 B.n709 B.n59 10.6151
R1834 B.n709 B.n708 10.6151
R1835 B.n708 B.n707 10.6151
R1836 B.n707 B.n66 10.6151
R1837 B.n701 B.n66 10.6151
R1838 B.n701 B.n700 10.6151
R1839 B.n699 B.n73 10.6151
R1840 B.n119 B.n73 10.6151
R1841 B.n120 B.n119 10.6151
R1842 B.n123 B.n120 10.6151
R1843 B.n124 B.n123 10.6151
R1844 B.n127 B.n124 10.6151
R1845 B.n128 B.n127 10.6151
R1846 B.n131 B.n128 10.6151
R1847 B.n132 B.n131 10.6151
R1848 B.n135 B.n132 10.6151
R1849 B.n136 B.n135 10.6151
R1850 B.n139 B.n136 10.6151
R1851 B.n140 B.n139 10.6151
R1852 B.n143 B.n140 10.6151
R1853 B.n144 B.n143 10.6151
R1854 B.n147 B.n144 10.6151
R1855 B.n148 B.n147 10.6151
R1856 B.n151 B.n148 10.6151
R1857 B.n152 B.n151 10.6151
R1858 B.n155 B.n152 10.6151
R1859 B.n156 B.n155 10.6151
R1860 B.n159 B.n156 10.6151
R1861 B.n160 B.n159 10.6151
R1862 B.n163 B.n160 10.6151
R1863 B.n164 B.n163 10.6151
R1864 B.n167 B.n164 10.6151
R1865 B.n168 B.n167 10.6151
R1866 B.n171 B.n168 10.6151
R1867 B.n172 B.n171 10.6151
R1868 B.n175 B.n172 10.6151
R1869 B.n176 B.n175 10.6151
R1870 B.n180 B.n179 10.6151
R1871 B.n183 B.n180 10.6151
R1872 B.n184 B.n183 10.6151
R1873 B.n187 B.n184 10.6151
R1874 B.n188 B.n187 10.6151
R1875 B.n191 B.n188 10.6151
R1876 B.n192 B.n191 10.6151
R1877 B.n195 B.n192 10.6151
R1878 B.n196 B.n195 10.6151
R1879 B.n200 B.n199 10.6151
R1880 B.n203 B.n200 10.6151
R1881 B.n204 B.n203 10.6151
R1882 B.n207 B.n204 10.6151
R1883 B.n208 B.n207 10.6151
R1884 B.n211 B.n208 10.6151
R1885 B.n212 B.n211 10.6151
R1886 B.n215 B.n212 10.6151
R1887 B.n216 B.n215 10.6151
R1888 B.n219 B.n216 10.6151
R1889 B.n220 B.n219 10.6151
R1890 B.n223 B.n220 10.6151
R1891 B.n224 B.n223 10.6151
R1892 B.n227 B.n224 10.6151
R1893 B.n228 B.n227 10.6151
R1894 B.n231 B.n228 10.6151
R1895 B.n232 B.n231 10.6151
R1896 B.n235 B.n232 10.6151
R1897 B.n236 B.n235 10.6151
R1898 B.n239 B.n236 10.6151
R1899 B.n240 B.n239 10.6151
R1900 B.n243 B.n240 10.6151
R1901 B.n244 B.n243 10.6151
R1902 B.n247 B.n244 10.6151
R1903 B.n248 B.n247 10.6151
R1904 B.n251 B.n248 10.6151
R1905 B.n252 B.n251 10.6151
R1906 B.n255 B.n252 10.6151
R1907 B.n257 B.n255 10.6151
R1908 B.n258 B.n257 10.6151
R1909 B.n693 B.n258 10.6151
R1910 B.n461 B.n460 9.36635
R1911 B.n439 B.n438 9.36635
R1912 B.n176 B.n117 9.36635
R1913 B.n199 B.n114 9.36635
R1914 B.n780 B.n0 8.11757
R1915 B.n780 B.n1 8.11757
R1916 B.n460 B.n459 1.24928
R1917 B.n440 B.n439 1.24928
R1918 B.n179 B.n117 1.24928
R1919 B.n196 B.n114 1.24928
R1920 VP.n36 VP.n35 181.852
R1921 VP.n62 VP.n61 181.852
R1922 VP.n34 VP.n33 181.852
R1923 VP.n15 VP.t0 175.512
R1924 VP.n16 VP.n13 161.3
R1925 VP.n18 VP.n17 161.3
R1926 VP.n19 VP.n12 161.3
R1927 VP.n21 VP.n20 161.3
R1928 VP.n22 VP.n11 161.3
R1929 VP.n24 VP.n23 161.3
R1930 VP.n25 VP.n10 161.3
R1931 VP.n28 VP.n27 161.3
R1932 VP.n29 VP.n9 161.3
R1933 VP.n31 VP.n30 161.3
R1934 VP.n32 VP.n8 161.3
R1935 VP.n60 VP.n0 161.3
R1936 VP.n59 VP.n58 161.3
R1937 VP.n57 VP.n1 161.3
R1938 VP.n56 VP.n55 161.3
R1939 VP.n53 VP.n2 161.3
R1940 VP.n52 VP.n51 161.3
R1941 VP.n50 VP.n3 161.3
R1942 VP.n49 VP.n48 161.3
R1943 VP.n47 VP.n4 161.3
R1944 VP.n46 VP.n45 161.3
R1945 VP.n44 VP.n5 161.3
R1946 VP.n43 VP.n42 161.3
R1947 VP.n40 VP.n6 161.3
R1948 VP.n39 VP.n38 161.3
R1949 VP.n37 VP.n7 161.3
R1950 VP.n48 VP.t7 145.095
R1951 VP.n35 VP.t5 145.095
R1952 VP.n41 VP.t8 145.095
R1953 VP.n54 VP.t4 145.095
R1954 VP.n61 VP.t1 145.095
R1955 VP.n20 VP.t9 145.095
R1956 VP.n33 VP.t6 145.095
R1957 VP.n26 VP.t2 145.095
R1958 VP.n14 VP.t3 145.095
R1959 VP.n40 VP.n39 56.5193
R1960 VP.n59 VP.n1 56.5193
R1961 VP.n31 VP.n9 56.5193
R1962 VP.n15 VP.n14 51.5804
R1963 VP.n47 VP.n46 50.6917
R1964 VP.n52 VP.n3 50.6917
R1965 VP.n24 VP.n11 50.6917
R1966 VP.n19 VP.n18 50.6917
R1967 VP.n36 VP.n34 44.3073
R1968 VP.n46 VP.n5 30.2951
R1969 VP.n53 VP.n52 30.2951
R1970 VP.n25 VP.n24 30.2951
R1971 VP.n18 VP.n13 30.2951
R1972 VP.n39 VP.n7 24.4675
R1973 VP.n42 VP.n40 24.4675
R1974 VP.n48 VP.n47 24.4675
R1975 VP.n48 VP.n3 24.4675
R1976 VP.n55 VP.n1 24.4675
R1977 VP.n60 VP.n59 24.4675
R1978 VP.n32 VP.n31 24.4675
R1979 VP.n27 VP.n9 24.4675
R1980 VP.n20 VP.n19 24.4675
R1981 VP.n20 VP.n11 24.4675
R1982 VP.n16 VP.n15 18.3855
R1983 VP.n41 VP.n5 14.1914
R1984 VP.n54 VP.n53 14.1914
R1985 VP.n26 VP.n25 14.1914
R1986 VP.n14 VP.n13 14.1914
R1987 VP.n42 VP.n41 10.2766
R1988 VP.n55 VP.n54 10.2766
R1989 VP.n27 VP.n26 10.2766
R1990 VP.n35 VP.n7 3.91522
R1991 VP.n61 VP.n60 3.91522
R1992 VP.n33 VP.n32 3.91522
R1993 VP.n17 VP.n16 0.189894
R1994 VP.n17 VP.n12 0.189894
R1995 VP.n21 VP.n12 0.189894
R1996 VP.n22 VP.n21 0.189894
R1997 VP.n23 VP.n22 0.189894
R1998 VP.n23 VP.n10 0.189894
R1999 VP.n28 VP.n10 0.189894
R2000 VP.n29 VP.n28 0.189894
R2001 VP.n30 VP.n29 0.189894
R2002 VP.n30 VP.n8 0.189894
R2003 VP.n34 VP.n8 0.189894
R2004 VP.n37 VP.n36 0.189894
R2005 VP.n38 VP.n37 0.189894
R2006 VP.n38 VP.n6 0.189894
R2007 VP.n43 VP.n6 0.189894
R2008 VP.n44 VP.n43 0.189894
R2009 VP.n45 VP.n44 0.189894
R2010 VP.n45 VP.n4 0.189894
R2011 VP.n49 VP.n4 0.189894
R2012 VP.n50 VP.n49 0.189894
R2013 VP.n51 VP.n50 0.189894
R2014 VP.n51 VP.n2 0.189894
R2015 VP.n56 VP.n2 0.189894
R2016 VP.n57 VP.n56 0.189894
R2017 VP.n58 VP.n57 0.189894
R2018 VP.n58 VP.n0 0.189894
R2019 VP.n62 VP.n0 0.189894
R2020 VP VP.n62 0.0516364
R2021 VDD1.n42 VDD1.n0 289.615
R2022 VDD1.n91 VDD1.n49 289.615
R2023 VDD1.n43 VDD1.n42 185
R2024 VDD1.n41 VDD1.n40 185
R2025 VDD1.n4 VDD1.n3 185
R2026 VDD1.n35 VDD1.n34 185
R2027 VDD1.n33 VDD1.n32 185
R2028 VDD1.n8 VDD1.n7 185
R2029 VDD1.n27 VDD1.n26 185
R2030 VDD1.n25 VDD1.n24 185
R2031 VDD1.n12 VDD1.n11 185
R2032 VDD1.n19 VDD1.n18 185
R2033 VDD1.n17 VDD1.n16 185
R2034 VDD1.n66 VDD1.n65 185
R2035 VDD1.n68 VDD1.n67 185
R2036 VDD1.n61 VDD1.n60 185
R2037 VDD1.n74 VDD1.n73 185
R2038 VDD1.n76 VDD1.n75 185
R2039 VDD1.n57 VDD1.n56 185
R2040 VDD1.n82 VDD1.n81 185
R2041 VDD1.n84 VDD1.n83 185
R2042 VDD1.n53 VDD1.n52 185
R2043 VDD1.n90 VDD1.n89 185
R2044 VDD1.n92 VDD1.n91 185
R2045 VDD1.n15 VDD1.t9 147.659
R2046 VDD1.n64 VDD1.t4 147.659
R2047 VDD1.n42 VDD1.n41 104.615
R2048 VDD1.n41 VDD1.n3 104.615
R2049 VDD1.n34 VDD1.n3 104.615
R2050 VDD1.n34 VDD1.n33 104.615
R2051 VDD1.n33 VDD1.n7 104.615
R2052 VDD1.n26 VDD1.n7 104.615
R2053 VDD1.n26 VDD1.n25 104.615
R2054 VDD1.n25 VDD1.n11 104.615
R2055 VDD1.n18 VDD1.n11 104.615
R2056 VDD1.n18 VDD1.n17 104.615
R2057 VDD1.n67 VDD1.n66 104.615
R2058 VDD1.n67 VDD1.n60 104.615
R2059 VDD1.n74 VDD1.n60 104.615
R2060 VDD1.n75 VDD1.n74 104.615
R2061 VDD1.n75 VDD1.n56 104.615
R2062 VDD1.n82 VDD1.n56 104.615
R2063 VDD1.n83 VDD1.n82 104.615
R2064 VDD1.n83 VDD1.n52 104.615
R2065 VDD1.n90 VDD1.n52 104.615
R2066 VDD1.n91 VDD1.n90 104.615
R2067 VDD1.n99 VDD1.n98 63.2945
R2068 VDD1.n101 VDD1.n100 62.1927
R2069 VDD1.n48 VDD1.n47 62.1927
R2070 VDD1.n97 VDD1.n96 62.1925
R2071 VDD1.n17 VDD1.t9 52.3082
R2072 VDD1.n66 VDD1.t4 52.3082
R2073 VDD1.n48 VDD1.n46 48.6618
R2074 VDD1.n97 VDD1.n95 48.6618
R2075 VDD1.n101 VDD1.n99 39.9772
R2076 VDD1.n16 VDD1.n15 15.6677
R2077 VDD1.n65 VDD1.n64 15.6677
R2078 VDD1.n19 VDD1.n14 12.8005
R2079 VDD1.n68 VDD1.n63 12.8005
R2080 VDD1.n20 VDD1.n12 12.0247
R2081 VDD1.n69 VDD1.n61 12.0247
R2082 VDD1.n24 VDD1.n23 11.249
R2083 VDD1.n73 VDD1.n72 11.249
R2084 VDD1.n27 VDD1.n10 10.4732
R2085 VDD1.n76 VDD1.n59 10.4732
R2086 VDD1.n28 VDD1.n8 9.69747
R2087 VDD1.n77 VDD1.n57 9.69747
R2088 VDD1.n46 VDD1.n45 9.45567
R2089 VDD1.n95 VDD1.n94 9.45567
R2090 VDD1.n2 VDD1.n1 9.3005
R2091 VDD1.n45 VDD1.n44 9.3005
R2092 VDD1.n39 VDD1.n38 9.3005
R2093 VDD1.n37 VDD1.n36 9.3005
R2094 VDD1.n6 VDD1.n5 9.3005
R2095 VDD1.n31 VDD1.n30 9.3005
R2096 VDD1.n29 VDD1.n28 9.3005
R2097 VDD1.n10 VDD1.n9 9.3005
R2098 VDD1.n23 VDD1.n22 9.3005
R2099 VDD1.n21 VDD1.n20 9.3005
R2100 VDD1.n14 VDD1.n13 9.3005
R2101 VDD1.n88 VDD1.n87 9.3005
R2102 VDD1.n51 VDD1.n50 9.3005
R2103 VDD1.n94 VDD1.n93 9.3005
R2104 VDD1.n55 VDD1.n54 9.3005
R2105 VDD1.n80 VDD1.n79 9.3005
R2106 VDD1.n78 VDD1.n77 9.3005
R2107 VDD1.n59 VDD1.n58 9.3005
R2108 VDD1.n72 VDD1.n71 9.3005
R2109 VDD1.n70 VDD1.n69 9.3005
R2110 VDD1.n63 VDD1.n62 9.3005
R2111 VDD1.n86 VDD1.n85 9.3005
R2112 VDD1.n46 VDD1.n0 8.92171
R2113 VDD1.n32 VDD1.n31 8.92171
R2114 VDD1.n81 VDD1.n80 8.92171
R2115 VDD1.n95 VDD1.n49 8.92171
R2116 VDD1.n44 VDD1.n43 8.14595
R2117 VDD1.n35 VDD1.n6 8.14595
R2118 VDD1.n84 VDD1.n55 8.14595
R2119 VDD1.n93 VDD1.n92 8.14595
R2120 VDD1.n40 VDD1.n2 7.3702
R2121 VDD1.n36 VDD1.n4 7.3702
R2122 VDD1.n85 VDD1.n53 7.3702
R2123 VDD1.n89 VDD1.n51 7.3702
R2124 VDD1.n40 VDD1.n39 6.59444
R2125 VDD1.n39 VDD1.n4 6.59444
R2126 VDD1.n88 VDD1.n53 6.59444
R2127 VDD1.n89 VDD1.n88 6.59444
R2128 VDD1.n43 VDD1.n2 5.81868
R2129 VDD1.n36 VDD1.n35 5.81868
R2130 VDD1.n85 VDD1.n84 5.81868
R2131 VDD1.n92 VDD1.n51 5.81868
R2132 VDD1.n44 VDD1.n0 5.04292
R2133 VDD1.n32 VDD1.n6 5.04292
R2134 VDD1.n81 VDD1.n55 5.04292
R2135 VDD1.n93 VDD1.n49 5.04292
R2136 VDD1.n15 VDD1.n13 4.38563
R2137 VDD1.n64 VDD1.n62 4.38563
R2138 VDD1.n31 VDD1.n8 4.26717
R2139 VDD1.n80 VDD1.n57 4.26717
R2140 VDD1.n28 VDD1.n27 3.49141
R2141 VDD1.n77 VDD1.n76 3.49141
R2142 VDD1.n24 VDD1.n10 2.71565
R2143 VDD1.n73 VDD1.n59 2.71565
R2144 VDD1.n100 VDD1.t7 2.25306
R2145 VDD1.n100 VDD1.t3 2.25306
R2146 VDD1.n47 VDD1.t6 2.25306
R2147 VDD1.n47 VDD1.t0 2.25306
R2148 VDD1.n98 VDD1.t5 2.25306
R2149 VDD1.n98 VDD1.t8 2.25306
R2150 VDD1.n96 VDD1.t1 2.25306
R2151 VDD1.n96 VDD1.t2 2.25306
R2152 VDD1.n23 VDD1.n12 1.93989
R2153 VDD1.n72 VDD1.n61 1.93989
R2154 VDD1.n20 VDD1.n19 1.16414
R2155 VDD1.n69 VDD1.n68 1.16414
R2156 VDD1 VDD1.n101 1.09964
R2157 VDD1 VDD1.n48 0.444466
R2158 VDD1.n16 VDD1.n14 0.388379
R2159 VDD1.n65 VDD1.n63 0.388379
R2160 VDD1.n99 VDD1.n97 0.33093
R2161 VDD1.n45 VDD1.n1 0.155672
R2162 VDD1.n38 VDD1.n1 0.155672
R2163 VDD1.n38 VDD1.n37 0.155672
R2164 VDD1.n37 VDD1.n5 0.155672
R2165 VDD1.n30 VDD1.n5 0.155672
R2166 VDD1.n30 VDD1.n29 0.155672
R2167 VDD1.n29 VDD1.n9 0.155672
R2168 VDD1.n22 VDD1.n9 0.155672
R2169 VDD1.n22 VDD1.n21 0.155672
R2170 VDD1.n21 VDD1.n13 0.155672
R2171 VDD1.n70 VDD1.n62 0.155672
R2172 VDD1.n71 VDD1.n70 0.155672
R2173 VDD1.n71 VDD1.n58 0.155672
R2174 VDD1.n78 VDD1.n58 0.155672
R2175 VDD1.n79 VDD1.n78 0.155672
R2176 VDD1.n79 VDD1.n54 0.155672
R2177 VDD1.n86 VDD1.n54 0.155672
R2178 VDD1.n87 VDD1.n86 0.155672
R2179 VDD1.n87 VDD1.n50 0.155672
R2180 VDD1.n94 VDD1.n50 0.155672
C0 VTAIL VN 7.14159f
C1 VP VTAIL 7.15593f
C2 VDD1 VTAIL 8.97096f
C3 VP VN 6.12781f
C4 VDD1 VN 0.150779f
C5 VDD1 VP 7.12919f
C6 VDD2 VTAIL 9.01369f
C7 VDD2 VN 6.84532f
C8 VP VDD2 0.437932f
C9 VDD1 VDD2 1.43288f
C10 VDD2 B 5.310319f
C11 VDD1 B 5.274548f
C12 VTAIL B 6.041904f
C13 VN B 12.50644f
C14 VP B 10.949032f
C15 VDD1.n0 B 0.033241f
C16 VDD1.n1 B 0.022881f
C17 VDD1.n2 B 0.012295f
C18 VDD1.n3 B 0.029061f
C19 VDD1.n4 B 0.013018f
C20 VDD1.n5 B 0.022881f
C21 VDD1.n6 B 0.012295f
C22 VDD1.n7 B 0.029061f
C23 VDD1.n8 B 0.013018f
C24 VDD1.n9 B 0.022881f
C25 VDD1.n10 B 0.012295f
C26 VDD1.n11 B 0.029061f
C27 VDD1.n12 B 0.013018f
C28 VDD1.n13 B 0.837423f
C29 VDD1.n14 B 0.012295f
C30 VDD1.t9 B 0.047441f
C31 VDD1.n15 B 0.11363f
C32 VDD1.n16 B 0.017167f
C33 VDD1.n17 B 0.021796f
C34 VDD1.n18 B 0.029061f
C35 VDD1.n19 B 0.013018f
C36 VDD1.n20 B 0.012295f
C37 VDD1.n21 B 0.022881f
C38 VDD1.n22 B 0.022881f
C39 VDD1.n23 B 0.012295f
C40 VDD1.n24 B 0.013018f
C41 VDD1.n25 B 0.029061f
C42 VDD1.n26 B 0.029061f
C43 VDD1.n27 B 0.013018f
C44 VDD1.n28 B 0.012295f
C45 VDD1.n29 B 0.022881f
C46 VDD1.n30 B 0.022881f
C47 VDD1.n31 B 0.012295f
C48 VDD1.n32 B 0.013018f
C49 VDD1.n33 B 0.029061f
C50 VDD1.n34 B 0.029061f
C51 VDD1.n35 B 0.013018f
C52 VDD1.n36 B 0.012295f
C53 VDD1.n37 B 0.022881f
C54 VDD1.n38 B 0.022881f
C55 VDD1.n39 B 0.012295f
C56 VDD1.n40 B 0.013018f
C57 VDD1.n41 B 0.029061f
C58 VDD1.n42 B 0.064823f
C59 VDD1.n43 B 0.013018f
C60 VDD1.n44 B 0.012295f
C61 VDD1.n45 B 0.050074f
C62 VDD1.n46 B 0.057155f
C63 VDD1.t6 B 0.158932f
C64 VDD1.t0 B 0.158932f
C65 VDD1.n47 B 1.37727f
C66 VDD1.n48 B 0.490975f
C67 VDD1.n49 B 0.033241f
C68 VDD1.n50 B 0.022881f
C69 VDD1.n51 B 0.012295f
C70 VDD1.n52 B 0.029061f
C71 VDD1.n53 B 0.013018f
C72 VDD1.n54 B 0.022881f
C73 VDD1.n55 B 0.012295f
C74 VDD1.n56 B 0.029061f
C75 VDD1.n57 B 0.013018f
C76 VDD1.n58 B 0.022881f
C77 VDD1.n59 B 0.012295f
C78 VDD1.n60 B 0.029061f
C79 VDD1.n61 B 0.013018f
C80 VDD1.n62 B 0.837423f
C81 VDD1.n63 B 0.012295f
C82 VDD1.t4 B 0.047441f
C83 VDD1.n64 B 0.11363f
C84 VDD1.n65 B 0.017167f
C85 VDD1.n66 B 0.021796f
C86 VDD1.n67 B 0.029061f
C87 VDD1.n68 B 0.013018f
C88 VDD1.n69 B 0.012295f
C89 VDD1.n70 B 0.022881f
C90 VDD1.n71 B 0.022881f
C91 VDD1.n72 B 0.012295f
C92 VDD1.n73 B 0.013018f
C93 VDD1.n74 B 0.029061f
C94 VDD1.n75 B 0.029061f
C95 VDD1.n76 B 0.013018f
C96 VDD1.n77 B 0.012295f
C97 VDD1.n78 B 0.022881f
C98 VDD1.n79 B 0.022881f
C99 VDD1.n80 B 0.012295f
C100 VDD1.n81 B 0.013018f
C101 VDD1.n82 B 0.029061f
C102 VDD1.n83 B 0.029061f
C103 VDD1.n84 B 0.013018f
C104 VDD1.n85 B 0.012295f
C105 VDD1.n86 B 0.022881f
C106 VDD1.n87 B 0.022881f
C107 VDD1.n88 B 0.012295f
C108 VDD1.n89 B 0.013018f
C109 VDD1.n90 B 0.029061f
C110 VDD1.n91 B 0.064823f
C111 VDD1.n92 B 0.013018f
C112 VDD1.n93 B 0.012295f
C113 VDD1.n94 B 0.050074f
C114 VDD1.n95 B 0.057155f
C115 VDD1.t1 B 0.158932f
C116 VDD1.t2 B 0.158932f
C117 VDD1.n96 B 1.37727f
C118 VDD1.n97 B 0.484216f
C119 VDD1.t5 B 0.158932f
C120 VDD1.t8 B 0.158932f
C121 VDD1.n98 B 1.3842f
C122 VDD1.n99 B 2.02347f
C123 VDD1.t7 B 0.158932f
C124 VDD1.t3 B 0.158932f
C125 VDD1.n100 B 1.37727f
C126 VDD1.n101 B 2.24878f
C127 VP.n0 B 0.031542f
C128 VP.t1 B 1.0914f
C129 VP.n1 B 0.040336f
C130 VP.n2 B 0.031542f
C131 VP.t4 B 1.0914f
C132 VP.n3 B 0.057585f
C133 VP.n4 B 0.031542f
C134 VP.t7 B 1.0914f
C135 VP.n5 B 0.05084f
C136 VP.n6 B 0.031542f
C137 VP.n7 B 0.034407f
C138 VP.n8 B 0.031542f
C139 VP.t6 B 1.0914f
C140 VP.n9 B 0.040336f
C141 VP.n10 B 0.031542f
C142 VP.t2 B 1.0914f
C143 VP.n11 B 0.057585f
C144 VP.n12 B 0.031542f
C145 VP.t9 B 1.0914f
C146 VP.n13 B 0.05084f
C147 VP.t0 B 1.18234f
C148 VP.t3 B 1.0914f
C149 VP.n14 B 0.466844f
C150 VP.n15 B 0.482379f
C151 VP.n16 B 0.195308f
C152 VP.n17 B 0.031542f
C153 VP.n18 B 0.030269f
C154 VP.n19 B 0.057585f
C155 VP.n20 B 0.436925f
C156 VP.n21 B 0.031542f
C157 VP.n22 B 0.031542f
C158 VP.n23 B 0.031542f
C159 VP.n24 B 0.030269f
C160 VP.n25 B 0.05084f
C161 VP.n26 B 0.407162f
C162 VP.n27 B 0.041953f
C163 VP.n28 B 0.031542f
C164 VP.n29 B 0.031542f
C165 VP.n30 B 0.031542f
C166 VP.n31 B 0.051762f
C167 VP.n32 B 0.034407f
C168 VP.n33 B 0.461364f
C169 VP.n34 B 1.42803f
C170 VP.t5 B 1.0914f
C171 VP.n35 B 0.461364f
C172 VP.n36 B 1.45362f
C173 VP.n37 B 0.031542f
C174 VP.n38 B 0.031542f
C175 VP.n39 B 0.051762f
C176 VP.n40 B 0.040336f
C177 VP.t8 B 1.0914f
C178 VP.n41 B 0.407162f
C179 VP.n42 B 0.041953f
C180 VP.n43 B 0.031542f
C181 VP.n44 B 0.031542f
C182 VP.n45 B 0.031542f
C183 VP.n46 B 0.030269f
C184 VP.n47 B 0.057585f
C185 VP.n48 B 0.436925f
C186 VP.n49 B 0.031542f
C187 VP.n50 B 0.031542f
C188 VP.n51 B 0.031542f
C189 VP.n52 B 0.030269f
C190 VP.n53 B 0.05084f
C191 VP.n54 B 0.407162f
C192 VP.n55 B 0.041953f
C193 VP.n56 B 0.031542f
C194 VP.n57 B 0.031542f
C195 VP.n58 B 0.031542f
C196 VP.n59 B 0.051762f
C197 VP.n60 B 0.034407f
C198 VP.n61 B 0.461364f
C199 VP.n62 B 0.03135f
C200 VTAIL.t9 B 0.176432f
C201 VTAIL.t11 B 0.176432f
C202 VTAIL.n0 B 1.45209f
C203 VTAIL.n1 B 0.457884f
C204 VTAIL.n2 B 0.036902f
C205 VTAIL.n3 B 0.0254f
C206 VTAIL.n4 B 0.013649f
C207 VTAIL.n5 B 0.032261f
C208 VTAIL.n6 B 0.014452f
C209 VTAIL.n7 B 0.0254f
C210 VTAIL.n8 B 0.013649f
C211 VTAIL.n9 B 0.032261f
C212 VTAIL.n10 B 0.014452f
C213 VTAIL.n11 B 0.0254f
C214 VTAIL.n12 B 0.013649f
C215 VTAIL.n13 B 0.032261f
C216 VTAIL.n14 B 0.014452f
C217 VTAIL.n15 B 0.92963f
C218 VTAIL.n16 B 0.013649f
C219 VTAIL.t5 B 0.052665f
C220 VTAIL.n17 B 0.126141f
C221 VTAIL.n18 B 0.019058f
C222 VTAIL.n19 B 0.024196f
C223 VTAIL.n20 B 0.032261f
C224 VTAIL.n21 B 0.014452f
C225 VTAIL.n22 B 0.013649f
C226 VTAIL.n23 B 0.0254f
C227 VTAIL.n24 B 0.0254f
C228 VTAIL.n25 B 0.013649f
C229 VTAIL.n26 B 0.014452f
C230 VTAIL.n27 B 0.032261f
C231 VTAIL.n28 B 0.032261f
C232 VTAIL.n29 B 0.014452f
C233 VTAIL.n30 B 0.013649f
C234 VTAIL.n31 B 0.0254f
C235 VTAIL.n32 B 0.0254f
C236 VTAIL.n33 B 0.013649f
C237 VTAIL.n34 B 0.014452f
C238 VTAIL.n35 B 0.032261f
C239 VTAIL.n36 B 0.032261f
C240 VTAIL.n37 B 0.014452f
C241 VTAIL.n38 B 0.013649f
C242 VTAIL.n39 B 0.0254f
C243 VTAIL.n40 B 0.0254f
C244 VTAIL.n41 B 0.013649f
C245 VTAIL.n42 B 0.014452f
C246 VTAIL.n43 B 0.032261f
C247 VTAIL.n44 B 0.071961f
C248 VTAIL.n45 B 0.014452f
C249 VTAIL.n46 B 0.013649f
C250 VTAIL.n47 B 0.055588f
C251 VTAIL.n48 B 0.040385f
C252 VTAIL.n49 B 0.247829f
C253 VTAIL.t2 B 0.176432f
C254 VTAIL.t0 B 0.176432f
C255 VTAIL.n50 B 1.45209f
C256 VTAIL.n51 B 0.50939f
C257 VTAIL.t8 B 0.176432f
C258 VTAIL.t19 B 0.176432f
C259 VTAIL.n52 B 1.45209f
C260 VTAIL.n53 B 1.6009f
C261 VTAIL.t17 B 0.176432f
C262 VTAIL.t10 B 0.176432f
C263 VTAIL.n54 B 1.45209f
C264 VTAIL.n55 B 1.60089f
C265 VTAIL.t14 B 0.176432f
C266 VTAIL.t18 B 0.176432f
C267 VTAIL.n56 B 1.45209f
C268 VTAIL.n57 B 0.50938f
C269 VTAIL.n58 B 0.036902f
C270 VTAIL.n59 B 0.0254f
C271 VTAIL.n60 B 0.013649f
C272 VTAIL.n61 B 0.032261f
C273 VTAIL.n62 B 0.014452f
C274 VTAIL.n63 B 0.0254f
C275 VTAIL.n64 B 0.013649f
C276 VTAIL.n65 B 0.032261f
C277 VTAIL.n66 B 0.014452f
C278 VTAIL.n67 B 0.0254f
C279 VTAIL.n68 B 0.013649f
C280 VTAIL.n69 B 0.032261f
C281 VTAIL.n70 B 0.014452f
C282 VTAIL.n71 B 0.92963f
C283 VTAIL.n72 B 0.013649f
C284 VTAIL.t12 B 0.052665f
C285 VTAIL.n73 B 0.126141f
C286 VTAIL.n74 B 0.019058f
C287 VTAIL.n75 B 0.024196f
C288 VTAIL.n76 B 0.032261f
C289 VTAIL.n77 B 0.014452f
C290 VTAIL.n78 B 0.013649f
C291 VTAIL.n79 B 0.0254f
C292 VTAIL.n80 B 0.0254f
C293 VTAIL.n81 B 0.013649f
C294 VTAIL.n82 B 0.014452f
C295 VTAIL.n83 B 0.032261f
C296 VTAIL.n84 B 0.032261f
C297 VTAIL.n85 B 0.014452f
C298 VTAIL.n86 B 0.013649f
C299 VTAIL.n87 B 0.0254f
C300 VTAIL.n88 B 0.0254f
C301 VTAIL.n89 B 0.013649f
C302 VTAIL.n90 B 0.014452f
C303 VTAIL.n91 B 0.032261f
C304 VTAIL.n92 B 0.032261f
C305 VTAIL.n93 B 0.014452f
C306 VTAIL.n94 B 0.013649f
C307 VTAIL.n95 B 0.0254f
C308 VTAIL.n96 B 0.0254f
C309 VTAIL.n97 B 0.013649f
C310 VTAIL.n98 B 0.014452f
C311 VTAIL.n99 B 0.032261f
C312 VTAIL.n100 B 0.071961f
C313 VTAIL.n101 B 0.014452f
C314 VTAIL.n102 B 0.013649f
C315 VTAIL.n103 B 0.055588f
C316 VTAIL.n104 B 0.040385f
C317 VTAIL.n105 B 0.247829f
C318 VTAIL.t7 B 0.176432f
C319 VTAIL.t1 B 0.176432f
C320 VTAIL.n106 B 1.45209f
C321 VTAIL.n107 B 0.484686f
C322 VTAIL.t3 B 0.176432f
C323 VTAIL.t6 B 0.176432f
C324 VTAIL.n108 B 1.45209f
C325 VTAIL.n109 B 0.50938f
C326 VTAIL.n110 B 0.036902f
C327 VTAIL.n111 B 0.0254f
C328 VTAIL.n112 B 0.013649f
C329 VTAIL.n113 B 0.032261f
C330 VTAIL.n114 B 0.014452f
C331 VTAIL.n115 B 0.0254f
C332 VTAIL.n116 B 0.013649f
C333 VTAIL.n117 B 0.032261f
C334 VTAIL.n118 B 0.014452f
C335 VTAIL.n119 B 0.0254f
C336 VTAIL.n120 B 0.013649f
C337 VTAIL.n121 B 0.032261f
C338 VTAIL.n122 B 0.014452f
C339 VTAIL.n123 B 0.92963f
C340 VTAIL.n124 B 0.013649f
C341 VTAIL.t4 B 0.052665f
C342 VTAIL.n125 B 0.126141f
C343 VTAIL.n126 B 0.019058f
C344 VTAIL.n127 B 0.024196f
C345 VTAIL.n128 B 0.032261f
C346 VTAIL.n129 B 0.014452f
C347 VTAIL.n130 B 0.013649f
C348 VTAIL.n131 B 0.0254f
C349 VTAIL.n132 B 0.0254f
C350 VTAIL.n133 B 0.013649f
C351 VTAIL.n134 B 0.014452f
C352 VTAIL.n135 B 0.032261f
C353 VTAIL.n136 B 0.032261f
C354 VTAIL.n137 B 0.014452f
C355 VTAIL.n138 B 0.013649f
C356 VTAIL.n139 B 0.0254f
C357 VTAIL.n140 B 0.0254f
C358 VTAIL.n141 B 0.013649f
C359 VTAIL.n142 B 0.014452f
C360 VTAIL.n143 B 0.032261f
C361 VTAIL.n144 B 0.032261f
C362 VTAIL.n145 B 0.014452f
C363 VTAIL.n146 B 0.013649f
C364 VTAIL.n147 B 0.0254f
C365 VTAIL.n148 B 0.0254f
C366 VTAIL.n149 B 0.013649f
C367 VTAIL.n150 B 0.014452f
C368 VTAIL.n151 B 0.032261f
C369 VTAIL.n152 B 0.071961f
C370 VTAIL.n153 B 0.014452f
C371 VTAIL.n154 B 0.013649f
C372 VTAIL.n155 B 0.055588f
C373 VTAIL.n156 B 0.040385f
C374 VTAIL.n157 B 1.23774f
C375 VTAIL.n158 B 0.036902f
C376 VTAIL.n159 B 0.0254f
C377 VTAIL.n160 B 0.013649f
C378 VTAIL.n161 B 0.032261f
C379 VTAIL.n162 B 0.014452f
C380 VTAIL.n163 B 0.0254f
C381 VTAIL.n164 B 0.013649f
C382 VTAIL.n165 B 0.032261f
C383 VTAIL.n166 B 0.014452f
C384 VTAIL.n167 B 0.0254f
C385 VTAIL.n168 B 0.013649f
C386 VTAIL.n169 B 0.032261f
C387 VTAIL.n170 B 0.014452f
C388 VTAIL.n171 B 0.92963f
C389 VTAIL.n172 B 0.013649f
C390 VTAIL.t15 B 0.052665f
C391 VTAIL.n173 B 0.126141f
C392 VTAIL.n174 B 0.019058f
C393 VTAIL.n175 B 0.024196f
C394 VTAIL.n176 B 0.032261f
C395 VTAIL.n177 B 0.014452f
C396 VTAIL.n178 B 0.013649f
C397 VTAIL.n179 B 0.0254f
C398 VTAIL.n180 B 0.0254f
C399 VTAIL.n181 B 0.013649f
C400 VTAIL.n182 B 0.014452f
C401 VTAIL.n183 B 0.032261f
C402 VTAIL.n184 B 0.032261f
C403 VTAIL.n185 B 0.014452f
C404 VTAIL.n186 B 0.013649f
C405 VTAIL.n187 B 0.0254f
C406 VTAIL.n188 B 0.0254f
C407 VTAIL.n189 B 0.013649f
C408 VTAIL.n190 B 0.014452f
C409 VTAIL.n191 B 0.032261f
C410 VTAIL.n192 B 0.032261f
C411 VTAIL.n193 B 0.014452f
C412 VTAIL.n194 B 0.013649f
C413 VTAIL.n195 B 0.0254f
C414 VTAIL.n196 B 0.0254f
C415 VTAIL.n197 B 0.013649f
C416 VTAIL.n198 B 0.014452f
C417 VTAIL.n199 B 0.032261f
C418 VTAIL.n200 B 0.071961f
C419 VTAIL.n201 B 0.014452f
C420 VTAIL.n202 B 0.013649f
C421 VTAIL.n203 B 0.055588f
C422 VTAIL.n204 B 0.040385f
C423 VTAIL.n205 B 1.23774f
C424 VTAIL.t16 B 0.176432f
C425 VTAIL.t13 B 0.176432f
C426 VTAIL.n206 B 1.45209f
C427 VTAIL.n207 B 0.409906f
C428 VDD2.n0 B 0.032794f
C429 VDD2.n1 B 0.022573f
C430 VDD2.n2 B 0.01213f
C431 VDD2.n3 B 0.02867f
C432 VDD2.n4 B 0.012843f
C433 VDD2.n5 B 0.022573f
C434 VDD2.n6 B 0.01213f
C435 VDD2.n7 B 0.02867f
C436 VDD2.n8 B 0.012843f
C437 VDD2.n9 B 0.022573f
C438 VDD2.n10 B 0.01213f
C439 VDD2.n11 B 0.02867f
C440 VDD2.n12 B 0.012843f
C441 VDD2.n13 B 0.826155f
C442 VDD2.n14 B 0.01213f
C443 VDD2.t7 B 0.046803f
C444 VDD2.n15 B 0.112101f
C445 VDD2.n16 B 0.016936f
C446 VDD2.n17 B 0.021503f
C447 VDD2.n18 B 0.02867f
C448 VDD2.n19 B 0.012843f
C449 VDD2.n20 B 0.01213f
C450 VDD2.n21 B 0.022573f
C451 VDD2.n22 B 0.022573f
C452 VDD2.n23 B 0.01213f
C453 VDD2.n24 B 0.012843f
C454 VDD2.n25 B 0.02867f
C455 VDD2.n26 B 0.02867f
C456 VDD2.n27 B 0.012843f
C457 VDD2.n28 B 0.01213f
C458 VDD2.n29 B 0.022573f
C459 VDD2.n30 B 0.022573f
C460 VDD2.n31 B 0.01213f
C461 VDD2.n32 B 0.012843f
C462 VDD2.n33 B 0.02867f
C463 VDD2.n34 B 0.02867f
C464 VDD2.n35 B 0.012843f
C465 VDD2.n36 B 0.01213f
C466 VDD2.n37 B 0.022573f
C467 VDD2.n38 B 0.022573f
C468 VDD2.n39 B 0.01213f
C469 VDD2.n40 B 0.012843f
C470 VDD2.n41 B 0.02867f
C471 VDD2.n42 B 0.063951f
C472 VDD2.n43 B 0.012843f
C473 VDD2.n44 B 0.01213f
C474 VDD2.n45 B 0.049401f
C475 VDD2.n46 B 0.056386f
C476 VDD2.t5 B 0.156794f
C477 VDD2.t2 B 0.156794f
C478 VDD2.n47 B 1.35874f
C479 VDD2.n48 B 0.477701f
C480 VDD2.t0 B 0.156794f
C481 VDD2.t1 B 0.156794f
C482 VDD2.n49 B 1.36557f
C483 VDD2.n50 B 1.91169f
C484 VDD2.n51 B 0.032794f
C485 VDD2.n52 B 0.022573f
C486 VDD2.n53 B 0.01213f
C487 VDD2.n54 B 0.02867f
C488 VDD2.n55 B 0.012843f
C489 VDD2.n56 B 0.022573f
C490 VDD2.n57 B 0.01213f
C491 VDD2.n58 B 0.02867f
C492 VDD2.n59 B 0.012843f
C493 VDD2.n60 B 0.022573f
C494 VDD2.n61 B 0.01213f
C495 VDD2.n62 B 0.02867f
C496 VDD2.n63 B 0.012843f
C497 VDD2.n64 B 0.826155f
C498 VDD2.n65 B 0.01213f
C499 VDD2.t4 B 0.046803f
C500 VDD2.n66 B 0.112101f
C501 VDD2.n67 B 0.016936f
C502 VDD2.n68 B 0.021503f
C503 VDD2.n69 B 0.02867f
C504 VDD2.n70 B 0.012843f
C505 VDD2.n71 B 0.01213f
C506 VDD2.n72 B 0.022573f
C507 VDD2.n73 B 0.022573f
C508 VDD2.n74 B 0.01213f
C509 VDD2.n75 B 0.012843f
C510 VDD2.n76 B 0.02867f
C511 VDD2.n77 B 0.02867f
C512 VDD2.n78 B 0.012843f
C513 VDD2.n79 B 0.01213f
C514 VDD2.n80 B 0.022573f
C515 VDD2.n81 B 0.022573f
C516 VDD2.n82 B 0.01213f
C517 VDD2.n83 B 0.012843f
C518 VDD2.n84 B 0.02867f
C519 VDD2.n85 B 0.02867f
C520 VDD2.n86 B 0.012843f
C521 VDD2.n87 B 0.01213f
C522 VDD2.n88 B 0.022573f
C523 VDD2.n89 B 0.022573f
C524 VDD2.n90 B 0.01213f
C525 VDD2.n91 B 0.012843f
C526 VDD2.n92 B 0.02867f
C527 VDD2.n93 B 0.063951f
C528 VDD2.n94 B 0.012843f
C529 VDD2.n95 B 0.01213f
C530 VDD2.n96 B 0.049401f
C531 VDD2.n97 B 0.051499f
C532 VDD2.n98 B 1.98194f
C533 VDD2.t8 B 0.156794f
C534 VDD2.t6 B 0.156794f
C535 VDD2.n99 B 1.35874f
C536 VDD2.n100 B 0.335141f
C537 VDD2.t3 B 0.156794f
C538 VDD2.t9 B 0.156794f
C539 VDD2.n101 B 1.36555f
C540 VN.n0 B 0.030856f
C541 VN.t3 B 1.06768f
C542 VN.n1 B 0.039459f
C543 VN.n2 B 0.030856f
C544 VN.t5 B 1.06768f
C545 VN.n3 B 0.056334f
C546 VN.n4 B 0.030856f
C547 VN.t2 B 1.06768f
C548 VN.n5 B 0.049735f
C549 VN.t9 B 1.15664f
C550 VN.t7 B 1.06768f
C551 VN.n6 B 0.456697f
C552 VN.n7 B 0.471895f
C553 VN.n8 B 0.191063f
C554 VN.n9 B 0.030856f
C555 VN.n10 B 0.029611f
C556 VN.n11 B 0.056334f
C557 VN.n12 B 0.427429f
C558 VN.n13 B 0.030856f
C559 VN.n14 B 0.030856f
C560 VN.n15 B 0.030856f
C561 VN.n16 B 0.029611f
C562 VN.n17 B 0.049735f
C563 VN.n18 B 0.398313f
C564 VN.n19 B 0.041041f
C565 VN.n20 B 0.030856f
C566 VN.n21 B 0.030856f
C567 VN.n22 B 0.030856f
C568 VN.n23 B 0.050637f
C569 VN.n24 B 0.033659f
C570 VN.n25 B 0.451337f
C571 VN.n26 B 0.030669f
C572 VN.n27 B 0.030856f
C573 VN.t1 B 1.06768f
C574 VN.n28 B 0.039459f
C575 VN.n29 B 0.030856f
C576 VN.t8 B 1.06768f
C577 VN.n30 B 0.056334f
C578 VN.n31 B 0.030856f
C579 VN.t4 B 1.06768f
C580 VN.n32 B 0.049735f
C581 VN.t6 B 1.15664f
C582 VN.t0 B 1.06768f
C583 VN.n33 B 0.456697f
C584 VN.n34 B 0.471895f
C585 VN.n35 B 0.191063f
C586 VN.n36 B 0.030856f
C587 VN.n37 B 0.029611f
C588 VN.n38 B 0.056334f
C589 VN.n39 B 0.427429f
C590 VN.n40 B 0.030856f
C591 VN.n41 B 0.030856f
C592 VN.n42 B 0.030856f
C593 VN.n43 B 0.029611f
C594 VN.n44 B 0.049735f
C595 VN.n45 B 0.398313f
C596 VN.n46 B 0.041041f
C597 VN.n47 B 0.030856f
C598 VN.n48 B 0.030856f
C599 VN.n49 B 0.030856f
C600 VN.n50 B 0.050637f
C601 VN.n51 B 0.033659f
C602 VN.n52 B 0.451337f
C603 VN.n53 B 1.41718f
.ends

