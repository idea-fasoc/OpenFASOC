* NGSPICE file created from diff_pair_sample_0594.ext - technology: sky130A

.subckt diff_pair_sample_0594 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t8 w_n4000_n4480# sky130_fd_pr__pfet_01v8 ad=2.8974 pd=17.89 as=2.8974 ps=17.89 w=17.56 l=2.7
X1 B.t11 B.t9 B.t10 w_n4000_n4480# sky130_fd_pr__pfet_01v8 ad=6.8484 pd=35.9 as=0 ps=0 w=17.56 l=2.7
X2 VDD2.t7 VN.t0 VTAIL.t4 w_n4000_n4480# sky130_fd_pr__pfet_01v8 ad=2.8974 pd=17.89 as=2.8974 ps=17.89 w=17.56 l=2.7
X3 VTAIL.t9 VP.t1 VDD1.t6 w_n4000_n4480# sky130_fd_pr__pfet_01v8 ad=2.8974 pd=17.89 as=2.8974 ps=17.89 w=17.56 l=2.7
X4 VTAIL.t11 VP.t2 VDD1.t5 w_n4000_n4480# sky130_fd_pr__pfet_01v8 ad=2.8974 pd=17.89 as=2.8974 ps=17.89 w=17.56 l=2.7
X5 B.t8 B.t6 B.t7 w_n4000_n4480# sky130_fd_pr__pfet_01v8 ad=6.8484 pd=35.9 as=0 ps=0 w=17.56 l=2.7
X6 VDD1.t4 VP.t3 VTAIL.t12 w_n4000_n4480# sky130_fd_pr__pfet_01v8 ad=2.8974 pd=17.89 as=6.8484 ps=35.9 w=17.56 l=2.7
X7 VTAIL.t5 VN.t1 VDD2.t6 w_n4000_n4480# sky130_fd_pr__pfet_01v8 ad=6.8484 pd=35.9 as=2.8974 ps=17.89 w=17.56 l=2.7
X8 VTAIL.t2 VN.t2 VDD2.t5 w_n4000_n4480# sky130_fd_pr__pfet_01v8 ad=6.8484 pd=35.9 as=2.8974 ps=17.89 w=17.56 l=2.7
X9 VDD1.t3 VP.t4 VTAIL.t14 w_n4000_n4480# sky130_fd_pr__pfet_01v8 ad=2.8974 pd=17.89 as=2.8974 ps=17.89 w=17.56 l=2.7
X10 VTAIL.t3 VN.t3 VDD2.t4 w_n4000_n4480# sky130_fd_pr__pfet_01v8 ad=2.8974 pd=17.89 as=2.8974 ps=17.89 w=17.56 l=2.7
X11 VDD2.t3 VN.t4 VTAIL.t1 w_n4000_n4480# sky130_fd_pr__pfet_01v8 ad=2.8974 pd=17.89 as=6.8484 ps=35.9 w=17.56 l=2.7
X12 VDD1.t2 VP.t5 VTAIL.t13 w_n4000_n4480# sky130_fd_pr__pfet_01v8 ad=2.8974 pd=17.89 as=6.8484 ps=35.9 w=17.56 l=2.7
X13 B.t5 B.t3 B.t4 w_n4000_n4480# sky130_fd_pr__pfet_01v8 ad=6.8484 pd=35.9 as=0 ps=0 w=17.56 l=2.7
X14 VTAIL.t7 VN.t5 VDD2.t2 w_n4000_n4480# sky130_fd_pr__pfet_01v8 ad=2.8974 pd=17.89 as=2.8974 ps=17.89 w=17.56 l=2.7
X15 VTAIL.t15 VP.t6 VDD1.t1 w_n4000_n4480# sky130_fd_pr__pfet_01v8 ad=6.8484 pd=35.9 as=2.8974 ps=17.89 w=17.56 l=2.7
X16 VTAIL.t10 VP.t7 VDD1.t0 w_n4000_n4480# sky130_fd_pr__pfet_01v8 ad=6.8484 pd=35.9 as=2.8974 ps=17.89 w=17.56 l=2.7
X17 B.t2 B.t0 B.t1 w_n4000_n4480# sky130_fd_pr__pfet_01v8 ad=6.8484 pd=35.9 as=0 ps=0 w=17.56 l=2.7
X18 VDD2.t1 VN.t6 VTAIL.t0 w_n4000_n4480# sky130_fd_pr__pfet_01v8 ad=2.8974 pd=17.89 as=6.8484 ps=35.9 w=17.56 l=2.7
X19 VDD2.t0 VN.t7 VTAIL.t6 w_n4000_n4480# sky130_fd_pr__pfet_01v8 ad=2.8974 pd=17.89 as=2.8974 ps=17.89 w=17.56 l=2.7
R0 VP.n19 VP.t7 187.621
R1 VP.n21 VP.n20 161.3
R2 VP.n22 VP.n17 161.3
R3 VP.n24 VP.n23 161.3
R4 VP.n25 VP.n16 161.3
R5 VP.n27 VP.n26 161.3
R6 VP.n28 VP.n15 161.3
R7 VP.n30 VP.n29 161.3
R8 VP.n32 VP.n31 161.3
R9 VP.n33 VP.n13 161.3
R10 VP.n35 VP.n34 161.3
R11 VP.n36 VP.n12 161.3
R12 VP.n38 VP.n37 161.3
R13 VP.n39 VP.n11 161.3
R14 VP.n72 VP.n0 161.3
R15 VP.n71 VP.n70 161.3
R16 VP.n69 VP.n1 161.3
R17 VP.n68 VP.n67 161.3
R18 VP.n66 VP.n2 161.3
R19 VP.n65 VP.n64 161.3
R20 VP.n63 VP.n62 161.3
R21 VP.n61 VP.n4 161.3
R22 VP.n60 VP.n59 161.3
R23 VP.n58 VP.n5 161.3
R24 VP.n57 VP.n56 161.3
R25 VP.n55 VP.n6 161.3
R26 VP.n54 VP.n53 161.3
R27 VP.n52 VP.n51 161.3
R28 VP.n50 VP.n8 161.3
R29 VP.n49 VP.n48 161.3
R30 VP.n47 VP.n9 161.3
R31 VP.n46 VP.n45 161.3
R32 VP.n44 VP.n10 161.3
R33 VP.n43 VP.t6 156.739
R34 VP.n7 VP.t4 156.739
R35 VP.n3 VP.t1 156.739
R36 VP.n73 VP.t5 156.739
R37 VP.n40 VP.t3 156.739
R38 VP.n14 VP.t2 156.739
R39 VP.n18 VP.t0 156.739
R40 VP.n43 VP.n42 108.695
R41 VP.n74 VP.n73 108.695
R42 VP.n41 VP.n40 108.695
R43 VP.n19 VP.n18 72.8488
R44 VP.n42 VP.n41 55.4997
R45 VP.n49 VP.n9 43.4833
R46 VP.n67 VP.n1 43.4833
R47 VP.n34 VP.n12 43.4833
R48 VP.n56 VP.n5 40.577
R49 VP.n60 VP.n5 40.577
R50 VP.n27 VP.n16 40.577
R51 VP.n23 VP.n16 40.577
R52 VP.n50 VP.n49 37.6707
R53 VP.n67 VP.n66 37.6707
R54 VP.n34 VP.n33 37.6707
R55 VP.n45 VP.n44 24.5923
R56 VP.n45 VP.n9 24.5923
R57 VP.n51 VP.n50 24.5923
R58 VP.n55 VP.n54 24.5923
R59 VP.n56 VP.n55 24.5923
R60 VP.n61 VP.n60 24.5923
R61 VP.n62 VP.n61 24.5923
R62 VP.n66 VP.n65 24.5923
R63 VP.n71 VP.n1 24.5923
R64 VP.n72 VP.n71 24.5923
R65 VP.n38 VP.n12 24.5923
R66 VP.n39 VP.n38 24.5923
R67 VP.n28 VP.n27 24.5923
R68 VP.n29 VP.n28 24.5923
R69 VP.n33 VP.n32 24.5923
R70 VP.n22 VP.n21 24.5923
R71 VP.n23 VP.n22 24.5923
R72 VP.n51 VP.n7 23.8546
R73 VP.n65 VP.n3 23.8546
R74 VP.n32 VP.n14 23.8546
R75 VP.n20 VP.n19 7.34013
R76 VP.n44 VP.n43 2.21377
R77 VP.n73 VP.n72 2.21377
R78 VP.n40 VP.n39 2.21377
R79 VP.n54 VP.n7 0.738255
R80 VP.n62 VP.n3 0.738255
R81 VP.n29 VP.n14 0.738255
R82 VP.n21 VP.n18 0.738255
R83 VP.n41 VP.n11 0.278335
R84 VP.n42 VP.n10 0.278335
R85 VP.n74 VP.n0 0.278335
R86 VP.n20 VP.n17 0.189894
R87 VP.n24 VP.n17 0.189894
R88 VP.n25 VP.n24 0.189894
R89 VP.n26 VP.n25 0.189894
R90 VP.n26 VP.n15 0.189894
R91 VP.n30 VP.n15 0.189894
R92 VP.n31 VP.n30 0.189894
R93 VP.n31 VP.n13 0.189894
R94 VP.n35 VP.n13 0.189894
R95 VP.n36 VP.n35 0.189894
R96 VP.n37 VP.n36 0.189894
R97 VP.n37 VP.n11 0.189894
R98 VP.n46 VP.n10 0.189894
R99 VP.n47 VP.n46 0.189894
R100 VP.n48 VP.n47 0.189894
R101 VP.n48 VP.n8 0.189894
R102 VP.n52 VP.n8 0.189894
R103 VP.n53 VP.n52 0.189894
R104 VP.n53 VP.n6 0.189894
R105 VP.n57 VP.n6 0.189894
R106 VP.n58 VP.n57 0.189894
R107 VP.n59 VP.n58 0.189894
R108 VP.n59 VP.n4 0.189894
R109 VP.n63 VP.n4 0.189894
R110 VP.n64 VP.n63 0.189894
R111 VP.n64 VP.n2 0.189894
R112 VP.n68 VP.n2 0.189894
R113 VP.n69 VP.n68 0.189894
R114 VP.n70 VP.n69 0.189894
R115 VP.n70 VP.n0 0.189894
R116 VP VP.n74 0.153485
R117 VTAIL.n786 VTAIL.n694 756.745
R118 VTAIL.n94 VTAIL.n2 756.745
R119 VTAIL.n192 VTAIL.n100 756.745
R120 VTAIL.n292 VTAIL.n200 756.745
R121 VTAIL.n688 VTAIL.n596 756.745
R122 VTAIL.n588 VTAIL.n496 756.745
R123 VTAIL.n490 VTAIL.n398 756.745
R124 VTAIL.n390 VTAIL.n298 756.745
R125 VTAIL.n727 VTAIL.n726 585
R126 VTAIL.n729 VTAIL.n728 585
R127 VTAIL.n722 VTAIL.n721 585
R128 VTAIL.n735 VTAIL.n734 585
R129 VTAIL.n737 VTAIL.n736 585
R130 VTAIL.n718 VTAIL.n717 585
R131 VTAIL.n743 VTAIL.n742 585
R132 VTAIL.n745 VTAIL.n744 585
R133 VTAIL.n714 VTAIL.n713 585
R134 VTAIL.n751 VTAIL.n750 585
R135 VTAIL.n753 VTAIL.n752 585
R136 VTAIL.n710 VTAIL.n709 585
R137 VTAIL.n759 VTAIL.n758 585
R138 VTAIL.n761 VTAIL.n760 585
R139 VTAIL.n706 VTAIL.n705 585
R140 VTAIL.n768 VTAIL.n767 585
R141 VTAIL.n769 VTAIL.n704 585
R142 VTAIL.n771 VTAIL.n770 585
R143 VTAIL.n702 VTAIL.n701 585
R144 VTAIL.n777 VTAIL.n776 585
R145 VTAIL.n779 VTAIL.n778 585
R146 VTAIL.n698 VTAIL.n697 585
R147 VTAIL.n785 VTAIL.n784 585
R148 VTAIL.n787 VTAIL.n786 585
R149 VTAIL.n35 VTAIL.n34 585
R150 VTAIL.n37 VTAIL.n36 585
R151 VTAIL.n30 VTAIL.n29 585
R152 VTAIL.n43 VTAIL.n42 585
R153 VTAIL.n45 VTAIL.n44 585
R154 VTAIL.n26 VTAIL.n25 585
R155 VTAIL.n51 VTAIL.n50 585
R156 VTAIL.n53 VTAIL.n52 585
R157 VTAIL.n22 VTAIL.n21 585
R158 VTAIL.n59 VTAIL.n58 585
R159 VTAIL.n61 VTAIL.n60 585
R160 VTAIL.n18 VTAIL.n17 585
R161 VTAIL.n67 VTAIL.n66 585
R162 VTAIL.n69 VTAIL.n68 585
R163 VTAIL.n14 VTAIL.n13 585
R164 VTAIL.n76 VTAIL.n75 585
R165 VTAIL.n77 VTAIL.n12 585
R166 VTAIL.n79 VTAIL.n78 585
R167 VTAIL.n10 VTAIL.n9 585
R168 VTAIL.n85 VTAIL.n84 585
R169 VTAIL.n87 VTAIL.n86 585
R170 VTAIL.n6 VTAIL.n5 585
R171 VTAIL.n93 VTAIL.n92 585
R172 VTAIL.n95 VTAIL.n94 585
R173 VTAIL.n133 VTAIL.n132 585
R174 VTAIL.n135 VTAIL.n134 585
R175 VTAIL.n128 VTAIL.n127 585
R176 VTAIL.n141 VTAIL.n140 585
R177 VTAIL.n143 VTAIL.n142 585
R178 VTAIL.n124 VTAIL.n123 585
R179 VTAIL.n149 VTAIL.n148 585
R180 VTAIL.n151 VTAIL.n150 585
R181 VTAIL.n120 VTAIL.n119 585
R182 VTAIL.n157 VTAIL.n156 585
R183 VTAIL.n159 VTAIL.n158 585
R184 VTAIL.n116 VTAIL.n115 585
R185 VTAIL.n165 VTAIL.n164 585
R186 VTAIL.n167 VTAIL.n166 585
R187 VTAIL.n112 VTAIL.n111 585
R188 VTAIL.n174 VTAIL.n173 585
R189 VTAIL.n175 VTAIL.n110 585
R190 VTAIL.n177 VTAIL.n176 585
R191 VTAIL.n108 VTAIL.n107 585
R192 VTAIL.n183 VTAIL.n182 585
R193 VTAIL.n185 VTAIL.n184 585
R194 VTAIL.n104 VTAIL.n103 585
R195 VTAIL.n191 VTAIL.n190 585
R196 VTAIL.n193 VTAIL.n192 585
R197 VTAIL.n233 VTAIL.n232 585
R198 VTAIL.n235 VTAIL.n234 585
R199 VTAIL.n228 VTAIL.n227 585
R200 VTAIL.n241 VTAIL.n240 585
R201 VTAIL.n243 VTAIL.n242 585
R202 VTAIL.n224 VTAIL.n223 585
R203 VTAIL.n249 VTAIL.n248 585
R204 VTAIL.n251 VTAIL.n250 585
R205 VTAIL.n220 VTAIL.n219 585
R206 VTAIL.n257 VTAIL.n256 585
R207 VTAIL.n259 VTAIL.n258 585
R208 VTAIL.n216 VTAIL.n215 585
R209 VTAIL.n265 VTAIL.n264 585
R210 VTAIL.n267 VTAIL.n266 585
R211 VTAIL.n212 VTAIL.n211 585
R212 VTAIL.n274 VTAIL.n273 585
R213 VTAIL.n275 VTAIL.n210 585
R214 VTAIL.n277 VTAIL.n276 585
R215 VTAIL.n208 VTAIL.n207 585
R216 VTAIL.n283 VTAIL.n282 585
R217 VTAIL.n285 VTAIL.n284 585
R218 VTAIL.n204 VTAIL.n203 585
R219 VTAIL.n291 VTAIL.n290 585
R220 VTAIL.n293 VTAIL.n292 585
R221 VTAIL.n689 VTAIL.n688 585
R222 VTAIL.n687 VTAIL.n686 585
R223 VTAIL.n600 VTAIL.n599 585
R224 VTAIL.n681 VTAIL.n680 585
R225 VTAIL.n679 VTAIL.n678 585
R226 VTAIL.n604 VTAIL.n603 585
R227 VTAIL.n608 VTAIL.n606 585
R228 VTAIL.n673 VTAIL.n672 585
R229 VTAIL.n671 VTAIL.n670 585
R230 VTAIL.n610 VTAIL.n609 585
R231 VTAIL.n665 VTAIL.n664 585
R232 VTAIL.n663 VTAIL.n662 585
R233 VTAIL.n614 VTAIL.n613 585
R234 VTAIL.n657 VTAIL.n656 585
R235 VTAIL.n655 VTAIL.n654 585
R236 VTAIL.n618 VTAIL.n617 585
R237 VTAIL.n649 VTAIL.n648 585
R238 VTAIL.n647 VTAIL.n646 585
R239 VTAIL.n622 VTAIL.n621 585
R240 VTAIL.n641 VTAIL.n640 585
R241 VTAIL.n639 VTAIL.n638 585
R242 VTAIL.n626 VTAIL.n625 585
R243 VTAIL.n633 VTAIL.n632 585
R244 VTAIL.n631 VTAIL.n630 585
R245 VTAIL.n589 VTAIL.n588 585
R246 VTAIL.n587 VTAIL.n586 585
R247 VTAIL.n500 VTAIL.n499 585
R248 VTAIL.n581 VTAIL.n580 585
R249 VTAIL.n579 VTAIL.n578 585
R250 VTAIL.n504 VTAIL.n503 585
R251 VTAIL.n508 VTAIL.n506 585
R252 VTAIL.n573 VTAIL.n572 585
R253 VTAIL.n571 VTAIL.n570 585
R254 VTAIL.n510 VTAIL.n509 585
R255 VTAIL.n565 VTAIL.n564 585
R256 VTAIL.n563 VTAIL.n562 585
R257 VTAIL.n514 VTAIL.n513 585
R258 VTAIL.n557 VTAIL.n556 585
R259 VTAIL.n555 VTAIL.n554 585
R260 VTAIL.n518 VTAIL.n517 585
R261 VTAIL.n549 VTAIL.n548 585
R262 VTAIL.n547 VTAIL.n546 585
R263 VTAIL.n522 VTAIL.n521 585
R264 VTAIL.n541 VTAIL.n540 585
R265 VTAIL.n539 VTAIL.n538 585
R266 VTAIL.n526 VTAIL.n525 585
R267 VTAIL.n533 VTAIL.n532 585
R268 VTAIL.n531 VTAIL.n530 585
R269 VTAIL.n491 VTAIL.n490 585
R270 VTAIL.n489 VTAIL.n488 585
R271 VTAIL.n402 VTAIL.n401 585
R272 VTAIL.n483 VTAIL.n482 585
R273 VTAIL.n481 VTAIL.n480 585
R274 VTAIL.n406 VTAIL.n405 585
R275 VTAIL.n410 VTAIL.n408 585
R276 VTAIL.n475 VTAIL.n474 585
R277 VTAIL.n473 VTAIL.n472 585
R278 VTAIL.n412 VTAIL.n411 585
R279 VTAIL.n467 VTAIL.n466 585
R280 VTAIL.n465 VTAIL.n464 585
R281 VTAIL.n416 VTAIL.n415 585
R282 VTAIL.n459 VTAIL.n458 585
R283 VTAIL.n457 VTAIL.n456 585
R284 VTAIL.n420 VTAIL.n419 585
R285 VTAIL.n451 VTAIL.n450 585
R286 VTAIL.n449 VTAIL.n448 585
R287 VTAIL.n424 VTAIL.n423 585
R288 VTAIL.n443 VTAIL.n442 585
R289 VTAIL.n441 VTAIL.n440 585
R290 VTAIL.n428 VTAIL.n427 585
R291 VTAIL.n435 VTAIL.n434 585
R292 VTAIL.n433 VTAIL.n432 585
R293 VTAIL.n391 VTAIL.n390 585
R294 VTAIL.n389 VTAIL.n388 585
R295 VTAIL.n302 VTAIL.n301 585
R296 VTAIL.n383 VTAIL.n382 585
R297 VTAIL.n381 VTAIL.n380 585
R298 VTAIL.n306 VTAIL.n305 585
R299 VTAIL.n310 VTAIL.n308 585
R300 VTAIL.n375 VTAIL.n374 585
R301 VTAIL.n373 VTAIL.n372 585
R302 VTAIL.n312 VTAIL.n311 585
R303 VTAIL.n367 VTAIL.n366 585
R304 VTAIL.n365 VTAIL.n364 585
R305 VTAIL.n316 VTAIL.n315 585
R306 VTAIL.n359 VTAIL.n358 585
R307 VTAIL.n357 VTAIL.n356 585
R308 VTAIL.n320 VTAIL.n319 585
R309 VTAIL.n351 VTAIL.n350 585
R310 VTAIL.n349 VTAIL.n348 585
R311 VTAIL.n324 VTAIL.n323 585
R312 VTAIL.n343 VTAIL.n342 585
R313 VTAIL.n341 VTAIL.n340 585
R314 VTAIL.n328 VTAIL.n327 585
R315 VTAIL.n335 VTAIL.n334 585
R316 VTAIL.n333 VTAIL.n332 585
R317 VTAIL.n725 VTAIL.t0 327.466
R318 VTAIL.n33 VTAIL.t2 327.466
R319 VTAIL.n131 VTAIL.t13 327.466
R320 VTAIL.n231 VTAIL.t15 327.466
R321 VTAIL.n629 VTAIL.t12 327.466
R322 VTAIL.n529 VTAIL.t10 327.466
R323 VTAIL.n431 VTAIL.t1 327.466
R324 VTAIL.n331 VTAIL.t5 327.466
R325 VTAIL.n728 VTAIL.n727 171.744
R326 VTAIL.n728 VTAIL.n721 171.744
R327 VTAIL.n735 VTAIL.n721 171.744
R328 VTAIL.n736 VTAIL.n735 171.744
R329 VTAIL.n736 VTAIL.n717 171.744
R330 VTAIL.n743 VTAIL.n717 171.744
R331 VTAIL.n744 VTAIL.n743 171.744
R332 VTAIL.n744 VTAIL.n713 171.744
R333 VTAIL.n751 VTAIL.n713 171.744
R334 VTAIL.n752 VTAIL.n751 171.744
R335 VTAIL.n752 VTAIL.n709 171.744
R336 VTAIL.n759 VTAIL.n709 171.744
R337 VTAIL.n760 VTAIL.n759 171.744
R338 VTAIL.n760 VTAIL.n705 171.744
R339 VTAIL.n768 VTAIL.n705 171.744
R340 VTAIL.n769 VTAIL.n768 171.744
R341 VTAIL.n770 VTAIL.n769 171.744
R342 VTAIL.n770 VTAIL.n701 171.744
R343 VTAIL.n777 VTAIL.n701 171.744
R344 VTAIL.n778 VTAIL.n777 171.744
R345 VTAIL.n778 VTAIL.n697 171.744
R346 VTAIL.n785 VTAIL.n697 171.744
R347 VTAIL.n786 VTAIL.n785 171.744
R348 VTAIL.n36 VTAIL.n35 171.744
R349 VTAIL.n36 VTAIL.n29 171.744
R350 VTAIL.n43 VTAIL.n29 171.744
R351 VTAIL.n44 VTAIL.n43 171.744
R352 VTAIL.n44 VTAIL.n25 171.744
R353 VTAIL.n51 VTAIL.n25 171.744
R354 VTAIL.n52 VTAIL.n51 171.744
R355 VTAIL.n52 VTAIL.n21 171.744
R356 VTAIL.n59 VTAIL.n21 171.744
R357 VTAIL.n60 VTAIL.n59 171.744
R358 VTAIL.n60 VTAIL.n17 171.744
R359 VTAIL.n67 VTAIL.n17 171.744
R360 VTAIL.n68 VTAIL.n67 171.744
R361 VTAIL.n68 VTAIL.n13 171.744
R362 VTAIL.n76 VTAIL.n13 171.744
R363 VTAIL.n77 VTAIL.n76 171.744
R364 VTAIL.n78 VTAIL.n77 171.744
R365 VTAIL.n78 VTAIL.n9 171.744
R366 VTAIL.n85 VTAIL.n9 171.744
R367 VTAIL.n86 VTAIL.n85 171.744
R368 VTAIL.n86 VTAIL.n5 171.744
R369 VTAIL.n93 VTAIL.n5 171.744
R370 VTAIL.n94 VTAIL.n93 171.744
R371 VTAIL.n134 VTAIL.n133 171.744
R372 VTAIL.n134 VTAIL.n127 171.744
R373 VTAIL.n141 VTAIL.n127 171.744
R374 VTAIL.n142 VTAIL.n141 171.744
R375 VTAIL.n142 VTAIL.n123 171.744
R376 VTAIL.n149 VTAIL.n123 171.744
R377 VTAIL.n150 VTAIL.n149 171.744
R378 VTAIL.n150 VTAIL.n119 171.744
R379 VTAIL.n157 VTAIL.n119 171.744
R380 VTAIL.n158 VTAIL.n157 171.744
R381 VTAIL.n158 VTAIL.n115 171.744
R382 VTAIL.n165 VTAIL.n115 171.744
R383 VTAIL.n166 VTAIL.n165 171.744
R384 VTAIL.n166 VTAIL.n111 171.744
R385 VTAIL.n174 VTAIL.n111 171.744
R386 VTAIL.n175 VTAIL.n174 171.744
R387 VTAIL.n176 VTAIL.n175 171.744
R388 VTAIL.n176 VTAIL.n107 171.744
R389 VTAIL.n183 VTAIL.n107 171.744
R390 VTAIL.n184 VTAIL.n183 171.744
R391 VTAIL.n184 VTAIL.n103 171.744
R392 VTAIL.n191 VTAIL.n103 171.744
R393 VTAIL.n192 VTAIL.n191 171.744
R394 VTAIL.n234 VTAIL.n233 171.744
R395 VTAIL.n234 VTAIL.n227 171.744
R396 VTAIL.n241 VTAIL.n227 171.744
R397 VTAIL.n242 VTAIL.n241 171.744
R398 VTAIL.n242 VTAIL.n223 171.744
R399 VTAIL.n249 VTAIL.n223 171.744
R400 VTAIL.n250 VTAIL.n249 171.744
R401 VTAIL.n250 VTAIL.n219 171.744
R402 VTAIL.n257 VTAIL.n219 171.744
R403 VTAIL.n258 VTAIL.n257 171.744
R404 VTAIL.n258 VTAIL.n215 171.744
R405 VTAIL.n265 VTAIL.n215 171.744
R406 VTAIL.n266 VTAIL.n265 171.744
R407 VTAIL.n266 VTAIL.n211 171.744
R408 VTAIL.n274 VTAIL.n211 171.744
R409 VTAIL.n275 VTAIL.n274 171.744
R410 VTAIL.n276 VTAIL.n275 171.744
R411 VTAIL.n276 VTAIL.n207 171.744
R412 VTAIL.n283 VTAIL.n207 171.744
R413 VTAIL.n284 VTAIL.n283 171.744
R414 VTAIL.n284 VTAIL.n203 171.744
R415 VTAIL.n291 VTAIL.n203 171.744
R416 VTAIL.n292 VTAIL.n291 171.744
R417 VTAIL.n688 VTAIL.n687 171.744
R418 VTAIL.n687 VTAIL.n599 171.744
R419 VTAIL.n680 VTAIL.n599 171.744
R420 VTAIL.n680 VTAIL.n679 171.744
R421 VTAIL.n679 VTAIL.n603 171.744
R422 VTAIL.n608 VTAIL.n603 171.744
R423 VTAIL.n672 VTAIL.n608 171.744
R424 VTAIL.n672 VTAIL.n671 171.744
R425 VTAIL.n671 VTAIL.n609 171.744
R426 VTAIL.n664 VTAIL.n609 171.744
R427 VTAIL.n664 VTAIL.n663 171.744
R428 VTAIL.n663 VTAIL.n613 171.744
R429 VTAIL.n656 VTAIL.n613 171.744
R430 VTAIL.n656 VTAIL.n655 171.744
R431 VTAIL.n655 VTAIL.n617 171.744
R432 VTAIL.n648 VTAIL.n617 171.744
R433 VTAIL.n648 VTAIL.n647 171.744
R434 VTAIL.n647 VTAIL.n621 171.744
R435 VTAIL.n640 VTAIL.n621 171.744
R436 VTAIL.n640 VTAIL.n639 171.744
R437 VTAIL.n639 VTAIL.n625 171.744
R438 VTAIL.n632 VTAIL.n625 171.744
R439 VTAIL.n632 VTAIL.n631 171.744
R440 VTAIL.n588 VTAIL.n587 171.744
R441 VTAIL.n587 VTAIL.n499 171.744
R442 VTAIL.n580 VTAIL.n499 171.744
R443 VTAIL.n580 VTAIL.n579 171.744
R444 VTAIL.n579 VTAIL.n503 171.744
R445 VTAIL.n508 VTAIL.n503 171.744
R446 VTAIL.n572 VTAIL.n508 171.744
R447 VTAIL.n572 VTAIL.n571 171.744
R448 VTAIL.n571 VTAIL.n509 171.744
R449 VTAIL.n564 VTAIL.n509 171.744
R450 VTAIL.n564 VTAIL.n563 171.744
R451 VTAIL.n563 VTAIL.n513 171.744
R452 VTAIL.n556 VTAIL.n513 171.744
R453 VTAIL.n556 VTAIL.n555 171.744
R454 VTAIL.n555 VTAIL.n517 171.744
R455 VTAIL.n548 VTAIL.n517 171.744
R456 VTAIL.n548 VTAIL.n547 171.744
R457 VTAIL.n547 VTAIL.n521 171.744
R458 VTAIL.n540 VTAIL.n521 171.744
R459 VTAIL.n540 VTAIL.n539 171.744
R460 VTAIL.n539 VTAIL.n525 171.744
R461 VTAIL.n532 VTAIL.n525 171.744
R462 VTAIL.n532 VTAIL.n531 171.744
R463 VTAIL.n490 VTAIL.n489 171.744
R464 VTAIL.n489 VTAIL.n401 171.744
R465 VTAIL.n482 VTAIL.n401 171.744
R466 VTAIL.n482 VTAIL.n481 171.744
R467 VTAIL.n481 VTAIL.n405 171.744
R468 VTAIL.n410 VTAIL.n405 171.744
R469 VTAIL.n474 VTAIL.n410 171.744
R470 VTAIL.n474 VTAIL.n473 171.744
R471 VTAIL.n473 VTAIL.n411 171.744
R472 VTAIL.n466 VTAIL.n411 171.744
R473 VTAIL.n466 VTAIL.n465 171.744
R474 VTAIL.n465 VTAIL.n415 171.744
R475 VTAIL.n458 VTAIL.n415 171.744
R476 VTAIL.n458 VTAIL.n457 171.744
R477 VTAIL.n457 VTAIL.n419 171.744
R478 VTAIL.n450 VTAIL.n419 171.744
R479 VTAIL.n450 VTAIL.n449 171.744
R480 VTAIL.n449 VTAIL.n423 171.744
R481 VTAIL.n442 VTAIL.n423 171.744
R482 VTAIL.n442 VTAIL.n441 171.744
R483 VTAIL.n441 VTAIL.n427 171.744
R484 VTAIL.n434 VTAIL.n427 171.744
R485 VTAIL.n434 VTAIL.n433 171.744
R486 VTAIL.n390 VTAIL.n389 171.744
R487 VTAIL.n389 VTAIL.n301 171.744
R488 VTAIL.n382 VTAIL.n301 171.744
R489 VTAIL.n382 VTAIL.n381 171.744
R490 VTAIL.n381 VTAIL.n305 171.744
R491 VTAIL.n310 VTAIL.n305 171.744
R492 VTAIL.n374 VTAIL.n310 171.744
R493 VTAIL.n374 VTAIL.n373 171.744
R494 VTAIL.n373 VTAIL.n311 171.744
R495 VTAIL.n366 VTAIL.n311 171.744
R496 VTAIL.n366 VTAIL.n365 171.744
R497 VTAIL.n365 VTAIL.n315 171.744
R498 VTAIL.n358 VTAIL.n315 171.744
R499 VTAIL.n358 VTAIL.n357 171.744
R500 VTAIL.n357 VTAIL.n319 171.744
R501 VTAIL.n350 VTAIL.n319 171.744
R502 VTAIL.n350 VTAIL.n349 171.744
R503 VTAIL.n349 VTAIL.n323 171.744
R504 VTAIL.n342 VTAIL.n323 171.744
R505 VTAIL.n342 VTAIL.n341 171.744
R506 VTAIL.n341 VTAIL.n327 171.744
R507 VTAIL.n334 VTAIL.n327 171.744
R508 VTAIL.n334 VTAIL.n333 171.744
R509 VTAIL.n727 VTAIL.t0 85.8723
R510 VTAIL.n35 VTAIL.t2 85.8723
R511 VTAIL.n133 VTAIL.t13 85.8723
R512 VTAIL.n233 VTAIL.t15 85.8723
R513 VTAIL.n631 VTAIL.t12 85.8723
R514 VTAIL.n531 VTAIL.t10 85.8723
R515 VTAIL.n433 VTAIL.t1 85.8723
R516 VTAIL.n333 VTAIL.t5 85.8723
R517 VTAIL.n595 VTAIL.n594 53.1192
R518 VTAIL.n397 VTAIL.n396 53.1192
R519 VTAIL.n1 VTAIL.n0 53.119
R520 VTAIL.n199 VTAIL.n198 53.119
R521 VTAIL.n791 VTAIL.n790 32.9611
R522 VTAIL.n99 VTAIL.n98 32.9611
R523 VTAIL.n197 VTAIL.n196 32.9611
R524 VTAIL.n297 VTAIL.n296 32.9611
R525 VTAIL.n693 VTAIL.n692 32.9611
R526 VTAIL.n593 VTAIL.n592 32.9611
R527 VTAIL.n495 VTAIL.n494 32.9611
R528 VTAIL.n395 VTAIL.n394 32.9611
R529 VTAIL.n791 VTAIL.n693 30.1169
R530 VTAIL.n395 VTAIL.n297 30.1169
R531 VTAIL.n726 VTAIL.n725 16.3895
R532 VTAIL.n34 VTAIL.n33 16.3895
R533 VTAIL.n132 VTAIL.n131 16.3895
R534 VTAIL.n232 VTAIL.n231 16.3895
R535 VTAIL.n630 VTAIL.n629 16.3895
R536 VTAIL.n530 VTAIL.n529 16.3895
R537 VTAIL.n432 VTAIL.n431 16.3895
R538 VTAIL.n332 VTAIL.n331 16.3895
R539 VTAIL.n771 VTAIL.n702 13.1884
R540 VTAIL.n79 VTAIL.n10 13.1884
R541 VTAIL.n177 VTAIL.n108 13.1884
R542 VTAIL.n277 VTAIL.n208 13.1884
R543 VTAIL.n606 VTAIL.n604 13.1884
R544 VTAIL.n506 VTAIL.n504 13.1884
R545 VTAIL.n408 VTAIL.n406 13.1884
R546 VTAIL.n308 VTAIL.n306 13.1884
R547 VTAIL.n729 VTAIL.n724 12.8005
R548 VTAIL.n772 VTAIL.n704 12.8005
R549 VTAIL.n776 VTAIL.n775 12.8005
R550 VTAIL.n37 VTAIL.n32 12.8005
R551 VTAIL.n80 VTAIL.n12 12.8005
R552 VTAIL.n84 VTAIL.n83 12.8005
R553 VTAIL.n135 VTAIL.n130 12.8005
R554 VTAIL.n178 VTAIL.n110 12.8005
R555 VTAIL.n182 VTAIL.n181 12.8005
R556 VTAIL.n235 VTAIL.n230 12.8005
R557 VTAIL.n278 VTAIL.n210 12.8005
R558 VTAIL.n282 VTAIL.n281 12.8005
R559 VTAIL.n678 VTAIL.n677 12.8005
R560 VTAIL.n674 VTAIL.n673 12.8005
R561 VTAIL.n633 VTAIL.n628 12.8005
R562 VTAIL.n578 VTAIL.n577 12.8005
R563 VTAIL.n574 VTAIL.n573 12.8005
R564 VTAIL.n533 VTAIL.n528 12.8005
R565 VTAIL.n480 VTAIL.n479 12.8005
R566 VTAIL.n476 VTAIL.n475 12.8005
R567 VTAIL.n435 VTAIL.n430 12.8005
R568 VTAIL.n380 VTAIL.n379 12.8005
R569 VTAIL.n376 VTAIL.n375 12.8005
R570 VTAIL.n335 VTAIL.n330 12.8005
R571 VTAIL.n730 VTAIL.n722 12.0247
R572 VTAIL.n767 VTAIL.n766 12.0247
R573 VTAIL.n779 VTAIL.n700 12.0247
R574 VTAIL.n38 VTAIL.n30 12.0247
R575 VTAIL.n75 VTAIL.n74 12.0247
R576 VTAIL.n87 VTAIL.n8 12.0247
R577 VTAIL.n136 VTAIL.n128 12.0247
R578 VTAIL.n173 VTAIL.n172 12.0247
R579 VTAIL.n185 VTAIL.n106 12.0247
R580 VTAIL.n236 VTAIL.n228 12.0247
R581 VTAIL.n273 VTAIL.n272 12.0247
R582 VTAIL.n285 VTAIL.n206 12.0247
R583 VTAIL.n681 VTAIL.n602 12.0247
R584 VTAIL.n670 VTAIL.n607 12.0247
R585 VTAIL.n634 VTAIL.n626 12.0247
R586 VTAIL.n581 VTAIL.n502 12.0247
R587 VTAIL.n570 VTAIL.n507 12.0247
R588 VTAIL.n534 VTAIL.n526 12.0247
R589 VTAIL.n483 VTAIL.n404 12.0247
R590 VTAIL.n472 VTAIL.n409 12.0247
R591 VTAIL.n436 VTAIL.n428 12.0247
R592 VTAIL.n383 VTAIL.n304 12.0247
R593 VTAIL.n372 VTAIL.n309 12.0247
R594 VTAIL.n336 VTAIL.n328 12.0247
R595 VTAIL.n734 VTAIL.n733 11.249
R596 VTAIL.n765 VTAIL.n706 11.249
R597 VTAIL.n780 VTAIL.n698 11.249
R598 VTAIL.n42 VTAIL.n41 11.249
R599 VTAIL.n73 VTAIL.n14 11.249
R600 VTAIL.n88 VTAIL.n6 11.249
R601 VTAIL.n140 VTAIL.n139 11.249
R602 VTAIL.n171 VTAIL.n112 11.249
R603 VTAIL.n186 VTAIL.n104 11.249
R604 VTAIL.n240 VTAIL.n239 11.249
R605 VTAIL.n271 VTAIL.n212 11.249
R606 VTAIL.n286 VTAIL.n204 11.249
R607 VTAIL.n682 VTAIL.n600 11.249
R608 VTAIL.n669 VTAIL.n610 11.249
R609 VTAIL.n638 VTAIL.n637 11.249
R610 VTAIL.n582 VTAIL.n500 11.249
R611 VTAIL.n569 VTAIL.n510 11.249
R612 VTAIL.n538 VTAIL.n537 11.249
R613 VTAIL.n484 VTAIL.n402 11.249
R614 VTAIL.n471 VTAIL.n412 11.249
R615 VTAIL.n440 VTAIL.n439 11.249
R616 VTAIL.n384 VTAIL.n302 11.249
R617 VTAIL.n371 VTAIL.n312 11.249
R618 VTAIL.n340 VTAIL.n339 11.249
R619 VTAIL.n737 VTAIL.n720 10.4732
R620 VTAIL.n762 VTAIL.n761 10.4732
R621 VTAIL.n784 VTAIL.n783 10.4732
R622 VTAIL.n45 VTAIL.n28 10.4732
R623 VTAIL.n70 VTAIL.n69 10.4732
R624 VTAIL.n92 VTAIL.n91 10.4732
R625 VTAIL.n143 VTAIL.n126 10.4732
R626 VTAIL.n168 VTAIL.n167 10.4732
R627 VTAIL.n190 VTAIL.n189 10.4732
R628 VTAIL.n243 VTAIL.n226 10.4732
R629 VTAIL.n268 VTAIL.n267 10.4732
R630 VTAIL.n290 VTAIL.n289 10.4732
R631 VTAIL.n686 VTAIL.n685 10.4732
R632 VTAIL.n666 VTAIL.n665 10.4732
R633 VTAIL.n641 VTAIL.n624 10.4732
R634 VTAIL.n586 VTAIL.n585 10.4732
R635 VTAIL.n566 VTAIL.n565 10.4732
R636 VTAIL.n541 VTAIL.n524 10.4732
R637 VTAIL.n488 VTAIL.n487 10.4732
R638 VTAIL.n468 VTAIL.n467 10.4732
R639 VTAIL.n443 VTAIL.n426 10.4732
R640 VTAIL.n388 VTAIL.n387 10.4732
R641 VTAIL.n368 VTAIL.n367 10.4732
R642 VTAIL.n343 VTAIL.n326 10.4732
R643 VTAIL.n738 VTAIL.n718 9.69747
R644 VTAIL.n758 VTAIL.n708 9.69747
R645 VTAIL.n787 VTAIL.n696 9.69747
R646 VTAIL.n46 VTAIL.n26 9.69747
R647 VTAIL.n66 VTAIL.n16 9.69747
R648 VTAIL.n95 VTAIL.n4 9.69747
R649 VTAIL.n144 VTAIL.n124 9.69747
R650 VTAIL.n164 VTAIL.n114 9.69747
R651 VTAIL.n193 VTAIL.n102 9.69747
R652 VTAIL.n244 VTAIL.n224 9.69747
R653 VTAIL.n264 VTAIL.n214 9.69747
R654 VTAIL.n293 VTAIL.n202 9.69747
R655 VTAIL.n689 VTAIL.n598 9.69747
R656 VTAIL.n662 VTAIL.n612 9.69747
R657 VTAIL.n642 VTAIL.n622 9.69747
R658 VTAIL.n589 VTAIL.n498 9.69747
R659 VTAIL.n562 VTAIL.n512 9.69747
R660 VTAIL.n542 VTAIL.n522 9.69747
R661 VTAIL.n491 VTAIL.n400 9.69747
R662 VTAIL.n464 VTAIL.n414 9.69747
R663 VTAIL.n444 VTAIL.n424 9.69747
R664 VTAIL.n391 VTAIL.n300 9.69747
R665 VTAIL.n364 VTAIL.n314 9.69747
R666 VTAIL.n344 VTAIL.n324 9.69747
R667 VTAIL.n790 VTAIL.n789 9.45567
R668 VTAIL.n98 VTAIL.n97 9.45567
R669 VTAIL.n196 VTAIL.n195 9.45567
R670 VTAIL.n296 VTAIL.n295 9.45567
R671 VTAIL.n692 VTAIL.n691 9.45567
R672 VTAIL.n592 VTAIL.n591 9.45567
R673 VTAIL.n494 VTAIL.n493 9.45567
R674 VTAIL.n394 VTAIL.n393 9.45567
R675 VTAIL.n789 VTAIL.n788 9.3005
R676 VTAIL.n696 VTAIL.n695 9.3005
R677 VTAIL.n783 VTAIL.n782 9.3005
R678 VTAIL.n781 VTAIL.n780 9.3005
R679 VTAIL.n700 VTAIL.n699 9.3005
R680 VTAIL.n775 VTAIL.n774 9.3005
R681 VTAIL.n747 VTAIL.n746 9.3005
R682 VTAIL.n716 VTAIL.n715 9.3005
R683 VTAIL.n741 VTAIL.n740 9.3005
R684 VTAIL.n739 VTAIL.n738 9.3005
R685 VTAIL.n720 VTAIL.n719 9.3005
R686 VTAIL.n733 VTAIL.n732 9.3005
R687 VTAIL.n731 VTAIL.n730 9.3005
R688 VTAIL.n724 VTAIL.n723 9.3005
R689 VTAIL.n749 VTAIL.n748 9.3005
R690 VTAIL.n712 VTAIL.n711 9.3005
R691 VTAIL.n755 VTAIL.n754 9.3005
R692 VTAIL.n757 VTAIL.n756 9.3005
R693 VTAIL.n708 VTAIL.n707 9.3005
R694 VTAIL.n763 VTAIL.n762 9.3005
R695 VTAIL.n765 VTAIL.n764 9.3005
R696 VTAIL.n766 VTAIL.n703 9.3005
R697 VTAIL.n773 VTAIL.n772 9.3005
R698 VTAIL.n97 VTAIL.n96 9.3005
R699 VTAIL.n4 VTAIL.n3 9.3005
R700 VTAIL.n91 VTAIL.n90 9.3005
R701 VTAIL.n89 VTAIL.n88 9.3005
R702 VTAIL.n8 VTAIL.n7 9.3005
R703 VTAIL.n83 VTAIL.n82 9.3005
R704 VTAIL.n55 VTAIL.n54 9.3005
R705 VTAIL.n24 VTAIL.n23 9.3005
R706 VTAIL.n49 VTAIL.n48 9.3005
R707 VTAIL.n47 VTAIL.n46 9.3005
R708 VTAIL.n28 VTAIL.n27 9.3005
R709 VTAIL.n41 VTAIL.n40 9.3005
R710 VTAIL.n39 VTAIL.n38 9.3005
R711 VTAIL.n32 VTAIL.n31 9.3005
R712 VTAIL.n57 VTAIL.n56 9.3005
R713 VTAIL.n20 VTAIL.n19 9.3005
R714 VTAIL.n63 VTAIL.n62 9.3005
R715 VTAIL.n65 VTAIL.n64 9.3005
R716 VTAIL.n16 VTAIL.n15 9.3005
R717 VTAIL.n71 VTAIL.n70 9.3005
R718 VTAIL.n73 VTAIL.n72 9.3005
R719 VTAIL.n74 VTAIL.n11 9.3005
R720 VTAIL.n81 VTAIL.n80 9.3005
R721 VTAIL.n195 VTAIL.n194 9.3005
R722 VTAIL.n102 VTAIL.n101 9.3005
R723 VTAIL.n189 VTAIL.n188 9.3005
R724 VTAIL.n187 VTAIL.n186 9.3005
R725 VTAIL.n106 VTAIL.n105 9.3005
R726 VTAIL.n181 VTAIL.n180 9.3005
R727 VTAIL.n153 VTAIL.n152 9.3005
R728 VTAIL.n122 VTAIL.n121 9.3005
R729 VTAIL.n147 VTAIL.n146 9.3005
R730 VTAIL.n145 VTAIL.n144 9.3005
R731 VTAIL.n126 VTAIL.n125 9.3005
R732 VTAIL.n139 VTAIL.n138 9.3005
R733 VTAIL.n137 VTAIL.n136 9.3005
R734 VTAIL.n130 VTAIL.n129 9.3005
R735 VTAIL.n155 VTAIL.n154 9.3005
R736 VTAIL.n118 VTAIL.n117 9.3005
R737 VTAIL.n161 VTAIL.n160 9.3005
R738 VTAIL.n163 VTAIL.n162 9.3005
R739 VTAIL.n114 VTAIL.n113 9.3005
R740 VTAIL.n169 VTAIL.n168 9.3005
R741 VTAIL.n171 VTAIL.n170 9.3005
R742 VTAIL.n172 VTAIL.n109 9.3005
R743 VTAIL.n179 VTAIL.n178 9.3005
R744 VTAIL.n295 VTAIL.n294 9.3005
R745 VTAIL.n202 VTAIL.n201 9.3005
R746 VTAIL.n289 VTAIL.n288 9.3005
R747 VTAIL.n287 VTAIL.n286 9.3005
R748 VTAIL.n206 VTAIL.n205 9.3005
R749 VTAIL.n281 VTAIL.n280 9.3005
R750 VTAIL.n253 VTAIL.n252 9.3005
R751 VTAIL.n222 VTAIL.n221 9.3005
R752 VTAIL.n247 VTAIL.n246 9.3005
R753 VTAIL.n245 VTAIL.n244 9.3005
R754 VTAIL.n226 VTAIL.n225 9.3005
R755 VTAIL.n239 VTAIL.n238 9.3005
R756 VTAIL.n237 VTAIL.n236 9.3005
R757 VTAIL.n230 VTAIL.n229 9.3005
R758 VTAIL.n255 VTAIL.n254 9.3005
R759 VTAIL.n218 VTAIL.n217 9.3005
R760 VTAIL.n261 VTAIL.n260 9.3005
R761 VTAIL.n263 VTAIL.n262 9.3005
R762 VTAIL.n214 VTAIL.n213 9.3005
R763 VTAIL.n269 VTAIL.n268 9.3005
R764 VTAIL.n271 VTAIL.n270 9.3005
R765 VTAIL.n272 VTAIL.n209 9.3005
R766 VTAIL.n279 VTAIL.n278 9.3005
R767 VTAIL.n616 VTAIL.n615 9.3005
R768 VTAIL.n659 VTAIL.n658 9.3005
R769 VTAIL.n661 VTAIL.n660 9.3005
R770 VTAIL.n612 VTAIL.n611 9.3005
R771 VTAIL.n667 VTAIL.n666 9.3005
R772 VTAIL.n669 VTAIL.n668 9.3005
R773 VTAIL.n607 VTAIL.n605 9.3005
R774 VTAIL.n675 VTAIL.n674 9.3005
R775 VTAIL.n691 VTAIL.n690 9.3005
R776 VTAIL.n598 VTAIL.n597 9.3005
R777 VTAIL.n685 VTAIL.n684 9.3005
R778 VTAIL.n683 VTAIL.n682 9.3005
R779 VTAIL.n602 VTAIL.n601 9.3005
R780 VTAIL.n677 VTAIL.n676 9.3005
R781 VTAIL.n653 VTAIL.n652 9.3005
R782 VTAIL.n651 VTAIL.n650 9.3005
R783 VTAIL.n620 VTAIL.n619 9.3005
R784 VTAIL.n645 VTAIL.n644 9.3005
R785 VTAIL.n643 VTAIL.n642 9.3005
R786 VTAIL.n624 VTAIL.n623 9.3005
R787 VTAIL.n637 VTAIL.n636 9.3005
R788 VTAIL.n635 VTAIL.n634 9.3005
R789 VTAIL.n628 VTAIL.n627 9.3005
R790 VTAIL.n516 VTAIL.n515 9.3005
R791 VTAIL.n559 VTAIL.n558 9.3005
R792 VTAIL.n561 VTAIL.n560 9.3005
R793 VTAIL.n512 VTAIL.n511 9.3005
R794 VTAIL.n567 VTAIL.n566 9.3005
R795 VTAIL.n569 VTAIL.n568 9.3005
R796 VTAIL.n507 VTAIL.n505 9.3005
R797 VTAIL.n575 VTAIL.n574 9.3005
R798 VTAIL.n591 VTAIL.n590 9.3005
R799 VTAIL.n498 VTAIL.n497 9.3005
R800 VTAIL.n585 VTAIL.n584 9.3005
R801 VTAIL.n583 VTAIL.n582 9.3005
R802 VTAIL.n502 VTAIL.n501 9.3005
R803 VTAIL.n577 VTAIL.n576 9.3005
R804 VTAIL.n553 VTAIL.n552 9.3005
R805 VTAIL.n551 VTAIL.n550 9.3005
R806 VTAIL.n520 VTAIL.n519 9.3005
R807 VTAIL.n545 VTAIL.n544 9.3005
R808 VTAIL.n543 VTAIL.n542 9.3005
R809 VTAIL.n524 VTAIL.n523 9.3005
R810 VTAIL.n537 VTAIL.n536 9.3005
R811 VTAIL.n535 VTAIL.n534 9.3005
R812 VTAIL.n528 VTAIL.n527 9.3005
R813 VTAIL.n418 VTAIL.n417 9.3005
R814 VTAIL.n461 VTAIL.n460 9.3005
R815 VTAIL.n463 VTAIL.n462 9.3005
R816 VTAIL.n414 VTAIL.n413 9.3005
R817 VTAIL.n469 VTAIL.n468 9.3005
R818 VTAIL.n471 VTAIL.n470 9.3005
R819 VTAIL.n409 VTAIL.n407 9.3005
R820 VTAIL.n477 VTAIL.n476 9.3005
R821 VTAIL.n493 VTAIL.n492 9.3005
R822 VTAIL.n400 VTAIL.n399 9.3005
R823 VTAIL.n487 VTAIL.n486 9.3005
R824 VTAIL.n485 VTAIL.n484 9.3005
R825 VTAIL.n404 VTAIL.n403 9.3005
R826 VTAIL.n479 VTAIL.n478 9.3005
R827 VTAIL.n455 VTAIL.n454 9.3005
R828 VTAIL.n453 VTAIL.n452 9.3005
R829 VTAIL.n422 VTAIL.n421 9.3005
R830 VTAIL.n447 VTAIL.n446 9.3005
R831 VTAIL.n445 VTAIL.n444 9.3005
R832 VTAIL.n426 VTAIL.n425 9.3005
R833 VTAIL.n439 VTAIL.n438 9.3005
R834 VTAIL.n437 VTAIL.n436 9.3005
R835 VTAIL.n430 VTAIL.n429 9.3005
R836 VTAIL.n318 VTAIL.n317 9.3005
R837 VTAIL.n361 VTAIL.n360 9.3005
R838 VTAIL.n363 VTAIL.n362 9.3005
R839 VTAIL.n314 VTAIL.n313 9.3005
R840 VTAIL.n369 VTAIL.n368 9.3005
R841 VTAIL.n371 VTAIL.n370 9.3005
R842 VTAIL.n309 VTAIL.n307 9.3005
R843 VTAIL.n377 VTAIL.n376 9.3005
R844 VTAIL.n393 VTAIL.n392 9.3005
R845 VTAIL.n300 VTAIL.n299 9.3005
R846 VTAIL.n387 VTAIL.n386 9.3005
R847 VTAIL.n385 VTAIL.n384 9.3005
R848 VTAIL.n304 VTAIL.n303 9.3005
R849 VTAIL.n379 VTAIL.n378 9.3005
R850 VTAIL.n355 VTAIL.n354 9.3005
R851 VTAIL.n353 VTAIL.n352 9.3005
R852 VTAIL.n322 VTAIL.n321 9.3005
R853 VTAIL.n347 VTAIL.n346 9.3005
R854 VTAIL.n345 VTAIL.n344 9.3005
R855 VTAIL.n326 VTAIL.n325 9.3005
R856 VTAIL.n339 VTAIL.n338 9.3005
R857 VTAIL.n337 VTAIL.n336 9.3005
R858 VTAIL.n330 VTAIL.n329 9.3005
R859 VTAIL.n742 VTAIL.n741 8.92171
R860 VTAIL.n757 VTAIL.n710 8.92171
R861 VTAIL.n788 VTAIL.n694 8.92171
R862 VTAIL.n50 VTAIL.n49 8.92171
R863 VTAIL.n65 VTAIL.n18 8.92171
R864 VTAIL.n96 VTAIL.n2 8.92171
R865 VTAIL.n148 VTAIL.n147 8.92171
R866 VTAIL.n163 VTAIL.n116 8.92171
R867 VTAIL.n194 VTAIL.n100 8.92171
R868 VTAIL.n248 VTAIL.n247 8.92171
R869 VTAIL.n263 VTAIL.n216 8.92171
R870 VTAIL.n294 VTAIL.n200 8.92171
R871 VTAIL.n690 VTAIL.n596 8.92171
R872 VTAIL.n661 VTAIL.n614 8.92171
R873 VTAIL.n646 VTAIL.n645 8.92171
R874 VTAIL.n590 VTAIL.n496 8.92171
R875 VTAIL.n561 VTAIL.n514 8.92171
R876 VTAIL.n546 VTAIL.n545 8.92171
R877 VTAIL.n492 VTAIL.n398 8.92171
R878 VTAIL.n463 VTAIL.n416 8.92171
R879 VTAIL.n448 VTAIL.n447 8.92171
R880 VTAIL.n392 VTAIL.n298 8.92171
R881 VTAIL.n363 VTAIL.n316 8.92171
R882 VTAIL.n348 VTAIL.n347 8.92171
R883 VTAIL.n745 VTAIL.n716 8.14595
R884 VTAIL.n754 VTAIL.n753 8.14595
R885 VTAIL.n53 VTAIL.n24 8.14595
R886 VTAIL.n62 VTAIL.n61 8.14595
R887 VTAIL.n151 VTAIL.n122 8.14595
R888 VTAIL.n160 VTAIL.n159 8.14595
R889 VTAIL.n251 VTAIL.n222 8.14595
R890 VTAIL.n260 VTAIL.n259 8.14595
R891 VTAIL.n658 VTAIL.n657 8.14595
R892 VTAIL.n649 VTAIL.n620 8.14595
R893 VTAIL.n558 VTAIL.n557 8.14595
R894 VTAIL.n549 VTAIL.n520 8.14595
R895 VTAIL.n460 VTAIL.n459 8.14595
R896 VTAIL.n451 VTAIL.n422 8.14595
R897 VTAIL.n360 VTAIL.n359 8.14595
R898 VTAIL.n351 VTAIL.n322 8.14595
R899 VTAIL.n746 VTAIL.n714 7.3702
R900 VTAIL.n750 VTAIL.n712 7.3702
R901 VTAIL.n54 VTAIL.n22 7.3702
R902 VTAIL.n58 VTAIL.n20 7.3702
R903 VTAIL.n152 VTAIL.n120 7.3702
R904 VTAIL.n156 VTAIL.n118 7.3702
R905 VTAIL.n252 VTAIL.n220 7.3702
R906 VTAIL.n256 VTAIL.n218 7.3702
R907 VTAIL.n654 VTAIL.n616 7.3702
R908 VTAIL.n650 VTAIL.n618 7.3702
R909 VTAIL.n554 VTAIL.n516 7.3702
R910 VTAIL.n550 VTAIL.n518 7.3702
R911 VTAIL.n456 VTAIL.n418 7.3702
R912 VTAIL.n452 VTAIL.n420 7.3702
R913 VTAIL.n356 VTAIL.n318 7.3702
R914 VTAIL.n352 VTAIL.n320 7.3702
R915 VTAIL.n749 VTAIL.n714 6.59444
R916 VTAIL.n750 VTAIL.n749 6.59444
R917 VTAIL.n57 VTAIL.n22 6.59444
R918 VTAIL.n58 VTAIL.n57 6.59444
R919 VTAIL.n155 VTAIL.n120 6.59444
R920 VTAIL.n156 VTAIL.n155 6.59444
R921 VTAIL.n255 VTAIL.n220 6.59444
R922 VTAIL.n256 VTAIL.n255 6.59444
R923 VTAIL.n654 VTAIL.n653 6.59444
R924 VTAIL.n653 VTAIL.n618 6.59444
R925 VTAIL.n554 VTAIL.n553 6.59444
R926 VTAIL.n553 VTAIL.n518 6.59444
R927 VTAIL.n456 VTAIL.n455 6.59444
R928 VTAIL.n455 VTAIL.n420 6.59444
R929 VTAIL.n356 VTAIL.n355 6.59444
R930 VTAIL.n355 VTAIL.n320 6.59444
R931 VTAIL.n746 VTAIL.n745 5.81868
R932 VTAIL.n753 VTAIL.n712 5.81868
R933 VTAIL.n54 VTAIL.n53 5.81868
R934 VTAIL.n61 VTAIL.n20 5.81868
R935 VTAIL.n152 VTAIL.n151 5.81868
R936 VTAIL.n159 VTAIL.n118 5.81868
R937 VTAIL.n252 VTAIL.n251 5.81868
R938 VTAIL.n259 VTAIL.n218 5.81868
R939 VTAIL.n657 VTAIL.n616 5.81868
R940 VTAIL.n650 VTAIL.n649 5.81868
R941 VTAIL.n557 VTAIL.n516 5.81868
R942 VTAIL.n550 VTAIL.n549 5.81868
R943 VTAIL.n459 VTAIL.n418 5.81868
R944 VTAIL.n452 VTAIL.n451 5.81868
R945 VTAIL.n359 VTAIL.n318 5.81868
R946 VTAIL.n352 VTAIL.n351 5.81868
R947 VTAIL.n742 VTAIL.n716 5.04292
R948 VTAIL.n754 VTAIL.n710 5.04292
R949 VTAIL.n790 VTAIL.n694 5.04292
R950 VTAIL.n50 VTAIL.n24 5.04292
R951 VTAIL.n62 VTAIL.n18 5.04292
R952 VTAIL.n98 VTAIL.n2 5.04292
R953 VTAIL.n148 VTAIL.n122 5.04292
R954 VTAIL.n160 VTAIL.n116 5.04292
R955 VTAIL.n196 VTAIL.n100 5.04292
R956 VTAIL.n248 VTAIL.n222 5.04292
R957 VTAIL.n260 VTAIL.n216 5.04292
R958 VTAIL.n296 VTAIL.n200 5.04292
R959 VTAIL.n692 VTAIL.n596 5.04292
R960 VTAIL.n658 VTAIL.n614 5.04292
R961 VTAIL.n646 VTAIL.n620 5.04292
R962 VTAIL.n592 VTAIL.n496 5.04292
R963 VTAIL.n558 VTAIL.n514 5.04292
R964 VTAIL.n546 VTAIL.n520 5.04292
R965 VTAIL.n494 VTAIL.n398 5.04292
R966 VTAIL.n460 VTAIL.n416 5.04292
R967 VTAIL.n448 VTAIL.n422 5.04292
R968 VTAIL.n394 VTAIL.n298 5.04292
R969 VTAIL.n360 VTAIL.n316 5.04292
R970 VTAIL.n348 VTAIL.n322 5.04292
R971 VTAIL.n741 VTAIL.n718 4.26717
R972 VTAIL.n758 VTAIL.n757 4.26717
R973 VTAIL.n788 VTAIL.n787 4.26717
R974 VTAIL.n49 VTAIL.n26 4.26717
R975 VTAIL.n66 VTAIL.n65 4.26717
R976 VTAIL.n96 VTAIL.n95 4.26717
R977 VTAIL.n147 VTAIL.n124 4.26717
R978 VTAIL.n164 VTAIL.n163 4.26717
R979 VTAIL.n194 VTAIL.n193 4.26717
R980 VTAIL.n247 VTAIL.n224 4.26717
R981 VTAIL.n264 VTAIL.n263 4.26717
R982 VTAIL.n294 VTAIL.n293 4.26717
R983 VTAIL.n690 VTAIL.n689 4.26717
R984 VTAIL.n662 VTAIL.n661 4.26717
R985 VTAIL.n645 VTAIL.n622 4.26717
R986 VTAIL.n590 VTAIL.n589 4.26717
R987 VTAIL.n562 VTAIL.n561 4.26717
R988 VTAIL.n545 VTAIL.n522 4.26717
R989 VTAIL.n492 VTAIL.n491 4.26717
R990 VTAIL.n464 VTAIL.n463 4.26717
R991 VTAIL.n447 VTAIL.n424 4.26717
R992 VTAIL.n392 VTAIL.n391 4.26717
R993 VTAIL.n364 VTAIL.n363 4.26717
R994 VTAIL.n347 VTAIL.n324 4.26717
R995 VTAIL.n725 VTAIL.n723 3.70982
R996 VTAIL.n33 VTAIL.n31 3.70982
R997 VTAIL.n131 VTAIL.n129 3.70982
R998 VTAIL.n231 VTAIL.n229 3.70982
R999 VTAIL.n629 VTAIL.n627 3.70982
R1000 VTAIL.n529 VTAIL.n527 3.70982
R1001 VTAIL.n431 VTAIL.n429 3.70982
R1002 VTAIL.n331 VTAIL.n329 3.70982
R1003 VTAIL.n738 VTAIL.n737 3.49141
R1004 VTAIL.n761 VTAIL.n708 3.49141
R1005 VTAIL.n784 VTAIL.n696 3.49141
R1006 VTAIL.n46 VTAIL.n45 3.49141
R1007 VTAIL.n69 VTAIL.n16 3.49141
R1008 VTAIL.n92 VTAIL.n4 3.49141
R1009 VTAIL.n144 VTAIL.n143 3.49141
R1010 VTAIL.n167 VTAIL.n114 3.49141
R1011 VTAIL.n190 VTAIL.n102 3.49141
R1012 VTAIL.n244 VTAIL.n243 3.49141
R1013 VTAIL.n267 VTAIL.n214 3.49141
R1014 VTAIL.n290 VTAIL.n202 3.49141
R1015 VTAIL.n686 VTAIL.n598 3.49141
R1016 VTAIL.n665 VTAIL.n612 3.49141
R1017 VTAIL.n642 VTAIL.n641 3.49141
R1018 VTAIL.n586 VTAIL.n498 3.49141
R1019 VTAIL.n565 VTAIL.n512 3.49141
R1020 VTAIL.n542 VTAIL.n541 3.49141
R1021 VTAIL.n488 VTAIL.n400 3.49141
R1022 VTAIL.n467 VTAIL.n414 3.49141
R1023 VTAIL.n444 VTAIL.n443 3.49141
R1024 VTAIL.n388 VTAIL.n300 3.49141
R1025 VTAIL.n367 VTAIL.n314 3.49141
R1026 VTAIL.n344 VTAIL.n343 3.49141
R1027 VTAIL.n734 VTAIL.n720 2.71565
R1028 VTAIL.n762 VTAIL.n706 2.71565
R1029 VTAIL.n783 VTAIL.n698 2.71565
R1030 VTAIL.n42 VTAIL.n28 2.71565
R1031 VTAIL.n70 VTAIL.n14 2.71565
R1032 VTAIL.n91 VTAIL.n6 2.71565
R1033 VTAIL.n140 VTAIL.n126 2.71565
R1034 VTAIL.n168 VTAIL.n112 2.71565
R1035 VTAIL.n189 VTAIL.n104 2.71565
R1036 VTAIL.n240 VTAIL.n226 2.71565
R1037 VTAIL.n268 VTAIL.n212 2.71565
R1038 VTAIL.n289 VTAIL.n204 2.71565
R1039 VTAIL.n685 VTAIL.n600 2.71565
R1040 VTAIL.n666 VTAIL.n610 2.71565
R1041 VTAIL.n638 VTAIL.n624 2.71565
R1042 VTAIL.n585 VTAIL.n500 2.71565
R1043 VTAIL.n566 VTAIL.n510 2.71565
R1044 VTAIL.n538 VTAIL.n524 2.71565
R1045 VTAIL.n487 VTAIL.n402 2.71565
R1046 VTAIL.n468 VTAIL.n412 2.71565
R1047 VTAIL.n440 VTAIL.n426 2.71565
R1048 VTAIL.n387 VTAIL.n302 2.71565
R1049 VTAIL.n368 VTAIL.n312 2.71565
R1050 VTAIL.n340 VTAIL.n326 2.71565
R1051 VTAIL.n397 VTAIL.n395 2.61257
R1052 VTAIL.n495 VTAIL.n397 2.61257
R1053 VTAIL.n595 VTAIL.n593 2.61257
R1054 VTAIL.n693 VTAIL.n595 2.61257
R1055 VTAIL.n297 VTAIL.n199 2.61257
R1056 VTAIL.n199 VTAIL.n197 2.61257
R1057 VTAIL.n99 VTAIL.n1 2.61257
R1058 VTAIL VTAIL.n791 2.55438
R1059 VTAIL.n733 VTAIL.n722 1.93989
R1060 VTAIL.n767 VTAIL.n765 1.93989
R1061 VTAIL.n780 VTAIL.n779 1.93989
R1062 VTAIL.n41 VTAIL.n30 1.93989
R1063 VTAIL.n75 VTAIL.n73 1.93989
R1064 VTAIL.n88 VTAIL.n87 1.93989
R1065 VTAIL.n139 VTAIL.n128 1.93989
R1066 VTAIL.n173 VTAIL.n171 1.93989
R1067 VTAIL.n186 VTAIL.n185 1.93989
R1068 VTAIL.n239 VTAIL.n228 1.93989
R1069 VTAIL.n273 VTAIL.n271 1.93989
R1070 VTAIL.n286 VTAIL.n285 1.93989
R1071 VTAIL.n682 VTAIL.n681 1.93989
R1072 VTAIL.n670 VTAIL.n669 1.93989
R1073 VTAIL.n637 VTAIL.n626 1.93989
R1074 VTAIL.n582 VTAIL.n581 1.93989
R1075 VTAIL.n570 VTAIL.n569 1.93989
R1076 VTAIL.n537 VTAIL.n526 1.93989
R1077 VTAIL.n484 VTAIL.n483 1.93989
R1078 VTAIL.n472 VTAIL.n471 1.93989
R1079 VTAIL.n439 VTAIL.n428 1.93989
R1080 VTAIL.n384 VTAIL.n383 1.93989
R1081 VTAIL.n372 VTAIL.n371 1.93989
R1082 VTAIL.n339 VTAIL.n328 1.93989
R1083 VTAIL.n0 VTAIL.t6 1.85158
R1084 VTAIL.n0 VTAIL.t3 1.85158
R1085 VTAIL.n198 VTAIL.t14 1.85158
R1086 VTAIL.n198 VTAIL.t9 1.85158
R1087 VTAIL.n594 VTAIL.t8 1.85158
R1088 VTAIL.n594 VTAIL.t11 1.85158
R1089 VTAIL.n396 VTAIL.t4 1.85158
R1090 VTAIL.n396 VTAIL.t7 1.85158
R1091 VTAIL.n730 VTAIL.n729 1.16414
R1092 VTAIL.n766 VTAIL.n704 1.16414
R1093 VTAIL.n776 VTAIL.n700 1.16414
R1094 VTAIL.n38 VTAIL.n37 1.16414
R1095 VTAIL.n74 VTAIL.n12 1.16414
R1096 VTAIL.n84 VTAIL.n8 1.16414
R1097 VTAIL.n136 VTAIL.n135 1.16414
R1098 VTAIL.n172 VTAIL.n110 1.16414
R1099 VTAIL.n182 VTAIL.n106 1.16414
R1100 VTAIL.n236 VTAIL.n235 1.16414
R1101 VTAIL.n272 VTAIL.n210 1.16414
R1102 VTAIL.n282 VTAIL.n206 1.16414
R1103 VTAIL.n678 VTAIL.n602 1.16414
R1104 VTAIL.n673 VTAIL.n607 1.16414
R1105 VTAIL.n634 VTAIL.n633 1.16414
R1106 VTAIL.n578 VTAIL.n502 1.16414
R1107 VTAIL.n573 VTAIL.n507 1.16414
R1108 VTAIL.n534 VTAIL.n533 1.16414
R1109 VTAIL.n480 VTAIL.n404 1.16414
R1110 VTAIL.n475 VTAIL.n409 1.16414
R1111 VTAIL.n436 VTAIL.n435 1.16414
R1112 VTAIL.n380 VTAIL.n304 1.16414
R1113 VTAIL.n375 VTAIL.n309 1.16414
R1114 VTAIL.n336 VTAIL.n335 1.16414
R1115 VTAIL.n593 VTAIL.n495 0.470328
R1116 VTAIL.n197 VTAIL.n99 0.470328
R1117 VTAIL.n726 VTAIL.n724 0.388379
R1118 VTAIL.n772 VTAIL.n771 0.388379
R1119 VTAIL.n775 VTAIL.n702 0.388379
R1120 VTAIL.n34 VTAIL.n32 0.388379
R1121 VTAIL.n80 VTAIL.n79 0.388379
R1122 VTAIL.n83 VTAIL.n10 0.388379
R1123 VTAIL.n132 VTAIL.n130 0.388379
R1124 VTAIL.n178 VTAIL.n177 0.388379
R1125 VTAIL.n181 VTAIL.n108 0.388379
R1126 VTAIL.n232 VTAIL.n230 0.388379
R1127 VTAIL.n278 VTAIL.n277 0.388379
R1128 VTAIL.n281 VTAIL.n208 0.388379
R1129 VTAIL.n677 VTAIL.n604 0.388379
R1130 VTAIL.n674 VTAIL.n606 0.388379
R1131 VTAIL.n630 VTAIL.n628 0.388379
R1132 VTAIL.n577 VTAIL.n504 0.388379
R1133 VTAIL.n574 VTAIL.n506 0.388379
R1134 VTAIL.n530 VTAIL.n528 0.388379
R1135 VTAIL.n479 VTAIL.n406 0.388379
R1136 VTAIL.n476 VTAIL.n408 0.388379
R1137 VTAIL.n432 VTAIL.n430 0.388379
R1138 VTAIL.n379 VTAIL.n306 0.388379
R1139 VTAIL.n376 VTAIL.n308 0.388379
R1140 VTAIL.n332 VTAIL.n330 0.388379
R1141 VTAIL.n731 VTAIL.n723 0.155672
R1142 VTAIL.n732 VTAIL.n731 0.155672
R1143 VTAIL.n732 VTAIL.n719 0.155672
R1144 VTAIL.n739 VTAIL.n719 0.155672
R1145 VTAIL.n740 VTAIL.n739 0.155672
R1146 VTAIL.n740 VTAIL.n715 0.155672
R1147 VTAIL.n747 VTAIL.n715 0.155672
R1148 VTAIL.n748 VTAIL.n747 0.155672
R1149 VTAIL.n748 VTAIL.n711 0.155672
R1150 VTAIL.n755 VTAIL.n711 0.155672
R1151 VTAIL.n756 VTAIL.n755 0.155672
R1152 VTAIL.n756 VTAIL.n707 0.155672
R1153 VTAIL.n763 VTAIL.n707 0.155672
R1154 VTAIL.n764 VTAIL.n763 0.155672
R1155 VTAIL.n764 VTAIL.n703 0.155672
R1156 VTAIL.n773 VTAIL.n703 0.155672
R1157 VTAIL.n774 VTAIL.n773 0.155672
R1158 VTAIL.n774 VTAIL.n699 0.155672
R1159 VTAIL.n781 VTAIL.n699 0.155672
R1160 VTAIL.n782 VTAIL.n781 0.155672
R1161 VTAIL.n782 VTAIL.n695 0.155672
R1162 VTAIL.n789 VTAIL.n695 0.155672
R1163 VTAIL.n39 VTAIL.n31 0.155672
R1164 VTAIL.n40 VTAIL.n39 0.155672
R1165 VTAIL.n40 VTAIL.n27 0.155672
R1166 VTAIL.n47 VTAIL.n27 0.155672
R1167 VTAIL.n48 VTAIL.n47 0.155672
R1168 VTAIL.n48 VTAIL.n23 0.155672
R1169 VTAIL.n55 VTAIL.n23 0.155672
R1170 VTAIL.n56 VTAIL.n55 0.155672
R1171 VTAIL.n56 VTAIL.n19 0.155672
R1172 VTAIL.n63 VTAIL.n19 0.155672
R1173 VTAIL.n64 VTAIL.n63 0.155672
R1174 VTAIL.n64 VTAIL.n15 0.155672
R1175 VTAIL.n71 VTAIL.n15 0.155672
R1176 VTAIL.n72 VTAIL.n71 0.155672
R1177 VTAIL.n72 VTAIL.n11 0.155672
R1178 VTAIL.n81 VTAIL.n11 0.155672
R1179 VTAIL.n82 VTAIL.n81 0.155672
R1180 VTAIL.n82 VTAIL.n7 0.155672
R1181 VTAIL.n89 VTAIL.n7 0.155672
R1182 VTAIL.n90 VTAIL.n89 0.155672
R1183 VTAIL.n90 VTAIL.n3 0.155672
R1184 VTAIL.n97 VTAIL.n3 0.155672
R1185 VTAIL.n137 VTAIL.n129 0.155672
R1186 VTAIL.n138 VTAIL.n137 0.155672
R1187 VTAIL.n138 VTAIL.n125 0.155672
R1188 VTAIL.n145 VTAIL.n125 0.155672
R1189 VTAIL.n146 VTAIL.n145 0.155672
R1190 VTAIL.n146 VTAIL.n121 0.155672
R1191 VTAIL.n153 VTAIL.n121 0.155672
R1192 VTAIL.n154 VTAIL.n153 0.155672
R1193 VTAIL.n154 VTAIL.n117 0.155672
R1194 VTAIL.n161 VTAIL.n117 0.155672
R1195 VTAIL.n162 VTAIL.n161 0.155672
R1196 VTAIL.n162 VTAIL.n113 0.155672
R1197 VTAIL.n169 VTAIL.n113 0.155672
R1198 VTAIL.n170 VTAIL.n169 0.155672
R1199 VTAIL.n170 VTAIL.n109 0.155672
R1200 VTAIL.n179 VTAIL.n109 0.155672
R1201 VTAIL.n180 VTAIL.n179 0.155672
R1202 VTAIL.n180 VTAIL.n105 0.155672
R1203 VTAIL.n187 VTAIL.n105 0.155672
R1204 VTAIL.n188 VTAIL.n187 0.155672
R1205 VTAIL.n188 VTAIL.n101 0.155672
R1206 VTAIL.n195 VTAIL.n101 0.155672
R1207 VTAIL.n237 VTAIL.n229 0.155672
R1208 VTAIL.n238 VTAIL.n237 0.155672
R1209 VTAIL.n238 VTAIL.n225 0.155672
R1210 VTAIL.n245 VTAIL.n225 0.155672
R1211 VTAIL.n246 VTAIL.n245 0.155672
R1212 VTAIL.n246 VTAIL.n221 0.155672
R1213 VTAIL.n253 VTAIL.n221 0.155672
R1214 VTAIL.n254 VTAIL.n253 0.155672
R1215 VTAIL.n254 VTAIL.n217 0.155672
R1216 VTAIL.n261 VTAIL.n217 0.155672
R1217 VTAIL.n262 VTAIL.n261 0.155672
R1218 VTAIL.n262 VTAIL.n213 0.155672
R1219 VTAIL.n269 VTAIL.n213 0.155672
R1220 VTAIL.n270 VTAIL.n269 0.155672
R1221 VTAIL.n270 VTAIL.n209 0.155672
R1222 VTAIL.n279 VTAIL.n209 0.155672
R1223 VTAIL.n280 VTAIL.n279 0.155672
R1224 VTAIL.n280 VTAIL.n205 0.155672
R1225 VTAIL.n287 VTAIL.n205 0.155672
R1226 VTAIL.n288 VTAIL.n287 0.155672
R1227 VTAIL.n288 VTAIL.n201 0.155672
R1228 VTAIL.n295 VTAIL.n201 0.155672
R1229 VTAIL.n691 VTAIL.n597 0.155672
R1230 VTAIL.n684 VTAIL.n597 0.155672
R1231 VTAIL.n684 VTAIL.n683 0.155672
R1232 VTAIL.n683 VTAIL.n601 0.155672
R1233 VTAIL.n676 VTAIL.n601 0.155672
R1234 VTAIL.n676 VTAIL.n675 0.155672
R1235 VTAIL.n675 VTAIL.n605 0.155672
R1236 VTAIL.n668 VTAIL.n605 0.155672
R1237 VTAIL.n668 VTAIL.n667 0.155672
R1238 VTAIL.n667 VTAIL.n611 0.155672
R1239 VTAIL.n660 VTAIL.n611 0.155672
R1240 VTAIL.n660 VTAIL.n659 0.155672
R1241 VTAIL.n659 VTAIL.n615 0.155672
R1242 VTAIL.n652 VTAIL.n615 0.155672
R1243 VTAIL.n652 VTAIL.n651 0.155672
R1244 VTAIL.n651 VTAIL.n619 0.155672
R1245 VTAIL.n644 VTAIL.n619 0.155672
R1246 VTAIL.n644 VTAIL.n643 0.155672
R1247 VTAIL.n643 VTAIL.n623 0.155672
R1248 VTAIL.n636 VTAIL.n623 0.155672
R1249 VTAIL.n636 VTAIL.n635 0.155672
R1250 VTAIL.n635 VTAIL.n627 0.155672
R1251 VTAIL.n591 VTAIL.n497 0.155672
R1252 VTAIL.n584 VTAIL.n497 0.155672
R1253 VTAIL.n584 VTAIL.n583 0.155672
R1254 VTAIL.n583 VTAIL.n501 0.155672
R1255 VTAIL.n576 VTAIL.n501 0.155672
R1256 VTAIL.n576 VTAIL.n575 0.155672
R1257 VTAIL.n575 VTAIL.n505 0.155672
R1258 VTAIL.n568 VTAIL.n505 0.155672
R1259 VTAIL.n568 VTAIL.n567 0.155672
R1260 VTAIL.n567 VTAIL.n511 0.155672
R1261 VTAIL.n560 VTAIL.n511 0.155672
R1262 VTAIL.n560 VTAIL.n559 0.155672
R1263 VTAIL.n559 VTAIL.n515 0.155672
R1264 VTAIL.n552 VTAIL.n515 0.155672
R1265 VTAIL.n552 VTAIL.n551 0.155672
R1266 VTAIL.n551 VTAIL.n519 0.155672
R1267 VTAIL.n544 VTAIL.n519 0.155672
R1268 VTAIL.n544 VTAIL.n543 0.155672
R1269 VTAIL.n543 VTAIL.n523 0.155672
R1270 VTAIL.n536 VTAIL.n523 0.155672
R1271 VTAIL.n536 VTAIL.n535 0.155672
R1272 VTAIL.n535 VTAIL.n527 0.155672
R1273 VTAIL.n493 VTAIL.n399 0.155672
R1274 VTAIL.n486 VTAIL.n399 0.155672
R1275 VTAIL.n486 VTAIL.n485 0.155672
R1276 VTAIL.n485 VTAIL.n403 0.155672
R1277 VTAIL.n478 VTAIL.n403 0.155672
R1278 VTAIL.n478 VTAIL.n477 0.155672
R1279 VTAIL.n477 VTAIL.n407 0.155672
R1280 VTAIL.n470 VTAIL.n407 0.155672
R1281 VTAIL.n470 VTAIL.n469 0.155672
R1282 VTAIL.n469 VTAIL.n413 0.155672
R1283 VTAIL.n462 VTAIL.n413 0.155672
R1284 VTAIL.n462 VTAIL.n461 0.155672
R1285 VTAIL.n461 VTAIL.n417 0.155672
R1286 VTAIL.n454 VTAIL.n417 0.155672
R1287 VTAIL.n454 VTAIL.n453 0.155672
R1288 VTAIL.n453 VTAIL.n421 0.155672
R1289 VTAIL.n446 VTAIL.n421 0.155672
R1290 VTAIL.n446 VTAIL.n445 0.155672
R1291 VTAIL.n445 VTAIL.n425 0.155672
R1292 VTAIL.n438 VTAIL.n425 0.155672
R1293 VTAIL.n438 VTAIL.n437 0.155672
R1294 VTAIL.n437 VTAIL.n429 0.155672
R1295 VTAIL.n393 VTAIL.n299 0.155672
R1296 VTAIL.n386 VTAIL.n299 0.155672
R1297 VTAIL.n386 VTAIL.n385 0.155672
R1298 VTAIL.n385 VTAIL.n303 0.155672
R1299 VTAIL.n378 VTAIL.n303 0.155672
R1300 VTAIL.n378 VTAIL.n377 0.155672
R1301 VTAIL.n377 VTAIL.n307 0.155672
R1302 VTAIL.n370 VTAIL.n307 0.155672
R1303 VTAIL.n370 VTAIL.n369 0.155672
R1304 VTAIL.n369 VTAIL.n313 0.155672
R1305 VTAIL.n362 VTAIL.n313 0.155672
R1306 VTAIL.n362 VTAIL.n361 0.155672
R1307 VTAIL.n361 VTAIL.n317 0.155672
R1308 VTAIL.n354 VTAIL.n317 0.155672
R1309 VTAIL.n354 VTAIL.n353 0.155672
R1310 VTAIL.n353 VTAIL.n321 0.155672
R1311 VTAIL.n346 VTAIL.n321 0.155672
R1312 VTAIL.n346 VTAIL.n345 0.155672
R1313 VTAIL.n345 VTAIL.n325 0.155672
R1314 VTAIL.n338 VTAIL.n325 0.155672
R1315 VTAIL.n338 VTAIL.n337 0.155672
R1316 VTAIL.n337 VTAIL.n329 0.155672
R1317 VTAIL VTAIL.n1 0.0586897
R1318 VDD1 VDD1.n0 71.1622
R1319 VDD1.n3 VDD1.n2 71.0485
R1320 VDD1.n3 VDD1.n1 71.0485
R1321 VDD1.n5 VDD1.n4 69.7978
R1322 VDD1.n5 VDD1.n3 51.1906
R1323 VDD1.n4 VDD1.t5 1.85158
R1324 VDD1.n4 VDD1.t4 1.85158
R1325 VDD1.n0 VDD1.t0 1.85158
R1326 VDD1.n0 VDD1.t7 1.85158
R1327 VDD1.n2 VDD1.t6 1.85158
R1328 VDD1.n2 VDD1.t2 1.85158
R1329 VDD1.n1 VDD1.t1 1.85158
R1330 VDD1.n1 VDD1.t3 1.85158
R1331 VDD1 VDD1.n5 1.24834
R1332 B.n505 B.n504 585
R1333 B.n503 B.n148 585
R1334 B.n502 B.n501 585
R1335 B.n500 B.n149 585
R1336 B.n499 B.n498 585
R1337 B.n497 B.n150 585
R1338 B.n496 B.n495 585
R1339 B.n494 B.n151 585
R1340 B.n493 B.n492 585
R1341 B.n491 B.n152 585
R1342 B.n490 B.n489 585
R1343 B.n488 B.n153 585
R1344 B.n487 B.n486 585
R1345 B.n485 B.n154 585
R1346 B.n484 B.n483 585
R1347 B.n482 B.n155 585
R1348 B.n481 B.n480 585
R1349 B.n479 B.n156 585
R1350 B.n478 B.n477 585
R1351 B.n476 B.n157 585
R1352 B.n475 B.n474 585
R1353 B.n473 B.n158 585
R1354 B.n472 B.n471 585
R1355 B.n470 B.n159 585
R1356 B.n469 B.n468 585
R1357 B.n467 B.n160 585
R1358 B.n466 B.n465 585
R1359 B.n464 B.n161 585
R1360 B.n463 B.n462 585
R1361 B.n461 B.n162 585
R1362 B.n460 B.n459 585
R1363 B.n458 B.n163 585
R1364 B.n457 B.n456 585
R1365 B.n455 B.n164 585
R1366 B.n454 B.n453 585
R1367 B.n452 B.n165 585
R1368 B.n451 B.n450 585
R1369 B.n449 B.n166 585
R1370 B.n448 B.n447 585
R1371 B.n446 B.n167 585
R1372 B.n445 B.n444 585
R1373 B.n443 B.n168 585
R1374 B.n442 B.n441 585
R1375 B.n440 B.n169 585
R1376 B.n439 B.n438 585
R1377 B.n437 B.n170 585
R1378 B.n436 B.n435 585
R1379 B.n434 B.n171 585
R1380 B.n433 B.n432 585
R1381 B.n431 B.n172 585
R1382 B.n430 B.n429 585
R1383 B.n428 B.n173 585
R1384 B.n427 B.n426 585
R1385 B.n425 B.n174 585
R1386 B.n424 B.n423 585
R1387 B.n422 B.n175 585
R1388 B.n421 B.n420 585
R1389 B.n419 B.n176 585
R1390 B.n418 B.n417 585
R1391 B.n413 B.n177 585
R1392 B.n412 B.n411 585
R1393 B.n410 B.n178 585
R1394 B.n409 B.n408 585
R1395 B.n407 B.n179 585
R1396 B.n406 B.n405 585
R1397 B.n404 B.n180 585
R1398 B.n403 B.n402 585
R1399 B.n400 B.n181 585
R1400 B.n399 B.n398 585
R1401 B.n397 B.n184 585
R1402 B.n396 B.n395 585
R1403 B.n394 B.n185 585
R1404 B.n393 B.n392 585
R1405 B.n391 B.n186 585
R1406 B.n390 B.n389 585
R1407 B.n388 B.n187 585
R1408 B.n387 B.n386 585
R1409 B.n385 B.n188 585
R1410 B.n384 B.n383 585
R1411 B.n382 B.n189 585
R1412 B.n381 B.n380 585
R1413 B.n379 B.n190 585
R1414 B.n378 B.n377 585
R1415 B.n376 B.n191 585
R1416 B.n375 B.n374 585
R1417 B.n373 B.n192 585
R1418 B.n372 B.n371 585
R1419 B.n370 B.n193 585
R1420 B.n369 B.n368 585
R1421 B.n367 B.n194 585
R1422 B.n366 B.n365 585
R1423 B.n364 B.n195 585
R1424 B.n363 B.n362 585
R1425 B.n361 B.n196 585
R1426 B.n360 B.n359 585
R1427 B.n358 B.n197 585
R1428 B.n357 B.n356 585
R1429 B.n355 B.n198 585
R1430 B.n354 B.n353 585
R1431 B.n352 B.n199 585
R1432 B.n351 B.n350 585
R1433 B.n349 B.n200 585
R1434 B.n348 B.n347 585
R1435 B.n346 B.n201 585
R1436 B.n345 B.n344 585
R1437 B.n343 B.n202 585
R1438 B.n342 B.n341 585
R1439 B.n340 B.n203 585
R1440 B.n339 B.n338 585
R1441 B.n337 B.n204 585
R1442 B.n336 B.n335 585
R1443 B.n334 B.n205 585
R1444 B.n333 B.n332 585
R1445 B.n331 B.n206 585
R1446 B.n330 B.n329 585
R1447 B.n328 B.n207 585
R1448 B.n327 B.n326 585
R1449 B.n325 B.n208 585
R1450 B.n324 B.n323 585
R1451 B.n322 B.n209 585
R1452 B.n321 B.n320 585
R1453 B.n319 B.n210 585
R1454 B.n318 B.n317 585
R1455 B.n316 B.n211 585
R1456 B.n315 B.n314 585
R1457 B.n506 B.n147 585
R1458 B.n508 B.n507 585
R1459 B.n509 B.n146 585
R1460 B.n511 B.n510 585
R1461 B.n512 B.n145 585
R1462 B.n514 B.n513 585
R1463 B.n515 B.n144 585
R1464 B.n517 B.n516 585
R1465 B.n518 B.n143 585
R1466 B.n520 B.n519 585
R1467 B.n521 B.n142 585
R1468 B.n523 B.n522 585
R1469 B.n524 B.n141 585
R1470 B.n526 B.n525 585
R1471 B.n527 B.n140 585
R1472 B.n529 B.n528 585
R1473 B.n530 B.n139 585
R1474 B.n532 B.n531 585
R1475 B.n533 B.n138 585
R1476 B.n535 B.n534 585
R1477 B.n536 B.n137 585
R1478 B.n538 B.n537 585
R1479 B.n539 B.n136 585
R1480 B.n541 B.n540 585
R1481 B.n542 B.n135 585
R1482 B.n544 B.n543 585
R1483 B.n545 B.n134 585
R1484 B.n547 B.n546 585
R1485 B.n548 B.n133 585
R1486 B.n550 B.n549 585
R1487 B.n551 B.n132 585
R1488 B.n553 B.n552 585
R1489 B.n554 B.n131 585
R1490 B.n556 B.n555 585
R1491 B.n557 B.n130 585
R1492 B.n559 B.n558 585
R1493 B.n560 B.n129 585
R1494 B.n562 B.n561 585
R1495 B.n563 B.n128 585
R1496 B.n565 B.n564 585
R1497 B.n566 B.n127 585
R1498 B.n568 B.n567 585
R1499 B.n569 B.n126 585
R1500 B.n571 B.n570 585
R1501 B.n572 B.n125 585
R1502 B.n574 B.n573 585
R1503 B.n575 B.n124 585
R1504 B.n577 B.n576 585
R1505 B.n578 B.n123 585
R1506 B.n580 B.n579 585
R1507 B.n581 B.n122 585
R1508 B.n583 B.n582 585
R1509 B.n584 B.n121 585
R1510 B.n586 B.n585 585
R1511 B.n587 B.n120 585
R1512 B.n589 B.n588 585
R1513 B.n590 B.n119 585
R1514 B.n592 B.n591 585
R1515 B.n593 B.n118 585
R1516 B.n595 B.n594 585
R1517 B.n596 B.n117 585
R1518 B.n598 B.n597 585
R1519 B.n599 B.n116 585
R1520 B.n601 B.n600 585
R1521 B.n602 B.n115 585
R1522 B.n604 B.n603 585
R1523 B.n605 B.n114 585
R1524 B.n607 B.n606 585
R1525 B.n608 B.n113 585
R1526 B.n610 B.n609 585
R1527 B.n611 B.n112 585
R1528 B.n613 B.n612 585
R1529 B.n614 B.n111 585
R1530 B.n616 B.n615 585
R1531 B.n617 B.n110 585
R1532 B.n619 B.n618 585
R1533 B.n620 B.n109 585
R1534 B.n622 B.n621 585
R1535 B.n623 B.n108 585
R1536 B.n625 B.n624 585
R1537 B.n626 B.n107 585
R1538 B.n628 B.n627 585
R1539 B.n629 B.n106 585
R1540 B.n631 B.n630 585
R1541 B.n632 B.n105 585
R1542 B.n634 B.n633 585
R1543 B.n635 B.n104 585
R1544 B.n637 B.n636 585
R1545 B.n638 B.n103 585
R1546 B.n640 B.n639 585
R1547 B.n641 B.n102 585
R1548 B.n643 B.n642 585
R1549 B.n644 B.n101 585
R1550 B.n646 B.n645 585
R1551 B.n647 B.n100 585
R1552 B.n649 B.n648 585
R1553 B.n650 B.n99 585
R1554 B.n652 B.n651 585
R1555 B.n653 B.n98 585
R1556 B.n655 B.n654 585
R1557 B.n656 B.n97 585
R1558 B.n658 B.n657 585
R1559 B.n659 B.n96 585
R1560 B.n661 B.n660 585
R1561 B.n662 B.n95 585
R1562 B.n664 B.n663 585
R1563 B.n853 B.n28 585
R1564 B.n852 B.n851 585
R1565 B.n850 B.n29 585
R1566 B.n849 B.n848 585
R1567 B.n847 B.n30 585
R1568 B.n846 B.n845 585
R1569 B.n844 B.n31 585
R1570 B.n843 B.n842 585
R1571 B.n841 B.n32 585
R1572 B.n840 B.n839 585
R1573 B.n838 B.n33 585
R1574 B.n837 B.n836 585
R1575 B.n835 B.n34 585
R1576 B.n834 B.n833 585
R1577 B.n832 B.n35 585
R1578 B.n831 B.n830 585
R1579 B.n829 B.n36 585
R1580 B.n828 B.n827 585
R1581 B.n826 B.n37 585
R1582 B.n825 B.n824 585
R1583 B.n823 B.n38 585
R1584 B.n822 B.n821 585
R1585 B.n820 B.n39 585
R1586 B.n819 B.n818 585
R1587 B.n817 B.n40 585
R1588 B.n816 B.n815 585
R1589 B.n814 B.n41 585
R1590 B.n813 B.n812 585
R1591 B.n811 B.n42 585
R1592 B.n810 B.n809 585
R1593 B.n808 B.n43 585
R1594 B.n807 B.n806 585
R1595 B.n805 B.n44 585
R1596 B.n804 B.n803 585
R1597 B.n802 B.n45 585
R1598 B.n801 B.n800 585
R1599 B.n799 B.n46 585
R1600 B.n798 B.n797 585
R1601 B.n796 B.n47 585
R1602 B.n795 B.n794 585
R1603 B.n793 B.n48 585
R1604 B.n792 B.n791 585
R1605 B.n790 B.n49 585
R1606 B.n789 B.n788 585
R1607 B.n787 B.n50 585
R1608 B.n786 B.n785 585
R1609 B.n784 B.n51 585
R1610 B.n783 B.n782 585
R1611 B.n781 B.n52 585
R1612 B.n780 B.n779 585
R1613 B.n778 B.n53 585
R1614 B.n777 B.n776 585
R1615 B.n775 B.n54 585
R1616 B.n774 B.n773 585
R1617 B.n772 B.n55 585
R1618 B.n771 B.n770 585
R1619 B.n769 B.n56 585
R1620 B.n768 B.n767 585
R1621 B.n765 B.n57 585
R1622 B.n764 B.n763 585
R1623 B.n762 B.n60 585
R1624 B.n761 B.n760 585
R1625 B.n759 B.n61 585
R1626 B.n758 B.n757 585
R1627 B.n756 B.n62 585
R1628 B.n755 B.n754 585
R1629 B.n753 B.n63 585
R1630 B.n751 B.n750 585
R1631 B.n749 B.n66 585
R1632 B.n748 B.n747 585
R1633 B.n746 B.n67 585
R1634 B.n745 B.n744 585
R1635 B.n743 B.n68 585
R1636 B.n742 B.n741 585
R1637 B.n740 B.n69 585
R1638 B.n739 B.n738 585
R1639 B.n737 B.n70 585
R1640 B.n736 B.n735 585
R1641 B.n734 B.n71 585
R1642 B.n733 B.n732 585
R1643 B.n731 B.n72 585
R1644 B.n730 B.n729 585
R1645 B.n728 B.n73 585
R1646 B.n727 B.n726 585
R1647 B.n725 B.n74 585
R1648 B.n724 B.n723 585
R1649 B.n722 B.n75 585
R1650 B.n721 B.n720 585
R1651 B.n719 B.n76 585
R1652 B.n718 B.n717 585
R1653 B.n716 B.n77 585
R1654 B.n715 B.n714 585
R1655 B.n713 B.n78 585
R1656 B.n712 B.n711 585
R1657 B.n710 B.n79 585
R1658 B.n709 B.n708 585
R1659 B.n707 B.n80 585
R1660 B.n706 B.n705 585
R1661 B.n704 B.n81 585
R1662 B.n703 B.n702 585
R1663 B.n701 B.n82 585
R1664 B.n700 B.n699 585
R1665 B.n698 B.n83 585
R1666 B.n697 B.n696 585
R1667 B.n695 B.n84 585
R1668 B.n694 B.n693 585
R1669 B.n692 B.n85 585
R1670 B.n691 B.n690 585
R1671 B.n689 B.n86 585
R1672 B.n688 B.n687 585
R1673 B.n686 B.n87 585
R1674 B.n685 B.n684 585
R1675 B.n683 B.n88 585
R1676 B.n682 B.n681 585
R1677 B.n680 B.n89 585
R1678 B.n679 B.n678 585
R1679 B.n677 B.n90 585
R1680 B.n676 B.n675 585
R1681 B.n674 B.n91 585
R1682 B.n673 B.n672 585
R1683 B.n671 B.n92 585
R1684 B.n670 B.n669 585
R1685 B.n668 B.n93 585
R1686 B.n667 B.n666 585
R1687 B.n665 B.n94 585
R1688 B.n855 B.n854 585
R1689 B.n856 B.n27 585
R1690 B.n858 B.n857 585
R1691 B.n859 B.n26 585
R1692 B.n861 B.n860 585
R1693 B.n862 B.n25 585
R1694 B.n864 B.n863 585
R1695 B.n865 B.n24 585
R1696 B.n867 B.n866 585
R1697 B.n868 B.n23 585
R1698 B.n870 B.n869 585
R1699 B.n871 B.n22 585
R1700 B.n873 B.n872 585
R1701 B.n874 B.n21 585
R1702 B.n876 B.n875 585
R1703 B.n877 B.n20 585
R1704 B.n879 B.n878 585
R1705 B.n880 B.n19 585
R1706 B.n882 B.n881 585
R1707 B.n883 B.n18 585
R1708 B.n885 B.n884 585
R1709 B.n886 B.n17 585
R1710 B.n888 B.n887 585
R1711 B.n889 B.n16 585
R1712 B.n891 B.n890 585
R1713 B.n892 B.n15 585
R1714 B.n894 B.n893 585
R1715 B.n895 B.n14 585
R1716 B.n897 B.n896 585
R1717 B.n898 B.n13 585
R1718 B.n900 B.n899 585
R1719 B.n901 B.n12 585
R1720 B.n903 B.n902 585
R1721 B.n904 B.n11 585
R1722 B.n906 B.n905 585
R1723 B.n907 B.n10 585
R1724 B.n909 B.n908 585
R1725 B.n910 B.n9 585
R1726 B.n912 B.n911 585
R1727 B.n913 B.n8 585
R1728 B.n915 B.n914 585
R1729 B.n916 B.n7 585
R1730 B.n918 B.n917 585
R1731 B.n919 B.n6 585
R1732 B.n921 B.n920 585
R1733 B.n922 B.n5 585
R1734 B.n924 B.n923 585
R1735 B.n925 B.n4 585
R1736 B.n927 B.n926 585
R1737 B.n928 B.n3 585
R1738 B.n930 B.n929 585
R1739 B.n931 B.n0 585
R1740 B.n2 B.n1 585
R1741 B.n238 B.n237 585
R1742 B.n240 B.n239 585
R1743 B.n241 B.n236 585
R1744 B.n243 B.n242 585
R1745 B.n244 B.n235 585
R1746 B.n246 B.n245 585
R1747 B.n247 B.n234 585
R1748 B.n249 B.n248 585
R1749 B.n250 B.n233 585
R1750 B.n252 B.n251 585
R1751 B.n253 B.n232 585
R1752 B.n255 B.n254 585
R1753 B.n256 B.n231 585
R1754 B.n258 B.n257 585
R1755 B.n259 B.n230 585
R1756 B.n261 B.n260 585
R1757 B.n262 B.n229 585
R1758 B.n264 B.n263 585
R1759 B.n265 B.n228 585
R1760 B.n267 B.n266 585
R1761 B.n268 B.n227 585
R1762 B.n270 B.n269 585
R1763 B.n271 B.n226 585
R1764 B.n273 B.n272 585
R1765 B.n274 B.n225 585
R1766 B.n276 B.n275 585
R1767 B.n277 B.n224 585
R1768 B.n279 B.n278 585
R1769 B.n280 B.n223 585
R1770 B.n282 B.n281 585
R1771 B.n283 B.n222 585
R1772 B.n285 B.n284 585
R1773 B.n286 B.n221 585
R1774 B.n288 B.n287 585
R1775 B.n289 B.n220 585
R1776 B.n291 B.n290 585
R1777 B.n292 B.n219 585
R1778 B.n294 B.n293 585
R1779 B.n295 B.n218 585
R1780 B.n297 B.n296 585
R1781 B.n298 B.n217 585
R1782 B.n300 B.n299 585
R1783 B.n301 B.n216 585
R1784 B.n303 B.n302 585
R1785 B.n304 B.n215 585
R1786 B.n306 B.n305 585
R1787 B.n307 B.n214 585
R1788 B.n309 B.n308 585
R1789 B.n310 B.n213 585
R1790 B.n312 B.n311 585
R1791 B.n313 B.n212 585
R1792 B.n314 B.n313 569.379
R1793 B.n504 B.n147 569.379
R1794 B.n665 B.n664 569.379
R1795 B.n854 B.n853 569.379
R1796 B.n414 B.t4 534.605
R1797 B.n64 B.t8 534.605
R1798 B.n182 B.t10 534.605
R1799 B.n58 B.t2 534.605
R1800 B.n415 B.t5 475.841
R1801 B.n65 B.t7 475.841
R1802 B.n183 B.t11 475.841
R1803 B.n59 B.t1 475.841
R1804 B.n182 B.t9 364.933
R1805 B.n414 B.t3 364.933
R1806 B.n64 B.t6 364.933
R1807 B.n58 B.t0 364.933
R1808 B.n933 B.n932 256.663
R1809 B.n932 B.n931 235.042
R1810 B.n932 B.n2 235.042
R1811 B.n314 B.n211 163.367
R1812 B.n318 B.n211 163.367
R1813 B.n319 B.n318 163.367
R1814 B.n320 B.n319 163.367
R1815 B.n320 B.n209 163.367
R1816 B.n324 B.n209 163.367
R1817 B.n325 B.n324 163.367
R1818 B.n326 B.n325 163.367
R1819 B.n326 B.n207 163.367
R1820 B.n330 B.n207 163.367
R1821 B.n331 B.n330 163.367
R1822 B.n332 B.n331 163.367
R1823 B.n332 B.n205 163.367
R1824 B.n336 B.n205 163.367
R1825 B.n337 B.n336 163.367
R1826 B.n338 B.n337 163.367
R1827 B.n338 B.n203 163.367
R1828 B.n342 B.n203 163.367
R1829 B.n343 B.n342 163.367
R1830 B.n344 B.n343 163.367
R1831 B.n344 B.n201 163.367
R1832 B.n348 B.n201 163.367
R1833 B.n349 B.n348 163.367
R1834 B.n350 B.n349 163.367
R1835 B.n350 B.n199 163.367
R1836 B.n354 B.n199 163.367
R1837 B.n355 B.n354 163.367
R1838 B.n356 B.n355 163.367
R1839 B.n356 B.n197 163.367
R1840 B.n360 B.n197 163.367
R1841 B.n361 B.n360 163.367
R1842 B.n362 B.n361 163.367
R1843 B.n362 B.n195 163.367
R1844 B.n366 B.n195 163.367
R1845 B.n367 B.n366 163.367
R1846 B.n368 B.n367 163.367
R1847 B.n368 B.n193 163.367
R1848 B.n372 B.n193 163.367
R1849 B.n373 B.n372 163.367
R1850 B.n374 B.n373 163.367
R1851 B.n374 B.n191 163.367
R1852 B.n378 B.n191 163.367
R1853 B.n379 B.n378 163.367
R1854 B.n380 B.n379 163.367
R1855 B.n380 B.n189 163.367
R1856 B.n384 B.n189 163.367
R1857 B.n385 B.n384 163.367
R1858 B.n386 B.n385 163.367
R1859 B.n386 B.n187 163.367
R1860 B.n390 B.n187 163.367
R1861 B.n391 B.n390 163.367
R1862 B.n392 B.n391 163.367
R1863 B.n392 B.n185 163.367
R1864 B.n396 B.n185 163.367
R1865 B.n397 B.n396 163.367
R1866 B.n398 B.n397 163.367
R1867 B.n398 B.n181 163.367
R1868 B.n403 B.n181 163.367
R1869 B.n404 B.n403 163.367
R1870 B.n405 B.n404 163.367
R1871 B.n405 B.n179 163.367
R1872 B.n409 B.n179 163.367
R1873 B.n410 B.n409 163.367
R1874 B.n411 B.n410 163.367
R1875 B.n411 B.n177 163.367
R1876 B.n418 B.n177 163.367
R1877 B.n419 B.n418 163.367
R1878 B.n420 B.n419 163.367
R1879 B.n420 B.n175 163.367
R1880 B.n424 B.n175 163.367
R1881 B.n425 B.n424 163.367
R1882 B.n426 B.n425 163.367
R1883 B.n426 B.n173 163.367
R1884 B.n430 B.n173 163.367
R1885 B.n431 B.n430 163.367
R1886 B.n432 B.n431 163.367
R1887 B.n432 B.n171 163.367
R1888 B.n436 B.n171 163.367
R1889 B.n437 B.n436 163.367
R1890 B.n438 B.n437 163.367
R1891 B.n438 B.n169 163.367
R1892 B.n442 B.n169 163.367
R1893 B.n443 B.n442 163.367
R1894 B.n444 B.n443 163.367
R1895 B.n444 B.n167 163.367
R1896 B.n448 B.n167 163.367
R1897 B.n449 B.n448 163.367
R1898 B.n450 B.n449 163.367
R1899 B.n450 B.n165 163.367
R1900 B.n454 B.n165 163.367
R1901 B.n455 B.n454 163.367
R1902 B.n456 B.n455 163.367
R1903 B.n456 B.n163 163.367
R1904 B.n460 B.n163 163.367
R1905 B.n461 B.n460 163.367
R1906 B.n462 B.n461 163.367
R1907 B.n462 B.n161 163.367
R1908 B.n466 B.n161 163.367
R1909 B.n467 B.n466 163.367
R1910 B.n468 B.n467 163.367
R1911 B.n468 B.n159 163.367
R1912 B.n472 B.n159 163.367
R1913 B.n473 B.n472 163.367
R1914 B.n474 B.n473 163.367
R1915 B.n474 B.n157 163.367
R1916 B.n478 B.n157 163.367
R1917 B.n479 B.n478 163.367
R1918 B.n480 B.n479 163.367
R1919 B.n480 B.n155 163.367
R1920 B.n484 B.n155 163.367
R1921 B.n485 B.n484 163.367
R1922 B.n486 B.n485 163.367
R1923 B.n486 B.n153 163.367
R1924 B.n490 B.n153 163.367
R1925 B.n491 B.n490 163.367
R1926 B.n492 B.n491 163.367
R1927 B.n492 B.n151 163.367
R1928 B.n496 B.n151 163.367
R1929 B.n497 B.n496 163.367
R1930 B.n498 B.n497 163.367
R1931 B.n498 B.n149 163.367
R1932 B.n502 B.n149 163.367
R1933 B.n503 B.n502 163.367
R1934 B.n504 B.n503 163.367
R1935 B.n664 B.n95 163.367
R1936 B.n660 B.n95 163.367
R1937 B.n660 B.n659 163.367
R1938 B.n659 B.n658 163.367
R1939 B.n658 B.n97 163.367
R1940 B.n654 B.n97 163.367
R1941 B.n654 B.n653 163.367
R1942 B.n653 B.n652 163.367
R1943 B.n652 B.n99 163.367
R1944 B.n648 B.n99 163.367
R1945 B.n648 B.n647 163.367
R1946 B.n647 B.n646 163.367
R1947 B.n646 B.n101 163.367
R1948 B.n642 B.n101 163.367
R1949 B.n642 B.n641 163.367
R1950 B.n641 B.n640 163.367
R1951 B.n640 B.n103 163.367
R1952 B.n636 B.n103 163.367
R1953 B.n636 B.n635 163.367
R1954 B.n635 B.n634 163.367
R1955 B.n634 B.n105 163.367
R1956 B.n630 B.n105 163.367
R1957 B.n630 B.n629 163.367
R1958 B.n629 B.n628 163.367
R1959 B.n628 B.n107 163.367
R1960 B.n624 B.n107 163.367
R1961 B.n624 B.n623 163.367
R1962 B.n623 B.n622 163.367
R1963 B.n622 B.n109 163.367
R1964 B.n618 B.n109 163.367
R1965 B.n618 B.n617 163.367
R1966 B.n617 B.n616 163.367
R1967 B.n616 B.n111 163.367
R1968 B.n612 B.n111 163.367
R1969 B.n612 B.n611 163.367
R1970 B.n611 B.n610 163.367
R1971 B.n610 B.n113 163.367
R1972 B.n606 B.n113 163.367
R1973 B.n606 B.n605 163.367
R1974 B.n605 B.n604 163.367
R1975 B.n604 B.n115 163.367
R1976 B.n600 B.n115 163.367
R1977 B.n600 B.n599 163.367
R1978 B.n599 B.n598 163.367
R1979 B.n598 B.n117 163.367
R1980 B.n594 B.n117 163.367
R1981 B.n594 B.n593 163.367
R1982 B.n593 B.n592 163.367
R1983 B.n592 B.n119 163.367
R1984 B.n588 B.n119 163.367
R1985 B.n588 B.n587 163.367
R1986 B.n587 B.n586 163.367
R1987 B.n586 B.n121 163.367
R1988 B.n582 B.n121 163.367
R1989 B.n582 B.n581 163.367
R1990 B.n581 B.n580 163.367
R1991 B.n580 B.n123 163.367
R1992 B.n576 B.n123 163.367
R1993 B.n576 B.n575 163.367
R1994 B.n575 B.n574 163.367
R1995 B.n574 B.n125 163.367
R1996 B.n570 B.n125 163.367
R1997 B.n570 B.n569 163.367
R1998 B.n569 B.n568 163.367
R1999 B.n568 B.n127 163.367
R2000 B.n564 B.n127 163.367
R2001 B.n564 B.n563 163.367
R2002 B.n563 B.n562 163.367
R2003 B.n562 B.n129 163.367
R2004 B.n558 B.n129 163.367
R2005 B.n558 B.n557 163.367
R2006 B.n557 B.n556 163.367
R2007 B.n556 B.n131 163.367
R2008 B.n552 B.n131 163.367
R2009 B.n552 B.n551 163.367
R2010 B.n551 B.n550 163.367
R2011 B.n550 B.n133 163.367
R2012 B.n546 B.n133 163.367
R2013 B.n546 B.n545 163.367
R2014 B.n545 B.n544 163.367
R2015 B.n544 B.n135 163.367
R2016 B.n540 B.n135 163.367
R2017 B.n540 B.n539 163.367
R2018 B.n539 B.n538 163.367
R2019 B.n538 B.n137 163.367
R2020 B.n534 B.n137 163.367
R2021 B.n534 B.n533 163.367
R2022 B.n533 B.n532 163.367
R2023 B.n532 B.n139 163.367
R2024 B.n528 B.n139 163.367
R2025 B.n528 B.n527 163.367
R2026 B.n527 B.n526 163.367
R2027 B.n526 B.n141 163.367
R2028 B.n522 B.n141 163.367
R2029 B.n522 B.n521 163.367
R2030 B.n521 B.n520 163.367
R2031 B.n520 B.n143 163.367
R2032 B.n516 B.n143 163.367
R2033 B.n516 B.n515 163.367
R2034 B.n515 B.n514 163.367
R2035 B.n514 B.n145 163.367
R2036 B.n510 B.n145 163.367
R2037 B.n510 B.n509 163.367
R2038 B.n509 B.n508 163.367
R2039 B.n508 B.n147 163.367
R2040 B.n853 B.n852 163.367
R2041 B.n852 B.n29 163.367
R2042 B.n848 B.n29 163.367
R2043 B.n848 B.n847 163.367
R2044 B.n847 B.n846 163.367
R2045 B.n846 B.n31 163.367
R2046 B.n842 B.n31 163.367
R2047 B.n842 B.n841 163.367
R2048 B.n841 B.n840 163.367
R2049 B.n840 B.n33 163.367
R2050 B.n836 B.n33 163.367
R2051 B.n836 B.n835 163.367
R2052 B.n835 B.n834 163.367
R2053 B.n834 B.n35 163.367
R2054 B.n830 B.n35 163.367
R2055 B.n830 B.n829 163.367
R2056 B.n829 B.n828 163.367
R2057 B.n828 B.n37 163.367
R2058 B.n824 B.n37 163.367
R2059 B.n824 B.n823 163.367
R2060 B.n823 B.n822 163.367
R2061 B.n822 B.n39 163.367
R2062 B.n818 B.n39 163.367
R2063 B.n818 B.n817 163.367
R2064 B.n817 B.n816 163.367
R2065 B.n816 B.n41 163.367
R2066 B.n812 B.n41 163.367
R2067 B.n812 B.n811 163.367
R2068 B.n811 B.n810 163.367
R2069 B.n810 B.n43 163.367
R2070 B.n806 B.n43 163.367
R2071 B.n806 B.n805 163.367
R2072 B.n805 B.n804 163.367
R2073 B.n804 B.n45 163.367
R2074 B.n800 B.n45 163.367
R2075 B.n800 B.n799 163.367
R2076 B.n799 B.n798 163.367
R2077 B.n798 B.n47 163.367
R2078 B.n794 B.n47 163.367
R2079 B.n794 B.n793 163.367
R2080 B.n793 B.n792 163.367
R2081 B.n792 B.n49 163.367
R2082 B.n788 B.n49 163.367
R2083 B.n788 B.n787 163.367
R2084 B.n787 B.n786 163.367
R2085 B.n786 B.n51 163.367
R2086 B.n782 B.n51 163.367
R2087 B.n782 B.n781 163.367
R2088 B.n781 B.n780 163.367
R2089 B.n780 B.n53 163.367
R2090 B.n776 B.n53 163.367
R2091 B.n776 B.n775 163.367
R2092 B.n775 B.n774 163.367
R2093 B.n774 B.n55 163.367
R2094 B.n770 B.n55 163.367
R2095 B.n770 B.n769 163.367
R2096 B.n769 B.n768 163.367
R2097 B.n768 B.n57 163.367
R2098 B.n763 B.n57 163.367
R2099 B.n763 B.n762 163.367
R2100 B.n762 B.n761 163.367
R2101 B.n761 B.n61 163.367
R2102 B.n757 B.n61 163.367
R2103 B.n757 B.n756 163.367
R2104 B.n756 B.n755 163.367
R2105 B.n755 B.n63 163.367
R2106 B.n750 B.n63 163.367
R2107 B.n750 B.n749 163.367
R2108 B.n749 B.n748 163.367
R2109 B.n748 B.n67 163.367
R2110 B.n744 B.n67 163.367
R2111 B.n744 B.n743 163.367
R2112 B.n743 B.n742 163.367
R2113 B.n742 B.n69 163.367
R2114 B.n738 B.n69 163.367
R2115 B.n738 B.n737 163.367
R2116 B.n737 B.n736 163.367
R2117 B.n736 B.n71 163.367
R2118 B.n732 B.n71 163.367
R2119 B.n732 B.n731 163.367
R2120 B.n731 B.n730 163.367
R2121 B.n730 B.n73 163.367
R2122 B.n726 B.n73 163.367
R2123 B.n726 B.n725 163.367
R2124 B.n725 B.n724 163.367
R2125 B.n724 B.n75 163.367
R2126 B.n720 B.n75 163.367
R2127 B.n720 B.n719 163.367
R2128 B.n719 B.n718 163.367
R2129 B.n718 B.n77 163.367
R2130 B.n714 B.n77 163.367
R2131 B.n714 B.n713 163.367
R2132 B.n713 B.n712 163.367
R2133 B.n712 B.n79 163.367
R2134 B.n708 B.n79 163.367
R2135 B.n708 B.n707 163.367
R2136 B.n707 B.n706 163.367
R2137 B.n706 B.n81 163.367
R2138 B.n702 B.n81 163.367
R2139 B.n702 B.n701 163.367
R2140 B.n701 B.n700 163.367
R2141 B.n700 B.n83 163.367
R2142 B.n696 B.n83 163.367
R2143 B.n696 B.n695 163.367
R2144 B.n695 B.n694 163.367
R2145 B.n694 B.n85 163.367
R2146 B.n690 B.n85 163.367
R2147 B.n690 B.n689 163.367
R2148 B.n689 B.n688 163.367
R2149 B.n688 B.n87 163.367
R2150 B.n684 B.n87 163.367
R2151 B.n684 B.n683 163.367
R2152 B.n683 B.n682 163.367
R2153 B.n682 B.n89 163.367
R2154 B.n678 B.n89 163.367
R2155 B.n678 B.n677 163.367
R2156 B.n677 B.n676 163.367
R2157 B.n676 B.n91 163.367
R2158 B.n672 B.n91 163.367
R2159 B.n672 B.n671 163.367
R2160 B.n671 B.n670 163.367
R2161 B.n670 B.n93 163.367
R2162 B.n666 B.n93 163.367
R2163 B.n666 B.n665 163.367
R2164 B.n854 B.n27 163.367
R2165 B.n858 B.n27 163.367
R2166 B.n859 B.n858 163.367
R2167 B.n860 B.n859 163.367
R2168 B.n860 B.n25 163.367
R2169 B.n864 B.n25 163.367
R2170 B.n865 B.n864 163.367
R2171 B.n866 B.n865 163.367
R2172 B.n866 B.n23 163.367
R2173 B.n870 B.n23 163.367
R2174 B.n871 B.n870 163.367
R2175 B.n872 B.n871 163.367
R2176 B.n872 B.n21 163.367
R2177 B.n876 B.n21 163.367
R2178 B.n877 B.n876 163.367
R2179 B.n878 B.n877 163.367
R2180 B.n878 B.n19 163.367
R2181 B.n882 B.n19 163.367
R2182 B.n883 B.n882 163.367
R2183 B.n884 B.n883 163.367
R2184 B.n884 B.n17 163.367
R2185 B.n888 B.n17 163.367
R2186 B.n889 B.n888 163.367
R2187 B.n890 B.n889 163.367
R2188 B.n890 B.n15 163.367
R2189 B.n894 B.n15 163.367
R2190 B.n895 B.n894 163.367
R2191 B.n896 B.n895 163.367
R2192 B.n896 B.n13 163.367
R2193 B.n900 B.n13 163.367
R2194 B.n901 B.n900 163.367
R2195 B.n902 B.n901 163.367
R2196 B.n902 B.n11 163.367
R2197 B.n906 B.n11 163.367
R2198 B.n907 B.n906 163.367
R2199 B.n908 B.n907 163.367
R2200 B.n908 B.n9 163.367
R2201 B.n912 B.n9 163.367
R2202 B.n913 B.n912 163.367
R2203 B.n914 B.n913 163.367
R2204 B.n914 B.n7 163.367
R2205 B.n918 B.n7 163.367
R2206 B.n919 B.n918 163.367
R2207 B.n920 B.n919 163.367
R2208 B.n920 B.n5 163.367
R2209 B.n924 B.n5 163.367
R2210 B.n925 B.n924 163.367
R2211 B.n926 B.n925 163.367
R2212 B.n926 B.n3 163.367
R2213 B.n930 B.n3 163.367
R2214 B.n931 B.n930 163.367
R2215 B.n237 B.n2 163.367
R2216 B.n240 B.n237 163.367
R2217 B.n241 B.n240 163.367
R2218 B.n242 B.n241 163.367
R2219 B.n242 B.n235 163.367
R2220 B.n246 B.n235 163.367
R2221 B.n247 B.n246 163.367
R2222 B.n248 B.n247 163.367
R2223 B.n248 B.n233 163.367
R2224 B.n252 B.n233 163.367
R2225 B.n253 B.n252 163.367
R2226 B.n254 B.n253 163.367
R2227 B.n254 B.n231 163.367
R2228 B.n258 B.n231 163.367
R2229 B.n259 B.n258 163.367
R2230 B.n260 B.n259 163.367
R2231 B.n260 B.n229 163.367
R2232 B.n264 B.n229 163.367
R2233 B.n265 B.n264 163.367
R2234 B.n266 B.n265 163.367
R2235 B.n266 B.n227 163.367
R2236 B.n270 B.n227 163.367
R2237 B.n271 B.n270 163.367
R2238 B.n272 B.n271 163.367
R2239 B.n272 B.n225 163.367
R2240 B.n276 B.n225 163.367
R2241 B.n277 B.n276 163.367
R2242 B.n278 B.n277 163.367
R2243 B.n278 B.n223 163.367
R2244 B.n282 B.n223 163.367
R2245 B.n283 B.n282 163.367
R2246 B.n284 B.n283 163.367
R2247 B.n284 B.n221 163.367
R2248 B.n288 B.n221 163.367
R2249 B.n289 B.n288 163.367
R2250 B.n290 B.n289 163.367
R2251 B.n290 B.n219 163.367
R2252 B.n294 B.n219 163.367
R2253 B.n295 B.n294 163.367
R2254 B.n296 B.n295 163.367
R2255 B.n296 B.n217 163.367
R2256 B.n300 B.n217 163.367
R2257 B.n301 B.n300 163.367
R2258 B.n302 B.n301 163.367
R2259 B.n302 B.n215 163.367
R2260 B.n306 B.n215 163.367
R2261 B.n307 B.n306 163.367
R2262 B.n308 B.n307 163.367
R2263 B.n308 B.n213 163.367
R2264 B.n312 B.n213 163.367
R2265 B.n313 B.n312 163.367
R2266 B.n401 B.n183 59.5399
R2267 B.n416 B.n415 59.5399
R2268 B.n752 B.n65 59.5399
R2269 B.n766 B.n59 59.5399
R2270 B.n183 B.n182 58.7641
R2271 B.n415 B.n414 58.7641
R2272 B.n65 B.n64 58.7641
R2273 B.n59 B.n58 58.7641
R2274 B.n855 B.n28 36.9956
R2275 B.n663 B.n94 36.9956
R2276 B.n506 B.n505 36.9956
R2277 B.n315 B.n212 36.9956
R2278 B B.n933 18.0485
R2279 B.n856 B.n855 10.6151
R2280 B.n857 B.n856 10.6151
R2281 B.n857 B.n26 10.6151
R2282 B.n861 B.n26 10.6151
R2283 B.n862 B.n861 10.6151
R2284 B.n863 B.n862 10.6151
R2285 B.n863 B.n24 10.6151
R2286 B.n867 B.n24 10.6151
R2287 B.n868 B.n867 10.6151
R2288 B.n869 B.n868 10.6151
R2289 B.n869 B.n22 10.6151
R2290 B.n873 B.n22 10.6151
R2291 B.n874 B.n873 10.6151
R2292 B.n875 B.n874 10.6151
R2293 B.n875 B.n20 10.6151
R2294 B.n879 B.n20 10.6151
R2295 B.n880 B.n879 10.6151
R2296 B.n881 B.n880 10.6151
R2297 B.n881 B.n18 10.6151
R2298 B.n885 B.n18 10.6151
R2299 B.n886 B.n885 10.6151
R2300 B.n887 B.n886 10.6151
R2301 B.n887 B.n16 10.6151
R2302 B.n891 B.n16 10.6151
R2303 B.n892 B.n891 10.6151
R2304 B.n893 B.n892 10.6151
R2305 B.n893 B.n14 10.6151
R2306 B.n897 B.n14 10.6151
R2307 B.n898 B.n897 10.6151
R2308 B.n899 B.n898 10.6151
R2309 B.n899 B.n12 10.6151
R2310 B.n903 B.n12 10.6151
R2311 B.n904 B.n903 10.6151
R2312 B.n905 B.n904 10.6151
R2313 B.n905 B.n10 10.6151
R2314 B.n909 B.n10 10.6151
R2315 B.n910 B.n909 10.6151
R2316 B.n911 B.n910 10.6151
R2317 B.n911 B.n8 10.6151
R2318 B.n915 B.n8 10.6151
R2319 B.n916 B.n915 10.6151
R2320 B.n917 B.n916 10.6151
R2321 B.n917 B.n6 10.6151
R2322 B.n921 B.n6 10.6151
R2323 B.n922 B.n921 10.6151
R2324 B.n923 B.n922 10.6151
R2325 B.n923 B.n4 10.6151
R2326 B.n927 B.n4 10.6151
R2327 B.n928 B.n927 10.6151
R2328 B.n929 B.n928 10.6151
R2329 B.n929 B.n0 10.6151
R2330 B.n851 B.n28 10.6151
R2331 B.n851 B.n850 10.6151
R2332 B.n850 B.n849 10.6151
R2333 B.n849 B.n30 10.6151
R2334 B.n845 B.n30 10.6151
R2335 B.n845 B.n844 10.6151
R2336 B.n844 B.n843 10.6151
R2337 B.n843 B.n32 10.6151
R2338 B.n839 B.n32 10.6151
R2339 B.n839 B.n838 10.6151
R2340 B.n838 B.n837 10.6151
R2341 B.n837 B.n34 10.6151
R2342 B.n833 B.n34 10.6151
R2343 B.n833 B.n832 10.6151
R2344 B.n832 B.n831 10.6151
R2345 B.n831 B.n36 10.6151
R2346 B.n827 B.n36 10.6151
R2347 B.n827 B.n826 10.6151
R2348 B.n826 B.n825 10.6151
R2349 B.n825 B.n38 10.6151
R2350 B.n821 B.n38 10.6151
R2351 B.n821 B.n820 10.6151
R2352 B.n820 B.n819 10.6151
R2353 B.n819 B.n40 10.6151
R2354 B.n815 B.n40 10.6151
R2355 B.n815 B.n814 10.6151
R2356 B.n814 B.n813 10.6151
R2357 B.n813 B.n42 10.6151
R2358 B.n809 B.n42 10.6151
R2359 B.n809 B.n808 10.6151
R2360 B.n808 B.n807 10.6151
R2361 B.n807 B.n44 10.6151
R2362 B.n803 B.n44 10.6151
R2363 B.n803 B.n802 10.6151
R2364 B.n802 B.n801 10.6151
R2365 B.n801 B.n46 10.6151
R2366 B.n797 B.n46 10.6151
R2367 B.n797 B.n796 10.6151
R2368 B.n796 B.n795 10.6151
R2369 B.n795 B.n48 10.6151
R2370 B.n791 B.n48 10.6151
R2371 B.n791 B.n790 10.6151
R2372 B.n790 B.n789 10.6151
R2373 B.n789 B.n50 10.6151
R2374 B.n785 B.n50 10.6151
R2375 B.n785 B.n784 10.6151
R2376 B.n784 B.n783 10.6151
R2377 B.n783 B.n52 10.6151
R2378 B.n779 B.n52 10.6151
R2379 B.n779 B.n778 10.6151
R2380 B.n778 B.n777 10.6151
R2381 B.n777 B.n54 10.6151
R2382 B.n773 B.n54 10.6151
R2383 B.n773 B.n772 10.6151
R2384 B.n772 B.n771 10.6151
R2385 B.n771 B.n56 10.6151
R2386 B.n767 B.n56 10.6151
R2387 B.n765 B.n764 10.6151
R2388 B.n764 B.n60 10.6151
R2389 B.n760 B.n60 10.6151
R2390 B.n760 B.n759 10.6151
R2391 B.n759 B.n758 10.6151
R2392 B.n758 B.n62 10.6151
R2393 B.n754 B.n62 10.6151
R2394 B.n754 B.n753 10.6151
R2395 B.n751 B.n66 10.6151
R2396 B.n747 B.n66 10.6151
R2397 B.n747 B.n746 10.6151
R2398 B.n746 B.n745 10.6151
R2399 B.n745 B.n68 10.6151
R2400 B.n741 B.n68 10.6151
R2401 B.n741 B.n740 10.6151
R2402 B.n740 B.n739 10.6151
R2403 B.n739 B.n70 10.6151
R2404 B.n735 B.n70 10.6151
R2405 B.n735 B.n734 10.6151
R2406 B.n734 B.n733 10.6151
R2407 B.n733 B.n72 10.6151
R2408 B.n729 B.n72 10.6151
R2409 B.n729 B.n728 10.6151
R2410 B.n728 B.n727 10.6151
R2411 B.n727 B.n74 10.6151
R2412 B.n723 B.n74 10.6151
R2413 B.n723 B.n722 10.6151
R2414 B.n722 B.n721 10.6151
R2415 B.n721 B.n76 10.6151
R2416 B.n717 B.n76 10.6151
R2417 B.n717 B.n716 10.6151
R2418 B.n716 B.n715 10.6151
R2419 B.n715 B.n78 10.6151
R2420 B.n711 B.n78 10.6151
R2421 B.n711 B.n710 10.6151
R2422 B.n710 B.n709 10.6151
R2423 B.n709 B.n80 10.6151
R2424 B.n705 B.n80 10.6151
R2425 B.n705 B.n704 10.6151
R2426 B.n704 B.n703 10.6151
R2427 B.n703 B.n82 10.6151
R2428 B.n699 B.n82 10.6151
R2429 B.n699 B.n698 10.6151
R2430 B.n698 B.n697 10.6151
R2431 B.n697 B.n84 10.6151
R2432 B.n693 B.n84 10.6151
R2433 B.n693 B.n692 10.6151
R2434 B.n692 B.n691 10.6151
R2435 B.n691 B.n86 10.6151
R2436 B.n687 B.n86 10.6151
R2437 B.n687 B.n686 10.6151
R2438 B.n686 B.n685 10.6151
R2439 B.n685 B.n88 10.6151
R2440 B.n681 B.n88 10.6151
R2441 B.n681 B.n680 10.6151
R2442 B.n680 B.n679 10.6151
R2443 B.n679 B.n90 10.6151
R2444 B.n675 B.n90 10.6151
R2445 B.n675 B.n674 10.6151
R2446 B.n674 B.n673 10.6151
R2447 B.n673 B.n92 10.6151
R2448 B.n669 B.n92 10.6151
R2449 B.n669 B.n668 10.6151
R2450 B.n668 B.n667 10.6151
R2451 B.n667 B.n94 10.6151
R2452 B.n663 B.n662 10.6151
R2453 B.n662 B.n661 10.6151
R2454 B.n661 B.n96 10.6151
R2455 B.n657 B.n96 10.6151
R2456 B.n657 B.n656 10.6151
R2457 B.n656 B.n655 10.6151
R2458 B.n655 B.n98 10.6151
R2459 B.n651 B.n98 10.6151
R2460 B.n651 B.n650 10.6151
R2461 B.n650 B.n649 10.6151
R2462 B.n649 B.n100 10.6151
R2463 B.n645 B.n100 10.6151
R2464 B.n645 B.n644 10.6151
R2465 B.n644 B.n643 10.6151
R2466 B.n643 B.n102 10.6151
R2467 B.n639 B.n102 10.6151
R2468 B.n639 B.n638 10.6151
R2469 B.n638 B.n637 10.6151
R2470 B.n637 B.n104 10.6151
R2471 B.n633 B.n104 10.6151
R2472 B.n633 B.n632 10.6151
R2473 B.n632 B.n631 10.6151
R2474 B.n631 B.n106 10.6151
R2475 B.n627 B.n106 10.6151
R2476 B.n627 B.n626 10.6151
R2477 B.n626 B.n625 10.6151
R2478 B.n625 B.n108 10.6151
R2479 B.n621 B.n108 10.6151
R2480 B.n621 B.n620 10.6151
R2481 B.n620 B.n619 10.6151
R2482 B.n619 B.n110 10.6151
R2483 B.n615 B.n110 10.6151
R2484 B.n615 B.n614 10.6151
R2485 B.n614 B.n613 10.6151
R2486 B.n613 B.n112 10.6151
R2487 B.n609 B.n112 10.6151
R2488 B.n609 B.n608 10.6151
R2489 B.n608 B.n607 10.6151
R2490 B.n607 B.n114 10.6151
R2491 B.n603 B.n114 10.6151
R2492 B.n603 B.n602 10.6151
R2493 B.n602 B.n601 10.6151
R2494 B.n601 B.n116 10.6151
R2495 B.n597 B.n116 10.6151
R2496 B.n597 B.n596 10.6151
R2497 B.n596 B.n595 10.6151
R2498 B.n595 B.n118 10.6151
R2499 B.n591 B.n118 10.6151
R2500 B.n591 B.n590 10.6151
R2501 B.n590 B.n589 10.6151
R2502 B.n589 B.n120 10.6151
R2503 B.n585 B.n120 10.6151
R2504 B.n585 B.n584 10.6151
R2505 B.n584 B.n583 10.6151
R2506 B.n583 B.n122 10.6151
R2507 B.n579 B.n122 10.6151
R2508 B.n579 B.n578 10.6151
R2509 B.n578 B.n577 10.6151
R2510 B.n577 B.n124 10.6151
R2511 B.n573 B.n124 10.6151
R2512 B.n573 B.n572 10.6151
R2513 B.n572 B.n571 10.6151
R2514 B.n571 B.n126 10.6151
R2515 B.n567 B.n126 10.6151
R2516 B.n567 B.n566 10.6151
R2517 B.n566 B.n565 10.6151
R2518 B.n565 B.n128 10.6151
R2519 B.n561 B.n128 10.6151
R2520 B.n561 B.n560 10.6151
R2521 B.n560 B.n559 10.6151
R2522 B.n559 B.n130 10.6151
R2523 B.n555 B.n130 10.6151
R2524 B.n555 B.n554 10.6151
R2525 B.n554 B.n553 10.6151
R2526 B.n553 B.n132 10.6151
R2527 B.n549 B.n132 10.6151
R2528 B.n549 B.n548 10.6151
R2529 B.n548 B.n547 10.6151
R2530 B.n547 B.n134 10.6151
R2531 B.n543 B.n134 10.6151
R2532 B.n543 B.n542 10.6151
R2533 B.n542 B.n541 10.6151
R2534 B.n541 B.n136 10.6151
R2535 B.n537 B.n136 10.6151
R2536 B.n537 B.n536 10.6151
R2537 B.n536 B.n535 10.6151
R2538 B.n535 B.n138 10.6151
R2539 B.n531 B.n138 10.6151
R2540 B.n531 B.n530 10.6151
R2541 B.n530 B.n529 10.6151
R2542 B.n529 B.n140 10.6151
R2543 B.n525 B.n140 10.6151
R2544 B.n525 B.n524 10.6151
R2545 B.n524 B.n523 10.6151
R2546 B.n523 B.n142 10.6151
R2547 B.n519 B.n142 10.6151
R2548 B.n519 B.n518 10.6151
R2549 B.n518 B.n517 10.6151
R2550 B.n517 B.n144 10.6151
R2551 B.n513 B.n144 10.6151
R2552 B.n513 B.n512 10.6151
R2553 B.n512 B.n511 10.6151
R2554 B.n511 B.n146 10.6151
R2555 B.n507 B.n146 10.6151
R2556 B.n507 B.n506 10.6151
R2557 B.n238 B.n1 10.6151
R2558 B.n239 B.n238 10.6151
R2559 B.n239 B.n236 10.6151
R2560 B.n243 B.n236 10.6151
R2561 B.n244 B.n243 10.6151
R2562 B.n245 B.n244 10.6151
R2563 B.n245 B.n234 10.6151
R2564 B.n249 B.n234 10.6151
R2565 B.n250 B.n249 10.6151
R2566 B.n251 B.n250 10.6151
R2567 B.n251 B.n232 10.6151
R2568 B.n255 B.n232 10.6151
R2569 B.n256 B.n255 10.6151
R2570 B.n257 B.n256 10.6151
R2571 B.n257 B.n230 10.6151
R2572 B.n261 B.n230 10.6151
R2573 B.n262 B.n261 10.6151
R2574 B.n263 B.n262 10.6151
R2575 B.n263 B.n228 10.6151
R2576 B.n267 B.n228 10.6151
R2577 B.n268 B.n267 10.6151
R2578 B.n269 B.n268 10.6151
R2579 B.n269 B.n226 10.6151
R2580 B.n273 B.n226 10.6151
R2581 B.n274 B.n273 10.6151
R2582 B.n275 B.n274 10.6151
R2583 B.n275 B.n224 10.6151
R2584 B.n279 B.n224 10.6151
R2585 B.n280 B.n279 10.6151
R2586 B.n281 B.n280 10.6151
R2587 B.n281 B.n222 10.6151
R2588 B.n285 B.n222 10.6151
R2589 B.n286 B.n285 10.6151
R2590 B.n287 B.n286 10.6151
R2591 B.n287 B.n220 10.6151
R2592 B.n291 B.n220 10.6151
R2593 B.n292 B.n291 10.6151
R2594 B.n293 B.n292 10.6151
R2595 B.n293 B.n218 10.6151
R2596 B.n297 B.n218 10.6151
R2597 B.n298 B.n297 10.6151
R2598 B.n299 B.n298 10.6151
R2599 B.n299 B.n216 10.6151
R2600 B.n303 B.n216 10.6151
R2601 B.n304 B.n303 10.6151
R2602 B.n305 B.n304 10.6151
R2603 B.n305 B.n214 10.6151
R2604 B.n309 B.n214 10.6151
R2605 B.n310 B.n309 10.6151
R2606 B.n311 B.n310 10.6151
R2607 B.n311 B.n212 10.6151
R2608 B.n316 B.n315 10.6151
R2609 B.n317 B.n316 10.6151
R2610 B.n317 B.n210 10.6151
R2611 B.n321 B.n210 10.6151
R2612 B.n322 B.n321 10.6151
R2613 B.n323 B.n322 10.6151
R2614 B.n323 B.n208 10.6151
R2615 B.n327 B.n208 10.6151
R2616 B.n328 B.n327 10.6151
R2617 B.n329 B.n328 10.6151
R2618 B.n329 B.n206 10.6151
R2619 B.n333 B.n206 10.6151
R2620 B.n334 B.n333 10.6151
R2621 B.n335 B.n334 10.6151
R2622 B.n335 B.n204 10.6151
R2623 B.n339 B.n204 10.6151
R2624 B.n340 B.n339 10.6151
R2625 B.n341 B.n340 10.6151
R2626 B.n341 B.n202 10.6151
R2627 B.n345 B.n202 10.6151
R2628 B.n346 B.n345 10.6151
R2629 B.n347 B.n346 10.6151
R2630 B.n347 B.n200 10.6151
R2631 B.n351 B.n200 10.6151
R2632 B.n352 B.n351 10.6151
R2633 B.n353 B.n352 10.6151
R2634 B.n353 B.n198 10.6151
R2635 B.n357 B.n198 10.6151
R2636 B.n358 B.n357 10.6151
R2637 B.n359 B.n358 10.6151
R2638 B.n359 B.n196 10.6151
R2639 B.n363 B.n196 10.6151
R2640 B.n364 B.n363 10.6151
R2641 B.n365 B.n364 10.6151
R2642 B.n365 B.n194 10.6151
R2643 B.n369 B.n194 10.6151
R2644 B.n370 B.n369 10.6151
R2645 B.n371 B.n370 10.6151
R2646 B.n371 B.n192 10.6151
R2647 B.n375 B.n192 10.6151
R2648 B.n376 B.n375 10.6151
R2649 B.n377 B.n376 10.6151
R2650 B.n377 B.n190 10.6151
R2651 B.n381 B.n190 10.6151
R2652 B.n382 B.n381 10.6151
R2653 B.n383 B.n382 10.6151
R2654 B.n383 B.n188 10.6151
R2655 B.n387 B.n188 10.6151
R2656 B.n388 B.n387 10.6151
R2657 B.n389 B.n388 10.6151
R2658 B.n389 B.n186 10.6151
R2659 B.n393 B.n186 10.6151
R2660 B.n394 B.n393 10.6151
R2661 B.n395 B.n394 10.6151
R2662 B.n395 B.n184 10.6151
R2663 B.n399 B.n184 10.6151
R2664 B.n400 B.n399 10.6151
R2665 B.n402 B.n180 10.6151
R2666 B.n406 B.n180 10.6151
R2667 B.n407 B.n406 10.6151
R2668 B.n408 B.n407 10.6151
R2669 B.n408 B.n178 10.6151
R2670 B.n412 B.n178 10.6151
R2671 B.n413 B.n412 10.6151
R2672 B.n417 B.n413 10.6151
R2673 B.n421 B.n176 10.6151
R2674 B.n422 B.n421 10.6151
R2675 B.n423 B.n422 10.6151
R2676 B.n423 B.n174 10.6151
R2677 B.n427 B.n174 10.6151
R2678 B.n428 B.n427 10.6151
R2679 B.n429 B.n428 10.6151
R2680 B.n429 B.n172 10.6151
R2681 B.n433 B.n172 10.6151
R2682 B.n434 B.n433 10.6151
R2683 B.n435 B.n434 10.6151
R2684 B.n435 B.n170 10.6151
R2685 B.n439 B.n170 10.6151
R2686 B.n440 B.n439 10.6151
R2687 B.n441 B.n440 10.6151
R2688 B.n441 B.n168 10.6151
R2689 B.n445 B.n168 10.6151
R2690 B.n446 B.n445 10.6151
R2691 B.n447 B.n446 10.6151
R2692 B.n447 B.n166 10.6151
R2693 B.n451 B.n166 10.6151
R2694 B.n452 B.n451 10.6151
R2695 B.n453 B.n452 10.6151
R2696 B.n453 B.n164 10.6151
R2697 B.n457 B.n164 10.6151
R2698 B.n458 B.n457 10.6151
R2699 B.n459 B.n458 10.6151
R2700 B.n459 B.n162 10.6151
R2701 B.n463 B.n162 10.6151
R2702 B.n464 B.n463 10.6151
R2703 B.n465 B.n464 10.6151
R2704 B.n465 B.n160 10.6151
R2705 B.n469 B.n160 10.6151
R2706 B.n470 B.n469 10.6151
R2707 B.n471 B.n470 10.6151
R2708 B.n471 B.n158 10.6151
R2709 B.n475 B.n158 10.6151
R2710 B.n476 B.n475 10.6151
R2711 B.n477 B.n476 10.6151
R2712 B.n477 B.n156 10.6151
R2713 B.n481 B.n156 10.6151
R2714 B.n482 B.n481 10.6151
R2715 B.n483 B.n482 10.6151
R2716 B.n483 B.n154 10.6151
R2717 B.n487 B.n154 10.6151
R2718 B.n488 B.n487 10.6151
R2719 B.n489 B.n488 10.6151
R2720 B.n489 B.n152 10.6151
R2721 B.n493 B.n152 10.6151
R2722 B.n494 B.n493 10.6151
R2723 B.n495 B.n494 10.6151
R2724 B.n495 B.n150 10.6151
R2725 B.n499 B.n150 10.6151
R2726 B.n500 B.n499 10.6151
R2727 B.n501 B.n500 10.6151
R2728 B.n501 B.n148 10.6151
R2729 B.n505 B.n148 10.6151
R2730 B.n933 B.n0 8.11757
R2731 B.n933 B.n1 8.11757
R2732 B.n766 B.n765 6.5566
R2733 B.n753 B.n752 6.5566
R2734 B.n402 B.n401 6.5566
R2735 B.n417 B.n416 6.5566
R2736 B.n767 B.n766 4.05904
R2737 B.n752 B.n751 4.05904
R2738 B.n401 B.n400 4.05904
R2739 B.n416 B.n176 4.05904
R2740 VN.n8 VN.t2 187.621
R2741 VN.n39 VN.t4 187.621
R2742 VN.n59 VN.n31 161.3
R2743 VN.n58 VN.n57 161.3
R2744 VN.n56 VN.n32 161.3
R2745 VN.n55 VN.n54 161.3
R2746 VN.n53 VN.n33 161.3
R2747 VN.n52 VN.n51 161.3
R2748 VN.n50 VN.n49 161.3
R2749 VN.n48 VN.n35 161.3
R2750 VN.n47 VN.n46 161.3
R2751 VN.n45 VN.n36 161.3
R2752 VN.n44 VN.n43 161.3
R2753 VN.n42 VN.n37 161.3
R2754 VN.n41 VN.n40 161.3
R2755 VN.n28 VN.n0 161.3
R2756 VN.n27 VN.n26 161.3
R2757 VN.n25 VN.n1 161.3
R2758 VN.n24 VN.n23 161.3
R2759 VN.n22 VN.n2 161.3
R2760 VN.n21 VN.n20 161.3
R2761 VN.n19 VN.n18 161.3
R2762 VN.n17 VN.n4 161.3
R2763 VN.n16 VN.n15 161.3
R2764 VN.n14 VN.n5 161.3
R2765 VN.n13 VN.n12 161.3
R2766 VN.n11 VN.n6 161.3
R2767 VN.n10 VN.n9 161.3
R2768 VN.n7 VN.t7 156.739
R2769 VN.n3 VN.t3 156.739
R2770 VN.n29 VN.t6 156.739
R2771 VN.n38 VN.t5 156.739
R2772 VN.n34 VN.t0 156.739
R2773 VN.n60 VN.t1 156.739
R2774 VN.n30 VN.n29 108.695
R2775 VN.n61 VN.n60 108.695
R2776 VN.n8 VN.n7 72.8488
R2777 VN.n39 VN.n38 72.8488
R2778 VN VN.n61 55.7785
R2779 VN.n23 VN.n1 43.4833
R2780 VN.n54 VN.n32 43.4833
R2781 VN.n12 VN.n5 40.577
R2782 VN.n16 VN.n5 40.577
R2783 VN.n43 VN.n36 40.577
R2784 VN.n47 VN.n36 40.577
R2785 VN.n23 VN.n22 37.6707
R2786 VN.n54 VN.n53 37.6707
R2787 VN.n11 VN.n10 24.5923
R2788 VN.n12 VN.n11 24.5923
R2789 VN.n17 VN.n16 24.5923
R2790 VN.n18 VN.n17 24.5923
R2791 VN.n22 VN.n21 24.5923
R2792 VN.n27 VN.n1 24.5923
R2793 VN.n28 VN.n27 24.5923
R2794 VN.n43 VN.n42 24.5923
R2795 VN.n42 VN.n41 24.5923
R2796 VN.n53 VN.n52 24.5923
R2797 VN.n49 VN.n48 24.5923
R2798 VN.n48 VN.n47 24.5923
R2799 VN.n59 VN.n58 24.5923
R2800 VN.n58 VN.n32 24.5923
R2801 VN.n21 VN.n3 23.8546
R2802 VN.n52 VN.n34 23.8546
R2803 VN.n40 VN.n39 7.34013
R2804 VN.n9 VN.n8 7.34013
R2805 VN.n29 VN.n28 2.21377
R2806 VN.n60 VN.n59 2.21377
R2807 VN.n10 VN.n7 0.738255
R2808 VN.n18 VN.n3 0.738255
R2809 VN.n41 VN.n38 0.738255
R2810 VN.n49 VN.n34 0.738255
R2811 VN.n61 VN.n31 0.278335
R2812 VN.n30 VN.n0 0.278335
R2813 VN.n57 VN.n31 0.189894
R2814 VN.n57 VN.n56 0.189894
R2815 VN.n56 VN.n55 0.189894
R2816 VN.n55 VN.n33 0.189894
R2817 VN.n51 VN.n33 0.189894
R2818 VN.n51 VN.n50 0.189894
R2819 VN.n50 VN.n35 0.189894
R2820 VN.n46 VN.n35 0.189894
R2821 VN.n46 VN.n45 0.189894
R2822 VN.n45 VN.n44 0.189894
R2823 VN.n44 VN.n37 0.189894
R2824 VN.n40 VN.n37 0.189894
R2825 VN.n9 VN.n6 0.189894
R2826 VN.n13 VN.n6 0.189894
R2827 VN.n14 VN.n13 0.189894
R2828 VN.n15 VN.n14 0.189894
R2829 VN.n15 VN.n4 0.189894
R2830 VN.n19 VN.n4 0.189894
R2831 VN.n20 VN.n19 0.189894
R2832 VN.n20 VN.n2 0.189894
R2833 VN.n24 VN.n2 0.189894
R2834 VN.n25 VN.n24 0.189894
R2835 VN.n26 VN.n25 0.189894
R2836 VN.n26 VN.n0 0.189894
R2837 VN VN.n30 0.153485
R2838 VDD2.n2 VDD2.n1 71.0485
R2839 VDD2.n2 VDD2.n0 71.0485
R2840 VDD2 VDD2.n5 71.0456
R2841 VDD2.n4 VDD2.n3 69.798
R2842 VDD2.n4 VDD2.n2 50.6075
R2843 VDD2.n5 VDD2.t2 1.85158
R2844 VDD2.n5 VDD2.t3 1.85158
R2845 VDD2.n3 VDD2.t6 1.85158
R2846 VDD2.n3 VDD2.t7 1.85158
R2847 VDD2.n1 VDD2.t4 1.85158
R2848 VDD2.n1 VDD2.t1 1.85158
R2849 VDD2.n0 VDD2.t5 1.85158
R2850 VDD2.n0 VDD2.t0 1.85158
R2851 VDD2 VDD2.n4 1.36472
C0 VDD2 VP 0.53026f
C1 VDD1 VN 0.151857f
C2 VDD1 VTAIL 9.932151f
C3 VDD2 VN 12.6147f
C4 VDD2 VTAIL 9.98724f
C5 VDD1 VDD2 1.82674f
C6 B w_n4000_n4480# 11.8278f
C7 VP w_n4000_n4480# 8.793389f
C8 B VP 2.18917f
C9 VN w_n4000_n4480# 8.273809f
C10 VTAIL w_n4000_n4480# 5.45698f
C11 VN B 1.31765f
C12 VDD1 w_n4000_n4480# 2.13039f
C13 VTAIL B 6.86395f
C14 VN VP 8.81094f
C15 VTAIL VP 12.8038f
C16 VDD2 w_n4000_n4480# 2.24929f
C17 VDD1 B 1.82868f
C18 VDD1 VP 12.9917f
C19 VDD2 B 1.92785f
C20 VN VTAIL 12.789701f
C21 VDD2 VSUBS 2.052599f
C22 VDD1 VSUBS 2.71392f
C23 VTAIL VSUBS 1.605149f
C24 VN VSUBS 7.08182f
C25 VP VSUBS 3.88267f
C26 B VSUBS 5.586854f
C27 w_n4000_n4480# VSUBS 0.219216p
C28 VDD2.t5 VSUBS 0.369865f
C29 VDD2.t0 VSUBS 0.369865f
C30 VDD2.n0 VSUBS 3.08143f
C31 VDD2.t4 VSUBS 0.369865f
C32 VDD2.t1 VSUBS 0.369865f
C33 VDD2.n1 VSUBS 3.08143f
C34 VDD2.n2 VSUBS 4.526f
C35 VDD2.t6 VSUBS 0.369865f
C36 VDD2.t7 VSUBS 0.369865f
C37 VDD2.n3 VSUBS 3.06624f
C38 VDD2.n4 VSUBS 3.93225f
C39 VDD2.t2 VSUBS 0.369865f
C40 VDD2.t3 VSUBS 0.369865f
C41 VDD2.n5 VSUBS 3.08139f
C42 VN.n0 VSUBS 0.033912f
C43 VN.t6 VSUBS 3.35302f
C44 VN.n1 VSUBS 0.049953f
C45 VN.n2 VSUBS 0.025724f
C46 VN.t3 VSUBS 3.35302f
C47 VN.n3 VSUBS 1.16285f
C48 VN.n4 VSUBS 0.025724f
C49 VN.n5 VSUBS 0.020776f
C50 VN.n6 VSUBS 0.025724f
C51 VN.t7 VSUBS 3.35302f
C52 VN.n7 VSUBS 1.22941f
C53 VN.t2 VSUBS 3.5706f
C54 VN.n8 VSUBS 1.21447f
C55 VN.n9 VSUBS 0.25076f
C56 VN.n10 VSUBS 0.024859f
C57 VN.n11 VSUBS 0.047702f
C58 VN.n12 VSUBS 0.050856f
C59 VN.n13 VSUBS 0.025724f
C60 VN.n14 VSUBS 0.025724f
C61 VN.n15 VSUBS 0.025724f
C62 VN.n16 VSUBS 0.050856f
C63 VN.n17 VSUBS 0.047702f
C64 VN.n18 VSUBS 0.024859f
C65 VN.n19 VSUBS 0.025724f
C66 VN.n20 VSUBS 0.025724f
C67 VN.n21 VSUBS 0.046995f
C68 VN.n22 VSUBS 0.051463f
C69 VN.n23 VSUBS 0.021073f
C70 VN.n24 VSUBS 0.025724f
C71 VN.n25 VSUBS 0.025724f
C72 VN.n26 VSUBS 0.025724f
C73 VN.n27 VSUBS 0.047702f
C74 VN.n28 VSUBS 0.026272f
C75 VN.n29 VSUBS 1.24133f
C76 VN.n30 VSUBS 0.047259f
C77 VN.n31 VSUBS 0.033912f
C78 VN.t1 VSUBS 3.35302f
C79 VN.n32 VSUBS 0.049953f
C80 VN.n33 VSUBS 0.025724f
C81 VN.t0 VSUBS 3.35302f
C82 VN.n34 VSUBS 1.16285f
C83 VN.n35 VSUBS 0.025724f
C84 VN.n36 VSUBS 0.020776f
C85 VN.n37 VSUBS 0.025724f
C86 VN.t5 VSUBS 3.35302f
C87 VN.n38 VSUBS 1.22941f
C88 VN.t4 VSUBS 3.5706f
C89 VN.n39 VSUBS 1.21447f
C90 VN.n40 VSUBS 0.25076f
C91 VN.n41 VSUBS 0.024859f
C92 VN.n42 VSUBS 0.047702f
C93 VN.n43 VSUBS 0.050856f
C94 VN.n44 VSUBS 0.025724f
C95 VN.n45 VSUBS 0.025724f
C96 VN.n46 VSUBS 0.025724f
C97 VN.n47 VSUBS 0.050856f
C98 VN.n48 VSUBS 0.047702f
C99 VN.n49 VSUBS 0.024859f
C100 VN.n50 VSUBS 0.025724f
C101 VN.n51 VSUBS 0.025724f
C102 VN.n52 VSUBS 0.046995f
C103 VN.n53 VSUBS 0.051463f
C104 VN.n54 VSUBS 0.021073f
C105 VN.n55 VSUBS 0.025724f
C106 VN.n56 VSUBS 0.025724f
C107 VN.n57 VSUBS 0.025724f
C108 VN.n58 VSUBS 0.047702f
C109 VN.n59 VSUBS 0.026272f
C110 VN.n60 VSUBS 1.24133f
C111 VN.n61 VSUBS 1.68074f
C112 B.n0 VSUBS 0.00597f
C113 B.n1 VSUBS 0.00597f
C114 B.n2 VSUBS 0.008829f
C115 B.n3 VSUBS 0.006766f
C116 B.n4 VSUBS 0.006766f
C117 B.n5 VSUBS 0.006766f
C118 B.n6 VSUBS 0.006766f
C119 B.n7 VSUBS 0.006766f
C120 B.n8 VSUBS 0.006766f
C121 B.n9 VSUBS 0.006766f
C122 B.n10 VSUBS 0.006766f
C123 B.n11 VSUBS 0.006766f
C124 B.n12 VSUBS 0.006766f
C125 B.n13 VSUBS 0.006766f
C126 B.n14 VSUBS 0.006766f
C127 B.n15 VSUBS 0.006766f
C128 B.n16 VSUBS 0.006766f
C129 B.n17 VSUBS 0.006766f
C130 B.n18 VSUBS 0.006766f
C131 B.n19 VSUBS 0.006766f
C132 B.n20 VSUBS 0.006766f
C133 B.n21 VSUBS 0.006766f
C134 B.n22 VSUBS 0.006766f
C135 B.n23 VSUBS 0.006766f
C136 B.n24 VSUBS 0.006766f
C137 B.n25 VSUBS 0.006766f
C138 B.n26 VSUBS 0.006766f
C139 B.n27 VSUBS 0.006766f
C140 B.n28 VSUBS 0.017496f
C141 B.n29 VSUBS 0.006766f
C142 B.n30 VSUBS 0.006766f
C143 B.n31 VSUBS 0.006766f
C144 B.n32 VSUBS 0.006766f
C145 B.n33 VSUBS 0.006766f
C146 B.n34 VSUBS 0.006766f
C147 B.n35 VSUBS 0.006766f
C148 B.n36 VSUBS 0.006766f
C149 B.n37 VSUBS 0.006766f
C150 B.n38 VSUBS 0.006766f
C151 B.n39 VSUBS 0.006766f
C152 B.n40 VSUBS 0.006766f
C153 B.n41 VSUBS 0.006766f
C154 B.n42 VSUBS 0.006766f
C155 B.n43 VSUBS 0.006766f
C156 B.n44 VSUBS 0.006766f
C157 B.n45 VSUBS 0.006766f
C158 B.n46 VSUBS 0.006766f
C159 B.n47 VSUBS 0.006766f
C160 B.n48 VSUBS 0.006766f
C161 B.n49 VSUBS 0.006766f
C162 B.n50 VSUBS 0.006766f
C163 B.n51 VSUBS 0.006766f
C164 B.n52 VSUBS 0.006766f
C165 B.n53 VSUBS 0.006766f
C166 B.n54 VSUBS 0.006766f
C167 B.n55 VSUBS 0.006766f
C168 B.n56 VSUBS 0.006766f
C169 B.n57 VSUBS 0.006766f
C170 B.t1 VSUBS 0.329118f
C171 B.t2 VSUBS 0.362454f
C172 B.t0 VSUBS 2.04176f
C173 B.n58 VSUBS 0.558786f
C174 B.n59 VSUBS 0.312927f
C175 B.n60 VSUBS 0.006766f
C176 B.n61 VSUBS 0.006766f
C177 B.n62 VSUBS 0.006766f
C178 B.n63 VSUBS 0.006766f
C179 B.t7 VSUBS 0.329121f
C180 B.t8 VSUBS 0.362457f
C181 B.t6 VSUBS 2.04176f
C182 B.n64 VSUBS 0.558783f
C183 B.n65 VSUBS 0.312923f
C184 B.n66 VSUBS 0.006766f
C185 B.n67 VSUBS 0.006766f
C186 B.n68 VSUBS 0.006766f
C187 B.n69 VSUBS 0.006766f
C188 B.n70 VSUBS 0.006766f
C189 B.n71 VSUBS 0.006766f
C190 B.n72 VSUBS 0.006766f
C191 B.n73 VSUBS 0.006766f
C192 B.n74 VSUBS 0.006766f
C193 B.n75 VSUBS 0.006766f
C194 B.n76 VSUBS 0.006766f
C195 B.n77 VSUBS 0.006766f
C196 B.n78 VSUBS 0.006766f
C197 B.n79 VSUBS 0.006766f
C198 B.n80 VSUBS 0.006766f
C199 B.n81 VSUBS 0.006766f
C200 B.n82 VSUBS 0.006766f
C201 B.n83 VSUBS 0.006766f
C202 B.n84 VSUBS 0.006766f
C203 B.n85 VSUBS 0.006766f
C204 B.n86 VSUBS 0.006766f
C205 B.n87 VSUBS 0.006766f
C206 B.n88 VSUBS 0.006766f
C207 B.n89 VSUBS 0.006766f
C208 B.n90 VSUBS 0.006766f
C209 B.n91 VSUBS 0.006766f
C210 B.n92 VSUBS 0.006766f
C211 B.n93 VSUBS 0.006766f
C212 B.n94 VSUBS 0.017496f
C213 B.n95 VSUBS 0.006766f
C214 B.n96 VSUBS 0.006766f
C215 B.n97 VSUBS 0.006766f
C216 B.n98 VSUBS 0.006766f
C217 B.n99 VSUBS 0.006766f
C218 B.n100 VSUBS 0.006766f
C219 B.n101 VSUBS 0.006766f
C220 B.n102 VSUBS 0.006766f
C221 B.n103 VSUBS 0.006766f
C222 B.n104 VSUBS 0.006766f
C223 B.n105 VSUBS 0.006766f
C224 B.n106 VSUBS 0.006766f
C225 B.n107 VSUBS 0.006766f
C226 B.n108 VSUBS 0.006766f
C227 B.n109 VSUBS 0.006766f
C228 B.n110 VSUBS 0.006766f
C229 B.n111 VSUBS 0.006766f
C230 B.n112 VSUBS 0.006766f
C231 B.n113 VSUBS 0.006766f
C232 B.n114 VSUBS 0.006766f
C233 B.n115 VSUBS 0.006766f
C234 B.n116 VSUBS 0.006766f
C235 B.n117 VSUBS 0.006766f
C236 B.n118 VSUBS 0.006766f
C237 B.n119 VSUBS 0.006766f
C238 B.n120 VSUBS 0.006766f
C239 B.n121 VSUBS 0.006766f
C240 B.n122 VSUBS 0.006766f
C241 B.n123 VSUBS 0.006766f
C242 B.n124 VSUBS 0.006766f
C243 B.n125 VSUBS 0.006766f
C244 B.n126 VSUBS 0.006766f
C245 B.n127 VSUBS 0.006766f
C246 B.n128 VSUBS 0.006766f
C247 B.n129 VSUBS 0.006766f
C248 B.n130 VSUBS 0.006766f
C249 B.n131 VSUBS 0.006766f
C250 B.n132 VSUBS 0.006766f
C251 B.n133 VSUBS 0.006766f
C252 B.n134 VSUBS 0.006766f
C253 B.n135 VSUBS 0.006766f
C254 B.n136 VSUBS 0.006766f
C255 B.n137 VSUBS 0.006766f
C256 B.n138 VSUBS 0.006766f
C257 B.n139 VSUBS 0.006766f
C258 B.n140 VSUBS 0.006766f
C259 B.n141 VSUBS 0.006766f
C260 B.n142 VSUBS 0.006766f
C261 B.n143 VSUBS 0.006766f
C262 B.n144 VSUBS 0.006766f
C263 B.n145 VSUBS 0.006766f
C264 B.n146 VSUBS 0.006766f
C265 B.n147 VSUBS 0.016928f
C266 B.n148 VSUBS 0.006766f
C267 B.n149 VSUBS 0.006766f
C268 B.n150 VSUBS 0.006766f
C269 B.n151 VSUBS 0.006766f
C270 B.n152 VSUBS 0.006766f
C271 B.n153 VSUBS 0.006766f
C272 B.n154 VSUBS 0.006766f
C273 B.n155 VSUBS 0.006766f
C274 B.n156 VSUBS 0.006766f
C275 B.n157 VSUBS 0.006766f
C276 B.n158 VSUBS 0.006766f
C277 B.n159 VSUBS 0.006766f
C278 B.n160 VSUBS 0.006766f
C279 B.n161 VSUBS 0.006766f
C280 B.n162 VSUBS 0.006766f
C281 B.n163 VSUBS 0.006766f
C282 B.n164 VSUBS 0.006766f
C283 B.n165 VSUBS 0.006766f
C284 B.n166 VSUBS 0.006766f
C285 B.n167 VSUBS 0.006766f
C286 B.n168 VSUBS 0.006766f
C287 B.n169 VSUBS 0.006766f
C288 B.n170 VSUBS 0.006766f
C289 B.n171 VSUBS 0.006766f
C290 B.n172 VSUBS 0.006766f
C291 B.n173 VSUBS 0.006766f
C292 B.n174 VSUBS 0.006766f
C293 B.n175 VSUBS 0.006766f
C294 B.n176 VSUBS 0.004676f
C295 B.n177 VSUBS 0.006766f
C296 B.n178 VSUBS 0.006766f
C297 B.n179 VSUBS 0.006766f
C298 B.n180 VSUBS 0.006766f
C299 B.n181 VSUBS 0.006766f
C300 B.t11 VSUBS 0.329118f
C301 B.t10 VSUBS 0.362454f
C302 B.t9 VSUBS 2.04176f
C303 B.n182 VSUBS 0.558786f
C304 B.n183 VSUBS 0.312927f
C305 B.n184 VSUBS 0.006766f
C306 B.n185 VSUBS 0.006766f
C307 B.n186 VSUBS 0.006766f
C308 B.n187 VSUBS 0.006766f
C309 B.n188 VSUBS 0.006766f
C310 B.n189 VSUBS 0.006766f
C311 B.n190 VSUBS 0.006766f
C312 B.n191 VSUBS 0.006766f
C313 B.n192 VSUBS 0.006766f
C314 B.n193 VSUBS 0.006766f
C315 B.n194 VSUBS 0.006766f
C316 B.n195 VSUBS 0.006766f
C317 B.n196 VSUBS 0.006766f
C318 B.n197 VSUBS 0.006766f
C319 B.n198 VSUBS 0.006766f
C320 B.n199 VSUBS 0.006766f
C321 B.n200 VSUBS 0.006766f
C322 B.n201 VSUBS 0.006766f
C323 B.n202 VSUBS 0.006766f
C324 B.n203 VSUBS 0.006766f
C325 B.n204 VSUBS 0.006766f
C326 B.n205 VSUBS 0.006766f
C327 B.n206 VSUBS 0.006766f
C328 B.n207 VSUBS 0.006766f
C329 B.n208 VSUBS 0.006766f
C330 B.n209 VSUBS 0.006766f
C331 B.n210 VSUBS 0.006766f
C332 B.n211 VSUBS 0.006766f
C333 B.n212 VSUBS 0.016928f
C334 B.n213 VSUBS 0.006766f
C335 B.n214 VSUBS 0.006766f
C336 B.n215 VSUBS 0.006766f
C337 B.n216 VSUBS 0.006766f
C338 B.n217 VSUBS 0.006766f
C339 B.n218 VSUBS 0.006766f
C340 B.n219 VSUBS 0.006766f
C341 B.n220 VSUBS 0.006766f
C342 B.n221 VSUBS 0.006766f
C343 B.n222 VSUBS 0.006766f
C344 B.n223 VSUBS 0.006766f
C345 B.n224 VSUBS 0.006766f
C346 B.n225 VSUBS 0.006766f
C347 B.n226 VSUBS 0.006766f
C348 B.n227 VSUBS 0.006766f
C349 B.n228 VSUBS 0.006766f
C350 B.n229 VSUBS 0.006766f
C351 B.n230 VSUBS 0.006766f
C352 B.n231 VSUBS 0.006766f
C353 B.n232 VSUBS 0.006766f
C354 B.n233 VSUBS 0.006766f
C355 B.n234 VSUBS 0.006766f
C356 B.n235 VSUBS 0.006766f
C357 B.n236 VSUBS 0.006766f
C358 B.n237 VSUBS 0.006766f
C359 B.n238 VSUBS 0.006766f
C360 B.n239 VSUBS 0.006766f
C361 B.n240 VSUBS 0.006766f
C362 B.n241 VSUBS 0.006766f
C363 B.n242 VSUBS 0.006766f
C364 B.n243 VSUBS 0.006766f
C365 B.n244 VSUBS 0.006766f
C366 B.n245 VSUBS 0.006766f
C367 B.n246 VSUBS 0.006766f
C368 B.n247 VSUBS 0.006766f
C369 B.n248 VSUBS 0.006766f
C370 B.n249 VSUBS 0.006766f
C371 B.n250 VSUBS 0.006766f
C372 B.n251 VSUBS 0.006766f
C373 B.n252 VSUBS 0.006766f
C374 B.n253 VSUBS 0.006766f
C375 B.n254 VSUBS 0.006766f
C376 B.n255 VSUBS 0.006766f
C377 B.n256 VSUBS 0.006766f
C378 B.n257 VSUBS 0.006766f
C379 B.n258 VSUBS 0.006766f
C380 B.n259 VSUBS 0.006766f
C381 B.n260 VSUBS 0.006766f
C382 B.n261 VSUBS 0.006766f
C383 B.n262 VSUBS 0.006766f
C384 B.n263 VSUBS 0.006766f
C385 B.n264 VSUBS 0.006766f
C386 B.n265 VSUBS 0.006766f
C387 B.n266 VSUBS 0.006766f
C388 B.n267 VSUBS 0.006766f
C389 B.n268 VSUBS 0.006766f
C390 B.n269 VSUBS 0.006766f
C391 B.n270 VSUBS 0.006766f
C392 B.n271 VSUBS 0.006766f
C393 B.n272 VSUBS 0.006766f
C394 B.n273 VSUBS 0.006766f
C395 B.n274 VSUBS 0.006766f
C396 B.n275 VSUBS 0.006766f
C397 B.n276 VSUBS 0.006766f
C398 B.n277 VSUBS 0.006766f
C399 B.n278 VSUBS 0.006766f
C400 B.n279 VSUBS 0.006766f
C401 B.n280 VSUBS 0.006766f
C402 B.n281 VSUBS 0.006766f
C403 B.n282 VSUBS 0.006766f
C404 B.n283 VSUBS 0.006766f
C405 B.n284 VSUBS 0.006766f
C406 B.n285 VSUBS 0.006766f
C407 B.n286 VSUBS 0.006766f
C408 B.n287 VSUBS 0.006766f
C409 B.n288 VSUBS 0.006766f
C410 B.n289 VSUBS 0.006766f
C411 B.n290 VSUBS 0.006766f
C412 B.n291 VSUBS 0.006766f
C413 B.n292 VSUBS 0.006766f
C414 B.n293 VSUBS 0.006766f
C415 B.n294 VSUBS 0.006766f
C416 B.n295 VSUBS 0.006766f
C417 B.n296 VSUBS 0.006766f
C418 B.n297 VSUBS 0.006766f
C419 B.n298 VSUBS 0.006766f
C420 B.n299 VSUBS 0.006766f
C421 B.n300 VSUBS 0.006766f
C422 B.n301 VSUBS 0.006766f
C423 B.n302 VSUBS 0.006766f
C424 B.n303 VSUBS 0.006766f
C425 B.n304 VSUBS 0.006766f
C426 B.n305 VSUBS 0.006766f
C427 B.n306 VSUBS 0.006766f
C428 B.n307 VSUBS 0.006766f
C429 B.n308 VSUBS 0.006766f
C430 B.n309 VSUBS 0.006766f
C431 B.n310 VSUBS 0.006766f
C432 B.n311 VSUBS 0.006766f
C433 B.n312 VSUBS 0.006766f
C434 B.n313 VSUBS 0.016928f
C435 B.n314 VSUBS 0.017496f
C436 B.n315 VSUBS 0.017496f
C437 B.n316 VSUBS 0.006766f
C438 B.n317 VSUBS 0.006766f
C439 B.n318 VSUBS 0.006766f
C440 B.n319 VSUBS 0.006766f
C441 B.n320 VSUBS 0.006766f
C442 B.n321 VSUBS 0.006766f
C443 B.n322 VSUBS 0.006766f
C444 B.n323 VSUBS 0.006766f
C445 B.n324 VSUBS 0.006766f
C446 B.n325 VSUBS 0.006766f
C447 B.n326 VSUBS 0.006766f
C448 B.n327 VSUBS 0.006766f
C449 B.n328 VSUBS 0.006766f
C450 B.n329 VSUBS 0.006766f
C451 B.n330 VSUBS 0.006766f
C452 B.n331 VSUBS 0.006766f
C453 B.n332 VSUBS 0.006766f
C454 B.n333 VSUBS 0.006766f
C455 B.n334 VSUBS 0.006766f
C456 B.n335 VSUBS 0.006766f
C457 B.n336 VSUBS 0.006766f
C458 B.n337 VSUBS 0.006766f
C459 B.n338 VSUBS 0.006766f
C460 B.n339 VSUBS 0.006766f
C461 B.n340 VSUBS 0.006766f
C462 B.n341 VSUBS 0.006766f
C463 B.n342 VSUBS 0.006766f
C464 B.n343 VSUBS 0.006766f
C465 B.n344 VSUBS 0.006766f
C466 B.n345 VSUBS 0.006766f
C467 B.n346 VSUBS 0.006766f
C468 B.n347 VSUBS 0.006766f
C469 B.n348 VSUBS 0.006766f
C470 B.n349 VSUBS 0.006766f
C471 B.n350 VSUBS 0.006766f
C472 B.n351 VSUBS 0.006766f
C473 B.n352 VSUBS 0.006766f
C474 B.n353 VSUBS 0.006766f
C475 B.n354 VSUBS 0.006766f
C476 B.n355 VSUBS 0.006766f
C477 B.n356 VSUBS 0.006766f
C478 B.n357 VSUBS 0.006766f
C479 B.n358 VSUBS 0.006766f
C480 B.n359 VSUBS 0.006766f
C481 B.n360 VSUBS 0.006766f
C482 B.n361 VSUBS 0.006766f
C483 B.n362 VSUBS 0.006766f
C484 B.n363 VSUBS 0.006766f
C485 B.n364 VSUBS 0.006766f
C486 B.n365 VSUBS 0.006766f
C487 B.n366 VSUBS 0.006766f
C488 B.n367 VSUBS 0.006766f
C489 B.n368 VSUBS 0.006766f
C490 B.n369 VSUBS 0.006766f
C491 B.n370 VSUBS 0.006766f
C492 B.n371 VSUBS 0.006766f
C493 B.n372 VSUBS 0.006766f
C494 B.n373 VSUBS 0.006766f
C495 B.n374 VSUBS 0.006766f
C496 B.n375 VSUBS 0.006766f
C497 B.n376 VSUBS 0.006766f
C498 B.n377 VSUBS 0.006766f
C499 B.n378 VSUBS 0.006766f
C500 B.n379 VSUBS 0.006766f
C501 B.n380 VSUBS 0.006766f
C502 B.n381 VSUBS 0.006766f
C503 B.n382 VSUBS 0.006766f
C504 B.n383 VSUBS 0.006766f
C505 B.n384 VSUBS 0.006766f
C506 B.n385 VSUBS 0.006766f
C507 B.n386 VSUBS 0.006766f
C508 B.n387 VSUBS 0.006766f
C509 B.n388 VSUBS 0.006766f
C510 B.n389 VSUBS 0.006766f
C511 B.n390 VSUBS 0.006766f
C512 B.n391 VSUBS 0.006766f
C513 B.n392 VSUBS 0.006766f
C514 B.n393 VSUBS 0.006766f
C515 B.n394 VSUBS 0.006766f
C516 B.n395 VSUBS 0.006766f
C517 B.n396 VSUBS 0.006766f
C518 B.n397 VSUBS 0.006766f
C519 B.n398 VSUBS 0.006766f
C520 B.n399 VSUBS 0.006766f
C521 B.n400 VSUBS 0.004676f
C522 B.n401 VSUBS 0.015675f
C523 B.n402 VSUBS 0.005472f
C524 B.n403 VSUBS 0.006766f
C525 B.n404 VSUBS 0.006766f
C526 B.n405 VSUBS 0.006766f
C527 B.n406 VSUBS 0.006766f
C528 B.n407 VSUBS 0.006766f
C529 B.n408 VSUBS 0.006766f
C530 B.n409 VSUBS 0.006766f
C531 B.n410 VSUBS 0.006766f
C532 B.n411 VSUBS 0.006766f
C533 B.n412 VSUBS 0.006766f
C534 B.n413 VSUBS 0.006766f
C535 B.t5 VSUBS 0.329121f
C536 B.t4 VSUBS 0.362457f
C537 B.t3 VSUBS 2.04176f
C538 B.n414 VSUBS 0.558783f
C539 B.n415 VSUBS 0.312923f
C540 B.n416 VSUBS 0.015675f
C541 B.n417 VSUBS 0.005472f
C542 B.n418 VSUBS 0.006766f
C543 B.n419 VSUBS 0.006766f
C544 B.n420 VSUBS 0.006766f
C545 B.n421 VSUBS 0.006766f
C546 B.n422 VSUBS 0.006766f
C547 B.n423 VSUBS 0.006766f
C548 B.n424 VSUBS 0.006766f
C549 B.n425 VSUBS 0.006766f
C550 B.n426 VSUBS 0.006766f
C551 B.n427 VSUBS 0.006766f
C552 B.n428 VSUBS 0.006766f
C553 B.n429 VSUBS 0.006766f
C554 B.n430 VSUBS 0.006766f
C555 B.n431 VSUBS 0.006766f
C556 B.n432 VSUBS 0.006766f
C557 B.n433 VSUBS 0.006766f
C558 B.n434 VSUBS 0.006766f
C559 B.n435 VSUBS 0.006766f
C560 B.n436 VSUBS 0.006766f
C561 B.n437 VSUBS 0.006766f
C562 B.n438 VSUBS 0.006766f
C563 B.n439 VSUBS 0.006766f
C564 B.n440 VSUBS 0.006766f
C565 B.n441 VSUBS 0.006766f
C566 B.n442 VSUBS 0.006766f
C567 B.n443 VSUBS 0.006766f
C568 B.n444 VSUBS 0.006766f
C569 B.n445 VSUBS 0.006766f
C570 B.n446 VSUBS 0.006766f
C571 B.n447 VSUBS 0.006766f
C572 B.n448 VSUBS 0.006766f
C573 B.n449 VSUBS 0.006766f
C574 B.n450 VSUBS 0.006766f
C575 B.n451 VSUBS 0.006766f
C576 B.n452 VSUBS 0.006766f
C577 B.n453 VSUBS 0.006766f
C578 B.n454 VSUBS 0.006766f
C579 B.n455 VSUBS 0.006766f
C580 B.n456 VSUBS 0.006766f
C581 B.n457 VSUBS 0.006766f
C582 B.n458 VSUBS 0.006766f
C583 B.n459 VSUBS 0.006766f
C584 B.n460 VSUBS 0.006766f
C585 B.n461 VSUBS 0.006766f
C586 B.n462 VSUBS 0.006766f
C587 B.n463 VSUBS 0.006766f
C588 B.n464 VSUBS 0.006766f
C589 B.n465 VSUBS 0.006766f
C590 B.n466 VSUBS 0.006766f
C591 B.n467 VSUBS 0.006766f
C592 B.n468 VSUBS 0.006766f
C593 B.n469 VSUBS 0.006766f
C594 B.n470 VSUBS 0.006766f
C595 B.n471 VSUBS 0.006766f
C596 B.n472 VSUBS 0.006766f
C597 B.n473 VSUBS 0.006766f
C598 B.n474 VSUBS 0.006766f
C599 B.n475 VSUBS 0.006766f
C600 B.n476 VSUBS 0.006766f
C601 B.n477 VSUBS 0.006766f
C602 B.n478 VSUBS 0.006766f
C603 B.n479 VSUBS 0.006766f
C604 B.n480 VSUBS 0.006766f
C605 B.n481 VSUBS 0.006766f
C606 B.n482 VSUBS 0.006766f
C607 B.n483 VSUBS 0.006766f
C608 B.n484 VSUBS 0.006766f
C609 B.n485 VSUBS 0.006766f
C610 B.n486 VSUBS 0.006766f
C611 B.n487 VSUBS 0.006766f
C612 B.n488 VSUBS 0.006766f
C613 B.n489 VSUBS 0.006766f
C614 B.n490 VSUBS 0.006766f
C615 B.n491 VSUBS 0.006766f
C616 B.n492 VSUBS 0.006766f
C617 B.n493 VSUBS 0.006766f
C618 B.n494 VSUBS 0.006766f
C619 B.n495 VSUBS 0.006766f
C620 B.n496 VSUBS 0.006766f
C621 B.n497 VSUBS 0.006766f
C622 B.n498 VSUBS 0.006766f
C623 B.n499 VSUBS 0.006766f
C624 B.n500 VSUBS 0.006766f
C625 B.n501 VSUBS 0.006766f
C626 B.n502 VSUBS 0.006766f
C627 B.n503 VSUBS 0.006766f
C628 B.n504 VSUBS 0.017496f
C629 B.n505 VSUBS 0.016791f
C630 B.n506 VSUBS 0.017634f
C631 B.n507 VSUBS 0.006766f
C632 B.n508 VSUBS 0.006766f
C633 B.n509 VSUBS 0.006766f
C634 B.n510 VSUBS 0.006766f
C635 B.n511 VSUBS 0.006766f
C636 B.n512 VSUBS 0.006766f
C637 B.n513 VSUBS 0.006766f
C638 B.n514 VSUBS 0.006766f
C639 B.n515 VSUBS 0.006766f
C640 B.n516 VSUBS 0.006766f
C641 B.n517 VSUBS 0.006766f
C642 B.n518 VSUBS 0.006766f
C643 B.n519 VSUBS 0.006766f
C644 B.n520 VSUBS 0.006766f
C645 B.n521 VSUBS 0.006766f
C646 B.n522 VSUBS 0.006766f
C647 B.n523 VSUBS 0.006766f
C648 B.n524 VSUBS 0.006766f
C649 B.n525 VSUBS 0.006766f
C650 B.n526 VSUBS 0.006766f
C651 B.n527 VSUBS 0.006766f
C652 B.n528 VSUBS 0.006766f
C653 B.n529 VSUBS 0.006766f
C654 B.n530 VSUBS 0.006766f
C655 B.n531 VSUBS 0.006766f
C656 B.n532 VSUBS 0.006766f
C657 B.n533 VSUBS 0.006766f
C658 B.n534 VSUBS 0.006766f
C659 B.n535 VSUBS 0.006766f
C660 B.n536 VSUBS 0.006766f
C661 B.n537 VSUBS 0.006766f
C662 B.n538 VSUBS 0.006766f
C663 B.n539 VSUBS 0.006766f
C664 B.n540 VSUBS 0.006766f
C665 B.n541 VSUBS 0.006766f
C666 B.n542 VSUBS 0.006766f
C667 B.n543 VSUBS 0.006766f
C668 B.n544 VSUBS 0.006766f
C669 B.n545 VSUBS 0.006766f
C670 B.n546 VSUBS 0.006766f
C671 B.n547 VSUBS 0.006766f
C672 B.n548 VSUBS 0.006766f
C673 B.n549 VSUBS 0.006766f
C674 B.n550 VSUBS 0.006766f
C675 B.n551 VSUBS 0.006766f
C676 B.n552 VSUBS 0.006766f
C677 B.n553 VSUBS 0.006766f
C678 B.n554 VSUBS 0.006766f
C679 B.n555 VSUBS 0.006766f
C680 B.n556 VSUBS 0.006766f
C681 B.n557 VSUBS 0.006766f
C682 B.n558 VSUBS 0.006766f
C683 B.n559 VSUBS 0.006766f
C684 B.n560 VSUBS 0.006766f
C685 B.n561 VSUBS 0.006766f
C686 B.n562 VSUBS 0.006766f
C687 B.n563 VSUBS 0.006766f
C688 B.n564 VSUBS 0.006766f
C689 B.n565 VSUBS 0.006766f
C690 B.n566 VSUBS 0.006766f
C691 B.n567 VSUBS 0.006766f
C692 B.n568 VSUBS 0.006766f
C693 B.n569 VSUBS 0.006766f
C694 B.n570 VSUBS 0.006766f
C695 B.n571 VSUBS 0.006766f
C696 B.n572 VSUBS 0.006766f
C697 B.n573 VSUBS 0.006766f
C698 B.n574 VSUBS 0.006766f
C699 B.n575 VSUBS 0.006766f
C700 B.n576 VSUBS 0.006766f
C701 B.n577 VSUBS 0.006766f
C702 B.n578 VSUBS 0.006766f
C703 B.n579 VSUBS 0.006766f
C704 B.n580 VSUBS 0.006766f
C705 B.n581 VSUBS 0.006766f
C706 B.n582 VSUBS 0.006766f
C707 B.n583 VSUBS 0.006766f
C708 B.n584 VSUBS 0.006766f
C709 B.n585 VSUBS 0.006766f
C710 B.n586 VSUBS 0.006766f
C711 B.n587 VSUBS 0.006766f
C712 B.n588 VSUBS 0.006766f
C713 B.n589 VSUBS 0.006766f
C714 B.n590 VSUBS 0.006766f
C715 B.n591 VSUBS 0.006766f
C716 B.n592 VSUBS 0.006766f
C717 B.n593 VSUBS 0.006766f
C718 B.n594 VSUBS 0.006766f
C719 B.n595 VSUBS 0.006766f
C720 B.n596 VSUBS 0.006766f
C721 B.n597 VSUBS 0.006766f
C722 B.n598 VSUBS 0.006766f
C723 B.n599 VSUBS 0.006766f
C724 B.n600 VSUBS 0.006766f
C725 B.n601 VSUBS 0.006766f
C726 B.n602 VSUBS 0.006766f
C727 B.n603 VSUBS 0.006766f
C728 B.n604 VSUBS 0.006766f
C729 B.n605 VSUBS 0.006766f
C730 B.n606 VSUBS 0.006766f
C731 B.n607 VSUBS 0.006766f
C732 B.n608 VSUBS 0.006766f
C733 B.n609 VSUBS 0.006766f
C734 B.n610 VSUBS 0.006766f
C735 B.n611 VSUBS 0.006766f
C736 B.n612 VSUBS 0.006766f
C737 B.n613 VSUBS 0.006766f
C738 B.n614 VSUBS 0.006766f
C739 B.n615 VSUBS 0.006766f
C740 B.n616 VSUBS 0.006766f
C741 B.n617 VSUBS 0.006766f
C742 B.n618 VSUBS 0.006766f
C743 B.n619 VSUBS 0.006766f
C744 B.n620 VSUBS 0.006766f
C745 B.n621 VSUBS 0.006766f
C746 B.n622 VSUBS 0.006766f
C747 B.n623 VSUBS 0.006766f
C748 B.n624 VSUBS 0.006766f
C749 B.n625 VSUBS 0.006766f
C750 B.n626 VSUBS 0.006766f
C751 B.n627 VSUBS 0.006766f
C752 B.n628 VSUBS 0.006766f
C753 B.n629 VSUBS 0.006766f
C754 B.n630 VSUBS 0.006766f
C755 B.n631 VSUBS 0.006766f
C756 B.n632 VSUBS 0.006766f
C757 B.n633 VSUBS 0.006766f
C758 B.n634 VSUBS 0.006766f
C759 B.n635 VSUBS 0.006766f
C760 B.n636 VSUBS 0.006766f
C761 B.n637 VSUBS 0.006766f
C762 B.n638 VSUBS 0.006766f
C763 B.n639 VSUBS 0.006766f
C764 B.n640 VSUBS 0.006766f
C765 B.n641 VSUBS 0.006766f
C766 B.n642 VSUBS 0.006766f
C767 B.n643 VSUBS 0.006766f
C768 B.n644 VSUBS 0.006766f
C769 B.n645 VSUBS 0.006766f
C770 B.n646 VSUBS 0.006766f
C771 B.n647 VSUBS 0.006766f
C772 B.n648 VSUBS 0.006766f
C773 B.n649 VSUBS 0.006766f
C774 B.n650 VSUBS 0.006766f
C775 B.n651 VSUBS 0.006766f
C776 B.n652 VSUBS 0.006766f
C777 B.n653 VSUBS 0.006766f
C778 B.n654 VSUBS 0.006766f
C779 B.n655 VSUBS 0.006766f
C780 B.n656 VSUBS 0.006766f
C781 B.n657 VSUBS 0.006766f
C782 B.n658 VSUBS 0.006766f
C783 B.n659 VSUBS 0.006766f
C784 B.n660 VSUBS 0.006766f
C785 B.n661 VSUBS 0.006766f
C786 B.n662 VSUBS 0.006766f
C787 B.n663 VSUBS 0.016928f
C788 B.n664 VSUBS 0.016928f
C789 B.n665 VSUBS 0.017496f
C790 B.n666 VSUBS 0.006766f
C791 B.n667 VSUBS 0.006766f
C792 B.n668 VSUBS 0.006766f
C793 B.n669 VSUBS 0.006766f
C794 B.n670 VSUBS 0.006766f
C795 B.n671 VSUBS 0.006766f
C796 B.n672 VSUBS 0.006766f
C797 B.n673 VSUBS 0.006766f
C798 B.n674 VSUBS 0.006766f
C799 B.n675 VSUBS 0.006766f
C800 B.n676 VSUBS 0.006766f
C801 B.n677 VSUBS 0.006766f
C802 B.n678 VSUBS 0.006766f
C803 B.n679 VSUBS 0.006766f
C804 B.n680 VSUBS 0.006766f
C805 B.n681 VSUBS 0.006766f
C806 B.n682 VSUBS 0.006766f
C807 B.n683 VSUBS 0.006766f
C808 B.n684 VSUBS 0.006766f
C809 B.n685 VSUBS 0.006766f
C810 B.n686 VSUBS 0.006766f
C811 B.n687 VSUBS 0.006766f
C812 B.n688 VSUBS 0.006766f
C813 B.n689 VSUBS 0.006766f
C814 B.n690 VSUBS 0.006766f
C815 B.n691 VSUBS 0.006766f
C816 B.n692 VSUBS 0.006766f
C817 B.n693 VSUBS 0.006766f
C818 B.n694 VSUBS 0.006766f
C819 B.n695 VSUBS 0.006766f
C820 B.n696 VSUBS 0.006766f
C821 B.n697 VSUBS 0.006766f
C822 B.n698 VSUBS 0.006766f
C823 B.n699 VSUBS 0.006766f
C824 B.n700 VSUBS 0.006766f
C825 B.n701 VSUBS 0.006766f
C826 B.n702 VSUBS 0.006766f
C827 B.n703 VSUBS 0.006766f
C828 B.n704 VSUBS 0.006766f
C829 B.n705 VSUBS 0.006766f
C830 B.n706 VSUBS 0.006766f
C831 B.n707 VSUBS 0.006766f
C832 B.n708 VSUBS 0.006766f
C833 B.n709 VSUBS 0.006766f
C834 B.n710 VSUBS 0.006766f
C835 B.n711 VSUBS 0.006766f
C836 B.n712 VSUBS 0.006766f
C837 B.n713 VSUBS 0.006766f
C838 B.n714 VSUBS 0.006766f
C839 B.n715 VSUBS 0.006766f
C840 B.n716 VSUBS 0.006766f
C841 B.n717 VSUBS 0.006766f
C842 B.n718 VSUBS 0.006766f
C843 B.n719 VSUBS 0.006766f
C844 B.n720 VSUBS 0.006766f
C845 B.n721 VSUBS 0.006766f
C846 B.n722 VSUBS 0.006766f
C847 B.n723 VSUBS 0.006766f
C848 B.n724 VSUBS 0.006766f
C849 B.n725 VSUBS 0.006766f
C850 B.n726 VSUBS 0.006766f
C851 B.n727 VSUBS 0.006766f
C852 B.n728 VSUBS 0.006766f
C853 B.n729 VSUBS 0.006766f
C854 B.n730 VSUBS 0.006766f
C855 B.n731 VSUBS 0.006766f
C856 B.n732 VSUBS 0.006766f
C857 B.n733 VSUBS 0.006766f
C858 B.n734 VSUBS 0.006766f
C859 B.n735 VSUBS 0.006766f
C860 B.n736 VSUBS 0.006766f
C861 B.n737 VSUBS 0.006766f
C862 B.n738 VSUBS 0.006766f
C863 B.n739 VSUBS 0.006766f
C864 B.n740 VSUBS 0.006766f
C865 B.n741 VSUBS 0.006766f
C866 B.n742 VSUBS 0.006766f
C867 B.n743 VSUBS 0.006766f
C868 B.n744 VSUBS 0.006766f
C869 B.n745 VSUBS 0.006766f
C870 B.n746 VSUBS 0.006766f
C871 B.n747 VSUBS 0.006766f
C872 B.n748 VSUBS 0.006766f
C873 B.n749 VSUBS 0.006766f
C874 B.n750 VSUBS 0.006766f
C875 B.n751 VSUBS 0.004676f
C876 B.n752 VSUBS 0.015675f
C877 B.n753 VSUBS 0.005472f
C878 B.n754 VSUBS 0.006766f
C879 B.n755 VSUBS 0.006766f
C880 B.n756 VSUBS 0.006766f
C881 B.n757 VSUBS 0.006766f
C882 B.n758 VSUBS 0.006766f
C883 B.n759 VSUBS 0.006766f
C884 B.n760 VSUBS 0.006766f
C885 B.n761 VSUBS 0.006766f
C886 B.n762 VSUBS 0.006766f
C887 B.n763 VSUBS 0.006766f
C888 B.n764 VSUBS 0.006766f
C889 B.n765 VSUBS 0.005472f
C890 B.n766 VSUBS 0.015675f
C891 B.n767 VSUBS 0.004676f
C892 B.n768 VSUBS 0.006766f
C893 B.n769 VSUBS 0.006766f
C894 B.n770 VSUBS 0.006766f
C895 B.n771 VSUBS 0.006766f
C896 B.n772 VSUBS 0.006766f
C897 B.n773 VSUBS 0.006766f
C898 B.n774 VSUBS 0.006766f
C899 B.n775 VSUBS 0.006766f
C900 B.n776 VSUBS 0.006766f
C901 B.n777 VSUBS 0.006766f
C902 B.n778 VSUBS 0.006766f
C903 B.n779 VSUBS 0.006766f
C904 B.n780 VSUBS 0.006766f
C905 B.n781 VSUBS 0.006766f
C906 B.n782 VSUBS 0.006766f
C907 B.n783 VSUBS 0.006766f
C908 B.n784 VSUBS 0.006766f
C909 B.n785 VSUBS 0.006766f
C910 B.n786 VSUBS 0.006766f
C911 B.n787 VSUBS 0.006766f
C912 B.n788 VSUBS 0.006766f
C913 B.n789 VSUBS 0.006766f
C914 B.n790 VSUBS 0.006766f
C915 B.n791 VSUBS 0.006766f
C916 B.n792 VSUBS 0.006766f
C917 B.n793 VSUBS 0.006766f
C918 B.n794 VSUBS 0.006766f
C919 B.n795 VSUBS 0.006766f
C920 B.n796 VSUBS 0.006766f
C921 B.n797 VSUBS 0.006766f
C922 B.n798 VSUBS 0.006766f
C923 B.n799 VSUBS 0.006766f
C924 B.n800 VSUBS 0.006766f
C925 B.n801 VSUBS 0.006766f
C926 B.n802 VSUBS 0.006766f
C927 B.n803 VSUBS 0.006766f
C928 B.n804 VSUBS 0.006766f
C929 B.n805 VSUBS 0.006766f
C930 B.n806 VSUBS 0.006766f
C931 B.n807 VSUBS 0.006766f
C932 B.n808 VSUBS 0.006766f
C933 B.n809 VSUBS 0.006766f
C934 B.n810 VSUBS 0.006766f
C935 B.n811 VSUBS 0.006766f
C936 B.n812 VSUBS 0.006766f
C937 B.n813 VSUBS 0.006766f
C938 B.n814 VSUBS 0.006766f
C939 B.n815 VSUBS 0.006766f
C940 B.n816 VSUBS 0.006766f
C941 B.n817 VSUBS 0.006766f
C942 B.n818 VSUBS 0.006766f
C943 B.n819 VSUBS 0.006766f
C944 B.n820 VSUBS 0.006766f
C945 B.n821 VSUBS 0.006766f
C946 B.n822 VSUBS 0.006766f
C947 B.n823 VSUBS 0.006766f
C948 B.n824 VSUBS 0.006766f
C949 B.n825 VSUBS 0.006766f
C950 B.n826 VSUBS 0.006766f
C951 B.n827 VSUBS 0.006766f
C952 B.n828 VSUBS 0.006766f
C953 B.n829 VSUBS 0.006766f
C954 B.n830 VSUBS 0.006766f
C955 B.n831 VSUBS 0.006766f
C956 B.n832 VSUBS 0.006766f
C957 B.n833 VSUBS 0.006766f
C958 B.n834 VSUBS 0.006766f
C959 B.n835 VSUBS 0.006766f
C960 B.n836 VSUBS 0.006766f
C961 B.n837 VSUBS 0.006766f
C962 B.n838 VSUBS 0.006766f
C963 B.n839 VSUBS 0.006766f
C964 B.n840 VSUBS 0.006766f
C965 B.n841 VSUBS 0.006766f
C966 B.n842 VSUBS 0.006766f
C967 B.n843 VSUBS 0.006766f
C968 B.n844 VSUBS 0.006766f
C969 B.n845 VSUBS 0.006766f
C970 B.n846 VSUBS 0.006766f
C971 B.n847 VSUBS 0.006766f
C972 B.n848 VSUBS 0.006766f
C973 B.n849 VSUBS 0.006766f
C974 B.n850 VSUBS 0.006766f
C975 B.n851 VSUBS 0.006766f
C976 B.n852 VSUBS 0.006766f
C977 B.n853 VSUBS 0.017496f
C978 B.n854 VSUBS 0.016928f
C979 B.n855 VSUBS 0.016928f
C980 B.n856 VSUBS 0.006766f
C981 B.n857 VSUBS 0.006766f
C982 B.n858 VSUBS 0.006766f
C983 B.n859 VSUBS 0.006766f
C984 B.n860 VSUBS 0.006766f
C985 B.n861 VSUBS 0.006766f
C986 B.n862 VSUBS 0.006766f
C987 B.n863 VSUBS 0.006766f
C988 B.n864 VSUBS 0.006766f
C989 B.n865 VSUBS 0.006766f
C990 B.n866 VSUBS 0.006766f
C991 B.n867 VSUBS 0.006766f
C992 B.n868 VSUBS 0.006766f
C993 B.n869 VSUBS 0.006766f
C994 B.n870 VSUBS 0.006766f
C995 B.n871 VSUBS 0.006766f
C996 B.n872 VSUBS 0.006766f
C997 B.n873 VSUBS 0.006766f
C998 B.n874 VSUBS 0.006766f
C999 B.n875 VSUBS 0.006766f
C1000 B.n876 VSUBS 0.006766f
C1001 B.n877 VSUBS 0.006766f
C1002 B.n878 VSUBS 0.006766f
C1003 B.n879 VSUBS 0.006766f
C1004 B.n880 VSUBS 0.006766f
C1005 B.n881 VSUBS 0.006766f
C1006 B.n882 VSUBS 0.006766f
C1007 B.n883 VSUBS 0.006766f
C1008 B.n884 VSUBS 0.006766f
C1009 B.n885 VSUBS 0.006766f
C1010 B.n886 VSUBS 0.006766f
C1011 B.n887 VSUBS 0.006766f
C1012 B.n888 VSUBS 0.006766f
C1013 B.n889 VSUBS 0.006766f
C1014 B.n890 VSUBS 0.006766f
C1015 B.n891 VSUBS 0.006766f
C1016 B.n892 VSUBS 0.006766f
C1017 B.n893 VSUBS 0.006766f
C1018 B.n894 VSUBS 0.006766f
C1019 B.n895 VSUBS 0.006766f
C1020 B.n896 VSUBS 0.006766f
C1021 B.n897 VSUBS 0.006766f
C1022 B.n898 VSUBS 0.006766f
C1023 B.n899 VSUBS 0.006766f
C1024 B.n900 VSUBS 0.006766f
C1025 B.n901 VSUBS 0.006766f
C1026 B.n902 VSUBS 0.006766f
C1027 B.n903 VSUBS 0.006766f
C1028 B.n904 VSUBS 0.006766f
C1029 B.n905 VSUBS 0.006766f
C1030 B.n906 VSUBS 0.006766f
C1031 B.n907 VSUBS 0.006766f
C1032 B.n908 VSUBS 0.006766f
C1033 B.n909 VSUBS 0.006766f
C1034 B.n910 VSUBS 0.006766f
C1035 B.n911 VSUBS 0.006766f
C1036 B.n912 VSUBS 0.006766f
C1037 B.n913 VSUBS 0.006766f
C1038 B.n914 VSUBS 0.006766f
C1039 B.n915 VSUBS 0.006766f
C1040 B.n916 VSUBS 0.006766f
C1041 B.n917 VSUBS 0.006766f
C1042 B.n918 VSUBS 0.006766f
C1043 B.n919 VSUBS 0.006766f
C1044 B.n920 VSUBS 0.006766f
C1045 B.n921 VSUBS 0.006766f
C1046 B.n922 VSUBS 0.006766f
C1047 B.n923 VSUBS 0.006766f
C1048 B.n924 VSUBS 0.006766f
C1049 B.n925 VSUBS 0.006766f
C1050 B.n926 VSUBS 0.006766f
C1051 B.n927 VSUBS 0.006766f
C1052 B.n928 VSUBS 0.006766f
C1053 B.n929 VSUBS 0.006766f
C1054 B.n930 VSUBS 0.006766f
C1055 B.n931 VSUBS 0.008829f
C1056 B.n932 VSUBS 0.009405f
C1057 B.n933 VSUBS 0.018702f
C1058 VDD1.t0 VSUBS 0.371373f
C1059 VDD1.t7 VSUBS 0.371373f
C1060 VDD1.n0 VSUBS 3.09555f
C1061 VDD1.t1 VSUBS 0.371373f
C1062 VDD1.t3 VSUBS 0.371373f
C1063 VDD1.n1 VSUBS 3.094f
C1064 VDD1.t6 VSUBS 0.371373f
C1065 VDD1.t2 VSUBS 0.371373f
C1066 VDD1.n2 VSUBS 3.094f
C1067 VDD1.n3 VSUBS 4.5999f
C1068 VDD1.t5 VSUBS 0.371373f
C1069 VDD1.t4 VSUBS 0.371373f
C1070 VDD1.n4 VSUBS 3.07873f
C1071 VDD1.n5 VSUBS 3.98168f
C1072 VTAIL.t6 VSUBS 0.329786f
C1073 VTAIL.t3 VSUBS 0.329786f
C1074 VTAIL.n0 VSUBS 2.58955f
C1075 VTAIL.n1 VSUBS 0.781071f
C1076 VTAIL.n2 VSUBS 0.026014f
C1077 VTAIL.n3 VSUBS 0.023766f
C1078 VTAIL.n4 VSUBS 0.012771f
C1079 VTAIL.n5 VSUBS 0.030185f
C1080 VTAIL.n6 VSUBS 0.013522f
C1081 VTAIL.n7 VSUBS 0.023766f
C1082 VTAIL.n8 VSUBS 0.012771f
C1083 VTAIL.n9 VSUBS 0.030185f
C1084 VTAIL.n10 VSUBS 0.013146f
C1085 VTAIL.n11 VSUBS 0.023766f
C1086 VTAIL.n12 VSUBS 0.013522f
C1087 VTAIL.n13 VSUBS 0.030185f
C1088 VTAIL.n14 VSUBS 0.013522f
C1089 VTAIL.n15 VSUBS 0.023766f
C1090 VTAIL.n16 VSUBS 0.012771f
C1091 VTAIL.n17 VSUBS 0.030185f
C1092 VTAIL.n18 VSUBS 0.013522f
C1093 VTAIL.n19 VSUBS 0.023766f
C1094 VTAIL.n20 VSUBS 0.012771f
C1095 VTAIL.n21 VSUBS 0.030185f
C1096 VTAIL.n22 VSUBS 0.013522f
C1097 VTAIL.n23 VSUBS 0.023766f
C1098 VTAIL.n24 VSUBS 0.012771f
C1099 VTAIL.n25 VSUBS 0.030185f
C1100 VTAIL.n26 VSUBS 0.013522f
C1101 VTAIL.n27 VSUBS 0.023766f
C1102 VTAIL.n28 VSUBS 0.012771f
C1103 VTAIL.n29 VSUBS 0.030185f
C1104 VTAIL.n30 VSUBS 0.013522f
C1105 VTAIL.n31 VSUBS 1.7937f
C1106 VTAIL.n32 VSUBS 0.012771f
C1107 VTAIL.t2 VSUBS 0.064772f
C1108 VTAIL.n33 VSUBS 0.185474f
C1109 VTAIL.n34 VSUBS 0.019203f
C1110 VTAIL.n35 VSUBS 0.022639f
C1111 VTAIL.n36 VSUBS 0.030185f
C1112 VTAIL.n37 VSUBS 0.013522f
C1113 VTAIL.n38 VSUBS 0.012771f
C1114 VTAIL.n39 VSUBS 0.023766f
C1115 VTAIL.n40 VSUBS 0.023766f
C1116 VTAIL.n41 VSUBS 0.012771f
C1117 VTAIL.n42 VSUBS 0.013522f
C1118 VTAIL.n43 VSUBS 0.030185f
C1119 VTAIL.n44 VSUBS 0.030185f
C1120 VTAIL.n45 VSUBS 0.013522f
C1121 VTAIL.n46 VSUBS 0.012771f
C1122 VTAIL.n47 VSUBS 0.023766f
C1123 VTAIL.n48 VSUBS 0.023766f
C1124 VTAIL.n49 VSUBS 0.012771f
C1125 VTAIL.n50 VSUBS 0.013522f
C1126 VTAIL.n51 VSUBS 0.030185f
C1127 VTAIL.n52 VSUBS 0.030185f
C1128 VTAIL.n53 VSUBS 0.013522f
C1129 VTAIL.n54 VSUBS 0.012771f
C1130 VTAIL.n55 VSUBS 0.023766f
C1131 VTAIL.n56 VSUBS 0.023766f
C1132 VTAIL.n57 VSUBS 0.012771f
C1133 VTAIL.n58 VSUBS 0.013522f
C1134 VTAIL.n59 VSUBS 0.030185f
C1135 VTAIL.n60 VSUBS 0.030185f
C1136 VTAIL.n61 VSUBS 0.013522f
C1137 VTAIL.n62 VSUBS 0.012771f
C1138 VTAIL.n63 VSUBS 0.023766f
C1139 VTAIL.n64 VSUBS 0.023766f
C1140 VTAIL.n65 VSUBS 0.012771f
C1141 VTAIL.n66 VSUBS 0.013522f
C1142 VTAIL.n67 VSUBS 0.030185f
C1143 VTAIL.n68 VSUBS 0.030185f
C1144 VTAIL.n69 VSUBS 0.013522f
C1145 VTAIL.n70 VSUBS 0.012771f
C1146 VTAIL.n71 VSUBS 0.023766f
C1147 VTAIL.n72 VSUBS 0.023766f
C1148 VTAIL.n73 VSUBS 0.012771f
C1149 VTAIL.n74 VSUBS 0.012771f
C1150 VTAIL.n75 VSUBS 0.013522f
C1151 VTAIL.n76 VSUBS 0.030185f
C1152 VTAIL.n77 VSUBS 0.030185f
C1153 VTAIL.n78 VSUBS 0.030185f
C1154 VTAIL.n79 VSUBS 0.013146f
C1155 VTAIL.n80 VSUBS 0.012771f
C1156 VTAIL.n81 VSUBS 0.023766f
C1157 VTAIL.n82 VSUBS 0.023766f
C1158 VTAIL.n83 VSUBS 0.012771f
C1159 VTAIL.n84 VSUBS 0.013522f
C1160 VTAIL.n85 VSUBS 0.030185f
C1161 VTAIL.n86 VSUBS 0.030185f
C1162 VTAIL.n87 VSUBS 0.013522f
C1163 VTAIL.n88 VSUBS 0.012771f
C1164 VTAIL.n89 VSUBS 0.023766f
C1165 VTAIL.n90 VSUBS 0.023766f
C1166 VTAIL.n91 VSUBS 0.012771f
C1167 VTAIL.n92 VSUBS 0.013522f
C1168 VTAIL.n93 VSUBS 0.030185f
C1169 VTAIL.n94 VSUBS 0.072737f
C1170 VTAIL.n95 VSUBS 0.013522f
C1171 VTAIL.n96 VSUBS 0.012771f
C1172 VTAIL.n97 VSUBS 0.056232f
C1173 VTAIL.n98 VSUBS 0.036603f
C1174 VTAIL.n99 VSUBS 0.257039f
C1175 VTAIL.n100 VSUBS 0.026014f
C1176 VTAIL.n101 VSUBS 0.023766f
C1177 VTAIL.n102 VSUBS 0.012771f
C1178 VTAIL.n103 VSUBS 0.030185f
C1179 VTAIL.n104 VSUBS 0.013522f
C1180 VTAIL.n105 VSUBS 0.023766f
C1181 VTAIL.n106 VSUBS 0.012771f
C1182 VTAIL.n107 VSUBS 0.030185f
C1183 VTAIL.n108 VSUBS 0.013146f
C1184 VTAIL.n109 VSUBS 0.023766f
C1185 VTAIL.n110 VSUBS 0.013522f
C1186 VTAIL.n111 VSUBS 0.030185f
C1187 VTAIL.n112 VSUBS 0.013522f
C1188 VTAIL.n113 VSUBS 0.023766f
C1189 VTAIL.n114 VSUBS 0.012771f
C1190 VTAIL.n115 VSUBS 0.030185f
C1191 VTAIL.n116 VSUBS 0.013522f
C1192 VTAIL.n117 VSUBS 0.023766f
C1193 VTAIL.n118 VSUBS 0.012771f
C1194 VTAIL.n119 VSUBS 0.030185f
C1195 VTAIL.n120 VSUBS 0.013522f
C1196 VTAIL.n121 VSUBS 0.023766f
C1197 VTAIL.n122 VSUBS 0.012771f
C1198 VTAIL.n123 VSUBS 0.030185f
C1199 VTAIL.n124 VSUBS 0.013522f
C1200 VTAIL.n125 VSUBS 0.023766f
C1201 VTAIL.n126 VSUBS 0.012771f
C1202 VTAIL.n127 VSUBS 0.030185f
C1203 VTAIL.n128 VSUBS 0.013522f
C1204 VTAIL.n129 VSUBS 1.7937f
C1205 VTAIL.n130 VSUBS 0.012771f
C1206 VTAIL.t13 VSUBS 0.064772f
C1207 VTAIL.n131 VSUBS 0.185474f
C1208 VTAIL.n132 VSUBS 0.019203f
C1209 VTAIL.n133 VSUBS 0.022639f
C1210 VTAIL.n134 VSUBS 0.030185f
C1211 VTAIL.n135 VSUBS 0.013522f
C1212 VTAIL.n136 VSUBS 0.012771f
C1213 VTAIL.n137 VSUBS 0.023766f
C1214 VTAIL.n138 VSUBS 0.023766f
C1215 VTAIL.n139 VSUBS 0.012771f
C1216 VTAIL.n140 VSUBS 0.013522f
C1217 VTAIL.n141 VSUBS 0.030185f
C1218 VTAIL.n142 VSUBS 0.030185f
C1219 VTAIL.n143 VSUBS 0.013522f
C1220 VTAIL.n144 VSUBS 0.012771f
C1221 VTAIL.n145 VSUBS 0.023766f
C1222 VTAIL.n146 VSUBS 0.023766f
C1223 VTAIL.n147 VSUBS 0.012771f
C1224 VTAIL.n148 VSUBS 0.013522f
C1225 VTAIL.n149 VSUBS 0.030185f
C1226 VTAIL.n150 VSUBS 0.030185f
C1227 VTAIL.n151 VSUBS 0.013522f
C1228 VTAIL.n152 VSUBS 0.012771f
C1229 VTAIL.n153 VSUBS 0.023766f
C1230 VTAIL.n154 VSUBS 0.023766f
C1231 VTAIL.n155 VSUBS 0.012771f
C1232 VTAIL.n156 VSUBS 0.013522f
C1233 VTAIL.n157 VSUBS 0.030185f
C1234 VTAIL.n158 VSUBS 0.030185f
C1235 VTAIL.n159 VSUBS 0.013522f
C1236 VTAIL.n160 VSUBS 0.012771f
C1237 VTAIL.n161 VSUBS 0.023766f
C1238 VTAIL.n162 VSUBS 0.023766f
C1239 VTAIL.n163 VSUBS 0.012771f
C1240 VTAIL.n164 VSUBS 0.013522f
C1241 VTAIL.n165 VSUBS 0.030185f
C1242 VTAIL.n166 VSUBS 0.030185f
C1243 VTAIL.n167 VSUBS 0.013522f
C1244 VTAIL.n168 VSUBS 0.012771f
C1245 VTAIL.n169 VSUBS 0.023766f
C1246 VTAIL.n170 VSUBS 0.023766f
C1247 VTAIL.n171 VSUBS 0.012771f
C1248 VTAIL.n172 VSUBS 0.012771f
C1249 VTAIL.n173 VSUBS 0.013522f
C1250 VTAIL.n174 VSUBS 0.030185f
C1251 VTAIL.n175 VSUBS 0.030185f
C1252 VTAIL.n176 VSUBS 0.030185f
C1253 VTAIL.n177 VSUBS 0.013146f
C1254 VTAIL.n178 VSUBS 0.012771f
C1255 VTAIL.n179 VSUBS 0.023766f
C1256 VTAIL.n180 VSUBS 0.023766f
C1257 VTAIL.n181 VSUBS 0.012771f
C1258 VTAIL.n182 VSUBS 0.013522f
C1259 VTAIL.n183 VSUBS 0.030185f
C1260 VTAIL.n184 VSUBS 0.030185f
C1261 VTAIL.n185 VSUBS 0.013522f
C1262 VTAIL.n186 VSUBS 0.012771f
C1263 VTAIL.n187 VSUBS 0.023766f
C1264 VTAIL.n188 VSUBS 0.023766f
C1265 VTAIL.n189 VSUBS 0.012771f
C1266 VTAIL.n190 VSUBS 0.013522f
C1267 VTAIL.n191 VSUBS 0.030185f
C1268 VTAIL.n192 VSUBS 0.072737f
C1269 VTAIL.n193 VSUBS 0.013522f
C1270 VTAIL.n194 VSUBS 0.012771f
C1271 VTAIL.n195 VSUBS 0.056232f
C1272 VTAIL.n196 VSUBS 0.036603f
C1273 VTAIL.n197 VSUBS 0.257039f
C1274 VTAIL.t14 VSUBS 0.329786f
C1275 VTAIL.t9 VSUBS 0.329786f
C1276 VTAIL.n198 VSUBS 2.58955f
C1277 VTAIL.n199 VSUBS 0.976644f
C1278 VTAIL.n200 VSUBS 0.026014f
C1279 VTAIL.n201 VSUBS 0.023766f
C1280 VTAIL.n202 VSUBS 0.012771f
C1281 VTAIL.n203 VSUBS 0.030185f
C1282 VTAIL.n204 VSUBS 0.013522f
C1283 VTAIL.n205 VSUBS 0.023766f
C1284 VTAIL.n206 VSUBS 0.012771f
C1285 VTAIL.n207 VSUBS 0.030185f
C1286 VTAIL.n208 VSUBS 0.013146f
C1287 VTAIL.n209 VSUBS 0.023766f
C1288 VTAIL.n210 VSUBS 0.013522f
C1289 VTAIL.n211 VSUBS 0.030185f
C1290 VTAIL.n212 VSUBS 0.013522f
C1291 VTAIL.n213 VSUBS 0.023766f
C1292 VTAIL.n214 VSUBS 0.012771f
C1293 VTAIL.n215 VSUBS 0.030185f
C1294 VTAIL.n216 VSUBS 0.013522f
C1295 VTAIL.n217 VSUBS 0.023766f
C1296 VTAIL.n218 VSUBS 0.012771f
C1297 VTAIL.n219 VSUBS 0.030185f
C1298 VTAIL.n220 VSUBS 0.013522f
C1299 VTAIL.n221 VSUBS 0.023766f
C1300 VTAIL.n222 VSUBS 0.012771f
C1301 VTAIL.n223 VSUBS 0.030185f
C1302 VTAIL.n224 VSUBS 0.013522f
C1303 VTAIL.n225 VSUBS 0.023766f
C1304 VTAIL.n226 VSUBS 0.012771f
C1305 VTAIL.n227 VSUBS 0.030185f
C1306 VTAIL.n228 VSUBS 0.013522f
C1307 VTAIL.n229 VSUBS 1.7937f
C1308 VTAIL.n230 VSUBS 0.012771f
C1309 VTAIL.t15 VSUBS 0.064772f
C1310 VTAIL.n231 VSUBS 0.185474f
C1311 VTAIL.n232 VSUBS 0.019203f
C1312 VTAIL.n233 VSUBS 0.022639f
C1313 VTAIL.n234 VSUBS 0.030185f
C1314 VTAIL.n235 VSUBS 0.013522f
C1315 VTAIL.n236 VSUBS 0.012771f
C1316 VTAIL.n237 VSUBS 0.023766f
C1317 VTAIL.n238 VSUBS 0.023766f
C1318 VTAIL.n239 VSUBS 0.012771f
C1319 VTAIL.n240 VSUBS 0.013522f
C1320 VTAIL.n241 VSUBS 0.030185f
C1321 VTAIL.n242 VSUBS 0.030185f
C1322 VTAIL.n243 VSUBS 0.013522f
C1323 VTAIL.n244 VSUBS 0.012771f
C1324 VTAIL.n245 VSUBS 0.023766f
C1325 VTAIL.n246 VSUBS 0.023766f
C1326 VTAIL.n247 VSUBS 0.012771f
C1327 VTAIL.n248 VSUBS 0.013522f
C1328 VTAIL.n249 VSUBS 0.030185f
C1329 VTAIL.n250 VSUBS 0.030185f
C1330 VTAIL.n251 VSUBS 0.013522f
C1331 VTAIL.n252 VSUBS 0.012771f
C1332 VTAIL.n253 VSUBS 0.023766f
C1333 VTAIL.n254 VSUBS 0.023766f
C1334 VTAIL.n255 VSUBS 0.012771f
C1335 VTAIL.n256 VSUBS 0.013522f
C1336 VTAIL.n257 VSUBS 0.030185f
C1337 VTAIL.n258 VSUBS 0.030185f
C1338 VTAIL.n259 VSUBS 0.013522f
C1339 VTAIL.n260 VSUBS 0.012771f
C1340 VTAIL.n261 VSUBS 0.023766f
C1341 VTAIL.n262 VSUBS 0.023766f
C1342 VTAIL.n263 VSUBS 0.012771f
C1343 VTAIL.n264 VSUBS 0.013522f
C1344 VTAIL.n265 VSUBS 0.030185f
C1345 VTAIL.n266 VSUBS 0.030185f
C1346 VTAIL.n267 VSUBS 0.013522f
C1347 VTAIL.n268 VSUBS 0.012771f
C1348 VTAIL.n269 VSUBS 0.023766f
C1349 VTAIL.n270 VSUBS 0.023766f
C1350 VTAIL.n271 VSUBS 0.012771f
C1351 VTAIL.n272 VSUBS 0.012771f
C1352 VTAIL.n273 VSUBS 0.013522f
C1353 VTAIL.n274 VSUBS 0.030185f
C1354 VTAIL.n275 VSUBS 0.030185f
C1355 VTAIL.n276 VSUBS 0.030185f
C1356 VTAIL.n277 VSUBS 0.013146f
C1357 VTAIL.n278 VSUBS 0.012771f
C1358 VTAIL.n279 VSUBS 0.023766f
C1359 VTAIL.n280 VSUBS 0.023766f
C1360 VTAIL.n281 VSUBS 0.012771f
C1361 VTAIL.n282 VSUBS 0.013522f
C1362 VTAIL.n283 VSUBS 0.030185f
C1363 VTAIL.n284 VSUBS 0.030185f
C1364 VTAIL.n285 VSUBS 0.013522f
C1365 VTAIL.n286 VSUBS 0.012771f
C1366 VTAIL.n287 VSUBS 0.023766f
C1367 VTAIL.n288 VSUBS 0.023766f
C1368 VTAIL.n289 VSUBS 0.012771f
C1369 VTAIL.n290 VSUBS 0.013522f
C1370 VTAIL.n291 VSUBS 0.030185f
C1371 VTAIL.n292 VSUBS 0.072737f
C1372 VTAIL.n293 VSUBS 0.013522f
C1373 VTAIL.n294 VSUBS 0.012771f
C1374 VTAIL.n295 VSUBS 0.056232f
C1375 VTAIL.n296 VSUBS 0.036603f
C1376 VTAIL.n297 VSUBS 1.90317f
C1377 VTAIL.n298 VSUBS 0.026014f
C1378 VTAIL.n299 VSUBS 0.023766f
C1379 VTAIL.n300 VSUBS 0.012771f
C1380 VTAIL.n301 VSUBS 0.030185f
C1381 VTAIL.n302 VSUBS 0.013522f
C1382 VTAIL.n303 VSUBS 0.023766f
C1383 VTAIL.n304 VSUBS 0.012771f
C1384 VTAIL.n305 VSUBS 0.030185f
C1385 VTAIL.n306 VSUBS 0.013146f
C1386 VTAIL.n307 VSUBS 0.023766f
C1387 VTAIL.n308 VSUBS 0.013146f
C1388 VTAIL.n309 VSUBS 0.012771f
C1389 VTAIL.n310 VSUBS 0.030185f
C1390 VTAIL.n311 VSUBS 0.030185f
C1391 VTAIL.n312 VSUBS 0.013522f
C1392 VTAIL.n313 VSUBS 0.023766f
C1393 VTAIL.n314 VSUBS 0.012771f
C1394 VTAIL.n315 VSUBS 0.030185f
C1395 VTAIL.n316 VSUBS 0.013522f
C1396 VTAIL.n317 VSUBS 0.023766f
C1397 VTAIL.n318 VSUBS 0.012771f
C1398 VTAIL.n319 VSUBS 0.030185f
C1399 VTAIL.n320 VSUBS 0.013522f
C1400 VTAIL.n321 VSUBS 0.023766f
C1401 VTAIL.n322 VSUBS 0.012771f
C1402 VTAIL.n323 VSUBS 0.030185f
C1403 VTAIL.n324 VSUBS 0.013522f
C1404 VTAIL.n325 VSUBS 0.023766f
C1405 VTAIL.n326 VSUBS 0.012771f
C1406 VTAIL.n327 VSUBS 0.030185f
C1407 VTAIL.n328 VSUBS 0.013522f
C1408 VTAIL.n329 VSUBS 1.7937f
C1409 VTAIL.n330 VSUBS 0.012771f
C1410 VTAIL.t5 VSUBS 0.064772f
C1411 VTAIL.n331 VSUBS 0.185474f
C1412 VTAIL.n332 VSUBS 0.019203f
C1413 VTAIL.n333 VSUBS 0.022639f
C1414 VTAIL.n334 VSUBS 0.030185f
C1415 VTAIL.n335 VSUBS 0.013522f
C1416 VTAIL.n336 VSUBS 0.012771f
C1417 VTAIL.n337 VSUBS 0.023766f
C1418 VTAIL.n338 VSUBS 0.023766f
C1419 VTAIL.n339 VSUBS 0.012771f
C1420 VTAIL.n340 VSUBS 0.013522f
C1421 VTAIL.n341 VSUBS 0.030185f
C1422 VTAIL.n342 VSUBS 0.030185f
C1423 VTAIL.n343 VSUBS 0.013522f
C1424 VTAIL.n344 VSUBS 0.012771f
C1425 VTAIL.n345 VSUBS 0.023766f
C1426 VTAIL.n346 VSUBS 0.023766f
C1427 VTAIL.n347 VSUBS 0.012771f
C1428 VTAIL.n348 VSUBS 0.013522f
C1429 VTAIL.n349 VSUBS 0.030185f
C1430 VTAIL.n350 VSUBS 0.030185f
C1431 VTAIL.n351 VSUBS 0.013522f
C1432 VTAIL.n352 VSUBS 0.012771f
C1433 VTAIL.n353 VSUBS 0.023766f
C1434 VTAIL.n354 VSUBS 0.023766f
C1435 VTAIL.n355 VSUBS 0.012771f
C1436 VTAIL.n356 VSUBS 0.013522f
C1437 VTAIL.n357 VSUBS 0.030185f
C1438 VTAIL.n358 VSUBS 0.030185f
C1439 VTAIL.n359 VSUBS 0.013522f
C1440 VTAIL.n360 VSUBS 0.012771f
C1441 VTAIL.n361 VSUBS 0.023766f
C1442 VTAIL.n362 VSUBS 0.023766f
C1443 VTAIL.n363 VSUBS 0.012771f
C1444 VTAIL.n364 VSUBS 0.013522f
C1445 VTAIL.n365 VSUBS 0.030185f
C1446 VTAIL.n366 VSUBS 0.030185f
C1447 VTAIL.n367 VSUBS 0.013522f
C1448 VTAIL.n368 VSUBS 0.012771f
C1449 VTAIL.n369 VSUBS 0.023766f
C1450 VTAIL.n370 VSUBS 0.023766f
C1451 VTAIL.n371 VSUBS 0.012771f
C1452 VTAIL.n372 VSUBS 0.013522f
C1453 VTAIL.n373 VSUBS 0.030185f
C1454 VTAIL.n374 VSUBS 0.030185f
C1455 VTAIL.n375 VSUBS 0.013522f
C1456 VTAIL.n376 VSUBS 0.012771f
C1457 VTAIL.n377 VSUBS 0.023766f
C1458 VTAIL.n378 VSUBS 0.023766f
C1459 VTAIL.n379 VSUBS 0.012771f
C1460 VTAIL.n380 VSUBS 0.013522f
C1461 VTAIL.n381 VSUBS 0.030185f
C1462 VTAIL.n382 VSUBS 0.030185f
C1463 VTAIL.n383 VSUBS 0.013522f
C1464 VTAIL.n384 VSUBS 0.012771f
C1465 VTAIL.n385 VSUBS 0.023766f
C1466 VTAIL.n386 VSUBS 0.023766f
C1467 VTAIL.n387 VSUBS 0.012771f
C1468 VTAIL.n388 VSUBS 0.013522f
C1469 VTAIL.n389 VSUBS 0.030185f
C1470 VTAIL.n390 VSUBS 0.072737f
C1471 VTAIL.n391 VSUBS 0.013522f
C1472 VTAIL.n392 VSUBS 0.012771f
C1473 VTAIL.n393 VSUBS 0.056232f
C1474 VTAIL.n394 VSUBS 0.036603f
C1475 VTAIL.n395 VSUBS 1.90317f
C1476 VTAIL.t4 VSUBS 0.329786f
C1477 VTAIL.t7 VSUBS 0.329786f
C1478 VTAIL.n396 VSUBS 2.58956f
C1479 VTAIL.n397 VSUBS 0.976629f
C1480 VTAIL.n398 VSUBS 0.026014f
C1481 VTAIL.n399 VSUBS 0.023766f
C1482 VTAIL.n400 VSUBS 0.012771f
C1483 VTAIL.n401 VSUBS 0.030185f
C1484 VTAIL.n402 VSUBS 0.013522f
C1485 VTAIL.n403 VSUBS 0.023766f
C1486 VTAIL.n404 VSUBS 0.012771f
C1487 VTAIL.n405 VSUBS 0.030185f
C1488 VTAIL.n406 VSUBS 0.013146f
C1489 VTAIL.n407 VSUBS 0.023766f
C1490 VTAIL.n408 VSUBS 0.013146f
C1491 VTAIL.n409 VSUBS 0.012771f
C1492 VTAIL.n410 VSUBS 0.030185f
C1493 VTAIL.n411 VSUBS 0.030185f
C1494 VTAIL.n412 VSUBS 0.013522f
C1495 VTAIL.n413 VSUBS 0.023766f
C1496 VTAIL.n414 VSUBS 0.012771f
C1497 VTAIL.n415 VSUBS 0.030185f
C1498 VTAIL.n416 VSUBS 0.013522f
C1499 VTAIL.n417 VSUBS 0.023766f
C1500 VTAIL.n418 VSUBS 0.012771f
C1501 VTAIL.n419 VSUBS 0.030185f
C1502 VTAIL.n420 VSUBS 0.013522f
C1503 VTAIL.n421 VSUBS 0.023766f
C1504 VTAIL.n422 VSUBS 0.012771f
C1505 VTAIL.n423 VSUBS 0.030185f
C1506 VTAIL.n424 VSUBS 0.013522f
C1507 VTAIL.n425 VSUBS 0.023766f
C1508 VTAIL.n426 VSUBS 0.012771f
C1509 VTAIL.n427 VSUBS 0.030185f
C1510 VTAIL.n428 VSUBS 0.013522f
C1511 VTAIL.n429 VSUBS 1.7937f
C1512 VTAIL.n430 VSUBS 0.012771f
C1513 VTAIL.t1 VSUBS 0.064772f
C1514 VTAIL.n431 VSUBS 0.185474f
C1515 VTAIL.n432 VSUBS 0.019203f
C1516 VTAIL.n433 VSUBS 0.022639f
C1517 VTAIL.n434 VSUBS 0.030185f
C1518 VTAIL.n435 VSUBS 0.013522f
C1519 VTAIL.n436 VSUBS 0.012771f
C1520 VTAIL.n437 VSUBS 0.023766f
C1521 VTAIL.n438 VSUBS 0.023766f
C1522 VTAIL.n439 VSUBS 0.012771f
C1523 VTAIL.n440 VSUBS 0.013522f
C1524 VTAIL.n441 VSUBS 0.030185f
C1525 VTAIL.n442 VSUBS 0.030185f
C1526 VTAIL.n443 VSUBS 0.013522f
C1527 VTAIL.n444 VSUBS 0.012771f
C1528 VTAIL.n445 VSUBS 0.023766f
C1529 VTAIL.n446 VSUBS 0.023766f
C1530 VTAIL.n447 VSUBS 0.012771f
C1531 VTAIL.n448 VSUBS 0.013522f
C1532 VTAIL.n449 VSUBS 0.030185f
C1533 VTAIL.n450 VSUBS 0.030185f
C1534 VTAIL.n451 VSUBS 0.013522f
C1535 VTAIL.n452 VSUBS 0.012771f
C1536 VTAIL.n453 VSUBS 0.023766f
C1537 VTAIL.n454 VSUBS 0.023766f
C1538 VTAIL.n455 VSUBS 0.012771f
C1539 VTAIL.n456 VSUBS 0.013522f
C1540 VTAIL.n457 VSUBS 0.030185f
C1541 VTAIL.n458 VSUBS 0.030185f
C1542 VTAIL.n459 VSUBS 0.013522f
C1543 VTAIL.n460 VSUBS 0.012771f
C1544 VTAIL.n461 VSUBS 0.023766f
C1545 VTAIL.n462 VSUBS 0.023766f
C1546 VTAIL.n463 VSUBS 0.012771f
C1547 VTAIL.n464 VSUBS 0.013522f
C1548 VTAIL.n465 VSUBS 0.030185f
C1549 VTAIL.n466 VSUBS 0.030185f
C1550 VTAIL.n467 VSUBS 0.013522f
C1551 VTAIL.n468 VSUBS 0.012771f
C1552 VTAIL.n469 VSUBS 0.023766f
C1553 VTAIL.n470 VSUBS 0.023766f
C1554 VTAIL.n471 VSUBS 0.012771f
C1555 VTAIL.n472 VSUBS 0.013522f
C1556 VTAIL.n473 VSUBS 0.030185f
C1557 VTAIL.n474 VSUBS 0.030185f
C1558 VTAIL.n475 VSUBS 0.013522f
C1559 VTAIL.n476 VSUBS 0.012771f
C1560 VTAIL.n477 VSUBS 0.023766f
C1561 VTAIL.n478 VSUBS 0.023766f
C1562 VTAIL.n479 VSUBS 0.012771f
C1563 VTAIL.n480 VSUBS 0.013522f
C1564 VTAIL.n481 VSUBS 0.030185f
C1565 VTAIL.n482 VSUBS 0.030185f
C1566 VTAIL.n483 VSUBS 0.013522f
C1567 VTAIL.n484 VSUBS 0.012771f
C1568 VTAIL.n485 VSUBS 0.023766f
C1569 VTAIL.n486 VSUBS 0.023766f
C1570 VTAIL.n487 VSUBS 0.012771f
C1571 VTAIL.n488 VSUBS 0.013522f
C1572 VTAIL.n489 VSUBS 0.030185f
C1573 VTAIL.n490 VSUBS 0.072737f
C1574 VTAIL.n491 VSUBS 0.013522f
C1575 VTAIL.n492 VSUBS 0.012771f
C1576 VTAIL.n493 VSUBS 0.056232f
C1577 VTAIL.n494 VSUBS 0.036603f
C1578 VTAIL.n495 VSUBS 0.257039f
C1579 VTAIL.n496 VSUBS 0.026014f
C1580 VTAIL.n497 VSUBS 0.023766f
C1581 VTAIL.n498 VSUBS 0.012771f
C1582 VTAIL.n499 VSUBS 0.030185f
C1583 VTAIL.n500 VSUBS 0.013522f
C1584 VTAIL.n501 VSUBS 0.023766f
C1585 VTAIL.n502 VSUBS 0.012771f
C1586 VTAIL.n503 VSUBS 0.030185f
C1587 VTAIL.n504 VSUBS 0.013146f
C1588 VTAIL.n505 VSUBS 0.023766f
C1589 VTAIL.n506 VSUBS 0.013146f
C1590 VTAIL.n507 VSUBS 0.012771f
C1591 VTAIL.n508 VSUBS 0.030185f
C1592 VTAIL.n509 VSUBS 0.030185f
C1593 VTAIL.n510 VSUBS 0.013522f
C1594 VTAIL.n511 VSUBS 0.023766f
C1595 VTAIL.n512 VSUBS 0.012771f
C1596 VTAIL.n513 VSUBS 0.030185f
C1597 VTAIL.n514 VSUBS 0.013522f
C1598 VTAIL.n515 VSUBS 0.023766f
C1599 VTAIL.n516 VSUBS 0.012771f
C1600 VTAIL.n517 VSUBS 0.030185f
C1601 VTAIL.n518 VSUBS 0.013522f
C1602 VTAIL.n519 VSUBS 0.023766f
C1603 VTAIL.n520 VSUBS 0.012771f
C1604 VTAIL.n521 VSUBS 0.030185f
C1605 VTAIL.n522 VSUBS 0.013522f
C1606 VTAIL.n523 VSUBS 0.023766f
C1607 VTAIL.n524 VSUBS 0.012771f
C1608 VTAIL.n525 VSUBS 0.030185f
C1609 VTAIL.n526 VSUBS 0.013522f
C1610 VTAIL.n527 VSUBS 1.7937f
C1611 VTAIL.n528 VSUBS 0.012771f
C1612 VTAIL.t10 VSUBS 0.064772f
C1613 VTAIL.n529 VSUBS 0.185474f
C1614 VTAIL.n530 VSUBS 0.019203f
C1615 VTAIL.n531 VSUBS 0.022639f
C1616 VTAIL.n532 VSUBS 0.030185f
C1617 VTAIL.n533 VSUBS 0.013522f
C1618 VTAIL.n534 VSUBS 0.012771f
C1619 VTAIL.n535 VSUBS 0.023766f
C1620 VTAIL.n536 VSUBS 0.023766f
C1621 VTAIL.n537 VSUBS 0.012771f
C1622 VTAIL.n538 VSUBS 0.013522f
C1623 VTAIL.n539 VSUBS 0.030185f
C1624 VTAIL.n540 VSUBS 0.030185f
C1625 VTAIL.n541 VSUBS 0.013522f
C1626 VTAIL.n542 VSUBS 0.012771f
C1627 VTAIL.n543 VSUBS 0.023766f
C1628 VTAIL.n544 VSUBS 0.023766f
C1629 VTAIL.n545 VSUBS 0.012771f
C1630 VTAIL.n546 VSUBS 0.013522f
C1631 VTAIL.n547 VSUBS 0.030185f
C1632 VTAIL.n548 VSUBS 0.030185f
C1633 VTAIL.n549 VSUBS 0.013522f
C1634 VTAIL.n550 VSUBS 0.012771f
C1635 VTAIL.n551 VSUBS 0.023766f
C1636 VTAIL.n552 VSUBS 0.023766f
C1637 VTAIL.n553 VSUBS 0.012771f
C1638 VTAIL.n554 VSUBS 0.013522f
C1639 VTAIL.n555 VSUBS 0.030185f
C1640 VTAIL.n556 VSUBS 0.030185f
C1641 VTAIL.n557 VSUBS 0.013522f
C1642 VTAIL.n558 VSUBS 0.012771f
C1643 VTAIL.n559 VSUBS 0.023766f
C1644 VTAIL.n560 VSUBS 0.023766f
C1645 VTAIL.n561 VSUBS 0.012771f
C1646 VTAIL.n562 VSUBS 0.013522f
C1647 VTAIL.n563 VSUBS 0.030185f
C1648 VTAIL.n564 VSUBS 0.030185f
C1649 VTAIL.n565 VSUBS 0.013522f
C1650 VTAIL.n566 VSUBS 0.012771f
C1651 VTAIL.n567 VSUBS 0.023766f
C1652 VTAIL.n568 VSUBS 0.023766f
C1653 VTAIL.n569 VSUBS 0.012771f
C1654 VTAIL.n570 VSUBS 0.013522f
C1655 VTAIL.n571 VSUBS 0.030185f
C1656 VTAIL.n572 VSUBS 0.030185f
C1657 VTAIL.n573 VSUBS 0.013522f
C1658 VTAIL.n574 VSUBS 0.012771f
C1659 VTAIL.n575 VSUBS 0.023766f
C1660 VTAIL.n576 VSUBS 0.023766f
C1661 VTAIL.n577 VSUBS 0.012771f
C1662 VTAIL.n578 VSUBS 0.013522f
C1663 VTAIL.n579 VSUBS 0.030185f
C1664 VTAIL.n580 VSUBS 0.030185f
C1665 VTAIL.n581 VSUBS 0.013522f
C1666 VTAIL.n582 VSUBS 0.012771f
C1667 VTAIL.n583 VSUBS 0.023766f
C1668 VTAIL.n584 VSUBS 0.023766f
C1669 VTAIL.n585 VSUBS 0.012771f
C1670 VTAIL.n586 VSUBS 0.013522f
C1671 VTAIL.n587 VSUBS 0.030185f
C1672 VTAIL.n588 VSUBS 0.072737f
C1673 VTAIL.n589 VSUBS 0.013522f
C1674 VTAIL.n590 VSUBS 0.012771f
C1675 VTAIL.n591 VSUBS 0.056232f
C1676 VTAIL.n592 VSUBS 0.036603f
C1677 VTAIL.n593 VSUBS 0.257039f
C1678 VTAIL.t8 VSUBS 0.329786f
C1679 VTAIL.t11 VSUBS 0.329786f
C1680 VTAIL.n594 VSUBS 2.58956f
C1681 VTAIL.n595 VSUBS 0.976629f
C1682 VTAIL.n596 VSUBS 0.026014f
C1683 VTAIL.n597 VSUBS 0.023766f
C1684 VTAIL.n598 VSUBS 0.012771f
C1685 VTAIL.n599 VSUBS 0.030185f
C1686 VTAIL.n600 VSUBS 0.013522f
C1687 VTAIL.n601 VSUBS 0.023766f
C1688 VTAIL.n602 VSUBS 0.012771f
C1689 VTAIL.n603 VSUBS 0.030185f
C1690 VTAIL.n604 VSUBS 0.013146f
C1691 VTAIL.n605 VSUBS 0.023766f
C1692 VTAIL.n606 VSUBS 0.013146f
C1693 VTAIL.n607 VSUBS 0.012771f
C1694 VTAIL.n608 VSUBS 0.030185f
C1695 VTAIL.n609 VSUBS 0.030185f
C1696 VTAIL.n610 VSUBS 0.013522f
C1697 VTAIL.n611 VSUBS 0.023766f
C1698 VTAIL.n612 VSUBS 0.012771f
C1699 VTAIL.n613 VSUBS 0.030185f
C1700 VTAIL.n614 VSUBS 0.013522f
C1701 VTAIL.n615 VSUBS 0.023766f
C1702 VTAIL.n616 VSUBS 0.012771f
C1703 VTAIL.n617 VSUBS 0.030185f
C1704 VTAIL.n618 VSUBS 0.013522f
C1705 VTAIL.n619 VSUBS 0.023766f
C1706 VTAIL.n620 VSUBS 0.012771f
C1707 VTAIL.n621 VSUBS 0.030185f
C1708 VTAIL.n622 VSUBS 0.013522f
C1709 VTAIL.n623 VSUBS 0.023766f
C1710 VTAIL.n624 VSUBS 0.012771f
C1711 VTAIL.n625 VSUBS 0.030185f
C1712 VTAIL.n626 VSUBS 0.013522f
C1713 VTAIL.n627 VSUBS 1.7937f
C1714 VTAIL.n628 VSUBS 0.012771f
C1715 VTAIL.t12 VSUBS 0.064772f
C1716 VTAIL.n629 VSUBS 0.185474f
C1717 VTAIL.n630 VSUBS 0.019203f
C1718 VTAIL.n631 VSUBS 0.022639f
C1719 VTAIL.n632 VSUBS 0.030185f
C1720 VTAIL.n633 VSUBS 0.013522f
C1721 VTAIL.n634 VSUBS 0.012771f
C1722 VTAIL.n635 VSUBS 0.023766f
C1723 VTAIL.n636 VSUBS 0.023766f
C1724 VTAIL.n637 VSUBS 0.012771f
C1725 VTAIL.n638 VSUBS 0.013522f
C1726 VTAIL.n639 VSUBS 0.030185f
C1727 VTAIL.n640 VSUBS 0.030185f
C1728 VTAIL.n641 VSUBS 0.013522f
C1729 VTAIL.n642 VSUBS 0.012771f
C1730 VTAIL.n643 VSUBS 0.023766f
C1731 VTAIL.n644 VSUBS 0.023766f
C1732 VTAIL.n645 VSUBS 0.012771f
C1733 VTAIL.n646 VSUBS 0.013522f
C1734 VTAIL.n647 VSUBS 0.030185f
C1735 VTAIL.n648 VSUBS 0.030185f
C1736 VTAIL.n649 VSUBS 0.013522f
C1737 VTAIL.n650 VSUBS 0.012771f
C1738 VTAIL.n651 VSUBS 0.023766f
C1739 VTAIL.n652 VSUBS 0.023766f
C1740 VTAIL.n653 VSUBS 0.012771f
C1741 VTAIL.n654 VSUBS 0.013522f
C1742 VTAIL.n655 VSUBS 0.030185f
C1743 VTAIL.n656 VSUBS 0.030185f
C1744 VTAIL.n657 VSUBS 0.013522f
C1745 VTAIL.n658 VSUBS 0.012771f
C1746 VTAIL.n659 VSUBS 0.023766f
C1747 VTAIL.n660 VSUBS 0.023766f
C1748 VTAIL.n661 VSUBS 0.012771f
C1749 VTAIL.n662 VSUBS 0.013522f
C1750 VTAIL.n663 VSUBS 0.030185f
C1751 VTAIL.n664 VSUBS 0.030185f
C1752 VTAIL.n665 VSUBS 0.013522f
C1753 VTAIL.n666 VSUBS 0.012771f
C1754 VTAIL.n667 VSUBS 0.023766f
C1755 VTAIL.n668 VSUBS 0.023766f
C1756 VTAIL.n669 VSUBS 0.012771f
C1757 VTAIL.n670 VSUBS 0.013522f
C1758 VTAIL.n671 VSUBS 0.030185f
C1759 VTAIL.n672 VSUBS 0.030185f
C1760 VTAIL.n673 VSUBS 0.013522f
C1761 VTAIL.n674 VSUBS 0.012771f
C1762 VTAIL.n675 VSUBS 0.023766f
C1763 VTAIL.n676 VSUBS 0.023766f
C1764 VTAIL.n677 VSUBS 0.012771f
C1765 VTAIL.n678 VSUBS 0.013522f
C1766 VTAIL.n679 VSUBS 0.030185f
C1767 VTAIL.n680 VSUBS 0.030185f
C1768 VTAIL.n681 VSUBS 0.013522f
C1769 VTAIL.n682 VSUBS 0.012771f
C1770 VTAIL.n683 VSUBS 0.023766f
C1771 VTAIL.n684 VSUBS 0.023766f
C1772 VTAIL.n685 VSUBS 0.012771f
C1773 VTAIL.n686 VSUBS 0.013522f
C1774 VTAIL.n687 VSUBS 0.030185f
C1775 VTAIL.n688 VSUBS 0.072737f
C1776 VTAIL.n689 VSUBS 0.013522f
C1777 VTAIL.n690 VSUBS 0.012771f
C1778 VTAIL.n691 VSUBS 0.056232f
C1779 VTAIL.n692 VSUBS 0.036603f
C1780 VTAIL.n693 VSUBS 1.90317f
C1781 VTAIL.n694 VSUBS 0.026014f
C1782 VTAIL.n695 VSUBS 0.023766f
C1783 VTAIL.n696 VSUBS 0.012771f
C1784 VTAIL.n697 VSUBS 0.030185f
C1785 VTAIL.n698 VSUBS 0.013522f
C1786 VTAIL.n699 VSUBS 0.023766f
C1787 VTAIL.n700 VSUBS 0.012771f
C1788 VTAIL.n701 VSUBS 0.030185f
C1789 VTAIL.n702 VSUBS 0.013146f
C1790 VTAIL.n703 VSUBS 0.023766f
C1791 VTAIL.n704 VSUBS 0.013522f
C1792 VTAIL.n705 VSUBS 0.030185f
C1793 VTAIL.n706 VSUBS 0.013522f
C1794 VTAIL.n707 VSUBS 0.023766f
C1795 VTAIL.n708 VSUBS 0.012771f
C1796 VTAIL.n709 VSUBS 0.030185f
C1797 VTAIL.n710 VSUBS 0.013522f
C1798 VTAIL.n711 VSUBS 0.023766f
C1799 VTAIL.n712 VSUBS 0.012771f
C1800 VTAIL.n713 VSUBS 0.030185f
C1801 VTAIL.n714 VSUBS 0.013522f
C1802 VTAIL.n715 VSUBS 0.023766f
C1803 VTAIL.n716 VSUBS 0.012771f
C1804 VTAIL.n717 VSUBS 0.030185f
C1805 VTAIL.n718 VSUBS 0.013522f
C1806 VTAIL.n719 VSUBS 0.023766f
C1807 VTAIL.n720 VSUBS 0.012771f
C1808 VTAIL.n721 VSUBS 0.030185f
C1809 VTAIL.n722 VSUBS 0.013522f
C1810 VTAIL.n723 VSUBS 1.7937f
C1811 VTAIL.n724 VSUBS 0.012771f
C1812 VTAIL.t0 VSUBS 0.064772f
C1813 VTAIL.n725 VSUBS 0.185474f
C1814 VTAIL.n726 VSUBS 0.019203f
C1815 VTAIL.n727 VSUBS 0.022639f
C1816 VTAIL.n728 VSUBS 0.030185f
C1817 VTAIL.n729 VSUBS 0.013522f
C1818 VTAIL.n730 VSUBS 0.012771f
C1819 VTAIL.n731 VSUBS 0.023766f
C1820 VTAIL.n732 VSUBS 0.023766f
C1821 VTAIL.n733 VSUBS 0.012771f
C1822 VTAIL.n734 VSUBS 0.013522f
C1823 VTAIL.n735 VSUBS 0.030185f
C1824 VTAIL.n736 VSUBS 0.030185f
C1825 VTAIL.n737 VSUBS 0.013522f
C1826 VTAIL.n738 VSUBS 0.012771f
C1827 VTAIL.n739 VSUBS 0.023766f
C1828 VTAIL.n740 VSUBS 0.023766f
C1829 VTAIL.n741 VSUBS 0.012771f
C1830 VTAIL.n742 VSUBS 0.013522f
C1831 VTAIL.n743 VSUBS 0.030185f
C1832 VTAIL.n744 VSUBS 0.030185f
C1833 VTAIL.n745 VSUBS 0.013522f
C1834 VTAIL.n746 VSUBS 0.012771f
C1835 VTAIL.n747 VSUBS 0.023766f
C1836 VTAIL.n748 VSUBS 0.023766f
C1837 VTAIL.n749 VSUBS 0.012771f
C1838 VTAIL.n750 VSUBS 0.013522f
C1839 VTAIL.n751 VSUBS 0.030185f
C1840 VTAIL.n752 VSUBS 0.030185f
C1841 VTAIL.n753 VSUBS 0.013522f
C1842 VTAIL.n754 VSUBS 0.012771f
C1843 VTAIL.n755 VSUBS 0.023766f
C1844 VTAIL.n756 VSUBS 0.023766f
C1845 VTAIL.n757 VSUBS 0.012771f
C1846 VTAIL.n758 VSUBS 0.013522f
C1847 VTAIL.n759 VSUBS 0.030185f
C1848 VTAIL.n760 VSUBS 0.030185f
C1849 VTAIL.n761 VSUBS 0.013522f
C1850 VTAIL.n762 VSUBS 0.012771f
C1851 VTAIL.n763 VSUBS 0.023766f
C1852 VTAIL.n764 VSUBS 0.023766f
C1853 VTAIL.n765 VSUBS 0.012771f
C1854 VTAIL.n766 VSUBS 0.012771f
C1855 VTAIL.n767 VSUBS 0.013522f
C1856 VTAIL.n768 VSUBS 0.030185f
C1857 VTAIL.n769 VSUBS 0.030185f
C1858 VTAIL.n770 VSUBS 0.030185f
C1859 VTAIL.n771 VSUBS 0.013146f
C1860 VTAIL.n772 VSUBS 0.012771f
C1861 VTAIL.n773 VSUBS 0.023766f
C1862 VTAIL.n774 VSUBS 0.023766f
C1863 VTAIL.n775 VSUBS 0.012771f
C1864 VTAIL.n776 VSUBS 0.013522f
C1865 VTAIL.n777 VSUBS 0.030185f
C1866 VTAIL.n778 VSUBS 0.030185f
C1867 VTAIL.n779 VSUBS 0.013522f
C1868 VTAIL.n780 VSUBS 0.012771f
C1869 VTAIL.n781 VSUBS 0.023766f
C1870 VTAIL.n782 VSUBS 0.023766f
C1871 VTAIL.n783 VSUBS 0.012771f
C1872 VTAIL.n784 VSUBS 0.013522f
C1873 VTAIL.n785 VSUBS 0.030185f
C1874 VTAIL.n786 VSUBS 0.072737f
C1875 VTAIL.n787 VSUBS 0.013522f
C1876 VTAIL.n788 VSUBS 0.012771f
C1877 VTAIL.n789 VSUBS 0.056232f
C1878 VTAIL.n790 VSUBS 0.036603f
C1879 VTAIL.n791 VSUBS 1.89871f
C1880 VP.n0 VSUBS 0.036417f
C1881 VP.t5 VSUBS 3.60066f
C1882 VP.n1 VSUBS 0.053642f
C1883 VP.n2 VSUBS 0.027623f
C1884 VP.t1 VSUBS 3.60066f
C1885 VP.n3 VSUBS 1.24873f
C1886 VP.n4 VSUBS 0.027623f
C1887 VP.n5 VSUBS 0.02231f
C1888 VP.n6 VSUBS 0.027623f
C1889 VP.t4 VSUBS 3.60066f
C1890 VP.n7 VSUBS 1.24873f
C1891 VP.n8 VSUBS 0.027623f
C1892 VP.n9 VSUBS 0.053642f
C1893 VP.n10 VSUBS 0.036417f
C1894 VP.t6 VSUBS 3.60066f
C1895 VP.n11 VSUBS 0.036417f
C1896 VP.t3 VSUBS 3.60066f
C1897 VP.n12 VSUBS 0.053642f
C1898 VP.n13 VSUBS 0.027623f
C1899 VP.t2 VSUBS 3.60066f
C1900 VP.n14 VSUBS 1.24873f
C1901 VP.n15 VSUBS 0.027623f
C1902 VP.n16 VSUBS 0.02231f
C1903 VP.n17 VSUBS 0.027623f
C1904 VP.t0 VSUBS 3.60066f
C1905 VP.n18 VSUBS 1.32021f
C1906 VP.t7 VSUBS 3.83431f
C1907 VP.n19 VSUBS 1.30416f
C1908 VP.n20 VSUBS 0.269279f
C1909 VP.n21 VSUBS 0.026695f
C1910 VP.n22 VSUBS 0.051225f
C1911 VP.n23 VSUBS 0.054612f
C1912 VP.n24 VSUBS 0.027623f
C1913 VP.n25 VSUBS 0.027623f
C1914 VP.n26 VSUBS 0.027623f
C1915 VP.n27 VSUBS 0.054612f
C1916 VP.n28 VSUBS 0.051225f
C1917 VP.n29 VSUBS 0.026695f
C1918 VP.n30 VSUBS 0.027623f
C1919 VP.n31 VSUBS 0.027623f
C1920 VP.n32 VSUBS 0.050466f
C1921 VP.n33 VSUBS 0.055264f
C1922 VP.n34 VSUBS 0.022629f
C1923 VP.n35 VSUBS 0.027623f
C1924 VP.n36 VSUBS 0.027623f
C1925 VP.n37 VSUBS 0.027623f
C1926 VP.n38 VSUBS 0.051225f
C1927 VP.n39 VSUBS 0.028213f
C1928 VP.n40 VSUBS 1.33301f
C1929 VP.n41 VSUBS 1.79026f
C1930 VP.n42 VSUBS 1.80821f
C1931 VP.n43 VSUBS 1.33301f
C1932 VP.n44 VSUBS 0.028213f
C1933 VP.n45 VSUBS 0.051225f
C1934 VP.n46 VSUBS 0.027623f
C1935 VP.n47 VSUBS 0.027623f
C1936 VP.n48 VSUBS 0.027623f
C1937 VP.n49 VSUBS 0.022629f
C1938 VP.n50 VSUBS 0.055264f
C1939 VP.n51 VSUBS 0.050466f
C1940 VP.n52 VSUBS 0.027623f
C1941 VP.n53 VSUBS 0.027623f
C1942 VP.n54 VSUBS 0.026695f
C1943 VP.n55 VSUBS 0.051225f
C1944 VP.n56 VSUBS 0.054612f
C1945 VP.n57 VSUBS 0.027623f
C1946 VP.n58 VSUBS 0.027623f
C1947 VP.n59 VSUBS 0.027623f
C1948 VP.n60 VSUBS 0.054612f
C1949 VP.n61 VSUBS 0.051225f
C1950 VP.n62 VSUBS 0.026695f
C1951 VP.n63 VSUBS 0.027623f
C1952 VP.n64 VSUBS 0.027623f
C1953 VP.n65 VSUBS 0.050466f
C1954 VP.n66 VSUBS 0.055264f
C1955 VP.n67 VSUBS 0.022629f
C1956 VP.n68 VSUBS 0.027623f
C1957 VP.n69 VSUBS 0.027623f
C1958 VP.n70 VSUBS 0.027623f
C1959 VP.n71 VSUBS 0.051225f
C1960 VP.n72 VSUBS 0.028213f
C1961 VP.n73 VSUBS 1.33301f
C1962 VP.n74 VSUBS 0.050749f
.ends

