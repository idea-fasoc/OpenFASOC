* NGSPICE file created from diff_pair_sample_1557.ext - technology: sky130A

.subckt diff_pair_sample_1557 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.8413 pd=17.55 as=6.7158 ps=35.22 w=17.22 l=0.37
X1 VDD2.t2 VN.t1 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.8413 pd=17.55 as=6.7158 ps=35.22 w=17.22 l=0.37
X2 VTAIL.t3 VP.t0 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=6.7158 pd=35.22 as=2.8413 ps=17.55 w=17.22 l=0.37
X3 VTAIL.t7 VN.t2 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=6.7158 pd=35.22 as=2.8413 ps=17.55 w=17.22 l=0.37
X4 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=6.7158 pd=35.22 as=0 ps=0 w=17.22 l=0.37
X5 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=6.7158 pd=35.22 as=0 ps=0 w=17.22 l=0.37
X6 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.7158 pd=35.22 as=0 ps=0 w=17.22 l=0.37
X7 VTAIL.t0 VP.t1 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=6.7158 pd=35.22 as=2.8413 ps=17.55 w=17.22 l=0.37
X8 VDD1.t1 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.8413 pd=17.55 as=6.7158 ps=35.22 w=17.22 l=0.37
X9 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.7158 pd=35.22 as=0 ps=0 w=17.22 l=0.37
X10 VTAIL.t4 VN.t3 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.7158 pd=35.22 as=2.8413 ps=17.55 w=17.22 l=0.37
X11 VDD1.t0 VP.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.8413 pd=17.55 as=6.7158 ps=35.22 w=17.22 l=0.37
R0 VN.n0 VN.t1 1251.9
R1 VN.n0 VN.t2 1251.9
R2 VN.n1 VN.t0 1251.9
R3 VN.n1 VN.t3 1251.9
R4 VN VN.n1 205.189
R5 VN VN.n0 161.351
R6 VTAIL.n5 VTAIL.t3 46.3367
R7 VTAIL.n4 VTAIL.t6 46.3367
R8 VTAIL.n3 VTAIL.t4 46.3367
R9 VTAIL.n7 VTAIL.t5 46.3366
R10 VTAIL.n0 VTAIL.t7 46.3366
R11 VTAIL.n1 VTAIL.t1 46.3366
R12 VTAIL.n2 VTAIL.t0 46.3366
R13 VTAIL.n6 VTAIL.t2 46.3366
R14 VTAIL.n7 VTAIL.n6 27.8324
R15 VTAIL.n3 VTAIL.n2 27.8324
R16 VTAIL.n4 VTAIL.n3 0.603948
R17 VTAIL.n6 VTAIL.n5 0.603948
R18 VTAIL.n2 VTAIL.n1 0.603948
R19 VTAIL.n5 VTAIL.n4 0.470328
R20 VTAIL.n1 VTAIL.n0 0.470328
R21 VTAIL VTAIL.n0 0.360414
R22 VTAIL VTAIL.n7 0.244034
R23 VDD2.n2 VDD2.n0 102.252
R24 VDD2.n2 VDD2.n1 61.8655
R25 VDD2.n1 VDD2.t0 1.15033
R26 VDD2.n1 VDD2.t3 1.15033
R27 VDD2.n0 VDD2.t1 1.15033
R28 VDD2.n0 VDD2.t2 1.15033
R29 VDD2 VDD2.n2 0.0586897
R30 B.n160 B.t4 1332.27
R31 B.n152 B.t15 1332.27
R32 B.n59 B.t12 1332.27
R33 B.n67 B.t8 1332.27
R34 B.n499 B.n498 585
R35 B.n501 B.n96 585
R36 B.n504 B.n503 585
R37 B.n505 B.n95 585
R38 B.n507 B.n506 585
R39 B.n509 B.n94 585
R40 B.n512 B.n511 585
R41 B.n513 B.n93 585
R42 B.n515 B.n514 585
R43 B.n517 B.n92 585
R44 B.n520 B.n519 585
R45 B.n521 B.n91 585
R46 B.n523 B.n522 585
R47 B.n525 B.n90 585
R48 B.n528 B.n527 585
R49 B.n529 B.n89 585
R50 B.n531 B.n530 585
R51 B.n533 B.n88 585
R52 B.n536 B.n535 585
R53 B.n537 B.n87 585
R54 B.n539 B.n538 585
R55 B.n541 B.n86 585
R56 B.n544 B.n543 585
R57 B.n545 B.n85 585
R58 B.n547 B.n546 585
R59 B.n549 B.n84 585
R60 B.n552 B.n551 585
R61 B.n553 B.n83 585
R62 B.n555 B.n554 585
R63 B.n557 B.n82 585
R64 B.n560 B.n559 585
R65 B.n561 B.n81 585
R66 B.n563 B.n562 585
R67 B.n565 B.n80 585
R68 B.n568 B.n567 585
R69 B.n569 B.n79 585
R70 B.n571 B.n570 585
R71 B.n573 B.n78 585
R72 B.n576 B.n575 585
R73 B.n577 B.n77 585
R74 B.n579 B.n578 585
R75 B.n581 B.n76 585
R76 B.n584 B.n583 585
R77 B.n585 B.n75 585
R78 B.n587 B.n586 585
R79 B.n589 B.n74 585
R80 B.n592 B.n591 585
R81 B.n593 B.n73 585
R82 B.n595 B.n594 585
R83 B.n597 B.n72 585
R84 B.n600 B.n599 585
R85 B.n601 B.n71 585
R86 B.n603 B.n602 585
R87 B.n605 B.n70 585
R88 B.n608 B.n607 585
R89 B.n609 B.n66 585
R90 B.n611 B.n610 585
R91 B.n613 B.n65 585
R92 B.n616 B.n615 585
R93 B.n617 B.n64 585
R94 B.n619 B.n618 585
R95 B.n621 B.n63 585
R96 B.n624 B.n623 585
R97 B.n625 B.n62 585
R98 B.n627 B.n626 585
R99 B.n629 B.n61 585
R100 B.n632 B.n631 585
R101 B.n634 B.n58 585
R102 B.n636 B.n635 585
R103 B.n638 B.n57 585
R104 B.n641 B.n640 585
R105 B.n642 B.n56 585
R106 B.n644 B.n643 585
R107 B.n646 B.n55 585
R108 B.n649 B.n648 585
R109 B.n650 B.n54 585
R110 B.n652 B.n651 585
R111 B.n654 B.n53 585
R112 B.n657 B.n656 585
R113 B.n658 B.n52 585
R114 B.n660 B.n659 585
R115 B.n662 B.n51 585
R116 B.n665 B.n664 585
R117 B.n666 B.n50 585
R118 B.n668 B.n667 585
R119 B.n670 B.n49 585
R120 B.n673 B.n672 585
R121 B.n674 B.n48 585
R122 B.n676 B.n675 585
R123 B.n678 B.n47 585
R124 B.n681 B.n680 585
R125 B.n682 B.n46 585
R126 B.n684 B.n683 585
R127 B.n686 B.n45 585
R128 B.n689 B.n688 585
R129 B.n690 B.n44 585
R130 B.n692 B.n691 585
R131 B.n694 B.n43 585
R132 B.n697 B.n696 585
R133 B.n698 B.n42 585
R134 B.n700 B.n699 585
R135 B.n702 B.n41 585
R136 B.n705 B.n704 585
R137 B.n706 B.n40 585
R138 B.n708 B.n707 585
R139 B.n710 B.n39 585
R140 B.n713 B.n712 585
R141 B.n714 B.n38 585
R142 B.n716 B.n715 585
R143 B.n718 B.n37 585
R144 B.n721 B.n720 585
R145 B.n722 B.n36 585
R146 B.n724 B.n723 585
R147 B.n726 B.n35 585
R148 B.n729 B.n728 585
R149 B.n730 B.n34 585
R150 B.n732 B.n731 585
R151 B.n734 B.n33 585
R152 B.n737 B.n736 585
R153 B.n738 B.n32 585
R154 B.n740 B.n739 585
R155 B.n742 B.n31 585
R156 B.n745 B.n744 585
R157 B.n746 B.n30 585
R158 B.n497 B.n28 585
R159 B.n749 B.n28 585
R160 B.n496 B.n27 585
R161 B.n750 B.n27 585
R162 B.n495 B.n26 585
R163 B.n751 B.n26 585
R164 B.n494 B.n493 585
R165 B.n493 B.n22 585
R166 B.n492 B.n21 585
R167 B.n757 B.n21 585
R168 B.n491 B.n20 585
R169 B.n758 B.n20 585
R170 B.n490 B.n19 585
R171 B.n759 B.n19 585
R172 B.n489 B.n488 585
R173 B.n488 B.n15 585
R174 B.n487 B.n14 585
R175 B.n765 B.n14 585
R176 B.n486 B.n13 585
R177 B.n766 B.n13 585
R178 B.n485 B.n12 585
R179 B.n767 B.n12 585
R180 B.n484 B.n483 585
R181 B.n483 B.n11 585
R182 B.n482 B.n7 585
R183 B.n773 B.n7 585
R184 B.n481 B.n6 585
R185 B.n774 B.n6 585
R186 B.n480 B.n5 585
R187 B.n775 B.n5 585
R188 B.n479 B.n478 585
R189 B.n478 B.n4 585
R190 B.n477 B.n97 585
R191 B.n477 B.n476 585
R192 B.n466 B.n98 585
R193 B.n469 B.n98 585
R194 B.n468 B.n467 585
R195 B.n470 B.n468 585
R196 B.n465 B.n102 585
R197 B.n106 B.n102 585
R198 B.n464 B.n463 585
R199 B.n463 B.n462 585
R200 B.n104 B.n103 585
R201 B.n105 B.n104 585
R202 B.n455 B.n454 585
R203 B.n456 B.n455 585
R204 B.n453 B.n111 585
R205 B.n111 B.n110 585
R206 B.n452 B.n451 585
R207 B.n451 B.n450 585
R208 B.n113 B.n112 585
R209 B.n114 B.n113 585
R210 B.n443 B.n442 585
R211 B.n444 B.n443 585
R212 B.n441 B.n119 585
R213 B.n119 B.n118 585
R214 B.n440 B.n439 585
R215 B.n439 B.n438 585
R216 B.n435 B.n123 585
R217 B.n434 B.n433 585
R218 B.n431 B.n124 585
R219 B.n431 B.n122 585
R220 B.n430 B.n429 585
R221 B.n428 B.n427 585
R222 B.n426 B.n126 585
R223 B.n424 B.n423 585
R224 B.n422 B.n127 585
R225 B.n421 B.n420 585
R226 B.n418 B.n128 585
R227 B.n416 B.n415 585
R228 B.n414 B.n129 585
R229 B.n413 B.n412 585
R230 B.n410 B.n130 585
R231 B.n408 B.n407 585
R232 B.n406 B.n131 585
R233 B.n405 B.n404 585
R234 B.n402 B.n132 585
R235 B.n400 B.n399 585
R236 B.n398 B.n133 585
R237 B.n397 B.n396 585
R238 B.n394 B.n134 585
R239 B.n392 B.n391 585
R240 B.n390 B.n135 585
R241 B.n389 B.n388 585
R242 B.n386 B.n136 585
R243 B.n384 B.n383 585
R244 B.n382 B.n137 585
R245 B.n381 B.n380 585
R246 B.n378 B.n138 585
R247 B.n376 B.n375 585
R248 B.n374 B.n139 585
R249 B.n373 B.n372 585
R250 B.n370 B.n140 585
R251 B.n368 B.n367 585
R252 B.n366 B.n141 585
R253 B.n365 B.n364 585
R254 B.n362 B.n142 585
R255 B.n360 B.n359 585
R256 B.n358 B.n143 585
R257 B.n357 B.n356 585
R258 B.n354 B.n144 585
R259 B.n352 B.n351 585
R260 B.n350 B.n145 585
R261 B.n349 B.n348 585
R262 B.n346 B.n146 585
R263 B.n344 B.n343 585
R264 B.n342 B.n147 585
R265 B.n341 B.n340 585
R266 B.n338 B.n148 585
R267 B.n336 B.n335 585
R268 B.n334 B.n149 585
R269 B.n333 B.n332 585
R270 B.n330 B.n150 585
R271 B.n328 B.n327 585
R272 B.n326 B.n151 585
R273 B.n325 B.n324 585
R274 B.n322 B.n321 585
R275 B.n320 B.n319 585
R276 B.n318 B.n156 585
R277 B.n316 B.n315 585
R278 B.n314 B.n157 585
R279 B.n313 B.n312 585
R280 B.n310 B.n158 585
R281 B.n308 B.n307 585
R282 B.n306 B.n159 585
R283 B.n305 B.n304 585
R284 B.n302 B.n301 585
R285 B.n300 B.n299 585
R286 B.n298 B.n164 585
R287 B.n296 B.n295 585
R288 B.n294 B.n165 585
R289 B.n293 B.n292 585
R290 B.n290 B.n166 585
R291 B.n288 B.n287 585
R292 B.n286 B.n167 585
R293 B.n285 B.n284 585
R294 B.n282 B.n168 585
R295 B.n280 B.n279 585
R296 B.n278 B.n169 585
R297 B.n277 B.n276 585
R298 B.n274 B.n170 585
R299 B.n272 B.n271 585
R300 B.n270 B.n171 585
R301 B.n269 B.n268 585
R302 B.n266 B.n172 585
R303 B.n264 B.n263 585
R304 B.n262 B.n173 585
R305 B.n261 B.n260 585
R306 B.n258 B.n174 585
R307 B.n256 B.n255 585
R308 B.n254 B.n175 585
R309 B.n253 B.n252 585
R310 B.n250 B.n176 585
R311 B.n248 B.n247 585
R312 B.n246 B.n177 585
R313 B.n245 B.n244 585
R314 B.n242 B.n178 585
R315 B.n240 B.n239 585
R316 B.n238 B.n179 585
R317 B.n237 B.n236 585
R318 B.n234 B.n180 585
R319 B.n232 B.n231 585
R320 B.n230 B.n181 585
R321 B.n229 B.n228 585
R322 B.n226 B.n182 585
R323 B.n224 B.n223 585
R324 B.n222 B.n183 585
R325 B.n221 B.n220 585
R326 B.n218 B.n184 585
R327 B.n216 B.n215 585
R328 B.n214 B.n185 585
R329 B.n213 B.n212 585
R330 B.n210 B.n186 585
R331 B.n208 B.n207 585
R332 B.n206 B.n187 585
R333 B.n205 B.n204 585
R334 B.n202 B.n188 585
R335 B.n200 B.n199 585
R336 B.n198 B.n189 585
R337 B.n197 B.n196 585
R338 B.n194 B.n190 585
R339 B.n192 B.n191 585
R340 B.n121 B.n120 585
R341 B.n122 B.n121 585
R342 B.n437 B.n436 585
R343 B.n438 B.n437 585
R344 B.n117 B.n116 585
R345 B.n118 B.n117 585
R346 B.n446 B.n445 585
R347 B.n445 B.n444 585
R348 B.n447 B.n115 585
R349 B.n115 B.n114 585
R350 B.n449 B.n448 585
R351 B.n450 B.n449 585
R352 B.n109 B.n108 585
R353 B.n110 B.n109 585
R354 B.n458 B.n457 585
R355 B.n457 B.n456 585
R356 B.n459 B.n107 585
R357 B.n107 B.n105 585
R358 B.n461 B.n460 585
R359 B.n462 B.n461 585
R360 B.n101 B.n100 585
R361 B.n106 B.n101 585
R362 B.n472 B.n471 585
R363 B.n471 B.n470 585
R364 B.n473 B.n99 585
R365 B.n469 B.n99 585
R366 B.n475 B.n474 585
R367 B.n476 B.n475 585
R368 B.n2 B.n0 585
R369 B.n4 B.n2 585
R370 B.n3 B.n1 585
R371 B.n774 B.n3 585
R372 B.n772 B.n771 585
R373 B.n773 B.n772 585
R374 B.n770 B.n8 585
R375 B.n11 B.n8 585
R376 B.n769 B.n768 585
R377 B.n768 B.n767 585
R378 B.n10 B.n9 585
R379 B.n766 B.n10 585
R380 B.n764 B.n763 585
R381 B.n765 B.n764 585
R382 B.n762 B.n16 585
R383 B.n16 B.n15 585
R384 B.n761 B.n760 585
R385 B.n760 B.n759 585
R386 B.n18 B.n17 585
R387 B.n758 B.n18 585
R388 B.n756 B.n755 585
R389 B.n757 B.n756 585
R390 B.n754 B.n23 585
R391 B.n23 B.n22 585
R392 B.n753 B.n752 585
R393 B.n752 B.n751 585
R394 B.n25 B.n24 585
R395 B.n750 B.n25 585
R396 B.n748 B.n747 585
R397 B.n749 B.n748 585
R398 B.n777 B.n776 585
R399 B.n776 B.n775 585
R400 B.n437 B.n123 516.524
R401 B.n748 B.n30 516.524
R402 B.n439 B.n121 516.524
R403 B.n499 B.n28 516.524
R404 B.n500 B.n29 256.663
R405 B.n502 B.n29 256.663
R406 B.n508 B.n29 256.663
R407 B.n510 B.n29 256.663
R408 B.n516 B.n29 256.663
R409 B.n518 B.n29 256.663
R410 B.n524 B.n29 256.663
R411 B.n526 B.n29 256.663
R412 B.n532 B.n29 256.663
R413 B.n534 B.n29 256.663
R414 B.n540 B.n29 256.663
R415 B.n542 B.n29 256.663
R416 B.n548 B.n29 256.663
R417 B.n550 B.n29 256.663
R418 B.n556 B.n29 256.663
R419 B.n558 B.n29 256.663
R420 B.n564 B.n29 256.663
R421 B.n566 B.n29 256.663
R422 B.n572 B.n29 256.663
R423 B.n574 B.n29 256.663
R424 B.n580 B.n29 256.663
R425 B.n582 B.n29 256.663
R426 B.n588 B.n29 256.663
R427 B.n590 B.n29 256.663
R428 B.n596 B.n29 256.663
R429 B.n598 B.n29 256.663
R430 B.n604 B.n29 256.663
R431 B.n606 B.n29 256.663
R432 B.n612 B.n29 256.663
R433 B.n614 B.n29 256.663
R434 B.n620 B.n29 256.663
R435 B.n622 B.n29 256.663
R436 B.n628 B.n29 256.663
R437 B.n630 B.n29 256.663
R438 B.n637 B.n29 256.663
R439 B.n639 B.n29 256.663
R440 B.n645 B.n29 256.663
R441 B.n647 B.n29 256.663
R442 B.n653 B.n29 256.663
R443 B.n655 B.n29 256.663
R444 B.n661 B.n29 256.663
R445 B.n663 B.n29 256.663
R446 B.n669 B.n29 256.663
R447 B.n671 B.n29 256.663
R448 B.n677 B.n29 256.663
R449 B.n679 B.n29 256.663
R450 B.n685 B.n29 256.663
R451 B.n687 B.n29 256.663
R452 B.n693 B.n29 256.663
R453 B.n695 B.n29 256.663
R454 B.n701 B.n29 256.663
R455 B.n703 B.n29 256.663
R456 B.n709 B.n29 256.663
R457 B.n711 B.n29 256.663
R458 B.n717 B.n29 256.663
R459 B.n719 B.n29 256.663
R460 B.n725 B.n29 256.663
R461 B.n727 B.n29 256.663
R462 B.n733 B.n29 256.663
R463 B.n735 B.n29 256.663
R464 B.n741 B.n29 256.663
R465 B.n743 B.n29 256.663
R466 B.n432 B.n122 256.663
R467 B.n125 B.n122 256.663
R468 B.n425 B.n122 256.663
R469 B.n419 B.n122 256.663
R470 B.n417 B.n122 256.663
R471 B.n411 B.n122 256.663
R472 B.n409 B.n122 256.663
R473 B.n403 B.n122 256.663
R474 B.n401 B.n122 256.663
R475 B.n395 B.n122 256.663
R476 B.n393 B.n122 256.663
R477 B.n387 B.n122 256.663
R478 B.n385 B.n122 256.663
R479 B.n379 B.n122 256.663
R480 B.n377 B.n122 256.663
R481 B.n371 B.n122 256.663
R482 B.n369 B.n122 256.663
R483 B.n363 B.n122 256.663
R484 B.n361 B.n122 256.663
R485 B.n355 B.n122 256.663
R486 B.n353 B.n122 256.663
R487 B.n347 B.n122 256.663
R488 B.n345 B.n122 256.663
R489 B.n339 B.n122 256.663
R490 B.n337 B.n122 256.663
R491 B.n331 B.n122 256.663
R492 B.n329 B.n122 256.663
R493 B.n323 B.n122 256.663
R494 B.n155 B.n122 256.663
R495 B.n317 B.n122 256.663
R496 B.n311 B.n122 256.663
R497 B.n309 B.n122 256.663
R498 B.n303 B.n122 256.663
R499 B.n163 B.n122 256.663
R500 B.n297 B.n122 256.663
R501 B.n291 B.n122 256.663
R502 B.n289 B.n122 256.663
R503 B.n283 B.n122 256.663
R504 B.n281 B.n122 256.663
R505 B.n275 B.n122 256.663
R506 B.n273 B.n122 256.663
R507 B.n267 B.n122 256.663
R508 B.n265 B.n122 256.663
R509 B.n259 B.n122 256.663
R510 B.n257 B.n122 256.663
R511 B.n251 B.n122 256.663
R512 B.n249 B.n122 256.663
R513 B.n243 B.n122 256.663
R514 B.n241 B.n122 256.663
R515 B.n235 B.n122 256.663
R516 B.n233 B.n122 256.663
R517 B.n227 B.n122 256.663
R518 B.n225 B.n122 256.663
R519 B.n219 B.n122 256.663
R520 B.n217 B.n122 256.663
R521 B.n211 B.n122 256.663
R522 B.n209 B.n122 256.663
R523 B.n203 B.n122 256.663
R524 B.n201 B.n122 256.663
R525 B.n195 B.n122 256.663
R526 B.n193 B.n122 256.663
R527 B.n437 B.n117 163.367
R528 B.n445 B.n117 163.367
R529 B.n445 B.n115 163.367
R530 B.n449 B.n115 163.367
R531 B.n449 B.n109 163.367
R532 B.n457 B.n109 163.367
R533 B.n457 B.n107 163.367
R534 B.n461 B.n107 163.367
R535 B.n461 B.n101 163.367
R536 B.n471 B.n101 163.367
R537 B.n471 B.n99 163.367
R538 B.n475 B.n99 163.367
R539 B.n475 B.n2 163.367
R540 B.n776 B.n2 163.367
R541 B.n776 B.n3 163.367
R542 B.n772 B.n3 163.367
R543 B.n772 B.n8 163.367
R544 B.n768 B.n8 163.367
R545 B.n768 B.n10 163.367
R546 B.n764 B.n10 163.367
R547 B.n764 B.n16 163.367
R548 B.n760 B.n16 163.367
R549 B.n760 B.n18 163.367
R550 B.n756 B.n18 163.367
R551 B.n756 B.n23 163.367
R552 B.n752 B.n23 163.367
R553 B.n752 B.n25 163.367
R554 B.n748 B.n25 163.367
R555 B.n433 B.n431 163.367
R556 B.n431 B.n430 163.367
R557 B.n427 B.n426 163.367
R558 B.n424 B.n127 163.367
R559 B.n420 B.n418 163.367
R560 B.n416 B.n129 163.367
R561 B.n412 B.n410 163.367
R562 B.n408 B.n131 163.367
R563 B.n404 B.n402 163.367
R564 B.n400 B.n133 163.367
R565 B.n396 B.n394 163.367
R566 B.n392 B.n135 163.367
R567 B.n388 B.n386 163.367
R568 B.n384 B.n137 163.367
R569 B.n380 B.n378 163.367
R570 B.n376 B.n139 163.367
R571 B.n372 B.n370 163.367
R572 B.n368 B.n141 163.367
R573 B.n364 B.n362 163.367
R574 B.n360 B.n143 163.367
R575 B.n356 B.n354 163.367
R576 B.n352 B.n145 163.367
R577 B.n348 B.n346 163.367
R578 B.n344 B.n147 163.367
R579 B.n340 B.n338 163.367
R580 B.n336 B.n149 163.367
R581 B.n332 B.n330 163.367
R582 B.n328 B.n151 163.367
R583 B.n324 B.n322 163.367
R584 B.n319 B.n318 163.367
R585 B.n316 B.n157 163.367
R586 B.n312 B.n310 163.367
R587 B.n308 B.n159 163.367
R588 B.n304 B.n302 163.367
R589 B.n299 B.n298 163.367
R590 B.n296 B.n165 163.367
R591 B.n292 B.n290 163.367
R592 B.n288 B.n167 163.367
R593 B.n284 B.n282 163.367
R594 B.n280 B.n169 163.367
R595 B.n276 B.n274 163.367
R596 B.n272 B.n171 163.367
R597 B.n268 B.n266 163.367
R598 B.n264 B.n173 163.367
R599 B.n260 B.n258 163.367
R600 B.n256 B.n175 163.367
R601 B.n252 B.n250 163.367
R602 B.n248 B.n177 163.367
R603 B.n244 B.n242 163.367
R604 B.n240 B.n179 163.367
R605 B.n236 B.n234 163.367
R606 B.n232 B.n181 163.367
R607 B.n228 B.n226 163.367
R608 B.n224 B.n183 163.367
R609 B.n220 B.n218 163.367
R610 B.n216 B.n185 163.367
R611 B.n212 B.n210 163.367
R612 B.n208 B.n187 163.367
R613 B.n204 B.n202 163.367
R614 B.n200 B.n189 163.367
R615 B.n196 B.n194 163.367
R616 B.n192 B.n121 163.367
R617 B.n439 B.n119 163.367
R618 B.n443 B.n119 163.367
R619 B.n443 B.n113 163.367
R620 B.n451 B.n113 163.367
R621 B.n451 B.n111 163.367
R622 B.n455 B.n111 163.367
R623 B.n455 B.n104 163.367
R624 B.n463 B.n104 163.367
R625 B.n463 B.n102 163.367
R626 B.n468 B.n102 163.367
R627 B.n468 B.n98 163.367
R628 B.n477 B.n98 163.367
R629 B.n478 B.n477 163.367
R630 B.n478 B.n5 163.367
R631 B.n6 B.n5 163.367
R632 B.n7 B.n6 163.367
R633 B.n483 B.n7 163.367
R634 B.n483 B.n12 163.367
R635 B.n13 B.n12 163.367
R636 B.n14 B.n13 163.367
R637 B.n488 B.n14 163.367
R638 B.n488 B.n19 163.367
R639 B.n20 B.n19 163.367
R640 B.n21 B.n20 163.367
R641 B.n493 B.n21 163.367
R642 B.n493 B.n26 163.367
R643 B.n27 B.n26 163.367
R644 B.n28 B.n27 163.367
R645 B.n744 B.n742 163.367
R646 B.n740 B.n32 163.367
R647 B.n736 B.n734 163.367
R648 B.n732 B.n34 163.367
R649 B.n728 B.n726 163.367
R650 B.n724 B.n36 163.367
R651 B.n720 B.n718 163.367
R652 B.n716 B.n38 163.367
R653 B.n712 B.n710 163.367
R654 B.n708 B.n40 163.367
R655 B.n704 B.n702 163.367
R656 B.n700 B.n42 163.367
R657 B.n696 B.n694 163.367
R658 B.n692 B.n44 163.367
R659 B.n688 B.n686 163.367
R660 B.n684 B.n46 163.367
R661 B.n680 B.n678 163.367
R662 B.n676 B.n48 163.367
R663 B.n672 B.n670 163.367
R664 B.n668 B.n50 163.367
R665 B.n664 B.n662 163.367
R666 B.n660 B.n52 163.367
R667 B.n656 B.n654 163.367
R668 B.n652 B.n54 163.367
R669 B.n648 B.n646 163.367
R670 B.n644 B.n56 163.367
R671 B.n640 B.n638 163.367
R672 B.n636 B.n58 163.367
R673 B.n631 B.n629 163.367
R674 B.n627 B.n62 163.367
R675 B.n623 B.n621 163.367
R676 B.n619 B.n64 163.367
R677 B.n615 B.n613 163.367
R678 B.n611 B.n66 163.367
R679 B.n607 B.n605 163.367
R680 B.n603 B.n71 163.367
R681 B.n599 B.n597 163.367
R682 B.n595 B.n73 163.367
R683 B.n591 B.n589 163.367
R684 B.n587 B.n75 163.367
R685 B.n583 B.n581 163.367
R686 B.n579 B.n77 163.367
R687 B.n575 B.n573 163.367
R688 B.n571 B.n79 163.367
R689 B.n567 B.n565 163.367
R690 B.n563 B.n81 163.367
R691 B.n559 B.n557 163.367
R692 B.n555 B.n83 163.367
R693 B.n551 B.n549 163.367
R694 B.n547 B.n85 163.367
R695 B.n543 B.n541 163.367
R696 B.n539 B.n87 163.367
R697 B.n535 B.n533 163.367
R698 B.n531 B.n89 163.367
R699 B.n527 B.n525 163.367
R700 B.n523 B.n91 163.367
R701 B.n519 B.n517 163.367
R702 B.n515 B.n93 163.367
R703 B.n511 B.n509 163.367
R704 B.n507 B.n95 163.367
R705 B.n503 B.n501 163.367
R706 B.n160 B.t7 85.1396
R707 B.n67 B.t10 85.1396
R708 B.n152 B.t17 85.1169
R709 B.n59 B.t13 85.1169
R710 B.n432 B.n123 71.676
R711 B.n430 B.n125 71.676
R712 B.n426 B.n425 71.676
R713 B.n419 B.n127 71.676
R714 B.n418 B.n417 71.676
R715 B.n411 B.n129 71.676
R716 B.n410 B.n409 71.676
R717 B.n403 B.n131 71.676
R718 B.n402 B.n401 71.676
R719 B.n395 B.n133 71.676
R720 B.n394 B.n393 71.676
R721 B.n387 B.n135 71.676
R722 B.n386 B.n385 71.676
R723 B.n379 B.n137 71.676
R724 B.n378 B.n377 71.676
R725 B.n371 B.n139 71.676
R726 B.n370 B.n369 71.676
R727 B.n363 B.n141 71.676
R728 B.n362 B.n361 71.676
R729 B.n355 B.n143 71.676
R730 B.n354 B.n353 71.676
R731 B.n347 B.n145 71.676
R732 B.n346 B.n345 71.676
R733 B.n339 B.n147 71.676
R734 B.n338 B.n337 71.676
R735 B.n331 B.n149 71.676
R736 B.n330 B.n329 71.676
R737 B.n323 B.n151 71.676
R738 B.n322 B.n155 71.676
R739 B.n318 B.n317 71.676
R740 B.n311 B.n157 71.676
R741 B.n310 B.n309 71.676
R742 B.n303 B.n159 71.676
R743 B.n302 B.n163 71.676
R744 B.n298 B.n297 71.676
R745 B.n291 B.n165 71.676
R746 B.n290 B.n289 71.676
R747 B.n283 B.n167 71.676
R748 B.n282 B.n281 71.676
R749 B.n275 B.n169 71.676
R750 B.n274 B.n273 71.676
R751 B.n267 B.n171 71.676
R752 B.n266 B.n265 71.676
R753 B.n259 B.n173 71.676
R754 B.n258 B.n257 71.676
R755 B.n251 B.n175 71.676
R756 B.n250 B.n249 71.676
R757 B.n243 B.n177 71.676
R758 B.n242 B.n241 71.676
R759 B.n235 B.n179 71.676
R760 B.n234 B.n233 71.676
R761 B.n227 B.n181 71.676
R762 B.n226 B.n225 71.676
R763 B.n219 B.n183 71.676
R764 B.n218 B.n217 71.676
R765 B.n211 B.n185 71.676
R766 B.n210 B.n209 71.676
R767 B.n203 B.n187 71.676
R768 B.n202 B.n201 71.676
R769 B.n195 B.n189 71.676
R770 B.n194 B.n193 71.676
R771 B.n743 B.n30 71.676
R772 B.n742 B.n741 71.676
R773 B.n735 B.n32 71.676
R774 B.n734 B.n733 71.676
R775 B.n727 B.n34 71.676
R776 B.n726 B.n725 71.676
R777 B.n719 B.n36 71.676
R778 B.n718 B.n717 71.676
R779 B.n711 B.n38 71.676
R780 B.n710 B.n709 71.676
R781 B.n703 B.n40 71.676
R782 B.n702 B.n701 71.676
R783 B.n695 B.n42 71.676
R784 B.n694 B.n693 71.676
R785 B.n687 B.n44 71.676
R786 B.n686 B.n685 71.676
R787 B.n679 B.n46 71.676
R788 B.n678 B.n677 71.676
R789 B.n671 B.n48 71.676
R790 B.n670 B.n669 71.676
R791 B.n663 B.n50 71.676
R792 B.n662 B.n661 71.676
R793 B.n655 B.n52 71.676
R794 B.n654 B.n653 71.676
R795 B.n647 B.n54 71.676
R796 B.n646 B.n645 71.676
R797 B.n639 B.n56 71.676
R798 B.n638 B.n637 71.676
R799 B.n630 B.n58 71.676
R800 B.n629 B.n628 71.676
R801 B.n622 B.n62 71.676
R802 B.n621 B.n620 71.676
R803 B.n614 B.n64 71.676
R804 B.n613 B.n612 71.676
R805 B.n606 B.n66 71.676
R806 B.n605 B.n604 71.676
R807 B.n598 B.n71 71.676
R808 B.n597 B.n596 71.676
R809 B.n590 B.n73 71.676
R810 B.n589 B.n588 71.676
R811 B.n582 B.n75 71.676
R812 B.n581 B.n580 71.676
R813 B.n574 B.n77 71.676
R814 B.n573 B.n572 71.676
R815 B.n566 B.n79 71.676
R816 B.n565 B.n564 71.676
R817 B.n558 B.n81 71.676
R818 B.n557 B.n556 71.676
R819 B.n550 B.n83 71.676
R820 B.n549 B.n548 71.676
R821 B.n542 B.n85 71.676
R822 B.n541 B.n540 71.676
R823 B.n534 B.n87 71.676
R824 B.n533 B.n532 71.676
R825 B.n526 B.n89 71.676
R826 B.n525 B.n524 71.676
R827 B.n518 B.n91 71.676
R828 B.n517 B.n516 71.676
R829 B.n510 B.n93 71.676
R830 B.n509 B.n508 71.676
R831 B.n502 B.n95 71.676
R832 B.n501 B.n500 71.676
R833 B.n500 B.n499 71.676
R834 B.n503 B.n502 71.676
R835 B.n508 B.n507 71.676
R836 B.n511 B.n510 71.676
R837 B.n516 B.n515 71.676
R838 B.n519 B.n518 71.676
R839 B.n524 B.n523 71.676
R840 B.n527 B.n526 71.676
R841 B.n532 B.n531 71.676
R842 B.n535 B.n534 71.676
R843 B.n540 B.n539 71.676
R844 B.n543 B.n542 71.676
R845 B.n548 B.n547 71.676
R846 B.n551 B.n550 71.676
R847 B.n556 B.n555 71.676
R848 B.n559 B.n558 71.676
R849 B.n564 B.n563 71.676
R850 B.n567 B.n566 71.676
R851 B.n572 B.n571 71.676
R852 B.n575 B.n574 71.676
R853 B.n580 B.n579 71.676
R854 B.n583 B.n582 71.676
R855 B.n588 B.n587 71.676
R856 B.n591 B.n590 71.676
R857 B.n596 B.n595 71.676
R858 B.n599 B.n598 71.676
R859 B.n604 B.n603 71.676
R860 B.n607 B.n606 71.676
R861 B.n612 B.n611 71.676
R862 B.n615 B.n614 71.676
R863 B.n620 B.n619 71.676
R864 B.n623 B.n622 71.676
R865 B.n628 B.n627 71.676
R866 B.n631 B.n630 71.676
R867 B.n637 B.n636 71.676
R868 B.n640 B.n639 71.676
R869 B.n645 B.n644 71.676
R870 B.n648 B.n647 71.676
R871 B.n653 B.n652 71.676
R872 B.n656 B.n655 71.676
R873 B.n661 B.n660 71.676
R874 B.n664 B.n663 71.676
R875 B.n669 B.n668 71.676
R876 B.n672 B.n671 71.676
R877 B.n677 B.n676 71.676
R878 B.n680 B.n679 71.676
R879 B.n685 B.n684 71.676
R880 B.n688 B.n687 71.676
R881 B.n693 B.n692 71.676
R882 B.n696 B.n695 71.676
R883 B.n701 B.n700 71.676
R884 B.n704 B.n703 71.676
R885 B.n709 B.n708 71.676
R886 B.n712 B.n711 71.676
R887 B.n717 B.n716 71.676
R888 B.n720 B.n719 71.676
R889 B.n725 B.n724 71.676
R890 B.n728 B.n727 71.676
R891 B.n733 B.n732 71.676
R892 B.n736 B.n735 71.676
R893 B.n741 B.n740 71.676
R894 B.n744 B.n743 71.676
R895 B.n433 B.n432 71.676
R896 B.n427 B.n125 71.676
R897 B.n425 B.n424 71.676
R898 B.n420 B.n419 71.676
R899 B.n417 B.n416 71.676
R900 B.n412 B.n411 71.676
R901 B.n409 B.n408 71.676
R902 B.n404 B.n403 71.676
R903 B.n401 B.n400 71.676
R904 B.n396 B.n395 71.676
R905 B.n393 B.n392 71.676
R906 B.n388 B.n387 71.676
R907 B.n385 B.n384 71.676
R908 B.n380 B.n379 71.676
R909 B.n377 B.n376 71.676
R910 B.n372 B.n371 71.676
R911 B.n369 B.n368 71.676
R912 B.n364 B.n363 71.676
R913 B.n361 B.n360 71.676
R914 B.n356 B.n355 71.676
R915 B.n353 B.n352 71.676
R916 B.n348 B.n347 71.676
R917 B.n345 B.n344 71.676
R918 B.n340 B.n339 71.676
R919 B.n337 B.n336 71.676
R920 B.n332 B.n331 71.676
R921 B.n329 B.n328 71.676
R922 B.n324 B.n323 71.676
R923 B.n319 B.n155 71.676
R924 B.n317 B.n316 71.676
R925 B.n312 B.n311 71.676
R926 B.n309 B.n308 71.676
R927 B.n304 B.n303 71.676
R928 B.n299 B.n163 71.676
R929 B.n297 B.n296 71.676
R930 B.n292 B.n291 71.676
R931 B.n289 B.n288 71.676
R932 B.n284 B.n283 71.676
R933 B.n281 B.n280 71.676
R934 B.n276 B.n275 71.676
R935 B.n273 B.n272 71.676
R936 B.n268 B.n267 71.676
R937 B.n265 B.n264 71.676
R938 B.n260 B.n259 71.676
R939 B.n257 B.n256 71.676
R940 B.n252 B.n251 71.676
R941 B.n249 B.n248 71.676
R942 B.n244 B.n243 71.676
R943 B.n241 B.n240 71.676
R944 B.n236 B.n235 71.676
R945 B.n233 B.n232 71.676
R946 B.n228 B.n227 71.676
R947 B.n225 B.n224 71.676
R948 B.n220 B.n219 71.676
R949 B.n217 B.n216 71.676
R950 B.n212 B.n211 71.676
R951 B.n209 B.n208 71.676
R952 B.n204 B.n203 71.676
R953 B.n201 B.n200 71.676
R954 B.n196 B.n195 71.676
R955 B.n193 B.n192 71.676
R956 B.n161 B.t6 71.5639
R957 B.n68 B.t11 71.5639
R958 B.n153 B.t16 71.5412
R959 B.n60 B.t14 71.5412
R960 B.n438 B.n122 69.865
R961 B.n749 B.n29 69.865
R962 B.n162 B.n161 59.5399
R963 B.n154 B.n153 59.5399
R964 B.n633 B.n60 59.5399
R965 B.n69 B.n68 59.5399
R966 B.n747 B.n746 33.5615
R967 B.n498 B.n497 33.5615
R968 B.n440 B.n120 33.5615
R969 B.n436 B.n435 33.5615
R970 B.n438 B.n118 33.2228
R971 B.n444 B.n118 33.2228
R972 B.n444 B.n114 33.2228
R973 B.n450 B.n114 33.2228
R974 B.n456 B.n110 33.2228
R975 B.n456 B.n105 33.2228
R976 B.n462 B.n105 33.2228
R977 B.n462 B.n106 33.2228
R978 B.n470 B.n469 33.2228
R979 B.n476 B.n4 33.2228
R980 B.n775 B.n4 33.2228
R981 B.n775 B.n774 33.2228
R982 B.n774 B.n773 33.2228
R983 B.n767 B.n11 33.2228
R984 B.n766 B.n765 33.2228
R985 B.n765 B.n15 33.2228
R986 B.n759 B.n15 33.2228
R987 B.n759 B.n758 33.2228
R988 B.n757 B.n22 33.2228
R989 B.n751 B.n22 33.2228
R990 B.n751 B.n750 33.2228
R991 B.n750 B.n749 33.2228
R992 B.t5 B.n110 31.7571
R993 B.n758 B.t9 31.7571
R994 B.n470 B.t0 22.963
R995 B.n767 B.t2 22.963
R996 B.n476 B.t1 21.0087
R997 B.n773 B.t3 21.0087
R998 B B.n777 18.0485
R999 B.n161 B.n160 13.5763
R1000 B.n153 B.n152 13.5763
R1001 B.n60 B.n59 13.5763
R1002 B.n68 B.n67 13.5763
R1003 B.n469 B.t1 12.2146
R1004 B.n11 B.t3 12.2146
R1005 B.n746 B.n745 10.6151
R1006 B.n745 B.n31 10.6151
R1007 B.n739 B.n31 10.6151
R1008 B.n739 B.n738 10.6151
R1009 B.n738 B.n737 10.6151
R1010 B.n737 B.n33 10.6151
R1011 B.n731 B.n33 10.6151
R1012 B.n731 B.n730 10.6151
R1013 B.n730 B.n729 10.6151
R1014 B.n729 B.n35 10.6151
R1015 B.n723 B.n35 10.6151
R1016 B.n723 B.n722 10.6151
R1017 B.n722 B.n721 10.6151
R1018 B.n721 B.n37 10.6151
R1019 B.n715 B.n37 10.6151
R1020 B.n715 B.n714 10.6151
R1021 B.n714 B.n713 10.6151
R1022 B.n713 B.n39 10.6151
R1023 B.n707 B.n39 10.6151
R1024 B.n707 B.n706 10.6151
R1025 B.n706 B.n705 10.6151
R1026 B.n705 B.n41 10.6151
R1027 B.n699 B.n41 10.6151
R1028 B.n699 B.n698 10.6151
R1029 B.n698 B.n697 10.6151
R1030 B.n697 B.n43 10.6151
R1031 B.n691 B.n43 10.6151
R1032 B.n691 B.n690 10.6151
R1033 B.n690 B.n689 10.6151
R1034 B.n689 B.n45 10.6151
R1035 B.n683 B.n45 10.6151
R1036 B.n683 B.n682 10.6151
R1037 B.n682 B.n681 10.6151
R1038 B.n681 B.n47 10.6151
R1039 B.n675 B.n47 10.6151
R1040 B.n675 B.n674 10.6151
R1041 B.n674 B.n673 10.6151
R1042 B.n673 B.n49 10.6151
R1043 B.n667 B.n49 10.6151
R1044 B.n667 B.n666 10.6151
R1045 B.n666 B.n665 10.6151
R1046 B.n665 B.n51 10.6151
R1047 B.n659 B.n51 10.6151
R1048 B.n659 B.n658 10.6151
R1049 B.n658 B.n657 10.6151
R1050 B.n657 B.n53 10.6151
R1051 B.n651 B.n53 10.6151
R1052 B.n651 B.n650 10.6151
R1053 B.n650 B.n649 10.6151
R1054 B.n649 B.n55 10.6151
R1055 B.n643 B.n55 10.6151
R1056 B.n643 B.n642 10.6151
R1057 B.n642 B.n641 10.6151
R1058 B.n641 B.n57 10.6151
R1059 B.n635 B.n57 10.6151
R1060 B.n635 B.n634 10.6151
R1061 B.n632 B.n61 10.6151
R1062 B.n626 B.n61 10.6151
R1063 B.n626 B.n625 10.6151
R1064 B.n625 B.n624 10.6151
R1065 B.n624 B.n63 10.6151
R1066 B.n618 B.n63 10.6151
R1067 B.n618 B.n617 10.6151
R1068 B.n617 B.n616 10.6151
R1069 B.n616 B.n65 10.6151
R1070 B.n610 B.n609 10.6151
R1071 B.n609 B.n608 10.6151
R1072 B.n608 B.n70 10.6151
R1073 B.n602 B.n70 10.6151
R1074 B.n602 B.n601 10.6151
R1075 B.n601 B.n600 10.6151
R1076 B.n600 B.n72 10.6151
R1077 B.n594 B.n72 10.6151
R1078 B.n594 B.n593 10.6151
R1079 B.n593 B.n592 10.6151
R1080 B.n592 B.n74 10.6151
R1081 B.n586 B.n74 10.6151
R1082 B.n586 B.n585 10.6151
R1083 B.n585 B.n584 10.6151
R1084 B.n584 B.n76 10.6151
R1085 B.n578 B.n76 10.6151
R1086 B.n578 B.n577 10.6151
R1087 B.n577 B.n576 10.6151
R1088 B.n576 B.n78 10.6151
R1089 B.n570 B.n78 10.6151
R1090 B.n570 B.n569 10.6151
R1091 B.n569 B.n568 10.6151
R1092 B.n568 B.n80 10.6151
R1093 B.n562 B.n80 10.6151
R1094 B.n562 B.n561 10.6151
R1095 B.n561 B.n560 10.6151
R1096 B.n560 B.n82 10.6151
R1097 B.n554 B.n82 10.6151
R1098 B.n554 B.n553 10.6151
R1099 B.n553 B.n552 10.6151
R1100 B.n552 B.n84 10.6151
R1101 B.n546 B.n84 10.6151
R1102 B.n546 B.n545 10.6151
R1103 B.n545 B.n544 10.6151
R1104 B.n544 B.n86 10.6151
R1105 B.n538 B.n86 10.6151
R1106 B.n538 B.n537 10.6151
R1107 B.n537 B.n536 10.6151
R1108 B.n536 B.n88 10.6151
R1109 B.n530 B.n88 10.6151
R1110 B.n530 B.n529 10.6151
R1111 B.n529 B.n528 10.6151
R1112 B.n528 B.n90 10.6151
R1113 B.n522 B.n90 10.6151
R1114 B.n522 B.n521 10.6151
R1115 B.n521 B.n520 10.6151
R1116 B.n520 B.n92 10.6151
R1117 B.n514 B.n92 10.6151
R1118 B.n514 B.n513 10.6151
R1119 B.n513 B.n512 10.6151
R1120 B.n512 B.n94 10.6151
R1121 B.n506 B.n94 10.6151
R1122 B.n506 B.n505 10.6151
R1123 B.n505 B.n504 10.6151
R1124 B.n504 B.n96 10.6151
R1125 B.n498 B.n96 10.6151
R1126 B.n441 B.n440 10.6151
R1127 B.n442 B.n441 10.6151
R1128 B.n442 B.n112 10.6151
R1129 B.n452 B.n112 10.6151
R1130 B.n453 B.n452 10.6151
R1131 B.n454 B.n453 10.6151
R1132 B.n454 B.n103 10.6151
R1133 B.n464 B.n103 10.6151
R1134 B.n465 B.n464 10.6151
R1135 B.n467 B.n465 10.6151
R1136 B.n467 B.n466 10.6151
R1137 B.n466 B.n97 10.6151
R1138 B.n479 B.n97 10.6151
R1139 B.n480 B.n479 10.6151
R1140 B.n481 B.n480 10.6151
R1141 B.n482 B.n481 10.6151
R1142 B.n484 B.n482 10.6151
R1143 B.n485 B.n484 10.6151
R1144 B.n486 B.n485 10.6151
R1145 B.n487 B.n486 10.6151
R1146 B.n489 B.n487 10.6151
R1147 B.n490 B.n489 10.6151
R1148 B.n491 B.n490 10.6151
R1149 B.n492 B.n491 10.6151
R1150 B.n494 B.n492 10.6151
R1151 B.n495 B.n494 10.6151
R1152 B.n496 B.n495 10.6151
R1153 B.n497 B.n496 10.6151
R1154 B.n435 B.n434 10.6151
R1155 B.n434 B.n124 10.6151
R1156 B.n429 B.n124 10.6151
R1157 B.n429 B.n428 10.6151
R1158 B.n428 B.n126 10.6151
R1159 B.n423 B.n126 10.6151
R1160 B.n423 B.n422 10.6151
R1161 B.n422 B.n421 10.6151
R1162 B.n421 B.n128 10.6151
R1163 B.n415 B.n128 10.6151
R1164 B.n415 B.n414 10.6151
R1165 B.n414 B.n413 10.6151
R1166 B.n413 B.n130 10.6151
R1167 B.n407 B.n130 10.6151
R1168 B.n407 B.n406 10.6151
R1169 B.n406 B.n405 10.6151
R1170 B.n405 B.n132 10.6151
R1171 B.n399 B.n132 10.6151
R1172 B.n399 B.n398 10.6151
R1173 B.n398 B.n397 10.6151
R1174 B.n397 B.n134 10.6151
R1175 B.n391 B.n134 10.6151
R1176 B.n391 B.n390 10.6151
R1177 B.n390 B.n389 10.6151
R1178 B.n389 B.n136 10.6151
R1179 B.n383 B.n136 10.6151
R1180 B.n383 B.n382 10.6151
R1181 B.n382 B.n381 10.6151
R1182 B.n381 B.n138 10.6151
R1183 B.n375 B.n138 10.6151
R1184 B.n375 B.n374 10.6151
R1185 B.n374 B.n373 10.6151
R1186 B.n373 B.n140 10.6151
R1187 B.n367 B.n140 10.6151
R1188 B.n367 B.n366 10.6151
R1189 B.n366 B.n365 10.6151
R1190 B.n365 B.n142 10.6151
R1191 B.n359 B.n142 10.6151
R1192 B.n359 B.n358 10.6151
R1193 B.n358 B.n357 10.6151
R1194 B.n357 B.n144 10.6151
R1195 B.n351 B.n144 10.6151
R1196 B.n351 B.n350 10.6151
R1197 B.n350 B.n349 10.6151
R1198 B.n349 B.n146 10.6151
R1199 B.n343 B.n146 10.6151
R1200 B.n343 B.n342 10.6151
R1201 B.n342 B.n341 10.6151
R1202 B.n341 B.n148 10.6151
R1203 B.n335 B.n148 10.6151
R1204 B.n335 B.n334 10.6151
R1205 B.n334 B.n333 10.6151
R1206 B.n333 B.n150 10.6151
R1207 B.n327 B.n150 10.6151
R1208 B.n327 B.n326 10.6151
R1209 B.n326 B.n325 10.6151
R1210 B.n321 B.n320 10.6151
R1211 B.n320 B.n156 10.6151
R1212 B.n315 B.n156 10.6151
R1213 B.n315 B.n314 10.6151
R1214 B.n314 B.n313 10.6151
R1215 B.n313 B.n158 10.6151
R1216 B.n307 B.n158 10.6151
R1217 B.n307 B.n306 10.6151
R1218 B.n306 B.n305 10.6151
R1219 B.n301 B.n300 10.6151
R1220 B.n300 B.n164 10.6151
R1221 B.n295 B.n164 10.6151
R1222 B.n295 B.n294 10.6151
R1223 B.n294 B.n293 10.6151
R1224 B.n293 B.n166 10.6151
R1225 B.n287 B.n166 10.6151
R1226 B.n287 B.n286 10.6151
R1227 B.n286 B.n285 10.6151
R1228 B.n285 B.n168 10.6151
R1229 B.n279 B.n168 10.6151
R1230 B.n279 B.n278 10.6151
R1231 B.n278 B.n277 10.6151
R1232 B.n277 B.n170 10.6151
R1233 B.n271 B.n170 10.6151
R1234 B.n271 B.n270 10.6151
R1235 B.n270 B.n269 10.6151
R1236 B.n269 B.n172 10.6151
R1237 B.n263 B.n172 10.6151
R1238 B.n263 B.n262 10.6151
R1239 B.n262 B.n261 10.6151
R1240 B.n261 B.n174 10.6151
R1241 B.n255 B.n174 10.6151
R1242 B.n255 B.n254 10.6151
R1243 B.n254 B.n253 10.6151
R1244 B.n253 B.n176 10.6151
R1245 B.n247 B.n176 10.6151
R1246 B.n247 B.n246 10.6151
R1247 B.n246 B.n245 10.6151
R1248 B.n245 B.n178 10.6151
R1249 B.n239 B.n178 10.6151
R1250 B.n239 B.n238 10.6151
R1251 B.n238 B.n237 10.6151
R1252 B.n237 B.n180 10.6151
R1253 B.n231 B.n180 10.6151
R1254 B.n231 B.n230 10.6151
R1255 B.n230 B.n229 10.6151
R1256 B.n229 B.n182 10.6151
R1257 B.n223 B.n182 10.6151
R1258 B.n223 B.n222 10.6151
R1259 B.n222 B.n221 10.6151
R1260 B.n221 B.n184 10.6151
R1261 B.n215 B.n184 10.6151
R1262 B.n215 B.n214 10.6151
R1263 B.n214 B.n213 10.6151
R1264 B.n213 B.n186 10.6151
R1265 B.n207 B.n186 10.6151
R1266 B.n207 B.n206 10.6151
R1267 B.n206 B.n205 10.6151
R1268 B.n205 B.n188 10.6151
R1269 B.n199 B.n188 10.6151
R1270 B.n199 B.n198 10.6151
R1271 B.n198 B.n197 10.6151
R1272 B.n197 B.n190 10.6151
R1273 B.n191 B.n190 10.6151
R1274 B.n191 B.n120 10.6151
R1275 B.n436 B.n116 10.6151
R1276 B.n446 B.n116 10.6151
R1277 B.n447 B.n446 10.6151
R1278 B.n448 B.n447 10.6151
R1279 B.n448 B.n108 10.6151
R1280 B.n458 B.n108 10.6151
R1281 B.n459 B.n458 10.6151
R1282 B.n460 B.n459 10.6151
R1283 B.n460 B.n100 10.6151
R1284 B.n472 B.n100 10.6151
R1285 B.n473 B.n472 10.6151
R1286 B.n474 B.n473 10.6151
R1287 B.n474 B.n0 10.6151
R1288 B.n771 B.n1 10.6151
R1289 B.n771 B.n770 10.6151
R1290 B.n770 B.n769 10.6151
R1291 B.n769 B.n9 10.6151
R1292 B.n763 B.n9 10.6151
R1293 B.n763 B.n762 10.6151
R1294 B.n762 B.n761 10.6151
R1295 B.n761 B.n17 10.6151
R1296 B.n755 B.n17 10.6151
R1297 B.n755 B.n754 10.6151
R1298 B.n754 B.n753 10.6151
R1299 B.n753 B.n24 10.6151
R1300 B.n747 B.n24 10.6151
R1301 B.n106 B.t0 10.2603
R1302 B.t2 B.n766 10.2603
R1303 B.n634 B.n633 8.74196
R1304 B.n610 B.n69 8.74196
R1305 B.n325 B.n154 8.74196
R1306 B.n301 B.n162 8.74196
R1307 B.n777 B.n0 2.81026
R1308 B.n777 B.n1 2.81026
R1309 B.n633 B.n632 1.87367
R1310 B.n69 B.n65 1.87367
R1311 B.n321 B.n154 1.87367
R1312 B.n305 B.n162 1.87367
R1313 B.n450 B.t5 1.46619
R1314 B.t9 B.n757 1.46619
R1315 VP.n1 VP.t2 1251.9
R1316 VP.n1 VP.t1 1251.9
R1317 VP.n0 VP.t3 1251.9
R1318 VP.n0 VP.t0 1251.9
R1319 VP.n2 VP.n0 204.809
R1320 VP.n2 VP.n1 161.3
R1321 VP VP.n2 0.0516364
R1322 VDD1 VDD1.n1 102.778
R1323 VDD1 VDD1.n0 61.9237
R1324 VDD1.n0 VDD1.t3 1.15033
R1325 VDD1.n0 VDD1.t0 1.15033
R1326 VDD1.n1 VDD1.t2 1.15033
R1327 VDD1.n1 VDD1.t1 1.15033
C0 VDD2 VTAIL 11.937799f
C1 VDD1 VP 3.30855f
C2 VDD1 VN 0.148459f
C3 VTAIL VDD1 11.898499f
C4 VDD2 VDD1 0.49323f
C5 VN VP 5.54055f
C6 VTAIL VP 2.49012f
C7 VTAIL VN 2.47602f
C8 VDD2 VP 0.253881f
C9 VDD2 VN 3.2033f
C10 VDD2 B 2.923644f
C11 VDD1 B 7.66451f
C12 VTAIL B 11.479221f
C13 VN B 9.370379f
C14 VP B 4.555239f
C15 VDD1.t3 B 0.433322f
C16 VDD1.t0 B 0.433322f
C17 VDD1.n0 B 3.94236f
C18 VDD1.t2 B 0.433322f
C19 VDD1.t1 B 0.433322f
C20 VDD1.n1 B 4.85323f
C21 VP.t0 B 1.0876f
C22 VP.t3 B 1.0876f
C23 VP.n0 B 1.37525f
C24 VP.t1 B 1.0876f
C25 VP.t2 B 1.0876f
C26 VP.n1 B 0.815681f
C27 VP.n2 B 4.72425f
C28 VDD2.t1 B 0.433828f
C29 VDD2.t2 B 0.433828f
C30 VDD2.n0 B 4.82649f
C31 VDD2.t0 B 0.433828f
C32 VDD2.t3 B 0.433828f
C33 VDD2.n1 B 3.94665f
C34 VDD2.n2 B 4.5227f
C35 VTAIL.t7 B 2.74835f
C36 VTAIL.n0 B 0.286579f
C37 VTAIL.t1 B 2.74835f
C38 VTAIL.n1 B 0.300551f
C39 VTAIL.t0 B 2.74835f
C40 VTAIL.n2 B 1.40276f
C41 VTAIL.t4 B 2.74836f
C42 VTAIL.n3 B 1.40274f
C43 VTAIL.t6 B 2.74836f
C44 VTAIL.n4 B 0.300534f
C45 VTAIL.t3 B 2.74836f
C46 VTAIL.n5 B 0.300534f
C47 VTAIL.t2 B 2.74835f
C48 VTAIL.n6 B 1.40276f
C49 VTAIL.t5 B 2.74835f
C50 VTAIL.n7 B 1.38211f
C51 VN.t2 B 1.07002f
C52 VN.t1 B 1.07002f
C53 VN.n0 B 0.802519f
C54 VN.t3 B 1.07002f
C55 VN.t0 B 1.07002f
C56 VN.n1 B 1.36504f
.ends

