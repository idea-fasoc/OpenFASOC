* NGSPICE file created from diff_pair_sample_0784.ext - technology: sky130A

.subckt diff_pair_sample_0784 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=7.683 pd=40.18 as=0 ps=0 w=19.7 l=3.06
X1 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=7.683 pd=40.18 as=0 ps=0 w=19.7 l=3.06
X2 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=7.683 pd=40.18 as=0 ps=0 w=19.7 l=3.06
X3 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=7.683 pd=40.18 as=0 ps=0 w=19.7 l=3.06
X4 VDD2.t1 VN.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=7.683 pd=40.18 as=7.683 ps=40.18 w=19.7 l=3.06
X5 VDD2.t0 VN.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=7.683 pd=40.18 as=7.683 ps=40.18 w=19.7 l=3.06
X6 VDD1.t1 VP.t0 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=7.683 pd=40.18 as=7.683 ps=40.18 w=19.7 l=3.06
X7 VDD1.t0 VP.t1 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=7.683 pd=40.18 as=7.683 ps=40.18 w=19.7 l=3.06
R0 B.n926 B.n925 585
R1 B.n400 B.n123 585
R2 B.n399 B.n398 585
R3 B.n397 B.n396 585
R4 B.n395 B.n394 585
R5 B.n393 B.n392 585
R6 B.n391 B.n390 585
R7 B.n389 B.n388 585
R8 B.n387 B.n386 585
R9 B.n385 B.n384 585
R10 B.n383 B.n382 585
R11 B.n381 B.n380 585
R12 B.n379 B.n378 585
R13 B.n377 B.n376 585
R14 B.n375 B.n374 585
R15 B.n373 B.n372 585
R16 B.n371 B.n370 585
R17 B.n369 B.n368 585
R18 B.n367 B.n366 585
R19 B.n365 B.n364 585
R20 B.n363 B.n362 585
R21 B.n361 B.n360 585
R22 B.n359 B.n358 585
R23 B.n357 B.n356 585
R24 B.n355 B.n354 585
R25 B.n353 B.n352 585
R26 B.n351 B.n350 585
R27 B.n349 B.n348 585
R28 B.n347 B.n346 585
R29 B.n345 B.n344 585
R30 B.n343 B.n342 585
R31 B.n341 B.n340 585
R32 B.n339 B.n338 585
R33 B.n337 B.n336 585
R34 B.n335 B.n334 585
R35 B.n333 B.n332 585
R36 B.n331 B.n330 585
R37 B.n329 B.n328 585
R38 B.n327 B.n326 585
R39 B.n325 B.n324 585
R40 B.n323 B.n322 585
R41 B.n321 B.n320 585
R42 B.n319 B.n318 585
R43 B.n317 B.n316 585
R44 B.n315 B.n314 585
R45 B.n313 B.n312 585
R46 B.n311 B.n310 585
R47 B.n309 B.n308 585
R48 B.n307 B.n306 585
R49 B.n305 B.n304 585
R50 B.n303 B.n302 585
R51 B.n301 B.n300 585
R52 B.n299 B.n298 585
R53 B.n297 B.n296 585
R54 B.n295 B.n294 585
R55 B.n293 B.n292 585
R56 B.n291 B.n290 585
R57 B.n289 B.n288 585
R58 B.n287 B.n286 585
R59 B.n285 B.n284 585
R60 B.n283 B.n282 585
R61 B.n281 B.n280 585
R62 B.n279 B.n278 585
R63 B.n277 B.n276 585
R64 B.n275 B.n274 585
R65 B.n273 B.n272 585
R66 B.n271 B.n270 585
R67 B.n269 B.n268 585
R68 B.n267 B.n266 585
R69 B.n265 B.n264 585
R70 B.n263 B.n262 585
R71 B.n261 B.n260 585
R72 B.n259 B.n258 585
R73 B.n257 B.n256 585
R74 B.n255 B.n254 585
R75 B.n253 B.n252 585
R76 B.n251 B.n250 585
R77 B.n249 B.n248 585
R78 B.n247 B.n246 585
R79 B.n245 B.n244 585
R80 B.n243 B.n242 585
R81 B.n241 B.n240 585
R82 B.n239 B.n238 585
R83 B.n237 B.n236 585
R84 B.n235 B.n234 585
R85 B.n233 B.n232 585
R86 B.n231 B.n230 585
R87 B.n229 B.n228 585
R88 B.n227 B.n226 585
R89 B.n225 B.n224 585
R90 B.n223 B.n222 585
R91 B.n221 B.n220 585
R92 B.n219 B.n218 585
R93 B.n217 B.n216 585
R94 B.n215 B.n214 585
R95 B.n213 B.n212 585
R96 B.n211 B.n210 585
R97 B.n209 B.n208 585
R98 B.n207 B.n206 585
R99 B.n205 B.n204 585
R100 B.n203 B.n202 585
R101 B.n201 B.n200 585
R102 B.n199 B.n198 585
R103 B.n197 B.n196 585
R104 B.n195 B.n194 585
R105 B.n193 B.n192 585
R106 B.n191 B.n190 585
R107 B.n189 B.n188 585
R108 B.n187 B.n186 585
R109 B.n185 B.n184 585
R110 B.n183 B.n182 585
R111 B.n181 B.n180 585
R112 B.n179 B.n178 585
R113 B.n177 B.n176 585
R114 B.n175 B.n174 585
R115 B.n173 B.n172 585
R116 B.n171 B.n170 585
R117 B.n169 B.n168 585
R118 B.n167 B.n166 585
R119 B.n165 B.n164 585
R120 B.n163 B.n162 585
R121 B.n161 B.n160 585
R122 B.n159 B.n158 585
R123 B.n157 B.n156 585
R124 B.n155 B.n154 585
R125 B.n153 B.n152 585
R126 B.n151 B.n150 585
R127 B.n149 B.n148 585
R128 B.n147 B.n146 585
R129 B.n145 B.n144 585
R130 B.n143 B.n142 585
R131 B.n141 B.n140 585
R132 B.n139 B.n138 585
R133 B.n137 B.n136 585
R134 B.n135 B.n134 585
R135 B.n133 B.n132 585
R136 B.n131 B.n130 585
R137 B.n53 B.n52 585
R138 B.n924 B.n54 585
R139 B.n929 B.n54 585
R140 B.n923 B.n922 585
R141 B.n922 B.n50 585
R142 B.n921 B.n49 585
R143 B.n935 B.n49 585
R144 B.n920 B.n48 585
R145 B.n936 B.n48 585
R146 B.n919 B.n47 585
R147 B.n937 B.n47 585
R148 B.n918 B.n917 585
R149 B.n917 B.n43 585
R150 B.n916 B.n42 585
R151 B.n943 B.n42 585
R152 B.n915 B.n41 585
R153 B.n944 B.n41 585
R154 B.n914 B.n40 585
R155 B.n945 B.n40 585
R156 B.n913 B.n912 585
R157 B.n912 B.n36 585
R158 B.n911 B.n35 585
R159 B.n951 B.n35 585
R160 B.n910 B.n34 585
R161 B.n952 B.n34 585
R162 B.n909 B.n33 585
R163 B.n953 B.n33 585
R164 B.n908 B.n907 585
R165 B.n907 B.n29 585
R166 B.n906 B.n28 585
R167 B.n959 B.n28 585
R168 B.n905 B.n27 585
R169 B.n960 B.n27 585
R170 B.n904 B.n26 585
R171 B.n961 B.n26 585
R172 B.n903 B.n902 585
R173 B.n902 B.n22 585
R174 B.n901 B.n21 585
R175 B.n967 B.n21 585
R176 B.n900 B.n20 585
R177 B.n968 B.n20 585
R178 B.n899 B.n19 585
R179 B.n969 B.n19 585
R180 B.n898 B.n897 585
R181 B.n897 B.n18 585
R182 B.n896 B.n14 585
R183 B.n975 B.n14 585
R184 B.n895 B.n13 585
R185 B.n976 B.n13 585
R186 B.n894 B.n12 585
R187 B.n977 B.n12 585
R188 B.n893 B.n892 585
R189 B.n892 B.n8 585
R190 B.n891 B.n7 585
R191 B.n983 B.n7 585
R192 B.n890 B.n6 585
R193 B.n984 B.n6 585
R194 B.n889 B.n5 585
R195 B.n985 B.n5 585
R196 B.n888 B.n887 585
R197 B.n887 B.n4 585
R198 B.n886 B.n401 585
R199 B.n886 B.n885 585
R200 B.n876 B.n402 585
R201 B.n403 B.n402 585
R202 B.n878 B.n877 585
R203 B.n879 B.n878 585
R204 B.n875 B.n408 585
R205 B.n408 B.n407 585
R206 B.n874 B.n873 585
R207 B.n873 B.n872 585
R208 B.n410 B.n409 585
R209 B.n865 B.n410 585
R210 B.n864 B.n863 585
R211 B.n866 B.n864 585
R212 B.n862 B.n415 585
R213 B.n415 B.n414 585
R214 B.n861 B.n860 585
R215 B.n860 B.n859 585
R216 B.n417 B.n416 585
R217 B.n418 B.n417 585
R218 B.n852 B.n851 585
R219 B.n853 B.n852 585
R220 B.n850 B.n423 585
R221 B.n423 B.n422 585
R222 B.n849 B.n848 585
R223 B.n848 B.n847 585
R224 B.n425 B.n424 585
R225 B.n426 B.n425 585
R226 B.n840 B.n839 585
R227 B.n841 B.n840 585
R228 B.n838 B.n431 585
R229 B.n431 B.n430 585
R230 B.n837 B.n836 585
R231 B.n836 B.n835 585
R232 B.n433 B.n432 585
R233 B.n434 B.n433 585
R234 B.n828 B.n827 585
R235 B.n829 B.n828 585
R236 B.n826 B.n439 585
R237 B.n439 B.n438 585
R238 B.n825 B.n824 585
R239 B.n824 B.n823 585
R240 B.n441 B.n440 585
R241 B.n442 B.n441 585
R242 B.n816 B.n815 585
R243 B.n817 B.n816 585
R244 B.n814 B.n447 585
R245 B.n447 B.n446 585
R246 B.n813 B.n812 585
R247 B.n812 B.n811 585
R248 B.n449 B.n448 585
R249 B.n450 B.n449 585
R250 B.n804 B.n803 585
R251 B.n805 B.n804 585
R252 B.n453 B.n452 585
R253 B.n528 B.n526 585
R254 B.n529 B.n525 585
R255 B.n529 B.n454 585
R256 B.n532 B.n531 585
R257 B.n533 B.n524 585
R258 B.n535 B.n534 585
R259 B.n537 B.n523 585
R260 B.n540 B.n539 585
R261 B.n541 B.n522 585
R262 B.n543 B.n542 585
R263 B.n545 B.n521 585
R264 B.n548 B.n547 585
R265 B.n549 B.n520 585
R266 B.n551 B.n550 585
R267 B.n553 B.n519 585
R268 B.n556 B.n555 585
R269 B.n557 B.n518 585
R270 B.n559 B.n558 585
R271 B.n561 B.n517 585
R272 B.n564 B.n563 585
R273 B.n565 B.n516 585
R274 B.n567 B.n566 585
R275 B.n569 B.n515 585
R276 B.n572 B.n571 585
R277 B.n573 B.n514 585
R278 B.n575 B.n574 585
R279 B.n577 B.n513 585
R280 B.n580 B.n579 585
R281 B.n581 B.n512 585
R282 B.n583 B.n582 585
R283 B.n585 B.n511 585
R284 B.n588 B.n587 585
R285 B.n589 B.n510 585
R286 B.n591 B.n590 585
R287 B.n593 B.n509 585
R288 B.n596 B.n595 585
R289 B.n597 B.n508 585
R290 B.n599 B.n598 585
R291 B.n601 B.n507 585
R292 B.n604 B.n603 585
R293 B.n605 B.n506 585
R294 B.n607 B.n606 585
R295 B.n609 B.n505 585
R296 B.n612 B.n611 585
R297 B.n613 B.n504 585
R298 B.n615 B.n614 585
R299 B.n617 B.n503 585
R300 B.n620 B.n619 585
R301 B.n621 B.n502 585
R302 B.n623 B.n622 585
R303 B.n625 B.n501 585
R304 B.n628 B.n627 585
R305 B.n629 B.n500 585
R306 B.n631 B.n630 585
R307 B.n633 B.n499 585
R308 B.n636 B.n635 585
R309 B.n637 B.n498 585
R310 B.n639 B.n638 585
R311 B.n641 B.n497 585
R312 B.n644 B.n643 585
R313 B.n645 B.n496 585
R314 B.n647 B.n646 585
R315 B.n649 B.n495 585
R316 B.n652 B.n651 585
R317 B.n654 B.n492 585
R318 B.n656 B.n655 585
R319 B.n658 B.n491 585
R320 B.n661 B.n660 585
R321 B.n662 B.n490 585
R322 B.n664 B.n663 585
R323 B.n666 B.n489 585
R324 B.n669 B.n668 585
R325 B.n670 B.n488 585
R326 B.n675 B.n674 585
R327 B.n677 B.n487 585
R328 B.n680 B.n679 585
R329 B.n681 B.n486 585
R330 B.n683 B.n682 585
R331 B.n685 B.n485 585
R332 B.n688 B.n687 585
R333 B.n689 B.n484 585
R334 B.n691 B.n690 585
R335 B.n693 B.n483 585
R336 B.n696 B.n695 585
R337 B.n697 B.n482 585
R338 B.n699 B.n698 585
R339 B.n701 B.n481 585
R340 B.n704 B.n703 585
R341 B.n705 B.n480 585
R342 B.n707 B.n706 585
R343 B.n709 B.n479 585
R344 B.n712 B.n711 585
R345 B.n713 B.n478 585
R346 B.n715 B.n714 585
R347 B.n717 B.n477 585
R348 B.n720 B.n719 585
R349 B.n721 B.n476 585
R350 B.n723 B.n722 585
R351 B.n725 B.n475 585
R352 B.n728 B.n727 585
R353 B.n729 B.n474 585
R354 B.n731 B.n730 585
R355 B.n733 B.n473 585
R356 B.n736 B.n735 585
R357 B.n737 B.n472 585
R358 B.n739 B.n738 585
R359 B.n741 B.n471 585
R360 B.n744 B.n743 585
R361 B.n745 B.n470 585
R362 B.n747 B.n746 585
R363 B.n749 B.n469 585
R364 B.n752 B.n751 585
R365 B.n753 B.n468 585
R366 B.n755 B.n754 585
R367 B.n757 B.n467 585
R368 B.n760 B.n759 585
R369 B.n761 B.n466 585
R370 B.n763 B.n762 585
R371 B.n765 B.n465 585
R372 B.n768 B.n767 585
R373 B.n769 B.n464 585
R374 B.n771 B.n770 585
R375 B.n773 B.n463 585
R376 B.n776 B.n775 585
R377 B.n777 B.n462 585
R378 B.n779 B.n778 585
R379 B.n781 B.n461 585
R380 B.n784 B.n783 585
R381 B.n785 B.n460 585
R382 B.n787 B.n786 585
R383 B.n789 B.n459 585
R384 B.n792 B.n791 585
R385 B.n793 B.n458 585
R386 B.n795 B.n794 585
R387 B.n797 B.n457 585
R388 B.n798 B.n456 585
R389 B.n801 B.n800 585
R390 B.n802 B.n455 585
R391 B.n455 B.n454 585
R392 B.n807 B.n806 585
R393 B.n806 B.n805 585
R394 B.n808 B.n451 585
R395 B.n451 B.n450 585
R396 B.n810 B.n809 585
R397 B.n811 B.n810 585
R398 B.n445 B.n444 585
R399 B.n446 B.n445 585
R400 B.n819 B.n818 585
R401 B.n818 B.n817 585
R402 B.n820 B.n443 585
R403 B.n443 B.n442 585
R404 B.n822 B.n821 585
R405 B.n823 B.n822 585
R406 B.n437 B.n436 585
R407 B.n438 B.n437 585
R408 B.n831 B.n830 585
R409 B.n830 B.n829 585
R410 B.n832 B.n435 585
R411 B.n435 B.n434 585
R412 B.n834 B.n833 585
R413 B.n835 B.n834 585
R414 B.n429 B.n428 585
R415 B.n430 B.n429 585
R416 B.n843 B.n842 585
R417 B.n842 B.n841 585
R418 B.n844 B.n427 585
R419 B.n427 B.n426 585
R420 B.n846 B.n845 585
R421 B.n847 B.n846 585
R422 B.n421 B.n420 585
R423 B.n422 B.n421 585
R424 B.n855 B.n854 585
R425 B.n854 B.n853 585
R426 B.n856 B.n419 585
R427 B.n419 B.n418 585
R428 B.n858 B.n857 585
R429 B.n859 B.n858 585
R430 B.n413 B.n412 585
R431 B.n414 B.n413 585
R432 B.n868 B.n867 585
R433 B.n867 B.n866 585
R434 B.n869 B.n411 585
R435 B.n865 B.n411 585
R436 B.n871 B.n870 585
R437 B.n872 B.n871 585
R438 B.n406 B.n405 585
R439 B.n407 B.n406 585
R440 B.n881 B.n880 585
R441 B.n880 B.n879 585
R442 B.n882 B.n404 585
R443 B.n404 B.n403 585
R444 B.n884 B.n883 585
R445 B.n885 B.n884 585
R446 B.n2 B.n0 585
R447 B.n4 B.n2 585
R448 B.n3 B.n1 585
R449 B.n984 B.n3 585
R450 B.n982 B.n981 585
R451 B.n983 B.n982 585
R452 B.n980 B.n9 585
R453 B.n9 B.n8 585
R454 B.n979 B.n978 585
R455 B.n978 B.n977 585
R456 B.n11 B.n10 585
R457 B.n976 B.n11 585
R458 B.n974 B.n973 585
R459 B.n975 B.n974 585
R460 B.n972 B.n15 585
R461 B.n18 B.n15 585
R462 B.n971 B.n970 585
R463 B.n970 B.n969 585
R464 B.n17 B.n16 585
R465 B.n968 B.n17 585
R466 B.n966 B.n965 585
R467 B.n967 B.n966 585
R468 B.n964 B.n23 585
R469 B.n23 B.n22 585
R470 B.n963 B.n962 585
R471 B.n962 B.n961 585
R472 B.n25 B.n24 585
R473 B.n960 B.n25 585
R474 B.n958 B.n957 585
R475 B.n959 B.n958 585
R476 B.n956 B.n30 585
R477 B.n30 B.n29 585
R478 B.n955 B.n954 585
R479 B.n954 B.n953 585
R480 B.n32 B.n31 585
R481 B.n952 B.n32 585
R482 B.n950 B.n949 585
R483 B.n951 B.n950 585
R484 B.n948 B.n37 585
R485 B.n37 B.n36 585
R486 B.n947 B.n946 585
R487 B.n946 B.n945 585
R488 B.n39 B.n38 585
R489 B.n944 B.n39 585
R490 B.n942 B.n941 585
R491 B.n943 B.n942 585
R492 B.n940 B.n44 585
R493 B.n44 B.n43 585
R494 B.n939 B.n938 585
R495 B.n938 B.n937 585
R496 B.n46 B.n45 585
R497 B.n936 B.n46 585
R498 B.n934 B.n933 585
R499 B.n935 B.n934 585
R500 B.n932 B.n51 585
R501 B.n51 B.n50 585
R502 B.n931 B.n930 585
R503 B.n930 B.n929 585
R504 B.n987 B.n986 585
R505 B.n986 B.n985 585
R506 B.n806 B.n453 516.524
R507 B.n930 B.n53 516.524
R508 B.n804 B.n455 516.524
R509 B.n926 B.n54 516.524
R510 B.n671 B.t15 480.856
R511 B.n124 B.t4 480.856
R512 B.n493 B.t12 480.856
R513 B.n127 B.t7 480.856
R514 B.n672 B.t14 415.111
R515 B.n125 B.t5 415.111
R516 B.n494 B.t11 415.111
R517 B.n128 B.t8 415.111
R518 B.n671 B.t13 363.803
R519 B.n493 B.t9 363.803
R520 B.n127 B.t6 363.803
R521 B.n124 B.t2 363.803
R522 B.n928 B.n927 256.663
R523 B.n928 B.n122 256.663
R524 B.n928 B.n121 256.663
R525 B.n928 B.n120 256.663
R526 B.n928 B.n119 256.663
R527 B.n928 B.n118 256.663
R528 B.n928 B.n117 256.663
R529 B.n928 B.n116 256.663
R530 B.n928 B.n115 256.663
R531 B.n928 B.n114 256.663
R532 B.n928 B.n113 256.663
R533 B.n928 B.n112 256.663
R534 B.n928 B.n111 256.663
R535 B.n928 B.n110 256.663
R536 B.n928 B.n109 256.663
R537 B.n928 B.n108 256.663
R538 B.n928 B.n107 256.663
R539 B.n928 B.n106 256.663
R540 B.n928 B.n105 256.663
R541 B.n928 B.n104 256.663
R542 B.n928 B.n103 256.663
R543 B.n928 B.n102 256.663
R544 B.n928 B.n101 256.663
R545 B.n928 B.n100 256.663
R546 B.n928 B.n99 256.663
R547 B.n928 B.n98 256.663
R548 B.n928 B.n97 256.663
R549 B.n928 B.n96 256.663
R550 B.n928 B.n95 256.663
R551 B.n928 B.n94 256.663
R552 B.n928 B.n93 256.663
R553 B.n928 B.n92 256.663
R554 B.n928 B.n91 256.663
R555 B.n928 B.n90 256.663
R556 B.n928 B.n89 256.663
R557 B.n928 B.n88 256.663
R558 B.n928 B.n87 256.663
R559 B.n928 B.n86 256.663
R560 B.n928 B.n85 256.663
R561 B.n928 B.n84 256.663
R562 B.n928 B.n83 256.663
R563 B.n928 B.n82 256.663
R564 B.n928 B.n81 256.663
R565 B.n928 B.n80 256.663
R566 B.n928 B.n79 256.663
R567 B.n928 B.n78 256.663
R568 B.n928 B.n77 256.663
R569 B.n928 B.n76 256.663
R570 B.n928 B.n75 256.663
R571 B.n928 B.n74 256.663
R572 B.n928 B.n73 256.663
R573 B.n928 B.n72 256.663
R574 B.n928 B.n71 256.663
R575 B.n928 B.n70 256.663
R576 B.n928 B.n69 256.663
R577 B.n928 B.n68 256.663
R578 B.n928 B.n67 256.663
R579 B.n928 B.n66 256.663
R580 B.n928 B.n65 256.663
R581 B.n928 B.n64 256.663
R582 B.n928 B.n63 256.663
R583 B.n928 B.n62 256.663
R584 B.n928 B.n61 256.663
R585 B.n928 B.n60 256.663
R586 B.n928 B.n59 256.663
R587 B.n928 B.n58 256.663
R588 B.n928 B.n57 256.663
R589 B.n928 B.n56 256.663
R590 B.n928 B.n55 256.663
R591 B.n527 B.n454 256.663
R592 B.n530 B.n454 256.663
R593 B.n536 B.n454 256.663
R594 B.n538 B.n454 256.663
R595 B.n544 B.n454 256.663
R596 B.n546 B.n454 256.663
R597 B.n552 B.n454 256.663
R598 B.n554 B.n454 256.663
R599 B.n560 B.n454 256.663
R600 B.n562 B.n454 256.663
R601 B.n568 B.n454 256.663
R602 B.n570 B.n454 256.663
R603 B.n576 B.n454 256.663
R604 B.n578 B.n454 256.663
R605 B.n584 B.n454 256.663
R606 B.n586 B.n454 256.663
R607 B.n592 B.n454 256.663
R608 B.n594 B.n454 256.663
R609 B.n600 B.n454 256.663
R610 B.n602 B.n454 256.663
R611 B.n608 B.n454 256.663
R612 B.n610 B.n454 256.663
R613 B.n616 B.n454 256.663
R614 B.n618 B.n454 256.663
R615 B.n624 B.n454 256.663
R616 B.n626 B.n454 256.663
R617 B.n632 B.n454 256.663
R618 B.n634 B.n454 256.663
R619 B.n640 B.n454 256.663
R620 B.n642 B.n454 256.663
R621 B.n648 B.n454 256.663
R622 B.n650 B.n454 256.663
R623 B.n657 B.n454 256.663
R624 B.n659 B.n454 256.663
R625 B.n665 B.n454 256.663
R626 B.n667 B.n454 256.663
R627 B.n676 B.n454 256.663
R628 B.n678 B.n454 256.663
R629 B.n684 B.n454 256.663
R630 B.n686 B.n454 256.663
R631 B.n692 B.n454 256.663
R632 B.n694 B.n454 256.663
R633 B.n700 B.n454 256.663
R634 B.n702 B.n454 256.663
R635 B.n708 B.n454 256.663
R636 B.n710 B.n454 256.663
R637 B.n716 B.n454 256.663
R638 B.n718 B.n454 256.663
R639 B.n724 B.n454 256.663
R640 B.n726 B.n454 256.663
R641 B.n732 B.n454 256.663
R642 B.n734 B.n454 256.663
R643 B.n740 B.n454 256.663
R644 B.n742 B.n454 256.663
R645 B.n748 B.n454 256.663
R646 B.n750 B.n454 256.663
R647 B.n756 B.n454 256.663
R648 B.n758 B.n454 256.663
R649 B.n764 B.n454 256.663
R650 B.n766 B.n454 256.663
R651 B.n772 B.n454 256.663
R652 B.n774 B.n454 256.663
R653 B.n780 B.n454 256.663
R654 B.n782 B.n454 256.663
R655 B.n788 B.n454 256.663
R656 B.n790 B.n454 256.663
R657 B.n796 B.n454 256.663
R658 B.n799 B.n454 256.663
R659 B.n806 B.n451 163.367
R660 B.n810 B.n451 163.367
R661 B.n810 B.n445 163.367
R662 B.n818 B.n445 163.367
R663 B.n818 B.n443 163.367
R664 B.n822 B.n443 163.367
R665 B.n822 B.n437 163.367
R666 B.n830 B.n437 163.367
R667 B.n830 B.n435 163.367
R668 B.n834 B.n435 163.367
R669 B.n834 B.n429 163.367
R670 B.n842 B.n429 163.367
R671 B.n842 B.n427 163.367
R672 B.n846 B.n427 163.367
R673 B.n846 B.n421 163.367
R674 B.n854 B.n421 163.367
R675 B.n854 B.n419 163.367
R676 B.n858 B.n419 163.367
R677 B.n858 B.n413 163.367
R678 B.n867 B.n413 163.367
R679 B.n867 B.n411 163.367
R680 B.n871 B.n411 163.367
R681 B.n871 B.n406 163.367
R682 B.n880 B.n406 163.367
R683 B.n880 B.n404 163.367
R684 B.n884 B.n404 163.367
R685 B.n884 B.n2 163.367
R686 B.n986 B.n2 163.367
R687 B.n986 B.n3 163.367
R688 B.n982 B.n3 163.367
R689 B.n982 B.n9 163.367
R690 B.n978 B.n9 163.367
R691 B.n978 B.n11 163.367
R692 B.n974 B.n11 163.367
R693 B.n974 B.n15 163.367
R694 B.n970 B.n15 163.367
R695 B.n970 B.n17 163.367
R696 B.n966 B.n17 163.367
R697 B.n966 B.n23 163.367
R698 B.n962 B.n23 163.367
R699 B.n962 B.n25 163.367
R700 B.n958 B.n25 163.367
R701 B.n958 B.n30 163.367
R702 B.n954 B.n30 163.367
R703 B.n954 B.n32 163.367
R704 B.n950 B.n32 163.367
R705 B.n950 B.n37 163.367
R706 B.n946 B.n37 163.367
R707 B.n946 B.n39 163.367
R708 B.n942 B.n39 163.367
R709 B.n942 B.n44 163.367
R710 B.n938 B.n44 163.367
R711 B.n938 B.n46 163.367
R712 B.n934 B.n46 163.367
R713 B.n934 B.n51 163.367
R714 B.n930 B.n51 163.367
R715 B.n529 B.n528 163.367
R716 B.n531 B.n529 163.367
R717 B.n535 B.n524 163.367
R718 B.n539 B.n537 163.367
R719 B.n543 B.n522 163.367
R720 B.n547 B.n545 163.367
R721 B.n551 B.n520 163.367
R722 B.n555 B.n553 163.367
R723 B.n559 B.n518 163.367
R724 B.n563 B.n561 163.367
R725 B.n567 B.n516 163.367
R726 B.n571 B.n569 163.367
R727 B.n575 B.n514 163.367
R728 B.n579 B.n577 163.367
R729 B.n583 B.n512 163.367
R730 B.n587 B.n585 163.367
R731 B.n591 B.n510 163.367
R732 B.n595 B.n593 163.367
R733 B.n599 B.n508 163.367
R734 B.n603 B.n601 163.367
R735 B.n607 B.n506 163.367
R736 B.n611 B.n609 163.367
R737 B.n615 B.n504 163.367
R738 B.n619 B.n617 163.367
R739 B.n623 B.n502 163.367
R740 B.n627 B.n625 163.367
R741 B.n631 B.n500 163.367
R742 B.n635 B.n633 163.367
R743 B.n639 B.n498 163.367
R744 B.n643 B.n641 163.367
R745 B.n647 B.n496 163.367
R746 B.n651 B.n649 163.367
R747 B.n656 B.n492 163.367
R748 B.n660 B.n658 163.367
R749 B.n664 B.n490 163.367
R750 B.n668 B.n666 163.367
R751 B.n675 B.n488 163.367
R752 B.n679 B.n677 163.367
R753 B.n683 B.n486 163.367
R754 B.n687 B.n685 163.367
R755 B.n691 B.n484 163.367
R756 B.n695 B.n693 163.367
R757 B.n699 B.n482 163.367
R758 B.n703 B.n701 163.367
R759 B.n707 B.n480 163.367
R760 B.n711 B.n709 163.367
R761 B.n715 B.n478 163.367
R762 B.n719 B.n717 163.367
R763 B.n723 B.n476 163.367
R764 B.n727 B.n725 163.367
R765 B.n731 B.n474 163.367
R766 B.n735 B.n733 163.367
R767 B.n739 B.n472 163.367
R768 B.n743 B.n741 163.367
R769 B.n747 B.n470 163.367
R770 B.n751 B.n749 163.367
R771 B.n755 B.n468 163.367
R772 B.n759 B.n757 163.367
R773 B.n763 B.n466 163.367
R774 B.n767 B.n765 163.367
R775 B.n771 B.n464 163.367
R776 B.n775 B.n773 163.367
R777 B.n779 B.n462 163.367
R778 B.n783 B.n781 163.367
R779 B.n787 B.n460 163.367
R780 B.n791 B.n789 163.367
R781 B.n795 B.n458 163.367
R782 B.n798 B.n797 163.367
R783 B.n800 B.n455 163.367
R784 B.n804 B.n449 163.367
R785 B.n812 B.n449 163.367
R786 B.n812 B.n447 163.367
R787 B.n816 B.n447 163.367
R788 B.n816 B.n441 163.367
R789 B.n824 B.n441 163.367
R790 B.n824 B.n439 163.367
R791 B.n828 B.n439 163.367
R792 B.n828 B.n433 163.367
R793 B.n836 B.n433 163.367
R794 B.n836 B.n431 163.367
R795 B.n840 B.n431 163.367
R796 B.n840 B.n425 163.367
R797 B.n848 B.n425 163.367
R798 B.n848 B.n423 163.367
R799 B.n852 B.n423 163.367
R800 B.n852 B.n417 163.367
R801 B.n860 B.n417 163.367
R802 B.n860 B.n415 163.367
R803 B.n864 B.n415 163.367
R804 B.n864 B.n410 163.367
R805 B.n873 B.n410 163.367
R806 B.n873 B.n408 163.367
R807 B.n878 B.n408 163.367
R808 B.n878 B.n402 163.367
R809 B.n886 B.n402 163.367
R810 B.n887 B.n886 163.367
R811 B.n887 B.n5 163.367
R812 B.n6 B.n5 163.367
R813 B.n7 B.n6 163.367
R814 B.n892 B.n7 163.367
R815 B.n892 B.n12 163.367
R816 B.n13 B.n12 163.367
R817 B.n14 B.n13 163.367
R818 B.n897 B.n14 163.367
R819 B.n897 B.n19 163.367
R820 B.n20 B.n19 163.367
R821 B.n21 B.n20 163.367
R822 B.n902 B.n21 163.367
R823 B.n902 B.n26 163.367
R824 B.n27 B.n26 163.367
R825 B.n28 B.n27 163.367
R826 B.n907 B.n28 163.367
R827 B.n907 B.n33 163.367
R828 B.n34 B.n33 163.367
R829 B.n35 B.n34 163.367
R830 B.n912 B.n35 163.367
R831 B.n912 B.n40 163.367
R832 B.n41 B.n40 163.367
R833 B.n42 B.n41 163.367
R834 B.n917 B.n42 163.367
R835 B.n917 B.n47 163.367
R836 B.n48 B.n47 163.367
R837 B.n49 B.n48 163.367
R838 B.n922 B.n49 163.367
R839 B.n922 B.n54 163.367
R840 B.n132 B.n131 163.367
R841 B.n136 B.n135 163.367
R842 B.n140 B.n139 163.367
R843 B.n144 B.n143 163.367
R844 B.n148 B.n147 163.367
R845 B.n152 B.n151 163.367
R846 B.n156 B.n155 163.367
R847 B.n160 B.n159 163.367
R848 B.n164 B.n163 163.367
R849 B.n168 B.n167 163.367
R850 B.n172 B.n171 163.367
R851 B.n176 B.n175 163.367
R852 B.n180 B.n179 163.367
R853 B.n184 B.n183 163.367
R854 B.n188 B.n187 163.367
R855 B.n192 B.n191 163.367
R856 B.n196 B.n195 163.367
R857 B.n200 B.n199 163.367
R858 B.n204 B.n203 163.367
R859 B.n208 B.n207 163.367
R860 B.n212 B.n211 163.367
R861 B.n216 B.n215 163.367
R862 B.n220 B.n219 163.367
R863 B.n224 B.n223 163.367
R864 B.n228 B.n227 163.367
R865 B.n232 B.n231 163.367
R866 B.n236 B.n235 163.367
R867 B.n240 B.n239 163.367
R868 B.n244 B.n243 163.367
R869 B.n248 B.n247 163.367
R870 B.n252 B.n251 163.367
R871 B.n256 B.n255 163.367
R872 B.n260 B.n259 163.367
R873 B.n264 B.n263 163.367
R874 B.n268 B.n267 163.367
R875 B.n272 B.n271 163.367
R876 B.n276 B.n275 163.367
R877 B.n280 B.n279 163.367
R878 B.n284 B.n283 163.367
R879 B.n288 B.n287 163.367
R880 B.n292 B.n291 163.367
R881 B.n296 B.n295 163.367
R882 B.n300 B.n299 163.367
R883 B.n304 B.n303 163.367
R884 B.n308 B.n307 163.367
R885 B.n312 B.n311 163.367
R886 B.n316 B.n315 163.367
R887 B.n320 B.n319 163.367
R888 B.n324 B.n323 163.367
R889 B.n328 B.n327 163.367
R890 B.n332 B.n331 163.367
R891 B.n336 B.n335 163.367
R892 B.n340 B.n339 163.367
R893 B.n344 B.n343 163.367
R894 B.n348 B.n347 163.367
R895 B.n352 B.n351 163.367
R896 B.n356 B.n355 163.367
R897 B.n360 B.n359 163.367
R898 B.n364 B.n363 163.367
R899 B.n368 B.n367 163.367
R900 B.n372 B.n371 163.367
R901 B.n376 B.n375 163.367
R902 B.n380 B.n379 163.367
R903 B.n384 B.n383 163.367
R904 B.n388 B.n387 163.367
R905 B.n392 B.n391 163.367
R906 B.n396 B.n395 163.367
R907 B.n398 B.n123 163.367
R908 B.n527 B.n453 71.676
R909 B.n531 B.n530 71.676
R910 B.n536 B.n535 71.676
R911 B.n539 B.n538 71.676
R912 B.n544 B.n543 71.676
R913 B.n547 B.n546 71.676
R914 B.n552 B.n551 71.676
R915 B.n555 B.n554 71.676
R916 B.n560 B.n559 71.676
R917 B.n563 B.n562 71.676
R918 B.n568 B.n567 71.676
R919 B.n571 B.n570 71.676
R920 B.n576 B.n575 71.676
R921 B.n579 B.n578 71.676
R922 B.n584 B.n583 71.676
R923 B.n587 B.n586 71.676
R924 B.n592 B.n591 71.676
R925 B.n595 B.n594 71.676
R926 B.n600 B.n599 71.676
R927 B.n603 B.n602 71.676
R928 B.n608 B.n607 71.676
R929 B.n611 B.n610 71.676
R930 B.n616 B.n615 71.676
R931 B.n619 B.n618 71.676
R932 B.n624 B.n623 71.676
R933 B.n627 B.n626 71.676
R934 B.n632 B.n631 71.676
R935 B.n635 B.n634 71.676
R936 B.n640 B.n639 71.676
R937 B.n643 B.n642 71.676
R938 B.n648 B.n647 71.676
R939 B.n651 B.n650 71.676
R940 B.n657 B.n656 71.676
R941 B.n660 B.n659 71.676
R942 B.n665 B.n664 71.676
R943 B.n668 B.n667 71.676
R944 B.n676 B.n675 71.676
R945 B.n679 B.n678 71.676
R946 B.n684 B.n683 71.676
R947 B.n687 B.n686 71.676
R948 B.n692 B.n691 71.676
R949 B.n695 B.n694 71.676
R950 B.n700 B.n699 71.676
R951 B.n703 B.n702 71.676
R952 B.n708 B.n707 71.676
R953 B.n711 B.n710 71.676
R954 B.n716 B.n715 71.676
R955 B.n719 B.n718 71.676
R956 B.n724 B.n723 71.676
R957 B.n727 B.n726 71.676
R958 B.n732 B.n731 71.676
R959 B.n735 B.n734 71.676
R960 B.n740 B.n739 71.676
R961 B.n743 B.n742 71.676
R962 B.n748 B.n747 71.676
R963 B.n751 B.n750 71.676
R964 B.n756 B.n755 71.676
R965 B.n759 B.n758 71.676
R966 B.n764 B.n763 71.676
R967 B.n767 B.n766 71.676
R968 B.n772 B.n771 71.676
R969 B.n775 B.n774 71.676
R970 B.n780 B.n779 71.676
R971 B.n783 B.n782 71.676
R972 B.n788 B.n787 71.676
R973 B.n791 B.n790 71.676
R974 B.n796 B.n795 71.676
R975 B.n799 B.n798 71.676
R976 B.n55 B.n53 71.676
R977 B.n132 B.n56 71.676
R978 B.n136 B.n57 71.676
R979 B.n140 B.n58 71.676
R980 B.n144 B.n59 71.676
R981 B.n148 B.n60 71.676
R982 B.n152 B.n61 71.676
R983 B.n156 B.n62 71.676
R984 B.n160 B.n63 71.676
R985 B.n164 B.n64 71.676
R986 B.n168 B.n65 71.676
R987 B.n172 B.n66 71.676
R988 B.n176 B.n67 71.676
R989 B.n180 B.n68 71.676
R990 B.n184 B.n69 71.676
R991 B.n188 B.n70 71.676
R992 B.n192 B.n71 71.676
R993 B.n196 B.n72 71.676
R994 B.n200 B.n73 71.676
R995 B.n204 B.n74 71.676
R996 B.n208 B.n75 71.676
R997 B.n212 B.n76 71.676
R998 B.n216 B.n77 71.676
R999 B.n220 B.n78 71.676
R1000 B.n224 B.n79 71.676
R1001 B.n228 B.n80 71.676
R1002 B.n232 B.n81 71.676
R1003 B.n236 B.n82 71.676
R1004 B.n240 B.n83 71.676
R1005 B.n244 B.n84 71.676
R1006 B.n248 B.n85 71.676
R1007 B.n252 B.n86 71.676
R1008 B.n256 B.n87 71.676
R1009 B.n260 B.n88 71.676
R1010 B.n264 B.n89 71.676
R1011 B.n268 B.n90 71.676
R1012 B.n272 B.n91 71.676
R1013 B.n276 B.n92 71.676
R1014 B.n280 B.n93 71.676
R1015 B.n284 B.n94 71.676
R1016 B.n288 B.n95 71.676
R1017 B.n292 B.n96 71.676
R1018 B.n296 B.n97 71.676
R1019 B.n300 B.n98 71.676
R1020 B.n304 B.n99 71.676
R1021 B.n308 B.n100 71.676
R1022 B.n312 B.n101 71.676
R1023 B.n316 B.n102 71.676
R1024 B.n320 B.n103 71.676
R1025 B.n324 B.n104 71.676
R1026 B.n328 B.n105 71.676
R1027 B.n332 B.n106 71.676
R1028 B.n336 B.n107 71.676
R1029 B.n340 B.n108 71.676
R1030 B.n344 B.n109 71.676
R1031 B.n348 B.n110 71.676
R1032 B.n352 B.n111 71.676
R1033 B.n356 B.n112 71.676
R1034 B.n360 B.n113 71.676
R1035 B.n364 B.n114 71.676
R1036 B.n368 B.n115 71.676
R1037 B.n372 B.n116 71.676
R1038 B.n376 B.n117 71.676
R1039 B.n380 B.n118 71.676
R1040 B.n384 B.n119 71.676
R1041 B.n388 B.n120 71.676
R1042 B.n392 B.n121 71.676
R1043 B.n396 B.n122 71.676
R1044 B.n927 B.n123 71.676
R1045 B.n927 B.n926 71.676
R1046 B.n398 B.n122 71.676
R1047 B.n395 B.n121 71.676
R1048 B.n391 B.n120 71.676
R1049 B.n387 B.n119 71.676
R1050 B.n383 B.n118 71.676
R1051 B.n379 B.n117 71.676
R1052 B.n375 B.n116 71.676
R1053 B.n371 B.n115 71.676
R1054 B.n367 B.n114 71.676
R1055 B.n363 B.n113 71.676
R1056 B.n359 B.n112 71.676
R1057 B.n355 B.n111 71.676
R1058 B.n351 B.n110 71.676
R1059 B.n347 B.n109 71.676
R1060 B.n343 B.n108 71.676
R1061 B.n339 B.n107 71.676
R1062 B.n335 B.n106 71.676
R1063 B.n331 B.n105 71.676
R1064 B.n327 B.n104 71.676
R1065 B.n323 B.n103 71.676
R1066 B.n319 B.n102 71.676
R1067 B.n315 B.n101 71.676
R1068 B.n311 B.n100 71.676
R1069 B.n307 B.n99 71.676
R1070 B.n303 B.n98 71.676
R1071 B.n299 B.n97 71.676
R1072 B.n295 B.n96 71.676
R1073 B.n291 B.n95 71.676
R1074 B.n287 B.n94 71.676
R1075 B.n283 B.n93 71.676
R1076 B.n279 B.n92 71.676
R1077 B.n275 B.n91 71.676
R1078 B.n271 B.n90 71.676
R1079 B.n267 B.n89 71.676
R1080 B.n263 B.n88 71.676
R1081 B.n259 B.n87 71.676
R1082 B.n255 B.n86 71.676
R1083 B.n251 B.n85 71.676
R1084 B.n247 B.n84 71.676
R1085 B.n243 B.n83 71.676
R1086 B.n239 B.n82 71.676
R1087 B.n235 B.n81 71.676
R1088 B.n231 B.n80 71.676
R1089 B.n227 B.n79 71.676
R1090 B.n223 B.n78 71.676
R1091 B.n219 B.n77 71.676
R1092 B.n215 B.n76 71.676
R1093 B.n211 B.n75 71.676
R1094 B.n207 B.n74 71.676
R1095 B.n203 B.n73 71.676
R1096 B.n199 B.n72 71.676
R1097 B.n195 B.n71 71.676
R1098 B.n191 B.n70 71.676
R1099 B.n187 B.n69 71.676
R1100 B.n183 B.n68 71.676
R1101 B.n179 B.n67 71.676
R1102 B.n175 B.n66 71.676
R1103 B.n171 B.n65 71.676
R1104 B.n167 B.n64 71.676
R1105 B.n163 B.n63 71.676
R1106 B.n159 B.n62 71.676
R1107 B.n155 B.n61 71.676
R1108 B.n151 B.n60 71.676
R1109 B.n147 B.n59 71.676
R1110 B.n143 B.n58 71.676
R1111 B.n139 B.n57 71.676
R1112 B.n135 B.n56 71.676
R1113 B.n131 B.n55 71.676
R1114 B.n528 B.n527 71.676
R1115 B.n530 B.n524 71.676
R1116 B.n537 B.n536 71.676
R1117 B.n538 B.n522 71.676
R1118 B.n545 B.n544 71.676
R1119 B.n546 B.n520 71.676
R1120 B.n553 B.n552 71.676
R1121 B.n554 B.n518 71.676
R1122 B.n561 B.n560 71.676
R1123 B.n562 B.n516 71.676
R1124 B.n569 B.n568 71.676
R1125 B.n570 B.n514 71.676
R1126 B.n577 B.n576 71.676
R1127 B.n578 B.n512 71.676
R1128 B.n585 B.n584 71.676
R1129 B.n586 B.n510 71.676
R1130 B.n593 B.n592 71.676
R1131 B.n594 B.n508 71.676
R1132 B.n601 B.n600 71.676
R1133 B.n602 B.n506 71.676
R1134 B.n609 B.n608 71.676
R1135 B.n610 B.n504 71.676
R1136 B.n617 B.n616 71.676
R1137 B.n618 B.n502 71.676
R1138 B.n625 B.n624 71.676
R1139 B.n626 B.n500 71.676
R1140 B.n633 B.n632 71.676
R1141 B.n634 B.n498 71.676
R1142 B.n641 B.n640 71.676
R1143 B.n642 B.n496 71.676
R1144 B.n649 B.n648 71.676
R1145 B.n650 B.n492 71.676
R1146 B.n658 B.n657 71.676
R1147 B.n659 B.n490 71.676
R1148 B.n666 B.n665 71.676
R1149 B.n667 B.n488 71.676
R1150 B.n677 B.n676 71.676
R1151 B.n678 B.n486 71.676
R1152 B.n685 B.n684 71.676
R1153 B.n686 B.n484 71.676
R1154 B.n693 B.n692 71.676
R1155 B.n694 B.n482 71.676
R1156 B.n701 B.n700 71.676
R1157 B.n702 B.n480 71.676
R1158 B.n709 B.n708 71.676
R1159 B.n710 B.n478 71.676
R1160 B.n717 B.n716 71.676
R1161 B.n718 B.n476 71.676
R1162 B.n725 B.n724 71.676
R1163 B.n726 B.n474 71.676
R1164 B.n733 B.n732 71.676
R1165 B.n734 B.n472 71.676
R1166 B.n741 B.n740 71.676
R1167 B.n742 B.n470 71.676
R1168 B.n749 B.n748 71.676
R1169 B.n750 B.n468 71.676
R1170 B.n757 B.n756 71.676
R1171 B.n758 B.n466 71.676
R1172 B.n765 B.n764 71.676
R1173 B.n766 B.n464 71.676
R1174 B.n773 B.n772 71.676
R1175 B.n774 B.n462 71.676
R1176 B.n781 B.n780 71.676
R1177 B.n782 B.n460 71.676
R1178 B.n789 B.n788 71.676
R1179 B.n790 B.n458 71.676
R1180 B.n797 B.n796 71.676
R1181 B.n800 B.n799 71.676
R1182 B.n672 B.n671 65.746
R1183 B.n494 B.n493 65.746
R1184 B.n128 B.n127 65.746
R1185 B.n125 B.n124 65.746
R1186 B.n673 B.n672 59.5399
R1187 B.n653 B.n494 59.5399
R1188 B.n129 B.n128 59.5399
R1189 B.n126 B.n125 59.5399
R1190 B.n805 B.n454 55.9364
R1191 B.n929 B.n928 55.9364
R1192 B.n931 B.n52 33.5615
R1193 B.n925 B.n924 33.5615
R1194 B.n803 B.n802 33.5615
R1195 B.n807 B.n452 33.5615
R1196 B.n805 B.n450 29.9504
R1197 B.n811 B.n450 29.9504
R1198 B.n811 B.n446 29.9504
R1199 B.n817 B.n446 29.9504
R1200 B.n817 B.n442 29.9504
R1201 B.n823 B.n442 29.9504
R1202 B.n823 B.n438 29.9504
R1203 B.n829 B.n438 29.9504
R1204 B.n835 B.n434 29.9504
R1205 B.n835 B.n430 29.9504
R1206 B.n841 B.n430 29.9504
R1207 B.n841 B.n426 29.9504
R1208 B.n847 B.n426 29.9504
R1209 B.n847 B.n422 29.9504
R1210 B.n853 B.n422 29.9504
R1211 B.n853 B.n418 29.9504
R1212 B.n859 B.n418 29.9504
R1213 B.n859 B.n414 29.9504
R1214 B.n866 B.n414 29.9504
R1215 B.n866 B.n865 29.9504
R1216 B.n872 B.n407 29.9504
R1217 B.n879 B.n407 29.9504
R1218 B.n879 B.n403 29.9504
R1219 B.n885 B.n403 29.9504
R1220 B.n885 B.n4 29.9504
R1221 B.n985 B.n4 29.9504
R1222 B.n985 B.n984 29.9504
R1223 B.n984 B.n983 29.9504
R1224 B.n983 B.n8 29.9504
R1225 B.n977 B.n8 29.9504
R1226 B.n977 B.n976 29.9504
R1227 B.n976 B.n975 29.9504
R1228 B.n969 B.n18 29.9504
R1229 B.n969 B.n968 29.9504
R1230 B.n968 B.n967 29.9504
R1231 B.n967 B.n22 29.9504
R1232 B.n961 B.n22 29.9504
R1233 B.n961 B.n960 29.9504
R1234 B.n960 B.n959 29.9504
R1235 B.n959 B.n29 29.9504
R1236 B.n953 B.n29 29.9504
R1237 B.n953 B.n952 29.9504
R1238 B.n952 B.n951 29.9504
R1239 B.n951 B.n36 29.9504
R1240 B.n945 B.n944 29.9504
R1241 B.n944 B.n943 29.9504
R1242 B.n943 B.n43 29.9504
R1243 B.n937 B.n43 29.9504
R1244 B.n937 B.n936 29.9504
R1245 B.n936 B.n935 29.9504
R1246 B.n935 B.n50 29.9504
R1247 B.n929 B.n50 29.9504
R1248 B.t10 B.n434 22.9034
R1249 B.t3 B.n36 22.9034
R1250 B B.n987 18.0485
R1251 B.n872 B.t1 17.6181
R1252 B.n975 B.t0 17.6181
R1253 B.n865 B.t1 12.3328
R1254 B.n18 B.t0 12.3328
R1255 B.n130 B.n52 10.6151
R1256 B.n133 B.n130 10.6151
R1257 B.n134 B.n133 10.6151
R1258 B.n137 B.n134 10.6151
R1259 B.n138 B.n137 10.6151
R1260 B.n141 B.n138 10.6151
R1261 B.n142 B.n141 10.6151
R1262 B.n145 B.n142 10.6151
R1263 B.n146 B.n145 10.6151
R1264 B.n149 B.n146 10.6151
R1265 B.n150 B.n149 10.6151
R1266 B.n153 B.n150 10.6151
R1267 B.n154 B.n153 10.6151
R1268 B.n157 B.n154 10.6151
R1269 B.n158 B.n157 10.6151
R1270 B.n161 B.n158 10.6151
R1271 B.n162 B.n161 10.6151
R1272 B.n165 B.n162 10.6151
R1273 B.n166 B.n165 10.6151
R1274 B.n169 B.n166 10.6151
R1275 B.n170 B.n169 10.6151
R1276 B.n173 B.n170 10.6151
R1277 B.n174 B.n173 10.6151
R1278 B.n177 B.n174 10.6151
R1279 B.n178 B.n177 10.6151
R1280 B.n181 B.n178 10.6151
R1281 B.n182 B.n181 10.6151
R1282 B.n185 B.n182 10.6151
R1283 B.n186 B.n185 10.6151
R1284 B.n189 B.n186 10.6151
R1285 B.n190 B.n189 10.6151
R1286 B.n193 B.n190 10.6151
R1287 B.n194 B.n193 10.6151
R1288 B.n197 B.n194 10.6151
R1289 B.n198 B.n197 10.6151
R1290 B.n201 B.n198 10.6151
R1291 B.n202 B.n201 10.6151
R1292 B.n205 B.n202 10.6151
R1293 B.n206 B.n205 10.6151
R1294 B.n209 B.n206 10.6151
R1295 B.n210 B.n209 10.6151
R1296 B.n213 B.n210 10.6151
R1297 B.n214 B.n213 10.6151
R1298 B.n217 B.n214 10.6151
R1299 B.n218 B.n217 10.6151
R1300 B.n221 B.n218 10.6151
R1301 B.n222 B.n221 10.6151
R1302 B.n225 B.n222 10.6151
R1303 B.n226 B.n225 10.6151
R1304 B.n229 B.n226 10.6151
R1305 B.n230 B.n229 10.6151
R1306 B.n233 B.n230 10.6151
R1307 B.n234 B.n233 10.6151
R1308 B.n237 B.n234 10.6151
R1309 B.n238 B.n237 10.6151
R1310 B.n241 B.n238 10.6151
R1311 B.n242 B.n241 10.6151
R1312 B.n245 B.n242 10.6151
R1313 B.n246 B.n245 10.6151
R1314 B.n249 B.n246 10.6151
R1315 B.n250 B.n249 10.6151
R1316 B.n253 B.n250 10.6151
R1317 B.n254 B.n253 10.6151
R1318 B.n258 B.n257 10.6151
R1319 B.n261 B.n258 10.6151
R1320 B.n262 B.n261 10.6151
R1321 B.n265 B.n262 10.6151
R1322 B.n266 B.n265 10.6151
R1323 B.n269 B.n266 10.6151
R1324 B.n270 B.n269 10.6151
R1325 B.n273 B.n270 10.6151
R1326 B.n274 B.n273 10.6151
R1327 B.n278 B.n277 10.6151
R1328 B.n281 B.n278 10.6151
R1329 B.n282 B.n281 10.6151
R1330 B.n285 B.n282 10.6151
R1331 B.n286 B.n285 10.6151
R1332 B.n289 B.n286 10.6151
R1333 B.n290 B.n289 10.6151
R1334 B.n293 B.n290 10.6151
R1335 B.n294 B.n293 10.6151
R1336 B.n297 B.n294 10.6151
R1337 B.n298 B.n297 10.6151
R1338 B.n301 B.n298 10.6151
R1339 B.n302 B.n301 10.6151
R1340 B.n305 B.n302 10.6151
R1341 B.n306 B.n305 10.6151
R1342 B.n309 B.n306 10.6151
R1343 B.n310 B.n309 10.6151
R1344 B.n313 B.n310 10.6151
R1345 B.n314 B.n313 10.6151
R1346 B.n317 B.n314 10.6151
R1347 B.n318 B.n317 10.6151
R1348 B.n321 B.n318 10.6151
R1349 B.n322 B.n321 10.6151
R1350 B.n325 B.n322 10.6151
R1351 B.n326 B.n325 10.6151
R1352 B.n329 B.n326 10.6151
R1353 B.n330 B.n329 10.6151
R1354 B.n333 B.n330 10.6151
R1355 B.n334 B.n333 10.6151
R1356 B.n337 B.n334 10.6151
R1357 B.n338 B.n337 10.6151
R1358 B.n341 B.n338 10.6151
R1359 B.n342 B.n341 10.6151
R1360 B.n345 B.n342 10.6151
R1361 B.n346 B.n345 10.6151
R1362 B.n349 B.n346 10.6151
R1363 B.n350 B.n349 10.6151
R1364 B.n353 B.n350 10.6151
R1365 B.n354 B.n353 10.6151
R1366 B.n357 B.n354 10.6151
R1367 B.n358 B.n357 10.6151
R1368 B.n361 B.n358 10.6151
R1369 B.n362 B.n361 10.6151
R1370 B.n365 B.n362 10.6151
R1371 B.n366 B.n365 10.6151
R1372 B.n369 B.n366 10.6151
R1373 B.n370 B.n369 10.6151
R1374 B.n373 B.n370 10.6151
R1375 B.n374 B.n373 10.6151
R1376 B.n377 B.n374 10.6151
R1377 B.n378 B.n377 10.6151
R1378 B.n381 B.n378 10.6151
R1379 B.n382 B.n381 10.6151
R1380 B.n385 B.n382 10.6151
R1381 B.n386 B.n385 10.6151
R1382 B.n389 B.n386 10.6151
R1383 B.n390 B.n389 10.6151
R1384 B.n393 B.n390 10.6151
R1385 B.n394 B.n393 10.6151
R1386 B.n397 B.n394 10.6151
R1387 B.n399 B.n397 10.6151
R1388 B.n400 B.n399 10.6151
R1389 B.n925 B.n400 10.6151
R1390 B.n803 B.n448 10.6151
R1391 B.n813 B.n448 10.6151
R1392 B.n814 B.n813 10.6151
R1393 B.n815 B.n814 10.6151
R1394 B.n815 B.n440 10.6151
R1395 B.n825 B.n440 10.6151
R1396 B.n826 B.n825 10.6151
R1397 B.n827 B.n826 10.6151
R1398 B.n827 B.n432 10.6151
R1399 B.n837 B.n432 10.6151
R1400 B.n838 B.n837 10.6151
R1401 B.n839 B.n838 10.6151
R1402 B.n839 B.n424 10.6151
R1403 B.n849 B.n424 10.6151
R1404 B.n850 B.n849 10.6151
R1405 B.n851 B.n850 10.6151
R1406 B.n851 B.n416 10.6151
R1407 B.n861 B.n416 10.6151
R1408 B.n862 B.n861 10.6151
R1409 B.n863 B.n862 10.6151
R1410 B.n863 B.n409 10.6151
R1411 B.n874 B.n409 10.6151
R1412 B.n875 B.n874 10.6151
R1413 B.n877 B.n875 10.6151
R1414 B.n877 B.n876 10.6151
R1415 B.n876 B.n401 10.6151
R1416 B.n888 B.n401 10.6151
R1417 B.n889 B.n888 10.6151
R1418 B.n890 B.n889 10.6151
R1419 B.n891 B.n890 10.6151
R1420 B.n893 B.n891 10.6151
R1421 B.n894 B.n893 10.6151
R1422 B.n895 B.n894 10.6151
R1423 B.n896 B.n895 10.6151
R1424 B.n898 B.n896 10.6151
R1425 B.n899 B.n898 10.6151
R1426 B.n900 B.n899 10.6151
R1427 B.n901 B.n900 10.6151
R1428 B.n903 B.n901 10.6151
R1429 B.n904 B.n903 10.6151
R1430 B.n905 B.n904 10.6151
R1431 B.n906 B.n905 10.6151
R1432 B.n908 B.n906 10.6151
R1433 B.n909 B.n908 10.6151
R1434 B.n910 B.n909 10.6151
R1435 B.n911 B.n910 10.6151
R1436 B.n913 B.n911 10.6151
R1437 B.n914 B.n913 10.6151
R1438 B.n915 B.n914 10.6151
R1439 B.n916 B.n915 10.6151
R1440 B.n918 B.n916 10.6151
R1441 B.n919 B.n918 10.6151
R1442 B.n920 B.n919 10.6151
R1443 B.n921 B.n920 10.6151
R1444 B.n923 B.n921 10.6151
R1445 B.n924 B.n923 10.6151
R1446 B.n526 B.n452 10.6151
R1447 B.n526 B.n525 10.6151
R1448 B.n532 B.n525 10.6151
R1449 B.n533 B.n532 10.6151
R1450 B.n534 B.n533 10.6151
R1451 B.n534 B.n523 10.6151
R1452 B.n540 B.n523 10.6151
R1453 B.n541 B.n540 10.6151
R1454 B.n542 B.n541 10.6151
R1455 B.n542 B.n521 10.6151
R1456 B.n548 B.n521 10.6151
R1457 B.n549 B.n548 10.6151
R1458 B.n550 B.n549 10.6151
R1459 B.n550 B.n519 10.6151
R1460 B.n556 B.n519 10.6151
R1461 B.n557 B.n556 10.6151
R1462 B.n558 B.n557 10.6151
R1463 B.n558 B.n517 10.6151
R1464 B.n564 B.n517 10.6151
R1465 B.n565 B.n564 10.6151
R1466 B.n566 B.n565 10.6151
R1467 B.n566 B.n515 10.6151
R1468 B.n572 B.n515 10.6151
R1469 B.n573 B.n572 10.6151
R1470 B.n574 B.n573 10.6151
R1471 B.n574 B.n513 10.6151
R1472 B.n580 B.n513 10.6151
R1473 B.n581 B.n580 10.6151
R1474 B.n582 B.n581 10.6151
R1475 B.n582 B.n511 10.6151
R1476 B.n588 B.n511 10.6151
R1477 B.n589 B.n588 10.6151
R1478 B.n590 B.n589 10.6151
R1479 B.n590 B.n509 10.6151
R1480 B.n596 B.n509 10.6151
R1481 B.n597 B.n596 10.6151
R1482 B.n598 B.n597 10.6151
R1483 B.n598 B.n507 10.6151
R1484 B.n604 B.n507 10.6151
R1485 B.n605 B.n604 10.6151
R1486 B.n606 B.n605 10.6151
R1487 B.n606 B.n505 10.6151
R1488 B.n612 B.n505 10.6151
R1489 B.n613 B.n612 10.6151
R1490 B.n614 B.n613 10.6151
R1491 B.n614 B.n503 10.6151
R1492 B.n620 B.n503 10.6151
R1493 B.n621 B.n620 10.6151
R1494 B.n622 B.n621 10.6151
R1495 B.n622 B.n501 10.6151
R1496 B.n628 B.n501 10.6151
R1497 B.n629 B.n628 10.6151
R1498 B.n630 B.n629 10.6151
R1499 B.n630 B.n499 10.6151
R1500 B.n636 B.n499 10.6151
R1501 B.n637 B.n636 10.6151
R1502 B.n638 B.n637 10.6151
R1503 B.n638 B.n497 10.6151
R1504 B.n644 B.n497 10.6151
R1505 B.n645 B.n644 10.6151
R1506 B.n646 B.n645 10.6151
R1507 B.n646 B.n495 10.6151
R1508 B.n652 B.n495 10.6151
R1509 B.n655 B.n654 10.6151
R1510 B.n655 B.n491 10.6151
R1511 B.n661 B.n491 10.6151
R1512 B.n662 B.n661 10.6151
R1513 B.n663 B.n662 10.6151
R1514 B.n663 B.n489 10.6151
R1515 B.n669 B.n489 10.6151
R1516 B.n670 B.n669 10.6151
R1517 B.n674 B.n670 10.6151
R1518 B.n680 B.n487 10.6151
R1519 B.n681 B.n680 10.6151
R1520 B.n682 B.n681 10.6151
R1521 B.n682 B.n485 10.6151
R1522 B.n688 B.n485 10.6151
R1523 B.n689 B.n688 10.6151
R1524 B.n690 B.n689 10.6151
R1525 B.n690 B.n483 10.6151
R1526 B.n696 B.n483 10.6151
R1527 B.n697 B.n696 10.6151
R1528 B.n698 B.n697 10.6151
R1529 B.n698 B.n481 10.6151
R1530 B.n704 B.n481 10.6151
R1531 B.n705 B.n704 10.6151
R1532 B.n706 B.n705 10.6151
R1533 B.n706 B.n479 10.6151
R1534 B.n712 B.n479 10.6151
R1535 B.n713 B.n712 10.6151
R1536 B.n714 B.n713 10.6151
R1537 B.n714 B.n477 10.6151
R1538 B.n720 B.n477 10.6151
R1539 B.n721 B.n720 10.6151
R1540 B.n722 B.n721 10.6151
R1541 B.n722 B.n475 10.6151
R1542 B.n728 B.n475 10.6151
R1543 B.n729 B.n728 10.6151
R1544 B.n730 B.n729 10.6151
R1545 B.n730 B.n473 10.6151
R1546 B.n736 B.n473 10.6151
R1547 B.n737 B.n736 10.6151
R1548 B.n738 B.n737 10.6151
R1549 B.n738 B.n471 10.6151
R1550 B.n744 B.n471 10.6151
R1551 B.n745 B.n744 10.6151
R1552 B.n746 B.n745 10.6151
R1553 B.n746 B.n469 10.6151
R1554 B.n752 B.n469 10.6151
R1555 B.n753 B.n752 10.6151
R1556 B.n754 B.n753 10.6151
R1557 B.n754 B.n467 10.6151
R1558 B.n760 B.n467 10.6151
R1559 B.n761 B.n760 10.6151
R1560 B.n762 B.n761 10.6151
R1561 B.n762 B.n465 10.6151
R1562 B.n768 B.n465 10.6151
R1563 B.n769 B.n768 10.6151
R1564 B.n770 B.n769 10.6151
R1565 B.n770 B.n463 10.6151
R1566 B.n776 B.n463 10.6151
R1567 B.n777 B.n776 10.6151
R1568 B.n778 B.n777 10.6151
R1569 B.n778 B.n461 10.6151
R1570 B.n784 B.n461 10.6151
R1571 B.n785 B.n784 10.6151
R1572 B.n786 B.n785 10.6151
R1573 B.n786 B.n459 10.6151
R1574 B.n792 B.n459 10.6151
R1575 B.n793 B.n792 10.6151
R1576 B.n794 B.n793 10.6151
R1577 B.n794 B.n457 10.6151
R1578 B.n457 B.n456 10.6151
R1579 B.n801 B.n456 10.6151
R1580 B.n802 B.n801 10.6151
R1581 B.n808 B.n807 10.6151
R1582 B.n809 B.n808 10.6151
R1583 B.n809 B.n444 10.6151
R1584 B.n819 B.n444 10.6151
R1585 B.n820 B.n819 10.6151
R1586 B.n821 B.n820 10.6151
R1587 B.n821 B.n436 10.6151
R1588 B.n831 B.n436 10.6151
R1589 B.n832 B.n831 10.6151
R1590 B.n833 B.n832 10.6151
R1591 B.n833 B.n428 10.6151
R1592 B.n843 B.n428 10.6151
R1593 B.n844 B.n843 10.6151
R1594 B.n845 B.n844 10.6151
R1595 B.n845 B.n420 10.6151
R1596 B.n855 B.n420 10.6151
R1597 B.n856 B.n855 10.6151
R1598 B.n857 B.n856 10.6151
R1599 B.n857 B.n412 10.6151
R1600 B.n868 B.n412 10.6151
R1601 B.n869 B.n868 10.6151
R1602 B.n870 B.n869 10.6151
R1603 B.n870 B.n405 10.6151
R1604 B.n881 B.n405 10.6151
R1605 B.n882 B.n881 10.6151
R1606 B.n883 B.n882 10.6151
R1607 B.n883 B.n0 10.6151
R1608 B.n981 B.n1 10.6151
R1609 B.n981 B.n980 10.6151
R1610 B.n980 B.n979 10.6151
R1611 B.n979 B.n10 10.6151
R1612 B.n973 B.n10 10.6151
R1613 B.n973 B.n972 10.6151
R1614 B.n972 B.n971 10.6151
R1615 B.n971 B.n16 10.6151
R1616 B.n965 B.n16 10.6151
R1617 B.n965 B.n964 10.6151
R1618 B.n964 B.n963 10.6151
R1619 B.n963 B.n24 10.6151
R1620 B.n957 B.n24 10.6151
R1621 B.n957 B.n956 10.6151
R1622 B.n956 B.n955 10.6151
R1623 B.n955 B.n31 10.6151
R1624 B.n949 B.n31 10.6151
R1625 B.n949 B.n948 10.6151
R1626 B.n948 B.n947 10.6151
R1627 B.n947 B.n38 10.6151
R1628 B.n941 B.n38 10.6151
R1629 B.n941 B.n940 10.6151
R1630 B.n940 B.n939 10.6151
R1631 B.n939 B.n45 10.6151
R1632 B.n933 B.n45 10.6151
R1633 B.n933 B.n932 10.6151
R1634 B.n932 B.n931 10.6151
R1635 B.n254 B.n129 9.36635
R1636 B.n277 B.n126 9.36635
R1637 B.n653 B.n652 9.36635
R1638 B.n673 B.n487 9.36635
R1639 B.n829 B.t10 7.04755
R1640 B.n945 B.t3 7.04755
R1641 B.n987 B.n0 2.81026
R1642 B.n987 B.n1 2.81026
R1643 B.n257 B.n129 1.24928
R1644 B.n274 B.n126 1.24928
R1645 B.n654 B.n653 1.24928
R1646 B.n674 B.n673 1.24928
R1647 VN VN.t0 248.004
R1648 VN VN.t1 196.724
R1649 VTAIL.n434 VTAIL.n330 289.615
R1650 VTAIL.n104 VTAIL.n0 289.615
R1651 VTAIL.n324 VTAIL.n220 289.615
R1652 VTAIL.n214 VTAIL.n110 289.615
R1653 VTAIL.n367 VTAIL.n366 185
R1654 VTAIL.n369 VTAIL.n368 185
R1655 VTAIL.n362 VTAIL.n361 185
R1656 VTAIL.n375 VTAIL.n374 185
R1657 VTAIL.n377 VTAIL.n376 185
R1658 VTAIL.n358 VTAIL.n357 185
R1659 VTAIL.n383 VTAIL.n382 185
R1660 VTAIL.n385 VTAIL.n384 185
R1661 VTAIL.n354 VTAIL.n353 185
R1662 VTAIL.n391 VTAIL.n390 185
R1663 VTAIL.n393 VTAIL.n392 185
R1664 VTAIL.n350 VTAIL.n349 185
R1665 VTAIL.n399 VTAIL.n398 185
R1666 VTAIL.n401 VTAIL.n400 185
R1667 VTAIL.n346 VTAIL.n345 185
R1668 VTAIL.n408 VTAIL.n407 185
R1669 VTAIL.n409 VTAIL.n344 185
R1670 VTAIL.n411 VTAIL.n410 185
R1671 VTAIL.n342 VTAIL.n341 185
R1672 VTAIL.n417 VTAIL.n416 185
R1673 VTAIL.n419 VTAIL.n418 185
R1674 VTAIL.n338 VTAIL.n337 185
R1675 VTAIL.n425 VTAIL.n424 185
R1676 VTAIL.n427 VTAIL.n426 185
R1677 VTAIL.n334 VTAIL.n333 185
R1678 VTAIL.n433 VTAIL.n432 185
R1679 VTAIL.n435 VTAIL.n434 185
R1680 VTAIL.n37 VTAIL.n36 185
R1681 VTAIL.n39 VTAIL.n38 185
R1682 VTAIL.n32 VTAIL.n31 185
R1683 VTAIL.n45 VTAIL.n44 185
R1684 VTAIL.n47 VTAIL.n46 185
R1685 VTAIL.n28 VTAIL.n27 185
R1686 VTAIL.n53 VTAIL.n52 185
R1687 VTAIL.n55 VTAIL.n54 185
R1688 VTAIL.n24 VTAIL.n23 185
R1689 VTAIL.n61 VTAIL.n60 185
R1690 VTAIL.n63 VTAIL.n62 185
R1691 VTAIL.n20 VTAIL.n19 185
R1692 VTAIL.n69 VTAIL.n68 185
R1693 VTAIL.n71 VTAIL.n70 185
R1694 VTAIL.n16 VTAIL.n15 185
R1695 VTAIL.n78 VTAIL.n77 185
R1696 VTAIL.n79 VTAIL.n14 185
R1697 VTAIL.n81 VTAIL.n80 185
R1698 VTAIL.n12 VTAIL.n11 185
R1699 VTAIL.n87 VTAIL.n86 185
R1700 VTAIL.n89 VTAIL.n88 185
R1701 VTAIL.n8 VTAIL.n7 185
R1702 VTAIL.n95 VTAIL.n94 185
R1703 VTAIL.n97 VTAIL.n96 185
R1704 VTAIL.n4 VTAIL.n3 185
R1705 VTAIL.n103 VTAIL.n102 185
R1706 VTAIL.n105 VTAIL.n104 185
R1707 VTAIL.n325 VTAIL.n324 185
R1708 VTAIL.n323 VTAIL.n322 185
R1709 VTAIL.n224 VTAIL.n223 185
R1710 VTAIL.n317 VTAIL.n316 185
R1711 VTAIL.n315 VTAIL.n314 185
R1712 VTAIL.n228 VTAIL.n227 185
R1713 VTAIL.n309 VTAIL.n308 185
R1714 VTAIL.n307 VTAIL.n306 185
R1715 VTAIL.n232 VTAIL.n231 185
R1716 VTAIL.n236 VTAIL.n234 185
R1717 VTAIL.n301 VTAIL.n300 185
R1718 VTAIL.n299 VTAIL.n298 185
R1719 VTAIL.n238 VTAIL.n237 185
R1720 VTAIL.n293 VTAIL.n292 185
R1721 VTAIL.n291 VTAIL.n290 185
R1722 VTAIL.n242 VTAIL.n241 185
R1723 VTAIL.n285 VTAIL.n284 185
R1724 VTAIL.n283 VTAIL.n282 185
R1725 VTAIL.n246 VTAIL.n245 185
R1726 VTAIL.n277 VTAIL.n276 185
R1727 VTAIL.n275 VTAIL.n274 185
R1728 VTAIL.n250 VTAIL.n249 185
R1729 VTAIL.n269 VTAIL.n268 185
R1730 VTAIL.n267 VTAIL.n266 185
R1731 VTAIL.n254 VTAIL.n253 185
R1732 VTAIL.n261 VTAIL.n260 185
R1733 VTAIL.n259 VTAIL.n258 185
R1734 VTAIL.n215 VTAIL.n214 185
R1735 VTAIL.n213 VTAIL.n212 185
R1736 VTAIL.n114 VTAIL.n113 185
R1737 VTAIL.n207 VTAIL.n206 185
R1738 VTAIL.n205 VTAIL.n204 185
R1739 VTAIL.n118 VTAIL.n117 185
R1740 VTAIL.n199 VTAIL.n198 185
R1741 VTAIL.n197 VTAIL.n196 185
R1742 VTAIL.n122 VTAIL.n121 185
R1743 VTAIL.n126 VTAIL.n124 185
R1744 VTAIL.n191 VTAIL.n190 185
R1745 VTAIL.n189 VTAIL.n188 185
R1746 VTAIL.n128 VTAIL.n127 185
R1747 VTAIL.n183 VTAIL.n182 185
R1748 VTAIL.n181 VTAIL.n180 185
R1749 VTAIL.n132 VTAIL.n131 185
R1750 VTAIL.n175 VTAIL.n174 185
R1751 VTAIL.n173 VTAIL.n172 185
R1752 VTAIL.n136 VTAIL.n135 185
R1753 VTAIL.n167 VTAIL.n166 185
R1754 VTAIL.n165 VTAIL.n164 185
R1755 VTAIL.n140 VTAIL.n139 185
R1756 VTAIL.n159 VTAIL.n158 185
R1757 VTAIL.n157 VTAIL.n156 185
R1758 VTAIL.n144 VTAIL.n143 185
R1759 VTAIL.n151 VTAIL.n150 185
R1760 VTAIL.n149 VTAIL.n148 185
R1761 VTAIL.n365 VTAIL.t3 147.659
R1762 VTAIL.n35 VTAIL.t0 147.659
R1763 VTAIL.n257 VTAIL.t1 147.659
R1764 VTAIL.n147 VTAIL.t2 147.659
R1765 VTAIL.n368 VTAIL.n367 104.615
R1766 VTAIL.n368 VTAIL.n361 104.615
R1767 VTAIL.n375 VTAIL.n361 104.615
R1768 VTAIL.n376 VTAIL.n375 104.615
R1769 VTAIL.n376 VTAIL.n357 104.615
R1770 VTAIL.n383 VTAIL.n357 104.615
R1771 VTAIL.n384 VTAIL.n383 104.615
R1772 VTAIL.n384 VTAIL.n353 104.615
R1773 VTAIL.n391 VTAIL.n353 104.615
R1774 VTAIL.n392 VTAIL.n391 104.615
R1775 VTAIL.n392 VTAIL.n349 104.615
R1776 VTAIL.n399 VTAIL.n349 104.615
R1777 VTAIL.n400 VTAIL.n399 104.615
R1778 VTAIL.n400 VTAIL.n345 104.615
R1779 VTAIL.n408 VTAIL.n345 104.615
R1780 VTAIL.n409 VTAIL.n408 104.615
R1781 VTAIL.n410 VTAIL.n409 104.615
R1782 VTAIL.n410 VTAIL.n341 104.615
R1783 VTAIL.n417 VTAIL.n341 104.615
R1784 VTAIL.n418 VTAIL.n417 104.615
R1785 VTAIL.n418 VTAIL.n337 104.615
R1786 VTAIL.n425 VTAIL.n337 104.615
R1787 VTAIL.n426 VTAIL.n425 104.615
R1788 VTAIL.n426 VTAIL.n333 104.615
R1789 VTAIL.n433 VTAIL.n333 104.615
R1790 VTAIL.n434 VTAIL.n433 104.615
R1791 VTAIL.n38 VTAIL.n37 104.615
R1792 VTAIL.n38 VTAIL.n31 104.615
R1793 VTAIL.n45 VTAIL.n31 104.615
R1794 VTAIL.n46 VTAIL.n45 104.615
R1795 VTAIL.n46 VTAIL.n27 104.615
R1796 VTAIL.n53 VTAIL.n27 104.615
R1797 VTAIL.n54 VTAIL.n53 104.615
R1798 VTAIL.n54 VTAIL.n23 104.615
R1799 VTAIL.n61 VTAIL.n23 104.615
R1800 VTAIL.n62 VTAIL.n61 104.615
R1801 VTAIL.n62 VTAIL.n19 104.615
R1802 VTAIL.n69 VTAIL.n19 104.615
R1803 VTAIL.n70 VTAIL.n69 104.615
R1804 VTAIL.n70 VTAIL.n15 104.615
R1805 VTAIL.n78 VTAIL.n15 104.615
R1806 VTAIL.n79 VTAIL.n78 104.615
R1807 VTAIL.n80 VTAIL.n79 104.615
R1808 VTAIL.n80 VTAIL.n11 104.615
R1809 VTAIL.n87 VTAIL.n11 104.615
R1810 VTAIL.n88 VTAIL.n87 104.615
R1811 VTAIL.n88 VTAIL.n7 104.615
R1812 VTAIL.n95 VTAIL.n7 104.615
R1813 VTAIL.n96 VTAIL.n95 104.615
R1814 VTAIL.n96 VTAIL.n3 104.615
R1815 VTAIL.n103 VTAIL.n3 104.615
R1816 VTAIL.n104 VTAIL.n103 104.615
R1817 VTAIL.n324 VTAIL.n323 104.615
R1818 VTAIL.n323 VTAIL.n223 104.615
R1819 VTAIL.n316 VTAIL.n223 104.615
R1820 VTAIL.n316 VTAIL.n315 104.615
R1821 VTAIL.n315 VTAIL.n227 104.615
R1822 VTAIL.n308 VTAIL.n227 104.615
R1823 VTAIL.n308 VTAIL.n307 104.615
R1824 VTAIL.n307 VTAIL.n231 104.615
R1825 VTAIL.n236 VTAIL.n231 104.615
R1826 VTAIL.n300 VTAIL.n236 104.615
R1827 VTAIL.n300 VTAIL.n299 104.615
R1828 VTAIL.n299 VTAIL.n237 104.615
R1829 VTAIL.n292 VTAIL.n237 104.615
R1830 VTAIL.n292 VTAIL.n291 104.615
R1831 VTAIL.n291 VTAIL.n241 104.615
R1832 VTAIL.n284 VTAIL.n241 104.615
R1833 VTAIL.n284 VTAIL.n283 104.615
R1834 VTAIL.n283 VTAIL.n245 104.615
R1835 VTAIL.n276 VTAIL.n245 104.615
R1836 VTAIL.n276 VTAIL.n275 104.615
R1837 VTAIL.n275 VTAIL.n249 104.615
R1838 VTAIL.n268 VTAIL.n249 104.615
R1839 VTAIL.n268 VTAIL.n267 104.615
R1840 VTAIL.n267 VTAIL.n253 104.615
R1841 VTAIL.n260 VTAIL.n253 104.615
R1842 VTAIL.n260 VTAIL.n259 104.615
R1843 VTAIL.n214 VTAIL.n213 104.615
R1844 VTAIL.n213 VTAIL.n113 104.615
R1845 VTAIL.n206 VTAIL.n113 104.615
R1846 VTAIL.n206 VTAIL.n205 104.615
R1847 VTAIL.n205 VTAIL.n117 104.615
R1848 VTAIL.n198 VTAIL.n117 104.615
R1849 VTAIL.n198 VTAIL.n197 104.615
R1850 VTAIL.n197 VTAIL.n121 104.615
R1851 VTAIL.n126 VTAIL.n121 104.615
R1852 VTAIL.n190 VTAIL.n126 104.615
R1853 VTAIL.n190 VTAIL.n189 104.615
R1854 VTAIL.n189 VTAIL.n127 104.615
R1855 VTAIL.n182 VTAIL.n127 104.615
R1856 VTAIL.n182 VTAIL.n181 104.615
R1857 VTAIL.n181 VTAIL.n131 104.615
R1858 VTAIL.n174 VTAIL.n131 104.615
R1859 VTAIL.n174 VTAIL.n173 104.615
R1860 VTAIL.n173 VTAIL.n135 104.615
R1861 VTAIL.n166 VTAIL.n135 104.615
R1862 VTAIL.n166 VTAIL.n165 104.615
R1863 VTAIL.n165 VTAIL.n139 104.615
R1864 VTAIL.n158 VTAIL.n139 104.615
R1865 VTAIL.n158 VTAIL.n157 104.615
R1866 VTAIL.n157 VTAIL.n143 104.615
R1867 VTAIL.n150 VTAIL.n143 104.615
R1868 VTAIL.n150 VTAIL.n149 104.615
R1869 VTAIL.n367 VTAIL.t3 52.3082
R1870 VTAIL.n37 VTAIL.t0 52.3082
R1871 VTAIL.n259 VTAIL.t1 52.3082
R1872 VTAIL.n149 VTAIL.t2 52.3082
R1873 VTAIL.n219 VTAIL.n109 35.1945
R1874 VTAIL.n439 VTAIL.n438 32.5732
R1875 VTAIL.n109 VTAIL.n108 32.5732
R1876 VTAIL.n329 VTAIL.n328 32.5732
R1877 VTAIL.n219 VTAIL.n218 32.5732
R1878 VTAIL.n439 VTAIL.n329 32.2721
R1879 VTAIL.n366 VTAIL.n365 15.6677
R1880 VTAIL.n36 VTAIL.n35 15.6677
R1881 VTAIL.n258 VTAIL.n257 15.6677
R1882 VTAIL.n148 VTAIL.n147 15.6677
R1883 VTAIL.n411 VTAIL.n342 13.1884
R1884 VTAIL.n81 VTAIL.n12 13.1884
R1885 VTAIL.n234 VTAIL.n232 13.1884
R1886 VTAIL.n124 VTAIL.n122 13.1884
R1887 VTAIL.n369 VTAIL.n364 12.8005
R1888 VTAIL.n412 VTAIL.n344 12.8005
R1889 VTAIL.n416 VTAIL.n415 12.8005
R1890 VTAIL.n39 VTAIL.n34 12.8005
R1891 VTAIL.n82 VTAIL.n14 12.8005
R1892 VTAIL.n86 VTAIL.n85 12.8005
R1893 VTAIL.n306 VTAIL.n305 12.8005
R1894 VTAIL.n302 VTAIL.n301 12.8005
R1895 VTAIL.n261 VTAIL.n256 12.8005
R1896 VTAIL.n196 VTAIL.n195 12.8005
R1897 VTAIL.n192 VTAIL.n191 12.8005
R1898 VTAIL.n151 VTAIL.n146 12.8005
R1899 VTAIL.n370 VTAIL.n362 12.0247
R1900 VTAIL.n407 VTAIL.n406 12.0247
R1901 VTAIL.n419 VTAIL.n340 12.0247
R1902 VTAIL.n40 VTAIL.n32 12.0247
R1903 VTAIL.n77 VTAIL.n76 12.0247
R1904 VTAIL.n89 VTAIL.n10 12.0247
R1905 VTAIL.n309 VTAIL.n230 12.0247
R1906 VTAIL.n298 VTAIL.n235 12.0247
R1907 VTAIL.n262 VTAIL.n254 12.0247
R1908 VTAIL.n199 VTAIL.n120 12.0247
R1909 VTAIL.n188 VTAIL.n125 12.0247
R1910 VTAIL.n152 VTAIL.n144 12.0247
R1911 VTAIL.n374 VTAIL.n373 11.249
R1912 VTAIL.n405 VTAIL.n346 11.249
R1913 VTAIL.n420 VTAIL.n338 11.249
R1914 VTAIL.n44 VTAIL.n43 11.249
R1915 VTAIL.n75 VTAIL.n16 11.249
R1916 VTAIL.n90 VTAIL.n8 11.249
R1917 VTAIL.n310 VTAIL.n228 11.249
R1918 VTAIL.n297 VTAIL.n238 11.249
R1919 VTAIL.n266 VTAIL.n265 11.249
R1920 VTAIL.n200 VTAIL.n118 11.249
R1921 VTAIL.n187 VTAIL.n128 11.249
R1922 VTAIL.n156 VTAIL.n155 11.249
R1923 VTAIL.n377 VTAIL.n360 10.4732
R1924 VTAIL.n402 VTAIL.n401 10.4732
R1925 VTAIL.n424 VTAIL.n423 10.4732
R1926 VTAIL.n47 VTAIL.n30 10.4732
R1927 VTAIL.n72 VTAIL.n71 10.4732
R1928 VTAIL.n94 VTAIL.n93 10.4732
R1929 VTAIL.n314 VTAIL.n313 10.4732
R1930 VTAIL.n294 VTAIL.n293 10.4732
R1931 VTAIL.n269 VTAIL.n252 10.4732
R1932 VTAIL.n204 VTAIL.n203 10.4732
R1933 VTAIL.n184 VTAIL.n183 10.4732
R1934 VTAIL.n159 VTAIL.n142 10.4732
R1935 VTAIL.n378 VTAIL.n358 9.69747
R1936 VTAIL.n398 VTAIL.n348 9.69747
R1937 VTAIL.n427 VTAIL.n336 9.69747
R1938 VTAIL.n48 VTAIL.n28 9.69747
R1939 VTAIL.n68 VTAIL.n18 9.69747
R1940 VTAIL.n97 VTAIL.n6 9.69747
R1941 VTAIL.n317 VTAIL.n226 9.69747
R1942 VTAIL.n290 VTAIL.n240 9.69747
R1943 VTAIL.n270 VTAIL.n250 9.69747
R1944 VTAIL.n207 VTAIL.n116 9.69747
R1945 VTAIL.n180 VTAIL.n130 9.69747
R1946 VTAIL.n160 VTAIL.n140 9.69747
R1947 VTAIL.n438 VTAIL.n437 9.45567
R1948 VTAIL.n108 VTAIL.n107 9.45567
R1949 VTAIL.n328 VTAIL.n327 9.45567
R1950 VTAIL.n218 VTAIL.n217 9.45567
R1951 VTAIL.n437 VTAIL.n436 9.3005
R1952 VTAIL.n431 VTAIL.n430 9.3005
R1953 VTAIL.n429 VTAIL.n428 9.3005
R1954 VTAIL.n336 VTAIL.n335 9.3005
R1955 VTAIL.n423 VTAIL.n422 9.3005
R1956 VTAIL.n421 VTAIL.n420 9.3005
R1957 VTAIL.n340 VTAIL.n339 9.3005
R1958 VTAIL.n415 VTAIL.n414 9.3005
R1959 VTAIL.n387 VTAIL.n386 9.3005
R1960 VTAIL.n356 VTAIL.n355 9.3005
R1961 VTAIL.n381 VTAIL.n380 9.3005
R1962 VTAIL.n379 VTAIL.n378 9.3005
R1963 VTAIL.n360 VTAIL.n359 9.3005
R1964 VTAIL.n373 VTAIL.n372 9.3005
R1965 VTAIL.n371 VTAIL.n370 9.3005
R1966 VTAIL.n364 VTAIL.n363 9.3005
R1967 VTAIL.n389 VTAIL.n388 9.3005
R1968 VTAIL.n352 VTAIL.n351 9.3005
R1969 VTAIL.n395 VTAIL.n394 9.3005
R1970 VTAIL.n397 VTAIL.n396 9.3005
R1971 VTAIL.n348 VTAIL.n347 9.3005
R1972 VTAIL.n403 VTAIL.n402 9.3005
R1973 VTAIL.n405 VTAIL.n404 9.3005
R1974 VTAIL.n406 VTAIL.n343 9.3005
R1975 VTAIL.n413 VTAIL.n412 9.3005
R1976 VTAIL.n332 VTAIL.n331 9.3005
R1977 VTAIL.n107 VTAIL.n106 9.3005
R1978 VTAIL.n101 VTAIL.n100 9.3005
R1979 VTAIL.n99 VTAIL.n98 9.3005
R1980 VTAIL.n6 VTAIL.n5 9.3005
R1981 VTAIL.n93 VTAIL.n92 9.3005
R1982 VTAIL.n91 VTAIL.n90 9.3005
R1983 VTAIL.n10 VTAIL.n9 9.3005
R1984 VTAIL.n85 VTAIL.n84 9.3005
R1985 VTAIL.n57 VTAIL.n56 9.3005
R1986 VTAIL.n26 VTAIL.n25 9.3005
R1987 VTAIL.n51 VTAIL.n50 9.3005
R1988 VTAIL.n49 VTAIL.n48 9.3005
R1989 VTAIL.n30 VTAIL.n29 9.3005
R1990 VTAIL.n43 VTAIL.n42 9.3005
R1991 VTAIL.n41 VTAIL.n40 9.3005
R1992 VTAIL.n34 VTAIL.n33 9.3005
R1993 VTAIL.n59 VTAIL.n58 9.3005
R1994 VTAIL.n22 VTAIL.n21 9.3005
R1995 VTAIL.n65 VTAIL.n64 9.3005
R1996 VTAIL.n67 VTAIL.n66 9.3005
R1997 VTAIL.n18 VTAIL.n17 9.3005
R1998 VTAIL.n73 VTAIL.n72 9.3005
R1999 VTAIL.n75 VTAIL.n74 9.3005
R2000 VTAIL.n76 VTAIL.n13 9.3005
R2001 VTAIL.n83 VTAIL.n82 9.3005
R2002 VTAIL.n2 VTAIL.n1 9.3005
R2003 VTAIL.n244 VTAIL.n243 9.3005
R2004 VTAIL.n287 VTAIL.n286 9.3005
R2005 VTAIL.n289 VTAIL.n288 9.3005
R2006 VTAIL.n240 VTAIL.n239 9.3005
R2007 VTAIL.n295 VTAIL.n294 9.3005
R2008 VTAIL.n297 VTAIL.n296 9.3005
R2009 VTAIL.n235 VTAIL.n233 9.3005
R2010 VTAIL.n303 VTAIL.n302 9.3005
R2011 VTAIL.n327 VTAIL.n326 9.3005
R2012 VTAIL.n222 VTAIL.n221 9.3005
R2013 VTAIL.n321 VTAIL.n320 9.3005
R2014 VTAIL.n319 VTAIL.n318 9.3005
R2015 VTAIL.n226 VTAIL.n225 9.3005
R2016 VTAIL.n313 VTAIL.n312 9.3005
R2017 VTAIL.n311 VTAIL.n310 9.3005
R2018 VTAIL.n230 VTAIL.n229 9.3005
R2019 VTAIL.n305 VTAIL.n304 9.3005
R2020 VTAIL.n281 VTAIL.n280 9.3005
R2021 VTAIL.n279 VTAIL.n278 9.3005
R2022 VTAIL.n248 VTAIL.n247 9.3005
R2023 VTAIL.n273 VTAIL.n272 9.3005
R2024 VTAIL.n271 VTAIL.n270 9.3005
R2025 VTAIL.n252 VTAIL.n251 9.3005
R2026 VTAIL.n265 VTAIL.n264 9.3005
R2027 VTAIL.n263 VTAIL.n262 9.3005
R2028 VTAIL.n256 VTAIL.n255 9.3005
R2029 VTAIL.n134 VTAIL.n133 9.3005
R2030 VTAIL.n177 VTAIL.n176 9.3005
R2031 VTAIL.n179 VTAIL.n178 9.3005
R2032 VTAIL.n130 VTAIL.n129 9.3005
R2033 VTAIL.n185 VTAIL.n184 9.3005
R2034 VTAIL.n187 VTAIL.n186 9.3005
R2035 VTAIL.n125 VTAIL.n123 9.3005
R2036 VTAIL.n193 VTAIL.n192 9.3005
R2037 VTAIL.n217 VTAIL.n216 9.3005
R2038 VTAIL.n112 VTAIL.n111 9.3005
R2039 VTAIL.n211 VTAIL.n210 9.3005
R2040 VTAIL.n209 VTAIL.n208 9.3005
R2041 VTAIL.n116 VTAIL.n115 9.3005
R2042 VTAIL.n203 VTAIL.n202 9.3005
R2043 VTAIL.n201 VTAIL.n200 9.3005
R2044 VTAIL.n120 VTAIL.n119 9.3005
R2045 VTAIL.n195 VTAIL.n194 9.3005
R2046 VTAIL.n171 VTAIL.n170 9.3005
R2047 VTAIL.n169 VTAIL.n168 9.3005
R2048 VTAIL.n138 VTAIL.n137 9.3005
R2049 VTAIL.n163 VTAIL.n162 9.3005
R2050 VTAIL.n161 VTAIL.n160 9.3005
R2051 VTAIL.n142 VTAIL.n141 9.3005
R2052 VTAIL.n155 VTAIL.n154 9.3005
R2053 VTAIL.n153 VTAIL.n152 9.3005
R2054 VTAIL.n146 VTAIL.n145 9.3005
R2055 VTAIL.n382 VTAIL.n381 8.92171
R2056 VTAIL.n397 VTAIL.n350 8.92171
R2057 VTAIL.n428 VTAIL.n334 8.92171
R2058 VTAIL.n52 VTAIL.n51 8.92171
R2059 VTAIL.n67 VTAIL.n20 8.92171
R2060 VTAIL.n98 VTAIL.n4 8.92171
R2061 VTAIL.n318 VTAIL.n224 8.92171
R2062 VTAIL.n289 VTAIL.n242 8.92171
R2063 VTAIL.n274 VTAIL.n273 8.92171
R2064 VTAIL.n208 VTAIL.n114 8.92171
R2065 VTAIL.n179 VTAIL.n132 8.92171
R2066 VTAIL.n164 VTAIL.n163 8.92171
R2067 VTAIL.n385 VTAIL.n356 8.14595
R2068 VTAIL.n394 VTAIL.n393 8.14595
R2069 VTAIL.n432 VTAIL.n431 8.14595
R2070 VTAIL.n55 VTAIL.n26 8.14595
R2071 VTAIL.n64 VTAIL.n63 8.14595
R2072 VTAIL.n102 VTAIL.n101 8.14595
R2073 VTAIL.n322 VTAIL.n321 8.14595
R2074 VTAIL.n286 VTAIL.n285 8.14595
R2075 VTAIL.n277 VTAIL.n248 8.14595
R2076 VTAIL.n212 VTAIL.n211 8.14595
R2077 VTAIL.n176 VTAIL.n175 8.14595
R2078 VTAIL.n167 VTAIL.n138 8.14595
R2079 VTAIL.n386 VTAIL.n354 7.3702
R2080 VTAIL.n390 VTAIL.n352 7.3702
R2081 VTAIL.n435 VTAIL.n332 7.3702
R2082 VTAIL.n438 VTAIL.n330 7.3702
R2083 VTAIL.n56 VTAIL.n24 7.3702
R2084 VTAIL.n60 VTAIL.n22 7.3702
R2085 VTAIL.n105 VTAIL.n2 7.3702
R2086 VTAIL.n108 VTAIL.n0 7.3702
R2087 VTAIL.n328 VTAIL.n220 7.3702
R2088 VTAIL.n325 VTAIL.n222 7.3702
R2089 VTAIL.n282 VTAIL.n244 7.3702
R2090 VTAIL.n278 VTAIL.n246 7.3702
R2091 VTAIL.n218 VTAIL.n110 7.3702
R2092 VTAIL.n215 VTAIL.n112 7.3702
R2093 VTAIL.n172 VTAIL.n134 7.3702
R2094 VTAIL.n168 VTAIL.n136 7.3702
R2095 VTAIL.n389 VTAIL.n354 6.59444
R2096 VTAIL.n390 VTAIL.n389 6.59444
R2097 VTAIL.n436 VTAIL.n435 6.59444
R2098 VTAIL.n436 VTAIL.n330 6.59444
R2099 VTAIL.n59 VTAIL.n24 6.59444
R2100 VTAIL.n60 VTAIL.n59 6.59444
R2101 VTAIL.n106 VTAIL.n105 6.59444
R2102 VTAIL.n106 VTAIL.n0 6.59444
R2103 VTAIL.n326 VTAIL.n220 6.59444
R2104 VTAIL.n326 VTAIL.n325 6.59444
R2105 VTAIL.n282 VTAIL.n281 6.59444
R2106 VTAIL.n281 VTAIL.n246 6.59444
R2107 VTAIL.n216 VTAIL.n110 6.59444
R2108 VTAIL.n216 VTAIL.n215 6.59444
R2109 VTAIL.n172 VTAIL.n171 6.59444
R2110 VTAIL.n171 VTAIL.n136 6.59444
R2111 VTAIL.n386 VTAIL.n385 5.81868
R2112 VTAIL.n393 VTAIL.n352 5.81868
R2113 VTAIL.n432 VTAIL.n332 5.81868
R2114 VTAIL.n56 VTAIL.n55 5.81868
R2115 VTAIL.n63 VTAIL.n22 5.81868
R2116 VTAIL.n102 VTAIL.n2 5.81868
R2117 VTAIL.n322 VTAIL.n222 5.81868
R2118 VTAIL.n285 VTAIL.n244 5.81868
R2119 VTAIL.n278 VTAIL.n277 5.81868
R2120 VTAIL.n212 VTAIL.n112 5.81868
R2121 VTAIL.n175 VTAIL.n134 5.81868
R2122 VTAIL.n168 VTAIL.n167 5.81868
R2123 VTAIL.n382 VTAIL.n356 5.04292
R2124 VTAIL.n394 VTAIL.n350 5.04292
R2125 VTAIL.n431 VTAIL.n334 5.04292
R2126 VTAIL.n52 VTAIL.n26 5.04292
R2127 VTAIL.n64 VTAIL.n20 5.04292
R2128 VTAIL.n101 VTAIL.n4 5.04292
R2129 VTAIL.n321 VTAIL.n224 5.04292
R2130 VTAIL.n286 VTAIL.n242 5.04292
R2131 VTAIL.n274 VTAIL.n248 5.04292
R2132 VTAIL.n211 VTAIL.n114 5.04292
R2133 VTAIL.n176 VTAIL.n132 5.04292
R2134 VTAIL.n164 VTAIL.n138 5.04292
R2135 VTAIL.n365 VTAIL.n363 4.38563
R2136 VTAIL.n35 VTAIL.n33 4.38563
R2137 VTAIL.n257 VTAIL.n255 4.38563
R2138 VTAIL.n147 VTAIL.n145 4.38563
R2139 VTAIL.n381 VTAIL.n358 4.26717
R2140 VTAIL.n398 VTAIL.n397 4.26717
R2141 VTAIL.n428 VTAIL.n427 4.26717
R2142 VTAIL.n51 VTAIL.n28 4.26717
R2143 VTAIL.n68 VTAIL.n67 4.26717
R2144 VTAIL.n98 VTAIL.n97 4.26717
R2145 VTAIL.n318 VTAIL.n317 4.26717
R2146 VTAIL.n290 VTAIL.n289 4.26717
R2147 VTAIL.n273 VTAIL.n250 4.26717
R2148 VTAIL.n208 VTAIL.n207 4.26717
R2149 VTAIL.n180 VTAIL.n179 4.26717
R2150 VTAIL.n163 VTAIL.n140 4.26717
R2151 VTAIL.n378 VTAIL.n377 3.49141
R2152 VTAIL.n401 VTAIL.n348 3.49141
R2153 VTAIL.n424 VTAIL.n336 3.49141
R2154 VTAIL.n48 VTAIL.n47 3.49141
R2155 VTAIL.n71 VTAIL.n18 3.49141
R2156 VTAIL.n94 VTAIL.n6 3.49141
R2157 VTAIL.n314 VTAIL.n226 3.49141
R2158 VTAIL.n293 VTAIL.n240 3.49141
R2159 VTAIL.n270 VTAIL.n269 3.49141
R2160 VTAIL.n204 VTAIL.n116 3.49141
R2161 VTAIL.n183 VTAIL.n130 3.49141
R2162 VTAIL.n160 VTAIL.n159 3.49141
R2163 VTAIL.n374 VTAIL.n360 2.71565
R2164 VTAIL.n402 VTAIL.n346 2.71565
R2165 VTAIL.n423 VTAIL.n338 2.71565
R2166 VTAIL.n44 VTAIL.n30 2.71565
R2167 VTAIL.n72 VTAIL.n16 2.71565
R2168 VTAIL.n93 VTAIL.n8 2.71565
R2169 VTAIL.n313 VTAIL.n228 2.71565
R2170 VTAIL.n294 VTAIL.n238 2.71565
R2171 VTAIL.n266 VTAIL.n252 2.71565
R2172 VTAIL.n203 VTAIL.n118 2.71565
R2173 VTAIL.n184 VTAIL.n128 2.71565
R2174 VTAIL.n156 VTAIL.n142 2.71565
R2175 VTAIL.n373 VTAIL.n362 1.93989
R2176 VTAIL.n407 VTAIL.n405 1.93989
R2177 VTAIL.n420 VTAIL.n419 1.93989
R2178 VTAIL.n43 VTAIL.n32 1.93989
R2179 VTAIL.n77 VTAIL.n75 1.93989
R2180 VTAIL.n90 VTAIL.n89 1.93989
R2181 VTAIL.n310 VTAIL.n309 1.93989
R2182 VTAIL.n298 VTAIL.n297 1.93989
R2183 VTAIL.n265 VTAIL.n254 1.93989
R2184 VTAIL.n200 VTAIL.n199 1.93989
R2185 VTAIL.n188 VTAIL.n187 1.93989
R2186 VTAIL.n155 VTAIL.n144 1.93989
R2187 VTAIL.n329 VTAIL.n219 1.93153
R2188 VTAIL VTAIL.n109 1.25912
R2189 VTAIL.n370 VTAIL.n369 1.16414
R2190 VTAIL.n406 VTAIL.n344 1.16414
R2191 VTAIL.n416 VTAIL.n340 1.16414
R2192 VTAIL.n40 VTAIL.n39 1.16414
R2193 VTAIL.n76 VTAIL.n14 1.16414
R2194 VTAIL.n86 VTAIL.n10 1.16414
R2195 VTAIL.n306 VTAIL.n230 1.16414
R2196 VTAIL.n301 VTAIL.n235 1.16414
R2197 VTAIL.n262 VTAIL.n261 1.16414
R2198 VTAIL.n196 VTAIL.n120 1.16414
R2199 VTAIL.n191 VTAIL.n125 1.16414
R2200 VTAIL.n152 VTAIL.n151 1.16414
R2201 VTAIL VTAIL.n439 0.672914
R2202 VTAIL.n366 VTAIL.n364 0.388379
R2203 VTAIL.n412 VTAIL.n411 0.388379
R2204 VTAIL.n415 VTAIL.n342 0.388379
R2205 VTAIL.n36 VTAIL.n34 0.388379
R2206 VTAIL.n82 VTAIL.n81 0.388379
R2207 VTAIL.n85 VTAIL.n12 0.388379
R2208 VTAIL.n305 VTAIL.n232 0.388379
R2209 VTAIL.n302 VTAIL.n234 0.388379
R2210 VTAIL.n258 VTAIL.n256 0.388379
R2211 VTAIL.n195 VTAIL.n122 0.388379
R2212 VTAIL.n192 VTAIL.n124 0.388379
R2213 VTAIL.n148 VTAIL.n146 0.388379
R2214 VTAIL.n371 VTAIL.n363 0.155672
R2215 VTAIL.n372 VTAIL.n371 0.155672
R2216 VTAIL.n372 VTAIL.n359 0.155672
R2217 VTAIL.n379 VTAIL.n359 0.155672
R2218 VTAIL.n380 VTAIL.n379 0.155672
R2219 VTAIL.n380 VTAIL.n355 0.155672
R2220 VTAIL.n387 VTAIL.n355 0.155672
R2221 VTAIL.n388 VTAIL.n387 0.155672
R2222 VTAIL.n388 VTAIL.n351 0.155672
R2223 VTAIL.n395 VTAIL.n351 0.155672
R2224 VTAIL.n396 VTAIL.n395 0.155672
R2225 VTAIL.n396 VTAIL.n347 0.155672
R2226 VTAIL.n403 VTAIL.n347 0.155672
R2227 VTAIL.n404 VTAIL.n403 0.155672
R2228 VTAIL.n404 VTAIL.n343 0.155672
R2229 VTAIL.n413 VTAIL.n343 0.155672
R2230 VTAIL.n414 VTAIL.n413 0.155672
R2231 VTAIL.n414 VTAIL.n339 0.155672
R2232 VTAIL.n421 VTAIL.n339 0.155672
R2233 VTAIL.n422 VTAIL.n421 0.155672
R2234 VTAIL.n422 VTAIL.n335 0.155672
R2235 VTAIL.n429 VTAIL.n335 0.155672
R2236 VTAIL.n430 VTAIL.n429 0.155672
R2237 VTAIL.n430 VTAIL.n331 0.155672
R2238 VTAIL.n437 VTAIL.n331 0.155672
R2239 VTAIL.n41 VTAIL.n33 0.155672
R2240 VTAIL.n42 VTAIL.n41 0.155672
R2241 VTAIL.n42 VTAIL.n29 0.155672
R2242 VTAIL.n49 VTAIL.n29 0.155672
R2243 VTAIL.n50 VTAIL.n49 0.155672
R2244 VTAIL.n50 VTAIL.n25 0.155672
R2245 VTAIL.n57 VTAIL.n25 0.155672
R2246 VTAIL.n58 VTAIL.n57 0.155672
R2247 VTAIL.n58 VTAIL.n21 0.155672
R2248 VTAIL.n65 VTAIL.n21 0.155672
R2249 VTAIL.n66 VTAIL.n65 0.155672
R2250 VTAIL.n66 VTAIL.n17 0.155672
R2251 VTAIL.n73 VTAIL.n17 0.155672
R2252 VTAIL.n74 VTAIL.n73 0.155672
R2253 VTAIL.n74 VTAIL.n13 0.155672
R2254 VTAIL.n83 VTAIL.n13 0.155672
R2255 VTAIL.n84 VTAIL.n83 0.155672
R2256 VTAIL.n84 VTAIL.n9 0.155672
R2257 VTAIL.n91 VTAIL.n9 0.155672
R2258 VTAIL.n92 VTAIL.n91 0.155672
R2259 VTAIL.n92 VTAIL.n5 0.155672
R2260 VTAIL.n99 VTAIL.n5 0.155672
R2261 VTAIL.n100 VTAIL.n99 0.155672
R2262 VTAIL.n100 VTAIL.n1 0.155672
R2263 VTAIL.n107 VTAIL.n1 0.155672
R2264 VTAIL.n327 VTAIL.n221 0.155672
R2265 VTAIL.n320 VTAIL.n221 0.155672
R2266 VTAIL.n320 VTAIL.n319 0.155672
R2267 VTAIL.n319 VTAIL.n225 0.155672
R2268 VTAIL.n312 VTAIL.n225 0.155672
R2269 VTAIL.n312 VTAIL.n311 0.155672
R2270 VTAIL.n311 VTAIL.n229 0.155672
R2271 VTAIL.n304 VTAIL.n229 0.155672
R2272 VTAIL.n304 VTAIL.n303 0.155672
R2273 VTAIL.n303 VTAIL.n233 0.155672
R2274 VTAIL.n296 VTAIL.n233 0.155672
R2275 VTAIL.n296 VTAIL.n295 0.155672
R2276 VTAIL.n295 VTAIL.n239 0.155672
R2277 VTAIL.n288 VTAIL.n239 0.155672
R2278 VTAIL.n288 VTAIL.n287 0.155672
R2279 VTAIL.n287 VTAIL.n243 0.155672
R2280 VTAIL.n280 VTAIL.n243 0.155672
R2281 VTAIL.n280 VTAIL.n279 0.155672
R2282 VTAIL.n279 VTAIL.n247 0.155672
R2283 VTAIL.n272 VTAIL.n247 0.155672
R2284 VTAIL.n272 VTAIL.n271 0.155672
R2285 VTAIL.n271 VTAIL.n251 0.155672
R2286 VTAIL.n264 VTAIL.n251 0.155672
R2287 VTAIL.n264 VTAIL.n263 0.155672
R2288 VTAIL.n263 VTAIL.n255 0.155672
R2289 VTAIL.n217 VTAIL.n111 0.155672
R2290 VTAIL.n210 VTAIL.n111 0.155672
R2291 VTAIL.n210 VTAIL.n209 0.155672
R2292 VTAIL.n209 VTAIL.n115 0.155672
R2293 VTAIL.n202 VTAIL.n115 0.155672
R2294 VTAIL.n202 VTAIL.n201 0.155672
R2295 VTAIL.n201 VTAIL.n119 0.155672
R2296 VTAIL.n194 VTAIL.n119 0.155672
R2297 VTAIL.n194 VTAIL.n193 0.155672
R2298 VTAIL.n193 VTAIL.n123 0.155672
R2299 VTAIL.n186 VTAIL.n123 0.155672
R2300 VTAIL.n186 VTAIL.n185 0.155672
R2301 VTAIL.n185 VTAIL.n129 0.155672
R2302 VTAIL.n178 VTAIL.n129 0.155672
R2303 VTAIL.n178 VTAIL.n177 0.155672
R2304 VTAIL.n177 VTAIL.n133 0.155672
R2305 VTAIL.n170 VTAIL.n133 0.155672
R2306 VTAIL.n170 VTAIL.n169 0.155672
R2307 VTAIL.n169 VTAIL.n137 0.155672
R2308 VTAIL.n162 VTAIL.n137 0.155672
R2309 VTAIL.n162 VTAIL.n161 0.155672
R2310 VTAIL.n161 VTAIL.n141 0.155672
R2311 VTAIL.n154 VTAIL.n141 0.155672
R2312 VTAIL.n154 VTAIL.n153 0.155672
R2313 VTAIL.n153 VTAIL.n145 0.155672
R2314 VDD2.n213 VDD2.n109 289.615
R2315 VDD2.n104 VDD2.n0 289.615
R2316 VDD2.n214 VDD2.n213 185
R2317 VDD2.n212 VDD2.n211 185
R2318 VDD2.n113 VDD2.n112 185
R2319 VDD2.n206 VDD2.n205 185
R2320 VDD2.n204 VDD2.n203 185
R2321 VDD2.n117 VDD2.n116 185
R2322 VDD2.n198 VDD2.n197 185
R2323 VDD2.n196 VDD2.n195 185
R2324 VDD2.n121 VDD2.n120 185
R2325 VDD2.n125 VDD2.n123 185
R2326 VDD2.n190 VDD2.n189 185
R2327 VDD2.n188 VDD2.n187 185
R2328 VDD2.n127 VDD2.n126 185
R2329 VDD2.n182 VDD2.n181 185
R2330 VDD2.n180 VDD2.n179 185
R2331 VDD2.n131 VDD2.n130 185
R2332 VDD2.n174 VDD2.n173 185
R2333 VDD2.n172 VDD2.n171 185
R2334 VDD2.n135 VDD2.n134 185
R2335 VDD2.n166 VDD2.n165 185
R2336 VDD2.n164 VDD2.n163 185
R2337 VDD2.n139 VDD2.n138 185
R2338 VDD2.n158 VDD2.n157 185
R2339 VDD2.n156 VDD2.n155 185
R2340 VDD2.n143 VDD2.n142 185
R2341 VDD2.n150 VDD2.n149 185
R2342 VDD2.n148 VDD2.n147 185
R2343 VDD2.n37 VDD2.n36 185
R2344 VDD2.n39 VDD2.n38 185
R2345 VDD2.n32 VDD2.n31 185
R2346 VDD2.n45 VDD2.n44 185
R2347 VDD2.n47 VDD2.n46 185
R2348 VDD2.n28 VDD2.n27 185
R2349 VDD2.n53 VDD2.n52 185
R2350 VDD2.n55 VDD2.n54 185
R2351 VDD2.n24 VDD2.n23 185
R2352 VDD2.n61 VDD2.n60 185
R2353 VDD2.n63 VDD2.n62 185
R2354 VDD2.n20 VDD2.n19 185
R2355 VDD2.n69 VDD2.n68 185
R2356 VDD2.n71 VDD2.n70 185
R2357 VDD2.n16 VDD2.n15 185
R2358 VDD2.n78 VDD2.n77 185
R2359 VDD2.n79 VDD2.n14 185
R2360 VDD2.n81 VDD2.n80 185
R2361 VDD2.n12 VDD2.n11 185
R2362 VDD2.n87 VDD2.n86 185
R2363 VDD2.n89 VDD2.n88 185
R2364 VDD2.n8 VDD2.n7 185
R2365 VDD2.n95 VDD2.n94 185
R2366 VDD2.n97 VDD2.n96 185
R2367 VDD2.n4 VDD2.n3 185
R2368 VDD2.n103 VDD2.n102 185
R2369 VDD2.n105 VDD2.n104 185
R2370 VDD2.n146 VDD2.t1 147.659
R2371 VDD2.n35 VDD2.t0 147.659
R2372 VDD2.n213 VDD2.n212 104.615
R2373 VDD2.n212 VDD2.n112 104.615
R2374 VDD2.n205 VDD2.n112 104.615
R2375 VDD2.n205 VDD2.n204 104.615
R2376 VDD2.n204 VDD2.n116 104.615
R2377 VDD2.n197 VDD2.n116 104.615
R2378 VDD2.n197 VDD2.n196 104.615
R2379 VDD2.n196 VDD2.n120 104.615
R2380 VDD2.n125 VDD2.n120 104.615
R2381 VDD2.n189 VDD2.n125 104.615
R2382 VDD2.n189 VDD2.n188 104.615
R2383 VDD2.n188 VDD2.n126 104.615
R2384 VDD2.n181 VDD2.n126 104.615
R2385 VDD2.n181 VDD2.n180 104.615
R2386 VDD2.n180 VDD2.n130 104.615
R2387 VDD2.n173 VDD2.n130 104.615
R2388 VDD2.n173 VDD2.n172 104.615
R2389 VDD2.n172 VDD2.n134 104.615
R2390 VDD2.n165 VDD2.n134 104.615
R2391 VDD2.n165 VDD2.n164 104.615
R2392 VDD2.n164 VDD2.n138 104.615
R2393 VDD2.n157 VDD2.n138 104.615
R2394 VDD2.n157 VDD2.n156 104.615
R2395 VDD2.n156 VDD2.n142 104.615
R2396 VDD2.n149 VDD2.n142 104.615
R2397 VDD2.n149 VDD2.n148 104.615
R2398 VDD2.n38 VDD2.n37 104.615
R2399 VDD2.n38 VDD2.n31 104.615
R2400 VDD2.n45 VDD2.n31 104.615
R2401 VDD2.n46 VDD2.n45 104.615
R2402 VDD2.n46 VDD2.n27 104.615
R2403 VDD2.n53 VDD2.n27 104.615
R2404 VDD2.n54 VDD2.n53 104.615
R2405 VDD2.n54 VDD2.n23 104.615
R2406 VDD2.n61 VDD2.n23 104.615
R2407 VDD2.n62 VDD2.n61 104.615
R2408 VDD2.n62 VDD2.n19 104.615
R2409 VDD2.n69 VDD2.n19 104.615
R2410 VDD2.n70 VDD2.n69 104.615
R2411 VDD2.n70 VDD2.n15 104.615
R2412 VDD2.n78 VDD2.n15 104.615
R2413 VDD2.n79 VDD2.n78 104.615
R2414 VDD2.n80 VDD2.n79 104.615
R2415 VDD2.n80 VDD2.n11 104.615
R2416 VDD2.n87 VDD2.n11 104.615
R2417 VDD2.n88 VDD2.n87 104.615
R2418 VDD2.n88 VDD2.n7 104.615
R2419 VDD2.n95 VDD2.n7 104.615
R2420 VDD2.n96 VDD2.n95 104.615
R2421 VDD2.n96 VDD2.n3 104.615
R2422 VDD2.n103 VDD2.n3 104.615
R2423 VDD2.n104 VDD2.n103 104.615
R2424 VDD2.n218 VDD2.n108 95.739
R2425 VDD2.n148 VDD2.t1 52.3082
R2426 VDD2.n37 VDD2.t0 52.3082
R2427 VDD2.n218 VDD2.n217 49.252
R2428 VDD2.n147 VDD2.n146 15.6677
R2429 VDD2.n36 VDD2.n35 15.6677
R2430 VDD2.n123 VDD2.n121 13.1884
R2431 VDD2.n81 VDD2.n12 13.1884
R2432 VDD2.n195 VDD2.n194 12.8005
R2433 VDD2.n191 VDD2.n190 12.8005
R2434 VDD2.n150 VDD2.n145 12.8005
R2435 VDD2.n39 VDD2.n34 12.8005
R2436 VDD2.n82 VDD2.n14 12.8005
R2437 VDD2.n86 VDD2.n85 12.8005
R2438 VDD2.n198 VDD2.n119 12.0247
R2439 VDD2.n187 VDD2.n124 12.0247
R2440 VDD2.n151 VDD2.n143 12.0247
R2441 VDD2.n40 VDD2.n32 12.0247
R2442 VDD2.n77 VDD2.n76 12.0247
R2443 VDD2.n89 VDD2.n10 12.0247
R2444 VDD2.n199 VDD2.n117 11.249
R2445 VDD2.n186 VDD2.n127 11.249
R2446 VDD2.n155 VDD2.n154 11.249
R2447 VDD2.n44 VDD2.n43 11.249
R2448 VDD2.n75 VDD2.n16 11.249
R2449 VDD2.n90 VDD2.n8 11.249
R2450 VDD2.n203 VDD2.n202 10.4732
R2451 VDD2.n183 VDD2.n182 10.4732
R2452 VDD2.n158 VDD2.n141 10.4732
R2453 VDD2.n47 VDD2.n30 10.4732
R2454 VDD2.n72 VDD2.n71 10.4732
R2455 VDD2.n94 VDD2.n93 10.4732
R2456 VDD2.n206 VDD2.n115 9.69747
R2457 VDD2.n179 VDD2.n129 9.69747
R2458 VDD2.n159 VDD2.n139 9.69747
R2459 VDD2.n48 VDD2.n28 9.69747
R2460 VDD2.n68 VDD2.n18 9.69747
R2461 VDD2.n97 VDD2.n6 9.69747
R2462 VDD2.n217 VDD2.n216 9.45567
R2463 VDD2.n108 VDD2.n107 9.45567
R2464 VDD2.n133 VDD2.n132 9.3005
R2465 VDD2.n176 VDD2.n175 9.3005
R2466 VDD2.n178 VDD2.n177 9.3005
R2467 VDD2.n129 VDD2.n128 9.3005
R2468 VDD2.n184 VDD2.n183 9.3005
R2469 VDD2.n186 VDD2.n185 9.3005
R2470 VDD2.n124 VDD2.n122 9.3005
R2471 VDD2.n192 VDD2.n191 9.3005
R2472 VDD2.n216 VDD2.n215 9.3005
R2473 VDD2.n111 VDD2.n110 9.3005
R2474 VDD2.n210 VDD2.n209 9.3005
R2475 VDD2.n208 VDD2.n207 9.3005
R2476 VDD2.n115 VDD2.n114 9.3005
R2477 VDD2.n202 VDD2.n201 9.3005
R2478 VDD2.n200 VDD2.n199 9.3005
R2479 VDD2.n119 VDD2.n118 9.3005
R2480 VDD2.n194 VDD2.n193 9.3005
R2481 VDD2.n170 VDD2.n169 9.3005
R2482 VDD2.n168 VDD2.n167 9.3005
R2483 VDD2.n137 VDD2.n136 9.3005
R2484 VDD2.n162 VDD2.n161 9.3005
R2485 VDD2.n160 VDD2.n159 9.3005
R2486 VDD2.n141 VDD2.n140 9.3005
R2487 VDD2.n154 VDD2.n153 9.3005
R2488 VDD2.n152 VDD2.n151 9.3005
R2489 VDD2.n145 VDD2.n144 9.3005
R2490 VDD2.n107 VDD2.n106 9.3005
R2491 VDD2.n101 VDD2.n100 9.3005
R2492 VDD2.n99 VDD2.n98 9.3005
R2493 VDD2.n6 VDD2.n5 9.3005
R2494 VDD2.n93 VDD2.n92 9.3005
R2495 VDD2.n91 VDD2.n90 9.3005
R2496 VDD2.n10 VDD2.n9 9.3005
R2497 VDD2.n85 VDD2.n84 9.3005
R2498 VDD2.n57 VDD2.n56 9.3005
R2499 VDD2.n26 VDD2.n25 9.3005
R2500 VDD2.n51 VDD2.n50 9.3005
R2501 VDD2.n49 VDD2.n48 9.3005
R2502 VDD2.n30 VDD2.n29 9.3005
R2503 VDD2.n43 VDD2.n42 9.3005
R2504 VDD2.n41 VDD2.n40 9.3005
R2505 VDD2.n34 VDD2.n33 9.3005
R2506 VDD2.n59 VDD2.n58 9.3005
R2507 VDD2.n22 VDD2.n21 9.3005
R2508 VDD2.n65 VDD2.n64 9.3005
R2509 VDD2.n67 VDD2.n66 9.3005
R2510 VDD2.n18 VDD2.n17 9.3005
R2511 VDD2.n73 VDD2.n72 9.3005
R2512 VDD2.n75 VDD2.n74 9.3005
R2513 VDD2.n76 VDD2.n13 9.3005
R2514 VDD2.n83 VDD2.n82 9.3005
R2515 VDD2.n2 VDD2.n1 9.3005
R2516 VDD2.n207 VDD2.n113 8.92171
R2517 VDD2.n178 VDD2.n131 8.92171
R2518 VDD2.n163 VDD2.n162 8.92171
R2519 VDD2.n52 VDD2.n51 8.92171
R2520 VDD2.n67 VDD2.n20 8.92171
R2521 VDD2.n98 VDD2.n4 8.92171
R2522 VDD2.n211 VDD2.n210 8.14595
R2523 VDD2.n175 VDD2.n174 8.14595
R2524 VDD2.n166 VDD2.n137 8.14595
R2525 VDD2.n55 VDD2.n26 8.14595
R2526 VDD2.n64 VDD2.n63 8.14595
R2527 VDD2.n102 VDD2.n101 8.14595
R2528 VDD2.n217 VDD2.n109 7.3702
R2529 VDD2.n214 VDD2.n111 7.3702
R2530 VDD2.n171 VDD2.n133 7.3702
R2531 VDD2.n167 VDD2.n135 7.3702
R2532 VDD2.n56 VDD2.n24 7.3702
R2533 VDD2.n60 VDD2.n22 7.3702
R2534 VDD2.n105 VDD2.n2 7.3702
R2535 VDD2.n108 VDD2.n0 7.3702
R2536 VDD2.n215 VDD2.n109 6.59444
R2537 VDD2.n215 VDD2.n214 6.59444
R2538 VDD2.n171 VDD2.n170 6.59444
R2539 VDD2.n170 VDD2.n135 6.59444
R2540 VDD2.n59 VDD2.n24 6.59444
R2541 VDD2.n60 VDD2.n59 6.59444
R2542 VDD2.n106 VDD2.n105 6.59444
R2543 VDD2.n106 VDD2.n0 6.59444
R2544 VDD2.n211 VDD2.n111 5.81868
R2545 VDD2.n174 VDD2.n133 5.81868
R2546 VDD2.n167 VDD2.n166 5.81868
R2547 VDD2.n56 VDD2.n55 5.81868
R2548 VDD2.n63 VDD2.n22 5.81868
R2549 VDD2.n102 VDD2.n2 5.81868
R2550 VDD2.n210 VDD2.n113 5.04292
R2551 VDD2.n175 VDD2.n131 5.04292
R2552 VDD2.n163 VDD2.n137 5.04292
R2553 VDD2.n52 VDD2.n26 5.04292
R2554 VDD2.n64 VDD2.n20 5.04292
R2555 VDD2.n101 VDD2.n4 5.04292
R2556 VDD2.n146 VDD2.n144 4.38563
R2557 VDD2.n35 VDD2.n33 4.38563
R2558 VDD2.n207 VDD2.n206 4.26717
R2559 VDD2.n179 VDD2.n178 4.26717
R2560 VDD2.n162 VDD2.n139 4.26717
R2561 VDD2.n51 VDD2.n28 4.26717
R2562 VDD2.n68 VDD2.n67 4.26717
R2563 VDD2.n98 VDD2.n97 4.26717
R2564 VDD2.n203 VDD2.n115 3.49141
R2565 VDD2.n182 VDD2.n129 3.49141
R2566 VDD2.n159 VDD2.n158 3.49141
R2567 VDD2.n48 VDD2.n47 3.49141
R2568 VDD2.n71 VDD2.n18 3.49141
R2569 VDD2.n94 VDD2.n6 3.49141
R2570 VDD2.n202 VDD2.n117 2.71565
R2571 VDD2.n183 VDD2.n127 2.71565
R2572 VDD2.n155 VDD2.n141 2.71565
R2573 VDD2.n44 VDD2.n30 2.71565
R2574 VDD2.n72 VDD2.n16 2.71565
R2575 VDD2.n93 VDD2.n8 2.71565
R2576 VDD2.n199 VDD2.n198 1.93989
R2577 VDD2.n187 VDD2.n186 1.93989
R2578 VDD2.n154 VDD2.n143 1.93989
R2579 VDD2.n43 VDD2.n32 1.93989
R2580 VDD2.n77 VDD2.n75 1.93989
R2581 VDD2.n90 VDD2.n89 1.93989
R2582 VDD2.n195 VDD2.n119 1.16414
R2583 VDD2.n190 VDD2.n124 1.16414
R2584 VDD2.n151 VDD2.n150 1.16414
R2585 VDD2.n40 VDD2.n39 1.16414
R2586 VDD2.n76 VDD2.n14 1.16414
R2587 VDD2.n86 VDD2.n10 1.16414
R2588 VDD2 VDD2.n218 0.789293
R2589 VDD2.n194 VDD2.n121 0.388379
R2590 VDD2.n191 VDD2.n123 0.388379
R2591 VDD2.n147 VDD2.n145 0.388379
R2592 VDD2.n36 VDD2.n34 0.388379
R2593 VDD2.n82 VDD2.n81 0.388379
R2594 VDD2.n85 VDD2.n12 0.388379
R2595 VDD2.n216 VDD2.n110 0.155672
R2596 VDD2.n209 VDD2.n110 0.155672
R2597 VDD2.n209 VDD2.n208 0.155672
R2598 VDD2.n208 VDD2.n114 0.155672
R2599 VDD2.n201 VDD2.n114 0.155672
R2600 VDD2.n201 VDD2.n200 0.155672
R2601 VDD2.n200 VDD2.n118 0.155672
R2602 VDD2.n193 VDD2.n118 0.155672
R2603 VDD2.n193 VDD2.n192 0.155672
R2604 VDD2.n192 VDD2.n122 0.155672
R2605 VDD2.n185 VDD2.n122 0.155672
R2606 VDD2.n185 VDD2.n184 0.155672
R2607 VDD2.n184 VDD2.n128 0.155672
R2608 VDD2.n177 VDD2.n128 0.155672
R2609 VDD2.n177 VDD2.n176 0.155672
R2610 VDD2.n176 VDD2.n132 0.155672
R2611 VDD2.n169 VDD2.n132 0.155672
R2612 VDD2.n169 VDD2.n168 0.155672
R2613 VDD2.n168 VDD2.n136 0.155672
R2614 VDD2.n161 VDD2.n136 0.155672
R2615 VDD2.n161 VDD2.n160 0.155672
R2616 VDD2.n160 VDD2.n140 0.155672
R2617 VDD2.n153 VDD2.n140 0.155672
R2618 VDD2.n153 VDD2.n152 0.155672
R2619 VDD2.n152 VDD2.n144 0.155672
R2620 VDD2.n41 VDD2.n33 0.155672
R2621 VDD2.n42 VDD2.n41 0.155672
R2622 VDD2.n42 VDD2.n29 0.155672
R2623 VDD2.n49 VDD2.n29 0.155672
R2624 VDD2.n50 VDD2.n49 0.155672
R2625 VDD2.n50 VDD2.n25 0.155672
R2626 VDD2.n57 VDD2.n25 0.155672
R2627 VDD2.n58 VDD2.n57 0.155672
R2628 VDD2.n58 VDD2.n21 0.155672
R2629 VDD2.n65 VDD2.n21 0.155672
R2630 VDD2.n66 VDD2.n65 0.155672
R2631 VDD2.n66 VDD2.n17 0.155672
R2632 VDD2.n73 VDD2.n17 0.155672
R2633 VDD2.n74 VDD2.n73 0.155672
R2634 VDD2.n74 VDD2.n13 0.155672
R2635 VDD2.n83 VDD2.n13 0.155672
R2636 VDD2.n84 VDD2.n83 0.155672
R2637 VDD2.n84 VDD2.n9 0.155672
R2638 VDD2.n91 VDD2.n9 0.155672
R2639 VDD2.n92 VDD2.n91 0.155672
R2640 VDD2.n92 VDD2.n5 0.155672
R2641 VDD2.n99 VDD2.n5 0.155672
R2642 VDD2.n100 VDD2.n99 0.155672
R2643 VDD2.n100 VDD2.n1 0.155672
R2644 VDD2.n107 VDD2.n1 0.155672
R2645 VP.n0 VP.t0 248.001
R2646 VP.n0 VP.t1 196.292
R2647 VP VP.n0 0.431812
R2648 VDD1.n104 VDD1.n0 289.615
R2649 VDD1.n213 VDD1.n109 289.615
R2650 VDD1.n105 VDD1.n104 185
R2651 VDD1.n103 VDD1.n102 185
R2652 VDD1.n4 VDD1.n3 185
R2653 VDD1.n97 VDD1.n96 185
R2654 VDD1.n95 VDD1.n94 185
R2655 VDD1.n8 VDD1.n7 185
R2656 VDD1.n89 VDD1.n88 185
R2657 VDD1.n87 VDD1.n86 185
R2658 VDD1.n12 VDD1.n11 185
R2659 VDD1.n16 VDD1.n14 185
R2660 VDD1.n81 VDD1.n80 185
R2661 VDD1.n79 VDD1.n78 185
R2662 VDD1.n18 VDD1.n17 185
R2663 VDD1.n73 VDD1.n72 185
R2664 VDD1.n71 VDD1.n70 185
R2665 VDD1.n22 VDD1.n21 185
R2666 VDD1.n65 VDD1.n64 185
R2667 VDD1.n63 VDD1.n62 185
R2668 VDD1.n26 VDD1.n25 185
R2669 VDD1.n57 VDD1.n56 185
R2670 VDD1.n55 VDD1.n54 185
R2671 VDD1.n30 VDD1.n29 185
R2672 VDD1.n49 VDD1.n48 185
R2673 VDD1.n47 VDD1.n46 185
R2674 VDD1.n34 VDD1.n33 185
R2675 VDD1.n41 VDD1.n40 185
R2676 VDD1.n39 VDD1.n38 185
R2677 VDD1.n146 VDD1.n145 185
R2678 VDD1.n148 VDD1.n147 185
R2679 VDD1.n141 VDD1.n140 185
R2680 VDD1.n154 VDD1.n153 185
R2681 VDD1.n156 VDD1.n155 185
R2682 VDD1.n137 VDD1.n136 185
R2683 VDD1.n162 VDD1.n161 185
R2684 VDD1.n164 VDD1.n163 185
R2685 VDD1.n133 VDD1.n132 185
R2686 VDD1.n170 VDD1.n169 185
R2687 VDD1.n172 VDD1.n171 185
R2688 VDD1.n129 VDD1.n128 185
R2689 VDD1.n178 VDD1.n177 185
R2690 VDD1.n180 VDD1.n179 185
R2691 VDD1.n125 VDD1.n124 185
R2692 VDD1.n187 VDD1.n186 185
R2693 VDD1.n188 VDD1.n123 185
R2694 VDD1.n190 VDD1.n189 185
R2695 VDD1.n121 VDD1.n120 185
R2696 VDD1.n196 VDD1.n195 185
R2697 VDD1.n198 VDD1.n197 185
R2698 VDD1.n117 VDD1.n116 185
R2699 VDD1.n204 VDD1.n203 185
R2700 VDD1.n206 VDD1.n205 185
R2701 VDD1.n113 VDD1.n112 185
R2702 VDD1.n212 VDD1.n211 185
R2703 VDD1.n214 VDD1.n213 185
R2704 VDD1.n37 VDD1.t1 147.659
R2705 VDD1.n144 VDD1.t0 147.659
R2706 VDD1.n104 VDD1.n103 104.615
R2707 VDD1.n103 VDD1.n3 104.615
R2708 VDD1.n96 VDD1.n3 104.615
R2709 VDD1.n96 VDD1.n95 104.615
R2710 VDD1.n95 VDD1.n7 104.615
R2711 VDD1.n88 VDD1.n7 104.615
R2712 VDD1.n88 VDD1.n87 104.615
R2713 VDD1.n87 VDD1.n11 104.615
R2714 VDD1.n16 VDD1.n11 104.615
R2715 VDD1.n80 VDD1.n16 104.615
R2716 VDD1.n80 VDD1.n79 104.615
R2717 VDD1.n79 VDD1.n17 104.615
R2718 VDD1.n72 VDD1.n17 104.615
R2719 VDD1.n72 VDD1.n71 104.615
R2720 VDD1.n71 VDD1.n21 104.615
R2721 VDD1.n64 VDD1.n21 104.615
R2722 VDD1.n64 VDD1.n63 104.615
R2723 VDD1.n63 VDD1.n25 104.615
R2724 VDD1.n56 VDD1.n25 104.615
R2725 VDD1.n56 VDD1.n55 104.615
R2726 VDD1.n55 VDD1.n29 104.615
R2727 VDD1.n48 VDD1.n29 104.615
R2728 VDD1.n48 VDD1.n47 104.615
R2729 VDD1.n47 VDD1.n33 104.615
R2730 VDD1.n40 VDD1.n33 104.615
R2731 VDD1.n40 VDD1.n39 104.615
R2732 VDD1.n147 VDD1.n146 104.615
R2733 VDD1.n147 VDD1.n140 104.615
R2734 VDD1.n154 VDD1.n140 104.615
R2735 VDD1.n155 VDD1.n154 104.615
R2736 VDD1.n155 VDD1.n136 104.615
R2737 VDD1.n162 VDD1.n136 104.615
R2738 VDD1.n163 VDD1.n162 104.615
R2739 VDD1.n163 VDD1.n132 104.615
R2740 VDD1.n170 VDD1.n132 104.615
R2741 VDD1.n171 VDD1.n170 104.615
R2742 VDD1.n171 VDD1.n128 104.615
R2743 VDD1.n178 VDD1.n128 104.615
R2744 VDD1.n179 VDD1.n178 104.615
R2745 VDD1.n179 VDD1.n124 104.615
R2746 VDD1.n187 VDD1.n124 104.615
R2747 VDD1.n188 VDD1.n187 104.615
R2748 VDD1.n189 VDD1.n188 104.615
R2749 VDD1.n189 VDD1.n120 104.615
R2750 VDD1.n196 VDD1.n120 104.615
R2751 VDD1.n197 VDD1.n196 104.615
R2752 VDD1.n197 VDD1.n116 104.615
R2753 VDD1.n204 VDD1.n116 104.615
R2754 VDD1.n205 VDD1.n204 104.615
R2755 VDD1.n205 VDD1.n112 104.615
R2756 VDD1.n212 VDD1.n112 104.615
R2757 VDD1.n213 VDD1.n212 104.615
R2758 VDD1 VDD1.n217 96.9945
R2759 VDD1.n39 VDD1.t1 52.3082
R2760 VDD1.n146 VDD1.t0 52.3082
R2761 VDD1 VDD1.n108 50.0408
R2762 VDD1.n38 VDD1.n37 15.6677
R2763 VDD1.n145 VDD1.n144 15.6677
R2764 VDD1.n14 VDD1.n12 13.1884
R2765 VDD1.n190 VDD1.n121 13.1884
R2766 VDD1.n86 VDD1.n85 12.8005
R2767 VDD1.n82 VDD1.n81 12.8005
R2768 VDD1.n41 VDD1.n36 12.8005
R2769 VDD1.n148 VDD1.n143 12.8005
R2770 VDD1.n191 VDD1.n123 12.8005
R2771 VDD1.n195 VDD1.n194 12.8005
R2772 VDD1.n89 VDD1.n10 12.0247
R2773 VDD1.n78 VDD1.n15 12.0247
R2774 VDD1.n42 VDD1.n34 12.0247
R2775 VDD1.n149 VDD1.n141 12.0247
R2776 VDD1.n186 VDD1.n185 12.0247
R2777 VDD1.n198 VDD1.n119 12.0247
R2778 VDD1.n90 VDD1.n8 11.249
R2779 VDD1.n77 VDD1.n18 11.249
R2780 VDD1.n46 VDD1.n45 11.249
R2781 VDD1.n153 VDD1.n152 11.249
R2782 VDD1.n184 VDD1.n125 11.249
R2783 VDD1.n199 VDD1.n117 11.249
R2784 VDD1.n94 VDD1.n93 10.4732
R2785 VDD1.n74 VDD1.n73 10.4732
R2786 VDD1.n49 VDD1.n32 10.4732
R2787 VDD1.n156 VDD1.n139 10.4732
R2788 VDD1.n181 VDD1.n180 10.4732
R2789 VDD1.n203 VDD1.n202 10.4732
R2790 VDD1.n97 VDD1.n6 9.69747
R2791 VDD1.n70 VDD1.n20 9.69747
R2792 VDD1.n50 VDD1.n30 9.69747
R2793 VDD1.n157 VDD1.n137 9.69747
R2794 VDD1.n177 VDD1.n127 9.69747
R2795 VDD1.n206 VDD1.n115 9.69747
R2796 VDD1.n108 VDD1.n107 9.45567
R2797 VDD1.n217 VDD1.n216 9.45567
R2798 VDD1.n24 VDD1.n23 9.3005
R2799 VDD1.n67 VDD1.n66 9.3005
R2800 VDD1.n69 VDD1.n68 9.3005
R2801 VDD1.n20 VDD1.n19 9.3005
R2802 VDD1.n75 VDD1.n74 9.3005
R2803 VDD1.n77 VDD1.n76 9.3005
R2804 VDD1.n15 VDD1.n13 9.3005
R2805 VDD1.n83 VDD1.n82 9.3005
R2806 VDD1.n107 VDD1.n106 9.3005
R2807 VDD1.n2 VDD1.n1 9.3005
R2808 VDD1.n101 VDD1.n100 9.3005
R2809 VDD1.n99 VDD1.n98 9.3005
R2810 VDD1.n6 VDD1.n5 9.3005
R2811 VDD1.n93 VDD1.n92 9.3005
R2812 VDD1.n91 VDD1.n90 9.3005
R2813 VDD1.n10 VDD1.n9 9.3005
R2814 VDD1.n85 VDD1.n84 9.3005
R2815 VDD1.n61 VDD1.n60 9.3005
R2816 VDD1.n59 VDD1.n58 9.3005
R2817 VDD1.n28 VDD1.n27 9.3005
R2818 VDD1.n53 VDD1.n52 9.3005
R2819 VDD1.n51 VDD1.n50 9.3005
R2820 VDD1.n32 VDD1.n31 9.3005
R2821 VDD1.n45 VDD1.n44 9.3005
R2822 VDD1.n43 VDD1.n42 9.3005
R2823 VDD1.n36 VDD1.n35 9.3005
R2824 VDD1.n216 VDD1.n215 9.3005
R2825 VDD1.n210 VDD1.n209 9.3005
R2826 VDD1.n208 VDD1.n207 9.3005
R2827 VDD1.n115 VDD1.n114 9.3005
R2828 VDD1.n202 VDD1.n201 9.3005
R2829 VDD1.n200 VDD1.n199 9.3005
R2830 VDD1.n119 VDD1.n118 9.3005
R2831 VDD1.n194 VDD1.n193 9.3005
R2832 VDD1.n166 VDD1.n165 9.3005
R2833 VDD1.n135 VDD1.n134 9.3005
R2834 VDD1.n160 VDD1.n159 9.3005
R2835 VDD1.n158 VDD1.n157 9.3005
R2836 VDD1.n139 VDD1.n138 9.3005
R2837 VDD1.n152 VDD1.n151 9.3005
R2838 VDD1.n150 VDD1.n149 9.3005
R2839 VDD1.n143 VDD1.n142 9.3005
R2840 VDD1.n168 VDD1.n167 9.3005
R2841 VDD1.n131 VDD1.n130 9.3005
R2842 VDD1.n174 VDD1.n173 9.3005
R2843 VDD1.n176 VDD1.n175 9.3005
R2844 VDD1.n127 VDD1.n126 9.3005
R2845 VDD1.n182 VDD1.n181 9.3005
R2846 VDD1.n184 VDD1.n183 9.3005
R2847 VDD1.n185 VDD1.n122 9.3005
R2848 VDD1.n192 VDD1.n191 9.3005
R2849 VDD1.n111 VDD1.n110 9.3005
R2850 VDD1.n98 VDD1.n4 8.92171
R2851 VDD1.n69 VDD1.n22 8.92171
R2852 VDD1.n54 VDD1.n53 8.92171
R2853 VDD1.n161 VDD1.n160 8.92171
R2854 VDD1.n176 VDD1.n129 8.92171
R2855 VDD1.n207 VDD1.n113 8.92171
R2856 VDD1.n102 VDD1.n101 8.14595
R2857 VDD1.n66 VDD1.n65 8.14595
R2858 VDD1.n57 VDD1.n28 8.14595
R2859 VDD1.n164 VDD1.n135 8.14595
R2860 VDD1.n173 VDD1.n172 8.14595
R2861 VDD1.n211 VDD1.n210 8.14595
R2862 VDD1.n108 VDD1.n0 7.3702
R2863 VDD1.n105 VDD1.n2 7.3702
R2864 VDD1.n62 VDD1.n24 7.3702
R2865 VDD1.n58 VDD1.n26 7.3702
R2866 VDD1.n165 VDD1.n133 7.3702
R2867 VDD1.n169 VDD1.n131 7.3702
R2868 VDD1.n214 VDD1.n111 7.3702
R2869 VDD1.n217 VDD1.n109 7.3702
R2870 VDD1.n106 VDD1.n0 6.59444
R2871 VDD1.n106 VDD1.n105 6.59444
R2872 VDD1.n62 VDD1.n61 6.59444
R2873 VDD1.n61 VDD1.n26 6.59444
R2874 VDD1.n168 VDD1.n133 6.59444
R2875 VDD1.n169 VDD1.n168 6.59444
R2876 VDD1.n215 VDD1.n214 6.59444
R2877 VDD1.n215 VDD1.n109 6.59444
R2878 VDD1.n102 VDD1.n2 5.81868
R2879 VDD1.n65 VDD1.n24 5.81868
R2880 VDD1.n58 VDD1.n57 5.81868
R2881 VDD1.n165 VDD1.n164 5.81868
R2882 VDD1.n172 VDD1.n131 5.81868
R2883 VDD1.n211 VDD1.n111 5.81868
R2884 VDD1.n101 VDD1.n4 5.04292
R2885 VDD1.n66 VDD1.n22 5.04292
R2886 VDD1.n54 VDD1.n28 5.04292
R2887 VDD1.n161 VDD1.n135 5.04292
R2888 VDD1.n173 VDD1.n129 5.04292
R2889 VDD1.n210 VDD1.n113 5.04292
R2890 VDD1.n37 VDD1.n35 4.38563
R2891 VDD1.n144 VDD1.n142 4.38563
R2892 VDD1.n98 VDD1.n97 4.26717
R2893 VDD1.n70 VDD1.n69 4.26717
R2894 VDD1.n53 VDD1.n30 4.26717
R2895 VDD1.n160 VDD1.n137 4.26717
R2896 VDD1.n177 VDD1.n176 4.26717
R2897 VDD1.n207 VDD1.n206 4.26717
R2898 VDD1.n94 VDD1.n6 3.49141
R2899 VDD1.n73 VDD1.n20 3.49141
R2900 VDD1.n50 VDD1.n49 3.49141
R2901 VDD1.n157 VDD1.n156 3.49141
R2902 VDD1.n180 VDD1.n127 3.49141
R2903 VDD1.n203 VDD1.n115 3.49141
R2904 VDD1.n93 VDD1.n8 2.71565
R2905 VDD1.n74 VDD1.n18 2.71565
R2906 VDD1.n46 VDD1.n32 2.71565
R2907 VDD1.n153 VDD1.n139 2.71565
R2908 VDD1.n181 VDD1.n125 2.71565
R2909 VDD1.n202 VDD1.n117 2.71565
R2910 VDD1.n90 VDD1.n89 1.93989
R2911 VDD1.n78 VDD1.n77 1.93989
R2912 VDD1.n45 VDD1.n34 1.93989
R2913 VDD1.n152 VDD1.n141 1.93989
R2914 VDD1.n186 VDD1.n184 1.93989
R2915 VDD1.n199 VDD1.n198 1.93989
R2916 VDD1.n86 VDD1.n10 1.16414
R2917 VDD1.n81 VDD1.n15 1.16414
R2918 VDD1.n42 VDD1.n41 1.16414
R2919 VDD1.n149 VDD1.n148 1.16414
R2920 VDD1.n185 VDD1.n123 1.16414
R2921 VDD1.n195 VDD1.n119 1.16414
R2922 VDD1.n85 VDD1.n12 0.388379
R2923 VDD1.n82 VDD1.n14 0.388379
R2924 VDD1.n38 VDD1.n36 0.388379
R2925 VDD1.n145 VDD1.n143 0.388379
R2926 VDD1.n191 VDD1.n190 0.388379
R2927 VDD1.n194 VDD1.n121 0.388379
R2928 VDD1.n107 VDD1.n1 0.155672
R2929 VDD1.n100 VDD1.n1 0.155672
R2930 VDD1.n100 VDD1.n99 0.155672
R2931 VDD1.n99 VDD1.n5 0.155672
R2932 VDD1.n92 VDD1.n5 0.155672
R2933 VDD1.n92 VDD1.n91 0.155672
R2934 VDD1.n91 VDD1.n9 0.155672
R2935 VDD1.n84 VDD1.n9 0.155672
R2936 VDD1.n84 VDD1.n83 0.155672
R2937 VDD1.n83 VDD1.n13 0.155672
R2938 VDD1.n76 VDD1.n13 0.155672
R2939 VDD1.n76 VDD1.n75 0.155672
R2940 VDD1.n75 VDD1.n19 0.155672
R2941 VDD1.n68 VDD1.n19 0.155672
R2942 VDD1.n68 VDD1.n67 0.155672
R2943 VDD1.n67 VDD1.n23 0.155672
R2944 VDD1.n60 VDD1.n23 0.155672
R2945 VDD1.n60 VDD1.n59 0.155672
R2946 VDD1.n59 VDD1.n27 0.155672
R2947 VDD1.n52 VDD1.n27 0.155672
R2948 VDD1.n52 VDD1.n51 0.155672
R2949 VDD1.n51 VDD1.n31 0.155672
R2950 VDD1.n44 VDD1.n31 0.155672
R2951 VDD1.n44 VDD1.n43 0.155672
R2952 VDD1.n43 VDD1.n35 0.155672
R2953 VDD1.n150 VDD1.n142 0.155672
R2954 VDD1.n151 VDD1.n150 0.155672
R2955 VDD1.n151 VDD1.n138 0.155672
R2956 VDD1.n158 VDD1.n138 0.155672
R2957 VDD1.n159 VDD1.n158 0.155672
R2958 VDD1.n159 VDD1.n134 0.155672
R2959 VDD1.n166 VDD1.n134 0.155672
R2960 VDD1.n167 VDD1.n166 0.155672
R2961 VDD1.n167 VDD1.n130 0.155672
R2962 VDD1.n174 VDD1.n130 0.155672
R2963 VDD1.n175 VDD1.n174 0.155672
R2964 VDD1.n175 VDD1.n126 0.155672
R2965 VDD1.n182 VDD1.n126 0.155672
R2966 VDD1.n183 VDD1.n182 0.155672
R2967 VDD1.n183 VDD1.n122 0.155672
R2968 VDD1.n192 VDD1.n122 0.155672
R2969 VDD1.n193 VDD1.n192 0.155672
R2970 VDD1.n193 VDD1.n118 0.155672
R2971 VDD1.n200 VDD1.n118 0.155672
R2972 VDD1.n201 VDD1.n200 0.155672
R2973 VDD1.n201 VDD1.n114 0.155672
R2974 VDD1.n208 VDD1.n114 0.155672
R2975 VDD1.n209 VDD1.n208 0.155672
R2976 VDD1.n209 VDD1.n110 0.155672
R2977 VDD1.n216 VDD1.n110 0.155672
C0 VDD1 VDD2 0.731235f
C1 VDD1 VN 0.148667f
C2 VDD2 VN 4.51002f
C3 VP VDD1 4.71111f
C4 VP VDD2 0.353259f
C5 VDD1 VTAIL 7.12336f
C6 VDD2 VTAIL 7.17598f
C7 VP VN 7.09169f
C8 VN VTAIL 3.85841f
C9 VP VTAIL 3.87276f
C10 VDD2 B 5.970544f
C11 VDD1 B 9.343901f
C12 VTAIL B 10.730593f
C13 VN B 12.95328f
C14 VP B 7.478579f
C15 VDD1.n0 B 0.029409f
C16 VDD1.n1 B 0.019965f
C17 VDD1.n2 B 0.010728f
C18 VDD1.n3 B 0.025358f
C19 VDD1.n4 B 0.011359f
C20 VDD1.n5 B 0.019965f
C21 VDD1.n6 B 0.010728f
C22 VDD1.n7 B 0.025358f
C23 VDD1.n8 B 0.011359f
C24 VDD1.n9 B 0.019965f
C25 VDD1.n10 B 0.010728f
C26 VDD1.n11 B 0.025358f
C27 VDD1.n12 B 0.011044f
C28 VDD1.n13 B 0.019965f
C29 VDD1.n14 B 0.011044f
C30 VDD1.n15 B 0.010728f
C31 VDD1.n16 B 0.025358f
C32 VDD1.n17 B 0.025358f
C33 VDD1.n18 B 0.011359f
C34 VDD1.n19 B 0.019965f
C35 VDD1.n20 B 0.010728f
C36 VDD1.n21 B 0.025358f
C37 VDD1.n22 B 0.011359f
C38 VDD1.n23 B 0.019965f
C39 VDD1.n24 B 0.010728f
C40 VDD1.n25 B 0.025358f
C41 VDD1.n26 B 0.011359f
C42 VDD1.n27 B 0.019965f
C43 VDD1.n28 B 0.010728f
C44 VDD1.n29 B 0.025358f
C45 VDD1.n30 B 0.011359f
C46 VDD1.n31 B 0.019965f
C47 VDD1.n32 B 0.010728f
C48 VDD1.n33 B 0.025358f
C49 VDD1.n34 B 0.011359f
C50 VDD1.n35 B 1.72899f
C51 VDD1.n36 B 0.010728f
C52 VDD1.t1 B 0.042134f
C53 VDD1.n37 B 0.153742f
C54 VDD1.n38 B 0.014979f
C55 VDD1.n39 B 0.019018f
C56 VDD1.n40 B 0.025358f
C57 VDD1.n41 B 0.011359f
C58 VDD1.n42 B 0.010728f
C59 VDD1.n43 B 0.019965f
C60 VDD1.n44 B 0.019965f
C61 VDD1.n45 B 0.010728f
C62 VDD1.n46 B 0.011359f
C63 VDD1.n47 B 0.025358f
C64 VDD1.n48 B 0.025358f
C65 VDD1.n49 B 0.011359f
C66 VDD1.n50 B 0.010728f
C67 VDD1.n51 B 0.019965f
C68 VDD1.n52 B 0.019965f
C69 VDD1.n53 B 0.010728f
C70 VDD1.n54 B 0.011359f
C71 VDD1.n55 B 0.025358f
C72 VDD1.n56 B 0.025358f
C73 VDD1.n57 B 0.011359f
C74 VDD1.n58 B 0.010728f
C75 VDD1.n59 B 0.019965f
C76 VDD1.n60 B 0.019965f
C77 VDD1.n61 B 0.010728f
C78 VDD1.n62 B 0.011359f
C79 VDD1.n63 B 0.025358f
C80 VDD1.n64 B 0.025358f
C81 VDD1.n65 B 0.011359f
C82 VDD1.n66 B 0.010728f
C83 VDD1.n67 B 0.019965f
C84 VDD1.n68 B 0.019965f
C85 VDD1.n69 B 0.010728f
C86 VDD1.n70 B 0.011359f
C87 VDD1.n71 B 0.025358f
C88 VDD1.n72 B 0.025358f
C89 VDD1.n73 B 0.011359f
C90 VDD1.n74 B 0.010728f
C91 VDD1.n75 B 0.019965f
C92 VDD1.n76 B 0.019965f
C93 VDD1.n77 B 0.010728f
C94 VDD1.n78 B 0.011359f
C95 VDD1.n79 B 0.025358f
C96 VDD1.n80 B 0.025358f
C97 VDD1.n81 B 0.011359f
C98 VDD1.n82 B 0.010728f
C99 VDD1.n83 B 0.019965f
C100 VDD1.n84 B 0.019965f
C101 VDD1.n85 B 0.010728f
C102 VDD1.n86 B 0.011359f
C103 VDD1.n87 B 0.025358f
C104 VDD1.n88 B 0.025358f
C105 VDD1.n89 B 0.011359f
C106 VDD1.n90 B 0.010728f
C107 VDD1.n91 B 0.019965f
C108 VDD1.n92 B 0.019965f
C109 VDD1.n93 B 0.010728f
C110 VDD1.n94 B 0.011359f
C111 VDD1.n95 B 0.025358f
C112 VDD1.n96 B 0.025358f
C113 VDD1.n97 B 0.011359f
C114 VDD1.n98 B 0.010728f
C115 VDD1.n99 B 0.019965f
C116 VDD1.n100 B 0.019965f
C117 VDD1.n101 B 0.010728f
C118 VDD1.n102 B 0.011359f
C119 VDD1.n103 B 0.025358f
C120 VDD1.n104 B 0.057277f
C121 VDD1.n105 B 0.011359f
C122 VDD1.n106 B 0.010728f
C123 VDD1.n107 B 0.046693f
C124 VDD1.n108 B 0.047502f
C125 VDD1.n109 B 0.029409f
C126 VDD1.n110 B 0.019965f
C127 VDD1.n111 B 0.010728f
C128 VDD1.n112 B 0.025358f
C129 VDD1.n113 B 0.011359f
C130 VDD1.n114 B 0.019965f
C131 VDD1.n115 B 0.010728f
C132 VDD1.n116 B 0.025358f
C133 VDD1.n117 B 0.011359f
C134 VDD1.n118 B 0.019965f
C135 VDD1.n119 B 0.010728f
C136 VDD1.n120 B 0.025358f
C137 VDD1.n121 B 0.011044f
C138 VDD1.n122 B 0.019965f
C139 VDD1.n123 B 0.011359f
C140 VDD1.n124 B 0.025358f
C141 VDD1.n125 B 0.011359f
C142 VDD1.n126 B 0.019965f
C143 VDD1.n127 B 0.010728f
C144 VDD1.n128 B 0.025358f
C145 VDD1.n129 B 0.011359f
C146 VDD1.n130 B 0.019965f
C147 VDD1.n131 B 0.010728f
C148 VDD1.n132 B 0.025358f
C149 VDD1.n133 B 0.011359f
C150 VDD1.n134 B 0.019965f
C151 VDD1.n135 B 0.010728f
C152 VDD1.n136 B 0.025358f
C153 VDD1.n137 B 0.011359f
C154 VDD1.n138 B 0.019965f
C155 VDD1.n139 B 0.010728f
C156 VDD1.n140 B 0.025358f
C157 VDD1.n141 B 0.011359f
C158 VDD1.n142 B 1.72899f
C159 VDD1.n143 B 0.010728f
C160 VDD1.t0 B 0.042134f
C161 VDD1.n144 B 0.153742f
C162 VDD1.n145 B 0.014979f
C163 VDD1.n146 B 0.019018f
C164 VDD1.n147 B 0.025358f
C165 VDD1.n148 B 0.011359f
C166 VDD1.n149 B 0.010728f
C167 VDD1.n150 B 0.019965f
C168 VDD1.n151 B 0.019965f
C169 VDD1.n152 B 0.010728f
C170 VDD1.n153 B 0.011359f
C171 VDD1.n154 B 0.025358f
C172 VDD1.n155 B 0.025358f
C173 VDD1.n156 B 0.011359f
C174 VDD1.n157 B 0.010728f
C175 VDD1.n158 B 0.019965f
C176 VDD1.n159 B 0.019965f
C177 VDD1.n160 B 0.010728f
C178 VDD1.n161 B 0.011359f
C179 VDD1.n162 B 0.025358f
C180 VDD1.n163 B 0.025358f
C181 VDD1.n164 B 0.011359f
C182 VDD1.n165 B 0.010728f
C183 VDD1.n166 B 0.019965f
C184 VDD1.n167 B 0.019965f
C185 VDD1.n168 B 0.010728f
C186 VDD1.n169 B 0.011359f
C187 VDD1.n170 B 0.025358f
C188 VDD1.n171 B 0.025358f
C189 VDD1.n172 B 0.011359f
C190 VDD1.n173 B 0.010728f
C191 VDD1.n174 B 0.019965f
C192 VDD1.n175 B 0.019965f
C193 VDD1.n176 B 0.010728f
C194 VDD1.n177 B 0.011359f
C195 VDD1.n178 B 0.025358f
C196 VDD1.n179 B 0.025358f
C197 VDD1.n180 B 0.011359f
C198 VDD1.n181 B 0.010728f
C199 VDD1.n182 B 0.019965f
C200 VDD1.n183 B 0.019965f
C201 VDD1.n184 B 0.010728f
C202 VDD1.n185 B 0.010728f
C203 VDD1.n186 B 0.011359f
C204 VDD1.n187 B 0.025358f
C205 VDD1.n188 B 0.025358f
C206 VDD1.n189 B 0.025358f
C207 VDD1.n190 B 0.011044f
C208 VDD1.n191 B 0.010728f
C209 VDD1.n192 B 0.019965f
C210 VDD1.n193 B 0.019965f
C211 VDD1.n194 B 0.010728f
C212 VDD1.n195 B 0.011359f
C213 VDD1.n196 B 0.025358f
C214 VDD1.n197 B 0.025358f
C215 VDD1.n198 B 0.011359f
C216 VDD1.n199 B 0.010728f
C217 VDD1.n200 B 0.019965f
C218 VDD1.n201 B 0.019965f
C219 VDD1.n202 B 0.010728f
C220 VDD1.n203 B 0.011359f
C221 VDD1.n204 B 0.025358f
C222 VDD1.n205 B 0.025358f
C223 VDD1.n206 B 0.011359f
C224 VDD1.n207 B 0.010728f
C225 VDD1.n208 B 0.019965f
C226 VDD1.n209 B 0.019965f
C227 VDD1.n210 B 0.010728f
C228 VDD1.n211 B 0.011359f
C229 VDD1.n212 B 0.025358f
C230 VDD1.n213 B 0.057277f
C231 VDD1.n214 B 0.011359f
C232 VDD1.n215 B 0.010728f
C233 VDD1.n216 B 0.046693f
C234 VDD1.n217 B 0.892347f
C235 VP.t1 B 4.79239f
C236 VP.t0 B 5.42799f
C237 VP.n0 B 5.39844f
C238 VDD2.n0 B 0.029344f
C239 VDD2.n1 B 0.01992f
C240 VDD2.n2 B 0.010704f
C241 VDD2.n3 B 0.025301f
C242 VDD2.n4 B 0.011334f
C243 VDD2.n5 B 0.01992f
C244 VDD2.n6 B 0.010704f
C245 VDD2.n7 B 0.025301f
C246 VDD2.n8 B 0.011334f
C247 VDD2.n9 B 0.01992f
C248 VDD2.n10 B 0.010704f
C249 VDD2.n11 B 0.025301f
C250 VDD2.n12 B 0.011019f
C251 VDD2.n13 B 0.01992f
C252 VDD2.n14 B 0.011334f
C253 VDD2.n15 B 0.025301f
C254 VDD2.n16 B 0.011334f
C255 VDD2.n17 B 0.01992f
C256 VDD2.n18 B 0.010704f
C257 VDD2.n19 B 0.025301f
C258 VDD2.n20 B 0.011334f
C259 VDD2.n21 B 0.01992f
C260 VDD2.n22 B 0.010704f
C261 VDD2.n23 B 0.025301f
C262 VDD2.n24 B 0.011334f
C263 VDD2.n25 B 0.01992f
C264 VDD2.n26 B 0.010704f
C265 VDD2.n27 B 0.025301f
C266 VDD2.n28 B 0.011334f
C267 VDD2.n29 B 0.01992f
C268 VDD2.n30 B 0.010704f
C269 VDD2.n31 B 0.025301f
C270 VDD2.n32 B 0.011334f
C271 VDD2.n33 B 1.72511f
C272 VDD2.n34 B 0.010704f
C273 VDD2.t0 B 0.042039f
C274 VDD2.n35 B 0.153397f
C275 VDD2.n36 B 0.014946f
C276 VDD2.n37 B 0.018976f
C277 VDD2.n38 B 0.025301f
C278 VDD2.n39 B 0.011334f
C279 VDD2.n40 B 0.010704f
C280 VDD2.n41 B 0.01992f
C281 VDD2.n42 B 0.01992f
C282 VDD2.n43 B 0.010704f
C283 VDD2.n44 B 0.011334f
C284 VDD2.n45 B 0.025301f
C285 VDD2.n46 B 0.025301f
C286 VDD2.n47 B 0.011334f
C287 VDD2.n48 B 0.010704f
C288 VDD2.n49 B 0.01992f
C289 VDD2.n50 B 0.01992f
C290 VDD2.n51 B 0.010704f
C291 VDD2.n52 B 0.011334f
C292 VDD2.n53 B 0.025301f
C293 VDD2.n54 B 0.025301f
C294 VDD2.n55 B 0.011334f
C295 VDD2.n56 B 0.010704f
C296 VDD2.n57 B 0.01992f
C297 VDD2.n58 B 0.01992f
C298 VDD2.n59 B 0.010704f
C299 VDD2.n60 B 0.011334f
C300 VDD2.n61 B 0.025301f
C301 VDD2.n62 B 0.025301f
C302 VDD2.n63 B 0.011334f
C303 VDD2.n64 B 0.010704f
C304 VDD2.n65 B 0.01992f
C305 VDD2.n66 B 0.01992f
C306 VDD2.n67 B 0.010704f
C307 VDD2.n68 B 0.011334f
C308 VDD2.n69 B 0.025301f
C309 VDD2.n70 B 0.025301f
C310 VDD2.n71 B 0.011334f
C311 VDD2.n72 B 0.010704f
C312 VDD2.n73 B 0.01992f
C313 VDD2.n74 B 0.01992f
C314 VDD2.n75 B 0.010704f
C315 VDD2.n76 B 0.010704f
C316 VDD2.n77 B 0.011334f
C317 VDD2.n78 B 0.025301f
C318 VDD2.n79 B 0.025301f
C319 VDD2.n80 B 0.025301f
C320 VDD2.n81 B 0.011019f
C321 VDD2.n82 B 0.010704f
C322 VDD2.n83 B 0.01992f
C323 VDD2.n84 B 0.01992f
C324 VDD2.n85 B 0.010704f
C325 VDD2.n86 B 0.011334f
C326 VDD2.n87 B 0.025301f
C327 VDD2.n88 B 0.025301f
C328 VDD2.n89 B 0.011334f
C329 VDD2.n90 B 0.010704f
C330 VDD2.n91 B 0.01992f
C331 VDD2.n92 B 0.01992f
C332 VDD2.n93 B 0.010704f
C333 VDD2.n94 B 0.011334f
C334 VDD2.n95 B 0.025301f
C335 VDD2.n96 B 0.025301f
C336 VDD2.n97 B 0.011334f
C337 VDD2.n98 B 0.010704f
C338 VDD2.n99 B 0.01992f
C339 VDD2.n100 B 0.01992f
C340 VDD2.n101 B 0.010704f
C341 VDD2.n102 B 0.011334f
C342 VDD2.n103 B 0.025301f
C343 VDD2.n104 B 0.057149f
C344 VDD2.n105 B 0.011334f
C345 VDD2.n106 B 0.010704f
C346 VDD2.n107 B 0.046589f
C347 VDD2.n108 B 0.843102f
C348 VDD2.n109 B 0.029344f
C349 VDD2.n110 B 0.01992f
C350 VDD2.n111 B 0.010704f
C351 VDD2.n112 B 0.025301f
C352 VDD2.n113 B 0.011334f
C353 VDD2.n114 B 0.01992f
C354 VDD2.n115 B 0.010704f
C355 VDD2.n116 B 0.025301f
C356 VDD2.n117 B 0.011334f
C357 VDD2.n118 B 0.01992f
C358 VDD2.n119 B 0.010704f
C359 VDD2.n120 B 0.025301f
C360 VDD2.n121 B 0.011019f
C361 VDD2.n122 B 0.01992f
C362 VDD2.n123 B 0.011019f
C363 VDD2.n124 B 0.010704f
C364 VDD2.n125 B 0.025301f
C365 VDD2.n126 B 0.025301f
C366 VDD2.n127 B 0.011334f
C367 VDD2.n128 B 0.01992f
C368 VDD2.n129 B 0.010704f
C369 VDD2.n130 B 0.025301f
C370 VDD2.n131 B 0.011334f
C371 VDD2.n132 B 0.01992f
C372 VDD2.n133 B 0.010704f
C373 VDD2.n134 B 0.025301f
C374 VDD2.n135 B 0.011334f
C375 VDD2.n136 B 0.01992f
C376 VDD2.n137 B 0.010704f
C377 VDD2.n138 B 0.025301f
C378 VDD2.n139 B 0.011334f
C379 VDD2.n140 B 0.01992f
C380 VDD2.n141 B 0.010704f
C381 VDD2.n142 B 0.025301f
C382 VDD2.n143 B 0.011334f
C383 VDD2.n144 B 1.72511f
C384 VDD2.n145 B 0.010704f
C385 VDD2.t1 B 0.042039f
C386 VDD2.n146 B 0.153397f
C387 VDD2.n147 B 0.014946f
C388 VDD2.n148 B 0.018976f
C389 VDD2.n149 B 0.025301f
C390 VDD2.n150 B 0.011334f
C391 VDD2.n151 B 0.010704f
C392 VDD2.n152 B 0.01992f
C393 VDD2.n153 B 0.01992f
C394 VDD2.n154 B 0.010704f
C395 VDD2.n155 B 0.011334f
C396 VDD2.n156 B 0.025301f
C397 VDD2.n157 B 0.025301f
C398 VDD2.n158 B 0.011334f
C399 VDD2.n159 B 0.010704f
C400 VDD2.n160 B 0.01992f
C401 VDD2.n161 B 0.01992f
C402 VDD2.n162 B 0.010704f
C403 VDD2.n163 B 0.011334f
C404 VDD2.n164 B 0.025301f
C405 VDD2.n165 B 0.025301f
C406 VDD2.n166 B 0.011334f
C407 VDD2.n167 B 0.010704f
C408 VDD2.n168 B 0.01992f
C409 VDD2.n169 B 0.01992f
C410 VDD2.n170 B 0.010704f
C411 VDD2.n171 B 0.011334f
C412 VDD2.n172 B 0.025301f
C413 VDD2.n173 B 0.025301f
C414 VDD2.n174 B 0.011334f
C415 VDD2.n175 B 0.010704f
C416 VDD2.n176 B 0.01992f
C417 VDD2.n177 B 0.01992f
C418 VDD2.n178 B 0.010704f
C419 VDD2.n179 B 0.011334f
C420 VDD2.n180 B 0.025301f
C421 VDD2.n181 B 0.025301f
C422 VDD2.n182 B 0.011334f
C423 VDD2.n183 B 0.010704f
C424 VDD2.n184 B 0.01992f
C425 VDD2.n185 B 0.01992f
C426 VDD2.n186 B 0.010704f
C427 VDD2.n187 B 0.011334f
C428 VDD2.n188 B 0.025301f
C429 VDD2.n189 B 0.025301f
C430 VDD2.n190 B 0.011334f
C431 VDD2.n191 B 0.010704f
C432 VDD2.n192 B 0.01992f
C433 VDD2.n193 B 0.01992f
C434 VDD2.n194 B 0.010704f
C435 VDD2.n195 B 0.011334f
C436 VDD2.n196 B 0.025301f
C437 VDD2.n197 B 0.025301f
C438 VDD2.n198 B 0.011334f
C439 VDD2.n199 B 0.010704f
C440 VDD2.n200 B 0.01992f
C441 VDD2.n201 B 0.01992f
C442 VDD2.n202 B 0.010704f
C443 VDD2.n203 B 0.011334f
C444 VDD2.n204 B 0.025301f
C445 VDD2.n205 B 0.025301f
C446 VDD2.n206 B 0.011334f
C447 VDD2.n207 B 0.010704f
C448 VDD2.n208 B 0.01992f
C449 VDD2.n209 B 0.01992f
C450 VDD2.n210 B 0.010704f
C451 VDD2.n211 B 0.011334f
C452 VDD2.n212 B 0.025301f
C453 VDD2.n213 B 0.057149f
C454 VDD2.n214 B 0.011334f
C455 VDD2.n215 B 0.010704f
C456 VDD2.n216 B 0.046589f
C457 VDD2.n217 B 0.045988f
C458 VDD2.n218 B 3.1249f
C459 VTAIL.n0 B 0.029023f
C460 VTAIL.n1 B 0.019702f
C461 VTAIL.n2 B 0.010587f
C462 VTAIL.n3 B 0.025024f
C463 VTAIL.n4 B 0.01121f
C464 VTAIL.n5 B 0.019702f
C465 VTAIL.n6 B 0.010587f
C466 VTAIL.n7 B 0.025024f
C467 VTAIL.n8 B 0.01121f
C468 VTAIL.n9 B 0.019702f
C469 VTAIL.n10 B 0.010587f
C470 VTAIL.n11 B 0.025024f
C471 VTAIL.n12 B 0.010899f
C472 VTAIL.n13 B 0.019702f
C473 VTAIL.n14 B 0.01121f
C474 VTAIL.n15 B 0.025024f
C475 VTAIL.n16 B 0.01121f
C476 VTAIL.n17 B 0.019702f
C477 VTAIL.n18 B 0.010587f
C478 VTAIL.n19 B 0.025024f
C479 VTAIL.n20 B 0.01121f
C480 VTAIL.n21 B 0.019702f
C481 VTAIL.n22 B 0.010587f
C482 VTAIL.n23 B 0.025024f
C483 VTAIL.n24 B 0.01121f
C484 VTAIL.n25 B 0.019702f
C485 VTAIL.n26 B 0.010587f
C486 VTAIL.n27 B 0.025024f
C487 VTAIL.n28 B 0.01121f
C488 VTAIL.n29 B 0.019702f
C489 VTAIL.n30 B 0.010587f
C490 VTAIL.n31 B 0.025024f
C491 VTAIL.n32 B 0.01121f
C492 VTAIL.n33 B 1.70626f
C493 VTAIL.n34 B 0.010587f
C494 VTAIL.t0 B 0.04158f
C495 VTAIL.n35 B 0.15172f
C496 VTAIL.n36 B 0.014783f
C497 VTAIL.n37 B 0.018768f
C498 VTAIL.n38 B 0.025024f
C499 VTAIL.n39 B 0.01121f
C500 VTAIL.n40 B 0.010587f
C501 VTAIL.n41 B 0.019702f
C502 VTAIL.n42 B 0.019702f
C503 VTAIL.n43 B 0.010587f
C504 VTAIL.n44 B 0.01121f
C505 VTAIL.n45 B 0.025024f
C506 VTAIL.n46 B 0.025024f
C507 VTAIL.n47 B 0.01121f
C508 VTAIL.n48 B 0.010587f
C509 VTAIL.n49 B 0.019702f
C510 VTAIL.n50 B 0.019702f
C511 VTAIL.n51 B 0.010587f
C512 VTAIL.n52 B 0.01121f
C513 VTAIL.n53 B 0.025024f
C514 VTAIL.n54 B 0.025024f
C515 VTAIL.n55 B 0.01121f
C516 VTAIL.n56 B 0.010587f
C517 VTAIL.n57 B 0.019702f
C518 VTAIL.n58 B 0.019702f
C519 VTAIL.n59 B 0.010587f
C520 VTAIL.n60 B 0.01121f
C521 VTAIL.n61 B 0.025024f
C522 VTAIL.n62 B 0.025024f
C523 VTAIL.n63 B 0.01121f
C524 VTAIL.n64 B 0.010587f
C525 VTAIL.n65 B 0.019702f
C526 VTAIL.n66 B 0.019702f
C527 VTAIL.n67 B 0.010587f
C528 VTAIL.n68 B 0.01121f
C529 VTAIL.n69 B 0.025024f
C530 VTAIL.n70 B 0.025024f
C531 VTAIL.n71 B 0.01121f
C532 VTAIL.n72 B 0.010587f
C533 VTAIL.n73 B 0.019702f
C534 VTAIL.n74 B 0.019702f
C535 VTAIL.n75 B 0.010587f
C536 VTAIL.n76 B 0.010587f
C537 VTAIL.n77 B 0.01121f
C538 VTAIL.n78 B 0.025024f
C539 VTAIL.n79 B 0.025024f
C540 VTAIL.n80 B 0.025024f
C541 VTAIL.n81 B 0.010899f
C542 VTAIL.n82 B 0.010587f
C543 VTAIL.n83 B 0.019702f
C544 VTAIL.n84 B 0.019702f
C545 VTAIL.n85 B 0.010587f
C546 VTAIL.n86 B 0.01121f
C547 VTAIL.n87 B 0.025024f
C548 VTAIL.n88 B 0.025024f
C549 VTAIL.n89 B 0.01121f
C550 VTAIL.n90 B 0.010587f
C551 VTAIL.n91 B 0.019702f
C552 VTAIL.n92 B 0.019702f
C553 VTAIL.n93 B 0.010587f
C554 VTAIL.n94 B 0.01121f
C555 VTAIL.n95 B 0.025024f
C556 VTAIL.n96 B 0.025024f
C557 VTAIL.n97 B 0.01121f
C558 VTAIL.n98 B 0.010587f
C559 VTAIL.n99 B 0.019702f
C560 VTAIL.n100 B 0.019702f
C561 VTAIL.n101 B 0.010587f
C562 VTAIL.n102 B 0.01121f
C563 VTAIL.n103 B 0.025024f
C564 VTAIL.n104 B 0.056524f
C565 VTAIL.n105 B 0.01121f
C566 VTAIL.n106 B 0.010587f
C567 VTAIL.n107 B 0.046079f
C568 VTAIL.n108 B 0.031886f
C569 VTAIL.n109 B 1.81389f
C570 VTAIL.n110 B 0.029023f
C571 VTAIL.n111 B 0.019702f
C572 VTAIL.n112 B 0.010587f
C573 VTAIL.n113 B 0.025024f
C574 VTAIL.n114 B 0.01121f
C575 VTAIL.n115 B 0.019702f
C576 VTAIL.n116 B 0.010587f
C577 VTAIL.n117 B 0.025024f
C578 VTAIL.n118 B 0.01121f
C579 VTAIL.n119 B 0.019702f
C580 VTAIL.n120 B 0.010587f
C581 VTAIL.n121 B 0.025024f
C582 VTAIL.n122 B 0.010899f
C583 VTAIL.n123 B 0.019702f
C584 VTAIL.n124 B 0.010899f
C585 VTAIL.n125 B 0.010587f
C586 VTAIL.n126 B 0.025024f
C587 VTAIL.n127 B 0.025024f
C588 VTAIL.n128 B 0.01121f
C589 VTAIL.n129 B 0.019702f
C590 VTAIL.n130 B 0.010587f
C591 VTAIL.n131 B 0.025024f
C592 VTAIL.n132 B 0.01121f
C593 VTAIL.n133 B 0.019702f
C594 VTAIL.n134 B 0.010587f
C595 VTAIL.n135 B 0.025024f
C596 VTAIL.n136 B 0.01121f
C597 VTAIL.n137 B 0.019702f
C598 VTAIL.n138 B 0.010587f
C599 VTAIL.n139 B 0.025024f
C600 VTAIL.n140 B 0.01121f
C601 VTAIL.n141 B 0.019702f
C602 VTAIL.n142 B 0.010587f
C603 VTAIL.n143 B 0.025024f
C604 VTAIL.n144 B 0.01121f
C605 VTAIL.n145 B 1.70626f
C606 VTAIL.n146 B 0.010587f
C607 VTAIL.t2 B 0.04158f
C608 VTAIL.n147 B 0.15172f
C609 VTAIL.n148 B 0.014783f
C610 VTAIL.n149 B 0.018768f
C611 VTAIL.n150 B 0.025024f
C612 VTAIL.n151 B 0.01121f
C613 VTAIL.n152 B 0.010587f
C614 VTAIL.n153 B 0.019702f
C615 VTAIL.n154 B 0.019702f
C616 VTAIL.n155 B 0.010587f
C617 VTAIL.n156 B 0.01121f
C618 VTAIL.n157 B 0.025024f
C619 VTAIL.n158 B 0.025024f
C620 VTAIL.n159 B 0.01121f
C621 VTAIL.n160 B 0.010587f
C622 VTAIL.n161 B 0.019702f
C623 VTAIL.n162 B 0.019702f
C624 VTAIL.n163 B 0.010587f
C625 VTAIL.n164 B 0.01121f
C626 VTAIL.n165 B 0.025024f
C627 VTAIL.n166 B 0.025024f
C628 VTAIL.n167 B 0.01121f
C629 VTAIL.n168 B 0.010587f
C630 VTAIL.n169 B 0.019702f
C631 VTAIL.n170 B 0.019702f
C632 VTAIL.n171 B 0.010587f
C633 VTAIL.n172 B 0.01121f
C634 VTAIL.n173 B 0.025024f
C635 VTAIL.n174 B 0.025024f
C636 VTAIL.n175 B 0.01121f
C637 VTAIL.n176 B 0.010587f
C638 VTAIL.n177 B 0.019702f
C639 VTAIL.n178 B 0.019702f
C640 VTAIL.n179 B 0.010587f
C641 VTAIL.n180 B 0.01121f
C642 VTAIL.n181 B 0.025024f
C643 VTAIL.n182 B 0.025024f
C644 VTAIL.n183 B 0.01121f
C645 VTAIL.n184 B 0.010587f
C646 VTAIL.n185 B 0.019702f
C647 VTAIL.n186 B 0.019702f
C648 VTAIL.n187 B 0.010587f
C649 VTAIL.n188 B 0.01121f
C650 VTAIL.n189 B 0.025024f
C651 VTAIL.n190 B 0.025024f
C652 VTAIL.n191 B 0.01121f
C653 VTAIL.n192 B 0.010587f
C654 VTAIL.n193 B 0.019702f
C655 VTAIL.n194 B 0.019702f
C656 VTAIL.n195 B 0.010587f
C657 VTAIL.n196 B 0.01121f
C658 VTAIL.n197 B 0.025024f
C659 VTAIL.n198 B 0.025024f
C660 VTAIL.n199 B 0.01121f
C661 VTAIL.n200 B 0.010587f
C662 VTAIL.n201 B 0.019702f
C663 VTAIL.n202 B 0.019702f
C664 VTAIL.n203 B 0.010587f
C665 VTAIL.n204 B 0.01121f
C666 VTAIL.n205 B 0.025024f
C667 VTAIL.n206 B 0.025024f
C668 VTAIL.n207 B 0.01121f
C669 VTAIL.n208 B 0.010587f
C670 VTAIL.n209 B 0.019702f
C671 VTAIL.n210 B 0.019702f
C672 VTAIL.n211 B 0.010587f
C673 VTAIL.n212 B 0.01121f
C674 VTAIL.n213 B 0.025024f
C675 VTAIL.n214 B 0.056524f
C676 VTAIL.n215 B 0.01121f
C677 VTAIL.n216 B 0.010587f
C678 VTAIL.n217 B 0.046079f
C679 VTAIL.n218 B 0.031886f
C680 VTAIL.n219 B 1.85658f
C681 VTAIL.n220 B 0.029023f
C682 VTAIL.n221 B 0.019702f
C683 VTAIL.n222 B 0.010587f
C684 VTAIL.n223 B 0.025024f
C685 VTAIL.n224 B 0.01121f
C686 VTAIL.n225 B 0.019702f
C687 VTAIL.n226 B 0.010587f
C688 VTAIL.n227 B 0.025024f
C689 VTAIL.n228 B 0.01121f
C690 VTAIL.n229 B 0.019702f
C691 VTAIL.n230 B 0.010587f
C692 VTAIL.n231 B 0.025024f
C693 VTAIL.n232 B 0.010899f
C694 VTAIL.n233 B 0.019702f
C695 VTAIL.n234 B 0.010899f
C696 VTAIL.n235 B 0.010587f
C697 VTAIL.n236 B 0.025024f
C698 VTAIL.n237 B 0.025024f
C699 VTAIL.n238 B 0.01121f
C700 VTAIL.n239 B 0.019702f
C701 VTAIL.n240 B 0.010587f
C702 VTAIL.n241 B 0.025024f
C703 VTAIL.n242 B 0.01121f
C704 VTAIL.n243 B 0.019702f
C705 VTAIL.n244 B 0.010587f
C706 VTAIL.n245 B 0.025024f
C707 VTAIL.n246 B 0.01121f
C708 VTAIL.n247 B 0.019702f
C709 VTAIL.n248 B 0.010587f
C710 VTAIL.n249 B 0.025024f
C711 VTAIL.n250 B 0.01121f
C712 VTAIL.n251 B 0.019702f
C713 VTAIL.n252 B 0.010587f
C714 VTAIL.n253 B 0.025024f
C715 VTAIL.n254 B 0.01121f
C716 VTAIL.n255 B 1.70626f
C717 VTAIL.n256 B 0.010587f
C718 VTAIL.t1 B 0.04158f
C719 VTAIL.n257 B 0.15172f
C720 VTAIL.n258 B 0.014783f
C721 VTAIL.n259 B 0.018768f
C722 VTAIL.n260 B 0.025024f
C723 VTAIL.n261 B 0.01121f
C724 VTAIL.n262 B 0.010587f
C725 VTAIL.n263 B 0.019702f
C726 VTAIL.n264 B 0.019702f
C727 VTAIL.n265 B 0.010587f
C728 VTAIL.n266 B 0.01121f
C729 VTAIL.n267 B 0.025024f
C730 VTAIL.n268 B 0.025024f
C731 VTAIL.n269 B 0.01121f
C732 VTAIL.n270 B 0.010587f
C733 VTAIL.n271 B 0.019702f
C734 VTAIL.n272 B 0.019702f
C735 VTAIL.n273 B 0.010587f
C736 VTAIL.n274 B 0.01121f
C737 VTAIL.n275 B 0.025024f
C738 VTAIL.n276 B 0.025024f
C739 VTAIL.n277 B 0.01121f
C740 VTAIL.n278 B 0.010587f
C741 VTAIL.n279 B 0.019702f
C742 VTAIL.n280 B 0.019702f
C743 VTAIL.n281 B 0.010587f
C744 VTAIL.n282 B 0.01121f
C745 VTAIL.n283 B 0.025024f
C746 VTAIL.n284 B 0.025024f
C747 VTAIL.n285 B 0.01121f
C748 VTAIL.n286 B 0.010587f
C749 VTAIL.n287 B 0.019702f
C750 VTAIL.n288 B 0.019702f
C751 VTAIL.n289 B 0.010587f
C752 VTAIL.n290 B 0.01121f
C753 VTAIL.n291 B 0.025024f
C754 VTAIL.n292 B 0.025024f
C755 VTAIL.n293 B 0.01121f
C756 VTAIL.n294 B 0.010587f
C757 VTAIL.n295 B 0.019702f
C758 VTAIL.n296 B 0.019702f
C759 VTAIL.n297 B 0.010587f
C760 VTAIL.n298 B 0.01121f
C761 VTAIL.n299 B 0.025024f
C762 VTAIL.n300 B 0.025024f
C763 VTAIL.n301 B 0.01121f
C764 VTAIL.n302 B 0.010587f
C765 VTAIL.n303 B 0.019702f
C766 VTAIL.n304 B 0.019702f
C767 VTAIL.n305 B 0.010587f
C768 VTAIL.n306 B 0.01121f
C769 VTAIL.n307 B 0.025024f
C770 VTAIL.n308 B 0.025024f
C771 VTAIL.n309 B 0.01121f
C772 VTAIL.n310 B 0.010587f
C773 VTAIL.n311 B 0.019702f
C774 VTAIL.n312 B 0.019702f
C775 VTAIL.n313 B 0.010587f
C776 VTAIL.n314 B 0.01121f
C777 VTAIL.n315 B 0.025024f
C778 VTAIL.n316 B 0.025024f
C779 VTAIL.n317 B 0.01121f
C780 VTAIL.n318 B 0.010587f
C781 VTAIL.n319 B 0.019702f
C782 VTAIL.n320 B 0.019702f
C783 VTAIL.n321 B 0.010587f
C784 VTAIL.n322 B 0.01121f
C785 VTAIL.n323 B 0.025024f
C786 VTAIL.n324 B 0.056524f
C787 VTAIL.n325 B 0.01121f
C788 VTAIL.n326 B 0.010587f
C789 VTAIL.n327 B 0.046079f
C790 VTAIL.n328 B 0.031886f
C791 VTAIL.n329 B 1.67105f
C792 VTAIL.n330 B 0.029023f
C793 VTAIL.n331 B 0.019702f
C794 VTAIL.n332 B 0.010587f
C795 VTAIL.n333 B 0.025024f
C796 VTAIL.n334 B 0.01121f
C797 VTAIL.n335 B 0.019702f
C798 VTAIL.n336 B 0.010587f
C799 VTAIL.n337 B 0.025024f
C800 VTAIL.n338 B 0.01121f
C801 VTAIL.n339 B 0.019702f
C802 VTAIL.n340 B 0.010587f
C803 VTAIL.n341 B 0.025024f
C804 VTAIL.n342 B 0.010899f
C805 VTAIL.n343 B 0.019702f
C806 VTAIL.n344 B 0.01121f
C807 VTAIL.n345 B 0.025024f
C808 VTAIL.n346 B 0.01121f
C809 VTAIL.n347 B 0.019702f
C810 VTAIL.n348 B 0.010587f
C811 VTAIL.n349 B 0.025024f
C812 VTAIL.n350 B 0.01121f
C813 VTAIL.n351 B 0.019702f
C814 VTAIL.n352 B 0.010587f
C815 VTAIL.n353 B 0.025024f
C816 VTAIL.n354 B 0.01121f
C817 VTAIL.n355 B 0.019702f
C818 VTAIL.n356 B 0.010587f
C819 VTAIL.n357 B 0.025024f
C820 VTAIL.n358 B 0.01121f
C821 VTAIL.n359 B 0.019702f
C822 VTAIL.n360 B 0.010587f
C823 VTAIL.n361 B 0.025024f
C824 VTAIL.n362 B 0.01121f
C825 VTAIL.n363 B 1.70626f
C826 VTAIL.n364 B 0.010587f
C827 VTAIL.t3 B 0.04158f
C828 VTAIL.n365 B 0.15172f
C829 VTAIL.n366 B 0.014783f
C830 VTAIL.n367 B 0.018768f
C831 VTAIL.n368 B 0.025024f
C832 VTAIL.n369 B 0.01121f
C833 VTAIL.n370 B 0.010587f
C834 VTAIL.n371 B 0.019702f
C835 VTAIL.n372 B 0.019702f
C836 VTAIL.n373 B 0.010587f
C837 VTAIL.n374 B 0.01121f
C838 VTAIL.n375 B 0.025024f
C839 VTAIL.n376 B 0.025024f
C840 VTAIL.n377 B 0.01121f
C841 VTAIL.n378 B 0.010587f
C842 VTAIL.n379 B 0.019702f
C843 VTAIL.n380 B 0.019702f
C844 VTAIL.n381 B 0.010587f
C845 VTAIL.n382 B 0.01121f
C846 VTAIL.n383 B 0.025024f
C847 VTAIL.n384 B 0.025024f
C848 VTAIL.n385 B 0.01121f
C849 VTAIL.n386 B 0.010587f
C850 VTAIL.n387 B 0.019702f
C851 VTAIL.n388 B 0.019702f
C852 VTAIL.n389 B 0.010587f
C853 VTAIL.n390 B 0.01121f
C854 VTAIL.n391 B 0.025024f
C855 VTAIL.n392 B 0.025024f
C856 VTAIL.n393 B 0.01121f
C857 VTAIL.n394 B 0.010587f
C858 VTAIL.n395 B 0.019702f
C859 VTAIL.n396 B 0.019702f
C860 VTAIL.n397 B 0.010587f
C861 VTAIL.n398 B 0.01121f
C862 VTAIL.n399 B 0.025024f
C863 VTAIL.n400 B 0.025024f
C864 VTAIL.n401 B 0.01121f
C865 VTAIL.n402 B 0.010587f
C866 VTAIL.n403 B 0.019702f
C867 VTAIL.n404 B 0.019702f
C868 VTAIL.n405 B 0.010587f
C869 VTAIL.n406 B 0.010587f
C870 VTAIL.n407 B 0.01121f
C871 VTAIL.n408 B 0.025024f
C872 VTAIL.n409 B 0.025024f
C873 VTAIL.n410 B 0.025024f
C874 VTAIL.n411 B 0.010899f
C875 VTAIL.n412 B 0.010587f
C876 VTAIL.n413 B 0.019702f
C877 VTAIL.n414 B 0.019702f
C878 VTAIL.n415 B 0.010587f
C879 VTAIL.n416 B 0.01121f
C880 VTAIL.n417 B 0.025024f
C881 VTAIL.n418 B 0.025024f
C882 VTAIL.n419 B 0.01121f
C883 VTAIL.n420 B 0.010587f
C884 VTAIL.n421 B 0.019702f
C885 VTAIL.n422 B 0.019702f
C886 VTAIL.n423 B 0.010587f
C887 VTAIL.n424 B 0.01121f
C888 VTAIL.n425 B 0.025024f
C889 VTAIL.n426 B 0.025024f
C890 VTAIL.n427 B 0.01121f
C891 VTAIL.n428 B 0.010587f
C892 VTAIL.n429 B 0.019702f
C893 VTAIL.n430 B 0.019702f
C894 VTAIL.n431 B 0.010587f
C895 VTAIL.n432 B 0.01121f
C896 VTAIL.n433 B 0.025024f
C897 VTAIL.n434 B 0.056524f
C898 VTAIL.n435 B 0.01121f
C899 VTAIL.n436 B 0.010587f
C900 VTAIL.n437 B 0.046079f
C901 VTAIL.n438 B 0.031886f
C902 VTAIL.n439 B 1.59114f
C903 VN.t1 B 4.72333f
C904 VN.t0 B 5.34726f
.ends

