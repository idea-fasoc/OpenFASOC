* NGSPICE file created from diff_pair_sample_0228.ext - technology: sky130A

.subckt diff_pair_sample_0228 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1898_n3346# sky130_fd_pr__pfet_01v8 ad=4.6371 pd=24.56 as=0 ps=0 w=11.89 l=1.99
X1 B.t8 B.t6 B.t7 w_n1898_n3346# sky130_fd_pr__pfet_01v8 ad=4.6371 pd=24.56 as=0 ps=0 w=11.89 l=1.99
X2 VDD2.t1 VN.t0 VTAIL.t3 w_n1898_n3346# sky130_fd_pr__pfet_01v8 ad=4.6371 pd=24.56 as=4.6371 ps=24.56 w=11.89 l=1.99
X3 VDD2.t0 VN.t1 VTAIL.t2 w_n1898_n3346# sky130_fd_pr__pfet_01v8 ad=4.6371 pd=24.56 as=4.6371 ps=24.56 w=11.89 l=1.99
X4 B.t5 B.t3 B.t4 w_n1898_n3346# sky130_fd_pr__pfet_01v8 ad=4.6371 pd=24.56 as=0 ps=0 w=11.89 l=1.99
X5 VDD1.t1 VP.t0 VTAIL.t0 w_n1898_n3346# sky130_fd_pr__pfet_01v8 ad=4.6371 pd=24.56 as=4.6371 ps=24.56 w=11.89 l=1.99
X6 VDD1.t0 VP.t1 VTAIL.t1 w_n1898_n3346# sky130_fd_pr__pfet_01v8 ad=4.6371 pd=24.56 as=4.6371 ps=24.56 w=11.89 l=1.99
X7 B.t2 B.t0 B.t1 w_n1898_n3346# sky130_fd_pr__pfet_01v8 ad=4.6371 pd=24.56 as=0 ps=0 w=11.89 l=1.99
R0 B.n314 B.n85 585
R1 B.n313 B.n312 585
R2 B.n311 B.n86 585
R3 B.n310 B.n309 585
R4 B.n308 B.n87 585
R5 B.n307 B.n306 585
R6 B.n305 B.n88 585
R7 B.n304 B.n303 585
R8 B.n302 B.n89 585
R9 B.n301 B.n300 585
R10 B.n299 B.n90 585
R11 B.n298 B.n297 585
R12 B.n296 B.n91 585
R13 B.n295 B.n294 585
R14 B.n293 B.n92 585
R15 B.n292 B.n291 585
R16 B.n290 B.n93 585
R17 B.n289 B.n288 585
R18 B.n287 B.n94 585
R19 B.n286 B.n285 585
R20 B.n284 B.n95 585
R21 B.n283 B.n282 585
R22 B.n281 B.n96 585
R23 B.n280 B.n279 585
R24 B.n278 B.n97 585
R25 B.n277 B.n276 585
R26 B.n275 B.n98 585
R27 B.n274 B.n273 585
R28 B.n272 B.n99 585
R29 B.n271 B.n270 585
R30 B.n269 B.n100 585
R31 B.n268 B.n267 585
R32 B.n266 B.n101 585
R33 B.n265 B.n264 585
R34 B.n263 B.n102 585
R35 B.n262 B.n261 585
R36 B.n260 B.n103 585
R37 B.n259 B.n258 585
R38 B.n257 B.n104 585
R39 B.n256 B.n255 585
R40 B.n254 B.n105 585
R41 B.n252 B.n251 585
R42 B.n250 B.n108 585
R43 B.n249 B.n248 585
R44 B.n247 B.n109 585
R45 B.n246 B.n245 585
R46 B.n244 B.n110 585
R47 B.n243 B.n242 585
R48 B.n241 B.n111 585
R49 B.n240 B.n239 585
R50 B.n238 B.n112 585
R51 B.n237 B.n236 585
R52 B.n232 B.n113 585
R53 B.n231 B.n230 585
R54 B.n229 B.n114 585
R55 B.n228 B.n227 585
R56 B.n226 B.n115 585
R57 B.n225 B.n224 585
R58 B.n223 B.n116 585
R59 B.n222 B.n221 585
R60 B.n220 B.n117 585
R61 B.n219 B.n218 585
R62 B.n217 B.n118 585
R63 B.n216 B.n215 585
R64 B.n214 B.n119 585
R65 B.n213 B.n212 585
R66 B.n211 B.n120 585
R67 B.n210 B.n209 585
R68 B.n208 B.n121 585
R69 B.n207 B.n206 585
R70 B.n205 B.n122 585
R71 B.n204 B.n203 585
R72 B.n202 B.n123 585
R73 B.n201 B.n200 585
R74 B.n199 B.n124 585
R75 B.n198 B.n197 585
R76 B.n196 B.n125 585
R77 B.n195 B.n194 585
R78 B.n193 B.n126 585
R79 B.n192 B.n191 585
R80 B.n190 B.n127 585
R81 B.n189 B.n188 585
R82 B.n187 B.n128 585
R83 B.n186 B.n185 585
R84 B.n184 B.n129 585
R85 B.n183 B.n182 585
R86 B.n181 B.n130 585
R87 B.n180 B.n179 585
R88 B.n178 B.n131 585
R89 B.n177 B.n176 585
R90 B.n175 B.n132 585
R91 B.n174 B.n173 585
R92 B.n316 B.n315 585
R93 B.n317 B.n84 585
R94 B.n319 B.n318 585
R95 B.n320 B.n83 585
R96 B.n322 B.n321 585
R97 B.n323 B.n82 585
R98 B.n325 B.n324 585
R99 B.n326 B.n81 585
R100 B.n328 B.n327 585
R101 B.n329 B.n80 585
R102 B.n331 B.n330 585
R103 B.n332 B.n79 585
R104 B.n334 B.n333 585
R105 B.n335 B.n78 585
R106 B.n337 B.n336 585
R107 B.n338 B.n77 585
R108 B.n340 B.n339 585
R109 B.n341 B.n76 585
R110 B.n343 B.n342 585
R111 B.n344 B.n75 585
R112 B.n346 B.n345 585
R113 B.n347 B.n74 585
R114 B.n349 B.n348 585
R115 B.n350 B.n73 585
R116 B.n352 B.n351 585
R117 B.n353 B.n72 585
R118 B.n355 B.n354 585
R119 B.n356 B.n71 585
R120 B.n358 B.n357 585
R121 B.n359 B.n70 585
R122 B.n361 B.n360 585
R123 B.n362 B.n69 585
R124 B.n364 B.n363 585
R125 B.n365 B.n68 585
R126 B.n367 B.n366 585
R127 B.n368 B.n67 585
R128 B.n370 B.n369 585
R129 B.n371 B.n66 585
R130 B.n373 B.n372 585
R131 B.n374 B.n65 585
R132 B.n376 B.n375 585
R133 B.n377 B.n64 585
R134 B.n379 B.n378 585
R135 B.n380 B.n63 585
R136 B.n520 B.n519 585
R137 B.n518 B.n13 585
R138 B.n517 B.n516 585
R139 B.n515 B.n14 585
R140 B.n514 B.n513 585
R141 B.n512 B.n15 585
R142 B.n511 B.n510 585
R143 B.n509 B.n16 585
R144 B.n508 B.n507 585
R145 B.n506 B.n17 585
R146 B.n505 B.n504 585
R147 B.n503 B.n18 585
R148 B.n502 B.n501 585
R149 B.n500 B.n19 585
R150 B.n499 B.n498 585
R151 B.n497 B.n20 585
R152 B.n496 B.n495 585
R153 B.n494 B.n21 585
R154 B.n493 B.n492 585
R155 B.n491 B.n22 585
R156 B.n490 B.n489 585
R157 B.n488 B.n23 585
R158 B.n487 B.n486 585
R159 B.n485 B.n24 585
R160 B.n484 B.n483 585
R161 B.n482 B.n25 585
R162 B.n481 B.n480 585
R163 B.n479 B.n26 585
R164 B.n478 B.n477 585
R165 B.n476 B.n27 585
R166 B.n475 B.n474 585
R167 B.n473 B.n28 585
R168 B.n472 B.n471 585
R169 B.n470 B.n29 585
R170 B.n469 B.n468 585
R171 B.n467 B.n30 585
R172 B.n466 B.n465 585
R173 B.n464 B.n31 585
R174 B.n463 B.n462 585
R175 B.n461 B.n32 585
R176 B.n460 B.n459 585
R177 B.n457 B.n33 585
R178 B.n456 B.n455 585
R179 B.n454 B.n36 585
R180 B.n453 B.n452 585
R181 B.n451 B.n37 585
R182 B.n450 B.n449 585
R183 B.n448 B.n38 585
R184 B.n447 B.n446 585
R185 B.n445 B.n39 585
R186 B.n444 B.n443 585
R187 B.n442 B.n441 585
R188 B.n440 B.n43 585
R189 B.n439 B.n438 585
R190 B.n437 B.n44 585
R191 B.n436 B.n435 585
R192 B.n434 B.n45 585
R193 B.n433 B.n432 585
R194 B.n431 B.n46 585
R195 B.n430 B.n429 585
R196 B.n428 B.n47 585
R197 B.n427 B.n426 585
R198 B.n425 B.n48 585
R199 B.n424 B.n423 585
R200 B.n422 B.n49 585
R201 B.n421 B.n420 585
R202 B.n419 B.n50 585
R203 B.n418 B.n417 585
R204 B.n416 B.n51 585
R205 B.n415 B.n414 585
R206 B.n413 B.n52 585
R207 B.n412 B.n411 585
R208 B.n410 B.n53 585
R209 B.n409 B.n408 585
R210 B.n407 B.n54 585
R211 B.n406 B.n405 585
R212 B.n404 B.n55 585
R213 B.n403 B.n402 585
R214 B.n401 B.n56 585
R215 B.n400 B.n399 585
R216 B.n398 B.n57 585
R217 B.n397 B.n396 585
R218 B.n395 B.n58 585
R219 B.n394 B.n393 585
R220 B.n392 B.n59 585
R221 B.n391 B.n390 585
R222 B.n389 B.n60 585
R223 B.n388 B.n387 585
R224 B.n386 B.n61 585
R225 B.n385 B.n384 585
R226 B.n383 B.n62 585
R227 B.n382 B.n381 585
R228 B.n521 B.n12 585
R229 B.n523 B.n522 585
R230 B.n524 B.n11 585
R231 B.n526 B.n525 585
R232 B.n527 B.n10 585
R233 B.n529 B.n528 585
R234 B.n530 B.n9 585
R235 B.n532 B.n531 585
R236 B.n533 B.n8 585
R237 B.n535 B.n534 585
R238 B.n536 B.n7 585
R239 B.n538 B.n537 585
R240 B.n539 B.n6 585
R241 B.n541 B.n540 585
R242 B.n542 B.n5 585
R243 B.n544 B.n543 585
R244 B.n545 B.n4 585
R245 B.n547 B.n546 585
R246 B.n548 B.n3 585
R247 B.n550 B.n549 585
R248 B.n551 B.n0 585
R249 B.n2 B.n1 585
R250 B.n144 B.n143 585
R251 B.n145 B.n142 585
R252 B.n147 B.n146 585
R253 B.n148 B.n141 585
R254 B.n150 B.n149 585
R255 B.n151 B.n140 585
R256 B.n153 B.n152 585
R257 B.n154 B.n139 585
R258 B.n156 B.n155 585
R259 B.n157 B.n138 585
R260 B.n159 B.n158 585
R261 B.n160 B.n137 585
R262 B.n162 B.n161 585
R263 B.n163 B.n136 585
R264 B.n165 B.n164 585
R265 B.n166 B.n135 585
R266 B.n168 B.n167 585
R267 B.n169 B.n134 585
R268 B.n171 B.n170 585
R269 B.n172 B.n133 585
R270 B.n174 B.n133 554.963
R271 B.n316 B.n85 554.963
R272 B.n382 B.n63 554.963
R273 B.n521 B.n520 554.963
R274 B.n233 B.t3 350.889
R275 B.n106 B.t6 350.889
R276 B.n40 B.t0 350.889
R277 B.n34 B.t9 350.889
R278 B.n553 B.n552 256.663
R279 B.n552 B.n551 235.042
R280 B.n552 B.n2 235.042
R281 B.n175 B.n174 163.367
R282 B.n176 B.n175 163.367
R283 B.n176 B.n131 163.367
R284 B.n180 B.n131 163.367
R285 B.n181 B.n180 163.367
R286 B.n182 B.n181 163.367
R287 B.n182 B.n129 163.367
R288 B.n186 B.n129 163.367
R289 B.n187 B.n186 163.367
R290 B.n188 B.n187 163.367
R291 B.n188 B.n127 163.367
R292 B.n192 B.n127 163.367
R293 B.n193 B.n192 163.367
R294 B.n194 B.n193 163.367
R295 B.n194 B.n125 163.367
R296 B.n198 B.n125 163.367
R297 B.n199 B.n198 163.367
R298 B.n200 B.n199 163.367
R299 B.n200 B.n123 163.367
R300 B.n204 B.n123 163.367
R301 B.n205 B.n204 163.367
R302 B.n206 B.n205 163.367
R303 B.n206 B.n121 163.367
R304 B.n210 B.n121 163.367
R305 B.n211 B.n210 163.367
R306 B.n212 B.n211 163.367
R307 B.n212 B.n119 163.367
R308 B.n216 B.n119 163.367
R309 B.n217 B.n216 163.367
R310 B.n218 B.n217 163.367
R311 B.n218 B.n117 163.367
R312 B.n222 B.n117 163.367
R313 B.n223 B.n222 163.367
R314 B.n224 B.n223 163.367
R315 B.n224 B.n115 163.367
R316 B.n228 B.n115 163.367
R317 B.n229 B.n228 163.367
R318 B.n230 B.n229 163.367
R319 B.n230 B.n113 163.367
R320 B.n237 B.n113 163.367
R321 B.n238 B.n237 163.367
R322 B.n239 B.n238 163.367
R323 B.n239 B.n111 163.367
R324 B.n243 B.n111 163.367
R325 B.n244 B.n243 163.367
R326 B.n245 B.n244 163.367
R327 B.n245 B.n109 163.367
R328 B.n249 B.n109 163.367
R329 B.n250 B.n249 163.367
R330 B.n251 B.n250 163.367
R331 B.n251 B.n105 163.367
R332 B.n256 B.n105 163.367
R333 B.n257 B.n256 163.367
R334 B.n258 B.n257 163.367
R335 B.n258 B.n103 163.367
R336 B.n262 B.n103 163.367
R337 B.n263 B.n262 163.367
R338 B.n264 B.n263 163.367
R339 B.n264 B.n101 163.367
R340 B.n268 B.n101 163.367
R341 B.n269 B.n268 163.367
R342 B.n270 B.n269 163.367
R343 B.n270 B.n99 163.367
R344 B.n274 B.n99 163.367
R345 B.n275 B.n274 163.367
R346 B.n276 B.n275 163.367
R347 B.n276 B.n97 163.367
R348 B.n280 B.n97 163.367
R349 B.n281 B.n280 163.367
R350 B.n282 B.n281 163.367
R351 B.n282 B.n95 163.367
R352 B.n286 B.n95 163.367
R353 B.n287 B.n286 163.367
R354 B.n288 B.n287 163.367
R355 B.n288 B.n93 163.367
R356 B.n292 B.n93 163.367
R357 B.n293 B.n292 163.367
R358 B.n294 B.n293 163.367
R359 B.n294 B.n91 163.367
R360 B.n298 B.n91 163.367
R361 B.n299 B.n298 163.367
R362 B.n300 B.n299 163.367
R363 B.n300 B.n89 163.367
R364 B.n304 B.n89 163.367
R365 B.n305 B.n304 163.367
R366 B.n306 B.n305 163.367
R367 B.n306 B.n87 163.367
R368 B.n310 B.n87 163.367
R369 B.n311 B.n310 163.367
R370 B.n312 B.n311 163.367
R371 B.n312 B.n85 163.367
R372 B.n378 B.n63 163.367
R373 B.n378 B.n377 163.367
R374 B.n377 B.n376 163.367
R375 B.n376 B.n65 163.367
R376 B.n372 B.n65 163.367
R377 B.n372 B.n371 163.367
R378 B.n371 B.n370 163.367
R379 B.n370 B.n67 163.367
R380 B.n366 B.n67 163.367
R381 B.n366 B.n365 163.367
R382 B.n365 B.n364 163.367
R383 B.n364 B.n69 163.367
R384 B.n360 B.n69 163.367
R385 B.n360 B.n359 163.367
R386 B.n359 B.n358 163.367
R387 B.n358 B.n71 163.367
R388 B.n354 B.n71 163.367
R389 B.n354 B.n353 163.367
R390 B.n353 B.n352 163.367
R391 B.n352 B.n73 163.367
R392 B.n348 B.n73 163.367
R393 B.n348 B.n347 163.367
R394 B.n347 B.n346 163.367
R395 B.n346 B.n75 163.367
R396 B.n342 B.n75 163.367
R397 B.n342 B.n341 163.367
R398 B.n341 B.n340 163.367
R399 B.n340 B.n77 163.367
R400 B.n336 B.n77 163.367
R401 B.n336 B.n335 163.367
R402 B.n335 B.n334 163.367
R403 B.n334 B.n79 163.367
R404 B.n330 B.n79 163.367
R405 B.n330 B.n329 163.367
R406 B.n329 B.n328 163.367
R407 B.n328 B.n81 163.367
R408 B.n324 B.n81 163.367
R409 B.n324 B.n323 163.367
R410 B.n323 B.n322 163.367
R411 B.n322 B.n83 163.367
R412 B.n318 B.n83 163.367
R413 B.n318 B.n317 163.367
R414 B.n317 B.n316 163.367
R415 B.n520 B.n13 163.367
R416 B.n516 B.n13 163.367
R417 B.n516 B.n515 163.367
R418 B.n515 B.n514 163.367
R419 B.n514 B.n15 163.367
R420 B.n510 B.n15 163.367
R421 B.n510 B.n509 163.367
R422 B.n509 B.n508 163.367
R423 B.n508 B.n17 163.367
R424 B.n504 B.n17 163.367
R425 B.n504 B.n503 163.367
R426 B.n503 B.n502 163.367
R427 B.n502 B.n19 163.367
R428 B.n498 B.n19 163.367
R429 B.n498 B.n497 163.367
R430 B.n497 B.n496 163.367
R431 B.n496 B.n21 163.367
R432 B.n492 B.n21 163.367
R433 B.n492 B.n491 163.367
R434 B.n491 B.n490 163.367
R435 B.n490 B.n23 163.367
R436 B.n486 B.n23 163.367
R437 B.n486 B.n485 163.367
R438 B.n485 B.n484 163.367
R439 B.n484 B.n25 163.367
R440 B.n480 B.n25 163.367
R441 B.n480 B.n479 163.367
R442 B.n479 B.n478 163.367
R443 B.n478 B.n27 163.367
R444 B.n474 B.n27 163.367
R445 B.n474 B.n473 163.367
R446 B.n473 B.n472 163.367
R447 B.n472 B.n29 163.367
R448 B.n468 B.n29 163.367
R449 B.n468 B.n467 163.367
R450 B.n467 B.n466 163.367
R451 B.n466 B.n31 163.367
R452 B.n462 B.n31 163.367
R453 B.n462 B.n461 163.367
R454 B.n461 B.n460 163.367
R455 B.n460 B.n33 163.367
R456 B.n455 B.n33 163.367
R457 B.n455 B.n454 163.367
R458 B.n454 B.n453 163.367
R459 B.n453 B.n37 163.367
R460 B.n449 B.n37 163.367
R461 B.n449 B.n448 163.367
R462 B.n448 B.n447 163.367
R463 B.n447 B.n39 163.367
R464 B.n443 B.n39 163.367
R465 B.n443 B.n442 163.367
R466 B.n442 B.n43 163.367
R467 B.n438 B.n43 163.367
R468 B.n438 B.n437 163.367
R469 B.n437 B.n436 163.367
R470 B.n436 B.n45 163.367
R471 B.n432 B.n45 163.367
R472 B.n432 B.n431 163.367
R473 B.n431 B.n430 163.367
R474 B.n430 B.n47 163.367
R475 B.n426 B.n47 163.367
R476 B.n426 B.n425 163.367
R477 B.n425 B.n424 163.367
R478 B.n424 B.n49 163.367
R479 B.n420 B.n49 163.367
R480 B.n420 B.n419 163.367
R481 B.n419 B.n418 163.367
R482 B.n418 B.n51 163.367
R483 B.n414 B.n51 163.367
R484 B.n414 B.n413 163.367
R485 B.n413 B.n412 163.367
R486 B.n412 B.n53 163.367
R487 B.n408 B.n53 163.367
R488 B.n408 B.n407 163.367
R489 B.n407 B.n406 163.367
R490 B.n406 B.n55 163.367
R491 B.n402 B.n55 163.367
R492 B.n402 B.n401 163.367
R493 B.n401 B.n400 163.367
R494 B.n400 B.n57 163.367
R495 B.n396 B.n57 163.367
R496 B.n396 B.n395 163.367
R497 B.n395 B.n394 163.367
R498 B.n394 B.n59 163.367
R499 B.n390 B.n59 163.367
R500 B.n390 B.n389 163.367
R501 B.n389 B.n388 163.367
R502 B.n388 B.n61 163.367
R503 B.n384 B.n61 163.367
R504 B.n384 B.n383 163.367
R505 B.n383 B.n382 163.367
R506 B.n522 B.n521 163.367
R507 B.n522 B.n11 163.367
R508 B.n526 B.n11 163.367
R509 B.n527 B.n526 163.367
R510 B.n528 B.n527 163.367
R511 B.n528 B.n9 163.367
R512 B.n532 B.n9 163.367
R513 B.n533 B.n532 163.367
R514 B.n534 B.n533 163.367
R515 B.n534 B.n7 163.367
R516 B.n538 B.n7 163.367
R517 B.n539 B.n538 163.367
R518 B.n540 B.n539 163.367
R519 B.n540 B.n5 163.367
R520 B.n544 B.n5 163.367
R521 B.n545 B.n544 163.367
R522 B.n546 B.n545 163.367
R523 B.n546 B.n3 163.367
R524 B.n550 B.n3 163.367
R525 B.n551 B.n550 163.367
R526 B.n144 B.n2 163.367
R527 B.n145 B.n144 163.367
R528 B.n146 B.n145 163.367
R529 B.n146 B.n141 163.367
R530 B.n150 B.n141 163.367
R531 B.n151 B.n150 163.367
R532 B.n152 B.n151 163.367
R533 B.n152 B.n139 163.367
R534 B.n156 B.n139 163.367
R535 B.n157 B.n156 163.367
R536 B.n158 B.n157 163.367
R537 B.n158 B.n137 163.367
R538 B.n162 B.n137 163.367
R539 B.n163 B.n162 163.367
R540 B.n164 B.n163 163.367
R541 B.n164 B.n135 163.367
R542 B.n168 B.n135 163.367
R543 B.n169 B.n168 163.367
R544 B.n170 B.n169 163.367
R545 B.n170 B.n133 163.367
R546 B.n106 B.t7 158.525
R547 B.n40 B.t2 158.525
R548 B.n233 B.t4 158.512
R549 B.n34 B.t11 158.512
R550 B.n107 B.t8 113.531
R551 B.n41 B.t1 113.531
R552 B.n234 B.t5 113.517
R553 B.n35 B.t10 113.517
R554 B.n235 B.n234 59.5399
R555 B.n253 B.n107 59.5399
R556 B.n42 B.n41 59.5399
R557 B.n458 B.n35 59.5399
R558 B.n234 B.n233 44.9944
R559 B.n107 B.n106 44.9944
R560 B.n41 B.n40 44.9944
R561 B.n35 B.n34 44.9944
R562 B.n315 B.n314 36.059
R563 B.n519 B.n12 36.059
R564 B.n381 B.n380 36.059
R565 B.n173 B.n172 36.059
R566 B B.n553 18.0485
R567 B.n523 B.n12 10.6151
R568 B.n524 B.n523 10.6151
R569 B.n525 B.n524 10.6151
R570 B.n525 B.n10 10.6151
R571 B.n529 B.n10 10.6151
R572 B.n530 B.n529 10.6151
R573 B.n531 B.n530 10.6151
R574 B.n531 B.n8 10.6151
R575 B.n535 B.n8 10.6151
R576 B.n536 B.n535 10.6151
R577 B.n537 B.n536 10.6151
R578 B.n537 B.n6 10.6151
R579 B.n541 B.n6 10.6151
R580 B.n542 B.n541 10.6151
R581 B.n543 B.n542 10.6151
R582 B.n543 B.n4 10.6151
R583 B.n547 B.n4 10.6151
R584 B.n548 B.n547 10.6151
R585 B.n549 B.n548 10.6151
R586 B.n549 B.n0 10.6151
R587 B.n519 B.n518 10.6151
R588 B.n518 B.n517 10.6151
R589 B.n517 B.n14 10.6151
R590 B.n513 B.n14 10.6151
R591 B.n513 B.n512 10.6151
R592 B.n512 B.n511 10.6151
R593 B.n511 B.n16 10.6151
R594 B.n507 B.n16 10.6151
R595 B.n507 B.n506 10.6151
R596 B.n506 B.n505 10.6151
R597 B.n505 B.n18 10.6151
R598 B.n501 B.n18 10.6151
R599 B.n501 B.n500 10.6151
R600 B.n500 B.n499 10.6151
R601 B.n499 B.n20 10.6151
R602 B.n495 B.n20 10.6151
R603 B.n495 B.n494 10.6151
R604 B.n494 B.n493 10.6151
R605 B.n493 B.n22 10.6151
R606 B.n489 B.n22 10.6151
R607 B.n489 B.n488 10.6151
R608 B.n488 B.n487 10.6151
R609 B.n487 B.n24 10.6151
R610 B.n483 B.n24 10.6151
R611 B.n483 B.n482 10.6151
R612 B.n482 B.n481 10.6151
R613 B.n481 B.n26 10.6151
R614 B.n477 B.n26 10.6151
R615 B.n477 B.n476 10.6151
R616 B.n476 B.n475 10.6151
R617 B.n475 B.n28 10.6151
R618 B.n471 B.n28 10.6151
R619 B.n471 B.n470 10.6151
R620 B.n470 B.n469 10.6151
R621 B.n469 B.n30 10.6151
R622 B.n465 B.n30 10.6151
R623 B.n465 B.n464 10.6151
R624 B.n464 B.n463 10.6151
R625 B.n463 B.n32 10.6151
R626 B.n459 B.n32 10.6151
R627 B.n457 B.n456 10.6151
R628 B.n456 B.n36 10.6151
R629 B.n452 B.n36 10.6151
R630 B.n452 B.n451 10.6151
R631 B.n451 B.n450 10.6151
R632 B.n450 B.n38 10.6151
R633 B.n446 B.n38 10.6151
R634 B.n446 B.n445 10.6151
R635 B.n445 B.n444 10.6151
R636 B.n441 B.n440 10.6151
R637 B.n440 B.n439 10.6151
R638 B.n439 B.n44 10.6151
R639 B.n435 B.n44 10.6151
R640 B.n435 B.n434 10.6151
R641 B.n434 B.n433 10.6151
R642 B.n433 B.n46 10.6151
R643 B.n429 B.n46 10.6151
R644 B.n429 B.n428 10.6151
R645 B.n428 B.n427 10.6151
R646 B.n427 B.n48 10.6151
R647 B.n423 B.n48 10.6151
R648 B.n423 B.n422 10.6151
R649 B.n422 B.n421 10.6151
R650 B.n421 B.n50 10.6151
R651 B.n417 B.n50 10.6151
R652 B.n417 B.n416 10.6151
R653 B.n416 B.n415 10.6151
R654 B.n415 B.n52 10.6151
R655 B.n411 B.n52 10.6151
R656 B.n411 B.n410 10.6151
R657 B.n410 B.n409 10.6151
R658 B.n409 B.n54 10.6151
R659 B.n405 B.n54 10.6151
R660 B.n405 B.n404 10.6151
R661 B.n404 B.n403 10.6151
R662 B.n403 B.n56 10.6151
R663 B.n399 B.n56 10.6151
R664 B.n399 B.n398 10.6151
R665 B.n398 B.n397 10.6151
R666 B.n397 B.n58 10.6151
R667 B.n393 B.n58 10.6151
R668 B.n393 B.n392 10.6151
R669 B.n392 B.n391 10.6151
R670 B.n391 B.n60 10.6151
R671 B.n387 B.n60 10.6151
R672 B.n387 B.n386 10.6151
R673 B.n386 B.n385 10.6151
R674 B.n385 B.n62 10.6151
R675 B.n381 B.n62 10.6151
R676 B.n380 B.n379 10.6151
R677 B.n379 B.n64 10.6151
R678 B.n375 B.n64 10.6151
R679 B.n375 B.n374 10.6151
R680 B.n374 B.n373 10.6151
R681 B.n373 B.n66 10.6151
R682 B.n369 B.n66 10.6151
R683 B.n369 B.n368 10.6151
R684 B.n368 B.n367 10.6151
R685 B.n367 B.n68 10.6151
R686 B.n363 B.n68 10.6151
R687 B.n363 B.n362 10.6151
R688 B.n362 B.n361 10.6151
R689 B.n361 B.n70 10.6151
R690 B.n357 B.n70 10.6151
R691 B.n357 B.n356 10.6151
R692 B.n356 B.n355 10.6151
R693 B.n355 B.n72 10.6151
R694 B.n351 B.n72 10.6151
R695 B.n351 B.n350 10.6151
R696 B.n350 B.n349 10.6151
R697 B.n349 B.n74 10.6151
R698 B.n345 B.n74 10.6151
R699 B.n345 B.n344 10.6151
R700 B.n344 B.n343 10.6151
R701 B.n343 B.n76 10.6151
R702 B.n339 B.n76 10.6151
R703 B.n339 B.n338 10.6151
R704 B.n338 B.n337 10.6151
R705 B.n337 B.n78 10.6151
R706 B.n333 B.n78 10.6151
R707 B.n333 B.n332 10.6151
R708 B.n332 B.n331 10.6151
R709 B.n331 B.n80 10.6151
R710 B.n327 B.n80 10.6151
R711 B.n327 B.n326 10.6151
R712 B.n326 B.n325 10.6151
R713 B.n325 B.n82 10.6151
R714 B.n321 B.n82 10.6151
R715 B.n321 B.n320 10.6151
R716 B.n320 B.n319 10.6151
R717 B.n319 B.n84 10.6151
R718 B.n315 B.n84 10.6151
R719 B.n143 B.n1 10.6151
R720 B.n143 B.n142 10.6151
R721 B.n147 B.n142 10.6151
R722 B.n148 B.n147 10.6151
R723 B.n149 B.n148 10.6151
R724 B.n149 B.n140 10.6151
R725 B.n153 B.n140 10.6151
R726 B.n154 B.n153 10.6151
R727 B.n155 B.n154 10.6151
R728 B.n155 B.n138 10.6151
R729 B.n159 B.n138 10.6151
R730 B.n160 B.n159 10.6151
R731 B.n161 B.n160 10.6151
R732 B.n161 B.n136 10.6151
R733 B.n165 B.n136 10.6151
R734 B.n166 B.n165 10.6151
R735 B.n167 B.n166 10.6151
R736 B.n167 B.n134 10.6151
R737 B.n171 B.n134 10.6151
R738 B.n172 B.n171 10.6151
R739 B.n173 B.n132 10.6151
R740 B.n177 B.n132 10.6151
R741 B.n178 B.n177 10.6151
R742 B.n179 B.n178 10.6151
R743 B.n179 B.n130 10.6151
R744 B.n183 B.n130 10.6151
R745 B.n184 B.n183 10.6151
R746 B.n185 B.n184 10.6151
R747 B.n185 B.n128 10.6151
R748 B.n189 B.n128 10.6151
R749 B.n190 B.n189 10.6151
R750 B.n191 B.n190 10.6151
R751 B.n191 B.n126 10.6151
R752 B.n195 B.n126 10.6151
R753 B.n196 B.n195 10.6151
R754 B.n197 B.n196 10.6151
R755 B.n197 B.n124 10.6151
R756 B.n201 B.n124 10.6151
R757 B.n202 B.n201 10.6151
R758 B.n203 B.n202 10.6151
R759 B.n203 B.n122 10.6151
R760 B.n207 B.n122 10.6151
R761 B.n208 B.n207 10.6151
R762 B.n209 B.n208 10.6151
R763 B.n209 B.n120 10.6151
R764 B.n213 B.n120 10.6151
R765 B.n214 B.n213 10.6151
R766 B.n215 B.n214 10.6151
R767 B.n215 B.n118 10.6151
R768 B.n219 B.n118 10.6151
R769 B.n220 B.n219 10.6151
R770 B.n221 B.n220 10.6151
R771 B.n221 B.n116 10.6151
R772 B.n225 B.n116 10.6151
R773 B.n226 B.n225 10.6151
R774 B.n227 B.n226 10.6151
R775 B.n227 B.n114 10.6151
R776 B.n231 B.n114 10.6151
R777 B.n232 B.n231 10.6151
R778 B.n236 B.n232 10.6151
R779 B.n240 B.n112 10.6151
R780 B.n241 B.n240 10.6151
R781 B.n242 B.n241 10.6151
R782 B.n242 B.n110 10.6151
R783 B.n246 B.n110 10.6151
R784 B.n247 B.n246 10.6151
R785 B.n248 B.n247 10.6151
R786 B.n248 B.n108 10.6151
R787 B.n252 B.n108 10.6151
R788 B.n255 B.n254 10.6151
R789 B.n255 B.n104 10.6151
R790 B.n259 B.n104 10.6151
R791 B.n260 B.n259 10.6151
R792 B.n261 B.n260 10.6151
R793 B.n261 B.n102 10.6151
R794 B.n265 B.n102 10.6151
R795 B.n266 B.n265 10.6151
R796 B.n267 B.n266 10.6151
R797 B.n267 B.n100 10.6151
R798 B.n271 B.n100 10.6151
R799 B.n272 B.n271 10.6151
R800 B.n273 B.n272 10.6151
R801 B.n273 B.n98 10.6151
R802 B.n277 B.n98 10.6151
R803 B.n278 B.n277 10.6151
R804 B.n279 B.n278 10.6151
R805 B.n279 B.n96 10.6151
R806 B.n283 B.n96 10.6151
R807 B.n284 B.n283 10.6151
R808 B.n285 B.n284 10.6151
R809 B.n285 B.n94 10.6151
R810 B.n289 B.n94 10.6151
R811 B.n290 B.n289 10.6151
R812 B.n291 B.n290 10.6151
R813 B.n291 B.n92 10.6151
R814 B.n295 B.n92 10.6151
R815 B.n296 B.n295 10.6151
R816 B.n297 B.n296 10.6151
R817 B.n297 B.n90 10.6151
R818 B.n301 B.n90 10.6151
R819 B.n302 B.n301 10.6151
R820 B.n303 B.n302 10.6151
R821 B.n303 B.n88 10.6151
R822 B.n307 B.n88 10.6151
R823 B.n308 B.n307 10.6151
R824 B.n309 B.n308 10.6151
R825 B.n309 B.n86 10.6151
R826 B.n313 B.n86 10.6151
R827 B.n314 B.n313 10.6151
R828 B.n459 B.n458 9.36635
R829 B.n441 B.n42 9.36635
R830 B.n236 B.n235 9.36635
R831 B.n254 B.n253 9.36635
R832 B.n553 B.n0 8.11757
R833 B.n553 B.n1 8.11757
R834 B.n458 B.n457 1.24928
R835 B.n444 B.n42 1.24928
R836 B.n235 B.n112 1.24928
R837 B.n253 B.n252 1.24928
R838 VN VN.t1 246.002
R839 VN VN.t0 203.096
R840 VTAIL.n1 VTAIL.t2 62.8712
R841 VTAIL.n3 VTAIL.t3 62.8709
R842 VTAIL.n0 VTAIL.t0 62.8709
R843 VTAIL.n2 VTAIL.t1 62.8709
R844 VTAIL.n1 VTAIL.n0 26.6169
R845 VTAIL.n3 VTAIL.n2 24.6169
R846 VTAIL.n2 VTAIL.n1 1.47033
R847 VTAIL VTAIL.n0 1.02852
R848 VTAIL VTAIL.n3 0.44231
R849 VDD2.n0 VDD2.t1 117.46
R850 VDD2.n0 VDD2.t0 79.5497
R851 VDD2 VDD2.n0 0.55869
R852 VP.n0 VP.t1 245.81
R853 VP.n0 VP.t0 202.856
R854 VP VP.n0 0.241678
R855 VDD1 VDD1.t1 118.484
R856 VDD1 VDD1.t0 80.1079
C0 VP VDD2 0.307479f
C1 VN B 0.94555f
C2 w_n1898_n3346# VDD2 1.7239f
C3 VP VN 5.14701f
C4 VN w_n1898_n3346# 2.56289f
C5 VP B 1.33842f
C6 B w_n1898_n3346# 8.11953f
C7 VP w_n1898_n3346# 2.80335f
C8 VDD1 VTAIL 4.9883f
C9 VDD2 VTAIL 5.03406f
C10 VN VTAIL 2.25605f
C11 B VTAIL 3.3724f
C12 VP VTAIL 2.2704f
C13 w_n1898_n3346# VTAIL 2.75964f
C14 VDD2 VDD1 0.60217f
C15 VN VDD1 0.147842f
C16 B VDD1 1.61282f
C17 VP VDD1 2.7895f
C18 w_n1898_n3346# VDD1 1.70532f
C19 VN VDD2 2.63275f
C20 B VDD2 1.6375f
C21 VDD2 VSUBS 0.835153f
C22 VDD1 VSUBS 4.304768f
C23 VTAIL VSUBS 0.928233f
C24 VN VSUBS 7.6739f
C25 VP VSUBS 1.50146f
C26 B VSUBS 3.430091f
C27 w_n1898_n3346# VSUBS 78.189995f
C28 VDD1.t0 VSUBS 1.95897f
C29 VDD1.t1 VSUBS 2.4993f
C30 VP.t1 VSUBS 3.94397f
C31 VP.t0 VSUBS 3.40685f
C32 VP.n0 VSUBS 5.57076f
C33 VDD2.t1 VSUBS 2.42949f
C34 VDD2.t0 VSUBS 1.92401f
C35 VDD2.n0 VSUBS 3.14539f
C36 VTAIL.t0 VSUBS 2.65273f
C37 VTAIL.n0 VSUBS 2.60004f
C38 VTAIL.t2 VSUBS 2.65274f
C39 VTAIL.n1 VSUBS 2.6418f
C40 VTAIL.t1 VSUBS 2.65273f
C41 VTAIL.n2 VSUBS 2.45273f
C42 VTAIL.t3 VSUBS 2.65273f
C43 VTAIL.n3 VSUBS 2.35553f
C44 VN.t0 VSUBS 3.28664f
C45 VN.t1 VSUBS 3.8089f
C46 B.n0 VSUBS 0.005682f
C47 B.n1 VSUBS 0.005682f
C48 B.n2 VSUBS 0.008403f
C49 B.n3 VSUBS 0.006439f
C50 B.n4 VSUBS 0.006439f
C51 B.n5 VSUBS 0.006439f
C52 B.n6 VSUBS 0.006439f
C53 B.n7 VSUBS 0.006439f
C54 B.n8 VSUBS 0.006439f
C55 B.n9 VSUBS 0.006439f
C56 B.n10 VSUBS 0.006439f
C57 B.n11 VSUBS 0.006439f
C58 B.n12 VSUBS 0.015669f
C59 B.n13 VSUBS 0.006439f
C60 B.n14 VSUBS 0.006439f
C61 B.n15 VSUBS 0.006439f
C62 B.n16 VSUBS 0.006439f
C63 B.n17 VSUBS 0.006439f
C64 B.n18 VSUBS 0.006439f
C65 B.n19 VSUBS 0.006439f
C66 B.n20 VSUBS 0.006439f
C67 B.n21 VSUBS 0.006439f
C68 B.n22 VSUBS 0.006439f
C69 B.n23 VSUBS 0.006439f
C70 B.n24 VSUBS 0.006439f
C71 B.n25 VSUBS 0.006439f
C72 B.n26 VSUBS 0.006439f
C73 B.n27 VSUBS 0.006439f
C74 B.n28 VSUBS 0.006439f
C75 B.n29 VSUBS 0.006439f
C76 B.n30 VSUBS 0.006439f
C77 B.n31 VSUBS 0.006439f
C78 B.n32 VSUBS 0.006439f
C79 B.n33 VSUBS 0.006439f
C80 B.t10 VSUBS 0.356074f
C81 B.t11 VSUBS 0.371553f
C82 B.t9 VSUBS 0.973332f
C83 B.n34 VSUBS 0.181382f
C84 B.n35 VSUBS 0.063716f
C85 B.n36 VSUBS 0.006439f
C86 B.n37 VSUBS 0.006439f
C87 B.n38 VSUBS 0.006439f
C88 B.n39 VSUBS 0.006439f
C89 B.t1 VSUBS 0.356068f
C90 B.t2 VSUBS 0.371547f
C91 B.t0 VSUBS 0.973332f
C92 B.n40 VSUBS 0.181388f
C93 B.n41 VSUBS 0.063722f
C94 B.n42 VSUBS 0.014919f
C95 B.n43 VSUBS 0.006439f
C96 B.n44 VSUBS 0.006439f
C97 B.n45 VSUBS 0.006439f
C98 B.n46 VSUBS 0.006439f
C99 B.n47 VSUBS 0.006439f
C100 B.n48 VSUBS 0.006439f
C101 B.n49 VSUBS 0.006439f
C102 B.n50 VSUBS 0.006439f
C103 B.n51 VSUBS 0.006439f
C104 B.n52 VSUBS 0.006439f
C105 B.n53 VSUBS 0.006439f
C106 B.n54 VSUBS 0.006439f
C107 B.n55 VSUBS 0.006439f
C108 B.n56 VSUBS 0.006439f
C109 B.n57 VSUBS 0.006439f
C110 B.n58 VSUBS 0.006439f
C111 B.n59 VSUBS 0.006439f
C112 B.n60 VSUBS 0.006439f
C113 B.n61 VSUBS 0.006439f
C114 B.n62 VSUBS 0.006439f
C115 B.n63 VSUBS 0.015669f
C116 B.n64 VSUBS 0.006439f
C117 B.n65 VSUBS 0.006439f
C118 B.n66 VSUBS 0.006439f
C119 B.n67 VSUBS 0.006439f
C120 B.n68 VSUBS 0.006439f
C121 B.n69 VSUBS 0.006439f
C122 B.n70 VSUBS 0.006439f
C123 B.n71 VSUBS 0.006439f
C124 B.n72 VSUBS 0.006439f
C125 B.n73 VSUBS 0.006439f
C126 B.n74 VSUBS 0.006439f
C127 B.n75 VSUBS 0.006439f
C128 B.n76 VSUBS 0.006439f
C129 B.n77 VSUBS 0.006439f
C130 B.n78 VSUBS 0.006439f
C131 B.n79 VSUBS 0.006439f
C132 B.n80 VSUBS 0.006439f
C133 B.n81 VSUBS 0.006439f
C134 B.n82 VSUBS 0.006439f
C135 B.n83 VSUBS 0.006439f
C136 B.n84 VSUBS 0.006439f
C137 B.n85 VSUBS 0.016526f
C138 B.n86 VSUBS 0.006439f
C139 B.n87 VSUBS 0.006439f
C140 B.n88 VSUBS 0.006439f
C141 B.n89 VSUBS 0.006439f
C142 B.n90 VSUBS 0.006439f
C143 B.n91 VSUBS 0.006439f
C144 B.n92 VSUBS 0.006439f
C145 B.n93 VSUBS 0.006439f
C146 B.n94 VSUBS 0.006439f
C147 B.n95 VSUBS 0.006439f
C148 B.n96 VSUBS 0.006439f
C149 B.n97 VSUBS 0.006439f
C150 B.n98 VSUBS 0.006439f
C151 B.n99 VSUBS 0.006439f
C152 B.n100 VSUBS 0.006439f
C153 B.n101 VSUBS 0.006439f
C154 B.n102 VSUBS 0.006439f
C155 B.n103 VSUBS 0.006439f
C156 B.n104 VSUBS 0.006439f
C157 B.n105 VSUBS 0.006439f
C158 B.t8 VSUBS 0.356068f
C159 B.t7 VSUBS 0.371547f
C160 B.t6 VSUBS 0.973332f
C161 B.n106 VSUBS 0.181388f
C162 B.n107 VSUBS 0.063722f
C163 B.n108 VSUBS 0.006439f
C164 B.n109 VSUBS 0.006439f
C165 B.n110 VSUBS 0.006439f
C166 B.n111 VSUBS 0.006439f
C167 B.n112 VSUBS 0.003598f
C168 B.n113 VSUBS 0.006439f
C169 B.n114 VSUBS 0.006439f
C170 B.n115 VSUBS 0.006439f
C171 B.n116 VSUBS 0.006439f
C172 B.n117 VSUBS 0.006439f
C173 B.n118 VSUBS 0.006439f
C174 B.n119 VSUBS 0.006439f
C175 B.n120 VSUBS 0.006439f
C176 B.n121 VSUBS 0.006439f
C177 B.n122 VSUBS 0.006439f
C178 B.n123 VSUBS 0.006439f
C179 B.n124 VSUBS 0.006439f
C180 B.n125 VSUBS 0.006439f
C181 B.n126 VSUBS 0.006439f
C182 B.n127 VSUBS 0.006439f
C183 B.n128 VSUBS 0.006439f
C184 B.n129 VSUBS 0.006439f
C185 B.n130 VSUBS 0.006439f
C186 B.n131 VSUBS 0.006439f
C187 B.n132 VSUBS 0.006439f
C188 B.n133 VSUBS 0.015669f
C189 B.n134 VSUBS 0.006439f
C190 B.n135 VSUBS 0.006439f
C191 B.n136 VSUBS 0.006439f
C192 B.n137 VSUBS 0.006439f
C193 B.n138 VSUBS 0.006439f
C194 B.n139 VSUBS 0.006439f
C195 B.n140 VSUBS 0.006439f
C196 B.n141 VSUBS 0.006439f
C197 B.n142 VSUBS 0.006439f
C198 B.n143 VSUBS 0.006439f
C199 B.n144 VSUBS 0.006439f
C200 B.n145 VSUBS 0.006439f
C201 B.n146 VSUBS 0.006439f
C202 B.n147 VSUBS 0.006439f
C203 B.n148 VSUBS 0.006439f
C204 B.n149 VSUBS 0.006439f
C205 B.n150 VSUBS 0.006439f
C206 B.n151 VSUBS 0.006439f
C207 B.n152 VSUBS 0.006439f
C208 B.n153 VSUBS 0.006439f
C209 B.n154 VSUBS 0.006439f
C210 B.n155 VSUBS 0.006439f
C211 B.n156 VSUBS 0.006439f
C212 B.n157 VSUBS 0.006439f
C213 B.n158 VSUBS 0.006439f
C214 B.n159 VSUBS 0.006439f
C215 B.n160 VSUBS 0.006439f
C216 B.n161 VSUBS 0.006439f
C217 B.n162 VSUBS 0.006439f
C218 B.n163 VSUBS 0.006439f
C219 B.n164 VSUBS 0.006439f
C220 B.n165 VSUBS 0.006439f
C221 B.n166 VSUBS 0.006439f
C222 B.n167 VSUBS 0.006439f
C223 B.n168 VSUBS 0.006439f
C224 B.n169 VSUBS 0.006439f
C225 B.n170 VSUBS 0.006439f
C226 B.n171 VSUBS 0.006439f
C227 B.n172 VSUBS 0.015669f
C228 B.n173 VSUBS 0.016526f
C229 B.n174 VSUBS 0.016526f
C230 B.n175 VSUBS 0.006439f
C231 B.n176 VSUBS 0.006439f
C232 B.n177 VSUBS 0.006439f
C233 B.n178 VSUBS 0.006439f
C234 B.n179 VSUBS 0.006439f
C235 B.n180 VSUBS 0.006439f
C236 B.n181 VSUBS 0.006439f
C237 B.n182 VSUBS 0.006439f
C238 B.n183 VSUBS 0.006439f
C239 B.n184 VSUBS 0.006439f
C240 B.n185 VSUBS 0.006439f
C241 B.n186 VSUBS 0.006439f
C242 B.n187 VSUBS 0.006439f
C243 B.n188 VSUBS 0.006439f
C244 B.n189 VSUBS 0.006439f
C245 B.n190 VSUBS 0.006439f
C246 B.n191 VSUBS 0.006439f
C247 B.n192 VSUBS 0.006439f
C248 B.n193 VSUBS 0.006439f
C249 B.n194 VSUBS 0.006439f
C250 B.n195 VSUBS 0.006439f
C251 B.n196 VSUBS 0.006439f
C252 B.n197 VSUBS 0.006439f
C253 B.n198 VSUBS 0.006439f
C254 B.n199 VSUBS 0.006439f
C255 B.n200 VSUBS 0.006439f
C256 B.n201 VSUBS 0.006439f
C257 B.n202 VSUBS 0.006439f
C258 B.n203 VSUBS 0.006439f
C259 B.n204 VSUBS 0.006439f
C260 B.n205 VSUBS 0.006439f
C261 B.n206 VSUBS 0.006439f
C262 B.n207 VSUBS 0.006439f
C263 B.n208 VSUBS 0.006439f
C264 B.n209 VSUBS 0.006439f
C265 B.n210 VSUBS 0.006439f
C266 B.n211 VSUBS 0.006439f
C267 B.n212 VSUBS 0.006439f
C268 B.n213 VSUBS 0.006439f
C269 B.n214 VSUBS 0.006439f
C270 B.n215 VSUBS 0.006439f
C271 B.n216 VSUBS 0.006439f
C272 B.n217 VSUBS 0.006439f
C273 B.n218 VSUBS 0.006439f
C274 B.n219 VSUBS 0.006439f
C275 B.n220 VSUBS 0.006439f
C276 B.n221 VSUBS 0.006439f
C277 B.n222 VSUBS 0.006439f
C278 B.n223 VSUBS 0.006439f
C279 B.n224 VSUBS 0.006439f
C280 B.n225 VSUBS 0.006439f
C281 B.n226 VSUBS 0.006439f
C282 B.n227 VSUBS 0.006439f
C283 B.n228 VSUBS 0.006439f
C284 B.n229 VSUBS 0.006439f
C285 B.n230 VSUBS 0.006439f
C286 B.n231 VSUBS 0.006439f
C287 B.n232 VSUBS 0.006439f
C288 B.t5 VSUBS 0.356074f
C289 B.t4 VSUBS 0.371553f
C290 B.t3 VSUBS 0.973332f
C291 B.n233 VSUBS 0.181382f
C292 B.n234 VSUBS 0.063716f
C293 B.n235 VSUBS 0.014919f
C294 B.n236 VSUBS 0.00606f
C295 B.n237 VSUBS 0.006439f
C296 B.n238 VSUBS 0.006439f
C297 B.n239 VSUBS 0.006439f
C298 B.n240 VSUBS 0.006439f
C299 B.n241 VSUBS 0.006439f
C300 B.n242 VSUBS 0.006439f
C301 B.n243 VSUBS 0.006439f
C302 B.n244 VSUBS 0.006439f
C303 B.n245 VSUBS 0.006439f
C304 B.n246 VSUBS 0.006439f
C305 B.n247 VSUBS 0.006439f
C306 B.n248 VSUBS 0.006439f
C307 B.n249 VSUBS 0.006439f
C308 B.n250 VSUBS 0.006439f
C309 B.n251 VSUBS 0.006439f
C310 B.n252 VSUBS 0.003598f
C311 B.n253 VSUBS 0.014919f
C312 B.n254 VSUBS 0.00606f
C313 B.n255 VSUBS 0.006439f
C314 B.n256 VSUBS 0.006439f
C315 B.n257 VSUBS 0.006439f
C316 B.n258 VSUBS 0.006439f
C317 B.n259 VSUBS 0.006439f
C318 B.n260 VSUBS 0.006439f
C319 B.n261 VSUBS 0.006439f
C320 B.n262 VSUBS 0.006439f
C321 B.n263 VSUBS 0.006439f
C322 B.n264 VSUBS 0.006439f
C323 B.n265 VSUBS 0.006439f
C324 B.n266 VSUBS 0.006439f
C325 B.n267 VSUBS 0.006439f
C326 B.n268 VSUBS 0.006439f
C327 B.n269 VSUBS 0.006439f
C328 B.n270 VSUBS 0.006439f
C329 B.n271 VSUBS 0.006439f
C330 B.n272 VSUBS 0.006439f
C331 B.n273 VSUBS 0.006439f
C332 B.n274 VSUBS 0.006439f
C333 B.n275 VSUBS 0.006439f
C334 B.n276 VSUBS 0.006439f
C335 B.n277 VSUBS 0.006439f
C336 B.n278 VSUBS 0.006439f
C337 B.n279 VSUBS 0.006439f
C338 B.n280 VSUBS 0.006439f
C339 B.n281 VSUBS 0.006439f
C340 B.n282 VSUBS 0.006439f
C341 B.n283 VSUBS 0.006439f
C342 B.n284 VSUBS 0.006439f
C343 B.n285 VSUBS 0.006439f
C344 B.n286 VSUBS 0.006439f
C345 B.n287 VSUBS 0.006439f
C346 B.n288 VSUBS 0.006439f
C347 B.n289 VSUBS 0.006439f
C348 B.n290 VSUBS 0.006439f
C349 B.n291 VSUBS 0.006439f
C350 B.n292 VSUBS 0.006439f
C351 B.n293 VSUBS 0.006439f
C352 B.n294 VSUBS 0.006439f
C353 B.n295 VSUBS 0.006439f
C354 B.n296 VSUBS 0.006439f
C355 B.n297 VSUBS 0.006439f
C356 B.n298 VSUBS 0.006439f
C357 B.n299 VSUBS 0.006439f
C358 B.n300 VSUBS 0.006439f
C359 B.n301 VSUBS 0.006439f
C360 B.n302 VSUBS 0.006439f
C361 B.n303 VSUBS 0.006439f
C362 B.n304 VSUBS 0.006439f
C363 B.n305 VSUBS 0.006439f
C364 B.n306 VSUBS 0.006439f
C365 B.n307 VSUBS 0.006439f
C366 B.n308 VSUBS 0.006439f
C367 B.n309 VSUBS 0.006439f
C368 B.n310 VSUBS 0.006439f
C369 B.n311 VSUBS 0.006439f
C370 B.n312 VSUBS 0.006439f
C371 B.n313 VSUBS 0.006439f
C372 B.n314 VSUBS 0.015837f
C373 B.n315 VSUBS 0.016358f
C374 B.n316 VSUBS 0.015669f
C375 B.n317 VSUBS 0.006439f
C376 B.n318 VSUBS 0.006439f
C377 B.n319 VSUBS 0.006439f
C378 B.n320 VSUBS 0.006439f
C379 B.n321 VSUBS 0.006439f
C380 B.n322 VSUBS 0.006439f
C381 B.n323 VSUBS 0.006439f
C382 B.n324 VSUBS 0.006439f
C383 B.n325 VSUBS 0.006439f
C384 B.n326 VSUBS 0.006439f
C385 B.n327 VSUBS 0.006439f
C386 B.n328 VSUBS 0.006439f
C387 B.n329 VSUBS 0.006439f
C388 B.n330 VSUBS 0.006439f
C389 B.n331 VSUBS 0.006439f
C390 B.n332 VSUBS 0.006439f
C391 B.n333 VSUBS 0.006439f
C392 B.n334 VSUBS 0.006439f
C393 B.n335 VSUBS 0.006439f
C394 B.n336 VSUBS 0.006439f
C395 B.n337 VSUBS 0.006439f
C396 B.n338 VSUBS 0.006439f
C397 B.n339 VSUBS 0.006439f
C398 B.n340 VSUBS 0.006439f
C399 B.n341 VSUBS 0.006439f
C400 B.n342 VSUBS 0.006439f
C401 B.n343 VSUBS 0.006439f
C402 B.n344 VSUBS 0.006439f
C403 B.n345 VSUBS 0.006439f
C404 B.n346 VSUBS 0.006439f
C405 B.n347 VSUBS 0.006439f
C406 B.n348 VSUBS 0.006439f
C407 B.n349 VSUBS 0.006439f
C408 B.n350 VSUBS 0.006439f
C409 B.n351 VSUBS 0.006439f
C410 B.n352 VSUBS 0.006439f
C411 B.n353 VSUBS 0.006439f
C412 B.n354 VSUBS 0.006439f
C413 B.n355 VSUBS 0.006439f
C414 B.n356 VSUBS 0.006439f
C415 B.n357 VSUBS 0.006439f
C416 B.n358 VSUBS 0.006439f
C417 B.n359 VSUBS 0.006439f
C418 B.n360 VSUBS 0.006439f
C419 B.n361 VSUBS 0.006439f
C420 B.n362 VSUBS 0.006439f
C421 B.n363 VSUBS 0.006439f
C422 B.n364 VSUBS 0.006439f
C423 B.n365 VSUBS 0.006439f
C424 B.n366 VSUBS 0.006439f
C425 B.n367 VSUBS 0.006439f
C426 B.n368 VSUBS 0.006439f
C427 B.n369 VSUBS 0.006439f
C428 B.n370 VSUBS 0.006439f
C429 B.n371 VSUBS 0.006439f
C430 B.n372 VSUBS 0.006439f
C431 B.n373 VSUBS 0.006439f
C432 B.n374 VSUBS 0.006439f
C433 B.n375 VSUBS 0.006439f
C434 B.n376 VSUBS 0.006439f
C435 B.n377 VSUBS 0.006439f
C436 B.n378 VSUBS 0.006439f
C437 B.n379 VSUBS 0.006439f
C438 B.n380 VSUBS 0.015669f
C439 B.n381 VSUBS 0.016526f
C440 B.n382 VSUBS 0.016526f
C441 B.n383 VSUBS 0.006439f
C442 B.n384 VSUBS 0.006439f
C443 B.n385 VSUBS 0.006439f
C444 B.n386 VSUBS 0.006439f
C445 B.n387 VSUBS 0.006439f
C446 B.n388 VSUBS 0.006439f
C447 B.n389 VSUBS 0.006439f
C448 B.n390 VSUBS 0.006439f
C449 B.n391 VSUBS 0.006439f
C450 B.n392 VSUBS 0.006439f
C451 B.n393 VSUBS 0.006439f
C452 B.n394 VSUBS 0.006439f
C453 B.n395 VSUBS 0.006439f
C454 B.n396 VSUBS 0.006439f
C455 B.n397 VSUBS 0.006439f
C456 B.n398 VSUBS 0.006439f
C457 B.n399 VSUBS 0.006439f
C458 B.n400 VSUBS 0.006439f
C459 B.n401 VSUBS 0.006439f
C460 B.n402 VSUBS 0.006439f
C461 B.n403 VSUBS 0.006439f
C462 B.n404 VSUBS 0.006439f
C463 B.n405 VSUBS 0.006439f
C464 B.n406 VSUBS 0.006439f
C465 B.n407 VSUBS 0.006439f
C466 B.n408 VSUBS 0.006439f
C467 B.n409 VSUBS 0.006439f
C468 B.n410 VSUBS 0.006439f
C469 B.n411 VSUBS 0.006439f
C470 B.n412 VSUBS 0.006439f
C471 B.n413 VSUBS 0.006439f
C472 B.n414 VSUBS 0.006439f
C473 B.n415 VSUBS 0.006439f
C474 B.n416 VSUBS 0.006439f
C475 B.n417 VSUBS 0.006439f
C476 B.n418 VSUBS 0.006439f
C477 B.n419 VSUBS 0.006439f
C478 B.n420 VSUBS 0.006439f
C479 B.n421 VSUBS 0.006439f
C480 B.n422 VSUBS 0.006439f
C481 B.n423 VSUBS 0.006439f
C482 B.n424 VSUBS 0.006439f
C483 B.n425 VSUBS 0.006439f
C484 B.n426 VSUBS 0.006439f
C485 B.n427 VSUBS 0.006439f
C486 B.n428 VSUBS 0.006439f
C487 B.n429 VSUBS 0.006439f
C488 B.n430 VSUBS 0.006439f
C489 B.n431 VSUBS 0.006439f
C490 B.n432 VSUBS 0.006439f
C491 B.n433 VSUBS 0.006439f
C492 B.n434 VSUBS 0.006439f
C493 B.n435 VSUBS 0.006439f
C494 B.n436 VSUBS 0.006439f
C495 B.n437 VSUBS 0.006439f
C496 B.n438 VSUBS 0.006439f
C497 B.n439 VSUBS 0.006439f
C498 B.n440 VSUBS 0.006439f
C499 B.n441 VSUBS 0.00606f
C500 B.n442 VSUBS 0.006439f
C501 B.n443 VSUBS 0.006439f
C502 B.n444 VSUBS 0.003598f
C503 B.n445 VSUBS 0.006439f
C504 B.n446 VSUBS 0.006439f
C505 B.n447 VSUBS 0.006439f
C506 B.n448 VSUBS 0.006439f
C507 B.n449 VSUBS 0.006439f
C508 B.n450 VSUBS 0.006439f
C509 B.n451 VSUBS 0.006439f
C510 B.n452 VSUBS 0.006439f
C511 B.n453 VSUBS 0.006439f
C512 B.n454 VSUBS 0.006439f
C513 B.n455 VSUBS 0.006439f
C514 B.n456 VSUBS 0.006439f
C515 B.n457 VSUBS 0.003598f
C516 B.n458 VSUBS 0.014919f
C517 B.n459 VSUBS 0.00606f
C518 B.n460 VSUBS 0.006439f
C519 B.n461 VSUBS 0.006439f
C520 B.n462 VSUBS 0.006439f
C521 B.n463 VSUBS 0.006439f
C522 B.n464 VSUBS 0.006439f
C523 B.n465 VSUBS 0.006439f
C524 B.n466 VSUBS 0.006439f
C525 B.n467 VSUBS 0.006439f
C526 B.n468 VSUBS 0.006439f
C527 B.n469 VSUBS 0.006439f
C528 B.n470 VSUBS 0.006439f
C529 B.n471 VSUBS 0.006439f
C530 B.n472 VSUBS 0.006439f
C531 B.n473 VSUBS 0.006439f
C532 B.n474 VSUBS 0.006439f
C533 B.n475 VSUBS 0.006439f
C534 B.n476 VSUBS 0.006439f
C535 B.n477 VSUBS 0.006439f
C536 B.n478 VSUBS 0.006439f
C537 B.n479 VSUBS 0.006439f
C538 B.n480 VSUBS 0.006439f
C539 B.n481 VSUBS 0.006439f
C540 B.n482 VSUBS 0.006439f
C541 B.n483 VSUBS 0.006439f
C542 B.n484 VSUBS 0.006439f
C543 B.n485 VSUBS 0.006439f
C544 B.n486 VSUBS 0.006439f
C545 B.n487 VSUBS 0.006439f
C546 B.n488 VSUBS 0.006439f
C547 B.n489 VSUBS 0.006439f
C548 B.n490 VSUBS 0.006439f
C549 B.n491 VSUBS 0.006439f
C550 B.n492 VSUBS 0.006439f
C551 B.n493 VSUBS 0.006439f
C552 B.n494 VSUBS 0.006439f
C553 B.n495 VSUBS 0.006439f
C554 B.n496 VSUBS 0.006439f
C555 B.n497 VSUBS 0.006439f
C556 B.n498 VSUBS 0.006439f
C557 B.n499 VSUBS 0.006439f
C558 B.n500 VSUBS 0.006439f
C559 B.n501 VSUBS 0.006439f
C560 B.n502 VSUBS 0.006439f
C561 B.n503 VSUBS 0.006439f
C562 B.n504 VSUBS 0.006439f
C563 B.n505 VSUBS 0.006439f
C564 B.n506 VSUBS 0.006439f
C565 B.n507 VSUBS 0.006439f
C566 B.n508 VSUBS 0.006439f
C567 B.n509 VSUBS 0.006439f
C568 B.n510 VSUBS 0.006439f
C569 B.n511 VSUBS 0.006439f
C570 B.n512 VSUBS 0.006439f
C571 B.n513 VSUBS 0.006439f
C572 B.n514 VSUBS 0.006439f
C573 B.n515 VSUBS 0.006439f
C574 B.n516 VSUBS 0.006439f
C575 B.n517 VSUBS 0.006439f
C576 B.n518 VSUBS 0.006439f
C577 B.n519 VSUBS 0.016526f
C578 B.n520 VSUBS 0.016526f
C579 B.n521 VSUBS 0.015669f
C580 B.n522 VSUBS 0.006439f
C581 B.n523 VSUBS 0.006439f
C582 B.n524 VSUBS 0.006439f
C583 B.n525 VSUBS 0.006439f
C584 B.n526 VSUBS 0.006439f
C585 B.n527 VSUBS 0.006439f
C586 B.n528 VSUBS 0.006439f
C587 B.n529 VSUBS 0.006439f
C588 B.n530 VSUBS 0.006439f
C589 B.n531 VSUBS 0.006439f
C590 B.n532 VSUBS 0.006439f
C591 B.n533 VSUBS 0.006439f
C592 B.n534 VSUBS 0.006439f
C593 B.n535 VSUBS 0.006439f
C594 B.n536 VSUBS 0.006439f
C595 B.n537 VSUBS 0.006439f
C596 B.n538 VSUBS 0.006439f
C597 B.n539 VSUBS 0.006439f
C598 B.n540 VSUBS 0.006439f
C599 B.n541 VSUBS 0.006439f
C600 B.n542 VSUBS 0.006439f
C601 B.n543 VSUBS 0.006439f
C602 B.n544 VSUBS 0.006439f
C603 B.n545 VSUBS 0.006439f
C604 B.n546 VSUBS 0.006439f
C605 B.n547 VSUBS 0.006439f
C606 B.n548 VSUBS 0.006439f
C607 B.n549 VSUBS 0.006439f
C608 B.n550 VSUBS 0.006439f
C609 B.n551 VSUBS 0.008403f
C610 B.n552 VSUBS 0.008951f
C611 B.n553 VSUBS 0.0178f
.ends

