* NGSPICE file created from tg_sample_0003.ext - technology: sky130A

.subckt tg_sample_0003 VIN VGN VGP VSS VCC VOUT
X0 VOUT.t27 VOUT.t26 VOUT.t27 VCC.t16 sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=0 ps=0 w=6 l=0.15
X1 VOUT.t25 VOUT.t24 VOUT.t25 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0 ps=0 w=3 l=0.15
X2 VOUT.t23 VOUT.t21 VOUT.t22 VSS.t2 sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X3 VCC.t13 VCC.t11 VCC.t12 VCC.t5 sky130_fd_pr__pfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X4 VCC.t10 VCC.t8 VCC.t9 VCC.t1 sky130_fd_pr__pfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X5 VOUT.t20 VOUT.t19 VOUT.t20 VCC.t15 sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=0 ps=0 w=6 l=0.15
X6 VOUT.t18 VOUT.t16 VOUT.t17 VCC.t14 sky130_fd_pr__pfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X7 VOUT.t15 VOUT.t13 VOUT.t14 VSS.t2 sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X8 VSS.t16 VSS.t14 VSS.t15 VSS.t8 sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X9 VOUT.t12 VOUT.t11 VOUT.t12 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0 ps=0 w=3 l=0.15
X10 VSS.t13 VSS.t11 VSS.t12 VSS.t4 sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X11 VSS.t10 VSS.t7 VSS.t9 VSS.t8 sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X12 VCC.t7 VCC.t4 VCC.t6 VCC.t5 sky130_fd_pr__pfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X13 VCC.t3 VCC.t0 VCC.t2 VCC.t1 sky130_fd_pr__pfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X14 VOUT.t10 VOUT.t9 VOUT.t10 VCC.t16 sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=0 ps=0 w=6 l=0.15
X15 VSS.t6 VSS.t3 VSS.t5 VSS.t4 sky130_fd_pr__nfet_01v8 ad=1.425 pd=6.95 as=0 ps=0 w=3 l=0.15
X16 VOUT.t8 VOUT.t7 VOUT.t8 VCC.t15 sky130_fd_pr__pfet_01v8 ad=1.5 pd=6.5 as=0 ps=0 w=6 l=0.15
X17 VOUT.t6 VOUT.t5 VOUT.t6 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0 ps=0 w=3 l=0.15
X18 VOUT.t4 VOUT.t2 VOUT.t3 VCC.t14 sky130_fd_pr__pfet_01v8 ad=2.85 pd=12.95 as=0 ps=0 w=6 l=0.15
X19 VOUT.t1 VOUT.t0 VOUT.t1 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.75 pd=3.5 as=0 ps=0 w=3 l=0.15
R0 VOUT.n17 VOUT.t2 1231.29
R1 VOUT.n19 VOUT.t7 1231.29
R2 VOUT.n8 VOUT.t16 1231.29
R3 VOUT.n10 VOUT.t19 1231.29
R4 VOUT.n18 VOUT.t9 1172.87
R5 VOUT.n9 VOUT.t26 1172.87
R6 VOUT.n14 VOUT.t0 749.292
R7 VOUT.n12 VOUT.t13 749.292
R8 VOUT.n2 VOUT.t24 749.292
R9 VOUT.n0 VOUT.t21 749.292
R10 VOUT.n13 VOUT.t11 690.867
R11 VOUT.n1 VOUT.t5 690.867
R12 VOUT.n15 VOUT.n12 161.489
R13 VOUT.n20 VOUT.n17 161.489
R14 VOUT.n11 VOUT.n8 161.489
R15 VOUT.n3 VOUT.n0 161.489
R16 VOUT.n15 VOUT.n14 161.3
R17 VOUT.n20 VOUT.n19 161.3
R18 VOUT.n11 VOUT.n10 161.3
R19 VOUT.n3 VOUT.n2 161.3
R20 VOUT.n27 VOUT.t20 101.062
R21 VOUT.n29 VOUT.t8 101.062
R22 VOUT.n27 VOUT.n26 92.2941
R23 VOUT.n30 VOUT.n29 92.2941
R24 VOUT.t1 VOUT.n6 90.3335
R25 VOUT.n40 VOUT.t25 90.3335
R26 VOUT.n32 VOUT.t4 83.8236
R27 VOUT.n23 VOUT.t18 83.8236
R28 VOUT.n34 VOUT.n6 79.7731
R29 VOUT.n41 VOUT.n40 79.7731
R30 VOUT.n32 VOUT.n31 76.1756
R31 VOUT.n25 VOUT.n24 75.6153
R32 VOUT.n36 VOUT.t15 73.0943
R33 VOUT.n5 VOUT.t23 73.0943
R34 VOUT.n36 VOUT.n35 63.6547
R35 VOUT.n43 VOUT.n42 63.0943
R36 VOUT.n14 VOUT.n13 36.5157
R37 VOUT.n13 VOUT.n12 36.5157
R38 VOUT.n19 VOUT.n18 36.5157
R39 VOUT.n18 VOUT.n17 36.5157
R40 VOUT.n10 VOUT.n9 36.5157
R41 VOUT.n9 VOUT.n8 36.5157
R42 VOUT.n2 VOUT.n1 36.5157
R43 VOUT.n1 VOUT.n0 36.5157
R44 VOUT.n29 VOUT.n28 14.1815
R45 VOUT.n39 VOUT.n6 12.8884
R46 VOUT.n35 VOUT.t1 10.0005
R47 VOUT.n35 VOUT.t12 10.0005
R48 VOUT.t12 VOUT.n34 10.0005
R49 VOUT.n34 VOUT.t14 10.0005
R50 VOUT.t6 VOUT.n41 10.0005
R51 VOUT.n41 VOUT.t22 10.0005
R52 VOUT.n42 VOUT.t25 10.0005
R53 VOUT.n42 VOUT.t6 10.0005
R54 VOUT.n26 VOUT.t27 8.20883
R55 VOUT.n26 VOUT.t17 8.20883
R56 VOUT.n31 VOUT.t8 8.20883
R57 VOUT.n31 VOUT.t10 8.20883
R58 VOUT.n25 VOUT.t20 8.20883
R59 VOUT.t27 VOUT.n25 8.20883
R60 VOUT.t10 VOUT.n30 8.20883
R61 VOUT.n30 VOUT.t3 8.20883
R62 VOUT.n22 VGP 7.46916
R63 VOUT.n21 VOUT.n16 6.47081
R64 VOUT.n4 VGN 6.3328
R65 VOUT.n24 VOUT.n22 5.12119
R66 VOUT.n23 VOUT.n7 5.06539
R67 VOUT.n38 VOUT.n5 5.06539
R68 VOUT.n16 VOUT.n15 4.9702
R69 VOUT.n21 VOUT.n20 4.9702
R70 VOUT.n33 VOUT.n32 4.88412
R71 VOUT.n37 VOUT.n36 4.88412
R72 VIN VOUT.n4 4.83671
R73 VOUT.n39 VOUT.n38 4.5005
R74 VOUT.n28 VOUT.n7 4.5005
R75 VOUT.n33 VOUT.n7 2.44427
R76 VOUT.n37 VOUT.n33 1.68416
R77 VOUT.n38 VOUT.n37 1.48273
R78 VOUT.n40 VOUT.n39 0.62119
R79 VOUT.n24 VOUT.n23 0.560845
R80 VOUT.n43 VOUT.n5 0.560845
R81 VOUT VOUT.n27 0.401362
R82 VIN VOUT.n43 0.284983
R83 VOUT.n22 VOUT.n21 0.243269
R84 VOUT.n16 VOUT.n4 0.243269
R85 VOUT.n28 VOUT 0.220328
R86 VGP VOUT.n11 0.129288
R87 VGN VOUT.n3 0.129288
R88 VCC.n38 VCC.t0 1220.43
R89 VCC.n40 VCC.t8 1220.43
R90 VCC.n97 VCC.t11 1220.43
R91 VCC.n95 VCC.t4 1220.43
R92 VCC.n336 VCC.n10 339.512
R93 VCC.n240 VCC.n239 339.512
R94 VCC.n100 VCC.n63 339.512
R95 VCC.n196 VCC.n64 339.512
R96 VCC.n239 VCC.n238 185
R97 VCC.n239 VCC.n13 185
R98 VCC.n237 VCC.n44 185
R99 VCC.n228 VCC.n44 185
R100 VCC.n49 VCC.n45 185
R101 VCC.n229 VCC.n49 185
R102 VCC.n233 VCC.n232 185
R103 VCC.n232 VCC.n231 185
R104 VCC.n48 VCC.n47 185
R105 VCC.n227 VCC.n48 185
R106 VCC.n225 VCC.n224 185
R107 VCC.n226 VCC.n225 185
R108 VCC.n52 VCC.n51 185
R109 VCC.n51 VCC.n50 185
R110 VCC.n220 VCC.n219 185
R111 VCC.n219 VCC.n218 185
R112 VCC.n55 VCC.n54 185
R113 VCC.n215 VCC.n55 185
R114 VCC.n213 VCC.n212 185
R115 VCC.n214 VCC.n213 185
R116 VCC.n60 VCC.n59 185
R117 VCC.n59 VCC.n58 185
R118 VCC.n208 VCC.n207 185
R119 VCC.n207 VCC.n206 185
R120 VCC.n63 VCC.n62 185
R121 VCC.n93 VCC.n63 185
R122 VCC.n66 VCC.n64 185
R123 VCC.n93 VCC.n64 185
R124 VCC.n205 VCC.n204 185
R125 VCC.n206 VCC.n205 185
R126 VCC.n67 VCC.n65 185
R127 VCC.n65 VCC.n58 185
R128 VCC.n200 VCC.n56 185
R129 VCC.n214 VCC.n56 185
R130 VCC.n216 VCC.n57 185
R131 VCC.n216 VCC.n215 185
R132 VCC.n217 VCC.n2 185
R133 VCC.n218 VCC.n217 185
R134 VCC.n347 VCC.n3 185
R135 VCC.n50 VCC.n3 185
R136 VCC.n346 VCC.n4 185
R137 VCC.n226 VCC.n4 185
R138 VCC.n345 VCC.n5 185
R139 VCC.n227 VCC.n5 185
R140 VCC.n230 VCC.n6 185
R141 VCC.n231 VCC.n230 185
R142 VCC.n341 VCC.n8 185
R143 VCC.n229 VCC.n8 185
R144 VCC.n340 VCC.n9 185
R145 VCC.n228 VCC.n9 185
R146 VCC.n339 VCC.n10 185
R147 VCC.n13 VCC.n10 185
R148 VCC.n241 VCC.n240 185
R149 VCC.n243 VCC.n242 185
R150 VCC.n245 VCC.n244 185
R151 VCC.n247 VCC.n246 185
R152 VCC.n249 VCC.n248 185
R153 VCC.n251 VCC.n250 185
R154 VCC.n253 VCC.n252 185
R155 VCC.n255 VCC.n254 185
R156 VCC.n257 VCC.n256 185
R157 VCC.n259 VCC.n258 185
R158 VCC.n261 VCC.n260 185
R159 VCC.n263 VCC.n262 185
R160 VCC.n265 VCC.n264 185
R161 VCC.n267 VCC.n266 185
R162 VCC.n269 VCC.n268 185
R163 VCC.n271 VCC.n270 185
R164 VCC.n273 VCC.n272 185
R165 VCC.n275 VCC.n274 185
R166 VCC.n277 VCC.n276 185
R167 VCC.n279 VCC.n278 185
R168 VCC.n281 VCC.n280 185
R169 VCC.n283 VCC.n282 185
R170 VCC.n285 VCC.n284 185
R171 VCC.n287 VCC.n286 185
R172 VCC.n289 VCC.n288 185
R173 VCC.n291 VCC.n290 185
R174 VCC.n293 VCC.n292 185
R175 VCC.n295 VCC.n294 185
R176 VCC.n297 VCC.n296 185
R177 VCC.n299 VCC.n298 185
R178 VCC.n301 VCC.n300 185
R179 VCC.n303 VCC.n302 185
R180 VCC.n305 VCC.n304 185
R181 VCC.n307 VCC.n306 185
R182 VCC.n309 VCC.n308 185
R183 VCC.n311 VCC.n310 185
R184 VCC.n313 VCC.n312 185
R185 VCC.n315 VCC.n314 185
R186 VCC.n317 VCC.n316 185
R187 VCC.n319 VCC.n318 185
R188 VCC.n321 VCC.n320 185
R189 VCC.n323 VCC.n322 185
R190 VCC.n325 VCC.n324 185
R191 VCC.n327 VCC.n326 185
R192 VCC.n329 VCC.n328 185
R193 VCC.n330 VCC.n37 185
R194 VCC.n333 VCC.n332 185
R195 VCC.n12 VCC.n11 185
R196 VCC.n337 VCC.n336 185
R197 VCC.n336 VCC.n335 185
R198 VCC.n197 VCC.n196 185
R199 VCC.n69 VCC.n68 185
R200 VCC.n193 VCC.n192 185
R201 VCC.n194 VCC.n193 185
R202 VCC.n190 VCC.n94 185
R203 VCC.n189 VCC.n188 185
R204 VCC.n187 VCC.n186 185
R205 VCC.n185 VCC.n184 185
R206 VCC.n183 VCC.n182 185
R207 VCC.n181 VCC.n180 185
R208 VCC.n179 VCC.n178 185
R209 VCC.n177 VCC.n176 185
R210 VCC.n175 VCC.n174 185
R211 VCC.n173 VCC.n172 185
R212 VCC.n171 VCC.n170 185
R213 VCC.n169 VCC.n168 185
R214 VCC.n167 VCC.n166 185
R215 VCC.n165 VCC.n164 185
R216 VCC.n163 VCC.n162 185
R217 VCC.n161 VCC.n160 185
R218 VCC.n159 VCC.n158 185
R219 VCC.n157 VCC.n156 185
R220 VCC.n155 VCC.n154 185
R221 VCC.n153 VCC.n152 185
R222 VCC.n151 VCC.n150 185
R223 VCC.n149 VCC.n148 185
R224 VCC.n147 VCC.n146 185
R225 VCC.n145 VCC.n144 185
R226 VCC.n143 VCC.n142 185
R227 VCC.n141 VCC.n140 185
R228 VCC.n139 VCC.n138 185
R229 VCC.n137 VCC.n136 185
R230 VCC.n135 VCC.n134 185
R231 VCC.n133 VCC.n132 185
R232 VCC.n131 VCC.n130 185
R233 VCC.n129 VCC.n128 185
R234 VCC.n127 VCC.n126 185
R235 VCC.n125 VCC.n124 185
R236 VCC.n123 VCC.n122 185
R237 VCC.n121 VCC.n120 185
R238 VCC.n119 VCC.n118 185
R239 VCC.n117 VCC.n116 185
R240 VCC.n115 VCC.n114 185
R241 VCC.n113 VCC.n112 185
R242 VCC.n111 VCC.n110 185
R243 VCC.n109 VCC.n108 185
R244 VCC.n107 VCC.n106 185
R245 VCC.n105 VCC.n104 185
R246 VCC.n103 VCC.n102 185
R247 VCC.n101 VCC.n100 185
R248 VCC.n207 VCC.n63 146.341
R249 VCC.n207 VCC.n59 146.341
R250 VCC.n213 VCC.n59 146.341
R251 VCC.n213 VCC.n55 146.341
R252 VCC.n219 VCC.n55 146.341
R253 VCC.n219 VCC.n51 146.341
R254 VCC.n225 VCC.n51 146.341
R255 VCC.n225 VCC.n48 146.341
R256 VCC.n232 VCC.n48 146.341
R257 VCC.n232 VCC.n49 146.341
R258 VCC.n49 VCC.n44 146.341
R259 VCC.n239 VCC.n44 146.341
R260 VCC.n205 VCC.n64 146.341
R261 VCC.n205 VCC.n65 146.341
R262 VCC.n65 VCC.n56 146.341
R263 VCC.n216 VCC.n56 146.341
R264 VCC.n217 VCC.n216 146.341
R265 VCC.n217 VCC.n3 146.341
R266 VCC.n4 VCC.n3 146.341
R267 VCC.n5 VCC.n4 146.341
R268 VCC.n230 VCC.n5 146.341
R269 VCC.n230 VCC.n8 146.341
R270 VCC.n9 VCC.n8 146.341
R271 VCC.n10 VCC.n9 146.341
R272 VCC.n38 VCC.t2 130.923
R273 VCC.n40 VCC.t9 130.923
R274 VCC.n97 VCC.t13 130.923
R275 VCC.n95 VCC.t7 130.923
R276 VCC.n39 VCC.t3 118.317
R277 VCC.n41 VCC.t10 118.317
R278 VCC.n98 VCC.t12 118.317
R279 VCC.n96 VCC.t6 118.317
R280 VCC.n336 VCC.n12 99.5127
R281 VCC.n333 VCC.n37 99.5127
R282 VCC.n328 VCC.n327 99.5127
R283 VCC.n324 VCC.n323 99.5127
R284 VCC.n320 VCC.n319 99.5127
R285 VCC.n316 VCC.n315 99.5127
R286 VCC.n312 VCC.n311 99.5127
R287 VCC.n308 VCC.n307 99.5127
R288 VCC.n304 VCC.n303 99.5127
R289 VCC.n300 VCC.n299 99.5127
R290 VCC.n296 VCC.n295 99.5127
R291 VCC.n292 VCC.n291 99.5127
R292 VCC.n288 VCC.n287 99.5127
R293 VCC.n284 VCC.n283 99.5127
R294 VCC.n280 VCC.n279 99.5127
R295 VCC.n276 VCC.n275 99.5127
R296 VCC.n272 VCC.n271 99.5127
R297 VCC.n268 VCC.n267 99.5127
R298 VCC.n264 VCC.n263 99.5127
R299 VCC.n260 VCC.n259 99.5127
R300 VCC.n256 VCC.n255 99.5127
R301 VCC.n252 VCC.n251 99.5127
R302 VCC.n248 VCC.n247 99.5127
R303 VCC.n244 VCC.n243 99.5127
R304 VCC.n193 VCC.n69 99.5127
R305 VCC.n193 VCC.n94 99.5127
R306 VCC.n188 VCC.n187 99.5127
R307 VCC.n184 VCC.n183 99.5127
R308 VCC.n180 VCC.n179 99.5127
R309 VCC.n176 VCC.n175 99.5127
R310 VCC.n172 VCC.n171 99.5127
R311 VCC.n168 VCC.n167 99.5127
R312 VCC.n164 VCC.n163 99.5127
R313 VCC.n160 VCC.n159 99.5127
R314 VCC.n156 VCC.n155 99.5127
R315 VCC.n152 VCC.n151 99.5127
R316 VCC.n148 VCC.n147 99.5127
R317 VCC.n144 VCC.n143 99.5127
R318 VCC.n140 VCC.n139 99.5127
R319 VCC.n136 VCC.n135 99.5127
R320 VCC.n132 VCC.n131 99.5127
R321 VCC.n128 VCC.n127 99.5127
R322 VCC.n124 VCC.n123 99.5127
R323 VCC.n120 VCC.n119 99.5127
R324 VCC.n116 VCC.n115 99.5127
R325 VCC.n112 VCC.n111 99.5127
R326 VCC.n108 VCC.n107 99.5127
R327 VCC.n104 VCC.n103 99.5127
R328 VCC.n335 VCC.n14 72.8958
R329 VCC.n335 VCC.n15 72.8958
R330 VCC.n335 VCC.n16 72.8958
R331 VCC.n335 VCC.n17 72.8958
R332 VCC.n335 VCC.n18 72.8958
R333 VCC.n335 VCC.n19 72.8958
R334 VCC.n335 VCC.n20 72.8958
R335 VCC.n335 VCC.n21 72.8958
R336 VCC.n335 VCC.n22 72.8958
R337 VCC.n335 VCC.n23 72.8958
R338 VCC.n335 VCC.n24 72.8958
R339 VCC.n335 VCC.n25 72.8958
R340 VCC.n335 VCC.n26 72.8958
R341 VCC.n335 VCC.n27 72.8958
R342 VCC.n335 VCC.n28 72.8958
R343 VCC.n335 VCC.n29 72.8958
R344 VCC.n335 VCC.n30 72.8958
R345 VCC.n335 VCC.n31 72.8958
R346 VCC.n335 VCC.n32 72.8958
R347 VCC.n335 VCC.n33 72.8958
R348 VCC.n335 VCC.n34 72.8958
R349 VCC.n335 VCC.n35 72.8958
R350 VCC.n335 VCC.n36 72.8958
R351 VCC.n335 VCC.n334 72.8958
R352 VCC.n195 VCC.n194 72.8958
R353 VCC.n194 VCC.n70 72.8958
R354 VCC.n194 VCC.n71 72.8958
R355 VCC.n194 VCC.n72 72.8958
R356 VCC.n194 VCC.n73 72.8958
R357 VCC.n194 VCC.n74 72.8958
R358 VCC.n194 VCC.n75 72.8958
R359 VCC.n194 VCC.n76 72.8958
R360 VCC.n194 VCC.n77 72.8958
R361 VCC.n194 VCC.n78 72.8958
R362 VCC.n194 VCC.n79 72.8958
R363 VCC.n194 VCC.n80 72.8958
R364 VCC.n194 VCC.n81 72.8958
R365 VCC.n194 VCC.n82 72.8958
R366 VCC.n194 VCC.n83 72.8958
R367 VCC.n194 VCC.n84 72.8958
R368 VCC.n194 VCC.n85 72.8958
R369 VCC.n194 VCC.n86 72.8958
R370 VCC.n194 VCC.n87 72.8958
R371 VCC.n194 VCC.n88 72.8958
R372 VCC.n194 VCC.n89 72.8958
R373 VCC.n194 VCC.n90 72.8958
R374 VCC.n194 VCC.n91 72.8958
R375 VCC.n194 VCC.n92 72.8958
R376 VCC.n194 VCC.n93 41.9653
R377 VCC.n335 VCC.n13 41.9653
R378 VCC.n331 VCC.n39 40.146
R379 VCC.n42 VCC.n41 40.146
R380 VCC.n334 VCC.n333 39.2114
R381 VCC.n328 VCC.n36 39.2114
R382 VCC.n324 VCC.n35 39.2114
R383 VCC.n320 VCC.n34 39.2114
R384 VCC.n316 VCC.n33 39.2114
R385 VCC.n312 VCC.n32 39.2114
R386 VCC.n308 VCC.n31 39.2114
R387 VCC.n304 VCC.n30 39.2114
R388 VCC.n300 VCC.n29 39.2114
R389 VCC.n296 VCC.n28 39.2114
R390 VCC.n292 VCC.n27 39.2114
R391 VCC.n288 VCC.n26 39.2114
R392 VCC.n284 VCC.n25 39.2114
R393 VCC.n280 VCC.n24 39.2114
R394 VCC.n276 VCC.n23 39.2114
R395 VCC.n272 VCC.n22 39.2114
R396 VCC.n268 VCC.n21 39.2114
R397 VCC.n264 VCC.n20 39.2114
R398 VCC.n260 VCC.n19 39.2114
R399 VCC.n256 VCC.n18 39.2114
R400 VCC.n252 VCC.n17 39.2114
R401 VCC.n248 VCC.n16 39.2114
R402 VCC.n244 VCC.n15 39.2114
R403 VCC.n240 VCC.n14 39.2114
R404 VCC.n196 VCC.n195 39.2114
R405 VCC.n94 VCC.n70 39.2114
R406 VCC.n187 VCC.n71 39.2114
R407 VCC.n183 VCC.n72 39.2114
R408 VCC.n179 VCC.n73 39.2114
R409 VCC.n175 VCC.n74 39.2114
R410 VCC.n171 VCC.n75 39.2114
R411 VCC.n167 VCC.n76 39.2114
R412 VCC.n163 VCC.n77 39.2114
R413 VCC.n159 VCC.n78 39.2114
R414 VCC.n155 VCC.n79 39.2114
R415 VCC.n151 VCC.n80 39.2114
R416 VCC.n147 VCC.n81 39.2114
R417 VCC.n143 VCC.n82 39.2114
R418 VCC.n139 VCC.n83 39.2114
R419 VCC.n135 VCC.n84 39.2114
R420 VCC.n131 VCC.n85 39.2114
R421 VCC.n127 VCC.n86 39.2114
R422 VCC.n123 VCC.n87 39.2114
R423 VCC.n119 VCC.n88 39.2114
R424 VCC.n115 VCC.n89 39.2114
R425 VCC.n111 VCC.n90 39.2114
R426 VCC.n107 VCC.n91 39.2114
R427 VCC.n103 VCC.n92 39.2114
R428 VCC.n243 VCC.n14 39.2114
R429 VCC.n247 VCC.n15 39.2114
R430 VCC.n251 VCC.n16 39.2114
R431 VCC.n255 VCC.n17 39.2114
R432 VCC.n259 VCC.n18 39.2114
R433 VCC.n263 VCC.n19 39.2114
R434 VCC.n267 VCC.n20 39.2114
R435 VCC.n271 VCC.n21 39.2114
R436 VCC.n275 VCC.n22 39.2114
R437 VCC.n279 VCC.n23 39.2114
R438 VCC.n283 VCC.n24 39.2114
R439 VCC.n287 VCC.n25 39.2114
R440 VCC.n291 VCC.n26 39.2114
R441 VCC.n295 VCC.n27 39.2114
R442 VCC.n299 VCC.n28 39.2114
R443 VCC.n303 VCC.n29 39.2114
R444 VCC.n307 VCC.n30 39.2114
R445 VCC.n311 VCC.n31 39.2114
R446 VCC.n315 VCC.n32 39.2114
R447 VCC.n319 VCC.n33 39.2114
R448 VCC.n323 VCC.n34 39.2114
R449 VCC.n327 VCC.n35 39.2114
R450 VCC.n37 VCC.n36 39.2114
R451 VCC.n334 VCC.n12 39.2114
R452 VCC.n195 VCC.n69 39.2114
R453 VCC.n188 VCC.n70 39.2114
R454 VCC.n184 VCC.n71 39.2114
R455 VCC.n180 VCC.n72 39.2114
R456 VCC.n176 VCC.n73 39.2114
R457 VCC.n172 VCC.n74 39.2114
R458 VCC.n168 VCC.n75 39.2114
R459 VCC.n164 VCC.n76 39.2114
R460 VCC.n160 VCC.n77 39.2114
R461 VCC.n156 VCC.n78 39.2114
R462 VCC.n152 VCC.n79 39.2114
R463 VCC.n148 VCC.n80 39.2114
R464 VCC.n144 VCC.n81 39.2114
R465 VCC.n140 VCC.n82 39.2114
R466 VCC.n136 VCC.n83 39.2114
R467 VCC.n132 VCC.n84 39.2114
R468 VCC.n128 VCC.n85 39.2114
R469 VCC.n124 VCC.n86 39.2114
R470 VCC.n120 VCC.n87 39.2114
R471 VCC.n116 VCC.n88 39.2114
R472 VCC.n112 VCC.n89 39.2114
R473 VCC.n108 VCC.n90 39.2114
R474 VCC.n104 VCC.n91 39.2114
R475 VCC.n100 VCC.n92 39.2114
R476 VCC.n99 VCC.n98 29.2853
R477 VCC.n191 VCC.n96 29.2853
R478 VCC.n338 VCC.n337 26.7197
R479 VCC.n241 VCC.n43 26.7197
R480 VCC.n198 VCC.n197 26.7197
R481 VCC.n101 VCC.n61 26.7197
R482 VCC.n206 VCC.n58 25.7458
R483 VCC.n214 VCC.n58 25.7458
R484 VCC.n215 VCC.n214 25.7458
R485 VCC.n226 VCC.n50 25.7458
R486 VCC.n231 VCC.n227 25.7458
R487 VCC.n231 VCC.n229 25.7458
R488 VCC.n228 VCC.n13 25.7458
R489 VCC.n227 VCC.t14 25.2309
R490 VCC.n93 VCC.t5 24.201
R491 VCC.n208 VCC.n62 19.3944
R492 VCC.n208 VCC.n60 19.3944
R493 VCC.n212 VCC.n60 19.3944
R494 VCC.n212 VCC.n54 19.3944
R495 VCC.n220 VCC.n54 19.3944
R496 VCC.n220 VCC.n52 19.3944
R497 VCC.n224 VCC.n52 19.3944
R498 VCC.n224 VCC.n47 19.3944
R499 VCC.n233 VCC.n47 19.3944
R500 VCC.n233 VCC.n45 19.3944
R501 VCC.n237 VCC.n45 19.3944
R502 VCC.n238 VCC.n237 19.3944
R503 VCC.n204 VCC.n66 19.3944
R504 VCC.n204 VCC.n67 19.3944
R505 VCC.n200 VCC.n67 19.3944
R506 VCC.n200 VCC.n57 19.3944
R507 VCC.n57 VCC.n2 19.3944
R508 VCC.n347 VCC.n2 19.3944
R509 VCC.n347 VCC.n346 19.3944
R510 VCC.n346 VCC.n345 19.3944
R511 VCC.n345 VCC.n6 19.3944
R512 VCC.n341 VCC.n6 19.3944
R513 VCC.n341 VCC.n340 19.3944
R514 VCC.n340 VCC.n339 19.3944
R515 VCC.n218 VCC.t16 18.5371
R516 VCC.n218 VCC.t15 14.9327
R517 VCC.n229 VCC.t1 12.8731
R518 VCC.t1 VCC.n228 12.8731
R519 VCC.n39 VCC.n38 12.6066
R520 VCC.n41 VCC.n40 12.6066
R521 VCC.n98 VCC.n97 12.6066
R522 VCC.n96 VCC.n95 12.6066
R523 VCC.n215 VCC.t15 10.8135
R524 VCC.n337 VCC.n11 10.6151
R525 VCC.n332 VCC.n11 10.6151
R526 VCC.n330 VCC.n329 10.6151
R527 VCC.n329 VCC.n326 10.6151
R528 VCC.n326 VCC.n325 10.6151
R529 VCC.n325 VCC.n322 10.6151
R530 VCC.n322 VCC.n321 10.6151
R531 VCC.n321 VCC.n318 10.6151
R532 VCC.n318 VCC.n317 10.6151
R533 VCC.n317 VCC.n314 10.6151
R534 VCC.n314 VCC.n313 10.6151
R535 VCC.n313 VCC.n310 10.6151
R536 VCC.n310 VCC.n309 10.6151
R537 VCC.n309 VCC.n306 10.6151
R538 VCC.n306 VCC.n305 10.6151
R539 VCC.n305 VCC.n302 10.6151
R540 VCC.n302 VCC.n301 10.6151
R541 VCC.n301 VCC.n298 10.6151
R542 VCC.n298 VCC.n297 10.6151
R543 VCC.n297 VCC.n294 10.6151
R544 VCC.n294 VCC.n293 10.6151
R545 VCC.n293 VCC.n290 10.6151
R546 VCC.n290 VCC.n289 10.6151
R547 VCC.n289 VCC.n286 10.6151
R548 VCC.n286 VCC.n285 10.6151
R549 VCC.n282 VCC.n281 10.6151
R550 VCC.n281 VCC.n278 10.6151
R551 VCC.n278 VCC.n277 10.6151
R552 VCC.n277 VCC.n274 10.6151
R553 VCC.n274 VCC.n273 10.6151
R554 VCC.n273 VCC.n270 10.6151
R555 VCC.n270 VCC.n269 10.6151
R556 VCC.n269 VCC.n266 10.6151
R557 VCC.n266 VCC.n265 10.6151
R558 VCC.n265 VCC.n262 10.6151
R559 VCC.n262 VCC.n261 10.6151
R560 VCC.n261 VCC.n258 10.6151
R561 VCC.n258 VCC.n257 10.6151
R562 VCC.n257 VCC.n254 10.6151
R563 VCC.n254 VCC.n253 10.6151
R564 VCC.n253 VCC.n250 10.6151
R565 VCC.n250 VCC.n249 10.6151
R566 VCC.n249 VCC.n246 10.6151
R567 VCC.n246 VCC.n245 10.6151
R568 VCC.n245 VCC.n242 10.6151
R569 VCC.n242 VCC.n241 10.6151
R570 VCC.n197 VCC.n68 10.6151
R571 VCC.n192 VCC.n68 10.6151
R572 VCC.n190 VCC.n189 10.6151
R573 VCC.n189 VCC.n186 10.6151
R574 VCC.n186 VCC.n185 10.6151
R575 VCC.n185 VCC.n182 10.6151
R576 VCC.n182 VCC.n181 10.6151
R577 VCC.n181 VCC.n178 10.6151
R578 VCC.n178 VCC.n177 10.6151
R579 VCC.n177 VCC.n174 10.6151
R580 VCC.n174 VCC.n173 10.6151
R581 VCC.n173 VCC.n170 10.6151
R582 VCC.n170 VCC.n169 10.6151
R583 VCC.n169 VCC.n166 10.6151
R584 VCC.n166 VCC.n165 10.6151
R585 VCC.n165 VCC.n162 10.6151
R586 VCC.n162 VCC.n161 10.6151
R587 VCC.n161 VCC.n158 10.6151
R588 VCC.n158 VCC.n157 10.6151
R589 VCC.n157 VCC.n154 10.6151
R590 VCC.n154 VCC.n153 10.6151
R591 VCC.n153 VCC.n150 10.6151
R592 VCC.n150 VCC.n149 10.6151
R593 VCC.n149 VCC.n146 10.6151
R594 VCC.n146 VCC.n145 10.6151
R595 VCC.n142 VCC.n141 10.6151
R596 VCC.n141 VCC.n138 10.6151
R597 VCC.n138 VCC.n137 10.6151
R598 VCC.n137 VCC.n134 10.6151
R599 VCC.n134 VCC.n133 10.6151
R600 VCC.n133 VCC.n130 10.6151
R601 VCC.n130 VCC.n129 10.6151
R602 VCC.n129 VCC.n126 10.6151
R603 VCC.n126 VCC.n125 10.6151
R604 VCC.n125 VCC.n122 10.6151
R605 VCC.n122 VCC.n121 10.6151
R606 VCC.n121 VCC.n118 10.6151
R607 VCC.n118 VCC.n117 10.6151
R608 VCC.n117 VCC.n114 10.6151
R609 VCC.n114 VCC.n113 10.6151
R610 VCC.n113 VCC.n110 10.6151
R611 VCC.n110 VCC.n109 10.6151
R612 VCC.n109 VCC.n106 10.6151
R613 VCC.n106 VCC.n105 10.6151
R614 VCC.n105 VCC.n102 10.6151
R615 VCC.n102 VCC.n101 10.6151
R616 VCC.n346 VCC.n0 9.3005
R617 VCC.n345 VCC.n344 9.3005
R618 VCC.n343 VCC.n6 9.3005
R619 VCC.n342 VCC.n341 9.3005
R620 VCC.n340 VCC.n7 9.3005
R621 VCC.n339 VCC.n338 9.3005
R622 VCC.n209 VCC.n208 9.3005
R623 VCC.n210 VCC.n60 9.3005
R624 VCC.n212 VCC.n211 9.3005
R625 VCC.n54 VCC.n53 9.3005
R626 VCC.n221 VCC.n220 9.3005
R627 VCC.n222 VCC.n52 9.3005
R628 VCC.n224 VCC.n223 9.3005
R629 VCC.n47 VCC.n46 9.3005
R630 VCC.n234 VCC.n233 9.3005
R631 VCC.n235 VCC.n45 9.3005
R632 VCC.n237 VCC.n236 9.3005
R633 VCC.n238 VCC.n43 9.3005
R634 VCC.n62 VCC.n61 9.3005
R635 VCC.n198 VCC.n66 9.3005
R636 VCC.n204 VCC.n203 9.3005
R637 VCC.n202 VCC.n67 9.3005
R638 VCC.n201 VCC.n200 9.3005
R639 VCC.n199 VCC.n57 9.3005
R640 VCC.n2 VCC.n1 9.3005
R641 VCC.n348 VCC.n347 9.3005
R642 VCC.n331 VCC.n330 9.21026
R643 VCC.n191 VCC.n190 9.21026
R644 VCC.t16 VCC.n50 7.20917
R645 VCC.n282 VCC.n42 6.0883
R646 VCC.n142 VCC.n99 6.0883
R647 VCC.n285 VCC.n42 4.52733
R648 VCC.n145 VCC.n99 4.52733
R649 VCC.n206 VCC.t5 1.54522
R650 VCC.n332 VCC.n331 1.40538
R651 VCC.n192 VCC.n191 1.40538
R652 VCC.t14 VCC.n226 0.515405
R653 VCC.n344 VCC.n0 0.152939
R654 VCC.n344 VCC.n343 0.152939
R655 VCC.n343 VCC.n342 0.152939
R656 VCC.n342 VCC.n7 0.152939
R657 VCC.n338 VCC.n7 0.152939
R658 VCC.n209 VCC.n61 0.152939
R659 VCC.n210 VCC.n209 0.152939
R660 VCC.n211 VCC.n210 0.152939
R661 VCC.n211 VCC.n53 0.152939
R662 VCC.n221 VCC.n53 0.152939
R663 VCC.n222 VCC.n221 0.152939
R664 VCC.n223 VCC.n222 0.152939
R665 VCC.n223 VCC.n46 0.152939
R666 VCC.n234 VCC.n46 0.152939
R667 VCC.n235 VCC.n234 0.152939
R668 VCC.n236 VCC.n235 0.152939
R669 VCC.n236 VCC.n43 0.152939
R670 VCC.n203 VCC.n198 0.152939
R671 VCC.n203 VCC.n202 0.152939
R672 VCC.n202 VCC.n201 0.152939
R673 VCC.n201 VCC.n199 0.152939
R674 VCC.n199 VCC.n1 0.152939
R675 VCC.n348 VCC.n1 0.13922
R676 VCC VCC.n0 0.0767195
R677 VCC VCC.n348 0.063
R678 VSS.n31 VSS.t3 738.433
R679 VSS.n29 VSS.t11 738.433
R680 VSS.n80 VSS.t14 738.433
R681 VSS.n78 VSS.t7 738.433
R682 VSS.n141 VSS.n54 631.841
R683 VSS.n144 VSS.n55 631.841
R684 VSS.n188 VSS.n187 631.841
R685 VSS.n251 VSS.n10 631.841
R686 VSS.n54 VSS.n53 585
R687 VSS.n75 VSS.n54 585
R688 VSS.n156 VSS.n155 585
R689 VSS.n155 VSS.n154 585
R690 VSS.n51 VSS.n50 585
R691 VSS.n50 VSS.n49 585
R692 VSS.n161 VSS.n160 585
R693 VSS.n162 VSS.n161 585
R694 VSS.n46 VSS.n45 585
R695 VSS.n163 VSS.n46 585
R696 VSS.n168 VSS.n167 585
R697 VSS.n167 VSS.n166 585
R698 VSS.n43 VSS.n42 585
R699 VSS.n42 VSS.n41 585
R700 VSS.n173 VSS.n172 585
R701 VSS.n174 VSS.n173 585
R702 VSS.n39 VSS.n38 585
R703 VSS.n175 VSS.n39 585
R704 VSS.n181 VSS.n180 585
R705 VSS.n180 VSS.n179 585
R706 VSS.n40 VSS.n36 585
R707 VSS.n178 VSS.n40 585
R708 VSS.n185 VSS.n35 585
R709 VSS.n177 VSS.n35 585
R710 VSS.n187 VSS.n186 585
R711 VSS.n187 VSS.n13 585
R712 VSS.n254 VSS.n10 585
R713 VSS.n13 VSS.n10 585
R714 VSS.n255 VSS.n9 585
R715 VSS.n177 VSS.n9 585
R716 VSS.n256 VSS.n8 585
R717 VSS.n178 VSS.n8 585
R718 VSS.n176 VSS.n6 585
R719 VSS.n179 VSS.n176 585
R720 VSS.n260 VSS.n5 585
R721 VSS.n175 VSS.n5 585
R722 VSS.n261 VSS.n4 585
R723 VSS.n174 VSS.n4 585
R724 VSS.n262 VSS.n3 585
R725 VSS.n41 VSS.n3 585
R726 VSS.n165 VSS.n2 585
R727 VSS.n166 VSS.n165 585
R728 VSS.n164 VSS.n48 585
R729 VSS.n164 VSS.n163 585
R730 VSS.n148 VSS.n47 585
R731 VSS.n162 VSS.n47 585
R732 VSS.n58 VSS.n56 585
R733 VSS.n56 VSS.n49 585
R734 VSS.n153 VSS.n152 585
R735 VSS.n154 VSS.n153 585
R736 VSS.n57 VSS.n55 585
R737 VSS.n75 VSS.n55 585
R738 VSS.n252 VSS.n251 585
R739 VSS.n12 VSS.n11 585
R740 VSS.n247 VSS.n246 585
R741 VSS.n244 VSS.n28 585
R742 VSS.n243 VSS.n242 585
R743 VSS.n241 VSS.n240 585
R744 VSS.n239 VSS.n238 585
R745 VSS.n237 VSS.n236 585
R746 VSS.n235 VSS.n234 585
R747 VSS.n233 VSS.n232 585
R748 VSS.n231 VSS.n230 585
R749 VSS.n229 VSS.n228 585
R750 VSS.n227 VSS.n226 585
R751 VSS.n225 VSS.n224 585
R752 VSS.n223 VSS.n222 585
R753 VSS.n221 VSS.n220 585
R754 VSS.n219 VSS.n218 585
R755 VSS.n217 VSS.n216 585
R756 VSS.n215 VSS.n214 585
R757 VSS.n213 VSS.n212 585
R758 VSS.n211 VSS.n210 585
R759 VSS.n209 VSS.n208 585
R760 VSS.n207 VSS.n206 585
R761 VSS.n205 VSS.n204 585
R762 VSS.n203 VSS.n202 585
R763 VSS.n201 VSS.n200 585
R764 VSS.n199 VSS.n198 585
R765 VSS.n197 VSS.n196 585
R766 VSS.n195 VSS.n194 585
R767 VSS.n193 VSS.n192 585
R768 VSS.n191 VSS.n190 585
R769 VSS.n189 VSS.n188 585
R770 VSS.n141 VSS.n140 585
R771 VSS.n139 VSS.n77 585
R772 VSS.n138 VSS.n76 585
R773 VSS.n143 VSS.n76 585
R774 VSS.n137 VSS.n136 585
R775 VSS.n135 VSS.n134 585
R776 VSS.n133 VSS.n132 585
R777 VSS.n131 VSS.n130 585
R778 VSS.n129 VSS.n128 585
R779 VSS.n127 VSS.n126 585
R780 VSS.n125 VSS.n124 585
R781 VSS.n123 VSS.n122 585
R782 VSS.n121 VSS.n120 585
R783 VSS.n119 VSS.n118 585
R784 VSS.n117 VSS.n116 585
R785 VSS.n114 VSS.n113 585
R786 VSS.n112 VSS.n111 585
R787 VSS.n110 VSS.n109 585
R788 VSS.n108 VSS.n107 585
R789 VSS.n106 VSS.n105 585
R790 VSS.n104 VSS.n103 585
R791 VSS.n102 VSS.n101 585
R792 VSS.n100 VSS.n99 585
R793 VSS.n98 VSS.n97 585
R794 VSS.n96 VSS.n95 585
R795 VSS.n94 VSS.n93 585
R796 VSS.n92 VSS.n91 585
R797 VSS.n90 VSS.n89 585
R798 VSS.n88 VSS.n87 585
R799 VSS.n86 VSS.n85 585
R800 VSS.n84 VSS.n83 585
R801 VSS.n60 VSS.n59 585
R802 VSS.n145 VSS.n144 585
R803 VSS.n144 VSS.n143 585
R804 VSS.n143 VSS.n75 321.329
R805 VSS.n249 VSS.n13 321.329
R806 VSS.n250 VSS.n249 256.663
R807 VSS.n249 VSS.n248 256.663
R808 VSS.n249 VSS.n27 256.663
R809 VSS.n249 VSS.n26 256.663
R810 VSS.n249 VSS.n25 256.663
R811 VSS.n249 VSS.n24 256.663
R812 VSS.n249 VSS.n23 256.663
R813 VSS.n249 VSS.n22 256.663
R814 VSS.n249 VSS.n21 256.663
R815 VSS.n249 VSS.n20 256.663
R816 VSS.n249 VSS.n19 256.663
R817 VSS.n249 VSS.n18 256.663
R818 VSS.n249 VSS.n17 256.663
R819 VSS.n249 VSS.n16 256.663
R820 VSS.n249 VSS.n15 256.663
R821 VSS.n249 VSS.n14 256.663
R822 VSS.n143 VSS.n142 256.663
R823 VSS.n143 VSS.n61 256.663
R824 VSS.n143 VSS.n62 256.663
R825 VSS.n143 VSS.n63 256.663
R826 VSS.n143 VSS.n64 256.663
R827 VSS.n143 VSS.n65 256.663
R828 VSS.n143 VSS.n66 256.663
R829 VSS.n143 VSS.n67 256.663
R830 VSS.n143 VSS.n68 256.663
R831 VSS.n143 VSS.n69 256.663
R832 VSS.n143 VSS.n70 256.663
R833 VSS.n143 VSS.n71 256.663
R834 VSS.n143 VSS.n72 256.663
R835 VSS.n143 VSS.n73 256.663
R836 VSS.n143 VSS.n74 256.663
R837 VSS.n155 VSS.n54 240.244
R838 VSS.n155 VSS.n50 240.244
R839 VSS.n161 VSS.n50 240.244
R840 VSS.n161 VSS.n46 240.244
R841 VSS.n167 VSS.n46 240.244
R842 VSS.n167 VSS.n42 240.244
R843 VSS.n173 VSS.n42 240.244
R844 VSS.n173 VSS.n39 240.244
R845 VSS.n180 VSS.n39 240.244
R846 VSS.n180 VSS.n40 240.244
R847 VSS.n40 VSS.n35 240.244
R848 VSS.n187 VSS.n35 240.244
R849 VSS.n153 VSS.n55 240.244
R850 VSS.n153 VSS.n56 240.244
R851 VSS.n56 VSS.n47 240.244
R852 VSS.n164 VSS.n47 240.244
R853 VSS.n165 VSS.n164 240.244
R854 VSS.n165 VSS.n3 240.244
R855 VSS.n4 VSS.n3 240.244
R856 VSS.n5 VSS.n4 240.244
R857 VSS.n176 VSS.n5 240.244
R858 VSS.n176 VSS.n8 240.244
R859 VSS.n9 VSS.n8 240.244
R860 VSS.n10 VSS.n9 240.244
R861 VSS.n154 VSS.n49 170.016
R862 VSS.n162 VSS.n49 170.016
R863 VSS.n163 VSS.n162 170.016
R864 VSS.n174 VSS.n41 170.016
R865 VSS.n179 VSS.n175 170.016
R866 VSS.n179 VSS.n178 170.016
R867 VSS.n177 VSS.n13 170.016
R868 VSS.n175 VSS.t2 166.615
R869 VSS.n77 VSS.n76 163.367
R870 VSS.n136 VSS.n76 163.367
R871 VSS.n134 VSS.n133 163.367
R872 VSS.n130 VSS.n129 163.367
R873 VSS.n126 VSS.n125 163.367
R874 VSS.n122 VSS.n121 163.367
R875 VSS.n118 VSS.n117 163.367
R876 VSS.n113 VSS.n112 163.367
R877 VSS.n109 VSS.n108 163.367
R878 VSS.n105 VSS.n104 163.367
R879 VSS.n101 VSS.n100 163.367
R880 VSS.n97 VSS.n96 163.367
R881 VSS.n93 VSS.n92 163.367
R882 VSS.n89 VSS.n88 163.367
R883 VSS.n85 VSS.n84 163.367
R884 VSS.n144 VSS.n60 163.367
R885 VSS.n192 VSS.n191 163.367
R886 VSS.n196 VSS.n195 163.367
R887 VSS.n200 VSS.n199 163.367
R888 VSS.n204 VSS.n203 163.367
R889 VSS.n208 VSS.n207 163.367
R890 VSS.n212 VSS.n211 163.367
R891 VSS.n216 VSS.n215 163.367
R892 VSS.n220 VSS.n219 163.367
R893 VSS.n224 VSS.n223 163.367
R894 VSS.n228 VSS.n227 163.367
R895 VSS.n232 VSS.n231 163.367
R896 VSS.n236 VSS.n235 163.367
R897 VSS.n240 VSS.n239 163.367
R898 VSS.n242 VSS.n28 163.367
R899 VSS.n247 VSS.n12 163.367
R900 VSS.n75 VSS.t8 159.815
R901 VSS.n166 VSS.t1 122.412
R902 VSS.n166 VSS.t0 98.6095
R903 VSS.n31 VSS.t5 96.619
R904 VSS.n29 VSS.t12 96.619
R905 VSS.n80 VSS.t16 96.619
R906 VSS.n78 VSS.t10 96.619
R907 VSS.n178 VSS.t4 85.0082
R908 VSS.t4 VSS.n177 85.0082
R909 VSS.n32 VSS.t6 84.013
R910 VSS.n30 VSS.t13 84.013
R911 VSS.n81 VSS.t15 84.013
R912 VSS.n79 VSS.t9 84.013
R913 VSS.n142 VSS.n141 71.676
R914 VSS.n136 VSS.n61 71.676
R915 VSS.n133 VSS.n62 71.676
R916 VSS.n129 VSS.n63 71.676
R917 VSS.n125 VSS.n64 71.676
R918 VSS.n121 VSS.n65 71.676
R919 VSS.n117 VSS.n66 71.676
R920 VSS.n112 VSS.n67 71.676
R921 VSS.n108 VSS.n68 71.676
R922 VSS.n104 VSS.n69 71.676
R923 VSS.n100 VSS.n70 71.676
R924 VSS.n96 VSS.n71 71.676
R925 VSS.n92 VSS.n72 71.676
R926 VSS.n88 VSS.n73 71.676
R927 VSS.n84 VSS.n74 71.676
R928 VSS.n191 VSS.n14 71.676
R929 VSS.n195 VSS.n15 71.676
R930 VSS.n199 VSS.n16 71.676
R931 VSS.n203 VSS.n17 71.676
R932 VSS.n207 VSS.n18 71.676
R933 VSS.n211 VSS.n19 71.676
R934 VSS.n215 VSS.n20 71.676
R935 VSS.n219 VSS.n21 71.676
R936 VSS.n223 VSS.n22 71.676
R937 VSS.n227 VSS.n23 71.676
R938 VSS.n231 VSS.n24 71.676
R939 VSS.n235 VSS.n25 71.676
R940 VSS.n239 VSS.n26 71.676
R941 VSS.n242 VSS.n27 71.676
R942 VSS.n248 VSS.n247 71.676
R943 VSS.n251 VSS.n250 71.676
R944 VSS.n250 VSS.n12 71.676
R945 VSS.n248 VSS.n28 71.676
R946 VSS.n240 VSS.n27 71.676
R947 VSS.n236 VSS.n26 71.676
R948 VSS.n232 VSS.n25 71.676
R949 VSS.n228 VSS.n24 71.676
R950 VSS.n224 VSS.n23 71.676
R951 VSS.n220 VSS.n22 71.676
R952 VSS.n216 VSS.n21 71.676
R953 VSS.n212 VSS.n20 71.676
R954 VSS.n208 VSS.n19 71.676
R955 VSS.n204 VSS.n18 71.676
R956 VSS.n200 VSS.n17 71.676
R957 VSS.n196 VSS.n16 71.676
R958 VSS.n192 VSS.n15 71.676
R959 VSS.n188 VSS.n14 71.676
R960 VSS.n142 VSS.n77 71.676
R961 VSS.n134 VSS.n61 71.676
R962 VSS.n130 VSS.n62 71.676
R963 VSS.n126 VSS.n63 71.676
R964 VSS.n122 VSS.n64 71.676
R965 VSS.n118 VSS.n65 71.676
R966 VSS.n113 VSS.n66 71.676
R967 VSS.n109 VSS.n67 71.676
R968 VSS.n105 VSS.n68 71.676
R969 VSS.n101 VSS.n69 71.676
R970 VSS.n97 VSS.n70 71.676
R971 VSS.n93 VSS.n71 71.676
R972 VSS.n89 VSS.n72 71.676
R973 VSS.n85 VSS.n73 71.676
R974 VSS.n74 VSS.n60 71.676
R975 VSS.n163 VSS.t0 71.407
R976 VSS.t1 VSS.n41 47.6048
R977 VSS.n33 VSS.n32 45.1884
R978 VSS.n245 VSS.n30 45.1884
R979 VSS.n82 VSS.n81 34.3278
R980 VSS.n115 VSS.n79 34.3278
R981 VSS.n189 VSS.n34 27.5398
R982 VSS.n253 VSS.n252 27.5398
R983 VSS.n140 VSS.n52 27.5398
R984 VSS.n146 VSS.n145 27.5398
R985 VSS.n156 VSS.n53 19.3944
R986 VSS.n156 VSS.n51 19.3944
R987 VSS.n160 VSS.n51 19.3944
R988 VSS.n160 VSS.n45 19.3944
R989 VSS.n168 VSS.n45 19.3944
R990 VSS.n168 VSS.n43 19.3944
R991 VSS.n172 VSS.n43 19.3944
R992 VSS.n172 VSS.n38 19.3944
R993 VSS.n181 VSS.n38 19.3944
R994 VSS.n181 VSS.n36 19.3944
R995 VSS.n185 VSS.n36 19.3944
R996 VSS.n186 VSS.n185 19.3944
R997 VSS.n152 VSS.n57 19.3944
R998 VSS.n152 VSS.n58 19.3944
R999 VSS.n148 VSS.n58 19.3944
R1000 VSS.n148 VSS.n48 19.3944
R1001 VSS.n48 VSS.n2 19.3944
R1002 VSS.n262 VSS.n2 19.3944
R1003 VSS.n262 VSS.n261 19.3944
R1004 VSS.n261 VSS.n260 19.3944
R1005 VSS.n260 VSS.n6 19.3944
R1006 VSS.n256 VSS.n6 19.3944
R1007 VSS.n256 VSS.n255 19.3944
R1008 VSS.n255 VSS.n254 19.3944
R1009 VSS.n32 VSS.n31 12.6066
R1010 VSS.n30 VSS.n29 12.6066
R1011 VSS.n81 VSS.n80 12.6066
R1012 VSS.n79 VSS.n78 12.6066
R1013 VSS.n190 VSS.n189 10.6151
R1014 VSS.n193 VSS.n190 10.6151
R1015 VSS.n194 VSS.n193 10.6151
R1016 VSS.n197 VSS.n194 10.6151
R1017 VSS.n198 VSS.n197 10.6151
R1018 VSS.n201 VSS.n198 10.6151
R1019 VSS.n202 VSS.n201 10.6151
R1020 VSS.n205 VSS.n202 10.6151
R1021 VSS.n206 VSS.n205 10.6151
R1022 VSS.n209 VSS.n206 10.6151
R1023 VSS.n210 VSS.n209 10.6151
R1024 VSS.n213 VSS.n210 10.6151
R1025 VSS.n214 VSS.n213 10.6151
R1026 VSS.n218 VSS.n217 10.6151
R1027 VSS.n221 VSS.n218 10.6151
R1028 VSS.n222 VSS.n221 10.6151
R1029 VSS.n225 VSS.n222 10.6151
R1030 VSS.n226 VSS.n225 10.6151
R1031 VSS.n229 VSS.n226 10.6151
R1032 VSS.n230 VSS.n229 10.6151
R1033 VSS.n233 VSS.n230 10.6151
R1034 VSS.n234 VSS.n233 10.6151
R1035 VSS.n237 VSS.n234 10.6151
R1036 VSS.n238 VSS.n237 10.6151
R1037 VSS.n241 VSS.n238 10.6151
R1038 VSS.n243 VSS.n241 10.6151
R1039 VSS.n244 VSS.n243 10.6151
R1040 VSS.n246 VSS.n11 10.6151
R1041 VSS.n252 VSS.n11 10.6151
R1042 VSS.n140 VSS.n139 10.6151
R1043 VSS.n139 VSS.n138 10.6151
R1044 VSS.n138 VSS.n137 10.6151
R1045 VSS.n137 VSS.n135 10.6151
R1046 VSS.n135 VSS.n132 10.6151
R1047 VSS.n132 VSS.n131 10.6151
R1048 VSS.n131 VSS.n128 10.6151
R1049 VSS.n128 VSS.n127 10.6151
R1050 VSS.n127 VSS.n124 10.6151
R1051 VSS.n124 VSS.n123 10.6151
R1052 VSS.n123 VSS.n120 10.6151
R1053 VSS.n120 VSS.n119 10.6151
R1054 VSS.n119 VSS.n116 10.6151
R1055 VSS.n114 VSS.n111 10.6151
R1056 VSS.n111 VSS.n110 10.6151
R1057 VSS.n110 VSS.n107 10.6151
R1058 VSS.n107 VSS.n106 10.6151
R1059 VSS.n106 VSS.n103 10.6151
R1060 VSS.n103 VSS.n102 10.6151
R1061 VSS.n102 VSS.n99 10.6151
R1062 VSS.n99 VSS.n98 10.6151
R1063 VSS.n98 VSS.n95 10.6151
R1064 VSS.n95 VSS.n94 10.6151
R1065 VSS.n94 VSS.n91 10.6151
R1066 VSS.n91 VSS.n90 10.6151
R1067 VSS.n90 VSS.n87 10.6151
R1068 VSS.n87 VSS.n86 10.6151
R1069 VSS.n83 VSS.n59 10.6151
R1070 VSS.n145 VSS.n59 10.6151
R1071 VSS.n154 VSS.t8 10.2014
R1072 VSS.n217 VSS.n33 9.83465
R1073 VSS.n115 VSS.n114 9.83465
R1074 VSS.n261 VSS.n0 9.3005
R1075 VSS.n260 VSS.n259 9.3005
R1076 VSS.n258 VSS.n6 9.3005
R1077 VSS.n257 VSS.n256 9.3005
R1078 VSS.n255 VSS.n7 9.3005
R1079 VSS.n254 VSS.n253 9.3005
R1080 VSS.n53 VSS.n52 9.3005
R1081 VSS.n157 VSS.n156 9.3005
R1082 VSS.n158 VSS.n51 9.3005
R1083 VSS.n160 VSS.n159 9.3005
R1084 VSS.n45 VSS.n44 9.3005
R1085 VSS.n169 VSS.n168 9.3005
R1086 VSS.n170 VSS.n43 9.3005
R1087 VSS.n172 VSS.n171 9.3005
R1088 VSS.n38 VSS.n37 9.3005
R1089 VSS.n182 VSS.n181 9.3005
R1090 VSS.n183 VSS.n36 9.3005
R1091 VSS.n185 VSS.n184 9.3005
R1092 VSS.n186 VSS.n34 9.3005
R1093 VSS.n152 VSS.n151 9.3005
R1094 VSS.n150 VSS.n58 9.3005
R1095 VSS.n149 VSS.n148 9.3005
R1096 VSS.n147 VSS.n48 9.3005
R1097 VSS.n2 VSS.n1 9.3005
R1098 VSS.n146 VSS.n57 9.3005
R1099 VSS.n263 VSS.n262 9.3005
R1100 VSS.n245 VSS.n244 5.77611
R1101 VSS.n86 VSS.n82 5.77611
R1102 VSS.n246 VSS.n245 4.83952
R1103 VSS.n83 VSS.n82 4.83952
R1104 VSS.t2 VSS.n174 3.40081
R1105 VSS.n214 VSS.n33 0.780988
R1106 VSS.n116 VSS.n115 0.780988
R1107 VSS.n259 VSS.n0 0.152939
R1108 VSS.n259 VSS.n258 0.152939
R1109 VSS.n258 VSS.n257 0.152939
R1110 VSS.n257 VSS.n7 0.152939
R1111 VSS.n253 VSS.n7 0.152939
R1112 VSS.n157 VSS.n52 0.152939
R1113 VSS.n158 VSS.n157 0.152939
R1114 VSS.n159 VSS.n158 0.152939
R1115 VSS.n159 VSS.n44 0.152939
R1116 VSS.n169 VSS.n44 0.152939
R1117 VSS.n170 VSS.n169 0.152939
R1118 VSS.n171 VSS.n170 0.152939
R1119 VSS.n171 VSS.n37 0.152939
R1120 VSS.n182 VSS.n37 0.152939
R1121 VSS.n183 VSS.n182 0.152939
R1122 VSS.n184 VSS.n183 0.152939
R1123 VSS.n184 VSS.n34 0.152939
R1124 VSS.n151 VSS.n146 0.152939
R1125 VSS.n151 VSS.n150 0.152939
R1126 VSS.n150 VSS.n149 0.152939
R1127 VSS.n149 VSS.n147 0.152939
R1128 VSS.n147 VSS.n1 0.152939
R1129 VSS.n263 VSS.n1 0.13922
R1130 VSS VSS.n0 0.0767195
R1131 VSS VSS.n263 0.063
C0 VCC VOUT 5.95364f
C1 VOUT VSS 6.306905f
C2 VGP VSS 0.042695f
C3 VGN VSS 0.030294f
C4 VIN VSS 0.020764f
C5 VCC VSS 21.049017f
C6 VCC.n0 VSS 0.00367f
C7 VCC.n1 VSS 0.004894f
C8 VCC.n2 VSS 0.003939f
C9 VCC.n3 VSS 0.004894f
C10 VCC.n4 VSS 0.004894f
C11 VCC.n5 VSS 0.004894f
C12 VCC.n6 VSS 0.003939f
C13 VCC.n7 VSS 0.004894f
C14 VCC.n8 VSS 0.004894f
C15 VCC.n9 VSS 0.004894f
C16 VCC.n10 VSS 0.00872f
C17 VCC.n11 VSS 0.003328f
C18 VCC.n12 VSS 0.003328f
C19 VCC.n13 VSS 0.289581f
C20 VCC.n37 VSS 0.003328f
C21 VCC.t3 VSS 0.09327f
C22 VCC.t2 VSS 0.095829f
C23 VCC.t0 VSS 0.016842f
C24 VCC.n38 VSS 0.033821f
C25 VCC.n39 VSS 0.029355f
C26 VCC.t10 VSS 0.09327f
C27 VCC.t9 VSS 0.095829f
C28 VCC.t8 VSS 0.016842f
C29 VCC.n40 VSS 0.033821f
C30 VCC.n41 VSS 0.029355f
C31 VCC.n42 VSS 0.00574f
C32 VCC.n43 VSS 0.015393f
C33 VCC.n44 VSS 0.004894f
C34 VCC.n45 VSS 0.003939f
C35 VCC.n46 VSS 0.004894f
C36 VCC.n47 VSS 0.003939f
C37 VCC.n48 VSS 0.004894f
C38 VCC.n49 VSS 0.004894f
C39 VCC.n50 VSS 0.140937f
C40 VCC.n51 VSS 0.004894f
C41 VCC.n52 VSS 0.003939f
C42 VCC.n53 VSS 0.004894f
C43 VCC.n54 VSS 0.003939f
C44 VCC.n55 VSS 0.004894f
C45 VCC.t15 VSS 0.110107f
C46 VCC.t16 VSS 0.110107f
C47 VCC.n56 VSS 0.004894f
C48 VCC.n57 VSS 0.003939f
C49 VCC.n58 VSS 0.220213f
C50 VCC.n59 VSS 0.004894f
C51 VCC.n60 VSS 0.003939f
C52 VCC.n61 VSS 0.015393f
C53 VCC.n62 VSS 0.003269f
C54 VCC.n63 VSS 0.00872f
C55 VCC.t5 VSS 0.110107f
C56 VCC.n64 VSS 0.00872f
C57 VCC.n65 VSS 0.004894f
C58 VCC.n66 VSS 0.003269f
C59 VCC.n67 VSS 0.003939f
C60 VCC.n68 VSS 0.003328f
C61 VCC.n69 VSS 0.003328f
C62 VCC.n93 VSS 0.282974f
C63 VCC.n94 VSS 0.003328f
C64 VCC.t6 VSS 0.09327f
C65 VCC.t7 VSS 0.095829f
C66 VCC.t4 VSS 0.016842f
C67 VCC.n95 VSS 0.033821f
C68 VCC.n96 VSS 0.028252f
C69 VCC.t12 VSS 0.09327f
C70 VCC.t13 VSS 0.095829f
C71 VCC.t11 VSS 0.016842f
C72 VCC.n97 VSS 0.033821f
C73 VCC.n98 VSS 0.028252f
C74 VCC.n99 VSS 0.004638f
C75 VCC.n100 VSS 0.00875f
C76 VCC.n101 VSS 0.00609f
C77 VCC.n102 VSS 0.003328f
C78 VCC.n103 VSS 0.003328f
C79 VCC.n104 VSS 0.003328f
C80 VCC.n105 VSS 0.003328f
C81 VCC.n106 VSS 0.003328f
C82 VCC.n107 VSS 0.003328f
C83 VCC.n108 VSS 0.003328f
C84 VCC.n109 VSS 0.003328f
C85 VCC.n110 VSS 0.003328f
C86 VCC.n111 VSS 0.003328f
C87 VCC.n112 VSS 0.003328f
C88 VCC.n113 VSS 0.003328f
C89 VCC.n114 VSS 0.003328f
C90 VCC.n115 VSS 0.003328f
C91 VCC.n116 VSS 0.003328f
C92 VCC.n117 VSS 0.003328f
C93 VCC.n118 VSS 0.003328f
C94 VCC.n119 VSS 0.003328f
C95 VCC.n120 VSS 0.003328f
C96 VCC.n121 VSS 0.003328f
C97 VCC.n122 VSS 0.003328f
C98 VCC.n123 VSS 0.003328f
C99 VCC.n124 VSS 0.003328f
C100 VCC.n125 VSS 0.003328f
C101 VCC.n126 VSS 0.003328f
C102 VCC.n127 VSS 0.003328f
C103 VCC.n128 VSS 0.003328f
C104 VCC.n129 VSS 0.003328f
C105 VCC.n130 VSS 0.003328f
C106 VCC.n131 VSS 0.003328f
C107 VCC.n132 VSS 0.003328f
C108 VCC.n133 VSS 0.003328f
C109 VCC.n134 VSS 0.003328f
C110 VCC.n135 VSS 0.003328f
C111 VCC.n136 VSS 0.003328f
C112 VCC.n137 VSS 0.003328f
C113 VCC.n138 VSS 0.003328f
C114 VCC.n139 VSS 0.003328f
C115 VCC.n140 VSS 0.003328f
C116 VCC.n141 VSS 0.003328f
C117 VCC.n142 VSS 0.002618f
C118 VCC.n143 VSS 0.003328f
C119 VCC.n144 VSS 0.003328f
C120 VCC.n145 VSS 0.002373f
C121 VCC.n146 VSS 0.003328f
C122 VCC.n147 VSS 0.003328f
C123 VCC.n148 VSS 0.003328f
C124 VCC.n149 VSS 0.003328f
C125 VCC.n150 VSS 0.003328f
C126 VCC.n151 VSS 0.003328f
C127 VCC.n152 VSS 0.003328f
C128 VCC.n153 VSS 0.003328f
C129 VCC.n154 VSS 0.003328f
C130 VCC.n155 VSS 0.003328f
C131 VCC.n156 VSS 0.003328f
C132 VCC.n157 VSS 0.003328f
C133 VCC.n158 VSS 0.003328f
C134 VCC.n159 VSS 0.003328f
C135 VCC.n160 VSS 0.003328f
C136 VCC.n161 VSS 0.003328f
C137 VCC.n162 VSS 0.003328f
C138 VCC.n163 VSS 0.003328f
C139 VCC.n164 VSS 0.003328f
C140 VCC.n165 VSS 0.003328f
C141 VCC.n166 VSS 0.003328f
C142 VCC.n167 VSS 0.003328f
C143 VCC.n168 VSS 0.003328f
C144 VCC.n169 VSS 0.003328f
C145 VCC.n170 VSS 0.003328f
C146 VCC.n171 VSS 0.003328f
C147 VCC.n172 VSS 0.003328f
C148 VCC.n173 VSS 0.003328f
C149 VCC.n174 VSS 0.003328f
C150 VCC.n175 VSS 0.003328f
C151 VCC.n176 VSS 0.003328f
C152 VCC.n177 VSS 0.003328f
C153 VCC.n178 VSS 0.003328f
C154 VCC.n179 VSS 0.003328f
C155 VCC.n180 VSS 0.003328f
C156 VCC.n181 VSS 0.003328f
C157 VCC.n182 VSS 0.003328f
C158 VCC.n183 VSS 0.003328f
C159 VCC.n184 VSS 0.003328f
C160 VCC.n185 VSS 0.003328f
C161 VCC.n186 VSS 0.003328f
C162 VCC.n187 VSS 0.003328f
C163 VCC.n188 VSS 0.003328f
C164 VCC.n189 VSS 0.003328f
C165 VCC.n190 VSS 0.003107f
C166 VCC.n191 VSS 0.004638f
C167 VCC.n192 VSS 0.001884f
C168 VCC.n193 VSS 0.003328f
C169 VCC.n194 VSS 0.406294f
C170 VCC.n196 VSS 0.00875f
C171 VCC.n197 VSS 0.00609f
C172 VCC.n198 VSS 0.015393f
C173 VCC.n199 VSS 0.004894f
C174 VCC.n200 VSS 0.003939f
C175 VCC.n201 VSS 0.004894f
C176 VCC.n202 VSS 0.004894f
C177 VCC.n203 VSS 0.004894f
C178 VCC.n204 VSS 0.003939f
C179 VCC.n205 VSS 0.004894f
C180 VCC.n206 VSS 0.116713f
C181 VCC.n207 VSS 0.004894f
C182 VCC.n208 VSS 0.003939f
C183 VCC.n209 VSS 0.004894f
C184 VCC.n210 VSS 0.004894f
C185 VCC.n211 VSS 0.004894f
C186 VCC.n212 VSS 0.003939f
C187 VCC.n213 VSS 0.004894f
C188 VCC.n214 VSS 0.220213f
C189 VCC.n215 VSS 0.156352f
C190 VCC.n216 VSS 0.004894f
C191 VCC.n217 VSS 0.004894f
C192 VCC.n218 VSS 0.143139f
C193 VCC.n219 VSS 0.004894f
C194 VCC.n220 VSS 0.003939f
C195 VCC.n221 VSS 0.004894f
C196 VCC.n222 VSS 0.004894f
C197 VCC.n223 VSS 0.004894f
C198 VCC.n224 VSS 0.003939f
C199 VCC.n225 VSS 0.004894f
C200 VCC.n226 VSS 0.112309f
C201 VCC.t14 VSS 0.110107f
C202 VCC.n227 VSS 0.218011f
C203 VCC.n228 VSS 0.16516f
C204 VCC.t1 VSS 0.110107f
C205 VCC.n229 VSS 0.16516f
C206 VCC.n230 VSS 0.004894f
C207 VCC.n231 VSS 0.220213f
C208 VCC.n232 VSS 0.004894f
C209 VCC.n233 VSS 0.003939f
C210 VCC.n234 VSS 0.004894f
C211 VCC.n235 VSS 0.004894f
C212 VCC.n236 VSS 0.004894f
C213 VCC.n237 VSS 0.003939f
C214 VCC.n238 VSS 0.003269f
C215 VCC.n239 VSS 0.00872f
C216 VCC.n240 VSS 0.00875f
C217 VCC.n241 VSS 0.00609f
C218 VCC.n242 VSS 0.003328f
C219 VCC.n243 VSS 0.003328f
C220 VCC.n244 VSS 0.003328f
C221 VCC.n245 VSS 0.003328f
C222 VCC.n246 VSS 0.003328f
C223 VCC.n247 VSS 0.003328f
C224 VCC.n248 VSS 0.003328f
C225 VCC.n249 VSS 0.003328f
C226 VCC.n250 VSS 0.003328f
C227 VCC.n251 VSS 0.003328f
C228 VCC.n252 VSS 0.003328f
C229 VCC.n253 VSS 0.003328f
C230 VCC.n254 VSS 0.003328f
C231 VCC.n255 VSS 0.003328f
C232 VCC.n256 VSS 0.003328f
C233 VCC.n257 VSS 0.003328f
C234 VCC.n258 VSS 0.003328f
C235 VCC.n259 VSS 0.003328f
C236 VCC.n260 VSS 0.003328f
C237 VCC.n261 VSS 0.003328f
C238 VCC.n262 VSS 0.003328f
C239 VCC.n263 VSS 0.003328f
C240 VCC.n264 VSS 0.003328f
C241 VCC.n265 VSS 0.003328f
C242 VCC.n266 VSS 0.003328f
C243 VCC.n267 VSS 0.003328f
C244 VCC.n268 VSS 0.003328f
C245 VCC.n269 VSS 0.003328f
C246 VCC.n270 VSS 0.003328f
C247 VCC.n271 VSS 0.003328f
C248 VCC.n272 VSS 0.003328f
C249 VCC.n273 VSS 0.003328f
C250 VCC.n274 VSS 0.003328f
C251 VCC.n275 VSS 0.003328f
C252 VCC.n276 VSS 0.003328f
C253 VCC.n277 VSS 0.003328f
C254 VCC.n278 VSS 0.003328f
C255 VCC.n279 VSS 0.003328f
C256 VCC.n280 VSS 0.003328f
C257 VCC.n281 VSS 0.003328f
C258 VCC.n282 VSS 0.002618f
C259 VCC.n283 VSS 0.003328f
C260 VCC.n284 VSS 0.003328f
C261 VCC.n285 VSS 0.002373f
C262 VCC.n286 VSS 0.003328f
C263 VCC.n287 VSS 0.003328f
C264 VCC.n288 VSS 0.003328f
C265 VCC.n289 VSS 0.003328f
C266 VCC.n290 VSS 0.003328f
C267 VCC.n291 VSS 0.003328f
C268 VCC.n292 VSS 0.003328f
C269 VCC.n293 VSS 0.003328f
C270 VCC.n294 VSS 0.003328f
C271 VCC.n295 VSS 0.003328f
C272 VCC.n296 VSS 0.003328f
C273 VCC.n297 VSS 0.003328f
C274 VCC.n298 VSS 0.003328f
C275 VCC.n299 VSS 0.003328f
C276 VCC.n300 VSS 0.003328f
C277 VCC.n301 VSS 0.003328f
C278 VCC.n302 VSS 0.003328f
C279 VCC.n303 VSS 0.003328f
C280 VCC.n304 VSS 0.003328f
C281 VCC.n305 VSS 0.003328f
C282 VCC.n306 VSS 0.003328f
C283 VCC.n307 VSS 0.003328f
C284 VCC.n308 VSS 0.003328f
C285 VCC.n309 VSS 0.003328f
C286 VCC.n310 VSS 0.003328f
C287 VCC.n311 VSS 0.003328f
C288 VCC.n312 VSS 0.003328f
C289 VCC.n313 VSS 0.003328f
C290 VCC.n314 VSS 0.003328f
C291 VCC.n315 VSS 0.003328f
C292 VCC.n316 VSS 0.003328f
C293 VCC.n317 VSS 0.003328f
C294 VCC.n318 VSS 0.003328f
C295 VCC.n319 VSS 0.003328f
C296 VCC.n320 VSS 0.003328f
C297 VCC.n321 VSS 0.003328f
C298 VCC.n322 VSS 0.003328f
C299 VCC.n323 VSS 0.003328f
C300 VCC.n324 VSS 0.003328f
C301 VCC.n325 VSS 0.003328f
C302 VCC.n326 VSS 0.003328f
C303 VCC.n327 VSS 0.003328f
C304 VCC.n328 VSS 0.003328f
C305 VCC.n329 VSS 0.003328f
C306 VCC.n330 VSS 0.003107f
C307 VCC.n331 VSS 0.00574f
C308 VCC.n332 VSS 0.001884f
C309 VCC.n333 VSS 0.003328f
C310 VCC.n335 VSS 0.406294f
C311 VCC.n336 VSS 0.00875f
C312 VCC.n337 VSS 0.00609f
C313 VCC.n338 VSS 0.015393f
C314 VCC.n339 VSS 0.003269f
C315 VCC.n340 VSS 0.003939f
C316 VCC.n341 VSS 0.003939f
C317 VCC.n342 VSS 0.004894f
C318 VCC.n343 VSS 0.004894f
C319 VCC.n344 VSS 0.004894f
C320 VCC.n345 VSS 0.003939f
C321 VCC.n346 VSS 0.003939f
C322 VCC.n347 VSS 0.003939f
C323 VCC.n348 VSS 0.004476f
C324 VOUT.t21 VSS 0.017102f
C325 VOUT.n0 VSS 0.016075f
C326 VOUT.t24 VSS 0.017102f
C327 VOUT.t5 VSS 0.01619f
C328 VOUT.n1 VSS 0.011315f
C329 VOUT.n2 VSS 0.016056f
C330 VOUT.n3 VSS 0.027049f
C331 VOUT.n4 VSS 0.078678f
C332 VOUT.t23 VSS 0.10253f
C333 VOUT.n5 VSS 0.082471f
C334 VOUT.t25 VSS 0.131722f
C335 VOUT.t22 VSS 0.017408f
C336 VOUT.n6 VSS 0.189468f
C337 VOUT.n7 VSS 0.08597f
C338 VOUT.t8 VSS 0.257314f
C339 VOUT.t20 VSS 0.257314f
C340 VOUT.t16 VSS 0.03266f
C341 VOUT.n8 VSS 0.021406f
C342 VOUT.t19 VSS 0.03266f
C343 VOUT.t26 VSS 0.031857f
C344 VOUT.n9 VSS 0.016538f
C345 VOUT.n10 VSS 0.021388f
C346 VOUT.n11 VSS 0.027049f
C347 VOUT.t13 VSS 0.017102f
C348 VOUT.n12 VSS 0.016075f
C349 VOUT.t0 VSS 0.017102f
C350 VOUT.t11 VSS 0.01619f
C351 VOUT.n13 VSS 0.011315f
C352 VOUT.n14 VSS 0.016056f
C353 VOUT.n15 VSS 0.048038f
C354 VOUT.n16 VSS 0.122651f
C355 VOUT.t2 VSS 0.03266f
C356 VOUT.n17 VSS 0.021406f
C357 VOUT.t7 VSS 0.03266f
C358 VOUT.t9 VSS 0.031857f
C359 VOUT.n18 VSS 0.016538f
C360 VOUT.n19 VSS 0.021388f
C361 VOUT.n20 VSS 0.048038f
C362 VOUT.n21 VSS 0.122651f
C363 VOUT.n22 VSS 0.113388f
C364 VOUT.t18 VSS 0.203109f
C365 VOUT.n23 VSS 0.134386f
C366 VOUT.n24 VSS 0.122158f
C367 VOUT.n25 VSS 0.158709f
C368 VOUT.t27 VSS 0.069632f
C369 VOUT.t17 VSS 0.034816f
C370 VOUT.n26 VSS 0.175881f
C371 VOUT.n27 VSS 0.199306f
C372 VOUT.n28 VSS 0.095832f
C373 VOUT.n29 VSS 0.293335f
C374 VOUT.t3 VSS 0.034816f
C375 VOUT.n30 VSS 0.175881f
C376 VOUT.t10 VSS 0.069632f
C377 VOUT.n31 VSS 0.15951f
C378 VOUT.t4 VSS 0.203109f
C379 VOUT.n32 VSS 0.242019f
C380 VOUT.n33 VSS 0.100345f
C381 VOUT.t1 VSS 0.131722f
C382 VOUT.t14 VSS 0.017408f
C383 VOUT.n34 VSS 0.094698f
C384 VOUT.t12 VSS 0.034816f
C385 VOUT.n35 VSS 0.085229f
C386 VOUT.t15 VSS 0.10253f
C387 VOUT.n36 VSS 0.143225f
C388 VOUT.n37 VSS 0.073189f
C389 VOUT.n38 VSS 0.058814f
C390 VOUT.n39 VSS 0.0815f
C391 VOUT.n40 VSS 0.11857f
C392 VOUT.n41 VSS 0.094698f
C393 VOUT.t6 VSS 0.034816f
C394 VOUT.n42 VSS 0.084686f
C395 VOUT.n43 VSS 0.055411f
.ends

