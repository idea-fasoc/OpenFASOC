* NGSPICE file created from diff_pair_sample_1544.ext - technology: sky130A

.subckt diff_pair_sample_1544 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.09735 pd=0.92 as=0.2301 ps=1.96 w=0.59 l=1.67
X1 VTAIL.t3 VP.t1 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2301 pd=1.96 as=0.09735 ps=0.92 w=0.59 l=1.67
X2 VDD1.t1 VP.t2 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.09735 pd=0.92 as=0.2301 ps=1.96 w=0.59 l=1.67
X3 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=0.2301 pd=1.96 as=0 ps=0 w=0.59 l=1.67
X4 VTAIL.t7 VN.t0 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2301 pd=1.96 as=0.09735 ps=0.92 w=0.59 l=1.67
X5 VTAIL.t5 VP.t3 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2301 pd=1.96 as=0.09735 ps=0.92 w=0.59 l=1.67
X6 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=0.2301 pd=1.96 as=0 ps=0 w=0.59 l=1.67
X7 VDD2.t2 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.09735 pd=0.92 as=0.2301 ps=1.96 w=0.59 l=1.67
X8 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2301 pd=1.96 as=0 ps=0 w=0.59 l=1.67
X9 VTAIL.t0 VN.t2 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2301 pd=1.96 as=0.09735 ps=0.92 w=0.59 l=1.67
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2301 pd=1.96 as=0 ps=0 w=0.59 l=1.67
X11 VDD2.t0 VN.t3 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.09735 pd=0.92 as=0.2301 ps=1.96 w=0.59 l=1.67
R0 VP.n8 VP.n0 161.3
R1 VP.n7 VP.n6 161.3
R2 VP.n5 VP.n1 161.3
R3 VP.n4 VP.n3 86.2894
R4 VP.n10 VP.n9 86.2894
R5 VP.n4 VP.n2 44.37
R6 VP.n2 VP.t3 43.0851
R7 VP.n2 VP.t2 42.6674
R8 VP.n7 VP.n1 40.4934
R9 VP.n8 VP.n7 40.4934
R10 VP.n3 VP.n1 24.4675
R11 VP.n9 VP.n8 24.4675
R12 VP.n9 VP.t0 8.51487
R13 VP.n3 VP.t1 8.51487
R14 VP.n5 VP.n4 0.278367
R15 VP.n10 VP.n0 0.278367
R16 VP.n6 VP.n5 0.189894
R17 VP.n6 VP.n0 0.189894
R18 VP VP.n10 0.153454
R19 VTAIL.n7 VTAIL.t6 250.55
R20 VTAIL.n0 VTAIL.t0 250.55
R21 VTAIL.n1 VTAIL.t2 250.55
R22 VTAIL.n2 VTAIL.t3 250.55
R23 VTAIL.n6 VTAIL.t4 250.55
R24 VTAIL.n5 VTAIL.t5 250.55
R25 VTAIL.n4 VTAIL.t1 250.55
R26 VTAIL.n3 VTAIL.t7 250.55
R27 VTAIL.n7 VTAIL.n6 14.5996
R28 VTAIL.n3 VTAIL.n2 14.5996
R29 VTAIL.n4 VTAIL.n3 1.72464
R30 VTAIL.n6 VTAIL.n5 1.72464
R31 VTAIL.n2 VTAIL.n1 1.72464
R32 VTAIL VTAIL.n0 0.920759
R33 VTAIL VTAIL.n7 0.804379
R34 VTAIL.n5 VTAIL.n4 0.470328
R35 VTAIL.n1 VTAIL.n0 0.470328
R36 VDD1 VDD1.n1 263.591
R37 VDD1 VDD1.n0 233.728
R38 VDD1.n0 VDD1.t0 33.5598
R39 VDD1.n0 VDD1.t1 33.5598
R40 VDD1.n1 VDD1.t2 33.5598
R41 VDD1.n1 VDD1.t3 33.5598
R42 B.n346 B.n345 585
R43 B.n117 B.n62 585
R44 B.n116 B.n115 585
R45 B.n114 B.n113 585
R46 B.n112 B.n111 585
R47 B.n110 B.n109 585
R48 B.n108 B.n107 585
R49 B.n106 B.n105 585
R50 B.n104 B.n103 585
R51 B.n102 B.n101 585
R52 B.n100 B.n99 585
R53 B.n98 B.n97 585
R54 B.n96 B.n95 585
R55 B.n94 B.n93 585
R56 B.n92 B.n91 585
R57 B.n90 B.n89 585
R58 B.n88 B.n87 585
R59 B.n86 B.n85 585
R60 B.n84 B.n83 585
R61 B.n82 B.n81 585
R62 B.n80 B.n79 585
R63 B.n78 B.n77 585
R64 B.n76 B.n75 585
R65 B.n74 B.n73 585
R66 B.n72 B.n71 585
R67 B.n70 B.n69 585
R68 B.n344 B.n49 585
R69 B.n349 B.n49 585
R70 B.n343 B.n48 585
R71 B.n350 B.n48 585
R72 B.n342 B.n341 585
R73 B.n341 B.n44 585
R74 B.n340 B.n43 585
R75 B.n356 B.n43 585
R76 B.n339 B.n42 585
R77 B.n357 B.n42 585
R78 B.n338 B.n41 585
R79 B.n358 B.n41 585
R80 B.n337 B.n336 585
R81 B.n336 B.n37 585
R82 B.n335 B.n36 585
R83 B.n364 B.n36 585
R84 B.n334 B.n35 585
R85 B.n365 B.n35 585
R86 B.n333 B.n34 585
R87 B.n366 B.n34 585
R88 B.n332 B.n331 585
R89 B.n331 B.n30 585
R90 B.n330 B.n29 585
R91 B.n372 B.n29 585
R92 B.n329 B.n28 585
R93 B.n373 B.n28 585
R94 B.n328 B.n27 585
R95 B.n374 B.n27 585
R96 B.n327 B.n326 585
R97 B.n326 B.n23 585
R98 B.n325 B.n22 585
R99 B.n380 B.n22 585
R100 B.n324 B.n21 585
R101 B.n381 B.n21 585
R102 B.n323 B.n20 585
R103 B.n382 B.n20 585
R104 B.n322 B.n321 585
R105 B.n321 B.n16 585
R106 B.n320 B.n15 585
R107 B.n388 B.n15 585
R108 B.n319 B.n14 585
R109 B.n389 B.n14 585
R110 B.n318 B.n13 585
R111 B.n390 B.n13 585
R112 B.n317 B.n316 585
R113 B.n316 B.n12 585
R114 B.n315 B.n314 585
R115 B.n315 B.n8 585
R116 B.n313 B.n7 585
R117 B.n397 B.n7 585
R118 B.n312 B.n6 585
R119 B.n398 B.n6 585
R120 B.n311 B.n5 585
R121 B.n399 B.n5 585
R122 B.n310 B.n309 585
R123 B.n309 B.n4 585
R124 B.n308 B.n118 585
R125 B.n308 B.n307 585
R126 B.n298 B.n119 585
R127 B.n120 B.n119 585
R128 B.n300 B.n299 585
R129 B.n301 B.n300 585
R130 B.n297 B.n124 585
R131 B.n128 B.n124 585
R132 B.n296 B.n295 585
R133 B.n295 B.n294 585
R134 B.n126 B.n125 585
R135 B.n127 B.n126 585
R136 B.n287 B.n286 585
R137 B.n288 B.n287 585
R138 B.n285 B.n133 585
R139 B.n133 B.n132 585
R140 B.n284 B.n283 585
R141 B.n283 B.n282 585
R142 B.n135 B.n134 585
R143 B.n136 B.n135 585
R144 B.n275 B.n274 585
R145 B.n276 B.n275 585
R146 B.n273 B.n141 585
R147 B.n141 B.n140 585
R148 B.n272 B.n271 585
R149 B.n271 B.n270 585
R150 B.n143 B.n142 585
R151 B.n144 B.n143 585
R152 B.n263 B.n262 585
R153 B.n264 B.n263 585
R154 B.n261 B.n149 585
R155 B.n149 B.n148 585
R156 B.n260 B.n259 585
R157 B.n259 B.n258 585
R158 B.n151 B.n150 585
R159 B.n152 B.n151 585
R160 B.n251 B.n250 585
R161 B.n252 B.n251 585
R162 B.n249 B.n157 585
R163 B.n157 B.n156 585
R164 B.n248 B.n247 585
R165 B.n247 B.n246 585
R166 B.n159 B.n158 585
R167 B.n160 B.n159 585
R168 B.n239 B.n238 585
R169 B.n240 B.n239 585
R170 B.n237 B.n165 585
R171 B.n165 B.n164 585
R172 B.n232 B.n231 585
R173 B.n230 B.n180 585
R174 B.n229 B.n179 585
R175 B.n234 B.n179 585
R176 B.n228 B.n227 585
R177 B.n226 B.n225 585
R178 B.n224 B.n223 585
R179 B.n222 B.n221 585
R180 B.n220 B.n219 585
R181 B.n217 B.n216 585
R182 B.n215 B.n214 585
R183 B.n213 B.n212 585
R184 B.n211 B.n210 585
R185 B.n209 B.n208 585
R186 B.n207 B.n206 585
R187 B.n205 B.n204 585
R188 B.n203 B.n202 585
R189 B.n201 B.n200 585
R190 B.n199 B.n198 585
R191 B.n196 B.n195 585
R192 B.n194 B.n193 585
R193 B.n192 B.n191 585
R194 B.n190 B.n189 585
R195 B.n188 B.n187 585
R196 B.n186 B.n185 585
R197 B.n167 B.n166 585
R198 B.n236 B.n235 585
R199 B.n235 B.n234 585
R200 B.n163 B.n162 585
R201 B.n164 B.n163 585
R202 B.n242 B.n241 585
R203 B.n241 B.n240 585
R204 B.n243 B.n161 585
R205 B.n161 B.n160 585
R206 B.n245 B.n244 585
R207 B.n246 B.n245 585
R208 B.n155 B.n154 585
R209 B.n156 B.n155 585
R210 B.n254 B.n253 585
R211 B.n253 B.n252 585
R212 B.n255 B.n153 585
R213 B.n153 B.n152 585
R214 B.n257 B.n256 585
R215 B.n258 B.n257 585
R216 B.n147 B.n146 585
R217 B.n148 B.n147 585
R218 B.n266 B.n265 585
R219 B.n265 B.n264 585
R220 B.n267 B.n145 585
R221 B.n145 B.n144 585
R222 B.n269 B.n268 585
R223 B.n270 B.n269 585
R224 B.n139 B.n138 585
R225 B.n140 B.n139 585
R226 B.n278 B.n277 585
R227 B.n277 B.n276 585
R228 B.n279 B.n137 585
R229 B.n137 B.n136 585
R230 B.n281 B.n280 585
R231 B.n282 B.n281 585
R232 B.n131 B.n130 585
R233 B.n132 B.n131 585
R234 B.n290 B.n289 585
R235 B.n289 B.n288 585
R236 B.n291 B.n129 585
R237 B.n129 B.n127 585
R238 B.n293 B.n292 585
R239 B.n294 B.n293 585
R240 B.n123 B.n122 585
R241 B.n128 B.n123 585
R242 B.n303 B.n302 585
R243 B.n302 B.n301 585
R244 B.n304 B.n121 585
R245 B.n121 B.n120 585
R246 B.n306 B.n305 585
R247 B.n307 B.n306 585
R248 B.n3 B.n0 585
R249 B.n4 B.n3 585
R250 B.n396 B.n1 585
R251 B.n397 B.n396 585
R252 B.n395 B.n394 585
R253 B.n395 B.n8 585
R254 B.n393 B.n9 585
R255 B.n12 B.n9 585
R256 B.n392 B.n391 585
R257 B.n391 B.n390 585
R258 B.n11 B.n10 585
R259 B.n389 B.n11 585
R260 B.n387 B.n386 585
R261 B.n388 B.n387 585
R262 B.n385 B.n17 585
R263 B.n17 B.n16 585
R264 B.n384 B.n383 585
R265 B.n383 B.n382 585
R266 B.n19 B.n18 585
R267 B.n381 B.n19 585
R268 B.n379 B.n378 585
R269 B.n380 B.n379 585
R270 B.n377 B.n24 585
R271 B.n24 B.n23 585
R272 B.n376 B.n375 585
R273 B.n375 B.n374 585
R274 B.n26 B.n25 585
R275 B.n373 B.n26 585
R276 B.n371 B.n370 585
R277 B.n372 B.n371 585
R278 B.n369 B.n31 585
R279 B.n31 B.n30 585
R280 B.n368 B.n367 585
R281 B.n367 B.n366 585
R282 B.n33 B.n32 585
R283 B.n365 B.n33 585
R284 B.n363 B.n362 585
R285 B.n364 B.n363 585
R286 B.n361 B.n38 585
R287 B.n38 B.n37 585
R288 B.n360 B.n359 585
R289 B.n359 B.n358 585
R290 B.n40 B.n39 585
R291 B.n357 B.n40 585
R292 B.n355 B.n354 585
R293 B.n356 B.n355 585
R294 B.n353 B.n45 585
R295 B.n45 B.n44 585
R296 B.n352 B.n351 585
R297 B.n351 B.n350 585
R298 B.n47 B.n46 585
R299 B.n349 B.n47 585
R300 B.n400 B.n399 585
R301 B.n398 B.n2 585
R302 B.n69 B.n47 516.524
R303 B.n346 B.n49 516.524
R304 B.n235 B.n165 516.524
R305 B.n232 B.n163 516.524
R306 B.n66 B.t13 278.488
R307 B.n63 B.t16 278.488
R308 B.n183 B.t10 278.488
R309 B.n181 B.t7 278.488
R310 B.n234 B.n164 264.45
R311 B.n349 B.n348 264.45
R312 B.n348 B.n347 256.663
R313 B.n348 B.n61 256.663
R314 B.n348 B.n60 256.663
R315 B.n348 B.n59 256.663
R316 B.n348 B.n58 256.663
R317 B.n348 B.n57 256.663
R318 B.n348 B.n56 256.663
R319 B.n348 B.n55 256.663
R320 B.n348 B.n54 256.663
R321 B.n348 B.n53 256.663
R322 B.n348 B.n52 256.663
R323 B.n348 B.n51 256.663
R324 B.n348 B.n50 256.663
R325 B.n234 B.n233 256.663
R326 B.n234 B.n168 256.663
R327 B.n234 B.n169 256.663
R328 B.n234 B.n170 256.663
R329 B.n234 B.n171 256.663
R330 B.n234 B.n172 256.663
R331 B.n234 B.n173 256.663
R332 B.n234 B.n174 256.663
R333 B.n234 B.n175 256.663
R334 B.n234 B.n176 256.663
R335 B.n234 B.n177 256.663
R336 B.n234 B.n178 256.663
R337 B.n402 B.n401 256.663
R338 B.n67 B.t14 239.7
R339 B.n64 B.t17 239.7
R340 B.n184 B.t9 239.7
R341 B.n182 B.t6 239.7
R342 B.n66 B.t11 207.919
R343 B.n63 B.t15 207.919
R344 B.n183 B.t8 207.919
R345 B.n181 B.t4 207.919
R346 B.n73 B.n72 163.367
R347 B.n77 B.n76 163.367
R348 B.n81 B.n80 163.367
R349 B.n85 B.n84 163.367
R350 B.n89 B.n88 163.367
R351 B.n93 B.n92 163.367
R352 B.n97 B.n96 163.367
R353 B.n101 B.n100 163.367
R354 B.n105 B.n104 163.367
R355 B.n109 B.n108 163.367
R356 B.n113 B.n112 163.367
R357 B.n115 B.n62 163.367
R358 B.n239 B.n165 163.367
R359 B.n239 B.n159 163.367
R360 B.n247 B.n159 163.367
R361 B.n247 B.n157 163.367
R362 B.n251 B.n157 163.367
R363 B.n251 B.n151 163.367
R364 B.n259 B.n151 163.367
R365 B.n259 B.n149 163.367
R366 B.n263 B.n149 163.367
R367 B.n263 B.n143 163.367
R368 B.n271 B.n143 163.367
R369 B.n271 B.n141 163.367
R370 B.n275 B.n141 163.367
R371 B.n275 B.n135 163.367
R372 B.n283 B.n135 163.367
R373 B.n283 B.n133 163.367
R374 B.n287 B.n133 163.367
R375 B.n287 B.n126 163.367
R376 B.n295 B.n126 163.367
R377 B.n295 B.n124 163.367
R378 B.n300 B.n124 163.367
R379 B.n300 B.n119 163.367
R380 B.n308 B.n119 163.367
R381 B.n309 B.n308 163.367
R382 B.n309 B.n5 163.367
R383 B.n6 B.n5 163.367
R384 B.n7 B.n6 163.367
R385 B.n315 B.n7 163.367
R386 B.n316 B.n315 163.367
R387 B.n316 B.n13 163.367
R388 B.n14 B.n13 163.367
R389 B.n15 B.n14 163.367
R390 B.n321 B.n15 163.367
R391 B.n321 B.n20 163.367
R392 B.n21 B.n20 163.367
R393 B.n22 B.n21 163.367
R394 B.n326 B.n22 163.367
R395 B.n326 B.n27 163.367
R396 B.n28 B.n27 163.367
R397 B.n29 B.n28 163.367
R398 B.n331 B.n29 163.367
R399 B.n331 B.n34 163.367
R400 B.n35 B.n34 163.367
R401 B.n36 B.n35 163.367
R402 B.n336 B.n36 163.367
R403 B.n336 B.n41 163.367
R404 B.n42 B.n41 163.367
R405 B.n43 B.n42 163.367
R406 B.n341 B.n43 163.367
R407 B.n341 B.n48 163.367
R408 B.n49 B.n48 163.367
R409 B.n180 B.n179 163.367
R410 B.n227 B.n179 163.367
R411 B.n225 B.n224 163.367
R412 B.n221 B.n220 163.367
R413 B.n216 B.n215 163.367
R414 B.n212 B.n211 163.367
R415 B.n208 B.n207 163.367
R416 B.n204 B.n203 163.367
R417 B.n200 B.n199 163.367
R418 B.n195 B.n194 163.367
R419 B.n191 B.n190 163.367
R420 B.n187 B.n186 163.367
R421 B.n235 B.n167 163.367
R422 B.n241 B.n163 163.367
R423 B.n241 B.n161 163.367
R424 B.n245 B.n161 163.367
R425 B.n245 B.n155 163.367
R426 B.n253 B.n155 163.367
R427 B.n253 B.n153 163.367
R428 B.n257 B.n153 163.367
R429 B.n257 B.n147 163.367
R430 B.n265 B.n147 163.367
R431 B.n265 B.n145 163.367
R432 B.n269 B.n145 163.367
R433 B.n269 B.n139 163.367
R434 B.n277 B.n139 163.367
R435 B.n277 B.n137 163.367
R436 B.n281 B.n137 163.367
R437 B.n281 B.n131 163.367
R438 B.n289 B.n131 163.367
R439 B.n289 B.n129 163.367
R440 B.n293 B.n129 163.367
R441 B.n293 B.n123 163.367
R442 B.n302 B.n123 163.367
R443 B.n302 B.n121 163.367
R444 B.n306 B.n121 163.367
R445 B.n306 B.n3 163.367
R446 B.n400 B.n3 163.367
R447 B.n396 B.n2 163.367
R448 B.n396 B.n395 163.367
R449 B.n395 B.n9 163.367
R450 B.n391 B.n9 163.367
R451 B.n391 B.n11 163.367
R452 B.n387 B.n11 163.367
R453 B.n387 B.n17 163.367
R454 B.n383 B.n17 163.367
R455 B.n383 B.n19 163.367
R456 B.n379 B.n19 163.367
R457 B.n379 B.n24 163.367
R458 B.n375 B.n24 163.367
R459 B.n375 B.n26 163.367
R460 B.n371 B.n26 163.367
R461 B.n371 B.n31 163.367
R462 B.n367 B.n31 163.367
R463 B.n367 B.n33 163.367
R464 B.n363 B.n33 163.367
R465 B.n363 B.n38 163.367
R466 B.n359 B.n38 163.367
R467 B.n359 B.n40 163.367
R468 B.n355 B.n40 163.367
R469 B.n355 B.n45 163.367
R470 B.n351 B.n45 163.367
R471 B.n351 B.n47 163.367
R472 B.n240 B.n164 127.537
R473 B.n240 B.n160 127.537
R474 B.n246 B.n160 127.537
R475 B.n246 B.n156 127.537
R476 B.n252 B.n156 127.537
R477 B.n258 B.n152 127.537
R478 B.n258 B.n148 127.537
R479 B.n264 B.n148 127.537
R480 B.n264 B.n144 127.537
R481 B.n270 B.n144 127.537
R482 B.n270 B.n140 127.537
R483 B.n276 B.n140 127.537
R484 B.n276 B.n136 127.537
R485 B.n282 B.n136 127.537
R486 B.n288 B.n132 127.537
R487 B.n288 B.n127 127.537
R488 B.n294 B.n127 127.537
R489 B.n294 B.n128 127.537
R490 B.n301 B.n120 127.537
R491 B.n307 B.n120 127.537
R492 B.n307 B.n4 127.537
R493 B.n399 B.n4 127.537
R494 B.n399 B.n398 127.537
R495 B.n398 B.n397 127.537
R496 B.n397 B.n8 127.537
R497 B.n12 B.n8 127.537
R498 B.n390 B.n12 127.537
R499 B.n389 B.n388 127.537
R500 B.n388 B.n16 127.537
R501 B.n382 B.n16 127.537
R502 B.n382 B.n381 127.537
R503 B.n380 B.n23 127.537
R504 B.n374 B.n23 127.537
R505 B.n374 B.n373 127.537
R506 B.n373 B.n372 127.537
R507 B.n372 B.n30 127.537
R508 B.n366 B.n30 127.537
R509 B.n366 B.n365 127.537
R510 B.n365 B.n364 127.537
R511 B.n364 B.n37 127.537
R512 B.n358 B.n357 127.537
R513 B.n357 B.n356 127.537
R514 B.n356 B.n44 127.537
R515 B.n350 B.n44 127.537
R516 B.n350 B.n349 127.537
R517 B.n252 B.t5 125.662
R518 B.n358 B.t12 125.662
R519 B.n128 B.t1 121.91
R520 B.t0 B.n389 121.91
R521 B.t3 B.n132 118.159
R522 B.n381 B.t2 118.159
R523 B.n69 B.n50 71.676
R524 B.n73 B.n51 71.676
R525 B.n77 B.n52 71.676
R526 B.n81 B.n53 71.676
R527 B.n85 B.n54 71.676
R528 B.n89 B.n55 71.676
R529 B.n93 B.n56 71.676
R530 B.n97 B.n57 71.676
R531 B.n101 B.n58 71.676
R532 B.n105 B.n59 71.676
R533 B.n109 B.n60 71.676
R534 B.n113 B.n61 71.676
R535 B.n347 B.n62 71.676
R536 B.n347 B.n346 71.676
R537 B.n115 B.n61 71.676
R538 B.n112 B.n60 71.676
R539 B.n108 B.n59 71.676
R540 B.n104 B.n58 71.676
R541 B.n100 B.n57 71.676
R542 B.n96 B.n56 71.676
R543 B.n92 B.n55 71.676
R544 B.n88 B.n54 71.676
R545 B.n84 B.n53 71.676
R546 B.n80 B.n52 71.676
R547 B.n76 B.n51 71.676
R548 B.n72 B.n50 71.676
R549 B.n233 B.n232 71.676
R550 B.n227 B.n168 71.676
R551 B.n224 B.n169 71.676
R552 B.n220 B.n170 71.676
R553 B.n215 B.n171 71.676
R554 B.n211 B.n172 71.676
R555 B.n207 B.n173 71.676
R556 B.n203 B.n174 71.676
R557 B.n199 B.n175 71.676
R558 B.n194 B.n176 71.676
R559 B.n190 B.n177 71.676
R560 B.n186 B.n178 71.676
R561 B.n233 B.n180 71.676
R562 B.n225 B.n168 71.676
R563 B.n221 B.n169 71.676
R564 B.n216 B.n170 71.676
R565 B.n212 B.n171 71.676
R566 B.n208 B.n172 71.676
R567 B.n204 B.n173 71.676
R568 B.n200 B.n174 71.676
R569 B.n195 B.n175 71.676
R570 B.n191 B.n176 71.676
R571 B.n187 B.n177 71.676
R572 B.n178 B.n167 71.676
R573 B.n401 B.n400 71.676
R574 B.n401 B.n2 71.676
R575 B.n68 B.n67 59.5399
R576 B.n65 B.n64 59.5399
R577 B.n197 B.n184 59.5399
R578 B.n218 B.n182 59.5399
R579 B.n67 B.n66 38.7884
R580 B.n64 B.n63 38.7884
R581 B.n184 B.n183 38.7884
R582 B.n182 B.n181 38.7884
R583 B.n231 B.n162 33.5615
R584 B.n237 B.n236 33.5615
R585 B.n345 B.n344 33.5615
R586 B.n70 B.n46 33.5615
R587 B B.n402 18.0485
R588 B.n242 B.n162 10.6151
R589 B.n243 B.n242 10.6151
R590 B.n244 B.n243 10.6151
R591 B.n244 B.n154 10.6151
R592 B.n254 B.n154 10.6151
R593 B.n255 B.n254 10.6151
R594 B.n256 B.n255 10.6151
R595 B.n256 B.n146 10.6151
R596 B.n266 B.n146 10.6151
R597 B.n267 B.n266 10.6151
R598 B.n268 B.n267 10.6151
R599 B.n268 B.n138 10.6151
R600 B.n278 B.n138 10.6151
R601 B.n279 B.n278 10.6151
R602 B.n280 B.n279 10.6151
R603 B.n280 B.n130 10.6151
R604 B.n290 B.n130 10.6151
R605 B.n291 B.n290 10.6151
R606 B.n292 B.n291 10.6151
R607 B.n292 B.n122 10.6151
R608 B.n303 B.n122 10.6151
R609 B.n304 B.n303 10.6151
R610 B.n305 B.n304 10.6151
R611 B.n305 B.n0 10.6151
R612 B.n231 B.n230 10.6151
R613 B.n230 B.n229 10.6151
R614 B.n229 B.n228 10.6151
R615 B.n228 B.n226 10.6151
R616 B.n226 B.n223 10.6151
R617 B.n223 B.n222 10.6151
R618 B.n222 B.n219 10.6151
R619 B.n217 B.n214 10.6151
R620 B.n214 B.n213 10.6151
R621 B.n213 B.n210 10.6151
R622 B.n210 B.n209 10.6151
R623 B.n209 B.n206 10.6151
R624 B.n206 B.n205 10.6151
R625 B.n205 B.n202 10.6151
R626 B.n202 B.n201 10.6151
R627 B.n201 B.n198 10.6151
R628 B.n196 B.n193 10.6151
R629 B.n193 B.n192 10.6151
R630 B.n192 B.n189 10.6151
R631 B.n189 B.n188 10.6151
R632 B.n188 B.n185 10.6151
R633 B.n185 B.n166 10.6151
R634 B.n236 B.n166 10.6151
R635 B.n238 B.n237 10.6151
R636 B.n238 B.n158 10.6151
R637 B.n248 B.n158 10.6151
R638 B.n249 B.n248 10.6151
R639 B.n250 B.n249 10.6151
R640 B.n250 B.n150 10.6151
R641 B.n260 B.n150 10.6151
R642 B.n261 B.n260 10.6151
R643 B.n262 B.n261 10.6151
R644 B.n262 B.n142 10.6151
R645 B.n272 B.n142 10.6151
R646 B.n273 B.n272 10.6151
R647 B.n274 B.n273 10.6151
R648 B.n274 B.n134 10.6151
R649 B.n284 B.n134 10.6151
R650 B.n285 B.n284 10.6151
R651 B.n286 B.n285 10.6151
R652 B.n286 B.n125 10.6151
R653 B.n296 B.n125 10.6151
R654 B.n297 B.n296 10.6151
R655 B.n299 B.n297 10.6151
R656 B.n299 B.n298 10.6151
R657 B.n298 B.n118 10.6151
R658 B.n310 B.n118 10.6151
R659 B.n311 B.n310 10.6151
R660 B.n312 B.n311 10.6151
R661 B.n313 B.n312 10.6151
R662 B.n314 B.n313 10.6151
R663 B.n317 B.n314 10.6151
R664 B.n318 B.n317 10.6151
R665 B.n319 B.n318 10.6151
R666 B.n320 B.n319 10.6151
R667 B.n322 B.n320 10.6151
R668 B.n323 B.n322 10.6151
R669 B.n324 B.n323 10.6151
R670 B.n325 B.n324 10.6151
R671 B.n327 B.n325 10.6151
R672 B.n328 B.n327 10.6151
R673 B.n329 B.n328 10.6151
R674 B.n330 B.n329 10.6151
R675 B.n332 B.n330 10.6151
R676 B.n333 B.n332 10.6151
R677 B.n334 B.n333 10.6151
R678 B.n335 B.n334 10.6151
R679 B.n337 B.n335 10.6151
R680 B.n338 B.n337 10.6151
R681 B.n339 B.n338 10.6151
R682 B.n340 B.n339 10.6151
R683 B.n342 B.n340 10.6151
R684 B.n343 B.n342 10.6151
R685 B.n344 B.n343 10.6151
R686 B.n394 B.n1 10.6151
R687 B.n394 B.n393 10.6151
R688 B.n393 B.n392 10.6151
R689 B.n392 B.n10 10.6151
R690 B.n386 B.n10 10.6151
R691 B.n386 B.n385 10.6151
R692 B.n385 B.n384 10.6151
R693 B.n384 B.n18 10.6151
R694 B.n378 B.n18 10.6151
R695 B.n378 B.n377 10.6151
R696 B.n377 B.n376 10.6151
R697 B.n376 B.n25 10.6151
R698 B.n370 B.n25 10.6151
R699 B.n370 B.n369 10.6151
R700 B.n369 B.n368 10.6151
R701 B.n368 B.n32 10.6151
R702 B.n362 B.n32 10.6151
R703 B.n362 B.n361 10.6151
R704 B.n361 B.n360 10.6151
R705 B.n360 B.n39 10.6151
R706 B.n354 B.n39 10.6151
R707 B.n354 B.n353 10.6151
R708 B.n353 B.n352 10.6151
R709 B.n352 B.n46 10.6151
R710 B.n71 B.n70 10.6151
R711 B.n74 B.n71 10.6151
R712 B.n75 B.n74 10.6151
R713 B.n78 B.n75 10.6151
R714 B.n79 B.n78 10.6151
R715 B.n82 B.n79 10.6151
R716 B.n83 B.n82 10.6151
R717 B.n87 B.n86 10.6151
R718 B.n90 B.n87 10.6151
R719 B.n91 B.n90 10.6151
R720 B.n94 B.n91 10.6151
R721 B.n95 B.n94 10.6151
R722 B.n98 B.n95 10.6151
R723 B.n99 B.n98 10.6151
R724 B.n102 B.n99 10.6151
R725 B.n103 B.n102 10.6151
R726 B.n107 B.n106 10.6151
R727 B.n110 B.n107 10.6151
R728 B.n111 B.n110 10.6151
R729 B.n114 B.n111 10.6151
R730 B.n116 B.n114 10.6151
R731 B.n117 B.n116 10.6151
R732 B.n345 B.n117 10.6151
R733 B.n282 B.t3 9.37816
R734 B.t2 B.n380 9.37816
R735 B.n219 B.n218 9.36635
R736 B.n197 B.n196 9.36635
R737 B.n83 B.n68 9.36635
R738 B.n106 B.n65 9.36635
R739 B.n402 B.n0 8.11757
R740 B.n402 B.n1 8.11757
R741 B.n301 B.t1 5.6271
R742 B.n390 B.t0 5.6271
R743 B.t5 B.n152 1.87603
R744 B.t12 B.n37 1.87603
R745 B.n218 B.n217 1.24928
R746 B.n198 B.n197 1.24928
R747 B.n86 B.n68 1.24928
R748 B.n103 B.n65 1.24928
R749 VN VN.n1 44.6488
R750 VN.n0 VN.t2 43.0851
R751 VN.n1 VN.t1 43.0851
R752 VN.n0 VN.t3 42.6674
R753 VN.n1 VN.t0 42.6674
R754 VN VN.n0 9.63747
R755 VDD2.n2 VDD2.n0 263.065
R756 VDD2.n2 VDD2.n1 233.671
R757 VDD2.n1 VDD2.t3 33.5598
R758 VDD2.n1 VDD2.t2 33.5598
R759 VDD2.n0 VDD2.t1 33.5598
R760 VDD2.n0 VDD2.t0 33.5598
R761 VDD2 VDD2.n2 0.0586897
C0 VDD1 VTAIL 2.18345f
C1 VDD1 VP 0.703551f
C2 VDD1 VDD2 0.799994f
C3 VDD1 VN 0.155694f
C4 VTAIL VP 1.045f
C5 VTAIL VDD2 2.23142f
C6 VTAIL VN 1.03089f
C7 VDD2 VP 0.344224f
C8 VN VP 3.42133f
C9 VN VDD2 0.51724f
C10 VDD2 B 2.32444f
C11 VDD1 B 4.43362f
C12 VTAIL B 2.408174f
C13 VN B 7.50167f
C14 VP B 5.955934f
C15 VDD2.t1 B 0.011399f
C16 VDD2.t0 B 0.011399f
C17 VDD2.n0 B 0.10367f
C18 VDD2.t3 B 0.011399f
C19 VDD2.t2 B 0.011399f
C20 VDD2.n1 B 0.029192f
C21 VDD2.n2 B 1.88045f
C22 VN.t2 B 0.200571f
C23 VN.t3 B 0.198774f
C24 VN.n0 B 0.131357f
C25 VN.t1 B 0.200571f
C26 VN.t0 B 0.198774f
C27 VN.n1 B 1.03553f
C28 VDD1.t0 B 0.010949f
C29 VDD1.t1 B 0.010949f
C30 VDD1.n0 B 0.028091f
C31 VDD1.t2 B 0.010949f
C32 VDD1.t3 B 0.010949f
C33 VDD1.n1 B 0.106184f
C34 VTAIL.t0 B 0.055317f
C35 VTAIL.n0 B 0.163811f
C36 VTAIL.t2 B 0.055317f
C37 VTAIL.n1 B 0.233932f
C38 VTAIL.t3 B 0.055317f
C39 VTAIL.n2 B 0.755435f
C40 VTAIL.t7 B 0.055317f
C41 VTAIL.n3 B 0.755435f
C42 VTAIL.t1 B 0.055317f
C43 VTAIL.n4 B 0.233932f
C44 VTAIL.t5 B 0.055317f
C45 VTAIL.n5 B 0.233932f
C46 VTAIL.t4 B 0.055317f
C47 VTAIL.n6 B 0.755435f
C48 VTAIL.t6 B 0.055317f
C49 VTAIL.n7 B 0.675162f
C50 VP.n0 B 0.042283f
C51 VP.t0 B 0.038525f
C52 VP.n1 B 0.063742f
C53 VP.t2 B 0.20141f
C54 VP.t3 B 0.20323f
C55 VP.n2 B 1.03321f
C56 VP.t1 B 0.038525f
C57 VP.n3 B 0.149906f
C58 VP.n4 B 1.24875f
C59 VP.n5 B 0.042283f
C60 VP.n6 B 0.032072f
C61 VP.n7 B 0.025927f
C62 VP.n8 B 0.063742f
C63 VP.n9 B 0.149906f
C64 VP.n10 B 0.033243f
.ends

