// Decoder output to apply to DCO
//

module decode_dco(
    input prop_gain,
    output dc_swval,
    input freq_val,

);

endmodule : decode_dco
