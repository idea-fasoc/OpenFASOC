* NGSPICE file created from diff_pair_sample_0129.ext - technology: sky130A

.subckt diff_pair_sample_0129 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t2 w_n3130_n3088# sky130_fd_pr__pfet_01v8 ad=1.749 pd=10.93 as=1.749 ps=10.93 w=10.6 l=1.83
X1 VDD2.t7 VN.t0 VTAIL.t3 w_n3130_n3088# sky130_fd_pr__pfet_01v8 ad=1.749 pd=10.93 as=1.749 ps=10.93 w=10.6 l=1.83
X2 B.t11 B.t9 B.t10 w_n3130_n3088# sky130_fd_pr__pfet_01v8 ad=4.134 pd=21.98 as=0 ps=0 w=10.6 l=1.83
X3 VTAIL.t1 VN.t1 VDD2.t6 w_n3130_n3088# sky130_fd_pr__pfet_01v8 ad=1.749 pd=10.93 as=1.749 ps=10.93 w=10.6 l=1.83
X4 VTAIL.t14 VP.t1 VDD1.t1 w_n3130_n3088# sky130_fd_pr__pfet_01v8 ad=4.134 pd=21.98 as=1.749 ps=10.93 w=10.6 l=1.83
X5 VDD2.t5 VN.t2 VTAIL.t4 w_n3130_n3088# sky130_fd_pr__pfet_01v8 ad=1.749 pd=10.93 as=4.134 ps=21.98 w=10.6 l=1.83
X6 VDD1.t0 VP.t2 VTAIL.t13 w_n3130_n3088# sky130_fd_pr__pfet_01v8 ad=1.749 pd=10.93 as=1.749 ps=10.93 w=10.6 l=1.83
X7 VDD1.t4 VP.t3 VTAIL.t12 w_n3130_n3088# sky130_fd_pr__pfet_01v8 ad=1.749 pd=10.93 as=4.134 ps=21.98 w=10.6 l=1.83
X8 VDD2.t4 VN.t3 VTAIL.t5 w_n3130_n3088# sky130_fd_pr__pfet_01v8 ad=1.749 pd=10.93 as=1.749 ps=10.93 w=10.6 l=1.83
X9 VDD1.t3 VP.t4 VTAIL.t11 w_n3130_n3088# sky130_fd_pr__pfet_01v8 ad=1.749 pd=10.93 as=1.749 ps=10.93 w=10.6 l=1.83
X10 B.t8 B.t6 B.t7 w_n3130_n3088# sky130_fd_pr__pfet_01v8 ad=4.134 pd=21.98 as=0 ps=0 w=10.6 l=1.83
X11 VDD1.t7 VP.t5 VTAIL.t10 w_n3130_n3088# sky130_fd_pr__pfet_01v8 ad=1.749 pd=10.93 as=4.134 ps=21.98 w=10.6 l=1.83
X12 VTAIL.t6 VN.t4 VDD2.t3 w_n3130_n3088# sky130_fd_pr__pfet_01v8 ad=1.749 pd=10.93 as=1.749 ps=10.93 w=10.6 l=1.83
X13 VDD2.t2 VN.t5 VTAIL.t0 w_n3130_n3088# sky130_fd_pr__pfet_01v8 ad=1.749 pd=10.93 as=4.134 ps=21.98 w=10.6 l=1.83
X14 VTAIL.t9 VP.t6 VDD1.t6 w_n3130_n3088# sky130_fd_pr__pfet_01v8 ad=4.134 pd=21.98 as=1.749 ps=10.93 w=10.6 l=1.83
X15 VTAIL.t7 VN.t6 VDD2.t1 w_n3130_n3088# sky130_fd_pr__pfet_01v8 ad=4.134 pd=21.98 as=1.749 ps=10.93 w=10.6 l=1.83
X16 VTAIL.t8 VP.t7 VDD1.t5 w_n3130_n3088# sky130_fd_pr__pfet_01v8 ad=1.749 pd=10.93 as=1.749 ps=10.93 w=10.6 l=1.83
X17 VTAIL.t2 VN.t7 VDD2.t0 w_n3130_n3088# sky130_fd_pr__pfet_01v8 ad=4.134 pd=21.98 as=1.749 ps=10.93 w=10.6 l=1.83
X18 B.t5 B.t3 B.t4 w_n3130_n3088# sky130_fd_pr__pfet_01v8 ad=4.134 pd=21.98 as=0 ps=0 w=10.6 l=1.83
X19 B.t2 B.t0 B.t1 w_n3130_n3088# sky130_fd_pr__pfet_01v8 ad=4.134 pd=21.98 as=0 ps=0 w=10.6 l=1.83
R0 VP.n10 VP.t1 171.28
R1 VP.n13 VP.n12 161.3
R2 VP.n14 VP.n9 161.3
R3 VP.n16 VP.n15 161.3
R4 VP.n17 VP.n8 161.3
R5 VP.n20 VP.n19 161.3
R6 VP.n21 VP.n7 161.3
R7 VP.n23 VP.n22 161.3
R8 VP.n24 VP.n6 161.3
R9 VP.n48 VP.n0 161.3
R10 VP.n47 VP.n46 161.3
R11 VP.n45 VP.n1 161.3
R12 VP.n44 VP.n43 161.3
R13 VP.n41 VP.n2 161.3
R14 VP.n40 VP.n39 161.3
R15 VP.n38 VP.n3 161.3
R16 VP.n37 VP.n36 161.3
R17 VP.n34 VP.n4 161.3
R18 VP.n33 VP.n32 161.3
R19 VP.n31 VP.n5 161.3
R20 VP.n30 VP.n29 161.3
R21 VP.n28 VP.t6 139.596
R22 VP.n35 VP.t2 139.596
R23 VP.n42 VP.t0 139.596
R24 VP.n49 VP.t5 139.596
R25 VP.n25 VP.t3 139.596
R26 VP.n18 VP.t7 139.596
R27 VP.n11 VP.t4 139.596
R28 VP.n28 VP.n27 86.8082
R29 VP.n50 VP.n49 86.8082
R30 VP.n26 VP.n25 86.8082
R31 VP.n40 VP.n3 56.5617
R32 VP.n16 VP.n9 56.5617
R33 VP.n11 VP.n10 53.8128
R34 VP.n33 VP.n5 49.296
R35 VP.n47 VP.n1 49.296
R36 VP.n23 VP.n7 49.296
R37 VP.n27 VP.n26 46.28
R38 VP.n29 VP.n5 31.8581
R39 VP.n48 VP.n47 31.8581
R40 VP.n24 VP.n23 31.8581
R41 VP.n34 VP.n33 24.5923
R42 VP.n36 VP.n3 24.5923
R43 VP.n41 VP.n40 24.5923
R44 VP.n43 VP.n1 24.5923
R45 VP.n17 VP.n16 24.5923
R46 VP.n19 VP.n7 24.5923
R47 VP.n12 VP.n9 24.5923
R48 VP.n29 VP.n28 24.1005
R49 VP.n49 VP.n48 24.1005
R50 VP.n25 VP.n24 24.1005
R51 VP.n36 VP.n35 16.2311
R52 VP.n42 VP.n41 16.2311
R53 VP.n18 VP.n17 16.2311
R54 VP.n12 VP.n11 16.2311
R55 VP.n13 VP.n10 12.6399
R56 VP.n35 VP.n34 8.36172
R57 VP.n43 VP.n42 8.36172
R58 VP.n19 VP.n18 8.36172
R59 VP.n26 VP.n6 0.278335
R60 VP.n30 VP.n27 0.278335
R61 VP.n50 VP.n0 0.278335
R62 VP.n14 VP.n13 0.189894
R63 VP.n15 VP.n14 0.189894
R64 VP.n15 VP.n8 0.189894
R65 VP.n20 VP.n8 0.189894
R66 VP.n21 VP.n20 0.189894
R67 VP.n22 VP.n21 0.189894
R68 VP.n22 VP.n6 0.189894
R69 VP.n31 VP.n30 0.189894
R70 VP.n32 VP.n31 0.189894
R71 VP.n32 VP.n4 0.189894
R72 VP.n37 VP.n4 0.189894
R73 VP.n38 VP.n37 0.189894
R74 VP.n39 VP.n38 0.189894
R75 VP.n39 VP.n2 0.189894
R76 VP.n44 VP.n2 0.189894
R77 VP.n45 VP.n44 0.189894
R78 VP.n46 VP.n45 0.189894
R79 VP.n46 VP.n0 0.189894
R80 VP VP.n50 0.153485
R81 VDD1 VDD1.n0 75.3039
R82 VDD1.n3 VDD1.n2 75.1902
R83 VDD1.n3 VDD1.n1 75.1902
R84 VDD1.n5 VDD1.n4 74.3145
R85 VDD1.n5 VDD1.n3 41.8156
R86 VDD1.n4 VDD1.t5 3.06701
R87 VDD1.n4 VDD1.t4 3.06701
R88 VDD1.n0 VDD1.t1 3.06701
R89 VDD1.n0 VDD1.t3 3.06701
R90 VDD1.n2 VDD1.t2 3.06701
R91 VDD1.n2 VDD1.t7 3.06701
R92 VDD1.n1 VDD1.t6 3.06701
R93 VDD1.n1 VDD1.t0 3.06701
R94 VDD1 VDD1.n5 0.873345
R95 VTAIL.n466 VTAIL.n414 756.745
R96 VTAIL.n54 VTAIL.n2 756.745
R97 VTAIL.n112 VTAIL.n60 756.745
R98 VTAIL.n172 VTAIL.n120 756.745
R99 VTAIL.n408 VTAIL.n356 756.745
R100 VTAIL.n348 VTAIL.n296 756.745
R101 VTAIL.n290 VTAIL.n238 756.745
R102 VTAIL.n230 VTAIL.n178 756.745
R103 VTAIL.n433 VTAIL.n432 585
R104 VTAIL.n430 VTAIL.n429 585
R105 VTAIL.n439 VTAIL.n438 585
R106 VTAIL.n441 VTAIL.n440 585
R107 VTAIL.n426 VTAIL.n425 585
R108 VTAIL.n447 VTAIL.n446 585
R109 VTAIL.n450 VTAIL.n449 585
R110 VTAIL.n448 VTAIL.n422 585
R111 VTAIL.n455 VTAIL.n421 585
R112 VTAIL.n457 VTAIL.n456 585
R113 VTAIL.n459 VTAIL.n458 585
R114 VTAIL.n418 VTAIL.n417 585
R115 VTAIL.n465 VTAIL.n464 585
R116 VTAIL.n467 VTAIL.n466 585
R117 VTAIL.n21 VTAIL.n20 585
R118 VTAIL.n18 VTAIL.n17 585
R119 VTAIL.n27 VTAIL.n26 585
R120 VTAIL.n29 VTAIL.n28 585
R121 VTAIL.n14 VTAIL.n13 585
R122 VTAIL.n35 VTAIL.n34 585
R123 VTAIL.n38 VTAIL.n37 585
R124 VTAIL.n36 VTAIL.n10 585
R125 VTAIL.n43 VTAIL.n9 585
R126 VTAIL.n45 VTAIL.n44 585
R127 VTAIL.n47 VTAIL.n46 585
R128 VTAIL.n6 VTAIL.n5 585
R129 VTAIL.n53 VTAIL.n52 585
R130 VTAIL.n55 VTAIL.n54 585
R131 VTAIL.n79 VTAIL.n78 585
R132 VTAIL.n76 VTAIL.n75 585
R133 VTAIL.n85 VTAIL.n84 585
R134 VTAIL.n87 VTAIL.n86 585
R135 VTAIL.n72 VTAIL.n71 585
R136 VTAIL.n93 VTAIL.n92 585
R137 VTAIL.n96 VTAIL.n95 585
R138 VTAIL.n94 VTAIL.n68 585
R139 VTAIL.n101 VTAIL.n67 585
R140 VTAIL.n103 VTAIL.n102 585
R141 VTAIL.n105 VTAIL.n104 585
R142 VTAIL.n64 VTAIL.n63 585
R143 VTAIL.n111 VTAIL.n110 585
R144 VTAIL.n113 VTAIL.n112 585
R145 VTAIL.n139 VTAIL.n138 585
R146 VTAIL.n136 VTAIL.n135 585
R147 VTAIL.n145 VTAIL.n144 585
R148 VTAIL.n147 VTAIL.n146 585
R149 VTAIL.n132 VTAIL.n131 585
R150 VTAIL.n153 VTAIL.n152 585
R151 VTAIL.n156 VTAIL.n155 585
R152 VTAIL.n154 VTAIL.n128 585
R153 VTAIL.n161 VTAIL.n127 585
R154 VTAIL.n163 VTAIL.n162 585
R155 VTAIL.n165 VTAIL.n164 585
R156 VTAIL.n124 VTAIL.n123 585
R157 VTAIL.n171 VTAIL.n170 585
R158 VTAIL.n173 VTAIL.n172 585
R159 VTAIL.n409 VTAIL.n408 585
R160 VTAIL.n407 VTAIL.n406 585
R161 VTAIL.n360 VTAIL.n359 585
R162 VTAIL.n401 VTAIL.n400 585
R163 VTAIL.n399 VTAIL.n398 585
R164 VTAIL.n397 VTAIL.n363 585
R165 VTAIL.n367 VTAIL.n364 585
R166 VTAIL.n392 VTAIL.n391 585
R167 VTAIL.n390 VTAIL.n389 585
R168 VTAIL.n369 VTAIL.n368 585
R169 VTAIL.n384 VTAIL.n383 585
R170 VTAIL.n382 VTAIL.n381 585
R171 VTAIL.n373 VTAIL.n372 585
R172 VTAIL.n376 VTAIL.n375 585
R173 VTAIL.n349 VTAIL.n348 585
R174 VTAIL.n347 VTAIL.n346 585
R175 VTAIL.n300 VTAIL.n299 585
R176 VTAIL.n341 VTAIL.n340 585
R177 VTAIL.n339 VTAIL.n338 585
R178 VTAIL.n337 VTAIL.n303 585
R179 VTAIL.n307 VTAIL.n304 585
R180 VTAIL.n332 VTAIL.n331 585
R181 VTAIL.n330 VTAIL.n329 585
R182 VTAIL.n309 VTAIL.n308 585
R183 VTAIL.n324 VTAIL.n323 585
R184 VTAIL.n322 VTAIL.n321 585
R185 VTAIL.n313 VTAIL.n312 585
R186 VTAIL.n316 VTAIL.n315 585
R187 VTAIL.n291 VTAIL.n290 585
R188 VTAIL.n289 VTAIL.n288 585
R189 VTAIL.n242 VTAIL.n241 585
R190 VTAIL.n283 VTAIL.n282 585
R191 VTAIL.n281 VTAIL.n280 585
R192 VTAIL.n279 VTAIL.n245 585
R193 VTAIL.n249 VTAIL.n246 585
R194 VTAIL.n274 VTAIL.n273 585
R195 VTAIL.n272 VTAIL.n271 585
R196 VTAIL.n251 VTAIL.n250 585
R197 VTAIL.n266 VTAIL.n265 585
R198 VTAIL.n264 VTAIL.n263 585
R199 VTAIL.n255 VTAIL.n254 585
R200 VTAIL.n258 VTAIL.n257 585
R201 VTAIL.n231 VTAIL.n230 585
R202 VTAIL.n229 VTAIL.n228 585
R203 VTAIL.n182 VTAIL.n181 585
R204 VTAIL.n223 VTAIL.n222 585
R205 VTAIL.n221 VTAIL.n220 585
R206 VTAIL.n219 VTAIL.n185 585
R207 VTAIL.n189 VTAIL.n186 585
R208 VTAIL.n214 VTAIL.n213 585
R209 VTAIL.n212 VTAIL.n211 585
R210 VTAIL.n191 VTAIL.n190 585
R211 VTAIL.n206 VTAIL.n205 585
R212 VTAIL.n204 VTAIL.n203 585
R213 VTAIL.n195 VTAIL.n194 585
R214 VTAIL.n198 VTAIL.n197 585
R215 VTAIL.t12 VTAIL.n374 329.038
R216 VTAIL.t14 VTAIL.n314 329.038
R217 VTAIL.t4 VTAIL.n256 329.038
R218 VTAIL.t2 VTAIL.n196 329.038
R219 VTAIL.t0 VTAIL.n431 329.038
R220 VTAIL.t7 VTAIL.n19 329.038
R221 VTAIL.t10 VTAIL.n77 329.038
R222 VTAIL.t9 VTAIL.n137 329.038
R223 VTAIL.n432 VTAIL.n429 171.744
R224 VTAIL.n439 VTAIL.n429 171.744
R225 VTAIL.n440 VTAIL.n439 171.744
R226 VTAIL.n440 VTAIL.n425 171.744
R227 VTAIL.n447 VTAIL.n425 171.744
R228 VTAIL.n449 VTAIL.n447 171.744
R229 VTAIL.n449 VTAIL.n448 171.744
R230 VTAIL.n448 VTAIL.n421 171.744
R231 VTAIL.n457 VTAIL.n421 171.744
R232 VTAIL.n458 VTAIL.n457 171.744
R233 VTAIL.n458 VTAIL.n417 171.744
R234 VTAIL.n465 VTAIL.n417 171.744
R235 VTAIL.n466 VTAIL.n465 171.744
R236 VTAIL.n20 VTAIL.n17 171.744
R237 VTAIL.n27 VTAIL.n17 171.744
R238 VTAIL.n28 VTAIL.n27 171.744
R239 VTAIL.n28 VTAIL.n13 171.744
R240 VTAIL.n35 VTAIL.n13 171.744
R241 VTAIL.n37 VTAIL.n35 171.744
R242 VTAIL.n37 VTAIL.n36 171.744
R243 VTAIL.n36 VTAIL.n9 171.744
R244 VTAIL.n45 VTAIL.n9 171.744
R245 VTAIL.n46 VTAIL.n45 171.744
R246 VTAIL.n46 VTAIL.n5 171.744
R247 VTAIL.n53 VTAIL.n5 171.744
R248 VTAIL.n54 VTAIL.n53 171.744
R249 VTAIL.n78 VTAIL.n75 171.744
R250 VTAIL.n85 VTAIL.n75 171.744
R251 VTAIL.n86 VTAIL.n85 171.744
R252 VTAIL.n86 VTAIL.n71 171.744
R253 VTAIL.n93 VTAIL.n71 171.744
R254 VTAIL.n95 VTAIL.n93 171.744
R255 VTAIL.n95 VTAIL.n94 171.744
R256 VTAIL.n94 VTAIL.n67 171.744
R257 VTAIL.n103 VTAIL.n67 171.744
R258 VTAIL.n104 VTAIL.n103 171.744
R259 VTAIL.n104 VTAIL.n63 171.744
R260 VTAIL.n111 VTAIL.n63 171.744
R261 VTAIL.n112 VTAIL.n111 171.744
R262 VTAIL.n138 VTAIL.n135 171.744
R263 VTAIL.n145 VTAIL.n135 171.744
R264 VTAIL.n146 VTAIL.n145 171.744
R265 VTAIL.n146 VTAIL.n131 171.744
R266 VTAIL.n153 VTAIL.n131 171.744
R267 VTAIL.n155 VTAIL.n153 171.744
R268 VTAIL.n155 VTAIL.n154 171.744
R269 VTAIL.n154 VTAIL.n127 171.744
R270 VTAIL.n163 VTAIL.n127 171.744
R271 VTAIL.n164 VTAIL.n163 171.744
R272 VTAIL.n164 VTAIL.n123 171.744
R273 VTAIL.n171 VTAIL.n123 171.744
R274 VTAIL.n172 VTAIL.n171 171.744
R275 VTAIL.n408 VTAIL.n407 171.744
R276 VTAIL.n407 VTAIL.n359 171.744
R277 VTAIL.n400 VTAIL.n359 171.744
R278 VTAIL.n400 VTAIL.n399 171.744
R279 VTAIL.n399 VTAIL.n363 171.744
R280 VTAIL.n367 VTAIL.n363 171.744
R281 VTAIL.n391 VTAIL.n367 171.744
R282 VTAIL.n391 VTAIL.n390 171.744
R283 VTAIL.n390 VTAIL.n368 171.744
R284 VTAIL.n383 VTAIL.n368 171.744
R285 VTAIL.n383 VTAIL.n382 171.744
R286 VTAIL.n382 VTAIL.n372 171.744
R287 VTAIL.n375 VTAIL.n372 171.744
R288 VTAIL.n348 VTAIL.n347 171.744
R289 VTAIL.n347 VTAIL.n299 171.744
R290 VTAIL.n340 VTAIL.n299 171.744
R291 VTAIL.n340 VTAIL.n339 171.744
R292 VTAIL.n339 VTAIL.n303 171.744
R293 VTAIL.n307 VTAIL.n303 171.744
R294 VTAIL.n331 VTAIL.n307 171.744
R295 VTAIL.n331 VTAIL.n330 171.744
R296 VTAIL.n330 VTAIL.n308 171.744
R297 VTAIL.n323 VTAIL.n308 171.744
R298 VTAIL.n323 VTAIL.n322 171.744
R299 VTAIL.n322 VTAIL.n312 171.744
R300 VTAIL.n315 VTAIL.n312 171.744
R301 VTAIL.n290 VTAIL.n289 171.744
R302 VTAIL.n289 VTAIL.n241 171.744
R303 VTAIL.n282 VTAIL.n241 171.744
R304 VTAIL.n282 VTAIL.n281 171.744
R305 VTAIL.n281 VTAIL.n245 171.744
R306 VTAIL.n249 VTAIL.n245 171.744
R307 VTAIL.n273 VTAIL.n249 171.744
R308 VTAIL.n273 VTAIL.n272 171.744
R309 VTAIL.n272 VTAIL.n250 171.744
R310 VTAIL.n265 VTAIL.n250 171.744
R311 VTAIL.n265 VTAIL.n264 171.744
R312 VTAIL.n264 VTAIL.n254 171.744
R313 VTAIL.n257 VTAIL.n254 171.744
R314 VTAIL.n230 VTAIL.n229 171.744
R315 VTAIL.n229 VTAIL.n181 171.744
R316 VTAIL.n222 VTAIL.n181 171.744
R317 VTAIL.n222 VTAIL.n221 171.744
R318 VTAIL.n221 VTAIL.n185 171.744
R319 VTAIL.n189 VTAIL.n185 171.744
R320 VTAIL.n213 VTAIL.n189 171.744
R321 VTAIL.n213 VTAIL.n212 171.744
R322 VTAIL.n212 VTAIL.n190 171.744
R323 VTAIL.n205 VTAIL.n190 171.744
R324 VTAIL.n205 VTAIL.n204 171.744
R325 VTAIL.n204 VTAIL.n194 171.744
R326 VTAIL.n197 VTAIL.n194 171.744
R327 VTAIL.n432 VTAIL.t0 85.8723
R328 VTAIL.n20 VTAIL.t7 85.8723
R329 VTAIL.n78 VTAIL.t10 85.8723
R330 VTAIL.n138 VTAIL.t9 85.8723
R331 VTAIL.n375 VTAIL.t12 85.8723
R332 VTAIL.n315 VTAIL.t14 85.8723
R333 VTAIL.n257 VTAIL.t4 85.8723
R334 VTAIL.n197 VTAIL.t2 85.8723
R335 VTAIL.n355 VTAIL.n354 57.6359
R336 VTAIL.n237 VTAIL.n236 57.6359
R337 VTAIL.n1 VTAIL.n0 57.6357
R338 VTAIL.n119 VTAIL.n118 57.6357
R339 VTAIL.n471 VTAIL.n470 30.6338
R340 VTAIL.n59 VTAIL.n58 30.6338
R341 VTAIL.n117 VTAIL.n116 30.6338
R342 VTAIL.n177 VTAIL.n176 30.6338
R343 VTAIL.n413 VTAIL.n412 30.6338
R344 VTAIL.n353 VTAIL.n352 30.6338
R345 VTAIL.n295 VTAIL.n294 30.6338
R346 VTAIL.n235 VTAIL.n234 30.6338
R347 VTAIL.n471 VTAIL.n413 23.3669
R348 VTAIL.n235 VTAIL.n177 23.3669
R349 VTAIL.n456 VTAIL.n455 13.1884
R350 VTAIL.n44 VTAIL.n43 13.1884
R351 VTAIL.n102 VTAIL.n101 13.1884
R352 VTAIL.n162 VTAIL.n161 13.1884
R353 VTAIL.n398 VTAIL.n397 13.1884
R354 VTAIL.n338 VTAIL.n337 13.1884
R355 VTAIL.n280 VTAIL.n279 13.1884
R356 VTAIL.n220 VTAIL.n219 13.1884
R357 VTAIL.n454 VTAIL.n422 12.8005
R358 VTAIL.n459 VTAIL.n420 12.8005
R359 VTAIL.n42 VTAIL.n10 12.8005
R360 VTAIL.n47 VTAIL.n8 12.8005
R361 VTAIL.n100 VTAIL.n68 12.8005
R362 VTAIL.n105 VTAIL.n66 12.8005
R363 VTAIL.n160 VTAIL.n128 12.8005
R364 VTAIL.n165 VTAIL.n126 12.8005
R365 VTAIL.n401 VTAIL.n362 12.8005
R366 VTAIL.n396 VTAIL.n364 12.8005
R367 VTAIL.n341 VTAIL.n302 12.8005
R368 VTAIL.n336 VTAIL.n304 12.8005
R369 VTAIL.n283 VTAIL.n244 12.8005
R370 VTAIL.n278 VTAIL.n246 12.8005
R371 VTAIL.n223 VTAIL.n184 12.8005
R372 VTAIL.n218 VTAIL.n186 12.8005
R373 VTAIL.n451 VTAIL.n450 12.0247
R374 VTAIL.n460 VTAIL.n418 12.0247
R375 VTAIL.n39 VTAIL.n38 12.0247
R376 VTAIL.n48 VTAIL.n6 12.0247
R377 VTAIL.n97 VTAIL.n96 12.0247
R378 VTAIL.n106 VTAIL.n64 12.0247
R379 VTAIL.n157 VTAIL.n156 12.0247
R380 VTAIL.n166 VTAIL.n124 12.0247
R381 VTAIL.n402 VTAIL.n360 12.0247
R382 VTAIL.n393 VTAIL.n392 12.0247
R383 VTAIL.n342 VTAIL.n300 12.0247
R384 VTAIL.n333 VTAIL.n332 12.0247
R385 VTAIL.n284 VTAIL.n242 12.0247
R386 VTAIL.n275 VTAIL.n274 12.0247
R387 VTAIL.n224 VTAIL.n182 12.0247
R388 VTAIL.n215 VTAIL.n214 12.0247
R389 VTAIL.n446 VTAIL.n424 11.249
R390 VTAIL.n464 VTAIL.n463 11.249
R391 VTAIL.n34 VTAIL.n12 11.249
R392 VTAIL.n52 VTAIL.n51 11.249
R393 VTAIL.n92 VTAIL.n70 11.249
R394 VTAIL.n110 VTAIL.n109 11.249
R395 VTAIL.n152 VTAIL.n130 11.249
R396 VTAIL.n170 VTAIL.n169 11.249
R397 VTAIL.n406 VTAIL.n405 11.249
R398 VTAIL.n389 VTAIL.n366 11.249
R399 VTAIL.n346 VTAIL.n345 11.249
R400 VTAIL.n329 VTAIL.n306 11.249
R401 VTAIL.n288 VTAIL.n287 11.249
R402 VTAIL.n271 VTAIL.n248 11.249
R403 VTAIL.n228 VTAIL.n227 11.249
R404 VTAIL.n211 VTAIL.n188 11.249
R405 VTAIL.n433 VTAIL.n431 10.7239
R406 VTAIL.n21 VTAIL.n19 10.7239
R407 VTAIL.n79 VTAIL.n77 10.7239
R408 VTAIL.n139 VTAIL.n137 10.7239
R409 VTAIL.n376 VTAIL.n374 10.7239
R410 VTAIL.n316 VTAIL.n314 10.7239
R411 VTAIL.n258 VTAIL.n256 10.7239
R412 VTAIL.n198 VTAIL.n196 10.7239
R413 VTAIL.n445 VTAIL.n426 10.4732
R414 VTAIL.n467 VTAIL.n416 10.4732
R415 VTAIL.n33 VTAIL.n14 10.4732
R416 VTAIL.n55 VTAIL.n4 10.4732
R417 VTAIL.n91 VTAIL.n72 10.4732
R418 VTAIL.n113 VTAIL.n62 10.4732
R419 VTAIL.n151 VTAIL.n132 10.4732
R420 VTAIL.n173 VTAIL.n122 10.4732
R421 VTAIL.n409 VTAIL.n358 10.4732
R422 VTAIL.n388 VTAIL.n369 10.4732
R423 VTAIL.n349 VTAIL.n298 10.4732
R424 VTAIL.n328 VTAIL.n309 10.4732
R425 VTAIL.n291 VTAIL.n240 10.4732
R426 VTAIL.n270 VTAIL.n251 10.4732
R427 VTAIL.n231 VTAIL.n180 10.4732
R428 VTAIL.n210 VTAIL.n191 10.4732
R429 VTAIL.n442 VTAIL.n441 9.69747
R430 VTAIL.n468 VTAIL.n414 9.69747
R431 VTAIL.n30 VTAIL.n29 9.69747
R432 VTAIL.n56 VTAIL.n2 9.69747
R433 VTAIL.n88 VTAIL.n87 9.69747
R434 VTAIL.n114 VTAIL.n60 9.69747
R435 VTAIL.n148 VTAIL.n147 9.69747
R436 VTAIL.n174 VTAIL.n120 9.69747
R437 VTAIL.n410 VTAIL.n356 9.69747
R438 VTAIL.n385 VTAIL.n384 9.69747
R439 VTAIL.n350 VTAIL.n296 9.69747
R440 VTAIL.n325 VTAIL.n324 9.69747
R441 VTAIL.n292 VTAIL.n238 9.69747
R442 VTAIL.n267 VTAIL.n266 9.69747
R443 VTAIL.n232 VTAIL.n178 9.69747
R444 VTAIL.n207 VTAIL.n206 9.69747
R445 VTAIL.n470 VTAIL.n469 9.45567
R446 VTAIL.n58 VTAIL.n57 9.45567
R447 VTAIL.n116 VTAIL.n115 9.45567
R448 VTAIL.n176 VTAIL.n175 9.45567
R449 VTAIL.n412 VTAIL.n411 9.45567
R450 VTAIL.n352 VTAIL.n351 9.45567
R451 VTAIL.n294 VTAIL.n293 9.45567
R452 VTAIL.n234 VTAIL.n233 9.45567
R453 VTAIL.n469 VTAIL.n468 9.3005
R454 VTAIL.n416 VTAIL.n415 9.3005
R455 VTAIL.n463 VTAIL.n462 9.3005
R456 VTAIL.n461 VTAIL.n460 9.3005
R457 VTAIL.n420 VTAIL.n419 9.3005
R458 VTAIL.n435 VTAIL.n434 9.3005
R459 VTAIL.n437 VTAIL.n436 9.3005
R460 VTAIL.n428 VTAIL.n427 9.3005
R461 VTAIL.n443 VTAIL.n442 9.3005
R462 VTAIL.n445 VTAIL.n444 9.3005
R463 VTAIL.n424 VTAIL.n423 9.3005
R464 VTAIL.n452 VTAIL.n451 9.3005
R465 VTAIL.n454 VTAIL.n453 9.3005
R466 VTAIL.n57 VTAIL.n56 9.3005
R467 VTAIL.n4 VTAIL.n3 9.3005
R468 VTAIL.n51 VTAIL.n50 9.3005
R469 VTAIL.n49 VTAIL.n48 9.3005
R470 VTAIL.n8 VTAIL.n7 9.3005
R471 VTAIL.n23 VTAIL.n22 9.3005
R472 VTAIL.n25 VTAIL.n24 9.3005
R473 VTAIL.n16 VTAIL.n15 9.3005
R474 VTAIL.n31 VTAIL.n30 9.3005
R475 VTAIL.n33 VTAIL.n32 9.3005
R476 VTAIL.n12 VTAIL.n11 9.3005
R477 VTAIL.n40 VTAIL.n39 9.3005
R478 VTAIL.n42 VTAIL.n41 9.3005
R479 VTAIL.n115 VTAIL.n114 9.3005
R480 VTAIL.n62 VTAIL.n61 9.3005
R481 VTAIL.n109 VTAIL.n108 9.3005
R482 VTAIL.n107 VTAIL.n106 9.3005
R483 VTAIL.n66 VTAIL.n65 9.3005
R484 VTAIL.n81 VTAIL.n80 9.3005
R485 VTAIL.n83 VTAIL.n82 9.3005
R486 VTAIL.n74 VTAIL.n73 9.3005
R487 VTAIL.n89 VTAIL.n88 9.3005
R488 VTAIL.n91 VTAIL.n90 9.3005
R489 VTAIL.n70 VTAIL.n69 9.3005
R490 VTAIL.n98 VTAIL.n97 9.3005
R491 VTAIL.n100 VTAIL.n99 9.3005
R492 VTAIL.n175 VTAIL.n174 9.3005
R493 VTAIL.n122 VTAIL.n121 9.3005
R494 VTAIL.n169 VTAIL.n168 9.3005
R495 VTAIL.n167 VTAIL.n166 9.3005
R496 VTAIL.n126 VTAIL.n125 9.3005
R497 VTAIL.n141 VTAIL.n140 9.3005
R498 VTAIL.n143 VTAIL.n142 9.3005
R499 VTAIL.n134 VTAIL.n133 9.3005
R500 VTAIL.n149 VTAIL.n148 9.3005
R501 VTAIL.n151 VTAIL.n150 9.3005
R502 VTAIL.n130 VTAIL.n129 9.3005
R503 VTAIL.n158 VTAIL.n157 9.3005
R504 VTAIL.n160 VTAIL.n159 9.3005
R505 VTAIL.n378 VTAIL.n377 9.3005
R506 VTAIL.n380 VTAIL.n379 9.3005
R507 VTAIL.n371 VTAIL.n370 9.3005
R508 VTAIL.n386 VTAIL.n385 9.3005
R509 VTAIL.n388 VTAIL.n387 9.3005
R510 VTAIL.n366 VTAIL.n365 9.3005
R511 VTAIL.n394 VTAIL.n393 9.3005
R512 VTAIL.n396 VTAIL.n395 9.3005
R513 VTAIL.n411 VTAIL.n410 9.3005
R514 VTAIL.n358 VTAIL.n357 9.3005
R515 VTAIL.n405 VTAIL.n404 9.3005
R516 VTAIL.n403 VTAIL.n402 9.3005
R517 VTAIL.n362 VTAIL.n361 9.3005
R518 VTAIL.n318 VTAIL.n317 9.3005
R519 VTAIL.n320 VTAIL.n319 9.3005
R520 VTAIL.n311 VTAIL.n310 9.3005
R521 VTAIL.n326 VTAIL.n325 9.3005
R522 VTAIL.n328 VTAIL.n327 9.3005
R523 VTAIL.n306 VTAIL.n305 9.3005
R524 VTAIL.n334 VTAIL.n333 9.3005
R525 VTAIL.n336 VTAIL.n335 9.3005
R526 VTAIL.n351 VTAIL.n350 9.3005
R527 VTAIL.n298 VTAIL.n297 9.3005
R528 VTAIL.n345 VTAIL.n344 9.3005
R529 VTAIL.n343 VTAIL.n342 9.3005
R530 VTAIL.n302 VTAIL.n301 9.3005
R531 VTAIL.n260 VTAIL.n259 9.3005
R532 VTAIL.n262 VTAIL.n261 9.3005
R533 VTAIL.n253 VTAIL.n252 9.3005
R534 VTAIL.n268 VTAIL.n267 9.3005
R535 VTAIL.n270 VTAIL.n269 9.3005
R536 VTAIL.n248 VTAIL.n247 9.3005
R537 VTAIL.n276 VTAIL.n275 9.3005
R538 VTAIL.n278 VTAIL.n277 9.3005
R539 VTAIL.n293 VTAIL.n292 9.3005
R540 VTAIL.n240 VTAIL.n239 9.3005
R541 VTAIL.n287 VTAIL.n286 9.3005
R542 VTAIL.n285 VTAIL.n284 9.3005
R543 VTAIL.n244 VTAIL.n243 9.3005
R544 VTAIL.n200 VTAIL.n199 9.3005
R545 VTAIL.n202 VTAIL.n201 9.3005
R546 VTAIL.n193 VTAIL.n192 9.3005
R547 VTAIL.n208 VTAIL.n207 9.3005
R548 VTAIL.n210 VTAIL.n209 9.3005
R549 VTAIL.n188 VTAIL.n187 9.3005
R550 VTAIL.n216 VTAIL.n215 9.3005
R551 VTAIL.n218 VTAIL.n217 9.3005
R552 VTAIL.n233 VTAIL.n232 9.3005
R553 VTAIL.n180 VTAIL.n179 9.3005
R554 VTAIL.n227 VTAIL.n226 9.3005
R555 VTAIL.n225 VTAIL.n224 9.3005
R556 VTAIL.n184 VTAIL.n183 9.3005
R557 VTAIL.n438 VTAIL.n428 8.92171
R558 VTAIL.n26 VTAIL.n16 8.92171
R559 VTAIL.n84 VTAIL.n74 8.92171
R560 VTAIL.n144 VTAIL.n134 8.92171
R561 VTAIL.n381 VTAIL.n371 8.92171
R562 VTAIL.n321 VTAIL.n311 8.92171
R563 VTAIL.n263 VTAIL.n253 8.92171
R564 VTAIL.n203 VTAIL.n193 8.92171
R565 VTAIL.n437 VTAIL.n430 8.14595
R566 VTAIL.n25 VTAIL.n18 8.14595
R567 VTAIL.n83 VTAIL.n76 8.14595
R568 VTAIL.n143 VTAIL.n136 8.14595
R569 VTAIL.n380 VTAIL.n373 8.14595
R570 VTAIL.n320 VTAIL.n313 8.14595
R571 VTAIL.n262 VTAIL.n255 8.14595
R572 VTAIL.n202 VTAIL.n195 8.14595
R573 VTAIL.n434 VTAIL.n433 7.3702
R574 VTAIL.n22 VTAIL.n21 7.3702
R575 VTAIL.n80 VTAIL.n79 7.3702
R576 VTAIL.n140 VTAIL.n139 7.3702
R577 VTAIL.n377 VTAIL.n376 7.3702
R578 VTAIL.n317 VTAIL.n316 7.3702
R579 VTAIL.n259 VTAIL.n258 7.3702
R580 VTAIL.n199 VTAIL.n198 7.3702
R581 VTAIL.n434 VTAIL.n430 5.81868
R582 VTAIL.n22 VTAIL.n18 5.81868
R583 VTAIL.n80 VTAIL.n76 5.81868
R584 VTAIL.n140 VTAIL.n136 5.81868
R585 VTAIL.n377 VTAIL.n373 5.81868
R586 VTAIL.n317 VTAIL.n313 5.81868
R587 VTAIL.n259 VTAIL.n255 5.81868
R588 VTAIL.n199 VTAIL.n195 5.81868
R589 VTAIL.n438 VTAIL.n437 5.04292
R590 VTAIL.n26 VTAIL.n25 5.04292
R591 VTAIL.n84 VTAIL.n83 5.04292
R592 VTAIL.n144 VTAIL.n143 5.04292
R593 VTAIL.n381 VTAIL.n380 5.04292
R594 VTAIL.n321 VTAIL.n320 5.04292
R595 VTAIL.n263 VTAIL.n262 5.04292
R596 VTAIL.n203 VTAIL.n202 5.04292
R597 VTAIL.n441 VTAIL.n428 4.26717
R598 VTAIL.n470 VTAIL.n414 4.26717
R599 VTAIL.n29 VTAIL.n16 4.26717
R600 VTAIL.n58 VTAIL.n2 4.26717
R601 VTAIL.n87 VTAIL.n74 4.26717
R602 VTAIL.n116 VTAIL.n60 4.26717
R603 VTAIL.n147 VTAIL.n134 4.26717
R604 VTAIL.n176 VTAIL.n120 4.26717
R605 VTAIL.n412 VTAIL.n356 4.26717
R606 VTAIL.n384 VTAIL.n371 4.26717
R607 VTAIL.n352 VTAIL.n296 4.26717
R608 VTAIL.n324 VTAIL.n311 4.26717
R609 VTAIL.n294 VTAIL.n238 4.26717
R610 VTAIL.n266 VTAIL.n253 4.26717
R611 VTAIL.n234 VTAIL.n178 4.26717
R612 VTAIL.n206 VTAIL.n193 4.26717
R613 VTAIL.n442 VTAIL.n426 3.49141
R614 VTAIL.n468 VTAIL.n467 3.49141
R615 VTAIL.n30 VTAIL.n14 3.49141
R616 VTAIL.n56 VTAIL.n55 3.49141
R617 VTAIL.n88 VTAIL.n72 3.49141
R618 VTAIL.n114 VTAIL.n113 3.49141
R619 VTAIL.n148 VTAIL.n132 3.49141
R620 VTAIL.n174 VTAIL.n173 3.49141
R621 VTAIL.n410 VTAIL.n409 3.49141
R622 VTAIL.n385 VTAIL.n369 3.49141
R623 VTAIL.n350 VTAIL.n349 3.49141
R624 VTAIL.n325 VTAIL.n309 3.49141
R625 VTAIL.n292 VTAIL.n291 3.49141
R626 VTAIL.n267 VTAIL.n251 3.49141
R627 VTAIL.n232 VTAIL.n231 3.49141
R628 VTAIL.n207 VTAIL.n191 3.49141
R629 VTAIL.n0 VTAIL.t3 3.06701
R630 VTAIL.n0 VTAIL.t1 3.06701
R631 VTAIL.n118 VTAIL.t13 3.06701
R632 VTAIL.n118 VTAIL.t15 3.06701
R633 VTAIL.n354 VTAIL.t11 3.06701
R634 VTAIL.n354 VTAIL.t8 3.06701
R635 VTAIL.n236 VTAIL.t5 3.06701
R636 VTAIL.n236 VTAIL.t6 3.06701
R637 VTAIL.n446 VTAIL.n445 2.71565
R638 VTAIL.n464 VTAIL.n416 2.71565
R639 VTAIL.n34 VTAIL.n33 2.71565
R640 VTAIL.n52 VTAIL.n4 2.71565
R641 VTAIL.n92 VTAIL.n91 2.71565
R642 VTAIL.n110 VTAIL.n62 2.71565
R643 VTAIL.n152 VTAIL.n151 2.71565
R644 VTAIL.n170 VTAIL.n122 2.71565
R645 VTAIL.n406 VTAIL.n358 2.71565
R646 VTAIL.n389 VTAIL.n388 2.71565
R647 VTAIL.n346 VTAIL.n298 2.71565
R648 VTAIL.n329 VTAIL.n328 2.71565
R649 VTAIL.n288 VTAIL.n240 2.71565
R650 VTAIL.n271 VTAIL.n270 2.71565
R651 VTAIL.n228 VTAIL.n180 2.71565
R652 VTAIL.n211 VTAIL.n210 2.71565
R653 VTAIL.n435 VTAIL.n431 2.41282
R654 VTAIL.n23 VTAIL.n19 2.41282
R655 VTAIL.n81 VTAIL.n77 2.41282
R656 VTAIL.n141 VTAIL.n137 2.41282
R657 VTAIL.n378 VTAIL.n374 2.41282
R658 VTAIL.n318 VTAIL.n314 2.41282
R659 VTAIL.n260 VTAIL.n256 2.41282
R660 VTAIL.n200 VTAIL.n196 2.41282
R661 VTAIL.n450 VTAIL.n424 1.93989
R662 VTAIL.n463 VTAIL.n418 1.93989
R663 VTAIL.n38 VTAIL.n12 1.93989
R664 VTAIL.n51 VTAIL.n6 1.93989
R665 VTAIL.n96 VTAIL.n70 1.93989
R666 VTAIL.n109 VTAIL.n64 1.93989
R667 VTAIL.n156 VTAIL.n130 1.93989
R668 VTAIL.n169 VTAIL.n124 1.93989
R669 VTAIL.n405 VTAIL.n360 1.93989
R670 VTAIL.n392 VTAIL.n366 1.93989
R671 VTAIL.n345 VTAIL.n300 1.93989
R672 VTAIL.n332 VTAIL.n306 1.93989
R673 VTAIL.n287 VTAIL.n242 1.93989
R674 VTAIL.n274 VTAIL.n248 1.93989
R675 VTAIL.n227 VTAIL.n182 1.93989
R676 VTAIL.n214 VTAIL.n188 1.93989
R677 VTAIL.n237 VTAIL.n235 1.86257
R678 VTAIL.n295 VTAIL.n237 1.86257
R679 VTAIL.n355 VTAIL.n353 1.86257
R680 VTAIL.n413 VTAIL.n355 1.86257
R681 VTAIL.n177 VTAIL.n119 1.86257
R682 VTAIL.n119 VTAIL.n117 1.86257
R683 VTAIL.n59 VTAIL.n1 1.86257
R684 VTAIL VTAIL.n471 1.80438
R685 VTAIL.n451 VTAIL.n422 1.16414
R686 VTAIL.n460 VTAIL.n459 1.16414
R687 VTAIL.n39 VTAIL.n10 1.16414
R688 VTAIL.n48 VTAIL.n47 1.16414
R689 VTAIL.n97 VTAIL.n68 1.16414
R690 VTAIL.n106 VTAIL.n105 1.16414
R691 VTAIL.n157 VTAIL.n128 1.16414
R692 VTAIL.n166 VTAIL.n165 1.16414
R693 VTAIL.n402 VTAIL.n401 1.16414
R694 VTAIL.n393 VTAIL.n364 1.16414
R695 VTAIL.n342 VTAIL.n341 1.16414
R696 VTAIL.n333 VTAIL.n304 1.16414
R697 VTAIL.n284 VTAIL.n283 1.16414
R698 VTAIL.n275 VTAIL.n246 1.16414
R699 VTAIL.n224 VTAIL.n223 1.16414
R700 VTAIL.n215 VTAIL.n186 1.16414
R701 VTAIL.n353 VTAIL.n295 0.470328
R702 VTAIL.n117 VTAIL.n59 0.470328
R703 VTAIL.n455 VTAIL.n454 0.388379
R704 VTAIL.n456 VTAIL.n420 0.388379
R705 VTAIL.n43 VTAIL.n42 0.388379
R706 VTAIL.n44 VTAIL.n8 0.388379
R707 VTAIL.n101 VTAIL.n100 0.388379
R708 VTAIL.n102 VTAIL.n66 0.388379
R709 VTAIL.n161 VTAIL.n160 0.388379
R710 VTAIL.n162 VTAIL.n126 0.388379
R711 VTAIL.n398 VTAIL.n362 0.388379
R712 VTAIL.n397 VTAIL.n396 0.388379
R713 VTAIL.n338 VTAIL.n302 0.388379
R714 VTAIL.n337 VTAIL.n336 0.388379
R715 VTAIL.n280 VTAIL.n244 0.388379
R716 VTAIL.n279 VTAIL.n278 0.388379
R717 VTAIL.n220 VTAIL.n184 0.388379
R718 VTAIL.n219 VTAIL.n218 0.388379
R719 VTAIL.n436 VTAIL.n435 0.155672
R720 VTAIL.n436 VTAIL.n427 0.155672
R721 VTAIL.n443 VTAIL.n427 0.155672
R722 VTAIL.n444 VTAIL.n443 0.155672
R723 VTAIL.n444 VTAIL.n423 0.155672
R724 VTAIL.n452 VTAIL.n423 0.155672
R725 VTAIL.n453 VTAIL.n452 0.155672
R726 VTAIL.n453 VTAIL.n419 0.155672
R727 VTAIL.n461 VTAIL.n419 0.155672
R728 VTAIL.n462 VTAIL.n461 0.155672
R729 VTAIL.n462 VTAIL.n415 0.155672
R730 VTAIL.n469 VTAIL.n415 0.155672
R731 VTAIL.n24 VTAIL.n23 0.155672
R732 VTAIL.n24 VTAIL.n15 0.155672
R733 VTAIL.n31 VTAIL.n15 0.155672
R734 VTAIL.n32 VTAIL.n31 0.155672
R735 VTAIL.n32 VTAIL.n11 0.155672
R736 VTAIL.n40 VTAIL.n11 0.155672
R737 VTAIL.n41 VTAIL.n40 0.155672
R738 VTAIL.n41 VTAIL.n7 0.155672
R739 VTAIL.n49 VTAIL.n7 0.155672
R740 VTAIL.n50 VTAIL.n49 0.155672
R741 VTAIL.n50 VTAIL.n3 0.155672
R742 VTAIL.n57 VTAIL.n3 0.155672
R743 VTAIL.n82 VTAIL.n81 0.155672
R744 VTAIL.n82 VTAIL.n73 0.155672
R745 VTAIL.n89 VTAIL.n73 0.155672
R746 VTAIL.n90 VTAIL.n89 0.155672
R747 VTAIL.n90 VTAIL.n69 0.155672
R748 VTAIL.n98 VTAIL.n69 0.155672
R749 VTAIL.n99 VTAIL.n98 0.155672
R750 VTAIL.n99 VTAIL.n65 0.155672
R751 VTAIL.n107 VTAIL.n65 0.155672
R752 VTAIL.n108 VTAIL.n107 0.155672
R753 VTAIL.n108 VTAIL.n61 0.155672
R754 VTAIL.n115 VTAIL.n61 0.155672
R755 VTAIL.n142 VTAIL.n141 0.155672
R756 VTAIL.n142 VTAIL.n133 0.155672
R757 VTAIL.n149 VTAIL.n133 0.155672
R758 VTAIL.n150 VTAIL.n149 0.155672
R759 VTAIL.n150 VTAIL.n129 0.155672
R760 VTAIL.n158 VTAIL.n129 0.155672
R761 VTAIL.n159 VTAIL.n158 0.155672
R762 VTAIL.n159 VTAIL.n125 0.155672
R763 VTAIL.n167 VTAIL.n125 0.155672
R764 VTAIL.n168 VTAIL.n167 0.155672
R765 VTAIL.n168 VTAIL.n121 0.155672
R766 VTAIL.n175 VTAIL.n121 0.155672
R767 VTAIL.n411 VTAIL.n357 0.155672
R768 VTAIL.n404 VTAIL.n357 0.155672
R769 VTAIL.n404 VTAIL.n403 0.155672
R770 VTAIL.n403 VTAIL.n361 0.155672
R771 VTAIL.n395 VTAIL.n361 0.155672
R772 VTAIL.n395 VTAIL.n394 0.155672
R773 VTAIL.n394 VTAIL.n365 0.155672
R774 VTAIL.n387 VTAIL.n365 0.155672
R775 VTAIL.n387 VTAIL.n386 0.155672
R776 VTAIL.n386 VTAIL.n370 0.155672
R777 VTAIL.n379 VTAIL.n370 0.155672
R778 VTAIL.n379 VTAIL.n378 0.155672
R779 VTAIL.n351 VTAIL.n297 0.155672
R780 VTAIL.n344 VTAIL.n297 0.155672
R781 VTAIL.n344 VTAIL.n343 0.155672
R782 VTAIL.n343 VTAIL.n301 0.155672
R783 VTAIL.n335 VTAIL.n301 0.155672
R784 VTAIL.n335 VTAIL.n334 0.155672
R785 VTAIL.n334 VTAIL.n305 0.155672
R786 VTAIL.n327 VTAIL.n305 0.155672
R787 VTAIL.n327 VTAIL.n326 0.155672
R788 VTAIL.n326 VTAIL.n310 0.155672
R789 VTAIL.n319 VTAIL.n310 0.155672
R790 VTAIL.n319 VTAIL.n318 0.155672
R791 VTAIL.n293 VTAIL.n239 0.155672
R792 VTAIL.n286 VTAIL.n239 0.155672
R793 VTAIL.n286 VTAIL.n285 0.155672
R794 VTAIL.n285 VTAIL.n243 0.155672
R795 VTAIL.n277 VTAIL.n243 0.155672
R796 VTAIL.n277 VTAIL.n276 0.155672
R797 VTAIL.n276 VTAIL.n247 0.155672
R798 VTAIL.n269 VTAIL.n247 0.155672
R799 VTAIL.n269 VTAIL.n268 0.155672
R800 VTAIL.n268 VTAIL.n252 0.155672
R801 VTAIL.n261 VTAIL.n252 0.155672
R802 VTAIL.n261 VTAIL.n260 0.155672
R803 VTAIL.n233 VTAIL.n179 0.155672
R804 VTAIL.n226 VTAIL.n179 0.155672
R805 VTAIL.n226 VTAIL.n225 0.155672
R806 VTAIL.n225 VTAIL.n183 0.155672
R807 VTAIL.n217 VTAIL.n183 0.155672
R808 VTAIL.n217 VTAIL.n216 0.155672
R809 VTAIL.n216 VTAIL.n187 0.155672
R810 VTAIL.n209 VTAIL.n187 0.155672
R811 VTAIL.n209 VTAIL.n208 0.155672
R812 VTAIL.n208 VTAIL.n192 0.155672
R813 VTAIL.n201 VTAIL.n192 0.155672
R814 VTAIL.n201 VTAIL.n200 0.155672
R815 VTAIL VTAIL.n1 0.0586897
R816 VN.n4 VN.t6 171.28
R817 VN.n25 VN.t2 171.28
R818 VN.n39 VN.n21 161.3
R819 VN.n38 VN.n37 161.3
R820 VN.n36 VN.n22 161.3
R821 VN.n35 VN.n34 161.3
R822 VN.n32 VN.n23 161.3
R823 VN.n31 VN.n30 161.3
R824 VN.n29 VN.n24 161.3
R825 VN.n28 VN.n27 161.3
R826 VN.n18 VN.n0 161.3
R827 VN.n17 VN.n16 161.3
R828 VN.n15 VN.n1 161.3
R829 VN.n14 VN.n13 161.3
R830 VN.n11 VN.n2 161.3
R831 VN.n10 VN.n9 161.3
R832 VN.n8 VN.n3 161.3
R833 VN.n7 VN.n6 161.3
R834 VN.n5 VN.t0 139.596
R835 VN.n12 VN.t1 139.596
R836 VN.n19 VN.t5 139.596
R837 VN.n26 VN.t4 139.596
R838 VN.n33 VN.t3 139.596
R839 VN.n40 VN.t7 139.596
R840 VN.n20 VN.n19 86.8082
R841 VN.n41 VN.n40 86.8082
R842 VN.n10 VN.n3 56.5617
R843 VN.n31 VN.n24 56.5617
R844 VN.n5 VN.n4 53.8128
R845 VN.n26 VN.n25 53.8128
R846 VN.n17 VN.n1 49.296
R847 VN.n38 VN.n22 49.296
R848 VN VN.n41 46.5588
R849 VN.n18 VN.n17 31.8581
R850 VN.n39 VN.n38 31.8581
R851 VN.n6 VN.n3 24.5923
R852 VN.n11 VN.n10 24.5923
R853 VN.n13 VN.n1 24.5923
R854 VN.n27 VN.n24 24.5923
R855 VN.n34 VN.n22 24.5923
R856 VN.n32 VN.n31 24.5923
R857 VN.n19 VN.n18 24.1005
R858 VN.n40 VN.n39 24.1005
R859 VN.n6 VN.n5 16.2311
R860 VN.n12 VN.n11 16.2311
R861 VN.n27 VN.n26 16.2311
R862 VN.n33 VN.n32 16.2311
R863 VN.n28 VN.n25 12.6399
R864 VN.n7 VN.n4 12.6399
R865 VN.n13 VN.n12 8.36172
R866 VN.n34 VN.n33 8.36172
R867 VN.n41 VN.n21 0.278335
R868 VN.n20 VN.n0 0.278335
R869 VN.n37 VN.n21 0.189894
R870 VN.n37 VN.n36 0.189894
R871 VN.n36 VN.n35 0.189894
R872 VN.n35 VN.n23 0.189894
R873 VN.n30 VN.n23 0.189894
R874 VN.n30 VN.n29 0.189894
R875 VN.n29 VN.n28 0.189894
R876 VN.n8 VN.n7 0.189894
R877 VN.n9 VN.n8 0.189894
R878 VN.n9 VN.n2 0.189894
R879 VN.n14 VN.n2 0.189894
R880 VN.n15 VN.n14 0.189894
R881 VN.n16 VN.n15 0.189894
R882 VN.n16 VN.n0 0.189894
R883 VN VN.n20 0.153485
R884 VDD2.n2 VDD2.n1 75.1902
R885 VDD2.n2 VDD2.n0 75.1902
R886 VDD2 VDD2.n5 75.1873
R887 VDD2.n4 VDD2.n3 74.3146
R888 VDD2.n4 VDD2.n2 41.2325
R889 VDD2.n5 VDD2.t3 3.06701
R890 VDD2.n5 VDD2.t5 3.06701
R891 VDD2.n3 VDD2.t0 3.06701
R892 VDD2.n3 VDD2.t4 3.06701
R893 VDD2.n1 VDD2.t6 3.06701
R894 VDD2.n1 VDD2.t2 3.06701
R895 VDD2.n0 VDD2.t1 3.06701
R896 VDD2.n0 VDD2.t7 3.06701
R897 VDD2 VDD2.n4 0.989724
R898 B.n485 B.n68 585
R899 B.n487 B.n486 585
R900 B.n488 B.n67 585
R901 B.n490 B.n489 585
R902 B.n491 B.n66 585
R903 B.n493 B.n492 585
R904 B.n494 B.n65 585
R905 B.n496 B.n495 585
R906 B.n497 B.n64 585
R907 B.n499 B.n498 585
R908 B.n500 B.n63 585
R909 B.n502 B.n501 585
R910 B.n503 B.n62 585
R911 B.n505 B.n504 585
R912 B.n506 B.n61 585
R913 B.n508 B.n507 585
R914 B.n509 B.n60 585
R915 B.n511 B.n510 585
R916 B.n512 B.n59 585
R917 B.n514 B.n513 585
R918 B.n515 B.n58 585
R919 B.n517 B.n516 585
R920 B.n518 B.n57 585
R921 B.n520 B.n519 585
R922 B.n521 B.n56 585
R923 B.n523 B.n522 585
R924 B.n524 B.n55 585
R925 B.n526 B.n525 585
R926 B.n527 B.n54 585
R927 B.n529 B.n528 585
R928 B.n530 B.n53 585
R929 B.n532 B.n531 585
R930 B.n533 B.n52 585
R931 B.n535 B.n534 585
R932 B.n536 B.n51 585
R933 B.n538 B.n537 585
R934 B.n539 B.n50 585
R935 B.n541 B.n540 585
R936 B.n543 B.n47 585
R937 B.n545 B.n544 585
R938 B.n546 B.n46 585
R939 B.n548 B.n547 585
R940 B.n549 B.n45 585
R941 B.n551 B.n550 585
R942 B.n552 B.n44 585
R943 B.n554 B.n553 585
R944 B.n555 B.n41 585
R945 B.n558 B.n557 585
R946 B.n559 B.n40 585
R947 B.n561 B.n560 585
R948 B.n562 B.n39 585
R949 B.n564 B.n563 585
R950 B.n565 B.n38 585
R951 B.n567 B.n566 585
R952 B.n568 B.n37 585
R953 B.n570 B.n569 585
R954 B.n571 B.n36 585
R955 B.n573 B.n572 585
R956 B.n574 B.n35 585
R957 B.n576 B.n575 585
R958 B.n577 B.n34 585
R959 B.n579 B.n578 585
R960 B.n580 B.n33 585
R961 B.n582 B.n581 585
R962 B.n583 B.n32 585
R963 B.n585 B.n584 585
R964 B.n586 B.n31 585
R965 B.n588 B.n587 585
R966 B.n589 B.n30 585
R967 B.n591 B.n590 585
R968 B.n592 B.n29 585
R969 B.n594 B.n593 585
R970 B.n595 B.n28 585
R971 B.n597 B.n596 585
R972 B.n598 B.n27 585
R973 B.n600 B.n599 585
R974 B.n601 B.n26 585
R975 B.n603 B.n602 585
R976 B.n604 B.n25 585
R977 B.n606 B.n605 585
R978 B.n607 B.n24 585
R979 B.n609 B.n608 585
R980 B.n610 B.n23 585
R981 B.n612 B.n611 585
R982 B.n613 B.n22 585
R983 B.n484 B.n483 585
R984 B.n482 B.n69 585
R985 B.n481 B.n480 585
R986 B.n479 B.n70 585
R987 B.n478 B.n477 585
R988 B.n476 B.n71 585
R989 B.n475 B.n474 585
R990 B.n473 B.n72 585
R991 B.n472 B.n471 585
R992 B.n470 B.n73 585
R993 B.n469 B.n468 585
R994 B.n467 B.n74 585
R995 B.n466 B.n465 585
R996 B.n464 B.n75 585
R997 B.n463 B.n462 585
R998 B.n461 B.n76 585
R999 B.n460 B.n459 585
R1000 B.n458 B.n77 585
R1001 B.n457 B.n456 585
R1002 B.n455 B.n78 585
R1003 B.n454 B.n453 585
R1004 B.n452 B.n79 585
R1005 B.n451 B.n450 585
R1006 B.n449 B.n80 585
R1007 B.n448 B.n447 585
R1008 B.n446 B.n81 585
R1009 B.n445 B.n444 585
R1010 B.n443 B.n82 585
R1011 B.n442 B.n441 585
R1012 B.n440 B.n83 585
R1013 B.n439 B.n438 585
R1014 B.n437 B.n84 585
R1015 B.n436 B.n435 585
R1016 B.n434 B.n85 585
R1017 B.n433 B.n432 585
R1018 B.n431 B.n86 585
R1019 B.n430 B.n429 585
R1020 B.n428 B.n87 585
R1021 B.n427 B.n426 585
R1022 B.n425 B.n88 585
R1023 B.n424 B.n423 585
R1024 B.n422 B.n89 585
R1025 B.n421 B.n420 585
R1026 B.n419 B.n90 585
R1027 B.n418 B.n417 585
R1028 B.n416 B.n91 585
R1029 B.n415 B.n414 585
R1030 B.n413 B.n92 585
R1031 B.n412 B.n411 585
R1032 B.n410 B.n93 585
R1033 B.n409 B.n408 585
R1034 B.n407 B.n94 585
R1035 B.n406 B.n405 585
R1036 B.n404 B.n95 585
R1037 B.n403 B.n402 585
R1038 B.n401 B.n96 585
R1039 B.n400 B.n399 585
R1040 B.n398 B.n97 585
R1041 B.n397 B.n396 585
R1042 B.n395 B.n98 585
R1043 B.n394 B.n393 585
R1044 B.n392 B.n99 585
R1045 B.n391 B.n390 585
R1046 B.n389 B.n100 585
R1047 B.n388 B.n387 585
R1048 B.n386 B.n101 585
R1049 B.n385 B.n384 585
R1050 B.n383 B.n102 585
R1051 B.n382 B.n381 585
R1052 B.n380 B.n103 585
R1053 B.n379 B.n378 585
R1054 B.n377 B.n104 585
R1055 B.n376 B.n375 585
R1056 B.n374 B.n105 585
R1057 B.n373 B.n372 585
R1058 B.n371 B.n106 585
R1059 B.n370 B.n369 585
R1060 B.n368 B.n107 585
R1061 B.n367 B.n366 585
R1062 B.n365 B.n108 585
R1063 B.n364 B.n363 585
R1064 B.n235 B.n234 585
R1065 B.n236 B.n155 585
R1066 B.n238 B.n237 585
R1067 B.n239 B.n154 585
R1068 B.n241 B.n240 585
R1069 B.n242 B.n153 585
R1070 B.n244 B.n243 585
R1071 B.n245 B.n152 585
R1072 B.n247 B.n246 585
R1073 B.n248 B.n151 585
R1074 B.n250 B.n249 585
R1075 B.n251 B.n150 585
R1076 B.n253 B.n252 585
R1077 B.n254 B.n149 585
R1078 B.n256 B.n255 585
R1079 B.n257 B.n148 585
R1080 B.n259 B.n258 585
R1081 B.n260 B.n147 585
R1082 B.n262 B.n261 585
R1083 B.n263 B.n146 585
R1084 B.n265 B.n264 585
R1085 B.n266 B.n145 585
R1086 B.n268 B.n267 585
R1087 B.n269 B.n144 585
R1088 B.n271 B.n270 585
R1089 B.n272 B.n143 585
R1090 B.n274 B.n273 585
R1091 B.n275 B.n142 585
R1092 B.n277 B.n276 585
R1093 B.n278 B.n141 585
R1094 B.n280 B.n279 585
R1095 B.n281 B.n140 585
R1096 B.n283 B.n282 585
R1097 B.n284 B.n139 585
R1098 B.n286 B.n285 585
R1099 B.n287 B.n138 585
R1100 B.n289 B.n288 585
R1101 B.n290 B.n135 585
R1102 B.n293 B.n292 585
R1103 B.n294 B.n134 585
R1104 B.n296 B.n295 585
R1105 B.n297 B.n133 585
R1106 B.n299 B.n298 585
R1107 B.n300 B.n132 585
R1108 B.n302 B.n301 585
R1109 B.n303 B.n131 585
R1110 B.n305 B.n304 585
R1111 B.n307 B.n306 585
R1112 B.n308 B.n127 585
R1113 B.n310 B.n309 585
R1114 B.n311 B.n126 585
R1115 B.n313 B.n312 585
R1116 B.n314 B.n125 585
R1117 B.n316 B.n315 585
R1118 B.n317 B.n124 585
R1119 B.n319 B.n318 585
R1120 B.n320 B.n123 585
R1121 B.n322 B.n321 585
R1122 B.n323 B.n122 585
R1123 B.n325 B.n324 585
R1124 B.n326 B.n121 585
R1125 B.n328 B.n327 585
R1126 B.n329 B.n120 585
R1127 B.n331 B.n330 585
R1128 B.n332 B.n119 585
R1129 B.n334 B.n333 585
R1130 B.n335 B.n118 585
R1131 B.n337 B.n336 585
R1132 B.n338 B.n117 585
R1133 B.n340 B.n339 585
R1134 B.n341 B.n116 585
R1135 B.n343 B.n342 585
R1136 B.n344 B.n115 585
R1137 B.n346 B.n345 585
R1138 B.n347 B.n114 585
R1139 B.n349 B.n348 585
R1140 B.n350 B.n113 585
R1141 B.n352 B.n351 585
R1142 B.n353 B.n112 585
R1143 B.n355 B.n354 585
R1144 B.n356 B.n111 585
R1145 B.n358 B.n357 585
R1146 B.n359 B.n110 585
R1147 B.n361 B.n360 585
R1148 B.n362 B.n109 585
R1149 B.n233 B.n156 585
R1150 B.n232 B.n231 585
R1151 B.n230 B.n157 585
R1152 B.n229 B.n228 585
R1153 B.n227 B.n158 585
R1154 B.n226 B.n225 585
R1155 B.n224 B.n159 585
R1156 B.n223 B.n222 585
R1157 B.n221 B.n160 585
R1158 B.n220 B.n219 585
R1159 B.n218 B.n161 585
R1160 B.n217 B.n216 585
R1161 B.n215 B.n162 585
R1162 B.n214 B.n213 585
R1163 B.n212 B.n163 585
R1164 B.n211 B.n210 585
R1165 B.n209 B.n164 585
R1166 B.n208 B.n207 585
R1167 B.n206 B.n165 585
R1168 B.n205 B.n204 585
R1169 B.n203 B.n166 585
R1170 B.n202 B.n201 585
R1171 B.n200 B.n167 585
R1172 B.n199 B.n198 585
R1173 B.n197 B.n168 585
R1174 B.n196 B.n195 585
R1175 B.n194 B.n169 585
R1176 B.n193 B.n192 585
R1177 B.n191 B.n170 585
R1178 B.n190 B.n189 585
R1179 B.n188 B.n171 585
R1180 B.n187 B.n186 585
R1181 B.n185 B.n172 585
R1182 B.n184 B.n183 585
R1183 B.n182 B.n173 585
R1184 B.n181 B.n180 585
R1185 B.n179 B.n174 585
R1186 B.n178 B.n177 585
R1187 B.n176 B.n175 585
R1188 B.n2 B.n0 585
R1189 B.n673 B.n1 585
R1190 B.n672 B.n671 585
R1191 B.n670 B.n3 585
R1192 B.n669 B.n668 585
R1193 B.n667 B.n4 585
R1194 B.n666 B.n665 585
R1195 B.n664 B.n5 585
R1196 B.n663 B.n662 585
R1197 B.n661 B.n6 585
R1198 B.n660 B.n659 585
R1199 B.n658 B.n7 585
R1200 B.n657 B.n656 585
R1201 B.n655 B.n8 585
R1202 B.n654 B.n653 585
R1203 B.n652 B.n9 585
R1204 B.n651 B.n650 585
R1205 B.n649 B.n10 585
R1206 B.n648 B.n647 585
R1207 B.n646 B.n11 585
R1208 B.n645 B.n644 585
R1209 B.n643 B.n12 585
R1210 B.n642 B.n641 585
R1211 B.n640 B.n13 585
R1212 B.n639 B.n638 585
R1213 B.n637 B.n14 585
R1214 B.n636 B.n635 585
R1215 B.n634 B.n15 585
R1216 B.n633 B.n632 585
R1217 B.n631 B.n16 585
R1218 B.n630 B.n629 585
R1219 B.n628 B.n17 585
R1220 B.n627 B.n626 585
R1221 B.n625 B.n18 585
R1222 B.n624 B.n623 585
R1223 B.n622 B.n19 585
R1224 B.n621 B.n620 585
R1225 B.n619 B.n20 585
R1226 B.n618 B.n617 585
R1227 B.n616 B.n21 585
R1228 B.n615 B.n614 585
R1229 B.n675 B.n674 585
R1230 B.n234 B.n233 444.452
R1231 B.n614 B.n613 444.452
R1232 B.n364 B.n109 444.452
R1233 B.n485 B.n484 444.452
R1234 B.n128 B.t2 392.156
R1235 B.n48 B.t4 392.156
R1236 B.n136 B.t8 392.156
R1237 B.n42 B.t10 392.156
R1238 B.n129 B.t1 350.264
R1239 B.n49 B.t5 350.264
R1240 B.n137 B.t7 350.264
R1241 B.n43 B.t11 350.264
R1242 B.n128 B.t0 346.084
R1243 B.n136 B.t6 346.084
R1244 B.n42 B.t9 346.084
R1245 B.n48 B.t3 346.084
R1246 B.n233 B.n232 163.367
R1247 B.n232 B.n157 163.367
R1248 B.n228 B.n157 163.367
R1249 B.n228 B.n227 163.367
R1250 B.n227 B.n226 163.367
R1251 B.n226 B.n159 163.367
R1252 B.n222 B.n159 163.367
R1253 B.n222 B.n221 163.367
R1254 B.n221 B.n220 163.367
R1255 B.n220 B.n161 163.367
R1256 B.n216 B.n161 163.367
R1257 B.n216 B.n215 163.367
R1258 B.n215 B.n214 163.367
R1259 B.n214 B.n163 163.367
R1260 B.n210 B.n163 163.367
R1261 B.n210 B.n209 163.367
R1262 B.n209 B.n208 163.367
R1263 B.n208 B.n165 163.367
R1264 B.n204 B.n165 163.367
R1265 B.n204 B.n203 163.367
R1266 B.n203 B.n202 163.367
R1267 B.n202 B.n167 163.367
R1268 B.n198 B.n167 163.367
R1269 B.n198 B.n197 163.367
R1270 B.n197 B.n196 163.367
R1271 B.n196 B.n169 163.367
R1272 B.n192 B.n169 163.367
R1273 B.n192 B.n191 163.367
R1274 B.n191 B.n190 163.367
R1275 B.n190 B.n171 163.367
R1276 B.n186 B.n171 163.367
R1277 B.n186 B.n185 163.367
R1278 B.n185 B.n184 163.367
R1279 B.n184 B.n173 163.367
R1280 B.n180 B.n173 163.367
R1281 B.n180 B.n179 163.367
R1282 B.n179 B.n178 163.367
R1283 B.n178 B.n175 163.367
R1284 B.n175 B.n2 163.367
R1285 B.n674 B.n2 163.367
R1286 B.n674 B.n673 163.367
R1287 B.n673 B.n672 163.367
R1288 B.n672 B.n3 163.367
R1289 B.n668 B.n3 163.367
R1290 B.n668 B.n667 163.367
R1291 B.n667 B.n666 163.367
R1292 B.n666 B.n5 163.367
R1293 B.n662 B.n5 163.367
R1294 B.n662 B.n661 163.367
R1295 B.n661 B.n660 163.367
R1296 B.n660 B.n7 163.367
R1297 B.n656 B.n7 163.367
R1298 B.n656 B.n655 163.367
R1299 B.n655 B.n654 163.367
R1300 B.n654 B.n9 163.367
R1301 B.n650 B.n9 163.367
R1302 B.n650 B.n649 163.367
R1303 B.n649 B.n648 163.367
R1304 B.n648 B.n11 163.367
R1305 B.n644 B.n11 163.367
R1306 B.n644 B.n643 163.367
R1307 B.n643 B.n642 163.367
R1308 B.n642 B.n13 163.367
R1309 B.n638 B.n13 163.367
R1310 B.n638 B.n637 163.367
R1311 B.n637 B.n636 163.367
R1312 B.n636 B.n15 163.367
R1313 B.n632 B.n15 163.367
R1314 B.n632 B.n631 163.367
R1315 B.n631 B.n630 163.367
R1316 B.n630 B.n17 163.367
R1317 B.n626 B.n17 163.367
R1318 B.n626 B.n625 163.367
R1319 B.n625 B.n624 163.367
R1320 B.n624 B.n19 163.367
R1321 B.n620 B.n19 163.367
R1322 B.n620 B.n619 163.367
R1323 B.n619 B.n618 163.367
R1324 B.n618 B.n21 163.367
R1325 B.n614 B.n21 163.367
R1326 B.n234 B.n155 163.367
R1327 B.n238 B.n155 163.367
R1328 B.n239 B.n238 163.367
R1329 B.n240 B.n239 163.367
R1330 B.n240 B.n153 163.367
R1331 B.n244 B.n153 163.367
R1332 B.n245 B.n244 163.367
R1333 B.n246 B.n245 163.367
R1334 B.n246 B.n151 163.367
R1335 B.n250 B.n151 163.367
R1336 B.n251 B.n250 163.367
R1337 B.n252 B.n251 163.367
R1338 B.n252 B.n149 163.367
R1339 B.n256 B.n149 163.367
R1340 B.n257 B.n256 163.367
R1341 B.n258 B.n257 163.367
R1342 B.n258 B.n147 163.367
R1343 B.n262 B.n147 163.367
R1344 B.n263 B.n262 163.367
R1345 B.n264 B.n263 163.367
R1346 B.n264 B.n145 163.367
R1347 B.n268 B.n145 163.367
R1348 B.n269 B.n268 163.367
R1349 B.n270 B.n269 163.367
R1350 B.n270 B.n143 163.367
R1351 B.n274 B.n143 163.367
R1352 B.n275 B.n274 163.367
R1353 B.n276 B.n275 163.367
R1354 B.n276 B.n141 163.367
R1355 B.n280 B.n141 163.367
R1356 B.n281 B.n280 163.367
R1357 B.n282 B.n281 163.367
R1358 B.n282 B.n139 163.367
R1359 B.n286 B.n139 163.367
R1360 B.n287 B.n286 163.367
R1361 B.n288 B.n287 163.367
R1362 B.n288 B.n135 163.367
R1363 B.n293 B.n135 163.367
R1364 B.n294 B.n293 163.367
R1365 B.n295 B.n294 163.367
R1366 B.n295 B.n133 163.367
R1367 B.n299 B.n133 163.367
R1368 B.n300 B.n299 163.367
R1369 B.n301 B.n300 163.367
R1370 B.n301 B.n131 163.367
R1371 B.n305 B.n131 163.367
R1372 B.n306 B.n305 163.367
R1373 B.n306 B.n127 163.367
R1374 B.n310 B.n127 163.367
R1375 B.n311 B.n310 163.367
R1376 B.n312 B.n311 163.367
R1377 B.n312 B.n125 163.367
R1378 B.n316 B.n125 163.367
R1379 B.n317 B.n316 163.367
R1380 B.n318 B.n317 163.367
R1381 B.n318 B.n123 163.367
R1382 B.n322 B.n123 163.367
R1383 B.n323 B.n322 163.367
R1384 B.n324 B.n323 163.367
R1385 B.n324 B.n121 163.367
R1386 B.n328 B.n121 163.367
R1387 B.n329 B.n328 163.367
R1388 B.n330 B.n329 163.367
R1389 B.n330 B.n119 163.367
R1390 B.n334 B.n119 163.367
R1391 B.n335 B.n334 163.367
R1392 B.n336 B.n335 163.367
R1393 B.n336 B.n117 163.367
R1394 B.n340 B.n117 163.367
R1395 B.n341 B.n340 163.367
R1396 B.n342 B.n341 163.367
R1397 B.n342 B.n115 163.367
R1398 B.n346 B.n115 163.367
R1399 B.n347 B.n346 163.367
R1400 B.n348 B.n347 163.367
R1401 B.n348 B.n113 163.367
R1402 B.n352 B.n113 163.367
R1403 B.n353 B.n352 163.367
R1404 B.n354 B.n353 163.367
R1405 B.n354 B.n111 163.367
R1406 B.n358 B.n111 163.367
R1407 B.n359 B.n358 163.367
R1408 B.n360 B.n359 163.367
R1409 B.n360 B.n109 163.367
R1410 B.n365 B.n364 163.367
R1411 B.n366 B.n365 163.367
R1412 B.n366 B.n107 163.367
R1413 B.n370 B.n107 163.367
R1414 B.n371 B.n370 163.367
R1415 B.n372 B.n371 163.367
R1416 B.n372 B.n105 163.367
R1417 B.n376 B.n105 163.367
R1418 B.n377 B.n376 163.367
R1419 B.n378 B.n377 163.367
R1420 B.n378 B.n103 163.367
R1421 B.n382 B.n103 163.367
R1422 B.n383 B.n382 163.367
R1423 B.n384 B.n383 163.367
R1424 B.n384 B.n101 163.367
R1425 B.n388 B.n101 163.367
R1426 B.n389 B.n388 163.367
R1427 B.n390 B.n389 163.367
R1428 B.n390 B.n99 163.367
R1429 B.n394 B.n99 163.367
R1430 B.n395 B.n394 163.367
R1431 B.n396 B.n395 163.367
R1432 B.n396 B.n97 163.367
R1433 B.n400 B.n97 163.367
R1434 B.n401 B.n400 163.367
R1435 B.n402 B.n401 163.367
R1436 B.n402 B.n95 163.367
R1437 B.n406 B.n95 163.367
R1438 B.n407 B.n406 163.367
R1439 B.n408 B.n407 163.367
R1440 B.n408 B.n93 163.367
R1441 B.n412 B.n93 163.367
R1442 B.n413 B.n412 163.367
R1443 B.n414 B.n413 163.367
R1444 B.n414 B.n91 163.367
R1445 B.n418 B.n91 163.367
R1446 B.n419 B.n418 163.367
R1447 B.n420 B.n419 163.367
R1448 B.n420 B.n89 163.367
R1449 B.n424 B.n89 163.367
R1450 B.n425 B.n424 163.367
R1451 B.n426 B.n425 163.367
R1452 B.n426 B.n87 163.367
R1453 B.n430 B.n87 163.367
R1454 B.n431 B.n430 163.367
R1455 B.n432 B.n431 163.367
R1456 B.n432 B.n85 163.367
R1457 B.n436 B.n85 163.367
R1458 B.n437 B.n436 163.367
R1459 B.n438 B.n437 163.367
R1460 B.n438 B.n83 163.367
R1461 B.n442 B.n83 163.367
R1462 B.n443 B.n442 163.367
R1463 B.n444 B.n443 163.367
R1464 B.n444 B.n81 163.367
R1465 B.n448 B.n81 163.367
R1466 B.n449 B.n448 163.367
R1467 B.n450 B.n449 163.367
R1468 B.n450 B.n79 163.367
R1469 B.n454 B.n79 163.367
R1470 B.n455 B.n454 163.367
R1471 B.n456 B.n455 163.367
R1472 B.n456 B.n77 163.367
R1473 B.n460 B.n77 163.367
R1474 B.n461 B.n460 163.367
R1475 B.n462 B.n461 163.367
R1476 B.n462 B.n75 163.367
R1477 B.n466 B.n75 163.367
R1478 B.n467 B.n466 163.367
R1479 B.n468 B.n467 163.367
R1480 B.n468 B.n73 163.367
R1481 B.n472 B.n73 163.367
R1482 B.n473 B.n472 163.367
R1483 B.n474 B.n473 163.367
R1484 B.n474 B.n71 163.367
R1485 B.n478 B.n71 163.367
R1486 B.n479 B.n478 163.367
R1487 B.n480 B.n479 163.367
R1488 B.n480 B.n69 163.367
R1489 B.n484 B.n69 163.367
R1490 B.n613 B.n612 163.367
R1491 B.n612 B.n23 163.367
R1492 B.n608 B.n23 163.367
R1493 B.n608 B.n607 163.367
R1494 B.n607 B.n606 163.367
R1495 B.n606 B.n25 163.367
R1496 B.n602 B.n25 163.367
R1497 B.n602 B.n601 163.367
R1498 B.n601 B.n600 163.367
R1499 B.n600 B.n27 163.367
R1500 B.n596 B.n27 163.367
R1501 B.n596 B.n595 163.367
R1502 B.n595 B.n594 163.367
R1503 B.n594 B.n29 163.367
R1504 B.n590 B.n29 163.367
R1505 B.n590 B.n589 163.367
R1506 B.n589 B.n588 163.367
R1507 B.n588 B.n31 163.367
R1508 B.n584 B.n31 163.367
R1509 B.n584 B.n583 163.367
R1510 B.n583 B.n582 163.367
R1511 B.n582 B.n33 163.367
R1512 B.n578 B.n33 163.367
R1513 B.n578 B.n577 163.367
R1514 B.n577 B.n576 163.367
R1515 B.n576 B.n35 163.367
R1516 B.n572 B.n35 163.367
R1517 B.n572 B.n571 163.367
R1518 B.n571 B.n570 163.367
R1519 B.n570 B.n37 163.367
R1520 B.n566 B.n37 163.367
R1521 B.n566 B.n565 163.367
R1522 B.n565 B.n564 163.367
R1523 B.n564 B.n39 163.367
R1524 B.n560 B.n39 163.367
R1525 B.n560 B.n559 163.367
R1526 B.n559 B.n558 163.367
R1527 B.n558 B.n41 163.367
R1528 B.n553 B.n41 163.367
R1529 B.n553 B.n552 163.367
R1530 B.n552 B.n551 163.367
R1531 B.n551 B.n45 163.367
R1532 B.n547 B.n45 163.367
R1533 B.n547 B.n546 163.367
R1534 B.n546 B.n545 163.367
R1535 B.n545 B.n47 163.367
R1536 B.n540 B.n47 163.367
R1537 B.n540 B.n539 163.367
R1538 B.n539 B.n538 163.367
R1539 B.n538 B.n51 163.367
R1540 B.n534 B.n51 163.367
R1541 B.n534 B.n533 163.367
R1542 B.n533 B.n532 163.367
R1543 B.n532 B.n53 163.367
R1544 B.n528 B.n53 163.367
R1545 B.n528 B.n527 163.367
R1546 B.n527 B.n526 163.367
R1547 B.n526 B.n55 163.367
R1548 B.n522 B.n55 163.367
R1549 B.n522 B.n521 163.367
R1550 B.n521 B.n520 163.367
R1551 B.n520 B.n57 163.367
R1552 B.n516 B.n57 163.367
R1553 B.n516 B.n515 163.367
R1554 B.n515 B.n514 163.367
R1555 B.n514 B.n59 163.367
R1556 B.n510 B.n59 163.367
R1557 B.n510 B.n509 163.367
R1558 B.n509 B.n508 163.367
R1559 B.n508 B.n61 163.367
R1560 B.n504 B.n61 163.367
R1561 B.n504 B.n503 163.367
R1562 B.n503 B.n502 163.367
R1563 B.n502 B.n63 163.367
R1564 B.n498 B.n63 163.367
R1565 B.n498 B.n497 163.367
R1566 B.n497 B.n496 163.367
R1567 B.n496 B.n65 163.367
R1568 B.n492 B.n65 163.367
R1569 B.n492 B.n491 163.367
R1570 B.n491 B.n490 163.367
R1571 B.n490 B.n67 163.367
R1572 B.n486 B.n67 163.367
R1573 B.n486 B.n485 163.367
R1574 B.n130 B.n129 59.5399
R1575 B.n291 B.n137 59.5399
R1576 B.n556 B.n43 59.5399
R1577 B.n542 B.n49 59.5399
R1578 B.n129 B.n128 41.8914
R1579 B.n137 B.n136 41.8914
R1580 B.n43 B.n42 41.8914
R1581 B.n49 B.n48 41.8914
R1582 B.n483 B.n68 28.8785
R1583 B.n615 B.n22 28.8785
R1584 B.n363 B.n362 28.8785
R1585 B.n235 B.n156 28.8785
R1586 B B.n675 18.0485
R1587 B.n611 B.n22 10.6151
R1588 B.n611 B.n610 10.6151
R1589 B.n610 B.n609 10.6151
R1590 B.n609 B.n24 10.6151
R1591 B.n605 B.n24 10.6151
R1592 B.n605 B.n604 10.6151
R1593 B.n604 B.n603 10.6151
R1594 B.n603 B.n26 10.6151
R1595 B.n599 B.n26 10.6151
R1596 B.n599 B.n598 10.6151
R1597 B.n598 B.n597 10.6151
R1598 B.n597 B.n28 10.6151
R1599 B.n593 B.n28 10.6151
R1600 B.n593 B.n592 10.6151
R1601 B.n592 B.n591 10.6151
R1602 B.n591 B.n30 10.6151
R1603 B.n587 B.n30 10.6151
R1604 B.n587 B.n586 10.6151
R1605 B.n586 B.n585 10.6151
R1606 B.n585 B.n32 10.6151
R1607 B.n581 B.n32 10.6151
R1608 B.n581 B.n580 10.6151
R1609 B.n580 B.n579 10.6151
R1610 B.n579 B.n34 10.6151
R1611 B.n575 B.n34 10.6151
R1612 B.n575 B.n574 10.6151
R1613 B.n574 B.n573 10.6151
R1614 B.n573 B.n36 10.6151
R1615 B.n569 B.n36 10.6151
R1616 B.n569 B.n568 10.6151
R1617 B.n568 B.n567 10.6151
R1618 B.n567 B.n38 10.6151
R1619 B.n563 B.n38 10.6151
R1620 B.n563 B.n562 10.6151
R1621 B.n562 B.n561 10.6151
R1622 B.n561 B.n40 10.6151
R1623 B.n557 B.n40 10.6151
R1624 B.n555 B.n554 10.6151
R1625 B.n554 B.n44 10.6151
R1626 B.n550 B.n44 10.6151
R1627 B.n550 B.n549 10.6151
R1628 B.n549 B.n548 10.6151
R1629 B.n548 B.n46 10.6151
R1630 B.n544 B.n46 10.6151
R1631 B.n544 B.n543 10.6151
R1632 B.n541 B.n50 10.6151
R1633 B.n537 B.n50 10.6151
R1634 B.n537 B.n536 10.6151
R1635 B.n536 B.n535 10.6151
R1636 B.n535 B.n52 10.6151
R1637 B.n531 B.n52 10.6151
R1638 B.n531 B.n530 10.6151
R1639 B.n530 B.n529 10.6151
R1640 B.n529 B.n54 10.6151
R1641 B.n525 B.n54 10.6151
R1642 B.n525 B.n524 10.6151
R1643 B.n524 B.n523 10.6151
R1644 B.n523 B.n56 10.6151
R1645 B.n519 B.n56 10.6151
R1646 B.n519 B.n518 10.6151
R1647 B.n518 B.n517 10.6151
R1648 B.n517 B.n58 10.6151
R1649 B.n513 B.n58 10.6151
R1650 B.n513 B.n512 10.6151
R1651 B.n512 B.n511 10.6151
R1652 B.n511 B.n60 10.6151
R1653 B.n507 B.n60 10.6151
R1654 B.n507 B.n506 10.6151
R1655 B.n506 B.n505 10.6151
R1656 B.n505 B.n62 10.6151
R1657 B.n501 B.n62 10.6151
R1658 B.n501 B.n500 10.6151
R1659 B.n500 B.n499 10.6151
R1660 B.n499 B.n64 10.6151
R1661 B.n495 B.n64 10.6151
R1662 B.n495 B.n494 10.6151
R1663 B.n494 B.n493 10.6151
R1664 B.n493 B.n66 10.6151
R1665 B.n489 B.n66 10.6151
R1666 B.n489 B.n488 10.6151
R1667 B.n488 B.n487 10.6151
R1668 B.n487 B.n68 10.6151
R1669 B.n363 B.n108 10.6151
R1670 B.n367 B.n108 10.6151
R1671 B.n368 B.n367 10.6151
R1672 B.n369 B.n368 10.6151
R1673 B.n369 B.n106 10.6151
R1674 B.n373 B.n106 10.6151
R1675 B.n374 B.n373 10.6151
R1676 B.n375 B.n374 10.6151
R1677 B.n375 B.n104 10.6151
R1678 B.n379 B.n104 10.6151
R1679 B.n380 B.n379 10.6151
R1680 B.n381 B.n380 10.6151
R1681 B.n381 B.n102 10.6151
R1682 B.n385 B.n102 10.6151
R1683 B.n386 B.n385 10.6151
R1684 B.n387 B.n386 10.6151
R1685 B.n387 B.n100 10.6151
R1686 B.n391 B.n100 10.6151
R1687 B.n392 B.n391 10.6151
R1688 B.n393 B.n392 10.6151
R1689 B.n393 B.n98 10.6151
R1690 B.n397 B.n98 10.6151
R1691 B.n398 B.n397 10.6151
R1692 B.n399 B.n398 10.6151
R1693 B.n399 B.n96 10.6151
R1694 B.n403 B.n96 10.6151
R1695 B.n404 B.n403 10.6151
R1696 B.n405 B.n404 10.6151
R1697 B.n405 B.n94 10.6151
R1698 B.n409 B.n94 10.6151
R1699 B.n410 B.n409 10.6151
R1700 B.n411 B.n410 10.6151
R1701 B.n411 B.n92 10.6151
R1702 B.n415 B.n92 10.6151
R1703 B.n416 B.n415 10.6151
R1704 B.n417 B.n416 10.6151
R1705 B.n417 B.n90 10.6151
R1706 B.n421 B.n90 10.6151
R1707 B.n422 B.n421 10.6151
R1708 B.n423 B.n422 10.6151
R1709 B.n423 B.n88 10.6151
R1710 B.n427 B.n88 10.6151
R1711 B.n428 B.n427 10.6151
R1712 B.n429 B.n428 10.6151
R1713 B.n429 B.n86 10.6151
R1714 B.n433 B.n86 10.6151
R1715 B.n434 B.n433 10.6151
R1716 B.n435 B.n434 10.6151
R1717 B.n435 B.n84 10.6151
R1718 B.n439 B.n84 10.6151
R1719 B.n440 B.n439 10.6151
R1720 B.n441 B.n440 10.6151
R1721 B.n441 B.n82 10.6151
R1722 B.n445 B.n82 10.6151
R1723 B.n446 B.n445 10.6151
R1724 B.n447 B.n446 10.6151
R1725 B.n447 B.n80 10.6151
R1726 B.n451 B.n80 10.6151
R1727 B.n452 B.n451 10.6151
R1728 B.n453 B.n452 10.6151
R1729 B.n453 B.n78 10.6151
R1730 B.n457 B.n78 10.6151
R1731 B.n458 B.n457 10.6151
R1732 B.n459 B.n458 10.6151
R1733 B.n459 B.n76 10.6151
R1734 B.n463 B.n76 10.6151
R1735 B.n464 B.n463 10.6151
R1736 B.n465 B.n464 10.6151
R1737 B.n465 B.n74 10.6151
R1738 B.n469 B.n74 10.6151
R1739 B.n470 B.n469 10.6151
R1740 B.n471 B.n470 10.6151
R1741 B.n471 B.n72 10.6151
R1742 B.n475 B.n72 10.6151
R1743 B.n476 B.n475 10.6151
R1744 B.n477 B.n476 10.6151
R1745 B.n477 B.n70 10.6151
R1746 B.n481 B.n70 10.6151
R1747 B.n482 B.n481 10.6151
R1748 B.n483 B.n482 10.6151
R1749 B.n236 B.n235 10.6151
R1750 B.n237 B.n236 10.6151
R1751 B.n237 B.n154 10.6151
R1752 B.n241 B.n154 10.6151
R1753 B.n242 B.n241 10.6151
R1754 B.n243 B.n242 10.6151
R1755 B.n243 B.n152 10.6151
R1756 B.n247 B.n152 10.6151
R1757 B.n248 B.n247 10.6151
R1758 B.n249 B.n248 10.6151
R1759 B.n249 B.n150 10.6151
R1760 B.n253 B.n150 10.6151
R1761 B.n254 B.n253 10.6151
R1762 B.n255 B.n254 10.6151
R1763 B.n255 B.n148 10.6151
R1764 B.n259 B.n148 10.6151
R1765 B.n260 B.n259 10.6151
R1766 B.n261 B.n260 10.6151
R1767 B.n261 B.n146 10.6151
R1768 B.n265 B.n146 10.6151
R1769 B.n266 B.n265 10.6151
R1770 B.n267 B.n266 10.6151
R1771 B.n267 B.n144 10.6151
R1772 B.n271 B.n144 10.6151
R1773 B.n272 B.n271 10.6151
R1774 B.n273 B.n272 10.6151
R1775 B.n273 B.n142 10.6151
R1776 B.n277 B.n142 10.6151
R1777 B.n278 B.n277 10.6151
R1778 B.n279 B.n278 10.6151
R1779 B.n279 B.n140 10.6151
R1780 B.n283 B.n140 10.6151
R1781 B.n284 B.n283 10.6151
R1782 B.n285 B.n284 10.6151
R1783 B.n285 B.n138 10.6151
R1784 B.n289 B.n138 10.6151
R1785 B.n290 B.n289 10.6151
R1786 B.n292 B.n134 10.6151
R1787 B.n296 B.n134 10.6151
R1788 B.n297 B.n296 10.6151
R1789 B.n298 B.n297 10.6151
R1790 B.n298 B.n132 10.6151
R1791 B.n302 B.n132 10.6151
R1792 B.n303 B.n302 10.6151
R1793 B.n304 B.n303 10.6151
R1794 B.n308 B.n307 10.6151
R1795 B.n309 B.n308 10.6151
R1796 B.n309 B.n126 10.6151
R1797 B.n313 B.n126 10.6151
R1798 B.n314 B.n313 10.6151
R1799 B.n315 B.n314 10.6151
R1800 B.n315 B.n124 10.6151
R1801 B.n319 B.n124 10.6151
R1802 B.n320 B.n319 10.6151
R1803 B.n321 B.n320 10.6151
R1804 B.n321 B.n122 10.6151
R1805 B.n325 B.n122 10.6151
R1806 B.n326 B.n325 10.6151
R1807 B.n327 B.n326 10.6151
R1808 B.n327 B.n120 10.6151
R1809 B.n331 B.n120 10.6151
R1810 B.n332 B.n331 10.6151
R1811 B.n333 B.n332 10.6151
R1812 B.n333 B.n118 10.6151
R1813 B.n337 B.n118 10.6151
R1814 B.n338 B.n337 10.6151
R1815 B.n339 B.n338 10.6151
R1816 B.n339 B.n116 10.6151
R1817 B.n343 B.n116 10.6151
R1818 B.n344 B.n343 10.6151
R1819 B.n345 B.n344 10.6151
R1820 B.n345 B.n114 10.6151
R1821 B.n349 B.n114 10.6151
R1822 B.n350 B.n349 10.6151
R1823 B.n351 B.n350 10.6151
R1824 B.n351 B.n112 10.6151
R1825 B.n355 B.n112 10.6151
R1826 B.n356 B.n355 10.6151
R1827 B.n357 B.n356 10.6151
R1828 B.n357 B.n110 10.6151
R1829 B.n361 B.n110 10.6151
R1830 B.n362 B.n361 10.6151
R1831 B.n231 B.n156 10.6151
R1832 B.n231 B.n230 10.6151
R1833 B.n230 B.n229 10.6151
R1834 B.n229 B.n158 10.6151
R1835 B.n225 B.n158 10.6151
R1836 B.n225 B.n224 10.6151
R1837 B.n224 B.n223 10.6151
R1838 B.n223 B.n160 10.6151
R1839 B.n219 B.n160 10.6151
R1840 B.n219 B.n218 10.6151
R1841 B.n218 B.n217 10.6151
R1842 B.n217 B.n162 10.6151
R1843 B.n213 B.n162 10.6151
R1844 B.n213 B.n212 10.6151
R1845 B.n212 B.n211 10.6151
R1846 B.n211 B.n164 10.6151
R1847 B.n207 B.n164 10.6151
R1848 B.n207 B.n206 10.6151
R1849 B.n206 B.n205 10.6151
R1850 B.n205 B.n166 10.6151
R1851 B.n201 B.n166 10.6151
R1852 B.n201 B.n200 10.6151
R1853 B.n200 B.n199 10.6151
R1854 B.n199 B.n168 10.6151
R1855 B.n195 B.n168 10.6151
R1856 B.n195 B.n194 10.6151
R1857 B.n194 B.n193 10.6151
R1858 B.n193 B.n170 10.6151
R1859 B.n189 B.n170 10.6151
R1860 B.n189 B.n188 10.6151
R1861 B.n188 B.n187 10.6151
R1862 B.n187 B.n172 10.6151
R1863 B.n183 B.n172 10.6151
R1864 B.n183 B.n182 10.6151
R1865 B.n182 B.n181 10.6151
R1866 B.n181 B.n174 10.6151
R1867 B.n177 B.n174 10.6151
R1868 B.n177 B.n176 10.6151
R1869 B.n176 B.n0 10.6151
R1870 B.n671 B.n1 10.6151
R1871 B.n671 B.n670 10.6151
R1872 B.n670 B.n669 10.6151
R1873 B.n669 B.n4 10.6151
R1874 B.n665 B.n4 10.6151
R1875 B.n665 B.n664 10.6151
R1876 B.n664 B.n663 10.6151
R1877 B.n663 B.n6 10.6151
R1878 B.n659 B.n6 10.6151
R1879 B.n659 B.n658 10.6151
R1880 B.n658 B.n657 10.6151
R1881 B.n657 B.n8 10.6151
R1882 B.n653 B.n8 10.6151
R1883 B.n653 B.n652 10.6151
R1884 B.n652 B.n651 10.6151
R1885 B.n651 B.n10 10.6151
R1886 B.n647 B.n10 10.6151
R1887 B.n647 B.n646 10.6151
R1888 B.n646 B.n645 10.6151
R1889 B.n645 B.n12 10.6151
R1890 B.n641 B.n12 10.6151
R1891 B.n641 B.n640 10.6151
R1892 B.n640 B.n639 10.6151
R1893 B.n639 B.n14 10.6151
R1894 B.n635 B.n14 10.6151
R1895 B.n635 B.n634 10.6151
R1896 B.n634 B.n633 10.6151
R1897 B.n633 B.n16 10.6151
R1898 B.n629 B.n16 10.6151
R1899 B.n629 B.n628 10.6151
R1900 B.n628 B.n627 10.6151
R1901 B.n627 B.n18 10.6151
R1902 B.n623 B.n18 10.6151
R1903 B.n623 B.n622 10.6151
R1904 B.n622 B.n621 10.6151
R1905 B.n621 B.n20 10.6151
R1906 B.n617 B.n20 10.6151
R1907 B.n617 B.n616 10.6151
R1908 B.n616 B.n615 10.6151
R1909 B.n556 B.n555 6.5566
R1910 B.n543 B.n542 6.5566
R1911 B.n292 B.n291 6.5566
R1912 B.n304 B.n130 6.5566
R1913 B.n557 B.n556 4.05904
R1914 B.n542 B.n541 4.05904
R1915 B.n291 B.n290 4.05904
R1916 B.n307 B.n130 4.05904
R1917 B.n675 B.n0 2.81026
R1918 B.n675 B.n1 2.81026
C0 B w_n3130_n3088# 8.543961f
C1 VP VDD2 0.437864f
C2 VTAIL VDD1 7.6054f
C3 VP VN 6.45841f
C4 VDD2 VN 7.13297f
C5 B VTAIL 4.16145f
C6 VP w_n3130_n3088# 6.52881f
C7 B VDD1 1.37764f
C8 w_n3130_n3088# VDD2 1.74483f
C9 w_n3130_n3088# VN 6.12474f
C10 VP VTAIL 7.34967f
C11 VTAIL VDD2 7.65465f
C12 VP VDD1 7.41936f
C13 VDD1 VDD2 1.37535f
C14 VTAIL VN 7.335569f
C15 VDD1 VN 0.150466f
C16 VP B 1.70593f
C17 B VDD2 1.44944f
C18 w_n3130_n3088# VTAIL 3.84503f
C19 w_n3130_n3088# VDD1 1.66243f
C20 B VN 1.03268f
C21 VDD2 VSUBS 1.556806f
C22 VDD1 VSUBS 2.065977f
C23 VTAIL VSUBS 1.136676f
C24 VN VSUBS 5.72305f
C25 VP VSUBS 2.755351f
C26 B VSUBS 4.023837f
C27 w_n3130_n3088# VSUBS 0.119253p
C28 B.n0 VSUBS 0.00466f
C29 B.n1 VSUBS 0.00466f
C30 B.n2 VSUBS 0.007369f
C31 B.n3 VSUBS 0.007369f
C32 B.n4 VSUBS 0.007369f
C33 B.n5 VSUBS 0.007369f
C34 B.n6 VSUBS 0.007369f
C35 B.n7 VSUBS 0.007369f
C36 B.n8 VSUBS 0.007369f
C37 B.n9 VSUBS 0.007369f
C38 B.n10 VSUBS 0.007369f
C39 B.n11 VSUBS 0.007369f
C40 B.n12 VSUBS 0.007369f
C41 B.n13 VSUBS 0.007369f
C42 B.n14 VSUBS 0.007369f
C43 B.n15 VSUBS 0.007369f
C44 B.n16 VSUBS 0.007369f
C45 B.n17 VSUBS 0.007369f
C46 B.n18 VSUBS 0.007369f
C47 B.n19 VSUBS 0.007369f
C48 B.n20 VSUBS 0.007369f
C49 B.n21 VSUBS 0.007369f
C50 B.n22 VSUBS 0.016471f
C51 B.n23 VSUBS 0.007369f
C52 B.n24 VSUBS 0.007369f
C53 B.n25 VSUBS 0.007369f
C54 B.n26 VSUBS 0.007369f
C55 B.n27 VSUBS 0.007369f
C56 B.n28 VSUBS 0.007369f
C57 B.n29 VSUBS 0.007369f
C58 B.n30 VSUBS 0.007369f
C59 B.n31 VSUBS 0.007369f
C60 B.n32 VSUBS 0.007369f
C61 B.n33 VSUBS 0.007369f
C62 B.n34 VSUBS 0.007369f
C63 B.n35 VSUBS 0.007369f
C64 B.n36 VSUBS 0.007369f
C65 B.n37 VSUBS 0.007369f
C66 B.n38 VSUBS 0.007369f
C67 B.n39 VSUBS 0.007369f
C68 B.n40 VSUBS 0.007369f
C69 B.n41 VSUBS 0.007369f
C70 B.t11 VSUBS 0.189672f
C71 B.t10 VSUBS 0.214288f
C72 B.t9 VSUBS 0.914567f
C73 B.n42 VSUBS 0.341301f
C74 B.n43 VSUBS 0.240952f
C75 B.n44 VSUBS 0.007369f
C76 B.n45 VSUBS 0.007369f
C77 B.n46 VSUBS 0.007369f
C78 B.n47 VSUBS 0.007369f
C79 B.t5 VSUBS 0.189675f
C80 B.t4 VSUBS 0.214291f
C81 B.t3 VSUBS 0.914567f
C82 B.n48 VSUBS 0.341298f
C83 B.n49 VSUBS 0.240949f
C84 B.n50 VSUBS 0.007369f
C85 B.n51 VSUBS 0.007369f
C86 B.n52 VSUBS 0.007369f
C87 B.n53 VSUBS 0.007369f
C88 B.n54 VSUBS 0.007369f
C89 B.n55 VSUBS 0.007369f
C90 B.n56 VSUBS 0.007369f
C91 B.n57 VSUBS 0.007369f
C92 B.n58 VSUBS 0.007369f
C93 B.n59 VSUBS 0.007369f
C94 B.n60 VSUBS 0.007369f
C95 B.n61 VSUBS 0.007369f
C96 B.n62 VSUBS 0.007369f
C97 B.n63 VSUBS 0.007369f
C98 B.n64 VSUBS 0.007369f
C99 B.n65 VSUBS 0.007369f
C100 B.n66 VSUBS 0.007369f
C101 B.n67 VSUBS 0.007369f
C102 B.n68 VSUBS 0.015486f
C103 B.n69 VSUBS 0.007369f
C104 B.n70 VSUBS 0.007369f
C105 B.n71 VSUBS 0.007369f
C106 B.n72 VSUBS 0.007369f
C107 B.n73 VSUBS 0.007369f
C108 B.n74 VSUBS 0.007369f
C109 B.n75 VSUBS 0.007369f
C110 B.n76 VSUBS 0.007369f
C111 B.n77 VSUBS 0.007369f
C112 B.n78 VSUBS 0.007369f
C113 B.n79 VSUBS 0.007369f
C114 B.n80 VSUBS 0.007369f
C115 B.n81 VSUBS 0.007369f
C116 B.n82 VSUBS 0.007369f
C117 B.n83 VSUBS 0.007369f
C118 B.n84 VSUBS 0.007369f
C119 B.n85 VSUBS 0.007369f
C120 B.n86 VSUBS 0.007369f
C121 B.n87 VSUBS 0.007369f
C122 B.n88 VSUBS 0.007369f
C123 B.n89 VSUBS 0.007369f
C124 B.n90 VSUBS 0.007369f
C125 B.n91 VSUBS 0.007369f
C126 B.n92 VSUBS 0.007369f
C127 B.n93 VSUBS 0.007369f
C128 B.n94 VSUBS 0.007369f
C129 B.n95 VSUBS 0.007369f
C130 B.n96 VSUBS 0.007369f
C131 B.n97 VSUBS 0.007369f
C132 B.n98 VSUBS 0.007369f
C133 B.n99 VSUBS 0.007369f
C134 B.n100 VSUBS 0.007369f
C135 B.n101 VSUBS 0.007369f
C136 B.n102 VSUBS 0.007369f
C137 B.n103 VSUBS 0.007369f
C138 B.n104 VSUBS 0.007369f
C139 B.n105 VSUBS 0.007369f
C140 B.n106 VSUBS 0.007369f
C141 B.n107 VSUBS 0.007369f
C142 B.n108 VSUBS 0.007369f
C143 B.n109 VSUBS 0.016471f
C144 B.n110 VSUBS 0.007369f
C145 B.n111 VSUBS 0.007369f
C146 B.n112 VSUBS 0.007369f
C147 B.n113 VSUBS 0.007369f
C148 B.n114 VSUBS 0.007369f
C149 B.n115 VSUBS 0.007369f
C150 B.n116 VSUBS 0.007369f
C151 B.n117 VSUBS 0.007369f
C152 B.n118 VSUBS 0.007369f
C153 B.n119 VSUBS 0.007369f
C154 B.n120 VSUBS 0.007369f
C155 B.n121 VSUBS 0.007369f
C156 B.n122 VSUBS 0.007369f
C157 B.n123 VSUBS 0.007369f
C158 B.n124 VSUBS 0.007369f
C159 B.n125 VSUBS 0.007369f
C160 B.n126 VSUBS 0.007369f
C161 B.n127 VSUBS 0.007369f
C162 B.t1 VSUBS 0.189675f
C163 B.t2 VSUBS 0.214291f
C164 B.t0 VSUBS 0.914567f
C165 B.n128 VSUBS 0.341298f
C166 B.n129 VSUBS 0.240949f
C167 B.n130 VSUBS 0.017074f
C168 B.n131 VSUBS 0.007369f
C169 B.n132 VSUBS 0.007369f
C170 B.n133 VSUBS 0.007369f
C171 B.n134 VSUBS 0.007369f
C172 B.n135 VSUBS 0.007369f
C173 B.t7 VSUBS 0.189672f
C174 B.t8 VSUBS 0.214288f
C175 B.t6 VSUBS 0.914567f
C176 B.n136 VSUBS 0.341301f
C177 B.n137 VSUBS 0.240952f
C178 B.n138 VSUBS 0.007369f
C179 B.n139 VSUBS 0.007369f
C180 B.n140 VSUBS 0.007369f
C181 B.n141 VSUBS 0.007369f
C182 B.n142 VSUBS 0.007369f
C183 B.n143 VSUBS 0.007369f
C184 B.n144 VSUBS 0.007369f
C185 B.n145 VSUBS 0.007369f
C186 B.n146 VSUBS 0.007369f
C187 B.n147 VSUBS 0.007369f
C188 B.n148 VSUBS 0.007369f
C189 B.n149 VSUBS 0.007369f
C190 B.n150 VSUBS 0.007369f
C191 B.n151 VSUBS 0.007369f
C192 B.n152 VSUBS 0.007369f
C193 B.n153 VSUBS 0.007369f
C194 B.n154 VSUBS 0.007369f
C195 B.n155 VSUBS 0.007369f
C196 B.n156 VSUBS 0.01539f
C197 B.n157 VSUBS 0.007369f
C198 B.n158 VSUBS 0.007369f
C199 B.n159 VSUBS 0.007369f
C200 B.n160 VSUBS 0.007369f
C201 B.n161 VSUBS 0.007369f
C202 B.n162 VSUBS 0.007369f
C203 B.n163 VSUBS 0.007369f
C204 B.n164 VSUBS 0.007369f
C205 B.n165 VSUBS 0.007369f
C206 B.n166 VSUBS 0.007369f
C207 B.n167 VSUBS 0.007369f
C208 B.n168 VSUBS 0.007369f
C209 B.n169 VSUBS 0.007369f
C210 B.n170 VSUBS 0.007369f
C211 B.n171 VSUBS 0.007369f
C212 B.n172 VSUBS 0.007369f
C213 B.n173 VSUBS 0.007369f
C214 B.n174 VSUBS 0.007369f
C215 B.n175 VSUBS 0.007369f
C216 B.n176 VSUBS 0.007369f
C217 B.n177 VSUBS 0.007369f
C218 B.n178 VSUBS 0.007369f
C219 B.n179 VSUBS 0.007369f
C220 B.n180 VSUBS 0.007369f
C221 B.n181 VSUBS 0.007369f
C222 B.n182 VSUBS 0.007369f
C223 B.n183 VSUBS 0.007369f
C224 B.n184 VSUBS 0.007369f
C225 B.n185 VSUBS 0.007369f
C226 B.n186 VSUBS 0.007369f
C227 B.n187 VSUBS 0.007369f
C228 B.n188 VSUBS 0.007369f
C229 B.n189 VSUBS 0.007369f
C230 B.n190 VSUBS 0.007369f
C231 B.n191 VSUBS 0.007369f
C232 B.n192 VSUBS 0.007369f
C233 B.n193 VSUBS 0.007369f
C234 B.n194 VSUBS 0.007369f
C235 B.n195 VSUBS 0.007369f
C236 B.n196 VSUBS 0.007369f
C237 B.n197 VSUBS 0.007369f
C238 B.n198 VSUBS 0.007369f
C239 B.n199 VSUBS 0.007369f
C240 B.n200 VSUBS 0.007369f
C241 B.n201 VSUBS 0.007369f
C242 B.n202 VSUBS 0.007369f
C243 B.n203 VSUBS 0.007369f
C244 B.n204 VSUBS 0.007369f
C245 B.n205 VSUBS 0.007369f
C246 B.n206 VSUBS 0.007369f
C247 B.n207 VSUBS 0.007369f
C248 B.n208 VSUBS 0.007369f
C249 B.n209 VSUBS 0.007369f
C250 B.n210 VSUBS 0.007369f
C251 B.n211 VSUBS 0.007369f
C252 B.n212 VSUBS 0.007369f
C253 B.n213 VSUBS 0.007369f
C254 B.n214 VSUBS 0.007369f
C255 B.n215 VSUBS 0.007369f
C256 B.n216 VSUBS 0.007369f
C257 B.n217 VSUBS 0.007369f
C258 B.n218 VSUBS 0.007369f
C259 B.n219 VSUBS 0.007369f
C260 B.n220 VSUBS 0.007369f
C261 B.n221 VSUBS 0.007369f
C262 B.n222 VSUBS 0.007369f
C263 B.n223 VSUBS 0.007369f
C264 B.n224 VSUBS 0.007369f
C265 B.n225 VSUBS 0.007369f
C266 B.n226 VSUBS 0.007369f
C267 B.n227 VSUBS 0.007369f
C268 B.n228 VSUBS 0.007369f
C269 B.n229 VSUBS 0.007369f
C270 B.n230 VSUBS 0.007369f
C271 B.n231 VSUBS 0.007369f
C272 B.n232 VSUBS 0.007369f
C273 B.n233 VSUBS 0.01539f
C274 B.n234 VSUBS 0.016471f
C275 B.n235 VSUBS 0.016471f
C276 B.n236 VSUBS 0.007369f
C277 B.n237 VSUBS 0.007369f
C278 B.n238 VSUBS 0.007369f
C279 B.n239 VSUBS 0.007369f
C280 B.n240 VSUBS 0.007369f
C281 B.n241 VSUBS 0.007369f
C282 B.n242 VSUBS 0.007369f
C283 B.n243 VSUBS 0.007369f
C284 B.n244 VSUBS 0.007369f
C285 B.n245 VSUBS 0.007369f
C286 B.n246 VSUBS 0.007369f
C287 B.n247 VSUBS 0.007369f
C288 B.n248 VSUBS 0.007369f
C289 B.n249 VSUBS 0.007369f
C290 B.n250 VSUBS 0.007369f
C291 B.n251 VSUBS 0.007369f
C292 B.n252 VSUBS 0.007369f
C293 B.n253 VSUBS 0.007369f
C294 B.n254 VSUBS 0.007369f
C295 B.n255 VSUBS 0.007369f
C296 B.n256 VSUBS 0.007369f
C297 B.n257 VSUBS 0.007369f
C298 B.n258 VSUBS 0.007369f
C299 B.n259 VSUBS 0.007369f
C300 B.n260 VSUBS 0.007369f
C301 B.n261 VSUBS 0.007369f
C302 B.n262 VSUBS 0.007369f
C303 B.n263 VSUBS 0.007369f
C304 B.n264 VSUBS 0.007369f
C305 B.n265 VSUBS 0.007369f
C306 B.n266 VSUBS 0.007369f
C307 B.n267 VSUBS 0.007369f
C308 B.n268 VSUBS 0.007369f
C309 B.n269 VSUBS 0.007369f
C310 B.n270 VSUBS 0.007369f
C311 B.n271 VSUBS 0.007369f
C312 B.n272 VSUBS 0.007369f
C313 B.n273 VSUBS 0.007369f
C314 B.n274 VSUBS 0.007369f
C315 B.n275 VSUBS 0.007369f
C316 B.n276 VSUBS 0.007369f
C317 B.n277 VSUBS 0.007369f
C318 B.n278 VSUBS 0.007369f
C319 B.n279 VSUBS 0.007369f
C320 B.n280 VSUBS 0.007369f
C321 B.n281 VSUBS 0.007369f
C322 B.n282 VSUBS 0.007369f
C323 B.n283 VSUBS 0.007369f
C324 B.n284 VSUBS 0.007369f
C325 B.n285 VSUBS 0.007369f
C326 B.n286 VSUBS 0.007369f
C327 B.n287 VSUBS 0.007369f
C328 B.n288 VSUBS 0.007369f
C329 B.n289 VSUBS 0.007369f
C330 B.n290 VSUBS 0.005093f
C331 B.n291 VSUBS 0.017074f
C332 B.n292 VSUBS 0.00596f
C333 B.n293 VSUBS 0.007369f
C334 B.n294 VSUBS 0.007369f
C335 B.n295 VSUBS 0.007369f
C336 B.n296 VSUBS 0.007369f
C337 B.n297 VSUBS 0.007369f
C338 B.n298 VSUBS 0.007369f
C339 B.n299 VSUBS 0.007369f
C340 B.n300 VSUBS 0.007369f
C341 B.n301 VSUBS 0.007369f
C342 B.n302 VSUBS 0.007369f
C343 B.n303 VSUBS 0.007369f
C344 B.n304 VSUBS 0.00596f
C345 B.n305 VSUBS 0.007369f
C346 B.n306 VSUBS 0.007369f
C347 B.n307 VSUBS 0.005093f
C348 B.n308 VSUBS 0.007369f
C349 B.n309 VSUBS 0.007369f
C350 B.n310 VSUBS 0.007369f
C351 B.n311 VSUBS 0.007369f
C352 B.n312 VSUBS 0.007369f
C353 B.n313 VSUBS 0.007369f
C354 B.n314 VSUBS 0.007369f
C355 B.n315 VSUBS 0.007369f
C356 B.n316 VSUBS 0.007369f
C357 B.n317 VSUBS 0.007369f
C358 B.n318 VSUBS 0.007369f
C359 B.n319 VSUBS 0.007369f
C360 B.n320 VSUBS 0.007369f
C361 B.n321 VSUBS 0.007369f
C362 B.n322 VSUBS 0.007369f
C363 B.n323 VSUBS 0.007369f
C364 B.n324 VSUBS 0.007369f
C365 B.n325 VSUBS 0.007369f
C366 B.n326 VSUBS 0.007369f
C367 B.n327 VSUBS 0.007369f
C368 B.n328 VSUBS 0.007369f
C369 B.n329 VSUBS 0.007369f
C370 B.n330 VSUBS 0.007369f
C371 B.n331 VSUBS 0.007369f
C372 B.n332 VSUBS 0.007369f
C373 B.n333 VSUBS 0.007369f
C374 B.n334 VSUBS 0.007369f
C375 B.n335 VSUBS 0.007369f
C376 B.n336 VSUBS 0.007369f
C377 B.n337 VSUBS 0.007369f
C378 B.n338 VSUBS 0.007369f
C379 B.n339 VSUBS 0.007369f
C380 B.n340 VSUBS 0.007369f
C381 B.n341 VSUBS 0.007369f
C382 B.n342 VSUBS 0.007369f
C383 B.n343 VSUBS 0.007369f
C384 B.n344 VSUBS 0.007369f
C385 B.n345 VSUBS 0.007369f
C386 B.n346 VSUBS 0.007369f
C387 B.n347 VSUBS 0.007369f
C388 B.n348 VSUBS 0.007369f
C389 B.n349 VSUBS 0.007369f
C390 B.n350 VSUBS 0.007369f
C391 B.n351 VSUBS 0.007369f
C392 B.n352 VSUBS 0.007369f
C393 B.n353 VSUBS 0.007369f
C394 B.n354 VSUBS 0.007369f
C395 B.n355 VSUBS 0.007369f
C396 B.n356 VSUBS 0.007369f
C397 B.n357 VSUBS 0.007369f
C398 B.n358 VSUBS 0.007369f
C399 B.n359 VSUBS 0.007369f
C400 B.n360 VSUBS 0.007369f
C401 B.n361 VSUBS 0.007369f
C402 B.n362 VSUBS 0.016471f
C403 B.n363 VSUBS 0.01539f
C404 B.n364 VSUBS 0.01539f
C405 B.n365 VSUBS 0.007369f
C406 B.n366 VSUBS 0.007369f
C407 B.n367 VSUBS 0.007369f
C408 B.n368 VSUBS 0.007369f
C409 B.n369 VSUBS 0.007369f
C410 B.n370 VSUBS 0.007369f
C411 B.n371 VSUBS 0.007369f
C412 B.n372 VSUBS 0.007369f
C413 B.n373 VSUBS 0.007369f
C414 B.n374 VSUBS 0.007369f
C415 B.n375 VSUBS 0.007369f
C416 B.n376 VSUBS 0.007369f
C417 B.n377 VSUBS 0.007369f
C418 B.n378 VSUBS 0.007369f
C419 B.n379 VSUBS 0.007369f
C420 B.n380 VSUBS 0.007369f
C421 B.n381 VSUBS 0.007369f
C422 B.n382 VSUBS 0.007369f
C423 B.n383 VSUBS 0.007369f
C424 B.n384 VSUBS 0.007369f
C425 B.n385 VSUBS 0.007369f
C426 B.n386 VSUBS 0.007369f
C427 B.n387 VSUBS 0.007369f
C428 B.n388 VSUBS 0.007369f
C429 B.n389 VSUBS 0.007369f
C430 B.n390 VSUBS 0.007369f
C431 B.n391 VSUBS 0.007369f
C432 B.n392 VSUBS 0.007369f
C433 B.n393 VSUBS 0.007369f
C434 B.n394 VSUBS 0.007369f
C435 B.n395 VSUBS 0.007369f
C436 B.n396 VSUBS 0.007369f
C437 B.n397 VSUBS 0.007369f
C438 B.n398 VSUBS 0.007369f
C439 B.n399 VSUBS 0.007369f
C440 B.n400 VSUBS 0.007369f
C441 B.n401 VSUBS 0.007369f
C442 B.n402 VSUBS 0.007369f
C443 B.n403 VSUBS 0.007369f
C444 B.n404 VSUBS 0.007369f
C445 B.n405 VSUBS 0.007369f
C446 B.n406 VSUBS 0.007369f
C447 B.n407 VSUBS 0.007369f
C448 B.n408 VSUBS 0.007369f
C449 B.n409 VSUBS 0.007369f
C450 B.n410 VSUBS 0.007369f
C451 B.n411 VSUBS 0.007369f
C452 B.n412 VSUBS 0.007369f
C453 B.n413 VSUBS 0.007369f
C454 B.n414 VSUBS 0.007369f
C455 B.n415 VSUBS 0.007369f
C456 B.n416 VSUBS 0.007369f
C457 B.n417 VSUBS 0.007369f
C458 B.n418 VSUBS 0.007369f
C459 B.n419 VSUBS 0.007369f
C460 B.n420 VSUBS 0.007369f
C461 B.n421 VSUBS 0.007369f
C462 B.n422 VSUBS 0.007369f
C463 B.n423 VSUBS 0.007369f
C464 B.n424 VSUBS 0.007369f
C465 B.n425 VSUBS 0.007369f
C466 B.n426 VSUBS 0.007369f
C467 B.n427 VSUBS 0.007369f
C468 B.n428 VSUBS 0.007369f
C469 B.n429 VSUBS 0.007369f
C470 B.n430 VSUBS 0.007369f
C471 B.n431 VSUBS 0.007369f
C472 B.n432 VSUBS 0.007369f
C473 B.n433 VSUBS 0.007369f
C474 B.n434 VSUBS 0.007369f
C475 B.n435 VSUBS 0.007369f
C476 B.n436 VSUBS 0.007369f
C477 B.n437 VSUBS 0.007369f
C478 B.n438 VSUBS 0.007369f
C479 B.n439 VSUBS 0.007369f
C480 B.n440 VSUBS 0.007369f
C481 B.n441 VSUBS 0.007369f
C482 B.n442 VSUBS 0.007369f
C483 B.n443 VSUBS 0.007369f
C484 B.n444 VSUBS 0.007369f
C485 B.n445 VSUBS 0.007369f
C486 B.n446 VSUBS 0.007369f
C487 B.n447 VSUBS 0.007369f
C488 B.n448 VSUBS 0.007369f
C489 B.n449 VSUBS 0.007369f
C490 B.n450 VSUBS 0.007369f
C491 B.n451 VSUBS 0.007369f
C492 B.n452 VSUBS 0.007369f
C493 B.n453 VSUBS 0.007369f
C494 B.n454 VSUBS 0.007369f
C495 B.n455 VSUBS 0.007369f
C496 B.n456 VSUBS 0.007369f
C497 B.n457 VSUBS 0.007369f
C498 B.n458 VSUBS 0.007369f
C499 B.n459 VSUBS 0.007369f
C500 B.n460 VSUBS 0.007369f
C501 B.n461 VSUBS 0.007369f
C502 B.n462 VSUBS 0.007369f
C503 B.n463 VSUBS 0.007369f
C504 B.n464 VSUBS 0.007369f
C505 B.n465 VSUBS 0.007369f
C506 B.n466 VSUBS 0.007369f
C507 B.n467 VSUBS 0.007369f
C508 B.n468 VSUBS 0.007369f
C509 B.n469 VSUBS 0.007369f
C510 B.n470 VSUBS 0.007369f
C511 B.n471 VSUBS 0.007369f
C512 B.n472 VSUBS 0.007369f
C513 B.n473 VSUBS 0.007369f
C514 B.n474 VSUBS 0.007369f
C515 B.n475 VSUBS 0.007369f
C516 B.n476 VSUBS 0.007369f
C517 B.n477 VSUBS 0.007369f
C518 B.n478 VSUBS 0.007369f
C519 B.n479 VSUBS 0.007369f
C520 B.n480 VSUBS 0.007369f
C521 B.n481 VSUBS 0.007369f
C522 B.n482 VSUBS 0.007369f
C523 B.n483 VSUBS 0.016375f
C524 B.n484 VSUBS 0.01539f
C525 B.n485 VSUBS 0.016471f
C526 B.n486 VSUBS 0.007369f
C527 B.n487 VSUBS 0.007369f
C528 B.n488 VSUBS 0.007369f
C529 B.n489 VSUBS 0.007369f
C530 B.n490 VSUBS 0.007369f
C531 B.n491 VSUBS 0.007369f
C532 B.n492 VSUBS 0.007369f
C533 B.n493 VSUBS 0.007369f
C534 B.n494 VSUBS 0.007369f
C535 B.n495 VSUBS 0.007369f
C536 B.n496 VSUBS 0.007369f
C537 B.n497 VSUBS 0.007369f
C538 B.n498 VSUBS 0.007369f
C539 B.n499 VSUBS 0.007369f
C540 B.n500 VSUBS 0.007369f
C541 B.n501 VSUBS 0.007369f
C542 B.n502 VSUBS 0.007369f
C543 B.n503 VSUBS 0.007369f
C544 B.n504 VSUBS 0.007369f
C545 B.n505 VSUBS 0.007369f
C546 B.n506 VSUBS 0.007369f
C547 B.n507 VSUBS 0.007369f
C548 B.n508 VSUBS 0.007369f
C549 B.n509 VSUBS 0.007369f
C550 B.n510 VSUBS 0.007369f
C551 B.n511 VSUBS 0.007369f
C552 B.n512 VSUBS 0.007369f
C553 B.n513 VSUBS 0.007369f
C554 B.n514 VSUBS 0.007369f
C555 B.n515 VSUBS 0.007369f
C556 B.n516 VSUBS 0.007369f
C557 B.n517 VSUBS 0.007369f
C558 B.n518 VSUBS 0.007369f
C559 B.n519 VSUBS 0.007369f
C560 B.n520 VSUBS 0.007369f
C561 B.n521 VSUBS 0.007369f
C562 B.n522 VSUBS 0.007369f
C563 B.n523 VSUBS 0.007369f
C564 B.n524 VSUBS 0.007369f
C565 B.n525 VSUBS 0.007369f
C566 B.n526 VSUBS 0.007369f
C567 B.n527 VSUBS 0.007369f
C568 B.n528 VSUBS 0.007369f
C569 B.n529 VSUBS 0.007369f
C570 B.n530 VSUBS 0.007369f
C571 B.n531 VSUBS 0.007369f
C572 B.n532 VSUBS 0.007369f
C573 B.n533 VSUBS 0.007369f
C574 B.n534 VSUBS 0.007369f
C575 B.n535 VSUBS 0.007369f
C576 B.n536 VSUBS 0.007369f
C577 B.n537 VSUBS 0.007369f
C578 B.n538 VSUBS 0.007369f
C579 B.n539 VSUBS 0.007369f
C580 B.n540 VSUBS 0.007369f
C581 B.n541 VSUBS 0.005093f
C582 B.n542 VSUBS 0.017074f
C583 B.n543 VSUBS 0.00596f
C584 B.n544 VSUBS 0.007369f
C585 B.n545 VSUBS 0.007369f
C586 B.n546 VSUBS 0.007369f
C587 B.n547 VSUBS 0.007369f
C588 B.n548 VSUBS 0.007369f
C589 B.n549 VSUBS 0.007369f
C590 B.n550 VSUBS 0.007369f
C591 B.n551 VSUBS 0.007369f
C592 B.n552 VSUBS 0.007369f
C593 B.n553 VSUBS 0.007369f
C594 B.n554 VSUBS 0.007369f
C595 B.n555 VSUBS 0.00596f
C596 B.n556 VSUBS 0.017074f
C597 B.n557 VSUBS 0.005093f
C598 B.n558 VSUBS 0.007369f
C599 B.n559 VSUBS 0.007369f
C600 B.n560 VSUBS 0.007369f
C601 B.n561 VSUBS 0.007369f
C602 B.n562 VSUBS 0.007369f
C603 B.n563 VSUBS 0.007369f
C604 B.n564 VSUBS 0.007369f
C605 B.n565 VSUBS 0.007369f
C606 B.n566 VSUBS 0.007369f
C607 B.n567 VSUBS 0.007369f
C608 B.n568 VSUBS 0.007369f
C609 B.n569 VSUBS 0.007369f
C610 B.n570 VSUBS 0.007369f
C611 B.n571 VSUBS 0.007369f
C612 B.n572 VSUBS 0.007369f
C613 B.n573 VSUBS 0.007369f
C614 B.n574 VSUBS 0.007369f
C615 B.n575 VSUBS 0.007369f
C616 B.n576 VSUBS 0.007369f
C617 B.n577 VSUBS 0.007369f
C618 B.n578 VSUBS 0.007369f
C619 B.n579 VSUBS 0.007369f
C620 B.n580 VSUBS 0.007369f
C621 B.n581 VSUBS 0.007369f
C622 B.n582 VSUBS 0.007369f
C623 B.n583 VSUBS 0.007369f
C624 B.n584 VSUBS 0.007369f
C625 B.n585 VSUBS 0.007369f
C626 B.n586 VSUBS 0.007369f
C627 B.n587 VSUBS 0.007369f
C628 B.n588 VSUBS 0.007369f
C629 B.n589 VSUBS 0.007369f
C630 B.n590 VSUBS 0.007369f
C631 B.n591 VSUBS 0.007369f
C632 B.n592 VSUBS 0.007369f
C633 B.n593 VSUBS 0.007369f
C634 B.n594 VSUBS 0.007369f
C635 B.n595 VSUBS 0.007369f
C636 B.n596 VSUBS 0.007369f
C637 B.n597 VSUBS 0.007369f
C638 B.n598 VSUBS 0.007369f
C639 B.n599 VSUBS 0.007369f
C640 B.n600 VSUBS 0.007369f
C641 B.n601 VSUBS 0.007369f
C642 B.n602 VSUBS 0.007369f
C643 B.n603 VSUBS 0.007369f
C644 B.n604 VSUBS 0.007369f
C645 B.n605 VSUBS 0.007369f
C646 B.n606 VSUBS 0.007369f
C647 B.n607 VSUBS 0.007369f
C648 B.n608 VSUBS 0.007369f
C649 B.n609 VSUBS 0.007369f
C650 B.n610 VSUBS 0.007369f
C651 B.n611 VSUBS 0.007369f
C652 B.n612 VSUBS 0.007369f
C653 B.n613 VSUBS 0.016471f
C654 B.n614 VSUBS 0.01539f
C655 B.n615 VSUBS 0.01539f
C656 B.n616 VSUBS 0.007369f
C657 B.n617 VSUBS 0.007369f
C658 B.n618 VSUBS 0.007369f
C659 B.n619 VSUBS 0.007369f
C660 B.n620 VSUBS 0.007369f
C661 B.n621 VSUBS 0.007369f
C662 B.n622 VSUBS 0.007369f
C663 B.n623 VSUBS 0.007369f
C664 B.n624 VSUBS 0.007369f
C665 B.n625 VSUBS 0.007369f
C666 B.n626 VSUBS 0.007369f
C667 B.n627 VSUBS 0.007369f
C668 B.n628 VSUBS 0.007369f
C669 B.n629 VSUBS 0.007369f
C670 B.n630 VSUBS 0.007369f
C671 B.n631 VSUBS 0.007369f
C672 B.n632 VSUBS 0.007369f
C673 B.n633 VSUBS 0.007369f
C674 B.n634 VSUBS 0.007369f
C675 B.n635 VSUBS 0.007369f
C676 B.n636 VSUBS 0.007369f
C677 B.n637 VSUBS 0.007369f
C678 B.n638 VSUBS 0.007369f
C679 B.n639 VSUBS 0.007369f
C680 B.n640 VSUBS 0.007369f
C681 B.n641 VSUBS 0.007369f
C682 B.n642 VSUBS 0.007369f
C683 B.n643 VSUBS 0.007369f
C684 B.n644 VSUBS 0.007369f
C685 B.n645 VSUBS 0.007369f
C686 B.n646 VSUBS 0.007369f
C687 B.n647 VSUBS 0.007369f
C688 B.n648 VSUBS 0.007369f
C689 B.n649 VSUBS 0.007369f
C690 B.n650 VSUBS 0.007369f
C691 B.n651 VSUBS 0.007369f
C692 B.n652 VSUBS 0.007369f
C693 B.n653 VSUBS 0.007369f
C694 B.n654 VSUBS 0.007369f
C695 B.n655 VSUBS 0.007369f
C696 B.n656 VSUBS 0.007369f
C697 B.n657 VSUBS 0.007369f
C698 B.n658 VSUBS 0.007369f
C699 B.n659 VSUBS 0.007369f
C700 B.n660 VSUBS 0.007369f
C701 B.n661 VSUBS 0.007369f
C702 B.n662 VSUBS 0.007369f
C703 B.n663 VSUBS 0.007369f
C704 B.n664 VSUBS 0.007369f
C705 B.n665 VSUBS 0.007369f
C706 B.n666 VSUBS 0.007369f
C707 B.n667 VSUBS 0.007369f
C708 B.n668 VSUBS 0.007369f
C709 B.n669 VSUBS 0.007369f
C710 B.n670 VSUBS 0.007369f
C711 B.n671 VSUBS 0.007369f
C712 B.n672 VSUBS 0.007369f
C713 B.n673 VSUBS 0.007369f
C714 B.n674 VSUBS 0.007369f
C715 B.n675 VSUBS 0.016686f
C716 VDD2.t1 VSUBS 0.206698f
C717 VDD2.t7 VSUBS 0.206698f
C718 VDD2.n0 VSUBS 1.58056f
C719 VDD2.t6 VSUBS 0.206698f
C720 VDD2.t2 VSUBS 0.206698f
C721 VDD2.n1 VSUBS 1.58056f
C722 VDD2.n2 VSUBS 3.21246f
C723 VDD2.t0 VSUBS 0.206698f
C724 VDD2.t4 VSUBS 0.206698f
C725 VDD2.n3 VSUBS 1.57259f
C726 VDD2.n4 VSUBS 2.79525f
C727 VDD2.t3 VSUBS 0.206698f
C728 VDD2.t5 VSUBS 0.206698f
C729 VDD2.n5 VSUBS 1.58052f
C730 VN.n0 VSUBS 0.047368f
C731 VN.t5 VSUBS 1.89182f
C732 VN.n1 VSUBS 0.066299f
C733 VN.n2 VSUBS 0.03593f
C734 VN.t1 VSUBS 1.89182f
C735 VN.n3 VSUBS 0.05223f
C736 VN.t6 VSUBS 2.04966f
C737 VN.n4 VSUBS 0.772145f
C738 VN.t0 VSUBS 1.89182f
C739 VN.n5 VSUBS 0.769645f
C740 VN.n6 VSUBS 0.055445f
C741 VN.n7 VSUBS 0.263467f
C742 VN.n8 VSUBS 0.03593f
C743 VN.n9 VSUBS 0.03593f
C744 VN.n10 VSUBS 0.05223f
C745 VN.n11 VSUBS 0.055445f
C746 VN.n12 VSUBS 0.683975f
C747 VN.n13 VSUBS 0.04492f
C748 VN.n14 VSUBS 0.03593f
C749 VN.n15 VSUBS 0.03593f
C750 VN.n16 VSUBS 0.03593f
C751 VN.n17 VSUBS 0.032909f
C752 VN.n18 VSUBS 0.071223f
C753 VN.n19 VSUBS 0.793256f
C754 VN.n20 VSUBS 0.038271f
C755 VN.n21 VSUBS 0.047368f
C756 VN.t7 VSUBS 1.89182f
C757 VN.n22 VSUBS 0.066299f
C758 VN.n23 VSUBS 0.03593f
C759 VN.t3 VSUBS 1.89182f
C760 VN.n24 VSUBS 0.05223f
C761 VN.t2 VSUBS 2.04966f
C762 VN.n25 VSUBS 0.772145f
C763 VN.t4 VSUBS 1.89182f
C764 VN.n26 VSUBS 0.769645f
C765 VN.n27 VSUBS 0.055445f
C766 VN.n28 VSUBS 0.263467f
C767 VN.n29 VSUBS 0.03593f
C768 VN.n30 VSUBS 0.03593f
C769 VN.n31 VSUBS 0.05223f
C770 VN.n32 VSUBS 0.055445f
C771 VN.n33 VSUBS 0.683975f
C772 VN.n34 VSUBS 0.04492f
C773 VN.n35 VSUBS 0.03593f
C774 VN.n36 VSUBS 0.03593f
C775 VN.n37 VSUBS 0.03593f
C776 VN.n38 VSUBS 0.032909f
C777 VN.n39 VSUBS 0.071223f
C778 VN.n40 VSUBS 0.793256f
C779 VN.n41 VSUBS 1.77904f
C780 VTAIL.t3 VSUBS 0.209052f
C781 VTAIL.t1 VSUBS 0.209052f
C782 VTAIL.n0 VSUBS 1.45812f
C783 VTAIL.n1 VSUBS 0.715051f
C784 VTAIL.n2 VSUBS 0.025626f
C785 VTAIL.n3 VSUBS 0.024957f
C786 VTAIL.n4 VSUBS 0.013411f
C787 VTAIL.n5 VSUBS 0.031699f
C788 VTAIL.n6 VSUBS 0.0142f
C789 VTAIL.n7 VSUBS 0.024957f
C790 VTAIL.n8 VSUBS 0.013411f
C791 VTAIL.n9 VSUBS 0.031699f
C792 VTAIL.n10 VSUBS 0.0142f
C793 VTAIL.n11 VSUBS 0.024957f
C794 VTAIL.n12 VSUBS 0.013411f
C795 VTAIL.n13 VSUBS 0.031699f
C796 VTAIL.n14 VSUBS 0.0142f
C797 VTAIL.n15 VSUBS 0.024957f
C798 VTAIL.n16 VSUBS 0.013411f
C799 VTAIL.n17 VSUBS 0.031699f
C800 VTAIL.n18 VSUBS 0.0142f
C801 VTAIL.n19 VSUBS 0.180759f
C802 VTAIL.t7 VSUBS 0.068194f
C803 VTAIL.n20 VSUBS 0.023774f
C804 VTAIL.n21 VSUBS 0.023845f
C805 VTAIL.n22 VSUBS 0.013411f
C806 VTAIL.n23 VSUBS 1.07312f
C807 VTAIL.n24 VSUBS 0.024957f
C808 VTAIL.n25 VSUBS 0.013411f
C809 VTAIL.n26 VSUBS 0.0142f
C810 VTAIL.n27 VSUBS 0.031699f
C811 VTAIL.n28 VSUBS 0.031699f
C812 VTAIL.n29 VSUBS 0.0142f
C813 VTAIL.n30 VSUBS 0.013411f
C814 VTAIL.n31 VSUBS 0.024957f
C815 VTAIL.n32 VSUBS 0.024957f
C816 VTAIL.n33 VSUBS 0.013411f
C817 VTAIL.n34 VSUBS 0.0142f
C818 VTAIL.n35 VSUBS 0.031699f
C819 VTAIL.n36 VSUBS 0.031699f
C820 VTAIL.n37 VSUBS 0.031699f
C821 VTAIL.n38 VSUBS 0.0142f
C822 VTAIL.n39 VSUBS 0.013411f
C823 VTAIL.n40 VSUBS 0.024957f
C824 VTAIL.n41 VSUBS 0.024957f
C825 VTAIL.n42 VSUBS 0.013411f
C826 VTAIL.n43 VSUBS 0.013805f
C827 VTAIL.n44 VSUBS 0.013805f
C828 VTAIL.n45 VSUBS 0.031699f
C829 VTAIL.n46 VSUBS 0.031699f
C830 VTAIL.n47 VSUBS 0.0142f
C831 VTAIL.n48 VSUBS 0.013411f
C832 VTAIL.n49 VSUBS 0.024957f
C833 VTAIL.n50 VSUBS 0.024957f
C834 VTAIL.n51 VSUBS 0.013411f
C835 VTAIL.n52 VSUBS 0.0142f
C836 VTAIL.n53 VSUBS 0.031699f
C837 VTAIL.n54 VSUBS 0.070618f
C838 VTAIL.n55 VSUBS 0.0142f
C839 VTAIL.n56 VSUBS 0.013411f
C840 VTAIL.n57 VSUBS 0.05496f
C841 VTAIL.n58 VSUBS 0.035155f
C842 VTAIL.n59 VSUBS 0.207303f
C843 VTAIL.n60 VSUBS 0.025626f
C844 VTAIL.n61 VSUBS 0.024957f
C845 VTAIL.n62 VSUBS 0.013411f
C846 VTAIL.n63 VSUBS 0.031699f
C847 VTAIL.n64 VSUBS 0.0142f
C848 VTAIL.n65 VSUBS 0.024957f
C849 VTAIL.n66 VSUBS 0.013411f
C850 VTAIL.n67 VSUBS 0.031699f
C851 VTAIL.n68 VSUBS 0.0142f
C852 VTAIL.n69 VSUBS 0.024957f
C853 VTAIL.n70 VSUBS 0.013411f
C854 VTAIL.n71 VSUBS 0.031699f
C855 VTAIL.n72 VSUBS 0.0142f
C856 VTAIL.n73 VSUBS 0.024957f
C857 VTAIL.n74 VSUBS 0.013411f
C858 VTAIL.n75 VSUBS 0.031699f
C859 VTAIL.n76 VSUBS 0.0142f
C860 VTAIL.n77 VSUBS 0.180759f
C861 VTAIL.t10 VSUBS 0.068194f
C862 VTAIL.n78 VSUBS 0.023774f
C863 VTAIL.n79 VSUBS 0.023845f
C864 VTAIL.n80 VSUBS 0.013411f
C865 VTAIL.n81 VSUBS 1.07312f
C866 VTAIL.n82 VSUBS 0.024957f
C867 VTAIL.n83 VSUBS 0.013411f
C868 VTAIL.n84 VSUBS 0.0142f
C869 VTAIL.n85 VSUBS 0.031699f
C870 VTAIL.n86 VSUBS 0.031699f
C871 VTAIL.n87 VSUBS 0.0142f
C872 VTAIL.n88 VSUBS 0.013411f
C873 VTAIL.n89 VSUBS 0.024957f
C874 VTAIL.n90 VSUBS 0.024957f
C875 VTAIL.n91 VSUBS 0.013411f
C876 VTAIL.n92 VSUBS 0.0142f
C877 VTAIL.n93 VSUBS 0.031699f
C878 VTAIL.n94 VSUBS 0.031699f
C879 VTAIL.n95 VSUBS 0.031699f
C880 VTAIL.n96 VSUBS 0.0142f
C881 VTAIL.n97 VSUBS 0.013411f
C882 VTAIL.n98 VSUBS 0.024957f
C883 VTAIL.n99 VSUBS 0.024957f
C884 VTAIL.n100 VSUBS 0.013411f
C885 VTAIL.n101 VSUBS 0.013805f
C886 VTAIL.n102 VSUBS 0.013805f
C887 VTAIL.n103 VSUBS 0.031699f
C888 VTAIL.n104 VSUBS 0.031699f
C889 VTAIL.n105 VSUBS 0.0142f
C890 VTAIL.n106 VSUBS 0.013411f
C891 VTAIL.n107 VSUBS 0.024957f
C892 VTAIL.n108 VSUBS 0.024957f
C893 VTAIL.n109 VSUBS 0.013411f
C894 VTAIL.n110 VSUBS 0.0142f
C895 VTAIL.n111 VSUBS 0.031699f
C896 VTAIL.n112 VSUBS 0.070618f
C897 VTAIL.n113 VSUBS 0.0142f
C898 VTAIL.n114 VSUBS 0.013411f
C899 VTAIL.n115 VSUBS 0.05496f
C900 VTAIL.n116 VSUBS 0.035155f
C901 VTAIL.n117 VSUBS 0.207303f
C902 VTAIL.t13 VSUBS 0.209052f
C903 VTAIL.t15 VSUBS 0.209052f
C904 VTAIL.n118 VSUBS 1.45812f
C905 VTAIL.n119 VSUBS 0.860115f
C906 VTAIL.n120 VSUBS 0.025626f
C907 VTAIL.n121 VSUBS 0.024957f
C908 VTAIL.n122 VSUBS 0.013411f
C909 VTAIL.n123 VSUBS 0.031699f
C910 VTAIL.n124 VSUBS 0.0142f
C911 VTAIL.n125 VSUBS 0.024957f
C912 VTAIL.n126 VSUBS 0.013411f
C913 VTAIL.n127 VSUBS 0.031699f
C914 VTAIL.n128 VSUBS 0.0142f
C915 VTAIL.n129 VSUBS 0.024957f
C916 VTAIL.n130 VSUBS 0.013411f
C917 VTAIL.n131 VSUBS 0.031699f
C918 VTAIL.n132 VSUBS 0.0142f
C919 VTAIL.n133 VSUBS 0.024957f
C920 VTAIL.n134 VSUBS 0.013411f
C921 VTAIL.n135 VSUBS 0.031699f
C922 VTAIL.n136 VSUBS 0.0142f
C923 VTAIL.n137 VSUBS 0.180759f
C924 VTAIL.t9 VSUBS 0.068194f
C925 VTAIL.n138 VSUBS 0.023774f
C926 VTAIL.n139 VSUBS 0.023845f
C927 VTAIL.n140 VSUBS 0.013411f
C928 VTAIL.n141 VSUBS 1.07312f
C929 VTAIL.n142 VSUBS 0.024957f
C930 VTAIL.n143 VSUBS 0.013411f
C931 VTAIL.n144 VSUBS 0.0142f
C932 VTAIL.n145 VSUBS 0.031699f
C933 VTAIL.n146 VSUBS 0.031699f
C934 VTAIL.n147 VSUBS 0.0142f
C935 VTAIL.n148 VSUBS 0.013411f
C936 VTAIL.n149 VSUBS 0.024957f
C937 VTAIL.n150 VSUBS 0.024957f
C938 VTAIL.n151 VSUBS 0.013411f
C939 VTAIL.n152 VSUBS 0.0142f
C940 VTAIL.n153 VSUBS 0.031699f
C941 VTAIL.n154 VSUBS 0.031699f
C942 VTAIL.n155 VSUBS 0.031699f
C943 VTAIL.n156 VSUBS 0.0142f
C944 VTAIL.n157 VSUBS 0.013411f
C945 VTAIL.n158 VSUBS 0.024957f
C946 VTAIL.n159 VSUBS 0.024957f
C947 VTAIL.n160 VSUBS 0.013411f
C948 VTAIL.n161 VSUBS 0.013805f
C949 VTAIL.n162 VSUBS 0.013805f
C950 VTAIL.n163 VSUBS 0.031699f
C951 VTAIL.n164 VSUBS 0.031699f
C952 VTAIL.n165 VSUBS 0.0142f
C953 VTAIL.n166 VSUBS 0.013411f
C954 VTAIL.n167 VSUBS 0.024957f
C955 VTAIL.n168 VSUBS 0.024957f
C956 VTAIL.n169 VSUBS 0.013411f
C957 VTAIL.n170 VSUBS 0.0142f
C958 VTAIL.n171 VSUBS 0.031699f
C959 VTAIL.n172 VSUBS 0.070618f
C960 VTAIL.n173 VSUBS 0.0142f
C961 VTAIL.n174 VSUBS 0.013411f
C962 VTAIL.n175 VSUBS 0.05496f
C963 VTAIL.n176 VSUBS 0.035155f
C964 VTAIL.n177 VSUBS 1.39313f
C965 VTAIL.n178 VSUBS 0.025626f
C966 VTAIL.n179 VSUBS 0.024957f
C967 VTAIL.n180 VSUBS 0.013411f
C968 VTAIL.n181 VSUBS 0.031699f
C969 VTAIL.n182 VSUBS 0.0142f
C970 VTAIL.n183 VSUBS 0.024957f
C971 VTAIL.n184 VSUBS 0.013411f
C972 VTAIL.n185 VSUBS 0.031699f
C973 VTAIL.n186 VSUBS 0.0142f
C974 VTAIL.n187 VSUBS 0.024957f
C975 VTAIL.n188 VSUBS 0.013411f
C976 VTAIL.n189 VSUBS 0.031699f
C977 VTAIL.n190 VSUBS 0.031699f
C978 VTAIL.n191 VSUBS 0.0142f
C979 VTAIL.n192 VSUBS 0.024957f
C980 VTAIL.n193 VSUBS 0.013411f
C981 VTAIL.n194 VSUBS 0.031699f
C982 VTAIL.n195 VSUBS 0.0142f
C983 VTAIL.n196 VSUBS 0.180759f
C984 VTAIL.t2 VSUBS 0.068194f
C985 VTAIL.n197 VSUBS 0.023774f
C986 VTAIL.n198 VSUBS 0.023845f
C987 VTAIL.n199 VSUBS 0.013411f
C988 VTAIL.n200 VSUBS 1.07312f
C989 VTAIL.n201 VSUBS 0.024957f
C990 VTAIL.n202 VSUBS 0.013411f
C991 VTAIL.n203 VSUBS 0.0142f
C992 VTAIL.n204 VSUBS 0.031699f
C993 VTAIL.n205 VSUBS 0.031699f
C994 VTAIL.n206 VSUBS 0.0142f
C995 VTAIL.n207 VSUBS 0.013411f
C996 VTAIL.n208 VSUBS 0.024957f
C997 VTAIL.n209 VSUBS 0.024957f
C998 VTAIL.n210 VSUBS 0.013411f
C999 VTAIL.n211 VSUBS 0.0142f
C1000 VTAIL.n212 VSUBS 0.031699f
C1001 VTAIL.n213 VSUBS 0.031699f
C1002 VTAIL.n214 VSUBS 0.0142f
C1003 VTAIL.n215 VSUBS 0.013411f
C1004 VTAIL.n216 VSUBS 0.024957f
C1005 VTAIL.n217 VSUBS 0.024957f
C1006 VTAIL.n218 VSUBS 0.013411f
C1007 VTAIL.n219 VSUBS 0.013805f
C1008 VTAIL.n220 VSUBS 0.013805f
C1009 VTAIL.n221 VSUBS 0.031699f
C1010 VTAIL.n222 VSUBS 0.031699f
C1011 VTAIL.n223 VSUBS 0.0142f
C1012 VTAIL.n224 VSUBS 0.013411f
C1013 VTAIL.n225 VSUBS 0.024957f
C1014 VTAIL.n226 VSUBS 0.024957f
C1015 VTAIL.n227 VSUBS 0.013411f
C1016 VTAIL.n228 VSUBS 0.0142f
C1017 VTAIL.n229 VSUBS 0.031699f
C1018 VTAIL.n230 VSUBS 0.070618f
C1019 VTAIL.n231 VSUBS 0.0142f
C1020 VTAIL.n232 VSUBS 0.013411f
C1021 VTAIL.n233 VSUBS 0.05496f
C1022 VTAIL.n234 VSUBS 0.035155f
C1023 VTAIL.n235 VSUBS 1.39313f
C1024 VTAIL.t5 VSUBS 0.209052f
C1025 VTAIL.t6 VSUBS 0.209052f
C1026 VTAIL.n236 VSUBS 1.45813f
C1027 VTAIL.n237 VSUBS 0.860104f
C1028 VTAIL.n238 VSUBS 0.025626f
C1029 VTAIL.n239 VSUBS 0.024957f
C1030 VTAIL.n240 VSUBS 0.013411f
C1031 VTAIL.n241 VSUBS 0.031699f
C1032 VTAIL.n242 VSUBS 0.0142f
C1033 VTAIL.n243 VSUBS 0.024957f
C1034 VTAIL.n244 VSUBS 0.013411f
C1035 VTAIL.n245 VSUBS 0.031699f
C1036 VTAIL.n246 VSUBS 0.0142f
C1037 VTAIL.n247 VSUBS 0.024957f
C1038 VTAIL.n248 VSUBS 0.013411f
C1039 VTAIL.n249 VSUBS 0.031699f
C1040 VTAIL.n250 VSUBS 0.031699f
C1041 VTAIL.n251 VSUBS 0.0142f
C1042 VTAIL.n252 VSUBS 0.024957f
C1043 VTAIL.n253 VSUBS 0.013411f
C1044 VTAIL.n254 VSUBS 0.031699f
C1045 VTAIL.n255 VSUBS 0.0142f
C1046 VTAIL.n256 VSUBS 0.180759f
C1047 VTAIL.t4 VSUBS 0.068194f
C1048 VTAIL.n257 VSUBS 0.023774f
C1049 VTAIL.n258 VSUBS 0.023845f
C1050 VTAIL.n259 VSUBS 0.013411f
C1051 VTAIL.n260 VSUBS 1.07312f
C1052 VTAIL.n261 VSUBS 0.024957f
C1053 VTAIL.n262 VSUBS 0.013411f
C1054 VTAIL.n263 VSUBS 0.0142f
C1055 VTAIL.n264 VSUBS 0.031699f
C1056 VTAIL.n265 VSUBS 0.031699f
C1057 VTAIL.n266 VSUBS 0.0142f
C1058 VTAIL.n267 VSUBS 0.013411f
C1059 VTAIL.n268 VSUBS 0.024957f
C1060 VTAIL.n269 VSUBS 0.024957f
C1061 VTAIL.n270 VSUBS 0.013411f
C1062 VTAIL.n271 VSUBS 0.0142f
C1063 VTAIL.n272 VSUBS 0.031699f
C1064 VTAIL.n273 VSUBS 0.031699f
C1065 VTAIL.n274 VSUBS 0.0142f
C1066 VTAIL.n275 VSUBS 0.013411f
C1067 VTAIL.n276 VSUBS 0.024957f
C1068 VTAIL.n277 VSUBS 0.024957f
C1069 VTAIL.n278 VSUBS 0.013411f
C1070 VTAIL.n279 VSUBS 0.013805f
C1071 VTAIL.n280 VSUBS 0.013805f
C1072 VTAIL.n281 VSUBS 0.031699f
C1073 VTAIL.n282 VSUBS 0.031699f
C1074 VTAIL.n283 VSUBS 0.0142f
C1075 VTAIL.n284 VSUBS 0.013411f
C1076 VTAIL.n285 VSUBS 0.024957f
C1077 VTAIL.n286 VSUBS 0.024957f
C1078 VTAIL.n287 VSUBS 0.013411f
C1079 VTAIL.n288 VSUBS 0.0142f
C1080 VTAIL.n289 VSUBS 0.031699f
C1081 VTAIL.n290 VSUBS 0.070618f
C1082 VTAIL.n291 VSUBS 0.0142f
C1083 VTAIL.n292 VSUBS 0.013411f
C1084 VTAIL.n293 VSUBS 0.05496f
C1085 VTAIL.n294 VSUBS 0.035155f
C1086 VTAIL.n295 VSUBS 0.207303f
C1087 VTAIL.n296 VSUBS 0.025626f
C1088 VTAIL.n297 VSUBS 0.024957f
C1089 VTAIL.n298 VSUBS 0.013411f
C1090 VTAIL.n299 VSUBS 0.031699f
C1091 VTAIL.n300 VSUBS 0.0142f
C1092 VTAIL.n301 VSUBS 0.024957f
C1093 VTAIL.n302 VSUBS 0.013411f
C1094 VTAIL.n303 VSUBS 0.031699f
C1095 VTAIL.n304 VSUBS 0.0142f
C1096 VTAIL.n305 VSUBS 0.024957f
C1097 VTAIL.n306 VSUBS 0.013411f
C1098 VTAIL.n307 VSUBS 0.031699f
C1099 VTAIL.n308 VSUBS 0.031699f
C1100 VTAIL.n309 VSUBS 0.0142f
C1101 VTAIL.n310 VSUBS 0.024957f
C1102 VTAIL.n311 VSUBS 0.013411f
C1103 VTAIL.n312 VSUBS 0.031699f
C1104 VTAIL.n313 VSUBS 0.0142f
C1105 VTAIL.n314 VSUBS 0.180759f
C1106 VTAIL.t14 VSUBS 0.068194f
C1107 VTAIL.n315 VSUBS 0.023774f
C1108 VTAIL.n316 VSUBS 0.023845f
C1109 VTAIL.n317 VSUBS 0.013411f
C1110 VTAIL.n318 VSUBS 1.07312f
C1111 VTAIL.n319 VSUBS 0.024957f
C1112 VTAIL.n320 VSUBS 0.013411f
C1113 VTAIL.n321 VSUBS 0.0142f
C1114 VTAIL.n322 VSUBS 0.031699f
C1115 VTAIL.n323 VSUBS 0.031699f
C1116 VTAIL.n324 VSUBS 0.0142f
C1117 VTAIL.n325 VSUBS 0.013411f
C1118 VTAIL.n326 VSUBS 0.024957f
C1119 VTAIL.n327 VSUBS 0.024957f
C1120 VTAIL.n328 VSUBS 0.013411f
C1121 VTAIL.n329 VSUBS 0.0142f
C1122 VTAIL.n330 VSUBS 0.031699f
C1123 VTAIL.n331 VSUBS 0.031699f
C1124 VTAIL.n332 VSUBS 0.0142f
C1125 VTAIL.n333 VSUBS 0.013411f
C1126 VTAIL.n334 VSUBS 0.024957f
C1127 VTAIL.n335 VSUBS 0.024957f
C1128 VTAIL.n336 VSUBS 0.013411f
C1129 VTAIL.n337 VSUBS 0.013805f
C1130 VTAIL.n338 VSUBS 0.013805f
C1131 VTAIL.n339 VSUBS 0.031699f
C1132 VTAIL.n340 VSUBS 0.031699f
C1133 VTAIL.n341 VSUBS 0.0142f
C1134 VTAIL.n342 VSUBS 0.013411f
C1135 VTAIL.n343 VSUBS 0.024957f
C1136 VTAIL.n344 VSUBS 0.024957f
C1137 VTAIL.n345 VSUBS 0.013411f
C1138 VTAIL.n346 VSUBS 0.0142f
C1139 VTAIL.n347 VSUBS 0.031699f
C1140 VTAIL.n348 VSUBS 0.070618f
C1141 VTAIL.n349 VSUBS 0.0142f
C1142 VTAIL.n350 VSUBS 0.013411f
C1143 VTAIL.n351 VSUBS 0.05496f
C1144 VTAIL.n352 VSUBS 0.035155f
C1145 VTAIL.n353 VSUBS 0.207303f
C1146 VTAIL.t11 VSUBS 0.209052f
C1147 VTAIL.t8 VSUBS 0.209052f
C1148 VTAIL.n354 VSUBS 1.45813f
C1149 VTAIL.n355 VSUBS 0.860104f
C1150 VTAIL.n356 VSUBS 0.025626f
C1151 VTAIL.n357 VSUBS 0.024957f
C1152 VTAIL.n358 VSUBS 0.013411f
C1153 VTAIL.n359 VSUBS 0.031699f
C1154 VTAIL.n360 VSUBS 0.0142f
C1155 VTAIL.n361 VSUBS 0.024957f
C1156 VTAIL.n362 VSUBS 0.013411f
C1157 VTAIL.n363 VSUBS 0.031699f
C1158 VTAIL.n364 VSUBS 0.0142f
C1159 VTAIL.n365 VSUBS 0.024957f
C1160 VTAIL.n366 VSUBS 0.013411f
C1161 VTAIL.n367 VSUBS 0.031699f
C1162 VTAIL.n368 VSUBS 0.031699f
C1163 VTAIL.n369 VSUBS 0.0142f
C1164 VTAIL.n370 VSUBS 0.024957f
C1165 VTAIL.n371 VSUBS 0.013411f
C1166 VTAIL.n372 VSUBS 0.031699f
C1167 VTAIL.n373 VSUBS 0.0142f
C1168 VTAIL.n374 VSUBS 0.180759f
C1169 VTAIL.t12 VSUBS 0.068194f
C1170 VTAIL.n375 VSUBS 0.023774f
C1171 VTAIL.n376 VSUBS 0.023845f
C1172 VTAIL.n377 VSUBS 0.013411f
C1173 VTAIL.n378 VSUBS 1.07312f
C1174 VTAIL.n379 VSUBS 0.024957f
C1175 VTAIL.n380 VSUBS 0.013411f
C1176 VTAIL.n381 VSUBS 0.0142f
C1177 VTAIL.n382 VSUBS 0.031699f
C1178 VTAIL.n383 VSUBS 0.031699f
C1179 VTAIL.n384 VSUBS 0.0142f
C1180 VTAIL.n385 VSUBS 0.013411f
C1181 VTAIL.n386 VSUBS 0.024957f
C1182 VTAIL.n387 VSUBS 0.024957f
C1183 VTAIL.n388 VSUBS 0.013411f
C1184 VTAIL.n389 VSUBS 0.0142f
C1185 VTAIL.n390 VSUBS 0.031699f
C1186 VTAIL.n391 VSUBS 0.031699f
C1187 VTAIL.n392 VSUBS 0.0142f
C1188 VTAIL.n393 VSUBS 0.013411f
C1189 VTAIL.n394 VSUBS 0.024957f
C1190 VTAIL.n395 VSUBS 0.024957f
C1191 VTAIL.n396 VSUBS 0.013411f
C1192 VTAIL.n397 VSUBS 0.013805f
C1193 VTAIL.n398 VSUBS 0.013805f
C1194 VTAIL.n399 VSUBS 0.031699f
C1195 VTAIL.n400 VSUBS 0.031699f
C1196 VTAIL.n401 VSUBS 0.0142f
C1197 VTAIL.n402 VSUBS 0.013411f
C1198 VTAIL.n403 VSUBS 0.024957f
C1199 VTAIL.n404 VSUBS 0.024957f
C1200 VTAIL.n405 VSUBS 0.013411f
C1201 VTAIL.n406 VSUBS 0.0142f
C1202 VTAIL.n407 VSUBS 0.031699f
C1203 VTAIL.n408 VSUBS 0.070618f
C1204 VTAIL.n409 VSUBS 0.0142f
C1205 VTAIL.n410 VSUBS 0.013411f
C1206 VTAIL.n411 VSUBS 0.05496f
C1207 VTAIL.n412 VSUBS 0.035155f
C1208 VTAIL.n413 VSUBS 1.39313f
C1209 VTAIL.n414 VSUBS 0.025626f
C1210 VTAIL.n415 VSUBS 0.024957f
C1211 VTAIL.n416 VSUBS 0.013411f
C1212 VTAIL.n417 VSUBS 0.031699f
C1213 VTAIL.n418 VSUBS 0.0142f
C1214 VTAIL.n419 VSUBS 0.024957f
C1215 VTAIL.n420 VSUBS 0.013411f
C1216 VTAIL.n421 VSUBS 0.031699f
C1217 VTAIL.n422 VSUBS 0.0142f
C1218 VTAIL.n423 VSUBS 0.024957f
C1219 VTAIL.n424 VSUBS 0.013411f
C1220 VTAIL.n425 VSUBS 0.031699f
C1221 VTAIL.n426 VSUBS 0.0142f
C1222 VTAIL.n427 VSUBS 0.024957f
C1223 VTAIL.n428 VSUBS 0.013411f
C1224 VTAIL.n429 VSUBS 0.031699f
C1225 VTAIL.n430 VSUBS 0.0142f
C1226 VTAIL.n431 VSUBS 0.180759f
C1227 VTAIL.t0 VSUBS 0.068194f
C1228 VTAIL.n432 VSUBS 0.023774f
C1229 VTAIL.n433 VSUBS 0.023845f
C1230 VTAIL.n434 VSUBS 0.013411f
C1231 VTAIL.n435 VSUBS 1.07312f
C1232 VTAIL.n436 VSUBS 0.024957f
C1233 VTAIL.n437 VSUBS 0.013411f
C1234 VTAIL.n438 VSUBS 0.0142f
C1235 VTAIL.n439 VSUBS 0.031699f
C1236 VTAIL.n440 VSUBS 0.031699f
C1237 VTAIL.n441 VSUBS 0.0142f
C1238 VTAIL.n442 VSUBS 0.013411f
C1239 VTAIL.n443 VSUBS 0.024957f
C1240 VTAIL.n444 VSUBS 0.024957f
C1241 VTAIL.n445 VSUBS 0.013411f
C1242 VTAIL.n446 VSUBS 0.0142f
C1243 VTAIL.n447 VSUBS 0.031699f
C1244 VTAIL.n448 VSUBS 0.031699f
C1245 VTAIL.n449 VSUBS 0.031699f
C1246 VTAIL.n450 VSUBS 0.0142f
C1247 VTAIL.n451 VSUBS 0.013411f
C1248 VTAIL.n452 VSUBS 0.024957f
C1249 VTAIL.n453 VSUBS 0.024957f
C1250 VTAIL.n454 VSUBS 0.013411f
C1251 VTAIL.n455 VSUBS 0.013805f
C1252 VTAIL.n456 VSUBS 0.013805f
C1253 VTAIL.n457 VSUBS 0.031699f
C1254 VTAIL.n458 VSUBS 0.031699f
C1255 VTAIL.n459 VSUBS 0.0142f
C1256 VTAIL.n460 VSUBS 0.013411f
C1257 VTAIL.n461 VSUBS 0.024957f
C1258 VTAIL.n462 VSUBS 0.024957f
C1259 VTAIL.n463 VSUBS 0.013411f
C1260 VTAIL.n464 VSUBS 0.0142f
C1261 VTAIL.n465 VSUBS 0.031699f
C1262 VTAIL.n466 VSUBS 0.070618f
C1263 VTAIL.n467 VSUBS 0.0142f
C1264 VTAIL.n468 VSUBS 0.013411f
C1265 VTAIL.n469 VSUBS 0.05496f
C1266 VTAIL.n470 VSUBS 0.035155f
C1267 VTAIL.n471 VSUBS 1.38845f
C1268 VDD1.t1 VSUBS 0.208209f
C1269 VDD1.t3 VSUBS 0.208209f
C1270 VDD1.n0 VSUBS 1.59326f
C1271 VDD1.t6 VSUBS 0.208209f
C1272 VDD1.t0 VSUBS 0.208209f
C1273 VDD1.n1 VSUBS 1.59211f
C1274 VDD1.t2 VSUBS 0.208209f
C1275 VDD1.t7 VSUBS 0.208209f
C1276 VDD1.n2 VSUBS 1.59211f
C1277 VDD1.n3 VSUBS 3.28823f
C1278 VDD1.t5 VSUBS 0.208209f
C1279 VDD1.t4 VSUBS 0.208209f
C1280 VDD1.n4 VSUBS 1.58408f
C1281 VDD1.n5 VSUBS 2.84588f
C1282 VP.n0 VSUBS 0.048687f
C1283 VP.t5 VSUBS 1.94451f
C1284 VP.n1 VSUBS 0.068146f
C1285 VP.n2 VSUBS 0.036931f
C1286 VP.t0 VSUBS 1.94451f
C1287 VP.n3 VSUBS 0.053685f
C1288 VP.n4 VSUBS 0.036931f
C1289 VP.t2 VSUBS 1.94451f
C1290 VP.n5 VSUBS 0.033826f
C1291 VP.n6 VSUBS 0.048687f
C1292 VP.t3 VSUBS 1.94451f
C1293 VP.n7 VSUBS 0.068146f
C1294 VP.n8 VSUBS 0.036931f
C1295 VP.t7 VSUBS 1.94451f
C1296 VP.n9 VSUBS 0.053685f
C1297 VP.t1 VSUBS 2.10674f
C1298 VP.n10 VSUBS 0.793648f
C1299 VP.t4 VSUBS 1.94451f
C1300 VP.n11 VSUBS 0.791078f
C1301 VP.n12 VSUBS 0.05699f
C1302 VP.n13 VSUBS 0.270805f
C1303 VP.n14 VSUBS 0.036931f
C1304 VP.n15 VSUBS 0.036931f
C1305 VP.n16 VSUBS 0.053685f
C1306 VP.n17 VSUBS 0.05699f
C1307 VP.n18 VSUBS 0.703023f
C1308 VP.n19 VSUBS 0.046171f
C1309 VP.n20 VSUBS 0.036931f
C1310 VP.n21 VSUBS 0.036931f
C1311 VP.n22 VSUBS 0.036931f
C1312 VP.n23 VSUBS 0.033826f
C1313 VP.n24 VSUBS 0.073206f
C1314 VP.n25 VSUBS 0.815348f
C1315 VP.n26 VSUBS 1.80848f
C1316 VP.n27 VSUBS 1.83725f
C1317 VP.t6 VSUBS 1.94451f
C1318 VP.n28 VSUBS 0.815348f
C1319 VP.n29 VSUBS 0.073206f
C1320 VP.n30 VSUBS 0.048687f
C1321 VP.n31 VSUBS 0.036931f
C1322 VP.n32 VSUBS 0.036931f
C1323 VP.n33 VSUBS 0.068146f
C1324 VP.n34 VSUBS 0.046171f
C1325 VP.n35 VSUBS 0.703023f
C1326 VP.n36 VSUBS 0.05699f
C1327 VP.n37 VSUBS 0.036931f
C1328 VP.n38 VSUBS 0.036931f
C1329 VP.n39 VSUBS 0.036931f
C1330 VP.n40 VSUBS 0.053685f
C1331 VP.n41 VSUBS 0.05699f
C1332 VP.n42 VSUBS 0.703023f
C1333 VP.n43 VSUBS 0.046171f
C1334 VP.n44 VSUBS 0.036931f
C1335 VP.n45 VSUBS 0.036931f
C1336 VP.n46 VSUBS 0.036931f
C1337 VP.n47 VSUBS 0.033826f
C1338 VP.n48 VSUBS 0.073206f
C1339 VP.n49 VSUBS 0.815348f
C1340 VP.n50 VSUBS 0.039336f
.ends

