* NGSPICE file created from diff_pair_sample_0656.ext - technology: sky130A

.subckt diff_pair_sample_0656 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=0.29535 pd=2.12 as=0.29535 ps=2.12 w=1.79 l=3.15
X1 VTAIL.t6 VN.t0 VDD2.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=0.29535 pd=2.12 as=0.29535 ps=2.12 w=1.79 l=3.15
X2 VTAIL.t5 VN.t1 VDD2.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.6981 pd=4.36 as=0.29535 ps=2.12 w=1.79 l=3.15
X3 VDD1.t6 VP.t1 VTAIL.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=0.29535 pd=2.12 as=0.29535 ps=2.12 w=1.79 l=3.15
X4 VDD2.t5 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.29535 pd=2.12 as=0.6981 ps=4.36 w=1.79 l=3.15
X5 VDD2.t4 VN.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.29535 pd=2.12 as=0.29535 ps=2.12 w=1.79 l=3.15
X6 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=0.6981 pd=4.36 as=0 ps=0 w=1.79 l=3.15
X7 VTAIL.t3 VN.t4 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.6981 pd=4.36 as=0.29535 ps=2.12 w=1.79 l=3.15
X8 VDD1.t3 VP.t2 VTAIL.t13 B.t2 sky130_fd_pr__nfet_01v8 ad=0.29535 pd=2.12 as=0.6981 ps=4.36 w=1.79 l=3.15
X9 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=0.6981 pd=4.36 as=0 ps=0 w=1.79 l=3.15
X10 VDD2.t2 VN.t5 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.29535 pd=2.12 as=0.29535 ps=2.12 w=1.79 l=3.15
X11 VDD1.t4 VP.t3 VTAIL.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=0.29535 pd=2.12 as=0.6981 ps=4.36 w=1.79 l=3.15
X12 VTAIL.t11 VP.t4 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.6981 pd=4.36 as=0.29535 ps=2.12 w=1.79 l=3.15
X13 VTAIL.t10 VP.t5 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.29535 pd=2.12 as=0.29535 ps=2.12 w=1.79 l=3.15
X14 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=0.6981 pd=4.36 as=0 ps=0 w=1.79 l=3.15
X15 VDD2.t1 VN.t6 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.29535 pd=2.12 as=0.6981 ps=4.36 w=1.79 l=3.15
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.6981 pd=4.36 as=0 ps=0 w=1.79 l=3.15
X17 VDD1.t2 VP.t6 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=0.29535 pd=2.12 as=0.29535 ps=2.12 w=1.79 l=3.15
X18 VTAIL.t0 VN.t7 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.29535 pd=2.12 as=0.29535 ps=2.12 w=1.79 l=3.15
X19 VTAIL.t8 VP.t7 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.6981 pd=4.36 as=0.29535 ps=2.12 w=1.79 l=3.15
R0 VP.n21 VP.n18 161.3
R1 VP.n23 VP.n22 161.3
R2 VP.n24 VP.n17 161.3
R3 VP.n26 VP.n25 161.3
R4 VP.n27 VP.n16 161.3
R5 VP.n29 VP.n28 161.3
R6 VP.n31 VP.n30 161.3
R7 VP.n32 VP.n14 161.3
R8 VP.n34 VP.n33 161.3
R9 VP.n35 VP.n13 161.3
R10 VP.n37 VP.n36 161.3
R11 VP.n38 VP.n12 161.3
R12 VP.n40 VP.n39 161.3
R13 VP.n75 VP.n74 161.3
R14 VP.n73 VP.n1 161.3
R15 VP.n72 VP.n71 161.3
R16 VP.n70 VP.n2 161.3
R17 VP.n69 VP.n68 161.3
R18 VP.n67 VP.n3 161.3
R19 VP.n66 VP.n65 161.3
R20 VP.n64 VP.n63 161.3
R21 VP.n62 VP.n5 161.3
R22 VP.n61 VP.n60 161.3
R23 VP.n59 VP.n6 161.3
R24 VP.n58 VP.n57 161.3
R25 VP.n56 VP.n7 161.3
R26 VP.n54 VP.n53 161.3
R27 VP.n52 VP.n8 161.3
R28 VP.n51 VP.n50 161.3
R29 VP.n49 VP.n9 161.3
R30 VP.n48 VP.n47 161.3
R31 VP.n46 VP.n10 161.3
R32 VP.n45 VP.n44 161.3
R33 VP.n43 VP.n42 67.0684
R34 VP.n76 VP.n0 67.0684
R35 VP.n41 VP.n11 67.0684
R36 VP.n49 VP.n48 56.5193
R37 VP.n61 VP.n6 56.5193
R38 VP.n72 VP.n2 56.5193
R39 VP.n37 VP.n13 56.5193
R40 VP.n26 VP.n17 56.5193
R41 VP.n20 VP.n19 50.0328
R42 VP.n19 VP.t7 47.0991
R43 VP.n42 VP.n41 45.9387
R44 VP.n44 VP.n10 24.4675
R45 VP.n48 VP.n10 24.4675
R46 VP.n50 VP.n49 24.4675
R47 VP.n50 VP.n8 24.4675
R48 VP.n54 VP.n8 24.4675
R49 VP.n57 VP.n56 24.4675
R50 VP.n57 VP.n6 24.4675
R51 VP.n62 VP.n61 24.4675
R52 VP.n63 VP.n62 24.4675
R53 VP.n67 VP.n66 24.4675
R54 VP.n68 VP.n67 24.4675
R55 VP.n68 VP.n2 24.4675
R56 VP.n73 VP.n72 24.4675
R57 VP.n74 VP.n73 24.4675
R58 VP.n38 VP.n37 24.4675
R59 VP.n39 VP.n38 24.4675
R60 VP.n27 VP.n26 24.4675
R61 VP.n28 VP.n27 24.4675
R62 VP.n32 VP.n31 24.4675
R63 VP.n33 VP.n32 24.4675
R64 VP.n33 VP.n13 24.4675
R65 VP.n22 VP.n21 24.4675
R66 VP.n22 VP.n17 24.4675
R67 VP.n56 VP.n55 23.9782
R68 VP.n63 VP.n4 23.9782
R69 VP.n28 VP.n15 23.9782
R70 VP.n21 VP.n20 23.9782
R71 VP.n44 VP.n43 22.9995
R72 VP.n74 VP.n0 22.9995
R73 VP.n39 VP.n11 22.9995
R74 VP.n43 VP.t4 13.6954
R75 VP.n55 VP.t6 13.6954
R76 VP.n4 VP.t5 13.6954
R77 VP.n0 VP.t3 13.6954
R78 VP.n11 VP.t2 13.6954
R79 VP.n15 VP.t0 13.6954
R80 VP.n20 VP.t1 13.6954
R81 VP.n19 VP.n18 3.77028
R82 VP.n55 VP.n54 0.48984
R83 VP.n66 VP.n4 0.48984
R84 VP.n31 VP.n15 0.48984
R85 VP.n41 VP.n40 0.354971
R86 VP.n45 VP.n42 0.354971
R87 VP.n76 VP.n75 0.354971
R88 VP VP.n76 0.26696
R89 VP.n23 VP.n18 0.189894
R90 VP.n24 VP.n23 0.189894
R91 VP.n25 VP.n24 0.189894
R92 VP.n25 VP.n16 0.189894
R93 VP.n29 VP.n16 0.189894
R94 VP.n30 VP.n29 0.189894
R95 VP.n30 VP.n14 0.189894
R96 VP.n34 VP.n14 0.189894
R97 VP.n35 VP.n34 0.189894
R98 VP.n36 VP.n35 0.189894
R99 VP.n36 VP.n12 0.189894
R100 VP.n40 VP.n12 0.189894
R101 VP.n46 VP.n45 0.189894
R102 VP.n47 VP.n46 0.189894
R103 VP.n47 VP.n9 0.189894
R104 VP.n51 VP.n9 0.189894
R105 VP.n52 VP.n51 0.189894
R106 VP.n53 VP.n52 0.189894
R107 VP.n53 VP.n7 0.189894
R108 VP.n58 VP.n7 0.189894
R109 VP.n59 VP.n58 0.189894
R110 VP.n60 VP.n59 0.189894
R111 VP.n60 VP.n5 0.189894
R112 VP.n64 VP.n5 0.189894
R113 VP.n65 VP.n64 0.189894
R114 VP.n65 VP.n3 0.189894
R115 VP.n69 VP.n3 0.189894
R116 VP.n70 VP.n69 0.189894
R117 VP.n71 VP.n70 0.189894
R118 VP.n71 VP.n1 0.189894
R119 VP.n75 VP.n1 0.189894
R120 VDD1 VDD1.n0 103.175
R121 VDD1.n3 VDD1.n2 103.061
R122 VDD1.n3 VDD1.n1 103.061
R123 VDD1.n5 VDD1.n4 101.618
R124 VDD1.n5 VDD1.n3 39.3414
R125 VDD1.n4 VDD1.t0 11.062
R126 VDD1.n4 VDD1.t3 11.062
R127 VDD1.n0 VDD1.t7 11.062
R128 VDD1.n0 VDD1.t6 11.062
R129 VDD1.n2 VDD1.t1 11.062
R130 VDD1.n2 VDD1.t4 11.062
R131 VDD1.n1 VDD1.t5 11.062
R132 VDD1.n1 VDD1.t2 11.062
R133 VDD1 VDD1.n5 1.44231
R134 VTAIL.n66 VTAIL.n64 289.615
R135 VTAIL.n4 VTAIL.n2 289.615
R136 VTAIL.n12 VTAIL.n10 289.615
R137 VTAIL.n22 VTAIL.n20 289.615
R138 VTAIL.n58 VTAIL.n56 289.615
R139 VTAIL.n48 VTAIL.n46 289.615
R140 VTAIL.n40 VTAIL.n38 289.615
R141 VTAIL.n30 VTAIL.n28 289.615
R142 VTAIL.n67 VTAIL.n66 185
R143 VTAIL.n5 VTAIL.n4 185
R144 VTAIL.n13 VTAIL.n12 185
R145 VTAIL.n23 VTAIL.n22 185
R146 VTAIL.n59 VTAIL.n58 185
R147 VTAIL.n49 VTAIL.n48 185
R148 VTAIL.n41 VTAIL.n40 185
R149 VTAIL.n31 VTAIL.n30 185
R150 VTAIL.t2 VTAIL.n65 164.876
R151 VTAIL.t3 VTAIL.n3 164.876
R152 VTAIL.t12 VTAIL.n11 164.876
R153 VTAIL.t11 VTAIL.n21 164.876
R154 VTAIL.t13 VTAIL.n57 164.876
R155 VTAIL.t8 VTAIL.n47 164.876
R156 VTAIL.t1 VTAIL.n39 164.876
R157 VTAIL.t5 VTAIL.n29 164.876
R158 VTAIL.n55 VTAIL.n54 84.9382
R159 VTAIL.n37 VTAIL.n36 84.9382
R160 VTAIL.n1 VTAIL.n0 84.9382
R161 VTAIL.n19 VTAIL.n18 84.9382
R162 VTAIL.n66 VTAIL.t2 52.3082
R163 VTAIL.n4 VTAIL.t3 52.3082
R164 VTAIL.n12 VTAIL.t12 52.3082
R165 VTAIL.n22 VTAIL.t11 52.3082
R166 VTAIL.n58 VTAIL.t13 52.3082
R167 VTAIL.n48 VTAIL.t8 52.3082
R168 VTAIL.n40 VTAIL.t1 52.3082
R169 VTAIL.n30 VTAIL.t5 52.3082
R170 VTAIL.n71 VTAIL.n70 34.3187
R171 VTAIL.n9 VTAIL.n8 34.3187
R172 VTAIL.n17 VTAIL.n16 34.3187
R173 VTAIL.n27 VTAIL.n26 34.3187
R174 VTAIL.n63 VTAIL.n62 34.3187
R175 VTAIL.n53 VTAIL.n52 34.3187
R176 VTAIL.n45 VTAIL.n44 34.3187
R177 VTAIL.n35 VTAIL.n34 34.3187
R178 VTAIL.n71 VTAIL.n63 16.91
R179 VTAIL.n35 VTAIL.n27 16.91
R180 VTAIL.n67 VTAIL.n65 14.7318
R181 VTAIL.n5 VTAIL.n3 14.7318
R182 VTAIL.n13 VTAIL.n11 14.7318
R183 VTAIL.n23 VTAIL.n21 14.7318
R184 VTAIL.n59 VTAIL.n57 14.7318
R185 VTAIL.n49 VTAIL.n47 14.7318
R186 VTAIL.n41 VTAIL.n39 14.7318
R187 VTAIL.n31 VTAIL.n29 14.7318
R188 VTAIL.n68 VTAIL.n64 12.8005
R189 VTAIL.n6 VTAIL.n2 12.8005
R190 VTAIL.n14 VTAIL.n10 12.8005
R191 VTAIL.n24 VTAIL.n20 12.8005
R192 VTAIL.n60 VTAIL.n56 12.8005
R193 VTAIL.n50 VTAIL.n46 12.8005
R194 VTAIL.n42 VTAIL.n38 12.8005
R195 VTAIL.n32 VTAIL.n28 12.8005
R196 VTAIL.n0 VTAIL.t7 11.062
R197 VTAIL.n0 VTAIL.t6 11.062
R198 VTAIL.n18 VTAIL.t9 11.062
R199 VTAIL.n18 VTAIL.t10 11.062
R200 VTAIL.n54 VTAIL.t14 11.062
R201 VTAIL.n54 VTAIL.t15 11.062
R202 VTAIL.n36 VTAIL.t4 11.062
R203 VTAIL.n36 VTAIL.t0 11.062
R204 VTAIL.n70 VTAIL.n69 9.45567
R205 VTAIL.n8 VTAIL.n7 9.45567
R206 VTAIL.n16 VTAIL.n15 9.45567
R207 VTAIL.n26 VTAIL.n25 9.45567
R208 VTAIL.n62 VTAIL.n61 9.45567
R209 VTAIL.n52 VTAIL.n51 9.45567
R210 VTAIL.n44 VTAIL.n43 9.45567
R211 VTAIL.n34 VTAIL.n33 9.45567
R212 VTAIL.n69 VTAIL.n68 9.3005
R213 VTAIL.n7 VTAIL.n6 9.3005
R214 VTAIL.n15 VTAIL.n14 9.3005
R215 VTAIL.n25 VTAIL.n24 9.3005
R216 VTAIL.n61 VTAIL.n60 9.3005
R217 VTAIL.n51 VTAIL.n50 9.3005
R218 VTAIL.n43 VTAIL.n42 9.3005
R219 VTAIL.n33 VTAIL.n32 9.3005
R220 VTAIL.n69 VTAIL.n65 5.62509
R221 VTAIL.n7 VTAIL.n3 5.62509
R222 VTAIL.n15 VTAIL.n11 5.62509
R223 VTAIL.n25 VTAIL.n21 5.62509
R224 VTAIL.n61 VTAIL.n57 5.62509
R225 VTAIL.n51 VTAIL.n47 5.62509
R226 VTAIL.n43 VTAIL.n39 5.62509
R227 VTAIL.n33 VTAIL.n29 5.62509
R228 VTAIL.n37 VTAIL.n35 3.0005
R229 VTAIL.n45 VTAIL.n37 3.0005
R230 VTAIL.n55 VTAIL.n53 3.0005
R231 VTAIL.n63 VTAIL.n55 3.0005
R232 VTAIL.n27 VTAIL.n19 3.0005
R233 VTAIL.n19 VTAIL.n17 3.0005
R234 VTAIL.n9 VTAIL.n1 3.0005
R235 VTAIL VTAIL.n71 2.94231
R236 VTAIL.n70 VTAIL.n64 1.16414
R237 VTAIL.n8 VTAIL.n2 1.16414
R238 VTAIL.n16 VTAIL.n10 1.16414
R239 VTAIL.n26 VTAIL.n20 1.16414
R240 VTAIL.n62 VTAIL.n56 1.16414
R241 VTAIL.n52 VTAIL.n46 1.16414
R242 VTAIL.n44 VTAIL.n38 1.16414
R243 VTAIL.n34 VTAIL.n28 1.16414
R244 VTAIL.n53 VTAIL.n45 0.470328
R245 VTAIL.n17 VTAIL.n9 0.470328
R246 VTAIL.n68 VTAIL.n67 0.388379
R247 VTAIL.n6 VTAIL.n5 0.388379
R248 VTAIL.n14 VTAIL.n13 0.388379
R249 VTAIL.n24 VTAIL.n23 0.388379
R250 VTAIL.n60 VTAIL.n59 0.388379
R251 VTAIL.n50 VTAIL.n49 0.388379
R252 VTAIL.n42 VTAIL.n41 0.388379
R253 VTAIL.n32 VTAIL.n31 0.388379
R254 VTAIL VTAIL.n1 0.0586897
R255 B.n651 B.n650 585
R256 B.n652 B.n651 585
R257 B.n192 B.n126 585
R258 B.n191 B.n190 585
R259 B.n189 B.n188 585
R260 B.n187 B.n186 585
R261 B.n185 B.n184 585
R262 B.n183 B.n182 585
R263 B.n181 B.n180 585
R264 B.n179 B.n178 585
R265 B.n177 B.n176 585
R266 B.n175 B.n174 585
R267 B.n173 B.n172 585
R268 B.n170 B.n169 585
R269 B.n168 B.n167 585
R270 B.n166 B.n165 585
R271 B.n164 B.n163 585
R272 B.n162 B.n161 585
R273 B.n160 B.n159 585
R274 B.n158 B.n157 585
R275 B.n156 B.n155 585
R276 B.n154 B.n153 585
R277 B.n152 B.n151 585
R278 B.n150 B.n149 585
R279 B.n148 B.n147 585
R280 B.n146 B.n145 585
R281 B.n144 B.n143 585
R282 B.n142 B.n141 585
R283 B.n140 B.n139 585
R284 B.n138 B.n137 585
R285 B.n136 B.n135 585
R286 B.n134 B.n133 585
R287 B.n110 B.n109 585
R288 B.n655 B.n654 585
R289 B.n649 B.n127 585
R290 B.n127 B.n107 585
R291 B.n648 B.n106 585
R292 B.n659 B.n106 585
R293 B.n647 B.n105 585
R294 B.n660 B.n105 585
R295 B.n646 B.n104 585
R296 B.n661 B.n104 585
R297 B.n645 B.n644 585
R298 B.n644 B.n100 585
R299 B.n643 B.n99 585
R300 B.n667 B.n99 585
R301 B.n642 B.n98 585
R302 B.n668 B.n98 585
R303 B.n641 B.n97 585
R304 B.n669 B.n97 585
R305 B.n640 B.n639 585
R306 B.n639 B.n96 585
R307 B.n638 B.n92 585
R308 B.n675 B.n92 585
R309 B.n637 B.n91 585
R310 B.n676 B.n91 585
R311 B.n636 B.n90 585
R312 B.n677 B.n90 585
R313 B.n635 B.n634 585
R314 B.n634 B.n86 585
R315 B.n633 B.n85 585
R316 B.n683 B.n85 585
R317 B.n632 B.n84 585
R318 B.n684 B.n84 585
R319 B.n631 B.n83 585
R320 B.n685 B.n83 585
R321 B.n630 B.n629 585
R322 B.n629 B.n79 585
R323 B.n628 B.n78 585
R324 B.n691 B.n78 585
R325 B.n627 B.n77 585
R326 B.n692 B.n77 585
R327 B.n626 B.n76 585
R328 B.n693 B.n76 585
R329 B.n625 B.n624 585
R330 B.n624 B.n72 585
R331 B.n623 B.n71 585
R332 B.n699 B.n71 585
R333 B.n622 B.n70 585
R334 B.n700 B.n70 585
R335 B.n621 B.n69 585
R336 B.n701 B.n69 585
R337 B.n620 B.n619 585
R338 B.n619 B.n65 585
R339 B.n618 B.n64 585
R340 B.n707 B.n64 585
R341 B.n617 B.n63 585
R342 B.n708 B.n63 585
R343 B.n616 B.n62 585
R344 B.n709 B.n62 585
R345 B.n615 B.n614 585
R346 B.n614 B.n58 585
R347 B.n613 B.n57 585
R348 B.n715 B.n57 585
R349 B.n612 B.n56 585
R350 B.n716 B.n56 585
R351 B.n611 B.n55 585
R352 B.n717 B.n55 585
R353 B.n610 B.n609 585
R354 B.n609 B.n54 585
R355 B.n608 B.n50 585
R356 B.n723 B.n50 585
R357 B.n607 B.n49 585
R358 B.n724 B.n49 585
R359 B.n606 B.n48 585
R360 B.n725 B.n48 585
R361 B.n605 B.n604 585
R362 B.n604 B.n44 585
R363 B.n603 B.n43 585
R364 B.n731 B.n43 585
R365 B.n602 B.n42 585
R366 B.n732 B.n42 585
R367 B.n601 B.n41 585
R368 B.n733 B.n41 585
R369 B.n600 B.n599 585
R370 B.n599 B.n37 585
R371 B.n598 B.n36 585
R372 B.n739 B.n36 585
R373 B.n597 B.n35 585
R374 B.n740 B.n35 585
R375 B.n596 B.n34 585
R376 B.n741 B.n34 585
R377 B.n595 B.n594 585
R378 B.n594 B.n30 585
R379 B.n593 B.n29 585
R380 B.n747 B.n29 585
R381 B.n592 B.n28 585
R382 B.n748 B.n28 585
R383 B.n591 B.n27 585
R384 B.n749 B.n27 585
R385 B.n590 B.n589 585
R386 B.n589 B.n23 585
R387 B.n588 B.n22 585
R388 B.n755 B.n22 585
R389 B.n587 B.n21 585
R390 B.n756 B.n21 585
R391 B.n586 B.n20 585
R392 B.n757 B.n20 585
R393 B.n585 B.n584 585
R394 B.n584 B.n19 585
R395 B.n583 B.n15 585
R396 B.n763 B.n15 585
R397 B.n582 B.n14 585
R398 B.n764 B.n14 585
R399 B.n581 B.n13 585
R400 B.n765 B.n13 585
R401 B.n580 B.n579 585
R402 B.n579 B.n12 585
R403 B.n578 B.n577 585
R404 B.n578 B.n8 585
R405 B.n576 B.n7 585
R406 B.n772 B.n7 585
R407 B.n575 B.n6 585
R408 B.n773 B.n6 585
R409 B.n574 B.n5 585
R410 B.n774 B.n5 585
R411 B.n573 B.n572 585
R412 B.n572 B.n4 585
R413 B.n571 B.n193 585
R414 B.n571 B.n570 585
R415 B.n561 B.n194 585
R416 B.n195 B.n194 585
R417 B.n563 B.n562 585
R418 B.n564 B.n563 585
R419 B.n560 B.n200 585
R420 B.n200 B.n199 585
R421 B.n559 B.n558 585
R422 B.n558 B.n557 585
R423 B.n202 B.n201 585
R424 B.n550 B.n202 585
R425 B.n549 B.n548 585
R426 B.n551 B.n549 585
R427 B.n547 B.n207 585
R428 B.n207 B.n206 585
R429 B.n546 B.n545 585
R430 B.n545 B.n544 585
R431 B.n209 B.n208 585
R432 B.n210 B.n209 585
R433 B.n537 B.n536 585
R434 B.n538 B.n537 585
R435 B.n535 B.n215 585
R436 B.n215 B.n214 585
R437 B.n534 B.n533 585
R438 B.n533 B.n532 585
R439 B.n217 B.n216 585
R440 B.n218 B.n217 585
R441 B.n525 B.n524 585
R442 B.n526 B.n525 585
R443 B.n523 B.n222 585
R444 B.n226 B.n222 585
R445 B.n522 B.n521 585
R446 B.n521 B.n520 585
R447 B.n224 B.n223 585
R448 B.n225 B.n224 585
R449 B.n513 B.n512 585
R450 B.n514 B.n513 585
R451 B.n511 B.n231 585
R452 B.n231 B.n230 585
R453 B.n510 B.n509 585
R454 B.n509 B.n508 585
R455 B.n233 B.n232 585
R456 B.n234 B.n233 585
R457 B.n501 B.n500 585
R458 B.n502 B.n501 585
R459 B.n499 B.n239 585
R460 B.n239 B.n238 585
R461 B.n498 B.n497 585
R462 B.n497 B.n496 585
R463 B.n241 B.n240 585
R464 B.n489 B.n241 585
R465 B.n488 B.n487 585
R466 B.n490 B.n488 585
R467 B.n486 B.n246 585
R468 B.n246 B.n245 585
R469 B.n485 B.n484 585
R470 B.n484 B.n483 585
R471 B.n248 B.n247 585
R472 B.n249 B.n248 585
R473 B.n476 B.n475 585
R474 B.n477 B.n476 585
R475 B.n474 B.n254 585
R476 B.n254 B.n253 585
R477 B.n473 B.n472 585
R478 B.n472 B.n471 585
R479 B.n256 B.n255 585
R480 B.n257 B.n256 585
R481 B.n464 B.n463 585
R482 B.n465 B.n464 585
R483 B.n462 B.n261 585
R484 B.n265 B.n261 585
R485 B.n461 B.n460 585
R486 B.n460 B.n459 585
R487 B.n263 B.n262 585
R488 B.n264 B.n263 585
R489 B.n452 B.n451 585
R490 B.n453 B.n452 585
R491 B.n450 B.n270 585
R492 B.n270 B.n269 585
R493 B.n449 B.n448 585
R494 B.n448 B.n447 585
R495 B.n272 B.n271 585
R496 B.n273 B.n272 585
R497 B.n440 B.n439 585
R498 B.n441 B.n440 585
R499 B.n438 B.n278 585
R500 B.n278 B.n277 585
R501 B.n437 B.n436 585
R502 B.n436 B.n435 585
R503 B.n280 B.n279 585
R504 B.n281 B.n280 585
R505 B.n428 B.n427 585
R506 B.n429 B.n428 585
R507 B.n426 B.n286 585
R508 B.n286 B.n285 585
R509 B.n425 B.n424 585
R510 B.n424 B.n423 585
R511 B.n288 B.n287 585
R512 B.n416 B.n288 585
R513 B.n415 B.n414 585
R514 B.n417 B.n415 585
R515 B.n413 B.n293 585
R516 B.n293 B.n292 585
R517 B.n412 B.n411 585
R518 B.n411 B.n410 585
R519 B.n295 B.n294 585
R520 B.n296 B.n295 585
R521 B.n403 B.n402 585
R522 B.n404 B.n403 585
R523 B.n401 B.n301 585
R524 B.n301 B.n300 585
R525 B.n400 B.n399 585
R526 B.n399 B.n398 585
R527 B.n303 B.n302 585
R528 B.n304 B.n303 585
R529 B.n394 B.n393 585
R530 B.n307 B.n306 585
R531 B.n390 B.n389 585
R532 B.n391 B.n390 585
R533 B.n388 B.n323 585
R534 B.n387 B.n386 585
R535 B.n385 B.n384 585
R536 B.n383 B.n382 585
R537 B.n381 B.n380 585
R538 B.n379 B.n378 585
R539 B.n377 B.n376 585
R540 B.n375 B.n374 585
R541 B.n373 B.n372 585
R542 B.n370 B.n369 585
R543 B.n368 B.n367 585
R544 B.n366 B.n365 585
R545 B.n364 B.n363 585
R546 B.n362 B.n361 585
R547 B.n360 B.n359 585
R548 B.n358 B.n357 585
R549 B.n356 B.n355 585
R550 B.n354 B.n353 585
R551 B.n352 B.n351 585
R552 B.n350 B.n349 585
R553 B.n348 B.n347 585
R554 B.n346 B.n345 585
R555 B.n344 B.n343 585
R556 B.n342 B.n341 585
R557 B.n340 B.n339 585
R558 B.n338 B.n337 585
R559 B.n336 B.n335 585
R560 B.n334 B.n333 585
R561 B.n332 B.n331 585
R562 B.n330 B.n329 585
R563 B.n395 B.n305 585
R564 B.n305 B.n304 585
R565 B.n397 B.n396 585
R566 B.n398 B.n397 585
R567 B.n299 B.n298 585
R568 B.n300 B.n299 585
R569 B.n406 B.n405 585
R570 B.n405 B.n404 585
R571 B.n407 B.n297 585
R572 B.n297 B.n296 585
R573 B.n409 B.n408 585
R574 B.n410 B.n409 585
R575 B.n291 B.n290 585
R576 B.n292 B.n291 585
R577 B.n419 B.n418 585
R578 B.n418 B.n417 585
R579 B.n420 B.n289 585
R580 B.n416 B.n289 585
R581 B.n422 B.n421 585
R582 B.n423 B.n422 585
R583 B.n284 B.n283 585
R584 B.n285 B.n284 585
R585 B.n431 B.n430 585
R586 B.n430 B.n429 585
R587 B.n432 B.n282 585
R588 B.n282 B.n281 585
R589 B.n434 B.n433 585
R590 B.n435 B.n434 585
R591 B.n276 B.n275 585
R592 B.n277 B.n276 585
R593 B.n443 B.n442 585
R594 B.n442 B.n441 585
R595 B.n444 B.n274 585
R596 B.n274 B.n273 585
R597 B.n446 B.n445 585
R598 B.n447 B.n446 585
R599 B.n268 B.n267 585
R600 B.n269 B.n268 585
R601 B.n455 B.n454 585
R602 B.n454 B.n453 585
R603 B.n456 B.n266 585
R604 B.n266 B.n264 585
R605 B.n458 B.n457 585
R606 B.n459 B.n458 585
R607 B.n260 B.n259 585
R608 B.n265 B.n260 585
R609 B.n467 B.n466 585
R610 B.n466 B.n465 585
R611 B.n468 B.n258 585
R612 B.n258 B.n257 585
R613 B.n470 B.n469 585
R614 B.n471 B.n470 585
R615 B.n252 B.n251 585
R616 B.n253 B.n252 585
R617 B.n479 B.n478 585
R618 B.n478 B.n477 585
R619 B.n480 B.n250 585
R620 B.n250 B.n249 585
R621 B.n482 B.n481 585
R622 B.n483 B.n482 585
R623 B.n244 B.n243 585
R624 B.n245 B.n244 585
R625 B.n492 B.n491 585
R626 B.n491 B.n490 585
R627 B.n493 B.n242 585
R628 B.n489 B.n242 585
R629 B.n495 B.n494 585
R630 B.n496 B.n495 585
R631 B.n237 B.n236 585
R632 B.n238 B.n237 585
R633 B.n504 B.n503 585
R634 B.n503 B.n502 585
R635 B.n505 B.n235 585
R636 B.n235 B.n234 585
R637 B.n507 B.n506 585
R638 B.n508 B.n507 585
R639 B.n229 B.n228 585
R640 B.n230 B.n229 585
R641 B.n516 B.n515 585
R642 B.n515 B.n514 585
R643 B.n517 B.n227 585
R644 B.n227 B.n225 585
R645 B.n519 B.n518 585
R646 B.n520 B.n519 585
R647 B.n221 B.n220 585
R648 B.n226 B.n221 585
R649 B.n528 B.n527 585
R650 B.n527 B.n526 585
R651 B.n529 B.n219 585
R652 B.n219 B.n218 585
R653 B.n531 B.n530 585
R654 B.n532 B.n531 585
R655 B.n213 B.n212 585
R656 B.n214 B.n213 585
R657 B.n540 B.n539 585
R658 B.n539 B.n538 585
R659 B.n541 B.n211 585
R660 B.n211 B.n210 585
R661 B.n543 B.n542 585
R662 B.n544 B.n543 585
R663 B.n205 B.n204 585
R664 B.n206 B.n205 585
R665 B.n553 B.n552 585
R666 B.n552 B.n551 585
R667 B.n554 B.n203 585
R668 B.n550 B.n203 585
R669 B.n556 B.n555 585
R670 B.n557 B.n556 585
R671 B.n198 B.n197 585
R672 B.n199 B.n198 585
R673 B.n566 B.n565 585
R674 B.n565 B.n564 585
R675 B.n567 B.n196 585
R676 B.n196 B.n195 585
R677 B.n569 B.n568 585
R678 B.n570 B.n569 585
R679 B.n3 B.n0 585
R680 B.n4 B.n3 585
R681 B.n771 B.n1 585
R682 B.n772 B.n771 585
R683 B.n770 B.n769 585
R684 B.n770 B.n8 585
R685 B.n768 B.n9 585
R686 B.n12 B.n9 585
R687 B.n767 B.n766 585
R688 B.n766 B.n765 585
R689 B.n11 B.n10 585
R690 B.n764 B.n11 585
R691 B.n762 B.n761 585
R692 B.n763 B.n762 585
R693 B.n760 B.n16 585
R694 B.n19 B.n16 585
R695 B.n759 B.n758 585
R696 B.n758 B.n757 585
R697 B.n18 B.n17 585
R698 B.n756 B.n18 585
R699 B.n754 B.n753 585
R700 B.n755 B.n754 585
R701 B.n752 B.n24 585
R702 B.n24 B.n23 585
R703 B.n751 B.n750 585
R704 B.n750 B.n749 585
R705 B.n26 B.n25 585
R706 B.n748 B.n26 585
R707 B.n746 B.n745 585
R708 B.n747 B.n746 585
R709 B.n744 B.n31 585
R710 B.n31 B.n30 585
R711 B.n743 B.n742 585
R712 B.n742 B.n741 585
R713 B.n33 B.n32 585
R714 B.n740 B.n33 585
R715 B.n738 B.n737 585
R716 B.n739 B.n738 585
R717 B.n736 B.n38 585
R718 B.n38 B.n37 585
R719 B.n735 B.n734 585
R720 B.n734 B.n733 585
R721 B.n40 B.n39 585
R722 B.n732 B.n40 585
R723 B.n730 B.n729 585
R724 B.n731 B.n730 585
R725 B.n728 B.n45 585
R726 B.n45 B.n44 585
R727 B.n727 B.n726 585
R728 B.n726 B.n725 585
R729 B.n47 B.n46 585
R730 B.n724 B.n47 585
R731 B.n722 B.n721 585
R732 B.n723 B.n722 585
R733 B.n720 B.n51 585
R734 B.n54 B.n51 585
R735 B.n719 B.n718 585
R736 B.n718 B.n717 585
R737 B.n53 B.n52 585
R738 B.n716 B.n53 585
R739 B.n714 B.n713 585
R740 B.n715 B.n714 585
R741 B.n712 B.n59 585
R742 B.n59 B.n58 585
R743 B.n711 B.n710 585
R744 B.n710 B.n709 585
R745 B.n61 B.n60 585
R746 B.n708 B.n61 585
R747 B.n706 B.n705 585
R748 B.n707 B.n706 585
R749 B.n704 B.n66 585
R750 B.n66 B.n65 585
R751 B.n703 B.n702 585
R752 B.n702 B.n701 585
R753 B.n68 B.n67 585
R754 B.n700 B.n68 585
R755 B.n698 B.n697 585
R756 B.n699 B.n698 585
R757 B.n696 B.n73 585
R758 B.n73 B.n72 585
R759 B.n695 B.n694 585
R760 B.n694 B.n693 585
R761 B.n75 B.n74 585
R762 B.n692 B.n75 585
R763 B.n690 B.n689 585
R764 B.n691 B.n690 585
R765 B.n688 B.n80 585
R766 B.n80 B.n79 585
R767 B.n687 B.n686 585
R768 B.n686 B.n685 585
R769 B.n82 B.n81 585
R770 B.n684 B.n82 585
R771 B.n682 B.n681 585
R772 B.n683 B.n682 585
R773 B.n680 B.n87 585
R774 B.n87 B.n86 585
R775 B.n679 B.n678 585
R776 B.n678 B.n677 585
R777 B.n89 B.n88 585
R778 B.n676 B.n89 585
R779 B.n674 B.n673 585
R780 B.n675 B.n674 585
R781 B.n672 B.n93 585
R782 B.n96 B.n93 585
R783 B.n671 B.n670 585
R784 B.n670 B.n669 585
R785 B.n95 B.n94 585
R786 B.n668 B.n95 585
R787 B.n666 B.n665 585
R788 B.n667 B.n666 585
R789 B.n664 B.n101 585
R790 B.n101 B.n100 585
R791 B.n663 B.n662 585
R792 B.n662 B.n661 585
R793 B.n103 B.n102 585
R794 B.n660 B.n103 585
R795 B.n658 B.n657 585
R796 B.n659 B.n658 585
R797 B.n656 B.n108 585
R798 B.n108 B.n107 585
R799 B.n775 B.n774 585
R800 B.n773 B.n2 585
R801 B.n654 B.n108 444.452
R802 B.n651 B.n127 444.452
R803 B.n329 B.n303 444.452
R804 B.n393 B.n305 444.452
R805 B.n652 B.n125 256.663
R806 B.n652 B.n124 256.663
R807 B.n652 B.n123 256.663
R808 B.n652 B.n122 256.663
R809 B.n652 B.n121 256.663
R810 B.n652 B.n120 256.663
R811 B.n652 B.n119 256.663
R812 B.n652 B.n118 256.663
R813 B.n652 B.n117 256.663
R814 B.n652 B.n116 256.663
R815 B.n652 B.n115 256.663
R816 B.n652 B.n114 256.663
R817 B.n652 B.n113 256.663
R818 B.n652 B.n112 256.663
R819 B.n652 B.n111 256.663
R820 B.n653 B.n652 256.663
R821 B.n392 B.n391 256.663
R822 B.n391 B.n308 256.663
R823 B.n391 B.n309 256.663
R824 B.n391 B.n310 256.663
R825 B.n391 B.n311 256.663
R826 B.n391 B.n312 256.663
R827 B.n391 B.n313 256.663
R828 B.n391 B.n314 256.663
R829 B.n391 B.n315 256.663
R830 B.n391 B.n316 256.663
R831 B.n391 B.n317 256.663
R832 B.n391 B.n318 256.663
R833 B.n391 B.n319 256.663
R834 B.n391 B.n320 256.663
R835 B.n391 B.n321 256.663
R836 B.n391 B.n322 256.663
R837 B.n777 B.n776 256.663
R838 B.n130 B.t8 222.445
R839 B.n128 B.t19 222.445
R840 B.n326 B.t16 222.445
R841 B.n324 B.t12 222.445
R842 B.n128 B.t20 186.436
R843 B.n326 B.t18 186.436
R844 B.n130 B.t10 186.436
R845 B.n324 B.t15 186.436
R846 B.n391 B.n304 169.71
R847 B.n652 B.n107 169.71
R848 B.n133 B.n110 163.367
R849 B.n137 B.n136 163.367
R850 B.n141 B.n140 163.367
R851 B.n145 B.n144 163.367
R852 B.n149 B.n148 163.367
R853 B.n153 B.n152 163.367
R854 B.n157 B.n156 163.367
R855 B.n161 B.n160 163.367
R856 B.n165 B.n164 163.367
R857 B.n169 B.n168 163.367
R858 B.n174 B.n173 163.367
R859 B.n178 B.n177 163.367
R860 B.n182 B.n181 163.367
R861 B.n186 B.n185 163.367
R862 B.n190 B.n189 163.367
R863 B.n651 B.n126 163.367
R864 B.n399 B.n303 163.367
R865 B.n399 B.n301 163.367
R866 B.n403 B.n301 163.367
R867 B.n403 B.n295 163.367
R868 B.n411 B.n295 163.367
R869 B.n411 B.n293 163.367
R870 B.n415 B.n293 163.367
R871 B.n415 B.n288 163.367
R872 B.n424 B.n288 163.367
R873 B.n424 B.n286 163.367
R874 B.n428 B.n286 163.367
R875 B.n428 B.n280 163.367
R876 B.n436 B.n280 163.367
R877 B.n436 B.n278 163.367
R878 B.n440 B.n278 163.367
R879 B.n440 B.n272 163.367
R880 B.n448 B.n272 163.367
R881 B.n448 B.n270 163.367
R882 B.n452 B.n270 163.367
R883 B.n452 B.n263 163.367
R884 B.n460 B.n263 163.367
R885 B.n460 B.n261 163.367
R886 B.n464 B.n261 163.367
R887 B.n464 B.n256 163.367
R888 B.n472 B.n256 163.367
R889 B.n472 B.n254 163.367
R890 B.n476 B.n254 163.367
R891 B.n476 B.n248 163.367
R892 B.n484 B.n248 163.367
R893 B.n484 B.n246 163.367
R894 B.n488 B.n246 163.367
R895 B.n488 B.n241 163.367
R896 B.n497 B.n241 163.367
R897 B.n497 B.n239 163.367
R898 B.n501 B.n239 163.367
R899 B.n501 B.n233 163.367
R900 B.n509 B.n233 163.367
R901 B.n509 B.n231 163.367
R902 B.n513 B.n231 163.367
R903 B.n513 B.n224 163.367
R904 B.n521 B.n224 163.367
R905 B.n521 B.n222 163.367
R906 B.n525 B.n222 163.367
R907 B.n525 B.n217 163.367
R908 B.n533 B.n217 163.367
R909 B.n533 B.n215 163.367
R910 B.n537 B.n215 163.367
R911 B.n537 B.n209 163.367
R912 B.n545 B.n209 163.367
R913 B.n545 B.n207 163.367
R914 B.n549 B.n207 163.367
R915 B.n549 B.n202 163.367
R916 B.n558 B.n202 163.367
R917 B.n558 B.n200 163.367
R918 B.n563 B.n200 163.367
R919 B.n563 B.n194 163.367
R920 B.n571 B.n194 163.367
R921 B.n572 B.n571 163.367
R922 B.n572 B.n5 163.367
R923 B.n6 B.n5 163.367
R924 B.n7 B.n6 163.367
R925 B.n578 B.n7 163.367
R926 B.n579 B.n578 163.367
R927 B.n579 B.n13 163.367
R928 B.n14 B.n13 163.367
R929 B.n15 B.n14 163.367
R930 B.n584 B.n15 163.367
R931 B.n584 B.n20 163.367
R932 B.n21 B.n20 163.367
R933 B.n22 B.n21 163.367
R934 B.n589 B.n22 163.367
R935 B.n589 B.n27 163.367
R936 B.n28 B.n27 163.367
R937 B.n29 B.n28 163.367
R938 B.n594 B.n29 163.367
R939 B.n594 B.n34 163.367
R940 B.n35 B.n34 163.367
R941 B.n36 B.n35 163.367
R942 B.n599 B.n36 163.367
R943 B.n599 B.n41 163.367
R944 B.n42 B.n41 163.367
R945 B.n43 B.n42 163.367
R946 B.n604 B.n43 163.367
R947 B.n604 B.n48 163.367
R948 B.n49 B.n48 163.367
R949 B.n50 B.n49 163.367
R950 B.n609 B.n50 163.367
R951 B.n609 B.n55 163.367
R952 B.n56 B.n55 163.367
R953 B.n57 B.n56 163.367
R954 B.n614 B.n57 163.367
R955 B.n614 B.n62 163.367
R956 B.n63 B.n62 163.367
R957 B.n64 B.n63 163.367
R958 B.n619 B.n64 163.367
R959 B.n619 B.n69 163.367
R960 B.n70 B.n69 163.367
R961 B.n71 B.n70 163.367
R962 B.n624 B.n71 163.367
R963 B.n624 B.n76 163.367
R964 B.n77 B.n76 163.367
R965 B.n78 B.n77 163.367
R966 B.n629 B.n78 163.367
R967 B.n629 B.n83 163.367
R968 B.n84 B.n83 163.367
R969 B.n85 B.n84 163.367
R970 B.n634 B.n85 163.367
R971 B.n634 B.n90 163.367
R972 B.n91 B.n90 163.367
R973 B.n92 B.n91 163.367
R974 B.n639 B.n92 163.367
R975 B.n639 B.n97 163.367
R976 B.n98 B.n97 163.367
R977 B.n99 B.n98 163.367
R978 B.n644 B.n99 163.367
R979 B.n644 B.n104 163.367
R980 B.n105 B.n104 163.367
R981 B.n106 B.n105 163.367
R982 B.n127 B.n106 163.367
R983 B.n390 B.n307 163.367
R984 B.n390 B.n323 163.367
R985 B.n386 B.n385 163.367
R986 B.n382 B.n381 163.367
R987 B.n378 B.n377 163.367
R988 B.n374 B.n373 163.367
R989 B.n369 B.n368 163.367
R990 B.n365 B.n364 163.367
R991 B.n361 B.n360 163.367
R992 B.n357 B.n356 163.367
R993 B.n353 B.n352 163.367
R994 B.n349 B.n348 163.367
R995 B.n345 B.n344 163.367
R996 B.n341 B.n340 163.367
R997 B.n337 B.n336 163.367
R998 B.n333 B.n332 163.367
R999 B.n397 B.n305 163.367
R1000 B.n397 B.n299 163.367
R1001 B.n405 B.n299 163.367
R1002 B.n405 B.n297 163.367
R1003 B.n409 B.n297 163.367
R1004 B.n409 B.n291 163.367
R1005 B.n418 B.n291 163.367
R1006 B.n418 B.n289 163.367
R1007 B.n422 B.n289 163.367
R1008 B.n422 B.n284 163.367
R1009 B.n430 B.n284 163.367
R1010 B.n430 B.n282 163.367
R1011 B.n434 B.n282 163.367
R1012 B.n434 B.n276 163.367
R1013 B.n442 B.n276 163.367
R1014 B.n442 B.n274 163.367
R1015 B.n446 B.n274 163.367
R1016 B.n446 B.n268 163.367
R1017 B.n454 B.n268 163.367
R1018 B.n454 B.n266 163.367
R1019 B.n458 B.n266 163.367
R1020 B.n458 B.n260 163.367
R1021 B.n466 B.n260 163.367
R1022 B.n466 B.n258 163.367
R1023 B.n470 B.n258 163.367
R1024 B.n470 B.n252 163.367
R1025 B.n478 B.n252 163.367
R1026 B.n478 B.n250 163.367
R1027 B.n482 B.n250 163.367
R1028 B.n482 B.n244 163.367
R1029 B.n491 B.n244 163.367
R1030 B.n491 B.n242 163.367
R1031 B.n495 B.n242 163.367
R1032 B.n495 B.n237 163.367
R1033 B.n503 B.n237 163.367
R1034 B.n503 B.n235 163.367
R1035 B.n507 B.n235 163.367
R1036 B.n507 B.n229 163.367
R1037 B.n515 B.n229 163.367
R1038 B.n515 B.n227 163.367
R1039 B.n519 B.n227 163.367
R1040 B.n519 B.n221 163.367
R1041 B.n527 B.n221 163.367
R1042 B.n527 B.n219 163.367
R1043 B.n531 B.n219 163.367
R1044 B.n531 B.n213 163.367
R1045 B.n539 B.n213 163.367
R1046 B.n539 B.n211 163.367
R1047 B.n543 B.n211 163.367
R1048 B.n543 B.n205 163.367
R1049 B.n552 B.n205 163.367
R1050 B.n552 B.n203 163.367
R1051 B.n556 B.n203 163.367
R1052 B.n556 B.n198 163.367
R1053 B.n565 B.n198 163.367
R1054 B.n565 B.n196 163.367
R1055 B.n569 B.n196 163.367
R1056 B.n569 B.n3 163.367
R1057 B.n775 B.n3 163.367
R1058 B.n771 B.n2 163.367
R1059 B.n771 B.n770 163.367
R1060 B.n770 B.n9 163.367
R1061 B.n766 B.n9 163.367
R1062 B.n766 B.n11 163.367
R1063 B.n762 B.n11 163.367
R1064 B.n762 B.n16 163.367
R1065 B.n758 B.n16 163.367
R1066 B.n758 B.n18 163.367
R1067 B.n754 B.n18 163.367
R1068 B.n754 B.n24 163.367
R1069 B.n750 B.n24 163.367
R1070 B.n750 B.n26 163.367
R1071 B.n746 B.n26 163.367
R1072 B.n746 B.n31 163.367
R1073 B.n742 B.n31 163.367
R1074 B.n742 B.n33 163.367
R1075 B.n738 B.n33 163.367
R1076 B.n738 B.n38 163.367
R1077 B.n734 B.n38 163.367
R1078 B.n734 B.n40 163.367
R1079 B.n730 B.n40 163.367
R1080 B.n730 B.n45 163.367
R1081 B.n726 B.n45 163.367
R1082 B.n726 B.n47 163.367
R1083 B.n722 B.n47 163.367
R1084 B.n722 B.n51 163.367
R1085 B.n718 B.n51 163.367
R1086 B.n718 B.n53 163.367
R1087 B.n714 B.n53 163.367
R1088 B.n714 B.n59 163.367
R1089 B.n710 B.n59 163.367
R1090 B.n710 B.n61 163.367
R1091 B.n706 B.n61 163.367
R1092 B.n706 B.n66 163.367
R1093 B.n702 B.n66 163.367
R1094 B.n702 B.n68 163.367
R1095 B.n698 B.n68 163.367
R1096 B.n698 B.n73 163.367
R1097 B.n694 B.n73 163.367
R1098 B.n694 B.n75 163.367
R1099 B.n690 B.n75 163.367
R1100 B.n690 B.n80 163.367
R1101 B.n686 B.n80 163.367
R1102 B.n686 B.n82 163.367
R1103 B.n682 B.n82 163.367
R1104 B.n682 B.n87 163.367
R1105 B.n678 B.n87 163.367
R1106 B.n678 B.n89 163.367
R1107 B.n674 B.n89 163.367
R1108 B.n674 B.n93 163.367
R1109 B.n670 B.n93 163.367
R1110 B.n670 B.n95 163.367
R1111 B.n666 B.n95 163.367
R1112 B.n666 B.n101 163.367
R1113 B.n662 B.n101 163.367
R1114 B.n662 B.n103 163.367
R1115 B.n658 B.n103 163.367
R1116 B.n658 B.n108 163.367
R1117 B.n129 B.t21 118.945
R1118 B.n327 B.t17 118.945
R1119 B.n131 B.t11 118.945
R1120 B.n325 B.t14 118.945
R1121 B.n398 B.n304 105.874
R1122 B.n398 B.n300 105.874
R1123 B.n404 B.n300 105.874
R1124 B.n404 B.n296 105.874
R1125 B.n410 B.n296 105.874
R1126 B.n410 B.n292 105.874
R1127 B.n417 B.n292 105.874
R1128 B.n417 B.n416 105.874
R1129 B.n423 B.n285 105.874
R1130 B.n429 B.n285 105.874
R1131 B.n429 B.n281 105.874
R1132 B.n435 B.n281 105.874
R1133 B.n435 B.n277 105.874
R1134 B.n441 B.n277 105.874
R1135 B.n441 B.n273 105.874
R1136 B.n447 B.n273 105.874
R1137 B.n447 B.n269 105.874
R1138 B.n453 B.n269 105.874
R1139 B.n453 B.n264 105.874
R1140 B.n459 B.n264 105.874
R1141 B.n459 B.n265 105.874
R1142 B.n465 B.n257 105.874
R1143 B.n471 B.n257 105.874
R1144 B.n471 B.n253 105.874
R1145 B.n477 B.n253 105.874
R1146 B.n477 B.n249 105.874
R1147 B.n483 B.n249 105.874
R1148 B.n483 B.n245 105.874
R1149 B.n490 B.n245 105.874
R1150 B.n490 B.n489 105.874
R1151 B.n496 B.n238 105.874
R1152 B.n502 B.n238 105.874
R1153 B.n502 B.n234 105.874
R1154 B.n508 B.n234 105.874
R1155 B.n508 B.n230 105.874
R1156 B.n514 B.n230 105.874
R1157 B.n514 B.n225 105.874
R1158 B.n520 B.n225 105.874
R1159 B.n520 B.n226 105.874
R1160 B.n526 B.n218 105.874
R1161 B.n532 B.n218 105.874
R1162 B.n532 B.n214 105.874
R1163 B.n538 B.n214 105.874
R1164 B.n538 B.n210 105.874
R1165 B.n544 B.n210 105.874
R1166 B.n544 B.n206 105.874
R1167 B.n551 B.n206 105.874
R1168 B.n551 B.n550 105.874
R1169 B.n557 B.n199 105.874
R1170 B.n564 B.n199 105.874
R1171 B.n564 B.n195 105.874
R1172 B.n570 B.n195 105.874
R1173 B.n570 B.n4 105.874
R1174 B.n774 B.n4 105.874
R1175 B.n774 B.n773 105.874
R1176 B.n773 B.n772 105.874
R1177 B.n772 B.n8 105.874
R1178 B.n12 B.n8 105.874
R1179 B.n765 B.n12 105.874
R1180 B.n765 B.n764 105.874
R1181 B.n764 B.n763 105.874
R1182 B.n757 B.n19 105.874
R1183 B.n757 B.n756 105.874
R1184 B.n756 B.n755 105.874
R1185 B.n755 B.n23 105.874
R1186 B.n749 B.n23 105.874
R1187 B.n749 B.n748 105.874
R1188 B.n748 B.n747 105.874
R1189 B.n747 B.n30 105.874
R1190 B.n741 B.n30 105.874
R1191 B.n740 B.n739 105.874
R1192 B.n739 B.n37 105.874
R1193 B.n733 B.n37 105.874
R1194 B.n733 B.n732 105.874
R1195 B.n732 B.n731 105.874
R1196 B.n731 B.n44 105.874
R1197 B.n725 B.n44 105.874
R1198 B.n725 B.n724 105.874
R1199 B.n724 B.n723 105.874
R1200 B.n717 B.n54 105.874
R1201 B.n717 B.n716 105.874
R1202 B.n716 B.n715 105.874
R1203 B.n715 B.n58 105.874
R1204 B.n709 B.n58 105.874
R1205 B.n709 B.n708 105.874
R1206 B.n708 B.n707 105.874
R1207 B.n707 B.n65 105.874
R1208 B.n701 B.n65 105.874
R1209 B.n700 B.n699 105.874
R1210 B.n699 B.n72 105.874
R1211 B.n693 B.n72 105.874
R1212 B.n693 B.n692 105.874
R1213 B.n692 B.n691 105.874
R1214 B.n691 B.n79 105.874
R1215 B.n685 B.n79 105.874
R1216 B.n685 B.n684 105.874
R1217 B.n684 B.n683 105.874
R1218 B.n683 B.n86 105.874
R1219 B.n677 B.n86 105.874
R1220 B.n677 B.n676 105.874
R1221 B.n676 B.n675 105.874
R1222 B.n669 B.n96 105.874
R1223 B.n669 B.n668 105.874
R1224 B.n668 B.n667 105.874
R1225 B.n667 B.n100 105.874
R1226 B.n661 B.n100 105.874
R1227 B.n661 B.n660 105.874
R1228 B.n660 B.n659 105.874
R1229 B.n659 B.n107 105.874
R1230 B.n465 B.t5 98.0897
R1231 B.n701 B.t2 98.0897
R1232 B.n550 B.t1 82.52
R1233 B.n19 B.t3 82.52
R1234 B.n496 B.t4 73.1781
R1235 B.n723 B.t6 73.1781
R1236 B.n654 B.n653 71.676
R1237 B.n133 B.n111 71.676
R1238 B.n137 B.n112 71.676
R1239 B.n141 B.n113 71.676
R1240 B.n145 B.n114 71.676
R1241 B.n149 B.n115 71.676
R1242 B.n153 B.n116 71.676
R1243 B.n157 B.n117 71.676
R1244 B.n161 B.n118 71.676
R1245 B.n165 B.n119 71.676
R1246 B.n169 B.n120 71.676
R1247 B.n174 B.n121 71.676
R1248 B.n178 B.n122 71.676
R1249 B.n182 B.n123 71.676
R1250 B.n186 B.n124 71.676
R1251 B.n190 B.n125 71.676
R1252 B.n126 B.n125 71.676
R1253 B.n189 B.n124 71.676
R1254 B.n185 B.n123 71.676
R1255 B.n181 B.n122 71.676
R1256 B.n177 B.n121 71.676
R1257 B.n173 B.n120 71.676
R1258 B.n168 B.n119 71.676
R1259 B.n164 B.n118 71.676
R1260 B.n160 B.n117 71.676
R1261 B.n156 B.n116 71.676
R1262 B.n152 B.n115 71.676
R1263 B.n148 B.n114 71.676
R1264 B.n144 B.n113 71.676
R1265 B.n140 B.n112 71.676
R1266 B.n136 B.n111 71.676
R1267 B.n653 B.n110 71.676
R1268 B.n393 B.n392 71.676
R1269 B.n323 B.n308 71.676
R1270 B.n385 B.n309 71.676
R1271 B.n381 B.n310 71.676
R1272 B.n377 B.n311 71.676
R1273 B.n373 B.n312 71.676
R1274 B.n368 B.n313 71.676
R1275 B.n364 B.n314 71.676
R1276 B.n360 B.n315 71.676
R1277 B.n356 B.n316 71.676
R1278 B.n352 B.n317 71.676
R1279 B.n348 B.n318 71.676
R1280 B.n344 B.n319 71.676
R1281 B.n340 B.n320 71.676
R1282 B.n336 B.n321 71.676
R1283 B.n332 B.n322 71.676
R1284 B.n392 B.n307 71.676
R1285 B.n386 B.n308 71.676
R1286 B.n382 B.n309 71.676
R1287 B.n378 B.n310 71.676
R1288 B.n374 B.n311 71.676
R1289 B.n369 B.n312 71.676
R1290 B.n365 B.n313 71.676
R1291 B.n361 B.n314 71.676
R1292 B.n357 B.n315 71.676
R1293 B.n353 B.n316 71.676
R1294 B.n349 B.n317 71.676
R1295 B.n345 B.n318 71.676
R1296 B.n341 B.n319 71.676
R1297 B.n337 B.n320 71.676
R1298 B.n333 B.n321 71.676
R1299 B.n329 B.n322 71.676
R1300 B.n776 B.n775 71.676
R1301 B.n776 B.n2 71.676
R1302 B.n131 B.n130 67.4914
R1303 B.n129 B.n128 67.4914
R1304 B.n327 B.n326 67.4914
R1305 B.n325 B.n324 67.4914
R1306 B.n416 B.t13 66.9503
R1307 B.n96 B.t9 66.9503
R1308 B.n132 B.n131 59.5399
R1309 B.n171 B.n129 59.5399
R1310 B.n328 B.n327 59.5399
R1311 B.n371 B.n325 59.5399
R1312 B.n226 B.t0 57.6084
R1313 B.t7 B.n740 57.6084
R1314 B.n526 B.t0 48.2666
R1315 B.n741 B.t7 48.2666
R1316 B.n423 B.t13 38.9248
R1317 B.n675 B.t9 38.9248
R1318 B.n489 B.t4 32.6969
R1319 B.n54 B.t6 32.6969
R1320 B.n395 B.n394 28.8785
R1321 B.n330 B.n302 28.8785
R1322 B.n656 B.n655 28.8785
R1323 B.n650 B.n649 28.8785
R1324 B.n557 B.t1 23.3551
R1325 B.n763 B.t3 23.3551
R1326 B B.n777 18.0485
R1327 B.n396 B.n395 10.6151
R1328 B.n396 B.n298 10.6151
R1329 B.n406 B.n298 10.6151
R1330 B.n407 B.n406 10.6151
R1331 B.n408 B.n407 10.6151
R1332 B.n408 B.n290 10.6151
R1333 B.n419 B.n290 10.6151
R1334 B.n420 B.n419 10.6151
R1335 B.n421 B.n420 10.6151
R1336 B.n421 B.n283 10.6151
R1337 B.n431 B.n283 10.6151
R1338 B.n432 B.n431 10.6151
R1339 B.n433 B.n432 10.6151
R1340 B.n433 B.n275 10.6151
R1341 B.n443 B.n275 10.6151
R1342 B.n444 B.n443 10.6151
R1343 B.n445 B.n444 10.6151
R1344 B.n445 B.n267 10.6151
R1345 B.n455 B.n267 10.6151
R1346 B.n456 B.n455 10.6151
R1347 B.n457 B.n456 10.6151
R1348 B.n457 B.n259 10.6151
R1349 B.n467 B.n259 10.6151
R1350 B.n468 B.n467 10.6151
R1351 B.n469 B.n468 10.6151
R1352 B.n469 B.n251 10.6151
R1353 B.n479 B.n251 10.6151
R1354 B.n480 B.n479 10.6151
R1355 B.n481 B.n480 10.6151
R1356 B.n481 B.n243 10.6151
R1357 B.n492 B.n243 10.6151
R1358 B.n493 B.n492 10.6151
R1359 B.n494 B.n493 10.6151
R1360 B.n494 B.n236 10.6151
R1361 B.n504 B.n236 10.6151
R1362 B.n505 B.n504 10.6151
R1363 B.n506 B.n505 10.6151
R1364 B.n506 B.n228 10.6151
R1365 B.n516 B.n228 10.6151
R1366 B.n517 B.n516 10.6151
R1367 B.n518 B.n517 10.6151
R1368 B.n518 B.n220 10.6151
R1369 B.n528 B.n220 10.6151
R1370 B.n529 B.n528 10.6151
R1371 B.n530 B.n529 10.6151
R1372 B.n530 B.n212 10.6151
R1373 B.n540 B.n212 10.6151
R1374 B.n541 B.n540 10.6151
R1375 B.n542 B.n541 10.6151
R1376 B.n542 B.n204 10.6151
R1377 B.n553 B.n204 10.6151
R1378 B.n554 B.n553 10.6151
R1379 B.n555 B.n554 10.6151
R1380 B.n555 B.n197 10.6151
R1381 B.n566 B.n197 10.6151
R1382 B.n567 B.n566 10.6151
R1383 B.n568 B.n567 10.6151
R1384 B.n568 B.n0 10.6151
R1385 B.n394 B.n306 10.6151
R1386 B.n389 B.n306 10.6151
R1387 B.n389 B.n388 10.6151
R1388 B.n388 B.n387 10.6151
R1389 B.n387 B.n384 10.6151
R1390 B.n384 B.n383 10.6151
R1391 B.n383 B.n380 10.6151
R1392 B.n380 B.n379 10.6151
R1393 B.n379 B.n376 10.6151
R1394 B.n376 B.n375 10.6151
R1395 B.n375 B.n372 10.6151
R1396 B.n370 B.n367 10.6151
R1397 B.n367 B.n366 10.6151
R1398 B.n366 B.n363 10.6151
R1399 B.n363 B.n362 10.6151
R1400 B.n362 B.n359 10.6151
R1401 B.n359 B.n358 10.6151
R1402 B.n358 B.n355 10.6151
R1403 B.n355 B.n354 10.6151
R1404 B.n351 B.n350 10.6151
R1405 B.n350 B.n347 10.6151
R1406 B.n347 B.n346 10.6151
R1407 B.n346 B.n343 10.6151
R1408 B.n343 B.n342 10.6151
R1409 B.n342 B.n339 10.6151
R1410 B.n339 B.n338 10.6151
R1411 B.n338 B.n335 10.6151
R1412 B.n335 B.n334 10.6151
R1413 B.n334 B.n331 10.6151
R1414 B.n331 B.n330 10.6151
R1415 B.n400 B.n302 10.6151
R1416 B.n401 B.n400 10.6151
R1417 B.n402 B.n401 10.6151
R1418 B.n402 B.n294 10.6151
R1419 B.n412 B.n294 10.6151
R1420 B.n413 B.n412 10.6151
R1421 B.n414 B.n413 10.6151
R1422 B.n414 B.n287 10.6151
R1423 B.n425 B.n287 10.6151
R1424 B.n426 B.n425 10.6151
R1425 B.n427 B.n426 10.6151
R1426 B.n427 B.n279 10.6151
R1427 B.n437 B.n279 10.6151
R1428 B.n438 B.n437 10.6151
R1429 B.n439 B.n438 10.6151
R1430 B.n439 B.n271 10.6151
R1431 B.n449 B.n271 10.6151
R1432 B.n450 B.n449 10.6151
R1433 B.n451 B.n450 10.6151
R1434 B.n451 B.n262 10.6151
R1435 B.n461 B.n262 10.6151
R1436 B.n462 B.n461 10.6151
R1437 B.n463 B.n462 10.6151
R1438 B.n463 B.n255 10.6151
R1439 B.n473 B.n255 10.6151
R1440 B.n474 B.n473 10.6151
R1441 B.n475 B.n474 10.6151
R1442 B.n475 B.n247 10.6151
R1443 B.n485 B.n247 10.6151
R1444 B.n486 B.n485 10.6151
R1445 B.n487 B.n486 10.6151
R1446 B.n487 B.n240 10.6151
R1447 B.n498 B.n240 10.6151
R1448 B.n499 B.n498 10.6151
R1449 B.n500 B.n499 10.6151
R1450 B.n500 B.n232 10.6151
R1451 B.n510 B.n232 10.6151
R1452 B.n511 B.n510 10.6151
R1453 B.n512 B.n511 10.6151
R1454 B.n512 B.n223 10.6151
R1455 B.n522 B.n223 10.6151
R1456 B.n523 B.n522 10.6151
R1457 B.n524 B.n523 10.6151
R1458 B.n524 B.n216 10.6151
R1459 B.n534 B.n216 10.6151
R1460 B.n535 B.n534 10.6151
R1461 B.n536 B.n535 10.6151
R1462 B.n536 B.n208 10.6151
R1463 B.n546 B.n208 10.6151
R1464 B.n547 B.n546 10.6151
R1465 B.n548 B.n547 10.6151
R1466 B.n548 B.n201 10.6151
R1467 B.n559 B.n201 10.6151
R1468 B.n560 B.n559 10.6151
R1469 B.n562 B.n560 10.6151
R1470 B.n562 B.n561 10.6151
R1471 B.n561 B.n193 10.6151
R1472 B.n573 B.n193 10.6151
R1473 B.n574 B.n573 10.6151
R1474 B.n575 B.n574 10.6151
R1475 B.n576 B.n575 10.6151
R1476 B.n577 B.n576 10.6151
R1477 B.n580 B.n577 10.6151
R1478 B.n581 B.n580 10.6151
R1479 B.n582 B.n581 10.6151
R1480 B.n583 B.n582 10.6151
R1481 B.n585 B.n583 10.6151
R1482 B.n586 B.n585 10.6151
R1483 B.n587 B.n586 10.6151
R1484 B.n588 B.n587 10.6151
R1485 B.n590 B.n588 10.6151
R1486 B.n591 B.n590 10.6151
R1487 B.n592 B.n591 10.6151
R1488 B.n593 B.n592 10.6151
R1489 B.n595 B.n593 10.6151
R1490 B.n596 B.n595 10.6151
R1491 B.n597 B.n596 10.6151
R1492 B.n598 B.n597 10.6151
R1493 B.n600 B.n598 10.6151
R1494 B.n601 B.n600 10.6151
R1495 B.n602 B.n601 10.6151
R1496 B.n603 B.n602 10.6151
R1497 B.n605 B.n603 10.6151
R1498 B.n606 B.n605 10.6151
R1499 B.n607 B.n606 10.6151
R1500 B.n608 B.n607 10.6151
R1501 B.n610 B.n608 10.6151
R1502 B.n611 B.n610 10.6151
R1503 B.n612 B.n611 10.6151
R1504 B.n613 B.n612 10.6151
R1505 B.n615 B.n613 10.6151
R1506 B.n616 B.n615 10.6151
R1507 B.n617 B.n616 10.6151
R1508 B.n618 B.n617 10.6151
R1509 B.n620 B.n618 10.6151
R1510 B.n621 B.n620 10.6151
R1511 B.n622 B.n621 10.6151
R1512 B.n623 B.n622 10.6151
R1513 B.n625 B.n623 10.6151
R1514 B.n626 B.n625 10.6151
R1515 B.n627 B.n626 10.6151
R1516 B.n628 B.n627 10.6151
R1517 B.n630 B.n628 10.6151
R1518 B.n631 B.n630 10.6151
R1519 B.n632 B.n631 10.6151
R1520 B.n633 B.n632 10.6151
R1521 B.n635 B.n633 10.6151
R1522 B.n636 B.n635 10.6151
R1523 B.n637 B.n636 10.6151
R1524 B.n638 B.n637 10.6151
R1525 B.n640 B.n638 10.6151
R1526 B.n641 B.n640 10.6151
R1527 B.n642 B.n641 10.6151
R1528 B.n643 B.n642 10.6151
R1529 B.n645 B.n643 10.6151
R1530 B.n646 B.n645 10.6151
R1531 B.n647 B.n646 10.6151
R1532 B.n648 B.n647 10.6151
R1533 B.n649 B.n648 10.6151
R1534 B.n769 B.n1 10.6151
R1535 B.n769 B.n768 10.6151
R1536 B.n768 B.n767 10.6151
R1537 B.n767 B.n10 10.6151
R1538 B.n761 B.n10 10.6151
R1539 B.n761 B.n760 10.6151
R1540 B.n760 B.n759 10.6151
R1541 B.n759 B.n17 10.6151
R1542 B.n753 B.n17 10.6151
R1543 B.n753 B.n752 10.6151
R1544 B.n752 B.n751 10.6151
R1545 B.n751 B.n25 10.6151
R1546 B.n745 B.n25 10.6151
R1547 B.n745 B.n744 10.6151
R1548 B.n744 B.n743 10.6151
R1549 B.n743 B.n32 10.6151
R1550 B.n737 B.n32 10.6151
R1551 B.n737 B.n736 10.6151
R1552 B.n736 B.n735 10.6151
R1553 B.n735 B.n39 10.6151
R1554 B.n729 B.n39 10.6151
R1555 B.n729 B.n728 10.6151
R1556 B.n728 B.n727 10.6151
R1557 B.n727 B.n46 10.6151
R1558 B.n721 B.n46 10.6151
R1559 B.n721 B.n720 10.6151
R1560 B.n720 B.n719 10.6151
R1561 B.n719 B.n52 10.6151
R1562 B.n713 B.n52 10.6151
R1563 B.n713 B.n712 10.6151
R1564 B.n712 B.n711 10.6151
R1565 B.n711 B.n60 10.6151
R1566 B.n705 B.n60 10.6151
R1567 B.n705 B.n704 10.6151
R1568 B.n704 B.n703 10.6151
R1569 B.n703 B.n67 10.6151
R1570 B.n697 B.n67 10.6151
R1571 B.n697 B.n696 10.6151
R1572 B.n696 B.n695 10.6151
R1573 B.n695 B.n74 10.6151
R1574 B.n689 B.n74 10.6151
R1575 B.n689 B.n688 10.6151
R1576 B.n688 B.n687 10.6151
R1577 B.n687 B.n81 10.6151
R1578 B.n681 B.n81 10.6151
R1579 B.n681 B.n680 10.6151
R1580 B.n680 B.n679 10.6151
R1581 B.n679 B.n88 10.6151
R1582 B.n673 B.n88 10.6151
R1583 B.n673 B.n672 10.6151
R1584 B.n672 B.n671 10.6151
R1585 B.n671 B.n94 10.6151
R1586 B.n665 B.n94 10.6151
R1587 B.n665 B.n664 10.6151
R1588 B.n664 B.n663 10.6151
R1589 B.n663 B.n102 10.6151
R1590 B.n657 B.n102 10.6151
R1591 B.n657 B.n656 10.6151
R1592 B.n655 B.n109 10.6151
R1593 B.n134 B.n109 10.6151
R1594 B.n135 B.n134 10.6151
R1595 B.n138 B.n135 10.6151
R1596 B.n139 B.n138 10.6151
R1597 B.n142 B.n139 10.6151
R1598 B.n143 B.n142 10.6151
R1599 B.n146 B.n143 10.6151
R1600 B.n147 B.n146 10.6151
R1601 B.n150 B.n147 10.6151
R1602 B.n151 B.n150 10.6151
R1603 B.n155 B.n154 10.6151
R1604 B.n158 B.n155 10.6151
R1605 B.n159 B.n158 10.6151
R1606 B.n162 B.n159 10.6151
R1607 B.n163 B.n162 10.6151
R1608 B.n166 B.n163 10.6151
R1609 B.n167 B.n166 10.6151
R1610 B.n170 B.n167 10.6151
R1611 B.n175 B.n172 10.6151
R1612 B.n176 B.n175 10.6151
R1613 B.n179 B.n176 10.6151
R1614 B.n180 B.n179 10.6151
R1615 B.n183 B.n180 10.6151
R1616 B.n184 B.n183 10.6151
R1617 B.n187 B.n184 10.6151
R1618 B.n188 B.n187 10.6151
R1619 B.n191 B.n188 10.6151
R1620 B.n192 B.n191 10.6151
R1621 B.n650 B.n192 10.6151
R1622 B.n777 B.n0 8.11757
R1623 B.n777 B.n1 8.11757
R1624 B.n265 B.t5 7.78535
R1625 B.t2 B.n700 7.78535
R1626 B.n371 B.n370 6.5566
R1627 B.n354 B.n328 6.5566
R1628 B.n154 B.n132 6.5566
R1629 B.n171 B.n170 6.5566
R1630 B.n372 B.n371 4.05904
R1631 B.n351 B.n328 4.05904
R1632 B.n151 B.n132 4.05904
R1633 B.n172 B.n171 4.05904
R1634 VN.n60 VN.n59 161.3
R1635 VN.n58 VN.n32 161.3
R1636 VN.n57 VN.n56 161.3
R1637 VN.n55 VN.n33 161.3
R1638 VN.n54 VN.n53 161.3
R1639 VN.n52 VN.n34 161.3
R1640 VN.n51 VN.n50 161.3
R1641 VN.n49 VN.n48 161.3
R1642 VN.n47 VN.n36 161.3
R1643 VN.n46 VN.n45 161.3
R1644 VN.n44 VN.n37 161.3
R1645 VN.n43 VN.n42 161.3
R1646 VN.n41 VN.n38 161.3
R1647 VN.n29 VN.n28 161.3
R1648 VN.n27 VN.n1 161.3
R1649 VN.n26 VN.n25 161.3
R1650 VN.n24 VN.n2 161.3
R1651 VN.n23 VN.n22 161.3
R1652 VN.n21 VN.n3 161.3
R1653 VN.n20 VN.n19 161.3
R1654 VN.n18 VN.n17 161.3
R1655 VN.n16 VN.n5 161.3
R1656 VN.n15 VN.n14 161.3
R1657 VN.n13 VN.n6 161.3
R1658 VN.n12 VN.n11 161.3
R1659 VN.n10 VN.n7 161.3
R1660 VN.n30 VN.n0 67.0684
R1661 VN.n61 VN.n31 67.0684
R1662 VN.n15 VN.n6 56.5193
R1663 VN.n26 VN.n2 56.5193
R1664 VN.n46 VN.n37 56.5193
R1665 VN.n57 VN.n33 56.5193
R1666 VN.n40 VN.n39 50.0328
R1667 VN.n9 VN.n8 50.0328
R1668 VN.n8 VN.t4 47.0994
R1669 VN.n39 VN.t6 47.0993
R1670 VN VN.n61 46.1041
R1671 VN.n11 VN.n10 24.4675
R1672 VN.n11 VN.n6 24.4675
R1673 VN.n16 VN.n15 24.4675
R1674 VN.n17 VN.n16 24.4675
R1675 VN.n21 VN.n20 24.4675
R1676 VN.n22 VN.n21 24.4675
R1677 VN.n22 VN.n2 24.4675
R1678 VN.n27 VN.n26 24.4675
R1679 VN.n28 VN.n27 24.4675
R1680 VN.n42 VN.n37 24.4675
R1681 VN.n42 VN.n41 24.4675
R1682 VN.n53 VN.n33 24.4675
R1683 VN.n53 VN.n52 24.4675
R1684 VN.n52 VN.n51 24.4675
R1685 VN.n48 VN.n47 24.4675
R1686 VN.n47 VN.n46 24.4675
R1687 VN.n59 VN.n58 24.4675
R1688 VN.n58 VN.n57 24.4675
R1689 VN.n10 VN.n9 23.9782
R1690 VN.n17 VN.n4 23.9782
R1691 VN.n41 VN.n40 23.9782
R1692 VN.n48 VN.n35 23.9782
R1693 VN.n28 VN.n0 22.9995
R1694 VN.n59 VN.n31 22.9995
R1695 VN.n9 VN.t5 13.6954
R1696 VN.n4 VN.t0 13.6954
R1697 VN.n0 VN.t2 13.6954
R1698 VN.n40 VN.t7 13.6954
R1699 VN.n35 VN.t3 13.6954
R1700 VN.n31 VN.t1 13.6954
R1701 VN.n39 VN.n38 3.77031
R1702 VN.n8 VN.n7 3.77031
R1703 VN.n20 VN.n4 0.48984
R1704 VN.n51 VN.n35 0.48984
R1705 VN.n61 VN.n60 0.354971
R1706 VN.n30 VN.n29 0.354971
R1707 VN VN.n30 0.26696
R1708 VN.n60 VN.n32 0.189894
R1709 VN.n56 VN.n32 0.189894
R1710 VN.n56 VN.n55 0.189894
R1711 VN.n55 VN.n54 0.189894
R1712 VN.n54 VN.n34 0.189894
R1713 VN.n50 VN.n34 0.189894
R1714 VN.n50 VN.n49 0.189894
R1715 VN.n49 VN.n36 0.189894
R1716 VN.n45 VN.n36 0.189894
R1717 VN.n45 VN.n44 0.189894
R1718 VN.n44 VN.n43 0.189894
R1719 VN.n43 VN.n38 0.189894
R1720 VN.n12 VN.n7 0.189894
R1721 VN.n13 VN.n12 0.189894
R1722 VN.n14 VN.n13 0.189894
R1723 VN.n14 VN.n5 0.189894
R1724 VN.n18 VN.n5 0.189894
R1725 VN.n19 VN.n18 0.189894
R1726 VN.n19 VN.n3 0.189894
R1727 VN.n23 VN.n3 0.189894
R1728 VN.n24 VN.n23 0.189894
R1729 VN.n25 VN.n24 0.189894
R1730 VN.n25 VN.n1 0.189894
R1731 VN.n29 VN.n1 0.189894
R1732 VDD2.n2 VDD2.n1 103.061
R1733 VDD2.n2 VDD2.n0 103.061
R1734 VDD2 VDD2.n5 103.058
R1735 VDD2.n4 VDD2.n3 101.618
R1736 VDD2.n4 VDD2.n2 38.7584
R1737 VDD2.n5 VDD2.t0 11.062
R1738 VDD2.n5 VDD2.t1 11.062
R1739 VDD2.n3 VDD2.t6 11.062
R1740 VDD2.n3 VDD2.t4 11.062
R1741 VDD2.n1 VDD2.t7 11.062
R1742 VDD2.n1 VDD2.t5 11.062
R1743 VDD2.n0 VDD2.t3 11.062
R1744 VDD2.n0 VDD2.t2 11.062
R1745 VDD2 VDD2.n4 1.55869
C0 VN VP 6.45018f
C1 VTAIL VP 3.15574f
C2 VDD1 VP 2.16254f
C3 VTAIL VN 3.14163f
C4 VDD1 VN 0.158902f
C5 VDD2 VP 0.585815f
C6 VDD1 VTAIL 5.1496f
C7 VDD2 VN 1.73912f
C8 VDD2 VTAIL 5.20771f
C9 VDD2 VDD1 2.0648f
C10 VDD2 B 5.077915f
C11 VDD1 B 5.77898f
C12 VTAIL B 4.182696f
C13 VN B 16.65725f
C14 VP B 15.277349f
C15 VDD2.t3 B 0.035752f
C16 VDD2.t2 B 0.035752f
C17 VDD2.n0 B 0.236532f
C18 VDD2.t7 B 0.035752f
C19 VDD2.t5 B 0.035752f
C20 VDD2.n1 B 0.236532f
C21 VDD2.n2 B 2.94875f
C22 VDD2.t6 B 0.035752f
C23 VDD2.t4 B 0.035752f
C24 VDD2.n3 B 0.228848f
C25 VDD2.n4 B 2.34256f
C26 VDD2.t0 B 0.035752f
C27 VDD2.t1 B 0.035752f
C28 VDD2.n5 B 0.236509f
C29 VN.t2 B 0.317849f
C30 VN.n0 B 0.260431f
C31 VN.n1 B 0.024718f
C32 VN.n2 B 0.034706f
C33 VN.n3 B 0.024718f
C34 VN.t0 B 0.317849f
C35 VN.n4 B 0.152938f
C36 VN.n5 B 0.024718f
C37 VN.n6 B 0.036084f
C38 VN.n7 B 0.281182f
C39 VN.t5 B 0.317849f
C40 VN.t4 B 0.554945f
C41 VN.n8 B 0.244892f
C42 VN.n9 B 0.246106f
C43 VN.n10 B 0.045613f
C44 VN.n11 B 0.046068f
C45 VN.n12 B 0.024718f
C46 VN.n13 B 0.024718f
C47 VN.n14 B 0.024718f
C48 VN.n15 B 0.036084f
C49 VN.n16 B 0.046068f
C50 VN.n17 B 0.045613f
C51 VN.n18 B 0.024718f
C52 VN.n19 B 0.024718f
C53 VN.n20 B 0.023779f
C54 VN.n21 B 0.046068f
C55 VN.n22 B 0.046068f
C56 VN.n23 B 0.024718f
C57 VN.n24 B 0.024718f
C58 VN.n25 B 0.024718f
C59 VN.n26 B 0.037461f
C60 VN.n27 B 0.046068f
C61 VN.n28 B 0.044703f
C62 VN.n29 B 0.039894f
C63 VN.n30 B 0.048876f
C64 VN.t1 B 0.317849f
C65 VN.n31 B 0.260431f
C66 VN.n32 B 0.024718f
C67 VN.n33 B 0.034706f
C68 VN.n34 B 0.024718f
C69 VN.t3 B 0.317849f
C70 VN.n35 B 0.152938f
C71 VN.n36 B 0.024718f
C72 VN.n37 B 0.036084f
C73 VN.n38 B 0.281182f
C74 VN.t7 B 0.317849f
C75 VN.t6 B 0.554945f
C76 VN.n39 B 0.244892f
C77 VN.n40 B 0.246106f
C78 VN.n41 B 0.045613f
C79 VN.n42 B 0.046068f
C80 VN.n43 B 0.024718f
C81 VN.n44 B 0.024718f
C82 VN.n45 B 0.024718f
C83 VN.n46 B 0.036084f
C84 VN.n47 B 0.046068f
C85 VN.n48 B 0.045613f
C86 VN.n49 B 0.024718f
C87 VN.n50 B 0.024718f
C88 VN.n51 B 0.023779f
C89 VN.n52 B 0.046068f
C90 VN.n53 B 0.046068f
C91 VN.n54 B 0.024718f
C92 VN.n55 B 0.024718f
C93 VN.n56 B 0.024718f
C94 VN.n57 B 0.037461f
C95 VN.n58 B 0.046068f
C96 VN.n59 B 0.044703f
C97 VN.n60 B 0.039894f
C98 VN.n61 B 1.24316f
C99 VTAIL.t7 B 0.047771f
C100 VTAIL.t6 B 0.047771f
C101 VTAIL.n0 B 0.260958f
C102 VTAIL.n1 B 0.566423f
C103 VTAIL.n2 B 0.044508f
C104 VTAIL.n3 B 0.104299f
C105 VTAIL.t3 B 0.074726f
C106 VTAIL.n4 B 0.076898f
C107 VTAIL.n5 B 0.022357f
C108 VTAIL.n6 B 0.018148f
C109 VTAIL.n7 B 0.20358f
C110 VTAIL.n8 B 0.048641f
C111 VTAIL.n9 B 0.409306f
C112 VTAIL.n10 B 0.044508f
C113 VTAIL.n11 B 0.104299f
C114 VTAIL.t12 B 0.074726f
C115 VTAIL.n12 B 0.076898f
C116 VTAIL.n13 B 0.022357f
C117 VTAIL.n14 B 0.018148f
C118 VTAIL.n15 B 0.20358f
C119 VTAIL.n16 B 0.048641f
C120 VTAIL.n17 B 0.409306f
C121 VTAIL.t9 B 0.047771f
C122 VTAIL.t10 B 0.047771f
C123 VTAIL.n18 B 0.260958f
C124 VTAIL.n19 B 0.886556f
C125 VTAIL.n20 B 0.044508f
C126 VTAIL.n21 B 0.104299f
C127 VTAIL.t11 B 0.074726f
C128 VTAIL.n22 B 0.076898f
C129 VTAIL.n23 B 0.022357f
C130 VTAIL.n24 B 0.018148f
C131 VTAIL.n25 B 0.20358f
C132 VTAIL.n26 B 0.048641f
C133 VTAIL.n27 B 1.31132f
C134 VTAIL.n28 B 0.044508f
C135 VTAIL.n29 B 0.104299f
C136 VTAIL.t5 B 0.074726f
C137 VTAIL.n30 B 0.076898f
C138 VTAIL.n31 B 0.022357f
C139 VTAIL.n32 B 0.018148f
C140 VTAIL.n33 B 0.20358f
C141 VTAIL.n34 B 0.048641f
C142 VTAIL.n35 B 1.31132f
C143 VTAIL.t4 B 0.047771f
C144 VTAIL.t0 B 0.047771f
C145 VTAIL.n36 B 0.26096f
C146 VTAIL.n37 B 0.886555f
C147 VTAIL.n38 B 0.044508f
C148 VTAIL.n39 B 0.104299f
C149 VTAIL.t1 B 0.074726f
C150 VTAIL.n40 B 0.076898f
C151 VTAIL.n41 B 0.022357f
C152 VTAIL.n42 B 0.018148f
C153 VTAIL.n43 B 0.20358f
C154 VTAIL.n44 B 0.048641f
C155 VTAIL.n45 B 0.409306f
C156 VTAIL.n46 B 0.044508f
C157 VTAIL.n47 B 0.104299f
C158 VTAIL.t8 B 0.074726f
C159 VTAIL.n48 B 0.076898f
C160 VTAIL.n49 B 0.022357f
C161 VTAIL.n50 B 0.018148f
C162 VTAIL.n51 B 0.20358f
C163 VTAIL.n52 B 0.048641f
C164 VTAIL.n53 B 0.409306f
C165 VTAIL.t14 B 0.047771f
C166 VTAIL.t15 B 0.047771f
C167 VTAIL.n54 B 0.26096f
C168 VTAIL.n55 B 0.886555f
C169 VTAIL.n56 B 0.044508f
C170 VTAIL.n57 B 0.104299f
C171 VTAIL.t13 B 0.074726f
C172 VTAIL.n58 B 0.076898f
C173 VTAIL.n59 B 0.022357f
C174 VTAIL.n60 B 0.018148f
C175 VTAIL.n61 B 0.20358f
C176 VTAIL.n62 B 0.048641f
C177 VTAIL.n63 B 1.31132f
C178 VTAIL.n64 B 0.044508f
C179 VTAIL.n65 B 0.104299f
C180 VTAIL.t2 B 0.074726f
C181 VTAIL.n66 B 0.076898f
C182 VTAIL.n67 B 0.022357f
C183 VTAIL.n68 B 0.018148f
C184 VTAIL.n69 B 0.20358f
C185 VTAIL.n70 B 0.048641f
C186 VTAIL.n71 B 1.30499f
C187 VDD1.t7 B 0.045455f
C188 VDD1.t6 B 0.045455f
C189 VDD1.n0 B 0.301657f
C190 VDD1.t5 B 0.045455f
C191 VDD1.t2 B 0.045455f
C192 VDD1.n1 B 0.30073f
C193 VDD1.t1 B 0.045455f
C194 VDD1.t4 B 0.045455f
C195 VDD1.n2 B 0.30073f
C196 VDD1.n3 B 3.8159f
C197 VDD1.t0 B 0.045455f
C198 VDD1.t3 B 0.045455f
C199 VDD1.n4 B 0.29096f
C200 VDD1.n5 B 3.01819f
C201 VP.t3 B 0.395431f
C202 VP.n0 B 0.323999f
C203 VP.n1 B 0.030751f
C204 VP.n2 B 0.043177f
C205 VP.n3 B 0.030751f
C206 VP.t5 B 0.395431f
C207 VP.n4 B 0.190268f
C208 VP.n5 B 0.030751f
C209 VP.n6 B 0.044891f
C210 VP.n7 B 0.030751f
C211 VP.t6 B 0.395431f
C212 VP.n8 B 0.057312f
C213 VP.n9 B 0.030751f
C214 VP.n10 B 0.057312f
C215 VP.t2 B 0.395431f
C216 VP.n11 B 0.323999f
C217 VP.n12 B 0.030751f
C218 VP.n13 B 0.043177f
C219 VP.n14 B 0.030751f
C220 VP.t0 B 0.395431f
C221 VP.n15 B 0.190268f
C222 VP.n16 B 0.030751f
C223 VP.n17 B 0.044891f
C224 VP.n18 B 0.349815f
C225 VP.t1 B 0.395431f
C226 VP.t7 B 0.690398f
C227 VP.n19 B 0.304667f
C228 VP.n20 B 0.306178f
C229 VP.n21 B 0.056746f
C230 VP.n22 B 0.057312f
C231 VP.n23 B 0.030751f
C232 VP.n24 B 0.030751f
C233 VP.n25 B 0.030751f
C234 VP.n26 B 0.044891f
C235 VP.n27 B 0.057312f
C236 VP.n28 B 0.056746f
C237 VP.n29 B 0.030751f
C238 VP.n30 B 0.030751f
C239 VP.n31 B 0.029583f
C240 VP.n32 B 0.057312f
C241 VP.n33 B 0.057312f
C242 VP.n34 B 0.030751f
C243 VP.n35 B 0.030751f
C244 VP.n36 B 0.030751f
C245 VP.n37 B 0.046605f
C246 VP.n38 B 0.057312f
C247 VP.n39 B 0.055614f
C248 VP.n40 B 0.049632f
C249 VP.n41 B 1.53364f
C250 VP.n42 B 1.55771f
C251 VP.t4 B 0.395431f
C252 VP.n43 B 0.323999f
C253 VP.n44 B 0.055614f
C254 VP.n45 B 0.049632f
C255 VP.n46 B 0.030751f
C256 VP.n47 B 0.030751f
C257 VP.n48 B 0.046605f
C258 VP.n49 B 0.043177f
C259 VP.n50 B 0.057312f
C260 VP.n51 B 0.030751f
C261 VP.n52 B 0.030751f
C262 VP.n53 B 0.030751f
C263 VP.n54 B 0.029583f
C264 VP.n55 B 0.190268f
C265 VP.n56 B 0.056746f
C266 VP.n57 B 0.057312f
C267 VP.n58 B 0.030751f
C268 VP.n59 B 0.030751f
C269 VP.n60 B 0.030751f
C270 VP.n61 B 0.044891f
C271 VP.n62 B 0.057312f
C272 VP.n63 B 0.056746f
C273 VP.n64 B 0.030751f
C274 VP.n65 B 0.030751f
C275 VP.n66 B 0.029583f
C276 VP.n67 B 0.057312f
C277 VP.n68 B 0.057312f
C278 VP.n69 B 0.030751f
C279 VP.n70 B 0.030751f
C280 VP.n71 B 0.030751f
C281 VP.n72 B 0.046605f
C282 VP.n73 B 0.057312f
C283 VP.n74 B 0.055614f
C284 VP.n75 B 0.049632f
C285 VP.n76 B 0.060806f
.ends

