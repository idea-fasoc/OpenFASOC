* NGSPICE file created from diff_pair_sample_1720.ext - technology: sky130A

.subckt diff_pair_sample_1720 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=1.89585 pd=11.82 as=4.4811 ps=23.76 w=11.49 l=0.33
X1 VDD2.t3 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.89585 pd=11.82 as=4.4811 ps=23.76 w=11.49 l=0.33
X2 VTAIL.t3 VN.t1 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=4.4811 pd=23.76 as=1.89585 ps=11.82 w=11.49 l=0.33
X3 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=4.4811 pd=23.76 as=0 ps=0 w=11.49 l=0.33
X4 VTAIL.t0 VN.t2 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=4.4811 pd=23.76 as=1.89585 ps=11.82 w=11.49 l=0.33
X5 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=4.4811 pd=23.76 as=0 ps=0 w=11.49 l=0.33
X6 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.4811 pd=23.76 as=0 ps=0 w=11.49 l=0.33
X7 VTAIL.t4 VP.t1 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=4.4811 pd=23.76 as=1.89585 ps=11.82 w=11.49 l=0.33
X8 VTAIL.t6 VP.t2 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=4.4811 pd=23.76 as=1.89585 ps=11.82 w=11.49 l=0.33
X9 VDD2.t0 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.89585 pd=11.82 as=4.4811 ps=23.76 w=11.49 l=0.33
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=4.4811 pd=23.76 as=0 ps=0 w=11.49 l=0.33
X11 VDD1.t0 VP.t3 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.89585 pd=11.82 as=4.4811 ps=23.76 w=11.49 l=0.33
R0 VP.n1 VP.t3 982.989
R1 VP.n1 VP.t1 982.989
R2 VP.n0 VP.t2 982.989
R3 VP.n0 VP.t0 982.989
R4 VP.n2 VP.n0 200.315
R5 VP.n2 VP.n1 161.3
R6 VP VP.n2 0.0516364
R7 VTAIL.n490 VTAIL.n434 289.615
R8 VTAIL.n56 VTAIL.n0 289.615
R9 VTAIL.n118 VTAIL.n62 289.615
R10 VTAIL.n180 VTAIL.n124 289.615
R11 VTAIL.n428 VTAIL.n372 289.615
R12 VTAIL.n366 VTAIL.n310 289.615
R13 VTAIL.n304 VTAIL.n248 289.615
R14 VTAIL.n242 VTAIL.n186 289.615
R15 VTAIL.n455 VTAIL.n454 185
R16 VTAIL.n457 VTAIL.n456 185
R17 VTAIL.n450 VTAIL.n449 185
R18 VTAIL.n463 VTAIL.n462 185
R19 VTAIL.n465 VTAIL.n464 185
R20 VTAIL.n446 VTAIL.n445 185
R21 VTAIL.n472 VTAIL.n471 185
R22 VTAIL.n473 VTAIL.n444 185
R23 VTAIL.n475 VTAIL.n474 185
R24 VTAIL.n442 VTAIL.n441 185
R25 VTAIL.n481 VTAIL.n480 185
R26 VTAIL.n483 VTAIL.n482 185
R27 VTAIL.n438 VTAIL.n437 185
R28 VTAIL.n489 VTAIL.n488 185
R29 VTAIL.n491 VTAIL.n490 185
R30 VTAIL.n21 VTAIL.n20 185
R31 VTAIL.n23 VTAIL.n22 185
R32 VTAIL.n16 VTAIL.n15 185
R33 VTAIL.n29 VTAIL.n28 185
R34 VTAIL.n31 VTAIL.n30 185
R35 VTAIL.n12 VTAIL.n11 185
R36 VTAIL.n38 VTAIL.n37 185
R37 VTAIL.n39 VTAIL.n10 185
R38 VTAIL.n41 VTAIL.n40 185
R39 VTAIL.n8 VTAIL.n7 185
R40 VTAIL.n47 VTAIL.n46 185
R41 VTAIL.n49 VTAIL.n48 185
R42 VTAIL.n4 VTAIL.n3 185
R43 VTAIL.n55 VTAIL.n54 185
R44 VTAIL.n57 VTAIL.n56 185
R45 VTAIL.n83 VTAIL.n82 185
R46 VTAIL.n85 VTAIL.n84 185
R47 VTAIL.n78 VTAIL.n77 185
R48 VTAIL.n91 VTAIL.n90 185
R49 VTAIL.n93 VTAIL.n92 185
R50 VTAIL.n74 VTAIL.n73 185
R51 VTAIL.n100 VTAIL.n99 185
R52 VTAIL.n101 VTAIL.n72 185
R53 VTAIL.n103 VTAIL.n102 185
R54 VTAIL.n70 VTAIL.n69 185
R55 VTAIL.n109 VTAIL.n108 185
R56 VTAIL.n111 VTAIL.n110 185
R57 VTAIL.n66 VTAIL.n65 185
R58 VTAIL.n117 VTAIL.n116 185
R59 VTAIL.n119 VTAIL.n118 185
R60 VTAIL.n145 VTAIL.n144 185
R61 VTAIL.n147 VTAIL.n146 185
R62 VTAIL.n140 VTAIL.n139 185
R63 VTAIL.n153 VTAIL.n152 185
R64 VTAIL.n155 VTAIL.n154 185
R65 VTAIL.n136 VTAIL.n135 185
R66 VTAIL.n162 VTAIL.n161 185
R67 VTAIL.n163 VTAIL.n134 185
R68 VTAIL.n165 VTAIL.n164 185
R69 VTAIL.n132 VTAIL.n131 185
R70 VTAIL.n171 VTAIL.n170 185
R71 VTAIL.n173 VTAIL.n172 185
R72 VTAIL.n128 VTAIL.n127 185
R73 VTAIL.n179 VTAIL.n178 185
R74 VTAIL.n181 VTAIL.n180 185
R75 VTAIL.n429 VTAIL.n428 185
R76 VTAIL.n427 VTAIL.n426 185
R77 VTAIL.n376 VTAIL.n375 185
R78 VTAIL.n421 VTAIL.n420 185
R79 VTAIL.n419 VTAIL.n418 185
R80 VTAIL.n380 VTAIL.n379 185
R81 VTAIL.n384 VTAIL.n382 185
R82 VTAIL.n413 VTAIL.n412 185
R83 VTAIL.n411 VTAIL.n410 185
R84 VTAIL.n386 VTAIL.n385 185
R85 VTAIL.n405 VTAIL.n404 185
R86 VTAIL.n403 VTAIL.n402 185
R87 VTAIL.n390 VTAIL.n389 185
R88 VTAIL.n397 VTAIL.n396 185
R89 VTAIL.n395 VTAIL.n394 185
R90 VTAIL.n367 VTAIL.n366 185
R91 VTAIL.n365 VTAIL.n364 185
R92 VTAIL.n314 VTAIL.n313 185
R93 VTAIL.n359 VTAIL.n358 185
R94 VTAIL.n357 VTAIL.n356 185
R95 VTAIL.n318 VTAIL.n317 185
R96 VTAIL.n322 VTAIL.n320 185
R97 VTAIL.n351 VTAIL.n350 185
R98 VTAIL.n349 VTAIL.n348 185
R99 VTAIL.n324 VTAIL.n323 185
R100 VTAIL.n343 VTAIL.n342 185
R101 VTAIL.n341 VTAIL.n340 185
R102 VTAIL.n328 VTAIL.n327 185
R103 VTAIL.n335 VTAIL.n334 185
R104 VTAIL.n333 VTAIL.n332 185
R105 VTAIL.n305 VTAIL.n304 185
R106 VTAIL.n303 VTAIL.n302 185
R107 VTAIL.n252 VTAIL.n251 185
R108 VTAIL.n297 VTAIL.n296 185
R109 VTAIL.n295 VTAIL.n294 185
R110 VTAIL.n256 VTAIL.n255 185
R111 VTAIL.n260 VTAIL.n258 185
R112 VTAIL.n289 VTAIL.n288 185
R113 VTAIL.n287 VTAIL.n286 185
R114 VTAIL.n262 VTAIL.n261 185
R115 VTAIL.n281 VTAIL.n280 185
R116 VTAIL.n279 VTAIL.n278 185
R117 VTAIL.n266 VTAIL.n265 185
R118 VTAIL.n273 VTAIL.n272 185
R119 VTAIL.n271 VTAIL.n270 185
R120 VTAIL.n243 VTAIL.n242 185
R121 VTAIL.n241 VTAIL.n240 185
R122 VTAIL.n190 VTAIL.n189 185
R123 VTAIL.n235 VTAIL.n234 185
R124 VTAIL.n233 VTAIL.n232 185
R125 VTAIL.n194 VTAIL.n193 185
R126 VTAIL.n198 VTAIL.n196 185
R127 VTAIL.n227 VTAIL.n226 185
R128 VTAIL.n225 VTAIL.n224 185
R129 VTAIL.n200 VTAIL.n199 185
R130 VTAIL.n219 VTAIL.n218 185
R131 VTAIL.n217 VTAIL.n216 185
R132 VTAIL.n204 VTAIL.n203 185
R133 VTAIL.n211 VTAIL.n210 185
R134 VTAIL.n209 VTAIL.n208 185
R135 VTAIL.n453 VTAIL.t1 149.524
R136 VTAIL.n19 VTAIL.t3 149.524
R137 VTAIL.n81 VTAIL.t5 149.524
R138 VTAIL.n143 VTAIL.t4 149.524
R139 VTAIL.n393 VTAIL.t7 149.524
R140 VTAIL.n331 VTAIL.t6 149.524
R141 VTAIL.n269 VTAIL.t2 149.524
R142 VTAIL.n207 VTAIL.t0 149.524
R143 VTAIL.n456 VTAIL.n455 104.615
R144 VTAIL.n456 VTAIL.n449 104.615
R145 VTAIL.n463 VTAIL.n449 104.615
R146 VTAIL.n464 VTAIL.n463 104.615
R147 VTAIL.n464 VTAIL.n445 104.615
R148 VTAIL.n472 VTAIL.n445 104.615
R149 VTAIL.n473 VTAIL.n472 104.615
R150 VTAIL.n474 VTAIL.n473 104.615
R151 VTAIL.n474 VTAIL.n441 104.615
R152 VTAIL.n481 VTAIL.n441 104.615
R153 VTAIL.n482 VTAIL.n481 104.615
R154 VTAIL.n482 VTAIL.n437 104.615
R155 VTAIL.n489 VTAIL.n437 104.615
R156 VTAIL.n490 VTAIL.n489 104.615
R157 VTAIL.n22 VTAIL.n21 104.615
R158 VTAIL.n22 VTAIL.n15 104.615
R159 VTAIL.n29 VTAIL.n15 104.615
R160 VTAIL.n30 VTAIL.n29 104.615
R161 VTAIL.n30 VTAIL.n11 104.615
R162 VTAIL.n38 VTAIL.n11 104.615
R163 VTAIL.n39 VTAIL.n38 104.615
R164 VTAIL.n40 VTAIL.n39 104.615
R165 VTAIL.n40 VTAIL.n7 104.615
R166 VTAIL.n47 VTAIL.n7 104.615
R167 VTAIL.n48 VTAIL.n47 104.615
R168 VTAIL.n48 VTAIL.n3 104.615
R169 VTAIL.n55 VTAIL.n3 104.615
R170 VTAIL.n56 VTAIL.n55 104.615
R171 VTAIL.n84 VTAIL.n83 104.615
R172 VTAIL.n84 VTAIL.n77 104.615
R173 VTAIL.n91 VTAIL.n77 104.615
R174 VTAIL.n92 VTAIL.n91 104.615
R175 VTAIL.n92 VTAIL.n73 104.615
R176 VTAIL.n100 VTAIL.n73 104.615
R177 VTAIL.n101 VTAIL.n100 104.615
R178 VTAIL.n102 VTAIL.n101 104.615
R179 VTAIL.n102 VTAIL.n69 104.615
R180 VTAIL.n109 VTAIL.n69 104.615
R181 VTAIL.n110 VTAIL.n109 104.615
R182 VTAIL.n110 VTAIL.n65 104.615
R183 VTAIL.n117 VTAIL.n65 104.615
R184 VTAIL.n118 VTAIL.n117 104.615
R185 VTAIL.n146 VTAIL.n145 104.615
R186 VTAIL.n146 VTAIL.n139 104.615
R187 VTAIL.n153 VTAIL.n139 104.615
R188 VTAIL.n154 VTAIL.n153 104.615
R189 VTAIL.n154 VTAIL.n135 104.615
R190 VTAIL.n162 VTAIL.n135 104.615
R191 VTAIL.n163 VTAIL.n162 104.615
R192 VTAIL.n164 VTAIL.n163 104.615
R193 VTAIL.n164 VTAIL.n131 104.615
R194 VTAIL.n171 VTAIL.n131 104.615
R195 VTAIL.n172 VTAIL.n171 104.615
R196 VTAIL.n172 VTAIL.n127 104.615
R197 VTAIL.n179 VTAIL.n127 104.615
R198 VTAIL.n180 VTAIL.n179 104.615
R199 VTAIL.n428 VTAIL.n427 104.615
R200 VTAIL.n427 VTAIL.n375 104.615
R201 VTAIL.n420 VTAIL.n375 104.615
R202 VTAIL.n420 VTAIL.n419 104.615
R203 VTAIL.n419 VTAIL.n379 104.615
R204 VTAIL.n384 VTAIL.n379 104.615
R205 VTAIL.n412 VTAIL.n384 104.615
R206 VTAIL.n412 VTAIL.n411 104.615
R207 VTAIL.n411 VTAIL.n385 104.615
R208 VTAIL.n404 VTAIL.n385 104.615
R209 VTAIL.n404 VTAIL.n403 104.615
R210 VTAIL.n403 VTAIL.n389 104.615
R211 VTAIL.n396 VTAIL.n389 104.615
R212 VTAIL.n396 VTAIL.n395 104.615
R213 VTAIL.n366 VTAIL.n365 104.615
R214 VTAIL.n365 VTAIL.n313 104.615
R215 VTAIL.n358 VTAIL.n313 104.615
R216 VTAIL.n358 VTAIL.n357 104.615
R217 VTAIL.n357 VTAIL.n317 104.615
R218 VTAIL.n322 VTAIL.n317 104.615
R219 VTAIL.n350 VTAIL.n322 104.615
R220 VTAIL.n350 VTAIL.n349 104.615
R221 VTAIL.n349 VTAIL.n323 104.615
R222 VTAIL.n342 VTAIL.n323 104.615
R223 VTAIL.n342 VTAIL.n341 104.615
R224 VTAIL.n341 VTAIL.n327 104.615
R225 VTAIL.n334 VTAIL.n327 104.615
R226 VTAIL.n334 VTAIL.n333 104.615
R227 VTAIL.n304 VTAIL.n303 104.615
R228 VTAIL.n303 VTAIL.n251 104.615
R229 VTAIL.n296 VTAIL.n251 104.615
R230 VTAIL.n296 VTAIL.n295 104.615
R231 VTAIL.n295 VTAIL.n255 104.615
R232 VTAIL.n260 VTAIL.n255 104.615
R233 VTAIL.n288 VTAIL.n260 104.615
R234 VTAIL.n288 VTAIL.n287 104.615
R235 VTAIL.n287 VTAIL.n261 104.615
R236 VTAIL.n280 VTAIL.n261 104.615
R237 VTAIL.n280 VTAIL.n279 104.615
R238 VTAIL.n279 VTAIL.n265 104.615
R239 VTAIL.n272 VTAIL.n265 104.615
R240 VTAIL.n272 VTAIL.n271 104.615
R241 VTAIL.n242 VTAIL.n241 104.615
R242 VTAIL.n241 VTAIL.n189 104.615
R243 VTAIL.n234 VTAIL.n189 104.615
R244 VTAIL.n234 VTAIL.n233 104.615
R245 VTAIL.n233 VTAIL.n193 104.615
R246 VTAIL.n198 VTAIL.n193 104.615
R247 VTAIL.n226 VTAIL.n198 104.615
R248 VTAIL.n226 VTAIL.n225 104.615
R249 VTAIL.n225 VTAIL.n199 104.615
R250 VTAIL.n218 VTAIL.n199 104.615
R251 VTAIL.n218 VTAIL.n217 104.615
R252 VTAIL.n217 VTAIL.n203 104.615
R253 VTAIL.n210 VTAIL.n203 104.615
R254 VTAIL.n210 VTAIL.n209 104.615
R255 VTAIL.n455 VTAIL.t1 52.3082
R256 VTAIL.n21 VTAIL.t3 52.3082
R257 VTAIL.n83 VTAIL.t5 52.3082
R258 VTAIL.n145 VTAIL.t4 52.3082
R259 VTAIL.n395 VTAIL.t7 52.3082
R260 VTAIL.n333 VTAIL.t6 52.3082
R261 VTAIL.n271 VTAIL.t2 52.3082
R262 VTAIL.n209 VTAIL.t0 52.3082
R263 VTAIL.n495 VTAIL.n494 33.9308
R264 VTAIL.n61 VTAIL.n60 33.9308
R265 VTAIL.n123 VTAIL.n122 33.9308
R266 VTAIL.n185 VTAIL.n184 33.9308
R267 VTAIL.n433 VTAIL.n432 33.9308
R268 VTAIL.n371 VTAIL.n370 33.9308
R269 VTAIL.n309 VTAIL.n308 33.9308
R270 VTAIL.n247 VTAIL.n246 33.9308
R271 VTAIL.n495 VTAIL.n433 22.8583
R272 VTAIL.n247 VTAIL.n185 22.8583
R273 VTAIL.n475 VTAIL.n442 13.1884
R274 VTAIL.n41 VTAIL.n8 13.1884
R275 VTAIL.n103 VTAIL.n70 13.1884
R276 VTAIL.n165 VTAIL.n132 13.1884
R277 VTAIL.n382 VTAIL.n380 13.1884
R278 VTAIL.n320 VTAIL.n318 13.1884
R279 VTAIL.n258 VTAIL.n256 13.1884
R280 VTAIL.n196 VTAIL.n194 13.1884
R281 VTAIL.n476 VTAIL.n444 12.8005
R282 VTAIL.n480 VTAIL.n479 12.8005
R283 VTAIL.n42 VTAIL.n10 12.8005
R284 VTAIL.n46 VTAIL.n45 12.8005
R285 VTAIL.n104 VTAIL.n72 12.8005
R286 VTAIL.n108 VTAIL.n107 12.8005
R287 VTAIL.n166 VTAIL.n134 12.8005
R288 VTAIL.n170 VTAIL.n169 12.8005
R289 VTAIL.n418 VTAIL.n417 12.8005
R290 VTAIL.n414 VTAIL.n413 12.8005
R291 VTAIL.n356 VTAIL.n355 12.8005
R292 VTAIL.n352 VTAIL.n351 12.8005
R293 VTAIL.n294 VTAIL.n293 12.8005
R294 VTAIL.n290 VTAIL.n289 12.8005
R295 VTAIL.n232 VTAIL.n231 12.8005
R296 VTAIL.n228 VTAIL.n227 12.8005
R297 VTAIL.n471 VTAIL.n470 12.0247
R298 VTAIL.n483 VTAIL.n440 12.0247
R299 VTAIL.n37 VTAIL.n36 12.0247
R300 VTAIL.n49 VTAIL.n6 12.0247
R301 VTAIL.n99 VTAIL.n98 12.0247
R302 VTAIL.n111 VTAIL.n68 12.0247
R303 VTAIL.n161 VTAIL.n160 12.0247
R304 VTAIL.n173 VTAIL.n130 12.0247
R305 VTAIL.n421 VTAIL.n378 12.0247
R306 VTAIL.n410 VTAIL.n383 12.0247
R307 VTAIL.n359 VTAIL.n316 12.0247
R308 VTAIL.n348 VTAIL.n321 12.0247
R309 VTAIL.n297 VTAIL.n254 12.0247
R310 VTAIL.n286 VTAIL.n259 12.0247
R311 VTAIL.n235 VTAIL.n192 12.0247
R312 VTAIL.n224 VTAIL.n197 12.0247
R313 VTAIL.n469 VTAIL.n446 11.249
R314 VTAIL.n484 VTAIL.n438 11.249
R315 VTAIL.n35 VTAIL.n12 11.249
R316 VTAIL.n50 VTAIL.n4 11.249
R317 VTAIL.n97 VTAIL.n74 11.249
R318 VTAIL.n112 VTAIL.n66 11.249
R319 VTAIL.n159 VTAIL.n136 11.249
R320 VTAIL.n174 VTAIL.n128 11.249
R321 VTAIL.n422 VTAIL.n376 11.249
R322 VTAIL.n409 VTAIL.n386 11.249
R323 VTAIL.n360 VTAIL.n314 11.249
R324 VTAIL.n347 VTAIL.n324 11.249
R325 VTAIL.n298 VTAIL.n252 11.249
R326 VTAIL.n285 VTAIL.n262 11.249
R327 VTAIL.n236 VTAIL.n190 11.249
R328 VTAIL.n223 VTAIL.n200 11.249
R329 VTAIL.n466 VTAIL.n465 10.4732
R330 VTAIL.n488 VTAIL.n487 10.4732
R331 VTAIL.n32 VTAIL.n31 10.4732
R332 VTAIL.n54 VTAIL.n53 10.4732
R333 VTAIL.n94 VTAIL.n93 10.4732
R334 VTAIL.n116 VTAIL.n115 10.4732
R335 VTAIL.n156 VTAIL.n155 10.4732
R336 VTAIL.n178 VTAIL.n177 10.4732
R337 VTAIL.n426 VTAIL.n425 10.4732
R338 VTAIL.n406 VTAIL.n405 10.4732
R339 VTAIL.n364 VTAIL.n363 10.4732
R340 VTAIL.n344 VTAIL.n343 10.4732
R341 VTAIL.n302 VTAIL.n301 10.4732
R342 VTAIL.n282 VTAIL.n281 10.4732
R343 VTAIL.n240 VTAIL.n239 10.4732
R344 VTAIL.n220 VTAIL.n219 10.4732
R345 VTAIL.n454 VTAIL.n453 10.2747
R346 VTAIL.n20 VTAIL.n19 10.2747
R347 VTAIL.n82 VTAIL.n81 10.2747
R348 VTAIL.n144 VTAIL.n143 10.2747
R349 VTAIL.n394 VTAIL.n393 10.2747
R350 VTAIL.n332 VTAIL.n331 10.2747
R351 VTAIL.n270 VTAIL.n269 10.2747
R352 VTAIL.n208 VTAIL.n207 10.2747
R353 VTAIL.n462 VTAIL.n448 9.69747
R354 VTAIL.n491 VTAIL.n436 9.69747
R355 VTAIL.n28 VTAIL.n14 9.69747
R356 VTAIL.n57 VTAIL.n2 9.69747
R357 VTAIL.n90 VTAIL.n76 9.69747
R358 VTAIL.n119 VTAIL.n64 9.69747
R359 VTAIL.n152 VTAIL.n138 9.69747
R360 VTAIL.n181 VTAIL.n126 9.69747
R361 VTAIL.n429 VTAIL.n374 9.69747
R362 VTAIL.n402 VTAIL.n388 9.69747
R363 VTAIL.n367 VTAIL.n312 9.69747
R364 VTAIL.n340 VTAIL.n326 9.69747
R365 VTAIL.n305 VTAIL.n250 9.69747
R366 VTAIL.n278 VTAIL.n264 9.69747
R367 VTAIL.n243 VTAIL.n188 9.69747
R368 VTAIL.n216 VTAIL.n202 9.69747
R369 VTAIL.n494 VTAIL.n493 9.45567
R370 VTAIL.n60 VTAIL.n59 9.45567
R371 VTAIL.n122 VTAIL.n121 9.45567
R372 VTAIL.n184 VTAIL.n183 9.45567
R373 VTAIL.n432 VTAIL.n431 9.45567
R374 VTAIL.n370 VTAIL.n369 9.45567
R375 VTAIL.n308 VTAIL.n307 9.45567
R376 VTAIL.n246 VTAIL.n245 9.45567
R377 VTAIL.n493 VTAIL.n492 9.3005
R378 VTAIL.n436 VTAIL.n435 9.3005
R379 VTAIL.n487 VTAIL.n486 9.3005
R380 VTAIL.n485 VTAIL.n484 9.3005
R381 VTAIL.n440 VTAIL.n439 9.3005
R382 VTAIL.n479 VTAIL.n478 9.3005
R383 VTAIL.n452 VTAIL.n451 9.3005
R384 VTAIL.n459 VTAIL.n458 9.3005
R385 VTAIL.n461 VTAIL.n460 9.3005
R386 VTAIL.n448 VTAIL.n447 9.3005
R387 VTAIL.n467 VTAIL.n466 9.3005
R388 VTAIL.n469 VTAIL.n468 9.3005
R389 VTAIL.n470 VTAIL.n443 9.3005
R390 VTAIL.n477 VTAIL.n476 9.3005
R391 VTAIL.n59 VTAIL.n58 9.3005
R392 VTAIL.n2 VTAIL.n1 9.3005
R393 VTAIL.n53 VTAIL.n52 9.3005
R394 VTAIL.n51 VTAIL.n50 9.3005
R395 VTAIL.n6 VTAIL.n5 9.3005
R396 VTAIL.n45 VTAIL.n44 9.3005
R397 VTAIL.n18 VTAIL.n17 9.3005
R398 VTAIL.n25 VTAIL.n24 9.3005
R399 VTAIL.n27 VTAIL.n26 9.3005
R400 VTAIL.n14 VTAIL.n13 9.3005
R401 VTAIL.n33 VTAIL.n32 9.3005
R402 VTAIL.n35 VTAIL.n34 9.3005
R403 VTAIL.n36 VTAIL.n9 9.3005
R404 VTAIL.n43 VTAIL.n42 9.3005
R405 VTAIL.n121 VTAIL.n120 9.3005
R406 VTAIL.n64 VTAIL.n63 9.3005
R407 VTAIL.n115 VTAIL.n114 9.3005
R408 VTAIL.n113 VTAIL.n112 9.3005
R409 VTAIL.n68 VTAIL.n67 9.3005
R410 VTAIL.n107 VTAIL.n106 9.3005
R411 VTAIL.n80 VTAIL.n79 9.3005
R412 VTAIL.n87 VTAIL.n86 9.3005
R413 VTAIL.n89 VTAIL.n88 9.3005
R414 VTAIL.n76 VTAIL.n75 9.3005
R415 VTAIL.n95 VTAIL.n94 9.3005
R416 VTAIL.n97 VTAIL.n96 9.3005
R417 VTAIL.n98 VTAIL.n71 9.3005
R418 VTAIL.n105 VTAIL.n104 9.3005
R419 VTAIL.n183 VTAIL.n182 9.3005
R420 VTAIL.n126 VTAIL.n125 9.3005
R421 VTAIL.n177 VTAIL.n176 9.3005
R422 VTAIL.n175 VTAIL.n174 9.3005
R423 VTAIL.n130 VTAIL.n129 9.3005
R424 VTAIL.n169 VTAIL.n168 9.3005
R425 VTAIL.n142 VTAIL.n141 9.3005
R426 VTAIL.n149 VTAIL.n148 9.3005
R427 VTAIL.n151 VTAIL.n150 9.3005
R428 VTAIL.n138 VTAIL.n137 9.3005
R429 VTAIL.n157 VTAIL.n156 9.3005
R430 VTAIL.n159 VTAIL.n158 9.3005
R431 VTAIL.n160 VTAIL.n133 9.3005
R432 VTAIL.n167 VTAIL.n166 9.3005
R433 VTAIL.n392 VTAIL.n391 9.3005
R434 VTAIL.n399 VTAIL.n398 9.3005
R435 VTAIL.n401 VTAIL.n400 9.3005
R436 VTAIL.n388 VTAIL.n387 9.3005
R437 VTAIL.n407 VTAIL.n406 9.3005
R438 VTAIL.n409 VTAIL.n408 9.3005
R439 VTAIL.n383 VTAIL.n381 9.3005
R440 VTAIL.n415 VTAIL.n414 9.3005
R441 VTAIL.n431 VTAIL.n430 9.3005
R442 VTAIL.n374 VTAIL.n373 9.3005
R443 VTAIL.n425 VTAIL.n424 9.3005
R444 VTAIL.n423 VTAIL.n422 9.3005
R445 VTAIL.n378 VTAIL.n377 9.3005
R446 VTAIL.n417 VTAIL.n416 9.3005
R447 VTAIL.n330 VTAIL.n329 9.3005
R448 VTAIL.n337 VTAIL.n336 9.3005
R449 VTAIL.n339 VTAIL.n338 9.3005
R450 VTAIL.n326 VTAIL.n325 9.3005
R451 VTAIL.n345 VTAIL.n344 9.3005
R452 VTAIL.n347 VTAIL.n346 9.3005
R453 VTAIL.n321 VTAIL.n319 9.3005
R454 VTAIL.n353 VTAIL.n352 9.3005
R455 VTAIL.n369 VTAIL.n368 9.3005
R456 VTAIL.n312 VTAIL.n311 9.3005
R457 VTAIL.n363 VTAIL.n362 9.3005
R458 VTAIL.n361 VTAIL.n360 9.3005
R459 VTAIL.n316 VTAIL.n315 9.3005
R460 VTAIL.n355 VTAIL.n354 9.3005
R461 VTAIL.n268 VTAIL.n267 9.3005
R462 VTAIL.n275 VTAIL.n274 9.3005
R463 VTAIL.n277 VTAIL.n276 9.3005
R464 VTAIL.n264 VTAIL.n263 9.3005
R465 VTAIL.n283 VTAIL.n282 9.3005
R466 VTAIL.n285 VTAIL.n284 9.3005
R467 VTAIL.n259 VTAIL.n257 9.3005
R468 VTAIL.n291 VTAIL.n290 9.3005
R469 VTAIL.n307 VTAIL.n306 9.3005
R470 VTAIL.n250 VTAIL.n249 9.3005
R471 VTAIL.n301 VTAIL.n300 9.3005
R472 VTAIL.n299 VTAIL.n298 9.3005
R473 VTAIL.n254 VTAIL.n253 9.3005
R474 VTAIL.n293 VTAIL.n292 9.3005
R475 VTAIL.n206 VTAIL.n205 9.3005
R476 VTAIL.n213 VTAIL.n212 9.3005
R477 VTAIL.n215 VTAIL.n214 9.3005
R478 VTAIL.n202 VTAIL.n201 9.3005
R479 VTAIL.n221 VTAIL.n220 9.3005
R480 VTAIL.n223 VTAIL.n222 9.3005
R481 VTAIL.n197 VTAIL.n195 9.3005
R482 VTAIL.n229 VTAIL.n228 9.3005
R483 VTAIL.n245 VTAIL.n244 9.3005
R484 VTAIL.n188 VTAIL.n187 9.3005
R485 VTAIL.n239 VTAIL.n238 9.3005
R486 VTAIL.n237 VTAIL.n236 9.3005
R487 VTAIL.n192 VTAIL.n191 9.3005
R488 VTAIL.n231 VTAIL.n230 9.3005
R489 VTAIL.n461 VTAIL.n450 8.92171
R490 VTAIL.n492 VTAIL.n434 8.92171
R491 VTAIL.n27 VTAIL.n16 8.92171
R492 VTAIL.n58 VTAIL.n0 8.92171
R493 VTAIL.n89 VTAIL.n78 8.92171
R494 VTAIL.n120 VTAIL.n62 8.92171
R495 VTAIL.n151 VTAIL.n140 8.92171
R496 VTAIL.n182 VTAIL.n124 8.92171
R497 VTAIL.n430 VTAIL.n372 8.92171
R498 VTAIL.n401 VTAIL.n390 8.92171
R499 VTAIL.n368 VTAIL.n310 8.92171
R500 VTAIL.n339 VTAIL.n328 8.92171
R501 VTAIL.n306 VTAIL.n248 8.92171
R502 VTAIL.n277 VTAIL.n266 8.92171
R503 VTAIL.n244 VTAIL.n186 8.92171
R504 VTAIL.n215 VTAIL.n204 8.92171
R505 VTAIL.n458 VTAIL.n457 8.14595
R506 VTAIL.n24 VTAIL.n23 8.14595
R507 VTAIL.n86 VTAIL.n85 8.14595
R508 VTAIL.n148 VTAIL.n147 8.14595
R509 VTAIL.n398 VTAIL.n397 8.14595
R510 VTAIL.n336 VTAIL.n335 8.14595
R511 VTAIL.n274 VTAIL.n273 8.14595
R512 VTAIL.n212 VTAIL.n211 8.14595
R513 VTAIL.n454 VTAIL.n452 7.3702
R514 VTAIL.n20 VTAIL.n18 7.3702
R515 VTAIL.n82 VTAIL.n80 7.3702
R516 VTAIL.n144 VTAIL.n142 7.3702
R517 VTAIL.n394 VTAIL.n392 7.3702
R518 VTAIL.n332 VTAIL.n330 7.3702
R519 VTAIL.n270 VTAIL.n268 7.3702
R520 VTAIL.n208 VTAIL.n206 7.3702
R521 VTAIL.n457 VTAIL.n452 5.81868
R522 VTAIL.n23 VTAIL.n18 5.81868
R523 VTAIL.n85 VTAIL.n80 5.81868
R524 VTAIL.n147 VTAIL.n142 5.81868
R525 VTAIL.n397 VTAIL.n392 5.81868
R526 VTAIL.n335 VTAIL.n330 5.81868
R527 VTAIL.n273 VTAIL.n268 5.81868
R528 VTAIL.n211 VTAIL.n206 5.81868
R529 VTAIL.n458 VTAIL.n450 5.04292
R530 VTAIL.n494 VTAIL.n434 5.04292
R531 VTAIL.n24 VTAIL.n16 5.04292
R532 VTAIL.n60 VTAIL.n0 5.04292
R533 VTAIL.n86 VTAIL.n78 5.04292
R534 VTAIL.n122 VTAIL.n62 5.04292
R535 VTAIL.n148 VTAIL.n140 5.04292
R536 VTAIL.n184 VTAIL.n124 5.04292
R537 VTAIL.n432 VTAIL.n372 5.04292
R538 VTAIL.n398 VTAIL.n390 5.04292
R539 VTAIL.n370 VTAIL.n310 5.04292
R540 VTAIL.n336 VTAIL.n328 5.04292
R541 VTAIL.n308 VTAIL.n248 5.04292
R542 VTAIL.n274 VTAIL.n266 5.04292
R543 VTAIL.n246 VTAIL.n186 5.04292
R544 VTAIL.n212 VTAIL.n204 5.04292
R545 VTAIL.n462 VTAIL.n461 4.26717
R546 VTAIL.n492 VTAIL.n491 4.26717
R547 VTAIL.n28 VTAIL.n27 4.26717
R548 VTAIL.n58 VTAIL.n57 4.26717
R549 VTAIL.n90 VTAIL.n89 4.26717
R550 VTAIL.n120 VTAIL.n119 4.26717
R551 VTAIL.n152 VTAIL.n151 4.26717
R552 VTAIL.n182 VTAIL.n181 4.26717
R553 VTAIL.n430 VTAIL.n429 4.26717
R554 VTAIL.n402 VTAIL.n401 4.26717
R555 VTAIL.n368 VTAIL.n367 4.26717
R556 VTAIL.n340 VTAIL.n339 4.26717
R557 VTAIL.n306 VTAIL.n305 4.26717
R558 VTAIL.n278 VTAIL.n277 4.26717
R559 VTAIL.n244 VTAIL.n243 4.26717
R560 VTAIL.n216 VTAIL.n215 4.26717
R561 VTAIL.n465 VTAIL.n448 3.49141
R562 VTAIL.n488 VTAIL.n436 3.49141
R563 VTAIL.n31 VTAIL.n14 3.49141
R564 VTAIL.n54 VTAIL.n2 3.49141
R565 VTAIL.n93 VTAIL.n76 3.49141
R566 VTAIL.n116 VTAIL.n64 3.49141
R567 VTAIL.n155 VTAIL.n138 3.49141
R568 VTAIL.n178 VTAIL.n126 3.49141
R569 VTAIL.n426 VTAIL.n374 3.49141
R570 VTAIL.n405 VTAIL.n388 3.49141
R571 VTAIL.n364 VTAIL.n312 3.49141
R572 VTAIL.n343 VTAIL.n326 3.49141
R573 VTAIL.n302 VTAIL.n250 3.49141
R574 VTAIL.n281 VTAIL.n264 3.49141
R575 VTAIL.n240 VTAIL.n188 3.49141
R576 VTAIL.n219 VTAIL.n202 3.49141
R577 VTAIL.n453 VTAIL.n451 2.84303
R578 VTAIL.n19 VTAIL.n17 2.84303
R579 VTAIL.n81 VTAIL.n79 2.84303
R580 VTAIL.n143 VTAIL.n141 2.84303
R581 VTAIL.n393 VTAIL.n391 2.84303
R582 VTAIL.n331 VTAIL.n329 2.84303
R583 VTAIL.n269 VTAIL.n267 2.84303
R584 VTAIL.n207 VTAIL.n205 2.84303
R585 VTAIL.n466 VTAIL.n446 2.71565
R586 VTAIL.n487 VTAIL.n438 2.71565
R587 VTAIL.n32 VTAIL.n12 2.71565
R588 VTAIL.n53 VTAIL.n4 2.71565
R589 VTAIL.n94 VTAIL.n74 2.71565
R590 VTAIL.n115 VTAIL.n66 2.71565
R591 VTAIL.n156 VTAIL.n136 2.71565
R592 VTAIL.n177 VTAIL.n128 2.71565
R593 VTAIL.n425 VTAIL.n376 2.71565
R594 VTAIL.n406 VTAIL.n386 2.71565
R595 VTAIL.n363 VTAIL.n314 2.71565
R596 VTAIL.n344 VTAIL.n324 2.71565
R597 VTAIL.n301 VTAIL.n252 2.71565
R598 VTAIL.n282 VTAIL.n262 2.71565
R599 VTAIL.n239 VTAIL.n190 2.71565
R600 VTAIL.n220 VTAIL.n200 2.71565
R601 VTAIL.n471 VTAIL.n469 1.93989
R602 VTAIL.n484 VTAIL.n483 1.93989
R603 VTAIL.n37 VTAIL.n35 1.93989
R604 VTAIL.n50 VTAIL.n49 1.93989
R605 VTAIL.n99 VTAIL.n97 1.93989
R606 VTAIL.n112 VTAIL.n111 1.93989
R607 VTAIL.n161 VTAIL.n159 1.93989
R608 VTAIL.n174 VTAIL.n173 1.93989
R609 VTAIL.n422 VTAIL.n421 1.93989
R610 VTAIL.n410 VTAIL.n409 1.93989
R611 VTAIL.n360 VTAIL.n359 1.93989
R612 VTAIL.n348 VTAIL.n347 1.93989
R613 VTAIL.n298 VTAIL.n297 1.93989
R614 VTAIL.n286 VTAIL.n285 1.93989
R615 VTAIL.n236 VTAIL.n235 1.93989
R616 VTAIL.n224 VTAIL.n223 1.93989
R617 VTAIL.n470 VTAIL.n444 1.16414
R618 VTAIL.n480 VTAIL.n440 1.16414
R619 VTAIL.n36 VTAIL.n10 1.16414
R620 VTAIL.n46 VTAIL.n6 1.16414
R621 VTAIL.n98 VTAIL.n72 1.16414
R622 VTAIL.n108 VTAIL.n68 1.16414
R623 VTAIL.n160 VTAIL.n134 1.16414
R624 VTAIL.n170 VTAIL.n130 1.16414
R625 VTAIL.n418 VTAIL.n378 1.16414
R626 VTAIL.n413 VTAIL.n383 1.16414
R627 VTAIL.n356 VTAIL.n316 1.16414
R628 VTAIL.n351 VTAIL.n321 1.16414
R629 VTAIL.n294 VTAIL.n254 1.16414
R630 VTAIL.n289 VTAIL.n259 1.16414
R631 VTAIL.n232 VTAIL.n192 1.16414
R632 VTAIL.n227 VTAIL.n197 1.16414
R633 VTAIL.n309 VTAIL.n247 0.569465
R634 VTAIL.n433 VTAIL.n371 0.569465
R635 VTAIL.n185 VTAIL.n123 0.569465
R636 VTAIL.n371 VTAIL.n309 0.470328
R637 VTAIL.n123 VTAIL.n61 0.470328
R638 VTAIL.n476 VTAIL.n475 0.388379
R639 VTAIL.n479 VTAIL.n442 0.388379
R640 VTAIL.n42 VTAIL.n41 0.388379
R641 VTAIL.n45 VTAIL.n8 0.388379
R642 VTAIL.n104 VTAIL.n103 0.388379
R643 VTAIL.n107 VTAIL.n70 0.388379
R644 VTAIL.n166 VTAIL.n165 0.388379
R645 VTAIL.n169 VTAIL.n132 0.388379
R646 VTAIL.n417 VTAIL.n380 0.388379
R647 VTAIL.n414 VTAIL.n382 0.388379
R648 VTAIL.n355 VTAIL.n318 0.388379
R649 VTAIL.n352 VTAIL.n320 0.388379
R650 VTAIL.n293 VTAIL.n256 0.388379
R651 VTAIL.n290 VTAIL.n258 0.388379
R652 VTAIL.n231 VTAIL.n194 0.388379
R653 VTAIL.n228 VTAIL.n196 0.388379
R654 VTAIL VTAIL.n61 0.343172
R655 VTAIL VTAIL.n495 0.226793
R656 VTAIL.n459 VTAIL.n451 0.155672
R657 VTAIL.n460 VTAIL.n459 0.155672
R658 VTAIL.n460 VTAIL.n447 0.155672
R659 VTAIL.n467 VTAIL.n447 0.155672
R660 VTAIL.n468 VTAIL.n467 0.155672
R661 VTAIL.n468 VTAIL.n443 0.155672
R662 VTAIL.n477 VTAIL.n443 0.155672
R663 VTAIL.n478 VTAIL.n477 0.155672
R664 VTAIL.n478 VTAIL.n439 0.155672
R665 VTAIL.n485 VTAIL.n439 0.155672
R666 VTAIL.n486 VTAIL.n485 0.155672
R667 VTAIL.n486 VTAIL.n435 0.155672
R668 VTAIL.n493 VTAIL.n435 0.155672
R669 VTAIL.n25 VTAIL.n17 0.155672
R670 VTAIL.n26 VTAIL.n25 0.155672
R671 VTAIL.n26 VTAIL.n13 0.155672
R672 VTAIL.n33 VTAIL.n13 0.155672
R673 VTAIL.n34 VTAIL.n33 0.155672
R674 VTAIL.n34 VTAIL.n9 0.155672
R675 VTAIL.n43 VTAIL.n9 0.155672
R676 VTAIL.n44 VTAIL.n43 0.155672
R677 VTAIL.n44 VTAIL.n5 0.155672
R678 VTAIL.n51 VTAIL.n5 0.155672
R679 VTAIL.n52 VTAIL.n51 0.155672
R680 VTAIL.n52 VTAIL.n1 0.155672
R681 VTAIL.n59 VTAIL.n1 0.155672
R682 VTAIL.n87 VTAIL.n79 0.155672
R683 VTAIL.n88 VTAIL.n87 0.155672
R684 VTAIL.n88 VTAIL.n75 0.155672
R685 VTAIL.n95 VTAIL.n75 0.155672
R686 VTAIL.n96 VTAIL.n95 0.155672
R687 VTAIL.n96 VTAIL.n71 0.155672
R688 VTAIL.n105 VTAIL.n71 0.155672
R689 VTAIL.n106 VTAIL.n105 0.155672
R690 VTAIL.n106 VTAIL.n67 0.155672
R691 VTAIL.n113 VTAIL.n67 0.155672
R692 VTAIL.n114 VTAIL.n113 0.155672
R693 VTAIL.n114 VTAIL.n63 0.155672
R694 VTAIL.n121 VTAIL.n63 0.155672
R695 VTAIL.n149 VTAIL.n141 0.155672
R696 VTAIL.n150 VTAIL.n149 0.155672
R697 VTAIL.n150 VTAIL.n137 0.155672
R698 VTAIL.n157 VTAIL.n137 0.155672
R699 VTAIL.n158 VTAIL.n157 0.155672
R700 VTAIL.n158 VTAIL.n133 0.155672
R701 VTAIL.n167 VTAIL.n133 0.155672
R702 VTAIL.n168 VTAIL.n167 0.155672
R703 VTAIL.n168 VTAIL.n129 0.155672
R704 VTAIL.n175 VTAIL.n129 0.155672
R705 VTAIL.n176 VTAIL.n175 0.155672
R706 VTAIL.n176 VTAIL.n125 0.155672
R707 VTAIL.n183 VTAIL.n125 0.155672
R708 VTAIL.n431 VTAIL.n373 0.155672
R709 VTAIL.n424 VTAIL.n373 0.155672
R710 VTAIL.n424 VTAIL.n423 0.155672
R711 VTAIL.n423 VTAIL.n377 0.155672
R712 VTAIL.n416 VTAIL.n377 0.155672
R713 VTAIL.n416 VTAIL.n415 0.155672
R714 VTAIL.n415 VTAIL.n381 0.155672
R715 VTAIL.n408 VTAIL.n381 0.155672
R716 VTAIL.n408 VTAIL.n407 0.155672
R717 VTAIL.n407 VTAIL.n387 0.155672
R718 VTAIL.n400 VTAIL.n387 0.155672
R719 VTAIL.n400 VTAIL.n399 0.155672
R720 VTAIL.n399 VTAIL.n391 0.155672
R721 VTAIL.n369 VTAIL.n311 0.155672
R722 VTAIL.n362 VTAIL.n311 0.155672
R723 VTAIL.n362 VTAIL.n361 0.155672
R724 VTAIL.n361 VTAIL.n315 0.155672
R725 VTAIL.n354 VTAIL.n315 0.155672
R726 VTAIL.n354 VTAIL.n353 0.155672
R727 VTAIL.n353 VTAIL.n319 0.155672
R728 VTAIL.n346 VTAIL.n319 0.155672
R729 VTAIL.n346 VTAIL.n345 0.155672
R730 VTAIL.n345 VTAIL.n325 0.155672
R731 VTAIL.n338 VTAIL.n325 0.155672
R732 VTAIL.n338 VTAIL.n337 0.155672
R733 VTAIL.n337 VTAIL.n329 0.155672
R734 VTAIL.n307 VTAIL.n249 0.155672
R735 VTAIL.n300 VTAIL.n249 0.155672
R736 VTAIL.n300 VTAIL.n299 0.155672
R737 VTAIL.n299 VTAIL.n253 0.155672
R738 VTAIL.n292 VTAIL.n253 0.155672
R739 VTAIL.n292 VTAIL.n291 0.155672
R740 VTAIL.n291 VTAIL.n257 0.155672
R741 VTAIL.n284 VTAIL.n257 0.155672
R742 VTAIL.n284 VTAIL.n283 0.155672
R743 VTAIL.n283 VTAIL.n263 0.155672
R744 VTAIL.n276 VTAIL.n263 0.155672
R745 VTAIL.n276 VTAIL.n275 0.155672
R746 VTAIL.n275 VTAIL.n267 0.155672
R747 VTAIL.n245 VTAIL.n187 0.155672
R748 VTAIL.n238 VTAIL.n187 0.155672
R749 VTAIL.n238 VTAIL.n237 0.155672
R750 VTAIL.n237 VTAIL.n191 0.155672
R751 VTAIL.n230 VTAIL.n191 0.155672
R752 VTAIL.n230 VTAIL.n229 0.155672
R753 VTAIL.n229 VTAIL.n195 0.155672
R754 VTAIL.n222 VTAIL.n195 0.155672
R755 VTAIL.n222 VTAIL.n221 0.155672
R756 VTAIL.n221 VTAIL.n201 0.155672
R757 VTAIL.n214 VTAIL.n201 0.155672
R758 VTAIL.n214 VTAIL.n213 0.155672
R759 VTAIL.n213 VTAIL.n205 0.155672
R760 VDD1 VDD1.n1 99.7041
R761 VDD1 VDD1.n0 63.8934
R762 VDD1.n0 VDD1.t1 1.72374
R763 VDD1.n0 VDD1.t3 1.72374
R764 VDD1.n1 VDD1.t2 1.72374
R765 VDD1.n1 VDD1.t0 1.72374
R766 B.n135 B.t15 1051.73
R767 B.n127 B.t8 1051.73
R768 B.n51 B.t4 1051.73
R769 B.n57 B.t12 1051.73
R770 B.n397 B.n396 585
R771 B.n399 B.n79 585
R772 B.n402 B.n401 585
R773 B.n403 B.n78 585
R774 B.n405 B.n404 585
R775 B.n407 B.n77 585
R776 B.n410 B.n409 585
R777 B.n411 B.n76 585
R778 B.n413 B.n412 585
R779 B.n415 B.n75 585
R780 B.n418 B.n417 585
R781 B.n419 B.n74 585
R782 B.n421 B.n420 585
R783 B.n423 B.n73 585
R784 B.n426 B.n425 585
R785 B.n427 B.n72 585
R786 B.n429 B.n428 585
R787 B.n431 B.n71 585
R788 B.n434 B.n433 585
R789 B.n435 B.n70 585
R790 B.n437 B.n436 585
R791 B.n439 B.n69 585
R792 B.n442 B.n441 585
R793 B.n443 B.n68 585
R794 B.n445 B.n444 585
R795 B.n447 B.n67 585
R796 B.n450 B.n449 585
R797 B.n451 B.n66 585
R798 B.n453 B.n452 585
R799 B.n455 B.n65 585
R800 B.n458 B.n457 585
R801 B.n459 B.n64 585
R802 B.n461 B.n460 585
R803 B.n463 B.n63 585
R804 B.n466 B.n465 585
R805 B.n467 B.n62 585
R806 B.n469 B.n468 585
R807 B.n471 B.n61 585
R808 B.n473 B.n472 585
R809 B.n475 B.n474 585
R810 B.n478 B.n477 585
R811 B.n479 B.n56 585
R812 B.n481 B.n480 585
R813 B.n483 B.n55 585
R814 B.n486 B.n485 585
R815 B.n487 B.n54 585
R816 B.n489 B.n488 585
R817 B.n491 B.n53 585
R818 B.n494 B.n493 585
R819 B.n495 B.n50 585
R820 B.n498 B.n497 585
R821 B.n500 B.n49 585
R822 B.n503 B.n502 585
R823 B.n504 B.n48 585
R824 B.n506 B.n505 585
R825 B.n508 B.n47 585
R826 B.n511 B.n510 585
R827 B.n512 B.n46 585
R828 B.n514 B.n513 585
R829 B.n516 B.n45 585
R830 B.n519 B.n518 585
R831 B.n520 B.n44 585
R832 B.n522 B.n521 585
R833 B.n524 B.n43 585
R834 B.n527 B.n526 585
R835 B.n528 B.n42 585
R836 B.n530 B.n529 585
R837 B.n532 B.n41 585
R838 B.n535 B.n534 585
R839 B.n536 B.n40 585
R840 B.n538 B.n537 585
R841 B.n540 B.n39 585
R842 B.n543 B.n542 585
R843 B.n544 B.n38 585
R844 B.n546 B.n545 585
R845 B.n548 B.n37 585
R846 B.n551 B.n550 585
R847 B.n552 B.n36 585
R848 B.n554 B.n553 585
R849 B.n556 B.n35 585
R850 B.n559 B.n558 585
R851 B.n560 B.n34 585
R852 B.n562 B.n561 585
R853 B.n564 B.n33 585
R854 B.n567 B.n566 585
R855 B.n568 B.n32 585
R856 B.n570 B.n569 585
R857 B.n572 B.n31 585
R858 B.n575 B.n574 585
R859 B.n576 B.n30 585
R860 B.n395 B.n28 585
R861 B.n579 B.n28 585
R862 B.n394 B.n27 585
R863 B.n580 B.n27 585
R864 B.n393 B.n26 585
R865 B.n581 B.n26 585
R866 B.n392 B.n391 585
R867 B.n391 B.n22 585
R868 B.n390 B.n21 585
R869 B.n587 B.n21 585
R870 B.n389 B.n20 585
R871 B.n588 B.n20 585
R872 B.n388 B.n19 585
R873 B.n589 B.n19 585
R874 B.n387 B.n386 585
R875 B.n386 B.n15 585
R876 B.n385 B.n14 585
R877 B.n595 B.n14 585
R878 B.n384 B.n13 585
R879 B.n596 B.n13 585
R880 B.n383 B.n12 585
R881 B.n597 B.n12 585
R882 B.n382 B.n381 585
R883 B.n381 B.n11 585
R884 B.n380 B.n7 585
R885 B.n603 B.n7 585
R886 B.n379 B.n6 585
R887 B.n604 B.n6 585
R888 B.n378 B.n5 585
R889 B.n605 B.n5 585
R890 B.n377 B.n376 585
R891 B.n376 B.n4 585
R892 B.n375 B.n80 585
R893 B.n375 B.n374 585
R894 B.n364 B.n81 585
R895 B.n367 B.n81 585
R896 B.n366 B.n365 585
R897 B.n368 B.n366 585
R898 B.n363 B.n85 585
R899 B.n89 B.n85 585
R900 B.n362 B.n361 585
R901 B.n361 B.n360 585
R902 B.n87 B.n86 585
R903 B.n88 B.n87 585
R904 B.n353 B.n352 585
R905 B.n354 B.n353 585
R906 B.n351 B.n94 585
R907 B.n94 B.n93 585
R908 B.n350 B.n349 585
R909 B.n349 B.n348 585
R910 B.n96 B.n95 585
R911 B.n97 B.n96 585
R912 B.n341 B.n340 585
R913 B.n342 B.n341 585
R914 B.n339 B.n102 585
R915 B.n102 B.n101 585
R916 B.n338 B.n337 585
R917 B.n337 B.n336 585
R918 B.n333 B.n106 585
R919 B.n332 B.n331 585
R920 B.n329 B.n107 585
R921 B.n329 B.n105 585
R922 B.n328 B.n327 585
R923 B.n326 B.n325 585
R924 B.n324 B.n109 585
R925 B.n322 B.n321 585
R926 B.n320 B.n110 585
R927 B.n319 B.n318 585
R928 B.n316 B.n111 585
R929 B.n314 B.n313 585
R930 B.n312 B.n112 585
R931 B.n311 B.n310 585
R932 B.n308 B.n113 585
R933 B.n306 B.n305 585
R934 B.n304 B.n114 585
R935 B.n303 B.n302 585
R936 B.n300 B.n115 585
R937 B.n298 B.n297 585
R938 B.n296 B.n116 585
R939 B.n295 B.n294 585
R940 B.n292 B.n117 585
R941 B.n290 B.n289 585
R942 B.n288 B.n118 585
R943 B.n287 B.n286 585
R944 B.n284 B.n119 585
R945 B.n282 B.n281 585
R946 B.n280 B.n120 585
R947 B.n279 B.n278 585
R948 B.n276 B.n121 585
R949 B.n274 B.n273 585
R950 B.n272 B.n122 585
R951 B.n271 B.n270 585
R952 B.n268 B.n123 585
R953 B.n266 B.n265 585
R954 B.n264 B.n124 585
R955 B.n263 B.n262 585
R956 B.n260 B.n125 585
R957 B.n258 B.n257 585
R958 B.n256 B.n126 585
R959 B.n254 B.n253 585
R960 B.n251 B.n129 585
R961 B.n249 B.n248 585
R962 B.n247 B.n130 585
R963 B.n246 B.n245 585
R964 B.n243 B.n131 585
R965 B.n241 B.n240 585
R966 B.n239 B.n132 585
R967 B.n238 B.n237 585
R968 B.n235 B.n133 585
R969 B.n233 B.n232 585
R970 B.n231 B.n134 585
R971 B.n230 B.n229 585
R972 B.n227 B.n138 585
R973 B.n225 B.n224 585
R974 B.n223 B.n139 585
R975 B.n222 B.n221 585
R976 B.n219 B.n140 585
R977 B.n217 B.n216 585
R978 B.n215 B.n141 585
R979 B.n214 B.n213 585
R980 B.n211 B.n142 585
R981 B.n209 B.n208 585
R982 B.n207 B.n143 585
R983 B.n206 B.n205 585
R984 B.n203 B.n144 585
R985 B.n201 B.n200 585
R986 B.n199 B.n145 585
R987 B.n198 B.n197 585
R988 B.n195 B.n146 585
R989 B.n193 B.n192 585
R990 B.n191 B.n147 585
R991 B.n190 B.n189 585
R992 B.n187 B.n148 585
R993 B.n185 B.n184 585
R994 B.n183 B.n149 585
R995 B.n182 B.n181 585
R996 B.n179 B.n150 585
R997 B.n177 B.n176 585
R998 B.n175 B.n151 585
R999 B.n174 B.n173 585
R1000 B.n171 B.n152 585
R1001 B.n169 B.n168 585
R1002 B.n167 B.n153 585
R1003 B.n166 B.n165 585
R1004 B.n163 B.n154 585
R1005 B.n161 B.n160 585
R1006 B.n159 B.n155 585
R1007 B.n158 B.n157 585
R1008 B.n104 B.n103 585
R1009 B.n105 B.n104 585
R1010 B.n335 B.n334 585
R1011 B.n336 B.n335 585
R1012 B.n100 B.n99 585
R1013 B.n101 B.n100 585
R1014 B.n344 B.n343 585
R1015 B.n343 B.n342 585
R1016 B.n345 B.n98 585
R1017 B.n98 B.n97 585
R1018 B.n347 B.n346 585
R1019 B.n348 B.n347 585
R1020 B.n92 B.n91 585
R1021 B.n93 B.n92 585
R1022 B.n356 B.n355 585
R1023 B.n355 B.n354 585
R1024 B.n357 B.n90 585
R1025 B.n90 B.n88 585
R1026 B.n359 B.n358 585
R1027 B.n360 B.n359 585
R1028 B.n84 B.n83 585
R1029 B.n89 B.n84 585
R1030 B.n370 B.n369 585
R1031 B.n369 B.n368 585
R1032 B.n371 B.n82 585
R1033 B.n367 B.n82 585
R1034 B.n373 B.n372 585
R1035 B.n374 B.n373 585
R1036 B.n2 B.n0 585
R1037 B.n4 B.n2 585
R1038 B.n3 B.n1 585
R1039 B.n604 B.n3 585
R1040 B.n602 B.n601 585
R1041 B.n603 B.n602 585
R1042 B.n600 B.n8 585
R1043 B.n11 B.n8 585
R1044 B.n599 B.n598 585
R1045 B.n598 B.n597 585
R1046 B.n10 B.n9 585
R1047 B.n596 B.n10 585
R1048 B.n594 B.n593 585
R1049 B.n595 B.n594 585
R1050 B.n592 B.n16 585
R1051 B.n16 B.n15 585
R1052 B.n591 B.n590 585
R1053 B.n590 B.n589 585
R1054 B.n18 B.n17 585
R1055 B.n588 B.n18 585
R1056 B.n586 B.n585 585
R1057 B.n587 B.n586 585
R1058 B.n584 B.n23 585
R1059 B.n23 B.n22 585
R1060 B.n583 B.n582 585
R1061 B.n582 B.n581 585
R1062 B.n25 B.n24 585
R1063 B.n580 B.n25 585
R1064 B.n578 B.n577 585
R1065 B.n579 B.n578 585
R1066 B.n607 B.n606 585
R1067 B.n606 B.n605 585
R1068 B.n335 B.n106 482.89
R1069 B.n578 B.n30 482.89
R1070 B.n337 B.n104 482.89
R1071 B.n397 B.n28 482.89
R1072 B.n135 B.t17 286.392
R1073 B.n57 B.t13 286.392
R1074 B.n127 B.t11 286.392
R1075 B.n51 B.t6 286.392
R1076 B.n136 B.t16 273.592
R1077 B.n58 B.t14 273.592
R1078 B.n128 B.t10 273.592
R1079 B.n52 B.t7 273.592
R1080 B.n398 B.n29 256.663
R1081 B.n400 B.n29 256.663
R1082 B.n406 B.n29 256.663
R1083 B.n408 B.n29 256.663
R1084 B.n414 B.n29 256.663
R1085 B.n416 B.n29 256.663
R1086 B.n422 B.n29 256.663
R1087 B.n424 B.n29 256.663
R1088 B.n430 B.n29 256.663
R1089 B.n432 B.n29 256.663
R1090 B.n438 B.n29 256.663
R1091 B.n440 B.n29 256.663
R1092 B.n446 B.n29 256.663
R1093 B.n448 B.n29 256.663
R1094 B.n454 B.n29 256.663
R1095 B.n456 B.n29 256.663
R1096 B.n462 B.n29 256.663
R1097 B.n464 B.n29 256.663
R1098 B.n470 B.n29 256.663
R1099 B.n60 B.n29 256.663
R1100 B.n476 B.n29 256.663
R1101 B.n482 B.n29 256.663
R1102 B.n484 B.n29 256.663
R1103 B.n490 B.n29 256.663
R1104 B.n492 B.n29 256.663
R1105 B.n499 B.n29 256.663
R1106 B.n501 B.n29 256.663
R1107 B.n507 B.n29 256.663
R1108 B.n509 B.n29 256.663
R1109 B.n515 B.n29 256.663
R1110 B.n517 B.n29 256.663
R1111 B.n523 B.n29 256.663
R1112 B.n525 B.n29 256.663
R1113 B.n531 B.n29 256.663
R1114 B.n533 B.n29 256.663
R1115 B.n539 B.n29 256.663
R1116 B.n541 B.n29 256.663
R1117 B.n547 B.n29 256.663
R1118 B.n549 B.n29 256.663
R1119 B.n555 B.n29 256.663
R1120 B.n557 B.n29 256.663
R1121 B.n563 B.n29 256.663
R1122 B.n565 B.n29 256.663
R1123 B.n571 B.n29 256.663
R1124 B.n573 B.n29 256.663
R1125 B.n330 B.n105 256.663
R1126 B.n108 B.n105 256.663
R1127 B.n323 B.n105 256.663
R1128 B.n317 B.n105 256.663
R1129 B.n315 B.n105 256.663
R1130 B.n309 B.n105 256.663
R1131 B.n307 B.n105 256.663
R1132 B.n301 B.n105 256.663
R1133 B.n299 B.n105 256.663
R1134 B.n293 B.n105 256.663
R1135 B.n291 B.n105 256.663
R1136 B.n285 B.n105 256.663
R1137 B.n283 B.n105 256.663
R1138 B.n277 B.n105 256.663
R1139 B.n275 B.n105 256.663
R1140 B.n269 B.n105 256.663
R1141 B.n267 B.n105 256.663
R1142 B.n261 B.n105 256.663
R1143 B.n259 B.n105 256.663
R1144 B.n252 B.n105 256.663
R1145 B.n250 B.n105 256.663
R1146 B.n244 B.n105 256.663
R1147 B.n242 B.n105 256.663
R1148 B.n236 B.n105 256.663
R1149 B.n234 B.n105 256.663
R1150 B.n228 B.n105 256.663
R1151 B.n226 B.n105 256.663
R1152 B.n220 B.n105 256.663
R1153 B.n218 B.n105 256.663
R1154 B.n212 B.n105 256.663
R1155 B.n210 B.n105 256.663
R1156 B.n204 B.n105 256.663
R1157 B.n202 B.n105 256.663
R1158 B.n196 B.n105 256.663
R1159 B.n194 B.n105 256.663
R1160 B.n188 B.n105 256.663
R1161 B.n186 B.n105 256.663
R1162 B.n180 B.n105 256.663
R1163 B.n178 B.n105 256.663
R1164 B.n172 B.n105 256.663
R1165 B.n170 B.n105 256.663
R1166 B.n164 B.n105 256.663
R1167 B.n162 B.n105 256.663
R1168 B.n156 B.n105 256.663
R1169 B.n335 B.n100 163.367
R1170 B.n343 B.n100 163.367
R1171 B.n343 B.n98 163.367
R1172 B.n347 B.n98 163.367
R1173 B.n347 B.n92 163.367
R1174 B.n355 B.n92 163.367
R1175 B.n355 B.n90 163.367
R1176 B.n359 B.n90 163.367
R1177 B.n359 B.n84 163.367
R1178 B.n369 B.n84 163.367
R1179 B.n369 B.n82 163.367
R1180 B.n373 B.n82 163.367
R1181 B.n373 B.n2 163.367
R1182 B.n606 B.n2 163.367
R1183 B.n606 B.n3 163.367
R1184 B.n602 B.n3 163.367
R1185 B.n602 B.n8 163.367
R1186 B.n598 B.n8 163.367
R1187 B.n598 B.n10 163.367
R1188 B.n594 B.n10 163.367
R1189 B.n594 B.n16 163.367
R1190 B.n590 B.n16 163.367
R1191 B.n590 B.n18 163.367
R1192 B.n586 B.n18 163.367
R1193 B.n586 B.n23 163.367
R1194 B.n582 B.n23 163.367
R1195 B.n582 B.n25 163.367
R1196 B.n578 B.n25 163.367
R1197 B.n331 B.n329 163.367
R1198 B.n329 B.n328 163.367
R1199 B.n325 B.n324 163.367
R1200 B.n322 B.n110 163.367
R1201 B.n318 B.n316 163.367
R1202 B.n314 B.n112 163.367
R1203 B.n310 B.n308 163.367
R1204 B.n306 B.n114 163.367
R1205 B.n302 B.n300 163.367
R1206 B.n298 B.n116 163.367
R1207 B.n294 B.n292 163.367
R1208 B.n290 B.n118 163.367
R1209 B.n286 B.n284 163.367
R1210 B.n282 B.n120 163.367
R1211 B.n278 B.n276 163.367
R1212 B.n274 B.n122 163.367
R1213 B.n270 B.n268 163.367
R1214 B.n266 B.n124 163.367
R1215 B.n262 B.n260 163.367
R1216 B.n258 B.n126 163.367
R1217 B.n253 B.n251 163.367
R1218 B.n249 B.n130 163.367
R1219 B.n245 B.n243 163.367
R1220 B.n241 B.n132 163.367
R1221 B.n237 B.n235 163.367
R1222 B.n233 B.n134 163.367
R1223 B.n229 B.n227 163.367
R1224 B.n225 B.n139 163.367
R1225 B.n221 B.n219 163.367
R1226 B.n217 B.n141 163.367
R1227 B.n213 B.n211 163.367
R1228 B.n209 B.n143 163.367
R1229 B.n205 B.n203 163.367
R1230 B.n201 B.n145 163.367
R1231 B.n197 B.n195 163.367
R1232 B.n193 B.n147 163.367
R1233 B.n189 B.n187 163.367
R1234 B.n185 B.n149 163.367
R1235 B.n181 B.n179 163.367
R1236 B.n177 B.n151 163.367
R1237 B.n173 B.n171 163.367
R1238 B.n169 B.n153 163.367
R1239 B.n165 B.n163 163.367
R1240 B.n161 B.n155 163.367
R1241 B.n157 B.n104 163.367
R1242 B.n337 B.n102 163.367
R1243 B.n341 B.n102 163.367
R1244 B.n341 B.n96 163.367
R1245 B.n349 B.n96 163.367
R1246 B.n349 B.n94 163.367
R1247 B.n353 B.n94 163.367
R1248 B.n353 B.n87 163.367
R1249 B.n361 B.n87 163.367
R1250 B.n361 B.n85 163.367
R1251 B.n366 B.n85 163.367
R1252 B.n366 B.n81 163.367
R1253 B.n375 B.n81 163.367
R1254 B.n376 B.n375 163.367
R1255 B.n376 B.n5 163.367
R1256 B.n6 B.n5 163.367
R1257 B.n7 B.n6 163.367
R1258 B.n381 B.n7 163.367
R1259 B.n381 B.n12 163.367
R1260 B.n13 B.n12 163.367
R1261 B.n14 B.n13 163.367
R1262 B.n386 B.n14 163.367
R1263 B.n386 B.n19 163.367
R1264 B.n20 B.n19 163.367
R1265 B.n21 B.n20 163.367
R1266 B.n391 B.n21 163.367
R1267 B.n391 B.n26 163.367
R1268 B.n27 B.n26 163.367
R1269 B.n28 B.n27 163.367
R1270 B.n574 B.n572 163.367
R1271 B.n570 B.n32 163.367
R1272 B.n566 B.n564 163.367
R1273 B.n562 B.n34 163.367
R1274 B.n558 B.n556 163.367
R1275 B.n554 B.n36 163.367
R1276 B.n550 B.n548 163.367
R1277 B.n546 B.n38 163.367
R1278 B.n542 B.n540 163.367
R1279 B.n538 B.n40 163.367
R1280 B.n534 B.n532 163.367
R1281 B.n530 B.n42 163.367
R1282 B.n526 B.n524 163.367
R1283 B.n522 B.n44 163.367
R1284 B.n518 B.n516 163.367
R1285 B.n514 B.n46 163.367
R1286 B.n510 B.n508 163.367
R1287 B.n506 B.n48 163.367
R1288 B.n502 B.n500 163.367
R1289 B.n498 B.n50 163.367
R1290 B.n493 B.n491 163.367
R1291 B.n489 B.n54 163.367
R1292 B.n485 B.n483 163.367
R1293 B.n481 B.n56 163.367
R1294 B.n477 B.n475 163.367
R1295 B.n472 B.n471 163.367
R1296 B.n469 B.n62 163.367
R1297 B.n465 B.n463 163.367
R1298 B.n461 B.n64 163.367
R1299 B.n457 B.n455 163.367
R1300 B.n453 B.n66 163.367
R1301 B.n449 B.n447 163.367
R1302 B.n445 B.n68 163.367
R1303 B.n441 B.n439 163.367
R1304 B.n437 B.n70 163.367
R1305 B.n433 B.n431 163.367
R1306 B.n429 B.n72 163.367
R1307 B.n425 B.n423 163.367
R1308 B.n421 B.n74 163.367
R1309 B.n417 B.n415 163.367
R1310 B.n413 B.n76 163.367
R1311 B.n409 B.n407 163.367
R1312 B.n405 B.n78 163.367
R1313 B.n401 B.n399 163.367
R1314 B.n336 B.n105 77.9868
R1315 B.n579 B.n29 77.9868
R1316 B.n330 B.n106 71.676
R1317 B.n328 B.n108 71.676
R1318 B.n324 B.n323 71.676
R1319 B.n317 B.n110 71.676
R1320 B.n316 B.n315 71.676
R1321 B.n309 B.n112 71.676
R1322 B.n308 B.n307 71.676
R1323 B.n301 B.n114 71.676
R1324 B.n300 B.n299 71.676
R1325 B.n293 B.n116 71.676
R1326 B.n292 B.n291 71.676
R1327 B.n285 B.n118 71.676
R1328 B.n284 B.n283 71.676
R1329 B.n277 B.n120 71.676
R1330 B.n276 B.n275 71.676
R1331 B.n269 B.n122 71.676
R1332 B.n268 B.n267 71.676
R1333 B.n261 B.n124 71.676
R1334 B.n260 B.n259 71.676
R1335 B.n252 B.n126 71.676
R1336 B.n251 B.n250 71.676
R1337 B.n244 B.n130 71.676
R1338 B.n243 B.n242 71.676
R1339 B.n236 B.n132 71.676
R1340 B.n235 B.n234 71.676
R1341 B.n228 B.n134 71.676
R1342 B.n227 B.n226 71.676
R1343 B.n220 B.n139 71.676
R1344 B.n219 B.n218 71.676
R1345 B.n212 B.n141 71.676
R1346 B.n211 B.n210 71.676
R1347 B.n204 B.n143 71.676
R1348 B.n203 B.n202 71.676
R1349 B.n196 B.n145 71.676
R1350 B.n195 B.n194 71.676
R1351 B.n188 B.n147 71.676
R1352 B.n187 B.n186 71.676
R1353 B.n180 B.n149 71.676
R1354 B.n179 B.n178 71.676
R1355 B.n172 B.n151 71.676
R1356 B.n171 B.n170 71.676
R1357 B.n164 B.n153 71.676
R1358 B.n163 B.n162 71.676
R1359 B.n156 B.n155 71.676
R1360 B.n573 B.n30 71.676
R1361 B.n572 B.n571 71.676
R1362 B.n565 B.n32 71.676
R1363 B.n564 B.n563 71.676
R1364 B.n557 B.n34 71.676
R1365 B.n556 B.n555 71.676
R1366 B.n549 B.n36 71.676
R1367 B.n548 B.n547 71.676
R1368 B.n541 B.n38 71.676
R1369 B.n540 B.n539 71.676
R1370 B.n533 B.n40 71.676
R1371 B.n532 B.n531 71.676
R1372 B.n525 B.n42 71.676
R1373 B.n524 B.n523 71.676
R1374 B.n517 B.n44 71.676
R1375 B.n516 B.n515 71.676
R1376 B.n509 B.n46 71.676
R1377 B.n508 B.n507 71.676
R1378 B.n501 B.n48 71.676
R1379 B.n500 B.n499 71.676
R1380 B.n492 B.n50 71.676
R1381 B.n491 B.n490 71.676
R1382 B.n484 B.n54 71.676
R1383 B.n483 B.n482 71.676
R1384 B.n476 B.n56 71.676
R1385 B.n475 B.n60 71.676
R1386 B.n471 B.n470 71.676
R1387 B.n464 B.n62 71.676
R1388 B.n463 B.n462 71.676
R1389 B.n456 B.n64 71.676
R1390 B.n455 B.n454 71.676
R1391 B.n448 B.n66 71.676
R1392 B.n447 B.n446 71.676
R1393 B.n440 B.n68 71.676
R1394 B.n439 B.n438 71.676
R1395 B.n432 B.n70 71.676
R1396 B.n431 B.n430 71.676
R1397 B.n424 B.n72 71.676
R1398 B.n423 B.n422 71.676
R1399 B.n416 B.n74 71.676
R1400 B.n415 B.n414 71.676
R1401 B.n408 B.n76 71.676
R1402 B.n407 B.n406 71.676
R1403 B.n400 B.n78 71.676
R1404 B.n399 B.n398 71.676
R1405 B.n398 B.n397 71.676
R1406 B.n401 B.n400 71.676
R1407 B.n406 B.n405 71.676
R1408 B.n409 B.n408 71.676
R1409 B.n414 B.n413 71.676
R1410 B.n417 B.n416 71.676
R1411 B.n422 B.n421 71.676
R1412 B.n425 B.n424 71.676
R1413 B.n430 B.n429 71.676
R1414 B.n433 B.n432 71.676
R1415 B.n438 B.n437 71.676
R1416 B.n441 B.n440 71.676
R1417 B.n446 B.n445 71.676
R1418 B.n449 B.n448 71.676
R1419 B.n454 B.n453 71.676
R1420 B.n457 B.n456 71.676
R1421 B.n462 B.n461 71.676
R1422 B.n465 B.n464 71.676
R1423 B.n470 B.n469 71.676
R1424 B.n472 B.n60 71.676
R1425 B.n477 B.n476 71.676
R1426 B.n482 B.n481 71.676
R1427 B.n485 B.n484 71.676
R1428 B.n490 B.n489 71.676
R1429 B.n493 B.n492 71.676
R1430 B.n499 B.n498 71.676
R1431 B.n502 B.n501 71.676
R1432 B.n507 B.n506 71.676
R1433 B.n510 B.n509 71.676
R1434 B.n515 B.n514 71.676
R1435 B.n518 B.n517 71.676
R1436 B.n523 B.n522 71.676
R1437 B.n526 B.n525 71.676
R1438 B.n531 B.n530 71.676
R1439 B.n534 B.n533 71.676
R1440 B.n539 B.n538 71.676
R1441 B.n542 B.n541 71.676
R1442 B.n547 B.n546 71.676
R1443 B.n550 B.n549 71.676
R1444 B.n555 B.n554 71.676
R1445 B.n558 B.n557 71.676
R1446 B.n563 B.n562 71.676
R1447 B.n566 B.n565 71.676
R1448 B.n571 B.n570 71.676
R1449 B.n574 B.n573 71.676
R1450 B.n331 B.n330 71.676
R1451 B.n325 B.n108 71.676
R1452 B.n323 B.n322 71.676
R1453 B.n318 B.n317 71.676
R1454 B.n315 B.n314 71.676
R1455 B.n310 B.n309 71.676
R1456 B.n307 B.n306 71.676
R1457 B.n302 B.n301 71.676
R1458 B.n299 B.n298 71.676
R1459 B.n294 B.n293 71.676
R1460 B.n291 B.n290 71.676
R1461 B.n286 B.n285 71.676
R1462 B.n283 B.n282 71.676
R1463 B.n278 B.n277 71.676
R1464 B.n275 B.n274 71.676
R1465 B.n270 B.n269 71.676
R1466 B.n267 B.n266 71.676
R1467 B.n262 B.n261 71.676
R1468 B.n259 B.n258 71.676
R1469 B.n253 B.n252 71.676
R1470 B.n250 B.n249 71.676
R1471 B.n245 B.n244 71.676
R1472 B.n242 B.n241 71.676
R1473 B.n237 B.n236 71.676
R1474 B.n234 B.n233 71.676
R1475 B.n229 B.n228 71.676
R1476 B.n226 B.n225 71.676
R1477 B.n221 B.n220 71.676
R1478 B.n218 B.n217 71.676
R1479 B.n213 B.n212 71.676
R1480 B.n210 B.n209 71.676
R1481 B.n205 B.n204 71.676
R1482 B.n202 B.n201 71.676
R1483 B.n197 B.n196 71.676
R1484 B.n194 B.n193 71.676
R1485 B.n189 B.n188 71.676
R1486 B.n186 B.n185 71.676
R1487 B.n181 B.n180 71.676
R1488 B.n178 B.n177 71.676
R1489 B.n173 B.n172 71.676
R1490 B.n170 B.n169 71.676
R1491 B.n165 B.n164 71.676
R1492 B.n162 B.n161 71.676
R1493 B.n157 B.n156 71.676
R1494 B.n137 B.n136 59.5399
R1495 B.n255 B.n128 59.5399
R1496 B.n496 B.n52 59.5399
R1497 B.n59 B.n58 59.5399
R1498 B.n336 B.n101 44.5641
R1499 B.n342 B.n101 44.5641
R1500 B.n342 B.n97 44.5641
R1501 B.n348 B.n97 44.5641
R1502 B.n354 B.n93 44.5641
R1503 B.n354 B.n88 44.5641
R1504 B.n360 B.n88 44.5641
R1505 B.n360 B.n89 44.5641
R1506 B.n368 B.n367 44.5641
R1507 B.n374 B.n4 44.5641
R1508 B.n605 B.n4 44.5641
R1509 B.n605 B.n604 44.5641
R1510 B.n604 B.n603 44.5641
R1511 B.n597 B.n11 44.5641
R1512 B.n596 B.n595 44.5641
R1513 B.n595 B.n15 44.5641
R1514 B.n589 B.n15 44.5641
R1515 B.n589 B.n588 44.5641
R1516 B.n587 B.n22 44.5641
R1517 B.n581 B.n22 44.5641
R1518 B.n581 B.n580 44.5641
R1519 B.n580 B.n579 44.5641
R1520 B.n577 B.n576 31.3761
R1521 B.n396 B.n395 31.3761
R1522 B.n338 B.n103 31.3761
R1523 B.n334 B.n333 31.3761
R1524 B.t9 B.n93 29.4911
R1525 B.n588 B.t5 29.4911
R1526 B.n374 B.t2 25.559
R1527 B.n603 B.t3 25.559
R1528 B.n368 B.t0 22.9376
R1529 B.n597 B.t1 22.9376
R1530 B.n89 B.t0 21.627
R1531 B.t1 B.n596 21.627
R1532 B.n367 B.t2 19.0056
R1533 B.n11 B.t3 19.0056
R1534 B B.n607 18.0485
R1535 B.n348 B.t9 15.0735
R1536 B.t5 B.n587 15.0735
R1537 B.n136 B.n135 12.8005
R1538 B.n128 B.n127 12.8005
R1539 B.n52 B.n51 12.8005
R1540 B.n58 B.n57 12.8005
R1541 B.n576 B.n575 10.6151
R1542 B.n575 B.n31 10.6151
R1543 B.n569 B.n31 10.6151
R1544 B.n569 B.n568 10.6151
R1545 B.n568 B.n567 10.6151
R1546 B.n567 B.n33 10.6151
R1547 B.n561 B.n33 10.6151
R1548 B.n561 B.n560 10.6151
R1549 B.n560 B.n559 10.6151
R1550 B.n559 B.n35 10.6151
R1551 B.n553 B.n35 10.6151
R1552 B.n553 B.n552 10.6151
R1553 B.n552 B.n551 10.6151
R1554 B.n551 B.n37 10.6151
R1555 B.n545 B.n37 10.6151
R1556 B.n545 B.n544 10.6151
R1557 B.n544 B.n543 10.6151
R1558 B.n543 B.n39 10.6151
R1559 B.n537 B.n39 10.6151
R1560 B.n537 B.n536 10.6151
R1561 B.n536 B.n535 10.6151
R1562 B.n535 B.n41 10.6151
R1563 B.n529 B.n41 10.6151
R1564 B.n529 B.n528 10.6151
R1565 B.n528 B.n527 10.6151
R1566 B.n527 B.n43 10.6151
R1567 B.n521 B.n43 10.6151
R1568 B.n521 B.n520 10.6151
R1569 B.n520 B.n519 10.6151
R1570 B.n519 B.n45 10.6151
R1571 B.n513 B.n45 10.6151
R1572 B.n513 B.n512 10.6151
R1573 B.n512 B.n511 10.6151
R1574 B.n511 B.n47 10.6151
R1575 B.n505 B.n47 10.6151
R1576 B.n505 B.n504 10.6151
R1577 B.n504 B.n503 10.6151
R1578 B.n503 B.n49 10.6151
R1579 B.n497 B.n49 10.6151
R1580 B.n495 B.n494 10.6151
R1581 B.n494 B.n53 10.6151
R1582 B.n488 B.n53 10.6151
R1583 B.n488 B.n487 10.6151
R1584 B.n487 B.n486 10.6151
R1585 B.n486 B.n55 10.6151
R1586 B.n480 B.n55 10.6151
R1587 B.n480 B.n479 10.6151
R1588 B.n479 B.n478 10.6151
R1589 B.n474 B.n473 10.6151
R1590 B.n473 B.n61 10.6151
R1591 B.n468 B.n61 10.6151
R1592 B.n468 B.n467 10.6151
R1593 B.n467 B.n466 10.6151
R1594 B.n466 B.n63 10.6151
R1595 B.n460 B.n63 10.6151
R1596 B.n460 B.n459 10.6151
R1597 B.n459 B.n458 10.6151
R1598 B.n458 B.n65 10.6151
R1599 B.n452 B.n65 10.6151
R1600 B.n452 B.n451 10.6151
R1601 B.n451 B.n450 10.6151
R1602 B.n450 B.n67 10.6151
R1603 B.n444 B.n67 10.6151
R1604 B.n444 B.n443 10.6151
R1605 B.n443 B.n442 10.6151
R1606 B.n442 B.n69 10.6151
R1607 B.n436 B.n69 10.6151
R1608 B.n436 B.n435 10.6151
R1609 B.n435 B.n434 10.6151
R1610 B.n434 B.n71 10.6151
R1611 B.n428 B.n71 10.6151
R1612 B.n428 B.n427 10.6151
R1613 B.n427 B.n426 10.6151
R1614 B.n426 B.n73 10.6151
R1615 B.n420 B.n73 10.6151
R1616 B.n420 B.n419 10.6151
R1617 B.n419 B.n418 10.6151
R1618 B.n418 B.n75 10.6151
R1619 B.n412 B.n75 10.6151
R1620 B.n412 B.n411 10.6151
R1621 B.n411 B.n410 10.6151
R1622 B.n410 B.n77 10.6151
R1623 B.n404 B.n77 10.6151
R1624 B.n404 B.n403 10.6151
R1625 B.n403 B.n402 10.6151
R1626 B.n402 B.n79 10.6151
R1627 B.n396 B.n79 10.6151
R1628 B.n339 B.n338 10.6151
R1629 B.n340 B.n339 10.6151
R1630 B.n340 B.n95 10.6151
R1631 B.n350 B.n95 10.6151
R1632 B.n351 B.n350 10.6151
R1633 B.n352 B.n351 10.6151
R1634 B.n352 B.n86 10.6151
R1635 B.n362 B.n86 10.6151
R1636 B.n363 B.n362 10.6151
R1637 B.n365 B.n363 10.6151
R1638 B.n365 B.n364 10.6151
R1639 B.n364 B.n80 10.6151
R1640 B.n377 B.n80 10.6151
R1641 B.n378 B.n377 10.6151
R1642 B.n379 B.n378 10.6151
R1643 B.n380 B.n379 10.6151
R1644 B.n382 B.n380 10.6151
R1645 B.n383 B.n382 10.6151
R1646 B.n384 B.n383 10.6151
R1647 B.n385 B.n384 10.6151
R1648 B.n387 B.n385 10.6151
R1649 B.n388 B.n387 10.6151
R1650 B.n389 B.n388 10.6151
R1651 B.n390 B.n389 10.6151
R1652 B.n392 B.n390 10.6151
R1653 B.n393 B.n392 10.6151
R1654 B.n394 B.n393 10.6151
R1655 B.n395 B.n394 10.6151
R1656 B.n333 B.n332 10.6151
R1657 B.n332 B.n107 10.6151
R1658 B.n327 B.n107 10.6151
R1659 B.n327 B.n326 10.6151
R1660 B.n326 B.n109 10.6151
R1661 B.n321 B.n109 10.6151
R1662 B.n321 B.n320 10.6151
R1663 B.n320 B.n319 10.6151
R1664 B.n319 B.n111 10.6151
R1665 B.n313 B.n111 10.6151
R1666 B.n313 B.n312 10.6151
R1667 B.n312 B.n311 10.6151
R1668 B.n311 B.n113 10.6151
R1669 B.n305 B.n113 10.6151
R1670 B.n305 B.n304 10.6151
R1671 B.n304 B.n303 10.6151
R1672 B.n303 B.n115 10.6151
R1673 B.n297 B.n115 10.6151
R1674 B.n297 B.n296 10.6151
R1675 B.n296 B.n295 10.6151
R1676 B.n295 B.n117 10.6151
R1677 B.n289 B.n117 10.6151
R1678 B.n289 B.n288 10.6151
R1679 B.n288 B.n287 10.6151
R1680 B.n287 B.n119 10.6151
R1681 B.n281 B.n119 10.6151
R1682 B.n281 B.n280 10.6151
R1683 B.n280 B.n279 10.6151
R1684 B.n279 B.n121 10.6151
R1685 B.n273 B.n121 10.6151
R1686 B.n273 B.n272 10.6151
R1687 B.n272 B.n271 10.6151
R1688 B.n271 B.n123 10.6151
R1689 B.n265 B.n123 10.6151
R1690 B.n265 B.n264 10.6151
R1691 B.n264 B.n263 10.6151
R1692 B.n263 B.n125 10.6151
R1693 B.n257 B.n125 10.6151
R1694 B.n257 B.n256 10.6151
R1695 B.n254 B.n129 10.6151
R1696 B.n248 B.n129 10.6151
R1697 B.n248 B.n247 10.6151
R1698 B.n247 B.n246 10.6151
R1699 B.n246 B.n131 10.6151
R1700 B.n240 B.n131 10.6151
R1701 B.n240 B.n239 10.6151
R1702 B.n239 B.n238 10.6151
R1703 B.n238 B.n133 10.6151
R1704 B.n232 B.n231 10.6151
R1705 B.n231 B.n230 10.6151
R1706 B.n230 B.n138 10.6151
R1707 B.n224 B.n138 10.6151
R1708 B.n224 B.n223 10.6151
R1709 B.n223 B.n222 10.6151
R1710 B.n222 B.n140 10.6151
R1711 B.n216 B.n140 10.6151
R1712 B.n216 B.n215 10.6151
R1713 B.n215 B.n214 10.6151
R1714 B.n214 B.n142 10.6151
R1715 B.n208 B.n142 10.6151
R1716 B.n208 B.n207 10.6151
R1717 B.n207 B.n206 10.6151
R1718 B.n206 B.n144 10.6151
R1719 B.n200 B.n144 10.6151
R1720 B.n200 B.n199 10.6151
R1721 B.n199 B.n198 10.6151
R1722 B.n198 B.n146 10.6151
R1723 B.n192 B.n146 10.6151
R1724 B.n192 B.n191 10.6151
R1725 B.n191 B.n190 10.6151
R1726 B.n190 B.n148 10.6151
R1727 B.n184 B.n148 10.6151
R1728 B.n184 B.n183 10.6151
R1729 B.n183 B.n182 10.6151
R1730 B.n182 B.n150 10.6151
R1731 B.n176 B.n150 10.6151
R1732 B.n176 B.n175 10.6151
R1733 B.n175 B.n174 10.6151
R1734 B.n174 B.n152 10.6151
R1735 B.n168 B.n152 10.6151
R1736 B.n168 B.n167 10.6151
R1737 B.n167 B.n166 10.6151
R1738 B.n166 B.n154 10.6151
R1739 B.n160 B.n154 10.6151
R1740 B.n160 B.n159 10.6151
R1741 B.n159 B.n158 10.6151
R1742 B.n158 B.n103 10.6151
R1743 B.n334 B.n99 10.6151
R1744 B.n344 B.n99 10.6151
R1745 B.n345 B.n344 10.6151
R1746 B.n346 B.n345 10.6151
R1747 B.n346 B.n91 10.6151
R1748 B.n356 B.n91 10.6151
R1749 B.n357 B.n356 10.6151
R1750 B.n358 B.n357 10.6151
R1751 B.n358 B.n83 10.6151
R1752 B.n370 B.n83 10.6151
R1753 B.n371 B.n370 10.6151
R1754 B.n372 B.n371 10.6151
R1755 B.n372 B.n0 10.6151
R1756 B.n601 B.n1 10.6151
R1757 B.n601 B.n600 10.6151
R1758 B.n600 B.n599 10.6151
R1759 B.n599 B.n9 10.6151
R1760 B.n593 B.n9 10.6151
R1761 B.n593 B.n592 10.6151
R1762 B.n592 B.n591 10.6151
R1763 B.n591 B.n17 10.6151
R1764 B.n585 B.n17 10.6151
R1765 B.n585 B.n584 10.6151
R1766 B.n584 B.n583 10.6151
R1767 B.n583 B.n24 10.6151
R1768 B.n577 B.n24 10.6151
R1769 B.n497 B.n496 8.74196
R1770 B.n474 B.n59 8.74196
R1771 B.n256 B.n255 8.74196
R1772 B.n232 B.n137 8.74196
R1773 B.n607 B.n0 2.81026
R1774 B.n607 B.n1 2.81026
R1775 B.n496 B.n495 1.87367
R1776 B.n478 B.n59 1.87367
R1777 B.n255 B.n254 1.87367
R1778 B.n137 B.n133 1.87367
R1779 VN.n0 VN.t3 982.989
R1780 VN.n0 VN.t1 982.989
R1781 VN.n1 VN.t2 982.989
R1782 VN.n1 VN.t0 982.989
R1783 VN VN.n1 200.696
R1784 VN VN.n0 161.351
R1785 VDD2.n2 VDD2.n0 99.1793
R1786 VDD2.n2 VDD2.n1 63.8352
R1787 VDD2.n1 VDD2.t1 1.72374
R1788 VDD2.n1 VDD2.t3 1.72374
R1789 VDD2.n0 VDD2.t2 1.72374
R1790 VDD2.n0 VDD2.t0 1.72374
R1791 VDD2 VDD2.n2 0.0586897
C0 VN VDD2 2.10143f
C1 VDD1 VDD2 0.484781f
C2 VP VTAIL 1.62298f
C3 VN VP 4.45418f
C4 VDD1 VP 2.20418f
C5 VN VTAIL 1.60887f
C6 VDD1 VTAIL 8.75684f
C7 VP VDD2 0.251002f
C8 VDD1 VN 0.148089f
C9 VDD2 VTAIL 8.79583f
C10 VDD2 B 2.453267f
C11 VDD1 B 6.46572f
C12 VTAIL B 8.243614f
C13 VN B 7.44429f
C14 VP B 4.076684f
C15 VDD2.t2 B 0.293706f
C16 VDD2.t0 B 0.293706f
C17 VDD2.n0 B 3.25293f
C18 VDD2.t1 B 0.293706f
C19 VDD2.t3 B 0.293706f
C20 VDD2.n1 B 2.61216f
C21 VDD2.n2 B 3.79382f
C22 VN.t1 B 0.527328f
C23 VN.t3 B 0.527328f
C24 VN.n0 B 0.419998f
C25 VN.t2 B 0.527328f
C26 VN.t0 B 0.527328f
C27 VN.n1 B 0.773473f
C28 VDD1.t1 B 0.293187f
C29 VDD1.t3 B 0.293187f
C30 VDD1.n0 B 2.60785f
C31 VDD1.t2 B 0.293187f
C32 VDD1.t0 B 0.293187f
C33 VDD1.n1 B 3.27695f
C34 VTAIL.n0 B 0.022842f
C35 VTAIL.n1 B 0.01587f
C36 VTAIL.n2 B 0.008528f
C37 VTAIL.n3 B 0.020156f
C38 VTAIL.n4 B 0.009029f
C39 VTAIL.n5 B 0.01587f
C40 VTAIL.n6 B 0.008528f
C41 VTAIL.n7 B 0.020156f
C42 VTAIL.n8 B 0.008779f
C43 VTAIL.n9 B 0.01587f
C44 VTAIL.n10 B 0.009029f
C45 VTAIL.n11 B 0.020156f
C46 VTAIL.n12 B 0.009029f
C47 VTAIL.n13 B 0.01587f
C48 VTAIL.n14 B 0.008528f
C49 VTAIL.n15 B 0.020156f
C50 VTAIL.n16 B 0.009029f
C51 VTAIL.n17 B 0.764602f
C52 VTAIL.n18 B 0.008528f
C53 VTAIL.t3 B 0.034f
C54 VTAIL.n19 B 0.111312f
C55 VTAIL.n20 B 0.014249f
C56 VTAIL.n21 B 0.015117f
C57 VTAIL.n22 B 0.020156f
C58 VTAIL.n23 B 0.009029f
C59 VTAIL.n24 B 0.008528f
C60 VTAIL.n25 B 0.01587f
C61 VTAIL.n26 B 0.01587f
C62 VTAIL.n27 B 0.008528f
C63 VTAIL.n28 B 0.009029f
C64 VTAIL.n29 B 0.020156f
C65 VTAIL.n30 B 0.020156f
C66 VTAIL.n31 B 0.009029f
C67 VTAIL.n32 B 0.008528f
C68 VTAIL.n33 B 0.01587f
C69 VTAIL.n34 B 0.01587f
C70 VTAIL.n35 B 0.008528f
C71 VTAIL.n36 B 0.008528f
C72 VTAIL.n37 B 0.009029f
C73 VTAIL.n38 B 0.020156f
C74 VTAIL.n39 B 0.020156f
C75 VTAIL.n40 B 0.020156f
C76 VTAIL.n41 B 0.008779f
C77 VTAIL.n42 B 0.008528f
C78 VTAIL.n43 B 0.01587f
C79 VTAIL.n44 B 0.01587f
C80 VTAIL.n45 B 0.008528f
C81 VTAIL.n46 B 0.009029f
C82 VTAIL.n47 B 0.020156f
C83 VTAIL.n48 B 0.020156f
C84 VTAIL.n49 B 0.009029f
C85 VTAIL.n50 B 0.008528f
C86 VTAIL.n51 B 0.01587f
C87 VTAIL.n52 B 0.01587f
C88 VTAIL.n53 B 0.008528f
C89 VTAIL.n54 B 0.009029f
C90 VTAIL.n55 B 0.020156f
C91 VTAIL.n56 B 0.044582f
C92 VTAIL.n57 B 0.009029f
C93 VTAIL.n58 B 0.008528f
C94 VTAIL.n59 B 0.038633f
C95 VTAIL.n60 B 0.025101f
C96 VTAIL.n61 B 0.056205f
C97 VTAIL.n62 B 0.022842f
C98 VTAIL.n63 B 0.01587f
C99 VTAIL.n64 B 0.008528f
C100 VTAIL.n65 B 0.020156f
C101 VTAIL.n66 B 0.009029f
C102 VTAIL.n67 B 0.01587f
C103 VTAIL.n68 B 0.008528f
C104 VTAIL.n69 B 0.020156f
C105 VTAIL.n70 B 0.008779f
C106 VTAIL.n71 B 0.01587f
C107 VTAIL.n72 B 0.009029f
C108 VTAIL.n73 B 0.020156f
C109 VTAIL.n74 B 0.009029f
C110 VTAIL.n75 B 0.01587f
C111 VTAIL.n76 B 0.008528f
C112 VTAIL.n77 B 0.020156f
C113 VTAIL.n78 B 0.009029f
C114 VTAIL.n79 B 0.764602f
C115 VTAIL.n80 B 0.008528f
C116 VTAIL.t5 B 0.034f
C117 VTAIL.n81 B 0.111312f
C118 VTAIL.n82 B 0.014249f
C119 VTAIL.n83 B 0.015117f
C120 VTAIL.n84 B 0.020156f
C121 VTAIL.n85 B 0.009029f
C122 VTAIL.n86 B 0.008528f
C123 VTAIL.n87 B 0.01587f
C124 VTAIL.n88 B 0.01587f
C125 VTAIL.n89 B 0.008528f
C126 VTAIL.n90 B 0.009029f
C127 VTAIL.n91 B 0.020156f
C128 VTAIL.n92 B 0.020156f
C129 VTAIL.n93 B 0.009029f
C130 VTAIL.n94 B 0.008528f
C131 VTAIL.n95 B 0.01587f
C132 VTAIL.n96 B 0.01587f
C133 VTAIL.n97 B 0.008528f
C134 VTAIL.n98 B 0.008528f
C135 VTAIL.n99 B 0.009029f
C136 VTAIL.n100 B 0.020156f
C137 VTAIL.n101 B 0.020156f
C138 VTAIL.n102 B 0.020156f
C139 VTAIL.n103 B 0.008779f
C140 VTAIL.n104 B 0.008528f
C141 VTAIL.n105 B 0.01587f
C142 VTAIL.n106 B 0.01587f
C143 VTAIL.n107 B 0.008528f
C144 VTAIL.n108 B 0.009029f
C145 VTAIL.n109 B 0.020156f
C146 VTAIL.n110 B 0.020156f
C147 VTAIL.n111 B 0.009029f
C148 VTAIL.n112 B 0.008528f
C149 VTAIL.n113 B 0.01587f
C150 VTAIL.n114 B 0.01587f
C151 VTAIL.n115 B 0.008528f
C152 VTAIL.n116 B 0.009029f
C153 VTAIL.n117 B 0.020156f
C154 VTAIL.n118 B 0.044582f
C155 VTAIL.n119 B 0.009029f
C156 VTAIL.n120 B 0.008528f
C157 VTAIL.n121 B 0.038633f
C158 VTAIL.n122 B 0.025101f
C159 VTAIL.n123 B 0.067776f
C160 VTAIL.n124 B 0.022842f
C161 VTAIL.n125 B 0.01587f
C162 VTAIL.n126 B 0.008528f
C163 VTAIL.n127 B 0.020156f
C164 VTAIL.n128 B 0.009029f
C165 VTAIL.n129 B 0.01587f
C166 VTAIL.n130 B 0.008528f
C167 VTAIL.n131 B 0.020156f
C168 VTAIL.n132 B 0.008779f
C169 VTAIL.n133 B 0.01587f
C170 VTAIL.n134 B 0.009029f
C171 VTAIL.n135 B 0.020156f
C172 VTAIL.n136 B 0.009029f
C173 VTAIL.n137 B 0.01587f
C174 VTAIL.n138 B 0.008528f
C175 VTAIL.n139 B 0.020156f
C176 VTAIL.n140 B 0.009029f
C177 VTAIL.n141 B 0.764602f
C178 VTAIL.n142 B 0.008528f
C179 VTAIL.t4 B 0.034f
C180 VTAIL.n143 B 0.111312f
C181 VTAIL.n144 B 0.014249f
C182 VTAIL.n145 B 0.015117f
C183 VTAIL.n146 B 0.020156f
C184 VTAIL.n147 B 0.009029f
C185 VTAIL.n148 B 0.008528f
C186 VTAIL.n149 B 0.01587f
C187 VTAIL.n150 B 0.01587f
C188 VTAIL.n151 B 0.008528f
C189 VTAIL.n152 B 0.009029f
C190 VTAIL.n153 B 0.020156f
C191 VTAIL.n154 B 0.020156f
C192 VTAIL.n155 B 0.009029f
C193 VTAIL.n156 B 0.008528f
C194 VTAIL.n157 B 0.01587f
C195 VTAIL.n158 B 0.01587f
C196 VTAIL.n159 B 0.008528f
C197 VTAIL.n160 B 0.008528f
C198 VTAIL.n161 B 0.009029f
C199 VTAIL.n162 B 0.020156f
C200 VTAIL.n163 B 0.020156f
C201 VTAIL.n164 B 0.020156f
C202 VTAIL.n165 B 0.008779f
C203 VTAIL.n166 B 0.008528f
C204 VTAIL.n167 B 0.01587f
C205 VTAIL.n168 B 0.01587f
C206 VTAIL.n169 B 0.008528f
C207 VTAIL.n170 B 0.009029f
C208 VTAIL.n171 B 0.020156f
C209 VTAIL.n172 B 0.020156f
C210 VTAIL.n173 B 0.009029f
C211 VTAIL.n174 B 0.008528f
C212 VTAIL.n175 B 0.01587f
C213 VTAIL.n176 B 0.01587f
C214 VTAIL.n177 B 0.008528f
C215 VTAIL.n178 B 0.009029f
C216 VTAIL.n179 B 0.020156f
C217 VTAIL.n180 B 0.044582f
C218 VTAIL.n181 B 0.009029f
C219 VTAIL.n182 B 0.008528f
C220 VTAIL.n183 B 0.038633f
C221 VTAIL.n184 B 0.025101f
C222 VTAIL.n185 B 0.79581f
C223 VTAIL.n186 B 0.022842f
C224 VTAIL.n187 B 0.01587f
C225 VTAIL.n188 B 0.008528f
C226 VTAIL.n189 B 0.020156f
C227 VTAIL.n190 B 0.009029f
C228 VTAIL.n191 B 0.01587f
C229 VTAIL.n192 B 0.008528f
C230 VTAIL.n193 B 0.020156f
C231 VTAIL.n194 B 0.008779f
C232 VTAIL.n195 B 0.01587f
C233 VTAIL.n196 B 0.008779f
C234 VTAIL.n197 B 0.008528f
C235 VTAIL.n198 B 0.020156f
C236 VTAIL.n199 B 0.020156f
C237 VTAIL.n200 B 0.009029f
C238 VTAIL.n201 B 0.01587f
C239 VTAIL.n202 B 0.008528f
C240 VTAIL.n203 B 0.020156f
C241 VTAIL.n204 B 0.009029f
C242 VTAIL.n205 B 0.764602f
C243 VTAIL.n206 B 0.008528f
C244 VTAIL.t0 B 0.034f
C245 VTAIL.n207 B 0.111312f
C246 VTAIL.n208 B 0.014249f
C247 VTAIL.n209 B 0.015117f
C248 VTAIL.n210 B 0.020156f
C249 VTAIL.n211 B 0.009029f
C250 VTAIL.n212 B 0.008528f
C251 VTAIL.n213 B 0.01587f
C252 VTAIL.n214 B 0.01587f
C253 VTAIL.n215 B 0.008528f
C254 VTAIL.n216 B 0.009029f
C255 VTAIL.n217 B 0.020156f
C256 VTAIL.n218 B 0.020156f
C257 VTAIL.n219 B 0.009029f
C258 VTAIL.n220 B 0.008528f
C259 VTAIL.n221 B 0.01587f
C260 VTAIL.n222 B 0.01587f
C261 VTAIL.n223 B 0.008528f
C262 VTAIL.n224 B 0.009029f
C263 VTAIL.n225 B 0.020156f
C264 VTAIL.n226 B 0.020156f
C265 VTAIL.n227 B 0.009029f
C266 VTAIL.n228 B 0.008528f
C267 VTAIL.n229 B 0.01587f
C268 VTAIL.n230 B 0.01587f
C269 VTAIL.n231 B 0.008528f
C270 VTAIL.n232 B 0.009029f
C271 VTAIL.n233 B 0.020156f
C272 VTAIL.n234 B 0.020156f
C273 VTAIL.n235 B 0.009029f
C274 VTAIL.n236 B 0.008528f
C275 VTAIL.n237 B 0.01587f
C276 VTAIL.n238 B 0.01587f
C277 VTAIL.n239 B 0.008528f
C278 VTAIL.n240 B 0.009029f
C279 VTAIL.n241 B 0.020156f
C280 VTAIL.n242 B 0.044582f
C281 VTAIL.n243 B 0.009029f
C282 VTAIL.n244 B 0.008528f
C283 VTAIL.n245 B 0.038633f
C284 VTAIL.n246 B 0.025101f
C285 VTAIL.n247 B 0.79581f
C286 VTAIL.n248 B 0.022842f
C287 VTAIL.n249 B 0.01587f
C288 VTAIL.n250 B 0.008528f
C289 VTAIL.n251 B 0.020156f
C290 VTAIL.n252 B 0.009029f
C291 VTAIL.n253 B 0.01587f
C292 VTAIL.n254 B 0.008528f
C293 VTAIL.n255 B 0.020156f
C294 VTAIL.n256 B 0.008779f
C295 VTAIL.n257 B 0.01587f
C296 VTAIL.n258 B 0.008779f
C297 VTAIL.n259 B 0.008528f
C298 VTAIL.n260 B 0.020156f
C299 VTAIL.n261 B 0.020156f
C300 VTAIL.n262 B 0.009029f
C301 VTAIL.n263 B 0.01587f
C302 VTAIL.n264 B 0.008528f
C303 VTAIL.n265 B 0.020156f
C304 VTAIL.n266 B 0.009029f
C305 VTAIL.n267 B 0.764602f
C306 VTAIL.n268 B 0.008528f
C307 VTAIL.t2 B 0.034f
C308 VTAIL.n269 B 0.111312f
C309 VTAIL.n270 B 0.014249f
C310 VTAIL.n271 B 0.015117f
C311 VTAIL.n272 B 0.020156f
C312 VTAIL.n273 B 0.009029f
C313 VTAIL.n274 B 0.008528f
C314 VTAIL.n275 B 0.01587f
C315 VTAIL.n276 B 0.01587f
C316 VTAIL.n277 B 0.008528f
C317 VTAIL.n278 B 0.009029f
C318 VTAIL.n279 B 0.020156f
C319 VTAIL.n280 B 0.020156f
C320 VTAIL.n281 B 0.009029f
C321 VTAIL.n282 B 0.008528f
C322 VTAIL.n283 B 0.01587f
C323 VTAIL.n284 B 0.01587f
C324 VTAIL.n285 B 0.008528f
C325 VTAIL.n286 B 0.009029f
C326 VTAIL.n287 B 0.020156f
C327 VTAIL.n288 B 0.020156f
C328 VTAIL.n289 B 0.009029f
C329 VTAIL.n290 B 0.008528f
C330 VTAIL.n291 B 0.01587f
C331 VTAIL.n292 B 0.01587f
C332 VTAIL.n293 B 0.008528f
C333 VTAIL.n294 B 0.009029f
C334 VTAIL.n295 B 0.020156f
C335 VTAIL.n296 B 0.020156f
C336 VTAIL.n297 B 0.009029f
C337 VTAIL.n298 B 0.008528f
C338 VTAIL.n299 B 0.01587f
C339 VTAIL.n300 B 0.01587f
C340 VTAIL.n301 B 0.008528f
C341 VTAIL.n302 B 0.009029f
C342 VTAIL.n303 B 0.020156f
C343 VTAIL.n304 B 0.044582f
C344 VTAIL.n305 B 0.009029f
C345 VTAIL.n306 B 0.008528f
C346 VTAIL.n307 B 0.038633f
C347 VTAIL.n308 B 0.025101f
C348 VTAIL.n309 B 0.067776f
C349 VTAIL.n310 B 0.022842f
C350 VTAIL.n311 B 0.01587f
C351 VTAIL.n312 B 0.008528f
C352 VTAIL.n313 B 0.020156f
C353 VTAIL.n314 B 0.009029f
C354 VTAIL.n315 B 0.01587f
C355 VTAIL.n316 B 0.008528f
C356 VTAIL.n317 B 0.020156f
C357 VTAIL.n318 B 0.008779f
C358 VTAIL.n319 B 0.01587f
C359 VTAIL.n320 B 0.008779f
C360 VTAIL.n321 B 0.008528f
C361 VTAIL.n322 B 0.020156f
C362 VTAIL.n323 B 0.020156f
C363 VTAIL.n324 B 0.009029f
C364 VTAIL.n325 B 0.01587f
C365 VTAIL.n326 B 0.008528f
C366 VTAIL.n327 B 0.020156f
C367 VTAIL.n328 B 0.009029f
C368 VTAIL.n329 B 0.764602f
C369 VTAIL.n330 B 0.008528f
C370 VTAIL.t6 B 0.034f
C371 VTAIL.n331 B 0.111312f
C372 VTAIL.n332 B 0.014249f
C373 VTAIL.n333 B 0.015117f
C374 VTAIL.n334 B 0.020156f
C375 VTAIL.n335 B 0.009029f
C376 VTAIL.n336 B 0.008528f
C377 VTAIL.n337 B 0.01587f
C378 VTAIL.n338 B 0.01587f
C379 VTAIL.n339 B 0.008528f
C380 VTAIL.n340 B 0.009029f
C381 VTAIL.n341 B 0.020156f
C382 VTAIL.n342 B 0.020156f
C383 VTAIL.n343 B 0.009029f
C384 VTAIL.n344 B 0.008528f
C385 VTAIL.n345 B 0.01587f
C386 VTAIL.n346 B 0.01587f
C387 VTAIL.n347 B 0.008528f
C388 VTAIL.n348 B 0.009029f
C389 VTAIL.n349 B 0.020156f
C390 VTAIL.n350 B 0.020156f
C391 VTAIL.n351 B 0.009029f
C392 VTAIL.n352 B 0.008528f
C393 VTAIL.n353 B 0.01587f
C394 VTAIL.n354 B 0.01587f
C395 VTAIL.n355 B 0.008528f
C396 VTAIL.n356 B 0.009029f
C397 VTAIL.n357 B 0.020156f
C398 VTAIL.n358 B 0.020156f
C399 VTAIL.n359 B 0.009029f
C400 VTAIL.n360 B 0.008528f
C401 VTAIL.n361 B 0.01587f
C402 VTAIL.n362 B 0.01587f
C403 VTAIL.n363 B 0.008528f
C404 VTAIL.n364 B 0.009029f
C405 VTAIL.n365 B 0.020156f
C406 VTAIL.n366 B 0.044582f
C407 VTAIL.n367 B 0.009029f
C408 VTAIL.n368 B 0.008528f
C409 VTAIL.n369 B 0.038633f
C410 VTAIL.n370 B 0.025101f
C411 VTAIL.n371 B 0.067776f
C412 VTAIL.n372 B 0.022842f
C413 VTAIL.n373 B 0.01587f
C414 VTAIL.n374 B 0.008528f
C415 VTAIL.n375 B 0.020156f
C416 VTAIL.n376 B 0.009029f
C417 VTAIL.n377 B 0.01587f
C418 VTAIL.n378 B 0.008528f
C419 VTAIL.n379 B 0.020156f
C420 VTAIL.n380 B 0.008779f
C421 VTAIL.n381 B 0.01587f
C422 VTAIL.n382 B 0.008779f
C423 VTAIL.n383 B 0.008528f
C424 VTAIL.n384 B 0.020156f
C425 VTAIL.n385 B 0.020156f
C426 VTAIL.n386 B 0.009029f
C427 VTAIL.n387 B 0.01587f
C428 VTAIL.n388 B 0.008528f
C429 VTAIL.n389 B 0.020156f
C430 VTAIL.n390 B 0.009029f
C431 VTAIL.n391 B 0.764602f
C432 VTAIL.n392 B 0.008528f
C433 VTAIL.t7 B 0.034f
C434 VTAIL.n393 B 0.111312f
C435 VTAIL.n394 B 0.014249f
C436 VTAIL.n395 B 0.015117f
C437 VTAIL.n396 B 0.020156f
C438 VTAIL.n397 B 0.009029f
C439 VTAIL.n398 B 0.008528f
C440 VTAIL.n399 B 0.01587f
C441 VTAIL.n400 B 0.01587f
C442 VTAIL.n401 B 0.008528f
C443 VTAIL.n402 B 0.009029f
C444 VTAIL.n403 B 0.020156f
C445 VTAIL.n404 B 0.020156f
C446 VTAIL.n405 B 0.009029f
C447 VTAIL.n406 B 0.008528f
C448 VTAIL.n407 B 0.01587f
C449 VTAIL.n408 B 0.01587f
C450 VTAIL.n409 B 0.008528f
C451 VTAIL.n410 B 0.009029f
C452 VTAIL.n411 B 0.020156f
C453 VTAIL.n412 B 0.020156f
C454 VTAIL.n413 B 0.009029f
C455 VTAIL.n414 B 0.008528f
C456 VTAIL.n415 B 0.01587f
C457 VTAIL.n416 B 0.01587f
C458 VTAIL.n417 B 0.008528f
C459 VTAIL.n418 B 0.009029f
C460 VTAIL.n419 B 0.020156f
C461 VTAIL.n420 B 0.020156f
C462 VTAIL.n421 B 0.009029f
C463 VTAIL.n422 B 0.008528f
C464 VTAIL.n423 B 0.01587f
C465 VTAIL.n424 B 0.01587f
C466 VTAIL.n425 B 0.008528f
C467 VTAIL.n426 B 0.009029f
C468 VTAIL.n427 B 0.020156f
C469 VTAIL.n428 B 0.044582f
C470 VTAIL.n429 B 0.009029f
C471 VTAIL.n430 B 0.008528f
C472 VTAIL.n431 B 0.038633f
C473 VTAIL.n432 B 0.025101f
C474 VTAIL.n433 B 0.79581f
C475 VTAIL.n434 B 0.022842f
C476 VTAIL.n435 B 0.01587f
C477 VTAIL.n436 B 0.008528f
C478 VTAIL.n437 B 0.020156f
C479 VTAIL.n438 B 0.009029f
C480 VTAIL.n439 B 0.01587f
C481 VTAIL.n440 B 0.008528f
C482 VTAIL.n441 B 0.020156f
C483 VTAIL.n442 B 0.008779f
C484 VTAIL.n443 B 0.01587f
C485 VTAIL.n444 B 0.009029f
C486 VTAIL.n445 B 0.020156f
C487 VTAIL.n446 B 0.009029f
C488 VTAIL.n447 B 0.01587f
C489 VTAIL.n448 B 0.008528f
C490 VTAIL.n449 B 0.020156f
C491 VTAIL.n450 B 0.009029f
C492 VTAIL.n451 B 0.764602f
C493 VTAIL.n452 B 0.008528f
C494 VTAIL.t1 B 0.034f
C495 VTAIL.n453 B 0.111312f
C496 VTAIL.n454 B 0.014249f
C497 VTAIL.n455 B 0.015117f
C498 VTAIL.n456 B 0.020156f
C499 VTAIL.n457 B 0.009029f
C500 VTAIL.n458 B 0.008528f
C501 VTAIL.n459 B 0.01587f
C502 VTAIL.n460 B 0.01587f
C503 VTAIL.n461 B 0.008528f
C504 VTAIL.n462 B 0.009029f
C505 VTAIL.n463 B 0.020156f
C506 VTAIL.n464 B 0.020156f
C507 VTAIL.n465 B 0.009029f
C508 VTAIL.n466 B 0.008528f
C509 VTAIL.n467 B 0.01587f
C510 VTAIL.n468 B 0.01587f
C511 VTAIL.n469 B 0.008528f
C512 VTAIL.n470 B 0.008528f
C513 VTAIL.n471 B 0.009029f
C514 VTAIL.n472 B 0.020156f
C515 VTAIL.n473 B 0.020156f
C516 VTAIL.n474 B 0.020156f
C517 VTAIL.n475 B 0.008779f
C518 VTAIL.n476 B 0.008528f
C519 VTAIL.n477 B 0.01587f
C520 VTAIL.n478 B 0.01587f
C521 VTAIL.n479 B 0.008528f
C522 VTAIL.n480 B 0.009029f
C523 VTAIL.n481 B 0.020156f
C524 VTAIL.n482 B 0.020156f
C525 VTAIL.n483 B 0.009029f
C526 VTAIL.n484 B 0.008528f
C527 VTAIL.n485 B 0.01587f
C528 VTAIL.n486 B 0.01587f
C529 VTAIL.n487 B 0.008528f
C530 VTAIL.n488 B 0.009029f
C531 VTAIL.n489 B 0.020156f
C532 VTAIL.n490 B 0.044582f
C533 VTAIL.n491 B 0.009029f
C534 VTAIL.n492 B 0.008528f
C535 VTAIL.n493 B 0.038633f
C536 VTAIL.n494 B 0.025101f
C537 VTAIL.n495 B 0.778287f
C538 VP.t2 B 0.540873f
C539 VP.t0 B 0.540873f
C540 VP.n0 B 0.784165f
C541 VP.t1 B 0.540873f
C542 VP.t3 B 0.540873f
C543 VP.n1 B 0.430769f
C544 VP.n2 B 3.2955f
.ends

