* NGSPICE file created from diff_pair_sample_1542.ext - technology: sky130A

.subckt diff_pair_sample_1542 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t9 w_n3680_n1438# sky130_fd_pr__pfet_01v8 ad=0.38775 pd=2.68 as=0.9165 ps=5.48 w=2.35 l=2.38
X1 VDD1.t6 VP.t1 VTAIL.t12 w_n3680_n1438# sky130_fd_pr__pfet_01v8 ad=0.38775 pd=2.68 as=0.38775 ps=2.68 w=2.35 l=2.38
X2 VTAIL.t3 VN.t0 VDD2.t7 w_n3680_n1438# sky130_fd_pr__pfet_01v8 ad=0.38775 pd=2.68 as=0.38775 ps=2.68 w=2.35 l=2.38
X3 VTAIL.t7 VN.t1 VDD2.t6 w_n3680_n1438# sky130_fd_pr__pfet_01v8 ad=0.9165 pd=5.48 as=0.38775 ps=2.68 w=2.35 l=2.38
X4 VDD2.t5 VN.t2 VTAIL.t1 w_n3680_n1438# sky130_fd_pr__pfet_01v8 ad=0.38775 pd=2.68 as=0.9165 ps=5.48 w=2.35 l=2.38
X5 VTAIL.t11 VP.t2 VDD1.t5 w_n3680_n1438# sky130_fd_pr__pfet_01v8 ad=0.9165 pd=5.48 as=0.38775 ps=2.68 w=2.35 l=2.38
X6 VDD1.t4 VP.t3 VTAIL.t13 w_n3680_n1438# sky130_fd_pr__pfet_01v8 ad=0.38775 pd=2.68 as=0.9165 ps=5.48 w=2.35 l=2.38
X7 VDD1.t3 VP.t4 VTAIL.t10 w_n3680_n1438# sky130_fd_pr__pfet_01v8 ad=0.38775 pd=2.68 as=0.38775 ps=2.68 w=2.35 l=2.38
X8 VDD2.t4 VN.t3 VTAIL.t2 w_n3680_n1438# sky130_fd_pr__pfet_01v8 ad=0.38775 pd=2.68 as=0.9165 ps=5.48 w=2.35 l=2.38
X9 VTAIL.t14 VP.t5 VDD1.t2 w_n3680_n1438# sky130_fd_pr__pfet_01v8 ad=0.38775 pd=2.68 as=0.38775 ps=2.68 w=2.35 l=2.38
X10 B.t11 B.t9 B.t10 w_n3680_n1438# sky130_fd_pr__pfet_01v8 ad=0.9165 pd=5.48 as=0 ps=0 w=2.35 l=2.38
X11 VDD2.t3 VN.t4 VTAIL.t6 w_n3680_n1438# sky130_fd_pr__pfet_01v8 ad=0.38775 pd=2.68 as=0.38775 ps=2.68 w=2.35 l=2.38
X12 VTAIL.t15 VP.t6 VDD1.t1 w_n3680_n1438# sky130_fd_pr__pfet_01v8 ad=0.38775 pd=2.68 as=0.38775 ps=2.68 w=2.35 l=2.38
X13 VTAIL.t5 VN.t5 VDD2.t2 w_n3680_n1438# sky130_fd_pr__pfet_01v8 ad=0.9165 pd=5.48 as=0.38775 ps=2.68 w=2.35 l=2.38
X14 VTAIL.t8 VP.t7 VDD1.t0 w_n3680_n1438# sky130_fd_pr__pfet_01v8 ad=0.9165 pd=5.48 as=0.38775 ps=2.68 w=2.35 l=2.38
X15 B.t8 B.t6 B.t7 w_n3680_n1438# sky130_fd_pr__pfet_01v8 ad=0.9165 pd=5.48 as=0 ps=0 w=2.35 l=2.38
X16 VDD2.t1 VN.t6 VTAIL.t0 w_n3680_n1438# sky130_fd_pr__pfet_01v8 ad=0.38775 pd=2.68 as=0.38775 ps=2.68 w=2.35 l=2.38
X17 B.t5 B.t3 B.t4 w_n3680_n1438# sky130_fd_pr__pfet_01v8 ad=0.9165 pd=5.48 as=0 ps=0 w=2.35 l=2.38
X18 VTAIL.t4 VN.t7 VDD2.t0 w_n3680_n1438# sky130_fd_pr__pfet_01v8 ad=0.38775 pd=2.68 as=0.38775 ps=2.68 w=2.35 l=2.38
X19 B.t2 B.t0 B.t1 w_n3680_n1438# sky130_fd_pr__pfet_01v8 ad=0.9165 pd=5.48 as=0 ps=0 w=2.35 l=2.38
R0 VP.n16 VP.n13 161.3
R1 VP.n18 VP.n17 161.3
R2 VP.n19 VP.n12 161.3
R3 VP.n21 VP.n20 161.3
R4 VP.n22 VP.n11 161.3
R5 VP.n24 VP.n23 161.3
R6 VP.n26 VP.n10 161.3
R7 VP.n28 VP.n27 161.3
R8 VP.n29 VP.n9 161.3
R9 VP.n31 VP.n30 161.3
R10 VP.n32 VP.n8 161.3
R11 VP.n62 VP.n0 161.3
R12 VP.n61 VP.n60 161.3
R13 VP.n59 VP.n1 161.3
R14 VP.n58 VP.n57 161.3
R15 VP.n56 VP.n2 161.3
R16 VP.n54 VP.n53 161.3
R17 VP.n52 VP.n3 161.3
R18 VP.n51 VP.n50 161.3
R19 VP.n49 VP.n4 161.3
R20 VP.n48 VP.n47 161.3
R21 VP.n46 VP.n5 161.3
R22 VP.n45 VP.n44 161.3
R23 VP.n42 VP.n6 161.3
R24 VP.n41 VP.n40 161.3
R25 VP.n39 VP.n7 161.3
R26 VP.n38 VP.n37 161.3
R27 VP.n36 VP.n35 95.3422
R28 VP.n64 VP.n63 95.3422
R29 VP.n34 VP.n33 95.3422
R30 VP.n15 VP.n14 66.9989
R31 VP.n50 VP.n49 56.5193
R32 VP.n20 VP.n19 56.5193
R33 VP.n15 VP.t7 56.4278
R34 VP.n42 VP.n41 44.3785
R35 VP.n57 VP.n1 44.3785
R36 VP.n27 VP.n9 44.3785
R37 VP.n35 VP.n34 42.6056
R38 VP.n41 VP.n7 36.6083
R39 VP.n61 VP.n1 36.6083
R40 VP.n31 VP.n9 36.6083
R41 VP.n37 VP.n7 24.4675
R42 VP.n44 VP.n42 24.4675
R43 VP.n48 VP.n5 24.4675
R44 VP.n49 VP.n48 24.4675
R45 VP.n50 VP.n3 24.4675
R46 VP.n54 VP.n3 24.4675
R47 VP.n57 VP.n56 24.4675
R48 VP.n62 VP.n61 24.4675
R49 VP.n32 VP.n31 24.4675
R50 VP.n20 VP.n11 24.4675
R51 VP.n24 VP.n11 24.4675
R52 VP.n27 VP.n26 24.4675
R53 VP.n18 VP.n13 24.4675
R54 VP.n19 VP.n18 24.4675
R55 VP.n36 VP.t2 23.7967
R56 VP.n43 VP.t1 23.7967
R57 VP.n55 VP.t5 23.7967
R58 VP.n63 VP.t3 23.7967
R59 VP.n33 VP.t0 23.7967
R60 VP.n25 VP.t6 23.7967
R61 VP.n14 VP.t4 23.7967
R62 VP.n44 VP.n43 19.3294
R63 VP.n56 VP.n55 19.3294
R64 VP.n26 VP.n25 19.3294
R65 VP.n37 VP.n36 15.4147
R66 VP.n63 VP.n62 15.4147
R67 VP.n33 VP.n32 15.4147
R68 VP.n16 VP.n15 9.45072
R69 VP.n43 VP.n5 5.13857
R70 VP.n55 VP.n54 5.13857
R71 VP.n25 VP.n24 5.13857
R72 VP.n14 VP.n13 5.13857
R73 VP.n34 VP.n8 0.278367
R74 VP.n38 VP.n35 0.278367
R75 VP.n64 VP.n0 0.278367
R76 VP.n17 VP.n16 0.189894
R77 VP.n17 VP.n12 0.189894
R78 VP.n21 VP.n12 0.189894
R79 VP.n22 VP.n21 0.189894
R80 VP.n23 VP.n22 0.189894
R81 VP.n23 VP.n10 0.189894
R82 VP.n28 VP.n10 0.189894
R83 VP.n29 VP.n28 0.189894
R84 VP.n30 VP.n29 0.189894
R85 VP.n30 VP.n8 0.189894
R86 VP.n39 VP.n38 0.189894
R87 VP.n40 VP.n39 0.189894
R88 VP.n40 VP.n6 0.189894
R89 VP.n45 VP.n6 0.189894
R90 VP.n46 VP.n45 0.189894
R91 VP.n47 VP.n46 0.189894
R92 VP.n47 VP.n4 0.189894
R93 VP.n51 VP.n4 0.189894
R94 VP.n52 VP.n51 0.189894
R95 VP.n53 VP.n52 0.189894
R96 VP.n53 VP.n2 0.189894
R97 VP.n58 VP.n2 0.189894
R98 VP.n59 VP.n58 0.189894
R99 VP.n60 VP.n59 0.189894
R100 VP.n60 VP.n0 0.189894
R101 VP VP.n64 0.153454
R102 VTAIL.n11 VTAIL.t8 168.7
R103 VTAIL.n10 VTAIL.t2 168.7
R104 VTAIL.n7 VTAIL.t7 168.7
R105 VTAIL.n14 VTAIL.t9 168.7
R106 VTAIL.n15 VTAIL.t1 168.698
R107 VTAIL.n2 VTAIL.t5 168.698
R108 VTAIL.n3 VTAIL.t13 168.698
R109 VTAIL.n6 VTAIL.t11 168.698
R110 VTAIL.n13 VTAIL.n12 154.868
R111 VTAIL.n9 VTAIL.n8 154.868
R112 VTAIL.n1 VTAIL.n0 154.868
R113 VTAIL.n5 VTAIL.n4 154.868
R114 VTAIL.n15 VTAIL.n14 16.7289
R115 VTAIL.n7 VTAIL.n6 16.7289
R116 VTAIL.n0 VTAIL.t0 13.8324
R117 VTAIL.n0 VTAIL.t4 13.8324
R118 VTAIL.n4 VTAIL.t12 13.8324
R119 VTAIL.n4 VTAIL.t14 13.8324
R120 VTAIL.n12 VTAIL.t10 13.8324
R121 VTAIL.n12 VTAIL.t15 13.8324
R122 VTAIL.n8 VTAIL.t6 13.8324
R123 VTAIL.n8 VTAIL.t3 13.8324
R124 VTAIL.n9 VTAIL.n7 2.33671
R125 VTAIL.n10 VTAIL.n9 2.33671
R126 VTAIL.n13 VTAIL.n11 2.33671
R127 VTAIL.n14 VTAIL.n13 2.33671
R128 VTAIL.n6 VTAIL.n5 2.33671
R129 VTAIL.n5 VTAIL.n3 2.33671
R130 VTAIL.n2 VTAIL.n1 2.33671
R131 VTAIL VTAIL.n15 2.27852
R132 VTAIL.n11 VTAIL.n10 0.470328
R133 VTAIL.n3 VTAIL.n2 0.470328
R134 VTAIL VTAIL.n1 0.0586897
R135 VDD1 VDD1.n0 172.773
R136 VDD1.n3 VDD1.n2 172.659
R137 VDD1.n3 VDD1.n1 172.659
R138 VDD1.n5 VDD1.n4 171.546
R139 VDD1.n5 VDD1.n3 36.8371
R140 VDD1.n4 VDD1.t1 13.8324
R141 VDD1.n4 VDD1.t7 13.8324
R142 VDD1.n0 VDD1.t0 13.8324
R143 VDD1.n0 VDD1.t3 13.8324
R144 VDD1.n2 VDD1.t2 13.8324
R145 VDD1.n2 VDD1.t4 13.8324
R146 VDD1.n1 VDD1.t5 13.8324
R147 VDD1.n1 VDD1.t6 13.8324
R148 VDD1 VDD1.n5 1.11041
R149 VN.n51 VN.n27 161.3
R150 VN.n50 VN.n49 161.3
R151 VN.n48 VN.n28 161.3
R152 VN.n47 VN.n46 161.3
R153 VN.n45 VN.n29 161.3
R154 VN.n43 VN.n42 161.3
R155 VN.n41 VN.n30 161.3
R156 VN.n40 VN.n39 161.3
R157 VN.n38 VN.n31 161.3
R158 VN.n37 VN.n36 161.3
R159 VN.n35 VN.n32 161.3
R160 VN.n24 VN.n0 161.3
R161 VN.n23 VN.n22 161.3
R162 VN.n21 VN.n1 161.3
R163 VN.n20 VN.n19 161.3
R164 VN.n18 VN.n2 161.3
R165 VN.n16 VN.n15 161.3
R166 VN.n14 VN.n3 161.3
R167 VN.n13 VN.n12 161.3
R168 VN.n11 VN.n4 161.3
R169 VN.n10 VN.n9 161.3
R170 VN.n8 VN.n5 161.3
R171 VN.n26 VN.n25 95.3422
R172 VN.n53 VN.n52 95.3422
R173 VN.n7 VN.n6 66.9989
R174 VN.n34 VN.n33 66.9989
R175 VN.n12 VN.n11 56.5193
R176 VN.n39 VN.n38 56.5193
R177 VN.n7 VN.t5 56.4278
R178 VN.n34 VN.t3 56.4278
R179 VN.n19 VN.n1 44.3785
R180 VN.n46 VN.n28 44.3785
R181 VN VN.n53 42.8845
R182 VN.n23 VN.n1 36.6083
R183 VN.n50 VN.n28 36.6083
R184 VN.n10 VN.n5 24.4675
R185 VN.n11 VN.n10 24.4675
R186 VN.n12 VN.n3 24.4675
R187 VN.n16 VN.n3 24.4675
R188 VN.n19 VN.n18 24.4675
R189 VN.n24 VN.n23 24.4675
R190 VN.n38 VN.n37 24.4675
R191 VN.n37 VN.n32 24.4675
R192 VN.n46 VN.n45 24.4675
R193 VN.n43 VN.n30 24.4675
R194 VN.n39 VN.n30 24.4675
R195 VN.n51 VN.n50 24.4675
R196 VN.n6 VN.t6 23.7967
R197 VN.n17 VN.t7 23.7967
R198 VN.n25 VN.t2 23.7967
R199 VN.n33 VN.t0 23.7967
R200 VN.n44 VN.t4 23.7967
R201 VN.n52 VN.t1 23.7967
R202 VN.n18 VN.n17 19.3294
R203 VN.n45 VN.n44 19.3294
R204 VN.n25 VN.n24 15.4147
R205 VN.n52 VN.n51 15.4147
R206 VN.n35 VN.n34 9.45072
R207 VN.n8 VN.n7 9.45072
R208 VN.n6 VN.n5 5.13857
R209 VN.n17 VN.n16 5.13857
R210 VN.n33 VN.n32 5.13857
R211 VN.n44 VN.n43 5.13857
R212 VN.n53 VN.n27 0.278367
R213 VN.n26 VN.n0 0.278367
R214 VN.n49 VN.n27 0.189894
R215 VN.n49 VN.n48 0.189894
R216 VN.n48 VN.n47 0.189894
R217 VN.n47 VN.n29 0.189894
R218 VN.n42 VN.n29 0.189894
R219 VN.n42 VN.n41 0.189894
R220 VN.n41 VN.n40 0.189894
R221 VN.n40 VN.n31 0.189894
R222 VN.n36 VN.n31 0.189894
R223 VN.n36 VN.n35 0.189894
R224 VN.n9 VN.n8 0.189894
R225 VN.n9 VN.n4 0.189894
R226 VN.n13 VN.n4 0.189894
R227 VN.n14 VN.n13 0.189894
R228 VN.n15 VN.n14 0.189894
R229 VN.n15 VN.n2 0.189894
R230 VN.n20 VN.n2 0.189894
R231 VN.n21 VN.n20 0.189894
R232 VN.n22 VN.n21 0.189894
R233 VN.n22 VN.n0 0.189894
R234 VN VN.n26 0.153454
R235 VDD2.n2 VDD2.n1 172.659
R236 VDD2.n2 VDD2.n0 172.659
R237 VDD2 VDD2.n5 172.655
R238 VDD2.n4 VDD2.n3 171.546
R239 VDD2.n4 VDD2.n2 36.2541
R240 VDD2.n5 VDD2.t7 13.8324
R241 VDD2.n5 VDD2.t4 13.8324
R242 VDD2.n3 VDD2.t6 13.8324
R243 VDD2.n3 VDD2.t3 13.8324
R244 VDD2.n1 VDD2.t0 13.8324
R245 VDD2.n1 VDD2.t5 13.8324
R246 VDD2.n0 VDD2.t2 13.8324
R247 VDD2.n0 VDD2.t1 13.8324
R248 VDD2 VDD2.n4 1.22679
R249 B.n416 B.n415 585
R250 B.n417 B.n48 585
R251 B.n419 B.n418 585
R252 B.n420 B.n47 585
R253 B.n422 B.n421 585
R254 B.n423 B.n46 585
R255 B.n425 B.n424 585
R256 B.n426 B.n45 585
R257 B.n428 B.n427 585
R258 B.n429 B.n44 585
R259 B.n431 B.n430 585
R260 B.n432 B.n43 585
R261 B.n434 B.n433 585
R262 B.n436 B.n40 585
R263 B.n438 B.n437 585
R264 B.n439 B.n39 585
R265 B.n441 B.n440 585
R266 B.n442 B.n38 585
R267 B.n444 B.n443 585
R268 B.n445 B.n37 585
R269 B.n447 B.n446 585
R270 B.n448 B.n33 585
R271 B.n450 B.n449 585
R272 B.n451 B.n32 585
R273 B.n453 B.n452 585
R274 B.n454 B.n31 585
R275 B.n456 B.n455 585
R276 B.n457 B.n30 585
R277 B.n459 B.n458 585
R278 B.n460 B.n29 585
R279 B.n462 B.n461 585
R280 B.n463 B.n28 585
R281 B.n465 B.n464 585
R282 B.n466 B.n27 585
R283 B.n468 B.n467 585
R284 B.n469 B.n26 585
R285 B.n414 B.n49 585
R286 B.n413 B.n412 585
R287 B.n411 B.n50 585
R288 B.n410 B.n409 585
R289 B.n408 B.n51 585
R290 B.n407 B.n406 585
R291 B.n405 B.n52 585
R292 B.n404 B.n403 585
R293 B.n402 B.n53 585
R294 B.n401 B.n400 585
R295 B.n399 B.n54 585
R296 B.n398 B.n397 585
R297 B.n396 B.n55 585
R298 B.n395 B.n394 585
R299 B.n393 B.n56 585
R300 B.n392 B.n391 585
R301 B.n390 B.n57 585
R302 B.n389 B.n388 585
R303 B.n387 B.n58 585
R304 B.n386 B.n385 585
R305 B.n384 B.n59 585
R306 B.n383 B.n382 585
R307 B.n381 B.n60 585
R308 B.n380 B.n379 585
R309 B.n378 B.n61 585
R310 B.n377 B.n376 585
R311 B.n375 B.n62 585
R312 B.n374 B.n373 585
R313 B.n372 B.n63 585
R314 B.n371 B.n370 585
R315 B.n369 B.n64 585
R316 B.n368 B.n367 585
R317 B.n366 B.n65 585
R318 B.n365 B.n364 585
R319 B.n363 B.n66 585
R320 B.n362 B.n361 585
R321 B.n360 B.n67 585
R322 B.n359 B.n358 585
R323 B.n357 B.n68 585
R324 B.n356 B.n355 585
R325 B.n354 B.n69 585
R326 B.n353 B.n352 585
R327 B.n351 B.n70 585
R328 B.n350 B.n349 585
R329 B.n348 B.n71 585
R330 B.n347 B.n346 585
R331 B.n345 B.n72 585
R332 B.n344 B.n343 585
R333 B.n342 B.n73 585
R334 B.n341 B.n340 585
R335 B.n339 B.n74 585
R336 B.n338 B.n337 585
R337 B.n336 B.n75 585
R338 B.n335 B.n334 585
R339 B.n333 B.n76 585
R340 B.n332 B.n331 585
R341 B.n330 B.n77 585
R342 B.n329 B.n328 585
R343 B.n327 B.n78 585
R344 B.n326 B.n325 585
R345 B.n324 B.n79 585
R346 B.n323 B.n322 585
R347 B.n321 B.n80 585
R348 B.n320 B.n319 585
R349 B.n318 B.n81 585
R350 B.n317 B.n316 585
R351 B.n315 B.n82 585
R352 B.n314 B.n313 585
R353 B.n312 B.n83 585
R354 B.n311 B.n310 585
R355 B.n309 B.n84 585
R356 B.n308 B.n307 585
R357 B.n306 B.n85 585
R358 B.n305 B.n304 585
R359 B.n303 B.n86 585
R360 B.n302 B.n301 585
R361 B.n300 B.n87 585
R362 B.n299 B.n298 585
R363 B.n297 B.n88 585
R364 B.n296 B.n295 585
R365 B.n294 B.n89 585
R366 B.n293 B.n292 585
R367 B.n291 B.n90 585
R368 B.n290 B.n289 585
R369 B.n288 B.n91 585
R370 B.n287 B.n286 585
R371 B.n285 B.n92 585
R372 B.n284 B.n283 585
R373 B.n282 B.n93 585
R374 B.n281 B.n280 585
R375 B.n279 B.n94 585
R376 B.n278 B.n277 585
R377 B.n276 B.n95 585
R378 B.n275 B.n274 585
R379 B.n273 B.n96 585
R380 B.n272 B.n271 585
R381 B.n270 B.n97 585
R382 B.n215 B.n214 585
R383 B.n216 B.n119 585
R384 B.n218 B.n217 585
R385 B.n219 B.n118 585
R386 B.n221 B.n220 585
R387 B.n222 B.n117 585
R388 B.n224 B.n223 585
R389 B.n225 B.n116 585
R390 B.n227 B.n226 585
R391 B.n228 B.n115 585
R392 B.n230 B.n229 585
R393 B.n231 B.n114 585
R394 B.n233 B.n232 585
R395 B.n235 B.n234 585
R396 B.n236 B.n110 585
R397 B.n238 B.n237 585
R398 B.n239 B.n109 585
R399 B.n241 B.n240 585
R400 B.n242 B.n108 585
R401 B.n244 B.n243 585
R402 B.n245 B.n107 585
R403 B.n247 B.n246 585
R404 B.n248 B.n104 585
R405 B.n251 B.n250 585
R406 B.n252 B.n103 585
R407 B.n254 B.n253 585
R408 B.n255 B.n102 585
R409 B.n257 B.n256 585
R410 B.n258 B.n101 585
R411 B.n260 B.n259 585
R412 B.n261 B.n100 585
R413 B.n263 B.n262 585
R414 B.n264 B.n99 585
R415 B.n266 B.n265 585
R416 B.n267 B.n98 585
R417 B.n269 B.n268 585
R418 B.n213 B.n120 585
R419 B.n212 B.n211 585
R420 B.n210 B.n121 585
R421 B.n209 B.n208 585
R422 B.n207 B.n122 585
R423 B.n206 B.n205 585
R424 B.n204 B.n123 585
R425 B.n203 B.n202 585
R426 B.n201 B.n124 585
R427 B.n200 B.n199 585
R428 B.n198 B.n125 585
R429 B.n197 B.n196 585
R430 B.n195 B.n126 585
R431 B.n194 B.n193 585
R432 B.n192 B.n127 585
R433 B.n191 B.n190 585
R434 B.n189 B.n128 585
R435 B.n188 B.n187 585
R436 B.n186 B.n129 585
R437 B.n185 B.n184 585
R438 B.n183 B.n130 585
R439 B.n182 B.n181 585
R440 B.n180 B.n131 585
R441 B.n179 B.n178 585
R442 B.n177 B.n132 585
R443 B.n176 B.n175 585
R444 B.n174 B.n133 585
R445 B.n173 B.n172 585
R446 B.n171 B.n134 585
R447 B.n170 B.n169 585
R448 B.n168 B.n135 585
R449 B.n167 B.n166 585
R450 B.n165 B.n136 585
R451 B.n164 B.n163 585
R452 B.n162 B.n137 585
R453 B.n161 B.n160 585
R454 B.n159 B.n138 585
R455 B.n158 B.n157 585
R456 B.n156 B.n139 585
R457 B.n155 B.n154 585
R458 B.n153 B.n140 585
R459 B.n152 B.n151 585
R460 B.n150 B.n141 585
R461 B.n149 B.n148 585
R462 B.n147 B.n142 585
R463 B.n146 B.n145 585
R464 B.n144 B.n143 585
R465 B.n2 B.n0 585
R466 B.n541 B.n1 585
R467 B.n540 B.n539 585
R468 B.n538 B.n3 585
R469 B.n537 B.n536 585
R470 B.n535 B.n4 585
R471 B.n534 B.n533 585
R472 B.n532 B.n5 585
R473 B.n531 B.n530 585
R474 B.n529 B.n6 585
R475 B.n528 B.n527 585
R476 B.n526 B.n7 585
R477 B.n525 B.n524 585
R478 B.n523 B.n8 585
R479 B.n522 B.n521 585
R480 B.n520 B.n9 585
R481 B.n519 B.n518 585
R482 B.n517 B.n10 585
R483 B.n516 B.n515 585
R484 B.n514 B.n11 585
R485 B.n513 B.n512 585
R486 B.n511 B.n12 585
R487 B.n510 B.n509 585
R488 B.n508 B.n13 585
R489 B.n507 B.n506 585
R490 B.n505 B.n14 585
R491 B.n504 B.n503 585
R492 B.n502 B.n15 585
R493 B.n501 B.n500 585
R494 B.n499 B.n16 585
R495 B.n498 B.n497 585
R496 B.n496 B.n17 585
R497 B.n495 B.n494 585
R498 B.n493 B.n18 585
R499 B.n492 B.n491 585
R500 B.n490 B.n19 585
R501 B.n489 B.n488 585
R502 B.n487 B.n20 585
R503 B.n486 B.n485 585
R504 B.n484 B.n21 585
R505 B.n483 B.n482 585
R506 B.n481 B.n22 585
R507 B.n480 B.n479 585
R508 B.n478 B.n23 585
R509 B.n477 B.n476 585
R510 B.n475 B.n24 585
R511 B.n474 B.n473 585
R512 B.n472 B.n25 585
R513 B.n471 B.n470 585
R514 B.n543 B.n542 585
R515 B.n215 B.n120 497.305
R516 B.n470 B.n469 497.305
R517 B.n270 B.n269 497.305
R518 B.n415 B.n414 497.305
R519 B.n105 B.t0 231.486
R520 B.n111 B.t6 231.486
R521 B.n34 B.t9 231.486
R522 B.n41 B.t3 231.486
R523 B.n105 B.t2 227.371
R524 B.n41 B.t4 227.371
R525 B.n111 B.t8 227.371
R526 B.n34 B.t10 227.371
R527 B.n106 B.t1 174.815
R528 B.n42 B.t5 174.815
R529 B.n112 B.t7 174.814
R530 B.n35 B.t11 174.814
R531 B.n211 B.n120 163.367
R532 B.n211 B.n210 163.367
R533 B.n210 B.n209 163.367
R534 B.n209 B.n122 163.367
R535 B.n205 B.n122 163.367
R536 B.n205 B.n204 163.367
R537 B.n204 B.n203 163.367
R538 B.n203 B.n124 163.367
R539 B.n199 B.n124 163.367
R540 B.n199 B.n198 163.367
R541 B.n198 B.n197 163.367
R542 B.n197 B.n126 163.367
R543 B.n193 B.n126 163.367
R544 B.n193 B.n192 163.367
R545 B.n192 B.n191 163.367
R546 B.n191 B.n128 163.367
R547 B.n187 B.n128 163.367
R548 B.n187 B.n186 163.367
R549 B.n186 B.n185 163.367
R550 B.n185 B.n130 163.367
R551 B.n181 B.n130 163.367
R552 B.n181 B.n180 163.367
R553 B.n180 B.n179 163.367
R554 B.n179 B.n132 163.367
R555 B.n175 B.n132 163.367
R556 B.n175 B.n174 163.367
R557 B.n174 B.n173 163.367
R558 B.n173 B.n134 163.367
R559 B.n169 B.n134 163.367
R560 B.n169 B.n168 163.367
R561 B.n168 B.n167 163.367
R562 B.n167 B.n136 163.367
R563 B.n163 B.n136 163.367
R564 B.n163 B.n162 163.367
R565 B.n162 B.n161 163.367
R566 B.n161 B.n138 163.367
R567 B.n157 B.n138 163.367
R568 B.n157 B.n156 163.367
R569 B.n156 B.n155 163.367
R570 B.n155 B.n140 163.367
R571 B.n151 B.n140 163.367
R572 B.n151 B.n150 163.367
R573 B.n150 B.n149 163.367
R574 B.n149 B.n142 163.367
R575 B.n145 B.n142 163.367
R576 B.n145 B.n144 163.367
R577 B.n144 B.n2 163.367
R578 B.n542 B.n2 163.367
R579 B.n542 B.n541 163.367
R580 B.n541 B.n540 163.367
R581 B.n540 B.n3 163.367
R582 B.n536 B.n3 163.367
R583 B.n536 B.n535 163.367
R584 B.n535 B.n534 163.367
R585 B.n534 B.n5 163.367
R586 B.n530 B.n5 163.367
R587 B.n530 B.n529 163.367
R588 B.n529 B.n528 163.367
R589 B.n528 B.n7 163.367
R590 B.n524 B.n7 163.367
R591 B.n524 B.n523 163.367
R592 B.n523 B.n522 163.367
R593 B.n522 B.n9 163.367
R594 B.n518 B.n9 163.367
R595 B.n518 B.n517 163.367
R596 B.n517 B.n516 163.367
R597 B.n516 B.n11 163.367
R598 B.n512 B.n11 163.367
R599 B.n512 B.n511 163.367
R600 B.n511 B.n510 163.367
R601 B.n510 B.n13 163.367
R602 B.n506 B.n13 163.367
R603 B.n506 B.n505 163.367
R604 B.n505 B.n504 163.367
R605 B.n504 B.n15 163.367
R606 B.n500 B.n15 163.367
R607 B.n500 B.n499 163.367
R608 B.n499 B.n498 163.367
R609 B.n498 B.n17 163.367
R610 B.n494 B.n17 163.367
R611 B.n494 B.n493 163.367
R612 B.n493 B.n492 163.367
R613 B.n492 B.n19 163.367
R614 B.n488 B.n19 163.367
R615 B.n488 B.n487 163.367
R616 B.n487 B.n486 163.367
R617 B.n486 B.n21 163.367
R618 B.n482 B.n21 163.367
R619 B.n482 B.n481 163.367
R620 B.n481 B.n480 163.367
R621 B.n480 B.n23 163.367
R622 B.n476 B.n23 163.367
R623 B.n476 B.n475 163.367
R624 B.n475 B.n474 163.367
R625 B.n474 B.n25 163.367
R626 B.n470 B.n25 163.367
R627 B.n216 B.n215 163.367
R628 B.n217 B.n216 163.367
R629 B.n217 B.n118 163.367
R630 B.n221 B.n118 163.367
R631 B.n222 B.n221 163.367
R632 B.n223 B.n222 163.367
R633 B.n223 B.n116 163.367
R634 B.n227 B.n116 163.367
R635 B.n228 B.n227 163.367
R636 B.n229 B.n228 163.367
R637 B.n229 B.n114 163.367
R638 B.n233 B.n114 163.367
R639 B.n234 B.n233 163.367
R640 B.n234 B.n110 163.367
R641 B.n238 B.n110 163.367
R642 B.n239 B.n238 163.367
R643 B.n240 B.n239 163.367
R644 B.n240 B.n108 163.367
R645 B.n244 B.n108 163.367
R646 B.n245 B.n244 163.367
R647 B.n246 B.n245 163.367
R648 B.n246 B.n104 163.367
R649 B.n251 B.n104 163.367
R650 B.n252 B.n251 163.367
R651 B.n253 B.n252 163.367
R652 B.n253 B.n102 163.367
R653 B.n257 B.n102 163.367
R654 B.n258 B.n257 163.367
R655 B.n259 B.n258 163.367
R656 B.n259 B.n100 163.367
R657 B.n263 B.n100 163.367
R658 B.n264 B.n263 163.367
R659 B.n265 B.n264 163.367
R660 B.n265 B.n98 163.367
R661 B.n269 B.n98 163.367
R662 B.n271 B.n270 163.367
R663 B.n271 B.n96 163.367
R664 B.n275 B.n96 163.367
R665 B.n276 B.n275 163.367
R666 B.n277 B.n276 163.367
R667 B.n277 B.n94 163.367
R668 B.n281 B.n94 163.367
R669 B.n282 B.n281 163.367
R670 B.n283 B.n282 163.367
R671 B.n283 B.n92 163.367
R672 B.n287 B.n92 163.367
R673 B.n288 B.n287 163.367
R674 B.n289 B.n288 163.367
R675 B.n289 B.n90 163.367
R676 B.n293 B.n90 163.367
R677 B.n294 B.n293 163.367
R678 B.n295 B.n294 163.367
R679 B.n295 B.n88 163.367
R680 B.n299 B.n88 163.367
R681 B.n300 B.n299 163.367
R682 B.n301 B.n300 163.367
R683 B.n301 B.n86 163.367
R684 B.n305 B.n86 163.367
R685 B.n306 B.n305 163.367
R686 B.n307 B.n306 163.367
R687 B.n307 B.n84 163.367
R688 B.n311 B.n84 163.367
R689 B.n312 B.n311 163.367
R690 B.n313 B.n312 163.367
R691 B.n313 B.n82 163.367
R692 B.n317 B.n82 163.367
R693 B.n318 B.n317 163.367
R694 B.n319 B.n318 163.367
R695 B.n319 B.n80 163.367
R696 B.n323 B.n80 163.367
R697 B.n324 B.n323 163.367
R698 B.n325 B.n324 163.367
R699 B.n325 B.n78 163.367
R700 B.n329 B.n78 163.367
R701 B.n330 B.n329 163.367
R702 B.n331 B.n330 163.367
R703 B.n331 B.n76 163.367
R704 B.n335 B.n76 163.367
R705 B.n336 B.n335 163.367
R706 B.n337 B.n336 163.367
R707 B.n337 B.n74 163.367
R708 B.n341 B.n74 163.367
R709 B.n342 B.n341 163.367
R710 B.n343 B.n342 163.367
R711 B.n343 B.n72 163.367
R712 B.n347 B.n72 163.367
R713 B.n348 B.n347 163.367
R714 B.n349 B.n348 163.367
R715 B.n349 B.n70 163.367
R716 B.n353 B.n70 163.367
R717 B.n354 B.n353 163.367
R718 B.n355 B.n354 163.367
R719 B.n355 B.n68 163.367
R720 B.n359 B.n68 163.367
R721 B.n360 B.n359 163.367
R722 B.n361 B.n360 163.367
R723 B.n361 B.n66 163.367
R724 B.n365 B.n66 163.367
R725 B.n366 B.n365 163.367
R726 B.n367 B.n366 163.367
R727 B.n367 B.n64 163.367
R728 B.n371 B.n64 163.367
R729 B.n372 B.n371 163.367
R730 B.n373 B.n372 163.367
R731 B.n373 B.n62 163.367
R732 B.n377 B.n62 163.367
R733 B.n378 B.n377 163.367
R734 B.n379 B.n378 163.367
R735 B.n379 B.n60 163.367
R736 B.n383 B.n60 163.367
R737 B.n384 B.n383 163.367
R738 B.n385 B.n384 163.367
R739 B.n385 B.n58 163.367
R740 B.n389 B.n58 163.367
R741 B.n390 B.n389 163.367
R742 B.n391 B.n390 163.367
R743 B.n391 B.n56 163.367
R744 B.n395 B.n56 163.367
R745 B.n396 B.n395 163.367
R746 B.n397 B.n396 163.367
R747 B.n397 B.n54 163.367
R748 B.n401 B.n54 163.367
R749 B.n402 B.n401 163.367
R750 B.n403 B.n402 163.367
R751 B.n403 B.n52 163.367
R752 B.n407 B.n52 163.367
R753 B.n408 B.n407 163.367
R754 B.n409 B.n408 163.367
R755 B.n409 B.n50 163.367
R756 B.n413 B.n50 163.367
R757 B.n414 B.n413 163.367
R758 B.n469 B.n468 163.367
R759 B.n468 B.n27 163.367
R760 B.n464 B.n27 163.367
R761 B.n464 B.n463 163.367
R762 B.n463 B.n462 163.367
R763 B.n462 B.n29 163.367
R764 B.n458 B.n29 163.367
R765 B.n458 B.n457 163.367
R766 B.n457 B.n456 163.367
R767 B.n456 B.n31 163.367
R768 B.n452 B.n31 163.367
R769 B.n452 B.n451 163.367
R770 B.n451 B.n450 163.367
R771 B.n450 B.n33 163.367
R772 B.n446 B.n33 163.367
R773 B.n446 B.n445 163.367
R774 B.n445 B.n444 163.367
R775 B.n444 B.n38 163.367
R776 B.n440 B.n38 163.367
R777 B.n440 B.n439 163.367
R778 B.n439 B.n438 163.367
R779 B.n438 B.n40 163.367
R780 B.n433 B.n40 163.367
R781 B.n433 B.n432 163.367
R782 B.n432 B.n431 163.367
R783 B.n431 B.n44 163.367
R784 B.n427 B.n44 163.367
R785 B.n427 B.n426 163.367
R786 B.n426 B.n425 163.367
R787 B.n425 B.n46 163.367
R788 B.n421 B.n46 163.367
R789 B.n421 B.n420 163.367
R790 B.n420 B.n419 163.367
R791 B.n419 B.n48 163.367
R792 B.n415 B.n48 163.367
R793 B.n249 B.n106 59.5399
R794 B.n113 B.n112 59.5399
R795 B.n36 B.n35 59.5399
R796 B.n435 B.n42 59.5399
R797 B.n106 B.n105 52.5581
R798 B.n112 B.n111 52.5581
R799 B.n35 B.n34 52.5581
R800 B.n42 B.n41 52.5581
R801 B.n471 B.n26 32.3127
R802 B.n416 B.n49 32.3127
R803 B.n268 B.n97 32.3127
R804 B.n214 B.n213 32.3127
R805 B B.n543 18.0485
R806 B.n467 B.n26 10.6151
R807 B.n467 B.n466 10.6151
R808 B.n466 B.n465 10.6151
R809 B.n465 B.n28 10.6151
R810 B.n461 B.n28 10.6151
R811 B.n461 B.n460 10.6151
R812 B.n460 B.n459 10.6151
R813 B.n459 B.n30 10.6151
R814 B.n455 B.n30 10.6151
R815 B.n455 B.n454 10.6151
R816 B.n454 B.n453 10.6151
R817 B.n453 B.n32 10.6151
R818 B.n449 B.n448 10.6151
R819 B.n448 B.n447 10.6151
R820 B.n447 B.n37 10.6151
R821 B.n443 B.n37 10.6151
R822 B.n443 B.n442 10.6151
R823 B.n442 B.n441 10.6151
R824 B.n441 B.n39 10.6151
R825 B.n437 B.n39 10.6151
R826 B.n437 B.n436 10.6151
R827 B.n434 B.n43 10.6151
R828 B.n430 B.n43 10.6151
R829 B.n430 B.n429 10.6151
R830 B.n429 B.n428 10.6151
R831 B.n428 B.n45 10.6151
R832 B.n424 B.n45 10.6151
R833 B.n424 B.n423 10.6151
R834 B.n423 B.n422 10.6151
R835 B.n422 B.n47 10.6151
R836 B.n418 B.n47 10.6151
R837 B.n418 B.n417 10.6151
R838 B.n417 B.n416 10.6151
R839 B.n272 B.n97 10.6151
R840 B.n273 B.n272 10.6151
R841 B.n274 B.n273 10.6151
R842 B.n274 B.n95 10.6151
R843 B.n278 B.n95 10.6151
R844 B.n279 B.n278 10.6151
R845 B.n280 B.n279 10.6151
R846 B.n280 B.n93 10.6151
R847 B.n284 B.n93 10.6151
R848 B.n285 B.n284 10.6151
R849 B.n286 B.n285 10.6151
R850 B.n286 B.n91 10.6151
R851 B.n290 B.n91 10.6151
R852 B.n291 B.n290 10.6151
R853 B.n292 B.n291 10.6151
R854 B.n292 B.n89 10.6151
R855 B.n296 B.n89 10.6151
R856 B.n297 B.n296 10.6151
R857 B.n298 B.n297 10.6151
R858 B.n298 B.n87 10.6151
R859 B.n302 B.n87 10.6151
R860 B.n303 B.n302 10.6151
R861 B.n304 B.n303 10.6151
R862 B.n304 B.n85 10.6151
R863 B.n308 B.n85 10.6151
R864 B.n309 B.n308 10.6151
R865 B.n310 B.n309 10.6151
R866 B.n310 B.n83 10.6151
R867 B.n314 B.n83 10.6151
R868 B.n315 B.n314 10.6151
R869 B.n316 B.n315 10.6151
R870 B.n316 B.n81 10.6151
R871 B.n320 B.n81 10.6151
R872 B.n321 B.n320 10.6151
R873 B.n322 B.n321 10.6151
R874 B.n322 B.n79 10.6151
R875 B.n326 B.n79 10.6151
R876 B.n327 B.n326 10.6151
R877 B.n328 B.n327 10.6151
R878 B.n328 B.n77 10.6151
R879 B.n332 B.n77 10.6151
R880 B.n333 B.n332 10.6151
R881 B.n334 B.n333 10.6151
R882 B.n334 B.n75 10.6151
R883 B.n338 B.n75 10.6151
R884 B.n339 B.n338 10.6151
R885 B.n340 B.n339 10.6151
R886 B.n340 B.n73 10.6151
R887 B.n344 B.n73 10.6151
R888 B.n345 B.n344 10.6151
R889 B.n346 B.n345 10.6151
R890 B.n346 B.n71 10.6151
R891 B.n350 B.n71 10.6151
R892 B.n351 B.n350 10.6151
R893 B.n352 B.n351 10.6151
R894 B.n352 B.n69 10.6151
R895 B.n356 B.n69 10.6151
R896 B.n357 B.n356 10.6151
R897 B.n358 B.n357 10.6151
R898 B.n358 B.n67 10.6151
R899 B.n362 B.n67 10.6151
R900 B.n363 B.n362 10.6151
R901 B.n364 B.n363 10.6151
R902 B.n364 B.n65 10.6151
R903 B.n368 B.n65 10.6151
R904 B.n369 B.n368 10.6151
R905 B.n370 B.n369 10.6151
R906 B.n370 B.n63 10.6151
R907 B.n374 B.n63 10.6151
R908 B.n375 B.n374 10.6151
R909 B.n376 B.n375 10.6151
R910 B.n376 B.n61 10.6151
R911 B.n380 B.n61 10.6151
R912 B.n381 B.n380 10.6151
R913 B.n382 B.n381 10.6151
R914 B.n382 B.n59 10.6151
R915 B.n386 B.n59 10.6151
R916 B.n387 B.n386 10.6151
R917 B.n388 B.n387 10.6151
R918 B.n388 B.n57 10.6151
R919 B.n392 B.n57 10.6151
R920 B.n393 B.n392 10.6151
R921 B.n394 B.n393 10.6151
R922 B.n394 B.n55 10.6151
R923 B.n398 B.n55 10.6151
R924 B.n399 B.n398 10.6151
R925 B.n400 B.n399 10.6151
R926 B.n400 B.n53 10.6151
R927 B.n404 B.n53 10.6151
R928 B.n405 B.n404 10.6151
R929 B.n406 B.n405 10.6151
R930 B.n406 B.n51 10.6151
R931 B.n410 B.n51 10.6151
R932 B.n411 B.n410 10.6151
R933 B.n412 B.n411 10.6151
R934 B.n412 B.n49 10.6151
R935 B.n214 B.n119 10.6151
R936 B.n218 B.n119 10.6151
R937 B.n219 B.n218 10.6151
R938 B.n220 B.n219 10.6151
R939 B.n220 B.n117 10.6151
R940 B.n224 B.n117 10.6151
R941 B.n225 B.n224 10.6151
R942 B.n226 B.n225 10.6151
R943 B.n226 B.n115 10.6151
R944 B.n230 B.n115 10.6151
R945 B.n231 B.n230 10.6151
R946 B.n232 B.n231 10.6151
R947 B.n236 B.n235 10.6151
R948 B.n237 B.n236 10.6151
R949 B.n237 B.n109 10.6151
R950 B.n241 B.n109 10.6151
R951 B.n242 B.n241 10.6151
R952 B.n243 B.n242 10.6151
R953 B.n243 B.n107 10.6151
R954 B.n247 B.n107 10.6151
R955 B.n248 B.n247 10.6151
R956 B.n250 B.n103 10.6151
R957 B.n254 B.n103 10.6151
R958 B.n255 B.n254 10.6151
R959 B.n256 B.n255 10.6151
R960 B.n256 B.n101 10.6151
R961 B.n260 B.n101 10.6151
R962 B.n261 B.n260 10.6151
R963 B.n262 B.n261 10.6151
R964 B.n262 B.n99 10.6151
R965 B.n266 B.n99 10.6151
R966 B.n267 B.n266 10.6151
R967 B.n268 B.n267 10.6151
R968 B.n213 B.n212 10.6151
R969 B.n212 B.n121 10.6151
R970 B.n208 B.n121 10.6151
R971 B.n208 B.n207 10.6151
R972 B.n207 B.n206 10.6151
R973 B.n206 B.n123 10.6151
R974 B.n202 B.n123 10.6151
R975 B.n202 B.n201 10.6151
R976 B.n201 B.n200 10.6151
R977 B.n200 B.n125 10.6151
R978 B.n196 B.n125 10.6151
R979 B.n196 B.n195 10.6151
R980 B.n195 B.n194 10.6151
R981 B.n194 B.n127 10.6151
R982 B.n190 B.n127 10.6151
R983 B.n190 B.n189 10.6151
R984 B.n189 B.n188 10.6151
R985 B.n188 B.n129 10.6151
R986 B.n184 B.n129 10.6151
R987 B.n184 B.n183 10.6151
R988 B.n183 B.n182 10.6151
R989 B.n182 B.n131 10.6151
R990 B.n178 B.n131 10.6151
R991 B.n178 B.n177 10.6151
R992 B.n177 B.n176 10.6151
R993 B.n176 B.n133 10.6151
R994 B.n172 B.n133 10.6151
R995 B.n172 B.n171 10.6151
R996 B.n171 B.n170 10.6151
R997 B.n170 B.n135 10.6151
R998 B.n166 B.n135 10.6151
R999 B.n166 B.n165 10.6151
R1000 B.n165 B.n164 10.6151
R1001 B.n164 B.n137 10.6151
R1002 B.n160 B.n137 10.6151
R1003 B.n160 B.n159 10.6151
R1004 B.n159 B.n158 10.6151
R1005 B.n158 B.n139 10.6151
R1006 B.n154 B.n139 10.6151
R1007 B.n154 B.n153 10.6151
R1008 B.n153 B.n152 10.6151
R1009 B.n152 B.n141 10.6151
R1010 B.n148 B.n141 10.6151
R1011 B.n148 B.n147 10.6151
R1012 B.n147 B.n146 10.6151
R1013 B.n146 B.n143 10.6151
R1014 B.n143 B.n0 10.6151
R1015 B.n539 B.n1 10.6151
R1016 B.n539 B.n538 10.6151
R1017 B.n538 B.n537 10.6151
R1018 B.n537 B.n4 10.6151
R1019 B.n533 B.n4 10.6151
R1020 B.n533 B.n532 10.6151
R1021 B.n532 B.n531 10.6151
R1022 B.n531 B.n6 10.6151
R1023 B.n527 B.n6 10.6151
R1024 B.n527 B.n526 10.6151
R1025 B.n526 B.n525 10.6151
R1026 B.n525 B.n8 10.6151
R1027 B.n521 B.n8 10.6151
R1028 B.n521 B.n520 10.6151
R1029 B.n520 B.n519 10.6151
R1030 B.n519 B.n10 10.6151
R1031 B.n515 B.n10 10.6151
R1032 B.n515 B.n514 10.6151
R1033 B.n514 B.n513 10.6151
R1034 B.n513 B.n12 10.6151
R1035 B.n509 B.n12 10.6151
R1036 B.n509 B.n508 10.6151
R1037 B.n508 B.n507 10.6151
R1038 B.n507 B.n14 10.6151
R1039 B.n503 B.n14 10.6151
R1040 B.n503 B.n502 10.6151
R1041 B.n502 B.n501 10.6151
R1042 B.n501 B.n16 10.6151
R1043 B.n497 B.n16 10.6151
R1044 B.n497 B.n496 10.6151
R1045 B.n496 B.n495 10.6151
R1046 B.n495 B.n18 10.6151
R1047 B.n491 B.n18 10.6151
R1048 B.n491 B.n490 10.6151
R1049 B.n490 B.n489 10.6151
R1050 B.n489 B.n20 10.6151
R1051 B.n485 B.n20 10.6151
R1052 B.n485 B.n484 10.6151
R1053 B.n484 B.n483 10.6151
R1054 B.n483 B.n22 10.6151
R1055 B.n479 B.n22 10.6151
R1056 B.n479 B.n478 10.6151
R1057 B.n478 B.n477 10.6151
R1058 B.n477 B.n24 10.6151
R1059 B.n473 B.n24 10.6151
R1060 B.n473 B.n472 10.6151
R1061 B.n472 B.n471 10.6151
R1062 B.n36 B.n32 9.36635
R1063 B.n435 B.n434 9.36635
R1064 B.n232 B.n113 9.36635
R1065 B.n250 B.n249 9.36635
R1066 B.n543 B.n0 2.81026
R1067 B.n543 B.n1 2.81026
R1068 B.n449 B.n36 1.24928
R1069 B.n436 B.n435 1.24928
R1070 B.n235 B.n113 1.24928
R1071 B.n249 B.n248 1.24928
C0 VDD1 B 1.32268f
C1 VP w_n3680_n1438# 7.72458f
C2 VN VP 5.61229f
C3 VDD1 VP 2.38417f
C4 VDD2 VTAIL 4.69712f
C5 VDD2 w_n3680_n1438# 1.71981f
C6 w_n3680_n1438# VTAIL 1.97257f
C7 VN VDD2 2.04074f
C8 VN VTAIL 3.02216f
C9 VDD1 VDD2 1.66038f
C10 VDD1 VTAIL 4.64418f
C11 VN w_n3680_n1438# 7.251f
C12 VP B 1.861f
C13 VDD1 w_n3680_n1438# 1.61499f
C14 VDD1 VN 0.156452f
C15 VDD2 B 1.41207f
C16 B VTAIL 1.67838f
C17 B w_n3680_n1438# 7.10991f
C18 VN B 1.06302f
C19 VP VDD2 0.502358f
C20 VP VTAIL 3.03626f
C21 VDD2 VSUBS 1.324207f
C22 VDD1 VSUBS 1.948145f
C23 VTAIL VSUBS 0.523595f
C24 VN VSUBS 6.41461f
C25 VP VSUBS 2.781084f
C26 B VSUBS 3.706382f
C27 w_n3680_n1438# VSUBS 67.344f
C28 B.n0 VSUBS 0.005207f
C29 B.n1 VSUBS 0.005207f
C30 B.n2 VSUBS 0.008235f
C31 B.n3 VSUBS 0.008235f
C32 B.n4 VSUBS 0.008235f
C33 B.n5 VSUBS 0.008235f
C34 B.n6 VSUBS 0.008235f
C35 B.n7 VSUBS 0.008235f
C36 B.n8 VSUBS 0.008235f
C37 B.n9 VSUBS 0.008235f
C38 B.n10 VSUBS 0.008235f
C39 B.n11 VSUBS 0.008235f
C40 B.n12 VSUBS 0.008235f
C41 B.n13 VSUBS 0.008235f
C42 B.n14 VSUBS 0.008235f
C43 B.n15 VSUBS 0.008235f
C44 B.n16 VSUBS 0.008235f
C45 B.n17 VSUBS 0.008235f
C46 B.n18 VSUBS 0.008235f
C47 B.n19 VSUBS 0.008235f
C48 B.n20 VSUBS 0.008235f
C49 B.n21 VSUBS 0.008235f
C50 B.n22 VSUBS 0.008235f
C51 B.n23 VSUBS 0.008235f
C52 B.n24 VSUBS 0.008235f
C53 B.n25 VSUBS 0.008235f
C54 B.n26 VSUBS 0.019554f
C55 B.n27 VSUBS 0.008235f
C56 B.n28 VSUBS 0.008235f
C57 B.n29 VSUBS 0.008235f
C58 B.n30 VSUBS 0.008235f
C59 B.n31 VSUBS 0.008235f
C60 B.n32 VSUBS 0.007751f
C61 B.n33 VSUBS 0.008235f
C62 B.t11 VSUBS 0.061707f
C63 B.t10 VSUBS 0.075471f
C64 B.t9 VSUBS 0.321947f
C65 B.n34 VSUBS 0.087085f
C66 B.n35 VSUBS 0.07129f
C67 B.n36 VSUBS 0.019079f
C68 B.n37 VSUBS 0.008235f
C69 B.n38 VSUBS 0.008235f
C70 B.n39 VSUBS 0.008235f
C71 B.n40 VSUBS 0.008235f
C72 B.t5 VSUBS 0.061707f
C73 B.t4 VSUBS 0.075471f
C74 B.t3 VSUBS 0.321947f
C75 B.n41 VSUBS 0.087085f
C76 B.n42 VSUBS 0.07129f
C77 B.n43 VSUBS 0.008235f
C78 B.n44 VSUBS 0.008235f
C79 B.n45 VSUBS 0.008235f
C80 B.n46 VSUBS 0.008235f
C81 B.n47 VSUBS 0.008235f
C82 B.n48 VSUBS 0.008235f
C83 B.n49 VSUBS 0.019698f
C84 B.n50 VSUBS 0.008235f
C85 B.n51 VSUBS 0.008235f
C86 B.n52 VSUBS 0.008235f
C87 B.n53 VSUBS 0.008235f
C88 B.n54 VSUBS 0.008235f
C89 B.n55 VSUBS 0.008235f
C90 B.n56 VSUBS 0.008235f
C91 B.n57 VSUBS 0.008235f
C92 B.n58 VSUBS 0.008235f
C93 B.n59 VSUBS 0.008235f
C94 B.n60 VSUBS 0.008235f
C95 B.n61 VSUBS 0.008235f
C96 B.n62 VSUBS 0.008235f
C97 B.n63 VSUBS 0.008235f
C98 B.n64 VSUBS 0.008235f
C99 B.n65 VSUBS 0.008235f
C100 B.n66 VSUBS 0.008235f
C101 B.n67 VSUBS 0.008235f
C102 B.n68 VSUBS 0.008235f
C103 B.n69 VSUBS 0.008235f
C104 B.n70 VSUBS 0.008235f
C105 B.n71 VSUBS 0.008235f
C106 B.n72 VSUBS 0.008235f
C107 B.n73 VSUBS 0.008235f
C108 B.n74 VSUBS 0.008235f
C109 B.n75 VSUBS 0.008235f
C110 B.n76 VSUBS 0.008235f
C111 B.n77 VSUBS 0.008235f
C112 B.n78 VSUBS 0.008235f
C113 B.n79 VSUBS 0.008235f
C114 B.n80 VSUBS 0.008235f
C115 B.n81 VSUBS 0.008235f
C116 B.n82 VSUBS 0.008235f
C117 B.n83 VSUBS 0.008235f
C118 B.n84 VSUBS 0.008235f
C119 B.n85 VSUBS 0.008235f
C120 B.n86 VSUBS 0.008235f
C121 B.n87 VSUBS 0.008235f
C122 B.n88 VSUBS 0.008235f
C123 B.n89 VSUBS 0.008235f
C124 B.n90 VSUBS 0.008235f
C125 B.n91 VSUBS 0.008235f
C126 B.n92 VSUBS 0.008235f
C127 B.n93 VSUBS 0.008235f
C128 B.n94 VSUBS 0.008235f
C129 B.n95 VSUBS 0.008235f
C130 B.n96 VSUBS 0.008235f
C131 B.n97 VSUBS 0.018714f
C132 B.n98 VSUBS 0.008235f
C133 B.n99 VSUBS 0.008235f
C134 B.n100 VSUBS 0.008235f
C135 B.n101 VSUBS 0.008235f
C136 B.n102 VSUBS 0.008235f
C137 B.n103 VSUBS 0.008235f
C138 B.n104 VSUBS 0.008235f
C139 B.t1 VSUBS 0.061707f
C140 B.t2 VSUBS 0.075471f
C141 B.t0 VSUBS 0.321947f
C142 B.n105 VSUBS 0.087085f
C143 B.n106 VSUBS 0.07129f
C144 B.n107 VSUBS 0.008235f
C145 B.n108 VSUBS 0.008235f
C146 B.n109 VSUBS 0.008235f
C147 B.n110 VSUBS 0.008235f
C148 B.t7 VSUBS 0.061707f
C149 B.t8 VSUBS 0.075471f
C150 B.t6 VSUBS 0.321947f
C151 B.n111 VSUBS 0.087085f
C152 B.n112 VSUBS 0.07129f
C153 B.n113 VSUBS 0.019079f
C154 B.n114 VSUBS 0.008235f
C155 B.n115 VSUBS 0.008235f
C156 B.n116 VSUBS 0.008235f
C157 B.n117 VSUBS 0.008235f
C158 B.n118 VSUBS 0.008235f
C159 B.n119 VSUBS 0.008235f
C160 B.n120 VSUBS 0.018714f
C161 B.n121 VSUBS 0.008235f
C162 B.n122 VSUBS 0.008235f
C163 B.n123 VSUBS 0.008235f
C164 B.n124 VSUBS 0.008235f
C165 B.n125 VSUBS 0.008235f
C166 B.n126 VSUBS 0.008235f
C167 B.n127 VSUBS 0.008235f
C168 B.n128 VSUBS 0.008235f
C169 B.n129 VSUBS 0.008235f
C170 B.n130 VSUBS 0.008235f
C171 B.n131 VSUBS 0.008235f
C172 B.n132 VSUBS 0.008235f
C173 B.n133 VSUBS 0.008235f
C174 B.n134 VSUBS 0.008235f
C175 B.n135 VSUBS 0.008235f
C176 B.n136 VSUBS 0.008235f
C177 B.n137 VSUBS 0.008235f
C178 B.n138 VSUBS 0.008235f
C179 B.n139 VSUBS 0.008235f
C180 B.n140 VSUBS 0.008235f
C181 B.n141 VSUBS 0.008235f
C182 B.n142 VSUBS 0.008235f
C183 B.n143 VSUBS 0.008235f
C184 B.n144 VSUBS 0.008235f
C185 B.n145 VSUBS 0.008235f
C186 B.n146 VSUBS 0.008235f
C187 B.n147 VSUBS 0.008235f
C188 B.n148 VSUBS 0.008235f
C189 B.n149 VSUBS 0.008235f
C190 B.n150 VSUBS 0.008235f
C191 B.n151 VSUBS 0.008235f
C192 B.n152 VSUBS 0.008235f
C193 B.n153 VSUBS 0.008235f
C194 B.n154 VSUBS 0.008235f
C195 B.n155 VSUBS 0.008235f
C196 B.n156 VSUBS 0.008235f
C197 B.n157 VSUBS 0.008235f
C198 B.n158 VSUBS 0.008235f
C199 B.n159 VSUBS 0.008235f
C200 B.n160 VSUBS 0.008235f
C201 B.n161 VSUBS 0.008235f
C202 B.n162 VSUBS 0.008235f
C203 B.n163 VSUBS 0.008235f
C204 B.n164 VSUBS 0.008235f
C205 B.n165 VSUBS 0.008235f
C206 B.n166 VSUBS 0.008235f
C207 B.n167 VSUBS 0.008235f
C208 B.n168 VSUBS 0.008235f
C209 B.n169 VSUBS 0.008235f
C210 B.n170 VSUBS 0.008235f
C211 B.n171 VSUBS 0.008235f
C212 B.n172 VSUBS 0.008235f
C213 B.n173 VSUBS 0.008235f
C214 B.n174 VSUBS 0.008235f
C215 B.n175 VSUBS 0.008235f
C216 B.n176 VSUBS 0.008235f
C217 B.n177 VSUBS 0.008235f
C218 B.n178 VSUBS 0.008235f
C219 B.n179 VSUBS 0.008235f
C220 B.n180 VSUBS 0.008235f
C221 B.n181 VSUBS 0.008235f
C222 B.n182 VSUBS 0.008235f
C223 B.n183 VSUBS 0.008235f
C224 B.n184 VSUBS 0.008235f
C225 B.n185 VSUBS 0.008235f
C226 B.n186 VSUBS 0.008235f
C227 B.n187 VSUBS 0.008235f
C228 B.n188 VSUBS 0.008235f
C229 B.n189 VSUBS 0.008235f
C230 B.n190 VSUBS 0.008235f
C231 B.n191 VSUBS 0.008235f
C232 B.n192 VSUBS 0.008235f
C233 B.n193 VSUBS 0.008235f
C234 B.n194 VSUBS 0.008235f
C235 B.n195 VSUBS 0.008235f
C236 B.n196 VSUBS 0.008235f
C237 B.n197 VSUBS 0.008235f
C238 B.n198 VSUBS 0.008235f
C239 B.n199 VSUBS 0.008235f
C240 B.n200 VSUBS 0.008235f
C241 B.n201 VSUBS 0.008235f
C242 B.n202 VSUBS 0.008235f
C243 B.n203 VSUBS 0.008235f
C244 B.n204 VSUBS 0.008235f
C245 B.n205 VSUBS 0.008235f
C246 B.n206 VSUBS 0.008235f
C247 B.n207 VSUBS 0.008235f
C248 B.n208 VSUBS 0.008235f
C249 B.n209 VSUBS 0.008235f
C250 B.n210 VSUBS 0.008235f
C251 B.n211 VSUBS 0.008235f
C252 B.n212 VSUBS 0.008235f
C253 B.n213 VSUBS 0.018714f
C254 B.n214 VSUBS 0.019554f
C255 B.n215 VSUBS 0.019554f
C256 B.n216 VSUBS 0.008235f
C257 B.n217 VSUBS 0.008235f
C258 B.n218 VSUBS 0.008235f
C259 B.n219 VSUBS 0.008235f
C260 B.n220 VSUBS 0.008235f
C261 B.n221 VSUBS 0.008235f
C262 B.n222 VSUBS 0.008235f
C263 B.n223 VSUBS 0.008235f
C264 B.n224 VSUBS 0.008235f
C265 B.n225 VSUBS 0.008235f
C266 B.n226 VSUBS 0.008235f
C267 B.n227 VSUBS 0.008235f
C268 B.n228 VSUBS 0.008235f
C269 B.n229 VSUBS 0.008235f
C270 B.n230 VSUBS 0.008235f
C271 B.n231 VSUBS 0.008235f
C272 B.n232 VSUBS 0.007751f
C273 B.n233 VSUBS 0.008235f
C274 B.n234 VSUBS 0.008235f
C275 B.n235 VSUBS 0.004602f
C276 B.n236 VSUBS 0.008235f
C277 B.n237 VSUBS 0.008235f
C278 B.n238 VSUBS 0.008235f
C279 B.n239 VSUBS 0.008235f
C280 B.n240 VSUBS 0.008235f
C281 B.n241 VSUBS 0.008235f
C282 B.n242 VSUBS 0.008235f
C283 B.n243 VSUBS 0.008235f
C284 B.n244 VSUBS 0.008235f
C285 B.n245 VSUBS 0.008235f
C286 B.n246 VSUBS 0.008235f
C287 B.n247 VSUBS 0.008235f
C288 B.n248 VSUBS 0.004602f
C289 B.n249 VSUBS 0.019079f
C290 B.n250 VSUBS 0.007751f
C291 B.n251 VSUBS 0.008235f
C292 B.n252 VSUBS 0.008235f
C293 B.n253 VSUBS 0.008235f
C294 B.n254 VSUBS 0.008235f
C295 B.n255 VSUBS 0.008235f
C296 B.n256 VSUBS 0.008235f
C297 B.n257 VSUBS 0.008235f
C298 B.n258 VSUBS 0.008235f
C299 B.n259 VSUBS 0.008235f
C300 B.n260 VSUBS 0.008235f
C301 B.n261 VSUBS 0.008235f
C302 B.n262 VSUBS 0.008235f
C303 B.n263 VSUBS 0.008235f
C304 B.n264 VSUBS 0.008235f
C305 B.n265 VSUBS 0.008235f
C306 B.n266 VSUBS 0.008235f
C307 B.n267 VSUBS 0.008235f
C308 B.n268 VSUBS 0.019554f
C309 B.n269 VSUBS 0.019554f
C310 B.n270 VSUBS 0.018714f
C311 B.n271 VSUBS 0.008235f
C312 B.n272 VSUBS 0.008235f
C313 B.n273 VSUBS 0.008235f
C314 B.n274 VSUBS 0.008235f
C315 B.n275 VSUBS 0.008235f
C316 B.n276 VSUBS 0.008235f
C317 B.n277 VSUBS 0.008235f
C318 B.n278 VSUBS 0.008235f
C319 B.n279 VSUBS 0.008235f
C320 B.n280 VSUBS 0.008235f
C321 B.n281 VSUBS 0.008235f
C322 B.n282 VSUBS 0.008235f
C323 B.n283 VSUBS 0.008235f
C324 B.n284 VSUBS 0.008235f
C325 B.n285 VSUBS 0.008235f
C326 B.n286 VSUBS 0.008235f
C327 B.n287 VSUBS 0.008235f
C328 B.n288 VSUBS 0.008235f
C329 B.n289 VSUBS 0.008235f
C330 B.n290 VSUBS 0.008235f
C331 B.n291 VSUBS 0.008235f
C332 B.n292 VSUBS 0.008235f
C333 B.n293 VSUBS 0.008235f
C334 B.n294 VSUBS 0.008235f
C335 B.n295 VSUBS 0.008235f
C336 B.n296 VSUBS 0.008235f
C337 B.n297 VSUBS 0.008235f
C338 B.n298 VSUBS 0.008235f
C339 B.n299 VSUBS 0.008235f
C340 B.n300 VSUBS 0.008235f
C341 B.n301 VSUBS 0.008235f
C342 B.n302 VSUBS 0.008235f
C343 B.n303 VSUBS 0.008235f
C344 B.n304 VSUBS 0.008235f
C345 B.n305 VSUBS 0.008235f
C346 B.n306 VSUBS 0.008235f
C347 B.n307 VSUBS 0.008235f
C348 B.n308 VSUBS 0.008235f
C349 B.n309 VSUBS 0.008235f
C350 B.n310 VSUBS 0.008235f
C351 B.n311 VSUBS 0.008235f
C352 B.n312 VSUBS 0.008235f
C353 B.n313 VSUBS 0.008235f
C354 B.n314 VSUBS 0.008235f
C355 B.n315 VSUBS 0.008235f
C356 B.n316 VSUBS 0.008235f
C357 B.n317 VSUBS 0.008235f
C358 B.n318 VSUBS 0.008235f
C359 B.n319 VSUBS 0.008235f
C360 B.n320 VSUBS 0.008235f
C361 B.n321 VSUBS 0.008235f
C362 B.n322 VSUBS 0.008235f
C363 B.n323 VSUBS 0.008235f
C364 B.n324 VSUBS 0.008235f
C365 B.n325 VSUBS 0.008235f
C366 B.n326 VSUBS 0.008235f
C367 B.n327 VSUBS 0.008235f
C368 B.n328 VSUBS 0.008235f
C369 B.n329 VSUBS 0.008235f
C370 B.n330 VSUBS 0.008235f
C371 B.n331 VSUBS 0.008235f
C372 B.n332 VSUBS 0.008235f
C373 B.n333 VSUBS 0.008235f
C374 B.n334 VSUBS 0.008235f
C375 B.n335 VSUBS 0.008235f
C376 B.n336 VSUBS 0.008235f
C377 B.n337 VSUBS 0.008235f
C378 B.n338 VSUBS 0.008235f
C379 B.n339 VSUBS 0.008235f
C380 B.n340 VSUBS 0.008235f
C381 B.n341 VSUBS 0.008235f
C382 B.n342 VSUBS 0.008235f
C383 B.n343 VSUBS 0.008235f
C384 B.n344 VSUBS 0.008235f
C385 B.n345 VSUBS 0.008235f
C386 B.n346 VSUBS 0.008235f
C387 B.n347 VSUBS 0.008235f
C388 B.n348 VSUBS 0.008235f
C389 B.n349 VSUBS 0.008235f
C390 B.n350 VSUBS 0.008235f
C391 B.n351 VSUBS 0.008235f
C392 B.n352 VSUBS 0.008235f
C393 B.n353 VSUBS 0.008235f
C394 B.n354 VSUBS 0.008235f
C395 B.n355 VSUBS 0.008235f
C396 B.n356 VSUBS 0.008235f
C397 B.n357 VSUBS 0.008235f
C398 B.n358 VSUBS 0.008235f
C399 B.n359 VSUBS 0.008235f
C400 B.n360 VSUBS 0.008235f
C401 B.n361 VSUBS 0.008235f
C402 B.n362 VSUBS 0.008235f
C403 B.n363 VSUBS 0.008235f
C404 B.n364 VSUBS 0.008235f
C405 B.n365 VSUBS 0.008235f
C406 B.n366 VSUBS 0.008235f
C407 B.n367 VSUBS 0.008235f
C408 B.n368 VSUBS 0.008235f
C409 B.n369 VSUBS 0.008235f
C410 B.n370 VSUBS 0.008235f
C411 B.n371 VSUBS 0.008235f
C412 B.n372 VSUBS 0.008235f
C413 B.n373 VSUBS 0.008235f
C414 B.n374 VSUBS 0.008235f
C415 B.n375 VSUBS 0.008235f
C416 B.n376 VSUBS 0.008235f
C417 B.n377 VSUBS 0.008235f
C418 B.n378 VSUBS 0.008235f
C419 B.n379 VSUBS 0.008235f
C420 B.n380 VSUBS 0.008235f
C421 B.n381 VSUBS 0.008235f
C422 B.n382 VSUBS 0.008235f
C423 B.n383 VSUBS 0.008235f
C424 B.n384 VSUBS 0.008235f
C425 B.n385 VSUBS 0.008235f
C426 B.n386 VSUBS 0.008235f
C427 B.n387 VSUBS 0.008235f
C428 B.n388 VSUBS 0.008235f
C429 B.n389 VSUBS 0.008235f
C430 B.n390 VSUBS 0.008235f
C431 B.n391 VSUBS 0.008235f
C432 B.n392 VSUBS 0.008235f
C433 B.n393 VSUBS 0.008235f
C434 B.n394 VSUBS 0.008235f
C435 B.n395 VSUBS 0.008235f
C436 B.n396 VSUBS 0.008235f
C437 B.n397 VSUBS 0.008235f
C438 B.n398 VSUBS 0.008235f
C439 B.n399 VSUBS 0.008235f
C440 B.n400 VSUBS 0.008235f
C441 B.n401 VSUBS 0.008235f
C442 B.n402 VSUBS 0.008235f
C443 B.n403 VSUBS 0.008235f
C444 B.n404 VSUBS 0.008235f
C445 B.n405 VSUBS 0.008235f
C446 B.n406 VSUBS 0.008235f
C447 B.n407 VSUBS 0.008235f
C448 B.n408 VSUBS 0.008235f
C449 B.n409 VSUBS 0.008235f
C450 B.n410 VSUBS 0.008235f
C451 B.n411 VSUBS 0.008235f
C452 B.n412 VSUBS 0.008235f
C453 B.n413 VSUBS 0.008235f
C454 B.n414 VSUBS 0.018714f
C455 B.n415 VSUBS 0.019554f
C456 B.n416 VSUBS 0.01857f
C457 B.n417 VSUBS 0.008235f
C458 B.n418 VSUBS 0.008235f
C459 B.n419 VSUBS 0.008235f
C460 B.n420 VSUBS 0.008235f
C461 B.n421 VSUBS 0.008235f
C462 B.n422 VSUBS 0.008235f
C463 B.n423 VSUBS 0.008235f
C464 B.n424 VSUBS 0.008235f
C465 B.n425 VSUBS 0.008235f
C466 B.n426 VSUBS 0.008235f
C467 B.n427 VSUBS 0.008235f
C468 B.n428 VSUBS 0.008235f
C469 B.n429 VSUBS 0.008235f
C470 B.n430 VSUBS 0.008235f
C471 B.n431 VSUBS 0.008235f
C472 B.n432 VSUBS 0.008235f
C473 B.n433 VSUBS 0.008235f
C474 B.n434 VSUBS 0.007751f
C475 B.n435 VSUBS 0.019079f
C476 B.n436 VSUBS 0.004602f
C477 B.n437 VSUBS 0.008235f
C478 B.n438 VSUBS 0.008235f
C479 B.n439 VSUBS 0.008235f
C480 B.n440 VSUBS 0.008235f
C481 B.n441 VSUBS 0.008235f
C482 B.n442 VSUBS 0.008235f
C483 B.n443 VSUBS 0.008235f
C484 B.n444 VSUBS 0.008235f
C485 B.n445 VSUBS 0.008235f
C486 B.n446 VSUBS 0.008235f
C487 B.n447 VSUBS 0.008235f
C488 B.n448 VSUBS 0.008235f
C489 B.n449 VSUBS 0.004602f
C490 B.n450 VSUBS 0.008235f
C491 B.n451 VSUBS 0.008235f
C492 B.n452 VSUBS 0.008235f
C493 B.n453 VSUBS 0.008235f
C494 B.n454 VSUBS 0.008235f
C495 B.n455 VSUBS 0.008235f
C496 B.n456 VSUBS 0.008235f
C497 B.n457 VSUBS 0.008235f
C498 B.n458 VSUBS 0.008235f
C499 B.n459 VSUBS 0.008235f
C500 B.n460 VSUBS 0.008235f
C501 B.n461 VSUBS 0.008235f
C502 B.n462 VSUBS 0.008235f
C503 B.n463 VSUBS 0.008235f
C504 B.n464 VSUBS 0.008235f
C505 B.n465 VSUBS 0.008235f
C506 B.n466 VSUBS 0.008235f
C507 B.n467 VSUBS 0.008235f
C508 B.n468 VSUBS 0.008235f
C509 B.n469 VSUBS 0.019554f
C510 B.n470 VSUBS 0.018714f
C511 B.n471 VSUBS 0.018714f
C512 B.n472 VSUBS 0.008235f
C513 B.n473 VSUBS 0.008235f
C514 B.n474 VSUBS 0.008235f
C515 B.n475 VSUBS 0.008235f
C516 B.n476 VSUBS 0.008235f
C517 B.n477 VSUBS 0.008235f
C518 B.n478 VSUBS 0.008235f
C519 B.n479 VSUBS 0.008235f
C520 B.n480 VSUBS 0.008235f
C521 B.n481 VSUBS 0.008235f
C522 B.n482 VSUBS 0.008235f
C523 B.n483 VSUBS 0.008235f
C524 B.n484 VSUBS 0.008235f
C525 B.n485 VSUBS 0.008235f
C526 B.n486 VSUBS 0.008235f
C527 B.n487 VSUBS 0.008235f
C528 B.n488 VSUBS 0.008235f
C529 B.n489 VSUBS 0.008235f
C530 B.n490 VSUBS 0.008235f
C531 B.n491 VSUBS 0.008235f
C532 B.n492 VSUBS 0.008235f
C533 B.n493 VSUBS 0.008235f
C534 B.n494 VSUBS 0.008235f
C535 B.n495 VSUBS 0.008235f
C536 B.n496 VSUBS 0.008235f
C537 B.n497 VSUBS 0.008235f
C538 B.n498 VSUBS 0.008235f
C539 B.n499 VSUBS 0.008235f
C540 B.n500 VSUBS 0.008235f
C541 B.n501 VSUBS 0.008235f
C542 B.n502 VSUBS 0.008235f
C543 B.n503 VSUBS 0.008235f
C544 B.n504 VSUBS 0.008235f
C545 B.n505 VSUBS 0.008235f
C546 B.n506 VSUBS 0.008235f
C547 B.n507 VSUBS 0.008235f
C548 B.n508 VSUBS 0.008235f
C549 B.n509 VSUBS 0.008235f
C550 B.n510 VSUBS 0.008235f
C551 B.n511 VSUBS 0.008235f
C552 B.n512 VSUBS 0.008235f
C553 B.n513 VSUBS 0.008235f
C554 B.n514 VSUBS 0.008235f
C555 B.n515 VSUBS 0.008235f
C556 B.n516 VSUBS 0.008235f
C557 B.n517 VSUBS 0.008235f
C558 B.n518 VSUBS 0.008235f
C559 B.n519 VSUBS 0.008235f
C560 B.n520 VSUBS 0.008235f
C561 B.n521 VSUBS 0.008235f
C562 B.n522 VSUBS 0.008235f
C563 B.n523 VSUBS 0.008235f
C564 B.n524 VSUBS 0.008235f
C565 B.n525 VSUBS 0.008235f
C566 B.n526 VSUBS 0.008235f
C567 B.n527 VSUBS 0.008235f
C568 B.n528 VSUBS 0.008235f
C569 B.n529 VSUBS 0.008235f
C570 B.n530 VSUBS 0.008235f
C571 B.n531 VSUBS 0.008235f
C572 B.n532 VSUBS 0.008235f
C573 B.n533 VSUBS 0.008235f
C574 B.n534 VSUBS 0.008235f
C575 B.n535 VSUBS 0.008235f
C576 B.n536 VSUBS 0.008235f
C577 B.n537 VSUBS 0.008235f
C578 B.n538 VSUBS 0.008235f
C579 B.n539 VSUBS 0.008235f
C580 B.n540 VSUBS 0.008235f
C581 B.n541 VSUBS 0.008235f
C582 B.n542 VSUBS 0.008235f
C583 B.n543 VSUBS 0.018647f
C584 VDD2.t2 VSUBS 0.044741f
C585 VDD2.t1 VSUBS 0.044741f
C586 VDD2.n0 VSUBS 0.204811f
C587 VDD2.t0 VSUBS 0.044741f
C588 VDD2.t5 VSUBS 0.044741f
C589 VDD2.n1 VSUBS 0.204811f
C590 VDD2.n2 VSUBS 2.6553f
C591 VDD2.t6 VSUBS 0.044741f
C592 VDD2.t3 VSUBS 0.044741f
C593 VDD2.n3 VSUBS 0.201178f
C594 VDD2.n4 VSUBS 2.13035f
C595 VDD2.t7 VSUBS 0.044741f
C596 VDD2.t4 VSUBS 0.044741f
C597 VDD2.n5 VSUBS 0.204798f
C598 VN.n0 VSUBS 0.06789f
C599 VN.t2 VSUBS 0.692641f
C600 VN.n1 VSUBS 0.042696f
C601 VN.n2 VSUBS 0.051494f
C602 VN.t7 VSUBS 0.692641f
C603 VN.n3 VSUBS 0.095972f
C604 VN.n4 VSUBS 0.051494f
C605 VN.n5 VSUBS 0.058538f
C606 VN.t5 VSUBS 1.04594f
C607 VN.t6 VSUBS 0.692641f
C608 VN.n6 VSUBS 0.444175f
C609 VN.n7 VSUBS 0.437151f
C610 VN.n8 VSUBS 0.447547f
C611 VN.n9 VSUBS 0.051494f
C612 VN.n10 VSUBS 0.095972f
C613 VN.n11 VSUBS 0.075172f
C614 VN.n12 VSUBS 0.075172f
C615 VN.n13 VSUBS 0.051494f
C616 VN.n14 VSUBS 0.051494f
C617 VN.n15 VSUBS 0.051494f
C618 VN.n16 VSUBS 0.058538f
C619 VN.n17 VSUBS 0.316419f
C620 VN.n18 VSUBS 0.086019f
C621 VN.n19 VSUBS 0.099794f
C622 VN.n20 VSUBS 0.051494f
C623 VN.n21 VSUBS 0.051494f
C624 VN.n22 VSUBS 0.051494f
C625 VN.n23 VSUBS 0.103825f
C626 VN.n24 VSUBS 0.078438f
C627 VN.n25 VSUBS 0.489659f
C628 VN.n26 VSUBS 0.072969f
C629 VN.n27 VSUBS 0.06789f
C630 VN.t1 VSUBS 0.692641f
C631 VN.n28 VSUBS 0.042696f
C632 VN.n29 VSUBS 0.051494f
C633 VN.t4 VSUBS 0.692641f
C634 VN.n30 VSUBS 0.095972f
C635 VN.n31 VSUBS 0.051494f
C636 VN.n32 VSUBS 0.058538f
C637 VN.t3 VSUBS 1.04594f
C638 VN.t0 VSUBS 0.692641f
C639 VN.n33 VSUBS 0.444175f
C640 VN.n34 VSUBS 0.437151f
C641 VN.n35 VSUBS 0.447547f
C642 VN.n36 VSUBS 0.051494f
C643 VN.n37 VSUBS 0.095972f
C644 VN.n38 VSUBS 0.075172f
C645 VN.n39 VSUBS 0.075172f
C646 VN.n40 VSUBS 0.051494f
C647 VN.n41 VSUBS 0.051494f
C648 VN.n42 VSUBS 0.051494f
C649 VN.n43 VSUBS 0.058538f
C650 VN.n44 VSUBS 0.316419f
C651 VN.n45 VSUBS 0.086019f
C652 VN.n46 VSUBS 0.099794f
C653 VN.n47 VSUBS 0.051494f
C654 VN.n48 VSUBS 0.051494f
C655 VN.n49 VSUBS 0.051494f
C656 VN.n50 VSUBS 0.103825f
C657 VN.n51 VSUBS 0.078438f
C658 VN.n52 VSUBS 0.489659f
C659 VN.n53 VSUBS 2.26023f
C660 VDD1.t0 VSUBS 0.046131f
C661 VDD1.t3 VSUBS 0.046131f
C662 VDD1.n0 VSUBS 0.211618f
C663 VDD1.t5 VSUBS 0.046131f
C664 VDD1.t6 VSUBS 0.046131f
C665 VDD1.n1 VSUBS 0.211177f
C666 VDD1.t2 VSUBS 0.046131f
C667 VDD1.t4 VSUBS 0.046131f
C668 VDD1.n2 VSUBS 0.211177f
C669 VDD1.n3 VSUBS 2.78992f
C670 VDD1.t1 VSUBS 0.046131f
C671 VDD1.t7 VSUBS 0.046131f
C672 VDD1.n4 VSUBS 0.207431f
C673 VDD1.n5 VSUBS 2.22692f
C674 VTAIL.t0 VSUBS 0.054777f
C675 VTAIL.t4 VSUBS 0.054777f
C676 VTAIL.n0 VSUBS 0.20922f
C677 VTAIL.n1 VSUBS 0.574536f
C678 VTAIL.t5 VSUBS 0.333701f
C679 VTAIL.n2 VSUBS 0.638573f
C680 VTAIL.t13 VSUBS 0.333701f
C681 VTAIL.n3 VSUBS 0.638573f
C682 VTAIL.t12 VSUBS 0.054777f
C683 VTAIL.t14 VSUBS 0.054777f
C684 VTAIL.n4 VSUBS 0.20922f
C685 VTAIL.n5 VSUBS 0.791053f
C686 VTAIL.t11 VSUBS 0.333701f
C687 VTAIL.n6 VSUBS 1.4092f
C688 VTAIL.t7 VSUBS 0.333702f
C689 VTAIL.n7 VSUBS 1.4092f
C690 VTAIL.t6 VSUBS 0.054777f
C691 VTAIL.t3 VSUBS 0.054777f
C692 VTAIL.n8 VSUBS 0.209222f
C693 VTAIL.n9 VSUBS 0.791052f
C694 VTAIL.t2 VSUBS 0.333702f
C695 VTAIL.n10 VSUBS 0.638572f
C696 VTAIL.t8 VSUBS 0.333702f
C697 VTAIL.n11 VSUBS 0.638572f
C698 VTAIL.t10 VSUBS 0.054777f
C699 VTAIL.t15 VSUBS 0.054777f
C700 VTAIL.n12 VSUBS 0.209222f
C701 VTAIL.n13 VSUBS 0.791052f
C702 VTAIL.t9 VSUBS 0.333702f
C703 VTAIL.n14 VSUBS 1.4092f
C704 VTAIL.t1 VSUBS 0.333701f
C705 VTAIL.n15 VSUBS 1.40367f
C706 VP.n0 VSUBS 0.071212f
C707 VP.t3 VSUBS 0.726534f
C708 VP.n1 VSUBS 0.044785f
C709 VP.n2 VSUBS 0.054014f
C710 VP.t5 VSUBS 0.726534f
C711 VP.n3 VSUBS 0.100668f
C712 VP.n4 VSUBS 0.054014f
C713 VP.n5 VSUBS 0.061402f
C714 VP.n6 VSUBS 0.054014f
C715 VP.n7 VSUBS 0.108906f
C716 VP.n8 VSUBS 0.071212f
C717 VP.t0 VSUBS 0.726534f
C718 VP.n9 VSUBS 0.044785f
C719 VP.n10 VSUBS 0.054014f
C720 VP.t6 VSUBS 0.726534f
C721 VP.n11 VSUBS 0.100668f
C722 VP.n12 VSUBS 0.054014f
C723 VP.n13 VSUBS 0.061402f
C724 VP.t7 VSUBS 1.09712f
C725 VP.t4 VSUBS 0.726534f
C726 VP.n14 VSUBS 0.465911f
C727 VP.n15 VSUBS 0.458542f
C728 VP.n16 VSUBS 0.469448f
C729 VP.n17 VSUBS 0.054014f
C730 VP.n18 VSUBS 0.100668f
C731 VP.n19 VSUBS 0.07885f
C732 VP.n20 VSUBS 0.07885f
C733 VP.n21 VSUBS 0.054014f
C734 VP.n22 VSUBS 0.054014f
C735 VP.n23 VSUBS 0.054014f
C736 VP.n24 VSUBS 0.061402f
C737 VP.n25 VSUBS 0.331903f
C738 VP.n26 VSUBS 0.090228f
C739 VP.n27 VSUBS 0.104678f
C740 VP.n28 VSUBS 0.054014f
C741 VP.n29 VSUBS 0.054014f
C742 VP.n30 VSUBS 0.054014f
C743 VP.n31 VSUBS 0.108906f
C744 VP.n32 VSUBS 0.082276f
C745 VP.n33 VSUBS 0.51362f
C746 VP.n34 VSUBS 2.34101f
C747 VP.n35 VSUBS 2.38658f
C748 VP.t2 VSUBS 0.726534f
C749 VP.n36 VSUBS 0.51362f
C750 VP.n37 VSUBS 0.082276f
C751 VP.n38 VSUBS 0.071212f
C752 VP.n39 VSUBS 0.054014f
C753 VP.n40 VSUBS 0.054014f
C754 VP.n41 VSUBS 0.044785f
C755 VP.n42 VSUBS 0.104678f
C756 VP.t1 VSUBS 0.726534f
C757 VP.n43 VSUBS 0.331903f
C758 VP.n44 VSUBS 0.090228f
C759 VP.n45 VSUBS 0.054014f
C760 VP.n46 VSUBS 0.054014f
C761 VP.n47 VSUBS 0.054014f
C762 VP.n48 VSUBS 0.100668f
C763 VP.n49 VSUBS 0.07885f
C764 VP.n50 VSUBS 0.07885f
C765 VP.n51 VSUBS 0.054014f
C766 VP.n52 VSUBS 0.054014f
C767 VP.n53 VSUBS 0.054014f
C768 VP.n54 VSUBS 0.061402f
C769 VP.n55 VSUBS 0.331903f
C770 VP.n56 VSUBS 0.090228f
C771 VP.n57 VSUBS 0.104678f
C772 VP.n58 VSUBS 0.054014f
C773 VP.n59 VSUBS 0.054014f
C774 VP.n60 VSUBS 0.054014f
C775 VP.n61 VSUBS 0.108906f
C776 VP.n62 VSUBS 0.082276f
C777 VP.n63 VSUBS 0.51362f
C778 VP.n64 VSUBS 0.07654f
.ends

