* NGSPICE file created from diff_pair_sample_0606.ext - technology: sky130A

.subckt diff_pair_sample_0606 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2177 pd=7.71 as=2.8782 ps=15.54 w=7.38 l=0.72
X1 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=2.8782 pd=15.54 as=0 ps=0 w=7.38 l=0.72
X2 VTAIL.t7 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.8782 pd=15.54 as=1.2177 ps=7.71 w=7.38 l=0.72
X3 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=2.8782 pd=15.54 as=0 ps=0 w=7.38 l=0.72
X4 VDD2.t3 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2177 pd=7.71 as=2.8782 ps=15.54 w=7.38 l=0.72
X5 VDD2.t2 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2177 pd=7.71 as=2.8782 ps=15.54 w=7.38 l=0.72
X6 VTAIL.t2 VN.t2 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.8782 pd=15.54 as=1.2177 ps=7.71 w=7.38 l=0.72
X7 VDD1.t1 VP.t2 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2177 pd=7.71 as=2.8782 ps=15.54 w=7.38 l=0.72
X8 VTAIL.t1 VN.t3 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.8782 pd=15.54 as=1.2177 ps=7.71 w=7.38 l=0.72
X9 VTAIL.t6 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.8782 pd=15.54 as=1.2177 ps=7.71 w=7.38 l=0.72
X10 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.8782 pd=15.54 as=0 ps=0 w=7.38 l=0.72
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.8782 pd=15.54 as=0 ps=0 w=7.38 l=0.72
R0 VP.n1 VP.t3 322.582
R1 VP.n1 VP.t0 322.531
R2 VP.n3 VP.t1 301.586
R3 VP.n5 VP.t2 301.586
R4 VP.n6 VP.n5 161.3
R5 VP.n4 VP.n0 161.3
R6 VP.n3 VP.n2 161.3
R7 VP.n2 VP.n1 81.6469
R8 VP.n4 VP.n3 24.1005
R9 VP.n5 VP.n4 24.1005
R10 VP.n2 VP.n0 0.189894
R11 VP.n6 VP.n0 0.189894
R12 VP VP.n6 0.0516364
R13 VTAIL.n314 VTAIL.n280 289.615
R14 VTAIL.n34 VTAIL.n0 289.615
R15 VTAIL.n74 VTAIL.n40 289.615
R16 VTAIL.n114 VTAIL.n80 289.615
R17 VTAIL.n274 VTAIL.n240 289.615
R18 VTAIL.n234 VTAIL.n200 289.615
R19 VTAIL.n194 VTAIL.n160 289.615
R20 VTAIL.n154 VTAIL.n120 289.615
R21 VTAIL.n292 VTAIL.n291 185
R22 VTAIL.n297 VTAIL.n296 185
R23 VTAIL.n299 VTAIL.n298 185
R24 VTAIL.n288 VTAIL.n287 185
R25 VTAIL.n305 VTAIL.n304 185
R26 VTAIL.n307 VTAIL.n306 185
R27 VTAIL.n284 VTAIL.n283 185
R28 VTAIL.n313 VTAIL.n312 185
R29 VTAIL.n315 VTAIL.n314 185
R30 VTAIL.n12 VTAIL.n11 185
R31 VTAIL.n17 VTAIL.n16 185
R32 VTAIL.n19 VTAIL.n18 185
R33 VTAIL.n8 VTAIL.n7 185
R34 VTAIL.n25 VTAIL.n24 185
R35 VTAIL.n27 VTAIL.n26 185
R36 VTAIL.n4 VTAIL.n3 185
R37 VTAIL.n33 VTAIL.n32 185
R38 VTAIL.n35 VTAIL.n34 185
R39 VTAIL.n52 VTAIL.n51 185
R40 VTAIL.n57 VTAIL.n56 185
R41 VTAIL.n59 VTAIL.n58 185
R42 VTAIL.n48 VTAIL.n47 185
R43 VTAIL.n65 VTAIL.n64 185
R44 VTAIL.n67 VTAIL.n66 185
R45 VTAIL.n44 VTAIL.n43 185
R46 VTAIL.n73 VTAIL.n72 185
R47 VTAIL.n75 VTAIL.n74 185
R48 VTAIL.n92 VTAIL.n91 185
R49 VTAIL.n97 VTAIL.n96 185
R50 VTAIL.n99 VTAIL.n98 185
R51 VTAIL.n88 VTAIL.n87 185
R52 VTAIL.n105 VTAIL.n104 185
R53 VTAIL.n107 VTAIL.n106 185
R54 VTAIL.n84 VTAIL.n83 185
R55 VTAIL.n113 VTAIL.n112 185
R56 VTAIL.n115 VTAIL.n114 185
R57 VTAIL.n275 VTAIL.n274 185
R58 VTAIL.n273 VTAIL.n272 185
R59 VTAIL.n244 VTAIL.n243 185
R60 VTAIL.n267 VTAIL.n266 185
R61 VTAIL.n265 VTAIL.n264 185
R62 VTAIL.n248 VTAIL.n247 185
R63 VTAIL.n259 VTAIL.n258 185
R64 VTAIL.n257 VTAIL.n256 185
R65 VTAIL.n252 VTAIL.n251 185
R66 VTAIL.n235 VTAIL.n234 185
R67 VTAIL.n233 VTAIL.n232 185
R68 VTAIL.n204 VTAIL.n203 185
R69 VTAIL.n227 VTAIL.n226 185
R70 VTAIL.n225 VTAIL.n224 185
R71 VTAIL.n208 VTAIL.n207 185
R72 VTAIL.n219 VTAIL.n218 185
R73 VTAIL.n217 VTAIL.n216 185
R74 VTAIL.n212 VTAIL.n211 185
R75 VTAIL.n195 VTAIL.n194 185
R76 VTAIL.n193 VTAIL.n192 185
R77 VTAIL.n164 VTAIL.n163 185
R78 VTAIL.n187 VTAIL.n186 185
R79 VTAIL.n185 VTAIL.n184 185
R80 VTAIL.n168 VTAIL.n167 185
R81 VTAIL.n179 VTAIL.n178 185
R82 VTAIL.n177 VTAIL.n176 185
R83 VTAIL.n172 VTAIL.n171 185
R84 VTAIL.n155 VTAIL.n154 185
R85 VTAIL.n153 VTAIL.n152 185
R86 VTAIL.n124 VTAIL.n123 185
R87 VTAIL.n147 VTAIL.n146 185
R88 VTAIL.n145 VTAIL.n144 185
R89 VTAIL.n128 VTAIL.n127 185
R90 VTAIL.n139 VTAIL.n138 185
R91 VTAIL.n137 VTAIL.n136 185
R92 VTAIL.n132 VTAIL.n131 185
R93 VTAIL.n293 VTAIL.t0 147.659
R94 VTAIL.n13 VTAIL.t1 147.659
R95 VTAIL.n53 VTAIL.t4 147.659
R96 VTAIL.n93 VTAIL.t7 147.659
R97 VTAIL.n253 VTAIL.t5 147.659
R98 VTAIL.n213 VTAIL.t6 147.659
R99 VTAIL.n173 VTAIL.t3 147.659
R100 VTAIL.n133 VTAIL.t2 147.659
R101 VTAIL.n297 VTAIL.n291 104.615
R102 VTAIL.n298 VTAIL.n297 104.615
R103 VTAIL.n298 VTAIL.n287 104.615
R104 VTAIL.n305 VTAIL.n287 104.615
R105 VTAIL.n306 VTAIL.n305 104.615
R106 VTAIL.n306 VTAIL.n283 104.615
R107 VTAIL.n313 VTAIL.n283 104.615
R108 VTAIL.n314 VTAIL.n313 104.615
R109 VTAIL.n17 VTAIL.n11 104.615
R110 VTAIL.n18 VTAIL.n17 104.615
R111 VTAIL.n18 VTAIL.n7 104.615
R112 VTAIL.n25 VTAIL.n7 104.615
R113 VTAIL.n26 VTAIL.n25 104.615
R114 VTAIL.n26 VTAIL.n3 104.615
R115 VTAIL.n33 VTAIL.n3 104.615
R116 VTAIL.n34 VTAIL.n33 104.615
R117 VTAIL.n57 VTAIL.n51 104.615
R118 VTAIL.n58 VTAIL.n57 104.615
R119 VTAIL.n58 VTAIL.n47 104.615
R120 VTAIL.n65 VTAIL.n47 104.615
R121 VTAIL.n66 VTAIL.n65 104.615
R122 VTAIL.n66 VTAIL.n43 104.615
R123 VTAIL.n73 VTAIL.n43 104.615
R124 VTAIL.n74 VTAIL.n73 104.615
R125 VTAIL.n97 VTAIL.n91 104.615
R126 VTAIL.n98 VTAIL.n97 104.615
R127 VTAIL.n98 VTAIL.n87 104.615
R128 VTAIL.n105 VTAIL.n87 104.615
R129 VTAIL.n106 VTAIL.n105 104.615
R130 VTAIL.n106 VTAIL.n83 104.615
R131 VTAIL.n113 VTAIL.n83 104.615
R132 VTAIL.n114 VTAIL.n113 104.615
R133 VTAIL.n274 VTAIL.n273 104.615
R134 VTAIL.n273 VTAIL.n243 104.615
R135 VTAIL.n266 VTAIL.n243 104.615
R136 VTAIL.n266 VTAIL.n265 104.615
R137 VTAIL.n265 VTAIL.n247 104.615
R138 VTAIL.n258 VTAIL.n247 104.615
R139 VTAIL.n258 VTAIL.n257 104.615
R140 VTAIL.n257 VTAIL.n251 104.615
R141 VTAIL.n234 VTAIL.n233 104.615
R142 VTAIL.n233 VTAIL.n203 104.615
R143 VTAIL.n226 VTAIL.n203 104.615
R144 VTAIL.n226 VTAIL.n225 104.615
R145 VTAIL.n225 VTAIL.n207 104.615
R146 VTAIL.n218 VTAIL.n207 104.615
R147 VTAIL.n218 VTAIL.n217 104.615
R148 VTAIL.n217 VTAIL.n211 104.615
R149 VTAIL.n194 VTAIL.n193 104.615
R150 VTAIL.n193 VTAIL.n163 104.615
R151 VTAIL.n186 VTAIL.n163 104.615
R152 VTAIL.n186 VTAIL.n185 104.615
R153 VTAIL.n185 VTAIL.n167 104.615
R154 VTAIL.n178 VTAIL.n167 104.615
R155 VTAIL.n178 VTAIL.n177 104.615
R156 VTAIL.n177 VTAIL.n171 104.615
R157 VTAIL.n154 VTAIL.n153 104.615
R158 VTAIL.n153 VTAIL.n123 104.615
R159 VTAIL.n146 VTAIL.n123 104.615
R160 VTAIL.n146 VTAIL.n145 104.615
R161 VTAIL.n145 VTAIL.n127 104.615
R162 VTAIL.n138 VTAIL.n127 104.615
R163 VTAIL.n138 VTAIL.n137 104.615
R164 VTAIL.n137 VTAIL.n131 104.615
R165 VTAIL.t0 VTAIL.n291 52.3082
R166 VTAIL.t1 VTAIL.n11 52.3082
R167 VTAIL.t4 VTAIL.n51 52.3082
R168 VTAIL.t7 VTAIL.n91 52.3082
R169 VTAIL.t5 VTAIL.n251 52.3082
R170 VTAIL.t6 VTAIL.n211 52.3082
R171 VTAIL.t3 VTAIL.n171 52.3082
R172 VTAIL.t2 VTAIL.n131 52.3082
R173 VTAIL.n319 VTAIL.n318 31.0217
R174 VTAIL.n39 VTAIL.n38 31.0217
R175 VTAIL.n79 VTAIL.n78 31.0217
R176 VTAIL.n119 VTAIL.n118 31.0217
R177 VTAIL.n279 VTAIL.n278 31.0217
R178 VTAIL.n239 VTAIL.n238 31.0217
R179 VTAIL.n199 VTAIL.n198 31.0217
R180 VTAIL.n159 VTAIL.n158 31.0217
R181 VTAIL.n319 VTAIL.n279 19.6341
R182 VTAIL.n159 VTAIL.n119 19.6341
R183 VTAIL.n293 VTAIL.n292 15.6677
R184 VTAIL.n13 VTAIL.n12 15.6677
R185 VTAIL.n53 VTAIL.n52 15.6677
R186 VTAIL.n93 VTAIL.n92 15.6677
R187 VTAIL.n253 VTAIL.n252 15.6677
R188 VTAIL.n213 VTAIL.n212 15.6677
R189 VTAIL.n173 VTAIL.n172 15.6677
R190 VTAIL.n133 VTAIL.n132 15.6677
R191 VTAIL.n296 VTAIL.n295 12.8005
R192 VTAIL.n16 VTAIL.n15 12.8005
R193 VTAIL.n56 VTAIL.n55 12.8005
R194 VTAIL.n96 VTAIL.n95 12.8005
R195 VTAIL.n256 VTAIL.n255 12.8005
R196 VTAIL.n216 VTAIL.n215 12.8005
R197 VTAIL.n176 VTAIL.n175 12.8005
R198 VTAIL.n136 VTAIL.n135 12.8005
R199 VTAIL.n299 VTAIL.n290 12.0247
R200 VTAIL.n19 VTAIL.n10 12.0247
R201 VTAIL.n59 VTAIL.n50 12.0247
R202 VTAIL.n99 VTAIL.n90 12.0247
R203 VTAIL.n259 VTAIL.n250 12.0247
R204 VTAIL.n219 VTAIL.n210 12.0247
R205 VTAIL.n179 VTAIL.n170 12.0247
R206 VTAIL.n139 VTAIL.n130 12.0247
R207 VTAIL.n300 VTAIL.n288 11.249
R208 VTAIL.n20 VTAIL.n8 11.249
R209 VTAIL.n60 VTAIL.n48 11.249
R210 VTAIL.n100 VTAIL.n88 11.249
R211 VTAIL.n260 VTAIL.n248 11.249
R212 VTAIL.n220 VTAIL.n208 11.249
R213 VTAIL.n180 VTAIL.n168 11.249
R214 VTAIL.n140 VTAIL.n128 11.249
R215 VTAIL.n304 VTAIL.n303 10.4732
R216 VTAIL.n24 VTAIL.n23 10.4732
R217 VTAIL.n64 VTAIL.n63 10.4732
R218 VTAIL.n104 VTAIL.n103 10.4732
R219 VTAIL.n264 VTAIL.n263 10.4732
R220 VTAIL.n224 VTAIL.n223 10.4732
R221 VTAIL.n184 VTAIL.n183 10.4732
R222 VTAIL.n144 VTAIL.n143 10.4732
R223 VTAIL.n307 VTAIL.n286 9.69747
R224 VTAIL.n27 VTAIL.n6 9.69747
R225 VTAIL.n67 VTAIL.n46 9.69747
R226 VTAIL.n107 VTAIL.n86 9.69747
R227 VTAIL.n267 VTAIL.n246 9.69747
R228 VTAIL.n227 VTAIL.n206 9.69747
R229 VTAIL.n187 VTAIL.n166 9.69747
R230 VTAIL.n147 VTAIL.n126 9.69747
R231 VTAIL.n318 VTAIL.n317 9.45567
R232 VTAIL.n38 VTAIL.n37 9.45567
R233 VTAIL.n78 VTAIL.n77 9.45567
R234 VTAIL.n118 VTAIL.n117 9.45567
R235 VTAIL.n278 VTAIL.n277 9.45567
R236 VTAIL.n238 VTAIL.n237 9.45567
R237 VTAIL.n198 VTAIL.n197 9.45567
R238 VTAIL.n158 VTAIL.n157 9.45567
R239 VTAIL.n317 VTAIL.n316 9.3005
R240 VTAIL.n311 VTAIL.n310 9.3005
R241 VTAIL.n309 VTAIL.n308 9.3005
R242 VTAIL.n286 VTAIL.n285 9.3005
R243 VTAIL.n303 VTAIL.n302 9.3005
R244 VTAIL.n301 VTAIL.n300 9.3005
R245 VTAIL.n290 VTAIL.n289 9.3005
R246 VTAIL.n295 VTAIL.n294 9.3005
R247 VTAIL.n282 VTAIL.n281 9.3005
R248 VTAIL.n37 VTAIL.n36 9.3005
R249 VTAIL.n31 VTAIL.n30 9.3005
R250 VTAIL.n29 VTAIL.n28 9.3005
R251 VTAIL.n6 VTAIL.n5 9.3005
R252 VTAIL.n23 VTAIL.n22 9.3005
R253 VTAIL.n21 VTAIL.n20 9.3005
R254 VTAIL.n10 VTAIL.n9 9.3005
R255 VTAIL.n15 VTAIL.n14 9.3005
R256 VTAIL.n2 VTAIL.n1 9.3005
R257 VTAIL.n77 VTAIL.n76 9.3005
R258 VTAIL.n71 VTAIL.n70 9.3005
R259 VTAIL.n69 VTAIL.n68 9.3005
R260 VTAIL.n46 VTAIL.n45 9.3005
R261 VTAIL.n63 VTAIL.n62 9.3005
R262 VTAIL.n61 VTAIL.n60 9.3005
R263 VTAIL.n50 VTAIL.n49 9.3005
R264 VTAIL.n55 VTAIL.n54 9.3005
R265 VTAIL.n42 VTAIL.n41 9.3005
R266 VTAIL.n117 VTAIL.n116 9.3005
R267 VTAIL.n111 VTAIL.n110 9.3005
R268 VTAIL.n109 VTAIL.n108 9.3005
R269 VTAIL.n86 VTAIL.n85 9.3005
R270 VTAIL.n103 VTAIL.n102 9.3005
R271 VTAIL.n101 VTAIL.n100 9.3005
R272 VTAIL.n90 VTAIL.n89 9.3005
R273 VTAIL.n95 VTAIL.n94 9.3005
R274 VTAIL.n82 VTAIL.n81 9.3005
R275 VTAIL.n277 VTAIL.n276 9.3005
R276 VTAIL.n242 VTAIL.n241 9.3005
R277 VTAIL.n271 VTAIL.n270 9.3005
R278 VTAIL.n269 VTAIL.n268 9.3005
R279 VTAIL.n246 VTAIL.n245 9.3005
R280 VTAIL.n263 VTAIL.n262 9.3005
R281 VTAIL.n261 VTAIL.n260 9.3005
R282 VTAIL.n250 VTAIL.n249 9.3005
R283 VTAIL.n255 VTAIL.n254 9.3005
R284 VTAIL.n237 VTAIL.n236 9.3005
R285 VTAIL.n202 VTAIL.n201 9.3005
R286 VTAIL.n231 VTAIL.n230 9.3005
R287 VTAIL.n229 VTAIL.n228 9.3005
R288 VTAIL.n206 VTAIL.n205 9.3005
R289 VTAIL.n223 VTAIL.n222 9.3005
R290 VTAIL.n221 VTAIL.n220 9.3005
R291 VTAIL.n210 VTAIL.n209 9.3005
R292 VTAIL.n215 VTAIL.n214 9.3005
R293 VTAIL.n197 VTAIL.n196 9.3005
R294 VTAIL.n162 VTAIL.n161 9.3005
R295 VTAIL.n191 VTAIL.n190 9.3005
R296 VTAIL.n189 VTAIL.n188 9.3005
R297 VTAIL.n166 VTAIL.n165 9.3005
R298 VTAIL.n183 VTAIL.n182 9.3005
R299 VTAIL.n181 VTAIL.n180 9.3005
R300 VTAIL.n170 VTAIL.n169 9.3005
R301 VTAIL.n175 VTAIL.n174 9.3005
R302 VTAIL.n157 VTAIL.n156 9.3005
R303 VTAIL.n122 VTAIL.n121 9.3005
R304 VTAIL.n151 VTAIL.n150 9.3005
R305 VTAIL.n149 VTAIL.n148 9.3005
R306 VTAIL.n126 VTAIL.n125 9.3005
R307 VTAIL.n143 VTAIL.n142 9.3005
R308 VTAIL.n141 VTAIL.n140 9.3005
R309 VTAIL.n130 VTAIL.n129 9.3005
R310 VTAIL.n135 VTAIL.n134 9.3005
R311 VTAIL.n308 VTAIL.n284 8.92171
R312 VTAIL.n28 VTAIL.n4 8.92171
R313 VTAIL.n68 VTAIL.n44 8.92171
R314 VTAIL.n108 VTAIL.n84 8.92171
R315 VTAIL.n268 VTAIL.n244 8.92171
R316 VTAIL.n228 VTAIL.n204 8.92171
R317 VTAIL.n188 VTAIL.n164 8.92171
R318 VTAIL.n148 VTAIL.n124 8.92171
R319 VTAIL.n312 VTAIL.n311 8.14595
R320 VTAIL.n32 VTAIL.n31 8.14595
R321 VTAIL.n72 VTAIL.n71 8.14595
R322 VTAIL.n112 VTAIL.n111 8.14595
R323 VTAIL.n272 VTAIL.n271 8.14595
R324 VTAIL.n232 VTAIL.n231 8.14595
R325 VTAIL.n192 VTAIL.n191 8.14595
R326 VTAIL.n152 VTAIL.n151 8.14595
R327 VTAIL.n315 VTAIL.n282 7.3702
R328 VTAIL.n318 VTAIL.n280 7.3702
R329 VTAIL.n35 VTAIL.n2 7.3702
R330 VTAIL.n38 VTAIL.n0 7.3702
R331 VTAIL.n75 VTAIL.n42 7.3702
R332 VTAIL.n78 VTAIL.n40 7.3702
R333 VTAIL.n115 VTAIL.n82 7.3702
R334 VTAIL.n118 VTAIL.n80 7.3702
R335 VTAIL.n278 VTAIL.n240 7.3702
R336 VTAIL.n275 VTAIL.n242 7.3702
R337 VTAIL.n238 VTAIL.n200 7.3702
R338 VTAIL.n235 VTAIL.n202 7.3702
R339 VTAIL.n198 VTAIL.n160 7.3702
R340 VTAIL.n195 VTAIL.n162 7.3702
R341 VTAIL.n158 VTAIL.n120 7.3702
R342 VTAIL.n155 VTAIL.n122 7.3702
R343 VTAIL.n316 VTAIL.n315 6.59444
R344 VTAIL.n316 VTAIL.n280 6.59444
R345 VTAIL.n36 VTAIL.n35 6.59444
R346 VTAIL.n36 VTAIL.n0 6.59444
R347 VTAIL.n76 VTAIL.n75 6.59444
R348 VTAIL.n76 VTAIL.n40 6.59444
R349 VTAIL.n116 VTAIL.n115 6.59444
R350 VTAIL.n116 VTAIL.n80 6.59444
R351 VTAIL.n276 VTAIL.n240 6.59444
R352 VTAIL.n276 VTAIL.n275 6.59444
R353 VTAIL.n236 VTAIL.n200 6.59444
R354 VTAIL.n236 VTAIL.n235 6.59444
R355 VTAIL.n196 VTAIL.n160 6.59444
R356 VTAIL.n196 VTAIL.n195 6.59444
R357 VTAIL.n156 VTAIL.n120 6.59444
R358 VTAIL.n156 VTAIL.n155 6.59444
R359 VTAIL.n312 VTAIL.n282 5.81868
R360 VTAIL.n32 VTAIL.n2 5.81868
R361 VTAIL.n72 VTAIL.n42 5.81868
R362 VTAIL.n112 VTAIL.n82 5.81868
R363 VTAIL.n272 VTAIL.n242 5.81868
R364 VTAIL.n232 VTAIL.n202 5.81868
R365 VTAIL.n192 VTAIL.n162 5.81868
R366 VTAIL.n152 VTAIL.n122 5.81868
R367 VTAIL.n311 VTAIL.n284 5.04292
R368 VTAIL.n31 VTAIL.n4 5.04292
R369 VTAIL.n71 VTAIL.n44 5.04292
R370 VTAIL.n111 VTAIL.n84 5.04292
R371 VTAIL.n271 VTAIL.n244 5.04292
R372 VTAIL.n231 VTAIL.n204 5.04292
R373 VTAIL.n191 VTAIL.n164 5.04292
R374 VTAIL.n151 VTAIL.n124 5.04292
R375 VTAIL.n254 VTAIL.n253 4.38565
R376 VTAIL.n214 VTAIL.n213 4.38565
R377 VTAIL.n174 VTAIL.n173 4.38565
R378 VTAIL.n134 VTAIL.n133 4.38565
R379 VTAIL.n294 VTAIL.n293 4.38565
R380 VTAIL.n14 VTAIL.n13 4.38565
R381 VTAIL.n54 VTAIL.n53 4.38565
R382 VTAIL.n94 VTAIL.n93 4.38565
R383 VTAIL.n308 VTAIL.n307 4.26717
R384 VTAIL.n28 VTAIL.n27 4.26717
R385 VTAIL.n68 VTAIL.n67 4.26717
R386 VTAIL.n108 VTAIL.n107 4.26717
R387 VTAIL.n268 VTAIL.n267 4.26717
R388 VTAIL.n228 VTAIL.n227 4.26717
R389 VTAIL.n188 VTAIL.n187 4.26717
R390 VTAIL.n148 VTAIL.n147 4.26717
R391 VTAIL.n304 VTAIL.n286 3.49141
R392 VTAIL.n24 VTAIL.n6 3.49141
R393 VTAIL.n64 VTAIL.n46 3.49141
R394 VTAIL.n104 VTAIL.n86 3.49141
R395 VTAIL.n264 VTAIL.n246 3.49141
R396 VTAIL.n224 VTAIL.n206 3.49141
R397 VTAIL.n184 VTAIL.n166 3.49141
R398 VTAIL.n144 VTAIL.n126 3.49141
R399 VTAIL.n303 VTAIL.n288 2.71565
R400 VTAIL.n23 VTAIL.n8 2.71565
R401 VTAIL.n63 VTAIL.n48 2.71565
R402 VTAIL.n103 VTAIL.n88 2.71565
R403 VTAIL.n263 VTAIL.n248 2.71565
R404 VTAIL.n223 VTAIL.n208 2.71565
R405 VTAIL.n183 VTAIL.n168 2.71565
R406 VTAIL.n143 VTAIL.n128 2.71565
R407 VTAIL.n300 VTAIL.n299 1.93989
R408 VTAIL.n20 VTAIL.n19 1.93989
R409 VTAIL.n60 VTAIL.n59 1.93989
R410 VTAIL.n100 VTAIL.n99 1.93989
R411 VTAIL.n260 VTAIL.n259 1.93989
R412 VTAIL.n220 VTAIL.n219 1.93989
R413 VTAIL.n180 VTAIL.n179 1.93989
R414 VTAIL.n140 VTAIL.n139 1.93989
R415 VTAIL.n296 VTAIL.n290 1.16414
R416 VTAIL.n16 VTAIL.n10 1.16414
R417 VTAIL.n56 VTAIL.n50 1.16414
R418 VTAIL.n96 VTAIL.n90 1.16414
R419 VTAIL.n256 VTAIL.n250 1.16414
R420 VTAIL.n216 VTAIL.n210 1.16414
R421 VTAIL.n176 VTAIL.n170 1.16414
R422 VTAIL.n136 VTAIL.n130 1.16414
R423 VTAIL.n199 VTAIL.n159 0.905672
R424 VTAIL.n279 VTAIL.n239 0.905672
R425 VTAIL.n119 VTAIL.n79 0.905672
R426 VTAIL VTAIL.n39 0.511276
R427 VTAIL.n239 VTAIL.n199 0.470328
R428 VTAIL.n79 VTAIL.n39 0.470328
R429 VTAIL VTAIL.n319 0.394897
R430 VTAIL.n295 VTAIL.n292 0.388379
R431 VTAIL.n15 VTAIL.n12 0.388379
R432 VTAIL.n55 VTAIL.n52 0.388379
R433 VTAIL.n95 VTAIL.n92 0.388379
R434 VTAIL.n255 VTAIL.n252 0.388379
R435 VTAIL.n215 VTAIL.n212 0.388379
R436 VTAIL.n175 VTAIL.n172 0.388379
R437 VTAIL.n135 VTAIL.n132 0.388379
R438 VTAIL.n294 VTAIL.n289 0.155672
R439 VTAIL.n301 VTAIL.n289 0.155672
R440 VTAIL.n302 VTAIL.n301 0.155672
R441 VTAIL.n302 VTAIL.n285 0.155672
R442 VTAIL.n309 VTAIL.n285 0.155672
R443 VTAIL.n310 VTAIL.n309 0.155672
R444 VTAIL.n310 VTAIL.n281 0.155672
R445 VTAIL.n317 VTAIL.n281 0.155672
R446 VTAIL.n14 VTAIL.n9 0.155672
R447 VTAIL.n21 VTAIL.n9 0.155672
R448 VTAIL.n22 VTAIL.n21 0.155672
R449 VTAIL.n22 VTAIL.n5 0.155672
R450 VTAIL.n29 VTAIL.n5 0.155672
R451 VTAIL.n30 VTAIL.n29 0.155672
R452 VTAIL.n30 VTAIL.n1 0.155672
R453 VTAIL.n37 VTAIL.n1 0.155672
R454 VTAIL.n54 VTAIL.n49 0.155672
R455 VTAIL.n61 VTAIL.n49 0.155672
R456 VTAIL.n62 VTAIL.n61 0.155672
R457 VTAIL.n62 VTAIL.n45 0.155672
R458 VTAIL.n69 VTAIL.n45 0.155672
R459 VTAIL.n70 VTAIL.n69 0.155672
R460 VTAIL.n70 VTAIL.n41 0.155672
R461 VTAIL.n77 VTAIL.n41 0.155672
R462 VTAIL.n94 VTAIL.n89 0.155672
R463 VTAIL.n101 VTAIL.n89 0.155672
R464 VTAIL.n102 VTAIL.n101 0.155672
R465 VTAIL.n102 VTAIL.n85 0.155672
R466 VTAIL.n109 VTAIL.n85 0.155672
R467 VTAIL.n110 VTAIL.n109 0.155672
R468 VTAIL.n110 VTAIL.n81 0.155672
R469 VTAIL.n117 VTAIL.n81 0.155672
R470 VTAIL.n277 VTAIL.n241 0.155672
R471 VTAIL.n270 VTAIL.n241 0.155672
R472 VTAIL.n270 VTAIL.n269 0.155672
R473 VTAIL.n269 VTAIL.n245 0.155672
R474 VTAIL.n262 VTAIL.n245 0.155672
R475 VTAIL.n262 VTAIL.n261 0.155672
R476 VTAIL.n261 VTAIL.n249 0.155672
R477 VTAIL.n254 VTAIL.n249 0.155672
R478 VTAIL.n237 VTAIL.n201 0.155672
R479 VTAIL.n230 VTAIL.n201 0.155672
R480 VTAIL.n230 VTAIL.n229 0.155672
R481 VTAIL.n229 VTAIL.n205 0.155672
R482 VTAIL.n222 VTAIL.n205 0.155672
R483 VTAIL.n222 VTAIL.n221 0.155672
R484 VTAIL.n221 VTAIL.n209 0.155672
R485 VTAIL.n214 VTAIL.n209 0.155672
R486 VTAIL.n197 VTAIL.n161 0.155672
R487 VTAIL.n190 VTAIL.n161 0.155672
R488 VTAIL.n190 VTAIL.n189 0.155672
R489 VTAIL.n189 VTAIL.n165 0.155672
R490 VTAIL.n182 VTAIL.n165 0.155672
R491 VTAIL.n182 VTAIL.n181 0.155672
R492 VTAIL.n181 VTAIL.n169 0.155672
R493 VTAIL.n174 VTAIL.n169 0.155672
R494 VTAIL.n157 VTAIL.n121 0.155672
R495 VTAIL.n150 VTAIL.n121 0.155672
R496 VTAIL.n150 VTAIL.n149 0.155672
R497 VTAIL.n149 VTAIL.n125 0.155672
R498 VTAIL.n142 VTAIL.n125 0.155672
R499 VTAIL.n142 VTAIL.n141 0.155672
R500 VTAIL.n141 VTAIL.n129 0.155672
R501 VTAIL.n134 VTAIL.n129 0.155672
R502 VDD1 VDD1.n1 97.3539
R503 VDD1 VDD1.n0 64.0949
R504 VDD1.n0 VDD1.t0 2.68343
R505 VDD1.n0 VDD1.t3 2.68343
R506 VDD1.n1 VDD1.t2 2.68343
R507 VDD1.n1 VDD1.t1 2.68343
R508 B.n482 B.n481 585
R509 B.n203 B.n68 585
R510 B.n202 B.n201 585
R511 B.n200 B.n199 585
R512 B.n198 B.n197 585
R513 B.n196 B.n195 585
R514 B.n194 B.n193 585
R515 B.n192 B.n191 585
R516 B.n190 B.n189 585
R517 B.n188 B.n187 585
R518 B.n186 B.n185 585
R519 B.n184 B.n183 585
R520 B.n182 B.n181 585
R521 B.n180 B.n179 585
R522 B.n178 B.n177 585
R523 B.n176 B.n175 585
R524 B.n174 B.n173 585
R525 B.n172 B.n171 585
R526 B.n170 B.n169 585
R527 B.n168 B.n167 585
R528 B.n166 B.n165 585
R529 B.n164 B.n163 585
R530 B.n162 B.n161 585
R531 B.n160 B.n159 585
R532 B.n158 B.n157 585
R533 B.n156 B.n155 585
R534 B.n154 B.n153 585
R535 B.n152 B.n151 585
R536 B.n150 B.n149 585
R537 B.n148 B.n147 585
R538 B.n146 B.n145 585
R539 B.n144 B.n143 585
R540 B.n142 B.n141 585
R541 B.n140 B.n139 585
R542 B.n138 B.n137 585
R543 B.n136 B.n135 585
R544 B.n134 B.n133 585
R545 B.n132 B.n131 585
R546 B.n130 B.n129 585
R547 B.n128 B.n127 585
R548 B.n126 B.n125 585
R549 B.n124 B.n123 585
R550 B.n122 B.n121 585
R551 B.n120 B.n119 585
R552 B.n118 B.n117 585
R553 B.n116 B.n115 585
R554 B.n114 B.n113 585
R555 B.n112 B.n111 585
R556 B.n110 B.n109 585
R557 B.n108 B.n107 585
R558 B.n106 B.n105 585
R559 B.n104 B.n103 585
R560 B.n102 B.n101 585
R561 B.n100 B.n99 585
R562 B.n98 B.n97 585
R563 B.n96 B.n95 585
R564 B.n94 B.n93 585
R565 B.n92 B.n91 585
R566 B.n90 B.n89 585
R567 B.n88 B.n87 585
R568 B.n86 B.n85 585
R569 B.n84 B.n83 585
R570 B.n82 B.n81 585
R571 B.n80 B.n79 585
R572 B.n78 B.n77 585
R573 B.n76 B.n75 585
R574 B.n480 B.n35 585
R575 B.n485 B.n35 585
R576 B.n479 B.n34 585
R577 B.n486 B.n34 585
R578 B.n478 B.n477 585
R579 B.n477 B.n30 585
R580 B.n476 B.n29 585
R581 B.n492 B.n29 585
R582 B.n475 B.n28 585
R583 B.n493 B.n28 585
R584 B.n474 B.n27 585
R585 B.n494 B.n27 585
R586 B.n473 B.n472 585
R587 B.n472 B.n23 585
R588 B.n471 B.n22 585
R589 B.n500 B.n22 585
R590 B.n470 B.n21 585
R591 B.n501 B.n21 585
R592 B.n469 B.n20 585
R593 B.n502 B.n20 585
R594 B.n468 B.n467 585
R595 B.n467 B.n16 585
R596 B.n466 B.n15 585
R597 B.n508 B.n15 585
R598 B.n465 B.n14 585
R599 B.n509 B.n14 585
R600 B.n464 B.n13 585
R601 B.n510 B.n13 585
R602 B.n463 B.n462 585
R603 B.n462 B.n12 585
R604 B.n461 B.n460 585
R605 B.n461 B.n8 585
R606 B.n459 B.n7 585
R607 B.n517 B.n7 585
R608 B.n458 B.n6 585
R609 B.n518 B.n6 585
R610 B.n457 B.n5 585
R611 B.n519 B.n5 585
R612 B.n456 B.n455 585
R613 B.n455 B.n4 585
R614 B.n454 B.n204 585
R615 B.n454 B.n453 585
R616 B.n443 B.n205 585
R617 B.n446 B.n205 585
R618 B.n445 B.n444 585
R619 B.n447 B.n445 585
R620 B.n442 B.n210 585
R621 B.n210 B.n209 585
R622 B.n441 B.n440 585
R623 B.n440 B.n439 585
R624 B.n212 B.n211 585
R625 B.n213 B.n212 585
R626 B.n432 B.n431 585
R627 B.n433 B.n432 585
R628 B.n430 B.n218 585
R629 B.n218 B.n217 585
R630 B.n429 B.n428 585
R631 B.n428 B.n427 585
R632 B.n220 B.n219 585
R633 B.n221 B.n220 585
R634 B.n420 B.n419 585
R635 B.n421 B.n420 585
R636 B.n418 B.n225 585
R637 B.n229 B.n225 585
R638 B.n417 B.n416 585
R639 B.n416 B.n415 585
R640 B.n227 B.n226 585
R641 B.n228 B.n227 585
R642 B.n408 B.n407 585
R643 B.n409 B.n408 585
R644 B.n406 B.n234 585
R645 B.n234 B.n233 585
R646 B.n401 B.n400 585
R647 B.n399 B.n269 585
R648 B.n398 B.n268 585
R649 B.n403 B.n268 585
R650 B.n397 B.n396 585
R651 B.n395 B.n394 585
R652 B.n393 B.n392 585
R653 B.n391 B.n390 585
R654 B.n389 B.n388 585
R655 B.n387 B.n386 585
R656 B.n385 B.n384 585
R657 B.n383 B.n382 585
R658 B.n381 B.n380 585
R659 B.n379 B.n378 585
R660 B.n377 B.n376 585
R661 B.n375 B.n374 585
R662 B.n373 B.n372 585
R663 B.n371 B.n370 585
R664 B.n369 B.n368 585
R665 B.n367 B.n366 585
R666 B.n365 B.n364 585
R667 B.n363 B.n362 585
R668 B.n361 B.n360 585
R669 B.n359 B.n358 585
R670 B.n357 B.n356 585
R671 B.n355 B.n354 585
R672 B.n353 B.n352 585
R673 B.n351 B.n350 585
R674 B.n349 B.n348 585
R675 B.n346 B.n345 585
R676 B.n344 B.n343 585
R677 B.n342 B.n341 585
R678 B.n340 B.n339 585
R679 B.n338 B.n337 585
R680 B.n336 B.n335 585
R681 B.n334 B.n333 585
R682 B.n332 B.n331 585
R683 B.n330 B.n329 585
R684 B.n328 B.n327 585
R685 B.n325 B.n324 585
R686 B.n323 B.n322 585
R687 B.n321 B.n320 585
R688 B.n319 B.n318 585
R689 B.n317 B.n316 585
R690 B.n315 B.n314 585
R691 B.n313 B.n312 585
R692 B.n311 B.n310 585
R693 B.n309 B.n308 585
R694 B.n307 B.n306 585
R695 B.n305 B.n304 585
R696 B.n303 B.n302 585
R697 B.n301 B.n300 585
R698 B.n299 B.n298 585
R699 B.n297 B.n296 585
R700 B.n295 B.n294 585
R701 B.n293 B.n292 585
R702 B.n291 B.n290 585
R703 B.n289 B.n288 585
R704 B.n287 B.n286 585
R705 B.n285 B.n284 585
R706 B.n283 B.n282 585
R707 B.n281 B.n280 585
R708 B.n279 B.n278 585
R709 B.n277 B.n276 585
R710 B.n275 B.n274 585
R711 B.n236 B.n235 585
R712 B.n405 B.n404 585
R713 B.n404 B.n403 585
R714 B.n232 B.n231 585
R715 B.n233 B.n232 585
R716 B.n411 B.n410 585
R717 B.n410 B.n409 585
R718 B.n412 B.n230 585
R719 B.n230 B.n228 585
R720 B.n414 B.n413 585
R721 B.n415 B.n414 585
R722 B.n224 B.n223 585
R723 B.n229 B.n224 585
R724 B.n423 B.n422 585
R725 B.n422 B.n421 585
R726 B.n424 B.n222 585
R727 B.n222 B.n221 585
R728 B.n426 B.n425 585
R729 B.n427 B.n426 585
R730 B.n216 B.n215 585
R731 B.n217 B.n216 585
R732 B.n435 B.n434 585
R733 B.n434 B.n433 585
R734 B.n436 B.n214 585
R735 B.n214 B.n213 585
R736 B.n438 B.n437 585
R737 B.n439 B.n438 585
R738 B.n208 B.n207 585
R739 B.n209 B.n208 585
R740 B.n449 B.n448 585
R741 B.n448 B.n447 585
R742 B.n450 B.n206 585
R743 B.n446 B.n206 585
R744 B.n452 B.n451 585
R745 B.n453 B.n452 585
R746 B.n3 B.n0 585
R747 B.n4 B.n3 585
R748 B.n516 B.n1 585
R749 B.n517 B.n516 585
R750 B.n515 B.n514 585
R751 B.n515 B.n8 585
R752 B.n513 B.n9 585
R753 B.n12 B.n9 585
R754 B.n512 B.n511 585
R755 B.n511 B.n510 585
R756 B.n11 B.n10 585
R757 B.n509 B.n11 585
R758 B.n507 B.n506 585
R759 B.n508 B.n507 585
R760 B.n505 B.n17 585
R761 B.n17 B.n16 585
R762 B.n504 B.n503 585
R763 B.n503 B.n502 585
R764 B.n19 B.n18 585
R765 B.n501 B.n19 585
R766 B.n499 B.n498 585
R767 B.n500 B.n499 585
R768 B.n497 B.n24 585
R769 B.n24 B.n23 585
R770 B.n496 B.n495 585
R771 B.n495 B.n494 585
R772 B.n26 B.n25 585
R773 B.n493 B.n26 585
R774 B.n491 B.n490 585
R775 B.n492 B.n491 585
R776 B.n489 B.n31 585
R777 B.n31 B.n30 585
R778 B.n488 B.n487 585
R779 B.n487 B.n486 585
R780 B.n33 B.n32 585
R781 B.n485 B.n33 585
R782 B.n520 B.n519 585
R783 B.n518 B.n2 585
R784 B.n72 B.t4 449.752
R785 B.n69 B.t15 449.752
R786 B.n272 B.t8 449.752
R787 B.n270 B.t12 449.752
R788 B.n75 B.n33 449.257
R789 B.n482 B.n35 449.257
R790 B.n404 B.n234 449.257
R791 B.n401 B.n232 449.257
R792 B.n484 B.n483 256.663
R793 B.n484 B.n67 256.663
R794 B.n484 B.n66 256.663
R795 B.n484 B.n65 256.663
R796 B.n484 B.n64 256.663
R797 B.n484 B.n63 256.663
R798 B.n484 B.n62 256.663
R799 B.n484 B.n61 256.663
R800 B.n484 B.n60 256.663
R801 B.n484 B.n59 256.663
R802 B.n484 B.n58 256.663
R803 B.n484 B.n57 256.663
R804 B.n484 B.n56 256.663
R805 B.n484 B.n55 256.663
R806 B.n484 B.n54 256.663
R807 B.n484 B.n53 256.663
R808 B.n484 B.n52 256.663
R809 B.n484 B.n51 256.663
R810 B.n484 B.n50 256.663
R811 B.n484 B.n49 256.663
R812 B.n484 B.n48 256.663
R813 B.n484 B.n47 256.663
R814 B.n484 B.n46 256.663
R815 B.n484 B.n45 256.663
R816 B.n484 B.n44 256.663
R817 B.n484 B.n43 256.663
R818 B.n484 B.n42 256.663
R819 B.n484 B.n41 256.663
R820 B.n484 B.n40 256.663
R821 B.n484 B.n39 256.663
R822 B.n484 B.n38 256.663
R823 B.n484 B.n37 256.663
R824 B.n484 B.n36 256.663
R825 B.n403 B.n402 256.663
R826 B.n403 B.n237 256.663
R827 B.n403 B.n238 256.663
R828 B.n403 B.n239 256.663
R829 B.n403 B.n240 256.663
R830 B.n403 B.n241 256.663
R831 B.n403 B.n242 256.663
R832 B.n403 B.n243 256.663
R833 B.n403 B.n244 256.663
R834 B.n403 B.n245 256.663
R835 B.n403 B.n246 256.663
R836 B.n403 B.n247 256.663
R837 B.n403 B.n248 256.663
R838 B.n403 B.n249 256.663
R839 B.n403 B.n250 256.663
R840 B.n403 B.n251 256.663
R841 B.n403 B.n252 256.663
R842 B.n403 B.n253 256.663
R843 B.n403 B.n254 256.663
R844 B.n403 B.n255 256.663
R845 B.n403 B.n256 256.663
R846 B.n403 B.n257 256.663
R847 B.n403 B.n258 256.663
R848 B.n403 B.n259 256.663
R849 B.n403 B.n260 256.663
R850 B.n403 B.n261 256.663
R851 B.n403 B.n262 256.663
R852 B.n403 B.n263 256.663
R853 B.n403 B.n264 256.663
R854 B.n403 B.n265 256.663
R855 B.n403 B.n266 256.663
R856 B.n403 B.n267 256.663
R857 B.n522 B.n521 256.663
R858 B.n69 B.t16 223.113
R859 B.n272 B.t11 223.113
R860 B.n72 B.t6 223.113
R861 B.n270 B.t14 223.113
R862 B.n70 B.t17 202.75
R863 B.n273 B.t10 202.75
R864 B.n73 B.t7 202.75
R865 B.n271 B.t13 202.75
R866 B.n79 B.n78 163.367
R867 B.n83 B.n82 163.367
R868 B.n87 B.n86 163.367
R869 B.n91 B.n90 163.367
R870 B.n95 B.n94 163.367
R871 B.n99 B.n98 163.367
R872 B.n103 B.n102 163.367
R873 B.n107 B.n106 163.367
R874 B.n111 B.n110 163.367
R875 B.n115 B.n114 163.367
R876 B.n119 B.n118 163.367
R877 B.n123 B.n122 163.367
R878 B.n127 B.n126 163.367
R879 B.n131 B.n130 163.367
R880 B.n135 B.n134 163.367
R881 B.n139 B.n138 163.367
R882 B.n143 B.n142 163.367
R883 B.n147 B.n146 163.367
R884 B.n151 B.n150 163.367
R885 B.n155 B.n154 163.367
R886 B.n159 B.n158 163.367
R887 B.n163 B.n162 163.367
R888 B.n167 B.n166 163.367
R889 B.n171 B.n170 163.367
R890 B.n175 B.n174 163.367
R891 B.n179 B.n178 163.367
R892 B.n183 B.n182 163.367
R893 B.n187 B.n186 163.367
R894 B.n191 B.n190 163.367
R895 B.n195 B.n194 163.367
R896 B.n199 B.n198 163.367
R897 B.n201 B.n68 163.367
R898 B.n408 B.n234 163.367
R899 B.n408 B.n227 163.367
R900 B.n416 B.n227 163.367
R901 B.n416 B.n225 163.367
R902 B.n420 B.n225 163.367
R903 B.n420 B.n220 163.367
R904 B.n428 B.n220 163.367
R905 B.n428 B.n218 163.367
R906 B.n432 B.n218 163.367
R907 B.n432 B.n212 163.367
R908 B.n440 B.n212 163.367
R909 B.n440 B.n210 163.367
R910 B.n445 B.n210 163.367
R911 B.n445 B.n205 163.367
R912 B.n454 B.n205 163.367
R913 B.n455 B.n454 163.367
R914 B.n455 B.n5 163.367
R915 B.n6 B.n5 163.367
R916 B.n7 B.n6 163.367
R917 B.n461 B.n7 163.367
R918 B.n462 B.n461 163.367
R919 B.n462 B.n13 163.367
R920 B.n14 B.n13 163.367
R921 B.n15 B.n14 163.367
R922 B.n467 B.n15 163.367
R923 B.n467 B.n20 163.367
R924 B.n21 B.n20 163.367
R925 B.n22 B.n21 163.367
R926 B.n472 B.n22 163.367
R927 B.n472 B.n27 163.367
R928 B.n28 B.n27 163.367
R929 B.n29 B.n28 163.367
R930 B.n477 B.n29 163.367
R931 B.n477 B.n34 163.367
R932 B.n35 B.n34 163.367
R933 B.n269 B.n268 163.367
R934 B.n396 B.n268 163.367
R935 B.n394 B.n393 163.367
R936 B.n390 B.n389 163.367
R937 B.n386 B.n385 163.367
R938 B.n382 B.n381 163.367
R939 B.n378 B.n377 163.367
R940 B.n374 B.n373 163.367
R941 B.n370 B.n369 163.367
R942 B.n366 B.n365 163.367
R943 B.n362 B.n361 163.367
R944 B.n358 B.n357 163.367
R945 B.n354 B.n353 163.367
R946 B.n350 B.n349 163.367
R947 B.n345 B.n344 163.367
R948 B.n341 B.n340 163.367
R949 B.n337 B.n336 163.367
R950 B.n333 B.n332 163.367
R951 B.n329 B.n328 163.367
R952 B.n324 B.n323 163.367
R953 B.n320 B.n319 163.367
R954 B.n316 B.n315 163.367
R955 B.n312 B.n311 163.367
R956 B.n308 B.n307 163.367
R957 B.n304 B.n303 163.367
R958 B.n300 B.n299 163.367
R959 B.n296 B.n295 163.367
R960 B.n292 B.n291 163.367
R961 B.n288 B.n287 163.367
R962 B.n284 B.n283 163.367
R963 B.n280 B.n279 163.367
R964 B.n276 B.n275 163.367
R965 B.n404 B.n236 163.367
R966 B.n410 B.n232 163.367
R967 B.n410 B.n230 163.367
R968 B.n414 B.n230 163.367
R969 B.n414 B.n224 163.367
R970 B.n422 B.n224 163.367
R971 B.n422 B.n222 163.367
R972 B.n426 B.n222 163.367
R973 B.n426 B.n216 163.367
R974 B.n434 B.n216 163.367
R975 B.n434 B.n214 163.367
R976 B.n438 B.n214 163.367
R977 B.n438 B.n208 163.367
R978 B.n448 B.n208 163.367
R979 B.n448 B.n206 163.367
R980 B.n452 B.n206 163.367
R981 B.n452 B.n3 163.367
R982 B.n520 B.n3 163.367
R983 B.n516 B.n2 163.367
R984 B.n516 B.n515 163.367
R985 B.n515 B.n9 163.367
R986 B.n511 B.n9 163.367
R987 B.n511 B.n11 163.367
R988 B.n507 B.n11 163.367
R989 B.n507 B.n17 163.367
R990 B.n503 B.n17 163.367
R991 B.n503 B.n19 163.367
R992 B.n499 B.n19 163.367
R993 B.n499 B.n24 163.367
R994 B.n495 B.n24 163.367
R995 B.n495 B.n26 163.367
R996 B.n491 B.n26 163.367
R997 B.n491 B.n31 163.367
R998 B.n487 B.n31 163.367
R999 B.n487 B.n33 163.367
R1000 B.n403 B.n233 99.961
R1001 B.n485 B.n484 99.961
R1002 B.n75 B.n36 71.676
R1003 B.n79 B.n37 71.676
R1004 B.n83 B.n38 71.676
R1005 B.n87 B.n39 71.676
R1006 B.n91 B.n40 71.676
R1007 B.n95 B.n41 71.676
R1008 B.n99 B.n42 71.676
R1009 B.n103 B.n43 71.676
R1010 B.n107 B.n44 71.676
R1011 B.n111 B.n45 71.676
R1012 B.n115 B.n46 71.676
R1013 B.n119 B.n47 71.676
R1014 B.n123 B.n48 71.676
R1015 B.n127 B.n49 71.676
R1016 B.n131 B.n50 71.676
R1017 B.n135 B.n51 71.676
R1018 B.n139 B.n52 71.676
R1019 B.n143 B.n53 71.676
R1020 B.n147 B.n54 71.676
R1021 B.n151 B.n55 71.676
R1022 B.n155 B.n56 71.676
R1023 B.n159 B.n57 71.676
R1024 B.n163 B.n58 71.676
R1025 B.n167 B.n59 71.676
R1026 B.n171 B.n60 71.676
R1027 B.n175 B.n61 71.676
R1028 B.n179 B.n62 71.676
R1029 B.n183 B.n63 71.676
R1030 B.n187 B.n64 71.676
R1031 B.n191 B.n65 71.676
R1032 B.n195 B.n66 71.676
R1033 B.n199 B.n67 71.676
R1034 B.n483 B.n68 71.676
R1035 B.n483 B.n482 71.676
R1036 B.n201 B.n67 71.676
R1037 B.n198 B.n66 71.676
R1038 B.n194 B.n65 71.676
R1039 B.n190 B.n64 71.676
R1040 B.n186 B.n63 71.676
R1041 B.n182 B.n62 71.676
R1042 B.n178 B.n61 71.676
R1043 B.n174 B.n60 71.676
R1044 B.n170 B.n59 71.676
R1045 B.n166 B.n58 71.676
R1046 B.n162 B.n57 71.676
R1047 B.n158 B.n56 71.676
R1048 B.n154 B.n55 71.676
R1049 B.n150 B.n54 71.676
R1050 B.n146 B.n53 71.676
R1051 B.n142 B.n52 71.676
R1052 B.n138 B.n51 71.676
R1053 B.n134 B.n50 71.676
R1054 B.n130 B.n49 71.676
R1055 B.n126 B.n48 71.676
R1056 B.n122 B.n47 71.676
R1057 B.n118 B.n46 71.676
R1058 B.n114 B.n45 71.676
R1059 B.n110 B.n44 71.676
R1060 B.n106 B.n43 71.676
R1061 B.n102 B.n42 71.676
R1062 B.n98 B.n41 71.676
R1063 B.n94 B.n40 71.676
R1064 B.n90 B.n39 71.676
R1065 B.n86 B.n38 71.676
R1066 B.n82 B.n37 71.676
R1067 B.n78 B.n36 71.676
R1068 B.n402 B.n401 71.676
R1069 B.n396 B.n237 71.676
R1070 B.n393 B.n238 71.676
R1071 B.n389 B.n239 71.676
R1072 B.n385 B.n240 71.676
R1073 B.n381 B.n241 71.676
R1074 B.n377 B.n242 71.676
R1075 B.n373 B.n243 71.676
R1076 B.n369 B.n244 71.676
R1077 B.n365 B.n245 71.676
R1078 B.n361 B.n246 71.676
R1079 B.n357 B.n247 71.676
R1080 B.n353 B.n248 71.676
R1081 B.n349 B.n249 71.676
R1082 B.n344 B.n250 71.676
R1083 B.n340 B.n251 71.676
R1084 B.n336 B.n252 71.676
R1085 B.n332 B.n253 71.676
R1086 B.n328 B.n254 71.676
R1087 B.n323 B.n255 71.676
R1088 B.n319 B.n256 71.676
R1089 B.n315 B.n257 71.676
R1090 B.n311 B.n258 71.676
R1091 B.n307 B.n259 71.676
R1092 B.n303 B.n260 71.676
R1093 B.n299 B.n261 71.676
R1094 B.n295 B.n262 71.676
R1095 B.n291 B.n263 71.676
R1096 B.n287 B.n264 71.676
R1097 B.n283 B.n265 71.676
R1098 B.n279 B.n266 71.676
R1099 B.n275 B.n267 71.676
R1100 B.n402 B.n269 71.676
R1101 B.n394 B.n237 71.676
R1102 B.n390 B.n238 71.676
R1103 B.n386 B.n239 71.676
R1104 B.n382 B.n240 71.676
R1105 B.n378 B.n241 71.676
R1106 B.n374 B.n242 71.676
R1107 B.n370 B.n243 71.676
R1108 B.n366 B.n244 71.676
R1109 B.n362 B.n245 71.676
R1110 B.n358 B.n246 71.676
R1111 B.n354 B.n247 71.676
R1112 B.n350 B.n248 71.676
R1113 B.n345 B.n249 71.676
R1114 B.n341 B.n250 71.676
R1115 B.n337 B.n251 71.676
R1116 B.n333 B.n252 71.676
R1117 B.n329 B.n253 71.676
R1118 B.n324 B.n254 71.676
R1119 B.n320 B.n255 71.676
R1120 B.n316 B.n256 71.676
R1121 B.n312 B.n257 71.676
R1122 B.n308 B.n258 71.676
R1123 B.n304 B.n259 71.676
R1124 B.n300 B.n260 71.676
R1125 B.n296 B.n261 71.676
R1126 B.n292 B.n262 71.676
R1127 B.n288 B.n263 71.676
R1128 B.n284 B.n264 71.676
R1129 B.n280 B.n265 71.676
R1130 B.n276 B.n266 71.676
R1131 B.n267 B.n236 71.676
R1132 B.n521 B.n520 71.676
R1133 B.n521 B.n2 71.676
R1134 B.n74 B.n73 59.5399
R1135 B.n71 B.n70 59.5399
R1136 B.n326 B.n273 59.5399
R1137 B.n347 B.n271 59.5399
R1138 B.n409 B.n233 59.1076
R1139 B.n409 B.n228 59.1076
R1140 B.n415 B.n228 59.1076
R1141 B.n415 B.n229 59.1076
R1142 B.n421 B.n221 59.1076
R1143 B.n427 B.n221 59.1076
R1144 B.n427 B.n217 59.1076
R1145 B.n433 B.n217 59.1076
R1146 B.n433 B.n213 59.1076
R1147 B.n439 B.n213 59.1076
R1148 B.n447 B.n209 59.1076
R1149 B.n447 B.n446 59.1076
R1150 B.n453 B.n4 59.1076
R1151 B.n519 B.n4 59.1076
R1152 B.n519 B.n518 59.1076
R1153 B.n518 B.n517 59.1076
R1154 B.n517 B.n8 59.1076
R1155 B.n510 B.n12 59.1076
R1156 B.n510 B.n509 59.1076
R1157 B.n508 B.n16 59.1076
R1158 B.n502 B.n16 59.1076
R1159 B.n502 B.n501 59.1076
R1160 B.n501 B.n500 59.1076
R1161 B.n500 B.n23 59.1076
R1162 B.n494 B.n23 59.1076
R1163 B.n493 B.n492 59.1076
R1164 B.n492 B.n30 59.1076
R1165 B.n486 B.n30 59.1076
R1166 B.n486 B.n485 59.1076
R1167 B.n229 B.t9 57.3691
R1168 B.t5 B.n493 57.3691
R1169 B.t2 B.n209 43.4616
R1170 B.n509 B.t0 43.4616
R1171 B.n453 B.t3 38.2463
R1172 B.t1 B.n8 38.2463
R1173 B.n400 B.n231 29.1907
R1174 B.n406 B.n405 29.1907
R1175 B.n481 B.n480 29.1907
R1176 B.n76 B.n32 29.1907
R1177 B.n446 B.t3 20.8618
R1178 B.n12 B.t1 20.8618
R1179 B.n73 B.n72 20.3641
R1180 B.n70 B.n69 20.3641
R1181 B.n273 B.n272 20.3641
R1182 B.n271 B.n270 20.3641
R1183 B B.n522 18.0485
R1184 B.n439 B.t2 15.6465
R1185 B.t0 B.n508 15.6465
R1186 B.n411 B.n231 10.6151
R1187 B.n412 B.n411 10.6151
R1188 B.n413 B.n412 10.6151
R1189 B.n413 B.n223 10.6151
R1190 B.n423 B.n223 10.6151
R1191 B.n424 B.n423 10.6151
R1192 B.n425 B.n424 10.6151
R1193 B.n425 B.n215 10.6151
R1194 B.n435 B.n215 10.6151
R1195 B.n436 B.n435 10.6151
R1196 B.n437 B.n436 10.6151
R1197 B.n437 B.n207 10.6151
R1198 B.n449 B.n207 10.6151
R1199 B.n450 B.n449 10.6151
R1200 B.n451 B.n450 10.6151
R1201 B.n451 B.n0 10.6151
R1202 B.n400 B.n399 10.6151
R1203 B.n399 B.n398 10.6151
R1204 B.n398 B.n397 10.6151
R1205 B.n397 B.n395 10.6151
R1206 B.n395 B.n392 10.6151
R1207 B.n392 B.n391 10.6151
R1208 B.n391 B.n388 10.6151
R1209 B.n388 B.n387 10.6151
R1210 B.n387 B.n384 10.6151
R1211 B.n384 B.n383 10.6151
R1212 B.n383 B.n380 10.6151
R1213 B.n380 B.n379 10.6151
R1214 B.n379 B.n376 10.6151
R1215 B.n376 B.n375 10.6151
R1216 B.n375 B.n372 10.6151
R1217 B.n372 B.n371 10.6151
R1218 B.n371 B.n368 10.6151
R1219 B.n368 B.n367 10.6151
R1220 B.n367 B.n364 10.6151
R1221 B.n364 B.n363 10.6151
R1222 B.n363 B.n360 10.6151
R1223 B.n360 B.n359 10.6151
R1224 B.n359 B.n356 10.6151
R1225 B.n356 B.n355 10.6151
R1226 B.n355 B.n352 10.6151
R1227 B.n352 B.n351 10.6151
R1228 B.n351 B.n348 10.6151
R1229 B.n346 B.n343 10.6151
R1230 B.n343 B.n342 10.6151
R1231 B.n342 B.n339 10.6151
R1232 B.n339 B.n338 10.6151
R1233 B.n338 B.n335 10.6151
R1234 B.n335 B.n334 10.6151
R1235 B.n334 B.n331 10.6151
R1236 B.n331 B.n330 10.6151
R1237 B.n330 B.n327 10.6151
R1238 B.n325 B.n322 10.6151
R1239 B.n322 B.n321 10.6151
R1240 B.n321 B.n318 10.6151
R1241 B.n318 B.n317 10.6151
R1242 B.n317 B.n314 10.6151
R1243 B.n314 B.n313 10.6151
R1244 B.n313 B.n310 10.6151
R1245 B.n310 B.n309 10.6151
R1246 B.n309 B.n306 10.6151
R1247 B.n306 B.n305 10.6151
R1248 B.n305 B.n302 10.6151
R1249 B.n302 B.n301 10.6151
R1250 B.n301 B.n298 10.6151
R1251 B.n298 B.n297 10.6151
R1252 B.n297 B.n294 10.6151
R1253 B.n294 B.n293 10.6151
R1254 B.n293 B.n290 10.6151
R1255 B.n290 B.n289 10.6151
R1256 B.n289 B.n286 10.6151
R1257 B.n286 B.n285 10.6151
R1258 B.n285 B.n282 10.6151
R1259 B.n282 B.n281 10.6151
R1260 B.n281 B.n278 10.6151
R1261 B.n278 B.n277 10.6151
R1262 B.n277 B.n274 10.6151
R1263 B.n274 B.n235 10.6151
R1264 B.n405 B.n235 10.6151
R1265 B.n407 B.n406 10.6151
R1266 B.n407 B.n226 10.6151
R1267 B.n417 B.n226 10.6151
R1268 B.n418 B.n417 10.6151
R1269 B.n419 B.n418 10.6151
R1270 B.n419 B.n219 10.6151
R1271 B.n429 B.n219 10.6151
R1272 B.n430 B.n429 10.6151
R1273 B.n431 B.n430 10.6151
R1274 B.n431 B.n211 10.6151
R1275 B.n441 B.n211 10.6151
R1276 B.n442 B.n441 10.6151
R1277 B.n444 B.n442 10.6151
R1278 B.n444 B.n443 10.6151
R1279 B.n443 B.n204 10.6151
R1280 B.n456 B.n204 10.6151
R1281 B.n457 B.n456 10.6151
R1282 B.n458 B.n457 10.6151
R1283 B.n459 B.n458 10.6151
R1284 B.n460 B.n459 10.6151
R1285 B.n463 B.n460 10.6151
R1286 B.n464 B.n463 10.6151
R1287 B.n465 B.n464 10.6151
R1288 B.n466 B.n465 10.6151
R1289 B.n468 B.n466 10.6151
R1290 B.n469 B.n468 10.6151
R1291 B.n470 B.n469 10.6151
R1292 B.n471 B.n470 10.6151
R1293 B.n473 B.n471 10.6151
R1294 B.n474 B.n473 10.6151
R1295 B.n475 B.n474 10.6151
R1296 B.n476 B.n475 10.6151
R1297 B.n478 B.n476 10.6151
R1298 B.n479 B.n478 10.6151
R1299 B.n480 B.n479 10.6151
R1300 B.n514 B.n1 10.6151
R1301 B.n514 B.n513 10.6151
R1302 B.n513 B.n512 10.6151
R1303 B.n512 B.n10 10.6151
R1304 B.n506 B.n10 10.6151
R1305 B.n506 B.n505 10.6151
R1306 B.n505 B.n504 10.6151
R1307 B.n504 B.n18 10.6151
R1308 B.n498 B.n18 10.6151
R1309 B.n498 B.n497 10.6151
R1310 B.n497 B.n496 10.6151
R1311 B.n496 B.n25 10.6151
R1312 B.n490 B.n25 10.6151
R1313 B.n490 B.n489 10.6151
R1314 B.n489 B.n488 10.6151
R1315 B.n488 B.n32 10.6151
R1316 B.n77 B.n76 10.6151
R1317 B.n80 B.n77 10.6151
R1318 B.n81 B.n80 10.6151
R1319 B.n84 B.n81 10.6151
R1320 B.n85 B.n84 10.6151
R1321 B.n88 B.n85 10.6151
R1322 B.n89 B.n88 10.6151
R1323 B.n92 B.n89 10.6151
R1324 B.n93 B.n92 10.6151
R1325 B.n96 B.n93 10.6151
R1326 B.n97 B.n96 10.6151
R1327 B.n100 B.n97 10.6151
R1328 B.n101 B.n100 10.6151
R1329 B.n104 B.n101 10.6151
R1330 B.n105 B.n104 10.6151
R1331 B.n108 B.n105 10.6151
R1332 B.n109 B.n108 10.6151
R1333 B.n112 B.n109 10.6151
R1334 B.n113 B.n112 10.6151
R1335 B.n116 B.n113 10.6151
R1336 B.n117 B.n116 10.6151
R1337 B.n120 B.n117 10.6151
R1338 B.n121 B.n120 10.6151
R1339 B.n124 B.n121 10.6151
R1340 B.n125 B.n124 10.6151
R1341 B.n128 B.n125 10.6151
R1342 B.n129 B.n128 10.6151
R1343 B.n133 B.n132 10.6151
R1344 B.n136 B.n133 10.6151
R1345 B.n137 B.n136 10.6151
R1346 B.n140 B.n137 10.6151
R1347 B.n141 B.n140 10.6151
R1348 B.n144 B.n141 10.6151
R1349 B.n145 B.n144 10.6151
R1350 B.n148 B.n145 10.6151
R1351 B.n149 B.n148 10.6151
R1352 B.n153 B.n152 10.6151
R1353 B.n156 B.n153 10.6151
R1354 B.n157 B.n156 10.6151
R1355 B.n160 B.n157 10.6151
R1356 B.n161 B.n160 10.6151
R1357 B.n164 B.n161 10.6151
R1358 B.n165 B.n164 10.6151
R1359 B.n168 B.n165 10.6151
R1360 B.n169 B.n168 10.6151
R1361 B.n172 B.n169 10.6151
R1362 B.n173 B.n172 10.6151
R1363 B.n176 B.n173 10.6151
R1364 B.n177 B.n176 10.6151
R1365 B.n180 B.n177 10.6151
R1366 B.n181 B.n180 10.6151
R1367 B.n184 B.n181 10.6151
R1368 B.n185 B.n184 10.6151
R1369 B.n188 B.n185 10.6151
R1370 B.n189 B.n188 10.6151
R1371 B.n192 B.n189 10.6151
R1372 B.n193 B.n192 10.6151
R1373 B.n196 B.n193 10.6151
R1374 B.n197 B.n196 10.6151
R1375 B.n200 B.n197 10.6151
R1376 B.n202 B.n200 10.6151
R1377 B.n203 B.n202 10.6151
R1378 B.n481 B.n203 10.6151
R1379 B.n348 B.n347 9.36635
R1380 B.n326 B.n325 9.36635
R1381 B.n129 B.n74 9.36635
R1382 B.n152 B.n71 9.36635
R1383 B.n522 B.n0 8.11757
R1384 B.n522 B.n1 8.11757
R1385 B.n421 B.t9 1.73894
R1386 B.n494 B.t5 1.73894
R1387 B.n347 B.n346 1.24928
R1388 B.n327 B.n326 1.24928
R1389 B.n132 B.n74 1.24928
R1390 B.n149 B.n71 1.24928
R1391 VN.n0 VN.t3 322.582
R1392 VN.n1 VN.t1 322.582
R1393 VN.n0 VN.t0 322.531
R1394 VN.n1 VN.t2 322.531
R1395 VN VN.n1 82.0276
R1396 VN VN.n0 44.7132
R1397 VDD2.n2 VDD2.n0 96.8291
R1398 VDD2.n2 VDD2.n1 64.0367
R1399 VDD2.n1 VDD2.t1 2.68343
R1400 VDD2.n1 VDD2.t2 2.68343
R1401 VDD2.n0 VDD2.t0 2.68343
R1402 VDD2.n0 VDD2.t3 2.68343
R1403 VDD2 VDD2.n2 0.0586897
C0 VTAIL VN 1.87381f
C1 VDD1 VTAIL 4.70313f
C2 VDD2 VP 0.274818f
C3 VP VN 3.97974f
C4 VP VDD1 2.20618f
C5 VDD2 VN 2.07906f
C6 VP VTAIL 1.88792f
C7 VDD2 VDD1 0.571013f
C8 VDD1 VN 0.147441f
C9 VDD2 VTAIL 4.74473f
C10 VDD2 B 2.348435f
C11 VDD1 B 5.44409f
C12 VTAIL B 6.171957f
C13 VN B 6.85029f
C14 VP B 4.623044f
C15 VDD2.t0 B 0.162103f
C16 VDD2.t3 B 0.162103f
C17 VDD2.n0 B 1.82215f
C18 VDD2.t1 B 0.162103f
C19 VDD2.t2 B 0.162103f
C20 VDD2.n1 B 1.38248f
C21 VDD2.n2 B 2.8599f
C22 VN.t3 B 0.59659f
C23 VN.t0 B 0.596544f
C24 VN.n0 B 0.478131f
C25 VN.t1 B 0.59659f
C26 VN.t2 B 0.596544f
C27 VN.n1 B 1.097f
C28 VDD1.t0 B 0.162041f
C29 VDD1.t3 B 0.162041f
C30 VDD1.n0 B 1.38225f
C31 VDD1.t2 B 0.162041f
C32 VDD1.t1 B 0.162041f
C33 VDD1.n1 B 1.84556f
C34 VTAIL.n0 B 0.017597f
C35 VTAIL.n1 B 0.0124f
C36 VTAIL.n2 B 0.006663f
C37 VTAIL.n3 B 0.01575f
C38 VTAIL.n4 B 0.007055f
C39 VTAIL.n5 B 0.0124f
C40 VTAIL.n6 B 0.006663f
C41 VTAIL.n7 B 0.01575f
C42 VTAIL.n8 B 0.007055f
C43 VTAIL.n9 B 0.0124f
C44 VTAIL.n10 B 0.006663f
C45 VTAIL.n11 B 0.011812f
C46 VTAIL.n12 B 0.009304f
C47 VTAIL.t1 B 0.025667f
C48 VTAIL.n13 B 0.057231f
C49 VTAIL.n14 B 0.373666f
C50 VTAIL.n15 B 0.006663f
C51 VTAIL.n16 B 0.007055f
C52 VTAIL.n17 B 0.01575f
C53 VTAIL.n18 B 0.01575f
C54 VTAIL.n19 B 0.007055f
C55 VTAIL.n20 B 0.006663f
C56 VTAIL.n21 B 0.0124f
C57 VTAIL.n22 B 0.0124f
C58 VTAIL.n23 B 0.006663f
C59 VTAIL.n24 B 0.007055f
C60 VTAIL.n25 B 0.01575f
C61 VTAIL.n26 B 0.01575f
C62 VTAIL.n27 B 0.007055f
C63 VTAIL.n28 B 0.006663f
C64 VTAIL.n29 B 0.0124f
C65 VTAIL.n30 B 0.0124f
C66 VTAIL.n31 B 0.006663f
C67 VTAIL.n32 B 0.007055f
C68 VTAIL.n33 B 0.01575f
C69 VTAIL.n34 B 0.034392f
C70 VTAIL.n35 B 0.007055f
C71 VTAIL.n36 B 0.006663f
C72 VTAIL.n37 B 0.027646f
C73 VTAIL.n38 B 0.019242f
C74 VTAIL.n39 B 0.049199f
C75 VTAIL.n40 B 0.017597f
C76 VTAIL.n41 B 0.0124f
C77 VTAIL.n42 B 0.006663f
C78 VTAIL.n43 B 0.01575f
C79 VTAIL.n44 B 0.007055f
C80 VTAIL.n45 B 0.0124f
C81 VTAIL.n46 B 0.006663f
C82 VTAIL.n47 B 0.01575f
C83 VTAIL.n48 B 0.007055f
C84 VTAIL.n49 B 0.0124f
C85 VTAIL.n50 B 0.006663f
C86 VTAIL.n51 B 0.011812f
C87 VTAIL.n52 B 0.009304f
C88 VTAIL.t4 B 0.025667f
C89 VTAIL.n53 B 0.057231f
C90 VTAIL.n54 B 0.373666f
C91 VTAIL.n55 B 0.006663f
C92 VTAIL.n56 B 0.007055f
C93 VTAIL.n57 B 0.01575f
C94 VTAIL.n58 B 0.01575f
C95 VTAIL.n59 B 0.007055f
C96 VTAIL.n60 B 0.006663f
C97 VTAIL.n61 B 0.0124f
C98 VTAIL.n62 B 0.0124f
C99 VTAIL.n63 B 0.006663f
C100 VTAIL.n64 B 0.007055f
C101 VTAIL.n65 B 0.01575f
C102 VTAIL.n66 B 0.01575f
C103 VTAIL.n67 B 0.007055f
C104 VTAIL.n68 B 0.006663f
C105 VTAIL.n69 B 0.0124f
C106 VTAIL.n70 B 0.0124f
C107 VTAIL.n71 B 0.006663f
C108 VTAIL.n72 B 0.007055f
C109 VTAIL.n73 B 0.01575f
C110 VTAIL.n74 B 0.034392f
C111 VTAIL.n75 B 0.007055f
C112 VTAIL.n76 B 0.006663f
C113 VTAIL.n77 B 0.027646f
C114 VTAIL.n78 B 0.019242f
C115 VTAIL.n79 B 0.064958f
C116 VTAIL.n80 B 0.017597f
C117 VTAIL.n81 B 0.0124f
C118 VTAIL.n82 B 0.006663f
C119 VTAIL.n83 B 0.01575f
C120 VTAIL.n84 B 0.007055f
C121 VTAIL.n85 B 0.0124f
C122 VTAIL.n86 B 0.006663f
C123 VTAIL.n87 B 0.01575f
C124 VTAIL.n88 B 0.007055f
C125 VTAIL.n89 B 0.0124f
C126 VTAIL.n90 B 0.006663f
C127 VTAIL.n91 B 0.011812f
C128 VTAIL.n92 B 0.009304f
C129 VTAIL.t7 B 0.025667f
C130 VTAIL.n93 B 0.057231f
C131 VTAIL.n94 B 0.373666f
C132 VTAIL.n95 B 0.006663f
C133 VTAIL.n96 B 0.007055f
C134 VTAIL.n97 B 0.01575f
C135 VTAIL.n98 B 0.01575f
C136 VTAIL.n99 B 0.007055f
C137 VTAIL.n100 B 0.006663f
C138 VTAIL.n101 B 0.0124f
C139 VTAIL.n102 B 0.0124f
C140 VTAIL.n103 B 0.006663f
C141 VTAIL.n104 B 0.007055f
C142 VTAIL.n105 B 0.01575f
C143 VTAIL.n106 B 0.01575f
C144 VTAIL.n107 B 0.007055f
C145 VTAIL.n108 B 0.006663f
C146 VTAIL.n109 B 0.0124f
C147 VTAIL.n110 B 0.0124f
C148 VTAIL.n111 B 0.006663f
C149 VTAIL.n112 B 0.007055f
C150 VTAIL.n113 B 0.01575f
C151 VTAIL.n114 B 0.034392f
C152 VTAIL.n115 B 0.007055f
C153 VTAIL.n116 B 0.006663f
C154 VTAIL.n117 B 0.027646f
C155 VTAIL.n118 B 0.019242f
C156 VTAIL.n119 B 0.505002f
C157 VTAIL.n120 B 0.017597f
C158 VTAIL.n121 B 0.0124f
C159 VTAIL.n122 B 0.006663f
C160 VTAIL.n123 B 0.01575f
C161 VTAIL.n124 B 0.007055f
C162 VTAIL.n125 B 0.0124f
C163 VTAIL.n126 B 0.006663f
C164 VTAIL.n127 B 0.01575f
C165 VTAIL.n128 B 0.007055f
C166 VTAIL.n129 B 0.0124f
C167 VTAIL.n130 B 0.006663f
C168 VTAIL.n131 B 0.011812f
C169 VTAIL.n132 B 0.009304f
C170 VTAIL.t2 B 0.025667f
C171 VTAIL.n133 B 0.057231f
C172 VTAIL.n134 B 0.373666f
C173 VTAIL.n135 B 0.006663f
C174 VTAIL.n136 B 0.007055f
C175 VTAIL.n137 B 0.01575f
C176 VTAIL.n138 B 0.01575f
C177 VTAIL.n139 B 0.007055f
C178 VTAIL.n140 B 0.006663f
C179 VTAIL.n141 B 0.0124f
C180 VTAIL.n142 B 0.0124f
C181 VTAIL.n143 B 0.006663f
C182 VTAIL.n144 B 0.007055f
C183 VTAIL.n145 B 0.01575f
C184 VTAIL.n146 B 0.01575f
C185 VTAIL.n147 B 0.007055f
C186 VTAIL.n148 B 0.006663f
C187 VTAIL.n149 B 0.0124f
C188 VTAIL.n150 B 0.0124f
C189 VTAIL.n151 B 0.006663f
C190 VTAIL.n152 B 0.007055f
C191 VTAIL.n153 B 0.01575f
C192 VTAIL.n154 B 0.034392f
C193 VTAIL.n155 B 0.007055f
C194 VTAIL.n156 B 0.006663f
C195 VTAIL.n157 B 0.027646f
C196 VTAIL.n158 B 0.019242f
C197 VTAIL.n159 B 0.505002f
C198 VTAIL.n160 B 0.017597f
C199 VTAIL.n161 B 0.0124f
C200 VTAIL.n162 B 0.006663f
C201 VTAIL.n163 B 0.01575f
C202 VTAIL.n164 B 0.007055f
C203 VTAIL.n165 B 0.0124f
C204 VTAIL.n166 B 0.006663f
C205 VTAIL.n167 B 0.01575f
C206 VTAIL.n168 B 0.007055f
C207 VTAIL.n169 B 0.0124f
C208 VTAIL.n170 B 0.006663f
C209 VTAIL.n171 B 0.011812f
C210 VTAIL.n172 B 0.009304f
C211 VTAIL.t3 B 0.025667f
C212 VTAIL.n173 B 0.057231f
C213 VTAIL.n174 B 0.373666f
C214 VTAIL.n175 B 0.006663f
C215 VTAIL.n176 B 0.007055f
C216 VTAIL.n177 B 0.01575f
C217 VTAIL.n178 B 0.01575f
C218 VTAIL.n179 B 0.007055f
C219 VTAIL.n180 B 0.006663f
C220 VTAIL.n181 B 0.0124f
C221 VTAIL.n182 B 0.0124f
C222 VTAIL.n183 B 0.006663f
C223 VTAIL.n184 B 0.007055f
C224 VTAIL.n185 B 0.01575f
C225 VTAIL.n186 B 0.01575f
C226 VTAIL.n187 B 0.007055f
C227 VTAIL.n188 B 0.006663f
C228 VTAIL.n189 B 0.0124f
C229 VTAIL.n190 B 0.0124f
C230 VTAIL.n191 B 0.006663f
C231 VTAIL.n192 B 0.007055f
C232 VTAIL.n193 B 0.01575f
C233 VTAIL.n194 B 0.034392f
C234 VTAIL.n195 B 0.007055f
C235 VTAIL.n196 B 0.006663f
C236 VTAIL.n197 B 0.027646f
C237 VTAIL.n198 B 0.019242f
C238 VTAIL.n199 B 0.064958f
C239 VTAIL.n200 B 0.017597f
C240 VTAIL.n201 B 0.0124f
C241 VTAIL.n202 B 0.006663f
C242 VTAIL.n203 B 0.01575f
C243 VTAIL.n204 B 0.007055f
C244 VTAIL.n205 B 0.0124f
C245 VTAIL.n206 B 0.006663f
C246 VTAIL.n207 B 0.01575f
C247 VTAIL.n208 B 0.007055f
C248 VTAIL.n209 B 0.0124f
C249 VTAIL.n210 B 0.006663f
C250 VTAIL.n211 B 0.011812f
C251 VTAIL.n212 B 0.009304f
C252 VTAIL.t6 B 0.025667f
C253 VTAIL.n213 B 0.057231f
C254 VTAIL.n214 B 0.373666f
C255 VTAIL.n215 B 0.006663f
C256 VTAIL.n216 B 0.007055f
C257 VTAIL.n217 B 0.01575f
C258 VTAIL.n218 B 0.01575f
C259 VTAIL.n219 B 0.007055f
C260 VTAIL.n220 B 0.006663f
C261 VTAIL.n221 B 0.0124f
C262 VTAIL.n222 B 0.0124f
C263 VTAIL.n223 B 0.006663f
C264 VTAIL.n224 B 0.007055f
C265 VTAIL.n225 B 0.01575f
C266 VTAIL.n226 B 0.01575f
C267 VTAIL.n227 B 0.007055f
C268 VTAIL.n228 B 0.006663f
C269 VTAIL.n229 B 0.0124f
C270 VTAIL.n230 B 0.0124f
C271 VTAIL.n231 B 0.006663f
C272 VTAIL.n232 B 0.007055f
C273 VTAIL.n233 B 0.01575f
C274 VTAIL.n234 B 0.034392f
C275 VTAIL.n235 B 0.007055f
C276 VTAIL.n236 B 0.006663f
C277 VTAIL.n237 B 0.027646f
C278 VTAIL.n238 B 0.019242f
C279 VTAIL.n239 B 0.064958f
C280 VTAIL.n240 B 0.017597f
C281 VTAIL.n241 B 0.0124f
C282 VTAIL.n242 B 0.006663f
C283 VTAIL.n243 B 0.01575f
C284 VTAIL.n244 B 0.007055f
C285 VTAIL.n245 B 0.0124f
C286 VTAIL.n246 B 0.006663f
C287 VTAIL.n247 B 0.01575f
C288 VTAIL.n248 B 0.007055f
C289 VTAIL.n249 B 0.0124f
C290 VTAIL.n250 B 0.006663f
C291 VTAIL.n251 B 0.011812f
C292 VTAIL.n252 B 0.009304f
C293 VTAIL.t5 B 0.025667f
C294 VTAIL.n253 B 0.057231f
C295 VTAIL.n254 B 0.373666f
C296 VTAIL.n255 B 0.006663f
C297 VTAIL.n256 B 0.007055f
C298 VTAIL.n257 B 0.01575f
C299 VTAIL.n258 B 0.01575f
C300 VTAIL.n259 B 0.007055f
C301 VTAIL.n260 B 0.006663f
C302 VTAIL.n261 B 0.0124f
C303 VTAIL.n262 B 0.0124f
C304 VTAIL.n263 B 0.006663f
C305 VTAIL.n264 B 0.007055f
C306 VTAIL.n265 B 0.01575f
C307 VTAIL.n266 B 0.01575f
C308 VTAIL.n267 B 0.007055f
C309 VTAIL.n268 B 0.006663f
C310 VTAIL.n269 B 0.0124f
C311 VTAIL.n270 B 0.0124f
C312 VTAIL.n271 B 0.006663f
C313 VTAIL.n272 B 0.007055f
C314 VTAIL.n273 B 0.01575f
C315 VTAIL.n274 B 0.034392f
C316 VTAIL.n275 B 0.007055f
C317 VTAIL.n276 B 0.006663f
C318 VTAIL.n277 B 0.027646f
C319 VTAIL.n278 B 0.019242f
C320 VTAIL.n279 B 0.505002f
C321 VTAIL.n280 B 0.017597f
C322 VTAIL.n281 B 0.0124f
C323 VTAIL.n282 B 0.006663f
C324 VTAIL.n283 B 0.01575f
C325 VTAIL.n284 B 0.007055f
C326 VTAIL.n285 B 0.0124f
C327 VTAIL.n286 B 0.006663f
C328 VTAIL.n287 B 0.01575f
C329 VTAIL.n288 B 0.007055f
C330 VTAIL.n289 B 0.0124f
C331 VTAIL.n290 B 0.006663f
C332 VTAIL.n291 B 0.011812f
C333 VTAIL.n292 B 0.009304f
C334 VTAIL.t0 B 0.025667f
C335 VTAIL.n293 B 0.057231f
C336 VTAIL.n294 B 0.373666f
C337 VTAIL.n295 B 0.006663f
C338 VTAIL.n296 B 0.007055f
C339 VTAIL.n297 B 0.01575f
C340 VTAIL.n298 B 0.01575f
C341 VTAIL.n299 B 0.007055f
C342 VTAIL.n300 B 0.006663f
C343 VTAIL.n301 B 0.0124f
C344 VTAIL.n302 B 0.0124f
C345 VTAIL.n303 B 0.006663f
C346 VTAIL.n304 B 0.007055f
C347 VTAIL.n305 B 0.01575f
C348 VTAIL.n306 B 0.01575f
C349 VTAIL.n307 B 0.007055f
C350 VTAIL.n308 B 0.006663f
C351 VTAIL.n309 B 0.0124f
C352 VTAIL.n310 B 0.0124f
C353 VTAIL.n311 B 0.006663f
C354 VTAIL.n312 B 0.007055f
C355 VTAIL.n313 B 0.01575f
C356 VTAIL.n314 B 0.034392f
C357 VTAIL.n315 B 0.007055f
C358 VTAIL.n316 B 0.006663f
C359 VTAIL.n317 B 0.027646f
C360 VTAIL.n318 B 0.019242f
C361 VTAIL.n319 B 0.484594f
C362 VP.n0 B 0.038835f
C363 VP.t0 B 0.611662f
C364 VP.t3 B 0.611709f
C365 VP.n1 B 1.10962f
C366 VP.n2 B 2.06965f
C367 VP.t1 B 0.594761f
C368 VP.n3 B 0.257446f
C369 VP.n4 B 0.008813f
C370 VP.t2 B 0.594761f
C371 VP.n5 B 0.257446f
C372 VP.n6 B 0.030096f
.ends

