* NGSPICE file created from diff_pair_sample_1612.ext - technology: sky130A

.subckt diff_pair_sample_1612 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t7 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=3.8
X1 VDD1.t4 VP.t1 VTAIL.t18 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=2.0553 pd=11.32 as=0.86955 ps=5.6 w=5.27 l=3.8
X2 B.t11 B.t9 B.t10 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=2.0553 pd=11.32 as=0 ps=0 w=5.27 l=3.8
X3 VTAIL.t9 VN.t0 VDD2.t9 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=3.8
X4 VTAIL.t17 VP.t2 VDD1.t8 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=3.8
X5 VDD2.t8 VN.t1 VTAIL.t0 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=2.0553 pd=11.32 as=0.86955 ps=5.6 w=5.27 l=3.8
X6 VDD1.t3 VP.t3 VTAIL.t16 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=3.8
X7 B.t8 B.t6 B.t7 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=2.0553 pd=11.32 as=0 ps=0 w=5.27 l=3.8
X8 VDD2.t7 VN.t2 VTAIL.t4 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=0.86955 pd=5.6 as=2.0553 ps=11.32 w=5.27 l=3.8
X9 VTAIL.t2 VN.t3 VDD2.t6 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=3.8
X10 B.t5 B.t3 B.t4 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=2.0553 pd=11.32 as=0 ps=0 w=5.27 l=3.8
X11 B.t2 B.t0 B.t1 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=2.0553 pd=11.32 as=0 ps=0 w=5.27 l=3.8
X12 VDD2.t5 VN.t4 VTAIL.t3 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=3.8
X13 VDD2.t4 VN.t5 VTAIL.t7 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=0.86955 pd=5.6 as=2.0553 ps=11.32 w=5.27 l=3.8
X14 VTAIL.t15 VP.t4 VDD1.t5 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=3.8
X15 VTAIL.t5 VN.t6 VDD2.t3 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=3.8
X16 VDD1.t2 VP.t5 VTAIL.t14 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=0.86955 pd=5.6 as=2.0553 ps=11.32 w=5.27 l=3.8
X17 VTAIL.t13 VP.t6 VDD1.t1 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=3.8
X18 VDD2.t2 VN.t7 VTAIL.t1 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=2.0553 pd=11.32 as=0.86955 ps=5.6 w=5.27 l=3.8
X19 VDD1.t6 VP.t7 VTAIL.t12 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=3.8
X20 VDD1.t0 VP.t8 VTAIL.t11 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=0.86955 pd=5.6 as=2.0553 ps=11.32 w=5.27 l=3.8
X21 VDD1.t9 VP.t9 VTAIL.t10 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=2.0553 pd=11.32 as=0.86955 ps=5.6 w=5.27 l=3.8
X22 VTAIL.t6 VN.t8 VDD2.t1 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=3.8
X23 VDD2.t0 VN.t9 VTAIL.t8 w_n5926_n2022# sky130_fd_pr__pfet_01v8 ad=0.86955 pd=5.6 as=0.86955 ps=5.6 w=5.27 l=3.8
R0 VP.n34 VP.n33 161.3
R1 VP.n35 VP.n30 161.3
R2 VP.n37 VP.n36 161.3
R3 VP.n38 VP.n29 161.3
R4 VP.n40 VP.n39 161.3
R5 VP.n41 VP.n28 161.3
R6 VP.n43 VP.n42 161.3
R7 VP.n44 VP.n27 161.3
R8 VP.n47 VP.n46 161.3
R9 VP.n48 VP.n26 161.3
R10 VP.n50 VP.n49 161.3
R11 VP.n51 VP.n25 161.3
R12 VP.n53 VP.n52 161.3
R13 VP.n54 VP.n24 161.3
R14 VP.n56 VP.n55 161.3
R15 VP.n57 VP.n23 161.3
R16 VP.n60 VP.n59 161.3
R17 VP.n61 VP.n22 161.3
R18 VP.n63 VP.n62 161.3
R19 VP.n64 VP.n21 161.3
R20 VP.n66 VP.n65 161.3
R21 VP.n67 VP.n20 161.3
R22 VP.n69 VP.n68 161.3
R23 VP.n70 VP.n19 161.3
R24 VP.n72 VP.n71 161.3
R25 VP.n129 VP.n128 161.3
R26 VP.n127 VP.n1 161.3
R27 VP.n126 VP.n125 161.3
R28 VP.n124 VP.n2 161.3
R29 VP.n123 VP.n122 161.3
R30 VP.n121 VP.n3 161.3
R31 VP.n120 VP.n119 161.3
R32 VP.n118 VP.n4 161.3
R33 VP.n117 VP.n116 161.3
R34 VP.n114 VP.n5 161.3
R35 VP.n113 VP.n112 161.3
R36 VP.n111 VP.n6 161.3
R37 VP.n110 VP.n109 161.3
R38 VP.n108 VP.n7 161.3
R39 VP.n107 VP.n106 161.3
R40 VP.n105 VP.n8 161.3
R41 VP.n104 VP.n103 161.3
R42 VP.n101 VP.n9 161.3
R43 VP.n100 VP.n99 161.3
R44 VP.n98 VP.n10 161.3
R45 VP.n97 VP.n96 161.3
R46 VP.n95 VP.n11 161.3
R47 VP.n94 VP.n93 161.3
R48 VP.n92 VP.n12 161.3
R49 VP.n91 VP.n90 161.3
R50 VP.n88 VP.n13 161.3
R51 VP.n87 VP.n86 161.3
R52 VP.n85 VP.n14 161.3
R53 VP.n84 VP.n83 161.3
R54 VP.n82 VP.n15 161.3
R55 VP.n81 VP.n80 161.3
R56 VP.n79 VP.n16 161.3
R57 VP.n78 VP.n77 161.3
R58 VP.n76 VP.n17 161.3
R59 VP.n75 VP.n74 89.5781
R60 VP.n130 VP.n0 89.5781
R61 VP.n73 VP.n18 89.5781
R62 VP.n31 VP.t9 65.6269
R63 VP.n96 VP.n95 56.5193
R64 VP.n109 VP.n108 56.5193
R65 VP.n52 VP.n51 56.5193
R66 VP.n39 VP.n38 56.5193
R67 VP.n32 VP.n31 56.4597
R68 VP.n74 VP.n73 54.5561
R69 VP.n83 VP.n82 45.8354
R70 VP.n122 VP.n121 45.8354
R71 VP.n65 VP.n64 45.8354
R72 VP.n82 VP.n81 35.1514
R73 VP.n122 VP.n2 35.1514
R74 VP.n65 VP.n20 35.1514
R75 VP.n75 VP.t1 33.4234
R76 VP.n89 VP.t2 33.4234
R77 VP.n102 VP.t3 33.4234
R78 VP.n115 VP.t6 33.4234
R79 VP.n0 VP.t5 33.4234
R80 VP.n18 VP.t8 33.4234
R81 VP.n58 VP.t4 33.4234
R82 VP.n45 VP.t7 33.4234
R83 VP.n32 VP.t0 33.4234
R84 VP.n77 VP.n76 24.4675
R85 VP.n77 VP.n16 24.4675
R86 VP.n81 VP.n16 24.4675
R87 VP.n83 VP.n14 24.4675
R88 VP.n87 VP.n14 24.4675
R89 VP.n88 VP.n87 24.4675
R90 VP.n90 VP.n12 24.4675
R91 VP.n94 VP.n12 24.4675
R92 VP.n95 VP.n94 24.4675
R93 VP.n96 VP.n10 24.4675
R94 VP.n100 VP.n10 24.4675
R95 VP.n101 VP.n100 24.4675
R96 VP.n103 VP.n8 24.4675
R97 VP.n107 VP.n8 24.4675
R98 VP.n108 VP.n107 24.4675
R99 VP.n109 VP.n6 24.4675
R100 VP.n113 VP.n6 24.4675
R101 VP.n114 VP.n113 24.4675
R102 VP.n116 VP.n4 24.4675
R103 VP.n120 VP.n4 24.4675
R104 VP.n121 VP.n120 24.4675
R105 VP.n126 VP.n2 24.4675
R106 VP.n127 VP.n126 24.4675
R107 VP.n128 VP.n127 24.4675
R108 VP.n69 VP.n20 24.4675
R109 VP.n70 VP.n69 24.4675
R110 VP.n71 VP.n70 24.4675
R111 VP.n52 VP.n24 24.4675
R112 VP.n56 VP.n24 24.4675
R113 VP.n57 VP.n56 24.4675
R114 VP.n59 VP.n22 24.4675
R115 VP.n63 VP.n22 24.4675
R116 VP.n64 VP.n63 24.4675
R117 VP.n39 VP.n28 24.4675
R118 VP.n43 VP.n28 24.4675
R119 VP.n44 VP.n43 24.4675
R120 VP.n46 VP.n26 24.4675
R121 VP.n50 VP.n26 24.4675
R122 VP.n51 VP.n50 24.4675
R123 VP.n33 VP.n30 24.4675
R124 VP.n37 VP.n30 24.4675
R125 VP.n38 VP.n37 24.4675
R126 VP.n90 VP.n89 18.5954
R127 VP.n115 VP.n114 18.5954
R128 VP.n58 VP.n57 18.5954
R129 VP.n33 VP.n32 18.5954
R130 VP.n102 VP.n101 12.234
R131 VP.n103 VP.n102 12.234
R132 VP.n45 VP.n44 12.234
R133 VP.n46 VP.n45 12.234
R134 VP.n89 VP.n88 5.87258
R135 VP.n116 VP.n115 5.87258
R136 VP.n59 VP.n58 5.87258
R137 VP.n34 VP.n31 2.51719
R138 VP.n76 VP.n75 0.48984
R139 VP.n128 VP.n0 0.48984
R140 VP.n71 VP.n18 0.48984
R141 VP.n73 VP.n72 0.354971
R142 VP.n74 VP.n17 0.354971
R143 VP.n130 VP.n129 0.354971
R144 VP VP.n130 0.26696
R145 VP.n35 VP.n34 0.189894
R146 VP.n36 VP.n35 0.189894
R147 VP.n36 VP.n29 0.189894
R148 VP.n40 VP.n29 0.189894
R149 VP.n41 VP.n40 0.189894
R150 VP.n42 VP.n41 0.189894
R151 VP.n42 VP.n27 0.189894
R152 VP.n47 VP.n27 0.189894
R153 VP.n48 VP.n47 0.189894
R154 VP.n49 VP.n48 0.189894
R155 VP.n49 VP.n25 0.189894
R156 VP.n53 VP.n25 0.189894
R157 VP.n54 VP.n53 0.189894
R158 VP.n55 VP.n54 0.189894
R159 VP.n55 VP.n23 0.189894
R160 VP.n60 VP.n23 0.189894
R161 VP.n61 VP.n60 0.189894
R162 VP.n62 VP.n61 0.189894
R163 VP.n62 VP.n21 0.189894
R164 VP.n66 VP.n21 0.189894
R165 VP.n67 VP.n66 0.189894
R166 VP.n68 VP.n67 0.189894
R167 VP.n68 VP.n19 0.189894
R168 VP.n72 VP.n19 0.189894
R169 VP.n78 VP.n17 0.189894
R170 VP.n79 VP.n78 0.189894
R171 VP.n80 VP.n79 0.189894
R172 VP.n80 VP.n15 0.189894
R173 VP.n84 VP.n15 0.189894
R174 VP.n85 VP.n84 0.189894
R175 VP.n86 VP.n85 0.189894
R176 VP.n86 VP.n13 0.189894
R177 VP.n91 VP.n13 0.189894
R178 VP.n92 VP.n91 0.189894
R179 VP.n93 VP.n92 0.189894
R180 VP.n93 VP.n11 0.189894
R181 VP.n97 VP.n11 0.189894
R182 VP.n98 VP.n97 0.189894
R183 VP.n99 VP.n98 0.189894
R184 VP.n99 VP.n9 0.189894
R185 VP.n104 VP.n9 0.189894
R186 VP.n105 VP.n104 0.189894
R187 VP.n106 VP.n105 0.189894
R188 VP.n106 VP.n7 0.189894
R189 VP.n110 VP.n7 0.189894
R190 VP.n111 VP.n110 0.189894
R191 VP.n112 VP.n111 0.189894
R192 VP.n112 VP.n5 0.189894
R193 VP.n117 VP.n5 0.189894
R194 VP.n118 VP.n117 0.189894
R195 VP.n119 VP.n118 0.189894
R196 VP.n119 VP.n3 0.189894
R197 VP.n123 VP.n3 0.189894
R198 VP.n124 VP.n123 0.189894
R199 VP.n125 VP.n124 0.189894
R200 VP.n125 VP.n1 0.189894
R201 VP.n129 VP.n1 0.189894
R202 VDD1.n22 VDD1.n0 756.745
R203 VDD1.n51 VDD1.n29 756.745
R204 VDD1.n23 VDD1.n22 585
R205 VDD1.n21 VDD1.n20 585
R206 VDD1.n4 VDD1.n3 585
R207 VDD1.n15 VDD1.n14 585
R208 VDD1.n13 VDD1.n12 585
R209 VDD1.n8 VDD1.n7 585
R210 VDD1.n37 VDD1.n36 585
R211 VDD1.n42 VDD1.n41 585
R212 VDD1.n44 VDD1.n43 585
R213 VDD1.n33 VDD1.n32 585
R214 VDD1.n50 VDD1.n49 585
R215 VDD1.n52 VDD1.n51 585
R216 VDD1.n9 VDD1.t9 327.856
R217 VDD1.n38 VDD1.t4 327.856
R218 VDD1.n22 VDD1.n21 171.744
R219 VDD1.n21 VDD1.n3 171.744
R220 VDD1.n14 VDD1.n3 171.744
R221 VDD1.n14 VDD1.n13 171.744
R222 VDD1.n13 VDD1.n7 171.744
R223 VDD1.n42 VDD1.n36 171.744
R224 VDD1.n43 VDD1.n42 171.744
R225 VDD1.n43 VDD1.n32 171.744
R226 VDD1.n50 VDD1.n32 171.744
R227 VDD1.n51 VDD1.n50 171.744
R228 VDD1.n59 VDD1.n58 99.7517
R229 VDD1.n28 VDD1.n27 97.137
R230 VDD1.n61 VDD1.n60 97.1368
R231 VDD1.n57 VDD1.n56 97.1368
R232 VDD1.t9 VDD1.n7 85.8723
R233 VDD1.t4 VDD1.n36 85.8723
R234 VDD1.n28 VDD1.n26 52.2305
R235 VDD1.n57 VDD1.n55 52.2305
R236 VDD1.n61 VDD1.n59 47.5332
R237 VDD1.n9 VDD1.n8 16.381
R238 VDD1.n38 VDD1.n37 16.381
R239 VDD1.n12 VDD1.n11 12.8005
R240 VDD1.n41 VDD1.n40 12.8005
R241 VDD1.n15 VDD1.n6 12.0247
R242 VDD1.n44 VDD1.n35 12.0247
R243 VDD1.n16 VDD1.n4 11.249
R244 VDD1.n45 VDD1.n33 11.249
R245 VDD1.n20 VDD1.n19 10.4732
R246 VDD1.n49 VDD1.n48 10.4732
R247 VDD1.n23 VDD1.n2 9.69747
R248 VDD1.n52 VDD1.n31 9.69747
R249 VDD1.n26 VDD1.n25 9.45567
R250 VDD1.n55 VDD1.n54 9.45567
R251 VDD1.n25 VDD1.n24 9.3005
R252 VDD1.n2 VDD1.n1 9.3005
R253 VDD1.n19 VDD1.n18 9.3005
R254 VDD1.n17 VDD1.n16 9.3005
R255 VDD1.n6 VDD1.n5 9.3005
R256 VDD1.n11 VDD1.n10 9.3005
R257 VDD1.n54 VDD1.n53 9.3005
R258 VDD1.n31 VDD1.n30 9.3005
R259 VDD1.n48 VDD1.n47 9.3005
R260 VDD1.n46 VDD1.n45 9.3005
R261 VDD1.n35 VDD1.n34 9.3005
R262 VDD1.n40 VDD1.n39 9.3005
R263 VDD1.n24 VDD1.n0 8.92171
R264 VDD1.n53 VDD1.n29 8.92171
R265 VDD1.n60 VDD1.t5 6.16843
R266 VDD1.n60 VDD1.t0 6.16843
R267 VDD1.n27 VDD1.t7 6.16843
R268 VDD1.n27 VDD1.t6 6.16843
R269 VDD1.n58 VDD1.t1 6.16843
R270 VDD1.n58 VDD1.t2 6.16843
R271 VDD1.n56 VDD1.t8 6.16843
R272 VDD1.n56 VDD1.t3 6.16843
R273 VDD1.n26 VDD1.n0 5.04292
R274 VDD1.n55 VDD1.n29 5.04292
R275 VDD1.n24 VDD1.n23 4.26717
R276 VDD1.n53 VDD1.n52 4.26717
R277 VDD1.n10 VDD1.n9 3.71853
R278 VDD1.n39 VDD1.n38 3.71853
R279 VDD1.n20 VDD1.n2 3.49141
R280 VDD1.n49 VDD1.n31 3.49141
R281 VDD1.n19 VDD1.n4 2.71565
R282 VDD1.n48 VDD1.n33 2.71565
R283 VDD1 VDD1.n61 2.61257
R284 VDD1.n16 VDD1.n15 1.93989
R285 VDD1.n45 VDD1.n44 1.93989
R286 VDD1.n12 VDD1.n6 1.16414
R287 VDD1.n41 VDD1.n35 1.16414
R288 VDD1 VDD1.n28 0.948776
R289 VDD1.n59 VDD1.n57 0.83524
R290 VDD1.n11 VDD1.n8 0.388379
R291 VDD1.n40 VDD1.n37 0.388379
R292 VDD1.n25 VDD1.n1 0.155672
R293 VDD1.n18 VDD1.n1 0.155672
R294 VDD1.n18 VDD1.n17 0.155672
R295 VDD1.n17 VDD1.n5 0.155672
R296 VDD1.n10 VDD1.n5 0.155672
R297 VDD1.n39 VDD1.n34 0.155672
R298 VDD1.n46 VDD1.n34 0.155672
R299 VDD1.n47 VDD1.n46 0.155672
R300 VDD1.n47 VDD1.n30 0.155672
R301 VDD1.n54 VDD1.n30 0.155672
R302 VTAIL.n120 VTAIL.n98 756.745
R303 VTAIL.n24 VTAIL.n2 756.745
R304 VTAIL.n92 VTAIL.n70 756.745
R305 VTAIL.n60 VTAIL.n38 756.745
R306 VTAIL.n106 VTAIL.n105 585
R307 VTAIL.n111 VTAIL.n110 585
R308 VTAIL.n113 VTAIL.n112 585
R309 VTAIL.n102 VTAIL.n101 585
R310 VTAIL.n119 VTAIL.n118 585
R311 VTAIL.n121 VTAIL.n120 585
R312 VTAIL.n10 VTAIL.n9 585
R313 VTAIL.n15 VTAIL.n14 585
R314 VTAIL.n17 VTAIL.n16 585
R315 VTAIL.n6 VTAIL.n5 585
R316 VTAIL.n23 VTAIL.n22 585
R317 VTAIL.n25 VTAIL.n24 585
R318 VTAIL.n93 VTAIL.n92 585
R319 VTAIL.n91 VTAIL.n90 585
R320 VTAIL.n74 VTAIL.n73 585
R321 VTAIL.n85 VTAIL.n84 585
R322 VTAIL.n83 VTAIL.n82 585
R323 VTAIL.n78 VTAIL.n77 585
R324 VTAIL.n61 VTAIL.n60 585
R325 VTAIL.n59 VTAIL.n58 585
R326 VTAIL.n42 VTAIL.n41 585
R327 VTAIL.n53 VTAIL.n52 585
R328 VTAIL.n51 VTAIL.n50 585
R329 VTAIL.n46 VTAIL.n45 585
R330 VTAIL.n107 VTAIL.t7 327.856
R331 VTAIL.n11 VTAIL.t14 327.856
R332 VTAIL.n79 VTAIL.t11 327.856
R333 VTAIL.n47 VTAIL.t4 327.856
R334 VTAIL.n111 VTAIL.n105 171.744
R335 VTAIL.n112 VTAIL.n111 171.744
R336 VTAIL.n112 VTAIL.n101 171.744
R337 VTAIL.n119 VTAIL.n101 171.744
R338 VTAIL.n120 VTAIL.n119 171.744
R339 VTAIL.n15 VTAIL.n9 171.744
R340 VTAIL.n16 VTAIL.n15 171.744
R341 VTAIL.n16 VTAIL.n5 171.744
R342 VTAIL.n23 VTAIL.n5 171.744
R343 VTAIL.n24 VTAIL.n23 171.744
R344 VTAIL.n92 VTAIL.n91 171.744
R345 VTAIL.n91 VTAIL.n73 171.744
R346 VTAIL.n84 VTAIL.n73 171.744
R347 VTAIL.n84 VTAIL.n83 171.744
R348 VTAIL.n83 VTAIL.n77 171.744
R349 VTAIL.n60 VTAIL.n59 171.744
R350 VTAIL.n59 VTAIL.n41 171.744
R351 VTAIL.n52 VTAIL.n41 171.744
R352 VTAIL.n52 VTAIL.n51 171.744
R353 VTAIL.n51 VTAIL.n45 171.744
R354 VTAIL.t7 VTAIL.n105 85.8723
R355 VTAIL.t14 VTAIL.n9 85.8723
R356 VTAIL.t11 VTAIL.n77 85.8723
R357 VTAIL.t4 VTAIL.n45 85.8723
R358 VTAIL.n69 VTAIL.n68 80.4582
R359 VTAIL.n67 VTAIL.n66 80.4582
R360 VTAIL.n37 VTAIL.n36 80.4582
R361 VTAIL.n35 VTAIL.n34 80.4582
R362 VTAIL.n127 VTAIL.n126 80.458
R363 VTAIL.n1 VTAIL.n0 80.458
R364 VTAIL.n31 VTAIL.n30 80.458
R365 VTAIL.n33 VTAIL.n32 80.458
R366 VTAIL.n125 VTAIL.n124 31.9914
R367 VTAIL.n29 VTAIL.n28 31.9914
R368 VTAIL.n97 VTAIL.n96 31.9914
R369 VTAIL.n65 VTAIL.n64 31.9914
R370 VTAIL.n35 VTAIL.n33 24.0307
R371 VTAIL.n125 VTAIL.n97 20.4703
R372 VTAIL.n107 VTAIL.n106 16.381
R373 VTAIL.n11 VTAIL.n10 16.381
R374 VTAIL.n79 VTAIL.n78 16.381
R375 VTAIL.n47 VTAIL.n46 16.381
R376 VTAIL.n110 VTAIL.n109 12.8005
R377 VTAIL.n14 VTAIL.n13 12.8005
R378 VTAIL.n82 VTAIL.n81 12.8005
R379 VTAIL.n50 VTAIL.n49 12.8005
R380 VTAIL.n113 VTAIL.n104 12.0247
R381 VTAIL.n17 VTAIL.n8 12.0247
R382 VTAIL.n85 VTAIL.n76 12.0247
R383 VTAIL.n53 VTAIL.n44 12.0247
R384 VTAIL.n114 VTAIL.n102 11.249
R385 VTAIL.n18 VTAIL.n6 11.249
R386 VTAIL.n86 VTAIL.n74 11.249
R387 VTAIL.n54 VTAIL.n42 11.249
R388 VTAIL.n118 VTAIL.n117 10.4732
R389 VTAIL.n22 VTAIL.n21 10.4732
R390 VTAIL.n90 VTAIL.n89 10.4732
R391 VTAIL.n58 VTAIL.n57 10.4732
R392 VTAIL.n121 VTAIL.n100 9.69747
R393 VTAIL.n25 VTAIL.n4 9.69747
R394 VTAIL.n93 VTAIL.n72 9.69747
R395 VTAIL.n61 VTAIL.n40 9.69747
R396 VTAIL.n124 VTAIL.n123 9.45567
R397 VTAIL.n28 VTAIL.n27 9.45567
R398 VTAIL.n96 VTAIL.n95 9.45567
R399 VTAIL.n64 VTAIL.n63 9.45567
R400 VTAIL.n123 VTAIL.n122 9.3005
R401 VTAIL.n100 VTAIL.n99 9.3005
R402 VTAIL.n117 VTAIL.n116 9.3005
R403 VTAIL.n115 VTAIL.n114 9.3005
R404 VTAIL.n104 VTAIL.n103 9.3005
R405 VTAIL.n109 VTAIL.n108 9.3005
R406 VTAIL.n27 VTAIL.n26 9.3005
R407 VTAIL.n4 VTAIL.n3 9.3005
R408 VTAIL.n21 VTAIL.n20 9.3005
R409 VTAIL.n19 VTAIL.n18 9.3005
R410 VTAIL.n8 VTAIL.n7 9.3005
R411 VTAIL.n13 VTAIL.n12 9.3005
R412 VTAIL.n95 VTAIL.n94 9.3005
R413 VTAIL.n72 VTAIL.n71 9.3005
R414 VTAIL.n89 VTAIL.n88 9.3005
R415 VTAIL.n87 VTAIL.n86 9.3005
R416 VTAIL.n76 VTAIL.n75 9.3005
R417 VTAIL.n81 VTAIL.n80 9.3005
R418 VTAIL.n63 VTAIL.n62 9.3005
R419 VTAIL.n40 VTAIL.n39 9.3005
R420 VTAIL.n57 VTAIL.n56 9.3005
R421 VTAIL.n55 VTAIL.n54 9.3005
R422 VTAIL.n44 VTAIL.n43 9.3005
R423 VTAIL.n49 VTAIL.n48 9.3005
R424 VTAIL.n122 VTAIL.n98 8.92171
R425 VTAIL.n26 VTAIL.n2 8.92171
R426 VTAIL.n94 VTAIL.n70 8.92171
R427 VTAIL.n62 VTAIL.n38 8.92171
R428 VTAIL.n126 VTAIL.t8 6.16843
R429 VTAIL.n126 VTAIL.t5 6.16843
R430 VTAIL.n0 VTAIL.t0 6.16843
R431 VTAIL.n0 VTAIL.t9 6.16843
R432 VTAIL.n30 VTAIL.t16 6.16843
R433 VTAIL.n30 VTAIL.t13 6.16843
R434 VTAIL.n32 VTAIL.t18 6.16843
R435 VTAIL.n32 VTAIL.t17 6.16843
R436 VTAIL.n68 VTAIL.t12 6.16843
R437 VTAIL.n68 VTAIL.t15 6.16843
R438 VTAIL.n66 VTAIL.t10 6.16843
R439 VTAIL.n66 VTAIL.t19 6.16843
R440 VTAIL.n36 VTAIL.t3 6.16843
R441 VTAIL.n36 VTAIL.t2 6.16843
R442 VTAIL.n34 VTAIL.t1 6.16843
R443 VTAIL.n34 VTAIL.t6 6.16843
R444 VTAIL.n124 VTAIL.n98 5.04292
R445 VTAIL.n28 VTAIL.n2 5.04292
R446 VTAIL.n96 VTAIL.n70 5.04292
R447 VTAIL.n64 VTAIL.n38 5.04292
R448 VTAIL.n122 VTAIL.n121 4.26717
R449 VTAIL.n26 VTAIL.n25 4.26717
R450 VTAIL.n94 VTAIL.n93 4.26717
R451 VTAIL.n62 VTAIL.n61 4.26717
R452 VTAIL.n80 VTAIL.n79 3.71853
R453 VTAIL.n48 VTAIL.n47 3.71853
R454 VTAIL.n108 VTAIL.n107 3.71853
R455 VTAIL.n12 VTAIL.n11 3.71853
R456 VTAIL.n37 VTAIL.n35 3.56084
R457 VTAIL.n65 VTAIL.n37 3.56084
R458 VTAIL.n69 VTAIL.n67 3.56084
R459 VTAIL.n97 VTAIL.n69 3.56084
R460 VTAIL.n33 VTAIL.n31 3.56084
R461 VTAIL.n31 VTAIL.n29 3.56084
R462 VTAIL.n127 VTAIL.n125 3.56084
R463 VTAIL.n118 VTAIL.n100 3.49141
R464 VTAIL.n22 VTAIL.n4 3.49141
R465 VTAIL.n90 VTAIL.n72 3.49141
R466 VTAIL.n58 VTAIL.n40 3.49141
R467 VTAIL VTAIL.n1 2.72895
R468 VTAIL.n117 VTAIL.n102 2.71565
R469 VTAIL.n21 VTAIL.n6 2.71565
R470 VTAIL.n89 VTAIL.n74 2.71565
R471 VTAIL.n57 VTAIL.n42 2.71565
R472 VTAIL.n67 VTAIL.n65 2.2505
R473 VTAIL.n29 VTAIL.n1 2.2505
R474 VTAIL.n114 VTAIL.n113 1.93989
R475 VTAIL.n18 VTAIL.n17 1.93989
R476 VTAIL.n86 VTAIL.n85 1.93989
R477 VTAIL.n54 VTAIL.n53 1.93989
R478 VTAIL.n110 VTAIL.n104 1.16414
R479 VTAIL.n14 VTAIL.n8 1.16414
R480 VTAIL.n82 VTAIL.n76 1.16414
R481 VTAIL.n50 VTAIL.n44 1.16414
R482 VTAIL VTAIL.n127 0.832397
R483 VTAIL.n109 VTAIL.n106 0.388379
R484 VTAIL.n13 VTAIL.n10 0.388379
R485 VTAIL.n81 VTAIL.n78 0.388379
R486 VTAIL.n49 VTAIL.n46 0.388379
R487 VTAIL.n108 VTAIL.n103 0.155672
R488 VTAIL.n115 VTAIL.n103 0.155672
R489 VTAIL.n116 VTAIL.n115 0.155672
R490 VTAIL.n116 VTAIL.n99 0.155672
R491 VTAIL.n123 VTAIL.n99 0.155672
R492 VTAIL.n12 VTAIL.n7 0.155672
R493 VTAIL.n19 VTAIL.n7 0.155672
R494 VTAIL.n20 VTAIL.n19 0.155672
R495 VTAIL.n20 VTAIL.n3 0.155672
R496 VTAIL.n27 VTAIL.n3 0.155672
R497 VTAIL.n95 VTAIL.n71 0.155672
R498 VTAIL.n88 VTAIL.n71 0.155672
R499 VTAIL.n88 VTAIL.n87 0.155672
R500 VTAIL.n87 VTAIL.n75 0.155672
R501 VTAIL.n80 VTAIL.n75 0.155672
R502 VTAIL.n63 VTAIL.n39 0.155672
R503 VTAIL.n56 VTAIL.n39 0.155672
R504 VTAIL.n56 VTAIL.n55 0.155672
R505 VTAIL.n55 VTAIL.n43 0.155672
R506 VTAIL.n48 VTAIL.n43 0.155672
R507 B.n672 B.n73 585
R508 B.n674 B.n673 585
R509 B.n675 B.n72 585
R510 B.n677 B.n676 585
R511 B.n678 B.n71 585
R512 B.n680 B.n679 585
R513 B.n681 B.n70 585
R514 B.n683 B.n682 585
R515 B.n684 B.n69 585
R516 B.n686 B.n685 585
R517 B.n687 B.n68 585
R518 B.n689 B.n688 585
R519 B.n690 B.n67 585
R520 B.n692 B.n691 585
R521 B.n693 B.n66 585
R522 B.n695 B.n694 585
R523 B.n696 B.n65 585
R524 B.n698 B.n697 585
R525 B.n699 B.n64 585
R526 B.n701 B.n700 585
R527 B.n702 B.n63 585
R528 B.n704 B.n703 585
R529 B.n706 B.n705 585
R530 B.n707 B.n59 585
R531 B.n709 B.n708 585
R532 B.n710 B.n58 585
R533 B.n712 B.n711 585
R534 B.n713 B.n57 585
R535 B.n715 B.n714 585
R536 B.n716 B.n56 585
R537 B.n718 B.n717 585
R538 B.n720 B.n53 585
R539 B.n722 B.n721 585
R540 B.n723 B.n52 585
R541 B.n725 B.n724 585
R542 B.n726 B.n51 585
R543 B.n728 B.n727 585
R544 B.n729 B.n50 585
R545 B.n731 B.n730 585
R546 B.n732 B.n49 585
R547 B.n734 B.n733 585
R548 B.n735 B.n48 585
R549 B.n737 B.n736 585
R550 B.n738 B.n47 585
R551 B.n740 B.n739 585
R552 B.n741 B.n46 585
R553 B.n743 B.n742 585
R554 B.n744 B.n45 585
R555 B.n746 B.n745 585
R556 B.n747 B.n44 585
R557 B.n749 B.n748 585
R558 B.n750 B.n43 585
R559 B.n752 B.n751 585
R560 B.n671 B.n670 585
R561 B.n669 B.n74 585
R562 B.n668 B.n667 585
R563 B.n666 B.n75 585
R564 B.n665 B.n664 585
R565 B.n663 B.n76 585
R566 B.n662 B.n661 585
R567 B.n660 B.n77 585
R568 B.n659 B.n658 585
R569 B.n657 B.n78 585
R570 B.n656 B.n655 585
R571 B.n654 B.n79 585
R572 B.n653 B.n652 585
R573 B.n651 B.n80 585
R574 B.n650 B.n649 585
R575 B.n648 B.n81 585
R576 B.n647 B.n646 585
R577 B.n645 B.n82 585
R578 B.n644 B.n643 585
R579 B.n642 B.n83 585
R580 B.n641 B.n640 585
R581 B.n639 B.n84 585
R582 B.n638 B.n637 585
R583 B.n636 B.n85 585
R584 B.n635 B.n634 585
R585 B.n633 B.n86 585
R586 B.n632 B.n631 585
R587 B.n630 B.n87 585
R588 B.n629 B.n628 585
R589 B.n627 B.n88 585
R590 B.n626 B.n625 585
R591 B.n624 B.n89 585
R592 B.n623 B.n622 585
R593 B.n621 B.n90 585
R594 B.n620 B.n619 585
R595 B.n618 B.n91 585
R596 B.n617 B.n616 585
R597 B.n615 B.n92 585
R598 B.n614 B.n613 585
R599 B.n612 B.n93 585
R600 B.n611 B.n610 585
R601 B.n609 B.n94 585
R602 B.n608 B.n607 585
R603 B.n606 B.n95 585
R604 B.n605 B.n604 585
R605 B.n603 B.n96 585
R606 B.n602 B.n601 585
R607 B.n600 B.n97 585
R608 B.n599 B.n598 585
R609 B.n597 B.n98 585
R610 B.n596 B.n595 585
R611 B.n594 B.n99 585
R612 B.n593 B.n592 585
R613 B.n591 B.n100 585
R614 B.n590 B.n589 585
R615 B.n588 B.n101 585
R616 B.n587 B.n586 585
R617 B.n585 B.n102 585
R618 B.n584 B.n583 585
R619 B.n582 B.n103 585
R620 B.n581 B.n580 585
R621 B.n579 B.n104 585
R622 B.n578 B.n577 585
R623 B.n576 B.n105 585
R624 B.n575 B.n574 585
R625 B.n573 B.n106 585
R626 B.n572 B.n571 585
R627 B.n570 B.n107 585
R628 B.n569 B.n568 585
R629 B.n567 B.n108 585
R630 B.n566 B.n565 585
R631 B.n564 B.n109 585
R632 B.n563 B.n562 585
R633 B.n561 B.n110 585
R634 B.n560 B.n559 585
R635 B.n558 B.n111 585
R636 B.n557 B.n556 585
R637 B.n555 B.n112 585
R638 B.n554 B.n553 585
R639 B.n552 B.n113 585
R640 B.n551 B.n550 585
R641 B.n549 B.n114 585
R642 B.n548 B.n547 585
R643 B.n546 B.n115 585
R644 B.n545 B.n544 585
R645 B.n543 B.n116 585
R646 B.n542 B.n541 585
R647 B.n540 B.n117 585
R648 B.n539 B.n538 585
R649 B.n537 B.n118 585
R650 B.n536 B.n535 585
R651 B.n534 B.n119 585
R652 B.n533 B.n532 585
R653 B.n531 B.n120 585
R654 B.n530 B.n529 585
R655 B.n528 B.n121 585
R656 B.n527 B.n526 585
R657 B.n525 B.n122 585
R658 B.n524 B.n523 585
R659 B.n522 B.n123 585
R660 B.n521 B.n520 585
R661 B.n519 B.n124 585
R662 B.n518 B.n517 585
R663 B.n516 B.n125 585
R664 B.n515 B.n514 585
R665 B.n513 B.n126 585
R666 B.n512 B.n511 585
R667 B.n510 B.n127 585
R668 B.n509 B.n508 585
R669 B.n507 B.n128 585
R670 B.n506 B.n505 585
R671 B.n504 B.n129 585
R672 B.n503 B.n502 585
R673 B.n501 B.n130 585
R674 B.n500 B.n499 585
R675 B.n498 B.n131 585
R676 B.n497 B.n496 585
R677 B.n495 B.n132 585
R678 B.n494 B.n493 585
R679 B.n492 B.n133 585
R680 B.n491 B.n490 585
R681 B.n489 B.n134 585
R682 B.n488 B.n487 585
R683 B.n486 B.n135 585
R684 B.n485 B.n484 585
R685 B.n483 B.n136 585
R686 B.n482 B.n481 585
R687 B.n480 B.n137 585
R688 B.n479 B.n478 585
R689 B.n477 B.n138 585
R690 B.n476 B.n475 585
R691 B.n474 B.n139 585
R692 B.n473 B.n472 585
R693 B.n471 B.n140 585
R694 B.n470 B.n469 585
R695 B.n468 B.n141 585
R696 B.n467 B.n466 585
R697 B.n465 B.n142 585
R698 B.n464 B.n463 585
R699 B.n462 B.n143 585
R700 B.n461 B.n460 585
R701 B.n459 B.n144 585
R702 B.n458 B.n457 585
R703 B.n456 B.n145 585
R704 B.n455 B.n454 585
R705 B.n453 B.n146 585
R706 B.n452 B.n451 585
R707 B.n450 B.n147 585
R708 B.n449 B.n448 585
R709 B.n447 B.n148 585
R710 B.n446 B.n445 585
R711 B.n444 B.n149 585
R712 B.n443 B.n442 585
R713 B.n441 B.n150 585
R714 B.n440 B.n439 585
R715 B.n438 B.n151 585
R716 B.n437 B.n436 585
R717 B.n435 B.n152 585
R718 B.n434 B.n433 585
R719 B.n432 B.n153 585
R720 B.n431 B.n430 585
R721 B.n429 B.n154 585
R722 B.n428 B.n427 585
R723 B.n347 B.n346 585
R724 B.n348 B.n185 585
R725 B.n350 B.n349 585
R726 B.n351 B.n184 585
R727 B.n353 B.n352 585
R728 B.n354 B.n183 585
R729 B.n356 B.n355 585
R730 B.n357 B.n182 585
R731 B.n359 B.n358 585
R732 B.n360 B.n181 585
R733 B.n362 B.n361 585
R734 B.n363 B.n180 585
R735 B.n365 B.n364 585
R736 B.n366 B.n179 585
R737 B.n368 B.n367 585
R738 B.n369 B.n178 585
R739 B.n371 B.n370 585
R740 B.n372 B.n177 585
R741 B.n374 B.n373 585
R742 B.n375 B.n176 585
R743 B.n377 B.n376 585
R744 B.n378 B.n173 585
R745 B.n381 B.n380 585
R746 B.n382 B.n172 585
R747 B.n384 B.n383 585
R748 B.n385 B.n171 585
R749 B.n387 B.n386 585
R750 B.n388 B.n170 585
R751 B.n390 B.n389 585
R752 B.n391 B.n169 585
R753 B.n393 B.n392 585
R754 B.n395 B.n394 585
R755 B.n396 B.n165 585
R756 B.n398 B.n397 585
R757 B.n399 B.n164 585
R758 B.n401 B.n400 585
R759 B.n402 B.n163 585
R760 B.n404 B.n403 585
R761 B.n405 B.n162 585
R762 B.n407 B.n406 585
R763 B.n408 B.n161 585
R764 B.n410 B.n409 585
R765 B.n411 B.n160 585
R766 B.n413 B.n412 585
R767 B.n414 B.n159 585
R768 B.n416 B.n415 585
R769 B.n417 B.n158 585
R770 B.n419 B.n418 585
R771 B.n420 B.n157 585
R772 B.n422 B.n421 585
R773 B.n423 B.n156 585
R774 B.n425 B.n424 585
R775 B.n426 B.n155 585
R776 B.n345 B.n186 585
R777 B.n344 B.n343 585
R778 B.n342 B.n187 585
R779 B.n341 B.n340 585
R780 B.n339 B.n188 585
R781 B.n338 B.n337 585
R782 B.n336 B.n189 585
R783 B.n335 B.n334 585
R784 B.n333 B.n190 585
R785 B.n332 B.n331 585
R786 B.n330 B.n191 585
R787 B.n329 B.n328 585
R788 B.n327 B.n192 585
R789 B.n326 B.n325 585
R790 B.n324 B.n193 585
R791 B.n323 B.n322 585
R792 B.n321 B.n194 585
R793 B.n320 B.n319 585
R794 B.n318 B.n195 585
R795 B.n317 B.n316 585
R796 B.n315 B.n196 585
R797 B.n314 B.n313 585
R798 B.n312 B.n197 585
R799 B.n311 B.n310 585
R800 B.n309 B.n198 585
R801 B.n308 B.n307 585
R802 B.n306 B.n199 585
R803 B.n305 B.n304 585
R804 B.n303 B.n200 585
R805 B.n302 B.n301 585
R806 B.n300 B.n201 585
R807 B.n299 B.n298 585
R808 B.n297 B.n202 585
R809 B.n296 B.n295 585
R810 B.n294 B.n203 585
R811 B.n293 B.n292 585
R812 B.n291 B.n204 585
R813 B.n290 B.n289 585
R814 B.n288 B.n205 585
R815 B.n287 B.n286 585
R816 B.n285 B.n206 585
R817 B.n284 B.n283 585
R818 B.n282 B.n207 585
R819 B.n281 B.n280 585
R820 B.n279 B.n208 585
R821 B.n278 B.n277 585
R822 B.n276 B.n209 585
R823 B.n275 B.n274 585
R824 B.n273 B.n210 585
R825 B.n272 B.n271 585
R826 B.n270 B.n211 585
R827 B.n269 B.n268 585
R828 B.n267 B.n212 585
R829 B.n266 B.n265 585
R830 B.n264 B.n213 585
R831 B.n263 B.n262 585
R832 B.n261 B.n214 585
R833 B.n260 B.n259 585
R834 B.n258 B.n215 585
R835 B.n257 B.n256 585
R836 B.n255 B.n216 585
R837 B.n254 B.n253 585
R838 B.n252 B.n217 585
R839 B.n251 B.n250 585
R840 B.n249 B.n218 585
R841 B.n248 B.n247 585
R842 B.n246 B.n219 585
R843 B.n245 B.n244 585
R844 B.n243 B.n220 585
R845 B.n242 B.n241 585
R846 B.n240 B.n221 585
R847 B.n239 B.n238 585
R848 B.n237 B.n222 585
R849 B.n236 B.n235 585
R850 B.n234 B.n223 585
R851 B.n233 B.n232 585
R852 B.n231 B.n224 585
R853 B.n230 B.n229 585
R854 B.n228 B.n225 585
R855 B.n227 B.n226 585
R856 B.n2 B.n0 585
R857 B.n873 B.n1 585
R858 B.n872 B.n871 585
R859 B.n870 B.n3 585
R860 B.n869 B.n868 585
R861 B.n867 B.n4 585
R862 B.n866 B.n865 585
R863 B.n864 B.n5 585
R864 B.n863 B.n862 585
R865 B.n861 B.n6 585
R866 B.n860 B.n859 585
R867 B.n858 B.n7 585
R868 B.n857 B.n856 585
R869 B.n855 B.n8 585
R870 B.n854 B.n853 585
R871 B.n852 B.n9 585
R872 B.n851 B.n850 585
R873 B.n849 B.n10 585
R874 B.n848 B.n847 585
R875 B.n846 B.n11 585
R876 B.n845 B.n844 585
R877 B.n843 B.n12 585
R878 B.n842 B.n841 585
R879 B.n840 B.n13 585
R880 B.n839 B.n838 585
R881 B.n837 B.n14 585
R882 B.n836 B.n835 585
R883 B.n834 B.n15 585
R884 B.n833 B.n832 585
R885 B.n831 B.n16 585
R886 B.n830 B.n829 585
R887 B.n828 B.n17 585
R888 B.n827 B.n826 585
R889 B.n825 B.n18 585
R890 B.n824 B.n823 585
R891 B.n822 B.n19 585
R892 B.n821 B.n820 585
R893 B.n819 B.n20 585
R894 B.n818 B.n817 585
R895 B.n816 B.n21 585
R896 B.n815 B.n814 585
R897 B.n813 B.n22 585
R898 B.n812 B.n811 585
R899 B.n810 B.n23 585
R900 B.n809 B.n808 585
R901 B.n807 B.n24 585
R902 B.n806 B.n805 585
R903 B.n804 B.n25 585
R904 B.n803 B.n802 585
R905 B.n801 B.n26 585
R906 B.n800 B.n799 585
R907 B.n798 B.n27 585
R908 B.n797 B.n796 585
R909 B.n795 B.n28 585
R910 B.n794 B.n793 585
R911 B.n792 B.n29 585
R912 B.n791 B.n790 585
R913 B.n789 B.n30 585
R914 B.n788 B.n787 585
R915 B.n786 B.n31 585
R916 B.n785 B.n784 585
R917 B.n783 B.n32 585
R918 B.n782 B.n781 585
R919 B.n780 B.n33 585
R920 B.n779 B.n778 585
R921 B.n777 B.n34 585
R922 B.n776 B.n775 585
R923 B.n774 B.n35 585
R924 B.n773 B.n772 585
R925 B.n771 B.n36 585
R926 B.n770 B.n769 585
R927 B.n768 B.n37 585
R928 B.n767 B.n766 585
R929 B.n765 B.n38 585
R930 B.n764 B.n763 585
R931 B.n762 B.n39 585
R932 B.n761 B.n760 585
R933 B.n759 B.n40 585
R934 B.n758 B.n757 585
R935 B.n756 B.n41 585
R936 B.n755 B.n754 585
R937 B.n753 B.n42 585
R938 B.n875 B.n874 585
R939 B.n346 B.n345 516.524
R940 B.n753 B.n752 516.524
R941 B.n428 B.n155 516.524
R942 B.n670 B.n73 516.524
R943 B.n166 B.t2 335.551
R944 B.n60 B.t4 335.551
R945 B.n174 B.t11 335.551
R946 B.n54 B.t7 335.551
R947 B.n167 B.t1 255.454
R948 B.n61 B.t5 255.454
R949 B.n175 B.t10 255.454
R950 B.n55 B.t8 255.454
R951 B.n166 B.t0 242.767
R952 B.n174 B.t9 242.767
R953 B.n54 B.t6 242.767
R954 B.n60 B.t3 242.767
R955 B.n345 B.n344 163.367
R956 B.n344 B.n187 163.367
R957 B.n340 B.n187 163.367
R958 B.n340 B.n339 163.367
R959 B.n339 B.n338 163.367
R960 B.n338 B.n189 163.367
R961 B.n334 B.n189 163.367
R962 B.n334 B.n333 163.367
R963 B.n333 B.n332 163.367
R964 B.n332 B.n191 163.367
R965 B.n328 B.n191 163.367
R966 B.n328 B.n327 163.367
R967 B.n327 B.n326 163.367
R968 B.n326 B.n193 163.367
R969 B.n322 B.n193 163.367
R970 B.n322 B.n321 163.367
R971 B.n321 B.n320 163.367
R972 B.n320 B.n195 163.367
R973 B.n316 B.n195 163.367
R974 B.n316 B.n315 163.367
R975 B.n315 B.n314 163.367
R976 B.n314 B.n197 163.367
R977 B.n310 B.n197 163.367
R978 B.n310 B.n309 163.367
R979 B.n309 B.n308 163.367
R980 B.n308 B.n199 163.367
R981 B.n304 B.n199 163.367
R982 B.n304 B.n303 163.367
R983 B.n303 B.n302 163.367
R984 B.n302 B.n201 163.367
R985 B.n298 B.n201 163.367
R986 B.n298 B.n297 163.367
R987 B.n297 B.n296 163.367
R988 B.n296 B.n203 163.367
R989 B.n292 B.n203 163.367
R990 B.n292 B.n291 163.367
R991 B.n291 B.n290 163.367
R992 B.n290 B.n205 163.367
R993 B.n286 B.n205 163.367
R994 B.n286 B.n285 163.367
R995 B.n285 B.n284 163.367
R996 B.n284 B.n207 163.367
R997 B.n280 B.n207 163.367
R998 B.n280 B.n279 163.367
R999 B.n279 B.n278 163.367
R1000 B.n278 B.n209 163.367
R1001 B.n274 B.n209 163.367
R1002 B.n274 B.n273 163.367
R1003 B.n273 B.n272 163.367
R1004 B.n272 B.n211 163.367
R1005 B.n268 B.n211 163.367
R1006 B.n268 B.n267 163.367
R1007 B.n267 B.n266 163.367
R1008 B.n266 B.n213 163.367
R1009 B.n262 B.n213 163.367
R1010 B.n262 B.n261 163.367
R1011 B.n261 B.n260 163.367
R1012 B.n260 B.n215 163.367
R1013 B.n256 B.n215 163.367
R1014 B.n256 B.n255 163.367
R1015 B.n255 B.n254 163.367
R1016 B.n254 B.n217 163.367
R1017 B.n250 B.n217 163.367
R1018 B.n250 B.n249 163.367
R1019 B.n249 B.n248 163.367
R1020 B.n248 B.n219 163.367
R1021 B.n244 B.n219 163.367
R1022 B.n244 B.n243 163.367
R1023 B.n243 B.n242 163.367
R1024 B.n242 B.n221 163.367
R1025 B.n238 B.n221 163.367
R1026 B.n238 B.n237 163.367
R1027 B.n237 B.n236 163.367
R1028 B.n236 B.n223 163.367
R1029 B.n232 B.n223 163.367
R1030 B.n232 B.n231 163.367
R1031 B.n231 B.n230 163.367
R1032 B.n230 B.n225 163.367
R1033 B.n226 B.n225 163.367
R1034 B.n226 B.n2 163.367
R1035 B.n874 B.n2 163.367
R1036 B.n874 B.n873 163.367
R1037 B.n873 B.n872 163.367
R1038 B.n872 B.n3 163.367
R1039 B.n868 B.n3 163.367
R1040 B.n868 B.n867 163.367
R1041 B.n867 B.n866 163.367
R1042 B.n866 B.n5 163.367
R1043 B.n862 B.n5 163.367
R1044 B.n862 B.n861 163.367
R1045 B.n861 B.n860 163.367
R1046 B.n860 B.n7 163.367
R1047 B.n856 B.n7 163.367
R1048 B.n856 B.n855 163.367
R1049 B.n855 B.n854 163.367
R1050 B.n854 B.n9 163.367
R1051 B.n850 B.n9 163.367
R1052 B.n850 B.n849 163.367
R1053 B.n849 B.n848 163.367
R1054 B.n848 B.n11 163.367
R1055 B.n844 B.n11 163.367
R1056 B.n844 B.n843 163.367
R1057 B.n843 B.n842 163.367
R1058 B.n842 B.n13 163.367
R1059 B.n838 B.n13 163.367
R1060 B.n838 B.n837 163.367
R1061 B.n837 B.n836 163.367
R1062 B.n836 B.n15 163.367
R1063 B.n832 B.n15 163.367
R1064 B.n832 B.n831 163.367
R1065 B.n831 B.n830 163.367
R1066 B.n830 B.n17 163.367
R1067 B.n826 B.n17 163.367
R1068 B.n826 B.n825 163.367
R1069 B.n825 B.n824 163.367
R1070 B.n824 B.n19 163.367
R1071 B.n820 B.n19 163.367
R1072 B.n820 B.n819 163.367
R1073 B.n819 B.n818 163.367
R1074 B.n818 B.n21 163.367
R1075 B.n814 B.n21 163.367
R1076 B.n814 B.n813 163.367
R1077 B.n813 B.n812 163.367
R1078 B.n812 B.n23 163.367
R1079 B.n808 B.n23 163.367
R1080 B.n808 B.n807 163.367
R1081 B.n807 B.n806 163.367
R1082 B.n806 B.n25 163.367
R1083 B.n802 B.n25 163.367
R1084 B.n802 B.n801 163.367
R1085 B.n801 B.n800 163.367
R1086 B.n800 B.n27 163.367
R1087 B.n796 B.n27 163.367
R1088 B.n796 B.n795 163.367
R1089 B.n795 B.n794 163.367
R1090 B.n794 B.n29 163.367
R1091 B.n790 B.n29 163.367
R1092 B.n790 B.n789 163.367
R1093 B.n789 B.n788 163.367
R1094 B.n788 B.n31 163.367
R1095 B.n784 B.n31 163.367
R1096 B.n784 B.n783 163.367
R1097 B.n783 B.n782 163.367
R1098 B.n782 B.n33 163.367
R1099 B.n778 B.n33 163.367
R1100 B.n778 B.n777 163.367
R1101 B.n777 B.n776 163.367
R1102 B.n776 B.n35 163.367
R1103 B.n772 B.n35 163.367
R1104 B.n772 B.n771 163.367
R1105 B.n771 B.n770 163.367
R1106 B.n770 B.n37 163.367
R1107 B.n766 B.n37 163.367
R1108 B.n766 B.n765 163.367
R1109 B.n765 B.n764 163.367
R1110 B.n764 B.n39 163.367
R1111 B.n760 B.n39 163.367
R1112 B.n760 B.n759 163.367
R1113 B.n759 B.n758 163.367
R1114 B.n758 B.n41 163.367
R1115 B.n754 B.n41 163.367
R1116 B.n754 B.n753 163.367
R1117 B.n346 B.n185 163.367
R1118 B.n350 B.n185 163.367
R1119 B.n351 B.n350 163.367
R1120 B.n352 B.n351 163.367
R1121 B.n352 B.n183 163.367
R1122 B.n356 B.n183 163.367
R1123 B.n357 B.n356 163.367
R1124 B.n358 B.n357 163.367
R1125 B.n358 B.n181 163.367
R1126 B.n362 B.n181 163.367
R1127 B.n363 B.n362 163.367
R1128 B.n364 B.n363 163.367
R1129 B.n364 B.n179 163.367
R1130 B.n368 B.n179 163.367
R1131 B.n369 B.n368 163.367
R1132 B.n370 B.n369 163.367
R1133 B.n370 B.n177 163.367
R1134 B.n374 B.n177 163.367
R1135 B.n375 B.n374 163.367
R1136 B.n376 B.n375 163.367
R1137 B.n376 B.n173 163.367
R1138 B.n381 B.n173 163.367
R1139 B.n382 B.n381 163.367
R1140 B.n383 B.n382 163.367
R1141 B.n383 B.n171 163.367
R1142 B.n387 B.n171 163.367
R1143 B.n388 B.n387 163.367
R1144 B.n389 B.n388 163.367
R1145 B.n389 B.n169 163.367
R1146 B.n393 B.n169 163.367
R1147 B.n394 B.n393 163.367
R1148 B.n394 B.n165 163.367
R1149 B.n398 B.n165 163.367
R1150 B.n399 B.n398 163.367
R1151 B.n400 B.n399 163.367
R1152 B.n400 B.n163 163.367
R1153 B.n404 B.n163 163.367
R1154 B.n405 B.n404 163.367
R1155 B.n406 B.n405 163.367
R1156 B.n406 B.n161 163.367
R1157 B.n410 B.n161 163.367
R1158 B.n411 B.n410 163.367
R1159 B.n412 B.n411 163.367
R1160 B.n412 B.n159 163.367
R1161 B.n416 B.n159 163.367
R1162 B.n417 B.n416 163.367
R1163 B.n418 B.n417 163.367
R1164 B.n418 B.n157 163.367
R1165 B.n422 B.n157 163.367
R1166 B.n423 B.n422 163.367
R1167 B.n424 B.n423 163.367
R1168 B.n424 B.n155 163.367
R1169 B.n429 B.n428 163.367
R1170 B.n430 B.n429 163.367
R1171 B.n430 B.n153 163.367
R1172 B.n434 B.n153 163.367
R1173 B.n435 B.n434 163.367
R1174 B.n436 B.n435 163.367
R1175 B.n436 B.n151 163.367
R1176 B.n440 B.n151 163.367
R1177 B.n441 B.n440 163.367
R1178 B.n442 B.n441 163.367
R1179 B.n442 B.n149 163.367
R1180 B.n446 B.n149 163.367
R1181 B.n447 B.n446 163.367
R1182 B.n448 B.n447 163.367
R1183 B.n448 B.n147 163.367
R1184 B.n452 B.n147 163.367
R1185 B.n453 B.n452 163.367
R1186 B.n454 B.n453 163.367
R1187 B.n454 B.n145 163.367
R1188 B.n458 B.n145 163.367
R1189 B.n459 B.n458 163.367
R1190 B.n460 B.n459 163.367
R1191 B.n460 B.n143 163.367
R1192 B.n464 B.n143 163.367
R1193 B.n465 B.n464 163.367
R1194 B.n466 B.n465 163.367
R1195 B.n466 B.n141 163.367
R1196 B.n470 B.n141 163.367
R1197 B.n471 B.n470 163.367
R1198 B.n472 B.n471 163.367
R1199 B.n472 B.n139 163.367
R1200 B.n476 B.n139 163.367
R1201 B.n477 B.n476 163.367
R1202 B.n478 B.n477 163.367
R1203 B.n478 B.n137 163.367
R1204 B.n482 B.n137 163.367
R1205 B.n483 B.n482 163.367
R1206 B.n484 B.n483 163.367
R1207 B.n484 B.n135 163.367
R1208 B.n488 B.n135 163.367
R1209 B.n489 B.n488 163.367
R1210 B.n490 B.n489 163.367
R1211 B.n490 B.n133 163.367
R1212 B.n494 B.n133 163.367
R1213 B.n495 B.n494 163.367
R1214 B.n496 B.n495 163.367
R1215 B.n496 B.n131 163.367
R1216 B.n500 B.n131 163.367
R1217 B.n501 B.n500 163.367
R1218 B.n502 B.n501 163.367
R1219 B.n502 B.n129 163.367
R1220 B.n506 B.n129 163.367
R1221 B.n507 B.n506 163.367
R1222 B.n508 B.n507 163.367
R1223 B.n508 B.n127 163.367
R1224 B.n512 B.n127 163.367
R1225 B.n513 B.n512 163.367
R1226 B.n514 B.n513 163.367
R1227 B.n514 B.n125 163.367
R1228 B.n518 B.n125 163.367
R1229 B.n519 B.n518 163.367
R1230 B.n520 B.n519 163.367
R1231 B.n520 B.n123 163.367
R1232 B.n524 B.n123 163.367
R1233 B.n525 B.n524 163.367
R1234 B.n526 B.n525 163.367
R1235 B.n526 B.n121 163.367
R1236 B.n530 B.n121 163.367
R1237 B.n531 B.n530 163.367
R1238 B.n532 B.n531 163.367
R1239 B.n532 B.n119 163.367
R1240 B.n536 B.n119 163.367
R1241 B.n537 B.n536 163.367
R1242 B.n538 B.n537 163.367
R1243 B.n538 B.n117 163.367
R1244 B.n542 B.n117 163.367
R1245 B.n543 B.n542 163.367
R1246 B.n544 B.n543 163.367
R1247 B.n544 B.n115 163.367
R1248 B.n548 B.n115 163.367
R1249 B.n549 B.n548 163.367
R1250 B.n550 B.n549 163.367
R1251 B.n550 B.n113 163.367
R1252 B.n554 B.n113 163.367
R1253 B.n555 B.n554 163.367
R1254 B.n556 B.n555 163.367
R1255 B.n556 B.n111 163.367
R1256 B.n560 B.n111 163.367
R1257 B.n561 B.n560 163.367
R1258 B.n562 B.n561 163.367
R1259 B.n562 B.n109 163.367
R1260 B.n566 B.n109 163.367
R1261 B.n567 B.n566 163.367
R1262 B.n568 B.n567 163.367
R1263 B.n568 B.n107 163.367
R1264 B.n572 B.n107 163.367
R1265 B.n573 B.n572 163.367
R1266 B.n574 B.n573 163.367
R1267 B.n574 B.n105 163.367
R1268 B.n578 B.n105 163.367
R1269 B.n579 B.n578 163.367
R1270 B.n580 B.n579 163.367
R1271 B.n580 B.n103 163.367
R1272 B.n584 B.n103 163.367
R1273 B.n585 B.n584 163.367
R1274 B.n586 B.n585 163.367
R1275 B.n586 B.n101 163.367
R1276 B.n590 B.n101 163.367
R1277 B.n591 B.n590 163.367
R1278 B.n592 B.n591 163.367
R1279 B.n592 B.n99 163.367
R1280 B.n596 B.n99 163.367
R1281 B.n597 B.n596 163.367
R1282 B.n598 B.n597 163.367
R1283 B.n598 B.n97 163.367
R1284 B.n602 B.n97 163.367
R1285 B.n603 B.n602 163.367
R1286 B.n604 B.n603 163.367
R1287 B.n604 B.n95 163.367
R1288 B.n608 B.n95 163.367
R1289 B.n609 B.n608 163.367
R1290 B.n610 B.n609 163.367
R1291 B.n610 B.n93 163.367
R1292 B.n614 B.n93 163.367
R1293 B.n615 B.n614 163.367
R1294 B.n616 B.n615 163.367
R1295 B.n616 B.n91 163.367
R1296 B.n620 B.n91 163.367
R1297 B.n621 B.n620 163.367
R1298 B.n622 B.n621 163.367
R1299 B.n622 B.n89 163.367
R1300 B.n626 B.n89 163.367
R1301 B.n627 B.n626 163.367
R1302 B.n628 B.n627 163.367
R1303 B.n628 B.n87 163.367
R1304 B.n632 B.n87 163.367
R1305 B.n633 B.n632 163.367
R1306 B.n634 B.n633 163.367
R1307 B.n634 B.n85 163.367
R1308 B.n638 B.n85 163.367
R1309 B.n639 B.n638 163.367
R1310 B.n640 B.n639 163.367
R1311 B.n640 B.n83 163.367
R1312 B.n644 B.n83 163.367
R1313 B.n645 B.n644 163.367
R1314 B.n646 B.n645 163.367
R1315 B.n646 B.n81 163.367
R1316 B.n650 B.n81 163.367
R1317 B.n651 B.n650 163.367
R1318 B.n652 B.n651 163.367
R1319 B.n652 B.n79 163.367
R1320 B.n656 B.n79 163.367
R1321 B.n657 B.n656 163.367
R1322 B.n658 B.n657 163.367
R1323 B.n658 B.n77 163.367
R1324 B.n662 B.n77 163.367
R1325 B.n663 B.n662 163.367
R1326 B.n664 B.n663 163.367
R1327 B.n664 B.n75 163.367
R1328 B.n668 B.n75 163.367
R1329 B.n669 B.n668 163.367
R1330 B.n670 B.n669 163.367
R1331 B.n752 B.n43 163.367
R1332 B.n748 B.n43 163.367
R1333 B.n748 B.n747 163.367
R1334 B.n747 B.n746 163.367
R1335 B.n746 B.n45 163.367
R1336 B.n742 B.n45 163.367
R1337 B.n742 B.n741 163.367
R1338 B.n741 B.n740 163.367
R1339 B.n740 B.n47 163.367
R1340 B.n736 B.n47 163.367
R1341 B.n736 B.n735 163.367
R1342 B.n735 B.n734 163.367
R1343 B.n734 B.n49 163.367
R1344 B.n730 B.n49 163.367
R1345 B.n730 B.n729 163.367
R1346 B.n729 B.n728 163.367
R1347 B.n728 B.n51 163.367
R1348 B.n724 B.n51 163.367
R1349 B.n724 B.n723 163.367
R1350 B.n723 B.n722 163.367
R1351 B.n722 B.n53 163.367
R1352 B.n717 B.n53 163.367
R1353 B.n717 B.n716 163.367
R1354 B.n716 B.n715 163.367
R1355 B.n715 B.n57 163.367
R1356 B.n711 B.n57 163.367
R1357 B.n711 B.n710 163.367
R1358 B.n710 B.n709 163.367
R1359 B.n709 B.n59 163.367
R1360 B.n705 B.n59 163.367
R1361 B.n705 B.n704 163.367
R1362 B.n704 B.n63 163.367
R1363 B.n700 B.n63 163.367
R1364 B.n700 B.n699 163.367
R1365 B.n699 B.n698 163.367
R1366 B.n698 B.n65 163.367
R1367 B.n694 B.n65 163.367
R1368 B.n694 B.n693 163.367
R1369 B.n693 B.n692 163.367
R1370 B.n692 B.n67 163.367
R1371 B.n688 B.n67 163.367
R1372 B.n688 B.n687 163.367
R1373 B.n687 B.n686 163.367
R1374 B.n686 B.n69 163.367
R1375 B.n682 B.n69 163.367
R1376 B.n682 B.n681 163.367
R1377 B.n681 B.n680 163.367
R1378 B.n680 B.n71 163.367
R1379 B.n676 B.n71 163.367
R1380 B.n676 B.n675 163.367
R1381 B.n675 B.n674 163.367
R1382 B.n674 B.n73 163.367
R1383 B.n167 B.n166 80.0975
R1384 B.n175 B.n174 80.0975
R1385 B.n55 B.n54 80.0975
R1386 B.n61 B.n60 80.0975
R1387 B.n168 B.n167 59.5399
R1388 B.n379 B.n175 59.5399
R1389 B.n719 B.n55 59.5399
R1390 B.n62 B.n61 59.5399
R1391 B.n751 B.n42 33.5615
R1392 B.n672 B.n671 33.5615
R1393 B.n427 B.n426 33.5615
R1394 B.n347 B.n186 33.5615
R1395 B B.n875 18.0485
R1396 B.n751 B.n750 10.6151
R1397 B.n750 B.n749 10.6151
R1398 B.n749 B.n44 10.6151
R1399 B.n745 B.n44 10.6151
R1400 B.n745 B.n744 10.6151
R1401 B.n744 B.n743 10.6151
R1402 B.n743 B.n46 10.6151
R1403 B.n739 B.n46 10.6151
R1404 B.n739 B.n738 10.6151
R1405 B.n738 B.n737 10.6151
R1406 B.n737 B.n48 10.6151
R1407 B.n733 B.n48 10.6151
R1408 B.n733 B.n732 10.6151
R1409 B.n732 B.n731 10.6151
R1410 B.n731 B.n50 10.6151
R1411 B.n727 B.n50 10.6151
R1412 B.n727 B.n726 10.6151
R1413 B.n726 B.n725 10.6151
R1414 B.n725 B.n52 10.6151
R1415 B.n721 B.n52 10.6151
R1416 B.n721 B.n720 10.6151
R1417 B.n718 B.n56 10.6151
R1418 B.n714 B.n56 10.6151
R1419 B.n714 B.n713 10.6151
R1420 B.n713 B.n712 10.6151
R1421 B.n712 B.n58 10.6151
R1422 B.n708 B.n58 10.6151
R1423 B.n708 B.n707 10.6151
R1424 B.n707 B.n706 10.6151
R1425 B.n703 B.n702 10.6151
R1426 B.n702 B.n701 10.6151
R1427 B.n701 B.n64 10.6151
R1428 B.n697 B.n64 10.6151
R1429 B.n697 B.n696 10.6151
R1430 B.n696 B.n695 10.6151
R1431 B.n695 B.n66 10.6151
R1432 B.n691 B.n66 10.6151
R1433 B.n691 B.n690 10.6151
R1434 B.n690 B.n689 10.6151
R1435 B.n689 B.n68 10.6151
R1436 B.n685 B.n68 10.6151
R1437 B.n685 B.n684 10.6151
R1438 B.n684 B.n683 10.6151
R1439 B.n683 B.n70 10.6151
R1440 B.n679 B.n70 10.6151
R1441 B.n679 B.n678 10.6151
R1442 B.n678 B.n677 10.6151
R1443 B.n677 B.n72 10.6151
R1444 B.n673 B.n72 10.6151
R1445 B.n673 B.n672 10.6151
R1446 B.n427 B.n154 10.6151
R1447 B.n431 B.n154 10.6151
R1448 B.n432 B.n431 10.6151
R1449 B.n433 B.n432 10.6151
R1450 B.n433 B.n152 10.6151
R1451 B.n437 B.n152 10.6151
R1452 B.n438 B.n437 10.6151
R1453 B.n439 B.n438 10.6151
R1454 B.n439 B.n150 10.6151
R1455 B.n443 B.n150 10.6151
R1456 B.n444 B.n443 10.6151
R1457 B.n445 B.n444 10.6151
R1458 B.n445 B.n148 10.6151
R1459 B.n449 B.n148 10.6151
R1460 B.n450 B.n449 10.6151
R1461 B.n451 B.n450 10.6151
R1462 B.n451 B.n146 10.6151
R1463 B.n455 B.n146 10.6151
R1464 B.n456 B.n455 10.6151
R1465 B.n457 B.n456 10.6151
R1466 B.n457 B.n144 10.6151
R1467 B.n461 B.n144 10.6151
R1468 B.n462 B.n461 10.6151
R1469 B.n463 B.n462 10.6151
R1470 B.n463 B.n142 10.6151
R1471 B.n467 B.n142 10.6151
R1472 B.n468 B.n467 10.6151
R1473 B.n469 B.n468 10.6151
R1474 B.n469 B.n140 10.6151
R1475 B.n473 B.n140 10.6151
R1476 B.n474 B.n473 10.6151
R1477 B.n475 B.n474 10.6151
R1478 B.n475 B.n138 10.6151
R1479 B.n479 B.n138 10.6151
R1480 B.n480 B.n479 10.6151
R1481 B.n481 B.n480 10.6151
R1482 B.n481 B.n136 10.6151
R1483 B.n485 B.n136 10.6151
R1484 B.n486 B.n485 10.6151
R1485 B.n487 B.n486 10.6151
R1486 B.n487 B.n134 10.6151
R1487 B.n491 B.n134 10.6151
R1488 B.n492 B.n491 10.6151
R1489 B.n493 B.n492 10.6151
R1490 B.n493 B.n132 10.6151
R1491 B.n497 B.n132 10.6151
R1492 B.n498 B.n497 10.6151
R1493 B.n499 B.n498 10.6151
R1494 B.n499 B.n130 10.6151
R1495 B.n503 B.n130 10.6151
R1496 B.n504 B.n503 10.6151
R1497 B.n505 B.n504 10.6151
R1498 B.n505 B.n128 10.6151
R1499 B.n509 B.n128 10.6151
R1500 B.n510 B.n509 10.6151
R1501 B.n511 B.n510 10.6151
R1502 B.n511 B.n126 10.6151
R1503 B.n515 B.n126 10.6151
R1504 B.n516 B.n515 10.6151
R1505 B.n517 B.n516 10.6151
R1506 B.n517 B.n124 10.6151
R1507 B.n521 B.n124 10.6151
R1508 B.n522 B.n521 10.6151
R1509 B.n523 B.n522 10.6151
R1510 B.n523 B.n122 10.6151
R1511 B.n527 B.n122 10.6151
R1512 B.n528 B.n527 10.6151
R1513 B.n529 B.n528 10.6151
R1514 B.n529 B.n120 10.6151
R1515 B.n533 B.n120 10.6151
R1516 B.n534 B.n533 10.6151
R1517 B.n535 B.n534 10.6151
R1518 B.n535 B.n118 10.6151
R1519 B.n539 B.n118 10.6151
R1520 B.n540 B.n539 10.6151
R1521 B.n541 B.n540 10.6151
R1522 B.n541 B.n116 10.6151
R1523 B.n545 B.n116 10.6151
R1524 B.n546 B.n545 10.6151
R1525 B.n547 B.n546 10.6151
R1526 B.n547 B.n114 10.6151
R1527 B.n551 B.n114 10.6151
R1528 B.n552 B.n551 10.6151
R1529 B.n553 B.n552 10.6151
R1530 B.n553 B.n112 10.6151
R1531 B.n557 B.n112 10.6151
R1532 B.n558 B.n557 10.6151
R1533 B.n559 B.n558 10.6151
R1534 B.n559 B.n110 10.6151
R1535 B.n563 B.n110 10.6151
R1536 B.n564 B.n563 10.6151
R1537 B.n565 B.n564 10.6151
R1538 B.n565 B.n108 10.6151
R1539 B.n569 B.n108 10.6151
R1540 B.n570 B.n569 10.6151
R1541 B.n571 B.n570 10.6151
R1542 B.n571 B.n106 10.6151
R1543 B.n575 B.n106 10.6151
R1544 B.n576 B.n575 10.6151
R1545 B.n577 B.n576 10.6151
R1546 B.n577 B.n104 10.6151
R1547 B.n581 B.n104 10.6151
R1548 B.n582 B.n581 10.6151
R1549 B.n583 B.n582 10.6151
R1550 B.n583 B.n102 10.6151
R1551 B.n587 B.n102 10.6151
R1552 B.n588 B.n587 10.6151
R1553 B.n589 B.n588 10.6151
R1554 B.n589 B.n100 10.6151
R1555 B.n593 B.n100 10.6151
R1556 B.n594 B.n593 10.6151
R1557 B.n595 B.n594 10.6151
R1558 B.n595 B.n98 10.6151
R1559 B.n599 B.n98 10.6151
R1560 B.n600 B.n599 10.6151
R1561 B.n601 B.n600 10.6151
R1562 B.n601 B.n96 10.6151
R1563 B.n605 B.n96 10.6151
R1564 B.n606 B.n605 10.6151
R1565 B.n607 B.n606 10.6151
R1566 B.n607 B.n94 10.6151
R1567 B.n611 B.n94 10.6151
R1568 B.n612 B.n611 10.6151
R1569 B.n613 B.n612 10.6151
R1570 B.n613 B.n92 10.6151
R1571 B.n617 B.n92 10.6151
R1572 B.n618 B.n617 10.6151
R1573 B.n619 B.n618 10.6151
R1574 B.n619 B.n90 10.6151
R1575 B.n623 B.n90 10.6151
R1576 B.n624 B.n623 10.6151
R1577 B.n625 B.n624 10.6151
R1578 B.n625 B.n88 10.6151
R1579 B.n629 B.n88 10.6151
R1580 B.n630 B.n629 10.6151
R1581 B.n631 B.n630 10.6151
R1582 B.n631 B.n86 10.6151
R1583 B.n635 B.n86 10.6151
R1584 B.n636 B.n635 10.6151
R1585 B.n637 B.n636 10.6151
R1586 B.n637 B.n84 10.6151
R1587 B.n641 B.n84 10.6151
R1588 B.n642 B.n641 10.6151
R1589 B.n643 B.n642 10.6151
R1590 B.n643 B.n82 10.6151
R1591 B.n647 B.n82 10.6151
R1592 B.n648 B.n647 10.6151
R1593 B.n649 B.n648 10.6151
R1594 B.n649 B.n80 10.6151
R1595 B.n653 B.n80 10.6151
R1596 B.n654 B.n653 10.6151
R1597 B.n655 B.n654 10.6151
R1598 B.n655 B.n78 10.6151
R1599 B.n659 B.n78 10.6151
R1600 B.n660 B.n659 10.6151
R1601 B.n661 B.n660 10.6151
R1602 B.n661 B.n76 10.6151
R1603 B.n665 B.n76 10.6151
R1604 B.n666 B.n665 10.6151
R1605 B.n667 B.n666 10.6151
R1606 B.n667 B.n74 10.6151
R1607 B.n671 B.n74 10.6151
R1608 B.n348 B.n347 10.6151
R1609 B.n349 B.n348 10.6151
R1610 B.n349 B.n184 10.6151
R1611 B.n353 B.n184 10.6151
R1612 B.n354 B.n353 10.6151
R1613 B.n355 B.n354 10.6151
R1614 B.n355 B.n182 10.6151
R1615 B.n359 B.n182 10.6151
R1616 B.n360 B.n359 10.6151
R1617 B.n361 B.n360 10.6151
R1618 B.n361 B.n180 10.6151
R1619 B.n365 B.n180 10.6151
R1620 B.n366 B.n365 10.6151
R1621 B.n367 B.n366 10.6151
R1622 B.n367 B.n178 10.6151
R1623 B.n371 B.n178 10.6151
R1624 B.n372 B.n371 10.6151
R1625 B.n373 B.n372 10.6151
R1626 B.n373 B.n176 10.6151
R1627 B.n377 B.n176 10.6151
R1628 B.n378 B.n377 10.6151
R1629 B.n380 B.n172 10.6151
R1630 B.n384 B.n172 10.6151
R1631 B.n385 B.n384 10.6151
R1632 B.n386 B.n385 10.6151
R1633 B.n386 B.n170 10.6151
R1634 B.n390 B.n170 10.6151
R1635 B.n391 B.n390 10.6151
R1636 B.n392 B.n391 10.6151
R1637 B.n396 B.n395 10.6151
R1638 B.n397 B.n396 10.6151
R1639 B.n397 B.n164 10.6151
R1640 B.n401 B.n164 10.6151
R1641 B.n402 B.n401 10.6151
R1642 B.n403 B.n402 10.6151
R1643 B.n403 B.n162 10.6151
R1644 B.n407 B.n162 10.6151
R1645 B.n408 B.n407 10.6151
R1646 B.n409 B.n408 10.6151
R1647 B.n409 B.n160 10.6151
R1648 B.n413 B.n160 10.6151
R1649 B.n414 B.n413 10.6151
R1650 B.n415 B.n414 10.6151
R1651 B.n415 B.n158 10.6151
R1652 B.n419 B.n158 10.6151
R1653 B.n420 B.n419 10.6151
R1654 B.n421 B.n420 10.6151
R1655 B.n421 B.n156 10.6151
R1656 B.n425 B.n156 10.6151
R1657 B.n426 B.n425 10.6151
R1658 B.n343 B.n186 10.6151
R1659 B.n343 B.n342 10.6151
R1660 B.n342 B.n341 10.6151
R1661 B.n341 B.n188 10.6151
R1662 B.n337 B.n188 10.6151
R1663 B.n337 B.n336 10.6151
R1664 B.n336 B.n335 10.6151
R1665 B.n335 B.n190 10.6151
R1666 B.n331 B.n190 10.6151
R1667 B.n331 B.n330 10.6151
R1668 B.n330 B.n329 10.6151
R1669 B.n329 B.n192 10.6151
R1670 B.n325 B.n192 10.6151
R1671 B.n325 B.n324 10.6151
R1672 B.n324 B.n323 10.6151
R1673 B.n323 B.n194 10.6151
R1674 B.n319 B.n194 10.6151
R1675 B.n319 B.n318 10.6151
R1676 B.n318 B.n317 10.6151
R1677 B.n317 B.n196 10.6151
R1678 B.n313 B.n196 10.6151
R1679 B.n313 B.n312 10.6151
R1680 B.n312 B.n311 10.6151
R1681 B.n311 B.n198 10.6151
R1682 B.n307 B.n198 10.6151
R1683 B.n307 B.n306 10.6151
R1684 B.n306 B.n305 10.6151
R1685 B.n305 B.n200 10.6151
R1686 B.n301 B.n200 10.6151
R1687 B.n301 B.n300 10.6151
R1688 B.n300 B.n299 10.6151
R1689 B.n299 B.n202 10.6151
R1690 B.n295 B.n202 10.6151
R1691 B.n295 B.n294 10.6151
R1692 B.n294 B.n293 10.6151
R1693 B.n293 B.n204 10.6151
R1694 B.n289 B.n204 10.6151
R1695 B.n289 B.n288 10.6151
R1696 B.n288 B.n287 10.6151
R1697 B.n287 B.n206 10.6151
R1698 B.n283 B.n206 10.6151
R1699 B.n283 B.n282 10.6151
R1700 B.n282 B.n281 10.6151
R1701 B.n281 B.n208 10.6151
R1702 B.n277 B.n208 10.6151
R1703 B.n277 B.n276 10.6151
R1704 B.n276 B.n275 10.6151
R1705 B.n275 B.n210 10.6151
R1706 B.n271 B.n210 10.6151
R1707 B.n271 B.n270 10.6151
R1708 B.n270 B.n269 10.6151
R1709 B.n269 B.n212 10.6151
R1710 B.n265 B.n212 10.6151
R1711 B.n265 B.n264 10.6151
R1712 B.n264 B.n263 10.6151
R1713 B.n263 B.n214 10.6151
R1714 B.n259 B.n214 10.6151
R1715 B.n259 B.n258 10.6151
R1716 B.n258 B.n257 10.6151
R1717 B.n257 B.n216 10.6151
R1718 B.n253 B.n216 10.6151
R1719 B.n253 B.n252 10.6151
R1720 B.n252 B.n251 10.6151
R1721 B.n251 B.n218 10.6151
R1722 B.n247 B.n218 10.6151
R1723 B.n247 B.n246 10.6151
R1724 B.n246 B.n245 10.6151
R1725 B.n245 B.n220 10.6151
R1726 B.n241 B.n220 10.6151
R1727 B.n241 B.n240 10.6151
R1728 B.n240 B.n239 10.6151
R1729 B.n239 B.n222 10.6151
R1730 B.n235 B.n222 10.6151
R1731 B.n235 B.n234 10.6151
R1732 B.n234 B.n233 10.6151
R1733 B.n233 B.n224 10.6151
R1734 B.n229 B.n224 10.6151
R1735 B.n229 B.n228 10.6151
R1736 B.n228 B.n227 10.6151
R1737 B.n227 B.n0 10.6151
R1738 B.n871 B.n1 10.6151
R1739 B.n871 B.n870 10.6151
R1740 B.n870 B.n869 10.6151
R1741 B.n869 B.n4 10.6151
R1742 B.n865 B.n4 10.6151
R1743 B.n865 B.n864 10.6151
R1744 B.n864 B.n863 10.6151
R1745 B.n863 B.n6 10.6151
R1746 B.n859 B.n6 10.6151
R1747 B.n859 B.n858 10.6151
R1748 B.n858 B.n857 10.6151
R1749 B.n857 B.n8 10.6151
R1750 B.n853 B.n8 10.6151
R1751 B.n853 B.n852 10.6151
R1752 B.n852 B.n851 10.6151
R1753 B.n851 B.n10 10.6151
R1754 B.n847 B.n10 10.6151
R1755 B.n847 B.n846 10.6151
R1756 B.n846 B.n845 10.6151
R1757 B.n845 B.n12 10.6151
R1758 B.n841 B.n12 10.6151
R1759 B.n841 B.n840 10.6151
R1760 B.n840 B.n839 10.6151
R1761 B.n839 B.n14 10.6151
R1762 B.n835 B.n14 10.6151
R1763 B.n835 B.n834 10.6151
R1764 B.n834 B.n833 10.6151
R1765 B.n833 B.n16 10.6151
R1766 B.n829 B.n16 10.6151
R1767 B.n829 B.n828 10.6151
R1768 B.n828 B.n827 10.6151
R1769 B.n827 B.n18 10.6151
R1770 B.n823 B.n18 10.6151
R1771 B.n823 B.n822 10.6151
R1772 B.n822 B.n821 10.6151
R1773 B.n821 B.n20 10.6151
R1774 B.n817 B.n20 10.6151
R1775 B.n817 B.n816 10.6151
R1776 B.n816 B.n815 10.6151
R1777 B.n815 B.n22 10.6151
R1778 B.n811 B.n22 10.6151
R1779 B.n811 B.n810 10.6151
R1780 B.n810 B.n809 10.6151
R1781 B.n809 B.n24 10.6151
R1782 B.n805 B.n24 10.6151
R1783 B.n805 B.n804 10.6151
R1784 B.n804 B.n803 10.6151
R1785 B.n803 B.n26 10.6151
R1786 B.n799 B.n26 10.6151
R1787 B.n799 B.n798 10.6151
R1788 B.n798 B.n797 10.6151
R1789 B.n797 B.n28 10.6151
R1790 B.n793 B.n28 10.6151
R1791 B.n793 B.n792 10.6151
R1792 B.n792 B.n791 10.6151
R1793 B.n791 B.n30 10.6151
R1794 B.n787 B.n30 10.6151
R1795 B.n787 B.n786 10.6151
R1796 B.n786 B.n785 10.6151
R1797 B.n785 B.n32 10.6151
R1798 B.n781 B.n32 10.6151
R1799 B.n781 B.n780 10.6151
R1800 B.n780 B.n779 10.6151
R1801 B.n779 B.n34 10.6151
R1802 B.n775 B.n34 10.6151
R1803 B.n775 B.n774 10.6151
R1804 B.n774 B.n773 10.6151
R1805 B.n773 B.n36 10.6151
R1806 B.n769 B.n36 10.6151
R1807 B.n769 B.n768 10.6151
R1808 B.n768 B.n767 10.6151
R1809 B.n767 B.n38 10.6151
R1810 B.n763 B.n38 10.6151
R1811 B.n763 B.n762 10.6151
R1812 B.n762 B.n761 10.6151
R1813 B.n761 B.n40 10.6151
R1814 B.n757 B.n40 10.6151
R1815 B.n757 B.n756 10.6151
R1816 B.n756 B.n755 10.6151
R1817 B.n755 B.n42 10.6151
R1818 B.n719 B.n718 6.5566
R1819 B.n706 B.n62 6.5566
R1820 B.n380 B.n379 6.5566
R1821 B.n392 B.n168 6.5566
R1822 B.n720 B.n719 4.05904
R1823 B.n703 B.n62 4.05904
R1824 B.n379 B.n378 4.05904
R1825 B.n395 B.n168 4.05904
R1826 B.n875 B.n0 2.81026
R1827 B.n875 B.n1 2.81026
R1828 VN.n110 VN.n109 161.3
R1829 VN.n108 VN.n57 161.3
R1830 VN.n107 VN.n106 161.3
R1831 VN.n105 VN.n58 161.3
R1832 VN.n104 VN.n103 161.3
R1833 VN.n102 VN.n59 161.3
R1834 VN.n101 VN.n100 161.3
R1835 VN.n99 VN.n60 161.3
R1836 VN.n98 VN.n97 161.3
R1837 VN.n95 VN.n61 161.3
R1838 VN.n94 VN.n93 161.3
R1839 VN.n92 VN.n62 161.3
R1840 VN.n91 VN.n90 161.3
R1841 VN.n89 VN.n63 161.3
R1842 VN.n88 VN.n87 161.3
R1843 VN.n86 VN.n64 161.3
R1844 VN.n85 VN.n84 161.3
R1845 VN.n82 VN.n65 161.3
R1846 VN.n81 VN.n80 161.3
R1847 VN.n79 VN.n66 161.3
R1848 VN.n78 VN.n77 161.3
R1849 VN.n76 VN.n67 161.3
R1850 VN.n75 VN.n74 161.3
R1851 VN.n73 VN.n68 161.3
R1852 VN.n72 VN.n71 161.3
R1853 VN.n54 VN.n53 161.3
R1854 VN.n52 VN.n1 161.3
R1855 VN.n51 VN.n50 161.3
R1856 VN.n49 VN.n2 161.3
R1857 VN.n48 VN.n47 161.3
R1858 VN.n46 VN.n3 161.3
R1859 VN.n45 VN.n44 161.3
R1860 VN.n43 VN.n4 161.3
R1861 VN.n42 VN.n41 161.3
R1862 VN.n39 VN.n5 161.3
R1863 VN.n38 VN.n37 161.3
R1864 VN.n36 VN.n6 161.3
R1865 VN.n35 VN.n34 161.3
R1866 VN.n33 VN.n7 161.3
R1867 VN.n32 VN.n31 161.3
R1868 VN.n30 VN.n8 161.3
R1869 VN.n29 VN.n28 161.3
R1870 VN.n26 VN.n9 161.3
R1871 VN.n25 VN.n24 161.3
R1872 VN.n23 VN.n10 161.3
R1873 VN.n22 VN.n21 161.3
R1874 VN.n20 VN.n11 161.3
R1875 VN.n19 VN.n18 161.3
R1876 VN.n17 VN.n12 161.3
R1877 VN.n16 VN.n15 161.3
R1878 VN.n55 VN.n0 89.5781
R1879 VN.n111 VN.n56 89.5781
R1880 VN.n69 VN.t2 65.6271
R1881 VN.n13 VN.t1 65.6271
R1882 VN.n21 VN.n20 56.5193
R1883 VN.n34 VN.n33 56.5193
R1884 VN.n77 VN.n76 56.5193
R1885 VN.n90 VN.n89 56.5193
R1886 VN.n14 VN.n13 56.4597
R1887 VN.n70 VN.n69 56.4597
R1888 VN VN.n111 54.7215
R1889 VN.n47 VN.n46 45.8354
R1890 VN.n103 VN.n102 45.8354
R1891 VN.n47 VN.n2 35.1514
R1892 VN.n103 VN.n58 35.1514
R1893 VN.n14 VN.t0 33.4234
R1894 VN.n27 VN.t9 33.4234
R1895 VN.n40 VN.t6 33.4234
R1896 VN.n0 VN.t5 33.4234
R1897 VN.n70 VN.t3 33.4234
R1898 VN.n83 VN.t4 33.4234
R1899 VN.n96 VN.t8 33.4234
R1900 VN.n56 VN.t7 33.4234
R1901 VN.n15 VN.n12 24.4675
R1902 VN.n19 VN.n12 24.4675
R1903 VN.n20 VN.n19 24.4675
R1904 VN.n21 VN.n10 24.4675
R1905 VN.n25 VN.n10 24.4675
R1906 VN.n26 VN.n25 24.4675
R1907 VN.n28 VN.n8 24.4675
R1908 VN.n32 VN.n8 24.4675
R1909 VN.n33 VN.n32 24.4675
R1910 VN.n34 VN.n6 24.4675
R1911 VN.n38 VN.n6 24.4675
R1912 VN.n39 VN.n38 24.4675
R1913 VN.n41 VN.n4 24.4675
R1914 VN.n45 VN.n4 24.4675
R1915 VN.n46 VN.n45 24.4675
R1916 VN.n51 VN.n2 24.4675
R1917 VN.n52 VN.n51 24.4675
R1918 VN.n53 VN.n52 24.4675
R1919 VN.n76 VN.n75 24.4675
R1920 VN.n75 VN.n68 24.4675
R1921 VN.n71 VN.n68 24.4675
R1922 VN.n89 VN.n88 24.4675
R1923 VN.n88 VN.n64 24.4675
R1924 VN.n84 VN.n64 24.4675
R1925 VN.n82 VN.n81 24.4675
R1926 VN.n81 VN.n66 24.4675
R1927 VN.n77 VN.n66 24.4675
R1928 VN.n102 VN.n101 24.4675
R1929 VN.n101 VN.n60 24.4675
R1930 VN.n97 VN.n60 24.4675
R1931 VN.n95 VN.n94 24.4675
R1932 VN.n94 VN.n62 24.4675
R1933 VN.n90 VN.n62 24.4675
R1934 VN.n109 VN.n108 24.4675
R1935 VN.n108 VN.n107 24.4675
R1936 VN.n107 VN.n58 24.4675
R1937 VN.n15 VN.n14 18.5954
R1938 VN.n40 VN.n39 18.5954
R1939 VN.n71 VN.n70 18.5954
R1940 VN.n96 VN.n95 18.5954
R1941 VN.n27 VN.n26 12.234
R1942 VN.n28 VN.n27 12.234
R1943 VN.n84 VN.n83 12.234
R1944 VN.n83 VN.n82 12.234
R1945 VN.n41 VN.n40 5.87258
R1946 VN.n97 VN.n96 5.87258
R1947 VN.n72 VN.n69 2.5172
R1948 VN.n16 VN.n13 2.5172
R1949 VN.n53 VN.n0 0.48984
R1950 VN.n109 VN.n56 0.48984
R1951 VN.n111 VN.n110 0.354971
R1952 VN.n55 VN.n54 0.354971
R1953 VN VN.n55 0.26696
R1954 VN.n110 VN.n57 0.189894
R1955 VN.n106 VN.n57 0.189894
R1956 VN.n106 VN.n105 0.189894
R1957 VN.n105 VN.n104 0.189894
R1958 VN.n104 VN.n59 0.189894
R1959 VN.n100 VN.n59 0.189894
R1960 VN.n100 VN.n99 0.189894
R1961 VN.n99 VN.n98 0.189894
R1962 VN.n98 VN.n61 0.189894
R1963 VN.n93 VN.n61 0.189894
R1964 VN.n93 VN.n92 0.189894
R1965 VN.n92 VN.n91 0.189894
R1966 VN.n91 VN.n63 0.189894
R1967 VN.n87 VN.n63 0.189894
R1968 VN.n87 VN.n86 0.189894
R1969 VN.n86 VN.n85 0.189894
R1970 VN.n85 VN.n65 0.189894
R1971 VN.n80 VN.n65 0.189894
R1972 VN.n80 VN.n79 0.189894
R1973 VN.n79 VN.n78 0.189894
R1974 VN.n78 VN.n67 0.189894
R1975 VN.n74 VN.n67 0.189894
R1976 VN.n74 VN.n73 0.189894
R1977 VN.n73 VN.n72 0.189894
R1978 VN.n17 VN.n16 0.189894
R1979 VN.n18 VN.n17 0.189894
R1980 VN.n18 VN.n11 0.189894
R1981 VN.n22 VN.n11 0.189894
R1982 VN.n23 VN.n22 0.189894
R1983 VN.n24 VN.n23 0.189894
R1984 VN.n24 VN.n9 0.189894
R1985 VN.n29 VN.n9 0.189894
R1986 VN.n30 VN.n29 0.189894
R1987 VN.n31 VN.n30 0.189894
R1988 VN.n31 VN.n7 0.189894
R1989 VN.n35 VN.n7 0.189894
R1990 VN.n36 VN.n35 0.189894
R1991 VN.n37 VN.n36 0.189894
R1992 VN.n37 VN.n5 0.189894
R1993 VN.n42 VN.n5 0.189894
R1994 VN.n43 VN.n42 0.189894
R1995 VN.n44 VN.n43 0.189894
R1996 VN.n44 VN.n3 0.189894
R1997 VN.n48 VN.n3 0.189894
R1998 VN.n49 VN.n48 0.189894
R1999 VN.n50 VN.n49 0.189894
R2000 VN.n50 VN.n1 0.189894
R2001 VN.n54 VN.n1 0.189894
R2002 VDD2.n53 VDD2.n31 756.745
R2003 VDD2.n22 VDD2.n0 756.745
R2004 VDD2.n54 VDD2.n53 585
R2005 VDD2.n52 VDD2.n51 585
R2006 VDD2.n35 VDD2.n34 585
R2007 VDD2.n46 VDD2.n45 585
R2008 VDD2.n44 VDD2.n43 585
R2009 VDD2.n39 VDD2.n38 585
R2010 VDD2.n8 VDD2.n7 585
R2011 VDD2.n13 VDD2.n12 585
R2012 VDD2.n15 VDD2.n14 585
R2013 VDD2.n4 VDD2.n3 585
R2014 VDD2.n21 VDD2.n20 585
R2015 VDD2.n23 VDD2.n22 585
R2016 VDD2.n40 VDD2.t2 327.856
R2017 VDD2.n9 VDD2.t8 327.856
R2018 VDD2.n53 VDD2.n52 171.744
R2019 VDD2.n52 VDD2.n34 171.744
R2020 VDD2.n45 VDD2.n34 171.744
R2021 VDD2.n45 VDD2.n44 171.744
R2022 VDD2.n44 VDD2.n38 171.744
R2023 VDD2.n13 VDD2.n7 171.744
R2024 VDD2.n14 VDD2.n13 171.744
R2025 VDD2.n14 VDD2.n3 171.744
R2026 VDD2.n21 VDD2.n3 171.744
R2027 VDD2.n22 VDD2.n21 171.744
R2028 VDD2.n30 VDD2.n29 99.7517
R2029 VDD2 VDD2.n61 99.7489
R2030 VDD2.n60 VDD2.n59 97.137
R2031 VDD2.n28 VDD2.n27 97.1368
R2032 VDD2.t2 VDD2.n38 85.8723
R2033 VDD2.t8 VDD2.n7 85.8723
R2034 VDD2.n28 VDD2.n26 52.2305
R2035 VDD2.n58 VDD2.n57 48.6702
R2036 VDD2.n58 VDD2.n30 45.17
R2037 VDD2.n40 VDD2.n39 16.381
R2038 VDD2.n9 VDD2.n8 16.381
R2039 VDD2.n43 VDD2.n42 12.8005
R2040 VDD2.n12 VDD2.n11 12.8005
R2041 VDD2.n46 VDD2.n37 12.0247
R2042 VDD2.n15 VDD2.n6 12.0247
R2043 VDD2.n47 VDD2.n35 11.249
R2044 VDD2.n16 VDD2.n4 11.249
R2045 VDD2.n51 VDD2.n50 10.4732
R2046 VDD2.n20 VDD2.n19 10.4732
R2047 VDD2.n54 VDD2.n33 9.69747
R2048 VDD2.n23 VDD2.n2 9.69747
R2049 VDD2.n57 VDD2.n56 9.45567
R2050 VDD2.n26 VDD2.n25 9.45567
R2051 VDD2.n56 VDD2.n55 9.3005
R2052 VDD2.n33 VDD2.n32 9.3005
R2053 VDD2.n50 VDD2.n49 9.3005
R2054 VDD2.n48 VDD2.n47 9.3005
R2055 VDD2.n37 VDD2.n36 9.3005
R2056 VDD2.n42 VDD2.n41 9.3005
R2057 VDD2.n25 VDD2.n24 9.3005
R2058 VDD2.n2 VDD2.n1 9.3005
R2059 VDD2.n19 VDD2.n18 9.3005
R2060 VDD2.n17 VDD2.n16 9.3005
R2061 VDD2.n6 VDD2.n5 9.3005
R2062 VDD2.n11 VDD2.n10 9.3005
R2063 VDD2.n55 VDD2.n31 8.92171
R2064 VDD2.n24 VDD2.n0 8.92171
R2065 VDD2.n61 VDD2.t6 6.16843
R2066 VDD2.n61 VDD2.t7 6.16843
R2067 VDD2.n59 VDD2.t1 6.16843
R2068 VDD2.n59 VDD2.t5 6.16843
R2069 VDD2.n29 VDD2.t3 6.16843
R2070 VDD2.n29 VDD2.t4 6.16843
R2071 VDD2.n27 VDD2.t9 6.16843
R2072 VDD2.n27 VDD2.t0 6.16843
R2073 VDD2.n57 VDD2.n31 5.04292
R2074 VDD2.n26 VDD2.n0 5.04292
R2075 VDD2.n55 VDD2.n54 4.26717
R2076 VDD2.n24 VDD2.n23 4.26717
R2077 VDD2.n41 VDD2.n40 3.71853
R2078 VDD2.n10 VDD2.n9 3.71853
R2079 VDD2.n60 VDD2.n58 3.56084
R2080 VDD2.n51 VDD2.n33 3.49141
R2081 VDD2.n20 VDD2.n2 3.49141
R2082 VDD2.n50 VDD2.n35 2.71565
R2083 VDD2.n19 VDD2.n4 2.71565
R2084 VDD2.n47 VDD2.n46 1.93989
R2085 VDD2.n16 VDD2.n15 1.93989
R2086 VDD2.n43 VDD2.n37 1.16414
R2087 VDD2.n12 VDD2.n6 1.16414
R2088 VDD2 VDD2.n60 0.948776
R2089 VDD2.n30 VDD2.n28 0.83524
R2090 VDD2.n42 VDD2.n39 0.388379
R2091 VDD2.n11 VDD2.n8 0.388379
R2092 VDD2.n56 VDD2.n32 0.155672
R2093 VDD2.n49 VDD2.n32 0.155672
R2094 VDD2.n49 VDD2.n48 0.155672
R2095 VDD2.n48 VDD2.n36 0.155672
R2096 VDD2.n41 VDD2.n36 0.155672
R2097 VDD2.n10 VDD2.n5 0.155672
R2098 VDD2.n17 VDD2.n5 0.155672
R2099 VDD2.n18 VDD2.n17 0.155672
R2100 VDD2.n18 VDD2.n1 0.155672
R2101 VDD2.n25 VDD2.n1 0.155672
C0 VTAIL w_n5926_n2022# 2.46954f
C1 VTAIL VP 7.09903f
C2 w_n5926_n2022# VDD1 2.78278f
C3 VDD1 VP 5.88435f
C4 VTAIL VDD1 8.40481f
C5 VDD2 w_n5926_n2022# 2.98843f
C6 VDD2 VP 0.740374f
C7 VDD2 VTAIL 8.465799f
C8 VDD2 VDD1 2.95556f
C9 VN B 1.57581f
C10 w_n5926_n2022# B 10.696401f
C11 B VP 2.88602f
C12 VN w_n5926_n2022# 12.9438f
C13 VN VP 8.92399f
C14 VTAIL B 2.54901f
C15 VTAIL VN 7.08466f
C16 B VDD1 2.40241f
C17 VN VDD1 0.156081f
C18 VDD2 B 2.56726f
C19 VDD2 VN 5.30751f
C20 w_n5926_n2022# VP 13.719f
C21 VDD2 VSUBS 2.5864f
C22 VDD1 VSUBS 2.325829f
C23 VTAIL VSUBS 0.795755f
C24 VN VSUBS 9.41643f
C25 VP VSUBS 5.107214f
C26 B VSUBS 5.894802f
C27 w_n5926_n2022# VSUBS 0.149975p
C28 VDD2.n0 VSUBS 0.039358f
C29 VDD2.n1 VSUBS 0.036666f
C30 VDD2.n2 VSUBS 0.019703f
C31 VDD2.n3 VSUBS 0.04657f
C32 VDD2.n4 VSUBS 0.020862f
C33 VDD2.n5 VSUBS 0.036666f
C34 VDD2.n6 VSUBS 0.019703f
C35 VDD2.n7 VSUBS 0.034928f
C36 VDD2.n8 VSUBS 0.029581f
C37 VDD2.t8 VSUBS 0.100385f
C38 VDD2.n9 VSUBS 0.154644f
C39 VDD2.n10 VSUBS 0.718665f
C40 VDD2.n11 VSUBS 0.019703f
C41 VDD2.n12 VSUBS 0.020862f
C42 VDD2.n13 VSUBS 0.04657f
C43 VDD2.n14 VSUBS 0.04657f
C44 VDD2.n15 VSUBS 0.020862f
C45 VDD2.n16 VSUBS 0.019703f
C46 VDD2.n17 VSUBS 0.036666f
C47 VDD2.n18 VSUBS 0.036666f
C48 VDD2.n19 VSUBS 0.019703f
C49 VDD2.n20 VSUBS 0.020862f
C50 VDD2.n21 VSUBS 0.04657f
C51 VDD2.n22 VSUBS 0.109572f
C52 VDD2.n23 VSUBS 0.020862f
C53 VDD2.n24 VSUBS 0.019703f
C54 VDD2.n25 VSUBS 0.084251f
C55 VDD2.n26 VSUBS 0.113734f
C56 VDD2.t9 VSUBS 0.152696f
C57 VDD2.t0 VSUBS 0.152696f
C58 VDD2.n27 VSUBS 0.974064f
C59 VDD2.n28 VSUBS 1.54993f
C60 VDD2.t3 VSUBS 0.152696f
C61 VDD2.t4 VSUBS 0.152696f
C62 VDD2.n29 VSUBS 1.00858f
C63 VDD2.n30 VSUBS 4.846799f
C64 VDD2.n31 VSUBS 0.039358f
C65 VDD2.n32 VSUBS 0.036666f
C66 VDD2.n33 VSUBS 0.019703f
C67 VDD2.n34 VSUBS 0.04657f
C68 VDD2.n35 VSUBS 0.020862f
C69 VDD2.n36 VSUBS 0.036666f
C70 VDD2.n37 VSUBS 0.019703f
C71 VDD2.n38 VSUBS 0.034928f
C72 VDD2.n39 VSUBS 0.029581f
C73 VDD2.t2 VSUBS 0.100385f
C74 VDD2.n40 VSUBS 0.154644f
C75 VDD2.n41 VSUBS 0.718665f
C76 VDD2.n42 VSUBS 0.019703f
C77 VDD2.n43 VSUBS 0.020862f
C78 VDD2.n44 VSUBS 0.04657f
C79 VDD2.n45 VSUBS 0.04657f
C80 VDD2.n46 VSUBS 0.020862f
C81 VDD2.n47 VSUBS 0.019703f
C82 VDD2.n48 VSUBS 0.036666f
C83 VDD2.n49 VSUBS 0.036666f
C84 VDD2.n50 VSUBS 0.019703f
C85 VDD2.n51 VSUBS 0.020862f
C86 VDD2.n52 VSUBS 0.04657f
C87 VDD2.n53 VSUBS 0.109572f
C88 VDD2.n54 VSUBS 0.020862f
C89 VDD2.n55 VSUBS 0.019703f
C90 VDD2.n56 VSUBS 0.084251f
C91 VDD2.n57 VSUBS 0.080267f
C92 VDD2.n58 VSUBS 4.16157f
C93 VDD2.t1 VSUBS 0.152696f
C94 VDD2.t5 VSUBS 0.152696f
C95 VDD2.n59 VSUBS 0.974069f
C96 VDD2.n60 VSUBS 1.10483f
C97 VDD2.t6 VSUBS 0.152696f
C98 VDD2.t7 VSUBS 0.152696f
C99 VDD2.n61 VSUBS 1.00853f
C100 VN.t5 VSUBS 1.69544f
C101 VN.n0 VSUBS 0.750042f
C102 VN.n1 VSUBS 0.03225f
C103 VN.n2 VSUBS 0.065156f
C104 VN.n3 VSUBS 0.03225f
C105 VN.n4 VSUBS 0.060105f
C106 VN.n5 VSUBS 0.03225f
C107 VN.t6 VSUBS 1.69544f
C108 VN.n6 VSUBS 0.060105f
C109 VN.n7 VSUBS 0.03225f
C110 VN.n8 VSUBS 0.060105f
C111 VN.n9 VSUBS 0.03225f
C112 VN.t9 VSUBS 1.69544f
C113 VN.n10 VSUBS 0.060105f
C114 VN.n11 VSUBS 0.03225f
C115 VN.n12 VSUBS 0.060105f
C116 VN.t1 VSUBS 2.13197f
C117 VN.n13 VSUBS 0.743929f
C118 VN.t0 VSUBS 1.69544f
C119 VN.n14 VSUBS 0.75702f
C120 VN.n15 VSUBS 0.052984f
C121 VN.n16 VSUBS 0.416082f
C122 VN.n17 VSUBS 0.03225f
C123 VN.n18 VSUBS 0.03225f
C124 VN.n19 VSUBS 0.060105f
C125 VN.n20 VSUBS 0.041241f
C126 VN.n21 VSUBS 0.052923f
C127 VN.n22 VSUBS 0.03225f
C128 VN.n23 VSUBS 0.03225f
C129 VN.n24 VSUBS 0.03225f
C130 VN.n25 VSUBS 0.060105f
C131 VN.n26 VSUBS 0.045268f
C132 VN.n27 VSUBS 0.632983f
C133 VN.n28 VSUBS 0.045268f
C134 VN.n29 VSUBS 0.03225f
C135 VN.n30 VSUBS 0.03225f
C136 VN.n31 VSUBS 0.03225f
C137 VN.n32 VSUBS 0.060105f
C138 VN.n33 VSUBS 0.052923f
C139 VN.n34 VSUBS 0.041241f
C140 VN.n35 VSUBS 0.03225f
C141 VN.n36 VSUBS 0.03225f
C142 VN.n37 VSUBS 0.03225f
C143 VN.n38 VSUBS 0.060105f
C144 VN.n39 VSUBS 0.052984f
C145 VN.n40 VSUBS 0.632983f
C146 VN.n41 VSUBS 0.037553f
C147 VN.n42 VSUBS 0.03225f
C148 VN.n43 VSUBS 0.03225f
C149 VN.n44 VSUBS 0.03225f
C150 VN.n45 VSUBS 0.060105f
C151 VN.n46 VSUBS 0.061765f
C152 VN.n47 VSUBS 0.027347f
C153 VN.n48 VSUBS 0.03225f
C154 VN.n49 VSUBS 0.03225f
C155 VN.n50 VSUBS 0.03225f
C156 VN.n51 VSUBS 0.060105f
C157 VN.n52 VSUBS 0.060105f
C158 VN.n53 VSUBS 0.031025f
C159 VN.n54 VSUBS 0.05205f
C160 VN.n55 VSUBS 0.101248f
C161 VN.t7 VSUBS 1.69544f
C162 VN.n56 VSUBS 0.750042f
C163 VN.n57 VSUBS 0.03225f
C164 VN.n58 VSUBS 0.065156f
C165 VN.n59 VSUBS 0.03225f
C166 VN.n60 VSUBS 0.060105f
C167 VN.n61 VSUBS 0.03225f
C168 VN.t8 VSUBS 1.69544f
C169 VN.n62 VSUBS 0.060105f
C170 VN.n63 VSUBS 0.03225f
C171 VN.n64 VSUBS 0.060105f
C172 VN.n65 VSUBS 0.03225f
C173 VN.t4 VSUBS 1.69544f
C174 VN.n66 VSUBS 0.060105f
C175 VN.n67 VSUBS 0.03225f
C176 VN.n68 VSUBS 0.060105f
C177 VN.t2 VSUBS 2.13197f
C178 VN.n69 VSUBS 0.743929f
C179 VN.t3 VSUBS 1.69544f
C180 VN.n70 VSUBS 0.75702f
C181 VN.n71 VSUBS 0.052984f
C182 VN.n72 VSUBS 0.416082f
C183 VN.n73 VSUBS 0.03225f
C184 VN.n74 VSUBS 0.03225f
C185 VN.n75 VSUBS 0.060105f
C186 VN.n76 VSUBS 0.041241f
C187 VN.n77 VSUBS 0.052923f
C188 VN.n78 VSUBS 0.03225f
C189 VN.n79 VSUBS 0.03225f
C190 VN.n80 VSUBS 0.03225f
C191 VN.n81 VSUBS 0.060105f
C192 VN.n82 VSUBS 0.045268f
C193 VN.n83 VSUBS 0.632983f
C194 VN.n84 VSUBS 0.045268f
C195 VN.n85 VSUBS 0.03225f
C196 VN.n86 VSUBS 0.03225f
C197 VN.n87 VSUBS 0.03225f
C198 VN.n88 VSUBS 0.060105f
C199 VN.n89 VSUBS 0.052923f
C200 VN.n90 VSUBS 0.041241f
C201 VN.n91 VSUBS 0.03225f
C202 VN.n92 VSUBS 0.03225f
C203 VN.n93 VSUBS 0.03225f
C204 VN.n94 VSUBS 0.060105f
C205 VN.n95 VSUBS 0.052984f
C206 VN.n96 VSUBS 0.632983f
C207 VN.n97 VSUBS 0.037553f
C208 VN.n98 VSUBS 0.03225f
C209 VN.n99 VSUBS 0.03225f
C210 VN.n100 VSUBS 0.03225f
C211 VN.n101 VSUBS 0.060105f
C212 VN.n102 VSUBS 0.061765f
C213 VN.n103 VSUBS 0.027347f
C214 VN.n104 VSUBS 0.03225f
C215 VN.n105 VSUBS 0.03225f
C216 VN.n106 VSUBS 0.03225f
C217 VN.n107 VSUBS 0.060105f
C218 VN.n108 VSUBS 0.060105f
C219 VN.n109 VSUBS 0.031025f
C220 VN.n110 VSUBS 0.05205f
C221 VN.n111 VSUBS 2.11001f
C222 B.n0 VSUBS 0.007653f
C223 B.n1 VSUBS 0.007653f
C224 B.n2 VSUBS 0.012103f
C225 B.n3 VSUBS 0.012103f
C226 B.n4 VSUBS 0.012103f
C227 B.n5 VSUBS 0.012103f
C228 B.n6 VSUBS 0.012103f
C229 B.n7 VSUBS 0.012103f
C230 B.n8 VSUBS 0.012103f
C231 B.n9 VSUBS 0.012103f
C232 B.n10 VSUBS 0.012103f
C233 B.n11 VSUBS 0.012103f
C234 B.n12 VSUBS 0.012103f
C235 B.n13 VSUBS 0.012103f
C236 B.n14 VSUBS 0.012103f
C237 B.n15 VSUBS 0.012103f
C238 B.n16 VSUBS 0.012103f
C239 B.n17 VSUBS 0.012103f
C240 B.n18 VSUBS 0.012103f
C241 B.n19 VSUBS 0.012103f
C242 B.n20 VSUBS 0.012103f
C243 B.n21 VSUBS 0.012103f
C244 B.n22 VSUBS 0.012103f
C245 B.n23 VSUBS 0.012103f
C246 B.n24 VSUBS 0.012103f
C247 B.n25 VSUBS 0.012103f
C248 B.n26 VSUBS 0.012103f
C249 B.n27 VSUBS 0.012103f
C250 B.n28 VSUBS 0.012103f
C251 B.n29 VSUBS 0.012103f
C252 B.n30 VSUBS 0.012103f
C253 B.n31 VSUBS 0.012103f
C254 B.n32 VSUBS 0.012103f
C255 B.n33 VSUBS 0.012103f
C256 B.n34 VSUBS 0.012103f
C257 B.n35 VSUBS 0.012103f
C258 B.n36 VSUBS 0.012103f
C259 B.n37 VSUBS 0.012103f
C260 B.n38 VSUBS 0.012103f
C261 B.n39 VSUBS 0.012103f
C262 B.n40 VSUBS 0.012103f
C263 B.n41 VSUBS 0.012103f
C264 B.n42 VSUBS 0.028308f
C265 B.n43 VSUBS 0.012103f
C266 B.n44 VSUBS 0.012103f
C267 B.n45 VSUBS 0.012103f
C268 B.n46 VSUBS 0.012103f
C269 B.n47 VSUBS 0.012103f
C270 B.n48 VSUBS 0.012103f
C271 B.n49 VSUBS 0.012103f
C272 B.n50 VSUBS 0.012103f
C273 B.n51 VSUBS 0.012103f
C274 B.n52 VSUBS 0.012103f
C275 B.n53 VSUBS 0.012103f
C276 B.t8 VSUBS 0.133242f
C277 B.t7 VSUBS 0.189974f
C278 B.t6 VSUBS 1.67203f
C279 B.n54 VSUBS 0.316231f
C280 B.n55 VSUBS 0.254932f
C281 B.n56 VSUBS 0.012103f
C282 B.n57 VSUBS 0.012103f
C283 B.n58 VSUBS 0.012103f
C284 B.n59 VSUBS 0.012103f
C285 B.t5 VSUBS 0.133244f
C286 B.t4 VSUBS 0.189976f
C287 B.t3 VSUBS 1.67203f
C288 B.n60 VSUBS 0.316229f
C289 B.n61 VSUBS 0.254929f
C290 B.n62 VSUBS 0.028041f
C291 B.n63 VSUBS 0.012103f
C292 B.n64 VSUBS 0.012103f
C293 B.n65 VSUBS 0.012103f
C294 B.n66 VSUBS 0.012103f
C295 B.n67 VSUBS 0.012103f
C296 B.n68 VSUBS 0.012103f
C297 B.n69 VSUBS 0.012103f
C298 B.n70 VSUBS 0.012103f
C299 B.n71 VSUBS 0.012103f
C300 B.n72 VSUBS 0.012103f
C301 B.n73 VSUBS 0.02936f
C302 B.n74 VSUBS 0.012103f
C303 B.n75 VSUBS 0.012103f
C304 B.n76 VSUBS 0.012103f
C305 B.n77 VSUBS 0.012103f
C306 B.n78 VSUBS 0.012103f
C307 B.n79 VSUBS 0.012103f
C308 B.n80 VSUBS 0.012103f
C309 B.n81 VSUBS 0.012103f
C310 B.n82 VSUBS 0.012103f
C311 B.n83 VSUBS 0.012103f
C312 B.n84 VSUBS 0.012103f
C313 B.n85 VSUBS 0.012103f
C314 B.n86 VSUBS 0.012103f
C315 B.n87 VSUBS 0.012103f
C316 B.n88 VSUBS 0.012103f
C317 B.n89 VSUBS 0.012103f
C318 B.n90 VSUBS 0.012103f
C319 B.n91 VSUBS 0.012103f
C320 B.n92 VSUBS 0.012103f
C321 B.n93 VSUBS 0.012103f
C322 B.n94 VSUBS 0.012103f
C323 B.n95 VSUBS 0.012103f
C324 B.n96 VSUBS 0.012103f
C325 B.n97 VSUBS 0.012103f
C326 B.n98 VSUBS 0.012103f
C327 B.n99 VSUBS 0.012103f
C328 B.n100 VSUBS 0.012103f
C329 B.n101 VSUBS 0.012103f
C330 B.n102 VSUBS 0.012103f
C331 B.n103 VSUBS 0.012103f
C332 B.n104 VSUBS 0.012103f
C333 B.n105 VSUBS 0.012103f
C334 B.n106 VSUBS 0.012103f
C335 B.n107 VSUBS 0.012103f
C336 B.n108 VSUBS 0.012103f
C337 B.n109 VSUBS 0.012103f
C338 B.n110 VSUBS 0.012103f
C339 B.n111 VSUBS 0.012103f
C340 B.n112 VSUBS 0.012103f
C341 B.n113 VSUBS 0.012103f
C342 B.n114 VSUBS 0.012103f
C343 B.n115 VSUBS 0.012103f
C344 B.n116 VSUBS 0.012103f
C345 B.n117 VSUBS 0.012103f
C346 B.n118 VSUBS 0.012103f
C347 B.n119 VSUBS 0.012103f
C348 B.n120 VSUBS 0.012103f
C349 B.n121 VSUBS 0.012103f
C350 B.n122 VSUBS 0.012103f
C351 B.n123 VSUBS 0.012103f
C352 B.n124 VSUBS 0.012103f
C353 B.n125 VSUBS 0.012103f
C354 B.n126 VSUBS 0.012103f
C355 B.n127 VSUBS 0.012103f
C356 B.n128 VSUBS 0.012103f
C357 B.n129 VSUBS 0.012103f
C358 B.n130 VSUBS 0.012103f
C359 B.n131 VSUBS 0.012103f
C360 B.n132 VSUBS 0.012103f
C361 B.n133 VSUBS 0.012103f
C362 B.n134 VSUBS 0.012103f
C363 B.n135 VSUBS 0.012103f
C364 B.n136 VSUBS 0.012103f
C365 B.n137 VSUBS 0.012103f
C366 B.n138 VSUBS 0.012103f
C367 B.n139 VSUBS 0.012103f
C368 B.n140 VSUBS 0.012103f
C369 B.n141 VSUBS 0.012103f
C370 B.n142 VSUBS 0.012103f
C371 B.n143 VSUBS 0.012103f
C372 B.n144 VSUBS 0.012103f
C373 B.n145 VSUBS 0.012103f
C374 B.n146 VSUBS 0.012103f
C375 B.n147 VSUBS 0.012103f
C376 B.n148 VSUBS 0.012103f
C377 B.n149 VSUBS 0.012103f
C378 B.n150 VSUBS 0.012103f
C379 B.n151 VSUBS 0.012103f
C380 B.n152 VSUBS 0.012103f
C381 B.n153 VSUBS 0.012103f
C382 B.n154 VSUBS 0.012103f
C383 B.n155 VSUBS 0.02936f
C384 B.n156 VSUBS 0.012103f
C385 B.n157 VSUBS 0.012103f
C386 B.n158 VSUBS 0.012103f
C387 B.n159 VSUBS 0.012103f
C388 B.n160 VSUBS 0.012103f
C389 B.n161 VSUBS 0.012103f
C390 B.n162 VSUBS 0.012103f
C391 B.n163 VSUBS 0.012103f
C392 B.n164 VSUBS 0.012103f
C393 B.n165 VSUBS 0.012103f
C394 B.t1 VSUBS 0.133244f
C395 B.t2 VSUBS 0.189976f
C396 B.t0 VSUBS 1.67203f
C397 B.n166 VSUBS 0.316229f
C398 B.n167 VSUBS 0.254929f
C399 B.n168 VSUBS 0.028041f
C400 B.n169 VSUBS 0.012103f
C401 B.n170 VSUBS 0.012103f
C402 B.n171 VSUBS 0.012103f
C403 B.n172 VSUBS 0.012103f
C404 B.n173 VSUBS 0.012103f
C405 B.t10 VSUBS 0.133242f
C406 B.t11 VSUBS 0.189974f
C407 B.t9 VSUBS 1.67203f
C408 B.n174 VSUBS 0.316231f
C409 B.n175 VSUBS 0.254932f
C410 B.n176 VSUBS 0.012103f
C411 B.n177 VSUBS 0.012103f
C412 B.n178 VSUBS 0.012103f
C413 B.n179 VSUBS 0.012103f
C414 B.n180 VSUBS 0.012103f
C415 B.n181 VSUBS 0.012103f
C416 B.n182 VSUBS 0.012103f
C417 B.n183 VSUBS 0.012103f
C418 B.n184 VSUBS 0.012103f
C419 B.n185 VSUBS 0.012103f
C420 B.n186 VSUBS 0.028308f
C421 B.n187 VSUBS 0.012103f
C422 B.n188 VSUBS 0.012103f
C423 B.n189 VSUBS 0.012103f
C424 B.n190 VSUBS 0.012103f
C425 B.n191 VSUBS 0.012103f
C426 B.n192 VSUBS 0.012103f
C427 B.n193 VSUBS 0.012103f
C428 B.n194 VSUBS 0.012103f
C429 B.n195 VSUBS 0.012103f
C430 B.n196 VSUBS 0.012103f
C431 B.n197 VSUBS 0.012103f
C432 B.n198 VSUBS 0.012103f
C433 B.n199 VSUBS 0.012103f
C434 B.n200 VSUBS 0.012103f
C435 B.n201 VSUBS 0.012103f
C436 B.n202 VSUBS 0.012103f
C437 B.n203 VSUBS 0.012103f
C438 B.n204 VSUBS 0.012103f
C439 B.n205 VSUBS 0.012103f
C440 B.n206 VSUBS 0.012103f
C441 B.n207 VSUBS 0.012103f
C442 B.n208 VSUBS 0.012103f
C443 B.n209 VSUBS 0.012103f
C444 B.n210 VSUBS 0.012103f
C445 B.n211 VSUBS 0.012103f
C446 B.n212 VSUBS 0.012103f
C447 B.n213 VSUBS 0.012103f
C448 B.n214 VSUBS 0.012103f
C449 B.n215 VSUBS 0.012103f
C450 B.n216 VSUBS 0.012103f
C451 B.n217 VSUBS 0.012103f
C452 B.n218 VSUBS 0.012103f
C453 B.n219 VSUBS 0.012103f
C454 B.n220 VSUBS 0.012103f
C455 B.n221 VSUBS 0.012103f
C456 B.n222 VSUBS 0.012103f
C457 B.n223 VSUBS 0.012103f
C458 B.n224 VSUBS 0.012103f
C459 B.n225 VSUBS 0.012103f
C460 B.n226 VSUBS 0.012103f
C461 B.n227 VSUBS 0.012103f
C462 B.n228 VSUBS 0.012103f
C463 B.n229 VSUBS 0.012103f
C464 B.n230 VSUBS 0.012103f
C465 B.n231 VSUBS 0.012103f
C466 B.n232 VSUBS 0.012103f
C467 B.n233 VSUBS 0.012103f
C468 B.n234 VSUBS 0.012103f
C469 B.n235 VSUBS 0.012103f
C470 B.n236 VSUBS 0.012103f
C471 B.n237 VSUBS 0.012103f
C472 B.n238 VSUBS 0.012103f
C473 B.n239 VSUBS 0.012103f
C474 B.n240 VSUBS 0.012103f
C475 B.n241 VSUBS 0.012103f
C476 B.n242 VSUBS 0.012103f
C477 B.n243 VSUBS 0.012103f
C478 B.n244 VSUBS 0.012103f
C479 B.n245 VSUBS 0.012103f
C480 B.n246 VSUBS 0.012103f
C481 B.n247 VSUBS 0.012103f
C482 B.n248 VSUBS 0.012103f
C483 B.n249 VSUBS 0.012103f
C484 B.n250 VSUBS 0.012103f
C485 B.n251 VSUBS 0.012103f
C486 B.n252 VSUBS 0.012103f
C487 B.n253 VSUBS 0.012103f
C488 B.n254 VSUBS 0.012103f
C489 B.n255 VSUBS 0.012103f
C490 B.n256 VSUBS 0.012103f
C491 B.n257 VSUBS 0.012103f
C492 B.n258 VSUBS 0.012103f
C493 B.n259 VSUBS 0.012103f
C494 B.n260 VSUBS 0.012103f
C495 B.n261 VSUBS 0.012103f
C496 B.n262 VSUBS 0.012103f
C497 B.n263 VSUBS 0.012103f
C498 B.n264 VSUBS 0.012103f
C499 B.n265 VSUBS 0.012103f
C500 B.n266 VSUBS 0.012103f
C501 B.n267 VSUBS 0.012103f
C502 B.n268 VSUBS 0.012103f
C503 B.n269 VSUBS 0.012103f
C504 B.n270 VSUBS 0.012103f
C505 B.n271 VSUBS 0.012103f
C506 B.n272 VSUBS 0.012103f
C507 B.n273 VSUBS 0.012103f
C508 B.n274 VSUBS 0.012103f
C509 B.n275 VSUBS 0.012103f
C510 B.n276 VSUBS 0.012103f
C511 B.n277 VSUBS 0.012103f
C512 B.n278 VSUBS 0.012103f
C513 B.n279 VSUBS 0.012103f
C514 B.n280 VSUBS 0.012103f
C515 B.n281 VSUBS 0.012103f
C516 B.n282 VSUBS 0.012103f
C517 B.n283 VSUBS 0.012103f
C518 B.n284 VSUBS 0.012103f
C519 B.n285 VSUBS 0.012103f
C520 B.n286 VSUBS 0.012103f
C521 B.n287 VSUBS 0.012103f
C522 B.n288 VSUBS 0.012103f
C523 B.n289 VSUBS 0.012103f
C524 B.n290 VSUBS 0.012103f
C525 B.n291 VSUBS 0.012103f
C526 B.n292 VSUBS 0.012103f
C527 B.n293 VSUBS 0.012103f
C528 B.n294 VSUBS 0.012103f
C529 B.n295 VSUBS 0.012103f
C530 B.n296 VSUBS 0.012103f
C531 B.n297 VSUBS 0.012103f
C532 B.n298 VSUBS 0.012103f
C533 B.n299 VSUBS 0.012103f
C534 B.n300 VSUBS 0.012103f
C535 B.n301 VSUBS 0.012103f
C536 B.n302 VSUBS 0.012103f
C537 B.n303 VSUBS 0.012103f
C538 B.n304 VSUBS 0.012103f
C539 B.n305 VSUBS 0.012103f
C540 B.n306 VSUBS 0.012103f
C541 B.n307 VSUBS 0.012103f
C542 B.n308 VSUBS 0.012103f
C543 B.n309 VSUBS 0.012103f
C544 B.n310 VSUBS 0.012103f
C545 B.n311 VSUBS 0.012103f
C546 B.n312 VSUBS 0.012103f
C547 B.n313 VSUBS 0.012103f
C548 B.n314 VSUBS 0.012103f
C549 B.n315 VSUBS 0.012103f
C550 B.n316 VSUBS 0.012103f
C551 B.n317 VSUBS 0.012103f
C552 B.n318 VSUBS 0.012103f
C553 B.n319 VSUBS 0.012103f
C554 B.n320 VSUBS 0.012103f
C555 B.n321 VSUBS 0.012103f
C556 B.n322 VSUBS 0.012103f
C557 B.n323 VSUBS 0.012103f
C558 B.n324 VSUBS 0.012103f
C559 B.n325 VSUBS 0.012103f
C560 B.n326 VSUBS 0.012103f
C561 B.n327 VSUBS 0.012103f
C562 B.n328 VSUBS 0.012103f
C563 B.n329 VSUBS 0.012103f
C564 B.n330 VSUBS 0.012103f
C565 B.n331 VSUBS 0.012103f
C566 B.n332 VSUBS 0.012103f
C567 B.n333 VSUBS 0.012103f
C568 B.n334 VSUBS 0.012103f
C569 B.n335 VSUBS 0.012103f
C570 B.n336 VSUBS 0.012103f
C571 B.n337 VSUBS 0.012103f
C572 B.n338 VSUBS 0.012103f
C573 B.n339 VSUBS 0.012103f
C574 B.n340 VSUBS 0.012103f
C575 B.n341 VSUBS 0.012103f
C576 B.n342 VSUBS 0.012103f
C577 B.n343 VSUBS 0.012103f
C578 B.n344 VSUBS 0.012103f
C579 B.n345 VSUBS 0.028308f
C580 B.n346 VSUBS 0.02936f
C581 B.n347 VSUBS 0.02936f
C582 B.n348 VSUBS 0.012103f
C583 B.n349 VSUBS 0.012103f
C584 B.n350 VSUBS 0.012103f
C585 B.n351 VSUBS 0.012103f
C586 B.n352 VSUBS 0.012103f
C587 B.n353 VSUBS 0.012103f
C588 B.n354 VSUBS 0.012103f
C589 B.n355 VSUBS 0.012103f
C590 B.n356 VSUBS 0.012103f
C591 B.n357 VSUBS 0.012103f
C592 B.n358 VSUBS 0.012103f
C593 B.n359 VSUBS 0.012103f
C594 B.n360 VSUBS 0.012103f
C595 B.n361 VSUBS 0.012103f
C596 B.n362 VSUBS 0.012103f
C597 B.n363 VSUBS 0.012103f
C598 B.n364 VSUBS 0.012103f
C599 B.n365 VSUBS 0.012103f
C600 B.n366 VSUBS 0.012103f
C601 B.n367 VSUBS 0.012103f
C602 B.n368 VSUBS 0.012103f
C603 B.n369 VSUBS 0.012103f
C604 B.n370 VSUBS 0.012103f
C605 B.n371 VSUBS 0.012103f
C606 B.n372 VSUBS 0.012103f
C607 B.n373 VSUBS 0.012103f
C608 B.n374 VSUBS 0.012103f
C609 B.n375 VSUBS 0.012103f
C610 B.n376 VSUBS 0.012103f
C611 B.n377 VSUBS 0.012103f
C612 B.n378 VSUBS 0.008365f
C613 B.n379 VSUBS 0.028041f
C614 B.n380 VSUBS 0.009789f
C615 B.n381 VSUBS 0.012103f
C616 B.n382 VSUBS 0.012103f
C617 B.n383 VSUBS 0.012103f
C618 B.n384 VSUBS 0.012103f
C619 B.n385 VSUBS 0.012103f
C620 B.n386 VSUBS 0.012103f
C621 B.n387 VSUBS 0.012103f
C622 B.n388 VSUBS 0.012103f
C623 B.n389 VSUBS 0.012103f
C624 B.n390 VSUBS 0.012103f
C625 B.n391 VSUBS 0.012103f
C626 B.n392 VSUBS 0.009789f
C627 B.n393 VSUBS 0.012103f
C628 B.n394 VSUBS 0.012103f
C629 B.n395 VSUBS 0.008365f
C630 B.n396 VSUBS 0.012103f
C631 B.n397 VSUBS 0.012103f
C632 B.n398 VSUBS 0.012103f
C633 B.n399 VSUBS 0.012103f
C634 B.n400 VSUBS 0.012103f
C635 B.n401 VSUBS 0.012103f
C636 B.n402 VSUBS 0.012103f
C637 B.n403 VSUBS 0.012103f
C638 B.n404 VSUBS 0.012103f
C639 B.n405 VSUBS 0.012103f
C640 B.n406 VSUBS 0.012103f
C641 B.n407 VSUBS 0.012103f
C642 B.n408 VSUBS 0.012103f
C643 B.n409 VSUBS 0.012103f
C644 B.n410 VSUBS 0.012103f
C645 B.n411 VSUBS 0.012103f
C646 B.n412 VSUBS 0.012103f
C647 B.n413 VSUBS 0.012103f
C648 B.n414 VSUBS 0.012103f
C649 B.n415 VSUBS 0.012103f
C650 B.n416 VSUBS 0.012103f
C651 B.n417 VSUBS 0.012103f
C652 B.n418 VSUBS 0.012103f
C653 B.n419 VSUBS 0.012103f
C654 B.n420 VSUBS 0.012103f
C655 B.n421 VSUBS 0.012103f
C656 B.n422 VSUBS 0.012103f
C657 B.n423 VSUBS 0.012103f
C658 B.n424 VSUBS 0.012103f
C659 B.n425 VSUBS 0.012103f
C660 B.n426 VSUBS 0.02936f
C661 B.n427 VSUBS 0.028308f
C662 B.n428 VSUBS 0.028308f
C663 B.n429 VSUBS 0.012103f
C664 B.n430 VSUBS 0.012103f
C665 B.n431 VSUBS 0.012103f
C666 B.n432 VSUBS 0.012103f
C667 B.n433 VSUBS 0.012103f
C668 B.n434 VSUBS 0.012103f
C669 B.n435 VSUBS 0.012103f
C670 B.n436 VSUBS 0.012103f
C671 B.n437 VSUBS 0.012103f
C672 B.n438 VSUBS 0.012103f
C673 B.n439 VSUBS 0.012103f
C674 B.n440 VSUBS 0.012103f
C675 B.n441 VSUBS 0.012103f
C676 B.n442 VSUBS 0.012103f
C677 B.n443 VSUBS 0.012103f
C678 B.n444 VSUBS 0.012103f
C679 B.n445 VSUBS 0.012103f
C680 B.n446 VSUBS 0.012103f
C681 B.n447 VSUBS 0.012103f
C682 B.n448 VSUBS 0.012103f
C683 B.n449 VSUBS 0.012103f
C684 B.n450 VSUBS 0.012103f
C685 B.n451 VSUBS 0.012103f
C686 B.n452 VSUBS 0.012103f
C687 B.n453 VSUBS 0.012103f
C688 B.n454 VSUBS 0.012103f
C689 B.n455 VSUBS 0.012103f
C690 B.n456 VSUBS 0.012103f
C691 B.n457 VSUBS 0.012103f
C692 B.n458 VSUBS 0.012103f
C693 B.n459 VSUBS 0.012103f
C694 B.n460 VSUBS 0.012103f
C695 B.n461 VSUBS 0.012103f
C696 B.n462 VSUBS 0.012103f
C697 B.n463 VSUBS 0.012103f
C698 B.n464 VSUBS 0.012103f
C699 B.n465 VSUBS 0.012103f
C700 B.n466 VSUBS 0.012103f
C701 B.n467 VSUBS 0.012103f
C702 B.n468 VSUBS 0.012103f
C703 B.n469 VSUBS 0.012103f
C704 B.n470 VSUBS 0.012103f
C705 B.n471 VSUBS 0.012103f
C706 B.n472 VSUBS 0.012103f
C707 B.n473 VSUBS 0.012103f
C708 B.n474 VSUBS 0.012103f
C709 B.n475 VSUBS 0.012103f
C710 B.n476 VSUBS 0.012103f
C711 B.n477 VSUBS 0.012103f
C712 B.n478 VSUBS 0.012103f
C713 B.n479 VSUBS 0.012103f
C714 B.n480 VSUBS 0.012103f
C715 B.n481 VSUBS 0.012103f
C716 B.n482 VSUBS 0.012103f
C717 B.n483 VSUBS 0.012103f
C718 B.n484 VSUBS 0.012103f
C719 B.n485 VSUBS 0.012103f
C720 B.n486 VSUBS 0.012103f
C721 B.n487 VSUBS 0.012103f
C722 B.n488 VSUBS 0.012103f
C723 B.n489 VSUBS 0.012103f
C724 B.n490 VSUBS 0.012103f
C725 B.n491 VSUBS 0.012103f
C726 B.n492 VSUBS 0.012103f
C727 B.n493 VSUBS 0.012103f
C728 B.n494 VSUBS 0.012103f
C729 B.n495 VSUBS 0.012103f
C730 B.n496 VSUBS 0.012103f
C731 B.n497 VSUBS 0.012103f
C732 B.n498 VSUBS 0.012103f
C733 B.n499 VSUBS 0.012103f
C734 B.n500 VSUBS 0.012103f
C735 B.n501 VSUBS 0.012103f
C736 B.n502 VSUBS 0.012103f
C737 B.n503 VSUBS 0.012103f
C738 B.n504 VSUBS 0.012103f
C739 B.n505 VSUBS 0.012103f
C740 B.n506 VSUBS 0.012103f
C741 B.n507 VSUBS 0.012103f
C742 B.n508 VSUBS 0.012103f
C743 B.n509 VSUBS 0.012103f
C744 B.n510 VSUBS 0.012103f
C745 B.n511 VSUBS 0.012103f
C746 B.n512 VSUBS 0.012103f
C747 B.n513 VSUBS 0.012103f
C748 B.n514 VSUBS 0.012103f
C749 B.n515 VSUBS 0.012103f
C750 B.n516 VSUBS 0.012103f
C751 B.n517 VSUBS 0.012103f
C752 B.n518 VSUBS 0.012103f
C753 B.n519 VSUBS 0.012103f
C754 B.n520 VSUBS 0.012103f
C755 B.n521 VSUBS 0.012103f
C756 B.n522 VSUBS 0.012103f
C757 B.n523 VSUBS 0.012103f
C758 B.n524 VSUBS 0.012103f
C759 B.n525 VSUBS 0.012103f
C760 B.n526 VSUBS 0.012103f
C761 B.n527 VSUBS 0.012103f
C762 B.n528 VSUBS 0.012103f
C763 B.n529 VSUBS 0.012103f
C764 B.n530 VSUBS 0.012103f
C765 B.n531 VSUBS 0.012103f
C766 B.n532 VSUBS 0.012103f
C767 B.n533 VSUBS 0.012103f
C768 B.n534 VSUBS 0.012103f
C769 B.n535 VSUBS 0.012103f
C770 B.n536 VSUBS 0.012103f
C771 B.n537 VSUBS 0.012103f
C772 B.n538 VSUBS 0.012103f
C773 B.n539 VSUBS 0.012103f
C774 B.n540 VSUBS 0.012103f
C775 B.n541 VSUBS 0.012103f
C776 B.n542 VSUBS 0.012103f
C777 B.n543 VSUBS 0.012103f
C778 B.n544 VSUBS 0.012103f
C779 B.n545 VSUBS 0.012103f
C780 B.n546 VSUBS 0.012103f
C781 B.n547 VSUBS 0.012103f
C782 B.n548 VSUBS 0.012103f
C783 B.n549 VSUBS 0.012103f
C784 B.n550 VSUBS 0.012103f
C785 B.n551 VSUBS 0.012103f
C786 B.n552 VSUBS 0.012103f
C787 B.n553 VSUBS 0.012103f
C788 B.n554 VSUBS 0.012103f
C789 B.n555 VSUBS 0.012103f
C790 B.n556 VSUBS 0.012103f
C791 B.n557 VSUBS 0.012103f
C792 B.n558 VSUBS 0.012103f
C793 B.n559 VSUBS 0.012103f
C794 B.n560 VSUBS 0.012103f
C795 B.n561 VSUBS 0.012103f
C796 B.n562 VSUBS 0.012103f
C797 B.n563 VSUBS 0.012103f
C798 B.n564 VSUBS 0.012103f
C799 B.n565 VSUBS 0.012103f
C800 B.n566 VSUBS 0.012103f
C801 B.n567 VSUBS 0.012103f
C802 B.n568 VSUBS 0.012103f
C803 B.n569 VSUBS 0.012103f
C804 B.n570 VSUBS 0.012103f
C805 B.n571 VSUBS 0.012103f
C806 B.n572 VSUBS 0.012103f
C807 B.n573 VSUBS 0.012103f
C808 B.n574 VSUBS 0.012103f
C809 B.n575 VSUBS 0.012103f
C810 B.n576 VSUBS 0.012103f
C811 B.n577 VSUBS 0.012103f
C812 B.n578 VSUBS 0.012103f
C813 B.n579 VSUBS 0.012103f
C814 B.n580 VSUBS 0.012103f
C815 B.n581 VSUBS 0.012103f
C816 B.n582 VSUBS 0.012103f
C817 B.n583 VSUBS 0.012103f
C818 B.n584 VSUBS 0.012103f
C819 B.n585 VSUBS 0.012103f
C820 B.n586 VSUBS 0.012103f
C821 B.n587 VSUBS 0.012103f
C822 B.n588 VSUBS 0.012103f
C823 B.n589 VSUBS 0.012103f
C824 B.n590 VSUBS 0.012103f
C825 B.n591 VSUBS 0.012103f
C826 B.n592 VSUBS 0.012103f
C827 B.n593 VSUBS 0.012103f
C828 B.n594 VSUBS 0.012103f
C829 B.n595 VSUBS 0.012103f
C830 B.n596 VSUBS 0.012103f
C831 B.n597 VSUBS 0.012103f
C832 B.n598 VSUBS 0.012103f
C833 B.n599 VSUBS 0.012103f
C834 B.n600 VSUBS 0.012103f
C835 B.n601 VSUBS 0.012103f
C836 B.n602 VSUBS 0.012103f
C837 B.n603 VSUBS 0.012103f
C838 B.n604 VSUBS 0.012103f
C839 B.n605 VSUBS 0.012103f
C840 B.n606 VSUBS 0.012103f
C841 B.n607 VSUBS 0.012103f
C842 B.n608 VSUBS 0.012103f
C843 B.n609 VSUBS 0.012103f
C844 B.n610 VSUBS 0.012103f
C845 B.n611 VSUBS 0.012103f
C846 B.n612 VSUBS 0.012103f
C847 B.n613 VSUBS 0.012103f
C848 B.n614 VSUBS 0.012103f
C849 B.n615 VSUBS 0.012103f
C850 B.n616 VSUBS 0.012103f
C851 B.n617 VSUBS 0.012103f
C852 B.n618 VSUBS 0.012103f
C853 B.n619 VSUBS 0.012103f
C854 B.n620 VSUBS 0.012103f
C855 B.n621 VSUBS 0.012103f
C856 B.n622 VSUBS 0.012103f
C857 B.n623 VSUBS 0.012103f
C858 B.n624 VSUBS 0.012103f
C859 B.n625 VSUBS 0.012103f
C860 B.n626 VSUBS 0.012103f
C861 B.n627 VSUBS 0.012103f
C862 B.n628 VSUBS 0.012103f
C863 B.n629 VSUBS 0.012103f
C864 B.n630 VSUBS 0.012103f
C865 B.n631 VSUBS 0.012103f
C866 B.n632 VSUBS 0.012103f
C867 B.n633 VSUBS 0.012103f
C868 B.n634 VSUBS 0.012103f
C869 B.n635 VSUBS 0.012103f
C870 B.n636 VSUBS 0.012103f
C871 B.n637 VSUBS 0.012103f
C872 B.n638 VSUBS 0.012103f
C873 B.n639 VSUBS 0.012103f
C874 B.n640 VSUBS 0.012103f
C875 B.n641 VSUBS 0.012103f
C876 B.n642 VSUBS 0.012103f
C877 B.n643 VSUBS 0.012103f
C878 B.n644 VSUBS 0.012103f
C879 B.n645 VSUBS 0.012103f
C880 B.n646 VSUBS 0.012103f
C881 B.n647 VSUBS 0.012103f
C882 B.n648 VSUBS 0.012103f
C883 B.n649 VSUBS 0.012103f
C884 B.n650 VSUBS 0.012103f
C885 B.n651 VSUBS 0.012103f
C886 B.n652 VSUBS 0.012103f
C887 B.n653 VSUBS 0.012103f
C888 B.n654 VSUBS 0.012103f
C889 B.n655 VSUBS 0.012103f
C890 B.n656 VSUBS 0.012103f
C891 B.n657 VSUBS 0.012103f
C892 B.n658 VSUBS 0.012103f
C893 B.n659 VSUBS 0.012103f
C894 B.n660 VSUBS 0.012103f
C895 B.n661 VSUBS 0.012103f
C896 B.n662 VSUBS 0.012103f
C897 B.n663 VSUBS 0.012103f
C898 B.n664 VSUBS 0.012103f
C899 B.n665 VSUBS 0.012103f
C900 B.n666 VSUBS 0.012103f
C901 B.n667 VSUBS 0.012103f
C902 B.n668 VSUBS 0.012103f
C903 B.n669 VSUBS 0.012103f
C904 B.n670 VSUBS 0.028308f
C905 B.n671 VSUBS 0.029699f
C906 B.n672 VSUBS 0.027968f
C907 B.n673 VSUBS 0.012103f
C908 B.n674 VSUBS 0.012103f
C909 B.n675 VSUBS 0.012103f
C910 B.n676 VSUBS 0.012103f
C911 B.n677 VSUBS 0.012103f
C912 B.n678 VSUBS 0.012103f
C913 B.n679 VSUBS 0.012103f
C914 B.n680 VSUBS 0.012103f
C915 B.n681 VSUBS 0.012103f
C916 B.n682 VSUBS 0.012103f
C917 B.n683 VSUBS 0.012103f
C918 B.n684 VSUBS 0.012103f
C919 B.n685 VSUBS 0.012103f
C920 B.n686 VSUBS 0.012103f
C921 B.n687 VSUBS 0.012103f
C922 B.n688 VSUBS 0.012103f
C923 B.n689 VSUBS 0.012103f
C924 B.n690 VSUBS 0.012103f
C925 B.n691 VSUBS 0.012103f
C926 B.n692 VSUBS 0.012103f
C927 B.n693 VSUBS 0.012103f
C928 B.n694 VSUBS 0.012103f
C929 B.n695 VSUBS 0.012103f
C930 B.n696 VSUBS 0.012103f
C931 B.n697 VSUBS 0.012103f
C932 B.n698 VSUBS 0.012103f
C933 B.n699 VSUBS 0.012103f
C934 B.n700 VSUBS 0.012103f
C935 B.n701 VSUBS 0.012103f
C936 B.n702 VSUBS 0.012103f
C937 B.n703 VSUBS 0.008365f
C938 B.n704 VSUBS 0.012103f
C939 B.n705 VSUBS 0.012103f
C940 B.n706 VSUBS 0.009789f
C941 B.n707 VSUBS 0.012103f
C942 B.n708 VSUBS 0.012103f
C943 B.n709 VSUBS 0.012103f
C944 B.n710 VSUBS 0.012103f
C945 B.n711 VSUBS 0.012103f
C946 B.n712 VSUBS 0.012103f
C947 B.n713 VSUBS 0.012103f
C948 B.n714 VSUBS 0.012103f
C949 B.n715 VSUBS 0.012103f
C950 B.n716 VSUBS 0.012103f
C951 B.n717 VSUBS 0.012103f
C952 B.n718 VSUBS 0.009789f
C953 B.n719 VSUBS 0.028041f
C954 B.n720 VSUBS 0.008365f
C955 B.n721 VSUBS 0.012103f
C956 B.n722 VSUBS 0.012103f
C957 B.n723 VSUBS 0.012103f
C958 B.n724 VSUBS 0.012103f
C959 B.n725 VSUBS 0.012103f
C960 B.n726 VSUBS 0.012103f
C961 B.n727 VSUBS 0.012103f
C962 B.n728 VSUBS 0.012103f
C963 B.n729 VSUBS 0.012103f
C964 B.n730 VSUBS 0.012103f
C965 B.n731 VSUBS 0.012103f
C966 B.n732 VSUBS 0.012103f
C967 B.n733 VSUBS 0.012103f
C968 B.n734 VSUBS 0.012103f
C969 B.n735 VSUBS 0.012103f
C970 B.n736 VSUBS 0.012103f
C971 B.n737 VSUBS 0.012103f
C972 B.n738 VSUBS 0.012103f
C973 B.n739 VSUBS 0.012103f
C974 B.n740 VSUBS 0.012103f
C975 B.n741 VSUBS 0.012103f
C976 B.n742 VSUBS 0.012103f
C977 B.n743 VSUBS 0.012103f
C978 B.n744 VSUBS 0.012103f
C979 B.n745 VSUBS 0.012103f
C980 B.n746 VSUBS 0.012103f
C981 B.n747 VSUBS 0.012103f
C982 B.n748 VSUBS 0.012103f
C983 B.n749 VSUBS 0.012103f
C984 B.n750 VSUBS 0.012103f
C985 B.n751 VSUBS 0.02936f
C986 B.n752 VSUBS 0.02936f
C987 B.n753 VSUBS 0.028308f
C988 B.n754 VSUBS 0.012103f
C989 B.n755 VSUBS 0.012103f
C990 B.n756 VSUBS 0.012103f
C991 B.n757 VSUBS 0.012103f
C992 B.n758 VSUBS 0.012103f
C993 B.n759 VSUBS 0.012103f
C994 B.n760 VSUBS 0.012103f
C995 B.n761 VSUBS 0.012103f
C996 B.n762 VSUBS 0.012103f
C997 B.n763 VSUBS 0.012103f
C998 B.n764 VSUBS 0.012103f
C999 B.n765 VSUBS 0.012103f
C1000 B.n766 VSUBS 0.012103f
C1001 B.n767 VSUBS 0.012103f
C1002 B.n768 VSUBS 0.012103f
C1003 B.n769 VSUBS 0.012103f
C1004 B.n770 VSUBS 0.012103f
C1005 B.n771 VSUBS 0.012103f
C1006 B.n772 VSUBS 0.012103f
C1007 B.n773 VSUBS 0.012103f
C1008 B.n774 VSUBS 0.012103f
C1009 B.n775 VSUBS 0.012103f
C1010 B.n776 VSUBS 0.012103f
C1011 B.n777 VSUBS 0.012103f
C1012 B.n778 VSUBS 0.012103f
C1013 B.n779 VSUBS 0.012103f
C1014 B.n780 VSUBS 0.012103f
C1015 B.n781 VSUBS 0.012103f
C1016 B.n782 VSUBS 0.012103f
C1017 B.n783 VSUBS 0.012103f
C1018 B.n784 VSUBS 0.012103f
C1019 B.n785 VSUBS 0.012103f
C1020 B.n786 VSUBS 0.012103f
C1021 B.n787 VSUBS 0.012103f
C1022 B.n788 VSUBS 0.012103f
C1023 B.n789 VSUBS 0.012103f
C1024 B.n790 VSUBS 0.012103f
C1025 B.n791 VSUBS 0.012103f
C1026 B.n792 VSUBS 0.012103f
C1027 B.n793 VSUBS 0.012103f
C1028 B.n794 VSUBS 0.012103f
C1029 B.n795 VSUBS 0.012103f
C1030 B.n796 VSUBS 0.012103f
C1031 B.n797 VSUBS 0.012103f
C1032 B.n798 VSUBS 0.012103f
C1033 B.n799 VSUBS 0.012103f
C1034 B.n800 VSUBS 0.012103f
C1035 B.n801 VSUBS 0.012103f
C1036 B.n802 VSUBS 0.012103f
C1037 B.n803 VSUBS 0.012103f
C1038 B.n804 VSUBS 0.012103f
C1039 B.n805 VSUBS 0.012103f
C1040 B.n806 VSUBS 0.012103f
C1041 B.n807 VSUBS 0.012103f
C1042 B.n808 VSUBS 0.012103f
C1043 B.n809 VSUBS 0.012103f
C1044 B.n810 VSUBS 0.012103f
C1045 B.n811 VSUBS 0.012103f
C1046 B.n812 VSUBS 0.012103f
C1047 B.n813 VSUBS 0.012103f
C1048 B.n814 VSUBS 0.012103f
C1049 B.n815 VSUBS 0.012103f
C1050 B.n816 VSUBS 0.012103f
C1051 B.n817 VSUBS 0.012103f
C1052 B.n818 VSUBS 0.012103f
C1053 B.n819 VSUBS 0.012103f
C1054 B.n820 VSUBS 0.012103f
C1055 B.n821 VSUBS 0.012103f
C1056 B.n822 VSUBS 0.012103f
C1057 B.n823 VSUBS 0.012103f
C1058 B.n824 VSUBS 0.012103f
C1059 B.n825 VSUBS 0.012103f
C1060 B.n826 VSUBS 0.012103f
C1061 B.n827 VSUBS 0.012103f
C1062 B.n828 VSUBS 0.012103f
C1063 B.n829 VSUBS 0.012103f
C1064 B.n830 VSUBS 0.012103f
C1065 B.n831 VSUBS 0.012103f
C1066 B.n832 VSUBS 0.012103f
C1067 B.n833 VSUBS 0.012103f
C1068 B.n834 VSUBS 0.012103f
C1069 B.n835 VSUBS 0.012103f
C1070 B.n836 VSUBS 0.012103f
C1071 B.n837 VSUBS 0.012103f
C1072 B.n838 VSUBS 0.012103f
C1073 B.n839 VSUBS 0.012103f
C1074 B.n840 VSUBS 0.012103f
C1075 B.n841 VSUBS 0.012103f
C1076 B.n842 VSUBS 0.012103f
C1077 B.n843 VSUBS 0.012103f
C1078 B.n844 VSUBS 0.012103f
C1079 B.n845 VSUBS 0.012103f
C1080 B.n846 VSUBS 0.012103f
C1081 B.n847 VSUBS 0.012103f
C1082 B.n848 VSUBS 0.012103f
C1083 B.n849 VSUBS 0.012103f
C1084 B.n850 VSUBS 0.012103f
C1085 B.n851 VSUBS 0.012103f
C1086 B.n852 VSUBS 0.012103f
C1087 B.n853 VSUBS 0.012103f
C1088 B.n854 VSUBS 0.012103f
C1089 B.n855 VSUBS 0.012103f
C1090 B.n856 VSUBS 0.012103f
C1091 B.n857 VSUBS 0.012103f
C1092 B.n858 VSUBS 0.012103f
C1093 B.n859 VSUBS 0.012103f
C1094 B.n860 VSUBS 0.012103f
C1095 B.n861 VSUBS 0.012103f
C1096 B.n862 VSUBS 0.012103f
C1097 B.n863 VSUBS 0.012103f
C1098 B.n864 VSUBS 0.012103f
C1099 B.n865 VSUBS 0.012103f
C1100 B.n866 VSUBS 0.012103f
C1101 B.n867 VSUBS 0.012103f
C1102 B.n868 VSUBS 0.012103f
C1103 B.n869 VSUBS 0.012103f
C1104 B.n870 VSUBS 0.012103f
C1105 B.n871 VSUBS 0.012103f
C1106 B.n872 VSUBS 0.012103f
C1107 B.n873 VSUBS 0.012103f
C1108 B.n874 VSUBS 0.012103f
C1109 B.n875 VSUBS 0.027405f
C1110 VTAIL.t0 VSUBS 0.150931f
C1111 VTAIL.t9 VSUBS 0.150931f
C1112 VTAIL.n0 VSUBS 0.846996f
C1113 VTAIL.n1 VSUBS 1.21348f
C1114 VTAIL.n2 VSUBS 0.038903f
C1115 VTAIL.n3 VSUBS 0.036242f
C1116 VTAIL.n4 VSUBS 0.019475f
C1117 VTAIL.n5 VSUBS 0.046032f
C1118 VTAIL.n6 VSUBS 0.020621f
C1119 VTAIL.n7 VSUBS 0.036242f
C1120 VTAIL.n8 VSUBS 0.019475f
C1121 VTAIL.n9 VSUBS 0.034524f
C1122 VTAIL.n10 VSUBS 0.029239f
C1123 VTAIL.t14 VSUBS 0.099224f
C1124 VTAIL.n11 VSUBS 0.152856f
C1125 VTAIL.n12 VSUBS 0.710357f
C1126 VTAIL.n13 VSUBS 0.019475f
C1127 VTAIL.n14 VSUBS 0.020621f
C1128 VTAIL.n15 VSUBS 0.046032f
C1129 VTAIL.n16 VSUBS 0.046032f
C1130 VTAIL.n17 VSUBS 0.020621f
C1131 VTAIL.n18 VSUBS 0.019475f
C1132 VTAIL.n19 VSUBS 0.036242f
C1133 VTAIL.n20 VSUBS 0.036242f
C1134 VTAIL.n21 VSUBS 0.019475f
C1135 VTAIL.n22 VSUBS 0.020621f
C1136 VTAIL.n23 VSUBS 0.046032f
C1137 VTAIL.n24 VSUBS 0.108305f
C1138 VTAIL.n25 VSUBS 0.020621f
C1139 VTAIL.n26 VSUBS 0.019475f
C1140 VTAIL.n27 VSUBS 0.083277f
C1141 VTAIL.n28 VSUBS 0.054311f
C1142 VTAIL.n29 VSUBS 0.709207f
C1143 VTAIL.t16 VSUBS 0.150931f
C1144 VTAIL.t13 VSUBS 0.150931f
C1145 VTAIL.n30 VSUBS 0.846996f
C1146 VTAIL.n31 VSUBS 1.46365f
C1147 VTAIL.t18 VSUBS 0.150931f
C1148 VTAIL.t17 VSUBS 0.150931f
C1149 VTAIL.n32 VSUBS 0.846996f
C1150 VTAIL.n33 VSUBS 2.90228f
C1151 VTAIL.t1 VSUBS 0.150931f
C1152 VTAIL.t6 VSUBS 0.150931f
C1153 VTAIL.n34 VSUBS 0.847003f
C1154 VTAIL.n35 VSUBS 2.90227f
C1155 VTAIL.t3 VSUBS 0.150931f
C1156 VTAIL.t2 VSUBS 0.150931f
C1157 VTAIL.n36 VSUBS 0.847003f
C1158 VTAIL.n37 VSUBS 1.46364f
C1159 VTAIL.n38 VSUBS 0.038903f
C1160 VTAIL.n39 VSUBS 0.036242f
C1161 VTAIL.n40 VSUBS 0.019475f
C1162 VTAIL.n41 VSUBS 0.046032f
C1163 VTAIL.n42 VSUBS 0.020621f
C1164 VTAIL.n43 VSUBS 0.036242f
C1165 VTAIL.n44 VSUBS 0.019475f
C1166 VTAIL.n45 VSUBS 0.034524f
C1167 VTAIL.n46 VSUBS 0.029239f
C1168 VTAIL.t4 VSUBS 0.099224f
C1169 VTAIL.n47 VSUBS 0.152856f
C1170 VTAIL.n48 VSUBS 0.710357f
C1171 VTAIL.n49 VSUBS 0.019475f
C1172 VTAIL.n50 VSUBS 0.020621f
C1173 VTAIL.n51 VSUBS 0.046032f
C1174 VTAIL.n52 VSUBS 0.046032f
C1175 VTAIL.n53 VSUBS 0.020621f
C1176 VTAIL.n54 VSUBS 0.019475f
C1177 VTAIL.n55 VSUBS 0.036242f
C1178 VTAIL.n56 VSUBS 0.036242f
C1179 VTAIL.n57 VSUBS 0.019475f
C1180 VTAIL.n58 VSUBS 0.020621f
C1181 VTAIL.n59 VSUBS 0.046032f
C1182 VTAIL.n60 VSUBS 0.108305f
C1183 VTAIL.n61 VSUBS 0.020621f
C1184 VTAIL.n62 VSUBS 0.019475f
C1185 VTAIL.n63 VSUBS 0.083277f
C1186 VTAIL.n64 VSUBS 0.054311f
C1187 VTAIL.n65 VSUBS 0.709207f
C1188 VTAIL.t10 VSUBS 0.150931f
C1189 VTAIL.t19 VSUBS 0.150931f
C1190 VTAIL.n66 VSUBS 0.847003f
C1191 VTAIL.n67 VSUBS 1.31062f
C1192 VTAIL.t12 VSUBS 0.150931f
C1193 VTAIL.t15 VSUBS 0.150931f
C1194 VTAIL.n68 VSUBS 0.847003f
C1195 VTAIL.n69 VSUBS 1.46364f
C1196 VTAIL.n70 VSUBS 0.038903f
C1197 VTAIL.n71 VSUBS 0.036242f
C1198 VTAIL.n72 VSUBS 0.019475f
C1199 VTAIL.n73 VSUBS 0.046032f
C1200 VTAIL.n74 VSUBS 0.020621f
C1201 VTAIL.n75 VSUBS 0.036242f
C1202 VTAIL.n76 VSUBS 0.019475f
C1203 VTAIL.n77 VSUBS 0.034524f
C1204 VTAIL.n78 VSUBS 0.029239f
C1205 VTAIL.t11 VSUBS 0.099224f
C1206 VTAIL.n79 VSUBS 0.152856f
C1207 VTAIL.n80 VSUBS 0.710357f
C1208 VTAIL.n81 VSUBS 0.019475f
C1209 VTAIL.n82 VSUBS 0.020621f
C1210 VTAIL.n83 VSUBS 0.046032f
C1211 VTAIL.n84 VSUBS 0.046032f
C1212 VTAIL.n85 VSUBS 0.020621f
C1213 VTAIL.n86 VSUBS 0.019475f
C1214 VTAIL.n87 VSUBS 0.036242f
C1215 VTAIL.n88 VSUBS 0.036242f
C1216 VTAIL.n89 VSUBS 0.019475f
C1217 VTAIL.n90 VSUBS 0.020621f
C1218 VTAIL.n91 VSUBS 0.046032f
C1219 VTAIL.n92 VSUBS 0.108305f
C1220 VTAIL.n93 VSUBS 0.020621f
C1221 VTAIL.n94 VSUBS 0.019475f
C1222 VTAIL.n95 VSUBS 0.083277f
C1223 VTAIL.n96 VSUBS 0.054311f
C1224 VTAIL.n97 VSUBS 1.88508f
C1225 VTAIL.n98 VSUBS 0.038903f
C1226 VTAIL.n99 VSUBS 0.036242f
C1227 VTAIL.n100 VSUBS 0.019475f
C1228 VTAIL.n101 VSUBS 0.046032f
C1229 VTAIL.n102 VSUBS 0.020621f
C1230 VTAIL.n103 VSUBS 0.036242f
C1231 VTAIL.n104 VSUBS 0.019475f
C1232 VTAIL.n105 VSUBS 0.034524f
C1233 VTAIL.n106 VSUBS 0.029239f
C1234 VTAIL.t7 VSUBS 0.099224f
C1235 VTAIL.n107 VSUBS 0.152856f
C1236 VTAIL.n108 VSUBS 0.710357f
C1237 VTAIL.n109 VSUBS 0.019475f
C1238 VTAIL.n110 VSUBS 0.020621f
C1239 VTAIL.n111 VSUBS 0.046032f
C1240 VTAIL.n112 VSUBS 0.046032f
C1241 VTAIL.n113 VSUBS 0.020621f
C1242 VTAIL.n114 VSUBS 0.019475f
C1243 VTAIL.n115 VSUBS 0.036242f
C1244 VTAIL.n116 VSUBS 0.036242f
C1245 VTAIL.n117 VSUBS 0.019475f
C1246 VTAIL.n118 VSUBS 0.020621f
C1247 VTAIL.n119 VSUBS 0.046032f
C1248 VTAIL.n120 VSUBS 0.108305f
C1249 VTAIL.n121 VSUBS 0.020621f
C1250 VTAIL.n122 VSUBS 0.019475f
C1251 VTAIL.n123 VSUBS 0.083277f
C1252 VTAIL.n124 VSUBS 0.054311f
C1253 VTAIL.n125 VSUBS 1.88508f
C1254 VTAIL.t8 VSUBS 0.150931f
C1255 VTAIL.t5 VSUBS 0.150931f
C1256 VTAIL.n126 VSUBS 0.846996f
C1257 VTAIL.n127 VSUBS 1.14502f
C1258 VDD1.n0 VSUBS 0.039296f
C1259 VDD1.n1 VSUBS 0.036608f
C1260 VDD1.n2 VSUBS 0.019672f
C1261 VDD1.n3 VSUBS 0.046497f
C1262 VDD1.n4 VSUBS 0.020829f
C1263 VDD1.n5 VSUBS 0.036608f
C1264 VDD1.n6 VSUBS 0.019672f
C1265 VDD1.n7 VSUBS 0.034873f
C1266 VDD1.n8 VSUBS 0.029535f
C1267 VDD1.t9 VSUBS 0.100227f
C1268 VDD1.n9 VSUBS 0.154401f
C1269 VDD1.n10 VSUBS 0.717535f
C1270 VDD1.n11 VSUBS 0.019672f
C1271 VDD1.n12 VSUBS 0.020829f
C1272 VDD1.n13 VSUBS 0.046497f
C1273 VDD1.n14 VSUBS 0.046497f
C1274 VDD1.n15 VSUBS 0.020829f
C1275 VDD1.n16 VSUBS 0.019672f
C1276 VDD1.n17 VSUBS 0.036608f
C1277 VDD1.n18 VSUBS 0.036608f
C1278 VDD1.n19 VSUBS 0.019672f
C1279 VDD1.n20 VSUBS 0.020829f
C1280 VDD1.n21 VSUBS 0.046497f
C1281 VDD1.n22 VSUBS 0.109399f
C1282 VDD1.n23 VSUBS 0.020829f
C1283 VDD1.n24 VSUBS 0.019672f
C1284 VDD1.n25 VSUBS 0.084118f
C1285 VDD1.n26 VSUBS 0.113556f
C1286 VDD1.t7 VSUBS 0.152456f
C1287 VDD1.t6 VSUBS 0.152456f
C1288 VDD1.n27 VSUBS 0.972538f
C1289 VDD1.n28 VSUBS 1.55986f
C1290 VDD1.n29 VSUBS 0.039296f
C1291 VDD1.n30 VSUBS 0.036608f
C1292 VDD1.n31 VSUBS 0.019672f
C1293 VDD1.n32 VSUBS 0.046497f
C1294 VDD1.n33 VSUBS 0.020829f
C1295 VDD1.n34 VSUBS 0.036608f
C1296 VDD1.n35 VSUBS 0.019672f
C1297 VDD1.n36 VSUBS 0.034873f
C1298 VDD1.n37 VSUBS 0.029535f
C1299 VDD1.t4 VSUBS 0.100227f
C1300 VDD1.n38 VSUBS 0.154401f
C1301 VDD1.n39 VSUBS 0.717535f
C1302 VDD1.n40 VSUBS 0.019672f
C1303 VDD1.n41 VSUBS 0.020829f
C1304 VDD1.n42 VSUBS 0.046497f
C1305 VDD1.n43 VSUBS 0.046497f
C1306 VDD1.n44 VSUBS 0.020829f
C1307 VDD1.n45 VSUBS 0.019672f
C1308 VDD1.n46 VSUBS 0.036608f
C1309 VDD1.n47 VSUBS 0.036608f
C1310 VDD1.n48 VSUBS 0.019672f
C1311 VDD1.n49 VSUBS 0.020829f
C1312 VDD1.n50 VSUBS 0.046497f
C1313 VDD1.n51 VSUBS 0.109399f
C1314 VDD1.n52 VSUBS 0.020829f
C1315 VDD1.n53 VSUBS 0.019672f
C1316 VDD1.n54 VSUBS 0.084118f
C1317 VDD1.n55 VSUBS 0.113556f
C1318 VDD1.t8 VSUBS 0.152456f
C1319 VDD1.t3 VSUBS 0.152456f
C1320 VDD1.n56 VSUBS 0.972533f
C1321 VDD1.n57 VSUBS 1.54749f
C1322 VDD1.t1 VSUBS 0.152456f
C1323 VDD1.t2 VSUBS 0.152456f
C1324 VDD1.n58 VSUBS 1.007f
C1325 VDD1.n59 VSUBS 5.06148f
C1326 VDD1.t5 VSUBS 0.152456f
C1327 VDD1.t0 VSUBS 0.152456f
C1328 VDD1.n60 VSUBS 0.972533f
C1329 VDD1.n61 VSUBS 4.89186f
C1330 VP.t5 VSUBS 1.91115f
C1331 VP.n0 VSUBS 0.845467f
C1332 VP.n1 VSUBS 0.036353f
C1333 VP.n2 VSUBS 0.073446f
C1334 VP.n3 VSUBS 0.036353f
C1335 VP.n4 VSUBS 0.067752f
C1336 VP.n5 VSUBS 0.036353f
C1337 VP.t6 VSUBS 1.91115f
C1338 VP.n6 VSUBS 0.067752f
C1339 VP.n7 VSUBS 0.036353f
C1340 VP.n8 VSUBS 0.067752f
C1341 VP.n9 VSUBS 0.036353f
C1342 VP.t3 VSUBS 1.91115f
C1343 VP.n10 VSUBS 0.067752f
C1344 VP.n11 VSUBS 0.036353f
C1345 VP.n12 VSUBS 0.067752f
C1346 VP.n13 VSUBS 0.036353f
C1347 VP.t2 VSUBS 1.91115f
C1348 VP.n14 VSUBS 0.067752f
C1349 VP.n15 VSUBS 0.036353f
C1350 VP.n16 VSUBS 0.067752f
C1351 VP.n17 VSUBS 0.058672f
C1352 VP.t1 VSUBS 1.91115f
C1353 VP.t8 VSUBS 1.91115f
C1354 VP.n18 VSUBS 0.845467f
C1355 VP.n19 VSUBS 0.036353f
C1356 VP.n20 VSUBS 0.073446f
C1357 VP.n21 VSUBS 0.036353f
C1358 VP.n22 VSUBS 0.067752f
C1359 VP.n23 VSUBS 0.036353f
C1360 VP.t4 VSUBS 1.91115f
C1361 VP.n24 VSUBS 0.067752f
C1362 VP.n25 VSUBS 0.036353f
C1363 VP.n26 VSUBS 0.067752f
C1364 VP.n27 VSUBS 0.036353f
C1365 VP.t7 VSUBS 1.91115f
C1366 VP.n28 VSUBS 0.067752f
C1367 VP.n29 VSUBS 0.036353f
C1368 VP.n30 VSUBS 0.067752f
C1369 VP.t9 VSUBS 2.40321f
C1370 VP.n31 VSUBS 0.838577f
C1371 VP.t0 VSUBS 1.91115f
C1372 VP.n32 VSUBS 0.853332f
C1373 VP.n33 VSUBS 0.059724f
C1374 VP.n34 VSUBS 0.469019f
C1375 VP.n35 VSUBS 0.036353f
C1376 VP.n36 VSUBS 0.036353f
C1377 VP.n37 VSUBS 0.067752f
C1378 VP.n38 VSUBS 0.046487f
C1379 VP.n39 VSUBS 0.059656f
C1380 VP.n40 VSUBS 0.036353f
C1381 VP.n41 VSUBS 0.036353f
C1382 VP.n42 VSUBS 0.036353f
C1383 VP.n43 VSUBS 0.067752f
C1384 VP.n44 VSUBS 0.051027f
C1385 VP.n45 VSUBS 0.713514f
C1386 VP.n46 VSUBS 0.051027f
C1387 VP.n47 VSUBS 0.036353f
C1388 VP.n48 VSUBS 0.036353f
C1389 VP.n49 VSUBS 0.036353f
C1390 VP.n50 VSUBS 0.067752f
C1391 VP.n51 VSUBS 0.059656f
C1392 VP.n52 VSUBS 0.046487f
C1393 VP.n53 VSUBS 0.036353f
C1394 VP.n54 VSUBS 0.036353f
C1395 VP.n55 VSUBS 0.036353f
C1396 VP.n56 VSUBS 0.067752f
C1397 VP.n57 VSUBS 0.059724f
C1398 VP.n58 VSUBS 0.713514f
C1399 VP.n59 VSUBS 0.04233f
C1400 VP.n60 VSUBS 0.036353f
C1401 VP.n61 VSUBS 0.036353f
C1402 VP.n62 VSUBS 0.036353f
C1403 VP.n63 VSUBS 0.067752f
C1404 VP.n64 VSUBS 0.069623f
C1405 VP.n65 VSUBS 0.030826f
C1406 VP.n66 VSUBS 0.036353f
C1407 VP.n67 VSUBS 0.036353f
C1408 VP.n68 VSUBS 0.036353f
C1409 VP.n69 VSUBS 0.067752f
C1410 VP.n70 VSUBS 0.067752f
C1411 VP.n71 VSUBS 0.034972f
C1412 VP.n72 VSUBS 0.058672f
C1413 VP.n73 VSUBS 2.364f
C1414 VP.n74 VSUBS 2.38796f
C1415 VP.n75 VSUBS 0.845467f
C1416 VP.n76 VSUBS 0.034972f
C1417 VP.n77 VSUBS 0.067752f
C1418 VP.n78 VSUBS 0.036353f
C1419 VP.n79 VSUBS 0.036353f
C1420 VP.n80 VSUBS 0.036353f
C1421 VP.n81 VSUBS 0.073446f
C1422 VP.n82 VSUBS 0.030826f
C1423 VP.n83 VSUBS 0.069623f
C1424 VP.n84 VSUBS 0.036353f
C1425 VP.n85 VSUBS 0.036353f
C1426 VP.n86 VSUBS 0.036353f
C1427 VP.n87 VSUBS 0.067752f
C1428 VP.n88 VSUBS 0.04233f
C1429 VP.n89 VSUBS 0.713514f
C1430 VP.n90 VSUBS 0.059724f
C1431 VP.n91 VSUBS 0.036353f
C1432 VP.n92 VSUBS 0.036353f
C1433 VP.n93 VSUBS 0.036353f
C1434 VP.n94 VSUBS 0.067752f
C1435 VP.n95 VSUBS 0.046487f
C1436 VP.n96 VSUBS 0.059656f
C1437 VP.n97 VSUBS 0.036353f
C1438 VP.n98 VSUBS 0.036353f
C1439 VP.n99 VSUBS 0.036353f
C1440 VP.n100 VSUBS 0.067752f
C1441 VP.n101 VSUBS 0.051027f
C1442 VP.n102 VSUBS 0.713514f
C1443 VP.n103 VSUBS 0.051027f
C1444 VP.n104 VSUBS 0.036353f
C1445 VP.n105 VSUBS 0.036353f
C1446 VP.n106 VSUBS 0.036353f
C1447 VP.n107 VSUBS 0.067752f
C1448 VP.n108 VSUBS 0.059656f
C1449 VP.n109 VSUBS 0.046487f
C1450 VP.n110 VSUBS 0.036353f
C1451 VP.n111 VSUBS 0.036353f
C1452 VP.n112 VSUBS 0.036353f
C1453 VP.n113 VSUBS 0.067752f
C1454 VP.n114 VSUBS 0.059724f
C1455 VP.n115 VSUBS 0.713514f
C1456 VP.n116 VSUBS 0.04233f
C1457 VP.n117 VSUBS 0.036353f
C1458 VP.n118 VSUBS 0.036353f
C1459 VP.n119 VSUBS 0.036353f
C1460 VP.n120 VSUBS 0.067752f
C1461 VP.n121 VSUBS 0.069623f
C1462 VP.n122 VSUBS 0.030826f
C1463 VP.n123 VSUBS 0.036353f
C1464 VP.n124 VSUBS 0.036353f
C1465 VP.n125 VSUBS 0.036353f
C1466 VP.n126 VSUBS 0.067752f
C1467 VP.n127 VSUBS 0.067752f
C1468 VP.n128 VSUBS 0.034972f
C1469 VP.n129 VSUBS 0.058672f
C1470 VP.n130 VSUBS 0.11413f
.ends

