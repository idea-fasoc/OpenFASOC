* NGSPICE file created from diff_pair_sample_1516.ext - technology: sky130A

.subckt diff_pair_sample_1516 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=0.4953 pd=3.32 as=0 ps=0 w=1.27 l=3.82
X1 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=0.4953 pd=3.32 as=0 ps=0 w=1.27 l=3.82
X2 VDD1.t1 VP.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.4953 pd=3.32 as=0.4953 ps=3.32 w=1.27 l=3.82
X3 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.4953 pd=3.32 as=0 ps=0 w=1.27 l=3.82
X4 VDD2.t1 VN.t0 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.4953 pd=3.32 as=0.4953 ps=3.32 w=1.27 l=3.82
X5 VDD2.t0 VN.t1 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4953 pd=3.32 as=0.4953 ps=3.32 w=1.27 l=3.82
X6 VDD1.t0 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4953 pd=3.32 as=0.4953 ps=3.32 w=1.27 l=3.82
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.4953 pd=3.32 as=0 ps=0 w=1.27 l=3.82
R0 B.n421 B.n420 585
R1 B.n138 B.n77 585
R2 B.n137 B.n136 585
R3 B.n135 B.n134 585
R4 B.n133 B.n132 585
R5 B.n131 B.n130 585
R6 B.n129 B.n128 585
R7 B.n127 B.n126 585
R8 B.n125 B.n124 585
R9 B.n123 B.n122 585
R10 B.n121 B.n120 585
R11 B.n119 B.n118 585
R12 B.n117 B.n116 585
R13 B.n115 B.n114 585
R14 B.n113 B.n112 585
R15 B.n111 B.n110 585
R16 B.n109 B.n108 585
R17 B.n107 B.n106 585
R18 B.n105 B.n104 585
R19 B.n103 B.n102 585
R20 B.n101 B.n100 585
R21 B.n99 B.n98 585
R22 B.n97 B.n96 585
R23 B.n95 B.n94 585
R24 B.n93 B.n92 585
R25 B.n91 B.n90 585
R26 B.n89 B.n88 585
R27 B.n87 B.n86 585
R28 B.n85 B.n84 585
R29 B.n61 B.n60 585
R30 B.n419 B.n62 585
R31 B.n424 B.n62 585
R32 B.n418 B.n417 585
R33 B.n417 B.n58 585
R34 B.n416 B.n57 585
R35 B.n430 B.n57 585
R36 B.n415 B.n56 585
R37 B.n431 B.n56 585
R38 B.n414 B.n55 585
R39 B.n432 B.n55 585
R40 B.n413 B.n412 585
R41 B.n412 B.n51 585
R42 B.n411 B.n50 585
R43 B.n438 B.n50 585
R44 B.n410 B.n49 585
R45 B.n439 B.n49 585
R46 B.n409 B.n48 585
R47 B.n440 B.n48 585
R48 B.n408 B.n407 585
R49 B.n407 B.n47 585
R50 B.n406 B.n43 585
R51 B.n446 B.n43 585
R52 B.n405 B.n42 585
R53 B.n447 B.n42 585
R54 B.n404 B.n41 585
R55 B.n448 B.n41 585
R56 B.n403 B.n402 585
R57 B.n402 B.n37 585
R58 B.n401 B.n36 585
R59 B.n454 B.n36 585
R60 B.n400 B.n35 585
R61 B.n455 B.n35 585
R62 B.n399 B.n34 585
R63 B.n456 B.n34 585
R64 B.n398 B.n397 585
R65 B.n397 B.n30 585
R66 B.n396 B.n29 585
R67 B.n462 B.n29 585
R68 B.n395 B.n28 585
R69 B.n463 B.n28 585
R70 B.n394 B.n27 585
R71 B.n464 B.n27 585
R72 B.n393 B.n392 585
R73 B.n392 B.n23 585
R74 B.n391 B.n22 585
R75 B.n470 B.n22 585
R76 B.n390 B.n21 585
R77 B.n471 B.n21 585
R78 B.n389 B.n20 585
R79 B.n472 B.n20 585
R80 B.n388 B.n387 585
R81 B.n387 B.n16 585
R82 B.n386 B.n15 585
R83 B.n478 B.n15 585
R84 B.n385 B.n14 585
R85 B.n479 B.n14 585
R86 B.n384 B.n13 585
R87 B.n480 B.n13 585
R88 B.n383 B.n382 585
R89 B.n382 B.n12 585
R90 B.n381 B.n380 585
R91 B.n381 B.n8 585
R92 B.n379 B.n7 585
R93 B.n487 B.n7 585
R94 B.n378 B.n6 585
R95 B.n488 B.n6 585
R96 B.n377 B.n5 585
R97 B.n489 B.n5 585
R98 B.n376 B.n375 585
R99 B.n375 B.n4 585
R100 B.n374 B.n139 585
R101 B.n374 B.n373 585
R102 B.n364 B.n140 585
R103 B.n141 B.n140 585
R104 B.n366 B.n365 585
R105 B.n367 B.n366 585
R106 B.n363 B.n146 585
R107 B.n146 B.n145 585
R108 B.n362 B.n361 585
R109 B.n361 B.n360 585
R110 B.n148 B.n147 585
R111 B.n149 B.n148 585
R112 B.n353 B.n352 585
R113 B.n354 B.n353 585
R114 B.n351 B.n154 585
R115 B.n154 B.n153 585
R116 B.n350 B.n349 585
R117 B.n349 B.n348 585
R118 B.n156 B.n155 585
R119 B.n157 B.n156 585
R120 B.n341 B.n340 585
R121 B.n342 B.n341 585
R122 B.n339 B.n162 585
R123 B.n162 B.n161 585
R124 B.n338 B.n337 585
R125 B.n337 B.n336 585
R126 B.n164 B.n163 585
R127 B.n165 B.n164 585
R128 B.n329 B.n328 585
R129 B.n330 B.n329 585
R130 B.n327 B.n170 585
R131 B.n170 B.n169 585
R132 B.n326 B.n325 585
R133 B.n325 B.n324 585
R134 B.n172 B.n171 585
R135 B.n173 B.n172 585
R136 B.n317 B.n316 585
R137 B.n318 B.n317 585
R138 B.n315 B.n178 585
R139 B.n178 B.n177 585
R140 B.n314 B.n313 585
R141 B.n313 B.n312 585
R142 B.n180 B.n179 585
R143 B.n305 B.n180 585
R144 B.n304 B.n303 585
R145 B.n306 B.n304 585
R146 B.n302 B.n185 585
R147 B.n185 B.n184 585
R148 B.n301 B.n300 585
R149 B.n300 B.n299 585
R150 B.n187 B.n186 585
R151 B.n188 B.n187 585
R152 B.n292 B.n291 585
R153 B.n293 B.n292 585
R154 B.n290 B.n193 585
R155 B.n193 B.n192 585
R156 B.n289 B.n288 585
R157 B.n288 B.n287 585
R158 B.n195 B.n194 585
R159 B.n196 B.n195 585
R160 B.n280 B.n279 585
R161 B.n281 B.n280 585
R162 B.n199 B.n198 585
R163 B.n220 B.n218 585
R164 B.n221 B.n217 585
R165 B.n221 B.n200 585
R166 B.n224 B.n223 585
R167 B.n225 B.n216 585
R168 B.n227 B.n226 585
R169 B.n229 B.n215 585
R170 B.n232 B.n231 585
R171 B.n233 B.n214 585
R172 B.n238 B.n237 585
R173 B.n240 B.n213 585
R174 B.n243 B.n242 585
R175 B.n244 B.n212 585
R176 B.n246 B.n245 585
R177 B.n248 B.n211 585
R178 B.n251 B.n250 585
R179 B.n252 B.n210 585
R180 B.n254 B.n253 585
R181 B.n256 B.n209 585
R182 B.n259 B.n258 585
R183 B.n261 B.n206 585
R184 B.n263 B.n262 585
R185 B.n265 B.n205 585
R186 B.n268 B.n267 585
R187 B.n269 B.n204 585
R188 B.n271 B.n270 585
R189 B.n273 B.n203 585
R190 B.n274 B.n202 585
R191 B.n277 B.n276 585
R192 B.n278 B.n201 585
R193 B.n201 B.n200 585
R194 B.n283 B.n282 585
R195 B.n282 B.n281 585
R196 B.n284 B.n197 585
R197 B.n197 B.n196 585
R198 B.n286 B.n285 585
R199 B.n287 B.n286 585
R200 B.n191 B.n190 585
R201 B.n192 B.n191 585
R202 B.n295 B.n294 585
R203 B.n294 B.n293 585
R204 B.n296 B.n189 585
R205 B.n189 B.n188 585
R206 B.n298 B.n297 585
R207 B.n299 B.n298 585
R208 B.n183 B.n182 585
R209 B.n184 B.n183 585
R210 B.n308 B.n307 585
R211 B.n307 B.n306 585
R212 B.n309 B.n181 585
R213 B.n305 B.n181 585
R214 B.n311 B.n310 585
R215 B.n312 B.n311 585
R216 B.n176 B.n175 585
R217 B.n177 B.n176 585
R218 B.n320 B.n319 585
R219 B.n319 B.n318 585
R220 B.n321 B.n174 585
R221 B.n174 B.n173 585
R222 B.n323 B.n322 585
R223 B.n324 B.n323 585
R224 B.n168 B.n167 585
R225 B.n169 B.n168 585
R226 B.n332 B.n331 585
R227 B.n331 B.n330 585
R228 B.n333 B.n166 585
R229 B.n166 B.n165 585
R230 B.n335 B.n334 585
R231 B.n336 B.n335 585
R232 B.n160 B.n159 585
R233 B.n161 B.n160 585
R234 B.n344 B.n343 585
R235 B.n343 B.n342 585
R236 B.n345 B.n158 585
R237 B.n158 B.n157 585
R238 B.n347 B.n346 585
R239 B.n348 B.n347 585
R240 B.n152 B.n151 585
R241 B.n153 B.n152 585
R242 B.n356 B.n355 585
R243 B.n355 B.n354 585
R244 B.n357 B.n150 585
R245 B.n150 B.n149 585
R246 B.n359 B.n358 585
R247 B.n360 B.n359 585
R248 B.n144 B.n143 585
R249 B.n145 B.n144 585
R250 B.n369 B.n368 585
R251 B.n368 B.n367 585
R252 B.n370 B.n142 585
R253 B.n142 B.n141 585
R254 B.n372 B.n371 585
R255 B.n373 B.n372 585
R256 B.n3 B.n0 585
R257 B.n4 B.n3 585
R258 B.n486 B.n1 585
R259 B.n487 B.n486 585
R260 B.n485 B.n484 585
R261 B.n485 B.n8 585
R262 B.n483 B.n9 585
R263 B.n12 B.n9 585
R264 B.n482 B.n481 585
R265 B.n481 B.n480 585
R266 B.n11 B.n10 585
R267 B.n479 B.n11 585
R268 B.n477 B.n476 585
R269 B.n478 B.n477 585
R270 B.n475 B.n17 585
R271 B.n17 B.n16 585
R272 B.n474 B.n473 585
R273 B.n473 B.n472 585
R274 B.n19 B.n18 585
R275 B.n471 B.n19 585
R276 B.n469 B.n468 585
R277 B.n470 B.n469 585
R278 B.n467 B.n24 585
R279 B.n24 B.n23 585
R280 B.n466 B.n465 585
R281 B.n465 B.n464 585
R282 B.n26 B.n25 585
R283 B.n463 B.n26 585
R284 B.n461 B.n460 585
R285 B.n462 B.n461 585
R286 B.n459 B.n31 585
R287 B.n31 B.n30 585
R288 B.n458 B.n457 585
R289 B.n457 B.n456 585
R290 B.n33 B.n32 585
R291 B.n455 B.n33 585
R292 B.n453 B.n452 585
R293 B.n454 B.n453 585
R294 B.n451 B.n38 585
R295 B.n38 B.n37 585
R296 B.n450 B.n449 585
R297 B.n449 B.n448 585
R298 B.n40 B.n39 585
R299 B.n447 B.n40 585
R300 B.n445 B.n444 585
R301 B.n446 B.n445 585
R302 B.n443 B.n44 585
R303 B.n47 B.n44 585
R304 B.n442 B.n441 585
R305 B.n441 B.n440 585
R306 B.n46 B.n45 585
R307 B.n439 B.n46 585
R308 B.n437 B.n436 585
R309 B.n438 B.n437 585
R310 B.n435 B.n52 585
R311 B.n52 B.n51 585
R312 B.n434 B.n433 585
R313 B.n433 B.n432 585
R314 B.n54 B.n53 585
R315 B.n431 B.n54 585
R316 B.n429 B.n428 585
R317 B.n430 B.n429 585
R318 B.n427 B.n59 585
R319 B.n59 B.n58 585
R320 B.n426 B.n425 585
R321 B.n425 B.n424 585
R322 B.n490 B.n489 585
R323 B.n488 B.n2 585
R324 B.n425 B.n61 478.086
R325 B.n421 B.n62 478.086
R326 B.n280 B.n201 478.086
R327 B.n282 B.n199 478.086
R328 B.n423 B.n422 256.663
R329 B.n423 B.n76 256.663
R330 B.n423 B.n75 256.663
R331 B.n423 B.n74 256.663
R332 B.n423 B.n73 256.663
R333 B.n423 B.n72 256.663
R334 B.n423 B.n71 256.663
R335 B.n423 B.n70 256.663
R336 B.n423 B.n69 256.663
R337 B.n423 B.n68 256.663
R338 B.n423 B.n67 256.663
R339 B.n423 B.n66 256.663
R340 B.n423 B.n65 256.663
R341 B.n423 B.n64 256.663
R342 B.n423 B.n63 256.663
R343 B.n219 B.n200 256.663
R344 B.n222 B.n200 256.663
R345 B.n228 B.n200 256.663
R346 B.n230 B.n200 256.663
R347 B.n239 B.n200 256.663
R348 B.n241 B.n200 256.663
R349 B.n247 B.n200 256.663
R350 B.n249 B.n200 256.663
R351 B.n255 B.n200 256.663
R352 B.n257 B.n200 256.663
R353 B.n264 B.n200 256.663
R354 B.n266 B.n200 256.663
R355 B.n272 B.n200 256.663
R356 B.n275 B.n200 256.663
R357 B.n492 B.n491 256.663
R358 B.n81 B.t11 230.082
R359 B.n78 B.t8 230.082
R360 B.n207 B.t5 230.082
R361 B.n234 B.t15 230.082
R362 B.n281 B.n200 210.084
R363 B.n424 B.n423 210.084
R364 B.n81 B.t10 209.885
R365 B.n78 B.t6 209.885
R366 B.n207 B.t2 209.885
R367 B.n234 B.t13 209.885
R368 B.n86 B.n85 163.367
R369 B.n90 B.n89 163.367
R370 B.n94 B.n93 163.367
R371 B.n98 B.n97 163.367
R372 B.n102 B.n101 163.367
R373 B.n106 B.n105 163.367
R374 B.n110 B.n109 163.367
R375 B.n114 B.n113 163.367
R376 B.n118 B.n117 163.367
R377 B.n122 B.n121 163.367
R378 B.n126 B.n125 163.367
R379 B.n130 B.n129 163.367
R380 B.n134 B.n133 163.367
R381 B.n136 B.n77 163.367
R382 B.n280 B.n195 163.367
R383 B.n288 B.n195 163.367
R384 B.n288 B.n193 163.367
R385 B.n292 B.n193 163.367
R386 B.n292 B.n187 163.367
R387 B.n300 B.n187 163.367
R388 B.n300 B.n185 163.367
R389 B.n304 B.n185 163.367
R390 B.n304 B.n180 163.367
R391 B.n313 B.n180 163.367
R392 B.n313 B.n178 163.367
R393 B.n317 B.n178 163.367
R394 B.n317 B.n172 163.367
R395 B.n325 B.n172 163.367
R396 B.n325 B.n170 163.367
R397 B.n329 B.n170 163.367
R398 B.n329 B.n164 163.367
R399 B.n337 B.n164 163.367
R400 B.n337 B.n162 163.367
R401 B.n341 B.n162 163.367
R402 B.n341 B.n156 163.367
R403 B.n349 B.n156 163.367
R404 B.n349 B.n154 163.367
R405 B.n353 B.n154 163.367
R406 B.n353 B.n148 163.367
R407 B.n361 B.n148 163.367
R408 B.n361 B.n146 163.367
R409 B.n366 B.n146 163.367
R410 B.n366 B.n140 163.367
R411 B.n374 B.n140 163.367
R412 B.n375 B.n374 163.367
R413 B.n375 B.n5 163.367
R414 B.n6 B.n5 163.367
R415 B.n7 B.n6 163.367
R416 B.n381 B.n7 163.367
R417 B.n382 B.n381 163.367
R418 B.n382 B.n13 163.367
R419 B.n14 B.n13 163.367
R420 B.n15 B.n14 163.367
R421 B.n387 B.n15 163.367
R422 B.n387 B.n20 163.367
R423 B.n21 B.n20 163.367
R424 B.n22 B.n21 163.367
R425 B.n392 B.n22 163.367
R426 B.n392 B.n27 163.367
R427 B.n28 B.n27 163.367
R428 B.n29 B.n28 163.367
R429 B.n397 B.n29 163.367
R430 B.n397 B.n34 163.367
R431 B.n35 B.n34 163.367
R432 B.n36 B.n35 163.367
R433 B.n402 B.n36 163.367
R434 B.n402 B.n41 163.367
R435 B.n42 B.n41 163.367
R436 B.n43 B.n42 163.367
R437 B.n407 B.n43 163.367
R438 B.n407 B.n48 163.367
R439 B.n49 B.n48 163.367
R440 B.n50 B.n49 163.367
R441 B.n412 B.n50 163.367
R442 B.n412 B.n55 163.367
R443 B.n56 B.n55 163.367
R444 B.n57 B.n56 163.367
R445 B.n417 B.n57 163.367
R446 B.n417 B.n62 163.367
R447 B.n221 B.n220 163.367
R448 B.n223 B.n221 163.367
R449 B.n227 B.n216 163.367
R450 B.n231 B.n229 163.367
R451 B.n238 B.n214 163.367
R452 B.n242 B.n240 163.367
R453 B.n246 B.n212 163.367
R454 B.n250 B.n248 163.367
R455 B.n254 B.n210 163.367
R456 B.n258 B.n256 163.367
R457 B.n263 B.n206 163.367
R458 B.n267 B.n265 163.367
R459 B.n271 B.n204 163.367
R460 B.n274 B.n273 163.367
R461 B.n276 B.n201 163.367
R462 B.n282 B.n197 163.367
R463 B.n286 B.n197 163.367
R464 B.n286 B.n191 163.367
R465 B.n294 B.n191 163.367
R466 B.n294 B.n189 163.367
R467 B.n298 B.n189 163.367
R468 B.n298 B.n183 163.367
R469 B.n307 B.n183 163.367
R470 B.n307 B.n181 163.367
R471 B.n311 B.n181 163.367
R472 B.n311 B.n176 163.367
R473 B.n319 B.n176 163.367
R474 B.n319 B.n174 163.367
R475 B.n323 B.n174 163.367
R476 B.n323 B.n168 163.367
R477 B.n331 B.n168 163.367
R478 B.n331 B.n166 163.367
R479 B.n335 B.n166 163.367
R480 B.n335 B.n160 163.367
R481 B.n343 B.n160 163.367
R482 B.n343 B.n158 163.367
R483 B.n347 B.n158 163.367
R484 B.n347 B.n152 163.367
R485 B.n355 B.n152 163.367
R486 B.n355 B.n150 163.367
R487 B.n359 B.n150 163.367
R488 B.n359 B.n144 163.367
R489 B.n368 B.n144 163.367
R490 B.n368 B.n142 163.367
R491 B.n372 B.n142 163.367
R492 B.n372 B.n3 163.367
R493 B.n490 B.n3 163.367
R494 B.n486 B.n2 163.367
R495 B.n486 B.n485 163.367
R496 B.n485 B.n9 163.367
R497 B.n481 B.n9 163.367
R498 B.n481 B.n11 163.367
R499 B.n477 B.n11 163.367
R500 B.n477 B.n17 163.367
R501 B.n473 B.n17 163.367
R502 B.n473 B.n19 163.367
R503 B.n469 B.n19 163.367
R504 B.n469 B.n24 163.367
R505 B.n465 B.n24 163.367
R506 B.n465 B.n26 163.367
R507 B.n461 B.n26 163.367
R508 B.n461 B.n31 163.367
R509 B.n457 B.n31 163.367
R510 B.n457 B.n33 163.367
R511 B.n453 B.n33 163.367
R512 B.n453 B.n38 163.367
R513 B.n449 B.n38 163.367
R514 B.n449 B.n40 163.367
R515 B.n445 B.n40 163.367
R516 B.n445 B.n44 163.367
R517 B.n441 B.n44 163.367
R518 B.n441 B.n46 163.367
R519 B.n437 B.n46 163.367
R520 B.n437 B.n52 163.367
R521 B.n433 B.n52 163.367
R522 B.n433 B.n54 163.367
R523 B.n429 B.n54 163.367
R524 B.n429 B.n59 163.367
R525 B.n425 B.n59 163.367
R526 B.n82 B.t12 149.596
R527 B.n79 B.t9 149.596
R528 B.n208 B.t4 149.596
R529 B.n235 B.t14 149.596
R530 B.n281 B.n196 114.287
R531 B.n287 B.n196 114.287
R532 B.n287 B.n192 114.287
R533 B.n293 B.n192 114.287
R534 B.n293 B.n188 114.287
R535 B.n299 B.n188 114.287
R536 B.n299 B.n184 114.287
R537 B.n306 B.n184 114.287
R538 B.n306 B.n305 114.287
R539 B.n312 B.n177 114.287
R540 B.n318 B.n177 114.287
R541 B.n318 B.n173 114.287
R542 B.n324 B.n173 114.287
R543 B.n324 B.n169 114.287
R544 B.n330 B.n169 114.287
R545 B.n330 B.n165 114.287
R546 B.n336 B.n165 114.287
R547 B.n336 B.n161 114.287
R548 B.n342 B.n161 114.287
R549 B.n342 B.n157 114.287
R550 B.n348 B.n157 114.287
R551 B.n348 B.n153 114.287
R552 B.n354 B.n153 114.287
R553 B.n360 B.n149 114.287
R554 B.n360 B.n145 114.287
R555 B.n367 B.n145 114.287
R556 B.n367 B.n141 114.287
R557 B.n373 B.n141 114.287
R558 B.n373 B.n4 114.287
R559 B.n489 B.n4 114.287
R560 B.n489 B.n488 114.287
R561 B.n488 B.n487 114.287
R562 B.n487 B.n8 114.287
R563 B.n12 B.n8 114.287
R564 B.n480 B.n12 114.287
R565 B.n480 B.n479 114.287
R566 B.n479 B.n478 114.287
R567 B.n478 B.n16 114.287
R568 B.n472 B.n471 114.287
R569 B.n471 B.n470 114.287
R570 B.n470 B.n23 114.287
R571 B.n464 B.n23 114.287
R572 B.n464 B.n463 114.287
R573 B.n463 B.n462 114.287
R574 B.n462 B.n30 114.287
R575 B.n456 B.n30 114.287
R576 B.n456 B.n455 114.287
R577 B.n455 B.n454 114.287
R578 B.n454 B.n37 114.287
R579 B.n448 B.n37 114.287
R580 B.n448 B.n447 114.287
R581 B.n447 B.n446 114.287
R582 B.n440 B.n47 114.287
R583 B.n440 B.n439 114.287
R584 B.n439 B.n438 114.287
R585 B.n438 B.n51 114.287
R586 B.n432 B.n51 114.287
R587 B.n432 B.n431 114.287
R588 B.n431 B.n430 114.287
R589 B.n430 B.n58 114.287
R590 B.n424 B.n58 114.287
R591 B.n354 B.t0 90.7568
R592 B.n472 B.t1 90.7568
R593 B.n82 B.n81 80.4853
R594 B.n79 B.n78 80.4853
R595 B.n208 B.n207 80.4853
R596 B.n235 B.n234 80.4853
R597 B.n63 B.n61 71.676
R598 B.n86 B.n64 71.676
R599 B.n90 B.n65 71.676
R600 B.n94 B.n66 71.676
R601 B.n98 B.n67 71.676
R602 B.n102 B.n68 71.676
R603 B.n106 B.n69 71.676
R604 B.n110 B.n70 71.676
R605 B.n114 B.n71 71.676
R606 B.n118 B.n72 71.676
R607 B.n122 B.n73 71.676
R608 B.n126 B.n74 71.676
R609 B.n130 B.n75 71.676
R610 B.n134 B.n76 71.676
R611 B.n422 B.n77 71.676
R612 B.n422 B.n421 71.676
R613 B.n136 B.n76 71.676
R614 B.n133 B.n75 71.676
R615 B.n129 B.n74 71.676
R616 B.n125 B.n73 71.676
R617 B.n121 B.n72 71.676
R618 B.n117 B.n71 71.676
R619 B.n113 B.n70 71.676
R620 B.n109 B.n69 71.676
R621 B.n105 B.n68 71.676
R622 B.n101 B.n67 71.676
R623 B.n97 B.n66 71.676
R624 B.n93 B.n65 71.676
R625 B.n89 B.n64 71.676
R626 B.n85 B.n63 71.676
R627 B.n219 B.n199 71.676
R628 B.n223 B.n222 71.676
R629 B.n228 B.n227 71.676
R630 B.n231 B.n230 71.676
R631 B.n239 B.n238 71.676
R632 B.n242 B.n241 71.676
R633 B.n247 B.n246 71.676
R634 B.n250 B.n249 71.676
R635 B.n255 B.n254 71.676
R636 B.n258 B.n257 71.676
R637 B.n264 B.n263 71.676
R638 B.n267 B.n266 71.676
R639 B.n272 B.n271 71.676
R640 B.n275 B.n274 71.676
R641 B.n220 B.n219 71.676
R642 B.n222 B.n216 71.676
R643 B.n229 B.n228 71.676
R644 B.n230 B.n214 71.676
R645 B.n240 B.n239 71.676
R646 B.n241 B.n212 71.676
R647 B.n248 B.n247 71.676
R648 B.n249 B.n210 71.676
R649 B.n256 B.n255 71.676
R650 B.n257 B.n206 71.676
R651 B.n265 B.n264 71.676
R652 B.n266 B.n204 71.676
R653 B.n273 B.n272 71.676
R654 B.n276 B.n275 71.676
R655 B.n491 B.n490 71.676
R656 B.n491 B.n2 71.676
R657 B.n312 B.t3 70.5887
R658 B.n446 B.t7 70.5887
R659 B.n83 B.n82 59.5399
R660 B.n80 B.n79 59.5399
R661 B.n260 B.n208 59.5399
R662 B.n236 B.n235 59.5399
R663 B.n305 B.t3 43.698
R664 B.n47 B.t7 43.698
R665 B.n283 B.n198 31.0639
R666 B.n279 B.n278 31.0639
R667 B.n420 B.n419 31.0639
R668 B.n426 B.n60 31.0639
R669 B.t0 B.n149 23.5299
R670 B.t1 B.n16 23.5299
R671 B B.n492 18.0485
R672 B.n284 B.n283 10.6151
R673 B.n285 B.n284 10.6151
R674 B.n285 B.n190 10.6151
R675 B.n295 B.n190 10.6151
R676 B.n296 B.n295 10.6151
R677 B.n297 B.n296 10.6151
R678 B.n297 B.n182 10.6151
R679 B.n308 B.n182 10.6151
R680 B.n309 B.n308 10.6151
R681 B.n310 B.n309 10.6151
R682 B.n310 B.n175 10.6151
R683 B.n320 B.n175 10.6151
R684 B.n321 B.n320 10.6151
R685 B.n322 B.n321 10.6151
R686 B.n322 B.n167 10.6151
R687 B.n332 B.n167 10.6151
R688 B.n333 B.n332 10.6151
R689 B.n334 B.n333 10.6151
R690 B.n334 B.n159 10.6151
R691 B.n344 B.n159 10.6151
R692 B.n345 B.n344 10.6151
R693 B.n346 B.n345 10.6151
R694 B.n346 B.n151 10.6151
R695 B.n356 B.n151 10.6151
R696 B.n357 B.n356 10.6151
R697 B.n358 B.n357 10.6151
R698 B.n358 B.n143 10.6151
R699 B.n369 B.n143 10.6151
R700 B.n370 B.n369 10.6151
R701 B.n371 B.n370 10.6151
R702 B.n371 B.n0 10.6151
R703 B.n218 B.n198 10.6151
R704 B.n218 B.n217 10.6151
R705 B.n224 B.n217 10.6151
R706 B.n225 B.n224 10.6151
R707 B.n226 B.n225 10.6151
R708 B.n226 B.n215 10.6151
R709 B.n232 B.n215 10.6151
R710 B.n233 B.n232 10.6151
R711 B.n237 B.n233 10.6151
R712 B.n243 B.n213 10.6151
R713 B.n244 B.n243 10.6151
R714 B.n245 B.n244 10.6151
R715 B.n245 B.n211 10.6151
R716 B.n251 B.n211 10.6151
R717 B.n252 B.n251 10.6151
R718 B.n253 B.n252 10.6151
R719 B.n253 B.n209 10.6151
R720 B.n259 B.n209 10.6151
R721 B.n262 B.n261 10.6151
R722 B.n262 B.n205 10.6151
R723 B.n268 B.n205 10.6151
R724 B.n269 B.n268 10.6151
R725 B.n270 B.n269 10.6151
R726 B.n270 B.n203 10.6151
R727 B.n203 B.n202 10.6151
R728 B.n277 B.n202 10.6151
R729 B.n278 B.n277 10.6151
R730 B.n279 B.n194 10.6151
R731 B.n289 B.n194 10.6151
R732 B.n290 B.n289 10.6151
R733 B.n291 B.n290 10.6151
R734 B.n291 B.n186 10.6151
R735 B.n301 B.n186 10.6151
R736 B.n302 B.n301 10.6151
R737 B.n303 B.n302 10.6151
R738 B.n303 B.n179 10.6151
R739 B.n314 B.n179 10.6151
R740 B.n315 B.n314 10.6151
R741 B.n316 B.n315 10.6151
R742 B.n316 B.n171 10.6151
R743 B.n326 B.n171 10.6151
R744 B.n327 B.n326 10.6151
R745 B.n328 B.n327 10.6151
R746 B.n328 B.n163 10.6151
R747 B.n338 B.n163 10.6151
R748 B.n339 B.n338 10.6151
R749 B.n340 B.n339 10.6151
R750 B.n340 B.n155 10.6151
R751 B.n350 B.n155 10.6151
R752 B.n351 B.n350 10.6151
R753 B.n352 B.n351 10.6151
R754 B.n352 B.n147 10.6151
R755 B.n362 B.n147 10.6151
R756 B.n363 B.n362 10.6151
R757 B.n365 B.n363 10.6151
R758 B.n365 B.n364 10.6151
R759 B.n364 B.n139 10.6151
R760 B.n376 B.n139 10.6151
R761 B.n377 B.n376 10.6151
R762 B.n378 B.n377 10.6151
R763 B.n379 B.n378 10.6151
R764 B.n380 B.n379 10.6151
R765 B.n383 B.n380 10.6151
R766 B.n384 B.n383 10.6151
R767 B.n385 B.n384 10.6151
R768 B.n386 B.n385 10.6151
R769 B.n388 B.n386 10.6151
R770 B.n389 B.n388 10.6151
R771 B.n390 B.n389 10.6151
R772 B.n391 B.n390 10.6151
R773 B.n393 B.n391 10.6151
R774 B.n394 B.n393 10.6151
R775 B.n395 B.n394 10.6151
R776 B.n396 B.n395 10.6151
R777 B.n398 B.n396 10.6151
R778 B.n399 B.n398 10.6151
R779 B.n400 B.n399 10.6151
R780 B.n401 B.n400 10.6151
R781 B.n403 B.n401 10.6151
R782 B.n404 B.n403 10.6151
R783 B.n405 B.n404 10.6151
R784 B.n406 B.n405 10.6151
R785 B.n408 B.n406 10.6151
R786 B.n409 B.n408 10.6151
R787 B.n410 B.n409 10.6151
R788 B.n411 B.n410 10.6151
R789 B.n413 B.n411 10.6151
R790 B.n414 B.n413 10.6151
R791 B.n415 B.n414 10.6151
R792 B.n416 B.n415 10.6151
R793 B.n418 B.n416 10.6151
R794 B.n419 B.n418 10.6151
R795 B.n484 B.n1 10.6151
R796 B.n484 B.n483 10.6151
R797 B.n483 B.n482 10.6151
R798 B.n482 B.n10 10.6151
R799 B.n476 B.n10 10.6151
R800 B.n476 B.n475 10.6151
R801 B.n475 B.n474 10.6151
R802 B.n474 B.n18 10.6151
R803 B.n468 B.n18 10.6151
R804 B.n468 B.n467 10.6151
R805 B.n467 B.n466 10.6151
R806 B.n466 B.n25 10.6151
R807 B.n460 B.n25 10.6151
R808 B.n460 B.n459 10.6151
R809 B.n459 B.n458 10.6151
R810 B.n458 B.n32 10.6151
R811 B.n452 B.n32 10.6151
R812 B.n452 B.n451 10.6151
R813 B.n451 B.n450 10.6151
R814 B.n450 B.n39 10.6151
R815 B.n444 B.n39 10.6151
R816 B.n444 B.n443 10.6151
R817 B.n443 B.n442 10.6151
R818 B.n442 B.n45 10.6151
R819 B.n436 B.n45 10.6151
R820 B.n436 B.n435 10.6151
R821 B.n435 B.n434 10.6151
R822 B.n434 B.n53 10.6151
R823 B.n428 B.n53 10.6151
R824 B.n428 B.n427 10.6151
R825 B.n427 B.n426 10.6151
R826 B.n84 B.n60 10.6151
R827 B.n87 B.n84 10.6151
R828 B.n88 B.n87 10.6151
R829 B.n91 B.n88 10.6151
R830 B.n92 B.n91 10.6151
R831 B.n95 B.n92 10.6151
R832 B.n96 B.n95 10.6151
R833 B.n99 B.n96 10.6151
R834 B.n100 B.n99 10.6151
R835 B.n104 B.n103 10.6151
R836 B.n107 B.n104 10.6151
R837 B.n108 B.n107 10.6151
R838 B.n111 B.n108 10.6151
R839 B.n112 B.n111 10.6151
R840 B.n115 B.n112 10.6151
R841 B.n116 B.n115 10.6151
R842 B.n119 B.n116 10.6151
R843 B.n120 B.n119 10.6151
R844 B.n124 B.n123 10.6151
R845 B.n127 B.n124 10.6151
R846 B.n128 B.n127 10.6151
R847 B.n131 B.n128 10.6151
R848 B.n132 B.n131 10.6151
R849 B.n135 B.n132 10.6151
R850 B.n137 B.n135 10.6151
R851 B.n138 B.n137 10.6151
R852 B.n420 B.n138 10.6151
R853 B.n237 B.n236 9.36635
R854 B.n261 B.n260 9.36635
R855 B.n100 B.n83 9.36635
R856 B.n123 B.n80 9.36635
R857 B.n492 B.n0 8.11757
R858 B.n492 B.n1 8.11757
R859 B.n236 B.n213 1.24928
R860 B.n260 B.n259 1.24928
R861 B.n103 B.n83 1.24928
R862 B.n120 B.n80 1.24928
R863 VP.n0 VP.t1 82.8129
R864 VP.n0 VP.t0 43.0499
R865 VP VP.n0 0.621237
R866 VTAIL.n3 VTAIL.t0 155.714
R867 VTAIL.n0 VTAIL.t2 155.714
R868 VTAIL.n2 VTAIL.t3 155.714
R869 VTAIL.n1 VTAIL.t1 155.714
R870 VTAIL.n1 VTAIL.n0 20.6169
R871 VTAIL.n3 VTAIL.n2 17.0393
R872 VTAIL.n2 VTAIL.n1 2.25912
R873 VTAIL VTAIL.n0 1.42291
R874 VTAIL VTAIL.n3 0.836707
R875 VDD1 VDD1.t1 205.721
R876 VDD1 VDD1.t0 173.345
R877 VN VN.t0 82.6252
R878 VN VN.t1 43.6707
R879 VDD2.n0 VDD2.t0 204.303
R880 VDD2.n0 VDD2.t1 172.393
R881 VDD2 VDD2.n0 0.953086
C0 VP VDD1 0.780346f
C1 VP VN 4.05149f
C2 VDD1 VTAIL 2.64533f
C3 VTAIL VN 1.08947f
C4 VDD2 VP 0.392173f
C5 VDD2 VTAIL 2.70676f
C6 VDD1 VN 0.156049f
C7 VP VTAIL 1.10365f
C8 VDD2 VDD1 0.809674f
C9 VDD2 VN 0.546166f
C10 VDD2 B 2.923385f
C11 VDD1 B 5.187941f
C12 VTAIL B 2.988663f
C13 VN B 9.167769f
C14 VP B 6.923026f
C15 VDD2.t0 B 0.277167f
C16 VDD2.t1 B 0.130791f
C17 VDD2.n0 B 2.1185f
C18 VN.t1 B 0.606881f
C19 VN.t0 B 1.28106f
C20 VDD1.t0 B 0.123834f
C21 VDD1.t1 B 0.275844f
C22 VTAIL.t2 B 0.139947f
C23 VTAIL.n0 B 1.25879f
C24 VTAIL.t1 B 0.139947f
C25 VTAIL.n1 B 1.32353f
C26 VTAIL.t3 B 0.139947f
C27 VTAIL.n2 B 1.04658f
C28 VTAIL.t0 B 0.139947f
C29 VTAIL.n3 B 0.93647f
C30 VP.t1 B 1.29438f
C31 VP.t0 B 0.608465f
C32 VP.n0 B 2.07398f
.ends

