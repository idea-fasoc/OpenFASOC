* NGSPICE file created from diff_pair_sample_1179.ext - technology: sky130A

.subckt diff_pair_sample_1179 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=4.9764 pd=26.3 as=0 ps=0 w=12.76 l=3.89
X1 VTAIL.t11 VN.t0 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1054 pd=13.09 as=2.1054 ps=13.09 w=12.76 l=3.89
X2 VDD1.t5 VP.t0 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=4.9764 pd=26.3 as=2.1054 ps=13.09 w=12.76 l=3.89
X3 VDD2.t3 VN.t1 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=4.9764 pd=26.3 as=2.1054 ps=13.09 w=12.76 l=3.89
X4 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=4.9764 pd=26.3 as=0 ps=0 w=12.76 l=3.89
X5 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.9764 pd=26.3 as=0 ps=0 w=12.76 l=3.89
X6 VDD1.t4 VP.t1 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.1054 pd=13.09 as=4.9764 ps=26.3 w=12.76 l=3.89
X7 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.9764 pd=26.3 as=0 ps=0 w=12.76 l=3.89
X8 VTAIL.t5 VP.t2 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1054 pd=13.09 as=2.1054 ps=13.09 w=12.76 l=3.89
X9 VDD2.t4 VN.t2 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=4.9764 pd=26.3 as=2.1054 ps=13.09 w=12.76 l=3.89
X10 VDD2.t2 VN.t3 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1054 pd=13.09 as=4.9764 ps=26.3 w=12.76 l=3.89
X11 VTAIL.t1 VP.t3 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.1054 pd=13.09 as=2.1054 ps=13.09 w=12.76 l=3.89
X12 VDD1.t1 VP.t4 VTAIL.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=4.9764 pd=26.3 as=2.1054 ps=13.09 w=12.76 l=3.89
X13 VDD2.t5 VN.t4 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.1054 pd=13.09 as=4.9764 ps=26.3 w=12.76 l=3.89
X14 VDD1.t0 VP.t5 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1054 pd=13.09 as=4.9764 ps=26.3 w=12.76 l=3.89
X15 VTAIL.t6 VN.t5 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.1054 pd=13.09 as=2.1054 ps=13.09 w=12.76 l=3.89
R0 B.n958 B.n957 585
R1 B.n959 B.n958 585
R2 B.n351 B.n154 585
R3 B.n350 B.n349 585
R4 B.n348 B.n347 585
R5 B.n346 B.n345 585
R6 B.n344 B.n343 585
R7 B.n342 B.n341 585
R8 B.n340 B.n339 585
R9 B.n338 B.n337 585
R10 B.n336 B.n335 585
R11 B.n334 B.n333 585
R12 B.n332 B.n331 585
R13 B.n330 B.n329 585
R14 B.n328 B.n327 585
R15 B.n326 B.n325 585
R16 B.n324 B.n323 585
R17 B.n322 B.n321 585
R18 B.n320 B.n319 585
R19 B.n318 B.n317 585
R20 B.n316 B.n315 585
R21 B.n314 B.n313 585
R22 B.n312 B.n311 585
R23 B.n310 B.n309 585
R24 B.n308 B.n307 585
R25 B.n306 B.n305 585
R26 B.n304 B.n303 585
R27 B.n302 B.n301 585
R28 B.n300 B.n299 585
R29 B.n298 B.n297 585
R30 B.n296 B.n295 585
R31 B.n294 B.n293 585
R32 B.n292 B.n291 585
R33 B.n290 B.n289 585
R34 B.n288 B.n287 585
R35 B.n286 B.n285 585
R36 B.n284 B.n283 585
R37 B.n282 B.n281 585
R38 B.n280 B.n279 585
R39 B.n278 B.n277 585
R40 B.n276 B.n275 585
R41 B.n274 B.n273 585
R42 B.n272 B.n271 585
R43 B.n270 B.n269 585
R44 B.n268 B.n267 585
R45 B.n265 B.n264 585
R46 B.n263 B.n262 585
R47 B.n261 B.n260 585
R48 B.n259 B.n258 585
R49 B.n257 B.n256 585
R50 B.n255 B.n254 585
R51 B.n253 B.n252 585
R52 B.n251 B.n250 585
R53 B.n249 B.n248 585
R54 B.n247 B.n246 585
R55 B.n245 B.n244 585
R56 B.n243 B.n242 585
R57 B.n241 B.n240 585
R58 B.n239 B.n238 585
R59 B.n237 B.n236 585
R60 B.n235 B.n234 585
R61 B.n233 B.n232 585
R62 B.n231 B.n230 585
R63 B.n229 B.n228 585
R64 B.n227 B.n226 585
R65 B.n225 B.n224 585
R66 B.n223 B.n222 585
R67 B.n221 B.n220 585
R68 B.n219 B.n218 585
R69 B.n217 B.n216 585
R70 B.n215 B.n214 585
R71 B.n213 B.n212 585
R72 B.n211 B.n210 585
R73 B.n209 B.n208 585
R74 B.n207 B.n206 585
R75 B.n205 B.n204 585
R76 B.n203 B.n202 585
R77 B.n201 B.n200 585
R78 B.n199 B.n198 585
R79 B.n197 B.n196 585
R80 B.n195 B.n194 585
R81 B.n193 B.n192 585
R82 B.n191 B.n190 585
R83 B.n189 B.n188 585
R84 B.n187 B.n186 585
R85 B.n185 B.n184 585
R86 B.n183 B.n182 585
R87 B.n181 B.n180 585
R88 B.n179 B.n178 585
R89 B.n177 B.n176 585
R90 B.n175 B.n174 585
R91 B.n173 B.n172 585
R92 B.n171 B.n170 585
R93 B.n169 B.n168 585
R94 B.n167 B.n166 585
R95 B.n165 B.n164 585
R96 B.n163 B.n162 585
R97 B.n161 B.n160 585
R98 B.n956 B.n105 585
R99 B.n960 B.n105 585
R100 B.n955 B.n104 585
R101 B.n961 B.n104 585
R102 B.n954 B.n953 585
R103 B.n953 B.n100 585
R104 B.n952 B.n99 585
R105 B.n967 B.n99 585
R106 B.n951 B.n98 585
R107 B.n968 B.n98 585
R108 B.n950 B.n97 585
R109 B.n969 B.n97 585
R110 B.n949 B.n948 585
R111 B.n948 B.n93 585
R112 B.n947 B.n92 585
R113 B.n975 B.n92 585
R114 B.n946 B.n91 585
R115 B.n976 B.n91 585
R116 B.n945 B.n90 585
R117 B.n977 B.n90 585
R118 B.n944 B.n943 585
R119 B.n943 B.n86 585
R120 B.n942 B.n85 585
R121 B.n983 B.n85 585
R122 B.n941 B.n84 585
R123 B.n984 B.n84 585
R124 B.n940 B.n83 585
R125 B.n985 B.n83 585
R126 B.n939 B.n938 585
R127 B.n938 B.n79 585
R128 B.n937 B.n78 585
R129 B.n991 B.n78 585
R130 B.n936 B.n77 585
R131 B.n992 B.n77 585
R132 B.n935 B.n76 585
R133 B.n993 B.n76 585
R134 B.n934 B.n933 585
R135 B.n933 B.n72 585
R136 B.n932 B.n71 585
R137 B.n999 B.n71 585
R138 B.n931 B.n70 585
R139 B.n1000 B.n70 585
R140 B.n930 B.n69 585
R141 B.n1001 B.n69 585
R142 B.n929 B.n928 585
R143 B.n928 B.n65 585
R144 B.n927 B.n64 585
R145 B.n1007 B.n64 585
R146 B.n926 B.n63 585
R147 B.n1008 B.n63 585
R148 B.n925 B.n62 585
R149 B.n1009 B.n62 585
R150 B.n924 B.n923 585
R151 B.n923 B.n58 585
R152 B.n922 B.n57 585
R153 B.n1015 B.n57 585
R154 B.n921 B.n56 585
R155 B.n1016 B.n56 585
R156 B.n920 B.n55 585
R157 B.n1017 B.n55 585
R158 B.n919 B.n918 585
R159 B.n918 B.n51 585
R160 B.n917 B.n50 585
R161 B.n1023 B.n50 585
R162 B.n916 B.n49 585
R163 B.n1024 B.n49 585
R164 B.n915 B.n48 585
R165 B.n1025 B.n48 585
R166 B.n914 B.n913 585
R167 B.n913 B.n44 585
R168 B.n912 B.n43 585
R169 B.n1031 B.n43 585
R170 B.n911 B.n42 585
R171 B.n1032 B.n42 585
R172 B.n910 B.n41 585
R173 B.n1033 B.n41 585
R174 B.n909 B.n908 585
R175 B.n908 B.n37 585
R176 B.n907 B.n36 585
R177 B.n1039 B.n36 585
R178 B.n906 B.n35 585
R179 B.n1040 B.n35 585
R180 B.n905 B.n34 585
R181 B.n1041 B.n34 585
R182 B.n904 B.n903 585
R183 B.n903 B.n30 585
R184 B.n902 B.n29 585
R185 B.n1047 B.n29 585
R186 B.n901 B.n28 585
R187 B.n1048 B.n28 585
R188 B.n900 B.n27 585
R189 B.n1049 B.n27 585
R190 B.n899 B.n898 585
R191 B.n898 B.n23 585
R192 B.n897 B.n22 585
R193 B.n1055 B.n22 585
R194 B.n896 B.n21 585
R195 B.n1056 B.n21 585
R196 B.n895 B.n20 585
R197 B.n1057 B.n20 585
R198 B.n894 B.n893 585
R199 B.n893 B.n16 585
R200 B.n892 B.n15 585
R201 B.n1063 B.n15 585
R202 B.n891 B.n14 585
R203 B.n1064 B.n14 585
R204 B.n890 B.n13 585
R205 B.n1065 B.n13 585
R206 B.n889 B.n888 585
R207 B.n888 B.n12 585
R208 B.n887 B.n886 585
R209 B.n887 B.n8 585
R210 B.n885 B.n7 585
R211 B.n1072 B.n7 585
R212 B.n884 B.n6 585
R213 B.n1073 B.n6 585
R214 B.n883 B.n5 585
R215 B.n1074 B.n5 585
R216 B.n882 B.n881 585
R217 B.n881 B.n4 585
R218 B.n880 B.n352 585
R219 B.n880 B.n879 585
R220 B.n870 B.n353 585
R221 B.n354 B.n353 585
R222 B.n872 B.n871 585
R223 B.n873 B.n872 585
R224 B.n869 B.n359 585
R225 B.n359 B.n358 585
R226 B.n868 B.n867 585
R227 B.n867 B.n866 585
R228 B.n361 B.n360 585
R229 B.n362 B.n361 585
R230 B.n859 B.n858 585
R231 B.n860 B.n859 585
R232 B.n857 B.n367 585
R233 B.n367 B.n366 585
R234 B.n856 B.n855 585
R235 B.n855 B.n854 585
R236 B.n369 B.n368 585
R237 B.n370 B.n369 585
R238 B.n847 B.n846 585
R239 B.n848 B.n847 585
R240 B.n845 B.n375 585
R241 B.n375 B.n374 585
R242 B.n844 B.n843 585
R243 B.n843 B.n842 585
R244 B.n377 B.n376 585
R245 B.n378 B.n377 585
R246 B.n835 B.n834 585
R247 B.n836 B.n835 585
R248 B.n833 B.n383 585
R249 B.n383 B.n382 585
R250 B.n832 B.n831 585
R251 B.n831 B.n830 585
R252 B.n385 B.n384 585
R253 B.n386 B.n385 585
R254 B.n823 B.n822 585
R255 B.n824 B.n823 585
R256 B.n821 B.n391 585
R257 B.n391 B.n390 585
R258 B.n820 B.n819 585
R259 B.n819 B.n818 585
R260 B.n393 B.n392 585
R261 B.n394 B.n393 585
R262 B.n811 B.n810 585
R263 B.n812 B.n811 585
R264 B.n809 B.n399 585
R265 B.n399 B.n398 585
R266 B.n808 B.n807 585
R267 B.n807 B.n806 585
R268 B.n401 B.n400 585
R269 B.n402 B.n401 585
R270 B.n799 B.n798 585
R271 B.n800 B.n799 585
R272 B.n797 B.n407 585
R273 B.n407 B.n406 585
R274 B.n796 B.n795 585
R275 B.n795 B.n794 585
R276 B.n409 B.n408 585
R277 B.n410 B.n409 585
R278 B.n787 B.n786 585
R279 B.n788 B.n787 585
R280 B.n785 B.n414 585
R281 B.n418 B.n414 585
R282 B.n784 B.n783 585
R283 B.n783 B.n782 585
R284 B.n416 B.n415 585
R285 B.n417 B.n416 585
R286 B.n775 B.n774 585
R287 B.n776 B.n775 585
R288 B.n773 B.n423 585
R289 B.n423 B.n422 585
R290 B.n772 B.n771 585
R291 B.n771 B.n770 585
R292 B.n425 B.n424 585
R293 B.n426 B.n425 585
R294 B.n763 B.n762 585
R295 B.n764 B.n763 585
R296 B.n761 B.n431 585
R297 B.n431 B.n430 585
R298 B.n760 B.n759 585
R299 B.n759 B.n758 585
R300 B.n433 B.n432 585
R301 B.n434 B.n433 585
R302 B.n751 B.n750 585
R303 B.n752 B.n751 585
R304 B.n749 B.n439 585
R305 B.n439 B.n438 585
R306 B.n748 B.n747 585
R307 B.n747 B.n746 585
R308 B.n441 B.n440 585
R309 B.n442 B.n441 585
R310 B.n739 B.n738 585
R311 B.n740 B.n739 585
R312 B.n737 B.n447 585
R313 B.n447 B.n446 585
R314 B.n736 B.n735 585
R315 B.n735 B.n734 585
R316 B.n449 B.n448 585
R317 B.n450 B.n449 585
R318 B.n727 B.n726 585
R319 B.n728 B.n727 585
R320 B.n725 B.n455 585
R321 B.n455 B.n454 585
R322 B.n724 B.n723 585
R323 B.n723 B.n722 585
R324 B.n457 B.n456 585
R325 B.n458 B.n457 585
R326 B.n715 B.n714 585
R327 B.n716 B.n715 585
R328 B.n713 B.n463 585
R329 B.n463 B.n462 585
R330 B.n707 B.n706 585
R331 B.n705 B.n513 585
R332 B.n704 B.n512 585
R333 B.n709 B.n512 585
R334 B.n703 B.n702 585
R335 B.n701 B.n700 585
R336 B.n699 B.n698 585
R337 B.n697 B.n696 585
R338 B.n695 B.n694 585
R339 B.n693 B.n692 585
R340 B.n691 B.n690 585
R341 B.n689 B.n688 585
R342 B.n687 B.n686 585
R343 B.n685 B.n684 585
R344 B.n683 B.n682 585
R345 B.n681 B.n680 585
R346 B.n679 B.n678 585
R347 B.n677 B.n676 585
R348 B.n675 B.n674 585
R349 B.n673 B.n672 585
R350 B.n671 B.n670 585
R351 B.n669 B.n668 585
R352 B.n667 B.n666 585
R353 B.n665 B.n664 585
R354 B.n663 B.n662 585
R355 B.n661 B.n660 585
R356 B.n659 B.n658 585
R357 B.n657 B.n656 585
R358 B.n655 B.n654 585
R359 B.n653 B.n652 585
R360 B.n651 B.n650 585
R361 B.n649 B.n648 585
R362 B.n647 B.n646 585
R363 B.n645 B.n644 585
R364 B.n643 B.n642 585
R365 B.n641 B.n640 585
R366 B.n639 B.n638 585
R367 B.n637 B.n636 585
R368 B.n635 B.n634 585
R369 B.n633 B.n632 585
R370 B.n631 B.n630 585
R371 B.n629 B.n628 585
R372 B.n627 B.n626 585
R373 B.n625 B.n624 585
R374 B.n623 B.n622 585
R375 B.n620 B.n619 585
R376 B.n618 B.n617 585
R377 B.n616 B.n615 585
R378 B.n614 B.n613 585
R379 B.n612 B.n611 585
R380 B.n610 B.n609 585
R381 B.n608 B.n607 585
R382 B.n606 B.n605 585
R383 B.n604 B.n603 585
R384 B.n602 B.n601 585
R385 B.n600 B.n599 585
R386 B.n598 B.n597 585
R387 B.n596 B.n595 585
R388 B.n594 B.n593 585
R389 B.n592 B.n591 585
R390 B.n590 B.n589 585
R391 B.n588 B.n587 585
R392 B.n586 B.n585 585
R393 B.n584 B.n583 585
R394 B.n582 B.n581 585
R395 B.n580 B.n579 585
R396 B.n578 B.n577 585
R397 B.n576 B.n575 585
R398 B.n574 B.n573 585
R399 B.n572 B.n571 585
R400 B.n570 B.n569 585
R401 B.n568 B.n567 585
R402 B.n566 B.n565 585
R403 B.n564 B.n563 585
R404 B.n562 B.n561 585
R405 B.n560 B.n559 585
R406 B.n558 B.n557 585
R407 B.n556 B.n555 585
R408 B.n554 B.n553 585
R409 B.n552 B.n551 585
R410 B.n550 B.n549 585
R411 B.n548 B.n547 585
R412 B.n546 B.n545 585
R413 B.n544 B.n543 585
R414 B.n542 B.n541 585
R415 B.n540 B.n539 585
R416 B.n538 B.n537 585
R417 B.n536 B.n535 585
R418 B.n534 B.n533 585
R419 B.n532 B.n531 585
R420 B.n530 B.n529 585
R421 B.n528 B.n527 585
R422 B.n526 B.n525 585
R423 B.n524 B.n523 585
R424 B.n522 B.n521 585
R425 B.n520 B.n519 585
R426 B.n465 B.n464 585
R427 B.n712 B.n711 585
R428 B.n461 B.n460 585
R429 B.n462 B.n461 585
R430 B.n718 B.n717 585
R431 B.n717 B.n716 585
R432 B.n719 B.n459 585
R433 B.n459 B.n458 585
R434 B.n721 B.n720 585
R435 B.n722 B.n721 585
R436 B.n453 B.n452 585
R437 B.n454 B.n453 585
R438 B.n730 B.n729 585
R439 B.n729 B.n728 585
R440 B.n731 B.n451 585
R441 B.n451 B.n450 585
R442 B.n733 B.n732 585
R443 B.n734 B.n733 585
R444 B.n445 B.n444 585
R445 B.n446 B.n445 585
R446 B.n742 B.n741 585
R447 B.n741 B.n740 585
R448 B.n743 B.n443 585
R449 B.n443 B.n442 585
R450 B.n745 B.n744 585
R451 B.n746 B.n745 585
R452 B.n437 B.n436 585
R453 B.n438 B.n437 585
R454 B.n754 B.n753 585
R455 B.n753 B.n752 585
R456 B.n755 B.n435 585
R457 B.n435 B.n434 585
R458 B.n757 B.n756 585
R459 B.n758 B.n757 585
R460 B.n429 B.n428 585
R461 B.n430 B.n429 585
R462 B.n766 B.n765 585
R463 B.n765 B.n764 585
R464 B.n767 B.n427 585
R465 B.n427 B.n426 585
R466 B.n769 B.n768 585
R467 B.n770 B.n769 585
R468 B.n421 B.n420 585
R469 B.n422 B.n421 585
R470 B.n778 B.n777 585
R471 B.n777 B.n776 585
R472 B.n779 B.n419 585
R473 B.n419 B.n417 585
R474 B.n781 B.n780 585
R475 B.n782 B.n781 585
R476 B.n413 B.n412 585
R477 B.n418 B.n413 585
R478 B.n790 B.n789 585
R479 B.n789 B.n788 585
R480 B.n791 B.n411 585
R481 B.n411 B.n410 585
R482 B.n793 B.n792 585
R483 B.n794 B.n793 585
R484 B.n405 B.n404 585
R485 B.n406 B.n405 585
R486 B.n802 B.n801 585
R487 B.n801 B.n800 585
R488 B.n803 B.n403 585
R489 B.n403 B.n402 585
R490 B.n805 B.n804 585
R491 B.n806 B.n805 585
R492 B.n397 B.n396 585
R493 B.n398 B.n397 585
R494 B.n814 B.n813 585
R495 B.n813 B.n812 585
R496 B.n815 B.n395 585
R497 B.n395 B.n394 585
R498 B.n817 B.n816 585
R499 B.n818 B.n817 585
R500 B.n389 B.n388 585
R501 B.n390 B.n389 585
R502 B.n826 B.n825 585
R503 B.n825 B.n824 585
R504 B.n827 B.n387 585
R505 B.n387 B.n386 585
R506 B.n829 B.n828 585
R507 B.n830 B.n829 585
R508 B.n381 B.n380 585
R509 B.n382 B.n381 585
R510 B.n838 B.n837 585
R511 B.n837 B.n836 585
R512 B.n839 B.n379 585
R513 B.n379 B.n378 585
R514 B.n841 B.n840 585
R515 B.n842 B.n841 585
R516 B.n373 B.n372 585
R517 B.n374 B.n373 585
R518 B.n850 B.n849 585
R519 B.n849 B.n848 585
R520 B.n851 B.n371 585
R521 B.n371 B.n370 585
R522 B.n853 B.n852 585
R523 B.n854 B.n853 585
R524 B.n365 B.n364 585
R525 B.n366 B.n365 585
R526 B.n862 B.n861 585
R527 B.n861 B.n860 585
R528 B.n863 B.n363 585
R529 B.n363 B.n362 585
R530 B.n865 B.n864 585
R531 B.n866 B.n865 585
R532 B.n357 B.n356 585
R533 B.n358 B.n357 585
R534 B.n875 B.n874 585
R535 B.n874 B.n873 585
R536 B.n876 B.n355 585
R537 B.n355 B.n354 585
R538 B.n878 B.n877 585
R539 B.n879 B.n878 585
R540 B.n3 B.n0 585
R541 B.n4 B.n3 585
R542 B.n1071 B.n1 585
R543 B.n1072 B.n1071 585
R544 B.n1070 B.n1069 585
R545 B.n1070 B.n8 585
R546 B.n1068 B.n9 585
R547 B.n12 B.n9 585
R548 B.n1067 B.n1066 585
R549 B.n1066 B.n1065 585
R550 B.n11 B.n10 585
R551 B.n1064 B.n11 585
R552 B.n1062 B.n1061 585
R553 B.n1063 B.n1062 585
R554 B.n1060 B.n17 585
R555 B.n17 B.n16 585
R556 B.n1059 B.n1058 585
R557 B.n1058 B.n1057 585
R558 B.n19 B.n18 585
R559 B.n1056 B.n19 585
R560 B.n1054 B.n1053 585
R561 B.n1055 B.n1054 585
R562 B.n1052 B.n24 585
R563 B.n24 B.n23 585
R564 B.n1051 B.n1050 585
R565 B.n1050 B.n1049 585
R566 B.n26 B.n25 585
R567 B.n1048 B.n26 585
R568 B.n1046 B.n1045 585
R569 B.n1047 B.n1046 585
R570 B.n1044 B.n31 585
R571 B.n31 B.n30 585
R572 B.n1043 B.n1042 585
R573 B.n1042 B.n1041 585
R574 B.n33 B.n32 585
R575 B.n1040 B.n33 585
R576 B.n1038 B.n1037 585
R577 B.n1039 B.n1038 585
R578 B.n1036 B.n38 585
R579 B.n38 B.n37 585
R580 B.n1035 B.n1034 585
R581 B.n1034 B.n1033 585
R582 B.n40 B.n39 585
R583 B.n1032 B.n40 585
R584 B.n1030 B.n1029 585
R585 B.n1031 B.n1030 585
R586 B.n1028 B.n45 585
R587 B.n45 B.n44 585
R588 B.n1027 B.n1026 585
R589 B.n1026 B.n1025 585
R590 B.n47 B.n46 585
R591 B.n1024 B.n47 585
R592 B.n1022 B.n1021 585
R593 B.n1023 B.n1022 585
R594 B.n1020 B.n52 585
R595 B.n52 B.n51 585
R596 B.n1019 B.n1018 585
R597 B.n1018 B.n1017 585
R598 B.n54 B.n53 585
R599 B.n1016 B.n54 585
R600 B.n1014 B.n1013 585
R601 B.n1015 B.n1014 585
R602 B.n1012 B.n59 585
R603 B.n59 B.n58 585
R604 B.n1011 B.n1010 585
R605 B.n1010 B.n1009 585
R606 B.n61 B.n60 585
R607 B.n1008 B.n61 585
R608 B.n1006 B.n1005 585
R609 B.n1007 B.n1006 585
R610 B.n1004 B.n66 585
R611 B.n66 B.n65 585
R612 B.n1003 B.n1002 585
R613 B.n1002 B.n1001 585
R614 B.n68 B.n67 585
R615 B.n1000 B.n68 585
R616 B.n998 B.n997 585
R617 B.n999 B.n998 585
R618 B.n996 B.n73 585
R619 B.n73 B.n72 585
R620 B.n995 B.n994 585
R621 B.n994 B.n993 585
R622 B.n75 B.n74 585
R623 B.n992 B.n75 585
R624 B.n990 B.n989 585
R625 B.n991 B.n990 585
R626 B.n988 B.n80 585
R627 B.n80 B.n79 585
R628 B.n987 B.n986 585
R629 B.n986 B.n985 585
R630 B.n82 B.n81 585
R631 B.n984 B.n82 585
R632 B.n982 B.n981 585
R633 B.n983 B.n982 585
R634 B.n980 B.n87 585
R635 B.n87 B.n86 585
R636 B.n979 B.n978 585
R637 B.n978 B.n977 585
R638 B.n89 B.n88 585
R639 B.n976 B.n89 585
R640 B.n974 B.n973 585
R641 B.n975 B.n974 585
R642 B.n972 B.n94 585
R643 B.n94 B.n93 585
R644 B.n971 B.n970 585
R645 B.n970 B.n969 585
R646 B.n96 B.n95 585
R647 B.n968 B.n96 585
R648 B.n966 B.n965 585
R649 B.n967 B.n966 585
R650 B.n964 B.n101 585
R651 B.n101 B.n100 585
R652 B.n963 B.n962 585
R653 B.n962 B.n961 585
R654 B.n103 B.n102 585
R655 B.n960 B.n103 585
R656 B.n1075 B.n1074 585
R657 B.n1073 B.n2 585
R658 B.n160 B.n103 564.573
R659 B.n958 B.n105 564.573
R660 B.n711 B.n463 564.573
R661 B.n707 B.n461 564.573
R662 B.n155 B.t12 377.115
R663 B.n516 B.t9 377.115
R664 B.n157 B.t15 377.115
R665 B.n514 B.t19 377.115
R666 B.n156 B.t13 295.272
R667 B.n517 B.t8 295.272
R668 B.n158 B.t16 295.272
R669 B.n515 B.t18 295.272
R670 B.n157 B.t14 288.466
R671 B.n155 B.t10 288.466
R672 B.n516 B.t6 288.466
R673 B.n514 B.t17 288.466
R674 B.n959 B.n153 256.663
R675 B.n959 B.n152 256.663
R676 B.n959 B.n151 256.663
R677 B.n959 B.n150 256.663
R678 B.n959 B.n149 256.663
R679 B.n959 B.n148 256.663
R680 B.n959 B.n147 256.663
R681 B.n959 B.n146 256.663
R682 B.n959 B.n145 256.663
R683 B.n959 B.n144 256.663
R684 B.n959 B.n143 256.663
R685 B.n959 B.n142 256.663
R686 B.n959 B.n141 256.663
R687 B.n959 B.n140 256.663
R688 B.n959 B.n139 256.663
R689 B.n959 B.n138 256.663
R690 B.n959 B.n137 256.663
R691 B.n959 B.n136 256.663
R692 B.n959 B.n135 256.663
R693 B.n959 B.n134 256.663
R694 B.n959 B.n133 256.663
R695 B.n959 B.n132 256.663
R696 B.n959 B.n131 256.663
R697 B.n959 B.n130 256.663
R698 B.n959 B.n129 256.663
R699 B.n959 B.n128 256.663
R700 B.n959 B.n127 256.663
R701 B.n959 B.n126 256.663
R702 B.n959 B.n125 256.663
R703 B.n959 B.n124 256.663
R704 B.n959 B.n123 256.663
R705 B.n959 B.n122 256.663
R706 B.n959 B.n121 256.663
R707 B.n959 B.n120 256.663
R708 B.n959 B.n119 256.663
R709 B.n959 B.n118 256.663
R710 B.n959 B.n117 256.663
R711 B.n959 B.n116 256.663
R712 B.n959 B.n115 256.663
R713 B.n959 B.n114 256.663
R714 B.n959 B.n113 256.663
R715 B.n959 B.n112 256.663
R716 B.n959 B.n111 256.663
R717 B.n959 B.n110 256.663
R718 B.n959 B.n109 256.663
R719 B.n959 B.n108 256.663
R720 B.n959 B.n107 256.663
R721 B.n959 B.n106 256.663
R722 B.n709 B.n708 256.663
R723 B.n709 B.n466 256.663
R724 B.n709 B.n467 256.663
R725 B.n709 B.n468 256.663
R726 B.n709 B.n469 256.663
R727 B.n709 B.n470 256.663
R728 B.n709 B.n471 256.663
R729 B.n709 B.n472 256.663
R730 B.n709 B.n473 256.663
R731 B.n709 B.n474 256.663
R732 B.n709 B.n475 256.663
R733 B.n709 B.n476 256.663
R734 B.n709 B.n477 256.663
R735 B.n709 B.n478 256.663
R736 B.n709 B.n479 256.663
R737 B.n709 B.n480 256.663
R738 B.n709 B.n481 256.663
R739 B.n709 B.n482 256.663
R740 B.n709 B.n483 256.663
R741 B.n709 B.n484 256.663
R742 B.n709 B.n485 256.663
R743 B.n709 B.n486 256.663
R744 B.n709 B.n487 256.663
R745 B.n709 B.n488 256.663
R746 B.n709 B.n489 256.663
R747 B.n709 B.n490 256.663
R748 B.n709 B.n491 256.663
R749 B.n709 B.n492 256.663
R750 B.n709 B.n493 256.663
R751 B.n709 B.n494 256.663
R752 B.n709 B.n495 256.663
R753 B.n709 B.n496 256.663
R754 B.n709 B.n497 256.663
R755 B.n709 B.n498 256.663
R756 B.n709 B.n499 256.663
R757 B.n709 B.n500 256.663
R758 B.n709 B.n501 256.663
R759 B.n709 B.n502 256.663
R760 B.n709 B.n503 256.663
R761 B.n709 B.n504 256.663
R762 B.n709 B.n505 256.663
R763 B.n709 B.n506 256.663
R764 B.n709 B.n507 256.663
R765 B.n709 B.n508 256.663
R766 B.n709 B.n509 256.663
R767 B.n709 B.n510 256.663
R768 B.n709 B.n511 256.663
R769 B.n710 B.n709 256.663
R770 B.n1077 B.n1076 256.663
R771 B.n164 B.n163 163.367
R772 B.n168 B.n167 163.367
R773 B.n172 B.n171 163.367
R774 B.n176 B.n175 163.367
R775 B.n180 B.n179 163.367
R776 B.n184 B.n183 163.367
R777 B.n188 B.n187 163.367
R778 B.n192 B.n191 163.367
R779 B.n196 B.n195 163.367
R780 B.n200 B.n199 163.367
R781 B.n204 B.n203 163.367
R782 B.n208 B.n207 163.367
R783 B.n212 B.n211 163.367
R784 B.n216 B.n215 163.367
R785 B.n220 B.n219 163.367
R786 B.n224 B.n223 163.367
R787 B.n228 B.n227 163.367
R788 B.n232 B.n231 163.367
R789 B.n236 B.n235 163.367
R790 B.n240 B.n239 163.367
R791 B.n244 B.n243 163.367
R792 B.n248 B.n247 163.367
R793 B.n252 B.n251 163.367
R794 B.n256 B.n255 163.367
R795 B.n260 B.n259 163.367
R796 B.n264 B.n263 163.367
R797 B.n269 B.n268 163.367
R798 B.n273 B.n272 163.367
R799 B.n277 B.n276 163.367
R800 B.n281 B.n280 163.367
R801 B.n285 B.n284 163.367
R802 B.n289 B.n288 163.367
R803 B.n293 B.n292 163.367
R804 B.n297 B.n296 163.367
R805 B.n301 B.n300 163.367
R806 B.n305 B.n304 163.367
R807 B.n309 B.n308 163.367
R808 B.n313 B.n312 163.367
R809 B.n317 B.n316 163.367
R810 B.n321 B.n320 163.367
R811 B.n325 B.n324 163.367
R812 B.n329 B.n328 163.367
R813 B.n333 B.n332 163.367
R814 B.n337 B.n336 163.367
R815 B.n341 B.n340 163.367
R816 B.n345 B.n344 163.367
R817 B.n349 B.n348 163.367
R818 B.n958 B.n154 163.367
R819 B.n715 B.n463 163.367
R820 B.n715 B.n457 163.367
R821 B.n723 B.n457 163.367
R822 B.n723 B.n455 163.367
R823 B.n727 B.n455 163.367
R824 B.n727 B.n449 163.367
R825 B.n735 B.n449 163.367
R826 B.n735 B.n447 163.367
R827 B.n739 B.n447 163.367
R828 B.n739 B.n441 163.367
R829 B.n747 B.n441 163.367
R830 B.n747 B.n439 163.367
R831 B.n751 B.n439 163.367
R832 B.n751 B.n433 163.367
R833 B.n759 B.n433 163.367
R834 B.n759 B.n431 163.367
R835 B.n763 B.n431 163.367
R836 B.n763 B.n425 163.367
R837 B.n771 B.n425 163.367
R838 B.n771 B.n423 163.367
R839 B.n775 B.n423 163.367
R840 B.n775 B.n416 163.367
R841 B.n783 B.n416 163.367
R842 B.n783 B.n414 163.367
R843 B.n787 B.n414 163.367
R844 B.n787 B.n409 163.367
R845 B.n795 B.n409 163.367
R846 B.n795 B.n407 163.367
R847 B.n799 B.n407 163.367
R848 B.n799 B.n401 163.367
R849 B.n807 B.n401 163.367
R850 B.n807 B.n399 163.367
R851 B.n811 B.n399 163.367
R852 B.n811 B.n393 163.367
R853 B.n819 B.n393 163.367
R854 B.n819 B.n391 163.367
R855 B.n823 B.n391 163.367
R856 B.n823 B.n385 163.367
R857 B.n831 B.n385 163.367
R858 B.n831 B.n383 163.367
R859 B.n835 B.n383 163.367
R860 B.n835 B.n377 163.367
R861 B.n843 B.n377 163.367
R862 B.n843 B.n375 163.367
R863 B.n847 B.n375 163.367
R864 B.n847 B.n369 163.367
R865 B.n855 B.n369 163.367
R866 B.n855 B.n367 163.367
R867 B.n859 B.n367 163.367
R868 B.n859 B.n361 163.367
R869 B.n867 B.n361 163.367
R870 B.n867 B.n359 163.367
R871 B.n872 B.n359 163.367
R872 B.n872 B.n353 163.367
R873 B.n880 B.n353 163.367
R874 B.n881 B.n880 163.367
R875 B.n881 B.n5 163.367
R876 B.n6 B.n5 163.367
R877 B.n7 B.n6 163.367
R878 B.n887 B.n7 163.367
R879 B.n888 B.n887 163.367
R880 B.n888 B.n13 163.367
R881 B.n14 B.n13 163.367
R882 B.n15 B.n14 163.367
R883 B.n893 B.n15 163.367
R884 B.n893 B.n20 163.367
R885 B.n21 B.n20 163.367
R886 B.n22 B.n21 163.367
R887 B.n898 B.n22 163.367
R888 B.n898 B.n27 163.367
R889 B.n28 B.n27 163.367
R890 B.n29 B.n28 163.367
R891 B.n903 B.n29 163.367
R892 B.n903 B.n34 163.367
R893 B.n35 B.n34 163.367
R894 B.n36 B.n35 163.367
R895 B.n908 B.n36 163.367
R896 B.n908 B.n41 163.367
R897 B.n42 B.n41 163.367
R898 B.n43 B.n42 163.367
R899 B.n913 B.n43 163.367
R900 B.n913 B.n48 163.367
R901 B.n49 B.n48 163.367
R902 B.n50 B.n49 163.367
R903 B.n918 B.n50 163.367
R904 B.n918 B.n55 163.367
R905 B.n56 B.n55 163.367
R906 B.n57 B.n56 163.367
R907 B.n923 B.n57 163.367
R908 B.n923 B.n62 163.367
R909 B.n63 B.n62 163.367
R910 B.n64 B.n63 163.367
R911 B.n928 B.n64 163.367
R912 B.n928 B.n69 163.367
R913 B.n70 B.n69 163.367
R914 B.n71 B.n70 163.367
R915 B.n933 B.n71 163.367
R916 B.n933 B.n76 163.367
R917 B.n77 B.n76 163.367
R918 B.n78 B.n77 163.367
R919 B.n938 B.n78 163.367
R920 B.n938 B.n83 163.367
R921 B.n84 B.n83 163.367
R922 B.n85 B.n84 163.367
R923 B.n943 B.n85 163.367
R924 B.n943 B.n90 163.367
R925 B.n91 B.n90 163.367
R926 B.n92 B.n91 163.367
R927 B.n948 B.n92 163.367
R928 B.n948 B.n97 163.367
R929 B.n98 B.n97 163.367
R930 B.n99 B.n98 163.367
R931 B.n953 B.n99 163.367
R932 B.n953 B.n104 163.367
R933 B.n105 B.n104 163.367
R934 B.n513 B.n512 163.367
R935 B.n702 B.n512 163.367
R936 B.n700 B.n699 163.367
R937 B.n696 B.n695 163.367
R938 B.n692 B.n691 163.367
R939 B.n688 B.n687 163.367
R940 B.n684 B.n683 163.367
R941 B.n680 B.n679 163.367
R942 B.n676 B.n675 163.367
R943 B.n672 B.n671 163.367
R944 B.n668 B.n667 163.367
R945 B.n664 B.n663 163.367
R946 B.n660 B.n659 163.367
R947 B.n656 B.n655 163.367
R948 B.n652 B.n651 163.367
R949 B.n648 B.n647 163.367
R950 B.n644 B.n643 163.367
R951 B.n640 B.n639 163.367
R952 B.n636 B.n635 163.367
R953 B.n632 B.n631 163.367
R954 B.n628 B.n627 163.367
R955 B.n624 B.n623 163.367
R956 B.n619 B.n618 163.367
R957 B.n615 B.n614 163.367
R958 B.n611 B.n610 163.367
R959 B.n607 B.n606 163.367
R960 B.n603 B.n602 163.367
R961 B.n599 B.n598 163.367
R962 B.n595 B.n594 163.367
R963 B.n591 B.n590 163.367
R964 B.n587 B.n586 163.367
R965 B.n583 B.n582 163.367
R966 B.n579 B.n578 163.367
R967 B.n575 B.n574 163.367
R968 B.n571 B.n570 163.367
R969 B.n567 B.n566 163.367
R970 B.n563 B.n562 163.367
R971 B.n559 B.n558 163.367
R972 B.n555 B.n554 163.367
R973 B.n551 B.n550 163.367
R974 B.n547 B.n546 163.367
R975 B.n543 B.n542 163.367
R976 B.n539 B.n538 163.367
R977 B.n535 B.n534 163.367
R978 B.n531 B.n530 163.367
R979 B.n527 B.n526 163.367
R980 B.n523 B.n522 163.367
R981 B.n519 B.n465 163.367
R982 B.n717 B.n461 163.367
R983 B.n717 B.n459 163.367
R984 B.n721 B.n459 163.367
R985 B.n721 B.n453 163.367
R986 B.n729 B.n453 163.367
R987 B.n729 B.n451 163.367
R988 B.n733 B.n451 163.367
R989 B.n733 B.n445 163.367
R990 B.n741 B.n445 163.367
R991 B.n741 B.n443 163.367
R992 B.n745 B.n443 163.367
R993 B.n745 B.n437 163.367
R994 B.n753 B.n437 163.367
R995 B.n753 B.n435 163.367
R996 B.n757 B.n435 163.367
R997 B.n757 B.n429 163.367
R998 B.n765 B.n429 163.367
R999 B.n765 B.n427 163.367
R1000 B.n769 B.n427 163.367
R1001 B.n769 B.n421 163.367
R1002 B.n777 B.n421 163.367
R1003 B.n777 B.n419 163.367
R1004 B.n781 B.n419 163.367
R1005 B.n781 B.n413 163.367
R1006 B.n789 B.n413 163.367
R1007 B.n789 B.n411 163.367
R1008 B.n793 B.n411 163.367
R1009 B.n793 B.n405 163.367
R1010 B.n801 B.n405 163.367
R1011 B.n801 B.n403 163.367
R1012 B.n805 B.n403 163.367
R1013 B.n805 B.n397 163.367
R1014 B.n813 B.n397 163.367
R1015 B.n813 B.n395 163.367
R1016 B.n817 B.n395 163.367
R1017 B.n817 B.n389 163.367
R1018 B.n825 B.n389 163.367
R1019 B.n825 B.n387 163.367
R1020 B.n829 B.n387 163.367
R1021 B.n829 B.n381 163.367
R1022 B.n837 B.n381 163.367
R1023 B.n837 B.n379 163.367
R1024 B.n841 B.n379 163.367
R1025 B.n841 B.n373 163.367
R1026 B.n849 B.n373 163.367
R1027 B.n849 B.n371 163.367
R1028 B.n853 B.n371 163.367
R1029 B.n853 B.n365 163.367
R1030 B.n861 B.n365 163.367
R1031 B.n861 B.n363 163.367
R1032 B.n865 B.n363 163.367
R1033 B.n865 B.n357 163.367
R1034 B.n874 B.n357 163.367
R1035 B.n874 B.n355 163.367
R1036 B.n878 B.n355 163.367
R1037 B.n878 B.n3 163.367
R1038 B.n1075 B.n3 163.367
R1039 B.n1071 B.n2 163.367
R1040 B.n1071 B.n1070 163.367
R1041 B.n1070 B.n9 163.367
R1042 B.n1066 B.n9 163.367
R1043 B.n1066 B.n11 163.367
R1044 B.n1062 B.n11 163.367
R1045 B.n1062 B.n17 163.367
R1046 B.n1058 B.n17 163.367
R1047 B.n1058 B.n19 163.367
R1048 B.n1054 B.n19 163.367
R1049 B.n1054 B.n24 163.367
R1050 B.n1050 B.n24 163.367
R1051 B.n1050 B.n26 163.367
R1052 B.n1046 B.n26 163.367
R1053 B.n1046 B.n31 163.367
R1054 B.n1042 B.n31 163.367
R1055 B.n1042 B.n33 163.367
R1056 B.n1038 B.n33 163.367
R1057 B.n1038 B.n38 163.367
R1058 B.n1034 B.n38 163.367
R1059 B.n1034 B.n40 163.367
R1060 B.n1030 B.n40 163.367
R1061 B.n1030 B.n45 163.367
R1062 B.n1026 B.n45 163.367
R1063 B.n1026 B.n47 163.367
R1064 B.n1022 B.n47 163.367
R1065 B.n1022 B.n52 163.367
R1066 B.n1018 B.n52 163.367
R1067 B.n1018 B.n54 163.367
R1068 B.n1014 B.n54 163.367
R1069 B.n1014 B.n59 163.367
R1070 B.n1010 B.n59 163.367
R1071 B.n1010 B.n61 163.367
R1072 B.n1006 B.n61 163.367
R1073 B.n1006 B.n66 163.367
R1074 B.n1002 B.n66 163.367
R1075 B.n1002 B.n68 163.367
R1076 B.n998 B.n68 163.367
R1077 B.n998 B.n73 163.367
R1078 B.n994 B.n73 163.367
R1079 B.n994 B.n75 163.367
R1080 B.n990 B.n75 163.367
R1081 B.n990 B.n80 163.367
R1082 B.n986 B.n80 163.367
R1083 B.n986 B.n82 163.367
R1084 B.n982 B.n82 163.367
R1085 B.n982 B.n87 163.367
R1086 B.n978 B.n87 163.367
R1087 B.n978 B.n89 163.367
R1088 B.n974 B.n89 163.367
R1089 B.n974 B.n94 163.367
R1090 B.n970 B.n94 163.367
R1091 B.n970 B.n96 163.367
R1092 B.n966 B.n96 163.367
R1093 B.n966 B.n101 163.367
R1094 B.n962 B.n101 163.367
R1095 B.n962 B.n103 163.367
R1096 B.n709 B.n462 85.9999
R1097 B.n960 B.n959 85.9999
R1098 B.n158 B.n157 81.8429
R1099 B.n156 B.n155 81.8429
R1100 B.n517 B.n516 81.8429
R1101 B.n515 B.n514 81.8429
R1102 B.n160 B.n106 71.676
R1103 B.n164 B.n107 71.676
R1104 B.n168 B.n108 71.676
R1105 B.n172 B.n109 71.676
R1106 B.n176 B.n110 71.676
R1107 B.n180 B.n111 71.676
R1108 B.n184 B.n112 71.676
R1109 B.n188 B.n113 71.676
R1110 B.n192 B.n114 71.676
R1111 B.n196 B.n115 71.676
R1112 B.n200 B.n116 71.676
R1113 B.n204 B.n117 71.676
R1114 B.n208 B.n118 71.676
R1115 B.n212 B.n119 71.676
R1116 B.n216 B.n120 71.676
R1117 B.n220 B.n121 71.676
R1118 B.n224 B.n122 71.676
R1119 B.n228 B.n123 71.676
R1120 B.n232 B.n124 71.676
R1121 B.n236 B.n125 71.676
R1122 B.n240 B.n126 71.676
R1123 B.n244 B.n127 71.676
R1124 B.n248 B.n128 71.676
R1125 B.n252 B.n129 71.676
R1126 B.n256 B.n130 71.676
R1127 B.n260 B.n131 71.676
R1128 B.n264 B.n132 71.676
R1129 B.n269 B.n133 71.676
R1130 B.n273 B.n134 71.676
R1131 B.n277 B.n135 71.676
R1132 B.n281 B.n136 71.676
R1133 B.n285 B.n137 71.676
R1134 B.n289 B.n138 71.676
R1135 B.n293 B.n139 71.676
R1136 B.n297 B.n140 71.676
R1137 B.n301 B.n141 71.676
R1138 B.n305 B.n142 71.676
R1139 B.n309 B.n143 71.676
R1140 B.n313 B.n144 71.676
R1141 B.n317 B.n145 71.676
R1142 B.n321 B.n146 71.676
R1143 B.n325 B.n147 71.676
R1144 B.n329 B.n148 71.676
R1145 B.n333 B.n149 71.676
R1146 B.n337 B.n150 71.676
R1147 B.n341 B.n151 71.676
R1148 B.n345 B.n152 71.676
R1149 B.n349 B.n153 71.676
R1150 B.n154 B.n153 71.676
R1151 B.n348 B.n152 71.676
R1152 B.n344 B.n151 71.676
R1153 B.n340 B.n150 71.676
R1154 B.n336 B.n149 71.676
R1155 B.n332 B.n148 71.676
R1156 B.n328 B.n147 71.676
R1157 B.n324 B.n146 71.676
R1158 B.n320 B.n145 71.676
R1159 B.n316 B.n144 71.676
R1160 B.n312 B.n143 71.676
R1161 B.n308 B.n142 71.676
R1162 B.n304 B.n141 71.676
R1163 B.n300 B.n140 71.676
R1164 B.n296 B.n139 71.676
R1165 B.n292 B.n138 71.676
R1166 B.n288 B.n137 71.676
R1167 B.n284 B.n136 71.676
R1168 B.n280 B.n135 71.676
R1169 B.n276 B.n134 71.676
R1170 B.n272 B.n133 71.676
R1171 B.n268 B.n132 71.676
R1172 B.n263 B.n131 71.676
R1173 B.n259 B.n130 71.676
R1174 B.n255 B.n129 71.676
R1175 B.n251 B.n128 71.676
R1176 B.n247 B.n127 71.676
R1177 B.n243 B.n126 71.676
R1178 B.n239 B.n125 71.676
R1179 B.n235 B.n124 71.676
R1180 B.n231 B.n123 71.676
R1181 B.n227 B.n122 71.676
R1182 B.n223 B.n121 71.676
R1183 B.n219 B.n120 71.676
R1184 B.n215 B.n119 71.676
R1185 B.n211 B.n118 71.676
R1186 B.n207 B.n117 71.676
R1187 B.n203 B.n116 71.676
R1188 B.n199 B.n115 71.676
R1189 B.n195 B.n114 71.676
R1190 B.n191 B.n113 71.676
R1191 B.n187 B.n112 71.676
R1192 B.n183 B.n111 71.676
R1193 B.n179 B.n110 71.676
R1194 B.n175 B.n109 71.676
R1195 B.n171 B.n108 71.676
R1196 B.n167 B.n107 71.676
R1197 B.n163 B.n106 71.676
R1198 B.n708 B.n707 71.676
R1199 B.n702 B.n466 71.676
R1200 B.n699 B.n467 71.676
R1201 B.n695 B.n468 71.676
R1202 B.n691 B.n469 71.676
R1203 B.n687 B.n470 71.676
R1204 B.n683 B.n471 71.676
R1205 B.n679 B.n472 71.676
R1206 B.n675 B.n473 71.676
R1207 B.n671 B.n474 71.676
R1208 B.n667 B.n475 71.676
R1209 B.n663 B.n476 71.676
R1210 B.n659 B.n477 71.676
R1211 B.n655 B.n478 71.676
R1212 B.n651 B.n479 71.676
R1213 B.n647 B.n480 71.676
R1214 B.n643 B.n481 71.676
R1215 B.n639 B.n482 71.676
R1216 B.n635 B.n483 71.676
R1217 B.n631 B.n484 71.676
R1218 B.n627 B.n485 71.676
R1219 B.n623 B.n486 71.676
R1220 B.n618 B.n487 71.676
R1221 B.n614 B.n488 71.676
R1222 B.n610 B.n489 71.676
R1223 B.n606 B.n490 71.676
R1224 B.n602 B.n491 71.676
R1225 B.n598 B.n492 71.676
R1226 B.n594 B.n493 71.676
R1227 B.n590 B.n494 71.676
R1228 B.n586 B.n495 71.676
R1229 B.n582 B.n496 71.676
R1230 B.n578 B.n497 71.676
R1231 B.n574 B.n498 71.676
R1232 B.n570 B.n499 71.676
R1233 B.n566 B.n500 71.676
R1234 B.n562 B.n501 71.676
R1235 B.n558 B.n502 71.676
R1236 B.n554 B.n503 71.676
R1237 B.n550 B.n504 71.676
R1238 B.n546 B.n505 71.676
R1239 B.n542 B.n506 71.676
R1240 B.n538 B.n507 71.676
R1241 B.n534 B.n508 71.676
R1242 B.n530 B.n509 71.676
R1243 B.n526 B.n510 71.676
R1244 B.n522 B.n511 71.676
R1245 B.n710 B.n465 71.676
R1246 B.n708 B.n513 71.676
R1247 B.n700 B.n466 71.676
R1248 B.n696 B.n467 71.676
R1249 B.n692 B.n468 71.676
R1250 B.n688 B.n469 71.676
R1251 B.n684 B.n470 71.676
R1252 B.n680 B.n471 71.676
R1253 B.n676 B.n472 71.676
R1254 B.n672 B.n473 71.676
R1255 B.n668 B.n474 71.676
R1256 B.n664 B.n475 71.676
R1257 B.n660 B.n476 71.676
R1258 B.n656 B.n477 71.676
R1259 B.n652 B.n478 71.676
R1260 B.n648 B.n479 71.676
R1261 B.n644 B.n480 71.676
R1262 B.n640 B.n481 71.676
R1263 B.n636 B.n482 71.676
R1264 B.n632 B.n483 71.676
R1265 B.n628 B.n484 71.676
R1266 B.n624 B.n485 71.676
R1267 B.n619 B.n486 71.676
R1268 B.n615 B.n487 71.676
R1269 B.n611 B.n488 71.676
R1270 B.n607 B.n489 71.676
R1271 B.n603 B.n490 71.676
R1272 B.n599 B.n491 71.676
R1273 B.n595 B.n492 71.676
R1274 B.n591 B.n493 71.676
R1275 B.n587 B.n494 71.676
R1276 B.n583 B.n495 71.676
R1277 B.n579 B.n496 71.676
R1278 B.n575 B.n497 71.676
R1279 B.n571 B.n498 71.676
R1280 B.n567 B.n499 71.676
R1281 B.n563 B.n500 71.676
R1282 B.n559 B.n501 71.676
R1283 B.n555 B.n502 71.676
R1284 B.n551 B.n503 71.676
R1285 B.n547 B.n504 71.676
R1286 B.n543 B.n505 71.676
R1287 B.n539 B.n506 71.676
R1288 B.n535 B.n507 71.676
R1289 B.n531 B.n508 71.676
R1290 B.n527 B.n509 71.676
R1291 B.n523 B.n510 71.676
R1292 B.n519 B.n511 71.676
R1293 B.n711 B.n710 71.676
R1294 B.n1076 B.n1075 71.676
R1295 B.n1076 B.n2 71.676
R1296 B.n159 B.n158 59.5399
R1297 B.n266 B.n156 59.5399
R1298 B.n518 B.n517 59.5399
R1299 B.n621 B.n515 59.5399
R1300 B.n716 B.n462 41.4754
R1301 B.n716 B.n458 41.4754
R1302 B.n722 B.n458 41.4754
R1303 B.n722 B.n454 41.4754
R1304 B.n728 B.n454 41.4754
R1305 B.n728 B.n450 41.4754
R1306 B.n734 B.n450 41.4754
R1307 B.n734 B.n446 41.4754
R1308 B.n740 B.n446 41.4754
R1309 B.n746 B.n442 41.4754
R1310 B.n746 B.n438 41.4754
R1311 B.n752 B.n438 41.4754
R1312 B.n752 B.n434 41.4754
R1313 B.n758 B.n434 41.4754
R1314 B.n758 B.n430 41.4754
R1315 B.n764 B.n430 41.4754
R1316 B.n764 B.n426 41.4754
R1317 B.n770 B.n426 41.4754
R1318 B.n770 B.n422 41.4754
R1319 B.n776 B.n422 41.4754
R1320 B.n776 B.n417 41.4754
R1321 B.n782 B.n417 41.4754
R1322 B.n782 B.n418 41.4754
R1323 B.n788 B.n410 41.4754
R1324 B.n794 B.n410 41.4754
R1325 B.n794 B.n406 41.4754
R1326 B.n800 B.n406 41.4754
R1327 B.n800 B.n402 41.4754
R1328 B.n806 B.n402 41.4754
R1329 B.n806 B.n398 41.4754
R1330 B.n812 B.n398 41.4754
R1331 B.n812 B.n394 41.4754
R1332 B.n818 B.n394 41.4754
R1333 B.n818 B.n390 41.4754
R1334 B.n824 B.n390 41.4754
R1335 B.n830 B.n386 41.4754
R1336 B.n830 B.n382 41.4754
R1337 B.n836 B.n382 41.4754
R1338 B.n836 B.n378 41.4754
R1339 B.n842 B.n378 41.4754
R1340 B.n842 B.n374 41.4754
R1341 B.n848 B.n374 41.4754
R1342 B.n848 B.n370 41.4754
R1343 B.n854 B.n370 41.4754
R1344 B.n854 B.n366 41.4754
R1345 B.n860 B.n366 41.4754
R1346 B.n866 B.n362 41.4754
R1347 B.n866 B.n358 41.4754
R1348 B.n873 B.n358 41.4754
R1349 B.n873 B.n354 41.4754
R1350 B.n879 B.n354 41.4754
R1351 B.n879 B.n4 41.4754
R1352 B.n1074 B.n4 41.4754
R1353 B.n1074 B.n1073 41.4754
R1354 B.n1073 B.n1072 41.4754
R1355 B.n1072 B.n8 41.4754
R1356 B.n12 B.n8 41.4754
R1357 B.n1065 B.n12 41.4754
R1358 B.n1065 B.n1064 41.4754
R1359 B.n1064 B.n1063 41.4754
R1360 B.n1063 B.n16 41.4754
R1361 B.n1057 B.n1056 41.4754
R1362 B.n1056 B.n1055 41.4754
R1363 B.n1055 B.n23 41.4754
R1364 B.n1049 B.n23 41.4754
R1365 B.n1049 B.n1048 41.4754
R1366 B.n1048 B.n1047 41.4754
R1367 B.n1047 B.n30 41.4754
R1368 B.n1041 B.n30 41.4754
R1369 B.n1041 B.n1040 41.4754
R1370 B.n1040 B.n1039 41.4754
R1371 B.n1039 B.n37 41.4754
R1372 B.n1033 B.n1032 41.4754
R1373 B.n1032 B.n1031 41.4754
R1374 B.n1031 B.n44 41.4754
R1375 B.n1025 B.n44 41.4754
R1376 B.n1025 B.n1024 41.4754
R1377 B.n1024 B.n1023 41.4754
R1378 B.n1023 B.n51 41.4754
R1379 B.n1017 B.n51 41.4754
R1380 B.n1017 B.n1016 41.4754
R1381 B.n1016 B.n1015 41.4754
R1382 B.n1015 B.n58 41.4754
R1383 B.n1009 B.n58 41.4754
R1384 B.n1008 B.n1007 41.4754
R1385 B.n1007 B.n65 41.4754
R1386 B.n1001 B.n65 41.4754
R1387 B.n1001 B.n1000 41.4754
R1388 B.n1000 B.n999 41.4754
R1389 B.n999 B.n72 41.4754
R1390 B.n993 B.n72 41.4754
R1391 B.n993 B.n992 41.4754
R1392 B.n992 B.n991 41.4754
R1393 B.n991 B.n79 41.4754
R1394 B.n985 B.n79 41.4754
R1395 B.n985 B.n984 41.4754
R1396 B.n984 B.n983 41.4754
R1397 B.n983 B.n86 41.4754
R1398 B.n977 B.n976 41.4754
R1399 B.n976 B.n975 41.4754
R1400 B.n975 B.n93 41.4754
R1401 B.n969 B.n93 41.4754
R1402 B.n969 B.n968 41.4754
R1403 B.n968 B.n967 41.4754
R1404 B.n967 B.n100 41.4754
R1405 B.n961 B.n100 41.4754
R1406 B.n961 B.n960 41.4754
R1407 B.n706 B.n460 36.6834
R1408 B.n713 B.n712 36.6834
R1409 B.n957 B.n956 36.6834
R1410 B.n161 B.n102 36.6834
R1411 B.n418 B.t5 35.9861
R1412 B.t2 B.n1008 35.9861
R1413 B.t7 B.n442 31.1067
R1414 B.t11 B.n86 31.1067
R1415 B.t4 B.n386 29.8868
R1416 B.t0 B.n37 29.8868
R1417 B.n860 B.t3 28.667
R1418 B.n1057 B.t1 28.667
R1419 B B.n1077 18.0485
R1420 B.t3 B.n362 12.8089
R1421 B.t1 B.n16 12.8089
R1422 B.n824 B.t4 11.5891
R1423 B.n1033 B.t0 11.5891
R1424 B.n718 B.n460 10.6151
R1425 B.n719 B.n718 10.6151
R1426 B.n720 B.n719 10.6151
R1427 B.n720 B.n452 10.6151
R1428 B.n730 B.n452 10.6151
R1429 B.n731 B.n730 10.6151
R1430 B.n732 B.n731 10.6151
R1431 B.n732 B.n444 10.6151
R1432 B.n742 B.n444 10.6151
R1433 B.n743 B.n742 10.6151
R1434 B.n744 B.n743 10.6151
R1435 B.n744 B.n436 10.6151
R1436 B.n754 B.n436 10.6151
R1437 B.n755 B.n754 10.6151
R1438 B.n756 B.n755 10.6151
R1439 B.n756 B.n428 10.6151
R1440 B.n766 B.n428 10.6151
R1441 B.n767 B.n766 10.6151
R1442 B.n768 B.n767 10.6151
R1443 B.n768 B.n420 10.6151
R1444 B.n778 B.n420 10.6151
R1445 B.n779 B.n778 10.6151
R1446 B.n780 B.n779 10.6151
R1447 B.n780 B.n412 10.6151
R1448 B.n790 B.n412 10.6151
R1449 B.n791 B.n790 10.6151
R1450 B.n792 B.n791 10.6151
R1451 B.n792 B.n404 10.6151
R1452 B.n802 B.n404 10.6151
R1453 B.n803 B.n802 10.6151
R1454 B.n804 B.n803 10.6151
R1455 B.n804 B.n396 10.6151
R1456 B.n814 B.n396 10.6151
R1457 B.n815 B.n814 10.6151
R1458 B.n816 B.n815 10.6151
R1459 B.n816 B.n388 10.6151
R1460 B.n826 B.n388 10.6151
R1461 B.n827 B.n826 10.6151
R1462 B.n828 B.n827 10.6151
R1463 B.n828 B.n380 10.6151
R1464 B.n838 B.n380 10.6151
R1465 B.n839 B.n838 10.6151
R1466 B.n840 B.n839 10.6151
R1467 B.n840 B.n372 10.6151
R1468 B.n850 B.n372 10.6151
R1469 B.n851 B.n850 10.6151
R1470 B.n852 B.n851 10.6151
R1471 B.n852 B.n364 10.6151
R1472 B.n862 B.n364 10.6151
R1473 B.n863 B.n862 10.6151
R1474 B.n864 B.n863 10.6151
R1475 B.n864 B.n356 10.6151
R1476 B.n875 B.n356 10.6151
R1477 B.n876 B.n875 10.6151
R1478 B.n877 B.n876 10.6151
R1479 B.n877 B.n0 10.6151
R1480 B.n706 B.n705 10.6151
R1481 B.n705 B.n704 10.6151
R1482 B.n704 B.n703 10.6151
R1483 B.n703 B.n701 10.6151
R1484 B.n701 B.n698 10.6151
R1485 B.n698 B.n697 10.6151
R1486 B.n697 B.n694 10.6151
R1487 B.n694 B.n693 10.6151
R1488 B.n693 B.n690 10.6151
R1489 B.n690 B.n689 10.6151
R1490 B.n689 B.n686 10.6151
R1491 B.n686 B.n685 10.6151
R1492 B.n685 B.n682 10.6151
R1493 B.n682 B.n681 10.6151
R1494 B.n681 B.n678 10.6151
R1495 B.n678 B.n677 10.6151
R1496 B.n677 B.n674 10.6151
R1497 B.n674 B.n673 10.6151
R1498 B.n673 B.n670 10.6151
R1499 B.n670 B.n669 10.6151
R1500 B.n669 B.n666 10.6151
R1501 B.n666 B.n665 10.6151
R1502 B.n665 B.n662 10.6151
R1503 B.n662 B.n661 10.6151
R1504 B.n661 B.n658 10.6151
R1505 B.n658 B.n657 10.6151
R1506 B.n657 B.n654 10.6151
R1507 B.n654 B.n653 10.6151
R1508 B.n653 B.n650 10.6151
R1509 B.n650 B.n649 10.6151
R1510 B.n649 B.n646 10.6151
R1511 B.n646 B.n645 10.6151
R1512 B.n645 B.n642 10.6151
R1513 B.n642 B.n641 10.6151
R1514 B.n641 B.n638 10.6151
R1515 B.n638 B.n637 10.6151
R1516 B.n637 B.n634 10.6151
R1517 B.n634 B.n633 10.6151
R1518 B.n633 B.n630 10.6151
R1519 B.n630 B.n629 10.6151
R1520 B.n629 B.n626 10.6151
R1521 B.n626 B.n625 10.6151
R1522 B.n625 B.n622 10.6151
R1523 B.n620 B.n617 10.6151
R1524 B.n617 B.n616 10.6151
R1525 B.n616 B.n613 10.6151
R1526 B.n613 B.n612 10.6151
R1527 B.n612 B.n609 10.6151
R1528 B.n609 B.n608 10.6151
R1529 B.n608 B.n605 10.6151
R1530 B.n605 B.n604 10.6151
R1531 B.n601 B.n600 10.6151
R1532 B.n600 B.n597 10.6151
R1533 B.n597 B.n596 10.6151
R1534 B.n596 B.n593 10.6151
R1535 B.n593 B.n592 10.6151
R1536 B.n592 B.n589 10.6151
R1537 B.n589 B.n588 10.6151
R1538 B.n588 B.n585 10.6151
R1539 B.n585 B.n584 10.6151
R1540 B.n584 B.n581 10.6151
R1541 B.n581 B.n580 10.6151
R1542 B.n580 B.n577 10.6151
R1543 B.n577 B.n576 10.6151
R1544 B.n576 B.n573 10.6151
R1545 B.n573 B.n572 10.6151
R1546 B.n572 B.n569 10.6151
R1547 B.n569 B.n568 10.6151
R1548 B.n568 B.n565 10.6151
R1549 B.n565 B.n564 10.6151
R1550 B.n564 B.n561 10.6151
R1551 B.n561 B.n560 10.6151
R1552 B.n560 B.n557 10.6151
R1553 B.n557 B.n556 10.6151
R1554 B.n556 B.n553 10.6151
R1555 B.n553 B.n552 10.6151
R1556 B.n552 B.n549 10.6151
R1557 B.n549 B.n548 10.6151
R1558 B.n548 B.n545 10.6151
R1559 B.n545 B.n544 10.6151
R1560 B.n544 B.n541 10.6151
R1561 B.n541 B.n540 10.6151
R1562 B.n540 B.n537 10.6151
R1563 B.n537 B.n536 10.6151
R1564 B.n536 B.n533 10.6151
R1565 B.n533 B.n532 10.6151
R1566 B.n532 B.n529 10.6151
R1567 B.n529 B.n528 10.6151
R1568 B.n528 B.n525 10.6151
R1569 B.n525 B.n524 10.6151
R1570 B.n524 B.n521 10.6151
R1571 B.n521 B.n520 10.6151
R1572 B.n520 B.n464 10.6151
R1573 B.n712 B.n464 10.6151
R1574 B.n714 B.n713 10.6151
R1575 B.n714 B.n456 10.6151
R1576 B.n724 B.n456 10.6151
R1577 B.n725 B.n724 10.6151
R1578 B.n726 B.n725 10.6151
R1579 B.n726 B.n448 10.6151
R1580 B.n736 B.n448 10.6151
R1581 B.n737 B.n736 10.6151
R1582 B.n738 B.n737 10.6151
R1583 B.n738 B.n440 10.6151
R1584 B.n748 B.n440 10.6151
R1585 B.n749 B.n748 10.6151
R1586 B.n750 B.n749 10.6151
R1587 B.n750 B.n432 10.6151
R1588 B.n760 B.n432 10.6151
R1589 B.n761 B.n760 10.6151
R1590 B.n762 B.n761 10.6151
R1591 B.n762 B.n424 10.6151
R1592 B.n772 B.n424 10.6151
R1593 B.n773 B.n772 10.6151
R1594 B.n774 B.n773 10.6151
R1595 B.n774 B.n415 10.6151
R1596 B.n784 B.n415 10.6151
R1597 B.n785 B.n784 10.6151
R1598 B.n786 B.n785 10.6151
R1599 B.n786 B.n408 10.6151
R1600 B.n796 B.n408 10.6151
R1601 B.n797 B.n796 10.6151
R1602 B.n798 B.n797 10.6151
R1603 B.n798 B.n400 10.6151
R1604 B.n808 B.n400 10.6151
R1605 B.n809 B.n808 10.6151
R1606 B.n810 B.n809 10.6151
R1607 B.n810 B.n392 10.6151
R1608 B.n820 B.n392 10.6151
R1609 B.n821 B.n820 10.6151
R1610 B.n822 B.n821 10.6151
R1611 B.n822 B.n384 10.6151
R1612 B.n832 B.n384 10.6151
R1613 B.n833 B.n832 10.6151
R1614 B.n834 B.n833 10.6151
R1615 B.n834 B.n376 10.6151
R1616 B.n844 B.n376 10.6151
R1617 B.n845 B.n844 10.6151
R1618 B.n846 B.n845 10.6151
R1619 B.n846 B.n368 10.6151
R1620 B.n856 B.n368 10.6151
R1621 B.n857 B.n856 10.6151
R1622 B.n858 B.n857 10.6151
R1623 B.n858 B.n360 10.6151
R1624 B.n868 B.n360 10.6151
R1625 B.n869 B.n868 10.6151
R1626 B.n871 B.n869 10.6151
R1627 B.n871 B.n870 10.6151
R1628 B.n870 B.n352 10.6151
R1629 B.n882 B.n352 10.6151
R1630 B.n883 B.n882 10.6151
R1631 B.n884 B.n883 10.6151
R1632 B.n885 B.n884 10.6151
R1633 B.n886 B.n885 10.6151
R1634 B.n889 B.n886 10.6151
R1635 B.n890 B.n889 10.6151
R1636 B.n891 B.n890 10.6151
R1637 B.n892 B.n891 10.6151
R1638 B.n894 B.n892 10.6151
R1639 B.n895 B.n894 10.6151
R1640 B.n896 B.n895 10.6151
R1641 B.n897 B.n896 10.6151
R1642 B.n899 B.n897 10.6151
R1643 B.n900 B.n899 10.6151
R1644 B.n901 B.n900 10.6151
R1645 B.n902 B.n901 10.6151
R1646 B.n904 B.n902 10.6151
R1647 B.n905 B.n904 10.6151
R1648 B.n906 B.n905 10.6151
R1649 B.n907 B.n906 10.6151
R1650 B.n909 B.n907 10.6151
R1651 B.n910 B.n909 10.6151
R1652 B.n911 B.n910 10.6151
R1653 B.n912 B.n911 10.6151
R1654 B.n914 B.n912 10.6151
R1655 B.n915 B.n914 10.6151
R1656 B.n916 B.n915 10.6151
R1657 B.n917 B.n916 10.6151
R1658 B.n919 B.n917 10.6151
R1659 B.n920 B.n919 10.6151
R1660 B.n921 B.n920 10.6151
R1661 B.n922 B.n921 10.6151
R1662 B.n924 B.n922 10.6151
R1663 B.n925 B.n924 10.6151
R1664 B.n926 B.n925 10.6151
R1665 B.n927 B.n926 10.6151
R1666 B.n929 B.n927 10.6151
R1667 B.n930 B.n929 10.6151
R1668 B.n931 B.n930 10.6151
R1669 B.n932 B.n931 10.6151
R1670 B.n934 B.n932 10.6151
R1671 B.n935 B.n934 10.6151
R1672 B.n936 B.n935 10.6151
R1673 B.n937 B.n936 10.6151
R1674 B.n939 B.n937 10.6151
R1675 B.n940 B.n939 10.6151
R1676 B.n941 B.n940 10.6151
R1677 B.n942 B.n941 10.6151
R1678 B.n944 B.n942 10.6151
R1679 B.n945 B.n944 10.6151
R1680 B.n946 B.n945 10.6151
R1681 B.n947 B.n946 10.6151
R1682 B.n949 B.n947 10.6151
R1683 B.n950 B.n949 10.6151
R1684 B.n951 B.n950 10.6151
R1685 B.n952 B.n951 10.6151
R1686 B.n954 B.n952 10.6151
R1687 B.n955 B.n954 10.6151
R1688 B.n956 B.n955 10.6151
R1689 B.n1069 B.n1 10.6151
R1690 B.n1069 B.n1068 10.6151
R1691 B.n1068 B.n1067 10.6151
R1692 B.n1067 B.n10 10.6151
R1693 B.n1061 B.n10 10.6151
R1694 B.n1061 B.n1060 10.6151
R1695 B.n1060 B.n1059 10.6151
R1696 B.n1059 B.n18 10.6151
R1697 B.n1053 B.n18 10.6151
R1698 B.n1053 B.n1052 10.6151
R1699 B.n1052 B.n1051 10.6151
R1700 B.n1051 B.n25 10.6151
R1701 B.n1045 B.n25 10.6151
R1702 B.n1045 B.n1044 10.6151
R1703 B.n1044 B.n1043 10.6151
R1704 B.n1043 B.n32 10.6151
R1705 B.n1037 B.n32 10.6151
R1706 B.n1037 B.n1036 10.6151
R1707 B.n1036 B.n1035 10.6151
R1708 B.n1035 B.n39 10.6151
R1709 B.n1029 B.n39 10.6151
R1710 B.n1029 B.n1028 10.6151
R1711 B.n1028 B.n1027 10.6151
R1712 B.n1027 B.n46 10.6151
R1713 B.n1021 B.n46 10.6151
R1714 B.n1021 B.n1020 10.6151
R1715 B.n1020 B.n1019 10.6151
R1716 B.n1019 B.n53 10.6151
R1717 B.n1013 B.n53 10.6151
R1718 B.n1013 B.n1012 10.6151
R1719 B.n1012 B.n1011 10.6151
R1720 B.n1011 B.n60 10.6151
R1721 B.n1005 B.n60 10.6151
R1722 B.n1005 B.n1004 10.6151
R1723 B.n1004 B.n1003 10.6151
R1724 B.n1003 B.n67 10.6151
R1725 B.n997 B.n67 10.6151
R1726 B.n997 B.n996 10.6151
R1727 B.n996 B.n995 10.6151
R1728 B.n995 B.n74 10.6151
R1729 B.n989 B.n74 10.6151
R1730 B.n989 B.n988 10.6151
R1731 B.n988 B.n987 10.6151
R1732 B.n987 B.n81 10.6151
R1733 B.n981 B.n81 10.6151
R1734 B.n981 B.n980 10.6151
R1735 B.n980 B.n979 10.6151
R1736 B.n979 B.n88 10.6151
R1737 B.n973 B.n88 10.6151
R1738 B.n973 B.n972 10.6151
R1739 B.n972 B.n971 10.6151
R1740 B.n971 B.n95 10.6151
R1741 B.n965 B.n95 10.6151
R1742 B.n965 B.n964 10.6151
R1743 B.n964 B.n963 10.6151
R1744 B.n963 B.n102 10.6151
R1745 B.n162 B.n161 10.6151
R1746 B.n165 B.n162 10.6151
R1747 B.n166 B.n165 10.6151
R1748 B.n169 B.n166 10.6151
R1749 B.n170 B.n169 10.6151
R1750 B.n173 B.n170 10.6151
R1751 B.n174 B.n173 10.6151
R1752 B.n177 B.n174 10.6151
R1753 B.n178 B.n177 10.6151
R1754 B.n181 B.n178 10.6151
R1755 B.n182 B.n181 10.6151
R1756 B.n185 B.n182 10.6151
R1757 B.n186 B.n185 10.6151
R1758 B.n189 B.n186 10.6151
R1759 B.n190 B.n189 10.6151
R1760 B.n193 B.n190 10.6151
R1761 B.n194 B.n193 10.6151
R1762 B.n197 B.n194 10.6151
R1763 B.n198 B.n197 10.6151
R1764 B.n201 B.n198 10.6151
R1765 B.n202 B.n201 10.6151
R1766 B.n205 B.n202 10.6151
R1767 B.n206 B.n205 10.6151
R1768 B.n209 B.n206 10.6151
R1769 B.n210 B.n209 10.6151
R1770 B.n213 B.n210 10.6151
R1771 B.n214 B.n213 10.6151
R1772 B.n217 B.n214 10.6151
R1773 B.n218 B.n217 10.6151
R1774 B.n221 B.n218 10.6151
R1775 B.n222 B.n221 10.6151
R1776 B.n225 B.n222 10.6151
R1777 B.n226 B.n225 10.6151
R1778 B.n229 B.n226 10.6151
R1779 B.n230 B.n229 10.6151
R1780 B.n233 B.n230 10.6151
R1781 B.n234 B.n233 10.6151
R1782 B.n237 B.n234 10.6151
R1783 B.n238 B.n237 10.6151
R1784 B.n241 B.n238 10.6151
R1785 B.n242 B.n241 10.6151
R1786 B.n245 B.n242 10.6151
R1787 B.n246 B.n245 10.6151
R1788 B.n250 B.n249 10.6151
R1789 B.n253 B.n250 10.6151
R1790 B.n254 B.n253 10.6151
R1791 B.n257 B.n254 10.6151
R1792 B.n258 B.n257 10.6151
R1793 B.n261 B.n258 10.6151
R1794 B.n262 B.n261 10.6151
R1795 B.n265 B.n262 10.6151
R1796 B.n270 B.n267 10.6151
R1797 B.n271 B.n270 10.6151
R1798 B.n274 B.n271 10.6151
R1799 B.n275 B.n274 10.6151
R1800 B.n278 B.n275 10.6151
R1801 B.n279 B.n278 10.6151
R1802 B.n282 B.n279 10.6151
R1803 B.n283 B.n282 10.6151
R1804 B.n286 B.n283 10.6151
R1805 B.n287 B.n286 10.6151
R1806 B.n290 B.n287 10.6151
R1807 B.n291 B.n290 10.6151
R1808 B.n294 B.n291 10.6151
R1809 B.n295 B.n294 10.6151
R1810 B.n298 B.n295 10.6151
R1811 B.n299 B.n298 10.6151
R1812 B.n302 B.n299 10.6151
R1813 B.n303 B.n302 10.6151
R1814 B.n306 B.n303 10.6151
R1815 B.n307 B.n306 10.6151
R1816 B.n310 B.n307 10.6151
R1817 B.n311 B.n310 10.6151
R1818 B.n314 B.n311 10.6151
R1819 B.n315 B.n314 10.6151
R1820 B.n318 B.n315 10.6151
R1821 B.n319 B.n318 10.6151
R1822 B.n322 B.n319 10.6151
R1823 B.n323 B.n322 10.6151
R1824 B.n326 B.n323 10.6151
R1825 B.n327 B.n326 10.6151
R1826 B.n330 B.n327 10.6151
R1827 B.n331 B.n330 10.6151
R1828 B.n334 B.n331 10.6151
R1829 B.n335 B.n334 10.6151
R1830 B.n338 B.n335 10.6151
R1831 B.n339 B.n338 10.6151
R1832 B.n342 B.n339 10.6151
R1833 B.n343 B.n342 10.6151
R1834 B.n346 B.n343 10.6151
R1835 B.n347 B.n346 10.6151
R1836 B.n350 B.n347 10.6151
R1837 B.n351 B.n350 10.6151
R1838 B.n957 B.n351 10.6151
R1839 B.n740 B.t7 10.3692
R1840 B.n977 B.t11 10.3692
R1841 B.n1077 B.n0 8.11757
R1842 B.n1077 B.n1 8.11757
R1843 B.n621 B.n620 6.5566
R1844 B.n604 B.n518 6.5566
R1845 B.n249 B.n159 6.5566
R1846 B.n266 B.n265 6.5566
R1847 B.n788 B.t5 5.48983
R1848 B.n1009 B.t2 5.48983
R1849 B.n622 B.n621 4.05904
R1850 B.n601 B.n518 4.05904
R1851 B.n246 B.n159 4.05904
R1852 B.n267 B.n266 4.05904
R1853 VN.n37 VN.n20 161.3
R1854 VN.n36 VN.n35 161.3
R1855 VN.n34 VN.n21 161.3
R1856 VN.n33 VN.n32 161.3
R1857 VN.n31 VN.n22 161.3
R1858 VN.n30 VN.n29 161.3
R1859 VN.n28 VN.n23 161.3
R1860 VN.n27 VN.n26 161.3
R1861 VN.n17 VN.n0 161.3
R1862 VN.n16 VN.n15 161.3
R1863 VN.n14 VN.n1 161.3
R1864 VN.n13 VN.n12 161.3
R1865 VN.n11 VN.n2 161.3
R1866 VN.n10 VN.n9 161.3
R1867 VN.n8 VN.n3 161.3
R1868 VN.n7 VN.n6 161.3
R1869 VN.n4 VN.t1 111.249
R1870 VN.n24 VN.t4 111.249
R1871 VN.n5 VN.t0 79.0535
R1872 VN.n18 VN.t3 79.0535
R1873 VN.n25 VN.t5 79.0535
R1874 VN.n38 VN.t2 79.0535
R1875 VN.n5 VN.n4 63.0626
R1876 VN.n25 VN.n24 63.0626
R1877 VN.n19 VN.n18 59.2636
R1878 VN.n39 VN.n38 59.2636
R1879 VN VN.n39 54.6104
R1880 VN.n12 VN.n11 54.1398
R1881 VN.n32 VN.n31 54.1398
R1882 VN.n12 VN.n1 27.0143
R1883 VN.n32 VN.n21 27.0143
R1884 VN.n6 VN.n3 24.5923
R1885 VN.n10 VN.n3 24.5923
R1886 VN.n11 VN.n10 24.5923
R1887 VN.n16 VN.n1 24.5923
R1888 VN.n17 VN.n16 24.5923
R1889 VN.n31 VN.n30 24.5923
R1890 VN.n30 VN.n23 24.5923
R1891 VN.n26 VN.n23 24.5923
R1892 VN.n37 VN.n36 24.5923
R1893 VN.n36 VN.n21 24.5923
R1894 VN.n18 VN.n17 23.1168
R1895 VN.n38 VN.n37 23.1168
R1896 VN.n6 VN.n5 12.2964
R1897 VN.n26 VN.n25 12.2964
R1898 VN.n27 VN.n24 2.57552
R1899 VN.n7 VN.n4 2.57552
R1900 VN.n39 VN.n20 0.417304
R1901 VN.n19 VN.n0 0.417304
R1902 VN VN.n19 0.394524
R1903 VN.n35 VN.n20 0.189894
R1904 VN.n35 VN.n34 0.189894
R1905 VN.n34 VN.n33 0.189894
R1906 VN.n33 VN.n22 0.189894
R1907 VN.n29 VN.n22 0.189894
R1908 VN.n29 VN.n28 0.189894
R1909 VN.n28 VN.n27 0.189894
R1910 VN.n8 VN.n7 0.189894
R1911 VN.n9 VN.n8 0.189894
R1912 VN.n9 VN.n2 0.189894
R1913 VN.n13 VN.n2 0.189894
R1914 VN.n14 VN.n13 0.189894
R1915 VN.n15 VN.n14 0.189894
R1916 VN.n15 VN.n0 0.189894
R1917 VDD2.n135 VDD2.n71 289.615
R1918 VDD2.n64 VDD2.n0 289.615
R1919 VDD2.n136 VDD2.n135 185
R1920 VDD2.n134 VDD2.n133 185
R1921 VDD2.n75 VDD2.n74 185
R1922 VDD2.n128 VDD2.n127 185
R1923 VDD2.n126 VDD2.n125 185
R1924 VDD2.n79 VDD2.n78 185
R1925 VDD2.n120 VDD2.n119 185
R1926 VDD2.n118 VDD2.n117 185
R1927 VDD2.n116 VDD2.n82 185
R1928 VDD2.n86 VDD2.n83 185
R1929 VDD2.n111 VDD2.n110 185
R1930 VDD2.n109 VDD2.n108 185
R1931 VDD2.n88 VDD2.n87 185
R1932 VDD2.n103 VDD2.n102 185
R1933 VDD2.n101 VDD2.n100 185
R1934 VDD2.n92 VDD2.n91 185
R1935 VDD2.n95 VDD2.n94 185
R1936 VDD2.n23 VDD2.n22 185
R1937 VDD2.n20 VDD2.n19 185
R1938 VDD2.n29 VDD2.n28 185
R1939 VDD2.n31 VDD2.n30 185
R1940 VDD2.n16 VDD2.n15 185
R1941 VDD2.n37 VDD2.n36 185
R1942 VDD2.n40 VDD2.n39 185
R1943 VDD2.n38 VDD2.n12 185
R1944 VDD2.n45 VDD2.n11 185
R1945 VDD2.n47 VDD2.n46 185
R1946 VDD2.n49 VDD2.n48 185
R1947 VDD2.n8 VDD2.n7 185
R1948 VDD2.n55 VDD2.n54 185
R1949 VDD2.n57 VDD2.n56 185
R1950 VDD2.n4 VDD2.n3 185
R1951 VDD2.n63 VDD2.n62 185
R1952 VDD2.n65 VDD2.n64 185
R1953 VDD2.t4 VDD2.n93 149.524
R1954 VDD2.t3 VDD2.n21 149.524
R1955 VDD2.n135 VDD2.n134 104.615
R1956 VDD2.n134 VDD2.n74 104.615
R1957 VDD2.n127 VDD2.n74 104.615
R1958 VDD2.n127 VDD2.n126 104.615
R1959 VDD2.n126 VDD2.n78 104.615
R1960 VDD2.n119 VDD2.n78 104.615
R1961 VDD2.n119 VDD2.n118 104.615
R1962 VDD2.n118 VDD2.n82 104.615
R1963 VDD2.n86 VDD2.n82 104.615
R1964 VDD2.n110 VDD2.n86 104.615
R1965 VDD2.n110 VDD2.n109 104.615
R1966 VDD2.n109 VDD2.n87 104.615
R1967 VDD2.n102 VDD2.n87 104.615
R1968 VDD2.n102 VDD2.n101 104.615
R1969 VDD2.n101 VDD2.n91 104.615
R1970 VDD2.n94 VDD2.n91 104.615
R1971 VDD2.n22 VDD2.n19 104.615
R1972 VDD2.n29 VDD2.n19 104.615
R1973 VDD2.n30 VDD2.n29 104.615
R1974 VDD2.n30 VDD2.n15 104.615
R1975 VDD2.n37 VDD2.n15 104.615
R1976 VDD2.n39 VDD2.n37 104.615
R1977 VDD2.n39 VDD2.n38 104.615
R1978 VDD2.n38 VDD2.n11 104.615
R1979 VDD2.n47 VDD2.n11 104.615
R1980 VDD2.n48 VDD2.n47 104.615
R1981 VDD2.n48 VDD2.n7 104.615
R1982 VDD2.n55 VDD2.n7 104.615
R1983 VDD2.n56 VDD2.n55 104.615
R1984 VDD2.n56 VDD2.n3 104.615
R1985 VDD2.n63 VDD2.n3 104.615
R1986 VDD2.n64 VDD2.n63 104.615
R1987 VDD2.n70 VDD2.n69 61.0059
R1988 VDD2 VDD2.n141 61.0029
R1989 VDD2.n94 VDD2.t4 52.3082
R1990 VDD2.n22 VDD2.t3 52.3082
R1991 VDD2.n70 VDD2.n68 49.9857
R1992 VDD2.n140 VDD2.n139 47.3126
R1993 VDD2.n140 VDD2.n70 46.5386
R1994 VDD2.n117 VDD2.n116 13.1884
R1995 VDD2.n46 VDD2.n45 13.1884
R1996 VDD2.n120 VDD2.n81 12.8005
R1997 VDD2.n115 VDD2.n83 12.8005
R1998 VDD2.n44 VDD2.n12 12.8005
R1999 VDD2.n49 VDD2.n10 12.8005
R2000 VDD2.n121 VDD2.n79 12.0247
R2001 VDD2.n112 VDD2.n111 12.0247
R2002 VDD2.n41 VDD2.n40 12.0247
R2003 VDD2.n50 VDD2.n8 12.0247
R2004 VDD2.n125 VDD2.n124 11.249
R2005 VDD2.n108 VDD2.n85 11.249
R2006 VDD2.n36 VDD2.n14 11.249
R2007 VDD2.n54 VDD2.n53 11.249
R2008 VDD2.n128 VDD2.n77 10.4732
R2009 VDD2.n107 VDD2.n88 10.4732
R2010 VDD2.n35 VDD2.n16 10.4732
R2011 VDD2.n57 VDD2.n6 10.4732
R2012 VDD2.n95 VDD2.n93 10.2747
R2013 VDD2.n23 VDD2.n21 10.2747
R2014 VDD2.n129 VDD2.n75 9.69747
R2015 VDD2.n104 VDD2.n103 9.69747
R2016 VDD2.n32 VDD2.n31 9.69747
R2017 VDD2.n58 VDD2.n4 9.69747
R2018 VDD2.n139 VDD2.n138 9.45567
R2019 VDD2.n68 VDD2.n67 9.45567
R2020 VDD2.n97 VDD2.n96 9.3005
R2021 VDD2.n99 VDD2.n98 9.3005
R2022 VDD2.n90 VDD2.n89 9.3005
R2023 VDD2.n105 VDD2.n104 9.3005
R2024 VDD2.n107 VDD2.n106 9.3005
R2025 VDD2.n85 VDD2.n84 9.3005
R2026 VDD2.n113 VDD2.n112 9.3005
R2027 VDD2.n115 VDD2.n114 9.3005
R2028 VDD2.n138 VDD2.n137 9.3005
R2029 VDD2.n73 VDD2.n72 9.3005
R2030 VDD2.n132 VDD2.n131 9.3005
R2031 VDD2.n130 VDD2.n129 9.3005
R2032 VDD2.n77 VDD2.n76 9.3005
R2033 VDD2.n124 VDD2.n123 9.3005
R2034 VDD2.n122 VDD2.n121 9.3005
R2035 VDD2.n81 VDD2.n80 9.3005
R2036 VDD2.n2 VDD2.n1 9.3005
R2037 VDD2.n61 VDD2.n60 9.3005
R2038 VDD2.n59 VDD2.n58 9.3005
R2039 VDD2.n6 VDD2.n5 9.3005
R2040 VDD2.n53 VDD2.n52 9.3005
R2041 VDD2.n51 VDD2.n50 9.3005
R2042 VDD2.n10 VDD2.n9 9.3005
R2043 VDD2.n25 VDD2.n24 9.3005
R2044 VDD2.n27 VDD2.n26 9.3005
R2045 VDD2.n18 VDD2.n17 9.3005
R2046 VDD2.n33 VDD2.n32 9.3005
R2047 VDD2.n35 VDD2.n34 9.3005
R2048 VDD2.n14 VDD2.n13 9.3005
R2049 VDD2.n42 VDD2.n41 9.3005
R2050 VDD2.n44 VDD2.n43 9.3005
R2051 VDD2.n67 VDD2.n66 9.3005
R2052 VDD2.n133 VDD2.n132 8.92171
R2053 VDD2.n100 VDD2.n90 8.92171
R2054 VDD2.n28 VDD2.n18 8.92171
R2055 VDD2.n62 VDD2.n61 8.92171
R2056 VDD2.n136 VDD2.n73 8.14595
R2057 VDD2.n99 VDD2.n92 8.14595
R2058 VDD2.n27 VDD2.n20 8.14595
R2059 VDD2.n65 VDD2.n2 8.14595
R2060 VDD2.n137 VDD2.n71 7.3702
R2061 VDD2.n96 VDD2.n95 7.3702
R2062 VDD2.n24 VDD2.n23 7.3702
R2063 VDD2.n66 VDD2.n0 7.3702
R2064 VDD2.n139 VDD2.n71 6.59444
R2065 VDD2.n68 VDD2.n0 6.59444
R2066 VDD2.n137 VDD2.n136 5.81868
R2067 VDD2.n96 VDD2.n92 5.81868
R2068 VDD2.n24 VDD2.n20 5.81868
R2069 VDD2.n66 VDD2.n65 5.81868
R2070 VDD2.n133 VDD2.n73 5.04292
R2071 VDD2.n100 VDD2.n99 5.04292
R2072 VDD2.n28 VDD2.n27 5.04292
R2073 VDD2.n62 VDD2.n2 5.04292
R2074 VDD2.n132 VDD2.n75 4.26717
R2075 VDD2.n103 VDD2.n90 4.26717
R2076 VDD2.n31 VDD2.n18 4.26717
R2077 VDD2.n61 VDD2.n4 4.26717
R2078 VDD2.n129 VDD2.n128 3.49141
R2079 VDD2.n104 VDD2.n88 3.49141
R2080 VDD2.n32 VDD2.n16 3.49141
R2081 VDD2.n58 VDD2.n57 3.49141
R2082 VDD2.n97 VDD2.n93 2.84303
R2083 VDD2.n25 VDD2.n21 2.84303
R2084 VDD2 VDD2.n140 2.78714
R2085 VDD2.n125 VDD2.n77 2.71565
R2086 VDD2.n108 VDD2.n107 2.71565
R2087 VDD2.n36 VDD2.n35 2.71565
R2088 VDD2.n54 VDD2.n6 2.71565
R2089 VDD2.n124 VDD2.n79 1.93989
R2090 VDD2.n111 VDD2.n85 1.93989
R2091 VDD2.n40 VDD2.n14 1.93989
R2092 VDD2.n53 VDD2.n8 1.93989
R2093 VDD2.n141 VDD2.t1 1.55222
R2094 VDD2.n141 VDD2.t5 1.55222
R2095 VDD2.n69 VDD2.t0 1.55222
R2096 VDD2.n69 VDD2.t2 1.55222
R2097 VDD2.n121 VDD2.n120 1.16414
R2098 VDD2.n112 VDD2.n83 1.16414
R2099 VDD2.n41 VDD2.n12 1.16414
R2100 VDD2.n50 VDD2.n49 1.16414
R2101 VDD2.n117 VDD2.n81 0.388379
R2102 VDD2.n116 VDD2.n115 0.388379
R2103 VDD2.n45 VDD2.n44 0.388379
R2104 VDD2.n46 VDD2.n10 0.388379
R2105 VDD2.n138 VDD2.n72 0.155672
R2106 VDD2.n131 VDD2.n72 0.155672
R2107 VDD2.n131 VDD2.n130 0.155672
R2108 VDD2.n130 VDD2.n76 0.155672
R2109 VDD2.n123 VDD2.n76 0.155672
R2110 VDD2.n123 VDD2.n122 0.155672
R2111 VDD2.n122 VDD2.n80 0.155672
R2112 VDD2.n114 VDD2.n80 0.155672
R2113 VDD2.n114 VDD2.n113 0.155672
R2114 VDD2.n113 VDD2.n84 0.155672
R2115 VDD2.n106 VDD2.n84 0.155672
R2116 VDD2.n106 VDD2.n105 0.155672
R2117 VDD2.n105 VDD2.n89 0.155672
R2118 VDD2.n98 VDD2.n89 0.155672
R2119 VDD2.n98 VDD2.n97 0.155672
R2120 VDD2.n26 VDD2.n25 0.155672
R2121 VDD2.n26 VDD2.n17 0.155672
R2122 VDD2.n33 VDD2.n17 0.155672
R2123 VDD2.n34 VDD2.n33 0.155672
R2124 VDD2.n34 VDD2.n13 0.155672
R2125 VDD2.n42 VDD2.n13 0.155672
R2126 VDD2.n43 VDD2.n42 0.155672
R2127 VDD2.n43 VDD2.n9 0.155672
R2128 VDD2.n51 VDD2.n9 0.155672
R2129 VDD2.n52 VDD2.n51 0.155672
R2130 VDD2.n52 VDD2.n5 0.155672
R2131 VDD2.n59 VDD2.n5 0.155672
R2132 VDD2.n60 VDD2.n59 0.155672
R2133 VDD2.n60 VDD2.n1 0.155672
R2134 VDD2.n67 VDD2.n1 0.155672
R2135 VTAIL.n282 VTAIL.n218 289.615
R2136 VTAIL.n66 VTAIL.n2 289.615
R2137 VTAIL.n212 VTAIL.n148 289.615
R2138 VTAIL.n140 VTAIL.n76 289.615
R2139 VTAIL.n241 VTAIL.n240 185
R2140 VTAIL.n238 VTAIL.n237 185
R2141 VTAIL.n247 VTAIL.n246 185
R2142 VTAIL.n249 VTAIL.n248 185
R2143 VTAIL.n234 VTAIL.n233 185
R2144 VTAIL.n255 VTAIL.n254 185
R2145 VTAIL.n258 VTAIL.n257 185
R2146 VTAIL.n256 VTAIL.n230 185
R2147 VTAIL.n263 VTAIL.n229 185
R2148 VTAIL.n265 VTAIL.n264 185
R2149 VTAIL.n267 VTAIL.n266 185
R2150 VTAIL.n226 VTAIL.n225 185
R2151 VTAIL.n273 VTAIL.n272 185
R2152 VTAIL.n275 VTAIL.n274 185
R2153 VTAIL.n222 VTAIL.n221 185
R2154 VTAIL.n281 VTAIL.n280 185
R2155 VTAIL.n283 VTAIL.n282 185
R2156 VTAIL.n25 VTAIL.n24 185
R2157 VTAIL.n22 VTAIL.n21 185
R2158 VTAIL.n31 VTAIL.n30 185
R2159 VTAIL.n33 VTAIL.n32 185
R2160 VTAIL.n18 VTAIL.n17 185
R2161 VTAIL.n39 VTAIL.n38 185
R2162 VTAIL.n42 VTAIL.n41 185
R2163 VTAIL.n40 VTAIL.n14 185
R2164 VTAIL.n47 VTAIL.n13 185
R2165 VTAIL.n49 VTAIL.n48 185
R2166 VTAIL.n51 VTAIL.n50 185
R2167 VTAIL.n10 VTAIL.n9 185
R2168 VTAIL.n57 VTAIL.n56 185
R2169 VTAIL.n59 VTAIL.n58 185
R2170 VTAIL.n6 VTAIL.n5 185
R2171 VTAIL.n65 VTAIL.n64 185
R2172 VTAIL.n67 VTAIL.n66 185
R2173 VTAIL.n213 VTAIL.n212 185
R2174 VTAIL.n211 VTAIL.n210 185
R2175 VTAIL.n152 VTAIL.n151 185
R2176 VTAIL.n205 VTAIL.n204 185
R2177 VTAIL.n203 VTAIL.n202 185
R2178 VTAIL.n156 VTAIL.n155 185
R2179 VTAIL.n197 VTAIL.n196 185
R2180 VTAIL.n195 VTAIL.n194 185
R2181 VTAIL.n193 VTAIL.n159 185
R2182 VTAIL.n163 VTAIL.n160 185
R2183 VTAIL.n188 VTAIL.n187 185
R2184 VTAIL.n186 VTAIL.n185 185
R2185 VTAIL.n165 VTAIL.n164 185
R2186 VTAIL.n180 VTAIL.n179 185
R2187 VTAIL.n178 VTAIL.n177 185
R2188 VTAIL.n169 VTAIL.n168 185
R2189 VTAIL.n172 VTAIL.n171 185
R2190 VTAIL.n141 VTAIL.n140 185
R2191 VTAIL.n139 VTAIL.n138 185
R2192 VTAIL.n80 VTAIL.n79 185
R2193 VTAIL.n133 VTAIL.n132 185
R2194 VTAIL.n131 VTAIL.n130 185
R2195 VTAIL.n84 VTAIL.n83 185
R2196 VTAIL.n125 VTAIL.n124 185
R2197 VTAIL.n123 VTAIL.n122 185
R2198 VTAIL.n121 VTAIL.n87 185
R2199 VTAIL.n91 VTAIL.n88 185
R2200 VTAIL.n116 VTAIL.n115 185
R2201 VTAIL.n114 VTAIL.n113 185
R2202 VTAIL.n93 VTAIL.n92 185
R2203 VTAIL.n108 VTAIL.n107 185
R2204 VTAIL.n106 VTAIL.n105 185
R2205 VTAIL.n97 VTAIL.n96 185
R2206 VTAIL.n100 VTAIL.n99 185
R2207 VTAIL.t8 VTAIL.n239 149.524
R2208 VTAIL.t2 VTAIL.n23 149.524
R2209 VTAIL.t4 VTAIL.n170 149.524
R2210 VTAIL.t7 VTAIL.n98 149.524
R2211 VTAIL.n240 VTAIL.n237 104.615
R2212 VTAIL.n247 VTAIL.n237 104.615
R2213 VTAIL.n248 VTAIL.n247 104.615
R2214 VTAIL.n248 VTAIL.n233 104.615
R2215 VTAIL.n255 VTAIL.n233 104.615
R2216 VTAIL.n257 VTAIL.n255 104.615
R2217 VTAIL.n257 VTAIL.n256 104.615
R2218 VTAIL.n256 VTAIL.n229 104.615
R2219 VTAIL.n265 VTAIL.n229 104.615
R2220 VTAIL.n266 VTAIL.n265 104.615
R2221 VTAIL.n266 VTAIL.n225 104.615
R2222 VTAIL.n273 VTAIL.n225 104.615
R2223 VTAIL.n274 VTAIL.n273 104.615
R2224 VTAIL.n274 VTAIL.n221 104.615
R2225 VTAIL.n281 VTAIL.n221 104.615
R2226 VTAIL.n282 VTAIL.n281 104.615
R2227 VTAIL.n24 VTAIL.n21 104.615
R2228 VTAIL.n31 VTAIL.n21 104.615
R2229 VTAIL.n32 VTAIL.n31 104.615
R2230 VTAIL.n32 VTAIL.n17 104.615
R2231 VTAIL.n39 VTAIL.n17 104.615
R2232 VTAIL.n41 VTAIL.n39 104.615
R2233 VTAIL.n41 VTAIL.n40 104.615
R2234 VTAIL.n40 VTAIL.n13 104.615
R2235 VTAIL.n49 VTAIL.n13 104.615
R2236 VTAIL.n50 VTAIL.n49 104.615
R2237 VTAIL.n50 VTAIL.n9 104.615
R2238 VTAIL.n57 VTAIL.n9 104.615
R2239 VTAIL.n58 VTAIL.n57 104.615
R2240 VTAIL.n58 VTAIL.n5 104.615
R2241 VTAIL.n65 VTAIL.n5 104.615
R2242 VTAIL.n66 VTAIL.n65 104.615
R2243 VTAIL.n212 VTAIL.n211 104.615
R2244 VTAIL.n211 VTAIL.n151 104.615
R2245 VTAIL.n204 VTAIL.n151 104.615
R2246 VTAIL.n204 VTAIL.n203 104.615
R2247 VTAIL.n203 VTAIL.n155 104.615
R2248 VTAIL.n196 VTAIL.n155 104.615
R2249 VTAIL.n196 VTAIL.n195 104.615
R2250 VTAIL.n195 VTAIL.n159 104.615
R2251 VTAIL.n163 VTAIL.n159 104.615
R2252 VTAIL.n187 VTAIL.n163 104.615
R2253 VTAIL.n187 VTAIL.n186 104.615
R2254 VTAIL.n186 VTAIL.n164 104.615
R2255 VTAIL.n179 VTAIL.n164 104.615
R2256 VTAIL.n179 VTAIL.n178 104.615
R2257 VTAIL.n178 VTAIL.n168 104.615
R2258 VTAIL.n171 VTAIL.n168 104.615
R2259 VTAIL.n140 VTAIL.n139 104.615
R2260 VTAIL.n139 VTAIL.n79 104.615
R2261 VTAIL.n132 VTAIL.n79 104.615
R2262 VTAIL.n132 VTAIL.n131 104.615
R2263 VTAIL.n131 VTAIL.n83 104.615
R2264 VTAIL.n124 VTAIL.n83 104.615
R2265 VTAIL.n124 VTAIL.n123 104.615
R2266 VTAIL.n123 VTAIL.n87 104.615
R2267 VTAIL.n91 VTAIL.n87 104.615
R2268 VTAIL.n115 VTAIL.n91 104.615
R2269 VTAIL.n115 VTAIL.n114 104.615
R2270 VTAIL.n114 VTAIL.n92 104.615
R2271 VTAIL.n107 VTAIL.n92 104.615
R2272 VTAIL.n107 VTAIL.n106 104.615
R2273 VTAIL.n106 VTAIL.n96 104.615
R2274 VTAIL.n99 VTAIL.n96 104.615
R2275 VTAIL.n240 VTAIL.t8 52.3082
R2276 VTAIL.n24 VTAIL.t2 52.3082
R2277 VTAIL.n171 VTAIL.t4 52.3082
R2278 VTAIL.n99 VTAIL.t7 52.3082
R2279 VTAIL.n147 VTAIL.n146 43.473
R2280 VTAIL.n75 VTAIL.n74 43.473
R2281 VTAIL.n1 VTAIL.n0 43.473
R2282 VTAIL.n73 VTAIL.n72 43.473
R2283 VTAIL.n75 VTAIL.n73 30.6427
R2284 VTAIL.n287 VTAIL.n286 30.6338
R2285 VTAIL.n71 VTAIL.n70 30.6338
R2286 VTAIL.n217 VTAIL.n216 30.6338
R2287 VTAIL.n145 VTAIL.n144 30.6338
R2288 VTAIL.n287 VTAIL.n217 27.0048
R2289 VTAIL.n264 VTAIL.n263 13.1884
R2290 VTAIL.n48 VTAIL.n47 13.1884
R2291 VTAIL.n194 VTAIL.n193 13.1884
R2292 VTAIL.n122 VTAIL.n121 13.1884
R2293 VTAIL.n262 VTAIL.n230 12.8005
R2294 VTAIL.n267 VTAIL.n228 12.8005
R2295 VTAIL.n46 VTAIL.n14 12.8005
R2296 VTAIL.n51 VTAIL.n12 12.8005
R2297 VTAIL.n197 VTAIL.n158 12.8005
R2298 VTAIL.n192 VTAIL.n160 12.8005
R2299 VTAIL.n125 VTAIL.n86 12.8005
R2300 VTAIL.n120 VTAIL.n88 12.8005
R2301 VTAIL.n259 VTAIL.n258 12.0247
R2302 VTAIL.n268 VTAIL.n226 12.0247
R2303 VTAIL.n43 VTAIL.n42 12.0247
R2304 VTAIL.n52 VTAIL.n10 12.0247
R2305 VTAIL.n198 VTAIL.n156 12.0247
R2306 VTAIL.n189 VTAIL.n188 12.0247
R2307 VTAIL.n126 VTAIL.n84 12.0247
R2308 VTAIL.n117 VTAIL.n116 12.0247
R2309 VTAIL.n254 VTAIL.n232 11.249
R2310 VTAIL.n272 VTAIL.n271 11.249
R2311 VTAIL.n38 VTAIL.n16 11.249
R2312 VTAIL.n56 VTAIL.n55 11.249
R2313 VTAIL.n202 VTAIL.n201 11.249
R2314 VTAIL.n185 VTAIL.n162 11.249
R2315 VTAIL.n130 VTAIL.n129 11.249
R2316 VTAIL.n113 VTAIL.n90 11.249
R2317 VTAIL.n253 VTAIL.n234 10.4732
R2318 VTAIL.n275 VTAIL.n224 10.4732
R2319 VTAIL.n37 VTAIL.n18 10.4732
R2320 VTAIL.n59 VTAIL.n8 10.4732
R2321 VTAIL.n205 VTAIL.n154 10.4732
R2322 VTAIL.n184 VTAIL.n165 10.4732
R2323 VTAIL.n133 VTAIL.n82 10.4732
R2324 VTAIL.n112 VTAIL.n93 10.4732
R2325 VTAIL.n241 VTAIL.n239 10.2747
R2326 VTAIL.n25 VTAIL.n23 10.2747
R2327 VTAIL.n172 VTAIL.n170 10.2747
R2328 VTAIL.n100 VTAIL.n98 10.2747
R2329 VTAIL.n250 VTAIL.n249 9.69747
R2330 VTAIL.n276 VTAIL.n222 9.69747
R2331 VTAIL.n34 VTAIL.n33 9.69747
R2332 VTAIL.n60 VTAIL.n6 9.69747
R2333 VTAIL.n206 VTAIL.n152 9.69747
R2334 VTAIL.n181 VTAIL.n180 9.69747
R2335 VTAIL.n134 VTAIL.n80 9.69747
R2336 VTAIL.n109 VTAIL.n108 9.69747
R2337 VTAIL.n286 VTAIL.n285 9.45567
R2338 VTAIL.n70 VTAIL.n69 9.45567
R2339 VTAIL.n216 VTAIL.n215 9.45567
R2340 VTAIL.n144 VTAIL.n143 9.45567
R2341 VTAIL.n220 VTAIL.n219 9.3005
R2342 VTAIL.n279 VTAIL.n278 9.3005
R2343 VTAIL.n277 VTAIL.n276 9.3005
R2344 VTAIL.n224 VTAIL.n223 9.3005
R2345 VTAIL.n271 VTAIL.n270 9.3005
R2346 VTAIL.n269 VTAIL.n268 9.3005
R2347 VTAIL.n228 VTAIL.n227 9.3005
R2348 VTAIL.n243 VTAIL.n242 9.3005
R2349 VTAIL.n245 VTAIL.n244 9.3005
R2350 VTAIL.n236 VTAIL.n235 9.3005
R2351 VTAIL.n251 VTAIL.n250 9.3005
R2352 VTAIL.n253 VTAIL.n252 9.3005
R2353 VTAIL.n232 VTAIL.n231 9.3005
R2354 VTAIL.n260 VTAIL.n259 9.3005
R2355 VTAIL.n262 VTAIL.n261 9.3005
R2356 VTAIL.n285 VTAIL.n284 9.3005
R2357 VTAIL.n4 VTAIL.n3 9.3005
R2358 VTAIL.n63 VTAIL.n62 9.3005
R2359 VTAIL.n61 VTAIL.n60 9.3005
R2360 VTAIL.n8 VTAIL.n7 9.3005
R2361 VTAIL.n55 VTAIL.n54 9.3005
R2362 VTAIL.n53 VTAIL.n52 9.3005
R2363 VTAIL.n12 VTAIL.n11 9.3005
R2364 VTAIL.n27 VTAIL.n26 9.3005
R2365 VTAIL.n29 VTAIL.n28 9.3005
R2366 VTAIL.n20 VTAIL.n19 9.3005
R2367 VTAIL.n35 VTAIL.n34 9.3005
R2368 VTAIL.n37 VTAIL.n36 9.3005
R2369 VTAIL.n16 VTAIL.n15 9.3005
R2370 VTAIL.n44 VTAIL.n43 9.3005
R2371 VTAIL.n46 VTAIL.n45 9.3005
R2372 VTAIL.n69 VTAIL.n68 9.3005
R2373 VTAIL.n174 VTAIL.n173 9.3005
R2374 VTAIL.n176 VTAIL.n175 9.3005
R2375 VTAIL.n167 VTAIL.n166 9.3005
R2376 VTAIL.n182 VTAIL.n181 9.3005
R2377 VTAIL.n184 VTAIL.n183 9.3005
R2378 VTAIL.n162 VTAIL.n161 9.3005
R2379 VTAIL.n190 VTAIL.n189 9.3005
R2380 VTAIL.n192 VTAIL.n191 9.3005
R2381 VTAIL.n215 VTAIL.n214 9.3005
R2382 VTAIL.n150 VTAIL.n149 9.3005
R2383 VTAIL.n209 VTAIL.n208 9.3005
R2384 VTAIL.n207 VTAIL.n206 9.3005
R2385 VTAIL.n154 VTAIL.n153 9.3005
R2386 VTAIL.n201 VTAIL.n200 9.3005
R2387 VTAIL.n199 VTAIL.n198 9.3005
R2388 VTAIL.n158 VTAIL.n157 9.3005
R2389 VTAIL.n102 VTAIL.n101 9.3005
R2390 VTAIL.n104 VTAIL.n103 9.3005
R2391 VTAIL.n95 VTAIL.n94 9.3005
R2392 VTAIL.n110 VTAIL.n109 9.3005
R2393 VTAIL.n112 VTAIL.n111 9.3005
R2394 VTAIL.n90 VTAIL.n89 9.3005
R2395 VTAIL.n118 VTAIL.n117 9.3005
R2396 VTAIL.n120 VTAIL.n119 9.3005
R2397 VTAIL.n143 VTAIL.n142 9.3005
R2398 VTAIL.n78 VTAIL.n77 9.3005
R2399 VTAIL.n137 VTAIL.n136 9.3005
R2400 VTAIL.n135 VTAIL.n134 9.3005
R2401 VTAIL.n82 VTAIL.n81 9.3005
R2402 VTAIL.n129 VTAIL.n128 9.3005
R2403 VTAIL.n127 VTAIL.n126 9.3005
R2404 VTAIL.n86 VTAIL.n85 9.3005
R2405 VTAIL.n246 VTAIL.n236 8.92171
R2406 VTAIL.n280 VTAIL.n279 8.92171
R2407 VTAIL.n30 VTAIL.n20 8.92171
R2408 VTAIL.n64 VTAIL.n63 8.92171
R2409 VTAIL.n210 VTAIL.n209 8.92171
R2410 VTAIL.n177 VTAIL.n167 8.92171
R2411 VTAIL.n138 VTAIL.n137 8.92171
R2412 VTAIL.n105 VTAIL.n95 8.92171
R2413 VTAIL.n245 VTAIL.n238 8.14595
R2414 VTAIL.n283 VTAIL.n220 8.14595
R2415 VTAIL.n29 VTAIL.n22 8.14595
R2416 VTAIL.n67 VTAIL.n4 8.14595
R2417 VTAIL.n213 VTAIL.n150 8.14595
R2418 VTAIL.n176 VTAIL.n169 8.14595
R2419 VTAIL.n141 VTAIL.n78 8.14595
R2420 VTAIL.n104 VTAIL.n97 8.14595
R2421 VTAIL.n242 VTAIL.n241 7.3702
R2422 VTAIL.n284 VTAIL.n218 7.3702
R2423 VTAIL.n26 VTAIL.n25 7.3702
R2424 VTAIL.n68 VTAIL.n2 7.3702
R2425 VTAIL.n214 VTAIL.n148 7.3702
R2426 VTAIL.n173 VTAIL.n172 7.3702
R2427 VTAIL.n142 VTAIL.n76 7.3702
R2428 VTAIL.n101 VTAIL.n100 7.3702
R2429 VTAIL.n286 VTAIL.n218 6.59444
R2430 VTAIL.n70 VTAIL.n2 6.59444
R2431 VTAIL.n216 VTAIL.n148 6.59444
R2432 VTAIL.n144 VTAIL.n76 6.59444
R2433 VTAIL.n242 VTAIL.n238 5.81868
R2434 VTAIL.n284 VTAIL.n283 5.81868
R2435 VTAIL.n26 VTAIL.n22 5.81868
R2436 VTAIL.n68 VTAIL.n67 5.81868
R2437 VTAIL.n214 VTAIL.n213 5.81868
R2438 VTAIL.n173 VTAIL.n169 5.81868
R2439 VTAIL.n142 VTAIL.n141 5.81868
R2440 VTAIL.n101 VTAIL.n97 5.81868
R2441 VTAIL.n246 VTAIL.n245 5.04292
R2442 VTAIL.n280 VTAIL.n220 5.04292
R2443 VTAIL.n30 VTAIL.n29 5.04292
R2444 VTAIL.n64 VTAIL.n4 5.04292
R2445 VTAIL.n210 VTAIL.n150 5.04292
R2446 VTAIL.n177 VTAIL.n176 5.04292
R2447 VTAIL.n138 VTAIL.n78 5.04292
R2448 VTAIL.n105 VTAIL.n104 5.04292
R2449 VTAIL.n249 VTAIL.n236 4.26717
R2450 VTAIL.n279 VTAIL.n222 4.26717
R2451 VTAIL.n33 VTAIL.n20 4.26717
R2452 VTAIL.n63 VTAIL.n6 4.26717
R2453 VTAIL.n209 VTAIL.n152 4.26717
R2454 VTAIL.n180 VTAIL.n167 4.26717
R2455 VTAIL.n137 VTAIL.n80 4.26717
R2456 VTAIL.n108 VTAIL.n95 4.26717
R2457 VTAIL.n145 VTAIL.n75 3.63843
R2458 VTAIL.n217 VTAIL.n147 3.63843
R2459 VTAIL.n73 VTAIL.n71 3.63843
R2460 VTAIL.n250 VTAIL.n234 3.49141
R2461 VTAIL.n276 VTAIL.n275 3.49141
R2462 VTAIL.n34 VTAIL.n18 3.49141
R2463 VTAIL.n60 VTAIL.n59 3.49141
R2464 VTAIL.n206 VTAIL.n205 3.49141
R2465 VTAIL.n181 VTAIL.n165 3.49141
R2466 VTAIL.n134 VTAIL.n133 3.49141
R2467 VTAIL.n109 VTAIL.n93 3.49141
R2468 VTAIL.n243 VTAIL.n239 2.84303
R2469 VTAIL.n27 VTAIL.n23 2.84303
R2470 VTAIL.n174 VTAIL.n170 2.84303
R2471 VTAIL.n102 VTAIL.n98 2.84303
R2472 VTAIL.n254 VTAIL.n253 2.71565
R2473 VTAIL.n272 VTAIL.n224 2.71565
R2474 VTAIL.n38 VTAIL.n37 2.71565
R2475 VTAIL.n56 VTAIL.n8 2.71565
R2476 VTAIL.n202 VTAIL.n154 2.71565
R2477 VTAIL.n185 VTAIL.n184 2.71565
R2478 VTAIL.n130 VTAIL.n82 2.71565
R2479 VTAIL.n113 VTAIL.n112 2.71565
R2480 VTAIL VTAIL.n287 2.67076
R2481 VTAIL.n147 VTAIL.n145 2.28929
R2482 VTAIL.n71 VTAIL.n1 2.28929
R2483 VTAIL.n258 VTAIL.n232 1.93989
R2484 VTAIL.n271 VTAIL.n226 1.93989
R2485 VTAIL.n42 VTAIL.n16 1.93989
R2486 VTAIL.n55 VTAIL.n10 1.93989
R2487 VTAIL.n201 VTAIL.n156 1.93989
R2488 VTAIL.n188 VTAIL.n162 1.93989
R2489 VTAIL.n129 VTAIL.n84 1.93989
R2490 VTAIL.n116 VTAIL.n90 1.93989
R2491 VTAIL.n0 VTAIL.t10 1.55222
R2492 VTAIL.n0 VTAIL.t11 1.55222
R2493 VTAIL.n72 VTAIL.t3 1.55222
R2494 VTAIL.n72 VTAIL.t1 1.55222
R2495 VTAIL.n146 VTAIL.t0 1.55222
R2496 VTAIL.n146 VTAIL.t5 1.55222
R2497 VTAIL.n74 VTAIL.t9 1.55222
R2498 VTAIL.n74 VTAIL.t6 1.55222
R2499 VTAIL.n259 VTAIL.n230 1.16414
R2500 VTAIL.n268 VTAIL.n267 1.16414
R2501 VTAIL.n43 VTAIL.n14 1.16414
R2502 VTAIL.n52 VTAIL.n51 1.16414
R2503 VTAIL.n198 VTAIL.n197 1.16414
R2504 VTAIL.n189 VTAIL.n160 1.16414
R2505 VTAIL.n126 VTAIL.n125 1.16414
R2506 VTAIL.n117 VTAIL.n88 1.16414
R2507 VTAIL VTAIL.n1 0.968172
R2508 VTAIL.n263 VTAIL.n262 0.388379
R2509 VTAIL.n264 VTAIL.n228 0.388379
R2510 VTAIL.n47 VTAIL.n46 0.388379
R2511 VTAIL.n48 VTAIL.n12 0.388379
R2512 VTAIL.n194 VTAIL.n158 0.388379
R2513 VTAIL.n193 VTAIL.n192 0.388379
R2514 VTAIL.n122 VTAIL.n86 0.388379
R2515 VTAIL.n121 VTAIL.n120 0.388379
R2516 VTAIL.n244 VTAIL.n243 0.155672
R2517 VTAIL.n244 VTAIL.n235 0.155672
R2518 VTAIL.n251 VTAIL.n235 0.155672
R2519 VTAIL.n252 VTAIL.n251 0.155672
R2520 VTAIL.n252 VTAIL.n231 0.155672
R2521 VTAIL.n260 VTAIL.n231 0.155672
R2522 VTAIL.n261 VTAIL.n260 0.155672
R2523 VTAIL.n261 VTAIL.n227 0.155672
R2524 VTAIL.n269 VTAIL.n227 0.155672
R2525 VTAIL.n270 VTAIL.n269 0.155672
R2526 VTAIL.n270 VTAIL.n223 0.155672
R2527 VTAIL.n277 VTAIL.n223 0.155672
R2528 VTAIL.n278 VTAIL.n277 0.155672
R2529 VTAIL.n278 VTAIL.n219 0.155672
R2530 VTAIL.n285 VTAIL.n219 0.155672
R2531 VTAIL.n28 VTAIL.n27 0.155672
R2532 VTAIL.n28 VTAIL.n19 0.155672
R2533 VTAIL.n35 VTAIL.n19 0.155672
R2534 VTAIL.n36 VTAIL.n35 0.155672
R2535 VTAIL.n36 VTAIL.n15 0.155672
R2536 VTAIL.n44 VTAIL.n15 0.155672
R2537 VTAIL.n45 VTAIL.n44 0.155672
R2538 VTAIL.n45 VTAIL.n11 0.155672
R2539 VTAIL.n53 VTAIL.n11 0.155672
R2540 VTAIL.n54 VTAIL.n53 0.155672
R2541 VTAIL.n54 VTAIL.n7 0.155672
R2542 VTAIL.n61 VTAIL.n7 0.155672
R2543 VTAIL.n62 VTAIL.n61 0.155672
R2544 VTAIL.n62 VTAIL.n3 0.155672
R2545 VTAIL.n69 VTAIL.n3 0.155672
R2546 VTAIL.n215 VTAIL.n149 0.155672
R2547 VTAIL.n208 VTAIL.n149 0.155672
R2548 VTAIL.n208 VTAIL.n207 0.155672
R2549 VTAIL.n207 VTAIL.n153 0.155672
R2550 VTAIL.n200 VTAIL.n153 0.155672
R2551 VTAIL.n200 VTAIL.n199 0.155672
R2552 VTAIL.n199 VTAIL.n157 0.155672
R2553 VTAIL.n191 VTAIL.n157 0.155672
R2554 VTAIL.n191 VTAIL.n190 0.155672
R2555 VTAIL.n190 VTAIL.n161 0.155672
R2556 VTAIL.n183 VTAIL.n161 0.155672
R2557 VTAIL.n183 VTAIL.n182 0.155672
R2558 VTAIL.n182 VTAIL.n166 0.155672
R2559 VTAIL.n175 VTAIL.n166 0.155672
R2560 VTAIL.n175 VTAIL.n174 0.155672
R2561 VTAIL.n143 VTAIL.n77 0.155672
R2562 VTAIL.n136 VTAIL.n77 0.155672
R2563 VTAIL.n136 VTAIL.n135 0.155672
R2564 VTAIL.n135 VTAIL.n81 0.155672
R2565 VTAIL.n128 VTAIL.n81 0.155672
R2566 VTAIL.n128 VTAIL.n127 0.155672
R2567 VTAIL.n127 VTAIL.n85 0.155672
R2568 VTAIL.n119 VTAIL.n85 0.155672
R2569 VTAIL.n119 VTAIL.n118 0.155672
R2570 VTAIL.n118 VTAIL.n89 0.155672
R2571 VTAIL.n111 VTAIL.n89 0.155672
R2572 VTAIL.n111 VTAIL.n110 0.155672
R2573 VTAIL.n110 VTAIL.n94 0.155672
R2574 VTAIL.n103 VTAIL.n94 0.155672
R2575 VTAIL.n103 VTAIL.n102 0.155672
R2576 VP.n15 VP.n14 161.3
R2577 VP.n16 VP.n11 161.3
R2578 VP.n18 VP.n17 161.3
R2579 VP.n19 VP.n10 161.3
R2580 VP.n21 VP.n20 161.3
R2581 VP.n22 VP.n9 161.3
R2582 VP.n24 VP.n23 161.3
R2583 VP.n25 VP.n8 161.3
R2584 VP.n54 VP.n0 161.3
R2585 VP.n53 VP.n52 161.3
R2586 VP.n51 VP.n1 161.3
R2587 VP.n50 VP.n49 161.3
R2588 VP.n48 VP.n2 161.3
R2589 VP.n47 VP.n46 161.3
R2590 VP.n45 VP.n3 161.3
R2591 VP.n44 VP.n43 161.3
R2592 VP.n41 VP.n4 161.3
R2593 VP.n40 VP.n39 161.3
R2594 VP.n38 VP.n5 161.3
R2595 VP.n37 VP.n36 161.3
R2596 VP.n35 VP.n6 161.3
R2597 VP.n34 VP.n33 161.3
R2598 VP.n32 VP.n7 161.3
R2599 VP.n31 VP.n30 161.3
R2600 VP.n12 VP.t0 111.249
R2601 VP.n29 VP.t4 79.0535
R2602 VP.n42 VP.t3 79.0535
R2603 VP.n55 VP.t1 79.0535
R2604 VP.n26 VP.t5 79.0535
R2605 VP.n13 VP.t2 79.0535
R2606 VP.n13 VP.n12 63.0627
R2607 VP.n29 VP.n28 59.2636
R2608 VP.n56 VP.n55 59.2636
R2609 VP.n27 VP.n26 59.2636
R2610 VP.n28 VP.n27 54.5726
R2611 VP.n36 VP.n35 54.1398
R2612 VP.n49 VP.n48 54.1398
R2613 VP.n20 VP.n19 54.1398
R2614 VP.n35 VP.n34 27.0143
R2615 VP.n49 VP.n1 27.0143
R2616 VP.n20 VP.n9 27.0143
R2617 VP.n30 VP.n7 24.5923
R2618 VP.n34 VP.n7 24.5923
R2619 VP.n36 VP.n5 24.5923
R2620 VP.n40 VP.n5 24.5923
R2621 VP.n41 VP.n40 24.5923
R2622 VP.n43 VP.n3 24.5923
R2623 VP.n47 VP.n3 24.5923
R2624 VP.n48 VP.n47 24.5923
R2625 VP.n53 VP.n1 24.5923
R2626 VP.n54 VP.n53 24.5923
R2627 VP.n24 VP.n9 24.5923
R2628 VP.n25 VP.n24 24.5923
R2629 VP.n14 VP.n11 24.5923
R2630 VP.n18 VP.n11 24.5923
R2631 VP.n19 VP.n18 24.5923
R2632 VP.n30 VP.n29 23.1168
R2633 VP.n55 VP.n54 23.1168
R2634 VP.n26 VP.n25 23.1168
R2635 VP.n42 VP.n41 12.2964
R2636 VP.n43 VP.n42 12.2964
R2637 VP.n14 VP.n13 12.2964
R2638 VP.n15 VP.n12 2.57549
R2639 VP.n27 VP.n8 0.417304
R2640 VP.n31 VP.n28 0.417304
R2641 VP.n56 VP.n0 0.417304
R2642 VP VP.n56 0.394524
R2643 VP.n16 VP.n15 0.189894
R2644 VP.n17 VP.n16 0.189894
R2645 VP.n17 VP.n10 0.189894
R2646 VP.n21 VP.n10 0.189894
R2647 VP.n22 VP.n21 0.189894
R2648 VP.n23 VP.n22 0.189894
R2649 VP.n23 VP.n8 0.189894
R2650 VP.n32 VP.n31 0.189894
R2651 VP.n33 VP.n32 0.189894
R2652 VP.n33 VP.n6 0.189894
R2653 VP.n37 VP.n6 0.189894
R2654 VP.n38 VP.n37 0.189894
R2655 VP.n39 VP.n38 0.189894
R2656 VP.n39 VP.n4 0.189894
R2657 VP.n44 VP.n4 0.189894
R2658 VP.n45 VP.n44 0.189894
R2659 VP.n46 VP.n45 0.189894
R2660 VP.n46 VP.n2 0.189894
R2661 VP.n50 VP.n2 0.189894
R2662 VP.n51 VP.n50 0.189894
R2663 VP.n52 VP.n51 0.189894
R2664 VP.n52 VP.n0 0.189894
R2665 VDD1.n64 VDD1.n0 289.615
R2666 VDD1.n133 VDD1.n69 289.615
R2667 VDD1.n65 VDD1.n64 185
R2668 VDD1.n63 VDD1.n62 185
R2669 VDD1.n4 VDD1.n3 185
R2670 VDD1.n57 VDD1.n56 185
R2671 VDD1.n55 VDD1.n54 185
R2672 VDD1.n8 VDD1.n7 185
R2673 VDD1.n49 VDD1.n48 185
R2674 VDD1.n47 VDD1.n46 185
R2675 VDD1.n45 VDD1.n11 185
R2676 VDD1.n15 VDD1.n12 185
R2677 VDD1.n40 VDD1.n39 185
R2678 VDD1.n38 VDD1.n37 185
R2679 VDD1.n17 VDD1.n16 185
R2680 VDD1.n32 VDD1.n31 185
R2681 VDD1.n30 VDD1.n29 185
R2682 VDD1.n21 VDD1.n20 185
R2683 VDD1.n24 VDD1.n23 185
R2684 VDD1.n92 VDD1.n91 185
R2685 VDD1.n89 VDD1.n88 185
R2686 VDD1.n98 VDD1.n97 185
R2687 VDD1.n100 VDD1.n99 185
R2688 VDD1.n85 VDD1.n84 185
R2689 VDD1.n106 VDD1.n105 185
R2690 VDD1.n109 VDD1.n108 185
R2691 VDD1.n107 VDD1.n81 185
R2692 VDD1.n114 VDD1.n80 185
R2693 VDD1.n116 VDD1.n115 185
R2694 VDD1.n118 VDD1.n117 185
R2695 VDD1.n77 VDD1.n76 185
R2696 VDD1.n124 VDD1.n123 185
R2697 VDD1.n126 VDD1.n125 185
R2698 VDD1.n73 VDD1.n72 185
R2699 VDD1.n132 VDD1.n131 185
R2700 VDD1.n134 VDD1.n133 185
R2701 VDD1.t5 VDD1.n22 149.524
R2702 VDD1.t1 VDD1.n90 149.524
R2703 VDD1.n64 VDD1.n63 104.615
R2704 VDD1.n63 VDD1.n3 104.615
R2705 VDD1.n56 VDD1.n3 104.615
R2706 VDD1.n56 VDD1.n55 104.615
R2707 VDD1.n55 VDD1.n7 104.615
R2708 VDD1.n48 VDD1.n7 104.615
R2709 VDD1.n48 VDD1.n47 104.615
R2710 VDD1.n47 VDD1.n11 104.615
R2711 VDD1.n15 VDD1.n11 104.615
R2712 VDD1.n39 VDD1.n15 104.615
R2713 VDD1.n39 VDD1.n38 104.615
R2714 VDD1.n38 VDD1.n16 104.615
R2715 VDD1.n31 VDD1.n16 104.615
R2716 VDD1.n31 VDD1.n30 104.615
R2717 VDD1.n30 VDD1.n20 104.615
R2718 VDD1.n23 VDD1.n20 104.615
R2719 VDD1.n91 VDD1.n88 104.615
R2720 VDD1.n98 VDD1.n88 104.615
R2721 VDD1.n99 VDD1.n98 104.615
R2722 VDD1.n99 VDD1.n84 104.615
R2723 VDD1.n106 VDD1.n84 104.615
R2724 VDD1.n108 VDD1.n106 104.615
R2725 VDD1.n108 VDD1.n107 104.615
R2726 VDD1.n107 VDD1.n80 104.615
R2727 VDD1.n116 VDD1.n80 104.615
R2728 VDD1.n117 VDD1.n116 104.615
R2729 VDD1.n117 VDD1.n76 104.615
R2730 VDD1.n124 VDD1.n76 104.615
R2731 VDD1.n125 VDD1.n124 104.615
R2732 VDD1.n125 VDD1.n72 104.615
R2733 VDD1.n132 VDD1.n72 104.615
R2734 VDD1.n133 VDD1.n132 104.615
R2735 VDD1.n139 VDD1.n138 61.0059
R2736 VDD1.n141 VDD1.n140 60.1516
R2737 VDD1.n23 VDD1.t5 52.3082
R2738 VDD1.n91 VDD1.t1 52.3082
R2739 VDD1 VDD1.n68 50.0993
R2740 VDD1.n139 VDD1.n137 49.9857
R2741 VDD1.n141 VDD1.n139 48.9405
R2742 VDD1.n46 VDD1.n45 13.1884
R2743 VDD1.n115 VDD1.n114 13.1884
R2744 VDD1.n49 VDD1.n10 12.8005
R2745 VDD1.n44 VDD1.n12 12.8005
R2746 VDD1.n113 VDD1.n81 12.8005
R2747 VDD1.n118 VDD1.n79 12.8005
R2748 VDD1.n50 VDD1.n8 12.0247
R2749 VDD1.n41 VDD1.n40 12.0247
R2750 VDD1.n110 VDD1.n109 12.0247
R2751 VDD1.n119 VDD1.n77 12.0247
R2752 VDD1.n54 VDD1.n53 11.249
R2753 VDD1.n37 VDD1.n14 11.249
R2754 VDD1.n105 VDD1.n83 11.249
R2755 VDD1.n123 VDD1.n122 11.249
R2756 VDD1.n57 VDD1.n6 10.4732
R2757 VDD1.n36 VDD1.n17 10.4732
R2758 VDD1.n104 VDD1.n85 10.4732
R2759 VDD1.n126 VDD1.n75 10.4732
R2760 VDD1.n24 VDD1.n22 10.2747
R2761 VDD1.n92 VDD1.n90 10.2747
R2762 VDD1.n58 VDD1.n4 9.69747
R2763 VDD1.n33 VDD1.n32 9.69747
R2764 VDD1.n101 VDD1.n100 9.69747
R2765 VDD1.n127 VDD1.n73 9.69747
R2766 VDD1.n68 VDD1.n67 9.45567
R2767 VDD1.n137 VDD1.n136 9.45567
R2768 VDD1.n26 VDD1.n25 9.3005
R2769 VDD1.n28 VDD1.n27 9.3005
R2770 VDD1.n19 VDD1.n18 9.3005
R2771 VDD1.n34 VDD1.n33 9.3005
R2772 VDD1.n36 VDD1.n35 9.3005
R2773 VDD1.n14 VDD1.n13 9.3005
R2774 VDD1.n42 VDD1.n41 9.3005
R2775 VDD1.n44 VDD1.n43 9.3005
R2776 VDD1.n67 VDD1.n66 9.3005
R2777 VDD1.n2 VDD1.n1 9.3005
R2778 VDD1.n61 VDD1.n60 9.3005
R2779 VDD1.n59 VDD1.n58 9.3005
R2780 VDD1.n6 VDD1.n5 9.3005
R2781 VDD1.n53 VDD1.n52 9.3005
R2782 VDD1.n51 VDD1.n50 9.3005
R2783 VDD1.n10 VDD1.n9 9.3005
R2784 VDD1.n71 VDD1.n70 9.3005
R2785 VDD1.n130 VDD1.n129 9.3005
R2786 VDD1.n128 VDD1.n127 9.3005
R2787 VDD1.n75 VDD1.n74 9.3005
R2788 VDD1.n122 VDD1.n121 9.3005
R2789 VDD1.n120 VDD1.n119 9.3005
R2790 VDD1.n79 VDD1.n78 9.3005
R2791 VDD1.n94 VDD1.n93 9.3005
R2792 VDD1.n96 VDD1.n95 9.3005
R2793 VDD1.n87 VDD1.n86 9.3005
R2794 VDD1.n102 VDD1.n101 9.3005
R2795 VDD1.n104 VDD1.n103 9.3005
R2796 VDD1.n83 VDD1.n82 9.3005
R2797 VDD1.n111 VDD1.n110 9.3005
R2798 VDD1.n113 VDD1.n112 9.3005
R2799 VDD1.n136 VDD1.n135 9.3005
R2800 VDD1.n62 VDD1.n61 8.92171
R2801 VDD1.n29 VDD1.n19 8.92171
R2802 VDD1.n97 VDD1.n87 8.92171
R2803 VDD1.n131 VDD1.n130 8.92171
R2804 VDD1.n65 VDD1.n2 8.14595
R2805 VDD1.n28 VDD1.n21 8.14595
R2806 VDD1.n96 VDD1.n89 8.14595
R2807 VDD1.n134 VDD1.n71 8.14595
R2808 VDD1.n66 VDD1.n0 7.3702
R2809 VDD1.n25 VDD1.n24 7.3702
R2810 VDD1.n93 VDD1.n92 7.3702
R2811 VDD1.n135 VDD1.n69 7.3702
R2812 VDD1.n68 VDD1.n0 6.59444
R2813 VDD1.n137 VDD1.n69 6.59444
R2814 VDD1.n66 VDD1.n65 5.81868
R2815 VDD1.n25 VDD1.n21 5.81868
R2816 VDD1.n93 VDD1.n89 5.81868
R2817 VDD1.n135 VDD1.n134 5.81868
R2818 VDD1.n62 VDD1.n2 5.04292
R2819 VDD1.n29 VDD1.n28 5.04292
R2820 VDD1.n97 VDD1.n96 5.04292
R2821 VDD1.n131 VDD1.n71 5.04292
R2822 VDD1.n61 VDD1.n4 4.26717
R2823 VDD1.n32 VDD1.n19 4.26717
R2824 VDD1.n100 VDD1.n87 4.26717
R2825 VDD1.n130 VDD1.n73 4.26717
R2826 VDD1.n58 VDD1.n57 3.49141
R2827 VDD1.n33 VDD1.n17 3.49141
R2828 VDD1.n101 VDD1.n85 3.49141
R2829 VDD1.n127 VDD1.n126 3.49141
R2830 VDD1.n26 VDD1.n22 2.84303
R2831 VDD1.n94 VDD1.n90 2.84303
R2832 VDD1.n54 VDD1.n6 2.71565
R2833 VDD1.n37 VDD1.n36 2.71565
R2834 VDD1.n105 VDD1.n104 2.71565
R2835 VDD1.n123 VDD1.n75 2.71565
R2836 VDD1.n53 VDD1.n8 1.93989
R2837 VDD1.n40 VDD1.n14 1.93989
R2838 VDD1.n109 VDD1.n83 1.93989
R2839 VDD1.n122 VDD1.n77 1.93989
R2840 VDD1.n140 VDD1.t3 1.55222
R2841 VDD1.n140 VDD1.t0 1.55222
R2842 VDD1.n138 VDD1.t2 1.55222
R2843 VDD1.n138 VDD1.t4 1.55222
R2844 VDD1.n50 VDD1.n49 1.16414
R2845 VDD1.n41 VDD1.n12 1.16414
R2846 VDD1.n110 VDD1.n81 1.16414
R2847 VDD1.n119 VDD1.n118 1.16414
R2848 VDD1 VDD1.n141 0.851793
R2849 VDD1.n46 VDD1.n10 0.388379
R2850 VDD1.n45 VDD1.n44 0.388379
R2851 VDD1.n114 VDD1.n113 0.388379
R2852 VDD1.n115 VDD1.n79 0.388379
R2853 VDD1.n67 VDD1.n1 0.155672
R2854 VDD1.n60 VDD1.n1 0.155672
R2855 VDD1.n60 VDD1.n59 0.155672
R2856 VDD1.n59 VDD1.n5 0.155672
R2857 VDD1.n52 VDD1.n5 0.155672
R2858 VDD1.n52 VDD1.n51 0.155672
R2859 VDD1.n51 VDD1.n9 0.155672
R2860 VDD1.n43 VDD1.n9 0.155672
R2861 VDD1.n43 VDD1.n42 0.155672
R2862 VDD1.n42 VDD1.n13 0.155672
R2863 VDD1.n35 VDD1.n13 0.155672
R2864 VDD1.n35 VDD1.n34 0.155672
R2865 VDD1.n34 VDD1.n18 0.155672
R2866 VDD1.n27 VDD1.n18 0.155672
R2867 VDD1.n27 VDD1.n26 0.155672
R2868 VDD1.n95 VDD1.n94 0.155672
R2869 VDD1.n95 VDD1.n86 0.155672
R2870 VDD1.n102 VDD1.n86 0.155672
R2871 VDD1.n103 VDD1.n102 0.155672
R2872 VDD1.n103 VDD1.n82 0.155672
R2873 VDD1.n111 VDD1.n82 0.155672
R2874 VDD1.n112 VDD1.n111 0.155672
R2875 VDD1.n112 VDD1.n78 0.155672
R2876 VDD1.n120 VDD1.n78 0.155672
R2877 VDD1.n121 VDD1.n120 0.155672
R2878 VDD1.n121 VDD1.n74 0.155672
R2879 VDD1.n128 VDD1.n74 0.155672
R2880 VDD1.n129 VDD1.n128 0.155672
R2881 VDD1.n129 VDD1.n70 0.155672
R2882 VDD1.n136 VDD1.n70 0.155672
C0 VP VN 8.31715f
C1 VTAIL VDD2 8.50806f
C2 VP VDD2 0.567436f
C3 VN VDD2 7.59675f
C4 VTAIL VDD1 8.44768f
C5 VP VDD1 8.00888f
C6 VN VDD1 0.152883f
C7 VP VTAIL 8.045461f
C8 VN VTAIL 8.03052f
C9 VDD1 VDD2 1.91082f
C10 VDD2 B 7.111055f
C11 VDD1 B 7.295453f
C12 VTAIL B 8.938512f
C13 VN B 16.75733f
C14 VP B 15.480748f
C15 VDD1.n0 B 0.029777f
C16 VDD1.n1 B 0.021599f
C17 VDD1.n2 B 0.011607f
C18 VDD1.n3 B 0.027434f
C19 VDD1.n4 B 0.012289f
C20 VDD1.n5 B 0.021599f
C21 VDD1.n6 B 0.011607f
C22 VDD1.n7 B 0.027434f
C23 VDD1.n8 B 0.012289f
C24 VDD1.n9 B 0.021599f
C25 VDD1.n10 B 0.011607f
C26 VDD1.n11 B 0.027434f
C27 VDD1.n12 B 0.012289f
C28 VDD1.n13 B 0.021599f
C29 VDD1.n14 B 0.011607f
C30 VDD1.n15 B 0.027434f
C31 VDD1.n16 B 0.027434f
C32 VDD1.n17 B 0.012289f
C33 VDD1.n18 B 0.021599f
C34 VDD1.n19 B 0.011607f
C35 VDD1.n20 B 0.027434f
C36 VDD1.n21 B 0.012289f
C37 VDD1.n22 B 0.162032f
C38 VDD1.t5 B 0.046422f
C39 VDD1.n23 B 0.020575f
C40 VDD1.n24 B 0.019394f
C41 VDD1.n25 B 0.011607f
C42 VDD1.n26 B 1.16267f
C43 VDD1.n27 B 0.021599f
C44 VDD1.n28 B 0.011607f
C45 VDD1.n29 B 0.012289f
C46 VDD1.n30 B 0.027434f
C47 VDD1.n31 B 0.027434f
C48 VDD1.n32 B 0.012289f
C49 VDD1.n33 B 0.011607f
C50 VDD1.n34 B 0.021599f
C51 VDD1.n35 B 0.021599f
C52 VDD1.n36 B 0.011607f
C53 VDD1.n37 B 0.012289f
C54 VDD1.n38 B 0.027434f
C55 VDD1.n39 B 0.027434f
C56 VDD1.n40 B 0.012289f
C57 VDD1.n41 B 0.011607f
C58 VDD1.n42 B 0.021599f
C59 VDD1.n43 B 0.021599f
C60 VDD1.n44 B 0.011607f
C61 VDD1.n45 B 0.011948f
C62 VDD1.n46 B 0.011948f
C63 VDD1.n47 B 0.027434f
C64 VDD1.n48 B 0.027434f
C65 VDD1.n49 B 0.012289f
C66 VDD1.n50 B 0.011607f
C67 VDD1.n51 B 0.021599f
C68 VDD1.n52 B 0.021599f
C69 VDD1.n53 B 0.011607f
C70 VDD1.n54 B 0.012289f
C71 VDD1.n55 B 0.027434f
C72 VDD1.n56 B 0.027434f
C73 VDD1.n57 B 0.012289f
C74 VDD1.n58 B 0.011607f
C75 VDD1.n59 B 0.021599f
C76 VDD1.n60 B 0.021599f
C77 VDD1.n61 B 0.011607f
C78 VDD1.n62 B 0.012289f
C79 VDD1.n63 B 0.027434f
C80 VDD1.n64 B 0.058359f
C81 VDD1.n65 B 0.012289f
C82 VDD1.n66 B 0.011607f
C83 VDD1.n67 B 0.047565f
C84 VDD1.n68 B 0.060434f
C85 VDD1.n69 B 0.029777f
C86 VDD1.n70 B 0.021599f
C87 VDD1.n71 B 0.011607f
C88 VDD1.n72 B 0.027434f
C89 VDD1.n73 B 0.012289f
C90 VDD1.n74 B 0.021599f
C91 VDD1.n75 B 0.011607f
C92 VDD1.n76 B 0.027434f
C93 VDD1.n77 B 0.012289f
C94 VDD1.n78 B 0.021599f
C95 VDD1.n79 B 0.011607f
C96 VDD1.n80 B 0.027434f
C97 VDD1.n81 B 0.012289f
C98 VDD1.n82 B 0.021599f
C99 VDD1.n83 B 0.011607f
C100 VDD1.n84 B 0.027434f
C101 VDD1.n85 B 0.012289f
C102 VDD1.n86 B 0.021599f
C103 VDD1.n87 B 0.011607f
C104 VDD1.n88 B 0.027434f
C105 VDD1.n89 B 0.012289f
C106 VDD1.n90 B 0.162032f
C107 VDD1.t1 B 0.046422f
C108 VDD1.n91 B 0.020575f
C109 VDD1.n92 B 0.019394f
C110 VDD1.n93 B 0.011607f
C111 VDD1.n94 B 1.16267f
C112 VDD1.n95 B 0.021599f
C113 VDD1.n96 B 0.011607f
C114 VDD1.n97 B 0.012289f
C115 VDD1.n98 B 0.027434f
C116 VDD1.n99 B 0.027434f
C117 VDD1.n100 B 0.012289f
C118 VDD1.n101 B 0.011607f
C119 VDD1.n102 B 0.021599f
C120 VDD1.n103 B 0.021599f
C121 VDD1.n104 B 0.011607f
C122 VDD1.n105 B 0.012289f
C123 VDD1.n106 B 0.027434f
C124 VDD1.n107 B 0.027434f
C125 VDD1.n108 B 0.027434f
C126 VDD1.n109 B 0.012289f
C127 VDD1.n110 B 0.011607f
C128 VDD1.n111 B 0.021599f
C129 VDD1.n112 B 0.021599f
C130 VDD1.n113 B 0.011607f
C131 VDD1.n114 B 0.011948f
C132 VDD1.n115 B 0.011948f
C133 VDD1.n116 B 0.027434f
C134 VDD1.n117 B 0.027434f
C135 VDD1.n118 B 0.012289f
C136 VDD1.n119 B 0.011607f
C137 VDD1.n120 B 0.021599f
C138 VDD1.n121 B 0.021599f
C139 VDD1.n122 B 0.011607f
C140 VDD1.n123 B 0.012289f
C141 VDD1.n124 B 0.027434f
C142 VDD1.n125 B 0.027434f
C143 VDD1.n126 B 0.012289f
C144 VDD1.n127 B 0.011607f
C145 VDD1.n128 B 0.021599f
C146 VDD1.n129 B 0.021599f
C147 VDD1.n130 B 0.011607f
C148 VDD1.n131 B 0.012289f
C149 VDD1.n132 B 0.027434f
C150 VDD1.n133 B 0.058359f
C151 VDD1.n134 B 0.012289f
C152 VDD1.n135 B 0.011607f
C153 VDD1.n136 B 0.047565f
C154 VDD1.n137 B 0.059519f
C155 VDD1.t2 B 0.217794f
C156 VDD1.t4 B 0.217794f
C157 VDD1.n138 B 1.95294f
C158 VDD1.n139 B 2.9739f
C159 VDD1.t3 B 0.217794f
C160 VDD1.t0 B 0.217794f
C161 VDD1.n140 B 1.94589f
C162 VDD1.n141 B 2.7771f
C163 VP.n0 B 0.033904f
C164 VP.t1 B 2.44251f
C165 VP.n1 B 0.034766f
C166 VP.n2 B 0.01803f
C167 VP.n3 B 0.033435f
C168 VP.n4 B 0.01803f
C169 VP.t3 B 2.44251f
C170 VP.n5 B 0.033435f
C171 VP.n6 B 0.01803f
C172 VP.n7 B 0.033435f
C173 VP.n8 B 0.033904f
C174 VP.t5 B 2.44251f
C175 VP.n9 B 0.034766f
C176 VP.n10 B 0.01803f
C177 VP.n11 B 0.033435f
C178 VP.t0 B 2.73045f
C179 VP.n12 B 0.874566f
C180 VP.t2 B 2.44251f
C181 VP.n13 B 0.917374f
C182 VP.n14 B 0.025182f
C183 VP.n15 B 0.236103f
C184 VP.n16 B 0.01803f
C185 VP.n17 B 0.01803f
C186 VP.n18 B 0.033435f
C187 VP.n19 B 0.031453f
C188 VP.n20 B 0.019634f
C189 VP.n21 B 0.01803f
C190 VP.n22 B 0.01803f
C191 VP.n23 B 0.01803f
C192 VP.n24 B 0.033435f
C193 VP.n25 B 0.032444f
C194 VP.n26 B 0.933401f
C195 VP.n27 B 1.18126f
C196 VP.n28 B 1.19317f
C197 VP.t4 B 2.44251f
C198 VP.n29 B 0.933401f
C199 VP.n30 B 0.032444f
C200 VP.n31 B 0.033904f
C201 VP.n32 B 0.01803f
C202 VP.n33 B 0.01803f
C203 VP.n34 B 0.034766f
C204 VP.n35 B 0.019634f
C205 VP.n36 B 0.031453f
C206 VP.n37 B 0.01803f
C207 VP.n38 B 0.01803f
C208 VP.n39 B 0.01803f
C209 VP.n40 B 0.033435f
C210 VP.n41 B 0.025182f
C211 VP.n42 B 0.852515f
C212 VP.n43 B 0.025182f
C213 VP.n44 B 0.01803f
C214 VP.n45 B 0.01803f
C215 VP.n46 B 0.01803f
C216 VP.n47 B 0.033435f
C217 VP.n48 B 0.031453f
C218 VP.n49 B 0.019634f
C219 VP.n50 B 0.01803f
C220 VP.n51 B 0.01803f
C221 VP.n52 B 0.01803f
C222 VP.n53 B 0.033435f
C223 VP.n54 B 0.032444f
C224 VP.n55 B 0.933401f
C225 VP.n56 B 0.053897f
C226 VTAIL.t10 B 0.24439f
C227 VTAIL.t11 B 0.24439f
C228 VTAIL.n0 B 2.10719f
C229 VTAIL.n1 B 0.501269f
C230 VTAIL.n2 B 0.033413f
C231 VTAIL.n3 B 0.024237f
C232 VTAIL.n4 B 0.013024f
C233 VTAIL.n5 B 0.030784f
C234 VTAIL.n6 B 0.01379f
C235 VTAIL.n7 B 0.024237f
C236 VTAIL.n8 B 0.013024f
C237 VTAIL.n9 B 0.030784f
C238 VTAIL.n10 B 0.01379f
C239 VTAIL.n11 B 0.024237f
C240 VTAIL.n12 B 0.013024f
C241 VTAIL.n13 B 0.030784f
C242 VTAIL.n14 B 0.01379f
C243 VTAIL.n15 B 0.024237f
C244 VTAIL.n16 B 0.013024f
C245 VTAIL.n17 B 0.030784f
C246 VTAIL.n18 B 0.01379f
C247 VTAIL.n19 B 0.024237f
C248 VTAIL.n20 B 0.013024f
C249 VTAIL.n21 B 0.030784f
C250 VTAIL.n22 B 0.01379f
C251 VTAIL.n23 B 0.181817f
C252 VTAIL.t2 B 0.052091f
C253 VTAIL.n24 B 0.023088f
C254 VTAIL.n25 B 0.021762f
C255 VTAIL.n26 B 0.013024f
C256 VTAIL.n27 B 1.30464f
C257 VTAIL.n28 B 0.024237f
C258 VTAIL.n29 B 0.013024f
C259 VTAIL.n30 B 0.01379f
C260 VTAIL.n31 B 0.030784f
C261 VTAIL.n32 B 0.030784f
C262 VTAIL.n33 B 0.01379f
C263 VTAIL.n34 B 0.013024f
C264 VTAIL.n35 B 0.024237f
C265 VTAIL.n36 B 0.024237f
C266 VTAIL.n37 B 0.013024f
C267 VTAIL.n38 B 0.01379f
C268 VTAIL.n39 B 0.030784f
C269 VTAIL.n40 B 0.030784f
C270 VTAIL.n41 B 0.030784f
C271 VTAIL.n42 B 0.01379f
C272 VTAIL.n43 B 0.013024f
C273 VTAIL.n44 B 0.024237f
C274 VTAIL.n45 B 0.024237f
C275 VTAIL.n46 B 0.013024f
C276 VTAIL.n47 B 0.013407f
C277 VTAIL.n48 B 0.013407f
C278 VTAIL.n49 B 0.030784f
C279 VTAIL.n50 B 0.030784f
C280 VTAIL.n51 B 0.01379f
C281 VTAIL.n52 B 0.013024f
C282 VTAIL.n53 B 0.024237f
C283 VTAIL.n54 B 0.024237f
C284 VTAIL.n55 B 0.013024f
C285 VTAIL.n56 B 0.01379f
C286 VTAIL.n57 B 0.030784f
C287 VTAIL.n58 B 0.030784f
C288 VTAIL.n59 B 0.01379f
C289 VTAIL.n60 B 0.013024f
C290 VTAIL.n61 B 0.024237f
C291 VTAIL.n62 B 0.024237f
C292 VTAIL.n63 B 0.013024f
C293 VTAIL.n64 B 0.01379f
C294 VTAIL.n65 B 0.030784f
C295 VTAIL.n66 B 0.065485f
C296 VTAIL.n67 B 0.01379f
C297 VTAIL.n68 B 0.013024f
C298 VTAIL.n69 B 0.053374f
C299 VTAIL.n70 B 0.036439f
C300 VTAIL.n71 B 0.482066f
C301 VTAIL.t3 B 0.24439f
C302 VTAIL.t1 B 0.24439f
C303 VTAIL.n72 B 2.10719f
C304 VTAIL.n73 B 2.28758f
C305 VTAIL.t9 B 0.24439f
C306 VTAIL.t6 B 0.24439f
C307 VTAIL.n74 B 2.10719f
C308 VTAIL.n75 B 2.28758f
C309 VTAIL.n76 B 0.033413f
C310 VTAIL.n77 B 0.024237f
C311 VTAIL.n78 B 0.013024f
C312 VTAIL.n79 B 0.030784f
C313 VTAIL.n80 B 0.01379f
C314 VTAIL.n81 B 0.024237f
C315 VTAIL.n82 B 0.013024f
C316 VTAIL.n83 B 0.030784f
C317 VTAIL.n84 B 0.01379f
C318 VTAIL.n85 B 0.024237f
C319 VTAIL.n86 B 0.013024f
C320 VTAIL.n87 B 0.030784f
C321 VTAIL.n88 B 0.01379f
C322 VTAIL.n89 B 0.024237f
C323 VTAIL.n90 B 0.013024f
C324 VTAIL.n91 B 0.030784f
C325 VTAIL.n92 B 0.030784f
C326 VTAIL.n93 B 0.01379f
C327 VTAIL.n94 B 0.024237f
C328 VTAIL.n95 B 0.013024f
C329 VTAIL.n96 B 0.030784f
C330 VTAIL.n97 B 0.01379f
C331 VTAIL.n98 B 0.181817f
C332 VTAIL.t7 B 0.052091f
C333 VTAIL.n99 B 0.023088f
C334 VTAIL.n100 B 0.021762f
C335 VTAIL.n101 B 0.013024f
C336 VTAIL.n102 B 1.30464f
C337 VTAIL.n103 B 0.024237f
C338 VTAIL.n104 B 0.013024f
C339 VTAIL.n105 B 0.01379f
C340 VTAIL.n106 B 0.030784f
C341 VTAIL.n107 B 0.030784f
C342 VTAIL.n108 B 0.01379f
C343 VTAIL.n109 B 0.013024f
C344 VTAIL.n110 B 0.024237f
C345 VTAIL.n111 B 0.024237f
C346 VTAIL.n112 B 0.013024f
C347 VTAIL.n113 B 0.01379f
C348 VTAIL.n114 B 0.030784f
C349 VTAIL.n115 B 0.030784f
C350 VTAIL.n116 B 0.01379f
C351 VTAIL.n117 B 0.013024f
C352 VTAIL.n118 B 0.024237f
C353 VTAIL.n119 B 0.024237f
C354 VTAIL.n120 B 0.013024f
C355 VTAIL.n121 B 0.013407f
C356 VTAIL.n122 B 0.013407f
C357 VTAIL.n123 B 0.030784f
C358 VTAIL.n124 B 0.030784f
C359 VTAIL.n125 B 0.01379f
C360 VTAIL.n126 B 0.013024f
C361 VTAIL.n127 B 0.024237f
C362 VTAIL.n128 B 0.024237f
C363 VTAIL.n129 B 0.013024f
C364 VTAIL.n130 B 0.01379f
C365 VTAIL.n131 B 0.030784f
C366 VTAIL.n132 B 0.030784f
C367 VTAIL.n133 B 0.01379f
C368 VTAIL.n134 B 0.013024f
C369 VTAIL.n135 B 0.024237f
C370 VTAIL.n136 B 0.024237f
C371 VTAIL.n137 B 0.013024f
C372 VTAIL.n138 B 0.01379f
C373 VTAIL.n139 B 0.030784f
C374 VTAIL.n140 B 0.065485f
C375 VTAIL.n141 B 0.01379f
C376 VTAIL.n142 B 0.013024f
C377 VTAIL.n143 B 0.053374f
C378 VTAIL.n144 B 0.036439f
C379 VTAIL.n145 B 0.482066f
C380 VTAIL.t0 B 0.24439f
C381 VTAIL.t5 B 0.24439f
C382 VTAIL.n146 B 2.10719f
C383 VTAIL.n147 B 0.709805f
C384 VTAIL.n148 B 0.033413f
C385 VTAIL.n149 B 0.024237f
C386 VTAIL.n150 B 0.013024f
C387 VTAIL.n151 B 0.030784f
C388 VTAIL.n152 B 0.01379f
C389 VTAIL.n153 B 0.024237f
C390 VTAIL.n154 B 0.013024f
C391 VTAIL.n155 B 0.030784f
C392 VTAIL.n156 B 0.01379f
C393 VTAIL.n157 B 0.024237f
C394 VTAIL.n158 B 0.013024f
C395 VTAIL.n159 B 0.030784f
C396 VTAIL.n160 B 0.01379f
C397 VTAIL.n161 B 0.024237f
C398 VTAIL.n162 B 0.013024f
C399 VTAIL.n163 B 0.030784f
C400 VTAIL.n164 B 0.030784f
C401 VTAIL.n165 B 0.01379f
C402 VTAIL.n166 B 0.024237f
C403 VTAIL.n167 B 0.013024f
C404 VTAIL.n168 B 0.030784f
C405 VTAIL.n169 B 0.01379f
C406 VTAIL.n170 B 0.181817f
C407 VTAIL.t4 B 0.052091f
C408 VTAIL.n171 B 0.023088f
C409 VTAIL.n172 B 0.021762f
C410 VTAIL.n173 B 0.013024f
C411 VTAIL.n174 B 1.30464f
C412 VTAIL.n175 B 0.024237f
C413 VTAIL.n176 B 0.013024f
C414 VTAIL.n177 B 0.01379f
C415 VTAIL.n178 B 0.030784f
C416 VTAIL.n179 B 0.030784f
C417 VTAIL.n180 B 0.01379f
C418 VTAIL.n181 B 0.013024f
C419 VTAIL.n182 B 0.024237f
C420 VTAIL.n183 B 0.024237f
C421 VTAIL.n184 B 0.013024f
C422 VTAIL.n185 B 0.01379f
C423 VTAIL.n186 B 0.030784f
C424 VTAIL.n187 B 0.030784f
C425 VTAIL.n188 B 0.01379f
C426 VTAIL.n189 B 0.013024f
C427 VTAIL.n190 B 0.024237f
C428 VTAIL.n191 B 0.024237f
C429 VTAIL.n192 B 0.013024f
C430 VTAIL.n193 B 0.013407f
C431 VTAIL.n194 B 0.013407f
C432 VTAIL.n195 B 0.030784f
C433 VTAIL.n196 B 0.030784f
C434 VTAIL.n197 B 0.01379f
C435 VTAIL.n198 B 0.013024f
C436 VTAIL.n199 B 0.024237f
C437 VTAIL.n200 B 0.024237f
C438 VTAIL.n201 B 0.013024f
C439 VTAIL.n202 B 0.01379f
C440 VTAIL.n203 B 0.030784f
C441 VTAIL.n204 B 0.030784f
C442 VTAIL.n205 B 0.01379f
C443 VTAIL.n206 B 0.013024f
C444 VTAIL.n207 B 0.024237f
C445 VTAIL.n208 B 0.024237f
C446 VTAIL.n209 B 0.013024f
C447 VTAIL.n210 B 0.01379f
C448 VTAIL.n211 B 0.030784f
C449 VTAIL.n212 B 0.065485f
C450 VTAIL.n213 B 0.01379f
C451 VTAIL.n214 B 0.013024f
C452 VTAIL.n215 B 0.053374f
C453 VTAIL.n216 B 0.036439f
C454 VTAIL.n217 B 1.77573f
C455 VTAIL.n218 B 0.033413f
C456 VTAIL.n219 B 0.024237f
C457 VTAIL.n220 B 0.013024f
C458 VTAIL.n221 B 0.030784f
C459 VTAIL.n222 B 0.01379f
C460 VTAIL.n223 B 0.024237f
C461 VTAIL.n224 B 0.013024f
C462 VTAIL.n225 B 0.030784f
C463 VTAIL.n226 B 0.01379f
C464 VTAIL.n227 B 0.024237f
C465 VTAIL.n228 B 0.013024f
C466 VTAIL.n229 B 0.030784f
C467 VTAIL.n230 B 0.01379f
C468 VTAIL.n231 B 0.024237f
C469 VTAIL.n232 B 0.013024f
C470 VTAIL.n233 B 0.030784f
C471 VTAIL.n234 B 0.01379f
C472 VTAIL.n235 B 0.024237f
C473 VTAIL.n236 B 0.013024f
C474 VTAIL.n237 B 0.030784f
C475 VTAIL.n238 B 0.01379f
C476 VTAIL.n239 B 0.181817f
C477 VTAIL.t8 B 0.052091f
C478 VTAIL.n240 B 0.023088f
C479 VTAIL.n241 B 0.021762f
C480 VTAIL.n242 B 0.013024f
C481 VTAIL.n243 B 1.30464f
C482 VTAIL.n244 B 0.024237f
C483 VTAIL.n245 B 0.013024f
C484 VTAIL.n246 B 0.01379f
C485 VTAIL.n247 B 0.030784f
C486 VTAIL.n248 B 0.030784f
C487 VTAIL.n249 B 0.01379f
C488 VTAIL.n250 B 0.013024f
C489 VTAIL.n251 B 0.024237f
C490 VTAIL.n252 B 0.024237f
C491 VTAIL.n253 B 0.013024f
C492 VTAIL.n254 B 0.01379f
C493 VTAIL.n255 B 0.030784f
C494 VTAIL.n256 B 0.030784f
C495 VTAIL.n257 B 0.030784f
C496 VTAIL.n258 B 0.01379f
C497 VTAIL.n259 B 0.013024f
C498 VTAIL.n260 B 0.024237f
C499 VTAIL.n261 B 0.024237f
C500 VTAIL.n262 B 0.013024f
C501 VTAIL.n263 B 0.013407f
C502 VTAIL.n264 B 0.013407f
C503 VTAIL.n265 B 0.030784f
C504 VTAIL.n266 B 0.030784f
C505 VTAIL.n267 B 0.01379f
C506 VTAIL.n268 B 0.013024f
C507 VTAIL.n269 B 0.024237f
C508 VTAIL.n270 B 0.024237f
C509 VTAIL.n271 B 0.013024f
C510 VTAIL.n272 B 0.01379f
C511 VTAIL.n273 B 0.030784f
C512 VTAIL.n274 B 0.030784f
C513 VTAIL.n275 B 0.01379f
C514 VTAIL.n276 B 0.013024f
C515 VTAIL.n277 B 0.024237f
C516 VTAIL.n278 B 0.024237f
C517 VTAIL.n279 B 0.013024f
C518 VTAIL.n280 B 0.01379f
C519 VTAIL.n281 B 0.030784f
C520 VTAIL.n282 B 0.065485f
C521 VTAIL.n283 B 0.01379f
C522 VTAIL.n284 B 0.013024f
C523 VTAIL.n285 B 0.053374f
C524 VTAIL.n286 B 0.036439f
C525 VTAIL.n287 B 1.70016f
C526 VDD2.n0 B 0.029375f
C527 VDD2.n1 B 0.021308f
C528 VDD2.n2 B 0.01145f
C529 VDD2.n3 B 0.027064f
C530 VDD2.n4 B 0.012123f
C531 VDD2.n5 B 0.021308f
C532 VDD2.n6 B 0.01145f
C533 VDD2.n7 B 0.027064f
C534 VDD2.n8 B 0.012123f
C535 VDD2.n9 B 0.021308f
C536 VDD2.n10 B 0.01145f
C537 VDD2.n11 B 0.027064f
C538 VDD2.n12 B 0.012123f
C539 VDD2.n13 B 0.021308f
C540 VDD2.n14 B 0.01145f
C541 VDD2.n15 B 0.027064f
C542 VDD2.n16 B 0.012123f
C543 VDD2.n17 B 0.021308f
C544 VDD2.n18 B 0.01145f
C545 VDD2.n19 B 0.027064f
C546 VDD2.n20 B 0.012123f
C547 VDD2.n21 B 0.159845f
C548 VDD2.t3 B 0.045796f
C549 VDD2.n22 B 0.020298f
C550 VDD2.n23 B 0.019132f
C551 VDD2.n24 B 0.01145f
C552 VDD2.n25 B 1.14698f
C553 VDD2.n26 B 0.021308f
C554 VDD2.n27 B 0.01145f
C555 VDD2.n28 B 0.012123f
C556 VDD2.n29 B 0.027064f
C557 VDD2.n30 B 0.027064f
C558 VDD2.n31 B 0.012123f
C559 VDD2.n32 B 0.01145f
C560 VDD2.n33 B 0.021308f
C561 VDD2.n34 B 0.021308f
C562 VDD2.n35 B 0.01145f
C563 VDD2.n36 B 0.012123f
C564 VDD2.n37 B 0.027064f
C565 VDD2.n38 B 0.027064f
C566 VDD2.n39 B 0.027064f
C567 VDD2.n40 B 0.012123f
C568 VDD2.n41 B 0.01145f
C569 VDD2.n42 B 0.021308f
C570 VDD2.n43 B 0.021308f
C571 VDD2.n44 B 0.01145f
C572 VDD2.n45 B 0.011787f
C573 VDD2.n46 B 0.011787f
C574 VDD2.n47 B 0.027064f
C575 VDD2.n48 B 0.027064f
C576 VDD2.n49 B 0.012123f
C577 VDD2.n50 B 0.01145f
C578 VDD2.n51 B 0.021308f
C579 VDD2.n52 B 0.021308f
C580 VDD2.n53 B 0.01145f
C581 VDD2.n54 B 0.012123f
C582 VDD2.n55 B 0.027064f
C583 VDD2.n56 B 0.027064f
C584 VDD2.n57 B 0.012123f
C585 VDD2.n58 B 0.01145f
C586 VDD2.n59 B 0.021308f
C587 VDD2.n60 B 0.021308f
C588 VDD2.n61 B 0.01145f
C589 VDD2.n62 B 0.012123f
C590 VDD2.n63 B 0.027064f
C591 VDD2.n64 B 0.057571f
C592 VDD2.n65 B 0.012123f
C593 VDD2.n66 B 0.01145f
C594 VDD2.n67 B 0.046924f
C595 VDD2.n68 B 0.058716f
C596 VDD2.t0 B 0.214856f
C597 VDD2.t2 B 0.214856f
C598 VDD2.n69 B 1.92659f
C599 VDD2.n70 B 2.79794f
C600 VDD2.n71 B 0.029375f
C601 VDD2.n72 B 0.021308f
C602 VDD2.n73 B 0.01145f
C603 VDD2.n74 B 0.027064f
C604 VDD2.n75 B 0.012123f
C605 VDD2.n76 B 0.021308f
C606 VDD2.n77 B 0.01145f
C607 VDD2.n78 B 0.027064f
C608 VDD2.n79 B 0.012123f
C609 VDD2.n80 B 0.021308f
C610 VDD2.n81 B 0.01145f
C611 VDD2.n82 B 0.027064f
C612 VDD2.n83 B 0.012123f
C613 VDD2.n84 B 0.021308f
C614 VDD2.n85 B 0.01145f
C615 VDD2.n86 B 0.027064f
C616 VDD2.n87 B 0.027064f
C617 VDD2.n88 B 0.012123f
C618 VDD2.n89 B 0.021308f
C619 VDD2.n90 B 0.01145f
C620 VDD2.n91 B 0.027064f
C621 VDD2.n92 B 0.012123f
C622 VDD2.n93 B 0.159845f
C623 VDD2.t4 B 0.045796f
C624 VDD2.n94 B 0.020298f
C625 VDD2.n95 B 0.019132f
C626 VDD2.n96 B 0.01145f
C627 VDD2.n97 B 1.14698f
C628 VDD2.n98 B 0.021308f
C629 VDD2.n99 B 0.01145f
C630 VDD2.n100 B 0.012123f
C631 VDD2.n101 B 0.027064f
C632 VDD2.n102 B 0.027064f
C633 VDD2.n103 B 0.012123f
C634 VDD2.n104 B 0.01145f
C635 VDD2.n105 B 0.021308f
C636 VDD2.n106 B 0.021308f
C637 VDD2.n107 B 0.01145f
C638 VDD2.n108 B 0.012123f
C639 VDD2.n109 B 0.027064f
C640 VDD2.n110 B 0.027064f
C641 VDD2.n111 B 0.012123f
C642 VDD2.n112 B 0.01145f
C643 VDD2.n113 B 0.021308f
C644 VDD2.n114 B 0.021308f
C645 VDD2.n115 B 0.01145f
C646 VDD2.n116 B 0.011787f
C647 VDD2.n117 B 0.011787f
C648 VDD2.n118 B 0.027064f
C649 VDD2.n119 B 0.027064f
C650 VDD2.n120 B 0.012123f
C651 VDD2.n121 B 0.01145f
C652 VDD2.n122 B 0.021308f
C653 VDD2.n123 B 0.021308f
C654 VDD2.n124 B 0.01145f
C655 VDD2.n125 B 0.012123f
C656 VDD2.n126 B 0.027064f
C657 VDD2.n127 B 0.027064f
C658 VDD2.n128 B 0.012123f
C659 VDD2.n129 B 0.01145f
C660 VDD2.n130 B 0.021308f
C661 VDD2.n131 B 0.021308f
C662 VDD2.n132 B 0.01145f
C663 VDD2.n133 B 0.012123f
C664 VDD2.n134 B 0.027064f
C665 VDD2.n135 B 0.057571f
C666 VDD2.n136 B 0.012123f
C667 VDD2.n137 B 0.01145f
C668 VDD2.n138 B 0.046924f
C669 VDD2.n139 B 0.046768f
C670 VDD2.n140 B 2.532f
C671 VDD2.t1 B 0.214856f
C672 VDD2.t5 B 0.214856f
C673 VDD2.n141 B 1.92655f
C674 VN.n0 B 0.033311f
C675 VN.t3 B 2.3998f
C676 VN.n1 B 0.034159f
C677 VN.n2 B 0.017715f
C678 VN.n3 B 0.03285f
C679 VN.t1 B 2.68271f
C680 VN.n4 B 0.859271f
C681 VN.t0 B 2.3998f
C682 VN.n5 B 0.901333f
C683 VN.n6 B 0.024741f
C684 VN.n7 B 0.231974f
C685 VN.n8 B 0.017715f
C686 VN.n9 B 0.017715f
C687 VN.n10 B 0.03285f
C688 VN.n11 B 0.030903f
C689 VN.n12 B 0.01929f
C690 VN.n13 B 0.017715f
C691 VN.n14 B 0.017715f
C692 VN.n15 B 0.017715f
C693 VN.n16 B 0.03285f
C694 VN.n17 B 0.031877f
C695 VN.n18 B 0.91708f
C696 VN.n19 B 0.052954f
C697 VN.n20 B 0.033311f
C698 VN.t2 B 2.3998f
C699 VN.n21 B 0.034159f
C700 VN.n22 B 0.017715f
C701 VN.n23 B 0.03285f
C702 VN.t4 B 2.68271f
C703 VN.n24 B 0.859271f
C704 VN.t5 B 2.3998f
C705 VN.n25 B 0.901333f
C706 VN.n26 B 0.024741f
C707 VN.n27 B 0.231974f
C708 VN.n28 B 0.017715f
C709 VN.n29 B 0.017715f
C710 VN.n30 B 0.03285f
C711 VN.n31 B 0.030903f
C712 VN.n32 B 0.01929f
C713 VN.n33 B 0.017715f
C714 VN.n34 B 0.017715f
C715 VN.n35 B 0.017715f
C716 VN.n36 B 0.03285f
C717 VN.n37 B 0.031877f
C718 VN.n38 B 0.91708f
C719 VN.n39 B 1.16494f
.ends

