* NGSPICE file created from diff_pair_sample_1302.ext - technology: sky130A

.subckt diff_pair_sample_1302 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t7 w_n1550_n3126# sky130_fd_pr__pfet_01v8 ad=4.2081 pd=22.36 as=1.78035 ps=11.12 w=10.79 l=0.25
X1 B.t11 B.t9 B.t10 w_n1550_n3126# sky130_fd_pr__pfet_01v8 ad=4.2081 pd=22.36 as=0 ps=0 w=10.79 l=0.25
X2 VDD2.t7 VN.t0 VTAIL.t1 w_n1550_n3126# sky130_fd_pr__pfet_01v8 ad=1.78035 pd=11.12 as=1.78035 ps=11.12 w=10.79 l=0.25
X3 B.t8 B.t6 B.t7 w_n1550_n3126# sky130_fd_pr__pfet_01v8 ad=4.2081 pd=22.36 as=0 ps=0 w=10.79 l=0.25
X4 B.t5 B.t3 B.t4 w_n1550_n3126# sky130_fd_pr__pfet_01v8 ad=4.2081 pd=22.36 as=0 ps=0 w=10.79 l=0.25
X5 VTAIL.t14 VP.t1 VDD1.t3 w_n1550_n3126# sky130_fd_pr__pfet_01v8 ad=1.78035 pd=11.12 as=1.78035 ps=11.12 w=10.79 l=0.25
X6 VDD1.t2 VP.t2 VTAIL.t13 w_n1550_n3126# sky130_fd_pr__pfet_01v8 ad=1.78035 pd=11.12 as=1.78035 ps=11.12 w=10.79 l=0.25
X7 VDD2.t6 VN.t1 VTAIL.t3 w_n1550_n3126# sky130_fd_pr__pfet_01v8 ad=1.78035 pd=11.12 as=4.2081 ps=22.36 w=10.79 l=0.25
X8 VDD2.t5 VN.t2 VTAIL.t4 w_n1550_n3126# sky130_fd_pr__pfet_01v8 ad=1.78035 pd=11.12 as=1.78035 ps=11.12 w=10.79 l=0.25
X9 VDD2.t4 VN.t3 VTAIL.t5 w_n1550_n3126# sky130_fd_pr__pfet_01v8 ad=1.78035 pd=11.12 as=4.2081 ps=22.36 w=10.79 l=0.25
X10 VTAIL.t12 VP.t3 VDD1.t4 w_n1550_n3126# sky130_fd_pr__pfet_01v8 ad=1.78035 pd=11.12 as=1.78035 ps=11.12 w=10.79 l=0.25
X11 VTAIL.t6 VN.t4 VDD2.t3 w_n1550_n3126# sky130_fd_pr__pfet_01v8 ad=1.78035 pd=11.12 as=1.78035 ps=11.12 w=10.79 l=0.25
X12 VDD1.t0 VP.t4 VTAIL.t11 w_n1550_n3126# sky130_fd_pr__pfet_01v8 ad=1.78035 pd=11.12 as=4.2081 ps=22.36 w=10.79 l=0.25
X13 B.t2 B.t0 B.t1 w_n1550_n3126# sky130_fd_pr__pfet_01v8 ad=4.2081 pd=22.36 as=0 ps=0 w=10.79 l=0.25
X14 VDD1.t1 VP.t5 VTAIL.t10 w_n1550_n3126# sky130_fd_pr__pfet_01v8 ad=1.78035 pd=11.12 as=1.78035 ps=11.12 w=10.79 l=0.25
X15 VDD1.t6 VP.t6 VTAIL.t9 w_n1550_n3126# sky130_fd_pr__pfet_01v8 ad=1.78035 pd=11.12 as=4.2081 ps=22.36 w=10.79 l=0.25
X16 VTAIL.t0 VN.t5 VDD2.t2 w_n1550_n3126# sky130_fd_pr__pfet_01v8 ad=4.2081 pd=22.36 as=1.78035 ps=11.12 w=10.79 l=0.25
X17 VTAIL.t7 VN.t6 VDD2.t1 w_n1550_n3126# sky130_fd_pr__pfet_01v8 ad=4.2081 pd=22.36 as=1.78035 ps=11.12 w=10.79 l=0.25
X18 VTAIL.t2 VN.t7 VDD2.t0 w_n1550_n3126# sky130_fd_pr__pfet_01v8 ad=1.78035 pd=11.12 as=1.78035 ps=11.12 w=10.79 l=0.25
X19 VTAIL.t8 VP.t7 VDD1.t5 w_n1550_n3126# sky130_fd_pr__pfet_01v8 ad=4.2081 pd=22.36 as=1.78035 ps=11.12 w=10.79 l=0.25
R0 VP.n13 VP.t6 1220.48
R1 VP.n9 VP.t7 1220.48
R2 VP.n2 VP.t0 1220.48
R3 VP.n6 VP.t4 1220.48
R4 VP.n12 VP.t3 1166.44
R5 VP.n10 VP.t2 1166.44
R6 VP.n3 VP.t5 1166.44
R7 VP.n5 VP.t1 1166.44
R8 VP.n2 VP.n1 161.489
R9 VP.n14 VP.n13 161.3
R10 VP.n4 VP.n1 161.3
R11 VP.n7 VP.n6 161.3
R12 VP.n11 VP.n0 161.3
R13 VP.n9 VP.n8 161.3
R14 VP.n11 VP.n10 42.3581
R15 VP.n12 VP.n11 42.3581
R16 VP.n4 VP.n3 42.3581
R17 VP.n5 VP.n4 42.3581
R18 VP.n8 VP.n7 39.1066
R19 VP.n10 VP.n9 30.6732
R20 VP.n13 VP.n12 30.6732
R21 VP.n3 VP.n2 30.6732
R22 VP.n6 VP.n5 30.6732
R23 VP.n7 VP.n1 0.189894
R24 VP.n8 VP.n0 0.189894
R25 VP.n14 VP.n0 0.189894
R26 VP VP.n14 0.0516364
R27 VDD1 VDD1.n0 78.3077
R28 VDD1.n3 VDD1.n2 78.194
R29 VDD1.n3 VDD1.n1 78.194
R30 VDD1.n5 VDD1.n4 77.9993
R31 VDD1.n5 VDD1.n3 35.85
R32 VDD1.n4 VDD1.t3 3.01301
R33 VDD1.n4 VDD1.t0 3.01301
R34 VDD1.n0 VDD1.t7 3.01301
R35 VDD1.n0 VDD1.t1 3.01301
R36 VDD1.n2 VDD1.t4 3.01301
R37 VDD1.n2 VDD1.t6 3.01301
R38 VDD1.n1 VDD1.t5 3.01301
R39 VDD1.n1 VDD1.t2 3.01301
R40 VDD1 VDD1.n5 0.19231
R41 VTAIL.n466 VTAIL.n414 756.745
R42 VTAIL.n54 VTAIL.n2 756.745
R43 VTAIL.n112 VTAIL.n60 756.745
R44 VTAIL.n172 VTAIL.n120 756.745
R45 VTAIL.n408 VTAIL.n356 756.745
R46 VTAIL.n348 VTAIL.n296 756.745
R47 VTAIL.n290 VTAIL.n238 756.745
R48 VTAIL.n230 VTAIL.n178 756.745
R49 VTAIL.n433 VTAIL.n432 585
R50 VTAIL.n430 VTAIL.n429 585
R51 VTAIL.n439 VTAIL.n438 585
R52 VTAIL.n441 VTAIL.n440 585
R53 VTAIL.n426 VTAIL.n425 585
R54 VTAIL.n447 VTAIL.n446 585
R55 VTAIL.n450 VTAIL.n449 585
R56 VTAIL.n448 VTAIL.n422 585
R57 VTAIL.n455 VTAIL.n421 585
R58 VTAIL.n457 VTAIL.n456 585
R59 VTAIL.n459 VTAIL.n458 585
R60 VTAIL.n418 VTAIL.n417 585
R61 VTAIL.n465 VTAIL.n464 585
R62 VTAIL.n467 VTAIL.n466 585
R63 VTAIL.n21 VTAIL.n20 585
R64 VTAIL.n18 VTAIL.n17 585
R65 VTAIL.n27 VTAIL.n26 585
R66 VTAIL.n29 VTAIL.n28 585
R67 VTAIL.n14 VTAIL.n13 585
R68 VTAIL.n35 VTAIL.n34 585
R69 VTAIL.n38 VTAIL.n37 585
R70 VTAIL.n36 VTAIL.n10 585
R71 VTAIL.n43 VTAIL.n9 585
R72 VTAIL.n45 VTAIL.n44 585
R73 VTAIL.n47 VTAIL.n46 585
R74 VTAIL.n6 VTAIL.n5 585
R75 VTAIL.n53 VTAIL.n52 585
R76 VTAIL.n55 VTAIL.n54 585
R77 VTAIL.n79 VTAIL.n78 585
R78 VTAIL.n76 VTAIL.n75 585
R79 VTAIL.n85 VTAIL.n84 585
R80 VTAIL.n87 VTAIL.n86 585
R81 VTAIL.n72 VTAIL.n71 585
R82 VTAIL.n93 VTAIL.n92 585
R83 VTAIL.n96 VTAIL.n95 585
R84 VTAIL.n94 VTAIL.n68 585
R85 VTAIL.n101 VTAIL.n67 585
R86 VTAIL.n103 VTAIL.n102 585
R87 VTAIL.n105 VTAIL.n104 585
R88 VTAIL.n64 VTAIL.n63 585
R89 VTAIL.n111 VTAIL.n110 585
R90 VTAIL.n113 VTAIL.n112 585
R91 VTAIL.n139 VTAIL.n138 585
R92 VTAIL.n136 VTAIL.n135 585
R93 VTAIL.n145 VTAIL.n144 585
R94 VTAIL.n147 VTAIL.n146 585
R95 VTAIL.n132 VTAIL.n131 585
R96 VTAIL.n153 VTAIL.n152 585
R97 VTAIL.n156 VTAIL.n155 585
R98 VTAIL.n154 VTAIL.n128 585
R99 VTAIL.n161 VTAIL.n127 585
R100 VTAIL.n163 VTAIL.n162 585
R101 VTAIL.n165 VTAIL.n164 585
R102 VTAIL.n124 VTAIL.n123 585
R103 VTAIL.n171 VTAIL.n170 585
R104 VTAIL.n173 VTAIL.n172 585
R105 VTAIL.n409 VTAIL.n408 585
R106 VTAIL.n407 VTAIL.n406 585
R107 VTAIL.n360 VTAIL.n359 585
R108 VTAIL.n401 VTAIL.n400 585
R109 VTAIL.n399 VTAIL.n398 585
R110 VTAIL.n397 VTAIL.n363 585
R111 VTAIL.n367 VTAIL.n364 585
R112 VTAIL.n392 VTAIL.n391 585
R113 VTAIL.n390 VTAIL.n389 585
R114 VTAIL.n369 VTAIL.n368 585
R115 VTAIL.n384 VTAIL.n383 585
R116 VTAIL.n382 VTAIL.n381 585
R117 VTAIL.n373 VTAIL.n372 585
R118 VTAIL.n376 VTAIL.n375 585
R119 VTAIL.n349 VTAIL.n348 585
R120 VTAIL.n347 VTAIL.n346 585
R121 VTAIL.n300 VTAIL.n299 585
R122 VTAIL.n341 VTAIL.n340 585
R123 VTAIL.n339 VTAIL.n338 585
R124 VTAIL.n337 VTAIL.n303 585
R125 VTAIL.n307 VTAIL.n304 585
R126 VTAIL.n332 VTAIL.n331 585
R127 VTAIL.n330 VTAIL.n329 585
R128 VTAIL.n309 VTAIL.n308 585
R129 VTAIL.n324 VTAIL.n323 585
R130 VTAIL.n322 VTAIL.n321 585
R131 VTAIL.n313 VTAIL.n312 585
R132 VTAIL.n316 VTAIL.n315 585
R133 VTAIL.n291 VTAIL.n290 585
R134 VTAIL.n289 VTAIL.n288 585
R135 VTAIL.n242 VTAIL.n241 585
R136 VTAIL.n283 VTAIL.n282 585
R137 VTAIL.n281 VTAIL.n280 585
R138 VTAIL.n279 VTAIL.n245 585
R139 VTAIL.n249 VTAIL.n246 585
R140 VTAIL.n274 VTAIL.n273 585
R141 VTAIL.n272 VTAIL.n271 585
R142 VTAIL.n251 VTAIL.n250 585
R143 VTAIL.n266 VTAIL.n265 585
R144 VTAIL.n264 VTAIL.n263 585
R145 VTAIL.n255 VTAIL.n254 585
R146 VTAIL.n258 VTAIL.n257 585
R147 VTAIL.n231 VTAIL.n230 585
R148 VTAIL.n229 VTAIL.n228 585
R149 VTAIL.n182 VTAIL.n181 585
R150 VTAIL.n223 VTAIL.n222 585
R151 VTAIL.n221 VTAIL.n220 585
R152 VTAIL.n219 VTAIL.n185 585
R153 VTAIL.n189 VTAIL.n186 585
R154 VTAIL.n214 VTAIL.n213 585
R155 VTAIL.n212 VTAIL.n211 585
R156 VTAIL.n191 VTAIL.n190 585
R157 VTAIL.n206 VTAIL.n205 585
R158 VTAIL.n204 VTAIL.n203 585
R159 VTAIL.n195 VTAIL.n194 585
R160 VTAIL.n198 VTAIL.n197 585
R161 VTAIL.t11 VTAIL.n374 329.038
R162 VTAIL.t15 VTAIL.n314 329.038
R163 VTAIL.t3 VTAIL.n256 329.038
R164 VTAIL.t0 VTAIL.n196 329.038
R165 VTAIL.t5 VTAIL.n431 329.038
R166 VTAIL.t7 VTAIL.n19 329.038
R167 VTAIL.t9 VTAIL.n77 329.038
R168 VTAIL.t8 VTAIL.n137 329.038
R169 VTAIL.n432 VTAIL.n429 171.744
R170 VTAIL.n439 VTAIL.n429 171.744
R171 VTAIL.n440 VTAIL.n439 171.744
R172 VTAIL.n440 VTAIL.n425 171.744
R173 VTAIL.n447 VTAIL.n425 171.744
R174 VTAIL.n449 VTAIL.n447 171.744
R175 VTAIL.n449 VTAIL.n448 171.744
R176 VTAIL.n448 VTAIL.n421 171.744
R177 VTAIL.n457 VTAIL.n421 171.744
R178 VTAIL.n458 VTAIL.n457 171.744
R179 VTAIL.n458 VTAIL.n417 171.744
R180 VTAIL.n465 VTAIL.n417 171.744
R181 VTAIL.n466 VTAIL.n465 171.744
R182 VTAIL.n20 VTAIL.n17 171.744
R183 VTAIL.n27 VTAIL.n17 171.744
R184 VTAIL.n28 VTAIL.n27 171.744
R185 VTAIL.n28 VTAIL.n13 171.744
R186 VTAIL.n35 VTAIL.n13 171.744
R187 VTAIL.n37 VTAIL.n35 171.744
R188 VTAIL.n37 VTAIL.n36 171.744
R189 VTAIL.n36 VTAIL.n9 171.744
R190 VTAIL.n45 VTAIL.n9 171.744
R191 VTAIL.n46 VTAIL.n45 171.744
R192 VTAIL.n46 VTAIL.n5 171.744
R193 VTAIL.n53 VTAIL.n5 171.744
R194 VTAIL.n54 VTAIL.n53 171.744
R195 VTAIL.n78 VTAIL.n75 171.744
R196 VTAIL.n85 VTAIL.n75 171.744
R197 VTAIL.n86 VTAIL.n85 171.744
R198 VTAIL.n86 VTAIL.n71 171.744
R199 VTAIL.n93 VTAIL.n71 171.744
R200 VTAIL.n95 VTAIL.n93 171.744
R201 VTAIL.n95 VTAIL.n94 171.744
R202 VTAIL.n94 VTAIL.n67 171.744
R203 VTAIL.n103 VTAIL.n67 171.744
R204 VTAIL.n104 VTAIL.n103 171.744
R205 VTAIL.n104 VTAIL.n63 171.744
R206 VTAIL.n111 VTAIL.n63 171.744
R207 VTAIL.n112 VTAIL.n111 171.744
R208 VTAIL.n138 VTAIL.n135 171.744
R209 VTAIL.n145 VTAIL.n135 171.744
R210 VTAIL.n146 VTAIL.n145 171.744
R211 VTAIL.n146 VTAIL.n131 171.744
R212 VTAIL.n153 VTAIL.n131 171.744
R213 VTAIL.n155 VTAIL.n153 171.744
R214 VTAIL.n155 VTAIL.n154 171.744
R215 VTAIL.n154 VTAIL.n127 171.744
R216 VTAIL.n163 VTAIL.n127 171.744
R217 VTAIL.n164 VTAIL.n163 171.744
R218 VTAIL.n164 VTAIL.n123 171.744
R219 VTAIL.n171 VTAIL.n123 171.744
R220 VTAIL.n172 VTAIL.n171 171.744
R221 VTAIL.n408 VTAIL.n407 171.744
R222 VTAIL.n407 VTAIL.n359 171.744
R223 VTAIL.n400 VTAIL.n359 171.744
R224 VTAIL.n400 VTAIL.n399 171.744
R225 VTAIL.n399 VTAIL.n363 171.744
R226 VTAIL.n367 VTAIL.n363 171.744
R227 VTAIL.n391 VTAIL.n367 171.744
R228 VTAIL.n391 VTAIL.n390 171.744
R229 VTAIL.n390 VTAIL.n368 171.744
R230 VTAIL.n383 VTAIL.n368 171.744
R231 VTAIL.n383 VTAIL.n382 171.744
R232 VTAIL.n382 VTAIL.n372 171.744
R233 VTAIL.n375 VTAIL.n372 171.744
R234 VTAIL.n348 VTAIL.n347 171.744
R235 VTAIL.n347 VTAIL.n299 171.744
R236 VTAIL.n340 VTAIL.n299 171.744
R237 VTAIL.n340 VTAIL.n339 171.744
R238 VTAIL.n339 VTAIL.n303 171.744
R239 VTAIL.n307 VTAIL.n303 171.744
R240 VTAIL.n331 VTAIL.n307 171.744
R241 VTAIL.n331 VTAIL.n330 171.744
R242 VTAIL.n330 VTAIL.n308 171.744
R243 VTAIL.n323 VTAIL.n308 171.744
R244 VTAIL.n323 VTAIL.n322 171.744
R245 VTAIL.n322 VTAIL.n312 171.744
R246 VTAIL.n315 VTAIL.n312 171.744
R247 VTAIL.n290 VTAIL.n289 171.744
R248 VTAIL.n289 VTAIL.n241 171.744
R249 VTAIL.n282 VTAIL.n241 171.744
R250 VTAIL.n282 VTAIL.n281 171.744
R251 VTAIL.n281 VTAIL.n245 171.744
R252 VTAIL.n249 VTAIL.n245 171.744
R253 VTAIL.n273 VTAIL.n249 171.744
R254 VTAIL.n273 VTAIL.n272 171.744
R255 VTAIL.n272 VTAIL.n250 171.744
R256 VTAIL.n265 VTAIL.n250 171.744
R257 VTAIL.n265 VTAIL.n264 171.744
R258 VTAIL.n264 VTAIL.n254 171.744
R259 VTAIL.n257 VTAIL.n254 171.744
R260 VTAIL.n230 VTAIL.n229 171.744
R261 VTAIL.n229 VTAIL.n181 171.744
R262 VTAIL.n222 VTAIL.n181 171.744
R263 VTAIL.n222 VTAIL.n221 171.744
R264 VTAIL.n221 VTAIL.n185 171.744
R265 VTAIL.n189 VTAIL.n185 171.744
R266 VTAIL.n213 VTAIL.n189 171.744
R267 VTAIL.n213 VTAIL.n212 171.744
R268 VTAIL.n212 VTAIL.n190 171.744
R269 VTAIL.n205 VTAIL.n190 171.744
R270 VTAIL.n205 VTAIL.n204 171.744
R271 VTAIL.n204 VTAIL.n194 171.744
R272 VTAIL.n197 VTAIL.n194 171.744
R273 VTAIL.n432 VTAIL.t5 85.8723
R274 VTAIL.n20 VTAIL.t7 85.8723
R275 VTAIL.n78 VTAIL.t9 85.8723
R276 VTAIL.n138 VTAIL.t8 85.8723
R277 VTAIL.n375 VTAIL.t11 85.8723
R278 VTAIL.n315 VTAIL.t15 85.8723
R279 VTAIL.n257 VTAIL.t3 85.8723
R280 VTAIL.n197 VTAIL.t0 85.8723
R281 VTAIL.n355 VTAIL.n354 61.3207
R282 VTAIL.n237 VTAIL.n236 61.3207
R283 VTAIL.n1 VTAIL.n0 61.3205
R284 VTAIL.n119 VTAIL.n118 61.3205
R285 VTAIL.n471 VTAIL.n470 34.3187
R286 VTAIL.n59 VTAIL.n58 34.3187
R287 VTAIL.n117 VTAIL.n116 34.3187
R288 VTAIL.n177 VTAIL.n176 34.3187
R289 VTAIL.n413 VTAIL.n412 34.3187
R290 VTAIL.n353 VTAIL.n352 34.3187
R291 VTAIL.n295 VTAIL.n294 34.3187
R292 VTAIL.n235 VTAIL.n234 34.3187
R293 VTAIL.n471 VTAIL.n413 22.1686
R294 VTAIL.n235 VTAIL.n177 22.1686
R295 VTAIL.n456 VTAIL.n455 13.1884
R296 VTAIL.n44 VTAIL.n43 13.1884
R297 VTAIL.n102 VTAIL.n101 13.1884
R298 VTAIL.n162 VTAIL.n161 13.1884
R299 VTAIL.n398 VTAIL.n397 13.1884
R300 VTAIL.n338 VTAIL.n337 13.1884
R301 VTAIL.n280 VTAIL.n279 13.1884
R302 VTAIL.n220 VTAIL.n219 13.1884
R303 VTAIL.n454 VTAIL.n422 12.8005
R304 VTAIL.n459 VTAIL.n420 12.8005
R305 VTAIL.n42 VTAIL.n10 12.8005
R306 VTAIL.n47 VTAIL.n8 12.8005
R307 VTAIL.n100 VTAIL.n68 12.8005
R308 VTAIL.n105 VTAIL.n66 12.8005
R309 VTAIL.n160 VTAIL.n128 12.8005
R310 VTAIL.n165 VTAIL.n126 12.8005
R311 VTAIL.n401 VTAIL.n362 12.8005
R312 VTAIL.n396 VTAIL.n364 12.8005
R313 VTAIL.n341 VTAIL.n302 12.8005
R314 VTAIL.n336 VTAIL.n304 12.8005
R315 VTAIL.n283 VTAIL.n244 12.8005
R316 VTAIL.n278 VTAIL.n246 12.8005
R317 VTAIL.n223 VTAIL.n184 12.8005
R318 VTAIL.n218 VTAIL.n186 12.8005
R319 VTAIL.n451 VTAIL.n450 12.0247
R320 VTAIL.n460 VTAIL.n418 12.0247
R321 VTAIL.n39 VTAIL.n38 12.0247
R322 VTAIL.n48 VTAIL.n6 12.0247
R323 VTAIL.n97 VTAIL.n96 12.0247
R324 VTAIL.n106 VTAIL.n64 12.0247
R325 VTAIL.n157 VTAIL.n156 12.0247
R326 VTAIL.n166 VTAIL.n124 12.0247
R327 VTAIL.n402 VTAIL.n360 12.0247
R328 VTAIL.n393 VTAIL.n392 12.0247
R329 VTAIL.n342 VTAIL.n300 12.0247
R330 VTAIL.n333 VTAIL.n332 12.0247
R331 VTAIL.n284 VTAIL.n242 12.0247
R332 VTAIL.n275 VTAIL.n274 12.0247
R333 VTAIL.n224 VTAIL.n182 12.0247
R334 VTAIL.n215 VTAIL.n214 12.0247
R335 VTAIL.n446 VTAIL.n424 11.249
R336 VTAIL.n464 VTAIL.n463 11.249
R337 VTAIL.n34 VTAIL.n12 11.249
R338 VTAIL.n52 VTAIL.n51 11.249
R339 VTAIL.n92 VTAIL.n70 11.249
R340 VTAIL.n110 VTAIL.n109 11.249
R341 VTAIL.n152 VTAIL.n130 11.249
R342 VTAIL.n170 VTAIL.n169 11.249
R343 VTAIL.n406 VTAIL.n405 11.249
R344 VTAIL.n389 VTAIL.n366 11.249
R345 VTAIL.n346 VTAIL.n345 11.249
R346 VTAIL.n329 VTAIL.n306 11.249
R347 VTAIL.n288 VTAIL.n287 11.249
R348 VTAIL.n271 VTAIL.n248 11.249
R349 VTAIL.n228 VTAIL.n227 11.249
R350 VTAIL.n211 VTAIL.n188 11.249
R351 VTAIL.n433 VTAIL.n431 10.7239
R352 VTAIL.n21 VTAIL.n19 10.7239
R353 VTAIL.n79 VTAIL.n77 10.7239
R354 VTAIL.n139 VTAIL.n137 10.7239
R355 VTAIL.n376 VTAIL.n374 10.7239
R356 VTAIL.n316 VTAIL.n314 10.7239
R357 VTAIL.n258 VTAIL.n256 10.7239
R358 VTAIL.n198 VTAIL.n196 10.7239
R359 VTAIL.n445 VTAIL.n426 10.4732
R360 VTAIL.n467 VTAIL.n416 10.4732
R361 VTAIL.n33 VTAIL.n14 10.4732
R362 VTAIL.n55 VTAIL.n4 10.4732
R363 VTAIL.n91 VTAIL.n72 10.4732
R364 VTAIL.n113 VTAIL.n62 10.4732
R365 VTAIL.n151 VTAIL.n132 10.4732
R366 VTAIL.n173 VTAIL.n122 10.4732
R367 VTAIL.n409 VTAIL.n358 10.4732
R368 VTAIL.n388 VTAIL.n369 10.4732
R369 VTAIL.n349 VTAIL.n298 10.4732
R370 VTAIL.n328 VTAIL.n309 10.4732
R371 VTAIL.n291 VTAIL.n240 10.4732
R372 VTAIL.n270 VTAIL.n251 10.4732
R373 VTAIL.n231 VTAIL.n180 10.4732
R374 VTAIL.n210 VTAIL.n191 10.4732
R375 VTAIL.n442 VTAIL.n441 9.69747
R376 VTAIL.n468 VTAIL.n414 9.69747
R377 VTAIL.n30 VTAIL.n29 9.69747
R378 VTAIL.n56 VTAIL.n2 9.69747
R379 VTAIL.n88 VTAIL.n87 9.69747
R380 VTAIL.n114 VTAIL.n60 9.69747
R381 VTAIL.n148 VTAIL.n147 9.69747
R382 VTAIL.n174 VTAIL.n120 9.69747
R383 VTAIL.n410 VTAIL.n356 9.69747
R384 VTAIL.n385 VTAIL.n384 9.69747
R385 VTAIL.n350 VTAIL.n296 9.69747
R386 VTAIL.n325 VTAIL.n324 9.69747
R387 VTAIL.n292 VTAIL.n238 9.69747
R388 VTAIL.n267 VTAIL.n266 9.69747
R389 VTAIL.n232 VTAIL.n178 9.69747
R390 VTAIL.n207 VTAIL.n206 9.69747
R391 VTAIL.n470 VTAIL.n469 9.45567
R392 VTAIL.n58 VTAIL.n57 9.45567
R393 VTAIL.n116 VTAIL.n115 9.45567
R394 VTAIL.n176 VTAIL.n175 9.45567
R395 VTAIL.n412 VTAIL.n411 9.45567
R396 VTAIL.n352 VTAIL.n351 9.45567
R397 VTAIL.n294 VTAIL.n293 9.45567
R398 VTAIL.n234 VTAIL.n233 9.45567
R399 VTAIL.n469 VTAIL.n468 9.3005
R400 VTAIL.n416 VTAIL.n415 9.3005
R401 VTAIL.n463 VTAIL.n462 9.3005
R402 VTAIL.n461 VTAIL.n460 9.3005
R403 VTAIL.n420 VTAIL.n419 9.3005
R404 VTAIL.n435 VTAIL.n434 9.3005
R405 VTAIL.n437 VTAIL.n436 9.3005
R406 VTAIL.n428 VTAIL.n427 9.3005
R407 VTAIL.n443 VTAIL.n442 9.3005
R408 VTAIL.n445 VTAIL.n444 9.3005
R409 VTAIL.n424 VTAIL.n423 9.3005
R410 VTAIL.n452 VTAIL.n451 9.3005
R411 VTAIL.n454 VTAIL.n453 9.3005
R412 VTAIL.n57 VTAIL.n56 9.3005
R413 VTAIL.n4 VTAIL.n3 9.3005
R414 VTAIL.n51 VTAIL.n50 9.3005
R415 VTAIL.n49 VTAIL.n48 9.3005
R416 VTAIL.n8 VTAIL.n7 9.3005
R417 VTAIL.n23 VTAIL.n22 9.3005
R418 VTAIL.n25 VTAIL.n24 9.3005
R419 VTAIL.n16 VTAIL.n15 9.3005
R420 VTAIL.n31 VTAIL.n30 9.3005
R421 VTAIL.n33 VTAIL.n32 9.3005
R422 VTAIL.n12 VTAIL.n11 9.3005
R423 VTAIL.n40 VTAIL.n39 9.3005
R424 VTAIL.n42 VTAIL.n41 9.3005
R425 VTAIL.n115 VTAIL.n114 9.3005
R426 VTAIL.n62 VTAIL.n61 9.3005
R427 VTAIL.n109 VTAIL.n108 9.3005
R428 VTAIL.n107 VTAIL.n106 9.3005
R429 VTAIL.n66 VTAIL.n65 9.3005
R430 VTAIL.n81 VTAIL.n80 9.3005
R431 VTAIL.n83 VTAIL.n82 9.3005
R432 VTAIL.n74 VTAIL.n73 9.3005
R433 VTAIL.n89 VTAIL.n88 9.3005
R434 VTAIL.n91 VTAIL.n90 9.3005
R435 VTAIL.n70 VTAIL.n69 9.3005
R436 VTAIL.n98 VTAIL.n97 9.3005
R437 VTAIL.n100 VTAIL.n99 9.3005
R438 VTAIL.n175 VTAIL.n174 9.3005
R439 VTAIL.n122 VTAIL.n121 9.3005
R440 VTAIL.n169 VTAIL.n168 9.3005
R441 VTAIL.n167 VTAIL.n166 9.3005
R442 VTAIL.n126 VTAIL.n125 9.3005
R443 VTAIL.n141 VTAIL.n140 9.3005
R444 VTAIL.n143 VTAIL.n142 9.3005
R445 VTAIL.n134 VTAIL.n133 9.3005
R446 VTAIL.n149 VTAIL.n148 9.3005
R447 VTAIL.n151 VTAIL.n150 9.3005
R448 VTAIL.n130 VTAIL.n129 9.3005
R449 VTAIL.n158 VTAIL.n157 9.3005
R450 VTAIL.n160 VTAIL.n159 9.3005
R451 VTAIL.n378 VTAIL.n377 9.3005
R452 VTAIL.n380 VTAIL.n379 9.3005
R453 VTAIL.n371 VTAIL.n370 9.3005
R454 VTAIL.n386 VTAIL.n385 9.3005
R455 VTAIL.n388 VTAIL.n387 9.3005
R456 VTAIL.n366 VTAIL.n365 9.3005
R457 VTAIL.n394 VTAIL.n393 9.3005
R458 VTAIL.n396 VTAIL.n395 9.3005
R459 VTAIL.n411 VTAIL.n410 9.3005
R460 VTAIL.n358 VTAIL.n357 9.3005
R461 VTAIL.n405 VTAIL.n404 9.3005
R462 VTAIL.n403 VTAIL.n402 9.3005
R463 VTAIL.n362 VTAIL.n361 9.3005
R464 VTAIL.n318 VTAIL.n317 9.3005
R465 VTAIL.n320 VTAIL.n319 9.3005
R466 VTAIL.n311 VTAIL.n310 9.3005
R467 VTAIL.n326 VTAIL.n325 9.3005
R468 VTAIL.n328 VTAIL.n327 9.3005
R469 VTAIL.n306 VTAIL.n305 9.3005
R470 VTAIL.n334 VTAIL.n333 9.3005
R471 VTAIL.n336 VTAIL.n335 9.3005
R472 VTAIL.n351 VTAIL.n350 9.3005
R473 VTAIL.n298 VTAIL.n297 9.3005
R474 VTAIL.n345 VTAIL.n344 9.3005
R475 VTAIL.n343 VTAIL.n342 9.3005
R476 VTAIL.n302 VTAIL.n301 9.3005
R477 VTAIL.n260 VTAIL.n259 9.3005
R478 VTAIL.n262 VTAIL.n261 9.3005
R479 VTAIL.n253 VTAIL.n252 9.3005
R480 VTAIL.n268 VTAIL.n267 9.3005
R481 VTAIL.n270 VTAIL.n269 9.3005
R482 VTAIL.n248 VTAIL.n247 9.3005
R483 VTAIL.n276 VTAIL.n275 9.3005
R484 VTAIL.n278 VTAIL.n277 9.3005
R485 VTAIL.n293 VTAIL.n292 9.3005
R486 VTAIL.n240 VTAIL.n239 9.3005
R487 VTAIL.n287 VTAIL.n286 9.3005
R488 VTAIL.n285 VTAIL.n284 9.3005
R489 VTAIL.n244 VTAIL.n243 9.3005
R490 VTAIL.n200 VTAIL.n199 9.3005
R491 VTAIL.n202 VTAIL.n201 9.3005
R492 VTAIL.n193 VTAIL.n192 9.3005
R493 VTAIL.n208 VTAIL.n207 9.3005
R494 VTAIL.n210 VTAIL.n209 9.3005
R495 VTAIL.n188 VTAIL.n187 9.3005
R496 VTAIL.n216 VTAIL.n215 9.3005
R497 VTAIL.n218 VTAIL.n217 9.3005
R498 VTAIL.n233 VTAIL.n232 9.3005
R499 VTAIL.n180 VTAIL.n179 9.3005
R500 VTAIL.n227 VTAIL.n226 9.3005
R501 VTAIL.n225 VTAIL.n224 9.3005
R502 VTAIL.n184 VTAIL.n183 9.3005
R503 VTAIL.n438 VTAIL.n428 8.92171
R504 VTAIL.n26 VTAIL.n16 8.92171
R505 VTAIL.n84 VTAIL.n74 8.92171
R506 VTAIL.n144 VTAIL.n134 8.92171
R507 VTAIL.n381 VTAIL.n371 8.92171
R508 VTAIL.n321 VTAIL.n311 8.92171
R509 VTAIL.n263 VTAIL.n253 8.92171
R510 VTAIL.n203 VTAIL.n193 8.92171
R511 VTAIL.n437 VTAIL.n430 8.14595
R512 VTAIL.n25 VTAIL.n18 8.14595
R513 VTAIL.n83 VTAIL.n76 8.14595
R514 VTAIL.n143 VTAIL.n136 8.14595
R515 VTAIL.n380 VTAIL.n373 8.14595
R516 VTAIL.n320 VTAIL.n313 8.14595
R517 VTAIL.n262 VTAIL.n255 8.14595
R518 VTAIL.n202 VTAIL.n195 8.14595
R519 VTAIL.n434 VTAIL.n433 7.3702
R520 VTAIL.n22 VTAIL.n21 7.3702
R521 VTAIL.n80 VTAIL.n79 7.3702
R522 VTAIL.n140 VTAIL.n139 7.3702
R523 VTAIL.n377 VTAIL.n376 7.3702
R524 VTAIL.n317 VTAIL.n316 7.3702
R525 VTAIL.n259 VTAIL.n258 7.3702
R526 VTAIL.n199 VTAIL.n198 7.3702
R527 VTAIL.n434 VTAIL.n430 5.81868
R528 VTAIL.n22 VTAIL.n18 5.81868
R529 VTAIL.n80 VTAIL.n76 5.81868
R530 VTAIL.n140 VTAIL.n136 5.81868
R531 VTAIL.n377 VTAIL.n373 5.81868
R532 VTAIL.n317 VTAIL.n313 5.81868
R533 VTAIL.n259 VTAIL.n255 5.81868
R534 VTAIL.n199 VTAIL.n195 5.81868
R535 VTAIL.n438 VTAIL.n437 5.04292
R536 VTAIL.n26 VTAIL.n25 5.04292
R537 VTAIL.n84 VTAIL.n83 5.04292
R538 VTAIL.n144 VTAIL.n143 5.04292
R539 VTAIL.n381 VTAIL.n380 5.04292
R540 VTAIL.n321 VTAIL.n320 5.04292
R541 VTAIL.n263 VTAIL.n262 5.04292
R542 VTAIL.n203 VTAIL.n202 5.04292
R543 VTAIL.n441 VTAIL.n428 4.26717
R544 VTAIL.n470 VTAIL.n414 4.26717
R545 VTAIL.n29 VTAIL.n16 4.26717
R546 VTAIL.n58 VTAIL.n2 4.26717
R547 VTAIL.n87 VTAIL.n74 4.26717
R548 VTAIL.n116 VTAIL.n60 4.26717
R549 VTAIL.n147 VTAIL.n134 4.26717
R550 VTAIL.n176 VTAIL.n120 4.26717
R551 VTAIL.n412 VTAIL.n356 4.26717
R552 VTAIL.n384 VTAIL.n371 4.26717
R553 VTAIL.n352 VTAIL.n296 4.26717
R554 VTAIL.n324 VTAIL.n311 4.26717
R555 VTAIL.n294 VTAIL.n238 4.26717
R556 VTAIL.n266 VTAIL.n253 4.26717
R557 VTAIL.n234 VTAIL.n178 4.26717
R558 VTAIL.n206 VTAIL.n193 4.26717
R559 VTAIL.n442 VTAIL.n426 3.49141
R560 VTAIL.n468 VTAIL.n467 3.49141
R561 VTAIL.n30 VTAIL.n14 3.49141
R562 VTAIL.n56 VTAIL.n55 3.49141
R563 VTAIL.n88 VTAIL.n72 3.49141
R564 VTAIL.n114 VTAIL.n113 3.49141
R565 VTAIL.n148 VTAIL.n132 3.49141
R566 VTAIL.n174 VTAIL.n173 3.49141
R567 VTAIL.n410 VTAIL.n409 3.49141
R568 VTAIL.n385 VTAIL.n369 3.49141
R569 VTAIL.n350 VTAIL.n349 3.49141
R570 VTAIL.n325 VTAIL.n309 3.49141
R571 VTAIL.n292 VTAIL.n291 3.49141
R572 VTAIL.n267 VTAIL.n251 3.49141
R573 VTAIL.n232 VTAIL.n231 3.49141
R574 VTAIL.n207 VTAIL.n191 3.49141
R575 VTAIL.n0 VTAIL.t1 3.01301
R576 VTAIL.n0 VTAIL.t6 3.01301
R577 VTAIL.n118 VTAIL.t13 3.01301
R578 VTAIL.n118 VTAIL.t12 3.01301
R579 VTAIL.n354 VTAIL.t10 3.01301
R580 VTAIL.n354 VTAIL.t14 3.01301
R581 VTAIL.n236 VTAIL.t4 3.01301
R582 VTAIL.n236 VTAIL.t2 3.01301
R583 VTAIL.n446 VTAIL.n445 2.71565
R584 VTAIL.n464 VTAIL.n416 2.71565
R585 VTAIL.n34 VTAIL.n33 2.71565
R586 VTAIL.n52 VTAIL.n4 2.71565
R587 VTAIL.n92 VTAIL.n91 2.71565
R588 VTAIL.n110 VTAIL.n62 2.71565
R589 VTAIL.n152 VTAIL.n151 2.71565
R590 VTAIL.n170 VTAIL.n122 2.71565
R591 VTAIL.n406 VTAIL.n358 2.71565
R592 VTAIL.n389 VTAIL.n388 2.71565
R593 VTAIL.n346 VTAIL.n298 2.71565
R594 VTAIL.n329 VTAIL.n328 2.71565
R595 VTAIL.n288 VTAIL.n240 2.71565
R596 VTAIL.n271 VTAIL.n270 2.71565
R597 VTAIL.n228 VTAIL.n180 2.71565
R598 VTAIL.n211 VTAIL.n210 2.71565
R599 VTAIL.n435 VTAIL.n431 2.41282
R600 VTAIL.n23 VTAIL.n19 2.41282
R601 VTAIL.n81 VTAIL.n77 2.41282
R602 VTAIL.n141 VTAIL.n137 2.41282
R603 VTAIL.n378 VTAIL.n374 2.41282
R604 VTAIL.n318 VTAIL.n314 2.41282
R605 VTAIL.n260 VTAIL.n256 2.41282
R606 VTAIL.n200 VTAIL.n196 2.41282
R607 VTAIL.n450 VTAIL.n424 1.93989
R608 VTAIL.n463 VTAIL.n418 1.93989
R609 VTAIL.n38 VTAIL.n12 1.93989
R610 VTAIL.n51 VTAIL.n6 1.93989
R611 VTAIL.n96 VTAIL.n70 1.93989
R612 VTAIL.n109 VTAIL.n64 1.93989
R613 VTAIL.n156 VTAIL.n130 1.93989
R614 VTAIL.n169 VTAIL.n124 1.93989
R615 VTAIL.n405 VTAIL.n360 1.93989
R616 VTAIL.n392 VTAIL.n366 1.93989
R617 VTAIL.n345 VTAIL.n300 1.93989
R618 VTAIL.n332 VTAIL.n306 1.93989
R619 VTAIL.n287 VTAIL.n242 1.93989
R620 VTAIL.n274 VTAIL.n248 1.93989
R621 VTAIL.n227 VTAIL.n182 1.93989
R622 VTAIL.n214 VTAIL.n188 1.93989
R623 VTAIL.n451 VTAIL.n422 1.16414
R624 VTAIL.n460 VTAIL.n459 1.16414
R625 VTAIL.n39 VTAIL.n10 1.16414
R626 VTAIL.n48 VTAIL.n47 1.16414
R627 VTAIL.n97 VTAIL.n68 1.16414
R628 VTAIL.n106 VTAIL.n105 1.16414
R629 VTAIL.n157 VTAIL.n128 1.16414
R630 VTAIL.n166 VTAIL.n165 1.16414
R631 VTAIL.n402 VTAIL.n401 1.16414
R632 VTAIL.n393 VTAIL.n364 1.16414
R633 VTAIL.n342 VTAIL.n341 1.16414
R634 VTAIL.n333 VTAIL.n304 1.16414
R635 VTAIL.n284 VTAIL.n283 1.16414
R636 VTAIL.n275 VTAIL.n246 1.16414
R637 VTAIL.n224 VTAIL.n223 1.16414
R638 VTAIL.n215 VTAIL.n186 1.16414
R639 VTAIL.n237 VTAIL.n235 0.5005
R640 VTAIL.n295 VTAIL.n237 0.5005
R641 VTAIL.n355 VTAIL.n353 0.5005
R642 VTAIL.n413 VTAIL.n355 0.5005
R643 VTAIL.n177 VTAIL.n119 0.5005
R644 VTAIL.n119 VTAIL.n117 0.5005
R645 VTAIL.n59 VTAIL.n1 0.5005
R646 VTAIL.n353 VTAIL.n295 0.470328
R647 VTAIL.n117 VTAIL.n59 0.470328
R648 VTAIL VTAIL.n471 0.44231
R649 VTAIL.n455 VTAIL.n454 0.388379
R650 VTAIL.n456 VTAIL.n420 0.388379
R651 VTAIL.n43 VTAIL.n42 0.388379
R652 VTAIL.n44 VTAIL.n8 0.388379
R653 VTAIL.n101 VTAIL.n100 0.388379
R654 VTAIL.n102 VTAIL.n66 0.388379
R655 VTAIL.n161 VTAIL.n160 0.388379
R656 VTAIL.n162 VTAIL.n126 0.388379
R657 VTAIL.n398 VTAIL.n362 0.388379
R658 VTAIL.n397 VTAIL.n396 0.388379
R659 VTAIL.n338 VTAIL.n302 0.388379
R660 VTAIL.n337 VTAIL.n336 0.388379
R661 VTAIL.n280 VTAIL.n244 0.388379
R662 VTAIL.n279 VTAIL.n278 0.388379
R663 VTAIL.n220 VTAIL.n184 0.388379
R664 VTAIL.n219 VTAIL.n218 0.388379
R665 VTAIL.n436 VTAIL.n435 0.155672
R666 VTAIL.n436 VTAIL.n427 0.155672
R667 VTAIL.n443 VTAIL.n427 0.155672
R668 VTAIL.n444 VTAIL.n443 0.155672
R669 VTAIL.n444 VTAIL.n423 0.155672
R670 VTAIL.n452 VTAIL.n423 0.155672
R671 VTAIL.n453 VTAIL.n452 0.155672
R672 VTAIL.n453 VTAIL.n419 0.155672
R673 VTAIL.n461 VTAIL.n419 0.155672
R674 VTAIL.n462 VTAIL.n461 0.155672
R675 VTAIL.n462 VTAIL.n415 0.155672
R676 VTAIL.n469 VTAIL.n415 0.155672
R677 VTAIL.n24 VTAIL.n23 0.155672
R678 VTAIL.n24 VTAIL.n15 0.155672
R679 VTAIL.n31 VTAIL.n15 0.155672
R680 VTAIL.n32 VTAIL.n31 0.155672
R681 VTAIL.n32 VTAIL.n11 0.155672
R682 VTAIL.n40 VTAIL.n11 0.155672
R683 VTAIL.n41 VTAIL.n40 0.155672
R684 VTAIL.n41 VTAIL.n7 0.155672
R685 VTAIL.n49 VTAIL.n7 0.155672
R686 VTAIL.n50 VTAIL.n49 0.155672
R687 VTAIL.n50 VTAIL.n3 0.155672
R688 VTAIL.n57 VTAIL.n3 0.155672
R689 VTAIL.n82 VTAIL.n81 0.155672
R690 VTAIL.n82 VTAIL.n73 0.155672
R691 VTAIL.n89 VTAIL.n73 0.155672
R692 VTAIL.n90 VTAIL.n89 0.155672
R693 VTAIL.n90 VTAIL.n69 0.155672
R694 VTAIL.n98 VTAIL.n69 0.155672
R695 VTAIL.n99 VTAIL.n98 0.155672
R696 VTAIL.n99 VTAIL.n65 0.155672
R697 VTAIL.n107 VTAIL.n65 0.155672
R698 VTAIL.n108 VTAIL.n107 0.155672
R699 VTAIL.n108 VTAIL.n61 0.155672
R700 VTAIL.n115 VTAIL.n61 0.155672
R701 VTAIL.n142 VTAIL.n141 0.155672
R702 VTAIL.n142 VTAIL.n133 0.155672
R703 VTAIL.n149 VTAIL.n133 0.155672
R704 VTAIL.n150 VTAIL.n149 0.155672
R705 VTAIL.n150 VTAIL.n129 0.155672
R706 VTAIL.n158 VTAIL.n129 0.155672
R707 VTAIL.n159 VTAIL.n158 0.155672
R708 VTAIL.n159 VTAIL.n125 0.155672
R709 VTAIL.n167 VTAIL.n125 0.155672
R710 VTAIL.n168 VTAIL.n167 0.155672
R711 VTAIL.n168 VTAIL.n121 0.155672
R712 VTAIL.n175 VTAIL.n121 0.155672
R713 VTAIL.n411 VTAIL.n357 0.155672
R714 VTAIL.n404 VTAIL.n357 0.155672
R715 VTAIL.n404 VTAIL.n403 0.155672
R716 VTAIL.n403 VTAIL.n361 0.155672
R717 VTAIL.n395 VTAIL.n361 0.155672
R718 VTAIL.n395 VTAIL.n394 0.155672
R719 VTAIL.n394 VTAIL.n365 0.155672
R720 VTAIL.n387 VTAIL.n365 0.155672
R721 VTAIL.n387 VTAIL.n386 0.155672
R722 VTAIL.n386 VTAIL.n370 0.155672
R723 VTAIL.n379 VTAIL.n370 0.155672
R724 VTAIL.n379 VTAIL.n378 0.155672
R725 VTAIL.n351 VTAIL.n297 0.155672
R726 VTAIL.n344 VTAIL.n297 0.155672
R727 VTAIL.n344 VTAIL.n343 0.155672
R728 VTAIL.n343 VTAIL.n301 0.155672
R729 VTAIL.n335 VTAIL.n301 0.155672
R730 VTAIL.n335 VTAIL.n334 0.155672
R731 VTAIL.n334 VTAIL.n305 0.155672
R732 VTAIL.n327 VTAIL.n305 0.155672
R733 VTAIL.n327 VTAIL.n326 0.155672
R734 VTAIL.n326 VTAIL.n310 0.155672
R735 VTAIL.n319 VTAIL.n310 0.155672
R736 VTAIL.n319 VTAIL.n318 0.155672
R737 VTAIL.n293 VTAIL.n239 0.155672
R738 VTAIL.n286 VTAIL.n239 0.155672
R739 VTAIL.n286 VTAIL.n285 0.155672
R740 VTAIL.n285 VTAIL.n243 0.155672
R741 VTAIL.n277 VTAIL.n243 0.155672
R742 VTAIL.n277 VTAIL.n276 0.155672
R743 VTAIL.n276 VTAIL.n247 0.155672
R744 VTAIL.n269 VTAIL.n247 0.155672
R745 VTAIL.n269 VTAIL.n268 0.155672
R746 VTAIL.n268 VTAIL.n252 0.155672
R747 VTAIL.n261 VTAIL.n252 0.155672
R748 VTAIL.n261 VTAIL.n260 0.155672
R749 VTAIL.n233 VTAIL.n179 0.155672
R750 VTAIL.n226 VTAIL.n179 0.155672
R751 VTAIL.n226 VTAIL.n225 0.155672
R752 VTAIL.n225 VTAIL.n183 0.155672
R753 VTAIL.n217 VTAIL.n183 0.155672
R754 VTAIL.n217 VTAIL.n216 0.155672
R755 VTAIL.n216 VTAIL.n187 0.155672
R756 VTAIL.n209 VTAIL.n187 0.155672
R757 VTAIL.n209 VTAIL.n208 0.155672
R758 VTAIL.n208 VTAIL.n192 0.155672
R759 VTAIL.n201 VTAIL.n192 0.155672
R760 VTAIL.n201 VTAIL.n200 0.155672
R761 VTAIL VTAIL.n1 0.0586897
R762 B.n205 B.t0 1264.46
R763 B.n94 B.t6 1264.46
R764 B.n36 B.t9 1264.46
R765 B.n30 B.t3 1264.46
R766 B.n282 B.n281 585
R767 B.n280 B.n75 585
R768 B.n279 B.n278 585
R769 B.n277 B.n76 585
R770 B.n276 B.n275 585
R771 B.n274 B.n77 585
R772 B.n273 B.n272 585
R773 B.n271 B.n78 585
R774 B.n270 B.n269 585
R775 B.n268 B.n79 585
R776 B.n267 B.n266 585
R777 B.n265 B.n80 585
R778 B.n264 B.n263 585
R779 B.n262 B.n81 585
R780 B.n261 B.n260 585
R781 B.n259 B.n82 585
R782 B.n258 B.n257 585
R783 B.n256 B.n83 585
R784 B.n255 B.n254 585
R785 B.n253 B.n84 585
R786 B.n252 B.n251 585
R787 B.n250 B.n85 585
R788 B.n249 B.n248 585
R789 B.n247 B.n86 585
R790 B.n246 B.n245 585
R791 B.n244 B.n87 585
R792 B.n243 B.n242 585
R793 B.n241 B.n88 585
R794 B.n240 B.n239 585
R795 B.n238 B.n89 585
R796 B.n237 B.n236 585
R797 B.n235 B.n90 585
R798 B.n234 B.n233 585
R799 B.n232 B.n91 585
R800 B.n231 B.n230 585
R801 B.n229 B.n92 585
R802 B.n228 B.n227 585
R803 B.n226 B.n93 585
R804 B.n224 B.n223 585
R805 B.n222 B.n96 585
R806 B.n221 B.n220 585
R807 B.n219 B.n97 585
R808 B.n218 B.n217 585
R809 B.n216 B.n98 585
R810 B.n215 B.n214 585
R811 B.n213 B.n99 585
R812 B.n212 B.n211 585
R813 B.n210 B.n100 585
R814 B.n209 B.n208 585
R815 B.n204 B.n101 585
R816 B.n203 B.n202 585
R817 B.n201 B.n102 585
R818 B.n200 B.n199 585
R819 B.n198 B.n103 585
R820 B.n197 B.n196 585
R821 B.n195 B.n104 585
R822 B.n194 B.n193 585
R823 B.n192 B.n105 585
R824 B.n191 B.n190 585
R825 B.n189 B.n106 585
R826 B.n188 B.n187 585
R827 B.n186 B.n107 585
R828 B.n185 B.n184 585
R829 B.n183 B.n108 585
R830 B.n182 B.n181 585
R831 B.n180 B.n109 585
R832 B.n179 B.n178 585
R833 B.n177 B.n110 585
R834 B.n176 B.n175 585
R835 B.n174 B.n111 585
R836 B.n173 B.n172 585
R837 B.n171 B.n112 585
R838 B.n170 B.n169 585
R839 B.n168 B.n113 585
R840 B.n167 B.n166 585
R841 B.n165 B.n114 585
R842 B.n164 B.n163 585
R843 B.n162 B.n115 585
R844 B.n161 B.n160 585
R845 B.n159 B.n116 585
R846 B.n158 B.n157 585
R847 B.n156 B.n117 585
R848 B.n155 B.n154 585
R849 B.n153 B.n118 585
R850 B.n152 B.n151 585
R851 B.n150 B.n119 585
R852 B.n283 B.n74 585
R853 B.n285 B.n284 585
R854 B.n286 B.n73 585
R855 B.n288 B.n287 585
R856 B.n289 B.n72 585
R857 B.n291 B.n290 585
R858 B.n292 B.n71 585
R859 B.n294 B.n293 585
R860 B.n295 B.n70 585
R861 B.n297 B.n296 585
R862 B.n298 B.n69 585
R863 B.n300 B.n299 585
R864 B.n301 B.n68 585
R865 B.n303 B.n302 585
R866 B.n304 B.n67 585
R867 B.n306 B.n305 585
R868 B.n307 B.n66 585
R869 B.n309 B.n308 585
R870 B.n310 B.n65 585
R871 B.n312 B.n311 585
R872 B.n313 B.n64 585
R873 B.n315 B.n314 585
R874 B.n316 B.n63 585
R875 B.n318 B.n317 585
R876 B.n319 B.n62 585
R877 B.n321 B.n320 585
R878 B.n322 B.n61 585
R879 B.n324 B.n323 585
R880 B.n325 B.n60 585
R881 B.n327 B.n326 585
R882 B.n328 B.n59 585
R883 B.n330 B.n329 585
R884 B.n331 B.n58 585
R885 B.n333 B.n332 585
R886 B.n463 B.n10 585
R887 B.n462 B.n461 585
R888 B.n460 B.n11 585
R889 B.n459 B.n458 585
R890 B.n457 B.n12 585
R891 B.n456 B.n455 585
R892 B.n454 B.n13 585
R893 B.n453 B.n452 585
R894 B.n451 B.n14 585
R895 B.n450 B.n449 585
R896 B.n448 B.n15 585
R897 B.n447 B.n446 585
R898 B.n445 B.n16 585
R899 B.n444 B.n443 585
R900 B.n442 B.n17 585
R901 B.n441 B.n440 585
R902 B.n439 B.n18 585
R903 B.n438 B.n437 585
R904 B.n436 B.n19 585
R905 B.n435 B.n434 585
R906 B.n433 B.n20 585
R907 B.n432 B.n431 585
R908 B.n430 B.n21 585
R909 B.n429 B.n428 585
R910 B.n427 B.n22 585
R911 B.n426 B.n425 585
R912 B.n424 B.n23 585
R913 B.n423 B.n422 585
R914 B.n421 B.n24 585
R915 B.n420 B.n419 585
R916 B.n418 B.n25 585
R917 B.n417 B.n416 585
R918 B.n415 B.n26 585
R919 B.n414 B.n413 585
R920 B.n412 B.n27 585
R921 B.n411 B.n410 585
R922 B.n409 B.n28 585
R923 B.n408 B.n407 585
R924 B.n405 B.n29 585
R925 B.n404 B.n403 585
R926 B.n402 B.n32 585
R927 B.n401 B.n400 585
R928 B.n399 B.n33 585
R929 B.n398 B.n397 585
R930 B.n396 B.n34 585
R931 B.n395 B.n394 585
R932 B.n393 B.n35 585
R933 B.n392 B.n391 585
R934 B.n390 B.n389 585
R935 B.n388 B.n39 585
R936 B.n387 B.n386 585
R937 B.n385 B.n40 585
R938 B.n384 B.n383 585
R939 B.n382 B.n41 585
R940 B.n381 B.n380 585
R941 B.n379 B.n42 585
R942 B.n378 B.n377 585
R943 B.n376 B.n43 585
R944 B.n375 B.n374 585
R945 B.n373 B.n44 585
R946 B.n372 B.n371 585
R947 B.n370 B.n45 585
R948 B.n369 B.n368 585
R949 B.n367 B.n46 585
R950 B.n366 B.n365 585
R951 B.n364 B.n47 585
R952 B.n363 B.n362 585
R953 B.n361 B.n48 585
R954 B.n360 B.n359 585
R955 B.n358 B.n49 585
R956 B.n357 B.n356 585
R957 B.n355 B.n50 585
R958 B.n354 B.n353 585
R959 B.n352 B.n51 585
R960 B.n351 B.n350 585
R961 B.n349 B.n52 585
R962 B.n348 B.n347 585
R963 B.n346 B.n53 585
R964 B.n345 B.n344 585
R965 B.n343 B.n54 585
R966 B.n342 B.n341 585
R967 B.n340 B.n55 585
R968 B.n339 B.n338 585
R969 B.n337 B.n56 585
R970 B.n336 B.n335 585
R971 B.n334 B.n57 585
R972 B.n465 B.n464 585
R973 B.n466 B.n9 585
R974 B.n468 B.n467 585
R975 B.n469 B.n8 585
R976 B.n471 B.n470 585
R977 B.n472 B.n7 585
R978 B.n474 B.n473 585
R979 B.n475 B.n6 585
R980 B.n477 B.n476 585
R981 B.n478 B.n5 585
R982 B.n480 B.n479 585
R983 B.n481 B.n4 585
R984 B.n483 B.n482 585
R985 B.n484 B.n3 585
R986 B.n486 B.n485 585
R987 B.n487 B.n0 585
R988 B.n2 B.n1 585
R989 B.n128 B.n127 585
R990 B.n129 B.n126 585
R991 B.n131 B.n130 585
R992 B.n132 B.n125 585
R993 B.n134 B.n133 585
R994 B.n135 B.n124 585
R995 B.n137 B.n136 585
R996 B.n138 B.n123 585
R997 B.n140 B.n139 585
R998 B.n141 B.n122 585
R999 B.n143 B.n142 585
R1000 B.n144 B.n121 585
R1001 B.n146 B.n145 585
R1002 B.n147 B.n120 585
R1003 B.n149 B.n148 585
R1004 B.n148 B.n119 497.305
R1005 B.n283 B.n282 497.305
R1006 B.n332 B.n57 497.305
R1007 B.n464 B.n463 497.305
R1008 B.n94 B.t7 365.199
R1009 B.n36 B.t11 365.199
R1010 B.n205 B.t1 365.199
R1011 B.n30 B.t5 365.199
R1012 B.n95 B.t8 353.95
R1013 B.n37 B.t10 353.95
R1014 B.n206 B.t2 353.95
R1015 B.n31 B.t4 353.95
R1016 B.n489 B.n488 256.663
R1017 B.n488 B.n487 235.042
R1018 B.n488 B.n2 235.042
R1019 B.n152 B.n119 163.367
R1020 B.n153 B.n152 163.367
R1021 B.n154 B.n153 163.367
R1022 B.n154 B.n117 163.367
R1023 B.n158 B.n117 163.367
R1024 B.n159 B.n158 163.367
R1025 B.n160 B.n159 163.367
R1026 B.n160 B.n115 163.367
R1027 B.n164 B.n115 163.367
R1028 B.n165 B.n164 163.367
R1029 B.n166 B.n165 163.367
R1030 B.n166 B.n113 163.367
R1031 B.n170 B.n113 163.367
R1032 B.n171 B.n170 163.367
R1033 B.n172 B.n171 163.367
R1034 B.n172 B.n111 163.367
R1035 B.n176 B.n111 163.367
R1036 B.n177 B.n176 163.367
R1037 B.n178 B.n177 163.367
R1038 B.n178 B.n109 163.367
R1039 B.n182 B.n109 163.367
R1040 B.n183 B.n182 163.367
R1041 B.n184 B.n183 163.367
R1042 B.n184 B.n107 163.367
R1043 B.n188 B.n107 163.367
R1044 B.n189 B.n188 163.367
R1045 B.n190 B.n189 163.367
R1046 B.n190 B.n105 163.367
R1047 B.n194 B.n105 163.367
R1048 B.n195 B.n194 163.367
R1049 B.n196 B.n195 163.367
R1050 B.n196 B.n103 163.367
R1051 B.n200 B.n103 163.367
R1052 B.n201 B.n200 163.367
R1053 B.n202 B.n201 163.367
R1054 B.n202 B.n101 163.367
R1055 B.n209 B.n101 163.367
R1056 B.n210 B.n209 163.367
R1057 B.n211 B.n210 163.367
R1058 B.n211 B.n99 163.367
R1059 B.n215 B.n99 163.367
R1060 B.n216 B.n215 163.367
R1061 B.n217 B.n216 163.367
R1062 B.n217 B.n97 163.367
R1063 B.n221 B.n97 163.367
R1064 B.n222 B.n221 163.367
R1065 B.n223 B.n222 163.367
R1066 B.n223 B.n93 163.367
R1067 B.n228 B.n93 163.367
R1068 B.n229 B.n228 163.367
R1069 B.n230 B.n229 163.367
R1070 B.n230 B.n91 163.367
R1071 B.n234 B.n91 163.367
R1072 B.n235 B.n234 163.367
R1073 B.n236 B.n235 163.367
R1074 B.n236 B.n89 163.367
R1075 B.n240 B.n89 163.367
R1076 B.n241 B.n240 163.367
R1077 B.n242 B.n241 163.367
R1078 B.n242 B.n87 163.367
R1079 B.n246 B.n87 163.367
R1080 B.n247 B.n246 163.367
R1081 B.n248 B.n247 163.367
R1082 B.n248 B.n85 163.367
R1083 B.n252 B.n85 163.367
R1084 B.n253 B.n252 163.367
R1085 B.n254 B.n253 163.367
R1086 B.n254 B.n83 163.367
R1087 B.n258 B.n83 163.367
R1088 B.n259 B.n258 163.367
R1089 B.n260 B.n259 163.367
R1090 B.n260 B.n81 163.367
R1091 B.n264 B.n81 163.367
R1092 B.n265 B.n264 163.367
R1093 B.n266 B.n265 163.367
R1094 B.n266 B.n79 163.367
R1095 B.n270 B.n79 163.367
R1096 B.n271 B.n270 163.367
R1097 B.n272 B.n271 163.367
R1098 B.n272 B.n77 163.367
R1099 B.n276 B.n77 163.367
R1100 B.n277 B.n276 163.367
R1101 B.n278 B.n277 163.367
R1102 B.n278 B.n75 163.367
R1103 B.n282 B.n75 163.367
R1104 B.n332 B.n331 163.367
R1105 B.n331 B.n330 163.367
R1106 B.n330 B.n59 163.367
R1107 B.n326 B.n59 163.367
R1108 B.n326 B.n325 163.367
R1109 B.n325 B.n324 163.367
R1110 B.n324 B.n61 163.367
R1111 B.n320 B.n61 163.367
R1112 B.n320 B.n319 163.367
R1113 B.n319 B.n318 163.367
R1114 B.n318 B.n63 163.367
R1115 B.n314 B.n63 163.367
R1116 B.n314 B.n313 163.367
R1117 B.n313 B.n312 163.367
R1118 B.n312 B.n65 163.367
R1119 B.n308 B.n65 163.367
R1120 B.n308 B.n307 163.367
R1121 B.n307 B.n306 163.367
R1122 B.n306 B.n67 163.367
R1123 B.n302 B.n67 163.367
R1124 B.n302 B.n301 163.367
R1125 B.n301 B.n300 163.367
R1126 B.n300 B.n69 163.367
R1127 B.n296 B.n69 163.367
R1128 B.n296 B.n295 163.367
R1129 B.n295 B.n294 163.367
R1130 B.n294 B.n71 163.367
R1131 B.n290 B.n71 163.367
R1132 B.n290 B.n289 163.367
R1133 B.n289 B.n288 163.367
R1134 B.n288 B.n73 163.367
R1135 B.n284 B.n73 163.367
R1136 B.n284 B.n283 163.367
R1137 B.n463 B.n462 163.367
R1138 B.n462 B.n11 163.367
R1139 B.n458 B.n11 163.367
R1140 B.n458 B.n457 163.367
R1141 B.n457 B.n456 163.367
R1142 B.n456 B.n13 163.367
R1143 B.n452 B.n13 163.367
R1144 B.n452 B.n451 163.367
R1145 B.n451 B.n450 163.367
R1146 B.n450 B.n15 163.367
R1147 B.n446 B.n15 163.367
R1148 B.n446 B.n445 163.367
R1149 B.n445 B.n444 163.367
R1150 B.n444 B.n17 163.367
R1151 B.n440 B.n17 163.367
R1152 B.n440 B.n439 163.367
R1153 B.n439 B.n438 163.367
R1154 B.n438 B.n19 163.367
R1155 B.n434 B.n19 163.367
R1156 B.n434 B.n433 163.367
R1157 B.n433 B.n432 163.367
R1158 B.n432 B.n21 163.367
R1159 B.n428 B.n21 163.367
R1160 B.n428 B.n427 163.367
R1161 B.n427 B.n426 163.367
R1162 B.n426 B.n23 163.367
R1163 B.n422 B.n23 163.367
R1164 B.n422 B.n421 163.367
R1165 B.n421 B.n420 163.367
R1166 B.n420 B.n25 163.367
R1167 B.n416 B.n25 163.367
R1168 B.n416 B.n415 163.367
R1169 B.n415 B.n414 163.367
R1170 B.n414 B.n27 163.367
R1171 B.n410 B.n27 163.367
R1172 B.n410 B.n409 163.367
R1173 B.n409 B.n408 163.367
R1174 B.n408 B.n29 163.367
R1175 B.n403 B.n29 163.367
R1176 B.n403 B.n402 163.367
R1177 B.n402 B.n401 163.367
R1178 B.n401 B.n33 163.367
R1179 B.n397 B.n33 163.367
R1180 B.n397 B.n396 163.367
R1181 B.n396 B.n395 163.367
R1182 B.n395 B.n35 163.367
R1183 B.n391 B.n35 163.367
R1184 B.n391 B.n390 163.367
R1185 B.n390 B.n39 163.367
R1186 B.n386 B.n39 163.367
R1187 B.n386 B.n385 163.367
R1188 B.n385 B.n384 163.367
R1189 B.n384 B.n41 163.367
R1190 B.n380 B.n41 163.367
R1191 B.n380 B.n379 163.367
R1192 B.n379 B.n378 163.367
R1193 B.n378 B.n43 163.367
R1194 B.n374 B.n43 163.367
R1195 B.n374 B.n373 163.367
R1196 B.n373 B.n372 163.367
R1197 B.n372 B.n45 163.367
R1198 B.n368 B.n45 163.367
R1199 B.n368 B.n367 163.367
R1200 B.n367 B.n366 163.367
R1201 B.n366 B.n47 163.367
R1202 B.n362 B.n47 163.367
R1203 B.n362 B.n361 163.367
R1204 B.n361 B.n360 163.367
R1205 B.n360 B.n49 163.367
R1206 B.n356 B.n49 163.367
R1207 B.n356 B.n355 163.367
R1208 B.n355 B.n354 163.367
R1209 B.n354 B.n51 163.367
R1210 B.n350 B.n51 163.367
R1211 B.n350 B.n349 163.367
R1212 B.n349 B.n348 163.367
R1213 B.n348 B.n53 163.367
R1214 B.n344 B.n53 163.367
R1215 B.n344 B.n343 163.367
R1216 B.n343 B.n342 163.367
R1217 B.n342 B.n55 163.367
R1218 B.n338 B.n55 163.367
R1219 B.n338 B.n337 163.367
R1220 B.n337 B.n336 163.367
R1221 B.n336 B.n57 163.367
R1222 B.n464 B.n9 163.367
R1223 B.n468 B.n9 163.367
R1224 B.n469 B.n468 163.367
R1225 B.n470 B.n469 163.367
R1226 B.n470 B.n7 163.367
R1227 B.n474 B.n7 163.367
R1228 B.n475 B.n474 163.367
R1229 B.n476 B.n475 163.367
R1230 B.n476 B.n5 163.367
R1231 B.n480 B.n5 163.367
R1232 B.n481 B.n480 163.367
R1233 B.n482 B.n481 163.367
R1234 B.n482 B.n3 163.367
R1235 B.n486 B.n3 163.367
R1236 B.n487 B.n486 163.367
R1237 B.n128 B.n2 163.367
R1238 B.n129 B.n128 163.367
R1239 B.n130 B.n129 163.367
R1240 B.n130 B.n125 163.367
R1241 B.n134 B.n125 163.367
R1242 B.n135 B.n134 163.367
R1243 B.n136 B.n135 163.367
R1244 B.n136 B.n123 163.367
R1245 B.n140 B.n123 163.367
R1246 B.n141 B.n140 163.367
R1247 B.n142 B.n141 163.367
R1248 B.n142 B.n121 163.367
R1249 B.n146 B.n121 163.367
R1250 B.n147 B.n146 163.367
R1251 B.n148 B.n147 163.367
R1252 B.n207 B.n206 59.5399
R1253 B.n225 B.n95 59.5399
R1254 B.n38 B.n37 59.5399
R1255 B.n406 B.n31 59.5399
R1256 B.n465 B.n10 32.3127
R1257 B.n334 B.n333 32.3127
R1258 B.n281 B.n74 32.3127
R1259 B.n150 B.n149 32.3127
R1260 B B.n489 18.0485
R1261 B.n206 B.n205 11.249
R1262 B.n95 B.n94 11.249
R1263 B.n37 B.n36 11.249
R1264 B.n31 B.n30 11.249
R1265 B.n466 B.n465 10.6151
R1266 B.n467 B.n466 10.6151
R1267 B.n467 B.n8 10.6151
R1268 B.n471 B.n8 10.6151
R1269 B.n472 B.n471 10.6151
R1270 B.n473 B.n472 10.6151
R1271 B.n473 B.n6 10.6151
R1272 B.n477 B.n6 10.6151
R1273 B.n478 B.n477 10.6151
R1274 B.n479 B.n478 10.6151
R1275 B.n479 B.n4 10.6151
R1276 B.n483 B.n4 10.6151
R1277 B.n484 B.n483 10.6151
R1278 B.n485 B.n484 10.6151
R1279 B.n485 B.n0 10.6151
R1280 B.n461 B.n10 10.6151
R1281 B.n461 B.n460 10.6151
R1282 B.n460 B.n459 10.6151
R1283 B.n459 B.n12 10.6151
R1284 B.n455 B.n12 10.6151
R1285 B.n455 B.n454 10.6151
R1286 B.n454 B.n453 10.6151
R1287 B.n453 B.n14 10.6151
R1288 B.n449 B.n14 10.6151
R1289 B.n449 B.n448 10.6151
R1290 B.n448 B.n447 10.6151
R1291 B.n447 B.n16 10.6151
R1292 B.n443 B.n16 10.6151
R1293 B.n443 B.n442 10.6151
R1294 B.n442 B.n441 10.6151
R1295 B.n441 B.n18 10.6151
R1296 B.n437 B.n18 10.6151
R1297 B.n437 B.n436 10.6151
R1298 B.n436 B.n435 10.6151
R1299 B.n435 B.n20 10.6151
R1300 B.n431 B.n20 10.6151
R1301 B.n431 B.n430 10.6151
R1302 B.n430 B.n429 10.6151
R1303 B.n429 B.n22 10.6151
R1304 B.n425 B.n22 10.6151
R1305 B.n425 B.n424 10.6151
R1306 B.n424 B.n423 10.6151
R1307 B.n423 B.n24 10.6151
R1308 B.n419 B.n24 10.6151
R1309 B.n419 B.n418 10.6151
R1310 B.n418 B.n417 10.6151
R1311 B.n417 B.n26 10.6151
R1312 B.n413 B.n26 10.6151
R1313 B.n413 B.n412 10.6151
R1314 B.n412 B.n411 10.6151
R1315 B.n411 B.n28 10.6151
R1316 B.n407 B.n28 10.6151
R1317 B.n405 B.n404 10.6151
R1318 B.n404 B.n32 10.6151
R1319 B.n400 B.n32 10.6151
R1320 B.n400 B.n399 10.6151
R1321 B.n399 B.n398 10.6151
R1322 B.n398 B.n34 10.6151
R1323 B.n394 B.n34 10.6151
R1324 B.n394 B.n393 10.6151
R1325 B.n393 B.n392 10.6151
R1326 B.n389 B.n388 10.6151
R1327 B.n388 B.n387 10.6151
R1328 B.n387 B.n40 10.6151
R1329 B.n383 B.n40 10.6151
R1330 B.n383 B.n382 10.6151
R1331 B.n382 B.n381 10.6151
R1332 B.n381 B.n42 10.6151
R1333 B.n377 B.n42 10.6151
R1334 B.n377 B.n376 10.6151
R1335 B.n376 B.n375 10.6151
R1336 B.n375 B.n44 10.6151
R1337 B.n371 B.n44 10.6151
R1338 B.n371 B.n370 10.6151
R1339 B.n370 B.n369 10.6151
R1340 B.n369 B.n46 10.6151
R1341 B.n365 B.n46 10.6151
R1342 B.n365 B.n364 10.6151
R1343 B.n364 B.n363 10.6151
R1344 B.n363 B.n48 10.6151
R1345 B.n359 B.n48 10.6151
R1346 B.n359 B.n358 10.6151
R1347 B.n358 B.n357 10.6151
R1348 B.n357 B.n50 10.6151
R1349 B.n353 B.n50 10.6151
R1350 B.n353 B.n352 10.6151
R1351 B.n352 B.n351 10.6151
R1352 B.n351 B.n52 10.6151
R1353 B.n347 B.n52 10.6151
R1354 B.n347 B.n346 10.6151
R1355 B.n346 B.n345 10.6151
R1356 B.n345 B.n54 10.6151
R1357 B.n341 B.n54 10.6151
R1358 B.n341 B.n340 10.6151
R1359 B.n340 B.n339 10.6151
R1360 B.n339 B.n56 10.6151
R1361 B.n335 B.n56 10.6151
R1362 B.n335 B.n334 10.6151
R1363 B.n333 B.n58 10.6151
R1364 B.n329 B.n58 10.6151
R1365 B.n329 B.n328 10.6151
R1366 B.n328 B.n327 10.6151
R1367 B.n327 B.n60 10.6151
R1368 B.n323 B.n60 10.6151
R1369 B.n323 B.n322 10.6151
R1370 B.n322 B.n321 10.6151
R1371 B.n321 B.n62 10.6151
R1372 B.n317 B.n62 10.6151
R1373 B.n317 B.n316 10.6151
R1374 B.n316 B.n315 10.6151
R1375 B.n315 B.n64 10.6151
R1376 B.n311 B.n64 10.6151
R1377 B.n311 B.n310 10.6151
R1378 B.n310 B.n309 10.6151
R1379 B.n309 B.n66 10.6151
R1380 B.n305 B.n66 10.6151
R1381 B.n305 B.n304 10.6151
R1382 B.n304 B.n303 10.6151
R1383 B.n303 B.n68 10.6151
R1384 B.n299 B.n68 10.6151
R1385 B.n299 B.n298 10.6151
R1386 B.n298 B.n297 10.6151
R1387 B.n297 B.n70 10.6151
R1388 B.n293 B.n70 10.6151
R1389 B.n293 B.n292 10.6151
R1390 B.n292 B.n291 10.6151
R1391 B.n291 B.n72 10.6151
R1392 B.n287 B.n72 10.6151
R1393 B.n287 B.n286 10.6151
R1394 B.n286 B.n285 10.6151
R1395 B.n285 B.n74 10.6151
R1396 B.n127 B.n1 10.6151
R1397 B.n127 B.n126 10.6151
R1398 B.n131 B.n126 10.6151
R1399 B.n132 B.n131 10.6151
R1400 B.n133 B.n132 10.6151
R1401 B.n133 B.n124 10.6151
R1402 B.n137 B.n124 10.6151
R1403 B.n138 B.n137 10.6151
R1404 B.n139 B.n138 10.6151
R1405 B.n139 B.n122 10.6151
R1406 B.n143 B.n122 10.6151
R1407 B.n144 B.n143 10.6151
R1408 B.n145 B.n144 10.6151
R1409 B.n145 B.n120 10.6151
R1410 B.n149 B.n120 10.6151
R1411 B.n151 B.n150 10.6151
R1412 B.n151 B.n118 10.6151
R1413 B.n155 B.n118 10.6151
R1414 B.n156 B.n155 10.6151
R1415 B.n157 B.n156 10.6151
R1416 B.n157 B.n116 10.6151
R1417 B.n161 B.n116 10.6151
R1418 B.n162 B.n161 10.6151
R1419 B.n163 B.n162 10.6151
R1420 B.n163 B.n114 10.6151
R1421 B.n167 B.n114 10.6151
R1422 B.n168 B.n167 10.6151
R1423 B.n169 B.n168 10.6151
R1424 B.n169 B.n112 10.6151
R1425 B.n173 B.n112 10.6151
R1426 B.n174 B.n173 10.6151
R1427 B.n175 B.n174 10.6151
R1428 B.n175 B.n110 10.6151
R1429 B.n179 B.n110 10.6151
R1430 B.n180 B.n179 10.6151
R1431 B.n181 B.n180 10.6151
R1432 B.n181 B.n108 10.6151
R1433 B.n185 B.n108 10.6151
R1434 B.n186 B.n185 10.6151
R1435 B.n187 B.n186 10.6151
R1436 B.n187 B.n106 10.6151
R1437 B.n191 B.n106 10.6151
R1438 B.n192 B.n191 10.6151
R1439 B.n193 B.n192 10.6151
R1440 B.n193 B.n104 10.6151
R1441 B.n197 B.n104 10.6151
R1442 B.n198 B.n197 10.6151
R1443 B.n199 B.n198 10.6151
R1444 B.n199 B.n102 10.6151
R1445 B.n203 B.n102 10.6151
R1446 B.n204 B.n203 10.6151
R1447 B.n208 B.n204 10.6151
R1448 B.n212 B.n100 10.6151
R1449 B.n213 B.n212 10.6151
R1450 B.n214 B.n213 10.6151
R1451 B.n214 B.n98 10.6151
R1452 B.n218 B.n98 10.6151
R1453 B.n219 B.n218 10.6151
R1454 B.n220 B.n219 10.6151
R1455 B.n220 B.n96 10.6151
R1456 B.n224 B.n96 10.6151
R1457 B.n227 B.n226 10.6151
R1458 B.n227 B.n92 10.6151
R1459 B.n231 B.n92 10.6151
R1460 B.n232 B.n231 10.6151
R1461 B.n233 B.n232 10.6151
R1462 B.n233 B.n90 10.6151
R1463 B.n237 B.n90 10.6151
R1464 B.n238 B.n237 10.6151
R1465 B.n239 B.n238 10.6151
R1466 B.n239 B.n88 10.6151
R1467 B.n243 B.n88 10.6151
R1468 B.n244 B.n243 10.6151
R1469 B.n245 B.n244 10.6151
R1470 B.n245 B.n86 10.6151
R1471 B.n249 B.n86 10.6151
R1472 B.n250 B.n249 10.6151
R1473 B.n251 B.n250 10.6151
R1474 B.n251 B.n84 10.6151
R1475 B.n255 B.n84 10.6151
R1476 B.n256 B.n255 10.6151
R1477 B.n257 B.n256 10.6151
R1478 B.n257 B.n82 10.6151
R1479 B.n261 B.n82 10.6151
R1480 B.n262 B.n261 10.6151
R1481 B.n263 B.n262 10.6151
R1482 B.n263 B.n80 10.6151
R1483 B.n267 B.n80 10.6151
R1484 B.n268 B.n267 10.6151
R1485 B.n269 B.n268 10.6151
R1486 B.n269 B.n78 10.6151
R1487 B.n273 B.n78 10.6151
R1488 B.n274 B.n273 10.6151
R1489 B.n275 B.n274 10.6151
R1490 B.n275 B.n76 10.6151
R1491 B.n279 B.n76 10.6151
R1492 B.n280 B.n279 10.6151
R1493 B.n281 B.n280 10.6151
R1494 B.n407 B.n406 9.36635
R1495 B.n389 B.n38 9.36635
R1496 B.n208 B.n207 9.36635
R1497 B.n226 B.n225 9.36635
R1498 B.n489 B.n0 8.11757
R1499 B.n489 B.n1 8.11757
R1500 B.n406 B.n405 1.24928
R1501 B.n392 B.n38 1.24928
R1502 B.n207 B.n100 1.24928
R1503 B.n225 B.n224 1.24928
R1504 VN.n5 VN.t3 1220.48
R1505 VN.n1 VN.t6 1220.48
R1506 VN.n12 VN.t5 1220.48
R1507 VN.n8 VN.t1 1220.48
R1508 VN.n4 VN.t4 1166.44
R1509 VN.n2 VN.t0 1166.44
R1510 VN.n11 VN.t2 1166.44
R1511 VN.n9 VN.t7 1166.44
R1512 VN.n8 VN.n7 161.489
R1513 VN.n1 VN.n0 161.489
R1514 VN.n6 VN.n5 161.3
R1515 VN.n13 VN.n12 161.3
R1516 VN.n10 VN.n7 161.3
R1517 VN.n3 VN.n0 161.3
R1518 VN.n3 VN.n2 42.3581
R1519 VN.n4 VN.n3 42.3581
R1520 VN.n11 VN.n10 42.3581
R1521 VN.n10 VN.n9 42.3581
R1522 VN VN.n13 39.4872
R1523 VN.n2 VN.n1 30.6732
R1524 VN.n5 VN.n4 30.6732
R1525 VN.n12 VN.n11 30.6732
R1526 VN.n9 VN.n8 30.6732
R1527 VN.n13 VN.n7 0.189894
R1528 VN.n6 VN.n0 0.189894
R1529 VN VN.n6 0.0516364
R1530 VDD2.n2 VDD2.n1 78.194
R1531 VDD2.n2 VDD2.n0 78.194
R1532 VDD2 VDD2.n5 78.1911
R1533 VDD2.n4 VDD2.n3 77.9995
R1534 VDD2.n4 VDD2.n2 35.267
R1535 VDD2.n5 VDD2.t0 3.01301
R1536 VDD2.n5 VDD2.t6 3.01301
R1537 VDD2.n3 VDD2.t2 3.01301
R1538 VDD2.n3 VDD2.t5 3.01301
R1539 VDD2.n1 VDD2.t3 3.01301
R1540 VDD2.n1 VDD2.t4 3.01301
R1541 VDD2.n0 VDD2.t1 3.01301
R1542 VDD2.n0 VDD2.t7 3.01301
R1543 VDD2 VDD2.n4 0.30869
C0 VDD1 B 0.899923f
C1 VDD1 VN 0.14719f
C2 VDD2 B 0.923009f
C3 VTAIL VP 2.33049f
C4 VDD2 VN 2.7193f
C5 w_n1550_n3126# VDD1 1.07762f
C6 w_n1550_n3126# VDD2 1.09409f
C7 B VP 0.972509f
C8 VN VP 4.56201f
C9 w_n1550_n3126# VP 2.66692f
C10 VDD2 VDD1 0.606984f
C11 VTAIL B 3.14691f
C12 VTAIL VN 2.31638f
C13 w_n1550_n3126# VTAIL 3.95987f
C14 VDD1 VP 2.84122f
C15 VDD2 VP 0.269317f
C16 B VN 0.659332f
C17 w_n1550_n3126# B 6.21825f
C18 w_n1550_n3126# VN 2.47263f
C19 VDD1 VTAIL 16.1659f
C20 VDD2 VTAIL 16.204498f
C21 VDD2 VSUBS 1.343415f
C22 VDD1 VSUBS 1.555757f
C23 VTAIL VSUBS 0.644188f
C24 VN VSUBS 4.41172f
C25 VP VSUBS 1.15674f
C26 B VSUBS 2.267318f
C27 w_n1550_n3126# VSUBS 59.7618f
C28 VDD2.t1 VSUBS 0.299808f
C29 VDD2.t7 VSUBS 0.299808f
C30 VDD2.n0 VSUBS 2.30684f
C31 VDD2.t3 VSUBS 0.299808f
C32 VDD2.t4 VSUBS 0.299808f
C33 VDD2.n1 VSUBS 2.30684f
C34 VDD2.n2 VSUBS 3.27566f
C35 VDD2.t2 VSUBS 0.299808f
C36 VDD2.t5 VSUBS 0.299808f
C37 VDD2.n3 VSUBS 2.30503f
C38 VDD2.n4 VSUBS 3.21579f
C39 VDD2.t0 VSUBS 0.299808f
C40 VDD2.t6 VSUBS 0.299808f
C41 VDD2.n5 VSUBS 2.30681f
C42 VN.n0 VSUBS 0.164997f
C43 VN.t4 VSUBS 0.54737f
C44 VN.t0 VSUBS 0.54737f
C45 VN.t6 VSUBS 0.557558f
C46 VN.n1 VSUBS 0.247334f
C47 VN.n2 VSUBS 0.224777f
C48 VN.n3 VSUBS 0.027329f
C49 VN.n4 VSUBS 0.224777f
C50 VN.t3 VSUBS 0.557558f
C51 VN.n5 VSUBS 0.247224f
C52 VN.n6 VSUBS 0.05558f
C53 VN.n7 VSUBS 0.164997f
C54 VN.t5 VSUBS 0.557558f
C55 VN.t2 VSUBS 0.54737f
C56 VN.t7 VSUBS 0.54737f
C57 VN.t1 VSUBS 0.557558f
C58 VN.n8 VSUBS 0.247334f
C59 VN.n9 VSUBS 0.224777f
C60 VN.n10 VSUBS 0.027329f
C61 VN.n11 VSUBS 0.224777f
C62 VN.n12 VSUBS 0.247224f
C63 VN.n13 VSUBS 2.66763f
C64 B.n0 VSUBS 0.007773f
C65 B.n1 VSUBS 0.007773f
C66 B.n2 VSUBS 0.011496f
C67 B.n3 VSUBS 0.00881f
C68 B.n4 VSUBS 0.00881f
C69 B.n5 VSUBS 0.00881f
C70 B.n6 VSUBS 0.00881f
C71 B.n7 VSUBS 0.00881f
C72 B.n8 VSUBS 0.00881f
C73 B.n9 VSUBS 0.00881f
C74 B.n10 VSUBS 0.021226f
C75 B.n11 VSUBS 0.00881f
C76 B.n12 VSUBS 0.00881f
C77 B.n13 VSUBS 0.00881f
C78 B.n14 VSUBS 0.00881f
C79 B.n15 VSUBS 0.00881f
C80 B.n16 VSUBS 0.00881f
C81 B.n17 VSUBS 0.00881f
C82 B.n18 VSUBS 0.00881f
C83 B.n19 VSUBS 0.00881f
C84 B.n20 VSUBS 0.00881f
C85 B.n21 VSUBS 0.00881f
C86 B.n22 VSUBS 0.00881f
C87 B.n23 VSUBS 0.00881f
C88 B.n24 VSUBS 0.00881f
C89 B.n25 VSUBS 0.00881f
C90 B.n26 VSUBS 0.00881f
C91 B.n27 VSUBS 0.00881f
C92 B.n28 VSUBS 0.00881f
C93 B.n29 VSUBS 0.00881f
C94 B.t4 VSUBS 0.232298f
C95 B.t5 VSUBS 0.240625f
C96 B.t3 VSUBS 0.13295f
C97 B.n30 VSUBS 0.312469f
C98 B.n31 VSUBS 0.282909f
C99 B.n32 VSUBS 0.00881f
C100 B.n33 VSUBS 0.00881f
C101 B.n34 VSUBS 0.00881f
C102 B.n35 VSUBS 0.00881f
C103 B.t10 VSUBS 0.232301f
C104 B.t11 VSUBS 0.240628f
C105 B.t9 VSUBS 0.13295f
C106 B.n36 VSUBS 0.312466f
C107 B.n37 VSUBS 0.282905f
C108 B.n38 VSUBS 0.020411f
C109 B.n39 VSUBS 0.00881f
C110 B.n40 VSUBS 0.00881f
C111 B.n41 VSUBS 0.00881f
C112 B.n42 VSUBS 0.00881f
C113 B.n43 VSUBS 0.00881f
C114 B.n44 VSUBS 0.00881f
C115 B.n45 VSUBS 0.00881f
C116 B.n46 VSUBS 0.00881f
C117 B.n47 VSUBS 0.00881f
C118 B.n48 VSUBS 0.00881f
C119 B.n49 VSUBS 0.00881f
C120 B.n50 VSUBS 0.00881f
C121 B.n51 VSUBS 0.00881f
C122 B.n52 VSUBS 0.00881f
C123 B.n53 VSUBS 0.00881f
C124 B.n54 VSUBS 0.00881f
C125 B.n55 VSUBS 0.00881f
C126 B.n56 VSUBS 0.00881f
C127 B.n57 VSUBS 0.021226f
C128 B.n58 VSUBS 0.00881f
C129 B.n59 VSUBS 0.00881f
C130 B.n60 VSUBS 0.00881f
C131 B.n61 VSUBS 0.00881f
C132 B.n62 VSUBS 0.00881f
C133 B.n63 VSUBS 0.00881f
C134 B.n64 VSUBS 0.00881f
C135 B.n65 VSUBS 0.00881f
C136 B.n66 VSUBS 0.00881f
C137 B.n67 VSUBS 0.00881f
C138 B.n68 VSUBS 0.00881f
C139 B.n69 VSUBS 0.00881f
C140 B.n70 VSUBS 0.00881f
C141 B.n71 VSUBS 0.00881f
C142 B.n72 VSUBS 0.00881f
C143 B.n73 VSUBS 0.00881f
C144 B.n74 VSUBS 0.020764f
C145 B.n75 VSUBS 0.00881f
C146 B.n76 VSUBS 0.00881f
C147 B.n77 VSUBS 0.00881f
C148 B.n78 VSUBS 0.00881f
C149 B.n79 VSUBS 0.00881f
C150 B.n80 VSUBS 0.00881f
C151 B.n81 VSUBS 0.00881f
C152 B.n82 VSUBS 0.00881f
C153 B.n83 VSUBS 0.00881f
C154 B.n84 VSUBS 0.00881f
C155 B.n85 VSUBS 0.00881f
C156 B.n86 VSUBS 0.00881f
C157 B.n87 VSUBS 0.00881f
C158 B.n88 VSUBS 0.00881f
C159 B.n89 VSUBS 0.00881f
C160 B.n90 VSUBS 0.00881f
C161 B.n91 VSUBS 0.00881f
C162 B.n92 VSUBS 0.00881f
C163 B.n93 VSUBS 0.00881f
C164 B.t8 VSUBS 0.232301f
C165 B.t7 VSUBS 0.240628f
C166 B.t6 VSUBS 0.13295f
C167 B.n94 VSUBS 0.312466f
C168 B.n95 VSUBS 0.282905f
C169 B.n96 VSUBS 0.00881f
C170 B.n97 VSUBS 0.00881f
C171 B.n98 VSUBS 0.00881f
C172 B.n99 VSUBS 0.00881f
C173 B.n100 VSUBS 0.004923f
C174 B.n101 VSUBS 0.00881f
C175 B.n102 VSUBS 0.00881f
C176 B.n103 VSUBS 0.00881f
C177 B.n104 VSUBS 0.00881f
C178 B.n105 VSUBS 0.00881f
C179 B.n106 VSUBS 0.00881f
C180 B.n107 VSUBS 0.00881f
C181 B.n108 VSUBS 0.00881f
C182 B.n109 VSUBS 0.00881f
C183 B.n110 VSUBS 0.00881f
C184 B.n111 VSUBS 0.00881f
C185 B.n112 VSUBS 0.00881f
C186 B.n113 VSUBS 0.00881f
C187 B.n114 VSUBS 0.00881f
C188 B.n115 VSUBS 0.00881f
C189 B.n116 VSUBS 0.00881f
C190 B.n117 VSUBS 0.00881f
C191 B.n118 VSUBS 0.00881f
C192 B.n119 VSUBS 0.021226f
C193 B.n120 VSUBS 0.00881f
C194 B.n121 VSUBS 0.00881f
C195 B.n122 VSUBS 0.00881f
C196 B.n123 VSUBS 0.00881f
C197 B.n124 VSUBS 0.00881f
C198 B.n125 VSUBS 0.00881f
C199 B.n126 VSUBS 0.00881f
C200 B.n127 VSUBS 0.00881f
C201 B.n128 VSUBS 0.00881f
C202 B.n129 VSUBS 0.00881f
C203 B.n130 VSUBS 0.00881f
C204 B.n131 VSUBS 0.00881f
C205 B.n132 VSUBS 0.00881f
C206 B.n133 VSUBS 0.00881f
C207 B.n134 VSUBS 0.00881f
C208 B.n135 VSUBS 0.00881f
C209 B.n136 VSUBS 0.00881f
C210 B.n137 VSUBS 0.00881f
C211 B.n138 VSUBS 0.00881f
C212 B.n139 VSUBS 0.00881f
C213 B.n140 VSUBS 0.00881f
C214 B.n141 VSUBS 0.00881f
C215 B.n142 VSUBS 0.00881f
C216 B.n143 VSUBS 0.00881f
C217 B.n144 VSUBS 0.00881f
C218 B.n145 VSUBS 0.00881f
C219 B.n146 VSUBS 0.00881f
C220 B.n147 VSUBS 0.00881f
C221 B.n148 VSUBS 0.019712f
C222 B.n149 VSUBS 0.019712f
C223 B.n150 VSUBS 0.021226f
C224 B.n151 VSUBS 0.00881f
C225 B.n152 VSUBS 0.00881f
C226 B.n153 VSUBS 0.00881f
C227 B.n154 VSUBS 0.00881f
C228 B.n155 VSUBS 0.00881f
C229 B.n156 VSUBS 0.00881f
C230 B.n157 VSUBS 0.00881f
C231 B.n158 VSUBS 0.00881f
C232 B.n159 VSUBS 0.00881f
C233 B.n160 VSUBS 0.00881f
C234 B.n161 VSUBS 0.00881f
C235 B.n162 VSUBS 0.00881f
C236 B.n163 VSUBS 0.00881f
C237 B.n164 VSUBS 0.00881f
C238 B.n165 VSUBS 0.00881f
C239 B.n166 VSUBS 0.00881f
C240 B.n167 VSUBS 0.00881f
C241 B.n168 VSUBS 0.00881f
C242 B.n169 VSUBS 0.00881f
C243 B.n170 VSUBS 0.00881f
C244 B.n171 VSUBS 0.00881f
C245 B.n172 VSUBS 0.00881f
C246 B.n173 VSUBS 0.00881f
C247 B.n174 VSUBS 0.00881f
C248 B.n175 VSUBS 0.00881f
C249 B.n176 VSUBS 0.00881f
C250 B.n177 VSUBS 0.00881f
C251 B.n178 VSUBS 0.00881f
C252 B.n179 VSUBS 0.00881f
C253 B.n180 VSUBS 0.00881f
C254 B.n181 VSUBS 0.00881f
C255 B.n182 VSUBS 0.00881f
C256 B.n183 VSUBS 0.00881f
C257 B.n184 VSUBS 0.00881f
C258 B.n185 VSUBS 0.00881f
C259 B.n186 VSUBS 0.00881f
C260 B.n187 VSUBS 0.00881f
C261 B.n188 VSUBS 0.00881f
C262 B.n189 VSUBS 0.00881f
C263 B.n190 VSUBS 0.00881f
C264 B.n191 VSUBS 0.00881f
C265 B.n192 VSUBS 0.00881f
C266 B.n193 VSUBS 0.00881f
C267 B.n194 VSUBS 0.00881f
C268 B.n195 VSUBS 0.00881f
C269 B.n196 VSUBS 0.00881f
C270 B.n197 VSUBS 0.00881f
C271 B.n198 VSUBS 0.00881f
C272 B.n199 VSUBS 0.00881f
C273 B.n200 VSUBS 0.00881f
C274 B.n201 VSUBS 0.00881f
C275 B.n202 VSUBS 0.00881f
C276 B.n203 VSUBS 0.00881f
C277 B.n204 VSUBS 0.00881f
C278 B.t2 VSUBS 0.232298f
C279 B.t1 VSUBS 0.240625f
C280 B.t0 VSUBS 0.13295f
C281 B.n205 VSUBS 0.312469f
C282 B.n206 VSUBS 0.282909f
C283 B.n207 VSUBS 0.020411f
C284 B.n208 VSUBS 0.008291f
C285 B.n209 VSUBS 0.00881f
C286 B.n210 VSUBS 0.00881f
C287 B.n211 VSUBS 0.00881f
C288 B.n212 VSUBS 0.00881f
C289 B.n213 VSUBS 0.00881f
C290 B.n214 VSUBS 0.00881f
C291 B.n215 VSUBS 0.00881f
C292 B.n216 VSUBS 0.00881f
C293 B.n217 VSUBS 0.00881f
C294 B.n218 VSUBS 0.00881f
C295 B.n219 VSUBS 0.00881f
C296 B.n220 VSUBS 0.00881f
C297 B.n221 VSUBS 0.00881f
C298 B.n222 VSUBS 0.00881f
C299 B.n223 VSUBS 0.00881f
C300 B.n224 VSUBS 0.004923f
C301 B.n225 VSUBS 0.020411f
C302 B.n226 VSUBS 0.008291f
C303 B.n227 VSUBS 0.00881f
C304 B.n228 VSUBS 0.00881f
C305 B.n229 VSUBS 0.00881f
C306 B.n230 VSUBS 0.00881f
C307 B.n231 VSUBS 0.00881f
C308 B.n232 VSUBS 0.00881f
C309 B.n233 VSUBS 0.00881f
C310 B.n234 VSUBS 0.00881f
C311 B.n235 VSUBS 0.00881f
C312 B.n236 VSUBS 0.00881f
C313 B.n237 VSUBS 0.00881f
C314 B.n238 VSUBS 0.00881f
C315 B.n239 VSUBS 0.00881f
C316 B.n240 VSUBS 0.00881f
C317 B.n241 VSUBS 0.00881f
C318 B.n242 VSUBS 0.00881f
C319 B.n243 VSUBS 0.00881f
C320 B.n244 VSUBS 0.00881f
C321 B.n245 VSUBS 0.00881f
C322 B.n246 VSUBS 0.00881f
C323 B.n247 VSUBS 0.00881f
C324 B.n248 VSUBS 0.00881f
C325 B.n249 VSUBS 0.00881f
C326 B.n250 VSUBS 0.00881f
C327 B.n251 VSUBS 0.00881f
C328 B.n252 VSUBS 0.00881f
C329 B.n253 VSUBS 0.00881f
C330 B.n254 VSUBS 0.00881f
C331 B.n255 VSUBS 0.00881f
C332 B.n256 VSUBS 0.00881f
C333 B.n257 VSUBS 0.00881f
C334 B.n258 VSUBS 0.00881f
C335 B.n259 VSUBS 0.00881f
C336 B.n260 VSUBS 0.00881f
C337 B.n261 VSUBS 0.00881f
C338 B.n262 VSUBS 0.00881f
C339 B.n263 VSUBS 0.00881f
C340 B.n264 VSUBS 0.00881f
C341 B.n265 VSUBS 0.00881f
C342 B.n266 VSUBS 0.00881f
C343 B.n267 VSUBS 0.00881f
C344 B.n268 VSUBS 0.00881f
C345 B.n269 VSUBS 0.00881f
C346 B.n270 VSUBS 0.00881f
C347 B.n271 VSUBS 0.00881f
C348 B.n272 VSUBS 0.00881f
C349 B.n273 VSUBS 0.00881f
C350 B.n274 VSUBS 0.00881f
C351 B.n275 VSUBS 0.00881f
C352 B.n276 VSUBS 0.00881f
C353 B.n277 VSUBS 0.00881f
C354 B.n278 VSUBS 0.00881f
C355 B.n279 VSUBS 0.00881f
C356 B.n280 VSUBS 0.00881f
C357 B.n281 VSUBS 0.020174f
C358 B.n282 VSUBS 0.021226f
C359 B.n283 VSUBS 0.019712f
C360 B.n284 VSUBS 0.00881f
C361 B.n285 VSUBS 0.00881f
C362 B.n286 VSUBS 0.00881f
C363 B.n287 VSUBS 0.00881f
C364 B.n288 VSUBS 0.00881f
C365 B.n289 VSUBS 0.00881f
C366 B.n290 VSUBS 0.00881f
C367 B.n291 VSUBS 0.00881f
C368 B.n292 VSUBS 0.00881f
C369 B.n293 VSUBS 0.00881f
C370 B.n294 VSUBS 0.00881f
C371 B.n295 VSUBS 0.00881f
C372 B.n296 VSUBS 0.00881f
C373 B.n297 VSUBS 0.00881f
C374 B.n298 VSUBS 0.00881f
C375 B.n299 VSUBS 0.00881f
C376 B.n300 VSUBS 0.00881f
C377 B.n301 VSUBS 0.00881f
C378 B.n302 VSUBS 0.00881f
C379 B.n303 VSUBS 0.00881f
C380 B.n304 VSUBS 0.00881f
C381 B.n305 VSUBS 0.00881f
C382 B.n306 VSUBS 0.00881f
C383 B.n307 VSUBS 0.00881f
C384 B.n308 VSUBS 0.00881f
C385 B.n309 VSUBS 0.00881f
C386 B.n310 VSUBS 0.00881f
C387 B.n311 VSUBS 0.00881f
C388 B.n312 VSUBS 0.00881f
C389 B.n313 VSUBS 0.00881f
C390 B.n314 VSUBS 0.00881f
C391 B.n315 VSUBS 0.00881f
C392 B.n316 VSUBS 0.00881f
C393 B.n317 VSUBS 0.00881f
C394 B.n318 VSUBS 0.00881f
C395 B.n319 VSUBS 0.00881f
C396 B.n320 VSUBS 0.00881f
C397 B.n321 VSUBS 0.00881f
C398 B.n322 VSUBS 0.00881f
C399 B.n323 VSUBS 0.00881f
C400 B.n324 VSUBS 0.00881f
C401 B.n325 VSUBS 0.00881f
C402 B.n326 VSUBS 0.00881f
C403 B.n327 VSUBS 0.00881f
C404 B.n328 VSUBS 0.00881f
C405 B.n329 VSUBS 0.00881f
C406 B.n330 VSUBS 0.00881f
C407 B.n331 VSUBS 0.00881f
C408 B.n332 VSUBS 0.019712f
C409 B.n333 VSUBS 0.019712f
C410 B.n334 VSUBS 0.021226f
C411 B.n335 VSUBS 0.00881f
C412 B.n336 VSUBS 0.00881f
C413 B.n337 VSUBS 0.00881f
C414 B.n338 VSUBS 0.00881f
C415 B.n339 VSUBS 0.00881f
C416 B.n340 VSUBS 0.00881f
C417 B.n341 VSUBS 0.00881f
C418 B.n342 VSUBS 0.00881f
C419 B.n343 VSUBS 0.00881f
C420 B.n344 VSUBS 0.00881f
C421 B.n345 VSUBS 0.00881f
C422 B.n346 VSUBS 0.00881f
C423 B.n347 VSUBS 0.00881f
C424 B.n348 VSUBS 0.00881f
C425 B.n349 VSUBS 0.00881f
C426 B.n350 VSUBS 0.00881f
C427 B.n351 VSUBS 0.00881f
C428 B.n352 VSUBS 0.00881f
C429 B.n353 VSUBS 0.00881f
C430 B.n354 VSUBS 0.00881f
C431 B.n355 VSUBS 0.00881f
C432 B.n356 VSUBS 0.00881f
C433 B.n357 VSUBS 0.00881f
C434 B.n358 VSUBS 0.00881f
C435 B.n359 VSUBS 0.00881f
C436 B.n360 VSUBS 0.00881f
C437 B.n361 VSUBS 0.00881f
C438 B.n362 VSUBS 0.00881f
C439 B.n363 VSUBS 0.00881f
C440 B.n364 VSUBS 0.00881f
C441 B.n365 VSUBS 0.00881f
C442 B.n366 VSUBS 0.00881f
C443 B.n367 VSUBS 0.00881f
C444 B.n368 VSUBS 0.00881f
C445 B.n369 VSUBS 0.00881f
C446 B.n370 VSUBS 0.00881f
C447 B.n371 VSUBS 0.00881f
C448 B.n372 VSUBS 0.00881f
C449 B.n373 VSUBS 0.00881f
C450 B.n374 VSUBS 0.00881f
C451 B.n375 VSUBS 0.00881f
C452 B.n376 VSUBS 0.00881f
C453 B.n377 VSUBS 0.00881f
C454 B.n378 VSUBS 0.00881f
C455 B.n379 VSUBS 0.00881f
C456 B.n380 VSUBS 0.00881f
C457 B.n381 VSUBS 0.00881f
C458 B.n382 VSUBS 0.00881f
C459 B.n383 VSUBS 0.00881f
C460 B.n384 VSUBS 0.00881f
C461 B.n385 VSUBS 0.00881f
C462 B.n386 VSUBS 0.00881f
C463 B.n387 VSUBS 0.00881f
C464 B.n388 VSUBS 0.00881f
C465 B.n389 VSUBS 0.008291f
C466 B.n390 VSUBS 0.00881f
C467 B.n391 VSUBS 0.00881f
C468 B.n392 VSUBS 0.004923f
C469 B.n393 VSUBS 0.00881f
C470 B.n394 VSUBS 0.00881f
C471 B.n395 VSUBS 0.00881f
C472 B.n396 VSUBS 0.00881f
C473 B.n397 VSUBS 0.00881f
C474 B.n398 VSUBS 0.00881f
C475 B.n399 VSUBS 0.00881f
C476 B.n400 VSUBS 0.00881f
C477 B.n401 VSUBS 0.00881f
C478 B.n402 VSUBS 0.00881f
C479 B.n403 VSUBS 0.00881f
C480 B.n404 VSUBS 0.00881f
C481 B.n405 VSUBS 0.004923f
C482 B.n406 VSUBS 0.020411f
C483 B.n407 VSUBS 0.008291f
C484 B.n408 VSUBS 0.00881f
C485 B.n409 VSUBS 0.00881f
C486 B.n410 VSUBS 0.00881f
C487 B.n411 VSUBS 0.00881f
C488 B.n412 VSUBS 0.00881f
C489 B.n413 VSUBS 0.00881f
C490 B.n414 VSUBS 0.00881f
C491 B.n415 VSUBS 0.00881f
C492 B.n416 VSUBS 0.00881f
C493 B.n417 VSUBS 0.00881f
C494 B.n418 VSUBS 0.00881f
C495 B.n419 VSUBS 0.00881f
C496 B.n420 VSUBS 0.00881f
C497 B.n421 VSUBS 0.00881f
C498 B.n422 VSUBS 0.00881f
C499 B.n423 VSUBS 0.00881f
C500 B.n424 VSUBS 0.00881f
C501 B.n425 VSUBS 0.00881f
C502 B.n426 VSUBS 0.00881f
C503 B.n427 VSUBS 0.00881f
C504 B.n428 VSUBS 0.00881f
C505 B.n429 VSUBS 0.00881f
C506 B.n430 VSUBS 0.00881f
C507 B.n431 VSUBS 0.00881f
C508 B.n432 VSUBS 0.00881f
C509 B.n433 VSUBS 0.00881f
C510 B.n434 VSUBS 0.00881f
C511 B.n435 VSUBS 0.00881f
C512 B.n436 VSUBS 0.00881f
C513 B.n437 VSUBS 0.00881f
C514 B.n438 VSUBS 0.00881f
C515 B.n439 VSUBS 0.00881f
C516 B.n440 VSUBS 0.00881f
C517 B.n441 VSUBS 0.00881f
C518 B.n442 VSUBS 0.00881f
C519 B.n443 VSUBS 0.00881f
C520 B.n444 VSUBS 0.00881f
C521 B.n445 VSUBS 0.00881f
C522 B.n446 VSUBS 0.00881f
C523 B.n447 VSUBS 0.00881f
C524 B.n448 VSUBS 0.00881f
C525 B.n449 VSUBS 0.00881f
C526 B.n450 VSUBS 0.00881f
C527 B.n451 VSUBS 0.00881f
C528 B.n452 VSUBS 0.00881f
C529 B.n453 VSUBS 0.00881f
C530 B.n454 VSUBS 0.00881f
C531 B.n455 VSUBS 0.00881f
C532 B.n456 VSUBS 0.00881f
C533 B.n457 VSUBS 0.00881f
C534 B.n458 VSUBS 0.00881f
C535 B.n459 VSUBS 0.00881f
C536 B.n460 VSUBS 0.00881f
C537 B.n461 VSUBS 0.00881f
C538 B.n462 VSUBS 0.00881f
C539 B.n463 VSUBS 0.021226f
C540 B.n464 VSUBS 0.019712f
C541 B.n465 VSUBS 0.019712f
C542 B.n466 VSUBS 0.00881f
C543 B.n467 VSUBS 0.00881f
C544 B.n468 VSUBS 0.00881f
C545 B.n469 VSUBS 0.00881f
C546 B.n470 VSUBS 0.00881f
C547 B.n471 VSUBS 0.00881f
C548 B.n472 VSUBS 0.00881f
C549 B.n473 VSUBS 0.00881f
C550 B.n474 VSUBS 0.00881f
C551 B.n475 VSUBS 0.00881f
C552 B.n476 VSUBS 0.00881f
C553 B.n477 VSUBS 0.00881f
C554 B.n478 VSUBS 0.00881f
C555 B.n479 VSUBS 0.00881f
C556 B.n480 VSUBS 0.00881f
C557 B.n481 VSUBS 0.00881f
C558 B.n482 VSUBS 0.00881f
C559 B.n483 VSUBS 0.00881f
C560 B.n484 VSUBS 0.00881f
C561 B.n485 VSUBS 0.00881f
C562 B.n486 VSUBS 0.00881f
C563 B.n487 VSUBS 0.011496f
C564 B.n488 VSUBS 0.012246f
C565 B.n489 VSUBS 0.024353f
C566 VTAIL.t1 VSUBS 0.258514f
C567 VTAIL.t6 VSUBS 0.258514f
C568 VTAIL.n0 VSUBS 1.83967f
C569 VTAIL.n1 VSUBS 0.710599f
C570 VTAIL.n2 VSUBS 0.033572f
C571 VTAIL.n3 VSUBS 0.030319f
C572 VTAIL.n4 VSUBS 0.016292f
C573 VTAIL.n5 VSUBS 0.038508f
C574 VTAIL.n6 VSUBS 0.01725f
C575 VTAIL.n7 VSUBS 0.030319f
C576 VTAIL.n8 VSUBS 0.016292f
C577 VTAIL.n9 VSUBS 0.038508f
C578 VTAIL.n10 VSUBS 0.01725f
C579 VTAIL.n11 VSUBS 0.030319f
C580 VTAIL.n12 VSUBS 0.016292f
C581 VTAIL.n13 VSUBS 0.038508f
C582 VTAIL.n14 VSUBS 0.01725f
C583 VTAIL.n15 VSUBS 0.030319f
C584 VTAIL.n16 VSUBS 0.016292f
C585 VTAIL.n17 VSUBS 0.038508f
C586 VTAIL.n18 VSUBS 0.01725f
C587 VTAIL.n19 VSUBS 0.222201f
C588 VTAIL.t7 VSUBS 0.082871f
C589 VTAIL.n20 VSUBS 0.028881f
C590 VTAIL.n21 VSUBS 0.028968f
C591 VTAIL.n22 VSUBS 0.016292f
C592 VTAIL.n23 VSUBS 1.32888f
C593 VTAIL.n24 VSUBS 0.030319f
C594 VTAIL.n25 VSUBS 0.016292f
C595 VTAIL.n26 VSUBS 0.01725f
C596 VTAIL.n27 VSUBS 0.038508f
C597 VTAIL.n28 VSUBS 0.038508f
C598 VTAIL.n29 VSUBS 0.01725f
C599 VTAIL.n30 VSUBS 0.016292f
C600 VTAIL.n31 VSUBS 0.030319f
C601 VTAIL.n32 VSUBS 0.030319f
C602 VTAIL.n33 VSUBS 0.016292f
C603 VTAIL.n34 VSUBS 0.01725f
C604 VTAIL.n35 VSUBS 0.038508f
C605 VTAIL.n36 VSUBS 0.038508f
C606 VTAIL.n37 VSUBS 0.038508f
C607 VTAIL.n38 VSUBS 0.01725f
C608 VTAIL.n39 VSUBS 0.016292f
C609 VTAIL.n40 VSUBS 0.030319f
C610 VTAIL.n41 VSUBS 0.030319f
C611 VTAIL.n42 VSUBS 0.016292f
C612 VTAIL.n43 VSUBS 0.016771f
C613 VTAIL.n44 VSUBS 0.016771f
C614 VTAIL.n45 VSUBS 0.038508f
C615 VTAIL.n46 VSUBS 0.038508f
C616 VTAIL.n47 VSUBS 0.01725f
C617 VTAIL.n48 VSUBS 0.016292f
C618 VTAIL.n49 VSUBS 0.030319f
C619 VTAIL.n50 VSUBS 0.030319f
C620 VTAIL.n51 VSUBS 0.016292f
C621 VTAIL.n52 VSUBS 0.01725f
C622 VTAIL.n53 VSUBS 0.038508f
C623 VTAIL.n54 VSUBS 0.094105f
C624 VTAIL.n55 VSUBS 0.01725f
C625 VTAIL.n56 VSUBS 0.016292f
C626 VTAIL.n57 VSUBS 0.074636f
C627 VTAIL.n58 VSUBS 0.0475f
C628 VTAIL.n59 VSUBS 0.123215f
C629 VTAIL.n60 VSUBS 0.033572f
C630 VTAIL.n61 VSUBS 0.030319f
C631 VTAIL.n62 VSUBS 0.016292f
C632 VTAIL.n63 VSUBS 0.038508f
C633 VTAIL.n64 VSUBS 0.01725f
C634 VTAIL.n65 VSUBS 0.030319f
C635 VTAIL.n66 VSUBS 0.016292f
C636 VTAIL.n67 VSUBS 0.038508f
C637 VTAIL.n68 VSUBS 0.01725f
C638 VTAIL.n69 VSUBS 0.030319f
C639 VTAIL.n70 VSUBS 0.016292f
C640 VTAIL.n71 VSUBS 0.038508f
C641 VTAIL.n72 VSUBS 0.01725f
C642 VTAIL.n73 VSUBS 0.030319f
C643 VTAIL.n74 VSUBS 0.016292f
C644 VTAIL.n75 VSUBS 0.038508f
C645 VTAIL.n76 VSUBS 0.01725f
C646 VTAIL.n77 VSUBS 0.222201f
C647 VTAIL.t9 VSUBS 0.082871f
C648 VTAIL.n78 VSUBS 0.028881f
C649 VTAIL.n79 VSUBS 0.028968f
C650 VTAIL.n80 VSUBS 0.016292f
C651 VTAIL.n81 VSUBS 1.32888f
C652 VTAIL.n82 VSUBS 0.030319f
C653 VTAIL.n83 VSUBS 0.016292f
C654 VTAIL.n84 VSUBS 0.01725f
C655 VTAIL.n85 VSUBS 0.038508f
C656 VTAIL.n86 VSUBS 0.038508f
C657 VTAIL.n87 VSUBS 0.01725f
C658 VTAIL.n88 VSUBS 0.016292f
C659 VTAIL.n89 VSUBS 0.030319f
C660 VTAIL.n90 VSUBS 0.030319f
C661 VTAIL.n91 VSUBS 0.016292f
C662 VTAIL.n92 VSUBS 0.01725f
C663 VTAIL.n93 VSUBS 0.038508f
C664 VTAIL.n94 VSUBS 0.038508f
C665 VTAIL.n95 VSUBS 0.038508f
C666 VTAIL.n96 VSUBS 0.01725f
C667 VTAIL.n97 VSUBS 0.016292f
C668 VTAIL.n98 VSUBS 0.030319f
C669 VTAIL.n99 VSUBS 0.030319f
C670 VTAIL.n100 VSUBS 0.016292f
C671 VTAIL.n101 VSUBS 0.016771f
C672 VTAIL.n102 VSUBS 0.016771f
C673 VTAIL.n103 VSUBS 0.038508f
C674 VTAIL.n104 VSUBS 0.038508f
C675 VTAIL.n105 VSUBS 0.01725f
C676 VTAIL.n106 VSUBS 0.016292f
C677 VTAIL.n107 VSUBS 0.030319f
C678 VTAIL.n108 VSUBS 0.030319f
C679 VTAIL.n109 VSUBS 0.016292f
C680 VTAIL.n110 VSUBS 0.01725f
C681 VTAIL.n111 VSUBS 0.038508f
C682 VTAIL.n112 VSUBS 0.094105f
C683 VTAIL.n113 VSUBS 0.01725f
C684 VTAIL.n114 VSUBS 0.016292f
C685 VTAIL.n115 VSUBS 0.074636f
C686 VTAIL.n116 VSUBS 0.0475f
C687 VTAIL.n117 VSUBS 0.123215f
C688 VTAIL.t13 VSUBS 0.258514f
C689 VTAIL.t12 VSUBS 0.258514f
C690 VTAIL.n118 VSUBS 1.83967f
C691 VTAIL.n119 VSUBS 0.753761f
C692 VTAIL.n120 VSUBS 0.033572f
C693 VTAIL.n121 VSUBS 0.030319f
C694 VTAIL.n122 VSUBS 0.016292f
C695 VTAIL.n123 VSUBS 0.038508f
C696 VTAIL.n124 VSUBS 0.01725f
C697 VTAIL.n125 VSUBS 0.030319f
C698 VTAIL.n126 VSUBS 0.016292f
C699 VTAIL.n127 VSUBS 0.038508f
C700 VTAIL.n128 VSUBS 0.01725f
C701 VTAIL.n129 VSUBS 0.030319f
C702 VTAIL.n130 VSUBS 0.016292f
C703 VTAIL.n131 VSUBS 0.038508f
C704 VTAIL.n132 VSUBS 0.01725f
C705 VTAIL.n133 VSUBS 0.030319f
C706 VTAIL.n134 VSUBS 0.016292f
C707 VTAIL.n135 VSUBS 0.038508f
C708 VTAIL.n136 VSUBS 0.01725f
C709 VTAIL.n137 VSUBS 0.222201f
C710 VTAIL.t8 VSUBS 0.082871f
C711 VTAIL.n138 VSUBS 0.028881f
C712 VTAIL.n139 VSUBS 0.028968f
C713 VTAIL.n140 VSUBS 0.016292f
C714 VTAIL.n141 VSUBS 1.32888f
C715 VTAIL.n142 VSUBS 0.030319f
C716 VTAIL.n143 VSUBS 0.016292f
C717 VTAIL.n144 VSUBS 0.01725f
C718 VTAIL.n145 VSUBS 0.038508f
C719 VTAIL.n146 VSUBS 0.038508f
C720 VTAIL.n147 VSUBS 0.01725f
C721 VTAIL.n148 VSUBS 0.016292f
C722 VTAIL.n149 VSUBS 0.030319f
C723 VTAIL.n150 VSUBS 0.030319f
C724 VTAIL.n151 VSUBS 0.016292f
C725 VTAIL.n152 VSUBS 0.01725f
C726 VTAIL.n153 VSUBS 0.038508f
C727 VTAIL.n154 VSUBS 0.038508f
C728 VTAIL.n155 VSUBS 0.038508f
C729 VTAIL.n156 VSUBS 0.01725f
C730 VTAIL.n157 VSUBS 0.016292f
C731 VTAIL.n158 VSUBS 0.030319f
C732 VTAIL.n159 VSUBS 0.030319f
C733 VTAIL.n160 VSUBS 0.016292f
C734 VTAIL.n161 VSUBS 0.016771f
C735 VTAIL.n162 VSUBS 0.016771f
C736 VTAIL.n163 VSUBS 0.038508f
C737 VTAIL.n164 VSUBS 0.038508f
C738 VTAIL.n165 VSUBS 0.01725f
C739 VTAIL.n166 VSUBS 0.016292f
C740 VTAIL.n167 VSUBS 0.030319f
C741 VTAIL.n168 VSUBS 0.030319f
C742 VTAIL.n169 VSUBS 0.016292f
C743 VTAIL.n170 VSUBS 0.01725f
C744 VTAIL.n171 VSUBS 0.038508f
C745 VTAIL.n172 VSUBS 0.094105f
C746 VTAIL.n173 VSUBS 0.01725f
C747 VTAIL.n174 VSUBS 0.016292f
C748 VTAIL.n175 VSUBS 0.074636f
C749 VTAIL.n176 VSUBS 0.0475f
C750 VTAIL.n177 VSUBS 1.44672f
C751 VTAIL.n178 VSUBS 0.033572f
C752 VTAIL.n179 VSUBS 0.030319f
C753 VTAIL.n180 VSUBS 0.016292f
C754 VTAIL.n181 VSUBS 0.038508f
C755 VTAIL.n182 VSUBS 0.01725f
C756 VTAIL.n183 VSUBS 0.030319f
C757 VTAIL.n184 VSUBS 0.016292f
C758 VTAIL.n185 VSUBS 0.038508f
C759 VTAIL.n186 VSUBS 0.01725f
C760 VTAIL.n187 VSUBS 0.030319f
C761 VTAIL.n188 VSUBS 0.016292f
C762 VTAIL.n189 VSUBS 0.038508f
C763 VTAIL.n190 VSUBS 0.038508f
C764 VTAIL.n191 VSUBS 0.01725f
C765 VTAIL.n192 VSUBS 0.030319f
C766 VTAIL.n193 VSUBS 0.016292f
C767 VTAIL.n194 VSUBS 0.038508f
C768 VTAIL.n195 VSUBS 0.01725f
C769 VTAIL.n196 VSUBS 0.222201f
C770 VTAIL.t0 VSUBS 0.082871f
C771 VTAIL.n197 VSUBS 0.028881f
C772 VTAIL.n198 VSUBS 0.028968f
C773 VTAIL.n199 VSUBS 0.016292f
C774 VTAIL.n200 VSUBS 1.32888f
C775 VTAIL.n201 VSUBS 0.030319f
C776 VTAIL.n202 VSUBS 0.016292f
C777 VTAIL.n203 VSUBS 0.01725f
C778 VTAIL.n204 VSUBS 0.038508f
C779 VTAIL.n205 VSUBS 0.038508f
C780 VTAIL.n206 VSUBS 0.01725f
C781 VTAIL.n207 VSUBS 0.016292f
C782 VTAIL.n208 VSUBS 0.030319f
C783 VTAIL.n209 VSUBS 0.030319f
C784 VTAIL.n210 VSUBS 0.016292f
C785 VTAIL.n211 VSUBS 0.01725f
C786 VTAIL.n212 VSUBS 0.038508f
C787 VTAIL.n213 VSUBS 0.038508f
C788 VTAIL.n214 VSUBS 0.01725f
C789 VTAIL.n215 VSUBS 0.016292f
C790 VTAIL.n216 VSUBS 0.030319f
C791 VTAIL.n217 VSUBS 0.030319f
C792 VTAIL.n218 VSUBS 0.016292f
C793 VTAIL.n219 VSUBS 0.016771f
C794 VTAIL.n220 VSUBS 0.016771f
C795 VTAIL.n221 VSUBS 0.038508f
C796 VTAIL.n222 VSUBS 0.038508f
C797 VTAIL.n223 VSUBS 0.01725f
C798 VTAIL.n224 VSUBS 0.016292f
C799 VTAIL.n225 VSUBS 0.030319f
C800 VTAIL.n226 VSUBS 0.030319f
C801 VTAIL.n227 VSUBS 0.016292f
C802 VTAIL.n228 VSUBS 0.01725f
C803 VTAIL.n229 VSUBS 0.038508f
C804 VTAIL.n230 VSUBS 0.094105f
C805 VTAIL.n231 VSUBS 0.01725f
C806 VTAIL.n232 VSUBS 0.016292f
C807 VTAIL.n233 VSUBS 0.074636f
C808 VTAIL.n234 VSUBS 0.0475f
C809 VTAIL.n235 VSUBS 1.44672f
C810 VTAIL.t4 VSUBS 0.258514f
C811 VTAIL.t2 VSUBS 0.258514f
C812 VTAIL.n236 VSUBS 1.83968f
C813 VTAIL.n237 VSUBS 0.753749f
C814 VTAIL.n238 VSUBS 0.033572f
C815 VTAIL.n239 VSUBS 0.030319f
C816 VTAIL.n240 VSUBS 0.016292f
C817 VTAIL.n241 VSUBS 0.038508f
C818 VTAIL.n242 VSUBS 0.01725f
C819 VTAIL.n243 VSUBS 0.030319f
C820 VTAIL.n244 VSUBS 0.016292f
C821 VTAIL.n245 VSUBS 0.038508f
C822 VTAIL.n246 VSUBS 0.01725f
C823 VTAIL.n247 VSUBS 0.030319f
C824 VTAIL.n248 VSUBS 0.016292f
C825 VTAIL.n249 VSUBS 0.038508f
C826 VTAIL.n250 VSUBS 0.038508f
C827 VTAIL.n251 VSUBS 0.01725f
C828 VTAIL.n252 VSUBS 0.030319f
C829 VTAIL.n253 VSUBS 0.016292f
C830 VTAIL.n254 VSUBS 0.038508f
C831 VTAIL.n255 VSUBS 0.01725f
C832 VTAIL.n256 VSUBS 0.222201f
C833 VTAIL.t3 VSUBS 0.082871f
C834 VTAIL.n257 VSUBS 0.028881f
C835 VTAIL.n258 VSUBS 0.028968f
C836 VTAIL.n259 VSUBS 0.016292f
C837 VTAIL.n260 VSUBS 1.32888f
C838 VTAIL.n261 VSUBS 0.030319f
C839 VTAIL.n262 VSUBS 0.016292f
C840 VTAIL.n263 VSUBS 0.01725f
C841 VTAIL.n264 VSUBS 0.038508f
C842 VTAIL.n265 VSUBS 0.038508f
C843 VTAIL.n266 VSUBS 0.01725f
C844 VTAIL.n267 VSUBS 0.016292f
C845 VTAIL.n268 VSUBS 0.030319f
C846 VTAIL.n269 VSUBS 0.030319f
C847 VTAIL.n270 VSUBS 0.016292f
C848 VTAIL.n271 VSUBS 0.01725f
C849 VTAIL.n272 VSUBS 0.038508f
C850 VTAIL.n273 VSUBS 0.038508f
C851 VTAIL.n274 VSUBS 0.01725f
C852 VTAIL.n275 VSUBS 0.016292f
C853 VTAIL.n276 VSUBS 0.030319f
C854 VTAIL.n277 VSUBS 0.030319f
C855 VTAIL.n278 VSUBS 0.016292f
C856 VTAIL.n279 VSUBS 0.016771f
C857 VTAIL.n280 VSUBS 0.016771f
C858 VTAIL.n281 VSUBS 0.038508f
C859 VTAIL.n282 VSUBS 0.038508f
C860 VTAIL.n283 VSUBS 0.01725f
C861 VTAIL.n284 VSUBS 0.016292f
C862 VTAIL.n285 VSUBS 0.030319f
C863 VTAIL.n286 VSUBS 0.030319f
C864 VTAIL.n287 VSUBS 0.016292f
C865 VTAIL.n288 VSUBS 0.01725f
C866 VTAIL.n289 VSUBS 0.038508f
C867 VTAIL.n290 VSUBS 0.094105f
C868 VTAIL.n291 VSUBS 0.01725f
C869 VTAIL.n292 VSUBS 0.016292f
C870 VTAIL.n293 VSUBS 0.074636f
C871 VTAIL.n294 VSUBS 0.0475f
C872 VTAIL.n295 VSUBS 0.123215f
C873 VTAIL.n296 VSUBS 0.033572f
C874 VTAIL.n297 VSUBS 0.030319f
C875 VTAIL.n298 VSUBS 0.016292f
C876 VTAIL.n299 VSUBS 0.038508f
C877 VTAIL.n300 VSUBS 0.01725f
C878 VTAIL.n301 VSUBS 0.030319f
C879 VTAIL.n302 VSUBS 0.016292f
C880 VTAIL.n303 VSUBS 0.038508f
C881 VTAIL.n304 VSUBS 0.01725f
C882 VTAIL.n305 VSUBS 0.030319f
C883 VTAIL.n306 VSUBS 0.016292f
C884 VTAIL.n307 VSUBS 0.038508f
C885 VTAIL.n308 VSUBS 0.038508f
C886 VTAIL.n309 VSUBS 0.01725f
C887 VTAIL.n310 VSUBS 0.030319f
C888 VTAIL.n311 VSUBS 0.016292f
C889 VTAIL.n312 VSUBS 0.038508f
C890 VTAIL.n313 VSUBS 0.01725f
C891 VTAIL.n314 VSUBS 0.222201f
C892 VTAIL.t15 VSUBS 0.082871f
C893 VTAIL.n315 VSUBS 0.028881f
C894 VTAIL.n316 VSUBS 0.028968f
C895 VTAIL.n317 VSUBS 0.016292f
C896 VTAIL.n318 VSUBS 1.32888f
C897 VTAIL.n319 VSUBS 0.030319f
C898 VTAIL.n320 VSUBS 0.016292f
C899 VTAIL.n321 VSUBS 0.01725f
C900 VTAIL.n322 VSUBS 0.038508f
C901 VTAIL.n323 VSUBS 0.038508f
C902 VTAIL.n324 VSUBS 0.01725f
C903 VTAIL.n325 VSUBS 0.016292f
C904 VTAIL.n326 VSUBS 0.030319f
C905 VTAIL.n327 VSUBS 0.030319f
C906 VTAIL.n328 VSUBS 0.016292f
C907 VTAIL.n329 VSUBS 0.01725f
C908 VTAIL.n330 VSUBS 0.038508f
C909 VTAIL.n331 VSUBS 0.038508f
C910 VTAIL.n332 VSUBS 0.01725f
C911 VTAIL.n333 VSUBS 0.016292f
C912 VTAIL.n334 VSUBS 0.030319f
C913 VTAIL.n335 VSUBS 0.030319f
C914 VTAIL.n336 VSUBS 0.016292f
C915 VTAIL.n337 VSUBS 0.016771f
C916 VTAIL.n338 VSUBS 0.016771f
C917 VTAIL.n339 VSUBS 0.038508f
C918 VTAIL.n340 VSUBS 0.038508f
C919 VTAIL.n341 VSUBS 0.01725f
C920 VTAIL.n342 VSUBS 0.016292f
C921 VTAIL.n343 VSUBS 0.030319f
C922 VTAIL.n344 VSUBS 0.030319f
C923 VTAIL.n345 VSUBS 0.016292f
C924 VTAIL.n346 VSUBS 0.01725f
C925 VTAIL.n347 VSUBS 0.038508f
C926 VTAIL.n348 VSUBS 0.094105f
C927 VTAIL.n349 VSUBS 0.01725f
C928 VTAIL.n350 VSUBS 0.016292f
C929 VTAIL.n351 VSUBS 0.074636f
C930 VTAIL.n352 VSUBS 0.0475f
C931 VTAIL.n353 VSUBS 0.123215f
C932 VTAIL.t10 VSUBS 0.258514f
C933 VTAIL.t14 VSUBS 0.258514f
C934 VTAIL.n354 VSUBS 1.83968f
C935 VTAIL.n355 VSUBS 0.753749f
C936 VTAIL.n356 VSUBS 0.033572f
C937 VTAIL.n357 VSUBS 0.030319f
C938 VTAIL.n358 VSUBS 0.016292f
C939 VTAIL.n359 VSUBS 0.038508f
C940 VTAIL.n360 VSUBS 0.01725f
C941 VTAIL.n361 VSUBS 0.030319f
C942 VTAIL.n362 VSUBS 0.016292f
C943 VTAIL.n363 VSUBS 0.038508f
C944 VTAIL.n364 VSUBS 0.01725f
C945 VTAIL.n365 VSUBS 0.030319f
C946 VTAIL.n366 VSUBS 0.016292f
C947 VTAIL.n367 VSUBS 0.038508f
C948 VTAIL.n368 VSUBS 0.038508f
C949 VTAIL.n369 VSUBS 0.01725f
C950 VTAIL.n370 VSUBS 0.030319f
C951 VTAIL.n371 VSUBS 0.016292f
C952 VTAIL.n372 VSUBS 0.038508f
C953 VTAIL.n373 VSUBS 0.01725f
C954 VTAIL.n374 VSUBS 0.222201f
C955 VTAIL.t11 VSUBS 0.082871f
C956 VTAIL.n375 VSUBS 0.028881f
C957 VTAIL.n376 VSUBS 0.028968f
C958 VTAIL.n377 VSUBS 0.016292f
C959 VTAIL.n378 VSUBS 1.32888f
C960 VTAIL.n379 VSUBS 0.030319f
C961 VTAIL.n380 VSUBS 0.016292f
C962 VTAIL.n381 VSUBS 0.01725f
C963 VTAIL.n382 VSUBS 0.038508f
C964 VTAIL.n383 VSUBS 0.038508f
C965 VTAIL.n384 VSUBS 0.01725f
C966 VTAIL.n385 VSUBS 0.016292f
C967 VTAIL.n386 VSUBS 0.030319f
C968 VTAIL.n387 VSUBS 0.030319f
C969 VTAIL.n388 VSUBS 0.016292f
C970 VTAIL.n389 VSUBS 0.01725f
C971 VTAIL.n390 VSUBS 0.038508f
C972 VTAIL.n391 VSUBS 0.038508f
C973 VTAIL.n392 VSUBS 0.01725f
C974 VTAIL.n393 VSUBS 0.016292f
C975 VTAIL.n394 VSUBS 0.030319f
C976 VTAIL.n395 VSUBS 0.030319f
C977 VTAIL.n396 VSUBS 0.016292f
C978 VTAIL.n397 VSUBS 0.016771f
C979 VTAIL.n398 VSUBS 0.016771f
C980 VTAIL.n399 VSUBS 0.038508f
C981 VTAIL.n400 VSUBS 0.038508f
C982 VTAIL.n401 VSUBS 0.01725f
C983 VTAIL.n402 VSUBS 0.016292f
C984 VTAIL.n403 VSUBS 0.030319f
C985 VTAIL.n404 VSUBS 0.030319f
C986 VTAIL.n405 VSUBS 0.016292f
C987 VTAIL.n406 VSUBS 0.01725f
C988 VTAIL.n407 VSUBS 0.038508f
C989 VTAIL.n408 VSUBS 0.094105f
C990 VTAIL.n409 VSUBS 0.01725f
C991 VTAIL.n410 VSUBS 0.016292f
C992 VTAIL.n411 VSUBS 0.074636f
C993 VTAIL.n412 VSUBS 0.0475f
C994 VTAIL.n413 VSUBS 1.44672f
C995 VTAIL.n414 VSUBS 0.033572f
C996 VTAIL.n415 VSUBS 0.030319f
C997 VTAIL.n416 VSUBS 0.016292f
C998 VTAIL.n417 VSUBS 0.038508f
C999 VTAIL.n418 VSUBS 0.01725f
C1000 VTAIL.n419 VSUBS 0.030319f
C1001 VTAIL.n420 VSUBS 0.016292f
C1002 VTAIL.n421 VSUBS 0.038508f
C1003 VTAIL.n422 VSUBS 0.01725f
C1004 VTAIL.n423 VSUBS 0.030319f
C1005 VTAIL.n424 VSUBS 0.016292f
C1006 VTAIL.n425 VSUBS 0.038508f
C1007 VTAIL.n426 VSUBS 0.01725f
C1008 VTAIL.n427 VSUBS 0.030319f
C1009 VTAIL.n428 VSUBS 0.016292f
C1010 VTAIL.n429 VSUBS 0.038508f
C1011 VTAIL.n430 VSUBS 0.01725f
C1012 VTAIL.n431 VSUBS 0.222201f
C1013 VTAIL.t5 VSUBS 0.082871f
C1014 VTAIL.n432 VSUBS 0.028881f
C1015 VTAIL.n433 VSUBS 0.028968f
C1016 VTAIL.n434 VSUBS 0.016292f
C1017 VTAIL.n435 VSUBS 1.32888f
C1018 VTAIL.n436 VSUBS 0.030319f
C1019 VTAIL.n437 VSUBS 0.016292f
C1020 VTAIL.n438 VSUBS 0.01725f
C1021 VTAIL.n439 VSUBS 0.038508f
C1022 VTAIL.n440 VSUBS 0.038508f
C1023 VTAIL.n441 VSUBS 0.01725f
C1024 VTAIL.n442 VSUBS 0.016292f
C1025 VTAIL.n443 VSUBS 0.030319f
C1026 VTAIL.n444 VSUBS 0.030319f
C1027 VTAIL.n445 VSUBS 0.016292f
C1028 VTAIL.n446 VSUBS 0.01725f
C1029 VTAIL.n447 VSUBS 0.038508f
C1030 VTAIL.n448 VSUBS 0.038508f
C1031 VTAIL.n449 VSUBS 0.038508f
C1032 VTAIL.n450 VSUBS 0.01725f
C1033 VTAIL.n451 VSUBS 0.016292f
C1034 VTAIL.n452 VSUBS 0.030319f
C1035 VTAIL.n453 VSUBS 0.030319f
C1036 VTAIL.n454 VSUBS 0.016292f
C1037 VTAIL.n455 VSUBS 0.016771f
C1038 VTAIL.n456 VSUBS 0.016771f
C1039 VTAIL.n457 VSUBS 0.038508f
C1040 VTAIL.n458 VSUBS 0.038508f
C1041 VTAIL.n459 VSUBS 0.01725f
C1042 VTAIL.n460 VSUBS 0.016292f
C1043 VTAIL.n461 VSUBS 0.030319f
C1044 VTAIL.n462 VSUBS 0.030319f
C1045 VTAIL.n463 VSUBS 0.016292f
C1046 VTAIL.n464 VSUBS 0.01725f
C1047 VTAIL.n465 VSUBS 0.038508f
C1048 VTAIL.n466 VSUBS 0.094105f
C1049 VTAIL.n467 VSUBS 0.01725f
C1050 VTAIL.n468 VSUBS 0.016292f
C1051 VTAIL.n469 VSUBS 0.074636f
C1052 VTAIL.n470 VSUBS 0.0475f
C1053 VTAIL.n471 VSUBS 1.44103f
C1054 VDD1.t7 VSUBS 0.299337f
C1055 VDD1.t1 VSUBS 0.299337f
C1056 VDD1.n0 VSUBS 2.30433f
C1057 VDD1.t5 VSUBS 0.299337f
C1058 VDD1.t2 VSUBS 0.299337f
C1059 VDD1.n1 VSUBS 2.30322f
C1060 VDD1.t4 VSUBS 0.299337f
C1061 VDD1.t6 VSUBS 0.299337f
C1062 VDD1.n2 VSUBS 2.30322f
C1063 VDD1.n3 VSUBS 3.34606f
C1064 VDD1.t3 VSUBS 0.299337f
C1065 VDD1.t0 VSUBS 0.299337f
C1066 VDD1.n4 VSUBS 2.3014f
C1067 VDD1.n5 VSUBS 3.25171f
C1068 VP.n0 VSUBS 0.074116f
C1069 VP.t3 VSUBS 0.565654f
C1070 VP.t2 VSUBS 0.565654f
C1071 VP.t7 VSUBS 0.576183f
C1072 VP.n1 VSUBS 0.170509f
C1073 VP.t1 VSUBS 0.565654f
C1074 VP.t5 VSUBS 0.565654f
C1075 VP.t0 VSUBS 0.576183f
C1076 VP.n2 VSUBS 0.255596f
C1077 VP.n3 VSUBS 0.232285f
C1078 VP.n4 VSUBS 0.028242f
C1079 VP.n5 VSUBS 0.232285f
C1080 VP.t4 VSUBS 0.576183f
C1081 VP.n6 VSUBS 0.255483f
C1082 VP.n7 VSUBS 2.70786f
C1083 VP.n8 VSUBS 2.77599f
C1084 VP.n9 VSUBS 0.255483f
C1085 VP.n10 VSUBS 0.232285f
C1086 VP.n11 VSUBS 0.028242f
C1087 VP.n12 VSUBS 0.232285f
C1088 VP.t6 VSUBS 0.576183f
C1089 VP.n13 VSUBS 0.255483f
C1090 VP.n14 VSUBS 0.057437f
.ends

