* NGSPICE file created from diff_pair_sample_0522.ext - technology: sky130A

.subckt diff_pair_sample_0522 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1758_n1356# sky130_fd_pr__pfet_01v8 ad=0.7566 pd=4.66 as=0 ps=0 w=1.94 l=1.64
X1 VDD2.t1 VN.t0 VTAIL.t2 w_n1758_n1356# sky130_fd_pr__pfet_01v8 ad=0.7566 pd=4.66 as=0.7566 ps=4.66 w=1.94 l=1.64
X2 B.t8 B.t6 B.t7 w_n1758_n1356# sky130_fd_pr__pfet_01v8 ad=0.7566 pd=4.66 as=0 ps=0 w=1.94 l=1.64
X3 VDD1.t1 VP.t0 VTAIL.t1 w_n1758_n1356# sky130_fd_pr__pfet_01v8 ad=0.7566 pd=4.66 as=0.7566 ps=4.66 w=1.94 l=1.64
X4 VDD1.t0 VP.t1 VTAIL.t0 w_n1758_n1356# sky130_fd_pr__pfet_01v8 ad=0.7566 pd=4.66 as=0.7566 ps=4.66 w=1.94 l=1.64
X5 VDD2.t0 VN.t1 VTAIL.t3 w_n1758_n1356# sky130_fd_pr__pfet_01v8 ad=0.7566 pd=4.66 as=0.7566 ps=4.66 w=1.94 l=1.64
X6 B.t5 B.t3 B.t4 w_n1758_n1356# sky130_fd_pr__pfet_01v8 ad=0.7566 pd=4.66 as=0 ps=0 w=1.94 l=1.64
X7 B.t2 B.t0 B.t1 w_n1758_n1356# sky130_fd_pr__pfet_01v8 ad=0.7566 pd=4.66 as=0 ps=0 w=1.94 l=1.64
R0 B.n163 B.n162 585
R1 B.n161 B.n54 585
R2 B.n160 B.n159 585
R3 B.n158 B.n55 585
R4 B.n157 B.n156 585
R5 B.n155 B.n56 585
R6 B.n154 B.n153 585
R7 B.n152 B.n57 585
R8 B.n151 B.n150 585
R9 B.n149 B.n58 585
R10 B.n148 B.n147 585
R11 B.n146 B.n59 585
R12 B.n145 B.n144 585
R13 B.n140 B.n60 585
R14 B.n139 B.n138 585
R15 B.n137 B.n61 585
R16 B.n136 B.n135 585
R17 B.n134 B.n62 585
R18 B.n133 B.n132 585
R19 B.n131 B.n63 585
R20 B.n130 B.n129 585
R21 B.n128 B.n64 585
R22 B.n126 B.n125 585
R23 B.n124 B.n67 585
R24 B.n123 B.n122 585
R25 B.n121 B.n68 585
R26 B.n120 B.n119 585
R27 B.n118 B.n69 585
R28 B.n117 B.n116 585
R29 B.n115 B.n70 585
R30 B.n114 B.n113 585
R31 B.n112 B.n71 585
R32 B.n111 B.n110 585
R33 B.n109 B.n72 585
R34 B.n164 B.n53 585
R35 B.n166 B.n165 585
R36 B.n167 B.n52 585
R37 B.n169 B.n168 585
R38 B.n170 B.n51 585
R39 B.n172 B.n171 585
R40 B.n173 B.n50 585
R41 B.n175 B.n174 585
R42 B.n176 B.n49 585
R43 B.n178 B.n177 585
R44 B.n179 B.n48 585
R45 B.n181 B.n180 585
R46 B.n182 B.n47 585
R47 B.n184 B.n183 585
R48 B.n185 B.n46 585
R49 B.n187 B.n186 585
R50 B.n188 B.n45 585
R51 B.n190 B.n189 585
R52 B.n191 B.n44 585
R53 B.n193 B.n192 585
R54 B.n194 B.n43 585
R55 B.n196 B.n195 585
R56 B.n197 B.n42 585
R57 B.n199 B.n198 585
R58 B.n200 B.n41 585
R59 B.n202 B.n201 585
R60 B.n203 B.n40 585
R61 B.n205 B.n204 585
R62 B.n206 B.n39 585
R63 B.n208 B.n207 585
R64 B.n209 B.n38 585
R65 B.n211 B.n210 585
R66 B.n212 B.n37 585
R67 B.n214 B.n213 585
R68 B.n215 B.n36 585
R69 B.n217 B.n216 585
R70 B.n218 B.n35 585
R71 B.n220 B.n219 585
R72 B.n221 B.n34 585
R73 B.n223 B.n222 585
R74 B.n275 B.n274 585
R75 B.n273 B.n12 585
R76 B.n272 B.n271 585
R77 B.n270 B.n13 585
R78 B.n269 B.n268 585
R79 B.n267 B.n14 585
R80 B.n266 B.n265 585
R81 B.n264 B.n15 585
R82 B.n263 B.n262 585
R83 B.n261 B.n16 585
R84 B.n260 B.n259 585
R85 B.n258 B.n17 585
R86 B.n256 B.n255 585
R87 B.n254 B.n20 585
R88 B.n253 B.n252 585
R89 B.n251 B.n21 585
R90 B.n250 B.n249 585
R91 B.n248 B.n22 585
R92 B.n247 B.n246 585
R93 B.n245 B.n23 585
R94 B.n244 B.n243 585
R95 B.n242 B.n24 585
R96 B.n241 B.n240 585
R97 B.n239 B.n25 585
R98 B.n238 B.n237 585
R99 B.n236 B.n29 585
R100 B.n235 B.n234 585
R101 B.n233 B.n30 585
R102 B.n232 B.n231 585
R103 B.n230 B.n31 585
R104 B.n229 B.n228 585
R105 B.n227 B.n32 585
R106 B.n226 B.n225 585
R107 B.n224 B.n33 585
R108 B.n276 B.n11 585
R109 B.n278 B.n277 585
R110 B.n279 B.n10 585
R111 B.n281 B.n280 585
R112 B.n282 B.n9 585
R113 B.n284 B.n283 585
R114 B.n285 B.n8 585
R115 B.n287 B.n286 585
R116 B.n288 B.n7 585
R117 B.n290 B.n289 585
R118 B.n291 B.n6 585
R119 B.n293 B.n292 585
R120 B.n294 B.n5 585
R121 B.n296 B.n295 585
R122 B.n297 B.n4 585
R123 B.n299 B.n298 585
R124 B.n300 B.n3 585
R125 B.n302 B.n301 585
R126 B.n303 B.n0 585
R127 B.n2 B.n1 585
R128 B.n82 B.n81 585
R129 B.n84 B.n83 585
R130 B.n85 B.n80 585
R131 B.n87 B.n86 585
R132 B.n88 B.n79 585
R133 B.n90 B.n89 585
R134 B.n91 B.n78 585
R135 B.n93 B.n92 585
R136 B.n94 B.n77 585
R137 B.n96 B.n95 585
R138 B.n97 B.n76 585
R139 B.n99 B.n98 585
R140 B.n100 B.n75 585
R141 B.n102 B.n101 585
R142 B.n103 B.n74 585
R143 B.n105 B.n104 585
R144 B.n106 B.n73 585
R145 B.n108 B.n107 585
R146 B.n107 B.n72 502.111
R147 B.n164 B.n163 502.111
R148 B.n224 B.n223 502.111
R149 B.n274 B.n11 502.111
R150 B.n141 B.t7 285.38
R151 B.n26 B.t11 285.38
R152 B.n65 B.t4 285.38
R153 B.n18 B.t2 285.38
R154 B.n305 B.n304 256.663
R155 B.n142 B.t8 247.173
R156 B.n27 B.t10 247.173
R157 B.n66 B.t5 247.173
R158 B.n19 B.t1 247.173
R159 B.n304 B.n303 235.042
R160 B.n304 B.n2 235.042
R161 B.n65 B.t3 234.435
R162 B.n141 B.t6 234.435
R163 B.n26 B.t9 234.435
R164 B.n18 B.t0 234.435
R165 B.n111 B.n72 163.367
R166 B.n112 B.n111 163.367
R167 B.n113 B.n112 163.367
R168 B.n113 B.n70 163.367
R169 B.n117 B.n70 163.367
R170 B.n118 B.n117 163.367
R171 B.n119 B.n118 163.367
R172 B.n119 B.n68 163.367
R173 B.n123 B.n68 163.367
R174 B.n124 B.n123 163.367
R175 B.n125 B.n124 163.367
R176 B.n125 B.n64 163.367
R177 B.n130 B.n64 163.367
R178 B.n131 B.n130 163.367
R179 B.n132 B.n131 163.367
R180 B.n132 B.n62 163.367
R181 B.n136 B.n62 163.367
R182 B.n137 B.n136 163.367
R183 B.n138 B.n137 163.367
R184 B.n138 B.n60 163.367
R185 B.n145 B.n60 163.367
R186 B.n146 B.n145 163.367
R187 B.n147 B.n146 163.367
R188 B.n147 B.n58 163.367
R189 B.n151 B.n58 163.367
R190 B.n152 B.n151 163.367
R191 B.n153 B.n152 163.367
R192 B.n153 B.n56 163.367
R193 B.n157 B.n56 163.367
R194 B.n158 B.n157 163.367
R195 B.n159 B.n158 163.367
R196 B.n159 B.n54 163.367
R197 B.n163 B.n54 163.367
R198 B.n223 B.n34 163.367
R199 B.n219 B.n34 163.367
R200 B.n219 B.n218 163.367
R201 B.n218 B.n217 163.367
R202 B.n217 B.n36 163.367
R203 B.n213 B.n36 163.367
R204 B.n213 B.n212 163.367
R205 B.n212 B.n211 163.367
R206 B.n211 B.n38 163.367
R207 B.n207 B.n38 163.367
R208 B.n207 B.n206 163.367
R209 B.n206 B.n205 163.367
R210 B.n205 B.n40 163.367
R211 B.n201 B.n40 163.367
R212 B.n201 B.n200 163.367
R213 B.n200 B.n199 163.367
R214 B.n199 B.n42 163.367
R215 B.n195 B.n42 163.367
R216 B.n195 B.n194 163.367
R217 B.n194 B.n193 163.367
R218 B.n193 B.n44 163.367
R219 B.n189 B.n44 163.367
R220 B.n189 B.n188 163.367
R221 B.n188 B.n187 163.367
R222 B.n187 B.n46 163.367
R223 B.n183 B.n46 163.367
R224 B.n183 B.n182 163.367
R225 B.n182 B.n181 163.367
R226 B.n181 B.n48 163.367
R227 B.n177 B.n48 163.367
R228 B.n177 B.n176 163.367
R229 B.n176 B.n175 163.367
R230 B.n175 B.n50 163.367
R231 B.n171 B.n50 163.367
R232 B.n171 B.n170 163.367
R233 B.n170 B.n169 163.367
R234 B.n169 B.n52 163.367
R235 B.n165 B.n52 163.367
R236 B.n165 B.n164 163.367
R237 B.n274 B.n273 163.367
R238 B.n273 B.n272 163.367
R239 B.n272 B.n13 163.367
R240 B.n268 B.n13 163.367
R241 B.n268 B.n267 163.367
R242 B.n267 B.n266 163.367
R243 B.n266 B.n15 163.367
R244 B.n262 B.n15 163.367
R245 B.n262 B.n261 163.367
R246 B.n261 B.n260 163.367
R247 B.n260 B.n17 163.367
R248 B.n255 B.n17 163.367
R249 B.n255 B.n254 163.367
R250 B.n254 B.n253 163.367
R251 B.n253 B.n21 163.367
R252 B.n249 B.n21 163.367
R253 B.n249 B.n248 163.367
R254 B.n248 B.n247 163.367
R255 B.n247 B.n23 163.367
R256 B.n243 B.n23 163.367
R257 B.n243 B.n242 163.367
R258 B.n242 B.n241 163.367
R259 B.n241 B.n25 163.367
R260 B.n237 B.n25 163.367
R261 B.n237 B.n236 163.367
R262 B.n236 B.n235 163.367
R263 B.n235 B.n30 163.367
R264 B.n231 B.n30 163.367
R265 B.n231 B.n230 163.367
R266 B.n230 B.n229 163.367
R267 B.n229 B.n32 163.367
R268 B.n225 B.n32 163.367
R269 B.n225 B.n224 163.367
R270 B.n278 B.n11 163.367
R271 B.n279 B.n278 163.367
R272 B.n280 B.n279 163.367
R273 B.n280 B.n9 163.367
R274 B.n284 B.n9 163.367
R275 B.n285 B.n284 163.367
R276 B.n286 B.n285 163.367
R277 B.n286 B.n7 163.367
R278 B.n290 B.n7 163.367
R279 B.n291 B.n290 163.367
R280 B.n292 B.n291 163.367
R281 B.n292 B.n5 163.367
R282 B.n296 B.n5 163.367
R283 B.n297 B.n296 163.367
R284 B.n298 B.n297 163.367
R285 B.n298 B.n3 163.367
R286 B.n302 B.n3 163.367
R287 B.n303 B.n302 163.367
R288 B.n82 B.n2 163.367
R289 B.n83 B.n82 163.367
R290 B.n83 B.n80 163.367
R291 B.n87 B.n80 163.367
R292 B.n88 B.n87 163.367
R293 B.n89 B.n88 163.367
R294 B.n89 B.n78 163.367
R295 B.n93 B.n78 163.367
R296 B.n94 B.n93 163.367
R297 B.n95 B.n94 163.367
R298 B.n95 B.n76 163.367
R299 B.n99 B.n76 163.367
R300 B.n100 B.n99 163.367
R301 B.n101 B.n100 163.367
R302 B.n101 B.n74 163.367
R303 B.n105 B.n74 163.367
R304 B.n106 B.n105 163.367
R305 B.n107 B.n106 163.367
R306 B.n127 B.n66 59.5399
R307 B.n143 B.n142 59.5399
R308 B.n28 B.n27 59.5399
R309 B.n257 B.n19 59.5399
R310 B.n66 B.n65 38.2066
R311 B.n142 B.n141 38.2066
R312 B.n27 B.n26 38.2066
R313 B.n19 B.n18 38.2066
R314 B.n276 B.n275 32.6249
R315 B.n222 B.n33 32.6249
R316 B.n162 B.n53 32.6249
R317 B.n109 B.n108 32.6249
R318 B B.n305 18.0485
R319 B.n277 B.n276 10.6151
R320 B.n277 B.n10 10.6151
R321 B.n281 B.n10 10.6151
R322 B.n282 B.n281 10.6151
R323 B.n283 B.n282 10.6151
R324 B.n283 B.n8 10.6151
R325 B.n287 B.n8 10.6151
R326 B.n288 B.n287 10.6151
R327 B.n289 B.n288 10.6151
R328 B.n289 B.n6 10.6151
R329 B.n293 B.n6 10.6151
R330 B.n294 B.n293 10.6151
R331 B.n295 B.n294 10.6151
R332 B.n295 B.n4 10.6151
R333 B.n299 B.n4 10.6151
R334 B.n300 B.n299 10.6151
R335 B.n301 B.n300 10.6151
R336 B.n301 B.n0 10.6151
R337 B.n275 B.n12 10.6151
R338 B.n271 B.n12 10.6151
R339 B.n271 B.n270 10.6151
R340 B.n270 B.n269 10.6151
R341 B.n269 B.n14 10.6151
R342 B.n265 B.n14 10.6151
R343 B.n265 B.n264 10.6151
R344 B.n264 B.n263 10.6151
R345 B.n263 B.n16 10.6151
R346 B.n259 B.n16 10.6151
R347 B.n259 B.n258 10.6151
R348 B.n256 B.n20 10.6151
R349 B.n252 B.n20 10.6151
R350 B.n252 B.n251 10.6151
R351 B.n251 B.n250 10.6151
R352 B.n250 B.n22 10.6151
R353 B.n246 B.n22 10.6151
R354 B.n246 B.n245 10.6151
R355 B.n245 B.n244 10.6151
R356 B.n244 B.n24 10.6151
R357 B.n240 B.n239 10.6151
R358 B.n239 B.n238 10.6151
R359 B.n238 B.n29 10.6151
R360 B.n234 B.n29 10.6151
R361 B.n234 B.n233 10.6151
R362 B.n233 B.n232 10.6151
R363 B.n232 B.n31 10.6151
R364 B.n228 B.n31 10.6151
R365 B.n228 B.n227 10.6151
R366 B.n227 B.n226 10.6151
R367 B.n226 B.n33 10.6151
R368 B.n222 B.n221 10.6151
R369 B.n221 B.n220 10.6151
R370 B.n220 B.n35 10.6151
R371 B.n216 B.n35 10.6151
R372 B.n216 B.n215 10.6151
R373 B.n215 B.n214 10.6151
R374 B.n214 B.n37 10.6151
R375 B.n210 B.n37 10.6151
R376 B.n210 B.n209 10.6151
R377 B.n209 B.n208 10.6151
R378 B.n208 B.n39 10.6151
R379 B.n204 B.n39 10.6151
R380 B.n204 B.n203 10.6151
R381 B.n203 B.n202 10.6151
R382 B.n202 B.n41 10.6151
R383 B.n198 B.n41 10.6151
R384 B.n198 B.n197 10.6151
R385 B.n197 B.n196 10.6151
R386 B.n196 B.n43 10.6151
R387 B.n192 B.n43 10.6151
R388 B.n192 B.n191 10.6151
R389 B.n191 B.n190 10.6151
R390 B.n190 B.n45 10.6151
R391 B.n186 B.n45 10.6151
R392 B.n186 B.n185 10.6151
R393 B.n185 B.n184 10.6151
R394 B.n184 B.n47 10.6151
R395 B.n180 B.n47 10.6151
R396 B.n180 B.n179 10.6151
R397 B.n179 B.n178 10.6151
R398 B.n178 B.n49 10.6151
R399 B.n174 B.n49 10.6151
R400 B.n174 B.n173 10.6151
R401 B.n173 B.n172 10.6151
R402 B.n172 B.n51 10.6151
R403 B.n168 B.n51 10.6151
R404 B.n168 B.n167 10.6151
R405 B.n167 B.n166 10.6151
R406 B.n166 B.n53 10.6151
R407 B.n81 B.n1 10.6151
R408 B.n84 B.n81 10.6151
R409 B.n85 B.n84 10.6151
R410 B.n86 B.n85 10.6151
R411 B.n86 B.n79 10.6151
R412 B.n90 B.n79 10.6151
R413 B.n91 B.n90 10.6151
R414 B.n92 B.n91 10.6151
R415 B.n92 B.n77 10.6151
R416 B.n96 B.n77 10.6151
R417 B.n97 B.n96 10.6151
R418 B.n98 B.n97 10.6151
R419 B.n98 B.n75 10.6151
R420 B.n102 B.n75 10.6151
R421 B.n103 B.n102 10.6151
R422 B.n104 B.n103 10.6151
R423 B.n104 B.n73 10.6151
R424 B.n108 B.n73 10.6151
R425 B.n110 B.n109 10.6151
R426 B.n110 B.n71 10.6151
R427 B.n114 B.n71 10.6151
R428 B.n115 B.n114 10.6151
R429 B.n116 B.n115 10.6151
R430 B.n116 B.n69 10.6151
R431 B.n120 B.n69 10.6151
R432 B.n121 B.n120 10.6151
R433 B.n122 B.n121 10.6151
R434 B.n122 B.n67 10.6151
R435 B.n126 B.n67 10.6151
R436 B.n129 B.n128 10.6151
R437 B.n129 B.n63 10.6151
R438 B.n133 B.n63 10.6151
R439 B.n134 B.n133 10.6151
R440 B.n135 B.n134 10.6151
R441 B.n135 B.n61 10.6151
R442 B.n139 B.n61 10.6151
R443 B.n140 B.n139 10.6151
R444 B.n144 B.n140 10.6151
R445 B.n148 B.n59 10.6151
R446 B.n149 B.n148 10.6151
R447 B.n150 B.n149 10.6151
R448 B.n150 B.n57 10.6151
R449 B.n154 B.n57 10.6151
R450 B.n155 B.n154 10.6151
R451 B.n156 B.n155 10.6151
R452 B.n156 B.n55 10.6151
R453 B.n160 B.n55 10.6151
R454 B.n161 B.n160 10.6151
R455 B.n162 B.n161 10.6151
R456 B.n258 B.n257 9.36635
R457 B.n240 B.n28 9.36635
R458 B.n127 B.n126 9.36635
R459 B.n143 B.n59 9.36635
R460 B.n305 B.n0 8.11757
R461 B.n305 B.n1 8.11757
R462 B.n257 B.n256 1.24928
R463 B.n28 B.n24 1.24928
R464 B.n128 B.n127 1.24928
R465 B.n144 B.n143 1.24928
R466 VN VN.t1 122.076
R467 VN VN.t0 87.6361
R468 VTAIL.n26 VTAIL.n24 756.745
R469 VTAIL.n2 VTAIL.n0 756.745
R470 VTAIL.n18 VTAIL.n16 756.745
R471 VTAIL.n10 VTAIL.n8 756.745
R472 VTAIL.n27 VTAIL.n26 585
R473 VTAIL.n3 VTAIL.n2 585
R474 VTAIL.n19 VTAIL.n18 585
R475 VTAIL.n11 VTAIL.n10 585
R476 VTAIL.t2 VTAIL.n25 417.779
R477 VTAIL.t0 VTAIL.n1 417.779
R478 VTAIL.t1 VTAIL.n17 417.779
R479 VTAIL.t3 VTAIL.n9 417.779
R480 VTAIL.n26 VTAIL.t2 85.8723
R481 VTAIL.n2 VTAIL.t0 85.8723
R482 VTAIL.n18 VTAIL.t1 85.8723
R483 VTAIL.n10 VTAIL.t3 85.8723
R484 VTAIL.n31 VTAIL.n30 30.246
R485 VTAIL.n7 VTAIL.n6 30.246
R486 VTAIL.n23 VTAIL.n22 30.246
R487 VTAIL.n15 VTAIL.n14 30.246
R488 VTAIL.n15 VTAIL.n7 17.4358
R489 VTAIL.n31 VTAIL.n23 15.7376
R490 VTAIL.n27 VTAIL.n25 9.84608
R491 VTAIL.n3 VTAIL.n1 9.84608
R492 VTAIL.n19 VTAIL.n17 9.84608
R493 VTAIL.n11 VTAIL.n9 9.84608
R494 VTAIL.n30 VTAIL.n29 9.45567
R495 VTAIL.n6 VTAIL.n5 9.45567
R496 VTAIL.n22 VTAIL.n21 9.45567
R497 VTAIL.n14 VTAIL.n13 9.45567
R498 VTAIL.n29 VTAIL.n28 9.3005
R499 VTAIL.n5 VTAIL.n4 9.3005
R500 VTAIL.n21 VTAIL.n20 9.3005
R501 VTAIL.n13 VTAIL.n12 9.3005
R502 VTAIL.n30 VTAIL.n24 8.14595
R503 VTAIL.n6 VTAIL.n0 8.14595
R504 VTAIL.n22 VTAIL.n16 8.14595
R505 VTAIL.n14 VTAIL.n8 8.14595
R506 VTAIL.n28 VTAIL.n27 7.3702
R507 VTAIL.n4 VTAIL.n3 7.3702
R508 VTAIL.n20 VTAIL.n19 7.3702
R509 VTAIL.n12 VTAIL.n11 7.3702
R510 VTAIL.n28 VTAIL.n24 5.81868
R511 VTAIL.n4 VTAIL.n0 5.81868
R512 VTAIL.n20 VTAIL.n16 5.81868
R513 VTAIL.n12 VTAIL.n8 5.81868
R514 VTAIL.n13 VTAIL.n9 3.32369
R515 VTAIL.n29 VTAIL.n25 3.32369
R516 VTAIL.n5 VTAIL.n1 3.32369
R517 VTAIL.n21 VTAIL.n17 3.32369
R518 VTAIL.n23 VTAIL.n15 1.31947
R519 VTAIL VTAIL.n7 0.953086
R520 VTAIL VTAIL.n31 0.366879
R521 VDD2.n9 VDD2.n7 756.745
R522 VDD2.n2 VDD2.n0 756.745
R523 VDD2.n10 VDD2.n9 585
R524 VDD2.n3 VDD2.n2 585
R525 VDD2.t1 VDD2.n1 417.779
R526 VDD2.t0 VDD2.n8 417.779
R527 VDD2.n9 VDD2.t0 85.8723
R528 VDD2.n2 VDD2.t1 85.8723
R529 VDD2.n14 VDD2.n6 75.6532
R530 VDD2.n14 VDD2.n13 46.9247
R531 VDD2.n10 VDD2.n8 9.84608
R532 VDD2.n3 VDD2.n1 9.84608
R533 VDD2.n13 VDD2.n12 9.45567
R534 VDD2.n6 VDD2.n5 9.45567
R535 VDD2.n12 VDD2.n11 9.3005
R536 VDD2.n5 VDD2.n4 9.3005
R537 VDD2.n13 VDD2.n7 8.14595
R538 VDD2.n6 VDD2.n0 8.14595
R539 VDD2.n11 VDD2.n10 7.3702
R540 VDD2.n4 VDD2.n3 7.3702
R541 VDD2.n11 VDD2.n7 5.81868
R542 VDD2.n4 VDD2.n0 5.81868
R543 VDD2.n12 VDD2.n8 3.32369
R544 VDD2.n5 VDD2.n1 3.32369
R545 VDD2 VDD2.n14 0.483259
R546 VP.n0 VP.t0 121.885
R547 VP.n0 VP.t1 87.3949
R548 VP VP.n0 0.241678
R549 VDD1.n2 VDD1.n0 756.745
R550 VDD1.n9 VDD1.n7 756.745
R551 VDD1.n3 VDD1.n2 585
R552 VDD1.n10 VDD1.n9 585
R553 VDD1.t0 VDD1.n8 417.779
R554 VDD1.t1 VDD1.n1 417.779
R555 VDD1.n2 VDD1.t1 85.8723
R556 VDD1.n9 VDD1.t0 85.8723
R557 VDD1 VDD1.n13 76.6025
R558 VDD1 VDD1.n6 47.4075
R559 VDD1.n3 VDD1.n1 9.84608
R560 VDD1.n10 VDD1.n8 9.84608
R561 VDD1.n6 VDD1.n5 9.45567
R562 VDD1.n13 VDD1.n12 9.45567
R563 VDD1.n5 VDD1.n4 9.3005
R564 VDD1.n12 VDD1.n11 9.3005
R565 VDD1.n6 VDD1.n0 8.14595
R566 VDD1.n13 VDD1.n7 8.14595
R567 VDD1.n4 VDD1.n3 7.3702
R568 VDD1.n11 VDD1.n10 7.3702
R569 VDD1.n4 VDD1.n0 5.81868
R570 VDD1.n11 VDD1.n7 5.81868
R571 VDD1.n5 VDD1.n1 3.32369
R572 VDD1.n12 VDD1.n8 3.32369
C0 w_n1758_n1356# VN 2.13134f
C1 VDD2 VTAIL 2.16342f
C2 VDD1 VTAIL 2.11717f
C3 w_n1758_n1356# VDD2 0.966108f
C4 w_n1758_n1356# VDD1 0.952478f
C5 VP VTAIL 0.802403f
C6 VDD2 VN 0.620885f
C7 VN VDD1 0.154402f
C8 w_n1758_n1356# VP 2.34842f
C9 VN VP 3.15054f
C10 VDD2 VDD1 0.560209f
C11 B VTAIL 1.08747f
C12 VDD2 VP 0.299209f
C13 VDD1 VP 0.764157f
C14 B w_n1758_n1356# 4.95558f
C15 B VN 0.745955f
C16 w_n1758_n1356# VTAIL 1.23238f
C17 B VDD2 0.818566f
C18 B VDD1 0.796704f
C19 VN VTAIL 0.788249f
C20 B VP 1.10609f
C21 VDD2 VSUBS 0.467437f
C22 VDD1 VSUBS 1.842381f
C23 VTAIL VSUBS 0.330899f
C24 VN VSUBS 4.88481f
C25 VP VSUBS 0.935083f
C26 B VSUBS 2.213434f
C27 w_n1758_n1356# VSUBS 30.4415f
C28 VDD1.n0 VSUBS 0.017684f
C29 VDD1.n1 VSUBS 0.045676f
C30 VDD1.t1 VSUBS 0.045788f
C31 VDD1.n2 VSUBS 0.044439f
C32 VDD1.n3 VSUBS 0.01328f
C33 VDD1.n4 VSUBS 0.008615f
C34 VDD1.n5 VSUBS 0.107102f
C35 VDD1.n6 VSUBS 0.036493f
C36 VDD1.n7 VSUBS 0.017684f
C37 VDD1.n8 VSUBS 0.045676f
C38 VDD1.t0 VSUBS 0.045788f
C39 VDD1.n9 VSUBS 0.044439f
C40 VDD1.n10 VSUBS 0.01328f
C41 VDD1.n11 VSUBS 0.008615f
C42 VDD1.n12 VSUBS 0.107102f
C43 VDD1.n13 VSUBS 0.26073f
C44 VP.t0 VSUBS 1.31496f
C45 VP.t1 VSUBS 0.760577f
C46 VP.n0 VSUBS 3.34363f
C47 VDD2.n0 VSUBS 0.019064f
C48 VDD2.n1 VSUBS 0.049239f
C49 VDD2.t1 VSUBS 0.04936f
C50 VDD2.n2 VSUBS 0.047906f
C51 VDD2.n3 VSUBS 0.014316f
C52 VDD2.n4 VSUBS 0.009287f
C53 VDD2.n5 VSUBS 0.115458f
C54 VDD2.n6 VSUBS 0.258213f
C55 VDD2.n7 VSUBS 0.019064f
C56 VDD2.n8 VSUBS 0.049239f
C57 VDD2.t0 VSUBS 0.04936f
C58 VDD2.n9 VSUBS 0.047906f
C59 VDD2.n10 VSUBS 0.014316f
C60 VDD2.n11 VSUBS 0.009287f
C61 VDD2.n12 VSUBS 0.115458f
C62 VDD2.n13 VSUBS 0.038741f
C63 VDD2.n14 VSUBS 1.21914f
C64 VTAIL.n0 VSUBS 0.023077f
C65 VTAIL.n1 VSUBS 0.059604f
C66 VTAIL.t0 VSUBS 0.059751f
C67 VTAIL.n2 VSUBS 0.05799f
C68 VTAIL.n3 VSUBS 0.01733f
C69 VTAIL.n4 VSUBS 0.011242f
C70 VTAIL.n5 VSUBS 0.139764f
C71 VTAIL.n6 VSUBS 0.032427f
C72 VTAIL.n7 VSUBS 0.706359f
C73 VTAIL.n8 VSUBS 0.023077f
C74 VTAIL.n9 VSUBS 0.059604f
C75 VTAIL.t3 VSUBS 0.059751f
C76 VTAIL.n10 VSUBS 0.05799f
C77 VTAIL.n11 VSUBS 0.01733f
C78 VTAIL.n12 VSUBS 0.011242f
C79 VTAIL.n13 VSUBS 0.139764f
C80 VTAIL.n14 VSUBS 0.032427f
C81 VTAIL.n15 VSUBS 0.731057f
C82 VTAIL.n16 VSUBS 0.023077f
C83 VTAIL.n17 VSUBS 0.059604f
C84 VTAIL.t1 VSUBS 0.059751f
C85 VTAIL.n18 VSUBS 0.05799f
C86 VTAIL.n19 VSUBS 0.01733f
C87 VTAIL.n20 VSUBS 0.011242f
C88 VTAIL.n21 VSUBS 0.139764f
C89 VTAIL.n22 VSUBS 0.032427f
C90 VTAIL.n23 VSUBS 0.616574f
C91 VTAIL.n24 VSUBS 0.023077f
C92 VTAIL.n25 VSUBS 0.059604f
C93 VTAIL.t2 VSUBS 0.059751f
C94 VTAIL.n26 VSUBS 0.05799f
C95 VTAIL.n27 VSUBS 0.01733f
C96 VTAIL.n28 VSUBS 0.011242f
C97 VTAIL.n29 VSUBS 0.139764f
C98 VTAIL.n30 VSUBS 0.032427f
C99 VTAIL.n31 VSUBS 0.552359f
C100 VN.t0 VSUBS 0.722981f
C101 VN.t1 VSUBS 1.25849f
C102 B.n0 VSUBS 0.008273f
C103 B.n1 VSUBS 0.008273f
C104 B.n2 VSUBS 0.012235f
C105 B.n3 VSUBS 0.009376f
C106 B.n4 VSUBS 0.009376f
C107 B.n5 VSUBS 0.009376f
C108 B.n6 VSUBS 0.009376f
C109 B.n7 VSUBS 0.009376f
C110 B.n8 VSUBS 0.009376f
C111 B.n9 VSUBS 0.009376f
C112 B.n10 VSUBS 0.009376f
C113 B.n11 VSUBS 0.021044f
C114 B.n12 VSUBS 0.009376f
C115 B.n13 VSUBS 0.009376f
C116 B.n14 VSUBS 0.009376f
C117 B.n15 VSUBS 0.009376f
C118 B.n16 VSUBS 0.009376f
C119 B.n17 VSUBS 0.009376f
C120 B.t1 VSUBS 0.044198f
C121 B.t2 VSUBS 0.053555f
C122 B.t0 VSUBS 0.208488f
C123 B.n18 VSUBS 0.095231f
C124 B.n19 VSUBS 0.083267f
C125 B.n20 VSUBS 0.009376f
C126 B.n21 VSUBS 0.009376f
C127 B.n22 VSUBS 0.009376f
C128 B.n23 VSUBS 0.009376f
C129 B.n24 VSUBS 0.00524f
C130 B.n25 VSUBS 0.009376f
C131 B.t10 VSUBS 0.044198f
C132 B.t11 VSUBS 0.053555f
C133 B.t9 VSUBS 0.208488f
C134 B.n26 VSUBS 0.095231f
C135 B.n27 VSUBS 0.083267f
C136 B.n28 VSUBS 0.021723f
C137 B.n29 VSUBS 0.009376f
C138 B.n30 VSUBS 0.009376f
C139 B.n31 VSUBS 0.009376f
C140 B.n32 VSUBS 0.009376f
C141 B.n33 VSUBS 0.022803f
C142 B.n34 VSUBS 0.009376f
C143 B.n35 VSUBS 0.009376f
C144 B.n36 VSUBS 0.009376f
C145 B.n37 VSUBS 0.009376f
C146 B.n38 VSUBS 0.009376f
C147 B.n39 VSUBS 0.009376f
C148 B.n40 VSUBS 0.009376f
C149 B.n41 VSUBS 0.009376f
C150 B.n42 VSUBS 0.009376f
C151 B.n43 VSUBS 0.009376f
C152 B.n44 VSUBS 0.009376f
C153 B.n45 VSUBS 0.009376f
C154 B.n46 VSUBS 0.009376f
C155 B.n47 VSUBS 0.009376f
C156 B.n48 VSUBS 0.009376f
C157 B.n49 VSUBS 0.009376f
C158 B.n50 VSUBS 0.009376f
C159 B.n51 VSUBS 0.009376f
C160 B.n52 VSUBS 0.009376f
C161 B.n53 VSUBS 0.022153f
C162 B.n54 VSUBS 0.009376f
C163 B.n55 VSUBS 0.009376f
C164 B.n56 VSUBS 0.009376f
C165 B.n57 VSUBS 0.009376f
C166 B.n58 VSUBS 0.009376f
C167 B.n59 VSUBS 0.008825f
C168 B.n60 VSUBS 0.009376f
C169 B.n61 VSUBS 0.009376f
C170 B.n62 VSUBS 0.009376f
C171 B.n63 VSUBS 0.009376f
C172 B.n64 VSUBS 0.009376f
C173 B.t5 VSUBS 0.044198f
C174 B.t4 VSUBS 0.053555f
C175 B.t3 VSUBS 0.208488f
C176 B.n65 VSUBS 0.095231f
C177 B.n66 VSUBS 0.083267f
C178 B.n67 VSUBS 0.009376f
C179 B.n68 VSUBS 0.009376f
C180 B.n69 VSUBS 0.009376f
C181 B.n70 VSUBS 0.009376f
C182 B.n71 VSUBS 0.009376f
C183 B.n72 VSUBS 0.022803f
C184 B.n73 VSUBS 0.009376f
C185 B.n74 VSUBS 0.009376f
C186 B.n75 VSUBS 0.009376f
C187 B.n76 VSUBS 0.009376f
C188 B.n77 VSUBS 0.009376f
C189 B.n78 VSUBS 0.009376f
C190 B.n79 VSUBS 0.009376f
C191 B.n80 VSUBS 0.009376f
C192 B.n81 VSUBS 0.009376f
C193 B.n82 VSUBS 0.009376f
C194 B.n83 VSUBS 0.009376f
C195 B.n84 VSUBS 0.009376f
C196 B.n85 VSUBS 0.009376f
C197 B.n86 VSUBS 0.009376f
C198 B.n87 VSUBS 0.009376f
C199 B.n88 VSUBS 0.009376f
C200 B.n89 VSUBS 0.009376f
C201 B.n90 VSUBS 0.009376f
C202 B.n91 VSUBS 0.009376f
C203 B.n92 VSUBS 0.009376f
C204 B.n93 VSUBS 0.009376f
C205 B.n94 VSUBS 0.009376f
C206 B.n95 VSUBS 0.009376f
C207 B.n96 VSUBS 0.009376f
C208 B.n97 VSUBS 0.009376f
C209 B.n98 VSUBS 0.009376f
C210 B.n99 VSUBS 0.009376f
C211 B.n100 VSUBS 0.009376f
C212 B.n101 VSUBS 0.009376f
C213 B.n102 VSUBS 0.009376f
C214 B.n103 VSUBS 0.009376f
C215 B.n104 VSUBS 0.009376f
C216 B.n105 VSUBS 0.009376f
C217 B.n106 VSUBS 0.009376f
C218 B.n107 VSUBS 0.021044f
C219 B.n108 VSUBS 0.021044f
C220 B.n109 VSUBS 0.022803f
C221 B.n110 VSUBS 0.009376f
C222 B.n111 VSUBS 0.009376f
C223 B.n112 VSUBS 0.009376f
C224 B.n113 VSUBS 0.009376f
C225 B.n114 VSUBS 0.009376f
C226 B.n115 VSUBS 0.009376f
C227 B.n116 VSUBS 0.009376f
C228 B.n117 VSUBS 0.009376f
C229 B.n118 VSUBS 0.009376f
C230 B.n119 VSUBS 0.009376f
C231 B.n120 VSUBS 0.009376f
C232 B.n121 VSUBS 0.009376f
C233 B.n122 VSUBS 0.009376f
C234 B.n123 VSUBS 0.009376f
C235 B.n124 VSUBS 0.009376f
C236 B.n125 VSUBS 0.009376f
C237 B.n126 VSUBS 0.008825f
C238 B.n127 VSUBS 0.021723f
C239 B.n128 VSUBS 0.00524f
C240 B.n129 VSUBS 0.009376f
C241 B.n130 VSUBS 0.009376f
C242 B.n131 VSUBS 0.009376f
C243 B.n132 VSUBS 0.009376f
C244 B.n133 VSUBS 0.009376f
C245 B.n134 VSUBS 0.009376f
C246 B.n135 VSUBS 0.009376f
C247 B.n136 VSUBS 0.009376f
C248 B.n137 VSUBS 0.009376f
C249 B.n138 VSUBS 0.009376f
C250 B.n139 VSUBS 0.009376f
C251 B.n140 VSUBS 0.009376f
C252 B.t8 VSUBS 0.044198f
C253 B.t7 VSUBS 0.053555f
C254 B.t6 VSUBS 0.208488f
C255 B.n141 VSUBS 0.095231f
C256 B.n142 VSUBS 0.083267f
C257 B.n143 VSUBS 0.021723f
C258 B.n144 VSUBS 0.00524f
C259 B.n145 VSUBS 0.009376f
C260 B.n146 VSUBS 0.009376f
C261 B.n147 VSUBS 0.009376f
C262 B.n148 VSUBS 0.009376f
C263 B.n149 VSUBS 0.009376f
C264 B.n150 VSUBS 0.009376f
C265 B.n151 VSUBS 0.009376f
C266 B.n152 VSUBS 0.009376f
C267 B.n153 VSUBS 0.009376f
C268 B.n154 VSUBS 0.009376f
C269 B.n155 VSUBS 0.009376f
C270 B.n156 VSUBS 0.009376f
C271 B.n157 VSUBS 0.009376f
C272 B.n158 VSUBS 0.009376f
C273 B.n159 VSUBS 0.009376f
C274 B.n160 VSUBS 0.009376f
C275 B.n161 VSUBS 0.009376f
C276 B.n162 VSUBS 0.021694f
C277 B.n163 VSUBS 0.022803f
C278 B.n164 VSUBS 0.021044f
C279 B.n165 VSUBS 0.009376f
C280 B.n166 VSUBS 0.009376f
C281 B.n167 VSUBS 0.009376f
C282 B.n168 VSUBS 0.009376f
C283 B.n169 VSUBS 0.009376f
C284 B.n170 VSUBS 0.009376f
C285 B.n171 VSUBS 0.009376f
C286 B.n172 VSUBS 0.009376f
C287 B.n173 VSUBS 0.009376f
C288 B.n174 VSUBS 0.009376f
C289 B.n175 VSUBS 0.009376f
C290 B.n176 VSUBS 0.009376f
C291 B.n177 VSUBS 0.009376f
C292 B.n178 VSUBS 0.009376f
C293 B.n179 VSUBS 0.009376f
C294 B.n180 VSUBS 0.009376f
C295 B.n181 VSUBS 0.009376f
C296 B.n182 VSUBS 0.009376f
C297 B.n183 VSUBS 0.009376f
C298 B.n184 VSUBS 0.009376f
C299 B.n185 VSUBS 0.009376f
C300 B.n186 VSUBS 0.009376f
C301 B.n187 VSUBS 0.009376f
C302 B.n188 VSUBS 0.009376f
C303 B.n189 VSUBS 0.009376f
C304 B.n190 VSUBS 0.009376f
C305 B.n191 VSUBS 0.009376f
C306 B.n192 VSUBS 0.009376f
C307 B.n193 VSUBS 0.009376f
C308 B.n194 VSUBS 0.009376f
C309 B.n195 VSUBS 0.009376f
C310 B.n196 VSUBS 0.009376f
C311 B.n197 VSUBS 0.009376f
C312 B.n198 VSUBS 0.009376f
C313 B.n199 VSUBS 0.009376f
C314 B.n200 VSUBS 0.009376f
C315 B.n201 VSUBS 0.009376f
C316 B.n202 VSUBS 0.009376f
C317 B.n203 VSUBS 0.009376f
C318 B.n204 VSUBS 0.009376f
C319 B.n205 VSUBS 0.009376f
C320 B.n206 VSUBS 0.009376f
C321 B.n207 VSUBS 0.009376f
C322 B.n208 VSUBS 0.009376f
C323 B.n209 VSUBS 0.009376f
C324 B.n210 VSUBS 0.009376f
C325 B.n211 VSUBS 0.009376f
C326 B.n212 VSUBS 0.009376f
C327 B.n213 VSUBS 0.009376f
C328 B.n214 VSUBS 0.009376f
C329 B.n215 VSUBS 0.009376f
C330 B.n216 VSUBS 0.009376f
C331 B.n217 VSUBS 0.009376f
C332 B.n218 VSUBS 0.009376f
C333 B.n219 VSUBS 0.009376f
C334 B.n220 VSUBS 0.009376f
C335 B.n221 VSUBS 0.009376f
C336 B.n222 VSUBS 0.021044f
C337 B.n223 VSUBS 0.021044f
C338 B.n224 VSUBS 0.022803f
C339 B.n225 VSUBS 0.009376f
C340 B.n226 VSUBS 0.009376f
C341 B.n227 VSUBS 0.009376f
C342 B.n228 VSUBS 0.009376f
C343 B.n229 VSUBS 0.009376f
C344 B.n230 VSUBS 0.009376f
C345 B.n231 VSUBS 0.009376f
C346 B.n232 VSUBS 0.009376f
C347 B.n233 VSUBS 0.009376f
C348 B.n234 VSUBS 0.009376f
C349 B.n235 VSUBS 0.009376f
C350 B.n236 VSUBS 0.009376f
C351 B.n237 VSUBS 0.009376f
C352 B.n238 VSUBS 0.009376f
C353 B.n239 VSUBS 0.009376f
C354 B.n240 VSUBS 0.008825f
C355 B.n241 VSUBS 0.009376f
C356 B.n242 VSUBS 0.009376f
C357 B.n243 VSUBS 0.009376f
C358 B.n244 VSUBS 0.009376f
C359 B.n245 VSUBS 0.009376f
C360 B.n246 VSUBS 0.009376f
C361 B.n247 VSUBS 0.009376f
C362 B.n248 VSUBS 0.009376f
C363 B.n249 VSUBS 0.009376f
C364 B.n250 VSUBS 0.009376f
C365 B.n251 VSUBS 0.009376f
C366 B.n252 VSUBS 0.009376f
C367 B.n253 VSUBS 0.009376f
C368 B.n254 VSUBS 0.009376f
C369 B.n255 VSUBS 0.009376f
C370 B.n256 VSUBS 0.00524f
C371 B.n257 VSUBS 0.021723f
C372 B.n258 VSUBS 0.008825f
C373 B.n259 VSUBS 0.009376f
C374 B.n260 VSUBS 0.009376f
C375 B.n261 VSUBS 0.009376f
C376 B.n262 VSUBS 0.009376f
C377 B.n263 VSUBS 0.009376f
C378 B.n264 VSUBS 0.009376f
C379 B.n265 VSUBS 0.009376f
C380 B.n266 VSUBS 0.009376f
C381 B.n267 VSUBS 0.009376f
C382 B.n268 VSUBS 0.009376f
C383 B.n269 VSUBS 0.009376f
C384 B.n270 VSUBS 0.009376f
C385 B.n271 VSUBS 0.009376f
C386 B.n272 VSUBS 0.009376f
C387 B.n273 VSUBS 0.009376f
C388 B.n274 VSUBS 0.022803f
C389 B.n275 VSUBS 0.022803f
C390 B.n276 VSUBS 0.021044f
C391 B.n277 VSUBS 0.009376f
C392 B.n278 VSUBS 0.009376f
C393 B.n279 VSUBS 0.009376f
C394 B.n280 VSUBS 0.009376f
C395 B.n281 VSUBS 0.009376f
C396 B.n282 VSUBS 0.009376f
C397 B.n283 VSUBS 0.009376f
C398 B.n284 VSUBS 0.009376f
C399 B.n285 VSUBS 0.009376f
C400 B.n286 VSUBS 0.009376f
C401 B.n287 VSUBS 0.009376f
C402 B.n288 VSUBS 0.009376f
C403 B.n289 VSUBS 0.009376f
C404 B.n290 VSUBS 0.009376f
C405 B.n291 VSUBS 0.009376f
C406 B.n292 VSUBS 0.009376f
C407 B.n293 VSUBS 0.009376f
C408 B.n294 VSUBS 0.009376f
C409 B.n295 VSUBS 0.009376f
C410 B.n296 VSUBS 0.009376f
C411 B.n297 VSUBS 0.009376f
C412 B.n298 VSUBS 0.009376f
C413 B.n299 VSUBS 0.009376f
C414 B.n300 VSUBS 0.009376f
C415 B.n301 VSUBS 0.009376f
C416 B.n302 VSUBS 0.009376f
C417 B.n303 VSUBS 0.012235f
C418 B.n304 VSUBS 0.013034f
C419 B.n305 VSUBS 0.025919f
.ends

