* NGSPICE file created from diff_pair_sample_0293.ext - technology: sky130A

.subckt diff_pair_sample_0293 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t9 w_n2460_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.3498 ps=2.45 w=2.12 l=1.16
X1 B.t11 B.t9 B.t10 w_n2460_n1392# sky130_fd_pr__pfet_01v8 ad=0.8268 pd=5.02 as=0 ps=0 w=2.12 l=1.16
X2 VTAIL.t4 VN.t0 VDD2.t7 w_n2460_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.3498 ps=2.45 w=2.12 l=1.16
X3 B.t8 B.t6 B.t7 w_n2460_n1392# sky130_fd_pr__pfet_01v8 ad=0.8268 pd=5.02 as=0 ps=0 w=2.12 l=1.16
X4 VTAIL.t6 VN.t1 VDD2.t6 w_n2460_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.3498 ps=2.45 w=2.12 l=1.16
X5 VTAIL.t14 VP.t1 VDD1.t6 w_n2460_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.3498 ps=2.45 w=2.12 l=1.16
X6 VTAIL.t15 VP.t2 VDD1.t5 w_n2460_n1392# sky130_fd_pr__pfet_01v8 ad=0.8268 pd=5.02 as=0.3498 ps=2.45 w=2.12 l=1.16
X7 VDD2.t5 VN.t2 VTAIL.t1 w_n2460_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.8268 ps=5.02 w=2.12 l=1.16
X8 VDD1.t4 VP.t3 VTAIL.t12 w_n2460_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.8268 ps=5.02 w=2.12 l=1.16
X9 VDD1.t3 VP.t4 VTAIL.t10 w_n2460_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.8268 ps=5.02 w=2.12 l=1.16
X10 VDD2.t4 VN.t3 VTAIL.t3 w_n2460_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.3498 ps=2.45 w=2.12 l=1.16
X11 VTAIL.t8 VP.t5 VDD1.t2 w_n2460_n1392# sky130_fd_pr__pfet_01v8 ad=0.8268 pd=5.02 as=0.3498 ps=2.45 w=2.12 l=1.16
X12 B.t5 B.t3 B.t4 w_n2460_n1392# sky130_fd_pr__pfet_01v8 ad=0.8268 pd=5.02 as=0 ps=0 w=2.12 l=1.16
X13 VTAIL.t5 VN.t4 VDD2.t3 w_n2460_n1392# sky130_fd_pr__pfet_01v8 ad=0.8268 pd=5.02 as=0.3498 ps=2.45 w=2.12 l=1.16
X14 VTAIL.t0 VN.t5 VDD2.t2 w_n2460_n1392# sky130_fd_pr__pfet_01v8 ad=0.8268 pd=5.02 as=0.3498 ps=2.45 w=2.12 l=1.16
X15 B.t2 B.t0 B.t1 w_n2460_n1392# sky130_fd_pr__pfet_01v8 ad=0.8268 pd=5.02 as=0 ps=0 w=2.12 l=1.16
X16 VDD1.t1 VP.t6 VTAIL.t11 w_n2460_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.3498 ps=2.45 w=2.12 l=1.16
X17 VTAIL.t13 VP.t7 VDD1.t0 w_n2460_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.3498 ps=2.45 w=2.12 l=1.16
X18 VDD2.t1 VN.t6 VTAIL.t2 w_n2460_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.3498 ps=2.45 w=2.12 l=1.16
X19 VDD2.t0 VN.t7 VTAIL.t7 w_n2460_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.8268 ps=5.02 w=2.12 l=1.16
R0 VP.n23 VP.n5 174.334
R1 VP.n40 VP.n39 174.334
R2 VP.n22 VP.n21 174.334
R3 VP.n12 VP.n11 161.3
R4 VP.n13 VP.n8 161.3
R5 VP.n16 VP.n15 161.3
R6 VP.n17 VP.n7 161.3
R7 VP.n19 VP.n18 161.3
R8 VP.n20 VP.n6 161.3
R9 VP.n38 VP.n0 161.3
R10 VP.n37 VP.n36 161.3
R11 VP.n35 VP.n1 161.3
R12 VP.n34 VP.n33 161.3
R13 VP.n31 VP.n2 161.3
R14 VP.n30 VP.n29 161.3
R15 VP.n28 VP.n27 161.3
R16 VP.n26 VP.n4 161.3
R17 VP.n25 VP.n24 161.3
R18 VP.n10 VP.t2 73.7195
R19 VP.n10 VP.n9 51.8775
R20 VP.n5 VP.t5 44.0453
R21 VP.n3 VP.t6 44.0453
R22 VP.n32 VP.t1 44.0453
R23 VP.n39 VP.t4 44.0453
R24 VP.n21 VP.t3 44.0453
R25 VP.n14 VP.t7 44.0453
R26 VP.n9 VP.t0 44.0453
R27 VP.n27 VP.n26 41.5458
R28 VP.n37 VP.n1 41.5458
R29 VP.n19 VP.n7 41.5458
R30 VP.n31 VP.n30 40.577
R31 VP.n33 VP.n31 40.577
R32 VP.n15 VP.n13 40.577
R33 VP.n13 VP.n12 40.577
R34 VP.n26 VP.n25 39.6083
R35 VP.n38 VP.n37 39.6083
R36 VP.n20 VP.n19 39.6083
R37 VP.n23 VP.n22 36.5384
R38 VP.n11 VP.n10 27.1451
R39 VP.n27 VP.n3 12.5423
R40 VP.n32 VP.n1 12.5423
R41 VP.n14 VP.n7 12.5423
R42 VP.n30 VP.n3 12.0505
R43 VP.n33 VP.n32 12.0505
R44 VP.n15 VP.n14 12.0505
R45 VP.n12 VP.n9 12.0505
R46 VP.n25 VP.n5 11.5587
R47 VP.n39 VP.n38 11.5587
R48 VP.n21 VP.n20 11.5587
R49 VP.n11 VP.n8 0.189894
R50 VP.n16 VP.n8 0.189894
R51 VP.n17 VP.n16 0.189894
R52 VP.n18 VP.n17 0.189894
R53 VP.n18 VP.n6 0.189894
R54 VP.n22 VP.n6 0.189894
R55 VP.n24 VP.n23 0.189894
R56 VP.n24 VP.n4 0.189894
R57 VP.n28 VP.n4 0.189894
R58 VP.n29 VP.n28 0.189894
R59 VP.n29 VP.n2 0.189894
R60 VP.n34 VP.n2 0.189894
R61 VP.n35 VP.n34 0.189894
R62 VP.n36 VP.n35 0.189894
R63 VP.n36 VP.n0 0.189894
R64 VP.n40 VP.n0 0.189894
R65 VP VP.n40 0.0516364
R66 VTAIL.n15 VTAIL.t7 171.044
R67 VTAIL.n2 VTAIL.t0 171.044
R68 VTAIL.n3 VTAIL.t10 171.044
R69 VTAIL.n6 VTAIL.t8 171.044
R70 VTAIL.n14 VTAIL.t12 171.044
R71 VTAIL.n11 VTAIL.t15 171.044
R72 VTAIL.n10 VTAIL.t1 171.044
R73 VTAIL.n7 VTAIL.t5 171.044
R74 VTAIL.n13 VTAIL.n12 155.713
R75 VTAIL.n9 VTAIL.n8 155.713
R76 VTAIL.n1 VTAIL.n0 155.712
R77 VTAIL.n5 VTAIL.n4 155.712
R78 VTAIL.n15 VTAIL.n14 15.4789
R79 VTAIL.n7 VTAIL.n6 15.4789
R80 VTAIL.n0 VTAIL.t3 15.333
R81 VTAIL.n0 VTAIL.t4 15.333
R82 VTAIL.n4 VTAIL.t11 15.333
R83 VTAIL.n4 VTAIL.t14 15.333
R84 VTAIL.n12 VTAIL.t9 15.333
R85 VTAIL.n12 VTAIL.t13 15.333
R86 VTAIL.n8 VTAIL.t2 15.333
R87 VTAIL.n8 VTAIL.t6 15.333
R88 VTAIL.n9 VTAIL.n7 1.28498
R89 VTAIL.n10 VTAIL.n9 1.28498
R90 VTAIL.n13 VTAIL.n11 1.28498
R91 VTAIL.n14 VTAIL.n13 1.28498
R92 VTAIL.n6 VTAIL.n5 1.28498
R93 VTAIL.n5 VTAIL.n3 1.28498
R94 VTAIL.n2 VTAIL.n1 1.28498
R95 VTAIL VTAIL.n15 1.22679
R96 VTAIL.n11 VTAIL.n10 0.470328
R97 VTAIL.n3 VTAIL.n2 0.470328
R98 VTAIL VTAIL.n1 0.0586897
R99 VDD1 VDD1.n0 173.091
R100 VDD1.n3 VDD1.n2 172.977
R101 VDD1.n3 VDD1.n1 172.977
R102 VDD1.n5 VDD1.n4 172.391
R103 VDD1.n5 VDD1.n3 31.9061
R104 VDD1.n4 VDD1.t0 15.333
R105 VDD1.n4 VDD1.t4 15.333
R106 VDD1.n0 VDD1.t5 15.333
R107 VDD1.n0 VDD1.t7 15.333
R108 VDD1.n2 VDD1.t6 15.333
R109 VDD1.n2 VDD1.t3 15.333
R110 VDD1.n1 VDD1.t2 15.333
R111 VDD1.n1 VDD1.t1 15.333
R112 VDD1 VDD1.n5 0.584552
R113 B.n296 B.n295 585
R114 B.n297 B.n38 585
R115 B.n299 B.n298 585
R116 B.n300 B.n37 585
R117 B.n302 B.n301 585
R118 B.n303 B.n36 585
R119 B.n305 B.n304 585
R120 B.n306 B.n35 585
R121 B.n308 B.n307 585
R122 B.n309 B.n34 585
R123 B.n311 B.n310 585
R124 B.n312 B.n33 585
R125 B.n314 B.n313 585
R126 B.n316 B.n315 585
R127 B.n317 B.n29 585
R128 B.n319 B.n318 585
R129 B.n320 B.n28 585
R130 B.n322 B.n321 585
R131 B.n323 B.n27 585
R132 B.n325 B.n324 585
R133 B.n326 B.n26 585
R134 B.n328 B.n327 585
R135 B.n330 B.n23 585
R136 B.n332 B.n331 585
R137 B.n333 B.n22 585
R138 B.n335 B.n334 585
R139 B.n336 B.n21 585
R140 B.n338 B.n337 585
R141 B.n339 B.n20 585
R142 B.n341 B.n340 585
R143 B.n342 B.n19 585
R144 B.n344 B.n343 585
R145 B.n345 B.n18 585
R146 B.n347 B.n346 585
R147 B.n348 B.n17 585
R148 B.n294 B.n39 585
R149 B.n293 B.n292 585
R150 B.n291 B.n40 585
R151 B.n290 B.n289 585
R152 B.n288 B.n41 585
R153 B.n287 B.n286 585
R154 B.n285 B.n42 585
R155 B.n284 B.n283 585
R156 B.n282 B.n43 585
R157 B.n281 B.n280 585
R158 B.n279 B.n44 585
R159 B.n278 B.n277 585
R160 B.n276 B.n45 585
R161 B.n275 B.n274 585
R162 B.n273 B.n46 585
R163 B.n272 B.n271 585
R164 B.n270 B.n47 585
R165 B.n269 B.n268 585
R166 B.n267 B.n48 585
R167 B.n266 B.n265 585
R168 B.n264 B.n49 585
R169 B.n263 B.n262 585
R170 B.n261 B.n50 585
R171 B.n260 B.n259 585
R172 B.n258 B.n51 585
R173 B.n257 B.n256 585
R174 B.n255 B.n52 585
R175 B.n254 B.n253 585
R176 B.n252 B.n53 585
R177 B.n251 B.n250 585
R178 B.n249 B.n54 585
R179 B.n248 B.n247 585
R180 B.n246 B.n55 585
R181 B.n245 B.n244 585
R182 B.n243 B.n56 585
R183 B.n242 B.n241 585
R184 B.n240 B.n57 585
R185 B.n239 B.n238 585
R186 B.n237 B.n58 585
R187 B.n236 B.n235 585
R188 B.n234 B.n59 585
R189 B.n233 B.n232 585
R190 B.n231 B.n60 585
R191 B.n230 B.n229 585
R192 B.n228 B.n61 585
R193 B.n227 B.n226 585
R194 B.n225 B.n62 585
R195 B.n224 B.n223 585
R196 B.n222 B.n63 585
R197 B.n221 B.n220 585
R198 B.n219 B.n64 585
R199 B.n218 B.n217 585
R200 B.n216 B.n65 585
R201 B.n215 B.n214 585
R202 B.n213 B.n66 585
R203 B.n212 B.n211 585
R204 B.n210 B.n67 585
R205 B.n209 B.n208 585
R206 B.n207 B.n68 585
R207 B.n206 B.n205 585
R208 B.n204 B.n69 585
R209 B.n150 B.n91 585
R210 B.n152 B.n151 585
R211 B.n153 B.n90 585
R212 B.n155 B.n154 585
R213 B.n156 B.n89 585
R214 B.n158 B.n157 585
R215 B.n159 B.n88 585
R216 B.n161 B.n160 585
R217 B.n162 B.n87 585
R218 B.n164 B.n163 585
R219 B.n165 B.n86 585
R220 B.n167 B.n166 585
R221 B.n168 B.n83 585
R222 B.n171 B.n170 585
R223 B.n172 B.n82 585
R224 B.n174 B.n173 585
R225 B.n175 B.n81 585
R226 B.n177 B.n176 585
R227 B.n178 B.n80 585
R228 B.n180 B.n179 585
R229 B.n181 B.n79 585
R230 B.n183 B.n182 585
R231 B.n185 B.n184 585
R232 B.n186 B.n75 585
R233 B.n188 B.n187 585
R234 B.n189 B.n74 585
R235 B.n191 B.n190 585
R236 B.n192 B.n73 585
R237 B.n194 B.n193 585
R238 B.n195 B.n72 585
R239 B.n197 B.n196 585
R240 B.n198 B.n71 585
R241 B.n200 B.n199 585
R242 B.n201 B.n70 585
R243 B.n203 B.n202 585
R244 B.n149 B.n148 585
R245 B.n147 B.n92 585
R246 B.n146 B.n145 585
R247 B.n144 B.n93 585
R248 B.n143 B.n142 585
R249 B.n141 B.n94 585
R250 B.n140 B.n139 585
R251 B.n138 B.n95 585
R252 B.n137 B.n136 585
R253 B.n135 B.n96 585
R254 B.n134 B.n133 585
R255 B.n132 B.n97 585
R256 B.n131 B.n130 585
R257 B.n129 B.n98 585
R258 B.n128 B.n127 585
R259 B.n126 B.n99 585
R260 B.n125 B.n124 585
R261 B.n123 B.n100 585
R262 B.n122 B.n121 585
R263 B.n120 B.n101 585
R264 B.n119 B.n118 585
R265 B.n117 B.n102 585
R266 B.n116 B.n115 585
R267 B.n114 B.n103 585
R268 B.n113 B.n112 585
R269 B.n111 B.n104 585
R270 B.n110 B.n109 585
R271 B.n108 B.n105 585
R272 B.n107 B.n106 585
R273 B.n2 B.n0 585
R274 B.n393 B.n1 585
R275 B.n392 B.n391 585
R276 B.n390 B.n3 585
R277 B.n389 B.n388 585
R278 B.n387 B.n4 585
R279 B.n386 B.n385 585
R280 B.n384 B.n5 585
R281 B.n383 B.n382 585
R282 B.n381 B.n6 585
R283 B.n380 B.n379 585
R284 B.n378 B.n7 585
R285 B.n377 B.n376 585
R286 B.n375 B.n8 585
R287 B.n374 B.n373 585
R288 B.n372 B.n9 585
R289 B.n371 B.n370 585
R290 B.n369 B.n10 585
R291 B.n368 B.n367 585
R292 B.n366 B.n11 585
R293 B.n365 B.n364 585
R294 B.n363 B.n12 585
R295 B.n362 B.n361 585
R296 B.n360 B.n13 585
R297 B.n359 B.n358 585
R298 B.n357 B.n14 585
R299 B.n356 B.n355 585
R300 B.n354 B.n15 585
R301 B.n353 B.n352 585
R302 B.n351 B.n16 585
R303 B.n350 B.n349 585
R304 B.n395 B.n394 585
R305 B.n148 B.n91 478.086
R306 B.n350 B.n17 478.086
R307 B.n202 B.n69 478.086
R308 B.n296 B.n39 478.086
R309 B.n76 B.t0 247.947
R310 B.n84 B.t9 247.947
R311 B.n24 B.t3 247.947
R312 B.n30 B.t6 247.947
R313 B.n76 B.t2 200.751
R314 B.n30 B.t7 200.751
R315 B.n84 B.t11 200.75
R316 B.n24 B.t4 200.75
R317 B.n77 B.t1 171.855
R318 B.n31 B.t8 171.855
R319 B.n85 B.t10 171.853
R320 B.n25 B.t5 171.853
R321 B.n148 B.n147 163.367
R322 B.n147 B.n146 163.367
R323 B.n146 B.n93 163.367
R324 B.n142 B.n93 163.367
R325 B.n142 B.n141 163.367
R326 B.n141 B.n140 163.367
R327 B.n140 B.n95 163.367
R328 B.n136 B.n95 163.367
R329 B.n136 B.n135 163.367
R330 B.n135 B.n134 163.367
R331 B.n134 B.n97 163.367
R332 B.n130 B.n97 163.367
R333 B.n130 B.n129 163.367
R334 B.n129 B.n128 163.367
R335 B.n128 B.n99 163.367
R336 B.n124 B.n99 163.367
R337 B.n124 B.n123 163.367
R338 B.n123 B.n122 163.367
R339 B.n122 B.n101 163.367
R340 B.n118 B.n101 163.367
R341 B.n118 B.n117 163.367
R342 B.n117 B.n116 163.367
R343 B.n116 B.n103 163.367
R344 B.n112 B.n103 163.367
R345 B.n112 B.n111 163.367
R346 B.n111 B.n110 163.367
R347 B.n110 B.n105 163.367
R348 B.n106 B.n105 163.367
R349 B.n106 B.n2 163.367
R350 B.n394 B.n2 163.367
R351 B.n394 B.n393 163.367
R352 B.n393 B.n392 163.367
R353 B.n392 B.n3 163.367
R354 B.n388 B.n3 163.367
R355 B.n388 B.n387 163.367
R356 B.n387 B.n386 163.367
R357 B.n386 B.n5 163.367
R358 B.n382 B.n5 163.367
R359 B.n382 B.n381 163.367
R360 B.n381 B.n380 163.367
R361 B.n380 B.n7 163.367
R362 B.n376 B.n7 163.367
R363 B.n376 B.n375 163.367
R364 B.n375 B.n374 163.367
R365 B.n374 B.n9 163.367
R366 B.n370 B.n9 163.367
R367 B.n370 B.n369 163.367
R368 B.n369 B.n368 163.367
R369 B.n368 B.n11 163.367
R370 B.n364 B.n11 163.367
R371 B.n364 B.n363 163.367
R372 B.n363 B.n362 163.367
R373 B.n362 B.n13 163.367
R374 B.n358 B.n13 163.367
R375 B.n358 B.n357 163.367
R376 B.n357 B.n356 163.367
R377 B.n356 B.n15 163.367
R378 B.n352 B.n15 163.367
R379 B.n352 B.n351 163.367
R380 B.n351 B.n350 163.367
R381 B.n152 B.n91 163.367
R382 B.n153 B.n152 163.367
R383 B.n154 B.n153 163.367
R384 B.n154 B.n89 163.367
R385 B.n158 B.n89 163.367
R386 B.n159 B.n158 163.367
R387 B.n160 B.n159 163.367
R388 B.n160 B.n87 163.367
R389 B.n164 B.n87 163.367
R390 B.n165 B.n164 163.367
R391 B.n166 B.n165 163.367
R392 B.n166 B.n83 163.367
R393 B.n171 B.n83 163.367
R394 B.n172 B.n171 163.367
R395 B.n173 B.n172 163.367
R396 B.n173 B.n81 163.367
R397 B.n177 B.n81 163.367
R398 B.n178 B.n177 163.367
R399 B.n179 B.n178 163.367
R400 B.n179 B.n79 163.367
R401 B.n183 B.n79 163.367
R402 B.n184 B.n183 163.367
R403 B.n184 B.n75 163.367
R404 B.n188 B.n75 163.367
R405 B.n189 B.n188 163.367
R406 B.n190 B.n189 163.367
R407 B.n190 B.n73 163.367
R408 B.n194 B.n73 163.367
R409 B.n195 B.n194 163.367
R410 B.n196 B.n195 163.367
R411 B.n196 B.n71 163.367
R412 B.n200 B.n71 163.367
R413 B.n201 B.n200 163.367
R414 B.n202 B.n201 163.367
R415 B.n206 B.n69 163.367
R416 B.n207 B.n206 163.367
R417 B.n208 B.n207 163.367
R418 B.n208 B.n67 163.367
R419 B.n212 B.n67 163.367
R420 B.n213 B.n212 163.367
R421 B.n214 B.n213 163.367
R422 B.n214 B.n65 163.367
R423 B.n218 B.n65 163.367
R424 B.n219 B.n218 163.367
R425 B.n220 B.n219 163.367
R426 B.n220 B.n63 163.367
R427 B.n224 B.n63 163.367
R428 B.n225 B.n224 163.367
R429 B.n226 B.n225 163.367
R430 B.n226 B.n61 163.367
R431 B.n230 B.n61 163.367
R432 B.n231 B.n230 163.367
R433 B.n232 B.n231 163.367
R434 B.n232 B.n59 163.367
R435 B.n236 B.n59 163.367
R436 B.n237 B.n236 163.367
R437 B.n238 B.n237 163.367
R438 B.n238 B.n57 163.367
R439 B.n242 B.n57 163.367
R440 B.n243 B.n242 163.367
R441 B.n244 B.n243 163.367
R442 B.n244 B.n55 163.367
R443 B.n248 B.n55 163.367
R444 B.n249 B.n248 163.367
R445 B.n250 B.n249 163.367
R446 B.n250 B.n53 163.367
R447 B.n254 B.n53 163.367
R448 B.n255 B.n254 163.367
R449 B.n256 B.n255 163.367
R450 B.n256 B.n51 163.367
R451 B.n260 B.n51 163.367
R452 B.n261 B.n260 163.367
R453 B.n262 B.n261 163.367
R454 B.n262 B.n49 163.367
R455 B.n266 B.n49 163.367
R456 B.n267 B.n266 163.367
R457 B.n268 B.n267 163.367
R458 B.n268 B.n47 163.367
R459 B.n272 B.n47 163.367
R460 B.n273 B.n272 163.367
R461 B.n274 B.n273 163.367
R462 B.n274 B.n45 163.367
R463 B.n278 B.n45 163.367
R464 B.n279 B.n278 163.367
R465 B.n280 B.n279 163.367
R466 B.n280 B.n43 163.367
R467 B.n284 B.n43 163.367
R468 B.n285 B.n284 163.367
R469 B.n286 B.n285 163.367
R470 B.n286 B.n41 163.367
R471 B.n290 B.n41 163.367
R472 B.n291 B.n290 163.367
R473 B.n292 B.n291 163.367
R474 B.n292 B.n39 163.367
R475 B.n346 B.n17 163.367
R476 B.n346 B.n345 163.367
R477 B.n345 B.n344 163.367
R478 B.n344 B.n19 163.367
R479 B.n340 B.n19 163.367
R480 B.n340 B.n339 163.367
R481 B.n339 B.n338 163.367
R482 B.n338 B.n21 163.367
R483 B.n334 B.n21 163.367
R484 B.n334 B.n333 163.367
R485 B.n333 B.n332 163.367
R486 B.n332 B.n23 163.367
R487 B.n327 B.n23 163.367
R488 B.n327 B.n326 163.367
R489 B.n326 B.n325 163.367
R490 B.n325 B.n27 163.367
R491 B.n321 B.n27 163.367
R492 B.n321 B.n320 163.367
R493 B.n320 B.n319 163.367
R494 B.n319 B.n29 163.367
R495 B.n315 B.n29 163.367
R496 B.n315 B.n314 163.367
R497 B.n314 B.n33 163.367
R498 B.n310 B.n33 163.367
R499 B.n310 B.n309 163.367
R500 B.n309 B.n308 163.367
R501 B.n308 B.n35 163.367
R502 B.n304 B.n35 163.367
R503 B.n304 B.n303 163.367
R504 B.n303 B.n302 163.367
R505 B.n302 B.n37 163.367
R506 B.n298 B.n37 163.367
R507 B.n298 B.n297 163.367
R508 B.n297 B.n296 163.367
R509 B.n78 B.n77 59.5399
R510 B.n169 B.n85 59.5399
R511 B.n329 B.n25 59.5399
R512 B.n32 B.n31 59.5399
R513 B.n349 B.n348 31.0639
R514 B.n295 B.n294 31.0639
R515 B.n204 B.n203 31.0639
R516 B.n150 B.n149 31.0639
R517 B.n77 B.n76 28.8975
R518 B.n85 B.n84 28.8975
R519 B.n25 B.n24 28.8975
R520 B.n31 B.n30 28.8975
R521 B B.n395 18.0485
R522 B.n348 B.n347 10.6151
R523 B.n347 B.n18 10.6151
R524 B.n343 B.n18 10.6151
R525 B.n343 B.n342 10.6151
R526 B.n342 B.n341 10.6151
R527 B.n341 B.n20 10.6151
R528 B.n337 B.n20 10.6151
R529 B.n337 B.n336 10.6151
R530 B.n336 B.n335 10.6151
R531 B.n335 B.n22 10.6151
R532 B.n331 B.n22 10.6151
R533 B.n331 B.n330 10.6151
R534 B.n328 B.n26 10.6151
R535 B.n324 B.n26 10.6151
R536 B.n324 B.n323 10.6151
R537 B.n323 B.n322 10.6151
R538 B.n322 B.n28 10.6151
R539 B.n318 B.n28 10.6151
R540 B.n318 B.n317 10.6151
R541 B.n317 B.n316 10.6151
R542 B.n313 B.n312 10.6151
R543 B.n312 B.n311 10.6151
R544 B.n311 B.n34 10.6151
R545 B.n307 B.n34 10.6151
R546 B.n307 B.n306 10.6151
R547 B.n306 B.n305 10.6151
R548 B.n305 B.n36 10.6151
R549 B.n301 B.n36 10.6151
R550 B.n301 B.n300 10.6151
R551 B.n300 B.n299 10.6151
R552 B.n299 B.n38 10.6151
R553 B.n295 B.n38 10.6151
R554 B.n205 B.n204 10.6151
R555 B.n205 B.n68 10.6151
R556 B.n209 B.n68 10.6151
R557 B.n210 B.n209 10.6151
R558 B.n211 B.n210 10.6151
R559 B.n211 B.n66 10.6151
R560 B.n215 B.n66 10.6151
R561 B.n216 B.n215 10.6151
R562 B.n217 B.n216 10.6151
R563 B.n217 B.n64 10.6151
R564 B.n221 B.n64 10.6151
R565 B.n222 B.n221 10.6151
R566 B.n223 B.n222 10.6151
R567 B.n223 B.n62 10.6151
R568 B.n227 B.n62 10.6151
R569 B.n228 B.n227 10.6151
R570 B.n229 B.n228 10.6151
R571 B.n229 B.n60 10.6151
R572 B.n233 B.n60 10.6151
R573 B.n234 B.n233 10.6151
R574 B.n235 B.n234 10.6151
R575 B.n235 B.n58 10.6151
R576 B.n239 B.n58 10.6151
R577 B.n240 B.n239 10.6151
R578 B.n241 B.n240 10.6151
R579 B.n241 B.n56 10.6151
R580 B.n245 B.n56 10.6151
R581 B.n246 B.n245 10.6151
R582 B.n247 B.n246 10.6151
R583 B.n247 B.n54 10.6151
R584 B.n251 B.n54 10.6151
R585 B.n252 B.n251 10.6151
R586 B.n253 B.n252 10.6151
R587 B.n253 B.n52 10.6151
R588 B.n257 B.n52 10.6151
R589 B.n258 B.n257 10.6151
R590 B.n259 B.n258 10.6151
R591 B.n259 B.n50 10.6151
R592 B.n263 B.n50 10.6151
R593 B.n264 B.n263 10.6151
R594 B.n265 B.n264 10.6151
R595 B.n265 B.n48 10.6151
R596 B.n269 B.n48 10.6151
R597 B.n270 B.n269 10.6151
R598 B.n271 B.n270 10.6151
R599 B.n271 B.n46 10.6151
R600 B.n275 B.n46 10.6151
R601 B.n276 B.n275 10.6151
R602 B.n277 B.n276 10.6151
R603 B.n277 B.n44 10.6151
R604 B.n281 B.n44 10.6151
R605 B.n282 B.n281 10.6151
R606 B.n283 B.n282 10.6151
R607 B.n283 B.n42 10.6151
R608 B.n287 B.n42 10.6151
R609 B.n288 B.n287 10.6151
R610 B.n289 B.n288 10.6151
R611 B.n289 B.n40 10.6151
R612 B.n293 B.n40 10.6151
R613 B.n294 B.n293 10.6151
R614 B.n151 B.n150 10.6151
R615 B.n151 B.n90 10.6151
R616 B.n155 B.n90 10.6151
R617 B.n156 B.n155 10.6151
R618 B.n157 B.n156 10.6151
R619 B.n157 B.n88 10.6151
R620 B.n161 B.n88 10.6151
R621 B.n162 B.n161 10.6151
R622 B.n163 B.n162 10.6151
R623 B.n163 B.n86 10.6151
R624 B.n167 B.n86 10.6151
R625 B.n168 B.n167 10.6151
R626 B.n170 B.n82 10.6151
R627 B.n174 B.n82 10.6151
R628 B.n175 B.n174 10.6151
R629 B.n176 B.n175 10.6151
R630 B.n176 B.n80 10.6151
R631 B.n180 B.n80 10.6151
R632 B.n181 B.n180 10.6151
R633 B.n182 B.n181 10.6151
R634 B.n186 B.n185 10.6151
R635 B.n187 B.n186 10.6151
R636 B.n187 B.n74 10.6151
R637 B.n191 B.n74 10.6151
R638 B.n192 B.n191 10.6151
R639 B.n193 B.n192 10.6151
R640 B.n193 B.n72 10.6151
R641 B.n197 B.n72 10.6151
R642 B.n198 B.n197 10.6151
R643 B.n199 B.n198 10.6151
R644 B.n199 B.n70 10.6151
R645 B.n203 B.n70 10.6151
R646 B.n149 B.n92 10.6151
R647 B.n145 B.n92 10.6151
R648 B.n145 B.n144 10.6151
R649 B.n144 B.n143 10.6151
R650 B.n143 B.n94 10.6151
R651 B.n139 B.n94 10.6151
R652 B.n139 B.n138 10.6151
R653 B.n138 B.n137 10.6151
R654 B.n137 B.n96 10.6151
R655 B.n133 B.n96 10.6151
R656 B.n133 B.n132 10.6151
R657 B.n132 B.n131 10.6151
R658 B.n131 B.n98 10.6151
R659 B.n127 B.n98 10.6151
R660 B.n127 B.n126 10.6151
R661 B.n126 B.n125 10.6151
R662 B.n125 B.n100 10.6151
R663 B.n121 B.n100 10.6151
R664 B.n121 B.n120 10.6151
R665 B.n120 B.n119 10.6151
R666 B.n119 B.n102 10.6151
R667 B.n115 B.n102 10.6151
R668 B.n115 B.n114 10.6151
R669 B.n114 B.n113 10.6151
R670 B.n113 B.n104 10.6151
R671 B.n109 B.n104 10.6151
R672 B.n109 B.n108 10.6151
R673 B.n108 B.n107 10.6151
R674 B.n107 B.n0 10.6151
R675 B.n391 B.n1 10.6151
R676 B.n391 B.n390 10.6151
R677 B.n390 B.n389 10.6151
R678 B.n389 B.n4 10.6151
R679 B.n385 B.n4 10.6151
R680 B.n385 B.n384 10.6151
R681 B.n384 B.n383 10.6151
R682 B.n383 B.n6 10.6151
R683 B.n379 B.n6 10.6151
R684 B.n379 B.n378 10.6151
R685 B.n378 B.n377 10.6151
R686 B.n377 B.n8 10.6151
R687 B.n373 B.n8 10.6151
R688 B.n373 B.n372 10.6151
R689 B.n372 B.n371 10.6151
R690 B.n371 B.n10 10.6151
R691 B.n367 B.n10 10.6151
R692 B.n367 B.n366 10.6151
R693 B.n366 B.n365 10.6151
R694 B.n365 B.n12 10.6151
R695 B.n361 B.n12 10.6151
R696 B.n361 B.n360 10.6151
R697 B.n360 B.n359 10.6151
R698 B.n359 B.n14 10.6151
R699 B.n355 B.n14 10.6151
R700 B.n355 B.n354 10.6151
R701 B.n354 B.n353 10.6151
R702 B.n353 B.n16 10.6151
R703 B.n349 B.n16 10.6151
R704 B.n329 B.n328 6.5566
R705 B.n316 B.n32 6.5566
R706 B.n170 B.n169 6.5566
R707 B.n182 B.n78 6.5566
R708 B.n330 B.n329 4.05904
R709 B.n313 B.n32 4.05904
R710 B.n169 B.n168 4.05904
R711 B.n185 B.n78 4.05904
R712 B.n395 B.n0 2.81026
R713 B.n395 B.n1 2.81026
R714 VN.n16 VN.n15 174.334
R715 VN.n33 VN.n32 174.334
R716 VN.n31 VN.n17 161.3
R717 VN.n30 VN.n29 161.3
R718 VN.n28 VN.n18 161.3
R719 VN.n27 VN.n26 161.3
R720 VN.n25 VN.n19 161.3
R721 VN.n24 VN.n23 161.3
R722 VN.n14 VN.n0 161.3
R723 VN.n13 VN.n12 161.3
R724 VN.n11 VN.n1 161.3
R725 VN.n10 VN.n9 161.3
R726 VN.n7 VN.n2 161.3
R727 VN.n6 VN.n5 161.3
R728 VN.n4 VN.t5 73.7195
R729 VN.n22 VN.t2 73.7195
R730 VN.n4 VN.n3 51.8775
R731 VN.n22 VN.n21 51.8775
R732 VN.n3 VN.t3 44.0453
R733 VN.n8 VN.t0 44.0453
R734 VN.n15 VN.t7 44.0453
R735 VN.n21 VN.t1 44.0453
R736 VN.n20 VN.t6 44.0453
R737 VN.n32 VN.t4 44.0453
R738 VN.n13 VN.n1 41.5458
R739 VN.n30 VN.n18 41.5458
R740 VN.n7 VN.n6 40.577
R741 VN.n9 VN.n7 40.577
R742 VN.n25 VN.n24 40.577
R743 VN.n26 VN.n25 40.577
R744 VN.n14 VN.n13 39.6083
R745 VN.n31 VN.n30 39.6083
R746 VN VN.n33 36.9191
R747 VN.n23 VN.n22 27.1451
R748 VN.n5 VN.n4 27.1451
R749 VN.n8 VN.n1 12.5423
R750 VN.n20 VN.n18 12.5423
R751 VN.n6 VN.n3 12.0505
R752 VN.n9 VN.n8 12.0505
R753 VN.n24 VN.n21 12.0505
R754 VN.n26 VN.n20 12.0505
R755 VN.n15 VN.n14 11.5587
R756 VN.n32 VN.n31 11.5587
R757 VN.n33 VN.n17 0.189894
R758 VN.n29 VN.n17 0.189894
R759 VN.n29 VN.n28 0.189894
R760 VN.n28 VN.n27 0.189894
R761 VN.n27 VN.n19 0.189894
R762 VN.n23 VN.n19 0.189894
R763 VN.n5 VN.n2 0.189894
R764 VN.n10 VN.n2 0.189894
R765 VN.n11 VN.n10 0.189894
R766 VN.n12 VN.n11 0.189894
R767 VN.n12 VN.n0 0.189894
R768 VN.n16 VN.n0 0.189894
R769 VN VN.n16 0.0516364
R770 VDD2.n2 VDD2.n1 172.977
R771 VDD2.n2 VDD2.n0 172.977
R772 VDD2 VDD2.n5 172.975
R773 VDD2.n4 VDD2.n3 172.391
R774 VDD2.n4 VDD2.n2 31.3231
R775 VDD2.n5 VDD2.t6 15.333
R776 VDD2.n5 VDD2.t5 15.333
R777 VDD2.n3 VDD2.t3 15.333
R778 VDD2.n3 VDD2.t1 15.333
R779 VDD2.n1 VDD2.t7 15.333
R780 VDD2.n1 VDD2.t0 15.333
R781 VDD2.n0 VDD2.t2 15.333
R782 VDD2.n0 VDD2.t4 15.333
R783 VDD2 VDD2.n4 0.700931
C0 VDD2 w_n2460_n1392# 1.2473f
C1 B w_n2460_n1392# 5.14614f
C2 VDD2 VN 1.5696f
C3 VP w_n2460_n1392# 4.72467f
C4 B VN 0.76945f
C5 VP VN 4.07952f
C6 w_n2460_n1392# VTAIL 1.72677f
C7 VDD1 VDD2 1.05283f
C8 VN VTAIL 2.0339f
C9 B VDD1 0.943116f
C10 VDD1 VP 1.78616f
C11 B VDD2 0.994224f
C12 VP VDD2 0.372782f
C13 VDD1 VTAIL 3.72375f
C14 VN w_n2460_n1392# 4.41374f
C15 B VP 1.28931f
C16 VDD2 VTAIL 3.76851f
C17 B VTAIL 1.27388f
C18 VDD1 w_n2460_n1392# 1.19386f
C19 VP VTAIL 2.04801f
C20 VDD1 VN 0.154658f
C21 VDD2 VSUBS 0.810383f
C22 VDD1 VSUBS 1.177108f
C23 VTAIL VSUBS 0.40066f
C24 VN VSUBS 4.39869f
C25 VP VSUBS 1.579872f
C26 B VSUBS 2.428747f
C27 w_n2460_n1392# VSUBS 43.660103f
C28 VDD2.t2 VSUBS 0.029717f
C29 VDD2.t4 VSUBS 0.029717f
C30 VDD2.n0 VSUBS 0.136734f
C31 VDD2.t7 VSUBS 0.029717f
C32 VDD2.t0 VSUBS 0.029717f
C33 VDD2.n1 VSUBS 0.136734f
C34 VDD2.n2 VSUBS 1.41049f
C35 VDD2.t3 VSUBS 0.029717f
C36 VDD2.t1 VSUBS 0.029717f
C37 VDD2.n3 VSUBS 0.135692f
C38 VDD2.n4 VSUBS 1.22735f
C39 VDD2.t6 VSUBS 0.029717f
C40 VDD2.t5 VSUBS 0.029717f
C41 VDD2.n5 VSUBS 0.136725f
C42 VN.n0 VSUBS 0.055561f
C43 VN.t7 VSUBS 0.322712f
C44 VN.n1 VSUBS 0.084337f
C45 VN.n2 VSUBS 0.055561f
C46 VN.t3 VSUBS 0.322712f
C47 VN.n3 VSUBS 0.258181f
C48 VN.t5 VSUBS 0.458144f
C49 VN.n4 VSUBS 0.264245f
C50 VN.n5 VSUBS 0.286449f
C51 VN.n6 VSUBS 0.083905f
C52 VN.n7 VSUBS 0.044875f
C53 VN.t0 VSUBS 0.322712f
C54 VN.n8 VSUBS 0.178505f
C55 VN.n9 VSUBS 0.083905f
C56 VN.n10 VSUBS 0.055561f
C57 VN.n11 VSUBS 0.055561f
C58 VN.n12 VSUBS 0.055561f
C59 VN.n13 VSUBS 0.044946f
C60 VN.n14 VSUBS 0.083403f
C61 VN.n15 VSUBS 0.263952f
C62 VN.n16 VSUBS 0.049962f
C63 VN.n17 VSUBS 0.055561f
C64 VN.t4 VSUBS 0.322712f
C65 VN.n18 VSUBS 0.084337f
C66 VN.n19 VSUBS 0.055561f
C67 VN.t6 VSUBS 0.322712f
C68 VN.n20 VSUBS 0.178505f
C69 VN.t1 VSUBS 0.322712f
C70 VN.n21 VSUBS 0.258181f
C71 VN.t2 VSUBS 0.458144f
C72 VN.n22 VSUBS 0.264245f
C73 VN.n23 VSUBS 0.286449f
C74 VN.n24 VSUBS 0.083905f
C75 VN.n25 VSUBS 0.044875f
C76 VN.n26 VSUBS 0.083905f
C77 VN.n27 VSUBS 0.055561f
C78 VN.n28 VSUBS 0.055561f
C79 VN.n29 VSUBS 0.055561f
C80 VN.n30 VSUBS 0.044946f
C81 VN.n31 VSUBS 0.083403f
C82 VN.n32 VSUBS 0.263952f
C83 VN.n33 VSUBS 1.83956f
C84 B.n0 VSUBS 0.005355f
C85 B.n1 VSUBS 0.005355f
C86 B.n2 VSUBS 0.008468f
C87 B.n3 VSUBS 0.008468f
C88 B.n4 VSUBS 0.008468f
C89 B.n5 VSUBS 0.008468f
C90 B.n6 VSUBS 0.008468f
C91 B.n7 VSUBS 0.008468f
C92 B.n8 VSUBS 0.008468f
C93 B.n9 VSUBS 0.008468f
C94 B.n10 VSUBS 0.008468f
C95 B.n11 VSUBS 0.008468f
C96 B.n12 VSUBS 0.008468f
C97 B.n13 VSUBS 0.008468f
C98 B.n14 VSUBS 0.008468f
C99 B.n15 VSUBS 0.008468f
C100 B.n16 VSUBS 0.008468f
C101 B.n17 VSUBS 0.019832f
C102 B.n18 VSUBS 0.008468f
C103 B.n19 VSUBS 0.008468f
C104 B.n20 VSUBS 0.008468f
C105 B.n21 VSUBS 0.008468f
C106 B.n22 VSUBS 0.008468f
C107 B.n23 VSUBS 0.008468f
C108 B.t5 VSUBS 0.056153f
C109 B.t4 VSUBS 0.06369f
C110 B.t3 VSUBS 0.143483f
C111 B.n24 VSUBS 0.072277f
C112 B.n25 VSUBS 0.064436f
C113 B.n26 VSUBS 0.008468f
C114 B.n27 VSUBS 0.008468f
C115 B.n28 VSUBS 0.008468f
C116 B.n29 VSUBS 0.008468f
C117 B.t8 VSUBS 0.056153f
C118 B.t7 VSUBS 0.06369f
C119 B.t6 VSUBS 0.143483f
C120 B.n30 VSUBS 0.072277f
C121 B.n31 VSUBS 0.064436f
C122 B.n32 VSUBS 0.01962f
C123 B.n33 VSUBS 0.008468f
C124 B.n34 VSUBS 0.008468f
C125 B.n35 VSUBS 0.008468f
C126 B.n36 VSUBS 0.008468f
C127 B.n37 VSUBS 0.008468f
C128 B.n38 VSUBS 0.008468f
C129 B.n39 VSUBS 0.018524f
C130 B.n40 VSUBS 0.008468f
C131 B.n41 VSUBS 0.008468f
C132 B.n42 VSUBS 0.008468f
C133 B.n43 VSUBS 0.008468f
C134 B.n44 VSUBS 0.008468f
C135 B.n45 VSUBS 0.008468f
C136 B.n46 VSUBS 0.008468f
C137 B.n47 VSUBS 0.008468f
C138 B.n48 VSUBS 0.008468f
C139 B.n49 VSUBS 0.008468f
C140 B.n50 VSUBS 0.008468f
C141 B.n51 VSUBS 0.008468f
C142 B.n52 VSUBS 0.008468f
C143 B.n53 VSUBS 0.008468f
C144 B.n54 VSUBS 0.008468f
C145 B.n55 VSUBS 0.008468f
C146 B.n56 VSUBS 0.008468f
C147 B.n57 VSUBS 0.008468f
C148 B.n58 VSUBS 0.008468f
C149 B.n59 VSUBS 0.008468f
C150 B.n60 VSUBS 0.008468f
C151 B.n61 VSUBS 0.008468f
C152 B.n62 VSUBS 0.008468f
C153 B.n63 VSUBS 0.008468f
C154 B.n64 VSUBS 0.008468f
C155 B.n65 VSUBS 0.008468f
C156 B.n66 VSUBS 0.008468f
C157 B.n67 VSUBS 0.008468f
C158 B.n68 VSUBS 0.008468f
C159 B.n69 VSUBS 0.018524f
C160 B.n70 VSUBS 0.008468f
C161 B.n71 VSUBS 0.008468f
C162 B.n72 VSUBS 0.008468f
C163 B.n73 VSUBS 0.008468f
C164 B.n74 VSUBS 0.008468f
C165 B.n75 VSUBS 0.008468f
C166 B.t1 VSUBS 0.056153f
C167 B.t2 VSUBS 0.06369f
C168 B.t0 VSUBS 0.143483f
C169 B.n76 VSUBS 0.072277f
C170 B.n77 VSUBS 0.064436f
C171 B.n78 VSUBS 0.01962f
C172 B.n79 VSUBS 0.008468f
C173 B.n80 VSUBS 0.008468f
C174 B.n81 VSUBS 0.008468f
C175 B.n82 VSUBS 0.008468f
C176 B.n83 VSUBS 0.008468f
C177 B.t10 VSUBS 0.056153f
C178 B.t11 VSUBS 0.06369f
C179 B.t9 VSUBS 0.143483f
C180 B.n84 VSUBS 0.072277f
C181 B.n85 VSUBS 0.064436f
C182 B.n86 VSUBS 0.008468f
C183 B.n87 VSUBS 0.008468f
C184 B.n88 VSUBS 0.008468f
C185 B.n89 VSUBS 0.008468f
C186 B.n90 VSUBS 0.008468f
C187 B.n91 VSUBS 0.019832f
C188 B.n92 VSUBS 0.008468f
C189 B.n93 VSUBS 0.008468f
C190 B.n94 VSUBS 0.008468f
C191 B.n95 VSUBS 0.008468f
C192 B.n96 VSUBS 0.008468f
C193 B.n97 VSUBS 0.008468f
C194 B.n98 VSUBS 0.008468f
C195 B.n99 VSUBS 0.008468f
C196 B.n100 VSUBS 0.008468f
C197 B.n101 VSUBS 0.008468f
C198 B.n102 VSUBS 0.008468f
C199 B.n103 VSUBS 0.008468f
C200 B.n104 VSUBS 0.008468f
C201 B.n105 VSUBS 0.008468f
C202 B.n106 VSUBS 0.008468f
C203 B.n107 VSUBS 0.008468f
C204 B.n108 VSUBS 0.008468f
C205 B.n109 VSUBS 0.008468f
C206 B.n110 VSUBS 0.008468f
C207 B.n111 VSUBS 0.008468f
C208 B.n112 VSUBS 0.008468f
C209 B.n113 VSUBS 0.008468f
C210 B.n114 VSUBS 0.008468f
C211 B.n115 VSUBS 0.008468f
C212 B.n116 VSUBS 0.008468f
C213 B.n117 VSUBS 0.008468f
C214 B.n118 VSUBS 0.008468f
C215 B.n119 VSUBS 0.008468f
C216 B.n120 VSUBS 0.008468f
C217 B.n121 VSUBS 0.008468f
C218 B.n122 VSUBS 0.008468f
C219 B.n123 VSUBS 0.008468f
C220 B.n124 VSUBS 0.008468f
C221 B.n125 VSUBS 0.008468f
C222 B.n126 VSUBS 0.008468f
C223 B.n127 VSUBS 0.008468f
C224 B.n128 VSUBS 0.008468f
C225 B.n129 VSUBS 0.008468f
C226 B.n130 VSUBS 0.008468f
C227 B.n131 VSUBS 0.008468f
C228 B.n132 VSUBS 0.008468f
C229 B.n133 VSUBS 0.008468f
C230 B.n134 VSUBS 0.008468f
C231 B.n135 VSUBS 0.008468f
C232 B.n136 VSUBS 0.008468f
C233 B.n137 VSUBS 0.008468f
C234 B.n138 VSUBS 0.008468f
C235 B.n139 VSUBS 0.008468f
C236 B.n140 VSUBS 0.008468f
C237 B.n141 VSUBS 0.008468f
C238 B.n142 VSUBS 0.008468f
C239 B.n143 VSUBS 0.008468f
C240 B.n144 VSUBS 0.008468f
C241 B.n145 VSUBS 0.008468f
C242 B.n146 VSUBS 0.008468f
C243 B.n147 VSUBS 0.008468f
C244 B.n148 VSUBS 0.018524f
C245 B.n149 VSUBS 0.018524f
C246 B.n150 VSUBS 0.019832f
C247 B.n151 VSUBS 0.008468f
C248 B.n152 VSUBS 0.008468f
C249 B.n153 VSUBS 0.008468f
C250 B.n154 VSUBS 0.008468f
C251 B.n155 VSUBS 0.008468f
C252 B.n156 VSUBS 0.008468f
C253 B.n157 VSUBS 0.008468f
C254 B.n158 VSUBS 0.008468f
C255 B.n159 VSUBS 0.008468f
C256 B.n160 VSUBS 0.008468f
C257 B.n161 VSUBS 0.008468f
C258 B.n162 VSUBS 0.008468f
C259 B.n163 VSUBS 0.008468f
C260 B.n164 VSUBS 0.008468f
C261 B.n165 VSUBS 0.008468f
C262 B.n166 VSUBS 0.008468f
C263 B.n167 VSUBS 0.008468f
C264 B.n168 VSUBS 0.005853f
C265 B.n169 VSUBS 0.01962f
C266 B.n170 VSUBS 0.006849f
C267 B.n171 VSUBS 0.008468f
C268 B.n172 VSUBS 0.008468f
C269 B.n173 VSUBS 0.008468f
C270 B.n174 VSUBS 0.008468f
C271 B.n175 VSUBS 0.008468f
C272 B.n176 VSUBS 0.008468f
C273 B.n177 VSUBS 0.008468f
C274 B.n178 VSUBS 0.008468f
C275 B.n179 VSUBS 0.008468f
C276 B.n180 VSUBS 0.008468f
C277 B.n181 VSUBS 0.008468f
C278 B.n182 VSUBS 0.006849f
C279 B.n183 VSUBS 0.008468f
C280 B.n184 VSUBS 0.008468f
C281 B.n185 VSUBS 0.005853f
C282 B.n186 VSUBS 0.008468f
C283 B.n187 VSUBS 0.008468f
C284 B.n188 VSUBS 0.008468f
C285 B.n189 VSUBS 0.008468f
C286 B.n190 VSUBS 0.008468f
C287 B.n191 VSUBS 0.008468f
C288 B.n192 VSUBS 0.008468f
C289 B.n193 VSUBS 0.008468f
C290 B.n194 VSUBS 0.008468f
C291 B.n195 VSUBS 0.008468f
C292 B.n196 VSUBS 0.008468f
C293 B.n197 VSUBS 0.008468f
C294 B.n198 VSUBS 0.008468f
C295 B.n199 VSUBS 0.008468f
C296 B.n200 VSUBS 0.008468f
C297 B.n201 VSUBS 0.008468f
C298 B.n202 VSUBS 0.019832f
C299 B.n203 VSUBS 0.019832f
C300 B.n204 VSUBS 0.018524f
C301 B.n205 VSUBS 0.008468f
C302 B.n206 VSUBS 0.008468f
C303 B.n207 VSUBS 0.008468f
C304 B.n208 VSUBS 0.008468f
C305 B.n209 VSUBS 0.008468f
C306 B.n210 VSUBS 0.008468f
C307 B.n211 VSUBS 0.008468f
C308 B.n212 VSUBS 0.008468f
C309 B.n213 VSUBS 0.008468f
C310 B.n214 VSUBS 0.008468f
C311 B.n215 VSUBS 0.008468f
C312 B.n216 VSUBS 0.008468f
C313 B.n217 VSUBS 0.008468f
C314 B.n218 VSUBS 0.008468f
C315 B.n219 VSUBS 0.008468f
C316 B.n220 VSUBS 0.008468f
C317 B.n221 VSUBS 0.008468f
C318 B.n222 VSUBS 0.008468f
C319 B.n223 VSUBS 0.008468f
C320 B.n224 VSUBS 0.008468f
C321 B.n225 VSUBS 0.008468f
C322 B.n226 VSUBS 0.008468f
C323 B.n227 VSUBS 0.008468f
C324 B.n228 VSUBS 0.008468f
C325 B.n229 VSUBS 0.008468f
C326 B.n230 VSUBS 0.008468f
C327 B.n231 VSUBS 0.008468f
C328 B.n232 VSUBS 0.008468f
C329 B.n233 VSUBS 0.008468f
C330 B.n234 VSUBS 0.008468f
C331 B.n235 VSUBS 0.008468f
C332 B.n236 VSUBS 0.008468f
C333 B.n237 VSUBS 0.008468f
C334 B.n238 VSUBS 0.008468f
C335 B.n239 VSUBS 0.008468f
C336 B.n240 VSUBS 0.008468f
C337 B.n241 VSUBS 0.008468f
C338 B.n242 VSUBS 0.008468f
C339 B.n243 VSUBS 0.008468f
C340 B.n244 VSUBS 0.008468f
C341 B.n245 VSUBS 0.008468f
C342 B.n246 VSUBS 0.008468f
C343 B.n247 VSUBS 0.008468f
C344 B.n248 VSUBS 0.008468f
C345 B.n249 VSUBS 0.008468f
C346 B.n250 VSUBS 0.008468f
C347 B.n251 VSUBS 0.008468f
C348 B.n252 VSUBS 0.008468f
C349 B.n253 VSUBS 0.008468f
C350 B.n254 VSUBS 0.008468f
C351 B.n255 VSUBS 0.008468f
C352 B.n256 VSUBS 0.008468f
C353 B.n257 VSUBS 0.008468f
C354 B.n258 VSUBS 0.008468f
C355 B.n259 VSUBS 0.008468f
C356 B.n260 VSUBS 0.008468f
C357 B.n261 VSUBS 0.008468f
C358 B.n262 VSUBS 0.008468f
C359 B.n263 VSUBS 0.008468f
C360 B.n264 VSUBS 0.008468f
C361 B.n265 VSUBS 0.008468f
C362 B.n266 VSUBS 0.008468f
C363 B.n267 VSUBS 0.008468f
C364 B.n268 VSUBS 0.008468f
C365 B.n269 VSUBS 0.008468f
C366 B.n270 VSUBS 0.008468f
C367 B.n271 VSUBS 0.008468f
C368 B.n272 VSUBS 0.008468f
C369 B.n273 VSUBS 0.008468f
C370 B.n274 VSUBS 0.008468f
C371 B.n275 VSUBS 0.008468f
C372 B.n276 VSUBS 0.008468f
C373 B.n277 VSUBS 0.008468f
C374 B.n278 VSUBS 0.008468f
C375 B.n279 VSUBS 0.008468f
C376 B.n280 VSUBS 0.008468f
C377 B.n281 VSUBS 0.008468f
C378 B.n282 VSUBS 0.008468f
C379 B.n283 VSUBS 0.008468f
C380 B.n284 VSUBS 0.008468f
C381 B.n285 VSUBS 0.008468f
C382 B.n286 VSUBS 0.008468f
C383 B.n287 VSUBS 0.008468f
C384 B.n288 VSUBS 0.008468f
C385 B.n289 VSUBS 0.008468f
C386 B.n290 VSUBS 0.008468f
C387 B.n291 VSUBS 0.008468f
C388 B.n292 VSUBS 0.008468f
C389 B.n293 VSUBS 0.008468f
C390 B.n294 VSUBS 0.019576f
C391 B.n295 VSUBS 0.01878f
C392 B.n296 VSUBS 0.019832f
C393 B.n297 VSUBS 0.008468f
C394 B.n298 VSUBS 0.008468f
C395 B.n299 VSUBS 0.008468f
C396 B.n300 VSUBS 0.008468f
C397 B.n301 VSUBS 0.008468f
C398 B.n302 VSUBS 0.008468f
C399 B.n303 VSUBS 0.008468f
C400 B.n304 VSUBS 0.008468f
C401 B.n305 VSUBS 0.008468f
C402 B.n306 VSUBS 0.008468f
C403 B.n307 VSUBS 0.008468f
C404 B.n308 VSUBS 0.008468f
C405 B.n309 VSUBS 0.008468f
C406 B.n310 VSUBS 0.008468f
C407 B.n311 VSUBS 0.008468f
C408 B.n312 VSUBS 0.008468f
C409 B.n313 VSUBS 0.005853f
C410 B.n314 VSUBS 0.008468f
C411 B.n315 VSUBS 0.008468f
C412 B.n316 VSUBS 0.006849f
C413 B.n317 VSUBS 0.008468f
C414 B.n318 VSUBS 0.008468f
C415 B.n319 VSUBS 0.008468f
C416 B.n320 VSUBS 0.008468f
C417 B.n321 VSUBS 0.008468f
C418 B.n322 VSUBS 0.008468f
C419 B.n323 VSUBS 0.008468f
C420 B.n324 VSUBS 0.008468f
C421 B.n325 VSUBS 0.008468f
C422 B.n326 VSUBS 0.008468f
C423 B.n327 VSUBS 0.008468f
C424 B.n328 VSUBS 0.006849f
C425 B.n329 VSUBS 0.01962f
C426 B.n330 VSUBS 0.005853f
C427 B.n331 VSUBS 0.008468f
C428 B.n332 VSUBS 0.008468f
C429 B.n333 VSUBS 0.008468f
C430 B.n334 VSUBS 0.008468f
C431 B.n335 VSUBS 0.008468f
C432 B.n336 VSUBS 0.008468f
C433 B.n337 VSUBS 0.008468f
C434 B.n338 VSUBS 0.008468f
C435 B.n339 VSUBS 0.008468f
C436 B.n340 VSUBS 0.008468f
C437 B.n341 VSUBS 0.008468f
C438 B.n342 VSUBS 0.008468f
C439 B.n343 VSUBS 0.008468f
C440 B.n344 VSUBS 0.008468f
C441 B.n345 VSUBS 0.008468f
C442 B.n346 VSUBS 0.008468f
C443 B.n347 VSUBS 0.008468f
C444 B.n348 VSUBS 0.019832f
C445 B.n349 VSUBS 0.018524f
C446 B.n350 VSUBS 0.018524f
C447 B.n351 VSUBS 0.008468f
C448 B.n352 VSUBS 0.008468f
C449 B.n353 VSUBS 0.008468f
C450 B.n354 VSUBS 0.008468f
C451 B.n355 VSUBS 0.008468f
C452 B.n356 VSUBS 0.008468f
C453 B.n357 VSUBS 0.008468f
C454 B.n358 VSUBS 0.008468f
C455 B.n359 VSUBS 0.008468f
C456 B.n360 VSUBS 0.008468f
C457 B.n361 VSUBS 0.008468f
C458 B.n362 VSUBS 0.008468f
C459 B.n363 VSUBS 0.008468f
C460 B.n364 VSUBS 0.008468f
C461 B.n365 VSUBS 0.008468f
C462 B.n366 VSUBS 0.008468f
C463 B.n367 VSUBS 0.008468f
C464 B.n368 VSUBS 0.008468f
C465 B.n369 VSUBS 0.008468f
C466 B.n370 VSUBS 0.008468f
C467 B.n371 VSUBS 0.008468f
C468 B.n372 VSUBS 0.008468f
C469 B.n373 VSUBS 0.008468f
C470 B.n374 VSUBS 0.008468f
C471 B.n375 VSUBS 0.008468f
C472 B.n376 VSUBS 0.008468f
C473 B.n377 VSUBS 0.008468f
C474 B.n378 VSUBS 0.008468f
C475 B.n379 VSUBS 0.008468f
C476 B.n380 VSUBS 0.008468f
C477 B.n381 VSUBS 0.008468f
C478 B.n382 VSUBS 0.008468f
C479 B.n383 VSUBS 0.008468f
C480 B.n384 VSUBS 0.008468f
C481 B.n385 VSUBS 0.008468f
C482 B.n386 VSUBS 0.008468f
C483 B.n387 VSUBS 0.008468f
C484 B.n388 VSUBS 0.008468f
C485 B.n389 VSUBS 0.008468f
C486 B.n390 VSUBS 0.008468f
C487 B.n391 VSUBS 0.008468f
C488 B.n392 VSUBS 0.008468f
C489 B.n393 VSUBS 0.008468f
C490 B.n394 VSUBS 0.008468f
C491 B.n395 VSUBS 0.019175f
C492 VDD1.t5 VSUBS 0.028445f
C493 VDD1.t7 VSUBS 0.028445f
C494 VDD1.n0 VSUBS 0.131094f
C495 VDD1.t2 VSUBS 0.028445f
C496 VDD1.t1 VSUBS 0.028445f
C497 VDD1.n1 VSUBS 0.130879f
C498 VDD1.t6 VSUBS 0.028445f
C499 VDD1.t3 VSUBS 0.028445f
C500 VDD1.n2 VSUBS 0.130879f
C501 VDD1.n3 VSUBS 1.38624f
C502 VDD1.t0 VSUBS 0.028445f
C503 VDD1.t4 VSUBS 0.028445f
C504 VDD1.n4 VSUBS 0.129882f
C505 VDD1.n5 VSUBS 1.195f
C506 VTAIL.t3 VSUBS 0.045633f
C507 VTAIL.t4 VSUBS 0.045633f
C508 VTAIL.n0 VSUBS 0.177306f
C509 VTAIL.n1 VSUBS 0.407033f
C510 VTAIL.t0 VSUBS 0.2788f
C511 VTAIL.n2 VSUBS 0.466122f
C512 VTAIL.t10 VSUBS 0.2788f
C513 VTAIL.n3 VSUBS 0.466122f
C514 VTAIL.t11 VSUBS 0.045633f
C515 VTAIL.t14 VSUBS 0.045633f
C516 VTAIL.n4 VSUBS 0.177306f
C517 VTAIL.n5 VSUBS 0.514665f
C518 VTAIL.t8 VSUBS 0.2788f
C519 VTAIL.n6 VSUBS 1.06804f
C520 VTAIL.t5 VSUBS 0.278801f
C521 VTAIL.n7 VSUBS 1.06804f
C522 VTAIL.t2 VSUBS 0.045633f
C523 VTAIL.t6 VSUBS 0.045633f
C524 VTAIL.n8 VSUBS 0.177307f
C525 VTAIL.n9 VSUBS 0.514664f
C526 VTAIL.t1 VSUBS 0.278801f
C527 VTAIL.n10 VSUBS 0.466121f
C528 VTAIL.t15 VSUBS 0.278801f
C529 VTAIL.n11 VSUBS 0.466121f
C530 VTAIL.t9 VSUBS 0.045633f
C531 VTAIL.t13 VSUBS 0.045633f
C532 VTAIL.n12 VSUBS 0.177307f
C533 VTAIL.n13 VSUBS 0.514664f
C534 VTAIL.t12 VSUBS 0.2788f
C535 VTAIL.n14 VSUBS 1.06804f
C536 VTAIL.t7 VSUBS 0.2788f
C537 VTAIL.n15 VSUBS 1.06293f
C538 VP.n0 VSUBS 0.057577f
C539 VP.t4 VSUBS 0.33442f
C540 VP.n1 VSUBS 0.087396f
C541 VP.n2 VSUBS 0.057577f
C542 VP.t6 VSUBS 0.33442f
C543 VP.n3 VSUBS 0.184981f
C544 VP.n4 VSUBS 0.057577f
C545 VP.t5 VSUBS 0.33442f
C546 VP.n5 VSUBS 0.273528f
C547 VP.n6 VSUBS 0.057577f
C548 VP.t3 VSUBS 0.33442f
C549 VP.n7 VSUBS 0.087396f
C550 VP.n8 VSUBS 0.057577f
C551 VP.t0 VSUBS 0.33442f
C552 VP.n9 VSUBS 0.267548f
C553 VP.t2 VSUBS 0.474766f
C554 VP.n10 VSUBS 0.273831f
C555 VP.n11 VSUBS 0.296841f
C556 VP.n12 VSUBS 0.086949f
C557 VP.n13 VSUBS 0.046503f
C558 VP.t7 VSUBS 0.33442f
C559 VP.n14 VSUBS 0.184981f
C560 VP.n15 VSUBS 0.086949f
C561 VP.n16 VSUBS 0.057577f
C562 VP.n17 VSUBS 0.057577f
C563 VP.n18 VSUBS 0.057577f
C564 VP.n19 VSUBS 0.046576f
C565 VP.n20 VSUBS 0.086429f
C566 VP.n21 VSUBS 0.273528f
C567 VP.n22 VSUBS 1.86815f
C568 VP.n23 VSUBS 1.92496f
C569 VP.n24 VSUBS 0.057577f
C570 VP.n25 VSUBS 0.086429f
C571 VP.n26 VSUBS 0.046576f
C572 VP.n27 VSUBS 0.087396f
C573 VP.n28 VSUBS 0.057577f
C574 VP.n29 VSUBS 0.057577f
C575 VP.n30 VSUBS 0.086949f
C576 VP.n31 VSUBS 0.046503f
C577 VP.t1 VSUBS 0.33442f
C578 VP.n32 VSUBS 0.184981f
C579 VP.n33 VSUBS 0.086949f
C580 VP.n34 VSUBS 0.057577f
C581 VP.n35 VSUBS 0.057577f
C582 VP.n36 VSUBS 0.057577f
C583 VP.n37 VSUBS 0.046576f
C584 VP.n38 VSUBS 0.086429f
C585 VP.n39 VSUBS 0.273528f
C586 VP.n40 VSUBS 0.051775f
.ends

