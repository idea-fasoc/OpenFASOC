* NGSPICE file created from diff_pair_sample_0467.ext - technology: sky130A

.subckt diff_pair_sample_0467 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=5.3508 pd=28.22 as=0 ps=0 w=13.72 l=0.75
X1 VTAIL.t7 VN.t0 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=5.3508 pd=28.22 as=2.2638 ps=14.05 w=13.72 l=0.75
X2 VDD1.t3 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2638 pd=14.05 as=5.3508 ps=28.22 w=13.72 l=0.75
X3 VDD2.t1 VN.t1 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.2638 pd=14.05 as=5.3508 ps=28.22 w=13.72 l=0.75
X4 VDD1.t2 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.2638 pd=14.05 as=5.3508 ps=28.22 w=13.72 l=0.75
X5 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=5.3508 pd=28.22 as=0 ps=0 w=13.72 l=0.75
X6 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.3508 pd=28.22 as=0 ps=0 w=13.72 l=0.75
X7 VDD2.t2 VN.t2 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2638 pd=14.05 as=5.3508 ps=28.22 w=13.72 l=0.75
X8 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.3508 pd=28.22 as=0 ps=0 w=13.72 l=0.75
X9 VTAIL.t4 VN.t3 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=5.3508 pd=28.22 as=2.2638 ps=14.05 w=13.72 l=0.75
X10 VTAIL.t3 VP.t2 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=5.3508 pd=28.22 as=2.2638 ps=14.05 w=13.72 l=0.75
X11 VTAIL.t0 VP.t3 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.3508 pd=28.22 as=2.2638 ps=14.05 w=13.72 l=0.75
R0 B.n91 B.t15 643.26
R1 B.n88 B.t4 643.26
R2 B.n384 B.t12 643.26
R3 B.n381 B.t8 643.26
R4 B.n668 B.n667 585
R5 B.n669 B.n668 585
R6 B.n296 B.n87 585
R7 B.n295 B.n294 585
R8 B.n293 B.n292 585
R9 B.n291 B.n290 585
R10 B.n289 B.n288 585
R11 B.n287 B.n286 585
R12 B.n285 B.n284 585
R13 B.n283 B.n282 585
R14 B.n281 B.n280 585
R15 B.n279 B.n278 585
R16 B.n277 B.n276 585
R17 B.n275 B.n274 585
R18 B.n273 B.n272 585
R19 B.n271 B.n270 585
R20 B.n269 B.n268 585
R21 B.n267 B.n266 585
R22 B.n265 B.n264 585
R23 B.n263 B.n262 585
R24 B.n261 B.n260 585
R25 B.n259 B.n258 585
R26 B.n257 B.n256 585
R27 B.n255 B.n254 585
R28 B.n253 B.n252 585
R29 B.n251 B.n250 585
R30 B.n249 B.n248 585
R31 B.n247 B.n246 585
R32 B.n245 B.n244 585
R33 B.n243 B.n242 585
R34 B.n241 B.n240 585
R35 B.n239 B.n238 585
R36 B.n237 B.n236 585
R37 B.n235 B.n234 585
R38 B.n233 B.n232 585
R39 B.n231 B.n230 585
R40 B.n229 B.n228 585
R41 B.n227 B.n226 585
R42 B.n225 B.n224 585
R43 B.n223 B.n222 585
R44 B.n221 B.n220 585
R45 B.n219 B.n218 585
R46 B.n217 B.n216 585
R47 B.n215 B.n214 585
R48 B.n213 B.n212 585
R49 B.n211 B.n210 585
R50 B.n209 B.n208 585
R51 B.n207 B.n206 585
R52 B.n205 B.n204 585
R53 B.n203 B.n202 585
R54 B.n201 B.n200 585
R55 B.n199 B.n198 585
R56 B.n197 B.n196 585
R57 B.n195 B.n194 585
R58 B.n193 B.n192 585
R59 B.n191 B.n190 585
R60 B.n189 B.n188 585
R61 B.n186 B.n185 585
R62 B.n184 B.n183 585
R63 B.n182 B.n181 585
R64 B.n180 B.n179 585
R65 B.n178 B.n177 585
R66 B.n176 B.n175 585
R67 B.n174 B.n173 585
R68 B.n172 B.n171 585
R69 B.n170 B.n169 585
R70 B.n168 B.n167 585
R71 B.n166 B.n165 585
R72 B.n164 B.n163 585
R73 B.n162 B.n161 585
R74 B.n160 B.n159 585
R75 B.n158 B.n157 585
R76 B.n156 B.n155 585
R77 B.n154 B.n153 585
R78 B.n152 B.n151 585
R79 B.n150 B.n149 585
R80 B.n148 B.n147 585
R81 B.n146 B.n145 585
R82 B.n144 B.n143 585
R83 B.n142 B.n141 585
R84 B.n140 B.n139 585
R85 B.n138 B.n137 585
R86 B.n136 B.n135 585
R87 B.n134 B.n133 585
R88 B.n132 B.n131 585
R89 B.n130 B.n129 585
R90 B.n128 B.n127 585
R91 B.n126 B.n125 585
R92 B.n124 B.n123 585
R93 B.n122 B.n121 585
R94 B.n120 B.n119 585
R95 B.n118 B.n117 585
R96 B.n116 B.n115 585
R97 B.n114 B.n113 585
R98 B.n112 B.n111 585
R99 B.n110 B.n109 585
R100 B.n108 B.n107 585
R101 B.n106 B.n105 585
R102 B.n104 B.n103 585
R103 B.n102 B.n101 585
R104 B.n100 B.n99 585
R105 B.n98 B.n97 585
R106 B.n96 B.n95 585
R107 B.n94 B.n93 585
R108 B.n666 B.n35 585
R109 B.n670 B.n35 585
R110 B.n665 B.n34 585
R111 B.n671 B.n34 585
R112 B.n664 B.n663 585
R113 B.n663 B.n30 585
R114 B.n662 B.n29 585
R115 B.n677 B.n29 585
R116 B.n661 B.n28 585
R117 B.n678 B.n28 585
R118 B.n660 B.n27 585
R119 B.n679 B.n27 585
R120 B.n659 B.n658 585
R121 B.n658 B.n23 585
R122 B.n657 B.n22 585
R123 B.n685 B.n22 585
R124 B.n656 B.n21 585
R125 B.n686 B.n21 585
R126 B.n655 B.n20 585
R127 B.n687 B.n20 585
R128 B.n654 B.n653 585
R129 B.n653 B.n16 585
R130 B.n652 B.n15 585
R131 B.n693 B.n15 585
R132 B.n651 B.n14 585
R133 B.n694 B.n14 585
R134 B.n650 B.n13 585
R135 B.n695 B.n13 585
R136 B.n649 B.n648 585
R137 B.n648 B.n12 585
R138 B.n647 B.n646 585
R139 B.n647 B.n8 585
R140 B.n645 B.n7 585
R141 B.n702 B.n7 585
R142 B.n644 B.n6 585
R143 B.n703 B.n6 585
R144 B.n643 B.n5 585
R145 B.n704 B.n5 585
R146 B.n642 B.n641 585
R147 B.n641 B.n4 585
R148 B.n640 B.n297 585
R149 B.n640 B.n639 585
R150 B.n629 B.n298 585
R151 B.n632 B.n298 585
R152 B.n631 B.n630 585
R153 B.n633 B.n631 585
R154 B.n628 B.n303 585
R155 B.n303 B.n302 585
R156 B.n627 B.n626 585
R157 B.n626 B.n625 585
R158 B.n305 B.n304 585
R159 B.n306 B.n305 585
R160 B.n618 B.n617 585
R161 B.n619 B.n618 585
R162 B.n616 B.n311 585
R163 B.n311 B.n310 585
R164 B.n615 B.n614 585
R165 B.n614 B.n613 585
R166 B.n313 B.n312 585
R167 B.n314 B.n313 585
R168 B.n606 B.n605 585
R169 B.n607 B.n606 585
R170 B.n604 B.n318 585
R171 B.n322 B.n318 585
R172 B.n603 B.n602 585
R173 B.n602 B.n601 585
R174 B.n320 B.n319 585
R175 B.n321 B.n320 585
R176 B.n594 B.n593 585
R177 B.n595 B.n594 585
R178 B.n592 B.n327 585
R179 B.n327 B.n326 585
R180 B.n586 B.n585 585
R181 B.n584 B.n380 585
R182 B.n583 B.n379 585
R183 B.n588 B.n379 585
R184 B.n582 B.n581 585
R185 B.n580 B.n579 585
R186 B.n578 B.n577 585
R187 B.n576 B.n575 585
R188 B.n574 B.n573 585
R189 B.n572 B.n571 585
R190 B.n570 B.n569 585
R191 B.n568 B.n567 585
R192 B.n566 B.n565 585
R193 B.n564 B.n563 585
R194 B.n562 B.n561 585
R195 B.n560 B.n559 585
R196 B.n558 B.n557 585
R197 B.n556 B.n555 585
R198 B.n554 B.n553 585
R199 B.n552 B.n551 585
R200 B.n550 B.n549 585
R201 B.n548 B.n547 585
R202 B.n546 B.n545 585
R203 B.n544 B.n543 585
R204 B.n542 B.n541 585
R205 B.n540 B.n539 585
R206 B.n538 B.n537 585
R207 B.n536 B.n535 585
R208 B.n534 B.n533 585
R209 B.n532 B.n531 585
R210 B.n530 B.n529 585
R211 B.n528 B.n527 585
R212 B.n526 B.n525 585
R213 B.n524 B.n523 585
R214 B.n522 B.n521 585
R215 B.n520 B.n519 585
R216 B.n518 B.n517 585
R217 B.n516 B.n515 585
R218 B.n514 B.n513 585
R219 B.n512 B.n511 585
R220 B.n510 B.n509 585
R221 B.n508 B.n507 585
R222 B.n506 B.n505 585
R223 B.n504 B.n503 585
R224 B.n502 B.n501 585
R225 B.n500 B.n499 585
R226 B.n498 B.n497 585
R227 B.n496 B.n495 585
R228 B.n494 B.n493 585
R229 B.n492 B.n491 585
R230 B.n490 B.n489 585
R231 B.n488 B.n487 585
R232 B.n486 B.n485 585
R233 B.n484 B.n483 585
R234 B.n482 B.n481 585
R235 B.n480 B.n479 585
R236 B.n478 B.n477 585
R237 B.n475 B.n474 585
R238 B.n473 B.n472 585
R239 B.n471 B.n470 585
R240 B.n469 B.n468 585
R241 B.n467 B.n466 585
R242 B.n465 B.n464 585
R243 B.n463 B.n462 585
R244 B.n461 B.n460 585
R245 B.n459 B.n458 585
R246 B.n457 B.n456 585
R247 B.n455 B.n454 585
R248 B.n453 B.n452 585
R249 B.n451 B.n450 585
R250 B.n449 B.n448 585
R251 B.n447 B.n446 585
R252 B.n445 B.n444 585
R253 B.n443 B.n442 585
R254 B.n441 B.n440 585
R255 B.n439 B.n438 585
R256 B.n437 B.n436 585
R257 B.n435 B.n434 585
R258 B.n433 B.n432 585
R259 B.n431 B.n430 585
R260 B.n429 B.n428 585
R261 B.n427 B.n426 585
R262 B.n425 B.n424 585
R263 B.n423 B.n422 585
R264 B.n421 B.n420 585
R265 B.n419 B.n418 585
R266 B.n417 B.n416 585
R267 B.n415 B.n414 585
R268 B.n413 B.n412 585
R269 B.n411 B.n410 585
R270 B.n409 B.n408 585
R271 B.n407 B.n406 585
R272 B.n405 B.n404 585
R273 B.n403 B.n402 585
R274 B.n401 B.n400 585
R275 B.n399 B.n398 585
R276 B.n397 B.n396 585
R277 B.n395 B.n394 585
R278 B.n393 B.n392 585
R279 B.n391 B.n390 585
R280 B.n389 B.n388 585
R281 B.n387 B.n386 585
R282 B.n329 B.n328 585
R283 B.n591 B.n590 585
R284 B.n325 B.n324 585
R285 B.n326 B.n325 585
R286 B.n597 B.n596 585
R287 B.n596 B.n595 585
R288 B.n598 B.n323 585
R289 B.n323 B.n321 585
R290 B.n600 B.n599 585
R291 B.n601 B.n600 585
R292 B.n317 B.n316 585
R293 B.n322 B.n317 585
R294 B.n609 B.n608 585
R295 B.n608 B.n607 585
R296 B.n610 B.n315 585
R297 B.n315 B.n314 585
R298 B.n612 B.n611 585
R299 B.n613 B.n612 585
R300 B.n309 B.n308 585
R301 B.n310 B.n309 585
R302 B.n621 B.n620 585
R303 B.n620 B.n619 585
R304 B.n622 B.n307 585
R305 B.n307 B.n306 585
R306 B.n624 B.n623 585
R307 B.n625 B.n624 585
R308 B.n301 B.n300 585
R309 B.n302 B.n301 585
R310 B.n635 B.n634 585
R311 B.n634 B.n633 585
R312 B.n636 B.n299 585
R313 B.n632 B.n299 585
R314 B.n638 B.n637 585
R315 B.n639 B.n638 585
R316 B.n3 B.n0 585
R317 B.n4 B.n3 585
R318 B.n701 B.n1 585
R319 B.n702 B.n701 585
R320 B.n700 B.n699 585
R321 B.n700 B.n8 585
R322 B.n698 B.n9 585
R323 B.n12 B.n9 585
R324 B.n697 B.n696 585
R325 B.n696 B.n695 585
R326 B.n11 B.n10 585
R327 B.n694 B.n11 585
R328 B.n692 B.n691 585
R329 B.n693 B.n692 585
R330 B.n690 B.n17 585
R331 B.n17 B.n16 585
R332 B.n689 B.n688 585
R333 B.n688 B.n687 585
R334 B.n19 B.n18 585
R335 B.n686 B.n19 585
R336 B.n684 B.n683 585
R337 B.n685 B.n684 585
R338 B.n682 B.n24 585
R339 B.n24 B.n23 585
R340 B.n681 B.n680 585
R341 B.n680 B.n679 585
R342 B.n26 B.n25 585
R343 B.n678 B.n26 585
R344 B.n676 B.n675 585
R345 B.n677 B.n676 585
R346 B.n674 B.n31 585
R347 B.n31 B.n30 585
R348 B.n673 B.n672 585
R349 B.n672 B.n671 585
R350 B.n33 B.n32 585
R351 B.n670 B.n33 585
R352 B.n705 B.n704 585
R353 B.n703 B.n2 585
R354 B.n93 B.n33 516.524
R355 B.n668 B.n35 516.524
R356 B.n590 B.n327 516.524
R357 B.n586 B.n325 516.524
R358 B.n669 B.n86 256.663
R359 B.n669 B.n85 256.663
R360 B.n669 B.n84 256.663
R361 B.n669 B.n83 256.663
R362 B.n669 B.n82 256.663
R363 B.n669 B.n81 256.663
R364 B.n669 B.n80 256.663
R365 B.n669 B.n79 256.663
R366 B.n669 B.n78 256.663
R367 B.n669 B.n77 256.663
R368 B.n669 B.n76 256.663
R369 B.n669 B.n75 256.663
R370 B.n669 B.n74 256.663
R371 B.n669 B.n73 256.663
R372 B.n669 B.n72 256.663
R373 B.n669 B.n71 256.663
R374 B.n669 B.n70 256.663
R375 B.n669 B.n69 256.663
R376 B.n669 B.n68 256.663
R377 B.n669 B.n67 256.663
R378 B.n669 B.n66 256.663
R379 B.n669 B.n65 256.663
R380 B.n669 B.n64 256.663
R381 B.n669 B.n63 256.663
R382 B.n669 B.n62 256.663
R383 B.n669 B.n61 256.663
R384 B.n669 B.n60 256.663
R385 B.n669 B.n59 256.663
R386 B.n669 B.n58 256.663
R387 B.n669 B.n57 256.663
R388 B.n669 B.n56 256.663
R389 B.n669 B.n55 256.663
R390 B.n669 B.n54 256.663
R391 B.n669 B.n53 256.663
R392 B.n669 B.n52 256.663
R393 B.n669 B.n51 256.663
R394 B.n669 B.n50 256.663
R395 B.n669 B.n49 256.663
R396 B.n669 B.n48 256.663
R397 B.n669 B.n47 256.663
R398 B.n669 B.n46 256.663
R399 B.n669 B.n45 256.663
R400 B.n669 B.n44 256.663
R401 B.n669 B.n43 256.663
R402 B.n669 B.n42 256.663
R403 B.n669 B.n41 256.663
R404 B.n669 B.n40 256.663
R405 B.n669 B.n39 256.663
R406 B.n669 B.n38 256.663
R407 B.n669 B.n37 256.663
R408 B.n669 B.n36 256.663
R409 B.n588 B.n587 256.663
R410 B.n588 B.n330 256.663
R411 B.n588 B.n331 256.663
R412 B.n588 B.n332 256.663
R413 B.n588 B.n333 256.663
R414 B.n588 B.n334 256.663
R415 B.n588 B.n335 256.663
R416 B.n588 B.n336 256.663
R417 B.n588 B.n337 256.663
R418 B.n588 B.n338 256.663
R419 B.n588 B.n339 256.663
R420 B.n588 B.n340 256.663
R421 B.n588 B.n341 256.663
R422 B.n588 B.n342 256.663
R423 B.n588 B.n343 256.663
R424 B.n588 B.n344 256.663
R425 B.n588 B.n345 256.663
R426 B.n588 B.n346 256.663
R427 B.n588 B.n347 256.663
R428 B.n588 B.n348 256.663
R429 B.n588 B.n349 256.663
R430 B.n588 B.n350 256.663
R431 B.n588 B.n351 256.663
R432 B.n588 B.n352 256.663
R433 B.n588 B.n353 256.663
R434 B.n588 B.n354 256.663
R435 B.n588 B.n355 256.663
R436 B.n588 B.n356 256.663
R437 B.n588 B.n357 256.663
R438 B.n588 B.n358 256.663
R439 B.n588 B.n359 256.663
R440 B.n588 B.n360 256.663
R441 B.n588 B.n361 256.663
R442 B.n588 B.n362 256.663
R443 B.n588 B.n363 256.663
R444 B.n588 B.n364 256.663
R445 B.n588 B.n365 256.663
R446 B.n588 B.n366 256.663
R447 B.n588 B.n367 256.663
R448 B.n588 B.n368 256.663
R449 B.n588 B.n369 256.663
R450 B.n588 B.n370 256.663
R451 B.n588 B.n371 256.663
R452 B.n588 B.n372 256.663
R453 B.n588 B.n373 256.663
R454 B.n588 B.n374 256.663
R455 B.n588 B.n375 256.663
R456 B.n588 B.n376 256.663
R457 B.n588 B.n377 256.663
R458 B.n588 B.n378 256.663
R459 B.n589 B.n588 256.663
R460 B.n707 B.n706 256.663
R461 B.n97 B.n96 163.367
R462 B.n101 B.n100 163.367
R463 B.n105 B.n104 163.367
R464 B.n109 B.n108 163.367
R465 B.n113 B.n112 163.367
R466 B.n117 B.n116 163.367
R467 B.n121 B.n120 163.367
R468 B.n125 B.n124 163.367
R469 B.n129 B.n128 163.367
R470 B.n133 B.n132 163.367
R471 B.n137 B.n136 163.367
R472 B.n141 B.n140 163.367
R473 B.n145 B.n144 163.367
R474 B.n149 B.n148 163.367
R475 B.n153 B.n152 163.367
R476 B.n157 B.n156 163.367
R477 B.n161 B.n160 163.367
R478 B.n165 B.n164 163.367
R479 B.n169 B.n168 163.367
R480 B.n173 B.n172 163.367
R481 B.n177 B.n176 163.367
R482 B.n181 B.n180 163.367
R483 B.n185 B.n184 163.367
R484 B.n190 B.n189 163.367
R485 B.n194 B.n193 163.367
R486 B.n198 B.n197 163.367
R487 B.n202 B.n201 163.367
R488 B.n206 B.n205 163.367
R489 B.n210 B.n209 163.367
R490 B.n214 B.n213 163.367
R491 B.n218 B.n217 163.367
R492 B.n222 B.n221 163.367
R493 B.n226 B.n225 163.367
R494 B.n230 B.n229 163.367
R495 B.n234 B.n233 163.367
R496 B.n238 B.n237 163.367
R497 B.n242 B.n241 163.367
R498 B.n246 B.n245 163.367
R499 B.n250 B.n249 163.367
R500 B.n254 B.n253 163.367
R501 B.n258 B.n257 163.367
R502 B.n262 B.n261 163.367
R503 B.n266 B.n265 163.367
R504 B.n270 B.n269 163.367
R505 B.n274 B.n273 163.367
R506 B.n278 B.n277 163.367
R507 B.n282 B.n281 163.367
R508 B.n286 B.n285 163.367
R509 B.n290 B.n289 163.367
R510 B.n294 B.n293 163.367
R511 B.n668 B.n87 163.367
R512 B.n594 B.n327 163.367
R513 B.n594 B.n320 163.367
R514 B.n602 B.n320 163.367
R515 B.n602 B.n318 163.367
R516 B.n606 B.n318 163.367
R517 B.n606 B.n313 163.367
R518 B.n614 B.n313 163.367
R519 B.n614 B.n311 163.367
R520 B.n618 B.n311 163.367
R521 B.n618 B.n305 163.367
R522 B.n626 B.n305 163.367
R523 B.n626 B.n303 163.367
R524 B.n631 B.n303 163.367
R525 B.n631 B.n298 163.367
R526 B.n640 B.n298 163.367
R527 B.n641 B.n640 163.367
R528 B.n641 B.n5 163.367
R529 B.n6 B.n5 163.367
R530 B.n7 B.n6 163.367
R531 B.n647 B.n7 163.367
R532 B.n648 B.n647 163.367
R533 B.n648 B.n13 163.367
R534 B.n14 B.n13 163.367
R535 B.n15 B.n14 163.367
R536 B.n653 B.n15 163.367
R537 B.n653 B.n20 163.367
R538 B.n21 B.n20 163.367
R539 B.n22 B.n21 163.367
R540 B.n658 B.n22 163.367
R541 B.n658 B.n27 163.367
R542 B.n28 B.n27 163.367
R543 B.n29 B.n28 163.367
R544 B.n663 B.n29 163.367
R545 B.n663 B.n34 163.367
R546 B.n35 B.n34 163.367
R547 B.n380 B.n379 163.367
R548 B.n581 B.n379 163.367
R549 B.n579 B.n578 163.367
R550 B.n575 B.n574 163.367
R551 B.n571 B.n570 163.367
R552 B.n567 B.n566 163.367
R553 B.n563 B.n562 163.367
R554 B.n559 B.n558 163.367
R555 B.n555 B.n554 163.367
R556 B.n551 B.n550 163.367
R557 B.n547 B.n546 163.367
R558 B.n543 B.n542 163.367
R559 B.n539 B.n538 163.367
R560 B.n535 B.n534 163.367
R561 B.n531 B.n530 163.367
R562 B.n527 B.n526 163.367
R563 B.n523 B.n522 163.367
R564 B.n519 B.n518 163.367
R565 B.n515 B.n514 163.367
R566 B.n511 B.n510 163.367
R567 B.n507 B.n506 163.367
R568 B.n503 B.n502 163.367
R569 B.n499 B.n498 163.367
R570 B.n495 B.n494 163.367
R571 B.n491 B.n490 163.367
R572 B.n487 B.n486 163.367
R573 B.n483 B.n482 163.367
R574 B.n479 B.n478 163.367
R575 B.n474 B.n473 163.367
R576 B.n470 B.n469 163.367
R577 B.n466 B.n465 163.367
R578 B.n462 B.n461 163.367
R579 B.n458 B.n457 163.367
R580 B.n454 B.n453 163.367
R581 B.n450 B.n449 163.367
R582 B.n446 B.n445 163.367
R583 B.n442 B.n441 163.367
R584 B.n438 B.n437 163.367
R585 B.n434 B.n433 163.367
R586 B.n430 B.n429 163.367
R587 B.n426 B.n425 163.367
R588 B.n422 B.n421 163.367
R589 B.n418 B.n417 163.367
R590 B.n414 B.n413 163.367
R591 B.n410 B.n409 163.367
R592 B.n406 B.n405 163.367
R593 B.n402 B.n401 163.367
R594 B.n398 B.n397 163.367
R595 B.n394 B.n393 163.367
R596 B.n390 B.n389 163.367
R597 B.n386 B.n329 163.367
R598 B.n596 B.n325 163.367
R599 B.n596 B.n323 163.367
R600 B.n600 B.n323 163.367
R601 B.n600 B.n317 163.367
R602 B.n608 B.n317 163.367
R603 B.n608 B.n315 163.367
R604 B.n612 B.n315 163.367
R605 B.n612 B.n309 163.367
R606 B.n620 B.n309 163.367
R607 B.n620 B.n307 163.367
R608 B.n624 B.n307 163.367
R609 B.n624 B.n301 163.367
R610 B.n634 B.n301 163.367
R611 B.n634 B.n299 163.367
R612 B.n638 B.n299 163.367
R613 B.n638 B.n3 163.367
R614 B.n705 B.n3 163.367
R615 B.n701 B.n2 163.367
R616 B.n701 B.n700 163.367
R617 B.n700 B.n9 163.367
R618 B.n696 B.n9 163.367
R619 B.n696 B.n11 163.367
R620 B.n692 B.n11 163.367
R621 B.n692 B.n17 163.367
R622 B.n688 B.n17 163.367
R623 B.n688 B.n19 163.367
R624 B.n684 B.n19 163.367
R625 B.n684 B.n24 163.367
R626 B.n680 B.n24 163.367
R627 B.n680 B.n26 163.367
R628 B.n676 B.n26 163.367
R629 B.n676 B.n31 163.367
R630 B.n672 B.n31 163.367
R631 B.n672 B.n33 163.367
R632 B.n88 B.t6 90.8583
R633 B.n384 B.t14 90.8583
R634 B.n91 B.t16 90.8405
R635 B.n381 B.t11 90.8405
R636 B.n588 B.n326 77.0208
R637 B.n670 B.n669 77.0208
R638 B.n93 B.n36 71.676
R639 B.n97 B.n37 71.676
R640 B.n101 B.n38 71.676
R641 B.n105 B.n39 71.676
R642 B.n109 B.n40 71.676
R643 B.n113 B.n41 71.676
R644 B.n117 B.n42 71.676
R645 B.n121 B.n43 71.676
R646 B.n125 B.n44 71.676
R647 B.n129 B.n45 71.676
R648 B.n133 B.n46 71.676
R649 B.n137 B.n47 71.676
R650 B.n141 B.n48 71.676
R651 B.n145 B.n49 71.676
R652 B.n149 B.n50 71.676
R653 B.n153 B.n51 71.676
R654 B.n157 B.n52 71.676
R655 B.n161 B.n53 71.676
R656 B.n165 B.n54 71.676
R657 B.n169 B.n55 71.676
R658 B.n173 B.n56 71.676
R659 B.n177 B.n57 71.676
R660 B.n181 B.n58 71.676
R661 B.n185 B.n59 71.676
R662 B.n190 B.n60 71.676
R663 B.n194 B.n61 71.676
R664 B.n198 B.n62 71.676
R665 B.n202 B.n63 71.676
R666 B.n206 B.n64 71.676
R667 B.n210 B.n65 71.676
R668 B.n214 B.n66 71.676
R669 B.n218 B.n67 71.676
R670 B.n222 B.n68 71.676
R671 B.n226 B.n69 71.676
R672 B.n230 B.n70 71.676
R673 B.n234 B.n71 71.676
R674 B.n238 B.n72 71.676
R675 B.n242 B.n73 71.676
R676 B.n246 B.n74 71.676
R677 B.n250 B.n75 71.676
R678 B.n254 B.n76 71.676
R679 B.n258 B.n77 71.676
R680 B.n262 B.n78 71.676
R681 B.n266 B.n79 71.676
R682 B.n270 B.n80 71.676
R683 B.n274 B.n81 71.676
R684 B.n278 B.n82 71.676
R685 B.n282 B.n83 71.676
R686 B.n286 B.n84 71.676
R687 B.n290 B.n85 71.676
R688 B.n294 B.n86 71.676
R689 B.n87 B.n86 71.676
R690 B.n293 B.n85 71.676
R691 B.n289 B.n84 71.676
R692 B.n285 B.n83 71.676
R693 B.n281 B.n82 71.676
R694 B.n277 B.n81 71.676
R695 B.n273 B.n80 71.676
R696 B.n269 B.n79 71.676
R697 B.n265 B.n78 71.676
R698 B.n261 B.n77 71.676
R699 B.n257 B.n76 71.676
R700 B.n253 B.n75 71.676
R701 B.n249 B.n74 71.676
R702 B.n245 B.n73 71.676
R703 B.n241 B.n72 71.676
R704 B.n237 B.n71 71.676
R705 B.n233 B.n70 71.676
R706 B.n229 B.n69 71.676
R707 B.n225 B.n68 71.676
R708 B.n221 B.n67 71.676
R709 B.n217 B.n66 71.676
R710 B.n213 B.n65 71.676
R711 B.n209 B.n64 71.676
R712 B.n205 B.n63 71.676
R713 B.n201 B.n62 71.676
R714 B.n197 B.n61 71.676
R715 B.n193 B.n60 71.676
R716 B.n189 B.n59 71.676
R717 B.n184 B.n58 71.676
R718 B.n180 B.n57 71.676
R719 B.n176 B.n56 71.676
R720 B.n172 B.n55 71.676
R721 B.n168 B.n54 71.676
R722 B.n164 B.n53 71.676
R723 B.n160 B.n52 71.676
R724 B.n156 B.n51 71.676
R725 B.n152 B.n50 71.676
R726 B.n148 B.n49 71.676
R727 B.n144 B.n48 71.676
R728 B.n140 B.n47 71.676
R729 B.n136 B.n46 71.676
R730 B.n132 B.n45 71.676
R731 B.n128 B.n44 71.676
R732 B.n124 B.n43 71.676
R733 B.n120 B.n42 71.676
R734 B.n116 B.n41 71.676
R735 B.n112 B.n40 71.676
R736 B.n108 B.n39 71.676
R737 B.n104 B.n38 71.676
R738 B.n100 B.n37 71.676
R739 B.n96 B.n36 71.676
R740 B.n587 B.n586 71.676
R741 B.n581 B.n330 71.676
R742 B.n578 B.n331 71.676
R743 B.n574 B.n332 71.676
R744 B.n570 B.n333 71.676
R745 B.n566 B.n334 71.676
R746 B.n562 B.n335 71.676
R747 B.n558 B.n336 71.676
R748 B.n554 B.n337 71.676
R749 B.n550 B.n338 71.676
R750 B.n546 B.n339 71.676
R751 B.n542 B.n340 71.676
R752 B.n538 B.n341 71.676
R753 B.n534 B.n342 71.676
R754 B.n530 B.n343 71.676
R755 B.n526 B.n344 71.676
R756 B.n522 B.n345 71.676
R757 B.n518 B.n346 71.676
R758 B.n514 B.n347 71.676
R759 B.n510 B.n348 71.676
R760 B.n506 B.n349 71.676
R761 B.n502 B.n350 71.676
R762 B.n498 B.n351 71.676
R763 B.n494 B.n352 71.676
R764 B.n490 B.n353 71.676
R765 B.n486 B.n354 71.676
R766 B.n482 B.n355 71.676
R767 B.n478 B.n356 71.676
R768 B.n473 B.n357 71.676
R769 B.n469 B.n358 71.676
R770 B.n465 B.n359 71.676
R771 B.n461 B.n360 71.676
R772 B.n457 B.n361 71.676
R773 B.n453 B.n362 71.676
R774 B.n449 B.n363 71.676
R775 B.n445 B.n364 71.676
R776 B.n441 B.n365 71.676
R777 B.n437 B.n366 71.676
R778 B.n433 B.n367 71.676
R779 B.n429 B.n368 71.676
R780 B.n425 B.n369 71.676
R781 B.n421 B.n370 71.676
R782 B.n417 B.n371 71.676
R783 B.n413 B.n372 71.676
R784 B.n409 B.n373 71.676
R785 B.n405 B.n374 71.676
R786 B.n401 B.n375 71.676
R787 B.n397 B.n376 71.676
R788 B.n393 B.n377 71.676
R789 B.n389 B.n378 71.676
R790 B.n589 B.n329 71.676
R791 B.n587 B.n380 71.676
R792 B.n579 B.n330 71.676
R793 B.n575 B.n331 71.676
R794 B.n571 B.n332 71.676
R795 B.n567 B.n333 71.676
R796 B.n563 B.n334 71.676
R797 B.n559 B.n335 71.676
R798 B.n555 B.n336 71.676
R799 B.n551 B.n337 71.676
R800 B.n547 B.n338 71.676
R801 B.n543 B.n339 71.676
R802 B.n539 B.n340 71.676
R803 B.n535 B.n341 71.676
R804 B.n531 B.n342 71.676
R805 B.n527 B.n343 71.676
R806 B.n523 B.n344 71.676
R807 B.n519 B.n345 71.676
R808 B.n515 B.n346 71.676
R809 B.n511 B.n347 71.676
R810 B.n507 B.n348 71.676
R811 B.n503 B.n349 71.676
R812 B.n499 B.n350 71.676
R813 B.n495 B.n351 71.676
R814 B.n491 B.n352 71.676
R815 B.n487 B.n353 71.676
R816 B.n483 B.n354 71.676
R817 B.n479 B.n355 71.676
R818 B.n474 B.n356 71.676
R819 B.n470 B.n357 71.676
R820 B.n466 B.n358 71.676
R821 B.n462 B.n359 71.676
R822 B.n458 B.n360 71.676
R823 B.n454 B.n361 71.676
R824 B.n450 B.n362 71.676
R825 B.n446 B.n363 71.676
R826 B.n442 B.n364 71.676
R827 B.n438 B.n365 71.676
R828 B.n434 B.n366 71.676
R829 B.n430 B.n367 71.676
R830 B.n426 B.n368 71.676
R831 B.n422 B.n369 71.676
R832 B.n418 B.n370 71.676
R833 B.n414 B.n371 71.676
R834 B.n410 B.n372 71.676
R835 B.n406 B.n373 71.676
R836 B.n402 B.n374 71.676
R837 B.n398 B.n375 71.676
R838 B.n394 B.n376 71.676
R839 B.n390 B.n377 71.676
R840 B.n386 B.n378 71.676
R841 B.n590 B.n589 71.676
R842 B.n706 B.n705 71.676
R843 B.n706 B.n2 71.676
R844 B.n89 B.t7 69.9128
R845 B.n385 B.t13 69.9128
R846 B.n92 B.t17 69.8951
R847 B.n382 B.t10 69.8951
R848 B.n187 B.n92 59.5399
R849 B.n90 B.n89 59.5399
R850 B.n476 B.n385 59.5399
R851 B.n383 B.n382 59.5399
R852 B.n595 B.n326 39.3793
R853 B.n595 B.n321 39.3793
R854 B.n601 B.n321 39.3793
R855 B.n601 B.n322 39.3793
R856 B.n607 B.n314 39.3793
R857 B.n613 B.n314 39.3793
R858 B.n613 B.n310 39.3793
R859 B.n619 B.n310 39.3793
R860 B.n619 B.n306 39.3793
R861 B.n625 B.n306 39.3793
R862 B.n633 B.n302 39.3793
R863 B.n633 B.n632 39.3793
R864 B.n639 B.n4 39.3793
R865 B.n704 B.n4 39.3793
R866 B.n704 B.n703 39.3793
R867 B.n703 B.n702 39.3793
R868 B.n702 B.n8 39.3793
R869 B.n695 B.n12 39.3793
R870 B.n695 B.n694 39.3793
R871 B.n693 B.n16 39.3793
R872 B.n687 B.n16 39.3793
R873 B.n687 B.n686 39.3793
R874 B.n686 B.n685 39.3793
R875 B.n685 B.n23 39.3793
R876 B.n679 B.n23 39.3793
R877 B.n678 B.n677 39.3793
R878 B.n677 B.n30 39.3793
R879 B.n671 B.n30 39.3793
R880 B.n671 B.n670 39.3793
R881 B.t0 B.n302 34.1674
R882 B.n694 B.t2 34.1674
R883 B.n585 B.n324 33.5615
R884 B.n592 B.n591 33.5615
R885 B.n667 B.n666 33.5615
R886 B.n94 B.n32 33.5615
R887 B.n322 B.t9 29.5346
R888 B.t5 B.n678 29.5346
R889 B.n639 B.t1 27.2182
R890 B.t3 B.n8 27.2182
R891 B.n92 B.n91 20.946
R892 B.n89 B.n88 20.946
R893 B.n385 B.n384 20.946
R894 B.n382 B.n381 20.946
R895 B B.n707 18.0485
R896 B.n632 B.t1 12.1616
R897 B.n12 B.t3 12.1616
R898 B.n597 B.n324 10.6151
R899 B.n598 B.n597 10.6151
R900 B.n599 B.n598 10.6151
R901 B.n599 B.n316 10.6151
R902 B.n609 B.n316 10.6151
R903 B.n610 B.n609 10.6151
R904 B.n611 B.n610 10.6151
R905 B.n611 B.n308 10.6151
R906 B.n621 B.n308 10.6151
R907 B.n622 B.n621 10.6151
R908 B.n623 B.n622 10.6151
R909 B.n623 B.n300 10.6151
R910 B.n635 B.n300 10.6151
R911 B.n636 B.n635 10.6151
R912 B.n637 B.n636 10.6151
R913 B.n637 B.n0 10.6151
R914 B.n585 B.n584 10.6151
R915 B.n584 B.n583 10.6151
R916 B.n583 B.n582 10.6151
R917 B.n582 B.n580 10.6151
R918 B.n580 B.n577 10.6151
R919 B.n577 B.n576 10.6151
R920 B.n576 B.n573 10.6151
R921 B.n573 B.n572 10.6151
R922 B.n572 B.n569 10.6151
R923 B.n569 B.n568 10.6151
R924 B.n568 B.n565 10.6151
R925 B.n565 B.n564 10.6151
R926 B.n564 B.n561 10.6151
R927 B.n561 B.n560 10.6151
R928 B.n560 B.n557 10.6151
R929 B.n557 B.n556 10.6151
R930 B.n556 B.n553 10.6151
R931 B.n553 B.n552 10.6151
R932 B.n552 B.n549 10.6151
R933 B.n549 B.n548 10.6151
R934 B.n548 B.n545 10.6151
R935 B.n545 B.n544 10.6151
R936 B.n544 B.n541 10.6151
R937 B.n541 B.n540 10.6151
R938 B.n540 B.n537 10.6151
R939 B.n537 B.n536 10.6151
R940 B.n536 B.n533 10.6151
R941 B.n533 B.n532 10.6151
R942 B.n532 B.n529 10.6151
R943 B.n529 B.n528 10.6151
R944 B.n528 B.n525 10.6151
R945 B.n525 B.n524 10.6151
R946 B.n524 B.n521 10.6151
R947 B.n521 B.n520 10.6151
R948 B.n520 B.n517 10.6151
R949 B.n517 B.n516 10.6151
R950 B.n516 B.n513 10.6151
R951 B.n513 B.n512 10.6151
R952 B.n512 B.n509 10.6151
R953 B.n509 B.n508 10.6151
R954 B.n508 B.n505 10.6151
R955 B.n505 B.n504 10.6151
R956 B.n504 B.n501 10.6151
R957 B.n501 B.n500 10.6151
R958 B.n500 B.n497 10.6151
R959 B.n497 B.n496 10.6151
R960 B.n493 B.n492 10.6151
R961 B.n492 B.n489 10.6151
R962 B.n489 B.n488 10.6151
R963 B.n488 B.n485 10.6151
R964 B.n485 B.n484 10.6151
R965 B.n484 B.n481 10.6151
R966 B.n481 B.n480 10.6151
R967 B.n480 B.n477 10.6151
R968 B.n475 B.n472 10.6151
R969 B.n472 B.n471 10.6151
R970 B.n471 B.n468 10.6151
R971 B.n468 B.n467 10.6151
R972 B.n467 B.n464 10.6151
R973 B.n464 B.n463 10.6151
R974 B.n463 B.n460 10.6151
R975 B.n460 B.n459 10.6151
R976 B.n459 B.n456 10.6151
R977 B.n456 B.n455 10.6151
R978 B.n455 B.n452 10.6151
R979 B.n452 B.n451 10.6151
R980 B.n451 B.n448 10.6151
R981 B.n448 B.n447 10.6151
R982 B.n447 B.n444 10.6151
R983 B.n444 B.n443 10.6151
R984 B.n443 B.n440 10.6151
R985 B.n440 B.n439 10.6151
R986 B.n439 B.n436 10.6151
R987 B.n436 B.n435 10.6151
R988 B.n435 B.n432 10.6151
R989 B.n432 B.n431 10.6151
R990 B.n431 B.n428 10.6151
R991 B.n428 B.n427 10.6151
R992 B.n427 B.n424 10.6151
R993 B.n424 B.n423 10.6151
R994 B.n423 B.n420 10.6151
R995 B.n420 B.n419 10.6151
R996 B.n419 B.n416 10.6151
R997 B.n416 B.n415 10.6151
R998 B.n415 B.n412 10.6151
R999 B.n412 B.n411 10.6151
R1000 B.n411 B.n408 10.6151
R1001 B.n408 B.n407 10.6151
R1002 B.n407 B.n404 10.6151
R1003 B.n404 B.n403 10.6151
R1004 B.n403 B.n400 10.6151
R1005 B.n400 B.n399 10.6151
R1006 B.n399 B.n396 10.6151
R1007 B.n396 B.n395 10.6151
R1008 B.n395 B.n392 10.6151
R1009 B.n392 B.n391 10.6151
R1010 B.n391 B.n388 10.6151
R1011 B.n388 B.n387 10.6151
R1012 B.n387 B.n328 10.6151
R1013 B.n591 B.n328 10.6151
R1014 B.n593 B.n592 10.6151
R1015 B.n593 B.n319 10.6151
R1016 B.n603 B.n319 10.6151
R1017 B.n604 B.n603 10.6151
R1018 B.n605 B.n604 10.6151
R1019 B.n605 B.n312 10.6151
R1020 B.n615 B.n312 10.6151
R1021 B.n616 B.n615 10.6151
R1022 B.n617 B.n616 10.6151
R1023 B.n617 B.n304 10.6151
R1024 B.n627 B.n304 10.6151
R1025 B.n628 B.n627 10.6151
R1026 B.n630 B.n628 10.6151
R1027 B.n630 B.n629 10.6151
R1028 B.n629 B.n297 10.6151
R1029 B.n642 B.n297 10.6151
R1030 B.n643 B.n642 10.6151
R1031 B.n644 B.n643 10.6151
R1032 B.n645 B.n644 10.6151
R1033 B.n646 B.n645 10.6151
R1034 B.n649 B.n646 10.6151
R1035 B.n650 B.n649 10.6151
R1036 B.n651 B.n650 10.6151
R1037 B.n652 B.n651 10.6151
R1038 B.n654 B.n652 10.6151
R1039 B.n655 B.n654 10.6151
R1040 B.n656 B.n655 10.6151
R1041 B.n657 B.n656 10.6151
R1042 B.n659 B.n657 10.6151
R1043 B.n660 B.n659 10.6151
R1044 B.n661 B.n660 10.6151
R1045 B.n662 B.n661 10.6151
R1046 B.n664 B.n662 10.6151
R1047 B.n665 B.n664 10.6151
R1048 B.n666 B.n665 10.6151
R1049 B.n699 B.n1 10.6151
R1050 B.n699 B.n698 10.6151
R1051 B.n698 B.n697 10.6151
R1052 B.n697 B.n10 10.6151
R1053 B.n691 B.n10 10.6151
R1054 B.n691 B.n690 10.6151
R1055 B.n690 B.n689 10.6151
R1056 B.n689 B.n18 10.6151
R1057 B.n683 B.n18 10.6151
R1058 B.n683 B.n682 10.6151
R1059 B.n682 B.n681 10.6151
R1060 B.n681 B.n25 10.6151
R1061 B.n675 B.n25 10.6151
R1062 B.n675 B.n674 10.6151
R1063 B.n674 B.n673 10.6151
R1064 B.n673 B.n32 10.6151
R1065 B.n95 B.n94 10.6151
R1066 B.n98 B.n95 10.6151
R1067 B.n99 B.n98 10.6151
R1068 B.n102 B.n99 10.6151
R1069 B.n103 B.n102 10.6151
R1070 B.n106 B.n103 10.6151
R1071 B.n107 B.n106 10.6151
R1072 B.n110 B.n107 10.6151
R1073 B.n111 B.n110 10.6151
R1074 B.n114 B.n111 10.6151
R1075 B.n115 B.n114 10.6151
R1076 B.n118 B.n115 10.6151
R1077 B.n119 B.n118 10.6151
R1078 B.n122 B.n119 10.6151
R1079 B.n123 B.n122 10.6151
R1080 B.n126 B.n123 10.6151
R1081 B.n127 B.n126 10.6151
R1082 B.n130 B.n127 10.6151
R1083 B.n131 B.n130 10.6151
R1084 B.n134 B.n131 10.6151
R1085 B.n135 B.n134 10.6151
R1086 B.n138 B.n135 10.6151
R1087 B.n139 B.n138 10.6151
R1088 B.n142 B.n139 10.6151
R1089 B.n143 B.n142 10.6151
R1090 B.n146 B.n143 10.6151
R1091 B.n147 B.n146 10.6151
R1092 B.n150 B.n147 10.6151
R1093 B.n151 B.n150 10.6151
R1094 B.n154 B.n151 10.6151
R1095 B.n155 B.n154 10.6151
R1096 B.n158 B.n155 10.6151
R1097 B.n159 B.n158 10.6151
R1098 B.n162 B.n159 10.6151
R1099 B.n163 B.n162 10.6151
R1100 B.n166 B.n163 10.6151
R1101 B.n167 B.n166 10.6151
R1102 B.n170 B.n167 10.6151
R1103 B.n171 B.n170 10.6151
R1104 B.n174 B.n171 10.6151
R1105 B.n175 B.n174 10.6151
R1106 B.n178 B.n175 10.6151
R1107 B.n179 B.n178 10.6151
R1108 B.n182 B.n179 10.6151
R1109 B.n183 B.n182 10.6151
R1110 B.n186 B.n183 10.6151
R1111 B.n191 B.n188 10.6151
R1112 B.n192 B.n191 10.6151
R1113 B.n195 B.n192 10.6151
R1114 B.n196 B.n195 10.6151
R1115 B.n199 B.n196 10.6151
R1116 B.n200 B.n199 10.6151
R1117 B.n203 B.n200 10.6151
R1118 B.n204 B.n203 10.6151
R1119 B.n208 B.n207 10.6151
R1120 B.n211 B.n208 10.6151
R1121 B.n212 B.n211 10.6151
R1122 B.n215 B.n212 10.6151
R1123 B.n216 B.n215 10.6151
R1124 B.n219 B.n216 10.6151
R1125 B.n220 B.n219 10.6151
R1126 B.n223 B.n220 10.6151
R1127 B.n224 B.n223 10.6151
R1128 B.n227 B.n224 10.6151
R1129 B.n228 B.n227 10.6151
R1130 B.n231 B.n228 10.6151
R1131 B.n232 B.n231 10.6151
R1132 B.n235 B.n232 10.6151
R1133 B.n236 B.n235 10.6151
R1134 B.n239 B.n236 10.6151
R1135 B.n240 B.n239 10.6151
R1136 B.n243 B.n240 10.6151
R1137 B.n244 B.n243 10.6151
R1138 B.n247 B.n244 10.6151
R1139 B.n248 B.n247 10.6151
R1140 B.n251 B.n248 10.6151
R1141 B.n252 B.n251 10.6151
R1142 B.n255 B.n252 10.6151
R1143 B.n256 B.n255 10.6151
R1144 B.n259 B.n256 10.6151
R1145 B.n260 B.n259 10.6151
R1146 B.n263 B.n260 10.6151
R1147 B.n264 B.n263 10.6151
R1148 B.n267 B.n264 10.6151
R1149 B.n268 B.n267 10.6151
R1150 B.n271 B.n268 10.6151
R1151 B.n272 B.n271 10.6151
R1152 B.n275 B.n272 10.6151
R1153 B.n276 B.n275 10.6151
R1154 B.n279 B.n276 10.6151
R1155 B.n280 B.n279 10.6151
R1156 B.n283 B.n280 10.6151
R1157 B.n284 B.n283 10.6151
R1158 B.n287 B.n284 10.6151
R1159 B.n288 B.n287 10.6151
R1160 B.n291 B.n288 10.6151
R1161 B.n292 B.n291 10.6151
R1162 B.n295 B.n292 10.6151
R1163 B.n296 B.n295 10.6151
R1164 B.n667 B.n296 10.6151
R1165 B.n607 B.t9 9.8452
R1166 B.n679 B.t5 9.8452
R1167 B.n707 B.n0 8.11757
R1168 B.n707 B.n1 8.11757
R1169 B.n493 B.n383 6.5566
R1170 B.n477 B.n476 6.5566
R1171 B.n188 B.n187 6.5566
R1172 B.n204 B.n90 6.5566
R1173 B.n625 B.t0 5.2124
R1174 B.t2 B.n693 5.2124
R1175 B.n496 B.n383 4.05904
R1176 B.n476 B.n475 4.05904
R1177 B.n187 B.n186 4.05904
R1178 B.n207 B.n90 4.05904
R1179 VN.n0 VN.t0 514.886
R1180 VN.n1 VN.t2 514.886
R1181 VN.n0 VN.t1 514.837
R1182 VN.n1 VN.t3 514.837
R1183 VN VN.n1 86.9443
R1184 VN VN.n0 44.7132
R1185 VDD2.n2 VDD2.n0 102.505
R1186 VDD2.n2 VDD2.n1 64.17
R1187 VDD2.n1 VDD2.t3 1.44365
R1188 VDD2.n1 VDD2.t2 1.44365
R1189 VDD2.n0 VDD2.t0 1.44365
R1190 VDD2.n0 VDD2.t1 1.44365
R1191 VDD2 VDD2.n2 0.0586897
R1192 VTAIL.n5 VTAIL.t3 48.9345
R1193 VTAIL.n4 VTAIL.t5 48.9345
R1194 VTAIL.n3 VTAIL.t4 48.9345
R1195 VTAIL.n7 VTAIL.t6 48.9343
R1196 VTAIL.n0 VTAIL.t7 48.9343
R1197 VTAIL.n1 VTAIL.t1 48.9343
R1198 VTAIL.n2 VTAIL.t0 48.9343
R1199 VTAIL.n6 VTAIL.t2 48.9343
R1200 VTAIL.n7 VTAIL.n6 25.1255
R1201 VTAIL.n3 VTAIL.n2 25.1255
R1202 VTAIL.n4 VTAIL.n3 0.931535
R1203 VTAIL.n6 VTAIL.n5 0.931535
R1204 VTAIL.n2 VTAIL.n1 0.931535
R1205 VTAIL VTAIL.n0 0.524207
R1206 VTAIL.n5 VTAIL.n4 0.470328
R1207 VTAIL.n1 VTAIL.n0 0.470328
R1208 VTAIL VTAIL.n7 0.407828
R1209 VP.n1 VP.t2 514.886
R1210 VP.n1 VP.t1 514.837
R1211 VP.n3 VP.t3 493.889
R1212 VP.n5 VP.t0 493.889
R1213 VP.n6 VP.n5 161.3
R1214 VP.n4 VP.n0 161.3
R1215 VP.n3 VP.n2 161.3
R1216 VP.n2 VP.n1 86.5636
R1217 VP.n4 VP.n3 24.1005
R1218 VP.n5 VP.n4 24.1005
R1219 VP.n2 VP.n0 0.189894
R1220 VP.n6 VP.n0 0.189894
R1221 VP VP.n6 0.0516364
R1222 VDD1 VDD1.n1 103.031
R1223 VDD1 VDD1.n0 64.2282
R1224 VDD1.n0 VDD1.t1 1.44365
R1225 VDD1.n0 VDD1.t2 1.44365
R1226 VDD1.n1 VDD1.t0 1.44365
R1227 VDD1.n1 VDD1.t3 1.44365
C0 VDD1 VP 3.81534f
C1 VN VP 5.17943f
C2 VP VDD2 0.276059f
C3 VDD1 VN 0.146801f
C4 VDD1 VDD2 0.577924f
C5 VN VDD2 3.68635f
C6 VP VTAIL 3.24822f
C7 VDD1 VTAIL 7.36231f
C8 VN VTAIL 3.23412f
C9 VTAIL VDD2 7.40411f
C10 VDD2 B 2.862212f
C11 VDD1 B 6.76003f
C12 VTAIL B 9.816226f
C13 VN B 8.444321f
C14 VP B 5.118975f
C15 VDD1.t1 B 0.304065f
C16 VDD1.t2 B 0.304065f
C17 VDD1.n0 B 2.74053f
C18 VDD1.t0 B 0.304065f
C19 VDD1.t3 B 0.304065f
C20 VDD1.n1 B 3.41554f
C21 VP.n0 B 0.048694f
C22 VP.t1 B 1.44901f
C23 VP.t2 B 1.44907f
C24 VP.n1 B 2.09291f
C25 VP.n2 B 3.132f
C26 VP.t3 B 1.42637f
C27 VP.n3 B 0.552967f
C28 VP.n4 B 0.01105f
C29 VP.t0 B 1.42637f
C30 VP.n5 B 0.552967f
C31 VP.n6 B 0.037736f
C32 VTAIL.t7 B 1.94599f
C33 VTAIL.n0 B 0.255929f
C34 VTAIL.t1 B 1.94599f
C35 VTAIL.n1 B 0.277006f
C36 VTAIL.t0 B 1.94599f
C37 VTAIL.n2 B 1.13101f
C38 VTAIL.t4 B 1.94599f
C39 VTAIL.n3 B 1.13101f
C40 VTAIL.t5 B 1.94599f
C41 VTAIL.n4 B 0.277004f
C42 VTAIL.t3 B 1.94599f
C43 VTAIL.n5 B 0.277004f
C44 VTAIL.t2 B 1.94599f
C45 VTAIL.n6 B 1.13101f
C46 VTAIL.t6 B 1.94599f
C47 VTAIL.n7 B 1.10392f
C48 VDD2.t0 B 0.304163f
C49 VDD2.t1 B 0.304163f
C50 VDD2.n0 B 3.38975f
C51 VDD2.t3 B 0.304163f
C52 VDD2.t2 B 0.304163f
C53 VDD2.n1 B 2.74112f
C54 VDD2.n2 B 3.66228f
C55 VN.t0 B 1.42917f
C56 VN.t1 B 1.42911f
C57 VN.n0 B 1.05743f
C58 VN.t2 B 1.42917f
C59 VN.t3 B 1.42911f
C60 VN.n1 B 2.08421f
.ends

