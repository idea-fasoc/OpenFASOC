* NGSPICE file created from diff_pair_sample_0114.ext - technology: sky130A

.subckt diff_pair_sample_0114 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3666_n1348# sky130_fd_pr__pfet_01v8 ad=0.741 pd=4.58 as=0 ps=0 w=1.9 l=3.04
X1 VDD1.t5 VP.t0 VTAIL.t7 w_n3666_n1348# sky130_fd_pr__pfet_01v8 ad=0.3135 pd=2.23 as=0.741 ps=4.58 w=1.9 l=3.04
X2 B.t8 B.t6 B.t7 w_n3666_n1348# sky130_fd_pr__pfet_01v8 ad=0.741 pd=4.58 as=0 ps=0 w=1.9 l=3.04
X3 VDD1.t4 VP.t1 VTAIL.t6 w_n3666_n1348# sky130_fd_pr__pfet_01v8 ad=0.741 pd=4.58 as=0.3135 ps=2.23 w=1.9 l=3.04
X4 VTAIL.t10 VP.t2 VDD1.t3 w_n3666_n1348# sky130_fd_pr__pfet_01v8 ad=0.3135 pd=2.23 as=0.3135 ps=2.23 w=1.9 l=3.04
X5 VDD2.t5 VN.t0 VTAIL.t3 w_n3666_n1348# sky130_fd_pr__pfet_01v8 ad=0.3135 pd=2.23 as=0.741 ps=4.58 w=1.9 l=3.04
X6 VDD1.t2 VP.t3 VTAIL.t11 w_n3666_n1348# sky130_fd_pr__pfet_01v8 ad=0.3135 pd=2.23 as=0.741 ps=4.58 w=1.9 l=3.04
X7 VDD2.t4 VN.t1 VTAIL.t1 w_n3666_n1348# sky130_fd_pr__pfet_01v8 ad=0.3135 pd=2.23 as=0.741 ps=4.58 w=1.9 l=3.04
X8 VTAIL.t4 VN.t2 VDD2.t3 w_n3666_n1348# sky130_fd_pr__pfet_01v8 ad=0.3135 pd=2.23 as=0.3135 ps=2.23 w=1.9 l=3.04
X9 VTAIL.t9 VP.t4 VDD1.t1 w_n3666_n1348# sky130_fd_pr__pfet_01v8 ad=0.3135 pd=2.23 as=0.3135 ps=2.23 w=1.9 l=3.04
X10 B.t5 B.t3 B.t4 w_n3666_n1348# sky130_fd_pr__pfet_01v8 ad=0.741 pd=4.58 as=0 ps=0 w=1.9 l=3.04
X11 VTAIL.t5 VN.t3 VDD2.t2 w_n3666_n1348# sky130_fd_pr__pfet_01v8 ad=0.3135 pd=2.23 as=0.3135 ps=2.23 w=1.9 l=3.04
X12 B.t2 B.t0 B.t1 w_n3666_n1348# sky130_fd_pr__pfet_01v8 ad=0.741 pd=4.58 as=0 ps=0 w=1.9 l=3.04
X13 VDD1.t0 VP.t5 VTAIL.t8 w_n3666_n1348# sky130_fd_pr__pfet_01v8 ad=0.741 pd=4.58 as=0.3135 ps=2.23 w=1.9 l=3.04
X14 VDD2.t1 VN.t4 VTAIL.t2 w_n3666_n1348# sky130_fd_pr__pfet_01v8 ad=0.741 pd=4.58 as=0.3135 ps=2.23 w=1.9 l=3.04
X15 VDD2.t0 VN.t5 VTAIL.t0 w_n3666_n1348# sky130_fd_pr__pfet_01v8 ad=0.741 pd=4.58 as=0.3135 ps=2.23 w=1.9 l=3.04
R0 B.n258 B.n257 585
R1 B.n256 B.n95 585
R2 B.n255 B.n254 585
R3 B.n253 B.n96 585
R4 B.n252 B.n251 585
R5 B.n250 B.n97 585
R6 B.n249 B.n248 585
R7 B.n247 B.n98 585
R8 B.n246 B.n245 585
R9 B.n244 B.n99 585
R10 B.n243 B.n242 585
R11 B.n241 B.n100 585
R12 B.n240 B.n239 585
R13 B.n235 B.n101 585
R14 B.n234 B.n233 585
R15 B.n232 B.n102 585
R16 B.n231 B.n230 585
R17 B.n229 B.n103 585
R18 B.n228 B.n227 585
R19 B.n226 B.n104 585
R20 B.n225 B.n224 585
R21 B.n222 B.n105 585
R22 B.n221 B.n220 585
R23 B.n219 B.n108 585
R24 B.n218 B.n217 585
R25 B.n216 B.n109 585
R26 B.n215 B.n214 585
R27 B.n213 B.n110 585
R28 B.n212 B.n211 585
R29 B.n210 B.n111 585
R30 B.n209 B.n208 585
R31 B.n207 B.n112 585
R32 B.n206 B.n205 585
R33 B.n259 B.n94 585
R34 B.n261 B.n260 585
R35 B.n262 B.n93 585
R36 B.n264 B.n263 585
R37 B.n265 B.n92 585
R38 B.n267 B.n266 585
R39 B.n268 B.n91 585
R40 B.n270 B.n269 585
R41 B.n271 B.n90 585
R42 B.n273 B.n272 585
R43 B.n274 B.n89 585
R44 B.n276 B.n275 585
R45 B.n277 B.n88 585
R46 B.n279 B.n278 585
R47 B.n280 B.n87 585
R48 B.n282 B.n281 585
R49 B.n283 B.n86 585
R50 B.n285 B.n284 585
R51 B.n286 B.n85 585
R52 B.n288 B.n287 585
R53 B.n289 B.n84 585
R54 B.n291 B.n290 585
R55 B.n292 B.n83 585
R56 B.n294 B.n293 585
R57 B.n295 B.n82 585
R58 B.n297 B.n296 585
R59 B.n298 B.n81 585
R60 B.n300 B.n299 585
R61 B.n301 B.n80 585
R62 B.n303 B.n302 585
R63 B.n304 B.n79 585
R64 B.n306 B.n305 585
R65 B.n307 B.n78 585
R66 B.n309 B.n308 585
R67 B.n310 B.n77 585
R68 B.n312 B.n311 585
R69 B.n313 B.n76 585
R70 B.n315 B.n314 585
R71 B.n316 B.n75 585
R72 B.n318 B.n317 585
R73 B.n319 B.n74 585
R74 B.n321 B.n320 585
R75 B.n322 B.n73 585
R76 B.n324 B.n323 585
R77 B.n325 B.n72 585
R78 B.n327 B.n326 585
R79 B.n328 B.n71 585
R80 B.n330 B.n329 585
R81 B.n331 B.n70 585
R82 B.n333 B.n332 585
R83 B.n334 B.n69 585
R84 B.n336 B.n335 585
R85 B.n337 B.n68 585
R86 B.n339 B.n338 585
R87 B.n340 B.n67 585
R88 B.n342 B.n341 585
R89 B.n343 B.n66 585
R90 B.n345 B.n344 585
R91 B.n346 B.n65 585
R92 B.n348 B.n347 585
R93 B.n349 B.n64 585
R94 B.n351 B.n350 585
R95 B.n352 B.n63 585
R96 B.n354 B.n353 585
R97 B.n355 B.n62 585
R98 B.n357 B.n356 585
R99 B.n358 B.n61 585
R100 B.n360 B.n359 585
R101 B.n361 B.n60 585
R102 B.n363 B.n362 585
R103 B.n364 B.n59 585
R104 B.n366 B.n365 585
R105 B.n367 B.n58 585
R106 B.n369 B.n368 585
R107 B.n370 B.n57 585
R108 B.n372 B.n371 585
R109 B.n373 B.n56 585
R110 B.n375 B.n374 585
R111 B.n376 B.n55 585
R112 B.n378 B.n377 585
R113 B.n379 B.n54 585
R114 B.n381 B.n380 585
R115 B.n382 B.n53 585
R116 B.n384 B.n383 585
R117 B.n385 B.n52 585
R118 B.n387 B.n386 585
R119 B.n388 B.n51 585
R120 B.n390 B.n389 585
R121 B.n391 B.n50 585
R122 B.n393 B.n392 585
R123 B.n394 B.n49 585
R124 B.n396 B.n395 585
R125 B.n397 B.n48 585
R126 B.n399 B.n398 585
R127 B.n400 B.n47 585
R128 B.n402 B.n401 585
R129 B.n453 B.n452 585
R130 B.n451 B.n26 585
R131 B.n450 B.n449 585
R132 B.n448 B.n27 585
R133 B.n447 B.n446 585
R134 B.n445 B.n28 585
R135 B.n444 B.n443 585
R136 B.n442 B.n29 585
R137 B.n441 B.n440 585
R138 B.n439 B.n30 585
R139 B.n438 B.n437 585
R140 B.n436 B.n31 585
R141 B.n434 B.n433 585
R142 B.n432 B.n34 585
R143 B.n431 B.n430 585
R144 B.n429 B.n35 585
R145 B.n428 B.n427 585
R146 B.n426 B.n36 585
R147 B.n425 B.n424 585
R148 B.n423 B.n37 585
R149 B.n422 B.n421 585
R150 B.n420 B.n419 585
R151 B.n418 B.n41 585
R152 B.n417 B.n416 585
R153 B.n415 B.n42 585
R154 B.n414 B.n413 585
R155 B.n412 B.n43 585
R156 B.n411 B.n410 585
R157 B.n409 B.n44 585
R158 B.n408 B.n407 585
R159 B.n406 B.n45 585
R160 B.n405 B.n404 585
R161 B.n403 B.n46 585
R162 B.n454 B.n25 585
R163 B.n456 B.n455 585
R164 B.n457 B.n24 585
R165 B.n459 B.n458 585
R166 B.n460 B.n23 585
R167 B.n462 B.n461 585
R168 B.n463 B.n22 585
R169 B.n465 B.n464 585
R170 B.n466 B.n21 585
R171 B.n468 B.n467 585
R172 B.n469 B.n20 585
R173 B.n471 B.n470 585
R174 B.n472 B.n19 585
R175 B.n474 B.n473 585
R176 B.n475 B.n18 585
R177 B.n477 B.n476 585
R178 B.n478 B.n17 585
R179 B.n480 B.n479 585
R180 B.n481 B.n16 585
R181 B.n483 B.n482 585
R182 B.n484 B.n15 585
R183 B.n486 B.n485 585
R184 B.n487 B.n14 585
R185 B.n489 B.n488 585
R186 B.n490 B.n13 585
R187 B.n492 B.n491 585
R188 B.n493 B.n12 585
R189 B.n495 B.n494 585
R190 B.n496 B.n11 585
R191 B.n498 B.n497 585
R192 B.n499 B.n10 585
R193 B.n501 B.n500 585
R194 B.n502 B.n9 585
R195 B.n504 B.n503 585
R196 B.n505 B.n8 585
R197 B.n507 B.n506 585
R198 B.n508 B.n7 585
R199 B.n510 B.n509 585
R200 B.n511 B.n6 585
R201 B.n513 B.n512 585
R202 B.n514 B.n5 585
R203 B.n516 B.n515 585
R204 B.n517 B.n4 585
R205 B.n519 B.n518 585
R206 B.n520 B.n3 585
R207 B.n522 B.n521 585
R208 B.n523 B.n0 585
R209 B.n2 B.n1 585
R210 B.n137 B.n136 585
R211 B.n138 B.n135 585
R212 B.n140 B.n139 585
R213 B.n141 B.n134 585
R214 B.n143 B.n142 585
R215 B.n144 B.n133 585
R216 B.n146 B.n145 585
R217 B.n147 B.n132 585
R218 B.n149 B.n148 585
R219 B.n150 B.n131 585
R220 B.n152 B.n151 585
R221 B.n153 B.n130 585
R222 B.n155 B.n154 585
R223 B.n156 B.n129 585
R224 B.n158 B.n157 585
R225 B.n159 B.n128 585
R226 B.n161 B.n160 585
R227 B.n162 B.n127 585
R228 B.n164 B.n163 585
R229 B.n165 B.n126 585
R230 B.n167 B.n166 585
R231 B.n168 B.n125 585
R232 B.n170 B.n169 585
R233 B.n171 B.n124 585
R234 B.n173 B.n172 585
R235 B.n174 B.n123 585
R236 B.n176 B.n175 585
R237 B.n177 B.n122 585
R238 B.n179 B.n178 585
R239 B.n180 B.n121 585
R240 B.n182 B.n181 585
R241 B.n183 B.n120 585
R242 B.n185 B.n184 585
R243 B.n186 B.n119 585
R244 B.n188 B.n187 585
R245 B.n189 B.n118 585
R246 B.n191 B.n190 585
R247 B.n192 B.n117 585
R248 B.n194 B.n193 585
R249 B.n195 B.n116 585
R250 B.n197 B.n196 585
R251 B.n198 B.n115 585
R252 B.n200 B.n199 585
R253 B.n201 B.n114 585
R254 B.n203 B.n202 585
R255 B.n204 B.n113 585
R256 B.n206 B.n113 574.183
R257 B.n259 B.n258 574.183
R258 B.n403 B.n402 574.183
R259 B.n452 B.n25 574.183
R260 B.n236 B.t1 311.755
R261 B.n38 B.t8 311.755
R262 B.n106 B.t10 311.755
R263 B.n32 B.t5 311.755
R264 B.n525 B.n524 256.663
R265 B.n237 B.t2 246.399
R266 B.n39 B.t7 246.399
R267 B.n107 B.t11 246.399
R268 B.n33 B.t4 246.399
R269 B.n524 B.n523 235.042
R270 B.n524 B.n2 235.042
R271 B.n106 B.t9 223.69
R272 B.n236 B.t0 223.69
R273 B.n38 B.t6 223.69
R274 B.n32 B.t3 223.69
R275 B.n207 B.n206 163.367
R276 B.n208 B.n207 163.367
R277 B.n208 B.n111 163.367
R278 B.n212 B.n111 163.367
R279 B.n213 B.n212 163.367
R280 B.n214 B.n213 163.367
R281 B.n214 B.n109 163.367
R282 B.n218 B.n109 163.367
R283 B.n219 B.n218 163.367
R284 B.n220 B.n219 163.367
R285 B.n220 B.n105 163.367
R286 B.n225 B.n105 163.367
R287 B.n226 B.n225 163.367
R288 B.n227 B.n226 163.367
R289 B.n227 B.n103 163.367
R290 B.n231 B.n103 163.367
R291 B.n232 B.n231 163.367
R292 B.n233 B.n232 163.367
R293 B.n233 B.n101 163.367
R294 B.n240 B.n101 163.367
R295 B.n241 B.n240 163.367
R296 B.n242 B.n241 163.367
R297 B.n242 B.n99 163.367
R298 B.n246 B.n99 163.367
R299 B.n247 B.n246 163.367
R300 B.n248 B.n247 163.367
R301 B.n248 B.n97 163.367
R302 B.n252 B.n97 163.367
R303 B.n253 B.n252 163.367
R304 B.n254 B.n253 163.367
R305 B.n254 B.n95 163.367
R306 B.n258 B.n95 163.367
R307 B.n402 B.n47 163.367
R308 B.n398 B.n47 163.367
R309 B.n398 B.n397 163.367
R310 B.n397 B.n396 163.367
R311 B.n396 B.n49 163.367
R312 B.n392 B.n49 163.367
R313 B.n392 B.n391 163.367
R314 B.n391 B.n390 163.367
R315 B.n390 B.n51 163.367
R316 B.n386 B.n51 163.367
R317 B.n386 B.n385 163.367
R318 B.n385 B.n384 163.367
R319 B.n384 B.n53 163.367
R320 B.n380 B.n53 163.367
R321 B.n380 B.n379 163.367
R322 B.n379 B.n378 163.367
R323 B.n378 B.n55 163.367
R324 B.n374 B.n55 163.367
R325 B.n374 B.n373 163.367
R326 B.n373 B.n372 163.367
R327 B.n372 B.n57 163.367
R328 B.n368 B.n57 163.367
R329 B.n368 B.n367 163.367
R330 B.n367 B.n366 163.367
R331 B.n366 B.n59 163.367
R332 B.n362 B.n59 163.367
R333 B.n362 B.n361 163.367
R334 B.n361 B.n360 163.367
R335 B.n360 B.n61 163.367
R336 B.n356 B.n61 163.367
R337 B.n356 B.n355 163.367
R338 B.n355 B.n354 163.367
R339 B.n354 B.n63 163.367
R340 B.n350 B.n63 163.367
R341 B.n350 B.n349 163.367
R342 B.n349 B.n348 163.367
R343 B.n348 B.n65 163.367
R344 B.n344 B.n65 163.367
R345 B.n344 B.n343 163.367
R346 B.n343 B.n342 163.367
R347 B.n342 B.n67 163.367
R348 B.n338 B.n67 163.367
R349 B.n338 B.n337 163.367
R350 B.n337 B.n336 163.367
R351 B.n336 B.n69 163.367
R352 B.n332 B.n69 163.367
R353 B.n332 B.n331 163.367
R354 B.n331 B.n330 163.367
R355 B.n330 B.n71 163.367
R356 B.n326 B.n71 163.367
R357 B.n326 B.n325 163.367
R358 B.n325 B.n324 163.367
R359 B.n324 B.n73 163.367
R360 B.n320 B.n73 163.367
R361 B.n320 B.n319 163.367
R362 B.n319 B.n318 163.367
R363 B.n318 B.n75 163.367
R364 B.n314 B.n75 163.367
R365 B.n314 B.n313 163.367
R366 B.n313 B.n312 163.367
R367 B.n312 B.n77 163.367
R368 B.n308 B.n77 163.367
R369 B.n308 B.n307 163.367
R370 B.n307 B.n306 163.367
R371 B.n306 B.n79 163.367
R372 B.n302 B.n79 163.367
R373 B.n302 B.n301 163.367
R374 B.n301 B.n300 163.367
R375 B.n300 B.n81 163.367
R376 B.n296 B.n81 163.367
R377 B.n296 B.n295 163.367
R378 B.n295 B.n294 163.367
R379 B.n294 B.n83 163.367
R380 B.n290 B.n83 163.367
R381 B.n290 B.n289 163.367
R382 B.n289 B.n288 163.367
R383 B.n288 B.n85 163.367
R384 B.n284 B.n85 163.367
R385 B.n284 B.n283 163.367
R386 B.n283 B.n282 163.367
R387 B.n282 B.n87 163.367
R388 B.n278 B.n87 163.367
R389 B.n278 B.n277 163.367
R390 B.n277 B.n276 163.367
R391 B.n276 B.n89 163.367
R392 B.n272 B.n89 163.367
R393 B.n272 B.n271 163.367
R394 B.n271 B.n270 163.367
R395 B.n270 B.n91 163.367
R396 B.n266 B.n91 163.367
R397 B.n266 B.n265 163.367
R398 B.n265 B.n264 163.367
R399 B.n264 B.n93 163.367
R400 B.n260 B.n93 163.367
R401 B.n260 B.n259 163.367
R402 B.n452 B.n451 163.367
R403 B.n451 B.n450 163.367
R404 B.n450 B.n27 163.367
R405 B.n446 B.n27 163.367
R406 B.n446 B.n445 163.367
R407 B.n445 B.n444 163.367
R408 B.n444 B.n29 163.367
R409 B.n440 B.n29 163.367
R410 B.n440 B.n439 163.367
R411 B.n439 B.n438 163.367
R412 B.n438 B.n31 163.367
R413 B.n433 B.n31 163.367
R414 B.n433 B.n432 163.367
R415 B.n432 B.n431 163.367
R416 B.n431 B.n35 163.367
R417 B.n427 B.n35 163.367
R418 B.n427 B.n426 163.367
R419 B.n426 B.n425 163.367
R420 B.n425 B.n37 163.367
R421 B.n421 B.n37 163.367
R422 B.n421 B.n420 163.367
R423 B.n420 B.n41 163.367
R424 B.n416 B.n41 163.367
R425 B.n416 B.n415 163.367
R426 B.n415 B.n414 163.367
R427 B.n414 B.n43 163.367
R428 B.n410 B.n43 163.367
R429 B.n410 B.n409 163.367
R430 B.n409 B.n408 163.367
R431 B.n408 B.n45 163.367
R432 B.n404 B.n45 163.367
R433 B.n404 B.n403 163.367
R434 B.n456 B.n25 163.367
R435 B.n457 B.n456 163.367
R436 B.n458 B.n457 163.367
R437 B.n458 B.n23 163.367
R438 B.n462 B.n23 163.367
R439 B.n463 B.n462 163.367
R440 B.n464 B.n463 163.367
R441 B.n464 B.n21 163.367
R442 B.n468 B.n21 163.367
R443 B.n469 B.n468 163.367
R444 B.n470 B.n469 163.367
R445 B.n470 B.n19 163.367
R446 B.n474 B.n19 163.367
R447 B.n475 B.n474 163.367
R448 B.n476 B.n475 163.367
R449 B.n476 B.n17 163.367
R450 B.n480 B.n17 163.367
R451 B.n481 B.n480 163.367
R452 B.n482 B.n481 163.367
R453 B.n482 B.n15 163.367
R454 B.n486 B.n15 163.367
R455 B.n487 B.n486 163.367
R456 B.n488 B.n487 163.367
R457 B.n488 B.n13 163.367
R458 B.n492 B.n13 163.367
R459 B.n493 B.n492 163.367
R460 B.n494 B.n493 163.367
R461 B.n494 B.n11 163.367
R462 B.n498 B.n11 163.367
R463 B.n499 B.n498 163.367
R464 B.n500 B.n499 163.367
R465 B.n500 B.n9 163.367
R466 B.n504 B.n9 163.367
R467 B.n505 B.n504 163.367
R468 B.n506 B.n505 163.367
R469 B.n506 B.n7 163.367
R470 B.n510 B.n7 163.367
R471 B.n511 B.n510 163.367
R472 B.n512 B.n511 163.367
R473 B.n512 B.n5 163.367
R474 B.n516 B.n5 163.367
R475 B.n517 B.n516 163.367
R476 B.n518 B.n517 163.367
R477 B.n518 B.n3 163.367
R478 B.n522 B.n3 163.367
R479 B.n523 B.n522 163.367
R480 B.n136 B.n2 163.367
R481 B.n136 B.n135 163.367
R482 B.n140 B.n135 163.367
R483 B.n141 B.n140 163.367
R484 B.n142 B.n141 163.367
R485 B.n142 B.n133 163.367
R486 B.n146 B.n133 163.367
R487 B.n147 B.n146 163.367
R488 B.n148 B.n147 163.367
R489 B.n148 B.n131 163.367
R490 B.n152 B.n131 163.367
R491 B.n153 B.n152 163.367
R492 B.n154 B.n153 163.367
R493 B.n154 B.n129 163.367
R494 B.n158 B.n129 163.367
R495 B.n159 B.n158 163.367
R496 B.n160 B.n159 163.367
R497 B.n160 B.n127 163.367
R498 B.n164 B.n127 163.367
R499 B.n165 B.n164 163.367
R500 B.n166 B.n165 163.367
R501 B.n166 B.n125 163.367
R502 B.n170 B.n125 163.367
R503 B.n171 B.n170 163.367
R504 B.n172 B.n171 163.367
R505 B.n172 B.n123 163.367
R506 B.n176 B.n123 163.367
R507 B.n177 B.n176 163.367
R508 B.n178 B.n177 163.367
R509 B.n178 B.n121 163.367
R510 B.n182 B.n121 163.367
R511 B.n183 B.n182 163.367
R512 B.n184 B.n183 163.367
R513 B.n184 B.n119 163.367
R514 B.n188 B.n119 163.367
R515 B.n189 B.n188 163.367
R516 B.n190 B.n189 163.367
R517 B.n190 B.n117 163.367
R518 B.n194 B.n117 163.367
R519 B.n195 B.n194 163.367
R520 B.n196 B.n195 163.367
R521 B.n196 B.n115 163.367
R522 B.n200 B.n115 163.367
R523 B.n201 B.n200 163.367
R524 B.n202 B.n201 163.367
R525 B.n202 B.n113 163.367
R526 B.n107 B.n106 65.3581
R527 B.n237 B.n236 65.3581
R528 B.n39 B.n38 65.3581
R529 B.n33 B.n32 65.3581
R530 B.n223 B.n107 59.5399
R531 B.n238 B.n237 59.5399
R532 B.n40 B.n39 59.5399
R533 B.n435 B.n33 59.5399
R534 B.n454 B.n453 37.3078
R535 B.n401 B.n46 37.3078
R536 B.n257 B.n94 37.3078
R537 B.n205 B.n204 37.3078
R538 B B.n525 18.0485
R539 B.n455 B.n454 10.6151
R540 B.n455 B.n24 10.6151
R541 B.n459 B.n24 10.6151
R542 B.n460 B.n459 10.6151
R543 B.n461 B.n460 10.6151
R544 B.n461 B.n22 10.6151
R545 B.n465 B.n22 10.6151
R546 B.n466 B.n465 10.6151
R547 B.n467 B.n466 10.6151
R548 B.n467 B.n20 10.6151
R549 B.n471 B.n20 10.6151
R550 B.n472 B.n471 10.6151
R551 B.n473 B.n472 10.6151
R552 B.n473 B.n18 10.6151
R553 B.n477 B.n18 10.6151
R554 B.n478 B.n477 10.6151
R555 B.n479 B.n478 10.6151
R556 B.n479 B.n16 10.6151
R557 B.n483 B.n16 10.6151
R558 B.n484 B.n483 10.6151
R559 B.n485 B.n484 10.6151
R560 B.n485 B.n14 10.6151
R561 B.n489 B.n14 10.6151
R562 B.n490 B.n489 10.6151
R563 B.n491 B.n490 10.6151
R564 B.n491 B.n12 10.6151
R565 B.n495 B.n12 10.6151
R566 B.n496 B.n495 10.6151
R567 B.n497 B.n496 10.6151
R568 B.n497 B.n10 10.6151
R569 B.n501 B.n10 10.6151
R570 B.n502 B.n501 10.6151
R571 B.n503 B.n502 10.6151
R572 B.n503 B.n8 10.6151
R573 B.n507 B.n8 10.6151
R574 B.n508 B.n507 10.6151
R575 B.n509 B.n508 10.6151
R576 B.n509 B.n6 10.6151
R577 B.n513 B.n6 10.6151
R578 B.n514 B.n513 10.6151
R579 B.n515 B.n514 10.6151
R580 B.n515 B.n4 10.6151
R581 B.n519 B.n4 10.6151
R582 B.n520 B.n519 10.6151
R583 B.n521 B.n520 10.6151
R584 B.n521 B.n0 10.6151
R585 B.n453 B.n26 10.6151
R586 B.n449 B.n26 10.6151
R587 B.n449 B.n448 10.6151
R588 B.n448 B.n447 10.6151
R589 B.n447 B.n28 10.6151
R590 B.n443 B.n28 10.6151
R591 B.n443 B.n442 10.6151
R592 B.n442 B.n441 10.6151
R593 B.n441 B.n30 10.6151
R594 B.n437 B.n30 10.6151
R595 B.n437 B.n436 10.6151
R596 B.n434 B.n34 10.6151
R597 B.n430 B.n34 10.6151
R598 B.n430 B.n429 10.6151
R599 B.n429 B.n428 10.6151
R600 B.n428 B.n36 10.6151
R601 B.n424 B.n36 10.6151
R602 B.n424 B.n423 10.6151
R603 B.n423 B.n422 10.6151
R604 B.n419 B.n418 10.6151
R605 B.n418 B.n417 10.6151
R606 B.n417 B.n42 10.6151
R607 B.n413 B.n42 10.6151
R608 B.n413 B.n412 10.6151
R609 B.n412 B.n411 10.6151
R610 B.n411 B.n44 10.6151
R611 B.n407 B.n44 10.6151
R612 B.n407 B.n406 10.6151
R613 B.n406 B.n405 10.6151
R614 B.n405 B.n46 10.6151
R615 B.n401 B.n400 10.6151
R616 B.n400 B.n399 10.6151
R617 B.n399 B.n48 10.6151
R618 B.n395 B.n48 10.6151
R619 B.n395 B.n394 10.6151
R620 B.n394 B.n393 10.6151
R621 B.n393 B.n50 10.6151
R622 B.n389 B.n50 10.6151
R623 B.n389 B.n388 10.6151
R624 B.n388 B.n387 10.6151
R625 B.n387 B.n52 10.6151
R626 B.n383 B.n52 10.6151
R627 B.n383 B.n382 10.6151
R628 B.n382 B.n381 10.6151
R629 B.n381 B.n54 10.6151
R630 B.n377 B.n54 10.6151
R631 B.n377 B.n376 10.6151
R632 B.n376 B.n375 10.6151
R633 B.n375 B.n56 10.6151
R634 B.n371 B.n56 10.6151
R635 B.n371 B.n370 10.6151
R636 B.n370 B.n369 10.6151
R637 B.n369 B.n58 10.6151
R638 B.n365 B.n58 10.6151
R639 B.n365 B.n364 10.6151
R640 B.n364 B.n363 10.6151
R641 B.n363 B.n60 10.6151
R642 B.n359 B.n60 10.6151
R643 B.n359 B.n358 10.6151
R644 B.n358 B.n357 10.6151
R645 B.n357 B.n62 10.6151
R646 B.n353 B.n62 10.6151
R647 B.n353 B.n352 10.6151
R648 B.n352 B.n351 10.6151
R649 B.n351 B.n64 10.6151
R650 B.n347 B.n64 10.6151
R651 B.n347 B.n346 10.6151
R652 B.n346 B.n345 10.6151
R653 B.n345 B.n66 10.6151
R654 B.n341 B.n66 10.6151
R655 B.n341 B.n340 10.6151
R656 B.n340 B.n339 10.6151
R657 B.n339 B.n68 10.6151
R658 B.n335 B.n68 10.6151
R659 B.n335 B.n334 10.6151
R660 B.n334 B.n333 10.6151
R661 B.n333 B.n70 10.6151
R662 B.n329 B.n70 10.6151
R663 B.n329 B.n328 10.6151
R664 B.n328 B.n327 10.6151
R665 B.n327 B.n72 10.6151
R666 B.n323 B.n72 10.6151
R667 B.n323 B.n322 10.6151
R668 B.n322 B.n321 10.6151
R669 B.n321 B.n74 10.6151
R670 B.n317 B.n74 10.6151
R671 B.n317 B.n316 10.6151
R672 B.n316 B.n315 10.6151
R673 B.n315 B.n76 10.6151
R674 B.n311 B.n76 10.6151
R675 B.n311 B.n310 10.6151
R676 B.n310 B.n309 10.6151
R677 B.n309 B.n78 10.6151
R678 B.n305 B.n78 10.6151
R679 B.n305 B.n304 10.6151
R680 B.n304 B.n303 10.6151
R681 B.n303 B.n80 10.6151
R682 B.n299 B.n80 10.6151
R683 B.n299 B.n298 10.6151
R684 B.n298 B.n297 10.6151
R685 B.n297 B.n82 10.6151
R686 B.n293 B.n82 10.6151
R687 B.n293 B.n292 10.6151
R688 B.n292 B.n291 10.6151
R689 B.n291 B.n84 10.6151
R690 B.n287 B.n84 10.6151
R691 B.n287 B.n286 10.6151
R692 B.n286 B.n285 10.6151
R693 B.n285 B.n86 10.6151
R694 B.n281 B.n86 10.6151
R695 B.n281 B.n280 10.6151
R696 B.n280 B.n279 10.6151
R697 B.n279 B.n88 10.6151
R698 B.n275 B.n88 10.6151
R699 B.n275 B.n274 10.6151
R700 B.n274 B.n273 10.6151
R701 B.n273 B.n90 10.6151
R702 B.n269 B.n90 10.6151
R703 B.n269 B.n268 10.6151
R704 B.n268 B.n267 10.6151
R705 B.n267 B.n92 10.6151
R706 B.n263 B.n92 10.6151
R707 B.n263 B.n262 10.6151
R708 B.n262 B.n261 10.6151
R709 B.n261 B.n94 10.6151
R710 B.n137 B.n1 10.6151
R711 B.n138 B.n137 10.6151
R712 B.n139 B.n138 10.6151
R713 B.n139 B.n134 10.6151
R714 B.n143 B.n134 10.6151
R715 B.n144 B.n143 10.6151
R716 B.n145 B.n144 10.6151
R717 B.n145 B.n132 10.6151
R718 B.n149 B.n132 10.6151
R719 B.n150 B.n149 10.6151
R720 B.n151 B.n150 10.6151
R721 B.n151 B.n130 10.6151
R722 B.n155 B.n130 10.6151
R723 B.n156 B.n155 10.6151
R724 B.n157 B.n156 10.6151
R725 B.n157 B.n128 10.6151
R726 B.n161 B.n128 10.6151
R727 B.n162 B.n161 10.6151
R728 B.n163 B.n162 10.6151
R729 B.n163 B.n126 10.6151
R730 B.n167 B.n126 10.6151
R731 B.n168 B.n167 10.6151
R732 B.n169 B.n168 10.6151
R733 B.n169 B.n124 10.6151
R734 B.n173 B.n124 10.6151
R735 B.n174 B.n173 10.6151
R736 B.n175 B.n174 10.6151
R737 B.n175 B.n122 10.6151
R738 B.n179 B.n122 10.6151
R739 B.n180 B.n179 10.6151
R740 B.n181 B.n180 10.6151
R741 B.n181 B.n120 10.6151
R742 B.n185 B.n120 10.6151
R743 B.n186 B.n185 10.6151
R744 B.n187 B.n186 10.6151
R745 B.n187 B.n118 10.6151
R746 B.n191 B.n118 10.6151
R747 B.n192 B.n191 10.6151
R748 B.n193 B.n192 10.6151
R749 B.n193 B.n116 10.6151
R750 B.n197 B.n116 10.6151
R751 B.n198 B.n197 10.6151
R752 B.n199 B.n198 10.6151
R753 B.n199 B.n114 10.6151
R754 B.n203 B.n114 10.6151
R755 B.n204 B.n203 10.6151
R756 B.n205 B.n112 10.6151
R757 B.n209 B.n112 10.6151
R758 B.n210 B.n209 10.6151
R759 B.n211 B.n210 10.6151
R760 B.n211 B.n110 10.6151
R761 B.n215 B.n110 10.6151
R762 B.n216 B.n215 10.6151
R763 B.n217 B.n216 10.6151
R764 B.n217 B.n108 10.6151
R765 B.n221 B.n108 10.6151
R766 B.n222 B.n221 10.6151
R767 B.n224 B.n104 10.6151
R768 B.n228 B.n104 10.6151
R769 B.n229 B.n228 10.6151
R770 B.n230 B.n229 10.6151
R771 B.n230 B.n102 10.6151
R772 B.n234 B.n102 10.6151
R773 B.n235 B.n234 10.6151
R774 B.n239 B.n235 10.6151
R775 B.n243 B.n100 10.6151
R776 B.n244 B.n243 10.6151
R777 B.n245 B.n244 10.6151
R778 B.n245 B.n98 10.6151
R779 B.n249 B.n98 10.6151
R780 B.n250 B.n249 10.6151
R781 B.n251 B.n250 10.6151
R782 B.n251 B.n96 10.6151
R783 B.n255 B.n96 10.6151
R784 B.n256 B.n255 10.6151
R785 B.n257 B.n256 10.6151
R786 B.n525 B.n0 8.11757
R787 B.n525 B.n1 8.11757
R788 B.n435 B.n434 6.5566
R789 B.n422 B.n40 6.5566
R790 B.n224 B.n223 6.5566
R791 B.n239 B.n238 6.5566
R792 B.n436 B.n435 4.05904
R793 B.n419 B.n40 4.05904
R794 B.n223 B.n222 4.05904
R795 B.n238 B.n100 4.05904
R796 VP.n13 VP.n10 161.3
R797 VP.n15 VP.n14 161.3
R798 VP.n16 VP.n9 161.3
R799 VP.n18 VP.n17 161.3
R800 VP.n19 VP.n8 161.3
R801 VP.n21 VP.n20 161.3
R802 VP.n44 VP.n43 161.3
R803 VP.n42 VP.n1 161.3
R804 VP.n41 VP.n40 161.3
R805 VP.n39 VP.n2 161.3
R806 VP.n38 VP.n37 161.3
R807 VP.n36 VP.n3 161.3
R808 VP.n35 VP.n34 161.3
R809 VP.n33 VP.n4 161.3
R810 VP.n32 VP.n31 161.3
R811 VP.n30 VP.n5 161.3
R812 VP.n29 VP.n28 161.3
R813 VP.n27 VP.n6 161.3
R814 VP.n26 VP.n25 161.3
R815 VP.n24 VP.n23 72.0476
R816 VP.n45 VP.n0 72.0476
R817 VP.n22 VP.n7 72.0476
R818 VP.n30 VP.n29 56.5617
R819 VP.n41 VP.n2 56.5617
R820 VP.n18 VP.n9 56.5617
R821 VP.n12 VP.n11 49.4174
R822 VP.n11 VP.t5 48.4773
R823 VP.n23 VP.n22 42.8518
R824 VP.n25 VP.n6 24.5923
R825 VP.n29 VP.n6 24.5923
R826 VP.n31 VP.n30 24.5923
R827 VP.n31 VP.n4 24.5923
R828 VP.n35 VP.n4 24.5923
R829 VP.n36 VP.n35 24.5923
R830 VP.n37 VP.n36 24.5923
R831 VP.n37 VP.n2 24.5923
R832 VP.n42 VP.n41 24.5923
R833 VP.n43 VP.n42 24.5923
R834 VP.n19 VP.n18 24.5923
R835 VP.n20 VP.n19 24.5923
R836 VP.n13 VP.n12 24.5923
R837 VP.n14 VP.n13 24.5923
R838 VP.n14 VP.n9 24.5923
R839 VP.n25 VP.n24 18.1985
R840 VP.n43 VP.n0 18.1985
R841 VP.n20 VP.n7 18.1985
R842 VP.n35 VP.t4 15.063
R843 VP.n24 VP.t1 15.063
R844 VP.n0 VP.t3 15.063
R845 VP.n12 VP.t2 15.063
R846 VP.n7 VP.t0 15.063
R847 VP.n11 VP.n10 3.99106
R848 VP.n22 VP.n21 0.354861
R849 VP.n26 VP.n23 0.354861
R850 VP.n45 VP.n44 0.354861
R851 VP VP.n45 0.267071
R852 VP.n15 VP.n10 0.189894
R853 VP.n16 VP.n15 0.189894
R854 VP.n17 VP.n16 0.189894
R855 VP.n17 VP.n8 0.189894
R856 VP.n21 VP.n8 0.189894
R857 VP.n27 VP.n26 0.189894
R858 VP.n28 VP.n27 0.189894
R859 VP.n28 VP.n5 0.189894
R860 VP.n32 VP.n5 0.189894
R861 VP.n33 VP.n32 0.189894
R862 VP.n34 VP.n33 0.189894
R863 VP.n34 VP.n3 0.189894
R864 VP.n38 VP.n3 0.189894
R865 VP.n39 VP.n38 0.189894
R866 VP.n40 VP.n39 0.189894
R867 VP.n40 VP.n1 0.189894
R868 VP.n44 VP.n1 0.189894
R869 VTAIL.n34 VTAIL.n32 756.745
R870 VTAIL.n4 VTAIL.n2 756.745
R871 VTAIL.n26 VTAIL.n24 756.745
R872 VTAIL.n16 VTAIL.n14 756.745
R873 VTAIL.n35 VTAIL.n34 585
R874 VTAIL.n5 VTAIL.n4 585
R875 VTAIL.n27 VTAIL.n26 585
R876 VTAIL.n17 VTAIL.n16 585
R877 VTAIL.t3 VTAIL.n33 415.613
R878 VTAIL.t11 VTAIL.n3 415.613
R879 VTAIL.t7 VTAIL.n25 415.613
R880 VTAIL.t1 VTAIL.n15 415.613
R881 VTAIL.n23 VTAIL.n22 187.147
R882 VTAIL.n13 VTAIL.n12 187.147
R883 VTAIL.n1 VTAIL.n0 187.147
R884 VTAIL.n11 VTAIL.n10 187.147
R885 VTAIL.n34 VTAIL.t3 85.8723
R886 VTAIL.n4 VTAIL.t11 85.8723
R887 VTAIL.n26 VTAIL.t7 85.8723
R888 VTAIL.n16 VTAIL.t1 85.8723
R889 VTAIL.n39 VTAIL.n38 36.452
R890 VTAIL.n9 VTAIL.n8 36.452
R891 VTAIL.n31 VTAIL.n30 36.452
R892 VTAIL.n21 VTAIL.n20 36.452
R893 VTAIL.n13 VTAIL.n11 19.8152
R894 VTAIL.n0 VTAIL.t0 17.1084
R895 VTAIL.n0 VTAIL.t4 17.1084
R896 VTAIL.n10 VTAIL.t6 17.1084
R897 VTAIL.n10 VTAIL.t9 17.1084
R898 VTAIL.n22 VTAIL.t8 17.1084
R899 VTAIL.n22 VTAIL.t10 17.1084
R900 VTAIL.n12 VTAIL.t2 17.1084
R901 VTAIL.n12 VTAIL.t5 17.1084
R902 VTAIL.n39 VTAIL.n31 16.91
R903 VTAIL.n35 VTAIL.n33 14.9339
R904 VTAIL.n5 VTAIL.n3 14.9339
R905 VTAIL.n27 VTAIL.n25 14.9339
R906 VTAIL.n17 VTAIL.n15 14.9339
R907 VTAIL.n36 VTAIL.n32 12.8005
R908 VTAIL.n6 VTAIL.n2 12.8005
R909 VTAIL.n28 VTAIL.n24 12.8005
R910 VTAIL.n18 VTAIL.n14 12.8005
R911 VTAIL.n38 VTAIL.n37 9.45567
R912 VTAIL.n8 VTAIL.n7 9.45567
R913 VTAIL.n30 VTAIL.n29 9.45567
R914 VTAIL.n20 VTAIL.n19 9.45567
R915 VTAIL.n37 VTAIL.n36 9.3005
R916 VTAIL.n7 VTAIL.n6 9.3005
R917 VTAIL.n29 VTAIL.n28 9.3005
R918 VTAIL.n19 VTAIL.n18 9.3005
R919 VTAIL.n37 VTAIL.n33 5.44463
R920 VTAIL.n7 VTAIL.n3 5.44463
R921 VTAIL.n29 VTAIL.n25 5.44463
R922 VTAIL.n19 VTAIL.n15 5.44463
R923 VTAIL.n21 VTAIL.n13 2.90567
R924 VTAIL.n31 VTAIL.n23 2.90567
R925 VTAIL.n11 VTAIL.n9 2.90567
R926 VTAIL VTAIL.n39 2.12119
R927 VTAIL.n23 VTAIL.n21 1.92291
R928 VTAIL.n9 VTAIL.n1 1.92291
R929 VTAIL.n38 VTAIL.n32 1.16414
R930 VTAIL.n8 VTAIL.n2 1.16414
R931 VTAIL.n30 VTAIL.n24 1.16414
R932 VTAIL.n20 VTAIL.n14 1.16414
R933 VTAIL VTAIL.n1 0.784983
R934 VTAIL.n36 VTAIL.n35 0.388379
R935 VTAIL.n6 VTAIL.n5 0.388379
R936 VTAIL.n28 VTAIL.n27 0.388379
R937 VTAIL.n18 VTAIL.n17 0.388379
R938 VDD1.n2 VDD1.n0 756.745
R939 VDD1.n9 VDD1.n7 756.745
R940 VDD1.n3 VDD1.n2 585
R941 VDD1.n10 VDD1.n9 585
R942 VDD1.t4 VDD1.n8 415.613
R943 VDD1.t0 VDD1.n1 415.613
R944 VDD1.n15 VDD1.n14 204.496
R945 VDD1.n17 VDD1.n16 203.826
R946 VDD1.n2 VDD1.t0 85.8723
R947 VDD1.n9 VDD1.t4 85.8723
R948 VDD1 VDD1.n6 55.3679
R949 VDD1.n15 VDD1.n13 55.2543
R950 VDD1.n17 VDD1.n15 36.8306
R951 VDD1.n16 VDD1.t3 17.1084
R952 VDD1.n16 VDD1.t5 17.1084
R953 VDD1.n14 VDD1.t1 17.1084
R954 VDD1.n14 VDD1.t2 17.1084
R955 VDD1.n3 VDD1.n1 14.9339
R956 VDD1.n10 VDD1.n8 14.9339
R957 VDD1.n4 VDD1.n0 12.8005
R958 VDD1.n11 VDD1.n7 12.8005
R959 VDD1.n6 VDD1.n5 9.45567
R960 VDD1.n13 VDD1.n12 9.45567
R961 VDD1.n5 VDD1.n4 9.3005
R962 VDD1.n12 VDD1.n11 9.3005
R963 VDD1.n5 VDD1.n1 5.44463
R964 VDD1.n12 VDD1.n8 5.44463
R965 VDD1.n6 VDD1.n0 1.16414
R966 VDD1.n13 VDD1.n7 1.16414
R967 VDD1 VDD1.n17 0.668603
R968 VDD1.n4 VDD1.n3 0.388379
R969 VDD1.n11 VDD1.n10 0.388379
R970 VN.n30 VN.n29 161.3
R971 VN.n28 VN.n17 161.3
R972 VN.n27 VN.n26 161.3
R973 VN.n25 VN.n18 161.3
R974 VN.n24 VN.n23 161.3
R975 VN.n22 VN.n19 161.3
R976 VN.n14 VN.n13 161.3
R977 VN.n12 VN.n1 161.3
R978 VN.n11 VN.n10 161.3
R979 VN.n9 VN.n2 161.3
R980 VN.n8 VN.n7 161.3
R981 VN.n6 VN.n3 161.3
R982 VN.n15 VN.n0 72.0476
R983 VN.n31 VN.n16 72.0476
R984 VN.n11 VN.n2 56.5617
R985 VN.n27 VN.n18 56.5617
R986 VN.n5 VN.n4 49.4174
R987 VN.n21 VN.n20 49.4174
R988 VN.n20 VN.t1 48.4776
R989 VN.n4 VN.t5 48.4776
R990 VN VN.n31 43.0171
R991 VN.n6 VN.n5 24.5923
R992 VN.n7 VN.n6 24.5923
R993 VN.n7 VN.n2 24.5923
R994 VN.n12 VN.n11 24.5923
R995 VN.n13 VN.n12 24.5923
R996 VN.n23 VN.n18 24.5923
R997 VN.n23 VN.n22 24.5923
R998 VN.n22 VN.n21 24.5923
R999 VN.n29 VN.n28 24.5923
R1000 VN.n28 VN.n27 24.5923
R1001 VN.n13 VN.n0 18.1985
R1002 VN.n29 VN.n16 18.1985
R1003 VN.n5 VN.t2 15.063
R1004 VN.n0 VN.t0 15.063
R1005 VN.n21 VN.t3 15.063
R1006 VN.n16 VN.t4 15.063
R1007 VN.n20 VN.n19 3.99109
R1008 VN.n4 VN.n3 3.99108
R1009 VN.n31 VN.n30 0.354861
R1010 VN.n15 VN.n14 0.354861
R1011 VN VN.n15 0.267071
R1012 VN.n30 VN.n17 0.189894
R1013 VN.n26 VN.n17 0.189894
R1014 VN.n26 VN.n25 0.189894
R1015 VN.n25 VN.n24 0.189894
R1016 VN.n24 VN.n19 0.189894
R1017 VN.n8 VN.n3 0.189894
R1018 VN.n9 VN.n8 0.189894
R1019 VN.n10 VN.n9 0.189894
R1020 VN.n10 VN.n1 0.189894
R1021 VN.n14 VN.n1 0.189894
R1022 VDD2.n11 VDD2.n9 756.745
R1023 VDD2.n2 VDD2.n0 756.745
R1024 VDD2.n12 VDD2.n11 585
R1025 VDD2.n3 VDD2.n2 585
R1026 VDD2.t0 VDD2.n1 415.613
R1027 VDD2.t1 VDD2.n10 415.613
R1028 VDD2.n8 VDD2.n7 204.496
R1029 VDD2 VDD2.n17 204.494
R1030 VDD2.n11 VDD2.t1 85.8723
R1031 VDD2.n2 VDD2.t0 85.8723
R1032 VDD2.n8 VDD2.n6 55.2543
R1033 VDD2.n16 VDD2.n15 53.1308
R1034 VDD2.n16 VDD2.n8 34.795
R1035 VDD2.n17 VDD2.t2 17.1084
R1036 VDD2.n17 VDD2.t4 17.1084
R1037 VDD2.n7 VDD2.t3 17.1084
R1038 VDD2.n7 VDD2.t5 17.1084
R1039 VDD2.n12 VDD2.n10 14.9339
R1040 VDD2.n3 VDD2.n1 14.9339
R1041 VDD2.n13 VDD2.n9 12.8005
R1042 VDD2.n4 VDD2.n0 12.8005
R1043 VDD2.n15 VDD2.n14 9.45567
R1044 VDD2.n6 VDD2.n5 9.45567
R1045 VDD2.n14 VDD2.n13 9.3005
R1046 VDD2.n5 VDD2.n4 9.3005
R1047 VDD2.n14 VDD2.n10 5.44463
R1048 VDD2.n5 VDD2.n1 5.44463
R1049 VDD2 VDD2.n16 2.23757
R1050 VDD2.n15 VDD2.n9 1.16414
R1051 VDD2.n6 VDD2.n0 1.16414
R1052 VDD2.n13 VDD2.n12 0.388379
R1053 VDD2.n4 VDD2.n3 0.388379
C0 VTAIL B 1.42335f
C1 w_n3666_n1348# VDD2 1.79514f
C2 VP VN 5.48897f
C3 VDD1 w_n3666_n1348# 1.69677f
C4 VDD2 VN 1.42718f
C5 VP VDD2 0.503035f
C6 VDD1 VN 0.15828f
C7 w_n3666_n1348# B 7.506061f
C8 VDD1 VP 1.76896f
C9 VDD1 VDD2 1.57818f
C10 w_n3666_n1348# VTAIL 1.57559f
C11 B VN 1.13065f
C12 VP B 1.92545f
C13 B VDD2 1.48648f
C14 VTAIL VN 2.44305f
C15 VP VTAIL 2.45718f
C16 VDD1 B 1.40141f
C17 VTAIL VDD2 4.43662f
C18 VDD1 VTAIL 4.38041f
C19 w_n3666_n1348# VN 6.86571f
C20 VP w_n3666_n1348# 7.335979f
C21 VDD2 VSUBS 1.135835f
C22 VDD1 VSUBS 1.469708f
C23 VTAIL VSUBS 0.585515f
C24 VN VSUBS 6.2199f
C25 VP VSUBS 2.690371f
C26 B VSUBS 3.962801f
C27 w_n3666_n1348# VSUBS 63.128498f
C28 VDD2.n0 VSUBS 0.018525f
C29 VDD2.n1 VSUBS 0.049922f
C30 VDD2.t0 VSUBS 0.047731f
C31 VDD2.n2 VSUBS 0.046294f
C32 VDD2.n3 VSUBS 0.011506f
C33 VDD2.n4 VSUBS 0.009165f
C34 VDD2.n5 VSUBS 0.107002f
C35 VDD2.n6 VSUBS 0.043731f
C36 VDD2.t3 VSUBS 0.025609f
C37 VDD2.t5 VSUBS 0.025609f
C38 VDD2.n7 VSUBS 0.110256f
C39 VDD2.n8 VSUBS 1.58713f
C40 VDD2.n9 VSUBS 0.018525f
C41 VDD2.n10 VSUBS 0.049922f
C42 VDD2.t1 VSUBS 0.047731f
C43 VDD2.n11 VSUBS 0.046294f
C44 VDD2.n12 VSUBS 0.011506f
C45 VDD2.n13 VSUBS 0.009165f
C46 VDD2.n14 VSUBS 0.107002f
C47 VDD2.n15 VSUBS 0.037863f
C48 VDD2.n16 VSUBS 1.2883f
C49 VDD2.t2 VSUBS 0.025609f
C50 VDD2.t4 VSUBS 0.025609f
C51 VDD2.n17 VSUBS 0.110248f
C52 VN.t0 VSUBS 0.649157f
C53 VN.n0 VSUBS 0.493922f
C54 VN.n1 VSUBS 0.048636f
C55 VN.n2 VSUBS 0.061953f
C56 VN.n3 VSUBS 0.553028f
C57 VN.t2 VSUBS 0.649157f
C58 VN.t5 VSUBS 1.09219f
C59 VN.n4 VSUBS 0.47305f
C60 VN.n5 VSUBS 0.487f
C61 VN.n6 VSUBS 0.090191f
C62 VN.n7 VSUBS 0.090191f
C63 VN.n8 VSUBS 0.048636f
C64 VN.n9 VSUBS 0.048636f
C65 VN.n10 VSUBS 0.048636f
C66 VN.n11 VSUBS 0.079447f
C67 VN.n12 VSUBS 0.090191f
C68 VN.n13 VSUBS 0.078615f
C69 VN.n14 VSUBS 0.078485f
C70 VN.n15 VSUBS 0.105846f
C71 VN.t4 VSUBS 0.649157f
C72 VN.n16 VSUBS 0.493922f
C73 VN.n17 VSUBS 0.048636f
C74 VN.n18 VSUBS 0.061953f
C75 VN.n19 VSUBS 0.553028f
C76 VN.t3 VSUBS 0.649157f
C77 VN.t1 VSUBS 1.09219f
C78 VN.n20 VSUBS 0.47305f
C79 VN.n21 VSUBS 0.487f
C80 VN.n22 VSUBS 0.090191f
C81 VN.n23 VSUBS 0.090191f
C82 VN.n24 VSUBS 0.048636f
C83 VN.n25 VSUBS 0.048636f
C84 VN.n26 VSUBS 0.048636f
C85 VN.n27 VSUBS 0.079447f
C86 VN.n28 VSUBS 0.090191f
C87 VN.n29 VSUBS 0.078615f
C88 VN.n30 VSUBS 0.078485f
C89 VN.n31 VSUBS 2.20528f
C90 VDD1.n0 VSUBS 0.018264f
C91 VDD1.n1 VSUBS 0.049217f
C92 VDD1.t0 VSUBS 0.047057f
C93 VDD1.n2 VSUBS 0.04564f
C94 VDD1.n3 VSUBS 0.011343f
C95 VDD1.n4 VSUBS 0.009036f
C96 VDD1.n5 VSUBS 0.105492f
C97 VDD1.n6 VSUBS 0.043651f
C98 VDD1.n7 VSUBS 0.018264f
C99 VDD1.n8 VSUBS 0.049217f
C100 VDD1.t4 VSUBS 0.047057f
C101 VDD1.n9 VSUBS 0.04564f
C102 VDD1.n10 VSUBS 0.011343f
C103 VDD1.n11 VSUBS 0.009036f
C104 VDD1.n12 VSUBS 0.105492f
C105 VDD1.n13 VSUBS 0.043113f
C106 VDD1.t1 VSUBS 0.025248f
C107 VDD1.t2 VSUBS 0.025248f
C108 VDD1.n14 VSUBS 0.108699f
C109 VDD1.n15 VSUBS 1.64818f
C110 VDD1.t3 VSUBS 0.025248f
C111 VDD1.t5 VSUBS 0.025248f
C112 VDD1.n16 VSUBS 0.107464f
C113 VDD1.n17 VSUBS 1.46823f
C114 VTAIL.t0 VSUBS 0.053645f
C115 VTAIL.t4 VSUBS 0.053645f
C116 VTAIL.n0 VSUBS 0.195694f
C117 VTAIL.n1 VSUBS 0.668727f
C118 VTAIL.n2 VSUBS 0.038806f
C119 VTAIL.n3 VSUBS 0.104573f
C120 VTAIL.t11 VSUBS 0.099984f
C121 VTAIL.n4 VSUBS 0.096974f
C122 VTAIL.n5 VSUBS 0.024102f
C123 VTAIL.n6 VSUBS 0.019199f
C124 VTAIL.n7 VSUBS 0.224142f
C125 VTAIL.n8 VSUBS 0.054716f
C126 VTAIL.n9 VSUBS 0.592374f
C127 VTAIL.t6 VSUBS 0.053645f
C128 VTAIL.t9 VSUBS 0.053645f
C129 VTAIL.n10 VSUBS 0.195694f
C130 VTAIL.n11 VSUBS 2.03438f
C131 VTAIL.t2 VSUBS 0.053645f
C132 VTAIL.t5 VSUBS 0.053645f
C133 VTAIL.n12 VSUBS 0.195695f
C134 VTAIL.n13 VSUBS 2.03438f
C135 VTAIL.n14 VSUBS 0.038806f
C136 VTAIL.n15 VSUBS 0.104573f
C137 VTAIL.t1 VSUBS 0.099984f
C138 VTAIL.n16 VSUBS 0.096974f
C139 VTAIL.n17 VSUBS 0.024102f
C140 VTAIL.n18 VSUBS 0.019199f
C141 VTAIL.n19 VSUBS 0.224142f
C142 VTAIL.n20 VSUBS 0.054716f
C143 VTAIL.n21 VSUBS 0.592374f
C144 VTAIL.t8 VSUBS 0.053645f
C145 VTAIL.t10 VSUBS 0.053645f
C146 VTAIL.n22 VSUBS 0.195695f
C147 VTAIL.n23 VSUBS 0.912873f
C148 VTAIL.n24 VSUBS 0.038806f
C149 VTAIL.n25 VSUBS 0.104573f
C150 VTAIL.t7 VSUBS 0.099984f
C151 VTAIL.n26 VSUBS 0.096974f
C152 VTAIL.n27 VSUBS 0.024102f
C153 VTAIL.n28 VSUBS 0.019199f
C154 VTAIL.n29 VSUBS 0.224142f
C155 VTAIL.n30 VSUBS 0.054716f
C156 VTAIL.n31 VSUBS 1.37942f
C157 VTAIL.n32 VSUBS 0.038806f
C158 VTAIL.n33 VSUBS 0.104573f
C159 VTAIL.t3 VSUBS 0.099984f
C160 VTAIL.n34 VSUBS 0.096974f
C161 VTAIL.n35 VSUBS 0.024102f
C162 VTAIL.n36 VSUBS 0.019199f
C163 VTAIL.n37 VSUBS 0.224142f
C164 VTAIL.n38 VSUBS 0.054716f
C165 VTAIL.n39 VSUBS 1.2891f
C166 VP.t3 VSUBS 0.674202f
C167 VP.n0 VSUBS 0.512978f
C168 VP.n1 VSUBS 0.050513f
C169 VP.n2 VSUBS 0.064344f
C170 VP.n3 VSUBS 0.050513f
C171 VP.t4 VSUBS 0.674202f
C172 VP.n4 VSUBS 0.093671f
C173 VP.n5 VSUBS 0.050513f
C174 VP.n6 VSUBS 0.093671f
C175 VP.t0 VSUBS 0.674202f
C176 VP.n7 VSUBS 0.512978f
C177 VP.n8 VSUBS 0.050513f
C178 VP.n9 VSUBS 0.064344f
C179 VP.n10 VSUBS 0.574366f
C180 VP.t2 VSUBS 0.674202f
C181 VP.t5 VSUBS 1.13432f
C182 VP.n11 VSUBS 0.491302f
C183 VP.n12 VSUBS 0.505789f
C184 VP.n13 VSUBS 0.093671f
C185 VP.n14 VSUBS 0.093671f
C186 VP.n15 VSUBS 0.050513f
C187 VP.n16 VSUBS 0.050513f
C188 VP.n17 VSUBS 0.050513f
C189 VP.n18 VSUBS 0.082512f
C190 VP.n19 VSUBS 0.093671f
C191 VP.n20 VSUBS 0.081648f
C192 VP.n21 VSUBS 0.081513f
C193 VP.n22 VSUBS 2.26851f
C194 VP.n23 VSUBS 2.311f
C195 VP.t1 VSUBS 0.674202f
C196 VP.n24 VSUBS 0.512978f
C197 VP.n25 VSUBS 0.081648f
C198 VP.n26 VSUBS 0.081513f
C199 VP.n27 VSUBS 0.050513f
C200 VP.n28 VSUBS 0.050513f
C201 VP.n29 VSUBS 0.082512f
C202 VP.n30 VSUBS 0.064344f
C203 VP.n31 VSUBS 0.093671f
C204 VP.n32 VSUBS 0.050513f
C205 VP.n33 VSUBS 0.050513f
C206 VP.n34 VSUBS 0.050513f
C207 VP.n35 VSUBS 0.366221f
C208 VP.n36 VSUBS 0.093671f
C209 VP.n37 VSUBS 0.093671f
C210 VP.n38 VSUBS 0.050513f
C211 VP.n39 VSUBS 0.050513f
C212 VP.n40 VSUBS 0.050513f
C213 VP.n41 VSUBS 0.082512f
C214 VP.n42 VSUBS 0.093671f
C215 VP.n43 VSUBS 0.081648f
C216 VP.n44 VSUBS 0.081513f
C217 VP.n45 VSUBS 0.10993f
C218 B.n0 VSUBS 0.007852f
C219 B.n1 VSUBS 0.007852f
C220 B.n2 VSUBS 0.011612f
C221 B.n3 VSUBS 0.008898f
C222 B.n4 VSUBS 0.008898f
C223 B.n5 VSUBS 0.008898f
C224 B.n6 VSUBS 0.008898f
C225 B.n7 VSUBS 0.008898f
C226 B.n8 VSUBS 0.008898f
C227 B.n9 VSUBS 0.008898f
C228 B.n10 VSUBS 0.008898f
C229 B.n11 VSUBS 0.008898f
C230 B.n12 VSUBS 0.008898f
C231 B.n13 VSUBS 0.008898f
C232 B.n14 VSUBS 0.008898f
C233 B.n15 VSUBS 0.008898f
C234 B.n16 VSUBS 0.008898f
C235 B.n17 VSUBS 0.008898f
C236 B.n18 VSUBS 0.008898f
C237 B.n19 VSUBS 0.008898f
C238 B.n20 VSUBS 0.008898f
C239 B.n21 VSUBS 0.008898f
C240 B.n22 VSUBS 0.008898f
C241 B.n23 VSUBS 0.008898f
C242 B.n24 VSUBS 0.008898f
C243 B.n25 VSUBS 0.022287f
C244 B.n26 VSUBS 0.008898f
C245 B.n27 VSUBS 0.008898f
C246 B.n28 VSUBS 0.008898f
C247 B.n29 VSUBS 0.008898f
C248 B.n30 VSUBS 0.008898f
C249 B.n31 VSUBS 0.008898f
C250 B.t4 VSUBS 0.041034f
C251 B.t5 VSUBS 0.056292f
C252 B.t3 VSUBS 0.36309f
C253 B.n32 VSUBS 0.10558f
C254 B.n33 VSUBS 0.085471f
C255 B.n34 VSUBS 0.008898f
C256 B.n35 VSUBS 0.008898f
C257 B.n36 VSUBS 0.008898f
C258 B.n37 VSUBS 0.008898f
C259 B.t7 VSUBS 0.041034f
C260 B.t8 VSUBS 0.056292f
C261 B.t6 VSUBS 0.36309f
C262 B.n38 VSUBS 0.10558f
C263 B.n39 VSUBS 0.085471f
C264 B.n40 VSUBS 0.020617f
C265 B.n41 VSUBS 0.008898f
C266 B.n42 VSUBS 0.008898f
C267 B.n43 VSUBS 0.008898f
C268 B.n44 VSUBS 0.008898f
C269 B.n45 VSUBS 0.008898f
C270 B.n46 VSUBS 0.023252f
C271 B.n47 VSUBS 0.008898f
C272 B.n48 VSUBS 0.008898f
C273 B.n49 VSUBS 0.008898f
C274 B.n50 VSUBS 0.008898f
C275 B.n51 VSUBS 0.008898f
C276 B.n52 VSUBS 0.008898f
C277 B.n53 VSUBS 0.008898f
C278 B.n54 VSUBS 0.008898f
C279 B.n55 VSUBS 0.008898f
C280 B.n56 VSUBS 0.008898f
C281 B.n57 VSUBS 0.008898f
C282 B.n58 VSUBS 0.008898f
C283 B.n59 VSUBS 0.008898f
C284 B.n60 VSUBS 0.008898f
C285 B.n61 VSUBS 0.008898f
C286 B.n62 VSUBS 0.008898f
C287 B.n63 VSUBS 0.008898f
C288 B.n64 VSUBS 0.008898f
C289 B.n65 VSUBS 0.008898f
C290 B.n66 VSUBS 0.008898f
C291 B.n67 VSUBS 0.008898f
C292 B.n68 VSUBS 0.008898f
C293 B.n69 VSUBS 0.008898f
C294 B.n70 VSUBS 0.008898f
C295 B.n71 VSUBS 0.008898f
C296 B.n72 VSUBS 0.008898f
C297 B.n73 VSUBS 0.008898f
C298 B.n74 VSUBS 0.008898f
C299 B.n75 VSUBS 0.008898f
C300 B.n76 VSUBS 0.008898f
C301 B.n77 VSUBS 0.008898f
C302 B.n78 VSUBS 0.008898f
C303 B.n79 VSUBS 0.008898f
C304 B.n80 VSUBS 0.008898f
C305 B.n81 VSUBS 0.008898f
C306 B.n82 VSUBS 0.008898f
C307 B.n83 VSUBS 0.008898f
C308 B.n84 VSUBS 0.008898f
C309 B.n85 VSUBS 0.008898f
C310 B.n86 VSUBS 0.008898f
C311 B.n87 VSUBS 0.008898f
C312 B.n88 VSUBS 0.008898f
C313 B.n89 VSUBS 0.008898f
C314 B.n90 VSUBS 0.008898f
C315 B.n91 VSUBS 0.008898f
C316 B.n92 VSUBS 0.008898f
C317 B.n93 VSUBS 0.008898f
C318 B.n94 VSUBS 0.023207f
C319 B.n95 VSUBS 0.008898f
C320 B.n96 VSUBS 0.008898f
C321 B.n97 VSUBS 0.008898f
C322 B.n98 VSUBS 0.008898f
C323 B.n99 VSUBS 0.008898f
C324 B.n100 VSUBS 0.00615f
C325 B.n101 VSUBS 0.008898f
C326 B.n102 VSUBS 0.008898f
C327 B.n103 VSUBS 0.008898f
C328 B.n104 VSUBS 0.008898f
C329 B.n105 VSUBS 0.008898f
C330 B.t11 VSUBS 0.041034f
C331 B.t10 VSUBS 0.056292f
C332 B.t9 VSUBS 0.36309f
C333 B.n106 VSUBS 0.10558f
C334 B.n107 VSUBS 0.085471f
C335 B.n108 VSUBS 0.008898f
C336 B.n109 VSUBS 0.008898f
C337 B.n110 VSUBS 0.008898f
C338 B.n111 VSUBS 0.008898f
C339 B.n112 VSUBS 0.008898f
C340 B.n113 VSUBS 0.022287f
C341 B.n114 VSUBS 0.008898f
C342 B.n115 VSUBS 0.008898f
C343 B.n116 VSUBS 0.008898f
C344 B.n117 VSUBS 0.008898f
C345 B.n118 VSUBS 0.008898f
C346 B.n119 VSUBS 0.008898f
C347 B.n120 VSUBS 0.008898f
C348 B.n121 VSUBS 0.008898f
C349 B.n122 VSUBS 0.008898f
C350 B.n123 VSUBS 0.008898f
C351 B.n124 VSUBS 0.008898f
C352 B.n125 VSUBS 0.008898f
C353 B.n126 VSUBS 0.008898f
C354 B.n127 VSUBS 0.008898f
C355 B.n128 VSUBS 0.008898f
C356 B.n129 VSUBS 0.008898f
C357 B.n130 VSUBS 0.008898f
C358 B.n131 VSUBS 0.008898f
C359 B.n132 VSUBS 0.008898f
C360 B.n133 VSUBS 0.008898f
C361 B.n134 VSUBS 0.008898f
C362 B.n135 VSUBS 0.008898f
C363 B.n136 VSUBS 0.008898f
C364 B.n137 VSUBS 0.008898f
C365 B.n138 VSUBS 0.008898f
C366 B.n139 VSUBS 0.008898f
C367 B.n140 VSUBS 0.008898f
C368 B.n141 VSUBS 0.008898f
C369 B.n142 VSUBS 0.008898f
C370 B.n143 VSUBS 0.008898f
C371 B.n144 VSUBS 0.008898f
C372 B.n145 VSUBS 0.008898f
C373 B.n146 VSUBS 0.008898f
C374 B.n147 VSUBS 0.008898f
C375 B.n148 VSUBS 0.008898f
C376 B.n149 VSUBS 0.008898f
C377 B.n150 VSUBS 0.008898f
C378 B.n151 VSUBS 0.008898f
C379 B.n152 VSUBS 0.008898f
C380 B.n153 VSUBS 0.008898f
C381 B.n154 VSUBS 0.008898f
C382 B.n155 VSUBS 0.008898f
C383 B.n156 VSUBS 0.008898f
C384 B.n157 VSUBS 0.008898f
C385 B.n158 VSUBS 0.008898f
C386 B.n159 VSUBS 0.008898f
C387 B.n160 VSUBS 0.008898f
C388 B.n161 VSUBS 0.008898f
C389 B.n162 VSUBS 0.008898f
C390 B.n163 VSUBS 0.008898f
C391 B.n164 VSUBS 0.008898f
C392 B.n165 VSUBS 0.008898f
C393 B.n166 VSUBS 0.008898f
C394 B.n167 VSUBS 0.008898f
C395 B.n168 VSUBS 0.008898f
C396 B.n169 VSUBS 0.008898f
C397 B.n170 VSUBS 0.008898f
C398 B.n171 VSUBS 0.008898f
C399 B.n172 VSUBS 0.008898f
C400 B.n173 VSUBS 0.008898f
C401 B.n174 VSUBS 0.008898f
C402 B.n175 VSUBS 0.008898f
C403 B.n176 VSUBS 0.008898f
C404 B.n177 VSUBS 0.008898f
C405 B.n178 VSUBS 0.008898f
C406 B.n179 VSUBS 0.008898f
C407 B.n180 VSUBS 0.008898f
C408 B.n181 VSUBS 0.008898f
C409 B.n182 VSUBS 0.008898f
C410 B.n183 VSUBS 0.008898f
C411 B.n184 VSUBS 0.008898f
C412 B.n185 VSUBS 0.008898f
C413 B.n186 VSUBS 0.008898f
C414 B.n187 VSUBS 0.008898f
C415 B.n188 VSUBS 0.008898f
C416 B.n189 VSUBS 0.008898f
C417 B.n190 VSUBS 0.008898f
C418 B.n191 VSUBS 0.008898f
C419 B.n192 VSUBS 0.008898f
C420 B.n193 VSUBS 0.008898f
C421 B.n194 VSUBS 0.008898f
C422 B.n195 VSUBS 0.008898f
C423 B.n196 VSUBS 0.008898f
C424 B.n197 VSUBS 0.008898f
C425 B.n198 VSUBS 0.008898f
C426 B.n199 VSUBS 0.008898f
C427 B.n200 VSUBS 0.008898f
C428 B.n201 VSUBS 0.008898f
C429 B.n202 VSUBS 0.008898f
C430 B.n203 VSUBS 0.008898f
C431 B.n204 VSUBS 0.022287f
C432 B.n205 VSUBS 0.023252f
C433 B.n206 VSUBS 0.023252f
C434 B.n207 VSUBS 0.008898f
C435 B.n208 VSUBS 0.008898f
C436 B.n209 VSUBS 0.008898f
C437 B.n210 VSUBS 0.008898f
C438 B.n211 VSUBS 0.008898f
C439 B.n212 VSUBS 0.008898f
C440 B.n213 VSUBS 0.008898f
C441 B.n214 VSUBS 0.008898f
C442 B.n215 VSUBS 0.008898f
C443 B.n216 VSUBS 0.008898f
C444 B.n217 VSUBS 0.008898f
C445 B.n218 VSUBS 0.008898f
C446 B.n219 VSUBS 0.008898f
C447 B.n220 VSUBS 0.008898f
C448 B.n221 VSUBS 0.008898f
C449 B.n222 VSUBS 0.00615f
C450 B.n223 VSUBS 0.020617f
C451 B.n224 VSUBS 0.007197f
C452 B.n225 VSUBS 0.008898f
C453 B.n226 VSUBS 0.008898f
C454 B.n227 VSUBS 0.008898f
C455 B.n228 VSUBS 0.008898f
C456 B.n229 VSUBS 0.008898f
C457 B.n230 VSUBS 0.008898f
C458 B.n231 VSUBS 0.008898f
C459 B.n232 VSUBS 0.008898f
C460 B.n233 VSUBS 0.008898f
C461 B.n234 VSUBS 0.008898f
C462 B.n235 VSUBS 0.008898f
C463 B.t2 VSUBS 0.041034f
C464 B.t1 VSUBS 0.056292f
C465 B.t0 VSUBS 0.36309f
C466 B.n236 VSUBS 0.10558f
C467 B.n237 VSUBS 0.085471f
C468 B.n238 VSUBS 0.020617f
C469 B.n239 VSUBS 0.007197f
C470 B.n240 VSUBS 0.008898f
C471 B.n241 VSUBS 0.008898f
C472 B.n242 VSUBS 0.008898f
C473 B.n243 VSUBS 0.008898f
C474 B.n244 VSUBS 0.008898f
C475 B.n245 VSUBS 0.008898f
C476 B.n246 VSUBS 0.008898f
C477 B.n247 VSUBS 0.008898f
C478 B.n248 VSUBS 0.008898f
C479 B.n249 VSUBS 0.008898f
C480 B.n250 VSUBS 0.008898f
C481 B.n251 VSUBS 0.008898f
C482 B.n252 VSUBS 0.008898f
C483 B.n253 VSUBS 0.008898f
C484 B.n254 VSUBS 0.008898f
C485 B.n255 VSUBS 0.008898f
C486 B.n256 VSUBS 0.008898f
C487 B.n257 VSUBS 0.022332f
C488 B.n258 VSUBS 0.023252f
C489 B.n259 VSUBS 0.022287f
C490 B.n260 VSUBS 0.008898f
C491 B.n261 VSUBS 0.008898f
C492 B.n262 VSUBS 0.008898f
C493 B.n263 VSUBS 0.008898f
C494 B.n264 VSUBS 0.008898f
C495 B.n265 VSUBS 0.008898f
C496 B.n266 VSUBS 0.008898f
C497 B.n267 VSUBS 0.008898f
C498 B.n268 VSUBS 0.008898f
C499 B.n269 VSUBS 0.008898f
C500 B.n270 VSUBS 0.008898f
C501 B.n271 VSUBS 0.008898f
C502 B.n272 VSUBS 0.008898f
C503 B.n273 VSUBS 0.008898f
C504 B.n274 VSUBS 0.008898f
C505 B.n275 VSUBS 0.008898f
C506 B.n276 VSUBS 0.008898f
C507 B.n277 VSUBS 0.008898f
C508 B.n278 VSUBS 0.008898f
C509 B.n279 VSUBS 0.008898f
C510 B.n280 VSUBS 0.008898f
C511 B.n281 VSUBS 0.008898f
C512 B.n282 VSUBS 0.008898f
C513 B.n283 VSUBS 0.008898f
C514 B.n284 VSUBS 0.008898f
C515 B.n285 VSUBS 0.008898f
C516 B.n286 VSUBS 0.008898f
C517 B.n287 VSUBS 0.008898f
C518 B.n288 VSUBS 0.008898f
C519 B.n289 VSUBS 0.008898f
C520 B.n290 VSUBS 0.008898f
C521 B.n291 VSUBS 0.008898f
C522 B.n292 VSUBS 0.008898f
C523 B.n293 VSUBS 0.008898f
C524 B.n294 VSUBS 0.008898f
C525 B.n295 VSUBS 0.008898f
C526 B.n296 VSUBS 0.008898f
C527 B.n297 VSUBS 0.008898f
C528 B.n298 VSUBS 0.008898f
C529 B.n299 VSUBS 0.008898f
C530 B.n300 VSUBS 0.008898f
C531 B.n301 VSUBS 0.008898f
C532 B.n302 VSUBS 0.008898f
C533 B.n303 VSUBS 0.008898f
C534 B.n304 VSUBS 0.008898f
C535 B.n305 VSUBS 0.008898f
C536 B.n306 VSUBS 0.008898f
C537 B.n307 VSUBS 0.008898f
C538 B.n308 VSUBS 0.008898f
C539 B.n309 VSUBS 0.008898f
C540 B.n310 VSUBS 0.008898f
C541 B.n311 VSUBS 0.008898f
C542 B.n312 VSUBS 0.008898f
C543 B.n313 VSUBS 0.008898f
C544 B.n314 VSUBS 0.008898f
C545 B.n315 VSUBS 0.008898f
C546 B.n316 VSUBS 0.008898f
C547 B.n317 VSUBS 0.008898f
C548 B.n318 VSUBS 0.008898f
C549 B.n319 VSUBS 0.008898f
C550 B.n320 VSUBS 0.008898f
C551 B.n321 VSUBS 0.008898f
C552 B.n322 VSUBS 0.008898f
C553 B.n323 VSUBS 0.008898f
C554 B.n324 VSUBS 0.008898f
C555 B.n325 VSUBS 0.008898f
C556 B.n326 VSUBS 0.008898f
C557 B.n327 VSUBS 0.008898f
C558 B.n328 VSUBS 0.008898f
C559 B.n329 VSUBS 0.008898f
C560 B.n330 VSUBS 0.008898f
C561 B.n331 VSUBS 0.008898f
C562 B.n332 VSUBS 0.008898f
C563 B.n333 VSUBS 0.008898f
C564 B.n334 VSUBS 0.008898f
C565 B.n335 VSUBS 0.008898f
C566 B.n336 VSUBS 0.008898f
C567 B.n337 VSUBS 0.008898f
C568 B.n338 VSUBS 0.008898f
C569 B.n339 VSUBS 0.008898f
C570 B.n340 VSUBS 0.008898f
C571 B.n341 VSUBS 0.008898f
C572 B.n342 VSUBS 0.008898f
C573 B.n343 VSUBS 0.008898f
C574 B.n344 VSUBS 0.008898f
C575 B.n345 VSUBS 0.008898f
C576 B.n346 VSUBS 0.008898f
C577 B.n347 VSUBS 0.008898f
C578 B.n348 VSUBS 0.008898f
C579 B.n349 VSUBS 0.008898f
C580 B.n350 VSUBS 0.008898f
C581 B.n351 VSUBS 0.008898f
C582 B.n352 VSUBS 0.008898f
C583 B.n353 VSUBS 0.008898f
C584 B.n354 VSUBS 0.008898f
C585 B.n355 VSUBS 0.008898f
C586 B.n356 VSUBS 0.008898f
C587 B.n357 VSUBS 0.008898f
C588 B.n358 VSUBS 0.008898f
C589 B.n359 VSUBS 0.008898f
C590 B.n360 VSUBS 0.008898f
C591 B.n361 VSUBS 0.008898f
C592 B.n362 VSUBS 0.008898f
C593 B.n363 VSUBS 0.008898f
C594 B.n364 VSUBS 0.008898f
C595 B.n365 VSUBS 0.008898f
C596 B.n366 VSUBS 0.008898f
C597 B.n367 VSUBS 0.008898f
C598 B.n368 VSUBS 0.008898f
C599 B.n369 VSUBS 0.008898f
C600 B.n370 VSUBS 0.008898f
C601 B.n371 VSUBS 0.008898f
C602 B.n372 VSUBS 0.008898f
C603 B.n373 VSUBS 0.008898f
C604 B.n374 VSUBS 0.008898f
C605 B.n375 VSUBS 0.008898f
C606 B.n376 VSUBS 0.008898f
C607 B.n377 VSUBS 0.008898f
C608 B.n378 VSUBS 0.008898f
C609 B.n379 VSUBS 0.008898f
C610 B.n380 VSUBS 0.008898f
C611 B.n381 VSUBS 0.008898f
C612 B.n382 VSUBS 0.008898f
C613 B.n383 VSUBS 0.008898f
C614 B.n384 VSUBS 0.008898f
C615 B.n385 VSUBS 0.008898f
C616 B.n386 VSUBS 0.008898f
C617 B.n387 VSUBS 0.008898f
C618 B.n388 VSUBS 0.008898f
C619 B.n389 VSUBS 0.008898f
C620 B.n390 VSUBS 0.008898f
C621 B.n391 VSUBS 0.008898f
C622 B.n392 VSUBS 0.008898f
C623 B.n393 VSUBS 0.008898f
C624 B.n394 VSUBS 0.008898f
C625 B.n395 VSUBS 0.008898f
C626 B.n396 VSUBS 0.008898f
C627 B.n397 VSUBS 0.008898f
C628 B.n398 VSUBS 0.008898f
C629 B.n399 VSUBS 0.008898f
C630 B.n400 VSUBS 0.008898f
C631 B.n401 VSUBS 0.022287f
C632 B.n402 VSUBS 0.022287f
C633 B.n403 VSUBS 0.023252f
C634 B.n404 VSUBS 0.008898f
C635 B.n405 VSUBS 0.008898f
C636 B.n406 VSUBS 0.008898f
C637 B.n407 VSUBS 0.008898f
C638 B.n408 VSUBS 0.008898f
C639 B.n409 VSUBS 0.008898f
C640 B.n410 VSUBS 0.008898f
C641 B.n411 VSUBS 0.008898f
C642 B.n412 VSUBS 0.008898f
C643 B.n413 VSUBS 0.008898f
C644 B.n414 VSUBS 0.008898f
C645 B.n415 VSUBS 0.008898f
C646 B.n416 VSUBS 0.008898f
C647 B.n417 VSUBS 0.008898f
C648 B.n418 VSUBS 0.008898f
C649 B.n419 VSUBS 0.00615f
C650 B.n420 VSUBS 0.008898f
C651 B.n421 VSUBS 0.008898f
C652 B.n422 VSUBS 0.007197f
C653 B.n423 VSUBS 0.008898f
C654 B.n424 VSUBS 0.008898f
C655 B.n425 VSUBS 0.008898f
C656 B.n426 VSUBS 0.008898f
C657 B.n427 VSUBS 0.008898f
C658 B.n428 VSUBS 0.008898f
C659 B.n429 VSUBS 0.008898f
C660 B.n430 VSUBS 0.008898f
C661 B.n431 VSUBS 0.008898f
C662 B.n432 VSUBS 0.008898f
C663 B.n433 VSUBS 0.008898f
C664 B.n434 VSUBS 0.007197f
C665 B.n435 VSUBS 0.020617f
C666 B.n436 VSUBS 0.00615f
C667 B.n437 VSUBS 0.008898f
C668 B.n438 VSUBS 0.008898f
C669 B.n439 VSUBS 0.008898f
C670 B.n440 VSUBS 0.008898f
C671 B.n441 VSUBS 0.008898f
C672 B.n442 VSUBS 0.008898f
C673 B.n443 VSUBS 0.008898f
C674 B.n444 VSUBS 0.008898f
C675 B.n445 VSUBS 0.008898f
C676 B.n446 VSUBS 0.008898f
C677 B.n447 VSUBS 0.008898f
C678 B.n448 VSUBS 0.008898f
C679 B.n449 VSUBS 0.008898f
C680 B.n450 VSUBS 0.008898f
C681 B.n451 VSUBS 0.008898f
C682 B.n452 VSUBS 0.023252f
C683 B.n453 VSUBS 0.023252f
C684 B.n454 VSUBS 0.022287f
C685 B.n455 VSUBS 0.008898f
C686 B.n456 VSUBS 0.008898f
C687 B.n457 VSUBS 0.008898f
C688 B.n458 VSUBS 0.008898f
C689 B.n459 VSUBS 0.008898f
C690 B.n460 VSUBS 0.008898f
C691 B.n461 VSUBS 0.008898f
C692 B.n462 VSUBS 0.008898f
C693 B.n463 VSUBS 0.008898f
C694 B.n464 VSUBS 0.008898f
C695 B.n465 VSUBS 0.008898f
C696 B.n466 VSUBS 0.008898f
C697 B.n467 VSUBS 0.008898f
C698 B.n468 VSUBS 0.008898f
C699 B.n469 VSUBS 0.008898f
C700 B.n470 VSUBS 0.008898f
C701 B.n471 VSUBS 0.008898f
C702 B.n472 VSUBS 0.008898f
C703 B.n473 VSUBS 0.008898f
C704 B.n474 VSUBS 0.008898f
C705 B.n475 VSUBS 0.008898f
C706 B.n476 VSUBS 0.008898f
C707 B.n477 VSUBS 0.008898f
C708 B.n478 VSUBS 0.008898f
C709 B.n479 VSUBS 0.008898f
C710 B.n480 VSUBS 0.008898f
C711 B.n481 VSUBS 0.008898f
C712 B.n482 VSUBS 0.008898f
C713 B.n483 VSUBS 0.008898f
C714 B.n484 VSUBS 0.008898f
C715 B.n485 VSUBS 0.008898f
C716 B.n486 VSUBS 0.008898f
C717 B.n487 VSUBS 0.008898f
C718 B.n488 VSUBS 0.008898f
C719 B.n489 VSUBS 0.008898f
C720 B.n490 VSUBS 0.008898f
C721 B.n491 VSUBS 0.008898f
C722 B.n492 VSUBS 0.008898f
C723 B.n493 VSUBS 0.008898f
C724 B.n494 VSUBS 0.008898f
C725 B.n495 VSUBS 0.008898f
C726 B.n496 VSUBS 0.008898f
C727 B.n497 VSUBS 0.008898f
C728 B.n498 VSUBS 0.008898f
C729 B.n499 VSUBS 0.008898f
C730 B.n500 VSUBS 0.008898f
C731 B.n501 VSUBS 0.008898f
C732 B.n502 VSUBS 0.008898f
C733 B.n503 VSUBS 0.008898f
C734 B.n504 VSUBS 0.008898f
C735 B.n505 VSUBS 0.008898f
C736 B.n506 VSUBS 0.008898f
C737 B.n507 VSUBS 0.008898f
C738 B.n508 VSUBS 0.008898f
C739 B.n509 VSUBS 0.008898f
C740 B.n510 VSUBS 0.008898f
C741 B.n511 VSUBS 0.008898f
C742 B.n512 VSUBS 0.008898f
C743 B.n513 VSUBS 0.008898f
C744 B.n514 VSUBS 0.008898f
C745 B.n515 VSUBS 0.008898f
C746 B.n516 VSUBS 0.008898f
C747 B.n517 VSUBS 0.008898f
C748 B.n518 VSUBS 0.008898f
C749 B.n519 VSUBS 0.008898f
C750 B.n520 VSUBS 0.008898f
C751 B.n521 VSUBS 0.008898f
C752 B.n522 VSUBS 0.008898f
C753 B.n523 VSUBS 0.011612f
C754 B.n524 VSUBS 0.01237f
C755 B.n525 VSUBS 0.024598f
.ends

