* NGSPICE file created from diff_pair_sample_1441.ext - technology: sky130A

.subckt diff_pair_sample_1441 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=2.4387 pd=15.11 as=2.4387 ps=15.11 w=14.78 l=3.9
X1 VDD1.t6 VP.t1 VTAIL.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=2.4387 pd=15.11 as=5.7642 ps=30.34 w=14.78 l=3.9
X2 VDD2.t7 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.4387 pd=15.11 as=2.4387 ps=15.11 w=14.78 l=3.9
X3 VTAIL.t6 VN.t1 VDD2.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.4387 pd=15.11 as=2.4387 ps=15.11 w=14.78 l=3.9
X4 VDD2.t5 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.4387 pd=15.11 as=5.7642 ps=30.34 w=14.78 l=3.9
X5 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=5.7642 pd=30.34 as=0 ps=0 w=14.78 l=3.9
X6 VDD2.t4 VN.t3 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.4387 pd=15.11 as=2.4387 ps=15.11 w=14.78 l=3.9
X7 VTAIL.t8 VP.t2 VDD1.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=2.4387 pd=15.11 as=2.4387 ps=15.11 w=14.78 l=3.9
X8 VTAIL.t0 VN.t4 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=5.7642 pd=30.34 as=2.4387 ps=15.11 w=14.78 l=3.9
X9 VTAIL.t15 VP.t3 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=5.7642 pd=30.34 as=2.4387 ps=15.11 w=14.78 l=3.9
X10 VDD2.t2 VN.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.4387 pd=15.11 as=5.7642 ps=30.34 w=14.78 l=3.9
X11 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=5.7642 pd=30.34 as=0 ps=0 w=14.78 l=3.9
X12 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=5.7642 pd=30.34 as=0 ps=0 w=14.78 l=3.9
X13 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.7642 pd=30.34 as=0 ps=0 w=14.78 l=3.9
X14 VTAIL.t9 VP.t4 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=2.4387 pd=15.11 as=2.4387 ps=15.11 w=14.78 l=3.9
X15 VDD1.t2 VP.t5 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=2.4387 pd=15.11 as=2.4387 ps=15.11 w=14.78 l=3.9
X16 VDD1.t1 VP.t6 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=2.4387 pd=15.11 as=5.7642 ps=30.34 w=14.78 l=3.9
X17 VTAIL.t4 VN.t6 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.4387 pd=15.11 as=2.4387 ps=15.11 w=14.78 l=3.9
X18 VTAIL.t3 VN.t7 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=5.7642 pd=30.34 as=2.4387 ps=15.11 w=14.78 l=3.9
X19 VTAIL.t14 VP.t7 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.7642 pd=30.34 as=2.4387 ps=15.11 w=14.78 l=3.9
R0 VP.n26 VP.n25 161.3
R1 VP.n27 VP.n22 161.3
R2 VP.n29 VP.n28 161.3
R3 VP.n30 VP.n21 161.3
R4 VP.n32 VP.n31 161.3
R5 VP.n33 VP.n20 161.3
R6 VP.n35 VP.n34 161.3
R7 VP.n36 VP.n19 161.3
R8 VP.n39 VP.n38 161.3
R9 VP.n40 VP.n18 161.3
R10 VP.n42 VP.n41 161.3
R11 VP.n43 VP.n17 161.3
R12 VP.n45 VP.n44 161.3
R13 VP.n46 VP.n16 161.3
R14 VP.n48 VP.n47 161.3
R15 VP.n49 VP.n15 161.3
R16 VP.n51 VP.n50 161.3
R17 VP.n95 VP.n94 161.3
R18 VP.n93 VP.n1 161.3
R19 VP.n92 VP.n91 161.3
R20 VP.n90 VP.n2 161.3
R21 VP.n89 VP.n88 161.3
R22 VP.n87 VP.n3 161.3
R23 VP.n86 VP.n85 161.3
R24 VP.n84 VP.n4 161.3
R25 VP.n83 VP.n82 161.3
R26 VP.n80 VP.n5 161.3
R27 VP.n79 VP.n78 161.3
R28 VP.n77 VP.n6 161.3
R29 VP.n76 VP.n75 161.3
R30 VP.n74 VP.n7 161.3
R31 VP.n73 VP.n72 161.3
R32 VP.n71 VP.n8 161.3
R33 VP.n70 VP.n69 161.3
R34 VP.n67 VP.n9 161.3
R35 VP.n66 VP.n65 161.3
R36 VP.n64 VP.n10 161.3
R37 VP.n63 VP.n62 161.3
R38 VP.n61 VP.n11 161.3
R39 VP.n60 VP.n59 161.3
R40 VP.n58 VP.n12 161.3
R41 VP.n57 VP.n56 161.3
R42 VP.n55 VP.n13 161.3
R43 VP.n23 VP.t3 124.7
R44 VP.n54 VP.t7 91.3333
R45 VP.n68 VP.t5 91.3333
R46 VP.n81 VP.t2 91.3333
R47 VP.n0 VP.t6 91.3333
R48 VP.n14 VP.t1 91.3333
R49 VP.n37 VP.t4 91.3333
R50 VP.n24 VP.t0 91.3333
R51 VP.n54 VP.n53 85.5731
R52 VP.n96 VP.n0 85.5731
R53 VP.n52 VP.n14 85.5731
R54 VP.n53 VP.n52 59.1889
R55 VP.n24 VP.n23 57.3643
R56 VP.n75 VP.n74 56.5617
R57 VP.n31 VP.n30 56.5617
R58 VP.n62 VP.n61 42.5146
R59 VP.n88 VP.n87 42.5146
R60 VP.n44 VP.n43 42.5146
R61 VP.n61 VP.n60 38.6395
R62 VP.n88 VP.n2 38.6395
R63 VP.n44 VP.n16 38.6395
R64 VP.n56 VP.n55 24.5923
R65 VP.n56 VP.n12 24.5923
R66 VP.n60 VP.n12 24.5923
R67 VP.n62 VP.n10 24.5923
R68 VP.n66 VP.n10 24.5923
R69 VP.n67 VP.n66 24.5923
R70 VP.n69 VP.n8 24.5923
R71 VP.n73 VP.n8 24.5923
R72 VP.n74 VP.n73 24.5923
R73 VP.n75 VP.n6 24.5923
R74 VP.n79 VP.n6 24.5923
R75 VP.n80 VP.n79 24.5923
R76 VP.n82 VP.n4 24.5923
R77 VP.n86 VP.n4 24.5923
R78 VP.n87 VP.n86 24.5923
R79 VP.n92 VP.n2 24.5923
R80 VP.n93 VP.n92 24.5923
R81 VP.n94 VP.n93 24.5923
R82 VP.n48 VP.n16 24.5923
R83 VP.n49 VP.n48 24.5923
R84 VP.n50 VP.n49 24.5923
R85 VP.n31 VP.n20 24.5923
R86 VP.n35 VP.n20 24.5923
R87 VP.n36 VP.n35 24.5923
R88 VP.n38 VP.n18 24.5923
R89 VP.n42 VP.n18 24.5923
R90 VP.n43 VP.n42 24.5923
R91 VP.n25 VP.n22 24.5923
R92 VP.n29 VP.n22 24.5923
R93 VP.n30 VP.n29 24.5923
R94 VP.n69 VP.n68 17.9525
R95 VP.n81 VP.n80 17.9525
R96 VP.n37 VP.n36 17.9525
R97 VP.n25 VP.n24 17.9525
R98 VP.n68 VP.n67 6.6403
R99 VP.n82 VP.n81 6.6403
R100 VP.n38 VP.n37 6.6403
R101 VP.n55 VP.n54 4.67295
R102 VP.n94 VP.n0 4.67295
R103 VP.n50 VP.n14 4.67295
R104 VP.n26 VP.n23 2.41404
R105 VP.n52 VP.n51 0.354861
R106 VP.n53 VP.n13 0.354861
R107 VP.n96 VP.n95 0.354861
R108 VP VP.n96 0.267071
R109 VP.n27 VP.n26 0.189894
R110 VP.n28 VP.n27 0.189894
R111 VP.n28 VP.n21 0.189894
R112 VP.n32 VP.n21 0.189894
R113 VP.n33 VP.n32 0.189894
R114 VP.n34 VP.n33 0.189894
R115 VP.n34 VP.n19 0.189894
R116 VP.n39 VP.n19 0.189894
R117 VP.n40 VP.n39 0.189894
R118 VP.n41 VP.n40 0.189894
R119 VP.n41 VP.n17 0.189894
R120 VP.n45 VP.n17 0.189894
R121 VP.n46 VP.n45 0.189894
R122 VP.n47 VP.n46 0.189894
R123 VP.n47 VP.n15 0.189894
R124 VP.n51 VP.n15 0.189894
R125 VP.n57 VP.n13 0.189894
R126 VP.n58 VP.n57 0.189894
R127 VP.n59 VP.n58 0.189894
R128 VP.n59 VP.n11 0.189894
R129 VP.n63 VP.n11 0.189894
R130 VP.n64 VP.n63 0.189894
R131 VP.n65 VP.n64 0.189894
R132 VP.n65 VP.n9 0.189894
R133 VP.n70 VP.n9 0.189894
R134 VP.n71 VP.n70 0.189894
R135 VP.n72 VP.n71 0.189894
R136 VP.n72 VP.n7 0.189894
R137 VP.n76 VP.n7 0.189894
R138 VP.n77 VP.n76 0.189894
R139 VP.n78 VP.n77 0.189894
R140 VP.n78 VP.n5 0.189894
R141 VP.n83 VP.n5 0.189894
R142 VP.n84 VP.n83 0.189894
R143 VP.n85 VP.n84 0.189894
R144 VP.n85 VP.n3 0.189894
R145 VP.n89 VP.n3 0.189894
R146 VP.n90 VP.n89 0.189894
R147 VP.n91 VP.n90 0.189894
R148 VP.n91 VP.n1 0.189894
R149 VP.n95 VP.n1 0.189894
R150 VTAIL.n658 VTAIL.n582 289.615
R151 VTAIL.n78 VTAIL.n2 289.615
R152 VTAIL.n160 VTAIL.n84 289.615
R153 VTAIL.n244 VTAIL.n168 289.615
R154 VTAIL.n576 VTAIL.n500 289.615
R155 VTAIL.n492 VTAIL.n416 289.615
R156 VTAIL.n410 VTAIL.n334 289.615
R157 VTAIL.n326 VTAIL.n250 289.615
R158 VTAIL.n609 VTAIL.n608 185
R159 VTAIL.n606 VTAIL.n605 185
R160 VTAIL.n615 VTAIL.n614 185
R161 VTAIL.n617 VTAIL.n616 185
R162 VTAIL.n602 VTAIL.n601 185
R163 VTAIL.n623 VTAIL.n622 185
R164 VTAIL.n625 VTAIL.n624 185
R165 VTAIL.n598 VTAIL.n597 185
R166 VTAIL.n631 VTAIL.n630 185
R167 VTAIL.n633 VTAIL.n632 185
R168 VTAIL.n594 VTAIL.n593 185
R169 VTAIL.n639 VTAIL.n638 185
R170 VTAIL.n641 VTAIL.n640 185
R171 VTAIL.n590 VTAIL.n589 185
R172 VTAIL.n647 VTAIL.n646 185
R173 VTAIL.n650 VTAIL.n649 185
R174 VTAIL.n648 VTAIL.n586 185
R175 VTAIL.n655 VTAIL.n585 185
R176 VTAIL.n657 VTAIL.n656 185
R177 VTAIL.n659 VTAIL.n658 185
R178 VTAIL.n29 VTAIL.n28 185
R179 VTAIL.n26 VTAIL.n25 185
R180 VTAIL.n35 VTAIL.n34 185
R181 VTAIL.n37 VTAIL.n36 185
R182 VTAIL.n22 VTAIL.n21 185
R183 VTAIL.n43 VTAIL.n42 185
R184 VTAIL.n45 VTAIL.n44 185
R185 VTAIL.n18 VTAIL.n17 185
R186 VTAIL.n51 VTAIL.n50 185
R187 VTAIL.n53 VTAIL.n52 185
R188 VTAIL.n14 VTAIL.n13 185
R189 VTAIL.n59 VTAIL.n58 185
R190 VTAIL.n61 VTAIL.n60 185
R191 VTAIL.n10 VTAIL.n9 185
R192 VTAIL.n67 VTAIL.n66 185
R193 VTAIL.n70 VTAIL.n69 185
R194 VTAIL.n68 VTAIL.n6 185
R195 VTAIL.n75 VTAIL.n5 185
R196 VTAIL.n77 VTAIL.n76 185
R197 VTAIL.n79 VTAIL.n78 185
R198 VTAIL.n111 VTAIL.n110 185
R199 VTAIL.n108 VTAIL.n107 185
R200 VTAIL.n117 VTAIL.n116 185
R201 VTAIL.n119 VTAIL.n118 185
R202 VTAIL.n104 VTAIL.n103 185
R203 VTAIL.n125 VTAIL.n124 185
R204 VTAIL.n127 VTAIL.n126 185
R205 VTAIL.n100 VTAIL.n99 185
R206 VTAIL.n133 VTAIL.n132 185
R207 VTAIL.n135 VTAIL.n134 185
R208 VTAIL.n96 VTAIL.n95 185
R209 VTAIL.n141 VTAIL.n140 185
R210 VTAIL.n143 VTAIL.n142 185
R211 VTAIL.n92 VTAIL.n91 185
R212 VTAIL.n149 VTAIL.n148 185
R213 VTAIL.n152 VTAIL.n151 185
R214 VTAIL.n150 VTAIL.n88 185
R215 VTAIL.n157 VTAIL.n87 185
R216 VTAIL.n159 VTAIL.n158 185
R217 VTAIL.n161 VTAIL.n160 185
R218 VTAIL.n195 VTAIL.n194 185
R219 VTAIL.n192 VTAIL.n191 185
R220 VTAIL.n201 VTAIL.n200 185
R221 VTAIL.n203 VTAIL.n202 185
R222 VTAIL.n188 VTAIL.n187 185
R223 VTAIL.n209 VTAIL.n208 185
R224 VTAIL.n211 VTAIL.n210 185
R225 VTAIL.n184 VTAIL.n183 185
R226 VTAIL.n217 VTAIL.n216 185
R227 VTAIL.n219 VTAIL.n218 185
R228 VTAIL.n180 VTAIL.n179 185
R229 VTAIL.n225 VTAIL.n224 185
R230 VTAIL.n227 VTAIL.n226 185
R231 VTAIL.n176 VTAIL.n175 185
R232 VTAIL.n233 VTAIL.n232 185
R233 VTAIL.n236 VTAIL.n235 185
R234 VTAIL.n234 VTAIL.n172 185
R235 VTAIL.n241 VTAIL.n171 185
R236 VTAIL.n243 VTAIL.n242 185
R237 VTAIL.n245 VTAIL.n244 185
R238 VTAIL.n577 VTAIL.n576 185
R239 VTAIL.n575 VTAIL.n574 185
R240 VTAIL.n573 VTAIL.n503 185
R241 VTAIL.n507 VTAIL.n504 185
R242 VTAIL.n568 VTAIL.n567 185
R243 VTAIL.n566 VTAIL.n565 185
R244 VTAIL.n509 VTAIL.n508 185
R245 VTAIL.n560 VTAIL.n559 185
R246 VTAIL.n558 VTAIL.n557 185
R247 VTAIL.n513 VTAIL.n512 185
R248 VTAIL.n552 VTAIL.n551 185
R249 VTAIL.n550 VTAIL.n549 185
R250 VTAIL.n517 VTAIL.n516 185
R251 VTAIL.n544 VTAIL.n543 185
R252 VTAIL.n542 VTAIL.n541 185
R253 VTAIL.n521 VTAIL.n520 185
R254 VTAIL.n536 VTAIL.n535 185
R255 VTAIL.n534 VTAIL.n533 185
R256 VTAIL.n525 VTAIL.n524 185
R257 VTAIL.n528 VTAIL.n527 185
R258 VTAIL.n493 VTAIL.n492 185
R259 VTAIL.n491 VTAIL.n490 185
R260 VTAIL.n489 VTAIL.n419 185
R261 VTAIL.n423 VTAIL.n420 185
R262 VTAIL.n484 VTAIL.n483 185
R263 VTAIL.n482 VTAIL.n481 185
R264 VTAIL.n425 VTAIL.n424 185
R265 VTAIL.n476 VTAIL.n475 185
R266 VTAIL.n474 VTAIL.n473 185
R267 VTAIL.n429 VTAIL.n428 185
R268 VTAIL.n468 VTAIL.n467 185
R269 VTAIL.n466 VTAIL.n465 185
R270 VTAIL.n433 VTAIL.n432 185
R271 VTAIL.n460 VTAIL.n459 185
R272 VTAIL.n458 VTAIL.n457 185
R273 VTAIL.n437 VTAIL.n436 185
R274 VTAIL.n452 VTAIL.n451 185
R275 VTAIL.n450 VTAIL.n449 185
R276 VTAIL.n441 VTAIL.n440 185
R277 VTAIL.n444 VTAIL.n443 185
R278 VTAIL.n411 VTAIL.n410 185
R279 VTAIL.n409 VTAIL.n408 185
R280 VTAIL.n407 VTAIL.n337 185
R281 VTAIL.n341 VTAIL.n338 185
R282 VTAIL.n402 VTAIL.n401 185
R283 VTAIL.n400 VTAIL.n399 185
R284 VTAIL.n343 VTAIL.n342 185
R285 VTAIL.n394 VTAIL.n393 185
R286 VTAIL.n392 VTAIL.n391 185
R287 VTAIL.n347 VTAIL.n346 185
R288 VTAIL.n386 VTAIL.n385 185
R289 VTAIL.n384 VTAIL.n383 185
R290 VTAIL.n351 VTAIL.n350 185
R291 VTAIL.n378 VTAIL.n377 185
R292 VTAIL.n376 VTAIL.n375 185
R293 VTAIL.n355 VTAIL.n354 185
R294 VTAIL.n370 VTAIL.n369 185
R295 VTAIL.n368 VTAIL.n367 185
R296 VTAIL.n359 VTAIL.n358 185
R297 VTAIL.n362 VTAIL.n361 185
R298 VTAIL.n327 VTAIL.n326 185
R299 VTAIL.n325 VTAIL.n324 185
R300 VTAIL.n323 VTAIL.n253 185
R301 VTAIL.n257 VTAIL.n254 185
R302 VTAIL.n318 VTAIL.n317 185
R303 VTAIL.n316 VTAIL.n315 185
R304 VTAIL.n259 VTAIL.n258 185
R305 VTAIL.n310 VTAIL.n309 185
R306 VTAIL.n308 VTAIL.n307 185
R307 VTAIL.n263 VTAIL.n262 185
R308 VTAIL.n302 VTAIL.n301 185
R309 VTAIL.n300 VTAIL.n299 185
R310 VTAIL.n267 VTAIL.n266 185
R311 VTAIL.n294 VTAIL.n293 185
R312 VTAIL.n292 VTAIL.n291 185
R313 VTAIL.n271 VTAIL.n270 185
R314 VTAIL.n286 VTAIL.n285 185
R315 VTAIL.n284 VTAIL.n283 185
R316 VTAIL.n275 VTAIL.n274 185
R317 VTAIL.n278 VTAIL.n277 185
R318 VTAIL.t12 VTAIL.n526 147.659
R319 VTAIL.t15 VTAIL.n442 147.659
R320 VTAIL.t5 VTAIL.n360 147.659
R321 VTAIL.t0 VTAIL.n276 147.659
R322 VTAIL.t1 VTAIL.n607 147.659
R323 VTAIL.t3 VTAIL.n27 147.659
R324 VTAIL.t13 VTAIL.n109 147.659
R325 VTAIL.t14 VTAIL.n193 147.659
R326 VTAIL.n608 VTAIL.n605 104.615
R327 VTAIL.n615 VTAIL.n605 104.615
R328 VTAIL.n616 VTAIL.n615 104.615
R329 VTAIL.n616 VTAIL.n601 104.615
R330 VTAIL.n623 VTAIL.n601 104.615
R331 VTAIL.n624 VTAIL.n623 104.615
R332 VTAIL.n624 VTAIL.n597 104.615
R333 VTAIL.n631 VTAIL.n597 104.615
R334 VTAIL.n632 VTAIL.n631 104.615
R335 VTAIL.n632 VTAIL.n593 104.615
R336 VTAIL.n639 VTAIL.n593 104.615
R337 VTAIL.n640 VTAIL.n639 104.615
R338 VTAIL.n640 VTAIL.n589 104.615
R339 VTAIL.n647 VTAIL.n589 104.615
R340 VTAIL.n649 VTAIL.n647 104.615
R341 VTAIL.n649 VTAIL.n648 104.615
R342 VTAIL.n648 VTAIL.n585 104.615
R343 VTAIL.n657 VTAIL.n585 104.615
R344 VTAIL.n658 VTAIL.n657 104.615
R345 VTAIL.n28 VTAIL.n25 104.615
R346 VTAIL.n35 VTAIL.n25 104.615
R347 VTAIL.n36 VTAIL.n35 104.615
R348 VTAIL.n36 VTAIL.n21 104.615
R349 VTAIL.n43 VTAIL.n21 104.615
R350 VTAIL.n44 VTAIL.n43 104.615
R351 VTAIL.n44 VTAIL.n17 104.615
R352 VTAIL.n51 VTAIL.n17 104.615
R353 VTAIL.n52 VTAIL.n51 104.615
R354 VTAIL.n52 VTAIL.n13 104.615
R355 VTAIL.n59 VTAIL.n13 104.615
R356 VTAIL.n60 VTAIL.n59 104.615
R357 VTAIL.n60 VTAIL.n9 104.615
R358 VTAIL.n67 VTAIL.n9 104.615
R359 VTAIL.n69 VTAIL.n67 104.615
R360 VTAIL.n69 VTAIL.n68 104.615
R361 VTAIL.n68 VTAIL.n5 104.615
R362 VTAIL.n77 VTAIL.n5 104.615
R363 VTAIL.n78 VTAIL.n77 104.615
R364 VTAIL.n110 VTAIL.n107 104.615
R365 VTAIL.n117 VTAIL.n107 104.615
R366 VTAIL.n118 VTAIL.n117 104.615
R367 VTAIL.n118 VTAIL.n103 104.615
R368 VTAIL.n125 VTAIL.n103 104.615
R369 VTAIL.n126 VTAIL.n125 104.615
R370 VTAIL.n126 VTAIL.n99 104.615
R371 VTAIL.n133 VTAIL.n99 104.615
R372 VTAIL.n134 VTAIL.n133 104.615
R373 VTAIL.n134 VTAIL.n95 104.615
R374 VTAIL.n141 VTAIL.n95 104.615
R375 VTAIL.n142 VTAIL.n141 104.615
R376 VTAIL.n142 VTAIL.n91 104.615
R377 VTAIL.n149 VTAIL.n91 104.615
R378 VTAIL.n151 VTAIL.n149 104.615
R379 VTAIL.n151 VTAIL.n150 104.615
R380 VTAIL.n150 VTAIL.n87 104.615
R381 VTAIL.n159 VTAIL.n87 104.615
R382 VTAIL.n160 VTAIL.n159 104.615
R383 VTAIL.n194 VTAIL.n191 104.615
R384 VTAIL.n201 VTAIL.n191 104.615
R385 VTAIL.n202 VTAIL.n201 104.615
R386 VTAIL.n202 VTAIL.n187 104.615
R387 VTAIL.n209 VTAIL.n187 104.615
R388 VTAIL.n210 VTAIL.n209 104.615
R389 VTAIL.n210 VTAIL.n183 104.615
R390 VTAIL.n217 VTAIL.n183 104.615
R391 VTAIL.n218 VTAIL.n217 104.615
R392 VTAIL.n218 VTAIL.n179 104.615
R393 VTAIL.n225 VTAIL.n179 104.615
R394 VTAIL.n226 VTAIL.n225 104.615
R395 VTAIL.n226 VTAIL.n175 104.615
R396 VTAIL.n233 VTAIL.n175 104.615
R397 VTAIL.n235 VTAIL.n233 104.615
R398 VTAIL.n235 VTAIL.n234 104.615
R399 VTAIL.n234 VTAIL.n171 104.615
R400 VTAIL.n243 VTAIL.n171 104.615
R401 VTAIL.n244 VTAIL.n243 104.615
R402 VTAIL.n576 VTAIL.n575 104.615
R403 VTAIL.n575 VTAIL.n503 104.615
R404 VTAIL.n507 VTAIL.n503 104.615
R405 VTAIL.n567 VTAIL.n507 104.615
R406 VTAIL.n567 VTAIL.n566 104.615
R407 VTAIL.n566 VTAIL.n508 104.615
R408 VTAIL.n559 VTAIL.n508 104.615
R409 VTAIL.n559 VTAIL.n558 104.615
R410 VTAIL.n558 VTAIL.n512 104.615
R411 VTAIL.n551 VTAIL.n512 104.615
R412 VTAIL.n551 VTAIL.n550 104.615
R413 VTAIL.n550 VTAIL.n516 104.615
R414 VTAIL.n543 VTAIL.n516 104.615
R415 VTAIL.n543 VTAIL.n542 104.615
R416 VTAIL.n542 VTAIL.n520 104.615
R417 VTAIL.n535 VTAIL.n520 104.615
R418 VTAIL.n535 VTAIL.n534 104.615
R419 VTAIL.n534 VTAIL.n524 104.615
R420 VTAIL.n527 VTAIL.n524 104.615
R421 VTAIL.n492 VTAIL.n491 104.615
R422 VTAIL.n491 VTAIL.n419 104.615
R423 VTAIL.n423 VTAIL.n419 104.615
R424 VTAIL.n483 VTAIL.n423 104.615
R425 VTAIL.n483 VTAIL.n482 104.615
R426 VTAIL.n482 VTAIL.n424 104.615
R427 VTAIL.n475 VTAIL.n424 104.615
R428 VTAIL.n475 VTAIL.n474 104.615
R429 VTAIL.n474 VTAIL.n428 104.615
R430 VTAIL.n467 VTAIL.n428 104.615
R431 VTAIL.n467 VTAIL.n466 104.615
R432 VTAIL.n466 VTAIL.n432 104.615
R433 VTAIL.n459 VTAIL.n432 104.615
R434 VTAIL.n459 VTAIL.n458 104.615
R435 VTAIL.n458 VTAIL.n436 104.615
R436 VTAIL.n451 VTAIL.n436 104.615
R437 VTAIL.n451 VTAIL.n450 104.615
R438 VTAIL.n450 VTAIL.n440 104.615
R439 VTAIL.n443 VTAIL.n440 104.615
R440 VTAIL.n410 VTAIL.n409 104.615
R441 VTAIL.n409 VTAIL.n337 104.615
R442 VTAIL.n341 VTAIL.n337 104.615
R443 VTAIL.n401 VTAIL.n341 104.615
R444 VTAIL.n401 VTAIL.n400 104.615
R445 VTAIL.n400 VTAIL.n342 104.615
R446 VTAIL.n393 VTAIL.n342 104.615
R447 VTAIL.n393 VTAIL.n392 104.615
R448 VTAIL.n392 VTAIL.n346 104.615
R449 VTAIL.n385 VTAIL.n346 104.615
R450 VTAIL.n385 VTAIL.n384 104.615
R451 VTAIL.n384 VTAIL.n350 104.615
R452 VTAIL.n377 VTAIL.n350 104.615
R453 VTAIL.n377 VTAIL.n376 104.615
R454 VTAIL.n376 VTAIL.n354 104.615
R455 VTAIL.n369 VTAIL.n354 104.615
R456 VTAIL.n369 VTAIL.n368 104.615
R457 VTAIL.n368 VTAIL.n358 104.615
R458 VTAIL.n361 VTAIL.n358 104.615
R459 VTAIL.n326 VTAIL.n325 104.615
R460 VTAIL.n325 VTAIL.n253 104.615
R461 VTAIL.n257 VTAIL.n253 104.615
R462 VTAIL.n317 VTAIL.n257 104.615
R463 VTAIL.n317 VTAIL.n316 104.615
R464 VTAIL.n316 VTAIL.n258 104.615
R465 VTAIL.n309 VTAIL.n258 104.615
R466 VTAIL.n309 VTAIL.n308 104.615
R467 VTAIL.n308 VTAIL.n262 104.615
R468 VTAIL.n301 VTAIL.n262 104.615
R469 VTAIL.n301 VTAIL.n300 104.615
R470 VTAIL.n300 VTAIL.n266 104.615
R471 VTAIL.n293 VTAIL.n266 104.615
R472 VTAIL.n293 VTAIL.n292 104.615
R473 VTAIL.n292 VTAIL.n270 104.615
R474 VTAIL.n285 VTAIL.n270 104.615
R475 VTAIL.n285 VTAIL.n284 104.615
R476 VTAIL.n284 VTAIL.n274 104.615
R477 VTAIL.n277 VTAIL.n274 104.615
R478 VTAIL.n608 VTAIL.t1 52.3082
R479 VTAIL.n28 VTAIL.t3 52.3082
R480 VTAIL.n110 VTAIL.t13 52.3082
R481 VTAIL.n194 VTAIL.t14 52.3082
R482 VTAIL.n527 VTAIL.t12 52.3082
R483 VTAIL.n443 VTAIL.t15 52.3082
R484 VTAIL.n361 VTAIL.t5 52.3082
R485 VTAIL.n277 VTAIL.t0 52.3082
R486 VTAIL.n499 VTAIL.n498 46.9575
R487 VTAIL.n333 VTAIL.n332 46.9575
R488 VTAIL.n1 VTAIL.n0 46.9573
R489 VTAIL.n167 VTAIL.n166 46.9573
R490 VTAIL.n663 VTAIL.n662 34.9005
R491 VTAIL.n83 VTAIL.n82 34.9005
R492 VTAIL.n165 VTAIL.n164 34.9005
R493 VTAIL.n249 VTAIL.n248 34.9005
R494 VTAIL.n581 VTAIL.n580 34.9005
R495 VTAIL.n497 VTAIL.n496 34.9005
R496 VTAIL.n415 VTAIL.n414 34.9005
R497 VTAIL.n331 VTAIL.n330 34.9005
R498 VTAIL.n663 VTAIL.n581 28.7548
R499 VTAIL.n331 VTAIL.n249 28.7548
R500 VTAIL.n609 VTAIL.n607 15.6677
R501 VTAIL.n29 VTAIL.n27 15.6677
R502 VTAIL.n111 VTAIL.n109 15.6677
R503 VTAIL.n195 VTAIL.n193 15.6677
R504 VTAIL.n528 VTAIL.n526 15.6677
R505 VTAIL.n444 VTAIL.n442 15.6677
R506 VTAIL.n362 VTAIL.n360 15.6677
R507 VTAIL.n278 VTAIL.n276 15.6677
R508 VTAIL.n656 VTAIL.n655 13.1884
R509 VTAIL.n76 VTAIL.n75 13.1884
R510 VTAIL.n158 VTAIL.n157 13.1884
R511 VTAIL.n242 VTAIL.n241 13.1884
R512 VTAIL.n574 VTAIL.n573 13.1884
R513 VTAIL.n490 VTAIL.n489 13.1884
R514 VTAIL.n408 VTAIL.n407 13.1884
R515 VTAIL.n324 VTAIL.n323 13.1884
R516 VTAIL.n610 VTAIL.n606 12.8005
R517 VTAIL.n654 VTAIL.n586 12.8005
R518 VTAIL.n659 VTAIL.n584 12.8005
R519 VTAIL.n30 VTAIL.n26 12.8005
R520 VTAIL.n74 VTAIL.n6 12.8005
R521 VTAIL.n79 VTAIL.n4 12.8005
R522 VTAIL.n112 VTAIL.n108 12.8005
R523 VTAIL.n156 VTAIL.n88 12.8005
R524 VTAIL.n161 VTAIL.n86 12.8005
R525 VTAIL.n196 VTAIL.n192 12.8005
R526 VTAIL.n240 VTAIL.n172 12.8005
R527 VTAIL.n245 VTAIL.n170 12.8005
R528 VTAIL.n577 VTAIL.n502 12.8005
R529 VTAIL.n572 VTAIL.n504 12.8005
R530 VTAIL.n529 VTAIL.n525 12.8005
R531 VTAIL.n493 VTAIL.n418 12.8005
R532 VTAIL.n488 VTAIL.n420 12.8005
R533 VTAIL.n445 VTAIL.n441 12.8005
R534 VTAIL.n411 VTAIL.n336 12.8005
R535 VTAIL.n406 VTAIL.n338 12.8005
R536 VTAIL.n363 VTAIL.n359 12.8005
R537 VTAIL.n327 VTAIL.n252 12.8005
R538 VTAIL.n322 VTAIL.n254 12.8005
R539 VTAIL.n279 VTAIL.n275 12.8005
R540 VTAIL.n614 VTAIL.n613 12.0247
R541 VTAIL.n651 VTAIL.n650 12.0247
R542 VTAIL.n660 VTAIL.n582 12.0247
R543 VTAIL.n34 VTAIL.n33 12.0247
R544 VTAIL.n71 VTAIL.n70 12.0247
R545 VTAIL.n80 VTAIL.n2 12.0247
R546 VTAIL.n116 VTAIL.n115 12.0247
R547 VTAIL.n153 VTAIL.n152 12.0247
R548 VTAIL.n162 VTAIL.n84 12.0247
R549 VTAIL.n200 VTAIL.n199 12.0247
R550 VTAIL.n237 VTAIL.n236 12.0247
R551 VTAIL.n246 VTAIL.n168 12.0247
R552 VTAIL.n578 VTAIL.n500 12.0247
R553 VTAIL.n569 VTAIL.n568 12.0247
R554 VTAIL.n533 VTAIL.n532 12.0247
R555 VTAIL.n494 VTAIL.n416 12.0247
R556 VTAIL.n485 VTAIL.n484 12.0247
R557 VTAIL.n449 VTAIL.n448 12.0247
R558 VTAIL.n412 VTAIL.n334 12.0247
R559 VTAIL.n403 VTAIL.n402 12.0247
R560 VTAIL.n367 VTAIL.n366 12.0247
R561 VTAIL.n328 VTAIL.n250 12.0247
R562 VTAIL.n319 VTAIL.n318 12.0247
R563 VTAIL.n283 VTAIL.n282 12.0247
R564 VTAIL.n617 VTAIL.n604 11.249
R565 VTAIL.n646 VTAIL.n588 11.249
R566 VTAIL.n37 VTAIL.n24 11.249
R567 VTAIL.n66 VTAIL.n8 11.249
R568 VTAIL.n119 VTAIL.n106 11.249
R569 VTAIL.n148 VTAIL.n90 11.249
R570 VTAIL.n203 VTAIL.n190 11.249
R571 VTAIL.n232 VTAIL.n174 11.249
R572 VTAIL.n565 VTAIL.n506 11.249
R573 VTAIL.n536 VTAIL.n523 11.249
R574 VTAIL.n481 VTAIL.n422 11.249
R575 VTAIL.n452 VTAIL.n439 11.249
R576 VTAIL.n399 VTAIL.n340 11.249
R577 VTAIL.n370 VTAIL.n357 11.249
R578 VTAIL.n315 VTAIL.n256 11.249
R579 VTAIL.n286 VTAIL.n273 11.249
R580 VTAIL.n618 VTAIL.n602 10.4732
R581 VTAIL.n645 VTAIL.n590 10.4732
R582 VTAIL.n38 VTAIL.n22 10.4732
R583 VTAIL.n65 VTAIL.n10 10.4732
R584 VTAIL.n120 VTAIL.n104 10.4732
R585 VTAIL.n147 VTAIL.n92 10.4732
R586 VTAIL.n204 VTAIL.n188 10.4732
R587 VTAIL.n231 VTAIL.n176 10.4732
R588 VTAIL.n564 VTAIL.n509 10.4732
R589 VTAIL.n537 VTAIL.n521 10.4732
R590 VTAIL.n480 VTAIL.n425 10.4732
R591 VTAIL.n453 VTAIL.n437 10.4732
R592 VTAIL.n398 VTAIL.n343 10.4732
R593 VTAIL.n371 VTAIL.n355 10.4732
R594 VTAIL.n314 VTAIL.n259 10.4732
R595 VTAIL.n287 VTAIL.n271 10.4732
R596 VTAIL.n622 VTAIL.n621 9.69747
R597 VTAIL.n642 VTAIL.n641 9.69747
R598 VTAIL.n42 VTAIL.n41 9.69747
R599 VTAIL.n62 VTAIL.n61 9.69747
R600 VTAIL.n124 VTAIL.n123 9.69747
R601 VTAIL.n144 VTAIL.n143 9.69747
R602 VTAIL.n208 VTAIL.n207 9.69747
R603 VTAIL.n228 VTAIL.n227 9.69747
R604 VTAIL.n561 VTAIL.n560 9.69747
R605 VTAIL.n541 VTAIL.n540 9.69747
R606 VTAIL.n477 VTAIL.n476 9.69747
R607 VTAIL.n457 VTAIL.n456 9.69747
R608 VTAIL.n395 VTAIL.n394 9.69747
R609 VTAIL.n375 VTAIL.n374 9.69747
R610 VTAIL.n311 VTAIL.n310 9.69747
R611 VTAIL.n291 VTAIL.n290 9.69747
R612 VTAIL.n662 VTAIL.n661 9.45567
R613 VTAIL.n82 VTAIL.n81 9.45567
R614 VTAIL.n164 VTAIL.n163 9.45567
R615 VTAIL.n248 VTAIL.n247 9.45567
R616 VTAIL.n580 VTAIL.n579 9.45567
R617 VTAIL.n496 VTAIL.n495 9.45567
R618 VTAIL.n414 VTAIL.n413 9.45567
R619 VTAIL.n330 VTAIL.n329 9.45567
R620 VTAIL.n661 VTAIL.n660 9.3005
R621 VTAIL.n584 VTAIL.n583 9.3005
R622 VTAIL.n629 VTAIL.n628 9.3005
R623 VTAIL.n627 VTAIL.n626 9.3005
R624 VTAIL.n600 VTAIL.n599 9.3005
R625 VTAIL.n621 VTAIL.n620 9.3005
R626 VTAIL.n619 VTAIL.n618 9.3005
R627 VTAIL.n604 VTAIL.n603 9.3005
R628 VTAIL.n613 VTAIL.n612 9.3005
R629 VTAIL.n611 VTAIL.n610 9.3005
R630 VTAIL.n596 VTAIL.n595 9.3005
R631 VTAIL.n635 VTAIL.n634 9.3005
R632 VTAIL.n637 VTAIL.n636 9.3005
R633 VTAIL.n592 VTAIL.n591 9.3005
R634 VTAIL.n643 VTAIL.n642 9.3005
R635 VTAIL.n645 VTAIL.n644 9.3005
R636 VTAIL.n588 VTAIL.n587 9.3005
R637 VTAIL.n652 VTAIL.n651 9.3005
R638 VTAIL.n654 VTAIL.n653 9.3005
R639 VTAIL.n81 VTAIL.n80 9.3005
R640 VTAIL.n4 VTAIL.n3 9.3005
R641 VTAIL.n49 VTAIL.n48 9.3005
R642 VTAIL.n47 VTAIL.n46 9.3005
R643 VTAIL.n20 VTAIL.n19 9.3005
R644 VTAIL.n41 VTAIL.n40 9.3005
R645 VTAIL.n39 VTAIL.n38 9.3005
R646 VTAIL.n24 VTAIL.n23 9.3005
R647 VTAIL.n33 VTAIL.n32 9.3005
R648 VTAIL.n31 VTAIL.n30 9.3005
R649 VTAIL.n16 VTAIL.n15 9.3005
R650 VTAIL.n55 VTAIL.n54 9.3005
R651 VTAIL.n57 VTAIL.n56 9.3005
R652 VTAIL.n12 VTAIL.n11 9.3005
R653 VTAIL.n63 VTAIL.n62 9.3005
R654 VTAIL.n65 VTAIL.n64 9.3005
R655 VTAIL.n8 VTAIL.n7 9.3005
R656 VTAIL.n72 VTAIL.n71 9.3005
R657 VTAIL.n74 VTAIL.n73 9.3005
R658 VTAIL.n163 VTAIL.n162 9.3005
R659 VTAIL.n86 VTAIL.n85 9.3005
R660 VTAIL.n131 VTAIL.n130 9.3005
R661 VTAIL.n129 VTAIL.n128 9.3005
R662 VTAIL.n102 VTAIL.n101 9.3005
R663 VTAIL.n123 VTAIL.n122 9.3005
R664 VTAIL.n121 VTAIL.n120 9.3005
R665 VTAIL.n106 VTAIL.n105 9.3005
R666 VTAIL.n115 VTAIL.n114 9.3005
R667 VTAIL.n113 VTAIL.n112 9.3005
R668 VTAIL.n98 VTAIL.n97 9.3005
R669 VTAIL.n137 VTAIL.n136 9.3005
R670 VTAIL.n139 VTAIL.n138 9.3005
R671 VTAIL.n94 VTAIL.n93 9.3005
R672 VTAIL.n145 VTAIL.n144 9.3005
R673 VTAIL.n147 VTAIL.n146 9.3005
R674 VTAIL.n90 VTAIL.n89 9.3005
R675 VTAIL.n154 VTAIL.n153 9.3005
R676 VTAIL.n156 VTAIL.n155 9.3005
R677 VTAIL.n247 VTAIL.n246 9.3005
R678 VTAIL.n170 VTAIL.n169 9.3005
R679 VTAIL.n215 VTAIL.n214 9.3005
R680 VTAIL.n213 VTAIL.n212 9.3005
R681 VTAIL.n186 VTAIL.n185 9.3005
R682 VTAIL.n207 VTAIL.n206 9.3005
R683 VTAIL.n205 VTAIL.n204 9.3005
R684 VTAIL.n190 VTAIL.n189 9.3005
R685 VTAIL.n199 VTAIL.n198 9.3005
R686 VTAIL.n197 VTAIL.n196 9.3005
R687 VTAIL.n182 VTAIL.n181 9.3005
R688 VTAIL.n221 VTAIL.n220 9.3005
R689 VTAIL.n223 VTAIL.n222 9.3005
R690 VTAIL.n178 VTAIL.n177 9.3005
R691 VTAIL.n229 VTAIL.n228 9.3005
R692 VTAIL.n231 VTAIL.n230 9.3005
R693 VTAIL.n174 VTAIL.n173 9.3005
R694 VTAIL.n238 VTAIL.n237 9.3005
R695 VTAIL.n240 VTAIL.n239 9.3005
R696 VTAIL.n554 VTAIL.n553 9.3005
R697 VTAIL.n556 VTAIL.n555 9.3005
R698 VTAIL.n511 VTAIL.n510 9.3005
R699 VTAIL.n562 VTAIL.n561 9.3005
R700 VTAIL.n564 VTAIL.n563 9.3005
R701 VTAIL.n506 VTAIL.n505 9.3005
R702 VTAIL.n570 VTAIL.n569 9.3005
R703 VTAIL.n572 VTAIL.n571 9.3005
R704 VTAIL.n579 VTAIL.n578 9.3005
R705 VTAIL.n502 VTAIL.n501 9.3005
R706 VTAIL.n515 VTAIL.n514 9.3005
R707 VTAIL.n548 VTAIL.n547 9.3005
R708 VTAIL.n546 VTAIL.n545 9.3005
R709 VTAIL.n519 VTAIL.n518 9.3005
R710 VTAIL.n540 VTAIL.n539 9.3005
R711 VTAIL.n538 VTAIL.n537 9.3005
R712 VTAIL.n523 VTAIL.n522 9.3005
R713 VTAIL.n532 VTAIL.n531 9.3005
R714 VTAIL.n530 VTAIL.n529 9.3005
R715 VTAIL.n470 VTAIL.n469 9.3005
R716 VTAIL.n472 VTAIL.n471 9.3005
R717 VTAIL.n427 VTAIL.n426 9.3005
R718 VTAIL.n478 VTAIL.n477 9.3005
R719 VTAIL.n480 VTAIL.n479 9.3005
R720 VTAIL.n422 VTAIL.n421 9.3005
R721 VTAIL.n486 VTAIL.n485 9.3005
R722 VTAIL.n488 VTAIL.n487 9.3005
R723 VTAIL.n495 VTAIL.n494 9.3005
R724 VTAIL.n418 VTAIL.n417 9.3005
R725 VTAIL.n431 VTAIL.n430 9.3005
R726 VTAIL.n464 VTAIL.n463 9.3005
R727 VTAIL.n462 VTAIL.n461 9.3005
R728 VTAIL.n435 VTAIL.n434 9.3005
R729 VTAIL.n456 VTAIL.n455 9.3005
R730 VTAIL.n454 VTAIL.n453 9.3005
R731 VTAIL.n439 VTAIL.n438 9.3005
R732 VTAIL.n448 VTAIL.n447 9.3005
R733 VTAIL.n446 VTAIL.n445 9.3005
R734 VTAIL.n388 VTAIL.n387 9.3005
R735 VTAIL.n390 VTAIL.n389 9.3005
R736 VTAIL.n345 VTAIL.n344 9.3005
R737 VTAIL.n396 VTAIL.n395 9.3005
R738 VTAIL.n398 VTAIL.n397 9.3005
R739 VTAIL.n340 VTAIL.n339 9.3005
R740 VTAIL.n404 VTAIL.n403 9.3005
R741 VTAIL.n406 VTAIL.n405 9.3005
R742 VTAIL.n413 VTAIL.n412 9.3005
R743 VTAIL.n336 VTAIL.n335 9.3005
R744 VTAIL.n349 VTAIL.n348 9.3005
R745 VTAIL.n382 VTAIL.n381 9.3005
R746 VTAIL.n380 VTAIL.n379 9.3005
R747 VTAIL.n353 VTAIL.n352 9.3005
R748 VTAIL.n374 VTAIL.n373 9.3005
R749 VTAIL.n372 VTAIL.n371 9.3005
R750 VTAIL.n357 VTAIL.n356 9.3005
R751 VTAIL.n366 VTAIL.n365 9.3005
R752 VTAIL.n364 VTAIL.n363 9.3005
R753 VTAIL.n304 VTAIL.n303 9.3005
R754 VTAIL.n306 VTAIL.n305 9.3005
R755 VTAIL.n261 VTAIL.n260 9.3005
R756 VTAIL.n312 VTAIL.n311 9.3005
R757 VTAIL.n314 VTAIL.n313 9.3005
R758 VTAIL.n256 VTAIL.n255 9.3005
R759 VTAIL.n320 VTAIL.n319 9.3005
R760 VTAIL.n322 VTAIL.n321 9.3005
R761 VTAIL.n329 VTAIL.n328 9.3005
R762 VTAIL.n252 VTAIL.n251 9.3005
R763 VTAIL.n265 VTAIL.n264 9.3005
R764 VTAIL.n298 VTAIL.n297 9.3005
R765 VTAIL.n296 VTAIL.n295 9.3005
R766 VTAIL.n269 VTAIL.n268 9.3005
R767 VTAIL.n290 VTAIL.n289 9.3005
R768 VTAIL.n288 VTAIL.n287 9.3005
R769 VTAIL.n273 VTAIL.n272 9.3005
R770 VTAIL.n282 VTAIL.n281 9.3005
R771 VTAIL.n280 VTAIL.n279 9.3005
R772 VTAIL.n625 VTAIL.n600 8.92171
R773 VTAIL.n638 VTAIL.n592 8.92171
R774 VTAIL.n45 VTAIL.n20 8.92171
R775 VTAIL.n58 VTAIL.n12 8.92171
R776 VTAIL.n127 VTAIL.n102 8.92171
R777 VTAIL.n140 VTAIL.n94 8.92171
R778 VTAIL.n211 VTAIL.n186 8.92171
R779 VTAIL.n224 VTAIL.n178 8.92171
R780 VTAIL.n557 VTAIL.n511 8.92171
R781 VTAIL.n544 VTAIL.n519 8.92171
R782 VTAIL.n473 VTAIL.n427 8.92171
R783 VTAIL.n460 VTAIL.n435 8.92171
R784 VTAIL.n391 VTAIL.n345 8.92171
R785 VTAIL.n378 VTAIL.n353 8.92171
R786 VTAIL.n307 VTAIL.n261 8.92171
R787 VTAIL.n294 VTAIL.n269 8.92171
R788 VTAIL.n626 VTAIL.n598 8.14595
R789 VTAIL.n637 VTAIL.n594 8.14595
R790 VTAIL.n46 VTAIL.n18 8.14595
R791 VTAIL.n57 VTAIL.n14 8.14595
R792 VTAIL.n128 VTAIL.n100 8.14595
R793 VTAIL.n139 VTAIL.n96 8.14595
R794 VTAIL.n212 VTAIL.n184 8.14595
R795 VTAIL.n223 VTAIL.n180 8.14595
R796 VTAIL.n556 VTAIL.n513 8.14595
R797 VTAIL.n545 VTAIL.n517 8.14595
R798 VTAIL.n472 VTAIL.n429 8.14595
R799 VTAIL.n461 VTAIL.n433 8.14595
R800 VTAIL.n390 VTAIL.n347 8.14595
R801 VTAIL.n379 VTAIL.n351 8.14595
R802 VTAIL.n306 VTAIL.n263 8.14595
R803 VTAIL.n295 VTAIL.n267 8.14595
R804 VTAIL.n630 VTAIL.n629 7.3702
R805 VTAIL.n634 VTAIL.n633 7.3702
R806 VTAIL.n50 VTAIL.n49 7.3702
R807 VTAIL.n54 VTAIL.n53 7.3702
R808 VTAIL.n132 VTAIL.n131 7.3702
R809 VTAIL.n136 VTAIL.n135 7.3702
R810 VTAIL.n216 VTAIL.n215 7.3702
R811 VTAIL.n220 VTAIL.n219 7.3702
R812 VTAIL.n553 VTAIL.n552 7.3702
R813 VTAIL.n549 VTAIL.n548 7.3702
R814 VTAIL.n469 VTAIL.n468 7.3702
R815 VTAIL.n465 VTAIL.n464 7.3702
R816 VTAIL.n387 VTAIL.n386 7.3702
R817 VTAIL.n383 VTAIL.n382 7.3702
R818 VTAIL.n303 VTAIL.n302 7.3702
R819 VTAIL.n299 VTAIL.n298 7.3702
R820 VTAIL.n630 VTAIL.n596 6.59444
R821 VTAIL.n633 VTAIL.n596 6.59444
R822 VTAIL.n50 VTAIL.n16 6.59444
R823 VTAIL.n53 VTAIL.n16 6.59444
R824 VTAIL.n132 VTAIL.n98 6.59444
R825 VTAIL.n135 VTAIL.n98 6.59444
R826 VTAIL.n216 VTAIL.n182 6.59444
R827 VTAIL.n219 VTAIL.n182 6.59444
R828 VTAIL.n552 VTAIL.n515 6.59444
R829 VTAIL.n549 VTAIL.n515 6.59444
R830 VTAIL.n468 VTAIL.n431 6.59444
R831 VTAIL.n465 VTAIL.n431 6.59444
R832 VTAIL.n386 VTAIL.n349 6.59444
R833 VTAIL.n383 VTAIL.n349 6.59444
R834 VTAIL.n302 VTAIL.n265 6.59444
R835 VTAIL.n299 VTAIL.n265 6.59444
R836 VTAIL.n629 VTAIL.n598 5.81868
R837 VTAIL.n634 VTAIL.n594 5.81868
R838 VTAIL.n49 VTAIL.n18 5.81868
R839 VTAIL.n54 VTAIL.n14 5.81868
R840 VTAIL.n131 VTAIL.n100 5.81868
R841 VTAIL.n136 VTAIL.n96 5.81868
R842 VTAIL.n215 VTAIL.n184 5.81868
R843 VTAIL.n220 VTAIL.n180 5.81868
R844 VTAIL.n553 VTAIL.n513 5.81868
R845 VTAIL.n548 VTAIL.n517 5.81868
R846 VTAIL.n469 VTAIL.n429 5.81868
R847 VTAIL.n464 VTAIL.n433 5.81868
R848 VTAIL.n387 VTAIL.n347 5.81868
R849 VTAIL.n382 VTAIL.n351 5.81868
R850 VTAIL.n303 VTAIL.n263 5.81868
R851 VTAIL.n298 VTAIL.n267 5.81868
R852 VTAIL.n626 VTAIL.n625 5.04292
R853 VTAIL.n638 VTAIL.n637 5.04292
R854 VTAIL.n46 VTAIL.n45 5.04292
R855 VTAIL.n58 VTAIL.n57 5.04292
R856 VTAIL.n128 VTAIL.n127 5.04292
R857 VTAIL.n140 VTAIL.n139 5.04292
R858 VTAIL.n212 VTAIL.n211 5.04292
R859 VTAIL.n224 VTAIL.n223 5.04292
R860 VTAIL.n557 VTAIL.n556 5.04292
R861 VTAIL.n545 VTAIL.n544 5.04292
R862 VTAIL.n473 VTAIL.n472 5.04292
R863 VTAIL.n461 VTAIL.n460 5.04292
R864 VTAIL.n391 VTAIL.n390 5.04292
R865 VTAIL.n379 VTAIL.n378 5.04292
R866 VTAIL.n307 VTAIL.n306 5.04292
R867 VTAIL.n295 VTAIL.n294 5.04292
R868 VTAIL.n530 VTAIL.n526 4.38563
R869 VTAIL.n446 VTAIL.n442 4.38563
R870 VTAIL.n364 VTAIL.n360 4.38563
R871 VTAIL.n280 VTAIL.n276 4.38563
R872 VTAIL.n611 VTAIL.n607 4.38563
R873 VTAIL.n31 VTAIL.n27 4.38563
R874 VTAIL.n113 VTAIL.n109 4.38563
R875 VTAIL.n197 VTAIL.n193 4.38563
R876 VTAIL.n622 VTAIL.n600 4.26717
R877 VTAIL.n641 VTAIL.n592 4.26717
R878 VTAIL.n42 VTAIL.n20 4.26717
R879 VTAIL.n61 VTAIL.n12 4.26717
R880 VTAIL.n124 VTAIL.n102 4.26717
R881 VTAIL.n143 VTAIL.n94 4.26717
R882 VTAIL.n208 VTAIL.n186 4.26717
R883 VTAIL.n227 VTAIL.n178 4.26717
R884 VTAIL.n560 VTAIL.n511 4.26717
R885 VTAIL.n541 VTAIL.n519 4.26717
R886 VTAIL.n476 VTAIL.n427 4.26717
R887 VTAIL.n457 VTAIL.n435 4.26717
R888 VTAIL.n394 VTAIL.n345 4.26717
R889 VTAIL.n375 VTAIL.n353 4.26717
R890 VTAIL.n310 VTAIL.n261 4.26717
R891 VTAIL.n291 VTAIL.n269 4.26717
R892 VTAIL.n333 VTAIL.n331 3.64705
R893 VTAIL.n415 VTAIL.n333 3.64705
R894 VTAIL.n499 VTAIL.n497 3.64705
R895 VTAIL.n581 VTAIL.n499 3.64705
R896 VTAIL.n249 VTAIL.n167 3.64705
R897 VTAIL.n167 VTAIL.n165 3.64705
R898 VTAIL.n83 VTAIL.n1 3.64705
R899 VTAIL VTAIL.n663 3.58886
R900 VTAIL.n621 VTAIL.n602 3.49141
R901 VTAIL.n642 VTAIL.n590 3.49141
R902 VTAIL.n41 VTAIL.n22 3.49141
R903 VTAIL.n62 VTAIL.n10 3.49141
R904 VTAIL.n123 VTAIL.n104 3.49141
R905 VTAIL.n144 VTAIL.n92 3.49141
R906 VTAIL.n207 VTAIL.n188 3.49141
R907 VTAIL.n228 VTAIL.n176 3.49141
R908 VTAIL.n561 VTAIL.n509 3.49141
R909 VTAIL.n540 VTAIL.n521 3.49141
R910 VTAIL.n477 VTAIL.n425 3.49141
R911 VTAIL.n456 VTAIL.n437 3.49141
R912 VTAIL.n395 VTAIL.n343 3.49141
R913 VTAIL.n374 VTAIL.n355 3.49141
R914 VTAIL.n311 VTAIL.n259 3.49141
R915 VTAIL.n290 VTAIL.n271 3.49141
R916 VTAIL.n618 VTAIL.n617 2.71565
R917 VTAIL.n646 VTAIL.n645 2.71565
R918 VTAIL.n38 VTAIL.n37 2.71565
R919 VTAIL.n66 VTAIL.n65 2.71565
R920 VTAIL.n120 VTAIL.n119 2.71565
R921 VTAIL.n148 VTAIL.n147 2.71565
R922 VTAIL.n204 VTAIL.n203 2.71565
R923 VTAIL.n232 VTAIL.n231 2.71565
R924 VTAIL.n565 VTAIL.n564 2.71565
R925 VTAIL.n537 VTAIL.n536 2.71565
R926 VTAIL.n481 VTAIL.n480 2.71565
R927 VTAIL.n453 VTAIL.n452 2.71565
R928 VTAIL.n399 VTAIL.n398 2.71565
R929 VTAIL.n371 VTAIL.n370 2.71565
R930 VTAIL.n315 VTAIL.n314 2.71565
R931 VTAIL.n287 VTAIL.n286 2.71565
R932 VTAIL.n614 VTAIL.n604 1.93989
R933 VTAIL.n650 VTAIL.n588 1.93989
R934 VTAIL.n662 VTAIL.n582 1.93989
R935 VTAIL.n34 VTAIL.n24 1.93989
R936 VTAIL.n70 VTAIL.n8 1.93989
R937 VTAIL.n82 VTAIL.n2 1.93989
R938 VTAIL.n116 VTAIL.n106 1.93989
R939 VTAIL.n152 VTAIL.n90 1.93989
R940 VTAIL.n164 VTAIL.n84 1.93989
R941 VTAIL.n200 VTAIL.n190 1.93989
R942 VTAIL.n236 VTAIL.n174 1.93989
R943 VTAIL.n248 VTAIL.n168 1.93989
R944 VTAIL.n580 VTAIL.n500 1.93989
R945 VTAIL.n568 VTAIL.n506 1.93989
R946 VTAIL.n533 VTAIL.n523 1.93989
R947 VTAIL.n496 VTAIL.n416 1.93989
R948 VTAIL.n484 VTAIL.n422 1.93989
R949 VTAIL.n449 VTAIL.n439 1.93989
R950 VTAIL.n414 VTAIL.n334 1.93989
R951 VTAIL.n402 VTAIL.n340 1.93989
R952 VTAIL.n367 VTAIL.n357 1.93989
R953 VTAIL.n330 VTAIL.n250 1.93989
R954 VTAIL.n318 VTAIL.n256 1.93989
R955 VTAIL.n283 VTAIL.n273 1.93989
R956 VTAIL.n0 VTAIL.t7 1.34015
R957 VTAIL.n0 VTAIL.t4 1.34015
R958 VTAIL.n166 VTAIL.t11 1.34015
R959 VTAIL.n166 VTAIL.t8 1.34015
R960 VTAIL.n498 VTAIL.t10 1.34015
R961 VTAIL.n498 VTAIL.t9 1.34015
R962 VTAIL.n332 VTAIL.t2 1.34015
R963 VTAIL.n332 VTAIL.t6 1.34015
R964 VTAIL.n613 VTAIL.n606 1.16414
R965 VTAIL.n651 VTAIL.n586 1.16414
R966 VTAIL.n660 VTAIL.n659 1.16414
R967 VTAIL.n33 VTAIL.n26 1.16414
R968 VTAIL.n71 VTAIL.n6 1.16414
R969 VTAIL.n80 VTAIL.n79 1.16414
R970 VTAIL.n115 VTAIL.n108 1.16414
R971 VTAIL.n153 VTAIL.n88 1.16414
R972 VTAIL.n162 VTAIL.n161 1.16414
R973 VTAIL.n199 VTAIL.n192 1.16414
R974 VTAIL.n237 VTAIL.n172 1.16414
R975 VTAIL.n246 VTAIL.n245 1.16414
R976 VTAIL.n578 VTAIL.n577 1.16414
R977 VTAIL.n569 VTAIL.n504 1.16414
R978 VTAIL.n532 VTAIL.n525 1.16414
R979 VTAIL.n494 VTAIL.n493 1.16414
R980 VTAIL.n485 VTAIL.n420 1.16414
R981 VTAIL.n448 VTAIL.n441 1.16414
R982 VTAIL.n412 VTAIL.n411 1.16414
R983 VTAIL.n403 VTAIL.n338 1.16414
R984 VTAIL.n366 VTAIL.n359 1.16414
R985 VTAIL.n328 VTAIL.n327 1.16414
R986 VTAIL.n319 VTAIL.n254 1.16414
R987 VTAIL.n282 VTAIL.n275 1.16414
R988 VTAIL.n497 VTAIL.n415 0.470328
R989 VTAIL.n165 VTAIL.n83 0.470328
R990 VTAIL.n610 VTAIL.n609 0.388379
R991 VTAIL.n655 VTAIL.n654 0.388379
R992 VTAIL.n656 VTAIL.n584 0.388379
R993 VTAIL.n30 VTAIL.n29 0.388379
R994 VTAIL.n75 VTAIL.n74 0.388379
R995 VTAIL.n76 VTAIL.n4 0.388379
R996 VTAIL.n112 VTAIL.n111 0.388379
R997 VTAIL.n157 VTAIL.n156 0.388379
R998 VTAIL.n158 VTAIL.n86 0.388379
R999 VTAIL.n196 VTAIL.n195 0.388379
R1000 VTAIL.n241 VTAIL.n240 0.388379
R1001 VTAIL.n242 VTAIL.n170 0.388379
R1002 VTAIL.n574 VTAIL.n502 0.388379
R1003 VTAIL.n573 VTAIL.n572 0.388379
R1004 VTAIL.n529 VTAIL.n528 0.388379
R1005 VTAIL.n490 VTAIL.n418 0.388379
R1006 VTAIL.n489 VTAIL.n488 0.388379
R1007 VTAIL.n445 VTAIL.n444 0.388379
R1008 VTAIL.n408 VTAIL.n336 0.388379
R1009 VTAIL.n407 VTAIL.n406 0.388379
R1010 VTAIL.n363 VTAIL.n362 0.388379
R1011 VTAIL.n324 VTAIL.n252 0.388379
R1012 VTAIL.n323 VTAIL.n322 0.388379
R1013 VTAIL.n279 VTAIL.n278 0.388379
R1014 VTAIL.n612 VTAIL.n611 0.155672
R1015 VTAIL.n612 VTAIL.n603 0.155672
R1016 VTAIL.n619 VTAIL.n603 0.155672
R1017 VTAIL.n620 VTAIL.n619 0.155672
R1018 VTAIL.n620 VTAIL.n599 0.155672
R1019 VTAIL.n627 VTAIL.n599 0.155672
R1020 VTAIL.n628 VTAIL.n627 0.155672
R1021 VTAIL.n628 VTAIL.n595 0.155672
R1022 VTAIL.n635 VTAIL.n595 0.155672
R1023 VTAIL.n636 VTAIL.n635 0.155672
R1024 VTAIL.n636 VTAIL.n591 0.155672
R1025 VTAIL.n643 VTAIL.n591 0.155672
R1026 VTAIL.n644 VTAIL.n643 0.155672
R1027 VTAIL.n644 VTAIL.n587 0.155672
R1028 VTAIL.n652 VTAIL.n587 0.155672
R1029 VTAIL.n653 VTAIL.n652 0.155672
R1030 VTAIL.n653 VTAIL.n583 0.155672
R1031 VTAIL.n661 VTAIL.n583 0.155672
R1032 VTAIL.n32 VTAIL.n31 0.155672
R1033 VTAIL.n32 VTAIL.n23 0.155672
R1034 VTAIL.n39 VTAIL.n23 0.155672
R1035 VTAIL.n40 VTAIL.n39 0.155672
R1036 VTAIL.n40 VTAIL.n19 0.155672
R1037 VTAIL.n47 VTAIL.n19 0.155672
R1038 VTAIL.n48 VTAIL.n47 0.155672
R1039 VTAIL.n48 VTAIL.n15 0.155672
R1040 VTAIL.n55 VTAIL.n15 0.155672
R1041 VTAIL.n56 VTAIL.n55 0.155672
R1042 VTAIL.n56 VTAIL.n11 0.155672
R1043 VTAIL.n63 VTAIL.n11 0.155672
R1044 VTAIL.n64 VTAIL.n63 0.155672
R1045 VTAIL.n64 VTAIL.n7 0.155672
R1046 VTAIL.n72 VTAIL.n7 0.155672
R1047 VTAIL.n73 VTAIL.n72 0.155672
R1048 VTAIL.n73 VTAIL.n3 0.155672
R1049 VTAIL.n81 VTAIL.n3 0.155672
R1050 VTAIL.n114 VTAIL.n113 0.155672
R1051 VTAIL.n114 VTAIL.n105 0.155672
R1052 VTAIL.n121 VTAIL.n105 0.155672
R1053 VTAIL.n122 VTAIL.n121 0.155672
R1054 VTAIL.n122 VTAIL.n101 0.155672
R1055 VTAIL.n129 VTAIL.n101 0.155672
R1056 VTAIL.n130 VTAIL.n129 0.155672
R1057 VTAIL.n130 VTAIL.n97 0.155672
R1058 VTAIL.n137 VTAIL.n97 0.155672
R1059 VTAIL.n138 VTAIL.n137 0.155672
R1060 VTAIL.n138 VTAIL.n93 0.155672
R1061 VTAIL.n145 VTAIL.n93 0.155672
R1062 VTAIL.n146 VTAIL.n145 0.155672
R1063 VTAIL.n146 VTAIL.n89 0.155672
R1064 VTAIL.n154 VTAIL.n89 0.155672
R1065 VTAIL.n155 VTAIL.n154 0.155672
R1066 VTAIL.n155 VTAIL.n85 0.155672
R1067 VTAIL.n163 VTAIL.n85 0.155672
R1068 VTAIL.n198 VTAIL.n197 0.155672
R1069 VTAIL.n198 VTAIL.n189 0.155672
R1070 VTAIL.n205 VTAIL.n189 0.155672
R1071 VTAIL.n206 VTAIL.n205 0.155672
R1072 VTAIL.n206 VTAIL.n185 0.155672
R1073 VTAIL.n213 VTAIL.n185 0.155672
R1074 VTAIL.n214 VTAIL.n213 0.155672
R1075 VTAIL.n214 VTAIL.n181 0.155672
R1076 VTAIL.n221 VTAIL.n181 0.155672
R1077 VTAIL.n222 VTAIL.n221 0.155672
R1078 VTAIL.n222 VTAIL.n177 0.155672
R1079 VTAIL.n229 VTAIL.n177 0.155672
R1080 VTAIL.n230 VTAIL.n229 0.155672
R1081 VTAIL.n230 VTAIL.n173 0.155672
R1082 VTAIL.n238 VTAIL.n173 0.155672
R1083 VTAIL.n239 VTAIL.n238 0.155672
R1084 VTAIL.n239 VTAIL.n169 0.155672
R1085 VTAIL.n247 VTAIL.n169 0.155672
R1086 VTAIL.n579 VTAIL.n501 0.155672
R1087 VTAIL.n571 VTAIL.n501 0.155672
R1088 VTAIL.n571 VTAIL.n570 0.155672
R1089 VTAIL.n570 VTAIL.n505 0.155672
R1090 VTAIL.n563 VTAIL.n505 0.155672
R1091 VTAIL.n563 VTAIL.n562 0.155672
R1092 VTAIL.n562 VTAIL.n510 0.155672
R1093 VTAIL.n555 VTAIL.n510 0.155672
R1094 VTAIL.n555 VTAIL.n554 0.155672
R1095 VTAIL.n554 VTAIL.n514 0.155672
R1096 VTAIL.n547 VTAIL.n514 0.155672
R1097 VTAIL.n547 VTAIL.n546 0.155672
R1098 VTAIL.n546 VTAIL.n518 0.155672
R1099 VTAIL.n539 VTAIL.n518 0.155672
R1100 VTAIL.n539 VTAIL.n538 0.155672
R1101 VTAIL.n538 VTAIL.n522 0.155672
R1102 VTAIL.n531 VTAIL.n522 0.155672
R1103 VTAIL.n531 VTAIL.n530 0.155672
R1104 VTAIL.n495 VTAIL.n417 0.155672
R1105 VTAIL.n487 VTAIL.n417 0.155672
R1106 VTAIL.n487 VTAIL.n486 0.155672
R1107 VTAIL.n486 VTAIL.n421 0.155672
R1108 VTAIL.n479 VTAIL.n421 0.155672
R1109 VTAIL.n479 VTAIL.n478 0.155672
R1110 VTAIL.n478 VTAIL.n426 0.155672
R1111 VTAIL.n471 VTAIL.n426 0.155672
R1112 VTAIL.n471 VTAIL.n470 0.155672
R1113 VTAIL.n470 VTAIL.n430 0.155672
R1114 VTAIL.n463 VTAIL.n430 0.155672
R1115 VTAIL.n463 VTAIL.n462 0.155672
R1116 VTAIL.n462 VTAIL.n434 0.155672
R1117 VTAIL.n455 VTAIL.n434 0.155672
R1118 VTAIL.n455 VTAIL.n454 0.155672
R1119 VTAIL.n454 VTAIL.n438 0.155672
R1120 VTAIL.n447 VTAIL.n438 0.155672
R1121 VTAIL.n447 VTAIL.n446 0.155672
R1122 VTAIL.n413 VTAIL.n335 0.155672
R1123 VTAIL.n405 VTAIL.n335 0.155672
R1124 VTAIL.n405 VTAIL.n404 0.155672
R1125 VTAIL.n404 VTAIL.n339 0.155672
R1126 VTAIL.n397 VTAIL.n339 0.155672
R1127 VTAIL.n397 VTAIL.n396 0.155672
R1128 VTAIL.n396 VTAIL.n344 0.155672
R1129 VTAIL.n389 VTAIL.n344 0.155672
R1130 VTAIL.n389 VTAIL.n388 0.155672
R1131 VTAIL.n388 VTAIL.n348 0.155672
R1132 VTAIL.n381 VTAIL.n348 0.155672
R1133 VTAIL.n381 VTAIL.n380 0.155672
R1134 VTAIL.n380 VTAIL.n352 0.155672
R1135 VTAIL.n373 VTAIL.n352 0.155672
R1136 VTAIL.n373 VTAIL.n372 0.155672
R1137 VTAIL.n372 VTAIL.n356 0.155672
R1138 VTAIL.n365 VTAIL.n356 0.155672
R1139 VTAIL.n365 VTAIL.n364 0.155672
R1140 VTAIL.n329 VTAIL.n251 0.155672
R1141 VTAIL.n321 VTAIL.n251 0.155672
R1142 VTAIL.n321 VTAIL.n320 0.155672
R1143 VTAIL.n320 VTAIL.n255 0.155672
R1144 VTAIL.n313 VTAIL.n255 0.155672
R1145 VTAIL.n313 VTAIL.n312 0.155672
R1146 VTAIL.n312 VTAIL.n260 0.155672
R1147 VTAIL.n305 VTAIL.n260 0.155672
R1148 VTAIL.n305 VTAIL.n304 0.155672
R1149 VTAIL.n304 VTAIL.n264 0.155672
R1150 VTAIL.n297 VTAIL.n264 0.155672
R1151 VTAIL.n297 VTAIL.n296 0.155672
R1152 VTAIL.n296 VTAIL.n268 0.155672
R1153 VTAIL.n289 VTAIL.n268 0.155672
R1154 VTAIL.n289 VTAIL.n288 0.155672
R1155 VTAIL.n288 VTAIL.n272 0.155672
R1156 VTAIL.n281 VTAIL.n272 0.155672
R1157 VTAIL.n281 VTAIL.n280 0.155672
R1158 VTAIL VTAIL.n1 0.0586897
R1159 VDD1 VDD1.n0 65.5177
R1160 VDD1.n3 VDD1.n2 65.404
R1161 VDD1.n3 VDD1.n1 65.404
R1162 VDD1.n5 VDD1.n4 63.6361
R1163 VDD1.n5 VDD1.n3 53.4492
R1164 VDD1 VDD1.n5 1.76559
R1165 VDD1.n4 VDD1.t3 1.34015
R1166 VDD1.n4 VDD1.t6 1.34015
R1167 VDD1.n0 VDD1.t4 1.34015
R1168 VDD1.n0 VDD1.t7 1.34015
R1169 VDD1.n2 VDD1.t5 1.34015
R1170 VDD1.n2 VDD1.t1 1.34015
R1171 VDD1.n1 VDD1.t0 1.34015
R1172 VDD1.n1 VDD1.t2 1.34015
R1173 B.n905 B.n904 585
R1174 B.n905 B.n128 585
R1175 B.n908 B.n907 585
R1176 B.n909 B.n187 585
R1177 B.n911 B.n910 585
R1178 B.n913 B.n186 585
R1179 B.n916 B.n915 585
R1180 B.n917 B.n185 585
R1181 B.n919 B.n918 585
R1182 B.n921 B.n184 585
R1183 B.n924 B.n923 585
R1184 B.n925 B.n183 585
R1185 B.n927 B.n926 585
R1186 B.n929 B.n182 585
R1187 B.n932 B.n931 585
R1188 B.n933 B.n181 585
R1189 B.n935 B.n934 585
R1190 B.n937 B.n180 585
R1191 B.n940 B.n939 585
R1192 B.n941 B.n179 585
R1193 B.n943 B.n942 585
R1194 B.n945 B.n178 585
R1195 B.n948 B.n947 585
R1196 B.n949 B.n177 585
R1197 B.n951 B.n950 585
R1198 B.n953 B.n176 585
R1199 B.n956 B.n955 585
R1200 B.n957 B.n175 585
R1201 B.n959 B.n958 585
R1202 B.n961 B.n174 585
R1203 B.n964 B.n963 585
R1204 B.n965 B.n173 585
R1205 B.n967 B.n966 585
R1206 B.n969 B.n172 585
R1207 B.n972 B.n971 585
R1208 B.n973 B.n171 585
R1209 B.n975 B.n974 585
R1210 B.n977 B.n170 585
R1211 B.n980 B.n979 585
R1212 B.n981 B.n169 585
R1213 B.n983 B.n982 585
R1214 B.n985 B.n168 585
R1215 B.n988 B.n987 585
R1216 B.n989 B.n167 585
R1217 B.n991 B.n990 585
R1218 B.n993 B.n166 585
R1219 B.n996 B.n995 585
R1220 B.n997 B.n165 585
R1221 B.n999 B.n998 585
R1222 B.n1001 B.n164 585
R1223 B.n1004 B.n1003 585
R1224 B.n1006 B.n161 585
R1225 B.n1008 B.n1007 585
R1226 B.n1010 B.n160 585
R1227 B.n1013 B.n1012 585
R1228 B.n1014 B.n159 585
R1229 B.n1016 B.n1015 585
R1230 B.n1018 B.n158 585
R1231 B.n1020 B.n1019 585
R1232 B.n1022 B.n1021 585
R1233 B.n1025 B.n1024 585
R1234 B.n1026 B.n153 585
R1235 B.n1028 B.n1027 585
R1236 B.n1030 B.n152 585
R1237 B.n1033 B.n1032 585
R1238 B.n1034 B.n151 585
R1239 B.n1036 B.n1035 585
R1240 B.n1038 B.n150 585
R1241 B.n1041 B.n1040 585
R1242 B.n1042 B.n149 585
R1243 B.n1044 B.n1043 585
R1244 B.n1046 B.n148 585
R1245 B.n1049 B.n1048 585
R1246 B.n1050 B.n147 585
R1247 B.n1052 B.n1051 585
R1248 B.n1054 B.n146 585
R1249 B.n1057 B.n1056 585
R1250 B.n1058 B.n145 585
R1251 B.n1060 B.n1059 585
R1252 B.n1062 B.n144 585
R1253 B.n1065 B.n1064 585
R1254 B.n1066 B.n143 585
R1255 B.n1068 B.n1067 585
R1256 B.n1070 B.n142 585
R1257 B.n1073 B.n1072 585
R1258 B.n1074 B.n141 585
R1259 B.n1076 B.n1075 585
R1260 B.n1078 B.n140 585
R1261 B.n1081 B.n1080 585
R1262 B.n1082 B.n139 585
R1263 B.n1084 B.n1083 585
R1264 B.n1086 B.n138 585
R1265 B.n1089 B.n1088 585
R1266 B.n1090 B.n137 585
R1267 B.n1092 B.n1091 585
R1268 B.n1094 B.n136 585
R1269 B.n1097 B.n1096 585
R1270 B.n1098 B.n135 585
R1271 B.n1100 B.n1099 585
R1272 B.n1102 B.n134 585
R1273 B.n1105 B.n1104 585
R1274 B.n1106 B.n133 585
R1275 B.n1108 B.n1107 585
R1276 B.n1110 B.n132 585
R1277 B.n1113 B.n1112 585
R1278 B.n1114 B.n131 585
R1279 B.n1116 B.n1115 585
R1280 B.n1118 B.n130 585
R1281 B.n1121 B.n1120 585
R1282 B.n1122 B.n129 585
R1283 B.n903 B.n127 585
R1284 B.n1125 B.n127 585
R1285 B.n902 B.n126 585
R1286 B.n1126 B.n126 585
R1287 B.n901 B.n125 585
R1288 B.n1127 B.n125 585
R1289 B.n900 B.n899 585
R1290 B.n899 B.n121 585
R1291 B.n898 B.n120 585
R1292 B.n1133 B.n120 585
R1293 B.n897 B.n119 585
R1294 B.n1134 B.n119 585
R1295 B.n896 B.n118 585
R1296 B.n1135 B.n118 585
R1297 B.n895 B.n894 585
R1298 B.n894 B.n114 585
R1299 B.n893 B.n113 585
R1300 B.n1141 B.n113 585
R1301 B.n892 B.n112 585
R1302 B.n1142 B.n112 585
R1303 B.n891 B.n111 585
R1304 B.n1143 B.n111 585
R1305 B.n890 B.n889 585
R1306 B.n889 B.n107 585
R1307 B.n888 B.n106 585
R1308 B.n1149 B.n106 585
R1309 B.n887 B.n105 585
R1310 B.n1150 B.n105 585
R1311 B.n886 B.n104 585
R1312 B.n1151 B.n104 585
R1313 B.n885 B.n884 585
R1314 B.n884 B.n100 585
R1315 B.n883 B.n99 585
R1316 B.n1157 B.n99 585
R1317 B.n882 B.n98 585
R1318 B.n1158 B.n98 585
R1319 B.n881 B.n97 585
R1320 B.n1159 B.n97 585
R1321 B.n880 B.n879 585
R1322 B.n879 B.n93 585
R1323 B.n878 B.n92 585
R1324 B.n1165 B.n92 585
R1325 B.n877 B.n91 585
R1326 B.n1166 B.n91 585
R1327 B.n876 B.n90 585
R1328 B.n1167 B.n90 585
R1329 B.n875 B.n874 585
R1330 B.n874 B.n86 585
R1331 B.n873 B.n85 585
R1332 B.n1173 B.n85 585
R1333 B.n872 B.n84 585
R1334 B.n1174 B.n84 585
R1335 B.n871 B.n83 585
R1336 B.n1175 B.n83 585
R1337 B.n870 B.n869 585
R1338 B.n869 B.n79 585
R1339 B.n868 B.n78 585
R1340 B.n1181 B.n78 585
R1341 B.n867 B.n77 585
R1342 B.n1182 B.n77 585
R1343 B.n866 B.n76 585
R1344 B.n1183 B.n76 585
R1345 B.n865 B.n864 585
R1346 B.n864 B.n72 585
R1347 B.n863 B.n71 585
R1348 B.n1189 B.n71 585
R1349 B.n862 B.n70 585
R1350 B.n1190 B.n70 585
R1351 B.n861 B.n69 585
R1352 B.n1191 B.n69 585
R1353 B.n860 B.n859 585
R1354 B.n859 B.n65 585
R1355 B.n858 B.n64 585
R1356 B.n1197 B.n64 585
R1357 B.n857 B.n63 585
R1358 B.n1198 B.n63 585
R1359 B.n856 B.n62 585
R1360 B.n1199 B.n62 585
R1361 B.n855 B.n854 585
R1362 B.n854 B.n58 585
R1363 B.n853 B.n57 585
R1364 B.n1205 B.n57 585
R1365 B.n852 B.n56 585
R1366 B.n1206 B.n56 585
R1367 B.n851 B.n55 585
R1368 B.n1207 B.n55 585
R1369 B.n850 B.n849 585
R1370 B.n849 B.n51 585
R1371 B.n848 B.n50 585
R1372 B.n1213 B.n50 585
R1373 B.n847 B.n49 585
R1374 B.n1214 B.n49 585
R1375 B.n846 B.n48 585
R1376 B.n1215 B.n48 585
R1377 B.n845 B.n844 585
R1378 B.n844 B.n44 585
R1379 B.n843 B.n43 585
R1380 B.n1221 B.n43 585
R1381 B.n842 B.n42 585
R1382 B.n1222 B.n42 585
R1383 B.n841 B.n41 585
R1384 B.n1223 B.n41 585
R1385 B.n840 B.n839 585
R1386 B.n839 B.n37 585
R1387 B.n838 B.n36 585
R1388 B.n1229 B.n36 585
R1389 B.n837 B.n35 585
R1390 B.n1230 B.n35 585
R1391 B.n836 B.n34 585
R1392 B.n1231 B.n34 585
R1393 B.n835 B.n834 585
R1394 B.n834 B.n30 585
R1395 B.n833 B.n29 585
R1396 B.n1237 B.n29 585
R1397 B.n832 B.n28 585
R1398 B.n1238 B.n28 585
R1399 B.n831 B.n27 585
R1400 B.n1239 B.n27 585
R1401 B.n830 B.n829 585
R1402 B.n829 B.n23 585
R1403 B.n828 B.n22 585
R1404 B.n1245 B.n22 585
R1405 B.n827 B.n21 585
R1406 B.n1246 B.n21 585
R1407 B.n826 B.n20 585
R1408 B.n1247 B.n20 585
R1409 B.n825 B.n824 585
R1410 B.n824 B.n16 585
R1411 B.n823 B.n15 585
R1412 B.n1253 B.n15 585
R1413 B.n822 B.n14 585
R1414 B.n1254 B.n14 585
R1415 B.n821 B.n13 585
R1416 B.n1255 B.n13 585
R1417 B.n820 B.n819 585
R1418 B.n819 B.n12 585
R1419 B.n818 B.n817 585
R1420 B.n818 B.n8 585
R1421 B.n816 B.n7 585
R1422 B.n1262 B.n7 585
R1423 B.n815 B.n6 585
R1424 B.n1263 B.n6 585
R1425 B.n814 B.n5 585
R1426 B.n1264 B.n5 585
R1427 B.n813 B.n812 585
R1428 B.n812 B.n4 585
R1429 B.n811 B.n188 585
R1430 B.n811 B.n810 585
R1431 B.n801 B.n189 585
R1432 B.n190 B.n189 585
R1433 B.n803 B.n802 585
R1434 B.n804 B.n803 585
R1435 B.n800 B.n195 585
R1436 B.n195 B.n194 585
R1437 B.n799 B.n798 585
R1438 B.n798 B.n797 585
R1439 B.n197 B.n196 585
R1440 B.n198 B.n197 585
R1441 B.n790 B.n789 585
R1442 B.n791 B.n790 585
R1443 B.n788 B.n203 585
R1444 B.n203 B.n202 585
R1445 B.n787 B.n786 585
R1446 B.n786 B.n785 585
R1447 B.n205 B.n204 585
R1448 B.n206 B.n205 585
R1449 B.n778 B.n777 585
R1450 B.n779 B.n778 585
R1451 B.n776 B.n211 585
R1452 B.n211 B.n210 585
R1453 B.n775 B.n774 585
R1454 B.n774 B.n773 585
R1455 B.n213 B.n212 585
R1456 B.n214 B.n213 585
R1457 B.n766 B.n765 585
R1458 B.n767 B.n766 585
R1459 B.n764 B.n219 585
R1460 B.n219 B.n218 585
R1461 B.n763 B.n762 585
R1462 B.n762 B.n761 585
R1463 B.n221 B.n220 585
R1464 B.n222 B.n221 585
R1465 B.n754 B.n753 585
R1466 B.n755 B.n754 585
R1467 B.n752 B.n227 585
R1468 B.n227 B.n226 585
R1469 B.n751 B.n750 585
R1470 B.n750 B.n749 585
R1471 B.n229 B.n228 585
R1472 B.n230 B.n229 585
R1473 B.n742 B.n741 585
R1474 B.n743 B.n742 585
R1475 B.n740 B.n235 585
R1476 B.n235 B.n234 585
R1477 B.n739 B.n738 585
R1478 B.n738 B.n737 585
R1479 B.n237 B.n236 585
R1480 B.n238 B.n237 585
R1481 B.n730 B.n729 585
R1482 B.n731 B.n730 585
R1483 B.n728 B.n243 585
R1484 B.n243 B.n242 585
R1485 B.n727 B.n726 585
R1486 B.n726 B.n725 585
R1487 B.n245 B.n244 585
R1488 B.n246 B.n245 585
R1489 B.n718 B.n717 585
R1490 B.n719 B.n718 585
R1491 B.n716 B.n250 585
R1492 B.n254 B.n250 585
R1493 B.n715 B.n714 585
R1494 B.n714 B.n713 585
R1495 B.n252 B.n251 585
R1496 B.n253 B.n252 585
R1497 B.n706 B.n705 585
R1498 B.n707 B.n706 585
R1499 B.n704 B.n259 585
R1500 B.n259 B.n258 585
R1501 B.n703 B.n702 585
R1502 B.n702 B.n701 585
R1503 B.n261 B.n260 585
R1504 B.n262 B.n261 585
R1505 B.n694 B.n693 585
R1506 B.n695 B.n694 585
R1507 B.n692 B.n267 585
R1508 B.n267 B.n266 585
R1509 B.n691 B.n690 585
R1510 B.n690 B.n689 585
R1511 B.n269 B.n268 585
R1512 B.n270 B.n269 585
R1513 B.n682 B.n681 585
R1514 B.n683 B.n682 585
R1515 B.n680 B.n274 585
R1516 B.n278 B.n274 585
R1517 B.n679 B.n678 585
R1518 B.n678 B.n677 585
R1519 B.n276 B.n275 585
R1520 B.n277 B.n276 585
R1521 B.n670 B.n669 585
R1522 B.n671 B.n670 585
R1523 B.n668 B.n283 585
R1524 B.n283 B.n282 585
R1525 B.n667 B.n666 585
R1526 B.n666 B.n665 585
R1527 B.n285 B.n284 585
R1528 B.n286 B.n285 585
R1529 B.n658 B.n657 585
R1530 B.n659 B.n658 585
R1531 B.n656 B.n291 585
R1532 B.n291 B.n290 585
R1533 B.n655 B.n654 585
R1534 B.n654 B.n653 585
R1535 B.n293 B.n292 585
R1536 B.n294 B.n293 585
R1537 B.n646 B.n645 585
R1538 B.n647 B.n646 585
R1539 B.n644 B.n299 585
R1540 B.n299 B.n298 585
R1541 B.n643 B.n642 585
R1542 B.n642 B.n641 585
R1543 B.n301 B.n300 585
R1544 B.n302 B.n301 585
R1545 B.n634 B.n633 585
R1546 B.n635 B.n634 585
R1547 B.n632 B.n306 585
R1548 B.n310 B.n306 585
R1549 B.n631 B.n630 585
R1550 B.n630 B.n629 585
R1551 B.n308 B.n307 585
R1552 B.n309 B.n308 585
R1553 B.n622 B.n621 585
R1554 B.n623 B.n622 585
R1555 B.n620 B.n315 585
R1556 B.n315 B.n314 585
R1557 B.n619 B.n618 585
R1558 B.n618 B.n617 585
R1559 B.n317 B.n316 585
R1560 B.n318 B.n317 585
R1561 B.n610 B.n609 585
R1562 B.n611 B.n610 585
R1563 B.n608 B.n323 585
R1564 B.n323 B.n322 585
R1565 B.n607 B.n606 585
R1566 B.n606 B.n605 585
R1567 B.n602 B.n327 585
R1568 B.n601 B.n600 585
R1569 B.n598 B.n328 585
R1570 B.n598 B.n326 585
R1571 B.n597 B.n596 585
R1572 B.n595 B.n594 585
R1573 B.n593 B.n330 585
R1574 B.n591 B.n590 585
R1575 B.n589 B.n331 585
R1576 B.n588 B.n587 585
R1577 B.n585 B.n332 585
R1578 B.n583 B.n582 585
R1579 B.n581 B.n333 585
R1580 B.n580 B.n579 585
R1581 B.n577 B.n334 585
R1582 B.n575 B.n574 585
R1583 B.n573 B.n335 585
R1584 B.n572 B.n571 585
R1585 B.n569 B.n336 585
R1586 B.n567 B.n566 585
R1587 B.n565 B.n337 585
R1588 B.n564 B.n563 585
R1589 B.n561 B.n338 585
R1590 B.n559 B.n558 585
R1591 B.n557 B.n339 585
R1592 B.n556 B.n555 585
R1593 B.n553 B.n340 585
R1594 B.n551 B.n550 585
R1595 B.n549 B.n341 585
R1596 B.n548 B.n547 585
R1597 B.n545 B.n342 585
R1598 B.n543 B.n542 585
R1599 B.n541 B.n343 585
R1600 B.n540 B.n539 585
R1601 B.n537 B.n344 585
R1602 B.n535 B.n534 585
R1603 B.n533 B.n345 585
R1604 B.n532 B.n531 585
R1605 B.n529 B.n346 585
R1606 B.n527 B.n526 585
R1607 B.n525 B.n347 585
R1608 B.n524 B.n523 585
R1609 B.n521 B.n348 585
R1610 B.n519 B.n518 585
R1611 B.n517 B.n349 585
R1612 B.n516 B.n515 585
R1613 B.n513 B.n350 585
R1614 B.n511 B.n510 585
R1615 B.n509 B.n351 585
R1616 B.n508 B.n507 585
R1617 B.n505 B.n352 585
R1618 B.n503 B.n502 585
R1619 B.n501 B.n353 585
R1620 B.n500 B.n499 585
R1621 B.n497 B.n357 585
R1622 B.n495 B.n494 585
R1623 B.n493 B.n358 585
R1624 B.n492 B.n491 585
R1625 B.n489 B.n359 585
R1626 B.n487 B.n486 585
R1627 B.n484 B.n360 585
R1628 B.n483 B.n482 585
R1629 B.n480 B.n363 585
R1630 B.n478 B.n477 585
R1631 B.n476 B.n364 585
R1632 B.n475 B.n474 585
R1633 B.n472 B.n365 585
R1634 B.n470 B.n469 585
R1635 B.n468 B.n366 585
R1636 B.n467 B.n466 585
R1637 B.n464 B.n367 585
R1638 B.n462 B.n461 585
R1639 B.n460 B.n368 585
R1640 B.n459 B.n458 585
R1641 B.n456 B.n369 585
R1642 B.n454 B.n453 585
R1643 B.n452 B.n370 585
R1644 B.n451 B.n450 585
R1645 B.n448 B.n371 585
R1646 B.n446 B.n445 585
R1647 B.n444 B.n372 585
R1648 B.n443 B.n442 585
R1649 B.n440 B.n373 585
R1650 B.n438 B.n437 585
R1651 B.n436 B.n374 585
R1652 B.n435 B.n434 585
R1653 B.n432 B.n375 585
R1654 B.n430 B.n429 585
R1655 B.n428 B.n376 585
R1656 B.n427 B.n426 585
R1657 B.n424 B.n377 585
R1658 B.n422 B.n421 585
R1659 B.n420 B.n378 585
R1660 B.n419 B.n418 585
R1661 B.n416 B.n379 585
R1662 B.n414 B.n413 585
R1663 B.n412 B.n380 585
R1664 B.n411 B.n410 585
R1665 B.n408 B.n381 585
R1666 B.n406 B.n405 585
R1667 B.n404 B.n382 585
R1668 B.n403 B.n402 585
R1669 B.n400 B.n383 585
R1670 B.n398 B.n397 585
R1671 B.n396 B.n384 585
R1672 B.n395 B.n394 585
R1673 B.n392 B.n385 585
R1674 B.n390 B.n389 585
R1675 B.n388 B.n387 585
R1676 B.n325 B.n324 585
R1677 B.n604 B.n603 585
R1678 B.n605 B.n604 585
R1679 B.n321 B.n320 585
R1680 B.n322 B.n321 585
R1681 B.n613 B.n612 585
R1682 B.n612 B.n611 585
R1683 B.n614 B.n319 585
R1684 B.n319 B.n318 585
R1685 B.n616 B.n615 585
R1686 B.n617 B.n616 585
R1687 B.n313 B.n312 585
R1688 B.n314 B.n313 585
R1689 B.n625 B.n624 585
R1690 B.n624 B.n623 585
R1691 B.n626 B.n311 585
R1692 B.n311 B.n309 585
R1693 B.n628 B.n627 585
R1694 B.n629 B.n628 585
R1695 B.n305 B.n304 585
R1696 B.n310 B.n305 585
R1697 B.n637 B.n636 585
R1698 B.n636 B.n635 585
R1699 B.n638 B.n303 585
R1700 B.n303 B.n302 585
R1701 B.n640 B.n639 585
R1702 B.n641 B.n640 585
R1703 B.n297 B.n296 585
R1704 B.n298 B.n297 585
R1705 B.n649 B.n648 585
R1706 B.n648 B.n647 585
R1707 B.n650 B.n295 585
R1708 B.n295 B.n294 585
R1709 B.n652 B.n651 585
R1710 B.n653 B.n652 585
R1711 B.n289 B.n288 585
R1712 B.n290 B.n289 585
R1713 B.n661 B.n660 585
R1714 B.n660 B.n659 585
R1715 B.n662 B.n287 585
R1716 B.n287 B.n286 585
R1717 B.n664 B.n663 585
R1718 B.n665 B.n664 585
R1719 B.n281 B.n280 585
R1720 B.n282 B.n281 585
R1721 B.n673 B.n672 585
R1722 B.n672 B.n671 585
R1723 B.n674 B.n279 585
R1724 B.n279 B.n277 585
R1725 B.n676 B.n675 585
R1726 B.n677 B.n676 585
R1727 B.n273 B.n272 585
R1728 B.n278 B.n273 585
R1729 B.n685 B.n684 585
R1730 B.n684 B.n683 585
R1731 B.n686 B.n271 585
R1732 B.n271 B.n270 585
R1733 B.n688 B.n687 585
R1734 B.n689 B.n688 585
R1735 B.n265 B.n264 585
R1736 B.n266 B.n265 585
R1737 B.n697 B.n696 585
R1738 B.n696 B.n695 585
R1739 B.n698 B.n263 585
R1740 B.n263 B.n262 585
R1741 B.n700 B.n699 585
R1742 B.n701 B.n700 585
R1743 B.n257 B.n256 585
R1744 B.n258 B.n257 585
R1745 B.n709 B.n708 585
R1746 B.n708 B.n707 585
R1747 B.n710 B.n255 585
R1748 B.n255 B.n253 585
R1749 B.n712 B.n711 585
R1750 B.n713 B.n712 585
R1751 B.n249 B.n248 585
R1752 B.n254 B.n249 585
R1753 B.n721 B.n720 585
R1754 B.n720 B.n719 585
R1755 B.n722 B.n247 585
R1756 B.n247 B.n246 585
R1757 B.n724 B.n723 585
R1758 B.n725 B.n724 585
R1759 B.n241 B.n240 585
R1760 B.n242 B.n241 585
R1761 B.n733 B.n732 585
R1762 B.n732 B.n731 585
R1763 B.n734 B.n239 585
R1764 B.n239 B.n238 585
R1765 B.n736 B.n735 585
R1766 B.n737 B.n736 585
R1767 B.n233 B.n232 585
R1768 B.n234 B.n233 585
R1769 B.n745 B.n744 585
R1770 B.n744 B.n743 585
R1771 B.n746 B.n231 585
R1772 B.n231 B.n230 585
R1773 B.n748 B.n747 585
R1774 B.n749 B.n748 585
R1775 B.n225 B.n224 585
R1776 B.n226 B.n225 585
R1777 B.n757 B.n756 585
R1778 B.n756 B.n755 585
R1779 B.n758 B.n223 585
R1780 B.n223 B.n222 585
R1781 B.n760 B.n759 585
R1782 B.n761 B.n760 585
R1783 B.n217 B.n216 585
R1784 B.n218 B.n217 585
R1785 B.n769 B.n768 585
R1786 B.n768 B.n767 585
R1787 B.n770 B.n215 585
R1788 B.n215 B.n214 585
R1789 B.n772 B.n771 585
R1790 B.n773 B.n772 585
R1791 B.n209 B.n208 585
R1792 B.n210 B.n209 585
R1793 B.n781 B.n780 585
R1794 B.n780 B.n779 585
R1795 B.n782 B.n207 585
R1796 B.n207 B.n206 585
R1797 B.n784 B.n783 585
R1798 B.n785 B.n784 585
R1799 B.n201 B.n200 585
R1800 B.n202 B.n201 585
R1801 B.n793 B.n792 585
R1802 B.n792 B.n791 585
R1803 B.n794 B.n199 585
R1804 B.n199 B.n198 585
R1805 B.n796 B.n795 585
R1806 B.n797 B.n796 585
R1807 B.n193 B.n192 585
R1808 B.n194 B.n193 585
R1809 B.n806 B.n805 585
R1810 B.n805 B.n804 585
R1811 B.n807 B.n191 585
R1812 B.n191 B.n190 585
R1813 B.n809 B.n808 585
R1814 B.n810 B.n809 585
R1815 B.n3 B.n0 585
R1816 B.n4 B.n3 585
R1817 B.n1261 B.n1 585
R1818 B.n1262 B.n1261 585
R1819 B.n1260 B.n1259 585
R1820 B.n1260 B.n8 585
R1821 B.n1258 B.n9 585
R1822 B.n12 B.n9 585
R1823 B.n1257 B.n1256 585
R1824 B.n1256 B.n1255 585
R1825 B.n11 B.n10 585
R1826 B.n1254 B.n11 585
R1827 B.n1252 B.n1251 585
R1828 B.n1253 B.n1252 585
R1829 B.n1250 B.n17 585
R1830 B.n17 B.n16 585
R1831 B.n1249 B.n1248 585
R1832 B.n1248 B.n1247 585
R1833 B.n19 B.n18 585
R1834 B.n1246 B.n19 585
R1835 B.n1244 B.n1243 585
R1836 B.n1245 B.n1244 585
R1837 B.n1242 B.n24 585
R1838 B.n24 B.n23 585
R1839 B.n1241 B.n1240 585
R1840 B.n1240 B.n1239 585
R1841 B.n26 B.n25 585
R1842 B.n1238 B.n26 585
R1843 B.n1236 B.n1235 585
R1844 B.n1237 B.n1236 585
R1845 B.n1234 B.n31 585
R1846 B.n31 B.n30 585
R1847 B.n1233 B.n1232 585
R1848 B.n1232 B.n1231 585
R1849 B.n33 B.n32 585
R1850 B.n1230 B.n33 585
R1851 B.n1228 B.n1227 585
R1852 B.n1229 B.n1228 585
R1853 B.n1226 B.n38 585
R1854 B.n38 B.n37 585
R1855 B.n1225 B.n1224 585
R1856 B.n1224 B.n1223 585
R1857 B.n40 B.n39 585
R1858 B.n1222 B.n40 585
R1859 B.n1220 B.n1219 585
R1860 B.n1221 B.n1220 585
R1861 B.n1218 B.n45 585
R1862 B.n45 B.n44 585
R1863 B.n1217 B.n1216 585
R1864 B.n1216 B.n1215 585
R1865 B.n47 B.n46 585
R1866 B.n1214 B.n47 585
R1867 B.n1212 B.n1211 585
R1868 B.n1213 B.n1212 585
R1869 B.n1210 B.n52 585
R1870 B.n52 B.n51 585
R1871 B.n1209 B.n1208 585
R1872 B.n1208 B.n1207 585
R1873 B.n54 B.n53 585
R1874 B.n1206 B.n54 585
R1875 B.n1204 B.n1203 585
R1876 B.n1205 B.n1204 585
R1877 B.n1202 B.n59 585
R1878 B.n59 B.n58 585
R1879 B.n1201 B.n1200 585
R1880 B.n1200 B.n1199 585
R1881 B.n61 B.n60 585
R1882 B.n1198 B.n61 585
R1883 B.n1196 B.n1195 585
R1884 B.n1197 B.n1196 585
R1885 B.n1194 B.n66 585
R1886 B.n66 B.n65 585
R1887 B.n1193 B.n1192 585
R1888 B.n1192 B.n1191 585
R1889 B.n68 B.n67 585
R1890 B.n1190 B.n68 585
R1891 B.n1188 B.n1187 585
R1892 B.n1189 B.n1188 585
R1893 B.n1186 B.n73 585
R1894 B.n73 B.n72 585
R1895 B.n1185 B.n1184 585
R1896 B.n1184 B.n1183 585
R1897 B.n75 B.n74 585
R1898 B.n1182 B.n75 585
R1899 B.n1180 B.n1179 585
R1900 B.n1181 B.n1180 585
R1901 B.n1178 B.n80 585
R1902 B.n80 B.n79 585
R1903 B.n1177 B.n1176 585
R1904 B.n1176 B.n1175 585
R1905 B.n82 B.n81 585
R1906 B.n1174 B.n82 585
R1907 B.n1172 B.n1171 585
R1908 B.n1173 B.n1172 585
R1909 B.n1170 B.n87 585
R1910 B.n87 B.n86 585
R1911 B.n1169 B.n1168 585
R1912 B.n1168 B.n1167 585
R1913 B.n89 B.n88 585
R1914 B.n1166 B.n89 585
R1915 B.n1164 B.n1163 585
R1916 B.n1165 B.n1164 585
R1917 B.n1162 B.n94 585
R1918 B.n94 B.n93 585
R1919 B.n1161 B.n1160 585
R1920 B.n1160 B.n1159 585
R1921 B.n96 B.n95 585
R1922 B.n1158 B.n96 585
R1923 B.n1156 B.n1155 585
R1924 B.n1157 B.n1156 585
R1925 B.n1154 B.n101 585
R1926 B.n101 B.n100 585
R1927 B.n1153 B.n1152 585
R1928 B.n1152 B.n1151 585
R1929 B.n103 B.n102 585
R1930 B.n1150 B.n103 585
R1931 B.n1148 B.n1147 585
R1932 B.n1149 B.n1148 585
R1933 B.n1146 B.n108 585
R1934 B.n108 B.n107 585
R1935 B.n1145 B.n1144 585
R1936 B.n1144 B.n1143 585
R1937 B.n110 B.n109 585
R1938 B.n1142 B.n110 585
R1939 B.n1140 B.n1139 585
R1940 B.n1141 B.n1140 585
R1941 B.n1138 B.n115 585
R1942 B.n115 B.n114 585
R1943 B.n1137 B.n1136 585
R1944 B.n1136 B.n1135 585
R1945 B.n117 B.n116 585
R1946 B.n1134 B.n117 585
R1947 B.n1132 B.n1131 585
R1948 B.n1133 B.n1132 585
R1949 B.n1130 B.n122 585
R1950 B.n122 B.n121 585
R1951 B.n1129 B.n1128 585
R1952 B.n1128 B.n1127 585
R1953 B.n124 B.n123 585
R1954 B.n1126 B.n124 585
R1955 B.n1124 B.n1123 585
R1956 B.n1125 B.n1124 585
R1957 B.n1265 B.n1264 585
R1958 B.n1263 B.n2 585
R1959 B.n1124 B.n129 482.89
R1960 B.n905 B.n127 482.89
R1961 B.n606 B.n325 482.89
R1962 B.n604 B.n327 482.89
R1963 B.n162 B.t14 412.058
R1964 B.n361 B.t18 412.058
R1965 B.n154 B.t20 412.058
R1966 B.n354 B.t11 412.058
R1967 B.n163 B.t15 330.022
R1968 B.n362 B.t17 330.022
R1969 B.n155 B.t21 330.022
R1970 B.n355 B.t10 330.022
R1971 B.n154 B.t19 300.752
R1972 B.n162 B.t12 300.752
R1973 B.n361 B.t16 300.752
R1974 B.n354 B.t8 300.752
R1975 B.n906 B.n128 256.663
R1976 B.n912 B.n128 256.663
R1977 B.n914 B.n128 256.663
R1978 B.n920 B.n128 256.663
R1979 B.n922 B.n128 256.663
R1980 B.n928 B.n128 256.663
R1981 B.n930 B.n128 256.663
R1982 B.n936 B.n128 256.663
R1983 B.n938 B.n128 256.663
R1984 B.n944 B.n128 256.663
R1985 B.n946 B.n128 256.663
R1986 B.n952 B.n128 256.663
R1987 B.n954 B.n128 256.663
R1988 B.n960 B.n128 256.663
R1989 B.n962 B.n128 256.663
R1990 B.n968 B.n128 256.663
R1991 B.n970 B.n128 256.663
R1992 B.n976 B.n128 256.663
R1993 B.n978 B.n128 256.663
R1994 B.n984 B.n128 256.663
R1995 B.n986 B.n128 256.663
R1996 B.n992 B.n128 256.663
R1997 B.n994 B.n128 256.663
R1998 B.n1000 B.n128 256.663
R1999 B.n1002 B.n128 256.663
R2000 B.n1009 B.n128 256.663
R2001 B.n1011 B.n128 256.663
R2002 B.n1017 B.n128 256.663
R2003 B.n157 B.n128 256.663
R2004 B.n1023 B.n128 256.663
R2005 B.n1029 B.n128 256.663
R2006 B.n1031 B.n128 256.663
R2007 B.n1037 B.n128 256.663
R2008 B.n1039 B.n128 256.663
R2009 B.n1045 B.n128 256.663
R2010 B.n1047 B.n128 256.663
R2011 B.n1053 B.n128 256.663
R2012 B.n1055 B.n128 256.663
R2013 B.n1061 B.n128 256.663
R2014 B.n1063 B.n128 256.663
R2015 B.n1069 B.n128 256.663
R2016 B.n1071 B.n128 256.663
R2017 B.n1077 B.n128 256.663
R2018 B.n1079 B.n128 256.663
R2019 B.n1085 B.n128 256.663
R2020 B.n1087 B.n128 256.663
R2021 B.n1093 B.n128 256.663
R2022 B.n1095 B.n128 256.663
R2023 B.n1101 B.n128 256.663
R2024 B.n1103 B.n128 256.663
R2025 B.n1109 B.n128 256.663
R2026 B.n1111 B.n128 256.663
R2027 B.n1117 B.n128 256.663
R2028 B.n1119 B.n128 256.663
R2029 B.n599 B.n326 256.663
R2030 B.n329 B.n326 256.663
R2031 B.n592 B.n326 256.663
R2032 B.n586 B.n326 256.663
R2033 B.n584 B.n326 256.663
R2034 B.n578 B.n326 256.663
R2035 B.n576 B.n326 256.663
R2036 B.n570 B.n326 256.663
R2037 B.n568 B.n326 256.663
R2038 B.n562 B.n326 256.663
R2039 B.n560 B.n326 256.663
R2040 B.n554 B.n326 256.663
R2041 B.n552 B.n326 256.663
R2042 B.n546 B.n326 256.663
R2043 B.n544 B.n326 256.663
R2044 B.n538 B.n326 256.663
R2045 B.n536 B.n326 256.663
R2046 B.n530 B.n326 256.663
R2047 B.n528 B.n326 256.663
R2048 B.n522 B.n326 256.663
R2049 B.n520 B.n326 256.663
R2050 B.n514 B.n326 256.663
R2051 B.n512 B.n326 256.663
R2052 B.n506 B.n326 256.663
R2053 B.n504 B.n326 256.663
R2054 B.n498 B.n326 256.663
R2055 B.n496 B.n326 256.663
R2056 B.n490 B.n326 256.663
R2057 B.n488 B.n326 256.663
R2058 B.n481 B.n326 256.663
R2059 B.n479 B.n326 256.663
R2060 B.n473 B.n326 256.663
R2061 B.n471 B.n326 256.663
R2062 B.n465 B.n326 256.663
R2063 B.n463 B.n326 256.663
R2064 B.n457 B.n326 256.663
R2065 B.n455 B.n326 256.663
R2066 B.n449 B.n326 256.663
R2067 B.n447 B.n326 256.663
R2068 B.n441 B.n326 256.663
R2069 B.n439 B.n326 256.663
R2070 B.n433 B.n326 256.663
R2071 B.n431 B.n326 256.663
R2072 B.n425 B.n326 256.663
R2073 B.n423 B.n326 256.663
R2074 B.n417 B.n326 256.663
R2075 B.n415 B.n326 256.663
R2076 B.n409 B.n326 256.663
R2077 B.n407 B.n326 256.663
R2078 B.n401 B.n326 256.663
R2079 B.n399 B.n326 256.663
R2080 B.n393 B.n326 256.663
R2081 B.n391 B.n326 256.663
R2082 B.n386 B.n326 256.663
R2083 B.n1267 B.n1266 256.663
R2084 B.n1120 B.n1118 163.367
R2085 B.n1116 B.n131 163.367
R2086 B.n1112 B.n1110 163.367
R2087 B.n1108 B.n133 163.367
R2088 B.n1104 B.n1102 163.367
R2089 B.n1100 B.n135 163.367
R2090 B.n1096 B.n1094 163.367
R2091 B.n1092 B.n137 163.367
R2092 B.n1088 B.n1086 163.367
R2093 B.n1084 B.n139 163.367
R2094 B.n1080 B.n1078 163.367
R2095 B.n1076 B.n141 163.367
R2096 B.n1072 B.n1070 163.367
R2097 B.n1068 B.n143 163.367
R2098 B.n1064 B.n1062 163.367
R2099 B.n1060 B.n145 163.367
R2100 B.n1056 B.n1054 163.367
R2101 B.n1052 B.n147 163.367
R2102 B.n1048 B.n1046 163.367
R2103 B.n1044 B.n149 163.367
R2104 B.n1040 B.n1038 163.367
R2105 B.n1036 B.n151 163.367
R2106 B.n1032 B.n1030 163.367
R2107 B.n1028 B.n153 163.367
R2108 B.n1024 B.n1022 163.367
R2109 B.n1019 B.n1018 163.367
R2110 B.n1016 B.n159 163.367
R2111 B.n1012 B.n1010 163.367
R2112 B.n1008 B.n161 163.367
R2113 B.n1003 B.n1001 163.367
R2114 B.n999 B.n165 163.367
R2115 B.n995 B.n993 163.367
R2116 B.n991 B.n167 163.367
R2117 B.n987 B.n985 163.367
R2118 B.n983 B.n169 163.367
R2119 B.n979 B.n977 163.367
R2120 B.n975 B.n171 163.367
R2121 B.n971 B.n969 163.367
R2122 B.n967 B.n173 163.367
R2123 B.n963 B.n961 163.367
R2124 B.n959 B.n175 163.367
R2125 B.n955 B.n953 163.367
R2126 B.n951 B.n177 163.367
R2127 B.n947 B.n945 163.367
R2128 B.n943 B.n179 163.367
R2129 B.n939 B.n937 163.367
R2130 B.n935 B.n181 163.367
R2131 B.n931 B.n929 163.367
R2132 B.n927 B.n183 163.367
R2133 B.n923 B.n921 163.367
R2134 B.n919 B.n185 163.367
R2135 B.n915 B.n913 163.367
R2136 B.n911 B.n187 163.367
R2137 B.n907 B.n905 163.367
R2138 B.n606 B.n323 163.367
R2139 B.n610 B.n323 163.367
R2140 B.n610 B.n317 163.367
R2141 B.n618 B.n317 163.367
R2142 B.n618 B.n315 163.367
R2143 B.n622 B.n315 163.367
R2144 B.n622 B.n308 163.367
R2145 B.n630 B.n308 163.367
R2146 B.n630 B.n306 163.367
R2147 B.n634 B.n306 163.367
R2148 B.n634 B.n301 163.367
R2149 B.n642 B.n301 163.367
R2150 B.n642 B.n299 163.367
R2151 B.n646 B.n299 163.367
R2152 B.n646 B.n293 163.367
R2153 B.n654 B.n293 163.367
R2154 B.n654 B.n291 163.367
R2155 B.n658 B.n291 163.367
R2156 B.n658 B.n285 163.367
R2157 B.n666 B.n285 163.367
R2158 B.n666 B.n283 163.367
R2159 B.n670 B.n283 163.367
R2160 B.n670 B.n276 163.367
R2161 B.n678 B.n276 163.367
R2162 B.n678 B.n274 163.367
R2163 B.n682 B.n274 163.367
R2164 B.n682 B.n269 163.367
R2165 B.n690 B.n269 163.367
R2166 B.n690 B.n267 163.367
R2167 B.n694 B.n267 163.367
R2168 B.n694 B.n261 163.367
R2169 B.n702 B.n261 163.367
R2170 B.n702 B.n259 163.367
R2171 B.n706 B.n259 163.367
R2172 B.n706 B.n252 163.367
R2173 B.n714 B.n252 163.367
R2174 B.n714 B.n250 163.367
R2175 B.n718 B.n250 163.367
R2176 B.n718 B.n245 163.367
R2177 B.n726 B.n245 163.367
R2178 B.n726 B.n243 163.367
R2179 B.n730 B.n243 163.367
R2180 B.n730 B.n237 163.367
R2181 B.n738 B.n237 163.367
R2182 B.n738 B.n235 163.367
R2183 B.n742 B.n235 163.367
R2184 B.n742 B.n229 163.367
R2185 B.n750 B.n229 163.367
R2186 B.n750 B.n227 163.367
R2187 B.n754 B.n227 163.367
R2188 B.n754 B.n221 163.367
R2189 B.n762 B.n221 163.367
R2190 B.n762 B.n219 163.367
R2191 B.n766 B.n219 163.367
R2192 B.n766 B.n213 163.367
R2193 B.n774 B.n213 163.367
R2194 B.n774 B.n211 163.367
R2195 B.n778 B.n211 163.367
R2196 B.n778 B.n205 163.367
R2197 B.n786 B.n205 163.367
R2198 B.n786 B.n203 163.367
R2199 B.n790 B.n203 163.367
R2200 B.n790 B.n197 163.367
R2201 B.n798 B.n197 163.367
R2202 B.n798 B.n195 163.367
R2203 B.n803 B.n195 163.367
R2204 B.n803 B.n189 163.367
R2205 B.n811 B.n189 163.367
R2206 B.n812 B.n811 163.367
R2207 B.n812 B.n5 163.367
R2208 B.n6 B.n5 163.367
R2209 B.n7 B.n6 163.367
R2210 B.n818 B.n7 163.367
R2211 B.n819 B.n818 163.367
R2212 B.n819 B.n13 163.367
R2213 B.n14 B.n13 163.367
R2214 B.n15 B.n14 163.367
R2215 B.n824 B.n15 163.367
R2216 B.n824 B.n20 163.367
R2217 B.n21 B.n20 163.367
R2218 B.n22 B.n21 163.367
R2219 B.n829 B.n22 163.367
R2220 B.n829 B.n27 163.367
R2221 B.n28 B.n27 163.367
R2222 B.n29 B.n28 163.367
R2223 B.n834 B.n29 163.367
R2224 B.n834 B.n34 163.367
R2225 B.n35 B.n34 163.367
R2226 B.n36 B.n35 163.367
R2227 B.n839 B.n36 163.367
R2228 B.n839 B.n41 163.367
R2229 B.n42 B.n41 163.367
R2230 B.n43 B.n42 163.367
R2231 B.n844 B.n43 163.367
R2232 B.n844 B.n48 163.367
R2233 B.n49 B.n48 163.367
R2234 B.n50 B.n49 163.367
R2235 B.n849 B.n50 163.367
R2236 B.n849 B.n55 163.367
R2237 B.n56 B.n55 163.367
R2238 B.n57 B.n56 163.367
R2239 B.n854 B.n57 163.367
R2240 B.n854 B.n62 163.367
R2241 B.n63 B.n62 163.367
R2242 B.n64 B.n63 163.367
R2243 B.n859 B.n64 163.367
R2244 B.n859 B.n69 163.367
R2245 B.n70 B.n69 163.367
R2246 B.n71 B.n70 163.367
R2247 B.n864 B.n71 163.367
R2248 B.n864 B.n76 163.367
R2249 B.n77 B.n76 163.367
R2250 B.n78 B.n77 163.367
R2251 B.n869 B.n78 163.367
R2252 B.n869 B.n83 163.367
R2253 B.n84 B.n83 163.367
R2254 B.n85 B.n84 163.367
R2255 B.n874 B.n85 163.367
R2256 B.n874 B.n90 163.367
R2257 B.n91 B.n90 163.367
R2258 B.n92 B.n91 163.367
R2259 B.n879 B.n92 163.367
R2260 B.n879 B.n97 163.367
R2261 B.n98 B.n97 163.367
R2262 B.n99 B.n98 163.367
R2263 B.n884 B.n99 163.367
R2264 B.n884 B.n104 163.367
R2265 B.n105 B.n104 163.367
R2266 B.n106 B.n105 163.367
R2267 B.n889 B.n106 163.367
R2268 B.n889 B.n111 163.367
R2269 B.n112 B.n111 163.367
R2270 B.n113 B.n112 163.367
R2271 B.n894 B.n113 163.367
R2272 B.n894 B.n118 163.367
R2273 B.n119 B.n118 163.367
R2274 B.n120 B.n119 163.367
R2275 B.n899 B.n120 163.367
R2276 B.n899 B.n125 163.367
R2277 B.n126 B.n125 163.367
R2278 B.n127 B.n126 163.367
R2279 B.n600 B.n598 163.367
R2280 B.n598 B.n597 163.367
R2281 B.n594 B.n593 163.367
R2282 B.n591 B.n331 163.367
R2283 B.n587 B.n585 163.367
R2284 B.n583 B.n333 163.367
R2285 B.n579 B.n577 163.367
R2286 B.n575 B.n335 163.367
R2287 B.n571 B.n569 163.367
R2288 B.n567 B.n337 163.367
R2289 B.n563 B.n561 163.367
R2290 B.n559 B.n339 163.367
R2291 B.n555 B.n553 163.367
R2292 B.n551 B.n341 163.367
R2293 B.n547 B.n545 163.367
R2294 B.n543 B.n343 163.367
R2295 B.n539 B.n537 163.367
R2296 B.n535 B.n345 163.367
R2297 B.n531 B.n529 163.367
R2298 B.n527 B.n347 163.367
R2299 B.n523 B.n521 163.367
R2300 B.n519 B.n349 163.367
R2301 B.n515 B.n513 163.367
R2302 B.n511 B.n351 163.367
R2303 B.n507 B.n505 163.367
R2304 B.n503 B.n353 163.367
R2305 B.n499 B.n497 163.367
R2306 B.n495 B.n358 163.367
R2307 B.n491 B.n489 163.367
R2308 B.n487 B.n360 163.367
R2309 B.n482 B.n480 163.367
R2310 B.n478 B.n364 163.367
R2311 B.n474 B.n472 163.367
R2312 B.n470 B.n366 163.367
R2313 B.n466 B.n464 163.367
R2314 B.n462 B.n368 163.367
R2315 B.n458 B.n456 163.367
R2316 B.n454 B.n370 163.367
R2317 B.n450 B.n448 163.367
R2318 B.n446 B.n372 163.367
R2319 B.n442 B.n440 163.367
R2320 B.n438 B.n374 163.367
R2321 B.n434 B.n432 163.367
R2322 B.n430 B.n376 163.367
R2323 B.n426 B.n424 163.367
R2324 B.n422 B.n378 163.367
R2325 B.n418 B.n416 163.367
R2326 B.n414 B.n380 163.367
R2327 B.n410 B.n408 163.367
R2328 B.n406 B.n382 163.367
R2329 B.n402 B.n400 163.367
R2330 B.n398 B.n384 163.367
R2331 B.n394 B.n392 163.367
R2332 B.n390 B.n387 163.367
R2333 B.n604 B.n321 163.367
R2334 B.n612 B.n321 163.367
R2335 B.n612 B.n319 163.367
R2336 B.n616 B.n319 163.367
R2337 B.n616 B.n313 163.367
R2338 B.n624 B.n313 163.367
R2339 B.n624 B.n311 163.367
R2340 B.n628 B.n311 163.367
R2341 B.n628 B.n305 163.367
R2342 B.n636 B.n305 163.367
R2343 B.n636 B.n303 163.367
R2344 B.n640 B.n303 163.367
R2345 B.n640 B.n297 163.367
R2346 B.n648 B.n297 163.367
R2347 B.n648 B.n295 163.367
R2348 B.n652 B.n295 163.367
R2349 B.n652 B.n289 163.367
R2350 B.n660 B.n289 163.367
R2351 B.n660 B.n287 163.367
R2352 B.n664 B.n287 163.367
R2353 B.n664 B.n281 163.367
R2354 B.n672 B.n281 163.367
R2355 B.n672 B.n279 163.367
R2356 B.n676 B.n279 163.367
R2357 B.n676 B.n273 163.367
R2358 B.n684 B.n273 163.367
R2359 B.n684 B.n271 163.367
R2360 B.n688 B.n271 163.367
R2361 B.n688 B.n265 163.367
R2362 B.n696 B.n265 163.367
R2363 B.n696 B.n263 163.367
R2364 B.n700 B.n263 163.367
R2365 B.n700 B.n257 163.367
R2366 B.n708 B.n257 163.367
R2367 B.n708 B.n255 163.367
R2368 B.n712 B.n255 163.367
R2369 B.n712 B.n249 163.367
R2370 B.n720 B.n249 163.367
R2371 B.n720 B.n247 163.367
R2372 B.n724 B.n247 163.367
R2373 B.n724 B.n241 163.367
R2374 B.n732 B.n241 163.367
R2375 B.n732 B.n239 163.367
R2376 B.n736 B.n239 163.367
R2377 B.n736 B.n233 163.367
R2378 B.n744 B.n233 163.367
R2379 B.n744 B.n231 163.367
R2380 B.n748 B.n231 163.367
R2381 B.n748 B.n225 163.367
R2382 B.n756 B.n225 163.367
R2383 B.n756 B.n223 163.367
R2384 B.n760 B.n223 163.367
R2385 B.n760 B.n217 163.367
R2386 B.n768 B.n217 163.367
R2387 B.n768 B.n215 163.367
R2388 B.n772 B.n215 163.367
R2389 B.n772 B.n209 163.367
R2390 B.n780 B.n209 163.367
R2391 B.n780 B.n207 163.367
R2392 B.n784 B.n207 163.367
R2393 B.n784 B.n201 163.367
R2394 B.n792 B.n201 163.367
R2395 B.n792 B.n199 163.367
R2396 B.n796 B.n199 163.367
R2397 B.n796 B.n193 163.367
R2398 B.n805 B.n193 163.367
R2399 B.n805 B.n191 163.367
R2400 B.n809 B.n191 163.367
R2401 B.n809 B.n3 163.367
R2402 B.n1265 B.n3 163.367
R2403 B.n1261 B.n2 163.367
R2404 B.n1261 B.n1260 163.367
R2405 B.n1260 B.n9 163.367
R2406 B.n1256 B.n9 163.367
R2407 B.n1256 B.n11 163.367
R2408 B.n1252 B.n11 163.367
R2409 B.n1252 B.n17 163.367
R2410 B.n1248 B.n17 163.367
R2411 B.n1248 B.n19 163.367
R2412 B.n1244 B.n19 163.367
R2413 B.n1244 B.n24 163.367
R2414 B.n1240 B.n24 163.367
R2415 B.n1240 B.n26 163.367
R2416 B.n1236 B.n26 163.367
R2417 B.n1236 B.n31 163.367
R2418 B.n1232 B.n31 163.367
R2419 B.n1232 B.n33 163.367
R2420 B.n1228 B.n33 163.367
R2421 B.n1228 B.n38 163.367
R2422 B.n1224 B.n38 163.367
R2423 B.n1224 B.n40 163.367
R2424 B.n1220 B.n40 163.367
R2425 B.n1220 B.n45 163.367
R2426 B.n1216 B.n45 163.367
R2427 B.n1216 B.n47 163.367
R2428 B.n1212 B.n47 163.367
R2429 B.n1212 B.n52 163.367
R2430 B.n1208 B.n52 163.367
R2431 B.n1208 B.n54 163.367
R2432 B.n1204 B.n54 163.367
R2433 B.n1204 B.n59 163.367
R2434 B.n1200 B.n59 163.367
R2435 B.n1200 B.n61 163.367
R2436 B.n1196 B.n61 163.367
R2437 B.n1196 B.n66 163.367
R2438 B.n1192 B.n66 163.367
R2439 B.n1192 B.n68 163.367
R2440 B.n1188 B.n68 163.367
R2441 B.n1188 B.n73 163.367
R2442 B.n1184 B.n73 163.367
R2443 B.n1184 B.n75 163.367
R2444 B.n1180 B.n75 163.367
R2445 B.n1180 B.n80 163.367
R2446 B.n1176 B.n80 163.367
R2447 B.n1176 B.n82 163.367
R2448 B.n1172 B.n82 163.367
R2449 B.n1172 B.n87 163.367
R2450 B.n1168 B.n87 163.367
R2451 B.n1168 B.n89 163.367
R2452 B.n1164 B.n89 163.367
R2453 B.n1164 B.n94 163.367
R2454 B.n1160 B.n94 163.367
R2455 B.n1160 B.n96 163.367
R2456 B.n1156 B.n96 163.367
R2457 B.n1156 B.n101 163.367
R2458 B.n1152 B.n101 163.367
R2459 B.n1152 B.n103 163.367
R2460 B.n1148 B.n103 163.367
R2461 B.n1148 B.n108 163.367
R2462 B.n1144 B.n108 163.367
R2463 B.n1144 B.n110 163.367
R2464 B.n1140 B.n110 163.367
R2465 B.n1140 B.n115 163.367
R2466 B.n1136 B.n115 163.367
R2467 B.n1136 B.n117 163.367
R2468 B.n1132 B.n117 163.367
R2469 B.n1132 B.n122 163.367
R2470 B.n1128 B.n122 163.367
R2471 B.n1128 B.n124 163.367
R2472 B.n1124 B.n124 163.367
R2473 B.n155 B.n154 82.0369
R2474 B.n163 B.n162 82.0369
R2475 B.n362 B.n361 82.0369
R2476 B.n355 B.n354 82.0369
R2477 B.n1119 B.n129 71.676
R2478 B.n1118 B.n1117 71.676
R2479 B.n1111 B.n131 71.676
R2480 B.n1110 B.n1109 71.676
R2481 B.n1103 B.n133 71.676
R2482 B.n1102 B.n1101 71.676
R2483 B.n1095 B.n135 71.676
R2484 B.n1094 B.n1093 71.676
R2485 B.n1087 B.n137 71.676
R2486 B.n1086 B.n1085 71.676
R2487 B.n1079 B.n139 71.676
R2488 B.n1078 B.n1077 71.676
R2489 B.n1071 B.n141 71.676
R2490 B.n1070 B.n1069 71.676
R2491 B.n1063 B.n143 71.676
R2492 B.n1062 B.n1061 71.676
R2493 B.n1055 B.n145 71.676
R2494 B.n1054 B.n1053 71.676
R2495 B.n1047 B.n147 71.676
R2496 B.n1046 B.n1045 71.676
R2497 B.n1039 B.n149 71.676
R2498 B.n1038 B.n1037 71.676
R2499 B.n1031 B.n151 71.676
R2500 B.n1030 B.n1029 71.676
R2501 B.n1023 B.n153 71.676
R2502 B.n1022 B.n157 71.676
R2503 B.n1018 B.n1017 71.676
R2504 B.n1011 B.n159 71.676
R2505 B.n1010 B.n1009 71.676
R2506 B.n1002 B.n161 71.676
R2507 B.n1001 B.n1000 71.676
R2508 B.n994 B.n165 71.676
R2509 B.n993 B.n992 71.676
R2510 B.n986 B.n167 71.676
R2511 B.n985 B.n984 71.676
R2512 B.n978 B.n169 71.676
R2513 B.n977 B.n976 71.676
R2514 B.n970 B.n171 71.676
R2515 B.n969 B.n968 71.676
R2516 B.n962 B.n173 71.676
R2517 B.n961 B.n960 71.676
R2518 B.n954 B.n175 71.676
R2519 B.n953 B.n952 71.676
R2520 B.n946 B.n177 71.676
R2521 B.n945 B.n944 71.676
R2522 B.n938 B.n179 71.676
R2523 B.n937 B.n936 71.676
R2524 B.n930 B.n181 71.676
R2525 B.n929 B.n928 71.676
R2526 B.n922 B.n183 71.676
R2527 B.n921 B.n920 71.676
R2528 B.n914 B.n185 71.676
R2529 B.n913 B.n912 71.676
R2530 B.n906 B.n187 71.676
R2531 B.n907 B.n906 71.676
R2532 B.n912 B.n911 71.676
R2533 B.n915 B.n914 71.676
R2534 B.n920 B.n919 71.676
R2535 B.n923 B.n922 71.676
R2536 B.n928 B.n927 71.676
R2537 B.n931 B.n930 71.676
R2538 B.n936 B.n935 71.676
R2539 B.n939 B.n938 71.676
R2540 B.n944 B.n943 71.676
R2541 B.n947 B.n946 71.676
R2542 B.n952 B.n951 71.676
R2543 B.n955 B.n954 71.676
R2544 B.n960 B.n959 71.676
R2545 B.n963 B.n962 71.676
R2546 B.n968 B.n967 71.676
R2547 B.n971 B.n970 71.676
R2548 B.n976 B.n975 71.676
R2549 B.n979 B.n978 71.676
R2550 B.n984 B.n983 71.676
R2551 B.n987 B.n986 71.676
R2552 B.n992 B.n991 71.676
R2553 B.n995 B.n994 71.676
R2554 B.n1000 B.n999 71.676
R2555 B.n1003 B.n1002 71.676
R2556 B.n1009 B.n1008 71.676
R2557 B.n1012 B.n1011 71.676
R2558 B.n1017 B.n1016 71.676
R2559 B.n1019 B.n157 71.676
R2560 B.n1024 B.n1023 71.676
R2561 B.n1029 B.n1028 71.676
R2562 B.n1032 B.n1031 71.676
R2563 B.n1037 B.n1036 71.676
R2564 B.n1040 B.n1039 71.676
R2565 B.n1045 B.n1044 71.676
R2566 B.n1048 B.n1047 71.676
R2567 B.n1053 B.n1052 71.676
R2568 B.n1056 B.n1055 71.676
R2569 B.n1061 B.n1060 71.676
R2570 B.n1064 B.n1063 71.676
R2571 B.n1069 B.n1068 71.676
R2572 B.n1072 B.n1071 71.676
R2573 B.n1077 B.n1076 71.676
R2574 B.n1080 B.n1079 71.676
R2575 B.n1085 B.n1084 71.676
R2576 B.n1088 B.n1087 71.676
R2577 B.n1093 B.n1092 71.676
R2578 B.n1096 B.n1095 71.676
R2579 B.n1101 B.n1100 71.676
R2580 B.n1104 B.n1103 71.676
R2581 B.n1109 B.n1108 71.676
R2582 B.n1112 B.n1111 71.676
R2583 B.n1117 B.n1116 71.676
R2584 B.n1120 B.n1119 71.676
R2585 B.n599 B.n327 71.676
R2586 B.n597 B.n329 71.676
R2587 B.n593 B.n592 71.676
R2588 B.n586 B.n331 71.676
R2589 B.n585 B.n584 71.676
R2590 B.n578 B.n333 71.676
R2591 B.n577 B.n576 71.676
R2592 B.n570 B.n335 71.676
R2593 B.n569 B.n568 71.676
R2594 B.n562 B.n337 71.676
R2595 B.n561 B.n560 71.676
R2596 B.n554 B.n339 71.676
R2597 B.n553 B.n552 71.676
R2598 B.n546 B.n341 71.676
R2599 B.n545 B.n544 71.676
R2600 B.n538 B.n343 71.676
R2601 B.n537 B.n536 71.676
R2602 B.n530 B.n345 71.676
R2603 B.n529 B.n528 71.676
R2604 B.n522 B.n347 71.676
R2605 B.n521 B.n520 71.676
R2606 B.n514 B.n349 71.676
R2607 B.n513 B.n512 71.676
R2608 B.n506 B.n351 71.676
R2609 B.n505 B.n504 71.676
R2610 B.n498 B.n353 71.676
R2611 B.n497 B.n496 71.676
R2612 B.n490 B.n358 71.676
R2613 B.n489 B.n488 71.676
R2614 B.n481 B.n360 71.676
R2615 B.n480 B.n479 71.676
R2616 B.n473 B.n364 71.676
R2617 B.n472 B.n471 71.676
R2618 B.n465 B.n366 71.676
R2619 B.n464 B.n463 71.676
R2620 B.n457 B.n368 71.676
R2621 B.n456 B.n455 71.676
R2622 B.n449 B.n370 71.676
R2623 B.n448 B.n447 71.676
R2624 B.n441 B.n372 71.676
R2625 B.n440 B.n439 71.676
R2626 B.n433 B.n374 71.676
R2627 B.n432 B.n431 71.676
R2628 B.n425 B.n376 71.676
R2629 B.n424 B.n423 71.676
R2630 B.n417 B.n378 71.676
R2631 B.n416 B.n415 71.676
R2632 B.n409 B.n380 71.676
R2633 B.n408 B.n407 71.676
R2634 B.n401 B.n382 71.676
R2635 B.n400 B.n399 71.676
R2636 B.n393 B.n384 71.676
R2637 B.n392 B.n391 71.676
R2638 B.n387 B.n386 71.676
R2639 B.n600 B.n599 71.676
R2640 B.n594 B.n329 71.676
R2641 B.n592 B.n591 71.676
R2642 B.n587 B.n586 71.676
R2643 B.n584 B.n583 71.676
R2644 B.n579 B.n578 71.676
R2645 B.n576 B.n575 71.676
R2646 B.n571 B.n570 71.676
R2647 B.n568 B.n567 71.676
R2648 B.n563 B.n562 71.676
R2649 B.n560 B.n559 71.676
R2650 B.n555 B.n554 71.676
R2651 B.n552 B.n551 71.676
R2652 B.n547 B.n546 71.676
R2653 B.n544 B.n543 71.676
R2654 B.n539 B.n538 71.676
R2655 B.n536 B.n535 71.676
R2656 B.n531 B.n530 71.676
R2657 B.n528 B.n527 71.676
R2658 B.n523 B.n522 71.676
R2659 B.n520 B.n519 71.676
R2660 B.n515 B.n514 71.676
R2661 B.n512 B.n511 71.676
R2662 B.n507 B.n506 71.676
R2663 B.n504 B.n503 71.676
R2664 B.n499 B.n498 71.676
R2665 B.n496 B.n495 71.676
R2666 B.n491 B.n490 71.676
R2667 B.n488 B.n487 71.676
R2668 B.n482 B.n481 71.676
R2669 B.n479 B.n478 71.676
R2670 B.n474 B.n473 71.676
R2671 B.n471 B.n470 71.676
R2672 B.n466 B.n465 71.676
R2673 B.n463 B.n462 71.676
R2674 B.n458 B.n457 71.676
R2675 B.n455 B.n454 71.676
R2676 B.n450 B.n449 71.676
R2677 B.n447 B.n446 71.676
R2678 B.n442 B.n441 71.676
R2679 B.n439 B.n438 71.676
R2680 B.n434 B.n433 71.676
R2681 B.n431 B.n430 71.676
R2682 B.n426 B.n425 71.676
R2683 B.n423 B.n422 71.676
R2684 B.n418 B.n417 71.676
R2685 B.n415 B.n414 71.676
R2686 B.n410 B.n409 71.676
R2687 B.n407 B.n406 71.676
R2688 B.n402 B.n401 71.676
R2689 B.n399 B.n398 71.676
R2690 B.n394 B.n393 71.676
R2691 B.n391 B.n390 71.676
R2692 B.n386 B.n325 71.676
R2693 B.n1266 B.n1265 71.676
R2694 B.n1266 B.n2 71.676
R2695 B.n605 B.n326 60.8831
R2696 B.n1125 B.n128 60.8831
R2697 B.n156 B.n155 59.5399
R2698 B.n1005 B.n163 59.5399
R2699 B.n485 B.n362 59.5399
R2700 B.n356 B.n355 59.5399
R2701 B.n605 B.n322 37.2979
R2702 B.n611 B.n322 37.2979
R2703 B.n611 B.n318 37.2979
R2704 B.n617 B.n318 37.2979
R2705 B.n617 B.n314 37.2979
R2706 B.n623 B.n314 37.2979
R2707 B.n623 B.n309 37.2979
R2708 B.n629 B.n309 37.2979
R2709 B.n629 B.n310 37.2979
R2710 B.n635 B.n302 37.2979
R2711 B.n641 B.n302 37.2979
R2712 B.n641 B.n298 37.2979
R2713 B.n647 B.n298 37.2979
R2714 B.n647 B.n294 37.2979
R2715 B.n653 B.n294 37.2979
R2716 B.n653 B.n290 37.2979
R2717 B.n659 B.n290 37.2979
R2718 B.n659 B.n286 37.2979
R2719 B.n665 B.n286 37.2979
R2720 B.n665 B.n282 37.2979
R2721 B.n671 B.n282 37.2979
R2722 B.n671 B.n277 37.2979
R2723 B.n677 B.n277 37.2979
R2724 B.n677 B.n278 37.2979
R2725 B.n683 B.n270 37.2979
R2726 B.n689 B.n270 37.2979
R2727 B.n689 B.n266 37.2979
R2728 B.n695 B.n266 37.2979
R2729 B.n695 B.n262 37.2979
R2730 B.n701 B.n262 37.2979
R2731 B.n701 B.n258 37.2979
R2732 B.n707 B.n258 37.2979
R2733 B.n707 B.n253 37.2979
R2734 B.n713 B.n253 37.2979
R2735 B.n713 B.n254 37.2979
R2736 B.n719 B.n246 37.2979
R2737 B.n725 B.n246 37.2979
R2738 B.n725 B.n242 37.2979
R2739 B.n731 B.n242 37.2979
R2740 B.n731 B.n238 37.2979
R2741 B.n737 B.n238 37.2979
R2742 B.n737 B.n234 37.2979
R2743 B.n743 B.n234 37.2979
R2744 B.n743 B.n230 37.2979
R2745 B.n749 B.n230 37.2979
R2746 B.n749 B.n226 37.2979
R2747 B.n755 B.n226 37.2979
R2748 B.n761 B.n222 37.2979
R2749 B.n761 B.n218 37.2979
R2750 B.n767 B.n218 37.2979
R2751 B.n767 B.n214 37.2979
R2752 B.n773 B.n214 37.2979
R2753 B.n773 B.n210 37.2979
R2754 B.n779 B.n210 37.2979
R2755 B.n779 B.n206 37.2979
R2756 B.n785 B.n206 37.2979
R2757 B.n785 B.n202 37.2979
R2758 B.n791 B.n202 37.2979
R2759 B.n797 B.n198 37.2979
R2760 B.n797 B.n194 37.2979
R2761 B.n804 B.n194 37.2979
R2762 B.n804 B.n190 37.2979
R2763 B.n810 B.n190 37.2979
R2764 B.n810 B.n4 37.2979
R2765 B.n1264 B.n4 37.2979
R2766 B.n1264 B.n1263 37.2979
R2767 B.n1263 B.n1262 37.2979
R2768 B.n1262 B.n8 37.2979
R2769 B.n12 B.n8 37.2979
R2770 B.n1255 B.n12 37.2979
R2771 B.n1255 B.n1254 37.2979
R2772 B.n1254 B.n1253 37.2979
R2773 B.n1253 B.n16 37.2979
R2774 B.n1247 B.n1246 37.2979
R2775 B.n1246 B.n1245 37.2979
R2776 B.n1245 B.n23 37.2979
R2777 B.n1239 B.n23 37.2979
R2778 B.n1239 B.n1238 37.2979
R2779 B.n1238 B.n1237 37.2979
R2780 B.n1237 B.n30 37.2979
R2781 B.n1231 B.n30 37.2979
R2782 B.n1231 B.n1230 37.2979
R2783 B.n1230 B.n1229 37.2979
R2784 B.n1229 B.n37 37.2979
R2785 B.n1223 B.n1222 37.2979
R2786 B.n1222 B.n1221 37.2979
R2787 B.n1221 B.n44 37.2979
R2788 B.n1215 B.n44 37.2979
R2789 B.n1215 B.n1214 37.2979
R2790 B.n1214 B.n1213 37.2979
R2791 B.n1213 B.n51 37.2979
R2792 B.n1207 B.n51 37.2979
R2793 B.n1207 B.n1206 37.2979
R2794 B.n1206 B.n1205 37.2979
R2795 B.n1205 B.n58 37.2979
R2796 B.n1199 B.n58 37.2979
R2797 B.n1198 B.n1197 37.2979
R2798 B.n1197 B.n65 37.2979
R2799 B.n1191 B.n65 37.2979
R2800 B.n1191 B.n1190 37.2979
R2801 B.n1190 B.n1189 37.2979
R2802 B.n1189 B.n72 37.2979
R2803 B.n1183 B.n72 37.2979
R2804 B.n1183 B.n1182 37.2979
R2805 B.n1182 B.n1181 37.2979
R2806 B.n1181 B.n79 37.2979
R2807 B.n1175 B.n79 37.2979
R2808 B.n1174 B.n1173 37.2979
R2809 B.n1173 B.n86 37.2979
R2810 B.n1167 B.n86 37.2979
R2811 B.n1167 B.n1166 37.2979
R2812 B.n1166 B.n1165 37.2979
R2813 B.n1165 B.n93 37.2979
R2814 B.n1159 B.n93 37.2979
R2815 B.n1159 B.n1158 37.2979
R2816 B.n1158 B.n1157 37.2979
R2817 B.n1157 B.n100 37.2979
R2818 B.n1151 B.n100 37.2979
R2819 B.n1151 B.n1150 37.2979
R2820 B.n1150 B.n1149 37.2979
R2821 B.n1149 B.n107 37.2979
R2822 B.n1143 B.n107 37.2979
R2823 B.n1142 B.n1141 37.2979
R2824 B.n1141 B.n114 37.2979
R2825 B.n1135 B.n114 37.2979
R2826 B.n1135 B.n1134 37.2979
R2827 B.n1134 B.n1133 37.2979
R2828 B.n1133 B.n121 37.2979
R2829 B.n1127 B.n121 37.2979
R2830 B.n1127 B.n1126 37.2979
R2831 B.n1126 B.n1125 37.2979
R2832 B.n603 B.n602 31.3761
R2833 B.n607 B.n324 31.3761
R2834 B.n904 B.n903 31.3761
R2835 B.n1123 B.n1122 31.3761
R2836 B.n254 B.t2 29.619
R2837 B.t4 B.n1198 29.619
R2838 B.t6 B.n222 28.5221
R2839 B.t7 B.n37 28.5221
R2840 B.n310 B.t9 26.3281
R2841 B.t13 B.n1142 26.3281
R2842 B.n791 B.t5 25.2311
R2843 B.n1247 B.t3 25.2311
R2844 B.n683 B.t0 24.1341
R2845 B.n1175 B.t1 24.1341
R2846 B B.n1267 18.0485
R2847 B.n278 B.t0 13.1643
R2848 B.t1 B.n1174 13.1643
R2849 B.t5 B.n198 12.0673
R2850 B.t3 B.n16 12.0673
R2851 B.n635 B.t9 10.9703
R2852 B.n1143 B.t13 10.9703
R2853 B.n603 B.n320 10.6151
R2854 B.n613 B.n320 10.6151
R2855 B.n614 B.n613 10.6151
R2856 B.n615 B.n614 10.6151
R2857 B.n615 B.n312 10.6151
R2858 B.n625 B.n312 10.6151
R2859 B.n626 B.n625 10.6151
R2860 B.n627 B.n626 10.6151
R2861 B.n627 B.n304 10.6151
R2862 B.n637 B.n304 10.6151
R2863 B.n638 B.n637 10.6151
R2864 B.n639 B.n638 10.6151
R2865 B.n639 B.n296 10.6151
R2866 B.n649 B.n296 10.6151
R2867 B.n650 B.n649 10.6151
R2868 B.n651 B.n650 10.6151
R2869 B.n651 B.n288 10.6151
R2870 B.n661 B.n288 10.6151
R2871 B.n662 B.n661 10.6151
R2872 B.n663 B.n662 10.6151
R2873 B.n663 B.n280 10.6151
R2874 B.n673 B.n280 10.6151
R2875 B.n674 B.n673 10.6151
R2876 B.n675 B.n674 10.6151
R2877 B.n675 B.n272 10.6151
R2878 B.n685 B.n272 10.6151
R2879 B.n686 B.n685 10.6151
R2880 B.n687 B.n686 10.6151
R2881 B.n687 B.n264 10.6151
R2882 B.n697 B.n264 10.6151
R2883 B.n698 B.n697 10.6151
R2884 B.n699 B.n698 10.6151
R2885 B.n699 B.n256 10.6151
R2886 B.n709 B.n256 10.6151
R2887 B.n710 B.n709 10.6151
R2888 B.n711 B.n710 10.6151
R2889 B.n711 B.n248 10.6151
R2890 B.n721 B.n248 10.6151
R2891 B.n722 B.n721 10.6151
R2892 B.n723 B.n722 10.6151
R2893 B.n723 B.n240 10.6151
R2894 B.n733 B.n240 10.6151
R2895 B.n734 B.n733 10.6151
R2896 B.n735 B.n734 10.6151
R2897 B.n735 B.n232 10.6151
R2898 B.n745 B.n232 10.6151
R2899 B.n746 B.n745 10.6151
R2900 B.n747 B.n746 10.6151
R2901 B.n747 B.n224 10.6151
R2902 B.n757 B.n224 10.6151
R2903 B.n758 B.n757 10.6151
R2904 B.n759 B.n758 10.6151
R2905 B.n759 B.n216 10.6151
R2906 B.n769 B.n216 10.6151
R2907 B.n770 B.n769 10.6151
R2908 B.n771 B.n770 10.6151
R2909 B.n771 B.n208 10.6151
R2910 B.n781 B.n208 10.6151
R2911 B.n782 B.n781 10.6151
R2912 B.n783 B.n782 10.6151
R2913 B.n783 B.n200 10.6151
R2914 B.n793 B.n200 10.6151
R2915 B.n794 B.n793 10.6151
R2916 B.n795 B.n794 10.6151
R2917 B.n795 B.n192 10.6151
R2918 B.n806 B.n192 10.6151
R2919 B.n807 B.n806 10.6151
R2920 B.n808 B.n807 10.6151
R2921 B.n808 B.n0 10.6151
R2922 B.n602 B.n601 10.6151
R2923 B.n601 B.n328 10.6151
R2924 B.n596 B.n328 10.6151
R2925 B.n596 B.n595 10.6151
R2926 B.n595 B.n330 10.6151
R2927 B.n590 B.n330 10.6151
R2928 B.n590 B.n589 10.6151
R2929 B.n589 B.n588 10.6151
R2930 B.n588 B.n332 10.6151
R2931 B.n582 B.n332 10.6151
R2932 B.n582 B.n581 10.6151
R2933 B.n581 B.n580 10.6151
R2934 B.n580 B.n334 10.6151
R2935 B.n574 B.n334 10.6151
R2936 B.n574 B.n573 10.6151
R2937 B.n573 B.n572 10.6151
R2938 B.n572 B.n336 10.6151
R2939 B.n566 B.n336 10.6151
R2940 B.n566 B.n565 10.6151
R2941 B.n565 B.n564 10.6151
R2942 B.n564 B.n338 10.6151
R2943 B.n558 B.n338 10.6151
R2944 B.n558 B.n557 10.6151
R2945 B.n557 B.n556 10.6151
R2946 B.n556 B.n340 10.6151
R2947 B.n550 B.n340 10.6151
R2948 B.n550 B.n549 10.6151
R2949 B.n549 B.n548 10.6151
R2950 B.n548 B.n342 10.6151
R2951 B.n542 B.n342 10.6151
R2952 B.n542 B.n541 10.6151
R2953 B.n541 B.n540 10.6151
R2954 B.n540 B.n344 10.6151
R2955 B.n534 B.n344 10.6151
R2956 B.n534 B.n533 10.6151
R2957 B.n533 B.n532 10.6151
R2958 B.n532 B.n346 10.6151
R2959 B.n526 B.n346 10.6151
R2960 B.n526 B.n525 10.6151
R2961 B.n525 B.n524 10.6151
R2962 B.n524 B.n348 10.6151
R2963 B.n518 B.n348 10.6151
R2964 B.n518 B.n517 10.6151
R2965 B.n517 B.n516 10.6151
R2966 B.n516 B.n350 10.6151
R2967 B.n510 B.n350 10.6151
R2968 B.n510 B.n509 10.6151
R2969 B.n509 B.n508 10.6151
R2970 B.n508 B.n352 10.6151
R2971 B.n502 B.n501 10.6151
R2972 B.n501 B.n500 10.6151
R2973 B.n500 B.n357 10.6151
R2974 B.n494 B.n357 10.6151
R2975 B.n494 B.n493 10.6151
R2976 B.n493 B.n492 10.6151
R2977 B.n492 B.n359 10.6151
R2978 B.n486 B.n359 10.6151
R2979 B.n484 B.n483 10.6151
R2980 B.n483 B.n363 10.6151
R2981 B.n477 B.n363 10.6151
R2982 B.n477 B.n476 10.6151
R2983 B.n476 B.n475 10.6151
R2984 B.n475 B.n365 10.6151
R2985 B.n469 B.n365 10.6151
R2986 B.n469 B.n468 10.6151
R2987 B.n468 B.n467 10.6151
R2988 B.n467 B.n367 10.6151
R2989 B.n461 B.n367 10.6151
R2990 B.n461 B.n460 10.6151
R2991 B.n460 B.n459 10.6151
R2992 B.n459 B.n369 10.6151
R2993 B.n453 B.n369 10.6151
R2994 B.n453 B.n452 10.6151
R2995 B.n452 B.n451 10.6151
R2996 B.n451 B.n371 10.6151
R2997 B.n445 B.n371 10.6151
R2998 B.n445 B.n444 10.6151
R2999 B.n444 B.n443 10.6151
R3000 B.n443 B.n373 10.6151
R3001 B.n437 B.n373 10.6151
R3002 B.n437 B.n436 10.6151
R3003 B.n436 B.n435 10.6151
R3004 B.n435 B.n375 10.6151
R3005 B.n429 B.n375 10.6151
R3006 B.n429 B.n428 10.6151
R3007 B.n428 B.n427 10.6151
R3008 B.n427 B.n377 10.6151
R3009 B.n421 B.n377 10.6151
R3010 B.n421 B.n420 10.6151
R3011 B.n420 B.n419 10.6151
R3012 B.n419 B.n379 10.6151
R3013 B.n413 B.n379 10.6151
R3014 B.n413 B.n412 10.6151
R3015 B.n412 B.n411 10.6151
R3016 B.n411 B.n381 10.6151
R3017 B.n405 B.n381 10.6151
R3018 B.n405 B.n404 10.6151
R3019 B.n404 B.n403 10.6151
R3020 B.n403 B.n383 10.6151
R3021 B.n397 B.n383 10.6151
R3022 B.n397 B.n396 10.6151
R3023 B.n396 B.n395 10.6151
R3024 B.n395 B.n385 10.6151
R3025 B.n389 B.n385 10.6151
R3026 B.n389 B.n388 10.6151
R3027 B.n388 B.n324 10.6151
R3028 B.n608 B.n607 10.6151
R3029 B.n609 B.n608 10.6151
R3030 B.n609 B.n316 10.6151
R3031 B.n619 B.n316 10.6151
R3032 B.n620 B.n619 10.6151
R3033 B.n621 B.n620 10.6151
R3034 B.n621 B.n307 10.6151
R3035 B.n631 B.n307 10.6151
R3036 B.n632 B.n631 10.6151
R3037 B.n633 B.n632 10.6151
R3038 B.n633 B.n300 10.6151
R3039 B.n643 B.n300 10.6151
R3040 B.n644 B.n643 10.6151
R3041 B.n645 B.n644 10.6151
R3042 B.n645 B.n292 10.6151
R3043 B.n655 B.n292 10.6151
R3044 B.n656 B.n655 10.6151
R3045 B.n657 B.n656 10.6151
R3046 B.n657 B.n284 10.6151
R3047 B.n667 B.n284 10.6151
R3048 B.n668 B.n667 10.6151
R3049 B.n669 B.n668 10.6151
R3050 B.n669 B.n275 10.6151
R3051 B.n679 B.n275 10.6151
R3052 B.n680 B.n679 10.6151
R3053 B.n681 B.n680 10.6151
R3054 B.n681 B.n268 10.6151
R3055 B.n691 B.n268 10.6151
R3056 B.n692 B.n691 10.6151
R3057 B.n693 B.n692 10.6151
R3058 B.n693 B.n260 10.6151
R3059 B.n703 B.n260 10.6151
R3060 B.n704 B.n703 10.6151
R3061 B.n705 B.n704 10.6151
R3062 B.n705 B.n251 10.6151
R3063 B.n715 B.n251 10.6151
R3064 B.n716 B.n715 10.6151
R3065 B.n717 B.n716 10.6151
R3066 B.n717 B.n244 10.6151
R3067 B.n727 B.n244 10.6151
R3068 B.n728 B.n727 10.6151
R3069 B.n729 B.n728 10.6151
R3070 B.n729 B.n236 10.6151
R3071 B.n739 B.n236 10.6151
R3072 B.n740 B.n739 10.6151
R3073 B.n741 B.n740 10.6151
R3074 B.n741 B.n228 10.6151
R3075 B.n751 B.n228 10.6151
R3076 B.n752 B.n751 10.6151
R3077 B.n753 B.n752 10.6151
R3078 B.n753 B.n220 10.6151
R3079 B.n763 B.n220 10.6151
R3080 B.n764 B.n763 10.6151
R3081 B.n765 B.n764 10.6151
R3082 B.n765 B.n212 10.6151
R3083 B.n775 B.n212 10.6151
R3084 B.n776 B.n775 10.6151
R3085 B.n777 B.n776 10.6151
R3086 B.n777 B.n204 10.6151
R3087 B.n787 B.n204 10.6151
R3088 B.n788 B.n787 10.6151
R3089 B.n789 B.n788 10.6151
R3090 B.n789 B.n196 10.6151
R3091 B.n799 B.n196 10.6151
R3092 B.n800 B.n799 10.6151
R3093 B.n802 B.n800 10.6151
R3094 B.n802 B.n801 10.6151
R3095 B.n801 B.n188 10.6151
R3096 B.n813 B.n188 10.6151
R3097 B.n814 B.n813 10.6151
R3098 B.n815 B.n814 10.6151
R3099 B.n816 B.n815 10.6151
R3100 B.n817 B.n816 10.6151
R3101 B.n820 B.n817 10.6151
R3102 B.n821 B.n820 10.6151
R3103 B.n822 B.n821 10.6151
R3104 B.n823 B.n822 10.6151
R3105 B.n825 B.n823 10.6151
R3106 B.n826 B.n825 10.6151
R3107 B.n827 B.n826 10.6151
R3108 B.n828 B.n827 10.6151
R3109 B.n830 B.n828 10.6151
R3110 B.n831 B.n830 10.6151
R3111 B.n832 B.n831 10.6151
R3112 B.n833 B.n832 10.6151
R3113 B.n835 B.n833 10.6151
R3114 B.n836 B.n835 10.6151
R3115 B.n837 B.n836 10.6151
R3116 B.n838 B.n837 10.6151
R3117 B.n840 B.n838 10.6151
R3118 B.n841 B.n840 10.6151
R3119 B.n842 B.n841 10.6151
R3120 B.n843 B.n842 10.6151
R3121 B.n845 B.n843 10.6151
R3122 B.n846 B.n845 10.6151
R3123 B.n847 B.n846 10.6151
R3124 B.n848 B.n847 10.6151
R3125 B.n850 B.n848 10.6151
R3126 B.n851 B.n850 10.6151
R3127 B.n852 B.n851 10.6151
R3128 B.n853 B.n852 10.6151
R3129 B.n855 B.n853 10.6151
R3130 B.n856 B.n855 10.6151
R3131 B.n857 B.n856 10.6151
R3132 B.n858 B.n857 10.6151
R3133 B.n860 B.n858 10.6151
R3134 B.n861 B.n860 10.6151
R3135 B.n862 B.n861 10.6151
R3136 B.n863 B.n862 10.6151
R3137 B.n865 B.n863 10.6151
R3138 B.n866 B.n865 10.6151
R3139 B.n867 B.n866 10.6151
R3140 B.n868 B.n867 10.6151
R3141 B.n870 B.n868 10.6151
R3142 B.n871 B.n870 10.6151
R3143 B.n872 B.n871 10.6151
R3144 B.n873 B.n872 10.6151
R3145 B.n875 B.n873 10.6151
R3146 B.n876 B.n875 10.6151
R3147 B.n877 B.n876 10.6151
R3148 B.n878 B.n877 10.6151
R3149 B.n880 B.n878 10.6151
R3150 B.n881 B.n880 10.6151
R3151 B.n882 B.n881 10.6151
R3152 B.n883 B.n882 10.6151
R3153 B.n885 B.n883 10.6151
R3154 B.n886 B.n885 10.6151
R3155 B.n887 B.n886 10.6151
R3156 B.n888 B.n887 10.6151
R3157 B.n890 B.n888 10.6151
R3158 B.n891 B.n890 10.6151
R3159 B.n892 B.n891 10.6151
R3160 B.n893 B.n892 10.6151
R3161 B.n895 B.n893 10.6151
R3162 B.n896 B.n895 10.6151
R3163 B.n897 B.n896 10.6151
R3164 B.n898 B.n897 10.6151
R3165 B.n900 B.n898 10.6151
R3166 B.n901 B.n900 10.6151
R3167 B.n902 B.n901 10.6151
R3168 B.n903 B.n902 10.6151
R3169 B.n1259 B.n1 10.6151
R3170 B.n1259 B.n1258 10.6151
R3171 B.n1258 B.n1257 10.6151
R3172 B.n1257 B.n10 10.6151
R3173 B.n1251 B.n10 10.6151
R3174 B.n1251 B.n1250 10.6151
R3175 B.n1250 B.n1249 10.6151
R3176 B.n1249 B.n18 10.6151
R3177 B.n1243 B.n18 10.6151
R3178 B.n1243 B.n1242 10.6151
R3179 B.n1242 B.n1241 10.6151
R3180 B.n1241 B.n25 10.6151
R3181 B.n1235 B.n25 10.6151
R3182 B.n1235 B.n1234 10.6151
R3183 B.n1234 B.n1233 10.6151
R3184 B.n1233 B.n32 10.6151
R3185 B.n1227 B.n32 10.6151
R3186 B.n1227 B.n1226 10.6151
R3187 B.n1226 B.n1225 10.6151
R3188 B.n1225 B.n39 10.6151
R3189 B.n1219 B.n39 10.6151
R3190 B.n1219 B.n1218 10.6151
R3191 B.n1218 B.n1217 10.6151
R3192 B.n1217 B.n46 10.6151
R3193 B.n1211 B.n46 10.6151
R3194 B.n1211 B.n1210 10.6151
R3195 B.n1210 B.n1209 10.6151
R3196 B.n1209 B.n53 10.6151
R3197 B.n1203 B.n53 10.6151
R3198 B.n1203 B.n1202 10.6151
R3199 B.n1202 B.n1201 10.6151
R3200 B.n1201 B.n60 10.6151
R3201 B.n1195 B.n60 10.6151
R3202 B.n1195 B.n1194 10.6151
R3203 B.n1194 B.n1193 10.6151
R3204 B.n1193 B.n67 10.6151
R3205 B.n1187 B.n67 10.6151
R3206 B.n1187 B.n1186 10.6151
R3207 B.n1186 B.n1185 10.6151
R3208 B.n1185 B.n74 10.6151
R3209 B.n1179 B.n74 10.6151
R3210 B.n1179 B.n1178 10.6151
R3211 B.n1178 B.n1177 10.6151
R3212 B.n1177 B.n81 10.6151
R3213 B.n1171 B.n81 10.6151
R3214 B.n1171 B.n1170 10.6151
R3215 B.n1170 B.n1169 10.6151
R3216 B.n1169 B.n88 10.6151
R3217 B.n1163 B.n88 10.6151
R3218 B.n1163 B.n1162 10.6151
R3219 B.n1162 B.n1161 10.6151
R3220 B.n1161 B.n95 10.6151
R3221 B.n1155 B.n95 10.6151
R3222 B.n1155 B.n1154 10.6151
R3223 B.n1154 B.n1153 10.6151
R3224 B.n1153 B.n102 10.6151
R3225 B.n1147 B.n102 10.6151
R3226 B.n1147 B.n1146 10.6151
R3227 B.n1146 B.n1145 10.6151
R3228 B.n1145 B.n109 10.6151
R3229 B.n1139 B.n109 10.6151
R3230 B.n1139 B.n1138 10.6151
R3231 B.n1138 B.n1137 10.6151
R3232 B.n1137 B.n116 10.6151
R3233 B.n1131 B.n116 10.6151
R3234 B.n1131 B.n1130 10.6151
R3235 B.n1130 B.n1129 10.6151
R3236 B.n1129 B.n123 10.6151
R3237 B.n1123 B.n123 10.6151
R3238 B.n1122 B.n1121 10.6151
R3239 B.n1121 B.n130 10.6151
R3240 B.n1115 B.n130 10.6151
R3241 B.n1115 B.n1114 10.6151
R3242 B.n1114 B.n1113 10.6151
R3243 B.n1113 B.n132 10.6151
R3244 B.n1107 B.n132 10.6151
R3245 B.n1107 B.n1106 10.6151
R3246 B.n1106 B.n1105 10.6151
R3247 B.n1105 B.n134 10.6151
R3248 B.n1099 B.n134 10.6151
R3249 B.n1099 B.n1098 10.6151
R3250 B.n1098 B.n1097 10.6151
R3251 B.n1097 B.n136 10.6151
R3252 B.n1091 B.n136 10.6151
R3253 B.n1091 B.n1090 10.6151
R3254 B.n1090 B.n1089 10.6151
R3255 B.n1089 B.n138 10.6151
R3256 B.n1083 B.n138 10.6151
R3257 B.n1083 B.n1082 10.6151
R3258 B.n1082 B.n1081 10.6151
R3259 B.n1081 B.n140 10.6151
R3260 B.n1075 B.n140 10.6151
R3261 B.n1075 B.n1074 10.6151
R3262 B.n1074 B.n1073 10.6151
R3263 B.n1073 B.n142 10.6151
R3264 B.n1067 B.n142 10.6151
R3265 B.n1067 B.n1066 10.6151
R3266 B.n1066 B.n1065 10.6151
R3267 B.n1065 B.n144 10.6151
R3268 B.n1059 B.n144 10.6151
R3269 B.n1059 B.n1058 10.6151
R3270 B.n1058 B.n1057 10.6151
R3271 B.n1057 B.n146 10.6151
R3272 B.n1051 B.n146 10.6151
R3273 B.n1051 B.n1050 10.6151
R3274 B.n1050 B.n1049 10.6151
R3275 B.n1049 B.n148 10.6151
R3276 B.n1043 B.n148 10.6151
R3277 B.n1043 B.n1042 10.6151
R3278 B.n1042 B.n1041 10.6151
R3279 B.n1041 B.n150 10.6151
R3280 B.n1035 B.n150 10.6151
R3281 B.n1035 B.n1034 10.6151
R3282 B.n1034 B.n1033 10.6151
R3283 B.n1033 B.n152 10.6151
R3284 B.n1027 B.n152 10.6151
R3285 B.n1027 B.n1026 10.6151
R3286 B.n1026 B.n1025 10.6151
R3287 B.n1021 B.n1020 10.6151
R3288 B.n1020 B.n158 10.6151
R3289 B.n1015 B.n158 10.6151
R3290 B.n1015 B.n1014 10.6151
R3291 B.n1014 B.n1013 10.6151
R3292 B.n1013 B.n160 10.6151
R3293 B.n1007 B.n160 10.6151
R3294 B.n1007 B.n1006 10.6151
R3295 B.n1004 B.n164 10.6151
R3296 B.n998 B.n164 10.6151
R3297 B.n998 B.n997 10.6151
R3298 B.n997 B.n996 10.6151
R3299 B.n996 B.n166 10.6151
R3300 B.n990 B.n166 10.6151
R3301 B.n990 B.n989 10.6151
R3302 B.n989 B.n988 10.6151
R3303 B.n988 B.n168 10.6151
R3304 B.n982 B.n168 10.6151
R3305 B.n982 B.n981 10.6151
R3306 B.n981 B.n980 10.6151
R3307 B.n980 B.n170 10.6151
R3308 B.n974 B.n170 10.6151
R3309 B.n974 B.n973 10.6151
R3310 B.n973 B.n972 10.6151
R3311 B.n972 B.n172 10.6151
R3312 B.n966 B.n172 10.6151
R3313 B.n966 B.n965 10.6151
R3314 B.n965 B.n964 10.6151
R3315 B.n964 B.n174 10.6151
R3316 B.n958 B.n174 10.6151
R3317 B.n958 B.n957 10.6151
R3318 B.n957 B.n956 10.6151
R3319 B.n956 B.n176 10.6151
R3320 B.n950 B.n176 10.6151
R3321 B.n950 B.n949 10.6151
R3322 B.n949 B.n948 10.6151
R3323 B.n948 B.n178 10.6151
R3324 B.n942 B.n178 10.6151
R3325 B.n942 B.n941 10.6151
R3326 B.n941 B.n940 10.6151
R3327 B.n940 B.n180 10.6151
R3328 B.n934 B.n180 10.6151
R3329 B.n934 B.n933 10.6151
R3330 B.n933 B.n932 10.6151
R3331 B.n932 B.n182 10.6151
R3332 B.n926 B.n182 10.6151
R3333 B.n926 B.n925 10.6151
R3334 B.n925 B.n924 10.6151
R3335 B.n924 B.n184 10.6151
R3336 B.n918 B.n184 10.6151
R3337 B.n918 B.n917 10.6151
R3338 B.n917 B.n916 10.6151
R3339 B.n916 B.n186 10.6151
R3340 B.n910 B.n186 10.6151
R3341 B.n910 B.n909 10.6151
R3342 B.n909 B.n908 10.6151
R3343 B.n908 B.n904 10.6151
R3344 B.n755 B.t6 8.77637
R3345 B.n1223 B.t7 8.77637
R3346 B.n1267 B.n0 8.11757
R3347 B.n1267 B.n1 8.11757
R3348 B.n719 B.t2 7.67938
R3349 B.n1199 B.t4 7.67938
R3350 B.n502 B.n356 6.5566
R3351 B.n486 B.n485 6.5566
R3352 B.n1021 B.n156 6.5566
R3353 B.n1006 B.n1005 6.5566
R3354 B.n356 B.n352 4.05904
R3355 B.n485 B.n484 4.05904
R3356 B.n1025 B.n156 4.05904
R3357 B.n1005 B.n1004 4.05904
R3358 VN.n76 VN.n75 161.3
R3359 VN.n74 VN.n40 161.3
R3360 VN.n73 VN.n72 161.3
R3361 VN.n71 VN.n41 161.3
R3362 VN.n70 VN.n69 161.3
R3363 VN.n68 VN.n42 161.3
R3364 VN.n67 VN.n66 161.3
R3365 VN.n65 VN.n43 161.3
R3366 VN.n64 VN.n63 161.3
R3367 VN.n61 VN.n44 161.3
R3368 VN.n60 VN.n59 161.3
R3369 VN.n58 VN.n45 161.3
R3370 VN.n57 VN.n56 161.3
R3371 VN.n55 VN.n46 161.3
R3372 VN.n54 VN.n53 161.3
R3373 VN.n52 VN.n47 161.3
R3374 VN.n51 VN.n50 161.3
R3375 VN.n37 VN.n36 161.3
R3376 VN.n35 VN.n1 161.3
R3377 VN.n34 VN.n33 161.3
R3378 VN.n32 VN.n2 161.3
R3379 VN.n31 VN.n30 161.3
R3380 VN.n29 VN.n3 161.3
R3381 VN.n28 VN.n27 161.3
R3382 VN.n26 VN.n4 161.3
R3383 VN.n25 VN.n24 161.3
R3384 VN.n22 VN.n5 161.3
R3385 VN.n21 VN.n20 161.3
R3386 VN.n19 VN.n6 161.3
R3387 VN.n18 VN.n17 161.3
R3388 VN.n16 VN.n7 161.3
R3389 VN.n15 VN.n14 161.3
R3390 VN.n13 VN.n8 161.3
R3391 VN.n12 VN.n11 161.3
R3392 VN.n48 VN.t5 124.7
R3393 VN.n9 VN.t7 124.7
R3394 VN.n10 VN.t3 91.3333
R3395 VN.n23 VN.t6 91.3333
R3396 VN.n0 VN.t2 91.3333
R3397 VN.n49 VN.t1 91.3333
R3398 VN.n62 VN.t0 91.3333
R3399 VN.n39 VN.t4 91.3333
R3400 VN.n38 VN.n0 85.5731
R3401 VN.n77 VN.n39 85.5731
R3402 VN VN.n77 59.3542
R3403 VN.n49 VN.n48 57.3643
R3404 VN.n10 VN.n9 57.3643
R3405 VN.n17 VN.n16 56.5617
R3406 VN.n56 VN.n55 56.5617
R3407 VN.n30 VN.n29 42.5146
R3408 VN.n69 VN.n68 42.5146
R3409 VN.n30 VN.n2 38.6395
R3410 VN.n69 VN.n41 38.6395
R3411 VN.n11 VN.n8 24.5923
R3412 VN.n15 VN.n8 24.5923
R3413 VN.n16 VN.n15 24.5923
R3414 VN.n17 VN.n6 24.5923
R3415 VN.n21 VN.n6 24.5923
R3416 VN.n22 VN.n21 24.5923
R3417 VN.n24 VN.n4 24.5923
R3418 VN.n28 VN.n4 24.5923
R3419 VN.n29 VN.n28 24.5923
R3420 VN.n34 VN.n2 24.5923
R3421 VN.n35 VN.n34 24.5923
R3422 VN.n36 VN.n35 24.5923
R3423 VN.n55 VN.n54 24.5923
R3424 VN.n54 VN.n47 24.5923
R3425 VN.n50 VN.n47 24.5923
R3426 VN.n68 VN.n67 24.5923
R3427 VN.n67 VN.n43 24.5923
R3428 VN.n63 VN.n43 24.5923
R3429 VN.n61 VN.n60 24.5923
R3430 VN.n60 VN.n45 24.5923
R3431 VN.n56 VN.n45 24.5923
R3432 VN.n75 VN.n74 24.5923
R3433 VN.n74 VN.n73 24.5923
R3434 VN.n73 VN.n41 24.5923
R3435 VN.n11 VN.n10 17.9525
R3436 VN.n23 VN.n22 17.9525
R3437 VN.n50 VN.n49 17.9525
R3438 VN.n62 VN.n61 17.9525
R3439 VN.n24 VN.n23 6.6403
R3440 VN.n63 VN.n62 6.6403
R3441 VN.n36 VN.n0 4.67295
R3442 VN.n75 VN.n39 4.67295
R3443 VN.n51 VN.n48 2.41405
R3444 VN.n12 VN.n9 2.41405
R3445 VN.n77 VN.n76 0.354861
R3446 VN.n38 VN.n37 0.354861
R3447 VN VN.n38 0.267071
R3448 VN.n76 VN.n40 0.189894
R3449 VN.n72 VN.n40 0.189894
R3450 VN.n72 VN.n71 0.189894
R3451 VN.n71 VN.n70 0.189894
R3452 VN.n70 VN.n42 0.189894
R3453 VN.n66 VN.n42 0.189894
R3454 VN.n66 VN.n65 0.189894
R3455 VN.n65 VN.n64 0.189894
R3456 VN.n64 VN.n44 0.189894
R3457 VN.n59 VN.n44 0.189894
R3458 VN.n59 VN.n58 0.189894
R3459 VN.n58 VN.n57 0.189894
R3460 VN.n57 VN.n46 0.189894
R3461 VN.n53 VN.n46 0.189894
R3462 VN.n53 VN.n52 0.189894
R3463 VN.n52 VN.n51 0.189894
R3464 VN.n13 VN.n12 0.189894
R3465 VN.n14 VN.n13 0.189894
R3466 VN.n14 VN.n7 0.189894
R3467 VN.n18 VN.n7 0.189894
R3468 VN.n19 VN.n18 0.189894
R3469 VN.n20 VN.n19 0.189894
R3470 VN.n20 VN.n5 0.189894
R3471 VN.n25 VN.n5 0.189894
R3472 VN.n26 VN.n25 0.189894
R3473 VN.n27 VN.n26 0.189894
R3474 VN.n27 VN.n3 0.189894
R3475 VN.n31 VN.n3 0.189894
R3476 VN.n32 VN.n31 0.189894
R3477 VN.n33 VN.n32 0.189894
R3478 VN.n33 VN.n1 0.189894
R3479 VN.n37 VN.n1 0.189894
R3480 VDD2.n2 VDD2.n1 65.404
R3481 VDD2.n2 VDD2.n0 65.404
R3482 VDD2 VDD2.n5 65.4012
R3483 VDD2.n4 VDD2.n3 63.6362
R3484 VDD2.n4 VDD2.n2 52.8662
R3485 VDD2 VDD2.n4 1.88197
R3486 VDD2.n5 VDD2.t6 1.34015
R3487 VDD2.n5 VDD2.t2 1.34015
R3488 VDD2.n3 VDD2.t3 1.34015
R3489 VDD2.n3 VDD2.t7 1.34015
R3490 VDD2.n1 VDD2.t1 1.34015
R3491 VDD2.n1 VDD2.t5 1.34015
R3492 VDD2.n0 VDD2.t0 1.34015
R3493 VDD2.n0 VDD2.t4 1.34015
C0 VDD1 VTAIL 9.42897f
C1 VDD2 VN 11.3418f
C2 VP VN 9.757759f
C3 VDD2 VTAIL 9.49211f
C4 VDD1 VDD2 2.44979f
C5 VP VTAIL 12.042299f
C6 VDD1 VP 11.8437f
C7 VDD2 VP 0.657959f
C8 VN VTAIL 12.0282f
C9 VDD1 VN 0.154033f
C10 VDD2 B 6.896034f
C11 VDD1 B 7.47153f
C12 VTAIL B 13.043134f
C13 VN B 20.71874f
C14 VP B 19.368212f
C15 VDD2.t0 B 0.312484f
C16 VDD2.t4 B 0.312484f
C17 VDD2.n0 B 2.84444f
C18 VDD2.t1 B 0.312484f
C19 VDD2.t5 B 0.312484f
C20 VDD2.n1 B 2.84444f
C21 VDD2.n2 B 4.4925f
C22 VDD2.t3 B 0.312484f
C23 VDD2.t7 B 0.312484f
C24 VDD2.n3 B 2.8257f
C25 VDD2.n4 B 3.85996f
C26 VDD2.t6 B 0.312484f
C27 VDD2.t2 B 0.312484f
C28 VDD2.n5 B 2.84439f
C29 VN.t2 B 2.59472f
C30 VN.n0 B 0.964276f
C31 VN.n1 B 0.016433f
C32 VN.n2 B 0.032771f
C33 VN.n3 B 0.016433f
C34 VN.n4 B 0.030473f
C35 VN.n5 B 0.016433f
C36 VN.t6 B 2.59472f
C37 VN.n6 B 0.030473f
C38 VN.n7 B 0.016433f
C39 VN.n8 B 0.030473f
C40 VN.t7 B 2.87095f
C41 VN.n9 B 0.912371f
C42 VN.t3 B 2.59472f
C43 VN.n10 B 0.962666f
C44 VN.n11 B 0.026412f
C45 VN.n12 B 0.212392f
C46 VN.n13 B 0.016433f
C47 VN.n14 B 0.016433f
C48 VN.n15 B 0.030473f
C49 VN.n16 B 0.023888f
C50 VN.n17 B 0.023888f
C51 VN.n18 B 0.016433f
C52 VN.n19 B 0.016433f
C53 VN.n20 B 0.016433f
C54 VN.n21 B 0.030473f
C55 VN.n22 B 0.026412f
C56 VN.n23 B 0.899907f
C57 VN.n24 B 0.019491f
C58 VN.n25 B 0.016433f
C59 VN.n26 B 0.016433f
C60 VN.n27 B 0.016433f
C61 VN.n28 B 0.030473f
C62 VN.n29 B 0.032122f
C63 VN.n30 B 0.013356f
C64 VN.n31 B 0.016433f
C65 VN.n32 B 0.016433f
C66 VN.n33 B 0.016433f
C67 VN.n34 B 0.030473f
C68 VN.n35 B 0.030473f
C69 VN.n36 B 0.018288f
C70 VN.n37 B 0.026518f
C71 VN.n38 B 0.050407f
C72 VN.t4 B 2.59472f
C73 VN.n39 B 0.964276f
C74 VN.n40 B 0.016433f
C75 VN.n41 B 0.032771f
C76 VN.n42 B 0.016433f
C77 VN.n43 B 0.030473f
C78 VN.n44 B 0.016433f
C79 VN.t0 B 2.59472f
C80 VN.n45 B 0.030473f
C81 VN.n46 B 0.016433f
C82 VN.n47 B 0.030473f
C83 VN.t5 B 2.87095f
C84 VN.n48 B 0.912371f
C85 VN.t1 B 2.59472f
C86 VN.n49 B 0.962666f
C87 VN.n50 B 0.026412f
C88 VN.n51 B 0.212392f
C89 VN.n52 B 0.016433f
C90 VN.n53 B 0.016433f
C91 VN.n54 B 0.030473f
C92 VN.n55 B 0.023888f
C93 VN.n56 B 0.023888f
C94 VN.n57 B 0.016433f
C95 VN.n58 B 0.016433f
C96 VN.n59 B 0.016433f
C97 VN.n60 B 0.030473f
C98 VN.n61 B 0.026412f
C99 VN.n62 B 0.899907f
C100 VN.n63 B 0.019491f
C101 VN.n64 B 0.016433f
C102 VN.n65 B 0.016433f
C103 VN.n66 B 0.016433f
C104 VN.n67 B 0.030473f
C105 VN.n68 B 0.032122f
C106 VN.n69 B 0.013356f
C107 VN.n70 B 0.016433f
C108 VN.n71 B 0.016433f
C109 VN.n72 B 0.016433f
C110 VN.n73 B 0.030473f
C111 VN.n74 B 0.030473f
C112 VN.n75 B 0.018288f
C113 VN.n76 B 0.026518f
C114 VN.n77 B 1.19965f
C115 VDD1.t4 B 0.316523f
C116 VDD1.t7 B 0.316523f
C117 VDD1.n0 B 2.88268f
C118 VDD1.t0 B 0.316523f
C119 VDD1.t2 B 0.316523f
C120 VDD1.n1 B 2.88121f
C121 VDD1.t5 B 0.316523f
C122 VDD1.t1 B 0.316523f
C123 VDD1.n2 B 2.88121f
C124 VDD1.n3 B 4.60621f
C125 VDD1.t3 B 0.316523f
C126 VDD1.t6 B 0.316523f
C127 VDD1.n4 B 2.86222f
C128 VDD1.n5 B 3.94417f
C129 VTAIL.t7 B 0.232433f
C130 VTAIL.t4 B 0.232433f
C131 VTAIL.n0 B 2.04616f
C132 VTAIL.n1 B 0.426622f
C133 VTAIL.n2 B 0.027167f
C134 VTAIL.n3 B 0.019901f
C135 VTAIL.n4 B 0.010694f
C136 VTAIL.n5 B 0.025276f
C137 VTAIL.n6 B 0.011323f
C138 VTAIL.n7 B 0.019901f
C139 VTAIL.n8 B 0.010694f
C140 VTAIL.n9 B 0.025276f
C141 VTAIL.n10 B 0.011323f
C142 VTAIL.n11 B 0.019901f
C143 VTAIL.n12 B 0.010694f
C144 VTAIL.n13 B 0.025276f
C145 VTAIL.n14 B 0.011323f
C146 VTAIL.n15 B 0.019901f
C147 VTAIL.n16 B 0.010694f
C148 VTAIL.n17 B 0.025276f
C149 VTAIL.n18 B 0.011323f
C150 VTAIL.n19 B 0.019901f
C151 VTAIL.n20 B 0.010694f
C152 VTAIL.n21 B 0.025276f
C153 VTAIL.n22 B 0.011323f
C154 VTAIL.n23 B 0.019901f
C155 VTAIL.n24 B 0.010694f
C156 VTAIL.n25 B 0.025276f
C157 VTAIL.n26 B 0.011323f
C158 VTAIL.n27 B 0.128699f
C159 VTAIL.t3 B 0.041662f
C160 VTAIL.n28 B 0.018957f
C161 VTAIL.n29 B 0.014931f
C162 VTAIL.n30 B 0.010694f
C163 VTAIL.n31 B 1.2747f
C164 VTAIL.n32 B 0.019901f
C165 VTAIL.n33 B 0.010694f
C166 VTAIL.n34 B 0.011323f
C167 VTAIL.n35 B 0.025276f
C168 VTAIL.n36 B 0.025276f
C169 VTAIL.n37 B 0.011323f
C170 VTAIL.n38 B 0.010694f
C171 VTAIL.n39 B 0.019901f
C172 VTAIL.n40 B 0.019901f
C173 VTAIL.n41 B 0.010694f
C174 VTAIL.n42 B 0.011323f
C175 VTAIL.n43 B 0.025276f
C176 VTAIL.n44 B 0.025276f
C177 VTAIL.n45 B 0.011323f
C178 VTAIL.n46 B 0.010694f
C179 VTAIL.n47 B 0.019901f
C180 VTAIL.n48 B 0.019901f
C181 VTAIL.n49 B 0.010694f
C182 VTAIL.n50 B 0.011323f
C183 VTAIL.n51 B 0.025276f
C184 VTAIL.n52 B 0.025276f
C185 VTAIL.n53 B 0.011323f
C186 VTAIL.n54 B 0.010694f
C187 VTAIL.n55 B 0.019901f
C188 VTAIL.n56 B 0.019901f
C189 VTAIL.n57 B 0.010694f
C190 VTAIL.n58 B 0.011323f
C191 VTAIL.n59 B 0.025276f
C192 VTAIL.n60 B 0.025276f
C193 VTAIL.n61 B 0.011323f
C194 VTAIL.n62 B 0.010694f
C195 VTAIL.n63 B 0.019901f
C196 VTAIL.n64 B 0.019901f
C197 VTAIL.n65 B 0.010694f
C198 VTAIL.n66 B 0.011323f
C199 VTAIL.n67 B 0.025276f
C200 VTAIL.n68 B 0.025276f
C201 VTAIL.n69 B 0.025276f
C202 VTAIL.n70 B 0.011323f
C203 VTAIL.n71 B 0.010694f
C204 VTAIL.n72 B 0.019901f
C205 VTAIL.n73 B 0.019901f
C206 VTAIL.n74 B 0.010694f
C207 VTAIL.n75 B 0.011008f
C208 VTAIL.n76 B 0.011008f
C209 VTAIL.n77 B 0.025276f
C210 VTAIL.n78 B 0.053294f
C211 VTAIL.n79 B 0.011323f
C212 VTAIL.n80 B 0.010694f
C213 VTAIL.n81 B 0.049806f
C214 VTAIL.n82 B 0.029787f
C215 VTAIL.n83 B 0.28311f
C216 VTAIL.n84 B 0.027167f
C217 VTAIL.n85 B 0.019901f
C218 VTAIL.n86 B 0.010694f
C219 VTAIL.n87 B 0.025276f
C220 VTAIL.n88 B 0.011323f
C221 VTAIL.n89 B 0.019901f
C222 VTAIL.n90 B 0.010694f
C223 VTAIL.n91 B 0.025276f
C224 VTAIL.n92 B 0.011323f
C225 VTAIL.n93 B 0.019901f
C226 VTAIL.n94 B 0.010694f
C227 VTAIL.n95 B 0.025276f
C228 VTAIL.n96 B 0.011323f
C229 VTAIL.n97 B 0.019901f
C230 VTAIL.n98 B 0.010694f
C231 VTAIL.n99 B 0.025276f
C232 VTAIL.n100 B 0.011323f
C233 VTAIL.n101 B 0.019901f
C234 VTAIL.n102 B 0.010694f
C235 VTAIL.n103 B 0.025276f
C236 VTAIL.n104 B 0.011323f
C237 VTAIL.n105 B 0.019901f
C238 VTAIL.n106 B 0.010694f
C239 VTAIL.n107 B 0.025276f
C240 VTAIL.n108 B 0.011323f
C241 VTAIL.n109 B 0.128699f
C242 VTAIL.t13 B 0.041662f
C243 VTAIL.n110 B 0.018957f
C244 VTAIL.n111 B 0.014931f
C245 VTAIL.n112 B 0.010694f
C246 VTAIL.n113 B 1.2747f
C247 VTAIL.n114 B 0.019901f
C248 VTAIL.n115 B 0.010694f
C249 VTAIL.n116 B 0.011323f
C250 VTAIL.n117 B 0.025276f
C251 VTAIL.n118 B 0.025276f
C252 VTAIL.n119 B 0.011323f
C253 VTAIL.n120 B 0.010694f
C254 VTAIL.n121 B 0.019901f
C255 VTAIL.n122 B 0.019901f
C256 VTAIL.n123 B 0.010694f
C257 VTAIL.n124 B 0.011323f
C258 VTAIL.n125 B 0.025276f
C259 VTAIL.n126 B 0.025276f
C260 VTAIL.n127 B 0.011323f
C261 VTAIL.n128 B 0.010694f
C262 VTAIL.n129 B 0.019901f
C263 VTAIL.n130 B 0.019901f
C264 VTAIL.n131 B 0.010694f
C265 VTAIL.n132 B 0.011323f
C266 VTAIL.n133 B 0.025276f
C267 VTAIL.n134 B 0.025276f
C268 VTAIL.n135 B 0.011323f
C269 VTAIL.n136 B 0.010694f
C270 VTAIL.n137 B 0.019901f
C271 VTAIL.n138 B 0.019901f
C272 VTAIL.n139 B 0.010694f
C273 VTAIL.n140 B 0.011323f
C274 VTAIL.n141 B 0.025276f
C275 VTAIL.n142 B 0.025276f
C276 VTAIL.n143 B 0.011323f
C277 VTAIL.n144 B 0.010694f
C278 VTAIL.n145 B 0.019901f
C279 VTAIL.n146 B 0.019901f
C280 VTAIL.n147 B 0.010694f
C281 VTAIL.n148 B 0.011323f
C282 VTAIL.n149 B 0.025276f
C283 VTAIL.n150 B 0.025276f
C284 VTAIL.n151 B 0.025276f
C285 VTAIL.n152 B 0.011323f
C286 VTAIL.n153 B 0.010694f
C287 VTAIL.n154 B 0.019901f
C288 VTAIL.n155 B 0.019901f
C289 VTAIL.n156 B 0.010694f
C290 VTAIL.n157 B 0.011008f
C291 VTAIL.n158 B 0.011008f
C292 VTAIL.n159 B 0.025276f
C293 VTAIL.n160 B 0.053294f
C294 VTAIL.n161 B 0.011323f
C295 VTAIL.n162 B 0.010694f
C296 VTAIL.n163 B 0.049806f
C297 VTAIL.n164 B 0.029787f
C298 VTAIL.n165 B 0.28311f
C299 VTAIL.t11 B 0.232433f
C300 VTAIL.t8 B 0.232433f
C301 VTAIL.n166 B 2.04616f
C302 VTAIL.n167 B 0.656724f
C303 VTAIL.n168 B 0.027167f
C304 VTAIL.n169 B 0.019901f
C305 VTAIL.n170 B 0.010694f
C306 VTAIL.n171 B 0.025276f
C307 VTAIL.n172 B 0.011323f
C308 VTAIL.n173 B 0.019901f
C309 VTAIL.n174 B 0.010694f
C310 VTAIL.n175 B 0.025276f
C311 VTAIL.n176 B 0.011323f
C312 VTAIL.n177 B 0.019901f
C313 VTAIL.n178 B 0.010694f
C314 VTAIL.n179 B 0.025276f
C315 VTAIL.n180 B 0.011323f
C316 VTAIL.n181 B 0.019901f
C317 VTAIL.n182 B 0.010694f
C318 VTAIL.n183 B 0.025276f
C319 VTAIL.n184 B 0.011323f
C320 VTAIL.n185 B 0.019901f
C321 VTAIL.n186 B 0.010694f
C322 VTAIL.n187 B 0.025276f
C323 VTAIL.n188 B 0.011323f
C324 VTAIL.n189 B 0.019901f
C325 VTAIL.n190 B 0.010694f
C326 VTAIL.n191 B 0.025276f
C327 VTAIL.n192 B 0.011323f
C328 VTAIL.n193 B 0.128699f
C329 VTAIL.t14 B 0.041662f
C330 VTAIL.n194 B 0.018957f
C331 VTAIL.n195 B 0.014931f
C332 VTAIL.n196 B 0.010694f
C333 VTAIL.n197 B 1.2747f
C334 VTAIL.n198 B 0.019901f
C335 VTAIL.n199 B 0.010694f
C336 VTAIL.n200 B 0.011323f
C337 VTAIL.n201 B 0.025276f
C338 VTAIL.n202 B 0.025276f
C339 VTAIL.n203 B 0.011323f
C340 VTAIL.n204 B 0.010694f
C341 VTAIL.n205 B 0.019901f
C342 VTAIL.n206 B 0.019901f
C343 VTAIL.n207 B 0.010694f
C344 VTAIL.n208 B 0.011323f
C345 VTAIL.n209 B 0.025276f
C346 VTAIL.n210 B 0.025276f
C347 VTAIL.n211 B 0.011323f
C348 VTAIL.n212 B 0.010694f
C349 VTAIL.n213 B 0.019901f
C350 VTAIL.n214 B 0.019901f
C351 VTAIL.n215 B 0.010694f
C352 VTAIL.n216 B 0.011323f
C353 VTAIL.n217 B 0.025276f
C354 VTAIL.n218 B 0.025276f
C355 VTAIL.n219 B 0.011323f
C356 VTAIL.n220 B 0.010694f
C357 VTAIL.n221 B 0.019901f
C358 VTAIL.n222 B 0.019901f
C359 VTAIL.n223 B 0.010694f
C360 VTAIL.n224 B 0.011323f
C361 VTAIL.n225 B 0.025276f
C362 VTAIL.n226 B 0.025276f
C363 VTAIL.n227 B 0.011323f
C364 VTAIL.n228 B 0.010694f
C365 VTAIL.n229 B 0.019901f
C366 VTAIL.n230 B 0.019901f
C367 VTAIL.n231 B 0.010694f
C368 VTAIL.n232 B 0.011323f
C369 VTAIL.n233 B 0.025276f
C370 VTAIL.n234 B 0.025276f
C371 VTAIL.n235 B 0.025276f
C372 VTAIL.n236 B 0.011323f
C373 VTAIL.n237 B 0.010694f
C374 VTAIL.n238 B 0.019901f
C375 VTAIL.n239 B 0.019901f
C376 VTAIL.n240 B 0.010694f
C377 VTAIL.n241 B 0.011008f
C378 VTAIL.n242 B 0.011008f
C379 VTAIL.n243 B 0.025276f
C380 VTAIL.n244 B 0.053294f
C381 VTAIL.n245 B 0.011323f
C382 VTAIL.n246 B 0.010694f
C383 VTAIL.n247 B 0.049806f
C384 VTAIL.n248 B 0.029787f
C385 VTAIL.n249 B 1.57418f
C386 VTAIL.n250 B 0.027167f
C387 VTAIL.n251 B 0.019901f
C388 VTAIL.n252 B 0.010694f
C389 VTAIL.n253 B 0.025276f
C390 VTAIL.n254 B 0.011323f
C391 VTAIL.n255 B 0.019901f
C392 VTAIL.n256 B 0.010694f
C393 VTAIL.n257 B 0.025276f
C394 VTAIL.n258 B 0.025276f
C395 VTAIL.n259 B 0.011323f
C396 VTAIL.n260 B 0.019901f
C397 VTAIL.n261 B 0.010694f
C398 VTAIL.n262 B 0.025276f
C399 VTAIL.n263 B 0.011323f
C400 VTAIL.n264 B 0.019901f
C401 VTAIL.n265 B 0.010694f
C402 VTAIL.n266 B 0.025276f
C403 VTAIL.n267 B 0.011323f
C404 VTAIL.n268 B 0.019901f
C405 VTAIL.n269 B 0.010694f
C406 VTAIL.n270 B 0.025276f
C407 VTAIL.n271 B 0.011323f
C408 VTAIL.n272 B 0.019901f
C409 VTAIL.n273 B 0.010694f
C410 VTAIL.n274 B 0.025276f
C411 VTAIL.n275 B 0.011323f
C412 VTAIL.n276 B 0.128699f
C413 VTAIL.t0 B 0.041662f
C414 VTAIL.n277 B 0.018957f
C415 VTAIL.n278 B 0.014931f
C416 VTAIL.n279 B 0.010694f
C417 VTAIL.n280 B 1.2747f
C418 VTAIL.n281 B 0.019901f
C419 VTAIL.n282 B 0.010694f
C420 VTAIL.n283 B 0.011323f
C421 VTAIL.n284 B 0.025276f
C422 VTAIL.n285 B 0.025276f
C423 VTAIL.n286 B 0.011323f
C424 VTAIL.n287 B 0.010694f
C425 VTAIL.n288 B 0.019901f
C426 VTAIL.n289 B 0.019901f
C427 VTAIL.n290 B 0.010694f
C428 VTAIL.n291 B 0.011323f
C429 VTAIL.n292 B 0.025276f
C430 VTAIL.n293 B 0.025276f
C431 VTAIL.n294 B 0.011323f
C432 VTAIL.n295 B 0.010694f
C433 VTAIL.n296 B 0.019901f
C434 VTAIL.n297 B 0.019901f
C435 VTAIL.n298 B 0.010694f
C436 VTAIL.n299 B 0.011323f
C437 VTAIL.n300 B 0.025276f
C438 VTAIL.n301 B 0.025276f
C439 VTAIL.n302 B 0.011323f
C440 VTAIL.n303 B 0.010694f
C441 VTAIL.n304 B 0.019901f
C442 VTAIL.n305 B 0.019901f
C443 VTAIL.n306 B 0.010694f
C444 VTAIL.n307 B 0.011323f
C445 VTAIL.n308 B 0.025276f
C446 VTAIL.n309 B 0.025276f
C447 VTAIL.n310 B 0.011323f
C448 VTAIL.n311 B 0.010694f
C449 VTAIL.n312 B 0.019901f
C450 VTAIL.n313 B 0.019901f
C451 VTAIL.n314 B 0.010694f
C452 VTAIL.n315 B 0.011323f
C453 VTAIL.n316 B 0.025276f
C454 VTAIL.n317 B 0.025276f
C455 VTAIL.n318 B 0.011323f
C456 VTAIL.n319 B 0.010694f
C457 VTAIL.n320 B 0.019901f
C458 VTAIL.n321 B 0.019901f
C459 VTAIL.n322 B 0.010694f
C460 VTAIL.n323 B 0.011008f
C461 VTAIL.n324 B 0.011008f
C462 VTAIL.n325 B 0.025276f
C463 VTAIL.n326 B 0.053294f
C464 VTAIL.n327 B 0.011323f
C465 VTAIL.n328 B 0.010694f
C466 VTAIL.n329 B 0.049806f
C467 VTAIL.n330 B 0.029787f
C468 VTAIL.n331 B 1.57418f
C469 VTAIL.t2 B 0.232433f
C470 VTAIL.t6 B 0.232433f
C471 VTAIL.n332 B 2.04617f
C472 VTAIL.n333 B 0.656714f
C473 VTAIL.n334 B 0.027167f
C474 VTAIL.n335 B 0.019901f
C475 VTAIL.n336 B 0.010694f
C476 VTAIL.n337 B 0.025276f
C477 VTAIL.n338 B 0.011323f
C478 VTAIL.n339 B 0.019901f
C479 VTAIL.n340 B 0.010694f
C480 VTAIL.n341 B 0.025276f
C481 VTAIL.n342 B 0.025276f
C482 VTAIL.n343 B 0.011323f
C483 VTAIL.n344 B 0.019901f
C484 VTAIL.n345 B 0.010694f
C485 VTAIL.n346 B 0.025276f
C486 VTAIL.n347 B 0.011323f
C487 VTAIL.n348 B 0.019901f
C488 VTAIL.n349 B 0.010694f
C489 VTAIL.n350 B 0.025276f
C490 VTAIL.n351 B 0.011323f
C491 VTAIL.n352 B 0.019901f
C492 VTAIL.n353 B 0.010694f
C493 VTAIL.n354 B 0.025276f
C494 VTAIL.n355 B 0.011323f
C495 VTAIL.n356 B 0.019901f
C496 VTAIL.n357 B 0.010694f
C497 VTAIL.n358 B 0.025276f
C498 VTAIL.n359 B 0.011323f
C499 VTAIL.n360 B 0.128699f
C500 VTAIL.t5 B 0.041662f
C501 VTAIL.n361 B 0.018957f
C502 VTAIL.n362 B 0.014931f
C503 VTAIL.n363 B 0.010694f
C504 VTAIL.n364 B 1.2747f
C505 VTAIL.n365 B 0.019901f
C506 VTAIL.n366 B 0.010694f
C507 VTAIL.n367 B 0.011323f
C508 VTAIL.n368 B 0.025276f
C509 VTAIL.n369 B 0.025276f
C510 VTAIL.n370 B 0.011323f
C511 VTAIL.n371 B 0.010694f
C512 VTAIL.n372 B 0.019901f
C513 VTAIL.n373 B 0.019901f
C514 VTAIL.n374 B 0.010694f
C515 VTAIL.n375 B 0.011323f
C516 VTAIL.n376 B 0.025276f
C517 VTAIL.n377 B 0.025276f
C518 VTAIL.n378 B 0.011323f
C519 VTAIL.n379 B 0.010694f
C520 VTAIL.n380 B 0.019901f
C521 VTAIL.n381 B 0.019901f
C522 VTAIL.n382 B 0.010694f
C523 VTAIL.n383 B 0.011323f
C524 VTAIL.n384 B 0.025276f
C525 VTAIL.n385 B 0.025276f
C526 VTAIL.n386 B 0.011323f
C527 VTAIL.n387 B 0.010694f
C528 VTAIL.n388 B 0.019901f
C529 VTAIL.n389 B 0.019901f
C530 VTAIL.n390 B 0.010694f
C531 VTAIL.n391 B 0.011323f
C532 VTAIL.n392 B 0.025276f
C533 VTAIL.n393 B 0.025276f
C534 VTAIL.n394 B 0.011323f
C535 VTAIL.n395 B 0.010694f
C536 VTAIL.n396 B 0.019901f
C537 VTAIL.n397 B 0.019901f
C538 VTAIL.n398 B 0.010694f
C539 VTAIL.n399 B 0.011323f
C540 VTAIL.n400 B 0.025276f
C541 VTAIL.n401 B 0.025276f
C542 VTAIL.n402 B 0.011323f
C543 VTAIL.n403 B 0.010694f
C544 VTAIL.n404 B 0.019901f
C545 VTAIL.n405 B 0.019901f
C546 VTAIL.n406 B 0.010694f
C547 VTAIL.n407 B 0.011008f
C548 VTAIL.n408 B 0.011008f
C549 VTAIL.n409 B 0.025276f
C550 VTAIL.n410 B 0.053294f
C551 VTAIL.n411 B 0.011323f
C552 VTAIL.n412 B 0.010694f
C553 VTAIL.n413 B 0.049806f
C554 VTAIL.n414 B 0.029787f
C555 VTAIL.n415 B 0.28311f
C556 VTAIL.n416 B 0.027167f
C557 VTAIL.n417 B 0.019901f
C558 VTAIL.n418 B 0.010694f
C559 VTAIL.n419 B 0.025276f
C560 VTAIL.n420 B 0.011323f
C561 VTAIL.n421 B 0.019901f
C562 VTAIL.n422 B 0.010694f
C563 VTAIL.n423 B 0.025276f
C564 VTAIL.n424 B 0.025276f
C565 VTAIL.n425 B 0.011323f
C566 VTAIL.n426 B 0.019901f
C567 VTAIL.n427 B 0.010694f
C568 VTAIL.n428 B 0.025276f
C569 VTAIL.n429 B 0.011323f
C570 VTAIL.n430 B 0.019901f
C571 VTAIL.n431 B 0.010694f
C572 VTAIL.n432 B 0.025276f
C573 VTAIL.n433 B 0.011323f
C574 VTAIL.n434 B 0.019901f
C575 VTAIL.n435 B 0.010694f
C576 VTAIL.n436 B 0.025276f
C577 VTAIL.n437 B 0.011323f
C578 VTAIL.n438 B 0.019901f
C579 VTAIL.n439 B 0.010694f
C580 VTAIL.n440 B 0.025276f
C581 VTAIL.n441 B 0.011323f
C582 VTAIL.n442 B 0.128699f
C583 VTAIL.t15 B 0.041662f
C584 VTAIL.n443 B 0.018957f
C585 VTAIL.n444 B 0.014931f
C586 VTAIL.n445 B 0.010694f
C587 VTAIL.n446 B 1.2747f
C588 VTAIL.n447 B 0.019901f
C589 VTAIL.n448 B 0.010694f
C590 VTAIL.n449 B 0.011323f
C591 VTAIL.n450 B 0.025276f
C592 VTAIL.n451 B 0.025276f
C593 VTAIL.n452 B 0.011323f
C594 VTAIL.n453 B 0.010694f
C595 VTAIL.n454 B 0.019901f
C596 VTAIL.n455 B 0.019901f
C597 VTAIL.n456 B 0.010694f
C598 VTAIL.n457 B 0.011323f
C599 VTAIL.n458 B 0.025276f
C600 VTAIL.n459 B 0.025276f
C601 VTAIL.n460 B 0.011323f
C602 VTAIL.n461 B 0.010694f
C603 VTAIL.n462 B 0.019901f
C604 VTAIL.n463 B 0.019901f
C605 VTAIL.n464 B 0.010694f
C606 VTAIL.n465 B 0.011323f
C607 VTAIL.n466 B 0.025276f
C608 VTAIL.n467 B 0.025276f
C609 VTAIL.n468 B 0.011323f
C610 VTAIL.n469 B 0.010694f
C611 VTAIL.n470 B 0.019901f
C612 VTAIL.n471 B 0.019901f
C613 VTAIL.n472 B 0.010694f
C614 VTAIL.n473 B 0.011323f
C615 VTAIL.n474 B 0.025276f
C616 VTAIL.n475 B 0.025276f
C617 VTAIL.n476 B 0.011323f
C618 VTAIL.n477 B 0.010694f
C619 VTAIL.n478 B 0.019901f
C620 VTAIL.n479 B 0.019901f
C621 VTAIL.n480 B 0.010694f
C622 VTAIL.n481 B 0.011323f
C623 VTAIL.n482 B 0.025276f
C624 VTAIL.n483 B 0.025276f
C625 VTAIL.n484 B 0.011323f
C626 VTAIL.n485 B 0.010694f
C627 VTAIL.n486 B 0.019901f
C628 VTAIL.n487 B 0.019901f
C629 VTAIL.n488 B 0.010694f
C630 VTAIL.n489 B 0.011008f
C631 VTAIL.n490 B 0.011008f
C632 VTAIL.n491 B 0.025276f
C633 VTAIL.n492 B 0.053294f
C634 VTAIL.n493 B 0.011323f
C635 VTAIL.n494 B 0.010694f
C636 VTAIL.n495 B 0.049806f
C637 VTAIL.n496 B 0.029787f
C638 VTAIL.n497 B 0.28311f
C639 VTAIL.t10 B 0.232433f
C640 VTAIL.t9 B 0.232433f
C641 VTAIL.n498 B 2.04617f
C642 VTAIL.n499 B 0.656714f
C643 VTAIL.n500 B 0.027167f
C644 VTAIL.n501 B 0.019901f
C645 VTAIL.n502 B 0.010694f
C646 VTAIL.n503 B 0.025276f
C647 VTAIL.n504 B 0.011323f
C648 VTAIL.n505 B 0.019901f
C649 VTAIL.n506 B 0.010694f
C650 VTAIL.n507 B 0.025276f
C651 VTAIL.n508 B 0.025276f
C652 VTAIL.n509 B 0.011323f
C653 VTAIL.n510 B 0.019901f
C654 VTAIL.n511 B 0.010694f
C655 VTAIL.n512 B 0.025276f
C656 VTAIL.n513 B 0.011323f
C657 VTAIL.n514 B 0.019901f
C658 VTAIL.n515 B 0.010694f
C659 VTAIL.n516 B 0.025276f
C660 VTAIL.n517 B 0.011323f
C661 VTAIL.n518 B 0.019901f
C662 VTAIL.n519 B 0.010694f
C663 VTAIL.n520 B 0.025276f
C664 VTAIL.n521 B 0.011323f
C665 VTAIL.n522 B 0.019901f
C666 VTAIL.n523 B 0.010694f
C667 VTAIL.n524 B 0.025276f
C668 VTAIL.n525 B 0.011323f
C669 VTAIL.n526 B 0.128699f
C670 VTAIL.t12 B 0.041662f
C671 VTAIL.n527 B 0.018957f
C672 VTAIL.n528 B 0.014931f
C673 VTAIL.n529 B 0.010694f
C674 VTAIL.n530 B 1.2747f
C675 VTAIL.n531 B 0.019901f
C676 VTAIL.n532 B 0.010694f
C677 VTAIL.n533 B 0.011323f
C678 VTAIL.n534 B 0.025276f
C679 VTAIL.n535 B 0.025276f
C680 VTAIL.n536 B 0.011323f
C681 VTAIL.n537 B 0.010694f
C682 VTAIL.n538 B 0.019901f
C683 VTAIL.n539 B 0.019901f
C684 VTAIL.n540 B 0.010694f
C685 VTAIL.n541 B 0.011323f
C686 VTAIL.n542 B 0.025276f
C687 VTAIL.n543 B 0.025276f
C688 VTAIL.n544 B 0.011323f
C689 VTAIL.n545 B 0.010694f
C690 VTAIL.n546 B 0.019901f
C691 VTAIL.n547 B 0.019901f
C692 VTAIL.n548 B 0.010694f
C693 VTAIL.n549 B 0.011323f
C694 VTAIL.n550 B 0.025276f
C695 VTAIL.n551 B 0.025276f
C696 VTAIL.n552 B 0.011323f
C697 VTAIL.n553 B 0.010694f
C698 VTAIL.n554 B 0.019901f
C699 VTAIL.n555 B 0.019901f
C700 VTAIL.n556 B 0.010694f
C701 VTAIL.n557 B 0.011323f
C702 VTAIL.n558 B 0.025276f
C703 VTAIL.n559 B 0.025276f
C704 VTAIL.n560 B 0.011323f
C705 VTAIL.n561 B 0.010694f
C706 VTAIL.n562 B 0.019901f
C707 VTAIL.n563 B 0.019901f
C708 VTAIL.n564 B 0.010694f
C709 VTAIL.n565 B 0.011323f
C710 VTAIL.n566 B 0.025276f
C711 VTAIL.n567 B 0.025276f
C712 VTAIL.n568 B 0.011323f
C713 VTAIL.n569 B 0.010694f
C714 VTAIL.n570 B 0.019901f
C715 VTAIL.n571 B 0.019901f
C716 VTAIL.n572 B 0.010694f
C717 VTAIL.n573 B 0.011008f
C718 VTAIL.n574 B 0.011008f
C719 VTAIL.n575 B 0.025276f
C720 VTAIL.n576 B 0.053294f
C721 VTAIL.n577 B 0.011323f
C722 VTAIL.n578 B 0.010694f
C723 VTAIL.n579 B 0.049806f
C724 VTAIL.n580 B 0.029787f
C725 VTAIL.n581 B 1.57418f
C726 VTAIL.n582 B 0.027167f
C727 VTAIL.n583 B 0.019901f
C728 VTAIL.n584 B 0.010694f
C729 VTAIL.n585 B 0.025276f
C730 VTAIL.n586 B 0.011323f
C731 VTAIL.n587 B 0.019901f
C732 VTAIL.n588 B 0.010694f
C733 VTAIL.n589 B 0.025276f
C734 VTAIL.n590 B 0.011323f
C735 VTAIL.n591 B 0.019901f
C736 VTAIL.n592 B 0.010694f
C737 VTAIL.n593 B 0.025276f
C738 VTAIL.n594 B 0.011323f
C739 VTAIL.n595 B 0.019901f
C740 VTAIL.n596 B 0.010694f
C741 VTAIL.n597 B 0.025276f
C742 VTAIL.n598 B 0.011323f
C743 VTAIL.n599 B 0.019901f
C744 VTAIL.n600 B 0.010694f
C745 VTAIL.n601 B 0.025276f
C746 VTAIL.n602 B 0.011323f
C747 VTAIL.n603 B 0.019901f
C748 VTAIL.n604 B 0.010694f
C749 VTAIL.n605 B 0.025276f
C750 VTAIL.n606 B 0.011323f
C751 VTAIL.n607 B 0.128699f
C752 VTAIL.t1 B 0.041662f
C753 VTAIL.n608 B 0.018957f
C754 VTAIL.n609 B 0.014931f
C755 VTAIL.n610 B 0.010694f
C756 VTAIL.n611 B 1.2747f
C757 VTAIL.n612 B 0.019901f
C758 VTAIL.n613 B 0.010694f
C759 VTAIL.n614 B 0.011323f
C760 VTAIL.n615 B 0.025276f
C761 VTAIL.n616 B 0.025276f
C762 VTAIL.n617 B 0.011323f
C763 VTAIL.n618 B 0.010694f
C764 VTAIL.n619 B 0.019901f
C765 VTAIL.n620 B 0.019901f
C766 VTAIL.n621 B 0.010694f
C767 VTAIL.n622 B 0.011323f
C768 VTAIL.n623 B 0.025276f
C769 VTAIL.n624 B 0.025276f
C770 VTAIL.n625 B 0.011323f
C771 VTAIL.n626 B 0.010694f
C772 VTAIL.n627 B 0.019901f
C773 VTAIL.n628 B 0.019901f
C774 VTAIL.n629 B 0.010694f
C775 VTAIL.n630 B 0.011323f
C776 VTAIL.n631 B 0.025276f
C777 VTAIL.n632 B 0.025276f
C778 VTAIL.n633 B 0.011323f
C779 VTAIL.n634 B 0.010694f
C780 VTAIL.n635 B 0.019901f
C781 VTAIL.n636 B 0.019901f
C782 VTAIL.n637 B 0.010694f
C783 VTAIL.n638 B 0.011323f
C784 VTAIL.n639 B 0.025276f
C785 VTAIL.n640 B 0.025276f
C786 VTAIL.n641 B 0.011323f
C787 VTAIL.n642 B 0.010694f
C788 VTAIL.n643 B 0.019901f
C789 VTAIL.n644 B 0.019901f
C790 VTAIL.n645 B 0.010694f
C791 VTAIL.n646 B 0.011323f
C792 VTAIL.n647 B 0.025276f
C793 VTAIL.n648 B 0.025276f
C794 VTAIL.n649 B 0.025276f
C795 VTAIL.n650 B 0.011323f
C796 VTAIL.n651 B 0.010694f
C797 VTAIL.n652 B 0.019901f
C798 VTAIL.n653 B 0.019901f
C799 VTAIL.n654 B 0.010694f
C800 VTAIL.n655 B 0.011008f
C801 VTAIL.n656 B 0.011008f
C802 VTAIL.n657 B 0.025276f
C803 VTAIL.n658 B 0.053294f
C804 VTAIL.n659 B 0.011323f
C805 VTAIL.n660 B 0.010694f
C806 VTAIL.n661 B 0.049806f
C807 VTAIL.n662 B 0.029787f
C808 VTAIL.n663 B 1.57045f
C809 VP.t6 B 2.63575f
C810 VP.n0 B 0.979526f
C811 VP.n1 B 0.016693f
C812 VP.n2 B 0.033289f
C813 VP.n3 B 0.016693f
C814 VP.n4 B 0.030956f
C815 VP.n5 B 0.016693f
C816 VP.t2 B 2.63575f
C817 VP.n6 B 0.030956f
C818 VP.n7 B 0.016693f
C819 VP.n8 B 0.030956f
C820 VP.n9 B 0.016693f
C821 VP.t5 B 2.63575f
C822 VP.n10 B 0.030956f
C823 VP.n11 B 0.016693f
C824 VP.n12 B 0.030956f
C825 VP.n13 B 0.026938f
C826 VP.t7 B 2.63575f
C827 VP.t1 B 2.63575f
C828 VP.n14 B 0.979526f
C829 VP.n15 B 0.016693f
C830 VP.n16 B 0.033289f
C831 VP.n17 B 0.016693f
C832 VP.n18 B 0.030956f
C833 VP.n19 B 0.016693f
C834 VP.t4 B 2.63575f
C835 VP.n20 B 0.030956f
C836 VP.n21 B 0.016693f
C837 VP.n22 B 0.030956f
C838 VP.t3 B 2.91635f
C839 VP.n23 B 0.926801f
C840 VP.t0 B 2.63575f
C841 VP.n24 B 0.97789f
C842 VP.n25 B 0.026829f
C843 VP.n26 B 0.215751f
C844 VP.n27 B 0.016693f
C845 VP.n28 B 0.016693f
C846 VP.n29 B 0.030956f
C847 VP.n30 B 0.024266f
C848 VP.n31 B 0.024266f
C849 VP.n32 B 0.016693f
C850 VP.n33 B 0.016693f
C851 VP.n34 B 0.016693f
C852 VP.n35 B 0.030956f
C853 VP.n36 B 0.026829f
C854 VP.n37 B 0.914139f
C855 VP.n38 B 0.0198f
C856 VP.n39 B 0.016693f
C857 VP.n40 B 0.016693f
C858 VP.n41 B 0.016693f
C859 VP.n42 B 0.030956f
C860 VP.n43 B 0.03263f
C861 VP.n44 B 0.013568f
C862 VP.n45 B 0.016693f
C863 VP.n46 B 0.016693f
C864 VP.n47 B 0.016693f
C865 VP.n48 B 0.030956f
C866 VP.n49 B 0.030956f
C867 VP.n50 B 0.018577f
C868 VP.n51 B 0.026938f
C869 VP.n52 B 1.21217f
C870 VP.n53 B 1.22234f
C871 VP.n54 B 0.979526f
C872 VP.n55 B 0.018577f
C873 VP.n56 B 0.030956f
C874 VP.n57 B 0.016693f
C875 VP.n58 B 0.016693f
C876 VP.n59 B 0.016693f
C877 VP.n60 B 0.033289f
C878 VP.n61 B 0.013568f
C879 VP.n62 B 0.03263f
C880 VP.n63 B 0.016693f
C881 VP.n64 B 0.016693f
C882 VP.n65 B 0.016693f
C883 VP.n66 B 0.030956f
C884 VP.n67 B 0.0198f
C885 VP.n68 B 0.914139f
C886 VP.n69 B 0.026829f
C887 VP.n70 B 0.016693f
C888 VP.n71 B 0.016693f
C889 VP.n72 B 0.016693f
C890 VP.n73 B 0.030956f
C891 VP.n74 B 0.024266f
C892 VP.n75 B 0.024266f
C893 VP.n76 B 0.016693f
C894 VP.n77 B 0.016693f
C895 VP.n78 B 0.016693f
C896 VP.n79 B 0.030956f
C897 VP.n80 B 0.026829f
C898 VP.n81 B 0.914139f
C899 VP.n82 B 0.0198f
C900 VP.n83 B 0.016693f
C901 VP.n84 B 0.016693f
C902 VP.n85 B 0.016693f
C903 VP.n86 B 0.030956f
C904 VP.n87 B 0.03263f
C905 VP.n88 B 0.013568f
C906 VP.n89 B 0.016693f
C907 VP.n90 B 0.016693f
C908 VP.n91 B 0.016693f
C909 VP.n92 B 0.030956f
C910 VP.n93 B 0.030956f
C911 VP.n94 B 0.018577f
C912 VP.n95 B 0.026938f
C913 VP.n96 B 0.051204f
.ends

