* NGSPICE file created from diff_pair_sample_0620.ext - technology: sky130A

.subckt diff_pair_sample_0620 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=5.2572 pd=27.74 as=0 ps=0 w=13.48 l=3.41
X1 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=5.2572 pd=27.74 as=0 ps=0 w=13.48 l=3.41
X2 VTAIL.t7 VN.t0 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=5.2572 pd=27.74 as=2.2242 ps=13.81 w=13.48 l=3.41
X3 VTAIL.t3 VP.t0 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=5.2572 pd=27.74 as=2.2242 ps=13.81 w=13.48 l=3.41
X4 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.2572 pd=27.74 as=0 ps=0 w=13.48 l=3.41
X5 VTAIL.t0 VP.t1 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=5.2572 pd=27.74 as=2.2242 ps=13.81 w=13.48 l=3.41
X6 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.2572 pd=27.74 as=0 ps=0 w=13.48 l=3.41
X7 VDD1.t1 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2242 pd=13.81 as=5.2572 ps=27.74 w=13.48 l=3.41
X8 VDD2.t1 VN.t1 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.2242 pd=13.81 as=5.2572 ps=27.74 w=13.48 l=3.41
X9 VDD1.t0 VP.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.2242 pd=13.81 as=5.2572 ps=27.74 w=13.48 l=3.41
X10 VTAIL.t5 VN.t2 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=5.2572 pd=27.74 as=2.2242 ps=13.81 w=13.48 l=3.41
X11 VDD2.t3 VN.t3 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.2242 pd=13.81 as=5.2572 ps=27.74 w=13.48 l=3.41
R0 B.n851 B.n850 585
R1 B.n334 B.n127 585
R2 B.n333 B.n332 585
R3 B.n331 B.n330 585
R4 B.n329 B.n328 585
R5 B.n327 B.n326 585
R6 B.n325 B.n324 585
R7 B.n323 B.n322 585
R8 B.n321 B.n320 585
R9 B.n319 B.n318 585
R10 B.n317 B.n316 585
R11 B.n315 B.n314 585
R12 B.n313 B.n312 585
R13 B.n311 B.n310 585
R14 B.n309 B.n308 585
R15 B.n307 B.n306 585
R16 B.n305 B.n304 585
R17 B.n303 B.n302 585
R18 B.n301 B.n300 585
R19 B.n299 B.n298 585
R20 B.n297 B.n296 585
R21 B.n295 B.n294 585
R22 B.n293 B.n292 585
R23 B.n291 B.n290 585
R24 B.n289 B.n288 585
R25 B.n287 B.n286 585
R26 B.n285 B.n284 585
R27 B.n283 B.n282 585
R28 B.n281 B.n280 585
R29 B.n279 B.n278 585
R30 B.n277 B.n276 585
R31 B.n275 B.n274 585
R32 B.n273 B.n272 585
R33 B.n271 B.n270 585
R34 B.n269 B.n268 585
R35 B.n267 B.n266 585
R36 B.n265 B.n264 585
R37 B.n263 B.n262 585
R38 B.n261 B.n260 585
R39 B.n259 B.n258 585
R40 B.n257 B.n256 585
R41 B.n255 B.n254 585
R42 B.n253 B.n252 585
R43 B.n251 B.n250 585
R44 B.n249 B.n248 585
R45 B.n247 B.n246 585
R46 B.n245 B.n244 585
R47 B.n243 B.n242 585
R48 B.n241 B.n240 585
R49 B.n239 B.n238 585
R50 B.n237 B.n236 585
R51 B.n235 B.n234 585
R52 B.n233 B.n232 585
R53 B.n231 B.n230 585
R54 B.n229 B.n228 585
R55 B.n227 B.n226 585
R56 B.n225 B.n224 585
R57 B.n223 B.n222 585
R58 B.n221 B.n220 585
R59 B.n219 B.n218 585
R60 B.n217 B.n216 585
R61 B.n215 B.n214 585
R62 B.n213 B.n212 585
R63 B.n211 B.n210 585
R64 B.n209 B.n208 585
R65 B.n207 B.n206 585
R66 B.n205 B.n204 585
R67 B.n203 B.n202 585
R68 B.n201 B.n200 585
R69 B.n199 B.n198 585
R70 B.n197 B.n196 585
R71 B.n195 B.n194 585
R72 B.n193 B.n192 585
R73 B.n191 B.n190 585
R74 B.n189 B.n188 585
R75 B.n187 B.n186 585
R76 B.n185 B.n184 585
R77 B.n183 B.n182 585
R78 B.n181 B.n180 585
R79 B.n179 B.n178 585
R80 B.n177 B.n176 585
R81 B.n175 B.n174 585
R82 B.n173 B.n172 585
R83 B.n171 B.n170 585
R84 B.n169 B.n168 585
R85 B.n167 B.n166 585
R86 B.n165 B.n164 585
R87 B.n163 B.n162 585
R88 B.n161 B.n160 585
R89 B.n159 B.n158 585
R90 B.n157 B.n156 585
R91 B.n155 B.n154 585
R92 B.n153 B.n152 585
R93 B.n151 B.n150 585
R94 B.n149 B.n148 585
R95 B.n147 B.n146 585
R96 B.n145 B.n144 585
R97 B.n143 B.n142 585
R98 B.n141 B.n140 585
R99 B.n139 B.n138 585
R100 B.n137 B.n136 585
R101 B.n135 B.n134 585
R102 B.n849 B.n76 585
R103 B.n854 B.n76 585
R104 B.n848 B.n75 585
R105 B.n855 B.n75 585
R106 B.n847 B.n846 585
R107 B.n846 B.n71 585
R108 B.n845 B.n70 585
R109 B.n861 B.n70 585
R110 B.n844 B.n69 585
R111 B.n862 B.n69 585
R112 B.n843 B.n68 585
R113 B.n863 B.n68 585
R114 B.n842 B.n841 585
R115 B.n841 B.n64 585
R116 B.n840 B.n63 585
R117 B.n869 B.n63 585
R118 B.n839 B.n62 585
R119 B.n870 B.n62 585
R120 B.n838 B.n61 585
R121 B.n871 B.n61 585
R122 B.n837 B.n836 585
R123 B.n836 B.n57 585
R124 B.n835 B.n56 585
R125 B.n877 B.n56 585
R126 B.n834 B.n55 585
R127 B.n878 B.n55 585
R128 B.n833 B.n54 585
R129 B.n879 B.n54 585
R130 B.n832 B.n831 585
R131 B.n831 B.n50 585
R132 B.n830 B.n49 585
R133 B.n885 B.n49 585
R134 B.n829 B.n48 585
R135 B.n886 B.n48 585
R136 B.n828 B.n47 585
R137 B.n887 B.n47 585
R138 B.n827 B.n826 585
R139 B.n826 B.n43 585
R140 B.n825 B.n42 585
R141 B.n893 B.n42 585
R142 B.n824 B.n41 585
R143 B.n894 B.n41 585
R144 B.n823 B.n40 585
R145 B.n895 B.n40 585
R146 B.n822 B.n821 585
R147 B.n821 B.n39 585
R148 B.n820 B.n35 585
R149 B.n901 B.n35 585
R150 B.n819 B.n34 585
R151 B.n902 B.n34 585
R152 B.n818 B.n33 585
R153 B.n903 B.n33 585
R154 B.n817 B.n816 585
R155 B.n816 B.n29 585
R156 B.n815 B.n28 585
R157 B.n909 B.n28 585
R158 B.n814 B.n27 585
R159 B.n910 B.n27 585
R160 B.n813 B.n26 585
R161 B.n911 B.n26 585
R162 B.n812 B.n811 585
R163 B.n811 B.n22 585
R164 B.n810 B.n21 585
R165 B.n917 B.n21 585
R166 B.n809 B.n20 585
R167 B.n918 B.n20 585
R168 B.n808 B.n19 585
R169 B.n919 B.n19 585
R170 B.n807 B.n806 585
R171 B.n806 B.n15 585
R172 B.n805 B.n14 585
R173 B.n925 B.n14 585
R174 B.n804 B.n13 585
R175 B.n926 B.n13 585
R176 B.n803 B.n12 585
R177 B.n927 B.n12 585
R178 B.n802 B.n801 585
R179 B.n801 B.n8 585
R180 B.n800 B.n7 585
R181 B.n933 B.n7 585
R182 B.n799 B.n6 585
R183 B.n934 B.n6 585
R184 B.n798 B.n5 585
R185 B.n935 B.n5 585
R186 B.n797 B.n796 585
R187 B.n796 B.n4 585
R188 B.n795 B.n335 585
R189 B.n795 B.n794 585
R190 B.n785 B.n336 585
R191 B.n337 B.n336 585
R192 B.n787 B.n786 585
R193 B.n788 B.n787 585
R194 B.n784 B.n342 585
R195 B.n342 B.n341 585
R196 B.n783 B.n782 585
R197 B.n782 B.n781 585
R198 B.n344 B.n343 585
R199 B.n345 B.n344 585
R200 B.n774 B.n773 585
R201 B.n775 B.n774 585
R202 B.n772 B.n350 585
R203 B.n350 B.n349 585
R204 B.n771 B.n770 585
R205 B.n770 B.n769 585
R206 B.n352 B.n351 585
R207 B.n353 B.n352 585
R208 B.n762 B.n761 585
R209 B.n763 B.n762 585
R210 B.n760 B.n358 585
R211 B.n358 B.n357 585
R212 B.n759 B.n758 585
R213 B.n758 B.n757 585
R214 B.n360 B.n359 585
R215 B.n361 B.n360 585
R216 B.n750 B.n749 585
R217 B.n751 B.n750 585
R218 B.n748 B.n366 585
R219 B.n366 B.n365 585
R220 B.n747 B.n746 585
R221 B.n746 B.n745 585
R222 B.n368 B.n367 585
R223 B.n738 B.n368 585
R224 B.n737 B.n736 585
R225 B.n739 B.n737 585
R226 B.n735 B.n373 585
R227 B.n373 B.n372 585
R228 B.n734 B.n733 585
R229 B.n733 B.n732 585
R230 B.n375 B.n374 585
R231 B.n376 B.n375 585
R232 B.n725 B.n724 585
R233 B.n726 B.n725 585
R234 B.n723 B.n381 585
R235 B.n381 B.n380 585
R236 B.n722 B.n721 585
R237 B.n721 B.n720 585
R238 B.n383 B.n382 585
R239 B.n384 B.n383 585
R240 B.n713 B.n712 585
R241 B.n714 B.n713 585
R242 B.n711 B.n389 585
R243 B.n389 B.n388 585
R244 B.n710 B.n709 585
R245 B.n709 B.n708 585
R246 B.n391 B.n390 585
R247 B.n392 B.n391 585
R248 B.n701 B.n700 585
R249 B.n702 B.n701 585
R250 B.n699 B.n396 585
R251 B.n400 B.n396 585
R252 B.n698 B.n697 585
R253 B.n697 B.n696 585
R254 B.n398 B.n397 585
R255 B.n399 B.n398 585
R256 B.n689 B.n688 585
R257 B.n690 B.n689 585
R258 B.n687 B.n405 585
R259 B.n405 B.n404 585
R260 B.n686 B.n685 585
R261 B.n685 B.n684 585
R262 B.n407 B.n406 585
R263 B.n408 B.n407 585
R264 B.n677 B.n676 585
R265 B.n678 B.n677 585
R266 B.n675 B.n413 585
R267 B.n413 B.n412 585
R268 B.n670 B.n669 585
R269 B.n668 B.n466 585
R270 B.n667 B.n465 585
R271 B.n672 B.n465 585
R272 B.n666 B.n665 585
R273 B.n664 B.n663 585
R274 B.n662 B.n661 585
R275 B.n660 B.n659 585
R276 B.n658 B.n657 585
R277 B.n656 B.n655 585
R278 B.n654 B.n653 585
R279 B.n652 B.n651 585
R280 B.n650 B.n649 585
R281 B.n648 B.n647 585
R282 B.n646 B.n645 585
R283 B.n644 B.n643 585
R284 B.n642 B.n641 585
R285 B.n640 B.n639 585
R286 B.n638 B.n637 585
R287 B.n636 B.n635 585
R288 B.n634 B.n633 585
R289 B.n632 B.n631 585
R290 B.n630 B.n629 585
R291 B.n628 B.n627 585
R292 B.n626 B.n625 585
R293 B.n624 B.n623 585
R294 B.n622 B.n621 585
R295 B.n620 B.n619 585
R296 B.n618 B.n617 585
R297 B.n616 B.n615 585
R298 B.n614 B.n613 585
R299 B.n612 B.n611 585
R300 B.n610 B.n609 585
R301 B.n608 B.n607 585
R302 B.n606 B.n605 585
R303 B.n604 B.n603 585
R304 B.n602 B.n601 585
R305 B.n600 B.n599 585
R306 B.n598 B.n597 585
R307 B.n596 B.n595 585
R308 B.n594 B.n593 585
R309 B.n592 B.n591 585
R310 B.n590 B.n589 585
R311 B.n588 B.n587 585
R312 B.n586 B.n585 585
R313 B.n584 B.n583 585
R314 B.n582 B.n581 585
R315 B.n579 B.n578 585
R316 B.n577 B.n576 585
R317 B.n575 B.n574 585
R318 B.n573 B.n572 585
R319 B.n571 B.n570 585
R320 B.n569 B.n568 585
R321 B.n567 B.n566 585
R322 B.n565 B.n564 585
R323 B.n563 B.n562 585
R324 B.n561 B.n560 585
R325 B.n558 B.n557 585
R326 B.n556 B.n555 585
R327 B.n554 B.n553 585
R328 B.n552 B.n551 585
R329 B.n550 B.n549 585
R330 B.n548 B.n547 585
R331 B.n546 B.n545 585
R332 B.n544 B.n543 585
R333 B.n542 B.n541 585
R334 B.n540 B.n539 585
R335 B.n538 B.n537 585
R336 B.n536 B.n535 585
R337 B.n534 B.n533 585
R338 B.n532 B.n531 585
R339 B.n530 B.n529 585
R340 B.n528 B.n527 585
R341 B.n526 B.n525 585
R342 B.n524 B.n523 585
R343 B.n522 B.n521 585
R344 B.n520 B.n519 585
R345 B.n518 B.n517 585
R346 B.n516 B.n515 585
R347 B.n514 B.n513 585
R348 B.n512 B.n511 585
R349 B.n510 B.n509 585
R350 B.n508 B.n507 585
R351 B.n506 B.n505 585
R352 B.n504 B.n503 585
R353 B.n502 B.n501 585
R354 B.n500 B.n499 585
R355 B.n498 B.n497 585
R356 B.n496 B.n495 585
R357 B.n494 B.n493 585
R358 B.n492 B.n491 585
R359 B.n490 B.n489 585
R360 B.n488 B.n487 585
R361 B.n486 B.n485 585
R362 B.n484 B.n483 585
R363 B.n482 B.n481 585
R364 B.n480 B.n479 585
R365 B.n478 B.n477 585
R366 B.n476 B.n475 585
R367 B.n474 B.n473 585
R368 B.n472 B.n471 585
R369 B.n415 B.n414 585
R370 B.n674 B.n673 585
R371 B.n673 B.n672 585
R372 B.n411 B.n410 585
R373 B.n412 B.n411 585
R374 B.n680 B.n679 585
R375 B.n679 B.n678 585
R376 B.n681 B.n409 585
R377 B.n409 B.n408 585
R378 B.n683 B.n682 585
R379 B.n684 B.n683 585
R380 B.n403 B.n402 585
R381 B.n404 B.n403 585
R382 B.n692 B.n691 585
R383 B.n691 B.n690 585
R384 B.n693 B.n401 585
R385 B.n401 B.n399 585
R386 B.n695 B.n694 585
R387 B.n696 B.n695 585
R388 B.n395 B.n394 585
R389 B.n400 B.n395 585
R390 B.n704 B.n703 585
R391 B.n703 B.n702 585
R392 B.n705 B.n393 585
R393 B.n393 B.n392 585
R394 B.n707 B.n706 585
R395 B.n708 B.n707 585
R396 B.n387 B.n386 585
R397 B.n388 B.n387 585
R398 B.n716 B.n715 585
R399 B.n715 B.n714 585
R400 B.n717 B.n385 585
R401 B.n385 B.n384 585
R402 B.n719 B.n718 585
R403 B.n720 B.n719 585
R404 B.n379 B.n378 585
R405 B.n380 B.n379 585
R406 B.n728 B.n727 585
R407 B.n727 B.n726 585
R408 B.n729 B.n377 585
R409 B.n377 B.n376 585
R410 B.n731 B.n730 585
R411 B.n732 B.n731 585
R412 B.n371 B.n370 585
R413 B.n372 B.n371 585
R414 B.n741 B.n740 585
R415 B.n740 B.n739 585
R416 B.n742 B.n369 585
R417 B.n738 B.n369 585
R418 B.n744 B.n743 585
R419 B.n745 B.n744 585
R420 B.n364 B.n363 585
R421 B.n365 B.n364 585
R422 B.n753 B.n752 585
R423 B.n752 B.n751 585
R424 B.n754 B.n362 585
R425 B.n362 B.n361 585
R426 B.n756 B.n755 585
R427 B.n757 B.n756 585
R428 B.n356 B.n355 585
R429 B.n357 B.n356 585
R430 B.n765 B.n764 585
R431 B.n764 B.n763 585
R432 B.n766 B.n354 585
R433 B.n354 B.n353 585
R434 B.n768 B.n767 585
R435 B.n769 B.n768 585
R436 B.n348 B.n347 585
R437 B.n349 B.n348 585
R438 B.n777 B.n776 585
R439 B.n776 B.n775 585
R440 B.n778 B.n346 585
R441 B.n346 B.n345 585
R442 B.n780 B.n779 585
R443 B.n781 B.n780 585
R444 B.n340 B.n339 585
R445 B.n341 B.n340 585
R446 B.n790 B.n789 585
R447 B.n789 B.n788 585
R448 B.n791 B.n338 585
R449 B.n338 B.n337 585
R450 B.n793 B.n792 585
R451 B.n794 B.n793 585
R452 B.n2 B.n0 585
R453 B.n4 B.n2 585
R454 B.n3 B.n1 585
R455 B.n934 B.n3 585
R456 B.n932 B.n931 585
R457 B.n933 B.n932 585
R458 B.n930 B.n9 585
R459 B.n9 B.n8 585
R460 B.n929 B.n928 585
R461 B.n928 B.n927 585
R462 B.n11 B.n10 585
R463 B.n926 B.n11 585
R464 B.n924 B.n923 585
R465 B.n925 B.n924 585
R466 B.n922 B.n16 585
R467 B.n16 B.n15 585
R468 B.n921 B.n920 585
R469 B.n920 B.n919 585
R470 B.n18 B.n17 585
R471 B.n918 B.n18 585
R472 B.n916 B.n915 585
R473 B.n917 B.n916 585
R474 B.n914 B.n23 585
R475 B.n23 B.n22 585
R476 B.n913 B.n912 585
R477 B.n912 B.n911 585
R478 B.n25 B.n24 585
R479 B.n910 B.n25 585
R480 B.n908 B.n907 585
R481 B.n909 B.n908 585
R482 B.n906 B.n30 585
R483 B.n30 B.n29 585
R484 B.n905 B.n904 585
R485 B.n904 B.n903 585
R486 B.n32 B.n31 585
R487 B.n902 B.n32 585
R488 B.n900 B.n899 585
R489 B.n901 B.n900 585
R490 B.n898 B.n36 585
R491 B.n39 B.n36 585
R492 B.n897 B.n896 585
R493 B.n896 B.n895 585
R494 B.n38 B.n37 585
R495 B.n894 B.n38 585
R496 B.n892 B.n891 585
R497 B.n893 B.n892 585
R498 B.n890 B.n44 585
R499 B.n44 B.n43 585
R500 B.n889 B.n888 585
R501 B.n888 B.n887 585
R502 B.n46 B.n45 585
R503 B.n886 B.n46 585
R504 B.n884 B.n883 585
R505 B.n885 B.n884 585
R506 B.n882 B.n51 585
R507 B.n51 B.n50 585
R508 B.n881 B.n880 585
R509 B.n880 B.n879 585
R510 B.n53 B.n52 585
R511 B.n878 B.n53 585
R512 B.n876 B.n875 585
R513 B.n877 B.n876 585
R514 B.n874 B.n58 585
R515 B.n58 B.n57 585
R516 B.n873 B.n872 585
R517 B.n872 B.n871 585
R518 B.n60 B.n59 585
R519 B.n870 B.n60 585
R520 B.n868 B.n867 585
R521 B.n869 B.n868 585
R522 B.n866 B.n65 585
R523 B.n65 B.n64 585
R524 B.n865 B.n864 585
R525 B.n864 B.n863 585
R526 B.n67 B.n66 585
R527 B.n862 B.n67 585
R528 B.n860 B.n859 585
R529 B.n861 B.n860 585
R530 B.n858 B.n72 585
R531 B.n72 B.n71 585
R532 B.n857 B.n856 585
R533 B.n856 B.n855 585
R534 B.n74 B.n73 585
R535 B.n854 B.n74 585
R536 B.n937 B.n936 585
R537 B.n936 B.n935 585
R538 B.n670 B.n411 478.086
R539 B.n134 B.n74 478.086
R540 B.n673 B.n413 478.086
R541 B.n851 B.n76 478.086
R542 B.n469 B.t7 380.293
R543 B.n467 B.t14 380.293
R544 B.n131 B.t10 380.293
R545 B.n128 B.t16 380.293
R546 B.n470 B.t6 307.76
R547 B.n129 B.t17 307.76
R548 B.n468 B.t13 307.76
R549 B.n132 B.t11 307.76
R550 B.n469 B.t4 304.281
R551 B.n467 B.t12 304.281
R552 B.n131 B.t8 304.281
R553 B.n128 B.t15 304.281
R554 B.n853 B.n852 256.663
R555 B.n853 B.n126 256.663
R556 B.n853 B.n125 256.663
R557 B.n853 B.n124 256.663
R558 B.n853 B.n123 256.663
R559 B.n853 B.n122 256.663
R560 B.n853 B.n121 256.663
R561 B.n853 B.n120 256.663
R562 B.n853 B.n119 256.663
R563 B.n853 B.n118 256.663
R564 B.n853 B.n117 256.663
R565 B.n853 B.n116 256.663
R566 B.n853 B.n115 256.663
R567 B.n853 B.n114 256.663
R568 B.n853 B.n113 256.663
R569 B.n853 B.n112 256.663
R570 B.n853 B.n111 256.663
R571 B.n853 B.n110 256.663
R572 B.n853 B.n109 256.663
R573 B.n853 B.n108 256.663
R574 B.n853 B.n107 256.663
R575 B.n853 B.n106 256.663
R576 B.n853 B.n105 256.663
R577 B.n853 B.n104 256.663
R578 B.n853 B.n103 256.663
R579 B.n853 B.n102 256.663
R580 B.n853 B.n101 256.663
R581 B.n853 B.n100 256.663
R582 B.n853 B.n99 256.663
R583 B.n853 B.n98 256.663
R584 B.n853 B.n97 256.663
R585 B.n853 B.n96 256.663
R586 B.n853 B.n95 256.663
R587 B.n853 B.n94 256.663
R588 B.n853 B.n93 256.663
R589 B.n853 B.n92 256.663
R590 B.n853 B.n91 256.663
R591 B.n853 B.n90 256.663
R592 B.n853 B.n89 256.663
R593 B.n853 B.n88 256.663
R594 B.n853 B.n87 256.663
R595 B.n853 B.n86 256.663
R596 B.n853 B.n85 256.663
R597 B.n853 B.n84 256.663
R598 B.n853 B.n83 256.663
R599 B.n853 B.n82 256.663
R600 B.n853 B.n81 256.663
R601 B.n853 B.n80 256.663
R602 B.n853 B.n79 256.663
R603 B.n853 B.n78 256.663
R604 B.n853 B.n77 256.663
R605 B.n672 B.n671 256.663
R606 B.n672 B.n416 256.663
R607 B.n672 B.n417 256.663
R608 B.n672 B.n418 256.663
R609 B.n672 B.n419 256.663
R610 B.n672 B.n420 256.663
R611 B.n672 B.n421 256.663
R612 B.n672 B.n422 256.663
R613 B.n672 B.n423 256.663
R614 B.n672 B.n424 256.663
R615 B.n672 B.n425 256.663
R616 B.n672 B.n426 256.663
R617 B.n672 B.n427 256.663
R618 B.n672 B.n428 256.663
R619 B.n672 B.n429 256.663
R620 B.n672 B.n430 256.663
R621 B.n672 B.n431 256.663
R622 B.n672 B.n432 256.663
R623 B.n672 B.n433 256.663
R624 B.n672 B.n434 256.663
R625 B.n672 B.n435 256.663
R626 B.n672 B.n436 256.663
R627 B.n672 B.n437 256.663
R628 B.n672 B.n438 256.663
R629 B.n672 B.n439 256.663
R630 B.n672 B.n440 256.663
R631 B.n672 B.n441 256.663
R632 B.n672 B.n442 256.663
R633 B.n672 B.n443 256.663
R634 B.n672 B.n444 256.663
R635 B.n672 B.n445 256.663
R636 B.n672 B.n446 256.663
R637 B.n672 B.n447 256.663
R638 B.n672 B.n448 256.663
R639 B.n672 B.n449 256.663
R640 B.n672 B.n450 256.663
R641 B.n672 B.n451 256.663
R642 B.n672 B.n452 256.663
R643 B.n672 B.n453 256.663
R644 B.n672 B.n454 256.663
R645 B.n672 B.n455 256.663
R646 B.n672 B.n456 256.663
R647 B.n672 B.n457 256.663
R648 B.n672 B.n458 256.663
R649 B.n672 B.n459 256.663
R650 B.n672 B.n460 256.663
R651 B.n672 B.n461 256.663
R652 B.n672 B.n462 256.663
R653 B.n672 B.n463 256.663
R654 B.n672 B.n464 256.663
R655 B.n679 B.n411 163.367
R656 B.n679 B.n409 163.367
R657 B.n683 B.n409 163.367
R658 B.n683 B.n403 163.367
R659 B.n691 B.n403 163.367
R660 B.n691 B.n401 163.367
R661 B.n695 B.n401 163.367
R662 B.n695 B.n395 163.367
R663 B.n703 B.n395 163.367
R664 B.n703 B.n393 163.367
R665 B.n707 B.n393 163.367
R666 B.n707 B.n387 163.367
R667 B.n715 B.n387 163.367
R668 B.n715 B.n385 163.367
R669 B.n719 B.n385 163.367
R670 B.n719 B.n379 163.367
R671 B.n727 B.n379 163.367
R672 B.n727 B.n377 163.367
R673 B.n731 B.n377 163.367
R674 B.n731 B.n371 163.367
R675 B.n740 B.n371 163.367
R676 B.n740 B.n369 163.367
R677 B.n744 B.n369 163.367
R678 B.n744 B.n364 163.367
R679 B.n752 B.n364 163.367
R680 B.n752 B.n362 163.367
R681 B.n756 B.n362 163.367
R682 B.n756 B.n356 163.367
R683 B.n764 B.n356 163.367
R684 B.n764 B.n354 163.367
R685 B.n768 B.n354 163.367
R686 B.n768 B.n348 163.367
R687 B.n776 B.n348 163.367
R688 B.n776 B.n346 163.367
R689 B.n780 B.n346 163.367
R690 B.n780 B.n340 163.367
R691 B.n789 B.n340 163.367
R692 B.n789 B.n338 163.367
R693 B.n793 B.n338 163.367
R694 B.n793 B.n2 163.367
R695 B.n936 B.n2 163.367
R696 B.n936 B.n3 163.367
R697 B.n932 B.n3 163.367
R698 B.n932 B.n9 163.367
R699 B.n928 B.n9 163.367
R700 B.n928 B.n11 163.367
R701 B.n924 B.n11 163.367
R702 B.n924 B.n16 163.367
R703 B.n920 B.n16 163.367
R704 B.n920 B.n18 163.367
R705 B.n916 B.n18 163.367
R706 B.n916 B.n23 163.367
R707 B.n912 B.n23 163.367
R708 B.n912 B.n25 163.367
R709 B.n908 B.n25 163.367
R710 B.n908 B.n30 163.367
R711 B.n904 B.n30 163.367
R712 B.n904 B.n32 163.367
R713 B.n900 B.n32 163.367
R714 B.n900 B.n36 163.367
R715 B.n896 B.n36 163.367
R716 B.n896 B.n38 163.367
R717 B.n892 B.n38 163.367
R718 B.n892 B.n44 163.367
R719 B.n888 B.n44 163.367
R720 B.n888 B.n46 163.367
R721 B.n884 B.n46 163.367
R722 B.n884 B.n51 163.367
R723 B.n880 B.n51 163.367
R724 B.n880 B.n53 163.367
R725 B.n876 B.n53 163.367
R726 B.n876 B.n58 163.367
R727 B.n872 B.n58 163.367
R728 B.n872 B.n60 163.367
R729 B.n868 B.n60 163.367
R730 B.n868 B.n65 163.367
R731 B.n864 B.n65 163.367
R732 B.n864 B.n67 163.367
R733 B.n860 B.n67 163.367
R734 B.n860 B.n72 163.367
R735 B.n856 B.n72 163.367
R736 B.n856 B.n74 163.367
R737 B.n466 B.n465 163.367
R738 B.n665 B.n465 163.367
R739 B.n663 B.n662 163.367
R740 B.n659 B.n658 163.367
R741 B.n655 B.n654 163.367
R742 B.n651 B.n650 163.367
R743 B.n647 B.n646 163.367
R744 B.n643 B.n642 163.367
R745 B.n639 B.n638 163.367
R746 B.n635 B.n634 163.367
R747 B.n631 B.n630 163.367
R748 B.n627 B.n626 163.367
R749 B.n623 B.n622 163.367
R750 B.n619 B.n618 163.367
R751 B.n615 B.n614 163.367
R752 B.n611 B.n610 163.367
R753 B.n607 B.n606 163.367
R754 B.n603 B.n602 163.367
R755 B.n599 B.n598 163.367
R756 B.n595 B.n594 163.367
R757 B.n591 B.n590 163.367
R758 B.n587 B.n586 163.367
R759 B.n583 B.n582 163.367
R760 B.n578 B.n577 163.367
R761 B.n574 B.n573 163.367
R762 B.n570 B.n569 163.367
R763 B.n566 B.n565 163.367
R764 B.n562 B.n561 163.367
R765 B.n557 B.n556 163.367
R766 B.n553 B.n552 163.367
R767 B.n549 B.n548 163.367
R768 B.n545 B.n544 163.367
R769 B.n541 B.n540 163.367
R770 B.n537 B.n536 163.367
R771 B.n533 B.n532 163.367
R772 B.n529 B.n528 163.367
R773 B.n525 B.n524 163.367
R774 B.n521 B.n520 163.367
R775 B.n517 B.n516 163.367
R776 B.n513 B.n512 163.367
R777 B.n509 B.n508 163.367
R778 B.n505 B.n504 163.367
R779 B.n501 B.n500 163.367
R780 B.n497 B.n496 163.367
R781 B.n493 B.n492 163.367
R782 B.n489 B.n488 163.367
R783 B.n485 B.n484 163.367
R784 B.n481 B.n480 163.367
R785 B.n477 B.n476 163.367
R786 B.n473 B.n472 163.367
R787 B.n673 B.n415 163.367
R788 B.n677 B.n413 163.367
R789 B.n677 B.n407 163.367
R790 B.n685 B.n407 163.367
R791 B.n685 B.n405 163.367
R792 B.n689 B.n405 163.367
R793 B.n689 B.n398 163.367
R794 B.n697 B.n398 163.367
R795 B.n697 B.n396 163.367
R796 B.n701 B.n396 163.367
R797 B.n701 B.n391 163.367
R798 B.n709 B.n391 163.367
R799 B.n709 B.n389 163.367
R800 B.n713 B.n389 163.367
R801 B.n713 B.n383 163.367
R802 B.n721 B.n383 163.367
R803 B.n721 B.n381 163.367
R804 B.n725 B.n381 163.367
R805 B.n725 B.n375 163.367
R806 B.n733 B.n375 163.367
R807 B.n733 B.n373 163.367
R808 B.n737 B.n373 163.367
R809 B.n737 B.n368 163.367
R810 B.n746 B.n368 163.367
R811 B.n746 B.n366 163.367
R812 B.n750 B.n366 163.367
R813 B.n750 B.n360 163.367
R814 B.n758 B.n360 163.367
R815 B.n758 B.n358 163.367
R816 B.n762 B.n358 163.367
R817 B.n762 B.n352 163.367
R818 B.n770 B.n352 163.367
R819 B.n770 B.n350 163.367
R820 B.n774 B.n350 163.367
R821 B.n774 B.n344 163.367
R822 B.n782 B.n344 163.367
R823 B.n782 B.n342 163.367
R824 B.n787 B.n342 163.367
R825 B.n787 B.n336 163.367
R826 B.n795 B.n336 163.367
R827 B.n796 B.n795 163.367
R828 B.n796 B.n5 163.367
R829 B.n6 B.n5 163.367
R830 B.n7 B.n6 163.367
R831 B.n801 B.n7 163.367
R832 B.n801 B.n12 163.367
R833 B.n13 B.n12 163.367
R834 B.n14 B.n13 163.367
R835 B.n806 B.n14 163.367
R836 B.n806 B.n19 163.367
R837 B.n20 B.n19 163.367
R838 B.n21 B.n20 163.367
R839 B.n811 B.n21 163.367
R840 B.n811 B.n26 163.367
R841 B.n27 B.n26 163.367
R842 B.n28 B.n27 163.367
R843 B.n816 B.n28 163.367
R844 B.n816 B.n33 163.367
R845 B.n34 B.n33 163.367
R846 B.n35 B.n34 163.367
R847 B.n821 B.n35 163.367
R848 B.n821 B.n40 163.367
R849 B.n41 B.n40 163.367
R850 B.n42 B.n41 163.367
R851 B.n826 B.n42 163.367
R852 B.n826 B.n47 163.367
R853 B.n48 B.n47 163.367
R854 B.n49 B.n48 163.367
R855 B.n831 B.n49 163.367
R856 B.n831 B.n54 163.367
R857 B.n55 B.n54 163.367
R858 B.n56 B.n55 163.367
R859 B.n836 B.n56 163.367
R860 B.n836 B.n61 163.367
R861 B.n62 B.n61 163.367
R862 B.n63 B.n62 163.367
R863 B.n841 B.n63 163.367
R864 B.n841 B.n68 163.367
R865 B.n69 B.n68 163.367
R866 B.n70 B.n69 163.367
R867 B.n846 B.n70 163.367
R868 B.n846 B.n75 163.367
R869 B.n76 B.n75 163.367
R870 B.n138 B.n137 163.367
R871 B.n142 B.n141 163.367
R872 B.n146 B.n145 163.367
R873 B.n150 B.n149 163.367
R874 B.n154 B.n153 163.367
R875 B.n158 B.n157 163.367
R876 B.n162 B.n161 163.367
R877 B.n166 B.n165 163.367
R878 B.n170 B.n169 163.367
R879 B.n174 B.n173 163.367
R880 B.n178 B.n177 163.367
R881 B.n182 B.n181 163.367
R882 B.n186 B.n185 163.367
R883 B.n190 B.n189 163.367
R884 B.n194 B.n193 163.367
R885 B.n198 B.n197 163.367
R886 B.n202 B.n201 163.367
R887 B.n206 B.n205 163.367
R888 B.n210 B.n209 163.367
R889 B.n214 B.n213 163.367
R890 B.n218 B.n217 163.367
R891 B.n222 B.n221 163.367
R892 B.n226 B.n225 163.367
R893 B.n230 B.n229 163.367
R894 B.n234 B.n233 163.367
R895 B.n238 B.n237 163.367
R896 B.n242 B.n241 163.367
R897 B.n246 B.n245 163.367
R898 B.n250 B.n249 163.367
R899 B.n254 B.n253 163.367
R900 B.n258 B.n257 163.367
R901 B.n262 B.n261 163.367
R902 B.n266 B.n265 163.367
R903 B.n270 B.n269 163.367
R904 B.n274 B.n273 163.367
R905 B.n278 B.n277 163.367
R906 B.n282 B.n281 163.367
R907 B.n286 B.n285 163.367
R908 B.n290 B.n289 163.367
R909 B.n294 B.n293 163.367
R910 B.n298 B.n297 163.367
R911 B.n302 B.n301 163.367
R912 B.n306 B.n305 163.367
R913 B.n310 B.n309 163.367
R914 B.n314 B.n313 163.367
R915 B.n318 B.n317 163.367
R916 B.n322 B.n321 163.367
R917 B.n326 B.n325 163.367
R918 B.n330 B.n329 163.367
R919 B.n332 B.n127 163.367
R920 B.n672 B.n412 76.8333
R921 B.n854 B.n853 76.8333
R922 B.n470 B.n469 72.5338
R923 B.n468 B.n467 72.5338
R924 B.n132 B.n131 72.5338
R925 B.n129 B.n128 72.5338
R926 B.n671 B.n670 71.676
R927 B.n665 B.n416 71.676
R928 B.n662 B.n417 71.676
R929 B.n658 B.n418 71.676
R930 B.n654 B.n419 71.676
R931 B.n650 B.n420 71.676
R932 B.n646 B.n421 71.676
R933 B.n642 B.n422 71.676
R934 B.n638 B.n423 71.676
R935 B.n634 B.n424 71.676
R936 B.n630 B.n425 71.676
R937 B.n626 B.n426 71.676
R938 B.n622 B.n427 71.676
R939 B.n618 B.n428 71.676
R940 B.n614 B.n429 71.676
R941 B.n610 B.n430 71.676
R942 B.n606 B.n431 71.676
R943 B.n602 B.n432 71.676
R944 B.n598 B.n433 71.676
R945 B.n594 B.n434 71.676
R946 B.n590 B.n435 71.676
R947 B.n586 B.n436 71.676
R948 B.n582 B.n437 71.676
R949 B.n577 B.n438 71.676
R950 B.n573 B.n439 71.676
R951 B.n569 B.n440 71.676
R952 B.n565 B.n441 71.676
R953 B.n561 B.n442 71.676
R954 B.n556 B.n443 71.676
R955 B.n552 B.n444 71.676
R956 B.n548 B.n445 71.676
R957 B.n544 B.n446 71.676
R958 B.n540 B.n447 71.676
R959 B.n536 B.n448 71.676
R960 B.n532 B.n449 71.676
R961 B.n528 B.n450 71.676
R962 B.n524 B.n451 71.676
R963 B.n520 B.n452 71.676
R964 B.n516 B.n453 71.676
R965 B.n512 B.n454 71.676
R966 B.n508 B.n455 71.676
R967 B.n504 B.n456 71.676
R968 B.n500 B.n457 71.676
R969 B.n496 B.n458 71.676
R970 B.n492 B.n459 71.676
R971 B.n488 B.n460 71.676
R972 B.n484 B.n461 71.676
R973 B.n480 B.n462 71.676
R974 B.n476 B.n463 71.676
R975 B.n472 B.n464 71.676
R976 B.n134 B.n77 71.676
R977 B.n138 B.n78 71.676
R978 B.n142 B.n79 71.676
R979 B.n146 B.n80 71.676
R980 B.n150 B.n81 71.676
R981 B.n154 B.n82 71.676
R982 B.n158 B.n83 71.676
R983 B.n162 B.n84 71.676
R984 B.n166 B.n85 71.676
R985 B.n170 B.n86 71.676
R986 B.n174 B.n87 71.676
R987 B.n178 B.n88 71.676
R988 B.n182 B.n89 71.676
R989 B.n186 B.n90 71.676
R990 B.n190 B.n91 71.676
R991 B.n194 B.n92 71.676
R992 B.n198 B.n93 71.676
R993 B.n202 B.n94 71.676
R994 B.n206 B.n95 71.676
R995 B.n210 B.n96 71.676
R996 B.n214 B.n97 71.676
R997 B.n218 B.n98 71.676
R998 B.n222 B.n99 71.676
R999 B.n226 B.n100 71.676
R1000 B.n230 B.n101 71.676
R1001 B.n234 B.n102 71.676
R1002 B.n238 B.n103 71.676
R1003 B.n242 B.n104 71.676
R1004 B.n246 B.n105 71.676
R1005 B.n250 B.n106 71.676
R1006 B.n254 B.n107 71.676
R1007 B.n258 B.n108 71.676
R1008 B.n262 B.n109 71.676
R1009 B.n266 B.n110 71.676
R1010 B.n270 B.n111 71.676
R1011 B.n274 B.n112 71.676
R1012 B.n278 B.n113 71.676
R1013 B.n282 B.n114 71.676
R1014 B.n286 B.n115 71.676
R1015 B.n290 B.n116 71.676
R1016 B.n294 B.n117 71.676
R1017 B.n298 B.n118 71.676
R1018 B.n302 B.n119 71.676
R1019 B.n306 B.n120 71.676
R1020 B.n310 B.n121 71.676
R1021 B.n314 B.n122 71.676
R1022 B.n318 B.n123 71.676
R1023 B.n322 B.n124 71.676
R1024 B.n326 B.n125 71.676
R1025 B.n330 B.n126 71.676
R1026 B.n852 B.n127 71.676
R1027 B.n852 B.n851 71.676
R1028 B.n332 B.n126 71.676
R1029 B.n329 B.n125 71.676
R1030 B.n325 B.n124 71.676
R1031 B.n321 B.n123 71.676
R1032 B.n317 B.n122 71.676
R1033 B.n313 B.n121 71.676
R1034 B.n309 B.n120 71.676
R1035 B.n305 B.n119 71.676
R1036 B.n301 B.n118 71.676
R1037 B.n297 B.n117 71.676
R1038 B.n293 B.n116 71.676
R1039 B.n289 B.n115 71.676
R1040 B.n285 B.n114 71.676
R1041 B.n281 B.n113 71.676
R1042 B.n277 B.n112 71.676
R1043 B.n273 B.n111 71.676
R1044 B.n269 B.n110 71.676
R1045 B.n265 B.n109 71.676
R1046 B.n261 B.n108 71.676
R1047 B.n257 B.n107 71.676
R1048 B.n253 B.n106 71.676
R1049 B.n249 B.n105 71.676
R1050 B.n245 B.n104 71.676
R1051 B.n241 B.n103 71.676
R1052 B.n237 B.n102 71.676
R1053 B.n233 B.n101 71.676
R1054 B.n229 B.n100 71.676
R1055 B.n225 B.n99 71.676
R1056 B.n221 B.n98 71.676
R1057 B.n217 B.n97 71.676
R1058 B.n213 B.n96 71.676
R1059 B.n209 B.n95 71.676
R1060 B.n205 B.n94 71.676
R1061 B.n201 B.n93 71.676
R1062 B.n197 B.n92 71.676
R1063 B.n193 B.n91 71.676
R1064 B.n189 B.n90 71.676
R1065 B.n185 B.n89 71.676
R1066 B.n181 B.n88 71.676
R1067 B.n177 B.n87 71.676
R1068 B.n173 B.n86 71.676
R1069 B.n169 B.n85 71.676
R1070 B.n165 B.n84 71.676
R1071 B.n161 B.n83 71.676
R1072 B.n157 B.n82 71.676
R1073 B.n153 B.n81 71.676
R1074 B.n149 B.n80 71.676
R1075 B.n145 B.n79 71.676
R1076 B.n141 B.n78 71.676
R1077 B.n137 B.n77 71.676
R1078 B.n671 B.n466 71.676
R1079 B.n663 B.n416 71.676
R1080 B.n659 B.n417 71.676
R1081 B.n655 B.n418 71.676
R1082 B.n651 B.n419 71.676
R1083 B.n647 B.n420 71.676
R1084 B.n643 B.n421 71.676
R1085 B.n639 B.n422 71.676
R1086 B.n635 B.n423 71.676
R1087 B.n631 B.n424 71.676
R1088 B.n627 B.n425 71.676
R1089 B.n623 B.n426 71.676
R1090 B.n619 B.n427 71.676
R1091 B.n615 B.n428 71.676
R1092 B.n611 B.n429 71.676
R1093 B.n607 B.n430 71.676
R1094 B.n603 B.n431 71.676
R1095 B.n599 B.n432 71.676
R1096 B.n595 B.n433 71.676
R1097 B.n591 B.n434 71.676
R1098 B.n587 B.n435 71.676
R1099 B.n583 B.n436 71.676
R1100 B.n578 B.n437 71.676
R1101 B.n574 B.n438 71.676
R1102 B.n570 B.n439 71.676
R1103 B.n566 B.n440 71.676
R1104 B.n562 B.n441 71.676
R1105 B.n557 B.n442 71.676
R1106 B.n553 B.n443 71.676
R1107 B.n549 B.n444 71.676
R1108 B.n545 B.n445 71.676
R1109 B.n541 B.n446 71.676
R1110 B.n537 B.n447 71.676
R1111 B.n533 B.n448 71.676
R1112 B.n529 B.n449 71.676
R1113 B.n525 B.n450 71.676
R1114 B.n521 B.n451 71.676
R1115 B.n517 B.n452 71.676
R1116 B.n513 B.n453 71.676
R1117 B.n509 B.n454 71.676
R1118 B.n505 B.n455 71.676
R1119 B.n501 B.n456 71.676
R1120 B.n497 B.n457 71.676
R1121 B.n493 B.n458 71.676
R1122 B.n489 B.n459 71.676
R1123 B.n485 B.n460 71.676
R1124 B.n481 B.n461 71.676
R1125 B.n477 B.n462 71.676
R1126 B.n473 B.n463 71.676
R1127 B.n464 B.n415 71.676
R1128 B.n559 B.n470 59.5399
R1129 B.n580 B.n468 59.5399
R1130 B.n133 B.n132 59.5399
R1131 B.n130 B.n129 59.5399
R1132 B.n678 B.n412 39.8832
R1133 B.n678 B.n408 39.8832
R1134 B.n684 B.n408 39.8832
R1135 B.n684 B.n404 39.8832
R1136 B.n690 B.n404 39.8832
R1137 B.n690 B.n399 39.8832
R1138 B.n696 B.n399 39.8832
R1139 B.n696 B.n400 39.8832
R1140 B.n702 B.n392 39.8832
R1141 B.n708 B.n392 39.8832
R1142 B.n708 B.n388 39.8832
R1143 B.n714 B.n388 39.8832
R1144 B.n714 B.n384 39.8832
R1145 B.n720 B.n384 39.8832
R1146 B.n720 B.n380 39.8832
R1147 B.n726 B.n380 39.8832
R1148 B.n726 B.n376 39.8832
R1149 B.n732 B.n376 39.8832
R1150 B.n732 B.n372 39.8832
R1151 B.n739 B.n372 39.8832
R1152 B.n739 B.n738 39.8832
R1153 B.n745 B.n365 39.8832
R1154 B.n751 B.n365 39.8832
R1155 B.n751 B.n361 39.8832
R1156 B.n757 B.n361 39.8832
R1157 B.n757 B.n357 39.8832
R1158 B.n763 B.n357 39.8832
R1159 B.n763 B.n353 39.8832
R1160 B.n769 B.n353 39.8832
R1161 B.n769 B.n349 39.8832
R1162 B.n775 B.n349 39.8832
R1163 B.n781 B.n345 39.8832
R1164 B.n781 B.n341 39.8832
R1165 B.n788 B.n341 39.8832
R1166 B.n788 B.n337 39.8832
R1167 B.n794 B.n337 39.8832
R1168 B.n794 B.n4 39.8832
R1169 B.n935 B.n4 39.8832
R1170 B.n935 B.n934 39.8832
R1171 B.n934 B.n933 39.8832
R1172 B.n933 B.n8 39.8832
R1173 B.n927 B.n8 39.8832
R1174 B.n927 B.n926 39.8832
R1175 B.n926 B.n925 39.8832
R1176 B.n925 B.n15 39.8832
R1177 B.n919 B.n918 39.8832
R1178 B.n918 B.n917 39.8832
R1179 B.n917 B.n22 39.8832
R1180 B.n911 B.n22 39.8832
R1181 B.n911 B.n910 39.8832
R1182 B.n910 B.n909 39.8832
R1183 B.n909 B.n29 39.8832
R1184 B.n903 B.n29 39.8832
R1185 B.n903 B.n902 39.8832
R1186 B.n902 B.n901 39.8832
R1187 B.n895 B.n39 39.8832
R1188 B.n895 B.n894 39.8832
R1189 B.n894 B.n893 39.8832
R1190 B.n893 B.n43 39.8832
R1191 B.n887 B.n43 39.8832
R1192 B.n887 B.n886 39.8832
R1193 B.n886 B.n885 39.8832
R1194 B.n885 B.n50 39.8832
R1195 B.n879 B.n50 39.8832
R1196 B.n879 B.n878 39.8832
R1197 B.n878 B.n877 39.8832
R1198 B.n877 B.n57 39.8832
R1199 B.n871 B.n57 39.8832
R1200 B.n870 B.n869 39.8832
R1201 B.n869 B.n64 39.8832
R1202 B.n863 B.n64 39.8832
R1203 B.n863 B.n862 39.8832
R1204 B.n862 B.n861 39.8832
R1205 B.n861 B.n71 39.8832
R1206 B.n855 B.n71 39.8832
R1207 B.n855 B.n854 39.8832
R1208 B.n738 B.t0 35.7776
R1209 B.n775 B.t2 35.7776
R1210 B.n919 B.t3 35.7776
R1211 B.n39 B.t1 35.7776
R1212 B.n135 B.n73 31.0639
R1213 B.n850 B.n849 31.0639
R1214 B.n675 B.n674 31.0639
R1215 B.n669 B.n410 31.0639
R1216 B.n400 B.t5 27.5665
R1217 B.t9 B.n870 27.5665
R1218 B B.n937 18.0485
R1219 B.n702 B.t5 12.3172
R1220 B.n871 B.t9 12.3172
R1221 B.n136 B.n135 10.6151
R1222 B.n139 B.n136 10.6151
R1223 B.n140 B.n139 10.6151
R1224 B.n143 B.n140 10.6151
R1225 B.n144 B.n143 10.6151
R1226 B.n147 B.n144 10.6151
R1227 B.n148 B.n147 10.6151
R1228 B.n151 B.n148 10.6151
R1229 B.n152 B.n151 10.6151
R1230 B.n155 B.n152 10.6151
R1231 B.n156 B.n155 10.6151
R1232 B.n159 B.n156 10.6151
R1233 B.n160 B.n159 10.6151
R1234 B.n163 B.n160 10.6151
R1235 B.n164 B.n163 10.6151
R1236 B.n167 B.n164 10.6151
R1237 B.n168 B.n167 10.6151
R1238 B.n171 B.n168 10.6151
R1239 B.n172 B.n171 10.6151
R1240 B.n175 B.n172 10.6151
R1241 B.n176 B.n175 10.6151
R1242 B.n179 B.n176 10.6151
R1243 B.n180 B.n179 10.6151
R1244 B.n183 B.n180 10.6151
R1245 B.n184 B.n183 10.6151
R1246 B.n187 B.n184 10.6151
R1247 B.n188 B.n187 10.6151
R1248 B.n191 B.n188 10.6151
R1249 B.n192 B.n191 10.6151
R1250 B.n195 B.n192 10.6151
R1251 B.n196 B.n195 10.6151
R1252 B.n199 B.n196 10.6151
R1253 B.n200 B.n199 10.6151
R1254 B.n203 B.n200 10.6151
R1255 B.n204 B.n203 10.6151
R1256 B.n207 B.n204 10.6151
R1257 B.n208 B.n207 10.6151
R1258 B.n211 B.n208 10.6151
R1259 B.n212 B.n211 10.6151
R1260 B.n215 B.n212 10.6151
R1261 B.n216 B.n215 10.6151
R1262 B.n219 B.n216 10.6151
R1263 B.n220 B.n219 10.6151
R1264 B.n223 B.n220 10.6151
R1265 B.n224 B.n223 10.6151
R1266 B.n228 B.n227 10.6151
R1267 B.n231 B.n228 10.6151
R1268 B.n232 B.n231 10.6151
R1269 B.n235 B.n232 10.6151
R1270 B.n236 B.n235 10.6151
R1271 B.n239 B.n236 10.6151
R1272 B.n240 B.n239 10.6151
R1273 B.n243 B.n240 10.6151
R1274 B.n244 B.n243 10.6151
R1275 B.n248 B.n247 10.6151
R1276 B.n251 B.n248 10.6151
R1277 B.n252 B.n251 10.6151
R1278 B.n255 B.n252 10.6151
R1279 B.n256 B.n255 10.6151
R1280 B.n259 B.n256 10.6151
R1281 B.n260 B.n259 10.6151
R1282 B.n263 B.n260 10.6151
R1283 B.n264 B.n263 10.6151
R1284 B.n267 B.n264 10.6151
R1285 B.n268 B.n267 10.6151
R1286 B.n271 B.n268 10.6151
R1287 B.n272 B.n271 10.6151
R1288 B.n275 B.n272 10.6151
R1289 B.n276 B.n275 10.6151
R1290 B.n279 B.n276 10.6151
R1291 B.n280 B.n279 10.6151
R1292 B.n283 B.n280 10.6151
R1293 B.n284 B.n283 10.6151
R1294 B.n287 B.n284 10.6151
R1295 B.n288 B.n287 10.6151
R1296 B.n291 B.n288 10.6151
R1297 B.n292 B.n291 10.6151
R1298 B.n295 B.n292 10.6151
R1299 B.n296 B.n295 10.6151
R1300 B.n299 B.n296 10.6151
R1301 B.n300 B.n299 10.6151
R1302 B.n303 B.n300 10.6151
R1303 B.n304 B.n303 10.6151
R1304 B.n307 B.n304 10.6151
R1305 B.n308 B.n307 10.6151
R1306 B.n311 B.n308 10.6151
R1307 B.n312 B.n311 10.6151
R1308 B.n315 B.n312 10.6151
R1309 B.n316 B.n315 10.6151
R1310 B.n319 B.n316 10.6151
R1311 B.n320 B.n319 10.6151
R1312 B.n323 B.n320 10.6151
R1313 B.n324 B.n323 10.6151
R1314 B.n327 B.n324 10.6151
R1315 B.n328 B.n327 10.6151
R1316 B.n331 B.n328 10.6151
R1317 B.n333 B.n331 10.6151
R1318 B.n334 B.n333 10.6151
R1319 B.n850 B.n334 10.6151
R1320 B.n676 B.n675 10.6151
R1321 B.n676 B.n406 10.6151
R1322 B.n686 B.n406 10.6151
R1323 B.n687 B.n686 10.6151
R1324 B.n688 B.n687 10.6151
R1325 B.n688 B.n397 10.6151
R1326 B.n698 B.n397 10.6151
R1327 B.n699 B.n698 10.6151
R1328 B.n700 B.n699 10.6151
R1329 B.n700 B.n390 10.6151
R1330 B.n710 B.n390 10.6151
R1331 B.n711 B.n710 10.6151
R1332 B.n712 B.n711 10.6151
R1333 B.n712 B.n382 10.6151
R1334 B.n722 B.n382 10.6151
R1335 B.n723 B.n722 10.6151
R1336 B.n724 B.n723 10.6151
R1337 B.n724 B.n374 10.6151
R1338 B.n734 B.n374 10.6151
R1339 B.n735 B.n734 10.6151
R1340 B.n736 B.n735 10.6151
R1341 B.n736 B.n367 10.6151
R1342 B.n747 B.n367 10.6151
R1343 B.n748 B.n747 10.6151
R1344 B.n749 B.n748 10.6151
R1345 B.n749 B.n359 10.6151
R1346 B.n759 B.n359 10.6151
R1347 B.n760 B.n759 10.6151
R1348 B.n761 B.n760 10.6151
R1349 B.n761 B.n351 10.6151
R1350 B.n771 B.n351 10.6151
R1351 B.n772 B.n771 10.6151
R1352 B.n773 B.n772 10.6151
R1353 B.n773 B.n343 10.6151
R1354 B.n783 B.n343 10.6151
R1355 B.n784 B.n783 10.6151
R1356 B.n786 B.n784 10.6151
R1357 B.n786 B.n785 10.6151
R1358 B.n785 B.n335 10.6151
R1359 B.n797 B.n335 10.6151
R1360 B.n798 B.n797 10.6151
R1361 B.n799 B.n798 10.6151
R1362 B.n800 B.n799 10.6151
R1363 B.n802 B.n800 10.6151
R1364 B.n803 B.n802 10.6151
R1365 B.n804 B.n803 10.6151
R1366 B.n805 B.n804 10.6151
R1367 B.n807 B.n805 10.6151
R1368 B.n808 B.n807 10.6151
R1369 B.n809 B.n808 10.6151
R1370 B.n810 B.n809 10.6151
R1371 B.n812 B.n810 10.6151
R1372 B.n813 B.n812 10.6151
R1373 B.n814 B.n813 10.6151
R1374 B.n815 B.n814 10.6151
R1375 B.n817 B.n815 10.6151
R1376 B.n818 B.n817 10.6151
R1377 B.n819 B.n818 10.6151
R1378 B.n820 B.n819 10.6151
R1379 B.n822 B.n820 10.6151
R1380 B.n823 B.n822 10.6151
R1381 B.n824 B.n823 10.6151
R1382 B.n825 B.n824 10.6151
R1383 B.n827 B.n825 10.6151
R1384 B.n828 B.n827 10.6151
R1385 B.n829 B.n828 10.6151
R1386 B.n830 B.n829 10.6151
R1387 B.n832 B.n830 10.6151
R1388 B.n833 B.n832 10.6151
R1389 B.n834 B.n833 10.6151
R1390 B.n835 B.n834 10.6151
R1391 B.n837 B.n835 10.6151
R1392 B.n838 B.n837 10.6151
R1393 B.n839 B.n838 10.6151
R1394 B.n840 B.n839 10.6151
R1395 B.n842 B.n840 10.6151
R1396 B.n843 B.n842 10.6151
R1397 B.n844 B.n843 10.6151
R1398 B.n845 B.n844 10.6151
R1399 B.n847 B.n845 10.6151
R1400 B.n848 B.n847 10.6151
R1401 B.n849 B.n848 10.6151
R1402 B.n669 B.n668 10.6151
R1403 B.n668 B.n667 10.6151
R1404 B.n667 B.n666 10.6151
R1405 B.n666 B.n664 10.6151
R1406 B.n664 B.n661 10.6151
R1407 B.n661 B.n660 10.6151
R1408 B.n660 B.n657 10.6151
R1409 B.n657 B.n656 10.6151
R1410 B.n656 B.n653 10.6151
R1411 B.n653 B.n652 10.6151
R1412 B.n652 B.n649 10.6151
R1413 B.n649 B.n648 10.6151
R1414 B.n648 B.n645 10.6151
R1415 B.n645 B.n644 10.6151
R1416 B.n644 B.n641 10.6151
R1417 B.n641 B.n640 10.6151
R1418 B.n640 B.n637 10.6151
R1419 B.n637 B.n636 10.6151
R1420 B.n636 B.n633 10.6151
R1421 B.n633 B.n632 10.6151
R1422 B.n632 B.n629 10.6151
R1423 B.n629 B.n628 10.6151
R1424 B.n628 B.n625 10.6151
R1425 B.n625 B.n624 10.6151
R1426 B.n624 B.n621 10.6151
R1427 B.n621 B.n620 10.6151
R1428 B.n620 B.n617 10.6151
R1429 B.n617 B.n616 10.6151
R1430 B.n616 B.n613 10.6151
R1431 B.n613 B.n612 10.6151
R1432 B.n612 B.n609 10.6151
R1433 B.n609 B.n608 10.6151
R1434 B.n608 B.n605 10.6151
R1435 B.n605 B.n604 10.6151
R1436 B.n604 B.n601 10.6151
R1437 B.n601 B.n600 10.6151
R1438 B.n600 B.n597 10.6151
R1439 B.n597 B.n596 10.6151
R1440 B.n596 B.n593 10.6151
R1441 B.n593 B.n592 10.6151
R1442 B.n592 B.n589 10.6151
R1443 B.n589 B.n588 10.6151
R1444 B.n588 B.n585 10.6151
R1445 B.n585 B.n584 10.6151
R1446 B.n584 B.n581 10.6151
R1447 B.n579 B.n576 10.6151
R1448 B.n576 B.n575 10.6151
R1449 B.n575 B.n572 10.6151
R1450 B.n572 B.n571 10.6151
R1451 B.n571 B.n568 10.6151
R1452 B.n568 B.n567 10.6151
R1453 B.n567 B.n564 10.6151
R1454 B.n564 B.n563 10.6151
R1455 B.n563 B.n560 10.6151
R1456 B.n558 B.n555 10.6151
R1457 B.n555 B.n554 10.6151
R1458 B.n554 B.n551 10.6151
R1459 B.n551 B.n550 10.6151
R1460 B.n550 B.n547 10.6151
R1461 B.n547 B.n546 10.6151
R1462 B.n546 B.n543 10.6151
R1463 B.n543 B.n542 10.6151
R1464 B.n542 B.n539 10.6151
R1465 B.n539 B.n538 10.6151
R1466 B.n538 B.n535 10.6151
R1467 B.n535 B.n534 10.6151
R1468 B.n534 B.n531 10.6151
R1469 B.n531 B.n530 10.6151
R1470 B.n530 B.n527 10.6151
R1471 B.n527 B.n526 10.6151
R1472 B.n526 B.n523 10.6151
R1473 B.n523 B.n522 10.6151
R1474 B.n522 B.n519 10.6151
R1475 B.n519 B.n518 10.6151
R1476 B.n518 B.n515 10.6151
R1477 B.n515 B.n514 10.6151
R1478 B.n514 B.n511 10.6151
R1479 B.n511 B.n510 10.6151
R1480 B.n510 B.n507 10.6151
R1481 B.n507 B.n506 10.6151
R1482 B.n506 B.n503 10.6151
R1483 B.n503 B.n502 10.6151
R1484 B.n502 B.n499 10.6151
R1485 B.n499 B.n498 10.6151
R1486 B.n498 B.n495 10.6151
R1487 B.n495 B.n494 10.6151
R1488 B.n494 B.n491 10.6151
R1489 B.n491 B.n490 10.6151
R1490 B.n490 B.n487 10.6151
R1491 B.n487 B.n486 10.6151
R1492 B.n486 B.n483 10.6151
R1493 B.n483 B.n482 10.6151
R1494 B.n482 B.n479 10.6151
R1495 B.n479 B.n478 10.6151
R1496 B.n478 B.n475 10.6151
R1497 B.n475 B.n474 10.6151
R1498 B.n474 B.n471 10.6151
R1499 B.n471 B.n414 10.6151
R1500 B.n674 B.n414 10.6151
R1501 B.n680 B.n410 10.6151
R1502 B.n681 B.n680 10.6151
R1503 B.n682 B.n681 10.6151
R1504 B.n682 B.n402 10.6151
R1505 B.n692 B.n402 10.6151
R1506 B.n693 B.n692 10.6151
R1507 B.n694 B.n693 10.6151
R1508 B.n694 B.n394 10.6151
R1509 B.n704 B.n394 10.6151
R1510 B.n705 B.n704 10.6151
R1511 B.n706 B.n705 10.6151
R1512 B.n706 B.n386 10.6151
R1513 B.n716 B.n386 10.6151
R1514 B.n717 B.n716 10.6151
R1515 B.n718 B.n717 10.6151
R1516 B.n718 B.n378 10.6151
R1517 B.n728 B.n378 10.6151
R1518 B.n729 B.n728 10.6151
R1519 B.n730 B.n729 10.6151
R1520 B.n730 B.n370 10.6151
R1521 B.n741 B.n370 10.6151
R1522 B.n742 B.n741 10.6151
R1523 B.n743 B.n742 10.6151
R1524 B.n743 B.n363 10.6151
R1525 B.n753 B.n363 10.6151
R1526 B.n754 B.n753 10.6151
R1527 B.n755 B.n754 10.6151
R1528 B.n755 B.n355 10.6151
R1529 B.n765 B.n355 10.6151
R1530 B.n766 B.n765 10.6151
R1531 B.n767 B.n766 10.6151
R1532 B.n767 B.n347 10.6151
R1533 B.n777 B.n347 10.6151
R1534 B.n778 B.n777 10.6151
R1535 B.n779 B.n778 10.6151
R1536 B.n779 B.n339 10.6151
R1537 B.n790 B.n339 10.6151
R1538 B.n791 B.n790 10.6151
R1539 B.n792 B.n791 10.6151
R1540 B.n792 B.n0 10.6151
R1541 B.n931 B.n1 10.6151
R1542 B.n931 B.n930 10.6151
R1543 B.n930 B.n929 10.6151
R1544 B.n929 B.n10 10.6151
R1545 B.n923 B.n10 10.6151
R1546 B.n923 B.n922 10.6151
R1547 B.n922 B.n921 10.6151
R1548 B.n921 B.n17 10.6151
R1549 B.n915 B.n17 10.6151
R1550 B.n915 B.n914 10.6151
R1551 B.n914 B.n913 10.6151
R1552 B.n913 B.n24 10.6151
R1553 B.n907 B.n24 10.6151
R1554 B.n907 B.n906 10.6151
R1555 B.n906 B.n905 10.6151
R1556 B.n905 B.n31 10.6151
R1557 B.n899 B.n31 10.6151
R1558 B.n899 B.n898 10.6151
R1559 B.n898 B.n897 10.6151
R1560 B.n897 B.n37 10.6151
R1561 B.n891 B.n37 10.6151
R1562 B.n891 B.n890 10.6151
R1563 B.n890 B.n889 10.6151
R1564 B.n889 B.n45 10.6151
R1565 B.n883 B.n45 10.6151
R1566 B.n883 B.n882 10.6151
R1567 B.n882 B.n881 10.6151
R1568 B.n881 B.n52 10.6151
R1569 B.n875 B.n52 10.6151
R1570 B.n875 B.n874 10.6151
R1571 B.n874 B.n873 10.6151
R1572 B.n873 B.n59 10.6151
R1573 B.n867 B.n59 10.6151
R1574 B.n867 B.n866 10.6151
R1575 B.n866 B.n865 10.6151
R1576 B.n865 B.n66 10.6151
R1577 B.n859 B.n66 10.6151
R1578 B.n859 B.n858 10.6151
R1579 B.n858 B.n857 10.6151
R1580 B.n857 B.n73 10.6151
R1581 B.n224 B.n133 9.36635
R1582 B.n247 B.n130 9.36635
R1583 B.n581 B.n580 9.36635
R1584 B.n559 B.n558 9.36635
R1585 B.n745 B.t0 4.10607
R1586 B.t2 B.n345 4.10607
R1587 B.t3 B.n15 4.10607
R1588 B.n901 B.t1 4.10607
R1589 B.n937 B.n0 2.81026
R1590 B.n937 B.n1 2.81026
R1591 B.n227 B.n133 1.24928
R1592 B.n244 B.n130 1.24928
R1593 B.n580 B.n579 1.24928
R1594 B.n560 B.n559 1.24928
R1595 VN.n1 VN.t1 129.168
R1596 VN.n0 VN.t0 129.168
R1597 VN.n0 VN.t3 127.972
R1598 VN.n1 VN.t2 127.972
R1599 VN VN.n1 52.3444
R1600 VN VN.n0 2.30277
R1601 VDD2.n2 VDD2.n0 105.01
R1602 VDD2.n2 VDD2.n1 60.0025
R1603 VDD2.n1 VDD2.t2 1.46934
R1604 VDD2.n1 VDD2.t1 1.46934
R1605 VDD2.n0 VDD2.t0 1.46934
R1606 VDD2.n0 VDD2.t3 1.46934
R1607 VDD2 VDD2.n2 0.0586897
R1608 VTAIL.n586 VTAIL.n518 289.615
R1609 VTAIL.n68 VTAIL.n0 289.615
R1610 VTAIL.n142 VTAIL.n74 289.615
R1611 VTAIL.n216 VTAIL.n148 289.615
R1612 VTAIL.n512 VTAIL.n444 289.615
R1613 VTAIL.n438 VTAIL.n370 289.615
R1614 VTAIL.n364 VTAIL.n296 289.615
R1615 VTAIL.n290 VTAIL.n222 289.615
R1616 VTAIL.n543 VTAIL.n542 185
R1617 VTAIL.n545 VTAIL.n544 185
R1618 VTAIL.n538 VTAIL.n537 185
R1619 VTAIL.n551 VTAIL.n550 185
R1620 VTAIL.n553 VTAIL.n552 185
R1621 VTAIL.n534 VTAIL.n533 185
R1622 VTAIL.n560 VTAIL.n559 185
R1623 VTAIL.n561 VTAIL.n532 185
R1624 VTAIL.n563 VTAIL.n562 185
R1625 VTAIL.n530 VTAIL.n529 185
R1626 VTAIL.n569 VTAIL.n568 185
R1627 VTAIL.n571 VTAIL.n570 185
R1628 VTAIL.n526 VTAIL.n525 185
R1629 VTAIL.n577 VTAIL.n576 185
R1630 VTAIL.n579 VTAIL.n578 185
R1631 VTAIL.n522 VTAIL.n521 185
R1632 VTAIL.n585 VTAIL.n584 185
R1633 VTAIL.n587 VTAIL.n586 185
R1634 VTAIL.n25 VTAIL.n24 185
R1635 VTAIL.n27 VTAIL.n26 185
R1636 VTAIL.n20 VTAIL.n19 185
R1637 VTAIL.n33 VTAIL.n32 185
R1638 VTAIL.n35 VTAIL.n34 185
R1639 VTAIL.n16 VTAIL.n15 185
R1640 VTAIL.n42 VTAIL.n41 185
R1641 VTAIL.n43 VTAIL.n14 185
R1642 VTAIL.n45 VTAIL.n44 185
R1643 VTAIL.n12 VTAIL.n11 185
R1644 VTAIL.n51 VTAIL.n50 185
R1645 VTAIL.n53 VTAIL.n52 185
R1646 VTAIL.n8 VTAIL.n7 185
R1647 VTAIL.n59 VTAIL.n58 185
R1648 VTAIL.n61 VTAIL.n60 185
R1649 VTAIL.n4 VTAIL.n3 185
R1650 VTAIL.n67 VTAIL.n66 185
R1651 VTAIL.n69 VTAIL.n68 185
R1652 VTAIL.n99 VTAIL.n98 185
R1653 VTAIL.n101 VTAIL.n100 185
R1654 VTAIL.n94 VTAIL.n93 185
R1655 VTAIL.n107 VTAIL.n106 185
R1656 VTAIL.n109 VTAIL.n108 185
R1657 VTAIL.n90 VTAIL.n89 185
R1658 VTAIL.n116 VTAIL.n115 185
R1659 VTAIL.n117 VTAIL.n88 185
R1660 VTAIL.n119 VTAIL.n118 185
R1661 VTAIL.n86 VTAIL.n85 185
R1662 VTAIL.n125 VTAIL.n124 185
R1663 VTAIL.n127 VTAIL.n126 185
R1664 VTAIL.n82 VTAIL.n81 185
R1665 VTAIL.n133 VTAIL.n132 185
R1666 VTAIL.n135 VTAIL.n134 185
R1667 VTAIL.n78 VTAIL.n77 185
R1668 VTAIL.n141 VTAIL.n140 185
R1669 VTAIL.n143 VTAIL.n142 185
R1670 VTAIL.n173 VTAIL.n172 185
R1671 VTAIL.n175 VTAIL.n174 185
R1672 VTAIL.n168 VTAIL.n167 185
R1673 VTAIL.n181 VTAIL.n180 185
R1674 VTAIL.n183 VTAIL.n182 185
R1675 VTAIL.n164 VTAIL.n163 185
R1676 VTAIL.n190 VTAIL.n189 185
R1677 VTAIL.n191 VTAIL.n162 185
R1678 VTAIL.n193 VTAIL.n192 185
R1679 VTAIL.n160 VTAIL.n159 185
R1680 VTAIL.n199 VTAIL.n198 185
R1681 VTAIL.n201 VTAIL.n200 185
R1682 VTAIL.n156 VTAIL.n155 185
R1683 VTAIL.n207 VTAIL.n206 185
R1684 VTAIL.n209 VTAIL.n208 185
R1685 VTAIL.n152 VTAIL.n151 185
R1686 VTAIL.n215 VTAIL.n214 185
R1687 VTAIL.n217 VTAIL.n216 185
R1688 VTAIL.n513 VTAIL.n512 185
R1689 VTAIL.n511 VTAIL.n510 185
R1690 VTAIL.n448 VTAIL.n447 185
R1691 VTAIL.n505 VTAIL.n504 185
R1692 VTAIL.n503 VTAIL.n502 185
R1693 VTAIL.n452 VTAIL.n451 185
R1694 VTAIL.n497 VTAIL.n496 185
R1695 VTAIL.n495 VTAIL.n494 185
R1696 VTAIL.n456 VTAIL.n455 185
R1697 VTAIL.n460 VTAIL.n458 185
R1698 VTAIL.n489 VTAIL.n488 185
R1699 VTAIL.n487 VTAIL.n486 185
R1700 VTAIL.n462 VTAIL.n461 185
R1701 VTAIL.n481 VTAIL.n480 185
R1702 VTAIL.n479 VTAIL.n478 185
R1703 VTAIL.n466 VTAIL.n465 185
R1704 VTAIL.n473 VTAIL.n472 185
R1705 VTAIL.n471 VTAIL.n470 185
R1706 VTAIL.n439 VTAIL.n438 185
R1707 VTAIL.n437 VTAIL.n436 185
R1708 VTAIL.n374 VTAIL.n373 185
R1709 VTAIL.n431 VTAIL.n430 185
R1710 VTAIL.n429 VTAIL.n428 185
R1711 VTAIL.n378 VTAIL.n377 185
R1712 VTAIL.n423 VTAIL.n422 185
R1713 VTAIL.n421 VTAIL.n420 185
R1714 VTAIL.n382 VTAIL.n381 185
R1715 VTAIL.n386 VTAIL.n384 185
R1716 VTAIL.n415 VTAIL.n414 185
R1717 VTAIL.n413 VTAIL.n412 185
R1718 VTAIL.n388 VTAIL.n387 185
R1719 VTAIL.n407 VTAIL.n406 185
R1720 VTAIL.n405 VTAIL.n404 185
R1721 VTAIL.n392 VTAIL.n391 185
R1722 VTAIL.n399 VTAIL.n398 185
R1723 VTAIL.n397 VTAIL.n396 185
R1724 VTAIL.n365 VTAIL.n364 185
R1725 VTAIL.n363 VTAIL.n362 185
R1726 VTAIL.n300 VTAIL.n299 185
R1727 VTAIL.n357 VTAIL.n356 185
R1728 VTAIL.n355 VTAIL.n354 185
R1729 VTAIL.n304 VTAIL.n303 185
R1730 VTAIL.n349 VTAIL.n348 185
R1731 VTAIL.n347 VTAIL.n346 185
R1732 VTAIL.n308 VTAIL.n307 185
R1733 VTAIL.n312 VTAIL.n310 185
R1734 VTAIL.n341 VTAIL.n340 185
R1735 VTAIL.n339 VTAIL.n338 185
R1736 VTAIL.n314 VTAIL.n313 185
R1737 VTAIL.n333 VTAIL.n332 185
R1738 VTAIL.n331 VTAIL.n330 185
R1739 VTAIL.n318 VTAIL.n317 185
R1740 VTAIL.n325 VTAIL.n324 185
R1741 VTAIL.n323 VTAIL.n322 185
R1742 VTAIL.n291 VTAIL.n290 185
R1743 VTAIL.n289 VTAIL.n288 185
R1744 VTAIL.n226 VTAIL.n225 185
R1745 VTAIL.n283 VTAIL.n282 185
R1746 VTAIL.n281 VTAIL.n280 185
R1747 VTAIL.n230 VTAIL.n229 185
R1748 VTAIL.n275 VTAIL.n274 185
R1749 VTAIL.n273 VTAIL.n272 185
R1750 VTAIL.n234 VTAIL.n233 185
R1751 VTAIL.n238 VTAIL.n236 185
R1752 VTAIL.n267 VTAIL.n266 185
R1753 VTAIL.n265 VTAIL.n264 185
R1754 VTAIL.n240 VTAIL.n239 185
R1755 VTAIL.n259 VTAIL.n258 185
R1756 VTAIL.n257 VTAIL.n256 185
R1757 VTAIL.n244 VTAIL.n243 185
R1758 VTAIL.n251 VTAIL.n250 185
R1759 VTAIL.n249 VTAIL.n248 185
R1760 VTAIL.n541 VTAIL.t4 149.524
R1761 VTAIL.n23 VTAIL.t7 149.524
R1762 VTAIL.n97 VTAIL.t2 149.524
R1763 VTAIL.n171 VTAIL.t0 149.524
R1764 VTAIL.n469 VTAIL.t1 149.524
R1765 VTAIL.n395 VTAIL.t3 149.524
R1766 VTAIL.n321 VTAIL.t6 149.524
R1767 VTAIL.n247 VTAIL.t5 149.524
R1768 VTAIL.n544 VTAIL.n543 104.615
R1769 VTAIL.n544 VTAIL.n537 104.615
R1770 VTAIL.n551 VTAIL.n537 104.615
R1771 VTAIL.n552 VTAIL.n551 104.615
R1772 VTAIL.n552 VTAIL.n533 104.615
R1773 VTAIL.n560 VTAIL.n533 104.615
R1774 VTAIL.n561 VTAIL.n560 104.615
R1775 VTAIL.n562 VTAIL.n561 104.615
R1776 VTAIL.n562 VTAIL.n529 104.615
R1777 VTAIL.n569 VTAIL.n529 104.615
R1778 VTAIL.n570 VTAIL.n569 104.615
R1779 VTAIL.n570 VTAIL.n525 104.615
R1780 VTAIL.n577 VTAIL.n525 104.615
R1781 VTAIL.n578 VTAIL.n577 104.615
R1782 VTAIL.n578 VTAIL.n521 104.615
R1783 VTAIL.n585 VTAIL.n521 104.615
R1784 VTAIL.n586 VTAIL.n585 104.615
R1785 VTAIL.n26 VTAIL.n25 104.615
R1786 VTAIL.n26 VTAIL.n19 104.615
R1787 VTAIL.n33 VTAIL.n19 104.615
R1788 VTAIL.n34 VTAIL.n33 104.615
R1789 VTAIL.n34 VTAIL.n15 104.615
R1790 VTAIL.n42 VTAIL.n15 104.615
R1791 VTAIL.n43 VTAIL.n42 104.615
R1792 VTAIL.n44 VTAIL.n43 104.615
R1793 VTAIL.n44 VTAIL.n11 104.615
R1794 VTAIL.n51 VTAIL.n11 104.615
R1795 VTAIL.n52 VTAIL.n51 104.615
R1796 VTAIL.n52 VTAIL.n7 104.615
R1797 VTAIL.n59 VTAIL.n7 104.615
R1798 VTAIL.n60 VTAIL.n59 104.615
R1799 VTAIL.n60 VTAIL.n3 104.615
R1800 VTAIL.n67 VTAIL.n3 104.615
R1801 VTAIL.n68 VTAIL.n67 104.615
R1802 VTAIL.n100 VTAIL.n99 104.615
R1803 VTAIL.n100 VTAIL.n93 104.615
R1804 VTAIL.n107 VTAIL.n93 104.615
R1805 VTAIL.n108 VTAIL.n107 104.615
R1806 VTAIL.n108 VTAIL.n89 104.615
R1807 VTAIL.n116 VTAIL.n89 104.615
R1808 VTAIL.n117 VTAIL.n116 104.615
R1809 VTAIL.n118 VTAIL.n117 104.615
R1810 VTAIL.n118 VTAIL.n85 104.615
R1811 VTAIL.n125 VTAIL.n85 104.615
R1812 VTAIL.n126 VTAIL.n125 104.615
R1813 VTAIL.n126 VTAIL.n81 104.615
R1814 VTAIL.n133 VTAIL.n81 104.615
R1815 VTAIL.n134 VTAIL.n133 104.615
R1816 VTAIL.n134 VTAIL.n77 104.615
R1817 VTAIL.n141 VTAIL.n77 104.615
R1818 VTAIL.n142 VTAIL.n141 104.615
R1819 VTAIL.n174 VTAIL.n173 104.615
R1820 VTAIL.n174 VTAIL.n167 104.615
R1821 VTAIL.n181 VTAIL.n167 104.615
R1822 VTAIL.n182 VTAIL.n181 104.615
R1823 VTAIL.n182 VTAIL.n163 104.615
R1824 VTAIL.n190 VTAIL.n163 104.615
R1825 VTAIL.n191 VTAIL.n190 104.615
R1826 VTAIL.n192 VTAIL.n191 104.615
R1827 VTAIL.n192 VTAIL.n159 104.615
R1828 VTAIL.n199 VTAIL.n159 104.615
R1829 VTAIL.n200 VTAIL.n199 104.615
R1830 VTAIL.n200 VTAIL.n155 104.615
R1831 VTAIL.n207 VTAIL.n155 104.615
R1832 VTAIL.n208 VTAIL.n207 104.615
R1833 VTAIL.n208 VTAIL.n151 104.615
R1834 VTAIL.n215 VTAIL.n151 104.615
R1835 VTAIL.n216 VTAIL.n215 104.615
R1836 VTAIL.n512 VTAIL.n511 104.615
R1837 VTAIL.n511 VTAIL.n447 104.615
R1838 VTAIL.n504 VTAIL.n447 104.615
R1839 VTAIL.n504 VTAIL.n503 104.615
R1840 VTAIL.n503 VTAIL.n451 104.615
R1841 VTAIL.n496 VTAIL.n451 104.615
R1842 VTAIL.n496 VTAIL.n495 104.615
R1843 VTAIL.n495 VTAIL.n455 104.615
R1844 VTAIL.n460 VTAIL.n455 104.615
R1845 VTAIL.n488 VTAIL.n460 104.615
R1846 VTAIL.n488 VTAIL.n487 104.615
R1847 VTAIL.n487 VTAIL.n461 104.615
R1848 VTAIL.n480 VTAIL.n461 104.615
R1849 VTAIL.n480 VTAIL.n479 104.615
R1850 VTAIL.n479 VTAIL.n465 104.615
R1851 VTAIL.n472 VTAIL.n465 104.615
R1852 VTAIL.n472 VTAIL.n471 104.615
R1853 VTAIL.n438 VTAIL.n437 104.615
R1854 VTAIL.n437 VTAIL.n373 104.615
R1855 VTAIL.n430 VTAIL.n373 104.615
R1856 VTAIL.n430 VTAIL.n429 104.615
R1857 VTAIL.n429 VTAIL.n377 104.615
R1858 VTAIL.n422 VTAIL.n377 104.615
R1859 VTAIL.n422 VTAIL.n421 104.615
R1860 VTAIL.n421 VTAIL.n381 104.615
R1861 VTAIL.n386 VTAIL.n381 104.615
R1862 VTAIL.n414 VTAIL.n386 104.615
R1863 VTAIL.n414 VTAIL.n413 104.615
R1864 VTAIL.n413 VTAIL.n387 104.615
R1865 VTAIL.n406 VTAIL.n387 104.615
R1866 VTAIL.n406 VTAIL.n405 104.615
R1867 VTAIL.n405 VTAIL.n391 104.615
R1868 VTAIL.n398 VTAIL.n391 104.615
R1869 VTAIL.n398 VTAIL.n397 104.615
R1870 VTAIL.n364 VTAIL.n363 104.615
R1871 VTAIL.n363 VTAIL.n299 104.615
R1872 VTAIL.n356 VTAIL.n299 104.615
R1873 VTAIL.n356 VTAIL.n355 104.615
R1874 VTAIL.n355 VTAIL.n303 104.615
R1875 VTAIL.n348 VTAIL.n303 104.615
R1876 VTAIL.n348 VTAIL.n347 104.615
R1877 VTAIL.n347 VTAIL.n307 104.615
R1878 VTAIL.n312 VTAIL.n307 104.615
R1879 VTAIL.n340 VTAIL.n312 104.615
R1880 VTAIL.n340 VTAIL.n339 104.615
R1881 VTAIL.n339 VTAIL.n313 104.615
R1882 VTAIL.n332 VTAIL.n313 104.615
R1883 VTAIL.n332 VTAIL.n331 104.615
R1884 VTAIL.n331 VTAIL.n317 104.615
R1885 VTAIL.n324 VTAIL.n317 104.615
R1886 VTAIL.n324 VTAIL.n323 104.615
R1887 VTAIL.n290 VTAIL.n289 104.615
R1888 VTAIL.n289 VTAIL.n225 104.615
R1889 VTAIL.n282 VTAIL.n225 104.615
R1890 VTAIL.n282 VTAIL.n281 104.615
R1891 VTAIL.n281 VTAIL.n229 104.615
R1892 VTAIL.n274 VTAIL.n229 104.615
R1893 VTAIL.n274 VTAIL.n273 104.615
R1894 VTAIL.n273 VTAIL.n233 104.615
R1895 VTAIL.n238 VTAIL.n233 104.615
R1896 VTAIL.n266 VTAIL.n238 104.615
R1897 VTAIL.n266 VTAIL.n265 104.615
R1898 VTAIL.n265 VTAIL.n239 104.615
R1899 VTAIL.n258 VTAIL.n239 104.615
R1900 VTAIL.n258 VTAIL.n257 104.615
R1901 VTAIL.n257 VTAIL.n243 104.615
R1902 VTAIL.n250 VTAIL.n243 104.615
R1903 VTAIL.n250 VTAIL.n249 104.615
R1904 VTAIL.n543 VTAIL.t4 52.3082
R1905 VTAIL.n25 VTAIL.t7 52.3082
R1906 VTAIL.n99 VTAIL.t2 52.3082
R1907 VTAIL.n173 VTAIL.t0 52.3082
R1908 VTAIL.n471 VTAIL.t1 52.3082
R1909 VTAIL.n397 VTAIL.t3 52.3082
R1910 VTAIL.n323 VTAIL.t6 52.3082
R1911 VTAIL.n249 VTAIL.t5 52.3082
R1912 VTAIL.n591 VTAIL.n590 30.6338
R1913 VTAIL.n73 VTAIL.n72 30.6338
R1914 VTAIL.n147 VTAIL.n146 30.6338
R1915 VTAIL.n221 VTAIL.n220 30.6338
R1916 VTAIL.n517 VTAIL.n516 30.6338
R1917 VTAIL.n443 VTAIL.n442 30.6338
R1918 VTAIL.n369 VTAIL.n368 30.6338
R1919 VTAIL.n295 VTAIL.n294 30.6338
R1920 VTAIL.n591 VTAIL.n517 27.2117
R1921 VTAIL.n295 VTAIL.n221 27.2117
R1922 VTAIL.n563 VTAIL.n530 13.1884
R1923 VTAIL.n45 VTAIL.n12 13.1884
R1924 VTAIL.n119 VTAIL.n86 13.1884
R1925 VTAIL.n193 VTAIL.n160 13.1884
R1926 VTAIL.n458 VTAIL.n456 13.1884
R1927 VTAIL.n384 VTAIL.n382 13.1884
R1928 VTAIL.n310 VTAIL.n308 13.1884
R1929 VTAIL.n236 VTAIL.n234 13.1884
R1930 VTAIL.n564 VTAIL.n532 12.8005
R1931 VTAIL.n568 VTAIL.n567 12.8005
R1932 VTAIL.n46 VTAIL.n14 12.8005
R1933 VTAIL.n50 VTAIL.n49 12.8005
R1934 VTAIL.n120 VTAIL.n88 12.8005
R1935 VTAIL.n124 VTAIL.n123 12.8005
R1936 VTAIL.n194 VTAIL.n162 12.8005
R1937 VTAIL.n198 VTAIL.n197 12.8005
R1938 VTAIL.n494 VTAIL.n493 12.8005
R1939 VTAIL.n490 VTAIL.n489 12.8005
R1940 VTAIL.n420 VTAIL.n419 12.8005
R1941 VTAIL.n416 VTAIL.n415 12.8005
R1942 VTAIL.n346 VTAIL.n345 12.8005
R1943 VTAIL.n342 VTAIL.n341 12.8005
R1944 VTAIL.n272 VTAIL.n271 12.8005
R1945 VTAIL.n268 VTAIL.n267 12.8005
R1946 VTAIL.n559 VTAIL.n558 12.0247
R1947 VTAIL.n571 VTAIL.n528 12.0247
R1948 VTAIL.n41 VTAIL.n40 12.0247
R1949 VTAIL.n53 VTAIL.n10 12.0247
R1950 VTAIL.n115 VTAIL.n114 12.0247
R1951 VTAIL.n127 VTAIL.n84 12.0247
R1952 VTAIL.n189 VTAIL.n188 12.0247
R1953 VTAIL.n201 VTAIL.n158 12.0247
R1954 VTAIL.n497 VTAIL.n454 12.0247
R1955 VTAIL.n486 VTAIL.n459 12.0247
R1956 VTAIL.n423 VTAIL.n380 12.0247
R1957 VTAIL.n412 VTAIL.n385 12.0247
R1958 VTAIL.n349 VTAIL.n306 12.0247
R1959 VTAIL.n338 VTAIL.n311 12.0247
R1960 VTAIL.n275 VTAIL.n232 12.0247
R1961 VTAIL.n264 VTAIL.n237 12.0247
R1962 VTAIL.n557 VTAIL.n534 11.249
R1963 VTAIL.n572 VTAIL.n526 11.249
R1964 VTAIL.n39 VTAIL.n16 11.249
R1965 VTAIL.n54 VTAIL.n8 11.249
R1966 VTAIL.n113 VTAIL.n90 11.249
R1967 VTAIL.n128 VTAIL.n82 11.249
R1968 VTAIL.n187 VTAIL.n164 11.249
R1969 VTAIL.n202 VTAIL.n156 11.249
R1970 VTAIL.n498 VTAIL.n452 11.249
R1971 VTAIL.n485 VTAIL.n462 11.249
R1972 VTAIL.n424 VTAIL.n378 11.249
R1973 VTAIL.n411 VTAIL.n388 11.249
R1974 VTAIL.n350 VTAIL.n304 11.249
R1975 VTAIL.n337 VTAIL.n314 11.249
R1976 VTAIL.n276 VTAIL.n230 11.249
R1977 VTAIL.n263 VTAIL.n240 11.249
R1978 VTAIL.n554 VTAIL.n553 10.4732
R1979 VTAIL.n576 VTAIL.n575 10.4732
R1980 VTAIL.n36 VTAIL.n35 10.4732
R1981 VTAIL.n58 VTAIL.n57 10.4732
R1982 VTAIL.n110 VTAIL.n109 10.4732
R1983 VTAIL.n132 VTAIL.n131 10.4732
R1984 VTAIL.n184 VTAIL.n183 10.4732
R1985 VTAIL.n206 VTAIL.n205 10.4732
R1986 VTAIL.n502 VTAIL.n501 10.4732
R1987 VTAIL.n482 VTAIL.n481 10.4732
R1988 VTAIL.n428 VTAIL.n427 10.4732
R1989 VTAIL.n408 VTAIL.n407 10.4732
R1990 VTAIL.n354 VTAIL.n353 10.4732
R1991 VTAIL.n334 VTAIL.n333 10.4732
R1992 VTAIL.n280 VTAIL.n279 10.4732
R1993 VTAIL.n260 VTAIL.n259 10.4732
R1994 VTAIL.n542 VTAIL.n541 10.2747
R1995 VTAIL.n24 VTAIL.n23 10.2747
R1996 VTAIL.n98 VTAIL.n97 10.2747
R1997 VTAIL.n172 VTAIL.n171 10.2747
R1998 VTAIL.n470 VTAIL.n469 10.2747
R1999 VTAIL.n396 VTAIL.n395 10.2747
R2000 VTAIL.n322 VTAIL.n321 10.2747
R2001 VTAIL.n248 VTAIL.n247 10.2747
R2002 VTAIL.n550 VTAIL.n536 9.69747
R2003 VTAIL.n579 VTAIL.n524 9.69747
R2004 VTAIL.n32 VTAIL.n18 9.69747
R2005 VTAIL.n61 VTAIL.n6 9.69747
R2006 VTAIL.n106 VTAIL.n92 9.69747
R2007 VTAIL.n135 VTAIL.n80 9.69747
R2008 VTAIL.n180 VTAIL.n166 9.69747
R2009 VTAIL.n209 VTAIL.n154 9.69747
R2010 VTAIL.n505 VTAIL.n450 9.69747
R2011 VTAIL.n478 VTAIL.n464 9.69747
R2012 VTAIL.n431 VTAIL.n376 9.69747
R2013 VTAIL.n404 VTAIL.n390 9.69747
R2014 VTAIL.n357 VTAIL.n302 9.69747
R2015 VTAIL.n330 VTAIL.n316 9.69747
R2016 VTAIL.n283 VTAIL.n228 9.69747
R2017 VTAIL.n256 VTAIL.n242 9.69747
R2018 VTAIL.n590 VTAIL.n589 9.45567
R2019 VTAIL.n72 VTAIL.n71 9.45567
R2020 VTAIL.n146 VTAIL.n145 9.45567
R2021 VTAIL.n220 VTAIL.n219 9.45567
R2022 VTAIL.n516 VTAIL.n515 9.45567
R2023 VTAIL.n442 VTAIL.n441 9.45567
R2024 VTAIL.n368 VTAIL.n367 9.45567
R2025 VTAIL.n294 VTAIL.n293 9.45567
R2026 VTAIL.n589 VTAIL.n588 9.3005
R2027 VTAIL.n583 VTAIL.n582 9.3005
R2028 VTAIL.n581 VTAIL.n580 9.3005
R2029 VTAIL.n524 VTAIL.n523 9.3005
R2030 VTAIL.n575 VTAIL.n574 9.3005
R2031 VTAIL.n573 VTAIL.n572 9.3005
R2032 VTAIL.n528 VTAIL.n527 9.3005
R2033 VTAIL.n567 VTAIL.n566 9.3005
R2034 VTAIL.n540 VTAIL.n539 9.3005
R2035 VTAIL.n547 VTAIL.n546 9.3005
R2036 VTAIL.n549 VTAIL.n548 9.3005
R2037 VTAIL.n536 VTAIL.n535 9.3005
R2038 VTAIL.n555 VTAIL.n554 9.3005
R2039 VTAIL.n557 VTAIL.n556 9.3005
R2040 VTAIL.n558 VTAIL.n531 9.3005
R2041 VTAIL.n565 VTAIL.n564 9.3005
R2042 VTAIL.n520 VTAIL.n519 9.3005
R2043 VTAIL.n71 VTAIL.n70 9.3005
R2044 VTAIL.n65 VTAIL.n64 9.3005
R2045 VTAIL.n63 VTAIL.n62 9.3005
R2046 VTAIL.n6 VTAIL.n5 9.3005
R2047 VTAIL.n57 VTAIL.n56 9.3005
R2048 VTAIL.n55 VTAIL.n54 9.3005
R2049 VTAIL.n10 VTAIL.n9 9.3005
R2050 VTAIL.n49 VTAIL.n48 9.3005
R2051 VTAIL.n22 VTAIL.n21 9.3005
R2052 VTAIL.n29 VTAIL.n28 9.3005
R2053 VTAIL.n31 VTAIL.n30 9.3005
R2054 VTAIL.n18 VTAIL.n17 9.3005
R2055 VTAIL.n37 VTAIL.n36 9.3005
R2056 VTAIL.n39 VTAIL.n38 9.3005
R2057 VTAIL.n40 VTAIL.n13 9.3005
R2058 VTAIL.n47 VTAIL.n46 9.3005
R2059 VTAIL.n2 VTAIL.n1 9.3005
R2060 VTAIL.n145 VTAIL.n144 9.3005
R2061 VTAIL.n139 VTAIL.n138 9.3005
R2062 VTAIL.n137 VTAIL.n136 9.3005
R2063 VTAIL.n80 VTAIL.n79 9.3005
R2064 VTAIL.n131 VTAIL.n130 9.3005
R2065 VTAIL.n129 VTAIL.n128 9.3005
R2066 VTAIL.n84 VTAIL.n83 9.3005
R2067 VTAIL.n123 VTAIL.n122 9.3005
R2068 VTAIL.n96 VTAIL.n95 9.3005
R2069 VTAIL.n103 VTAIL.n102 9.3005
R2070 VTAIL.n105 VTAIL.n104 9.3005
R2071 VTAIL.n92 VTAIL.n91 9.3005
R2072 VTAIL.n111 VTAIL.n110 9.3005
R2073 VTAIL.n113 VTAIL.n112 9.3005
R2074 VTAIL.n114 VTAIL.n87 9.3005
R2075 VTAIL.n121 VTAIL.n120 9.3005
R2076 VTAIL.n76 VTAIL.n75 9.3005
R2077 VTAIL.n219 VTAIL.n218 9.3005
R2078 VTAIL.n213 VTAIL.n212 9.3005
R2079 VTAIL.n211 VTAIL.n210 9.3005
R2080 VTAIL.n154 VTAIL.n153 9.3005
R2081 VTAIL.n205 VTAIL.n204 9.3005
R2082 VTAIL.n203 VTAIL.n202 9.3005
R2083 VTAIL.n158 VTAIL.n157 9.3005
R2084 VTAIL.n197 VTAIL.n196 9.3005
R2085 VTAIL.n170 VTAIL.n169 9.3005
R2086 VTAIL.n177 VTAIL.n176 9.3005
R2087 VTAIL.n179 VTAIL.n178 9.3005
R2088 VTAIL.n166 VTAIL.n165 9.3005
R2089 VTAIL.n185 VTAIL.n184 9.3005
R2090 VTAIL.n187 VTAIL.n186 9.3005
R2091 VTAIL.n188 VTAIL.n161 9.3005
R2092 VTAIL.n195 VTAIL.n194 9.3005
R2093 VTAIL.n150 VTAIL.n149 9.3005
R2094 VTAIL.n468 VTAIL.n467 9.3005
R2095 VTAIL.n475 VTAIL.n474 9.3005
R2096 VTAIL.n477 VTAIL.n476 9.3005
R2097 VTAIL.n464 VTAIL.n463 9.3005
R2098 VTAIL.n483 VTAIL.n482 9.3005
R2099 VTAIL.n485 VTAIL.n484 9.3005
R2100 VTAIL.n459 VTAIL.n457 9.3005
R2101 VTAIL.n491 VTAIL.n490 9.3005
R2102 VTAIL.n515 VTAIL.n514 9.3005
R2103 VTAIL.n446 VTAIL.n445 9.3005
R2104 VTAIL.n509 VTAIL.n508 9.3005
R2105 VTAIL.n507 VTAIL.n506 9.3005
R2106 VTAIL.n450 VTAIL.n449 9.3005
R2107 VTAIL.n501 VTAIL.n500 9.3005
R2108 VTAIL.n499 VTAIL.n498 9.3005
R2109 VTAIL.n454 VTAIL.n453 9.3005
R2110 VTAIL.n493 VTAIL.n492 9.3005
R2111 VTAIL.n394 VTAIL.n393 9.3005
R2112 VTAIL.n401 VTAIL.n400 9.3005
R2113 VTAIL.n403 VTAIL.n402 9.3005
R2114 VTAIL.n390 VTAIL.n389 9.3005
R2115 VTAIL.n409 VTAIL.n408 9.3005
R2116 VTAIL.n411 VTAIL.n410 9.3005
R2117 VTAIL.n385 VTAIL.n383 9.3005
R2118 VTAIL.n417 VTAIL.n416 9.3005
R2119 VTAIL.n441 VTAIL.n440 9.3005
R2120 VTAIL.n372 VTAIL.n371 9.3005
R2121 VTAIL.n435 VTAIL.n434 9.3005
R2122 VTAIL.n433 VTAIL.n432 9.3005
R2123 VTAIL.n376 VTAIL.n375 9.3005
R2124 VTAIL.n427 VTAIL.n426 9.3005
R2125 VTAIL.n425 VTAIL.n424 9.3005
R2126 VTAIL.n380 VTAIL.n379 9.3005
R2127 VTAIL.n419 VTAIL.n418 9.3005
R2128 VTAIL.n320 VTAIL.n319 9.3005
R2129 VTAIL.n327 VTAIL.n326 9.3005
R2130 VTAIL.n329 VTAIL.n328 9.3005
R2131 VTAIL.n316 VTAIL.n315 9.3005
R2132 VTAIL.n335 VTAIL.n334 9.3005
R2133 VTAIL.n337 VTAIL.n336 9.3005
R2134 VTAIL.n311 VTAIL.n309 9.3005
R2135 VTAIL.n343 VTAIL.n342 9.3005
R2136 VTAIL.n367 VTAIL.n366 9.3005
R2137 VTAIL.n298 VTAIL.n297 9.3005
R2138 VTAIL.n361 VTAIL.n360 9.3005
R2139 VTAIL.n359 VTAIL.n358 9.3005
R2140 VTAIL.n302 VTAIL.n301 9.3005
R2141 VTAIL.n353 VTAIL.n352 9.3005
R2142 VTAIL.n351 VTAIL.n350 9.3005
R2143 VTAIL.n306 VTAIL.n305 9.3005
R2144 VTAIL.n345 VTAIL.n344 9.3005
R2145 VTAIL.n246 VTAIL.n245 9.3005
R2146 VTAIL.n253 VTAIL.n252 9.3005
R2147 VTAIL.n255 VTAIL.n254 9.3005
R2148 VTAIL.n242 VTAIL.n241 9.3005
R2149 VTAIL.n261 VTAIL.n260 9.3005
R2150 VTAIL.n263 VTAIL.n262 9.3005
R2151 VTAIL.n237 VTAIL.n235 9.3005
R2152 VTAIL.n269 VTAIL.n268 9.3005
R2153 VTAIL.n293 VTAIL.n292 9.3005
R2154 VTAIL.n224 VTAIL.n223 9.3005
R2155 VTAIL.n287 VTAIL.n286 9.3005
R2156 VTAIL.n285 VTAIL.n284 9.3005
R2157 VTAIL.n228 VTAIL.n227 9.3005
R2158 VTAIL.n279 VTAIL.n278 9.3005
R2159 VTAIL.n277 VTAIL.n276 9.3005
R2160 VTAIL.n232 VTAIL.n231 9.3005
R2161 VTAIL.n271 VTAIL.n270 9.3005
R2162 VTAIL.n549 VTAIL.n538 8.92171
R2163 VTAIL.n580 VTAIL.n522 8.92171
R2164 VTAIL.n31 VTAIL.n20 8.92171
R2165 VTAIL.n62 VTAIL.n4 8.92171
R2166 VTAIL.n105 VTAIL.n94 8.92171
R2167 VTAIL.n136 VTAIL.n78 8.92171
R2168 VTAIL.n179 VTAIL.n168 8.92171
R2169 VTAIL.n210 VTAIL.n152 8.92171
R2170 VTAIL.n506 VTAIL.n448 8.92171
R2171 VTAIL.n477 VTAIL.n466 8.92171
R2172 VTAIL.n432 VTAIL.n374 8.92171
R2173 VTAIL.n403 VTAIL.n392 8.92171
R2174 VTAIL.n358 VTAIL.n300 8.92171
R2175 VTAIL.n329 VTAIL.n318 8.92171
R2176 VTAIL.n284 VTAIL.n226 8.92171
R2177 VTAIL.n255 VTAIL.n244 8.92171
R2178 VTAIL.n546 VTAIL.n545 8.14595
R2179 VTAIL.n584 VTAIL.n583 8.14595
R2180 VTAIL.n28 VTAIL.n27 8.14595
R2181 VTAIL.n66 VTAIL.n65 8.14595
R2182 VTAIL.n102 VTAIL.n101 8.14595
R2183 VTAIL.n140 VTAIL.n139 8.14595
R2184 VTAIL.n176 VTAIL.n175 8.14595
R2185 VTAIL.n214 VTAIL.n213 8.14595
R2186 VTAIL.n510 VTAIL.n509 8.14595
R2187 VTAIL.n474 VTAIL.n473 8.14595
R2188 VTAIL.n436 VTAIL.n435 8.14595
R2189 VTAIL.n400 VTAIL.n399 8.14595
R2190 VTAIL.n362 VTAIL.n361 8.14595
R2191 VTAIL.n326 VTAIL.n325 8.14595
R2192 VTAIL.n288 VTAIL.n287 8.14595
R2193 VTAIL.n252 VTAIL.n251 8.14595
R2194 VTAIL.n542 VTAIL.n540 7.3702
R2195 VTAIL.n587 VTAIL.n520 7.3702
R2196 VTAIL.n590 VTAIL.n518 7.3702
R2197 VTAIL.n24 VTAIL.n22 7.3702
R2198 VTAIL.n69 VTAIL.n2 7.3702
R2199 VTAIL.n72 VTAIL.n0 7.3702
R2200 VTAIL.n98 VTAIL.n96 7.3702
R2201 VTAIL.n143 VTAIL.n76 7.3702
R2202 VTAIL.n146 VTAIL.n74 7.3702
R2203 VTAIL.n172 VTAIL.n170 7.3702
R2204 VTAIL.n217 VTAIL.n150 7.3702
R2205 VTAIL.n220 VTAIL.n148 7.3702
R2206 VTAIL.n516 VTAIL.n444 7.3702
R2207 VTAIL.n513 VTAIL.n446 7.3702
R2208 VTAIL.n470 VTAIL.n468 7.3702
R2209 VTAIL.n442 VTAIL.n370 7.3702
R2210 VTAIL.n439 VTAIL.n372 7.3702
R2211 VTAIL.n396 VTAIL.n394 7.3702
R2212 VTAIL.n368 VTAIL.n296 7.3702
R2213 VTAIL.n365 VTAIL.n298 7.3702
R2214 VTAIL.n322 VTAIL.n320 7.3702
R2215 VTAIL.n294 VTAIL.n222 7.3702
R2216 VTAIL.n291 VTAIL.n224 7.3702
R2217 VTAIL.n248 VTAIL.n246 7.3702
R2218 VTAIL.n588 VTAIL.n587 6.59444
R2219 VTAIL.n588 VTAIL.n518 6.59444
R2220 VTAIL.n70 VTAIL.n69 6.59444
R2221 VTAIL.n70 VTAIL.n0 6.59444
R2222 VTAIL.n144 VTAIL.n143 6.59444
R2223 VTAIL.n144 VTAIL.n74 6.59444
R2224 VTAIL.n218 VTAIL.n217 6.59444
R2225 VTAIL.n218 VTAIL.n148 6.59444
R2226 VTAIL.n514 VTAIL.n444 6.59444
R2227 VTAIL.n514 VTAIL.n513 6.59444
R2228 VTAIL.n440 VTAIL.n370 6.59444
R2229 VTAIL.n440 VTAIL.n439 6.59444
R2230 VTAIL.n366 VTAIL.n296 6.59444
R2231 VTAIL.n366 VTAIL.n365 6.59444
R2232 VTAIL.n292 VTAIL.n222 6.59444
R2233 VTAIL.n292 VTAIL.n291 6.59444
R2234 VTAIL.n545 VTAIL.n540 5.81868
R2235 VTAIL.n584 VTAIL.n520 5.81868
R2236 VTAIL.n27 VTAIL.n22 5.81868
R2237 VTAIL.n66 VTAIL.n2 5.81868
R2238 VTAIL.n101 VTAIL.n96 5.81868
R2239 VTAIL.n140 VTAIL.n76 5.81868
R2240 VTAIL.n175 VTAIL.n170 5.81868
R2241 VTAIL.n214 VTAIL.n150 5.81868
R2242 VTAIL.n510 VTAIL.n446 5.81868
R2243 VTAIL.n473 VTAIL.n468 5.81868
R2244 VTAIL.n436 VTAIL.n372 5.81868
R2245 VTAIL.n399 VTAIL.n394 5.81868
R2246 VTAIL.n362 VTAIL.n298 5.81868
R2247 VTAIL.n325 VTAIL.n320 5.81868
R2248 VTAIL.n288 VTAIL.n224 5.81868
R2249 VTAIL.n251 VTAIL.n246 5.81868
R2250 VTAIL.n546 VTAIL.n538 5.04292
R2251 VTAIL.n583 VTAIL.n522 5.04292
R2252 VTAIL.n28 VTAIL.n20 5.04292
R2253 VTAIL.n65 VTAIL.n4 5.04292
R2254 VTAIL.n102 VTAIL.n94 5.04292
R2255 VTAIL.n139 VTAIL.n78 5.04292
R2256 VTAIL.n176 VTAIL.n168 5.04292
R2257 VTAIL.n213 VTAIL.n152 5.04292
R2258 VTAIL.n509 VTAIL.n448 5.04292
R2259 VTAIL.n474 VTAIL.n466 5.04292
R2260 VTAIL.n435 VTAIL.n374 5.04292
R2261 VTAIL.n400 VTAIL.n392 5.04292
R2262 VTAIL.n361 VTAIL.n300 5.04292
R2263 VTAIL.n326 VTAIL.n318 5.04292
R2264 VTAIL.n287 VTAIL.n226 5.04292
R2265 VTAIL.n252 VTAIL.n244 5.04292
R2266 VTAIL.n550 VTAIL.n549 4.26717
R2267 VTAIL.n580 VTAIL.n579 4.26717
R2268 VTAIL.n32 VTAIL.n31 4.26717
R2269 VTAIL.n62 VTAIL.n61 4.26717
R2270 VTAIL.n106 VTAIL.n105 4.26717
R2271 VTAIL.n136 VTAIL.n135 4.26717
R2272 VTAIL.n180 VTAIL.n179 4.26717
R2273 VTAIL.n210 VTAIL.n209 4.26717
R2274 VTAIL.n506 VTAIL.n505 4.26717
R2275 VTAIL.n478 VTAIL.n477 4.26717
R2276 VTAIL.n432 VTAIL.n431 4.26717
R2277 VTAIL.n404 VTAIL.n403 4.26717
R2278 VTAIL.n358 VTAIL.n357 4.26717
R2279 VTAIL.n330 VTAIL.n329 4.26717
R2280 VTAIL.n284 VTAIL.n283 4.26717
R2281 VTAIL.n256 VTAIL.n255 4.26717
R2282 VTAIL.n553 VTAIL.n536 3.49141
R2283 VTAIL.n576 VTAIL.n524 3.49141
R2284 VTAIL.n35 VTAIL.n18 3.49141
R2285 VTAIL.n58 VTAIL.n6 3.49141
R2286 VTAIL.n109 VTAIL.n92 3.49141
R2287 VTAIL.n132 VTAIL.n80 3.49141
R2288 VTAIL.n183 VTAIL.n166 3.49141
R2289 VTAIL.n206 VTAIL.n154 3.49141
R2290 VTAIL.n502 VTAIL.n450 3.49141
R2291 VTAIL.n481 VTAIL.n464 3.49141
R2292 VTAIL.n428 VTAIL.n376 3.49141
R2293 VTAIL.n407 VTAIL.n390 3.49141
R2294 VTAIL.n354 VTAIL.n302 3.49141
R2295 VTAIL.n333 VTAIL.n316 3.49141
R2296 VTAIL.n280 VTAIL.n228 3.49141
R2297 VTAIL.n259 VTAIL.n242 3.49141
R2298 VTAIL.n369 VTAIL.n295 3.22464
R2299 VTAIL.n517 VTAIL.n443 3.22464
R2300 VTAIL.n221 VTAIL.n147 3.22464
R2301 VTAIL.n541 VTAIL.n539 2.84303
R2302 VTAIL.n23 VTAIL.n21 2.84303
R2303 VTAIL.n97 VTAIL.n95 2.84303
R2304 VTAIL.n171 VTAIL.n169 2.84303
R2305 VTAIL.n469 VTAIL.n467 2.84303
R2306 VTAIL.n395 VTAIL.n393 2.84303
R2307 VTAIL.n321 VTAIL.n319 2.84303
R2308 VTAIL.n247 VTAIL.n245 2.84303
R2309 VTAIL.n554 VTAIL.n534 2.71565
R2310 VTAIL.n575 VTAIL.n526 2.71565
R2311 VTAIL.n36 VTAIL.n16 2.71565
R2312 VTAIL.n57 VTAIL.n8 2.71565
R2313 VTAIL.n110 VTAIL.n90 2.71565
R2314 VTAIL.n131 VTAIL.n82 2.71565
R2315 VTAIL.n184 VTAIL.n164 2.71565
R2316 VTAIL.n205 VTAIL.n156 2.71565
R2317 VTAIL.n501 VTAIL.n452 2.71565
R2318 VTAIL.n482 VTAIL.n462 2.71565
R2319 VTAIL.n427 VTAIL.n378 2.71565
R2320 VTAIL.n408 VTAIL.n388 2.71565
R2321 VTAIL.n353 VTAIL.n304 2.71565
R2322 VTAIL.n334 VTAIL.n314 2.71565
R2323 VTAIL.n279 VTAIL.n230 2.71565
R2324 VTAIL.n260 VTAIL.n240 2.71565
R2325 VTAIL.n559 VTAIL.n557 1.93989
R2326 VTAIL.n572 VTAIL.n571 1.93989
R2327 VTAIL.n41 VTAIL.n39 1.93989
R2328 VTAIL.n54 VTAIL.n53 1.93989
R2329 VTAIL.n115 VTAIL.n113 1.93989
R2330 VTAIL.n128 VTAIL.n127 1.93989
R2331 VTAIL.n189 VTAIL.n187 1.93989
R2332 VTAIL.n202 VTAIL.n201 1.93989
R2333 VTAIL.n498 VTAIL.n497 1.93989
R2334 VTAIL.n486 VTAIL.n485 1.93989
R2335 VTAIL.n424 VTAIL.n423 1.93989
R2336 VTAIL.n412 VTAIL.n411 1.93989
R2337 VTAIL.n350 VTAIL.n349 1.93989
R2338 VTAIL.n338 VTAIL.n337 1.93989
R2339 VTAIL.n276 VTAIL.n275 1.93989
R2340 VTAIL.n264 VTAIL.n263 1.93989
R2341 VTAIL VTAIL.n73 1.67076
R2342 VTAIL VTAIL.n591 1.55438
R2343 VTAIL.n558 VTAIL.n532 1.16414
R2344 VTAIL.n568 VTAIL.n528 1.16414
R2345 VTAIL.n40 VTAIL.n14 1.16414
R2346 VTAIL.n50 VTAIL.n10 1.16414
R2347 VTAIL.n114 VTAIL.n88 1.16414
R2348 VTAIL.n124 VTAIL.n84 1.16414
R2349 VTAIL.n188 VTAIL.n162 1.16414
R2350 VTAIL.n198 VTAIL.n158 1.16414
R2351 VTAIL.n494 VTAIL.n454 1.16414
R2352 VTAIL.n489 VTAIL.n459 1.16414
R2353 VTAIL.n420 VTAIL.n380 1.16414
R2354 VTAIL.n415 VTAIL.n385 1.16414
R2355 VTAIL.n346 VTAIL.n306 1.16414
R2356 VTAIL.n341 VTAIL.n311 1.16414
R2357 VTAIL.n272 VTAIL.n232 1.16414
R2358 VTAIL.n267 VTAIL.n237 1.16414
R2359 VTAIL.n443 VTAIL.n369 0.470328
R2360 VTAIL.n147 VTAIL.n73 0.470328
R2361 VTAIL.n564 VTAIL.n563 0.388379
R2362 VTAIL.n567 VTAIL.n530 0.388379
R2363 VTAIL.n46 VTAIL.n45 0.388379
R2364 VTAIL.n49 VTAIL.n12 0.388379
R2365 VTAIL.n120 VTAIL.n119 0.388379
R2366 VTAIL.n123 VTAIL.n86 0.388379
R2367 VTAIL.n194 VTAIL.n193 0.388379
R2368 VTAIL.n197 VTAIL.n160 0.388379
R2369 VTAIL.n493 VTAIL.n456 0.388379
R2370 VTAIL.n490 VTAIL.n458 0.388379
R2371 VTAIL.n419 VTAIL.n382 0.388379
R2372 VTAIL.n416 VTAIL.n384 0.388379
R2373 VTAIL.n345 VTAIL.n308 0.388379
R2374 VTAIL.n342 VTAIL.n310 0.388379
R2375 VTAIL.n271 VTAIL.n234 0.388379
R2376 VTAIL.n268 VTAIL.n236 0.388379
R2377 VTAIL.n547 VTAIL.n539 0.155672
R2378 VTAIL.n548 VTAIL.n547 0.155672
R2379 VTAIL.n548 VTAIL.n535 0.155672
R2380 VTAIL.n555 VTAIL.n535 0.155672
R2381 VTAIL.n556 VTAIL.n555 0.155672
R2382 VTAIL.n556 VTAIL.n531 0.155672
R2383 VTAIL.n565 VTAIL.n531 0.155672
R2384 VTAIL.n566 VTAIL.n565 0.155672
R2385 VTAIL.n566 VTAIL.n527 0.155672
R2386 VTAIL.n573 VTAIL.n527 0.155672
R2387 VTAIL.n574 VTAIL.n573 0.155672
R2388 VTAIL.n574 VTAIL.n523 0.155672
R2389 VTAIL.n581 VTAIL.n523 0.155672
R2390 VTAIL.n582 VTAIL.n581 0.155672
R2391 VTAIL.n582 VTAIL.n519 0.155672
R2392 VTAIL.n589 VTAIL.n519 0.155672
R2393 VTAIL.n29 VTAIL.n21 0.155672
R2394 VTAIL.n30 VTAIL.n29 0.155672
R2395 VTAIL.n30 VTAIL.n17 0.155672
R2396 VTAIL.n37 VTAIL.n17 0.155672
R2397 VTAIL.n38 VTAIL.n37 0.155672
R2398 VTAIL.n38 VTAIL.n13 0.155672
R2399 VTAIL.n47 VTAIL.n13 0.155672
R2400 VTAIL.n48 VTAIL.n47 0.155672
R2401 VTAIL.n48 VTAIL.n9 0.155672
R2402 VTAIL.n55 VTAIL.n9 0.155672
R2403 VTAIL.n56 VTAIL.n55 0.155672
R2404 VTAIL.n56 VTAIL.n5 0.155672
R2405 VTAIL.n63 VTAIL.n5 0.155672
R2406 VTAIL.n64 VTAIL.n63 0.155672
R2407 VTAIL.n64 VTAIL.n1 0.155672
R2408 VTAIL.n71 VTAIL.n1 0.155672
R2409 VTAIL.n103 VTAIL.n95 0.155672
R2410 VTAIL.n104 VTAIL.n103 0.155672
R2411 VTAIL.n104 VTAIL.n91 0.155672
R2412 VTAIL.n111 VTAIL.n91 0.155672
R2413 VTAIL.n112 VTAIL.n111 0.155672
R2414 VTAIL.n112 VTAIL.n87 0.155672
R2415 VTAIL.n121 VTAIL.n87 0.155672
R2416 VTAIL.n122 VTAIL.n121 0.155672
R2417 VTAIL.n122 VTAIL.n83 0.155672
R2418 VTAIL.n129 VTAIL.n83 0.155672
R2419 VTAIL.n130 VTAIL.n129 0.155672
R2420 VTAIL.n130 VTAIL.n79 0.155672
R2421 VTAIL.n137 VTAIL.n79 0.155672
R2422 VTAIL.n138 VTAIL.n137 0.155672
R2423 VTAIL.n138 VTAIL.n75 0.155672
R2424 VTAIL.n145 VTAIL.n75 0.155672
R2425 VTAIL.n177 VTAIL.n169 0.155672
R2426 VTAIL.n178 VTAIL.n177 0.155672
R2427 VTAIL.n178 VTAIL.n165 0.155672
R2428 VTAIL.n185 VTAIL.n165 0.155672
R2429 VTAIL.n186 VTAIL.n185 0.155672
R2430 VTAIL.n186 VTAIL.n161 0.155672
R2431 VTAIL.n195 VTAIL.n161 0.155672
R2432 VTAIL.n196 VTAIL.n195 0.155672
R2433 VTAIL.n196 VTAIL.n157 0.155672
R2434 VTAIL.n203 VTAIL.n157 0.155672
R2435 VTAIL.n204 VTAIL.n203 0.155672
R2436 VTAIL.n204 VTAIL.n153 0.155672
R2437 VTAIL.n211 VTAIL.n153 0.155672
R2438 VTAIL.n212 VTAIL.n211 0.155672
R2439 VTAIL.n212 VTAIL.n149 0.155672
R2440 VTAIL.n219 VTAIL.n149 0.155672
R2441 VTAIL.n515 VTAIL.n445 0.155672
R2442 VTAIL.n508 VTAIL.n445 0.155672
R2443 VTAIL.n508 VTAIL.n507 0.155672
R2444 VTAIL.n507 VTAIL.n449 0.155672
R2445 VTAIL.n500 VTAIL.n449 0.155672
R2446 VTAIL.n500 VTAIL.n499 0.155672
R2447 VTAIL.n499 VTAIL.n453 0.155672
R2448 VTAIL.n492 VTAIL.n453 0.155672
R2449 VTAIL.n492 VTAIL.n491 0.155672
R2450 VTAIL.n491 VTAIL.n457 0.155672
R2451 VTAIL.n484 VTAIL.n457 0.155672
R2452 VTAIL.n484 VTAIL.n483 0.155672
R2453 VTAIL.n483 VTAIL.n463 0.155672
R2454 VTAIL.n476 VTAIL.n463 0.155672
R2455 VTAIL.n476 VTAIL.n475 0.155672
R2456 VTAIL.n475 VTAIL.n467 0.155672
R2457 VTAIL.n441 VTAIL.n371 0.155672
R2458 VTAIL.n434 VTAIL.n371 0.155672
R2459 VTAIL.n434 VTAIL.n433 0.155672
R2460 VTAIL.n433 VTAIL.n375 0.155672
R2461 VTAIL.n426 VTAIL.n375 0.155672
R2462 VTAIL.n426 VTAIL.n425 0.155672
R2463 VTAIL.n425 VTAIL.n379 0.155672
R2464 VTAIL.n418 VTAIL.n379 0.155672
R2465 VTAIL.n418 VTAIL.n417 0.155672
R2466 VTAIL.n417 VTAIL.n383 0.155672
R2467 VTAIL.n410 VTAIL.n383 0.155672
R2468 VTAIL.n410 VTAIL.n409 0.155672
R2469 VTAIL.n409 VTAIL.n389 0.155672
R2470 VTAIL.n402 VTAIL.n389 0.155672
R2471 VTAIL.n402 VTAIL.n401 0.155672
R2472 VTAIL.n401 VTAIL.n393 0.155672
R2473 VTAIL.n367 VTAIL.n297 0.155672
R2474 VTAIL.n360 VTAIL.n297 0.155672
R2475 VTAIL.n360 VTAIL.n359 0.155672
R2476 VTAIL.n359 VTAIL.n301 0.155672
R2477 VTAIL.n352 VTAIL.n301 0.155672
R2478 VTAIL.n352 VTAIL.n351 0.155672
R2479 VTAIL.n351 VTAIL.n305 0.155672
R2480 VTAIL.n344 VTAIL.n305 0.155672
R2481 VTAIL.n344 VTAIL.n343 0.155672
R2482 VTAIL.n343 VTAIL.n309 0.155672
R2483 VTAIL.n336 VTAIL.n309 0.155672
R2484 VTAIL.n336 VTAIL.n335 0.155672
R2485 VTAIL.n335 VTAIL.n315 0.155672
R2486 VTAIL.n328 VTAIL.n315 0.155672
R2487 VTAIL.n328 VTAIL.n327 0.155672
R2488 VTAIL.n327 VTAIL.n319 0.155672
R2489 VTAIL.n293 VTAIL.n223 0.155672
R2490 VTAIL.n286 VTAIL.n223 0.155672
R2491 VTAIL.n286 VTAIL.n285 0.155672
R2492 VTAIL.n285 VTAIL.n227 0.155672
R2493 VTAIL.n278 VTAIL.n227 0.155672
R2494 VTAIL.n278 VTAIL.n277 0.155672
R2495 VTAIL.n277 VTAIL.n231 0.155672
R2496 VTAIL.n270 VTAIL.n231 0.155672
R2497 VTAIL.n270 VTAIL.n269 0.155672
R2498 VTAIL.n269 VTAIL.n235 0.155672
R2499 VTAIL.n262 VTAIL.n235 0.155672
R2500 VTAIL.n262 VTAIL.n261 0.155672
R2501 VTAIL.n261 VTAIL.n241 0.155672
R2502 VTAIL.n254 VTAIL.n241 0.155672
R2503 VTAIL.n254 VTAIL.n253 0.155672
R2504 VTAIL.n253 VTAIL.n245 0.155672
R2505 VP.n19 VP.n18 161.3
R2506 VP.n17 VP.n1 161.3
R2507 VP.n16 VP.n15 161.3
R2508 VP.n14 VP.n2 161.3
R2509 VP.n13 VP.n12 161.3
R2510 VP.n11 VP.n3 161.3
R2511 VP.n10 VP.n9 161.3
R2512 VP.n8 VP.n4 161.3
R2513 VP.n5 VP.t0 129.168
R2514 VP.n5 VP.t2 127.972
R2515 VP.n6 VP.t1 95.2697
R2516 VP.n0 VP.t3 95.2697
R2517 VP.n7 VP.n6 84.0486
R2518 VP.n20 VP.n0 84.0486
R2519 VP.n12 VP.n2 56.4773
R2520 VP.n7 VP.n5 52.179
R2521 VP.n10 VP.n4 24.3439
R2522 VP.n11 VP.n10 24.3439
R2523 VP.n12 VP.n11 24.3439
R2524 VP.n16 VP.n2 24.3439
R2525 VP.n17 VP.n16 24.3439
R2526 VP.n18 VP.n17 24.3439
R2527 VP.n6 VP.n4 5.84292
R2528 VP.n18 VP.n0 5.84292
R2529 VP.n8 VP.n7 0.355081
R2530 VP.n20 VP.n19 0.355081
R2531 VP VP.n20 0.26685
R2532 VP.n9 VP.n8 0.189894
R2533 VP.n9 VP.n3 0.189894
R2534 VP.n13 VP.n3 0.189894
R2535 VP.n14 VP.n13 0.189894
R2536 VP.n15 VP.n14 0.189894
R2537 VP.n15 VP.n1 0.189894
R2538 VP.n19 VP.n1 0.189894
R2539 VDD1 VDD1.n1 105.535
R2540 VDD1 VDD1.n0 60.0607
R2541 VDD1.n0 VDD1.t3 1.46934
R2542 VDD1.n0 VDD1.t1 1.46934
R2543 VDD1.n1 VDD1.t2 1.46934
R2544 VDD1.n1 VDD1.t0 1.46934
C0 VDD1 VP 5.82369f
C1 VDD2 VTAIL 5.98939f
C2 VDD1 VN 0.149547f
C3 VDD2 VP 0.445662f
C4 VDD2 VN 5.52852f
C5 VTAIL VP 5.50725f
C6 VN VTAIL 5.49314f
C7 VDD1 VDD2 1.21812f
C8 VN VP 7.05845f
C9 VDD1 VTAIL 5.92975f
C10 VDD2 B 4.350386f
C11 VDD1 B 8.91256f
C12 VTAIL B 11.420152f
C13 VN B 12.387699f
C14 VP B 10.771137f
C15 VDD1.t3 B 0.289439f
C16 VDD1.t1 B 0.289439f
C17 VDD1.n0 B 2.59443f
C18 VDD1.t2 B 0.289439f
C19 VDD1.t0 B 0.289439f
C20 VDD1.n1 B 3.41773f
C21 VP.t3 B 2.6851f
C22 VP.n0 B 1.01365f
C23 VP.n1 B 0.021372f
C24 VP.n2 B 0.031335f
C25 VP.n3 B 0.021372f
C26 VP.n4 B 0.02501f
C27 VP.t0 B 2.9741f
C28 VP.t2 B 2.96422f
C29 VP.n5 B 3.19674f
C30 VP.t1 B 2.6851f
C31 VP.n6 B 1.01365f
C32 VP.n7 B 1.29931f
C33 VP.n8 B 0.0345f
C34 VP.n9 B 0.021372f
C35 VP.n10 B 0.040032f
C36 VP.n11 B 0.040032f
C37 VP.n12 B 0.031335f
C38 VP.n13 B 0.021372f
C39 VP.n14 B 0.021372f
C40 VP.n15 B 0.021372f
C41 VP.n16 B 0.040032f
C42 VP.n17 B 0.040032f
C43 VP.n18 B 0.02501f
C44 VP.n19 B 0.0345f
C45 VP.n20 B 0.059352f
C46 VTAIL.n0 B 0.023197f
C47 VTAIL.n1 B 0.016503f
C48 VTAIL.n2 B 0.008868f
C49 VTAIL.n3 B 0.020961f
C50 VTAIL.n4 B 0.00939f
C51 VTAIL.n5 B 0.016503f
C52 VTAIL.n6 B 0.008868f
C53 VTAIL.n7 B 0.020961f
C54 VTAIL.n8 B 0.00939f
C55 VTAIL.n9 B 0.016503f
C56 VTAIL.n10 B 0.008868f
C57 VTAIL.n11 B 0.020961f
C58 VTAIL.n12 B 0.009129f
C59 VTAIL.n13 B 0.016503f
C60 VTAIL.n14 B 0.00939f
C61 VTAIL.n15 B 0.020961f
C62 VTAIL.n16 B 0.00939f
C63 VTAIL.n17 B 0.016503f
C64 VTAIL.n18 B 0.008868f
C65 VTAIL.n19 B 0.020961f
C66 VTAIL.n20 B 0.00939f
C67 VTAIL.n21 B 0.941204f
C68 VTAIL.n22 B 0.008868f
C69 VTAIL.t7 B 0.035533f
C70 VTAIL.n23 B 0.128364f
C71 VTAIL.n24 B 0.014818f
C72 VTAIL.n25 B 0.015721f
C73 VTAIL.n26 B 0.020961f
C74 VTAIL.n27 B 0.00939f
C75 VTAIL.n28 B 0.008868f
C76 VTAIL.n29 B 0.016503f
C77 VTAIL.n30 B 0.016503f
C78 VTAIL.n31 B 0.008868f
C79 VTAIL.n32 B 0.00939f
C80 VTAIL.n33 B 0.020961f
C81 VTAIL.n34 B 0.020961f
C82 VTAIL.n35 B 0.00939f
C83 VTAIL.n36 B 0.008868f
C84 VTAIL.n37 B 0.016503f
C85 VTAIL.n38 B 0.016503f
C86 VTAIL.n39 B 0.008868f
C87 VTAIL.n40 B 0.008868f
C88 VTAIL.n41 B 0.00939f
C89 VTAIL.n42 B 0.020961f
C90 VTAIL.n43 B 0.020961f
C91 VTAIL.n44 B 0.020961f
C92 VTAIL.n45 B 0.009129f
C93 VTAIL.n46 B 0.008868f
C94 VTAIL.n47 B 0.016503f
C95 VTAIL.n48 B 0.016503f
C96 VTAIL.n49 B 0.008868f
C97 VTAIL.n50 B 0.00939f
C98 VTAIL.n51 B 0.020961f
C99 VTAIL.n52 B 0.020961f
C100 VTAIL.n53 B 0.00939f
C101 VTAIL.n54 B 0.008868f
C102 VTAIL.n55 B 0.016503f
C103 VTAIL.n56 B 0.016503f
C104 VTAIL.n57 B 0.008868f
C105 VTAIL.n58 B 0.00939f
C106 VTAIL.n59 B 0.020961f
C107 VTAIL.n60 B 0.020961f
C108 VTAIL.n61 B 0.00939f
C109 VTAIL.n62 B 0.008868f
C110 VTAIL.n63 B 0.016503f
C111 VTAIL.n64 B 0.016503f
C112 VTAIL.n65 B 0.008868f
C113 VTAIL.n66 B 0.00939f
C114 VTAIL.n67 B 0.020961f
C115 VTAIL.n68 B 0.045377f
C116 VTAIL.n69 B 0.00939f
C117 VTAIL.n70 B 0.008868f
C118 VTAIL.n71 B 0.036343f
C119 VTAIL.n72 B 0.025334f
C120 VTAIL.n73 B 0.126883f
C121 VTAIL.n74 B 0.023197f
C122 VTAIL.n75 B 0.016503f
C123 VTAIL.n76 B 0.008868f
C124 VTAIL.n77 B 0.020961f
C125 VTAIL.n78 B 0.00939f
C126 VTAIL.n79 B 0.016503f
C127 VTAIL.n80 B 0.008868f
C128 VTAIL.n81 B 0.020961f
C129 VTAIL.n82 B 0.00939f
C130 VTAIL.n83 B 0.016503f
C131 VTAIL.n84 B 0.008868f
C132 VTAIL.n85 B 0.020961f
C133 VTAIL.n86 B 0.009129f
C134 VTAIL.n87 B 0.016503f
C135 VTAIL.n88 B 0.00939f
C136 VTAIL.n89 B 0.020961f
C137 VTAIL.n90 B 0.00939f
C138 VTAIL.n91 B 0.016503f
C139 VTAIL.n92 B 0.008868f
C140 VTAIL.n93 B 0.020961f
C141 VTAIL.n94 B 0.00939f
C142 VTAIL.n95 B 0.941204f
C143 VTAIL.n96 B 0.008868f
C144 VTAIL.t2 B 0.035533f
C145 VTAIL.n97 B 0.128364f
C146 VTAIL.n98 B 0.014818f
C147 VTAIL.n99 B 0.015721f
C148 VTAIL.n100 B 0.020961f
C149 VTAIL.n101 B 0.00939f
C150 VTAIL.n102 B 0.008868f
C151 VTAIL.n103 B 0.016503f
C152 VTAIL.n104 B 0.016503f
C153 VTAIL.n105 B 0.008868f
C154 VTAIL.n106 B 0.00939f
C155 VTAIL.n107 B 0.020961f
C156 VTAIL.n108 B 0.020961f
C157 VTAIL.n109 B 0.00939f
C158 VTAIL.n110 B 0.008868f
C159 VTAIL.n111 B 0.016503f
C160 VTAIL.n112 B 0.016503f
C161 VTAIL.n113 B 0.008868f
C162 VTAIL.n114 B 0.008868f
C163 VTAIL.n115 B 0.00939f
C164 VTAIL.n116 B 0.020961f
C165 VTAIL.n117 B 0.020961f
C166 VTAIL.n118 B 0.020961f
C167 VTAIL.n119 B 0.009129f
C168 VTAIL.n120 B 0.008868f
C169 VTAIL.n121 B 0.016503f
C170 VTAIL.n122 B 0.016503f
C171 VTAIL.n123 B 0.008868f
C172 VTAIL.n124 B 0.00939f
C173 VTAIL.n125 B 0.020961f
C174 VTAIL.n126 B 0.020961f
C175 VTAIL.n127 B 0.00939f
C176 VTAIL.n128 B 0.008868f
C177 VTAIL.n129 B 0.016503f
C178 VTAIL.n130 B 0.016503f
C179 VTAIL.n131 B 0.008868f
C180 VTAIL.n132 B 0.00939f
C181 VTAIL.n133 B 0.020961f
C182 VTAIL.n134 B 0.020961f
C183 VTAIL.n135 B 0.00939f
C184 VTAIL.n136 B 0.008868f
C185 VTAIL.n137 B 0.016503f
C186 VTAIL.n138 B 0.016503f
C187 VTAIL.n139 B 0.008868f
C188 VTAIL.n140 B 0.00939f
C189 VTAIL.n141 B 0.020961f
C190 VTAIL.n142 B 0.045377f
C191 VTAIL.n143 B 0.00939f
C192 VTAIL.n144 B 0.008868f
C193 VTAIL.n145 B 0.036343f
C194 VTAIL.n146 B 0.025334f
C195 VTAIL.n147 B 0.209514f
C196 VTAIL.n148 B 0.023197f
C197 VTAIL.n149 B 0.016503f
C198 VTAIL.n150 B 0.008868f
C199 VTAIL.n151 B 0.020961f
C200 VTAIL.n152 B 0.00939f
C201 VTAIL.n153 B 0.016503f
C202 VTAIL.n154 B 0.008868f
C203 VTAIL.n155 B 0.020961f
C204 VTAIL.n156 B 0.00939f
C205 VTAIL.n157 B 0.016503f
C206 VTAIL.n158 B 0.008868f
C207 VTAIL.n159 B 0.020961f
C208 VTAIL.n160 B 0.009129f
C209 VTAIL.n161 B 0.016503f
C210 VTAIL.n162 B 0.00939f
C211 VTAIL.n163 B 0.020961f
C212 VTAIL.n164 B 0.00939f
C213 VTAIL.n165 B 0.016503f
C214 VTAIL.n166 B 0.008868f
C215 VTAIL.n167 B 0.020961f
C216 VTAIL.n168 B 0.00939f
C217 VTAIL.n169 B 0.941204f
C218 VTAIL.n170 B 0.008868f
C219 VTAIL.t0 B 0.035533f
C220 VTAIL.n171 B 0.128364f
C221 VTAIL.n172 B 0.014818f
C222 VTAIL.n173 B 0.015721f
C223 VTAIL.n174 B 0.020961f
C224 VTAIL.n175 B 0.00939f
C225 VTAIL.n176 B 0.008868f
C226 VTAIL.n177 B 0.016503f
C227 VTAIL.n178 B 0.016503f
C228 VTAIL.n179 B 0.008868f
C229 VTAIL.n180 B 0.00939f
C230 VTAIL.n181 B 0.020961f
C231 VTAIL.n182 B 0.020961f
C232 VTAIL.n183 B 0.00939f
C233 VTAIL.n184 B 0.008868f
C234 VTAIL.n185 B 0.016503f
C235 VTAIL.n186 B 0.016503f
C236 VTAIL.n187 B 0.008868f
C237 VTAIL.n188 B 0.008868f
C238 VTAIL.n189 B 0.00939f
C239 VTAIL.n190 B 0.020961f
C240 VTAIL.n191 B 0.020961f
C241 VTAIL.n192 B 0.020961f
C242 VTAIL.n193 B 0.009129f
C243 VTAIL.n194 B 0.008868f
C244 VTAIL.n195 B 0.016503f
C245 VTAIL.n196 B 0.016503f
C246 VTAIL.n197 B 0.008868f
C247 VTAIL.n198 B 0.00939f
C248 VTAIL.n199 B 0.020961f
C249 VTAIL.n200 B 0.020961f
C250 VTAIL.n201 B 0.00939f
C251 VTAIL.n202 B 0.008868f
C252 VTAIL.n203 B 0.016503f
C253 VTAIL.n204 B 0.016503f
C254 VTAIL.n205 B 0.008868f
C255 VTAIL.n206 B 0.00939f
C256 VTAIL.n207 B 0.020961f
C257 VTAIL.n208 B 0.020961f
C258 VTAIL.n209 B 0.00939f
C259 VTAIL.n210 B 0.008868f
C260 VTAIL.n211 B 0.016503f
C261 VTAIL.n212 B 0.016503f
C262 VTAIL.n213 B 0.008868f
C263 VTAIL.n214 B 0.00939f
C264 VTAIL.n215 B 0.020961f
C265 VTAIL.n216 B 0.045377f
C266 VTAIL.n217 B 0.00939f
C267 VTAIL.n218 B 0.008868f
C268 VTAIL.n219 B 0.036343f
C269 VTAIL.n220 B 0.025334f
C270 VTAIL.n221 B 1.19812f
C271 VTAIL.n222 B 0.023197f
C272 VTAIL.n223 B 0.016503f
C273 VTAIL.n224 B 0.008868f
C274 VTAIL.n225 B 0.020961f
C275 VTAIL.n226 B 0.00939f
C276 VTAIL.n227 B 0.016503f
C277 VTAIL.n228 B 0.008868f
C278 VTAIL.n229 B 0.020961f
C279 VTAIL.n230 B 0.00939f
C280 VTAIL.n231 B 0.016503f
C281 VTAIL.n232 B 0.008868f
C282 VTAIL.n233 B 0.020961f
C283 VTAIL.n234 B 0.009129f
C284 VTAIL.n235 B 0.016503f
C285 VTAIL.n236 B 0.009129f
C286 VTAIL.n237 B 0.008868f
C287 VTAIL.n238 B 0.020961f
C288 VTAIL.n239 B 0.020961f
C289 VTAIL.n240 B 0.00939f
C290 VTAIL.n241 B 0.016503f
C291 VTAIL.n242 B 0.008868f
C292 VTAIL.n243 B 0.020961f
C293 VTAIL.n244 B 0.00939f
C294 VTAIL.n245 B 0.941204f
C295 VTAIL.n246 B 0.008868f
C296 VTAIL.t5 B 0.035533f
C297 VTAIL.n247 B 0.128364f
C298 VTAIL.n248 B 0.014818f
C299 VTAIL.n249 B 0.015721f
C300 VTAIL.n250 B 0.020961f
C301 VTAIL.n251 B 0.00939f
C302 VTAIL.n252 B 0.008868f
C303 VTAIL.n253 B 0.016503f
C304 VTAIL.n254 B 0.016503f
C305 VTAIL.n255 B 0.008868f
C306 VTAIL.n256 B 0.00939f
C307 VTAIL.n257 B 0.020961f
C308 VTAIL.n258 B 0.020961f
C309 VTAIL.n259 B 0.00939f
C310 VTAIL.n260 B 0.008868f
C311 VTAIL.n261 B 0.016503f
C312 VTAIL.n262 B 0.016503f
C313 VTAIL.n263 B 0.008868f
C314 VTAIL.n264 B 0.00939f
C315 VTAIL.n265 B 0.020961f
C316 VTAIL.n266 B 0.020961f
C317 VTAIL.n267 B 0.00939f
C318 VTAIL.n268 B 0.008868f
C319 VTAIL.n269 B 0.016503f
C320 VTAIL.n270 B 0.016503f
C321 VTAIL.n271 B 0.008868f
C322 VTAIL.n272 B 0.00939f
C323 VTAIL.n273 B 0.020961f
C324 VTAIL.n274 B 0.020961f
C325 VTAIL.n275 B 0.00939f
C326 VTAIL.n276 B 0.008868f
C327 VTAIL.n277 B 0.016503f
C328 VTAIL.n278 B 0.016503f
C329 VTAIL.n279 B 0.008868f
C330 VTAIL.n280 B 0.00939f
C331 VTAIL.n281 B 0.020961f
C332 VTAIL.n282 B 0.020961f
C333 VTAIL.n283 B 0.00939f
C334 VTAIL.n284 B 0.008868f
C335 VTAIL.n285 B 0.016503f
C336 VTAIL.n286 B 0.016503f
C337 VTAIL.n287 B 0.008868f
C338 VTAIL.n288 B 0.00939f
C339 VTAIL.n289 B 0.020961f
C340 VTAIL.n290 B 0.045377f
C341 VTAIL.n291 B 0.00939f
C342 VTAIL.n292 B 0.008868f
C343 VTAIL.n293 B 0.036343f
C344 VTAIL.n294 B 0.025334f
C345 VTAIL.n295 B 1.19812f
C346 VTAIL.n296 B 0.023197f
C347 VTAIL.n297 B 0.016503f
C348 VTAIL.n298 B 0.008868f
C349 VTAIL.n299 B 0.020961f
C350 VTAIL.n300 B 0.00939f
C351 VTAIL.n301 B 0.016503f
C352 VTAIL.n302 B 0.008868f
C353 VTAIL.n303 B 0.020961f
C354 VTAIL.n304 B 0.00939f
C355 VTAIL.n305 B 0.016503f
C356 VTAIL.n306 B 0.008868f
C357 VTAIL.n307 B 0.020961f
C358 VTAIL.n308 B 0.009129f
C359 VTAIL.n309 B 0.016503f
C360 VTAIL.n310 B 0.009129f
C361 VTAIL.n311 B 0.008868f
C362 VTAIL.n312 B 0.020961f
C363 VTAIL.n313 B 0.020961f
C364 VTAIL.n314 B 0.00939f
C365 VTAIL.n315 B 0.016503f
C366 VTAIL.n316 B 0.008868f
C367 VTAIL.n317 B 0.020961f
C368 VTAIL.n318 B 0.00939f
C369 VTAIL.n319 B 0.941204f
C370 VTAIL.n320 B 0.008868f
C371 VTAIL.t6 B 0.035533f
C372 VTAIL.n321 B 0.128364f
C373 VTAIL.n322 B 0.014818f
C374 VTAIL.n323 B 0.015721f
C375 VTAIL.n324 B 0.020961f
C376 VTAIL.n325 B 0.00939f
C377 VTAIL.n326 B 0.008868f
C378 VTAIL.n327 B 0.016503f
C379 VTAIL.n328 B 0.016503f
C380 VTAIL.n329 B 0.008868f
C381 VTAIL.n330 B 0.00939f
C382 VTAIL.n331 B 0.020961f
C383 VTAIL.n332 B 0.020961f
C384 VTAIL.n333 B 0.00939f
C385 VTAIL.n334 B 0.008868f
C386 VTAIL.n335 B 0.016503f
C387 VTAIL.n336 B 0.016503f
C388 VTAIL.n337 B 0.008868f
C389 VTAIL.n338 B 0.00939f
C390 VTAIL.n339 B 0.020961f
C391 VTAIL.n340 B 0.020961f
C392 VTAIL.n341 B 0.00939f
C393 VTAIL.n342 B 0.008868f
C394 VTAIL.n343 B 0.016503f
C395 VTAIL.n344 B 0.016503f
C396 VTAIL.n345 B 0.008868f
C397 VTAIL.n346 B 0.00939f
C398 VTAIL.n347 B 0.020961f
C399 VTAIL.n348 B 0.020961f
C400 VTAIL.n349 B 0.00939f
C401 VTAIL.n350 B 0.008868f
C402 VTAIL.n351 B 0.016503f
C403 VTAIL.n352 B 0.016503f
C404 VTAIL.n353 B 0.008868f
C405 VTAIL.n354 B 0.00939f
C406 VTAIL.n355 B 0.020961f
C407 VTAIL.n356 B 0.020961f
C408 VTAIL.n357 B 0.00939f
C409 VTAIL.n358 B 0.008868f
C410 VTAIL.n359 B 0.016503f
C411 VTAIL.n360 B 0.016503f
C412 VTAIL.n361 B 0.008868f
C413 VTAIL.n362 B 0.00939f
C414 VTAIL.n363 B 0.020961f
C415 VTAIL.n364 B 0.045377f
C416 VTAIL.n365 B 0.00939f
C417 VTAIL.n366 B 0.008868f
C418 VTAIL.n367 B 0.036343f
C419 VTAIL.n368 B 0.025334f
C420 VTAIL.n369 B 0.209514f
C421 VTAIL.n370 B 0.023197f
C422 VTAIL.n371 B 0.016503f
C423 VTAIL.n372 B 0.008868f
C424 VTAIL.n373 B 0.020961f
C425 VTAIL.n374 B 0.00939f
C426 VTAIL.n375 B 0.016503f
C427 VTAIL.n376 B 0.008868f
C428 VTAIL.n377 B 0.020961f
C429 VTAIL.n378 B 0.00939f
C430 VTAIL.n379 B 0.016503f
C431 VTAIL.n380 B 0.008868f
C432 VTAIL.n381 B 0.020961f
C433 VTAIL.n382 B 0.009129f
C434 VTAIL.n383 B 0.016503f
C435 VTAIL.n384 B 0.009129f
C436 VTAIL.n385 B 0.008868f
C437 VTAIL.n386 B 0.020961f
C438 VTAIL.n387 B 0.020961f
C439 VTAIL.n388 B 0.00939f
C440 VTAIL.n389 B 0.016503f
C441 VTAIL.n390 B 0.008868f
C442 VTAIL.n391 B 0.020961f
C443 VTAIL.n392 B 0.00939f
C444 VTAIL.n393 B 0.941204f
C445 VTAIL.n394 B 0.008868f
C446 VTAIL.t3 B 0.035533f
C447 VTAIL.n395 B 0.128364f
C448 VTAIL.n396 B 0.014818f
C449 VTAIL.n397 B 0.015721f
C450 VTAIL.n398 B 0.020961f
C451 VTAIL.n399 B 0.00939f
C452 VTAIL.n400 B 0.008868f
C453 VTAIL.n401 B 0.016503f
C454 VTAIL.n402 B 0.016503f
C455 VTAIL.n403 B 0.008868f
C456 VTAIL.n404 B 0.00939f
C457 VTAIL.n405 B 0.020961f
C458 VTAIL.n406 B 0.020961f
C459 VTAIL.n407 B 0.00939f
C460 VTAIL.n408 B 0.008868f
C461 VTAIL.n409 B 0.016503f
C462 VTAIL.n410 B 0.016503f
C463 VTAIL.n411 B 0.008868f
C464 VTAIL.n412 B 0.00939f
C465 VTAIL.n413 B 0.020961f
C466 VTAIL.n414 B 0.020961f
C467 VTAIL.n415 B 0.00939f
C468 VTAIL.n416 B 0.008868f
C469 VTAIL.n417 B 0.016503f
C470 VTAIL.n418 B 0.016503f
C471 VTAIL.n419 B 0.008868f
C472 VTAIL.n420 B 0.00939f
C473 VTAIL.n421 B 0.020961f
C474 VTAIL.n422 B 0.020961f
C475 VTAIL.n423 B 0.00939f
C476 VTAIL.n424 B 0.008868f
C477 VTAIL.n425 B 0.016503f
C478 VTAIL.n426 B 0.016503f
C479 VTAIL.n427 B 0.008868f
C480 VTAIL.n428 B 0.00939f
C481 VTAIL.n429 B 0.020961f
C482 VTAIL.n430 B 0.020961f
C483 VTAIL.n431 B 0.00939f
C484 VTAIL.n432 B 0.008868f
C485 VTAIL.n433 B 0.016503f
C486 VTAIL.n434 B 0.016503f
C487 VTAIL.n435 B 0.008868f
C488 VTAIL.n436 B 0.00939f
C489 VTAIL.n437 B 0.020961f
C490 VTAIL.n438 B 0.045377f
C491 VTAIL.n439 B 0.00939f
C492 VTAIL.n440 B 0.008868f
C493 VTAIL.n441 B 0.036343f
C494 VTAIL.n442 B 0.025334f
C495 VTAIL.n443 B 0.209514f
C496 VTAIL.n444 B 0.023197f
C497 VTAIL.n445 B 0.016503f
C498 VTAIL.n446 B 0.008868f
C499 VTAIL.n447 B 0.020961f
C500 VTAIL.n448 B 0.00939f
C501 VTAIL.n449 B 0.016503f
C502 VTAIL.n450 B 0.008868f
C503 VTAIL.n451 B 0.020961f
C504 VTAIL.n452 B 0.00939f
C505 VTAIL.n453 B 0.016503f
C506 VTAIL.n454 B 0.008868f
C507 VTAIL.n455 B 0.020961f
C508 VTAIL.n456 B 0.009129f
C509 VTAIL.n457 B 0.016503f
C510 VTAIL.n458 B 0.009129f
C511 VTAIL.n459 B 0.008868f
C512 VTAIL.n460 B 0.020961f
C513 VTAIL.n461 B 0.020961f
C514 VTAIL.n462 B 0.00939f
C515 VTAIL.n463 B 0.016503f
C516 VTAIL.n464 B 0.008868f
C517 VTAIL.n465 B 0.020961f
C518 VTAIL.n466 B 0.00939f
C519 VTAIL.n467 B 0.941204f
C520 VTAIL.n468 B 0.008868f
C521 VTAIL.t1 B 0.035533f
C522 VTAIL.n469 B 0.128364f
C523 VTAIL.n470 B 0.014818f
C524 VTAIL.n471 B 0.015721f
C525 VTAIL.n472 B 0.020961f
C526 VTAIL.n473 B 0.00939f
C527 VTAIL.n474 B 0.008868f
C528 VTAIL.n475 B 0.016503f
C529 VTAIL.n476 B 0.016503f
C530 VTAIL.n477 B 0.008868f
C531 VTAIL.n478 B 0.00939f
C532 VTAIL.n479 B 0.020961f
C533 VTAIL.n480 B 0.020961f
C534 VTAIL.n481 B 0.00939f
C535 VTAIL.n482 B 0.008868f
C536 VTAIL.n483 B 0.016503f
C537 VTAIL.n484 B 0.016503f
C538 VTAIL.n485 B 0.008868f
C539 VTAIL.n486 B 0.00939f
C540 VTAIL.n487 B 0.020961f
C541 VTAIL.n488 B 0.020961f
C542 VTAIL.n489 B 0.00939f
C543 VTAIL.n490 B 0.008868f
C544 VTAIL.n491 B 0.016503f
C545 VTAIL.n492 B 0.016503f
C546 VTAIL.n493 B 0.008868f
C547 VTAIL.n494 B 0.00939f
C548 VTAIL.n495 B 0.020961f
C549 VTAIL.n496 B 0.020961f
C550 VTAIL.n497 B 0.00939f
C551 VTAIL.n498 B 0.008868f
C552 VTAIL.n499 B 0.016503f
C553 VTAIL.n500 B 0.016503f
C554 VTAIL.n501 B 0.008868f
C555 VTAIL.n502 B 0.00939f
C556 VTAIL.n503 B 0.020961f
C557 VTAIL.n504 B 0.020961f
C558 VTAIL.n505 B 0.00939f
C559 VTAIL.n506 B 0.008868f
C560 VTAIL.n507 B 0.016503f
C561 VTAIL.n508 B 0.016503f
C562 VTAIL.n509 B 0.008868f
C563 VTAIL.n510 B 0.00939f
C564 VTAIL.n511 B 0.020961f
C565 VTAIL.n512 B 0.045377f
C566 VTAIL.n513 B 0.00939f
C567 VTAIL.n514 B 0.008868f
C568 VTAIL.n515 B 0.036343f
C569 VTAIL.n516 B 0.025334f
C570 VTAIL.n517 B 1.19812f
C571 VTAIL.n518 B 0.023197f
C572 VTAIL.n519 B 0.016503f
C573 VTAIL.n520 B 0.008868f
C574 VTAIL.n521 B 0.020961f
C575 VTAIL.n522 B 0.00939f
C576 VTAIL.n523 B 0.016503f
C577 VTAIL.n524 B 0.008868f
C578 VTAIL.n525 B 0.020961f
C579 VTAIL.n526 B 0.00939f
C580 VTAIL.n527 B 0.016503f
C581 VTAIL.n528 B 0.008868f
C582 VTAIL.n529 B 0.020961f
C583 VTAIL.n530 B 0.009129f
C584 VTAIL.n531 B 0.016503f
C585 VTAIL.n532 B 0.00939f
C586 VTAIL.n533 B 0.020961f
C587 VTAIL.n534 B 0.00939f
C588 VTAIL.n535 B 0.016503f
C589 VTAIL.n536 B 0.008868f
C590 VTAIL.n537 B 0.020961f
C591 VTAIL.n538 B 0.00939f
C592 VTAIL.n539 B 0.941204f
C593 VTAIL.n540 B 0.008868f
C594 VTAIL.t4 B 0.035533f
C595 VTAIL.n541 B 0.128364f
C596 VTAIL.n542 B 0.014818f
C597 VTAIL.n543 B 0.015721f
C598 VTAIL.n544 B 0.020961f
C599 VTAIL.n545 B 0.00939f
C600 VTAIL.n546 B 0.008868f
C601 VTAIL.n547 B 0.016503f
C602 VTAIL.n548 B 0.016503f
C603 VTAIL.n549 B 0.008868f
C604 VTAIL.n550 B 0.00939f
C605 VTAIL.n551 B 0.020961f
C606 VTAIL.n552 B 0.020961f
C607 VTAIL.n553 B 0.00939f
C608 VTAIL.n554 B 0.008868f
C609 VTAIL.n555 B 0.016503f
C610 VTAIL.n556 B 0.016503f
C611 VTAIL.n557 B 0.008868f
C612 VTAIL.n558 B 0.008868f
C613 VTAIL.n559 B 0.00939f
C614 VTAIL.n560 B 0.020961f
C615 VTAIL.n561 B 0.020961f
C616 VTAIL.n562 B 0.020961f
C617 VTAIL.n563 B 0.009129f
C618 VTAIL.n564 B 0.008868f
C619 VTAIL.n565 B 0.016503f
C620 VTAIL.n566 B 0.016503f
C621 VTAIL.n567 B 0.008868f
C622 VTAIL.n568 B 0.00939f
C623 VTAIL.n569 B 0.020961f
C624 VTAIL.n570 B 0.020961f
C625 VTAIL.n571 B 0.00939f
C626 VTAIL.n572 B 0.008868f
C627 VTAIL.n573 B 0.016503f
C628 VTAIL.n574 B 0.016503f
C629 VTAIL.n575 B 0.008868f
C630 VTAIL.n576 B 0.00939f
C631 VTAIL.n577 B 0.020961f
C632 VTAIL.n578 B 0.020961f
C633 VTAIL.n579 B 0.00939f
C634 VTAIL.n580 B 0.008868f
C635 VTAIL.n581 B 0.016503f
C636 VTAIL.n582 B 0.016503f
C637 VTAIL.n583 B 0.008868f
C638 VTAIL.n584 B 0.00939f
C639 VTAIL.n585 B 0.020961f
C640 VTAIL.n586 B 0.045377f
C641 VTAIL.n587 B 0.00939f
C642 VTAIL.n588 B 0.008868f
C643 VTAIL.n589 B 0.036343f
C644 VTAIL.n590 B 0.025334f
C645 VTAIL.n591 B 1.1093f
C646 VDD2.t0 B 0.286952f
C647 VDD2.t3 B 0.286952f
C648 VDD2.n0 B 3.36025f
C649 VDD2.t2 B 0.286952f
C650 VDD2.t1 B 0.286952f
C651 VDD2.n1 B 2.57163f
C652 VDD2.n2 B 4.13465f
C653 VN.t3 B 2.91113f
C654 VN.t0 B 2.92084f
C655 VN.n0 B 1.78753f
C656 VN.t1 B 2.92084f
C657 VN.t2 B 2.91113f
C658 VN.n1 B 3.14792f
.ends

