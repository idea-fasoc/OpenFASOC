* NGSPICE file created from opamp_sample_0003.ext - technology: sky130A

.subckt opamp_sample_0003 GND VOUT VDD VN VP CS_BIAS DIFFPAIR_BIAS
X0 VDD.t157 a_n24758_8502.t18 VOUT.t78 VDD.t138 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X1 GND.t154 GND.t152 VP.t3 GND.t153 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X2 GND.t151 GND.t149 VN.t3 GND.t150 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X3 GND.t231 CS_BIAS.t32 VOUT.t104 GND.t171 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=1.2309 ps=4.39 w=3.73 l=5.83
X4 VDD.t71 VDD.t69 VDD.t70 VDD.t44 sky130_fd_pr__pfet_01v8 ad=2.7576 pd=9.1 as=0 ps=0 w=3.83 l=5.98
X5 VDD.t156 a_n24758_8502.t19 VOUT.t77 VDD.t102 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X6 VOUT.t105 CS_BIAS.t33 GND.t232 GND.t38 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X7 VDD.t155 a_n24758_8502.t20 VOUT.t53 VDD.t110 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X8 GND.t176 CS_BIAS.t34 VOUT.t27 GND.t175 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X9 VOUT.t52 a_n24758_8502.t21 VDD.t154 VDD.t118 sky130_fd_pr__pfet_01v8 ad=2.2104 pd=7.58 as=1.0131 ps=3.73 w=3.07 l=5.49
X10 GND.t148 GND.t145 GND.t147 GND.t146 sky130_fd_pr__nfet_01v8 ad=1.8072 pd=6.46 as=0 ps=0 w=2.51 l=2.32
X11 GND.t177 CS_BIAS.t35 VOUT.t28 GND.t175 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X12 GND.t144 GND.t142 GND.t143 GND.t46 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=0 ps=0 w=3.73 l=5.83
X13 VDD.t68 VDD.t66 VDD.t67 VDD.t63 sky130_fd_pr__pfet_01v8 ad=2.7576 pd=9.1 as=0 ps=0 w=3.83 l=5.98
X14 VOUT.t97 CS_BIAS.t36 GND.t222 GND.t4 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X15 VOUT.t98 CS_BIAS.t37 GND.t223 GND.t4 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X16 a_n24758_8502.t12 a_n11922_9718.t24 a_n6268_8041.t14 VDD.t91 sky130_fd_pr__pfet_01v8 ad=2.7576 pd=9.1 as=1.2639 ps=4.49 w=3.83 l=5.98
X17 VDD.t153 a_n24758_8502.t22 VOUT.t51 VDD.t126 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X18 a_n24758_8502.t10 VN.t4 a_n5140_n467.t24 GND.t199 sky130_fd_pr__nfet_01v8 ad=1.9668 pd=6.62 as=1.9668 ps=6.62 w=5.96 l=3.44
X19 a_n24758_8502.t0 VN.t5 a_n5140_n467.t23 GND.t11 sky130_fd_pr__nfet_01v8 ad=1.9668 pd=6.62 as=1.9668 ps=6.62 w=5.96 l=3.44
X20 VOUT.t50 a_n24758_8502.t23 VDD.t152 VDD.t104 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=2.2104 ps=7.58 w=3.07 l=5.49
X21 VOUT.t100 CS_BIAS.t38 GND.t227 GND.t159 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X22 VDD.t151 a_n24758_8502.t24 VOUT.t86 VDD.t141 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X23 VDD.t150 a_n24758_8502.t25 VOUT.t85 VDD.t110 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X24 GND.t228 CS_BIAS.t39 VOUT.t101 GND.t17 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X25 VOUT.t15 CS_BIAS.t40 GND.t160 GND.t159 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X26 VOUT.t16 CS_BIAS.t41 GND.t161 GND.t22 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=2.6856 ps=8.9 w=3.73 l=5.83
X27 VOUT.t18 CS_BIAS.t42 GND.t163 GND.t22 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=2.6856 ps=8.9 w=3.73 l=5.83
X28 VOUT.t84 a_n24758_8502.t26 VDD.t149 VDD.t118 sky130_fd_pr__pfet_01v8 ad=2.2104 pd=7.58 as=1.0131 ps=3.73 w=3.07 l=5.49
X29 a_n12066_9915.t7 a_n11922_9718.t25 VDD.t83 VDD.t82 sky130_fd_pr__pfet_01v8 ad=1.2639 pd=4.49 as=1.2639 ps=4.49 w=3.83 l=5.98
X30 VDD.t75 a_n11922_9718.t26 a_n6268_8041.t8 VDD.t74 sky130_fd_pr__pfet_01v8 ad=1.2639 pd=4.49 as=1.2639 ps=4.49 w=3.83 l=5.98
X31 VDD.t65 VDD.t62 VDD.t64 VDD.t63 sky130_fd_pr__pfet_01v8 ad=2.7576 pd=9.1 as=0 ps=0 w=3.83 l=5.98
X32 GND.t164 CS_BIAS.t43 VOUT.t19 GND.t17 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X33 VDD.t148 a_n24758_8502.t27 VOUT.t83 VDD.t126 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X34 GND.t141 GND.t139 GND.t140 GND.t130 sky130_fd_pr__nfet_01v8 ad=4.2912 pd=13.36 as=0 ps=0 w=5.96 l=3.44
X35 a_n11922_9718.t13 a_n11922_9718.t12 a_n12066_9915.t13 VDD.t72 sky130_fd_pr__pfet_01v8 ad=1.2639 pd=4.49 as=1.2639 ps=4.49 w=3.83 l=5.98
X36 VOUT.t82 a_n24758_8502.t28 VDD.t147 VDD.t128 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X37 GND.t138 GND.t136 GND.t137 GND.t46 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=0 ps=0 w=3.73 l=5.83
X38 VOUT.t91 CS_BIAS.t44 GND.t215 GND.t25 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X39 VOUT.t92 CS_BIAS.t45 GND.t216 GND.t27 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X40 VOUT.t7 CS_BIAS.t46 GND.t26 GND.t25 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X41 VOUT.t81 a_n24758_8502.t29 VDD.t146 VDD.t107 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X42 VOUT.t80 a_n24758_8502.t30 VDD.t145 VDD.t128 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X43 a_n11922_9718.t10 VP.t4 a_n5140_n467.t11 GND.t11 sky130_fd_pr__nfet_01v8 ad=1.9668 pd=6.62 as=1.9668 ps=6.62 w=5.96 l=3.44
X44 a_n11922_9718.t23 a_n11922_9718.t22 a_n12066_9915.t12 VDD.t2 sky130_fd_pr__pfet_01v8 ad=1.2639 pd=4.49 as=1.2639 ps=4.49 w=3.83 l=5.98
X45 GND.t135 GND.t133 GND.t134 GND.t74 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=0 ps=0 w=3.73 l=5.83
X46 a_n24758_8502.t11 VN.t6 a_n5140_n467.t22 GND.t168 sky130_fd_pr__nfet_01v8 ad=1.9668 pd=6.62 as=4.2912 ps=13.36 w=5.96 l=3.44
X47 VOUT.t8 CS_BIAS.t47 GND.t28 GND.t27 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X48 GND.t42 CS_BIAS.t48 VOUT.t12 GND.t41 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X49 a_n6268_8041.t7 a_n11922_9718.t27 VDD.t95 VDD.t94 sky130_fd_pr__pfet_01v8 ad=2.7576 pd=9.1 as=1.2639 ps=4.49 w=3.83 l=5.98
X50 GND.t43 CS_BIAS.t49 VOUT.t13 GND.t29 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X51 a_n5140_n467.t21 VN.t7 a_n24758_8502.t6 GND.t10 sky130_fd_pr__nfet_01v8 ad=4.2912 pd=13.36 as=1.9668 ps=6.62 w=5.96 l=3.44
X52 GND.t132 GND.t129 GND.t131 GND.t130 sky130_fd_pr__nfet_01v8 ad=4.2912 pd=13.36 as=0 ps=0 w=5.96 l=3.44
X53 GND.t183 CS_BIAS.t50 VOUT.t32 GND.t29 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X54 DIFFPAIR_BIAS.t7 DIFFPAIR_BIAS.t6 GND.t198 GND.t197 sky130_fd_pr__nfet_01v8 ad=1.8072 pd=6.46 as=1.8072 ps=6.46 w=2.51 l=2.32
X55 GND.t224 CS_BIAS.t30 CS_BIAS.t31 GND.t157 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X56 CS_BIAS.t29 CS_BIAS.t28 GND.t194 GND.t22 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=2.6856 ps=8.9 w=3.73 l=5.83
X57 VOUT.t33 CS_BIAS.t51 GND.t184 GND.t20 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=2.6856 ps=8.9 w=3.73 l=5.83
X58 VOUT.t106 a_n6268_8041.t0 sky130_fd_pr__cap_mim_m3_1 l=5.65 w=9.9
X59 VOUT.t25 CS_BIAS.t52 GND.t173 GND.t20 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=2.6856 ps=8.9 w=3.73 l=5.83
X60 VOUT.t79 a_n24758_8502.t31 VDD.t144 VDD.t112 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=2.2104 ps=7.58 w=3.07 l=5.49
X61 CS_BIAS.t27 CS_BIAS.t26 GND.t178 GND.t0 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X62 CS_BIAS.t25 CS_BIAS.t24 GND.t233 GND.t38 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X63 GND.t174 CS_BIAS.t53 VOUT.t26 GND.t41 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X64 GND.t128 GND.t126 GND.t127 GND.t70 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=0 ps=0 w=3.73 l=5.83
X65 a_n11922_9718.t8 VP.t5 a_n5140_n467.t10 GND.t168 sky130_fd_pr__nfet_01v8 ad=1.9668 pd=6.62 as=4.2912 ps=13.36 w=5.96 l=3.44
X66 a_n13678_9915# a_n13678_9915# a_n13678_9915# VDD.t80 sky130_fd_pr__pfet_01v8 ad=2.7576 pd=9.1 as=5.5152 ps=18.2 w=3.83 l=5.98
X67 VOUT.t107 a_n6268_8041.t0 sky130_fd_pr__cap_mim_m3_1 l=5.65 w=9.9
X68 GND.t125 GND.t123 GND.t124 GND.t70 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=0 ps=0 w=3.73 l=5.83
X69 VDD.t163 a_n11922_9718.t28 a_n12066_9915.t6 VDD.t162 sky130_fd_pr__pfet_01v8 ad=1.2639 pd=4.49 as=2.7576 ps=9.1 w=3.83 l=5.98
X70 VDD.t99 a_n11922_9718.t29 a_n12066_9915.t5 VDD.t98 sky130_fd_pr__pfet_01v8 ad=1.2639 pd=4.49 as=1.2639 ps=4.49 w=3.83 l=5.98
X71 VDD.t61 VDD.t59 VDD.t60 VDD.t33 sky130_fd_pr__pfet_01v8 ad=2.2104 pd=7.58 as=0 ps=0 w=3.07 l=5.49
X72 a_n5140_n467.t9 VP.t6 a_n11922_9718.t7 GND.t10 sky130_fd_pr__nfet_01v8 ad=4.2912 pd=13.36 as=1.9668 ps=6.62 w=5.96 l=3.44
X73 VDD.t143 a_n24758_8502.t32 VOUT.t56 VDD.t141 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X74 VDD.t58 VDD.t56 VDD.t57 VDD.t33 sky130_fd_pr__pfet_01v8 ad=2.2104 pd=7.58 as=0 ps=0 w=3.07 l=5.49
X75 VDD.t55 VDD.t53 VDD.t54 VDD.t29 sky130_fd_pr__pfet_01v8 ad=2.2104 pd=7.58 as=0 ps=0 w=3.07 l=5.49
X76 GND.t122 GND.t120 GND.t121 GND.t54 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=0 ps=0 w=3.73 l=5.83
X77 VDD.t86 a_n11922_9718.t30 a_n6268_8041.t6 VDD.t85 sky130_fd_pr__pfet_01v8 ad=1.2639 pd=4.49 as=2.7576 ps=9.1 w=3.83 l=5.98
X78 a_n5140_n467.t8 VP.t7 a_n11922_9718.t5 GND.t15 sky130_fd_pr__nfet_01v8 ad=1.9668 pd=6.62 as=1.9668 ps=6.62 w=5.96 l=3.44
X79 VDD.t142 a_n24758_8502.t33 VOUT.t55 VDD.t141 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X80 GND.t203 CS_BIAS.t54 VOUT.t43 GND.t157 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X81 GND.t204 CS_BIAS.t55 VOUT.t44 GND.t157 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X82 VDD.t52 VDD.t50 VDD.t51 VDD.t29 sky130_fd_pr__pfet_01v8 ad=2.2104 pd=7.58 as=0 ps=0 w=3.07 l=5.49
X83 VDD.t49 VDD.t47 VDD.t48 VDD.t40 sky130_fd_pr__pfet_01v8 ad=2.7576 pd=9.1 as=0 ps=0 w=3.83 l=5.98
X84 GND.t119 GND.t117 GND.t118 GND.t54 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=0 ps=0 w=3.73 l=5.83
X85 GND.t116 GND.t113 GND.t115 GND.t114 sky130_fd_pr__nfet_01v8 ad=1.8072 pd=6.46 as=0 ps=0 w=2.51 l=2.32
X86 VDD.t97 a_n11922_9718.t31 a_n6268_8041.t5 VDD.t96 sky130_fd_pr__pfet_01v8 ad=1.2639 pd=4.49 as=1.2639 ps=4.49 w=3.83 l=5.98
X87 VDD.t140 a_n24758_8502.t34 VOUT.t54 VDD.t138 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X88 a_n12066_9915.t4 a_n11922_9718.t32 VDD.t77 VDD.t76 sky130_fd_pr__pfet_01v8 ad=2.7576 pd=9.1 as=1.2639 ps=4.49 w=3.83 l=5.98
X89 VDD.t161 a_n11922_9718.t33 a_n6268_8041.t4 VDD.t160 sky130_fd_pr__pfet_01v8 ad=1.2639 pd=4.49 as=2.7576 ps=9.1 w=3.83 l=5.98
X90 a_12194_9915# a_12194_9915# a_12194_9915# VDD.t73 sky130_fd_pr__pfet_01v8 ad=2.7576 pd=9.1 as=5.5152 ps=18.2 w=3.83 l=5.98
X91 VN.t2 GND.t110 GND.t112 GND.t111 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X92 VDD.t46 VDD.t43 VDD.t45 VDD.t44 sky130_fd_pr__pfet_01v8 ad=2.7576 pd=9.1 as=0 ps=0 w=3.83 l=5.98
X93 GND.t192 CS_BIAS.t56 VOUT.t38 GND.t191 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X94 VDD.t139 a_n24758_8502.t35 VOUT.t73 VDD.t138 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X95 a_n6268_8041.t3 a_n11922_9718.t34 VDD.t79 VDD.t78 sky130_fd_pr__pfet_01v8 ad=2.7576 pd=9.1 as=1.2639 ps=4.49 w=3.83 l=5.98
X96 VP.t2 GND.t107 GND.t109 GND.t108 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X97 GND.t193 CS_BIAS.t57 VOUT.t39 GND.t157 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X98 GND.t106 GND.t104 GND.t105 GND.t70 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=0 ps=0 w=3.73 l=5.83
X99 VOUT.t5 CS_BIAS.t58 GND.t23 GND.t22 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=2.6856 ps=8.9 w=3.73 l=5.83
X100 a_n5140_n467.t20 VN.t8 a_n24758_8502.t2 GND.t15 sky130_fd_pr__nfet_01v8 ad=1.9668 pd=6.62 as=1.9668 ps=6.62 w=5.96 l=3.44
X101 GND.t225 CS_BIAS.t22 CS_BIAS.t23 GND.t171 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=1.2309 ps=4.39 w=3.73 l=5.83
X102 VOUT.t6 CS_BIAS.t59 GND.t24 GND.t0 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X103 VOUT.t0 CS_BIAS.t60 GND.t1 GND.t0 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X104 GND.t195 CS_BIAS.t20 CS_BIAS.t21 GND.t175 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X105 GND.t3 CS_BIAS.t61 VOUT.t1 GND.t2 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=1.2309 ps=4.39 w=3.73 l=5.83
X106 VOUT.t36 CS_BIAS.t62 GND.t189 GND.t38 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X107 VOUT.t37 CS_BIAS.t63 GND.t190 GND.t0 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X108 GND.t213 CS_BIAS.t64 VOUT.t89 GND.t171 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=1.2309 ps=4.39 w=3.73 l=5.83
X109 DIFFPAIR_BIAS.t5 DIFFPAIR_BIAS.t4 GND.t207 GND.t206 sky130_fd_pr__nfet_01v8 ad=1.8072 pd=6.46 as=1.8072 ps=6.46 w=2.51 l=2.32
X110 GND.t214 CS_BIAS.t65 VOUT.t90 GND.t171 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=1.2309 ps=4.39 w=3.73 l=5.83
X111 VDD.t42 VDD.t39 VDD.t41 VDD.t40 sky130_fd_pr__pfet_01v8 ad=2.7576 pd=9.1 as=0 ps=0 w=3.83 l=5.98
X112 GND.t103 GND.t101 GND.t102 GND.t74 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=0 ps=0 w=3.73 l=5.83
X113 VOUT.t72 a_n24758_8502.t36 VDD.t137 VDD.t114 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X114 VOUT.t10 CS_BIAS.t66 GND.t39 GND.t38 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X115 VOUT.t71 a_n24758_8502.t37 VDD.t136 VDD.t131 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X116 VOUT.t11 CS_BIAS.t67 GND.t40 GND.t38 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X117 DIFFPAIR_BIAS.t3 DIFFPAIR_BIAS.t2 GND.t7 GND.t6 sky130_fd_pr__nfet_01v8 ad=1.8072 pd=6.46 as=1.8072 ps=6.46 w=2.51 l=2.32
X118 CS_BIAS.t19 CS_BIAS.t18 GND.t5 GND.t4 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X119 VDD.t135 a_n24758_8502.t38 VOUT.t49 VDD.t122 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X120 a_n12066_9915.t11 a_n11922_9718.t14 a_n11922_9718.t15 VDD.t91 sky130_fd_pr__pfet_01v8 ad=2.7576 pd=9.1 as=1.2639 ps=4.49 w=3.83 l=5.98
X121 VOUT.t48 a_n24758_8502.t39 VDD.t134 VDD.t131 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X122 GND.t100 GND.t98 GND.t99 GND.t46 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=0 ps=0 w=3.73 l=5.83
X123 VDD.t38 VDD.t36 VDD.t37 VDD.t22 sky130_fd_pr__pfet_01v8 ad=2.2104 pd=7.58 as=0 ps=0 w=3.07 l=5.49
X124 a_n6268_8041.t2 a_n11922_9718.t35 VDD.t90 VDD.t89 sky130_fd_pr__pfet_01v8 ad=1.2639 pd=4.49 as=1.2639 ps=4.49 w=3.83 l=5.98
X125 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.t0 GND.t9 GND.t8 sky130_fd_pr__nfet_01v8 ad=1.8072 pd=6.46 as=1.8072 ps=6.46 w=2.51 l=2.32
X126 GND.t97 GND.t95 GND.t96 GND.t46 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=0 ps=0 w=3.73 l=5.83
X127 VOUT.t47 a_n24758_8502.t40 VDD.t133 VDD.t114 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X128 GND.t94 GND.t92 GND.t93 GND.t54 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=0 ps=0 w=3.73 l=5.83
X129 GND.t181 CS_BIAS.t68 VOUT.t30 GND.t175 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X130 a_n11922_9718.t4 VP.t8 a_n5140_n467.t7 GND.t14 sky130_fd_pr__nfet_01v8 ad=1.9668 pd=6.62 as=1.9668 ps=6.62 w=5.96 l=3.44
X131 VN.t1 GND.t89 GND.t91 GND.t90 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X132 VOUT.t31 CS_BIAS.t69 GND.t182 GND.t4 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X133 a_n24758_8502.t17 a_n11922_9718.t36 a_n6268_8041.t13 VDD.t84 sky130_fd_pr__pfet_01v8 ad=2.7576 pd=9.1 as=1.2639 ps=4.49 w=3.83 l=5.98
X134 a_n5140_n467.t12 DIFFPAIR_BIAS.t8 GND.t13 GND.t12 sky130_fd_pr__nfet_01v8 ad=1.8072 pd=6.46 as=1.8072 ps=6.46 w=2.51 l=2.32
X135 GND.t30 CS_BIAS.t16 CS_BIAS.t17 GND.t29 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X136 VOUT.t46 a_n24758_8502.t41 VDD.t132 VDD.t131 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X137 VP.t1 GND.t86 GND.t88 GND.t87 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X138 VOUT.t65 a_n24758_8502.t42 VDD.t130 VDD.t120 sky130_fd_pr__pfet_01v8 ad=2.2104 pd=7.58 as=1.0131 ps=3.73 w=3.07 l=5.49
X139 VOUT.t41 CS_BIAS.t70 GND.t201 GND.t159 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X140 VOUT.t42 CS_BIAS.t71 GND.t202 GND.t22 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=2.6856 ps=8.9 w=3.73 l=5.83
X141 VOUT.t64 a_n24758_8502.t43 VDD.t129 VDD.t128 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X142 VDD.t127 a_n24758_8502.t44 VOUT.t63 VDD.t126 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X143 VDD.t125 a_n24758_8502.t45 VOUT.t62 VDD.t122 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X144 GND.t220 CS_BIAS.t72 VOUT.t95 GND.t17 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X145 a_n6268_8041.t1 a_n11922_9718.t37 VDD.t101 VDD.t100 sky130_fd_pr__pfet_01v8 ad=1.2639 pd=4.49 as=1.2639 ps=4.49 w=3.83 l=5.98
X146 a_n5140_n467.t19 VN.t9 a_n24758_8502.t16 GND.t32 sky130_fd_pr__nfet_01v8 ad=1.9668 pd=6.62 as=1.9668 ps=6.62 w=5.96 l=3.44
X147 GND.t196 CS_BIAS.t14 CS_BIAS.t15 GND.t191 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X148 VOUT.t96 CS_BIAS.t73 GND.t221 GND.t25 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X149 GND.t205 CS_BIAS.t12 CS_BIAS.t13 GND.t2 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=1.2309 ps=4.39 w=3.73 l=5.83
X150 VOUT.t102 CS_BIAS.t74 GND.t229 GND.t25 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X151 VDD.t93 a_n11922_9718.t38 a_n12066_9915.t3 VDD.t92 sky130_fd_pr__pfet_01v8 ad=1.2639 pd=4.49 as=2.7576 ps=9.1 w=3.83 l=5.98
X152 VOUT.t61 a_n24758_8502.t46 VDD.t124 VDD.t120 sky130_fd_pr__pfet_01v8 ad=2.2104 pd=7.58 as=1.0131 ps=3.73 w=3.07 l=5.49
X153 VDD.t35 VDD.t32 VDD.t34 VDD.t33 sky130_fd_pr__pfet_01v8 ad=2.2104 pd=7.58 as=0 ps=0 w=3.07 l=5.49
X154 VDD.t123 a_n24758_8502.t47 VOUT.t60 VDD.t122 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X155 a_n12066_9915.t10 a_n11922_9718.t16 a_n11922_9718.t17 VDD.t3 sky130_fd_pr__pfet_01v8 ad=1.2639 pd=4.49 as=2.7576 ps=9.1 w=3.83 l=5.98
X156 a_n24758_8502.t1 VN.t10 a_n5140_n467.t18 GND.t14 sky130_fd_pr__nfet_01v8 ad=1.9668 pd=6.62 as=1.9668 ps=6.62 w=5.96 l=3.44
X157 VOUT.t108 a_n6268_8041.t0 sky130_fd_pr__cap_mim_m3_1 l=5.65 w=9.9
X158 CS_BIAS.t11 CS_BIAS.t10 GND.t179 GND.t159 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X159 GND.t85 GND.t83 GND.t84 GND.t70 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=0 ps=0 w=3.73 l=5.83
X160 a_n24758_8502.t4 VN.t11 a_n5140_n467.t17 GND.t155 sky130_fd_pr__nfet_01v8 ad=1.9668 pd=6.62 as=1.9668 ps=6.62 w=5.96 l=3.44
X161 VOUT.t67 a_n24758_8502.t48 VDD.t121 VDD.t120 sky130_fd_pr__pfet_01v8 ad=2.2104 pd=7.58 as=1.0131 ps=3.73 w=3.07 l=5.49
X162 GND.t82 GND.t80 GND.t81 GND.t74 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=0 ps=0 w=3.73 l=5.83
X163 VOUT.t103 CS_BIAS.t75 GND.t230 GND.t27 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X164 GND.t79 GND.t77 GND.t78 GND.t74 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=0 ps=0 w=3.73 l=5.83
X165 VOUT.t66 a_n24758_8502.t49 VDD.t119 VDD.t118 sky130_fd_pr__pfet_01v8 ad=2.2104 pd=7.58 as=1.0131 ps=3.73 w=3.07 l=5.49
X166 VDD.t117 a_n24758_8502.t50 VOUT.t59 VDD.t102 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X167 VOUT.t23 CS_BIAS.t76 GND.t170 GND.t27 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X168 GND.t172 CS_BIAS.t77 VOUT.t24 GND.t171 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=1.2309 ps=4.39 w=3.73 l=5.83
X169 GND.t187 CS_BIAS.t78 VOUT.t34 GND.t175 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X170 a_n5140_n467.t6 VP.t9 a_n11922_9718.t11 GND.t210 sky130_fd_pr__nfet_01v8 ad=4.2912 pd=13.36 as=1.9668 ps=6.62 w=5.96 l=3.44
X171 VDD.t31 VDD.t28 VDD.t30 VDD.t29 sky130_fd_pr__pfet_01v8 ad=2.2104 pd=7.58 as=0 ps=0 w=3.07 l=5.49
X172 VOUT.t109 a_n6268_8041.t0 sky130_fd_pr__cap_mim_m3_1 l=5.65 w=9.9
X173 a_n5140_n467.t5 VP.t10 a_n11922_9718.t9 GND.t32 sky130_fd_pr__nfet_01v8 ad=1.9668 pd=6.62 as=1.9668 ps=6.62 w=5.96 l=3.44
X174 a_n12066_9915.t9 a_n11922_9718.t18 a_n11922_9718.t19 VDD.t84 sky130_fd_pr__pfet_01v8 ad=2.7576 pd=9.1 as=1.2639 ps=4.49 w=3.83 l=5.98
X175 VOUT.t58 a_n24758_8502.t51 VDD.t116 VDD.t112 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=2.2104 ps=7.58 w=3.07 l=5.49
X176 GND.t185 CS_BIAS.t8 CS_BIAS.t9 GND.t17 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X177 GND.t188 CS_BIAS.t79 VOUT.t35 GND.t29 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X178 GND.t76 GND.t73 GND.t75 GND.t74 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=0 ps=0 w=3.73 l=5.83
X179 a_n6268_8041.t12 a_n11922_9718.t39 a_n24758_8502.t13 VDD.t2 sky130_fd_pr__pfet_01v8 ad=1.2639 pd=4.49 as=1.2639 ps=4.49 w=3.83 l=5.98
X180 VOUT.t57 a_n24758_8502.t52 VDD.t115 VDD.t114 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X181 a_n24758_8502.t9 a_n11922_9718.t40 a_n6268_8041.t11 VDD.t81 sky130_fd_pr__pfet_01v8 ad=1.2639 pd=4.49 as=2.7576 ps=9.1 w=3.83 l=5.98
X182 VDD.t27 VDD.t25 VDD.t26 VDD.t22 sky130_fd_pr__pfet_01v8 ad=2.2104 pd=7.58 as=0 ps=0 w=3.07 l=5.49
X183 VOUT.t3 CS_BIAS.t80 GND.t19 GND.t4 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X184 VOUT.t76 a_n24758_8502.t53 VDD.t113 VDD.t112 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=2.2104 ps=7.58 w=3.07 l=5.49
X185 VOUT.t4 CS_BIAS.t81 GND.t21 GND.t20 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=2.6856 ps=8.9 w=3.73 l=5.83
X186 a_n12066_9915.t2 a_n11922_9718.t41 VDD.t88 VDD.t87 sky130_fd_pr__pfet_01v8 ad=1.2639 pd=4.49 as=1.2639 ps=4.49 w=3.83 l=5.98
X187 CS_BIAS.t7 CS_BIAS.t6 GND.t44 GND.t20 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=2.6856 ps=8.9 w=3.73 l=5.83
X188 a_n5140_n467.t4 VP.t11 a_n11922_9718.t3 GND.t186 sky130_fd_pr__nfet_01v8 ad=1.9668 pd=6.62 as=1.9668 ps=6.62 w=5.96 l=3.44
X189 a_n11922_9718.t0 VP.t12 a_n5140_n467.t3 GND.t155 sky130_fd_pr__nfet_01v8 ad=1.9668 pd=6.62 as=1.9668 ps=6.62 w=5.96 l=3.44
X190 GND.t166 CS_BIAS.t82 VOUT.t20 GND.t41 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X191 a_n5140_n467.t27 DIFFPAIR_BIAS.t9 GND.t209 GND.t208 sky130_fd_pr__nfet_01v8 ad=1.8072 pd=6.46 as=1.8072 ps=6.46 w=2.51 l=2.32
X192 GND.t167 CS_BIAS.t83 VOUT.t21 GND.t41 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X193 VDD.t24 VDD.t21 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8 ad=2.2104 pd=7.58 as=0 ps=0 w=3.07 l=5.49
X194 VDD.t20 VDD.t18 VDD.t19 VDD.t9 sky130_fd_pr__pfet_01v8 ad=2.2104 pd=7.58 as=0 ps=0 w=3.07 l=5.49
X195 GND.t218 CS_BIAS.t84 VOUT.t93 GND.t29 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X196 GND.t72 GND.t69 GND.t71 GND.t70 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=0 ps=0 w=3.73 l=5.83
X197 GND.t68 GND.t66 GND.t67 GND.t50 sky130_fd_pr__nfet_01v8 ad=4.2912 pd=13.36 as=0 ps=0 w=5.96 l=3.44
X198 VDD.t17 VDD.t15 VDD.t16 VDD.t5 sky130_fd_pr__pfet_01v8 ad=2.7576 pd=9.1 as=0 ps=0 w=3.83 l=5.98
X199 GND.t65 GND.t63 VN.t0 GND.t64 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X200 a_n5140_n467.t16 VN.t12 a_n24758_8502.t15 GND.t210 sky130_fd_pr__nfet_01v8 ad=4.2912 pd=13.36 as=1.9668 ps=6.62 w=5.96 l=3.44
X201 VDD.t111 a_n24758_8502.t54 VOUT.t75 VDD.t110 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X202 a_n11922_9718.t6 VP.t13 a_n5140_n467.t2 GND.t156 sky130_fd_pr__nfet_01v8 ad=1.9668 pd=6.62 as=4.2912 ps=13.36 w=5.96 l=3.44
X203 GND.t219 CS_BIAS.t85 VOUT.t94 GND.t2 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=1.2309 ps=4.39 w=3.73 l=5.83
X204 a_n5140_n467.t26 DIFFPAIR_BIAS.t10 GND.t36 GND.t35 sky130_fd_pr__nfet_01v8 ad=1.8072 pd=6.46 as=1.8072 ps=6.46 w=2.51 l=2.32
X205 GND.t226 CS_BIAS.t86 VOUT.t99 GND.t191 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X206 a_n24758_8502.t14 a_n11922_9718.t42 a_n6268_8041.t10 VDD.t3 sky130_fd_pr__pfet_01v8 ad=1.2639 pd=4.49 as=2.7576 ps=9.1 w=3.83 l=5.98
X207 VOUT.t74 a_n24758_8502.t55 VDD.t109 VDD.t107 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X208 a_n12066_9915.t1 a_n11922_9718.t43 VDD.t159 VDD.t158 sky130_fd_pr__pfet_01v8 ad=2.7576 pd=9.1 as=1.2639 ps=4.49 w=3.83 l=5.98
X209 a_n5140_n467.t25 DIFFPAIR_BIAS.t11 GND.t34 GND.t33 sky130_fd_pr__nfet_01v8 ad=1.8072 pd=6.46 as=1.8072 ps=6.46 w=2.51 l=2.32
X210 a_n6268_8041.t9 a_n11922_9718.t44 a_n24758_8502.t7 VDD.t72 sky130_fd_pr__pfet_01v8 ad=1.2639 pd=4.49 as=1.2639 ps=4.49 w=3.83 l=5.98
X211 a_n5140_n467.t15 VN.t13 a_n24758_8502.t8 GND.t186 sky130_fd_pr__nfet_01v8 ad=1.9668 pd=6.62 as=1.9668 ps=6.62 w=5.96 l=3.44
X212 a_n5140_n467.t14 VN.t14 a_n24758_8502.t3 GND.t16 sky130_fd_pr__nfet_01v8 ad=1.9668 pd=6.62 as=1.9668 ps=6.62 w=5.96 l=3.44
X213 GND.t62 GND.t60 GND.t61 GND.t54 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=0 ps=0 w=3.73 l=5.83
X214 GND.t158 CS_BIAS.t87 VOUT.t14 GND.t157 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X215 GND.t59 GND.t57 VP.t0 GND.t58 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X216 GND.t56 GND.t53 GND.t55 GND.t54 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=0 ps=0 w=3.73 l=5.83
X217 VOUT.t17 CS_BIAS.t88 GND.t162 GND.t159 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X218 VOUT.t70 a_n24758_8502.t56 VDD.t108 VDD.t107 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X219 VDD.t14 VDD.t12 VDD.t13 VDD.t9 sky130_fd_pr__pfet_01v8 ad=2.2104 pd=7.58 as=0 ps=0 w=3.07 l=5.49
X220 GND.t52 GND.t49 GND.t51 GND.t50 sky130_fd_pr__nfet_01v8 ad=4.2912 pd=13.36 as=0 ps=0 w=5.96 l=3.44
X221 a_n12066_9915.t8 a_n11922_9718.t20 a_n11922_9718.t21 VDD.t81 sky130_fd_pr__pfet_01v8 ad=1.2639 pd=4.49 as=2.7576 ps=9.1 w=3.83 l=5.98
X222 GND.t48 GND.t45 GND.t47 GND.t46 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=0 ps=0 w=3.73 l=5.83
X223 a_n24758_8502.t5 VN.t15 a_n5140_n467.t13 GND.t156 sky130_fd_pr__nfet_01v8 ad=1.9668 pd=6.62 as=4.2912 ps=13.36 w=5.96 l=3.44
X224 CS_BIAS.t5 CS_BIAS.t4 GND.t31 GND.t25 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X225 CS_BIAS.t3 CS_BIAS.t2 GND.t217 GND.t27 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X226 VOUT.t69 a_n24758_8502.t57 VDD.t106 VDD.t104 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=2.2104 ps=7.58 w=3.07 l=5.49
X227 GND.t212 CS_BIAS.t89 VOUT.t88 GND.t191 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X228 GND.t211 CS_BIAS.t90 VOUT.t87 GND.t191 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X229 VDD.t11 VDD.t8 VDD.t10 VDD.t9 sky130_fd_pr__pfet_01v8 ad=2.2104 pd=7.58 as=0 ps=0 w=3.07 l=5.49
X230 GND.t18 CS_BIAS.t91 VOUT.t2 GND.t17 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X231 VDD.t7 VDD.t4 VDD.t6 VDD.t5 sky130_fd_pr__pfet_01v8 ad=2.7576 pd=9.1 as=0 ps=0 w=3.83 l=5.98
X232 VOUT.t68 a_n24758_8502.t58 VDD.t105 VDD.t104 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=2.2104 ps=7.58 w=3.07 l=5.49
X233 GND.t165 CS_BIAS.t0 CS_BIAS.t1 GND.t41 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X234 a_n11922_9718.t1 VP.t14 a_n5140_n467.t1 GND.t199 sky130_fd_pr__nfet_01v8 ad=1.9668 pd=6.62 as=1.9668 ps=6.62 w=5.96 l=3.44
X235 a_n5140_n467.t0 VP.t15 a_n11922_9718.t2 GND.t16 sky130_fd_pr__nfet_01v8 ad=1.9668 pd=6.62 as=1.9668 ps=6.62 w=5.96 l=3.44
X236 VOUT.t9 CS_BIAS.t92 GND.t37 GND.t0 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=1.2309 ps=4.39 w=3.73 l=5.83
X237 GND.t180 CS_BIAS.t93 VOUT.t29 GND.t2 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=1.2309 ps=4.39 w=3.73 l=5.83
X238 VOUT.t22 CS_BIAS.t94 GND.t169 GND.t20 sky130_fd_pr__nfet_01v8 ad=1.2309 pd=4.39 as=2.6856 ps=8.9 w=3.73 l=5.83
X239 VDD.t1 a_n11922_9718.t45 a_n12066_9915.t0 VDD.t0 sky130_fd_pr__pfet_01v8 ad=1.2639 pd=4.49 as=1.2639 ps=4.49 w=3.83 l=5.98
X240 VDD.t103 a_n24758_8502.t59 VOUT.t45 VDD.t102 sky130_fd_pr__pfet_01v8 ad=1.0131 pd=3.73 as=1.0131 ps=3.73 w=3.07 l=5.49
X241 GND.t200 CS_BIAS.t95 VOUT.t40 GND.t2 sky130_fd_pr__nfet_01v8 ad=2.6856 pd=8.9 as=1.2309 ps=4.39 w=3.73 l=5.83
R0 a_n24758_8502.n27 a_n24758_8502.t12 128.156
R1 a_n24758_8502.n25 a_n24758_8502.t17 126.249
R2 a_n24758_8502.n25 a_n24758_8502.n24 111.183
R3 a_n24758_8502.n27 a_n24758_8502.n26 109.275
R4 a_n24758_8502.n23 a_n24758_8502.n31 63.7938
R5 a_n24758_8502.n36 a_n24758_8502.n35 63.7936
R6 a_n24758_8502.n36 a_n24758_8502.n34 63.7936
R7 a_n24758_8502.n37 a_n24758_8502.n36 62.6158
R8 a_n24758_8502.n23 a_n24758_8502.n33 62.6156
R9 a_n24758_8502.n23 a_n24758_8502.n32 62.6156
R10 a_n24758_8502.n10 a_n24758_8502.t42 47.1791
R11 a_n24758_8502.n8 a_n24758_8502.t46 47.1791
R12 a_n24758_8502.n6 a_n24758_8502.t48 47.1791
R13 a_n24758_8502.n0 a_n24758_8502.t57 47.179
R14 a_n24758_8502.n2 a_n24758_8502.t58 47.179
R15 a_n24758_8502.n4 a_n24758_8502.t23 47.179
R16 a_n24758_8502.n28 a_n24758_8502.n25 36.8503
R17 a_n24758_8502.n36 a_n24758_8502.n23 35.5519
R18 a_n24758_8502.n28 a_n24758_8502.n27 26.581
R19 a_n24758_8502.n12 a_n24758_8502.n0 2.10367
R20 a_n24758_8502.n0 a_n24758_8502.n13 0.803298
R21 a_n24758_8502.n0 a_n24758_8502.n1 2.02685
R22 a_n24758_8502.n14 a_n24758_8502.n2 2.10367
R23 a_n24758_8502.n2 a_n24758_8502.n15 0.803298
R24 a_n24758_8502.n2 a_n24758_8502.n3 2.02685
R25 a_n24758_8502.n16 a_n24758_8502.n4 2.10367
R26 a_n24758_8502.n4 a_n24758_8502.n17 0.803298
R27 a_n24758_8502.n4 a_n24758_8502.n5 2.02685
R28 a_n24758_8502.n10 a_n24758_8502.n11 2.89029
R29 a_n24758_8502.n8 a_n24758_8502.n9 2.89029
R30 a_n24758_8502.n6 a_n24758_8502.n7 2.89029
R31 a_n24758_8502.n26 a_n24758_8502.t7 16.9744
R32 a_n24758_8502.n26 a_n24758_8502.t9 16.9744
R33 a_n24758_8502.n24 a_n24758_8502.t13 16.9744
R34 a_n24758_8502.n24 a_n24758_8502.t14 16.9744
R35 a_n24758_8502.n12 a_n24758_8502.t21 48.3076
R36 a_n24758_8502.n12 a_n24758_8502.t32 43.6901
R37 a_n24758_8502.n13 a_n24758_8502.t55 44.8511
R38 a_n24758_8502.n13 a_n24758_8502.t45 45.3701
R39 a_n24758_8502.n1 a_n24758_8502.t28 43.7845
R40 a_n24758_8502.n1 a_n24758_8502.t34 47.7133
R41 a_n24758_8502.n14 a_n24758_8502.t26 48.3076
R42 a_n24758_8502.n14 a_n24758_8502.t33 43.6901
R43 a_n24758_8502.n15 a_n24758_8502.t56 44.8511
R44 a_n24758_8502.n15 a_n24758_8502.t47 45.3701
R45 a_n24758_8502.n3 a_n24758_8502.t30 43.7845
R46 a_n24758_8502.n3 a_n24758_8502.t35 47.7133
R47 a_n24758_8502.n16 a_n24758_8502.t49 48.3076
R48 a_n24758_8502.n16 a_n24758_8502.t24 43.6901
R49 a_n24758_8502.n17 a_n24758_8502.t29 44.8511
R50 a_n24758_8502.n17 a_n24758_8502.t38 45.3701
R51 a_n24758_8502.n5 a_n24758_8502.t43 43.7845
R52 a_n24758_8502.n5 a_n24758_8502.t18 47.7133
R53 a_n24758_8502.n10 a_n24758_8502.t22 44.5164
R54 a_n24758_8502.n18 a_n24758_8502.t39 44.9233
R55 a_n24758_8502.n18 a_n24758_8502.t20 45.3689
R56 a_n24758_8502.n11 a_n24758_8502.t36 46.3106
R57 a_n24758_8502.n11 a_n24758_8502.t59 44.1175
R58 a_n24758_8502.n10 a_n24758_8502.t51 45.693
R59 a_n24758_8502.n8 a_n24758_8502.t27 44.5164
R60 a_n24758_8502.n19 a_n24758_8502.t41 44.9233
R61 a_n24758_8502.n19 a_n24758_8502.t25 45.3689
R62 a_n24758_8502.n9 a_n24758_8502.t40 46.3106
R63 a_n24758_8502.n9 a_n24758_8502.t19 44.1175
R64 a_n24758_8502.n8 a_n24758_8502.t53 45.693
R65 a_n24758_8502.n6 a_n24758_8502.t44 44.5164
R66 a_n24758_8502.n20 a_n24758_8502.t37 44.9233
R67 a_n24758_8502.n20 a_n24758_8502.t54 45.3689
R68 a_n24758_8502.n7 a_n24758_8502.t52 46.3106
R69 a_n24758_8502.n7 a_n24758_8502.t50 44.1175
R70 a_n24758_8502.n6 a_n24758_8502.t31 45.693
R71 a_n24758_8502.n30 a_n24758_8502.n28 11.4887
R72 a_n24758_8502.n29 a_n24758_8502.n22 8.91572
R73 a_n24758_8502.n29 a_n24758_8502.n21 8.10043
R74 a_n24758_8502.n21 a_n24758_8502.n4 7.86675
R75 a_n24758_8502.n22 a_n24758_8502.n6 7.86675
R76 a_n24758_8502.n33 a_n24758_8502.t2 6.6448
R77 a_n24758_8502.n33 a_n24758_8502.t5 6.6448
R78 a_n24758_8502.n32 a_n24758_8502.t8 6.6448
R79 a_n24758_8502.n32 a_n24758_8502.t1 6.6448
R80 a_n24758_8502.n31 a_n24758_8502.t15 6.6448
R81 a_n24758_8502.n31 a_n24758_8502.t10 6.6448
R82 a_n24758_8502.n35 a_n24758_8502.t16 6.6448
R83 a_n24758_8502.n35 a_n24758_8502.t11 6.6448
R84 a_n24758_8502.n34 a_n24758_8502.t6 6.6448
R85 a_n24758_8502.n34 a_n24758_8502.t4 6.6448
R86 a_n24758_8502.n37 a_n24758_8502.t3 6.6448
R87 a_n24758_8502.t0 a_n24758_8502.n37 6.6448
R88 a_n24758_8502.n21 a_n24758_8502.n2 5.44251
R89 a_n24758_8502.n22 a_n24758_8502.n8 5.44251
R90 a_n24758_8502.n30 a_n24758_8502.n29 3.4105
R91 a_n24758_8502.n23 a_n24758_8502.n30 13.5206
R92 a_n24758_8502.n22 a_n24758_8502.n10 7.86675
R93 a_n24758_8502.n21 a_n24758_8502.n0 7.86675
R94 a_n24758_8502.n18 a_n24758_8502.n10 5.39696
R95 a_n24758_8502.n19 a_n24758_8502.n8 5.39696
R96 a_n24758_8502.n20 a_n24758_8502.n6 5.39696
R97 VOUT.n41 VOUT.t66 146.114
R98 VOUT.n34 VOUT.t84 146.114
R99 VOUT.n28 VOUT.t52 146.114
R100 VOUT.n18 VOUT.t67 144.347
R101 VOUT.n11 VOUT.t61 144.347
R102 VOUT.n5 VOUT.t65 144.347
R103 VOUT.n15 VOUT.n13 124.939
R104 VOUT.n8 VOUT.n6 124.939
R105 VOUT.n2 VOUT.n0 124.939
R106 VOUT.n43 VOUT.n42 123.171
R107 VOUT.n41 VOUT.n40 123.171
R108 VOUT.n38 VOUT.n37 123.171
R109 VOUT.n36 VOUT.n35 123.171
R110 VOUT.n34 VOUT.n33 123.171
R111 VOUT.n32 VOUT.n31 123.171
R112 VOUT.n30 VOUT.n29 123.171
R113 VOUT.n28 VOUT.n27 123.171
R114 VOUT.n15 VOUT.n14 123.171
R115 VOUT.n17 VOUT.n16 123.171
R116 VOUT.n8 VOUT.n7 123.171
R117 VOUT.n10 VOUT.n9 123.171
R118 VOUT.n2 VOUT.n1 123.171
R119 VOUT.n4 VOUT.n3 123.171
R120 VOUT.n45 VOUT.n44 123.171
R121 VOUT.n73 VOUT.n71 72.7259
R122 VOUT.n65 VOUT.n63 72.7259
R123 VOUT.n57 VOUT.n55 72.7259
R124 VOUT.n50 VOUT.n48 72.7259
R125 VOUT.n105 VOUT.n103 72.7259
R126 VOUT.n97 VOUT.n95 72.7259
R127 VOUT.n89 VOUT.n87 72.7259
R128 VOUT.n82 VOUT.n80 72.7259
R129 VOUT.n77 VOUT.n76 70.8609
R130 VOUT.n75 VOUT.n74 70.8609
R131 VOUT.n73 VOUT.n72 70.8609
R132 VOUT.n69 VOUT.n68 70.8609
R133 VOUT.n67 VOUT.n66 70.8609
R134 VOUT.n65 VOUT.n64 70.8609
R135 VOUT.n61 VOUT.n60 70.8609
R136 VOUT.n59 VOUT.n58 70.8609
R137 VOUT.n57 VOUT.n56 70.8609
R138 VOUT.n54 VOUT.n53 70.8609
R139 VOUT.n52 VOUT.n51 70.8609
R140 VOUT.n50 VOUT.n49 70.8609
R141 VOUT.n105 VOUT.n104 70.8609
R142 VOUT.n107 VOUT.n106 70.8609
R143 VOUT.n109 VOUT.n108 70.8609
R144 VOUT.n97 VOUT.n96 70.8609
R145 VOUT.n99 VOUT.n98 70.8609
R146 VOUT.n101 VOUT.n100 70.8609
R147 VOUT.n89 VOUT.n88 70.8609
R148 VOUT.n91 VOUT.n90 70.8609
R149 VOUT.n93 VOUT.n92 70.8609
R150 VOUT.n82 VOUT.n81 70.8609
R151 VOUT.n84 VOUT.n83 70.8609
R152 VOUT.n86 VOUT.n85 70.8609
R153 VOUT.n44 VOUT.t78 21.1764
R154 VOUT.n44 VOUT.t50 21.1764
R155 VOUT.n42 VOUT.t49 21.1764
R156 VOUT.n42 VOUT.t64 21.1764
R157 VOUT.n40 VOUT.t86 21.1764
R158 VOUT.n40 VOUT.t81 21.1764
R159 VOUT.n37 VOUT.t73 21.1764
R160 VOUT.n37 VOUT.t68 21.1764
R161 VOUT.n35 VOUT.t60 21.1764
R162 VOUT.n35 VOUT.t80 21.1764
R163 VOUT.n33 VOUT.t55 21.1764
R164 VOUT.n33 VOUT.t70 21.1764
R165 VOUT.n31 VOUT.t54 21.1764
R166 VOUT.n31 VOUT.t69 21.1764
R167 VOUT.n29 VOUT.t62 21.1764
R168 VOUT.n29 VOUT.t82 21.1764
R169 VOUT.n27 VOUT.t56 21.1764
R170 VOUT.n27 VOUT.t74 21.1764
R171 VOUT.n13 VOUT.t59 21.1764
R172 VOUT.n13 VOUT.t79 21.1764
R173 VOUT.n14 VOUT.t75 21.1764
R174 VOUT.n14 VOUT.t57 21.1764
R175 VOUT.n16 VOUT.t63 21.1764
R176 VOUT.n16 VOUT.t71 21.1764
R177 VOUT.n6 VOUT.t77 21.1764
R178 VOUT.n6 VOUT.t76 21.1764
R179 VOUT.n7 VOUT.t85 21.1764
R180 VOUT.n7 VOUT.t47 21.1764
R181 VOUT.n9 VOUT.t83 21.1764
R182 VOUT.n9 VOUT.t46 21.1764
R183 VOUT.n0 VOUT.t45 21.1764
R184 VOUT.n0 VOUT.t58 21.1764
R185 VOUT.n1 VOUT.t53 21.1764
R186 VOUT.n1 VOUT.t72 21.1764
R187 VOUT.n3 VOUT.t51 21.1764
R188 VOUT.n3 VOUT.t48 21.1764
R189 VOUT.n76 VOUT.t13 10.6171
R190 VOUT.n76 VOUT.t33 10.6171
R191 VOUT.n74 VOUT.t101 10.6171
R192 VOUT.n74 VOUT.t10 10.6171
R193 VOUT.n72 VOUT.t43 10.6171
R194 VOUT.n72 VOUT.t97 10.6171
R195 VOUT.n71 VOUT.t29 10.6171
R196 VOUT.n71 VOUT.t103 10.6171
R197 VOUT.n68 VOUT.t35 10.6171
R198 VOUT.n68 VOUT.t4 10.6171
R199 VOUT.n66 VOUT.t95 10.6171
R200 VOUT.n66 VOUT.t105 10.6171
R201 VOUT.n64 VOUT.t14 10.6171
R202 VOUT.n64 VOUT.t31 10.6171
R203 VOUT.n63 VOUT.t1 10.6171
R204 VOUT.n63 VOUT.t8 10.6171
R205 VOUT.n60 VOUT.t32 10.6171
R206 VOUT.n60 VOUT.t25 10.6171
R207 VOUT.n58 VOUT.t19 10.6171
R208 VOUT.n58 VOUT.t11 10.6171
R209 VOUT.n56 VOUT.t44 10.6171
R210 VOUT.n56 VOUT.t98 10.6171
R211 VOUT.n55 VOUT.t40 10.6171
R212 VOUT.n55 VOUT.t23 10.6171
R213 VOUT.n53 VOUT.t93 10.6171
R214 VOUT.n53 VOUT.t22 10.6171
R215 VOUT.n51 VOUT.t2 10.6171
R216 VOUT.n51 VOUT.t36 10.6171
R217 VOUT.n49 VOUT.t39 10.6171
R218 VOUT.n49 VOUT.t3 10.6171
R219 VOUT.n48 VOUT.t94 10.6171
R220 VOUT.n48 VOUT.t92 10.6171
R221 VOUT.n103 VOUT.t87 10.6171
R222 VOUT.n103 VOUT.t18 10.6171
R223 VOUT.n104 VOUT.t27 10.6171
R224 VOUT.n104 VOUT.t96 10.6171
R225 VOUT.n106 VOUT.t20 10.6171
R226 VOUT.n106 VOUT.t100 10.6171
R227 VOUT.n108 VOUT.t89 10.6171
R228 VOUT.n108 VOUT.t6 10.6171
R229 VOUT.n95 VOUT.t38 10.6171
R230 VOUT.n95 VOUT.t42 10.6171
R231 VOUT.n96 VOUT.t30 10.6171
R232 VOUT.n96 VOUT.t91 10.6171
R233 VOUT.n98 VOUT.t26 10.6171
R234 VOUT.n98 VOUT.t41 10.6171
R235 VOUT.n100 VOUT.t104 10.6171
R236 VOUT.n100 VOUT.t9 10.6171
R237 VOUT.n87 VOUT.t88 10.6171
R238 VOUT.n87 VOUT.t16 10.6171
R239 VOUT.n88 VOUT.t28 10.6171
R240 VOUT.n88 VOUT.t102 10.6171
R241 VOUT.n90 VOUT.t21 10.6171
R242 VOUT.n90 VOUT.t15 10.6171
R243 VOUT.n92 VOUT.t90 10.6171
R244 VOUT.n92 VOUT.t0 10.6171
R245 VOUT.n80 VOUT.t99 10.6171
R246 VOUT.n80 VOUT.t5 10.6171
R247 VOUT.n81 VOUT.t34 10.6171
R248 VOUT.n81 VOUT.t7 10.6171
R249 VOUT.n83 VOUT.t12 10.6171
R250 VOUT.n83 VOUT.t17 10.6171
R251 VOUT.n85 VOUT.t24 10.6171
R252 VOUT.n85 VOUT.t37 10.6171
R253 VOUT.n79 VOUT.n47 9.4664
R254 VOUT.n47 VOUT.n20 7.93379
R255 VOUT.n62 VOUT.n54 6.77205
R256 VOUT.n94 VOUT.n86 6.77205
R257 VOUT.n39 VOUT.n32 6.62837
R258 VOUT.n111 VOUT.n79 6.14528
R259 VOUT.n12 VOUT.n5 5.74475
R260 VOUT.n78 VOUT.n77 5.74332
R261 VOUT.n70 VOUT.n69 5.74332
R262 VOUT.n62 VOUT.n61 5.74332
R263 VOUT.n110 VOUT.n109 5.74332
R264 VOUT.n102 VOUT.n101 5.74332
R265 VOUT.n94 VOUT.n93 5.74332
R266 VOUT.n46 VOUT.n45 5.69447
R267 VOUT.n39 VOUT.n38 5.69447
R268 VOUT.n47 VOUT.n46 4.93062
R269 VOUT.n20 VOUT.n19 4.93062
R270 VOUT.n19 VOUT.n18 4.81084
R271 VOUT.n12 VOUT.n11 4.81084
R272 VOUT.n112 VOUT.n20 4.80691
R273 VOUT.n112 VOUT.n111 4.64049
R274 VOUT.n79 VOUT.n78 4.48234
R275 VOUT.n111 VOUT.n110 4.48234
R276 VOUT.n26 VOUT 3.46675
R277 VOUT.n75 VOUT.n73 1.86544
R278 VOUT.n77 VOUT.n75 1.86544
R279 VOUT.n67 VOUT.n65 1.86544
R280 VOUT.n69 VOUT.n67 1.86544
R281 VOUT.n59 VOUT.n57 1.86544
R282 VOUT.n61 VOUT.n59 1.86544
R283 VOUT.n52 VOUT.n50 1.86544
R284 VOUT.n54 VOUT.n52 1.86544
R285 VOUT.n109 VOUT.n107 1.86544
R286 VOUT.n107 VOUT.n105 1.86544
R287 VOUT.n101 VOUT.n99 1.86544
R288 VOUT.n99 VOUT.n97 1.86544
R289 VOUT.n93 VOUT.n91 1.86544
R290 VOUT.n91 VOUT.n89 1.86544
R291 VOUT.n86 VOUT.n84 1.86544
R292 VOUT.n84 VOUT.n82 1.86544
R293 VOUT.n43 VOUT.n41 1.76774
R294 VOUT.n45 VOUT.n43 1.76774
R295 VOUT.n36 VOUT.n34 1.76774
R296 VOUT.n38 VOUT.n36 1.76774
R297 VOUT.n30 VOUT.n28 1.76774
R298 VOUT.n32 VOUT.n30 1.76774
R299 VOUT.n18 VOUT.n17 1.76774
R300 VOUT.n17 VOUT.n15 1.76774
R301 VOUT.n11 VOUT.n10 1.76774
R302 VOUT.n10 VOUT.n8 1.76774
R303 VOUT.n5 VOUT.n4 1.76774
R304 VOUT.n4 VOUT.n2 1.76774
R305 VOUT.n78 VOUT.n70 1.02924
R306 VOUT.n70 VOUT.n62 1.02924
R307 VOUT.n110 VOUT.n102 1.02924
R308 VOUT.n102 VOUT.n94 1.02924
R309 VOUT.n46 VOUT.n39 0.934408
R310 VOUT.n19 VOUT.n12 0.934408
R311 VOUT.n26 VOUT.n25 0.346423
R312 VOUT.n112 VOUT.n26 0.337725
R313 VOUT.n24 VOUT.n23 0.112999
R314 VOUT.n22 VOUT.n21 0.11058
R315 VOUT.n21 VOUT.t106 0.0671754
R316 VOUT.n22 VOUT.t107 0.0666091
R317 VOUT.n23 VOUT.t109 0.0664805
R318 VOUT.n24 VOUT.t108 0.0657554
R319 VOUT.n23 VOUT.n22 0.0595027
R320 VOUT.n25 VOUT.n21 0.0507907
R321 VOUT.n25 VOUT.n24 0.0111165
R322 VOUT VOUT.n112 0.0099
R323 VDD.n245 VDD.n196 500.488
R324 VDD.n4591 VDD.n198 500.488
R325 VDD.n4241 VDD.n537 500.488
R326 VDD.n543 VDD.n539 500.488
R327 VDD.n2843 VDD.n2842 500.488
R328 VDD.n2908 VDD.n1835 500.488
R329 VDD.n2247 VDD.n2223 500.488
R330 VDD.n2366 VDD.n2225 500.488
R331 VDD.n3818 VDD.n1035 323.416
R332 VDD.n4208 VDD.n696 323.416
R333 VDD.n4173 VDD.n4172 323.416
R334 VDD.n3598 VDD.n3387 323.416
R335 VDD.n3384 VDD.n1058 323.416
R336 VDD.n3344 VDD.n3343 323.416
R337 VDD.n1576 VDD.n1398 323.416
R338 VDD.n2963 VDD.n1400 323.416
R339 VDD.n4150 VDD.n4149 323.416
R340 VDD.n4218 VDD.n688 323.416
R341 VDD.n3612 VDD.n3599 323.416
R342 VDD.n3816 VDD.n3600 323.416
R343 VDD.n3329 VDD.n1037 323.416
R344 VDD.n3288 VDD.n3287 323.416
R345 VDD.n1626 VDD.n1399 323.416
R346 VDD.n2965 VDD.n1396 323.416
R347 VDD.t73 VDD.t78 261.51
R348 VDD.t162 VDD.t80 261.51
R349 VDD.n2906 VDD.t73 249.667
R350 VDD.n4242 VDD.t80 249.667
R351 VDD.n2304 VDD.t61 229.163
R352 VDD.n2326 VDD.t58 229.163
R353 VDD.n2260 VDD.t35 229.163
R354 VDD.n565 VDD.t55 229.163
R355 VDD.n575 VDD.t52 229.163
R356 VDD.n583 VDD.t31 229.163
R357 VDD.n218 VDD.t13 229.163
R358 VDD.n228 VDD.t10 229.163
R359 VDD.n237 VDD.t19 229.163
R360 VDD.n2871 VDD.t37 229.163
R361 VDD.n1814 VDD.t23 229.163
R362 VDD.n1832 VDD.t26 229.163
R363 VDD.n3609 VDD.t62 225.893
R364 VDD.n709 VDD.t39 225.893
R365 VDD.n3391 VDD.t66 225.893
R366 VDD.n684 VDD.t47 225.893
R367 VDD.n1409 VDD.t15 225.893
R368 VDD.n1061 VDD.t43 225.893
R369 VDD.n1623 VDD.t4 225.893
R370 VDD.n1079 VDD.t69 225.893
R371 VDD.n3609 VDD.t65 224.287
R372 VDD.n709 VDD.t41 224.287
R373 VDD.n3391 VDD.t68 224.287
R374 VDD.n684 VDD.t48 224.287
R375 VDD.n1409 VDD.t17 224.287
R376 VDD.n1061 VDD.t45 224.287
R377 VDD.n1623 VDD.t7 224.287
R378 VDD.n1079 VDD.t70 224.287
R379 VDD.n2304 VDD.t59 223.755
R380 VDD.n2326 VDD.t56 223.755
R381 VDD.n2260 VDD.t32 223.755
R382 VDD.n565 VDD.t53 223.755
R383 VDD.n575 VDD.t50 223.755
R384 VDD.n583 VDD.t28 223.755
R385 VDD.n218 VDD.t12 223.755
R386 VDD.n228 VDD.t8 223.755
R387 VDD.n237 VDD.t18 223.755
R388 VDD.n2871 VDD.t36 223.755
R389 VDD.n1814 VDD.t21 223.755
R390 VDD.n1832 VDD.t25 223.755
R391 VDD.t78 VDD.t74 215.438
R392 VDD.t74 VDD.t89 215.438
R393 VDD.t0 VDD.t87 215.438
R394 VDD.t87 VDD.t162 215.438
R395 VDD.n3330 VDD.n3329 185
R396 VDD.n3329 VDD.n1036 185
R397 VDD.n3331 VDD.n1069 185
R398 VDD.n3341 VDD.n1069 185
R399 VDD.n3332 VDD.n1077 185
R400 VDD.n1077 VDD.n1067 185
R401 VDD.n3334 VDD.n3333 185
R402 VDD.n3335 VDD.n3334 185
R403 VDD.n1078 VDD.n1076 185
R404 VDD.n1076 VDD.n1073 185
R405 VDD.n3268 VDD.n1086 185
R406 VDD.n3278 VDD.n1086 185
R407 VDD.n3269 VDD.n1094 185
R408 VDD.n1094 VDD.n1084 185
R409 VDD.n3271 VDD.n3270 185
R410 VDD.n3272 VDD.n3271 185
R411 VDD.n3267 VDD.n1093 185
R412 VDD.n1093 VDD.n1090 185
R413 VDD.n3266 VDD.n3265 185
R414 VDD.n3265 VDD.n3264 185
R415 VDD.n1096 VDD.n1095 185
R416 VDD.n1097 VDD.n1096 185
R417 VDD.n3257 VDD.n3256 185
R418 VDD.n3258 VDD.n3257 185
R419 VDD.n3255 VDD.n1105 185
R420 VDD.n1110 VDD.n1105 185
R421 VDD.n3254 VDD.n3253 185
R422 VDD.n3253 VDD.n3252 185
R423 VDD.n1107 VDD.n1106 185
R424 VDD.n1117 VDD.n1107 185
R425 VDD.n3245 VDD.n3244 185
R426 VDD.n3246 VDD.n3245 185
R427 VDD.n3243 VDD.n1118 185
R428 VDD.n1118 VDD.n1114 185
R429 VDD.n3242 VDD.n3241 185
R430 VDD.n3241 VDD.n3240 185
R431 VDD.n1120 VDD.n1119 185
R432 VDD.n1121 VDD.n1120 185
R433 VDD.n3233 VDD.n3232 185
R434 VDD.n3234 VDD.n3233 185
R435 VDD.n3231 VDD.n1130 185
R436 VDD.n1130 VDD.n1127 185
R437 VDD.n3230 VDD.n3229 185
R438 VDD.n3229 VDD.n3228 185
R439 VDD.n1132 VDD.n1131 185
R440 VDD.n1133 VDD.n1132 185
R441 VDD.n3221 VDD.n3220 185
R442 VDD.n3222 VDD.n3221 185
R443 VDD.n3219 VDD.n1142 185
R444 VDD.n1142 VDD.n1139 185
R445 VDD.n3218 VDD.n3217 185
R446 VDD.n3217 VDD.n3216 185
R447 VDD.n1144 VDD.n1143 185
R448 VDD.n1145 VDD.n1144 185
R449 VDD.n3209 VDD.n3208 185
R450 VDD.n3210 VDD.n3209 185
R451 VDD.n3207 VDD.n1154 185
R452 VDD.n1154 VDD.n1151 185
R453 VDD.n3206 VDD.n3205 185
R454 VDD.n3205 VDD.n3204 185
R455 VDD.n1156 VDD.n1155 185
R456 VDD.n1157 VDD.n1156 185
R457 VDD.n3197 VDD.n3196 185
R458 VDD.n3198 VDD.n3197 185
R459 VDD.n3195 VDD.n1166 185
R460 VDD.n1166 VDD.n1163 185
R461 VDD.n3194 VDD.n3193 185
R462 VDD.n3193 VDD.n3192 185
R463 VDD.n1168 VDD.n1167 185
R464 VDD.n1169 VDD.n1168 185
R465 VDD.n3185 VDD.n3184 185
R466 VDD.n3186 VDD.n3185 185
R467 VDD.n3183 VDD.n1178 185
R468 VDD.n1178 VDD.n1175 185
R469 VDD.n3182 VDD.n3181 185
R470 VDD.n3181 VDD.n3180 185
R471 VDD.n1180 VDD.n1179 185
R472 VDD.n1181 VDD.n1180 185
R473 VDD.n3173 VDD.n3172 185
R474 VDD.n3174 VDD.n3173 185
R475 VDD.n3171 VDD.n1190 185
R476 VDD.n1190 VDD.n1187 185
R477 VDD.n3170 VDD.n3169 185
R478 VDD.n3169 VDD.n3168 185
R479 VDD.n1192 VDD.n1191 185
R480 VDD.n1193 VDD.n1192 185
R481 VDD.n3161 VDD.n3160 185
R482 VDD.n3162 VDD.n3161 185
R483 VDD.n3159 VDD.n1202 185
R484 VDD.n1202 VDD.n1199 185
R485 VDD.n3158 VDD.n3157 185
R486 VDD.n3157 VDD.n3156 185
R487 VDD.n1204 VDD.n1203 185
R488 VDD.n1205 VDD.n1204 185
R489 VDD.n3149 VDD.n3148 185
R490 VDD.n3150 VDD.n3149 185
R491 VDD.n3147 VDD.n1214 185
R492 VDD.n1214 VDD.n1211 185
R493 VDD.n3146 VDD.n3145 185
R494 VDD.n3145 VDD.n3144 185
R495 VDD.n1216 VDD.n1215 185
R496 VDD.n1217 VDD.n1216 185
R497 VDD.n3137 VDD.n3136 185
R498 VDD.n3138 VDD.n3137 185
R499 VDD.n3135 VDD.n1226 185
R500 VDD.n1226 VDD.n1223 185
R501 VDD.n3134 VDD.n3133 185
R502 VDD.n3133 VDD.n3132 185
R503 VDD.n1228 VDD.n1227 185
R504 VDD.n1229 VDD.n1228 185
R505 VDD.n3125 VDD.n3124 185
R506 VDD.n3126 VDD.n3125 185
R507 VDD.n3123 VDD.n1238 185
R508 VDD.n1238 VDD.n1235 185
R509 VDD.n3122 VDD.n3121 185
R510 VDD.n3121 VDD.n3120 185
R511 VDD.n1240 VDD.n1239 185
R512 VDD.n1241 VDD.n1240 185
R513 VDD.n3113 VDD.n3112 185
R514 VDD.n3114 VDD.n3113 185
R515 VDD.n3111 VDD.n1250 185
R516 VDD.n1250 VDD.n1247 185
R517 VDD.n3110 VDD.n3109 185
R518 VDD.n3109 VDD.n3108 185
R519 VDD.n1252 VDD.n1251 185
R520 VDD.n1253 VDD.n1252 185
R521 VDD.n3101 VDD.n3100 185
R522 VDD.n3102 VDD.n3101 185
R523 VDD.n3099 VDD.n1262 185
R524 VDD.n1262 VDD.n1259 185
R525 VDD.n3098 VDD.n3097 185
R526 VDD.n3097 VDD.n3096 185
R527 VDD.n1264 VDD.n1263 185
R528 VDD.n1265 VDD.n1264 185
R529 VDD.n3089 VDD.n3088 185
R530 VDD.n3090 VDD.n3089 185
R531 VDD.n3087 VDD.n1274 185
R532 VDD.n1274 VDD.n1271 185
R533 VDD.n3086 VDD.n3085 185
R534 VDD.n3085 VDD.n3084 185
R535 VDD.n1276 VDD.n1275 185
R536 VDD.n1277 VDD.n1276 185
R537 VDD.n3077 VDD.n3076 185
R538 VDD.n3078 VDD.n3077 185
R539 VDD.n3075 VDD.n1285 185
R540 VDD.n1291 VDD.n1285 185
R541 VDD.n3074 VDD.n3073 185
R542 VDD.n3073 VDD.n3072 185
R543 VDD.n1287 VDD.n1286 185
R544 VDD.n1288 VDD.n1287 185
R545 VDD.n3065 VDD.n3064 185
R546 VDD.n3066 VDD.n3065 185
R547 VDD.n3063 VDD.n1298 185
R548 VDD.n1298 VDD.n1295 185
R549 VDD.n3062 VDD.n3061 185
R550 VDD.n3061 VDD.n3060 185
R551 VDD.n1300 VDD.n1299 185
R552 VDD.n1301 VDD.n1300 185
R553 VDD.n3053 VDD.n3052 185
R554 VDD.n3054 VDD.n3053 185
R555 VDD.n3051 VDD.n1310 185
R556 VDD.n1310 VDD.n1307 185
R557 VDD.n3050 VDD.n3049 185
R558 VDD.n3049 VDD.n3048 185
R559 VDD.n1312 VDD.n1311 185
R560 VDD.n1313 VDD.n1312 185
R561 VDD.n3041 VDD.n3040 185
R562 VDD.n3042 VDD.n3041 185
R563 VDD.n3039 VDD.n1322 185
R564 VDD.n1322 VDD.n1319 185
R565 VDD.n3038 VDD.n3037 185
R566 VDD.n3037 VDD.n3036 185
R567 VDD.n1324 VDD.n1323 185
R568 VDD.n1325 VDD.n1324 185
R569 VDD.n3029 VDD.n3028 185
R570 VDD.n3030 VDD.n3029 185
R571 VDD.n3027 VDD.n1334 185
R572 VDD.n1334 VDD.n1331 185
R573 VDD.n3026 VDD.n3025 185
R574 VDD.n3025 VDD.n3024 185
R575 VDD.n1336 VDD.n1335 185
R576 VDD.n1337 VDD.n1336 185
R577 VDD.n3017 VDD.n3016 185
R578 VDD.n3018 VDD.n3017 185
R579 VDD.n3015 VDD.n1346 185
R580 VDD.n1346 VDD.n1343 185
R581 VDD.n3014 VDD.n3013 185
R582 VDD.n3013 VDD.n3012 185
R583 VDD.n1348 VDD.n1347 185
R584 VDD.n1349 VDD.n1348 185
R585 VDD.n3005 VDD.n3004 185
R586 VDD.n3006 VDD.n3005 185
R587 VDD.n3003 VDD.n1358 185
R588 VDD.n1358 VDD.n1355 185
R589 VDD.n3002 VDD.n3001 185
R590 VDD.n3001 VDD.n3000 185
R591 VDD.n1360 VDD.n1359 185
R592 VDD.n1369 VDD.n1360 185
R593 VDD.n2993 VDD.n2992 185
R594 VDD.n2994 VDD.n2993 185
R595 VDD.n2991 VDD.n1370 185
R596 VDD.n1370 VDD.n1366 185
R597 VDD.n2990 VDD.n2989 185
R598 VDD.n2989 VDD.n2988 185
R599 VDD.n1372 VDD.n1371 185
R600 VDD.n1373 VDD.n1372 185
R601 VDD.n2981 VDD.n2980 185
R602 VDD.n2982 VDD.n2981 185
R603 VDD.n2979 VDD.n1382 185
R604 VDD.n1382 VDD.n1379 185
R605 VDD.n2978 VDD.n2977 185
R606 VDD.n2977 VDD.n2976 185
R607 VDD.n1384 VDD.n1383 185
R608 VDD.n1385 VDD.n1384 185
R609 VDD.n2969 VDD.n2968 185
R610 VDD.n2970 VDD.n2969 185
R611 VDD.n2967 VDD.n1394 185
R612 VDD.n1394 VDD.n1391 185
R613 VDD.n2966 VDD.n2965 185
R614 VDD.n2965 VDD.n2964 185
R615 VDD.n1396 VDD.n1395 185
R616 VDD.n1603 VDD.n1601 185
R617 VDD.n1606 VDD.n1605 185
R618 VDD.n1607 VDD.n1600 185
R619 VDD.n1609 VDD.n1608 185
R620 VDD.n1611 VDD.n1599 185
R621 VDD.n1614 VDD.n1613 185
R622 VDD.n1615 VDD.n1598 185
R623 VDD.n1617 VDD.n1616 185
R624 VDD.n1619 VDD.n1596 185
R625 VDD.n1803 VDD.n1802 185
R626 VDD.n1800 VDD.n1597 185
R627 VDD.n1799 VDD.n1798 185
R628 VDD.n1797 VDD.n1796 185
R629 VDD.n1795 VDD.n1621 185
R630 VDD.n1793 VDD.n1792 185
R631 VDD.n1791 VDD.n1622 185
R632 VDD.n1789 VDD.n1788 185
R633 VDD.n1786 VDD.n1625 185
R634 VDD.n1784 VDD.n1783 185
R635 VDD.n1782 VDD.n1626 185
R636 VDD.n1626 VDD.n1397 185
R637 VDD.n3289 VDD.n3288 185
R638 VDD.n3291 VDD.n3290 185
R639 VDD.n3293 VDD.n3292 185
R640 VDD.n3295 VDD.n3294 185
R641 VDD.n3297 VDD.n3296 185
R642 VDD.n3299 VDD.n3298 185
R643 VDD.n3301 VDD.n3300 185
R644 VDD.n3303 VDD.n3302 185
R645 VDD.n3305 VDD.n3304 185
R646 VDD.n3307 VDD.n3306 185
R647 VDD.n3309 VDD.n3308 185
R648 VDD.n3311 VDD.n3310 185
R649 VDD.n3313 VDD.n3312 185
R650 VDD.n3315 VDD.n3314 185
R651 VDD.n3317 VDD.n3316 185
R652 VDD.n3319 VDD.n3318 185
R653 VDD.n3321 VDD.n3320 185
R654 VDD.n3323 VDD.n3322 185
R655 VDD.n3325 VDD.n3324 185
R656 VDD.n3327 VDD.n3326 185
R657 VDD.n3328 VDD.n1037 185
R658 VDD.n3385 VDD.n1037 185
R659 VDD.n3287 VDD.n3286 185
R660 VDD.n3287 VDD.n1036 185
R661 VDD.n3285 VDD.n1068 185
R662 VDD.n3341 VDD.n1068 185
R663 VDD.n3284 VDD.n3283 185
R664 VDD.n3283 VDD.n1067 185
R665 VDD.n3282 VDD.n1075 185
R666 VDD.n3335 VDD.n1075 185
R667 VDD.n3281 VDD.n3280 185
R668 VDD.n3280 VDD.n1073 185
R669 VDD.n3279 VDD.n1082 185
R670 VDD.n3279 VDD.n3278 185
R671 VDD.n1627 VDD.n1083 185
R672 VDD.n1084 VDD.n1083 185
R673 VDD.n1628 VDD.n1092 185
R674 VDD.n3272 VDD.n1092 185
R675 VDD.n1630 VDD.n1629 185
R676 VDD.n1629 VDD.n1090 185
R677 VDD.n1631 VDD.n1099 185
R678 VDD.n3264 VDD.n1099 185
R679 VDD.n1633 VDD.n1632 185
R680 VDD.n1632 VDD.n1097 185
R681 VDD.n1634 VDD.n1104 185
R682 VDD.n3258 VDD.n1104 185
R683 VDD.n1636 VDD.n1635 185
R684 VDD.n1635 VDD.n1110 185
R685 VDD.n1637 VDD.n1109 185
R686 VDD.n3252 VDD.n1109 185
R687 VDD.n1639 VDD.n1638 185
R688 VDD.n1638 VDD.n1117 185
R689 VDD.n1640 VDD.n1116 185
R690 VDD.n3246 VDD.n1116 185
R691 VDD.n1642 VDD.n1641 185
R692 VDD.n1641 VDD.n1114 185
R693 VDD.n1643 VDD.n1123 185
R694 VDD.n3240 VDD.n1123 185
R695 VDD.n1645 VDD.n1644 185
R696 VDD.n1644 VDD.n1121 185
R697 VDD.n1646 VDD.n1129 185
R698 VDD.n3234 VDD.n1129 185
R699 VDD.n1648 VDD.n1647 185
R700 VDD.n1647 VDD.n1127 185
R701 VDD.n1649 VDD.n1135 185
R702 VDD.n3228 VDD.n1135 185
R703 VDD.n1651 VDD.n1650 185
R704 VDD.n1650 VDD.n1133 185
R705 VDD.n1652 VDD.n1141 185
R706 VDD.n3222 VDD.n1141 185
R707 VDD.n1654 VDD.n1653 185
R708 VDD.n1653 VDD.n1139 185
R709 VDD.n1655 VDD.n1147 185
R710 VDD.n3216 VDD.n1147 185
R711 VDD.n1657 VDD.n1656 185
R712 VDD.n1656 VDD.n1145 185
R713 VDD.n1658 VDD.n1153 185
R714 VDD.n3210 VDD.n1153 185
R715 VDD.n1660 VDD.n1659 185
R716 VDD.n1659 VDD.n1151 185
R717 VDD.n1661 VDD.n1159 185
R718 VDD.n3204 VDD.n1159 185
R719 VDD.n1663 VDD.n1662 185
R720 VDD.n1662 VDD.n1157 185
R721 VDD.n1664 VDD.n1165 185
R722 VDD.n3198 VDD.n1165 185
R723 VDD.n1666 VDD.n1665 185
R724 VDD.n1665 VDD.n1163 185
R725 VDD.n1667 VDD.n1171 185
R726 VDD.n3192 VDD.n1171 185
R727 VDD.n1669 VDD.n1668 185
R728 VDD.n1668 VDD.n1169 185
R729 VDD.n1670 VDD.n1177 185
R730 VDD.n3186 VDD.n1177 185
R731 VDD.n1672 VDD.n1671 185
R732 VDD.n1671 VDD.n1175 185
R733 VDD.n1673 VDD.n1183 185
R734 VDD.n3180 VDD.n1183 185
R735 VDD.n1675 VDD.n1674 185
R736 VDD.n1674 VDD.n1181 185
R737 VDD.n1676 VDD.n1189 185
R738 VDD.n3174 VDD.n1189 185
R739 VDD.n1678 VDD.n1677 185
R740 VDD.n1677 VDD.n1187 185
R741 VDD.n1679 VDD.n1195 185
R742 VDD.n3168 VDD.n1195 185
R743 VDD.n1681 VDD.n1680 185
R744 VDD.n1680 VDD.n1193 185
R745 VDD.n1682 VDD.n1201 185
R746 VDD.n3162 VDD.n1201 185
R747 VDD.n1684 VDD.n1683 185
R748 VDD.n1683 VDD.n1199 185
R749 VDD.n1685 VDD.n1207 185
R750 VDD.n3156 VDD.n1207 185
R751 VDD.n1687 VDD.n1686 185
R752 VDD.n1686 VDD.n1205 185
R753 VDD.n1688 VDD.n1213 185
R754 VDD.n3150 VDD.n1213 185
R755 VDD.n1690 VDD.n1689 185
R756 VDD.n1689 VDD.n1211 185
R757 VDD.n1691 VDD.n1219 185
R758 VDD.n3144 VDD.n1219 185
R759 VDD.n1693 VDD.n1692 185
R760 VDD.n1692 VDD.n1217 185
R761 VDD.n1694 VDD.n1225 185
R762 VDD.n3138 VDD.n1225 185
R763 VDD.n1696 VDD.n1695 185
R764 VDD.n1695 VDD.n1223 185
R765 VDD.n1697 VDD.n1231 185
R766 VDD.n3132 VDD.n1231 185
R767 VDD.n1699 VDD.n1698 185
R768 VDD.n1698 VDD.n1229 185
R769 VDD.n1700 VDD.n1237 185
R770 VDD.n3126 VDD.n1237 185
R771 VDD.n1702 VDD.n1701 185
R772 VDD.n1701 VDD.n1235 185
R773 VDD.n1703 VDD.n1243 185
R774 VDD.n3120 VDD.n1243 185
R775 VDD.n1705 VDD.n1704 185
R776 VDD.n1704 VDD.n1241 185
R777 VDD.n1706 VDD.n1249 185
R778 VDD.n3114 VDD.n1249 185
R779 VDD.n1708 VDD.n1707 185
R780 VDD.n1707 VDD.n1247 185
R781 VDD.n1709 VDD.n1255 185
R782 VDD.n3108 VDD.n1255 185
R783 VDD.n1711 VDD.n1710 185
R784 VDD.n1710 VDD.n1253 185
R785 VDD.n1712 VDD.n1261 185
R786 VDD.n3102 VDD.n1261 185
R787 VDD.n1714 VDD.n1713 185
R788 VDD.n1713 VDD.n1259 185
R789 VDD.n1715 VDD.n1267 185
R790 VDD.n3096 VDD.n1267 185
R791 VDD.n1717 VDD.n1716 185
R792 VDD.n1716 VDD.n1265 185
R793 VDD.n1718 VDD.n1273 185
R794 VDD.n3090 VDD.n1273 185
R795 VDD.n1720 VDD.n1719 185
R796 VDD.n1719 VDD.n1271 185
R797 VDD.n1721 VDD.n1279 185
R798 VDD.n3084 VDD.n1279 185
R799 VDD.n1723 VDD.n1722 185
R800 VDD.n1722 VDD.n1277 185
R801 VDD.n1724 VDD.n1284 185
R802 VDD.n3078 VDD.n1284 185
R803 VDD.n1726 VDD.n1725 185
R804 VDD.n1725 VDD.n1291 185
R805 VDD.n1727 VDD.n1290 185
R806 VDD.n3072 VDD.n1290 185
R807 VDD.n1729 VDD.n1728 185
R808 VDD.n1728 VDD.n1288 185
R809 VDD.n1730 VDD.n1297 185
R810 VDD.n3066 VDD.n1297 185
R811 VDD.n1732 VDD.n1731 185
R812 VDD.n1731 VDD.n1295 185
R813 VDD.n1733 VDD.n1303 185
R814 VDD.n3060 VDD.n1303 185
R815 VDD.n1735 VDD.n1734 185
R816 VDD.n1734 VDD.n1301 185
R817 VDD.n1736 VDD.n1309 185
R818 VDD.n3054 VDD.n1309 185
R819 VDD.n1738 VDD.n1737 185
R820 VDD.n1737 VDD.n1307 185
R821 VDD.n1739 VDD.n1315 185
R822 VDD.n3048 VDD.n1315 185
R823 VDD.n1741 VDD.n1740 185
R824 VDD.n1740 VDD.n1313 185
R825 VDD.n1742 VDD.n1321 185
R826 VDD.n3042 VDD.n1321 185
R827 VDD.n1744 VDD.n1743 185
R828 VDD.n1743 VDD.n1319 185
R829 VDD.n1745 VDD.n1327 185
R830 VDD.n3036 VDD.n1327 185
R831 VDD.n1747 VDD.n1746 185
R832 VDD.n1746 VDD.n1325 185
R833 VDD.n1748 VDD.n1333 185
R834 VDD.n3030 VDD.n1333 185
R835 VDD.n1750 VDD.n1749 185
R836 VDD.n1749 VDD.n1331 185
R837 VDD.n1751 VDD.n1339 185
R838 VDD.n3024 VDD.n1339 185
R839 VDD.n1753 VDD.n1752 185
R840 VDD.n1752 VDD.n1337 185
R841 VDD.n1754 VDD.n1345 185
R842 VDD.n3018 VDD.n1345 185
R843 VDD.n1756 VDD.n1755 185
R844 VDD.n1755 VDD.n1343 185
R845 VDD.n1757 VDD.n1351 185
R846 VDD.n3012 VDD.n1351 185
R847 VDD.n1759 VDD.n1758 185
R848 VDD.n1758 VDD.n1349 185
R849 VDD.n1760 VDD.n1357 185
R850 VDD.n3006 VDD.n1357 185
R851 VDD.n1762 VDD.n1761 185
R852 VDD.n1761 VDD.n1355 185
R853 VDD.n1763 VDD.n1362 185
R854 VDD.n3000 VDD.n1362 185
R855 VDD.n1765 VDD.n1764 185
R856 VDD.n1764 VDD.n1369 185
R857 VDD.n1766 VDD.n1368 185
R858 VDD.n2994 VDD.n1368 185
R859 VDD.n1768 VDD.n1767 185
R860 VDD.n1767 VDD.n1366 185
R861 VDD.n1769 VDD.n1375 185
R862 VDD.n2988 VDD.n1375 185
R863 VDD.n1771 VDD.n1770 185
R864 VDD.n1770 VDD.n1373 185
R865 VDD.n1772 VDD.n1381 185
R866 VDD.n2982 VDD.n1381 185
R867 VDD.n1774 VDD.n1773 185
R868 VDD.n1773 VDD.n1379 185
R869 VDD.n1775 VDD.n1387 185
R870 VDD.n2976 VDD.n1387 185
R871 VDD.n1777 VDD.n1776 185
R872 VDD.n1776 VDD.n1385 185
R873 VDD.n1778 VDD.n1393 185
R874 VDD.n2970 VDD.n1393 185
R875 VDD.n1780 VDD.n1779 185
R876 VDD.n1779 VDD.n1391 185
R877 VDD.n1781 VDD.n1399 185
R878 VDD.n2964 VDD.n1399 185
R879 VDD.n4151 VDD.n4150 185
R880 VDD.n4150 VDD.n693 185
R881 VDD.n4152 VDD.n694 185
R882 VDD.n4213 VDD.n694 185
R883 VDD.n4154 VDD.n4153 185
R884 VDD.n4153 VDD.n691 185
R885 VDD.n4155 VDD.n719 185
R886 VDD.n4165 VDD.n719 185
R887 VDD.n4156 VDD.n727 185
R888 VDD.n727 VDD.n717 185
R889 VDD.n4158 VDD.n4157 185
R890 VDD.n4159 VDD.n4158 185
R891 VDD.n4126 VDD.n726 185
R892 VDD.n726 VDD.n723 185
R893 VDD.n4125 VDD.n4124 185
R894 VDD.n4124 VDD.n4123 185
R895 VDD.n729 VDD.n728 185
R896 VDD.n730 VDD.n729 185
R897 VDD.n4116 VDD.n4115 185
R898 VDD.n4117 VDD.n4116 185
R899 VDD.n4114 VDD.n739 185
R900 VDD.n739 VDD.n736 185
R901 VDD.n4113 VDD.n4112 185
R902 VDD.n4112 VDD.n4111 185
R903 VDD.n741 VDD.n740 185
R904 VDD.n750 VDD.n741 185
R905 VDD.n4104 VDD.n4103 185
R906 VDD.n4105 VDD.n4104 185
R907 VDD.n4102 VDD.n751 185
R908 VDD.n751 VDD.n747 185
R909 VDD.n4101 VDD.n4100 185
R910 VDD.n4100 VDD.n4099 185
R911 VDD.n753 VDD.n752 185
R912 VDD.n754 VDD.n753 185
R913 VDD.n4092 VDD.n4091 185
R914 VDD.n4093 VDD.n4092 185
R915 VDD.n4090 VDD.n763 185
R916 VDD.n763 VDD.n760 185
R917 VDD.n4089 VDD.n4088 185
R918 VDD.n4088 VDD.n4087 185
R919 VDD.n765 VDD.n764 185
R920 VDD.n766 VDD.n765 185
R921 VDD.n4080 VDD.n4079 185
R922 VDD.n4081 VDD.n4080 185
R923 VDD.n4078 VDD.n775 185
R924 VDD.n775 VDD.n772 185
R925 VDD.n4077 VDD.n4076 185
R926 VDD.n4076 VDD.n4075 185
R927 VDD.n777 VDD.n776 185
R928 VDD.n778 VDD.n777 185
R929 VDD.n4068 VDD.n4067 185
R930 VDD.n4069 VDD.n4068 185
R931 VDD.n4066 VDD.n787 185
R932 VDD.n787 VDD.n784 185
R933 VDD.n4065 VDD.n4064 185
R934 VDD.n4064 VDD.n4063 185
R935 VDD.n789 VDD.n788 185
R936 VDD.n790 VDD.n789 185
R937 VDD.n4056 VDD.n4055 185
R938 VDD.n4057 VDD.n4056 185
R939 VDD.n4054 VDD.n799 185
R940 VDD.n799 VDD.n796 185
R941 VDD.n4053 VDD.n4052 185
R942 VDD.n4052 VDD.n4051 185
R943 VDD.n801 VDD.n800 185
R944 VDD.n802 VDD.n801 185
R945 VDD.n4044 VDD.n4043 185
R946 VDD.n4045 VDD.n4044 185
R947 VDD.n4042 VDD.n811 185
R948 VDD.n811 VDD.n808 185
R949 VDD.n4041 VDD.n4040 185
R950 VDD.n4040 VDD.n4039 185
R951 VDD.n813 VDD.n812 185
R952 VDD.n814 VDD.n813 185
R953 VDD.n4032 VDD.n4031 185
R954 VDD.n4033 VDD.n4032 185
R955 VDD.n4030 VDD.n822 185
R956 VDD.n828 VDD.n822 185
R957 VDD.n4029 VDD.n4028 185
R958 VDD.n4028 VDD.n4027 185
R959 VDD.n824 VDD.n823 185
R960 VDD.n825 VDD.n824 185
R961 VDD.n4020 VDD.n4019 185
R962 VDD.n4021 VDD.n4020 185
R963 VDD.n4018 VDD.n835 185
R964 VDD.n835 VDD.n832 185
R965 VDD.n4017 VDD.n4016 185
R966 VDD.n4016 VDD.n4015 185
R967 VDD.n837 VDD.n836 185
R968 VDD.n838 VDD.n837 185
R969 VDD.n4008 VDD.n4007 185
R970 VDD.n4009 VDD.n4008 185
R971 VDD.n4006 VDD.n847 185
R972 VDD.n847 VDD.n844 185
R973 VDD.n4005 VDD.n4004 185
R974 VDD.n4004 VDD.n4003 185
R975 VDD.n849 VDD.n848 185
R976 VDD.n850 VDD.n849 185
R977 VDD.n3996 VDD.n3995 185
R978 VDD.n3997 VDD.n3996 185
R979 VDD.n3994 VDD.n859 185
R980 VDD.n859 VDD.n856 185
R981 VDD.n3993 VDD.n3992 185
R982 VDD.n3992 VDD.n3991 185
R983 VDD.n861 VDD.n860 185
R984 VDD.n862 VDD.n861 185
R985 VDD.n3984 VDD.n3983 185
R986 VDD.n3985 VDD.n3984 185
R987 VDD.n3982 VDD.n871 185
R988 VDD.n871 VDD.n868 185
R989 VDD.n3981 VDD.n3980 185
R990 VDD.n3980 VDD.n3979 185
R991 VDD.n873 VDD.n872 185
R992 VDD.n874 VDD.n873 185
R993 VDD.n3972 VDD.n3971 185
R994 VDD.n3973 VDD.n3972 185
R995 VDD.n3970 VDD.n883 185
R996 VDD.n883 VDD.n880 185
R997 VDD.n3969 VDD.n3968 185
R998 VDD.n3968 VDD.n3967 185
R999 VDD.n885 VDD.n884 185
R1000 VDD.n886 VDD.n885 185
R1001 VDD.n3960 VDD.n3959 185
R1002 VDD.n3961 VDD.n3960 185
R1003 VDD.n3958 VDD.n895 185
R1004 VDD.n895 VDD.n892 185
R1005 VDD.n3957 VDD.n3956 185
R1006 VDD.n3956 VDD.n3955 185
R1007 VDD.n897 VDD.n896 185
R1008 VDD.n898 VDD.n897 185
R1009 VDD.n3948 VDD.n3947 185
R1010 VDD.n3949 VDD.n3948 185
R1011 VDD.n3946 VDD.n907 185
R1012 VDD.n907 VDD.n904 185
R1013 VDD.n3945 VDD.n3944 185
R1014 VDD.n3944 VDD.n3943 185
R1015 VDD.n909 VDD.n908 185
R1016 VDD.n910 VDD.n909 185
R1017 VDD.n3936 VDD.n3935 185
R1018 VDD.n3937 VDD.n3936 185
R1019 VDD.n3934 VDD.n919 185
R1020 VDD.n919 VDD.n916 185
R1021 VDD.n3933 VDD.n3932 185
R1022 VDD.n3932 VDD.n3931 185
R1023 VDD.n921 VDD.n920 185
R1024 VDD.n922 VDD.n921 185
R1025 VDD.n3924 VDD.n3923 185
R1026 VDD.n3925 VDD.n3924 185
R1027 VDD.n3922 VDD.n931 185
R1028 VDD.n931 VDD.n928 185
R1029 VDD.n3921 VDD.n3920 185
R1030 VDD.n3920 VDD.n3919 185
R1031 VDD.n933 VDD.n932 185
R1032 VDD.n934 VDD.n933 185
R1033 VDD.n3912 VDD.n3911 185
R1034 VDD.n3913 VDD.n3912 185
R1035 VDD.n3910 VDD.n943 185
R1036 VDD.n943 VDD.n940 185
R1037 VDD.n3909 VDD.n3908 185
R1038 VDD.n3908 VDD.n3907 185
R1039 VDD.n945 VDD.n944 185
R1040 VDD.n946 VDD.n945 185
R1041 VDD.n3900 VDD.n3899 185
R1042 VDD.n3901 VDD.n3900 185
R1043 VDD.n3898 VDD.n955 185
R1044 VDD.n955 VDD.n952 185
R1045 VDD.n3897 VDD.n3896 185
R1046 VDD.n3896 VDD.n3895 185
R1047 VDD.n957 VDD.n956 185
R1048 VDD.n958 VDD.n957 185
R1049 VDD.n3888 VDD.n3887 185
R1050 VDD.n3889 VDD.n3888 185
R1051 VDD.n3886 VDD.n967 185
R1052 VDD.n967 VDD.n964 185
R1053 VDD.n3885 VDD.n3884 185
R1054 VDD.n3884 VDD.n3883 185
R1055 VDD.n969 VDD.n968 185
R1056 VDD.n970 VDD.n969 185
R1057 VDD.n3876 VDD.n3875 185
R1058 VDD.n3877 VDD.n3876 185
R1059 VDD.n3874 VDD.n979 185
R1060 VDD.n979 VDD.n976 185
R1061 VDD.n3873 VDD.n3872 185
R1062 VDD.n3872 VDD.n3871 185
R1063 VDD.n981 VDD.n980 185
R1064 VDD.n982 VDD.n981 185
R1065 VDD.n3864 VDD.n3863 185
R1066 VDD.n3865 VDD.n3864 185
R1067 VDD.n3862 VDD.n991 185
R1068 VDD.n991 VDD.n988 185
R1069 VDD.n3861 VDD.n3860 185
R1070 VDD.n3860 VDD.n3859 185
R1071 VDD.n993 VDD.n992 185
R1072 VDD.n1001 VDD.n993 185
R1073 VDD.n3852 VDD.n3851 185
R1074 VDD.n3853 VDD.n3852 185
R1075 VDD.n3850 VDD.n1002 185
R1076 VDD.n1008 VDD.n1002 185
R1077 VDD.n3849 VDD.n3848 185
R1078 VDD.n3848 VDD.n3847 185
R1079 VDD.n1004 VDD.n1003 185
R1080 VDD.n1005 VDD.n1004 185
R1081 VDD.n3840 VDD.n3839 185
R1082 VDD.n3841 VDD.n3840 185
R1083 VDD.n3838 VDD.n1015 185
R1084 VDD.n1015 VDD.n1012 185
R1085 VDD.n3837 VDD.n3836 185
R1086 VDD.n3836 VDD.n3835 185
R1087 VDD.n1017 VDD.n1016 185
R1088 VDD.n1018 VDD.n1017 185
R1089 VDD.n3828 VDD.n3827 185
R1090 VDD.n3829 VDD.n3828 185
R1091 VDD.n3826 VDD.n1027 185
R1092 VDD.n1027 VDD.n1024 185
R1093 VDD.n3825 VDD.n3824 185
R1094 VDD.n3824 VDD.n3823 185
R1095 VDD.n1029 VDD.n1028 185
R1096 VDD.n1030 VDD.n1029 185
R1097 VDD.n3816 VDD.n3815 185
R1098 VDD.n3817 VDD.n3816 185
R1099 VDD.n3814 VDD.n3600 185
R1100 VDD.n3813 VDD.n3812 185
R1101 VDD.n3810 VDD.n3601 185
R1102 VDD.n3808 VDD.n3807 185
R1103 VDD.n3806 VDD.n3602 185
R1104 VDD.n3805 VDD.n3804 185
R1105 VDD.n3802 VDD.n3603 185
R1106 VDD.n3800 VDD.n3799 185
R1107 VDD.n3798 VDD.n3604 185
R1108 VDD.n3797 VDD.n3796 185
R1109 VDD.n3794 VDD.n3605 185
R1110 VDD.n3792 VDD.n3791 185
R1111 VDD.n3790 VDD.n3606 185
R1112 VDD.n3789 VDD.n3788 185
R1113 VDD.n3786 VDD.n3607 185
R1114 VDD.n3784 VDD.n3783 185
R1115 VDD.n3782 VDD.n3608 185
R1116 VDD.n3780 VDD.n3779 185
R1117 VDD.n3777 VDD.n3611 185
R1118 VDD.n3775 VDD.n3774 185
R1119 VDD.n3773 VDD.n3612 185
R1120 VDD.n3612 VDD.n3386 185
R1121 VDD.n4218 VDD.n4217 185
R1122 VDD.n4220 VDD.n686 185
R1123 VDD.n4222 VDD.n4221 185
R1124 VDD.n4223 VDD.n683 185
R1125 VDD.n4226 VDD.n4225 185
R1126 VDD.n4228 VDD.n681 185
R1127 VDD.n4230 VDD.n4229 185
R1128 VDD.n4231 VDD.n680 185
R1129 VDD.n4233 VDD.n4232 185
R1130 VDD.n4235 VDD.n677 185
R1131 VDD.n4237 VDD.n4236 185
R1132 VDD.n4134 VDD.n676 185
R1133 VDD.n4136 VDD.n4135 185
R1134 VDD.n4137 VDD.n4132 185
R1135 VDD.n4139 VDD.n4138 185
R1136 VDD.n4141 VDD.n4130 185
R1137 VDD.n4143 VDD.n4142 185
R1138 VDD.n4144 VDD.n4129 185
R1139 VDD.n4146 VDD.n4145 185
R1140 VDD.n4148 VDD.n4128 185
R1141 VDD.n4149 VDD.n4127 185
R1142 VDD.n4149 VDD.n679 185
R1143 VDD.n4216 VDD.n688 185
R1144 VDD.n693 VDD.n688 185
R1145 VDD.n4215 VDD.n4214 185
R1146 VDD.n4214 VDD.n4213 185
R1147 VDD.n690 VDD.n689 185
R1148 VDD.n691 VDD.n690 185
R1149 VDD.n3613 VDD.n718 185
R1150 VDD.n4165 VDD.n718 185
R1151 VDD.n3615 VDD.n3614 185
R1152 VDD.n3614 VDD.n717 185
R1153 VDD.n3616 VDD.n725 185
R1154 VDD.n4159 VDD.n725 185
R1155 VDD.n3618 VDD.n3617 185
R1156 VDD.n3617 VDD.n723 185
R1157 VDD.n3619 VDD.n732 185
R1158 VDD.n4123 VDD.n732 185
R1159 VDD.n3621 VDD.n3620 185
R1160 VDD.n3620 VDD.n730 185
R1161 VDD.n3622 VDD.n738 185
R1162 VDD.n4117 VDD.n738 185
R1163 VDD.n3624 VDD.n3623 185
R1164 VDD.n3623 VDD.n736 185
R1165 VDD.n3625 VDD.n743 185
R1166 VDD.n4111 VDD.n743 185
R1167 VDD.n3627 VDD.n3626 185
R1168 VDD.n3626 VDD.n750 185
R1169 VDD.n3628 VDD.n749 185
R1170 VDD.n4105 VDD.n749 185
R1171 VDD.n3630 VDD.n3629 185
R1172 VDD.n3629 VDD.n747 185
R1173 VDD.n3631 VDD.n756 185
R1174 VDD.n4099 VDD.n756 185
R1175 VDD.n3633 VDD.n3632 185
R1176 VDD.n3632 VDD.n754 185
R1177 VDD.n3634 VDD.n762 185
R1178 VDD.n4093 VDD.n762 185
R1179 VDD.n3636 VDD.n3635 185
R1180 VDD.n3635 VDD.n760 185
R1181 VDD.n3637 VDD.n768 185
R1182 VDD.n4087 VDD.n768 185
R1183 VDD.n3639 VDD.n3638 185
R1184 VDD.n3638 VDD.n766 185
R1185 VDD.n3640 VDD.n774 185
R1186 VDD.n4081 VDD.n774 185
R1187 VDD.n3642 VDD.n3641 185
R1188 VDD.n3641 VDD.n772 185
R1189 VDD.n3643 VDD.n780 185
R1190 VDD.n4075 VDD.n780 185
R1191 VDD.n3645 VDD.n3644 185
R1192 VDD.n3644 VDD.n778 185
R1193 VDD.n3646 VDD.n786 185
R1194 VDD.n4069 VDD.n786 185
R1195 VDD.n3648 VDD.n3647 185
R1196 VDD.n3647 VDD.n784 185
R1197 VDD.n3649 VDD.n792 185
R1198 VDD.n4063 VDD.n792 185
R1199 VDD.n3651 VDD.n3650 185
R1200 VDD.n3650 VDD.n790 185
R1201 VDD.n3652 VDD.n798 185
R1202 VDD.n4057 VDD.n798 185
R1203 VDD.n3654 VDD.n3653 185
R1204 VDD.n3653 VDD.n796 185
R1205 VDD.n3655 VDD.n804 185
R1206 VDD.n4051 VDD.n804 185
R1207 VDD.n3657 VDD.n3656 185
R1208 VDD.n3656 VDD.n802 185
R1209 VDD.n3658 VDD.n810 185
R1210 VDD.n4045 VDD.n810 185
R1211 VDD.n3660 VDD.n3659 185
R1212 VDD.n3659 VDD.n808 185
R1213 VDD.n3661 VDD.n816 185
R1214 VDD.n4039 VDD.n816 185
R1215 VDD.n3663 VDD.n3662 185
R1216 VDD.n3662 VDD.n814 185
R1217 VDD.n3664 VDD.n821 185
R1218 VDD.n4033 VDD.n821 185
R1219 VDD.n3666 VDD.n3665 185
R1220 VDD.n3665 VDD.n828 185
R1221 VDD.n3667 VDD.n827 185
R1222 VDD.n4027 VDD.n827 185
R1223 VDD.n3669 VDD.n3668 185
R1224 VDD.n3668 VDD.n825 185
R1225 VDD.n3670 VDD.n834 185
R1226 VDD.n4021 VDD.n834 185
R1227 VDD.n3672 VDD.n3671 185
R1228 VDD.n3671 VDD.n832 185
R1229 VDD.n3673 VDD.n840 185
R1230 VDD.n4015 VDD.n840 185
R1231 VDD.n3675 VDD.n3674 185
R1232 VDD.n3674 VDD.n838 185
R1233 VDD.n3676 VDD.n846 185
R1234 VDD.n4009 VDD.n846 185
R1235 VDD.n3678 VDD.n3677 185
R1236 VDD.n3677 VDD.n844 185
R1237 VDD.n3679 VDD.n852 185
R1238 VDD.n4003 VDD.n852 185
R1239 VDD.n3681 VDD.n3680 185
R1240 VDD.n3680 VDD.n850 185
R1241 VDD.n3682 VDD.n858 185
R1242 VDD.n3997 VDD.n858 185
R1243 VDD.n3684 VDD.n3683 185
R1244 VDD.n3683 VDD.n856 185
R1245 VDD.n3685 VDD.n864 185
R1246 VDD.n3991 VDD.n864 185
R1247 VDD.n3687 VDD.n3686 185
R1248 VDD.n3686 VDD.n862 185
R1249 VDD.n3688 VDD.n870 185
R1250 VDD.n3985 VDD.n870 185
R1251 VDD.n3690 VDD.n3689 185
R1252 VDD.n3689 VDD.n868 185
R1253 VDD.n3691 VDD.n876 185
R1254 VDD.n3979 VDD.n876 185
R1255 VDD.n3693 VDD.n3692 185
R1256 VDD.n3692 VDD.n874 185
R1257 VDD.n3694 VDD.n882 185
R1258 VDD.n3973 VDD.n882 185
R1259 VDD.n3696 VDD.n3695 185
R1260 VDD.n3695 VDD.n880 185
R1261 VDD.n3697 VDD.n888 185
R1262 VDD.n3967 VDD.n888 185
R1263 VDD.n3699 VDD.n3698 185
R1264 VDD.n3698 VDD.n886 185
R1265 VDD.n3700 VDD.n894 185
R1266 VDD.n3961 VDD.n894 185
R1267 VDD.n3702 VDD.n3701 185
R1268 VDD.n3701 VDD.n892 185
R1269 VDD.n3703 VDD.n900 185
R1270 VDD.n3955 VDD.n900 185
R1271 VDD.n3705 VDD.n3704 185
R1272 VDD.n3704 VDD.n898 185
R1273 VDD.n3706 VDD.n906 185
R1274 VDD.n3949 VDD.n906 185
R1275 VDD.n3708 VDD.n3707 185
R1276 VDD.n3707 VDD.n904 185
R1277 VDD.n3709 VDD.n912 185
R1278 VDD.n3943 VDD.n912 185
R1279 VDD.n3711 VDD.n3710 185
R1280 VDD.n3710 VDD.n910 185
R1281 VDD.n3712 VDD.n918 185
R1282 VDD.n3937 VDD.n918 185
R1283 VDD.n3714 VDD.n3713 185
R1284 VDD.n3713 VDD.n916 185
R1285 VDD.n3715 VDD.n924 185
R1286 VDD.n3931 VDD.n924 185
R1287 VDD.n3717 VDD.n3716 185
R1288 VDD.n3716 VDD.n922 185
R1289 VDD.n3718 VDD.n930 185
R1290 VDD.n3925 VDD.n930 185
R1291 VDD.n3720 VDD.n3719 185
R1292 VDD.n3719 VDD.n928 185
R1293 VDD.n3721 VDD.n936 185
R1294 VDD.n3919 VDD.n936 185
R1295 VDD.n3723 VDD.n3722 185
R1296 VDD.n3722 VDD.n934 185
R1297 VDD.n3724 VDD.n942 185
R1298 VDD.n3913 VDD.n942 185
R1299 VDD.n3726 VDD.n3725 185
R1300 VDD.n3725 VDD.n940 185
R1301 VDD.n3727 VDD.n948 185
R1302 VDD.n3907 VDD.n948 185
R1303 VDD.n3729 VDD.n3728 185
R1304 VDD.n3728 VDD.n946 185
R1305 VDD.n3730 VDD.n954 185
R1306 VDD.n3901 VDD.n954 185
R1307 VDD.n3732 VDD.n3731 185
R1308 VDD.n3731 VDD.n952 185
R1309 VDD.n3733 VDD.n960 185
R1310 VDD.n3895 VDD.n960 185
R1311 VDD.n3735 VDD.n3734 185
R1312 VDD.n3734 VDD.n958 185
R1313 VDD.n3736 VDD.n966 185
R1314 VDD.n3889 VDD.n966 185
R1315 VDD.n3738 VDD.n3737 185
R1316 VDD.n3737 VDD.n964 185
R1317 VDD.n3739 VDD.n972 185
R1318 VDD.n3883 VDD.n972 185
R1319 VDD.n3741 VDD.n3740 185
R1320 VDD.n3740 VDD.n970 185
R1321 VDD.n3742 VDD.n978 185
R1322 VDD.n3877 VDD.n978 185
R1323 VDD.n3744 VDD.n3743 185
R1324 VDD.n3743 VDD.n976 185
R1325 VDD.n3745 VDD.n984 185
R1326 VDD.n3871 VDD.n984 185
R1327 VDD.n3747 VDD.n3746 185
R1328 VDD.n3746 VDD.n982 185
R1329 VDD.n3748 VDD.n990 185
R1330 VDD.n3865 VDD.n990 185
R1331 VDD.n3750 VDD.n3749 185
R1332 VDD.n3749 VDD.n988 185
R1333 VDD.n3751 VDD.n995 185
R1334 VDD.n3859 VDD.n995 185
R1335 VDD.n3753 VDD.n3752 185
R1336 VDD.n3752 VDD.n1001 185
R1337 VDD.n3754 VDD.n1000 185
R1338 VDD.n3853 VDD.n1000 185
R1339 VDD.n3756 VDD.n3755 185
R1340 VDD.n3755 VDD.n1008 185
R1341 VDD.n3757 VDD.n1007 185
R1342 VDD.n3847 VDD.n1007 185
R1343 VDD.n3759 VDD.n3758 185
R1344 VDD.n3758 VDD.n1005 185
R1345 VDD.n3760 VDD.n1014 185
R1346 VDD.n3841 VDD.n1014 185
R1347 VDD.n3762 VDD.n3761 185
R1348 VDD.n3761 VDD.n1012 185
R1349 VDD.n3763 VDD.n1020 185
R1350 VDD.n3835 VDD.n1020 185
R1351 VDD.n3765 VDD.n3764 185
R1352 VDD.n3764 VDD.n1018 185
R1353 VDD.n3766 VDD.n1026 185
R1354 VDD.n3829 VDD.n1026 185
R1355 VDD.n3768 VDD.n3767 185
R1356 VDD.n3767 VDD.n1024 185
R1357 VDD.n3769 VDD.n1032 185
R1358 VDD.n3823 VDD.n1032 185
R1359 VDD.n3771 VDD.n3770 185
R1360 VDD.n3770 VDD.n1030 185
R1361 VDD.n3772 VDD.n3599 185
R1362 VDD.n3817 VDD.n3599 185
R1363 VDD.n1060 VDD.n1058 185
R1364 VDD.n1058 VDD.n1036 185
R1365 VDD.n3340 VDD.n3339 185
R1366 VDD.n3341 VDD.n3340 185
R1367 VDD.n3338 VDD.n1070 185
R1368 VDD.n1070 VDD.n1067 185
R1369 VDD.n3337 VDD.n3336 185
R1370 VDD.n3336 VDD.n3335 185
R1371 VDD.n1072 VDD.n1071 185
R1372 VDD.n1073 VDD.n1072 185
R1373 VDD.n3277 VDD.n3276 185
R1374 VDD.n3278 VDD.n3277 185
R1375 VDD.n3275 VDD.n1087 185
R1376 VDD.n1087 VDD.n1084 185
R1377 VDD.n3274 VDD.n3273 185
R1378 VDD.n3273 VDD.n3272 185
R1379 VDD.n1089 VDD.n1088 185
R1380 VDD.n1090 VDD.n1089 185
R1381 VDD.n3263 VDD.n3262 185
R1382 VDD.n3264 VDD.n3263 185
R1383 VDD.n3261 VDD.n1100 185
R1384 VDD.n1100 VDD.n1097 185
R1385 VDD.n3260 VDD.n3259 185
R1386 VDD.n3259 VDD.n3258 185
R1387 VDD.n1102 VDD.n1101 185
R1388 VDD.n1110 VDD.n1102 185
R1389 VDD.n3251 VDD.n3250 185
R1390 VDD.n3252 VDD.n3251 185
R1391 VDD.n3249 VDD.n1111 185
R1392 VDD.n1117 VDD.n1111 185
R1393 VDD.n3248 VDD.n3247 185
R1394 VDD.n3247 VDD.n3246 185
R1395 VDD.n1113 VDD.n1112 185
R1396 VDD.n1114 VDD.n1113 185
R1397 VDD.n3239 VDD.n3238 185
R1398 VDD.n3240 VDD.n3239 185
R1399 VDD.n3237 VDD.n1124 185
R1400 VDD.n1124 VDD.n1121 185
R1401 VDD.n3236 VDD.n3235 185
R1402 VDD.n3235 VDD.n3234 185
R1403 VDD.n1126 VDD.n1125 185
R1404 VDD.n1127 VDD.n1126 185
R1405 VDD.n3227 VDD.n3226 185
R1406 VDD.n3228 VDD.n3227 185
R1407 VDD.n3225 VDD.n1136 185
R1408 VDD.n1136 VDD.n1133 185
R1409 VDD.n3224 VDD.n3223 185
R1410 VDD.n3223 VDD.n3222 185
R1411 VDD.n1138 VDD.n1137 185
R1412 VDD.n1139 VDD.n1138 185
R1413 VDD.n3215 VDD.n3214 185
R1414 VDD.n3216 VDD.n3215 185
R1415 VDD.n3213 VDD.n1148 185
R1416 VDD.n1148 VDD.n1145 185
R1417 VDD.n3212 VDD.n3211 185
R1418 VDD.n3211 VDD.n3210 185
R1419 VDD.n1150 VDD.n1149 185
R1420 VDD.n1151 VDD.n1150 185
R1421 VDD.n3203 VDD.n3202 185
R1422 VDD.n3204 VDD.n3203 185
R1423 VDD.n3201 VDD.n1160 185
R1424 VDD.n1160 VDD.n1157 185
R1425 VDD.n3200 VDD.n3199 185
R1426 VDD.n3199 VDD.n3198 185
R1427 VDD.n1162 VDD.n1161 185
R1428 VDD.n1163 VDD.n1162 185
R1429 VDD.n3191 VDD.n3190 185
R1430 VDD.n3192 VDD.n3191 185
R1431 VDD.n3189 VDD.n1172 185
R1432 VDD.n1172 VDD.n1169 185
R1433 VDD.n3188 VDD.n3187 185
R1434 VDD.n3187 VDD.n3186 185
R1435 VDD.n1174 VDD.n1173 185
R1436 VDD.n1175 VDD.n1174 185
R1437 VDD.n3179 VDD.n3178 185
R1438 VDD.n3180 VDD.n3179 185
R1439 VDD.n3177 VDD.n1184 185
R1440 VDD.n1184 VDD.n1181 185
R1441 VDD.n3176 VDD.n3175 185
R1442 VDD.n3175 VDD.n3174 185
R1443 VDD.n1186 VDD.n1185 185
R1444 VDD.n1187 VDD.n1186 185
R1445 VDD.n3167 VDD.n3166 185
R1446 VDD.n3168 VDD.n3167 185
R1447 VDD.n3165 VDD.n1196 185
R1448 VDD.n1196 VDD.n1193 185
R1449 VDD.n3164 VDD.n3163 185
R1450 VDD.n3163 VDD.n3162 185
R1451 VDD.n1198 VDD.n1197 185
R1452 VDD.n1199 VDD.n1198 185
R1453 VDD.n3155 VDD.n3154 185
R1454 VDD.n3156 VDD.n3155 185
R1455 VDD.n3153 VDD.n1208 185
R1456 VDD.n1208 VDD.n1205 185
R1457 VDD.n3152 VDD.n3151 185
R1458 VDD.n3151 VDD.n3150 185
R1459 VDD.n1210 VDD.n1209 185
R1460 VDD.n1211 VDD.n1210 185
R1461 VDD.n3143 VDD.n3142 185
R1462 VDD.n3144 VDD.n3143 185
R1463 VDD.n3141 VDD.n1220 185
R1464 VDD.n1220 VDD.n1217 185
R1465 VDD.n3140 VDD.n3139 185
R1466 VDD.n3139 VDD.n3138 185
R1467 VDD.n1222 VDD.n1221 185
R1468 VDD.n1223 VDD.n1222 185
R1469 VDD.n3131 VDD.n3130 185
R1470 VDD.n3132 VDD.n3131 185
R1471 VDD.n3129 VDD.n1232 185
R1472 VDD.n1232 VDD.n1229 185
R1473 VDD.n3128 VDD.n3127 185
R1474 VDD.n3127 VDD.n3126 185
R1475 VDD.n1234 VDD.n1233 185
R1476 VDD.n1235 VDD.n1234 185
R1477 VDD.n3119 VDD.n3118 185
R1478 VDD.n3120 VDD.n3119 185
R1479 VDD.n3117 VDD.n1244 185
R1480 VDD.n1244 VDD.n1241 185
R1481 VDD.n3116 VDD.n3115 185
R1482 VDD.n3115 VDD.n3114 185
R1483 VDD.n1246 VDD.n1245 185
R1484 VDD.n1247 VDD.n1246 185
R1485 VDD.n3107 VDD.n3106 185
R1486 VDD.n3108 VDD.n3107 185
R1487 VDD.n3105 VDD.n1256 185
R1488 VDD.n1256 VDD.n1253 185
R1489 VDD.n3104 VDD.n3103 185
R1490 VDD.n3103 VDD.n3102 185
R1491 VDD.n1258 VDD.n1257 185
R1492 VDD.n1259 VDD.n1258 185
R1493 VDD.n3095 VDD.n3094 185
R1494 VDD.n3096 VDD.n3095 185
R1495 VDD.n3093 VDD.n1268 185
R1496 VDD.n1268 VDD.n1265 185
R1497 VDD.n3092 VDD.n3091 185
R1498 VDD.n3091 VDD.n3090 185
R1499 VDD.n1270 VDD.n1269 185
R1500 VDD.n1271 VDD.n1270 185
R1501 VDD.n3083 VDD.n3082 185
R1502 VDD.n3084 VDD.n3083 185
R1503 VDD.n3081 VDD.n1280 185
R1504 VDD.n1280 VDD.n1277 185
R1505 VDD.n3080 VDD.n3079 185
R1506 VDD.n3079 VDD.n3078 185
R1507 VDD.n1282 VDD.n1281 185
R1508 VDD.n1291 VDD.n1282 185
R1509 VDD.n3071 VDD.n3070 185
R1510 VDD.n3072 VDD.n3071 185
R1511 VDD.n3069 VDD.n1292 185
R1512 VDD.n1292 VDD.n1288 185
R1513 VDD.n3068 VDD.n3067 185
R1514 VDD.n3067 VDD.n3066 185
R1515 VDD.n1294 VDD.n1293 185
R1516 VDD.n1295 VDD.n1294 185
R1517 VDD.n3059 VDD.n3058 185
R1518 VDD.n3060 VDD.n3059 185
R1519 VDD.n3057 VDD.n1304 185
R1520 VDD.n1304 VDD.n1301 185
R1521 VDD.n3056 VDD.n3055 185
R1522 VDD.n3055 VDD.n3054 185
R1523 VDD.n1306 VDD.n1305 185
R1524 VDD.n1307 VDD.n1306 185
R1525 VDD.n3047 VDD.n3046 185
R1526 VDD.n3048 VDD.n3047 185
R1527 VDD.n3045 VDD.n1316 185
R1528 VDD.n1316 VDD.n1313 185
R1529 VDD.n3044 VDD.n3043 185
R1530 VDD.n3043 VDD.n3042 185
R1531 VDD.n1318 VDD.n1317 185
R1532 VDD.n1319 VDD.n1318 185
R1533 VDD.n3035 VDD.n3034 185
R1534 VDD.n3036 VDD.n3035 185
R1535 VDD.n3033 VDD.n1328 185
R1536 VDD.n1328 VDD.n1325 185
R1537 VDD.n3032 VDD.n3031 185
R1538 VDD.n3031 VDD.n3030 185
R1539 VDD.n1330 VDD.n1329 185
R1540 VDD.n1331 VDD.n1330 185
R1541 VDD.n3023 VDD.n3022 185
R1542 VDD.n3024 VDD.n3023 185
R1543 VDD.n3021 VDD.n1340 185
R1544 VDD.n1340 VDD.n1337 185
R1545 VDD.n3020 VDD.n3019 185
R1546 VDD.n3019 VDD.n3018 185
R1547 VDD.n1342 VDD.n1341 185
R1548 VDD.n1343 VDD.n1342 185
R1549 VDD.n3011 VDD.n3010 185
R1550 VDD.n3012 VDD.n3011 185
R1551 VDD.n3009 VDD.n1352 185
R1552 VDD.n1352 VDD.n1349 185
R1553 VDD.n3008 VDD.n3007 185
R1554 VDD.n3007 VDD.n3006 185
R1555 VDD.n1354 VDD.n1353 185
R1556 VDD.n1355 VDD.n1354 185
R1557 VDD.n2999 VDD.n2998 185
R1558 VDD.n3000 VDD.n2999 185
R1559 VDD.n2997 VDD.n1363 185
R1560 VDD.n1369 VDD.n1363 185
R1561 VDD.n2996 VDD.n2995 185
R1562 VDD.n2995 VDD.n2994 185
R1563 VDD.n1365 VDD.n1364 185
R1564 VDD.n1366 VDD.n1365 185
R1565 VDD.n2987 VDD.n2986 185
R1566 VDD.n2988 VDD.n2987 185
R1567 VDD.n2985 VDD.n1376 185
R1568 VDD.n1376 VDD.n1373 185
R1569 VDD.n2984 VDD.n2983 185
R1570 VDD.n2983 VDD.n2982 185
R1571 VDD.n1378 VDD.n1377 185
R1572 VDD.n1379 VDD.n1378 185
R1573 VDD.n2975 VDD.n2974 185
R1574 VDD.n2976 VDD.n2975 185
R1575 VDD.n2973 VDD.n1388 185
R1576 VDD.n1388 VDD.n1385 185
R1577 VDD.n2972 VDD.n2971 185
R1578 VDD.n2971 VDD.n2970 185
R1579 VDD.n1390 VDD.n1389 185
R1580 VDD.n1391 VDD.n1390 185
R1581 VDD.n2963 VDD.n2962 185
R1582 VDD.n2964 VDD.n2963 185
R1583 VDD.n2961 VDD.n1400 185
R1584 VDD.n2960 VDD.n2959 185
R1585 VDD.n2957 VDD.n1401 185
R1586 VDD.n2957 VDD.n1397 185
R1587 VDD.n2956 VDD.n2955 185
R1588 VDD.n2954 VDD.n2953 185
R1589 VDD.n2952 VDD.n1403 185
R1590 VDD.n2950 VDD.n2949 185
R1591 VDD.n2948 VDD.n1404 185
R1592 VDD.n2947 VDD.n2946 185
R1593 VDD.n2944 VDD.n1405 185
R1594 VDD.n2942 VDD.n2941 185
R1595 VDD.n1594 VDD.n1406 185
R1596 VDD.n1593 VDD.n1592 185
R1597 VDD.n1590 VDD.n1407 185
R1598 VDD.n1588 VDD.n1587 185
R1599 VDD.n1586 VDD.n1408 185
R1600 VDD.n1585 VDD.n1584 185
R1601 VDD.n1582 VDD.n1581 185
R1602 VDD.n1580 VDD.n1579 185
R1603 VDD.n1578 VDD.n1413 185
R1604 VDD.n1576 VDD.n1575 185
R1605 VDD.n3345 VDD.n3344 185
R1606 VDD.n3347 VDD.n3346 185
R1607 VDD.n3349 VDD.n3348 185
R1608 VDD.n3351 VDD.n3350 185
R1609 VDD.n3353 VDD.n3352 185
R1610 VDD.n3355 VDD.n3354 185
R1611 VDD.n3357 VDD.n3356 185
R1612 VDD.n3359 VDD.n3358 185
R1613 VDD.n3361 VDD.n3360 185
R1614 VDD.n3363 VDD.n3362 185
R1615 VDD.n3365 VDD.n3364 185
R1616 VDD.n3367 VDD.n3366 185
R1617 VDD.n3369 VDD.n3368 185
R1618 VDD.n3371 VDD.n3370 185
R1619 VDD.n3373 VDD.n3372 185
R1620 VDD.n3375 VDD.n3374 185
R1621 VDD.n3377 VDD.n3376 185
R1622 VDD.n3379 VDD.n3378 185
R1623 VDD.n3381 VDD.n3380 185
R1624 VDD.n3382 VDD.n1059 185
R1625 VDD.n3384 VDD.n3383 185
R1626 VDD.n3385 VDD.n3384 185
R1627 VDD.n3343 VDD.n1064 185
R1628 VDD.n3343 VDD.n1036 185
R1629 VDD.n3342 VDD.n1066 185
R1630 VDD.n3342 VDD.n3341 185
R1631 VDD.n1414 VDD.n1065 185
R1632 VDD.n1067 VDD.n1065 185
R1633 VDD.n1415 VDD.n1074 185
R1634 VDD.n3335 VDD.n1074 185
R1635 VDD.n1417 VDD.n1416 185
R1636 VDD.n1416 VDD.n1073 185
R1637 VDD.n1418 VDD.n1085 185
R1638 VDD.n3278 VDD.n1085 185
R1639 VDD.n1420 VDD.n1419 185
R1640 VDD.n1419 VDD.n1084 185
R1641 VDD.n1421 VDD.n1091 185
R1642 VDD.n3272 VDD.n1091 185
R1643 VDD.n1423 VDD.n1422 185
R1644 VDD.n1422 VDD.n1090 185
R1645 VDD.n1424 VDD.n1098 185
R1646 VDD.n3264 VDD.n1098 185
R1647 VDD.n1426 VDD.n1425 185
R1648 VDD.n1425 VDD.n1097 185
R1649 VDD.n1427 VDD.n1103 185
R1650 VDD.n3258 VDD.n1103 185
R1651 VDD.n1429 VDD.n1428 185
R1652 VDD.n1428 VDD.n1110 185
R1653 VDD.n1430 VDD.n1108 185
R1654 VDD.n3252 VDD.n1108 185
R1655 VDD.n1432 VDD.n1431 185
R1656 VDD.n1431 VDD.n1117 185
R1657 VDD.n1433 VDD.n1115 185
R1658 VDD.n3246 VDD.n1115 185
R1659 VDD.n1435 VDD.n1434 185
R1660 VDD.n1434 VDD.n1114 185
R1661 VDD.n1436 VDD.n1122 185
R1662 VDD.n3240 VDD.n1122 185
R1663 VDD.n1438 VDD.n1437 185
R1664 VDD.n1437 VDD.n1121 185
R1665 VDD.n1439 VDD.n1128 185
R1666 VDD.n3234 VDD.n1128 185
R1667 VDD.n1441 VDD.n1440 185
R1668 VDD.n1440 VDD.n1127 185
R1669 VDD.n1442 VDD.n1134 185
R1670 VDD.n3228 VDD.n1134 185
R1671 VDD.n1444 VDD.n1443 185
R1672 VDD.n1443 VDD.n1133 185
R1673 VDD.n1445 VDD.n1140 185
R1674 VDD.n3222 VDD.n1140 185
R1675 VDD.n1447 VDD.n1446 185
R1676 VDD.n1446 VDD.n1139 185
R1677 VDD.n1448 VDD.n1146 185
R1678 VDD.n3216 VDD.n1146 185
R1679 VDD.n1450 VDD.n1449 185
R1680 VDD.n1449 VDD.n1145 185
R1681 VDD.n1451 VDD.n1152 185
R1682 VDD.n3210 VDD.n1152 185
R1683 VDD.n1453 VDD.n1452 185
R1684 VDD.n1452 VDD.n1151 185
R1685 VDD.n1454 VDD.n1158 185
R1686 VDD.n3204 VDD.n1158 185
R1687 VDD.n1456 VDD.n1455 185
R1688 VDD.n1455 VDD.n1157 185
R1689 VDD.n1457 VDD.n1164 185
R1690 VDD.n3198 VDD.n1164 185
R1691 VDD.n1459 VDD.n1458 185
R1692 VDD.n1458 VDD.n1163 185
R1693 VDD.n1460 VDD.n1170 185
R1694 VDD.n3192 VDD.n1170 185
R1695 VDD.n1462 VDD.n1461 185
R1696 VDD.n1461 VDD.n1169 185
R1697 VDD.n1463 VDD.n1176 185
R1698 VDD.n3186 VDD.n1176 185
R1699 VDD.n1465 VDD.n1464 185
R1700 VDD.n1464 VDD.n1175 185
R1701 VDD.n1466 VDD.n1182 185
R1702 VDD.n3180 VDD.n1182 185
R1703 VDD.n1468 VDD.n1467 185
R1704 VDD.n1467 VDD.n1181 185
R1705 VDD.n1469 VDD.n1188 185
R1706 VDD.n3174 VDD.n1188 185
R1707 VDD.n1471 VDD.n1470 185
R1708 VDD.n1470 VDD.n1187 185
R1709 VDD.n1472 VDD.n1194 185
R1710 VDD.n3168 VDD.n1194 185
R1711 VDD.n1474 VDD.n1473 185
R1712 VDD.n1473 VDD.n1193 185
R1713 VDD.n1475 VDD.n1200 185
R1714 VDD.n3162 VDD.n1200 185
R1715 VDD.n1477 VDD.n1476 185
R1716 VDD.n1476 VDD.n1199 185
R1717 VDD.n1478 VDD.n1206 185
R1718 VDD.n3156 VDD.n1206 185
R1719 VDD.n1480 VDD.n1479 185
R1720 VDD.n1479 VDD.n1205 185
R1721 VDD.n1481 VDD.n1212 185
R1722 VDD.n3150 VDD.n1212 185
R1723 VDD.n1483 VDD.n1482 185
R1724 VDD.n1482 VDD.n1211 185
R1725 VDD.n1484 VDD.n1218 185
R1726 VDD.n3144 VDD.n1218 185
R1727 VDD.n1486 VDD.n1485 185
R1728 VDD.n1485 VDD.n1217 185
R1729 VDD.n1487 VDD.n1224 185
R1730 VDD.n3138 VDD.n1224 185
R1731 VDD.n1489 VDD.n1488 185
R1732 VDD.n1488 VDD.n1223 185
R1733 VDD.n1490 VDD.n1230 185
R1734 VDD.n3132 VDD.n1230 185
R1735 VDD.n1492 VDD.n1491 185
R1736 VDD.n1491 VDD.n1229 185
R1737 VDD.n1493 VDD.n1236 185
R1738 VDD.n3126 VDD.n1236 185
R1739 VDD.n1495 VDD.n1494 185
R1740 VDD.n1494 VDD.n1235 185
R1741 VDD.n1496 VDD.n1242 185
R1742 VDD.n3120 VDD.n1242 185
R1743 VDD.n1498 VDD.n1497 185
R1744 VDD.n1497 VDD.n1241 185
R1745 VDD.n1499 VDD.n1248 185
R1746 VDD.n3114 VDD.n1248 185
R1747 VDD.n1501 VDD.n1500 185
R1748 VDD.n1500 VDD.n1247 185
R1749 VDD.n1502 VDD.n1254 185
R1750 VDD.n3108 VDD.n1254 185
R1751 VDD.n1504 VDD.n1503 185
R1752 VDD.n1503 VDD.n1253 185
R1753 VDD.n1505 VDD.n1260 185
R1754 VDD.n3102 VDD.n1260 185
R1755 VDD.n1507 VDD.n1506 185
R1756 VDD.n1506 VDD.n1259 185
R1757 VDD.n1508 VDD.n1266 185
R1758 VDD.n3096 VDD.n1266 185
R1759 VDD.n1510 VDD.n1509 185
R1760 VDD.n1509 VDD.n1265 185
R1761 VDD.n1511 VDD.n1272 185
R1762 VDD.n3090 VDD.n1272 185
R1763 VDD.n1513 VDD.n1512 185
R1764 VDD.n1512 VDD.n1271 185
R1765 VDD.n1514 VDD.n1278 185
R1766 VDD.n3084 VDD.n1278 185
R1767 VDD.n1516 VDD.n1515 185
R1768 VDD.n1515 VDD.n1277 185
R1769 VDD.n1517 VDD.n1283 185
R1770 VDD.n3078 VDD.n1283 185
R1771 VDD.n1519 VDD.n1518 185
R1772 VDD.n1518 VDD.n1291 185
R1773 VDD.n1520 VDD.n1289 185
R1774 VDD.n3072 VDD.n1289 185
R1775 VDD.n1522 VDD.n1521 185
R1776 VDD.n1521 VDD.n1288 185
R1777 VDD.n1523 VDD.n1296 185
R1778 VDD.n3066 VDD.n1296 185
R1779 VDD.n1525 VDD.n1524 185
R1780 VDD.n1524 VDD.n1295 185
R1781 VDD.n1526 VDD.n1302 185
R1782 VDD.n3060 VDD.n1302 185
R1783 VDD.n1528 VDD.n1527 185
R1784 VDD.n1527 VDD.n1301 185
R1785 VDD.n1529 VDD.n1308 185
R1786 VDD.n3054 VDD.n1308 185
R1787 VDD.n1531 VDD.n1530 185
R1788 VDD.n1530 VDD.n1307 185
R1789 VDD.n1532 VDD.n1314 185
R1790 VDD.n3048 VDD.n1314 185
R1791 VDD.n1534 VDD.n1533 185
R1792 VDD.n1533 VDD.n1313 185
R1793 VDD.n1535 VDD.n1320 185
R1794 VDD.n3042 VDD.n1320 185
R1795 VDD.n1537 VDD.n1536 185
R1796 VDD.n1536 VDD.n1319 185
R1797 VDD.n1538 VDD.n1326 185
R1798 VDD.n3036 VDD.n1326 185
R1799 VDD.n1540 VDD.n1539 185
R1800 VDD.n1539 VDD.n1325 185
R1801 VDD.n1541 VDD.n1332 185
R1802 VDD.n3030 VDD.n1332 185
R1803 VDD.n1543 VDD.n1542 185
R1804 VDD.n1542 VDD.n1331 185
R1805 VDD.n1544 VDD.n1338 185
R1806 VDD.n3024 VDD.n1338 185
R1807 VDD.n1546 VDD.n1545 185
R1808 VDD.n1545 VDD.n1337 185
R1809 VDD.n1547 VDD.n1344 185
R1810 VDD.n3018 VDD.n1344 185
R1811 VDD.n1549 VDD.n1548 185
R1812 VDD.n1548 VDD.n1343 185
R1813 VDD.n1550 VDD.n1350 185
R1814 VDD.n3012 VDD.n1350 185
R1815 VDD.n1552 VDD.n1551 185
R1816 VDD.n1551 VDD.n1349 185
R1817 VDD.n1553 VDD.n1356 185
R1818 VDD.n3006 VDD.n1356 185
R1819 VDD.n1555 VDD.n1554 185
R1820 VDD.n1554 VDD.n1355 185
R1821 VDD.n1556 VDD.n1361 185
R1822 VDD.n3000 VDD.n1361 185
R1823 VDD.n1558 VDD.n1557 185
R1824 VDD.n1557 VDD.n1369 185
R1825 VDD.n1559 VDD.n1367 185
R1826 VDD.n2994 VDD.n1367 185
R1827 VDD.n1561 VDD.n1560 185
R1828 VDD.n1560 VDD.n1366 185
R1829 VDD.n1562 VDD.n1374 185
R1830 VDD.n2988 VDD.n1374 185
R1831 VDD.n1564 VDD.n1563 185
R1832 VDD.n1563 VDD.n1373 185
R1833 VDD.n1565 VDD.n1380 185
R1834 VDD.n2982 VDD.n1380 185
R1835 VDD.n1567 VDD.n1566 185
R1836 VDD.n1566 VDD.n1379 185
R1837 VDD.n1568 VDD.n1386 185
R1838 VDD.n2976 VDD.n1386 185
R1839 VDD.n1570 VDD.n1569 185
R1840 VDD.n1569 VDD.n1385 185
R1841 VDD.n1571 VDD.n1392 185
R1842 VDD.n2970 VDD.n1392 185
R1843 VDD.n1573 VDD.n1572 185
R1844 VDD.n1572 VDD.n1391 185
R1845 VDD.n1574 VDD.n1398 185
R1846 VDD.n2964 VDD.n1398 185
R1847 VDD.n196 VDD.n195 185
R1848 VDD.n4594 VDD.n196 185
R1849 VDD.n4597 VDD.n4596 185
R1850 VDD.n4596 VDD.n4595 185
R1851 VDD.n4598 VDD.n190 185
R1852 VDD.n190 VDD.n189 185
R1853 VDD.n4600 VDD.n4599 185
R1854 VDD.n4601 VDD.n4600 185
R1855 VDD.n184 VDD.n183 185
R1856 VDD.n4602 VDD.n184 185
R1857 VDD.n4605 VDD.n4604 185
R1858 VDD.n4604 VDD.n4603 185
R1859 VDD.n4606 VDD.n178 185
R1860 VDD.n185 VDD.n178 185
R1861 VDD.n4608 VDD.n4607 185
R1862 VDD.n4609 VDD.n4608 185
R1863 VDD.n174 VDD.n173 185
R1864 VDD.n4610 VDD.n174 185
R1865 VDD.n4613 VDD.n4612 185
R1866 VDD.n4612 VDD.n4611 185
R1867 VDD.n4614 VDD.n168 185
R1868 VDD.n168 VDD.n167 185
R1869 VDD.n4616 VDD.n4615 185
R1870 VDD.n4617 VDD.n4616 185
R1871 VDD.n163 VDD.n162 185
R1872 VDD.n4618 VDD.n163 185
R1873 VDD.n4621 VDD.n4620 185
R1874 VDD.n4620 VDD.n4619 185
R1875 VDD.n4622 VDD.n157 185
R1876 VDD.n157 VDD.n156 185
R1877 VDD.n4624 VDD.n4623 185
R1878 VDD.n4625 VDD.n4624 185
R1879 VDD.n152 VDD.n151 185
R1880 VDD.n4626 VDD.n152 185
R1881 VDD.n4629 VDD.n4628 185
R1882 VDD.n4628 VDD.n4627 185
R1883 VDD.n4630 VDD.n146 185
R1884 VDD.n146 VDD.n145 185
R1885 VDD.n4632 VDD.n4631 185
R1886 VDD.n4633 VDD.n4632 185
R1887 VDD.n141 VDD.n140 185
R1888 VDD.n4634 VDD.n141 185
R1889 VDD.n4637 VDD.n4636 185
R1890 VDD.n4636 VDD.n4635 185
R1891 VDD.n4638 VDD.n135 185
R1892 VDD.n135 VDD.n134 185
R1893 VDD.n4640 VDD.n4639 185
R1894 VDD.n4641 VDD.n4640 185
R1895 VDD.n130 VDD.n129 185
R1896 VDD.n4642 VDD.n130 185
R1897 VDD.n4645 VDD.n4644 185
R1898 VDD.n4644 VDD.n4643 185
R1899 VDD.n4646 VDD.n124 185
R1900 VDD.n124 VDD.n123 185
R1901 VDD.n4648 VDD.n4647 185
R1902 VDD.n4649 VDD.n4648 185
R1903 VDD.n119 VDD.n118 185
R1904 VDD.n4650 VDD.n119 185
R1905 VDD.n4653 VDD.n4652 185
R1906 VDD.n4652 VDD.n4651 185
R1907 VDD.n4654 VDD.n113 185
R1908 VDD.n113 VDD.n112 185
R1909 VDD.n4656 VDD.n4655 185
R1910 VDD.n4657 VDD.n4656 185
R1911 VDD.n108 VDD.n107 185
R1912 VDD.n4658 VDD.n108 185
R1913 VDD.n4661 VDD.n4660 185
R1914 VDD.n4660 VDD.n4659 185
R1915 VDD.n4662 VDD.n102 185
R1916 VDD.n102 VDD.n101 185
R1917 VDD.n4664 VDD.n4663 185
R1918 VDD.n4665 VDD.n4664 185
R1919 VDD.n97 VDD.n96 185
R1920 VDD.n4666 VDD.n97 185
R1921 VDD.n4669 VDD.n4668 185
R1922 VDD.n4668 VDD.n4667 185
R1923 VDD.n4670 VDD.n91 185
R1924 VDD.n91 VDD.n90 185
R1925 VDD.n4672 VDD.n4671 185
R1926 VDD.n4673 VDD.n4672 185
R1927 VDD.n86 VDD.n85 185
R1928 VDD.n4674 VDD.n86 185
R1929 VDD.n4677 VDD.n4676 185
R1930 VDD.n4676 VDD.n4675 185
R1931 VDD.n4678 VDD.n80 185
R1932 VDD.n80 VDD.n79 185
R1933 VDD.n4680 VDD.n4679 185
R1934 VDD.n4681 VDD.n4680 185
R1935 VDD.n74 VDD.n73 185
R1936 VDD.n4682 VDD.n74 185
R1937 VDD.n4685 VDD.n4684 185
R1938 VDD.n4684 VDD.n4683 185
R1939 VDD.n4686 VDD.n68 185
R1940 VDD.n75 VDD.n68 185
R1941 VDD.n4688 VDD.n4687 185
R1942 VDD.n4689 VDD.n4688 185
R1943 VDD.n64 VDD.n63 185
R1944 VDD.n4690 VDD.n64 185
R1945 VDD.n4693 VDD.n4692 185
R1946 VDD.n4692 VDD.n4691 185
R1947 VDD.n4694 VDD.n58 185
R1948 VDD.n58 VDD.n57 185
R1949 VDD.n4696 VDD.n4695 185
R1950 VDD.n4697 VDD.n4696 185
R1951 VDD.n53 VDD.n52 185
R1952 VDD.n4698 VDD.n53 185
R1953 VDD.n4701 VDD.n4700 185
R1954 VDD.n4700 VDD.n4699 185
R1955 VDD.n4702 VDD.n47 185
R1956 VDD.n47 VDD.n46 185
R1957 VDD.n4704 VDD.n4703 185
R1958 VDD.n4705 VDD.n4704 185
R1959 VDD.n41 VDD.n40 185
R1960 VDD.n4706 VDD.n41 185
R1961 VDD.n4709 VDD.n4708 185
R1962 VDD.n4708 VDD.n4707 185
R1963 VDD.n4710 VDD.n39 185
R1964 VDD.n42 VDD.n39 185
R1965 VDD.n4483 VDD.n38 185
R1966 VDD.n4484 VDD.n4483 185
R1967 VDD.n4482 VDD.n4481 185
R1968 VDD.n4482 VDD.n370 185
R1969 VDD.n372 VDD.n371 185
R1970 VDD.n4474 VDD.n371 185
R1971 VDD.n4477 VDD.n4476 185
R1972 VDD.n4476 VDD.n4475 185
R1973 VDD.n375 VDD.n374 185
R1974 VDD.n376 VDD.n375 185
R1975 VDD.n4461 VDD.n4460 185
R1976 VDD.n4462 VDD.n4461 185
R1977 VDD.n384 VDD.n383 185
R1978 VDD.n383 VDD.n382 185
R1979 VDD.n4456 VDD.n4455 185
R1980 VDD.n4455 VDD.n4454 185
R1981 VDD.n387 VDD.n386 185
R1982 VDD.n388 VDD.n387 185
R1983 VDD.n4443 VDD.n4442 185
R1984 VDD.n4444 VDD.n4443 185
R1985 VDD.n396 VDD.n395 185
R1986 VDD.n395 VDD.n394 185
R1987 VDD.n4438 VDD.n4437 185
R1988 VDD.n4437 VDD.n4436 185
R1989 VDD.n399 VDD.n398 185
R1990 VDD.n406 VDD.n399 185
R1991 VDD.n4427 VDD.n4426 185
R1992 VDD.n4428 VDD.n4427 185
R1993 VDD.n408 VDD.n407 185
R1994 VDD.n407 VDD.n405 185
R1995 VDD.n4422 VDD.n4421 185
R1996 VDD.n4421 VDD.n4420 185
R1997 VDD.n411 VDD.n410 185
R1998 VDD.n412 VDD.n411 185
R1999 VDD.n4411 VDD.n4410 185
R2000 VDD.n4412 VDD.n4411 185
R2001 VDD.n420 VDD.n419 185
R2002 VDD.n419 VDD.n418 185
R2003 VDD.n4406 VDD.n4405 185
R2004 VDD.n4405 VDD.n4404 185
R2005 VDD.n423 VDD.n422 185
R2006 VDD.n424 VDD.n423 185
R2007 VDD.n4395 VDD.n4394 185
R2008 VDD.n4396 VDD.n4395 185
R2009 VDD.n432 VDD.n431 185
R2010 VDD.n431 VDD.n430 185
R2011 VDD.n4390 VDD.n4389 185
R2012 VDD.n4389 VDD.n4388 185
R2013 VDD.n435 VDD.n434 185
R2014 VDD.n436 VDD.n435 185
R2015 VDD.n4379 VDD.n4378 185
R2016 VDD.n4380 VDD.n4379 185
R2017 VDD.n444 VDD.n443 185
R2018 VDD.n443 VDD.n442 185
R2019 VDD.n4374 VDD.n4373 185
R2020 VDD.n4373 VDD.n4372 185
R2021 VDD.n447 VDD.n446 185
R2022 VDD.n448 VDD.n447 185
R2023 VDD.n4363 VDD.n4362 185
R2024 VDD.n4364 VDD.n4363 185
R2025 VDD.n456 VDD.n455 185
R2026 VDD.n455 VDD.n454 185
R2027 VDD.n4358 VDD.n4357 185
R2028 VDD.n4357 VDD.n4356 185
R2029 VDD.n459 VDD.n458 185
R2030 VDD.n460 VDD.n459 185
R2031 VDD.n4347 VDD.n4346 185
R2032 VDD.n4348 VDD.n4347 185
R2033 VDD.n468 VDD.n467 185
R2034 VDD.n467 VDD.n466 185
R2035 VDD.n4342 VDD.n4341 185
R2036 VDD.n4341 VDD.n4340 185
R2037 VDD.n471 VDD.n470 185
R2038 VDD.n472 VDD.n471 185
R2039 VDD.n4331 VDD.n4330 185
R2040 VDD.n4332 VDD.n4331 185
R2041 VDD.n480 VDD.n479 185
R2042 VDD.n479 VDD.n478 185
R2043 VDD.n4326 VDD.n4325 185
R2044 VDD.n4325 VDD.n4324 185
R2045 VDD.n483 VDD.n482 185
R2046 VDD.n484 VDD.n483 185
R2047 VDD.n4315 VDD.n4314 185
R2048 VDD.n4316 VDD.n4315 185
R2049 VDD.n492 VDD.n491 185
R2050 VDD.n491 VDD.n490 185
R2051 VDD.n4310 VDD.n4309 185
R2052 VDD.n4309 VDD.n4308 185
R2053 VDD.n495 VDD.n494 185
R2054 VDD.n496 VDD.n495 185
R2055 VDD.n4299 VDD.n4298 185
R2056 VDD.n4300 VDD.n4299 185
R2057 VDD.n504 VDD.n503 185
R2058 VDD.n503 VDD.n502 185
R2059 VDD.n4294 VDD.n4293 185
R2060 VDD.n4293 VDD.n4292 185
R2061 VDD.n507 VDD.n506 185
R2062 VDD.n508 VDD.n507 185
R2063 VDD.n4283 VDD.n4282 185
R2064 VDD.n4284 VDD.n4283 185
R2065 VDD.n516 VDD.n515 185
R2066 VDD.n515 VDD.n514 185
R2067 VDD.n4278 VDD.n4277 185
R2068 VDD.n4277 VDD.n4276 185
R2069 VDD.n519 VDD.n518 185
R2070 VDD.n526 VDD.n519 185
R2071 VDD.n4267 VDD.n4266 185
R2072 VDD.n4268 VDD.n4267 185
R2073 VDD.n528 VDD.n527 185
R2074 VDD.n527 VDD.n525 185
R2075 VDD.n4262 VDD.n4261 185
R2076 VDD.n4261 VDD.n4260 185
R2077 VDD.n531 VDD.n530 185
R2078 VDD.n532 VDD.n531 185
R2079 VDD.n4251 VDD.n4250 185
R2080 VDD.n4252 VDD.n4251 185
R2081 VDD.n540 VDD.n539 185
R2082 VDD.n539 VDD.n538 185
R2083 VDD.n4246 VDD.n543 185
R2084 VDD.n4245 VDD.n4244 185
R2085 VDD.n546 VDD.n545 185
R2086 VDD.n4242 VDD.n546 185
R2087 VDD.n592 VDD.n591 185
R2088 VDD.n595 VDD.n594 185
R2089 VDD.n593 VDD.n588 185
R2090 VDD.n600 VDD.n599 185
R2091 VDD.n602 VDD.n601 185
R2092 VDD.n605 VDD.n604 185
R2093 VDD.n603 VDD.n586 185
R2094 VDD.n610 VDD.n609 185
R2095 VDD.n612 VDD.n611 185
R2096 VDD.n615 VDD.n614 185
R2097 VDD.n613 VDD.n581 185
R2098 VDD.n620 VDD.n619 185
R2099 VDD.n622 VDD.n621 185
R2100 VDD.n625 VDD.n624 185
R2101 VDD.n623 VDD.n579 185
R2102 VDD.n630 VDD.n629 185
R2103 VDD.n632 VDD.n631 185
R2104 VDD.n635 VDD.n634 185
R2105 VDD.n633 VDD.n577 185
R2106 VDD.n640 VDD.n639 185
R2107 VDD.n642 VDD.n641 185
R2108 VDD.n646 VDD.n645 185
R2109 VDD.n644 VDD.n573 185
R2110 VDD.n651 VDD.n650 185
R2111 VDD.n653 VDD.n652 185
R2112 VDD.n656 VDD.n655 185
R2113 VDD.n654 VDD.n571 185
R2114 VDD.n661 VDD.n660 185
R2115 VDD.n663 VDD.n662 185
R2116 VDD.n666 VDD.n665 185
R2117 VDD.n664 VDD.n569 185
R2118 VDD.n671 VDD.n670 185
R2119 VDD.n673 VDD.n672 185
R2120 VDD.n674 VDD.n564 185
R2121 VDD.n4241 VDD.n4240 185
R2122 VDD.n4242 VDD.n4241 185
R2123 VDD.n4591 VDD.n4590 185
R2124 VDD.n336 VDD.n217 185
R2125 VDD.n335 VDD.n334 185
R2126 VDD.n333 VDD.n332 185
R2127 VDD.n331 VDD.n222 185
R2128 VDD.n327 VDD.n326 185
R2129 VDD.n325 VDD.n324 185
R2130 VDD.n323 VDD.n322 185
R2131 VDD.n321 VDD.n224 185
R2132 VDD.n317 VDD.n316 185
R2133 VDD.n315 VDD.n314 185
R2134 VDD.n313 VDD.n312 185
R2135 VDD.n311 VDD.n226 185
R2136 VDD.n307 VDD.n306 185
R2137 VDD.n305 VDD.n304 185
R2138 VDD.n303 VDD.n302 185
R2139 VDD.n301 VDD.n231 185
R2140 VDD.n297 VDD.n296 185
R2141 VDD.n295 VDD.n294 185
R2142 VDD.n293 VDD.n292 185
R2143 VDD.n291 VDD.n233 185
R2144 VDD.n287 VDD.n286 185
R2145 VDD.n285 VDD.n284 185
R2146 VDD.n283 VDD.n282 185
R2147 VDD.n281 VDD.n235 185
R2148 VDD.n277 VDD.n276 185
R2149 VDD.n275 VDD.n274 185
R2150 VDD.n272 VDD.n271 185
R2151 VDD.n270 VDD.n239 185
R2152 VDD.n266 VDD.n265 185
R2153 VDD.n264 VDD.n263 185
R2154 VDD.n262 VDD.n261 185
R2155 VDD.n260 VDD.n241 185
R2156 VDD.n256 VDD.n255 185
R2157 VDD.n254 VDD.n253 185
R2158 VDD.n252 VDD.n251 185
R2159 VDD.n250 VDD.n243 185
R2160 VDD.n246 VDD.n245 185
R2161 VDD.n4587 VDD.n198 185
R2162 VDD.n4594 VDD.n198 185
R2163 VDD.n4586 VDD.n197 185
R2164 VDD.n4595 VDD.n197 185
R2165 VDD.n4585 VDD.n4584 185
R2166 VDD.n4584 VDD.n189 185
R2167 VDD.n339 VDD.n188 185
R2168 VDD.n4601 VDD.n188 185
R2169 VDD.n4580 VDD.n187 185
R2170 VDD.n4602 VDD.n187 185
R2171 VDD.n4579 VDD.n186 185
R2172 VDD.n4603 VDD.n186 185
R2173 VDD.n4578 VDD.n4577 185
R2174 VDD.n4577 VDD.n185 185
R2175 VDD.n341 VDD.n177 185
R2176 VDD.n4609 VDD.n177 185
R2177 VDD.n4573 VDD.n176 185
R2178 VDD.n4610 VDD.n176 185
R2179 VDD.n4572 VDD.n175 185
R2180 VDD.n4611 VDD.n175 185
R2181 VDD.n4571 VDD.n4570 185
R2182 VDD.n4570 VDD.n167 185
R2183 VDD.n343 VDD.n166 185
R2184 VDD.n4617 VDD.n166 185
R2185 VDD.n4566 VDD.n165 185
R2186 VDD.n4618 VDD.n165 185
R2187 VDD.n4565 VDD.n164 185
R2188 VDD.n4619 VDD.n164 185
R2189 VDD.n4564 VDD.n4563 185
R2190 VDD.n4563 VDD.n156 185
R2191 VDD.n345 VDD.n155 185
R2192 VDD.n4625 VDD.n155 185
R2193 VDD.n4559 VDD.n154 185
R2194 VDD.n4626 VDD.n154 185
R2195 VDD.n4558 VDD.n153 185
R2196 VDD.n4627 VDD.n153 185
R2197 VDD.n4557 VDD.n4556 185
R2198 VDD.n4556 VDD.n145 185
R2199 VDD.n347 VDD.n144 185
R2200 VDD.n4633 VDD.n144 185
R2201 VDD.n4552 VDD.n143 185
R2202 VDD.n4634 VDD.n143 185
R2203 VDD.n4551 VDD.n142 185
R2204 VDD.n4635 VDD.n142 185
R2205 VDD.n4550 VDD.n4549 185
R2206 VDD.n4549 VDD.n134 185
R2207 VDD.n349 VDD.n133 185
R2208 VDD.n4641 VDD.n133 185
R2209 VDD.n4545 VDD.n132 185
R2210 VDD.n4642 VDD.n132 185
R2211 VDD.n4544 VDD.n131 185
R2212 VDD.n4643 VDD.n131 185
R2213 VDD.n4543 VDD.n4542 185
R2214 VDD.n4542 VDD.n123 185
R2215 VDD.n351 VDD.n122 185
R2216 VDD.n4649 VDD.n122 185
R2217 VDD.n4538 VDD.n121 185
R2218 VDD.n4650 VDD.n121 185
R2219 VDD.n4537 VDD.n120 185
R2220 VDD.n4651 VDD.n120 185
R2221 VDD.n4536 VDD.n4535 185
R2222 VDD.n4535 VDD.n112 185
R2223 VDD.n353 VDD.n111 185
R2224 VDD.n4657 VDD.n111 185
R2225 VDD.n4531 VDD.n110 185
R2226 VDD.n4658 VDD.n110 185
R2227 VDD.n4530 VDD.n109 185
R2228 VDD.n4659 VDD.n109 185
R2229 VDD.n4529 VDD.n4528 185
R2230 VDD.n4528 VDD.n101 185
R2231 VDD.n355 VDD.n100 185
R2232 VDD.n4665 VDD.n100 185
R2233 VDD.n4524 VDD.n99 185
R2234 VDD.n4666 VDD.n99 185
R2235 VDD.n4523 VDD.n98 185
R2236 VDD.n4667 VDD.n98 185
R2237 VDD.n4522 VDD.n4521 185
R2238 VDD.n4521 VDD.n90 185
R2239 VDD.n357 VDD.n89 185
R2240 VDD.n4673 VDD.n89 185
R2241 VDD.n4517 VDD.n88 185
R2242 VDD.n4674 VDD.n88 185
R2243 VDD.n4516 VDD.n87 185
R2244 VDD.n4675 VDD.n87 185
R2245 VDD.n4515 VDD.n4514 185
R2246 VDD.n4514 VDD.n79 185
R2247 VDD.n359 VDD.n78 185
R2248 VDD.n4681 VDD.n78 185
R2249 VDD.n4510 VDD.n77 185
R2250 VDD.n4682 VDD.n77 185
R2251 VDD.n4509 VDD.n76 185
R2252 VDD.n4683 VDD.n76 185
R2253 VDD.n4508 VDD.n4507 185
R2254 VDD.n4507 VDD.n75 185
R2255 VDD.n361 VDD.n67 185
R2256 VDD.n4689 VDD.n67 185
R2257 VDD.n4503 VDD.n66 185
R2258 VDD.n4690 VDD.n66 185
R2259 VDD.n4502 VDD.n65 185
R2260 VDD.n4691 VDD.n65 185
R2261 VDD.n4501 VDD.n4500 185
R2262 VDD.n4500 VDD.n57 185
R2263 VDD.n363 VDD.n56 185
R2264 VDD.n4697 VDD.n56 185
R2265 VDD.n4496 VDD.n55 185
R2266 VDD.n4698 VDD.n55 185
R2267 VDD.n4495 VDD.n54 185
R2268 VDD.n4699 VDD.n54 185
R2269 VDD.n4494 VDD.n4493 185
R2270 VDD.n4493 VDD.n46 185
R2271 VDD.n365 VDD.n45 185
R2272 VDD.n4705 VDD.n45 185
R2273 VDD.n4489 VDD.n44 185
R2274 VDD.n4706 VDD.n44 185
R2275 VDD.n4488 VDD.n43 185
R2276 VDD.n4707 VDD.n43 185
R2277 VDD.n4487 VDD.n4486 185
R2278 VDD.n4486 VDD.n42 185
R2279 VDD.n4485 VDD.n367 185
R2280 VDD.n4485 VDD.n4484 185
R2281 VDD.n4471 VDD.n369 185
R2282 VDD.n370 VDD.n369 185
R2283 VDD.n4473 VDD.n4472 185
R2284 VDD.n4474 VDD.n4473 185
R2285 VDD.n378 VDD.n377 185
R2286 VDD.n4475 VDD.n377 185
R2287 VDD.n4465 VDD.n4464 185
R2288 VDD.n4464 VDD.n376 185
R2289 VDD.n4463 VDD.n380 185
R2290 VDD.n4463 VDD.n4462 185
R2291 VDD.n4451 VDD.n381 185
R2292 VDD.n382 VDD.n381 185
R2293 VDD.n4453 VDD.n4452 185
R2294 VDD.n4454 VDD.n4453 185
R2295 VDD.n390 VDD.n389 185
R2296 VDD.n389 VDD.n388 185
R2297 VDD.n4446 VDD.n4445 185
R2298 VDD.n4445 VDD.n4444 185
R2299 VDD.n393 VDD.n392 185
R2300 VDD.n394 VDD.n393 185
R2301 VDD.n4435 VDD.n4434 185
R2302 VDD.n4436 VDD.n4435 185
R2303 VDD.n401 VDD.n400 185
R2304 VDD.n406 VDD.n400 185
R2305 VDD.n4430 VDD.n4429 185
R2306 VDD.n4429 VDD.n4428 185
R2307 VDD.n404 VDD.n403 185
R2308 VDD.n405 VDD.n404 185
R2309 VDD.n4419 VDD.n4418 185
R2310 VDD.n4420 VDD.n4419 185
R2311 VDD.n414 VDD.n413 185
R2312 VDD.n413 VDD.n412 185
R2313 VDD.n4414 VDD.n4413 185
R2314 VDD.n4413 VDD.n4412 185
R2315 VDD.n417 VDD.n416 185
R2316 VDD.n418 VDD.n417 185
R2317 VDD.n4403 VDD.n4402 185
R2318 VDD.n4404 VDD.n4403 185
R2319 VDD.n426 VDD.n425 185
R2320 VDD.n425 VDD.n424 185
R2321 VDD.n4398 VDD.n4397 185
R2322 VDD.n4397 VDD.n4396 185
R2323 VDD.n429 VDD.n428 185
R2324 VDD.n430 VDD.n429 185
R2325 VDD.n4387 VDD.n4386 185
R2326 VDD.n4388 VDD.n4387 185
R2327 VDD.n438 VDD.n437 185
R2328 VDD.n437 VDD.n436 185
R2329 VDD.n4382 VDD.n4381 185
R2330 VDD.n4381 VDD.n4380 185
R2331 VDD.n441 VDD.n440 185
R2332 VDD.n442 VDD.n441 185
R2333 VDD.n4371 VDD.n4370 185
R2334 VDD.n4372 VDD.n4371 185
R2335 VDD.n450 VDD.n449 185
R2336 VDD.n449 VDD.n448 185
R2337 VDD.n4366 VDD.n4365 185
R2338 VDD.n4365 VDD.n4364 185
R2339 VDD.n453 VDD.n452 185
R2340 VDD.n454 VDD.n453 185
R2341 VDD.n4355 VDD.n4354 185
R2342 VDD.n4356 VDD.n4355 185
R2343 VDD.n462 VDD.n461 185
R2344 VDD.n461 VDD.n460 185
R2345 VDD.n4350 VDD.n4349 185
R2346 VDD.n4349 VDD.n4348 185
R2347 VDD.n465 VDD.n464 185
R2348 VDD.n466 VDD.n465 185
R2349 VDD.n4339 VDD.n4338 185
R2350 VDD.n4340 VDD.n4339 185
R2351 VDD.n474 VDD.n473 185
R2352 VDD.n473 VDD.n472 185
R2353 VDD.n4334 VDD.n4333 185
R2354 VDD.n4333 VDD.n4332 185
R2355 VDD.n477 VDD.n476 185
R2356 VDD.n478 VDD.n477 185
R2357 VDD.n4323 VDD.n4322 185
R2358 VDD.n4324 VDD.n4323 185
R2359 VDD.n486 VDD.n485 185
R2360 VDD.n485 VDD.n484 185
R2361 VDD.n4318 VDD.n4317 185
R2362 VDD.n4317 VDD.n4316 185
R2363 VDD.n489 VDD.n488 185
R2364 VDD.n490 VDD.n489 185
R2365 VDD.n4307 VDD.n4306 185
R2366 VDD.n4308 VDD.n4307 185
R2367 VDD.n498 VDD.n497 185
R2368 VDD.n497 VDD.n496 185
R2369 VDD.n4302 VDD.n4301 185
R2370 VDD.n4301 VDD.n4300 185
R2371 VDD.n501 VDD.n500 185
R2372 VDD.n502 VDD.n501 185
R2373 VDD.n4291 VDD.n4290 185
R2374 VDD.n4292 VDD.n4291 185
R2375 VDD.n510 VDD.n509 185
R2376 VDD.n509 VDD.n508 185
R2377 VDD.n4286 VDD.n4285 185
R2378 VDD.n4285 VDD.n4284 185
R2379 VDD.n513 VDD.n512 185
R2380 VDD.n514 VDD.n513 185
R2381 VDD.n4275 VDD.n4274 185
R2382 VDD.n4276 VDD.n4275 185
R2383 VDD.n521 VDD.n520 185
R2384 VDD.n526 VDD.n520 185
R2385 VDD.n4270 VDD.n4269 185
R2386 VDD.n4269 VDD.n4268 185
R2387 VDD.n524 VDD.n523 185
R2388 VDD.n525 VDD.n524 185
R2389 VDD.n4259 VDD.n4258 185
R2390 VDD.n4260 VDD.n4259 185
R2391 VDD.n534 VDD.n533 185
R2392 VDD.n533 VDD.n532 185
R2393 VDD.n4254 VDD.n4253 185
R2394 VDD.n4253 VDD.n4252 185
R2395 VDD.n537 VDD.n536 185
R2396 VDD.n538 VDD.n537 185
R2397 VDD.n1035 VDD.n1034 185
R2398 VDD.n3402 VDD.n3400 185
R2399 VDD.n3403 VDD.n3399 185
R2400 VDD.n3403 VDD.n3386 185
R2401 VDD.n3406 VDD.n3405 185
R2402 VDD.n3407 VDD.n3398 185
R2403 VDD.n3409 VDD.n3408 185
R2404 VDD.n3411 VDD.n3397 185
R2405 VDD.n3414 VDD.n3413 185
R2406 VDD.n3415 VDD.n3396 185
R2407 VDD.n3417 VDD.n3416 185
R2408 VDD.n3419 VDD.n3395 185
R2409 VDD.n3422 VDD.n3421 185
R2410 VDD.n3423 VDD.n3394 185
R2411 VDD.n3425 VDD.n3424 185
R2412 VDD.n3427 VDD.n3393 185
R2413 VDD.n3430 VDD.n3429 185
R2414 VDD.n3431 VDD.n3390 185
R2415 VDD.n3434 VDD.n3433 185
R2416 VDD.n3436 VDD.n3389 185
R2417 VDD.n3439 VDD.n3438 185
R2418 VDD.n3440 VDD.n3387 185
R2419 VDD.n4174 VDD.n4173 185
R2420 VDD.n4175 VDD.n714 185
R2421 VDD.n4177 VDD.n4176 185
R2422 VDD.n4179 VDD.n713 185
R2423 VDD.n4181 VDD.n4180 185
R2424 VDD.n4182 VDD.n708 185
R2425 VDD.n4184 VDD.n4183 185
R2426 VDD.n4186 VDD.n706 185
R2427 VDD.n4188 VDD.n4187 185
R2428 VDD.n4189 VDD.n705 185
R2429 VDD.n4191 VDD.n4190 185
R2430 VDD.n4193 VDD.n703 185
R2431 VDD.n4195 VDD.n4194 185
R2432 VDD.n4196 VDD.n702 185
R2433 VDD.n4198 VDD.n4197 185
R2434 VDD.n4200 VDD.n700 185
R2435 VDD.n4202 VDD.n4201 185
R2436 VDD.n4203 VDD.n699 185
R2437 VDD.n4205 VDD.n4204 185
R2438 VDD.n4207 VDD.n698 185
R2439 VDD.n4209 VDD.n4208 185
R2440 VDD.n4208 VDD.n679 185
R2441 VDD.n4172 VDD.n4170 185
R2442 VDD.n4172 VDD.n693 185
R2443 VDD.n4169 VDD.n692 185
R2444 VDD.n4213 VDD.n692 185
R2445 VDD.n4168 VDD.n4167 185
R2446 VDD.n4167 VDD.n691 185
R2447 VDD.n4166 VDD.n715 185
R2448 VDD.n4166 VDD.n4165 185
R2449 VDD.n3441 VDD.n716 185
R2450 VDD.n717 VDD.n716 185
R2451 VDD.n3442 VDD.n724 185
R2452 VDD.n4159 VDD.n724 185
R2453 VDD.n3444 VDD.n3443 185
R2454 VDD.n3443 VDD.n723 185
R2455 VDD.n3445 VDD.n731 185
R2456 VDD.n4123 VDD.n731 185
R2457 VDD.n3447 VDD.n3446 185
R2458 VDD.n3446 VDD.n730 185
R2459 VDD.n3448 VDD.n737 185
R2460 VDD.n4117 VDD.n737 185
R2461 VDD.n3450 VDD.n3449 185
R2462 VDD.n3449 VDD.n736 185
R2463 VDD.n3451 VDD.n742 185
R2464 VDD.n4111 VDD.n742 185
R2465 VDD.n3453 VDD.n3452 185
R2466 VDD.n3452 VDD.n750 185
R2467 VDD.n3454 VDD.n748 185
R2468 VDD.n4105 VDD.n748 185
R2469 VDD.n3456 VDD.n3455 185
R2470 VDD.n3455 VDD.n747 185
R2471 VDD.n3457 VDD.n755 185
R2472 VDD.n4099 VDD.n755 185
R2473 VDD.n3459 VDD.n3458 185
R2474 VDD.n3458 VDD.n754 185
R2475 VDD.n3460 VDD.n761 185
R2476 VDD.n4093 VDD.n761 185
R2477 VDD.n3462 VDD.n3461 185
R2478 VDD.n3461 VDD.n760 185
R2479 VDD.n3463 VDD.n767 185
R2480 VDD.n4087 VDD.n767 185
R2481 VDD.n3465 VDD.n3464 185
R2482 VDD.n3464 VDD.n766 185
R2483 VDD.n3466 VDD.n773 185
R2484 VDD.n4081 VDD.n773 185
R2485 VDD.n3468 VDD.n3467 185
R2486 VDD.n3467 VDD.n772 185
R2487 VDD.n3469 VDD.n779 185
R2488 VDD.n4075 VDD.n779 185
R2489 VDD.n3471 VDD.n3470 185
R2490 VDD.n3470 VDD.n778 185
R2491 VDD.n3472 VDD.n785 185
R2492 VDD.n4069 VDD.n785 185
R2493 VDD.n3474 VDD.n3473 185
R2494 VDD.n3473 VDD.n784 185
R2495 VDD.n3475 VDD.n791 185
R2496 VDD.n4063 VDD.n791 185
R2497 VDD.n3477 VDD.n3476 185
R2498 VDD.n3476 VDD.n790 185
R2499 VDD.n3478 VDD.n797 185
R2500 VDD.n4057 VDD.n797 185
R2501 VDD.n3480 VDD.n3479 185
R2502 VDD.n3479 VDD.n796 185
R2503 VDD.n3481 VDD.n803 185
R2504 VDD.n4051 VDD.n803 185
R2505 VDD.n3483 VDD.n3482 185
R2506 VDD.n3482 VDD.n802 185
R2507 VDD.n3484 VDD.n809 185
R2508 VDD.n4045 VDD.n809 185
R2509 VDD.n3486 VDD.n3485 185
R2510 VDD.n3485 VDD.n808 185
R2511 VDD.n3487 VDD.n815 185
R2512 VDD.n4039 VDD.n815 185
R2513 VDD.n3489 VDD.n3488 185
R2514 VDD.n3488 VDD.n814 185
R2515 VDD.n3490 VDD.n820 185
R2516 VDD.n4033 VDD.n820 185
R2517 VDD.n3492 VDD.n3491 185
R2518 VDD.n3491 VDD.n828 185
R2519 VDD.n3493 VDD.n826 185
R2520 VDD.n4027 VDD.n826 185
R2521 VDD.n3495 VDD.n3494 185
R2522 VDD.n3494 VDD.n825 185
R2523 VDD.n3496 VDD.n833 185
R2524 VDD.n4021 VDD.n833 185
R2525 VDD.n3498 VDD.n3497 185
R2526 VDD.n3497 VDD.n832 185
R2527 VDD.n3499 VDD.n839 185
R2528 VDD.n4015 VDD.n839 185
R2529 VDD.n3501 VDD.n3500 185
R2530 VDD.n3500 VDD.n838 185
R2531 VDD.n3502 VDD.n845 185
R2532 VDD.n4009 VDD.n845 185
R2533 VDD.n3504 VDD.n3503 185
R2534 VDD.n3503 VDD.n844 185
R2535 VDD.n3505 VDD.n851 185
R2536 VDD.n4003 VDD.n851 185
R2537 VDD.n3507 VDD.n3506 185
R2538 VDD.n3506 VDD.n850 185
R2539 VDD.n3508 VDD.n857 185
R2540 VDD.n3997 VDD.n857 185
R2541 VDD.n3510 VDD.n3509 185
R2542 VDD.n3509 VDD.n856 185
R2543 VDD.n3511 VDD.n863 185
R2544 VDD.n3991 VDD.n863 185
R2545 VDD.n3513 VDD.n3512 185
R2546 VDD.n3512 VDD.n862 185
R2547 VDD.n3514 VDD.n869 185
R2548 VDD.n3985 VDD.n869 185
R2549 VDD.n3516 VDD.n3515 185
R2550 VDD.n3515 VDD.n868 185
R2551 VDD.n3517 VDD.n875 185
R2552 VDD.n3979 VDD.n875 185
R2553 VDD.n3519 VDD.n3518 185
R2554 VDD.n3518 VDD.n874 185
R2555 VDD.n3520 VDD.n881 185
R2556 VDD.n3973 VDD.n881 185
R2557 VDD.n3522 VDD.n3521 185
R2558 VDD.n3521 VDD.n880 185
R2559 VDD.n3523 VDD.n887 185
R2560 VDD.n3967 VDD.n887 185
R2561 VDD.n3525 VDD.n3524 185
R2562 VDD.n3524 VDD.n886 185
R2563 VDD.n3526 VDD.n893 185
R2564 VDD.n3961 VDD.n893 185
R2565 VDD.n3528 VDD.n3527 185
R2566 VDD.n3527 VDD.n892 185
R2567 VDD.n3529 VDD.n899 185
R2568 VDD.n3955 VDD.n899 185
R2569 VDD.n3531 VDD.n3530 185
R2570 VDD.n3530 VDD.n898 185
R2571 VDD.n3532 VDD.n905 185
R2572 VDD.n3949 VDD.n905 185
R2573 VDD.n3534 VDD.n3533 185
R2574 VDD.n3533 VDD.n904 185
R2575 VDD.n3535 VDD.n911 185
R2576 VDD.n3943 VDD.n911 185
R2577 VDD.n3537 VDD.n3536 185
R2578 VDD.n3536 VDD.n910 185
R2579 VDD.n3538 VDD.n917 185
R2580 VDD.n3937 VDD.n917 185
R2581 VDD.n3540 VDD.n3539 185
R2582 VDD.n3539 VDD.n916 185
R2583 VDD.n3541 VDD.n923 185
R2584 VDD.n3931 VDD.n923 185
R2585 VDD.n3543 VDD.n3542 185
R2586 VDD.n3542 VDD.n922 185
R2587 VDD.n3544 VDD.n929 185
R2588 VDD.n3925 VDD.n929 185
R2589 VDD.n3546 VDD.n3545 185
R2590 VDD.n3545 VDD.n928 185
R2591 VDD.n3547 VDD.n935 185
R2592 VDD.n3919 VDD.n935 185
R2593 VDD.n3549 VDD.n3548 185
R2594 VDD.n3548 VDD.n934 185
R2595 VDD.n3550 VDD.n941 185
R2596 VDD.n3913 VDD.n941 185
R2597 VDD.n3552 VDD.n3551 185
R2598 VDD.n3551 VDD.n940 185
R2599 VDD.n3553 VDD.n947 185
R2600 VDD.n3907 VDD.n947 185
R2601 VDD.n3555 VDD.n3554 185
R2602 VDD.n3554 VDD.n946 185
R2603 VDD.n3556 VDD.n953 185
R2604 VDD.n3901 VDD.n953 185
R2605 VDD.n3558 VDD.n3557 185
R2606 VDD.n3557 VDD.n952 185
R2607 VDD.n3559 VDD.n959 185
R2608 VDD.n3895 VDD.n959 185
R2609 VDD.n3561 VDD.n3560 185
R2610 VDD.n3560 VDD.n958 185
R2611 VDD.n3562 VDD.n965 185
R2612 VDD.n3889 VDD.n965 185
R2613 VDD.n3564 VDD.n3563 185
R2614 VDD.n3563 VDD.n964 185
R2615 VDD.n3565 VDD.n971 185
R2616 VDD.n3883 VDD.n971 185
R2617 VDD.n3567 VDD.n3566 185
R2618 VDD.n3566 VDD.n970 185
R2619 VDD.n3568 VDD.n977 185
R2620 VDD.n3877 VDD.n977 185
R2621 VDD.n3570 VDD.n3569 185
R2622 VDD.n3569 VDD.n976 185
R2623 VDD.n3571 VDD.n983 185
R2624 VDD.n3871 VDD.n983 185
R2625 VDD.n3573 VDD.n3572 185
R2626 VDD.n3572 VDD.n982 185
R2627 VDD.n3574 VDD.n989 185
R2628 VDD.n3865 VDD.n989 185
R2629 VDD.n3576 VDD.n3575 185
R2630 VDD.n3575 VDD.n988 185
R2631 VDD.n3577 VDD.n994 185
R2632 VDD.n3859 VDD.n994 185
R2633 VDD.n3579 VDD.n3578 185
R2634 VDD.n3578 VDD.n1001 185
R2635 VDD.n3580 VDD.n999 185
R2636 VDD.n3853 VDD.n999 185
R2637 VDD.n3582 VDD.n3581 185
R2638 VDD.n3581 VDD.n1008 185
R2639 VDD.n3583 VDD.n1006 185
R2640 VDD.n3847 VDD.n1006 185
R2641 VDD.n3585 VDD.n3584 185
R2642 VDD.n3584 VDD.n1005 185
R2643 VDD.n3586 VDD.n1013 185
R2644 VDD.n3841 VDD.n1013 185
R2645 VDD.n3588 VDD.n3587 185
R2646 VDD.n3587 VDD.n1012 185
R2647 VDD.n3589 VDD.n1019 185
R2648 VDD.n3835 VDD.n1019 185
R2649 VDD.n3591 VDD.n3590 185
R2650 VDD.n3590 VDD.n1018 185
R2651 VDD.n3592 VDD.n1025 185
R2652 VDD.n3829 VDD.n1025 185
R2653 VDD.n3594 VDD.n3593 185
R2654 VDD.n3593 VDD.n1024 185
R2655 VDD.n3595 VDD.n1031 185
R2656 VDD.n3823 VDD.n1031 185
R2657 VDD.n3596 VDD.n3388 185
R2658 VDD.n3388 VDD.n1030 185
R2659 VDD.n3598 VDD.n3597 185
R2660 VDD.n3817 VDD.n3598 185
R2661 VDD.n3819 VDD.n3818 185
R2662 VDD.n3818 VDD.n3817 185
R2663 VDD.n3820 VDD.n1033 185
R2664 VDD.n1033 VDD.n1030 185
R2665 VDD.n3822 VDD.n3821 185
R2666 VDD.n3823 VDD.n3822 185
R2667 VDD.n1023 VDD.n1022 185
R2668 VDD.n1024 VDD.n1023 185
R2669 VDD.n3831 VDD.n3830 185
R2670 VDD.n3830 VDD.n3829 185
R2671 VDD.n3832 VDD.n1021 185
R2672 VDD.n1021 VDD.n1018 185
R2673 VDD.n3834 VDD.n3833 185
R2674 VDD.n3835 VDD.n3834 185
R2675 VDD.n1011 VDD.n1010 185
R2676 VDD.n1012 VDD.n1011 185
R2677 VDD.n3843 VDD.n3842 185
R2678 VDD.n3842 VDD.n3841 185
R2679 VDD.n3844 VDD.n1009 185
R2680 VDD.n1009 VDD.n1005 185
R2681 VDD.n3846 VDD.n3845 185
R2682 VDD.n3847 VDD.n3846 185
R2683 VDD.n998 VDD.n997 185
R2684 VDD.n1008 VDD.n998 185
R2685 VDD.n3855 VDD.n3854 185
R2686 VDD.n3854 VDD.n3853 185
R2687 VDD.n3856 VDD.n996 185
R2688 VDD.n1001 VDD.n996 185
R2689 VDD.n3858 VDD.n3857 185
R2690 VDD.n3859 VDD.n3858 185
R2691 VDD.n987 VDD.n986 185
R2692 VDD.n988 VDD.n987 185
R2693 VDD.n3867 VDD.n3866 185
R2694 VDD.n3866 VDD.n3865 185
R2695 VDD.n3868 VDD.n985 185
R2696 VDD.n985 VDD.n982 185
R2697 VDD.n3870 VDD.n3869 185
R2698 VDD.n3871 VDD.n3870 185
R2699 VDD.n975 VDD.n974 185
R2700 VDD.n976 VDD.n975 185
R2701 VDD.n3879 VDD.n3878 185
R2702 VDD.n3878 VDD.n3877 185
R2703 VDD.n3880 VDD.n973 185
R2704 VDD.n973 VDD.n970 185
R2705 VDD.n3882 VDD.n3881 185
R2706 VDD.n3883 VDD.n3882 185
R2707 VDD.n963 VDD.n962 185
R2708 VDD.n964 VDD.n963 185
R2709 VDD.n3891 VDD.n3890 185
R2710 VDD.n3890 VDD.n3889 185
R2711 VDD.n3892 VDD.n961 185
R2712 VDD.n961 VDD.n958 185
R2713 VDD.n3894 VDD.n3893 185
R2714 VDD.n3895 VDD.n3894 185
R2715 VDD.n951 VDD.n950 185
R2716 VDD.n952 VDD.n951 185
R2717 VDD.n3903 VDD.n3902 185
R2718 VDD.n3902 VDD.n3901 185
R2719 VDD.n3904 VDD.n949 185
R2720 VDD.n949 VDD.n946 185
R2721 VDD.n3906 VDD.n3905 185
R2722 VDD.n3907 VDD.n3906 185
R2723 VDD.n939 VDD.n938 185
R2724 VDD.n940 VDD.n939 185
R2725 VDD.n3915 VDD.n3914 185
R2726 VDD.n3914 VDD.n3913 185
R2727 VDD.n3916 VDD.n937 185
R2728 VDD.n937 VDD.n934 185
R2729 VDD.n3918 VDD.n3917 185
R2730 VDD.n3919 VDD.n3918 185
R2731 VDD.n927 VDD.n926 185
R2732 VDD.n928 VDD.n927 185
R2733 VDD.n3927 VDD.n3926 185
R2734 VDD.n3926 VDD.n3925 185
R2735 VDD.n3928 VDD.n925 185
R2736 VDD.n925 VDD.n922 185
R2737 VDD.n3930 VDD.n3929 185
R2738 VDD.n3931 VDD.n3930 185
R2739 VDD.n915 VDD.n914 185
R2740 VDD.n916 VDD.n915 185
R2741 VDD.n3939 VDD.n3938 185
R2742 VDD.n3938 VDD.n3937 185
R2743 VDD.n3940 VDD.n913 185
R2744 VDD.n913 VDD.n910 185
R2745 VDD.n3942 VDD.n3941 185
R2746 VDD.n3943 VDD.n3942 185
R2747 VDD.n903 VDD.n902 185
R2748 VDD.n904 VDD.n903 185
R2749 VDD.n3951 VDD.n3950 185
R2750 VDD.n3950 VDD.n3949 185
R2751 VDD.n3952 VDD.n901 185
R2752 VDD.n901 VDD.n898 185
R2753 VDD.n3954 VDD.n3953 185
R2754 VDD.n3955 VDD.n3954 185
R2755 VDD.n891 VDD.n890 185
R2756 VDD.n892 VDD.n891 185
R2757 VDD.n3963 VDD.n3962 185
R2758 VDD.n3962 VDD.n3961 185
R2759 VDD.n3964 VDD.n889 185
R2760 VDD.n889 VDD.n886 185
R2761 VDD.n3966 VDD.n3965 185
R2762 VDD.n3967 VDD.n3966 185
R2763 VDD.n879 VDD.n878 185
R2764 VDD.n880 VDD.n879 185
R2765 VDD.n3975 VDD.n3974 185
R2766 VDD.n3974 VDD.n3973 185
R2767 VDD.n3976 VDD.n877 185
R2768 VDD.n877 VDD.n874 185
R2769 VDD.n3978 VDD.n3977 185
R2770 VDD.n3979 VDD.n3978 185
R2771 VDD.n867 VDD.n866 185
R2772 VDD.n868 VDD.n867 185
R2773 VDD.n3987 VDD.n3986 185
R2774 VDD.n3986 VDD.n3985 185
R2775 VDD.n3988 VDD.n865 185
R2776 VDD.n865 VDD.n862 185
R2777 VDD.n3990 VDD.n3989 185
R2778 VDD.n3991 VDD.n3990 185
R2779 VDD.n855 VDD.n854 185
R2780 VDD.n856 VDD.n855 185
R2781 VDD.n3999 VDD.n3998 185
R2782 VDD.n3998 VDD.n3997 185
R2783 VDD.n4000 VDD.n853 185
R2784 VDD.n853 VDD.n850 185
R2785 VDD.n4002 VDD.n4001 185
R2786 VDD.n4003 VDD.n4002 185
R2787 VDD.n843 VDD.n842 185
R2788 VDD.n844 VDD.n843 185
R2789 VDD.n4011 VDD.n4010 185
R2790 VDD.n4010 VDD.n4009 185
R2791 VDD.n4012 VDD.n841 185
R2792 VDD.n841 VDD.n838 185
R2793 VDD.n4014 VDD.n4013 185
R2794 VDD.n4015 VDD.n4014 185
R2795 VDD.n831 VDD.n830 185
R2796 VDD.n832 VDD.n831 185
R2797 VDD.n4023 VDD.n4022 185
R2798 VDD.n4022 VDD.n4021 185
R2799 VDD.n4024 VDD.n829 185
R2800 VDD.n829 VDD.n825 185
R2801 VDD.n4026 VDD.n4025 185
R2802 VDD.n4027 VDD.n4026 185
R2803 VDD.n819 VDD.n818 185
R2804 VDD.n828 VDD.n819 185
R2805 VDD.n4035 VDD.n4034 185
R2806 VDD.n4034 VDD.n4033 185
R2807 VDD.n4036 VDD.n817 185
R2808 VDD.n817 VDD.n814 185
R2809 VDD.n4038 VDD.n4037 185
R2810 VDD.n4039 VDD.n4038 185
R2811 VDD.n807 VDD.n806 185
R2812 VDD.n808 VDD.n807 185
R2813 VDD.n4047 VDD.n4046 185
R2814 VDD.n4046 VDD.n4045 185
R2815 VDD.n4048 VDD.n805 185
R2816 VDD.n805 VDD.n802 185
R2817 VDD.n4050 VDD.n4049 185
R2818 VDD.n4051 VDD.n4050 185
R2819 VDD.n795 VDD.n794 185
R2820 VDD.n796 VDD.n795 185
R2821 VDD.n4059 VDD.n4058 185
R2822 VDD.n4058 VDD.n4057 185
R2823 VDD.n4060 VDD.n793 185
R2824 VDD.n793 VDD.n790 185
R2825 VDD.n4062 VDD.n4061 185
R2826 VDD.n4063 VDD.n4062 185
R2827 VDD.n783 VDD.n782 185
R2828 VDD.n784 VDD.n783 185
R2829 VDD.n4071 VDD.n4070 185
R2830 VDD.n4070 VDD.n4069 185
R2831 VDD.n4072 VDD.n781 185
R2832 VDD.n781 VDD.n778 185
R2833 VDD.n4074 VDD.n4073 185
R2834 VDD.n4075 VDD.n4074 185
R2835 VDD.n771 VDD.n770 185
R2836 VDD.n772 VDD.n771 185
R2837 VDD.n4083 VDD.n4082 185
R2838 VDD.n4082 VDD.n4081 185
R2839 VDD.n4084 VDD.n769 185
R2840 VDD.n769 VDD.n766 185
R2841 VDD.n4086 VDD.n4085 185
R2842 VDD.n4087 VDD.n4086 185
R2843 VDD.n759 VDD.n758 185
R2844 VDD.n760 VDD.n759 185
R2845 VDD.n4095 VDD.n4094 185
R2846 VDD.n4094 VDD.n4093 185
R2847 VDD.n4096 VDD.n757 185
R2848 VDD.n757 VDD.n754 185
R2849 VDD.n4098 VDD.n4097 185
R2850 VDD.n4099 VDD.n4098 185
R2851 VDD.n746 VDD.n745 185
R2852 VDD.n747 VDD.n746 185
R2853 VDD.n4107 VDD.n4106 185
R2854 VDD.n4106 VDD.n4105 185
R2855 VDD.n4108 VDD.n744 185
R2856 VDD.n750 VDD.n744 185
R2857 VDD.n4110 VDD.n4109 185
R2858 VDD.n4111 VDD.n4110 185
R2859 VDD.n735 VDD.n734 185
R2860 VDD.n736 VDD.n735 185
R2861 VDD.n4119 VDD.n4118 185
R2862 VDD.n4118 VDD.n4117 185
R2863 VDD.n4120 VDD.n733 185
R2864 VDD.n733 VDD.n730 185
R2865 VDD.n4122 VDD.n4121 185
R2866 VDD.n4123 VDD.n4122 185
R2867 VDD.n722 VDD.n721 185
R2868 VDD.n723 VDD.n722 185
R2869 VDD.n4161 VDD.n4160 185
R2870 VDD.n4160 VDD.n4159 185
R2871 VDD.n4162 VDD.n720 185
R2872 VDD.n720 VDD.n717 185
R2873 VDD.n4164 VDD.n4163 185
R2874 VDD.n4165 VDD.n4164 185
R2875 VDD.n697 VDD.n695 185
R2876 VDD.n695 VDD.n691 185
R2877 VDD.n4212 VDD.n4211 185
R2878 VDD.n4213 VDD.n4212 185
R2879 VDD.n4210 VDD.n696 185
R2880 VDD.n696 VDD.n693 185
R2881 VDD.n2909 VDD.n2908 185
R2882 VDD.n2911 VDD.n1831 185
R2883 VDD.n2912 VDD.n1830 185
R2884 VDD.n2904 VDD.n1828 185
R2885 VDD.n2916 VDD.n1827 185
R2886 VDD.n2917 VDD.n1826 185
R2887 VDD.n2918 VDD.n1825 185
R2888 VDD.n2901 VDD.n1823 185
R2889 VDD.n2922 VDD.n1822 185
R2890 VDD.n2923 VDD.n1821 185
R2891 VDD.n2924 VDD.n1820 185
R2892 VDD.n2898 VDD.n1818 185
R2893 VDD.n2928 VDD.n1817 185
R2894 VDD.n2929 VDD.n1816 185
R2895 VDD.n2931 VDD.n1813 185
R2896 VDD.n2895 VDD.n1811 185
R2897 VDD.n2935 VDD.n1810 185
R2898 VDD.n2936 VDD.n1809 185
R2899 VDD.n2937 VDD.n1808 185
R2900 VDD.n2892 VDD.n1807 185
R2901 VDD.n2891 VDD.n2890 185
R2902 VDD.n2884 VDD.n1846 185
R2903 VDD.n2886 VDD.n2885 185
R2904 VDD.n2883 VDD.n2882 185
R2905 VDD.n2881 VDD.n2880 185
R2906 VDD.n2874 VDD.n1848 185
R2907 VDD.n2876 VDD.n2875 185
R2908 VDD.n2870 VDD.n2869 185
R2909 VDD.n2868 VDD.n2867 185
R2910 VDD.n2861 VDD.n1850 185
R2911 VDD.n2863 VDD.n2862 185
R2912 VDD.n2860 VDD.n2859 185
R2913 VDD.n2858 VDD.n2857 185
R2914 VDD.n2851 VDD.n1852 185
R2915 VDD.n2853 VDD.n2852 185
R2916 VDD.n2850 VDD.n2849 185
R2917 VDD.n2848 VDD.n2847 185
R2918 VDD.n2844 VDD.n2843 185
R2919 VDD.n1862 VDD.n1835 185
R2920 VDD.n1836 VDD.n1835 185
R2921 VDD.n2833 VDD.n2832 185
R2922 VDD.n2834 VDD.n2833 185
R2923 VDD.n1861 VDD.n1860 185
R2924 VDD.n2835 VDD.n1860 185
R2925 VDD.n2826 VDD.n2825 185
R2926 VDD.n2825 VDD.n1859 185
R2927 VDD.n2824 VDD.n1864 185
R2928 VDD.n2824 VDD.n2823 185
R2929 VDD.n1874 VDD.n1865 185
R2930 VDD.n1866 VDD.n1865 185
R2931 VDD.n2814 VDD.n2813 185
R2932 VDD.n2815 VDD.n2814 185
R2933 VDD.n1873 VDD.n1872 185
R2934 VDD.n1879 VDD.n1872 185
R2935 VDD.n2808 VDD.n2807 185
R2936 VDD.n2807 VDD.n2806 185
R2937 VDD.n1877 VDD.n1876 185
R2938 VDD.n1878 VDD.n1877 185
R2939 VDD.n2797 VDD.n2796 185
R2940 VDD.n2798 VDD.n2797 185
R2941 VDD.n1887 VDD.n1886 185
R2942 VDD.n1886 VDD.n1885 185
R2943 VDD.n2792 VDD.n2791 185
R2944 VDD.n2791 VDD.n2790 185
R2945 VDD.n1890 VDD.n1889 185
R2946 VDD.n1891 VDD.n1890 185
R2947 VDD.n2781 VDD.n2780 185
R2948 VDD.n2782 VDD.n2781 185
R2949 VDD.n1899 VDD.n1898 185
R2950 VDD.n1898 VDD.n1897 185
R2951 VDD.n2776 VDD.n2775 185
R2952 VDD.n2775 VDD.n2774 185
R2953 VDD.n1902 VDD.n1901 185
R2954 VDD.n1903 VDD.n1902 185
R2955 VDD.n2765 VDD.n2764 185
R2956 VDD.n2766 VDD.n2765 185
R2957 VDD.n1911 VDD.n1910 185
R2958 VDD.n1910 VDD.n1909 185
R2959 VDD.n2760 VDD.n2759 185
R2960 VDD.n2759 VDD.n2758 185
R2961 VDD.n1914 VDD.n1913 185
R2962 VDD.n1915 VDD.n1914 185
R2963 VDD.n2749 VDD.n2748 185
R2964 VDD.n2750 VDD.n2749 185
R2965 VDD.n1923 VDD.n1922 185
R2966 VDD.n1922 VDD.n1921 185
R2967 VDD.n2744 VDD.n2743 185
R2968 VDD.n2743 VDD.n2742 185
R2969 VDD.n1926 VDD.n1925 185
R2970 VDD.n1927 VDD.n1926 185
R2971 VDD.n2733 VDD.n2732 185
R2972 VDD.n2734 VDD.n2733 185
R2973 VDD.n1935 VDD.n1934 185
R2974 VDD.n1934 VDD.n1933 185
R2975 VDD.n2728 VDD.n2727 185
R2976 VDD.n2727 VDD.n2726 185
R2977 VDD.n1938 VDD.n1937 185
R2978 VDD.n1939 VDD.n1938 185
R2979 VDD.n2717 VDD.n2716 185
R2980 VDD.n2718 VDD.n2717 185
R2981 VDD.n1947 VDD.n1946 185
R2982 VDD.n1946 VDD.n1945 185
R2983 VDD.n2712 VDD.n2711 185
R2984 VDD.n2711 VDD.n2710 185
R2985 VDD.n1950 VDD.n1949 185
R2986 VDD.n1951 VDD.n1950 185
R2987 VDD.n2701 VDD.n2700 185
R2988 VDD.n2702 VDD.n2701 185
R2989 VDD.n1959 VDD.n1958 185
R2990 VDD.n1958 VDD.n1957 185
R2991 VDD.n2696 VDD.n2695 185
R2992 VDD.n2695 VDD.n2694 185
R2993 VDD.n1962 VDD.n1961 185
R2994 VDD.n1963 VDD.n1962 185
R2995 VDD.n2685 VDD.n2684 185
R2996 VDD.n2686 VDD.n2685 185
R2997 VDD.n1971 VDD.n1970 185
R2998 VDD.n1970 VDD.n1969 185
R2999 VDD.n2680 VDD.n2679 185
R3000 VDD.n2679 VDD.n2678 185
R3001 VDD.n1974 VDD.n1973 185
R3002 VDD.n1975 VDD.n1974 185
R3003 VDD.n2669 VDD.n2668 185
R3004 VDD.n2670 VDD.n2669 185
R3005 VDD.n1983 VDD.n1982 185
R3006 VDD.n1982 VDD.n1981 185
R3007 VDD.n2664 VDD.n2663 185
R3008 VDD.n2663 VDD.n2662 185
R3009 VDD.n1986 VDD.n1985 185
R3010 VDD.n1987 VDD.n1986 185
R3011 VDD.n2653 VDD.n2652 185
R3012 VDD.n2654 VDD.n2653 185
R3013 VDD.n1994 VDD.n1993 185
R3014 VDD.n1999 VDD.n1993 185
R3015 VDD.n2648 VDD.n2647 185
R3016 VDD.n2647 VDD.n2646 185
R3017 VDD.n1997 VDD.n1996 185
R3018 VDD.n1998 VDD.n1997 185
R3019 VDD.n2637 VDD.n2636 185
R3020 VDD.n2638 VDD.n2637 185
R3021 VDD.n2007 VDD.n2006 185
R3022 VDD.n2006 VDD.n2005 185
R3023 VDD.n2632 VDD.n2631 185
R3024 VDD.n2631 VDD.n2630 185
R3025 VDD.n2010 VDD.n2009 185
R3026 VDD.n2011 VDD.n2010 185
R3027 VDD.n2621 VDD.n2620 185
R3028 VDD.n2622 VDD.n2621 185
R3029 VDD.n2019 VDD.n2018 185
R3030 VDD.n2018 VDD.n2017 185
R3031 VDD.n2616 VDD.n2615 185
R3032 VDD.n2615 VDD.n2614 185
R3033 VDD.n2022 VDD.n2021 185
R3034 VDD.n2023 VDD.n2022 185
R3035 VDD.n2605 VDD.n2604 185
R3036 VDD.n2606 VDD.n2605 185
R3037 VDD.n2051 VDD.n2050 185
R3038 VDD.n2056 VDD.n2050 185
R3039 VDD.n2600 VDD.n2599 185
R3040 VDD.n2599 VDD.n2598 185
R3041 VDD.n2054 VDD.n2053 185
R3042 VDD.n2055 VDD.n2054 185
R3043 VDD.n2588 VDD.n2587 185
R3044 VDD.n2589 VDD.n2588 185
R3045 VDD.n2064 VDD.n2063 185
R3046 VDD.n2063 VDD.n2062 185
R3047 VDD.n2583 VDD.n2582 185
R3048 VDD.n2582 VDD.n2581 185
R3049 VDD.n2067 VDD.n2066 185
R3050 VDD.n2068 VDD.n2067 185
R3051 VDD.n2572 VDD.n2571 185
R3052 VDD.n2573 VDD.n2572 185
R3053 VDD.n2076 VDD.n2075 185
R3054 VDD.n2075 VDD.n2074 185
R3055 VDD.n2567 VDD.n2566 185
R3056 VDD.n2566 VDD.n2565 185
R3057 VDD.n2079 VDD.n2078 185
R3058 VDD.n2080 VDD.n2079 185
R3059 VDD.n2556 VDD.n2555 185
R3060 VDD.n2557 VDD.n2556 185
R3061 VDD.n2087 VDD.n2086 185
R3062 VDD.n2092 VDD.n2086 185
R3063 VDD.n2551 VDD.n2550 185
R3064 VDD.n2550 VDD.n2549 185
R3065 VDD.n2090 VDD.n2089 185
R3066 VDD.n2091 VDD.n2090 185
R3067 VDD.n2540 VDD.n2539 185
R3068 VDD.n2541 VDD.n2540 185
R3069 VDD.n2100 VDD.n2099 185
R3070 VDD.n2099 VDD.n2098 185
R3071 VDD.n2535 VDD.n2534 185
R3072 VDD.n2534 VDD.n2533 185
R3073 VDD.n2103 VDD.n2102 185
R3074 VDD.n2104 VDD.n2103 185
R3075 VDD.n2524 VDD.n2523 185
R3076 VDD.n2525 VDD.n2524 185
R3077 VDD.n2112 VDD.n2111 185
R3078 VDD.n2111 VDD.n2110 185
R3079 VDD.n2519 VDD.n2518 185
R3080 VDD.n2518 VDD.n2517 185
R3081 VDD.n2115 VDD.n2114 185
R3082 VDD.n2116 VDD.n2115 185
R3083 VDD.n2508 VDD.n2507 185
R3084 VDD.n2509 VDD.n2508 185
R3085 VDD.n2124 VDD.n2123 185
R3086 VDD.n2123 VDD.n2122 185
R3087 VDD.n2503 VDD.n2502 185
R3088 VDD.n2502 VDD.n2501 185
R3089 VDD.n2127 VDD.n2126 185
R3090 VDD.n2128 VDD.n2127 185
R3091 VDD.n2492 VDD.n2491 185
R3092 VDD.n2493 VDD.n2492 185
R3093 VDD.n2136 VDD.n2135 185
R3094 VDD.n2135 VDD.n2134 185
R3095 VDD.n2487 VDD.n2486 185
R3096 VDD.n2486 VDD.n2485 185
R3097 VDD.n2139 VDD.n2138 185
R3098 VDD.n2140 VDD.n2139 185
R3099 VDD.n2476 VDD.n2475 185
R3100 VDD.n2477 VDD.n2476 185
R3101 VDD.n2148 VDD.n2147 185
R3102 VDD.n2147 VDD.n2146 185
R3103 VDD.n2471 VDD.n2470 185
R3104 VDD.n2470 VDD.n2469 185
R3105 VDD.n2151 VDD.n2150 185
R3106 VDD.n2152 VDD.n2151 185
R3107 VDD.n2460 VDD.n2459 185
R3108 VDD.n2461 VDD.n2460 185
R3109 VDD.n2160 VDD.n2159 185
R3110 VDD.n2159 VDD.n2158 185
R3111 VDD.n2455 VDD.n2454 185
R3112 VDD.n2454 VDD.n2453 185
R3113 VDD.n2163 VDD.n2162 185
R3114 VDD.n2164 VDD.n2163 185
R3115 VDD.n2444 VDD.n2443 185
R3116 VDD.n2445 VDD.n2444 185
R3117 VDD.n2172 VDD.n2171 185
R3118 VDD.n2171 VDD.n2170 185
R3119 VDD.n2439 VDD.n2438 185
R3120 VDD.n2438 VDD.n2437 185
R3121 VDD.n2175 VDD.n2174 185
R3122 VDD.n2176 VDD.n2175 185
R3123 VDD.n2428 VDD.n2427 185
R3124 VDD.n2429 VDD.n2428 185
R3125 VDD.n2184 VDD.n2183 185
R3126 VDD.n2183 VDD.n2182 185
R3127 VDD.n2423 VDD.n2422 185
R3128 VDD.n2422 VDD.n2421 185
R3129 VDD.n2187 VDD.n2186 185
R3130 VDD.n2188 VDD.n2187 185
R3131 VDD.n2412 VDD.n2411 185
R3132 VDD.n2413 VDD.n2412 185
R3133 VDD.n2196 VDD.n2195 185
R3134 VDD.n2195 VDD.n2194 185
R3135 VDD.n2407 VDD.n2406 185
R3136 VDD.n2406 VDD.n2405 185
R3137 VDD.n2199 VDD.n2198 185
R3138 VDD.n2200 VDD.n2199 185
R3139 VDD.n2396 VDD.n2395 185
R3140 VDD.n2397 VDD.n2396 185
R3141 VDD.n2207 VDD.n2206 185
R3142 VDD.n2212 VDD.n2206 185
R3143 VDD.n2391 VDD.n2390 185
R3144 VDD.n2390 VDD.n2389 185
R3145 VDD.n2210 VDD.n2209 185
R3146 VDD.n2211 VDD.n2210 185
R3147 VDD.n2380 VDD.n2379 185
R3148 VDD.n2381 VDD.n2380 185
R3149 VDD.n2220 VDD.n2219 185
R3150 VDD.n2219 VDD.n2218 185
R3151 VDD.n2375 VDD.n2374 185
R3152 VDD.n2374 VDD.n2373 185
R3153 VDD.n2223 VDD.n2222 185
R3154 VDD.n2224 VDD.n2223 185
R3155 VDD.n2367 VDD.n2366 185
R3156 VDD.n2229 VDD.n2228 185
R3157 VDD.n2363 VDD.n2362 185
R3158 VDD.n2364 VDD.n2363 185
R3159 VDD.n2249 VDD.n2248 185
R3160 VDD.n2358 VDD.n2251 185
R3161 VDD.n2357 VDD.n2252 185
R3162 VDD.n2356 VDD.n2253 185
R3163 VDD.n2255 VDD.n2254 185
R3164 VDD.n2352 VDD.n2257 185
R3165 VDD.n2351 VDD.n2258 185
R3166 VDD.n2350 VDD.n2259 185
R3167 VDD.n2347 VDD.n2264 185
R3168 VDD.n2346 VDD.n2265 185
R3169 VDD.n2345 VDD.n2266 185
R3170 VDD.n2269 VDD.n2267 185
R3171 VDD.n2341 VDD.n2270 185
R3172 VDD.n2340 VDD.n2271 185
R3173 VDD.n2339 VDD.n2272 185
R3174 VDD.n2275 VDD.n2273 185
R3175 VDD.n2335 VDD.n2276 185
R3176 VDD.n2334 VDD.n2277 185
R3177 VDD.n2333 VDD.n2278 185
R3178 VDD.n2281 VDD.n2279 185
R3179 VDD.n2329 VDD.n2282 185
R3180 VDD.n2325 VDD.n2283 185
R3181 VDD.n2324 VDD.n2284 185
R3182 VDD.n2287 VDD.n2285 185
R3183 VDD.n2320 VDD.n2288 185
R3184 VDD.n2319 VDD.n2289 185
R3185 VDD.n2318 VDD.n2290 185
R3186 VDD.n2293 VDD.n2291 185
R3187 VDD.n2314 VDD.n2294 185
R3188 VDD.n2313 VDD.n2295 185
R3189 VDD.n2312 VDD.n2296 185
R3190 VDD.n2299 VDD.n2297 185
R3191 VDD.n2308 VDD.n2300 185
R3192 VDD.n2307 VDD.n2301 185
R3193 VDD.n2303 VDD.n2247 185
R3194 VDD.n2364 VDD.n2247 185
R3195 VDD.n2842 VDD.n2841 185
R3196 VDD.n2842 VDD.n1836 185
R3197 VDD.n1855 VDD.n1854 185
R3198 VDD.n2834 VDD.n1854 185
R3199 VDD.n2837 VDD.n2836 185
R3200 VDD.n2836 VDD.n2835 185
R3201 VDD.n1858 VDD.n1857 185
R3202 VDD.n1859 VDD.n1858 185
R3203 VDD.n2822 VDD.n2821 185
R3204 VDD.n2823 VDD.n2822 185
R3205 VDD.n1868 VDD.n1867 185
R3206 VDD.n1867 VDD.n1866 185
R3207 VDD.n2817 VDD.n2816 185
R3208 VDD.n2816 VDD.n2815 185
R3209 VDD.n1871 VDD.n1870 185
R3210 VDD.n1879 VDD.n1871 185
R3211 VDD.n2805 VDD.n2804 185
R3212 VDD.n2806 VDD.n2805 185
R3213 VDD.n1881 VDD.n1880 185
R3214 VDD.n1880 VDD.n1878 185
R3215 VDD.n2800 VDD.n2799 185
R3216 VDD.n2799 VDD.n2798 185
R3217 VDD.n1884 VDD.n1883 185
R3218 VDD.n1885 VDD.n1884 185
R3219 VDD.n2789 VDD.n2788 185
R3220 VDD.n2790 VDD.n2789 185
R3221 VDD.n1893 VDD.n1892 185
R3222 VDD.n1892 VDD.n1891 185
R3223 VDD.n2784 VDD.n2783 185
R3224 VDD.n2783 VDD.n2782 185
R3225 VDD.n1896 VDD.n1895 185
R3226 VDD.n1897 VDD.n1896 185
R3227 VDD.n2773 VDD.n2772 185
R3228 VDD.n2774 VDD.n2773 185
R3229 VDD.n1905 VDD.n1904 185
R3230 VDD.n1904 VDD.n1903 185
R3231 VDD.n2768 VDD.n2767 185
R3232 VDD.n2767 VDD.n2766 185
R3233 VDD.n1908 VDD.n1907 185
R3234 VDD.n1909 VDD.n1908 185
R3235 VDD.n2757 VDD.n2756 185
R3236 VDD.n2758 VDD.n2757 185
R3237 VDD.n1917 VDD.n1916 185
R3238 VDD.n1916 VDD.n1915 185
R3239 VDD.n2752 VDD.n2751 185
R3240 VDD.n2751 VDD.n2750 185
R3241 VDD.n1920 VDD.n1919 185
R3242 VDD.n1921 VDD.n1920 185
R3243 VDD.n2741 VDD.n2740 185
R3244 VDD.n2742 VDD.n2741 185
R3245 VDD.n1929 VDD.n1928 185
R3246 VDD.n1928 VDD.n1927 185
R3247 VDD.n2736 VDD.n2735 185
R3248 VDD.n2735 VDD.n2734 185
R3249 VDD.n1932 VDD.n1931 185
R3250 VDD.n1933 VDD.n1932 185
R3251 VDD.n2725 VDD.n2724 185
R3252 VDD.n2726 VDD.n2725 185
R3253 VDD.n1941 VDD.n1940 185
R3254 VDD.n1940 VDD.n1939 185
R3255 VDD.n2720 VDD.n2719 185
R3256 VDD.n2719 VDD.n2718 185
R3257 VDD.n1944 VDD.n1943 185
R3258 VDD.n1945 VDD.n1944 185
R3259 VDD.n2709 VDD.n2708 185
R3260 VDD.n2710 VDD.n2709 185
R3261 VDD.n1953 VDD.n1952 185
R3262 VDD.n1952 VDD.n1951 185
R3263 VDD.n2704 VDD.n2703 185
R3264 VDD.n2703 VDD.n2702 185
R3265 VDD.n1956 VDD.n1955 185
R3266 VDD.n1957 VDD.n1956 185
R3267 VDD.n2693 VDD.n2692 185
R3268 VDD.n2694 VDD.n2693 185
R3269 VDD.n1965 VDD.n1964 185
R3270 VDD.n1964 VDD.n1963 185
R3271 VDD.n2688 VDD.n2687 185
R3272 VDD.n2687 VDD.n2686 185
R3273 VDD.n1968 VDD.n1967 185
R3274 VDD.n1969 VDD.n1968 185
R3275 VDD.n2677 VDD.n2676 185
R3276 VDD.n2678 VDD.n2677 185
R3277 VDD.n1977 VDD.n1976 185
R3278 VDD.n1976 VDD.n1975 185
R3279 VDD.n2672 VDD.n2671 185
R3280 VDD.n2671 VDD.n2670 185
R3281 VDD.n1980 VDD.n1979 185
R3282 VDD.n1981 VDD.n1980 185
R3283 VDD.n2661 VDD.n2660 185
R3284 VDD.n2662 VDD.n2661 185
R3285 VDD.n1989 VDD.n1988 185
R3286 VDD.n1988 VDD.n1987 185
R3287 VDD.n2656 VDD.n2655 185
R3288 VDD.n2655 VDD.n2654 185
R3289 VDD.n1992 VDD.n1991 185
R3290 VDD.n1999 VDD.n1992 185
R3291 VDD.n2645 VDD.n2644 185
R3292 VDD.n2646 VDD.n2645 185
R3293 VDD.n2001 VDD.n2000 185
R3294 VDD.n2000 VDD.n1998 185
R3295 VDD.n2640 VDD.n2639 185
R3296 VDD.n2639 VDD.n2638 185
R3297 VDD.n2004 VDD.n2003 185
R3298 VDD.n2005 VDD.n2004 185
R3299 VDD.n2629 VDD.n2628 185
R3300 VDD.n2630 VDD.n2629 185
R3301 VDD.n2013 VDD.n2012 185
R3302 VDD.n2012 VDD.n2011 185
R3303 VDD.n2624 VDD.n2623 185
R3304 VDD.n2623 VDD.n2622 185
R3305 VDD.n2016 VDD.n2015 185
R3306 VDD.n2017 VDD.n2016 185
R3307 VDD.n2613 VDD.n2612 185
R3308 VDD.n2614 VDD.n2613 185
R3309 VDD.n2025 VDD.n2024 185
R3310 VDD.n2024 VDD.n2023 185
R3311 VDD.n2608 VDD.n2607 185
R3312 VDD.n2607 VDD.n2606 185
R3313 VDD.n2049 VDD.n2048 185
R3314 VDD.n2056 VDD.n2049 185
R3315 VDD.n2597 VDD.n2596 185
R3316 VDD.n2598 VDD.n2597 185
R3317 VDD.n2058 VDD.n2057 185
R3318 VDD.n2057 VDD.n2055 185
R3319 VDD.n2591 VDD.n2590 185
R3320 VDD.n2590 VDD.n2589 185
R3321 VDD.n2061 VDD.n2060 185
R3322 VDD.n2062 VDD.n2061 185
R3323 VDD.n2580 VDD.n2579 185
R3324 VDD.n2581 VDD.n2580 185
R3325 VDD.n2070 VDD.n2069 185
R3326 VDD.n2069 VDD.n2068 185
R3327 VDD.n2575 VDD.n2574 185
R3328 VDD.n2574 VDD.n2573 185
R3329 VDD.n2073 VDD.n2072 185
R3330 VDD.n2074 VDD.n2073 185
R3331 VDD.n2564 VDD.n2563 185
R3332 VDD.n2565 VDD.n2564 185
R3333 VDD.n2082 VDD.n2081 185
R3334 VDD.n2081 VDD.n2080 185
R3335 VDD.n2559 VDD.n2558 185
R3336 VDD.n2558 VDD.n2557 185
R3337 VDD.n2085 VDD.n2084 185
R3338 VDD.n2092 VDD.n2085 185
R3339 VDD.n2548 VDD.n2547 185
R3340 VDD.n2549 VDD.n2548 185
R3341 VDD.n2094 VDD.n2093 185
R3342 VDD.n2093 VDD.n2091 185
R3343 VDD.n2543 VDD.n2542 185
R3344 VDD.n2542 VDD.n2541 185
R3345 VDD.n2097 VDD.n2096 185
R3346 VDD.n2098 VDD.n2097 185
R3347 VDD.n2532 VDD.n2531 185
R3348 VDD.n2533 VDD.n2532 185
R3349 VDD.n2106 VDD.n2105 185
R3350 VDD.n2105 VDD.n2104 185
R3351 VDD.n2527 VDD.n2526 185
R3352 VDD.n2526 VDD.n2525 185
R3353 VDD.n2109 VDD.n2108 185
R3354 VDD.n2110 VDD.n2109 185
R3355 VDD.n2516 VDD.n2515 185
R3356 VDD.n2517 VDD.n2516 185
R3357 VDD.n2118 VDD.n2117 185
R3358 VDD.n2117 VDD.n2116 185
R3359 VDD.n2511 VDD.n2510 185
R3360 VDD.n2510 VDD.n2509 185
R3361 VDD.n2121 VDD.n2120 185
R3362 VDD.n2122 VDD.n2121 185
R3363 VDD.n2500 VDD.n2499 185
R3364 VDD.n2501 VDD.n2500 185
R3365 VDD.n2130 VDD.n2129 185
R3366 VDD.n2129 VDD.n2128 185
R3367 VDD.n2495 VDD.n2494 185
R3368 VDD.n2494 VDD.n2493 185
R3369 VDD.n2133 VDD.n2132 185
R3370 VDD.n2134 VDD.n2133 185
R3371 VDD.n2484 VDD.n2483 185
R3372 VDD.n2485 VDD.n2484 185
R3373 VDD.n2142 VDD.n2141 185
R3374 VDD.n2141 VDD.n2140 185
R3375 VDD.n2479 VDD.n2478 185
R3376 VDD.n2478 VDD.n2477 185
R3377 VDD.n2145 VDD.n2144 185
R3378 VDD.n2146 VDD.n2145 185
R3379 VDD.n2468 VDD.n2467 185
R3380 VDD.n2469 VDD.n2468 185
R3381 VDD.n2154 VDD.n2153 185
R3382 VDD.n2153 VDD.n2152 185
R3383 VDD.n2463 VDD.n2462 185
R3384 VDD.n2462 VDD.n2461 185
R3385 VDD.n2157 VDD.n2156 185
R3386 VDD.n2158 VDD.n2157 185
R3387 VDD.n2452 VDD.n2451 185
R3388 VDD.n2453 VDD.n2452 185
R3389 VDD.n2166 VDD.n2165 185
R3390 VDD.n2165 VDD.n2164 185
R3391 VDD.n2447 VDD.n2446 185
R3392 VDD.n2446 VDD.n2445 185
R3393 VDD.n2169 VDD.n2168 185
R3394 VDD.n2170 VDD.n2169 185
R3395 VDD.n2436 VDD.n2435 185
R3396 VDD.n2437 VDD.n2436 185
R3397 VDD.n2178 VDD.n2177 185
R3398 VDD.n2177 VDD.n2176 185
R3399 VDD.n2431 VDD.n2430 185
R3400 VDD.n2430 VDD.n2429 185
R3401 VDD.n2181 VDD.n2180 185
R3402 VDD.n2182 VDD.n2181 185
R3403 VDD.n2420 VDD.n2419 185
R3404 VDD.n2421 VDD.n2420 185
R3405 VDD.n2190 VDD.n2189 185
R3406 VDD.n2189 VDD.n2188 185
R3407 VDD.n2415 VDD.n2414 185
R3408 VDD.n2414 VDD.n2413 185
R3409 VDD.n2193 VDD.n2192 185
R3410 VDD.n2194 VDD.n2193 185
R3411 VDD.n2404 VDD.n2403 185
R3412 VDD.n2405 VDD.n2404 185
R3413 VDD.n2202 VDD.n2201 185
R3414 VDD.n2201 VDD.n2200 185
R3415 VDD.n2399 VDD.n2398 185
R3416 VDD.n2398 VDD.n2397 185
R3417 VDD.n2205 VDD.n2204 185
R3418 VDD.n2212 VDD.n2205 185
R3419 VDD.n2388 VDD.n2387 185
R3420 VDD.n2389 VDD.n2388 185
R3421 VDD.n2214 VDD.n2213 185
R3422 VDD.n2213 VDD.n2211 185
R3423 VDD.n2383 VDD.n2382 185
R3424 VDD.n2382 VDD.n2381 185
R3425 VDD.n2217 VDD.n2216 185
R3426 VDD.n2218 VDD.n2217 185
R3427 VDD.n2372 VDD.n2371 185
R3428 VDD.n2373 VDD.n2372 185
R3429 VDD.n2226 VDD.n2225 185
R3430 VDD.n2225 VDD.n2224 185
R3431 VDD.n251 VDD.n250 146.341
R3432 VDD.n255 VDD.n254 146.341
R3433 VDD.n261 VDD.n260 146.341
R3434 VDD.n265 VDD.n264 146.341
R3435 VDD.n271 VDD.n270 146.341
R3436 VDD.n276 VDD.n275 146.341
R3437 VDD.n282 VDD.n281 146.341
R3438 VDD.n286 VDD.n285 146.341
R3439 VDD.n292 VDD.n291 146.341
R3440 VDD.n296 VDD.n295 146.341
R3441 VDD.n302 VDD.n301 146.341
R3442 VDD.n306 VDD.n305 146.341
R3443 VDD.n312 VDD.n311 146.341
R3444 VDD.n316 VDD.n315 146.341
R3445 VDD.n322 VDD.n321 146.341
R3446 VDD.n326 VDD.n325 146.341
R3447 VDD.n332 VDD.n331 146.341
R3448 VDD.n334 VDD.n217 146.341
R3449 VDD.n4253 VDD.n537 146.341
R3450 VDD.n4253 VDD.n533 146.341
R3451 VDD.n4259 VDD.n533 146.341
R3452 VDD.n4259 VDD.n524 146.341
R3453 VDD.n4269 VDD.n524 146.341
R3454 VDD.n4269 VDD.n520 146.341
R3455 VDD.n4275 VDD.n520 146.341
R3456 VDD.n4275 VDD.n513 146.341
R3457 VDD.n4285 VDD.n513 146.341
R3458 VDD.n4285 VDD.n509 146.341
R3459 VDD.n4291 VDD.n509 146.341
R3460 VDD.n4291 VDD.n501 146.341
R3461 VDD.n4301 VDD.n501 146.341
R3462 VDD.n4301 VDD.n497 146.341
R3463 VDD.n4307 VDD.n497 146.341
R3464 VDD.n4307 VDD.n489 146.341
R3465 VDD.n4317 VDD.n489 146.341
R3466 VDD.n4317 VDD.n485 146.341
R3467 VDD.n4323 VDD.n485 146.341
R3468 VDD.n4323 VDD.n477 146.341
R3469 VDD.n4333 VDD.n477 146.341
R3470 VDD.n4333 VDD.n473 146.341
R3471 VDD.n4339 VDD.n473 146.341
R3472 VDD.n4339 VDD.n465 146.341
R3473 VDD.n4349 VDD.n465 146.341
R3474 VDD.n4349 VDD.n461 146.341
R3475 VDD.n4355 VDD.n461 146.341
R3476 VDD.n4355 VDD.n453 146.341
R3477 VDD.n4365 VDD.n453 146.341
R3478 VDD.n4365 VDD.n449 146.341
R3479 VDD.n4371 VDD.n449 146.341
R3480 VDD.n4371 VDD.n441 146.341
R3481 VDD.n4381 VDD.n441 146.341
R3482 VDD.n4381 VDD.n437 146.341
R3483 VDD.n4387 VDD.n437 146.341
R3484 VDD.n4387 VDD.n429 146.341
R3485 VDD.n4397 VDD.n429 146.341
R3486 VDD.n4397 VDD.n425 146.341
R3487 VDD.n4403 VDD.n425 146.341
R3488 VDD.n4403 VDD.n417 146.341
R3489 VDD.n4413 VDD.n417 146.341
R3490 VDD.n4413 VDD.n413 146.341
R3491 VDD.n4419 VDD.n413 146.341
R3492 VDD.n4419 VDD.n404 146.341
R3493 VDD.n4429 VDD.n404 146.341
R3494 VDD.n4429 VDD.n400 146.341
R3495 VDD.n4435 VDD.n400 146.341
R3496 VDD.n4435 VDD.n393 146.341
R3497 VDD.n4445 VDD.n393 146.341
R3498 VDD.n4445 VDD.n389 146.341
R3499 VDD.n4453 VDD.n389 146.341
R3500 VDD.n4453 VDD.n381 146.341
R3501 VDD.n4463 VDD.n381 146.341
R3502 VDD.n4464 VDD.n4463 146.341
R3503 VDD.n4464 VDD.n377 146.341
R3504 VDD.n4473 VDD.n377 146.341
R3505 VDD.n4473 VDD.n369 146.341
R3506 VDD.n4485 VDD.n369 146.341
R3507 VDD.n4486 VDD.n4485 146.341
R3508 VDD.n4486 VDD.n43 146.341
R3509 VDD.n44 VDD.n43 146.341
R3510 VDD.n45 VDD.n44 146.341
R3511 VDD.n4493 VDD.n45 146.341
R3512 VDD.n4493 VDD.n54 146.341
R3513 VDD.n55 VDD.n54 146.341
R3514 VDD.n56 VDD.n55 146.341
R3515 VDD.n4500 VDD.n56 146.341
R3516 VDD.n4500 VDD.n65 146.341
R3517 VDD.n66 VDD.n65 146.341
R3518 VDD.n67 VDD.n66 146.341
R3519 VDD.n4507 VDD.n67 146.341
R3520 VDD.n4507 VDD.n76 146.341
R3521 VDD.n77 VDD.n76 146.341
R3522 VDD.n78 VDD.n77 146.341
R3523 VDD.n4514 VDD.n78 146.341
R3524 VDD.n4514 VDD.n87 146.341
R3525 VDD.n88 VDD.n87 146.341
R3526 VDD.n89 VDD.n88 146.341
R3527 VDD.n4521 VDD.n89 146.341
R3528 VDD.n4521 VDD.n98 146.341
R3529 VDD.n99 VDD.n98 146.341
R3530 VDD.n100 VDD.n99 146.341
R3531 VDD.n4528 VDD.n100 146.341
R3532 VDD.n4528 VDD.n109 146.341
R3533 VDD.n110 VDD.n109 146.341
R3534 VDD.n111 VDD.n110 146.341
R3535 VDD.n4535 VDD.n111 146.341
R3536 VDD.n4535 VDD.n120 146.341
R3537 VDD.n121 VDD.n120 146.341
R3538 VDD.n122 VDD.n121 146.341
R3539 VDD.n4542 VDD.n122 146.341
R3540 VDD.n4542 VDD.n131 146.341
R3541 VDD.n132 VDD.n131 146.341
R3542 VDD.n133 VDD.n132 146.341
R3543 VDD.n4549 VDD.n133 146.341
R3544 VDD.n4549 VDD.n142 146.341
R3545 VDD.n143 VDD.n142 146.341
R3546 VDD.n144 VDD.n143 146.341
R3547 VDD.n4556 VDD.n144 146.341
R3548 VDD.n4556 VDD.n153 146.341
R3549 VDD.n154 VDD.n153 146.341
R3550 VDD.n155 VDD.n154 146.341
R3551 VDD.n4563 VDD.n155 146.341
R3552 VDD.n4563 VDD.n164 146.341
R3553 VDD.n165 VDD.n164 146.341
R3554 VDD.n166 VDD.n165 146.341
R3555 VDD.n4570 VDD.n166 146.341
R3556 VDD.n4570 VDD.n175 146.341
R3557 VDD.n176 VDD.n175 146.341
R3558 VDD.n177 VDD.n176 146.341
R3559 VDD.n4577 VDD.n177 146.341
R3560 VDD.n4577 VDD.n186 146.341
R3561 VDD.n187 VDD.n186 146.341
R3562 VDD.n188 VDD.n187 146.341
R3563 VDD.n4584 VDD.n188 146.341
R3564 VDD.n4584 VDD.n197 146.341
R3565 VDD.n198 VDD.n197 146.341
R3566 VDD.n4244 VDD.n546 146.341
R3567 VDD.n591 VDD.n546 146.341
R3568 VDD.n594 VDD.n593 146.341
R3569 VDD.n601 VDD.n600 146.341
R3570 VDD.n604 VDD.n603 146.341
R3571 VDD.n611 VDD.n610 146.341
R3572 VDD.n614 VDD.n613 146.341
R3573 VDD.n621 VDD.n620 146.341
R3574 VDD.n624 VDD.n623 146.341
R3575 VDD.n631 VDD.n630 146.341
R3576 VDD.n634 VDD.n633 146.341
R3577 VDD.n641 VDD.n640 146.341
R3578 VDD.n645 VDD.n644 146.341
R3579 VDD.n652 VDD.n651 146.341
R3580 VDD.n655 VDD.n654 146.341
R3581 VDD.n662 VDD.n661 146.341
R3582 VDD.n665 VDD.n664 146.341
R3583 VDD.n672 VDD.n671 146.341
R3584 VDD.n4241 VDD.n564 146.341
R3585 VDD.n4251 VDD.n539 146.341
R3586 VDD.n4251 VDD.n531 146.341
R3587 VDD.n4261 VDD.n531 146.341
R3588 VDD.n4261 VDD.n527 146.341
R3589 VDD.n4267 VDD.n527 146.341
R3590 VDD.n4267 VDD.n519 146.341
R3591 VDD.n4277 VDD.n519 146.341
R3592 VDD.n4277 VDD.n515 146.341
R3593 VDD.n4283 VDD.n515 146.341
R3594 VDD.n4283 VDD.n507 146.341
R3595 VDD.n4293 VDD.n507 146.341
R3596 VDD.n4293 VDD.n503 146.341
R3597 VDD.n4299 VDD.n503 146.341
R3598 VDD.n4299 VDD.n495 146.341
R3599 VDD.n4309 VDD.n495 146.341
R3600 VDD.n4309 VDD.n491 146.341
R3601 VDD.n4315 VDD.n491 146.341
R3602 VDD.n4315 VDD.n483 146.341
R3603 VDD.n4325 VDD.n483 146.341
R3604 VDD.n4325 VDD.n479 146.341
R3605 VDD.n4331 VDD.n479 146.341
R3606 VDD.n4331 VDD.n471 146.341
R3607 VDD.n4341 VDD.n471 146.341
R3608 VDD.n4341 VDD.n467 146.341
R3609 VDD.n4347 VDD.n467 146.341
R3610 VDD.n4347 VDD.n459 146.341
R3611 VDD.n4357 VDD.n459 146.341
R3612 VDD.n4357 VDD.n455 146.341
R3613 VDD.n4363 VDD.n455 146.341
R3614 VDD.n4363 VDD.n447 146.341
R3615 VDD.n4373 VDD.n447 146.341
R3616 VDD.n4373 VDD.n443 146.341
R3617 VDD.n4379 VDD.n443 146.341
R3618 VDD.n4379 VDD.n435 146.341
R3619 VDD.n4389 VDD.n435 146.341
R3620 VDD.n4389 VDD.n431 146.341
R3621 VDD.n4395 VDD.n431 146.341
R3622 VDD.n4395 VDD.n423 146.341
R3623 VDD.n4405 VDD.n423 146.341
R3624 VDD.n4405 VDD.n419 146.341
R3625 VDD.n4411 VDD.n419 146.341
R3626 VDD.n4411 VDD.n411 146.341
R3627 VDD.n4421 VDD.n411 146.341
R3628 VDD.n4421 VDD.n407 146.341
R3629 VDD.n4427 VDD.n407 146.341
R3630 VDD.n4427 VDD.n399 146.341
R3631 VDD.n4437 VDD.n399 146.341
R3632 VDD.n4437 VDD.n395 146.341
R3633 VDD.n4443 VDD.n395 146.341
R3634 VDD.n4443 VDD.n387 146.341
R3635 VDD.n4455 VDD.n387 146.341
R3636 VDD.n4455 VDD.n383 146.341
R3637 VDD.n4461 VDD.n383 146.341
R3638 VDD.n4461 VDD.n375 146.341
R3639 VDD.n4476 VDD.n375 146.341
R3640 VDD.n4476 VDD.n371 146.341
R3641 VDD.n4482 VDD.n371 146.341
R3642 VDD.n4483 VDD.n4482 146.341
R3643 VDD.n4483 VDD.n39 146.341
R3644 VDD.n4708 VDD.n39 146.341
R3645 VDD.n4708 VDD.n41 146.341
R3646 VDD.n4704 VDD.n41 146.341
R3647 VDD.n4704 VDD.n47 146.341
R3648 VDD.n4700 VDD.n47 146.341
R3649 VDD.n4700 VDD.n53 146.341
R3650 VDD.n4696 VDD.n53 146.341
R3651 VDD.n4696 VDD.n58 146.341
R3652 VDD.n4692 VDD.n58 146.341
R3653 VDD.n4692 VDD.n64 146.341
R3654 VDD.n4688 VDD.n64 146.341
R3655 VDD.n4688 VDD.n68 146.341
R3656 VDD.n4684 VDD.n68 146.341
R3657 VDD.n4684 VDD.n74 146.341
R3658 VDD.n4680 VDD.n74 146.341
R3659 VDD.n4680 VDD.n80 146.341
R3660 VDD.n4676 VDD.n80 146.341
R3661 VDD.n4676 VDD.n86 146.341
R3662 VDD.n4672 VDD.n86 146.341
R3663 VDD.n4672 VDD.n91 146.341
R3664 VDD.n4668 VDD.n91 146.341
R3665 VDD.n4668 VDD.n97 146.341
R3666 VDD.n4664 VDD.n97 146.341
R3667 VDD.n4664 VDD.n102 146.341
R3668 VDD.n4660 VDD.n102 146.341
R3669 VDD.n4660 VDD.n108 146.341
R3670 VDD.n4656 VDD.n108 146.341
R3671 VDD.n4656 VDD.n113 146.341
R3672 VDD.n4652 VDD.n113 146.341
R3673 VDD.n4652 VDD.n119 146.341
R3674 VDD.n4648 VDD.n119 146.341
R3675 VDD.n4648 VDD.n124 146.341
R3676 VDD.n4644 VDD.n124 146.341
R3677 VDD.n4644 VDD.n130 146.341
R3678 VDD.n4640 VDD.n130 146.341
R3679 VDD.n4640 VDD.n135 146.341
R3680 VDD.n4636 VDD.n135 146.341
R3681 VDD.n4636 VDD.n141 146.341
R3682 VDD.n4632 VDD.n141 146.341
R3683 VDD.n4632 VDD.n146 146.341
R3684 VDD.n4628 VDD.n146 146.341
R3685 VDD.n4628 VDD.n152 146.341
R3686 VDD.n4624 VDD.n152 146.341
R3687 VDD.n4624 VDD.n157 146.341
R3688 VDD.n4620 VDD.n157 146.341
R3689 VDD.n4620 VDD.n163 146.341
R3690 VDD.n4616 VDD.n163 146.341
R3691 VDD.n4616 VDD.n168 146.341
R3692 VDD.n4612 VDD.n168 146.341
R3693 VDD.n4612 VDD.n174 146.341
R3694 VDD.n4608 VDD.n174 146.341
R3695 VDD.n4608 VDD.n178 146.341
R3696 VDD.n4604 VDD.n178 146.341
R3697 VDD.n4604 VDD.n184 146.341
R3698 VDD.n4600 VDD.n184 146.341
R3699 VDD.n4600 VDD.n190 146.341
R3700 VDD.n4596 VDD.n190 146.341
R3701 VDD.n4596 VDD.n196 146.341
R3702 VDD.n2849 VDD.n2848 146.341
R3703 VDD.n2852 VDD.n2851 146.341
R3704 VDD.n2859 VDD.n2858 146.341
R3705 VDD.n2862 VDD.n2861 146.341
R3706 VDD.n2869 VDD.n2868 146.341
R3707 VDD.n2875 VDD.n2874 146.341
R3708 VDD.n2882 VDD.n2881 146.341
R3709 VDD.n2885 VDD.n2884 146.341
R3710 VDD.n2892 VDD.n2891 146.341
R3711 VDD.n1809 VDD.n1808 146.341
R3712 VDD.n2895 VDD.n1810 146.341
R3713 VDD.n1816 VDD.n1813 146.341
R3714 VDD.n2898 VDD.n1817 146.341
R3715 VDD.n1821 VDD.n1820 146.341
R3716 VDD.n2901 VDD.n1822 146.341
R3717 VDD.n1826 VDD.n1825 146.341
R3718 VDD.n2904 VDD.n1827 146.341
R3719 VDD.n1831 VDD.n1830 146.341
R3720 VDD.n2374 VDD.n2223 146.341
R3721 VDD.n2374 VDD.n2219 146.341
R3722 VDD.n2380 VDD.n2219 146.341
R3723 VDD.n2380 VDD.n2210 146.341
R3724 VDD.n2390 VDD.n2210 146.341
R3725 VDD.n2390 VDD.n2206 146.341
R3726 VDD.n2396 VDD.n2206 146.341
R3727 VDD.n2396 VDD.n2199 146.341
R3728 VDD.n2406 VDD.n2199 146.341
R3729 VDD.n2406 VDD.n2195 146.341
R3730 VDD.n2412 VDD.n2195 146.341
R3731 VDD.n2412 VDD.n2187 146.341
R3732 VDD.n2422 VDD.n2187 146.341
R3733 VDD.n2422 VDD.n2183 146.341
R3734 VDD.n2428 VDD.n2183 146.341
R3735 VDD.n2428 VDD.n2175 146.341
R3736 VDD.n2438 VDD.n2175 146.341
R3737 VDD.n2438 VDD.n2171 146.341
R3738 VDD.n2444 VDD.n2171 146.341
R3739 VDD.n2444 VDD.n2163 146.341
R3740 VDD.n2454 VDD.n2163 146.341
R3741 VDD.n2454 VDD.n2159 146.341
R3742 VDD.n2460 VDD.n2159 146.341
R3743 VDD.n2460 VDD.n2151 146.341
R3744 VDD.n2470 VDD.n2151 146.341
R3745 VDD.n2470 VDD.n2147 146.341
R3746 VDD.n2476 VDD.n2147 146.341
R3747 VDD.n2476 VDD.n2139 146.341
R3748 VDD.n2486 VDD.n2139 146.341
R3749 VDD.n2486 VDD.n2135 146.341
R3750 VDD.n2492 VDD.n2135 146.341
R3751 VDD.n2492 VDD.n2127 146.341
R3752 VDD.n2502 VDD.n2127 146.341
R3753 VDD.n2502 VDD.n2123 146.341
R3754 VDD.n2508 VDD.n2123 146.341
R3755 VDD.n2508 VDD.n2115 146.341
R3756 VDD.n2518 VDD.n2115 146.341
R3757 VDD.n2518 VDD.n2111 146.341
R3758 VDD.n2524 VDD.n2111 146.341
R3759 VDD.n2524 VDD.n2103 146.341
R3760 VDD.n2534 VDD.n2103 146.341
R3761 VDD.n2534 VDD.n2099 146.341
R3762 VDD.n2540 VDD.n2099 146.341
R3763 VDD.n2540 VDD.n2090 146.341
R3764 VDD.n2550 VDD.n2090 146.341
R3765 VDD.n2550 VDD.n2086 146.341
R3766 VDD.n2556 VDD.n2086 146.341
R3767 VDD.n2556 VDD.n2079 146.341
R3768 VDD.n2566 VDD.n2079 146.341
R3769 VDD.n2566 VDD.n2075 146.341
R3770 VDD.n2572 VDD.n2075 146.341
R3771 VDD.n2572 VDD.n2067 146.341
R3772 VDD.n2582 VDD.n2067 146.341
R3773 VDD.n2582 VDD.n2063 146.341
R3774 VDD.n2588 VDD.n2063 146.341
R3775 VDD.n2588 VDD.n2054 146.341
R3776 VDD.n2599 VDD.n2054 146.341
R3777 VDD.n2599 VDD.n2050 146.341
R3778 VDD.n2605 VDD.n2050 146.341
R3779 VDD.n2605 VDD.n2022 146.341
R3780 VDD.n2615 VDD.n2022 146.341
R3781 VDD.n2615 VDD.n2018 146.341
R3782 VDD.n2621 VDD.n2018 146.341
R3783 VDD.n2621 VDD.n2010 146.341
R3784 VDD.n2631 VDD.n2010 146.341
R3785 VDD.n2631 VDD.n2006 146.341
R3786 VDD.n2637 VDD.n2006 146.341
R3787 VDD.n2637 VDD.n1997 146.341
R3788 VDD.n2647 VDD.n1997 146.341
R3789 VDD.n2647 VDD.n1993 146.341
R3790 VDD.n2653 VDD.n1993 146.341
R3791 VDD.n2653 VDD.n1986 146.341
R3792 VDD.n2663 VDD.n1986 146.341
R3793 VDD.n2663 VDD.n1982 146.341
R3794 VDD.n2669 VDD.n1982 146.341
R3795 VDD.n2669 VDD.n1974 146.341
R3796 VDD.n2679 VDD.n1974 146.341
R3797 VDD.n2679 VDD.n1970 146.341
R3798 VDD.n2685 VDD.n1970 146.341
R3799 VDD.n2685 VDD.n1962 146.341
R3800 VDD.n2695 VDD.n1962 146.341
R3801 VDD.n2695 VDD.n1958 146.341
R3802 VDD.n2701 VDD.n1958 146.341
R3803 VDD.n2701 VDD.n1950 146.341
R3804 VDD.n2711 VDD.n1950 146.341
R3805 VDD.n2711 VDD.n1946 146.341
R3806 VDD.n2717 VDD.n1946 146.341
R3807 VDD.n2717 VDD.n1938 146.341
R3808 VDD.n2727 VDD.n1938 146.341
R3809 VDD.n2727 VDD.n1934 146.341
R3810 VDD.n2733 VDD.n1934 146.341
R3811 VDD.n2733 VDD.n1926 146.341
R3812 VDD.n2743 VDD.n1926 146.341
R3813 VDD.n2743 VDD.n1922 146.341
R3814 VDD.n2749 VDD.n1922 146.341
R3815 VDD.n2749 VDD.n1914 146.341
R3816 VDD.n2759 VDD.n1914 146.341
R3817 VDD.n2759 VDD.n1910 146.341
R3818 VDD.n2765 VDD.n1910 146.341
R3819 VDD.n2765 VDD.n1902 146.341
R3820 VDD.n2775 VDD.n1902 146.341
R3821 VDD.n2775 VDD.n1898 146.341
R3822 VDD.n2781 VDD.n1898 146.341
R3823 VDD.n2781 VDD.n1890 146.341
R3824 VDD.n2791 VDD.n1890 146.341
R3825 VDD.n2791 VDD.n1886 146.341
R3826 VDD.n2797 VDD.n1886 146.341
R3827 VDD.n2797 VDD.n1877 146.341
R3828 VDD.n2807 VDD.n1877 146.341
R3829 VDD.n2807 VDD.n1872 146.341
R3830 VDD.n2814 VDD.n1872 146.341
R3831 VDD.n2814 VDD.n1865 146.341
R3832 VDD.n2824 VDD.n1865 146.341
R3833 VDD.n2825 VDD.n2824 146.341
R3834 VDD.n2825 VDD.n1860 146.341
R3835 VDD.n2833 VDD.n1860 146.341
R3836 VDD.n2833 VDD.n1835 146.341
R3837 VDD.n2363 VDD.n2229 146.341
R3838 VDD.n2363 VDD.n2248 146.341
R3839 VDD.n2252 VDD.n2251 146.341
R3840 VDD.n2254 VDD.n2253 146.341
R3841 VDD.n2258 VDD.n2257 146.341
R3842 VDD.n2264 VDD.n2259 146.341
R3843 VDD.n2266 VDD.n2265 146.341
R3844 VDD.n2270 VDD.n2269 146.341
R3845 VDD.n2272 VDD.n2271 146.341
R3846 VDD.n2276 VDD.n2275 146.341
R3847 VDD.n2278 VDD.n2277 146.341
R3848 VDD.n2282 VDD.n2281 146.341
R3849 VDD.n2284 VDD.n2283 146.341
R3850 VDD.n2288 VDD.n2287 146.341
R3851 VDD.n2290 VDD.n2289 146.341
R3852 VDD.n2294 VDD.n2293 146.341
R3853 VDD.n2296 VDD.n2295 146.341
R3854 VDD.n2300 VDD.n2299 146.341
R3855 VDD.n2301 VDD.n2247 146.341
R3856 VDD.n2372 VDD.n2225 146.341
R3857 VDD.n2372 VDD.n2217 146.341
R3858 VDD.n2382 VDD.n2217 146.341
R3859 VDD.n2382 VDD.n2213 146.341
R3860 VDD.n2388 VDD.n2213 146.341
R3861 VDD.n2388 VDD.n2205 146.341
R3862 VDD.n2398 VDD.n2205 146.341
R3863 VDD.n2398 VDD.n2201 146.341
R3864 VDD.n2404 VDD.n2201 146.341
R3865 VDD.n2404 VDD.n2193 146.341
R3866 VDD.n2414 VDD.n2193 146.341
R3867 VDD.n2414 VDD.n2189 146.341
R3868 VDD.n2420 VDD.n2189 146.341
R3869 VDD.n2420 VDD.n2181 146.341
R3870 VDD.n2430 VDD.n2181 146.341
R3871 VDD.n2430 VDD.n2177 146.341
R3872 VDD.n2436 VDD.n2177 146.341
R3873 VDD.n2436 VDD.n2169 146.341
R3874 VDD.n2446 VDD.n2169 146.341
R3875 VDD.n2446 VDD.n2165 146.341
R3876 VDD.n2452 VDD.n2165 146.341
R3877 VDD.n2452 VDD.n2157 146.341
R3878 VDD.n2462 VDD.n2157 146.341
R3879 VDD.n2462 VDD.n2153 146.341
R3880 VDD.n2468 VDD.n2153 146.341
R3881 VDD.n2468 VDD.n2145 146.341
R3882 VDD.n2478 VDD.n2145 146.341
R3883 VDD.n2478 VDD.n2141 146.341
R3884 VDD.n2484 VDD.n2141 146.341
R3885 VDD.n2484 VDD.n2133 146.341
R3886 VDD.n2494 VDD.n2133 146.341
R3887 VDD.n2494 VDD.n2129 146.341
R3888 VDD.n2500 VDD.n2129 146.341
R3889 VDD.n2500 VDD.n2121 146.341
R3890 VDD.n2510 VDD.n2121 146.341
R3891 VDD.n2510 VDD.n2117 146.341
R3892 VDD.n2516 VDD.n2117 146.341
R3893 VDD.n2516 VDD.n2109 146.341
R3894 VDD.n2526 VDD.n2109 146.341
R3895 VDD.n2526 VDD.n2105 146.341
R3896 VDD.n2532 VDD.n2105 146.341
R3897 VDD.n2532 VDD.n2097 146.341
R3898 VDD.n2542 VDD.n2097 146.341
R3899 VDD.n2542 VDD.n2093 146.341
R3900 VDD.n2548 VDD.n2093 146.341
R3901 VDD.n2548 VDD.n2085 146.341
R3902 VDD.n2558 VDD.n2085 146.341
R3903 VDD.n2558 VDD.n2081 146.341
R3904 VDD.n2564 VDD.n2081 146.341
R3905 VDD.n2564 VDD.n2073 146.341
R3906 VDD.n2574 VDD.n2073 146.341
R3907 VDD.n2574 VDD.n2069 146.341
R3908 VDD.n2580 VDD.n2069 146.341
R3909 VDD.n2580 VDD.n2061 146.341
R3910 VDD.n2590 VDD.n2061 146.341
R3911 VDD.n2590 VDD.n2057 146.341
R3912 VDD.n2597 VDD.n2057 146.341
R3913 VDD.n2597 VDD.n2049 146.341
R3914 VDD.n2607 VDD.n2049 146.341
R3915 VDD.n2607 VDD.n2024 146.341
R3916 VDD.n2613 VDD.n2024 146.341
R3917 VDD.n2613 VDD.n2016 146.341
R3918 VDD.n2623 VDD.n2016 146.341
R3919 VDD.n2623 VDD.n2012 146.341
R3920 VDD.n2629 VDD.n2012 146.341
R3921 VDD.n2629 VDD.n2004 146.341
R3922 VDD.n2639 VDD.n2004 146.341
R3923 VDD.n2639 VDD.n2000 146.341
R3924 VDD.n2645 VDD.n2000 146.341
R3925 VDD.n2645 VDD.n1992 146.341
R3926 VDD.n2655 VDD.n1992 146.341
R3927 VDD.n2655 VDD.n1988 146.341
R3928 VDD.n2661 VDD.n1988 146.341
R3929 VDD.n2661 VDD.n1980 146.341
R3930 VDD.n2671 VDD.n1980 146.341
R3931 VDD.n2671 VDD.n1976 146.341
R3932 VDD.n2677 VDD.n1976 146.341
R3933 VDD.n2677 VDD.n1968 146.341
R3934 VDD.n2687 VDD.n1968 146.341
R3935 VDD.n2687 VDD.n1964 146.341
R3936 VDD.n2693 VDD.n1964 146.341
R3937 VDD.n2693 VDD.n1956 146.341
R3938 VDD.n2703 VDD.n1956 146.341
R3939 VDD.n2703 VDD.n1952 146.341
R3940 VDD.n2709 VDD.n1952 146.341
R3941 VDD.n2709 VDD.n1944 146.341
R3942 VDD.n2719 VDD.n1944 146.341
R3943 VDD.n2719 VDD.n1940 146.341
R3944 VDD.n2725 VDD.n1940 146.341
R3945 VDD.n2725 VDD.n1932 146.341
R3946 VDD.n2735 VDD.n1932 146.341
R3947 VDD.n2735 VDD.n1928 146.341
R3948 VDD.n2741 VDD.n1928 146.341
R3949 VDD.n2741 VDD.n1920 146.341
R3950 VDD.n2751 VDD.n1920 146.341
R3951 VDD.n2751 VDD.n1916 146.341
R3952 VDD.n2757 VDD.n1916 146.341
R3953 VDD.n2757 VDD.n1908 146.341
R3954 VDD.n2767 VDD.n1908 146.341
R3955 VDD.n2767 VDD.n1904 146.341
R3956 VDD.n2773 VDD.n1904 146.341
R3957 VDD.n2773 VDD.n1896 146.341
R3958 VDD.n2783 VDD.n1896 146.341
R3959 VDD.n2783 VDD.n1892 146.341
R3960 VDD.n2789 VDD.n1892 146.341
R3961 VDD.n2789 VDD.n1884 146.341
R3962 VDD.n2799 VDD.n1884 146.341
R3963 VDD.n2799 VDD.n1880 146.341
R3964 VDD.n2805 VDD.n1880 146.341
R3965 VDD.n2805 VDD.n1871 146.341
R3966 VDD.n2816 VDD.n1871 146.341
R3967 VDD.n2816 VDD.n1867 146.341
R3968 VDD.n2822 VDD.n1867 146.341
R3969 VDD.n2822 VDD.n1858 146.341
R3970 VDD.n2836 VDD.n1858 146.341
R3971 VDD.n2836 VDD.n1854 146.341
R3972 VDD.n2842 VDD.n1854 146.341
R3973 VDD.n2040 VDD.t144 126.526
R3974 VDD.n2033 VDD.t113 126.526
R3975 VDD.n2027 VDD.t116 126.526
R3976 VDD.n34 VDD.t152 124.76
R3977 VDD.n27 VDD.t105 124.76
R3978 VDD.n21 VDD.t106 124.76
R3979 VDD.n2305 VDD.t60 122.692
R3980 VDD.n2327 VDD.t57 122.692
R3981 VDD.n2261 VDD.t34 122.692
R3982 VDD.n566 VDD.t54 122.692
R3983 VDD.n576 VDD.t51 122.692
R3984 VDD.n584 VDD.t30 122.692
R3985 VDD.n219 VDD.t14 122.692
R3986 VDD.n229 VDD.t11 122.692
R3987 VDD.n238 VDD.t20 122.692
R3988 VDD.n2872 VDD.t38 122.692
R3989 VDD.n1815 VDD.t24 122.692
R3990 VDD.n1833 VDD.t27 122.692
R3991 VDD.n3386 VDD.n3385 117.778
R3992 VDD.n3610 VDD.n3609 115.977
R3993 VDD.n710 VDD.n709 115.977
R3994 VDD.n3392 VDD.n3391 115.977
R3995 VDD.n685 VDD.n684 115.977
R3996 VDD.n1410 VDD.n1409 115.977
R3997 VDD.n1062 VDD.n1061 115.977
R3998 VDD.n1624 VDD.n1623 115.977
R3999 VDD.n1080 VDD.n1079 115.977
R4000 VDD.n9 VDD.n7 111.183
R4001 VDD.n2 VDD.n0 111.183
R4002 VDD.n9 VDD.n8 109.275
R4003 VDD.n11 VDD.n10 109.275
R4004 VDD.n13 VDD.n12 109.275
R4005 VDD.n6 VDD.n5 109.275
R4006 VDD.n4 VDD.n3 109.275
R4007 VDD.n2 VDD.n1 109.275
R4008 VDD.n3610 VDD.t64 108.311
R4009 VDD.n710 VDD.t42 108.311
R4010 VDD.n3392 VDD.t67 108.311
R4011 VDD.n685 VDD.t49 108.311
R4012 VDD.n1410 VDD.t16 108.311
R4013 VDD.n1062 VDD.t46 108.311
R4014 VDD.n1624 VDD.t6 108.311
R4015 VDD.n1080 VDD.t71 108.311
R4016 VDD.n2305 VDD.n2304 106.474
R4017 VDD.n2327 VDD.n2326 106.474
R4018 VDD.n2261 VDD.n2260 106.474
R4019 VDD.n566 VDD.n565 106.474
R4020 VDD.n576 VDD.n575 106.474
R4021 VDD.n584 VDD.n583 106.474
R4022 VDD.n219 VDD.n218 106.474
R4023 VDD.n229 VDD.n228 106.474
R4024 VDD.n238 VDD.n237 106.474
R4025 VDD.n2872 VDD.n2871 106.474
R4026 VDD.n1815 VDD.n1814 106.474
R4027 VDD.n1833 VDD.n1832 106.474
R4028 VDD.n31 VDD.n29 105.35
R4029 VDD.n24 VDD.n22 105.35
R4030 VDD.n18 VDD.n16 105.35
R4031 VDD.n33 VDD.n32 103.584
R4032 VDD.n31 VDD.n30 103.584
R4033 VDD.n26 VDD.n25 103.584
R4034 VDD.n24 VDD.n23 103.584
R4035 VDD.n20 VDD.n19 103.584
R4036 VDD.n18 VDD.n17 103.584
R4037 VDD.n2040 VDD.n2039 103.584
R4038 VDD.n2042 VDD.n2041 103.584
R4039 VDD.n2044 VDD.n2043 103.584
R4040 VDD.n2033 VDD.n2032 103.584
R4041 VDD.n2035 VDD.n2034 103.584
R4042 VDD.n2037 VDD.n2036 103.584
R4043 VDD.n2027 VDD.n2026 103.584
R4044 VDD.n2029 VDD.n2028 103.584
R4045 VDD.n2031 VDD.n2030 103.584
R4046 VDD.t89 VDD.n1397 103.014
R4047 VDD.n679 VDD.t0 103.014
R4048 VDD.n3818 VDD.n1033 99.5127
R4049 VDD.n3822 VDD.n1033 99.5127
R4050 VDD.n3822 VDD.n1023 99.5127
R4051 VDD.n3830 VDD.n1023 99.5127
R4052 VDD.n3830 VDD.n1021 99.5127
R4053 VDD.n3834 VDD.n1021 99.5127
R4054 VDD.n3834 VDD.n1011 99.5127
R4055 VDD.n3842 VDD.n1011 99.5127
R4056 VDD.n3842 VDD.n1009 99.5127
R4057 VDD.n3846 VDD.n1009 99.5127
R4058 VDD.n3846 VDD.n998 99.5127
R4059 VDD.n3854 VDD.n998 99.5127
R4060 VDD.n3854 VDD.n996 99.5127
R4061 VDD.n3858 VDD.n996 99.5127
R4062 VDD.n3858 VDD.n987 99.5127
R4063 VDD.n3866 VDD.n987 99.5127
R4064 VDD.n3866 VDD.n985 99.5127
R4065 VDD.n3870 VDD.n985 99.5127
R4066 VDD.n3870 VDD.n975 99.5127
R4067 VDD.n3878 VDD.n975 99.5127
R4068 VDD.n3878 VDD.n973 99.5127
R4069 VDD.n3882 VDD.n973 99.5127
R4070 VDD.n3882 VDD.n963 99.5127
R4071 VDD.n3890 VDD.n963 99.5127
R4072 VDD.n3890 VDD.n961 99.5127
R4073 VDD.n3894 VDD.n961 99.5127
R4074 VDD.n3894 VDD.n951 99.5127
R4075 VDD.n3902 VDD.n951 99.5127
R4076 VDD.n3902 VDD.n949 99.5127
R4077 VDD.n3906 VDD.n949 99.5127
R4078 VDD.n3906 VDD.n939 99.5127
R4079 VDD.n3914 VDD.n939 99.5127
R4080 VDD.n3914 VDD.n937 99.5127
R4081 VDD.n3918 VDD.n937 99.5127
R4082 VDD.n3918 VDD.n927 99.5127
R4083 VDD.n3926 VDD.n927 99.5127
R4084 VDD.n3926 VDD.n925 99.5127
R4085 VDD.n3930 VDD.n925 99.5127
R4086 VDD.n3930 VDD.n915 99.5127
R4087 VDD.n3938 VDD.n915 99.5127
R4088 VDD.n3938 VDD.n913 99.5127
R4089 VDD.n3942 VDD.n913 99.5127
R4090 VDD.n3942 VDD.n903 99.5127
R4091 VDD.n3950 VDD.n903 99.5127
R4092 VDD.n3950 VDD.n901 99.5127
R4093 VDD.n3954 VDD.n901 99.5127
R4094 VDD.n3954 VDD.n891 99.5127
R4095 VDD.n3962 VDD.n891 99.5127
R4096 VDD.n3962 VDD.n889 99.5127
R4097 VDD.n3966 VDD.n889 99.5127
R4098 VDD.n3966 VDD.n879 99.5127
R4099 VDD.n3974 VDD.n879 99.5127
R4100 VDD.n3974 VDD.n877 99.5127
R4101 VDD.n3978 VDD.n877 99.5127
R4102 VDD.n3978 VDD.n867 99.5127
R4103 VDD.n3986 VDD.n867 99.5127
R4104 VDD.n3986 VDD.n865 99.5127
R4105 VDD.n3990 VDD.n865 99.5127
R4106 VDD.n3990 VDD.n855 99.5127
R4107 VDD.n3998 VDD.n855 99.5127
R4108 VDD.n3998 VDD.n853 99.5127
R4109 VDD.n4002 VDD.n853 99.5127
R4110 VDD.n4002 VDD.n843 99.5127
R4111 VDD.n4010 VDD.n843 99.5127
R4112 VDD.n4010 VDD.n841 99.5127
R4113 VDD.n4014 VDD.n841 99.5127
R4114 VDD.n4014 VDD.n831 99.5127
R4115 VDD.n4022 VDD.n831 99.5127
R4116 VDD.n4022 VDD.n829 99.5127
R4117 VDD.n4026 VDD.n829 99.5127
R4118 VDD.n4026 VDD.n819 99.5127
R4119 VDD.n4034 VDD.n819 99.5127
R4120 VDD.n4034 VDD.n817 99.5127
R4121 VDD.n4038 VDD.n817 99.5127
R4122 VDD.n4038 VDD.n807 99.5127
R4123 VDD.n4046 VDD.n807 99.5127
R4124 VDD.n4046 VDD.n805 99.5127
R4125 VDD.n4050 VDD.n805 99.5127
R4126 VDD.n4050 VDD.n795 99.5127
R4127 VDD.n4058 VDD.n795 99.5127
R4128 VDD.n4058 VDD.n793 99.5127
R4129 VDD.n4062 VDD.n793 99.5127
R4130 VDD.n4062 VDD.n783 99.5127
R4131 VDD.n4070 VDD.n783 99.5127
R4132 VDD.n4070 VDD.n781 99.5127
R4133 VDD.n4074 VDD.n781 99.5127
R4134 VDD.n4074 VDD.n771 99.5127
R4135 VDD.n4082 VDD.n771 99.5127
R4136 VDD.n4082 VDD.n769 99.5127
R4137 VDD.n4086 VDD.n769 99.5127
R4138 VDD.n4086 VDD.n759 99.5127
R4139 VDD.n4094 VDD.n759 99.5127
R4140 VDD.n4094 VDD.n757 99.5127
R4141 VDD.n4098 VDD.n757 99.5127
R4142 VDD.n4098 VDD.n746 99.5127
R4143 VDD.n4106 VDD.n746 99.5127
R4144 VDD.n4106 VDD.n744 99.5127
R4145 VDD.n4110 VDD.n744 99.5127
R4146 VDD.n4110 VDD.n735 99.5127
R4147 VDD.n4118 VDD.n735 99.5127
R4148 VDD.n4118 VDD.n733 99.5127
R4149 VDD.n4122 VDD.n733 99.5127
R4150 VDD.n4122 VDD.n722 99.5127
R4151 VDD.n4160 VDD.n722 99.5127
R4152 VDD.n4160 VDD.n720 99.5127
R4153 VDD.n4164 VDD.n720 99.5127
R4154 VDD.n4164 VDD.n695 99.5127
R4155 VDD.n4212 VDD.n695 99.5127
R4156 VDD.n4212 VDD.n696 99.5127
R4157 VDD.n4208 VDD.n4207 99.5127
R4158 VDD.n4205 VDD.n699 99.5127
R4159 VDD.n4201 VDD.n4200 99.5127
R4160 VDD.n4198 VDD.n702 99.5127
R4161 VDD.n4194 VDD.n4193 99.5127
R4162 VDD.n4191 VDD.n705 99.5127
R4163 VDD.n4187 VDD.n4186 99.5127
R4164 VDD.n4184 VDD.n708 99.5127
R4165 VDD.n4180 VDD.n4179 99.5127
R4166 VDD.n4177 VDD.n714 99.5127
R4167 VDD.n3598 VDD.n3388 99.5127
R4168 VDD.n3388 VDD.n1031 99.5127
R4169 VDD.n3593 VDD.n1031 99.5127
R4170 VDD.n3593 VDD.n1025 99.5127
R4171 VDD.n3590 VDD.n1025 99.5127
R4172 VDD.n3590 VDD.n1019 99.5127
R4173 VDD.n3587 VDD.n1019 99.5127
R4174 VDD.n3587 VDD.n1013 99.5127
R4175 VDD.n3584 VDD.n1013 99.5127
R4176 VDD.n3584 VDD.n1006 99.5127
R4177 VDD.n3581 VDD.n1006 99.5127
R4178 VDD.n3581 VDD.n999 99.5127
R4179 VDD.n3578 VDD.n999 99.5127
R4180 VDD.n3578 VDD.n994 99.5127
R4181 VDD.n3575 VDD.n994 99.5127
R4182 VDD.n3575 VDD.n989 99.5127
R4183 VDD.n3572 VDD.n989 99.5127
R4184 VDD.n3572 VDD.n983 99.5127
R4185 VDD.n3569 VDD.n983 99.5127
R4186 VDD.n3569 VDD.n977 99.5127
R4187 VDD.n3566 VDD.n977 99.5127
R4188 VDD.n3566 VDD.n971 99.5127
R4189 VDD.n3563 VDD.n971 99.5127
R4190 VDD.n3563 VDD.n965 99.5127
R4191 VDD.n3560 VDD.n965 99.5127
R4192 VDD.n3560 VDD.n959 99.5127
R4193 VDD.n3557 VDD.n959 99.5127
R4194 VDD.n3557 VDD.n953 99.5127
R4195 VDD.n3554 VDD.n953 99.5127
R4196 VDD.n3554 VDD.n947 99.5127
R4197 VDD.n3551 VDD.n947 99.5127
R4198 VDD.n3551 VDD.n941 99.5127
R4199 VDD.n3548 VDD.n941 99.5127
R4200 VDD.n3548 VDD.n935 99.5127
R4201 VDD.n3545 VDD.n935 99.5127
R4202 VDD.n3545 VDD.n929 99.5127
R4203 VDD.n3542 VDD.n929 99.5127
R4204 VDD.n3542 VDD.n923 99.5127
R4205 VDD.n3539 VDD.n923 99.5127
R4206 VDD.n3539 VDD.n917 99.5127
R4207 VDD.n3536 VDD.n917 99.5127
R4208 VDD.n3536 VDD.n911 99.5127
R4209 VDD.n3533 VDD.n911 99.5127
R4210 VDD.n3533 VDD.n905 99.5127
R4211 VDD.n3530 VDD.n905 99.5127
R4212 VDD.n3530 VDD.n899 99.5127
R4213 VDD.n3527 VDD.n899 99.5127
R4214 VDD.n3527 VDD.n893 99.5127
R4215 VDD.n3524 VDD.n893 99.5127
R4216 VDD.n3524 VDD.n887 99.5127
R4217 VDD.n3521 VDD.n887 99.5127
R4218 VDD.n3521 VDD.n881 99.5127
R4219 VDD.n3518 VDD.n881 99.5127
R4220 VDD.n3518 VDD.n875 99.5127
R4221 VDD.n3515 VDD.n875 99.5127
R4222 VDD.n3515 VDD.n869 99.5127
R4223 VDD.n3512 VDD.n869 99.5127
R4224 VDD.n3512 VDD.n863 99.5127
R4225 VDD.n3509 VDD.n863 99.5127
R4226 VDD.n3509 VDD.n857 99.5127
R4227 VDD.n3506 VDD.n857 99.5127
R4228 VDD.n3506 VDD.n851 99.5127
R4229 VDD.n3503 VDD.n851 99.5127
R4230 VDD.n3503 VDD.n845 99.5127
R4231 VDD.n3500 VDD.n845 99.5127
R4232 VDD.n3500 VDD.n839 99.5127
R4233 VDD.n3497 VDD.n839 99.5127
R4234 VDD.n3497 VDD.n833 99.5127
R4235 VDD.n3494 VDD.n833 99.5127
R4236 VDD.n3494 VDD.n826 99.5127
R4237 VDD.n3491 VDD.n826 99.5127
R4238 VDD.n3491 VDD.n820 99.5127
R4239 VDD.n3488 VDD.n820 99.5127
R4240 VDD.n3488 VDD.n815 99.5127
R4241 VDD.n3485 VDD.n815 99.5127
R4242 VDD.n3485 VDD.n809 99.5127
R4243 VDD.n3482 VDD.n809 99.5127
R4244 VDD.n3482 VDD.n803 99.5127
R4245 VDD.n3479 VDD.n803 99.5127
R4246 VDD.n3479 VDD.n797 99.5127
R4247 VDD.n3476 VDD.n797 99.5127
R4248 VDD.n3476 VDD.n791 99.5127
R4249 VDD.n3473 VDD.n791 99.5127
R4250 VDD.n3473 VDD.n785 99.5127
R4251 VDD.n3470 VDD.n785 99.5127
R4252 VDD.n3470 VDD.n779 99.5127
R4253 VDD.n3467 VDD.n779 99.5127
R4254 VDD.n3467 VDD.n773 99.5127
R4255 VDD.n3464 VDD.n773 99.5127
R4256 VDD.n3464 VDD.n767 99.5127
R4257 VDD.n3461 VDD.n767 99.5127
R4258 VDD.n3461 VDD.n761 99.5127
R4259 VDD.n3458 VDD.n761 99.5127
R4260 VDD.n3458 VDD.n755 99.5127
R4261 VDD.n3455 VDD.n755 99.5127
R4262 VDD.n3455 VDD.n748 99.5127
R4263 VDD.n3452 VDD.n748 99.5127
R4264 VDD.n3452 VDD.n742 99.5127
R4265 VDD.n3449 VDD.n742 99.5127
R4266 VDD.n3449 VDD.n737 99.5127
R4267 VDD.n3446 VDD.n737 99.5127
R4268 VDD.n3446 VDD.n731 99.5127
R4269 VDD.n3443 VDD.n731 99.5127
R4270 VDD.n3443 VDD.n724 99.5127
R4271 VDD.n724 VDD.n716 99.5127
R4272 VDD.n4166 VDD.n716 99.5127
R4273 VDD.n4167 VDD.n4166 99.5127
R4274 VDD.n4167 VDD.n692 99.5127
R4275 VDD.n4172 VDD.n692 99.5127
R4276 VDD.n3403 VDD.n3402 99.5127
R4277 VDD.n3405 VDD.n3403 99.5127
R4278 VDD.n3409 VDD.n3398 99.5127
R4279 VDD.n3413 VDD.n3411 99.5127
R4280 VDD.n3417 VDD.n3396 99.5127
R4281 VDD.n3421 VDD.n3419 99.5127
R4282 VDD.n3425 VDD.n3394 99.5127
R4283 VDD.n3429 VDD.n3427 99.5127
R4284 VDD.n3434 VDD.n3390 99.5127
R4285 VDD.n3438 VDD.n3436 99.5127
R4286 VDD.n3384 VDD.n1059 99.5127
R4287 VDD.n3380 VDD.n3379 99.5127
R4288 VDD.n3376 VDD.n3375 99.5127
R4289 VDD.n3372 VDD.n3371 99.5127
R4290 VDD.n3368 VDD.n3367 99.5127
R4291 VDD.n3364 VDD.n3363 99.5127
R4292 VDD.n3360 VDD.n3359 99.5127
R4293 VDD.n3356 VDD.n3355 99.5127
R4294 VDD.n3352 VDD.n3351 99.5127
R4295 VDD.n3348 VDD.n3347 99.5127
R4296 VDD.n1572 VDD.n1398 99.5127
R4297 VDD.n1572 VDD.n1392 99.5127
R4298 VDD.n1569 VDD.n1392 99.5127
R4299 VDD.n1569 VDD.n1386 99.5127
R4300 VDD.n1566 VDD.n1386 99.5127
R4301 VDD.n1566 VDD.n1380 99.5127
R4302 VDD.n1563 VDD.n1380 99.5127
R4303 VDD.n1563 VDD.n1374 99.5127
R4304 VDD.n1560 VDD.n1374 99.5127
R4305 VDD.n1560 VDD.n1367 99.5127
R4306 VDD.n1557 VDD.n1367 99.5127
R4307 VDD.n1557 VDD.n1361 99.5127
R4308 VDD.n1554 VDD.n1361 99.5127
R4309 VDD.n1554 VDD.n1356 99.5127
R4310 VDD.n1551 VDD.n1356 99.5127
R4311 VDD.n1551 VDD.n1350 99.5127
R4312 VDD.n1548 VDD.n1350 99.5127
R4313 VDD.n1548 VDD.n1344 99.5127
R4314 VDD.n1545 VDD.n1344 99.5127
R4315 VDD.n1545 VDD.n1338 99.5127
R4316 VDD.n1542 VDD.n1338 99.5127
R4317 VDD.n1542 VDD.n1332 99.5127
R4318 VDD.n1539 VDD.n1332 99.5127
R4319 VDD.n1539 VDD.n1326 99.5127
R4320 VDD.n1536 VDD.n1326 99.5127
R4321 VDD.n1536 VDD.n1320 99.5127
R4322 VDD.n1533 VDD.n1320 99.5127
R4323 VDD.n1533 VDD.n1314 99.5127
R4324 VDD.n1530 VDD.n1314 99.5127
R4325 VDD.n1530 VDD.n1308 99.5127
R4326 VDD.n1527 VDD.n1308 99.5127
R4327 VDD.n1527 VDD.n1302 99.5127
R4328 VDD.n1524 VDD.n1302 99.5127
R4329 VDD.n1524 VDD.n1296 99.5127
R4330 VDD.n1521 VDD.n1296 99.5127
R4331 VDD.n1521 VDD.n1289 99.5127
R4332 VDD.n1518 VDD.n1289 99.5127
R4333 VDD.n1518 VDD.n1283 99.5127
R4334 VDD.n1515 VDD.n1283 99.5127
R4335 VDD.n1515 VDD.n1278 99.5127
R4336 VDD.n1512 VDD.n1278 99.5127
R4337 VDD.n1512 VDD.n1272 99.5127
R4338 VDD.n1509 VDD.n1272 99.5127
R4339 VDD.n1509 VDD.n1266 99.5127
R4340 VDD.n1506 VDD.n1266 99.5127
R4341 VDD.n1506 VDD.n1260 99.5127
R4342 VDD.n1503 VDD.n1260 99.5127
R4343 VDD.n1503 VDD.n1254 99.5127
R4344 VDD.n1500 VDD.n1254 99.5127
R4345 VDD.n1500 VDD.n1248 99.5127
R4346 VDD.n1497 VDD.n1248 99.5127
R4347 VDD.n1497 VDD.n1242 99.5127
R4348 VDD.n1494 VDD.n1242 99.5127
R4349 VDD.n1494 VDD.n1236 99.5127
R4350 VDD.n1491 VDD.n1236 99.5127
R4351 VDD.n1491 VDD.n1230 99.5127
R4352 VDD.n1488 VDD.n1230 99.5127
R4353 VDD.n1488 VDD.n1224 99.5127
R4354 VDD.n1485 VDD.n1224 99.5127
R4355 VDD.n1485 VDD.n1218 99.5127
R4356 VDD.n1482 VDD.n1218 99.5127
R4357 VDD.n1482 VDD.n1212 99.5127
R4358 VDD.n1479 VDD.n1212 99.5127
R4359 VDD.n1479 VDD.n1206 99.5127
R4360 VDD.n1476 VDD.n1206 99.5127
R4361 VDD.n1476 VDD.n1200 99.5127
R4362 VDD.n1473 VDD.n1200 99.5127
R4363 VDD.n1473 VDD.n1194 99.5127
R4364 VDD.n1470 VDD.n1194 99.5127
R4365 VDD.n1470 VDD.n1188 99.5127
R4366 VDD.n1467 VDD.n1188 99.5127
R4367 VDD.n1467 VDD.n1182 99.5127
R4368 VDD.n1464 VDD.n1182 99.5127
R4369 VDD.n1464 VDD.n1176 99.5127
R4370 VDD.n1461 VDD.n1176 99.5127
R4371 VDD.n1461 VDD.n1170 99.5127
R4372 VDD.n1458 VDD.n1170 99.5127
R4373 VDD.n1458 VDD.n1164 99.5127
R4374 VDD.n1455 VDD.n1164 99.5127
R4375 VDD.n1455 VDD.n1158 99.5127
R4376 VDD.n1452 VDD.n1158 99.5127
R4377 VDD.n1452 VDD.n1152 99.5127
R4378 VDD.n1449 VDD.n1152 99.5127
R4379 VDD.n1449 VDD.n1146 99.5127
R4380 VDD.n1446 VDD.n1146 99.5127
R4381 VDD.n1446 VDD.n1140 99.5127
R4382 VDD.n1443 VDD.n1140 99.5127
R4383 VDD.n1443 VDD.n1134 99.5127
R4384 VDD.n1440 VDD.n1134 99.5127
R4385 VDD.n1440 VDD.n1128 99.5127
R4386 VDD.n1437 VDD.n1128 99.5127
R4387 VDD.n1437 VDD.n1122 99.5127
R4388 VDD.n1434 VDD.n1122 99.5127
R4389 VDD.n1434 VDD.n1115 99.5127
R4390 VDD.n1431 VDD.n1115 99.5127
R4391 VDD.n1431 VDD.n1108 99.5127
R4392 VDD.n1428 VDD.n1108 99.5127
R4393 VDD.n1428 VDD.n1103 99.5127
R4394 VDD.n1425 VDD.n1103 99.5127
R4395 VDD.n1425 VDD.n1098 99.5127
R4396 VDD.n1422 VDD.n1098 99.5127
R4397 VDD.n1422 VDD.n1091 99.5127
R4398 VDD.n1419 VDD.n1091 99.5127
R4399 VDD.n1419 VDD.n1085 99.5127
R4400 VDD.n1416 VDD.n1085 99.5127
R4401 VDD.n1416 VDD.n1074 99.5127
R4402 VDD.n1074 VDD.n1065 99.5127
R4403 VDD.n3342 VDD.n1065 99.5127
R4404 VDD.n3343 VDD.n3342 99.5127
R4405 VDD.n2959 VDD.n2957 99.5127
R4406 VDD.n2957 VDD.n2956 99.5127
R4407 VDD.n2953 VDD.n2952 99.5127
R4408 VDD.n2950 VDD.n1404 99.5127
R4409 VDD.n2946 VDD.n2944 99.5127
R4410 VDD.n2942 VDD.n1406 99.5127
R4411 VDD.n1592 VDD.n1590 99.5127
R4412 VDD.n1588 VDD.n1408 99.5127
R4413 VDD.n1584 VDD.n1582 99.5127
R4414 VDD.n1579 VDD.n1578 99.5127
R4415 VDD.n2963 VDD.n1390 99.5127
R4416 VDD.n2971 VDD.n1390 99.5127
R4417 VDD.n2971 VDD.n1388 99.5127
R4418 VDD.n2975 VDD.n1388 99.5127
R4419 VDD.n2975 VDD.n1378 99.5127
R4420 VDD.n2983 VDD.n1378 99.5127
R4421 VDD.n2983 VDD.n1376 99.5127
R4422 VDD.n2987 VDD.n1376 99.5127
R4423 VDD.n2987 VDD.n1365 99.5127
R4424 VDD.n2995 VDD.n1365 99.5127
R4425 VDD.n2995 VDD.n1363 99.5127
R4426 VDD.n2999 VDD.n1363 99.5127
R4427 VDD.n2999 VDD.n1354 99.5127
R4428 VDD.n3007 VDD.n1354 99.5127
R4429 VDD.n3007 VDD.n1352 99.5127
R4430 VDD.n3011 VDD.n1352 99.5127
R4431 VDD.n3011 VDD.n1342 99.5127
R4432 VDD.n3019 VDD.n1342 99.5127
R4433 VDD.n3019 VDD.n1340 99.5127
R4434 VDD.n3023 VDD.n1340 99.5127
R4435 VDD.n3023 VDD.n1330 99.5127
R4436 VDD.n3031 VDD.n1330 99.5127
R4437 VDD.n3031 VDD.n1328 99.5127
R4438 VDD.n3035 VDD.n1328 99.5127
R4439 VDD.n3035 VDD.n1318 99.5127
R4440 VDD.n3043 VDD.n1318 99.5127
R4441 VDD.n3043 VDD.n1316 99.5127
R4442 VDD.n3047 VDD.n1316 99.5127
R4443 VDD.n3047 VDD.n1306 99.5127
R4444 VDD.n3055 VDD.n1306 99.5127
R4445 VDD.n3055 VDD.n1304 99.5127
R4446 VDD.n3059 VDD.n1304 99.5127
R4447 VDD.n3059 VDD.n1294 99.5127
R4448 VDD.n3067 VDD.n1294 99.5127
R4449 VDD.n3067 VDD.n1292 99.5127
R4450 VDD.n3071 VDD.n1292 99.5127
R4451 VDD.n3071 VDD.n1282 99.5127
R4452 VDD.n3079 VDD.n1282 99.5127
R4453 VDD.n3079 VDD.n1280 99.5127
R4454 VDD.n3083 VDD.n1280 99.5127
R4455 VDD.n3083 VDD.n1270 99.5127
R4456 VDD.n3091 VDD.n1270 99.5127
R4457 VDD.n3091 VDD.n1268 99.5127
R4458 VDD.n3095 VDD.n1268 99.5127
R4459 VDD.n3095 VDD.n1258 99.5127
R4460 VDD.n3103 VDD.n1258 99.5127
R4461 VDD.n3103 VDD.n1256 99.5127
R4462 VDD.n3107 VDD.n1256 99.5127
R4463 VDD.n3107 VDD.n1246 99.5127
R4464 VDD.n3115 VDD.n1246 99.5127
R4465 VDD.n3115 VDD.n1244 99.5127
R4466 VDD.n3119 VDD.n1244 99.5127
R4467 VDD.n3119 VDD.n1234 99.5127
R4468 VDD.n3127 VDD.n1234 99.5127
R4469 VDD.n3127 VDD.n1232 99.5127
R4470 VDD.n3131 VDD.n1232 99.5127
R4471 VDD.n3131 VDD.n1222 99.5127
R4472 VDD.n3139 VDD.n1222 99.5127
R4473 VDD.n3139 VDD.n1220 99.5127
R4474 VDD.n3143 VDD.n1220 99.5127
R4475 VDD.n3143 VDD.n1210 99.5127
R4476 VDD.n3151 VDD.n1210 99.5127
R4477 VDD.n3151 VDD.n1208 99.5127
R4478 VDD.n3155 VDD.n1208 99.5127
R4479 VDD.n3155 VDD.n1198 99.5127
R4480 VDD.n3163 VDD.n1198 99.5127
R4481 VDD.n3163 VDD.n1196 99.5127
R4482 VDD.n3167 VDD.n1196 99.5127
R4483 VDD.n3167 VDD.n1186 99.5127
R4484 VDD.n3175 VDD.n1186 99.5127
R4485 VDD.n3175 VDD.n1184 99.5127
R4486 VDD.n3179 VDD.n1184 99.5127
R4487 VDD.n3179 VDD.n1174 99.5127
R4488 VDD.n3187 VDD.n1174 99.5127
R4489 VDD.n3187 VDD.n1172 99.5127
R4490 VDD.n3191 VDD.n1172 99.5127
R4491 VDD.n3191 VDD.n1162 99.5127
R4492 VDD.n3199 VDD.n1162 99.5127
R4493 VDD.n3199 VDD.n1160 99.5127
R4494 VDD.n3203 VDD.n1160 99.5127
R4495 VDD.n3203 VDD.n1150 99.5127
R4496 VDD.n3211 VDD.n1150 99.5127
R4497 VDD.n3211 VDD.n1148 99.5127
R4498 VDD.n3215 VDD.n1148 99.5127
R4499 VDD.n3215 VDD.n1138 99.5127
R4500 VDD.n3223 VDD.n1138 99.5127
R4501 VDD.n3223 VDD.n1136 99.5127
R4502 VDD.n3227 VDD.n1136 99.5127
R4503 VDD.n3227 VDD.n1126 99.5127
R4504 VDD.n3235 VDD.n1126 99.5127
R4505 VDD.n3235 VDD.n1124 99.5127
R4506 VDD.n3239 VDD.n1124 99.5127
R4507 VDD.n3239 VDD.n1113 99.5127
R4508 VDD.n3247 VDD.n1113 99.5127
R4509 VDD.n3247 VDD.n1111 99.5127
R4510 VDD.n3251 VDD.n1111 99.5127
R4511 VDD.n3251 VDD.n1102 99.5127
R4512 VDD.n3259 VDD.n1102 99.5127
R4513 VDD.n3259 VDD.n1100 99.5127
R4514 VDD.n3263 VDD.n1100 99.5127
R4515 VDD.n3263 VDD.n1089 99.5127
R4516 VDD.n3273 VDD.n1089 99.5127
R4517 VDD.n3273 VDD.n1087 99.5127
R4518 VDD.n3277 VDD.n1087 99.5127
R4519 VDD.n3277 VDD.n1072 99.5127
R4520 VDD.n3336 VDD.n1072 99.5127
R4521 VDD.n3336 VDD.n1070 99.5127
R4522 VDD.n3340 VDD.n1070 99.5127
R4523 VDD.n3340 VDD.n1058 99.5127
R4524 VDD.n4149 VDD.n4148 99.5127
R4525 VDD.n4146 VDD.n4129 99.5127
R4526 VDD.n4142 VDD.n4141 99.5127
R4527 VDD.n4139 VDD.n4132 99.5127
R4528 VDD.n4135 VDD.n4134 99.5127
R4529 VDD.n4236 VDD.n4235 99.5127
R4530 VDD.n4233 VDD.n680 99.5127
R4531 VDD.n4229 VDD.n4228 99.5127
R4532 VDD.n4226 VDD.n683 99.5127
R4533 VDD.n4221 VDD.n4220 99.5127
R4534 VDD.n3770 VDD.n3599 99.5127
R4535 VDD.n3770 VDD.n1032 99.5127
R4536 VDD.n3767 VDD.n1032 99.5127
R4537 VDD.n3767 VDD.n1026 99.5127
R4538 VDD.n3764 VDD.n1026 99.5127
R4539 VDD.n3764 VDD.n1020 99.5127
R4540 VDD.n3761 VDD.n1020 99.5127
R4541 VDD.n3761 VDD.n1014 99.5127
R4542 VDD.n3758 VDD.n1014 99.5127
R4543 VDD.n3758 VDD.n1007 99.5127
R4544 VDD.n3755 VDD.n1007 99.5127
R4545 VDD.n3755 VDD.n1000 99.5127
R4546 VDD.n3752 VDD.n1000 99.5127
R4547 VDD.n3752 VDD.n995 99.5127
R4548 VDD.n3749 VDD.n995 99.5127
R4549 VDD.n3749 VDD.n990 99.5127
R4550 VDD.n3746 VDD.n990 99.5127
R4551 VDD.n3746 VDD.n984 99.5127
R4552 VDD.n3743 VDD.n984 99.5127
R4553 VDD.n3743 VDD.n978 99.5127
R4554 VDD.n3740 VDD.n978 99.5127
R4555 VDD.n3740 VDD.n972 99.5127
R4556 VDD.n3737 VDD.n972 99.5127
R4557 VDD.n3737 VDD.n966 99.5127
R4558 VDD.n3734 VDD.n966 99.5127
R4559 VDD.n3734 VDD.n960 99.5127
R4560 VDD.n3731 VDD.n960 99.5127
R4561 VDD.n3731 VDD.n954 99.5127
R4562 VDD.n3728 VDD.n954 99.5127
R4563 VDD.n3728 VDD.n948 99.5127
R4564 VDD.n3725 VDD.n948 99.5127
R4565 VDD.n3725 VDD.n942 99.5127
R4566 VDD.n3722 VDD.n942 99.5127
R4567 VDD.n3722 VDD.n936 99.5127
R4568 VDD.n3719 VDD.n936 99.5127
R4569 VDD.n3719 VDD.n930 99.5127
R4570 VDD.n3716 VDD.n930 99.5127
R4571 VDD.n3716 VDD.n924 99.5127
R4572 VDD.n3713 VDD.n924 99.5127
R4573 VDD.n3713 VDD.n918 99.5127
R4574 VDD.n3710 VDD.n918 99.5127
R4575 VDD.n3710 VDD.n912 99.5127
R4576 VDD.n3707 VDD.n912 99.5127
R4577 VDD.n3707 VDD.n906 99.5127
R4578 VDD.n3704 VDD.n906 99.5127
R4579 VDD.n3704 VDD.n900 99.5127
R4580 VDD.n3701 VDD.n900 99.5127
R4581 VDD.n3701 VDD.n894 99.5127
R4582 VDD.n3698 VDD.n894 99.5127
R4583 VDD.n3698 VDD.n888 99.5127
R4584 VDD.n3695 VDD.n888 99.5127
R4585 VDD.n3695 VDD.n882 99.5127
R4586 VDD.n3692 VDD.n882 99.5127
R4587 VDD.n3692 VDD.n876 99.5127
R4588 VDD.n3689 VDD.n876 99.5127
R4589 VDD.n3689 VDD.n870 99.5127
R4590 VDD.n3686 VDD.n870 99.5127
R4591 VDD.n3686 VDD.n864 99.5127
R4592 VDD.n3683 VDD.n864 99.5127
R4593 VDD.n3683 VDD.n858 99.5127
R4594 VDD.n3680 VDD.n858 99.5127
R4595 VDD.n3680 VDD.n852 99.5127
R4596 VDD.n3677 VDD.n852 99.5127
R4597 VDD.n3677 VDD.n846 99.5127
R4598 VDD.n3674 VDD.n846 99.5127
R4599 VDD.n3674 VDD.n840 99.5127
R4600 VDD.n3671 VDD.n840 99.5127
R4601 VDD.n3671 VDD.n834 99.5127
R4602 VDD.n3668 VDD.n834 99.5127
R4603 VDD.n3668 VDD.n827 99.5127
R4604 VDD.n3665 VDD.n827 99.5127
R4605 VDD.n3665 VDD.n821 99.5127
R4606 VDD.n3662 VDD.n821 99.5127
R4607 VDD.n3662 VDD.n816 99.5127
R4608 VDD.n3659 VDD.n816 99.5127
R4609 VDD.n3659 VDD.n810 99.5127
R4610 VDD.n3656 VDD.n810 99.5127
R4611 VDD.n3656 VDD.n804 99.5127
R4612 VDD.n3653 VDD.n804 99.5127
R4613 VDD.n3653 VDD.n798 99.5127
R4614 VDD.n3650 VDD.n798 99.5127
R4615 VDD.n3650 VDD.n792 99.5127
R4616 VDD.n3647 VDD.n792 99.5127
R4617 VDD.n3647 VDD.n786 99.5127
R4618 VDD.n3644 VDD.n786 99.5127
R4619 VDD.n3644 VDD.n780 99.5127
R4620 VDD.n3641 VDD.n780 99.5127
R4621 VDD.n3641 VDD.n774 99.5127
R4622 VDD.n3638 VDD.n774 99.5127
R4623 VDD.n3638 VDD.n768 99.5127
R4624 VDD.n3635 VDD.n768 99.5127
R4625 VDD.n3635 VDD.n762 99.5127
R4626 VDD.n3632 VDD.n762 99.5127
R4627 VDD.n3632 VDD.n756 99.5127
R4628 VDD.n3629 VDD.n756 99.5127
R4629 VDD.n3629 VDD.n749 99.5127
R4630 VDD.n3626 VDD.n749 99.5127
R4631 VDD.n3626 VDD.n743 99.5127
R4632 VDD.n3623 VDD.n743 99.5127
R4633 VDD.n3623 VDD.n738 99.5127
R4634 VDD.n3620 VDD.n738 99.5127
R4635 VDD.n3620 VDD.n732 99.5127
R4636 VDD.n3617 VDD.n732 99.5127
R4637 VDD.n3617 VDD.n725 99.5127
R4638 VDD.n3614 VDD.n725 99.5127
R4639 VDD.n3614 VDD.n718 99.5127
R4640 VDD.n718 VDD.n690 99.5127
R4641 VDD.n4214 VDD.n690 99.5127
R4642 VDD.n4214 VDD.n688 99.5127
R4643 VDD.n3812 VDD.n3810 99.5127
R4644 VDD.n3808 VDD.n3602 99.5127
R4645 VDD.n3804 VDD.n3802 99.5127
R4646 VDD.n3800 VDD.n3604 99.5127
R4647 VDD.n3796 VDD.n3794 99.5127
R4648 VDD.n3792 VDD.n3606 99.5127
R4649 VDD.n3788 VDD.n3786 99.5127
R4650 VDD.n3784 VDD.n3608 99.5127
R4651 VDD.n3779 VDD.n3777 99.5127
R4652 VDD.n3775 VDD.n3612 99.5127
R4653 VDD.n3816 VDD.n1029 99.5127
R4654 VDD.n3824 VDD.n1029 99.5127
R4655 VDD.n3824 VDD.n1027 99.5127
R4656 VDD.n3828 VDD.n1027 99.5127
R4657 VDD.n3828 VDD.n1017 99.5127
R4658 VDD.n3836 VDD.n1017 99.5127
R4659 VDD.n3836 VDD.n1015 99.5127
R4660 VDD.n3840 VDD.n1015 99.5127
R4661 VDD.n3840 VDD.n1004 99.5127
R4662 VDD.n3848 VDD.n1004 99.5127
R4663 VDD.n3848 VDD.n1002 99.5127
R4664 VDD.n3852 VDD.n1002 99.5127
R4665 VDD.n3852 VDD.n993 99.5127
R4666 VDD.n3860 VDD.n993 99.5127
R4667 VDD.n3860 VDD.n991 99.5127
R4668 VDD.n3864 VDD.n991 99.5127
R4669 VDD.n3864 VDD.n981 99.5127
R4670 VDD.n3872 VDD.n981 99.5127
R4671 VDD.n3872 VDD.n979 99.5127
R4672 VDD.n3876 VDD.n979 99.5127
R4673 VDD.n3876 VDD.n969 99.5127
R4674 VDD.n3884 VDD.n969 99.5127
R4675 VDD.n3884 VDD.n967 99.5127
R4676 VDD.n3888 VDD.n967 99.5127
R4677 VDD.n3888 VDD.n957 99.5127
R4678 VDD.n3896 VDD.n957 99.5127
R4679 VDD.n3896 VDD.n955 99.5127
R4680 VDD.n3900 VDD.n955 99.5127
R4681 VDD.n3900 VDD.n945 99.5127
R4682 VDD.n3908 VDD.n945 99.5127
R4683 VDD.n3908 VDD.n943 99.5127
R4684 VDD.n3912 VDD.n943 99.5127
R4685 VDD.n3912 VDD.n933 99.5127
R4686 VDD.n3920 VDD.n933 99.5127
R4687 VDD.n3920 VDD.n931 99.5127
R4688 VDD.n3924 VDD.n931 99.5127
R4689 VDD.n3924 VDD.n921 99.5127
R4690 VDD.n3932 VDD.n921 99.5127
R4691 VDD.n3932 VDD.n919 99.5127
R4692 VDD.n3936 VDD.n919 99.5127
R4693 VDD.n3936 VDD.n909 99.5127
R4694 VDD.n3944 VDD.n909 99.5127
R4695 VDD.n3944 VDD.n907 99.5127
R4696 VDD.n3948 VDD.n907 99.5127
R4697 VDD.n3948 VDD.n897 99.5127
R4698 VDD.n3956 VDD.n897 99.5127
R4699 VDD.n3956 VDD.n895 99.5127
R4700 VDD.n3960 VDD.n895 99.5127
R4701 VDD.n3960 VDD.n885 99.5127
R4702 VDD.n3968 VDD.n885 99.5127
R4703 VDD.n3968 VDD.n883 99.5127
R4704 VDD.n3972 VDD.n883 99.5127
R4705 VDD.n3972 VDD.n873 99.5127
R4706 VDD.n3980 VDD.n873 99.5127
R4707 VDD.n3980 VDD.n871 99.5127
R4708 VDD.n3984 VDD.n871 99.5127
R4709 VDD.n3984 VDD.n861 99.5127
R4710 VDD.n3992 VDD.n861 99.5127
R4711 VDD.n3992 VDD.n859 99.5127
R4712 VDD.n3996 VDD.n859 99.5127
R4713 VDD.n3996 VDD.n849 99.5127
R4714 VDD.n4004 VDD.n849 99.5127
R4715 VDD.n4004 VDD.n847 99.5127
R4716 VDD.n4008 VDD.n847 99.5127
R4717 VDD.n4008 VDD.n837 99.5127
R4718 VDD.n4016 VDD.n837 99.5127
R4719 VDD.n4016 VDD.n835 99.5127
R4720 VDD.n4020 VDD.n835 99.5127
R4721 VDD.n4020 VDD.n824 99.5127
R4722 VDD.n4028 VDD.n824 99.5127
R4723 VDD.n4028 VDD.n822 99.5127
R4724 VDD.n4032 VDD.n822 99.5127
R4725 VDD.n4032 VDD.n813 99.5127
R4726 VDD.n4040 VDD.n813 99.5127
R4727 VDD.n4040 VDD.n811 99.5127
R4728 VDD.n4044 VDD.n811 99.5127
R4729 VDD.n4044 VDD.n801 99.5127
R4730 VDD.n4052 VDD.n801 99.5127
R4731 VDD.n4052 VDD.n799 99.5127
R4732 VDD.n4056 VDD.n799 99.5127
R4733 VDD.n4056 VDD.n789 99.5127
R4734 VDD.n4064 VDD.n789 99.5127
R4735 VDD.n4064 VDD.n787 99.5127
R4736 VDD.n4068 VDD.n787 99.5127
R4737 VDD.n4068 VDD.n777 99.5127
R4738 VDD.n4076 VDD.n777 99.5127
R4739 VDD.n4076 VDD.n775 99.5127
R4740 VDD.n4080 VDD.n775 99.5127
R4741 VDD.n4080 VDD.n765 99.5127
R4742 VDD.n4088 VDD.n765 99.5127
R4743 VDD.n4088 VDD.n763 99.5127
R4744 VDD.n4092 VDD.n763 99.5127
R4745 VDD.n4092 VDD.n753 99.5127
R4746 VDD.n4100 VDD.n753 99.5127
R4747 VDD.n4100 VDD.n751 99.5127
R4748 VDD.n4104 VDD.n751 99.5127
R4749 VDD.n4104 VDD.n741 99.5127
R4750 VDD.n4112 VDD.n741 99.5127
R4751 VDD.n4112 VDD.n739 99.5127
R4752 VDD.n4116 VDD.n739 99.5127
R4753 VDD.n4116 VDD.n729 99.5127
R4754 VDD.n4124 VDD.n729 99.5127
R4755 VDD.n4124 VDD.n726 99.5127
R4756 VDD.n4158 VDD.n726 99.5127
R4757 VDD.n4158 VDD.n727 99.5127
R4758 VDD.n727 VDD.n719 99.5127
R4759 VDD.n4153 VDD.n719 99.5127
R4760 VDD.n4153 VDD.n694 99.5127
R4761 VDD.n4150 VDD.n694 99.5127
R4762 VDD.n3326 VDD.n1037 99.5127
R4763 VDD.n3324 VDD.n3323 99.5127
R4764 VDD.n3320 VDD.n3319 99.5127
R4765 VDD.n3316 VDD.n3315 99.5127
R4766 VDD.n3312 VDD.n3311 99.5127
R4767 VDD.n3308 VDD.n3307 99.5127
R4768 VDD.n3304 VDD.n3303 99.5127
R4769 VDD.n3300 VDD.n3299 99.5127
R4770 VDD.n3296 VDD.n3295 99.5127
R4771 VDD.n3292 VDD.n3291 99.5127
R4772 VDD.n1779 VDD.n1399 99.5127
R4773 VDD.n1779 VDD.n1393 99.5127
R4774 VDD.n1776 VDD.n1393 99.5127
R4775 VDD.n1776 VDD.n1387 99.5127
R4776 VDD.n1773 VDD.n1387 99.5127
R4777 VDD.n1773 VDD.n1381 99.5127
R4778 VDD.n1770 VDD.n1381 99.5127
R4779 VDD.n1770 VDD.n1375 99.5127
R4780 VDD.n1767 VDD.n1375 99.5127
R4781 VDD.n1767 VDD.n1368 99.5127
R4782 VDD.n1764 VDD.n1368 99.5127
R4783 VDD.n1764 VDD.n1362 99.5127
R4784 VDD.n1761 VDD.n1362 99.5127
R4785 VDD.n1761 VDD.n1357 99.5127
R4786 VDD.n1758 VDD.n1357 99.5127
R4787 VDD.n1758 VDD.n1351 99.5127
R4788 VDD.n1755 VDD.n1351 99.5127
R4789 VDD.n1755 VDD.n1345 99.5127
R4790 VDD.n1752 VDD.n1345 99.5127
R4791 VDD.n1752 VDD.n1339 99.5127
R4792 VDD.n1749 VDD.n1339 99.5127
R4793 VDD.n1749 VDD.n1333 99.5127
R4794 VDD.n1746 VDD.n1333 99.5127
R4795 VDD.n1746 VDD.n1327 99.5127
R4796 VDD.n1743 VDD.n1327 99.5127
R4797 VDD.n1743 VDD.n1321 99.5127
R4798 VDD.n1740 VDD.n1321 99.5127
R4799 VDD.n1740 VDD.n1315 99.5127
R4800 VDD.n1737 VDD.n1315 99.5127
R4801 VDD.n1737 VDD.n1309 99.5127
R4802 VDD.n1734 VDD.n1309 99.5127
R4803 VDD.n1734 VDD.n1303 99.5127
R4804 VDD.n1731 VDD.n1303 99.5127
R4805 VDD.n1731 VDD.n1297 99.5127
R4806 VDD.n1728 VDD.n1297 99.5127
R4807 VDD.n1728 VDD.n1290 99.5127
R4808 VDD.n1725 VDD.n1290 99.5127
R4809 VDD.n1725 VDD.n1284 99.5127
R4810 VDD.n1722 VDD.n1284 99.5127
R4811 VDD.n1722 VDD.n1279 99.5127
R4812 VDD.n1719 VDD.n1279 99.5127
R4813 VDD.n1719 VDD.n1273 99.5127
R4814 VDD.n1716 VDD.n1273 99.5127
R4815 VDD.n1716 VDD.n1267 99.5127
R4816 VDD.n1713 VDD.n1267 99.5127
R4817 VDD.n1713 VDD.n1261 99.5127
R4818 VDD.n1710 VDD.n1261 99.5127
R4819 VDD.n1710 VDD.n1255 99.5127
R4820 VDD.n1707 VDD.n1255 99.5127
R4821 VDD.n1707 VDD.n1249 99.5127
R4822 VDD.n1704 VDD.n1249 99.5127
R4823 VDD.n1704 VDD.n1243 99.5127
R4824 VDD.n1701 VDD.n1243 99.5127
R4825 VDD.n1701 VDD.n1237 99.5127
R4826 VDD.n1698 VDD.n1237 99.5127
R4827 VDD.n1698 VDD.n1231 99.5127
R4828 VDD.n1695 VDD.n1231 99.5127
R4829 VDD.n1695 VDD.n1225 99.5127
R4830 VDD.n1692 VDD.n1225 99.5127
R4831 VDD.n1692 VDD.n1219 99.5127
R4832 VDD.n1689 VDD.n1219 99.5127
R4833 VDD.n1689 VDD.n1213 99.5127
R4834 VDD.n1686 VDD.n1213 99.5127
R4835 VDD.n1686 VDD.n1207 99.5127
R4836 VDD.n1683 VDD.n1207 99.5127
R4837 VDD.n1683 VDD.n1201 99.5127
R4838 VDD.n1680 VDD.n1201 99.5127
R4839 VDD.n1680 VDD.n1195 99.5127
R4840 VDD.n1677 VDD.n1195 99.5127
R4841 VDD.n1677 VDD.n1189 99.5127
R4842 VDD.n1674 VDD.n1189 99.5127
R4843 VDD.n1674 VDD.n1183 99.5127
R4844 VDD.n1671 VDD.n1183 99.5127
R4845 VDD.n1671 VDD.n1177 99.5127
R4846 VDD.n1668 VDD.n1177 99.5127
R4847 VDD.n1668 VDD.n1171 99.5127
R4848 VDD.n1665 VDD.n1171 99.5127
R4849 VDD.n1665 VDD.n1165 99.5127
R4850 VDD.n1662 VDD.n1165 99.5127
R4851 VDD.n1662 VDD.n1159 99.5127
R4852 VDD.n1659 VDD.n1159 99.5127
R4853 VDD.n1659 VDD.n1153 99.5127
R4854 VDD.n1656 VDD.n1153 99.5127
R4855 VDD.n1656 VDD.n1147 99.5127
R4856 VDD.n1653 VDD.n1147 99.5127
R4857 VDD.n1653 VDD.n1141 99.5127
R4858 VDD.n1650 VDD.n1141 99.5127
R4859 VDD.n1650 VDD.n1135 99.5127
R4860 VDD.n1647 VDD.n1135 99.5127
R4861 VDD.n1647 VDD.n1129 99.5127
R4862 VDD.n1644 VDD.n1129 99.5127
R4863 VDD.n1644 VDD.n1123 99.5127
R4864 VDD.n1641 VDD.n1123 99.5127
R4865 VDD.n1641 VDD.n1116 99.5127
R4866 VDD.n1638 VDD.n1116 99.5127
R4867 VDD.n1638 VDD.n1109 99.5127
R4868 VDD.n1635 VDD.n1109 99.5127
R4869 VDD.n1635 VDD.n1104 99.5127
R4870 VDD.n1632 VDD.n1104 99.5127
R4871 VDD.n1632 VDD.n1099 99.5127
R4872 VDD.n1629 VDD.n1099 99.5127
R4873 VDD.n1629 VDD.n1092 99.5127
R4874 VDD.n1092 VDD.n1083 99.5127
R4875 VDD.n3279 VDD.n1083 99.5127
R4876 VDD.n3280 VDD.n3279 99.5127
R4877 VDD.n3280 VDD.n1075 99.5127
R4878 VDD.n3283 VDD.n1075 99.5127
R4879 VDD.n3283 VDD.n1068 99.5127
R4880 VDD.n3287 VDD.n1068 99.5127
R4881 VDD.n1605 VDD.n1603 99.5127
R4882 VDD.n1609 VDD.n1600 99.5127
R4883 VDD.n1613 VDD.n1611 99.5127
R4884 VDD.n1617 VDD.n1598 99.5127
R4885 VDD.n1802 VDD.n1619 99.5127
R4886 VDD.n1800 VDD.n1799 99.5127
R4887 VDD.n1796 VDD.n1795 99.5127
R4888 VDD.n1793 VDD.n1622 99.5127
R4889 VDD.n1788 VDD.n1786 99.5127
R4890 VDD.n1784 VDD.n1626 99.5127
R4891 VDD.n2965 VDD.n1394 99.5127
R4892 VDD.n2969 VDD.n1394 99.5127
R4893 VDD.n2969 VDD.n1384 99.5127
R4894 VDD.n2977 VDD.n1384 99.5127
R4895 VDD.n2977 VDD.n1382 99.5127
R4896 VDD.n2981 VDD.n1382 99.5127
R4897 VDD.n2981 VDD.n1372 99.5127
R4898 VDD.n2989 VDD.n1372 99.5127
R4899 VDD.n2989 VDD.n1370 99.5127
R4900 VDD.n2993 VDD.n1370 99.5127
R4901 VDD.n2993 VDD.n1360 99.5127
R4902 VDD.n3001 VDD.n1360 99.5127
R4903 VDD.n3001 VDD.n1358 99.5127
R4904 VDD.n3005 VDD.n1358 99.5127
R4905 VDD.n3005 VDD.n1348 99.5127
R4906 VDD.n3013 VDD.n1348 99.5127
R4907 VDD.n3013 VDD.n1346 99.5127
R4908 VDD.n3017 VDD.n1346 99.5127
R4909 VDD.n3017 VDD.n1336 99.5127
R4910 VDD.n3025 VDD.n1336 99.5127
R4911 VDD.n3025 VDD.n1334 99.5127
R4912 VDD.n3029 VDD.n1334 99.5127
R4913 VDD.n3029 VDD.n1324 99.5127
R4914 VDD.n3037 VDD.n1324 99.5127
R4915 VDD.n3037 VDD.n1322 99.5127
R4916 VDD.n3041 VDD.n1322 99.5127
R4917 VDD.n3041 VDD.n1312 99.5127
R4918 VDD.n3049 VDD.n1312 99.5127
R4919 VDD.n3049 VDD.n1310 99.5127
R4920 VDD.n3053 VDD.n1310 99.5127
R4921 VDD.n3053 VDD.n1300 99.5127
R4922 VDD.n3061 VDD.n1300 99.5127
R4923 VDD.n3061 VDD.n1298 99.5127
R4924 VDD.n3065 VDD.n1298 99.5127
R4925 VDD.n3065 VDD.n1287 99.5127
R4926 VDD.n3073 VDD.n1287 99.5127
R4927 VDD.n3073 VDD.n1285 99.5127
R4928 VDD.n3077 VDD.n1285 99.5127
R4929 VDD.n3077 VDD.n1276 99.5127
R4930 VDD.n3085 VDD.n1276 99.5127
R4931 VDD.n3085 VDD.n1274 99.5127
R4932 VDD.n3089 VDD.n1274 99.5127
R4933 VDD.n3089 VDD.n1264 99.5127
R4934 VDD.n3097 VDD.n1264 99.5127
R4935 VDD.n3097 VDD.n1262 99.5127
R4936 VDD.n3101 VDD.n1262 99.5127
R4937 VDD.n3101 VDD.n1252 99.5127
R4938 VDD.n3109 VDD.n1252 99.5127
R4939 VDD.n3109 VDD.n1250 99.5127
R4940 VDD.n3113 VDD.n1250 99.5127
R4941 VDD.n3113 VDD.n1240 99.5127
R4942 VDD.n3121 VDD.n1240 99.5127
R4943 VDD.n3121 VDD.n1238 99.5127
R4944 VDD.n3125 VDD.n1238 99.5127
R4945 VDD.n3125 VDD.n1228 99.5127
R4946 VDD.n3133 VDD.n1228 99.5127
R4947 VDD.n3133 VDD.n1226 99.5127
R4948 VDD.n3137 VDD.n1226 99.5127
R4949 VDD.n3137 VDD.n1216 99.5127
R4950 VDD.n3145 VDD.n1216 99.5127
R4951 VDD.n3145 VDD.n1214 99.5127
R4952 VDD.n3149 VDD.n1214 99.5127
R4953 VDD.n3149 VDD.n1204 99.5127
R4954 VDD.n3157 VDD.n1204 99.5127
R4955 VDD.n3157 VDD.n1202 99.5127
R4956 VDD.n3161 VDD.n1202 99.5127
R4957 VDD.n3161 VDD.n1192 99.5127
R4958 VDD.n3169 VDD.n1192 99.5127
R4959 VDD.n3169 VDD.n1190 99.5127
R4960 VDD.n3173 VDD.n1190 99.5127
R4961 VDD.n3173 VDD.n1180 99.5127
R4962 VDD.n3181 VDD.n1180 99.5127
R4963 VDD.n3181 VDD.n1178 99.5127
R4964 VDD.n3185 VDD.n1178 99.5127
R4965 VDD.n3185 VDD.n1168 99.5127
R4966 VDD.n3193 VDD.n1168 99.5127
R4967 VDD.n3193 VDD.n1166 99.5127
R4968 VDD.n3197 VDD.n1166 99.5127
R4969 VDD.n3197 VDD.n1156 99.5127
R4970 VDD.n3205 VDD.n1156 99.5127
R4971 VDD.n3205 VDD.n1154 99.5127
R4972 VDD.n3209 VDD.n1154 99.5127
R4973 VDD.n3209 VDD.n1144 99.5127
R4974 VDD.n3217 VDD.n1144 99.5127
R4975 VDD.n3217 VDD.n1142 99.5127
R4976 VDD.n3221 VDD.n1142 99.5127
R4977 VDD.n3221 VDD.n1132 99.5127
R4978 VDD.n3229 VDD.n1132 99.5127
R4979 VDD.n3229 VDD.n1130 99.5127
R4980 VDD.n3233 VDD.n1130 99.5127
R4981 VDD.n3233 VDD.n1120 99.5127
R4982 VDD.n3241 VDD.n1120 99.5127
R4983 VDD.n3241 VDD.n1118 99.5127
R4984 VDD.n3245 VDD.n1118 99.5127
R4985 VDD.n3245 VDD.n1107 99.5127
R4986 VDD.n3253 VDD.n1107 99.5127
R4987 VDD.n3253 VDD.n1105 99.5127
R4988 VDD.n3257 VDD.n1105 99.5127
R4989 VDD.n3257 VDD.n1096 99.5127
R4990 VDD.n3265 VDD.n1096 99.5127
R4991 VDD.n3265 VDD.n1093 99.5127
R4992 VDD.n3271 VDD.n1093 99.5127
R4993 VDD.n3271 VDD.n1094 99.5127
R4994 VDD.n1094 VDD.n1086 99.5127
R4995 VDD.n1086 VDD.n1076 99.5127
R4996 VDD.n3334 VDD.n1076 99.5127
R4997 VDD.n3334 VDD.n1077 99.5127
R4998 VDD.n1077 VDD.n1069 99.5127
R4999 VDD.n3329 VDD.n1069 99.5127
R5000 VDD.n1602 VDD.n1397 72.8958
R5001 VDD.n1604 VDD.n1397 72.8958
R5002 VDD.n1610 VDD.n1397 72.8958
R5003 VDD.n1612 VDD.n1397 72.8958
R5004 VDD.n1618 VDD.n1397 72.8958
R5005 VDD.n1801 VDD.n1397 72.8958
R5006 VDD.n1620 VDD.n1397 72.8958
R5007 VDD.n1794 VDD.n1397 72.8958
R5008 VDD.n1787 VDD.n1397 72.8958
R5009 VDD.n1785 VDD.n1397 72.8958
R5010 VDD.n3385 VDD.n1047 72.8958
R5011 VDD.n3385 VDD.n1046 72.8958
R5012 VDD.n3385 VDD.n1045 72.8958
R5013 VDD.n3385 VDD.n1044 72.8958
R5014 VDD.n3385 VDD.n1043 72.8958
R5015 VDD.n3385 VDD.n1042 72.8958
R5016 VDD.n3385 VDD.n1041 72.8958
R5017 VDD.n3385 VDD.n1040 72.8958
R5018 VDD.n3385 VDD.n1039 72.8958
R5019 VDD.n3385 VDD.n1038 72.8958
R5020 VDD.n3811 VDD.n3386 72.8958
R5021 VDD.n3809 VDD.n3386 72.8958
R5022 VDD.n3803 VDD.n3386 72.8958
R5023 VDD.n3801 VDD.n3386 72.8958
R5024 VDD.n3795 VDD.n3386 72.8958
R5025 VDD.n3793 VDD.n3386 72.8958
R5026 VDD.n3787 VDD.n3386 72.8958
R5027 VDD.n3785 VDD.n3386 72.8958
R5028 VDD.n3778 VDD.n3386 72.8958
R5029 VDD.n3776 VDD.n3386 72.8958
R5030 VDD.n4219 VDD.n679 72.8958
R5031 VDD.n687 VDD.n679 72.8958
R5032 VDD.n4227 VDD.n679 72.8958
R5033 VDD.n682 VDD.n679 72.8958
R5034 VDD.n4234 VDD.n679 72.8958
R5035 VDD.n679 VDD.n678 72.8958
R5036 VDD.n4133 VDD.n679 72.8958
R5037 VDD.n4140 VDD.n679 72.8958
R5038 VDD.n4131 VDD.n679 72.8958
R5039 VDD.n4147 VDD.n679 72.8958
R5040 VDD.n2958 VDD.n1397 72.8958
R5041 VDD.n1402 VDD.n1397 72.8958
R5042 VDD.n2951 VDD.n1397 72.8958
R5043 VDD.n2945 VDD.n1397 72.8958
R5044 VDD.n2943 VDD.n1397 72.8958
R5045 VDD.n1591 VDD.n1397 72.8958
R5046 VDD.n1589 VDD.n1397 72.8958
R5047 VDD.n1583 VDD.n1397 72.8958
R5048 VDD.n1412 VDD.n1397 72.8958
R5049 VDD.n1577 VDD.n1397 72.8958
R5050 VDD.n3385 VDD.n1048 72.8958
R5051 VDD.n3385 VDD.n1049 72.8958
R5052 VDD.n3385 VDD.n1050 72.8958
R5053 VDD.n3385 VDD.n1051 72.8958
R5054 VDD.n3385 VDD.n1052 72.8958
R5055 VDD.n3385 VDD.n1053 72.8958
R5056 VDD.n3385 VDD.n1054 72.8958
R5057 VDD.n3385 VDD.n1055 72.8958
R5058 VDD.n3385 VDD.n1056 72.8958
R5059 VDD.n3385 VDD.n1057 72.8958
R5060 VDD.n3401 VDD.n3386 72.8958
R5061 VDD.n3404 VDD.n3386 72.8958
R5062 VDD.n3410 VDD.n3386 72.8958
R5063 VDD.n3412 VDD.n3386 72.8958
R5064 VDD.n3418 VDD.n3386 72.8958
R5065 VDD.n3420 VDD.n3386 72.8958
R5066 VDD.n3426 VDD.n3386 72.8958
R5067 VDD.n3428 VDD.n3386 72.8958
R5068 VDD.n3435 VDD.n3386 72.8958
R5069 VDD.n3437 VDD.n3386 72.8958
R5070 VDD.n4171 VDD.n679 72.8958
R5071 VDD.n4178 VDD.n679 72.8958
R5072 VDD.n712 VDD.n679 72.8958
R5073 VDD.n4185 VDD.n679 72.8958
R5074 VDD.n707 VDD.n679 72.8958
R5075 VDD.n4192 VDD.n679 72.8958
R5076 VDD.n704 VDD.n679 72.8958
R5077 VDD.n4199 VDD.n679 72.8958
R5078 VDD.n701 VDD.n679 72.8958
R5079 VDD.n4206 VDD.n679 72.8958
R5080 VDD.n4243 VDD.n4242 66.2847
R5081 VDD.n4242 VDD.n547 66.2847
R5082 VDD.n4242 VDD.n548 66.2847
R5083 VDD.n4242 VDD.n549 66.2847
R5084 VDD.n4242 VDD.n550 66.2847
R5085 VDD.n4242 VDD.n551 66.2847
R5086 VDD.n4242 VDD.n552 66.2847
R5087 VDD.n4242 VDD.n553 66.2847
R5088 VDD.n4242 VDD.n554 66.2847
R5089 VDD.n4242 VDD.n555 66.2847
R5090 VDD.n4242 VDD.n556 66.2847
R5091 VDD.n4242 VDD.n557 66.2847
R5092 VDD.n4242 VDD.n558 66.2847
R5093 VDD.n4242 VDD.n559 66.2847
R5094 VDD.n4242 VDD.n560 66.2847
R5095 VDD.n4242 VDD.n561 66.2847
R5096 VDD.n4242 VDD.n562 66.2847
R5097 VDD.n4242 VDD.n563 66.2847
R5098 VDD.n4593 VDD.n4592 66.2847
R5099 VDD.n4593 VDD.n216 66.2847
R5100 VDD.n4593 VDD.n215 66.2847
R5101 VDD.n4593 VDD.n214 66.2847
R5102 VDD.n4593 VDD.n213 66.2847
R5103 VDD.n4593 VDD.n212 66.2847
R5104 VDD.n4593 VDD.n211 66.2847
R5105 VDD.n4593 VDD.n210 66.2847
R5106 VDD.n4593 VDD.n209 66.2847
R5107 VDD.n4593 VDD.n208 66.2847
R5108 VDD.n4593 VDD.n207 66.2847
R5109 VDD.n4593 VDD.n206 66.2847
R5110 VDD.n4593 VDD.n205 66.2847
R5111 VDD.n4593 VDD.n204 66.2847
R5112 VDD.n4593 VDD.n203 66.2847
R5113 VDD.n4593 VDD.n202 66.2847
R5114 VDD.n4593 VDD.n201 66.2847
R5115 VDD.n4593 VDD.n200 66.2847
R5116 VDD.n4593 VDD.n199 66.2847
R5117 VDD.n2907 VDD.n2906 66.2847
R5118 VDD.n2906 VDD.n2905 66.2847
R5119 VDD.n2906 VDD.n2903 66.2847
R5120 VDD.n2906 VDD.n2902 66.2847
R5121 VDD.n2906 VDD.n2900 66.2847
R5122 VDD.n2906 VDD.n2899 66.2847
R5123 VDD.n2906 VDD.n2897 66.2847
R5124 VDD.n2906 VDD.n2896 66.2847
R5125 VDD.n2906 VDD.n2894 66.2847
R5126 VDD.n2906 VDD.n2893 66.2847
R5127 VDD.n2906 VDD.n1845 66.2847
R5128 VDD.n2906 VDD.n1844 66.2847
R5129 VDD.n2906 VDD.n1843 66.2847
R5130 VDD.n2906 VDD.n1842 66.2847
R5131 VDD.n2906 VDD.n1841 66.2847
R5132 VDD.n2906 VDD.n1840 66.2847
R5133 VDD.n2906 VDD.n1839 66.2847
R5134 VDD.n2906 VDD.n1838 66.2847
R5135 VDD.n2906 VDD.n1837 66.2847
R5136 VDD.n2365 VDD.n2364 66.2847
R5137 VDD.n2364 VDD.n2230 66.2847
R5138 VDD.n2364 VDD.n2231 66.2847
R5139 VDD.n2364 VDD.n2232 66.2847
R5140 VDD.n2364 VDD.n2233 66.2847
R5141 VDD.n2364 VDD.n2234 66.2847
R5142 VDD.n2364 VDD.n2235 66.2847
R5143 VDD.n2364 VDD.n2236 66.2847
R5144 VDD.n2364 VDD.n2237 66.2847
R5145 VDD.n2364 VDD.n2238 66.2847
R5146 VDD.n2364 VDD.n2239 66.2847
R5147 VDD.n2364 VDD.n2240 66.2847
R5148 VDD.n2364 VDD.n2241 66.2847
R5149 VDD.n2364 VDD.n2242 66.2847
R5150 VDD.n2364 VDD.n2243 66.2847
R5151 VDD.n2364 VDD.n2244 66.2847
R5152 VDD.n2364 VDD.n2245 66.2847
R5153 VDD.n2364 VDD.n2246 66.2847
R5154 VDD.n250 VDD.n199 52.4337
R5155 VDD.n254 VDD.n200 52.4337
R5156 VDD.n260 VDD.n201 52.4337
R5157 VDD.n264 VDD.n202 52.4337
R5158 VDD.n270 VDD.n203 52.4337
R5159 VDD.n275 VDD.n204 52.4337
R5160 VDD.n281 VDD.n205 52.4337
R5161 VDD.n285 VDD.n206 52.4337
R5162 VDD.n291 VDD.n207 52.4337
R5163 VDD.n295 VDD.n208 52.4337
R5164 VDD.n301 VDD.n209 52.4337
R5165 VDD.n305 VDD.n210 52.4337
R5166 VDD.n311 VDD.n211 52.4337
R5167 VDD.n315 VDD.n212 52.4337
R5168 VDD.n321 VDD.n213 52.4337
R5169 VDD.n325 VDD.n214 52.4337
R5170 VDD.n331 VDD.n215 52.4337
R5171 VDD.n334 VDD.n216 52.4337
R5172 VDD.n4592 VDD.n4591 52.4337
R5173 VDD.n4243 VDD.n543 52.4337
R5174 VDD.n591 VDD.n547 52.4337
R5175 VDD.n593 VDD.n548 52.4337
R5176 VDD.n601 VDD.n549 52.4337
R5177 VDD.n603 VDD.n550 52.4337
R5178 VDD.n611 VDD.n551 52.4337
R5179 VDD.n613 VDD.n552 52.4337
R5180 VDD.n621 VDD.n553 52.4337
R5181 VDD.n623 VDD.n554 52.4337
R5182 VDD.n631 VDD.n555 52.4337
R5183 VDD.n633 VDD.n556 52.4337
R5184 VDD.n641 VDD.n557 52.4337
R5185 VDD.n644 VDD.n558 52.4337
R5186 VDD.n652 VDD.n559 52.4337
R5187 VDD.n654 VDD.n560 52.4337
R5188 VDD.n662 VDD.n561 52.4337
R5189 VDD.n664 VDD.n562 52.4337
R5190 VDD.n672 VDD.n563 52.4337
R5191 VDD.n4244 VDD.n4243 52.4337
R5192 VDD.n594 VDD.n547 52.4337
R5193 VDD.n600 VDD.n548 52.4337
R5194 VDD.n604 VDD.n549 52.4337
R5195 VDD.n610 VDD.n550 52.4337
R5196 VDD.n614 VDD.n551 52.4337
R5197 VDD.n620 VDD.n552 52.4337
R5198 VDD.n624 VDD.n553 52.4337
R5199 VDD.n630 VDD.n554 52.4337
R5200 VDD.n634 VDD.n555 52.4337
R5201 VDD.n640 VDD.n556 52.4337
R5202 VDD.n645 VDD.n557 52.4337
R5203 VDD.n651 VDD.n558 52.4337
R5204 VDD.n655 VDD.n559 52.4337
R5205 VDD.n661 VDD.n560 52.4337
R5206 VDD.n665 VDD.n561 52.4337
R5207 VDD.n671 VDD.n562 52.4337
R5208 VDD.n564 VDD.n563 52.4337
R5209 VDD.n4592 VDD.n217 52.4337
R5210 VDD.n332 VDD.n216 52.4337
R5211 VDD.n326 VDD.n215 52.4337
R5212 VDD.n322 VDD.n214 52.4337
R5213 VDD.n316 VDD.n213 52.4337
R5214 VDD.n312 VDD.n212 52.4337
R5215 VDD.n306 VDD.n211 52.4337
R5216 VDD.n302 VDD.n210 52.4337
R5217 VDD.n296 VDD.n209 52.4337
R5218 VDD.n292 VDD.n208 52.4337
R5219 VDD.n286 VDD.n207 52.4337
R5220 VDD.n282 VDD.n206 52.4337
R5221 VDD.n276 VDD.n205 52.4337
R5222 VDD.n271 VDD.n204 52.4337
R5223 VDD.n265 VDD.n203 52.4337
R5224 VDD.n261 VDD.n202 52.4337
R5225 VDD.n255 VDD.n201 52.4337
R5226 VDD.n251 VDD.n200 52.4337
R5227 VDD.n245 VDD.n199 52.4337
R5228 VDD.n2843 VDD.n1837 52.4337
R5229 VDD.n2849 VDD.n1838 52.4337
R5230 VDD.n2851 VDD.n1839 52.4337
R5231 VDD.n2859 VDD.n1840 52.4337
R5232 VDD.n2861 VDD.n1841 52.4337
R5233 VDD.n2869 VDD.n1842 52.4337
R5234 VDD.n2874 VDD.n1843 52.4337
R5235 VDD.n2882 VDD.n1844 52.4337
R5236 VDD.n2884 VDD.n1845 52.4337
R5237 VDD.n2893 VDD.n2892 52.4337
R5238 VDD.n2894 VDD.n1809 52.4337
R5239 VDD.n2896 VDD.n2895 52.4337
R5240 VDD.n2897 VDD.n1816 52.4337
R5241 VDD.n2899 VDD.n2898 52.4337
R5242 VDD.n2900 VDD.n1821 52.4337
R5243 VDD.n2902 VDD.n2901 52.4337
R5244 VDD.n2903 VDD.n1826 52.4337
R5245 VDD.n2905 VDD.n2904 52.4337
R5246 VDD.n2907 VDD.n1831 52.4337
R5247 VDD.n2908 VDD.n2907 52.4337
R5248 VDD.n2905 VDD.n1830 52.4337
R5249 VDD.n2903 VDD.n1827 52.4337
R5250 VDD.n2902 VDD.n1825 52.4337
R5251 VDD.n2900 VDD.n1822 52.4337
R5252 VDD.n2899 VDD.n1820 52.4337
R5253 VDD.n2897 VDD.n1817 52.4337
R5254 VDD.n2896 VDD.n1813 52.4337
R5255 VDD.n2894 VDD.n1810 52.4337
R5256 VDD.n2893 VDD.n1808 52.4337
R5257 VDD.n2891 VDD.n1845 52.4337
R5258 VDD.n2885 VDD.n1844 52.4337
R5259 VDD.n2881 VDD.n1843 52.4337
R5260 VDD.n2875 VDD.n1842 52.4337
R5261 VDD.n2868 VDD.n1841 52.4337
R5262 VDD.n2862 VDD.n1840 52.4337
R5263 VDD.n2858 VDD.n1839 52.4337
R5264 VDD.n2852 VDD.n1838 52.4337
R5265 VDD.n2848 VDD.n1837 52.4337
R5266 VDD.n2366 VDD.n2365 52.4337
R5267 VDD.n2248 VDD.n2230 52.4337
R5268 VDD.n2252 VDD.n2231 52.4337
R5269 VDD.n2254 VDD.n2232 52.4337
R5270 VDD.n2258 VDD.n2233 52.4337
R5271 VDD.n2264 VDD.n2234 52.4337
R5272 VDD.n2266 VDD.n2235 52.4337
R5273 VDD.n2270 VDD.n2236 52.4337
R5274 VDD.n2272 VDD.n2237 52.4337
R5275 VDD.n2276 VDD.n2238 52.4337
R5276 VDD.n2278 VDD.n2239 52.4337
R5277 VDD.n2282 VDD.n2240 52.4337
R5278 VDD.n2284 VDD.n2241 52.4337
R5279 VDD.n2288 VDD.n2242 52.4337
R5280 VDD.n2290 VDD.n2243 52.4337
R5281 VDD.n2294 VDD.n2244 52.4337
R5282 VDD.n2296 VDD.n2245 52.4337
R5283 VDD.n2300 VDD.n2246 52.4337
R5284 VDD.n2365 VDD.n2229 52.4337
R5285 VDD.n2251 VDD.n2230 52.4337
R5286 VDD.n2253 VDD.n2231 52.4337
R5287 VDD.n2257 VDD.n2232 52.4337
R5288 VDD.n2259 VDD.n2233 52.4337
R5289 VDD.n2265 VDD.n2234 52.4337
R5290 VDD.n2269 VDD.n2235 52.4337
R5291 VDD.n2271 VDD.n2236 52.4337
R5292 VDD.n2275 VDD.n2237 52.4337
R5293 VDD.n2277 VDD.n2238 52.4337
R5294 VDD.n2281 VDD.n2239 52.4337
R5295 VDD.n2283 VDD.n2240 52.4337
R5296 VDD.n2287 VDD.n2241 52.4337
R5297 VDD.n2289 VDD.n2242 52.4337
R5298 VDD.n2293 VDD.n2243 52.4337
R5299 VDD.n2295 VDD.n2244 52.4337
R5300 VDD.n2299 VDD.n2245 52.4337
R5301 VDD.n2301 VDD.n2246 52.4337
R5302 VDD.n4206 VDD.n4205 39.2114
R5303 VDD.n4201 VDD.n701 39.2114
R5304 VDD.n4199 VDD.n4198 39.2114
R5305 VDD.n4194 VDD.n704 39.2114
R5306 VDD.n4192 VDD.n4191 39.2114
R5307 VDD.n4187 VDD.n707 39.2114
R5308 VDD.n4185 VDD.n4184 39.2114
R5309 VDD.n4180 VDD.n712 39.2114
R5310 VDD.n4178 VDD.n4177 39.2114
R5311 VDD.n4173 VDD.n4171 39.2114
R5312 VDD.n3401 VDD.n1035 39.2114
R5313 VDD.n3405 VDD.n3404 39.2114
R5314 VDD.n3410 VDD.n3409 39.2114
R5315 VDD.n3413 VDD.n3412 39.2114
R5316 VDD.n3418 VDD.n3417 39.2114
R5317 VDD.n3421 VDD.n3420 39.2114
R5318 VDD.n3426 VDD.n3425 39.2114
R5319 VDD.n3429 VDD.n3428 39.2114
R5320 VDD.n3435 VDD.n3434 39.2114
R5321 VDD.n3438 VDD.n3437 39.2114
R5322 VDD.n3380 VDD.n1057 39.2114
R5323 VDD.n3376 VDD.n1056 39.2114
R5324 VDD.n3372 VDD.n1055 39.2114
R5325 VDD.n3368 VDD.n1054 39.2114
R5326 VDD.n3364 VDD.n1053 39.2114
R5327 VDD.n3360 VDD.n1052 39.2114
R5328 VDD.n3356 VDD.n1051 39.2114
R5329 VDD.n3352 VDD.n1050 39.2114
R5330 VDD.n3348 VDD.n1049 39.2114
R5331 VDD.n3344 VDD.n1048 39.2114
R5332 VDD.n2958 VDD.n1400 39.2114
R5333 VDD.n2956 VDD.n1402 39.2114
R5334 VDD.n2952 VDD.n2951 39.2114
R5335 VDD.n2945 VDD.n1404 39.2114
R5336 VDD.n2944 VDD.n2943 39.2114
R5337 VDD.n1591 VDD.n1406 39.2114
R5338 VDD.n1590 VDD.n1589 39.2114
R5339 VDD.n1583 VDD.n1408 39.2114
R5340 VDD.n1582 VDD.n1412 39.2114
R5341 VDD.n1578 VDD.n1577 39.2114
R5342 VDD.n4147 VDD.n4146 39.2114
R5343 VDD.n4142 VDD.n4131 39.2114
R5344 VDD.n4140 VDD.n4139 39.2114
R5345 VDD.n4135 VDD.n4133 39.2114
R5346 VDD.n4236 VDD.n678 39.2114
R5347 VDD.n4234 VDD.n4233 39.2114
R5348 VDD.n4229 VDD.n682 39.2114
R5349 VDD.n4227 VDD.n4226 39.2114
R5350 VDD.n4221 VDD.n687 39.2114
R5351 VDD.n4219 VDD.n4218 39.2114
R5352 VDD.n3811 VDD.n3600 39.2114
R5353 VDD.n3810 VDD.n3809 39.2114
R5354 VDD.n3803 VDD.n3602 39.2114
R5355 VDD.n3802 VDD.n3801 39.2114
R5356 VDD.n3795 VDD.n3604 39.2114
R5357 VDD.n3794 VDD.n3793 39.2114
R5358 VDD.n3787 VDD.n3606 39.2114
R5359 VDD.n3786 VDD.n3785 39.2114
R5360 VDD.n3778 VDD.n3608 39.2114
R5361 VDD.n3777 VDD.n3776 39.2114
R5362 VDD.n3324 VDD.n1038 39.2114
R5363 VDD.n3320 VDD.n1039 39.2114
R5364 VDD.n3316 VDD.n1040 39.2114
R5365 VDD.n3312 VDD.n1041 39.2114
R5366 VDD.n3308 VDD.n1042 39.2114
R5367 VDD.n3304 VDD.n1043 39.2114
R5368 VDD.n3300 VDD.n1044 39.2114
R5369 VDD.n3296 VDD.n1045 39.2114
R5370 VDD.n3292 VDD.n1046 39.2114
R5371 VDD.n3288 VDD.n1047 39.2114
R5372 VDD.n1602 VDD.n1396 39.2114
R5373 VDD.n1605 VDD.n1604 39.2114
R5374 VDD.n1610 VDD.n1609 39.2114
R5375 VDD.n1613 VDD.n1612 39.2114
R5376 VDD.n1618 VDD.n1617 39.2114
R5377 VDD.n1802 VDD.n1801 39.2114
R5378 VDD.n1799 VDD.n1620 39.2114
R5379 VDD.n1795 VDD.n1794 39.2114
R5380 VDD.n1787 VDD.n1622 39.2114
R5381 VDD.n1786 VDD.n1785 39.2114
R5382 VDD.n1603 VDD.n1602 39.2114
R5383 VDD.n1604 VDD.n1600 39.2114
R5384 VDD.n1611 VDD.n1610 39.2114
R5385 VDD.n1612 VDD.n1598 39.2114
R5386 VDD.n1619 VDD.n1618 39.2114
R5387 VDD.n1801 VDD.n1800 39.2114
R5388 VDD.n1796 VDD.n1620 39.2114
R5389 VDD.n1794 VDD.n1793 39.2114
R5390 VDD.n1788 VDD.n1787 39.2114
R5391 VDD.n1785 VDD.n1784 39.2114
R5392 VDD.n3291 VDD.n1047 39.2114
R5393 VDD.n3295 VDD.n1046 39.2114
R5394 VDD.n3299 VDD.n1045 39.2114
R5395 VDD.n3303 VDD.n1044 39.2114
R5396 VDD.n3307 VDD.n1043 39.2114
R5397 VDD.n3311 VDD.n1042 39.2114
R5398 VDD.n3315 VDD.n1041 39.2114
R5399 VDD.n3319 VDD.n1040 39.2114
R5400 VDD.n3323 VDD.n1039 39.2114
R5401 VDD.n3326 VDD.n1038 39.2114
R5402 VDD.n3812 VDD.n3811 39.2114
R5403 VDD.n3809 VDD.n3808 39.2114
R5404 VDD.n3804 VDD.n3803 39.2114
R5405 VDD.n3801 VDD.n3800 39.2114
R5406 VDD.n3796 VDD.n3795 39.2114
R5407 VDD.n3793 VDD.n3792 39.2114
R5408 VDD.n3788 VDD.n3787 39.2114
R5409 VDD.n3785 VDD.n3784 39.2114
R5410 VDD.n3779 VDD.n3778 39.2114
R5411 VDD.n3776 VDD.n3775 39.2114
R5412 VDD.n4220 VDD.n4219 39.2114
R5413 VDD.n687 VDD.n683 39.2114
R5414 VDD.n4228 VDD.n4227 39.2114
R5415 VDD.n682 VDD.n680 39.2114
R5416 VDD.n4235 VDD.n4234 39.2114
R5417 VDD.n4134 VDD.n678 39.2114
R5418 VDD.n4133 VDD.n4132 39.2114
R5419 VDD.n4141 VDD.n4140 39.2114
R5420 VDD.n4131 VDD.n4129 39.2114
R5421 VDD.n4148 VDD.n4147 39.2114
R5422 VDD.n2959 VDD.n2958 39.2114
R5423 VDD.n2953 VDD.n1402 39.2114
R5424 VDD.n2951 VDD.n2950 39.2114
R5425 VDD.n2946 VDD.n2945 39.2114
R5426 VDD.n2943 VDD.n2942 39.2114
R5427 VDD.n1592 VDD.n1591 39.2114
R5428 VDD.n1589 VDD.n1588 39.2114
R5429 VDD.n1584 VDD.n1583 39.2114
R5430 VDD.n1579 VDD.n1412 39.2114
R5431 VDD.n1577 VDD.n1576 39.2114
R5432 VDD.n3347 VDD.n1048 39.2114
R5433 VDD.n3351 VDD.n1049 39.2114
R5434 VDD.n3355 VDD.n1050 39.2114
R5435 VDD.n3359 VDD.n1051 39.2114
R5436 VDD.n3363 VDD.n1052 39.2114
R5437 VDD.n3367 VDD.n1053 39.2114
R5438 VDD.n3371 VDD.n1054 39.2114
R5439 VDD.n3375 VDD.n1055 39.2114
R5440 VDD.n3379 VDD.n1056 39.2114
R5441 VDD.n1059 VDD.n1057 39.2114
R5442 VDD.n3402 VDD.n3401 39.2114
R5443 VDD.n3404 VDD.n3398 39.2114
R5444 VDD.n3411 VDD.n3410 39.2114
R5445 VDD.n3412 VDD.n3396 39.2114
R5446 VDD.n3419 VDD.n3418 39.2114
R5447 VDD.n3420 VDD.n3394 39.2114
R5448 VDD.n3427 VDD.n3426 39.2114
R5449 VDD.n3428 VDD.n3390 39.2114
R5450 VDD.n3436 VDD.n3435 39.2114
R5451 VDD.n3437 VDD.n3387 39.2114
R5452 VDD.n4171 VDD.n714 39.2114
R5453 VDD.n4179 VDD.n4178 39.2114
R5454 VDD.n712 VDD.n708 39.2114
R5455 VDD.n4186 VDD.n4185 39.2114
R5456 VDD.n707 VDD.n705 39.2114
R5457 VDD.n4193 VDD.n4192 39.2114
R5458 VDD.n704 VDD.n702 39.2114
R5459 VDD.n4200 VDD.n4199 39.2114
R5460 VDD.n701 VDD.n699 39.2114
R5461 VDD.n4207 VDD.n4206 39.2114
R5462 VDD.n3597 VDD.n3440 34.4981
R5463 VDD.n4174 VDD.n4170 34.4981
R5464 VDD.n3819 VDD.n1034 34.4981
R5465 VDD.n4210 VDD.n4209 34.4981
R5466 VDD.n4151 VDD.n4127 34.4981
R5467 VDD.n4217 VDD.n4216 34.4981
R5468 VDD.n3773 VDD.n3772 34.4981
R5469 VDD.n3815 VDD.n3814 34.4981
R5470 VDD.n2962 VDD.n2961 34.4981
R5471 VDD.n3383 VDD.n1060 34.4981
R5472 VDD.n3345 VDD.n1064 34.4981
R5473 VDD.n1575 VDD.n1574 34.4981
R5474 VDD.n3330 VDD.n3328 34.4981
R5475 VDD.n3289 VDD.n3286 34.4981
R5476 VDD.n1782 VDD.n1781 34.4981
R5477 VDD.n2966 VDD.n1395 34.4981
R5478 VDD.n2364 VDD.n2224 31.4725
R5479 VDD.n2906 VDD.n1836 31.4725
R5480 VDD.n4242 VDD.n538 31.4725
R5481 VDD.n4594 VDD.n4593 31.4725
R5482 VDD.n2306 VDD.n2305 30.8369
R5483 VDD.n2328 VDD.n2327 30.8369
R5484 VDD.n2262 VDD.n2261 30.8369
R5485 VDD.n567 VDD.n566 30.8369
R5486 VDD.n643 VDD.n576 30.8369
R5487 VDD.n585 VDD.n584 30.8369
R5488 VDD.n220 VDD.n219 30.8369
R5489 VDD.n230 VDD.n229 30.8369
R5490 VDD.n273 VDD.n238 30.8369
R5491 VDD.n2873 VDD.n2872 30.8369
R5492 VDD.n2930 VDD.n1815 30.8369
R5493 VDD.n2910 VDD.n1833 30.8369
R5494 VDD.n3781 VDD.n3610 24.049
R5495 VDD.n711 VDD.n710 24.049
R5496 VDD.n3432 VDD.n3392 24.049
R5497 VDD.n4224 VDD.n685 24.049
R5498 VDD.n1411 VDD.n1410 24.049
R5499 VDD.n1063 VDD.n1062 24.049
R5500 VDD.n1790 VDD.n1624 24.049
R5501 VDD.n1081 VDD.n1080 24.049
R5502 VDD.n32 VDD.t129 21.1764
R5503 VDD.n32 VDD.t157 21.1764
R5504 VDD.n30 VDD.t146 21.1764
R5505 VDD.n30 VDD.t135 21.1764
R5506 VDD.n29 VDD.t119 21.1764
R5507 VDD.n29 VDD.t151 21.1764
R5508 VDD.n25 VDD.t145 21.1764
R5509 VDD.n25 VDD.t139 21.1764
R5510 VDD.n23 VDD.t108 21.1764
R5511 VDD.n23 VDD.t123 21.1764
R5512 VDD.n22 VDD.t149 21.1764
R5513 VDD.n22 VDD.t142 21.1764
R5514 VDD.n19 VDD.t147 21.1764
R5515 VDD.n19 VDD.t140 21.1764
R5516 VDD.n17 VDD.t109 21.1764
R5517 VDD.n17 VDD.t125 21.1764
R5518 VDD.n16 VDD.t154 21.1764
R5519 VDD.n16 VDD.t143 21.1764
R5520 VDD.n2039 VDD.t115 21.1764
R5521 VDD.n2039 VDD.t117 21.1764
R5522 VDD.n2041 VDD.t136 21.1764
R5523 VDD.n2041 VDD.t111 21.1764
R5524 VDD.n2043 VDD.t121 21.1764
R5525 VDD.n2043 VDD.t127 21.1764
R5526 VDD.n2032 VDD.t133 21.1764
R5527 VDD.n2032 VDD.t156 21.1764
R5528 VDD.n2034 VDD.t132 21.1764
R5529 VDD.n2034 VDD.t150 21.1764
R5530 VDD.n2036 VDD.t124 21.1764
R5531 VDD.n2036 VDD.t148 21.1764
R5532 VDD.n2026 VDD.t137 21.1764
R5533 VDD.n2026 VDD.t103 21.1764
R5534 VDD.n2028 VDD.t134 21.1764
R5535 VDD.n2028 VDD.t155 21.1764
R5536 VDD.n2030 VDD.t130 21.1764
R5537 VDD.n2030 VDD.t153 21.1764
R5538 VDD.n2964 VDD.n1397 20.9278
R5539 VDD.n3385 VDD.n1036 20.9278
R5540 VDD.n3817 VDD.n3386 20.9278
R5541 VDD.n693 VDD.n679 20.9278
R5542 VDD.n2325 VDD.n2324 19.3944
R5543 VDD.n2324 VDD.n2285 19.3944
R5544 VDD.n2320 VDD.n2285 19.3944
R5545 VDD.n2320 VDD.n2319 19.3944
R5546 VDD.n2319 VDD.n2318 19.3944
R5547 VDD.n2318 VDD.n2291 19.3944
R5548 VDD.n2314 VDD.n2291 19.3944
R5549 VDD.n2314 VDD.n2313 19.3944
R5550 VDD.n2313 VDD.n2312 19.3944
R5551 VDD.n2312 VDD.n2297 19.3944
R5552 VDD.n2308 VDD.n2297 19.3944
R5553 VDD.n2308 VDD.n2307 19.3944
R5554 VDD.n2347 VDD.n2346 19.3944
R5555 VDD.n2346 VDD.n2345 19.3944
R5556 VDD.n2345 VDD.n2267 19.3944
R5557 VDD.n2341 VDD.n2267 19.3944
R5558 VDD.n2341 VDD.n2340 19.3944
R5559 VDD.n2340 VDD.n2339 19.3944
R5560 VDD.n2339 VDD.n2273 19.3944
R5561 VDD.n2335 VDD.n2273 19.3944
R5562 VDD.n2335 VDD.n2334 19.3944
R5563 VDD.n2334 VDD.n2333 19.3944
R5564 VDD.n2333 VDD.n2279 19.3944
R5565 VDD.n2329 VDD.n2279 19.3944
R5566 VDD.n2367 VDD.n2228 19.3944
R5567 VDD.n2362 VDD.n2228 19.3944
R5568 VDD.n2362 VDD.n2249 19.3944
R5569 VDD.n2358 VDD.n2249 19.3944
R5570 VDD.n2358 VDD.n2357 19.3944
R5571 VDD.n2357 VDD.n2356 19.3944
R5572 VDD.n2356 VDD.n2255 19.3944
R5573 VDD.n2352 VDD.n2255 19.3944
R5574 VDD.n2352 VDD.n2351 19.3944
R5575 VDD.n2351 VDD.n2350 19.3944
R5576 VDD.n2375 VDD.n2222 19.3944
R5577 VDD.n2375 VDD.n2220 19.3944
R5578 VDD.n2379 VDD.n2220 19.3944
R5579 VDD.n2379 VDD.n2209 19.3944
R5580 VDD.n2391 VDD.n2209 19.3944
R5581 VDD.n2391 VDD.n2207 19.3944
R5582 VDD.n2395 VDD.n2207 19.3944
R5583 VDD.n2395 VDD.n2198 19.3944
R5584 VDD.n2407 VDD.n2198 19.3944
R5585 VDD.n2407 VDD.n2196 19.3944
R5586 VDD.n2411 VDD.n2196 19.3944
R5587 VDD.n2411 VDD.n2186 19.3944
R5588 VDD.n2423 VDD.n2186 19.3944
R5589 VDD.n2423 VDD.n2184 19.3944
R5590 VDD.n2427 VDD.n2184 19.3944
R5591 VDD.n2427 VDD.n2174 19.3944
R5592 VDD.n2439 VDD.n2174 19.3944
R5593 VDD.n2439 VDD.n2172 19.3944
R5594 VDD.n2443 VDD.n2172 19.3944
R5595 VDD.n2443 VDD.n2162 19.3944
R5596 VDD.n2455 VDD.n2162 19.3944
R5597 VDD.n2455 VDD.n2160 19.3944
R5598 VDD.n2459 VDD.n2160 19.3944
R5599 VDD.n2459 VDD.n2150 19.3944
R5600 VDD.n2471 VDD.n2150 19.3944
R5601 VDD.n2471 VDD.n2148 19.3944
R5602 VDD.n2475 VDD.n2148 19.3944
R5603 VDD.n2475 VDD.n2138 19.3944
R5604 VDD.n2487 VDD.n2138 19.3944
R5605 VDD.n2487 VDD.n2136 19.3944
R5606 VDD.n2491 VDD.n2136 19.3944
R5607 VDD.n2491 VDD.n2126 19.3944
R5608 VDD.n2503 VDD.n2126 19.3944
R5609 VDD.n2503 VDD.n2124 19.3944
R5610 VDD.n2507 VDD.n2124 19.3944
R5611 VDD.n2507 VDD.n2114 19.3944
R5612 VDD.n2519 VDD.n2114 19.3944
R5613 VDD.n2519 VDD.n2112 19.3944
R5614 VDD.n2523 VDD.n2112 19.3944
R5615 VDD.n2523 VDD.n2102 19.3944
R5616 VDD.n2535 VDD.n2102 19.3944
R5617 VDD.n2535 VDD.n2100 19.3944
R5618 VDD.n2539 VDD.n2100 19.3944
R5619 VDD.n2539 VDD.n2089 19.3944
R5620 VDD.n2551 VDD.n2089 19.3944
R5621 VDD.n2551 VDD.n2087 19.3944
R5622 VDD.n2555 VDD.n2087 19.3944
R5623 VDD.n2555 VDD.n2078 19.3944
R5624 VDD.n2567 VDD.n2078 19.3944
R5625 VDD.n2567 VDD.n2076 19.3944
R5626 VDD.n2571 VDD.n2076 19.3944
R5627 VDD.n2571 VDD.n2066 19.3944
R5628 VDD.n2583 VDD.n2066 19.3944
R5629 VDD.n2583 VDD.n2064 19.3944
R5630 VDD.n2587 VDD.n2064 19.3944
R5631 VDD.n2587 VDD.n2053 19.3944
R5632 VDD.n2600 VDD.n2053 19.3944
R5633 VDD.n2600 VDD.n2051 19.3944
R5634 VDD.n2604 VDD.n2051 19.3944
R5635 VDD.n2604 VDD.n2021 19.3944
R5636 VDD.n2616 VDD.n2021 19.3944
R5637 VDD.n2616 VDD.n2019 19.3944
R5638 VDD.n2620 VDD.n2019 19.3944
R5639 VDD.n2620 VDD.n2009 19.3944
R5640 VDD.n2632 VDD.n2009 19.3944
R5641 VDD.n2632 VDD.n2007 19.3944
R5642 VDD.n2636 VDD.n2007 19.3944
R5643 VDD.n2636 VDD.n1996 19.3944
R5644 VDD.n2648 VDD.n1996 19.3944
R5645 VDD.n2648 VDD.n1994 19.3944
R5646 VDD.n2652 VDD.n1994 19.3944
R5647 VDD.n2652 VDD.n1985 19.3944
R5648 VDD.n2664 VDD.n1985 19.3944
R5649 VDD.n2664 VDD.n1983 19.3944
R5650 VDD.n2668 VDD.n1983 19.3944
R5651 VDD.n2668 VDD.n1973 19.3944
R5652 VDD.n2680 VDD.n1973 19.3944
R5653 VDD.n2680 VDD.n1971 19.3944
R5654 VDD.n2684 VDD.n1971 19.3944
R5655 VDD.n2684 VDD.n1961 19.3944
R5656 VDD.n2696 VDD.n1961 19.3944
R5657 VDD.n2696 VDD.n1959 19.3944
R5658 VDD.n2700 VDD.n1959 19.3944
R5659 VDD.n2700 VDD.n1949 19.3944
R5660 VDD.n2712 VDD.n1949 19.3944
R5661 VDD.n2712 VDD.n1947 19.3944
R5662 VDD.n2716 VDD.n1947 19.3944
R5663 VDD.n2716 VDD.n1937 19.3944
R5664 VDD.n2728 VDD.n1937 19.3944
R5665 VDD.n2728 VDD.n1935 19.3944
R5666 VDD.n2732 VDD.n1935 19.3944
R5667 VDD.n2732 VDD.n1925 19.3944
R5668 VDD.n2744 VDD.n1925 19.3944
R5669 VDD.n2744 VDD.n1923 19.3944
R5670 VDD.n2748 VDD.n1923 19.3944
R5671 VDD.n2748 VDD.n1913 19.3944
R5672 VDD.n2760 VDD.n1913 19.3944
R5673 VDD.n2760 VDD.n1911 19.3944
R5674 VDD.n2764 VDD.n1911 19.3944
R5675 VDD.n2764 VDD.n1901 19.3944
R5676 VDD.n2776 VDD.n1901 19.3944
R5677 VDD.n2776 VDD.n1899 19.3944
R5678 VDD.n2780 VDD.n1899 19.3944
R5679 VDD.n2780 VDD.n1889 19.3944
R5680 VDD.n2792 VDD.n1889 19.3944
R5681 VDD.n2792 VDD.n1887 19.3944
R5682 VDD.n2796 VDD.n1887 19.3944
R5683 VDD.n2796 VDD.n1876 19.3944
R5684 VDD.n2808 VDD.n1876 19.3944
R5685 VDD.n2808 VDD.n1873 19.3944
R5686 VDD.n2813 VDD.n1873 19.3944
R5687 VDD.n2813 VDD.n1874 19.3944
R5688 VDD.n1874 VDD.n1864 19.3944
R5689 VDD.n2826 VDD.n1864 19.3944
R5690 VDD.n2826 VDD.n1861 19.3944
R5691 VDD.n2832 VDD.n1861 19.3944
R5692 VDD.n2832 VDD.n1862 19.3944
R5693 VDD.n646 VDD.n573 19.3944
R5694 VDD.n650 VDD.n573 19.3944
R5695 VDD.n653 VDD.n650 19.3944
R5696 VDD.n656 VDD.n653 19.3944
R5697 VDD.n656 VDD.n571 19.3944
R5698 VDD.n660 VDD.n571 19.3944
R5699 VDD.n663 VDD.n660 19.3944
R5700 VDD.n666 VDD.n663 19.3944
R5701 VDD.n666 VDD.n569 19.3944
R5702 VDD.n670 VDD.n569 19.3944
R5703 VDD.n673 VDD.n670 19.3944
R5704 VDD.n674 VDD.n673 19.3944
R5705 VDD.n615 VDD.n612 19.3944
R5706 VDD.n615 VDD.n581 19.3944
R5707 VDD.n619 VDD.n581 19.3944
R5708 VDD.n622 VDD.n619 19.3944
R5709 VDD.n625 VDD.n622 19.3944
R5710 VDD.n625 VDD.n579 19.3944
R5711 VDD.n629 VDD.n579 19.3944
R5712 VDD.n632 VDD.n629 19.3944
R5713 VDD.n635 VDD.n632 19.3944
R5714 VDD.n635 VDD.n577 19.3944
R5715 VDD.n639 VDD.n577 19.3944
R5716 VDD.n642 VDD.n639 19.3944
R5717 VDD.n4246 VDD.n4245 19.3944
R5718 VDD.n4245 VDD.n545 19.3944
R5719 VDD.n592 VDD.n545 19.3944
R5720 VDD.n595 VDD.n592 19.3944
R5721 VDD.n595 VDD.n588 19.3944
R5722 VDD.n599 VDD.n588 19.3944
R5723 VDD.n602 VDD.n599 19.3944
R5724 VDD.n605 VDD.n602 19.3944
R5725 VDD.n605 VDD.n586 19.3944
R5726 VDD.n609 VDD.n586 19.3944
R5727 VDD.n4250 VDD.n540 19.3944
R5728 VDD.n4250 VDD.n530 19.3944
R5729 VDD.n4262 VDD.n530 19.3944
R5730 VDD.n4262 VDD.n528 19.3944
R5731 VDD.n4266 VDD.n528 19.3944
R5732 VDD.n4266 VDD.n518 19.3944
R5733 VDD.n4278 VDD.n518 19.3944
R5734 VDD.n4278 VDD.n516 19.3944
R5735 VDD.n4282 VDD.n516 19.3944
R5736 VDD.n4282 VDD.n506 19.3944
R5737 VDD.n4294 VDD.n506 19.3944
R5738 VDD.n4294 VDD.n504 19.3944
R5739 VDD.n4298 VDD.n504 19.3944
R5740 VDD.n4298 VDD.n494 19.3944
R5741 VDD.n4310 VDD.n494 19.3944
R5742 VDD.n4310 VDD.n492 19.3944
R5743 VDD.n4314 VDD.n492 19.3944
R5744 VDD.n4314 VDD.n482 19.3944
R5745 VDD.n4326 VDD.n482 19.3944
R5746 VDD.n4326 VDD.n480 19.3944
R5747 VDD.n4330 VDD.n480 19.3944
R5748 VDD.n4330 VDD.n470 19.3944
R5749 VDD.n4342 VDD.n470 19.3944
R5750 VDD.n4342 VDD.n468 19.3944
R5751 VDD.n4346 VDD.n468 19.3944
R5752 VDD.n4346 VDD.n458 19.3944
R5753 VDD.n4358 VDD.n458 19.3944
R5754 VDD.n4358 VDD.n456 19.3944
R5755 VDD.n4362 VDD.n456 19.3944
R5756 VDD.n4362 VDD.n446 19.3944
R5757 VDD.n4374 VDD.n446 19.3944
R5758 VDD.n4374 VDD.n444 19.3944
R5759 VDD.n4378 VDD.n444 19.3944
R5760 VDD.n4378 VDD.n434 19.3944
R5761 VDD.n4390 VDD.n434 19.3944
R5762 VDD.n4390 VDD.n432 19.3944
R5763 VDD.n4394 VDD.n432 19.3944
R5764 VDD.n4394 VDD.n422 19.3944
R5765 VDD.n4406 VDD.n422 19.3944
R5766 VDD.n4406 VDD.n420 19.3944
R5767 VDD.n4410 VDD.n420 19.3944
R5768 VDD.n4410 VDD.n410 19.3944
R5769 VDD.n4422 VDD.n410 19.3944
R5770 VDD.n4422 VDD.n408 19.3944
R5771 VDD.n4426 VDD.n408 19.3944
R5772 VDD.n4426 VDD.n398 19.3944
R5773 VDD.n4438 VDD.n398 19.3944
R5774 VDD.n4438 VDD.n396 19.3944
R5775 VDD.n4442 VDD.n396 19.3944
R5776 VDD.n4442 VDD.n386 19.3944
R5777 VDD.n4456 VDD.n386 19.3944
R5778 VDD.n4456 VDD.n384 19.3944
R5779 VDD.n4460 VDD.n384 19.3944
R5780 VDD.n4460 VDD.n374 19.3944
R5781 VDD.n4477 VDD.n374 19.3944
R5782 VDD.n4477 VDD.n372 19.3944
R5783 VDD.n4481 VDD.n372 19.3944
R5784 VDD.n4481 VDD.n38 19.3944
R5785 VDD.n4710 VDD.n38 19.3944
R5786 VDD.n4710 VDD.n4709 19.3944
R5787 VDD.n4709 VDD.n40 19.3944
R5788 VDD.n4703 VDD.n40 19.3944
R5789 VDD.n4703 VDD.n4702 19.3944
R5790 VDD.n4702 VDD.n4701 19.3944
R5791 VDD.n4701 VDD.n52 19.3944
R5792 VDD.n4695 VDD.n52 19.3944
R5793 VDD.n4695 VDD.n4694 19.3944
R5794 VDD.n4694 VDD.n4693 19.3944
R5795 VDD.n4693 VDD.n63 19.3944
R5796 VDD.n4687 VDD.n63 19.3944
R5797 VDD.n4687 VDD.n4686 19.3944
R5798 VDD.n4686 VDD.n4685 19.3944
R5799 VDD.n4685 VDD.n73 19.3944
R5800 VDD.n4679 VDD.n73 19.3944
R5801 VDD.n4679 VDD.n4678 19.3944
R5802 VDD.n4678 VDD.n4677 19.3944
R5803 VDD.n4677 VDD.n85 19.3944
R5804 VDD.n4671 VDD.n85 19.3944
R5805 VDD.n4671 VDD.n4670 19.3944
R5806 VDD.n4670 VDD.n4669 19.3944
R5807 VDD.n4669 VDD.n96 19.3944
R5808 VDD.n4663 VDD.n96 19.3944
R5809 VDD.n4663 VDD.n4662 19.3944
R5810 VDD.n4662 VDD.n4661 19.3944
R5811 VDD.n4661 VDD.n107 19.3944
R5812 VDD.n4655 VDD.n107 19.3944
R5813 VDD.n4655 VDD.n4654 19.3944
R5814 VDD.n4654 VDD.n4653 19.3944
R5815 VDD.n4653 VDD.n118 19.3944
R5816 VDD.n4647 VDD.n118 19.3944
R5817 VDD.n4647 VDD.n4646 19.3944
R5818 VDD.n4646 VDD.n4645 19.3944
R5819 VDD.n4645 VDD.n129 19.3944
R5820 VDD.n4639 VDD.n129 19.3944
R5821 VDD.n4639 VDD.n4638 19.3944
R5822 VDD.n4638 VDD.n4637 19.3944
R5823 VDD.n4637 VDD.n140 19.3944
R5824 VDD.n4631 VDD.n140 19.3944
R5825 VDD.n4631 VDD.n4630 19.3944
R5826 VDD.n4630 VDD.n4629 19.3944
R5827 VDD.n4629 VDD.n151 19.3944
R5828 VDD.n4623 VDD.n151 19.3944
R5829 VDD.n4623 VDD.n4622 19.3944
R5830 VDD.n4622 VDD.n4621 19.3944
R5831 VDD.n4621 VDD.n162 19.3944
R5832 VDD.n4615 VDD.n162 19.3944
R5833 VDD.n4615 VDD.n4614 19.3944
R5834 VDD.n4614 VDD.n4613 19.3944
R5835 VDD.n4613 VDD.n173 19.3944
R5836 VDD.n4607 VDD.n173 19.3944
R5837 VDD.n4607 VDD.n4606 19.3944
R5838 VDD.n4606 VDD.n4605 19.3944
R5839 VDD.n4605 VDD.n183 19.3944
R5840 VDD.n4599 VDD.n183 19.3944
R5841 VDD.n4599 VDD.n4598 19.3944
R5842 VDD.n4598 VDD.n4597 19.3944
R5843 VDD.n4597 VDD.n195 19.3944
R5844 VDD.n307 VDD.n226 19.3944
R5845 VDD.n313 VDD.n226 19.3944
R5846 VDD.n314 VDD.n313 19.3944
R5847 VDD.n317 VDD.n314 19.3944
R5848 VDD.n317 VDD.n224 19.3944
R5849 VDD.n323 VDD.n224 19.3944
R5850 VDD.n324 VDD.n323 19.3944
R5851 VDD.n327 VDD.n324 19.3944
R5852 VDD.n327 VDD.n222 19.3944
R5853 VDD.n333 VDD.n222 19.3944
R5854 VDD.n335 VDD.n333 19.3944
R5855 VDD.n336 VDD.n335 19.3944
R5856 VDD.n277 VDD.n274 19.3944
R5857 VDD.n277 VDD.n235 19.3944
R5858 VDD.n283 VDD.n235 19.3944
R5859 VDD.n284 VDD.n283 19.3944
R5860 VDD.n287 VDD.n284 19.3944
R5861 VDD.n287 VDD.n233 19.3944
R5862 VDD.n293 VDD.n233 19.3944
R5863 VDD.n294 VDD.n293 19.3944
R5864 VDD.n297 VDD.n294 19.3944
R5865 VDD.n297 VDD.n231 19.3944
R5866 VDD.n303 VDD.n231 19.3944
R5867 VDD.n304 VDD.n303 19.3944
R5868 VDD.n246 VDD.n243 19.3944
R5869 VDD.n252 VDD.n243 19.3944
R5870 VDD.n253 VDD.n252 19.3944
R5871 VDD.n256 VDD.n253 19.3944
R5872 VDD.n256 VDD.n241 19.3944
R5873 VDD.n262 VDD.n241 19.3944
R5874 VDD.n263 VDD.n262 19.3944
R5875 VDD.n266 VDD.n263 19.3944
R5876 VDD.n266 VDD.n239 19.3944
R5877 VDD.n272 VDD.n239 19.3944
R5878 VDD.n4254 VDD.n536 19.3944
R5879 VDD.n4254 VDD.n534 19.3944
R5880 VDD.n4258 VDD.n534 19.3944
R5881 VDD.n4258 VDD.n523 19.3944
R5882 VDD.n4270 VDD.n523 19.3944
R5883 VDD.n4270 VDD.n521 19.3944
R5884 VDD.n4274 VDD.n521 19.3944
R5885 VDD.n4274 VDD.n512 19.3944
R5886 VDD.n4286 VDD.n512 19.3944
R5887 VDD.n4286 VDD.n510 19.3944
R5888 VDD.n4290 VDD.n510 19.3944
R5889 VDD.n4290 VDD.n500 19.3944
R5890 VDD.n4302 VDD.n500 19.3944
R5891 VDD.n4302 VDD.n498 19.3944
R5892 VDD.n4306 VDD.n498 19.3944
R5893 VDD.n4306 VDD.n488 19.3944
R5894 VDD.n4318 VDD.n488 19.3944
R5895 VDD.n4318 VDD.n486 19.3944
R5896 VDD.n4322 VDD.n486 19.3944
R5897 VDD.n4322 VDD.n476 19.3944
R5898 VDD.n4334 VDD.n476 19.3944
R5899 VDD.n4334 VDD.n474 19.3944
R5900 VDD.n4338 VDD.n474 19.3944
R5901 VDD.n4338 VDD.n464 19.3944
R5902 VDD.n4350 VDD.n464 19.3944
R5903 VDD.n4350 VDD.n462 19.3944
R5904 VDD.n4354 VDD.n462 19.3944
R5905 VDD.n4354 VDD.n452 19.3944
R5906 VDD.n4366 VDD.n452 19.3944
R5907 VDD.n4366 VDD.n450 19.3944
R5908 VDD.n4370 VDD.n450 19.3944
R5909 VDD.n4370 VDD.n440 19.3944
R5910 VDD.n4382 VDD.n440 19.3944
R5911 VDD.n4382 VDD.n438 19.3944
R5912 VDD.n4386 VDD.n438 19.3944
R5913 VDD.n4386 VDD.n428 19.3944
R5914 VDD.n4398 VDD.n428 19.3944
R5915 VDD.n4398 VDD.n426 19.3944
R5916 VDD.n4402 VDD.n426 19.3944
R5917 VDD.n4402 VDD.n416 19.3944
R5918 VDD.n4414 VDD.n416 19.3944
R5919 VDD.n4414 VDD.n414 19.3944
R5920 VDD.n4418 VDD.n414 19.3944
R5921 VDD.n4418 VDD.n403 19.3944
R5922 VDD.n4430 VDD.n403 19.3944
R5923 VDD.n4430 VDD.n401 19.3944
R5924 VDD.n4434 VDD.n401 19.3944
R5925 VDD.n4434 VDD.n392 19.3944
R5926 VDD.n4446 VDD.n392 19.3944
R5927 VDD.n4446 VDD.n390 19.3944
R5928 VDD.n4452 VDD.n390 19.3944
R5929 VDD.n4452 VDD.n4451 19.3944
R5930 VDD.n4451 VDD.n380 19.3944
R5931 VDD.n4465 VDD.n380 19.3944
R5932 VDD.n4465 VDD.n378 19.3944
R5933 VDD.n4472 VDD.n378 19.3944
R5934 VDD.n4472 VDD.n4471 19.3944
R5935 VDD.n4471 VDD.n367 19.3944
R5936 VDD.n4487 VDD.n367 19.3944
R5937 VDD.n4488 VDD.n4487 19.3944
R5938 VDD.n4489 VDD.n4488 19.3944
R5939 VDD.n4489 VDD.n365 19.3944
R5940 VDD.n4494 VDD.n365 19.3944
R5941 VDD.n4495 VDD.n4494 19.3944
R5942 VDD.n4496 VDD.n4495 19.3944
R5943 VDD.n4496 VDD.n363 19.3944
R5944 VDD.n4501 VDD.n363 19.3944
R5945 VDD.n4502 VDD.n4501 19.3944
R5946 VDD.n4503 VDD.n4502 19.3944
R5947 VDD.n4503 VDD.n361 19.3944
R5948 VDD.n4508 VDD.n361 19.3944
R5949 VDD.n4509 VDD.n4508 19.3944
R5950 VDD.n4510 VDD.n4509 19.3944
R5951 VDD.n4510 VDD.n359 19.3944
R5952 VDD.n4515 VDD.n359 19.3944
R5953 VDD.n4516 VDD.n4515 19.3944
R5954 VDD.n4517 VDD.n4516 19.3944
R5955 VDD.n4517 VDD.n357 19.3944
R5956 VDD.n4522 VDD.n357 19.3944
R5957 VDD.n4523 VDD.n4522 19.3944
R5958 VDD.n4524 VDD.n4523 19.3944
R5959 VDD.n4524 VDD.n355 19.3944
R5960 VDD.n4529 VDD.n355 19.3944
R5961 VDD.n4530 VDD.n4529 19.3944
R5962 VDD.n4531 VDD.n4530 19.3944
R5963 VDD.n4531 VDD.n353 19.3944
R5964 VDD.n4536 VDD.n353 19.3944
R5965 VDD.n4537 VDD.n4536 19.3944
R5966 VDD.n4538 VDD.n4537 19.3944
R5967 VDD.n4538 VDD.n351 19.3944
R5968 VDD.n4543 VDD.n351 19.3944
R5969 VDD.n4544 VDD.n4543 19.3944
R5970 VDD.n4545 VDD.n4544 19.3944
R5971 VDD.n4545 VDD.n349 19.3944
R5972 VDD.n4550 VDD.n349 19.3944
R5973 VDD.n4551 VDD.n4550 19.3944
R5974 VDD.n4552 VDD.n4551 19.3944
R5975 VDD.n4552 VDD.n347 19.3944
R5976 VDD.n4557 VDD.n347 19.3944
R5977 VDD.n4558 VDD.n4557 19.3944
R5978 VDD.n4559 VDD.n4558 19.3944
R5979 VDD.n4559 VDD.n345 19.3944
R5980 VDD.n4564 VDD.n345 19.3944
R5981 VDD.n4565 VDD.n4564 19.3944
R5982 VDD.n4566 VDD.n4565 19.3944
R5983 VDD.n4566 VDD.n343 19.3944
R5984 VDD.n4571 VDD.n343 19.3944
R5985 VDD.n4572 VDD.n4571 19.3944
R5986 VDD.n4573 VDD.n4572 19.3944
R5987 VDD.n4573 VDD.n341 19.3944
R5988 VDD.n4578 VDD.n341 19.3944
R5989 VDD.n4579 VDD.n4578 19.3944
R5990 VDD.n4580 VDD.n4579 19.3944
R5991 VDD.n4580 VDD.n339 19.3944
R5992 VDD.n4585 VDD.n339 19.3944
R5993 VDD.n4586 VDD.n4585 19.3944
R5994 VDD.n4587 VDD.n4586 19.3944
R5995 VDD.n2847 VDD.n2844 19.3944
R5996 VDD.n2850 VDD.n2847 19.3944
R5997 VDD.n2853 VDD.n2850 19.3944
R5998 VDD.n2853 VDD.n1852 19.3944
R5999 VDD.n2857 VDD.n1852 19.3944
R6000 VDD.n2860 VDD.n2857 19.3944
R6001 VDD.n2863 VDD.n2860 19.3944
R6002 VDD.n2863 VDD.n1850 19.3944
R6003 VDD.n2867 VDD.n1850 19.3944
R6004 VDD.n2870 VDD.n2867 19.3944
R6005 VDD.n2876 VDD.n1848 19.3944
R6006 VDD.n2880 VDD.n1848 19.3944
R6007 VDD.n2883 VDD.n2880 19.3944
R6008 VDD.n2886 VDD.n2883 19.3944
R6009 VDD.n2886 VDD.n1846 19.3944
R6010 VDD.n2890 VDD.n1846 19.3944
R6011 VDD.n2890 VDD.n1807 19.3944
R6012 VDD.n2937 VDD.n1807 19.3944
R6013 VDD.n2937 VDD.n2936 19.3944
R6014 VDD.n2936 VDD.n2935 19.3944
R6015 VDD.n2935 VDD.n1811 19.3944
R6016 VDD.n2931 VDD.n1811 19.3944
R6017 VDD.n2929 VDD.n2928 19.3944
R6018 VDD.n2928 VDD.n1818 19.3944
R6019 VDD.n2924 VDD.n1818 19.3944
R6020 VDD.n2924 VDD.n2923 19.3944
R6021 VDD.n2923 VDD.n2922 19.3944
R6022 VDD.n2922 VDD.n1823 19.3944
R6023 VDD.n2918 VDD.n1823 19.3944
R6024 VDD.n2918 VDD.n2917 19.3944
R6025 VDD.n2917 VDD.n2916 19.3944
R6026 VDD.n2916 VDD.n1828 19.3944
R6027 VDD.n2912 VDD.n1828 19.3944
R6028 VDD.n2912 VDD.n2911 19.3944
R6029 VDD.n2371 VDD.n2226 19.3944
R6030 VDD.n2371 VDD.n2216 19.3944
R6031 VDD.n2383 VDD.n2216 19.3944
R6032 VDD.n2383 VDD.n2214 19.3944
R6033 VDD.n2387 VDD.n2214 19.3944
R6034 VDD.n2387 VDD.n2204 19.3944
R6035 VDD.n2399 VDD.n2204 19.3944
R6036 VDD.n2399 VDD.n2202 19.3944
R6037 VDD.n2403 VDD.n2202 19.3944
R6038 VDD.n2403 VDD.n2192 19.3944
R6039 VDD.n2415 VDD.n2192 19.3944
R6040 VDD.n2415 VDD.n2190 19.3944
R6041 VDD.n2419 VDD.n2190 19.3944
R6042 VDD.n2419 VDD.n2180 19.3944
R6043 VDD.n2431 VDD.n2180 19.3944
R6044 VDD.n2431 VDD.n2178 19.3944
R6045 VDD.n2435 VDD.n2178 19.3944
R6046 VDD.n2435 VDD.n2168 19.3944
R6047 VDD.n2447 VDD.n2168 19.3944
R6048 VDD.n2447 VDD.n2166 19.3944
R6049 VDD.n2451 VDD.n2166 19.3944
R6050 VDD.n2451 VDD.n2156 19.3944
R6051 VDD.n2463 VDD.n2156 19.3944
R6052 VDD.n2463 VDD.n2154 19.3944
R6053 VDD.n2467 VDD.n2154 19.3944
R6054 VDD.n2467 VDD.n2144 19.3944
R6055 VDD.n2479 VDD.n2144 19.3944
R6056 VDD.n2479 VDD.n2142 19.3944
R6057 VDD.n2483 VDD.n2142 19.3944
R6058 VDD.n2483 VDD.n2132 19.3944
R6059 VDD.n2495 VDD.n2132 19.3944
R6060 VDD.n2495 VDD.n2130 19.3944
R6061 VDD.n2499 VDD.n2130 19.3944
R6062 VDD.n2499 VDD.n2120 19.3944
R6063 VDD.n2511 VDD.n2120 19.3944
R6064 VDD.n2511 VDD.n2118 19.3944
R6065 VDD.n2515 VDD.n2118 19.3944
R6066 VDD.n2515 VDD.n2108 19.3944
R6067 VDD.n2527 VDD.n2108 19.3944
R6068 VDD.n2527 VDD.n2106 19.3944
R6069 VDD.n2531 VDD.n2106 19.3944
R6070 VDD.n2531 VDD.n2096 19.3944
R6071 VDD.n2543 VDD.n2096 19.3944
R6072 VDD.n2543 VDD.n2094 19.3944
R6073 VDD.n2547 VDD.n2094 19.3944
R6074 VDD.n2547 VDD.n2084 19.3944
R6075 VDD.n2559 VDD.n2084 19.3944
R6076 VDD.n2559 VDD.n2082 19.3944
R6077 VDD.n2563 VDD.n2082 19.3944
R6078 VDD.n2563 VDD.n2072 19.3944
R6079 VDD.n2575 VDD.n2072 19.3944
R6080 VDD.n2575 VDD.n2070 19.3944
R6081 VDD.n2579 VDD.n2070 19.3944
R6082 VDD.n2579 VDD.n2060 19.3944
R6083 VDD.n2591 VDD.n2060 19.3944
R6084 VDD.n2591 VDD.n2058 19.3944
R6085 VDD.n2596 VDD.n2058 19.3944
R6086 VDD.n2596 VDD.n2048 19.3944
R6087 VDD.n2608 VDD.n2048 19.3944
R6088 VDD.n2608 VDD.n2025 19.3944
R6089 VDD.n2612 VDD.n2025 19.3944
R6090 VDD.n2612 VDD.n2015 19.3944
R6091 VDD.n2624 VDD.n2015 19.3944
R6092 VDD.n2624 VDD.n2013 19.3944
R6093 VDD.n2628 VDD.n2013 19.3944
R6094 VDD.n2628 VDD.n2003 19.3944
R6095 VDD.n2640 VDD.n2003 19.3944
R6096 VDD.n2640 VDD.n2001 19.3944
R6097 VDD.n2644 VDD.n2001 19.3944
R6098 VDD.n2644 VDD.n1991 19.3944
R6099 VDD.n2656 VDD.n1991 19.3944
R6100 VDD.n2656 VDD.n1989 19.3944
R6101 VDD.n2660 VDD.n1989 19.3944
R6102 VDD.n2660 VDD.n1979 19.3944
R6103 VDD.n2672 VDD.n1979 19.3944
R6104 VDD.n2672 VDD.n1977 19.3944
R6105 VDD.n2676 VDD.n1977 19.3944
R6106 VDD.n2676 VDD.n1967 19.3944
R6107 VDD.n2688 VDD.n1967 19.3944
R6108 VDD.n2688 VDD.n1965 19.3944
R6109 VDD.n2692 VDD.n1965 19.3944
R6110 VDD.n2692 VDD.n1955 19.3944
R6111 VDD.n2704 VDD.n1955 19.3944
R6112 VDD.n2704 VDD.n1953 19.3944
R6113 VDD.n2708 VDD.n1953 19.3944
R6114 VDD.n2708 VDD.n1943 19.3944
R6115 VDD.n2720 VDD.n1943 19.3944
R6116 VDD.n2720 VDD.n1941 19.3944
R6117 VDD.n2724 VDD.n1941 19.3944
R6118 VDD.n2724 VDD.n1931 19.3944
R6119 VDD.n2736 VDD.n1931 19.3944
R6120 VDD.n2736 VDD.n1929 19.3944
R6121 VDD.n2740 VDD.n1929 19.3944
R6122 VDD.n2740 VDD.n1919 19.3944
R6123 VDD.n2752 VDD.n1919 19.3944
R6124 VDD.n2752 VDD.n1917 19.3944
R6125 VDD.n2756 VDD.n1917 19.3944
R6126 VDD.n2756 VDD.n1907 19.3944
R6127 VDD.n2768 VDD.n1907 19.3944
R6128 VDD.n2768 VDD.n1905 19.3944
R6129 VDD.n2772 VDD.n1905 19.3944
R6130 VDD.n2772 VDD.n1895 19.3944
R6131 VDD.n2784 VDD.n1895 19.3944
R6132 VDD.n2784 VDD.n1893 19.3944
R6133 VDD.n2788 VDD.n1893 19.3944
R6134 VDD.n2788 VDD.n1883 19.3944
R6135 VDD.n2800 VDD.n1883 19.3944
R6136 VDD.n2800 VDD.n1881 19.3944
R6137 VDD.n2804 VDD.n1881 19.3944
R6138 VDD.n2804 VDD.n1870 19.3944
R6139 VDD.n2817 VDD.n1870 19.3944
R6140 VDD.n2817 VDD.n1868 19.3944
R6141 VDD.n2821 VDD.n1868 19.3944
R6142 VDD.n2821 VDD.n1857 19.3944
R6143 VDD.n2837 VDD.n1857 19.3944
R6144 VDD.n2837 VDD.n1855 19.3944
R6145 VDD.n2841 VDD.n1855 19.3944
R6146 VDD.n7 VDD.t88 16.9744
R6147 VDD.n7 VDD.t163 16.9744
R6148 VDD.n8 VDD.t159 16.9744
R6149 VDD.n8 VDD.t1 16.9744
R6150 VDD.n10 VDD.t83 16.9744
R6151 VDD.n10 VDD.t93 16.9744
R6152 VDD.n12 VDD.t77 16.9744
R6153 VDD.n12 VDD.t99 16.9744
R6154 VDD.n5 VDD.t101 16.9744
R6155 VDD.n5 VDD.t86 16.9744
R6156 VDD.n3 VDD.t95 16.9744
R6157 VDD.n3 VDD.t97 16.9744
R6158 VDD.n1 VDD.t90 16.9744
R6159 VDD.n1 VDD.t161 16.9744
R6160 VDD.n0 VDD.t79 16.9744
R6161 VDD.n0 VDD.t75 16.9744
R6162 VDD.n2373 VDD.n2224 16.2232
R6163 VDD.n2373 VDD.n2218 16.2232
R6164 VDD.n2381 VDD.n2218 16.2232
R6165 VDD.n2381 VDD.n2211 16.2232
R6166 VDD.n2389 VDD.n2211 16.2232
R6167 VDD.n2389 VDD.n2212 16.2232
R6168 VDD.n2397 VDD.n2200 16.2232
R6169 VDD.n2405 VDD.n2200 16.2232
R6170 VDD.n2405 VDD.n2194 16.2232
R6171 VDD.n2413 VDD.n2194 16.2232
R6172 VDD.n2413 VDD.n2188 16.2232
R6173 VDD.n2421 VDD.n2188 16.2232
R6174 VDD.n2421 VDD.n2182 16.2232
R6175 VDD.n2429 VDD.n2182 16.2232
R6176 VDD.n2429 VDD.n2176 16.2232
R6177 VDD.n2437 VDD.n2176 16.2232
R6178 VDD.n2437 VDD.n2170 16.2232
R6179 VDD.n2445 VDD.n2170 16.2232
R6180 VDD.n2445 VDD.n2164 16.2232
R6181 VDD.n2453 VDD.n2164 16.2232
R6182 VDD.n2461 VDD.n2158 16.2232
R6183 VDD.n2461 VDD.n2152 16.2232
R6184 VDD.n2469 VDD.n2152 16.2232
R6185 VDD.n2469 VDD.n2146 16.2232
R6186 VDD.n2477 VDD.n2146 16.2232
R6187 VDD.n2477 VDD.n2140 16.2232
R6188 VDD.n2485 VDD.n2140 16.2232
R6189 VDD.n2485 VDD.n2134 16.2232
R6190 VDD.n2493 VDD.n2134 16.2232
R6191 VDD.n2493 VDD.n2128 16.2232
R6192 VDD.n2501 VDD.n2128 16.2232
R6193 VDD.n2509 VDD.n2122 16.2232
R6194 VDD.n2509 VDD.n2116 16.2232
R6195 VDD.n2517 VDD.n2116 16.2232
R6196 VDD.n2517 VDD.n2110 16.2232
R6197 VDD.n2525 VDD.n2110 16.2232
R6198 VDD.n2525 VDD.n2104 16.2232
R6199 VDD.n2533 VDD.n2104 16.2232
R6200 VDD.n2533 VDD.n2098 16.2232
R6201 VDD.n2541 VDD.n2098 16.2232
R6202 VDD.n2541 VDD.n2091 16.2232
R6203 VDD.n2549 VDD.n2091 16.2232
R6204 VDD.n2549 VDD.n2092 16.2232
R6205 VDD.n2557 VDD.n2080 16.2232
R6206 VDD.n2565 VDD.n2080 16.2232
R6207 VDD.n2565 VDD.n2074 16.2232
R6208 VDD.n2573 VDD.n2074 16.2232
R6209 VDD.n2573 VDD.n2068 16.2232
R6210 VDD.n2581 VDD.n2068 16.2232
R6211 VDD.n2581 VDD.n2062 16.2232
R6212 VDD.n2589 VDD.n2062 16.2232
R6213 VDD.n2589 VDD.n2055 16.2232
R6214 VDD.n2598 VDD.n2055 16.2232
R6215 VDD.n2598 VDD.n2056 16.2232
R6216 VDD.n2606 VDD.n2023 16.2232
R6217 VDD.n2614 VDD.n2023 16.2232
R6218 VDD.n2614 VDD.n2017 16.2232
R6219 VDD.n2622 VDD.n2017 16.2232
R6220 VDD.n2622 VDD.n2011 16.2232
R6221 VDD.n2630 VDD.n2011 16.2232
R6222 VDD.n2630 VDD.n2005 16.2232
R6223 VDD.n2638 VDD.n2005 16.2232
R6224 VDD.n2638 VDD.n1998 16.2232
R6225 VDD.n2646 VDD.n1998 16.2232
R6226 VDD.n2646 VDD.n1999 16.2232
R6227 VDD.n2654 VDD.n1987 16.2232
R6228 VDD.n2662 VDD.n1987 16.2232
R6229 VDD.n2662 VDD.n1981 16.2232
R6230 VDD.n2670 VDD.n1981 16.2232
R6231 VDD.n2670 VDD.n1975 16.2232
R6232 VDD.n2678 VDD.n1975 16.2232
R6233 VDD.n2678 VDD.n1969 16.2232
R6234 VDD.n2686 VDD.n1969 16.2232
R6235 VDD.n2686 VDD.n1963 16.2232
R6236 VDD.n2694 VDD.n1963 16.2232
R6237 VDD.n2694 VDD.n1957 16.2232
R6238 VDD.n2702 VDD.n1957 16.2232
R6239 VDD.n2710 VDD.n1951 16.2232
R6240 VDD.n2710 VDD.n1945 16.2232
R6241 VDD.n2718 VDD.n1945 16.2232
R6242 VDD.n2718 VDD.n1939 16.2232
R6243 VDD.n2726 VDD.n1939 16.2232
R6244 VDD.n2726 VDD.n1933 16.2232
R6245 VDD.n2734 VDD.n1933 16.2232
R6246 VDD.n2734 VDD.n1927 16.2232
R6247 VDD.n2742 VDD.n1927 16.2232
R6248 VDD.n2742 VDD.n1921 16.2232
R6249 VDD.n2750 VDD.n1921 16.2232
R6250 VDD.n2758 VDD.n1915 16.2232
R6251 VDD.n2758 VDD.n1909 16.2232
R6252 VDD.n2766 VDD.n1909 16.2232
R6253 VDD.n2766 VDD.n1903 16.2232
R6254 VDD.n2774 VDD.n1903 16.2232
R6255 VDD.n2774 VDD.n1897 16.2232
R6256 VDD.n2782 VDD.n1897 16.2232
R6257 VDD.n2782 VDD.n1891 16.2232
R6258 VDD.n2790 VDD.n1891 16.2232
R6259 VDD.n2790 VDD.n1885 16.2232
R6260 VDD.n2798 VDD.n1885 16.2232
R6261 VDD.n2798 VDD.n1878 16.2232
R6262 VDD.n2806 VDD.n1878 16.2232
R6263 VDD.n2806 VDD.n1879 16.2232
R6264 VDD.n2815 VDD.n1866 16.2232
R6265 VDD.n2823 VDD.n1866 16.2232
R6266 VDD.n2823 VDD.n1859 16.2232
R6267 VDD.n2835 VDD.n1859 16.2232
R6268 VDD.n2835 VDD.n2834 16.2232
R6269 VDD.n2834 VDD.n1836 16.2232
R6270 VDD.n4252 VDD.n538 16.2232
R6271 VDD.n4252 VDD.n532 16.2232
R6272 VDD.n4260 VDD.n532 16.2232
R6273 VDD.n4260 VDD.n525 16.2232
R6274 VDD.n4268 VDD.n525 16.2232
R6275 VDD.n4268 VDD.n526 16.2232
R6276 VDD.n4276 VDD.n514 16.2232
R6277 VDD.n4284 VDD.n514 16.2232
R6278 VDD.n4284 VDD.n508 16.2232
R6279 VDD.n4292 VDD.n508 16.2232
R6280 VDD.n4292 VDD.n502 16.2232
R6281 VDD.n4300 VDD.n502 16.2232
R6282 VDD.n4300 VDD.n496 16.2232
R6283 VDD.n4308 VDD.n496 16.2232
R6284 VDD.n4308 VDD.n490 16.2232
R6285 VDD.n4316 VDD.n490 16.2232
R6286 VDD.n4316 VDD.n484 16.2232
R6287 VDD.n4324 VDD.n484 16.2232
R6288 VDD.n4324 VDD.n478 16.2232
R6289 VDD.n4332 VDD.n478 16.2232
R6290 VDD.n4340 VDD.n472 16.2232
R6291 VDD.n4340 VDD.n466 16.2232
R6292 VDD.n4348 VDD.n466 16.2232
R6293 VDD.n4348 VDD.n460 16.2232
R6294 VDD.n4356 VDD.n460 16.2232
R6295 VDD.n4356 VDD.n454 16.2232
R6296 VDD.n4364 VDD.n454 16.2232
R6297 VDD.n4364 VDD.n448 16.2232
R6298 VDD.n4372 VDD.n448 16.2232
R6299 VDD.n4372 VDD.n442 16.2232
R6300 VDD.n4380 VDD.n442 16.2232
R6301 VDD.n4388 VDD.n436 16.2232
R6302 VDD.n4388 VDD.n430 16.2232
R6303 VDD.n4396 VDD.n430 16.2232
R6304 VDD.n4396 VDD.n424 16.2232
R6305 VDD.n4404 VDD.n424 16.2232
R6306 VDD.n4404 VDD.n418 16.2232
R6307 VDD.n4412 VDD.n418 16.2232
R6308 VDD.n4412 VDD.n412 16.2232
R6309 VDD.n4420 VDD.n412 16.2232
R6310 VDD.n4420 VDD.n405 16.2232
R6311 VDD.n4428 VDD.n405 16.2232
R6312 VDD.n4428 VDD.n406 16.2232
R6313 VDD.n4436 VDD.n394 16.2232
R6314 VDD.n4444 VDD.n394 16.2232
R6315 VDD.n4444 VDD.n388 16.2232
R6316 VDD.n4454 VDD.n388 16.2232
R6317 VDD.n4454 VDD.n382 16.2232
R6318 VDD.n4462 VDD.n382 16.2232
R6319 VDD.n4462 VDD.n376 16.2232
R6320 VDD.n4475 VDD.n376 16.2232
R6321 VDD.n4475 VDD.n4474 16.2232
R6322 VDD.n4474 VDD.n370 16.2232
R6323 VDD.n4484 VDD.n370 16.2232
R6324 VDD.n4707 VDD.n42 16.2232
R6325 VDD.n4707 VDD.n4706 16.2232
R6326 VDD.n4706 VDD.n4705 16.2232
R6327 VDD.n4705 VDD.n46 16.2232
R6328 VDD.n4699 VDD.n46 16.2232
R6329 VDD.n4699 VDD.n4698 16.2232
R6330 VDD.n4698 VDD.n4697 16.2232
R6331 VDD.n4697 VDD.n57 16.2232
R6332 VDD.n4691 VDD.n57 16.2232
R6333 VDD.n4691 VDD.n4690 16.2232
R6334 VDD.n4690 VDD.n4689 16.2232
R6335 VDD.n4683 VDD.n75 16.2232
R6336 VDD.n4683 VDD.n4682 16.2232
R6337 VDD.n4682 VDD.n4681 16.2232
R6338 VDD.n4681 VDD.n79 16.2232
R6339 VDD.n4675 VDD.n79 16.2232
R6340 VDD.n4675 VDD.n4674 16.2232
R6341 VDD.n4674 VDD.n4673 16.2232
R6342 VDD.n4673 VDD.n90 16.2232
R6343 VDD.n4667 VDD.n90 16.2232
R6344 VDD.n4667 VDD.n4666 16.2232
R6345 VDD.n4666 VDD.n4665 16.2232
R6346 VDD.n4665 VDD.n101 16.2232
R6347 VDD.n4659 VDD.n4658 16.2232
R6348 VDD.n4658 VDD.n4657 16.2232
R6349 VDD.n4657 VDD.n112 16.2232
R6350 VDD.n4651 VDD.n112 16.2232
R6351 VDD.n4651 VDD.n4650 16.2232
R6352 VDD.n4650 VDD.n4649 16.2232
R6353 VDD.n4649 VDD.n123 16.2232
R6354 VDD.n4643 VDD.n123 16.2232
R6355 VDD.n4643 VDD.n4642 16.2232
R6356 VDD.n4642 VDD.n4641 16.2232
R6357 VDD.n4641 VDD.n134 16.2232
R6358 VDD.n4635 VDD.n4634 16.2232
R6359 VDD.n4634 VDD.n4633 16.2232
R6360 VDD.n4633 VDD.n145 16.2232
R6361 VDD.n4627 VDD.n145 16.2232
R6362 VDD.n4627 VDD.n4626 16.2232
R6363 VDD.n4626 VDD.n4625 16.2232
R6364 VDD.n4625 VDD.n156 16.2232
R6365 VDD.n4619 VDD.n156 16.2232
R6366 VDD.n4619 VDD.n4618 16.2232
R6367 VDD.n4618 VDD.n4617 16.2232
R6368 VDD.n4617 VDD.n167 16.2232
R6369 VDD.n4611 VDD.n167 16.2232
R6370 VDD.n4611 VDD.n4610 16.2232
R6371 VDD.n4610 VDD.n4609 16.2232
R6372 VDD.n4603 VDD.n185 16.2232
R6373 VDD.n4603 VDD.n4602 16.2232
R6374 VDD.n4602 VDD.n4601 16.2232
R6375 VDD.n4601 VDD.n189 16.2232
R6376 VDD.n4595 VDD.n189 16.2232
R6377 VDD.n4595 VDD.n4594 16.2232
R6378 VDD.n2501 VDD.t126 14.6009
R6379 VDD.t102 VDD.n1951 14.6009
R6380 VDD.n4380 VDD.t141 14.6009
R6381 VDD.n4659 VDD.t138 14.6009
R6382 VDD.n2557 VDD.t131 12.9786
R6383 VDD.n1999 VDD.t114 12.9786
R6384 VDD.n4436 VDD.t107 12.9786
R6385 VDD.n4689 VDD.t128 12.9786
R6386 VDD.n4190 VDD.n542 11.2946
R6387 VDD.n4238 VDD.n4237 11.2946
R6388 VDD.n2941 VDD.n2940 11.2942
R6389 VDD.n1804 VDD.n1803 11.2942
R6390 VDD.n2964 VDD.n1391 11.0319
R6391 VDD.n2970 VDD.n1391 11.0319
R6392 VDD.n2970 VDD.n1385 11.0319
R6393 VDD.n2976 VDD.n1385 11.0319
R6394 VDD.n2976 VDD.n1379 11.0319
R6395 VDD.n2982 VDD.n1379 11.0319
R6396 VDD.n2982 VDD.n1373 11.0319
R6397 VDD.n2988 VDD.n1373 11.0319
R6398 VDD.n2994 VDD.n1366 11.0319
R6399 VDD.n2994 VDD.n1369 11.0319
R6400 VDD.n3000 VDD.n1355 11.0319
R6401 VDD.n3006 VDD.n1355 11.0319
R6402 VDD.n3006 VDD.n1349 11.0319
R6403 VDD.n3012 VDD.n1349 11.0319
R6404 VDD.n3012 VDD.n1343 11.0319
R6405 VDD.n3018 VDD.n1343 11.0319
R6406 VDD.n3018 VDD.n1337 11.0319
R6407 VDD.n3024 VDD.n1337 11.0319
R6408 VDD.n3024 VDD.n1331 11.0319
R6409 VDD.n3030 VDD.n1331 11.0319
R6410 VDD.n3030 VDD.n1325 11.0319
R6411 VDD.n3036 VDD.n1325 11.0319
R6412 VDD.n3036 VDD.n1319 11.0319
R6413 VDD.n3042 VDD.n1319 11.0319
R6414 VDD.n3042 VDD.n1313 11.0319
R6415 VDD.n3048 VDD.n1313 11.0319
R6416 VDD.n3048 VDD.n1307 11.0319
R6417 VDD.n3054 VDD.n1307 11.0319
R6418 VDD.n3054 VDD.n1301 11.0319
R6419 VDD.n3060 VDD.n1301 11.0319
R6420 VDD.n3060 VDD.n1295 11.0319
R6421 VDD.n3066 VDD.n1295 11.0319
R6422 VDD.n3072 VDD.n1288 11.0319
R6423 VDD.n3072 VDD.n1291 11.0319
R6424 VDD.n3078 VDD.n1277 11.0319
R6425 VDD.n3084 VDD.n1277 11.0319
R6426 VDD.n3084 VDD.n1271 11.0319
R6427 VDD.n3090 VDD.n1271 11.0319
R6428 VDD.n3090 VDD.n1265 11.0319
R6429 VDD.n3096 VDD.n1265 11.0319
R6430 VDD.n3096 VDD.n1259 11.0319
R6431 VDD.n3102 VDD.n1259 11.0319
R6432 VDD.n3102 VDD.n1253 11.0319
R6433 VDD.n3108 VDD.n1253 11.0319
R6434 VDD.n3108 VDD.n1247 11.0319
R6435 VDD.n3114 VDD.n1247 11.0319
R6436 VDD.n3114 VDD.n1241 11.0319
R6437 VDD.n3120 VDD.n1241 11.0319
R6438 VDD.n3120 VDD.n1235 11.0319
R6439 VDD.n3126 VDD.n1235 11.0319
R6440 VDD.n3132 VDD.n1229 11.0319
R6441 VDD.n3138 VDD.n1223 11.0319
R6442 VDD.n3138 VDD.n1217 11.0319
R6443 VDD.n3144 VDD.n1217 11.0319
R6444 VDD.n3144 VDD.n1211 11.0319
R6445 VDD.n3150 VDD.n1211 11.0319
R6446 VDD.n3150 VDD.n1205 11.0319
R6447 VDD.n3156 VDD.n1205 11.0319
R6448 VDD.n3156 VDD.n1199 11.0319
R6449 VDD.n3162 VDD.n1199 11.0319
R6450 VDD.n3162 VDD.n1193 11.0319
R6451 VDD.n3168 VDD.n1193 11.0319
R6452 VDD.n3168 VDD.n1187 11.0319
R6453 VDD.n3174 VDD.n1187 11.0319
R6454 VDD.n3174 VDD.n1181 11.0319
R6455 VDD.n3180 VDD.n1181 11.0319
R6456 VDD.n3180 VDD.n1175 11.0319
R6457 VDD.n3186 VDD.n1175 11.0319
R6458 VDD.n3192 VDD.n1169 11.0319
R6459 VDD.n3198 VDD.n1163 11.0319
R6460 VDD.n3198 VDD.n1157 11.0319
R6461 VDD.n3204 VDD.n1157 11.0319
R6462 VDD.n3204 VDD.n1151 11.0319
R6463 VDD.n3210 VDD.n1151 11.0319
R6464 VDD.n3210 VDD.n1145 11.0319
R6465 VDD.n3216 VDD.n1145 11.0319
R6466 VDD.n3216 VDD.n1139 11.0319
R6467 VDD.n3222 VDD.n1139 11.0319
R6468 VDD.n3222 VDD.n1133 11.0319
R6469 VDD.n3228 VDD.n1133 11.0319
R6470 VDD.n3228 VDD.n1127 11.0319
R6471 VDD.n3234 VDD.n1127 11.0319
R6472 VDD.n3234 VDD.n1121 11.0319
R6473 VDD.n3240 VDD.n1121 11.0319
R6474 VDD.n3240 VDD.n1114 11.0319
R6475 VDD.n3246 VDD.n1114 11.0319
R6476 VDD.n3246 VDD.n1117 11.0319
R6477 VDD.n3252 VDD.n1110 11.0319
R6478 VDD.n3258 VDD.n1097 11.0319
R6479 VDD.n3264 VDD.n1097 11.0319
R6480 VDD.n3264 VDD.n1090 11.0319
R6481 VDD.n3272 VDD.n1090 11.0319
R6482 VDD.n3272 VDD.n1084 11.0319
R6483 VDD.n3278 VDD.n1084 11.0319
R6484 VDD.n3278 VDD.n1073 11.0319
R6485 VDD.n3335 VDD.n1073 11.0319
R6486 VDD.n3335 VDD.n1067 11.0319
R6487 VDD.n3341 VDD.n1067 11.0319
R6488 VDD.n3341 VDD.n1036 11.0319
R6489 VDD.n3817 VDD.n1030 11.0319
R6490 VDD.n3823 VDD.n1030 11.0319
R6491 VDD.n3823 VDD.n1024 11.0319
R6492 VDD.n3829 VDD.n1024 11.0319
R6493 VDD.n3829 VDD.n1018 11.0319
R6494 VDD.n3835 VDD.n1018 11.0319
R6495 VDD.n3835 VDD.n1012 11.0319
R6496 VDD.n3841 VDD.n1012 11.0319
R6497 VDD.n3841 VDD.n1005 11.0319
R6498 VDD.n3847 VDD.n1005 11.0319
R6499 VDD.n3847 VDD.n1008 11.0319
R6500 VDD.n3853 VDD.n1001 11.0319
R6501 VDD.n3859 VDD.n988 11.0319
R6502 VDD.n3865 VDD.n988 11.0319
R6503 VDD.n3865 VDD.n982 11.0319
R6504 VDD.n3871 VDD.n982 11.0319
R6505 VDD.n3871 VDD.n976 11.0319
R6506 VDD.n3877 VDD.n976 11.0319
R6507 VDD.n3877 VDD.n970 11.0319
R6508 VDD.n3883 VDD.n970 11.0319
R6509 VDD.n3883 VDD.n964 11.0319
R6510 VDD.n3889 VDD.n964 11.0319
R6511 VDD.n3889 VDD.n958 11.0319
R6512 VDD.n3895 VDD.n958 11.0319
R6513 VDD.n3895 VDD.n952 11.0319
R6514 VDD.n3901 VDD.n952 11.0319
R6515 VDD.n3901 VDD.n946 11.0319
R6516 VDD.n3907 VDD.n946 11.0319
R6517 VDD.n3907 VDD.n940 11.0319
R6518 VDD.n3913 VDD.n940 11.0319
R6519 VDD.n3919 VDD.n934 11.0319
R6520 VDD.n3925 VDD.n928 11.0319
R6521 VDD.n3925 VDD.n922 11.0319
R6522 VDD.n3931 VDD.n922 11.0319
R6523 VDD.n3931 VDD.n916 11.0319
R6524 VDD.n3937 VDD.n916 11.0319
R6525 VDD.n3937 VDD.n910 11.0319
R6526 VDD.n3943 VDD.n910 11.0319
R6527 VDD.n3943 VDD.n904 11.0319
R6528 VDD.n3949 VDD.n904 11.0319
R6529 VDD.n3949 VDD.n898 11.0319
R6530 VDD.n3955 VDD.n898 11.0319
R6531 VDD.n3955 VDD.n892 11.0319
R6532 VDD.n3961 VDD.n892 11.0319
R6533 VDD.n3961 VDD.n886 11.0319
R6534 VDD.n3967 VDD.n886 11.0319
R6535 VDD.n3967 VDD.n880 11.0319
R6536 VDD.n3973 VDD.n880 11.0319
R6537 VDD.n3979 VDD.n874 11.0319
R6538 VDD.n3985 VDD.n868 11.0319
R6539 VDD.n3985 VDD.n862 11.0319
R6540 VDD.n3991 VDD.n862 11.0319
R6541 VDD.n3991 VDD.n856 11.0319
R6542 VDD.n3997 VDD.n856 11.0319
R6543 VDD.n3997 VDD.n850 11.0319
R6544 VDD.n4003 VDD.n850 11.0319
R6545 VDD.n4003 VDD.n844 11.0319
R6546 VDD.n4009 VDD.n844 11.0319
R6547 VDD.n4009 VDD.n838 11.0319
R6548 VDD.n4015 VDD.n838 11.0319
R6549 VDD.n4015 VDD.n832 11.0319
R6550 VDD.n4021 VDD.n832 11.0319
R6551 VDD.n4021 VDD.n825 11.0319
R6552 VDD.n4027 VDD.n825 11.0319
R6553 VDD.n4027 VDD.n828 11.0319
R6554 VDD.n4033 VDD.n814 11.0319
R6555 VDD.n4039 VDD.n814 11.0319
R6556 VDD.n4045 VDD.n808 11.0319
R6557 VDD.n4045 VDD.n802 11.0319
R6558 VDD.n4051 VDD.n802 11.0319
R6559 VDD.n4051 VDD.n796 11.0319
R6560 VDD.n4057 VDD.n796 11.0319
R6561 VDD.n4057 VDD.n790 11.0319
R6562 VDD.n4063 VDD.n790 11.0319
R6563 VDD.n4063 VDD.n784 11.0319
R6564 VDD.n4069 VDD.n784 11.0319
R6565 VDD.n4069 VDD.n778 11.0319
R6566 VDD.n4075 VDD.n778 11.0319
R6567 VDD.n4075 VDD.n772 11.0319
R6568 VDD.n4081 VDD.n772 11.0319
R6569 VDD.n4081 VDD.n766 11.0319
R6570 VDD.n4087 VDD.n766 11.0319
R6571 VDD.n4087 VDD.n760 11.0319
R6572 VDD.n4093 VDD.n760 11.0319
R6573 VDD.n4093 VDD.n754 11.0319
R6574 VDD.n4099 VDD.n754 11.0319
R6575 VDD.n4099 VDD.n747 11.0319
R6576 VDD.n4105 VDD.n747 11.0319
R6577 VDD.n4105 VDD.n750 11.0319
R6578 VDD.n4111 VDD.n736 11.0319
R6579 VDD.n4117 VDD.n736 11.0319
R6580 VDD.n4123 VDD.n730 11.0319
R6581 VDD.n4123 VDD.n723 11.0319
R6582 VDD.n4159 VDD.n723 11.0319
R6583 VDD.n4159 VDD.n717 11.0319
R6584 VDD.n4165 VDD.n717 11.0319
R6585 VDD.n4165 VDD.n691 11.0319
R6586 VDD.n4213 VDD.n691 11.0319
R6587 VDD.n4213 VDD.n693 11.0319
R6588 VDD.n3066 VDD.t84 10.7075
R6589 VDD.t3 VDD.n1169 10.7075
R6590 VDD.n3919 VDD.t91 10.7075
R6591 VDD.t81 VDD.n808 10.7075
R6592 VDD.n3597 VDD.n3596 10.6151
R6593 VDD.n3596 VDD.n3595 10.6151
R6594 VDD.n3595 VDD.n3594 10.6151
R6595 VDD.n3594 VDD.n3592 10.6151
R6596 VDD.n3592 VDD.n3591 10.6151
R6597 VDD.n3591 VDD.n3589 10.6151
R6598 VDD.n3589 VDD.n3588 10.6151
R6599 VDD.n3588 VDD.n3586 10.6151
R6600 VDD.n3586 VDD.n3585 10.6151
R6601 VDD.n3585 VDD.n3583 10.6151
R6602 VDD.n3583 VDD.n3582 10.6151
R6603 VDD.n3582 VDD.n3580 10.6151
R6604 VDD.n3580 VDD.n3579 10.6151
R6605 VDD.n3579 VDD.n3577 10.6151
R6606 VDD.n3577 VDD.n3576 10.6151
R6607 VDD.n3576 VDD.n3574 10.6151
R6608 VDD.n3574 VDD.n3573 10.6151
R6609 VDD.n3573 VDD.n3571 10.6151
R6610 VDD.n3571 VDD.n3570 10.6151
R6611 VDD.n3570 VDD.n3568 10.6151
R6612 VDD.n3568 VDD.n3567 10.6151
R6613 VDD.n3567 VDD.n3565 10.6151
R6614 VDD.n3565 VDD.n3564 10.6151
R6615 VDD.n3564 VDD.n3562 10.6151
R6616 VDD.n3562 VDD.n3561 10.6151
R6617 VDD.n3561 VDD.n3559 10.6151
R6618 VDD.n3559 VDD.n3558 10.6151
R6619 VDD.n3558 VDD.n3556 10.6151
R6620 VDD.n3556 VDD.n3555 10.6151
R6621 VDD.n3555 VDD.n3553 10.6151
R6622 VDD.n3553 VDD.n3552 10.6151
R6623 VDD.n3552 VDD.n3550 10.6151
R6624 VDD.n3550 VDD.n3549 10.6151
R6625 VDD.n3549 VDD.n3547 10.6151
R6626 VDD.n3547 VDD.n3546 10.6151
R6627 VDD.n3546 VDD.n3544 10.6151
R6628 VDD.n3544 VDD.n3543 10.6151
R6629 VDD.n3543 VDD.n3541 10.6151
R6630 VDD.n3541 VDD.n3540 10.6151
R6631 VDD.n3540 VDD.n3538 10.6151
R6632 VDD.n3538 VDD.n3537 10.6151
R6633 VDD.n3537 VDD.n3535 10.6151
R6634 VDD.n3535 VDD.n3534 10.6151
R6635 VDD.n3534 VDD.n3532 10.6151
R6636 VDD.n3532 VDD.n3531 10.6151
R6637 VDD.n3531 VDD.n3529 10.6151
R6638 VDD.n3529 VDD.n3528 10.6151
R6639 VDD.n3528 VDD.n3526 10.6151
R6640 VDD.n3526 VDD.n3525 10.6151
R6641 VDD.n3525 VDD.n3523 10.6151
R6642 VDD.n3523 VDD.n3522 10.6151
R6643 VDD.n3522 VDD.n3520 10.6151
R6644 VDD.n3520 VDD.n3519 10.6151
R6645 VDD.n3519 VDD.n3517 10.6151
R6646 VDD.n3517 VDD.n3516 10.6151
R6647 VDD.n3516 VDD.n3514 10.6151
R6648 VDD.n3514 VDD.n3513 10.6151
R6649 VDD.n3513 VDD.n3511 10.6151
R6650 VDD.n3511 VDD.n3510 10.6151
R6651 VDD.n3510 VDD.n3508 10.6151
R6652 VDD.n3508 VDD.n3507 10.6151
R6653 VDD.n3507 VDD.n3505 10.6151
R6654 VDD.n3505 VDD.n3504 10.6151
R6655 VDD.n3504 VDD.n3502 10.6151
R6656 VDD.n3502 VDD.n3501 10.6151
R6657 VDD.n3501 VDD.n3499 10.6151
R6658 VDD.n3499 VDD.n3498 10.6151
R6659 VDD.n3498 VDD.n3496 10.6151
R6660 VDD.n3496 VDD.n3495 10.6151
R6661 VDD.n3495 VDD.n3493 10.6151
R6662 VDD.n3493 VDD.n3492 10.6151
R6663 VDD.n3492 VDD.n3490 10.6151
R6664 VDD.n3490 VDD.n3489 10.6151
R6665 VDD.n3489 VDD.n3487 10.6151
R6666 VDD.n3487 VDD.n3486 10.6151
R6667 VDD.n3486 VDD.n3484 10.6151
R6668 VDD.n3484 VDD.n3483 10.6151
R6669 VDD.n3483 VDD.n3481 10.6151
R6670 VDD.n3481 VDD.n3480 10.6151
R6671 VDD.n3480 VDD.n3478 10.6151
R6672 VDD.n3478 VDD.n3477 10.6151
R6673 VDD.n3477 VDD.n3475 10.6151
R6674 VDD.n3475 VDD.n3474 10.6151
R6675 VDD.n3474 VDD.n3472 10.6151
R6676 VDD.n3472 VDD.n3471 10.6151
R6677 VDD.n3471 VDD.n3469 10.6151
R6678 VDD.n3469 VDD.n3468 10.6151
R6679 VDD.n3468 VDD.n3466 10.6151
R6680 VDD.n3466 VDD.n3465 10.6151
R6681 VDD.n3465 VDD.n3463 10.6151
R6682 VDD.n3463 VDD.n3462 10.6151
R6683 VDD.n3462 VDD.n3460 10.6151
R6684 VDD.n3460 VDD.n3459 10.6151
R6685 VDD.n3459 VDD.n3457 10.6151
R6686 VDD.n3457 VDD.n3456 10.6151
R6687 VDD.n3456 VDD.n3454 10.6151
R6688 VDD.n3454 VDD.n3453 10.6151
R6689 VDD.n3453 VDD.n3451 10.6151
R6690 VDD.n3451 VDD.n3450 10.6151
R6691 VDD.n3450 VDD.n3448 10.6151
R6692 VDD.n3448 VDD.n3447 10.6151
R6693 VDD.n3447 VDD.n3445 10.6151
R6694 VDD.n3445 VDD.n3444 10.6151
R6695 VDD.n3444 VDD.n3442 10.6151
R6696 VDD.n3442 VDD.n3441 10.6151
R6697 VDD.n3441 VDD.n715 10.6151
R6698 VDD.n4168 VDD.n715 10.6151
R6699 VDD.n4169 VDD.n4168 10.6151
R6700 VDD.n4170 VDD.n4169 10.6151
R6701 VDD.n3400 VDD.n1034 10.6151
R6702 VDD.n3400 VDD.n3399 10.6151
R6703 VDD.n3406 VDD.n3399 10.6151
R6704 VDD.n3407 VDD.n3406 10.6151
R6705 VDD.n3408 VDD.n3407 10.6151
R6706 VDD.n3408 VDD.n3397 10.6151
R6707 VDD.n3414 VDD.n3397 10.6151
R6708 VDD.n3415 VDD.n3414 10.6151
R6709 VDD.n3416 VDD.n3415 10.6151
R6710 VDD.n3416 VDD.n3395 10.6151
R6711 VDD.n3422 VDD.n3395 10.6151
R6712 VDD.n3423 VDD.n3422 10.6151
R6713 VDD.n3424 VDD.n3423 10.6151
R6714 VDD.n3424 VDD.n3393 10.6151
R6715 VDD.n3430 VDD.n3393 10.6151
R6716 VDD.n3431 VDD.n3430 10.6151
R6717 VDD.n3433 VDD.n3389 10.6151
R6718 VDD.n3439 VDD.n3389 10.6151
R6719 VDD.n3440 VDD.n3439 10.6151
R6720 VDD.n3820 VDD.n3819 10.6151
R6721 VDD.n3821 VDD.n3820 10.6151
R6722 VDD.n3821 VDD.n1022 10.6151
R6723 VDD.n3831 VDD.n1022 10.6151
R6724 VDD.n3832 VDD.n3831 10.6151
R6725 VDD.n3833 VDD.n3832 10.6151
R6726 VDD.n3833 VDD.n1010 10.6151
R6727 VDD.n3843 VDD.n1010 10.6151
R6728 VDD.n3844 VDD.n3843 10.6151
R6729 VDD.n3845 VDD.n3844 10.6151
R6730 VDD.n3845 VDD.n997 10.6151
R6731 VDD.n3855 VDD.n997 10.6151
R6732 VDD.n3856 VDD.n3855 10.6151
R6733 VDD.n3857 VDD.n3856 10.6151
R6734 VDD.n3857 VDD.n986 10.6151
R6735 VDD.n3867 VDD.n986 10.6151
R6736 VDD.n3868 VDD.n3867 10.6151
R6737 VDD.n3869 VDD.n3868 10.6151
R6738 VDD.n3869 VDD.n974 10.6151
R6739 VDD.n3879 VDD.n974 10.6151
R6740 VDD.n3880 VDD.n3879 10.6151
R6741 VDD.n3881 VDD.n3880 10.6151
R6742 VDD.n3881 VDD.n962 10.6151
R6743 VDD.n3891 VDD.n962 10.6151
R6744 VDD.n3892 VDD.n3891 10.6151
R6745 VDD.n3893 VDD.n3892 10.6151
R6746 VDD.n3893 VDD.n950 10.6151
R6747 VDD.n3903 VDD.n950 10.6151
R6748 VDD.n3904 VDD.n3903 10.6151
R6749 VDD.n3905 VDD.n3904 10.6151
R6750 VDD.n3905 VDD.n938 10.6151
R6751 VDD.n3915 VDD.n938 10.6151
R6752 VDD.n3916 VDD.n3915 10.6151
R6753 VDD.n3917 VDD.n3916 10.6151
R6754 VDD.n3917 VDD.n926 10.6151
R6755 VDD.n3927 VDD.n926 10.6151
R6756 VDD.n3928 VDD.n3927 10.6151
R6757 VDD.n3929 VDD.n3928 10.6151
R6758 VDD.n3929 VDD.n914 10.6151
R6759 VDD.n3939 VDD.n914 10.6151
R6760 VDD.n3940 VDD.n3939 10.6151
R6761 VDD.n3941 VDD.n3940 10.6151
R6762 VDD.n3941 VDD.n902 10.6151
R6763 VDD.n3951 VDD.n902 10.6151
R6764 VDD.n3952 VDD.n3951 10.6151
R6765 VDD.n3953 VDD.n3952 10.6151
R6766 VDD.n3953 VDD.n890 10.6151
R6767 VDD.n3963 VDD.n890 10.6151
R6768 VDD.n3964 VDD.n3963 10.6151
R6769 VDD.n3965 VDD.n3964 10.6151
R6770 VDD.n3965 VDD.n878 10.6151
R6771 VDD.n3975 VDD.n878 10.6151
R6772 VDD.n3976 VDD.n3975 10.6151
R6773 VDD.n3977 VDD.n3976 10.6151
R6774 VDD.n3977 VDD.n866 10.6151
R6775 VDD.n3987 VDD.n866 10.6151
R6776 VDD.n3988 VDD.n3987 10.6151
R6777 VDD.n3989 VDD.n3988 10.6151
R6778 VDD.n3989 VDD.n854 10.6151
R6779 VDD.n3999 VDD.n854 10.6151
R6780 VDD.n4000 VDD.n3999 10.6151
R6781 VDD.n4001 VDD.n4000 10.6151
R6782 VDD.n4001 VDD.n842 10.6151
R6783 VDD.n4011 VDD.n842 10.6151
R6784 VDD.n4012 VDD.n4011 10.6151
R6785 VDD.n4013 VDD.n4012 10.6151
R6786 VDD.n4013 VDD.n830 10.6151
R6787 VDD.n4023 VDD.n830 10.6151
R6788 VDD.n4024 VDD.n4023 10.6151
R6789 VDD.n4025 VDD.n4024 10.6151
R6790 VDD.n4025 VDD.n818 10.6151
R6791 VDD.n4035 VDD.n818 10.6151
R6792 VDD.n4036 VDD.n4035 10.6151
R6793 VDD.n4037 VDD.n4036 10.6151
R6794 VDD.n4037 VDD.n806 10.6151
R6795 VDD.n4047 VDD.n806 10.6151
R6796 VDD.n4048 VDD.n4047 10.6151
R6797 VDD.n4049 VDD.n4048 10.6151
R6798 VDD.n4049 VDD.n794 10.6151
R6799 VDD.n4059 VDD.n794 10.6151
R6800 VDD.n4060 VDD.n4059 10.6151
R6801 VDD.n4061 VDD.n4060 10.6151
R6802 VDD.n4061 VDD.n782 10.6151
R6803 VDD.n4071 VDD.n782 10.6151
R6804 VDD.n4072 VDD.n4071 10.6151
R6805 VDD.n4073 VDD.n4072 10.6151
R6806 VDD.n4073 VDD.n770 10.6151
R6807 VDD.n4083 VDD.n770 10.6151
R6808 VDD.n4084 VDD.n4083 10.6151
R6809 VDD.n4085 VDD.n4084 10.6151
R6810 VDD.n4085 VDD.n758 10.6151
R6811 VDD.n4095 VDD.n758 10.6151
R6812 VDD.n4096 VDD.n4095 10.6151
R6813 VDD.n4097 VDD.n4096 10.6151
R6814 VDD.n4097 VDD.n745 10.6151
R6815 VDD.n4107 VDD.n745 10.6151
R6816 VDD.n4108 VDD.n4107 10.6151
R6817 VDD.n4109 VDD.n4108 10.6151
R6818 VDD.n4109 VDD.n734 10.6151
R6819 VDD.n4119 VDD.n734 10.6151
R6820 VDD.n4120 VDD.n4119 10.6151
R6821 VDD.n4121 VDD.n4120 10.6151
R6822 VDD.n4121 VDD.n721 10.6151
R6823 VDD.n4161 VDD.n721 10.6151
R6824 VDD.n4162 VDD.n4161 10.6151
R6825 VDD.n4163 VDD.n4162 10.6151
R6826 VDD.n4163 VDD.n697 10.6151
R6827 VDD.n4211 VDD.n697 10.6151
R6828 VDD.n4211 VDD.n4210 10.6151
R6829 VDD.n4209 VDD.n698 10.6151
R6830 VDD.n4204 VDD.n698 10.6151
R6831 VDD.n4204 VDD.n4203 10.6151
R6832 VDD.n4203 VDD.n4202 10.6151
R6833 VDD.n4202 VDD.n700 10.6151
R6834 VDD.n4197 VDD.n700 10.6151
R6835 VDD.n4197 VDD.n4196 10.6151
R6836 VDD.n4196 VDD.n4195 10.6151
R6837 VDD.n4195 VDD.n703 10.6151
R6838 VDD.n4190 VDD.n703 10.6151
R6839 VDD.n4190 VDD.n4189 10.6151
R6840 VDD.n4189 VDD.n4188 10.6151
R6841 VDD.n4188 VDD.n706 10.6151
R6842 VDD.n4183 VDD.n706 10.6151
R6843 VDD.n4183 VDD.n4182 10.6151
R6844 VDD.n4182 VDD.n4181 10.6151
R6845 VDD.n4176 VDD.n713 10.6151
R6846 VDD.n4176 VDD.n4175 10.6151
R6847 VDD.n4175 VDD.n4174 10.6151
R6848 VDD.n4128 VDD.n4127 10.6151
R6849 VDD.n4145 VDD.n4128 10.6151
R6850 VDD.n4145 VDD.n4144 10.6151
R6851 VDD.n4144 VDD.n4143 10.6151
R6852 VDD.n4143 VDD.n4130 10.6151
R6853 VDD.n4138 VDD.n4130 10.6151
R6854 VDD.n4138 VDD.n4137 10.6151
R6855 VDD.n4137 VDD.n4136 10.6151
R6856 VDD.n4136 VDD.n676 10.6151
R6857 VDD.n4237 VDD.n676 10.6151
R6858 VDD.n4237 VDD.n677 10.6151
R6859 VDD.n4232 VDD.n677 10.6151
R6860 VDD.n4232 VDD.n4231 10.6151
R6861 VDD.n4231 VDD.n4230 10.6151
R6862 VDD.n4230 VDD.n681 10.6151
R6863 VDD.n4225 VDD.n681 10.6151
R6864 VDD.n4223 VDD.n4222 10.6151
R6865 VDD.n4222 VDD.n686 10.6151
R6866 VDD.n4217 VDD.n686 10.6151
R6867 VDD.n3772 VDD.n3771 10.6151
R6868 VDD.n3771 VDD.n3769 10.6151
R6869 VDD.n3769 VDD.n3768 10.6151
R6870 VDD.n3768 VDD.n3766 10.6151
R6871 VDD.n3766 VDD.n3765 10.6151
R6872 VDD.n3765 VDD.n3763 10.6151
R6873 VDD.n3763 VDD.n3762 10.6151
R6874 VDD.n3762 VDD.n3760 10.6151
R6875 VDD.n3760 VDD.n3759 10.6151
R6876 VDD.n3759 VDD.n3757 10.6151
R6877 VDD.n3757 VDD.n3756 10.6151
R6878 VDD.n3756 VDD.n3754 10.6151
R6879 VDD.n3754 VDD.n3753 10.6151
R6880 VDD.n3753 VDD.n3751 10.6151
R6881 VDD.n3751 VDD.n3750 10.6151
R6882 VDD.n3750 VDD.n3748 10.6151
R6883 VDD.n3748 VDD.n3747 10.6151
R6884 VDD.n3747 VDD.n3745 10.6151
R6885 VDD.n3745 VDD.n3744 10.6151
R6886 VDD.n3744 VDD.n3742 10.6151
R6887 VDD.n3742 VDD.n3741 10.6151
R6888 VDD.n3741 VDD.n3739 10.6151
R6889 VDD.n3739 VDD.n3738 10.6151
R6890 VDD.n3738 VDD.n3736 10.6151
R6891 VDD.n3736 VDD.n3735 10.6151
R6892 VDD.n3735 VDD.n3733 10.6151
R6893 VDD.n3733 VDD.n3732 10.6151
R6894 VDD.n3732 VDD.n3730 10.6151
R6895 VDD.n3730 VDD.n3729 10.6151
R6896 VDD.n3729 VDD.n3727 10.6151
R6897 VDD.n3727 VDD.n3726 10.6151
R6898 VDD.n3726 VDD.n3724 10.6151
R6899 VDD.n3724 VDD.n3723 10.6151
R6900 VDD.n3723 VDD.n3721 10.6151
R6901 VDD.n3721 VDD.n3720 10.6151
R6902 VDD.n3720 VDD.n3718 10.6151
R6903 VDD.n3718 VDD.n3717 10.6151
R6904 VDD.n3717 VDD.n3715 10.6151
R6905 VDD.n3715 VDD.n3714 10.6151
R6906 VDD.n3714 VDD.n3712 10.6151
R6907 VDD.n3712 VDD.n3711 10.6151
R6908 VDD.n3711 VDD.n3709 10.6151
R6909 VDD.n3709 VDD.n3708 10.6151
R6910 VDD.n3708 VDD.n3706 10.6151
R6911 VDD.n3706 VDD.n3705 10.6151
R6912 VDD.n3705 VDD.n3703 10.6151
R6913 VDD.n3703 VDD.n3702 10.6151
R6914 VDD.n3702 VDD.n3700 10.6151
R6915 VDD.n3700 VDD.n3699 10.6151
R6916 VDD.n3699 VDD.n3697 10.6151
R6917 VDD.n3697 VDD.n3696 10.6151
R6918 VDD.n3696 VDD.n3694 10.6151
R6919 VDD.n3694 VDD.n3693 10.6151
R6920 VDD.n3693 VDD.n3691 10.6151
R6921 VDD.n3691 VDD.n3690 10.6151
R6922 VDD.n3690 VDD.n3688 10.6151
R6923 VDD.n3688 VDD.n3687 10.6151
R6924 VDD.n3687 VDD.n3685 10.6151
R6925 VDD.n3685 VDD.n3684 10.6151
R6926 VDD.n3684 VDD.n3682 10.6151
R6927 VDD.n3682 VDD.n3681 10.6151
R6928 VDD.n3681 VDD.n3679 10.6151
R6929 VDD.n3679 VDD.n3678 10.6151
R6930 VDD.n3678 VDD.n3676 10.6151
R6931 VDD.n3676 VDD.n3675 10.6151
R6932 VDD.n3675 VDD.n3673 10.6151
R6933 VDD.n3673 VDD.n3672 10.6151
R6934 VDD.n3672 VDD.n3670 10.6151
R6935 VDD.n3670 VDD.n3669 10.6151
R6936 VDD.n3669 VDD.n3667 10.6151
R6937 VDD.n3667 VDD.n3666 10.6151
R6938 VDD.n3666 VDD.n3664 10.6151
R6939 VDD.n3664 VDD.n3663 10.6151
R6940 VDD.n3663 VDD.n3661 10.6151
R6941 VDD.n3661 VDD.n3660 10.6151
R6942 VDD.n3660 VDD.n3658 10.6151
R6943 VDD.n3658 VDD.n3657 10.6151
R6944 VDD.n3657 VDD.n3655 10.6151
R6945 VDD.n3655 VDD.n3654 10.6151
R6946 VDD.n3654 VDD.n3652 10.6151
R6947 VDD.n3652 VDD.n3651 10.6151
R6948 VDD.n3651 VDD.n3649 10.6151
R6949 VDD.n3649 VDD.n3648 10.6151
R6950 VDD.n3648 VDD.n3646 10.6151
R6951 VDD.n3646 VDD.n3645 10.6151
R6952 VDD.n3645 VDD.n3643 10.6151
R6953 VDD.n3643 VDD.n3642 10.6151
R6954 VDD.n3642 VDD.n3640 10.6151
R6955 VDD.n3640 VDD.n3639 10.6151
R6956 VDD.n3639 VDD.n3637 10.6151
R6957 VDD.n3637 VDD.n3636 10.6151
R6958 VDD.n3636 VDD.n3634 10.6151
R6959 VDD.n3634 VDD.n3633 10.6151
R6960 VDD.n3633 VDD.n3631 10.6151
R6961 VDD.n3631 VDD.n3630 10.6151
R6962 VDD.n3630 VDD.n3628 10.6151
R6963 VDD.n3628 VDD.n3627 10.6151
R6964 VDD.n3627 VDD.n3625 10.6151
R6965 VDD.n3625 VDD.n3624 10.6151
R6966 VDD.n3624 VDD.n3622 10.6151
R6967 VDD.n3622 VDD.n3621 10.6151
R6968 VDD.n3621 VDD.n3619 10.6151
R6969 VDD.n3619 VDD.n3618 10.6151
R6970 VDD.n3618 VDD.n3616 10.6151
R6971 VDD.n3616 VDD.n3615 10.6151
R6972 VDD.n3615 VDD.n3613 10.6151
R6973 VDD.n3613 VDD.n689 10.6151
R6974 VDD.n4215 VDD.n689 10.6151
R6975 VDD.n4216 VDD.n4215 10.6151
R6976 VDD.n3814 VDD.n3813 10.6151
R6977 VDD.n3813 VDD.n3601 10.6151
R6978 VDD.n3807 VDD.n3601 10.6151
R6979 VDD.n3807 VDD.n3806 10.6151
R6980 VDD.n3806 VDD.n3805 10.6151
R6981 VDD.n3805 VDD.n3603 10.6151
R6982 VDD.n3799 VDD.n3603 10.6151
R6983 VDD.n3799 VDD.n3798 10.6151
R6984 VDD.n3798 VDD.n3797 10.6151
R6985 VDD.n3797 VDD.n3605 10.6151
R6986 VDD.n3791 VDD.n3605 10.6151
R6987 VDD.n3791 VDD.n3790 10.6151
R6988 VDD.n3790 VDD.n3789 10.6151
R6989 VDD.n3789 VDD.n3607 10.6151
R6990 VDD.n3783 VDD.n3607 10.6151
R6991 VDD.n3783 VDD.n3782 10.6151
R6992 VDD.n3780 VDD.n3611 10.6151
R6993 VDD.n3774 VDD.n3611 10.6151
R6994 VDD.n3774 VDD.n3773 10.6151
R6995 VDD.n3815 VDD.n1028 10.6151
R6996 VDD.n3825 VDD.n1028 10.6151
R6997 VDD.n3826 VDD.n3825 10.6151
R6998 VDD.n3827 VDD.n3826 10.6151
R6999 VDD.n3827 VDD.n1016 10.6151
R7000 VDD.n3837 VDD.n1016 10.6151
R7001 VDD.n3838 VDD.n3837 10.6151
R7002 VDD.n3839 VDD.n3838 10.6151
R7003 VDD.n3839 VDD.n1003 10.6151
R7004 VDD.n3849 VDD.n1003 10.6151
R7005 VDD.n3850 VDD.n3849 10.6151
R7006 VDD.n3851 VDD.n3850 10.6151
R7007 VDD.n3851 VDD.n992 10.6151
R7008 VDD.n3861 VDD.n992 10.6151
R7009 VDD.n3862 VDD.n3861 10.6151
R7010 VDD.n3863 VDD.n3862 10.6151
R7011 VDD.n3863 VDD.n980 10.6151
R7012 VDD.n3873 VDD.n980 10.6151
R7013 VDD.n3874 VDD.n3873 10.6151
R7014 VDD.n3875 VDD.n3874 10.6151
R7015 VDD.n3875 VDD.n968 10.6151
R7016 VDD.n3885 VDD.n968 10.6151
R7017 VDD.n3886 VDD.n3885 10.6151
R7018 VDD.n3887 VDD.n3886 10.6151
R7019 VDD.n3887 VDD.n956 10.6151
R7020 VDD.n3897 VDD.n956 10.6151
R7021 VDD.n3898 VDD.n3897 10.6151
R7022 VDD.n3899 VDD.n3898 10.6151
R7023 VDD.n3899 VDD.n944 10.6151
R7024 VDD.n3909 VDD.n944 10.6151
R7025 VDD.n3910 VDD.n3909 10.6151
R7026 VDD.n3911 VDD.n3910 10.6151
R7027 VDD.n3911 VDD.n932 10.6151
R7028 VDD.n3921 VDD.n932 10.6151
R7029 VDD.n3922 VDD.n3921 10.6151
R7030 VDD.n3923 VDD.n3922 10.6151
R7031 VDD.n3923 VDD.n920 10.6151
R7032 VDD.n3933 VDD.n920 10.6151
R7033 VDD.n3934 VDD.n3933 10.6151
R7034 VDD.n3935 VDD.n3934 10.6151
R7035 VDD.n3935 VDD.n908 10.6151
R7036 VDD.n3945 VDD.n908 10.6151
R7037 VDD.n3946 VDD.n3945 10.6151
R7038 VDD.n3947 VDD.n3946 10.6151
R7039 VDD.n3947 VDD.n896 10.6151
R7040 VDD.n3957 VDD.n896 10.6151
R7041 VDD.n3958 VDD.n3957 10.6151
R7042 VDD.n3959 VDD.n3958 10.6151
R7043 VDD.n3959 VDD.n884 10.6151
R7044 VDD.n3969 VDD.n884 10.6151
R7045 VDD.n3970 VDD.n3969 10.6151
R7046 VDD.n3971 VDD.n3970 10.6151
R7047 VDD.n3971 VDD.n872 10.6151
R7048 VDD.n3981 VDD.n872 10.6151
R7049 VDD.n3982 VDD.n3981 10.6151
R7050 VDD.n3983 VDD.n3982 10.6151
R7051 VDD.n3983 VDD.n860 10.6151
R7052 VDD.n3993 VDD.n860 10.6151
R7053 VDD.n3994 VDD.n3993 10.6151
R7054 VDD.n3995 VDD.n3994 10.6151
R7055 VDD.n3995 VDD.n848 10.6151
R7056 VDD.n4005 VDD.n848 10.6151
R7057 VDD.n4006 VDD.n4005 10.6151
R7058 VDD.n4007 VDD.n4006 10.6151
R7059 VDD.n4007 VDD.n836 10.6151
R7060 VDD.n4017 VDD.n836 10.6151
R7061 VDD.n4018 VDD.n4017 10.6151
R7062 VDD.n4019 VDD.n4018 10.6151
R7063 VDD.n4019 VDD.n823 10.6151
R7064 VDD.n4029 VDD.n823 10.6151
R7065 VDD.n4030 VDD.n4029 10.6151
R7066 VDD.n4031 VDD.n4030 10.6151
R7067 VDD.n4031 VDD.n812 10.6151
R7068 VDD.n4041 VDD.n812 10.6151
R7069 VDD.n4042 VDD.n4041 10.6151
R7070 VDD.n4043 VDD.n4042 10.6151
R7071 VDD.n4043 VDD.n800 10.6151
R7072 VDD.n4053 VDD.n800 10.6151
R7073 VDD.n4054 VDD.n4053 10.6151
R7074 VDD.n4055 VDD.n4054 10.6151
R7075 VDD.n4055 VDD.n788 10.6151
R7076 VDD.n4065 VDD.n788 10.6151
R7077 VDD.n4066 VDD.n4065 10.6151
R7078 VDD.n4067 VDD.n4066 10.6151
R7079 VDD.n4067 VDD.n776 10.6151
R7080 VDD.n4077 VDD.n776 10.6151
R7081 VDD.n4078 VDD.n4077 10.6151
R7082 VDD.n4079 VDD.n4078 10.6151
R7083 VDD.n4079 VDD.n764 10.6151
R7084 VDD.n4089 VDD.n764 10.6151
R7085 VDD.n4090 VDD.n4089 10.6151
R7086 VDD.n4091 VDD.n4090 10.6151
R7087 VDD.n4091 VDD.n752 10.6151
R7088 VDD.n4101 VDD.n752 10.6151
R7089 VDD.n4102 VDD.n4101 10.6151
R7090 VDD.n4103 VDD.n4102 10.6151
R7091 VDD.n4103 VDD.n740 10.6151
R7092 VDD.n4113 VDD.n740 10.6151
R7093 VDD.n4114 VDD.n4113 10.6151
R7094 VDD.n4115 VDD.n4114 10.6151
R7095 VDD.n4115 VDD.n728 10.6151
R7096 VDD.n4125 VDD.n728 10.6151
R7097 VDD.n4126 VDD.n4125 10.6151
R7098 VDD.n4157 VDD.n4126 10.6151
R7099 VDD.n4157 VDD.n4156 10.6151
R7100 VDD.n4156 VDD.n4155 10.6151
R7101 VDD.n4155 VDD.n4154 10.6151
R7102 VDD.n4154 VDD.n4152 10.6151
R7103 VDD.n4152 VDD.n4151 10.6151
R7104 VDD.n2962 VDD.n1389 10.6151
R7105 VDD.n2972 VDD.n1389 10.6151
R7106 VDD.n2973 VDD.n2972 10.6151
R7107 VDD.n2974 VDD.n2973 10.6151
R7108 VDD.n2974 VDD.n1377 10.6151
R7109 VDD.n2984 VDD.n1377 10.6151
R7110 VDD.n2985 VDD.n2984 10.6151
R7111 VDD.n2986 VDD.n2985 10.6151
R7112 VDD.n2986 VDD.n1364 10.6151
R7113 VDD.n2996 VDD.n1364 10.6151
R7114 VDD.n2997 VDD.n2996 10.6151
R7115 VDD.n2998 VDD.n2997 10.6151
R7116 VDD.n2998 VDD.n1353 10.6151
R7117 VDD.n3008 VDD.n1353 10.6151
R7118 VDD.n3009 VDD.n3008 10.6151
R7119 VDD.n3010 VDD.n3009 10.6151
R7120 VDD.n3010 VDD.n1341 10.6151
R7121 VDD.n3020 VDD.n1341 10.6151
R7122 VDD.n3021 VDD.n3020 10.6151
R7123 VDD.n3022 VDD.n3021 10.6151
R7124 VDD.n3022 VDD.n1329 10.6151
R7125 VDD.n3032 VDD.n1329 10.6151
R7126 VDD.n3033 VDD.n3032 10.6151
R7127 VDD.n3034 VDD.n3033 10.6151
R7128 VDD.n3034 VDD.n1317 10.6151
R7129 VDD.n3044 VDD.n1317 10.6151
R7130 VDD.n3045 VDD.n3044 10.6151
R7131 VDD.n3046 VDD.n3045 10.6151
R7132 VDD.n3046 VDD.n1305 10.6151
R7133 VDD.n3056 VDD.n1305 10.6151
R7134 VDD.n3057 VDD.n3056 10.6151
R7135 VDD.n3058 VDD.n3057 10.6151
R7136 VDD.n3058 VDD.n1293 10.6151
R7137 VDD.n3068 VDD.n1293 10.6151
R7138 VDD.n3069 VDD.n3068 10.6151
R7139 VDD.n3070 VDD.n3069 10.6151
R7140 VDD.n3070 VDD.n1281 10.6151
R7141 VDD.n3080 VDD.n1281 10.6151
R7142 VDD.n3081 VDD.n3080 10.6151
R7143 VDD.n3082 VDD.n3081 10.6151
R7144 VDD.n3082 VDD.n1269 10.6151
R7145 VDD.n3092 VDD.n1269 10.6151
R7146 VDD.n3093 VDD.n3092 10.6151
R7147 VDD.n3094 VDD.n3093 10.6151
R7148 VDD.n3094 VDD.n1257 10.6151
R7149 VDD.n3104 VDD.n1257 10.6151
R7150 VDD.n3105 VDD.n3104 10.6151
R7151 VDD.n3106 VDD.n3105 10.6151
R7152 VDD.n3106 VDD.n1245 10.6151
R7153 VDD.n3116 VDD.n1245 10.6151
R7154 VDD.n3117 VDD.n3116 10.6151
R7155 VDD.n3118 VDD.n3117 10.6151
R7156 VDD.n3118 VDD.n1233 10.6151
R7157 VDD.n3128 VDD.n1233 10.6151
R7158 VDD.n3129 VDD.n3128 10.6151
R7159 VDD.n3130 VDD.n3129 10.6151
R7160 VDD.n3130 VDD.n1221 10.6151
R7161 VDD.n3140 VDD.n1221 10.6151
R7162 VDD.n3141 VDD.n3140 10.6151
R7163 VDD.n3142 VDD.n3141 10.6151
R7164 VDD.n3142 VDD.n1209 10.6151
R7165 VDD.n3152 VDD.n1209 10.6151
R7166 VDD.n3153 VDD.n3152 10.6151
R7167 VDD.n3154 VDD.n3153 10.6151
R7168 VDD.n3154 VDD.n1197 10.6151
R7169 VDD.n3164 VDD.n1197 10.6151
R7170 VDD.n3165 VDD.n3164 10.6151
R7171 VDD.n3166 VDD.n3165 10.6151
R7172 VDD.n3166 VDD.n1185 10.6151
R7173 VDD.n3176 VDD.n1185 10.6151
R7174 VDD.n3177 VDD.n3176 10.6151
R7175 VDD.n3178 VDD.n3177 10.6151
R7176 VDD.n3178 VDD.n1173 10.6151
R7177 VDD.n3188 VDD.n1173 10.6151
R7178 VDD.n3189 VDD.n3188 10.6151
R7179 VDD.n3190 VDD.n3189 10.6151
R7180 VDD.n3190 VDD.n1161 10.6151
R7181 VDD.n3200 VDD.n1161 10.6151
R7182 VDD.n3201 VDD.n3200 10.6151
R7183 VDD.n3202 VDD.n3201 10.6151
R7184 VDD.n3202 VDD.n1149 10.6151
R7185 VDD.n3212 VDD.n1149 10.6151
R7186 VDD.n3213 VDD.n3212 10.6151
R7187 VDD.n3214 VDD.n3213 10.6151
R7188 VDD.n3214 VDD.n1137 10.6151
R7189 VDD.n3224 VDD.n1137 10.6151
R7190 VDD.n3225 VDD.n3224 10.6151
R7191 VDD.n3226 VDD.n3225 10.6151
R7192 VDD.n3226 VDD.n1125 10.6151
R7193 VDD.n3236 VDD.n1125 10.6151
R7194 VDD.n3237 VDD.n3236 10.6151
R7195 VDD.n3238 VDD.n3237 10.6151
R7196 VDD.n3238 VDD.n1112 10.6151
R7197 VDD.n3248 VDD.n1112 10.6151
R7198 VDD.n3249 VDD.n3248 10.6151
R7199 VDD.n3250 VDD.n3249 10.6151
R7200 VDD.n3250 VDD.n1101 10.6151
R7201 VDD.n3260 VDD.n1101 10.6151
R7202 VDD.n3261 VDD.n3260 10.6151
R7203 VDD.n3262 VDD.n3261 10.6151
R7204 VDD.n3262 VDD.n1088 10.6151
R7205 VDD.n3274 VDD.n1088 10.6151
R7206 VDD.n3275 VDD.n3274 10.6151
R7207 VDD.n3276 VDD.n3275 10.6151
R7208 VDD.n3276 VDD.n1071 10.6151
R7209 VDD.n3337 VDD.n1071 10.6151
R7210 VDD.n3338 VDD.n3337 10.6151
R7211 VDD.n3339 VDD.n3338 10.6151
R7212 VDD.n3339 VDD.n1060 10.6151
R7213 VDD.n3383 VDD.n3382 10.6151
R7214 VDD.n3382 VDD.n3381 10.6151
R7215 VDD.n3381 VDD.n3378 10.6151
R7216 VDD.n3378 VDD.n3377 10.6151
R7217 VDD.n3377 VDD.n3374 10.6151
R7218 VDD.n3374 VDD.n3373 10.6151
R7219 VDD.n3373 VDD.n3370 10.6151
R7220 VDD.n3370 VDD.n3369 10.6151
R7221 VDD.n3369 VDD.n3366 10.6151
R7222 VDD.n3366 VDD.n3365 10.6151
R7223 VDD.n3365 VDD.n3362 10.6151
R7224 VDD.n3362 VDD.n3361 10.6151
R7225 VDD.n3361 VDD.n3358 10.6151
R7226 VDD.n3358 VDD.n3357 10.6151
R7227 VDD.n3357 VDD.n3354 10.6151
R7228 VDD.n3354 VDD.n3353 10.6151
R7229 VDD.n3350 VDD.n3349 10.6151
R7230 VDD.n3349 VDD.n3346 10.6151
R7231 VDD.n3346 VDD.n3345 10.6151
R7232 VDD.n1574 VDD.n1573 10.6151
R7233 VDD.n1573 VDD.n1571 10.6151
R7234 VDD.n1571 VDD.n1570 10.6151
R7235 VDD.n1570 VDD.n1568 10.6151
R7236 VDD.n1568 VDD.n1567 10.6151
R7237 VDD.n1567 VDD.n1565 10.6151
R7238 VDD.n1565 VDD.n1564 10.6151
R7239 VDD.n1564 VDD.n1562 10.6151
R7240 VDD.n1562 VDD.n1561 10.6151
R7241 VDD.n1561 VDD.n1559 10.6151
R7242 VDD.n1559 VDD.n1558 10.6151
R7243 VDD.n1558 VDD.n1556 10.6151
R7244 VDD.n1556 VDD.n1555 10.6151
R7245 VDD.n1555 VDD.n1553 10.6151
R7246 VDD.n1553 VDD.n1552 10.6151
R7247 VDD.n1552 VDD.n1550 10.6151
R7248 VDD.n1550 VDD.n1549 10.6151
R7249 VDD.n1549 VDD.n1547 10.6151
R7250 VDD.n1547 VDD.n1546 10.6151
R7251 VDD.n1546 VDD.n1544 10.6151
R7252 VDD.n1544 VDD.n1543 10.6151
R7253 VDD.n1543 VDD.n1541 10.6151
R7254 VDD.n1541 VDD.n1540 10.6151
R7255 VDD.n1540 VDD.n1538 10.6151
R7256 VDD.n1538 VDD.n1537 10.6151
R7257 VDD.n1537 VDD.n1535 10.6151
R7258 VDD.n1535 VDD.n1534 10.6151
R7259 VDD.n1534 VDD.n1532 10.6151
R7260 VDD.n1532 VDD.n1531 10.6151
R7261 VDD.n1531 VDD.n1529 10.6151
R7262 VDD.n1529 VDD.n1528 10.6151
R7263 VDD.n1528 VDD.n1526 10.6151
R7264 VDD.n1526 VDD.n1525 10.6151
R7265 VDD.n1525 VDD.n1523 10.6151
R7266 VDD.n1523 VDD.n1522 10.6151
R7267 VDD.n1522 VDD.n1520 10.6151
R7268 VDD.n1520 VDD.n1519 10.6151
R7269 VDD.n1519 VDD.n1517 10.6151
R7270 VDD.n1517 VDD.n1516 10.6151
R7271 VDD.n1516 VDD.n1514 10.6151
R7272 VDD.n1514 VDD.n1513 10.6151
R7273 VDD.n1513 VDD.n1511 10.6151
R7274 VDD.n1511 VDD.n1510 10.6151
R7275 VDD.n1510 VDD.n1508 10.6151
R7276 VDD.n1508 VDD.n1507 10.6151
R7277 VDD.n1507 VDD.n1505 10.6151
R7278 VDD.n1505 VDD.n1504 10.6151
R7279 VDD.n1504 VDD.n1502 10.6151
R7280 VDD.n1502 VDD.n1501 10.6151
R7281 VDD.n1501 VDD.n1499 10.6151
R7282 VDD.n1499 VDD.n1498 10.6151
R7283 VDD.n1498 VDD.n1496 10.6151
R7284 VDD.n1496 VDD.n1495 10.6151
R7285 VDD.n1495 VDD.n1493 10.6151
R7286 VDD.n1493 VDD.n1492 10.6151
R7287 VDD.n1492 VDD.n1490 10.6151
R7288 VDD.n1490 VDD.n1489 10.6151
R7289 VDD.n1489 VDD.n1487 10.6151
R7290 VDD.n1487 VDD.n1486 10.6151
R7291 VDD.n1486 VDD.n1484 10.6151
R7292 VDD.n1484 VDD.n1483 10.6151
R7293 VDD.n1483 VDD.n1481 10.6151
R7294 VDD.n1481 VDD.n1480 10.6151
R7295 VDD.n1480 VDD.n1478 10.6151
R7296 VDD.n1478 VDD.n1477 10.6151
R7297 VDD.n1477 VDD.n1475 10.6151
R7298 VDD.n1475 VDD.n1474 10.6151
R7299 VDD.n1474 VDD.n1472 10.6151
R7300 VDD.n1472 VDD.n1471 10.6151
R7301 VDD.n1471 VDD.n1469 10.6151
R7302 VDD.n1469 VDD.n1468 10.6151
R7303 VDD.n1468 VDD.n1466 10.6151
R7304 VDD.n1466 VDD.n1465 10.6151
R7305 VDD.n1465 VDD.n1463 10.6151
R7306 VDD.n1463 VDD.n1462 10.6151
R7307 VDD.n1462 VDD.n1460 10.6151
R7308 VDD.n1460 VDD.n1459 10.6151
R7309 VDD.n1459 VDD.n1457 10.6151
R7310 VDD.n1457 VDD.n1456 10.6151
R7311 VDD.n1456 VDD.n1454 10.6151
R7312 VDD.n1454 VDD.n1453 10.6151
R7313 VDD.n1453 VDD.n1451 10.6151
R7314 VDD.n1451 VDD.n1450 10.6151
R7315 VDD.n1450 VDD.n1448 10.6151
R7316 VDD.n1448 VDD.n1447 10.6151
R7317 VDD.n1447 VDD.n1445 10.6151
R7318 VDD.n1445 VDD.n1444 10.6151
R7319 VDD.n1444 VDD.n1442 10.6151
R7320 VDD.n1442 VDD.n1441 10.6151
R7321 VDD.n1441 VDD.n1439 10.6151
R7322 VDD.n1439 VDD.n1438 10.6151
R7323 VDD.n1438 VDD.n1436 10.6151
R7324 VDD.n1436 VDD.n1435 10.6151
R7325 VDD.n1435 VDD.n1433 10.6151
R7326 VDD.n1433 VDD.n1432 10.6151
R7327 VDD.n1432 VDD.n1430 10.6151
R7328 VDD.n1430 VDD.n1429 10.6151
R7329 VDD.n1429 VDD.n1427 10.6151
R7330 VDD.n1427 VDD.n1426 10.6151
R7331 VDD.n1426 VDD.n1424 10.6151
R7332 VDD.n1424 VDD.n1423 10.6151
R7333 VDD.n1423 VDD.n1421 10.6151
R7334 VDD.n1421 VDD.n1420 10.6151
R7335 VDD.n1420 VDD.n1418 10.6151
R7336 VDD.n1418 VDD.n1417 10.6151
R7337 VDD.n1417 VDD.n1415 10.6151
R7338 VDD.n1415 VDD.n1414 10.6151
R7339 VDD.n1414 VDD.n1066 10.6151
R7340 VDD.n1066 VDD.n1064 10.6151
R7341 VDD.n2961 VDD.n2960 10.6151
R7342 VDD.n2960 VDD.n1401 10.6151
R7343 VDD.n2955 VDD.n1401 10.6151
R7344 VDD.n2955 VDD.n2954 10.6151
R7345 VDD.n2954 VDD.n1403 10.6151
R7346 VDD.n2949 VDD.n1403 10.6151
R7347 VDD.n2949 VDD.n2948 10.6151
R7348 VDD.n2948 VDD.n2947 10.6151
R7349 VDD.n2947 VDD.n1405 10.6151
R7350 VDD.n2941 VDD.n1405 10.6151
R7351 VDD.n2941 VDD.n1594 10.6151
R7352 VDD.n1594 VDD.n1593 10.6151
R7353 VDD.n1593 VDD.n1407 10.6151
R7354 VDD.n1587 VDD.n1407 10.6151
R7355 VDD.n1587 VDD.n1586 10.6151
R7356 VDD.n1586 VDD.n1585 10.6151
R7357 VDD.n1581 VDD.n1580 10.6151
R7358 VDD.n1580 VDD.n1413 10.6151
R7359 VDD.n1575 VDD.n1413 10.6151
R7360 VDD.n3328 VDD.n3327 10.6151
R7361 VDD.n3327 VDD.n3325 10.6151
R7362 VDD.n3325 VDD.n3322 10.6151
R7363 VDD.n3322 VDD.n3321 10.6151
R7364 VDD.n3321 VDD.n3318 10.6151
R7365 VDD.n3318 VDD.n3317 10.6151
R7366 VDD.n3317 VDD.n3314 10.6151
R7367 VDD.n3314 VDD.n3313 10.6151
R7368 VDD.n3313 VDD.n3310 10.6151
R7369 VDD.n3310 VDD.n3309 10.6151
R7370 VDD.n3309 VDD.n3306 10.6151
R7371 VDD.n3306 VDD.n3305 10.6151
R7372 VDD.n3305 VDD.n3302 10.6151
R7373 VDD.n3302 VDD.n3301 10.6151
R7374 VDD.n3301 VDD.n3298 10.6151
R7375 VDD.n3298 VDD.n3297 10.6151
R7376 VDD.n3294 VDD.n3293 10.6151
R7377 VDD.n3293 VDD.n3290 10.6151
R7378 VDD.n3290 VDD.n3289 10.6151
R7379 VDD.n1781 VDD.n1780 10.6151
R7380 VDD.n1780 VDD.n1778 10.6151
R7381 VDD.n1778 VDD.n1777 10.6151
R7382 VDD.n1777 VDD.n1775 10.6151
R7383 VDD.n1775 VDD.n1774 10.6151
R7384 VDD.n1774 VDD.n1772 10.6151
R7385 VDD.n1772 VDD.n1771 10.6151
R7386 VDD.n1771 VDD.n1769 10.6151
R7387 VDD.n1769 VDD.n1768 10.6151
R7388 VDD.n1768 VDD.n1766 10.6151
R7389 VDD.n1766 VDD.n1765 10.6151
R7390 VDD.n1765 VDD.n1763 10.6151
R7391 VDD.n1763 VDD.n1762 10.6151
R7392 VDD.n1762 VDD.n1760 10.6151
R7393 VDD.n1760 VDD.n1759 10.6151
R7394 VDD.n1759 VDD.n1757 10.6151
R7395 VDD.n1757 VDD.n1756 10.6151
R7396 VDD.n1756 VDD.n1754 10.6151
R7397 VDD.n1754 VDD.n1753 10.6151
R7398 VDD.n1753 VDD.n1751 10.6151
R7399 VDD.n1751 VDD.n1750 10.6151
R7400 VDD.n1750 VDD.n1748 10.6151
R7401 VDD.n1748 VDD.n1747 10.6151
R7402 VDD.n1747 VDD.n1745 10.6151
R7403 VDD.n1745 VDD.n1744 10.6151
R7404 VDD.n1744 VDD.n1742 10.6151
R7405 VDD.n1742 VDD.n1741 10.6151
R7406 VDD.n1741 VDD.n1739 10.6151
R7407 VDD.n1739 VDD.n1738 10.6151
R7408 VDD.n1738 VDD.n1736 10.6151
R7409 VDD.n1736 VDD.n1735 10.6151
R7410 VDD.n1735 VDD.n1733 10.6151
R7411 VDD.n1733 VDD.n1732 10.6151
R7412 VDD.n1732 VDD.n1730 10.6151
R7413 VDD.n1730 VDD.n1729 10.6151
R7414 VDD.n1729 VDD.n1727 10.6151
R7415 VDD.n1727 VDD.n1726 10.6151
R7416 VDD.n1726 VDD.n1724 10.6151
R7417 VDD.n1724 VDD.n1723 10.6151
R7418 VDD.n1723 VDD.n1721 10.6151
R7419 VDD.n1721 VDD.n1720 10.6151
R7420 VDD.n1720 VDD.n1718 10.6151
R7421 VDD.n1718 VDD.n1717 10.6151
R7422 VDD.n1717 VDD.n1715 10.6151
R7423 VDD.n1715 VDD.n1714 10.6151
R7424 VDD.n1714 VDD.n1712 10.6151
R7425 VDD.n1712 VDD.n1711 10.6151
R7426 VDD.n1711 VDD.n1709 10.6151
R7427 VDD.n1709 VDD.n1708 10.6151
R7428 VDD.n1708 VDD.n1706 10.6151
R7429 VDD.n1706 VDD.n1705 10.6151
R7430 VDD.n1705 VDD.n1703 10.6151
R7431 VDD.n1703 VDD.n1702 10.6151
R7432 VDD.n1702 VDD.n1700 10.6151
R7433 VDD.n1700 VDD.n1699 10.6151
R7434 VDD.n1699 VDD.n1697 10.6151
R7435 VDD.n1697 VDD.n1696 10.6151
R7436 VDD.n1696 VDD.n1694 10.6151
R7437 VDD.n1694 VDD.n1693 10.6151
R7438 VDD.n1693 VDD.n1691 10.6151
R7439 VDD.n1691 VDD.n1690 10.6151
R7440 VDD.n1690 VDD.n1688 10.6151
R7441 VDD.n1688 VDD.n1687 10.6151
R7442 VDD.n1687 VDD.n1685 10.6151
R7443 VDD.n1685 VDD.n1684 10.6151
R7444 VDD.n1684 VDD.n1682 10.6151
R7445 VDD.n1682 VDD.n1681 10.6151
R7446 VDD.n1681 VDD.n1679 10.6151
R7447 VDD.n1679 VDD.n1678 10.6151
R7448 VDD.n1678 VDD.n1676 10.6151
R7449 VDD.n1676 VDD.n1675 10.6151
R7450 VDD.n1675 VDD.n1673 10.6151
R7451 VDD.n1673 VDD.n1672 10.6151
R7452 VDD.n1672 VDD.n1670 10.6151
R7453 VDD.n1670 VDD.n1669 10.6151
R7454 VDD.n1669 VDD.n1667 10.6151
R7455 VDD.n1667 VDD.n1666 10.6151
R7456 VDD.n1666 VDD.n1664 10.6151
R7457 VDD.n1664 VDD.n1663 10.6151
R7458 VDD.n1663 VDD.n1661 10.6151
R7459 VDD.n1661 VDD.n1660 10.6151
R7460 VDD.n1660 VDD.n1658 10.6151
R7461 VDD.n1658 VDD.n1657 10.6151
R7462 VDD.n1657 VDD.n1655 10.6151
R7463 VDD.n1655 VDD.n1654 10.6151
R7464 VDD.n1654 VDD.n1652 10.6151
R7465 VDD.n1652 VDD.n1651 10.6151
R7466 VDD.n1651 VDD.n1649 10.6151
R7467 VDD.n1649 VDD.n1648 10.6151
R7468 VDD.n1648 VDD.n1646 10.6151
R7469 VDD.n1646 VDD.n1645 10.6151
R7470 VDD.n1645 VDD.n1643 10.6151
R7471 VDD.n1643 VDD.n1642 10.6151
R7472 VDD.n1642 VDD.n1640 10.6151
R7473 VDD.n1640 VDD.n1639 10.6151
R7474 VDD.n1639 VDD.n1637 10.6151
R7475 VDD.n1637 VDD.n1636 10.6151
R7476 VDD.n1636 VDD.n1634 10.6151
R7477 VDD.n1634 VDD.n1633 10.6151
R7478 VDD.n1633 VDD.n1631 10.6151
R7479 VDD.n1631 VDD.n1630 10.6151
R7480 VDD.n1630 VDD.n1628 10.6151
R7481 VDD.n1628 VDD.n1627 10.6151
R7482 VDD.n1627 VDD.n1082 10.6151
R7483 VDD.n3281 VDD.n1082 10.6151
R7484 VDD.n3282 VDD.n3281 10.6151
R7485 VDD.n3284 VDD.n3282 10.6151
R7486 VDD.n3285 VDD.n3284 10.6151
R7487 VDD.n3286 VDD.n3285 10.6151
R7488 VDD.n1601 VDD.n1395 10.6151
R7489 VDD.n1606 VDD.n1601 10.6151
R7490 VDD.n1607 VDD.n1606 10.6151
R7491 VDD.n1608 VDD.n1607 10.6151
R7492 VDD.n1608 VDD.n1599 10.6151
R7493 VDD.n1614 VDD.n1599 10.6151
R7494 VDD.n1615 VDD.n1614 10.6151
R7495 VDD.n1616 VDD.n1615 10.6151
R7496 VDD.n1616 VDD.n1596 10.6151
R7497 VDD.n1803 VDD.n1596 10.6151
R7498 VDD.n1803 VDD.n1597 10.6151
R7499 VDD.n1798 VDD.n1597 10.6151
R7500 VDD.n1798 VDD.n1797 10.6151
R7501 VDD.n1797 VDD.n1621 10.6151
R7502 VDD.n1792 VDD.n1621 10.6151
R7503 VDD.n1792 VDD.n1791 10.6151
R7504 VDD.n1789 VDD.n1625 10.6151
R7505 VDD.n1783 VDD.n1625 10.6151
R7506 VDD.n1783 VDD.n1782 10.6151
R7507 VDD.n2967 VDD.n2966 10.6151
R7508 VDD.n2968 VDD.n2967 10.6151
R7509 VDD.n2968 VDD.n1383 10.6151
R7510 VDD.n2978 VDD.n1383 10.6151
R7511 VDD.n2979 VDD.n2978 10.6151
R7512 VDD.n2980 VDD.n2979 10.6151
R7513 VDD.n2980 VDD.n1371 10.6151
R7514 VDD.n2990 VDD.n1371 10.6151
R7515 VDD.n2991 VDD.n2990 10.6151
R7516 VDD.n2992 VDD.n2991 10.6151
R7517 VDD.n2992 VDD.n1359 10.6151
R7518 VDD.n3002 VDD.n1359 10.6151
R7519 VDD.n3003 VDD.n3002 10.6151
R7520 VDD.n3004 VDD.n3003 10.6151
R7521 VDD.n3004 VDD.n1347 10.6151
R7522 VDD.n3014 VDD.n1347 10.6151
R7523 VDD.n3015 VDD.n3014 10.6151
R7524 VDD.n3016 VDD.n3015 10.6151
R7525 VDD.n3016 VDD.n1335 10.6151
R7526 VDD.n3026 VDD.n1335 10.6151
R7527 VDD.n3027 VDD.n3026 10.6151
R7528 VDD.n3028 VDD.n3027 10.6151
R7529 VDD.n3028 VDD.n1323 10.6151
R7530 VDD.n3038 VDD.n1323 10.6151
R7531 VDD.n3039 VDD.n3038 10.6151
R7532 VDD.n3040 VDD.n3039 10.6151
R7533 VDD.n3040 VDD.n1311 10.6151
R7534 VDD.n3050 VDD.n1311 10.6151
R7535 VDD.n3051 VDD.n3050 10.6151
R7536 VDD.n3052 VDD.n3051 10.6151
R7537 VDD.n3052 VDD.n1299 10.6151
R7538 VDD.n3062 VDD.n1299 10.6151
R7539 VDD.n3063 VDD.n3062 10.6151
R7540 VDD.n3064 VDD.n3063 10.6151
R7541 VDD.n3064 VDD.n1286 10.6151
R7542 VDD.n3074 VDD.n1286 10.6151
R7543 VDD.n3075 VDD.n3074 10.6151
R7544 VDD.n3076 VDD.n3075 10.6151
R7545 VDD.n3076 VDD.n1275 10.6151
R7546 VDD.n3086 VDD.n1275 10.6151
R7547 VDD.n3087 VDD.n3086 10.6151
R7548 VDD.n3088 VDD.n3087 10.6151
R7549 VDD.n3088 VDD.n1263 10.6151
R7550 VDD.n3098 VDD.n1263 10.6151
R7551 VDD.n3099 VDD.n3098 10.6151
R7552 VDD.n3100 VDD.n3099 10.6151
R7553 VDD.n3100 VDD.n1251 10.6151
R7554 VDD.n3110 VDD.n1251 10.6151
R7555 VDD.n3111 VDD.n3110 10.6151
R7556 VDD.n3112 VDD.n3111 10.6151
R7557 VDD.n3112 VDD.n1239 10.6151
R7558 VDD.n3122 VDD.n1239 10.6151
R7559 VDD.n3123 VDD.n3122 10.6151
R7560 VDD.n3124 VDD.n3123 10.6151
R7561 VDD.n3124 VDD.n1227 10.6151
R7562 VDD.n3134 VDD.n1227 10.6151
R7563 VDD.n3135 VDD.n3134 10.6151
R7564 VDD.n3136 VDD.n3135 10.6151
R7565 VDD.n3136 VDD.n1215 10.6151
R7566 VDD.n3146 VDD.n1215 10.6151
R7567 VDD.n3147 VDD.n3146 10.6151
R7568 VDD.n3148 VDD.n3147 10.6151
R7569 VDD.n3148 VDD.n1203 10.6151
R7570 VDD.n3158 VDD.n1203 10.6151
R7571 VDD.n3159 VDD.n3158 10.6151
R7572 VDD.n3160 VDD.n3159 10.6151
R7573 VDD.n3160 VDD.n1191 10.6151
R7574 VDD.n3170 VDD.n1191 10.6151
R7575 VDD.n3171 VDD.n3170 10.6151
R7576 VDD.n3172 VDD.n3171 10.6151
R7577 VDD.n3172 VDD.n1179 10.6151
R7578 VDD.n3182 VDD.n1179 10.6151
R7579 VDD.n3183 VDD.n3182 10.6151
R7580 VDD.n3184 VDD.n3183 10.6151
R7581 VDD.n3184 VDD.n1167 10.6151
R7582 VDD.n3194 VDD.n1167 10.6151
R7583 VDD.n3195 VDD.n3194 10.6151
R7584 VDD.n3196 VDD.n3195 10.6151
R7585 VDD.n3196 VDD.n1155 10.6151
R7586 VDD.n3206 VDD.n1155 10.6151
R7587 VDD.n3207 VDD.n3206 10.6151
R7588 VDD.n3208 VDD.n3207 10.6151
R7589 VDD.n3208 VDD.n1143 10.6151
R7590 VDD.n3218 VDD.n1143 10.6151
R7591 VDD.n3219 VDD.n3218 10.6151
R7592 VDD.n3220 VDD.n3219 10.6151
R7593 VDD.n3220 VDD.n1131 10.6151
R7594 VDD.n3230 VDD.n1131 10.6151
R7595 VDD.n3231 VDD.n3230 10.6151
R7596 VDD.n3232 VDD.n3231 10.6151
R7597 VDD.n3232 VDD.n1119 10.6151
R7598 VDD.n3242 VDD.n1119 10.6151
R7599 VDD.n3243 VDD.n3242 10.6151
R7600 VDD.n3244 VDD.n3243 10.6151
R7601 VDD.n3244 VDD.n1106 10.6151
R7602 VDD.n3254 VDD.n1106 10.6151
R7603 VDD.n3255 VDD.n3254 10.6151
R7604 VDD.n3256 VDD.n3255 10.6151
R7605 VDD.n3256 VDD.n1095 10.6151
R7606 VDD.n3266 VDD.n1095 10.6151
R7607 VDD.n3267 VDD.n3266 10.6151
R7608 VDD.n3270 VDD.n3267 10.6151
R7609 VDD.n3270 VDD.n3269 10.6151
R7610 VDD.n3269 VDD.n3268 10.6151
R7611 VDD.n3268 VDD.n1078 10.6151
R7612 VDD.n3333 VDD.n1078 10.6151
R7613 VDD.n3333 VDD.n3332 10.6151
R7614 VDD.n3332 VDD.n3331 10.6151
R7615 VDD.n3331 VDD.n3330 10.6151
R7616 VDD.n2453 VDD.t120 9.73411
R7617 VDD.t112 VDD.n1915 9.73411
R7618 VDD.n4332 VDD.t118 9.73411
R7619 VDD.n4635 VDD.t104 9.73411
R7620 VDD.n4255 VDD.n4254 9.3005
R7621 VDD.n4256 VDD.n534 9.3005
R7622 VDD.n4258 VDD.n4257 9.3005
R7623 VDD.n523 VDD.n522 9.3005
R7624 VDD.n4271 VDD.n4270 9.3005
R7625 VDD.n4272 VDD.n521 9.3005
R7626 VDD.n4274 VDD.n4273 9.3005
R7627 VDD.n512 VDD.n511 9.3005
R7628 VDD.n4287 VDD.n4286 9.3005
R7629 VDD.n4288 VDD.n510 9.3005
R7630 VDD.n4290 VDD.n4289 9.3005
R7631 VDD.n500 VDD.n499 9.3005
R7632 VDD.n4303 VDD.n4302 9.3005
R7633 VDD.n4304 VDD.n498 9.3005
R7634 VDD.n4306 VDD.n4305 9.3005
R7635 VDD.n488 VDD.n487 9.3005
R7636 VDD.n4319 VDD.n4318 9.3005
R7637 VDD.n4320 VDD.n486 9.3005
R7638 VDD.n4322 VDD.n4321 9.3005
R7639 VDD.n476 VDD.n475 9.3005
R7640 VDD.n4335 VDD.n4334 9.3005
R7641 VDD.n4336 VDD.n474 9.3005
R7642 VDD.n4338 VDD.n4337 9.3005
R7643 VDD.n464 VDD.n463 9.3005
R7644 VDD.n4351 VDD.n4350 9.3005
R7645 VDD.n4352 VDD.n462 9.3005
R7646 VDD.n4354 VDD.n4353 9.3005
R7647 VDD.n452 VDD.n451 9.3005
R7648 VDD.n4367 VDD.n4366 9.3005
R7649 VDD.n4368 VDD.n450 9.3005
R7650 VDD.n4370 VDD.n4369 9.3005
R7651 VDD.n440 VDD.n439 9.3005
R7652 VDD.n4383 VDD.n4382 9.3005
R7653 VDD.n4384 VDD.n438 9.3005
R7654 VDD.n4386 VDD.n4385 9.3005
R7655 VDD.n428 VDD.n427 9.3005
R7656 VDD.n4399 VDD.n4398 9.3005
R7657 VDD.n4400 VDD.n426 9.3005
R7658 VDD.n4402 VDD.n4401 9.3005
R7659 VDD.n416 VDD.n415 9.3005
R7660 VDD.n4415 VDD.n4414 9.3005
R7661 VDD.n4416 VDD.n414 9.3005
R7662 VDD.n4418 VDD.n4417 9.3005
R7663 VDD.n403 VDD.n402 9.3005
R7664 VDD.n4431 VDD.n4430 9.3005
R7665 VDD.n4432 VDD.n401 9.3005
R7666 VDD.n4434 VDD.n4433 9.3005
R7667 VDD.n392 VDD.n391 9.3005
R7668 VDD.n4447 VDD.n4446 9.3005
R7669 VDD.n4448 VDD.n390 9.3005
R7670 VDD.n4452 VDD.n4449 9.3005
R7671 VDD.n4451 VDD.n4450 9.3005
R7672 VDD.n380 VDD.n379 9.3005
R7673 VDD.n4466 VDD.n4465 9.3005
R7674 VDD.n4467 VDD.n378 9.3005
R7675 VDD.n4472 VDD.n4468 9.3005
R7676 VDD.n4471 VDD.n4470 9.3005
R7677 VDD.n4469 VDD.n367 9.3005
R7678 VDD.n4487 VDD.n368 9.3005
R7679 VDD.n4488 VDD.n366 9.3005
R7680 VDD.n4490 VDD.n4489 9.3005
R7681 VDD.n4491 VDD.n365 9.3005
R7682 VDD.n4494 VDD.n4492 9.3005
R7683 VDD.n4495 VDD.n364 9.3005
R7684 VDD.n4497 VDD.n4496 9.3005
R7685 VDD.n4498 VDD.n363 9.3005
R7686 VDD.n4501 VDD.n4499 9.3005
R7687 VDD.n4502 VDD.n362 9.3005
R7688 VDD.n4504 VDD.n4503 9.3005
R7689 VDD.n4505 VDD.n361 9.3005
R7690 VDD.n4508 VDD.n4506 9.3005
R7691 VDD.n4509 VDD.n360 9.3005
R7692 VDD.n4511 VDD.n4510 9.3005
R7693 VDD.n4512 VDD.n359 9.3005
R7694 VDD.n4515 VDD.n4513 9.3005
R7695 VDD.n4516 VDD.n358 9.3005
R7696 VDD.n4518 VDD.n4517 9.3005
R7697 VDD.n4519 VDD.n357 9.3005
R7698 VDD.n4522 VDD.n4520 9.3005
R7699 VDD.n4523 VDD.n356 9.3005
R7700 VDD.n4525 VDD.n4524 9.3005
R7701 VDD.n4526 VDD.n355 9.3005
R7702 VDD.n4529 VDD.n4527 9.3005
R7703 VDD.n4530 VDD.n354 9.3005
R7704 VDD.n4532 VDD.n4531 9.3005
R7705 VDD.n4533 VDD.n353 9.3005
R7706 VDD.n4536 VDD.n4534 9.3005
R7707 VDD.n4537 VDD.n352 9.3005
R7708 VDD.n4539 VDD.n4538 9.3005
R7709 VDD.n4540 VDD.n351 9.3005
R7710 VDD.n4543 VDD.n4541 9.3005
R7711 VDD.n4544 VDD.n350 9.3005
R7712 VDD.n4546 VDD.n4545 9.3005
R7713 VDD.n4547 VDD.n349 9.3005
R7714 VDD.n4550 VDD.n4548 9.3005
R7715 VDD.n4551 VDD.n348 9.3005
R7716 VDD.n4553 VDD.n4552 9.3005
R7717 VDD.n4554 VDD.n347 9.3005
R7718 VDD.n4557 VDD.n4555 9.3005
R7719 VDD.n4558 VDD.n346 9.3005
R7720 VDD.n4560 VDD.n4559 9.3005
R7721 VDD.n4561 VDD.n345 9.3005
R7722 VDD.n4564 VDD.n4562 9.3005
R7723 VDD.n4565 VDD.n344 9.3005
R7724 VDD.n4567 VDD.n4566 9.3005
R7725 VDD.n4568 VDD.n343 9.3005
R7726 VDD.n4571 VDD.n4569 9.3005
R7727 VDD.n4572 VDD.n342 9.3005
R7728 VDD.n4574 VDD.n4573 9.3005
R7729 VDD.n4575 VDD.n341 9.3005
R7730 VDD.n4578 VDD.n4576 9.3005
R7731 VDD.n4579 VDD.n340 9.3005
R7732 VDD.n4581 VDD.n4580 9.3005
R7733 VDD.n4582 VDD.n339 9.3005
R7734 VDD.n4585 VDD.n4583 9.3005
R7735 VDD.n4586 VDD.n338 9.3005
R7736 VDD.n4588 VDD.n4587 9.3005
R7737 VDD.n536 VDD.n535 9.3005
R7738 VDD.n248 VDD.n243 9.3005
R7739 VDD.n252 VDD.n249 9.3005
R7740 VDD.n253 VDD.n242 9.3005
R7741 VDD.n257 VDD.n256 9.3005
R7742 VDD.n258 VDD.n241 9.3005
R7743 VDD.n262 VDD.n259 9.3005
R7744 VDD.n263 VDD.n240 9.3005
R7745 VDD.n267 VDD.n266 9.3005
R7746 VDD.n268 VDD.n239 9.3005
R7747 VDD.n272 VDD.n269 9.3005
R7748 VDD.n274 VDD.n236 9.3005
R7749 VDD.n278 VDD.n277 9.3005
R7750 VDD.n279 VDD.n235 9.3005
R7751 VDD.n283 VDD.n280 9.3005
R7752 VDD.n284 VDD.n234 9.3005
R7753 VDD.n288 VDD.n287 9.3005
R7754 VDD.n289 VDD.n233 9.3005
R7755 VDD.n293 VDD.n290 9.3005
R7756 VDD.n294 VDD.n232 9.3005
R7757 VDD.n298 VDD.n297 9.3005
R7758 VDD.n299 VDD.n231 9.3005
R7759 VDD.n303 VDD.n300 9.3005
R7760 VDD.n304 VDD.n227 9.3005
R7761 VDD.n308 VDD.n307 9.3005
R7762 VDD.n309 VDD.n226 9.3005
R7763 VDD.n313 VDD.n310 9.3005
R7764 VDD.n314 VDD.n225 9.3005
R7765 VDD.n318 VDD.n317 9.3005
R7766 VDD.n319 VDD.n224 9.3005
R7767 VDD.n323 VDD.n320 9.3005
R7768 VDD.n324 VDD.n223 9.3005
R7769 VDD.n328 VDD.n327 9.3005
R7770 VDD.n329 VDD.n222 9.3005
R7771 VDD.n333 VDD.n330 9.3005
R7772 VDD.n335 VDD.n221 9.3005
R7773 VDD.n337 VDD.n336 9.3005
R7774 VDD.n4590 VDD.n4589 9.3005
R7775 VDD.n247 VDD.n246 9.3005
R7776 VDD.n4711 VDD.n4710 9.3005
R7777 VDD.n4709 VDD.n37 9.3005
R7778 VDD.n48 VDD.n40 9.3005
R7779 VDD.n4703 VDD.n49 9.3005
R7780 VDD.n4702 VDD.n50 9.3005
R7781 VDD.n4701 VDD.n51 9.3005
R7782 VDD.n59 VDD.n52 9.3005
R7783 VDD.n4695 VDD.n60 9.3005
R7784 VDD.n4694 VDD.n61 9.3005
R7785 VDD.n4693 VDD.n62 9.3005
R7786 VDD.n69 VDD.n63 9.3005
R7787 VDD.n4687 VDD.n70 9.3005
R7788 VDD.n4686 VDD.n71 9.3005
R7789 VDD.n4685 VDD.n72 9.3005
R7790 VDD.n81 VDD.n73 9.3005
R7791 VDD.n4679 VDD.n82 9.3005
R7792 VDD.n4678 VDD.n83 9.3005
R7793 VDD.n4677 VDD.n84 9.3005
R7794 VDD.n92 VDD.n85 9.3005
R7795 VDD.n4671 VDD.n93 9.3005
R7796 VDD.n4670 VDD.n94 9.3005
R7797 VDD.n4669 VDD.n95 9.3005
R7798 VDD.n103 VDD.n96 9.3005
R7799 VDD.n4663 VDD.n104 9.3005
R7800 VDD.n4662 VDD.n105 9.3005
R7801 VDD.n4661 VDD.n106 9.3005
R7802 VDD.n114 VDD.n107 9.3005
R7803 VDD.n4655 VDD.n115 9.3005
R7804 VDD.n4654 VDD.n116 9.3005
R7805 VDD.n4653 VDD.n117 9.3005
R7806 VDD.n125 VDD.n118 9.3005
R7807 VDD.n4647 VDD.n126 9.3005
R7808 VDD.n4646 VDD.n127 9.3005
R7809 VDD.n4645 VDD.n128 9.3005
R7810 VDD.n136 VDD.n129 9.3005
R7811 VDD.n4639 VDD.n137 9.3005
R7812 VDD.n4638 VDD.n138 9.3005
R7813 VDD.n4637 VDD.n139 9.3005
R7814 VDD.n147 VDD.n140 9.3005
R7815 VDD.n4631 VDD.n148 9.3005
R7816 VDD.n4630 VDD.n149 9.3005
R7817 VDD.n4629 VDD.n150 9.3005
R7818 VDD.n158 VDD.n151 9.3005
R7819 VDD.n4623 VDD.n159 9.3005
R7820 VDD.n4622 VDD.n160 9.3005
R7821 VDD.n4621 VDD.n161 9.3005
R7822 VDD.n169 VDD.n162 9.3005
R7823 VDD.n4615 VDD.n170 9.3005
R7824 VDD.n4614 VDD.n171 9.3005
R7825 VDD.n4613 VDD.n172 9.3005
R7826 VDD.n179 VDD.n173 9.3005
R7827 VDD.n4607 VDD.n180 9.3005
R7828 VDD.n4606 VDD.n181 9.3005
R7829 VDD.n4605 VDD.n182 9.3005
R7830 VDD.n191 VDD.n183 9.3005
R7831 VDD.n4599 VDD.n192 9.3005
R7832 VDD.n4598 VDD.n193 9.3005
R7833 VDD.n4597 VDD.n194 9.3005
R7834 VDD.n244 VDD.n195 9.3005
R7835 VDD.n4250 VDD.n4249 9.3005
R7836 VDD.n530 VDD.n529 9.3005
R7837 VDD.n4263 VDD.n4262 9.3005
R7838 VDD.n4264 VDD.n528 9.3005
R7839 VDD.n4266 VDD.n4265 9.3005
R7840 VDD.n518 VDD.n517 9.3005
R7841 VDD.n4279 VDD.n4278 9.3005
R7842 VDD.n4280 VDD.n516 9.3005
R7843 VDD.n4282 VDD.n4281 9.3005
R7844 VDD.n506 VDD.n505 9.3005
R7845 VDD.n4295 VDD.n4294 9.3005
R7846 VDD.n4296 VDD.n504 9.3005
R7847 VDD.n4298 VDD.n4297 9.3005
R7848 VDD.n494 VDD.n493 9.3005
R7849 VDD.n4311 VDD.n4310 9.3005
R7850 VDD.n4312 VDD.n492 9.3005
R7851 VDD.n4314 VDD.n4313 9.3005
R7852 VDD.n482 VDD.n481 9.3005
R7853 VDD.n4327 VDD.n4326 9.3005
R7854 VDD.n4328 VDD.n480 9.3005
R7855 VDD.n4330 VDD.n4329 9.3005
R7856 VDD.n470 VDD.n469 9.3005
R7857 VDD.n4343 VDD.n4342 9.3005
R7858 VDD.n4344 VDD.n468 9.3005
R7859 VDD.n4346 VDD.n4345 9.3005
R7860 VDD.n458 VDD.n457 9.3005
R7861 VDD.n4359 VDD.n4358 9.3005
R7862 VDD.n4360 VDD.n456 9.3005
R7863 VDD.n4362 VDD.n4361 9.3005
R7864 VDD.n446 VDD.n445 9.3005
R7865 VDD.n4375 VDD.n4374 9.3005
R7866 VDD.n4376 VDD.n444 9.3005
R7867 VDD.n4378 VDD.n4377 9.3005
R7868 VDD.n434 VDD.n433 9.3005
R7869 VDD.n4391 VDD.n4390 9.3005
R7870 VDD.n4392 VDD.n432 9.3005
R7871 VDD.n4394 VDD.n4393 9.3005
R7872 VDD.n422 VDD.n421 9.3005
R7873 VDD.n4407 VDD.n4406 9.3005
R7874 VDD.n4408 VDD.n420 9.3005
R7875 VDD.n4410 VDD.n4409 9.3005
R7876 VDD.n410 VDD.n409 9.3005
R7877 VDD.n4423 VDD.n4422 9.3005
R7878 VDD.n4424 VDD.n408 9.3005
R7879 VDD.n4426 VDD.n4425 9.3005
R7880 VDD.n398 VDD.n397 9.3005
R7881 VDD.n4439 VDD.n4438 9.3005
R7882 VDD.n4440 VDD.n396 9.3005
R7883 VDD.n4442 VDD.n4441 9.3005
R7884 VDD.n386 VDD.n385 9.3005
R7885 VDD.n4457 VDD.n4456 9.3005
R7886 VDD.n4458 VDD.n384 9.3005
R7887 VDD.n4460 VDD.n4459 9.3005
R7888 VDD.n374 VDD.n373 9.3005
R7889 VDD.n4478 VDD.n4477 9.3005
R7890 VDD.n4479 VDD.n372 9.3005
R7891 VDD.n4481 VDD.n4480 9.3005
R7892 VDD.n38 VDD.n36 9.3005
R7893 VDD.n4248 VDD.n540 9.3005
R7894 VDD.n4247 VDD.n4246 9.3005
R7895 VDD.n673 VDD.n568 9.3005
R7896 VDD.n670 VDD.n669 9.3005
R7897 VDD.n668 VDD.n569 9.3005
R7898 VDD.n667 VDD.n666 9.3005
R7899 VDD.n663 VDD.n570 9.3005
R7900 VDD.n660 VDD.n659 9.3005
R7901 VDD.n658 VDD.n571 9.3005
R7902 VDD.n657 VDD.n656 9.3005
R7903 VDD.n653 VDD.n572 9.3005
R7904 VDD.n650 VDD.n649 9.3005
R7905 VDD.n648 VDD.n573 9.3005
R7906 VDD.n647 VDD.n646 9.3005
R7907 VDD.n639 VDD.n638 9.3005
R7908 VDD.n637 VDD.n577 9.3005
R7909 VDD.n636 VDD.n635 9.3005
R7910 VDD.n632 VDD.n578 9.3005
R7911 VDD.n629 VDD.n628 9.3005
R7912 VDD.n627 VDD.n579 9.3005
R7913 VDD.n626 VDD.n625 9.3005
R7914 VDD.n622 VDD.n580 9.3005
R7915 VDD.n619 VDD.n618 9.3005
R7916 VDD.n617 VDD.n581 9.3005
R7917 VDD.n616 VDD.n615 9.3005
R7918 VDD.n612 VDD.n582 9.3005
R7919 VDD.n607 VDD.n586 9.3005
R7920 VDD.n606 VDD.n605 9.3005
R7921 VDD.n602 VDD.n587 9.3005
R7922 VDD.n599 VDD.n598 9.3005
R7923 VDD.n597 VDD.n588 9.3005
R7924 VDD.n596 VDD.n595 9.3005
R7925 VDD.n592 VDD.n590 9.3005
R7926 VDD.n589 VDD.n545 9.3005
R7927 VDD.n4245 VDD.n544 9.3005
R7928 VDD.n609 VDD.n608 9.3005
R7929 VDD.n642 VDD.n574 9.3005
R7930 VDD.n675 VDD.n674 9.3005
R7931 VDD.n4240 VDD.n4239 9.3005
R7932 VDD.n2609 VDD.n2608 9.3005
R7933 VDD.n2610 VDD.n2025 9.3005
R7934 VDD.n2612 VDD.n2611 9.3005
R7935 VDD.n2015 VDD.n2014 9.3005
R7936 VDD.n2625 VDD.n2624 9.3005
R7937 VDD.n2626 VDD.n2013 9.3005
R7938 VDD.n2628 VDD.n2627 9.3005
R7939 VDD.n2003 VDD.n2002 9.3005
R7940 VDD.n2641 VDD.n2640 9.3005
R7941 VDD.n2642 VDD.n2001 9.3005
R7942 VDD.n2644 VDD.n2643 9.3005
R7943 VDD.n1991 VDD.n1990 9.3005
R7944 VDD.n2657 VDD.n2656 9.3005
R7945 VDD.n2658 VDD.n1989 9.3005
R7946 VDD.n2660 VDD.n2659 9.3005
R7947 VDD.n1979 VDD.n1978 9.3005
R7948 VDD.n2673 VDD.n2672 9.3005
R7949 VDD.n2674 VDD.n1977 9.3005
R7950 VDD.n2676 VDD.n2675 9.3005
R7951 VDD.n1967 VDD.n1966 9.3005
R7952 VDD.n2689 VDD.n2688 9.3005
R7953 VDD.n2690 VDD.n1965 9.3005
R7954 VDD.n2692 VDD.n2691 9.3005
R7955 VDD.n1955 VDD.n1954 9.3005
R7956 VDD.n2705 VDD.n2704 9.3005
R7957 VDD.n2706 VDD.n1953 9.3005
R7958 VDD.n2708 VDD.n2707 9.3005
R7959 VDD.n1943 VDD.n1942 9.3005
R7960 VDD.n2721 VDD.n2720 9.3005
R7961 VDD.n2722 VDD.n1941 9.3005
R7962 VDD.n2724 VDD.n2723 9.3005
R7963 VDD.n1931 VDD.n1930 9.3005
R7964 VDD.n2737 VDD.n2736 9.3005
R7965 VDD.n2738 VDD.n1929 9.3005
R7966 VDD.n2740 VDD.n2739 9.3005
R7967 VDD.n1919 VDD.n1918 9.3005
R7968 VDD.n2753 VDD.n2752 9.3005
R7969 VDD.n2754 VDD.n1917 9.3005
R7970 VDD.n2756 VDD.n2755 9.3005
R7971 VDD.n1907 VDD.n1906 9.3005
R7972 VDD.n2769 VDD.n2768 9.3005
R7973 VDD.n2770 VDD.n1905 9.3005
R7974 VDD.n2772 VDD.n2771 9.3005
R7975 VDD.n1895 VDD.n1894 9.3005
R7976 VDD.n2785 VDD.n2784 9.3005
R7977 VDD.n2786 VDD.n1893 9.3005
R7978 VDD.n2788 VDD.n2787 9.3005
R7979 VDD.n1883 VDD.n1882 9.3005
R7980 VDD.n2801 VDD.n2800 9.3005
R7981 VDD.n2802 VDD.n1881 9.3005
R7982 VDD.n2804 VDD.n2803 9.3005
R7983 VDD.n1870 VDD.n1869 9.3005
R7984 VDD.n2818 VDD.n2817 9.3005
R7985 VDD.n2819 VDD.n1868 9.3005
R7986 VDD.n2821 VDD.n2820 9.3005
R7987 VDD.n1857 VDD.n1856 9.3005
R7988 VDD.n2838 VDD.n2837 9.3005
R7989 VDD.n2839 VDD.n1855 9.3005
R7990 VDD.n2841 VDD.n2840 9.3005
R7991 VDD.n2847 VDD.n2846 9.3005
R7992 VDD.n2850 VDD.n1853 9.3005
R7993 VDD.n2854 VDD.n2853 9.3005
R7994 VDD.n2855 VDD.n1852 9.3005
R7995 VDD.n2857 VDD.n2856 9.3005
R7996 VDD.n2860 VDD.n1851 9.3005
R7997 VDD.n2864 VDD.n2863 9.3005
R7998 VDD.n2865 VDD.n1850 9.3005
R7999 VDD.n2867 VDD.n2866 9.3005
R8000 VDD.n2870 VDD.n1849 9.3005
R8001 VDD.n2877 VDD.n2876 9.3005
R8002 VDD.n2878 VDD.n1848 9.3005
R8003 VDD.n2880 VDD.n2879 9.3005
R8004 VDD.n2883 VDD.n1847 9.3005
R8005 VDD.n2887 VDD.n2886 9.3005
R8006 VDD.n2888 VDD.n1846 9.3005
R8007 VDD.n2890 VDD.n2889 9.3005
R8008 VDD.n1807 VDD.n1805 9.3005
R8009 VDD.n2938 VDD.n2937 9.3005
R8010 VDD.n2936 VDD.n1806 9.3005
R8011 VDD.n2935 VDD.n2934 9.3005
R8012 VDD.n2933 VDD.n1811 9.3005
R8013 VDD.n2932 VDD.n2931 9.3005
R8014 VDD.n2929 VDD.n1812 9.3005
R8015 VDD.n2928 VDD.n2927 9.3005
R8016 VDD.n2926 VDD.n1818 9.3005
R8017 VDD.n2925 VDD.n2924 9.3005
R8018 VDD.n2923 VDD.n1819 9.3005
R8019 VDD.n2922 VDD.n2921 9.3005
R8020 VDD.n2920 VDD.n1823 9.3005
R8021 VDD.n2919 VDD.n2918 9.3005
R8022 VDD.n2917 VDD.n1824 9.3005
R8023 VDD.n2916 VDD.n2915 9.3005
R8024 VDD.n2914 VDD.n1828 9.3005
R8025 VDD.n2913 VDD.n2912 9.3005
R8026 VDD.n2911 VDD.n1829 9.3005
R8027 VDD.n2909 VDD.n1834 9.3005
R8028 VDD.n2845 VDD.n2844 9.3005
R8029 VDD.n2376 VDD.n2375 9.3005
R8030 VDD.n2377 VDD.n2220 9.3005
R8031 VDD.n2379 VDD.n2378 9.3005
R8032 VDD.n2209 VDD.n2208 9.3005
R8033 VDD.n2392 VDD.n2391 9.3005
R8034 VDD.n2393 VDD.n2207 9.3005
R8035 VDD.n2395 VDD.n2394 9.3005
R8036 VDD.n2198 VDD.n2197 9.3005
R8037 VDD.n2408 VDD.n2407 9.3005
R8038 VDD.n2409 VDD.n2196 9.3005
R8039 VDD.n2411 VDD.n2410 9.3005
R8040 VDD.n2186 VDD.n2185 9.3005
R8041 VDD.n2424 VDD.n2423 9.3005
R8042 VDD.n2425 VDD.n2184 9.3005
R8043 VDD.n2427 VDD.n2426 9.3005
R8044 VDD.n2174 VDD.n2173 9.3005
R8045 VDD.n2440 VDD.n2439 9.3005
R8046 VDD.n2441 VDD.n2172 9.3005
R8047 VDD.n2443 VDD.n2442 9.3005
R8048 VDD.n2162 VDD.n2161 9.3005
R8049 VDD.n2456 VDD.n2455 9.3005
R8050 VDD.n2457 VDD.n2160 9.3005
R8051 VDD.n2459 VDD.n2458 9.3005
R8052 VDD.n2150 VDD.n2149 9.3005
R8053 VDD.n2472 VDD.n2471 9.3005
R8054 VDD.n2473 VDD.n2148 9.3005
R8055 VDD.n2475 VDD.n2474 9.3005
R8056 VDD.n2138 VDD.n2137 9.3005
R8057 VDD.n2488 VDD.n2487 9.3005
R8058 VDD.n2489 VDD.n2136 9.3005
R8059 VDD.n2491 VDD.n2490 9.3005
R8060 VDD.n2126 VDD.n2125 9.3005
R8061 VDD.n2504 VDD.n2503 9.3005
R8062 VDD.n2505 VDD.n2124 9.3005
R8063 VDD.n2507 VDD.n2506 9.3005
R8064 VDD.n2114 VDD.n2113 9.3005
R8065 VDD.n2520 VDD.n2519 9.3005
R8066 VDD.n2521 VDD.n2112 9.3005
R8067 VDD.n2523 VDD.n2522 9.3005
R8068 VDD.n2102 VDD.n2101 9.3005
R8069 VDD.n2536 VDD.n2535 9.3005
R8070 VDD.n2537 VDD.n2100 9.3005
R8071 VDD.n2539 VDD.n2538 9.3005
R8072 VDD.n2089 VDD.n2088 9.3005
R8073 VDD.n2552 VDD.n2551 9.3005
R8074 VDD.n2553 VDD.n2087 9.3005
R8075 VDD.n2555 VDD.n2554 9.3005
R8076 VDD.n2078 VDD.n2077 9.3005
R8077 VDD.n2568 VDD.n2567 9.3005
R8078 VDD.n2569 VDD.n2076 9.3005
R8079 VDD.n2571 VDD.n2570 9.3005
R8080 VDD.n2066 VDD.n2065 9.3005
R8081 VDD.n2584 VDD.n2583 9.3005
R8082 VDD.n2585 VDD.n2064 9.3005
R8083 VDD.n2587 VDD.n2586 9.3005
R8084 VDD.n2053 VDD.n2052 9.3005
R8085 VDD.n2601 VDD.n2600 9.3005
R8086 VDD.n2602 VDD.n2051 9.3005
R8087 VDD.n2604 VDD.n2603 9.3005
R8088 VDD.n2021 VDD.n2020 9.3005
R8089 VDD.n2617 VDD.n2616 9.3005
R8090 VDD.n2618 VDD.n2019 9.3005
R8091 VDD.n2620 VDD.n2619 9.3005
R8092 VDD.n2009 VDD.n2008 9.3005
R8093 VDD.n2633 VDD.n2632 9.3005
R8094 VDD.n2634 VDD.n2007 9.3005
R8095 VDD.n2636 VDD.n2635 9.3005
R8096 VDD.n1996 VDD.n1995 9.3005
R8097 VDD.n2649 VDD.n2648 9.3005
R8098 VDD.n2650 VDD.n1994 9.3005
R8099 VDD.n2652 VDD.n2651 9.3005
R8100 VDD.n1985 VDD.n1984 9.3005
R8101 VDD.n2665 VDD.n2664 9.3005
R8102 VDD.n2666 VDD.n1983 9.3005
R8103 VDD.n2668 VDD.n2667 9.3005
R8104 VDD.n1973 VDD.n1972 9.3005
R8105 VDD.n2681 VDD.n2680 9.3005
R8106 VDD.n2682 VDD.n1971 9.3005
R8107 VDD.n2684 VDD.n2683 9.3005
R8108 VDD.n1961 VDD.n1960 9.3005
R8109 VDD.n2697 VDD.n2696 9.3005
R8110 VDD.n2698 VDD.n1959 9.3005
R8111 VDD.n2700 VDD.n2699 9.3005
R8112 VDD.n1949 VDD.n1948 9.3005
R8113 VDD.n2713 VDD.n2712 9.3005
R8114 VDD.n2714 VDD.n1947 9.3005
R8115 VDD.n2716 VDD.n2715 9.3005
R8116 VDD.n1937 VDD.n1936 9.3005
R8117 VDD.n2729 VDD.n2728 9.3005
R8118 VDD.n2730 VDD.n1935 9.3005
R8119 VDD.n2732 VDD.n2731 9.3005
R8120 VDD.n1925 VDD.n1924 9.3005
R8121 VDD.n2745 VDD.n2744 9.3005
R8122 VDD.n2746 VDD.n1923 9.3005
R8123 VDD.n2748 VDD.n2747 9.3005
R8124 VDD.n1913 VDD.n1912 9.3005
R8125 VDD.n2761 VDD.n2760 9.3005
R8126 VDD.n2762 VDD.n1911 9.3005
R8127 VDD.n2764 VDD.n2763 9.3005
R8128 VDD.n1901 VDD.n1900 9.3005
R8129 VDD.n2777 VDD.n2776 9.3005
R8130 VDD.n2778 VDD.n1899 9.3005
R8131 VDD.n2780 VDD.n2779 9.3005
R8132 VDD.n1889 VDD.n1888 9.3005
R8133 VDD.n2793 VDD.n2792 9.3005
R8134 VDD.n2794 VDD.n1887 9.3005
R8135 VDD.n2796 VDD.n2795 9.3005
R8136 VDD.n1876 VDD.n1875 9.3005
R8137 VDD.n2809 VDD.n2808 9.3005
R8138 VDD.n2810 VDD.n1873 9.3005
R8139 VDD.n2813 VDD.n2812 9.3005
R8140 VDD.n2811 VDD.n1874 9.3005
R8141 VDD.n1864 VDD.n1863 9.3005
R8142 VDD.n2827 VDD.n2826 9.3005
R8143 VDD.n2828 VDD.n1861 9.3005
R8144 VDD.n2832 VDD.n2831 9.3005
R8145 VDD.n2830 VDD.n1862 9.3005
R8146 VDD.n2222 VDD.n2221 9.3005
R8147 VDD.n2309 VDD.n2308 9.3005
R8148 VDD.n2310 VDD.n2297 9.3005
R8149 VDD.n2312 VDD.n2311 9.3005
R8150 VDD.n2313 VDD.n2292 9.3005
R8151 VDD.n2315 VDD.n2314 9.3005
R8152 VDD.n2316 VDD.n2291 9.3005
R8153 VDD.n2318 VDD.n2317 9.3005
R8154 VDD.n2319 VDD.n2286 9.3005
R8155 VDD.n2321 VDD.n2320 9.3005
R8156 VDD.n2322 VDD.n2285 9.3005
R8157 VDD.n2324 VDD.n2323 9.3005
R8158 VDD.n2325 VDD.n2280 9.3005
R8159 VDD.n2331 VDD.n2279 9.3005
R8160 VDD.n2333 VDD.n2332 9.3005
R8161 VDD.n2334 VDD.n2274 9.3005
R8162 VDD.n2336 VDD.n2335 9.3005
R8163 VDD.n2337 VDD.n2273 9.3005
R8164 VDD.n2339 VDD.n2338 9.3005
R8165 VDD.n2340 VDD.n2268 9.3005
R8166 VDD.n2342 VDD.n2341 9.3005
R8167 VDD.n2343 VDD.n2267 9.3005
R8168 VDD.n2345 VDD.n2344 9.3005
R8169 VDD.n2346 VDD.n2263 9.3005
R8170 VDD.n2348 VDD.n2347 9.3005
R8171 VDD.n2351 VDD.n2256 9.3005
R8172 VDD.n2353 VDD.n2352 9.3005
R8173 VDD.n2354 VDD.n2255 9.3005
R8174 VDD.n2356 VDD.n2355 9.3005
R8175 VDD.n2357 VDD.n2250 9.3005
R8176 VDD.n2359 VDD.n2358 9.3005
R8177 VDD.n2360 VDD.n2249 9.3005
R8178 VDD.n2362 VDD.n2361 9.3005
R8179 VDD.n2228 VDD.n2227 9.3005
R8180 VDD.n2368 VDD.n2367 9.3005
R8181 VDD.n2350 VDD.n2349 9.3005
R8182 VDD.n2330 VDD.n2329 9.3005
R8183 VDD.n2307 VDD.n2298 9.3005
R8184 VDD.n2303 VDD.n2302 9.3005
R8185 VDD.n2371 VDD.n2370 9.3005
R8186 VDD.n2216 VDD.n2215 9.3005
R8187 VDD.n2384 VDD.n2383 9.3005
R8188 VDD.n2385 VDD.n2214 9.3005
R8189 VDD.n2387 VDD.n2386 9.3005
R8190 VDD.n2204 VDD.n2203 9.3005
R8191 VDD.n2400 VDD.n2399 9.3005
R8192 VDD.n2401 VDD.n2202 9.3005
R8193 VDD.n2403 VDD.n2402 9.3005
R8194 VDD.n2192 VDD.n2191 9.3005
R8195 VDD.n2416 VDD.n2415 9.3005
R8196 VDD.n2417 VDD.n2190 9.3005
R8197 VDD.n2419 VDD.n2418 9.3005
R8198 VDD.n2180 VDD.n2179 9.3005
R8199 VDD.n2432 VDD.n2431 9.3005
R8200 VDD.n2433 VDD.n2178 9.3005
R8201 VDD.n2435 VDD.n2434 9.3005
R8202 VDD.n2168 VDD.n2167 9.3005
R8203 VDD.n2448 VDD.n2447 9.3005
R8204 VDD.n2449 VDD.n2166 9.3005
R8205 VDD.n2451 VDD.n2450 9.3005
R8206 VDD.n2156 VDD.n2155 9.3005
R8207 VDD.n2464 VDD.n2463 9.3005
R8208 VDD.n2465 VDD.n2154 9.3005
R8209 VDD.n2467 VDD.n2466 9.3005
R8210 VDD.n2144 VDD.n2143 9.3005
R8211 VDD.n2480 VDD.n2479 9.3005
R8212 VDD.n2481 VDD.n2142 9.3005
R8213 VDD.n2483 VDD.n2482 9.3005
R8214 VDD.n2132 VDD.n2131 9.3005
R8215 VDD.n2496 VDD.n2495 9.3005
R8216 VDD.n2497 VDD.n2130 9.3005
R8217 VDD.n2499 VDD.n2498 9.3005
R8218 VDD.n2120 VDD.n2119 9.3005
R8219 VDD.n2512 VDD.n2511 9.3005
R8220 VDD.n2513 VDD.n2118 9.3005
R8221 VDD.n2515 VDD.n2514 9.3005
R8222 VDD.n2108 VDD.n2107 9.3005
R8223 VDD.n2528 VDD.n2527 9.3005
R8224 VDD.n2529 VDD.n2106 9.3005
R8225 VDD.n2531 VDD.n2530 9.3005
R8226 VDD.n2096 VDD.n2095 9.3005
R8227 VDD.n2544 VDD.n2543 9.3005
R8228 VDD.n2545 VDD.n2094 9.3005
R8229 VDD.n2547 VDD.n2546 9.3005
R8230 VDD.n2084 VDD.n2083 9.3005
R8231 VDD.n2560 VDD.n2559 9.3005
R8232 VDD.n2561 VDD.n2082 9.3005
R8233 VDD.n2563 VDD.n2562 9.3005
R8234 VDD.n2072 VDD.n2071 9.3005
R8235 VDD.n2576 VDD.n2575 9.3005
R8236 VDD.n2577 VDD.n2070 9.3005
R8237 VDD.n2579 VDD.n2578 9.3005
R8238 VDD.n2060 VDD.n2059 9.3005
R8239 VDD.n2592 VDD.n2591 9.3005
R8240 VDD.n2593 VDD.n2058 9.3005
R8241 VDD.n2596 VDD.n2595 9.3005
R8242 VDD.n2594 VDD.n2048 9.3005
R8243 VDD.n2369 VDD.n2226 9.3005
R8244 VDD.n1117 VDD.t85 9.0852
R8245 VDD.n3859 VDD.t76 9.0852
R8246 VDD.n3432 VDD.n3431 9.05416
R8247 VDD.n4181 VDD.n711 9.05416
R8248 VDD.n4225 VDD.n4224 9.05416
R8249 VDD.n3782 VDD.n3781 9.05416
R8250 VDD.n3353 VDD.n1063 9.05416
R8251 VDD.n1585 VDD.n1411 9.05416
R8252 VDD.n3297 VDD.n1081 9.05416
R8253 VDD.n1791 VDD.n1790 9.05416
R8254 VDD.n2397 VDD.t33 8.76075
R8255 VDD.n1879 VDD.t22 8.76075
R8256 VDD.n4276 VDD.t29 8.76075
R8257 VDD.n4609 VDD.t9 8.76075
R8258 VDD.n3078 VDD.t94 8.43629
R8259 VDD.n3132 VDD.t96 8.43629
R8260 VDD.t82 VDD.n874 8.43629
R8261 VDD.n828 VDD.t92 8.43629
R8262 VDD.n15 VDD.n14 8.30123
R8263 VDD.n4713 VDD.n4712 8.1675
R8264 VDD.n2047 VDD.n2046 8.1675
R8265 VDD.n2056 VDD.t110 8.11184
R8266 VDD.n2606 VDD.t110 8.11184
R8267 VDD.n3000 VDD.t5 8.11184
R8268 VDD.n1110 VDD.t44 8.11184
R8269 VDD.n3853 VDD.t63 8.11184
R8270 VDD.n750 VDD.t40 8.11184
R8271 VDD.n4484 VDD.t122 8.11184
R8272 VDD.t122 VDD.n42 8.11184
R8273 VDD.t160 VDD.n1366 7.78739
R8274 VDD.t100 VDD.n1163 7.78739
R8275 VDD.n3913 VDD.t98 7.78739
R8276 VDD.n4117 VDD.t158 7.78739
R8277 VDD.n2212 VDD.t33 7.46293
R8278 VDD.n2815 VDD.t22 7.46293
R8279 VDD.n526 VDD.t29 7.46293
R8280 VDD.n185 VDD.t9 7.46293
R8281 VDD.t120 VDD.n2158 6.48957
R8282 VDD.n2750 VDD.t112 6.48957
R8283 VDD.t118 VDD.n472 6.48957
R8284 VDD.t104 VDD.n134 6.48957
R8285 VDD.n2038 VDD.n2031 6.45596
R8286 VDD.n2306 VDD.n2303 6.4005
R8287 VDD.n2328 VDD.n2325 6.4005
R8288 VDD.n2347 VDD.n2262 6.4005
R8289 VDD.n4240 VDD.n567 6.4005
R8290 VDD.n646 VDD.n643 6.4005
R8291 VDD.n612 VDD.n585 6.4005
R8292 VDD.n4590 VDD.n220 6.4005
R8293 VDD.n307 VDD.n230 6.4005
R8294 VDD.n274 VDD.n273 6.4005
R8295 VDD.n2876 VDD.n2873 6.4005
R8296 VDD.n2930 VDD.n2929 6.4005
R8297 VDD.n2910 VDD.n2909 6.4005
R8298 VDD.n4239 VDD.n541 6.02489
R8299 VDD.n4247 VDD.n541 5.87855
R8300 VDD.n28 VDD.n21 5.57234
R8301 VDD.n2045 VDD.n2044 5.52205
R8302 VDD.n2038 VDD.n2037 5.52205
R8303 VDD.n3126 VDD.t2 5.51621
R8304 VDD.t2 VDD.n1229 5.51621
R8305 VDD.n3979 VDD.t72 5.51621
R8306 VDD.t72 VDD.n868 5.51621
R8307 VDD.n2940 VDD.n2939 5.41513
R8308 VDD.n2939 VDD.n1804 5.41513
R8309 VDD.n4713 VDD.n35 5.28188
R8310 VDD.n2046 VDD.n2045 5.28188
R8311 VDD.n35 VDD.n34 4.63843
R8312 VDD.n28 VDD.n27 4.63843
R8313 VDD.n2092 VDD.t131 3.24504
R8314 VDD.n2654 VDD.t114 3.24504
R8315 VDD.n2988 VDD.t160 3.24504
R8316 VDD.n3192 VDD.t100 3.24504
R8317 VDD.t98 VDD.n934 3.24504
R8318 VDD.t158 VDD.n730 3.24504
R8319 VDD.n406 VDD.t107 3.24504
R8320 VDD.n75 VDD.t128 3.24504
R8321 VDD.n2046 VDD.n15 3.17598
R8322 VDD VDD.n4713 3.16814
R8323 VDD.n1369 VDD.t5 2.92058
R8324 VDD.n3258 VDD.t44 2.92058
R8325 VDD.n1008 VDD.t63 2.92058
R8326 VDD.n4111 VDD.t40 2.92058
R8327 VDD.n1291 VDD.t94 2.59613
R8328 VDD.t96 VDD.n1223 2.59613
R8329 VDD.n3973 VDD.t82 2.59613
R8330 VDD.n4033 VDD.t92 2.59613
R8331 VDD.n4 VDD.n2 2.36832
R8332 VDD.n11 VDD.n9 2.36832
R8333 VDD.n3252 VDD.t85 1.94722
R8334 VDD.n1001 VDD.t76 1.94722
R8335 VDD.n6 VDD.n4 1.90855
R8336 VDD.n13 VDD.n11 1.90855
R8337 VDD.n33 VDD.n31 1.76774
R8338 VDD.n34 VDD.n33 1.76774
R8339 VDD.n26 VDD.n24 1.76774
R8340 VDD.n27 VDD.n26 1.76774
R8341 VDD.n20 VDD.n18 1.76774
R8342 VDD.n21 VDD.n20 1.76774
R8343 VDD.n2044 VDD.n2042 1.76774
R8344 VDD.n2042 VDD.n2040 1.76774
R8345 VDD.n2037 VDD.n2035 1.76774
R8346 VDD.n2035 VDD.n2033 1.76774
R8347 VDD.n2031 VDD.n2029 1.76774
R8348 VDD.n2029 VDD.n2027 1.76774
R8349 VDD.t126 VDD.n2122 1.62277
R8350 VDD.n2702 VDD.t102 1.62277
R8351 VDD.t141 VDD.n436 1.62277
R8352 VDD.t138 VDD.n101 1.62277
R8353 VDD.n3433 VDD.n3432 1.56148
R8354 VDD.n713 VDD.n711 1.56148
R8355 VDD.n4224 VDD.n4223 1.56148
R8356 VDD.n3781 VDD.n3780 1.56148
R8357 VDD.n3350 VDD.n1063 1.56148
R8358 VDD.n1581 VDD.n1411 1.56148
R8359 VDD.n3294 VDD.n1081 1.56148
R8360 VDD.n1790 VDD.n1789 1.56148
R8361 VDD.n14 VDD.n6 1.47464
R8362 VDD.n14 VDD.n13 1.47464
R8363 VDD.n35 VDD.n28 0.934408
R8364 VDD.n2045 VDD.n2038 0.934408
R8365 VDD.n4248 VDD.n4247 0.572146
R8366 VDD.n2840 VDD.n1595 0.572146
R8367 VDD.n4589 VDD.n4588 0.521842
R8368 VDD.n247 VDD.n244 0.521842
R8369 VDD.n2302 VDD.n2221 0.521842
R8370 VDD.n2369 VDD.n2368 0.521842
R8371 VDD.n4239 VDD.n535 0.425805
R8372 VDD.n2830 VDD.n2829 0.425805
R8373 VDD.n2829 VDD.n1834 0.384646
R8374 VDD.t84 VDD.n1288 0.324954
R8375 VDD.n3186 VDD.t3 0.324954
R8376 VDD.t91 VDD.n928 0.324954
R8377 VDD.n4039 VDD.t81 0.324954
R8378 VDD.n589 VDD.n544 0.305378
R8379 VDD.n590 VDD.n589 0.305378
R8380 VDD.n596 VDD.n590 0.305378
R8381 VDD.n597 VDD.n596 0.305378
R8382 VDD.n598 VDD.n597 0.305378
R8383 VDD.n598 VDD.n587 0.305378
R8384 VDD.n606 VDD.n587 0.305378
R8385 VDD.n607 VDD.n606 0.305378
R8386 VDD.n608 VDD.n607 0.305378
R8387 VDD.n608 VDD.n582 0.305378
R8388 VDD.n616 VDD.n582 0.305378
R8389 VDD.n617 VDD.n616 0.305378
R8390 VDD.n618 VDD.n617 0.305378
R8391 VDD.n618 VDD.n580 0.305378
R8392 VDD.n626 VDD.n580 0.305378
R8393 VDD.n627 VDD.n626 0.305378
R8394 VDD.n628 VDD.n627 0.305378
R8395 VDD.n636 VDD.n578 0.305378
R8396 VDD.n637 VDD.n636 0.305378
R8397 VDD.n638 VDD.n637 0.305378
R8398 VDD.n638 VDD.n574 0.305378
R8399 VDD.n647 VDD.n574 0.305378
R8400 VDD.n648 VDD.n647 0.305378
R8401 VDD.n649 VDD.n648 0.305378
R8402 VDD.n649 VDD.n572 0.305378
R8403 VDD.n657 VDD.n572 0.305378
R8404 VDD.n658 VDD.n657 0.305378
R8405 VDD.n659 VDD.n658 0.305378
R8406 VDD.n659 VDD.n570 0.305378
R8407 VDD.n667 VDD.n570 0.305378
R8408 VDD.n668 VDD.n667 0.305378
R8409 VDD.n669 VDD.n668 0.305378
R8410 VDD.n669 VDD.n568 0.305378
R8411 VDD.n675 VDD.n568 0.305378
R8412 VDD.n2846 VDD.n2845 0.305378
R8413 VDD.n2846 VDD.n1853 0.305378
R8414 VDD.n2854 VDD.n1853 0.305378
R8415 VDD.n2855 VDD.n2854 0.305378
R8416 VDD.n2856 VDD.n2855 0.305378
R8417 VDD.n2856 VDD.n1851 0.305378
R8418 VDD.n2864 VDD.n1851 0.305378
R8419 VDD.n2865 VDD.n2864 0.305378
R8420 VDD.n2866 VDD.n2865 0.305378
R8421 VDD.n2866 VDD.n1849 0.305378
R8422 VDD.n2877 VDD.n1849 0.305378
R8423 VDD.n2878 VDD.n2877 0.305378
R8424 VDD.n2879 VDD.n2878 0.305378
R8425 VDD.n2879 VDD.n1847 0.305378
R8426 VDD.n2887 VDD.n1847 0.305378
R8427 VDD.n2888 VDD.n2887 0.305378
R8428 VDD.n2889 VDD.n2888 0.305378
R8429 VDD.n2889 VDD.n1805 0.305378
R8430 VDD.n2938 VDD.n1806 0.305378
R8431 VDD.n2934 VDD.n1806 0.305378
R8432 VDD.n2934 VDD.n2933 0.305378
R8433 VDD.n2933 VDD.n2932 0.305378
R8434 VDD.n2932 VDD.n1812 0.305378
R8435 VDD.n2927 VDD.n1812 0.305378
R8436 VDD.n2927 VDD.n2926 0.305378
R8437 VDD.n2926 VDD.n2925 0.305378
R8438 VDD.n2925 VDD.n1819 0.305378
R8439 VDD.n2921 VDD.n1819 0.305378
R8440 VDD.n2921 VDD.n2920 0.305378
R8441 VDD.n2920 VDD.n2919 0.305378
R8442 VDD.n2919 VDD.n1824 0.305378
R8443 VDD.n2915 VDD.n1824 0.305378
R8444 VDD.n2915 VDD.n2914 0.305378
R8445 VDD.n2914 VDD.n2913 0.305378
R8446 VDD.n2913 VDD.n1829 0.305378
R8447 VDD.n1834 VDD.n1829 0.305378
R8448 VDD.n2845 VDD.n1595 0.238305
R8449 VDD.n2307 VDD.n2306 0.194439
R8450 VDD.n2329 VDD.n2328 0.194439
R8451 VDD.n2350 VDD.n2262 0.194439
R8452 VDD.n674 VDD.n567 0.194439
R8453 VDD.n643 VDD.n642 0.194439
R8454 VDD.n609 VDD.n585 0.194439
R8455 VDD.n336 VDD.n220 0.194439
R8456 VDD.n304 VDD.n230 0.194439
R8457 VDD.n273 VDD.n272 0.194439
R8458 VDD.n2873 VDD.n2870 0.194439
R8459 VDD.n2931 VDD.n2930 0.194439
R8460 VDD.n2911 VDD.n2910 0.194439
R8461 VDD.n4255 VDD.n535 0.152939
R8462 VDD.n4256 VDD.n4255 0.152939
R8463 VDD.n4257 VDD.n4256 0.152939
R8464 VDD.n4257 VDD.n522 0.152939
R8465 VDD.n4271 VDD.n522 0.152939
R8466 VDD.n4272 VDD.n4271 0.152939
R8467 VDD.n4273 VDD.n4272 0.152939
R8468 VDD.n4273 VDD.n511 0.152939
R8469 VDD.n4287 VDD.n511 0.152939
R8470 VDD.n4288 VDD.n4287 0.152939
R8471 VDD.n4289 VDD.n4288 0.152939
R8472 VDD.n4289 VDD.n499 0.152939
R8473 VDD.n4303 VDD.n499 0.152939
R8474 VDD.n4304 VDD.n4303 0.152939
R8475 VDD.n4305 VDD.n4304 0.152939
R8476 VDD.n4305 VDD.n487 0.152939
R8477 VDD.n4319 VDD.n487 0.152939
R8478 VDD.n4320 VDD.n4319 0.152939
R8479 VDD.n4321 VDD.n4320 0.152939
R8480 VDD.n4321 VDD.n475 0.152939
R8481 VDD.n4335 VDD.n475 0.152939
R8482 VDD.n4336 VDD.n4335 0.152939
R8483 VDD.n4337 VDD.n4336 0.152939
R8484 VDD.n4337 VDD.n463 0.152939
R8485 VDD.n4351 VDD.n463 0.152939
R8486 VDD.n4352 VDD.n4351 0.152939
R8487 VDD.n4353 VDD.n4352 0.152939
R8488 VDD.n4353 VDD.n451 0.152939
R8489 VDD.n4367 VDD.n451 0.152939
R8490 VDD.n4368 VDD.n4367 0.152939
R8491 VDD.n4369 VDD.n4368 0.152939
R8492 VDD.n4369 VDD.n439 0.152939
R8493 VDD.n4383 VDD.n439 0.152939
R8494 VDD.n4384 VDD.n4383 0.152939
R8495 VDD.n4385 VDD.n4384 0.152939
R8496 VDD.n4385 VDD.n427 0.152939
R8497 VDD.n4399 VDD.n427 0.152939
R8498 VDD.n4400 VDD.n4399 0.152939
R8499 VDD.n4401 VDD.n4400 0.152939
R8500 VDD.n4401 VDD.n415 0.152939
R8501 VDD.n4415 VDD.n415 0.152939
R8502 VDD.n4416 VDD.n4415 0.152939
R8503 VDD.n4417 VDD.n4416 0.152939
R8504 VDD.n4417 VDD.n402 0.152939
R8505 VDD.n4431 VDD.n402 0.152939
R8506 VDD.n4432 VDD.n4431 0.152939
R8507 VDD.n4433 VDD.n4432 0.152939
R8508 VDD.n4433 VDD.n391 0.152939
R8509 VDD.n4447 VDD.n391 0.152939
R8510 VDD.n4448 VDD.n4447 0.152939
R8511 VDD.n4449 VDD.n4448 0.152939
R8512 VDD.n4450 VDD.n4449 0.152939
R8513 VDD.n4450 VDD.n379 0.152939
R8514 VDD.n4466 VDD.n379 0.152939
R8515 VDD.n4467 VDD.n4466 0.152939
R8516 VDD.n4468 VDD.n4467 0.152939
R8517 VDD.n4470 VDD.n4468 0.152939
R8518 VDD.n4470 VDD.n4469 0.152939
R8519 VDD.n4469 VDD.n368 0.152939
R8520 VDD.n368 VDD.n366 0.152939
R8521 VDD.n4490 VDD.n366 0.152939
R8522 VDD.n4491 VDD.n4490 0.152939
R8523 VDD.n4492 VDD.n4491 0.152939
R8524 VDD.n4492 VDD.n364 0.152939
R8525 VDD.n4497 VDD.n364 0.152939
R8526 VDD.n4498 VDD.n4497 0.152939
R8527 VDD.n4499 VDD.n4498 0.152939
R8528 VDD.n4499 VDD.n362 0.152939
R8529 VDD.n4504 VDD.n362 0.152939
R8530 VDD.n4505 VDD.n4504 0.152939
R8531 VDD.n4506 VDD.n4505 0.152939
R8532 VDD.n4506 VDD.n360 0.152939
R8533 VDD.n4511 VDD.n360 0.152939
R8534 VDD.n4512 VDD.n4511 0.152939
R8535 VDD.n4513 VDD.n4512 0.152939
R8536 VDD.n4513 VDD.n358 0.152939
R8537 VDD.n4518 VDD.n358 0.152939
R8538 VDD.n4519 VDD.n4518 0.152939
R8539 VDD.n4520 VDD.n4519 0.152939
R8540 VDD.n4520 VDD.n356 0.152939
R8541 VDD.n4525 VDD.n356 0.152939
R8542 VDD.n4526 VDD.n4525 0.152939
R8543 VDD.n4527 VDD.n4526 0.152939
R8544 VDD.n4527 VDD.n354 0.152939
R8545 VDD.n4532 VDD.n354 0.152939
R8546 VDD.n4533 VDD.n4532 0.152939
R8547 VDD.n4534 VDD.n4533 0.152939
R8548 VDD.n4534 VDD.n352 0.152939
R8549 VDD.n4539 VDD.n352 0.152939
R8550 VDD.n4540 VDD.n4539 0.152939
R8551 VDD.n4541 VDD.n4540 0.152939
R8552 VDD.n4541 VDD.n350 0.152939
R8553 VDD.n4546 VDD.n350 0.152939
R8554 VDD.n4547 VDD.n4546 0.152939
R8555 VDD.n4548 VDD.n4547 0.152939
R8556 VDD.n4548 VDD.n348 0.152939
R8557 VDD.n4553 VDD.n348 0.152939
R8558 VDD.n4554 VDD.n4553 0.152939
R8559 VDD.n4555 VDD.n4554 0.152939
R8560 VDD.n4555 VDD.n346 0.152939
R8561 VDD.n4560 VDD.n346 0.152939
R8562 VDD.n4561 VDD.n4560 0.152939
R8563 VDD.n4562 VDD.n4561 0.152939
R8564 VDD.n4562 VDD.n344 0.152939
R8565 VDD.n4567 VDD.n344 0.152939
R8566 VDD.n4568 VDD.n4567 0.152939
R8567 VDD.n4569 VDD.n4568 0.152939
R8568 VDD.n4569 VDD.n342 0.152939
R8569 VDD.n4574 VDD.n342 0.152939
R8570 VDD.n4575 VDD.n4574 0.152939
R8571 VDD.n4576 VDD.n4575 0.152939
R8572 VDD.n4576 VDD.n340 0.152939
R8573 VDD.n4581 VDD.n340 0.152939
R8574 VDD.n4582 VDD.n4581 0.152939
R8575 VDD.n4583 VDD.n4582 0.152939
R8576 VDD.n4583 VDD.n338 0.152939
R8577 VDD.n4588 VDD.n338 0.152939
R8578 VDD.n248 VDD.n247 0.152939
R8579 VDD.n249 VDD.n248 0.152939
R8580 VDD.n249 VDD.n242 0.152939
R8581 VDD.n257 VDD.n242 0.152939
R8582 VDD.n258 VDD.n257 0.152939
R8583 VDD.n259 VDD.n258 0.152939
R8584 VDD.n259 VDD.n240 0.152939
R8585 VDD.n267 VDD.n240 0.152939
R8586 VDD.n268 VDD.n267 0.152939
R8587 VDD.n269 VDD.n268 0.152939
R8588 VDD.n269 VDD.n236 0.152939
R8589 VDD.n278 VDD.n236 0.152939
R8590 VDD.n279 VDD.n278 0.152939
R8591 VDD.n280 VDD.n279 0.152939
R8592 VDD.n280 VDD.n234 0.152939
R8593 VDD.n288 VDD.n234 0.152939
R8594 VDD.n289 VDD.n288 0.152939
R8595 VDD.n290 VDD.n289 0.152939
R8596 VDD.n290 VDD.n232 0.152939
R8597 VDD.n298 VDD.n232 0.152939
R8598 VDD.n299 VDD.n298 0.152939
R8599 VDD.n300 VDD.n299 0.152939
R8600 VDD.n300 VDD.n227 0.152939
R8601 VDD.n308 VDD.n227 0.152939
R8602 VDD.n309 VDD.n308 0.152939
R8603 VDD.n310 VDD.n309 0.152939
R8604 VDD.n310 VDD.n225 0.152939
R8605 VDD.n318 VDD.n225 0.152939
R8606 VDD.n319 VDD.n318 0.152939
R8607 VDD.n320 VDD.n319 0.152939
R8608 VDD.n320 VDD.n223 0.152939
R8609 VDD.n328 VDD.n223 0.152939
R8610 VDD.n329 VDD.n328 0.152939
R8611 VDD.n330 VDD.n329 0.152939
R8612 VDD.n330 VDD.n221 0.152939
R8613 VDD.n337 VDD.n221 0.152939
R8614 VDD.n4589 VDD.n337 0.152939
R8615 VDD.n4711 VDD.n37 0.152939
R8616 VDD.n48 VDD.n37 0.152939
R8617 VDD.n49 VDD.n48 0.152939
R8618 VDD.n50 VDD.n49 0.152939
R8619 VDD.n51 VDD.n50 0.152939
R8620 VDD.n59 VDD.n51 0.152939
R8621 VDD.n60 VDD.n59 0.152939
R8622 VDD.n61 VDD.n60 0.152939
R8623 VDD.n62 VDD.n61 0.152939
R8624 VDD.n69 VDD.n62 0.152939
R8625 VDD.n70 VDD.n69 0.152939
R8626 VDD.n71 VDD.n70 0.152939
R8627 VDD.n72 VDD.n71 0.152939
R8628 VDD.n81 VDD.n72 0.152939
R8629 VDD.n82 VDD.n81 0.152939
R8630 VDD.n83 VDD.n82 0.152939
R8631 VDD.n84 VDD.n83 0.152939
R8632 VDD.n92 VDD.n84 0.152939
R8633 VDD.n93 VDD.n92 0.152939
R8634 VDD.n94 VDD.n93 0.152939
R8635 VDD.n95 VDD.n94 0.152939
R8636 VDD.n103 VDD.n95 0.152939
R8637 VDD.n104 VDD.n103 0.152939
R8638 VDD.n105 VDD.n104 0.152939
R8639 VDD.n106 VDD.n105 0.152939
R8640 VDD.n114 VDD.n106 0.152939
R8641 VDD.n115 VDD.n114 0.152939
R8642 VDD.n116 VDD.n115 0.152939
R8643 VDD.n117 VDD.n116 0.152939
R8644 VDD.n125 VDD.n117 0.152939
R8645 VDD.n126 VDD.n125 0.152939
R8646 VDD.n127 VDD.n126 0.152939
R8647 VDD.n128 VDD.n127 0.152939
R8648 VDD.n136 VDD.n128 0.152939
R8649 VDD.n137 VDD.n136 0.152939
R8650 VDD.n138 VDD.n137 0.152939
R8651 VDD.n139 VDD.n138 0.152939
R8652 VDD.n147 VDD.n139 0.152939
R8653 VDD.n148 VDD.n147 0.152939
R8654 VDD.n149 VDD.n148 0.152939
R8655 VDD.n150 VDD.n149 0.152939
R8656 VDD.n158 VDD.n150 0.152939
R8657 VDD.n159 VDD.n158 0.152939
R8658 VDD.n160 VDD.n159 0.152939
R8659 VDD.n161 VDD.n160 0.152939
R8660 VDD.n169 VDD.n161 0.152939
R8661 VDD.n170 VDD.n169 0.152939
R8662 VDD.n171 VDD.n170 0.152939
R8663 VDD.n172 VDD.n171 0.152939
R8664 VDD.n179 VDD.n172 0.152939
R8665 VDD.n180 VDD.n179 0.152939
R8666 VDD.n181 VDD.n180 0.152939
R8667 VDD.n182 VDD.n181 0.152939
R8668 VDD.n191 VDD.n182 0.152939
R8669 VDD.n192 VDD.n191 0.152939
R8670 VDD.n193 VDD.n192 0.152939
R8671 VDD.n194 VDD.n193 0.152939
R8672 VDD.n244 VDD.n194 0.152939
R8673 VDD.n4249 VDD.n4248 0.152939
R8674 VDD.n4249 VDD.n529 0.152939
R8675 VDD.n4263 VDD.n529 0.152939
R8676 VDD.n4264 VDD.n4263 0.152939
R8677 VDD.n4265 VDD.n4264 0.152939
R8678 VDD.n4265 VDD.n517 0.152939
R8679 VDD.n4279 VDD.n517 0.152939
R8680 VDD.n4280 VDD.n4279 0.152939
R8681 VDD.n4281 VDD.n4280 0.152939
R8682 VDD.n4281 VDD.n505 0.152939
R8683 VDD.n4295 VDD.n505 0.152939
R8684 VDD.n4296 VDD.n4295 0.152939
R8685 VDD.n4297 VDD.n4296 0.152939
R8686 VDD.n4297 VDD.n493 0.152939
R8687 VDD.n4311 VDD.n493 0.152939
R8688 VDD.n4312 VDD.n4311 0.152939
R8689 VDD.n4313 VDD.n4312 0.152939
R8690 VDD.n4313 VDD.n481 0.152939
R8691 VDD.n4327 VDD.n481 0.152939
R8692 VDD.n4328 VDD.n4327 0.152939
R8693 VDD.n4329 VDD.n4328 0.152939
R8694 VDD.n4329 VDD.n469 0.152939
R8695 VDD.n4343 VDD.n469 0.152939
R8696 VDD.n4344 VDD.n4343 0.152939
R8697 VDD.n4345 VDD.n4344 0.152939
R8698 VDD.n4345 VDD.n457 0.152939
R8699 VDD.n4359 VDD.n457 0.152939
R8700 VDD.n4360 VDD.n4359 0.152939
R8701 VDD.n4361 VDD.n4360 0.152939
R8702 VDD.n4361 VDD.n445 0.152939
R8703 VDD.n4375 VDD.n445 0.152939
R8704 VDD.n4376 VDD.n4375 0.152939
R8705 VDD.n4377 VDD.n4376 0.152939
R8706 VDD.n4377 VDD.n433 0.152939
R8707 VDD.n4391 VDD.n433 0.152939
R8708 VDD.n4392 VDD.n4391 0.152939
R8709 VDD.n4393 VDD.n4392 0.152939
R8710 VDD.n4393 VDD.n421 0.152939
R8711 VDD.n4407 VDD.n421 0.152939
R8712 VDD.n4408 VDD.n4407 0.152939
R8713 VDD.n4409 VDD.n4408 0.152939
R8714 VDD.n4409 VDD.n409 0.152939
R8715 VDD.n4423 VDD.n409 0.152939
R8716 VDD.n4424 VDD.n4423 0.152939
R8717 VDD.n4425 VDD.n4424 0.152939
R8718 VDD.n4425 VDD.n397 0.152939
R8719 VDD.n4439 VDD.n397 0.152939
R8720 VDD.n4440 VDD.n4439 0.152939
R8721 VDD.n4441 VDD.n4440 0.152939
R8722 VDD.n4441 VDD.n385 0.152939
R8723 VDD.n4457 VDD.n385 0.152939
R8724 VDD.n4458 VDD.n4457 0.152939
R8725 VDD.n4459 VDD.n4458 0.152939
R8726 VDD.n4459 VDD.n373 0.152939
R8727 VDD.n4478 VDD.n373 0.152939
R8728 VDD.n4479 VDD.n4478 0.152939
R8729 VDD.n4480 VDD.n4479 0.152939
R8730 VDD.n4480 VDD.n36 0.152939
R8731 VDD.n628 VDD.n541 0.152939
R8732 VDD.n578 VDD.n541 0.152939
R8733 VDD.n2610 VDD.n2609 0.152939
R8734 VDD.n2611 VDD.n2610 0.152939
R8735 VDD.n2611 VDD.n2014 0.152939
R8736 VDD.n2625 VDD.n2014 0.152939
R8737 VDD.n2626 VDD.n2625 0.152939
R8738 VDD.n2627 VDD.n2626 0.152939
R8739 VDD.n2627 VDD.n2002 0.152939
R8740 VDD.n2641 VDD.n2002 0.152939
R8741 VDD.n2642 VDD.n2641 0.152939
R8742 VDD.n2643 VDD.n2642 0.152939
R8743 VDD.n2643 VDD.n1990 0.152939
R8744 VDD.n2657 VDD.n1990 0.152939
R8745 VDD.n2658 VDD.n2657 0.152939
R8746 VDD.n2659 VDD.n2658 0.152939
R8747 VDD.n2659 VDD.n1978 0.152939
R8748 VDD.n2673 VDD.n1978 0.152939
R8749 VDD.n2674 VDD.n2673 0.152939
R8750 VDD.n2675 VDD.n2674 0.152939
R8751 VDD.n2675 VDD.n1966 0.152939
R8752 VDD.n2689 VDD.n1966 0.152939
R8753 VDD.n2690 VDD.n2689 0.152939
R8754 VDD.n2691 VDD.n2690 0.152939
R8755 VDD.n2691 VDD.n1954 0.152939
R8756 VDD.n2705 VDD.n1954 0.152939
R8757 VDD.n2706 VDD.n2705 0.152939
R8758 VDD.n2707 VDD.n2706 0.152939
R8759 VDD.n2707 VDD.n1942 0.152939
R8760 VDD.n2721 VDD.n1942 0.152939
R8761 VDD.n2722 VDD.n2721 0.152939
R8762 VDD.n2723 VDD.n2722 0.152939
R8763 VDD.n2723 VDD.n1930 0.152939
R8764 VDD.n2737 VDD.n1930 0.152939
R8765 VDD.n2738 VDD.n2737 0.152939
R8766 VDD.n2739 VDD.n2738 0.152939
R8767 VDD.n2739 VDD.n1918 0.152939
R8768 VDD.n2753 VDD.n1918 0.152939
R8769 VDD.n2754 VDD.n2753 0.152939
R8770 VDD.n2755 VDD.n2754 0.152939
R8771 VDD.n2755 VDD.n1906 0.152939
R8772 VDD.n2769 VDD.n1906 0.152939
R8773 VDD.n2770 VDD.n2769 0.152939
R8774 VDD.n2771 VDD.n2770 0.152939
R8775 VDD.n2771 VDD.n1894 0.152939
R8776 VDD.n2785 VDD.n1894 0.152939
R8777 VDD.n2786 VDD.n2785 0.152939
R8778 VDD.n2787 VDD.n2786 0.152939
R8779 VDD.n2787 VDD.n1882 0.152939
R8780 VDD.n2801 VDD.n1882 0.152939
R8781 VDD.n2802 VDD.n2801 0.152939
R8782 VDD.n2803 VDD.n2802 0.152939
R8783 VDD.n2803 VDD.n1869 0.152939
R8784 VDD.n2818 VDD.n1869 0.152939
R8785 VDD.n2819 VDD.n2818 0.152939
R8786 VDD.n2820 VDD.n2819 0.152939
R8787 VDD.n2820 VDD.n1856 0.152939
R8788 VDD.n2838 VDD.n1856 0.152939
R8789 VDD.n2839 VDD.n2838 0.152939
R8790 VDD.n2840 VDD.n2839 0.152939
R8791 VDD.n2939 VDD.n1805 0.152939
R8792 VDD.n2939 VDD.n2938 0.152939
R8793 VDD.n2376 VDD.n2221 0.152939
R8794 VDD.n2377 VDD.n2376 0.152939
R8795 VDD.n2378 VDD.n2377 0.152939
R8796 VDD.n2378 VDD.n2208 0.152939
R8797 VDD.n2392 VDD.n2208 0.152939
R8798 VDD.n2393 VDD.n2392 0.152939
R8799 VDD.n2394 VDD.n2393 0.152939
R8800 VDD.n2394 VDD.n2197 0.152939
R8801 VDD.n2408 VDD.n2197 0.152939
R8802 VDD.n2409 VDD.n2408 0.152939
R8803 VDD.n2410 VDD.n2409 0.152939
R8804 VDD.n2410 VDD.n2185 0.152939
R8805 VDD.n2424 VDD.n2185 0.152939
R8806 VDD.n2425 VDD.n2424 0.152939
R8807 VDD.n2426 VDD.n2425 0.152939
R8808 VDD.n2426 VDD.n2173 0.152939
R8809 VDD.n2440 VDD.n2173 0.152939
R8810 VDD.n2441 VDD.n2440 0.152939
R8811 VDD.n2442 VDD.n2441 0.152939
R8812 VDD.n2442 VDD.n2161 0.152939
R8813 VDD.n2456 VDD.n2161 0.152939
R8814 VDD.n2457 VDD.n2456 0.152939
R8815 VDD.n2458 VDD.n2457 0.152939
R8816 VDD.n2458 VDD.n2149 0.152939
R8817 VDD.n2472 VDD.n2149 0.152939
R8818 VDD.n2473 VDD.n2472 0.152939
R8819 VDD.n2474 VDD.n2473 0.152939
R8820 VDD.n2474 VDD.n2137 0.152939
R8821 VDD.n2488 VDD.n2137 0.152939
R8822 VDD.n2489 VDD.n2488 0.152939
R8823 VDD.n2490 VDD.n2489 0.152939
R8824 VDD.n2490 VDD.n2125 0.152939
R8825 VDD.n2504 VDD.n2125 0.152939
R8826 VDD.n2505 VDD.n2504 0.152939
R8827 VDD.n2506 VDD.n2505 0.152939
R8828 VDD.n2506 VDD.n2113 0.152939
R8829 VDD.n2520 VDD.n2113 0.152939
R8830 VDD.n2521 VDD.n2520 0.152939
R8831 VDD.n2522 VDD.n2521 0.152939
R8832 VDD.n2522 VDD.n2101 0.152939
R8833 VDD.n2536 VDD.n2101 0.152939
R8834 VDD.n2537 VDD.n2536 0.152939
R8835 VDD.n2538 VDD.n2537 0.152939
R8836 VDD.n2538 VDD.n2088 0.152939
R8837 VDD.n2552 VDD.n2088 0.152939
R8838 VDD.n2553 VDD.n2552 0.152939
R8839 VDD.n2554 VDD.n2553 0.152939
R8840 VDD.n2554 VDD.n2077 0.152939
R8841 VDD.n2568 VDD.n2077 0.152939
R8842 VDD.n2569 VDD.n2568 0.152939
R8843 VDD.n2570 VDD.n2569 0.152939
R8844 VDD.n2570 VDD.n2065 0.152939
R8845 VDD.n2584 VDD.n2065 0.152939
R8846 VDD.n2585 VDD.n2584 0.152939
R8847 VDD.n2586 VDD.n2585 0.152939
R8848 VDD.n2586 VDD.n2052 0.152939
R8849 VDD.n2601 VDD.n2052 0.152939
R8850 VDD.n2602 VDD.n2601 0.152939
R8851 VDD.n2603 VDD.n2602 0.152939
R8852 VDD.n2603 VDD.n2020 0.152939
R8853 VDD.n2617 VDD.n2020 0.152939
R8854 VDD.n2618 VDD.n2617 0.152939
R8855 VDD.n2619 VDD.n2618 0.152939
R8856 VDD.n2619 VDD.n2008 0.152939
R8857 VDD.n2633 VDD.n2008 0.152939
R8858 VDD.n2634 VDD.n2633 0.152939
R8859 VDD.n2635 VDD.n2634 0.152939
R8860 VDD.n2635 VDD.n1995 0.152939
R8861 VDD.n2649 VDD.n1995 0.152939
R8862 VDD.n2650 VDD.n2649 0.152939
R8863 VDD.n2651 VDD.n2650 0.152939
R8864 VDD.n2651 VDD.n1984 0.152939
R8865 VDD.n2665 VDD.n1984 0.152939
R8866 VDD.n2666 VDD.n2665 0.152939
R8867 VDD.n2667 VDD.n2666 0.152939
R8868 VDD.n2667 VDD.n1972 0.152939
R8869 VDD.n2681 VDD.n1972 0.152939
R8870 VDD.n2682 VDD.n2681 0.152939
R8871 VDD.n2683 VDD.n2682 0.152939
R8872 VDD.n2683 VDD.n1960 0.152939
R8873 VDD.n2697 VDD.n1960 0.152939
R8874 VDD.n2698 VDD.n2697 0.152939
R8875 VDD.n2699 VDD.n2698 0.152939
R8876 VDD.n2699 VDD.n1948 0.152939
R8877 VDD.n2713 VDD.n1948 0.152939
R8878 VDD.n2714 VDD.n2713 0.152939
R8879 VDD.n2715 VDD.n2714 0.152939
R8880 VDD.n2715 VDD.n1936 0.152939
R8881 VDD.n2729 VDD.n1936 0.152939
R8882 VDD.n2730 VDD.n2729 0.152939
R8883 VDD.n2731 VDD.n2730 0.152939
R8884 VDD.n2731 VDD.n1924 0.152939
R8885 VDD.n2745 VDD.n1924 0.152939
R8886 VDD.n2746 VDD.n2745 0.152939
R8887 VDD.n2747 VDD.n2746 0.152939
R8888 VDD.n2747 VDD.n1912 0.152939
R8889 VDD.n2761 VDD.n1912 0.152939
R8890 VDD.n2762 VDD.n2761 0.152939
R8891 VDD.n2763 VDD.n2762 0.152939
R8892 VDD.n2763 VDD.n1900 0.152939
R8893 VDD.n2777 VDD.n1900 0.152939
R8894 VDD.n2778 VDD.n2777 0.152939
R8895 VDD.n2779 VDD.n2778 0.152939
R8896 VDD.n2779 VDD.n1888 0.152939
R8897 VDD.n2793 VDD.n1888 0.152939
R8898 VDD.n2794 VDD.n2793 0.152939
R8899 VDD.n2795 VDD.n2794 0.152939
R8900 VDD.n2795 VDD.n1875 0.152939
R8901 VDD.n2809 VDD.n1875 0.152939
R8902 VDD.n2810 VDD.n2809 0.152939
R8903 VDD.n2812 VDD.n2810 0.152939
R8904 VDD.n2812 VDD.n2811 0.152939
R8905 VDD.n2811 VDD.n1863 0.152939
R8906 VDD.n2827 VDD.n1863 0.152939
R8907 VDD.n2828 VDD.n2827 0.152939
R8908 VDD.n2831 VDD.n2828 0.152939
R8909 VDD.n2831 VDD.n2830 0.152939
R8910 VDD.n2368 VDD.n2227 0.152939
R8911 VDD.n2361 VDD.n2227 0.152939
R8912 VDD.n2361 VDD.n2360 0.152939
R8913 VDD.n2360 VDD.n2359 0.152939
R8914 VDD.n2359 VDD.n2250 0.152939
R8915 VDD.n2355 VDD.n2250 0.152939
R8916 VDD.n2355 VDD.n2354 0.152939
R8917 VDD.n2354 VDD.n2353 0.152939
R8918 VDD.n2353 VDD.n2256 0.152939
R8919 VDD.n2349 VDD.n2256 0.152939
R8920 VDD.n2349 VDD.n2348 0.152939
R8921 VDD.n2348 VDD.n2263 0.152939
R8922 VDD.n2344 VDD.n2263 0.152939
R8923 VDD.n2344 VDD.n2343 0.152939
R8924 VDD.n2343 VDD.n2342 0.152939
R8925 VDD.n2342 VDD.n2268 0.152939
R8926 VDD.n2338 VDD.n2268 0.152939
R8927 VDD.n2338 VDD.n2337 0.152939
R8928 VDD.n2337 VDD.n2336 0.152939
R8929 VDD.n2336 VDD.n2274 0.152939
R8930 VDD.n2332 VDD.n2274 0.152939
R8931 VDD.n2332 VDD.n2331 0.152939
R8932 VDD.n2331 VDD.n2330 0.152939
R8933 VDD.n2330 VDD.n2280 0.152939
R8934 VDD.n2323 VDD.n2280 0.152939
R8935 VDD.n2323 VDD.n2322 0.152939
R8936 VDD.n2322 VDD.n2321 0.152939
R8937 VDD.n2321 VDD.n2286 0.152939
R8938 VDD.n2317 VDD.n2286 0.152939
R8939 VDD.n2317 VDD.n2316 0.152939
R8940 VDD.n2316 VDD.n2315 0.152939
R8941 VDD.n2315 VDD.n2292 0.152939
R8942 VDD.n2311 VDD.n2292 0.152939
R8943 VDD.n2311 VDD.n2310 0.152939
R8944 VDD.n2310 VDD.n2309 0.152939
R8945 VDD.n2309 VDD.n2298 0.152939
R8946 VDD.n2302 VDD.n2298 0.152939
R8947 VDD.n2370 VDD.n2369 0.152939
R8948 VDD.n2370 VDD.n2215 0.152939
R8949 VDD.n2384 VDD.n2215 0.152939
R8950 VDD.n2385 VDD.n2384 0.152939
R8951 VDD.n2386 VDD.n2385 0.152939
R8952 VDD.n2386 VDD.n2203 0.152939
R8953 VDD.n2400 VDD.n2203 0.152939
R8954 VDD.n2401 VDD.n2400 0.152939
R8955 VDD.n2402 VDD.n2401 0.152939
R8956 VDD.n2402 VDD.n2191 0.152939
R8957 VDD.n2416 VDD.n2191 0.152939
R8958 VDD.n2417 VDD.n2416 0.152939
R8959 VDD.n2418 VDD.n2417 0.152939
R8960 VDD.n2418 VDD.n2179 0.152939
R8961 VDD.n2432 VDD.n2179 0.152939
R8962 VDD.n2433 VDD.n2432 0.152939
R8963 VDD.n2434 VDD.n2433 0.152939
R8964 VDD.n2434 VDD.n2167 0.152939
R8965 VDD.n2448 VDD.n2167 0.152939
R8966 VDD.n2449 VDD.n2448 0.152939
R8967 VDD.n2450 VDD.n2449 0.152939
R8968 VDD.n2450 VDD.n2155 0.152939
R8969 VDD.n2464 VDD.n2155 0.152939
R8970 VDD.n2465 VDD.n2464 0.152939
R8971 VDD.n2466 VDD.n2465 0.152939
R8972 VDD.n2466 VDD.n2143 0.152939
R8973 VDD.n2480 VDD.n2143 0.152939
R8974 VDD.n2481 VDD.n2480 0.152939
R8975 VDD.n2482 VDD.n2481 0.152939
R8976 VDD.n2482 VDD.n2131 0.152939
R8977 VDD.n2496 VDD.n2131 0.152939
R8978 VDD.n2497 VDD.n2496 0.152939
R8979 VDD.n2498 VDD.n2497 0.152939
R8980 VDD.n2498 VDD.n2119 0.152939
R8981 VDD.n2512 VDD.n2119 0.152939
R8982 VDD.n2513 VDD.n2512 0.152939
R8983 VDD.n2514 VDD.n2513 0.152939
R8984 VDD.n2514 VDD.n2107 0.152939
R8985 VDD.n2528 VDD.n2107 0.152939
R8986 VDD.n2529 VDD.n2528 0.152939
R8987 VDD.n2530 VDD.n2529 0.152939
R8988 VDD.n2530 VDD.n2095 0.152939
R8989 VDD.n2544 VDD.n2095 0.152939
R8990 VDD.n2545 VDD.n2544 0.152939
R8991 VDD.n2546 VDD.n2545 0.152939
R8992 VDD.n2546 VDD.n2083 0.152939
R8993 VDD.n2560 VDD.n2083 0.152939
R8994 VDD.n2561 VDD.n2560 0.152939
R8995 VDD.n2562 VDD.n2561 0.152939
R8996 VDD.n2562 VDD.n2071 0.152939
R8997 VDD.n2576 VDD.n2071 0.152939
R8998 VDD.n2577 VDD.n2576 0.152939
R8999 VDD.n2578 VDD.n2577 0.152939
R9000 VDD.n2578 VDD.n2059 0.152939
R9001 VDD.n2592 VDD.n2059 0.152939
R9002 VDD.n2593 VDD.n2592 0.152939
R9003 VDD.n2595 VDD.n2593 0.152939
R9004 VDD.n2595 VDD.n2594 0.152939
R9005 VDD.n544 VDD.n542 0.0797683
R9006 VDD.n4238 VDD.n675 0.0797683
R9007 VDD.n4712 VDD.n4711 0.0695946
R9008 VDD.n4712 VDD.n36 0.0695946
R9009 VDD.n2609 VDD.n2047 0.0695946
R9010 VDD.n2594 VDD.n2047 0.0695946
R9011 VDD VDD.n15 0.00833333
R9012 VDD.n2940 VDD.n1595 0.0070625
R9013 VDD.n2829 VDD.n1804 0.0070625
R9014 VDD.n4247 VDD.n542 0.00675
R9015 VDD.n4239 VDD.n4238 0.00675
R9016 GND.n10385 GND.n10384 2287.73
R9017 GND.n8931 GND.n8930 1248.19
R9018 GND.n9051 GND.n1462 780.793
R9019 GND.n10386 GND.n662 780.793
R9020 GND.n10533 GND.n573 780.793
R9021 GND.n8929 GND.n1577 780.793
R9022 GND.n5816 GND.n4367 775.989
R9023 GND.n5868 GND.n4369 775.989
R9024 GND.n8007 GND.n8006 775.989
R9025 GND.n8054 GND.n3864 775.989
R9026 GND.n10913 GND.n444 751.963
R9027 GND.n10782 GND.n446 751.963
R9028 GND.n7533 GND.n5877 751.963
R9029 GND.n7645 GND.n4605 751.963
R9030 GND.n8309 GND.n2126 751.963
R9031 GND.n8481 GND.n2124 751.963
R9032 GND.n1803 GND.n1802 751.963
R9033 GND.n8814 GND.n1728 751.963
R9034 GND.n10911 GND.n449 737.549
R9035 GND.n10898 GND.n447 737.549
R9036 GND.n5883 GND.n5880 737.549
R9037 GND.n7531 GND.n5916 737.549
R9038 GND.n8700 GND.n8699 737.549
R9039 GND.n8479 GND.n8478 737.549
R9040 GND.n2948 GND.n1804 737.549
R9041 GND.n2146 GND.n2127 737.549
R9042 GND.n9052 GND.n1461 644.729
R9043 GND.n5916 GND.n5915 589.749
R9044 GND.n8478 GND.n8477 589.749
R9045 GND.n2146 GND.n2145 588.543
R9046 GND.n5884 GND.n5883 588.543
R9047 GND.n9047 GND.n1462 585
R9048 GND.n1462 GND.n1461 585
R9049 GND.n9046 GND.n9045 585
R9050 GND.n9045 GND.n9044 585
R9051 GND.n1465 GND.n1464 585
R9052 GND.n9043 GND.n1465 585
R9053 GND.n9041 GND.n9040 585
R9054 GND.n9042 GND.n9041 585
R9055 GND.n9039 GND.n1467 585
R9056 GND.n1467 GND.n1466 585
R9057 GND.n9038 GND.n9037 585
R9058 GND.n9037 GND.n9036 585
R9059 GND.n1473 GND.n1472 585
R9060 GND.n9035 GND.n1473 585
R9061 GND.n9033 GND.n9032 585
R9062 GND.n9034 GND.n9033 585
R9063 GND.n9031 GND.n1475 585
R9064 GND.n1475 GND.n1474 585
R9065 GND.n9030 GND.n9029 585
R9066 GND.n9029 GND.n9028 585
R9067 GND.n1481 GND.n1480 585
R9068 GND.n9027 GND.n1481 585
R9069 GND.n9025 GND.n9024 585
R9070 GND.n9026 GND.n9025 585
R9071 GND.n9023 GND.n1483 585
R9072 GND.n1483 GND.n1482 585
R9073 GND.n9022 GND.n9021 585
R9074 GND.n9021 GND.n9020 585
R9075 GND.n1489 GND.n1488 585
R9076 GND.n9019 GND.n1489 585
R9077 GND.n9017 GND.n9016 585
R9078 GND.n9018 GND.n9017 585
R9079 GND.n9015 GND.n1491 585
R9080 GND.n1491 GND.n1490 585
R9081 GND.n9014 GND.n9013 585
R9082 GND.n9013 GND.n9012 585
R9083 GND.n1497 GND.n1496 585
R9084 GND.n9011 GND.n1497 585
R9085 GND.n9009 GND.n9008 585
R9086 GND.n9010 GND.n9009 585
R9087 GND.n9007 GND.n1499 585
R9088 GND.n1499 GND.n1498 585
R9089 GND.n9006 GND.n9005 585
R9090 GND.n9005 GND.n9004 585
R9091 GND.n1505 GND.n1504 585
R9092 GND.n9003 GND.n1505 585
R9093 GND.n9001 GND.n9000 585
R9094 GND.n9002 GND.n9001 585
R9095 GND.n8999 GND.n1507 585
R9096 GND.n1507 GND.n1506 585
R9097 GND.n8998 GND.n8997 585
R9098 GND.n8997 GND.n8996 585
R9099 GND.n1513 GND.n1512 585
R9100 GND.n8995 GND.n1513 585
R9101 GND.n8993 GND.n8992 585
R9102 GND.n8994 GND.n8993 585
R9103 GND.n8991 GND.n1515 585
R9104 GND.n1515 GND.n1514 585
R9105 GND.n8990 GND.n8989 585
R9106 GND.n8989 GND.n8988 585
R9107 GND.n1521 GND.n1520 585
R9108 GND.n8987 GND.n1521 585
R9109 GND.n8985 GND.n8984 585
R9110 GND.n8986 GND.n8985 585
R9111 GND.n8983 GND.n1523 585
R9112 GND.n1523 GND.n1522 585
R9113 GND.n8982 GND.n8981 585
R9114 GND.n8981 GND.n8980 585
R9115 GND.n1529 GND.n1528 585
R9116 GND.n8979 GND.n1529 585
R9117 GND.n8977 GND.n8976 585
R9118 GND.n8978 GND.n8977 585
R9119 GND.n8975 GND.n1531 585
R9120 GND.n1531 GND.n1530 585
R9121 GND.n8974 GND.n8973 585
R9122 GND.n8973 GND.n8972 585
R9123 GND.n1537 GND.n1536 585
R9124 GND.n8971 GND.n1537 585
R9125 GND.n8969 GND.n8968 585
R9126 GND.n8970 GND.n8969 585
R9127 GND.n8967 GND.n1539 585
R9128 GND.n1539 GND.n1538 585
R9129 GND.n8966 GND.n8965 585
R9130 GND.n8965 GND.n8964 585
R9131 GND.n1545 GND.n1544 585
R9132 GND.n8963 GND.n1545 585
R9133 GND.n8961 GND.n8960 585
R9134 GND.n8962 GND.n8961 585
R9135 GND.n8959 GND.n1547 585
R9136 GND.n1547 GND.n1546 585
R9137 GND.n8958 GND.n8957 585
R9138 GND.n8957 GND.n8956 585
R9139 GND.n1553 GND.n1552 585
R9140 GND.n8955 GND.n1553 585
R9141 GND.n8953 GND.n8952 585
R9142 GND.n8954 GND.n8953 585
R9143 GND.n8951 GND.n1555 585
R9144 GND.n1555 GND.n1554 585
R9145 GND.n8950 GND.n8949 585
R9146 GND.n8949 GND.n8948 585
R9147 GND.n1561 GND.n1560 585
R9148 GND.n8947 GND.n1561 585
R9149 GND.n8945 GND.n8944 585
R9150 GND.n8946 GND.n8945 585
R9151 GND.n8943 GND.n1563 585
R9152 GND.n1563 GND.n1562 585
R9153 GND.n8942 GND.n8941 585
R9154 GND.n8941 GND.n8940 585
R9155 GND.n1569 GND.n1568 585
R9156 GND.n8939 GND.n1569 585
R9157 GND.n8937 GND.n8936 585
R9158 GND.n8938 GND.n8937 585
R9159 GND.n8935 GND.n1571 585
R9160 GND.n1571 GND.n1570 585
R9161 GND.n8934 GND.n8933 585
R9162 GND.n8933 GND.n8932 585
R9163 GND.n1577 GND.n1576 585
R9164 GND.n8931 GND.n1577 585
R9165 GND.n9051 GND.n9050 585
R9166 GND.n9052 GND.n9051 585
R9167 GND.n1460 GND.n1459 585
R9168 GND.n9053 GND.n1460 585
R9169 GND.n9056 GND.n9055 585
R9170 GND.n9055 GND.n9054 585
R9171 GND.n1457 GND.n1456 585
R9172 GND.n1456 GND.n1455 585
R9173 GND.n9061 GND.n9060 585
R9174 GND.n9062 GND.n9061 585
R9175 GND.n1454 GND.n1453 585
R9176 GND.n9063 GND.n1454 585
R9177 GND.n9066 GND.n9065 585
R9178 GND.n9065 GND.n9064 585
R9179 GND.n1451 GND.n1450 585
R9180 GND.n1450 GND.n1449 585
R9181 GND.n9071 GND.n9070 585
R9182 GND.n9072 GND.n9071 585
R9183 GND.n1448 GND.n1447 585
R9184 GND.n9073 GND.n1448 585
R9185 GND.n9076 GND.n9075 585
R9186 GND.n9075 GND.n9074 585
R9187 GND.n1445 GND.n1444 585
R9188 GND.n1444 GND.n1443 585
R9189 GND.n9081 GND.n9080 585
R9190 GND.n9082 GND.n9081 585
R9191 GND.n1442 GND.n1441 585
R9192 GND.n9083 GND.n1442 585
R9193 GND.n9086 GND.n9085 585
R9194 GND.n9085 GND.n9084 585
R9195 GND.n1439 GND.n1438 585
R9196 GND.n1438 GND.n1437 585
R9197 GND.n9091 GND.n9090 585
R9198 GND.n9092 GND.n9091 585
R9199 GND.n1436 GND.n1435 585
R9200 GND.n9093 GND.n1436 585
R9201 GND.n9096 GND.n9095 585
R9202 GND.n9095 GND.n9094 585
R9203 GND.n1433 GND.n1432 585
R9204 GND.n1432 GND.n1431 585
R9205 GND.n9101 GND.n9100 585
R9206 GND.n9102 GND.n9101 585
R9207 GND.n1430 GND.n1429 585
R9208 GND.n9103 GND.n1430 585
R9209 GND.n9106 GND.n9105 585
R9210 GND.n9105 GND.n9104 585
R9211 GND.n1427 GND.n1426 585
R9212 GND.n1426 GND.n1425 585
R9213 GND.n9111 GND.n9110 585
R9214 GND.n9112 GND.n9111 585
R9215 GND.n1424 GND.n1423 585
R9216 GND.n9113 GND.n1424 585
R9217 GND.n9116 GND.n9115 585
R9218 GND.n9115 GND.n9114 585
R9219 GND.n1421 GND.n1420 585
R9220 GND.n1420 GND.n1419 585
R9221 GND.n9121 GND.n9120 585
R9222 GND.n9122 GND.n9121 585
R9223 GND.n1418 GND.n1417 585
R9224 GND.n9123 GND.n1418 585
R9225 GND.n9126 GND.n9125 585
R9226 GND.n9125 GND.n9124 585
R9227 GND.n1415 GND.n1414 585
R9228 GND.n1414 GND.n1413 585
R9229 GND.n9131 GND.n9130 585
R9230 GND.n9132 GND.n9131 585
R9231 GND.n1412 GND.n1411 585
R9232 GND.n9133 GND.n1412 585
R9233 GND.n9136 GND.n9135 585
R9234 GND.n9135 GND.n9134 585
R9235 GND.n1409 GND.n1408 585
R9236 GND.n1408 GND.n1407 585
R9237 GND.n9141 GND.n9140 585
R9238 GND.n9142 GND.n9141 585
R9239 GND.n1406 GND.n1405 585
R9240 GND.n9143 GND.n1406 585
R9241 GND.n9146 GND.n9145 585
R9242 GND.n9145 GND.n9144 585
R9243 GND.n1403 GND.n1402 585
R9244 GND.n1402 GND.n1401 585
R9245 GND.n9151 GND.n9150 585
R9246 GND.n9152 GND.n9151 585
R9247 GND.n1400 GND.n1399 585
R9248 GND.n9153 GND.n1400 585
R9249 GND.n9156 GND.n9155 585
R9250 GND.n9155 GND.n9154 585
R9251 GND.n1397 GND.n1396 585
R9252 GND.n1396 GND.n1395 585
R9253 GND.n9161 GND.n9160 585
R9254 GND.n9162 GND.n9161 585
R9255 GND.n1394 GND.n1393 585
R9256 GND.n9163 GND.n1394 585
R9257 GND.n9166 GND.n9165 585
R9258 GND.n9165 GND.n9164 585
R9259 GND.n1391 GND.n1390 585
R9260 GND.n1390 GND.n1389 585
R9261 GND.n9171 GND.n9170 585
R9262 GND.n9172 GND.n9171 585
R9263 GND.n1388 GND.n1387 585
R9264 GND.n9173 GND.n1388 585
R9265 GND.n9176 GND.n9175 585
R9266 GND.n9175 GND.n9174 585
R9267 GND.n1385 GND.n1384 585
R9268 GND.n1384 GND.n1383 585
R9269 GND.n9181 GND.n9180 585
R9270 GND.n9182 GND.n9181 585
R9271 GND.n1382 GND.n1381 585
R9272 GND.n9183 GND.n1382 585
R9273 GND.n9186 GND.n9185 585
R9274 GND.n9185 GND.n9184 585
R9275 GND.n1379 GND.n1378 585
R9276 GND.n1378 GND.n1377 585
R9277 GND.n9191 GND.n9190 585
R9278 GND.n9192 GND.n9191 585
R9279 GND.n1376 GND.n1375 585
R9280 GND.n9193 GND.n1376 585
R9281 GND.n9196 GND.n9195 585
R9282 GND.n9195 GND.n9194 585
R9283 GND.n1373 GND.n1372 585
R9284 GND.n1372 GND.n1371 585
R9285 GND.n9201 GND.n9200 585
R9286 GND.n9202 GND.n9201 585
R9287 GND.n1370 GND.n1369 585
R9288 GND.n9203 GND.n1370 585
R9289 GND.n9206 GND.n9205 585
R9290 GND.n9205 GND.n9204 585
R9291 GND.n1367 GND.n1366 585
R9292 GND.n1366 GND.n1365 585
R9293 GND.n9211 GND.n9210 585
R9294 GND.n9212 GND.n9211 585
R9295 GND.n1364 GND.n1363 585
R9296 GND.n9213 GND.n1364 585
R9297 GND.n9216 GND.n9215 585
R9298 GND.n9215 GND.n9214 585
R9299 GND.n1361 GND.n1360 585
R9300 GND.n1360 GND.n1359 585
R9301 GND.n9221 GND.n9220 585
R9302 GND.n9222 GND.n9221 585
R9303 GND.n1358 GND.n1357 585
R9304 GND.n9223 GND.n1358 585
R9305 GND.n9226 GND.n9225 585
R9306 GND.n9225 GND.n9224 585
R9307 GND.n1355 GND.n1354 585
R9308 GND.n1354 GND.n1353 585
R9309 GND.n9231 GND.n9230 585
R9310 GND.n9232 GND.n9231 585
R9311 GND.n1352 GND.n1351 585
R9312 GND.n9233 GND.n1352 585
R9313 GND.n9236 GND.n9235 585
R9314 GND.n9235 GND.n9234 585
R9315 GND.n1349 GND.n1348 585
R9316 GND.n1348 GND.n1347 585
R9317 GND.n9241 GND.n9240 585
R9318 GND.n9242 GND.n9241 585
R9319 GND.n1346 GND.n1345 585
R9320 GND.n9243 GND.n1346 585
R9321 GND.n9246 GND.n9245 585
R9322 GND.n9245 GND.n9244 585
R9323 GND.n1343 GND.n1342 585
R9324 GND.n1342 GND.n1341 585
R9325 GND.n9251 GND.n9250 585
R9326 GND.n9252 GND.n9251 585
R9327 GND.n1340 GND.n1339 585
R9328 GND.n9253 GND.n1340 585
R9329 GND.n9256 GND.n9255 585
R9330 GND.n9255 GND.n9254 585
R9331 GND.n1337 GND.n1336 585
R9332 GND.n1336 GND.n1335 585
R9333 GND.n9261 GND.n9260 585
R9334 GND.n9262 GND.n9261 585
R9335 GND.n1334 GND.n1333 585
R9336 GND.n9263 GND.n1334 585
R9337 GND.n9266 GND.n9265 585
R9338 GND.n9265 GND.n9264 585
R9339 GND.n1331 GND.n1330 585
R9340 GND.n1330 GND.n1329 585
R9341 GND.n9271 GND.n9270 585
R9342 GND.n9272 GND.n9271 585
R9343 GND.n1328 GND.n1327 585
R9344 GND.n9273 GND.n1328 585
R9345 GND.n9276 GND.n9275 585
R9346 GND.n9275 GND.n9274 585
R9347 GND.n1325 GND.n1324 585
R9348 GND.n1324 GND.n1323 585
R9349 GND.n9281 GND.n9280 585
R9350 GND.n9282 GND.n9281 585
R9351 GND.n1322 GND.n1321 585
R9352 GND.n9283 GND.n1322 585
R9353 GND.n9286 GND.n9285 585
R9354 GND.n9285 GND.n9284 585
R9355 GND.n1319 GND.n1318 585
R9356 GND.n1318 GND.n1317 585
R9357 GND.n9291 GND.n9290 585
R9358 GND.n9292 GND.n9291 585
R9359 GND.n1316 GND.n1315 585
R9360 GND.n9293 GND.n1316 585
R9361 GND.n9296 GND.n9295 585
R9362 GND.n9295 GND.n9294 585
R9363 GND.n1313 GND.n1312 585
R9364 GND.n1312 GND.n1311 585
R9365 GND.n9301 GND.n9300 585
R9366 GND.n9302 GND.n9301 585
R9367 GND.n1310 GND.n1309 585
R9368 GND.n9303 GND.n1310 585
R9369 GND.n9306 GND.n9305 585
R9370 GND.n9305 GND.n9304 585
R9371 GND.n1307 GND.n1306 585
R9372 GND.n1306 GND.n1305 585
R9373 GND.n9311 GND.n9310 585
R9374 GND.n9312 GND.n9311 585
R9375 GND.n1304 GND.n1303 585
R9376 GND.n9313 GND.n1304 585
R9377 GND.n9316 GND.n9315 585
R9378 GND.n9315 GND.n9314 585
R9379 GND.n1301 GND.n1300 585
R9380 GND.n1300 GND.n1299 585
R9381 GND.n9321 GND.n9320 585
R9382 GND.n9322 GND.n9321 585
R9383 GND.n1298 GND.n1297 585
R9384 GND.n9323 GND.n1298 585
R9385 GND.n9326 GND.n9325 585
R9386 GND.n9325 GND.n9324 585
R9387 GND.n1295 GND.n1294 585
R9388 GND.n1294 GND.n1293 585
R9389 GND.n9331 GND.n9330 585
R9390 GND.n9332 GND.n9331 585
R9391 GND.n1292 GND.n1291 585
R9392 GND.n9333 GND.n1292 585
R9393 GND.n9336 GND.n9335 585
R9394 GND.n9335 GND.n9334 585
R9395 GND.n1289 GND.n1288 585
R9396 GND.n1288 GND.n1287 585
R9397 GND.n9341 GND.n9340 585
R9398 GND.n9342 GND.n9341 585
R9399 GND.n1286 GND.n1285 585
R9400 GND.n9343 GND.n1286 585
R9401 GND.n9346 GND.n9345 585
R9402 GND.n9345 GND.n9344 585
R9403 GND.n1283 GND.n1282 585
R9404 GND.n1282 GND.n1281 585
R9405 GND.n9351 GND.n9350 585
R9406 GND.n9352 GND.n9351 585
R9407 GND.n1280 GND.n1279 585
R9408 GND.n9353 GND.n1280 585
R9409 GND.n9356 GND.n9355 585
R9410 GND.n9355 GND.n9354 585
R9411 GND.n1277 GND.n1276 585
R9412 GND.n1276 GND.n1275 585
R9413 GND.n9361 GND.n9360 585
R9414 GND.n9362 GND.n9361 585
R9415 GND.n1274 GND.n1273 585
R9416 GND.n9363 GND.n1274 585
R9417 GND.n9366 GND.n9365 585
R9418 GND.n9365 GND.n9364 585
R9419 GND.n1271 GND.n1270 585
R9420 GND.n1270 GND.n1269 585
R9421 GND.n9371 GND.n9370 585
R9422 GND.n9372 GND.n9371 585
R9423 GND.n1268 GND.n1267 585
R9424 GND.n9373 GND.n1268 585
R9425 GND.n9376 GND.n9375 585
R9426 GND.n9375 GND.n9374 585
R9427 GND.n1265 GND.n1264 585
R9428 GND.n1264 GND.n1263 585
R9429 GND.n9381 GND.n9380 585
R9430 GND.n9382 GND.n9381 585
R9431 GND.n1262 GND.n1261 585
R9432 GND.n9383 GND.n1262 585
R9433 GND.n9386 GND.n9385 585
R9434 GND.n9385 GND.n9384 585
R9435 GND.n1259 GND.n1258 585
R9436 GND.n1258 GND.n1257 585
R9437 GND.n9391 GND.n9390 585
R9438 GND.n9392 GND.n9391 585
R9439 GND.n1256 GND.n1255 585
R9440 GND.n9393 GND.n1256 585
R9441 GND.n9396 GND.n9395 585
R9442 GND.n9395 GND.n9394 585
R9443 GND.n1253 GND.n1252 585
R9444 GND.n1252 GND.n1251 585
R9445 GND.n9401 GND.n9400 585
R9446 GND.n9402 GND.n9401 585
R9447 GND.n1250 GND.n1249 585
R9448 GND.n9403 GND.n1250 585
R9449 GND.n9406 GND.n9405 585
R9450 GND.n9405 GND.n9404 585
R9451 GND.n1247 GND.n1246 585
R9452 GND.n1246 GND.n1245 585
R9453 GND.n9411 GND.n9410 585
R9454 GND.n9412 GND.n9411 585
R9455 GND.n1244 GND.n1243 585
R9456 GND.n9413 GND.n1244 585
R9457 GND.n9416 GND.n9415 585
R9458 GND.n9415 GND.n9414 585
R9459 GND.n1241 GND.n1240 585
R9460 GND.n1240 GND.n1239 585
R9461 GND.n9421 GND.n9420 585
R9462 GND.n9422 GND.n9421 585
R9463 GND.n1238 GND.n1237 585
R9464 GND.n9423 GND.n1238 585
R9465 GND.n9426 GND.n9425 585
R9466 GND.n9425 GND.n9424 585
R9467 GND.n1235 GND.n1234 585
R9468 GND.n1234 GND.n1233 585
R9469 GND.n9431 GND.n9430 585
R9470 GND.n9432 GND.n9431 585
R9471 GND.n1232 GND.n1231 585
R9472 GND.n9433 GND.n1232 585
R9473 GND.n9436 GND.n9435 585
R9474 GND.n9435 GND.n9434 585
R9475 GND.n1229 GND.n1228 585
R9476 GND.n1228 GND.n1227 585
R9477 GND.n9441 GND.n9440 585
R9478 GND.n9442 GND.n9441 585
R9479 GND.n1226 GND.n1225 585
R9480 GND.n9443 GND.n1226 585
R9481 GND.n9446 GND.n9445 585
R9482 GND.n9445 GND.n9444 585
R9483 GND.n1223 GND.n1222 585
R9484 GND.n1222 GND.n1221 585
R9485 GND.n9451 GND.n9450 585
R9486 GND.n9452 GND.n9451 585
R9487 GND.n1220 GND.n1219 585
R9488 GND.n9453 GND.n1220 585
R9489 GND.n9456 GND.n9455 585
R9490 GND.n9455 GND.n9454 585
R9491 GND.n1217 GND.n1216 585
R9492 GND.n1216 GND.n1215 585
R9493 GND.n9461 GND.n9460 585
R9494 GND.n9462 GND.n9461 585
R9495 GND.n1214 GND.n1213 585
R9496 GND.n9463 GND.n1214 585
R9497 GND.n9466 GND.n9465 585
R9498 GND.n9465 GND.n9464 585
R9499 GND.n1211 GND.n1210 585
R9500 GND.n1210 GND.n1209 585
R9501 GND.n9471 GND.n9470 585
R9502 GND.n9472 GND.n9471 585
R9503 GND.n1208 GND.n1207 585
R9504 GND.n9473 GND.n1208 585
R9505 GND.n9476 GND.n9475 585
R9506 GND.n9475 GND.n9474 585
R9507 GND.n1205 GND.n1204 585
R9508 GND.n1204 GND.n1203 585
R9509 GND.n9481 GND.n9480 585
R9510 GND.n9482 GND.n9481 585
R9511 GND.n1202 GND.n1201 585
R9512 GND.n9483 GND.n1202 585
R9513 GND.n9486 GND.n9485 585
R9514 GND.n9485 GND.n9484 585
R9515 GND.n1199 GND.n1198 585
R9516 GND.n1198 GND.n1197 585
R9517 GND.n9491 GND.n9490 585
R9518 GND.n9492 GND.n9491 585
R9519 GND.n1196 GND.n1195 585
R9520 GND.n9493 GND.n1196 585
R9521 GND.n9496 GND.n9495 585
R9522 GND.n9495 GND.n9494 585
R9523 GND.n1193 GND.n1192 585
R9524 GND.n1192 GND.n1191 585
R9525 GND.n9501 GND.n9500 585
R9526 GND.n9502 GND.n9501 585
R9527 GND.n1190 GND.n1189 585
R9528 GND.n9503 GND.n1190 585
R9529 GND.n9506 GND.n9505 585
R9530 GND.n9505 GND.n9504 585
R9531 GND.n1187 GND.n1186 585
R9532 GND.n1186 GND.n1185 585
R9533 GND.n9511 GND.n9510 585
R9534 GND.n9512 GND.n9511 585
R9535 GND.n1184 GND.n1183 585
R9536 GND.n9513 GND.n1184 585
R9537 GND.n9516 GND.n9515 585
R9538 GND.n9515 GND.n9514 585
R9539 GND.n1181 GND.n1180 585
R9540 GND.n1180 GND.n1179 585
R9541 GND.n9521 GND.n9520 585
R9542 GND.n9522 GND.n9521 585
R9543 GND.n1178 GND.n1177 585
R9544 GND.n9523 GND.n1178 585
R9545 GND.n9526 GND.n9525 585
R9546 GND.n9525 GND.n9524 585
R9547 GND.n1175 GND.n1174 585
R9548 GND.n1174 GND.n1173 585
R9549 GND.n9531 GND.n9530 585
R9550 GND.n9532 GND.n9531 585
R9551 GND.n1172 GND.n1171 585
R9552 GND.n9533 GND.n1172 585
R9553 GND.n9536 GND.n9535 585
R9554 GND.n9535 GND.n9534 585
R9555 GND.n1169 GND.n1168 585
R9556 GND.n1168 GND.n1167 585
R9557 GND.n9541 GND.n9540 585
R9558 GND.n9542 GND.n9541 585
R9559 GND.n1166 GND.n1165 585
R9560 GND.n9543 GND.n1166 585
R9561 GND.n9546 GND.n9545 585
R9562 GND.n9545 GND.n9544 585
R9563 GND.n1163 GND.n1162 585
R9564 GND.n1162 GND.n1161 585
R9565 GND.n9551 GND.n9550 585
R9566 GND.n9552 GND.n9551 585
R9567 GND.n1160 GND.n1159 585
R9568 GND.n9553 GND.n1160 585
R9569 GND.n9556 GND.n9555 585
R9570 GND.n9555 GND.n9554 585
R9571 GND.n1157 GND.n1156 585
R9572 GND.n1156 GND.n1155 585
R9573 GND.n9561 GND.n9560 585
R9574 GND.n9562 GND.n9561 585
R9575 GND.n1154 GND.n1153 585
R9576 GND.n9563 GND.n1154 585
R9577 GND.n9566 GND.n9565 585
R9578 GND.n9565 GND.n9564 585
R9579 GND.n1151 GND.n1150 585
R9580 GND.n1150 GND.n1149 585
R9581 GND.n9571 GND.n9570 585
R9582 GND.n9572 GND.n9571 585
R9583 GND.n1148 GND.n1147 585
R9584 GND.n9573 GND.n1148 585
R9585 GND.n9576 GND.n9575 585
R9586 GND.n9575 GND.n9574 585
R9587 GND.n1145 GND.n1144 585
R9588 GND.n1144 GND.n1143 585
R9589 GND.n9581 GND.n9580 585
R9590 GND.n9582 GND.n9581 585
R9591 GND.n1142 GND.n1141 585
R9592 GND.n9583 GND.n1142 585
R9593 GND.n9586 GND.n9585 585
R9594 GND.n9585 GND.n9584 585
R9595 GND.n1139 GND.n1138 585
R9596 GND.n1138 GND.n1137 585
R9597 GND.n9591 GND.n9590 585
R9598 GND.n9592 GND.n9591 585
R9599 GND.n1136 GND.n1135 585
R9600 GND.n9593 GND.n1136 585
R9601 GND.n9596 GND.n9595 585
R9602 GND.n9595 GND.n9594 585
R9603 GND.n1133 GND.n1132 585
R9604 GND.n1132 GND.n1131 585
R9605 GND.n9601 GND.n9600 585
R9606 GND.n9602 GND.n9601 585
R9607 GND.n1130 GND.n1129 585
R9608 GND.n9603 GND.n1130 585
R9609 GND.n9606 GND.n9605 585
R9610 GND.n9605 GND.n9604 585
R9611 GND.n1127 GND.n1126 585
R9612 GND.n1126 GND.n1125 585
R9613 GND.n9611 GND.n9610 585
R9614 GND.n9612 GND.n9611 585
R9615 GND.n1124 GND.n1123 585
R9616 GND.n9613 GND.n1124 585
R9617 GND.n9616 GND.n9615 585
R9618 GND.n9615 GND.n9614 585
R9619 GND.n1121 GND.n1120 585
R9620 GND.n1120 GND.n1119 585
R9621 GND.n9621 GND.n9620 585
R9622 GND.n9622 GND.n9621 585
R9623 GND.n1118 GND.n1117 585
R9624 GND.n9623 GND.n1118 585
R9625 GND.n9626 GND.n9625 585
R9626 GND.n9625 GND.n9624 585
R9627 GND.n1115 GND.n1114 585
R9628 GND.n1114 GND.n1113 585
R9629 GND.n9631 GND.n9630 585
R9630 GND.n9632 GND.n9631 585
R9631 GND.n1112 GND.n1111 585
R9632 GND.n9633 GND.n1112 585
R9633 GND.n9636 GND.n9635 585
R9634 GND.n9635 GND.n9634 585
R9635 GND.n1109 GND.n1108 585
R9636 GND.n1108 GND.n1107 585
R9637 GND.n9641 GND.n9640 585
R9638 GND.n9642 GND.n9641 585
R9639 GND.n1106 GND.n1105 585
R9640 GND.n9643 GND.n1106 585
R9641 GND.n9646 GND.n9645 585
R9642 GND.n9645 GND.n9644 585
R9643 GND.n1103 GND.n1102 585
R9644 GND.n1102 GND.n1101 585
R9645 GND.n9651 GND.n9650 585
R9646 GND.n9652 GND.n9651 585
R9647 GND.n1100 GND.n1099 585
R9648 GND.n9653 GND.n1100 585
R9649 GND.n9656 GND.n9655 585
R9650 GND.n9655 GND.n9654 585
R9651 GND.n1097 GND.n1096 585
R9652 GND.n1096 GND.n1095 585
R9653 GND.n9661 GND.n9660 585
R9654 GND.n9662 GND.n9661 585
R9655 GND.n1094 GND.n1093 585
R9656 GND.n9663 GND.n1094 585
R9657 GND.n9666 GND.n9665 585
R9658 GND.n9665 GND.n9664 585
R9659 GND.n1091 GND.n1090 585
R9660 GND.n1090 GND.n1089 585
R9661 GND.n9671 GND.n9670 585
R9662 GND.n9672 GND.n9671 585
R9663 GND.n1088 GND.n1087 585
R9664 GND.n9673 GND.n1088 585
R9665 GND.n9676 GND.n9675 585
R9666 GND.n9675 GND.n9674 585
R9667 GND.n1085 GND.n1084 585
R9668 GND.n1084 GND.n1083 585
R9669 GND.n9681 GND.n9680 585
R9670 GND.n9682 GND.n9681 585
R9671 GND.n1082 GND.n1081 585
R9672 GND.n9683 GND.n1082 585
R9673 GND.n9686 GND.n9685 585
R9674 GND.n9685 GND.n9684 585
R9675 GND.n1079 GND.n1078 585
R9676 GND.n1078 GND.n1077 585
R9677 GND.n9691 GND.n9690 585
R9678 GND.n9692 GND.n9691 585
R9679 GND.n1076 GND.n1075 585
R9680 GND.n9693 GND.n1076 585
R9681 GND.n9696 GND.n9695 585
R9682 GND.n9695 GND.n9694 585
R9683 GND.n1073 GND.n1072 585
R9684 GND.n1072 GND.n1071 585
R9685 GND.n9701 GND.n9700 585
R9686 GND.n9702 GND.n9701 585
R9687 GND.n1070 GND.n1069 585
R9688 GND.n9703 GND.n1070 585
R9689 GND.n9706 GND.n9705 585
R9690 GND.n9705 GND.n9704 585
R9691 GND.n1067 GND.n1066 585
R9692 GND.n1066 GND.n1065 585
R9693 GND.n9711 GND.n9710 585
R9694 GND.n9712 GND.n9711 585
R9695 GND.n1064 GND.n1063 585
R9696 GND.n9713 GND.n1064 585
R9697 GND.n9716 GND.n9715 585
R9698 GND.n9715 GND.n9714 585
R9699 GND.n1061 GND.n1060 585
R9700 GND.n1060 GND.n1059 585
R9701 GND.n9721 GND.n9720 585
R9702 GND.n9722 GND.n9721 585
R9703 GND.n1058 GND.n1057 585
R9704 GND.n9723 GND.n1058 585
R9705 GND.n9726 GND.n9725 585
R9706 GND.n9725 GND.n9724 585
R9707 GND.n1055 GND.n1054 585
R9708 GND.n1054 GND.n1053 585
R9709 GND.n9731 GND.n9730 585
R9710 GND.n9732 GND.n9731 585
R9711 GND.n1052 GND.n1051 585
R9712 GND.n9733 GND.n1052 585
R9713 GND.n9736 GND.n9735 585
R9714 GND.n9735 GND.n9734 585
R9715 GND.n1049 GND.n1048 585
R9716 GND.n1048 GND.n1047 585
R9717 GND.n9741 GND.n9740 585
R9718 GND.n9742 GND.n9741 585
R9719 GND.n1046 GND.n1045 585
R9720 GND.n9743 GND.n1046 585
R9721 GND.n9746 GND.n9745 585
R9722 GND.n9745 GND.n9744 585
R9723 GND.n1043 GND.n1042 585
R9724 GND.n1042 GND.n1041 585
R9725 GND.n9751 GND.n9750 585
R9726 GND.n9752 GND.n9751 585
R9727 GND.n1040 GND.n1039 585
R9728 GND.n9753 GND.n1040 585
R9729 GND.n9756 GND.n9755 585
R9730 GND.n9755 GND.n9754 585
R9731 GND.n1037 GND.n1036 585
R9732 GND.n1036 GND.n1035 585
R9733 GND.n9761 GND.n9760 585
R9734 GND.n9762 GND.n9761 585
R9735 GND.n1034 GND.n1033 585
R9736 GND.n9763 GND.n1034 585
R9737 GND.n9766 GND.n9765 585
R9738 GND.n9765 GND.n9764 585
R9739 GND.n1031 GND.n1030 585
R9740 GND.n1030 GND.n1029 585
R9741 GND.n9771 GND.n9770 585
R9742 GND.n9772 GND.n9771 585
R9743 GND.n1028 GND.n1027 585
R9744 GND.n9773 GND.n1028 585
R9745 GND.n9776 GND.n9775 585
R9746 GND.n9775 GND.n9774 585
R9747 GND.n1025 GND.n1024 585
R9748 GND.n1024 GND.n1023 585
R9749 GND.n9781 GND.n9780 585
R9750 GND.n9782 GND.n9781 585
R9751 GND.n1022 GND.n1021 585
R9752 GND.n9783 GND.n1022 585
R9753 GND.n9786 GND.n9785 585
R9754 GND.n9785 GND.n9784 585
R9755 GND.n1019 GND.n1018 585
R9756 GND.n1018 GND.n1017 585
R9757 GND.n9791 GND.n9790 585
R9758 GND.n9792 GND.n9791 585
R9759 GND.n1016 GND.n1015 585
R9760 GND.n9793 GND.n1016 585
R9761 GND.n9796 GND.n9795 585
R9762 GND.n9795 GND.n9794 585
R9763 GND.n1013 GND.n1012 585
R9764 GND.n1012 GND.n1011 585
R9765 GND.n9801 GND.n9800 585
R9766 GND.n9802 GND.n9801 585
R9767 GND.n1010 GND.n1009 585
R9768 GND.n9803 GND.n1010 585
R9769 GND.n9806 GND.n9805 585
R9770 GND.n9805 GND.n9804 585
R9771 GND.n1007 GND.n1006 585
R9772 GND.n1006 GND.n1005 585
R9773 GND.n9811 GND.n9810 585
R9774 GND.n9812 GND.n9811 585
R9775 GND.n1004 GND.n1003 585
R9776 GND.n9813 GND.n1004 585
R9777 GND.n9816 GND.n9815 585
R9778 GND.n9815 GND.n9814 585
R9779 GND.n1001 GND.n1000 585
R9780 GND.n1000 GND.n999 585
R9781 GND.n9821 GND.n9820 585
R9782 GND.n9822 GND.n9821 585
R9783 GND.n998 GND.n997 585
R9784 GND.n9823 GND.n998 585
R9785 GND.n9826 GND.n9825 585
R9786 GND.n9825 GND.n9824 585
R9787 GND.n995 GND.n994 585
R9788 GND.n994 GND.n993 585
R9789 GND.n9831 GND.n9830 585
R9790 GND.n9832 GND.n9831 585
R9791 GND.n992 GND.n991 585
R9792 GND.n9833 GND.n992 585
R9793 GND.n9836 GND.n9835 585
R9794 GND.n9835 GND.n9834 585
R9795 GND.n989 GND.n988 585
R9796 GND.n988 GND.n987 585
R9797 GND.n9841 GND.n9840 585
R9798 GND.n9842 GND.n9841 585
R9799 GND.n986 GND.n985 585
R9800 GND.n9843 GND.n986 585
R9801 GND.n9846 GND.n9845 585
R9802 GND.n9845 GND.n9844 585
R9803 GND.n983 GND.n982 585
R9804 GND.n982 GND.n981 585
R9805 GND.n9851 GND.n9850 585
R9806 GND.n9852 GND.n9851 585
R9807 GND.n980 GND.n979 585
R9808 GND.n9853 GND.n980 585
R9809 GND.n9856 GND.n9855 585
R9810 GND.n9855 GND.n9854 585
R9811 GND.n977 GND.n976 585
R9812 GND.n976 GND.n975 585
R9813 GND.n9861 GND.n9860 585
R9814 GND.n9862 GND.n9861 585
R9815 GND.n974 GND.n973 585
R9816 GND.n9863 GND.n974 585
R9817 GND.n9866 GND.n9865 585
R9818 GND.n9865 GND.n9864 585
R9819 GND.n971 GND.n970 585
R9820 GND.n970 GND.n969 585
R9821 GND.n9871 GND.n9870 585
R9822 GND.n9872 GND.n9871 585
R9823 GND.n968 GND.n967 585
R9824 GND.n9873 GND.n968 585
R9825 GND.n9876 GND.n9875 585
R9826 GND.n9875 GND.n9874 585
R9827 GND.n965 GND.n964 585
R9828 GND.n964 GND.n963 585
R9829 GND.n9881 GND.n9880 585
R9830 GND.n9882 GND.n9881 585
R9831 GND.n962 GND.n961 585
R9832 GND.n9883 GND.n962 585
R9833 GND.n9886 GND.n9885 585
R9834 GND.n9885 GND.n9884 585
R9835 GND.n959 GND.n958 585
R9836 GND.n958 GND.n957 585
R9837 GND.n9891 GND.n9890 585
R9838 GND.n9892 GND.n9891 585
R9839 GND.n956 GND.n955 585
R9840 GND.n9893 GND.n956 585
R9841 GND.n9896 GND.n9895 585
R9842 GND.n9895 GND.n9894 585
R9843 GND.n953 GND.n952 585
R9844 GND.n952 GND.n951 585
R9845 GND.n9901 GND.n9900 585
R9846 GND.n9902 GND.n9901 585
R9847 GND.n950 GND.n949 585
R9848 GND.n9903 GND.n950 585
R9849 GND.n9906 GND.n9905 585
R9850 GND.n9905 GND.n9904 585
R9851 GND.n947 GND.n946 585
R9852 GND.n946 GND.n945 585
R9853 GND.n9911 GND.n9910 585
R9854 GND.n9912 GND.n9911 585
R9855 GND.n944 GND.n943 585
R9856 GND.n9913 GND.n944 585
R9857 GND.n9916 GND.n9915 585
R9858 GND.n9915 GND.n9914 585
R9859 GND.n941 GND.n940 585
R9860 GND.n940 GND.n939 585
R9861 GND.n9921 GND.n9920 585
R9862 GND.n9922 GND.n9921 585
R9863 GND.n938 GND.n937 585
R9864 GND.n9923 GND.n938 585
R9865 GND.n9926 GND.n9925 585
R9866 GND.n9925 GND.n9924 585
R9867 GND.n935 GND.n934 585
R9868 GND.n934 GND.n933 585
R9869 GND.n9931 GND.n9930 585
R9870 GND.n9932 GND.n9931 585
R9871 GND.n932 GND.n931 585
R9872 GND.n9933 GND.n932 585
R9873 GND.n9936 GND.n9935 585
R9874 GND.n9935 GND.n9934 585
R9875 GND.n929 GND.n928 585
R9876 GND.n928 GND.n927 585
R9877 GND.n9941 GND.n9940 585
R9878 GND.n9942 GND.n9941 585
R9879 GND.n926 GND.n925 585
R9880 GND.n9943 GND.n926 585
R9881 GND.n9946 GND.n9945 585
R9882 GND.n9945 GND.n9944 585
R9883 GND.n923 GND.n922 585
R9884 GND.n922 GND.n921 585
R9885 GND.n9951 GND.n9950 585
R9886 GND.n9952 GND.n9951 585
R9887 GND.n920 GND.n919 585
R9888 GND.n9953 GND.n920 585
R9889 GND.n9956 GND.n9955 585
R9890 GND.n9955 GND.n9954 585
R9891 GND.n917 GND.n916 585
R9892 GND.n916 GND.n915 585
R9893 GND.n9961 GND.n9960 585
R9894 GND.n9962 GND.n9961 585
R9895 GND.n914 GND.n913 585
R9896 GND.n9963 GND.n914 585
R9897 GND.n9966 GND.n9965 585
R9898 GND.n9965 GND.n9964 585
R9899 GND.n911 GND.n910 585
R9900 GND.n910 GND.n909 585
R9901 GND.n9971 GND.n9970 585
R9902 GND.n9972 GND.n9971 585
R9903 GND.n908 GND.n907 585
R9904 GND.n9973 GND.n908 585
R9905 GND.n9976 GND.n9975 585
R9906 GND.n9975 GND.n9974 585
R9907 GND.n905 GND.n904 585
R9908 GND.n904 GND.n903 585
R9909 GND.n9981 GND.n9980 585
R9910 GND.n9982 GND.n9981 585
R9911 GND.n902 GND.n901 585
R9912 GND.n9983 GND.n902 585
R9913 GND.n9986 GND.n9985 585
R9914 GND.n9985 GND.n9984 585
R9915 GND.n899 GND.n898 585
R9916 GND.n898 GND.n897 585
R9917 GND.n9991 GND.n9990 585
R9918 GND.n9992 GND.n9991 585
R9919 GND.n896 GND.n895 585
R9920 GND.n9993 GND.n896 585
R9921 GND.n9996 GND.n9995 585
R9922 GND.n9995 GND.n9994 585
R9923 GND.n893 GND.n892 585
R9924 GND.n892 GND.n891 585
R9925 GND.n10001 GND.n10000 585
R9926 GND.n10002 GND.n10001 585
R9927 GND.n890 GND.n889 585
R9928 GND.n10003 GND.n890 585
R9929 GND.n10006 GND.n10005 585
R9930 GND.n10005 GND.n10004 585
R9931 GND.n887 GND.n886 585
R9932 GND.n886 GND.n885 585
R9933 GND.n10011 GND.n10010 585
R9934 GND.n10012 GND.n10011 585
R9935 GND.n884 GND.n883 585
R9936 GND.n10013 GND.n884 585
R9937 GND.n10016 GND.n10015 585
R9938 GND.n10015 GND.n10014 585
R9939 GND.n881 GND.n880 585
R9940 GND.n880 GND.n879 585
R9941 GND.n10021 GND.n10020 585
R9942 GND.n10022 GND.n10021 585
R9943 GND.n878 GND.n877 585
R9944 GND.n10023 GND.n878 585
R9945 GND.n10026 GND.n10025 585
R9946 GND.n10025 GND.n10024 585
R9947 GND.n875 GND.n874 585
R9948 GND.n874 GND.n873 585
R9949 GND.n10031 GND.n10030 585
R9950 GND.n10032 GND.n10031 585
R9951 GND.n872 GND.n871 585
R9952 GND.n10033 GND.n872 585
R9953 GND.n10036 GND.n10035 585
R9954 GND.n10035 GND.n10034 585
R9955 GND.n869 GND.n868 585
R9956 GND.n868 GND.n867 585
R9957 GND.n10041 GND.n10040 585
R9958 GND.n10042 GND.n10041 585
R9959 GND.n866 GND.n865 585
R9960 GND.n10043 GND.n866 585
R9961 GND.n10046 GND.n10045 585
R9962 GND.n10045 GND.n10044 585
R9963 GND.n863 GND.n862 585
R9964 GND.n862 GND.n861 585
R9965 GND.n10051 GND.n10050 585
R9966 GND.n10052 GND.n10051 585
R9967 GND.n860 GND.n859 585
R9968 GND.n10053 GND.n860 585
R9969 GND.n10056 GND.n10055 585
R9970 GND.n10055 GND.n10054 585
R9971 GND.n857 GND.n856 585
R9972 GND.n856 GND.n855 585
R9973 GND.n10061 GND.n10060 585
R9974 GND.n10062 GND.n10061 585
R9975 GND.n854 GND.n853 585
R9976 GND.n10063 GND.n854 585
R9977 GND.n10066 GND.n10065 585
R9978 GND.n10065 GND.n10064 585
R9979 GND.n851 GND.n850 585
R9980 GND.n850 GND.n849 585
R9981 GND.n10071 GND.n10070 585
R9982 GND.n10072 GND.n10071 585
R9983 GND.n848 GND.n847 585
R9984 GND.n10073 GND.n848 585
R9985 GND.n10076 GND.n10075 585
R9986 GND.n10075 GND.n10074 585
R9987 GND.n845 GND.n844 585
R9988 GND.n844 GND.n843 585
R9989 GND.n10081 GND.n10080 585
R9990 GND.n10082 GND.n10081 585
R9991 GND.n842 GND.n841 585
R9992 GND.n10083 GND.n842 585
R9993 GND.n10086 GND.n10085 585
R9994 GND.n10085 GND.n10084 585
R9995 GND.n839 GND.n838 585
R9996 GND.n838 GND.n837 585
R9997 GND.n10091 GND.n10090 585
R9998 GND.n10092 GND.n10091 585
R9999 GND.n836 GND.n835 585
R10000 GND.n10093 GND.n836 585
R10001 GND.n10096 GND.n10095 585
R10002 GND.n10095 GND.n10094 585
R10003 GND.n833 GND.n832 585
R10004 GND.n832 GND.n831 585
R10005 GND.n10101 GND.n10100 585
R10006 GND.n10102 GND.n10101 585
R10007 GND.n830 GND.n829 585
R10008 GND.n10103 GND.n830 585
R10009 GND.n10106 GND.n10105 585
R10010 GND.n10105 GND.n10104 585
R10011 GND.n827 GND.n826 585
R10012 GND.n826 GND.n825 585
R10013 GND.n10111 GND.n10110 585
R10014 GND.n10112 GND.n10111 585
R10015 GND.n824 GND.n823 585
R10016 GND.n10113 GND.n824 585
R10017 GND.n10116 GND.n10115 585
R10018 GND.n10115 GND.n10114 585
R10019 GND.n821 GND.n820 585
R10020 GND.n820 GND.n819 585
R10021 GND.n10121 GND.n10120 585
R10022 GND.n10122 GND.n10121 585
R10023 GND.n818 GND.n817 585
R10024 GND.n10123 GND.n818 585
R10025 GND.n10126 GND.n10125 585
R10026 GND.n10125 GND.n10124 585
R10027 GND.n815 GND.n814 585
R10028 GND.n814 GND.n813 585
R10029 GND.n10131 GND.n10130 585
R10030 GND.n10132 GND.n10131 585
R10031 GND.n812 GND.n811 585
R10032 GND.n10133 GND.n812 585
R10033 GND.n10136 GND.n10135 585
R10034 GND.n10135 GND.n10134 585
R10035 GND.n809 GND.n808 585
R10036 GND.n808 GND.n807 585
R10037 GND.n10141 GND.n10140 585
R10038 GND.n10142 GND.n10141 585
R10039 GND.n806 GND.n805 585
R10040 GND.n10143 GND.n806 585
R10041 GND.n10146 GND.n10145 585
R10042 GND.n10145 GND.n10144 585
R10043 GND.n803 GND.n802 585
R10044 GND.n802 GND.n801 585
R10045 GND.n10151 GND.n10150 585
R10046 GND.n10152 GND.n10151 585
R10047 GND.n800 GND.n799 585
R10048 GND.n10153 GND.n800 585
R10049 GND.n10156 GND.n10155 585
R10050 GND.n10155 GND.n10154 585
R10051 GND.n797 GND.n796 585
R10052 GND.n796 GND.n795 585
R10053 GND.n10161 GND.n10160 585
R10054 GND.n10162 GND.n10161 585
R10055 GND.n794 GND.n793 585
R10056 GND.n10163 GND.n794 585
R10057 GND.n10166 GND.n10165 585
R10058 GND.n10165 GND.n10164 585
R10059 GND.n791 GND.n790 585
R10060 GND.n790 GND.n789 585
R10061 GND.n10171 GND.n10170 585
R10062 GND.n10172 GND.n10171 585
R10063 GND.n788 GND.n787 585
R10064 GND.n10173 GND.n788 585
R10065 GND.n10176 GND.n10175 585
R10066 GND.n10175 GND.n10174 585
R10067 GND.n785 GND.n784 585
R10068 GND.n784 GND.n783 585
R10069 GND.n10181 GND.n10180 585
R10070 GND.n10182 GND.n10181 585
R10071 GND.n782 GND.n781 585
R10072 GND.n10183 GND.n782 585
R10073 GND.n10186 GND.n10185 585
R10074 GND.n10185 GND.n10184 585
R10075 GND.n779 GND.n778 585
R10076 GND.n778 GND.n777 585
R10077 GND.n10191 GND.n10190 585
R10078 GND.n10192 GND.n10191 585
R10079 GND.n776 GND.n775 585
R10080 GND.n10193 GND.n776 585
R10081 GND.n10196 GND.n10195 585
R10082 GND.n10195 GND.n10194 585
R10083 GND.n773 GND.n772 585
R10084 GND.n772 GND.n771 585
R10085 GND.n10201 GND.n10200 585
R10086 GND.n10202 GND.n10201 585
R10087 GND.n770 GND.n769 585
R10088 GND.n10203 GND.n770 585
R10089 GND.n10206 GND.n10205 585
R10090 GND.n10205 GND.n10204 585
R10091 GND.n767 GND.n766 585
R10092 GND.n766 GND.n765 585
R10093 GND.n10211 GND.n10210 585
R10094 GND.n10212 GND.n10211 585
R10095 GND.n764 GND.n763 585
R10096 GND.n10213 GND.n764 585
R10097 GND.n10216 GND.n10215 585
R10098 GND.n10215 GND.n10214 585
R10099 GND.n761 GND.n760 585
R10100 GND.n760 GND.n759 585
R10101 GND.n10221 GND.n10220 585
R10102 GND.n10222 GND.n10221 585
R10103 GND.n758 GND.n757 585
R10104 GND.n10223 GND.n758 585
R10105 GND.n10226 GND.n10225 585
R10106 GND.n10225 GND.n10224 585
R10107 GND.n755 GND.n754 585
R10108 GND.n754 GND.n753 585
R10109 GND.n10231 GND.n10230 585
R10110 GND.n10232 GND.n10231 585
R10111 GND.n752 GND.n751 585
R10112 GND.n10233 GND.n752 585
R10113 GND.n10236 GND.n10235 585
R10114 GND.n10235 GND.n10234 585
R10115 GND.n749 GND.n748 585
R10116 GND.n748 GND.n747 585
R10117 GND.n10241 GND.n10240 585
R10118 GND.n10242 GND.n10241 585
R10119 GND.n746 GND.n745 585
R10120 GND.n10243 GND.n746 585
R10121 GND.n10246 GND.n10245 585
R10122 GND.n10245 GND.n10244 585
R10123 GND.n743 GND.n742 585
R10124 GND.n742 GND.n741 585
R10125 GND.n10251 GND.n10250 585
R10126 GND.n10252 GND.n10251 585
R10127 GND.n740 GND.n739 585
R10128 GND.n10253 GND.n740 585
R10129 GND.n10256 GND.n10255 585
R10130 GND.n10255 GND.n10254 585
R10131 GND.n737 GND.n736 585
R10132 GND.n736 GND.n735 585
R10133 GND.n10261 GND.n10260 585
R10134 GND.n10262 GND.n10261 585
R10135 GND.n734 GND.n733 585
R10136 GND.n10263 GND.n734 585
R10137 GND.n10266 GND.n10265 585
R10138 GND.n10265 GND.n10264 585
R10139 GND.n731 GND.n730 585
R10140 GND.n730 GND.n729 585
R10141 GND.n10271 GND.n10270 585
R10142 GND.n10272 GND.n10271 585
R10143 GND.n728 GND.n727 585
R10144 GND.n10273 GND.n728 585
R10145 GND.n10276 GND.n10275 585
R10146 GND.n10275 GND.n10274 585
R10147 GND.n725 GND.n724 585
R10148 GND.n724 GND.n723 585
R10149 GND.n10281 GND.n10280 585
R10150 GND.n10282 GND.n10281 585
R10151 GND.n722 GND.n721 585
R10152 GND.n10283 GND.n722 585
R10153 GND.n10286 GND.n10285 585
R10154 GND.n10285 GND.n10284 585
R10155 GND.n719 GND.n718 585
R10156 GND.n718 GND.n717 585
R10157 GND.n10291 GND.n10290 585
R10158 GND.n10292 GND.n10291 585
R10159 GND.n716 GND.n715 585
R10160 GND.n10293 GND.n716 585
R10161 GND.n10296 GND.n10295 585
R10162 GND.n10295 GND.n10294 585
R10163 GND.n713 GND.n712 585
R10164 GND.n712 GND.n711 585
R10165 GND.n10301 GND.n10300 585
R10166 GND.n10302 GND.n10301 585
R10167 GND.n710 GND.n709 585
R10168 GND.n10303 GND.n710 585
R10169 GND.n10306 GND.n10305 585
R10170 GND.n10305 GND.n10304 585
R10171 GND.n707 GND.n706 585
R10172 GND.n706 GND.n705 585
R10173 GND.n10311 GND.n10310 585
R10174 GND.n10312 GND.n10311 585
R10175 GND.n704 GND.n703 585
R10176 GND.n10313 GND.n704 585
R10177 GND.n10316 GND.n10315 585
R10178 GND.n10315 GND.n10314 585
R10179 GND.n701 GND.n700 585
R10180 GND.n700 GND.n699 585
R10181 GND.n10321 GND.n10320 585
R10182 GND.n10322 GND.n10321 585
R10183 GND.n698 GND.n697 585
R10184 GND.n10323 GND.n698 585
R10185 GND.n10326 GND.n10325 585
R10186 GND.n10325 GND.n10324 585
R10187 GND.n695 GND.n694 585
R10188 GND.n694 GND.n693 585
R10189 GND.n10331 GND.n10330 585
R10190 GND.n10332 GND.n10331 585
R10191 GND.n692 GND.n691 585
R10192 GND.n10333 GND.n692 585
R10193 GND.n10336 GND.n10335 585
R10194 GND.n10335 GND.n10334 585
R10195 GND.n689 GND.n688 585
R10196 GND.n688 GND.n687 585
R10197 GND.n10341 GND.n10340 585
R10198 GND.n10342 GND.n10341 585
R10199 GND.n686 GND.n685 585
R10200 GND.n10343 GND.n686 585
R10201 GND.n10346 GND.n10345 585
R10202 GND.n10345 GND.n10344 585
R10203 GND.n683 GND.n682 585
R10204 GND.n682 GND.n681 585
R10205 GND.n10351 GND.n10350 585
R10206 GND.n10352 GND.n10351 585
R10207 GND.n680 GND.n679 585
R10208 GND.n10353 GND.n680 585
R10209 GND.n10356 GND.n10355 585
R10210 GND.n10355 GND.n10354 585
R10211 GND.n677 GND.n676 585
R10212 GND.n676 GND.n675 585
R10213 GND.n10361 GND.n10360 585
R10214 GND.n10362 GND.n10361 585
R10215 GND.n674 GND.n673 585
R10216 GND.n10363 GND.n674 585
R10217 GND.n10366 GND.n10365 585
R10218 GND.n10365 GND.n10364 585
R10219 GND.n671 GND.n670 585
R10220 GND.n670 GND.n669 585
R10221 GND.n10371 GND.n10370 585
R10222 GND.n10372 GND.n10371 585
R10223 GND.n668 GND.n667 585
R10224 GND.n10373 GND.n668 585
R10225 GND.n10376 GND.n10375 585
R10226 GND.n10375 GND.n10374 585
R10227 GND.n665 GND.n664 585
R10228 GND.n664 GND.n663 585
R10229 GND.n10382 GND.n10381 585
R10230 GND.n10383 GND.n10382 585
R10231 GND.n10380 GND.n662 585
R10232 GND.n10384 GND.n662 585
R10233 GND.n10533 GND.n10532 585
R10234 GND.n10534 GND.n10533 585
R10235 GND.n576 GND.n575 585
R10236 GND.n575 GND.n574 585
R10237 GND.n10527 GND.n10526 585
R10238 GND.n10526 GND.n10525 585
R10239 GND.n579 GND.n578 585
R10240 GND.n10524 GND.n579 585
R10241 GND.n10522 GND.n10521 585
R10242 GND.n10523 GND.n10522 585
R10243 GND.n582 GND.n581 585
R10244 GND.n581 GND.n580 585
R10245 GND.n10517 GND.n10516 585
R10246 GND.n10516 GND.n10515 585
R10247 GND.n585 GND.n584 585
R10248 GND.n10514 GND.n585 585
R10249 GND.n10512 GND.n10511 585
R10250 GND.n10513 GND.n10512 585
R10251 GND.n588 GND.n587 585
R10252 GND.n587 GND.n586 585
R10253 GND.n10507 GND.n10506 585
R10254 GND.n10506 GND.n10505 585
R10255 GND.n591 GND.n590 585
R10256 GND.n10504 GND.n591 585
R10257 GND.n10502 GND.n10501 585
R10258 GND.n10503 GND.n10502 585
R10259 GND.n594 GND.n593 585
R10260 GND.n593 GND.n592 585
R10261 GND.n10497 GND.n10496 585
R10262 GND.n10496 GND.n10495 585
R10263 GND.n597 GND.n596 585
R10264 GND.n10494 GND.n597 585
R10265 GND.n10492 GND.n10491 585
R10266 GND.n10493 GND.n10492 585
R10267 GND.n600 GND.n599 585
R10268 GND.n599 GND.n598 585
R10269 GND.n10487 GND.n10486 585
R10270 GND.n10486 GND.n10485 585
R10271 GND.n603 GND.n602 585
R10272 GND.n10484 GND.n603 585
R10273 GND.n10482 GND.n10481 585
R10274 GND.n10483 GND.n10482 585
R10275 GND.n606 GND.n605 585
R10276 GND.n605 GND.n604 585
R10277 GND.n10477 GND.n10476 585
R10278 GND.n10476 GND.n10475 585
R10279 GND.n609 GND.n608 585
R10280 GND.n10474 GND.n609 585
R10281 GND.n10472 GND.n10471 585
R10282 GND.n10473 GND.n10472 585
R10283 GND.n612 GND.n611 585
R10284 GND.n611 GND.n610 585
R10285 GND.n10467 GND.n10466 585
R10286 GND.n10466 GND.n10465 585
R10287 GND.n615 GND.n614 585
R10288 GND.n10464 GND.n615 585
R10289 GND.n10462 GND.n10461 585
R10290 GND.n10463 GND.n10462 585
R10291 GND.n618 GND.n617 585
R10292 GND.n617 GND.n616 585
R10293 GND.n10457 GND.n10456 585
R10294 GND.n10456 GND.n10455 585
R10295 GND.n621 GND.n620 585
R10296 GND.n10454 GND.n621 585
R10297 GND.n10452 GND.n10451 585
R10298 GND.n10453 GND.n10452 585
R10299 GND.n624 GND.n623 585
R10300 GND.n623 GND.n622 585
R10301 GND.n10447 GND.n10446 585
R10302 GND.n10446 GND.n10445 585
R10303 GND.n627 GND.n626 585
R10304 GND.n10444 GND.n627 585
R10305 GND.n10442 GND.n10441 585
R10306 GND.n10443 GND.n10442 585
R10307 GND.n630 GND.n629 585
R10308 GND.n629 GND.n628 585
R10309 GND.n10437 GND.n10436 585
R10310 GND.n10436 GND.n10435 585
R10311 GND.n633 GND.n632 585
R10312 GND.n10434 GND.n633 585
R10313 GND.n10432 GND.n10431 585
R10314 GND.n10433 GND.n10432 585
R10315 GND.n636 GND.n635 585
R10316 GND.n635 GND.n634 585
R10317 GND.n10427 GND.n10426 585
R10318 GND.n10426 GND.n10425 585
R10319 GND.n639 GND.n638 585
R10320 GND.n10424 GND.n639 585
R10321 GND.n10422 GND.n10421 585
R10322 GND.n10423 GND.n10422 585
R10323 GND.n642 GND.n641 585
R10324 GND.n641 GND.n640 585
R10325 GND.n10417 GND.n10416 585
R10326 GND.n10416 GND.n10415 585
R10327 GND.n645 GND.n644 585
R10328 GND.n10414 GND.n645 585
R10329 GND.n10412 GND.n10411 585
R10330 GND.n10413 GND.n10412 585
R10331 GND.n648 GND.n647 585
R10332 GND.n647 GND.n646 585
R10333 GND.n10407 GND.n10406 585
R10334 GND.n10406 GND.n10405 585
R10335 GND.n651 GND.n650 585
R10336 GND.n10404 GND.n651 585
R10337 GND.n10402 GND.n10401 585
R10338 GND.n10403 GND.n10402 585
R10339 GND.n654 GND.n653 585
R10340 GND.n653 GND.n652 585
R10341 GND.n10397 GND.n10396 585
R10342 GND.n10396 GND.n10395 585
R10343 GND.n657 GND.n656 585
R10344 GND.n10394 GND.n657 585
R10345 GND.n10392 GND.n10391 585
R10346 GND.n10393 GND.n10392 585
R10347 GND.n660 GND.n659 585
R10348 GND.n659 GND.n658 585
R10349 GND.n10387 GND.n10386 585
R10350 GND.n10386 GND.n10385 585
R10351 GND.n10911 GND.n10910 585
R10352 GND.n10912 GND.n10911 585
R10353 GND.n434 GND.n433 585
R10354 GND.n10905 GND.n434 585
R10355 GND.n10920 GND.n10919 585
R10356 GND.n10919 GND.n10918 585
R10357 GND.n10921 GND.n429 585
R10358 GND.n7166 GND.n429 585
R10359 GND.n10923 GND.n10922 585
R10360 GND.n10924 GND.n10923 585
R10361 GND.n413 GND.n412 585
R10362 GND.n7172 GND.n413 585
R10363 GND.n10932 GND.n10931 585
R10364 GND.n10931 GND.n10930 585
R10365 GND.n10933 GND.n408 585
R10366 GND.n7178 GND.n408 585
R10367 GND.n10935 GND.n10934 585
R10368 GND.n10936 GND.n10935 585
R10369 GND.n392 GND.n391 585
R10370 GND.n7184 GND.n392 585
R10371 GND.n10944 GND.n10943 585
R10372 GND.n10943 GND.n10942 585
R10373 GND.n10945 GND.n387 585
R10374 GND.n7190 GND.n387 585
R10375 GND.n10947 GND.n10946 585
R10376 GND.n10948 GND.n10947 585
R10377 GND.n371 GND.n370 585
R10378 GND.n7196 GND.n371 585
R10379 GND.n10956 GND.n10955 585
R10380 GND.n10955 GND.n10954 585
R10381 GND.n10957 GND.n366 585
R10382 GND.n7202 GND.n366 585
R10383 GND.n10959 GND.n10958 585
R10384 GND.n10960 GND.n10959 585
R10385 GND.n350 GND.n349 585
R10386 GND.n7208 GND.n350 585
R10387 GND.n10968 GND.n10967 585
R10388 GND.n10967 GND.n10966 585
R10389 GND.n10969 GND.n345 585
R10390 GND.n7214 GND.n345 585
R10391 GND.n10971 GND.n10970 585
R10392 GND.n10972 GND.n10971 585
R10393 GND.n329 GND.n328 585
R10394 GND.n7220 GND.n329 585
R10395 GND.n10980 GND.n10979 585
R10396 GND.n10979 GND.n10978 585
R10397 GND.n10981 GND.n324 585
R10398 GND.n7226 GND.n324 585
R10399 GND.n10983 GND.n10982 585
R10400 GND.n10984 GND.n10983 585
R10401 GND.n308 GND.n307 585
R10402 GND.n7232 GND.n308 585
R10403 GND.n10992 GND.n10991 585
R10404 GND.n10991 GND.n10990 585
R10405 GND.n10993 GND.n303 585
R10406 GND.n7238 GND.n303 585
R10407 GND.n10995 GND.n10994 585
R10408 GND.n10996 GND.n10995 585
R10409 GND.n287 GND.n286 585
R10410 GND.n7244 GND.n287 585
R10411 GND.n11004 GND.n11003 585
R10412 GND.n11003 GND.n11002 585
R10413 GND.n11005 GND.n282 585
R10414 GND.n7250 GND.n282 585
R10415 GND.n11007 GND.n11006 585
R10416 GND.n11008 GND.n11007 585
R10417 GND.n266 GND.n265 585
R10418 GND.n7256 GND.n266 585
R10419 GND.n11016 GND.n11015 585
R10420 GND.n11015 GND.n11014 585
R10421 GND.n11017 GND.n261 585
R10422 GND.n7262 GND.n261 585
R10423 GND.n11019 GND.n11018 585
R10424 GND.n11020 GND.n11019 585
R10425 GND.n246 GND.n245 585
R10426 GND.n7268 GND.n246 585
R10427 GND.n11028 GND.n11027 585
R10428 GND.n11027 GND.n11026 585
R10429 GND.n11029 GND.n241 585
R10430 GND.n7101 GND.n241 585
R10431 GND.n11031 GND.n11030 585
R10432 GND.n11032 GND.n11031 585
R10433 GND.n225 GND.n224 585
R10434 GND.n7092 GND.n225 585
R10435 GND.n11040 GND.n11039 585
R10436 GND.n11039 GND.n11038 585
R10437 GND.n11041 GND.n220 585
R10438 GND.n7085 GND.n220 585
R10439 GND.n11043 GND.n11042 585
R10440 GND.n11044 GND.n11043 585
R10441 GND.n204 GND.n203 585
R10442 GND.n7077 GND.n204 585
R10443 GND.n11052 GND.n11051 585
R10444 GND.n11051 GND.n11050 585
R10445 GND.n11053 GND.n199 585
R10446 GND.n7070 GND.n199 585
R10447 GND.n11055 GND.n11054 585
R10448 GND.n11056 GND.n11055 585
R10449 GND.n183 GND.n182 585
R10450 GND.n7062 GND.n183 585
R10451 GND.n11064 GND.n11063 585
R10452 GND.n11063 GND.n11062 585
R10453 GND.n11065 GND.n178 585
R10454 GND.n7055 GND.n178 585
R10455 GND.n11067 GND.n11066 585
R10456 GND.n11068 GND.n11067 585
R10457 GND.n162 GND.n161 585
R10458 GND.n7047 GND.n162 585
R10459 GND.n11076 GND.n11075 585
R10460 GND.n11075 GND.n11074 585
R10461 GND.n11077 GND.n157 585
R10462 GND.n7040 GND.n157 585
R10463 GND.n11079 GND.n11078 585
R10464 GND.n11080 GND.n11079 585
R10465 GND.n141 GND.n140 585
R10466 GND.n7032 GND.n141 585
R10467 GND.n11088 GND.n11087 585
R10468 GND.n11087 GND.n11086 585
R10469 GND.n11089 GND.n136 585
R10470 GND.n7025 GND.n136 585
R10471 GND.n11091 GND.n11090 585
R10472 GND.n11092 GND.n11091 585
R10473 GND.n122 GND.n121 585
R10474 GND.n7017 GND.n122 585
R10475 GND.n11100 GND.n11099 585
R10476 GND.n11099 GND.n11098 585
R10477 GND.n11101 GND.n116 585
R10478 GND.n7312 GND.n116 585
R10479 GND.n11103 GND.n11102 585
R10480 GND.n11104 GND.n11103 585
R10481 GND.n117 GND.n115 585
R10482 GND.n7318 GND.n115 585
R10483 GND.n7007 GND.n7006 585
R10484 GND.n7006 GND.n6269 585
R10485 GND.n7005 GND.n6465 585
R10486 GND.n7005 GND.n7004 585
R10487 GND.n6998 GND.n95 585
R10488 GND.n11111 GND.n95 585
R10489 GND.n6997 GND.n6996 585
R10490 GND.n6996 GND.n6995 585
R10491 GND.n6470 GND.n6469 585
R10492 GND.n6470 GND.n6259 585
R10493 GND.n6250 GND.n6249 585
R10494 GND.n7333 GND.n6250 585
R10495 GND.n7339 GND.n7338 585
R10496 GND.n7338 GND.n7337 585
R10497 GND.n7340 GND.n6245 585
R10498 GND.n6985 GND.n6245 585
R10499 GND.n7342 GND.n7341 585
R10500 GND.n7343 GND.n7342 585
R10501 GND.n6230 GND.n6229 585
R10502 GND.n6970 GND.n6230 585
R10503 GND.n7351 GND.n7350 585
R10504 GND.n7350 GND.n7349 585
R10505 GND.n7352 GND.n6225 585
R10506 GND.n6963 GND.n6225 585
R10507 GND.n7354 GND.n7353 585
R10508 GND.n7355 GND.n7354 585
R10509 GND.n6209 GND.n6208 585
R10510 GND.n6955 GND.n6209 585
R10511 GND.n7363 GND.n7362 585
R10512 GND.n7362 GND.n7361 585
R10513 GND.n7364 GND.n6204 585
R10514 GND.n6948 GND.n6204 585
R10515 GND.n7366 GND.n7365 585
R10516 GND.n7367 GND.n7366 585
R10517 GND.n6188 GND.n6187 585
R10518 GND.n6940 GND.n6188 585
R10519 GND.n7375 GND.n7374 585
R10520 GND.n7374 GND.n7373 585
R10521 GND.n7376 GND.n6183 585
R10522 GND.n6933 GND.n6183 585
R10523 GND.n7378 GND.n7377 585
R10524 GND.n7379 GND.n7378 585
R10525 GND.n6168 GND.n6167 585
R10526 GND.n6925 GND.n6168 585
R10527 GND.n7387 GND.n7386 585
R10528 GND.n7386 GND.n7385 585
R10529 GND.n7388 GND.n6163 585
R10530 GND.n6918 GND.n6163 585
R10531 GND.n7390 GND.n7389 585
R10532 GND.n7391 GND.n7390 585
R10533 GND.n6147 GND.n6146 585
R10534 GND.n6910 GND.n6147 585
R10535 GND.n7399 GND.n7398 585
R10536 GND.n7398 GND.n7397 585
R10537 GND.n7400 GND.n6142 585
R10538 GND.n6903 GND.n6142 585
R10539 GND.n7402 GND.n7401 585
R10540 GND.n7403 GND.n7402 585
R10541 GND.n6126 GND.n6125 585
R10542 GND.n6895 GND.n6126 585
R10543 GND.n7411 GND.n7410 585
R10544 GND.n7410 GND.n7409 585
R10545 GND.n7412 GND.n6121 585
R10546 GND.n6888 GND.n6121 585
R10547 GND.n7414 GND.n7413 585
R10548 GND.n7415 GND.n7414 585
R10549 GND.n6105 GND.n6104 585
R10550 GND.n6880 GND.n6105 585
R10551 GND.n7423 GND.n7422 585
R10552 GND.n7422 GND.n7421 585
R10553 GND.n7424 GND.n6100 585
R10554 GND.n6873 GND.n6100 585
R10555 GND.n7426 GND.n7425 585
R10556 GND.n7427 GND.n7426 585
R10557 GND.n6084 GND.n6083 585
R10558 GND.n6865 GND.n6084 585
R10559 GND.n7435 GND.n7434 585
R10560 GND.n7434 GND.n7433 585
R10561 GND.n7436 GND.n6079 585
R10562 GND.n6858 GND.n6079 585
R10563 GND.n7438 GND.n7437 585
R10564 GND.n7439 GND.n7438 585
R10565 GND.n6063 GND.n6062 585
R10566 GND.n6850 GND.n6063 585
R10567 GND.n7447 GND.n7446 585
R10568 GND.n7446 GND.n7445 585
R10569 GND.n7448 GND.n6058 585
R10570 GND.n6843 GND.n6058 585
R10571 GND.n7450 GND.n7449 585
R10572 GND.n7451 GND.n7450 585
R10573 GND.n6042 GND.n6041 585
R10574 GND.n6835 GND.n6042 585
R10575 GND.n7459 GND.n7458 585
R10576 GND.n7458 GND.n7457 585
R10577 GND.n7460 GND.n6037 585
R10578 GND.n6828 GND.n6037 585
R10579 GND.n7462 GND.n7461 585
R10580 GND.n7463 GND.n7462 585
R10581 GND.n6022 GND.n6021 585
R10582 GND.n6820 GND.n6022 585
R10583 GND.n7471 GND.n7470 585
R10584 GND.n7470 GND.n7469 585
R10585 GND.n7472 GND.n6017 585
R10586 GND.n6813 GND.n6017 585
R10587 GND.n7474 GND.n7473 585
R10588 GND.n7475 GND.n7474 585
R10589 GND.n6001 GND.n6000 585
R10590 GND.n6805 GND.n6001 585
R10591 GND.n7483 GND.n7482 585
R10592 GND.n7482 GND.n7481 585
R10593 GND.n7484 GND.n5996 585
R10594 GND.n6798 GND.n5996 585
R10595 GND.n7486 GND.n7485 585
R10596 GND.n7487 GND.n7486 585
R10597 GND.n5980 GND.n5979 585
R10598 GND.n6790 GND.n5980 585
R10599 GND.n7495 GND.n7494 585
R10600 GND.n7494 GND.n7493 585
R10601 GND.n7496 GND.n5975 585
R10602 GND.n6783 GND.n5975 585
R10603 GND.n7498 GND.n7497 585
R10604 GND.n7499 GND.n7498 585
R10605 GND.n5959 GND.n5958 585
R10606 GND.n6775 GND.n5959 585
R10607 GND.n7507 GND.n7506 585
R10608 GND.n7506 GND.n7505 585
R10609 GND.n7508 GND.n5954 585
R10610 GND.n6768 GND.n5954 585
R10611 GND.n7510 GND.n7509 585
R10612 GND.n7511 GND.n7510 585
R10613 GND.n5939 GND.n5938 585
R10614 GND.n6760 GND.n5939 585
R10615 GND.n7519 GND.n7518 585
R10616 GND.n7518 GND.n7517 585
R10617 GND.n7520 GND.n5933 585
R10618 GND.n6753 GND.n5933 585
R10619 GND.n7522 GND.n7521 585
R10620 GND.n7523 GND.n7522 585
R10621 GND.n5934 GND.n5917 585
R10622 GND.n6745 GND.n5917 585
R10623 GND.n7530 GND.n5918 585
R10624 GND.n7530 GND.n7529 585
R10625 GND.n7531 GND.n5874 585
R10626 GND.n7532 GND.n7531 585
R10627 GND.n5914 GND.n5913 585
R10628 GND.n5912 GND.n5911 585
R10629 GND.n5909 GND.n5908 585
R10630 GND.n5907 GND.n5906 585
R10631 GND.n5904 GND.n5903 585
R10632 GND.n5902 GND.n5901 585
R10633 GND.n5899 GND.n5898 585
R10634 GND.n5897 GND.n5896 585
R10635 GND.n5894 GND.n5893 585
R10636 GND.n5892 GND.n5891 585
R10637 GND.n5889 GND.n5882 585
R10638 GND.n5888 GND.n5885 585
R10639 GND.n10899 GND.n10898 585
R10640 GND.n459 GND.n458 585
R10641 GND.n10665 GND.n10664 585
R10642 GND.n10667 GND.n10666 585
R10643 GND.n10669 GND.n10668 585
R10644 GND.n10671 GND.n10670 585
R10645 GND.n10673 GND.n10672 585
R10646 GND.n10675 GND.n10674 585
R10647 GND.n10677 GND.n10676 585
R10648 GND.n10679 GND.n10678 585
R10649 GND.n10681 GND.n10680 585
R10650 GND.n10654 GND.n10652 585
R10651 GND.n10686 GND.n10685 585
R10652 GND.n10653 GND.n449 585
R10653 GND.n10902 GND.n447 585
R10654 GND.n10912 GND.n447 585
R10655 GND.n10904 GND.n10903 585
R10656 GND.n10905 GND.n10904 585
R10657 GND.n453 GND.n437 585
R10658 GND.n10918 GND.n437 585
R10659 GND.n7168 GND.n7167 585
R10660 GND.n7167 GND.n7166 585
R10661 GND.n7169 GND.n427 585
R10662 GND.n10924 GND.n427 585
R10663 GND.n7171 GND.n7170 585
R10664 GND.n7172 GND.n7171 585
R10665 GND.n7156 GND.n416 585
R10666 GND.n10930 GND.n416 585
R10667 GND.n7180 GND.n7179 585
R10668 GND.n7179 GND.n7178 585
R10669 GND.n7181 GND.n406 585
R10670 GND.n10936 GND.n406 585
R10671 GND.n7183 GND.n7182 585
R10672 GND.n7184 GND.n7183 585
R10673 GND.n7149 GND.n395 585
R10674 GND.n10942 GND.n395 585
R10675 GND.n7192 GND.n7191 585
R10676 GND.n7191 GND.n7190 585
R10677 GND.n7193 GND.n385 585
R10678 GND.n10948 GND.n385 585
R10679 GND.n7195 GND.n7194 585
R10680 GND.n7196 GND.n7195 585
R10681 GND.n7142 GND.n374 585
R10682 GND.n10954 GND.n374 585
R10683 GND.n7204 GND.n7203 585
R10684 GND.n7203 GND.n7202 585
R10685 GND.n7205 GND.n364 585
R10686 GND.n10960 GND.n364 585
R10687 GND.n7207 GND.n7206 585
R10688 GND.n7208 GND.n7207 585
R10689 GND.n7135 GND.n353 585
R10690 GND.n10966 GND.n353 585
R10691 GND.n7216 GND.n7215 585
R10692 GND.n7215 GND.n7214 585
R10693 GND.n7217 GND.n343 585
R10694 GND.n10972 GND.n343 585
R10695 GND.n7219 GND.n7218 585
R10696 GND.n7220 GND.n7219 585
R10697 GND.n7128 GND.n332 585
R10698 GND.n10978 GND.n332 585
R10699 GND.n7228 GND.n7227 585
R10700 GND.n7227 GND.n7226 585
R10701 GND.n7229 GND.n322 585
R10702 GND.n10984 GND.n322 585
R10703 GND.n7231 GND.n7230 585
R10704 GND.n7232 GND.n7231 585
R10705 GND.n7121 GND.n311 585
R10706 GND.n10990 GND.n311 585
R10707 GND.n7240 GND.n7239 585
R10708 GND.n7239 GND.n7238 585
R10709 GND.n7241 GND.n301 585
R10710 GND.n10996 GND.n301 585
R10711 GND.n7243 GND.n7242 585
R10712 GND.n7244 GND.n7243 585
R10713 GND.n7114 GND.n290 585
R10714 GND.n11002 GND.n290 585
R10715 GND.n7252 GND.n7251 585
R10716 GND.n7251 GND.n7250 585
R10717 GND.n7253 GND.n280 585
R10718 GND.n11008 GND.n280 585
R10719 GND.n7255 GND.n7254 585
R10720 GND.n7256 GND.n7255 585
R10721 GND.n6439 GND.n269 585
R10722 GND.n11014 GND.n269 585
R10723 GND.n7264 GND.n7263 585
R10724 GND.n7263 GND.n7262 585
R10725 GND.n7265 GND.n259 585
R10726 GND.n11020 GND.n259 585
R10727 GND.n7267 GND.n7266 585
R10728 GND.n7268 GND.n7267 585
R10729 GND.n6435 GND.n249 585
R10730 GND.n11026 GND.n249 585
R10731 GND.n7100 GND.n7099 585
R10732 GND.n7101 GND.n7100 585
R10733 GND.n6441 GND.n239 585
R10734 GND.n11032 GND.n239 585
R10735 GND.n7094 GND.n7093 585
R10736 GND.n7093 GND.n7092 585
R10737 GND.n6443 GND.n228 585
R10738 GND.n11038 GND.n228 585
R10739 GND.n7084 GND.n7083 585
R10740 GND.n7085 GND.n7084 585
R10741 GND.n6445 GND.n218 585
R10742 GND.n11044 GND.n218 585
R10743 GND.n7079 GND.n7078 585
R10744 GND.n7078 GND.n7077 585
R10745 GND.n6447 GND.n207 585
R10746 GND.n11050 GND.n207 585
R10747 GND.n7069 GND.n7068 585
R10748 GND.n7070 GND.n7069 585
R10749 GND.n6449 GND.n197 585
R10750 GND.n11056 GND.n197 585
R10751 GND.n7064 GND.n7063 585
R10752 GND.n7063 GND.n7062 585
R10753 GND.n6451 GND.n186 585
R10754 GND.n11062 GND.n186 585
R10755 GND.n7054 GND.n7053 585
R10756 GND.n7055 GND.n7054 585
R10757 GND.n6453 GND.n176 585
R10758 GND.n11068 GND.n176 585
R10759 GND.n7049 GND.n7048 585
R10760 GND.n7048 GND.n7047 585
R10761 GND.n6455 GND.n165 585
R10762 GND.n11074 GND.n165 585
R10763 GND.n7039 GND.n7038 585
R10764 GND.n7040 GND.n7039 585
R10765 GND.n6457 GND.n155 585
R10766 GND.n11080 GND.n155 585
R10767 GND.n7034 GND.n7033 585
R10768 GND.n7033 GND.n7032 585
R10769 GND.n6459 GND.n144 585
R10770 GND.n11086 GND.n144 585
R10771 GND.n7024 GND.n7023 585
R10772 GND.n7025 GND.n7024 585
R10773 GND.n6461 GND.n134 585
R10774 GND.n11092 GND.n134 585
R10775 GND.n7019 GND.n7018 585
R10776 GND.n7018 GND.n7017 585
R10777 GND.n6277 GND.n124 585
R10778 GND.n11098 GND.n124 585
R10779 GND.n7314 GND.n7313 585
R10780 GND.n7313 GND.n7312 585
R10781 GND.n7315 GND.n113 585
R10782 GND.n11104 GND.n113 585
R10783 GND.n7317 GND.n7316 585
R10784 GND.n7318 GND.n7317 585
R10785 GND.n6272 GND.n6271 585
R10786 GND.n6271 GND.n6269 585
R10787 GND.n91 GND.n89 585
R10788 GND.n7004 GND.n91 585
R10789 GND.n11113 GND.n11112 585
R10790 GND.n11112 GND.n11111 585
R10791 GND.n90 GND.n88 585
R10792 GND.n6995 GND.n90 585
R10793 GND.n6980 GND.n6979 585
R10794 GND.n6979 GND.n6259 585
R10795 GND.n6981 GND.n6258 585
R10796 GND.n7333 GND.n6258 585
R10797 GND.n6982 GND.n6253 585
R10798 GND.n7337 GND.n6253 585
R10799 GND.n6984 GND.n6983 585
R10800 GND.n6985 GND.n6984 585
R10801 GND.n6473 GND.n6243 585
R10802 GND.n7343 GND.n6243 585
R10803 GND.n6972 GND.n6971 585
R10804 GND.n6971 GND.n6970 585
R10805 GND.n6475 GND.n6233 585
R10806 GND.n7349 GND.n6233 585
R10807 GND.n6962 GND.n6961 585
R10808 GND.n6963 GND.n6962 585
R10809 GND.n6477 GND.n6223 585
R10810 GND.n7355 GND.n6223 585
R10811 GND.n6957 GND.n6956 585
R10812 GND.n6956 GND.n6955 585
R10813 GND.n6479 GND.n6212 585
R10814 GND.n7361 GND.n6212 585
R10815 GND.n6947 GND.n6946 585
R10816 GND.n6948 GND.n6947 585
R10817 GND.n6481 GND.n6202 585
R10818 GND.n7367 GND.n6202 585
R10819 GND.n6942 GND.n6941 585
R10820 GND.n6941 GND.n6940 585
R10821 GND.n6483 GND.n6191 585
R10822 GND.n7373 GND.n6191 585
R10823 GND.n6932 GND.n6931 585
R10824 GND.n6933 GND.n6932 585
R10825 GND.n6485 GND.n6181 585
R10826 GND.n7379 GND.n6181 585
R10827 GND.n6927 GND.n6926 585
R10828 GND.n6926 GND.n6925 585
R10829 GND.n6487 GND.n6171 585
R10830 GND.n7385 GND.n6171 585
R10831 GND.n6917 GND.n6916 585
R10832 GND.n6918 GND.n6917 585
R10833 GND.n6490 GND.n6161 585
R10834 GND.n7391 GND.n6161 585
R10835 GND.n6912 GND.n6911 585
R10836 GND.n6911 GND.n6910 585
R10837 GND.n6492 GND.n6150 585
R10838 GND.n7397 GND.n6150 585
R10839 GND.n6902 GND.n6901 585
R10840 GND.n6903 GND.n6902 585
R10841 GND.n6494 GND.n6140 585
R10842 GND.n7403 GND.n6140 585
R10843 GND.n6897 GND.n6896 585
R10844 GND.n6896 GND.n6895 585
R10845 GND.n6496 GND.n6129 585
R10846 GND.n7409 GND.n6129 585
R10847 GND.n6887 GND.n6886 585
R10848 GND.n6888 GND.n6887 585
R10849 GND.n6498 GND.n6119 585
R10850 GND.n7415 GND.n6119 585
R10851 GND.n6882 GND.n6881 585
R10852 GND.n6881 GND.n6880 585
R10853 GND.n6500 GND.n6108 585
R10854 GND.n7421 GND.n6108 585
R10855 GND.n6872 GND.n6871 585
R10856 GND.n6873 GND.n6872 585
R10857 GND.n6502 GND.n6098 585
R10858 GND.n7427 GND.n6098 585
R10859 GND.n6867 GND.n6866 585
R10860 GND.n6866 GND.n6865 585
R10861 GND.n6504 GND.n6087 585
R10862 GND.n7433 GND.n6087 585
R10863 GND.n6857 GND.n6856 585
R10864 GND.n6858 GND.n6857 585
R10865 GND.n6506 GND.n6077 585
R10866 GND.n7439 GND.n6077 585
R10867 GND.n6852 GND.n6851 585
R10868 GND.n6851 GND.n6850 585
R10869 GND.n6508 GND.n6066 585
R10870 GND.n7445 GND.n6066 585
R10871 GND.n6842 GND.n6841 585
R10872 GND.n6843 GND.n6842 585
R10873 GND.n6510 GND.n6056 585
R10874 GND.n7451 GND.n6056 585
R10875 GND.n6837 GND.n6836 585
R10876 GND.n6836 GND.n6835 585
R10877 GND.n6512 GND.n6045 585
R10878 GND.n7457 GND.n6045 585
R10879 GND.n6827 GND.n6826 585
R10880 GND.n6828 GND.n6827 585
R10881 GND.n6515 GND.n6036 585
R10882 GND.n7463 GND.n6036 585
R10883 GND.n6822 GND.n6821 585
R10884 GND.n6821 GND.n6820 585
R10885 GND.n6517 GND.n6025 585
R10886 GND.n7469 GND.n6025 585
R10887 GND.n6812 GND.n6811 585
R10888 GND.n6813 GND.n6812 585
R10889 GND.n6519 GND.n6015 585
R10890 GND.n7475 GND.n6015 585
R10891 GND.n6807 GND.n6806 585
R10892 GND.n6806 GND.n6805 585
R10893 GND.n6521 GND.n6004 585
R10894 GND.n7481 GND.n6004 585
R10895 GND.n6797 GND.n6796 585
R10896 GND.n6798 GND.n6797 585
R10897 GND.n6523 GND.n5994 585
R10898 GND.n7487 GND.n5994 585
R10899 GND.n6792 GND.n6791 585
R10900 GND.n6791 GND.n6790 585
R10901 GND.n6525 GND.n5983 585
R10902 GND.n7493 GND.n5983 585
R10903 GND.n6782 GND.n6781 585
R10904 GND.n6783 GND.n6782 585
R10905 GND.n6527 GND.n5973 585
R10906 GND.n7499 GND.n5973 585
R10907 GND.n6777 GND.n6776 585
R10908 GND.n6776 GND.n6775 585
R10909 GND.n6529 GND.n5962 585
R10910 GND.n7505 GND.n5962 585
R10911 GND.n6767 GND.n6766 585
R10912 GND.n6768 GND.n6767 585
R10913 GND.n6733 GND.n5953 585
R10914 GND.n7511 GND.n5953 585
R10915 GND.n6762 GND.n6761 585
R10916 GND.n6761 GND.n6760 585
R10917 GND.n6735 GND.n5942 585
R10918 GND.n7517 GND.n5942 585
R10919 GND.n6752 GND.n6751 585
R10920 GND.n6753 GND.n6752 585
R10921 GND.n6737 GND.n5931 585
R10922 GND.n7523 GND.n5931 585
R10923 GND.n6747 GND.n6746 585
R10924 GND.n6746 GND.n6745 585
R10925 GND.n6741 GND.n5919 585
R10926 GND.n7529 GND.n5919 585
R10927 GND.n6740 GND.n5880 585
R10928 GND.n7532 GND.n5880 585
R10929 GND.n5812 GND.n4367 585
R10930 GND.n7738 GND.n4367 585
R10931 GND.n5811 GND.n5810 585
R10932 GND.n5810 GND.n5809 585
R10933 GND.n5808 GND.n4356 585
R10934 GND.n7744 GND.n4356 585
R10935 GND.n4867 GND.n4850 585
R10936 GND.n5793 GND.n4867 585
R10937 GND.n5804 GND.n4347 585
R10938 GND.n7750 GND.n4347 585
R10939 GND.n5803 GND.n5802 585
R10940 GND.n5802 GND.n5801 585
R10941 GND.n4852 GND.n4337 585
R10942 GND.n7756 GND.n4337 585
R10943 GND.n5733 GND.n5732 585
R10944 GND.n5732 GND.n4872 585
R10945 GND.n5734 GND.n4327 585
R10946 GND.n7762 GND.n4327 585
R10947 GND.n5736 GND.n5735 585
R10948 GND.n5735 GND.n4877 585
R10949 GND.n5737 GND.n4317 585
R10950 GND.n7768 GND.n4317 585
R10951 GND.n5739 GND.n5738 585
R10952 GND.n5738 GND.n4882 585
R10953 GND.n5740 GND.n4294 585
R10954 GND.n7774 GND.n4294 585
R10955 GND.n5742 GND.n5741 585
R10956 GND.n5743 GND.n5742 585
R10957 GND.n4886 GND.n4280 585
R10958 GND.n7780 GND.n4280 585
R10959 GND.n5721 GND.n5720 585
R10960 GND.n5720 GND.n4272 585
R10961 GND.n5719 GND.n5718 585
R10962 GND.n5719 GND.n4271 585
R10963 GND.n5717 GND.n4263 585
R10964 GND.n7793 GND.n4263 585
R10965 GND.n4890 GND.n4889 585
R10966 GND.n4889 GND.n4888 585
R10967 GND.n5713 GND.n4252 585
R10968 GND.n7799 GND.n4252 585
R10969 GND.n5712 GND.n5711 585
R10970 GND.n5711 GND.n5710 585
R10971 GND.n4892 GND.n4243 585
R10972 GND.n7805 GND.n4243 585
R10973 GND.n5633 GND.n5632 585
R10974 GND.n5632 GND.n5631 585
R10975 GND.n5634 GND.n4234 585
R10976 GND.n7811 GND.n4234 585
R10977 GND.n5636 GND.n5635 585
R10978 GND.n5635 GND.n4905 585
R10979 GND.n5637 GND.n4224 585
R10980 GND.n7817 GND.n4224 585
R10981 GND.n5639 GND.n5638 585
R10982 GND.n5638 GND.n4910 585
R10983 GND.n5640 GND.n4214 585
R10984 GND.n7823 GND.n4214 585
R10985 GND.n5642 GND.n5641 585
R10986 GND.n5641 GND.n4915 585
R10987 GND.n5643 GND.n4192 585
R10988 GND.n7829 GND.n4192 585
R10989 GND.n5645 GND.n5644 585
R10990 GND.n5646 GND.n5645 585
R10991 GND.n4920 GND.n4178 585
R10992 GND.n7835 GND.n4178 585
R10993 GND.n5618 GND.n5617 585
R10994 GND.n5617 GND.n4170 585
R10995 GND.n5616 GND.n5615 585
R10996 GND.n5616 GND.n4169 585
R10997 GND.n5614 GND.n4161 585
R10998 GND.n7848 GND.n4161 585
R10999 GND.n4924 GND.n4923 585
R11000 GND.n4923 GND.n4922 585
R11001 GND.n5610 GND.n4150 585
R11002 GND.n7854 GND.n4150 585
R11003 GND.n5609 GND.n5608 585
R11004 GND.n5608 GND.n5607 585
R11005 GND.n4926 GND.n4140 585
R11006 GND.n7860 GND.n4140 585
R11007 GND.n5529 GND.n5528 585
R11008 GND.n5528 GND.n4932 585
R11009 GND.n5530 GND.n4130 585
R11010 GND.n7866 GND.n4130 585
R11011 GND.n5532 GND.n5531 585
R11012 GND.n5531 GND.n4937 585
R11013 GND.n5533 GND.n4120 585
R11014 GND.n7872 GND.n4120 585
R11015 GND.n5535 GND.n5534 585
R11016 GND.n5534 GND.n4942 585
R11017 GND.n5536 GND.n4110 585
R11018 GND.n7878 GND.n4110 585
R11019 GND.n5538 GND.n5537 585
R11020 GND.n5537 GND.n4947 585
R11021 GND.n5539 GND.n4087 585
R11022 GND.n7884 GND.n4087 585
R11023 GND.n5541 GND.n5540 585
R11024 GND.n5542 GND.n5541 585
R11025 GND.n4951 GND.n4073 585
R11026 GND.n7890 GND.n4073 585
R11027 GND.n5515 GND.n5514 585
R11028 GND.n5514 GND.n4065 585
R11029 GND.n5513 GND.n5512 585
R11030 GND.n5513 GND.n4064 585
R11031 GND.n5511 GND.n4056 585
R11032 GND.n7903 GND.n4056 585
R11033 GND.n4955 GND.n4954 585
R11034 GND.n4954 GND.n4953 585
R11035 GND.n5507 GND.n4045 585
R11036 GND.n7909 GND.n4045 585
R11037 GND.n5506 GND.n5505 585
R11038 GND.n5505 GND.n5504 585
R11039 GND.n4957 GND.n4035 585
R11040 GND.n7915 GND.n4035 585
R11041 GND.n5386 GND.n5385 585
R11042 GND.n5385 GND.n4963 585
R11043 GND.n5387 GND.n4025 585
R11044 GND.n7921 GND.n4025 585
R11045 GND.n5389 GND.n5388 585
R11046 GND.n5388 GND.n4968 585
R11047 GND.n5390 GND.n4015 585
R11048 GND.n7927 GND.n4015 585
R11049 GND.n5392 GND.n5391 585
R11050 GND.n5391 GND.n4973 585
R11051 GND.n5393 GND.n4005 585
R11052 GND.n7933 GND.n4005 585
R11053 GND.n5395 GND.n5394 585
R11054 GND.n5394 GND.n4978 585
R11055 GND.n5396 GND.n3995 585
R11056 GND.n7939 GND.n3995 585
R11057 GND.n5399 GND.n5398 585
R11058 GND.n5398 GND.n5397 585
R11059 GND.n5400 GND.n3985 585
R11060 GND.n7945 GND.n3985 585
R11061 GND.n5402 GND.n5401 585
R11062 GND.n5401 GND.n4987 585
R11063 GND.n5403 GND.n3975 585
R11064 GND.n7951 GND.n3975 585
R11065 GND.n5404 GND.n4992 585
R11066 GND.n5430 GND.n4992 585
R11067 GND.n5405 GND.n3965 585
R11068 GND.n7957 GND.n3965 585
R11069 GND.n5407 GND.n5406 585
R11070 GND.n5406 GND.n4997 585
R11071 GND.n5408 GND.n3955 585
R11072 GND.n7963 GND.n3955 585
R11073 GND.n5410 GND.n5409 585
R11074 GND.n5411 GND.n5410 585
R11075 GND.n5003 GND.n3945 585
R11076 GND.n7969 GND.n3945 585
R11077 GND.n5364 GND.n5363 585
R11078 GND.n5363 GND.n5362 585
R11079 GND.n5005 GND.n3935 585
R11080 GND.n7975 GND.n3935 585
R11081 GND.n5350 GND.n5349 585
R11082 GND.n5351 GND.n5350 585
R11083 GND.n5012 GND.n3925 585
R11084 GND.n7981 GND.n3925 585
R11085 GND.n5345 GND.n5344 585
R11086 GND.n5344 GND.n5343 585
R11087 GND.n5014 GND.n3915 585
R11088 GND.n7987 GND.n3915 585
R11089 GND.n5331 GND.n5330 585
R11090 GND.n5332 GND.n5331 585
R11091 GND.n5021 GND.n3905 585
R11092 GND.n7993 GND.n3905 585
R11093 GND.n5326 GND.n5325 585
R11094 GND.n5325 GND.n5324 585
R11095 GND.n5029 GND.n3894 585
R11096 GND.n7999 GND.n3894 585
R11097 GND.n5028 GND.n5025 585
R11098 GND.n5025 GND.n5024 585
R11099 GND.n5023 GND.n3864 585
R11100 GND.n8005 GND.n3864 585
R11101 GND.n8054 GND.n8053 585
R11102 GND.n8052 GND.n3863 585
R11103 GND.n8051 GND.n3862 585
R11104 GND.n8056 GND.n3862 585
R11105 GND.n8050 GND.n8049 585
R11106 GND.n8048 GND.n8047 585
R11107 GND.n8046 GND.n8045 585
R11108 GND.n8044 GND.n3871 585
R11109 GND.n3873 GND.n3872 585
R11110 GND.n8041 GND.n8038 585
R11111 GND.n8040 GND.n8039 585
R11112 GND.n8036 GND.n8033 585
R11113 GND.n8035 GND.n8034 585
R11114 GND.n8031 GND.n8028 585
R11115 GND.n8030 GND.n8029 585
R11116 GND.n8026 GND.n8023 585
R11117 GND.n8025 GND.n8024 585
R11118 GND.n8021 GND.n8018 585
R11119 GND.n8020 GND.n8019 585
R11120 GND.n8016 GND.n8012 585
R11121 GND.n8011 GND.n3875 585
R11122 GND.n3877 GND.n3876 585
R11123 GND.n8009 GND.n3878 585
R11124 GND.n8008 GND.n8007 585
R11125 GND.n5868 GND.n4844 585
R11126 GND.n5871 GND.n5870 585
R11127 GND.n5867 GND.n4843 585
R11128 GND.n5865 GND.n5864 585
R11129 GND.n5862 GND.n5859 585
R11130 GND.n5857 GND.n5856 585
R11131 GND.n5855 GND.n5854 585
R11132 GND.n5852 GND.n5851 585
R11133 GND.n5850 GND.n5849 585
R11134 GND.n5847 GND.n5846 585
R11135 GND.n5845 GND.n5844 585
R11136 GND.n5842 GND.n5841 585
R11137 GND.n5840 GND.n5839 585
R11138 GND.n5837 GND.n5836 585
R11139 GND.n5835 GND.n4841 585
R11140 GND.n5833 GND.n5832 585
R11141 GND.n5831 GND.n5830 585
R11142 GND.n5829 GND.n5828 585
R11143 GND.n5827 GND.n4846 585
R11144 GND.n5825 GND.n5824 585
R11145 GND.n4848 GND.n4847 585
R11146 GND.n5819 GND.n5818 585
R11147 GND.n5816 GND.n5815 585
R11148 GND.n5816 GND.n4376 585
R11149 GND.n4832 GND.n4369 585
R11150 GND.n7738 GND.n4369 585
R11151 GND.n4354 GND.n4353 585
R11152 GND.n5809 GND.n4354 585
R11153 GND.n7746 GND.n7745 585
R11154 GND.n7745 GND.n7744 585
R11155 GND.n7747 GND.n4348 585
R11156 GND.n5793 GND.n4348 585
R11157 GND.n7749 GND.n7748 585
R11158 GND.n7750 GND.n7749 585
R11159 GND.n4335 GND.n4334 585
R11160 GND.n5801 GND.n4335 585
R11161 GND.n7758 GND.n7757 585
R11162 GND.n7757 GND.n7756 585
R11163 GND.n7759 GND.n4329 585
R11164 GND.n4872 GND.n4329 585
R11165 GND.n7761 GND.n7760 585
R11166 GND.n7762 GND.n7761 585
R11167 GND.n4315 GND.n4314 585
R11168 GND.n4877 GND.n4315 585
R11169 GND.n7770 GND.n7769 585
R11170 GND.n7769 GND.n7768 585
R11171 GND.n7771 GND.n4297 585
R11172 GND.n4882 GND.n4297 585
R11173 GND.n7773 GND.n7772 585
R11174 GND.n7774 GND.n7773 585
R11175 GND.n4298 GND.n4296 585
R11176 GND.n5743 GND.n4296 585
R11177 GND.n4308 GND.n4282 585
R11178 GND.n7780 GND.n4282 585
R11179 GND.n4307 GND.n4306 585
R11180 GND.n4306 GND.n4272 585
R11181 GND.n4305 GND.n4304 585
R11182 GND.n4305 GND.n4271 585
R11183 GND.n4300 GND.n4265 585
R11184 GND.n7793 GND.n4265 585
R11185 GND.n4250 GND.n4249 585
R11186 GND.n4888 GND.n4250 585
R11187 GND.n7801 GND.n7800 585
R11188 GND.n7800 GND.n7799 585
R11189 GND.n7802 GND.n4244 585
R11190 GND.n5710 GND.n4244 585
R11191 GND.n7804 GND.n7803 585
R11192 GND.n7805 GND.n7804 585
R11193 GND.n4232 GND.n4231 585
R11194 GND.n5631 GND.n4232 585
R11195 GND.n7813 GND.n7812 585
R11196 GND.n7812 GND.n7811 585
R11197 GND.n7814 GND.n4226 585
R11198 GND.n4905 GND.n4226 585
R11199 GND.n7816 GND.n7815 585
R11200 GND.n7817 GND.n7816 585
R11201 GND.n4212 GND.n4211 585
R11202 GND.n4910 GND.n4212 585
R11203 GND.n7825 GND.n7824 585
R11204 GND.n7824 GND.n7823 585
R11205 GND.n7826 GND.n4194 585
R11206 GND.n4915 GND.n4194 585
R11207 GND.n7828 GND.n7827 585
R11208 GND.n7829 GND.n7828 585
R11209 GND.n4195 GND.n4193 585
R11210 GND.n5646 GND.n4193 585
R11211 GND.n4205 GND.n4180 585
R11212 GND.n7835 GND.n4180 585
R11213 GND.n4204 GND.n4203 585
R11214 GND.n4203 GND.n4170 585
R11215 GND.n4202 GND.n4201 585
R11216 GND.n4202 GND.n4169 585
R11217 GND.n4197 GND.n4163 585
R11218 GND.n7848 GND.n4163 585
R11219 GND.n4148 GND.n4147 585
R11220 GND.n4922 GND.n4148 585
R11221 GND.n7856 GND.n7855 585
R11222 GND.n7855 GND.n7854 585
R11223 GND.n7857 GND.n4142 585
R11224 GND.n5607 GND.n4142 585
R11225 GND.n7859 GND.n7858 585
R11226 GND.n7860 GND.n7859 585
R11227 GND.n4128 GND.n4127 585
R11228 GND.n4932 GND.n4128 585
R11229 GND.n7868 GND.n7867 585
R11230 GND.n7867 GND.n7866 585
R11231 GND.n7869 GND.n4122 585
R11232 GND.n4937 GND.n4122 585
R11233 GND.n7871 GND.n7870 585
R11234 GND.n7872 GND.n7871 585
R11235 GND.n4108 GND.n4107 585
R11236 GND.n4942 GND.n4108 585
R11237 GND.n7880 GND.n7879 585
R11238 GND.n7879 GND.n7878 585
R11239 GND.n7881 GND.n4090 585
R11240 GND.n4947 GND.n4090 585
R11241 GND.n7883 GND.n7882 585
R11242 GND.n7884 GND.n7883 585
R11243 GND.n4091 GND.n4089 585
R11244 GND.n5542 GND.n4089 585
R11245 GND.n4101 GND.n4075 585
R11246 GND.n7890 GND.n4075 585
R11247 GND.n4100 GND.n4099 585
R11248 GND.n4099 GND.n4065 585
R11249 GND.n4098 GND.n4097 585
R11250 GND.n4098 GND.n4064 585
R11251 GND.n4093 GND.n4058 585
R11252 GND.n7903 GND.n4058 585
R11253 GND.n4043 GND.n4042 585
R11254 GND.n4953 GND.n4043 585
R11255 GND.n7911 GND.n7910 585
R11256 GND.n7910 GND.n7909 585
R11257 GND.n7912 GND.n4037 585
R11258 GND.n5504 GND.n4037 585
R11259 GND.n7914 GND.n7913 585
R11260 GND.n7915 GND.n7914 585
R11261 GND.n4023 GND.n4022 585
R11262 GND.n4963 GND.n4023 585
R11263 GND.n7923 GND.n7922 585
R11264 GND.n7922 GND.n7921 585
R11265 GND.n7924 GND.n4017 585
R11266 GND.n4968 GND.n4017 585
R11267 GND.n7926 GND.n7925 585
R11268 GND.n7927 GND.n7926 585
R11269 GND.n4003 GND.n4002 585
R11270 GND.n4973 GND.n4003 585
R11271 GND.n7935 GND.n7934 585
R11272 GND.n7934 GND.n7933 585
R11273 GND.n7936 GND.n3997 585
R11274 GND.n4978 GND.n3997 585
R11275 GND.n7938 GND.n7937 585
R11276 GND.n7939 GND.n7938 585
R11277 GND.n3983 GND.n3982 585
R11278 GND.n5397 GND.n3983 585
R11279 GND.n7947 GND.n7946 585
R11280 GND.n7946 GND.n7945 585
R11281 GND.n7948 GND.n3977 585
R11282 GND.n4987 GND.n3977 585
R11283 GND.n7950 GND.n7949 585
R11284 GND.n7951 GND.n7950 585
R11285 GND.n3963 GND.n3962 585
R11286 GND.n5430 GND.n3963 585
R11287 GND.n7959 GND.n7958 585
R11288 GND.n7958 GND.n7957 585
R11289 GND.n7960 GND.n3957 585
R11290 GND.n4997 GND.n3957 585
R11291 GND.n7962 GND.n7961 585
R11292 GND.n7963 GND.n7962 585
R11293 GND.n3943 GND.n3942 585
R11294 GND.n5411 GND.n3943 585
R11295 GND.n7971 GND.n7970 585
R11296 GND.n7970 GND.n7969 585
R11297 GND.n7972 GND.n3937 585
R11298 GND.n5362 GND.n3937 585
R11299 GND.n7974 GND.n7973 585
R11300 GND.n7975 GND.n7974 585
R11301 GND.n3923 GND.n3922 585
R11302 GND.n5351 GND.n3923 585
R11303 GND.n7983 GND.n7982 585
R11304 GND.n7982 GND.n7981 585
R11305 GND.n7984 GND.n3917 585
R11306 GND.n5343 GND.n3917 585
R11307 GND.n7986 GND.n7985 585
R11308 GND.n7987 GND.n7986 585
R11309 GND.n3904 GND.n3903 585
R11310 GND.n5332 GND.n3904 585
R11311 GND.n7995 GND.n7994 585
R11312 GND.n7994 GND.n7993 585
R11313 GND.n7996 GND.n3896 585
R11314 GND.n5324 GND.n3896 585
R11315 GND.n7998 GND.n7997 585
R11316 GND.n7999 GND.n7998 585
R11317 GND.n3897 GND.n3879 585
R11318 GND.n5024 GND.n3879 585
R11319 GND.n8006 GND.n3880 585
R11320 GND.n8006 GND.n8005 585
R11321 GND.n4726 GND.n4725 585
R11322 GND.n4726 GND.n4527 585
R11323 GND.n4724 GND.n4723 585
R11324 GND.n4723 GND.n4722 585
R11325 GND.n4513 GND.n4512 585
R11326 GND.n4516 GND.n4513 585
R11327 GND.n7667 GND.n7666 585
R11328 GND.n7666 GND.n7665 585
R11329 GND.n7668 GND.n4507 585
R11330 GND.n4514 GND.n4507 585
R11331 GND.n7670 GND.n7669 585
R11332 GND.n7671 GND.n7670 585
R11333 GND.n4511 GND.n4506 585
R11334 GND.n4506 GND.n4451 585
R11335 GND.n4510 GND.n4450 585
R11336 GND.n7677 GND.n4450 585
R11337 GND.n4509 GND.n4508 585
R11338 GND.n4508 GND.n4449 585
R11339 GND.n4439 GND.n4438 585
R11340 GND.n4498 GND.n4439 585
R11341 GND.n7686 GND.n7685 585
R11342 GND.n7685 GND.n7684 585
R11343 GND.n7687 GND.n4436 585
R11344 GND.n4440 GND.n4436 585
R11345 GND.n7689 GND.n7688 585
R11346 GND.n7690 GND.n7689 585
R11347 GND.n4437 GND.n4435 585
R11348 GND.n4435 GND.n4432 585
R11349 GND.n4488 GND.n4487 585
R11350 GND.n4489 GND.n4488 585
R11351 GND.n4421 GND.n4420 585
R11352 GND.n4424 GND.n4421 585
R11353 GND.n7700 GND.n7699 585
R11354 GND.n7699 GND.n7698 585
R11355 GND.n7701 GND.n4418 585
R11356 GND.n4422 GND.n4418 585
R11357 GND.n7703 GND.n7702 585
R11358 GND.n7704 GND.n7703 585
R11359 GND.n4419 GND.n4417 585
R11360 GND.n4417 GND.n4414 585
R11361 GND.n4475 GND.n4474 585
R11362 GND.n4476 GND.n4475 585
R11363 GND.n4403 GND.n4402 585
R11364 GND.n4406 GND.n4403 585
R11365 GND.n7714 GND.n7713 585
R11366 GND.n7713 GND.n7712 585
R11367 GND.n7715 GND.n4400 585
R11368 GND.n4404 GND.n4400 585
R11369 GND.n7717 GND.n7716 585
R11370 GND.n7718 GND.n7717 585
R11371 GND.n4401 GND.n4399 585
R11372 GND.n4399 GND.n4396 585
R11373 GND.n4462 GND.n4461 585
R11374 GND.n4463 GND.n4462 585
R11375 GND.n4381 GND.n4380 585
R11376 GND.n4384 GND.n4381 585
R11377 GND.n7728 GND.n7727 585
R11378 GND.n7727 GND.n7726 585
R11379 GND.n7729 GND.n4378 585
R11380 GND.n4382 GND.n4378 585
R11381 GND.n7731 GND.n7730 585
R11382 GND.n7732 GND.n7731 585
R11383 GND.n4379 GND.n4377 585
R11384 GND.n4377 GND.n4368 585
R11385 GND.n4859 GND.n4366 585
R11386 GND.n7738 GND.n4366 585
R11387 GND.n4861 GND.n4860 585
R11388 GND.n4860 GND.n4365 585
R11389 GND.n4862 GND.n4858 585
R11390 GND.n4858 GND.n4357 585
R11391 GND.n4864 GND.n4863 585
R11392 GND.n4864 GND.n4355 585
R11393 GND.n4865 GND.n4857 585
R11394 GND.n5792 GND.n4865 585
R11395 GND.n5796 GND.n5795 585
R11396 GND.n5795 GND.n5794 585
R11397 GND.n5797 GND.n4855 585
R11398 GND.n4855 GND.n4346 585
R11399 GND.n5799 GND.n5798 585
R11400 GND.n5800 GND.n5799 585
R11401 GND.n4856 GND.n4854 585
R11402 GND.n4854 GND.n4338 585
R11403 GND.n5775 GND.n4874 585
R11404 GND.n4874 GND.n4336 585
R11405 GND.n5777 GND.n5776 585
R11406 GND.n5778 GND.n5777 585
R11407 GND.n5774 GND.n4873 585
R11408 GND.n4873 GND.n4328 585
R11409 GND.n5773 GND.n5772 585
R11410 GND.n5772 GND.n4326 585
R11411 GND.n5771 GND.n4875 585
R11412 GND.n5771 GND.n5770 585
R11413 GND.n5757 GND.n4876 585
R11414 GND.n4876 GND.n4318 585
R11415 GND.n5758 GND.n4884 585
R11416 GND.n4884 GND.n4316 585
R11417 GND.n5760 GND.n5759 585
R11418 GND.n5761 GND.n5760 585
R11419 GND.n5756 GND.n4883 585
R11420 GND.n4883 GND.n4295 585
R11421 GND.n5755 GND.n5754 585
R11422 GND.n5754 GND.n4293 585
R11423 GND.n5753 GND.n4885 585
R11424 GND.n5753 GND.n5752 585
R11425 GND.n4277 GND.n4276 585
R11426 GND.n4281 GND.n4277 585
R11427 GND.n7783 GND.n7782 585
R11428 GND.n7782 GND.n7781 585
R11429 GND.n7784 GND.n4274 585
R11430 GND.n4278 GND.n4274 585
R11431 GND.n7786 GND.n7785 585
R11432 GND.n7787 GND.n7786 585
R11433 GND.n4275 GND.n4273 585
R11434 GND.n4273 GND.n4264 585
R11435 GND.n5701 GND.n4262 585
R11436 GND.n7793 GND.n4262 585
R11437 GND.n5703 GND.n5702 585
R11438 GND.n5703 GND.n4261 585
R11439 GND.n5705 GND.n5704 585
R11440 GND.n5704 GND.n4253 585
R11441 GND.n5706 GND.n4896 585
R11442 GND.n4896 GND.n4251 585
R11443 GND.n5708 GND.n5707 585
R11444 GND.n5709 GND.n5708 585
R11445 GND.n5700 GND.n4895 585
R11446 GND.n4895 GND.n4893 585
R11447 GND.n5699 GND.n5698 585
R11448 GND.n5698 GND.n5697 585
R11449 GND.n4898 GND.n4897 585
R11450 GND.n4899 GND.n4898 585
R11451 GND.n5679 GND.n5678 585
R11452 GND.n5678 GND.n4235 585
R11453 GND.n5680 GND.n4907 585
R11454 GND.n4907 GND.n4233 585
R11455 GND.n5682 GND.n5681 585
R11456 GND.n5683 GND.n5682 585
R11457 GND.n5677 GND.n4906 585
R11458 GND.n4906 GND.n4225 585
R11459 GND.n5676 GND.n5675 585
R11460 GND.n5675 GND.n4223 585
R11461 GND.n5674 GND.n4908 585
R11462 GND.n5674 GND.n5673 585
R11463 GND.n5660 GND.n4909 585
R11464 GND.n4909 GND.n4215 585
R11465 GND.n5661 GND.n4918 585
R11466 GND.n4918 GND.n4213 585
R11467 GND.n5663 GND.n5662 585
R11468 GND.n5664 GND.n5663 585
R11469 GND.n5659 GND.n4917 585
R11470 GND.n4917 GND.n4916 585
R11471 GND.n5658 GND.n5657 585
R11472 GND.n5657 GND.n4191 585
R11473 GND.n5656 GND.n4919 585
R11474 GND.n5656 GND.n5655 585
R11475 GND.n4175 GND.n4174 585
R11476 GND.n4179 GND.n4175 585
R11477 GND.n7838 GND.n7837 585
R11478 GND.n7837 GND.n7836 585
R11479 GND.n7839 GND.n4172 585
R11480 GND.n4176 GND.n4172 585
R11481 GND.n7841 GND.n7840 585
R11482 GND.n7842 GND.n7841 585
R11483 GND.n4173 GND.n4171 585
R11484 GND.n4171 GND.n4162 585
R11485 GND.n5598 GND.n4160 585
R11486 GND.n7848 GND.n4160 585
R11487 GND.n5600 GND.n5599 585
R11488 GND.n5600 GND.n4159 585
R11489 GND.n5602 GND.n5601 585
R11490 GND.n5601 GND.n4151 585
R11491 GND.n5603 GND.n4929 585
R11492 GND.n4929 GND.n4149 585
R11493 GND.n5605 GND.n5604 585
R11494 GND.n5606 GND.n5605 585
R11495 GND.n5597 GND.n4928 585
R11496 GND.n4928 GND.n4141 585
R11497 GND.n5596 GND.n5595 585
R11498 GND.n5595 GND.n4139 585
R11499 GND.n5594 GND.n4930 585
R11500 GND.n5594 GND.n5593 585
R11501 GND.n5574 GND.n4931 585
R11502 GND.n4931 GND.n4131 585
R11503 GND.n5575 GND.n4939 585
R11504 GND.n4939 GND.n4129 585
R11505 GND.n5577 GND.n5576 585
R11506 GND.n5578 GND.n5577 585
R11507 GND.n5573 GND.n4938 585
R11508 GND.n4938 GND.n4121 585
R11509 GND.n5572 GND.n5571 585
R11510 GND.n5571 GND.n4119 585
R11511 GND.n5570 GND.n4940 585
R11512 GND.n5570 GND.n5569 585
R11513 GND.n5556 GND.n4941 585
R11514 GND.n4941 GND.n4111 585
R11515 GND.n5557 GND.n4949 585
R11516 GND.n4949 GND.n4109 585
R11517 GND.n5559 GND.n5558 585
R11518 GND.n5560 GND.n5559 585
R11519 GND.n5555 GND.n4948 585
R11520 GND.n4948 GND.n4088 585
R11521 GND.n5554 GND.n5553 585
R11522 GND.n5553 GND.n4086 585
R11523 GND.n5552 GND.n4950 585
R11524 GND.n5552 GND.n5551 585
R11525 GND.n4070 GND.n4069 585
R11526 GND.n4074 GND.n4070 585
R11527 GND.n7893 GND.n7892 585
R11528 GND.n7892 GND.n7891 585
R11529 GND.n7894 GND.n4067 585
R11530 GND.n4071 GND.n4067 585
R11531 GND.n7896 GND.n7895 585
R11532 GND.n7897 GND.n7896 585
R11533 GND.n4068 GND.n4066 585
R11534 GND.n4066 GND.n4057 585
R11535 GND.n5495 GND.n4055 585
R11536 GND.n7903 GND.n4055 585
R11537 GND.n5497 GND.n5496 585
R11538 GND.n5497 GND.n4054 585
R11539 GND.n5499 GND.n5498 585
R11540 GND.n5498 GND.n4046 585
R11541 GND.n5500 GND.n4960 585
R11542 GND.n4960 GND.n4044 585
R11543 GND.n5502 GND.n5501 585
R11544 GND.n5503 GND.n5502 585
R11545 GND.n5494 GND.n4959 585
R11546 GND.n4959 GND.n4036 585
R11547 GND.n5493 GND.n5492 585
R11548 GND.n5492 GND.n4034 585
R11549 GND.n5491 GND.n4961 585
R11550 GND.n5491 GND.n5490 585
R11551 GND.n5471 GND.n4962 585
R11552 GND.n4962 GND.n4026 585
R11553 GND.n5472 GND.n4970 585
R11554 GND.n4970 GND.n4024 585
R11555 GND.n5474 GND.n5473 585
R11556 GND.n5475 GND.n5474 585
R11557 GND.n5470 GND.n4969 585
R11558 GND.n4969 GND.n4016 585
R11559 GND.n5469 GND.n5468 585
R11560 GND.n5468 GND.n4014 585
R11561 GND.n5467 GND.n4971 585
R11562 GND.n5467 GND.n5466 585
R11563 GND.n5453 GND.n4972 585
R11564 GND.n4972 GND.n4006 585
R11565 GND.n5454 GND.n4980 585
R11566 GND.n4980 GND.n4004 585
R11567 GND.n5456 GND.n5455 585
R11568 GND.n5457 GND.n5456 585
R11569 GND.n5452 GND.n4979 585
R11570 GND.n4979 GND.n3996 585
R11571 GND.n5451 GND.n5450 585
R11572 GND.n5450 GND.n3994 585
R11573 GND.n5449 GND.n4981 585
R11574 GND.n5449 GND.n5448 585
R11575 GND.n5435 GND.n4982 585
R11576 GND.n4982 GND.n3986 585
R11577 GND.n5436 GND.n4989 585
R11578 GND.n4989 GND.n3984 585
R11579 GND.n5438 GND.n5437 585
R11580 GND.n5439 GND.n5438 585
R11581 GND.n5434 GND.n4988 585
R11582 GND.n4988 GND.n3976 585
R11583 GND.n5433 GND.n5432 585
R11584 GND.n5432 GND.n3974 585
R11585 GND.n5431 GND.n4990 585
R11586 GND.n5431 GND.n5430 585
R11587 GND.n5417 GND.n4991 585
R11588 GND.n4991 GND.n3966 585
R11589 GND.n5418 GND.n4999 585
R11590 GND.n4999 GND.n3964 585
R11591 GND.n5420 GND.n5419 585
R11592 GND.n5421 GND.n5420 585
R11593 GND.n5416 GND.n4998 585
R11594 GND.n4998 GND.n3956 585
R11595 GND.n5415 GND.n5414 585
R11596 GND.n5414 GND.n3954 585
R11597 GND.n5413 GND.n5000 585
R11598 GND.n5413 GND.n5412 585
R11599 GND.n5357 GND.n5001 585
R11600 GND.n5001 GND.n3946 585
R11601 GND.n5358 GND.n5008 585
R11602 GND.n5008 GND.n3944 585
R11603 GND.n5360 GND.n5359 585
R11604 GND.n5361 GND.n5360 585
R11605 GND.n5356 GND.n5007 585
R11606 GND.n5007 GND.n3936 585
R11607 GND.n5355 GND.n5354 585
R11608 GND.n5354 GND.n3934 585
R11609 GND.n5353 GND.n5009 585
R11610 GND.n5353 GND.n5352 585
R11611 GND.n5338 GND.n5010 585
R11612 GND.n5010 GND.n3926 585
R11613 GND.n5339 GND.n5017 585
R11614 GND.n5017 GND.n3924 585
R11615 GND.n5341 GND.n5340 585
R11616 GND.n5342 GND.n5341 585
R11617 GND.n5337 GND.n5016 585
R11618 GND.n5016 GND.n3916 585
R11619 GND.n5336 GND.n5335 585
R11620 GND.n5335 GND.n3914 585
R11621 GND.n5334 GND.n5018 585
R11622 GND.n5334 GND.n5333 585
R11623 GND.n5320 GND.n5019 585
R11624 GND.n5019 GND.n3906 585
R11625 GND.n5322 GND.n5321 585
R11626 GND.n5323 GND.n5322 585
R11627 GND.n5319 GND.n5032 585
R11628 GND.n5032 GND.n5030 585
R11629 GND.n5318 GND.n5317 585
R11630 GND.n5317 GND.n3895 585
R11631 GND.n5316 GND.n5033 585
R11632 GND.n5316 GND.n3893 585
R11633 GND.n5315 GND.n5314 585
R11634 GND.n5315 GND.n3884 585
R11635 GND.n5313 GND.n3883 585
R11636 GND.n8005 GND.n3883 585
R11637 GND.n5312 GND.n5311 585
R11638 GND.n5311 GND.n3882 585
R11639 GND.n5310 GND.n5034 585
R11640 GND.n5310 GND.n3861 585
R11641 GND.n5309 GND.n5308 585
R11642 GND.n5309 GND.n3850 585
R11643 GND.n5307 GND.n5306 585
R11644 GND.n5306 GND.n5305 585
R11645 GND.n3839 GND.n3838 585
R11646 GND.n3842 GND.n3839 585
R11647 GND.n8066 GND.n8065 585
R11648 GND.n8065 GND.n8064 585
R11649 GND.n8067 GND.n3836 585
R11650 GND.n3840 GND.n3836 585
R11651 GND.n8069 GND.n8068 585
R11652 GND.n8070 GND.n8069 585
R11653 GND.n3837 GND.n3835 585
R11654 GND.n3835 GND.n3832 585
R11655 GND.n5252 GND.n5251 585
R11656 GND.n5253 GND.n5252 585
R11657 GND.n3821 GND.n3820 585
R11658 GND.n3824 GND.n3821 585
R11659 GND.n8080 GND.n8079 585
R11660 GND.n8079 GND.n8078 585
R11661 GND.n8081 GND.n3818 585
R11662 GND.n3822 GND.n3818 585
R11663 GND.n8083 GND.n8082 585
R11664 GND.n8084 GND.n8083 585
R11665 GND.n3819 GND.n3817 585
R11666 GND.n3817 GND.n3814 585
R11667 GND.n5239 GND.n5238 585
R11668 GND.n5240 GND.n5239 585
R11669 GND.n3803 GND.n3802 585
R11670 GND.n3806 GND.n3803 585
R11671 GND.n8094 GND.n8093 585
R11672 GND.n8093 GND.n8092 585
R11673 GND.n8095 GND.n3800 585
R11674 GND.n3804 GND.n3800 585
R11675 GND.n8097 GND.n8096 585
R11676 GND.n8098 GND.n8097 585
R11677 GND.n3801 GND.n3799 585
R11678 GND.n3799 GND.n3796 585
R11679 GND.n5226 GND.n5225 585
R11680 GND.n5227 GND.n5226 585
R11681 GND.n3786 GND.n3785 585
R11682 GND.n3788 GND.n3786 585
R11683 GND.n8108 GND.n8107 585
R11684 GND.n8107 GND.n8106 585
R11685 GND.n8109 GND.n3783 585
R11686 GND.n3783 GND.t64 585
R11687 GND.n8111 GND.n8110 585
R11688 GND.n8112 GND.n8111 585
R11689 GND.n3784 GND.n3782 585
R11690 GND.n3782 GND.n3780 585
R11691 GND.n5213 GND.n5212 585
R11692 GND.n5214 GND.n5213 585
R11693 GND.n3769 GND.n3768 585
R11694 GND.n3772 GND.n3769 585
R11695 GND.n8122 GND.n8121 585
R11696 GND.n8121 GND.n8120 585
R11697 GND.n8123 GND.n3753 585
R11698 GND.n3753 GND.n3751 585
R11699 GND.n8125 GND.n8124 585
R11700 GND.n8126 GND.n8125 585
R11701 GND.n5079 GND.n3752 585
R11702 GND.n5082 GND.n5081 585
R11703 GND.n5083 GND.n5078 585
R11704 GND.n5078 GND.n3749 585
R11705 GND.n5085 GND.n5084 585
R11706 GND.n5087 GND.n5077 585
R11707 GND.n5090 GND.n5089 585
R11708 GND.n5091 GND.n5076 585
R11709 GND.n5093 GND.n5092 585
R11710 GND.n5095 GND.n5075 585
R11711 GND.n5098 GND.n5097 585
R11712 GND.n5099 GND.n5074 585
R11713 GND.n5101 GND.n5100 585
R11714 GND.n5103 GND.n5073 585
R11715 GND.n5106 GND.n5105 585
R11716 GND.n5107 GND.n5072 585
R11717 GND.n5109 GND.n5108 585
R11718 GND.n5111 GND.n5071 585
R11719 GND.n5114 GND.n5113 585
R11720 GND.n5115 GND.n5070 585
R11721 GND.n5117 GND.n5116 585
R11722 GND.n5119 GND.n5069 585
R11723 GND.n5122 GND.n5121 585
R11724 GND.n5123 GND.n5068 585
R11725 GND.n5125 GND.n5124 585
R11726 GND.n5127 GND.n5067 585
R11727 GND.n5130 GND.n5129 585
R11728 GND.n5131 GND.n5064 585
R11729 GND.n5134 GND.n5133 585
R11730 GND.n5136 GND.n5063 585
R11731 GND.n5137 GND.n5062 585
R11732 GND.n5140 GND.n5139 585
R11733 GND.n5141 GND.n5061 585
R11734 GND.n5141 GND.n5059 585
R11735 GND.n5143 GND.n5142 585
R11736 GND.n5145 GND.n5058 585
R11737 GND.n5148 GND.n5147 585
R11738 GND.n5149 GND.n5055 585
R11739 GND.n5152 GND.n5151 585
R11740 GND.n5154 GND.n5054 585
R11741 GND.n5157 GND.n5156 585
R11742 GND.n5158 GND.n5053 585
R11743 GND.n5160 GND.n5159 585
R11744 GND.n5162 GND.n5052 585
R11745 GND.n5165 GND.n5164 585
R11746 GND.n5166 GND.n5051 585
R11747 GND.n5168 GND.n5167 585
R11748 GND.n5170 GND.n5050 585
R11749 GND.n5173 GND.n5172 585
R11750 GND.n5174 GND.n5049 585
R11751 GND.n5176 GND.n5175 585
R11752 GND.n5178 GND.n5048 585
R11753 GND.n5181 GND.n5180 585
R11754 GND.n5182 GND.n5047 585
R11755 GND.n5184 GND.n5183 585
R11756 GND.n5186 GND.n5046 585
R11757 GND.n5189 GND.n5188 585
R11758 GND.n5190 GND.n5045 585
R11759 GND.n5192 GND.n5191 585
R11760 GND.n5194 GND.n5044 585
R11761 GND.n5197 GND.n5196 585
R11762 GND.n5198 GND.n5043 585
R11763 GND.n5200 GND.n5199 585
R11764 GND.n5202 GND.n5042 585
R11765 GND.n5204 GND.n5203 585
R11766 GND.n5203 GND.n3749 585
R11767 GND.n4718 GND.n4717 585
R11768 GND.n4716 GND.n4715 585
R11769 GND.n4714 GND.n4713 585
R11770 GND.n4712 GND.n4711 585
R11771 GND.n4710 GND.n4709 585
R11772 GND.n4708 GND.n4707 585
R11773 GND.n4706 GND.n4705 585
R11774 GND.n4704 GND.n4703 585
R11775 GND.n4702 GND.n4701 585
R11776 GND.n4700 GND.n4699 585
R11777 GND.n4698 GND.n4697 585
R11778 GND.n4696 GND.n4695 585
R11779 GND.n4694 GND.n4693 585
R11780 GND.n4692 GND.n4691 585
R11781 GND.n4690 GND.n4689 585
R11782 GND.n4688 GND.n4687 585
R11783 GND.n4686 GND.n4685 585
R11784 GND.n4684 GND.n4683 585
R11785 GND.n4682 GND.n4681 585
R11786 GND.n4680 GND.n4679 585
R11787 GND.n4678 GND.n4677 585
R11788 GND.n4676 GND.n4675 585
R11789 GND.n4674 GND.n4673 585
R11790 GND.n4672 GND.n4671 585
R11791 GND.n4670 GND.n4669 585
R11792 GND.n4668 GND.n4667 585
R11793 GND.n4666 GND.n4665 585
R11794 GND.n4663 GND.n4662 585
R11795 GND.n4661 GND.n4660 585
R11796 GND.n4659 GND.n4658 585
R11797 GND.n4657 GND.n4634 585
R11798 GND.n4789 GND.n4788 585
R11799 GND.n4787 GND.n4786 585
R11800 GND.n4785 GND.n4784 585
R11801 GND.n4783 GND.n4782 585
R11802 GND.n4780 GND.n4779 585
R11803 GND.n4778 GND.n4777 585
R11804 GND.n4776 GND.n4775 585
R11805 GND.n4774 GND.n4773 585
R11806 GND.n4772 GND.n4771 585
R11807 GND.n4770 GND.n4769 585
R11808 GND.n4768 GND.n4767 585
R11809 GND.n4766 GND.n4765 585
R11810 GND.n4764 GND.n4763 585
R11811 GND.n4762 GND.n4761 585
R11812 GND.n4760 GND.n4759 585
R11813 GND.n4758 GND.n4757 585
R11814 GND.n4756 GND.n4755 585
R11815 GND.n4754 GND.n4753 585
R11816 GND.n4752 GND.n4751 585
R11817 GND.n4750 GND.n4749 585
R11818 GND.n4748 GND.n4747 585
R11819 GND.n4746 GND.n4745 585
R11820 GND.n4744 GND.n4743 585
R11821 GND.n4742 GND.n4741 585
R11822 GND.n4740 GND.n4739 585
R11823 GND.n4738 GND.n4737 585
R11824 GND.n4736 GND.n4735 585
R11825 GND.n4734 GND.n4733 585
R11826 GND.n4732 GND.n4731 585
R11827 GND.n4730 GND.n4729 585
R11828 GND.n4728 GND.n4727 585
R11829 GND.n4719 GND.n4652 585
R11830 GND.n4652 GND.n4527 585
R11831 GND.n4721 GND.n4720 585
R11832 GND.n4722 GND.n4721 585
R11833 GND.n4654 GND.n4651 585
R11834 GND.n4651 GND.n4516 585
R11835 GND.n4653 GND.n4515 585
R11836 GND.n7665 GND.n4515 585
R11837 GND.n4503 GND.n4502 585
R11838 GND.n4514 GND.n4503 585
R11839 GND.n7673 GND.n7672 585
R11840 GND.n7672 GND.n7671 585
R11841 GND.n7674 GND.n4453 585
R11842 GND.n4453 GND.n4451 585
R11843 GND.n7676 GND.n7675 585
R11844 GND.n7677 GND.n7676 585
R11845 GND.n4501 GND.n4452 585
R11846 GND.n4452 GND.n4449 585
R11847 GND.n4500 GND.n4499 585
R11848 GND.n4499 GND.n4498 585
R11849 GND.n4496 GND.n4441 585
R11850 GND.n7684 GND.n4441 585
R11851 GND.n4495 GND.n4494 585
R11852 GND.n4494 GND.n4440 585
R11853 GND.n4493 GND.n4433 585
R11854 GND.n7690 GND.n4433 585
R11855 GND.n4492 GND.n4491 585
R11856 GND.n4491 GND.n4432 585
R11857 GND.n4490 GND.n4454 585
R11858 GND.n4490 GND.n4489 585
R11859 GND.n4485 GND.n4484 585
R11860 GND.n4485 GND.n4424 585
R11861 GND.n4483 GND.n4423 585
R11862 GND.n7698 GND.n4423 585
R11863 GND.n4482 GND.n4481 585
R11864 GND.n4481 GND.n4422 585
R11865 GND.n4480 GND.n4415 585
R11866 GND.n7704 GND.n4415 585
R11867 GND.n4479 GND.n4478 585
R11868 GND.n4478 GND.n4414 585
R11869 GND.n4477 GND.n4455 585
R11870 GND.n4477 GND.n4476 585
R11871 GND.n4472 GND.n4471 585
R11872 GND.n4472 GND.n4406 585
R11873 GND.n4470 GND.n4405 585
R11874 GND.n7712 GND.n4405 585
R11875 GND.n4469 GND.n4468 585
R11876 GND.n4468 GND.n4404 585
R11877 GND.n4467 GND.n4397 585
R11878 GND.n7718 GND.n4397 585
R11879 GND.n4466 GND.n4465 585
R11880 GND.n4465 GND.n4396 585
R11881 GND.n4464 GND.n4456 585
R11882 GND.n4464 GND.n4463 585
R11883 GND.n4459 GND.n4458 585
R11884 GND.n4459 GND.n4384 585
R11885 GND.n4457 GND.n4383 585
R11886 GND.n7726 GND.n4383 585
R11887 GND.n4374 GND.n4373 585
R11888 GND.n4382 GND.n4374 585
R11889 GND.n7734 GND.n7733 585
R11890 GND.n7733 GND.n7732 585
R11891 GND.n7735 GND.n4371 585
R11892 GND.n4371 GND.n4368 585
R11893 GND.n7737 GND.n7736 585
R11894 GND.n7738 GND.n7737 585
R11895 GND.n4372 GND.n4370 585
R11896 GND.n4370 GND.n4365 585
R11897 GND.n5788 GND.n5787 585
R11898 GND.n5787 GND.n4357 585
R11899 GND.n5789 GND.n4868 585
R11900 GND.n4868 GND.n4355 585
R11901 GND.n5791 GND.n5790 585
R11902 GND.n5792 GND.n5791 585
R11903 GND.n5786 GND.n4866 585
R11904 GND.n5794 GND.n4866 585
R11905 GND.n5785 GND.n5784 585
R11906 GND.n5784 GND.n4346 585
R11907 GND.n5783 GND.n4853 585
R11908 GND.n5800 GND.n4853 585
R11909 GND.n5782 GND.n5781 585
R11910 GND.n5781 GND.n4338 585
R11911 GND.n5780 GND.n4869 585
R11912 GND.n5780 GND.n4336 585
R11913 GND.n5779 GND.n4871 585
R11914 GND.n5779 GND.n5778 585
R11915 GND.n5766 GND.n4870 585
R11916 GND.n4870 GND.n4328 585
R11917 GND.n5767 GND.n4879 585
R11918 GND.n4879 GND.n4326 585
R11919 GND.n5769 GND.n5768 585
R11920 GND.n5770 GND.n5769 585
R11921 GND.n5765 GND.n4878 585
R11922 GND.n4878 GND.n4318 585
R11923 GND.n5764 GND.n5763 585
R11924 GND.n5763 GND.n4316 585
R11925 GND.n5762 GND.n4880 585
R11926 GND.n5762 GND.n5761 585
R11927 GND.n5748 GND.n4881 585
R11928 GND.n4881 GND.n4295 585
R11929 GND.n5749 GND.n5745 585
R11930 GND.n5745 GND.n4293 585
R11931 GND.n5751 GND.n5750 585
R11932 GND.n5752 GND.n5751 585
R11933 GND.n5747 GND.n5744 585
R11934 GND.n5744 GND.n4281 585
R11935 GND.n5746 GND.n4279 585
R11936 GND.n7781 GND.n4279 585
R11937 GND.n4270 GND.n4269 585
R11938 GND.n4278 GND.n4270 585
R11939 GND.n7789 GND.n7788 585
R11940 GND.n7788 GND.n7787 585
R11941 GND.n7790 GND.n4267 585
R11942 GND.n4267 GND.n4264 585
R11943 GND.n7792 GND.n7791 585
R11944 GND.n7793 GND.n7792 585
R11945 GND.n4268 GND.n4266 585
R11946 GND.n4266 GND.n4261 585
R11947 GND.n5690 GND.n5689 585
R11948 GND.n5690 GND.n4253 585
R11949 GND.n5692 GND.n5691 585
R11950 GND.n5691 GND.n4251 585
R11951 GND.n5693 GND.n4894 585
R11952 GND.n5709 GND.n4894 585
R11953 GND.n5694 GND.n4901 585
R11954 GND.n4901 GND.n4893 585
R11955 GND.n5696 GND.n5695 585
R11956 GND.n5697 GND.n5696 585
R11957 GND.n5688 GND.n4900 585
R11958 GND.n4900 GND.n4899 585
R11959 GND.n5687 GND.n5686 585
R11960 GND.n5686 GND.n4235 585
R11961 GND.n5685 GND.n4902 585
R11962 GND.n5685 GND.n4233 585
R11963 GND.n5684 GND.n4904 585
R11964 GND.n5684 GND.n5683 585
R11965 GND.n5669 GND.n4903 585
R11966 GND.n4903 GND.n4225 585
R11967 GND.n5670 GND.n4912 585
R11968 GND.n4912 GND.n4223 585
R11969 GND.n5672 GND.n5671 585
R11970 GND.n5673 GND.n5672 585
R11971 GND.n5668 GND.n4911 585
R11972 GND.n4911 GND.n4215 585
R11973 GND.n5667 GND.n5666 585
R11974 GND.n5666 GND.n4213 585
R11975 GND.n5665 GND.n4913 585
R11976 GND.n5665 GND.n5664 585
R11977 GND.n5651 GND.n4914 585
R11978 GND.n4916 GND.n4914 585
R11979 GND.n5652 GND.n5648 585
R11980 GND.n5648 GND.n4191 585
R11981 GND.n5654 GND.n5653 585
R11982 GND.n5655 GND.n5654 585
R11983 GND.n5650 GND.n5647 585
R11984 GND.n5647 GND.n4179 585
R11985 GND.n5649 GND.n4177 585
R11986 GND.n7836 GND.n4177 585
R11987 GND.n4168 GND.n4167 585
R11988 GND.n4176 GND.n4168 585
R11989 GND.n7844 GND.n7843 585
R11990 GND.n7843 GND.n7842 585
R11991 GND.n7845 GND.n4165 585
R11992 GND.n4165 GND.n4162 585
R11993 GND.n7847 GND.n7846 585
R11994 GND.n7848 GND.n7847 585
R11995 GND.n4166 GND.n4164 585
R11996 GND.n4164 GND.n4159 585
R11997 GND.n5584 GND.n5583 585
R11998 GND.n5584 GND.n4151 585
R11999 GND.n5586 GND.n5585 585
R12000 GND.n5585 GND.n4149 585
R12001 GND.n5587 GND.n4927 585
R12002 GND.n5606 GND.n4927 585
R12003 GND.n5589 GND.n5588 585
R12004 GND.n5588 GND.n4141 585
R12005 GND.n5590 GND.n4934 585
R12006 GND.n4934 GND.n4139 585
R12007 GND.n5592 GND.n5591 585
R12008 GND.n5593 GND.n5592 585
R12009 GND.n5582 GND.n4933 585
R12010 GND.n4933 GND.n4131 585
R12011 GND.n5581 GND.n5580 585
R12012 GND.n5580 GND.n4129 585
R12013 GND.n5579 GND.n4935 585
R12014 GND.n5579 GND.n5578 585
R12015 GND.n5565 GND.n4936 585
R12016 GND.n4936 GND.n4121 585
R12017 GND.n5566 GND.n4944 585
R12018 GND.n4944 GND.n4119 585
R12019 GND.n5568 GND.n5567 585
R12020 GND.n5569 GND.n5568 585
R12021 GND.n5564 GND.n4943 585
R12022 GND.n4943 GND.n4111 585
R12023 GND.n5563 GND.n5562 585
R12024 GND.n5562 GND.n4109 585
R12025 GND.n5561 GND.n4945 585
R12026 GND.n5561 GND.n5560 585
R12027 GND.n5547 GND.n4946 585
R12028 GND.n4946 GND.n4088 585
R12029 GND.n5548 GND.n5544 585
R12030 GND.n5544 GND.n4086 585
R12031 GND.n5550 GND.n5549 585
R12032 GND.n5551 GND.n5550 585
R12033 GND.n5546 GND.n5543 585
R12034 GND.n5543 GND.n4074 585
R12035 GND.n5545 GND.n4072 585
R12036 GND.n7891 GND.n4072 585
R12037 GND.n4063 GND.n4062 585
R12038 GND.n4071 GND.n4063 585
R12039 GND.n7899 GND.n7898 585
R12040 GND.n7898 GND.n7897 585
R12041 GND.n7900 GND.n4060 585
R12042 GND.n4060 GND.n4057 585
R12043 GND.n7902 GND.n7901 585
R12044 GND.n7903 GND.n7902 585
R12045 GND.n4061 GND.n4059 585
R12046 GND.n4059 GND.n4054 585
R12047 GND.n5481 GND.n5480 585
R12048 GND.n5481 GND.n4046 585
R12049 GND.n5483 GND.n5482 585
R12050 GND.n5482 GND.n4044 585
R12051 GND.n5484 GND.n4958 585
R12052 GND.n5503 GND.n4958 585
R12053 GND.n5486 GND.n5485 585
R12054 GND.n5485 GND.n4036 585
R12055 GND.n5487 GND.n4965 585
R12056 GND.n4965 GND.n4034 585
R12057 GND.n5489 GND.n5488 585
R12058 GND.n5490 GND.n5489 585
R12059 GND.n5479 GND.n4964 585
R12060 GND.n4964 GND.n4026 585
R12061 GND.n5478 GND.n5477 585
R12062 GND.n5477 GND.n4024 585
R12063 GND.n5476 GND.n4966 585
R12064 GND.n5476 GND.n5475 585
R12065 GND.n5462 GND.n4967 585
R12066 GND.n4967 GND.n4016 585
R12067 GND.n5463 GND.n4975 585
R12068 GND.n4975 GND.n4014 585
R12069 GND.n5465 GND.n5464 585
R12070 GND.n5466 GND.n5465 585
R12071 GND.n5461 GND.n4974 585
R12072 GND.n4974 GND.n4006 585
R12073 GND.n5460 GND.n5459 585
R12074 GND.n5459 GND.n4004 585
R12075 GND.n5458 GND.n4976 585
R12076 GND.n5458 GND.n5457 585
R12077 GND.n5444 GND.n4977 585
R12078 GND.n4977 GND.n3996 585
R12079 GND.n5445 GND.n4984 585
R12080 GND.n4984 GND.n3994 585
R12081 GND.n5447 GND.n5446 585
R12082 GND.n5448 GND.n5447 585
R12083 GND.n5443 GND.n4983 585
R12084 GND.n4983 GND.n3986 585
R12085 GND.n5442 GND.n5441 585
R12086 GND.n5441 GND.n3984 585
R12087 GND.n5440 GND.n4985 585
R12088 GND.n5440 GND.n5439 585
R12089 GND.n5426 GND.n4986 585
R12090 GND.n4986 GND.n3976 585
R12091 GND.n5427 GND.n4994 585
R12092 GND.n4994 GND.n3974 585
R12093 GND.n5429 GND.n5428 585
R12094 GND.n5430 GND.n5429 585
R12095 GND.n5425 GND.n4993 585
R12096 GND.n4993 GND.n3966 585
R12097 GND.n5424 GND.n5423 585
R12098 GND.n5423 GND.n3964 585
R12099 GND.n5422 GND.n4995 585
R12100 GND.n5422 GND.n5421 585
R12101 GND.n5264 GND.n4996 585
R12102 GND.n4996 GND.n3956 585
R12103 GND.n5266 GND.n5265 585
R12104 GND.n5265 GND.n3954 585
R12105 GND.n5267 GND.n5002 585
R12106 GND.n5412 GND.n5002 585
R12107 GND.n5269 GND.n5268 585
R12108 GND.n5269 GND.n3946 585
R12109 GND.n5271 GND.n5270 585
R12110 GND.n5270 GND.n3944 585
R12111 GND.n5272 GND.n5006 585
R12112 GND.n5361 GND.n5006 585
R12113 GND.n5274 GND.n5273 585
R12114 GND.n5274 GND.n3936 585
R12115 GND.n5276 GND.n5275 585
R12116 GND.n5275 GND.n3934 585
R12117 GND.n5277 GND.n5011 585
R12118 GND.n5352 GND.n5011 585
R12119 GND.n5279 GND.n5278 585
R12120 GND.n5279 GND.n3926 585
R12121 GND.n5281 GND.n5280 585
R12122 GND.n5280 GND.n3924 585
R12123 GND.n5282 GND.n5015 585
R12124 GND.n5342 GND.n5015 585
R12125 GND.n5284 GND.n5283 585
R12126 GND.n5284 GND.n3916 585
R12127 GND.n5286 GND.n5285 585
R12128 GND.n5285 GND.n3914 585
R12129 GND.n5287 GND.n5020 585
R12130 GND.n5333 GND.n5020 585
R12131 GND.n5289 GND.n5288 585
R12132 GND.n5288 GND.n3906 585
R12133 GND.n5290 GND.n5031 585
R12134 GND.n5323 GND.n5031 585
R12135 GND.n5291 GND.n5263 585
R12136 GND.n5263 GND.n5030 585
R12137 GND.n5293 GND.n5292 585
R12138 GND.n5293 GND.n3895 585
R12139 GND.n5294 GND.n5262 585
R12140 GND.n5294 GND.n3893 585
R12141 GND.n5296 GND.n5295 585
R12142 GND.n5295 GND.n3884 585
R12143 GND.n5297 GND.n3885 585
R12144 GND.n8005 GND.n3885 585
R12145 GND.n5299 GND.n5298 585
R12146 GND.n5299 GND.n3882 585
R12147 GND.n5301 GND.n5300 585
R12148 GND.n5300 GND.n3861 585
R12149 GND.n5302 GND.n5037 585
R12150 GND.n5037 GND.n3850 585
R12151 GND.n5304 GND.n5303 585
R12152 GND.n5305 GND.n5304 585
R12153 GND.n5261 GND.n5036 585
R12154 GND.n5036 GND.n3842 585
R12155 GND.n5260 GND.n3841 585
R12156 GND.n8064 GND.n3841 585
R12157 GND.n5259 GND.n5258 585
R12158 GND.n5258 GND.n3840 585
R12159 GND.n5257 GND.n3833 585
R12160 GND.n8070 GND.n3833 585
R12161 GND.n5256 GND.n5255 585
R12162 GND.n5255 GND.n3832 585
R12163 GND.n5254 GND.n5038 585
R12164 GND.n5254 GND.n5253 585
R12165 GND.n5249 GND.n5248 585
R12166 GND.n5249 GND.n3824 585
R12167 GND.n5247 GND.n3823 585
R12168 GND.n8078 GND.n3823 585
R12169 GND.n5246 GND.n5245 585
R12170 GND.n5245 GND.n3822 585
R12171 GND.n5244 GND.n3815 585
R12172 GND.n8084 GND.n3815 585
R12173 GND.n5243 GND.n5242 585
R12174 GND.n5242 GND.n3814 585
R12175 GND.n5241 GND.n5039 585
R12176 GND.n5241 GND.n5240 585
R12177 GND.n5236 GND.n5235 585
R12178 GND.n5236 GND.n3806 585
R12179 GND.n5234 GND.n3805 585
R12180 GND.n8092 GND.n3805 585
R12181 GND.n5233 GND.n5232 585
R12182 GND.n5232 GND.n3804 585
R12183 GND.n5231 GND.n3797 585
R12184 GND.n8098 GND.n3797 585
R12185 GND.n5230 GND.n5229 585
R12186 GND.n5229 GND.n3796 585
R12187 GND.n5228 GND.n5040 585
R12188 GND.n5228 GND.n5227 585
R12189 GND.n5223 GND.n5222 585
R12190 GND.n5223 GND.n3788 585
R12191 GND.n5221 GND.n3787 585
R12192 GND.n8106 GND.n3787 585
R12193 GND.n5220 GND.n5219 585
R12194 GND.n5219 GND.t64 585
R12195 GND.n5218 GND.n3781 585
R12196 GND.n8112 GND.n3781 585
R12197 GND.n5217 GND.n5216 585
R12198 GND.n5216 GND.n3780 585
R12199 GND.n5215 GND.n5041 585
R12200 GND.n5215 GND.n5214 585
R12201 GND.n5210 GND.n5209 585
R12202 GND.n5210 GND.n3772 585
R12203 GND.n5208 GND.n3771 585
R12204 GND.n8120 GND.n3771 585
R12205 GND.n5207 GND.n5206 585
R12206 GND.n5206 GND.n3751 585
R12207 GND.n5205 GND.n3750 585
R12208 GND.n8126 GND.n3750 585
R12209 GND.n8307 GND.n2126 585
R12210 GND.n8480 GND.n2126 585
R12211 GND.n8306 GND.n8305 585
R12212 GND.n8305 GND.n8304 585
R12213 GND.n2213 GND.n2212 585
R12214 GND.n2222 GND.n2213 585
R12215 GND.n8293 GND.n8292 585
R12216 GND.n8294 GND.n8293 585
R12217 GND.n2227 GND.n2226 585
R12218 GND.n8282 GND.n2226 585
R12219 GND.n8287 GND.n8286 585
R12220 GND.n8286 GND.n8285 585
R12221 GND.n2230 GND.n2229 585
R12222 GND.n8280 GND.n2230 585
R12223 GND.n8267 GND.n2248 585
R12224 GND.n2248 GND.n2247 585
R12225 GND.n8269 GND.n8268 585
R12226 GND.n8270 GND.n8269 585
R12227 GND.n2249 GND.n2246 585
R12228 GND.n8257 GND.n2246 585
R12229 GND.n8262 GND.n8261 585
R12230 GND.n8261 GND.n8260 585
R12231 GND.n2252 GND.n2251 585
R12232 GND.n8254 GND.n2252 585
R12233 GND.n8241 GND.n2270 585
R12234 GND.n2270 GND.n2269 585
R12235 GND.n8243 GND.n8242 585
R12236 GND.n8244 GND.n8243 585
R12237 GND.n2271 GND.n2268 585
R12238 GND.n8230 GND.n2268 585
R12239 GND.n8236 GND.n8235 585
R12240 GND.n8235 GND.n8234 585
R12241 GND.n2274 GND.n2273 585
R12242 GND.n8228 GND.n2274 585
R12243 GND.n8215 GND.n2291 585
R12244 GND.n2291 GND.n2290 585
R12245 GND.n8217 GND.n8216 585
R12246 GND.n8218 GND.n8217 585
R12247 GND.n2292 GND.n2288 585
R12248 GND.n8205 GND.n2288 585
R12249 GND.n8210 GND.n8209 585
R12250 GND.n8209 GND.n8208 585
R12251 GND.n2295 GND.n2294 585
R12252 GND.n8202 GND.n2295 585
R12253 GND.n8189 GND.n2312 585
R12254 GND.n2312 GND.n2311 585
R12255 GND.n8191 GND.n8190 585
R12256 GND.n8192 GND.n8191 585
R12257 GND.n2313 GND.n2310 585
R12258 GND.n8179 GND.n2310 585
R12259 GND.n8184 GND.n8183 585
R12260 GND.n8183 GND.n8182 585
R12261 GND.n2316 GND.n2315 585
R12262 GND.n3691 GND.n2316 585
R12263 GND.n3678 GND.n2340 585
R12264 GND.n2340 GND.n2328 585
R12265 GND.n3680 GND.n3679 585
R12266 GND.n3681 GND.n3680 585
R12267 GND.n2341 GND.n2339 585
R12268 GND.n3668 GND.n2339 585
R12269 GND.n3673 GND.n3672 585
R12270 GND.n3672 GND.n3671 585
R12271 GND.n2344 GND.n2343 585
R12272 GND.n3665 GND.n2344 585
R12273 GND.n3652 GND.n2362 585
R12274 GND.n2362 GND.n2361 585
R12275 GND.n3654 GND.n3653 585
R12276 GND.n3655 GND.n3654 585
R12277 GND.n2363 GND.n2360 585
R12278 GND.n3641 GND.n2360 585
R12279 GND.n3647 GND.n3646 585
R12280 GND.n3646 GND.n3645 585
R12281 GND.n2366 GND.n2365 585
R12282 GND.n3639 GND.n2366 585
R12283 GND.n3626 GND.n2380 585
R12284 GND.n2605 GND.n2380 585
R12285 GND.n3628 GND.n3627 585
R12286 GND.n3629 GND.n3628 585
R12287 GND.n2381 GND.n2379 585
R12288 GND.n3616 GND.n2379 585
R12289 GND.n3621 GND.n3620 585
R12290 GND.n3620 GND.n3619 585
R12291 GND.n2384 GND.n2383 585
R12292 GND.n3613 GND.n2384 585
R12293 GND.n3600 GND.n2402 585
R12294 GND.n2402 GND.n2401 585
R12295 GND.n3602 GND.n3601 585
R12296 GND.n3603 GND.n3602 585
R12297 GND.n2403 GND.n2400 585
R12298 GND.n3590 GND.n2400 585
R12299 GND.n3595 GND.n3594 585
R12300 GND.n3594 GND.n3593 585
R12301 GND.n2406 GND.n2405 585
R12302 GND.n3588 GND.n2406 585
R12303 GND.n3575 GND.n2424 585
R12304 GND.n2424 GND.n2423 585
R12305 GND.n3577 GND.n3576 585
R12306 GND.n3578 GND.n3577 585
R12307 GND.n2425 GND.n2422 585
R12308 GND.n3565 GND.n2422 585
R12309 GND.n3570 GND.n3569 585
R12310 GND.n3569 GND.n3568 585
R12311 GND.n2428 GND.n2427 585
R12312 GND.n3562 GND.n2428 585
R12313 GND.n3549 GND.n2446 585
R12314 GND.n2446 GND.n2445 585
R12315 GND.n3551 GND.n3550 585
R12316 GND.n3552 GND.n3551 585
R12317 GND.n2447 GND.n2444 585
R12318 GND.n3538 GND.n2444 585
R12319 GND.n3544 GND.n3543 585
R12320 GND.n3543 GND.n3542 585
R12321 GND.n2450 GND.n2449 585
R12322 GND.n3536 GND.n2450 585
R12323 GND.n3523 GND.n2467 585
R12324 GND.n2467 GND.n2466 585
R12325 GND.n3525 GND.n3524 585
R12326 GND.n3526 GND.n3525 585
R12327 GND.n2468 GND.n2464 585
R12328 GND.n3513 GND.n2464 585
R12329 GND.n3518 GND.n3517 585
R12330 GND.n3517 GND.n3516 585
R12331 GND.n2471 GND.n2470 585
R12332 GND.n3510 GND.n2471 585
R12333 GND.n3497 GND.n2489 585
R12334 GND.n2489 GND.n2488 585
R12335 GND.n3499 GND.n3498 585
R12336 GND.n3500 GND.n3499 585
R12337 GND.n2490 GND.n2487 585
R12338 GND.n3461 GND.n2487 585
R12339 GND.n3457 GND.n3456 585
R12340 GND.n3458 GND.n3457 585
R12341 GND.n3455 GND.n3454 585
R12342 GND.n3455 GND.n2531 585
R12343 GND.n3453 GND.n2525 585
R12344 GND.n3470 GND.n2525 585
R12345 GND.n3475 GND.n3474 585
R12346 GND.n3474 GND.n3473 585
R12347 GND.n3477 GND.n3476 585
R12348 GND.n3478 GND.n3477 585
R12349 GND.n2524 GND.n2523 585
R12350 GND.n2524 GND.n2516 585
R12351 GND.n2522 GND.n2496 585
R12352 GND.n2522 GND.n2509 585
R12353 GND.n2500 GND.n2497 585
R12354 GND.n3487 GND.n2500 585
R12355 GND.n3492 GND.n3491 585
R12356 GND.n3491 GND.n3490 585
R12357 GND.n2499 GND.n2498 585
R12358 GND.n3064 GND.n2499 585
R12359 GND.n3429 GND.n3428 585
R12360 GND.n3430 GND.n3429 585
R12361 GND.n2665 GND.n2664 585
R12362 GND.n3419 GND.n2664 585
R12363 GND.n3424 GND.n3423 585
R12364 GND.n3423 GND.n3422 585
R12365 GND.n2668 GND.n2667 585
R12366 GND.n3417 GND.n2668 585
R12367 GND.n3405 GND.n2687 585
R12368 GND.n2687 GND.n2686 585
R12369 GND.n3407 GND.n3406 585
R12370 GND.n3408 GND.n3407 585
R12371 GND.n2688 GND.n2685 585
R12372 GND.n3395 GND.n2685 585
R12373 GND.n3400 GND.n3399 585
R12374 GND.n3399 GND.n3398 585
R12375 GND.n2691 GND.n2690 585
R12376 GND.n3392 GND.n2691 585
R12377 GND.n3380 GND.n2710 585
R12378 GND.n2710 GND.n2709 585
R12379 GND.n3382 GND.n3381 585
R12380 GND.n3383 GND.n3382 585
R12381 GND.n2711 GND.n2708 585
R12382 GND.n3369 GND.n2708 585
R12383 GND.n3375 GND.n3374 585
R12384 GND.n3374 GND.n3373 585
R12385 GND.n2714 GND.n2713 585
R12386 GND.n3367 GND.n2714 585
R12387 GND.n3355 GND.n2732 585
R12388 GND.n2732 GND.n2731 585
R12389 GND.n3357 GND.n3356 585
R12390 GND.n3358 GND.n3357 585
R12391 GND.n2733 GND.n2729 585
R12392 GND.n3345 GND.n2729 585
R12393 GND.n3350 GND.n3349 585
R12394 GND.n3349 GND.n3348 585
R12395 GND.n2736 GND.n2735 585
R12396 GND.n3342 GND.n2736 585
R12397 GND.n3330 GND.n2755 585
R12398 GND.n2755 GND.n2754 585
R12399 GND.n3332 GND.n3331 585
R12400 GND.n3333 GND.n3332 585
R12401 GND.n2756 GND.n2753 585
R12402 GND.n3320 GND.n2753 585
R12403 GND.n3325 GND.n3324 585
R12404 GND.n3324 GND.n3323 585
R12405 GND.n2759 GND.n2758 585
R12406 GND.n3318 GND.n2759 585
R12407 GND.n3306 GND.n2778 585
R12408 GND.n2778 GND.n2777 585
R12409 GND.n3308 GND.n3307 585
R12410 GND.n3309 GND.n3308 585
R12411 GND.n2779 GND.n2776 585
R12412 GND.n3296 GND.n2776 585
R12413 GND.n3301 GND.n3300 585
R12414 GND.n3300 GND.n3299 585
R12415 GND.n2782 GND.n2781 585
R12416 GND.n3293 GND.n2782 585
R12417 GND.n3281 GND.n2801 585
R12418 GND.n2801 GND.n2800 585
R12419 GND.n3283 GND.n3282 585
R12420 GND.n3284 GND.n3283 585
R12421 GND.n2802 GND.n2799 585
R12422 GND.n3270 GND.n2799 585
R12423 GND.n3276 GND.n3275 585
R12424 GND.n3275 GND.n3274 585
R12425 GND.n2805 GND.n2804 585
R12426 GND.n3268 GND.n2805 585
R12427 GND.n3256 GND.n2823 585
R12428 GND.n2823 GND.n2822 585
R12429 GND.n3258 GND.n3257 585
R12430 GND.n3259 GND.n3258 585
R12431 GND.n2824 GND.n2820 585
R12432 GND.n3246 GND.n2820 585
R12433 GND.n3251 GND.n3250 585
R12434 GND.n3250 GND.n3249 585
R12435 GND.n2827 GND.n2826 585
R12436 GND.n3243 GND.n2827 585
R12437 GND.n3231 GND.n2846 585
R12438 GND.n2846 GND.n2845 585
R12439 GND.n3233 GND.n3232 585
R12440 GND.n3234 GND.n3233 585
R12441 GND.n2847 GND.n2844 585
R12442 GND.n3221 GND.n2844 585
R12443 GND.n3226 GND.n3225 585
R12444 GND.n3225 GND.n3224 585
R12445 GND.n2850 GND.n2849 585
R12446 GND.n3219 GND.n2850 585
R12447 GND.n3207 GND.n2869 585
R12448 GND.n2869 GND.n2868 585
R12449 GND.n3209 GND.n3208 585
R12450 GND.n3210 GND.n3209 585
R12451 GND.n2870 GND.n2867 585
R12452 GND.n3197 GND.n2867 585
R12453 GND.n3202 GND.n3201 585
R12454 GND.n3201 GND.n3200 585
R12455 GND.n2873 GND.n2872 585
R12456 GND.n3194 GND.n2873 585
R12457 GND.n3182 GND.n2892 585
R12458 GND.n2892 GND.n2891 585
R12459 GND.n3184 GND.n3183 585
R12460 GND.n3185 GND.n3184 585
R12461 GND.n2893 GND.n2890 585
R12462 GND.n3171 GND.n2890 585
R12463 GND.n3177 GND.n3176 585
R12464 GND.n3176 GND.n3175 585
R12465 GND.n2896 GND.n2895 585
R12466 GND.n3169 GND.n2896 585
R12467 GND.n3157 GND.n3153 585
R12468 GND.n3153 GND.n3152 585
R12469 GND.n3159 GND.n3158 585
R12470 GND.n3160 GND.n3159 585
R12471 GND.n1835 GND.n1834 585
R12472 GND.n2964 GND.n1835 585
R12473 GND.n8686 GND.n8685 585
R12474 GND.n8685 GND.n8684 585
R12475 GND.n8687 GND.n1823 585
R12476 GND.n2907 GND.n1823 585
R12477 GND.n8689 GND.n8688 585
R12478 GND.n8690 GND.n8689 585
R12479 GND.n1824 GND.n1822 585
R12480 GND.n1822 GND.n1817 585
R12481 GND.n1828 GND.n1827 585
R12482 GND.n1827 GND.n1805 585
R12483 GND.n1826 GND.n1728 585
R12484 GND.n8698 GND.n1728 585
R12485 GND.n8814 GND.n8813 585
R12486 GND.n8812 GND.n1727 585
R12487 GND.n8811 GND.n1726 585
R12488 GND.n8816 GND.n1726 585
R12489 GND.n8810 GND.n8809 585
R12490 GND.n8808 GND.n8807 585
R12491 GND.n8806 GND.n8805 585
R12492 GND.n8804 GND.n8803 585
R12493 GND.n8802 GND.n8801 585
R12494 GND.n8800 GND.n8799 585
R12495 GND.n8798 GND.n8797 585
R12496 GND.n8796 GND.n8795 585
R12497 GND.n8794 GND.n8793 585
R12498 GND.n8792 GND.n1741 585
R12499 GND.n8791 GND.n8790 585
R12500 GND.n8789 GND.n8788 585
R12501 GND.n8787 GND.n8786 585
R12502 GND.n8785 GND.n8784 585
R12503 GND.n8783 GND.n8782 585
R12504 GND.n8781 GND.n8780 585
R12505 GND.n8779 GND.n8778 585
R12506 GND.n8777 GND.n8776 585
R12507 GND.n8775 GND.n8774 585
R12508 GND.n8773 GND.n8772 585
R12509 GND.n8771 GND.n8770 585
R12510 GND.n8769 GND.n8768 585
R12511 GND.n8767 GND.n8766 585
R12512 GND.n8765 GND.n8764 585
R12513 GND.n8763 GND.n8762 585
R12514 GND.n8761 GND.n8760 585
R12515 GND.n8759 GND.n8758 585
R12516 GND.n8757 GND.n8756 585
R12517 GND.n8755 GND.n8754 585
R12518 GND.n8753 GND.n8752 585
R12519 GND.n8751 GND.n8750 585
R12520 GND.n8749 GND.n8748 585
R12521 GND.n8747 GND.n8746 585
R12522 GND.n8745 GND.n8744 585
R12523 GND.n8743 GND.n8742 585
R12524 GND.n8741 GND.n8740 585
R12525 GND.n8739 GND.n8738 585
R12526 GND.n8737 GND.n8736 585
R12527 GND.n8735 GND.n8734 585
R12528 GND.n8733 GND.n8732 585
R12529 GND.n8731 GND.n8730 585
R12530 GND.n8729 GND.n8728 585
R12531 GND.n8727 GND.n8726 585
R12532 GND.n8725 GND.n8724 585
R12533 GND.n8723 GND.n8722 585
R12534 GND.n8721 GND.n8720 585
R12535 GND.n8719 GND.n8718 585
R12536 GND.n8717 GND.n8716 585
R12537 GND.n8715 GND.n8714 585
R12538 GND.n8713 GND.n8712 585
R12539 GND.n8711 GND.n8710 585
R12540 GND.n8709 GND.n8708 585
R12541 GND.n8707 GND.n8706 585
R12542 GND.n1802 GND.n1793 585
R12543 GND.n8411 GND.n2124 585
R12544 GND.n8412 GND.n8409 585
R12545 GND.n8413 GND.n8405 585
R12546 GND.n8414 GND.n8404 585
R12547 GND.n8403 GND.n8401 585
R12548 GND.n8418 GND.n8400 585
R12549 GND.n8419 GND.n8399 585
R12550 GND.n8420 GND.n8398 585
R12551 GND.n8397 GND.n8395 585
R12552 GND.n8424 GND.n8394 585
R12553 GND.n8425 GND.n8393 585
R12554 GND.n8426 GND.n8392 585
R12555 GND.n8391 GND.n8389 585
R12556 GND.n8430 GND.n8388 585
R12557 GND.n8431 GND.n8387 585
R12558 GND.n8432 GND.n8386 585
R12559 GND.n8385 GND.n8380 585
R12560 GND.n8436 GND.n8379 585
R12561 GND.n8437 GND.n8378 585
R12562 GND.n8438 GND.n8377 585
R12563 GND.n8376 GND.n8374 585
R12564 GND.n8442 GND.n8373 585
R12565 GND.n8443 GND.n8372 585
R12566 GND.n8444 GND.n8371 585
R12567 GND.n8370 GND.n8368 585
R12568 GND.n8448 GND.n8367 585
R12569 GND.n8449 GND.n8366 585
R12570 GND.n8450 GND.n8365 585
R12571 GND.n8364 GND.n2186 585
R12572 GND.n8455 GND.n8454 585
R12573 GND.n8457 GND.n8456 585
R12574 GND.n8360 GND.n8359 585
R12575 GND.n8358 GND.n8357 585
R12576 GND.n8356 GND.n2190 585
R12577 GND.n2189 GND.n2188 585
R12578 GND.n8352 GND.n8351 585
R12579 GND.n8350 GND.n8349 585
R12580 GND.n8348 GND.n2194 585
R12581 GND.n2193 GND.n2192 585
R12582 GND.n8344 GND.n8343 585
R12583 GND.n8342 GND.n8341 585
R12584 GND.n8340 GND.n2198 585
R12585 GND.n2197 GND.n2196 585
R12586 GND.n8336 GND.n8335 585
R12587 GND.n8334 GND.n8331 585
R12588 GND.n8330 GND.n2202 585
R12589 GND.n2201 GND.n2200 585
R12590 GND.n8326 GND.n8325 585
R12591 GND.n8324 GND.n8323 585
R12592 GND.n8322 GND.n2206 585
R12593 GND.n2205 GND.n2204 585
R12594 GND.n8318 GND.n8317 585
R12595 GND.n8316 GND.n8315 585
R12596 GND.n8314 GND.n2210 585
R12597 GND.n2209 GND.n2208 585
R12598 GND.n8310 GND.n8309 585
R12599 GND.n8482 GND.n8481 585
R12600 GND.n8481 GND.n8480 585
R12601 GND.n2123 GND.n2118 585
R12602 GND.n8304 GND.n2123 585
R12603 GND.n8486 GND.n2117 585
R12604 GND.n2222 GND.n2117 585
R12605 GND.n8487 GND.n2116 585
R12606 GND.n8294 GND.n2116 585
R12607 GND.n8488 GND.n2115 585
R12608 GND.n8282 GND.n2115 585
R12609 GND.n2232 GND.n2110 585
R12610 GND.n8285 GND.n2232 585
R12611 GND.n8492 GND.n2109 585
R12612 GND.n8280 GND.n2109 585
R12613 GND.n8493 GND.n2108 585
R12614 GND.n2247 GND.n2108 585
R12615 GND.n8494 GND.n2107 585
R12616 GND.n8270 GND.n2107 585
R12617 GND.n8256 GND.n2102 585
R12618 GND.n8257 GND.n8256 585
R12619 GND.n8498 GND.n2101 585
R12620 GND.n8260 GND.n2101 585
R12621 GND.n8499 GND.n2100 585
R12622 GND.n8254 GND.n2100 585
R12623 GND.n8500 GND.n2099 585
R12624 GND.n2269 GND.n2099 585
R12625 GND.n2265 GND.n2094 585
R12626 GND.n8244 GND.n2265 585
R12627 GND.n8504 GND.n2093 585
R12628 GND.n8230 GND.n2093 585
R12629 GND.n8505 GND.n2092 585
R12630 GND.n8234 GND.n2092 585
R12631 GND.n8506 GND.n2091 585
R12632 GND.n8228 GND.n2091 585
R12633 GND.n2289 GND.n2086 585
R12634 GND.n2290 GND.n2289 585
R12635 GND.n8510 GND.n2085 585
R12636 GND.n8218 GND.n2085 585
R12637 GND.n8511 GND.n2084 585
R12638 GND.n8205 GND.n2084 585
R12639 GND.n8512 GND.n2083 585
R12640 GND.n8208 GND.n2083 585
R12641 GND.n2301 GND.n2078 585
R12642 GND.n8202 GND.n2301 585
R12643 GND.n8516 GND.n2077 585
R12644 GND.n2311 GND.n2077 585
R12645 GND.n8517 GND.n2076 585
R12646 GND.n8192 GND.n2076 585
R12647 GND.n8518 GND.n2075 585
R12648 GND.n8179 GND.n2075 585
R12649 GND.n2318 GND.n2070 585
R12650 GND.n8182 GND.n2318 585
R12651 GND.n8522 GND.n2069 585
R12652 GND.n3691 GND.n2069 585
R12653 GND.n8523 GND.n2068 585
R12654 GND.n2328 GND.n2068 585
R12655 GND.n8524 GND.n2067 585
R12656 GND.n3681 GND.n2067 585
R12657 GND.n3667 GND.n2062 585
R12658 GND.n3668 GND.n3667 585
R12659 GND.n8528 GND.n2061 585
R12660 GND.n3671 GND.n2061 585
R12661 GND.n8529 GND.n2060 585
R12662 GND.n3665 GND.n2060 585
R12663 GND.n8530 GND.n2059 585
R12664 GND.n2361 GND.n2059 585
R12665 GND.n2357 GND.n2054 585
R12666 GND.n3655 GND.n2357 585
R12667 GND.n8534 GND.n2053 585
R12668 GND.n3641 GND.n2053 585
R12669 GND.n8535 GND.n2052 585
R12670 GND.n3645 GND.n2052 585
R12671 GND.n8536 GND.n2051 585
R12672 GND.n3639 GND.n2051 585
R12673 GND.n2604 GND.n2046 585
R12674 GND.n2605 GND.n2604 585
R12675 GND.n8540 GND.n2045 585
R12676 GND.n3629 GND.n2045 585
R12677 GND.n8541 GND.n2044 585
R12678 GND.n3616 GND.n2044 585
R12679 GND.n8542 GND.n2043 585
R12680 GND.n3619 GND.n2043 585
R12681 GND.n2390 GND.n2038 585
R12682 GND.n3613 GND.n2390 585
R12683 GND.n8546 GND.n2037 585
R12684 GND.n2401 GND.n2037 585
R12685 GND.n8547 GND.n2036 585
R12686 GND.n3603 GND.n2036 585
R12687 GND.n8548 GND.n2035 585
R12688 GND.n3590 GND.n2035 585
R12689 GND.n2408 GND.n2030 585
R12690 GND.n3593 GND.n2408 585
R12691 GND.n8552 GND.n2029 585
R12692 GND.n3588 GND.n2029 585
R12693 GND.n8553 GND.n2028 585
R12694 GND.n2423 GND.n2028 585
R12695 GND.n8554 GND.n2027 585
R12696 GND.n3578 GND.n2027 585
R12697 GND.n3564 GND.n2022 585
R12698 GND.n3565 GND.n3564 585
R12699 GND.n8558 GND.n2021 585
R12700 GND.n3568 GND.n2021 585
R12701 GND.n8559 GND.n2020 585
R12702 GND.n3562 GND.n2020 585
R12703 GND.n8560 GND.n2019 585
R12704 GND.n2445 GND.n2019 585
R12705 GND.n2441 GND.n2014 585
R12706 GND.n3552 GND.n2441 585
R12707 GND.n8564 GND.n2013 585
R12708 GND.n3538 GND.n2013 585
R12709 GND.n8565 GND.n2012 585
R12710 GND.n3542 GND.n2012 585
R12711 GND.n8566 GND.n2011 585
R12712 GND.n3536 GND.n2011 585
R12713 GND.n2465 GND.n2006 585
R12714 GND.n2466 GND.n2465 585
R12715 GND.n8570 GND.n2005 585
R12716 GND.n3526 GND.n2005 585
R12717 GND.n8571 GND.n2004 585
R12718 GND.n3513 GND.n2004 585
R12719 GND.n8572 GND.n2003 585
R12720 GND.n3516 GND.n2003 585
R12721 GND.n2477 GND.n1998 585
R12722 GND.n3510 GND.n2477 585
R12723 GND.n8576 GND.n1997 585
R12724 GND.n2488 GND.n1997 585
R12725 GND.n8577 GND.n1996 585
R12726 GND.n3500 GND.n1996 585
R12727 GND.n8578 GND.n1995 585
R12728 GND.n3461 GND.n1995 585
R12729 GND.n2650 GND.n1990 585
R12730 GND.n3458 GND.n2650 585
R12731 GND.n8582 GND.n1989 585
R12732 GND.n2531 GND.n1989 585
R12733 GND.n8583 GND.n1988 585
R12734 GND.n3470 GND.n1988 585
R12735 GND.n8584 GND.n1987 585
R12736 GND.n3473 GND.n1987 585
R12737 GND.n2517 GND.n1982 585
R12738 GND.n3478 GND.n2517 585
R12739 GND.n8588 GND.n1981 585
R12740 GND.n2516 GND.n1981 585
R12741 GND.n8589 GND.n1980 585
R12742 GND.n2509 GND.n1980 585
R12743 GND.n8590 GND.n1979 585
R12744 GND.n3487 GND.n1979 585
R12745 GND.n2502 GND.n1974 585
R12746 GND.n3490 GND.n2502 585
R12747 GND.n8594 GND.n1973 585
R12748 GND.n3064 GND.n1973 585
R12749 GND.n8595 GND.n1972 585
R12750 GND.n3430 GND.n1972 585
R12751 GND.n8596 GND.n1971 585
R12752 GND.n3419 GND.n1971 585
R12753 GND.n2670 GND.n1966 585
R12754 GND.n3422 GND.n2670 585
R12755 GND.n8600 GND.n1965 585
R12756 GND.n3417 GND.n1965 585
R12757 GND.n8601 GND.n1964 585
R12758 GND.n2686 GND.n1964 585
R12759 GND.n8602 GND.n1963 585
R12760 GND.n3408 GND.n1963 585
R12761 GND.n3394 GND.n1958 585
R12762 GND.n3395 GND.n3394 585
R12763 GND.n8606 GND.n1957 585
R12764 GND.n3398 GND.n1957 585
R12765 GND.n8607 GND.n1956 585
R12766 GND.n3392 GND.n1956 585
R12767 GND.n8608 GND.n1955 585
R12768 GND.n2709 GND.n1955 585
R12769 GND.n2705 GND.n1950 585
R12770 GND.n3383 GND.n2705 585
R12771 GND.n8612 GND.n1949 585
R12772 GND.n3369 GND.n1949 585
R12773 GND.n8613 GND.n1948 585
R12774 GND.n3373 GND.n1948 585
R12775 GND.n8614 GND.n1947 585
R12776 GND.n3367 GND.n1947 585
R12777 GND.n2730 GND.n1942 585
R12778 GND.n2731 GND.n2730 585
R12779 GND.n8618 GND.n1941 585
R12780 GND.n3358 GND.n1941 585
R12781 GND.n8619 GND.n1940 585
R12782 GND.n3345 GND.n1940 585
R12783 GND.n8620 GND.n1939 585
R12784 GND.n3348 GND.n1939 585
R12785 GND.n2742 GND.n1934 585
R12786 GND.n3342 GND.n2742 585
R12787 GND.n8624 GND.n1933 585
R12788 GND.n2754 GND.n1933 585
R12789 GND.n8625 GND.n1932 585
R12790 GND.n3333 GND.n1932 585
R12791 GND.n8626 GND.n1931 585
R12792 GND.n3320 GND.n1931 585
R12793 GND.n2761 GND.n1926 585
R12794 GND.n3323 GND.n2761 585
R12795 GND.n8630 GND.n1925 585
R12796 GND.n3318 GND.n1925 585
R12797 GND.n8631 GND.n1924 585
R12798 GND.n2777 GND.n1924 585
R12799 GND.n8632 GND.n1923 585
R12800 GND.n3309 GND.n1923 585
R12801 GND.n3295 GND.n1918 585
R12802 GND.n3296 GND.n3295 585
R12803 GND.n8636 GND.n1917 585
R12804 GND.n3299 GND.n1917 585
R12805 GND.n8637 GND.n1916 585
R12806 GND.n3293 GND.n1916 585
R12807 GND.n8638 GND.n1915 585
R12808 GND.n2800 GND.n1915 585
R12809 GND.n2796 GND.n1910 585
R12810 GND.n3284 GND.n2796 585
R12811 GND.n8642 GND.n1909 585
R12812 GND.n3270 GND.n1909 585
R12813 GND.n8643 GND.n1908 585
R12814 GND.n3274 GND.n1908 585
R12815 GND.n8644 GND.n1907 585
R12816 GND.n3268 GND.n1907 585
R12817 GND.n2821 GND.n1902 585
R12818 GND.n2822 GND.n2821 585
R12819 GND.n8648 GND.n1901 585
R12820 GND.n3259 GND.n1901 585
R12821 GND.n8649 GND.n1900 585
R12822 GND.n3246 GND.n1900 585
R12823 GND.n8650 GND.n1899 585
R12824 GND.n3249 GND.n1899 585
R12825 GND.n2833 GND.n1894 585
R12826 GND.n3243 GND.n2833 585
R12827 GND.n8654 GND.n1893 585
R12828 GND.n2845 GND.n1893 585
R12829 GND.n8655 GND.n1892 585
R12830 GND.n3234 GND.n1892 585
R12831 GND.n8656 GND.n1891 585
R12832 GND.n3221 GND.n1891 585
R12833 GND.n2852 GND.n1886 585
R12834 GND.n3224 GND.n2852 585
R12835 GND.n8660 GND.n1885 585
R12836 GND.n3219 GND.n1885 585
R12837 GND.n8661 GND.n1884 585
R12838 GND.n2868 GND.n1884 585
R12839 GND.n8662 GND.n1883 585
R12840 GND.n3210 GND.n1883 585
R12841 GND.n3196 GND.n1878 585
R12842 GND.n3197 GND.n3196 585
R12843 GND.n8666 GND.n1877 585
R12844 GND.n3200 GND.n1877 585
R12845 GND.n8667 GND.n1876 585
R12846 GND.n3194 GND.n1876 585
R12847 GND.n8668 GND.n1875 585
R12848 GND.n2891 GND.n1875 585
R12849 GND.n2887 GND.n1870 585
R12850 GND.n3185 GND.n2887 585
R12851 GND.n8672 GND.n1869 585
R12852 GND.n3171 GND.n1869 585
R12853 GND.n8673 GND.n1868 585
R12854 GND.n3175 GND.n1868 585
R12855 GND.n8674 GND.n1867 585
R12856 GND.n3169 GND.n1867 585
R12857 GND.n3151 GND.n1862 585
R12858 GND.n3152 GND.n3151 585
R12859 GND.n8678 GND.n1861 585
R12860 GND.n3160 GND.n1861 585
R12861 GND.n8679 GND.n1860 585
R12862 GND.n2964 GND.n1860 585
R12863 GND.n8680 GND.n1837 585
R12864 GND.n8684 GND.n1837 585
R12865 GND.n2906 GND.n1859 585
R12866 GND.n2907 GND.n2906 585
R12867 GND.n1858 GND.n1818 585
R12868 GND.n8690 GND.n1818 585
R12869 GND.n1849 GND.n1846 585
R12870 GND.n1849 GND.n1817 585
R12871 GND.n1851 GND.n1850 585
R12872 GND.n1850 GND.n1805 585
R12873 GND.n1848 GND.n1803 585
R12874 GND.n8698 GND.n1803 585
R12875 GND.n10914 GND.n10913 585
R12876 GND.n10913 GND.n10912 585
R12877 GND.n10915 GND.n439 585
R12878 GND.n10905 GND.n439 585
R12879 GND.n10917 GND.n10916 585
R12880 GND.n10918 GND.n10917 585
R12881 GND.n424 GND.n423 585
R12882 GND.n7166 GND.n424 585
R12883 GND.n10926 GND.n10925 585
R12884 GND.n10925 GND.n10924 585
R12885 GND.n10927 GND.n418 585
R12886 GND.n7172 GND.n418 585
R12887 GND.n10929 GND.n10928 585
R12888 GND.n10930 GND.n10929 585
R12889 GND.n403 GND.n402 585
R12890 GND.n7178 GND.n403 585
R12891 GND.n10938 GND.n10937 585
R12892 GND.n10937 GND.n10936 585
R12893 GND.n10939 GND.n397 585
R12894 GND.n7184 GND.n397 585
R12895 GND.n10941 GND.n10940 585
R12896 GND.n10942 GND.n10941 585
R12897 GND.n382 GND.n381 585
R12898 GND.n7190 GND.n382 585
R12899 GND.n10950 GND.n10949 585
R12900 GND.n10949 GND.n10948 585
R12901 GND.n10951 GND.n376 585
R12902 GND.n7196 GND.n376 585
R12903 GND.n10953 GND.n10952 585
R12904 GND.n10954 GND.n10953 585
R12905 GND.n361 GND.n360 585
R12906 GND.n7202 GND.n361 585
R12907 GND.n10962 GND.n10961 585
R12908 GND.n10961 GND.n10960 585
R12909 GND.n10963 GND.n355 585
R12910 GND.n7208 GND.n355 585
R12911 GND.n10965 GND.n10964 585
R12912 GND.n10966 GND.n10965 585
R12913 GND.n340 GND.n339 585
R12914 GND.n7214 GND.n340 585
R12915 GND.n10974 GND.n10973 585
R12916 GND.n10973 GND.n10972 585
R12917 GND.n10975 GND.n334 585
R12918 GND.n7220 GND.n334 585
R12919 GND.n10977 GND.n10976 585
R12920 GND.n10978 GND.n10977 585
R12921 GND.n319 GND.n318 585
R12922 GND.n7226 GND.n319 585
R12923 GND.n10986 GND.n10985 585
R12924 GND.n10985 GND.n10984 585
R12925 GND.n10987 GND.n313 585
R12926 GND.n7232 GND.n313 585
R12927 GND.n10989 GND.n10988 585
R12928 GND.n10990 GND.n10989 585
R12929 GND.n298 GND.n297 585
R12930 GND.n7238 GND.n298 585
R12931 GND.n10998 GND.n10997 585
R12932 GND.n10997 GND.n10996 585
R12933 GND.n10999 GND.n292 585
R12934 GND.n7244 GND.n292 585
R12935 GND.n11001 GND.n11000 585
R12936 GND.n11002 GND.n11001 585
R12937 GND.n277 GND.n276 585
R12938 GND.n7250 GND.n277 585
R12939 GND.n11010 GND.n11009 585
R12940 GND.n11009 GND.n11008 585
R12941 GND.n11011 GND.n271 585
R12942 GND.n7256 GND.n271 585
R12943 GND.n11013 GND.n11012 585
R12944 GND.n11014 GND.n11013 585
R12945 GND.n257 GND.n256 585
R12946 GND.n7262 GND.n257 585
R12947 GND.n11022 GND.n11021 585
R12948 GND.n11021 GND.n11020 585
R12949 GND.n11023 GND.n251 585
R12950 GND.n7268 GND.n251 585
R12951 GND.n11025 GND.n11024 585
R12952 GND.n11026 GND.n11025 585
R12953 GND.n236 GND.n235 585
R12954 GND.n7101 GND.n236 585
R12955 GND.n11034 GND.n11033 585
R12956 GND.n11033 GND.n11032 585
R12957 GND.n11035 GND.n230 585
R12958 GND.n7092 GND.n230 585
R12959 GND.n11037 GND.n11036 585
R12960 GND.n11038 GND.n11037 585
R12961 GND.n215 GND.n214 585
R12962 GND.n7085 GND.n215 585
R12963 GND.n11046 GND.n11045 585
R12964 GND.n11045 GND.n11044 585
R12965 GND.n11047 GND.n209 585
R12966 GND.n7077 GND.n209 585
R12967 GND.n11049 GND.n11048 585
R12968 GND.n11050 GND.n11049 585
R12969 GND.n194 GND.n193 585
R12970 GND.n7070 GND.n194 585
R12971 GND.n11058 GND.n11057 585
R12972 GND.n11057 GND.n11056 585
R12973 GND.n11059 GND.n188 585
R12974 GND.n7062 GND.n188 585
R12975 GND.n11061 GND.n11060 585
R12976 GND.n11062 GND.n11061 585
R12977 GND.n173 GND.n172 585
R12978 GND.n7055 GND.n173 585
R12979 GND.n11070 GND.n11069 585
R12980 GND.n11069 GND.n11068 585
R12981 GND.n11071 GND.n167 585
R12982 GND.n7047 GND.n167 585
R12983 GND.n11073 GND.n11072 585
R12984 GND.n11074 GND.n11073 585
R12985 GND.n152 GND.n151 585
R12986 GND.n7040 GND.n152 585
R12987 GND.n11082 GND.n11081 585
R12988 GND.n11081 GND.n11080 585
R12989 GND.n11083 GND.n146 585
R12990 GND.n7032 GND.n146 585
R12991 GND.n11085 GND.n11084 585
R12992 GND.n11086 GND.n11085 585
R12993 GND.n131 GND.n130 585
R12994 GND.n7025 GND.n131 585
R12995 GND.n11094 GND.n11093 585
R12996 GND.n11093 GND.n11092 585
R12997 GND.n11095 GND.n126 585
R12998 GND.n7017 GND.n126 585
R12999 GND.n11097 GND.n11096 585
R13000 GND.n11098 GND.n11097 585
R13001 GND.n110 GND.n108 585
R13002 GND.n7312 GND.n110 585
R13003 GND.n11106 GND.n11105 585
R13004 GND.n11105 GND.n11104 585
R13005 GND.n109 GND.n107 585
R13006 GND.n7318 GND.n109 585
R13007 GND.n6268 GND.n6267 585
R13008 GND.n6269 GND.n6268 585
R13009 GND.n99 GND.n97 585
R13010 GND.n7004 GND.n97 585
R13011 GND.n11110 GND.n11109 585
R13012 GND.n11111 GND.n11110 585
R13013 GND.n98 GND.n96 585
R13014 GND.n6995 GND.n96 585
R13015 GND.n6256 GND.n6255 585
R13016 GND.n6259 GND.n6256 585
R13017 GND.n7334 GND.n105 585
R13018 GND.n7334 GND.n7333 585
R13019 GND.n7336 GND.n7335 585
R13020 GND.n7337 GND.n7336 585
R13021 GND.n6240 GND.n6239 585
R13022 GND.n6985 GND.n6240 585
R13023 GND.n7345 GND.n7344 585
R13024 GND.n7344 GND.n7343 585
R13025 GND.n7346 GND.n6235 585
R13026 GND.n6970 GND.n6235 585
R13027 GND.n7348 GND.n7347 585
R13028 GND.n7349 GND.n7348 585
R13029 GND.n6220 GND.n6219 585
R13030 GND.n6963 GND.n6220 585
R13031 GND.n7357 GND.n7356 585
R13032 GND.n7356 GND.n7355 585
R13033 GND.n7358 GND.n6214 585
R13034 GND.n6955 GND.n6214 585
R13035 GND.n7360 GND.n7359 585
R13036 GND.n7361 GND.n7360 585
R13037 GND.n6199 GND.n6198 585
R13038 GND.n6948 GND.n6199 585
R13039 GND.n7369 GND.n7368 585
R13040 GND.n7368 GND.n7367 585
R13041 GND.n7370 GND.n6193 585
R13042 GND.n6940 GND.n6193 585
R13043 GND.n7372 GND.n7371 585
R13044 GND.n7373 GND.n7372 585
R13045 GND.n6178 GND.n6177 585
R13046 GND.n6933 GND.n6178 585
R13047 GND.n7381 GND.n7380 585
R13048 GND.n7380 GND.n7379 585
R13049 GND.n7382 GND.n6172 585
R13050 GND.n6925 GND.n6172 585
R13051 GND.n7384 GND.n7383 585
R13052 GND.n7385 GND.n7384 585
R13053 GND.n6158 GND.n6157 585
R13054 GND.n6918 GND.n6158 585
R13055 GND.n7393 GND.n7392 585
R13056 GND.n7392 GND.n7391 585
R13057 GND.n7394 GND.n6152 585
R13058 GND.n6910 GND.n6152 585
R13059 GND.n7396 GND.n7395 585
R13060 GND.n7397 GND.n7396 585
R13061 GND.n6137 GND.n6136 585
R13062 GND.n6903 GND.n6137 585
R13063 GND.n7405 GND.n7404 585
R13064 GND.n7404 GND.n7403 585
R13065 GND.n7406 GND.n6131 585
R13066 GND.n6895 GND.n6131 585
R13067 GND.n7408 GND.n7407 585
R13068 GND.n7409 GND.n7408 585
R13069 GND.n6116 GND.n6115 585
R13070 GND.n6888 GND.n6116 585
R13071 GND.n7417 GND.n7416 585
R13072 GND.n7416 GND.n7415 585
R13073 GND.n7418 GND.n6110 585
R13074 GND.n6880 GND.n6110 585
R13075 GND.n7420 GND.n7419 585
R13076 GND.n7421 GND.n7420 585
R13077 GND.n6095 GND.n6094 585
R13078 GND.n6873 GND.n6095 585
R13079 GND.n7429 GND.n7428 585
R13080 GND.n7428 GND.n7427 585
R13081 GND.n7430 GND.n6089 585
R13082 GND.n6865 GND.n6089 585
R13083 GND.n7432 GND.n7431 585
R13084 GND.n7433 GND.n7432 585
R13085 GND.n6074 GND.n6073 585
R13086 GND.n6858 GND.n6074 585
R13087 GND.n7441 GND.n7440 585
R13088 GND.n7440 GND.n7439 585
R13089 GND.n7442 GND.n6068 585
R13090 GND.n6850 GND.n6068 585
R13091 GND.n7444 GND.n7443 585
R13092 GND.n7445 GND.n7444 585
R13093 GND.n6053 GND.n6052 585
R13094 GND.n6843 GND.n6053 585
R13095 GND.n7453 GND.n7452 585
R13096 GND.n7452 GND.n7451 585
R13097 GND.n7454 GND.n6047 585
R13098 GND.n6835 GND.n6047 585
R13099 GND.n7456 GND.n7455 585
R13100 GND.n7457 GND.n7456 585
R13101 GND.n6033 GND.n6032 585
R13102 GND.n6828 GND.n6033 585
R13103 GND.n7465 GND.n7464 585
R13104 GND.n7464 GND.n7463 585
R13105 GND.n7466 GND.n6027 585
R13106 GND.n6820 GND.n6027 585
R13107 GND.n7468 GND.n7467 585
R13108 GND.n7469 GND.n7468 585
R13109 GND.n6012 GND.n6011 585
R13110 GND.n6813 GND.n6012 585
R13111 GND.n7477 GND.n7476 585
R13112 GND.n7476 GND.n7475 585
R13113 GND.n7478 GND.n6006 585
R13114 GND.n6805 GND.n6006 585
R13115 GND.n7480 GND.n7479 585
R13116 GND.n7481 GND.n7480 585
R13117 GND.n5991 GND.n5990 585
R13118 GND.n6798 GND.n5991 585
R13119 GND.n7489 GND.n7488 585
R13120 GND.n7488 GND.n7487 585
R13121 GND.n7490 GND.n5985 585
R13122 GND.n6790 GND.n5985 585
R13123 GND.n7492 GND.n7491 585
R13124 GND.n7493 GND.n7492 585
R13125 GND.n5970 GND.n5969 585
R13126 GND.n6783 GND.n5970 585
R13127 GND.n7501 GND.n7500 585
R13128 GND.n7500 GND.n7499 585
R13129 GND.n7502 GND.n5964 585
R13130 GND.n6775 GND.n5964 585
R13131 GND.n7504 GND.n7503 585
R13132 GND.n7505 GND.n7504 585
R13133 GND.n5950 GND.n5949 585
R13134 GND.n6768 GND.n5950 585
R13135 GND.n7513 GND.n7512 585
R13136 GND.n7512 GND.n7511 585
R13137 GND.n7514 GND.n5944 585
R13138 GND.n6760 GND.n5944 585
R13139 GND.n7516 GND.n7515 585
R13140 GND.n7517 GND.n7516 585
R13141 GND.n5928 GND.n5927 585
R13142 GND.n6753 GND.n5928 585
R13143 GND.n7525 GND.n7524 585
R13144 GND.n7524 GND.n7523 585
R13145 GND.n7526 GND.n5921 585
R13146 GND.n6745 GND.n5921 585
R13147 GND.n7528 GND.n7527 585
R13148 GND.n7529 GND.n7528 585
R13149 GND.n5922 GND.n4605 585
R13150 GND.n7532 GND.n4605 585
R13151 GND.n7645 GND.n7644 585
R13152 GND.n7643 GND.n4604 585
R13153 GND.n7642 GND.n4603 585
R13154 GND.n7647 GND.n4603 585
R13155 GND.n7641 GND.n7640 585
R13156 GND.n7639 GND.n7638 585
R13157 GND.n7637 GND.n7636 585
R13158 GND.n7635 GND.n7634 585
R13159 GND.n7633 GND.n7632 585
R13160 GND.n7631 GND.n7630 585
R13161 GND.n7629 GND.n7628 585
R13162 GND.n7627 GND.n7626 585
R13163 GND.n7625 GND.n7624 585
R13164 GND.n7623 GND.n4618 585
R13165 GND.n7622 GND.n7621 585
R13166 GND.n7620 GND.n7619 585
R13167 GND.n7618 GND.n7617 585
R13168 GND.n7616 GND.n7615 585
R13169 GND.n7614 GND.n7613 585
R13170 GND.n7612 GND.n7611 585
R13171 GND.n7610 GND.n7609 585
R13172 GND.n7608 GND.n7607 585
R13173 GND.n7606 GND.n7605 585
R13174 GND.n7604 GND.n7603 585
R13175 GND.n7602 GND.n7601 585
R13176 GND.n7600 GND.n7599 585
R13177 GND.n7598 GND.n7597 585
R13178 GND.n7597 GND.n4792 585
R13179 GND.n7596 GND.n7595 585
R13180 GND.n7594 GND.n7593 585
R13181 GND.n7592 GND.n7591 585
R13182 GND.n7590 GND.n7589 585
R13183 GND.n7588 GND.n7587 585
R13184 GND.n7586 GND.n7585 585
R13185 GND.n7584 GND.n7583 585
R13186 GND.n7582 GND.n7581 585
R13187 GND.n7580 GND.n7579 585
R13188 GND.n7578 GND.n7577 585
R13189 GND.n7576 GND.n7575 585
R13190 GND.n7574 GND.n7573 585
R13191 GND.n7572 GND.n7571 585
R13192 GND.n7570 GND.n7569 585
R13193 GND.n7568 GND.n7567 585
R13194 GND.n7566 GND.n7565 585
R13195 GND.n7564 GND.n7563 585
R13196 GND.n7562 GND.n7561 585
R13197 GND.n7560 GND.n7559 585
R13198 GND.n7558 GND.n7557 585
R13199 GND.n7556 GND.n7555 585
R13200 GND.n7554 GND.n7553 585
R13201 GND.n7552 GND.n7551 585
R13202 GND.n7550 GND.n7549 585
R13203 GND.n7548 GND.n7547 585
R13204 GND.n7546 GND.n7545 585
R13205 GND.n7544 GND.n7543 585
R13206 GND.n7542 GND.n7541 585
R13207 GND.n7540 GND.n7539 585
R13208 GND.n5877 GND.n4827 585
R13209 GND.n10783 GND.n10782 585
R13210 GND.n10789 GND.n10788 585
R13211 GND.n10791 GND.n10790 585
R13212 GND.n10793 GND.n10792 585
R13213 GND.n10795 GND.n10794 585
R13214 GND.n10797 GND.n10796 585
R13215 GND.n10799 GND.n10798 585
R13216 GND.n10801 GND.n10800 585
R13217 GND.n10803 GND.n10802 585
R13218 GND.n10805 GND.n10804 585
R13219 GND.n10807 GND.n10806 585
R13220 GND.n10809 GND.n10808 585
R13221 GND.n10811 GND.n10810 585
R13222 GND.n10813 GND.n10812 585
R13223 GND.n10815 GND.n10814 585
R13224 GND.n10817 GND.n10816 585
R13225 GND.n10819 GND.n10818 585
R13226 GND.n10821 GND.n10820 585
R13227 GND.n10823 GND.n10822 585
R13228 GND.n10825 GND.n10824 585
R13229 GND.n10827 GND.n10826 585
R13230 GND.n10829 GND.n10828 585
R13231 GND.n10831 GND.n10830 585
R13232 GND.n10833 GND.n10832 585
R13233 GND.n10835 GND.n10834 585
R13234 GND.n10837 GND.n10836 585
R13235 GND.n10839 GND.n10838 585
R13236 GND.n10841 GND.n10840 585
R13237 GND.n10843 GND.n10842 585
R13238 GND.n10845 GND.n10844 585
R13239 GND.n10847 GND.n10846 585
R13240 GND.n10849 GND.n10848 585
R13241 GND.n10851 GND.n10850 585
R13242 GND.n10853 GND.n10852 585
R13243 GND.n10855 GND.n10854 585
R13244 GND.n10857 GND.n10856 585
R13245 GND.n10859 GND.n10858 585
R13246 GND.n10861 GND.n10860 585
R13247 GND.n10863 GND.n10862 585
R13248 GND.n10865 GND.n10864 585
R13249 GND.n10867 GND.n10866 585
R13250 GND.n10869 GND.n10868 585
R13251 GND.n10871 GND.n10870 585
R13252 GND.n10734 GND.n10731 585
R13253 GND.n10875 GND.n10735 585
R13254 GND.n10877 GND.n10876 585
R13255 GND.n10879 GND.n10878 585
R13256 GND.n10881 GND.n10880 585
R13257 GND.n10883 GND.n10882 585
R13258 GND.n10885 GND.n10884 585
R13259 GND.n10887 GND.n10886 585
R13260 GND.n10889 GND.n10888 585
R13261 GND.n10891 GND.n10890 585
R13262 GND.n10892 GND.n10716 585
R13263 GND.n10894 GND.n10893 585
R13264 GND.n10717 GND.n10715 585
R13265 GND.n10718 GND.n444 585
R13266 GND.n10896 GND.n444 585
R13267 GND.n10908 GND.n446 585
R13268 GND.n10912 GND.n446 585
R13269 GND.n10907 GND.n10906 585
R13270 GND.n10906 GND.n10905 585
R13271 GND.n452 GND.n436 585
R13272 GND.n10918 GND.n436 585
R13273 GND.n7165 GND.n7164 585
R13274 GND.n7166 GND.n7165 585
R13275 GND.n7158 GND.n426 585
R13276 GND.n10924 GND.n426 585
R13277 GND.n7174 GND.n7173 585
R13278 GND.n7173 GND.n7172 585
R13279 GND.n7175 GND.n415 585
R13280 GND.n10930 GND.n415 585
R13281 GND.n7177 GND.n7176 585
R13282 GND.n7178 GND.n7177 585
R13283 GND.n7151 GND.n405 585
R13284 GND.n10936 GND.n405 585
R13285 GND.n7186 GND.n7185 585
R13286 GND.n7185 GND.n7184 585
R13287 GND.n7187 GND.n394 585
R13288 GND.n10942 GND.n394 585
R13289 GND.n7189 GND.n7188 585
R13290 GND.n7190 GND.n7189 585
R13291 GND.n7144 GND.n384 585
R13292 GND.n10948 GND.n384 585
R13293 GND.n7198 GND.n7197 585
R13294 GND.n7197 GND.n7196 585
R13295 GND.n7199 GND.n373 585
R13296 GND.n10954 GND.n373 585
R13297 GND.n7201 GND.n7200 585
R13298 GND.n7202 GND.n7201 585
R13299 GND.n7137 GND.n363 585
R13300 GND.n10960 GND.n363 585
R13301 GND.n7210 GND.n7209 585
R13302 GND.n7209 GND.n7208 585
R13303 GND.n7211 GND.n352 585
R13304 GND.n10966 GND.n352 585
R13305 GND.n7213 GND.n7212 585
R13306 GND.n7214 GND.n7213 585
R13307 GND.n7130 GND.n342 585
R13308 GND.n10972 GND.n342 585
R13309 GND.n7222 GND.n7221 585
R13310 GND.n7221 GND.n7220 585
R13311 GND.n7223 GND.n331 585
R13312 GND.n10978 GND.n331 585
R13313 GND.n7225 GND.n7224 585
R13314 GND.n7226 GND.n7225 585
R13315 GND.n7123 GND.n321 585
R13316 GND.n10984 GND.n321 585
R13317 GND.n7234 GND.n7233 585
R13318 GND.n7233 GND.n7232 585
R13319 GND.n7235 GND.n310 585
R13320 GND.n10990 GND.n310 585
R13321 GND.n7237 GND.n7236 585
R13322 GND.n7238 GND.n7237 585
R13323 GND.n7116 GND.n300 585
R13324 GND.n10996 GND.n300 585
R13325 GND.n7246 GND.n7245 585
R13326 GND.n7245 GND.n7244 585
R13327 GND.n7247 GND.n289 585
R13328 GND.n11002 GND.n289 585
R13329 GND.n7249 GND.n7248 585
R13330 GND.n7250 GND.n7249 585
R13331 GND.n7109 GND.n279 585
R13332 GND.n11008 GND.n279 585
R13333 GND.n7258 GND.n7257 585
R13334 GND.n7257 GND.n7256 585
R13335 GND.n7259 GND.n268 585
R13336 GND.n11014 GND.n268 585
R13337 GND.n7261 GND.n7260 585
R13338 GND.n7262 GND.n7261 585
R13339 GND.n7107 GND.n258 585
R13340 GND.n11020 GND.n258 585
R13341 GND.n7106 GND.n6434 585
R13342 GND.n7268 GND.n6434 585
R13343 GND.n7104 GND.n248 585
R13344 GND.n11026 GND.n248 585
R13345 GND.n7103 GND.n7102 585
R13346 GND.n7102 GND.n7101 585
R13347 GND.n6440 GND.n238 585
R13348 GND.n11032 GND.n238 585
R13349 GND.n7091 GND.n7090 585
R13350 GND.n7092 GND.n7091 585
R13351 GND.n7088 GND.n227 585
R13352 GND.n11038 GND.n227 585
R13353 GND.n7087 GND.n7086 585
R13354 GND.n7086 GND.n7085 585
R13355 GND.n6444 GND.n217 585
R13356 GND.n11044 GND.n217 585
R13357 GND.n7076 GND.n7075 585
R13358 GND.n7077 GND.n7076 585
R13359 GND.n7073 GND.n206 585
R13360 GND.n11050 GND.n206 585
R13361 GND.n7072 GND.n7071 585
R13362 GND.n7071 GND.n7070 585
R13363 GND.n6448 GND.n196 585
R13364 GND.n11056 GND.n196 585
R13365 GND.n7061 GND.n7060 585
R13366 GND.n7062 GND.n7061 585
R13367 GND.n7058 GND.n185 585
R13368 GND.n11062 GND.n185 585
R13369 GND.n7057 GND.n7056 585
R13370 GND.n7056 GND.n7055 585
R13371 GND.n6452 GND.n175 585
R13372 GND.n11068 GND.n175 585
R13373 GND.n7046 GND.n7045 585
R13374 GND.n7047 GND.n7046 585
R13375 GND.n7043 GND.n164 585
R13376 GND.n11074 GND.n164 585
R13377 GND.n7042 GND.n7041 585
R13378 GND.n7041 GND.n7040 585
R13379 GND.n6456 GND.n154 585
R13380 GND.n11080 GND.n154 585
R13381 GND.n7031 GND.n7030 585
R13382 GND.n7032 GND.n7031 585
R13383 GND.n7028 GND.n143 585
R13384 GND.n11086 GND.n143 585
R13385 GND.n7027 GND.n7026 585
R13386 GND.n7026 GND.n7025 585
R13387 GND.n6460 GND.n133 585
R13388 GND.n11092 GND.n133 585
R13389 GND.n7016 GND.n7015 585
R13390 GND.n7017 GND.n7016 585
R13391 GND.n7013 GND.n123 585
R13392 GND.n11098 GND.n123 585
R13393 GND.n7012 GND.n6278 585
R13394 GND.n7312 GND.n6278 585
R13395 GND.n7011 GND.n112 585
R13396 GND.n11104 GND.n112 585
R13397 GND.n7010 GND.n6270 585
R13398 GND.n7318 GND.n6270 585
R13399 GND.n6466 GND.n6463 585
R13400 GND.n6466 GND.n6269 585
R13401 GND.n7002 GND.n7001 585
R13402 GND.n7004 GND.n7002 585
R13403 GND.n7000 GND.n93 585
R13404 GND.n11111 GND.n93 585
R13405 GND.n6994 GND.n6467 585
R13406 GND.n6995 GND.n6994 585
R13407 GND.n6993 GND.n6992 585
R13408 GND.n6993 GND.n6259 585
R13409 GND.n6989 GND.n6257 585
R13410 GND.n7333 GND.n6257 585
R13411 GND.n6988 GND.n6252 585
R13412 GND.n7337 GND.n6252 585
R13413 GND.n6987 GND.n6986 585
R13414 GND.n6986 GND.n6985 585
R13415 GND.n6472 GND.n6242 585
R13416 GND.n7343 GND.n6242 585
R13417 GND.n6969 GND.n6968 585
R13418 GND.n6970 GND.n6969 585
R13419 GND.n6966 GND.n6232 585
R13420 GND.n7349 GND.n6232 585
R13421 GND.n6965 GND.n6964 585
R13422 GND.n6964 GND.n6963 585
R13423 GND.n6476 GND.n6222 585
R13424 GND.n7355 GND.n6222 585
R13425 GND.n6954 GND.n6953 585
R13426 GND.n6955 GND.n6954 585
R13427 GND.n6951 GND.n6211 585
R13428 GND.n7361 GND.n6211 585
R13429 GND.n6950 GND.n6949 585
R13430 GND.n6949 GND.n6948 585
R13431 GND.n6480 GND.n6201 585
R13432 GND.n7367 GND.n6201 585
R13433 GND.n6939 GND.n6938 585
R13434 GND.n6940 GND.n6939 585
R13435 GND.n6936 GND.n6190 585
R13436 GND.n7373 GND.n6190 585
R13437 GND.n6935 GND.n6934 585
R13438 GND.n6934 GND.n6933 585
R13439 GND.n6484 GND.n6180 585
R13440 GND.n7379 GND.n6180 585
R13441 GND.n6924 GND.n6923 585
R13442 GND.n6925 GND.n6924 585
R13443 GND.n6921 GND.n6170 585
R13444 GND.n7385 GND.n6170 585
R13445 GND.n6920 GND.n6919 585
R13446 GND.n6919 GND.n6918 585
R13447 GND.n6489 GND.n6160 585
R13448 GND.n7391 GND.n6160 585
R13449 GND.n6909 GND.n6908 585
R13450 GND.n6910 GND.n6909 585
R13451 GND.n6906 GND.n6149 585
R13452 GND.n7397 GND.n6149 585
R13453 GND.n6905 GND.n6904 585
R13454 GND.n6904 GND.n6903 585
R13455 GND.n6493 GND.n6139 585
R13456 GND.n7403 GND.n6139 585
R13457 GND.n6894 GND.n6893 585
R13458 GND.n6895 GND.n6894 585
R13459 GND.n6891 GND.n6128 585
R13460 GND.n7409 GND.n6128 585
R13461 GND.n6890 GND.n6889 585
R13462 GND.n6889 GND.n6888 585
R13463 GND.n6497 GND.n6118 585
R13464 GND.n7415 GND.n6118 585
R13465 GND.n6879 GND.n6878 585
R13466 GND.n6880 GND.n6879 585
R13467 GND.n6876 GND.n6107 585
R13468 GND.n7421 GND.n6107 585
R13469 GND.n6875 GND.n6874 585
R13470 GND.n6874 GND.n6873 585
R13471 GND.n6501 GND.n6097 585
R13472 GND.n7427 GND.n6097 585
R13473 GND.n6864 GND.n6863 585
R13474 GND.n6865 GND.n6864 585
R13475 GND.n6861 GND.n6086 585
R13476 GND.n7433 GND.n6086 585
R13477 GND.n6860 GND.n6859 585
R13478 GND.n6859 GND.n6858 585
R13479 GND.n6505 GND.n6076 585
R13480 GND.n7439 GND.n6076 585
R13481 GND.n6849 GND.n6848 585
R13482 GND.n6850 GND.n6849 585
R13483 GND.n6846 GND.n6065 585
R13484 GND.n7445 GND.n6065 585
R13485 GND.n6845 GND.n6844 585
R13486 GND.n6844 GND.n6843 585
R13487 GND.n6509 GND.n6055 585
R13488 GND.n7451 GND.n6055 585
R13489 GND.n6834 GND.n6833 585
R13490 GND.n6835 GND.n6834 585
R13491 GND.n6831 GND.n6044 585
R13492 GND.n7457 GND.n6044 585
R13493 GND.n6830 GND.n6829 585
R13494 GND.n6829 GND.n6828 585
R13495 GND.n6513 GND.n6035 585
R13496 GND.n7463 GND.n6035 585
R13497 GND.n6819 GND.n6818 585
R13498 GND.n6820 GND.n6819 585
R13499 GND.n6816 GND.n6024 585
R13500 GND.n7469 GND.n6024 585
R13501 GND.n6815 GND.n6814 585
R13502 GND.n6814 GND.n6813 585
R13503 GND.n6518 GND.n6014 585
R13504 GND.n7475 GND.n6014 585
R13505 GND.n6804 GND.n6803 585
R13506 GND.n6805 GND.n6804 585
R13507 GND.n6801 GND.n6003 585
R13508 GND.n7481 GND.n6003 585
R13509 GND.n6800 GND.n6799 585
R13510 GND.n6799 GND.n6798 585
R13511 GND.n6522 GND.n5993 585
R13512 GND.n7487 GND.n5993 585
R13513 GND.n6789 GND.n6788 585
R13514 GND.n6790 GND.n6789 585
R13515 GND.n6786 GND.n5982 585
R13516 GND.n7493 GND.n5982 585
R13517 GND.n6785 GND.n6784 585
R13518 GND.n6784 GND.n6783 585
R13519 GND.n6526 GND.n5972 585
R13520 GND.n7499 GND.n5972 585
R13521 GND.n6774 GND.n6773 585
R13522 GND.n6775 GND.n6774 585
R13523 GND.n6771 GND.n5961 585
R13524 GND.n7505 GND.n5961 585
R13525 GND.n6770 GND.n6769 585
R13526 GND.n6769 GND.n6768 585
R13527 GND.n6530 GND.n5952 585
R13528 GND.n7511 GND.n5952 585
R13529 GND.n6759 GND.n6758 585
R13530 GND.n6760 GND.n6759 585
R13531 GND.n6756 GND.n5941 585
R13532 GND.n7517 GND.n5941 585
R13533 GND.n6755 GND.n6754 585
R13534 GND.n6754 GND.n6753 585
R13535 GND.n6736 GND.n5930 585
R13536 GND.n7523 GND.n5930 585
R13537 GND.n6744 GND.n6743 585
R13538 GND.n6745 GND.n6744 585
R13539 GND.n5878 GND.n5876 585
R13540 GND.n7529 GND.n5878 585
R13541 GND.n7534 GND.n7533 585
R13542 GND.n7533 GND.n7532 585
R13543 GND.n573 GND.n572 585
R13544 GND.n10535 GND.n573 585
R13545 GND.n10538 GND.n10537 585
R13546 GND.n10537 GND.n10536 585
R13547 GND.n10539 GND.n567 585
R13548 GND.n567 GND.n566 585
R13549 GND.n10541 GND.n10540 585
R13550 GND.n10542 GND.n10541 585
R13551 GND.n565 GND.n564 585
R13552 GND.n10543 GND.n565 585
R13553 GND.n10546 GND.n10545 585
R13554 GND.n10545 GND.n10544 585
R13555 GND.n10547 GND.n559 585
R13556 GND.n559 GND.n558 585
R13557 GND.n10549 GND.n10548 585
R13558 GND.n10550 GND.n10549 585
R13559 GND.n557 GND.n556 585
R13560 GND.n10551 GND.n557 585
R13561 GND.n10554 GND.n10553 585
R13562 GND.n10553 GND.n10552 585
R13563 GND.n10555 GND.n551 585
R13564 GND.n551 GND.n550 585
R13565 GND.n10557 GND.n10556 585
R13566 GND.n10558 GND.n10557 585
R13567 GND.n549 GND.n548 585
R13568 GND.n10559 GND.n549 585
R13569 GND.n10562 GND.n10561 585
R13570 GND.n10561 GND.n10560 585
R13571 GND.n10563 GND.n543 585
R13572 GND.n543 GND.n542 585
R13573 GND.n10565 GND.n10564 585
R13574 GND.n10566 GND.n10565 585
R13575 GND.n541 GND.n540 585
R13576 GND.n10567 GND.n541 585
R13577 GND.n10570 GND.n10569 585
R13578 GND.n10569 GND.n10568 585
R13579 GND.n10571 GND.n535 585
R13580 GND.n535 GND.n534 585
R13581 GND.n10573 GND.n10572 585
R13582 GND.n10574 GND.n10573 585
R13583 GND.n533 GND.n532 585
R13584 GND.n10575 GND.n533 585
R13585 GND.n10578 GND.n10577 585
R13586 GND.n10577 GND.n10576 585
R13587 GND.n10579 GND.n527 585
R13588 GND.n527 GND.n526 585
R13589 GND.n10581 GND.n10580 585
R13590 GND.n10582 GND.n10581 585
R13591 GND.n525 GND.n524 585
R13592 GND.n10583 GND.n525 585
R13593 GND.n10586 GND.n10585 585
R13594 GND.n10585 GND.n10584 585
R13595 GND.n10587 GND.n519 585
R13596 GND.n519 GND.n518 585
R13597 GND.n10589 GND.n10588 585
R13598 GND.n10590 GND.n10589 585
R13599 GND.n517 GND.n516 585
R13600 GND.n10591 GND.n517 585
R13601 GND.n10594 GND.n10593 585
R13602 GND.n10593 GND.n10592 585
R13603 GND.n10595 GND.n511 585
R13604 GND.n511 GND.n510 585
R13605 GND.n10597 GND.n10596 585
R13606 GND.n10598 GND.n10597 585
R13607 GND.n509 GND.n508 585
R13608 GND.n10599 GND.n509 585
R13609 GND.n10602 GND.n10601 585
R13610 GND.n10601 GND.n10600 585
R13611 GND.n10603 GND.n503 585
R13612 GND.n503 GND.n502 585
R13613 GND.n10605 GND.n10604 585
R13614 GND.n10606 GND.n10605 585
R13615 GND.n501 GND.n500 585
R13616 GND.n10607 GND.n501 585
R13617 GND.n10610 GND.n10609 585
R13618 GND.n10609 GND.n10608 585
R13619 GND.n10611 GND.n495 585
R13620 GND.n495 GND.n494 585
R13621 GND.n10613 GND.n10612 585
R13622 GND.n10614 GND.n10613 585
R13623 GND.n493 GND.n492 585
R13624 GND.n10615 GND.n493 585
R13625 GND.n10618 GND.n10617 585
R13626 GND.n10617 GND.n10616 585
R13627 GND.n10619 GND.n487 585
R13628 GND.n487 GND.n486 585
R13629 GND.n10621 GND.n10620 585
R13630 GND.n10622 GND.n10621 585
R13631 GND.n485 GND.n484 585
R13632 GND.n10623 GND.n485 585
R13633 GND.n10626 GND.n10625 585
R13634 GND.n10625 GND.n10624 585
R13635 GND.n10627 GND.n479 585
R13636 GND.n479 GND.n478 585
R13637 GND.n10629 GND.n10628 585
R13638 GND.n10630 GND.n10629 585
R13639 GND.n477 GND.n476 585
R13640 GND.n10631 GND.n477 585
R13641 GND.n10634 GND.n10633 585
R13642 GND.n10633 GND.n10632 585
R13643 GND.n10635 GND.n471 585
R13644 GND.n471 GND.n470 585
R13645 GND.n10637 GND.n10636 585
R13646 GND.n10638 GND.n10637 585
R13647 GND.n469 GND.n468 585
R13648 GND.n10639 GND.n469 585
R13649 GND.n10642 GND.n10641 585
R13650 GND.n10641 GND.n10640 585
R13651 GND.n10643 GND.n463 585
R13652 GND.n463 GND.n461 585
R13653 GND.n10645 GND.n10644 585
R13654 GND.n10646 GND.n10645 585
R13655 GND.n464 GND.n462 585
R13656 GND.n462 GND.n460 585
R13657 GND.n6379 GND.n6378 585
R13658 GND.n6379 GND.n448 585
R13659 GND.n6381 GND.n6380 585
R13660 GND.n6380 GND.n445 585
R13661 GND.n6382 GND.n6371 585
R13662 GND.n6371 GND.n438 585
R13663 GND.n6384 GND.n6383 585
R13664 GND.n6384 GND.n435 585
R13665 GND.n6385 GND.n6370 585
R13666 GND.n6385 GND.n428 585
R13667 GND.n6387 GND.n6386 585
R13668 GND.n6386 GND.n425 585
R13669 GND.n6388 GND.n6365 585
R13670 GND.n6365 GND.n417 585
R13671 GND.n6390 GND.n6389 585
R13672 GND.n6390 GND.n414 585
R13673 GND.n6391 GND.n6364 585
R13674 GND.n6391 GND.n407 585
R13675 GND.n6393 GND.n6392 585
R13676 GND.n6392 GND.n404 585
R13677 GND.n6394 GND.n6359 585
R13678 GND.n6359 GND.n396 585
R13679 GND.n6396 GND.n6395 585
R13680 GND.n6396 GND.n393 585
R13681 GND.n6397 GND.n6358 585
R13682 GND.n6397 GND.n386 585
R13683 GND.n6399 GND.n6398 585
R13684 GND.n6398 GND.n383 585
R13685 GND.n6400 GND.n6353 585
R13686 GND.n6353 GND.n375 585
R13687 GND.n6402 GND.n6401 585
R13688 GND.n6402 GND.n372 585
R13689 GND.n6403 GND.n6352 585
R13690 GND.n6403 GND.n365 585
R13691 GND.n6405 GND.n6404 585
R13692 GND.n6404 GND.n362 585
R13693 GND.n6406 GND.n6347 585
R13694 GND.n6347 GND.n354 585
R13695 GND.n6408 GND.n6407 585
R13696 GND.n6408 GND.n351 585
R13697 GND.n6409 GND.n6346 585
R13698 GND.n6409 GND.n344 585
R13699 GND.n6411 GND.n6410 585
R13700 GND.n6410 GND.n341 585
R13701 GND.n6412 GND.n6341 585
R13702 GND.n6341 GND.n333 585
R13703 GND.n6414 GND.n6413 585
R13704 GND.n6414 GND.n330 585
R13705 GND.n6415 GND.n6340 585
R13706 GND.n6415 GND.n323 585
R13707 GND.n6417 GND.n6416 585
R13708 GND.n6416 GND.n320 585
R13709 GND.n6418 GND.n6335 585
R13710 GND.n6335 GND.n312 585
R13711 GND.n6420 GND.n6419 585
R13712 GND.n6420 GND.n309 585
R13713 GND.n6421 GND.n6334 585
R13714 GND.n6421 GND.n302 585
R13715 GND.n6423 GND.n6422 585
R13716 GND.n6422 GND.n299 585
R13717 GND.n6424 GND.n6329 585
R13718 GND.n6329 GND.n291 585
R13719 GND.n6426 GND.n6425 585
R13720 GND.n6426 GND.n288 585
R13721 GND.n6427 GND.n6328 585
R13722 GND.n6427 GND.n281 585
R13723 GND.n6429 GND.n6428 585
R13724 GND.n6428 GND.n278 585
R13725 GND.n6430 GND.n6323 585
R13726 GND.n6323 GND.n270 585
R13727 GND.n6432 GND.n6431 585
R13728 GND.n6432 GND.n267 585
R13729 GND.n6433 GND.n6322 585
R13730 GND.n6433 GND.n260 585
R13731 GND.n7271 GND.n7270 585
R13732 GND.n7270 GND.n7269 585
R13733 GND.n7272 GND.n6317 585
R13734 GND.n6317 GND.n250 585
R13735 GND.n7274 GND.n7273 585
R13736 GND.n7274 GND.n247 585
R13737 GND.n7275 GND.n6316 585
R13738 GND.n7275 GND.n240 585
R13739 GND.n7277 GND.n7276 585
R13740 GND.n7276 GND.n237 585
R13741 GND.n7278 GND.n6311 585
R13742 GND.n6311 GND.n229 585
R13743 GND.n7280 GND.n7279 585
R13744 GND.n7280 GND.n226 585
R13745 GND.n7281 GND.n6310 585
R13746 GND.n7281 GND.n219 585
R13747 GND.n7283 GND.n7282 585
R13748 GND.n7282 GND.n216 585
R13749 GND.n7284 GND.n6305 585
R13750 GND.n6305 GND.n208 585
R13751 GND.n7286 GND.n7285 585
R13752 GND.n7286 GND.n205 585
R13753 GND.n7287 GND.n6304 585
R13754 GND.n7287 GND.n198 585
R13755 GND.n7289 GND.n7288 585
R13756 GND.n7288 GND.n195 585
R13757 GND.n7290 GND.n6299 585
R13758 GND.n6299 GND.n187 585
R13759 GND.n7292 GND.n7291 585
R13760 GND.n7292 GND.n184 585
R13761 GND.n7293 GND.n6298 585
R13762 GND.n7293 GND.n177 585
R13763 GND.n7295 GND.n7294 585
R13764 GND.n7294 GND.n174 585
R13765 GND.n7296 GND.n6293 585
R13766 GND.n6293 GND.n166 585
R13767 GND.n7298 GND.n7297 585
R13768 GND.n7298 GND.n163 585
R13769 GND.n7299 GND.n6292 585
R13770 GND.n7299 GND.n156 585
R13771 GND.n7301 GND.n7300 585
R13772 GND.n7300 GND.n153 585
R13773 GND.n7302 GND.n6287 585
R13774 GND.n6287 GND.n145 585
R13775 GND.n7304 GND.n7303 585
R13776 GND.n7304 GND.n142 585
R13777 GND.n7305 GND.n6286 585
R13778 GND.n7305 GND.n135 585
R13779 GND.n7307 GND.n7306 585
R13780 GND.n7306 GND.n132 585
R13781 GND.n7308 GND.n6280 585
R13782 GND.n6280 GND.n125 585
R13783 GND.n7310 GND.n7309 585
R13784 GND.n7311 GND.n7310 585
R13785 GND.n6282 GND.n6279 585
R13786 GND.n6279 GND.n114 585
R13787 GND.n6266 GND.n6265 585
R13788 GND.n6266 GND.n111 585
R13789 GND.n7321 GND.n7320 585
R13790 GND.n7320 GND.n7319 585
R13791 GND.n7323 GND.n6264 585
R13792 GND.n7003 GND.n6264 585
R13793 GND.n7325 GND.n7324 585
R13794 GND.n7325 GND.n94 585
R13795 GND.n7327 GND.n7326 585
R13796 GND.n7326 GND.n92 585
R13797 GND.n7328 GND.n6261 585
R13798 GND.n6471 GND.n6261 585
R13799 GND.n7331 GND.n7330 585
R13800 GND.n7332 GND.n7331 585
R13801 GND.n6262 GND.n6260 585
R13802 GND.n6260 GND.n6254 585
R13803 GND.n6645 GND.n6643 585
R13804 GND.n6643 GND.n6251 585
R13805 GND.n6647 GND.n6646 585
R13806 GND.n6647 GND.n6244 585
R13807 GND.n6648 GND.n6642 585
R13808 GND.n6648 GND.n6241 585
R13809 GND.n6650 GND.n6649 585
R13810 GND.n6649 GND.n6234 585
R13811 GND.n6651 GND.n6636 585
R13812 GND.n6636 GND.n6231 585
R13813 GND.n6653 GND.n6652 585
R13814 GND.n6653 GND.n6224 585
R13815 GND.n6654 GND.n6635 585
R13816 GND.n6654 GND.n6221 585
R13817 GND.n6656 GND.n6655 585
R13818 GND.n6655 GND.n6213 585
R13819 GND.n6657 GND.n6630 585
R13820 GND.n6630 GND.n6210 585
R13821 GND.n6659 GND.n6658 585
R13822 GND.n6659 GND.n6203 585
R13823 GND.n6660 GND.n6629 585
R13824 GND.n6660 GND.n6200 585
R13825 GND.n6662 GND.n6661 585
R13826 GND.n6661 GND.n6192 585
R13827 GND.n6663 GND.n6624 585
R13828 GND.n6624 GND.n6189 585
R13829 GND.n6665 GND.n6664 585
R13830 GND.n6665 GND.n6182 585
R13831 GND.n6666 GND.n6623 585
R13832 GND.n6666 GND.n6179 585
R13833 GND.n6668 GND.n6667 585
R13834 GND.n6667 GND.n6488 585
R13835 GND.n6669 GND.n6618 585
R13836 GND.n6618 GND.n6169 585
R13837 GND.n6671 GND.n6670 585
R13838 GND.n6671 GND.n6162 585
R13839 GND.n6672 GND.n6617 585
R13840 GND.n6672 GND.n6159 585
R13841 GND.n6674 GND.n6673 585
R13842 GND.n6673 GND.n6151 585
R13843 GND.n6675 GND.n6612 585
R13844 GND.n6612 GND.n6148 585
R13845 GND.n6677 GND.n6676 585
R13846 GND.n6677 GND.n6141 585
R13847 GND.n6678 GND.n6611 585
R13848 GND.n6678 GND.n6138 585
R13849 GND.n6680 GND.n6679 585
R13850 GND.n6679 GND.n6130 585
R13851 GND.n6681 GND.n6606 585
R13852 GND.n6606 GND.n6127 585
R13853 GND.n6683 GND.n6682 585
R13854 GND.n6683 GND.n6120 585
R13855 GND.n6684 GND.n6605 585
R13856 GND.n6684 GND.n6117 585
R13857 GND.n6686 GND.n6685 585
R13858 GND.n6685 GND.n6109 585
R13859 GND.n6687 GND.n6600 585
R13860 GND.n6600 GND.n6106 585
R13861 GND.n6689 GND.n6688 585
R13862 GND.n6689 GND.n6099 585
R13863 GND.n6690 GND.n6599 585
R13864 GND.n6690 GND.n6096 585
R13865 GND.n6692 GND.n6691 585
R13866 GND.n6691 GND.n6088 585
R13867 GND.n6693 GND.n6594 585
R13868 GND.n6594 GND.n6085 585
R13869 GND.n6695 GND.n6694 585
R13870 GND.n6695 GND.n6078 585
R13871 GND.n6696 GND.n6593 585
R13872 GND.n6696 GND.n6075 585
R13873 GND.n6698 GND.n6697 585
R13874 GND.n6697 GND.n6067 585
R13875 GND.n6699 GND.n6588 585
R13876 GND.n6588 GND.n6064 585
R13877 GND.n6701 GND.n6700 585
R13878 GND.n6701 GND.n6057 585
R13879 GND.n6702 GND.n6587 585
R13880 GND.n6702 GND.n6054 585
R13881 GND.n6704 GND.n6703 585
R13882 GND.n6703 GND.n6046 585
R13883 GND.n6705 GND.n6582 585
R13884 GND.n6582 GND.n6043 585
R13885 GND.n6707 GND.n6706 585
R13886 GND.n6707 GND.n6514 585
R13887 GND.n6708 GND.n6581 585
R13888 GND.n6708 GND.n6034 585
R13889 GND.n6710 GND.n6709 585
R13890 GND.n6709 GND.n6026 585
R13891 GND.n6711 GND.n6576 585
R13892 GND.n6576 GND.n6023 585
R13893 GND.n6713 GND.n6712 585
R13894 GND.n6713 GND.n6016 585
R13895 GND.n6714 GND.n6575 585
R13896 GND.n6714 GND.n6013 585
R13897 GND.n6716 GND.n6715 585
R13898 GND.n6715 GND.n6005 585
R13899 GND.n6717 GND.n6570 585
R13900 GND.n6570 GND.n6002 585
R13901 GND.n6719 GND.n6718 585
R13902 GND.n6719 GND.n5995 585
R13903 GND.n6720 GND.n6569 585
R13904 GND.n6720 GND.n5992 585
R13905 GND.n6722 GND.n6721 585
R13906 GND.n6721 GND.n5984 585
R13907 GND.n6723 GND.n6564 585
R13908 GND.n6564 GND.n5981 585
R13909 GND.n6725 GND.n6724 585
R13910 GND.n6725 GND.n5974 585
R13911 GND.n6726 GND.n6563 585
R13912 GND.n6726 GND.n5971 585
R13913 GND.n6728 GND.n6727 585
R13914 GND.n6727 GND.n5963 585
R13915 GND.n6729 GND.n6532 585
R13916 GND.n6532 GND.n5960 585
R13917 GND.n6731 GND.n6730 585
R13918 GND.n6732 GND.n6731 585
R13919 GND.n6533 GND.n6531 585
R13920 GND.n6531 GND.n5951 585
R13921 GND.n6557 GND.n6556 585
R13922 GND.n6556 GND.n5943 585
R13923 GND.n6555 GND.n6535 585
R13924 GND.n6555 GND.n5940 585
R13925 GND.n6554 GND.n6553 585
R13926 GND.n6554 GND.n5932 585
R13927 GND.n6537 GND.n6536 585
R13928 GND.n6536 GND.n5929 585
R13929 GND.n6549 GND.n6548 585
R13930 GND.n6548 GND.n5920 585
R13931 GND.n6547 GND.n6539 585
R13932 GND.n6547 GND.n5881 585
R13933 GND.n6546 GND.n6545 585
R13934 GND.n6546 GND.n5879 585
R13935 GND.n6541 GND.n6540 585
R13936 GND.n6540 GND.n4602 585
R13937 GND.n4567 GND.n4566 585
R13938 GND.n7648 GND.n4567 585
R13939 GND.n7651 GND.n7650 585
R13940 GND.n7650 GND.n7649 585
R13941 GND.n7652 GND.n4561 585
R13942 GND.n4561 GND.n4560 585
R13943 GND.n7654 GND.n7653 585
R13944 GND.n7655 GND.n7654 585
R13945 GND.n4526 GND.n4525 585
R13946 GND.n7656 GND.n4526 585
R13947 GND.n7660 GND.n7659 585
R13948 GND.n7659 GND.n7658 585
R13949 GND.n7661 GND.n4518 585
R13950 GND.n4650 GND.n4518 585
R13951 GND.n7663 GND.n7662 585
R13952 GND.n7664 GND.n7663 585
R13953 GND.n4519 GND.n4517 585
R13954 GND.n4517 GND.n4505 585
R13955 GND.n4448 GND.n4447 585
R13956 GND.n4504 GND.n4448 585
R13957 GND.n7679 GND.n7678 585
R13958 GND.n7678 GND.n7677 585
R13959 GND.n7680 GND.n4442 585
R13960 GND.n4497 GND.n4442 585
R13961 GND.n7682 GND.n7681 585
R13962 GND.n7683 GND.n7682 585
R13963 GND.n4431 GND.n4430 585
R13964 GND.n4434 GND.n4431 585
R13965 GND.n7693 GND.n7692 585
R13966 GND.n7692 GND.n7691 585
R13967 GND.n7694 GND.n4425 585
R13968 GND.n4486 GND.n4425 585
R13969 GND.n7696 GND.n7695 585
R13970 GND.n7697 GND.n7696 585
R13971 GND.n4413 GND.n4412 585
R13972 GND.n4416 GND.n4413 585
R13973 GND.n7707 GND.n7706 585
R13974 GND.n7706 GND.n7705 585
R13975 GND.n7708 GND.n4407 585
R13976 GND.n4473 GND.n4407 585
R13977 GND.n7710 GND.n7709 585
R13978 GND.n7711 GND.n7710 585
R13979 GND.n4395 GND.n4394 585
R13980 GND.n4398 GND.n4395 585
R13981 GND.n7721 GND.n7720 585
R13982 GND.n7720 GND.n7719 585
R13983 GND.n7722 GND.n4387 585
R13984 GND.n4460 GND.n4387 585
R13985 GND.n7724 GND.n7723 585
R13986 GND.n7725 GND.n7724 585
R13987 GND.n4388 GND.n4386 585
R13988 GND.n4386 GND.n4385 585
R13989 GND.n4364 GND.n4363 585
R13990 GND.n4375 GND.n4364 585
R13991 GND.n7740 GND.n7739 585
R13992 GND.n7739 GND.n7738 585
R13993 GND.n7741 GND.n4358 585
R13994 GND.n5809 GND.n4358 585
R13995 GND.n7743 GND.n7742 585
R13996 GND.n7744 GND.n7743 585
R13997 GND.n4345 GND.n4344 585
R13998 GND.n5793 GND.n4345 585
R13999 GND.n7752 GND.n7751 585
R14000 GND.n7751 GND.n7750 585
R14001 GND.n7753 GND.n4339 585
R14002 GND.n5801 GND.n4339 585
R14003 GND.n7755 GND.n7754 585
R14004 GND.n7756 GND.n7755 585
R14005 GND.n4325 GND.n4324 585
R14006 GND.n4872 GND.n4325 585
R14007 GND.n7764 GND.n7763 585
R14008 GND.n7763 GND.n7762 585
R14009 GND.n7765 GND.n4319 585
R14010 GND.n4877 GND.n4319 585
R14011 GND.n7767 GND.n7766 585
R14012 GND.n7768 GND.n7767 585
R14013 GND.n4292 GND.n4291 585
R14014 GND.n4882 GND.n4292 585
R14015 GND.n7776 GND.n7775 585
R14016 GND.n7775 GND.n7774 585
R14017 GND.n7777 GND.n4284 585
R14018 GND.n5743 GND.n4284 585
R14019 GND.n7779 GND.n7778 585
R14020 GND.n7780 GND.n7779 585
R14021 GND.n4285 GND.n4283 585
R14022 GND.n4283 GND.n4272 585
R14023 GND.n4260 GND.n4259 585
R14024 GND.n4271 GND.n4260 585
R14025 GND.n7795 GND.n7794 585
R14026 GND.n7794 GND.n7793 585
R14027 GND.n7796 GND.n4254 585
R14028 GND.n4888 GND.n4254 585
R14029 GND.n7798 GND.n7797 585
R14030 GND.n7799 GND.n7798 585
R14031 GND.n4242 GND.n4241 585
R14032 GND.n5710 GND.n4242 585
R14033 GND.n7807 GND.n7806 585
R14034 GND.n7806 GND.n7805 585
R14035 GND.n7808 GND.n4236 585
R14036 GND.n5631 GND.n4236 585
R14037 GND.n7810 GND.n7809 585
R14038 GND.n7811 GND.n7810 585
R14039 GND.n4222 GND.n4221 585
R14040 GND.n4905 GND.n4222 585
R14041 GND.n7819 GND.n7818 585
R14042 GND.n7818 GND.n7817 585
R14043 GND.n7820 GND.n4216 585
R14044 GND.n4910 GND.n4216 585
R14045 GND.n7822 GND.n7821 585
R14046 GND.n7823 GND.n7822 585
R14047 GND.n4190 GND.n4189 585
R14048 GND.n4915 GND.n4190 585
R14049 GND.n7831 GND.n7830 585
R14050 GND.n7830 GND.n7829 585
R14051 GND.n7832 GND.n4182 585
R14052 GND.n5646 GND.n4182 585
R14053 GND.n7834 GND.n7833 585
R14054 GND.n7835 GND.n7834 585
R14055 GND.n4183 GND.n4181 585
R14056 GND.n4181 GND.n4170 585
R14057 GND.n4158 GND.n4157 585
R14058 GND.n4169 GND.n4158 585
R14059 GND.n7850 GND.n7849 585
R14060 GND.n7849 GND.n7848 585
R14061 GND.n7851 GND.n4152 585
R14062 GND.n4922 GND.n4152 585
R14063 GND.n7853 GND.n7852 585
R14064 GND.n7854 GND.n7853 585
R14065 GND.n4138 GND.n4137 585
R14066 GND.n5607 GND.n4138 585
R14067 GND.n7862 GND.n7861 585
R14068 GND.n7861 GND.n7860 585
R14069 GND.n7863 GND.n4132 585
R14070 GND.n4932 GND.n4132 585
R14071 GND.n7865 GND.n7864 585
R14072 GND.n7866 GND.n7865 585
R14073 GND.n4118 GND.n4117 585
R14074 GND.n4937 GND.n4118 585
R14075 GND.n7874 GND.n7873 585
R14076 GND.n7873 GND.n7872 585
R14077 GND.n7875 GND.n4112 585
R14078 GND.n4942 GND.n4112 585
R14079 GND.n7877 GND.n7876 585
R14080 GND.n7878 GND.n7877 585
R14081 GND.n4085 GND.n4084 585
R14082 GND.n4947 GND.n4085 585
R14083 GND.n7886 GND.n7885 585
R14084 GND.n7885 GND.n7884 585
R14085 GND.n7887 GND.n4077 585
R14086 GND.n5542 GND.n4077 585
R14087 GND.n7889 GND.n7888 585
R14088 GND.n7890 GND.n7889 585
R14089 GND.n4078 GND.n4076 585
R14090 GND.n4076 GND.n4065 585
R14091 GND.n4053 GND.n4052 585
R14092 GND.n4064 GND.n4053 585
R14093 GND.n7905 GND.n7904 585
R14094 GND.n7904 GND.n7903 585
R14095 GND.n7906 GND.n4047 585
R14096 GND.n4953 GND.n4047 585
R14097 GND.n7908 GND.n7907 585
R14098 GND.n7909 GND.n7908 585
R14099 GND.n4033 GND.n4032 585
R14100 GND.n5504 GND.n4033 585
R14101 GND.n7917 GND.n7916 585
R14102 GND.n7916 GND.n7915 585
R14103 GND.n7918 GND.n4027 585
R14104 GND.n4963 GND.n4027 585
R14105 GND.n7920 GND.n7919 585
R14106 GND.n7921 GND.n7920 585
R14107 GND.n4013 GND.n4012 585
R14108 GND.n4968 GND.n4013 585
R14109 GND.n7929 GND.n7928 585
R14110 GND.n7928 GND.n7927 585
R14111 GND.n7930 GND.n4007 585
R14112 GND.n4973 GND.n4007 585
R14113 GND.n7932 GND.n7931 585
R14114 GND.n7933 GND.n7932 585
R14115 GND.n3993 GND.n3992 585
R14116 GND.n4978 GND.n3993 585
R14117 GND.n7941 GND.n7940 585
R14118 GND.n7940 GND.n7939 585
R14119 GND.n7942 GND.n3987 585
R14120 GND.n5397 GND.n3987 585
R14121 GND.n7944 GND.n7943 585
R14122 GND.n7945 GND.n7944 585
R14123 GND.n3973 GND.n3972 585
R14124 GND.n4987 GND.n3973 585
R14125 GND.n7953 GND.n7952 585
R14126 GND.n7952 GND.n7951 585
R14127 GND.n7954 GND.n3967 585
R14128 GND.n5430 GND.n3967 585
R14129 GND.n7956 GND.n7955 585
R14130 GND.n7957 GND.n7956 585
R14131 GND.n3953 GND.n3952 585
R14132 GND.n4997 GND.n3953 585
R14133 GND.n7965 GND.n7964 585
R14134 GND.n7964 GND.n7963 585
R14135 GND.n7966 GND.n3947 585
R14136 GND.n5411 GND.n3947 585
R14137 GND.n7968 GND.n7967 585
R14138 GND.n7969 GND.n7968 585
R14139 GND.n3933 GND.n3932 585
R14140 GND.n5362 GND.n3933 585
R14141 GND.n7977 GND.n7976 585
R14142 GND.n7976 GND.n7975 585
R14143 GND.n7978 GND.n3927 585
R14144 GND.n5351 GND.n3927 585
R14145 GND.n7980 GND.n7979 585
R14146 GND.n7981 GND.n7980 585
R14147 GND.n3913 GND.n3912 585
R14148 GND.n5343 GND.n3913 585
R14149 GND.n7989 GND.n7988 585
R14150 GND.n7988 GND.n7987 585
R14151 GND.n7990 GND.n3907 585
R14152 GND.n5332 GND.n3907 585
R14153 GND.n7992 GND.n7991 585
R14154 GND.n7993 GND.n7992 585
R14155 GND.n3892 GND.n3891 585
R14156 GND.n5324 GND.n3892 585
R14157 GND.n8001 GND.n8000 585
R14158 GND.n8000 GND.n7999 585
R14159 GND.n8002 GND.n3886 585
R14160 GND.n5024 GND.n3886 585
R14161 GND.n8004 GND.n8003 585
R14162 GND.n8005 GND.n8004 585
R14163 GND.n3849 GND.n3848 585
R14164 GND.n3881 GND.n3849 585
R14165 GND.n8059 GND.n8058 585
R14166 GND.n8058 GND.n8057 585
R14167 GND.n8060 GND.n3843 585
R14168 GND.n5035 GND.n3843 585
R14169 GND.n8062 GND.n8061 585
R14170 GND.n8063 GND.n8062 585
R14171 GND.n3831 GND.n3830 585
R14172 GND.n3834 GND.n3831 585
R14173 GND.n8073 GND.n8072 585
R14174 GND.n8072 GND.n8071 585
R14175 GND.n8074 GND.n3825 585
R14176 GND.n5250 GND.n3825 585
R14177 GND.n8076 GND.n8075 585
R14178 GND.n8077 GND.n8076 585
R14179 GND.n3813 GND.n3812 585
R14180 GND.n3816 GND.n3813 585
R14181 GND.n8087 GND.n8086 585
R14182 GND.n8086 GND.n8085 585
R14183 GND.n8088 GND.n3807 585
R14184 GND.n5237 GND.n3807 585
R14185 GND.n8090 GND.n8089 585
R14186 GND.n8091 GND.n8090 585
R14187 GND.n3795 GND.n3794 585
R14188 GND.n3798 GND.n3795 585
R14189 GND.n8101 GND.n8100 585
R14190 GND.n8100 GND.n8099 585
R14191 GND.n8102 GND.n3789 585
R14192 GND.n5224 GND.n3789 585
R14193 GND.n8104 GND.n8103 585
R14194 GND.n8105 GND.n8104 585
R14195 GND.n3779 GND.n3778 585
R14196 GND.t64 GND.n3779 585
R14197 GND.n8115 GND.n8114 585
R14198 GND.n8114 GND.n8113 585
R14199 GND.n8116 GND.n3773 585
R14200 GND.n5211 GND.n3773 585
R14201 GND.n8118 GND.n8117 585
R14202 GND.n8119 GND.n8118 585
R14203 GND.n3748 GND.n3747 585
R14204 GND.n3770 GND.n3748 585
R14205 GND.n8129 GND.n8128 585
R14206 GND.n8128 GND.n8127 585
R14207 GND.n8130 GND.n3740 585
R14208 GND.n3740 GND.n3739 585
R14209 GND.n8132 GND.n8131 585
R14210 GND.n8133 GND.n8132 585
R14211 GND.n3741 GND.n3738 585
R14212 GND.n8134 GND.n3738 585
R14213 GND.n8136 GND.n3737 585
R14214 GND.n8136 GND.n8135 585
R14215 GND.n8138 GND.n8137 585
R14216 GND.n8137 GND.n2166 585
R14217 GND.n8139 GND.n3732 585
R14218 GND.n3732 GND.n2147 585
R14219 GND.n8141 GND.n8140 585
R14220 GND.n8141 GND.n2128 585
R14221 GND.n8142 GND.n3731 585
R14222 GND.n8142 GND.n2125 585
R14223 GND.n8144 GND.n8143 585
R14224 GND.n8143 GND.n2214 585
R14225 GND.n8145 GND.n3726 585
R14226 GND.n3726 GND.n2221 585
R14227 GND.n8147 GND.n8146 585
R14228 GND.n8147 GND.n2220 585
R14229 GND.n8148 GND.n3725 585
R14230 GND.n8148 GND.n2234 585
R14231 GND.n8150 GND.n8149 585
R14232 GND.n8149 GND.n2231 585
R14233 GND.n8151 GND.n3720 585
R14234 GND.n3720 GND.n2237 585
R14235 GND.n8153 GND.n8152 585
R14236 GND.n8153 GND.n2244 585
R14237 GND.n8154 GND.n3719 585
R14238 GND.n8154 GND.n2243 585
R14239 GND.n8156 GND.n8155 585
R14240 GND.n8155 GND.n2255 585
R14241 GND.n8157 GND.n3714 585
R14242 GND.n3714 GND.n2253 585
R14243 GND.n8159 GND.n8158 585
R14244 GND.n8159 GND.n2258 585
R14245 GND.n8160 GND.n3713 585
R14246 GND.n8160 GND.n2266 585
R14247 GND.n8162 GND.n8161 585
R14248 GND.n8161 GND.n2264 585
R14249 GND.n8163 GND.n3708 585
R14250 GND.n3708 GND.n2277 585
R14251 GND.n8165 GND.n8164 585
R14252 GND.n8165 GND.n2275 585
R14253 GND.n8166 GND.n3707 585
R14254 GND.n8166 GND.n2279 585
R14255 GND.n8168 GND.n8167 585
R14256 GND.n8167 GND.n2286 585
R14257 GND.n8169 GND.n3702 585
R14258 GND.n3702 GND.n2285 585
R14259 GND.n8171 GND.n8170 585
R14260 GND.n8171 GND.n2298 585
R14261 GND.n8172 GND.n3701 585
R14262 GND.n8172 GND.n2296 585
R14263 GND.n8174 GND.n8173 585
R14264 GND.n8173 GND.n2300 585
R14265 GND.n8175 GND.n2323 585
R14266 GND.n2323 GND.n2307 585
R14267 GND.n8177 GND.n8176 585
R14268 GND.n8178 GND.n8177 585
R14269 GND.n2324 GND.n2322 585
R14270 GND.n2322 GND.n2320 585
R14271 GND.n3695 GND.n3694 585
R14272 GND.n3694 GND.n2317 585
R14273 GND.n3693 GND.n2326 585
R14274 GND.n3693 GND.n3692 585
R14275 GND.n2590 GND.n2327 585
R14276 GND.n2335 GND.n2327 585
R14277 GND.n2592 GND.n2591 585
R14278 GND.n2592 GND.n2334 585
R14279 GND.n2594 GND.n2593 585
R14280 GND.n2593 GND.n2347 585
R14281 GND.n2595 GND.n2583 585
R14282 GND.n2583 GND.n2345 585
R14283 GND.n2597 GND.n2596 585
R14284 GND.n2597 GND.n2350 585
R14285 GND.n2598 GND.n2582 585
R14286 GND.n2598 GND.n2358 585
R14287 GND.n2600 GND.n2599 585
R14288 GND.n2599 GND.n2356 585
R14289 GND.n2601 GND.n2577 585
R14290 GND.n2577 GND.n2369 585
R14291 GND.n2603 GND.n2602 585
R14292 GND.n2603 GND.n2367 585
R14293 GND.n2607 GND.n2576 585
R14294 GND.n2607 GND.n2606 585
R14295 GND.n2609 GND.n2608 585
R14296 GND.n2608 GND.n2377 585
R14297 GND.n2610 GND.n2571 585
R14298 GND.n2571 GND.n2376 585
R14299 GND.n2612 GND.n2611 585
R14300 GND.n2612 GND.n2387 585
R14301 GND.n2613 GND.n2570 585
R14302 GND.n2613 GND.n2385 585
R14303 GND.n2615 GND.n2614 585
R14304 GND.n2614 GND.n2389 585
R14305 GND.n2616 GND.n2565 585
R14306 GND.n2565 GND.n2397 585
R14307 GND.n2618 GND.n2617 585
R14308 GND.n2618 GND.n2396 585
R14309 GND.n2619 GND.n2564 585
R14310 GND.n2619 GND.n2410 585
R14311 GND.n2621 GND.n2620 585
R14312 GND.n2620 GND.n2407 585
R14313 GND.n2622 GND.n2559 585
R14314 GND.n2559 GND.n2413 585
R14315 GND.n2624 GND.n2623 585
R14316 GND.n2624 GND.n2420 585
R14317 GND.n2625 GND.n2558 585
R14318 GND.n2625 GND.n2419 585
R14319 GND.n2627 GND.n2626 585
R14320 GND.n2626 GND.n2431 585
R14321 GND.n2628 GND.n2553 585
R14322 GND.n2553 GND.n2429 585
R14323 GND.n2630 GND.n2629 585
R14324 GND.n2630 GND.n2434 585
R14325 GND.n2631 GND.n2552 585
R14326 GND.n2631 GND.n2442 585
R14327 GND.n2633 GND.n2632 585
R14328 GND.n2632 GND.n2440 585
R14329 GND.n2634 GND.n2547 585
R14330 GND.n2547 GND.n2453 585
R14331 GND.n2636 GND.n2635 585
R14332 GND.n2636 GND.n2451 585
R14333 GND.n2637 GND.n2546 585
R14334 GND.n2637 GND.n2455 585
R14335 GND.n2639 GND.n2638 585
R14336 GND.n2638 GND.n2462 585
R14337 GND.n2640 GND.n2541 585
R14338 GND.n2541 GND.n2461 585
R14339 GND.n2642 GND.n2641 585
R14340 GND.n2642 GND.n2474 585
R14341 GND.n2643 GND.n2540 585
R14342 GND.n2643 GND.n2472 585
R14343 GND.n2645 GND.n2644 585
R14344 GND.n2644 GND.n2476 585
R14345 GND.n2646 GND.n2537 585
R14346 GND.n2537 GND.n2484 585
R14347 GND.n2648 GND.n2647 585
R14348 GND.n2648 GND.n2483 585
R14349 GND.n3464 GND.n3463 585
R14350 GND.n3463 GND.n3462 585
R14351 GND.n3465 GND.n2533 585
R14352 GND.n2649 GND.n2533 585
R14353 GND.n3468 GND.n3467 585
R14354 GND.n3469 GND.n3468 585
R14355 GND.n2535 GND.n2532 585
R14356 GND.n2532 GND.n2527 585
R14357 GND.n2514 GND.n2513 585
R14358 GND.n2519 GND.n2514 585
R14359 GND.n3481 GND.n3480 585
R14360 GND.n3480 GND.n3479 585
R14361 GND.n3483 GND.n2511 585
R14362 GND.n2515 GND.n2511 585
R14363 GND.n3485 GND.n3484 585
R14364 GND.n3486 GND.n3485 585
R14365 GND.n2512 GND.n2510 585
R14366 GND.n2510 GND.n2504 585
R14367 GND.n3063 GND.n3062 585
R14368 GND.n3063 GND.n2501 585
R14369 GND.n3066 GND.n3060 585
R14370 GND.n3066 GND.n3065 585
R14371 GND.n3068 GND.n3067 585
R14372 GND.n3067 GND.n2661 585
R14373 GND.n3069 GND.n3054 585
R14374 GND.n3054 GND.n2672 585
R14375 GND.n3071 GND.n3070 585
R14376 GND.n3071 GND.n2669 585
R14377 GND.n3072 GND.n3053 585
R14378 GND.n3072 GND.n2675 585
R14379 GND.n3074 GND.n3073 585
R14380 GND.n3073 GND.n2683 585
R14381 GND.n3075 GND.n3048 585
R14382 GND.n3048 GND.n2682 585
R14383 GND.n3077 GND.n3076 585
R14384 GND.n3077 GND.n2694 585
R14385 GND.n3078 GND.n3047 585
R14386 GND.n3078 GND.n2692 585
R14387 GND.n3080 GND.n3079 585
R14388 GND.n3079 GND.n2697 585
R14389 GND.n3081 GND.n3042 585
R14390 GND.n3042 GND.n2706 585
R14391 GND.n3083 GND.n3082 585
R14392 GND.n3083 GND.n2704 585
R14393 GND.n3084 GND.n3041 585
R14394 GND.n3084 GND.n2717 585
R14395 GND.n3086 GND.n3085 585
R14396 GND.n3085 GND.n2715 585
R14397 GND.n3087 GND.n3036 585
R14398 GND.n3036 GND.n2719 585
R14399 GND.n3089 GND.n3088 585
R14400 GND.n3089 GND.n2727 585
R14401 GND.n3090 GND.n3035 585
R14402 GND.n3090 GND.n2726 585
R14403 GND.n3092 GND.n3091 585
R14404 GND.n3091 GND.n2739 585
R14405 GND.n3093 GND.n3030 585
R14406 GND.n3030 GND.n2737 585
R14407 GND.n3095 GND.n3094 585
R14408 GND.n3095 GND.n2741 585
R14409 GND.n3096 GND.n3029 585
R14410 GND.n3096 GND.n2750 585
R14411 GND.n3098 GND.n3097 585
R14412 GND.n3097 GND.n2749 585
R14413 GND.n3099 GND.n3024 585
R14414 GND.n3024 GND.n2763 585
R14415 GND.n3101 GND.n3100 585
R14416 GND.n3101 GND.n2760 585
R14417 GND.n3102 GND.n3023 585
R14418 GND.n3102 GND.n2766 585
R14419 GND.n3104 GND.n3103 585
R14420 GND.n3103 GND.n2774 585
R14421 GND.n3105 GND.n3018 585
R14422 GND.n3018 GND.n2773 585
R14423 GND.n3107 GND.n3106 585
R14424 GND.n3107 GND.n2785 585
R14425 GND.n3108 GND.n3017 585
R14426 GND.n3108 GND.n2783 585
R14427 GND.n3110 GND.n3109 585
R14428 GND.n3109 GND.n2788 585
R14429 GND.n3111 GND.n3012 585
R14430 GND.n3012 GND.n2797 585
R14431 GND.n3113 GND.n3112 585
R14432 GND.n3113 GND.n2795 585
R14433 GND.n3114 GND.n3011 585
R14434 GND.n3114 GND.n2808 585
R14435 GND.n3116 GND.n3115 585
R14436 GND.n3115 GND.n2806 585
R14437 GND.n3117 GND.n3006 585
R14438 GND.n3006 GND.n2810 585
R14439 GND.n3119 GND.n3118 585
R14440 GND.n3119 GND.n2818 585
R14441 GND.n3120 GND.n3005 585
R14442 GND.n3120 GND.n2817 585
R14443 GND.n3122 GND.n3121 585
R14444 GND.n3121 GND.n2830 585
R14445 GND.n3123 GND.n3000 585
R14446 GND.n3000 GND.n2828 585
R14447 GND.n3125 GND.n3124 585
R14448 GND.n3125 GND.n2832 585
R14449 GND.n3126 GND.n2999 585
R14450 GND.n3126 GND.n2841 585
R14451 GND.n3128 GND.n3127 585
R14452 GND.n3127 GND.n2840 585
R14453 GND.n3129 GND.n2994 585
R14454 GND.n2994 GND.n2854 585
R14455 GND.n3131 GND.n3130 585
R14456 GND.n3131 GND.n2851 585
R14457 GND.n3132 GND.n2993 585
R14458 GND.n3132 GND.n2857 585
R14459 GND.n3134 GND.n3133 585
R14460 GND.n3133 GND.n2865 585
R14461 GND.n3135 GND.n2988 585
R14462 GND.n2988 GND.n2864 585
R14463 GND.n3137 GND.n3136 585
R14464 GND.n3137 GND.n2876 585
R14465 GND.n3138 GND.n2987 585
R14466 GND.n3138 GND.n2874 585
R14467 GND.n3140 GND.n3139 585
R14468 GND.n3139 GND.n2879 585
R14469 GND.n3141 GND.n2982 585
R14470 GND.n2982 GND.n2888 585
R14471 GND.n3143 GND.n3142 585
R14472 GND.n3143 GND.n2886 585
R14473 GND.n3144 GND.n2981 585
R14474 GND.n3144 GND.n2899 585
R14475 GND.n3146 GND.n3145 585
R14476 GND.n3145 GND.n2897 585
R14477 GND.n3147 GND.n2968 585
R14478 GND.n2968 GND.n2901 585
R14479 GND.n3149 GND.n3148 585
R14480 GND.n3150 GND.n3149 585
R14481 GND.n2969 GND.n2967 585
R14482 GND.n2967 GND.n2965 585
R14483 GND.n2975 GND.n2974 585
R14484 GND.n2974 GND.n1839 585
R14485 GND.n2973 GND.n2972 585
R14486 GND.n2973 GND.n1836 585
R14487 GND.n1815 GND.n1814 585
R14488 GND.n1820 GND.n1815 585
R14489 GND.n8693 GND.n8692 585
R14490 GND.n8692 GND.n8691 585
R14491 GND.n8694 GND.n1807 585
R14492 GND.n1816 GND.n1807 585
R14493 GND.n8696 GND.n8695 585
R14494 GND.n8697 GND.n8696 585
R14495 GND.n1808 GND.n1806 585
R14496 GND.n1806 GND.n1801 585
R14497 GND.n1690 GND.n1689 585
R14498 GND.n1725 GND.n1690 585
R14499 GND.n8819 GND.n8818 585
R14500 GND.n8818 GND.n8817 585
R14501 GND.n8820 GND.n1684 585
R14502 GND.n1684 GND.n1683 585
R14503 GND.n8822 GND.n8821 585
R14504 GND.n8823 GND.n8822 585
R14505 GND.n1682 GND.n1681 585
R14506 GND.n8824 GND.n1682 585
R14507 GND.n8827 GND.n8826 585
R14508 GND.n8826 GND.n8825 585
R14509 GND.n8828 GND.n1676 585
R14510 GND.n1676 GND.n1675 585
R14511 GND.n8830 GND.n8829 585
R14512 GND.n8831 GND.n8830 585
R14513 GND.n1674 GND.n1673 585
R14514 GND.n8832 GND.n1674 585
R14515 GND.n8835 GND.n8834 585
R14516 GND.n8834 GND.n8833 585
R14517 GND.n8836 GND.n1668 585
R14518 GND.n1668 GND.n1667 585
R14519 GND.n8838 GND.n8837 585
R14520 GND.n8839 GND.n8838 585
R14521 GND.n1666 GND.n1665 585
R14522 GND.n8840 GND.n1666 585
R14523 GND.n8843 GND.n8842 585
R14524 GND.n8842 GND.n8841 585
R14525 GND.n8844 GND.n1660 585
R14526 GND.n1660 GND.n1659 585
R14527 GND.n8846 GND.n8845 585
R14528 GND.n8847 GND.n8846 585
R14529 GND.n1658 GND.n1657 585
R14530 GND.n8848 GND.n1658 585
R14531 GND.n8851 GND.n8850 585
R14532 GND.n8850 GND.n8849 585
R14533 GND.n8852 GND.n1652 585
R14534 GND.n1652 GND.n1651 585
R14535 GND.n8854 GND.n8853 585
R14536 GND.n8855 GND.n8854 585
R14537 GND.n1650 GND.n1649 585
R14538 GND.n8856 GND.n1650 585
R14539 GND.n8859 GND.n8858 585
R14540 GND.n8858 GND.n8857 585
R14541 GND.n8860 GND.n1644 585
R14542 GND.n1644 GND.n1643 585
R14543 GND.n8862 GND.n8861 585
R14544 GND.n8863 GND.n8862 585
R14545 GND.n1642 GND.n1641 585
R14546 GND.n8864 GND.n1642 585
R14547 GND.n8867 GND.n8866 585
R14548 GND.n8866 GND.n8865 585
R14549 GND.n8868 GND.n1636 585
R14550 GND.n1636 GND.n1635 585
R14551 GND.n8870 GND.n8869 585
R14552 GND.n8871 GND.n8870 585
R14553 GND.n1634 GND.n1633 585
R14554 GND.n8872 GND.n1634 585
R14555 GND.n8875 GND.n8874 585
R14556 GND.n8874 GND.n8873 585
R14557 GND.n8876 GND.n1628 585
R14558 GND.n1628 GND.n1627 585
R14559 GND.n8878 GND.n8877 585
R14560 GND.n8879 GND.n8878 585
R14561 GND.n1626 GND.n1625 585
R14562 GND.n8880 GND.n1626 585
R14563 GND.n8883 GND.n8882 585
R14564 GND.n8882 GND.n8881 585
R14565 GND.n8884 GND.n1620 585
R14566 GND.n1620 GND.n1619 585
R14567 GND.n8886 GND.n8885 585
R14568 GND.n8887 GND.n8886 585
R14569 GND.n1618 GND.n1617 585
R14570 GND.n8888 GND.n1618 585
R14571 GND.n8891 GND.n8890 585
R14572 GND.n8890 GND.n8889 585
R14573 GND.n8892 GND.n1612 585
R14574 GND.n1612 GND.n1611 585
R14575 GND.n8894 GND.n8893 585
R14576 GND.n8895 GND.n8894 585
R14577 GND.n1610 GND.n1609 585
R14578 GND.n8896 GND.n1610 585
R14579 GND.n8899 GND.n8898 585
R14580 GND.n8898 GND.n8897 585
R14581 GND.n8900 GND.n1604 585
R14582 GND.n1604 GND.n1603 585
R14583 GND.n8902 GND.n8901 585
R14584 GND.n8903 GND.n8902 585
R14585 GND.n1602 GND.n1601 585
R14586 GND.n8904 GND.n1602 585
R14587 GND.n8907 GND.n8906 585
R14588 GND.n8906 GND.n8905 585
R14589 GND.n8908 GND.n1596 585
R14590 GND.n1596 GND.n1595 585
R14591 GND.n8910 GND.n8909 585
R14592 GND.n8911 GND.n8910 585
R14593 GND.n1594 GND.n1593 585
R14594 GND.n8912 GND.n1594 585
R14595 GND.n8915 GND.n8914 585
R14596 GND.n8914 GND.n8913 585
R14597 GND.n8916 GND.n1589 585
R14598 GND.n1589 GND.n1588 585
R14599 GND.n8918 GND.n8917 585
R14600 GND.n8919 GND.n8918 585
R14601 GND.n1586 GND.n1584 585
R14602 GND.n8920 GND.n1586 585
R14603 GND.n8923 GND.n8922 585
R14604 GND.n8922 GND.n8921 585
R14605 GND.n1585 GND.n1582 585
R14606 GND.n1587 GND.n1585 585
R14607 GND.n8927 GND.n1579 585
R14608 GND.n1579 GND.n1578 585
R14609 GND.n8929 GND.n8928 585
R14610 GND.n8930 GND.n8929 585
R14611 GND.n8479 GND.n2121 585
R14612 GND.n8480 GND.n8479 585
R14613 GND.n2129 GND.n2120 585
R14614 GND.n8304 GND.n2129 585
R14615 GND.n2223 GND.n2119 585
R14616 GND.n2223 GND.n2222 585
R14617 GND.n2225 GND.n2224 585
R14618 GND.n8294 GND.n2225 585
R14619 GND.n8283 GND.n2113 585
R14620 GND.n8283 GND.n8282 585
R14621 GND.n8284 GND.n2112 585
R14622 GND.n8285 GND.n8284 585
R14623 GND.n8281 GND.n2111 585
R14624 GND.n8281 GND.n8280 585
R14625 GND.n2236 GND.n2235 585
R14626 GND.n2247 GND.n2236 585
R14627 GND.n2245 GND.n2105 585
R14628 GND.n8270 GND.n2245 585
R14629 GND.n8258 GND.n2104 585
R14630 GND.n8258 GND.n8257 585
R14631 GND.n8259 GND.n2103 585
R14632 GND.n8260 GND.n8259 585
R14633 GND.n8255 GND.n2257 585
R14634 GND.n8255 GND.n8254 585
R14635 GND.n2256 GND.n2097 585
R14636 GND.n2269 GND.n2256 585
R14637 GND.n2267 GND.n2096 585
R14638 GND.n8244 GND.n2267 585
R14639 GND.n8231 GND.n2095 585
R14640 GND.n8231 GND.n8230 585
R14641 GND.n8233 GND.n8232 585
R14642 GND.n8234 GND.n8233 585
R14643 GND.n8229 GND.n2089 585
R14644 GND.n8229 GND.n8228 585
R14645 GND.n2278 GND.n2088 585
R14646 GND.n2290 GND.n2278 585
R14647 GND.n2287 GND.n2087 585
R14648 GND.n8218 GND.n2287 585
R14649 GND.n8206 GND.n8204 585
R14650 GND.n8206 GND.n8205 585
R14651 GND.n8207 GND.n2081 585
R14652 GND.n8208 GND.n8207 585
R14653 GND.n8203 GND.n2080 585
R14654 GND.n8203 GND.n8202 585
R14655 GND.n2299 GND.n2079 585
R14656 GND.n2311 GND.n2299 585
R14657 GND.n2309 GND.n2308 585
R14658 GND.n8192 GND.n2309 585
R14659 GND.n8180 GND.n2073 585
R14660 GND.n8180 GND.n8179 585
R14661 GND.n8181 GND.n2072 585
R14662 GND.n8182 GND.n8181 585
R14663 GND.n2321 GND.n2071 585
R14664 GND.n3691 GND.n2321 585
R14665 GND.n2337 GND.n2336 585
R14666 GND.n2337 GND.n2328 585
R14667 GND.n2338 GND.n2065 585
R14668 GND.n3681 GND.n2338 585
R14669 GND.n3669 GND.n2064 585
R14670 GND.n3669 GND.n3668 585
R14671 GND.n3670 GND.n2063 585
R14672 GND.n3671 GND.n3670 585
R14673 GND.n3666 GND.n2349 585
R14674 GND.n3666 GND.n3665 585
R14675 GND.n2348 GND.n2057 585
R14676 GND.n2361 GND.n2348 585
R14677 GND.n2359 GND.n2056 585
R14678 GND.n3655 GND.n2359 585
R14679 GND.n3642 GND.n2055 585
R14680 GND.n3642 GND.n3641 585
R14681 GND.n3644 GND.n3643 585
R14682 GND.n3645 GND.n3644 585
R14683 GND.n3640 GND.n2049 585
R14684 GND.n3640 GND.n3639 585
R14685 GND.n2370 GND.n2048 585
R14686 GND.n2605 GND.n2370 585
R14687 GND.n2378 GND.n2047 585
R14688 GND.n3629 GND.n2378 585
R14689 GND.n3617 GND.n3615 585
R14690 GND.n3617 GND.n3616 585
R14691 GND.n3618 GND.n2041 585
R14692 GND.n3619 GND.n3618 585
R14693 GND.n3614 GND.n2040 585
R14694 GND.n3614 GND.n3613 585
R14695 GND.n2388 GND.n2039 585
R14696 GND.n2401 GND.n2388 585
R14697 GND.n2399 GND.n2398 585
R14698 GND.n3603 GND.n2399 585
R14699 GND.n3591 GND.n2033 585
R14700 GND.n3591 GND.n3590 585
R14701 GND.n3592 GND.n2032 585
R14702 GND.n3593 GND.n3592 585
R14703 GND.n3589 GND.n2031 585
R14704 GND.n3589 GND.n3588 585
R14705 GND.n2412 GND.n2411 585
R14706 GND.n2423 GND.n2412 585
R14707 GND.n2421 GND.n2025 585
R14708 GND.n3578 GND.n2421 585
R14709 GND.n3566 GND.n2024 585
R14710 GND.n3566 GND.n3565 585
R14711 GND.n3567 GND.n2023 585
R14712 GND.n3568 GND.n3567 585
R14713 GND.n3563 GND.n2433 585
R14714 GND.n3563 GND.n3562 585
R14715 GND.n2432 GND.n2017 585
R14716 GND.n2445 GND.n2432 585
R14717 GND.n2443 GND.n2016 585
R14718 GND.n3552 GND.n2443 585
R14719 GND.n3539 GND.n2015 585
R14720 GND.n3539 GND.n3538 585
R14721 GND.n3541 GND.n3540 585
R14722 GND.n3542 GND.n3541 585
R14723 GND.n3537 GND.n2009 585
R14724 GND.n3537 GND.n3536 585
R14725 GND.n2454 GND.n2008 585
R14726 GND.n2466 GND.n2454 585
R14727 GND.n2463 GND.n2007 585
R14728 GND.n3526 GND.n2463 585
R14729 GND.n3514 GND.n3512 585
R14730 GND.n3514 GND.n3513 585
R14731 GND.n3515 GND.n2001 585
R14732 GND.n3516 GND.n3515 585
R14733 GND.n3511 GND.n2000 585
R14734 GND.n3511 GND.n3510 585
R14735 GND.n2475 GND.n1999 585
R14736 GND.n2488 GND.n2475 585
R14737 GND.n2486 GND.n2485 585
R14738 GND.n3500 GND.n2486 585
R14739 GND.n3460 GND.n1993 585
R14740 GND.n3461 GND.n3460 585
R14741 GND.n3459 GND.n1992 585
R14742 GND.n3459 GND.n3458 585
R14743 GND.n2528 GND.n1991 585
R14744 GND.n2531 GND.n2528 585
R14745 GND.n3471 GND.n2529 585
R14746 GND.n3471 GND.n3470 585
R14747 GND.n3472 GND.n1985 585
R14748 GND.n3473 GND.n3472 585
R14749 GND.n2521 GND.n1984 585
R14750 GND.n3478 GND.n2521 585
R14751 GND.n2520 GND.n1983 585
R14752 GND.n2520 GND.n2516 585
R14753 GND.n2507 GND.n2506 585
R14754 GND.n2509 GND.n2507 585
R14755 GND.n3488 GND.n1977 585
R14756 GND.n3488 GND.n3487 585
R14757 GND.n3489 GND.n1976 585
R14758 GND.n3490 GND.n3489 585
R14759 GND.n2505 GND.n1975 585
R14760 GND.n3064 GND.n2505 585
R14761 GND.n2663 GND.n2662 585
R14762 GND.n3430 GND.n2663 585
R14763 GND.n3420 GND.n1969 585
R14764 GND.n3420 GND.n3419 585
R14765 GND.n3421 GND.n1968 585
R14766 GND.n3422 GND.n3421 585
R14767 GND.n3418 GND.n1967 585
R14768 GND.n3418 GND.n3417 585
R14769 GND.n2674 GND.n2673 585
R14770 GND.n2686 GND.n2674 585
R14771 GND.n2684 GND.n1961 585
R14772 GND.n3408 GND.n2684 585
R14773 GND.n3396 GND.n1960 585
R14774 GND.n3396 GND.n3395 585
R14775 GND.n3397 GND.n1959 585
R14776 GND.n3398 GND.n3397 585
R14777 GND.n3393 GND.n2696 585
R14778 GND.n3393 GND.n3392 585
R14779 GND.n2695 GND.n1953 585
R14780 GND.n2709 GND.n2695 585
R14781 GND.n2707 GND.n1952 585
R14782 GND.n3383 GND.n2707 585
R14783 GND.n3370 GND.n1951 585
R14784 GND.n3370 GND.n3369 585
R14785 GND.n3372 GND.n3371 585
R14786 GND.n3373 GND.n3372 585
R14787 GND.n3368 GND.n1945 585
R14788 GND.n3368 GND.n3367 585
R14789 GND.n2718 GND.n1944 585
R14790 GND.n2731 GND.n2718 585
R14791 GND.n2728 GND.n1943 585
R14792 GND.n3358 GND.n2728 585
R14793 GND.n3346 GND.n3344 585
R14794 GND.n3346 GND.n3345 585
R14795 GND.n3347 GND.n1937 585
R14796 GND.n3348 GND.n3347 585
R14797 GND.n3343 GND.n1936 585
R14798 GND.n3343 GND.n3342 585
R14799 GND.n2740 GND.n1935 585
R14800 GND.n2754 GND.n2740 585
R14801 GND.n2752 GND.n2751 585
R14802 GND.n3333 GND.n2752 585
R14803 GND.n3321 GND.n1929 585
R14804 GND.n3321 GND.n3320 585
R14805 GND.n3322 GND.n1928 585
R14806 GND.n3323 GND.n3322 585
R14807 GND.n3319 GND.n1927 585
R14808 GND.n3319 GND.n3318 585
R14809 GND.n2765 GND.n2764 585
R14810 GND.n2777 GND.n2765 585
R14811 GND.n2775 GND.n1921 585
R14812 GND.n3309 GND.n2775 585
R14813 GND.n3297 GND.n1920 585
R14814 GND.n3297 GND.n3296 585
R14815 GND.n3298 GND.n1919 585
R14816 GND.n3299 GND.n3298 585
R14817 GND.n3294 GND.n2787 585
R14818 GND.n3294 GND.n3293 585
R14819 GND.n2786 GND.n1913 585
R14820 GND.n2800 GND.n2786 585
R14821 GND.n2798 GND.n1912 585
R14822 GND.n3284 GND.n2798 585
R14823 GND.n3271 GND.n1911 585
R14824 GND.n3271 GND.n3270 585
R14825 GND.n3273 GND.n3272 585
R14826 GND.n3274 GND.n3273 585
R14827 GND.n3269 GND.n1905 585
R14828 GND.n3269 GND.n3268 585
R14829 GND.n2809 GND.n1904 585
R14830 GND.n2822 GND.n2809 585
R14831 GND.n2819 GND.n1903 585
R14832 GND.n3259 GND.n2819 585
R14833 GND.n3247 GND.n3245 585
R14834 GND.n3247 GND.n3246 585
R14835 GND.n3248 GND.n1897 585
R14836 GND.n3249 GND.n3248 585
R14837 GND.n3244 GND.n1896 585
R14838 GND.n3244 GND.n3243 585
R14839 GND.n2831 GND.n1895 585
R14840 GND.n2845 GND.n2831 585
R14841 GND.n2843 GND.n2842 585
R14842 GND.n3234 GND.n2843 585
R14843 GND.n3222 GND.n1889 585
R14844 GND.n3222 GND.n3221 585
R14845 GND.n3223 GND.n1888 585
R14846 GND.n3224 GND.n3223 585
R14847 GND.n3220 GND.n1887 585
R14848 GND.n3220 GND.n3219 585
R14849 GND.n2856 GND.n2855 585
R14850 GND.n2868 GND.n2856 585
R14851 GND.n2866 GND.n1881 585
R14852 GND.n3210 GND.n2866 585
R14853 GND.n3198 GND.n1880 585
R14854 GND.n3198 GND.n3197 585
R14855 GND.n3199 GND.n1879 585
R14856 GND.n3200 GND.n3199 585
R14857 GND.n3195 GND.n2878 585
R14858 GND.n3195 GND.n3194 585
R14859 GND.n2877 GND.n1873 585
R14860 GND.n2891 GND.n2877 585
R14861 GND.n2889 GND.n1872 585
R14862 GND.n3185 GND.n2889 585
R14863 GND.n3172 GND.n1871 585
R14864 GND.n3172 GND.n3171 585
R14865 GND.n3174 GND.n3173 585
R14866 GND.n3175 GND.n3174 585
R14867 GND.n3170 GND.n1865 585
R14868 GND.n3170 GND.n3169 585
R14869 GND.n2900 GND.n1864 585
R14870 GND.n3152 GND.n2900 585
R14871 GND.n2966 GND.n1863 585
R14872 GND.n3160 GND.n2966 585
R14873 GND.n1843 GND.n1841 585
R14874 GND.n2964 GND.n1841 585
R14875 GND.n8683 GND.n8682 585
R14876 GND.n8684 GND.n8683 585
R14877 GND.n1842 GND.n1840 585
R14878 GND.n2907 GND.n1840 585
R14879 GND.n1856 GND.n1821 585
R14880 GND.n8690 GND.n1821 585
R14881 GND.n1855 GND.n1854 585
R14882 GND.n1854 GND.n1817 585
R14883 GND.n1853 GND.n1799 585
R14884 GND.n1805 GND.n1799 585
R14885 GND.n8699 GND.n1800 585
R14886 GND.n8699 GND.n8698 585
R14887 GND.n8701 GND.n8700 585
R14888 GND.n2921 GND.n1798 585
R14889 GND.n2923 GND.n2922 585
R14890 GND.n2927 GND.n2926 585
R14891 GND.n2929 GND.n2928 585
R14892 GND.n2932 GND.n2931 585
R14893 GND.n2930 GND.n2919 585
R14894 GND.n2937 GND.n2936 585
R14895 GND.n2939 GND.n2938 585
R14896 GND.n2942 GND.n2941 585
R14897 GND.n2940 GND.n2916 585
R14898 GND.n2946 GND.n2917 585
R14899 GND.n2947 GND.n2913 585
R14900 GND.n2949 GND.n2948 585
R14901 GND.n8301 GND.n2127 585
R14902 GND.n8480 GND.n2127 585
R14903 GND.n8303 GND.n8302 585
R14904 GND.n8304 GND.n8303 585
R14905 GND.n2216 GND.n2215 585
R14906 GND.n2222 GND.n2215 585
R14907 GND.n8296 GND.n8295 585
R14908 GND.n8295 GND.n8294 585
R14909 GND.n2219 GND.n2218 585
R14910 GND.n8282 GND.n2219 585
R14911 GND.n8277 GND.n2233 585
R14912 GND.n8285 GND.n2233 585
R14913 GND.n8279 GND.n8278 585
R14914 GND.n8280 GND.n8279 585
R14915 GND.n2239 GND.n2238 585
R14916 GND.n2247 GND.n2238 585
R14917 GND.n8272 GND.n8271 585
R14918 GND.n8271 GND.n8270 585
R14919 GND.n2242 GND.n2241 585
R14920 GND.n8257 GND.n2242 585
R14921 GND.n8251 GND.n2254 585
R14922 GND.n8260 GND.n2254 585
R14923 GND.n8253 GND.n8252 585
R14924 GND.n8254 GND.n8253 585
R14925 GND.n2260 GND.n2259 585
R14926 GND.n2269 GND.n2259 585
R14927 GND.n8246 GND.n8245 585
R14928 GND.n8245 GND.n8244 585
R14929 GND.n2263 GND.n2262 585
R14930 GND.n8230 GND.n2263 585
R14931 GND.n8225 GND.n2276 585
R14932 GND.n8234 GND.n2276 585
R14933 GND.n8227 GND.n8226 585
R14934 GND.n8228 GND.n8227 585
R14935 GND.n2281 GND.n2280 585
R14936 GND.n2290 GND.n2280 585
R14937 GND.n8220 GND.n8219 585
R14938 GND.n8219 GND.n8218 585
R14939 GND.n2284 GND.n2283 585
R14940 GND.n8205 GND.n2284 585
R14941 GND.n8199 GND.n2297 585
R14942 GND.n8208 GND.n2297 585
R14943 GND.n8201 GND.n8200 585
R14944 GND.n8202 GND.n8201 585
R14945 GND.n2303 GND.n2302 585
R14946 GND.n2311 GND.n2302 585
R14947 GND.n8194 GND.n8193 585
R14948 GND.n8193 GND.n8192 585
R14949 GND.n2306 GND.n2305 585
R14950 GND.n8179 GND.n2306 585
R14951 GND.n3688 GND.n2319 585
R14952 GND.n8182 GND.n2319 585
R14953 GND.n3690 GND.n3689 585
R14954 GND.n3691 GND.n3690 585
R14955 GND.n2330 GND.n2329 585
R14956 GND.n2329 GND.n2328 585
R14957 GND.n3683 GND.n3682 585
R14958 GND.n3682 GND.n3681 585
R14959 GND.n2333 GND.n2332 585
R14960 GND.n3668 GND.n2333 585
R14961 GND.n3662 GND.n2346 585
R14962 GND.n3671 GND.n2346 585
R14963 GND.n3664 GND.n3663 585
R14964 GND.n3665 GND.n3664 585
R14965 GND.n2352 GND.n2351 585
R14966 GND.n2361 GND.n2351 585
R14967 GND.n3657 GND.n3656 585
R14968 GND.n3656 GND.n3655 585
R14969 GND.n2355 GND.n2354 585
R14970 GND.n3641 GND.n2355 585
R14971 GND.n3636 GND.n2368 585
R14972 GND.n3645 GND.n2368 585
R14973 GND.n3638 GND.n3637 585
R14974 GND.n3639 GND.n3638 585
R14975 GND.n2372 GND.n2371 585
R14976 GND.n2605 GND.n2371 585
R14977 GND.n3631 GND.n3630 585
R14978 GND.n3630 GND.n3629 585
R14979 GND.n2375 GND.n2374 585
R14980 GND.n3616 GND.n2375 585
R14981 GND.n3610 GND.n2386 585
R14982 GND.n3619 GND.n2386 585
R14983 GND.n3612 GND.n3611 585
R14984 GND.n3613 GND.n3612 585
R14985 GND.n2392 GND.n2391 585
R14986 GND.n2401 GND.n2391 585
R14987 GND.n3605 GND.n3604 585
R14988 GND.n3604 GND.n3603 585
R14989 GND.n2395 GND.n2394 585
R14990 GND.n3590 GND.n2395 585
R14991 GND.n3585 GND.n2409 585
R14992 GND.n3593 GND.n2409 585
R14993 GND.n3587 GND.n3586 585
R14994 GND.n3588 GND.n3587 585
R14995 GND.n2415 GND.n2414 585
R14996 GND.n2423 GND.n2414 585
R14997 GND.n3580 GND.n3579 585
R14998 GND.n3579 GND.n3578 585
R14999 GND.n2418 GND.n2417 585
R15000 GND.n3565 GND.n2418 585
R15001 GND.n3559 GND.n2430 585
R15002 GND.n3568 GND.n2430 585
R15003 GND.n3561 GND.n3560 585
R15004 GND.n3562 GND.n3561 585
R15005 GND.n2436 GND.n2435 585
R15006 GND.n2445 GND.n2435 585
R15007 GND.n3554 GND.n3553 585
R15008 GND.n3553 GND.n3552 585
R15009 GND.n2439 GND.n2438 585
R15010 GND.n3538 GND.n2439 585
R15011 GND.n3533 GND.n2452 585
R15012 GND.n3542 GND.n2452 585
R15013 GND.n3535 GND.n3534 585
R15014 GND.n3536 GND.n3535 585
R15015 GND.n2457 GND.n2456 585
R15016 GND.n2466 GND.n2456 585
R15017 GND.n3528 GND.n3527 585
R15018 GND.n3527 GND.n3526 585
R15019 GND.n2460 GND.n2459 585
R15020 GND.n3513 GND.n2460 585
R15021 GND.n3507 GND.n2473 585
R15022 GND.n3516 GND.n2473 585
R15023 GND.n3509 GND.n3508 585
R15024 GND.n3510 GND.n3509 585
R15025 GND.n2479 GND.n2478 585
R15026 GND.n2488 GND.n2478 585
R15027 GND.n3502 GND.n3501 585
R15028 GND.n3501 GND.n3500 585
R15029 GND.n2482 GND.n2481 585
R15030 GND.n3461 GND.n2482 585
R15031 GND.n3452 GND.n3451 585
R15032 GND.n3458 GND.n3452 585
R15033 GND.n2652 GND.n2651 585
R15034 GND.n2651 GND.n2531 585
R15035 GND.n3447 GND.n2530 585
R15036 GND.n3470 GND.n2530 585
R15037 GND.n3446 GND.n2526 585
R15038 GND.n3473 GND.n2526 585
R15039 GND.n3445 GND.n2518 585
R15040 GND.n3478 GND.n2518 585
R15041 GND.n3438 GND.n2654 585
R15042 GND.n3438 GND.n2516 585
R15043 GND.n3440 GND.n3439 585
R15044 GND.n3439 GND.n2509 585
R15045 GND.n3437 GND.n2508 585
R15046 GND.n3487 GND.n2508 585
R15047 GND.n3436 GND.n2503 585
R15048 GND.n3490 GND.n2503 585
R15049 GND.n2660 GND.n2656 585
R15050 GND.n3064 GND.n2660 585
R15051 GND.n3432 GND.n3431 585
R15052 GND.n3431 GND.n3430 585
R15053 GND.n2659 GND.n2658 585
R15054 GND.n3419 GND.n2659 585
R15055 GND.n2678 GND.n2671 585
R15056 GND.n3422 GND.n2671 585
R15057 GND.n3416 GND.n3415 585
R15058 GND.n3417 GND.n3416 585
R15059 GND.n2677 GND.n2676 585
R15060 GND.n2686 GND.n2676 585
R15061 GND.n3410 GND.n3409 585
R15062 GND.n3409 GND.n3408 585
R15063 GND.n2681 GND.n2680 585
R15064 GND.n3395 GND.n2681 585
R15065 GND.n2700 GND.n2693 585
R15066 GND.n3398 GND.n2693 585
R15067 GND.n3391 GND.n3390 585
R15068 GND.n3392 GND.n3391 585
R15069 GND.n2699 GND.n2698 585
R15070 GND.n2709 GND.n2698 585
R15071 GND.n3385 GND.n3384 585
R15072 GND.n3384 GND.n3383 585
R15073 GND.n2703 GND.n2702 585
R15074 GND.n3369 GND.n2703 585
R15075 GND.n2722 GND.n2716 585
R15076 GND.n3373 GND.n2716 585
R15077 GND.n3366 GND.n3365 585
R15078 GND.n3367 GND.n3366 585
R15079 GND.n2721 GND.n2720 585
R15080 GND.n2731 GND.n2720 585
R15081 GND.n3360 GND.n3359 585
R15082 GND.n3359 GND.n3358 585
R15083 GND.n2725 GND.n2724 585
R15084 GND.n3345 GND.n2725 585
R15085 GND.n2745 GND.n2738 585
R15086 GND.n3348 GND.n2738 585
R15087 GND.n3341 GND.n3340 585
R15088 GND.n3342 GND.n3341 585
R15089 GND.n2744 GND.n2743 585
R15090 GND.n2754 GND.n2743 585
R15091 GND.n3335 GND.n3334 585
R15092 GND.n3334 GND.n3333 585
R15093 GND.n2748 GND.n2747 585
R15094 GND.n3320 GND.n2748 585
R15095 GND.n2769 GND.n2762 585
R15096 GND.n3323 GND.n2762 585
R15097 GND.n3317 GND.n3316 585
R15098 GND.n3318 GND.n3317 585
R15099 GND.n2768 GND.n2767 585
R15100 GND.n2777 GND.n2767 585
R15101 GND.n3311 GND.n3310 585
R15102 GND.n3310 GND.n3309 585
R15103 GND.n2772 GND.n2771 585
R15104 GND.n3296 GND.n2772 585
R15105 GND.n2791 GND.n2784 585
R15106 GND.n3299 GND.n2784 585
R15107 GND.n3292 GND.n3291 585
R15108 GND.n3293 GND.n3292 585
R15109 GND.n2790 GND.n2789 585
R15110 GND.n2800 GND.n2789 585
R15111 GND.n3286 GND.n3285 585
R15112 GND.n3285 GND.n3284 585
R15113 GND.n2794 GND.n2793 585
R15114 GND.n3270 GND.n2794 585
R15115 GND.n2813 GND.n2807 585
R15116 GND.n3274 GND.n2807 585
R15117 GND.n3267 GND.n3266 585
R15118 GND.n3268 GND.n3267 585
R15119 GND.n2812 GND.n2811 585
R15120 GND.n2822 GND.n2811 585
R15121 GND.n3261 GND.n3260 585
R15122 GND.n3260 GND.n3259 585
R15123 GND.n2816 GND.n2815 585
R15124 GND.n3246 GND.n2816 585
R15125 GND.n2836 GND.n2829 585
R15126 GND.n3249 GND.n2829 585
R15127 GND.n3242 GND.n3241 585
R15128 GND.n3243 GND.n3242 585
R15129 GND.n2835 GND.n2834 585
R15130 GND.n2845 GND.n2834 585
R15131 GND.n3236 GND.n3235 585
R15132 GND.n3235 GND.n3234 585
R15133 GND.n2839 GND.n2838 585
R15134 GND.n3221 GND.n2839 585
R15135 GND.n2860 GND.n2853 585
R15136 GND.n3224 GND.n2853 585
R15137 GND.n3218 GND.n3217 585
R15138 GND.n3219 GND.n3218 585
R15139 GND.n2859 GND.n2858 585
R15140 GND.n2868 GND.n2858 585
R15141 GND.n3212 GND.n3211 585
R15142 GND.n3211 GND.n3210 585
R15143 GND.n2863 GND.n2862 585
R15144 GND.n3197 GND.n2863 585
R15145 GND.n2882 GND.n2875 585
R15146 GND.n3200 GND.n2875 585
R15147 GND.n3193 GND.n3192 585
R15148 GND.n3194 GND.n3193 585
R15149 GND.n2881 GND.n2880 585
R15150 GND.n2891 GND.n2880 585
R15151 GND.n3187 GND.n3186 585
R15152 GND.n3186 GND.n3185 585
R15153 GND.n2885 GND.n2884 585
R15154 GND.n3171 GND.n2885 585
R15155 GND.n2904 GND.n2898 585
R15156 GND.n3175 GND.n2898 585
R15157 GND.n3168 GND.n3167 585
R15158 GND.n3169 GND.n3168 585
R15159 GND.n2903 GND.n2902 585
R15160 GND.n3152 GND.n2902 585
R15161 GND.n3162 GND.n3161 585
R15162 GND.n3161 GND.n3160 585
R15163 GND.n2963 GND.n2962 585
R15164 GND.n2964 GND.n2963 585
R15165 GND.n2961 GND.n1838 585
R15166 GND.n8684 GND.n1838 585
R15167 GND.n2909 GND.n2908 585
R15168 GND.n2908 GND.n2907 585
R15169 GND.n2957 GND.n1819 585
R15170 GND.n8690 GND.n1819 585
R15171 GND.n2956 GND.n2955 585
R15172 GND.n2955 GND.n1817 585
R15173 GND.n2954 GND.n2953 585
R15174 GND.n2954 GND.n1805 585
R15175 GND.n2911 GND.n1804 585
R15176 GND.n8698 GND.n1804 585
R15177 GND.n8460 GND.n8459 585
R15178 GND.n8461 GND.n2142 585
R15179 GND.n8463 GND.n2141 585
R15180 GND.n8464 GND.n2140 585
R15181 GND.n8466 GND.n2139 585
R15182 GND.n8467 GND.n2138 585
R15183 GND.n8469 GND.n2137 585
R15184 GND.n8470 GND.n2136 585
R15185 GND.n8472 GND.n2135 585
R15186 GND.n8473 GND.n2134 585
R15187 GND.n8475 GND.n2133 585
R15188 GND.n8476 GND.n2132 585
R15189 GND.n4727 GND.n4726 502.111
R15190 GND.n4717 GND.n4652 502.111
R15191 GND.n5203 GND.n3750 502.111
R15192 GND.n8125 GND.n3752 502.111
R15193 GND.n10535 GND.n10534 340.337
R15194 GND.n10385 GND.n658 301.784
R15195 GND.n10393 GND.n658 301.784
R15196 GND.n10394 GND.n10393 301.784
R15197 GND.n10395 GND.n10394 301.784
R15198 GND.n10395 GND.n652 301.784
R15199 GND.n10403 GND.n652 301.784
R15200 GND.n10404 GND.n10403 301.784
R15201 GND.n10405 GND.n10404 301.784
R15202 GND.n10405 GND.n646 301.784
R15203 GND.n10413 GND.n646 301.784
R15204 GND.n10414 GND.n10413 301.784
R15205 GND.n10415 GND.n10414 301.784
R15206 GND.n10415 GND.n640 301.784
R15207 GND.n10423 GND.n640 301.784
R15208 GND.n10424 GND.n10423 301.784
R15209 GND.n10425 GND.n10424 301.784
R15210 GND.n10425 GND.n634 301.784
R15211 GND.n10433 GND.n634 301.784
R15212 GND.n10434 GND.n10433 301.784
R15213 GND.n10435 GND.n10434 301.784
R15214 GND.n10435 GND.n628 301.784
R15215 GND.n10443 GND.n628 301.784
R15216 GND.n10444 GND.n10443 301.784
R15217 GND.n10445 GND.n10444 301.784
R15218 GND.n10445 GND.n622 301.784
R15219 GND.n10453 GND.n622 301.784
R15220 GND.n10454 GND.n10453 301.784
R15221 GND.n10455 GND.n10454 301.784
R15222 GND.n10455 GND.n616 301.784
R15223 GND.n10463 GND.n616 301.784
R15224 GND.n10464 GND.n10463 301.784
R15225 GND.n10465 GND.n10464 301.784
R15226 GND.n10465 GND.n610 301.784
R15227 GND.n10473 GND.n610 301.784
R15228 GND.n10474 GND.n10473 301.784
R15229 GND.n10475 GND.n10474 301.784
R15230 GND.n10475 GND.n604 301.784
R15231 GND.n10483 GND.n604 301.784
R15232 GND.n10484 GND.n10483 301.784
R15233 GND.n10485 GND.n10484 301.784
R15234 GND.n10485 GND.n598 301.784
R15235 GND.n10493 GND.n598 301.784
R15236 GND.n10494 GND.n10493 301.784
R15237 GND.n10495 GND.n10494 301.784
R15238 GND.n10495 GND.n592 301.784
R15239 GND.n10503 GND.n592 301.784
R15240 GND.n10504 GND.n10503 301.784
R15241 GND.n10505 GND.n10504 301.784
R15242 GND.n10505 GND.n586 301.784
R15243 GND.n10513 GND.n586 301.784
R15244 GND.n10514 GND.n10513 301.784
R15245 GND.n10515 GND.n10514 301.784
R15246 GND.n10515 GND.n580 301.784
R15247 GND.n10523 GND.n580 301.784
R15248 GND.n10524 GND.n10523 301.784
R15249 GND.n10525 GND.n10524 301.784
R15250 GND.n10525 GND.n574 301.784
R15251 GND.n10534 GND.n574 301.784
R15252 GND.n3759 GND.n3758 294.49
R15253 GND.n4642 GND.n4641 294.49
R15254 GND.n9053 GND.n9052 280.613
R15255 GND.n9054 GND.n9053 280.613
R15256 GND.n9054 GND.n1455 280.613
R15257 GND.n9062 GND.n1455 280.613
R15258 GND.n9063 GND.n9062 280.613
R15259 GND.n9064 GND.n9063 280.613
R15260 GND.n9064 GND.n1449 280.613
R15261 GND.n9072 GND.n1449 280.613
R15262 GND.n9073 GND.n9072 280.613
R15263 GND.n9074 GND.n9073 280.613
R15264 GND.n9074 GND.n1443 280.613
R15265 GND.n9082 GND.n1443 280.613
R15266 GND.n9083 GND.n9082 280.613
R15267 GND.n9084 GND.n9083 280.613
R15268 GND.n9084 GND.n1437 280.613
R15269 GND.n9092 GND.n1437 280.613
R15270 GND.n9093 GND.n9092 280.613
R15271 GND.n9094 GND.n9093 280.613
R15272 GND.n9094 GND.n1431 280.613
R15273 GND.n9102 GND.n1431 280.613
R15274 GND.n9103 GND.n9102 280.613
R15275 GND.n9104 GND.n9103 280.613
R15276 GND.n9104 GND.n1425 280.613
R15277 GND.n9112 GND.n1425 280.613
R15278 GND.n9113 GND.n9112 280.613
R15279 GND.n9114 GND.n9113 280.613
R15280 GND.n9114 GND.n1419 280.613
R15281 GND.n9122 GND.n1419 280.613
R15282 GND.n9123 GND.n9122 280.613
R15283 GND.n9124 GND.n9123 280.613
R15284 GND.n9124 GND.n1413 280.613
R15285 GND.n9132 GND.n1413 280.613
R15286 GND.n9133 GND.n9132 280.613
R15287 GND.n9134 GND.n9133 280.613
R15288 GND.n9134 GND.n1407 280.613
R15289 GND.n9142 GND.n1407 280.613
R15290 GND.n9143 GND.n9142 280.613
R15291 GND.n9144 GND.n9143 280.613
R15292 GND.n9144 GND.n1401 280.613
R15293 GND.n9152 GND.n1401 280.613
R15294 GND.n9153 GND.n9152 280.613
R15295 GND.n9154 GND.n9153 280.613
R15296 GND.n9154 GND.n1395 280.613
R15297 GND.n9162 GND.n1395 280.613
R15298 GND.n9163 GND.n9162 280.613
R15299 GND.n9164 GND.n9163 280.613
R15300 GND.n9164 GND.n1389 280.613
R15301 GND.n9172 GND.n1389 280.613
R15302 GND.n9173 GND.n9172 280.613
R15303 GND.n9174 GND.n9173 280.613
R15304 GND.n9174 GND.n1383 280.613
R15305 GND.n9182 GND.n1383 280.613
R15306 GND.n9183 GND.n9182 280.613
R15307 GND.n9184 GND.n9183 280.613
R15308 GND.n9184 GND.n1377 280.613
R15309 GND.n9192 GND.n1377 280.613
R15310 GND.n9193 GND.n9192 280.613
R15311 GND.n9194 GND.n9193 280.613
R15312 GND.n9194 GND.n1371 280.613
R15313 GND.n9202 GND.n1371 280.613
R15314 GND.n9203 GND.n9202 280.613
R15315 GND.n9204 GND.n9203 280.613
R15316 GND.n9204 GND.n1365 280.613
R15317 GND.n9212 GND.n1365 280.613
R15318 GND.n9213 GND.n9212 280.613
R15319 GND.n9214 GND.n9213 280.613
R15320 GND.n9214 GND.n1359 280.613
R15321 GND.n9222 GND.n1359 280.613
R15322 GND.n9223 GND.n9222 280.613
R15323 GND.n9224 GND.n9223 280.613
R15324 GND.n9224 GND.n1353 280.613
R15325 GND.n9232 GND.n1353 280.613
R15326 GND.n9233 GND.n9232 280.613
R15327 GND.n9234 GND.n9233 280.613
R15328 GND.n9234 GND.n1347 280.613
R15329 GND.n9242 GND.n1347 280.613
R15330 GND.n9243 GND.n9242 280.613
R15331 GND.n9244 GND.n9243 280.613
R15332 GND.n9244 GND.n1341 280.613
R15333 GND.n9252 GND.n1341 280.613
R15334 GND.n9253 GND.n9252 280.613
R15335 GND.n9254 GND.n9253 280.613
R15336 GND.n9254 GND.n1335 280.613
R15337 GND.n9262 GND.n1335 280.613
R15338 GND.n9263 GND.n9262 280.613
R15339 GND.n9264 GND.n9263 280.613
R15340 GND.n9264 GND.n1329 280.613
R15341 GND.n9272 GND.n1329 280.613
R15342 GND.n9273 GND.n9272 280.613
R15343 GND.n9274 GND.n9273 280.613
R15344 GND.n9274 GND.n1323 280.613
R15345 GND.n9282 GND.n1323 280.613
R15346 GND.n9283 GND.n9282 280.613
R15347 GND.n9284 GND.n9283 280.613
R15348 GND.n9284 GND.n1317 280.613
R15349 GND.n9292 GND.n1317 280.613
R15350 GND.n9293 GND.n9292 280.613
R15351 GND.n9294 GND.n9293 280.613
R15352 GND.n9294 GND.n1311 280.613
R15353 GND.n9302 GND.n1311 280.613
R15354 GND.n9303 GND.n9302 280.613
R15355 GND.n9304 GND.n9303 280.613
R15356 GND.n9304 GND.n1305 280.613
R15357 GND.n9312 GND.n1305 280.613
R15358 GND.n9313 GND.n9312 280.613
R15359 GND.n9314 GND.n9313 280.613
R15360 GND.n9314 GND.n1299 280.613
R15361 GND.n9322 GND.n1299 280.613
R15362 GND.n9323 GND.n9322 280.613
R15363 GND.n9324 GND.n9323 280.613
R15364 GND.n9324 GND.n1293 280.613
R15365 GND.n9332 GND.n1293 280.613
R15366 GND.n9333 GND.n9332 280.613
R15367 GND.n9334 GND.n9333 280.613
R15368 GND.n9334 GND.n1287 280.613
R15369 GND.n9342 GND.n1287 280.613
R15370 GND.n9343 GND.n9342 280.613
R15371 GND.n9344 GND.n9343 280.613
R15372 GND.n9344 GND.n1281 280.613
R15373 GND.n9352 GND.n1281 280.613
R15374 GND.n9353 GND.n9352 280.613
R15375 GND.n9354 GND.n9353 280.613
R15376 GND.n9354 GND.n1275 280.613
R15377 GND.n9362 GND.n1275 280.613
R15378 GND.n9363 GND.n9362 280.613
R15379 GND.n9364 GND.n9363 280.613
R15380 GND.n9364 GND.n1269 280.613
R15381 GND.n9372 GND.n1269 280.613
R15382 GND.n9373 GND.n9372 280.613
R15383 GND.n9374 GND.n9373 280.613
R15384 GND.n9374 GND.n1263 280.613
R15385 GND.n9382 GND.n1263 280.613
R15386 GND.n9383 GND.n9382 280.613
R15387 GND.n9384 GND.n9383 280.613
R15388 GND.n9384 GND.n1257 280.613
R15389 GND.n9392 GND.n1257 280.613
R15390 GND.n9393 GND.n9392 280.613
R15391 GND.n9394 GND.n9393 280.613
R15392 GND.n9394 GND.n1251 280.613
R15393 GND.n9402 GND.n1251 280.613
R15394 GND.n9403 GND.n9402 280.613
R15395 GND.n9404 GND.n9403 280.613
R15396 GND.n9404 GND.n1245 280.613
R15397 GND.n9412 GND.n1245 280.613
R15398 GND.n9413 GND.n9412 280.613
R15399 GND.n9414 GND.n9413 280.613
R15400 GND.n9414 GND.n1239 280.613
R15401 GND.n9422 GND.n1239 280.613
R15402 GND.n9423 GND.n9422 280.613
R15403 GND.n9424 GND.n9423 280.613
R15404 GND.n9424 GND.n1233 280.613
R15405 GND.n9432 GND.n1233 280.613
R15406 GND.n9433 GND.n9432 280.613
R15407 GND.n9434 GND.n9433 280.613
R15408 GND.n9434 GND.n1227 280.613
R15409 GND.n9442 GND.n1227 280.613
R15410 GND.n9443 GND.n9442 280.613
R15411 GND.n9444 GND.n9443 280.613
R15412 GND.n9444 GND.n1221 280.613
R15413 GND.n9452 GND.n1221 280.613
R15414 GND.n9453 GND.n9452 280.613
R15415 GND.n9454 GND.n9453 280.613
R15416 GND.n9454 GND.n1215 280.613
R15417 GND.n9462 GND.n1215 280.613
R15418 GND.n9463 GND.n9462 280.613
R15419 GND.n9464 GND.n9463 280.613
R15420 GND.n9464 GND.n1209 280.613
R15421 GND.n9472 GND.n1209 280.613
R15422 GND.n9473 GND.n9472 280.613
R15423 GND.n9474 GND.n9473 280.613
R15424 GND.n9474 GND.n1203 280.613
R15425 GND.n9482 GND.n1203 280.613
R15426 GND.n9483 GND.n9482 280.613
R15427 GND.n9484 GND.n9483 280.613
R15428 GND.n9484 GND.n1197 280.613
R15429 GND.n9492 GND.n1197 280.613
R15430 GND.n9493 GND.n9492 280.613
R15431 GND.n9494 GND.n9493 280.613
R15432 GND.n9494 GND.n1191 280.613
R15433 GND.n9502 GND.n1191 280.613
R15434 GND.n9503 GND.n9502 280.613
R15435 GND.n9504 GND.n9503 280.613
R15436 GND.n9504 GND.n1185 280.613
R15437 GND.n9512 GND.n1185 280.613
R15438 GND.n9513 GND.n9512 280.613
R15439 GND.n9514 GND.n9513 280.613
R15440 GND.n9514 GND.n1179 280.613
R15441 GND.n9522 GND.n1179 280.613
R15442 GND.n9523 GND.n9522 280.613
R15443 GND.n9524 GND.n9523 280.613
R15444 GND.n9524 GND.n1173 280.613
R15445 GND.n9532 GND.n1173 280.613
R15446 GND.n9533 GND.n9532 280.613
R15447 GND.n9534 GND.n9533 280.613
R15448 GND.n9534 GND.n1167 280.613
R15449 GND.n9542 GND.n1167 280.613
R15450 GND.n9543 GND.n9542 280.613
R15451 GND.n9544 GND.n9543 280.613
R15452 GND.n9544 GND.n1161 280.613
R15453 GND.n9552 GND.n1161 280.613
R15454 GND.n9553 GND.n9552 280.613
R15455 GND.n9554 GND.n9553 280.613
R15456 GND.n9554 GND.n1155 280.613
R15457 GND.n9562 GND.n1155 280.613
R15458 GND.n9563 GND.n9562 280.613
R15459 GND.n9564 GND.n9563 280.613
R15460 GND.n9564 GND.n1149 280.613
R15461 GND.n9572 GND.n1149 280.613
R15462 GND.n9573 GND.n9572 280.613
R15463 GND.n9574 GND.n9573 280.613
R15464 GND.n9574 GND.n1143 280.613
R15465 GND.n9582 GND.n1143 280.613
R15466 GND.n9583 GND.n9582 280.613
R15467 GND.n9584 GND.n9583 280.613
R15468 GND.n9584 GND.n1137 280.613
R15469 GND.n9592 GND.n1137 280.613
R15470 GND.n9593 GND.n9592 280.613
R15471 GND.n9594 GND.n9593 280.613
R15472 GND.n9594 GND.n1131 280.613
R15473 GND.n9602 GND.n1131 280.613
R15474 GND.n9603 GND.n9602 280.613
R15475 GND.n9604 GND.n9603 280.613
R15476 GND.n9604 GND.n1125 280.613
R15477 GND.n9612 GND.n1125 280.613
R15478 GND.n9613 GND.n9612 280.613
R15479 GND.n9614 GND.n9613 280.613
R15480 GND.n9614 GND.n1119 280.613
R15481 GND.n9622 GND.n1119 280.613
R15482 GND.n9623 GND.n9622 280.613
R15483 GND.n9624 GND.n9623 280.613
R15484 GND.n9624 GND.n1113 280.613
R15485 GND.n9632 GND.n1113 280.613
R15486 GND.n9633 GND.n9632 280.613
R15487 GND.n9634 GND.n9633 280.613
R15488 GND.n9634 GND.n1107 280.613
R15489 GND.n9642 GND.n1107 280.613
R15490 GND.n9643 GND.n9642 280.613
R15491 GND.n9644 GND.n9643 280.613
R15492 GND.n9644 GND.n1101 280.613
R15493 GND.n9652 GND.n1101 280.613
R15494 GND.n9653 GND.n9652 280.613
R15495 GND.n9654 GND.n9653 280.613
R15496 GND.n9654 GND.n1095 280.613
R15497 GND.n9662 GND.n1095 280.613
R15498 GND.n9663 GND.n9662 280.613
R15499 GND.n9664 GND.n9663 280.613
R15500 GND.n9664 GND.n1089 280.613
R15501 GND.n9672 GND.n1089 280.613
R15502 GND.n9673 GND.n9672 280.613
R15503 GND.n9674 GND.n9673 280.613
R15504 GND.n9674 GND.n1083 280.613
R15505 GND.n9682 GND.n1083 280.613
R15506 GND.n9683 GND.n9682 280.613
R15507 GND.n9684 GND.n9683 280.613
R15508 GND.n9684 GND.n1077 280.613
R15509 GND.n9692 GND.n1077 280.613
R15510 GND.n9693 GND.n9692 280.613
R15511 GND.n9694 GND.n9693 280.613
R15512 GND.n9694 GND.n1071 280.613
R15513 GND.n9702 GND.n1071 280.613
R15514 GND.n9703 GND.n9702 280.613
R15515 GND.n9704 GND.n9703 280.613
R15516 GND.n9704 GND.n1065 280.613
R15517 GND.n9712 GND.n1065 280.613
R15518 GND.n9713 GND.n9712 280.613
R15519 GND.n9714 GND.n9713 280.613
R15520 GND.n9714 GND.n1059 280.613
R15521 GND.n9722 GND.n1059 280.613
R15522 GND.n9723 GND.n9722 280.613
R15523 GND.n9724 GND.n9723 280.613
R15524 GND.n9724 GND.n1053 280.613
R15525 GND.n9732 GND.n1053 280.613
R15526 GND.n9733 GND.n9732 280.613
R15527 GND.n9734 GND.n9733 280.613
R15528 GND.n9734 GND.n1047 280.613
R15529 GND.n9742 GND.n1047 280.613
R15530 GND.n9743 GND.n9742 280.613
R15531 GND.n9744 GND.n9743 280.613
R15532 GND.n9744 GND.n1041 280.613
R15533 GND.n9752 GND.n1041 280.613
R15534 GND.n9753 GND.n9752 280.613
R15535 GND.n9754 GND.n9753 280.613
R15536 GND.n9754 GND.n1035 280.613
R15537 GND.n9762 GND.n1035 280.613
R15538 GND.n9763 GND.n9762 280.613
R15539 GND.n9764 GND.n9763 280.613
R15540 GND.n9764 GND.n1029 280.613
R15541 GND.n9772 GND.n1029 280.613
R15542 GND.n9773 GND.n9772 280.613
R15543 GND.n9774 GND.n9773 280.613
R15544 GND.n9774 GND.n1023 280.613
R15545 GND.n9782 GND.n1023 280.613
R15546 GND.n9783 GND.n9782 280.613
R15547 GND.n9784 GND.n9783 280.613
R15548 GND.n9784 GND.n1017 280.613
R15549 GND.n9792 GND.n1017 280.613
R15550 GND.n9793 GND.n9792 280.613
R15551 GND.n9794 GND.n9793 280.613
R15552 GND.n9794 GND.n1011 280.613
R15553 GND.n9802 GND.n1011 280.613
R15554 GND.n9803 GND.n9802 280.613
R15555 GND.n9804 GND.n9803 280.613
R15556 GND.n9804 GND.n1005 280.613
R15557 GND.n9812 GND.n1005 280.613
R15558 GND.n9813 GND.n9812 280.613
R15559 GND.n9814 GND.n9813 280.613
R15560 GND.n9814 GND.n999 280.613
R15561 GND.n9822 GND.n999 280.613
R15562 GND.n9823 GND.n9822 280.613
R15563 GND.n9824 GND.n9823 280.613
R15564 GND.n9824 GND.n993 280.613
R15565 GND.n9832 GND.n993 280.613
R15566 GND.n9833 GND.n9832 280.613
R15567 GND.n9834 GND.n9833 280.613
R15568 GND.n9834 GND.n987 280.613
R15569 GND.n9842 GND.n987 280.613
R15570 GND.n9843 GND.n9842 280.613
R15571 GND.n9844 GND.n9843 280.613
R15572 GND.n9844 GND.n981 280.613
R15573 GND.n9852 GND.n981 280.613
R15574 GND.n9853 GND.n9852 280.613
R15575 GND.n9854 GND.n9853 280.613
R15576 GND.n9854 GND.n975 280.613
R15577 GND.n9862 GND.n975 280.613
R15578 GND.n9863 GND.n9862 280.613
R15579 GND.n9864 GND.n9863 280.613
R15580 GND.n9864 GND.n969 280.613
R15581 GND.n9872 GND.n969 280.613
R15582 GND.n9873 GND.n9872 280.613
R15583 GND.n9874 GND.n9873 280.613
R15584 GND.n9874 GND.n963 280.613
R15585 GND.n9882 GND.n963 280.613
R15586 GND.n9883 GND.n9882 280.613
R15587 GND.n9884 GND.n9883 280.613
R15588 GND.n9884 GND.n957 280.613
R15589 GND.n9892 GND.n957 280.613
R15590 GND.n9893 GND.n9892 280.613
R15591 GND.n9894 GND.n9893 280.613
R15592 GND.n9894 GND.n951 280.613
R15593 GND.n9902 GND.n951 280.613
R15594 GND.n9903 GND.n9902 280.613
R15595 GND.n9904 GND.n9903 280.613
R15596 GND.n9904 GND.n945 280.613
R15597 GND.n9912 GND.n945 280.613
R15598 GND.n9913 GND.n9912 280.613
R15599 GND.n9914 GND.n9913 280.613
R15600 GND.n9914 GND.n939 280.613
R15601 GND.n9922 GND.n939 280.613
R15602 GND.n9923 GND.n9922 280.613
R15603 GND.n9924 GND.n9923 280.613
R15604 GND.n9924 GND.n933 280.613
R15605 GND.n9932 GND.n933 280.613
R15606 GND.n9933 GND.n9932 280.613
R15607 GND.n9934 GND.n9933 280.613
R15608 GND.n9934 GND.n927 280.613
R15609 GND.n9942 GND.n927 280.613
R15610 GND.n9943 GND.n9942 280.613
R15611 GND.n9944 GND.n9943 280.613
R15612 GND.n9944 GND.n921 280.613
R15613 GND.n9952 GND.n921 280.613
R15614 GND.n9953 GND.n9952 280.613
R15615 GND.n9954 GND.n9953 280.613
R15616 GND.n9954 GND.n915 280.613
R15617 GND.n9962 GND.n915 280.613
R15618 GND.n9963 GND.n9962 280.613
R15619 GND.n9964 GND.n9963 280.613
R15620 GND.n9964 GND.n909 280.613
R15621 GND.n9972 GND.n909 280.613
R15622 GND.n9973 GND.n9972 280.613
R15623 GND.n9974 GND.n9973 280.613
R15624 GND.n9974 GND.n903 280.613
R15625 GND.n9982 GND.n903 280.613
R15626 GND.n9983 GND.n9982 280.613
R15627 GND.n9984 GND.n9983 280.613
R15628 GND.n9984 GND.n897 280.613
R15629 GND.n9992 GND.n897 280.613
R15630 GND.n9993 GND.n9992 280.613
R15631 GND.n9994 GND.n9993 280.613
R15632 GND.n9994 GND.n891 280.613
R15633 GND.n10002 GND.n891 280.613
R15634 GND.n10003 GND.n10002 280.613
R15635 GND.n10004 GND.n10003 280.613
R15636 GND.n10004 GND.n885 280.613
R15637 GND.n10012 GND.n885 280.613
R15638 GND.n10013 GND.n10012 280.613
R15639 GND.n10014 GND.n10013 280.613
R15640 GND.n10014 GND.n879 280.613
R15641 GND.n10022 GND.n879 280.613
R15642 GND.n10023 GND.n10022 280.613
R15643 GND.n10024 GND.n10023 280.613
R15644 GND.n10024 GND.n873 280.613
R15645 GND.n10032 GND.n873 280.613
R15646 GND.n10033 GND.n10032 280.613
R15647 GND.n10034 GND.n10033 280.613
R15648 GND.n10034 GND.n867 280.613
R15649 GND.n10042 GND.n867 280.613
R15650 GND.n10043 GND.n10042 280.613
R15651 GND.n10044 GND.n10043 280.613
R15652 GND.n10044 GND.n861 280.613
R15653 GND.n10052 GND.n861 280.613
R15654 GND.n10053 GND.n10052 280.613
R15655 GND.n10054 GND.n10053 280.613
R15656 GND.n10054 GND.n855 280.613
R15657 GND.n10062 GND.n855 280.613
R15658 GND.n10063 GND.n10062 280.613
R15659 GND.n10064 GND.n10063 280.613
R15660 GND.n10064 GND.n849 280.613
R15661 GND.n10072 GND.n849 280.613
R15662 GND.n10073 GND.n10072 280.613
R15663 GND.n10074 GND.n10073 280.613
R15664 GND.n10074 GND.n843 280.613
R15665 GND.n10082 GND.n843 280.613
R15666 GND.n10083 GND.n10082 280.613
R15667 GND.n10084 GND.n10083 280.613
R15668 GND.n10084 GND.n837 280.613
R15669 GND.n10092 GND.n837 280.613
R15670 GND.n10093 GND.n10092 280.613
R15671 GND.n10094 GND.n10093 280.613
R15672 GND.n10094 GND.n831 280.613
R15673 GND.n10102 GND.n831 280.613
R15674 GND.n10103 GND.n10102 280.613
R15675 GND.n10104 GND.n10103 280.613
R15676 GND.n10104 GND.n825 280.613
R15677 GND.n10112 GND.n825 280.613
R15678 GND.n10113 GND.n10112 280.613
R15679 GND.n10114 GND.n10113 280.613
R15680 GND.n10114 GND.n819 280.613
R15681 GND.n10122 GND.n819 280.613
R15682 GND.n10123 GND.n10122 280.613
R15683 GND.n10124 GND.n10123 280.613
R15684 GND.n10124 GND.n813 280.613
R15685 GND.n10132 GND.n813 280.613
R15686 GND.n10133 GND.n10132 280.613
R15687 GND.n10134 GND.n10133 280.613
R15688 GND.n10134 GND.n807 280.613
R15689 GND.n10142 GND.n807 280.613
R15690 GND.n10143 GND.n10142 280.613
R15691 GND.n10144 GND.n10143 280.613
R15692 GND.n10144 GND.n801 280.613
R15693 GND.n10152 GND.n801 280.613
R15694 GND.n10153 GND.n10152 280.613
R15695 GND.n10154 GND.n10153 280.613
R15696 GND.n10154 GND.n795 280.613
R15697 GND.n10162 GND.n795 280.613
R15698 GND.n10163 GND.n10162 280.613
R15699 GND.n10164 GND.n10163 280.613
R15700 GND.n10164 GND.n789 280.613
R15701 GND.n10172 GND.n789 280.613
R15702 GND.n10173 GND.n10172 280.613
R15703 GND.n10174 GND.n10173 280.613
R15704 GND.n10174 GND.n783 280.613
R15705 GND.n10182 GND.n783 280.613
R15706 GND.n10183 GND.n10182 280.613
R15707 GND.n10184 GND.n10183 280.613
R15708 GND.n10184 GND.n777 280.613
R15709 GND.n10192 GND.n777 280.613
R15710 GND.n10193 GND.n10192 280.613
R15711 GND.n10194 GND.n10193 280.613
R15712 GND.n10194 GND.n771 280.613
R15713 GND.n10202 GND.n771 280.613
R15714 GND.n10203 GND.n10202 280.613
R15715 GND.n10204 GND.n10203 280.613
R15716 GND.n10204 GND.n765 280.613
R15717 GND.n10212 GND.n765 280.613
R15718 GND.n10213 GND.n10212 280.613
R15719 GND.n10214 GND.n10213 280.613
R15720 GND.n10214 GND.n759 280.613
R15721 GND.n10222 GND.n759 280.613
R15722 GND.n10223 GND.n10222 280.613
R15723 GND.n10224 GND.n10223 280.613
R15724 GND.n10224 GND.n753 280.613
R15725 GND.n10232 GND.n753 280.613
R15726 GND.n10233 GND.n10232 280.613
R15727 GND.n10234 GND.n10233 280.613
R15728 GND.n10234 GND.n747 280.613
R15729 GND.n10242 GND.n747 280.613
R15730 GND.n10243 GND.n10242 280.613
R15731 GND.n10244 GND.n10243 280.613
R15732 GND.n10244 GND.n741 280.613
R15733 GND.n10252 GND.n741 280.613
R15734 GND.n10253 GND.n10252 280.613
R15735 GND.n10254 GND.n10253 280.613
R15736 GND.n10254 GND.n735 280.613
R15737 GND.n10262 GND.n735 280.613
R15738 GND.n10263 GND.n10262 280.613
R15739 GND.n10264 GND.n10263 280.613
R15740 GND.n10264 GND.n729 280.613
R15741 GND.n10272 GND.n729 280.613
R15742 GND.n10273 GND.n10272 280.613
R15743 GND.n10274 GND.n10273 280.613
R15744 GND.n10274 GND.n723 280.613
R15745 GND.n10282 GND.n723 280.613
R15746 GND.n10283 GND.n10282 280.613
R15747 GND.n10284 GND.n10283 280.613
R15748 GND.n10284 GND.n717 280.613
R15749 GND.n10292 GND.n717 280.613
R15750 GND.n10293 GND.n10292 280.613
R15751 GND.n10294 GND.n10293 280.613
R15752 GND.n10294 GND.n711 280.613
R15753 GND.n10302 GND.n711 280.613
R15754 GND.n10303 GND.n10302 280.613
R15755 GND.n10304 GND.n10303 280.613
R15756 GND.n10304 GND.n705 280.613
R15757 GND.n10312 GND.n705 280.613
R15758 GND.n10313 GND.n10312 280.613
R15759 GND.n10314 GND.n10313 280.613
R15760 GND.n10314 GND.n699 280.613
R15761 GND.n10322 GND.n699 280.613
R15762 GND.n10323 GND.n10322 280.613
R15763 GND.n10324 GND.n10323 280.613
R15764 GND.n10324 GND.n693 280.613
R15765 GND.n10332 GND.n693 280.613
R15766 GND.n10333 GND.n10332 280.613
R15767 GND.n10334 GND.n10333 280.613
R15768 GND.n10334 GND.n687 280.613
R15769 GND.n10342 GND.n687 280.613
R15770 GND.n10343 GND.n10342 280.613
R15771 GND.n10344 GND.n10343 280.613
R15772 GND.n10344 GND.n681 280.613
R15773 GND.n10352 GND.n681 280.613
R15774 GND.n10353 GND.n10352 280.613
R15775 GND.n10354 GND.n10353 280.613
R15776 GND.n10354 GND.n675 280.613
R15777 GND.n10362 GND.n675 280.613
R15778 GND.n10363 GND.n10362 280.613
R15779 GND.n10364 GND.n10363 280.613
R15780 GND.n10364 GND.n669 280.613
R15781 GND.n10372 GND.n669 280.613
R15782 GND.n10373 GND.n10372 280.613
R15783 GND.n10374 GND.n10373 280.613
R15784 GND.n10374 GND.n663 280.613
R15785 GND.n10383 GND.n663 280.613
R15786 GND.n10384 GND.n10383 280.613
R15787 GND.n5080 GND.n3749 256.663
R15788 GND.n5086 GND.n3749 256.663
R15789 GND.n5088 GND.n3749 256.663
R15790 GND.n5094 GND.n3749 256.663
R15791 GND.n5096 GND.n3749 256.663
R15792 GND.n5102 GND.n3749 256.663
R15793 GND.n5104 GND.n3749 256.663
R15794 GND.n5110 GND.n3749 256.663
R15795 GND.n5112 GND.n3749 256.663
R15796 GND.n5118 GND.n3749 256.663
R15797 GND.n5120 GND.n3749 256.663
R15798 GND.n5126 GND.n3749 256.663
R15799 GND.n5128 GND.n3749 256.663
R15800 GND.n5135 GND.n3749 256.663
R15801 GND.n5138 GND.n3749 256.663
R15802 GND.n5060 GND.n3749 256.663
R15803 GND.n5144 GND.n3749 256.663
R15804 GND.n5146 GND.n3749 256.663
R15805 GND.n5153 GND.n3749 256.663
R15806 GND.n5155 GND.n3749 256.663
R15807 GND.n5161 GND.n3749 256.663
R15808 GND.n5163 GND.n3749 256.663
R15809 GND.n5169 GND.n3749 256.663
R15810 GND.n5171 GND.n3749 256.663
R15811 GND.n5177 GND.n3749 256.663
R15812 GND.n5179 GND.n3749 256.663
R15813 GND.n5185 GND.n3749 256.663
R15814 GND.n5187 GND.n3749 256.663
R15815 GND.n5193 GND.n3749 256.663
R15816 GND.n5195 GND.n3749 256.663
R15817 GND.n5201 GND.n3749 256.663
R15818 GND.n7657 GND.n4559 256.663
R15819 GND.n7657 GND.n4558 256.663
R15820 GND.n7657 GND.n4557 256.663
R15821 GND.n7657 GND.n4556 256.663
R15822 GND.n7657 GND.n4555 256.663
R15823 GND.n7657 GND.n4554 256.663
R15824 GND.n7657 GND.n4553 256.663
R15825 GND.n7657 GND.n4552 256.663
R15826 GND.n7657 GND.n4551 256.663
R15827 GND.n7657 GND.n4550 256.663
R15828 GND.n7657 GND.n4549 256.663
R15829 GND.n7657 GND.n4548 256.663
R15830 GND.n7657 GND.n4547 256.663
R15831 GND.n7657 GND.n4546 256.663
R15832 GND.n7657 GND.n4545 256.663
R15833 GND.n7657 GND.n4544 256.663
R15834 GND.n4791 GND.n4790 256.663
R15835 GND.n7657 GND.n4543 256.663
R15836 GND.n7657 GND.n4542 256.663
R15837 GND.n7657 GND.n4541 256.663
R15838 GND.n7657 GND.n4540 256.663
R15839 GND.n7657 GND.n4539 256.663
R15840 GND.n7657 GND.n4538 256.663
R15841 GND.n7657 GND.n4537 256.663
R15842 GND.n7657 GND.n4536 256.663
R15843 GND.n7657 GND.n4535 256.663
R15844 GND.n7657 GND.n4534 256.663
R15845 GND.n7657 GND.n4533 256.663
R15846 GND.n7657 GND.n4532 256.663
R15847 GND.n7657 GND.n4531 256.663
R15848 GND.n7657 GND.n4530 256.663
R15849 GND.n7657 GND.n4529 256.663
R15850 GND.n7657 GND.n4528 256.663
R15851 GND.n5065 GND.t129 250.794
R15852 GND.n5056 GND.t139 250.794
R15853 GND.n4655 GND.t66 250.794
R15854 GND.n4635 GND.t49 250.794
R15855 GND.n7647 GND.n4595 242.672
R15856 GND.n7647 GND.n4596 242.672
R15857 GND.n7647 GND.n4597 242.672
R15858 GND.n7647 GND.n4598 242.672
R15859 GND.n7647 GND.n4599 242.672
R15860 GND.n7647 GND.n4600 242.672
R15861 GND.n7647 GND.n4601 242.672
R15862 GND.n10897 GND.n10896 242.672
R15863 GND.n10896 GND.n10647 242.672
R15864 GND.n10896 GND.n10648 242.672
R15865 GND.n10896 GND.n10649 242.672
R15866 GND.n10896 GND.n10650 242.672
R15867 GND.n10896 GND.n10651 242.672
R15868 GND.n10896 GND.n10687 242.672
R15869 GND.n8056 GND.n8055 242.672
R15870 GND.n8056 GND.n3851 242.672
R15871 GND.n8056 GND.n3852 242.672
R15872 GND.n8056 GND.n3853 242.672
R15873 GND.n8056 GND.n3854 242.672
R15874 GND.n8056 GND.n3855 242.672
R15875 GND.n8056 GND.n3856 242.672
R15876 GND.n8056 GND.n3857 242.672
R15877 GND.n8056 GND.n3858 242.672
R15878 GND.n8056 GND.n3859 242.672
R15879 GND.n8056 GND.n3860 242.672
R15880 GND.n5869 GND.n4376 242.672
R15881 GND.n5866 GND.n4376 242.672
R15882 GND.n5858 GND.n4376 242.672
R15883 GND.n5853 GND.n4376 242.672
R15884 GND.n5848 GND.n4376 242.672
R15885 GND.n5843 GND.n4376 242.672
R15886 GND.n5838 GND.n4376 242.672
R15887 GND.n5834 GND.n4376 242.672
R15888 GND.n4845 GND.n4376 242.672
R15889 GND.n5826 GND.n4376 242.672
R15890 GND.n5817 GND.n4376 242.672
R15891 GND.n8816 GND.n8815 242.672
R15892 GND.n8816 GND.n1691 242.672
R15893 GND.n8816 GND.n1692 242.672
R15894 GND.n8816 GND.n1693 242.672
R15895 GND.n8816 GND.n1694 242.672
R15896 GND.n8816 GND.n1695 242.672
R15897 GND.n8816 GND.n1696 242.672
R15898 GND.n8816 GND.n1697 242.672
R15899 GND.n8816 GND.n1698 242.672
R15900 GND.n8816 GND.n1699 242.672
R15901 GND.n8816 GND.n1700 242.672
R15902 GND.n8816 GND.n1701 242.672
R15903 GND.n8816 GND.n1702 242.672
R15904 GND.n8816 GND.n1703 242.672
R15905 GND.n8816 GND.n1704 242.672
R15906 GND.n8816 GND.n1705 242.672
R15907 GND.n8816 GND.n1706 242.672
R15908 GND.n8816 GND.n1707 242.672
R15909 GND.n8816 GND.n1708 242.672
R15910 GND.n8816 GND.n1709 242.672
R15911 GND.n8816 GND.n1710 242.672
R15912 GND.n8816 GND.n1711 242.672
R15913 GND.n8816 GND.n1712 242.672
R15914 GND.n8816 GND.n1713 242.672
R15915 GND.n8816 GND.n1714 242.672
R15916 GND.n8816 GND.n1715 242.672
R15917 GND.n8816 GND.n1716 242.672
R15918 GND.n8816 GND.n1717 242.672
R15919 GND.n8457 GND.n2167 242.672
R15920 GND.n8457 GND.n2168 242.672
R15921 GND.n8457 GND.n2169 242.672
R15922 GND.n8457 GND.n2170 242.672
R15923 GND.n8457 GND.n2171 242.672
R15924 GND.n8457 GND.n2172 242.672
R15925 GND.n8457 GND.n2173 242.672
R15926 GND.n8457 GND.n2174 242.672
R15927 GND.n8457 GND.n2175 242.672
R15928 GND.n8457 GND.n2176 242.672
R15929 GND.n8457 GND.n2177 242.672
R15930 GND.n8457 GND.n2178 242.672
R15931 GND.n8457 GND.n2179 242.672
R15932 GND.n8457 GND.n2180 242.672
R15933 GND.n8457 GND.n2181 242.672
R15934 GND.n2185 GND.n2182 242.672
R15935 GND.n8457 GND.n2160 242.672
R15936 GND.n8457 GND.n2159 242.672
R15937 GND.n8457 GND.n2158 242.672
R15938 GND.n8457 GND.n2157 242.672
R15939 GND.n8457 GND.n2156 242.672
R15940 GND.n8457 GND.n2155 242.672
R15941 GND.n8457 GND.n2154 242.672
R15942 GND.n8457 GND.n2153 242.672
R15943 GND.n8457 GND.n2152 242.672
R15944 GND.n8457 GND.n2151 242.672
R15945 GND.n8457 GND.n2150 242.672
R15946 GND.n8457 GND.n2149 242.672
R15947 GND.n8457 GND.n2148 242.672
R15948 GND.n7647 GND.n7646 242.672
R15949 GND.n7647 GND.n4568 242.672
R15950 GND.n7647 GND.n4569 242.672
R15951 GND.n7647 GND.n4570 242.672
R15952 GND.n7647 GND.n4571 242.672
R15953 GND.n7647 GND.n4572 242.672
R15954 GND.n7647 GND.n4573 242.672
R15955 GND.n7647 GND.n4574 242.672
R15956 GND.n7647 GND.n4575 242.672
R15957 GND.n7647 GND.n4576 242.672
R15958 GND.n7647 GND.n4577 242.672
R15959 GND.n7647 GND.n4578 242.672
R15960 GND.n7647 GND.n4579 242.672
R15961 GND.n7647 GND.n4580 242.672
R15962 GND.n7647 GND.n4581 242.672
R15963 GND.n7647 GND.n4582 242.672
R15964 GND.n7647 GND.n4583 242.672
R15965 GND.n7647 GND.n4584 242.672
R15966 GND.n7647 GND.n4585 242.672
R15967 GND.n7647 GND.n4586 242.672
R15968 GND.n7647 GND.n4587 242.672
R15969 GND.n7647 GND.n4588 242.672
R15970 GND.n7647 GND.n4589 242.672
R15971 GND.n7647 GND.n4590 242.672
R15972 GND.n7647 GND.n4591 242.672
R15973 GND.n7647 GND.n4592 242.672
R15974 GND.n7647 GND.n4593 242.672
R15975 GND.n7647 GND.n4594 242.672
R15976 GND.n10896 GND.n10688 242.672
R15977 GND.n10896 GND.n10689 242.672
R15978 GND.n10896 GND.n10690 242.672
R15979 GND.n10896 GND.n10691 242.672
R15980 GND.n10896 GND.n10692 242.672
R15981 GND.n10896 GND.n10693 242.672
R15982 GND.n10896 GND.n10694 242.672
R15983 GND.n10896 GND.n10695 242.672
R15984 GND.n10896 GND.n10696 242.672
R15985 GND.n10896 GND.n10697 242.672
R15986 GND.n10896 GND.n10698 242.672
R15987 GND.n10896 GND.n10699 242.672
R15988 GND.n10896 GND.n10700 242.672
R15989 GND.n10896 GND.n10701 242.672
R15990 GND.n10896 GND.n10702 242.672
R15991 GND.n10896 GND.n10703 242.672
R15992 GND.n10896 GND.n10704 242.672
R15993 GND.n10896 GND.n10705 242.672
R15994 GND.n10896 GND.n10706 242.672
R15995 GND.n10896 GND.n10707 242.672
R15996 GND.n10896 GND.n10708 242.672
R15997 GND.n10896 GND.n10709 242.672
R15998 GND.n10896 GND.n10710 242.672
R15999 GND.n10896 GND.n10711 242.672
R16000 GND.n10896 GND.n10712 242.672
R16001 GND.n10896 GND.n10713 242.672
R16002 GND.n10896 GND.n10714 242.672
R16003 GND.n10896 GND.n10895 242.672
R16004 GND.n8816 GND.n1718 242.672
R16005 GND.n8816 GND.n1719 242.672
R16006 GND.n8816 GND.n1720 242.672
R16007 GND.n8816 GND.n1721 242.672
R16008 GND.n8816 GND.n1722 242.672
R16009 GND.n8816 GND.n1723 242.672
R16010 GND.n8816 GND.n1724 242.672
R16011 GND.n8458 GND.n8457 242.672
R16012 GND.n8457 GND.n2165 242.672
R16013 GND.n8457 GND.n2164 242.672
R16014 GND.n8457 GND.n2163 242.672
R16015 GND.n8457 GND.n2162 242.672
R16016 GND.n8457 GND.n2161 242.672
R16017 GND.n8457 GND.n2130 242.672
R16018 GND.n10715 GND.n444 240.244
R16019 GND.n10894 GND.n10716 240.244
R16020 GND.n10890 GND.n10889 240.244
R16021 GND.n10886 GND.n10885 240.244
R16022 GND.n10882 GND.n10881 240.244
R16023 GND.n10878 GND.n10877 240.244
R16024 GND.n10735 GND.n10734 240.244
R16025 GND.n10870 GND.n10869 240.244
R16026 GND.n10866 GND.n10865 240.244
R16027 GND.n10862 GND.n10861 240.244
R16028 GND.n10858 GND.n10857 240.244
R16029 GND.n10854 GND.n10853 240.244
R16030 GND.n10850 GND.n10849 240.244
R16031 GND.n10846 GND.n10845 240.244
R16032 GND.n10842 GND.n10841 240.244
R16033 GND.n10838 GND.n10837 240.244
R16034 GND.n10834 GND.n10833 240.244
R16035 GND.n10830 GND.n10829 240.244
R16036 GND.n10826 GND.n10825 240.244
R16037 GND.n10822 GND.n10821 240.244
R16038 GND.n10818 GND.n10817 240.244
R16039 GND.n10814 GND.n10813 240.244
R16040 GND.n10810 GND.n10809 240.244
R16041 GND.n10806 GND.n10805 240.244
R16042 GND.n10802 GND.n10801 240.244
R16043 GND.n10798 GND.n10797 240.244
R16044 GND.n10794 GND.n10793 240.244
R16045 GND.n10790 GND.n10789 240.244
R16046 GND.n7533 GND.n5878 240.244
R16047 GND.n6744 GND.n5878 240.244
R16048 GND.n6744 GND.n5930 240.244
R16049 GND.n6754 GND.n5930 240.244
R16050 GND.n6754 GND.n5941 240.244
R16051 GND.n6759 GND.n5941 240.244
R16052 GND.n6759 GND.n5952 240.244
R16053 GND.n6769 GND.n5952 240.244
R16054 GND.n6769 GND.n5961 240.244
R16055 GND.n6774 GND.n5961 240.244
R16056 GND.n6774 GND.n5972 240.244
R16057 GND.n6784 GND.n5972 240.244
R16058 GND.n6784 GND.n5982 240.244
R16059 GND.n6789 GND.n5982 240.244
R16060 GND.n6789 GND.n5993 240.244
R16061 GND.n6799 GND.n5993 240.244
R16062 GND.n6799 GND.n6003 240.244
R16063 GND.n6804 GND.n6003 240.244
R16064 GND.n6804 GND.n6014 240.244
R16065 GND.n6814 GND.n6014 240.244
R16066 GND.n6814 GND.n6024 240.244
R16067 GND.n6819 GND.n6024 240.244
R16068 GND.n6819 GND.n6035 240.244
R16069 GND.n6829 GND.n6035 240.244
R16070 GND.n6829 GND.n6044 240.244
R16071 GND.n6834 GND.n6044 240.244
R16072 GND.n6834 GND.n6055 240.244
R16073 GND.n6844 GND.n6055 240.244
R16074 GND.n6844 GND.n6065 240.244
R16075 GND.n6849 GND.n6065 240.244
R16076 GND.n6849 GND.n6076 240.244
R16077 GND.n6859 GND.n6076 240.244
R16078 GND.n6859 GND.n6086 240.244
R16079 GND.n6864 GND.n6086 240.244
R16080 GND.n6864 GND.n6097 240.244
R16081 GND.n6874 GND.n6097 240.244
R16082 GND.n6874 GND.n6107 240.244
R16083 GND.n6879 GND.n6107 240.244
R16084 GND.n6879 GND.n6118 240.244
R16085 GND.n6889 GND.n6118 240.244
R16086 GND.n6889 GND.n6128 240.244
R16087 GND.n6894 GND.n6128 240.244
R16088 GND.n6894 GND.n6139 240.244
R16089 GND.n6904 GND.n6139 240.244
R16090 GND.n6904 GND.n6149 240.244
R16091 GND.n6909 GND.n6149 240.244
R16092 GND.n6909 GND.n6160 240.244
R16093 GND.n6919 GND.n6160 240.244
R16094 GND.n6919 GND.n6170 240.244
R16095 GND.n6924 GND.n6170 240.244
R16096 GND.n6924 GND.n6180 240.244
R16097 GND.n6934 GND.n6180 240.244
R16098 GND.n6934 GND.n6190 240.244
R16099 GND.n6939 GND.n6190 240.244
R16100 GND.n6939 GND.n6201 240.244
R16101 GND.n6949 GND.n6201 240.244
R16102 GND.n6949 GND.n6211 240.244
R16103 GND.n6954 GND.n6211 240.244
R16104 GND.n6954 GND.n6222 240.244
R16105 GND.n6964 GND.n6222 240.244
R16106 GND.n6964 GND.n6232 240.244
R16107 GND.n6969 GND.n6232 240.244
R16108 GND.n6969 GND.n6242 240.244
R16109 GND.n6986 GND.n6242 240.244
R16110 GND.n6986 GND.n6252 240.244
R16111 GND.n6257 GND.n6252 240.244
R16112 GND.n6993 GND.n6257 240.244
R16113 GND.n6994 GND.n6993 240.244
R16114 GND.n6994 GND.n93 240.244
R16115 GND.n7002 GND.n93 240.244
R16116 GND.n7002 GND.n6466 240.244
R16117 GND.n6466 GND.n6270 240.244
R16118 GND.n6270 GND.n112 240.244
R16119 GND.n6278 GND.n112 240.244
R16120 GND.n6278 GND.n123 240.244
R16121 GND.n7016 GND.n123 240.244
R16122 GND.n7016 GND.n133 240.244
R16123 GND.n7026 GND.n133 240.244
R16124 GND.n7026 GND.n143 240.244
R16125 GND.n7031 GND.n143 240.244
R16126 GND.n7031 GND.n154 240.244
R16127 GND.n7041 GND.n154 240.244
R16128 GND.n7041 GND.n164 240.244
R16129 GND.n7046 GND.n164 240.244
R16130 GND.n7046 GND.n175 240.244
R16131 GND.n7056 GND.n175 240.244
R16132 GND.n7056 GND.n185 240.244
R16133 GND.n7061 GND.n185 240.244
R16134 GND.n7061 GND.n196 240.244
R16135 GND.n7071 GND.n196 240.244
R16136 GND.n7071 GND.n206 240.244
R16137 GND.n7076 GND.n206 240.244
R16138 GND.n7076 GND.n217 240.244
R16139 GND.n7086 GND.n217 240.244
R16140 GND.n7086 GND.n227 240.244
R16141 GND.n7091 GND.n227 240.244
R16142 GND.n7091 GND.n238 240.244
R16143 GND.n7102 GND.n238 240.244
R16144 GND.n7102 GND.n248 240.244
R16145 GND.n6434 GND.n248 240.244
R16146 GND.n6434 GND.n258 240.244
R16147 GND.n7261 GND.n258 240.244
R16148 GND.n7261 GND.n268 240.244
R16149 GND.n7257 GND.n268 240.244
R16150 GND.n7257 GND.n279 240.244
R16151 GND.n7249 GND.n279 240.244
R16152 GND.n7249 GND.n289 240.244
R16153 GND.n7245 GND.n289 240.244
R16154 GND.n7245 GND.n300 240.244
R16155 GND.n7237 GND.n300 240.244
R16156 GND.n7237 GND.n310 240.244
R16157 GND.n7233 GND.n310 240.244
R16158 GND.n7233 GND.n321 240.244
R16159 GND.n7225 GND.n321 240.244
R16160 GND.n7225 GND.n331 240.244
R16161 GND.n7221 GND.n331 240.244
R16162 GND.n7221 GND.n342 240.244
R16163 GND.n7213 GND.n342 240.244
R16164 GND.n7213 GND.n352 240.244
R16165 GND.n7209 GND.n352 240.244
R16166 GND.n7209 GND.n363 240.244
R16167 GND.n7201 GND.n363 240.244
R16168 GND.n7201 GND.n373 240.244
R16169 GND.n7197 GND.n373 240.244
R16170 GND.n7197 GND.n384 240.244
R16171 GND.n7189 GND.n384 240.244
R16172 GND.n7189 GND.n394 240.244
R16173 GND.n7185 GND.n394 240.244
R16174 GND.n7185 GND.n405 240.244
R16175 GND.n7177 GND.n405 240.244
R16176 GND.n7177 GND.n415 240.244
R16177 GND.n7173 GND.n415 240.244
R16178 GND.n7173 GND.n426 240.244
R16179 GND.n7165 GND.n426 240.244
R16180 GND.n7165 GND.n436 240.244
R16181 GND.n10906 GND.n436 240.244
R16182 GND.n10906 GND.n446 240.244
R16183 GND.n4604 GND.n4603 240.244
R16184 GND.n7640 GND.n4603 240.244
R16185 GND.n7638 GND.n7637 240.244
R16186 GND.n7634 GND.n7633 240.244
R16187 GND.n7630 GND.n7629 240.244
R16188 GND.n7626 GND.n7625 240.244
R16189 GND.n7621 GND.n4618 240.244
R16190 GND.n7619 GND.n7618 240.244
R16191 GND.n7615 GND.n7614 240.244
R16192 GND.n7611 GND.n7610 240.244
R16193 GND.n7607 GND.n7606 240.244
R16194 GND.n7603 GND.n7602 240.244
R16195 GND.n7599 GND.n7598 240.244
R16196 GND.n7595 GND.n4792 240.244
R16197 GND.n7593 GND.n7592 240.244
R16198 GND.n7589 GND.n7588 240.244
R16199 GND.n7585 GND.n7584 240.244
R16200 GND.n7581 GND.n7580 240.244
R16201 GND.n7577 GND.n7576 240.244
R16202 GND.n7573 GND.n7572 240.244
R16203 GND.n7569 GND.n7568 240.244
R16204 GND.n7565 GND.n7564 240.244
R16205 GND.n7561 GND.n7560 240.244
R16206 GND.n7557 GND.n7556 240.244
R16207 GND.n7553 GND.n7552 240.244
R16208 GND.n7549 GND.n7548 240.244
R16209 GND.n7545 GND.n7544 240.244
R16210 GND.n7541 GND.n7540 240.244
R16211 GND.n7528 GND.n4605 240.244
R16212 GND.n7528 GND.n5921 240.244
R16213 GND.n7524 GND.n5921 240.244
R16214 GND.n7524 GND.n5928 240.244
R16215 GND.n7516 GND.n5928 240.244
R16216 GND.n7516 GND.n5944 240.244
R16217 GND.n7512 GND.n5944 240.244
R16218 GND.n7512 GND.n5950 240.244
R16219 GND.n7504 GND.n5950 240.244
R16220 GND.n7504 GND.n5964 240.244
R16221 GND.n7500 GND.n5964 240.244
R16222 GND.n7500 GND.n5970 240.244
R16223 GND.n7492 GND.n5970 240.244
R16224 GND.n7492 GND.n5985 240.244
R16225 GND.n7488 GND.n5985 240.244
R16226 GND.n7488 GND.n5991 240.244
R16227 GND.n7480 GND.n5991 240.244
R16228 GND.n7480 GND.n6006 240.244
R16229 GND.n7476 GND.n6006 240.244
R16230 GND.n7476 GND.n6012 240.244
R16231 GND.n7468 GND.n6012 240.244
R16232 GND.n7468 GND.n6027 240.244
R16233 GND.n7464 GND.n6027 240.244
R16234 GND.n7464 GND.n6033 240.244
R16235 GND.n7456 GND.n6033 240.244
R16236 GND.n7456 GND.n6047 240.244
R16237 GND.n7452 GND.n6047 240.244
R16238 GND.n7452 GND.n6053 240.244
R16239 GND.n7444 GND.n6053 240.244
R16240 GND.n7444 GND.n6068 240.244
R16241 GND.n7440 GND.n6068 240.244
R16242 GND.n7440 GND.n6074 240.244
R16243 GND.n7432 GND.n6074 240.244
R16244 GND.n7432 GND.n6089 240.244
R16245 GND.n7428 GND.n6089 240.244
R16246 GND.n7428 GND.n6095 240.244
R16247 GND.n7420 GND.n6095 240.244
R16248 GND.n7420 GND.n6110 240.244
R16249 GND.n7416 GND.n6110 240.244
R16250 GND.n7416 GND.n6116 240.244
R16251 GND.n7408 GND.n6116 240.244
R16252 GND.n7408 GND.n6131 240.244
R16253 GND.n7404 GND.n6131 240.244
R16254 GND.n7404 GND.n6137 240.244
R16255 GND.n7396 GND.n6137 240.244
R16256 GND.n7396 GND.n6152 240.244
R16257 GND.n7392 GND.n6152 240.244
R16258 GND.n7392 GND.n6158 240.244
R16259 GND.n7384 GND.n6158 240.244
R16260 GND.n7384 GND.n6172 240.244
R16261 GND.n7380 GND.n6172 240.244
R16262 GND.n7380 GND.n6178 240.244
R16263 GND.n7372 GND.n6178 240.244
R16264 GND.n7372 GND.n6193 240.244
R16265 GND.n7368 GND.n6193 240.244
R16266 GND.n7368 GND.n6199 240.244
R16267 GND.n7360 GND.n6199 240.244
R16268 GND.n7360 GND.n6214 240.244
R16269 GND.n7356 GND.n6214 240.244
R16270 GND.n7356 GND.n6220 240.244
R16271 GND.n7348 GND.n6220 240.244
R16272 GND.n7348 GND.n6235 240.244
R16273 GND.n7344 GND.n6235 240.244
R16274 GND.n7344 GND.n6240 240.244
R16275 GND.n7336 GND.n6240 240.244
R16276 GND.n7336 GND.n7334 240.244
R16277 GND.n7334 GND.n6256 240.244
R16278 GND.n6256 GND.n96 240.244
R16279 GND.n11110 GND.n96 240.244
R16280 GND.n11110 GND.n97 240.244
R16281 GND.n6268 GND.n97 240.244
R16282 GND.n6268 GND.n109 240.244
R16283 GND.n11105 GND.n109 240.244
R16284 GND.n11105 GND.n110 240.244
R16285 GND.n11097 GND.n110 240.244
R16286 GND.n11097 GND.n126 240.244
R16287 GND.n11093 GND.n126 240.244
R16288 GND.n11093 GND.n131 240.244
R16289 GND.n11085 GND.n131 240.244
R16290 GND.n11085 GND.n146 240.244
R16291 GND.n11081 GND.n146 240.244
R16292 GND.n11081 GND.n152 240.244
R16293 GND.n11073 GND.n152 240.244
R16294 GND.n11073 GND.n167 240.244
R16295 GND.n11069 GND.n167 240.244
R16296 GND.n11069 GND.n173 240.244
R16297 GND.n11061 GND.n173 240.244
R16298 GND.n11061 GND.n188 240.244
R16299 GND.n11057 GND.n188 240.244
R16300 GND.n11057 GND.n194 240.244
R16301 GND.n11049 GND.n194 240.244
R16302 GND.n11049 GND.n209 240.244
R16303 GND.n11045 GND.n209 240.244
R16304 GND.n11045 GND.n215 240.244
R16305 GND.n11037 GND.n215 240.244
R16306 GND.n11037 GND.n230 240.244
R16307 GND.n11033 GND.n230 240.244
R16308 GND.n11033 GND.n236 240.244
R16309 GND.n11025 GND.n236 240.244
R16310 GND.n11025 GND.n251 240.244
R16311 GND.n11021 GND.n251 240.244
R16312 GND.n11021 GND.n257 240.244
R16313 GND.n11013 GND.n257 240.244
R16314 GND.n11013 GND.n271 240.244
R16315 GND.n11009 GND.n271 240.244
R16316 GND.n11009 GND.n277 240.244
R16317 GND.n11001 GND.n277 240.244
R16318 GND.n11001 GND.n292 240.244
R16319 GND.n10997 GND.n292 240.244
R16320 GND.n10997 GND.n298 240.244
R16321 GND.n10989 GND.n298 240.244
R16322 GND.n10989 GND.n313 240.244
R16323 GND.n10985 GND.n313 240.244
R16324 GND.n10985 GND.n319 240.244
R16325 GND.n10977 GND.n319 240.244
R16326 GND.n10977 GND.n334 240.244
R16327 GND.n10973 GND.n334 240.244
R16328 GND.n10973 GND.n340 240.244
R16329 GND.n10965 GND.n340 240.244
R16330 GND.n10965 GND.n355 240.244
R16331 GND.n10961 GND.n355 240.244
R16332 GND.n10961 GND.n361 240.244
R16333 GND.n10953 GND.n361 240.244
R16334 GND.n10953 GND.n376 240.244
R16335 GND.n10949 GND.n376 240.244
R16336 GND.n10949 GND.n382 240.244
R16337 GND.n10941 GND.n382 240.244
R16338 GND.n10941 GND.n397 240.244
R16339 GND.n10937 GND.n397 240.244
R16340 GND.n10937 GND.n403 240.244
R16341 GND.n10929 GND.n403 240.244
R16342 GND.n10929 GND.n418 240.244
R16343 GND.n10925 GND.n418 240.244
R16344 GND.n10925 GND.n424 240.244
R16345 GND.n10917 GND.n424 240.244
R16346 GND.n10917 GND.n439 240.244
R16347 GND.n10913 GND.n439 240.244
R16348 GND.n2210 GND.n2209 240.244
R16349 GND.n8317 GND.n8316 240.244
R16350 GND.n2206 GND.n2205 240.244
R16351 GND.n8325 GND.n8324 240.244
R16352 GND.n2202 GND.n2201 240.244
R16353 GND.n8335 GND.n8334 240.244
R16354 GND.n2198 GND.n2197 240.244
R16355 GND.n8343 GND.n8342 240.244
R16356 GND.n2194 GND.n2193 240.244
R16357 GND.n8351 GND.n8350 240.244
R16358 GND.n2190 GND.n2189 240.244
R16359 GND.n8359 GND.n8358 240.244
R16360 GND.n8456 GND.n8455 240.244
R16361 GND.n8365 GND.n8364 240.244
R16362 GND.n8367 GND.n8366 240.244
R16363 GND.n8371 GND.n8370 240.244
R16364 GND.n8373 GND.n8372 240.244
R16365 GND.n8377 GND.n8376 240.244
R16366 GND.n8379 GND.n8378 240.244
R16367 GND.n8386 GND.n8385 240.244
R16368 GND.n8388 GND.n8387 240.244
R16369 GND.n8392 GND.n8391 240.244
R16370 GND.n8394 GND.n8393 240.244
R16371 GND.n8398 GND.n8397 240.244
R16372 GND.n8400 GND.n8399 240.244
R16373 GND.n8404 GND.n8403 240.244
R16374 GND.n8409 GND.n8405 240.244
R16375 GND.n1850 GND.n1803 240.244
R16376 GND.n1850 GND.n1849 240.244
R16377 GND.n1849 GND.n1818 240.244
R16378 GND.n2906 GND.n1818 240.244
R16379 GND.n2906 GND.n1837 240.244
R16380 GND.n1860 GND.n1837 240.244
R16381 GND.n1861 GND.n1860 240.244
R16382 GND.n3151 GND.n1861 240.244
R16383 GND.n3151 GND.n1867 240.244
R16384 GND.n1868 GND.n1867 240.244
R16385 GND.n1869 GND.n1868 240.244
R16386 GND.n2887 GND.n1869 240.244
R16387 GND.n2887 GND.n1875 240.244
R16388 GND.n1876 GND.n1875 240.244
R16389 GND.n1877 GND.n1876 240.244
R16390 GND.n3196 GND.n1877 240.244
R16391 GND.n3196 GND.n1883 240.244
R16392 GND.n1884 GND.n1883 240.244
R16393 GND.n1885 GND.n1884 240.244
R16394 GND.n2852 GND.n1885 240.244
R16395 GND.n2852 GND.n1891 240.244
R16396 GND.n1892 GND.n1891 240.244
R16397 GND.n1893 GND.n1892 240.244
R16398 GND.n2833 GND.n1893 240.244
R16399 GND.n2833 GND.n1899 240.244
R16400 GND.n1900 GND.n1899 240.244
R16401 GND.n1901 GND.n1900 240.244
R16402 GND.n2821 GND.n1901 240.244
R16403 GND.n2821 GND.n1907 240.244
R16404 GND.n1908 GND.n1907 240.244
R16405 GND.n1909 GND.n1908 240.244
R16406 GND.n2796 GND.n1909 240.244
R16407 GND.n2796 GND.n1915 240.244
R16408 GND.n1916 GND.n1915 240.244
R16409 GND.n1917 GND.n1916 240.244
R16410 GND.n3295 GND.n1917 240.244
R16411 GND.n3295 GND.n1923 240.244
R16412 GND.n1924 GND.n1923 240.244
R16413 GND.n1925 GND.n1924 240.244
R16414 GND.n2761 GND.n1925 240.244
R16415 GND.n2761 GND.n1931 240.244
R16416 GND.n1932 GND.n1931 240.244
R16417 GND.n1933 GND.n1932 240.244
R16418 GND.n2742 GND.n1933 240.244
R16419 GND.n2742 GND.n1939 240.244
R16420 GND.n1940 GND.n1939 240.244
R16421 GND.n1941 GND.n1940 240.244
R16422 GND.n2730 GND.n1941 240.244
R16423 GND.n2730 GND.n1947 240.244
R16424 GND.n1948 GND.n1947 240.244
R16425 GND.n1949 GND.n1948 240.244
R16426 GND.n2705 GND.n1949 240.244
R16427 GND.n2705 GND.n1955 240.244
R16428 GND.n1956 GND.n1955 240.244
R16429 GND.n1957 GND.n1956 240.244
R16430 GND.n3394 GND.n1957 240.244
R16431 GND.n3394 GND.n1963 240.244
R16432 GND.n1964 GND.n1963 240.244
R16433 GND.n1965 GND.n1964 240.244
R16434 GND.n2670 GND.n1965 240.244
R16435 GND.n2670 GND.n1971 240.244
R16436 GND.n1972 GND.n1971 240.244
R16437 GND.n1973 GND.n1972 240.244
R16438 GND.n2502 GND.n1973 240.244
R16439 GND.n2502 GND.n1979 240.244
R16440 GND.n1980 GND.n1979 240.244
R16441 GND.n1981 GND.n1980 240.244
R16442 GND.n2517 GND.n1981 240.244
R16443 GND.n2517 GND.n1987 240.244
R16444 GND.n1988 GND.n1987 240.244
R16445 GND.n1989 GND.n1988 240.244
R16446 GND.n2650 GND.n1989 240.244
R16447 GND.n2650 GND.n1995 240.244
R16448 GND.n1996 GND.n1995 240.244
R16449 GND.n1997 GND.n1996 240.244
R16450 GND.n2477 GND.n1997 240.244
R16451 GND.n2477 GND.n2003 240.244
R16452 GND.n2004 GND.n2003 240.244
R16453 GND.n2005 GND.n2004 240.244
R16454 GND.n2465 GND.n2005 240.244
R16455 GND.n2465 GND.n2011 240.244
R16456 GND.n2012 GND.n2011 240.244
R16457 GND.n2013 GND.n2012 240.244
R16458 GND.n2441 GND.n2013 240.244
R16459 GND.n2441 GND.n2019 240.244
R16460 GND.n2020 GND.n2019 240.244
R16461 GND.n2021 GND.n2020 240.244
R16462 GND.n3564 GND.n2021 240.244
R16463 GND.n3564 GND.n2027 240.244
R16464 GND.n2028 GND.n2027 240.244
R16465 GND.n2029 GND.n2028 240.244
R16466 GND.n2408 GND.n2029 240.244
R16467 GND.n2408 GND.n2035 240.244
R16468 GND.n2036 GND.n2035 240.244
R16469 GND.n2037 GND.n2036 240.244
R16470 GND.n2390 GND.n2037 240.244
R16471 GND.n2390 GND.n2043 240.244
R16472 GND.n2044 GND.n2043 240.244
R16473 GND.n2045 GND.n2044 240.244
R16474 GND.n2604 GND.n2045 240.244
R16475 GND.n2604 GND.n2051 240.244
R16476 GND.n2052 GND.n2051 240.244
R16477 GND.n2053 GND.n2052 240.244
R16478 GND.n2357 GND.n2053 240.244
R16479 GND.n2357 GND.n2059 240.244
R16480 GND.n2060 GND.n2059 240.244
R16481 GND.n2061 GND.n2060 240.244
R16482 GND.n3667 GND.n2061 240.244
R16483 GND.n3667 GND.n2067 240.244
R16484 GND.n2068 GND.n2067 240.244
R16485 GND.n2069 GND.n2068 240.244
R16486 GND.n2318 GND.n2069 240.244
R16487 GND.n2318 GND.n2075 240.244
R16488 GND.n2076 GND.n2075 240.244
R16489 GND.n2077 GND.n2076 240.244
R16490 GND.n2301 GND.n2077 240.244
R16491 GND.n2301 GND.n2083 240.244
R16492 GND.n2084 GND.n2083 240.244
R16493 GND.n2085 GND.n2084 240.244
R16494 GND.n2289 GND.n2085 240.244
R16495 GND.n2289 GND.n2091 240.244
R16496 GND.n2092 GND.n2091 240.244
R16497 GND.n2093 GND.n2092 240.244
R16498 GND.n2265 GND.n2093 240.244
R16499 GND.n2265 GND.n2099 240.244
R16500 GND.n2100 GND.n2099 240.244
R16501 GND.n2101 GND.n2100 240.244
R16502 GND.n8256 GND.n2101 240.244
R16503 GND.n8256 GND.n2107 240.244
R16504 GND.n2108 GND.n2107 240.244
R16505 GND.n2109 GND.n2108 240.244
R16506 GND.n2232 GND.n2109 240.244
R16507 GND.n2232 GND.n2115 240.244
R16508 GND.n2116 GND.n2115 240.244
R16509 GND.n2117 GND.n2116 240.244
R16510 GND.n2123 GND.n2117 240.244
R16511 GND.n8481 GND.n2123 240.244
R16512 GND.n1727 GND.n1726 240.244
R16513 GND.n8809 GND.n1726 240.244
R16514 GND.n8807 GND.n8806 240.244
R16515 GND.n8803 GND.n8802 240.244
R16516 GND.n8799 GND.n8798 240.244
R16517 GND.n8795 GND.n8794 240.244
R16518 GND.n8790 GND.n1741 240.244
R16519 GND.n8788 GND.n8787 240.244
R16520 GND.n8784 GND.n8783 240.244
R16521 GND.n8780 GND.n8779 240.244
R16522 GND.n8776 GND.n8775 240.244
R16523 GND.n8772 GND.n8771 240.244
R16524 GND.n8768 GND.n8767 240.244
R16525 GND.n8764 GND.n8763 240.244
R16526 GND.n8760 GND.n8759 240.244
R16527 GND.n8756 GND.n8755 240.244
R16528 GND.n8752 GND.n8751 240.244
R16529 GND.n8748 GND.n8747 240.244
R16530 GND.n8744 GND.n8743 240.244
R16531 GND.n8740 GND.n8739 240.244
R16532 GND.n8736 GND.n8735 240.244
R16533 GND.n8732 GND.n8731 240.244
R16534 GND.n8728 GND.n8727 240.244
R16535 GND.n8724 GND.n8723 240.244
R16536 GND.n8720 GND.n8719 240.244
R16537 GND.n8716 GND.n8715 240.244
R16538 GND.n8712 GND.n8711 240.244
R16539 GND.n8708 GND.n8707 240.244
R16540 GND.n1827 GND.n1728 240.244
R16541 GND.n1827 GND.n1822 240.244
R16542 GND.n8689 GND.n1822 240.244
R16543 GND.n8689 GND.n1823 240.244
R16544 GND.n8685 GND.n1823 240.244
R16545 GND.n8685 GND.n1835 240.244
R16546 GND.n3159 GND.n1835 240.244
R16547 GND.n3159 GND.n3153 240.244
R16548 GND.n3153 GND.n2896 240.244
R16549 GND.n3176 GND.n2896 240.244
R16550 GND.n3176 GND.n2890 240.244
R16551 GND.n3184 GND.n2890 240.244
R16552 GND.n3184 GND.n2892 240.244
R16553 GND.n2892 GND.n2873 240.244
R16554 GND.n3201 GND.n2873 240.244
R16555 GND.n3201 GND.n2867 240.244
R16556 GND.n3209 GND.n2867 240.244
R16557 GND.n3209 GND.n2869 240.244
R16558 GND.n2869 GND.n2850 240.244
R16559 GND.n3225 GND.n2850 240.244
R16560 GND.n3225 GND.n2844 240.244
R16561 GND.n3233 GND.n2844 240.244
R16562 GND.n3233 GND.n2846 240.244
R16563 GND.n2846 GND.n2827 240.244
R16564 GND.n3250 GND.n2827 240.244
R16565 GND.n3250 GND.n2820 240.244
R16566 GND.n3258 GND.n2820 240.244
R16567 GND.n3258 GND.n2823 240.244
R16568 GND.n2823 GND.n2805 240.244
R16569 GND.n3275 GND.n2805 240.244
R16570 GND.n3275 GND.n2799 240.244
R16571 GND.n3283 GND.n2799 240.244
R16572 GND.n3283 GND.n2801 240.244
R16573 GND.n2801 GND.n2782 240.244
R16574 GND.n3300 GND.n2782 240.244
R16575 GND.n3300 GND.n2776 240.244
R16576 GND.n3308 GND.n2776 240.244
R16577 GND.n3308 GND.n2778 240.244
R16578 GND.n2778 GND.n2759 240.244
R16579 GND.n3324 GND.n2759 240.244
R16580 GND.n3324 GND.n2753 240.244
R16581 GND.n3332 GND.n2753 240.244
R16582 GND.n3332 GND.n2755 240.244
R16583 GND.n2755 GND.n2736 240.244
R16584 GND.n3349 GND.n2736 240.244
R16585 GND.n3349 GND.n2729 240.244
R16586 GND.n3357 GND.n2729 240.244
R16587 GND.n3357 GND.n2732 240.244
R16588 GND.n2732 GND.n2714 240.244
R16589 GND.n3374 GND.n2714 240.244
R16590 GND.n3374 GND.n2708 240.244
R16591 GND.n3382 GND.n2708 240.244
R16592 GND.n3382 GND.n2710 240.244
R16593 GND.n2710 GND.n2691 240.244
R16594 GND.n3399 GND.n2691 240.244
R16595 GND.n3399 GND.n2685 240.244
R16596 GND.n3407 GND.n2685 240.244
R16597 GND.n3407 GND.n2687 240.244
R16598 GND.n2687 GND.n2668 240.244
R16599 GND.n3423 GND.n2668 240.244
R16600 GND.n3423 GND.n2664 240.244
R16601 GND.n3429 GND.n2664 240.244
R16602 GND.n3429 GND.n2499 240.244
R16603 GND.n3491 GND.n2499 240.244
R16604 GND.n3491 GND.n2500 240.244
R16605 GND.n2522 GND.n2500 240.244
R16606 GND.n2524 GND.n2522 240.244
R16607 GND.n3477 GND.n2524 240.244
R16608 GND.n3477 GND.n3474 240.244
R16609 GND.n3474 GND.n2525 240.244
R16610 GND.n3455 GND.n2525 240.244
R16611 GND.n3457 GND.n3455 240.244
R16612 GND.n3457 GND.n2487 240.244
R16613 GND.n3499 GND.n2487 240.244
R16614 GND.n3499 GND.n2489 240.244
R16615 GND.n2489 GND.n2471 240.244
R16616 GND.n3517 GND.n2471 240.244
R16617 GND.n3517 GND.n2464 240.244
R16618 GND.n3525 GND.n2464 240.244
R16619 GND.n3525 GND.n2467 240.244
R16620 GND.n2467 GND.n2450 240.244
R16621 GND.n3543 GND.n2450 240.244
R16622 GND.n3543 GND.n2444 240.244
R16623 GND.n3551 GND.n2444 240.244
R16624 GND.n3551 GND.n2446 240.244
R16625 GND.n2446 GND.n2428 240.244
R16626 GND.n3569 GND.n2428 240.244
R16627 GND.n3569 GND.n2422 240.244
R16628 GND.n3577 GND.n2422 240.244
R16629 GND.n3577 GND.n2424 240.244
R16630 GND.n2424 GND.n2406 240.244
R16631 GND.n3594 GND.n2406 240.244
R16632 GND.n3594 GND.n2400 240.244
R16633 GND.n3602 GND.n2400 240.244
R16634 GND.n3602 GND.n2402 240.244
R16635 GND.n2402 GND.n2384 240.244
R16636 GND.n3620 GND.n2384 240.244
R16637 GND.n3620 GND.n2379 240.244
R16638 GND.n3628 GND.n2379 240.244
R16639 GND.n3628 GND.n2380 240.244
R16640 GND.n2380 GND.n2366 240.244
R16641 GND.n3646 GND.n2366 240.244
R16642 GND.n3646 GND.n2360 240.244
R16643 GND.n3654 GND.n2360 240.244
R16644 GND.n3654 GND.n2362 240.244
R16645 GND.n2362 GND.n2344 240.244
R16646 GND.n3672 GND.n2344 240.244
R16647 GND.n3672 GND.n2339 240.244
R16648 GND.n3680 GND.n2339 240.244
R16649 GND.n3680 GND.n2340 240.244
R16650 GND.n2340 GND.n2316 240.244
R16651 GND.n8183 GND.n2316 240.244
R16652 GND.n8183 GND.n2310 240.244
R16653 GND.n8191 GND.n2310 240.244
R16654 GND.n8191 GND.n2312 240.244
R16655 GND.n2312 GND.n2295 240.244
R16656 GND.n8209 GND.n2295 240.244
R16657 GND.n8209 GND.n2288 240.244
R16658 GND.n8217 GND.n2288 240.244
R16659 GND.n8217 GND.n2291 240.244
R16660 GND.n2291 GND.n2274 240.244
R16661 GND.n8235 GND.n2274 240.244
R16662 GND.n8235 GND.n2268 240.244
R16663 GND.n8243 GND.n2268 240.244
R16664 GND.n8243 GND.n2270 240.244
R16665 GND.n2270 GND.n2252 240.244
R16666 GND.n8261 GND.n2252 240.244
R16667 GND.n8261 GND.n2246 240.244
R16668 GND.n8269 GND.n2246 240.244
R16669 GND.n8269 GND.n2248 240.244
R16670 GND.n2248 GND.n2230 240.244
R16671 GND.n8286 GND.n2230 240.244
R16672 GND.n8286 GND.n2226 240.244
R16673 GND.n8293 GND.n2226 240.244
R16674 GND.n8293 GND.n2213 240.244
R16675 GND.n8305 GND.n2213 240.244
R16676 GND.n8305 GND.n2126 240.244
R16677 GND.n5818 GND.n5816 240.244
R16678 GND.n5825 GND.n4847 240.244
R16679 GND.n5828 GND.n5827 240.244
R16680 GND.n5833 GND.n5831 240.244
R16681 GND.n5837 GND.n5835 240.244
R16682 GND.n5842 GND.n5839 240.244
R16683 GND.n5847 GND.n5844 240.244
R16684 GND.n5852 GND.n5849 240.244
R16685 GND.n5857 GND.n5854 240.244
R16686 GND.n5865 GND.n5859 240.244
R16687 GND.n5870 GND.n5867 240.244
R16688 GND.n8006 GND.n3879 240.244
R16689 GND.n7998 GND.n3879 240.244
R16690 GND.n7998 GND.n3896 240.244
R16691 GND.n7994 GND.n3896 240.244
R16692 GND.n7994 GND.n3904 240.244
R16693 GND.n7986 GND.n3904 240.244
R16694 GND.n7986 GND.n3917 240.244
R16695 GND.n7982 GND.n3917 240.244
R16696 GND.n7982 GND.n3923 240.244
R16697 GND.n7974 GND.n3923 240.244
R16698 GND.n7974 GND.n3937 240.244
R16699 GND.n7970 GND.n3937 240.244
R16700 GND.n7970 GND.n3943 240.244
R16701 GND.n7962 GND.n3943 240.244
R16702 GND.n7962 GND.n3957 240.244
R16703 GND.n7958 GND.n3957 240.244
R16704 GND.n7958 GND.n3963 240.244
R16705 GND.n7950 GND.n3963 240.244
R16706 GND.n7950 GND.n3977 240.244
R16707 GND.n7946 GND.n3977 240.244
R16708 GND.n7946 GND.n3983 240.244
R16709 GND.n7938 GND.n3983 240.244
R16710 GND.n7938 GND.n3997 240.244
R16711 GND.n7934 GND.n3997 240.244
R16712 GND.n7934 GND.n4003 240.244
R16713 GND.n7926 GND.n4003 240.244
R16714 GND.n7926 GND.n4017 240.244
R16715 GND.n7922 GND.n4017 240.244
R16716 GND.n7922 GND.n4023 240.244
R16717 GND.n7914 GND.n4023 240.244
R16718 GND.n7914 GND.n4037 240.244
R16719 GND.n7910 GND.n4037 240.244
R16720 GND.n7910 GND.n4043 240.244
R16721 GND.n4058 GND.n4043 240.244
R16722 GND.n4098 GND.n4058 240.244
R16723 GND.n4099 GND.n4098 240.244
R16724 GND.n4099 GND.n4075 240.244
R16725 GND.n4089 GND.n4075 240.244
R16726 GND.n7883 GND.n4089 240.244
R16727 GND.n7883 GND.n4090 240.244
R16728 GND.n7879 GND.n4090 240.244
R16729 GND.n7879 GND.n4108 240.244
R16730 GND.n7871 GND.n4108 240.244
R16731 GND.n7871 GND.n4122 240.244
R16732 GND.n7867 GND.n4122 240.244
R16733 GND.n7867 GND.n4128 240.244
R16734 GND.n7859 GND.n4128 240.244
R16735 GND.n7859 GND.n4142 240.244
R16736 GND.n7855 GND.n4142 240.244
R16737 GND.n7855 GND.n4148 240.244
R16738 GND.n4163 GND.n4148 240.244
R16739 GND.n4202 GND.n4163 240.244
R16740 GND.n4203 GND.n4202 240.244
R16741 GND.n4203 GND.n4180 240.244
R16742 GND.n4193 GND.n4180 240.244
R16743 GND.n7828 GND.n4193 240.244
R16744 GND.n7828 GND.n4194 240.244
R16745 GND.n7824 GND.n4194 240.244
R16746 GND.n7824 GND.n4212 240.244
R16747 GND.n7816 GND.n4212 240.244
R16748 GND.n7816 GND.n4226 240.244
R16749 GND.n7812 GND.n4226 240.244
R16750 GND.n7812 GND.n4232 240.244
R16751 GND.n7804 GND.n4232 240.244
R16752 GND.n7804 GND.n4244 240.244
R16753 GND.n7800 GND.n4244 240.244
R16754 GND.n7800 GND.n4250 240.244
R16755 GND.n4265 GND.n4250 240.244
R16756 GND.n4305 GND.n4265 240.244
R16757 GND.n4306 GND.n4305 240.244
R16758 GND.n4306 GND.n4282 240.244
R16759 GND.n4296 GND.n4282 240.244
R16760 GND.n7773 GND.n4296 240.244
R16761 GND.n7773 GND.n4297 240.244
R16762 GND.n7769 GND.n4297 240.244
R16763 GND.n7769 GND.n4315 240.244
R16764 GND.n7761 GND.n4315 240.244
R16765 GND.n7761 GND.n4329 240.244
R16766 GND.n7757 GND.n4329 240.244
R16767 GND.n7757 GND.n4335 240.244
R16768 GND.n7749 GND.n4335 240.244
R16769 GND.n7749 GND.n4348 240.244
R16770 GND.n7745 GND.n4348 240.244
R16771 GND.n7745 GND.n4354 240.244
R16772 GND.n4369 GND.n4354 240.244
R16773 GND.n3863 GND.n3862 240.244
R16774 GND.n8049 GND.n3862 240.244
R16775 GND.n8047 GND.n8046 240.244
R16776 GND.n3872 GND.n3871 240.244
R16777 GND.n8039 GND.n8038 240.244
R16778 GND.n8034 GND.n8033 240.244
R16779 GND.n8029 GND.n8028 240.244
R16780 GND.n8024 GND.n8023 240.244
R16781 GND.n8019 GND.n8018 240.244
R16782 GND.n8012 GND.n8011 240.244
R16783 GND.n3878 GND.n3877 240.244
R16784 GND.n5025 GND.n3864 240.244
R16785 GND.n5025 GND.n3894 240.244
R16786 GND.n5325 GND.n3894 240.244
R16787 GND.n5325 GND.n3905 240.244
R16788 GND.n5331 GND.n3905 240.244
R16789 GND.n5331 GND.n3915 240.244
R16790 GND.n5344 GND.n3915 240.244
R16791 GND.n5344 GND.n3925 240.244
R16792 GND.n5350 GND.n3925 240.244
R16793 GND.n5350 GND.n3935 240.244
R16794 GND.n5363 GND.n3935 240.244
R16795 GND.n5363 GND.n3945 240.244
R16796 GND.n5410 GND.n3945 240.244
R16797 GND.n5410 GND.n3955 240.244
R16798 GND.n5406 GND.n3955 240.244
R16799 GND.n5406 GND.n3965 240.244
R16800 GND.n4992 GND.n3965 240.244
R16801 GND.n4992 GND.n3975 240.244
R16802 GND.n5401 GND.n3975 240.244
R16803 GND.n5401 GND.n3985 240.244
R16804 GND.n5398 GND.n3985 240.244
R16805 GND.n5398 GND.n3995 240.244
R16806 GND.n5394 GND.n3995 240.244
R16807 GND.n5394 GND.n4005 240.244
R16808 GND.n5391 GND.n4005 240.244
R16809 GND.n5391 GND.n4015 240.244
R16810 GND.n5388 GND.n4015 240.244
R16811 GND.n5388 GND.n4025 240.244
R16812 GND.n5385 GND.n4025 240.244
R16813 GND.n5385 GND.n4035 240.244
R16814 GND.n5505 GND.n4035 240.244
R16815 GND.n5505 GND.n4045 240.244
R16816 GND.n4954 GND.n4045 240.244
R16817 GND.n4954 GND.n4056 240.244
R16818 GND.n5513 GND.n4056 240.244
R16819 GND.n5514 GND.n5513 240.244
R16820 GND.n5514 GND.n4073 240.244
R16821 GND.n5541 GND.n4073 240.244
R16822 GND.n5541 GND.n4087 240.244
R16823 GND.n5537 GND.n4087 240.244
R16824 GND.n5537 GND.n4110 240.244
R16825 GND.n5534 GND.n4110 240.244
R16826 GND.n5534 GND.n4120 240.244
R16827 GND.n5531 GND.n4120 240.244
R16828 GND.n5531 GND.n4130 240.244
R16829 GND.n5528 GND.n4130 240.244
R16830 GND.n5528 GND.n4140 240.244
R16831 GND.n5608 GND.n4140 240.244
R16832 GND.n5608 GND.n4150 240.244
R16833 GND.n4923 GND.n4150 240.244
R16834 GND.n4923 GND.n4161 240.244
R16835 GND.n5616 GND.n4161 240.244
R16836 GND.n5617 GND.n5616 240.244
R16837 GND.n5617 GND.n4178 240.244
R16838 GND.n5645 GND.n4178 240.244
R16839 GND.n5645 GND.n4192 240.244
R16840 GND.n5641 GND.n4192 240.244
R16841 GND.n5641 GND.n4214 240.244
R16842 GND.n5638 GND.n4214 240.244
R16843 GND.n5638 GND.n4224 240.244
R16844 GND.n5635 GND.n4224 240.244
R16845 GND.n5635 GND.n4234 240.244
R16846 GND.n5632 GND.n4234 240.244
R16847 GND.n5632 GND.n4243 240.244
R16848 GND.n5711 GND.n4243 240.244
R16849 GND.n5711 GND.n4252 240.244
R16850 GND.n4889 GND.n4252 240.244
R16851 GND.n4889 GND.n4263 240.244
R16852 GND.n5719 GND.n4263 240.244
R16853 GND.n5720 GND.n5719 240.244
R16854 GND.n5720 GND.n4280 240.244
R16855 GND.n5742 GND.n4280 240.244
R16856 GND.n5742 GND.n4294 240.244
R16857 GND.n5738 GND.n4294 240.244
R16858 GND.n5738 GND.n4317 240.244
R16859 GND.n5735 GND.n4317 240.244
R16860 GND.n5735 GND.n4327 240.244
R16861 GND.n5732 GND.n4327 240.244
R16862 GND.n5732 GND.n4337 240.244
R16863 GND.n5802 GND.n4337 240.244
R16864 GND.n5802 GND.n4347 240.244
R16865 GND.n4867 GND.n4347 240.244
R16866 GND.n4867 GND.n4356 240.244
R16867 GND.n5810 GND.n4356 240.244
R16868 GND.n5810 GND.n4367 240.244
R16869 GND.n10686 GND.n10652 240.244
R16870 GND.n10680 GND.n10679 240.244
R16871 GND.n10676 GND.n10675 240.244
R16872 GND.n10672 GND.n10671 240.244
R16873 GND.n10668 GND.n10667 240.244
R16874 GND.n10664 GND.n459 240.244
R16875 GND.n5919 GND.n5880 240.244
R16876 GND.n6746 GND.n5919 240.244
R16877 GND.n6746 GND.n5931 240.244
R16878 GND.n6752 GND.n5931 240.244
R16879 GND.n6752 GND.n5942 240.244
R16880 GND.n6761 GND.n5942 240.244
R16881 GND.n6761 GND.n5953 240.244
R16882 GND.n6767 GND.n5953 240.244
R16883 GND.n6767 GND.n5962 240.244
R16884 GND.n6776 GND.n5962 240.244
R16885 GND.n6776 GND.n5973 240.244
R16886 GND.n6782 GND.n5973 240.244
R16887 GND.n6782 GND.n5983 240.244
R16888 GND.n6791 GND.n5983 240.244
R16889 GND.n6791 GND.n5994 240.244
R16890 GND.n6797 GND.n5994 240.244
R16891 GND.n6797 GND.n6004 240.244
R16892 GND.n6806 GND.n6004 240.244
R16893 GND.n6806 GND.n6015 240.244
R16894 GND.n6812 GND.n6015 240.244
R16895 GND.n6812 GND.n6025 240.244
R16896 GND.n6821 GND.n6025 240.244
R16897 GND.n6821 GND.n6036 240.244
R16898 GND.n6827 GND.n6036 240.244
R16899 GND.n6827 GND.n6045 240.244
R16900 GND.n6836 GND.n6045 240.244
R16901 GND.n6836 GND.n6056 240.244
R16902 GND.n6842 GND.n6056 240.244
R16903 GND.n6842 GND.n6066 240.244
R16904 GND.n6851 GND.n6066 240.244
R16905 GND.n6851 GND.n6077 240.244
R16906 GND.n6857 GND.n6077 240.244
R16907 GND.n6857 GND.n6087 240.244
R16908 GND.n6866 GND.n6087 240.244
R16909 GND.n6866 GND.n6098 240.244
R16910 GND.n6872 GND.n6098 240.244
R16911 GND.n6872 GND.n6108 240.244
R16912 GND.n6881 GND.n6108 240.244
R16913 GND.n6881 GND.n6119 240.244
R16914 GND.n6887 GND.n6119 240.244
R16915 GND.n6887 GND.n6129 240.244
R16916 GND.n6896 GND.n6129 240.244
R16917 GND.n6896 GND.n6140 240.244
R16918 GND.n6902 GND.n6140 240.244
R16919 GND.n6902 GND.n6150 240.244
R16920 GND.n6911 GND.n6150 240.244
R16921 GND.n6911 GND.n6161 240.244
R16922 GND.n6917 GND.n6161 240.244
R16923 GND.n6917 GND.n6171 240.244
R16924 GND.n6926 GND.n6171 240.244
R16925 GND.n6926 GND.n6181 240.244
R16926 GND.n6932 GND.n6181 240.244
R16927 GND.n6932 GND.n6191 240.244
R16928 GND.n6941 GND.n6191 240.244
R16929 GND.n6941 GND.n6202 240.244
R16930 GND.n6947 GND.n6202 240.244
R16931 GND.n6947 GND.n6212 240.244
R16932 GND.n6956 GND.n6212 240.244
R16933 GND.n6956 GND.n6223 240.244
R16934 GND.n6962 GND.n6223 240.244
R16935 GND.n6962 GND.n6233 240.244
R16936 GND.n6971 GND.n6233 240.244
R16937 GND.n6971 GND.n6243 240.244
R16938 GND.n6984 GND.n6243 240.244
R16939 GND.n6984 GND.n6253 240.244
R16940 GND.n6258 GND.n6253 240.244
R16941 GND.n6979 GND.n6258 240.244
R16942 GND.n6979 GND.n90 240.244
R16943 GND.n11112 GND.n90 240.244
R16944 GND.n11112 GND.n91 240.244
R16945 GND.n6271 GND.n91 240.244
R16946 GND.n7317 GND.n6271 240.244
R16947 GND.n7317 GND.n113 240.244
R16948 GND.n7313 GND.n113 240.244
R16949 GND.n7313 GND.n124 240.244
R16950 GND.n7018 GND.n124 240.244
R16951 GND.n7018 GND.n134 240.244
R16952 GND.n7024 GND.n134 240.244
R16953 GND.n7024 GND.n144 240.244
R16954 GND.n7033 GND.n144 240.244
R16955 GND.n7033 GND.n155 240.244
R16956 GND.n7039 GND.n155 240.244
R16957 GND.n7039 GND.n165 240.244
R16958 GND.n7048 GND.n165 240.244
R16959 GND.n7048 GND.n176 240.244
R16960 GND.n7054 GND.n176 240.244
R16961 GND.n7054 GND.n186 240.244
R16962 GND.n7063 GND.n186 240.244
R16963 GND.n7063 GND.n197 240.244
R16964 GND.n7069 GND.n197 240.244
R16965 GND.n7069 GND.n207 240.244
R16966 GND.n7078 GND.n207 240.244
R16967 GND.n7078 GND.n218 240.244
R16968 GND.n7084 GND.n218 240.244
R16969 GND.n7084 GND.n228 240.244
R16970 GND.n7093 GND.n228 240.244
R16971 GND.n7093 GND.n239 240.244
R16972 GND.n7100 GND.n239 240.244
R16973 GND.n7100 GND.n249 240.244
R16974 GND.n7267 GND.n249 240.244
R16975 GND.n7267 GND.n259 240.244
R16976 GND.n7263 GND.n259 240.244
R16977 GND.n7263 GND.n269 240.244
R16978 GND.n7255 GND.n269 240.244
R16979 GND.n7255 GND.n280 240.244
R16980 GND.n7251 GND.n280 240.244
R16981 GND.n7251 GND.n290 240.244
R16982 GND.n7243 GND.n290 240.244
R16983 GND.n7243 GND.n301 240.244
R16984 GND.n7239 GND.n301 240.244
R16985 GND.n7239 GND.n311 240.244
R16986 GND.n7231 GND.n311 240.244
R16987 GND.n7231 GND.n322 240.244
R16988 GND.n7227 GND.n322 240.244
R16989 GND.n7227 GND.n332 240.244
R16990 GND.n7219 GND.n332 240.244
R16991 GND.n7219 GND.n343 240.244
R16992 GND.n7215 GND.n343 240.244
R16993 GND.n7215 GND.n353 240.244
R16994 GND.n7207 GND.n353 240.244
R16995 GND.n7207 GND.n364 240.244
R16996 GND.n7203 GND.n364 240.244
R16997 GND.n7203 GND.n374 240.244
R16998 GND.n7195 GND.n374 240.244
R16999 GND.n7195 GND.n385 240.244
R17000 GND.n7191 GND.n385 240.244
R17001 GND.n7191 GND.n395 240.244
R17002 GND.n7183 GND.n395 240.244
R17003 GND.n7183 GND.n406 240.244
R17004 GND.n7179 GND.n406 240.244
R17005 GND.n7179 GND.n416 240.244
R17006 GND.n7171 GND.n416 240.244
R17007 GND.n7171 GND.n427 240.244
R17008 GND.n7167 GND.n427 240.244
R17009 GND.n7167 GND.n437 240.244
R17010 GND.n10904 GND.n437 240.244
R17011 GND.n10904 GND.n447 240.244
R17012 GND.n5913 GND.n5912 240.244
R17013 GND.n5908 GND.n5907 240.244
R17014 GND.n5903 GND.n5902 240.244
R17015 GND.n5898 GND.n5897 240.244
R17016 GND.n5893 GND.n5892 240.244
R17017 GND.n5885 GND.n5882 240.244
R17018 GND.n7531 GND.n7530 240.244
R17019 GND.n7530 GND.n5917 240.244
R17020 GND.n7522 GND.n5917 240.244
R17021 GND.n7522 GND.n5933 240.244
R17022 GND.n7518 GND.n5933 240.244
R17023 GND.n7518 GND.n5939 240.244
R17024 GND.n7510 GND.n5939 240.244
R17025 GND.n7510 GND.n5954 240.244
R17026 GND.n7506 GND.n5954 240.244
R17027 GND.n7506 GND.n5959 240.244
R17028 GND.n7498 GND.n5959 240.244
R17029 GND.n7498 GND.n5975 240.244
R17030 GND.n7494 GND.n5975 240.244
R17031 GND.n7494 GND.n5980 240.244
R17032 GND.n7486 GND.n5980 240.244
R17033 GND.n7486 GND.n5996 240.244
R17034 GND.n7482 GND.n5996 240.244
R17035 GND.n7482 GND.n6001 240.244
R17036 GND.n7474 GND.n6001 240.244
R17037 GND.n7474 GND.n6017 240.244
R17038 GND.n7470 GND.n6017 240.244
R17039 GND.n7470 GND.n6022 240.244
R17040 GND.n7462 GND.n6022 240.244
R17041 GND.n7462 GND.n6037 240.244
R17042 GND.n7458 GND.n6037 240.244
R17043 GND.n7458 GND.n6042 240.244
R17044 GND.n7450 GND.n6042 240.244
R17045 GND.n7450 GND.n6058 240.244
R17046 GND.n7446 GND.n6058 240.244
R17047 GND.n7446 GND.n6063 240.244
R17048 GND.n7438 GND.n6063 240.244
R17049 GND.n7438 GND.n6079 240.244
R17050 GND.n7434 GND.n6079 240.244
R17051 GND.n7434 GND.n6084 240.244
R17052 GND.n7426 GND.n6084 240.244
R17053 GND.n7426 GND.n6100 240.244
R17054 GND.n7422 GND.n6100 240.244
R17055 GND.n7422 GND.n6105 240.244
R17056 GND.n7414 GND.n6105 240.244
R17057 GND.n7414 GND.n6121 240.244
R17058 GND.n7410 GND.n6121 240.244
R17059 GND.n7410 GND.n6126 240.244
R17060 GND.n7402 GND.n6126 240.244
R17061 GND.n7402 GND.n6142 240.244
R17062 GND.n7398 GND.n6142 240.244
R17063 GND.n7398 GND.n6147 240.244
R17064 GND.n7390 GND.n6147 240.244
R17065 GND.n7390 GND.n6163 240.244
R17066 GND.n7386 GND.n6163 240.244
R17067 GND.n7386 GND.n6168 240.244
R17068 GND.n7378 GND.n6168 240.244
R17069 GND.n7378 GND.n6183 240.244
R17070 GND.n7374 GND.n6183 240.244
R17071 GND.n7374 GND.n6188 240.244
R17072 GND.n7366 GND.n6188 240.244
R17073 GND.n7366 GND.n6204 240.244
R17074 GND.n7362 GND.n6204 240.244
R17075 GND.n7362 GND.n6209 240.244
R17076 GND.n7354 GND.n6209 240.244
R17077 GND.n7354 GND.n6225 240.244
R17078 GND.n7350 GND.n6225 240.244
R17079 GND.n7350 GND.n6230 240.244
R17080 GND.n7342 GND.n6230 240.244
R17081 GND.n7342 GND.n6245 240.244
R17082 GND.n7338 GND.n6245 240.244
R17083 GND.n7338 GND.n6250 240.244
R17084 GND.n6470 GND.n6250 240.244
R17085 GND.n6996 GND.n6470 240.244
R17086 GND.n6996 GND.n95 240.244
R17087 GND.n7005 GND.n95 240.244
R17088 GND.n7006 GND.n7005 240.244
R17089 GND.n7006 GND.n115 240.244
R17090 GND.n11103 GND.n115 240.244
R17091 GND.n11103 GND.n116 240.244
R17092 GND.n11099 GND.n116 240.244
R17093 GND.n11099 GND.n122 240.244
R17094 GND.n11091 GND.n122 240.244
R17095 GND.n11091 GND.n136 240.244
R17096 GND.n11087 GND.n136 240.244
R17097 GND.n11087 GND.n141 240.244
R17098 GND.n11079 GND.n141 240.244
R17099 GND.n11079 GND.n157 240.244
R17100 GND.n11075 GND.n157 240.244
R17101 GND.n11075 GND.n162 240.244
R17102 GND.n11067 GND.n162 240.244
R17103 GND.n11067 GND.n178 240.244
R17104 GND.n11063 GND.n178 240.244
R17105 GND.n11063 GND.n183 240.244
R17106 GND.n11055 GND.n183 240.244
R17107 GND.n11055 GND.n199 240.244
R17108 GND.n11051 GND.n199 240.244
R17109 GND.n11051 GND.n204 240.244
R17110 GND.n11043 GND.n204 240.244
R17111 GND.n11043 GND.n220 240.244
R17112 GND.n11039 GND.n220 240.244
R17113 GND.n11039 GND.n225 240.244
R17114 GND.n11031 GND.n225 240.244
R17115 GND.n11031 GND.n241 240.244
R17116 GND.n11027 GND.n241 240.244
R17117 GND.n11027 GND.n246 240.244
R17118 GND.n11019 GND.n246 240.244
R17119 GND.n11019 GND.n261 240.244
R17120 GND.n11015 GND.n261 240.244
R17121 GND.n11015 GND.n266 240.244
R17122 GND.n11007 GND.n266 240.244
R17123 GND.n11007 GND.n282 240.244
R17124 GND.n11003 GND.n282 240.244
R17125 GND.n11003 GND.n287 240.244
R17126 GND.n10995 GND.n287 240.244
R17127 GND.n10995 GND.n303 240.244
R17128 GND.n10991 GND.n303 240.244
R17129 GND.n10991 GND.n308 240.244
R17130 GND.n10983 GND.n308 240.244
R17131 GND.n10983 GND.n324 240.244
R17132 GND.n10979 GND.n324 240.244
R17133 GND.n10979 GND.n329 240.244
R17134 GND.n10971 GND.n329 240.244
R17135 GND.n10971 GND.n345 240.244
R17136 GND.n10967 GND.n345 240.244
R17137 GND.n10967 GND.n350 240.244
R17138 GND.n10959 GND.n350 240.244
R17139 GND.n10959 GND.n366 240.244
R17140 GND.n10955 GND.n366 240.244
R17141 GND.n10955 GND.n371 240.244
R17142 GND.n10947 GND.n371 240.244
R17143 GND.n10947 GND.n387 240.244
R17144 GND.n10943 GND.n387 240.244
R17145 GND.n10943 GND.n392 240.244
R17146 GND.n10935 GND.n392 240.244
R17147 GND.n10935 GND.n408 240.244
R17148 GND.n10931 GND.n408 240.244
R17149 GND.n10931 GND.n413 240.244
R17150 GND.n10923 GND.n413 240.244
R17151 GND.n10923 GND.n429 240.244
R17152 GND.n10919 GND.n429 240.244
R17153 GND.n10919 GND.n434 240.244
R17154 GND.n10911 GND.n434 240.244
R17155 GND.n9051 GND.n1460 240.244
R17156 GND.n9055 GND.n1460 240.244
R17157 GND.n9055 GND.n1456 240.244
R17158 GND.n9061 GND.n1456 240.244
R17159 GND.n9061 GND.n1454 240.244
R17160 GND.n9065 GND.n1454 240.244
R17161 GND.n9065 GND.n1450 240.244
R17162 GND.n9071 GND.n1450 240.244
R17163 GND.n9071 GND.n1448 240.244
R17164 GND.n9075 GND.n1448 240.244
R17165 GND.n9075 GND.n1444 240.244
R17166 GND.n9081 GND.n1444 240.244
R17167 GND.n9081 GND.n1442 240.244
R17168 GND.n9085 GND.n1442 240.244
R17169 GND.n9085 GND.n1438 240.244
R17170 GND.n9091 GND.n1438 240.244
R17171 GND.n9091 GND.n1436 240.244
R17172 GND.n9095 GND.n1436 240.244
R17173 GND.n9095 GND.n1432 240.244
R17174 GND.n9101 GND.n1432 240.244
R17175 GND.n9101 GND.n1430 240.244
R17176 GND.n9105 GND.n1430 240.244
R17177 GND.n9105 GND.n1426 240.244
R17178 GND.n9111 GND.n1426 240.244
R17179 GND.n9111 GND.n1424 240.244
R17180 GND.n9115 GND.n1424 240.244
R17181 GND.n9115 GND.n1420 240.244
R17182 GND.n9121 GND.n1420 240.244
R17183 GND.n9121 GND.n1418 240.244
R17184 GND.n9125 GND.n1418 240.244
R17185 GND.n9125 GND.n1414 240.244
R17186 GND.n9131 GND.n1414 240.244
R17187 GND.n9131 GND.n1412 240.244
R17188 GND.n9135 GND.n1412 240.244
R17189 GND.n9135 GND.n1408 240.244
R17190 GND.n9141 GND.n1408 240.244
R17191 GND.n9141 GND.n1406 240.244
R17192 GND.n9145 GND.n1406 240.244
R17193 GND.n9145 GND.n1402 240.244
R17194 GND.n9151 GND.n1402 240.244
R17195 GND.n9151 GND.n1400 240.244
R17196 GND.n9155 GND.n1400 240.244
R17197 GND.n9155 GND.n1396 240.244
R17198 GND.n9161 GND.n1396 240.244
R17199 GND.n9161 GND.n1394 240.244
R17200 GND.n9165 GND.n1394 240.244
R17201 GND.n9165 GND.n1390 240.244
R17202 GND.n9171 GND.n1390 240.244
R17203 GND.n9171 GND.n1388 240.244
R17204 GND.n9175 GND.n1388 240.244
R17205 GND.n9175 GND.n1384 240.244
R17206 GND.n9181 GND.n1384 240.244
R17207 GND.n9181 GND.n1382 240.244
R17208 GND.n9185 GND.n1382 240.244
R17209 GND.n9185 GND.n1378 240.244
R17210 GND.n9191 GND.n1378 240.244
R17211 GND.n9191 GND.n1376 240.244
R17212 GND.n9195 GND.n1376 240.244
R17213 GND.n9195 GND.n1372 240.244
R17214 GND.n9201 GND.n1372 240.244
R17215 GND.n9201 GND.n1370 240.244
R17216 GND.n9205 GND.n1370 240.244
R17217 GND.n9205 GND.n1366 240.244
R17218 GND.n9211 GND.n1366 240.244
R17219 GND.n9211 GND.n1364 240.244
R17220 GND.n9215 GND.n1364 240.244
R17221 GND.n9215 GND.n1360 240.244
R17222 GND.n9221 GND.n1360 240.244
R17223 GND.n9221 GND.n1358 240.244
R17224 GND.n9225 GND.n1358 240.244
R17225 GND.n9225 GND.n1354 240.244
R17226 GND.n9231 GND.n1354 240.244
R17227 GND.n9231 GND.n1352 240.244
R17228 GND.n9235 GND.n1352 240.244
R17229 GND.n9235 GND.n1348 240.244
R17230 GND.n9241 GND.n1348 240.244
R17231 GND.n9241 GND.n1346 240.244
R17232 GND.n9245 GND.n1346 240.244
R17233 GND.n9245 GND.n1342 240.244
R17234 GND.n9251 GND.n1342 240.244
R17235 GND.n9251 GND.n1340 240.244
R17236 GND.n9255 GND.n1340 240.244
R17237 GND.n9255 GND.n1336 240.244
R17238 GND.n9261 GND.n1336 240.244
R17239 GND.n9261 GND.n1334 240.244
R17240 GND.n9265 GND.n1334 240.244
R17241 GND.n9265 GND.n1330 240.244
R17242 GND.n9271 GND.n1330 240.244
R17243 GND.n9271 GND.n1328 240.244
R17244 GND.n9275 GND.n1328 240.244
R17245 GND.n9275 GND.n1324 240.244
R17246 GND.n9281 GND.n1324 240.244
R17247 GND.n9281 GND.n1322 240.244
R17248 GND.n9285 GND.n1322 240.244
R17249 GND.n9285 GND.n1318 240.244
R17250 GND.n9291 GND.n1318 240.244
R17251 GND.n9291 GND.n1316 240.244
R17252 GND.n9295 GND.n1316 240.244
R17253 GND.n9295 GND.n1312 240.244
R17254 GND.n9301 GND.n1312 240.244
R17255 GND.n9301 GND.n1310 240.244
R17256 GND.n9305 GND.n1310 240.244
R17257 GND.n9305 GND.n1306 240.244
R17258 GND.n9311 GND.n1306 240.244
R17259 GND.n9311 GND.n1304 240.244
R17260 GND.n9315 GND.n1304 240.244
R17261 GND.n9315 GND.n1300 240.244
R17262 GND.n9321 GND.n1300 240.244
R17263 GND.n9321 GND.n1298 240.244
R17264 GND.n9325 GND.n1298 240.244
R17265 GND.n9325 GND.n1294 240.244
R17266 GND.n9331 GND.n1294 240.244
R17267 GND.n9331 GND.n1292 240.244
R17268 GND.n9335 GND.n1292 240.244
R17269 GND.n9335 GND.n1288 240.244
R17270 GND.n9341 GND.n1288 240.244
R17271 GND.n9341 GND.n1286 240.244
R17272 GND.n9345 GND.n1286 240.244
R17273 GND.n9345 GND.n1282 240.244
R17274 GND.n9351 GND.n1282 240.244
R17275 GND.n9351 GND.n1280 240.244
R17276 GND.n9355 GND.n1280 240.244
R17277 GND.n9355 GND.n1276 240.244
R17278 GND.n9361 GND.n1276 240.244
R17279 GND.n9361 GND.n1274 240.244
R17280 GND.n9365 GND.n1274 240.244
R17281 GND.n9365 GND.n1270 240.244
R17282 GND.n9371 GND.n1270 240.244
R17283 GND.n9371 GND.n1268 240.244
R17284 GND.n9375 GND.n1268 240.244
R17285 GND.n9375 GND.n1264 240.244
R17286 GND.n9381 GND.n1264 240.244
R17287 GND.n9381 GND.n1262 240.244
R17288 GND.n9385 GND.n1262 240.244
R17289 GND.n9385 GND.n1258 240.244
R17290 GND.n9391 GND.n1258 240.244
R17291 GND.n9391 GND.n1256 240.244
R17292 GND.n9395 GND.n1256 240.244
R17293 GND.n9395 GND.n1252 240.244
R17294 GND.n9401 GND.n1252 240.244
R17295 GND.n9401 GND.n1250 240.244
R17296 GND.n9405 GND.n1250 240.244
R17297 GND.n9405 GND.n1246 240.244
R17298 GND.n9411 GND.n1246 240.244
R17299 GND.n9411 GND.n1244 240.244
R17300 GND.n9415 GND.n1244 240.244
R17301 GND.n9415 GND.n1240 240.244
R17302 GND.n9421 GND.n1240 240.244
R17303 GND.n9421 GND.n1238 240.244
R17304 GND.n9425 GND.n1238 240.244
R17305 GND.n9425 GND.n1234 240.244
R17306 GND.n9431 GND.n1234 240.244
R17307 GND.n9431 GND.n1232 240.244
R17308 GND.n9435 GND.n1232 240.244
R17309 GND.n9435 GND.n1228 240.244
R17310 GND.n9441 GND.n1228 240.244
R17311 GND.n9441 GND.n1226 240.244
R17312 GND.n9445 GND.n1226 240.244
R17313 GND.n9445 GND.n1222 240.244
R17314 GND.n9451 GND.n1222 240.244
R17315 GND.n9451 GND.n1220 240.244
R17316 GND.n9455 GND.n1220 240.244
R17317 GND.n9455 GND.n1216 240.244
R17318 GND.n9461 GND.n1216 240.244
R17319 GND.n9461 GND.n1214 240.244
R17320 GND.n9465 GND.n1214 240.244
R17321 GND.n9465 GND.n1210 240.244
R17322 GND.n9471 GND.n1210 240.244
R17323 GND.n9471 GND.n1208 240.244
R17324 GND.n9475 GND.n1208 240.244
R17325 GND.n9475 GND.n1204 240.244
R17326 GND.n9481 GND.n1204 240.244
R17327 GND.n9481 GND.n1202 240.244
R17328 GND.n9485 GND.n1202 240.244
R17329 GND.n9485 GND.n1198 240.244
R17330 GND.n9491 GND.n1198 240.244
R17331 GND.n9491 GND.n1196 240.244
R17332 GND.n9495 GND.n1196 240.244
R17333 GND.n9495 GND.n1192 240.244
R17334 GND.n9501 GND.n1192 240.244
R17335 GND.n9501 GND.n1190 240.244
R17336 GND.n9505 GND.n1190 240.244
R17337 GND.n9505 GND.n1186 240.244
R17338 GND.n9511 GND.n1186 240.244
R17339 GND.n9511 GND.n1184 240.244
R17340 GND.n9515 GND.n1184 240.244
R17341 GND.n9515 GND.n1180 240.244
R17342 GND.n9521 GND.n1180 240.244
R17343 GND.n9521 GND.n1178 240.244
R17344 GND.n9525 GND.n1178 240.244
R17345 GND.n9525 GND.n1174 240.244
R17346 GND.n9531 GND.n1174 240.244
R17347 GND.n9531 GND.n1172 240.244
R17348 GND.n9535 GND.n1172 240.244
R17349 GND.n9535 GND.n1168 240.244
R17350 GND.n9541 GND.n1168 240.244
R17351 GND.n9541 GND.n1166 240.244
R17352 GND.n9545 GND.n1166 240.244
R17353 GND.n9545 GND.n1162 240.244
R17354 GND.n9551 GND.n1162 240.244
R17355 GND.n9551 GND.n1160 240.244
R17356 GND.n9555 GND.n1160 240.244
R17357 GND.n9555 GND.n1156 240.244
R17358 GND.n9561 GND.n1156 240.244
R17359 GND.n9561 GND.n1154 240.244
R17360 GND.n9565 GND.n1154 240.244
R17361 GND.n9565 GND.n1150 240.244
R17362 GND.n9571 GND.n1150 240.244
R17363 GND.n9571 GND.n1148 240.244
R17364 GND.n9575 GND.n1148 240.244
R17365 GND.n9575 GND.n1144 240.244
R17366 GND.n9581 GND.n1144 240.244
R17367 GND.n9581 GND.n1142 240.244
R17368 GND.n9585 GND.n1142 240.244
R17369 GND.n9585 GND.n1138 240.244
R17370 GND.n9591 GND.n1138 240.244
R17371 GND.n9591 GND.n1136 240.244
R17372 GND.n9595 GND.n1136 240.244
R17373 GND.n9595 GND.n1132 240.244
R17374 GND.n9601 GND.n1132 240.244
R17375 GND.n9601 GND.n1130 240.244
R17376 GND.n9605 GND.n1130 240.244
R17377 GND.n9605 GND.n1126 240.244
R17378 GND.n9611 GND.n1126 240.244
R17379 GND.n9611 GND.n1124 240.244
R17380 GND.n9615 GND.n1124 240.244
R17381 GND.n9615 GND.n1120 240.244
R17382 GND.n9621 GND.n1120 240.244
R17383 GND.n9621 GND.n1118 240.244
R17384 GND.n9625 GND.n1118 240.244
R17385 GND.n9625 GND.n1114 240.244
R17386 GND.n9631 GND.n1114 240.244
R17387 GND.n9631 GND.n1112 240.244
R17388 GND.n9635 GND.n1112 240.244
R17389 GND.n9635 GND.n1108 240.244
R17390 GND.n9641 GND.n1108 240.244
R17391 GND.n9641 GND.n1106 240.244
R17392 GND.n9645 GND.n1106 240.244
R17393 GND.n9645 GND.n1102 240.244
R17394 GND.n9651 GND.n1102 240.244
R17395 GND.n9651 GND.n1100 240.244
R17396 GND.n9655 GND.n1100 240.244
R17397 GND.n9655 GND.n1096 240.244
R17398 GND.n9661 GND.n1096 240.244
R17399 GND.n9661 GND.n1094 240.244
R17400 GND.n9665 GND.n1094 240.244
R17401 GND.n9665 GND.n1090 240.244
R17402 GND.n9671 GND.n1090 240.244
R17403 GND.n9671 GND.n1088 240.244
R17404 GND.n9675 GND.n1088 240.244
R17405 GND.n9675 GND.n1084 240.244
R17406 GND.n9681 GND.n1084 240.244
R17407 GND.n9681 GND.n1082 240.244
R17408 GND.n9685 GND.n1082 240.244
R17409 GND.n9685 GND.n1078 240.244
R17410 GND.n9691 GND.n1078 240.244
R17411 GND.n9691 GND.n1076 240.244
R17412 GND.n9695 GND.n1076 240.244
R17413 GND.n9695 GND.n1072 240.244
R17414 GND.n9701 GND.n1072 240.244
R17415 GND.n9701 GND.n1070 240.244
R17416 GND.n9705 GND.n1070 240.244
R17417 GND.n9705 GND.n1066 240.244
R17418 GND.n9711 GND.n1066 240.244
R17419 GND.n9711 GND.n1064 240.244
R17420 GND.n9715 GND.n1064 240.244
R17421 GND.n9715 GND.n1060 240.244
R17422 GND.n9721 GND.n1060 240.244
R17423 GND.n9721 GND.n1058 240.244
R17424 GND.n9725 GND.n1058 240.244
R17425 GND.n9725 GND.n1054 240.244
R17426 GND.n9731 GND.n1054 240.244
R17427 GND.n9731 GND.n1052 240.244
R17428 GND.n9735 GND.n1052 240.244
R17429 GND.n9735 GND.n1048 240.244
R17430 GND.n9741 GND.n1048 240.244
R17431 GND.n9741 GND.n1046 240.244
R17432 GND.n9745 GND.n1046 240.244
R17433 GND.n9745 GND.n1042 240.244
R17434 GND.n9751 GND.n1042 240.244
R17435 GND.n9751 GND.n1040 240.244
R17436 GND.n9755 GND.n1040 240.244
R17437 GND.n9755 GND.n1036 240.244
R17438 GND.n9761 GND.n1036 240.244
R17439 GND.n9761 GND.n1034 240.244
R17440 GND.n9765 GND.n1034 240.244
R17441 GND.n9765 GND.n1030 240.244
R17442 GND.n9771 GND.n1030 240.244
R17443 GND.n9771 GND.n1028 240.244
R17444 GND.n9775 GND.n1028 240.244
R17445 GND.n9775 GND.n1024 240.244
R17446 GND.n9781 GND.n1024 240.244
R17447 GND.n9781 GND.n1022 240.244
R17448 GND.n9785 GND.n1022 240.244
R17449 GND.n9785 GND.n1018 240.244
R17450 GND.n9791 GND.n1018 240.244
R17451 GND.n9791 GND.n1016 240.244
R17452 GND.n9795 GND.n1016 240.244
R17453 GND.n9795 GND.n1012 240.244
R17454 GND.n9801 GND.n1012 240.244
R17455 GND.n9801 GND.n1010 240.244
R17456 GND.n9805 GND.n1010 240.244
R17457 GND.n9805 GND.n1006 240.244
R17458 GND.n9811 GND.n1006 240.244
R17459 GND.n9811 GND.n1004 240.244
R17460 GND.n9815 GND.n1004 240.244
R17461 GND.n9815 GND.n1000 240.244
R17462 GND.n9821 GND.n1000 240.244
R17463 GND.n9821 GND.n998 240.244
R17464 GND.n9825 GND.n998 240.244
R17465 GND.n9825 GND.n994 240.244
R17466 GND.n9831 GND.n994 240.244
R17467 GND.n9831 GND.n992 240.244
R17468 GND.n9835 GND.n992 240.244
R17469 GND.n9835 GND.n988 240.244
R17470 GND.n9841 GND.n988 240.244
R17471 GND.n9841 GND.n986 240.244
R17472 GND.n9845 GND.n986 240.244
R17473 GND.n9845 GND.n982 240.244
R17474 GND.n9851 GND.n982 240.244
R17475 GND.n9851 GND.n980 240.244
R17476 GND.n9855 GND.n980 240.244
R17477 GND.n9855 GND.n976 240.244
R17478 GND.n9861 GND.n976 240.244
R17479 GND.n9861 GND.n974 240.244
R17480 GND.n9865 GND.n974 240.244
R17481 GND.n9865 GND.n970 240.244
R17482 GND.n9871 GND.n970 240.244
R17483 GND.n9871 GND.n968 240.244
R17484 GND.n9875 GND.n968 240.244
R17485 GND.n9875 GND.n964 240.244
R17486 GND.n9881 GND.n964 240.244
R17487 GND.n9881 GND.n962 240.244
R17488 GND.n9885 GND.n962 240.244
R17489 GND.n9885 GND.n958 240.244
R17490 GND.n9891 GND.n958 240.244
R17491 GND.n9891 GND.n956 240.244
R17492 GND.n9895 GND.n956 240.244
R17493 GND.n9895 GND.n952 240.244
R17494 GND.n9901 GND.n952 240.244
R17495 GND.n9901 GND.n950 240.244
R17496 GND.n9905 GND.n950 240.244
R17497 GND.n9905 GND.n946 240.244
R17498 GND.n9911 GND.n946 240.244
R17499 GND.n9911 GND.n944 240.244
R17500 GND.n9915 GND.n944 240.244
R17501 GND.n9915 GND.n940 240.244
R17502 GND.n9921 GND.n940 240.244
R17503 GND.n9921 GND.n938 240.244
R17504 GND.n9925 GND.n938 240.244
R17505 GND.n9925 GND.n934 240.244
R17506 GND.n9931 GND.n934 240.244
R17507 GND.n9931 GND.n932 240.244
R17508 GND.n9935 GND.n932 240.244
R17509 GND.n9935 GND.n928 240.244
R17510 GND.n9941 GND.n928 240.244
R17511 GND.n9941 GND.n926 240.244
R17512 GND.n9945 GND.n926 240.244
R17513 GND.n9945 GND.n922 240.244
R17514 GND.n9951 GND.n922 240.244
R17515 GND.n9951 GND.n920 240.244
R17516 GND.n9955 GND.n920 240.244
R17517 GND.n9955 GND.n916 240.244
R17518 GND.n9961 GND.n916 240.244
R17519 GND.n9961 GND.n914 240.244
R17520 GND.n9965 GND.n914 240.244
R17521 GND.n9965 GND.n910 240.244
R17522 GND.n9971 GND.n910 240.244
R17523 GND.n9971 GND.n908 240.244
R17524 GND.n9975 GND.n908 240.244
R17525 GND.n9975 GND.n904 240.244
R17526 GND.n9981 GND.n904 240.244
R17527 GND.n9981 GND.n902 240.244
R17528 GND.n9985 GND.n902 240.244
R17529 GND.n9985 GND.n898 240.244
R17530 GND.n9991 GND.n898 240.244
R17531 GND.n9991 GND.n896 240.244
R17532 GND.n9995 GND.n896 240.244
R17533 GND.n9995 GND.n892 240.244
R17534 GND.n10001 GND.n892 240.244
R17535 GND.n10001 GND.n890 240.244
R17536 GND.n10005 GND.n890 240.244
R17537 GND.n10005 GND.n886 240.244
R17538 GND.n10011 GND.n886 240.244
R17539 GND.n10011 GND.n884 240.244
R17540 GND.n10015 GND.n884 240.244
R17541 GND.n10015 GND.n880 240.244
R17542 GND.n10021 GND.n880 240.244
R17543 GND.n10021 GND.n878 240.244
R17544 GND.n10025 GND.n878 240.244
R17545 GND.n10025 GND.n874 240.244
R17546 GND.n10031 GND.n874 240.244
R17547 GND.n10031 GND.n872 240.244
R17548 GND.n10035 GND.n872 240.244
R17549 GND.n10035 GND.n868 240.244
R17550 GND.n10041 GND.n868 240.244
R17551 GND.n10041 GND.n866 240.244
R17552 GND.n10045 GND.n866 240.244
R17553 GND.n10045 GND.n862 240.244
R17554 GND.n10051 GND.n862 240.244
R17555 GND.n10051 GND.n860 240.244
R17556 GND.n10055 GND.n860 240.244
R17557 GND.n10055 GND.n856 240.244
R17558 GND.n10061 GND.n856 240.244
R17559 GND.n10061 GND.n854 240.244
R17560 GND.n10065 GND.n854 240.244
R17561 GND.n10065 GND.n850 240.244
R17562 GND.n10071 GND.n850 240.244
R17563 GND.n10071 GND.n848 240.244
R17564 GND.n10075 GND.n848 240.244
R17565 GND.n10075 GND.n844 240.244
R17566 GND.n10081 GND.n844 240.244
R17567 GND.n10081 GND.n842 240.244
R17568 GND.n10085 GND.n842 240.244
R17569 GND.n10085 GND.n838 240.244
R17570 GND.n10091 GND.n838 240.244
R17571 GND.n10091 GND.n836 240.244
R17572 GND.n10095 GND.n836 240.244
R17573 GND.n10095 GND.n832 240.244
R17574 GND.n10101 GND.n832 240.244
R17575 GND.n10101 GND.n830 240.244
R17576 GND.n10105 GND.n830 240.244
R17577 GND.n10105 GND.n826 240.244
R17578 GND.n10111 GND.n826 240.244
R17579 GND.n10111 GND.n824 240.244
R17580 GND.n10115 GND.n824 240.244
R17581 GND.n10115 GND.n820 240.244
R17582 GND.n10121 GND.n820 240.244
R17583 GND.n10121 GND.n818 240.244
R17584 GND.n10125 GND.n818 240.244
R17585 GND.n10125 GND.n814 240.244
R17586 GND.n10131 GND.n814 240.244
R17587 GND.n10131 GND.n812 240.244
R17588 GND.n10135 GND.n812 240.244
R17589 GND.n10135 GND.n808 240.244
R17590 GND.n10141 GND.n808 240.244
R17591 GND.n10141 GND.n806 240.244
R17592 GND.n10145 GND.n806 240.244
R17593 GND.n10145 GND.n802 240.244
R17594 GND.n10151 GND.n802 240.244
R17595 GND.n10151 GND.n800 240.244
R17596 GND.n10155 GND.n800 240.244
R17597 GND.n10155 GND.n796 240.244
R17598 GND.n10161 GND.n796 240.244
R17599 GND.n10161 GND.n794 240.244
R17600 GND.n10165 GND.n794 240.244
R17601 GND.n10165 GND.n790 240.244
R17602 GND.n10171 GND.n790 240.244
R17603 GND.n10171 GND.n788 240.244
R17604 GND.n10175 GND.n788 240.244
R17605 GND.n10175 GND.n784 240.244
R17606 GND.n10181 GND.n784 240.244
R17607 GND.n10181 GND.n782 240.244
R17608 GND.n10185 GND.n782 240.244
R17609 GND.n10185 GND.n778 240.244
R17610 GND.n10191 GND.n778 240.244
R17611 GND.n10191 GND.n776 240.244
R17612 GND.n10195 GND.n776 240.244
R17613 GND.n10195 GND.n772 240.244
R17614 GND.n10201 GND.n772 240.244
R17615 GND.n10201 GND.n770 240.244
R17616 GND.n10205 GND.n770 240.244
R17617 GND.n10205 GND.n766 240.244
R17618 GND.n10211 GND.n766 240.244
R17619 GND.n10211 GND.n764 240.244
R17620 GND.n10215 GND.n764 240.244
R17621 GND.n10215 GND.n760 240.244
R17622 GND.n10221 GND.n760 240.244
R17623 GND.n10221 GND.n758 240.244
R17624 GND.n10225 GND.n758 240.244
R17625 GND.n10225 GND.n754 240.244
R17626 GND.n10231 GND.n754 240.244
R17627 GND.n10231 GND.n752 240.244
R17628 GND.n10235 GND.n752 240.244
R17629 GND.n10235 GND.n748 240.244
R17630 GND.n10241 GND.n748 240.244
R17631 GND.n10241 GND.n746 240.244
R17632 GND.n10245 GND.n746 240.244
R17633 GND.n10245 GND.n742 240.244
R17634 GND.n10251 GND.n742 240.244
R17635 GND.n10251 GND.n740 240.244
R17636 GND.n10255 GND.n740 240.244
R17637 GND.n10255 GND.n736 240.244
R17638 GND.n10261 GND.n736 240.244
R17639 GND.n10261 GND.n734 240.244
R17640 GND.n10265 GND.n734 240.244
R17641 GND.n10265 GND.n730 240.244
R17642 GND.n10271 GND.n730 240.244
R17643 GND.n10271 GND.n728 240.244
R17644 GND.n10275 GND.n728 240.244
R17645 GND.n10275 GND.n724 240.244
R17646 GND.n10281 GND.n724 240.244
R17647 GND.n10281 GND.n722 240.244
R17648 GND.n10285 GND.n722 240.244
R17649 GND.n10285 GND.n718 240.244
R17650 GND.n10291 GND.n718 240.244
R17651 GND.n10291 GND.n716 240.244
R17652 GND.n10295 GND.n716 240.244
R17653 GND.n10295 GND.n712 240.244
R17654 GND.n10301 GND.n712 240.244
R17655 GND.n10301 GND.n710 240.244
R17656 GND.n10305 GND.n710 240.244
R17657 GND.n10305 GND.n706 240.244
R17658 GND.n10311 GND.n706 240.244
R17659 GND.n10311 GND.n704 240.244
R17660 GND.n10315 GND.n704 240.244
R17661 GND.n10315 GND.n700 240.244
R17662 GND.n10321 GND.n700 240.244
R17663 GND.n10321 GND.n698 240.244
R17664 GND.n10325 GND.n698 240.244
R17665 GND.n10325 GND.n694 240.244
R17666 GND.n10331 GND.n694 240.244
R17667 GND.n10331 GND.n692 240.244
R17668 GND.n10335 GND.n692 240.244
R17669 GND.n10335 GND.n688 240.244
R17670 GND.n10341 GND.n688 240.244
R17671 GND.n10341 GND.n686 240.244
R17672 GND.n10345 GND.n686 240.244
R17673 GND.n10345 GND.n682 240.244
R17674 GND.n10351 GND.n682 240.244
R17675 GND.n10351 GND.n680 240.244
R17676 GND.n10355 GND.n680 240.244
R17677 GND.n10355 GND.n676 240.244
R17678 GND.n10361 GND.n676 240.244
R17679 GND.n10361 GND.n674 240.244
R17680 GND.n10365 GND.n674 240.244
R17681 GND.n10365 GND.n670 240.244
R17682 GND.n10371 GND.n670 240.244
R17683 GND.n10371 GND.n668 240.244
R17684 GND.n10375 GND.n668 240.244
R17685 GND.n10375 GND.n664 240.244
R17686 GND.n10382 GND.n664 240.244
R17687 GND.n10382 GND.n662 240.244
R17688 GND.n10386 GND.n659 240.244
R17689 GND.n10392 GND.n659 240.244
R17690 GND.n10392 GND.n657 240.244
R17691 GND.n10396 GND.n657 240.244
R17692 GND.n10396 GND.n653 240.244
R17693 GND.n10402 GND.n653 240.244
R17694 GND.n10402 GND.n651 240.244
R17695 GND.n10406 GND.n651 240.244
R17696 GND.n10406 GND.n647 240.244
R17697 GND.n10412 GND.n647 240.244
R17698 GND.n10412 GND.n645 240.244
R17699 GND.n10416 GND.n645 240.244
R17700 GND.n10416 GND.n641 240.244
R17701 GND.n10422 GND.n641 240.244
R17702 GND.n10422 GND.n639 240.244
R17703 GND.n10426 GND.n639 240.244
R17704 GND.n10426 GND.n635 240.244
R17705 GND.n10432 GND.n635 240.244
R17706 GND.n10432 GND.n633 240.244
R17707 GND.n10436 GND.n633 240.244
R17708 GND.n10436 GND.n629 240.244
R17709 GND.n10442 GND.n629 240.244
R17710 GND.n10442 GND.n627 240.244
R17711 GND.n10446 GND.n627 240.244
R17712 GND.n10446 GND.n623 240.244
R17713 GND.n10452 GND.n623 240.244
R17714 GND.n10452 GND.n621 240.244
R17715 GND.n10456 GND.n621 240.244
R17716 GND.n10456 GND.n617 240.244
R17717 GND.n10462 GND.n617 240.244
R17718 GND.n10462 GND.n615 240.244
R17719 GND.n10466 GND.n615 240.244
R17720 GND.n10466 GND.n611 240.244
R17721 GND.n10472 GND.n611 240.244
R17722 GND.n10472 GND.n609 240.244
R17723 GND.n10476 GND.n609 240.244
R17724 GND.n10476 GND.n605 240.244
R17725 GND.n10482 GND.n605 240.244
R17726 GND.n10482 GND.n603 240.244
R17727 GND.n10486 GND.n603 240.244
R17728 GND.n10486 GND.n599 240.244
R17729 GND.n10492 GND.n599 240.244
R17730 GND.n10492 GND.n597 240.244
R17731 GND.n10496 GND.n597 240.244
R17732 GND.n10496 GND.n593 240.244
R17733 GND.n10502 GND.n593 240.244
R17734 GND.n10502 GND.n591 240.244
R17735 GND.n10506 GND.n591 240.244
R17736 GND.n10506 GND.n587 240.244
R17737 GND.n10512 GND.n587 240.244
R17738 GND.n10512 GND.n585 240.244
R17739 GND.n10516 GND.n585 240.244
R17740 GND.n10516 GND.n581 240.244
R17741 GND.n10522 GND.n581 240.244
R17742 GND.n10522 GND.n579 240.244
R17743 GND.n10526 GND.n579 240.244
R17744 GND.n10526 GND.n575 240.244
R17745 GND.n10533 GND.n575 240.244
R17746 GND.n8929 GND.n1579 240.244
R17747 GND.n1585 GND.n1579 240.244
R17748 GND.n8922 GND.n1585 240.244
R17749 GND.n8922 GND.n1586 240.244
R17750 GND.n8918 GND.n1586 240.244
R17751 GND.n8918 GND.n1589 240.244
R17752 GND.n8914 GND.n1589 240.244
R17753 GND.n8914 GND.n1594 240.244
R17754 GND.n8910 GND.n1594 240.244
R17755 GND.n8910 GND.n1596 240.244
R17756 GND.n8906 GND.n1596 240.244
R17757 GND.n8906 GND.n1602 240.244
R17758 GND.n8902 GND.n1602 240.244
R17759 GND.n8902 GND.n1604 240.244
R17760 GND.n8898 GND.n1604 240.244
R17761 GND.n8898 GND.n1610 240.244
R17762 GND.n8894 GND.n1610 240.244
R17763 GND.n8894 GND.n1612 240.244
R17764 GND.n8890 GND.n1612 240.244
R17765 GND.n8890 GND.n1618 240.244
R17766 GND.n8886 GND.n1618 240.244
R17767 GND.n8886 GND.n1620 240.244
R17768 GND.n8882 GND.n1620 240.244
R17769 GND.n8882 GND.n1626 240.244
R17770 GND.n8878 GND.n1626 240.244
R17771 GND.n8878 GND.n1628 240.244
R17772 GND.n8874 GND.n1628 240.244
R17773 GND.n8874 GND.n1634 240.244
R17774 GND.n8870 GND.n1634 240.244
R17775 GND.n8870 GND.n1636 240.244
R17776 GND.n8866 GND.n1636 240.244
R17777 GND.n8866 GND.n1642 240.244
R17778 GND.n8862 GND.n1642 240.244
R17779 GND.n8862 GND.n1644 240.244
R17780 GND.n8858 GND.n1644 240.244
R17781 GND.n8858 GND.n1650 240.244
R17782 GND.n8854 GND.n1650 240.244
R17783 GND.n8854 GND.n1652 240.244
R17784 GND.n8850 GND.n1652 240.244
R17785 GND.n8850 GND.n1658 240.244
R17786 GND.n8846 GND.n1658 240.244
R17787 GND.n8846 GND.n1660 240.244
R17788 GND.n8842 GND.n1660 240.244
R17789 GND.n8842 GND.n1666 240.244
R17790 GND.n8838 GND.n1666 240.244
R17791 GND.n8838 GND.n1668 240.244
R17792 GND.n8834 GND.n1668 240.244
R17793 GND.n8834 GND.n1674 240.244
R17794 GND.n8830 GND.n1674 240.244
R17795 GND.n8830 GND.n1676 240.244
R17796 GND.n8826 GND.n1676 240.244
R17797 GND.n8826 GND.n1682 240.244
R17798 GND.n8822 GND.n1682 240.244
R17799 GND.n8822 GND.n1684 240.244
R17800 GND.n8818 GND.n1684 240.244
R17801 GND.n8818 GND.n1690 240.244
R17802 GND.n1806 GND.n1690 240.244
R17803 GND.n8696 GND.n1806 240.244
R17804 GND.n8696 GND.n1807 240.244
R17805 GND.n8692 GND.n1807 240.244
R17806 GND.n8692 GND.n1815 240.244
R17807 GND.n2973 GND.n1815 240.244
R17808 GND.n2974 GND.n2973 240.244
R17809 GND.n2974 GND.n2967 240.244
R17810 GND.n3149 GND.n2967 240.244
R17811 GND.n3149 GND.n2968 240.244
R17812 GND.n3145 GND.n2968 240.244
R17813 GND.n3145 GND.n3144 240.244
R17814 GND.n3144 GND.n3143 240.244
R17815 GND.n3143 GND.n2982 240.244
R17816 GND.n3139 GND.n2982 240.244
R17817 GND.n3139 GND.n3138 240.244
R17818 GND.n3138 GND.n3137 240.244
R17819 GND.n3137 GND.n2988 240.244
R17820 GND.n3133 GND.n2988 240.244
R17821 GND.n3133 GND.n3132 240.244
R17822 GND.n3132 GND.n3131 240.244
R17823 GND.n3131 GND.n2994 240.244
R17824 GND.n3127 GND.n2994 240.244
R17825 GND.n3127 GND.n3126 240.244
R17826 GND.n3126 GND.n3125 240.244
R17827 GND.n3125 GND.n3000 240.244
R17828 GND.n3121 GND.n3000 240.244
R17829 GND.n3121 GND.n3120 240.244
R17830 GND.n3120 GND.n3119 240.244
R17831 GND.n3119 GND.n3006 240.244
R17832 GND.n3115 GND.n3006 240.244
R17833 GND.n3115 GND.n3114 240.244
R17834 GND.n3114 GND.n3113 240.244
R17835 GND.n3113 GND.n3012 240.244
R17836 GND.n3109 GND.n3012 240.244
R17837 GND.n3109 GND.n3108 240.244
R17838 GND.n3108 GND.n3107 240.244
R17839 GND.n3107 GND.n3018 240.244
R17840 GND.n3103 GND.n3018 240.244
R17841 GND.n3103 GND.n3102 240.244
R17842 GND.n3102 GND.n3101 240.244
R17843 GND.n3101 GND.n3024 240.244
R17844 GND.n3097 GND.n3024 240.244
R17845 GND.n3097 GND.n3096 240.244
R17846 GND.n3096 GND.n3095 240.244
R17847 GND.n3095 GND.n3030 240.244
R17848 GND.n3091 GND.n3030 240.244
R17849 GND.n3091 GND.n3090 240.244
R17850 GND.n3090 GND.n3089 240.244
R17851 GND.n3089 GND.n3036 240.244
R17852 GND.n3085 GND.n3036 240.244
R17853 GND.n3085 GND.n3084 240.244
R17854 GND.n3084 GND.n3083 240.244
R17855 GND.n3083 GND.n3042 240.244
R17856 GND.n3079 GND.n3042 240.244
R17857 GND.n3079 GND.n3078 240.244
R17858 GND.n3078 GND.n3077 240.244
R17859 GND.n3077 GND.n3048 240.244
R17860 GND.n3073 GND.n3048 240.244
R17861 GND.n3073 GND.n3072 240.244
R17862 GND.n3072 GND.n3071 240.244
R17863 GND.n3071 GND.n3054 240.244
R17864 GND.n3067 GND.n3054 240.244
R17865 GND.n3067 GND.n3066 240.244
R17866 GND.n3066 GND.n3063 240.244
R17867 GND.n3063 GND.n2510 240.244
R17868 GND.n3485 GND.n2510 240.244
R17869 GND.n3485 GND.n2511 240.244
R17870 GND.n3480 GND.n2511 240.244
R17871 GND.n3480 GND.n2514 240.244
R17872 GND.n2532 GND.n2514 240.244
R17873 GND.n3468 GND.n2532 240.244
R17874 GND.n3468 GND.n2533 240.244
R17875 GND.n3463 GND.n2533 240.244
R17876 GND.n3463 GND.n2648 240.244
R17877 GND.n2648 GND.n2537 240.244
R17878 GND.n2644 GND.n2537 240.244
R17879 GND.n2644 GND.n2643 240.244
R17880 GND.n2643 GND.n2642 240.244
R17881 GND.n2642 GND.n2541 240.244
R17882 GND.n2638 GND.n2541 240.244
R17883 GND.n2638 GND.n2637 240.244
R17884 GND.n2637 GND.n2636 240.244
R17885 GND.n2636 GND.n2547 240.244
R17886 GND.n2632 GND.n2547 240.244
R17887 GND.n2632 GND.n2631 240.244
R17888 GND.n2631 GND.n2630 240.244
R17889 GND.n2630 GND.n2553 240.244
R17890 GND.n2626 GND.n2553 240.244
R17891 GND.n2626 GND.n2625 240.244
R17892 GND.n2625 GND.n2624 240.244
R17893 GND.n2624 GND.n2559 240.244
R17894 GND.n2620 GND.n2559 240.244
R17895 GND.n2620 GND.n2619 240.244
R17896 GND.n2619 GND.n2618 240.244
R17897 GND.n2618 GND.n2565 240.244
R17898 GND.n2614 GND.n2565 240.244
R17899 GND.n2614 GND.n2613 240.244
R17900 GND.n2613 GND.n2612 240.244
R17901 GND.n2612 GND.n2571 240.244
R17902 GND.n2608 GND.n2571 240.244
R17903 GND.n2608 GND.n2607 240.244
R17904 GND.n2607 GND.n2603 240.244
R17905 GND.n2603 GND.n2577 240.244
R17906 GND.n2599 GND.n2577 240.244
R17907 GND.n2599 GND.n2598 240.244
R17908 GND.n2598 GND.n2597 240.244
R17909 GND.n2597 GND.n2583 240.244
R17910 GND.n2593 GND.n2583 240.244
R17911 GND.n2593 GND.n2592 240.244
R17912 GND.n2592 GND.n2327 240.244
R17913 GND.n3693 GND.n2327 240.244
R17914 GND.n3694 GND.n3693 240.244
R17915 GND.n3694 GND.n2322 240.244
R17916 GND.n8177 GND.n2322 240.244
R17917 GND.n8177 GND.n2323 240.244
R17918 GND.n8173 GND.n2323 240.244
R17919 GND.n8173 GND.n8172 240.244
R17920 GND.n8172 GND.n8171 240.244
R17921 GND.n8171 GND.n3702 240.244
R17922 GND.n8167 GND.n3702 240.244
R17923 GND.n8167 GND.n8166 240.244
R17924 GND.n8166 GND.n8165 240.244
R17925 GND.n8165 GND.n3708 240.244
R17926 GND.n8161 GND.n3708 240.244
R17927 GND.n8161 GND.n8160 240.244
R17928 GND.n8160 GND.n8159 240.244
R17929 GND.n8159 GND.n3714 240.244
R17930 GND.n8155 GND.n3714 240.244
R17931 GND.n8155 GND.n8154 240.244
R17932 GND.n8154 GND.n8153 240.244
R17933 GND.n8153 GND.n3720 240.244
R17934 GND.n8149 GND.n3720 240.244
R17935 GND.n8149 GND.n8148 240.244
R17936 GND.n8148 GND.n8147 240.244
R17937 GND.n8147 GND.n3726 240.244
R17938 GND.n8143 GND.n3726 240.244
R17939 GND.n8143 GND.n8142 240.244
R17940 GND.n8142 GND.n8141 240.244
R17941 GND.n8141 GND.n3732 240.244
R17942 GND.n8137 GND.n3732 240.244
R17943 GND.n8137 GND.n8136 240.244
R17944 GND.n8136 GND.n3738 240.244
R17945 GND.n8132 GND.n3738 240.244
R17946 GND.n8132 GND.n3740 240.244
R17947 GND.n8128 GND.n3740 240.244
R17948 GND.n8128 GND.n3748 240.244
R17949 GND.n8118 GND.n3748 240.244
R17950 GND.n8118 GND.n3773 240.244
R17951 GND.n8114 GND.n3773 240.244
R17952 GND.n8114 GND.n3779 240.244
R17953 GND.n8104 GND.n3779 240.244
R17954 GND.n8104 GND.n3789 240.244
R17955 GND.n8100 GND.n3789 240.244
R17956 GND.n8100 GND.n3795 240.244
R17957 GND.n8090 GND.n3795 240.244
R17958 GND.n8090 GND.n3807 240.244
R17959 GND.n8086 GND.n3807 240.244
R17960 GND.n8086 GND.n3813 240.244
R17961 GND.n8076 GND.n3813 240.244
R17962 GND.n8076 GND.n3825 240.244
R17963 GND.n8072 GND.n3825 240.244
R17964 GND.n8072 GND.n3831 240.244
R17965 GND.n8062 GND.n3831 240.244
R17966 GND.n8062 GND.n3843 240.244
R17967 GND.n8058 GND.n3843 240.244
R17968 GND.n8058 GND.n3849 240.244
R17969 GND.n8004 GND.n3849 240.244
R17970 GND.n8004 GND.n3886 240.244
R17971 GND.n8000 GND.n3886 240.244
R17972 GND.n8000 GND.n3892 240.244
R17973 GND.n7992 GND.n3892 240.244
R17974 GND.n7992 GND.n3907 240.244
R17975 GND.n7988 GND.n3907 240.244
R17976 GND.n7988 GND.n3913 240.244
R17977 GND.n7980 GND.n3913 240.244
R17978 GND.n7980 GND.n3927 240.244
R17979 GND.n7976 GND.n3927 240.244
R17980 GND.n7976 GND.n3933 240.244
R17981 GND.n7968 GND.n3933 240.244
R17982 GND.n7968 GND.n3947 240.244
R17983 GND.n7964 GND.n3947 240.244
R17984 GND.n7964 GND.n3953 240.244
R17985 GND.n7956 GND.n3953 240.244
R17986 GND.n7956 GND.n3967 240.244
R17987 GND.n7952 GND.n3967 240.244
R17988 GND.n7952 GND.n3973 240.244
R17989 GND.n7944 GND.n3973 240.244
R17990 GND.n7944 GND.n3987 240.244
R17991 GND.n7940 GND.n3987 240.244
R17992 GND.n7940 GND.n3993 240.244
R17993 GND.n7932 GND.n3993 240.244
R17994 GND.n7932 GND.n4007 240.244
R17995 GND.n7928 GND.n4007 240.244
R17996 GND.n7928 GND.n4013 240.244
R17997 GND.n7920 GND.n4013 240.244
R17998 GND.n7920 GND.n4027 240.244
R17999 GND.n7916 GND.n4027 240.244
R18000 GND.n7916 GND.n4033 240.244
R18001 GND.n7908 GND.n4033 240.244
R18002 GND.n7908 GND.n4047 240.244
R18003 GND.n7904 GND.n4047 240.244
R18004 GND.n7904 GND.n4053 240.244
R18005 GND.n4076 GND.n4053 240.244
R18006 GND.n7889 GND.n4076 240.244
R18007 GND.n7889 GND.n4077 240.244
R18008 GND.n7885 GND.n4077 240.244
R18009 GND.n7885 GND.n4085 240.244
R18010 GND.n7877 GND.n4085 240.244
R18011 GND.n7877 GND.n4112 240.244
R18012 GND.n7873 GND.n4112 240.244
R18013 GND.n7873 GND.n4118 240.244
R18014 GND.n7865 GND.n4118 240.244
R18015 GND.n7865 GND.n4132 240.244
R18016 GND.n7861 GND.n4132 240.244
R18017 GND.n7861 GND.n4138 240.244
R18018 GND.n7853 GND.n4138 240.244
R18019 GND.n7853 GND.n4152 240.244
R18020 GND.n7849 GND.n4152 240.244
R18021 GND.n7849 GND.n4158 240.244
R18022 GND.n4181 GND.n4158 240.244
R18023 GND.n7834 GND.n4181 240.244
R18024 GND.n7834 GND.n4182 240.244
R18025 GND.n7830 GND.n4182 240.244
R18026 GND.n7830 GND.n4190 240.244
R18027 GND.n7822 GND.n4190 240.244
R18028 GND.n7822 GND.n4216 240.244
R18029 GND.n7818 GND.n4216 240.244
R18030 GND.n7818 GND.n4222 240.244
R18031 GND.n7810 GND.n4222 240.244
R18032 GND.n7810 GND.n4236 240.244
R18033 GND.n7806 GND.n4236 240.244
R18034 GND.n7806 GND.n4242 240.244
R18035 GND.n7798 GND.n4242 240.244
R18036 GND.n7798 GND.n4254 240.244
R18037 GND.n7794 GND.n4254 240.244
R18038 GND.n7794 GND.n4260 240.244
R18039 GND.n4283 GND.n4260 240.244
R18040 GND.n7779 GND.n4283 240.244
R18041 GND.n7779 GND.n4284 240.244
R18042 GND.n7775 GND.n4284 240.244
R18043 GND.n7775 GND.n4292 240.244
R18044 GND.n7767 GND.n4292 240.244
R18045 GND.n7767 GND.n4319 240.244
R18046 GND.n7763 GND.n4319 240.244
R18047 GND.n7763 GND.n4325 240.244
R18048 GND.n7755 GND.n4325 240.244
R18049 GND.n7755 GND.n4339 240.244
R18050 GND.n7751 GND.n4339 240.244
R18051 GND.n7751 GND.n4345 240.244
R18052 GND.n7743 GND.n4345 240.244
R18053 GND.n7743 GND.n4358 240.244
R18054 GND.n7739 GND.n4358 240.244
R18055 GND.n7739 GND.n4364 240.244
R18056 GND.n4386 GND.n4364 240.244
R18057 GND.n7724 GND.n4386 240.244
R18058 GND.n7724 GND.n4387 240.244
R18059 GND.n7720 GND.n4387 240.244
R18060 GND.n7720 GND.n4395 240.244
R18061 GND.n7710 GND.n4395 240.244
R18062 GND.n7710 GND.n4407 240.244
R18063 GND.n7706 GND.n4407 240.244
R18064 GND.n7706 GND.n4413 240.244
R18065 GND.n7696 GND.n4413 240.244
R18066 GND.n7696 GND.n4425 240.244
R18067 GND.n7692 GND.n4425 240.244
R18068 GND.n7692 GND.n4431 240.244
R18069 GND.n7682 GND.n4431 240.244
R18070 GND.n7682 GND.n4442 240.244
R18071 GND.n7678 GND.n4442 240.244
R18072 GND.n7678 GND.n4448 240.244
R18073 GND.n4517 GND.n4448 240.244
R18074 GND.n7663 GND.n4517 240.244
R18075 GND.n7663 GND.n4518 240.244
R18076 GND.n7659 GND.n4518 240.244
R18077 GND.n7659 GND.n4526 240.244
R18078 GND.n7654 GND.n4526 240.244
R18079 GND.n7654 GND.n4561 240.244
R18080 GND.n7650 GND.n4561 240.244
R18081 GND.n7650 GND.n4567 240.244
R18082 GND.n6540 GND.n4567 240.244
R18083 GND.n6546 GND.n6540 240.244
R18084 GND.n6547 GND.n6546 240.244
R18085 GND.n6548 GND.n6547 240.244
R18086 GND.n6548 GND.n6536 240.244
R18087 GND.n6554 GND.n6536 240.244
R18088 GND.n6555 GND.n6554 240.244
R18089 GND.n6556 GND.n6555 240.244
R18090 GND.n6556 GND.n6531 240.244
R18091 GND.n6731 GND.n6531 240.244
R18092 GND.n6731 GND.n6532 240.244
R18093 GND.n6727 GND.n6532 240.244
R18094 GND.n6727 GND.n6726 240.244
R18095 GND.n6726 GND.n6725 240.244
R18096 GND.n6725 GND.n6564 240.244
R18097 GND.n6721 GND.n6564 240.244
R18098 GND.n6721 GND.n6720 240.244
R18099 GND.n6720 GND.n6719 240.244
R18100 GND.n6719 GND.n6570 240.244
R18101 GND.n6715 GND.n6570 240.244
R18102 GND.n6715 GND.n6714 240.244
R18103 GND.n6714 GND.n6713 240.244
R18104 GND.n6713 GND.n6576 240.244
R18105 GND.n6709 GND.n6576 240.244
R18106 GND.n6709 GND.n6708 240.244
R18107 GND.n6708 GND.n6707 240.244
R18108 GND.n6707 GND.n6582 240.244
R18109 GND.n6703 GND.n6582 240.244
R18110 GND.n6703 GND.n6702 240.244
R18111 GND.n6702 GND.n6701 240.244
R18112 GND.n6701 GND.n6588 240.244
R18113 GND.n6697 GND.n6588 240.244
R18114 GND.n6697 GND.n6696 240.244
R18115 GND.n6696 GND.n6695 240.244
R18116 GND.n6695 GND.n6594 240.244
R18117 GND.n6691 GND.n6594 240.244
R18118 GND.n6691 GND.n6690 240.244
R18119 GND.n6690 GND.n6689 240.244
R18120 GND.n6689 GND.n6600 240.244
R18121 GND.n6685 GND.n6600 240.244
R18122 GND.n6685 GND.n6684 240.244
R18123 GND.n6684 GND.n6683 240.244
R18124 GND.n6683 GND.n6606 240.244
R18125 GND.n6679 GND.n6606 240.244
R18126 GND.n6679 GND.n6678 240.244
R18127 GND.n6678 GND.n6677 240.244
R18128 GND.n6677 GND.n6612 240.244
R18129 GND.n6673 GND.n6612 240.244
R18130 GND.n6673 GND.n6672 240.244
R18131 GND.n6672 GND.n6671 240.244
R18132 GND.n6671 GND.n6618 240.244
R18133 GND.n6667 GND.n6618 240.244
R18134 GND.n6667 GND.n6666 240.244
R18135 GND.n6666 GND.n6665 240.244
R18136 GND.n6665 GND.n6624 240.244
R18137 GND.n6661 GND.n6624 240.244
R18138 GND.n6661 GND.n6660 240.244
R18139 GND.n6660 GND.n6659 240.244
R18140 GND.n6659 GND.n6630 240.244
R18141 GND.n6655 GND.n6630 240.244
R18142 GND.n6655 GND.n6654 240.244
R18143 GND.n6654 GND.n6653 240.244
R18144 GND.n6653 GND.n6636 240.244
R18145 GND.n6649 GND.n6636 240.244
R18146 GND.n6649 GND.n6648 240.244
R18147 GND.n6648 GND.n6647 240.244
R18148 GND.n6647 GND.n6643 240.244
R18149 GND.n6643 GND.n6260 240.244
R18150 GND.n7331 GND.n6260 240.244
R18151 GND.n7331 GND.n6261 240.244
R18152 GND.n7326 GND.n6261 240.244
R18153 GND.n7326 GND.n7325 240.244
R18154 GND.n7325 GND.n6264 240.244
R18155 GND.n7320 GND.n6264 240.244
R18156 GND.n7320 GND.n6266 240.244
R18157 GND.n6279 GND.n6266 240.244
R18158 GND.n7310 GND.n6279 240.244
R18159 GND.n7310 GND.n6280 240.244
R18160 GND.n7306 GND.n6280 240.244
R18161 GND.n7306 GND.n7305 240.244
R18162 GND.n7305 GND.n7304 240.244
R18163 GND.n7304 GND.n6287 240.244
R18164 GND.n7300 GND.n6287 240.244
R18165 GND.n7300 GND.n7299 240.244
R18166 GND.n7299 GND.n7298 240.244
R18167 GND.n7298 GND.n6293 240.244
R18168 GND.n7294 GND.n6293 240.244
R18169 GND.n7294 GND.n7293 240.244
R18170 GND.n7293 GND.n7292 240.244
R18171 GND.n7292 GND.n6299 240.244
R18172 GND.n7288 GND.n6299 240.244
R18173 GND.n7288 GND.n7287 240.244
R18174 GND.n7287 GND.n7286 240.244
R18175 GND.n7286 GND.n6305 240.244
R18176 GND.n7282 GND.n6305 240.244
R18177 GND.n7282 GND.n7281 240.244
R18178 GND.n7281 GND.n7280 240.244
R18179 GND.n7280 GND.n6311 240.244
R18180 GND.n7276 GND.n6311 240.244
R18181 GND.n7276 GND.n7275 240.244
R18182 GND.n7275 GND.n7274 240.244
R18183 GND.n7274 GND.n6317 240.244
R18184 GND.n7270 GND.n6317 240.244
R18185 GND.n7270 GND.n6433 240.244
R18186 GND.n6433 GND.n6432 240.244
R18187 GND.n6432 GND.n6323 240.244
R18188 GND.n6428 GND.n6323 240.244
R18189 GND.n6428 GND.n6427 240.244
R18190 GND.n6427 GND.n6426 240.244
R18191 GND.n6426 GND.n6329 240.244
R18192 GND.n6422 GND.n6329 240.244
R18193 GND.n6422 GND.n6421 240.244
R18194 GND.n6421 GND.n6420 240.244
R18195 GND.n6420 GND.n6335 240.244
R18196 GND.n6416 GND.n6335 240.244
R18197 GND.n6416 GND.n6415 240.244
R18198 GND.n6415 GND.n6414 240.244
R18199 GND.n6414 GND.n6341 240.244
R18200 GND.n6410 GND.n6341 240.244
R18201 GND.n6410 GND.n6409 240.244
R18202 GND.n6409 GND.n6408 240.244
R18203 GND.n6408 GND.n6347 240.244
R18204 GND.n6404 GND.n6347 240.244
R18205 GND.n6404 GND.n6403 240.244
R18206 GND.n6403 GND.n6402 240.244
R18207 GND.n6402 GND.n6353 240.244
R18208 GND.n6398 GND.n6353 240.244
R18209 GND.n6398 GND.n6397 240.244
R18210 GND.n6397 GND.n6396 240.244
R18211 GND.n6396 GND.n6359 240.244
R18212 GND.n6392 GND.n6359 240.244
R18213 GND.n6392 GND.n6391 240.244
R18214 GND.n6391 GND.n6390 240.244
R18215 GND.n6390 GND.n6365 240.244
R18216 GND.n6386 GND.n6365 240.244
R18217 GND.n6386 GND.n6385 240.244
R18218 GND.n6385 GND.n6384 240.244
R18219 GND.n6384 GND.n6371 240.244
R18220 GND.n6380 GND.n6371 240.244
R18221 GND.n6380 GND.n6379 240.244
R18222 GND.n6379 GND.n462 240.244
R18223 GND.n10645 GND.n462 240.244
R18224 GND.n10645 GND.n463 240.244
R18225 GND.n10641 GND.n463 240.244
R18226 GND.n10641 GND.n469 240.244
R18227 GND.n10637 GND.n469 240.244
R18228 GND.n10637 GND.n471 240.244
R18229 GND.n10633 GND.n471 240.244
R18230 GND.n10633 GND.n477 240.244
R18231 GND.n10629 GND.n477 240.244
R18232 GND.n10629 GND.n479 240.244
R18233 GND.n10625 GND.n479 240.244
R18234 GND.n10625 GND.n485 240.244
R18235 GND.n10621 GND.n485 240.244
R18236 GND.n10621 GND.n487 240.244
R18237 GND.n10617 GND.n487 240.244
R18238 GND.n10617 GND.n493 240.244
R18239 GND.n10613 GND.n493 240.244
R18240 GND.n10613 GND.n495 240.244
R18241 GND.n10609 GND.n495 240.244
R18242 GND.n10609 GND.n501 240.244
R18243 GND.n10605 GND.n501 240.244
R18244 GND.n10605 GND.n503 240.244
R18245 GND.n10601 GND.n503 240.244
R18246 GND.n10601 GND.n509 240.244
R18247 GND.n10597 GND.n509 240.244
R18248 GND.n10597 GND.n511 240.244
R18249 GND.n10593 GND.n511 240.244
R18250 GND.n10593 GND.n517 240.244
R18251 GND.n10589 GND.n517 240.244
R18252 GND.n10589 GND.n519 240.244
R18253 GND.n10585 GND.n519 240.244
R18254 GND.n10585 GND.n525 240.244
R18255 GND.n10581 GND.n525 240.244
R18256 GND.n10581 GND.n527 240.244
R18257 GND.n10577 GND.n527 240.244
R18258 GND.n10577 GND.n533 240.244
R18259 GND.n10573 GND.n533 240.244
R18260 GND.n10573 GND.n535 240.244
R18261 GND.n10569 GND.n535 240.244
R18262 GND.n10569 GND.n541 240.244
R18263 GND.n10565 GND.n541 240.244
R18264 GND.n10565 GND.n543 240.244
R18265 GND.n10561 GND.n543 240.244
R18266 GND.n10561 GND.n549 240.244
R18267 GND.n10557 GND.n549 240.244
R18268 GND.n10557 GND.n551 240.244
R18269 GND.n10553 GND.n551 240.244
R18270 GND.n10553 GND.n557 240.244
R18271 GND.n10549 GND.n557 240.244
R18272 GND.n10549 GND.n559 240.244
R18273 GND.n10545 GND.n559 240.244
R18274 GND.n10545 GND.n565 240.244
R18275 GND.n10541 GND.n565 240.244
R18276 GND.n10541 GND.n567 240.244
R18277 GND.n10537 GND.n567 240.244
R18278 GND.n10537 GND.n573 240.244
R18279 GND.n9045 GND.n1462 240.244
R18280 GND.n9045 GND.n1465 240.244
R18281 GND.n9041 GND.n1465 240.244
R18282 GND.n9041 GND.n1467 240.244
R18283 GND.n9037 GND.n1467 240.244
R18284 GND.n9037 GND.n1473 240.244
R18285 GND.n9033 GND.n1473 240.244
R18286 GND.n9033 GND.n1475 240.244
R18287 GND.n9029 GND.n1475 240.244
R18288 GND.n9029 GND.n1481 240.244
R18289 GND.n9025 GND.n1481 240.244
R18290 GND.n9025 GND.n1483 240.244
R18291 GND.n9021 GND.n1483 240.244
R18292 GND.n9021 GND.n1489 240.244
R18293 GND.n9017 GND.n1489 240.244
R18294 GND.n9017 GND.n1491 240.244
R18295 GND.n9013 GND.n1491 240.244
R18296 GND.n9013 GND.n1497 240.244
R18297 GND.n9009 GND.n1497 240.244
R18298 GND.n9009 GND.n1499 240.244
R18299 GND.n9005 GND.n1499 240.244
R18300 GND.n9005 GND.n1505 240.244
R18301 GND.n9001 GND.n1505 240.244
R18302 GND.n9001 GND.n1507 240.244
R18303 GND.n8997 GND.n1507 240.244
R18304 GND.n8997 GND.n1513 240.244
R18305 GND.n8993 GND.n1513 240.244
R18306 GND.n8993 GND.n1515 240.244
R18307 GND.n8989 GND.n1515 240.244
R18308 GND.n8989 GND.n1521 240.244
R18309 GND.n8985 GND.n1521 240.244
R18310 GND.n8985 GND.n1523 240.244
R18311 GND.n8981 GND.n1523 240.244
R18312 GND.n8981 GND.n1529 240.244
R18313 GND.n8977 GND.n1529 240.244
R18314 GND.n8977 GND.n1531 240.244
R18315 GND.n8973 GND.n1531 240.244
R18316 GND.n8973 GND.n1537 240.244
R18317 GND.n8969 GND.n1537 240.244
R18318 GND.n8969 GND.n1539 240.244
R18319 GND.n8965 GND.n1539 240.244
R18320 GND.n8965 GND.n1545 240.244
R18321 GND.n8961 GND.n1545 240.244
R18322 GND.n8961 GND.n1547 240.244
R18323 GND.n8957 GND.n1547 240.244
R18324 GND.n8957 GND.n1553 240.244
R18325 GND.n8953 GND.n1553 240.244
R18326 GND.n8953 GND.n1555 240.244
R18327 GND.n8949 GND.n1555 240.244
R18328 GND.n8949 GND.n1561 240.244
R18329 GND.n8945 GND.n1561 240.244
R18330 GND.n8945 GND.n1563 240.244
R18331 GND.n8941 GND.n1563 240.244
R18332 GND.n8941 GND.n1569 240.244
R18333 GND.n8937 GND.n1569 240.244
R18334 GND.n8937 GND.n1571 240.244
R18335 GND.n8933 GND.n1571 240.244
R18336 GND.n8933 GND.n1577 240.244
R18337 GND.n8699 GND.n1799 240.244
R18338 GND.n1854 GND.n1799 240.244
R18339 GND.n1854 GND.n1821 240.244
R18340 GND.n1840 GND.n1821 240.244
R18341 GND.n8683 GND.n1840 240.244
R18342 GND.n8683 GND.n1841 240.244
R18343 GND.n2966 GND.n1841 240.244
R18344 GND.n2966 GND.n2900 240.244
R18345 GND.n3170 GND.n2900 240.244
R18346 GND.n3174 GND.n3170 240.244
R18347 GND.n3174 GND.n3172 240.244
R18348 GND.n3172 GND.n2889 240.244
R18349 GND.n2889 GND.n2877 240.244
R18350 GND.n3195 GND.n2877 240.244
R18351 GND.n3199 GND.n3195 240.244
R18352 GND.n3199 GND.n3198 240.244
R18353 GND.n3198 GND.n2866 240.244
R18354 GND.n2866 GND.n2856 240.244
R18355 GND.n3220 GND.n2856 240.244
R18356 GND.n3223 GND.n3220 240.244
R18357 GND.n3223 GND.n3222 240.244
R18358 GND.n3222 GND.n2843 240.244
R18359 GND.n2843 GND.n2831 240.244
R18360 GND.n3244 GND.n2831 240.244
R18361 GND.n3248 GND.n3244 240.244
R18362 GND.n3248 GND.n3247 240.244
R18363 GND.n3247 GND.n2819 240.244
R18364 GND.n2819 GND.n2809 240.244
R18365 GND.n3269 GND.n2809 240.244
R18366 GND.n3273 GND.n3269 240.244
R18367 GND.n3273 GND.n3271 240.244
R18368 GND.n3271 GND.n2798 240.244
R18369 GND.n2798 GND.n2786 240.244
R18370 GND.n3294 GND.n2786 240.244
R18371 GND.n3298 GND.n3294 240.244
R18372 GND.n3298 GND.n3297 240.244
R18373 GND.n3297 GND.n2775 240.244
R18374 GND.n2775 GND.n2765 240.244
R18375 GND.n3319 GND.n2765 240.244
R18376 GND.n3322 GND.n3319 240.244
R18377 GND.n3322 GND.n3321 240.244
R18378 GND.n3321 GND.n2752 240.244
R18379 GND.n2752 GND.n2740 240.244
R18380 GND.n3343 GND.n2740 240.244
R18381 GND.n3347 GND.n3343 240.244
R18382 GND.n3347 GND.n3346 240.244
R18383 GND.n3346 GND.n2728 240.244
R18384 GND.n2728 GND.n2718 240.244
R18385 GND.n3368 GND.n2718 240.244
R18386 GND.n3372 GND.n3368 240.244
R18387 GND.n3372 GND.n3370 240.244
R18388 GND.n3370 GND.n2707 240.244
R18389 GND.n2707 GND.n2695 240.244
R18390 GND.n3393 GND.n2695 240.244
R18391 GND.n3397 GND.n3393 240.244
R18392 GND.n3397 GND.n3396 240.244
R18393 GND.n3396 GND.n2684 240.244
R18394 GND.n2684 GND.n2674 240.244
R18395 GND.n3418 GND.n2674 240.244
R18396 GND.n3421 GND.n3418 240.244
R18397 GND.n3421 GND.n3420 240.244
R18398 GND.n3420 GND.n2663 240.244
R18399 GND.n2663 GND.n2505 240.244
R18400 GND.n3489 GND.n2505 240.244
R18401 GND.n3489 GND.n3488 240.244
R18402 GND.n3488 GND.n2507 240.244
R18403 GND.n2520 GND.n2507 240.244
R18404 GND.n2521 GND.n2520 240.244
R18405 GND.n3472 GND.n2521 240.244
R18406 GND.n3472 GND.n3471 240.244
R18407 GND.n3471 GND.n2528 240.244
R18408 GND.n3459 GND.n2528 240.244
R18409 GND.n3460 GND.n3459 240.244
R18410 GND.n3460 GND.n2486 240.244
R18411 GND.n2486 GND.n2475 240.244
R18412 GND.n3511 GND.n2475 240.244
R18413 GND.n3515 GND.n3511 240.244
R18414 GND.n3515 GND.n3514 240.244
R18415 GND.n3514 GND.n2463 240.244
R18416 GND.n2463 GND.n2454 240.244
R18417 GND.n3537 GND.n2454 240.244
R18418 GND.n3541 GND.n3537 240.244
R18419 GND.n3541 GND.n3539 240.244
R18420 GND.n3539 GND.n2443 240.244
R18421 GND.n2443 GND.n2432 240.244
R18422 GND.n3563 GND.n2432 240.244
R18423 GND.n3567 GND.n3563 240.244
R18424 GND.n3567 GND.n3566 240.244
R18425 GND.n3566 GND.n2421 240.244
R18426 GND.n2421 GND.n2412 240.244
R18427 GND.n3589 GND.n2412 240.244
R18428 GND.n3592 GND.n3589 240.244
R18429 GND.n3592 GND.n3591 240.244
R18430 GND.n3591 GND.n2399 240.244
R18431 GND.n2399 GND.n2388 240.244
R18432 GND.n3614 GND.n2388 240.244
R18433 GND.n3618 GND.n3614 240.244
R18434 GND.n3618 GND.n3617 240.244
R18435 GND.n3617 GND.n2378 240.244
R18436 GND.n2378 GND.n2370 240.244
R18437 GND.n3640 GND.n2370 240.244
R18438 GND.n3644 GND.n3640 240.244
R18439 GND.n3644 GND.n3642 240.244
R18440 GND.n3642 GND.n2359 240.244
R18441 GND.n2359 GND.n2348 240.244
R18442 GND.n3666 GND.n2348 240.244
R18443 GND.n3670 GND.n3666 240.244
R18444 GND.n3670 GND.n3669 240.244
R18445 GND.n3669 GND.n2338 240.244
R18446 GND.n2338 GND.n2337 240.244
R18447 GND.n2337 GND.n2321 240.244
R18448 GND.n8181 GND.n2321 240.244
R18449 GND.n8181 GND.n8180 240.244
R18450 GND.n8180 GND.n2309 240.244
R18451 GND.n2309 GND.n2299 240.244
R18452 GND.n8203 GND.n2299 240.244
R18453 GND.n8207 GND.n8203 240.244
R18454 GND.n8207 GND.n8206 240.244
R18455 GND.n8206 GND.n2287 240.244
R18456 GND.n2287 GND.n2278 240.244
R18457 GND.n8229 GND.n2278 240.244
R18458 GND.n8233 GND.n8229 240.244
R18459 GND.n8233 GND.n8231 240.244
R18460 GND.n8231 GND.n2267 240.244
R18461 GND.n2267 GND.n2256 240.244
R18462 GND.n8255 GND.n2256 240.244
R18463 GND.n8259 GND.n8255 240.244
R18464 GND.n8259 GND.n8258 240.244
R18465 GND.n8258 GND.n2245 240.244
R18466 GND.n2245 GND.n2236 240.244
R18467 GND.n8281 GND.n2236 240.244
R18468 GND.n8284 GND.n8281 240.244
R18469 GND.n8284 GND.n8283 240.244
R18470 GND.n8283 GND.n2225 240.244
R18471 GND.n2225 GND.n2223 240.244
R18472 GND.n2223 GND.n2129 240.244
R18473 GND.n8479 GND.n2129 240.244
R18474 GND.n2922 GND.n2921 240.244
R18475 GND.n2928 GND.n2927 240.244
R18476 GND.n2931 GND.n2930 240.244
R18477 GND.n2938 GND.n2937 240.244
R18478 GND.n2941 GND.n2940 240.244
R18479 GND.n2917 GND.n2913 240.244
R18480 GND.n2954 GND.n1804 240.244
R18481 GND.n2955 GND.n2954 240.244
R18482 GND.n2955 GND.n1819 240.244
R18483 GND.n2908 GND.n1819 240.244
R18484 GND.n2908 GND.n1838 240.244
R18485 GND.n2963 GND.n1838 240.244
R18486 GND.n3161 GND.n2963 240.244
R18487 GND.n3161 GND.n2902 240.244
R18488 GND.n3168 GND.n2902 240.244
R18489 GND.n3168 GND.n2898 240.244
R18490 GND.n2898 GND.n2885 240.244
R18491 GND.n3186 GND.n2885 240.244
R18492 GND.n3186 GND.n2880 240.244
R18493 GND.n3193 GND.n2880 240.244
R18494 GND.n3193 GND.n2875 240.244
R18495 GND.n2875 GND.n2863 240.244
R18496 GND.n3211 GND.n2863 240.244
R18497 GND.n3211 GND.n2858 240.244
R18498 GND.n3218 GND.n2858 240.244
R18499 GND.n3218 GND.n2853 240.244
R18500 GND.n2853 GND.n2839 240.244
R18501 GND.n3235 GND.n2839 240.244
R18502 GND.n3235 GND.n2834 240.244
R18503 GND.n3242 GND.n2834 240.244
R18504 GND.n3242 GND.n2829 240.244
R18505 GND.n2829 GND.n2816 240.244
R18506 GND.n3260 GND.n2816 240.244
R18507 GND.n3260 GND.n2811 240.244
R18508 GND.n3267 GND.n2811 240.244
R18509 GND.n3267 GND.n2807 240.244
R18510 GND.n2807 GND.n2794 240.244
R18511 GND.n3285 GND.n2794 240.244
R18512 GND.n3285 GND.n2789 240.244
R18513 GND.n3292 GND.n2789 240.244
R18514 GND.n3292 GND.n2784 240.244
R18515 GND.n2784 GND.n2772 240.244
R18516 GND.n3310 GND.n2772 240.244
R18517 GND.n3310 GND.n2767 240.244
R18518 GND.n3317 GND.n2767 240.244
R18519 GND.n3317 GND.n2762 240.244
R18520 GND.n2762 GND.n2748 240.244
R18521 GND.n3334 GND.n2748 240.244
R18522 GND.n3334 GND.n2743 240.244
R18523 GND.n3341 GND.n2743 240.244
R18524 GND.n3341 GND.n2738 240.244
R18525 GND.n2738 GND.n2725 240.244
R18526 GND.n3359 GND.n2725 240.244
R18527 GND.n3359 GND.n2720 240.244
R18528 GND.n3366 GND.n2720 240.244
R18529 GND.n3366 GND.n2716 240.244
R18530 GND.n2716 GND.n2703 240.244
R18531 GND.n3384 GND.n2703 240.244
R18532 GND.n3384 GND.n2698 240.244
R18533 GND.n3391 GND.n2698 240.244
R18534 GND.n3391 GND.n2693 240.244
R18535 GND.n2693 GND.n2681 240.244
R18536 GND.n3409 GND.n2681 240.244
R18537 GND.n3409 GND.n2676 240.244
R18538 GND.n3416 GND.n2676 240.244
R18539 GND.n3416 GND.n2671 240.244
R18540 GND.n2671 GND.n2659 240.244
R18541 GND.n3431 GND.n2659 240.244
R18542 GND.n3431 GND.n2660 240.244
R18543 GND.n2660 GND.n2503 240.244
R18544 GND.n2508 GND.n2503 240.244
R18545 GND.n3439 GND.n2508 240.244
R18546 GND.n3439 GND.n3438 240.244
R18547 GND.n3438 GND.n2518 240.244
R18548 GND.n2526 GND.n2518 240.244
R18549 GND.n2530 GND.n2526 240.244
R18550 GND.n2651 GND.n2530 240.244
R18551 GND.n3452 GND.n2651 240.244
R18552 GND.n3452 GND.n2482 240.244
R18553 GND.n3501 GND.n2482 240.244
R18554 GND.n3501 GND.n2478 240.244
R18555 GND.n3509 GND.n2478 240.244
R18556 GND.n3509 GND.n2473 240.244
R18557 GND.n2473 GND.n2460 240.244
R18558 GND.n3527 GND.n2460 240.244
R18559 GND.n3527 GND.n2456 240.244
R18560 GND.n3535 GND.n2456 240.244
R18561 GND.n3535 GND.n2452 240.244
R18562 GND.n2452 GND.n2439 240.244
R18563 GND.n3553 GND.n2439 240.244
R18564 GND.n3553 GND.n2435 240.244
R18565 GND.n3561 GND.n2435 240.244
R18566 GND.n3561 GND.n2430 240.244
R18567 GND.n2430 GND.n2418 240.244
R18568 GND.n3579 GND.n2418 240.244
R18569 GND.n3579 GND.n2414 240.244
R18570 GND.n3587 GND.n2414 240.244
R18571 GND.n3587 GND.n2409 240.244
R18572 GND.n2409 GND.n2395 240.244
R18573 GND.n3604 GND.n2395 240.244
R18574 GND.n3604 GND.n2391 240.244
R18575 GND.n3612 GND.n2391 240.244
R18576 GND.n3612 GND.n2386 240.244
R18577 GND.n2386 GND.n2375 240.244
R18578 GND.n3630 GND.n2375 240.244
R18579 GND.n3630 GND.n2371 240.244
R18580 GND.n3638 GND.n2371 240.244
R18581 GND.n3638 GND.n2368 240.244
R18582 GND.n2368 GND.n2355 240.244
R18583 GND.n3656 GND.n2355 240.244
R18584 GND.n3656 GND.n2351 240.244
R18585 GND.n3664 GND.n2351 240.244
R18586 GND.n3664 GND.n2346 240.244
R18587 GND.n2346 GND.n2333 240.244
R18588 GND.n3682 GND.n2333 240.244
R18589 GND.n3682 GND.n2329 240.244
R18590 GND.n3690 GND.n2329 240.244
R18591 GND.n3690 GND.n2319 240.244
R18592 GND.n2319 GND.n2306 240.244
R18593 GND.n8193 GND.n2306 240.244
R18594 GND.n8193 GND.n2302 240.244
R18595 GND.n8201 GND.n2302 240.244
R18596 GND.n8201 GND.n2297 240.244
R18597 GND.n2297 GND.n2284 240.244
R18598 GND.n8219 GND.n2284 240.244
R18599 GND.n8219 GND.n2280 240.244
R18600 GND.n8227 GND.n2280 240.244
R18601 GND.n8227 GND.n2276 240.244
R18602 GND.n2276 GND.n2263 240.244
R18603 GND.n8245 GND.n2263 240.244
R18604 GND.n8245 GND.n2259 240.244
R18605 GND.n8253 GND.n2259 240.244
R18606 GND.n8253 GND.n2254 240.244
R18607 GND.n2254 GND.n2242 240.244
R18608 GND.n8271 GND.n2242 240.244
R18609 GND.n8271 GND.n2238 240.244
R18610 GND.n8279 GND.n2238 240.244
R18611 GND.n8279 GND.n2233 240.244
R18612 GND.n2233 GND.n2219 240.244
R18613 GND.n8295 GND.n2219 240.244
R18614 GND.n8295 GND.n2215 240.244
R18615 GND.n8303 GND.n2215 240.244
R18616 GND.n8303 GND.n2127 240.244
R18617 GND.n2133 GND.n2132 240.244
R18618 GND.n2135 GND.n2134 240.244
R18619 GND.n2137 GND.n2136 240.244
R18620 GND.n2139 GND.n2138 240.244
R18621 GND.n2141 GND.n2140 240.244
R18622 GND.n8459 GND.n2142 240.244
R18623 GND.n8013 GND.t113 233.655
R18624 GND.n5860 GND.t145 233.655
R18625 GND.n2914 GND.t104 225.825
R18626 GND.n8332 GND.t98 225.825
R18627 GND.n8382 GND.t95 225.825
R18628 GND.n8406 GND.t136 225.825
R18629 GND.n2183 GND.t142 225.825
R18630 GND.n4620 GND.t60 225.825
R18631 GND.n4794 GND.t117 225.825
R18632 GND.n4810 GND.t53 225.825
R18633 GND.n4828 GND.t92 225.825
R18634 GND.n10784 GND.t73 225.825
R18635 GND.n10765 GND.t77 225.825
R18636 GND.n10748 GND.t133 225.825
R18637 GND.n10732 GND.t80 225.825
R18638 GND.n456 GND.t101 225.825
R18639 GND.n5886 GND.t120 225.825
R18640 GND.n1743 GND.t126 225.825
R18641 GND.n1759 GND.t69 225.825
R18642 GND.n1776 GND.t123 225.825
R18643 GND.n1794 GND.t83 225.825
R18644 GND.n2143 GND.t45 225.825
R18645 GND.n2182 GND.n2160 199.319
R18646 GND.n3759 GND.n3757 186.49
R18647 GND.n4642 GND.n4640 186.49
R18648 GND.n4810 GND.t56 185.352
R18649 GND.n10784 GND.t75 185.352
R18650 GND.n2914 GND.t106 175.752
R18651 GND.n8332 GND.t99 175.752
R18652 GND.n8382 GND.t96 175.752
R18653 GND.n8406 GND.t137 175.752
R18654 GND.n2183 GND.t143 175.752
R18655 GND.n4620 GND.t62 175.752
R18656 GND.n4794 GND.t119 175.752
R18657 GND.n4828 GND.t94 175.752
R18658 GND.n10765 GND.t78 175.752
R18659 GND.n10748 GND.t134 175.752
R18660 GND.n10732 GND.t81 175.752
R18661 GND.n456 GND.t102 175.752
R18662 GND.n5886 GND.t122 175.752
R18663 GND.n1743 GND.t128 175.752
R18664 GND.n1759 GND.t72 175.752
R18665 GND.n1776 GND.t125 175.752
R18666 GND.n1794 GND.t85 175.752
R18667 GND.n2143 GND.t47 175.752
R18668 GND.n4731 GND.n4730 163.367
R18669 GND.n4735 GND.n4734 163.367
R18670 GND.n4739 GND.n4738 163.367
R18671 GND.n4743 GND.n4742 163.367
R18672 GND.n4747 GND.n4746 163.367
R18673 GND.n4751 GND.n4750 163.367
R18674 GND.n4755 GND.n4754 163.367
R18675 GND.n4759 GND.n4758 163.367
R18676 GND.n4763 GND.n4762 163.367
R18677 GND.n4767 GND.n4766 163.367
R18678 GND.n4771 GND.n4770 163.367
R18679 GND.n4775 GND.n4774 163.367
R18680 GND.n4779 GND.n4778 163.367
R18681 GND.n4784 GND.n4783 163.367
R18682 GND.n4788 GND.n4787 163.367
R18683 GND.n4658 GND.n4657 163.367
R18684 GND.n4662 GND.n4661 163.367
R18685 GND.n4667 GND.n4666 163.367
R18686 GND.n4671 GND.n4670 163.367
R18687 GND.n4675 GND.n4674 163.367
R18688 GND.n4679 GND.n4678 163.367
R18689 GND.n4683 GND.n4682 163.367
R18690 GND.n4687 GND.n4686 163.367
R18691 GND.n4691 GND.n4690 163.367
R18692 GND.n4695 GND.n4694 163.367
R18693 GND.n4699 GND.n4698 163.367
R18694 GND.n4703 GND.n4702 163.367
R18695 GND.n4707 GND.n4706 163.367
R18696 GND.n4711 GND.n4710 163.367
R18697 GND.n4715 GND.n4714 163.367
R18698 GND.n5206 GND.n3750 163.367
R18699 GND.n5206 GND.n3771 163.367
R18700 GND.n5210 GND.n3771 163.367
R18701 GND.n5215 GND.n5210 163.367
R18702 GND.n5216 GND.n5215 163.367
R18703 GND.n5216 GND.n3781 163.367
R18704 GND.n5219 GND.n3781 163.367
R18705 GND.n5219 GND.n3787 163.367
R18706 GND.n5223 GND.n3787 163.367
R18707 GND.n5228 GND.n5223 163.367
R18708 GND.n5229 GND.n5228 163.367
R18709 GND.n5229 GND.n3797 163.367
R18710 GND.n5232 GND.n3797 163.367
R18711 GND.n5232 GND.n3805 163.367
R18712 GND.n5236 GND.n3805 163.367
R18713 GND.n5241 GND.n5236 163.367
R18714 GND.n5242 GND.n5241 163.367
R18715 GND.n5242 GND.n3815 163.367
R18716 GND.n5245 GND.n3815 163.367
R18717 GND.n5245 GND.n3823 163.367
R18718 GND.n5249 GND.n3823 163.367
R18719 GND.n5254 GND.n5249 163.367
R18720 GND.n5255 GND.n5254 163.367
R18721 GND.n5255 GND.n3833 163.367
R18722 GND.n5258 GND.n3833 163.367
R18723 GND.n5258 GND.n3841 163.367
R18724 GND.n5036 GND.n3841 163.367
R18725 GND.n5304 GND.n5036 163.367
R18726 GND.n5304 GND.n5037 163.367
R18727 GND.n5300 GND.n5037 163.367
R18728 GND.n5300 GND.n5299 163.367
R18729 GND.n5299 GND.n3885 163.367
R18730 GND.n5295 GND.n3885 163.367
R18731 GND.n5295 GND.n5294 163.367
R18732 GND.n5294 GND.n5293 163.367
R18733 GND.n5293 GND.n5263 163.367
R18734 GND.n5263 GND.n5031 163.367
R18735 GND.n5288 GND.n5031 163.367
R18736 GND.n5288 GND.n5020 163.367
R18737 GND.n5285 GND.n5020 163.367
R18738 GND.n5285 GND.n5284 163.367
R18739 GND.n5284 GND.n5015 163.367
R18740 GND.n5280 GND.n5015 163.367
R18741 GND.n5280 GND.n5279 163.367
R18742 GND.n5279 GND.n5011 163.367
R18743 GND.n5275 GND.n5011 163.367
R18744 GND.n5275 GND.n5274 163.367
R18745 GND.n5274 GND.n5006 163.367
R18746 GND.n5270 GND.n5006 163.367
R18747 GND.n5270 GND.n5269 163.367
R18748 GND.n5269 GND.n5002 163.367
R18749 GND.n5265 GND.n5002 163.367
R18750 GND.n5265 GND.n4996 163.367
R18751 GND.n5422 GND.n4996 163.367
R18752 GND.n5423 GND.n5422 163.367
R18753 GND.n5423 GND.n4993 163.367
R18754 GND.n5429 GND.n4993 163.367
R18755 GND.n5429 GND.n4994 163.367
R18756 GND.n4994 GND.n4986 163.367
R18757 GND.n5440 GND.n4986 163.367
R18758 GND.n5441 GND.n5440 163.367
R18759 GND.n5441 GND.n4983 163.367
R18760 GND.n5447 GND.n4983 163.367
R18761 GND.n5447 GND.n4984 163.367
R18762 GND.n4984 GND.n4977 163.367
R18763 GND.n5458 GND.n4977 163.367
R18764 GND.n5459 GND.n5458 163.367
R18765 GND.n5459 GND.n4974 163.367
R18766 GND.n5465 GND.n4974 163.367
R18767 GND.n5465 GND.n4975 163.367
R18768 GND.n4975 GND.n4967 163.367
R18769 GND.n5476 GND.n4967 163.367
R18770 GND.n5477 GND.n5476 163.367
R18771 GND.n5477 GND.n4964 163.367
R18772 GND.n5489 GND.n4964 163.367
R18773 GND.n5489 GND.n4965 163.367
R18774 GND.n5485 GND.n4965 163.367
R18775 GND.n5485 GND.n4958 163.367
R18776 GND.n5482 GND.n4958 163.367
R18777 GND.n5482 GND.n5481 163.367
R18778 GND.n5481 GND.n4059 163.367
R18779 GND.n7902 GND.n4059 163.367
R18780 GND.n7902 GND.n4060 163.367
R18781 GND.n7898 GND.n4060 163.367
R18782 GND.n7898 GND.n4063 163.367
R18783 GND.n4072 GND.n4063 163.367
R18784 GND.n5543 GND.n4072 163.367
R18785 GND.n5550 GND.n5543 163.367
R18786 GND.n5550 GND.n5544 163.367
R18787 GND.n5544 GND.n4946 163.367
R18788 GND.n5561 GND.n4946 163.367
R18789 GND.n5562 GND.n5561 163.367
R18790 GND.n5562 GND.n4943 163.367
R18791 GND.n5568 GND.n4943 163.367
R18792 GND.n5568 GND.n4944 163.367
R18793 GND.n4944 GND.n4936 163.367
R18794 GND.n5579 GND.n4936 163.367
R18795 GND.n5580 GND.n5579 163.367
R18796 GND.n5580 GND.n4933 163.367
R18797 GND.n5592 GND.n4933 163.367
R18798 GND.n5592 GND.n4934 163.367
R18799 GND.n5588 GND.n4934 163.367
R18800 GND.n5588 GND.n4927 163.367
R18801 GND.n5585 GND.n4927 163.367
R18802 GND.n5585 GND.n5584 163.367
R18803 GND.n5584 GND.n4164 163.367
R18804 GND.n7847 GND.n4164 163.367
R18805 GND.n7847 GND.n4165 163.367
R18806 GND.n7843 GND.n4165 163.367
R18807 GND.n7843 GND.n4168 163.367
R18808 GND.n4177 GND.n4168 163.367
R18809 GND.n5647 GND.n4177 163.367
R18810 GND.n5654 GND.n5647 163.367
R18811 GND.n5654 GND.n5648 163.367
R18812 GND.n5648 GND.n4914 163.367
R18813 GND.n5665 GND.n4914 163.367
R18814 GND.n5666 GND.n5665 163.367
R18815 GND.n5666 GND.n4911 163.367
R18816 GND.n5672 GND.n4911 163.367
R18817 GND.n5672 GND.n4912 163.367
R18818 GND.n4912 GND.n4903 163.367
R18819 GND.n5684 GND.n4903 163.367
R18820 GND.n5685 GND.n5684 163.367
R18821 GND.n5686 GND.n5685 163.367
R18822 GND.n5686 GND.n4900 163.367
R18823 GND.n5696 GND.n4900 163.367
R18824 GND.n5696 GND.n4901 163.367
R18825 GND.n4901 GND.n4894 163.367
R18826 GND.n5691 GND.n4894 163.367
R18827 GND.n5691 GND.n5690 163.367
R18828 GND.n5690 GND.n4266 163.367
R18829 GND.n7792 GND.n4266 163.367
R18830 GND.n7792 GND.n4267 163.367
R18831 GND.n7788 GND.n4267 163.367
R18832 GND.n7788 GND.n4270 163.367
R18833 GND.n4279 GND.n4270 163.367
R18834 GND.n5744 GND.n4279 163.367
R18835 GND.n5751 GND.n5744 163.367
R18836 GND.n5751 GND.n5745 163.367
R18837 GND.n5745 GND.n4881 163.367
R18838 GND.n5762 GND.n4881 163.367
R18839 GND.n5763 GND.n5762 163.367
R18840 GND.n5763 GND.n4878 163.367
R18841 GND.n5769 GND.n4878 163.367
R18842 GND.n5769 GND.n4879 163.367
R18843 GND.n4879 GND.n4870 163.367
R18844 GND.n5779 GND.n4870 163.367
R18845 GND.n5780 GND.n5779 163.367
R18846 GND.n5781 GND.n5780 163.367
R18847 GND.n5781 GND.n4853 163.367
R18848 GND.n5784 GND.n4853 163.367
R18849 GND.n5784 GND.n4866 163.367
R18850 GND.n5791 GND.n4866 163.367
R18851 GND.n5791 GND.n4868 163.367
R18852 GND.n5787 GND.n4868 163.367
R18853 GND.n5787 GND.n4370 163.367
R18854 GND.n7737 GND.n4370 163.367
R18855 GND.n7737 GND.n4371 163.367
R18856 GND.n7733 GND.n4371 163.367
R18857 GND.n7733 GND.n4374 163.367
R18858 GND.n4383 GND.n4374 163.367
R18859 GND.n4459 GND.n4383 163.367
R18860 GND.n4464 GND.n4459 163.367
R18861 GND.n4465 GND.n4464 163.367
R18862 GND.n4465 GND.n4397 163.367
R18863 GND.n4468 GND.n4397 163.367
R18864 GND.n4468 GND.n4405 163.367
R18865 GND.n4472 GND.n4405 163.367
R18866 GND.n4477 GND.n4472 163.367
R18867 GND.n4478 GND.n4477 163.367
R18868 GND.n4478 GND.n4415 163.367
R18869 GND.n4481 GND.n4415 163.367
R18870 GND.n4481 GND.n4423 163.367
R18871 GND.n4485 GND.n4423 163.367
R18872 GND.n4490 GND.n4485 163.367
R18873 GND.n4491 GND.n4490 163.367
R18874 GND.n4491 GND.n4433 163.367
R18875 GND.n4494 GND.n4433 163.367
R18876 GND.n4494 GND.n4441 163.367
R18877 GND.n4499 GND.n4441 163.367
R18878 GND.n4499 GND.n4452 163.367
R18879 GND.n7676 GND.n4452 163.367
R18880 GND.n7676 GND.n4453 163.367
R18881 GND.n7672 GND.n4453 163.367
R18882 GND.n7672 GND.n4503 163.367
R18883 GND.n4515 GND.n4503 163.367
R18884 GND.n4651 GND.n4515 163.367
R18885 GND.n4721 GND.n4651 163.367
R18886 GND.n4721 GND.n4652 163.367
R18887 GND.n5081 GND.n5078 163.367
R18888 GND.n5085 GND.n5078 163.367
R18889 GND.n5089 GND.n5087 163.367
R18890 GND.n5093 GND.n5076 163.367
R18891 GND.n5097 GND.n5095 163.367
R18892 GND.n5101 GND.n5074 163.367
R18893 GND.n5105 GND.n5103 163.367
R18894 GND.n5109 GND.n5072 163.367
R18895 GND.n5113 GND.n5111 163.367
R18896 GND.n5117 GND.n5070 163.367
R18897 GND.n5121 GND.n5119 163.367
R18898 GND.n5125 GND.n5068 163.367
R18899 GND.n5129 GND.n5127 163.367
R18900 GND.n5134 GND.n5064 163.367
R18901 GND.n5137 GND.n5136 163.367
R18902 GND.n5139 GND.n5061 163.367
R18903 GND.n5143 GND.n5059 163.367
R18904 GND.n5147 GND.n5145 163.367
R18905 GND.n5152 GND.n5055 163.367
R18906 GND.n5156 GND.n5154 163.367
R18907 GND.n5160 GND.n5053 163.367
R18908 GND.n5164 GND.n5162 163.367
R18909 GND.n5168 GND.n5051 163.367
R18910 GND.n5172 GND.n5170 163.367
R18911 GND.n5176 GND.n5049 163.367
R18912 GND.n5180 GND.n5178 163.367
R18913 GND.n5184 GND.n5047 163.367
R18914 GND.n5188 GND.n5186 163.367
R18915 GND.n5192 GND.n5045 163.367
R18916 GND.n5196 GND.n5194 163.367
R18917 GND.n5200 GND.n5043 163.367
R18918 GND.n5203 GND.n5202 163.367
R18919 GND.n8125 GND.n3753 163.367
R18920 GND.n8121 GND.n3753 163.367
R18921 GND.n8121 GND.n3769 163.367
R18922 GND.n5213 GND.n3769 163.367
R18923 GND.n5213 GND.n3782 163.367
R18924 GND.n8111 GND.n3782 163.367
R18925 GND.n8111 GND.n3783 163.367
R18926 GND.n8107 GND.n3783 163.367
R18927 GND.n8107 GND.n3786 163.367
R18928 GND.n5226 GND.n3786 163.367
R18929 GND.n5226 GND.n3799 163.367
R18930 GND.n8097 GND.n3799 163.367
R18931 GND.n8097 GND.n3800 163.367
R18932 GND.n8093 GND.n3800 163.367
R18933 GND.n8093 GND.n3803 163.367
R18934 GND.n5239 GND.n3803 163.367
R18935 GND.n5239 GND.n3817 163.367
R18936 GND.n8083 GND.n3817 163.367
R18937 GND.n8083 GND.n3818 163.367
R18938 GND.n8079 GND.n3818 163.367
R18939 GND.n8079 GND.n3821 163.367
R18940 GND.n5252 GND.n3821 163.367
R18941 GND.n5252 GND.n3835 163.367
R18942 GND.n8069 GND.n3835 163.367
R18943 GND.n8069 GND.n3836 163.367
R18944 GND.n8065 GND.n3836 163.367
R18945 GND.n8065 GND.n3839 163.367
R18946 GND.n5306 GND.n3839 163.367
R18947 GND.n5309 GND.n5306 163.367
R18948 GND.n5310 GND.n5309 163.367
R18949 GND.n5311 GND.n5310 163.367
R18950 GND.n5311 GND.n3883 163.367
R18951 GND.n5315 GND.n3883 163.367
R18952 GND.n5316 GND.n5315 163.367
R18953 GND.n5317 GND.n5316 163.367
R18954 GND.n5317 GND.n5032 163.367
R18955 GND.n5322 GND.n5032 163.367
R18956 GND.n5322 GND.n5019 163.367
R18957 GND.n5334 GND.n5019 163.367
R18958 GND.n5335 GND.n5334 163.367
R18959 GND.n5335 GND.n5016 163.367
R18960 GND.n5341 GND.n5016 163.367
R18961 GND.n5341 GND.n5017 163.367
R18962 GND.n5017 GND.n5010 163.367
R18963 GND.n5353 GND.n5010 163.367
R18964 GND.n5354 GND.n5353 163.367
R18965 GND.n5354 GND.n5007 163.367
R18966 GND.n5360 GND.n5007 163.367
R18967 GND.n5360 GND.n5008 163.367
R18968 GND.n5008 GND.n5001 163.367
R18969 GND.n5413 GND.n5001 163.367
R18970 GND.n5414 GND.n5413 163.367
R18971 GND.n5414 GND.n4998 163.367
R18972 GND.n5420 GND.n4998 163.367
R18973 GND.n5420 GND.n4999 163.367
R18974 GND.n4999 GND.n4991 163.367
R18975 GND.n5431 GND.n4991 163.367
R18976 GND.n5432 GND.n5431 163.367
R18977 GND.n5432 GND.n4988 163.367
R18978 GND.n5438 GND.n4988 163.367
R18979 GND.n5438 GND.n4989 163.367
R18980 GND.n4989 GND.n4982 163.367
R18981 GND.n5449 GND.n4982 163.367
R18982 GND.n5450 GND.n5449 163.367
R18983 GND.n5450 GND.n4979 163.367
R18984 GND.n5456 GND.n4979 163.367
R18985 GND.n5456 GND.n4980 163.367
R18986 GND.n4980 GND.n4972 163.367
R18987 GND.n5467 GND.n4972 163.367
R18988 GND.n5468 GND.n5467 163.367
R18989 GND.n5468 GND.n4969 163.367
R18990 GND.n5474 GND.n4969 163.367
R18991 GND.n5474 GND.n4970 163.367
R18992 GND.n4970 GND.n4962 163.367
R18993 GND.n5491 GND.n4962 163.367
R18994 GND.n5492 GND.n5491 163.367
R18995 GND.n5492 GND.n4959 163.367
R18996 GND.n5502 GND.n4959 163.367
R18997 GND.n5502 GND.n4960 163.367
R18998 GND.n5498 GND.n4960 163.367
R18999 GND.n5498 GND.n5497 163.367
R19000 GND.n5497 GND.n4055 163.367
R19001 GND.n4066 GND.n4055 163.367
R19002 GND.n7896 GND.n4066 163.367
R19003 GND.n7896 GND.n4067 163.367
R19004 GND.n7892 GND.n4067 163.367
R19005 GND.n7892 GND.n4070 163.367
R19006 GND.n5552 GND.n4070 163.367
R19007 GND.n5553 GND.n5552 163.367
R19008 GND.n5553 GND.n4948 163.367
R19009 GND.n5559 GND.n4948 163.367
R19010 GND.n5559 GND.n4949 163.367
R19011 GND.n4949 GND.n4941 163.367
R19012 GND.n5570 GND.n4941 163.367
R19013 GND.n5571 GND.n5570 163.367
R19014 GND.n5571 GND.n4938 163.367
R19015 GND.n5577 GND.n4938 163.367
R19016 GND.n5577 GND.n4939 163.367
R19017 GND.n4939 GND.n4931 163.367
R19018 GND.n5594 GND.n4931 163.367
R19019 GND.n5595 GND.n5594 163.367
R19020 GND.n5595 GND.n4928 163.367
R19021 GND.n5605 GND.n4928 163.367
R19022 GND.n5605 GND.n4929 163.367
R19023 GND.n5601 GND.n4929 163.367
R19024 GND.n5601 GND.n5600 163.367
R19025 GND.n5600 GND.n4160 163.367
R19026 GND.n4171 GND.n4160 163.367
R19027 GND.n7841 GND.n4171 163.367
R19028 GND.n7841 GND.n4172 163.367
R19029 GND.n7837 GND.n4172 163.367
R19030 GND.n7837 GND.n4175 163.367
R19031 GND.n5656 GND.n4175 163.367
R19032 GND.n5657 GND.n5656 163.367
R19033 GND.n5657 GND.n4917 163.367
R19034 GND.n5663 GND.n4917 163.367
R19035 GND.n5663 GND.n4918 163.367
R19036 GND.n4918 GND.n4909 163.367
R19037 GND.n5674 GND.n4909 163.367
R19038 GND.n5675 GND.n5674 163.367
R19039 GND.n5675 GND.n4906 163.367
R19040 GND.n5682 GND.n4906 163.367
R19041 GND.n5682 GND.n4907 163.367
R19042 GND.n5678 GND.n4907 163.367
R19043 GND.n5678 GND.n4898 163.367
R19044 GND.n5698 GND.n4898 163.367
R19045 GND.n5698 GND.n4895 163.367
R19046 GND.n5708 GND.n4895 163.367
R19047 GND.n5708 GND.n4896 163.367
R19048 GND.n5704 GND.n4896 163.367
R19049 GND.n5704 GND.n5703 163.367
R19050 GND.n5703 GND.n4262 163.367
R19051 GND.n4273 GND.n4262 163.367
R19052 GND.n7786 GND.n4273 163.367
R19053 GND.n7786 GND.n4274 163.367
R19054 GND.n7782 GND.n4274 163.367
R19055 GND.n7782 GND.n4277 163.367
R19056 GND.n5753 GND.n4277 163.367
R19057 GND.n5754 GND.n5753 163.367
R19058 GND.n5754 GND.n4883 163.367
R19059 GND.n5760 GND.n4883 163.367
R19060 GND.n5760 GND.n4884 163.367
R19061 GND.n4884 GND.n4876 163.367
R19062 GND.n5771 GND.n4876 163.367
R19063 GND.n5772 GND.n5771 163.367
R19064 GND.n5772 GND.n4873 163.367
R19065 GND.n5777 GND.n4873 163.367
R19066 GND.n5777 GND.n4874 163.367
R19067 GND.n4874 GND.n4854 163.367
R19068 GND.n5799 GND.n4854 163.367
R19069 GND.n5799 GND.n4855 163.367
R19070 GND.n5795 GND.n4855 163.367
R19071 GND.n5795 GND.n4865 163.367
R19072 GND.n4865 GND.n4864 163.367
R19073 GND.n4864 GND.n4858 163.367
R19074 GND.n4860 GND.n4858 163.367
R19075 GND.n4860 GND.n4366 163.367
R19076 GND.n4377 GND.n4366 163.367
R19077 GND.n7731 GND.n4377 163.367
R19078 GND.n7731 GND.n4378 163.367
R19079 GND.n7727 GND.n4378 163.367
R19080 GND.n7727 GND.n4381 163.367
R19081 GND.n4462 GND.n4381 163.367
R19082 GND.n4462 GND.n4399 163.367
R19083 GND.n7717 GND.n4399 163.367
R19084 GND.n7717 GND.n4400 163.367
R19085 GND.n7713 GND.n4400 163.367
R19086 GND.n7713 GND.n4403 163.367
R19087 GND.n4475 GND.n4403 163.367
R19088 GND.n4475 GND.n4417 163.367
R19089 GND.n7703 GND.n4417 163.367
R19090 GND.n7703 GND.n4418 163.367
R19091 GND.n7699 GND.n4418 163.367
R19092 GND.n7699 GND.n4421 163.367
R19093 GND.n4488 GND.n4421 163.367
R19094 GND.n4488 GND.n4435 163.367
R19095 GND.n7689 GND.n4435 163.367
R19096 GND.n7689 GND.n4436 163.367
R19097 GND.n7685 GND.n4436 163.367
R19098 GND.n7685 GND.n4439 163.367
R19099 GND.n4508 GND.n4439 163.367
R19100 GND.n4508 GND.n4450 163.367
R19101 GND.n4506 GND.n4450 163.367
R19102 GND.n7670 GND.n4506 163.367
R19103 GND.n7670 GND.n4507 163.367
R19104 GND.n7666 GND.n4507 163.367
R19105 GND.n7666 GND.n4513 163.367
R19106 GND.n4723 GND.n4513 163.367
R19107 GND.n4726 GND.n4723 163.367
R19108 GND.n40 GND.t36 156.31
R19109 GND.n42 GND.t34 155.48
R19110 GND.n41 GND.t13 155.48
R19111 GND.n40 GND.t209 155.48
R19112 GND.n4639 GND.t86 153.965
R19113 GND.n4648 GND.n4647 152.776
R19114 GND.n3764 GND.n3754 152
R19115 GND.n3766 GND.n3765 152
R19116 GND.n4646 GND.n4637 152
R19117 GND.n4790 GND.n4543 143.351
R19118 GND.n4790 GND.n4544 143.351
R19119 GND.n3761 GND.t63 137.107
R19120 GND.n3765 GND.t110 126.766
R19121 GND.n3763 GND.t149 126.766
R19122 GND.n3762 GND.t89 126.766
R19123 GND.n4638 GND.t152 126.766
R19124 GND.n4645 GND.t107 126.766
R19125 GND.n4647 GND.t57 126.766
R19126 GND.n4811 GND.n4810 125.868
R19127 GND.n10785 GND.n10784 125.868
R19128 GND.n5056 GND.t141 121.709
R19129 GND.n4655 GND.t67 121.709
R19130 GND.n5065 GND.t132 121.703
R19131 GND.n4635 GND.t51 121.703
R19132 GND.n8013 GND.t116 116.615
R19133 GND.n5860 GND.t147 116.615
R19134 GND.n2915 GND.n2914 113.067
R19135 GND.n8333 GND.n8332 113.067
R19136 GND.n8383 GND.n8382 113.067
R19137 GND.n8407 GND.n8406 113.067
R19138 GND.n2184 GND.n2183 113.067
R19139 GND.n4621 GND.n4620 113.067
R19140 GND.n4795 GND.n4794 113.067
R19141 GND.n4829 GND.n4828 113.067
R19142 GND.n10766 GND.n10765 113.067
R19143 GND.n10749 GND.n10748 113.067
R19144 GND.n10733 GND.n10732 113.067
R19145 GND.n457 GND.n456 113.067
R19146 GND.n5887 GND.n5886 113.067
R19147 GND.n1744 GND.n1743 113.067
R19148 GND.n1760 GND.n1759 113.067
R19149 GND.n1777 GND.n1776 113.067
R19150 GND.n1795 GND.n1794 113.067
R19151 GND.n2144 GND.n2143 113.067
R19152 GND.n10895 GND.n10894 99.6594
R19153 GND.n10890 GND.n10714 99.6594
R19154 GND.n10886 GND.n10713 99.6594
R19155 GND.n10882 GND.n10712 99.6594
R19156 GND.n10878 GND.n10711 99.6594
R19157 GND.n10735 GND.n10710 99.6594
R19158 GND.n10870 GND.n10709 99.6594
R19159 GND.n10866 GND.n10708 99.6594
R19160 GND.n10862 GND.n10707 99.6594
R19161 GND.n10858 GND.n10706 99.6594
R19162 GND.n10854 GND.n10705 99.6594
R19163 GND.n10850 GND.n10704 99.6594
R19164 GND.n10846 GND.n10703 99.6594
R19165 GND.n10842 GND.n10702 99.6594
R19166 GND.n10838 GND.n10701 99.6594
R19167 GND.n10834 GND.n10700 99.6594
R19168 GND.n10830 GND.n10699 99.6594
R19169 GND.n10826 GND.n10698 99.6594
R19170 GND.n10822 GND.n10697 99.6594
R19171 GND.n10818 GND.n10696 99.6594
R19172 GND.n10814 GND.n10695 99.6594
R19173 GND.n10810 GND.n10694 99.6594
R19174 GND.n10806 GND.n10693 99.6594
R19175 GND.n10802 GND.n10692 99.6594
R19176 GND.n10798 GND.n10691 99.6594
R19177 GND.n10794 GND.n10690 99.6594
R19178 GND.n10790 GND.n10689 99.6594
R19179 GND.n10782 GND.n10688 99.6594
R19180 GND.n7646 GND.n7645 99.6594
R19181 GND.n7640 GND.n4568 99.6594
R19182 GND.n7637 GND.n4569 99.6594
R19183 GND.n7633 GND.n4570 99.6594
R19184 GND.n7629 GND.n4571 99.6594
R19185 GND.n7625 GND.n4572 99.6594
R19186 GND.n7621 GND.n4573 99.6594
R19187 GND.n7618 GND.n4574 99.6594
R19188 GND.n7614 GND.n4575 99.6594
R19189 GND.n7610 GND.n4576 99.6594
R19190 GND.n7606 GND.n4577 99.6594
R19191 GND.n7602 GND.n4578 99.6594
R19192 GND.n7598 GND.n4579 99.6594
R19193 GND.n7595 GND.n4580 99.6594
R19194 GND.n7592 GND.n4581 99.6594
R19195 GND.n7588 GND.n4582 99.6594
R19196 GND.n7584 GND.n4583 99.6594
R19197 GND.n7580 GND.n4584 99.6594
R19198 GND.n7576 GND.n4585 99.6594
R19199 GND.n7572 GND.n4586 99.6594
R19200 GND.n7568 GND.n4587 99.6594
R19201 GND.n7564 GND.n4588 99.6594
R19202 GND.n7560 GND.n4589 99.6594
R19203 GND.n7556 GND.n4590 99.6594
R19204 GND.n7552 GND.n4591 99.6594
R19205 GND.n7548 GND.n4592 99.6594
R19206 GND.n7544 GND.n4593 99.6594
R19207 GND.n7540 GND.n4594 99.6594
R19208 GND.n2209 GND.n2148 99.6594
R19209 GND.n8316 GND.n2149 99.6594
R19210 GND.n2205 GND.n2150 99.6594
R19211 GND.n8324 GND.n2151 99.6594
R19212 GND.n2201 GND.n2152 99.6594
R19213 GND.n8334 GND.n2153 99.6594
R19214 GND.n2197 GND.n2154 99.6594
R19215 GND.n8342 GND.n2155 99.6594
R19216 GND.n2193 GND.n2156 99.6594
R19217 GND.n8350 GND.n2157 99.6594
R19218 GND.n2189 GND.n2158 99.6594
R19219 GND.n8358 GND.n2159 99.6594
R19220 GND.n8456 GND.n2182 99.6594
R19221 GND.n8364 GND.n2181 99.6594
R19222 GND.n8366 GND.n2180 99.6594
R19223 GND.n8370 GND.n2179 99.6594
R19224 GND.n8372 GND.n2178 99.6594
R19225 GND.n8376 GND.n2177 99.6594
R19226 GND.n8378 GND.n2176 99.6594
R19227 GND.n8385 GND.n2175 99.6594
R19228 GND.n8387 GND.n2174 99.6594
R19229 GND.n8391 GND.n2173 99.6594
R19230 GND.n8393 GND.n2172 99.6594
R19231 GND.n8397 GND.n2171 99.6594
R19232 GND.n8399 GND.n2170 99.6594
R19233 GND.n8403 GND.n2169 99.6594
R19234 GND.n8405 GND.n2168 99.6594
R19235 GND.n2167 GND.n2124 99.6594
R19236 GND.n8815 GND.n8814 99.6594
R19237 GND.n8809 GND.n1691 99.6594
R19238 GND.n8806 GND.n1692 99.6594
R19239 GND.n8802 GND.n1693 99.6594
R19240 GND.n8798 GND.n1694 99.6594
R19241 GND.n8794 GND.n1695 99.6594
R19242 GND.n8790 GND.n1696 99.6594
R19243 GND.n8787 GND.n1697 99.6594
R19244 GND.n8783 GND.n1698 99.6594
R19245 GND.n8779 GND.n1699 99.6594
R19246 GND.n8775 GND.n1700 99.6594
R19247 GND.n8771 GND.n1701 99.6594
R19248 GND.n8767 GND.n1702 99.6594
R19249 GND.n8763 GND.n1703 99.6594
R19250 GND.n8759 GND.n1704 99.6594
R19251 GND.n8755 GND.n1705 99.6594
R19252 GND.n8751 GND.n1706 99.6594
R19253 GND.n8747 GND.n1707 99.6594
R19254 GND.n8743 GND.n1708 99.6594
R19255 GND.n8739 GND.n1709 99.6594
R19256 GND.n8735 GND.n1710 99.6594
R19257 GND.n8731 GND.n1711 99.6594
R19258 GND.n8727 GND.n1712 99.6594
R19259 GND.n8723 GND.n1713 99.6594
R19260 GND.n8719 GND.n1714 99.6594
R19261 GND.n8715 GND.n1715 99.6594
R19262 GND.n8711 GND.n1716 99.6594
R19263 GND.n8707 GND.n1717 99.6594
R19264 GND.n5817 GND.n4847 99.6594
R19265 GND.n5827 GND.n5826 99.6594
R19266 GND.n5831 GND.n4845 99.6594
R19267 GND.n5835 GND.n5834 99.6594
R19268 GND.n5839 GND.n5838 99.6594
R19269 GND.n5844 GND.n5843 99.6594
R19270 GND.n5849 GND.n5848 99.6594
R19271 GND.n5854 GND.n5853 99.6594
R19272 GND.n5859 GND.n5858 99.6594
R19273 GND.n5867 GND.n5866 99.6594
R19274 GND.n5869 GND.n5868 99.6594
R19275 GND.n8055 GND.n8054 99.6594
R19276 GND.n8049 GND.n3851 99.6594
R19277 GND.n8046 GND.n3852 99.6594
R19278 GND.n3872 GND.n3853 99.6594
R19279 GND.n8039 GND.n3854 99.6594
R19280 GND.n8034 GND.n3855 99.6594
R19281 GND.n8029 GND.n3856 99.6594
R19282 GND.n8024 GND.n3857 99.6594
R19283 GND.n8019 GND.n3858 99.6594
R19284 GND.n8011 GND.n3859 99.6594
R19285 GND.n3878 GND.n3860 99.6594
R19286 GND.n10687 GND.n10686 99.6594
R19287 GND.n10680 GND.n10651 99.6594
R19288 GND.n10676 GND.n10650 99.6594
R19289 GND.n10672 GND.n10649 99.6594
R19290 GND.n10668 GND.n10648 99.6594
R19291 GND.n10664 GND.n10647 99.6594
R19292 GND.n10898 GND.n10897 99.6594
R19293 GND.n5916 GND.n4595 99.6594
R19294 GND.n5912 GND.n4596 99.6594
R19295 GND.n5907 GND.n4597 99.6594
R19296 GND.n5902 GND.n4598 99.6594
R19297 GND.n5897 GND.n4599 99.6594
R19298 GND.n5892 GND.n4600 99.6594
R19299 GND.n5885 GND.n4601 99.6594
R19300 GND.n5913 GND.n4595 99.6594
R19301 GND.n5908 GND.n4596 99.6594
R19302 GND.n5903 GND.n4597 99.6594
R19303 GND.n5898 GND.n4598 99.6594
R19304 GND.n5893 GND.n4599 99.6594
R19305 GND.n5882 GND.n4600 99.6594
R19306 GND.n5883 GND.n4601 99.6594
R19307 GND.n10897 GND.n459 99.6594
R19308 GND.n10667 GND.n10647 99.6594
R19309 GND.n10671 GND.n10648 99.6594
R19310 GND.n10675 GND.n10649 99.6594
R19311 GND.n10679 GND.n10650 99.6594
R19312 GND.n10652 GND.n10651 99.6594
R19313 GND.n10687 GND.n449 99.6594
R19314 GND.n8055 GND.n3863 99.6594
R19315 GND.n8047 GND.n3851 99.6594
R19316 GND.n3871 GND.n3852 99.6594
R19317 GND.n8038 GND.n3853 99.6594
R19318 GND.n8033 GND.n3854 99.6594
R19319 GND.n8028 GND.n3855 99.6594
R19320 GND.n8023 GND.n3856 99.6594
R19321 GND.n8018 GND.n3857 99.6594
R19322 GND.n8012 GND.n3858 99.6594
R19323 GND.n3877 GND.n3859 99.6594
R19324 GND.n8007 GND.n3860 99.6594
R19325 GND.n5870 GND.n5869 99.6594
R19326 GND.n5866 GND.n5865 99.6594
R19327 GND.n5858 GND.n5857 99.6594
R19328 GND.n5853 GND.n5852 99.6594
R19329 GND.n5848 GND.n5847 99.6594
R19330 GND.n5843 GND.n5842 99.6594
R19331 GND.n5838 GND.n5837 99.6594
R19332 GND.n5834 GND.n5833 99.6594
R19333 GND.n5828 GND.n4845 99.6594
R19334 GND.n5826 GND.n5825 99.6594
R19335 GND.n5818 GND.n5817 99.6594
R19336 GND.n8815 GND.n1727 99.6594
R19337 GND.n8807 GND.n1691 99.6594
R19338 GND.n8803 GND.n1692 99.6594
R19339 GND.n8799 GND.n1693 99.6594
R19340 GND.n8795 GND.n1694 99.6594
R19341 GND.n1741 GND.n1695 99.6594
R19342 GND.n8788 GND.n1696 99.6594
R19343 GND.n8784 GND.n1697 99.6594
R19344 GND.n8780 GND.n1698 99.6594
R19345 GND.n8776 GND.n1699 99.6594
R19346 GND.n8772 GND.n1700 99.6594
R19347 GND.n8768 GND.n1701 99.6594
R19348 GND.n8764 GND.n1702 99.6594
R19349 GND.n8760 GND.n1703 99.6594
R19350 GND.n8756 GND.n1704 99.6594
R19351 GND.n8752 GND.n1705 99.6594
R19352 GND.n8748 GND.n1706 99.6594
R19353 GND.n8744 GND.n1707 99.6594
R19354 GND.n8740 GND.n1708 99.6594
R19355 GND.n8736 GND.n1709 99.6594
R19356 GND.n8732 GND.n1710 99.6594
R19357 GND.n8728 GND.n1711 99.6594
R19358 GND.n8724 GND.n1712 99.6594
R19359 GND.n8720 GND.n1713 99.6594
R19360 GND.n8716 GND.n1714 99.6594
R19361 GND.n8712 GND.n1715 99.6594
R19362 GND.n8708 GND.n1716 99.6594
R19363 GND.n1802 GND.n1717 99.6594
R19364 GND.n8409 GND.n2167 99.6594
R19365 GND.n8404 GND.n2168 99.6594
R19366 GND.n8400 GND.n2169 99.6594
R19367 GND.n8398 GND.n2170 99.6594
R19368 GND.n8394 GND.n2171 99.6594
R19369 GND.n8392 GND.n2172 99.6594
R19370 GND.n8388 GND.n2173 99.6594
R19371 GND.n8386 GND.n2174 99.6594
R19372 GND.n8379 GND.n2175 99.6594
R19373 GND.n8377 GND.n2176 99.6594
R19374 GND.n8373 GND.n2177 99.6594
R19375 GND.n8371 GND.n2178 99.6594
R19376 GND.n8367 GND.n2179 99.6594
R19377 GND.n8365 GND.n2180 99.6594
R19378 GND.n8455 GND.n2181 99.6594
R19379 GND.n8359 GND.n2160 99.6594
R19380 GND.n2190 GND.n2159 99.6594
R19381 GND.n8351 GND.n2158 99.6594
R19382 GND.n2194 GND.n2157 99.6594
R19383 GND.n8343 GND.n2156 99.6594
R19384 GND.n2198 GND.n2155 99.6594
R19385 GND.n8335 GND.n2154 99.6594
R19386 GND.n2202 GND.n2153 99.6594
R19387 GND.n8325 GND.n2152 99.6594
R19388 GND.n2206 GND.n2151 99.6594
R19389 GND.n8317 GND.n2150 99.6594
R19390 GND.n2210 GND.n2149 99.6594
R19391 GND.n8309 GND.n2148 99.6594
R19392 GND.n7646 GND.n4604 99.6594
R19393 GND.n7638 GND.n4568 99.6594
R19394 GND.n7634 GND.n4569 99.6594
R19395 GND.n7630 GND.n4570 99.6594
R19396 GND.n7626 GND.n4571 99.6594
R19397 GND.n4618 GND.n4572 99.6594
R19398 GND.n7619 GND.n4573 99.6594
R19399 GND.n7615 GND.n4574 99.6594
R19400 GND.n7611 GND.n4575 99.6594
R19401 GND.n7607 GND.n4576 99.6594
R19402 GND.n7603 GND.n4577 99.6594
R19403 GND.n7599 GND.n4578 99.6594
R19404 GND.n4792 GND.n4579 99.6594
R19405 GND.n7593 GND.n4580 99.6594
R19406 GND.n7589 GND.n4581 99.6594
R19407 GND.n7585 GND.n4582 99.6594
R19408 GND.n7581 GND.n4583 99.6594
R19409 GND.n7577 GND.n4584 99.6594
R19410 GND.n7573 GND.n4585 99.6594
R19411 GND.n7569 GND.n4586 99.6594
R19412 GND.n7565 GND.n4587 99.6594
R19413 GND.n7561 GND.n4588 99.6594
R19414 GND.n7557 GND.n4589 99.6594
R19415 GND.n7553 GND.n4590 99.6594
R19416 GND.n7549 GND.n4591 99.6594
R19417 GND.n7545 GND.n4592 99.6594
R19418 GND.n7541 GND.n4593 99.6594
R19419 GND.n5877 GND.n4594 99.6594
R19420 GND.n10789 GND.n10688 99.6594
R19421 GND.n10793 GND.n10689 99.6594
R19422 GND.n10797 GND.n10690 99.6594
R19423 GND.n10801 GND.n10691 99.6594
R19424 GND.n10805 GND.n10692 99.6594
R19425 GND.n10809 GND.n10693 99.6594
R19426 GND.n10813 GND.n10694 99.6594
R19427 GND.n10817 GND.n10695 99.6594
R19428 GND.n10821 GND.n10696 99.6594
R19429 GND.n10825 GND.n10697 99.6594
R19430 GND.n10829 GND.n10698 99.6594
R19431 GND.n10833 GND.n10699 99.6594
R19432 GND.n10837 GND.n10700 99.6594
R19433 GND.n10841 GND.n10701 99.6594
R19434 GND.n10845 GND.n10702 99.6594
R19435 GND.n10849 GND.n10703 99.6594
R19436 GND.n10853 GND.n10704 99.6594
R19437 GND.n10857 GND.n10705 99.6594
R19438 GND.n10861 GND.n10706 99.6594
R19439 GND.n10865 GND.n10707 99.6594
R19440 GND.n10869 GND.n10708 99.6594
R19441 GND.n10734 GND.n10709 99.6594
R19442 GND.n10877 GND.n10710 99.6594
R19443 GND.n10881 GND.n10711 99.6594
R19444 GND.n10885 GND.n10712 99.6594
R19445 GND.n10889 GND.n10713 99.6594
R19446 GND.n10716 GND.n10714 99.6594
R19447 GND.n10895 GND.n10715 99.6594
R19448 GND.n8700 GND.n1718 99.6594
R19449 GND.n2922 GND.n1719 99.6594
R19450 GND.n2928 GND.n1720 99.6594
R19451 GND.n2930 GND.n1721 99.6594
R19452 GND.n2938 GND.n1722 99.6594
R19453 GND.n2940 GND.n1723 99.6594
R19454 GND.n2913 GND.n1724 99.6594
R19455 GND.n2921 GND.n1718 99.6594
R19456 GND.n2927 GND.n1719 99.6594
R19457 GND.n2931 GND.n1720 99.6594
R19458 GND.n2937 GND.n1721 99.6594
R19459 GND.n2941 GND.n1722 99.6594
R19460 GND.n2917 GND.n1723 99.6594
R19461 GND.n2948 GND.n1724 99.6594
R19462 GND.n8478 GND.n2130 99.6594
R19463 GND.n2161 GND.n2133 99.6594
R19464 GND.n2162 GND.n2135 99.6594
R19465 GND.n2163 GND.n2137 99.6594
R19466 GND.n2164 GND.n2139 99.6594
R19467 GND.n2165 GND.n2141 99.6594
R19468 GND.n8459 GND.n8458 99.6594
R19469 GND.n8458 GND.n2146 99.6594
R19470 GND.n2165 GND.n2142 99.6594
R19471 GND.n2164 GND.n2140 99.6594
R19472 GND.n2163 GND.n2138 99.6594
R19473 GND.n2162 GND.n2136 99.6594
R19474 GND.n2161 GND.n2134 99.6594
R19475 GND.n2132 GND.n2130 99.6594
R19476 GND.n43 GND.t7 88.8196
R19477 GND.n45 GND.t207 87.9882
R19478 GND.n44 GND.t9 87.9882
R19479 GND.n43 GND.t198 87.9882
R19480 GND.n3761 GND.n3760 74.9819
R19481 GND.n3762 GND.n3756 72.8411
R19482 GND.n3763 GND.n3755 72.8411
R19483 GND.n4645 GND.n4644 72.8411
R19484 GND.n4730 GND.n4528 71.676
R19485 GND.n4734 GND.n4529 71.676
R19486 GND.n4738 GND.n4530 71.676
R19487 GND.n4742 GND.n4531 71.676
R19488 GND.n4746 GND.n4532 71.676
R19489 GND.n4750 GND.n4533 71.676
R19490 GND.n4754 GND.n4534 71.676
R19491 GND.n4758 GND.n4535 71.676
R19492 GND.n4762 GND.n4536 71.676
R19493 GND.n4766 GND.n4537 71.676
R19494 GND.n4770 GND.n4538 71.676
R19495 GND.n4774 GND.n4539 71.676
R19496 GND.n4778 GND.n4540 71.676
R19497 GND.n4783 GND.n4541 71.676
R19498 GND.n4787 GND.n4542 71.676
R19499 GND.n4657 GND.n4544 71.676
R19500 GND.n4661 GND.n4545 71.676
R19501 GND.n4666 GND.n4546 71.676
R19502 GND.n4670 GND.n4547 71.676
R19503 GND.n4674 GND.n4548 71.676
R19504 GND.n4678 GND.n4549 71.676
R19505 GND.n4682 GND.n4550 71.676
R19506 GND.n4686 GND.n4551 71.676
R19507 GND.n4690 GND.n4552 71.676
R19508 GND.n4694 GND.n4553 71.676
R19509 GND.n4698 GND.n4554 71.676
R19510 GND.n4702 GND.n4555 71.676
R19511 GND.n4706 GND.n4556 71.676
R19512 GND.n4710 GND.n4557 71.676
R19513 GND.n4714 GND.n4558 71.676
R19514 GND.n4717 GND.n4559 71.676
R19515 GND.n5080 GND.n3752 71.676
R19516 GND.n5086 GND.n5085 71.676
R19517 GND.n5089 GND.n5088 71.676
R19518 GND.n5094 GND.n5093 71.676
R19519 GND.n5097 GND.n5096 71.676
R19520 GND.n5102 GND.n5101 71.676
R19521 GND.n5105 GND.n5104 71.676
R19522 GND.n5110 GND.n5109 71.676
R19523 GND.n5113 GND.n5112 71.676
R19524 GND.n5118 GND.n5117 71.676
R19525 GND.n5121 GND.n5120 71.676
R19526 GND.n5126 GND.n5125 71.676
R19527 GND.n5129 GND.n5128 71.676
R19528 GND.n5135 GND.n5134 71.676
R19529 GND.n5138 GND.n5137 71.676
R19530 GND.n5061 GND.n5060 71.676
R19531 GND.n5144 GND.n5143 71.676
R19532 GND.n5147 GND.n5146 71.676
R19533 GND.n5153 GND.n5152 71.676
R19534 GND.n5156 GND.n5155 71.676
R19535 GND.n5161 GND.n5160 71.676
R19536 GND.n5164 GND.n5163 71.676
R19537 GND.n5169 GND.n5168 71.676
R19538 GND.n5172 GND.n5171 71.676
R19539 GND.n5177 GND.n5176 71.676
R19540 GND.n5180 GND.n5179 71.676
R19541 GND.n5185 GND.n5184 71.676
R19542 GND.n5188 GND.n5187 71.676
R19543 GND.n5193 GND.n5192 71.676
R19544 GND.n5196 GND.n5195 71.676
R19545 GND.n5201 GND.n5200 71.676
R19546 GND.n5081 GND.n5080 71.676
R19547 GND.n5087 GND.n5086 71.676
R19548 GND.n5088 GND.n5076 71.676
R19549 GND.n5095 GND.n5094 71.676
R19550 GND.n5096 GND.n5074 71.676
R19551 GND.n5103 GND.n5102 71.676
R19552 GND.n5104 GND.n5072 71.676
R19553 GND.n5111 GND.n5110 71.676
R19554 GND.n5112 GND.n5070 71.676
R19555 GND.n5119 GND.n5118 71.676
R19556 GND.n5120 GND.n5068 71.676
R19557 GND.n5127 GND.n5126 71.676
R19558 GND.n5128 GND.n5064 71.676
R19559 GND.n5136 GND.n5135 71.676
R19560 GND.n5139 GND.n5138 71.676
R19561 GND.n5060 GND.n5059 71.676
R19562 GND.n5145 GND.n5144 71.676
R19563 GND.n5146 GND.n5055 71.676
R19564 GND.n5154 GND.n5153 71.676
R19565 GND.n5155 GND.n5053 71.676
R19566 GND.n5162 GND.n5161 71.676
R19567 GND.n5163 GND.n5051 71.676
R19568 GND.n5170 GND.n5169 71.676
R19569 GND.n5171 GND.n5049 71.676
R19570 GND.n5178 GND.n5177 71.676
R19571 GND.n5179 GND.n5047 71.676
R19572 GND.n5186 GND.n5185 71.676
R19573 GND.n5187 GND.n5045 71.676
R19574 GND.n5194 GND.n5193 71.676
R19575 GND.n5195 GND.n5043 71.676
R19576 GND.n5202 GND.n5201 71.676
R19577 GND.n4715 GND.n4559 71.676
R19578 GND.n4711 GND.n4558 71.676
R19579 GND.n4707 GND.n4557 71.676
R19580 GND.n4703 GND.n4556 71.676
R19581 GND.n4699 GND.n4555 71.676
R19582 GND.n4695 GND.n4554 71.676
R19583 GND.n4691 GND.n4553 71.676
R19584 GND.n4687 GND.n4552 71.676
R19585 GND.n4683 GND.n4551 71.676
R19586 GND.n4679 GND.n4550 71.676
R19587 GND.n4675 GND.n4549 71.676
R19588 GND.n4671 GND.n4548 71.676
R19589 GND.n4667 GND.n4547 71.676
R19590 GND.n4662 GND.n4546 71.676
R19591 GND.n4658 GND.n4545 71.676
R19592 GND.n4788 GND.n4543 71.676
R19593 GND.n4784 GND.n4542 71.676
R19594 GND.n4779 GND.n4541 71.676
R19595 GND.n4775 GND.n4540 71.676
R19596 GND.n4771 GND.n4539 71.676
R19597 GND.n4767 GND.n4538 71.676
R19598 GND.n4763 GND.n4537 71.676
R19599 GND.n4759 GND.n4536 71.676
R19600 GND.n4755 GND.n4535 71.676
R19601 GND.n4751 GND.n4534 71.676
R19602 GND.n4747 GND.n4533 71.676
R19603 GND.n4743 GND.n4532 71.676
R19604 GND.n4739 GND.n4531 71.676
R19605 GND.n4735 GND.n4530 71.676
R19606 GND.n4731 GND.n4529 71.676
R19607 GND.n4727 GND.n4528 71.676
R19608 GND.n8014 GND.t115 71.6217
R19609 GND.n5861 GND.t148 71.6217
R19610 GND.n5066 GND.n5065 66.7156
R19611 GND.n5057 GND.n5056 66.7156
R19612 GND.n4656 GND.n4655 66.7156
R19613 GND.n4636 GND.n4635 66.7156
R19614 GND.n8 GND.t163 63.7546
R19615 GND.n15 GND.t202 63.7546
R19616 GND.n23 GND.t161 63.7546
R19617 GND.n31 GND.t23 63.7546
R19618 GND.n1 GND.t194 63.7546
R19619 GND.n48 GND.t180 63.7546
R19620 GND.n55 GND.t3 63.7546
R19621 GND.n63 GND.t200 63.7546
R19622 GND.n71 GND.t219 63.7546
R19623 GND.n79 GND.t205 63.7546
R19624 GND.n3767 GND.n3766 62.8652
R19625 GND.n2915 GND.t105 62.6855
R19626 GND.n8333 GND.t100 62.6855
R19627 GND.n8383 GND.t97 62.6855
R19628 GND.n8407 GND.t138 62.6855
R19629 GND.n2184 GND.t144 62.6855
R19630 GND.n4621 GND.t61 62.6855
R19631 GND.n4795 GND.t118 62.6855
R19632 GND.n4829 GND.t93 62.6855
R19633 GND.n10766 GND.t79 62.6855
R19634 GND.n10749 GND.t135 62.6855
R19635 GND.n10733 GND.t82 62.6855
R19636 GND.n457 GND.t103 62.6855
R19637 GND.n5887 GND.t121 62.6855
R19638 GND.n1744 GND.t127 62.6855
R19639 GND.n1760 GND.t71 62.6855
R19640 GND.n1777 GND.t124 62.6855
R19641 GND.n1795 GND.t84 62.6855
R19642 GND.n2144 GND.t48 62.6855
R19643 GND.n13 GND.t213 61.8897
R19644 GND.n20 GND.t231 61.8897
R19645 GND.n28 GND.t214 61.8897
R19646 GND.n36 GND.t172 61.8897
R19647 GND.n6 GND.t225 61.8897
R19648 GND.n53 GND.t184 61.8897
R19649 GND.n60 GND.t21 61.8897
R19650 GND.n68 GND.t173 61.8897
R19651 GND.n76 GND.t169 61.8897
R19652 GND.n84 GND.t44 61.8897
R19653 GND.n9044 GND.n1461 60.5899
R19654 GND.n9044 GND.n9043 60.5899
R19655 GND.n9043 GND.n9042 60.5899
R19656 GND.n9042 GND.n1466 60.5899
R19657 GND.n9036 GND.n1466 60.5899
R19658 GND.n9036 GND.n9035 60.5899
R19659 GND.n9035 GND.n9034 60.5899
R19660 GND.n9034 GND.n1474 60.5899
R19661 GND.n9028 GND.n1474 60.5899
R19662 GND.n9028 GND.n9027 60.5899
R19663 GND.n9027 GND.n9026 60.5899
R19664 GND.n9026 GND.n1482 60.5899
R19665 GND.n9020 GND.n1482 60.5899
R19666 GND.n9020 GND.n9019 60.5899
R19667 GND.n9019 GND.n9018 60.5899
R19668 GND.n9018 GND.n1490 60.5899
R19669 GND.n9012 GND.n1490 60.5899
R19670 GND.n9012 GND.n9011 60.5899
R19671 GND.n9011 GND.n9010 60.5899
R19672 GND.n9010 GND.n1498 60.5899
R19673 GND.n9004 GND.n1498 60.5899
R19674 GND.n9004 GND.n9003 60.5899
R19675 GND.n9003 GND.n9002 60.5899
R19676 GND.n9002 GND.n1506 60.5899
R19677 GND.n8996 GND.n1506 60.5899
R19678 GND.n8996 GND.n8995 60.5899
R19679 GND.n8995 GND.n8994 60.5899
R19680 GND.n8994 GND.n1514 60.5899
R19681 GND.n8988 GND.n1514 60.5899
R19682 GND.n8988 GND.n8987 60.5899
R19683 GND.n8987 GND.n8986 60.5899
R19684 GND.n8986 GND.n1522 60.5899
R19685 GND.n8980 GND.n1522 60.5899
R19686 GND.n8980 GND.n8979 60.5899
R19687 GND.n8979 GND.n8978 60.5899
R19688 GND.n8978 GND.n1530 60.5899
R19689 GND.n8972 GND.n1530 60.5899
R19690 GND.n8972 GND.n8971 60.5899
R19691 GND.n8971 GND.n8970 60.5899
R19692 GND.n8970 GND.n1538 60.5899
R19693 GND.n8964 GND.n1538 60.5899
R19694 GND.n8964 GND.n8963 60.5899
R19695 GND.n8963 GND.n8962 60.5899
R19696 GND.n8962 GND.n1546 60.5899
R19697 GND.n8956 GND.n1546 60.5899
R19698 GND.n8956 GND.n8955 60.5899
R19699 GND.n8955 GND.n8954 60.5899
R19700 GND.n8954 GND.n1554 60.5899
R19701 GND.n8948 GND.n1554 60.5899
R19702 GND.n8948 GND.n8947 60.5899
R19703 GND.n8947 GND.n8946 60.5899
R19704 GND.n8946 GND.n1562 60.5899
R19705 GND.n8940 GND.n1562 60.5899
R19706 GND.n8940 GND.n8939 60.5899
R19707 GND.n8939 GND.n8938 60.5899
R19708 GND.n8938 GND.n1570 60.5899
R19709 GND.n8932 GND.n1570 60.5899
R19710 GND.n8932 GND.n8931 60.5899
R19711 GND.n4811 GND.t55 59.4855
R19712 GND.n10785 GND.t76 59.4855
R19713 GND.n4644 GND.n4639 59.441
R19714 GND.n5057 GND.t140 54.9935
R19715 GND.n4656 GND.t68 54.9935
R19716 GND.n5066 GND.t131 54.9875
R19717 GND.n4636 GND.t52 54.9875
R19718 GND.n5132 GND.n5066 53.1399
R19719 GND.n5150 GND.n5057 53.1399
R19720 GND.n4664 GND.n4656 53.1399
R19721 GND.n4781 GND.n4636 53.1399
R19722 GND.n8 GND.n7 51.2731
R19723 GND.n10 GND.n9 51.2731
R19724 GND.n12 GND.n11 51.2731
R19725 GND.n15 GND.n14 51.2731
R19726 GND.n17 GND.n16 51.2731
R19727 GND.n19 GND.n18 51.2731
R19728 GND.n23 GND.n22 51.2731
R19729 GND.n25 GND.n24 51.2731
R19730 GND.n27 GND.n26 51.2731
R19731 GND.n31 GND.n30 51.2731
R19732 GND.n33 GND.n32 51.2731
R19733 GND.n35 GND.n34 51.2731
R19734 GND.n1 GND.n0 51.2731
R19735 GND.n3 GND.n2 51.2731
R19736 GND.n5 GND.n4 51.2731
R19737 GND.n52 GND.n51 51.2731
R19738 GND.n50 GND.n49 51.2731
R19739 GND.n48 GND.n47 51.2731
R19740 GND.n59 GND.n58 51.2731
R19741 GND.n57 GND.n56 51.2731
R19742 GND.n55 GND.n54 51.2731
R19743 GND.n67 GND.n66 51.2731
R19744 GND.n65 GND.n64 51.2731
R19745 GND.n63 GND.n62 51.2731
R19746 GND.n75 GND.n74 51.2731
R19747 GND.n73 GND.n72 51.2731
R19748 GND.n71 GND.n70 51.2731
R19749 GND.n83 GND.n82 51.2731
R19750 GND.n81 GND.n80 51.2731
R19751 GND.n79 GND.n78 51.2731
R19752 GND.n4812 GND.n4811 48.6793
R19753 GND.n10788 GND.n10785 48.6793
R19754 GND.n3763 GND.n3762 48.2005
R19755 GND.n4645 GND.n4638 48.2005
R19756 GND.n8014 GND.n8013 44.9944
R19757 GND.n5861 GND.n5860 44.9944
R19758 GND.n4649 GND.n4648 44.3322
R19759 GND.n3760 GND.n3759 41.6274
R19760 GND.n4643 GND.n4642 41.6274
R19761 GND.n3762 GND.n3761 36.5361
R19762 GND.n8015 GND.n8014 36.0732
R19763 GND.n5863 GND.n5861 36.0732
R19764 GND.n2947 GND.n2915 35.8793
R19765 GND.n8336 GND.n8333 35.8793
R19766 GND.n8384 GND.n8383 35.8793
R19767 GND.n8412 GND.n8407 35.8793
R19768 GND.n7623 GND.n4621 35.8793
R19769 GND.n7539 GND.n4829 35.8793
R19770 GND.n10767 GND.n10766 35.8793
R19771 GND.n10750 GND.n10749 35.8793
R19772 GND.n10875 GND.n10733 35.8793
R19773 GND.n458 GND.n457 35.8793
R19774 GND.n5888 GND.n5887 35.8793
R19775 GND.n8792 GND.n1744 35.8793
R19776 GND.n1761 GND.n1760 35.8793
R19777 GND.n1778 GND.n1777 35.8793
R19778 GND.n8706 GND.n1795 35.8793
R19779 GND.n8460 GND.n2144 35.8793
R19780 GND.n8930 GND.n1578 33.4453
R19781 GND.n1587 GND.n1578 33.4453
R19782 GND.n8921 GND.n1587 33.4453
R19783 GND.n8921 GND.n8920 33.4453
R19784 GND.n8920 GND.n8919 33.4453
R19785 GND.n8919 GND.n1588 33.4453
R19786 GND.n8913 GND.n1588 33.4453
R19787 GND.n8913 GND.n8912 33.4453
R19788 GND.n8912 GND.n8911 33.4453
R19789 GND.n8911 GND.n1595 33.4453
R19790 GND.n8905 GND.n1595 33.4453
R19791 GND.n8905 GND.n8904 33.4453
R19792 GND.n8904 GND.n8903 33.4453
R19793 GND.n8903 GND.n1603 33.4453
R19794 GND.n8897 GND.n1603 33.4453
R19795 GND.n8897 GND.n8896 33.4453
R19796 GND.n8896 GND.n8895 33.4453
R19797 GND.n8895 GND.n1611 33.4453
R19798 GND.n8889 GND.n1611 33.4453
R19799 GND.n8889 GND.n8888 33.4453
R19800 GND.n8888 GND.n8887 33.4453
R19801 GND.n8887 GND.n1619 33.4453
R19802 GND.n8881 GND.n1619 33.4453
R19803 GND.n8881 GND.n8880 33.4453
R19804 GND.n8880 GND.n8879 33.4453
R19805 GND.n8879 GND.n1627 33.4453
R19806 GND.n8873 GND.n1627 33.4453
R19807 GND.n8873 GND.n8872 33.4453
R19808 GND.n8872 GND.n8871 33.4453
R19809 GND.n8871 GND.n1635 33.4453
R19810 GND.n8865 GND.n1635 33.4453
R19811 GND.n8865 GND.n8864 33.4453
R19812 GND.n8864 GND.n8863 33.4453
R19813 GND.n8863 GND.n1643 33.4453
R19814 GND.n8857 GND.n1643 33.4453
R19815 GND.n8857 GND.n8856 33.4453
R19816 GND.n8856 GND.n8855 33.4453
R19817 GND.n8855 GND.n1651 33.4453
R19818 GND.n8849 GND.n1651 33.4453
R19819 GND.n8849 GND.n8848 33.4453
R19820 GND.n8848 GND.n8847 33.4453
R19821 GND.n8847 GND.n1659 33.4453
R19822 GND.n8841 GND.n1659 33.4453
R19823 GND.n8841 GND.n8840 33.4453
R19824 GND.n8840 GND.n8839 33.4453
R19825 GND.n8839 GND.n1667 33.4453
R19826 GND.n8833 GND.n1667 33.4453
R19827 GND.n8833 GND.n8832 33.4453
R19828 GND.n8832 GND.n8831 33.4453
R19829 GND.n8831 GND.n1675 33.4453
R19830 GND.n8825 GND.n1675 33.4453
R19831 GND.n8825 GND.n8824 33.4453
R19832 GND.n8824 GND.n8823 33.4453
R19833 GND.n8823 GND.n1683 33.4453
R19834 GND.n8817 GND.n1683 33.4453
R19835 GND.n1801 GND.n1725 33.4453
R19836 GND.n2147 GND.n2128 33.4453
R19837 GND.n8135 GND.n2166 33.4453
R19838 GND.n8135 GND.n8134 33.4453
R19839 GND.n8134 GND.n8133 33.4453
R19840 GND.n8133 GND.n3739 33.4453
R19841 GND.n7655 GND.n4560 33.4453
R19842 GND.n7649 GND.n4560 33.4453
R19843 GND.n7649 GND.n7648 33.4453
R19844 GND.n5879 GND.n4602 33.4453
R19845 GND.n460 GND.n448 33.4453
R19846 GND.n10646 GND.n461 33.4453
R19847 GND.n10640 GND.n461 33.4453
R19848 GND.n10640 GND.n10639 33.4453
R19849 GND.n10639 GND.n10638 33.4453
R19850 GND.n10638 GND.n470 33.4453
R19851 GND.n10632 GND.n470 33.4453
R19852 GND.n10632 GND.n10631 33.4453
R19853 GND.n10631 GND.n10630 33.4453
R19854 GND.n10630 GND.n478 33.4453
R19855 GND.n10624 GND.n478 33.4453
R19856 GND.n10624 GND.n10623 33.4453
R19857 GND.n10623 GND.n10622 33.4453
R19858 GND.n10622 GND.n486 33.4453
R19859 GND.n10616 GND.n486 33.4453
R19860 GND.n10616 GND.n10615 33.4453
R19861 GND.n10615 GND.n10614 33.4453
R19862 GND.n10614 GND.n494 33.4453
R19863 GND.n10608 GND.n494 33.4453
R19864 GND.n10608 GND.n10607 33.4453
R19865 GND.n10607 GND.n10606 33.4453
R19866 GND.n10606 GND.n502 33.4453
R19867 GND.n10600 GND.n502 33.4453
R19868 GND.n10600 GND.n10599 33.4453
R19869 GND.n10599 GND.n10598 33.4453
R19870 GND.n10598 GND.n510 33.4453
R19871 GND.n10592 GND.n510 33.4453
R19872 GND.n10592 GND.n10591 33.4453
R19873 GND.n10591 GND.n10590 33.4453
R19874 GND.n10590 GND.n518 33.4453
R19875 GND.n10584 GND.n518 33.4453
R19876 GND.n10584 GND.n10583 33.4453
R19877 GND.n10583 GND.n10582 33.4453
R19878 GND.n10582 GND.n526 33.4453
R19879 GND.n10576 GND.n526 33.4453
R19880 GND.n10576 GND.n10575 33.4453
R19881 GND.n10575 GND.n10574 33.4453
R19882 GND.n10574 GND.n534 33.4453
R19883 GND.n10568 GND.n534 33.4453
R19884 GND.n10568 GND.n10567 33.4453
R19885 GND.n10567 GND.n10566 33.4453
R19886 GND.n10566 GND.n542 33.4453
R19887 GND.n10560 GND.n542 33.4453
R19888 GND.n10560 GND.n10559 33.4453
R19889 GND.n10559 GND.n10558 33.4453
R19890 GND.n10558 GND.n550 33.4453
R19891 GND.n10552 GND.n550 33.4453
R19892 GND.n10552 GND.n10551 33.4453
R19893 GND.n10551 GND.n10550 33.4453
R19894 GND.n10550 GND.n558 33.4453
R19895 GND.n10544 GND.n558 33.4453
R19896 GND.n10544 GND.n10543 33.4453
R19897 GND.n10543 GND.n10542 33.4453
R19898 GND.n10542 GND.n566 33.4453
R19899 GND.n10536 GND.n566 33.4453
R19900 GND.n10536 GND.n10535 33.4453
R19901 GND.n4719 GND.n4718 32.6249
R19902 GND.n5205 GND.n5204 32.6249
R19903 GND.n8127 GND.n3749 32.442
R19904 GND.n7658 GND.n7657 32.442
R19905 GND.n5141 GND.n2185 30.5925
R19906 GND.n7597 GND.n4791 30.5925
R19907 GND.n2185 GND.n2184 30.5518
R19908 GND.n7597 GND.n4795 30.5518
R19909 GND.t58 GND.n7655 29.4319
R19910 GND.n3764 GND.n3763 27.0217
R19911 GND.n4646 GND.n4645 27.0217
R19912 GND.n3756 GND.n3755 25.8289
R19913 GND.n8817 GND.n8816 25.0841
R19914 GND.n8457 GND.n2166 25.0841
R19915 GND.n7648 GND.n7647 25.0841
R19916 GND.n10896 GND.n10646 25.0841
R19917 GND.n8126 GND.n3751 22.743
R19918 GND.n5214 GND.n3772 22.743
R19919 GND.n8112 GND.t64 22.743
R19920 GND.n8106 GND.t64 22.743
R19921 GND.n5227 GND.n3796 22.743
R19922 GND.n8092 GND.n3804 22.743
R19923 GND.n5240 GND.n3814 22.743
R19924 GND.n8078 GND.n3822 22.743
R19925 GND.n5253 GND.n3832 22.743
R19926 GND.n8064 GND.n3840 22.743
R19927 GND.n5305 GND.n3850 22.743
R19928 GND.n8005 GND.n3882 22.743
R19929 GND.n8005 GND.n3884 22.743
R19930 GND.n5030 GND.n3895 22.743
R19931 GND.n5342 GND.n3916 22.743
R19932 GND.n5352 GND.n3926 22.743
R19933 GND.n5361 GND.n3936 22.743
R19934 GND.n5421 GND.n3956 22.743
R19935 GND.n5430 GND.n3966 22.743
R19936 GND.n5430 GND.n3974 22.743
R19937 GND.n5439 GND.n3984 22.743
R19938 GND.n5448 GND.n3994 22.743
R19939 GND.n5457 GND.n4004 22.743
R19940 GND.n5466 GND.n4014 22.743
R19941 GND.n5475 GND.n4024 22.743
R19942 GND.n5503 GND.n4044 22.743
R19943 GND.n7903 GND.n4054 22.743
R19944 GND.n7903 GND.n4057 22.743
R19945 GND.n7891 GND.n4071 22.743
R19946 GND.n5560 GND.n4109 22.743
R19947 GND.n5569 GND.n4119 22.743
R19948 GND.n5578 GND.n4129 22.743
R19949 GND.n5606 GND.n4149 22.743
R19950 GND.n7848 GND.n4159 22.743
R19951 GND.n7848 GND.n4162 22.743
R19952 GND.n7836 GND.n4176 22.743
R19953 GND.n5664 GND.n4213 22.743
R19954 GND.n5673 GND.n4223 22.743
R19955 GND.n5683 GND.n4233 22.743
R19956 GND.n5697 GND.n4899 22.743
R19957 GND.n5709 GND.n4251 22.743
R19958 GND.n7793 GND.n4261 22.743
R19959 GND.n7793 GND.n4264 22.743
R19960 GND.n7781 GND.n4278 22.743
R19961 GND.n5761 GND.n4316 22.743
R19962 GND.n5770 GND.n4326 22.743
R19963 GND.n5778 GND.n4336 22.743
R19964 GND.n5792 GND.n4355 22.743
R19965 GND.n7738 GND.n4365 22.743
R19966 GND.n7738 GND.n4368 22.743
R19967 GND.n7726 GND.n4382 22.743
R19968 GND.n4463 GND.n4396 22.743
R19969 GND.n7712 GND.n4404 22.743
R19970 GND.n4476 GND.n4414 22.743
R19971 GND.n7698 GND.n4422 22.743
R19972 GND.n4489 GND.n4432 22.743
R19973 GND.n7684 GND.n4440 22.743
R19974 GND.n7677 GND.n4449 22.743
R19975 GND.n7677 GND.n4451 22.743
R19976 GND.n7665 GND.n4514 22.743
R19977 GND.n7999 GND.n3893 21.4052
R19978 GND.n4997 GND.n3964 21.4052
R19979 GND.n4987 GND.n3976 21.4052
R19980 GND.n7909 GND.n4046 21.4052
R19981 GND.n7897 GND.n4065 21.4052
R19982 GND.n7854 GND.n4151 21.4052
R19983 GND.n7842 GND.n4170 21.4052
R19984 GND.n7799 GND.n4253 21.4052
R19985 GND.n7787 GND.n4272 21.4052
R19986 GND.n7744 GND.n4357 21.4052
R19987 GND.n7671 GND.n4505 21.4052
R19988 GND.n3765 GND.n3764 21.1793
R19989 GND.n4647 GND.n4646 21.1793
R19990 GND.n8120 GND.n3770 20.0674
R19991 GND.n8098 GND.n3798 20.0674
R19992 GND.n8063 GND.n3842 20.0674
R19993 GND.n5411 GND.n3954 20.0674
R19994 GND.n7915 GND.n4036 20.0674
R19995 GND.n5542 GND.n4074 20.0674
R19996 GND.n7860 GND.n4141 20.0674
R19997 GND.n5646 GND.n4179 20.0674
R19998 GND.n5743 GND.n4281 20.0674
R19999 GND.n4460 GND.n4384 20.0674
R20000 GND.n7691 GND.n7690 20.0674
R20001 GND.n4650 GND.n4516 20.0674
R20002 GND.n3758 GND.t112 19.8005
R20003 GND.n3758 GND.t151 19.8005
R20004 GND.n3757 GND.t91 19.8005
R20005 GND.n3757 GND.t65 19.8005
R20006 GND.n4641 GND.t88 19.8005
R20007 GND.n4641 GND.t154 19.8005
R20008 GND.n4640 GND.t109 19.8005
R20009 GND.n4640 GND.t59 19.8005
R20010 GND.n3755 GND.n3754 19.5087
R20011 GND.t130 GND.n3788 19.3985
R20012 GND.n5333 GND.t155 19.3985
R20013 GND.n5800 GND.t15 19.3985
R20014 GND.n4498 GND.t50 19.3985
R20015 GND.n2953 GND.n2911 19.3944
R20016 GND.n2956 GND.n2953 19.3944
R20017 GND.n2957 GND.n2956 19.3944
R20018 GND.n2957 GND.n2909 19.3944
R20019 GND.n2961 GND.n2909 19.3944
R20020 GND.n2962 GND.n2961 19.3944
R20021 GND.n3162 GND.n2962 19.3944
R20022 GND.n3162 GND.n2903 19.3944
R20023 GND.n3167 GND.n2903 19.3944
R20024 GND.n3167 GND.n2904 19.3944
R20025 GND.n2904 GND.n2884 19.3944
R20026 GND.n3187 GND.n2884 19.3944
R20027 GND.n3187 GND.n2881 19.3944
R20028 GND.n3192 GND.n2881 19.3944
R20029 GND.n3192 GND.n2882 19.3944
R20030 GND.n2882 GND.n2862 19.3944
R20031 GND.n3212 GND.n2862 19.3944
R20032 GND.n3212 GND.n2859 19.3944
R20033 GND.n3217 GND.n2859 19.3944
R20034 GND.n3217 GND.n2860 19.3944
R20035 GND.n2860 GND.n2838 19.3944
R20036 GND.n3236 GND.n2838 19.3944
R20037 GND.n3236 GND.n2835 19.3944
R20038 GND.n3241 GND.n2835 19.3944
R20039 GND.n3241 GND.n2836 19.3944
R20040 GND.n2836 GND.n2815 19.3944
R20041 GND.n3261 GND.n2815 19.3944
R20042 GND.n3261 GND.n2812 19.3944
R20043 GND.n3266 GND.n2812 19.3944
R20044 GND.n3266 GND.n2813 19.3944
R20045 GND.n2813 GND.n2793 19.3944
R20046 GND.n3286 GND.n2793 19.3944
R20047 GND.n3286 GND.n2790 19.3944
R20048 GND.n3291 GND.n2790 19.3944
R20049 GND.n3291 GND.n2791 19.3944
R20050 GND.n2791 GND.n2771 19.3944
R20051 GND.n3311 GND.n2771 19.3944
R20052 GND.n3311 GND.n2768 19.3944
R20053 GND.n3316 GND.n2768 19.3944
R20054 GND.n3316 GND.n2769 19.3944
R20055 GND.n2769 GND.n2747 19.3944
R20056 GND.n3335 GND.n2747 19.3944
R20057 GND.n3335 GND.n2744 19.3944
R20058 GND.n3340 GND.n2744 19.3944
R20059 GND.n3340 GND.n2745 19.3944
R20060 GND.n2745 GND.n2724 19.3944
R20061 GND.n3360 GND.n2724 19.3944
R20062 GND.n3360 GND.n2721 19.3944
R20063 GND.n3365 GND.n2721 19.3944
R20064 GND.n3365 GND.n2722 19.3944
R20065 GND.n2722 GND.n2702 19.3944
R20066 GND.n3385 GND.n2702 19.3944
R20067 GND.n3385 GND.n2699 19.3944
R20068 GND.n3390 GND.n2699 19.3944
R20069 GND.n3390 GND.n2700 19.3944
R20070 GND.n2700 GND.n2680 19.3944
R20071 GND.n3410 GND.n2680 19.3944
R20072 GND.n3410 GND.n2677 19.3944
R20073 GND.n3415 GND.n2677 19.3944
R20074 GND.n3415 GND.n2678 19.3944
R20075 GND.n2678 GND.n2658 19.3944
R20076 GND.n3432 GND.n2658 19.3944
R20077 GND.n3432 GND.n2656 19.3944
R20078 GND.n3436 GND.n2656 19.3944
R20079 GND.n3437 GND.n3436 19.3944
R20080 GND.n3440 GND.n3437 19.3944
R20081 GND.n3440 GND.n2654 19.3944
R20082 GND.n3445 GND.n2654 19.3944
R20083 GND.n3446 GND.n3445 19.3944
R20084 GND.n3447 GND.n3446 19.3944
R20085 GND.n3447 GND.n2652 19.3944
R20086 GND.n3451 GND.n2652 19.3944
R20087 GND.n3451 GND.n2481 19.3944
R20088 GND.n3502 GND.n2481 19.3944
R20089 GND.n3502 GND.n2479 19.3944
R20090 GND.n3508 GND.n2479 19.3944
R20091 GND.n3508 GND.n3507 19.3944
R20092 GND.n3507 GND.n2459 19.3944
R20093 GND.n3528 GND.n2459 19.3944
R20094 GND.n3528 GND.n2457 19.3944
R20095 GND.n3534 GND.n2457 19.3944
R20096 GND.n3534 GND.n3533 19.3944
R20097 GND.n3533 GND.n2438 19.3944
R20098 GND.n3554 GND.n2438 19.3944
R20099 GND.n3554 GND.n2436 19.3944
R20100 GND.n3560 GND.n2436 19.3944
R20101 GND.n3560 GND.n3559 19.3944
R20102 GND.n3559 GND.n2417 19.3944
R20103 GND.n3580 GND.n2417 19.3944
R20104 GND.n3580 GND.n2415 19.3944
R20105 GND.n3586 GND.n2415 19.3944
R20106 GND.n3586 GND.n3585 19.3944
R20107 GND.n3585 GND.n2394 19.3944
R20108 GND.n3605 GND.n2394 19.3944
R20109 GND.n3605 GND.n2392 19.3944
R20110 GND.n3611 GND.n2392 19.3944
R20111 GND.n3611 GND.n3610 19.3944
R20112 GND.n3610 GND.n2374 19.3944
R20113 GND.n3631 GND.n2374 19.3944
R20114 GND.n3631 GND.n2372 19.3944
R20115 GND.n3637 GND.n2372 19.3944
R20116 GND.n3637 GND.n3636 19.3944
R20117 GND.n3636 GND.n2354 19.3944
R20118 GND.n3657 GND.n2354 19.3944
R20119 GND.n3657 GND.n2352 19.3944
R20120 GND.n3663 GND.n2352 19.3944
R20121 GND.n3663 GND.n3662 19.3944
R20122 GND.n3662 GND.n2332 19.3944
R20123 GND.n3683 GND.n2332 19.3944
R20124 GND.n3683 GND.n2330 19.3944
R20125 GND.n3689 GND.n2330 19.3944
R20126 GND.n3689 GND.n3688 19.3944
R20127 GND.n3688 GND.n2305 19.3944
R20128 GND.n8194 GND.n2305 19.3944
R20129 GND.n8194 GND.n2303 19.3944
R20130 GND.n8200 GND.n2303 19.3944
R20131 GND.n8200 GND.n8199 19.3944
R20132 GND.n8199 GND.n2283 19.3944
R20133 GND.n8220 GND.n2283 19.3944
R20134 GND.n8220 GND.n2281 19.3944
R20135 GND.n8226 GND.n2281 19.3944
R20136 GND.n8226 GND.n8225 19.3944
R20137 GND.n8225 GND.n2262 19.3944
R20138 GND.n8246 GND.n2262 19.3944
R20139 GND.n8246 GND.n2260 19.3944
R20140 GND.n8252 GND.n2260 19.3944
R20141 GND.n8252 GND.n8251 19.3944
R20142 GND.n8251 GND.n2241 19.3944
R20143 GND.n8272 GND.n2241 19.3944
R20144 GND.n8272 GND.n2239 19.3944
R20145 GND.n8278 GND.n2239 19.3944
R20146 GND.n8278 GND.n8277 19.3944
R20147 GND.n8277 GND.n2218 19.3944
R20148 GND.n8296 GND.n2218 19.3944
R20149 GND.n8296 GND.n2216 19.3944
R20150 GND.n8302 GND.n2216 19.3944
R20151 GND.n8302 GND.n8301 19.3944
R20152 GND.n8701 GND.n1798 19.3944
R20153 GND.n2923 GND.n1798 19.3944
R20154 GND.n2926 GND.n2923 19.3944
R20155 GND.n2929 GND.n2926 19.3944
R20156 GND.n2932 GND.n2929 19.3944
R20157 GND.n2932 GND.n2919 19.3944
R20158 GND.n2936 GND.n2919 19.3944
R20159 GND.n2939 GND.n2936 19.3944
R20160 GND.n2942 GND.n2939 19.3944
R20161 GND.n2942 GND.n2916 19.3944
R20162 GND.n2946 GND.n2916 19.3944
R20163 GND.n1851 GND.n1848 19.3944
R20164 GND.n1851 GND.n1846 19.3944
R20165 GND.n1858 GND.n1846 19.3944
R20166 GND.n1859 GND.n1858 19.3944
R20167 GND.n8680 GND.n1859 19.3944
R20168 GND.n8680 GND.n8679 19.3944
R20169 GND.n8679 GND.n8678 19.3944
R20170 GND.n8678 GND.n1862 19.3944
R20171 GND.n8674 GND.n1862 19.3944
R20172 GND.n8674 GND.n8673 19.3944
R20173 GND.n8673 GND.n8672 19.3944
R20174 GND.n8672 GND.n1870 19.3944
R20175 GND.n8668 GND.n1870 19.3944
R20176 GND.n8668 GND.n8667 19.3944
R20177 GND.n8667 GND.n8666 19.3944
R20178 GND.n8666 GND.n1878 19.3944
R20179 GND.n8662 GND.n1878 19.3944
R20180 GND.n8662 GND.n8661 19.3944
R20181 GND.n8661 GND.n8660 19.3944
R20182 GND.n8660 GND.n1886 19.3944
R20183 GND.n8656 GND.n1886 19.3944
R20184 GND.n8656 GND.n8655 19.3944
R20185 GND.n8655 GND.n8654 19.3944
R20186 GND.n8654 GND.n1894 19.3944
R20187 GND.n8650 GND.n1894 19.3944
R20188 GND.n8650 GND.n8649 19.3944
R20189 GND.n8649 GND.n8648 19.3944
R20190 GND.n8648 GND.n1902 19.3944
R20191 GND.n8644 GND.n1902 19.3944
R20192 GND.n8644 GND.n8643 19.3944
R20193 GND.n8643 GND.n8642 19.3944
R20194 GND.n8642 GND.n1910 19.3944
R20195 GND.n8638 GND.n1910 19.3944
R20196 GND.n8638 GND.n8637 19.3944
R20197 GND.n8637 GND.n8636 19.3944
R20198 GND.n8636 GND.n1918 19.3944
R20199 GND.n8632 GND.n1918 19.3944
R20200 GND.n8632 GND.n8631 19.3944
R20201 GND.n8631 GND.n8630 19.3944
R20202 GND.n8630 GND.n1926 19.3944
R20203 GND.n8626 GND.n1926 19.3944
R20204 GND.n8626 GND.n8625 19.3944
R20205 GND.n8625 GND.n8624 19.3944
R20206 GND.n8624 GND.n1934 19.3944
R20207 GND.n8620 GND.n1934 19.3944
R20208 GND.n8620 GND.n8619 19.3944
R20209 GND.n8619 GND.n8618 19.3944
R20210 GND.n8618 GND.n1942 19.3944
R20211 GND.n8614 GND.n1942 19.3944
R20212 GND.n8614 GND.n8613 19.3944
R20213 GND.n8613 GND.n8612 19.3944
R20214 GND.n8612 GND.n1950 19.3944
R20215 GND.n8608 GND.n1950 19.3944
R20216 GND.n8608 GND.n8607 19.3944
R20217 GND.n8607 GND.n8606 19.3944
R20218 GND.n8606 GND.n1958 19.3944
R20219 GND.n8602 GND.n1958 19.3944
R20220 GND.n8602 GND.n8601 19.3944
R20221 GND.n8601 GND.n8600 19.3944
R20222 GND.n8600 GND.n1966 19.3944
R20223 GND.n8596 GND.n1966 19.3944
R20224 GND.n8596 GND.n8595 19.3944
R20225 GND.n8595 GND.n8594 19.3944
R20226 GND.n8594 GND.n1974 19.3944
R20227 GND.n8590 GND.n1974 19.3944
R20228 GND.n8590 GND.n8589 19.3944
R20229 GND.n8589 GND.n8588 19.3944
R20230 GND.n8588 GND.n1982 19.3944
R20231 GND.n8584 GND.n1982 19.3944
R20232 GND.n8584 GND.n8583 19.3944
R20233 GND.n8583 GND.n8582 19.3944
R20234 GND.n8582 GND.n1990 19.3944
R20235 GND.n8578 GND.n1990 19.3944
R20236 GND.n8578 GND.n8577 19.3944
R20237 GND.n8577 GND.n8576 19.3944
R20238 GND.n8576 GND.n1998 19.3944
R20239 GND.n8572 GND.n1998 19.3944
R20240 GND.n8572 GND.n8571 19.3944
R20241 GND.n8571 GND.n8570 19.3944
R20242 GND.n8570 GND.n2006 19.3944
R20243 GND.n8566 GND.n2006 19.3944
R20244 GND.n8566 GND.n8565 19.3944
R20245 GND.n8565 GND.n8564 19.3944
R20246 GND.n8564 GND.n2014 19.3944
R20247 GND.n8560 GND.n2014 19.3944
R20248 GND.n8560 GND.n8559 19.3944
R20249 GND.n8559 GND.n8558 19.3944
R20250 GND.n8558 GND.n2022 19.3944
R20251 GND.n8554 GND.n2022 19.3944
R20252 GND.n8554 GND.n8553 19.3944
R20253 GND.n8553 GND.n8552 19.3944
R20254 GND.n8552 GND.n2030 19.3944
R20255 GND.n8548 GND.n2030 19.3944
R20256 GND.n8548 GND.n8547 19.3944
R20257 GND.n8547 GND.n8546 19.3944
R20258 GND.n8546 GND.n2038 19.3944
R20259 GND.n8542 GND.n2038 19.3944
R20260 GND.n8542 GND.n8541 19.3944
R20261 GND.n8541 GND.n8540 19.3944
R20262 GND.n8540 GND.n2046 19.3944
R20263 GND.n8536 GND.n2046 19.3944
R20264 GND.n8536 GND.n8535 19.3944
R20265 GND.n8535 GND.n8534 19.3944
R20266 GND.n8534 GND.n2054 19.3944
R20267 GND.n8530 GND.n2054 19.3944
R20268 GND.n8530 GND.n8529 19.3944
R20269 GND.n8529 GND.n8528 19.3944
R20270 GND.n8528 GND.n2062 19.3944
R20271 GND.n8524 GND.n2062 19.3944
R20272 GND.n8524 GND.n8523 19.3944
R20273 GND.n8523 GND.n8522 19.3944
R20274 GND.n8522 GND.n2070 19.3944
R20275 GND.n8518 GND.n2070 19.3944
R20276 GND.n8518 GND.n8517 19.3944
R20277 GND.n8517 GND.n8516 19.3944
R20278 GND.n8516 GND.n2078 19.3944
R20279 GND.n8512 GND.n2078 19.3944
R20280 GND.n8512 GND.n8511 19.3944
R20281 GND.n8511 GND.n8510 19.3944
R20282 GND.n8510 GND.n2086 19.3944
R20283 GND.n8506 GND.n2086 19.3944
R20284 GND.n8506 GND.n8505 19.3944
R20285 GND.n8505 GND.n8504 19.3944
R20286 GND.n8504 GND.n2094 19.3944
R20287 GND.n8500 GND.n2094 19.3944
R20288 GND.n8500 GND.n8499 19.3944
R20289 GND.n8499 GND.n8498 19.3944
R20290 GND.n8498 GND.n2102 19.3944
R20291 GND.n8494 GND.n2102 19.3944
R20292 GND.n8494 GND.n8493 19.3944
R20293 GND.n8493 GND.n8492 19.3944
R20294 GND.n8492 GND.n2110 19.3944
R20295 GND.n8488 GND.n2110 19.3944
R20296 GND.n8488 GND.n8487 19.3944
R20297 GND.n8487 GND.n8486 19.3944
R20298 GND.n8486 GND.n2118 19.3944
R20299 GND.n8482 GND.n2118 19.3944
R20300 GND.n8310 GND.n2208 19.3944
R20301 GND.n8314 GND.n2208 19.3944
R20302 GND.n8315 GND.n8314 19.3944
R20303 GND.n8318 GND.n8315 19.3944
R20304 GND.n8318 GND.n2204 19.3944
R20305 GND.n8322 GND.n2204 19.3944
R20306 GND.n8323 GND.n8322 19.3944
R20307 GND.n8326 GND.n8323 19.3944
R20308 GND.n8326 GND.n2200 19.3944
R20309 GND.n8330 GND.n2200 19.3944
R20310 GND.n8331 GND.n8330 19.3944
R20311 GND.n8340 GND.n2196 19.3944
R20312 GND.n8341 GND.n8340 19.3944
R20313 GND.n8344 GND.n8341 19.3944
R20314 GND.n8344 GND.n2192 19.3944
R20315 GND.n8348 GND.n2192 19.3944
R20316 GND.n8349 GND.n8348 19.3944
R20317 GND.n8352 GND.n8349 19.3944
R20318 GND.n8352 GND.n2188 19.3944
R20319 GND.n8356 GND.n2188 19.3944
R20320 GND.n8357 GND.n8356 19.3944
R20321 GND.n8360 GND.n8357 19.3944
R20322 GND.n8454 GND.n2186 19.3944
R20323 GND.n8450 GND.n2186 19.3944
R20324 GND.n8450 GND.n8449 19.3944
R20325 GND.n8449 GND.n8448 19.3944
R20326 GND.n8448 GND.n8368 19.3944
R20327 GND.n8444 GND.n8368 19.3944
R20328 GND.n8444 GND.n8443 19.3944
R20329 GND.n8443 GND.n8442 19.3944
R20330 GND.n8442 GND.n8374 19.3944
R20331 GND.n8438 GND.n8374 19.3944
R20332 GND.n8438 GND.n8437 19.3944
R20333 GND.n8437 GND.n8436 19.3944
R20334 GND.n8436 GND.n8380 19.3944
R20335 GND.n8432 GND.n8431 19.3944
R20336 GND.n8431 GND.n8430 19.3944
R20337 GND.n8430 GND.n8389 19.3944
R20338 GND.n8426 GND.n8389 19.3944
R20339 GND.n8426 GND.n8425 19.3944
R20340 GND.n8425 GND.n8424 19.3944
R20341 GND.n8424 GND.n8395 19.3944
R20342 GND.n8420 GND.n8395 19.3944
R20343 GND.n8420 GND.n8419 19.3944
R20344 GND.n8419 GND.n8418 19.3944
R20345 GND.n8418 GND.n8401 19.3944
R20346 GND.n8414 GND.n8401 19.3944
R20347 GND.n8414 GND.n8413 19.3944
R20348 GND.n10387 GND.n660 19.3944
R20349 GND.n10391 GND.n660 19.3944
R20350 GND.n10391 GND.n656 19.3944
R20351 GND.n10397 GND.n656 19.3944
R20352 GND.n10397 GND.n654 19.3944
R20353 GND.n10401 GND.n654 19.3944
R20354 GND.n10401 GND.n650 19.3944
R20355 GND.n10407 GND.n650 19.3944
R20356 GND.n10407 GND.n648 19.3944
R20357 GND.n10411 GND.n648 19.3944
R20358 GND.n10411 GND.n644 19.3944
R20359 GND.n10417 GND.n644 19.3944
R20360 GND.n10417 GND.n642 19.3944
R20361 GND.n10421 GND.n642 19.3944
R20362 GND.n10421 GND.n638 19.3944
R20363 GND.n10427 GND.n638 19.3944
R20364 GND.n10427 GND.n636 19.3944
R20365 GND.n10431 GND.n636 19.3944
R20366 GND.n10431 GND.n632 19.3944
R20367 GND.n10437 GND.n632 19.3944
R20368 GND.n10437 GND.n630 19.3944
R20369 GND.n10441 GND.n630 19.3944
R20370 GND.n10441 GND.n626 19.3944
R20371 GND.n10447 GND.n626 19.3944
R20372 GND.n10447 GND.n624 19.3944
R20373 GND.n10451 GND.n624 19.3944
R20374 GND.n10451 GND.n620 19.3944
R20375 GND.n10457 GND.n620 19.3944
R20376 GND.n10457 GND.n618 19.3944
R20377 GND.n10461 GND.n618 19.3944
R20378 GND.n10461 GND.n614 19.3944
R20379 GND.n10467 GND.n614 19.3944
R20380 GND.n10467 GND.n612 19.3944
R20381 GND.n10471 GND.n612 19.3944
R20382 GND.n10471 GND.n608 19.3944
R20383 GND.n10477 GND.n608 19.3944
R20384 GND.n10477 GND.n606 19.3944
R20385 GND.n10481 GND.n606 19.3944
R20386 GND.n10481 GND.n602 19.3944
R20387 GND.n10487 GND.n602 19.3944
R20388 GND.n10487 GND.n600 19.3944
R20389 GND.n10491 GND.n600 19.3944
R20390 GND.n10491 GND.n596 19.3944
R20391 GND.n10497 GND.n596 19.3944
R20392 GND.n10497 GND.n594 19.3944
R20393 GND.n10501 GND.n594 19.3944
R20394 GND.n10501 GND.n590 19.3944
R20395 GND.n10507 GND.n590 19.3944
R20396 GND.n10507 GND.n588 19.3944
R20397 GND.n10511 GND.n588 19.3944
R20398 GND.n10511 GND.n584 19.3944
R20399 GND.n10517 GND.n584 19.3944
R20400 GND.n10517 GND.n582 19.3944
R20401 GND.n10521 GND.n582 19.3944
R20402 GND.n10521 GND.n578 19.3944
R20403 GND.n10527 GND.n578 19.3944
R20404 GND.n10527 GND.n576 19.3944
R20405 GND.n10532 GND.n576 19.3944
R20406 GND.n9050 GND.n1459 19.3944
R20407 GND.n9056 GND.n1459 19.3944
R20408 GND.n9056 GND.n1457 19.3944
R20409 GND.n9060 GND.n1457 19.3944
R20410 GND.n9060 GND.n1453 19.3944
R20411 GND.n9066 GND.n1453 19.3944
R20412 GND.n9066 GND.n1451 19.3944
R20413 GND.n9070 GND.n1451 19.3944
R20414 GND.n9070 GND.n1447 19.3944
R20415 GND.n9076 GND.n1447 19.3944
R20416 GND.n9076 GND.n1445 19.3944
R20417 GND.n9080 GND.n1445 19.3944
R20418 GND.n9080 GND.n1441 19.3944
R20419 GND.n9086 GND.n1441 19.3944
R20420 GND.n9086 GND.n1439 19.3944
R20421 GND.n9090 GND.n1439 19.3944
R20422 GND.n9090 GND.n1435 19.3944
R20423 GND.n9096 GND.n1435 19.3944
R20424 GND.n9096 GND.n1433 19.3944
R20425 GND.n9100 GND.n1433 19.3944
R20426 GND.n9100 GND.n1429 19.3944
R20427 GND.n9106 GND.n1429 19.3944
R20428 GND.n9106 GND.n1427 19.3944
R20429 GND.n9110 GND.n1427 19.3944
R20430 GND.n9110 GND.n1423 19.3944
R20431 GND.n9116 GND.n1423 19.3944
R20432 GND.n9116 GND.n1421 19.3944
R20433 GND.n9120 GND.n1421 19.3944
R20434 GND.n9120 GND.n1417 19.3944
R20435 GND.n9126 GND.n1417 19.3944
R20436 GND.n9126 GND.n1415 19.3944
R20437 GND.n9130 GND.n1415 19.3944
R20438 GND.n9130 GND.n1411 19.3944
R20439 GND.n9136 GND.n1411 19.3944
R20440 GND.n9136 GND.n1409 19.3944
R20441 GND.n9140 GND.n1409 19.3944
R20442 GND.n9140 GND.n1405 19.3944
R20443 GND.n9146 GND.n1405 19.3944
R20444 GND.n9146 GND.n1403 19.3944
R20445 GND.n9150 GND.n1403 19.3944
R20446 GND.n9150 GND.n1399 19.3944
R20447 GND.n9156 GND.n1399 19.3944
R20448 GND.n9156 GND.n1397 19.3944
R20449 GND.n9160 GND.n1397 19.3944
R20450 GND.n9160 GND.n1393 19.3944
R20451 GND.n9166 GND.n1393 19.3944
R20452 GND.n9166 GND.n1391 19.3944
R20453 GND.n9170 GND.n1391 19.3944
R20454 GND.n9170 GND.n1387 19.3944
R20455 GND.n9176 GND.n1387 19.3944
R20456 GND.n9176 GND.n1385 19.3944
R20457 GND.n9180 GND.n1385 19.3944
R20458 GND.n9180 GND.n1381 19.3944
R20459 GND.n9186 GND.n1381 19.3944
R20460 GND.n9186 GND.n1379 19.3944
R20461 GND.n9190 GND.n1379 19.3944
R20462 GND.n9190 GND.n1375 19.3944
R20463 GND.n9196 GND.n1375 19.3944
R20464 GND.n9196 GND.n1373 19.3944
R20465 GND.n9200 GND.n1373 19.3944
R20466 GND.n9200 GND.n1369 19.3944
R20467 GND.n9206 GND.n1369 19.3944
R20468 GND.n9206 GND.n1367 19.3944
R20469 GND.n9210 GND.n1367 19.3944
R20470 GND.n9210 GND.n1363 19.3944
R20471 GND.n9216 GND.n1363 19.3944
R20472 GND.n9216 GND.n1361 19.3944
R20473 GND.n9220 GND.n1361 19.3944
R20474 GND.n9220 GND.n1357 19.3944
R20475 GND.n9226 GND.n1357 19.3944
R20476 GND.n9226 GND.n1355 19.3944
R20477 GND.n9230 GND.n1355 19.3944
R20478 GND.n9230 GND.n1351 19.3944
R20479 GND.n9236 GND.n1351 19.3944
R20480 GND.n9236 GND.n1349 19.3944
R20481 GND.n9240 GND.n1349 19.3944
R20482 GND.n9240 GND.n1345 19.3944
R20483 GND.n9246 GND.n1345 19.3944
R20484 GND.n9246 GND.n1343 19.3944
R20485 GND.n9250 GND.n1343 19.3944
R20486 GND.n9250 GND.n1339 19.3944
R20487 GND.n9256 GND.n1339 19.3944
R20488 GND.n9256 GND.n1337 19.3944
R20489 GND.n9260 GND.n1337 19.3944
R20490 GND.n9260 GND.n1333 19.3944
R20491 GND.n9266 GND.n1333 19.3944
R20492 GND.n9266 GND.n1331 19.3944
R20493 GND.n9270 GND.n1331 19.3944
R20494 GND.n9270 GND.n1327 19.3944
R20495 GND.n9276 GND.n1327 19.3944
R20496 GND.n9276 GND.n1325 19.3944
R20497 GND.n9280 GND.n1325 19.3944
R20498 GND.n9280 GND.n1321 19.3944
R20499 GND.n9286 GND.n1321 19.3944
R20500 GND.n9286 GND.n1319 19.3944
R20501 GND.n9290 GND.n1319 19.3944
R20502 GND.n9290 GND.n1315 19.3944
R20503 GND.n9296 GND.n1315 19.3944
R20504 GND.n9296 GND.n1313 19.3944
R20505 GND.n9300 GND.n1313 19.3944
R20506 GND.n9300 GND.n1309 19.3944
R20507 GND.n9306 GND.n1309 19.3944
R20508 GND.n9306 GND.n1307 19.3944
R20509 GND.n9310 GND.n1307 19.3944
R20510 GND.n9310 GND.n1303 19.3944
R20511 GND.n9316 GND.n1303 19.3944
R20512 GND.n9316 GND.n1301 19.3944
R20513 GND.n9320 GND.n1301 19.3944
R20514 GND.n9320 GND.n1297 19.3944
R20515 GND.n9326 GND.n1297 19.3944
R20516 GND.n9326 GND.n1295 19.3944
R20517 GND.n9330 GND.n1295 19.3944
R20518 GND.n9330 GND.n1291 19.3944
R20519 GND.n9336 GND.n1291 19.3944
R20520 GND.n9336 GND.n1289 19.3944
R20521 GND.n9340 GND.n1289 19.3944
R20522 GND.n9340 GND.n1285 19.3944
R20523 GND.n9346 GND.n1285 19.3944
R20524 GND.n9346 GND.n1283 19.3944
R20525 GND.n9350 GND.n1283 19.3944
R20526 GND.n9350 GND.n1279 19.3944
R20527 GND.n9356 GND.n1279 19.3944
R20528 GND.n9356 GND.n1277 19.3944
R20529 GND.n9360 GND.n1277 19.3944
R20530 GND.n9360 GND.n1273 19.3944
R20531 GND.n9366 GND.n1273 19.3944
R20532 GND.n9366 GND.n1271 19.3944
R20533 GND.n9370 GND.n1271 19.3944
R20534 GND.n9370 GND.n1267 19.3944
R20535 GND.n9376 GND.n1267 19.3944
R20536 GND.n9376 GND.n1265 19.3944
R20537 GND.n9380 GND.n1265 19.3944
R20538 GND.n9380 GND.n1261 19.3944
R20539 GND.n9386 GND.n1261 19.3944
R20540 GND.n9386 GND.n1259 19.3944
R20541 GND.n9390 GND.n1259 19.3944
R20542 GND.n9390 GND.n1255 19.3944
R20543 GND.n9396 GND.n1255 19.3944
R20544 GND.n9396 GND.n1253 19.3944
R20545 GND.n9400 GND.n1253 19.3944
R20546 GND.n9400 GND.n1249 19.3944
R20547 GND.n9406 GND.n1249 19.3944
R20548 GND.n9406 GND.n1247 19.3944
R20549 GND.n9410 GND.n1247 19.3944
R20550 GND.n9410 GND.n1243 19.3944
R20551 GND.n9416 GND.n1243 19.3944
R20552 GND.n9416 GND.n1241 19.3944
R20553 GND.n9420 GND.n1241 19.3944
R20554 GND.n9420 GND.n1237 19.3944
R20555 GND.n9426 GND.n1237 19.3944
R20556 GND.n9426 GND.n1235 19.3944
R20557 GND.n9430 GND.n1235 19.3944
R20558 GND.n9430 GND.n1231 19.3944
R20559 GND.n9436 GND.n1231 19.3944
R20560 GND.n9436 GND.n1229 19.3944
R20561 GND.n9440 GND.n1229 19.3944
R20562 GND.n9440 GND.n1225 19.3944
R20563 GND.n9446 GND.n1225 19.3944
R20564 GND.n9446 GND.n1223 19.3944
R20565 GND.n9450 GND.n1223 19.3944
R20566 GND.n9450 GND.n1219 19.3944
R20567 GND.n9456 GND.n1219 19.3944
R20568 GND.n9456 GND.n1217 19.3944
R20569 GND.n9460 GND.n1217 19.3944
R20570 GND.n9460 GND.n1213 19.3944
R20571 GND.n9466 GND.n1213 19.3944
R20572 GND.n9466 GND.n1211 19.3944
R20573 GND.n9470 GND.n1211 19.3944
R20574 GND.n9470 GND.n1207 19.3944
R20575 GND.n9476 GND.n1207 19.3944
R20576 GND.n9476 GND.n1205 19.3944
R20577 GND.n9480 GND.n1205 19.3944
R20578 GND.n9480 GND.n1201 19.3944
R20579 GND.n9486 GND.n1201 19.3944
R20580 GND.n9486 GND.n1199 19.3944
R20581 GND.n9490 GND.n1199 19.3944
R20582 GND.n9490 GND.n1195 19.3944
R20583 GND.n9496 GND.n1195 19.3944
R20584 GND.n9496 GND.n1193 19.3944
R20585 GND.n9500 GND.n1193 19.3944
R20586 GND.n9500 GND.n1189 19.3944
R20587 GND.n9506 GND.n1189 19.3944
R20588 GND.n9506 GND.n1187 19.3944
R20589 GND.n9510 GND.n1187 19.3944
R20590 GND.n9510 GND.n1183 19.3944
R20591 GND.n9516 GND.n1183 19.3944
R20592 GND.n9516 GND.n1181 19.3944
R20593 GND.n9520 GND.n1181 19.3944
R20594 GND.n9520 GND.n1177 19.3944
R20595 GND.n9526 GND.n1177 19.3944
R20596 GND.n9526 GND.n1175 19.3944
R20597 GND.n9530 GND.n1175 19.3944
R20598 GND.n9530 GND.n1171 19.3944
R20599 GND.n9536 GND.n1171 19.3944
R20600 GND.n9536 GND.n1169 19.3944
R20601 GND.n9540 GND.n1169 19.3944
R20602 GND.n9540 GND.n1165 19.3944
R20603 GND.n9546 GND.n1165 19.3944
R20604 GND.n9546 GND.n1163 19.3944
R20605 GND.n9550 GND.n1163 19.3944
R20606 GND.n9550 GND.n1159 19.3944
R20607 GND.n9556 GND.n1159 19.3944
R20608 GND.n9556 GND.n1157 19.3944
R20609 GND.n9560 GND.n1157 19.3944
R20610 GND.n9560 GND.n1153 19.3944
R20611 GND.n9566 GND.n1153 19.3944
R20612 GND.n9566 GND.n1151 19.3944
R20613 GND.n9570 GND.n1151 19.3944
R20614 GND.n9570 GND.n1147 19.3944
R20615 GND.n9576 GND.n1147 19.3944
R20616 GND.n9576 GND.n1145 19.3944
R20617 GND.n9580 GND.n1145 19.3944
R20618 GND.n9580 GND.n1141 19.3944
R20619 GND.n9586 GND.n1141 19.3944
R20620 GND.n9586 GND.n1139 19.3944
R20621 GND.n9590 GND.n1139 19.3944
R20622 GND.n9590 GND.n1135 19.3944
R20623 GND.n9596 GND.n1135 19.3944
R20624 GND.n9596 GND.n1133 19.3944
R20625 GND.n9600 GND.n1133 19.3944
R20626 GND.n9600 GND.n1129 19.3944
R20627 GND.n9606 GND.n1129 19.3944
R20628 GND.n9606 GND.n1127 19.3944
R20629 GND.n9610 GND.n1127 19.3944
R20630 GND.n9610 GND.n1123 19.3944
R20631 GND.n9616 GND.n1123 19.3944
R20632 GND.n9616 GND.n1121 19.3944
R20633 GND.n9620 GND.n1121 19.3944
R20634 GND.n9620 GND.n1117 19.3944
R20635 GND.n9626 GND.n1117 19.3944
R20636 GND.n9626 GND.n1115 19.3944
R20637 GND.n9630 GND.n1115 19.3944
R20638 GND.n9630 GND.n1111 19.3944
R20639 GND.n9636 GND.n1111 19.3944
R20640 GND.n9636 GND.n1109 19.3944
R20641 GND.n9640 GND.n1109 19.3944
R20642 GND.n9640 GND.n1105 19.3944
R20643 GND.n9646 GND.n1105 19.3944
R20644 GND.n9646 GND.n1103 19.3944
R20645 GND.n9650 GND.n1103 19.3944
R20646 GND.n9650 GND.n1099 19.3944
R20647 GND.n9656 GND.n1099 19.3944
R20648 GND.n9656 GND.n1097 19.3944
R20649 GND.n9660 GND.n1097 19.3944
R20650 GND.n9660 GND.n1093 19.3944
R20651 GND.n9666 GND.n1093 19.3944
R20652 GND.n9666 GND.n1091 19.3944
R20653 GND.n9670 GND.n1091 19.3944
R20654 GND.n9670 GND.n1087 19.3944
R20655 GND.n9676 GND.n1087 19.3944
R20656 GND.n9676 GND.n1085 19.3944
R20657 GND.n9680 GND.n1085 19.3944
R20658 GND.n9680 GND.n1081 19.3944
R20659 GND.n9686 GND.n1081 19.3944
R20660 GND.n9686 GND.n1079 19.3944
R20661 GND.n9690 GND.n1079 19.3944
R20662 GND.n9690 GND.n1075 19.3944
R20663 GND.n9696 GND.n1075 19.3944
R20664 GND.n9696 GND.n1073 19.3944
R20665 GND.n9700 GND.n1073 19.3944
R20666 GND.n9700 GND.n1069 19.3944
R20667 GND.n9706 GND.n1069 19.3944
R20668 GND.n9706 GND.n1067 19.3944
R20669 GND.n9710 GND.n1067 19.3944
R20670 GND.n9710 GND.n1063 19.3944
R20671 GND.n9716 GND.n1063 19.3944
R20672 GND.n9716 GND.n1061 19.3944
R20673 GND.n9720 GND.n1061 19.3944
R20674 GND.n9720 GND.n1057 19.3944
R20675 GND.n9726 GND.n1057 19.3944
R20676 GND.n9726 GND.n1055 19.3944
R20677 GND.n9730 GND.n1055 19.3944
R20678 GND.n9730 GND.n1051 19.3944
R20679 GND.n9736 GND.n1051 19.3944
R20680 GND.n9736 GND.n1049 19.3944
R20681 GND.n9740 GND.n1049 19.3944
R20682 GND.n9740 GND.n1045 19.3944
R20683 GND.n9746 GND.n1045 19.3944
R20684 GND.n9746 GND.n1043 19.3944
R20685 GND.n9750 GND.n1043 19.3944
R20686 GND.n9750 GND.n1039 19.3944
R20687 GND.n9756 GND.n1039 19.3944
R20688 GND.n9756 GND.n1037 19.3944
R20689 GND.n9760 GND.n1037 19.3944
R20690 GND.n9760 GND.n1033 19.3944
R20691 GND.n9766 GND.n1033 19.3944
R20692 GND.n9766 GND.n1031 19.3944
R20693 GND.n9770 GND.n1031 19.3944
R20694 GND.n9770 GND.n1027 19.3944
R20695 GND.n9776 GND.n1027 19.3944
R20696 GND.n9776 GND.n1025 19.3944
R20697 GND.n9780 GND.n1025 19.3944
R20698 GND.n9780 GND.n1021 19.3944
R20699 GND.n9786 GND.n1021 19.3944
R20700 GND.n9786 GND.n1019 19.3944
R20701 GND.n9790 GND.n1019 19.3944
R20702 GND.n9790 GND.n1015 19.3944
R20703 GND.n9796 GND.n1015 19.3944
R20704 GND.n9796 GND.n1013 19.3944
R20705 GND.n9800 GND.n1013 19.3944
R20706 GND.n9800 GND.n1009 19.3944
R20707 GND.n9806 GND.n1009 19.3944
R20708 GND.n9806 GND.n1007 19.3944
R20709 GND.n9810 GND.n1007 19.3944
R20710 GND.n9810 GND.n1003 19.3944
R20711 GND.n9816 GND.n1003 19.3944
R20712 GND.n9816 GND.n1001 19.3944
R20713 GND.n9820 GND.n1001 19.3944
R20714 GND.n9820 GND.n997 19.3944
R20715 GND.n9826 GND.n997 19.3944
R20716 GND.n9826 GND.n995 19.3944
R20717 GND.n9830 GND.n995 19.3944
R20718 GND.n9830 GND.n991 19.3944
R20719 GND.n9836 GND.n991 19.3944
R20720 GND.n9836 GND.n989 19.3944
R20721 GND.n9840 GND.n989 19.3944
R20722 GND.n9840 GND.n985 19.3944
R20723 GND.n9846 GND.n985 19.3944
R20724 GND.n9846 GND.n983 19.3944
R20725 GND.n9850 GND.n983 19.3944
R20726 GND.n9850 GND.n979 19.3944
R20727 GND.n9856 GND.n979 19.3944
R20728 GND.n9856 GND.n977 19.3944
R20729 GND.n9860 GND.n977 19.3944
R20730 GND.n9860 GND.n973 19.3944
R20731 GND.n9866 GND.n973 19.3944
R20732 GND.n9866 GND.n971 19.3944
R20733 GND.n9870 GND.n971 19.3944
R20734 GND.n9870 GND.n967 19.3944
R20735 GND.n9876 GND.n967 19.3944
R20736 GND.n9876 GND.n965 19.3944
R20737 GND.n9880 GND.n965 19.3944
R20738 GND.n9880 GND.n961 19.3944
R20739 GND.n9886 GND.n961 19.3944
R20740 GND.n9886 GND.n959 19.3944
R20741 GND.n9890 GND.n959 19.3944
R20742 GND.n9890 GND.n955 19.3944
R20743 GND.n9896 GND.n955 19.3944
R20744 GND.n9896 GND.n953 19.3944
R20745 GND.n9900 GND.n953 19.3944
R20746 GND.n9900 GND.n949 19.3944
R20747 GND.n9906 GND.n949 19.3944
R20748 GND.n9906 GND.n947 19.3944
R20749 GND.n9910 GND.n947 19.3944
R20750 GND.n9910 GND.n943 19.3944
R20751 GND.n9916 GND.n943 19.3944
R20752 GND.n9916 GND.n941 19.3944
R20753 GND.n9920 GND.n941 19.3944
R20754 GND.n9920 GND.n937 19.3944
R20755 GND.n9926 GND.n937 19.3944
R20756 GND.n9926 GND.n935 19.3944
R20757 GND.n9930 GND.n935 19.3944
R20758 GND.n9930 GND.n931 19.3944
R20759 GND.n9936 GND.n931 19.3944
R20760 GND.n9936 GND.n929 19.3944
R20761 GND.n9940 GND.n929 19.3944
R20762 GND.n9940 GND.n925 19.3944
R20763 GND.n9946 GND.n925 19.3944
R20764 GND.n9946 GND.n923 19.3944
R20765 GND.n9950 GND.n923 19.3944
R20766 GND.n9950 GND.n919 19.3944
R20767 GND.n9956 GND.n919 19.3944
R20768 GND.n9956 GND.n917 19.3944
R20769 GND.n9960 GND.n917 19.3944
R20770 GND.n9960 GND.n913 19.3944
R20771 GND.n9966 GND.n913 19.3944
R20772 GND.n9966 GND.n911 19.3944
R20773 GND.n9970 GND.n911 19.3944
R20774 GND.n9970 GND.n907 19.3944
R20775 GND.n9976 GND.n907 19.3944
R20776 GND.n9976 GND.n905 19.3944
R20777 GND.n9980 GND.n905 19.3944
R20778 GND.n9980 GND.n901 19.3944
R20779 GND.n9986 GND.n901 19.3944
R20780 GND.n9986 GND.n899 19.3944
R20781 GND.n9990 GND.n899 19.3944
R20782 GND.n9990 GND.n895 19.3944
R20783 GND.n9996 GND.n895 19.3944
R20784 GND.n9996 GND.n893 19.3944
R20785 GND.n10000 GND.n893 19.3944
R20786 GND.n10000 GND.n889 19.3944
R20787 GND.n10006 GND.n889 19.3944
R20788 GND.n10006 GND.n887 19.3944
R20789 GND.n10010 GND.n887 19.3944
R20790 GND.n10010 GND.n883 19.3944
R20791 GND.n10016 GND.n883 19.3944
R20792 GND.n10016 GND.n881 19.3944
R20793 GND.n10020 GND.n881 19.3944
R20794 GND.n10020 GND.n877 19.3944
R20795 GND.n10026 GND.n877 19.3944
R20796 GND.n10026 GND.n875 19.3944
R20797 GND.n10030 GND.n875 19.3944
R20798 GND.n10030 GND.n871 19.3944
R20799 GND.n10036 GND.n871 19.3944
R20800 GND.n10036 GND.n869 19.3944
R20801 GND.n10040 GND.n869 19.3944
R20802 GND.n10040 GND.n865 19.3944
R20803 GND.n10046 GND.n865 19.3944
R20804 GND.n10046 GND.n863 19.3944
R20805 GND.n10050 GND.n863 19.3944
R20806 GND.n10050 GND.n859 19.3944
R20807 GND.n10056 GND.n859 19.3944
R20808 GND.n10056 GND.n857 19.3944
R20809 GND.n10060 GND.n857 19.3944
R20810 GND.n10060 GND.n853 19.3944
R20811 GND.n10066 GND.n853 19.3944
R20812 GND.n10066 GND.n851 19.3944
R20813 GND.n10070 GND.n851 19.3944
R20814 GND.n10070 GND.n847 19.3944
R20815 GND.n10076 GND.n847 19.3944
R20816 GND.n10076 GND.n845 19.3944
R20817 GND.n10080 GND.n845 19.3944
R20818 GND.n10080 GND.n841 19.3944
R20819 GND.n10086 GND.n841 19.3944
R20820 GND.n10086 GND.n839 19.3944
R20821 GND.n10090 GND.n839 19.3944
R20822 GND.n10090 GND.n835 19.3944
R20823 GND.n10096 GND.n835 19.3944
R20824 GND.n10096 GND.n833 19.3944
R20825 GND.n10100 GND.n833 19.3944
R20826 GND.n10100 GND.n829 19.3944
R20827 GND.n10106 GND.n829 19.3944
R20828 GND.n10106 GND.n827 19.3944
R20829 GND.n10110 GND.n827 19.3944
R20830 GND.n10110 GND.n823 19.3944
R20831 GND.n10116 GND.n823 19.3944
R20832 GND.n10116 GND.n821 19.3944
R20833 GND.n10120 GND.n821 19.3944
R20834 GND.n10120 GND.n817 19.3944
R20835 GND.n10126 GND.n817 19.3944
R20836 GND.n10126 GND.n815 19.3944
R20837 GND.n10130 GND.n815 19.3944
R20838 GND.n10130 GND.n811 19.3944
R20839 GND.n10136 GND.n811 19.3944
R20840 GND.n10136 GND.n809 19.3944
R20841 GND.n10140 GND.n809 19.3944
R20842 GND.n10140 GND.n805 19.3944
R20843 GND.n10146 GND.n805 19.3944
R20844 GND.n10146 GND.n803 19.3944
R20845 GND.n10150 GND.n803 19.3944
R20846 GND.n10150 GND.n799 19.3944
R20847 GND.n10156 GND.n799 19.3944
R20848 GND.n10156 GND.n797 19.3944
R20849 GND.n10160 GND.n797 19.3944
R20850 GND.n10160 GND.n793 19.3944
R20851 GND.n10166 GND.n793 19.3944
R20852 GND.n10166 GND.n791 19.3944
R20853 GND.n10170 GND.n791 19.3944
R20854 GND.n10170 GND.n787 19.3944
R20855 GND.n10176 GND.n787 19.3944
R20856 GND.n10176 GND.n785 19.3944
R20857 GND.n10180 GND.n785 19.3944
R20858 GND.n10180 GND.n781 19.3944
R20859 GND.n10186 GND.n781 19.3944
R20860 GND.n10186 GND.n779 19.3944
R20861 GND.n10190 GND.n779 19.3944
R20862 GND.n10190 GND.n775 19.3944
R20863 GND.n10196 GND.n775 19.3944
R20864 GND.n10196 GND.n773 19.3944
R20865 GND.n10200 GND.n773 19.3944
R20866 GND.n10200 GND.n769 19.3944
R20867 GND.n10206 GND.n769 19.3944
R20868 GND.n10206 GND.n767 19.3944
R20869 GND.n10210 GND.n767 19.3944
R20870 GND.n10210 GND.n763 19.3944
R20871 GND.n10216 GND.n763 19.3944
R20872 GND.n10216 GND.n761 19.3944
R20873 GND.n10220 GND.n761 19.3944
R20874 GND.n10220 GND.n757 19.3944
R20875 GND.n10226 GND.n757 19.3944
R20876 GND.n10226 GND.n755 19.3944
R20877 GND.n10230 GND.n755 19.3944
R20878 GND.n10230 GND.n751 19.3944
R20879 GND.n10236 GND.n751 19.3944
R20880 GND.n10236 GND.n749 19.3944
R20881 GND.n10240 GND.n749 19.3944
R20882 GND.n10240 GND.n745 19.3944
R20883 GND.n10246 GND.n745 19.3944
R20884 GND.n10246 GND.n743 19.3944
R20885 GND.n10250 GND.n743 19.3944
R20886 GND.n10250 GND.n739 19.3944
R20887 GND.n10256 GND.n739 19.3944
R20888 GND.n10256 GND.n737 19.3944
R20889 GND.n10260 GND.n737 19.3944
R20890 GND.n10260 GND.n733 19.3944
R20891 GND.n10266 GND.n733 19.3944
R20892 GND.n10266 GND.n731 19.3944
R20893 GND.n10270 GND.n731 19.3944
R20894 GND.n10270 GND.n727 19.3944
R20895 GND.n10276 GND.n727 19.3944
R20896 GND.n10276 GND.n725 19.3944
R20897 GND.n10280 GND.n725 19.3944
R20898 GND.n10280 GND.n721 19.3944
R20899 GND.n10286 GND.n721 19.3944
R20900 GND.n10286 GND.n719 19.3944
R20901 GND.n10290 GND.n719 19.3944
R20902 GND.n10290 GND.n715 19.3944
R20903 GND.n10296 GND.n715 19.3944
R20904 GND.n10296 GND.n713 19.3944
R20905 GND.n10300 GND.n713 19.3944
R20906 GND.n10300 GND.n709 19.3944
R20907 GND.n10306 GND.n709 19.3944
R20908 GND.n10306 GND.n707 19.3944
R20909 GND.n10310 GND.n707 19.3944
R20910 GND.n10310 GND.n703 19.3944
R20911 GND.n10316 GND.n703 19.3944
R20912 GND.n10316 GND.n701 19.3944
R20913 GND.n10320 GND.n701 19.3944
R20914 GND.n10320 GND.n697 19.3944
R20915 GND.n10326 GND.n697 19.3944
R20916 GND.n10326 GND.n695 19.3944
R20917 GND.n10330 GND.n695 19.3944
R20918 GND.n10330 GND.n691 19.3944
R20919 GND.n10336 GND.n691 19.3944
R20920 GND.n10336 GND.n689 19.3944
R20921 GND.n10340 GND.n689 19.3944
R20922 GND.n10340 GND.n685 19.3944
R20923 GND.n10346 GND.n685 19.3944
R20924 GND.n10346 GND.n683 19.3944
R20925 GND.n10350 GND.n683 19.3944
R20926 GND.n10350 GND.n679 19.3944
R20927 GND.n10356 GND.n679 19.3944
R20928 GND.n10356 GND.n677 19.3944
R20929 GND.n10360 GND.n677 19.3944
R20930 GND.n10360 GND.n673 19.3944
R20931 GND.n10366 GND.n673 19.3944
R20932 GND.n10366 GND.n671 19.3944
R20933 GND.n10370 GND.n671 19.3944
R20934 GND.n10370 GND.n667 19.3944
R20935 GND.n10376 GND.n667 19.3944
R20936 GND.n10376 GND.n665 19.3944
R20937 GND.n10381 GND.n665 19.3944
R20938 GND.n10381 GND.n10380 19.3944
R20939 GND.n7644 GND.n7643 19.3944
R20940 GND.n7643 GND.n7642 19.3944
R20941 GND.n7642 GND.n7641 19.3944
R20942 GND.n7641 GND.n7639 19.3944
R20943 GND.n7639 GND.n7636 19.3944
R20944 GND.n7636 GND.n7635 19.3944
R20945 GND.n7635 GND.n7632 19.3944
R20946 GND.n7632 GND.n7631 19.3944
R20947 GND.n7631 GND.n7628 19.3944
R20948 GND.n7628 GND.n7627 19.3944
R20949 GND.n7627 GND.n7624 19.3944
R20950 GND.n7622 GND.n7620 19.3944
R20951 GND.n7620 GND.n7617 19.3944
R20952 GND.n7617 GND.n7616 19.3944
R20953 GND.n7616 GND.n7613 19.3944
R20954 GND.n7613 GND.n7612 19.3944
R20955 GND.n7612 GND.n7609 19.3944
R20956 GND.n7609 GND.n7608 19.3944
R20957 GND.n7608 GND.n7605 19.3944
R20958 GND.n7605 GND.n7604 19.3944
R20959 GND.n7604 GND.n7601 19.3944
R20960 GND.n7601 GND.n7600 19.3944
R20961 GND.n7596 GND.n7594 19.3944
R20962 GND.n7594 GND.n7591 19.3944
R20963 GND.n7591 GND.n7590 19.3944
R20964 GND.n7590 GND.n7587 19.3944
R20965 GND.n7587 GND.n7586 19.3944
R20966 GND.n7586 GND.n7583 19.3944
R20967 GND.n7583 GND.n7582 19.3944
R20968 GND.n7582 GND.n7579 19.3944
R20969 GND.n7579 GND.n7578 19.3944
R20970 GND.n7578 GND.n7575 19.3944
R20971 GND.n7575 GND.n7574 19.3944
R20972 GND.n7574 GND.n7571 19.3944
R20973 GND.n7571 GND.n7570 19.3944
R20974 GND.n7567 GND.n7566 19.3944
R20975 GND.n7566 GND.n7563 19.3944
R20976 GND.n7563 GND.n7562 19.3944
R20977 GND.n7562 GND.n7559 19.3944
R20978 GND.n7559 GND.n7558 19.3944
R20979 GND.n7558 GND.n7555 19.3944
R20980 GND.n7555 GND.n7554 19.3944
R20981 GND.n7554 GND.n7551 19.3944
R20982 GND.n7551 GND.n7550 19.3944
R20983 GND.n7550 GND.n7547 19.3944
R20984 GND.n7547 GND.n7546 19.3944
R20985 GND.n7546 GND.n7543 19.3944
R20986 GND.n7543 GND.n7542 19.3944
R20987 GND.n7534 GND.n5876 19.3944
R20988 GND.n6743 GND.n5876 19.3944
R20989 GND.n6743 GND.n6736 19.3944
R20990 GND.n6755 GND.n6736 19.3944
R20991 GND.n6756 GND.n6755 19.3944
R20992 GND.n6758 GND.n6756 19.3944
R20993 GND.n6758 GND.n6530 19.3944
R20994 GND.n6770 GND.n6530 19.3944
R20995 GND.n6771 GND.n6770 19.3944
R20996 GND.n6773 GND.n6771 19.3944
R20997 GND.n6773 GND.n6526 19.3944
R20998 GND.n6785 GND.n6526 19.3944
R20999 GND.n6786 GND.n6785 19.3944
R21000 GND.n6788 GND.n6786 19.3944
R21001 GND.n6788 GND.n6522 19.3944
R21002 GND.n6800 GND.n6522 19.3944
R21003 GND.n6801 GND.n6800 19.3944
R21004 GND.n6803 GND.n6801 19.3944
R21005 GND.n6803 GND.n6518 19.3944
R21006 GND.n6815 GND.n6518 19.3944
R21007 GND.n6816 GND.n6815 19.3944
R21008 GND.n6818 GND.n6816 19.3944
R21009 GND.n6818 GND.n6513 19.3944
R21010 GND.n6830 GND.n6513 19.3944
R21011 GND.n6831 GND.n6830 19.3944
R21012 GND.n6833 GND.n6831 19.3944
R21013 GND.n6833 GND.n6509 19.3944
R21014 GND.n6845 GND.n6509 19.3944
R21015 GND.n6846 GND.n6845 19.3944
R21016 GND.n6848 GND.n6846 19.3944
R21017 GND.n6848 GND.n6505 19.3944
R21018 GND.n6860 GND.n6505 19.3944
R21019 GND.n6861 GND.n6860 19.3944
R21020 GND.n6863 GND.n6861 19.3944
R21021 GND.n6863 GND.n6501 19.3944
R21022 GND.n6875 GND.n6501 19.3944
R21023 GND.n6876 GND.n6875 19.3944
R21024 GND.n6878 GND.n6876 19.3944
R21025 GND.n6878 GND.n6497 19.3944
R21026 GND.n6890 GND.n6497 19.3944
R21027 GND.n6891 GND.n6890 19.3944
R21028 GND.n6893 GND.n6891 19.3944
R21029 GND.n6893 GND.n6493 19.3944
R21030 GND.n6905 GND.n6493 19.3944
R21031 GND.n6906 GND.n6905 19.3944
R21032 GND.n6908 GND.n6906 19.3944
R21033 GND.n6908 GND.n6489 19.3944
R21034 GND.n6920 GND.n6489 19.3944
R21035 GND.n6921 GND.n6920 19.3944
R21036 GND.n6923 GND.n6921 19.3944
R21037 GND.n6923 GND.n6484 19.3944
R21038 GND.n6935 GND.n6484 19.3944
R21039 GND.n6936 GND.n6935 19.3944
R21040 GND.n6938 GND.n6936 19.3944
R21041 GND.n6938 GND.n6480 19.3944
R21042 GND.n6950 GND.n6480 19.3944
R21043 GND.n6951 GND.n6950 19.3944
R21044 GND.n6953 GND.n6951 19.3944
R21045 GND.n6953 GND.n6476 19.3944
R21046 GND.n6965 GND.n6476 19.3944
R21047 GND.n6966 GND.n6965 19.3944
R21048 GND.n6968 GND.n6966 19.3944
R21049 GND.n6968 GND.n6472 19.3944
R21050 GND.n6987 GND.n6472 19.3944
R21051 GND.n6988 GND.n6987 19.3944
R21052 GND.n6989 GND.n6988 19.3944
R21053 GND.n6992 GND.n6989 19.3944
R21054 GND.n6992 GND.n6467 19.3944
R21055 GND.n7000 GND.n6467 19.3944
R21056 GND.n7001 GND.n7000 19.3944
R21057 GND.n7001 GND.n6463 19.3944
R21058 GND.n7010 GND.n6463 19.3944
R21059 GND.n7011 GND.n7010 19.3944
R21060 GND.n7012 GND.n7011 19.3944
R21061 GND.n7013 GND.n7012 19.3944
R21062 GND.n7015 GND.n7013 19.3944
R21063 GND.n7015 GND.n6460 19.3944
R21064 GND.n7027 GND.n6460 19.3944
R21065 GND.n7028 GND.n7027 19.3944
R21066 GND.n7030 GND.n7028 19.3944
R21067 GND.n7030 GND.n6456 19.3944
R21068 GND.n7042 GND.n6456 19.3944
R21069 GND.n7043 GND.n7042 19.3944
R21070 GND.n7045 GND.n7043 19.3944
R21071 GND.n7045 GND.n6452 19.3944
R21072 GND.n7057 GND.n6452 19.3944
R21073 GND.n7058 GND.n7057 19.3944
R21074 GND.n7060 GND.n7058 19.3944
R21075 GND.n7060 GND.n6448 19.3944
R21076 GND.n7072 GND.n6448 19.3944
R21077 GND.n7073 GND.n7072 19.3944
R21078 GND.n7075 GND.n7073 19.3944
R21079 GND.n7075 GND.n6444 19.3944
R21080 GND.n7087 GND.n6444 19.3944
R21081 GND.n7088 GND.n7087 19.3944
R21082 GND.n7090 GND.n7088 19.3944
R21083 GND.n7090 GND.n6440 19.3944
R21084 GND.n7103 GND.n6440 19.3944
R21085 GND.n7104 GND.n7103 19.3944
R21086 GND.n7106 GND.n7104 19.3944
R21087 GND.n7107 GND.n7106 19.3944
R21088 GND.n7260 GND.n7107 19.3944
R21089 GND.n7260 GND.n7259 19.3944
R21090 GND.n7259 GND.n7258 19.3944
R21091 GND.n7258 GND.n7109 19.3944
R21092 GND.n7248 GND.n7109 19.3944
R21093 GND.n7248 GND.n7247 19.3944
R21094 GND.n7247 GND.n7246 19.3944
R21095 GND.n7246 GND.n7116 19.3944
R21096 GND.n7236 GND.n7116 19.3944
R21097 GND.n7236 GND.n7235 19.3944
R21098 GND.n7235 GND.n7234 19.3944
R21099 GND.n7234 GND.n7123 19.3944
R21100 GND.n7224 GND.n7123 19.3944
R21101 GND.n7224 GND.n7223 19.3944
R21102 GND.n7223 GND.n7222 19.3944
R21103 GND.n7222 GND.n7130 19.3944
R21104 GND.n7212 GND.n7130 19.3944
R21105 GND.n7212 GND.n7211 19.3944
R21106 GND.n7211 GND.n7210 19.3944
R21107 GND.n7210 GND.n7137 19.3944
R21108 GND.n7200 GND.n7137 19.3944
R21109 GND.n7200 GND.n7199 19.3944
R21110 GND.n7199 GND.n7198 19.3944
R21111 GND.n7198 GND.n7144 19.3944
R21112 GND.n7188 GND.n7144 19.3944
R21113 GND.n7188 GND.n7187 19.3944
R21114 GND.n7187 GND.n7186 19.3944
R21115 GND.n7186 GND.n7151 19.3944
R21116 GND.n7176 GND.n7151 19.3944
R21117 GND.n7176 GND.n7175 19.3944
R21118 GND.n7175 GND.n7174 19.3944
R21119 GND.n7174 GND.n7158 19.3944
R21120 GND.n7164 GND.n7158 19.3944
R21121 GND.n7164 GND.n452 19.3944
R21122 GND.n10907 GND.n452 19.3944
R21123 GND.n10908 GND.n10907 19.3944
R21124 GND.n5918 GND.n5874 19.3944
R21125 GND.n5934 GND.n5918 19.3944
R21126 GND.n7521 GND.n5934 19.3944
R21127 GND.n7521 GND.n7520 19.3944
R21128 GND.n7520 GND.n7519 19.3944
R21129 GND.n7519 GND.n5938 19.3944
R21130 GND.n7509 GND.n5938 19.3944
R21131 GND.n7509 GND.n7508 19.3944
R21132 GND.n7508 GND.n7507 19.3944
R21133 GND.n7507 GND.n5958 19.3944
R21134 GND.n7497 GND.n5958 19.3944
R21135 GND.n7497 GND.n7496 19.3944
R21136 GND.n7496 GND.n7495 19.3944
R21137 GND.n7495 GND.n5979 19.3944
R21138 GND.n7485 GND.n5979 19.3944
R21139 GND.n7485 GND.n7484 19.3944
R21140 GND.n7484 GND.n7483 19.3944
R21141 GND.n7483 GND.n6000 19.3944
R21142 GND.n7473 GND.n6000 19.3944
R21143 GND.n7473 GND.n7472 19.3944
R21144 GND.n7472 GND.n7471 19.3944
R21145 GND.n7471 GND.n6021 19.3944
R21146 GND.n7461 GND.n6021 19.3944
R21147 GND.n7461 GND.n7460 19.3944
R21148 GND.n7460 GND.n7459 19.3944
R21149 GND.n7459 GND.n6041 19.3944
R21150 GND.n7449 GND.n6041 19.3944
R21151 GND.n7449 GND.n7448 19.3944
R21152 GND.n7448 GND.n7447 19.3944
R21153 GND.n7447 GND.n6062 19.3944
R21154 GND.n7437 GND.n6062 19.3944
R21155 GND.n7437 GND.n7436 19.3944
R21156 GND.n7436 GND.n7435 19.3944
R21157 GND.n7435 GND.n6083 19.3944
R21158 GND.n7425 GND.n6083 19.3944
R21159 GND.n7425 GND.n7424 19.3944
R21160 GND.n7424 GND.n7423 19.3944
R21161 GND.n7423 GND.n6104 19.3944
R21162 GND.n7413 GND.n6104 19.3944
R21163 GND.n7413 GND.n7412 19.3944
R21164 GND.n7412 GND.n7411 19.3944
R21165 GND.n7411 GND.n6125 19.3944
R21166 GND.n7401 GND.n6125 19.3944
R21167 GND.n7401 GND.n7400 19.3944
R21168 GND.n7400 GND.n7399 19.3944
R21169 GND.n7399 GND.n6146 19.3944
R21170 GND.n7389 GND.n6146 19.3944
R21171 GND.n7389 GND.n7388 19.3944
R21172 GND.n7388 GND.n7387 19.3944
R21173 GND.n7387 GND.n6167 19.3944
R21174 GND.n7377 GND.n6167 19.3944
R21175 GND.n7377 GND.n7376 19.3944
R21176 GND.n7376 GND.n7375 19.3944
R21177 GND.n7375 GND.n6187 19.3944
R21178 GND.n7365 GND.n6187 19.3944
R21179 GND.n7365 GND.n7364 19.3944
R21180 GND.n7364 GND.n7363 19.3944
R21181 GND.n7363 GND.n6208 19.3944
R21182 GND.n7353 GND.n6208 19.3944
R21183 GND.n7353 GND.n7352 19.3944
R21184 GND.n7352 GND.n7351 19.3944
R21185 GND.n7351 GND.n6229 19.3944
R21186 GND.n7341 GND.n6229 19.3944
R21187 GND.n7341 GND.n7340 19.3944
R21188 GND.n7340 GND.n7339 19.3944
R21189 GND.n7339 GND.n6249 19.3944
R21190 GND.n6469 GND.n6249 19.3944
R21191 GND.n6997 GND.n6469 19.3944
R21192 GND.n6998 GND.n6997 19.3944
R21193 GND.n6998 GND.n6465 19.3944
R21194 GND.n7007 GND.n6465 19.3944
R21195 GND.n7007 GND.n117 19.3944
R21196 GND.n11102 GND.n117 19.3944
R21197 GND.n11102 GND.n11101 19.3944
R21198 GND.n11101 GND.n11100 19.3944
R21199 GND.n11100 GND.n121 19.3944
R21200 GND.n11090 GND.n121 19.3944
R21201 GND.n11090 GND.n11089 19.3944
R21202 GND.n11089 GND.n11088 19.3944
R21203 GND.n11088 GND.n140 19.3944
R21204 GND.n11078 GND.n140 19.3944
R21205 GND.n11078 GND.n11077 19.3944
R21206 GND.n11077 GND.n11076 19.3944
R21207 GND.n11076 GND.n161 19.3944
R21208 GND.n11066 GND.n161 19.3944
R21209 GND.n11066 GND.n11065 19.3944
R21210 GND.n11065 GND.n11064 19.3944
R21211 GND.n11064 GND.n182 19.3944
R21212 GND.n11054 GND.n182 19.3944
R21213 GND.n11054 GND.n11053 19.3944
R21214 GND.n11053 GND.n11052 19.3944
R21215 GND.n11052 GND.n203 19.3944
R21216 GND.n11042 GND.n203 19.3944
R21217 GND.n11042 GND.n11041 19.3944
R21218 GND.n11041 GND.n11040 19.3944
R21219 GND.n11040 GND.n224 19.3944
R21220 GND.n11030 GND.n224 19.3944
R21221 GND.n11030 GND.n11029 19.3944
R21222 GND.n11029 GND.n11028 19.3944
R21223 GND.n11028 GND.n245 19.3944
R21224 GND.n11018 GND.n245 19.3944
R21225 GND.n11018 GND.n11017 19.3944
R21226 GND.n11017 GND.n11016 19.3944
R21227 GND.n11016 GND.n265 19.3944
R21228 GND.n11006 GND.n265 19.3944
R21229 GND.n11006 GND.n11005 19.3944
R21230 GND.n11005 GND.n11004 19.3944
R21231 GND.n11004 GND.n286 19.3944
R21232 GND.n10994 GND.n286 19.3944
R21233 GND.n10994 GND.n10993 19.3944
R21234 GND.n10993 GND.n10992 19.3944
R21235 GND.n10992 GND.n307 19.3944
R21236 GND.n10982 GND.n307 19.3944
R21237 GND.n10982 GND.n10981 19.3944
R21238 GND.n10981 GND.n10980 19.3944
R21239 GND.n10980 GND.n328 19.3944
R21240 GND.n10970 GND.n328 19.3944
R21241 GND.n10970 GND.n10969 19.3944
R21242 GND.n10969 GND.n10968 19.3944
R21243 GND.n10968 GND.n349 19.3944
R21244 GND.n10958 GND.n349 19.3944
R21245 GND.n10958 GND.n10957 19.3944
R21246 GND.n10957 GND.n10956 19.3944
R21247 GND.n10956 GND.n370 19.3944
R21248 GND.n10946 GND.n370 19.3944
R21249 GND.n10946 GND.n10945 19.3944
R21250 GND.n10945 GND.n10944 19.3944
R21251 GND.n10944 GND.n391 19.3944
R21252 GND.n10934 GND.n391 19.3944
R21253 GND.n10934 GND.n10933 19.3944
R21254 GND.n10933 GND.n10932 19.3944
R21255 GND.n10932 GND.n412 19.3944
R21256 GND.n10922 GND.n412 19.3944
R21257 GND.n10922 GND.n10921 19.3944
R21258 GND.n10921 GND.n10920 19.3944
R21259 GND.n10920 GND.n433 19.3944
R21260 GND.n10910 GND.n433 19.3944
R21261 GND.n10816 GND.n10815 19.3944
R21262 GND.n10815 GND.n10812 19.3944
R21263 GND.n10812 GND.n10811 19.3944
R21264 GND.n10811 GND.n10808 19.3944
R21265 GND.n10808 GND.n10807 19.3944
R21266 GND.n10807 GND.n10804 19.3944
R21267 GND.n10804 GND.n10803 19.3944
R21268 GND.n10803 GND.n10800 19.3944
R21269 GND.n10800 GND.n10799 19.3944
R21270 GND.n10799 GND.n10796 19.3944
R21271 GND.n10796 GND.n10795 19.3944
R21272 GND.n10795 GND.n10792 19.3944
R21273 GND.n10792 GND.n10791 19.3944
R21274 GND.n10844 GND.n10843 19.3944
R21275 GND.n10843 GND.n10840 19.3944
R21276 GND.n10840 GND.n10839 19.3944
R21277 GND.n10839 GND.n10836 19.3944
R21278 GND.n10836 GND.n10835 19.3944
R21279 GND.n10835 GND.n10832 19.3944
R21280 GND.n10832 GND.n10831 19.3944
R21281 GND.n10831 GND.n10828 19.3944
R21282 GND.n10828 GND.n10827 19.3944
R21283 GND.n10827 GND.n10824 19.3944
R21284 GND.n10824 GND.n10823 19.3944
R21285 GND.n10823 GND.n10820 19.3944
R21286 GND.n10820 GND.n10819 19.3944
R21287 GND.n10871 GND.n10731 19.3944
R21288 GND.n10871 GND.n10868 19.3944
R21289 GND.n10868 GND.n10867 19.3944
R21290 GND.n10867 GND.n10864 19.3944
R21291 GND.n10864 GND.n10863 19.3944
R21292 GND.n10863 GND.n10860 19.3944
R21293 GND.n10860 GND.n10859 19.3944
R21294 GND.n10859 GND.n10856 19.3944
R21295 GND.n10856 GND.n10855 19.3944
R21296 GND.n10855 GND.n10852 19.3944
R21297 GND.n10852 GND.n10851 19.3944
R21298 GND.n10851 GND.n10848 19.3944
R21299 GND.n10848 GND.n10847 19.3944
R21300 GND.n10718 GND.n10717 19.3944
R21301 GND.n10893 GND.n10717 19.3944
R21302 GND.n10893 GND.n10892 19.3944
R21303 GND.n10892 GND.n10891 19.3944
R21304 GND.n10891 GND.n10888 19.3944
R21305 GND.n10888 GND.n10887 19.3944
R21306 GND.n10887 GND.n10884 19.3944
R21307 GND.n10884 GND.n10883 19.3944
R21308 GND.n10883 GND.n10880 19.3944
R21309 GND.n10880 GND.n10879 19.3944
R21310 GND.n10879 GND.n10876 19.3944
R21311 GND.n10685 GND.n10653 19.3944
R21312 GND.n10685 GND.n10654 19.3944
R21313 GND.n10681 GND.n10654 19.3944
R21314 GND.n10681 GND.n10678 19.3944
R21315 GND.n10678 GND.n10677 19.3944
R21316 GND.n10677 GND.n10674 19.3944
R21317 GND.n10674 GND.n10673 19.3944
R21318 GND.n10673 GND.n10670 19.3944
R21319 GND.n10670 GND.n10669 19.3944
R21320 GND.n10669 GND.n10666 19.3944
R21321 GND.n10666 GND.n10665 19.3944
R21322 GND.n6741 GND.n6740 19.3944
R21323 GND.n6747 GND.n6741 19.3944
R21324 GND.n6747 GND.n6737 19.3944
R21325 GND.n6751 GND.n6737 19.3944
R21326 GND.n6751 GND.n6735 19.3944
R21327 GND.n6762 GND.n6735 19.3944
R21328 GND.n6762 GND.n6733 19.3944
R21329 GND.n6766 GND.n6733 19.3944
R21330 GND.n6766 GND.n6529 19.3944
R21331 GND.n6777 GND.n6529 19.3944
R21332 GND.n6777 GND.n6527 19.3944
R21333 GND.n6781 GND.n6527 19.3944
R21334 GND.n6781 GND.n6525 19.3944
R21335 GND.n6792 GND.n6525 19.3944
R21336 GND.n6792 GND.n6523 19.3944
R21337 GND.n6796 GND.n6523 19.3944
R21338 GND.n6796 GND.n6521 19.3944
R21339 GND.n6807 GND.n6521 19.3944
R21340 GND.n6807 GND.n6519 19.3944
R21341 GND.n6811 GND.n6519 19.3944
R21342 GND.n6811 GND.n6517 19.3944
R21343 GND.n6822 GND.n6517 19.3944
R21344 GND.n6822 GND.n6515 19.3944
R21345 GND.n6826 GND.n6515 19.3944
R21346 GND.n6826 GND.n6512 19.3944
R21347 GND.n6837 GND.n6512 19.3944
R21348 GND.n6837 GND.n6510 19.3944
R21349 GND.n6841 GND.n6510 19.3944
R21350 GND.n6841 GND.n6508 19.3944
R21351 GND.n6852 GND.n6508 19.3944
R21352 GND.n6852 GND.n6506 19.3944
R21353 GND.n6856 GND.n6506 19.3944
R21354 GND.n6856 GND.n6504 19.3944
R21355 GND.n6867 GND.n6504 19.3944
R21356 GND.n6867 GND.n6502 19.3944
R21357 GND.n6871 GND.n6502 19.3944
R21358 GND.n6871 GND.n6500 19.3944
R21359 GND.n6882 GND.n6500 19.3944
R21360 GND.n6882 GND.n6498 19.3944
R21361 GND.n6886 GND.n6498 19.3944
R21362 GND.n6886 GND.n6496 19.3944
R21363 GND.n6897 GND.n6496 19.3944
R21364 GND.n6897 GND.n6494 19.3944
R21365 GND.n6901 GND.n6494 19.3944
R21366 GND.n6901 GND.n6492 19.3944
R21367 GND.n6912 GND.n6492 19.3944
R21368 GND.n6912 GND.n6490 19.3944
R21369 GND.n6916 GND.n6490 19.3944
R21370 GND.n6916 GND.n6487 19.3944
R21371 GND.n6927 GND.n6487 19.3944
R21372 GND.n6927 GND.n6485 19.3944
R21373 GND.n6931 GND.n6485 19.3944
R21374 GND.n6931 GND.n6483 19.3944
R21375 GND.n6942 GND.n6483 19.3944
R21376 GND.n6942 GND.n6481 19.3944
R21377 GND.n6946 GND.n6481 19.3944
R21378 GND.n6946 GND.n6479 19.3944
R21379 GND.n6957 GND.n6479 19.3944
R21380 GND.n6957 GND.n6477 19.3944
R21381 GND.n6961 GND.n6477 19.3944
R21382 GND.n6961 GND.n6475 19.3944
R21383 GND.n6972 GND.n6475 19.3944
R21384 GND.n6972 GND.n6473 19.3944
R21385 GND.n6983 GND.n6473 19.3944
R21386 GND.n6983 GND.n6982 19.3944
R21387 GND.n6982 GND.n6981 19.3944
R21388 GND.n6981 GND.n6980 19.3944
R21389 GND.n6980 GND.n88 19.3944
R21390 GND.n11113 GND.n88 19.3944
R21391 GND.n11113 GND.n89 19.3944
R21392 GND.n6272 GND.n89 19.3944
R21393 GND.n7316 GND.n6272 19.3944
R21394 GND.n7316 GND.n7315 19.3944
R21395 GND.n7315 GND.n7314 19.3944
R21396 GND.n7314 GND.n6277 19.3944
R21397 GND.n7019 GND.n6277 19.3944
R21398 GND.n7019 GND.n6461 19.3944
R21399 GND.n7023 GND.n6461 19.3944
R21400 GND.n7023 GND.n6459 19.3944
R21401 GND.n7034 GND.n6459 19.3944
R21402 GND.n7034 GND.n6457 19.3944
R21403 GND.n7038 GND.n6457 19.3944
R21404 GND.n7038 GND.n6455 19.3944
R21405 GND.n7049 GND.n6455 19.3944
R21406 GND.n7049 GND.n6453 19.3944
R21407 GND.n7053 GND.n6453 19.3944
R21408 GND.n7053 GND.n6451 19.3944
R21409 GND.n7064 GND.n6451 19.3944
R21410 GND.n7064 GND.n6449 19.3944
R21411 GND.n7068 GND.n6449 19.3944
R21412 GND.n7068 GND.n6447 19.3944
R21413 GND.n7079 GND.n6447 19.3944
R21414 GND.n7079 GND.n6445 19.3944
R21415 GND.n7083 GND.n6445 19.3944
R21416 GND.n7083 GND.n6443 19.3944
R21417 GND.n7094 GND.n6443 19.3944
R21418 GND.n7094 GND.n6441 19.3944
R21419 GND.n7099 GND.n6441 19.3944
R21420 GND.n7099 GND.n6435 19.3944
R21421 GND.n7266 GND.n6435 19.3944
R21422 GND.n7266 GND.n7265 19.3944
R21423 GND.n7265 GND.n7264 19.3944
R21424 GND.n7264 GND.n6439 19.3944
R21425 GND.n7254 GND.n6439 19.3944
R21426 GND.n7254 GND.n7253 19.3944
R21427 GND.n7253 GND.n7252 19.3944
R21428 GND.n7252 GND.n7114 19.3944
R21429 GND.n7242 GND.n7114 19.3944
R21430 GND.n7242 GND.n7241 19.3944
R21431 GND.n7241 GND.n7240 19.3944
R21432 GND.n7240 GND.n7121 19.3944
R21433 GND.n7230 GND.n7121 19.3944
R21434 GND.n7230 GND.n7229 19.3944
R21435 GND.n7229 GND.n7228 19.3944
R21436 GND.n7228 GND.n7128 19.3944
R21437 GND.n7218 GND.n7128 19.3944
R21438 GND.n7218 GND.n7217 19.3944
R21439 GND.n7217 GND.n7216 19.3944
R21440 GND.n7216 GND.n7135 19.3944
R21441 GND.n7206 GND.n7135 19.3944
R21442 GND.n7206 GND.n7205 19.3944
R21443 GND.n7205 GND.n7204 19.3944
R21444 GND.n7204 GND.n7142 19.3944
R21445 GND.n7194 GND.n7142 19.3944
R21446 GND.n7194 GND.n7193 19.3944
R21447 GND.n7193 GND.n7192 19.3944
R21448 GND.n7192 GND.n7149 19.3944
R21449 GND.n7182 GND.n7149 19.3944
R21450 GND.n7182 GND.n7181 19.3944
R21451 GND.n7181 GND.n7180 19.3944
R21452 GND.n7180 GND.n7156 19.3944
R21453 GND.n7170 GND.n7156 19.3944
R21454 GND.n7170 GND.n7169 19.3944
R21455 GND.n7169 GND.n7168 19.3944
R21456 GND.n7168 GND.n453 19.3944
R21457 GND.n10903 GND.n453 19.3944
R21458 GND.n10903 GND.n10902 19.3944
R21459 GND.n3897 GND.n3880 19.3944
R21460 GND.n7997 GND.n3897 19.3944
R21461 GND.n7997 GND.n7996 19.3944
R21462 GND.n7996 GND.n7995 19.3944
R21463 GND.n7995 GND.n3903 19.3944
R21464 GND.n7985 GND.n3903 19.3944
R21465 GND.n7985 GND.n7984 19.3944
R21466 GND.n7984 GND.n7983 19.3944
R21467 GND.n7983 GND.n3922 19.3944
R21468 GND.n7973 GND.n3922 19.3944
R21469 GND.n7973 GND.n7972 19.3944
R21470 GND.n7972 GND.n7971 19.3944
R21471 GND.n7971 GND.n3942 19.3944
R21472 GND.n7961 GND.n3942 19.3944
R21473 GND.n7961 GND.n7960 19.3944
R21474 GND.n7960 GND.n7959 19.3944
R21475 GND.n7959 GND.n3962 19.3944
R21476 GND.n7949 GND.n3962 19.3944
R21477 GND.n7949 GND.n7948 19.3944
R21478 GND.n7948 GND.n7947 19.3944
R21479 GND.n7947 GND.n3982 19.3944
R21480 GND.n7937 GND.n3982 19.3944
R21481 GND.n7937 GND.n7936 19.3944
R21482 GND.n7936 GND.n7935 19.3944
R21483 GND.n7935 GND.n4002 19.3944
R21484 GND.n7925 GND.n4002 19.3944
R21485 GND.n7925 GND.n7924 19.3944
R21486 GND.n7924 GND.n7923 19.3944
R21487 GND.n7923 GND.n4022 19.3944
R21488 GND.n7913 GND.n4022 19.3944
R21489 GND.n7913 GND.n7912 19.3944
R21490 GND.n7912 GND.n7911 19.3944
R21491 GND.n7911 GND.n4042 19.3944
R21492 GND.n4093 GND.n4042 19.3944
R21493 GND.n4097 GND.n4093 19.3944
R21494 GND.n4100 GND.n4097 19.3944
R21495 GND.n4101 GND.n4100 19.3944
R21496 GND.n4101 GND.n4091 19.3944
R21497 GND.n7882 GND.n4091 19.3944
R21498 GND.n7882 GND.n7881 19.3944
R21499 GND.n7881 GND.n7880 19.3944
R21500 GND.n7880 GND.n4107 19.3944
R21501 GND.n7870 GND.n4107 19.3944
R21502 GND.n7870 GND.n7869 19.3944
R21503 GND.n7869 GND.n7868 19.3944
R21504 GND.n7868 GND.n4127 19.3944
R21505 GND.n7858 GND.n4127 19.3944
R21506 GND.n7858 GND.n7857 19.3944
R21507 GND.n7857 GND.n7856 19.3944
R21508 GND.n7856 GND.n4147 19.3944
R21509 GND.n4197 GND.n4147 19.3944
R21510 GND.n4201 GND.n4197 19.3944
R21511 GND.n4204 GND.n4201 19.3944
R21512 GND.n4205 GND.n4204 19.3944
R21513 GND.n4205 GND.n4195 19.3944
R21514 GND.n7827 GND.n4195 19.3944
R21515 GND.n7827 GND.n7826 19.3944
R21516 GND.n7826 GND.n7825 19.3944
R21517 GND.n7825 GND.n4211 19.3944
R21518 GND.n7815 GND.n4211 19.3944
R21519 GND.n7815 GND.n7814 19.3944
R21520 GND.n7814 GND.n7813 19.3944
R21521 GND.n7813 GND.n4231 19.3944
R21522 GND.n7803 GND.n4231 19.3944
R21523 GND.n7803 GND.n7802 19.3944
R21524 GND.n7802 GND.n7801 19.3944
R21525 GND.n7801 GND.n4249 19.3944
R21526 GND.n4300 GND.n4249 19.3944
R21527 GND.n4304 GND.n4300 19.3944
R21528 GND.n4307 GND.n4304 19.3944
R21529 GND.n4308 GND.n4307 19.3944
R21530 GND.n4308 GND.n4298 19.3944
R21531 GND.n7772 GND.n4298 19.3944
R21532 GND.n7772 GND.n7771 19.3944
R21533 GND.n7771 GND.n7770 19.3944
R21534 GND.n7770 GND.n4314 19.3944
R21535 GND.n7760 GND.n4314 19.3944
R21536 GND.n7760 GND.n7759 19.3944
R21537 GND.n7759 GND.n7758 19.3944
R21538 GND.n7758 GND.n4334 19.3944
R21539 GND.n7748 GND.n4334 19.3944
R21540 GND.n7748 GND.n7747 19.3944
R21541 GND.n7747 GND.n7746 19.3944
R21542 GND.n7746 GND.n4353 19.3944
R21543 GND.n4832 GND.n4353 19.3944
R21544 GND.n5028 GND.n5023 19.3944
R21545 GND.n5029 GND.n5028 19.3944
R21546 GND.n5326 GND.n5029 19.3944
R21547 GND.n5326 GND.n5021 19.3944
R21548 GND.n5330 GND.n5021 19.3944
R21549 GND.n5330 GND.n5014 19.3944
R21550 GND.n5345 GND.n5014 19.3944
R21551 GND.n5345 GND.n5012 19.3944
R21552 GND.n5349 GND.n5012 19.3944
R21553 GND.n5349 GND.n5005 19.3944
R21554 GND.n5364 GND.n5005 19.3944
R21555 GND.n5364 GND.n5003 19.3944
R21556 GND.n5409 GND.n5003 19.3944
R21557 GND.n5409 GND.n5408 19.3944
R21558 GND.n5408 GND.n5407 19.3944
R21559 GND.n5407 GND.n5405 19.3944
R21560 GND.n5405 GND.n5404 19.3944
R21561 GND.n5404 GND.n5403 19.3944
R21562 GND.n5403 GND.n5402 19.3944
R21563 GND.n5402 GND.n5400 19.3944
R21564 GND.n5400 GND.n5399 19.3944
R21565 GND.n5399 GND.n5396 19.3944
R21566 GND.n5396 GND.n5395 19.3944
R21567 GND.n5395 GND.n5393 19.3944
R21568 GND.n5393 GND.n5392 19.3944
R21569 GND.n5392 GND.n5390 19.3944
R21570 GND.n5390 GND.n5389 19.3944
R21571 GND.n5389 GND.n5387 19.3944
R21572 GND.n5387 GND.n5386 19.3944
R21573 GND.n5386 GND.n4957 19.3944
R21574 GND.n5506 GND.n4957 19.3944
R21575 GND.n5507 GND.n5506 19.3944
R21576 GND.n5507 GND.n4955 19.3944
R21577 GND.n5511 GND.n4955 19.3944
R21578 GND.n5512 GND.n5511 19.3944
R21579 GND.n5515 GND.n5512 19.3944
R21580 GND.n5515 GND.n4951 19.3944
R21581 GND.n5540 GND.n4951 19.3944
R21582 GND.n5540 GND.n5539 19.3944
R21583 GND.n5539 GND.n5538 19.3944
R21584 GND.n5538 GND.n5536 19.3944
R21585 GND.n5536 GND.n5535 19.3944
R21586 GND.n5535 GND.n5533 19.3944
R21587 GND.n5533 GND.n5532 19.3944
R21588 GND.n5532 GND.n5530 19.3944
R21589 GND.n5530 GND.n5529 19.3944
R21590 GND.n5529 GND.n4926 19.3944
R21591 GND.n5609 GND.n4926 19.3944
R21592 GND.n5610 GND.n5609 19.3944
R21593 GND.n5610 GND.n4924 19.3944
R21594 GND.n5614 GND.n4924 19.3944
R21595 GND.n5615 GND.n5614 19.3944
R21596 GND.n5618 GND.n5615 19.3944
R21597 GND.n5618 GND.n4920 19.3944
R21598 GND.n5644 GND.n4920 19.3944
R21599 GND.n5644 GND.n5643 19.3944
R21600 GND.n5643 GND.n5642 19.3944
R21601 GND.n5642 GND.n5640 19.3944
R21602 GND.n5640 GND.n5639 19.3944
R21603 GND.n5639 GND.n5637 19.3944
R21604 GND.n5637 GND.n5636 19.3944
R21605 GND.n5636 GND.n5634 19.3944
R21606 GND.n5634 GND.n5633 19.3944
R21607 GND.n5633 GND.n4892 19.3944
R21608 GND.n5712 GND.n4892 19.3944
R21609 GND.n5713 GND.n5712 19.3944
R21610 GND.n5713 GND.n4890 19.3944
R21611 GND.n5717 GND.n4890 19.3944
R21612 GND.n5718 GND.n5717 19.3944
R21613 GND.n5721 GND.n5718 19.3944
R21614 GND.n5721 GND.n4886 19.3944
R21615 GND.n5741 GND.n4886 19.3944
R21616 GND.n5741 GND.n5740 19.3944
R21617 GND.n5740 GND.n5739 19.3944
R21618 GND.n5739 GND.n5737 19.3944
R21619 GND.n5737 GND.n5736 19.3944
R21620 GND.n5736 GND.n5734 19.3944
R21621 GND.n5734 GND.n5733 19.3944
R21622 GND.n5733 GND.n4852 19.3944
R21623 GND.n5803 GND.n4852 19.3944
R21624 GND.n5804 GND.n5803 19.3944
R21625 GND.n5804 GND.n4850 19.3944
R21626 GND.n5808 GND.n4850 19.3944
R21627 GND.n5811 GND.n5808 19.3944
R21628 GND.n5812 GND.n5811 19.3944
R21629 GND.n8053 GND.n8052 19.3944
R21630 GND.n8052 GND.n8051 19.3944
R21631 GND.n8051 GND.n8050 19.3944
R21632 GND.n8050 GND.n8048 19.3944
R21633 GND.n8048 GND.n8045 19.3944
R21634 GND.n8045 GND.n8044 19.3944
R21635 GND.n8044 GND.n3873 19.3944
R21636 GND.n8041 GND.n8040 19.3944
R21637 GND.n8036 GND.n8035 19.3944
R21638 GND.n8031 GND.n8030 19.3944
R21639 GND.n8026 GND.n8025 19.3944
R21640 GND.n8021 GND.n8020 19.3944
R21641 GND.n3876 GND.n3875 19.3944
R21642 GND.n8009 GND.n8008 19.3944
R21643 GND.n5871 GND.n4843 19.3944
R21644 GND.n5871 GND.n4844 19.3944
R21645 GND.n5819 GND.n5815 19.3944
R21646 GND.n5819 GND.n4848 19.3944
R21647 GND.n5824 GND.n4848 19.3944
R21648 GND.n5824 GND.n4846 19.3944
R21649 GND.n5829 GND.n4846 19.3944
R21650 GND.n5830 GND.n5829 19.3944
R21651 GND.n5832 GND.n4841 19.3944
R21652 GND.n5836 GND.n4841 19.3944
R21653 GND.n5841 GND.n5840 19.3944
R21654 GND.n5846 GND.n5845 19.3944
R21655 GND.n5851 GND.n5850 19.3944
R21656 GND.n5856 GND.n5855 19.3944
R21657 GND.n5914 GND.n5911 19.3944
R21658 GND.n5909 GND.n5906 19.3944
R21659 GND.n5904 GND.n5901 19.3944
R21660 GND.n5899 GND.n5896 19.3944
R21661 GND.n5894 GND.n5891 19.3944
R21662 GND.n7527 GND.n5922 19.3944
R21663 GND.n7527 GND.n7526 19.3944
R21664 GND.n7526 GND.n7525 19.3944
R21665 GND.n7525 GND.n5927 19.3944
R21666 GND.n7515 GND.n5927 19.3944
R21667 GND.n7515 GND.n7514 19.3944
R21668 GND.n7514 GND.n7513 19.3944
R21669 GND.n7513 GND.n5949 19.3944
R21670 GND.n7503 GND.n5949 19.3944
R21671 GND.n7503 GND.n7502 19.3944
R21672 GND.n7502 GND.n7501 19.3944
R21673 GND.n7501 GND.n5969 19.3944
R21674 GND.n7491 GND.n5969 19.3944
R21675 GND.n7491 GND.n7490 19.3944
R21676 GND.n7490 GND.n7489 19.3944
R21677 GND.n7489 GND.n5990 19.3944
R21678 GND.n7479 GND.n5990 19.3944
R21679 GND.n7479 GND.n7478 19.3944
R21680 GND.n7478 GND.n7477 19.3944
R21681 GND.n7477 GND.n6011 19.3944
R21682 GND.n7467 GND.n6011 19.3944
R21683 GND.n7467 GND.n7466 19.3944
R21684 GND.n7466 GND.n7465 19.3944
R21685 GND.n7465 GND.n6032 19.3944
R21686 GND.n7455 GND.n6032 19.3944
R21687 GND.n7455 GND.n7454 19.3944
R21688 GND.n7454 GND.n7453 19.3944
R21689 GND.n7453 GND.n6052 19.3944
R21690 GND.n7443 GND.n6052 19.3944
R21691 GND.n7443 GND.n7442 19.3944
R21692 GND.n7442 GND.n7441 19.3944
R21693 GND.n7441 GND.n6073 19.3944
R21694 GND.n7431 GND.n6073 19.3944
R21695 GND.n7431 GND.n7430 19.3944
R21696 GND.n7430 GND.n7429 19.3944
R21697 GND.n7429 GND.n6094 19.3944
R21698 GND.n7419 GND.n6094 19.3944
R21699 GND.n7419 GND.n7418 19.3944
R21700 GND.n7418 GND.n7417 19.3944
R21701 GND.n7417 GND.n6115 19.3944
R21702 GND.n7407 GND.n6115 19.3944
R21703 GND.n7407 GND.n7406 19.3944
R21704 GND.n7406 GND.n7405 19.3944
R21705 GND.n7405 GND.n6136 19.3944
R21706 GND.n7395 GND.n6136 19.3944
R21707 GND.n7395 GND.n7394 19.3944
R21708 GND.n7394 GND.n7393 19.3944
R21709 GND.n7393 GND.n6157 19.3944
R21710 GND.n7383 GND.n6157 19.3944
R21711 GND.n7383 GND.n7382 19.3944
R21712 GND.n7382 GND.n7381 19.3944
R21713 GND.n7381 GND.n6177 19.3944
R21714 GND.n7371 GND.n6177 19.3944
R21715 GND.n7371 GND.n7370 19.3944
R21716 GND.n7370 GND.n7369 19.3944
R21717 GND.n7369 GND.n6198 19.3944
R21718 GND.n7359 GND.n6198 19.3944
R21719 GND.n7359 GND.n7358 19.3944
R21720 GND.n7358 GND.n7357 19.3944
R21721 GND.n7357 GND.n6219 19.3944
R21722 GND.n7347 GND.n6219 19.3944
R21723 GND.n7347 GND.n7346 19.3944
R21724 GND.n7346 GND.n7345 19.3944
R21725 GND.n7345 GND.n6239 19.3944
R21726 GND.n7335 GND.n105 19.3944
R21727 GND.n6255 GND.n105 19.3944
R21728 GND.n11109 GND.n98 19.3944
R21729 GND.n6267 GND.n99 19.3944
R21730 GND.n11106 GND.n107 19.3944
R21731 GND.n11106 GND.n108 19.3944
R21732 GND.n11096 GND.n108 19.3944
R21733 GND.n11096 GND.n11095 19.3944
R21734 GND.n11095 GND.n11094 19.3944
R21735 GND.n11094 GND.n130 19.3944
R21736 GND.n11084 GND.n130 19.3944
R21737 GND.n11084 GND.n11083 19.3944
R21738 GND.n11083 GND.n11082 19.3944
R21739 GND.n11082 GND.n151 19.3944
R21740 GND.n11072 GND.n151 19.3944
R21741 GND.n11072 GND.n11071 19.3944
R21742 GND.n11071 GND.n11070 19.3944
R21743 GND.n11070 GND.n172 19.3944
R21744 GND.n11060 GND.n172 19.3944
R21745 GND.n11060 GND.n11059 19.3944
R21746 GND.n11059 GND.n11058 19.3944
R21747 GND.n11058 GND.n193 19.3944
R21748 GND.n11048 GND.n193 19.3944
R21749 GND.n11048 GND.n11047 19.3944
R21750 GND.n11047 GND.n11046 19.3944
R21751 GND.n11046 GND.n214 19.3944
R21752 GND.n11036 GND.n214 19.3944
R21753 GND.n11036 GND.n11035 19.3944
R21754 GND.n11035 GND.n11034 19.3944
R21755 GND.n11034 GND.n235 19.3944
R21756 GND.n11024 GND.n235 19.3944
R21757 GND.n11024 GND.n11023 19.3944
R21758 GND.n11023 GND.n11022 19.3944
R21759 GND.n11022 GND.n256 19.3944
R21760 GND.n11012 GND.n256 19.3944
R21761 GND.n11012 GND.n11011 19.3944
R21762 GND.n11011 GND.n11010 19.3944
R21763 GND.n11010 GND.n276 19.3944
R21764 GND.n11000 GND.n276 19.3944
R21765 GND.n11000 GND.n10999 19.3944
R21766 GND.n10999 GND.n10998 19.3944
R21767 GND.n10998 GND.n297 19.3944
R21768 GND.n10988 GND.n297 19.3944
R21769 GND.n10988 GND.n10987 19.3944
R21770 GND.n10987 GND.n10986 19.3944
R21771 GND.n10986 GND.n318 19.3944
R21772 GND.n10976 GND.n318 19.3944
R21773 GND.n10976 GND.n10975 19.3944
R21774 GND.n10975 GND.n10974 19.3944
R21775 GND.n10974 GND.n339 19.3944
R21776 GND.n10964 GND.n339 19.3944
R21777 GND.n10964 GND.n10963 19.3944
R21778 GND.n10963 GND.n10962 19.3944
R21779 GND.n10962 GND.n360 19.3944
R21780 GND.n10952 GND.n360 19.3944
R21781 GND.n10952 GND.n10951 19.3944
R21782 GND.n10951 GND.n10950 19.3944
R21783 GND.n10950 GND.n381 19.3944
R21784 GND.n10940 GND.n381 19.3944
R21785 GND.n10940 GND.n10939 19.3944
R21786 GND.n10939 GND.n10938 19.3944
R21787 GND.n10938 GND.n402 19.3944
R21788 GND.n10928 GND.n402 19.3944
R21789 GND.n10928 GND.n10927 19.3944
R21790 GND.n10927 GND.n10926 19.3944
R21791 GND.n10926 GND.n423 19.3944
R21792 GND.n10916 GND.n423 19.3944
R21793 GND.n10916 GND.n10915 19.3944
R21794 GND.n10915 GND.n10914 19.3944
R21795 GND.n8813 GND.n8812 19.3944
R21796 GND.n8812 GND.n8811 19.3944
R21797 GND.n8811 GND.n8810 19.3944
R21798 GND.n8810 GND.n8808 19.3944
R21799 GND.n8808 GND.n8805 19.3944
R21800 GND.n8805 GND.n8804 19.3944
R21801 GND.n8804 GND.n8801 19.3944
R21802 GND.n8801 GND.n8800 19.3944
R21803 GND.n8800 GND.n8797 19.3944
R21804 GND.n8797 GND.n8796 19.3944
R21805 GND.n8796 GND.n8793 19.3944
R21806 GND.n8791 GND.n8789 19.3944
R21807 GND.n8789 GND.n8786 19.3944
R21808 GND.n8786 GND.n8785 19.3944
R21809 GND.n8785 GND.n8782 19.3944
R21810 GND.n8782 GND.n8781 19.3944
R21811 GND.n8781 GND.n8778 19.3944
R21812 GND.n8778 GND.n8777 19.3944
R21813 GND.n8777 GND.n8774 19.3944
R21814 GND.n8774 GND.n8773 19.3944
R21815 GND.n8773 GND.n8770 19.3944
R21816 GND.n8770 GND.n8769 19.3944
R21817 GND.n8769 GND.n8766 19.3944
R21818 GND.n8766 GND.n8765 19.3944
R21819 GND.n8762 GND.n8761 19.3944
R21820 GND.n8761 GND.n8758 19.3944
R21821 GND.n8758 GND.n8757 19.3944
R21822 GND.n8757 GND.n8754 19.3944
R21823 GND.n8754 GND.n8753 19.3944
R21824 GND.n8753 GND.n8750 19.3944
R21825 GND.n8750 GND.n8749 19.3944
R21826 GND.n8749 GND.n8746 19.3944
R21827 GND.n8746 GND.n8745 19.3944
R21828 GND.n8745 GND.n8742 19.3944
R21829 GND.n8742 GND.n8741 19.3944
R21830 GND.n8741 GND.n8738 19.3944
R21831 GND.n8738 GND.n8737 19.3944
R21832 GND.n8734 GND.n8733 19.3944
R21833 GND.n8733 GND.n8730 19.3944
R21834 GND.n8730 GND.n8729 19.3944
R21835 GND.n8729 GND.n8726 19.3944
R21836 GND.n8726 GND.n8725 19.3944
R21837 GND.n8725 GND.n8722 19.3944
R21838 GND.n8722 GND.n8721 19.3944
R21839 GND.n8721 GND.n8718 19.3944
R21840 GND.n8718 GND.n8717 19.3944
R21841 GND.n8717 GND.n8714 19.3944
R21842 GND.n8714 GND.n8713 19.3944
R21843 GND.n8713 GND.n8710 19.3944
R21844 GND.n8710 GND.n8709 19.3944
R21845 GND.n1828 GND.n1826 19.3944
R21846 GND.n1828 GND.n1824 19.3944
R21847 GND.n8688 GND.n1824 19.3944
R21848 GND.n8688 GND.n8687 19.3944
R21849 GND.n8687 GND.n8686 19.3944
R21850 GND.n8686 GND.n1834 19.3944
R21851 GND.n3158 GND.n1834 19.3944
R21852 GND.n3158 GND.n3157 19.3944
R21853 GND.n3157 GND.n2895 19.3944
R21854 GND.n3177 GND.n2895 19.3944
R21855 GND.n3177 GND.n2893 19.3944
R21856 GND.n3183 GND.n2893 19.3944
R21857 GND.n3183 GND.n3182 19.3944
R21858 GND.n3182 GND.n2872 19.3944
R21859 GND.n3202 GND.n2872 19.3944
R21860 GND.n3202 GND.n2870 19.3944
R21861 GND.n3208 GND.n2870 19.3944
R21862 GND.n3208 GND.n3207 19.3944
R21863 GND.n3207 GND.n2849 19.3944
R21864 GND.n3226 GND.n2849 19.3944
R21865 GND.n3226 GND.n2847 19.3944
R21866 GND.n3232 GND.n2847 19.3944
R21867 GND.n3232 GND.n3231 19.3944
R21868 GND.n3231 GND.n2826 19.3944
R21869 GND.n3251 GND.n2826 19.3944
R21870 GND.n3251 GND.n2824 19.3944
R21871 GND.n3257 GND.n2824 19.3944
R21872 GND.n3257 GND.n3256 19.3944
R21873 GND.n3256 GND.n2804 19.3944
R21874 GND.n3276 GND.n2804 19.3944
R21875 GND.n3276 GND.n2802 19.3944
R21876 GND.n3282 GND.n2802 19.3944
R21877 GND.n3282 GND.n3281 19.3944
R21878 GND.n3281 GND.n2781 19.3944
R21879 GND.n3301 GND.n2781 19.3944
R21880 GND.n3301 GND.n2779 19.3944
R21881 GND.n3307 GND.n2779 19.3944
R21882 GND.n3307 GND.n3306 19.3944
R21883 GND.n3306 GND.n2758 19.3944
R21884 GND.n3325 GND.n2758 19.3944
R21885 GND.n3325 GND.n2756 19.3944
R21886 GND.n3331 GND.n2756 19.3944
R21887 GND.n3331 GND.n3330 19.3944
R21888 GND.n3330 GND.n2735 19.3944
R21889 GND.n3350 GND.n2735 19.3944
R21890 GND.n3350 GND.n2733 19.3944
R21891 GND.n3356 GND.n2733 19.3944
R21892 GND.n3356 GND.n3355 19.3944
R21893 GND.n3355 GND.n2713 19.3944
R21894 GND.n3375 GND.n2713 19.3944
R21895 GND.n3375 GND.n2711 19.3944
R21896 GND.n3381 GND.n2711 19.3944
R21897 GND.n3381 GND.n3380 19.3944
R21898 GND.n3380 GND.n2690 19.3944
R21899 GND.n3400 GND.n2690 19.3944
R21900 GND.n3400 GND.n2688 19.3944
R21901 GND.n3406 GND.n2688 19.3944
R21902 GND.n3406 GND.n3405 19.3944
R21903 GND.n3405 GND.n2667 19.3944
R21904 GND.n3424 GND.n2667 19.3944
R21905 GND.n3424 GND.n2665 19.3944
R21906 GND.n3428 GND.n2665 19.3944
R21907 GND.n3428 GND.n2498 19.3944
R21908 GND.n3492 GND.n2498 19.3944
R21909 GND.n2497 GND.n2496 19.3944
R21910 GND.n2523 GND.n2496 19.3944
R21911 GND.n3476 GND.n3475 19.3944
R21912 GND.n3454 GND.n3453 19.3944
R21913 GND.n3456 GND.n2490 19.3944
R21914 GND.n3498 GND.n2490 19.3944
R21915 GND.n3498 GND.n3497 19.3944
R21916 GND.n3497 GND.n2470 19.3944
R21917 GND.n3518 GND.n2470 19.3944
R21918 GND.n3518 GND.n2468 19.3944
R21919 GND.n3524 GND.n2468 19.3944
R21920 GND.n3524 GND.n3523 19.3944
R21921 GND.n3523 GND.n2449 19.3944
R21922 GND.n3544 GND.n2449 19.3944
R21923 GND.n3544 GND.n2447 19.3944
R21924 GND.n3550 GND.n2447 19.3944
R21925 GND.n3550 GND.n3549 19.3944
R21926 GND.n3549 GND.n2427 19.3944
R21927 GND.n3570 GND.n2427 19.3944
R21928 GND.n3570 GND.n2425 19.3944
R21929 GND.n3576 GND.n2425 19.3944
R21930 GND.n3576 GND.n3575 19.3944
R21931 GND.n3575 GND.n2405 19.3944
R21932 GND.n3595 GND.n2405 19.3944
R21933 GND.n3595 GND.n2403 19.3944
R21934 GND.n3601 GND.n2403 19.3944
R21935 GND.n3601 GND.n3600 19.3944
R21936 GND.n3600 GND.n2383 19.3944
R21937 GND.n3621 GND.n2383 19.3944
R21938 GND.n3621 GND.n2381 19.3944
R21939 GND.n3627 GND.n2381 19.3944
R21940 GND.n3627 GND.n3626 19.3944
R21941 GND.n3626 GND.n2365 19.3944
R21942 GND.n3647 GND.n2365 19.3944
R21943 GND.n3647 GND.n2363 19.3944
R21944 GND.n3653 GND.n2363 19.3944
R21945 GND.n3653 GND.n3652 19.3944
R21946 GND.n3652 GND.n2343 19.3944
R21947 GND.n3673 GND.n2343 19.3944
R21948 GND.n3673 GND.n2341 19.3944
R21949 GND.n3679 GND.n2341 19.3944
R21950 GND.n3679 GND.n3678 19.3944
R21951 GND.n3678 GND.n2315 19.3944
R21952 GND.n8184 GND.n2315 19.3944
R21953 GND.n8184 GND.n2313 19.3944
R21954 GND.n8190 GND.n2313 19.3944
R21955 GND.n8190 GND.n8189 19.3944
R21956 GND.n8189 GND.n2294 19.3944
R21957 GND.n8210 GND.n2294 19.3944
R21958 GND.n8210 GND.n2292 19.3944
R21959 GND.n8216 GND.n2292 19.3944
R21960 GND.n8216 GND.n8215 19.3944
R21961 GND.n8215 GND.n2273 19.3944
R21962 GND.n8236 GND.n2273 19.3944
R21963 GND.n8236 GND.n2271 19.3944
R21964 GND.n8242 GND.n2271 19.3944
R21965 GND.n8242 GND.n8241 19.3944
R21966 GND.n8241 GND.n2251 19.3944
R21967 GND.n8262 GND.n2251 19.3944
R21968 GND.n8262 GND.n2249 19.3944
R21969 GND.n8268 GND.n2249 19.3944
R21970 GND.n8268 GND.n8267 19.3944
R21971 GND.n8267 GND.n2229 19.3944
R21972 GND.n8287 GND.n2229 19.3944
R21973 GND.n8287 GND.n2227 19.3944
R21974 GND.n8292 GND.n2227 19.3944
R21975 GND.n8292 GND.n2212 19.3944
R21976 GND.n8306 GND.n2212 19.3944
R21977 GND.n8307 GND.n8306 19.3944
R21978 GND.n8928 GND.n8927 19.3944
R21979 GND.n8927 GND.n1582 19.3944
R21980 GND.n8923 GND.n1582 19.3944
R21981 GND.n8923 GND.n1584 19.3944
R21982 GND.n8917 GND.n1584 19.3944
R21983 GND.n8917 GND.n8916 19.3944
R21984 GND.n8916 GND.n8915 19.3944
R21985 GND.n8915 GND.n1593 19.3944
R21986 GND.n8909 GND.n1593 19.3944
R21987 GND.n8909 GND.n8908 19.3944
R21988 GND.n8908 GND.n8907 19.3944
R21989 GND.n8907 GND.n1601 19.3944
R21990 GND.n8901 GND.n1601 19.3944
R21991 GND.n8901 GND.n8900 19.3944
R21992 GND.n8900 GND.n8899 19.3944
R21993 GND.n8899 GND.n1609 19.3944
R21994 GND.n8893 GND.n1609 19.3944
R21995 GND.n8893 GND.n8892 19.3944
R21996 GND.n8892 GND.n8891 19.3944
R21997 GND.n8891 GND.n1617 19.3944
R21998 GND.n8885 GND.n1617 19.3944
R21999 GND.n8885 GND.n8884 19.3944
R22000 GND.n8884 GND.n8883 19.3944
R22001 GND.n8883 GND.n1625 19.3944
R22002 GND.n8877 GND.n1625 19.3944
R22003 GND.n8877 GND.n8876 19.3944
R22004 GND.n8876 GND.n8875 19.3944
R22005 GND.n8875 GND.n1633 19.3944
R22006 GND.n8869 GND.n1633 19.3944
R22007 GND.n8869 GND.n8868 19.3944
R22008 GND.n8868 GND.n8867 19.3944
R22009 GND.n8867 GND.n1641 19.3944
R22010 GND.n8861 GND.n1641 19.3944
R22011 GND.n8861 GND.n8860 19.3944
R22012 GND.n8860 GND.n8859 19.3944
R22013 GND.n8859 GND.n1649 19.3944
R22014 GND.n8853 GND.n1649 19.3944
R22015 GND.n8853 GND.n8852 19.3944
R22016 GND.n8852 GND.n8851 19.3944
R22017 GND.n8851 GND.n1657 19.3944
R22018 GND.n8845 GND.n1657 19.3944
R22019 GND.n8845 GND.n8844 19.3944
R22020 GND.n8844 GND.n8843 19.3944
R22021 GND.n8843 GND.n1665 19.3944
R22022 GND.n8837 GND.n1665 19.3944
R22023 GND.n8837 GND.n8836 19.3944
R22024 GND.n8836 GND.n8835 19.3944
R22025 GND.n8835 GND.n1673 19.3944
R22026 GND.n8829 GND.n1673 19.3944
R22027 GND.n8829 GND.n8828 19.3944
R22028 GND.n8828 GND.n8827 19.3944
R22029 GND.n8827 GND.n1681 19.3944
R22030 GND.n8821 GND.n1681 19.3944
R22031 GND.n8821 GND.n8820 19.3944
R22032 GND.n8820 GND.n8819 19.3944
R22033 GND.n8819 GND.n1689 19.3944
R22034 GND.n1808 GND.n1689 19.3944
R22035 GND.n8695 GND.n1808 19.3944
R22036 GND.n8695 GND.n8694 19.3944
R22037 GND.n8694 GND.n8693 19.3944
R22038 GND.n8693 GND.n1814 19.3944
R22039 GND.n2972 GND.n1814 19.3944
R22040 GND.n2975 GND.n2972 19.3944
R22041 GND.n2975 GND.n2969 19.3944
R22042 GND.n3148 GND.n2969 19.3944
R22043 GND.n3148 GND.n3147 19.3944
R22044 GND.n3147 GND.n3146 19.3944
R22045 GND.n3146 GND.n2981 19.3944
R22046 GND.n3142 GND.n2981 19.3944
R22047 GND.n3142 GND.n3141 19.3944
R22048 GND.n3141 GND.n3140 19.3944
R22049 GND.n3140 GND.n2987 19.3944
R22050 GND.n3136 GND.n2987 19.3944
R22051 GND.n3136 GND.n3135 19.3944
R22052 GND.n3135 GND.n3134 19.3944
R22053 GND.n3134 GND.n2993 19.3944
R22054 GND.n3130 GND.n2993 19.3944
R22055 GND.n3130 GND.n3129 19.3944
R22056 GND.n3129 GND.n3128 19.3944
R22057 GND.n3128 GND.n2999 19.3944
R22058 GND.n3124 GND.n2999 19.3944
R22059 GND.n3124 GND.n3123 19.3944
R22060 GND.n3123 GND.n3122 19.3944
R22061 GND.n3122 GND.n3005 19.3944
R22062 GND.n3118 GND.n3005 19.3944
R22063 GND.n3118 GND.n3117 19.3944
R22064 GND.n3117 GND.n3116 19.3944
R22065 GND.n3116 GND.n3011 19.3944
R22066 GND.n3112 GND.n3011 19.3944
R22067 GND.n3112 GND.n3111 19.3944
R22068 GND.n3111 GND.n3110 19.3944
R22069 GND.n3110 GND.n3017 19.3944
R22070 GND.n3106 GND.n3017 19.3944
R22071 GND.n3106 GND.n3105 19.3944
R22072 GND.n3105 GND.n3104 19.3944
R22073 GND.n3104 GND.n3023 19.3944
R22074 GND.n3100 GND.n3023 19.3944
R22075 GND.n3100 GND.n3099 19.3944
R22076 GND.n3099 GND.n3098 19.3944
R22077 GND.n3098 GND.n3029 19.3944
R22078 GND.n3094 GND.n3029 19.3944
R22079 GND.n3094 GND.n3093 19.3944
R22080 GND.n3093 GND.n3092 19.3944
R22081 GND.n3092 GND.n3035 19.3944
R22082 GND.n3088 GND.n3035 19.3944
R22083 GND.n3088 GND.n3087 19.3944
R22084 GND.n3087 GND.n3086 19.3944
R22085 GND.n3086 GND.n3041 19.3944
R22086 GND.n3082 GND.n3041 19.3944
R22087 GND.n3082 GND.n3081 19.3944
R22088 GND.n3081 GND.n3080 19.3944
R22089 GND.n3080 GND.n3047 19.3944
R22090 GND.n3076 GND.n3047 19.3944
R22091 GND.n3076 GND.n3075 19.3944
R22092 GND.n3075 GND.n3074 19.3944
R22093 GND.n3074 GND.n3053 19.3944
R22094 GND.n3070 GND.n3053 19.3944
R22095 GND.n3070 GND.n3069 19.3944
R22096 GND.n3069 GND.n3068 19.3944
R22097 GND.n3068 GND.n3060 19.3944
R22098 GND.n3062 GND.n3060 19.3944
R22099 GND.n3484 GND.n2512 19.3944
R22100 GND.n3484 GND.n3483 19.3944
R22101 GND.n3481 GND.n2513 19.3944
R22102 GND.n3467 GND.n2535 19.3944
R22103 GND.n3465 GND.n3464 19.3944
R22104 GND.n2647 GND.n2646 19.3944
R22105 GND.n2646 GND.n2645 19.3944
R22106 GND.n2645 GND.n2540 19.3944
R22107 GND.n2641 GND.n2540 19.3944
R22108 GND.n2641 GND.n2640 19.3944
R22109 GND.n2640 GND.n2639 19.3944
R22110 GND.n2639 GND.n2546 19.3944
R22111 GND.n2635 GND.n2546 19.3944
R22112 GND.n2635 GND.n2634 19.3944
R22113 GND.n2634 GND.n2633 19.3944
R22114 GND.n2633 GND.n2552 19.3944
R22115 GND.n2629 GND.n2552 19.3944
R22116 GND.n2629 GND.n2628 19.3944
R22117 GND.n2628 GND.n2627 19.3944
R22118 GND.n2627 GND.n2558 19.3944
R22119 GND.n2623 GND.n2558 19.3944
R22120 GND.n2623 GND.n2622 19.3944
R22121 GND.n2622 GND.n2621 19.3944
R22122 GND.n2621 GND.n2564 19.3944
R22123 GND.n2617 GND.n2564 19.3944
R22124 GND.n2617 GND.n2616 19.3944
R22125 GND.n2616 GND.n2615 19.3944
R22126 GND.n2615 GND.n2570 19.3944
R22127 GND.n2611 GND.n2570 19.3944
R22128 GND.n2611 GND.n2610 19.3944
R22129 GND.n2610 GND.n2609 19.3944
R22130 GND.n2609 GND.n2576 19.3944
R22131 GND.n2602 GND.n2576 19.3944
R22132 GND.n2602 GND.n2601 19.3944
R22133 GND.n2601 GND.n2600 19.3944
R22134 GND.n2600 GND.n2582 19.3944
R22135 GND.n2596 GND.n2582 19.3944
R22136 GND.n2596 GND.n2595 19.3944
R22137 GND.n2595 GND.n2594 19.3944
R22138 GND.n2594 GND.n2591 19.3944
R22139 GND.n2591 GND.n2590 19.3944
R22140 GND.n2590 GND.n2326 19.3944
R22141 GND.n3695 GND.n2326 19.3944
R22142 GND.n3695 GND.n2324 19.3944
R22143 GND.n8176 GND.n2324 19.3944
R22144 GND.n8176 GND.n8175 19.3944
R22145 GND.n8175 GND.n8174 19.3944
R22146 GND.n8174 GND.n3701 19.3944
R22147 GND.n8170 GND.n3701 19.3944
R22148 GND.n8170 GND.n8169 19.3944
R22149 GND.n8169 GND.n8168 19.3944
R22150 GND.n8168 GND.n3707 19.3944
R22151 GND.n8164 GND.n3707 19.3944
R22152 GND.n8164 GND.n8163 19.3944
R22153 GND.n8163 GND.n8162 19.3944
R22154 GND.n8162 GND.n3713 19.3944
R22155 GND.n8158 GND.n3713 19.3944
R22156 GND.n8158 GND.n8157 19.3944
R22157 GND.n8157 GND.n8156 19.3944
R22158 GND.n8156 GND.n3719 19.3944
R22159 GND.n8152 GND.n3719 19.3944
R22160 GND.n8152 GND.n8151 19.3944
R22161 GND.n8151 GND.n8150 19.3944
R22162 GND.n8150 GND.n3725 19.3944
R22163 GND.n8146 GND.n3725 19.3944
R22164 GND.n8146 GND.n8145 19.3944
R22165 GND.n8145 GND.n8144 19.3944
R22166 GND.n8144 GND.n3731 19.3944
R22167 GND.n8140 GND.n3731 19.3944
R22168 GND.n8140 GND.n8139 19.3944
R22169 GND.n8139 GND.n8138 19.3944
R22170 GND.n8138 GND.n3737 19.3944
R22171 GND.n3741 GND.n3737 19.3944
R22172 GND.n8131 GND.n3741 19.3944
R22173 GND.n8131 GND.n8130 19.3944
R22174 GND.n8130 GND.n8129 19.3944
R22175 GND.n8129 GND.n3747 19.3944
R22176 GND.n8117 GND.n3747 19.3944
R22177 GND.n8117 GND.n8116 19.3944
R22178 GND.n8116 GND.n8115 19.3944
R22179 GND.n8115 GND.n3778 19.3944
R22180 GND.n8103 GND.n3778 19.3944
R22181 GND.n8103 GND.n8102 19.3944
R22182 GND.n8102 GND.n8101 19.3944
R22183 GND.n8101 GND.n3794 19.3944
R22184 GND.n8089 GND.n3794 19.3944
R22185 GND.n8089 GND.n8088 19.3944
R22186 GND.n8088 GND.n8087 19.3944
R22187 GND.n8087 GND.n3812 19.3944
R22188 GND.n8075 GND.n3812 19.3944
R22189 GND.n8075 GND.n8074 19.3944
R22190 GND.n8074 GND.n8073 19.3944
R22191 GND.n8073 GND.n3830 19.3944
R22192 GND.n8061 GND.n3830 19.3944
R22193 GND.n8061 GND.n8060 19.3944
R22194 GND.n8060 GND.n8059 19.3944
R22195 GND.n8059 GND.n3848 19.3944
R22196 GND.n8003 GND.n3848 19.3944
R22197 GND.n8003 GND.n8002 19.3944
R22198 GND.n8002 GND.n8001 19.3944
R22199 GND.n8001 GND.n3891 19.3944
R22200 GND.n7991 GND.n3891 19.3944
R22201 GND.n7991 GND.n7990 19.3944
R22202 GND.n7990 GND.n7989 19.3944
R22203 GND.n7989 GND.n3912 19.3944
R22204 GND.n7979 GND.n3912 19.3944
R22205 GND.n7979 GND.n7978 19.3944
R22206 GND.n7978 GND.n7977 19.3944
R22207 GND.n7977 GND.n3932 19.3944
R22208 GND.n7967 GND.n3932 19.3944
R22209 GND.n7967 GND.n7966 19.3944
R22210 GND.n7966 GND.n7965 19.3944
R22211 GND.n7965 GND.n3952 19.3944
R22212 GND.n7955 GND.n3952 19.3944
R22213 GND.n7955 GND.n7954 19.3944
R22214 GND.n7954 GND.n7953 19.3944
R22215 GND.n7953 GND.n3972 19.3944
R22216 GND.n7943 GND.n3972 19.3944
R22217 GND.n7943 GND.n7942 19.3944
R22218 GND.n7942 GND.n7941 19.3944
R22219 GND.n7941 GND.n3992 19.3944
R22220 GND.n7931 GND.n3992 19.3944
R22221 GND.n7931 GND.n7930 19.3944
R22222 GND.n7930 GND.n7929 19.3944
R22223 GND.n7929 GND.n4012 19.3944
R22224 GND.n7919 GND.n4012 19.3944
R22225 GND.n7919 GND.n7918 19.3944
R22226 GND.n7918 GND.n7917 19.3944
R22227 GND.n7917 GND.n4032 19.3944
R22228 GND.n7907 GND.n4032 19.3944
R22229 GND.n7907 GND.n7906 19.3944
R22230 GND.n7906 GND.n7905 19.3944
R22231 GND.n7905 GND.n4052 19.3944
R22232 GND.n4078 GND.n4052 19.3944
R22233 GND.n7888 GND.n4078 19.3944
R22234 GND.n7888 GND.n7887 19.3944
R22235 GND.n7887 GND.n7886 19.3944
R22236 GND.n7886 GND.n4084 19.3944
R22237 GND.n7876 GND.n4084 19.3944
R22238 GND.n7876 GND.n7875 19.3944
R22239 GND.n7875 GND.n7874 19.3944
R22240 GND.n7874 GND.n4117 19.3944
R22241 GND.n7864 GND.n4117 19.3944
R22242 GND.n7864 GND.n7863 19.3944
R22243 GND.n7863 GND.n7862 19.3944
R22244 GND.n7862 GND.n4137 19.3944
R22245 GND.n7852 GND.n4137 19.3944
R22246 GND.n7852 GND.n7851 19.3944
R22247 GND.n7851 GND.n7850 19.3944
R22248 GND.n7850 GND.n4157 19.3944
R22249 GND.n4183 GND.n4157 19.3944
R22250 GND.n7833 GND.n4183 19.3944
R22251 GND.n7833 GND.n7832 19.3944
R22252 GND.n7832 GND.n7831 19.3944
R22253 GND.n7831 GND.n4189 19.3944
R22254 GND.n7821 GND.n4189 19.3944
R22255 GND.n7821 GND.n7820 19.3944
R22256 GND.n7820 GND.n7819 19.3944
R22257 GND.n7819 GND.n4221 19.3944
R22258 GND.n7809 GND.n4221 19.3944
R22259 GND.n7809 GND.n7808 19.3944
R22260 GND.n7808 GND.n7807 19.3944
R22261 GND.n7807 GND.n4241 19.3944
R22262 GND.n7797 GND.n4241 19.3944
R22263 GND.n7797 GND.n7796 19.3944
R22264 GND.n7796 GND.n7795 19.3944
R22265 GND.n7795 GND.n4259 19.3944
R22266 GND.n4285 GND.n4259 19.3944
R22267 GND.n7778 GND.n4285 19.3944
R22268 GND.n7778 GND.n7777 19.3944
R22269 GND.n7777 GND.n7776 19.3944
R22270 GND.n7776 GND.n4291 19.3944
R22271 GND.n7766 GND.n4291 19.3944
R22272 GND.n7766 GND.n7765 19.3944
R22273 GND.n7765 GND.n7764 19.3944
R22274 GND.n7764 GND.n4324 19.3944
R22275 GND.n7754 GND.n4324 19.3944
R22276 GND.n7754 GND.n7753 19.3944
R22277 GND.n7753 GND.n7752 19.3944
R22278 GND.n7752 GND.n4344 19.3944
R22279 GND.n7742 GND.n4344 19.3944
R22280 GND.n7742 GND.n7741 19.3944
R22281 GND.n7741 GND.n7740 19.3944
R22282 GND.n7740 GND.n4363 19.3944
R22283 GND.n4388 GND.n4363 19.3944
R22284 GND.n7723 GND.n4388 19.3944
R22285 GND.n7723 GND.n7722 19.3944
R22286 GND.n7722 GND.n7721 19.3944
R22287 GND.n7721 GND.n4394 19.3944
R22288 GND.n7709 GND.n4394 19.3944
R22289 GND.n7709 GND.n7708 19.3944
R22290 GND.n7708 GND.n7707 19.3944
R22291 GND.n7707 GND.n4412 19.3944
R22292 GND.n7695 GND.n4412 19.3944
R22293 GND.n7695 GND.n7694 19.3944
R22294 GND.n7694 GND.n7693 19.3944
R22295 GND.n7693 GND.n4430 19.3944
R22296 GND.n7681 GND.n4430 19.3944
R22297 GND.n7681 GND.n7680 19.3944
R22298 GND.n7680 GND.n7679 19.3944
R22299 GND.n7679 GND.n4447 19.3944
R22300 GND.n4519 GND.n4447 19.3944
R22301 GND.n7662 GND.n4519 19.3944
R22302 GND.n7662 GND.n7661 19.3944
R22303 GND.n7661 GND.n7660 19.3944
R22304 GND.n7660 GND.n4525 19.3944
R22305 GND.n7653 GND.n4525 19.3944
R22306 GND.n7653 GND.n7652 19.3944
R22307 GND.n7652 GND.n7651 19.3944
R22308 GND.n7651 GND.n4566 19.3944
R22309 GND.n6541 GND.n4566 19.3944
R22310 GND.n6545 GND.n6541 19.3944
R22311 GND.n6545 GND.n6539 19.3944
R22312 GND.n6549 GND.n6539 19.3944
R22313 GND.n6549 GND.n6537 19.3944
R22314 GND.n6553 GND.n6537 19.3944
R22315 GND.n6553 GND.n6535 19.3944
R22316 GND.n6557 GND.n6535 19.3944
R22317 GND.n6557 GND.n6533 19.3944
R22318 GND.n6730 GND.n6533 19.3944
R22319 GND.n6730 GND.n6729 19.3944
R22320 GND.n6729 GND.n6728 19.3944
R22321 GND.n6728 GND.n6563 19.3944
R22322 GND.n6724 GND.n6563 19.3944
R22323 GND.n6724 GND.n6723 19.3944
R22324 GND.n6723 GND.n6722 19.3944
R22325 GND.n6722 GND.n6569 19.3944
R22326 GND.n6718 GND.n6569 19.3944
R22327 GND.n6718 GND.n6717 19.3944
R22328 GND.n6717 GND.n6716 19.3944
R22329 GND.n6716 GND.n6575 19.3944
R22330 GND.n6712 GND.n6575 19.3944
R22331 GND.n6712 GND.n6711 19.3944
R22332 GND.n6711 GND.n6710 19.3944
R22333 GND.n6710 GND.n6581 19.3944
R22334 GND.n6706 GND.n6581 19.3944
R22335 GND.n6706 GND.n6705 19.3944
R22336 GND.n6705 GND.n6704 19.3944
R22337 GND.n6704 GND.n6587 19.3944
R22338 GND.n6700 GND.n6587 19.3944
R22339 GND.n6700 GND.n6699 19.3944
R22340 GND.n6699 GND.n6698 19.3944
R22341 GND.n6698 GND.n6593 19.3944
R22342 GND.n6694 GND.n6593 19.3944
R22343 GND.n6694 GND.n6693 19.3944
R22344 GND.n6693 GND.n6692 19.3944
R22345 GND.n6692 GND.n6599 19.3944
R22346 GND.n6688 GND.n6599 19.3944
R22347 GND.n6688 GND.n6687 19.3944
R22348 GND.n6687 GND.n6686 19.3944
R22349 GND.n6686 GND.n6605 19.3944
R22350 GND.n6682 GND.n6605 19.3944
R22351 GND.n6682 GND.n6681 19.3944
R22352 GND.n6681 GND.n6680 19.3944
R22353 GND.n6680 GND.n6611 19.3944
R22354 GND.n6676 GND.n6611 19.3944
R22355 GND.n6676 GND.n6675 19.3944
R22356 GND.n6675 GND.n6674 19.3944
R22357 GND.n6674 GND.n6617 19.3944
R22358 GND.n6670 GND.n6617 19.3944
R22359 GND.n6670 GND.n6669 19.3944
R22360 GND.n6669 GND.n6668 19.3944
R22361 GND.n6668 GND.n6623 19.3944
R22362 GND.n6664 GND.n6623 19.3944
R22363 GND.n6664 GND.n6663 19.3944
R22364 GND.n6663 GND.n6662 19.3944
R22365 GND.n6662 GND.n6629 19.3944
R22366 GND.n6658 GND.n6629 19.3944
R22367 GND.n6658 GND.n6657 19.3944
R22368 GND.n6657 GND.n6656 19.3944
R22369 GND.n6656 GND.n6635 19.3944
R22370 GND.n6652 GND.n6635 19.3944
R22371 GND.n6652 GND.n6651 19.3944
R22372 GND.n6651 GND.n6650 19.3944
R22373 GND.n6650 GND.n6642 19.3944
R22374 GND.n6646 GND.n6642 19.3944
R22375 GND.n6646 GND.n6645 19.3944
R22376 GND.n7330 GND.n6262 19.3944
R22377 GND.n7328 GND.n7327 19.3944
R22378 GND.n7324 GND.n7323 19.3944
R22379 GND.n7321 GND.n6265 19.3944
R22380 GND.n7309 GND.n6282 19.3944
R22381 GND.n7309 GND.n7308 19.3944
R22382 GND.n7308 GND.n7307 19.3944
R22383 GND.n7307 GND.n6286 19.3944
R22384 GND.n7303 GND.n6286 19.3944
R22385 GND.n7303 GND.n7302 19.3944
R22386 GND.n7302 GND.n7301 19.3944
R22387 GND.n7301 GND.n6292 19.3944
R22388 GND.n7297 GND.n6292 19.3944
R22389 GND.n7297 GND.n7296 19.3944
R22390 GND.n7296 GND.n7295 19.3944
R22391 GND.n7295 GND.n6298 19.3944
R22392 GND.n7291 GND.n6298 19.3944
R22393 GND.n7291 GND.n7290 19.3944
R22394 GND.n7290 GND.n7289 19.3944
R22395 GND.n7289 GND.n6304 19.3944
R22396 GND.n7285 GND.n6304 19.3944
R22397 GND.n7285 GND.n7284 19.3944
R22398 GND.n7284 GND.n7283 19.3944
R22399 GND.n7283 GND.n6310 19.3944
R22400 GND.n7279 GND.n6310 19.3944
R22401 GND.n7279 GND.n7278 19.3944
R22402 GND.n7278 GND.n7277 19.3944
R22403 GND.n7277 GND.n6316 19.3944
R22404 GND.n7273 GND.n6316 19.3944
R22405 GND.n7273 GND.n7272 19.3944
R22406 GND.n7272 GND.n7271 19.3944
R22407 GND.n7271 GND.n6322 19.3944
R22408 GND.n6431 GND.n6322 19.3944
R22409 GND.n6431 GND.n6430 19.3944
R22410 GND.n6430 GND.n6429 19.3944
R22411 GND.n6429 GND.n6328 19.3944
R22412 GND.n6425 GND.n6328 19.3944
R22413 GND.n6425 GND.n6424 19.3944
R22414 GND.n6424 GND.n6423 19.3944
R22415 GND.n6423 GND.n6334 19.3944
R22416 GND.n6419 GND.n6334 19.3944
R22417 GND.n6419 GND.n6418 19.3944
R22418 GND.n6418 GND.n6417 19.3944
R22419 GND.n6417 GND.n6340 19.3944
R22420 GND.n6413 GND.n6340 19.3944
R22421 GND.n6413 GND.n6412 19.3944
R22422 GND.n6412 GND.n6411 19.3944
R22423 GND.n6411 GND.n6346 19.3944
R22424 GND.n6407 GND.n6346 19.3944
R22425 GND.n6407 GND.n6406 19.3944
R22426 GND.n6406 GND.n6405 19.3944
R22427 GND.n6405 GND.n6352 19.3944
R22428 GND.n6401 GND.n6352 19.3944
R22429 GND.n6401 GND.n6400 19.3944
R22430 GND.n6400 GND.n6399 19.3944
R22431 GND.n6399 GND.n6358 19.3944
R22432 GND.n6395 GND.n6358 19.3944
R22433 GND.n6395 GND.n6394 19.3944
R22434 GND.n6394 GND.n6393 19.3944
R22435 GND.n6393 GND.n6364 19.3944
R22436 GND.n6389 GND.n6364 19.3944
R22437 GND.n6389 GND.n6388 19.3944
R22438 GND.n6388 GND.n6387 19.3944
R22439 GND.n6387 GND.n6370 19.3944
R22440 GND.n6383 GND.n6370 19.3944
R22441 GND.n6383 GND.n6382 19.3944
R22442 GND.n6382 GND.n6381 19.3944
R22443 GND.n6381 GND.n6378 19.3944
R22444 GND.n6378 GND.n464 19.3944
R22445 GND.n10644 GND.n464 19.3944
R22446 GND.n10644 GND.n10643 19.3944
R22447 GND.n10643 GND.n10642 19.3944
R22448 GND.n10642 GND.n468 19.3944
R22449 GND.n10636 GND.n468 19.3944
R22450 GND.n10636 GND.n10635 19.3944
R22451 GND.n10635 GND.n10634 19.3944
R22452 GND.n10634 GND.n476 19.3944
R22453 GND.n10628 GND.n476 19.3944
R22454 GND.n10628 GND.n10627 19.3944
R22455 GND.n10627 GND.n10626 19.3944
R22456 GND.n10626 GND.n484 19.3944
R22457 GND.n10620 GND.n484 19.3944
R22458 GND.n10620 GND.n10619 19.3944
R22459 GND.n10619 GND.n10618 19.3944
R22460 GND.n10618 GND.n492 19.3944
R22461 GND.n10612 GND.n492 19.3944
R22462 GND.n10612 GND.n10611 19.3944
R22463 GND.n10611 GND.n10610 19.3944
R22464 GND.n10610 GND.n500 19.3944
R22465 GND.n10604 GND.n500 19.3944
R22466 GND.n10604 GND.n10603 19.3944
R22467 GND.n10603 GND.n10602 19.3944
R22468 GND.n10602 GND.n508 19.3944
R22469 GND.n10596 GND.n508 19.3944
R22470 GND.n10596 GND.n10595 19.3944
R22471 GND.n10595 GND.n10594 19.3944
R22472 GND.n10594 GND.n516 19.3944
R22473 GND.n10588 GND.n516 19.3944
R22474 GND.n10588 GND.n10587 19.3944
R22475 GND.n10587 GND.n10586 19.3944
R22476 GND.n10586 GND.n524 19.3944
R22477 GND.n10580 GND.n524 19.3944
R22478 GND.n10580 GND.n10579 19.3944
R22479 GND.n10579 GND.n10578 19.3944
R22480 GND.n10578 GND.n532 19.3944
R22481 GND.n10572 GND.n532 19.3944
R22482 GND.n10572 GND.n10571 19.3944
R22483 GND.n10571 GND.n10570 19.3944
R22484 GND.n10570 GND.n540 19.3944
R22485 GND.n10564 GND.n540 19.3944
R22486 GND.n10564 GND.n10563 19.3944
R22487 GND.n10563 GND.n10562 19.3944
R22488 GND.n10562 GND.n548 19.3944
R22489 GND.n10556 GND.n548 19.3944
R22490 GND.n10556 GND.n10555 19.3944
R22491 GND.n10555 GND.n10554 19.3944
R22492 GND.n10554 GND.n556 19.3944
R22493 GND.n10548 GND.n556 19.3944
R22494 GND.n10548 GND.n10547 19.3944
R22495 GND.n10547 GND.n10546 19.3944
R22496 GND.n10546 GND.n564 19.3944
R22497 GND.n10540 GND.n564 19.3944
R22498 GND.n10540 GND.n10539 19.3944
R22499 GND.n10539 GND.n10538 19.3944
R22500 GND.n10538 GND.n572 19.3944
R22501 GND.n9047 GND.n9046 19.3944
R22502 GND.n9046 GND.n1464 19.3944
R22503 GND.n9040 GND.n1464 19.3944
R22504 GND.n9040 GND.n9039 19.3944
R22505 GND.n9039 GND.n9038 19.3944
R22506 GND.n9038 GND.n1472 19.3944
R22507 GND.n9032 GND.n1472 19.3944
R22508 GND.n9032 GND.n9031 19.3944
R22509 GND.n9031 GND.n9030 19.3944
R22510 GND.n9030 GND.n1480 19.3944
R22511 GND.n9024 GND.n1480 19.3944
R22512 GND.n9024 GND.n9023 19.3944
R22513 GND.n9023 GND.n9022 19.3944
R22514 GND.n9022 GND.n1488 19.3944
R22515 GND.n9016 GND.n1488 19.3944
R22516 GND.n9016 GND.n9015 19.3944
R22517 GND.n9015 GND.n9014 19.3944
R22518 GND.n9014 GND.n1496 19.3944
R22519 GND.n9008 GND.n1496 19.3944
R22520 GND.n9008 GND.n9007 19.3944
R22521 GND.n9007 GND.n9006 19.3944
R22522 GND.n9006 GND.n1504 19.3944
R22523 GND.n9000 GND.n1504 19.3944
R22524 GND.n9000 GND.n8999 19.3944
R22525 GND.n8999 GND.n8998 19.3944
R22526 GND.n8998 GND.n1512 19.3944
R22527 GND.n8992 GND.n1512 19.3944
R22528 GND.n8992 GND.n8991 19.3944
R22529 GND.n8991 GND.n8990 19.3944
R22530 GND.n8990 GND.n1520 19.3944
R22531 GND.n8984 GND.n1520 19.3944
R22532 GND.n8984 GND.n8983 19.3944
R22533 GND.n8983 GND.n8982 19.3944
R22534 GND.n8982 GND.n1528 19.3944
R22535 GND.n8976 GND.n1528 19.3944
R22536 GND.n8976 GND.n8975 19.3944
R22537 GND.n8975 GND.n8974 19.3944
R22538 GND.n8974 GND.n1536 19.3944
R22539 GND.n8968 GND.n1536 19.3944
R22540 GND.n8968 GND.n8967 19.3944
R22541 GND.n8967 GND.n8966 19.3944
R22542 GND.n8966 GND.n1544 19.3944
R22543 GND.n8960 GND.n1544 19.3944
R22544 GND.n8960 GND.n8959 19.3944
R22545 GND.n8959 GND.n8958 19.3944
R22546 GND.n8958 GND.n1552 19.3944
R22547 GND.n8952 GND.n1552 19.3944
R22548 GND.n8952 GND.n8951 19.3944
R22549 GND.n8951 GND.n8950 19.3944
R22550 GND.n8950 GND.n1560 19.3944
R22551 GND.n8944 GND.n1560 19.3944
R22552 GND.n8944 GND.n8943 19.3944
R22553 GND.n8943 GND.n8942 19.3944
R22554 GND.n8942 GND.n1568 19.3944
R22555 GND.n8936 GND.n1568 19.3944
R22556 GND.n8936 GND.n8935 19.3944
R22557 GND.n8935 GND.n8934 19.3944
R22558 GND.n8934 GND.n1576 19.3944
R22559 GND.n1853 GND.n1800 19.3944
R22560 GND.n1855 GND.n1853 19.3944
R22561 GND.n1856 GND.n1855 19.3944
R22562 GND.n1856 GND.n1842 19.3944
R22563 GND.n8682 GND.n1842 19.3944
R22564 GND.n8682 GND.n1843 19.3944
R22565 GND.n1863 GND.n1843 19.3944
R22566 GND.n1864 GND.n1863 19.3944
R22567 GND.n1865 GND.n1864 19.3944
R22568 GND.n3173 GND.n1865 19.3944
R22569 GND.n3173 GND.n1871 19.3944
R22570 GND.n1872 GND.n1871 19.3944
R22571 GND.n1873 GND.n1872 19.3944
R22572 GND.n2878 GND.n1873 19.3944
R22573 GND.n2878 GND.n1879 19.3944
R22574 GND.n1880 GND.n1879 19.3944
R22575 GND.n1881 GND.n1880 19.3944
R22576 GND.n2855 GND.n1881 19.3944
R22577 GND.n2855 GND.n1887 19.3944
R22578 GND.n1888 GND.n1887 19.3944
R22579 GND.n1889 GND.n1888 19.3944
R22580 GND.n2842 GND.n1889 19.3944
R22581 GND.n2842 GND.n1895 19.3944
R22582 GND.n1896 GND.n1895 19.3944
R22583 GND.n1897 GND.n1896 19.3944
R22584 GND.n3245 GND.n1897 19.3944
R22585 GND.n3245 GND.n1903 19.3944
R22586 GND.n1904 GND.n1903 19.3944
R22587 GND.n1905 GND.n1904 19.3944
R22588 GND.n3272 GND.n1905 19.3944
R22589 GND.n3272 GND.n1911 19.3944
R22590 GND.n1912 GND.n1911 19.3944
R22591 GND.n1913 GND.n1912 19.3944
R22592 GND.n2787 GND.n1913 19.3944
R22593 GND.n2787 GND.n1919 19.3944
R22594 GND.n1920 GND.n1919 19.3944
R22595 GND.n1921 GND.n1920 19.3944
R22596 GND.n2764 GND.n1921 19.3944
R22597 GND.n2764 GND.n1927 19.3944
R22598 GND.n1928 GND.n1927 19.3944
R22599 GND.n1929 GND.n1928 19.3944
R22600 GND.n2751 GND.n1929 19.3944
R22601 GND.n2751 GND.n1935 19.3944
R22602 GND.n1936 GND.n1935 19.3944
R22603 GND.n1937 GND.n1936 19.3944
R22604 GND.n3344 GND.n1937 19.3944
R22605 GND.n3344 GND.n1943 19.3944
R22606 GND.n1944 GND.n1943 19.3944
R22607 GND.n1945 GND.n1944 19.3944
R22608 GND.n3371 GND.n1945 19.3944
R22609 GND.n3371 GND.n1951 19.3944
R22610 GND.n1952 GND.n1951 19.3944
R22611 GND.n1953 GND.n1952 19.3944
R22612 GND.n2696 GND.n1953 19.3944
R22613 GND.n2696 GND.n1959 19.3944
R22614 GND.n1960 GND.n1959 19.3944
R22615 GND.n1961 GND.n1960 19.3944
R22616 GND.n2673 GND.n1961 19.3944
R22617 GND.n2673 GND.n1967 19.3944
R22618 GND.n1968 GND.n1967 19.3944
R22619 GND.n1969 GND.n1968 19.3944
R22620 GND.n2662 GND.n1969 19.3944
R22621 GND.n2662 GND.n1975 19.3944
R22622 GND.n1976 GND.n1975 19.3944
R22623 GND.n1977 GND.n1976 19.3944
R22624 GND.n2506 GND.n1977 19.3944
R22625 GND.n2506 GND.n1983 19.3944
R22626 GND.n1984 GND.n1983 19.3944
R22627 GND.n1985 GND.n1984 19.3944
R22628 GND.n2529 GND.n1985 19.3944
R22629 GND.n2529 GND.n1991 19.3944
R22630 GND.n1992 GND.n1991 19.3944
R22631 GND.n1993 GND.n1992 19.3944
R22632 GND.n2485 GND.n1993 19.3944
R22633 GND.n2485 GND.n1999 19.3944
R22634 GND.n2000 GND.n1999 19.3944
R22635 GND.n2001 GND.n2000 19.3944
R22636 GND.n3512 GND.n2001 19.3944
R22637 GND.n3512 GND.n2007 19.3944
R22638 GND.n2008 GND.n2007 19.3944
R22639 GND.n2009 GND.n2008 19.3944
R22640 GND.n3540 GND.n2009 19.3944
R22641 GND.n3540 GND.n2015 19.3944
R22642 GND.n2016 GND.n2015 19.3944
R22643 GND.n2017 GND.n2016 19.3944
R22644 GND.n2433 GND.n2017 19.3944
R22645 GND.n2433 GND.n2023 19.3944
R22646 GND.n2024 GND.n2023 19.3944
R22647 GND.n2025 GND.n2024 19.3944
R22648 GND.n2411 GND.n2025 19.3944
R22649 GND.n2411 GND.n2031 19.3944
R22650 GND.n2032 GND.n2031 19.3944
R22651 GND.n2033 GND.n2032 19.3944
R22652 GND.n2398 GND.n2033 19.3944
R22653 GND.n2398 GND.n2039 19.3944
R22654 GND.n2040 GND.n2039 19.3944
R22655 GND.n2041 GND.n2040 19.3944
R22656 GND.n3615 GND.n2041 19.3944
R22657 GND.n3615 GND.n2047 19.3944
R22658 GND.n2048 GND.n2047 19.3944
R22659 GND.n2049 GND.n2048 19.3944
R22660 GND.n3643 GND.n2049 19.3944
R22661 GND.n3643 GND.n2055 19.3944
R22662 GND.n2056 GND.n2055 19.3944
R22663 GND.n2057 GND.n2056 19.3944
R22664 GND.n2349 GND.n2057 19.3944
R22665 GND.n2349 GND.n2063 19.3944
R22666 GND.n2064 GND.n2063 19.3944
R22667 GND.n2065 GND.n2064 19.3944
R22668 GND.n2336 GND.n2065 19.3944
R22669 GND.n2336 GND.n2071 19.3944
R22670 GND.n2072 GND.n2071 19.3944
R22671 GND.n2073 GND.n2072 19.3944
R22672 GND.n2308 GND.n2073 19.3944
R22673 GND.n2308 GND.n2079 19.3944
R22674 GND.n2080 GND.n2079 19.3944
R22675 GND.n2081 GND.n2080 19.3944
R22676 GND.n8204 GND.n2081 19.3944
R22677 GND.n8204 GND.n2087 19.3944
R22678 GND.n2088 GND.n2087 19.3944
R22679 GND.n2089 GND.n2088 19.3944
R22680 GND.n8232 GND.n2089 19.3944
R22681 GND.n8232 GND.n2095 19.3944
R22682 GND.n2096 GND.n2095 19.3944
R22683 GND.n2097 GND.n2096 19.3944
R22684 GND.n2257 GND.n2097 19.3944
R22685 GND.n2257 GND.n2103 19.3944
R22686 GND.n2104 GND.n2103 19.3944
R22687 GND.n2105 GND.n2104 19.3944
R22688 GND.n2235 GND.n2105 19.3944
R22689 GND.n2235 GND.n2111 19.3944
R22690 GND.n2112 GND.n2111 19.3944
R22691 GND.n2113 GND.n2112 19.3944
R22692 GND.n2224 GND.n2113 19.3944
R22693 GND.n2224 GND.n2119 19.3944
R22694 GND.n2120 GND.n2119 19.3944
R22695 GND.n2121 GND.n2120 19.3944
R22696 GND.n8476 GND.n8475 19.3944
R22697 GND.n8473 GND.n8472 19.3944
R22698 GND.n8470 GND.n8469 19.3944
R22699 GND.n8467 GND.n8466 19.3944
R22700 GND.n8464 GND.n8463 19.3944
R22701 GND.n8124 GND.n3767 18.8883
R22702 GND.n4725 GND.n4649 18.8883
R22703 GND.n3760 GND.n3756 18.7329
R22704 GND.n4644 GND.n4643 18.7329
R22705 GND.n5237 GND.n3806 18.7296
R22706 GND.n8071 GND.n8070 18.7296
R22707 GND.n7987 GND.n3914 18.7296
R22708 GND.n5362 GND.n3944 18.7296
R22709 GND.n4978 GND.n3996 18.7296
R22710 GND.n7921 GND.n4026 18.7296
R22711 GND.n4947 GND.n4088 18.7296
R22712 GND.n7866 GND.n4131 18.7296
R22713 GND.n4916 GND.n4915 18.7296
R22714 GND.n7811 GND.n4235 18.7296
R22715 GND.n4882 GND.n4295 18.7296
R22716 GND.n7756 GND.n4338 18.7296
R22717 GND.n7718 GND.n4398 18.7296
R22718 GND.n7697 GND.n4424 18.7296
R22719 GND.n8360 GND.n2185 18.4247
R22720 GND.n7600 GND.n7597 18.4247
R22721 GND.t197 GND.n4086 18.3951
R22722 GND.n5593 GND.t12 18.3951
R22723 GND.n8084 GND.n3816 17.3918
R22724 GND.n8077 GND.n3824 17.3918
R22725 GND.n7981 GND.n3924 17.3918
R22726 GND.n5351 GND.n3934 17.3918
R22727 GND.n4973 GND.n4006 17.3918
R22728 GND.n7927 GND.n4016 17.3918
R22729 GND.n4942 GND.n4111 17.3918
R22730 GND.n7872 GND.n4121 17.3918
R22731 GND.n4910 GND.n4215 17.3918
R22732 GND.n7817 GND.n4225 17.3918
R22733 GND.n4877 GND.n4318 17.3918
R22734 GND.n7762 GND.n4328 17.3918
R22735 GND.n4473 GND.n4406 17.3918
R22736 GND.n7705 GND.n7704 17.3918
R22737 GND.n8698 GND.n1801 16.7229
R22738 GND.n8698 GND.n8697 16.7229
R22739 GND.n8697 GND.n1805 16.7229
R22740 GND.n1816 GND.n1805 16.7229
R22741 GND.n1817 GND.n1816 16.7229
R22742 GND.n8691 GND.n1817 16.7229
R22743 GND.n8691 GND.n8690 16.7229
R22744 GND.n8690 GND.n1820 16.7229
R22745 GND.n2907 GND.n1820 16.7229
R22746 GND.n2907 GND.n1836 16.7229
R22747 GND.n8684 GND.n1836 16.7229
R22748 GND.n8684 GND.n1839 16.7229
R22749 GND.n2964 GND.n1839 16.7229
R22750 GND.n2965 GND.n2964 16.7229
R22751 GND.n3160 GND.n2965 16.7229
R22752 GND.n3152 GND.n3150 16.7229
R22753 GND.n3152 GND.n2901 16.7229
R22754 GND.n3169 GND.n2901 16.7229
R22755 GND.n3169 GND.n2897 16.7229
R22756 GND.n3175 GND.n2897 16.7229
R22757 GND.n3175 GND.n2899 16.7229
R22758 GND.n3171 GND.n2899 16.7229
R22759 GND.n3171 GND.n2886 16.7229
R22760 GND.n3185 GND.n2886 16.7229
R22761 GND.n3185 GND.n2888 16.7229
R22762 GND.n2891 GND.n2888 16.7229
R22763 GND.n2891 GND.n2879 16.7229
R22764 GND.n3194 GND.n2879 16.7229
R22765 GND.n3194 GND.n2874 16.7229
R22766 GND.n3200 GND.n2874 16.7229
R22767 GND.n3200 GND.n2876 16.7229
R22768 GND.n3197 GND.n2876 16.7229
R22769 GND.n3197 GND.n2864 16.7229
R22770 GND.n3210 GND.n2864 16.7229
R22771 GND.n3210 GND.n2865 16.7229
R22772 GND.n2868 GND.n2865 16.7229
R22773 GND.n2868 GND.n2857 16.7229
R22774 GND.n3219 GND.n2857 16.7229
R22775 GND.n3219 GND.n2851 16.7229
R22776 GND.n3224 GND.n2851 16.7229
R22777 GND.n3224 GND.n2854 16.7229
R22778 GND.n3221 GND.n2854 16.7229
R22779 GND.n3221 GND.n2840 16.7229
R22780 GND.n3234 GND.n2840 16.7229
R22781 GND.n3234 GND.n2841 16.7229
R22782 GND.n2845 GND.n2841 16.7229
R22783 GND.n3243 GND.n2832 16.7229
R22784 GND.n3243 GND.n2828 16.7229
R22785 GND.n3249 GND.n2828 16.7229
R22786 GND.n3249 GND.n2830 16.7229
R22787 GND.n3246 GND.n2830 16.7229
R22788 GND.n3246 GND.n2817 16.7229
R22789 GND.n3259 GND.n2817 16.7229
R22790 GND.n3259 GND.n2818 16.7229
R22791 GND.n2822 GND.n2818 16.7229
R22792 GND.n2822 GND.n2810 16.7229
R22793 GND.n3268 GND.n2810 16.7229
R22794 GND.n3268 GND.n2806 16.7229
R22795 GND.n3274 GND.n2806 16.7229
R22796 GND.n3274 GND.n2808 16.7229
R22797 GND.n3270 GND.n2808 16.7229
R22798 GND.n3270 GND.n2795 16.7229
R22799 GND.n3284 GND.n2795 16.7229
R22800 GND.n3284 GND.n2797 16.7229
R22801 GND.n2800 GND.n2797 16.7229
R22802 GND.n2800 GND.n2788 16.7229
R22803 GND.n3293 GND.n2788 16.7229
R22804 GND.n3293 GND.n2783 16.7229
R22805 GND.n3299 GND.n2783 16.7229
R22806 GND.n3299 GND.n2785 16.7229
R22807 GND.n3296 GND.n2785 16.7229
R22808 GND.n3309 GND.n2773 16.7229
R22809 GND.n3309 GND.n2774 16.7229
R22810 GND.n2777 GND.n2774 16.7229
R22811 GND.n2777 GND.n2766 16.7229
R22812 GND.n3318 GND.n2766 16.7229
R22813 GND.n3318 GND.n2760 16.7229
R22814 GND.n3323 GND.n2760 16.7229
R22815 GND.n3323 GND.n2763 16.7229
R22816 GND.n3320 GND.n2763 16.7229
R22817 GND.n3320 GND.n2749 16.7229
R22818 GND.n3333 GND.n2749 16.7229
R22819 GND.n3333 GND.n2750 16.7229
R22820 GND.n2754 GND.n2750 16.7229
R22821 GND.n2754 GND.n2741 16.7229
R22822 GND.n3342 GND.n2741 16.7229
R22823 GND.n3342 GND.n2737 16.7229
R22824 GND.n3348 GND.n2737 16.7229
R22825 GND.n3348 GND.n2739 16.7229
R22826 GND.n3345 GND.n2739 16.7229
R22827 GND.n3345 GND.n2726 16.7229
R22828 GND.n3358 GND.n2726 16.7229
R22829 GND.n3358 GND.n2727 16.7229
R22830 GND.n2731 GND.n2727 16.7229
R22831 GND.n2731 GND.n2719 16.7229
R22832 GND.n3367 GND.n2719 16.7229
R22833 GND.n3373 GND.n2715 16.7229
R22834 GND.n3373 GND.n2717 16.7229
R22835 GND.n3369 GND.n2717 16.7229
R22836 GND.n3369 GND.n2704 16.7229
R22837 GND.n3383 GND.n2704 16.7229
R22838 GND.n3383 GND.n2706 16.7229
R22839 GND.n2709 GND.n2706 16.7229
R22840 GND.n2709 GND.n2697 16.7229
R22841 GND.n3392 GND.n2697 16.7229
R22842 GND.n3392 GND.n2692 16.7229
R22843 GND.n3398 GND.n2692 16.7229
R22844 GND.n3398 GND.n2694 16.7229
R22845 GND.n3395 GND.n2694 16.7229
R22846 GND.n3395 GND.n2682 16.7229
R22847 GND.n3408 GND.n2682 16.7229
R22848 GND.n3408 GND.n2683 16.7229
R22849 GND.n2686 GND.n2683 16.7229
R22850 GND.n2686 GND.n2675 16.7229
R22851 GND.n3417 GND.n2675 16.7229
R22852 GND.n3417 GND.n2669 16.7229
R22853 GND.n3422 GND.n2669 16.7229
R22854 GND.n3422 GND.n2672 16.7229
R22855 GND.n3419 GND.n2672 16.7229
R22856 GND.n3419 GND.n2661 16.7229
R22857 GND.n3430 GND.n2661 16.7229
R22858 GND.n3065 GND.n3064 16.7229
R22859 GND.n3064 GND.n2501 16.7229
R22860 GND.n3490 GND.n2501 16.7229
R22861 GND.n3490 GND.n2504 16.7229
R22862 GND.n3487 GND.n2504 16.7229
R22863 GND.n3487 GND.n3486 16.7229
R22864 GND.n3486 GND.n2509 16.7229
R22865 GND.n2515 GND.n2509 16.7229
R22866 GND.n2516 GND.n2515 16.7229
R22867 GND.n3479 GND.n2516 16.7229
R22868 GND.n3479 GND.n3478 16.7229
R22869 GND.n3478 GND.n2519 16.7229
R22870 GND.n3473 GND.n2519 16.7229
R22871 GND.n3473 GND.n2527 16.7229
R22872 GND.n3470 GND.n2527 16.7229
R22873 GND.n3470 GND.n3469 16.7229
R22874 GND.n3469 GND.n2531 16.7229
R22875 GND.n2649 GND.n2531 16.7229
R22876 GND.n3458 GND.n2649 16.7229
R22877 GND.n3462 GND.n3458 16.7229
R22878 GND.n3462 GND.n3461 16.7229
R22879 GND.n3461 GND.n2483 16.7229
R22880 GND.n3500 GND.n2483 16.7229
R22881 GND.n3500 GND.n2484 16.7229
R22882 GND.n2488 GND.n2476 16.7229
R22883 GND.n3510 GND.n2476 16.7229
R22884 GND.n3510 GND.n2472 16.7229
R22885 GND.n3516 GND.n2472 16.7229
R22886 GND.n3516 GND.n2474 16.7229
R22887 GND.n3513 GND.n2474 16.7229
R22888 GND.n3513 GND.n2461 16.7229
R22889 GND.n3526 GND.n2461 16.7229
R22890 GND.n3526 GND.n2462 16.7229
R22891 GND.n2466 GND.n2462 16.7229
R22892 GND.n2466 GND.n2455 16.7229
R22893 GND.n3536 GND.n2455 16.7229
R22894 GND.n3536 GND.n2451 16.7229
R22895 GND.n3542 GND.n2451 16.7229
R22896 GND.n3542 GND.n2453 16.7229
R22897 GND.n3538 GND.n2453 16.7229
R22898 GND.n3538 GND.n2440 16.7229
R22899 GND.n3552 GND.n2440 16.7229
R22900 GND.n3552 GND.n2442 16.7229
R22901 GND.n2445 GND.n2442 16.7229
R22902 GND.n2445 GND.n2434 16.7229
R22903 GND.n3562 GND.n2434 16.7229
R22904 GND.n3562 GND.n2429 16.7229
R22905 GND.n3568 GND.n2429 16.7229
R22906 GND.n3568 GND.n2431 16.7229
R22907 GND.n3565 GND.n2419 16.7229
R22908 GND.n3578 GND.n2419 16.7229
R22909 GND.n3578 GND.n2420 16.7229
R22910 GND.n2423 GND.n2420 16.7229
R22911 GND.n2423 GND.n2413 16.7229
R22912 GND.n3588 GND.n2413 16.7229
R22913 GND.n3588 GND.n2407 16.7229
R22914 GND.n3593 GND.n2407 16.7229
R22915 GND.n3593 GND.n2410 16.7229
R22916 GND.n3590 GND.n2410 16.7229
R22917 GND.n3590 GND.n2396 16.7229
R22918 GND.n3603 GND.n2396 16.7229
R22919 GND.n3603 GND.n2397 16.7229
R22920 GND.n2401 GND.n2397 16.7229
R22921 GND.n2401 GND.n2389 16.7229
R22922 GND.n3613 GND.n2389 16.7229
R22923 GND.n3613 GND.n2385 16.7229
R22924 GND.n3619 GND.n2385 16.7229
R22925 GND.n3619 GND.n2387 16.7229
R22926 GND.n3616 GND.n2387 16.7229
R22927 GND.n3616 GND.n2376 16.7229
R22928 GND.n3629 GND.n2376 16.7229
R22929 GND.n3629 GND.n2377 16.7229
R22930 GND.n2605 GND.n2377 16.7229
R22931 GND.n2606 GND.n2605 16.7229
R22932 GND.n3639 GND.n2367 16.7229
R22933 GND.n3645 GND.n2367 16.7229
R22934 GND.n3645 GND.n2369 16.7229
R22935 GND.n3641 GND.n2369 16.7229
R22936 GND.n3641 GND.n2356 16.7229
R22937 GND.n3655 GND.n2356 16.7229
R22938 GND.n3655 GND.n2358 16.7229
R22939 GND.n2361 GND.n2358 16.7229
R22940 GND.n2361 GND.n2350 16.7229
R22941 GND.n3665 GND.n2350 16.7229
R22942 GND.n3665 GND.n2345 16.7229
R22943 GND.n3671 GND.n2345 16.7229
R22944 GND.n3671 GND.n2347 16.7229
R22945 GND.n3668 GND.n2347 16.7229
R22946 GND.n3668 GND.n2334 16.7229
R22947 GND.n3681 GND.n2334 16.7229
R22948 GND.n3681 GND.n2335 16.7229
R22949 GND.n2335 GND.n2328 16.7229
R22950 GND.n3692 GND.n2328 16.7229
R22951 GND.n3692 GND.n3691 16.7229
R22952 GND.n3691 GND.n2317 16.7229
R22953 GND.n8182 GND.n2317 16.7229
R22954 GND.n8182 GND.n2320 16.7229
R22955 GND.n8179 GND.n2320 16.7229
R22956 GND.n8179 GND.n8178 16.7229
R22957 GND.n8192 GND.n2307 16.7229
R22958 GND.n2311 GND.n2307 16.7229
R22959 GND.n2311 GND.n2300 16.7229
R22960 GND.n8202 GND.n2300 16.7229
R22961 GND.n8202 GND.n2296 16.7229
R22962 GND.n8208 GND.n2296 16.7229
R22963 GND.n8208 GND.n2298 16.7229
R22964 GND.n8205 GND.n2298 16.7229
R22965 GND.n8205 GND.n2285 16.7229
R22966 GND.n8218 GND.n2285 16.7229
R22967 GND.n8218 GND.n2286 16.7229
R22968 GND.n2290 GND.n2286 16.7229
R22969 GND.n2290 GND.n2279 16.7229
R22970 GND.n8228 GND.n2279 16.7229
R22971 GND.n8228 GND.n2275 16.7229
R22972 GND.n8234 GND.n2275 16.7229
R22973 GND.n8234 GND.n2277 16.7229
R22974 GND.n8230 GND.n2277 16.7229
R22975 GND.n8230 GND.n2264 16.7229
R22976 GND.n8244 GND.n2264 16.7229
R22977 GND.n8244 GND.n2266 16.7229
R22978 GND.n2269 GND.n2266 16.7229
R22979 GND.n2269 GND.n2258 16.7229
R22980 GND.n8254 GND.n2258 16.7229
R22981 GND.n8254 GND.n2253 16.7229
R22982 GND.n8260 GND.n2253 16.7229
R22983 GND.n8260 GND.n2255 16.7229
R22984 GND.n8257 GND.n2255 16.7229
R22985 GND.n8257 GND.n2243 16.7229
R22986 GND.n8270 GND.n2243 16.7229
R22987 GND.n8270 GND.n2244 16.7229
R22988 GND.n2247 GND.n2237 16.7229
R22989 GND.n8280 GND.n2237 16.7229
R22990 GND.n8280 GND.n2231 16.7229
R22991 GND.n8285 GND.n2231 16.7229
R22992 GND.n8285 GND.n2234 16.7229
R22993 GND.n8282 GND.n2234 16.7229
R22994 GND.n8282 GND.n2220 16.7229
R22995 GND.n8294 GND.n2220 16.7229
R22996 GND.n8294 GND.n2221 16.7229
R22997 GND.n2222 GND.n2221 16.7229
R22998 GND.n2222 GND.n2214 16.7229
R22999 GND.n8304 GND.n2214 16.7229
R23000 GND.n8304 GND.n2125 16.7229
R23001 GND.n8480 GND.n2125 16.7229
R23002 GND.n8480 GND.n2128 16.7229
R23003 GND.n7532 GND.n5879 16.7229
R23004 GND.n7532 GND.n5881 16.7229
R23005 GND.n7529 GND.n5881 16.7229
R23006 GND.n7529 GND.n5920 16.7229
R23007 GND.n6745 GND.n5920 16.7229
R23008 GND.n6745 GND.n5929 16.7229
R23009 GND.n7523 GND.n5929 16.7229
R23010 GND.n7523 GND.n5932 16.7229
R23011 GND.n6753 GND.n5932 16.7229
R23012 GND.n6753 GND.n5940 16.7229
R23013 GND.n7517 GND.n5940 16.7229
R23014 GND.n7517 GND.n5943 16.7229
R23015 GND.n6760 GND.n5943 16.7229
R23016 GND.n6760 GND.n5951 16.7229
R23017 GND.n7511 GND.n5951 16.7229
R23018 GND.n6768 GND.n6732 16.7229
R23019 GND.n6768 GND.n5960 16.7229
R23020 GND.n7505 GND.n5960 16.7229
R23021 GND.n7505 GND.n5963 16.7229
R23022 GND.n6775 GND.n5963 16.7229
R23023 GND.n6775 GND.n5971 16.7229
R23024 GND.n7499 GND.n5971 16.7229
R23025 GND.n7499 GND.n5974 16.7229
R23026 GND.n6783 GND.n5974 16.7229
R23027 GND.n6783 GND.n5981 16.7229
R23028 GND.n7493 GND.n5981 16.7229
R23029 GND.n7493 GND.n5984 16.7229
R23030 GND.n6790 GND.n5984 16.7229
R23031 GND.n6790 GND.n5992 16.7229
R23032 GND.n7487 GND.n5992 16.7229
R23033 GND.n7487 GND.n5995 16.7229
R23034 GND.n6798 GND.n5995 16.7229
R23035 GND.n6798 GND.n6002 16.7229
R23036 GND.n7481 GND.n6002 16.7229
R23037 GND.n7481 GND.n6005 16.7229
R23038 GND.n6805 GND.n6005 16.7229
R23039 GND.n6805 GND.n6013 16.7229
R23040 GND.n7475 GND.n6013 16.7229
R23041 GND.n7475 GND.n6016 16.7229
R23042 GND.n6813 GND.n6016 16.7229
R23043 GND.n6813 GND.n6023 16.7229
R23044 GND.n7469 GND.n6023 16.7229
R23045 GND.n7469 GND.n6026 16.7229
R23046 GND.n6820 GND.n6026 16.7229
R23047 GND.n6820 GND.n6034 16.7229
R23048 GND.n7463 GND.n6034 16.7229
R23049 GND.n6828 GND.n6514 16.7229
R23050 GND.n6828 GND.n6043 16.7229
R23051 GND.n7457 GND.n6043 16.7229
R23052 GND.n7457 GND.n6046 16.7229
R23053 GND.n6835 GND.n6046 16.7229
R23054 GND.n6835 GND.n6054 16.7229
R23055 GND.n7451 GND.n6054 16.7229
R23056 GND.n7451 GND.n6057 16.7229
R23057 GND.n6843 GND.n6057 16.7229
R23058 GND.n6843 GND.n6064 16.7229
R23059 GND.n7445 GND.n6064 16.7229
R23060 GND.n7445 GND.n6067 16.7229
R23061 GND.n6850 GND.n6067 16.7229
R23062 GND.n6850 GND.n6075 16.7229
R23063 GND.n7439 GND.n6075 16.7229
R23064 GND.n7439 GND.n6078 16.7229
R23065 GND.n6858 GND.n6078 16.7229
R23066 GND.n6858 GND.n6085 16.7229
R23067 GND.n7433 GND.n6085 16.7229
R23068 GND.n7433 GND.n6088 16.7229
R23069 GND.n6865 GND.n6088 16.7229
R23070 GND.n6865 GND.n6096 16.7229
R23071 GND.n7427 GND.n6096 16.7229
R23072 GND.n7427 GND.n6099 16.7229
R23073 GND.n6873 GND.n6099 16.7229
R23074 GND.n7421 GND.n6106 16.7229
R23075 GND.n7421 GND.n6109 16.7229
R23076 GND.n6880 GND.n6109 16.7229
R23077 GND.n6880 GND.n6117 16.7229
R23078 GND.n7415 GND.n6117 16.7229
R23079 GND.n7415 GND.n6120 16.7229
R23080 GND.n6888 GND.n6120 16.7229
R23081 GND.n6888 GND.n6127 16.7229
R23082 GND.n7409 GND.n6127 16.7229
R23083 GND.n7409 GND.n6130 16.7229
R23084 GND.n6895 GND.n6130 16.7229
R23085 GND.n6895 GND.n6138 16.7229
R23086 GND.n7403 GND.n6138 16.7229
R23087 GND.n7403 GND.n6141 16.7229
R23088 GND.n6903 GND.n6141 16.7229
R23089 GND.n6903 GND.n6148 16.7229
R23090 GND.n7397 GND.n6148 16.7229
R23091 GND.n7397 GND.n6151 16.7229
R23092 GND.n6910 GND.n6151 16.7229
R23093 GND.n6910 GND.n6159 16.7229
R23094 GND.n7391 GND.n6159 16.7229
R23095 GND.n7391 GND.n6162 16.7229
R23096 GND.n6918 GND.n6162 16.7229
R23097 GND.n6918 GND.n6169 16.7229
R23098 GND.n7385 GND.n6169 16.7229
R23099 GND.n6925 GND.n6488 16.7229
R23100 GND.n6925 GND.n6179 16.7229
R23101 GND.n7379 GND.n6179 16.7229
R23102 GND.n7379 GND.n6182 16.7229
R23103 GND.n6933 GND.n6182 16.7229
R23104 GND.n6933 GND.n6189 16.7229
R23105 GND.n7373 GND.n6189 16.7229
R23106 GND.n7373 GND.n6192 16.7229
R23107 GND.n6940 GND.n6192 16.7229
R23108 GND.n6940 GND.n6200 16.7229
R23109 GND.n7367 GND.n6200 16.7229
R23110 GND.n7367 GND.n6203 16.7229
R23111 GND.n6948 GND.n6203 16.7229
R23112 GND.n6948 GND.n6210 16.7229
R23113 GND.n7361 GND.n6210 16.7229
R23114 GND.n7361 GND.n6213 16.7229
R23115 GND.n6955 GND.n6213 16.7229
R23116 GND.n6955 GND.n6221 16.7229
R23117 GND.n7355 GND.n6221 16.7229
R23118 GND.n7355 GND.n6224 16.7229
R23119 GND.n6963 GND.n6224 16.7229
R23120 GND.n6963 GND.n6231 16.7229
R23121 GND.n7349 GND.n6231 16.7229
R23122 GND.n7349 GND.n6234 16.7229
R23123 GND.n6970 GND.n6234 16.7229
R23124 GND.n7343 GND.n6241 16.7229
R23125 GND.n7343 GND.n6244 16.7229
R23126 GND.n6985 GND.n6244 16.7229
R23127 GND.n6985 GND.n6251 16.7229
R23128 GND.n7337 GND.n6251 16.7229
R23129 GND.n7337 GND.n6254 16.7229
R23130 GND.n7333 GND.n6254 16.7229
R23131 GND.n7333 GND.n7332 16.7229
R23132 GND.n7332 GND.n6259 16.7229
R23133 GND.n6471 GND.n6259 16.7229
R23134 GND.n6995 GND.n6471 16.7229
R23135 GND.n6995 GND.n92 16.7229
R23136 GND.n11111 GND.n92 16.7229
R23137 GND.n11111 GND.n94 16.7229
R23138 GND.n7004 GND.n94 16.7229
R23139 GND.n7004 GND.n7003 16.7229
R23140 GND.n7003 GND.n6269 16.7229
R23141 GND.n7319 GND.n6269 16.7229
R23142 GND.n7319 GND.n7318 16.7229
R23143 GND.n7318 GND.n111 16.7229
R23144 GND.n11104 GND.n111 16.7229
R23145 GND.n11104 GND.n114 16.7229
R23146 GND.n7312 GND.n114 16.7229
R23147 GND.n7312 GND.n7311 16.7229
R23148 GND.n11098 GND.n125 16.7229
R23149 GND.n7017 GND.n125 16.7229
R23150 GND.n7017 GND.n132 16.7229
R23151 GND.n11092 GND.n132 16.7229
R23152 GND.n11092 GND.n135 16.7229
R23153 GND.n7025 GND.n135 16.7229
R23154 GND.n7025 GND.n142 16.7229
R23155 GND.n11086 GND.n142 16.7229
R23156 GND.n11086 GND.n145 16.7229
R23157 GND.n7032 GND.n145 16.7229
R23158 GND.n7032 GND.n153 16.7229
R23159 GND.n11080 GND.n153 16.7229
R23160 GND.n11080 GND.n156 16.7229
R23161 GND.n7040 GND.n156 16.7229
R23162 GND.n7040 GND.n163 16.7229
R23163 GND.n11074 GND.n163 16.7229
R23164 GND.n11074 GND.n166 16.7229
R23165 GND.n7047 GND.n166 16.7229
R23166 GND.n7047 GND.n174 16.7229
R23167 GND.n11068 GND.n174 16.7229
R23168 GND.n11068 GND.n177 16.7229
R23169 GND.n7055 GND.n177 16.7229
R23170 GND.n7055 GND.n184 16.7229
R23171 GND.n11062 GND.n184 16.7229
R23172 GND.n11062 GND.n187 16.7229
R23173 GND.n7062 GND.n195 16.7229
R23174 GND.n11056 GND.n195 16.7229
R23175 GND.n11056 GND.n198 16.7229
R23176 GND.n7070 GND.n198 16.7229
R23177 GND.n7070 GND.n205 16.7229
R23178 GND.n11050 GND.n205 16.7229
R23179 GND.n11050 GND.n208 16.7229
R23180 GND.n7077 GND.n208 16.7229
R23181 GND.n7077 GND.n216 16.7229
R23182 GND.n11044 GND.n216 16.7229
R23183 GND.n11044 GND.n219 16.7229
R23184 GND.n7085 GND.n219 16.7229
R23185 GND.n7085 GND.n226 16.7229
R23186 GND.n11038 GND.n226 16.7229
R23187 GND.n11038 GND.n229 16.7229
R23188 GND.n7092 GND.n229 16.7229
R23189 GND.n7092 GND.n237 16.7229
R23190 GND.n11032 GND.n237 16.7229
R23191 GND.n11032 GND.n240 16.7229
R23192 GND.n7101 GND.n240 16.7229
R23193 GND.n7101 GND.n247 16.7229
R23194 GND.n11026 GND.n247 16.7229
R23195 GND.n11026 GND.n250 16.7229
R23196 GND.n7268 GND.n250 16.7229
R23197 GND.n7269 GND.n7268 16.7229
R23198 GND.n11020 GND.n260 16.7229
R23199 GND.n7262 GND.n260 16.7229
R23200 GND.n7262 GND.n267 16.7229
R23201 GND.n11014 GND.n267 16.7229
R23202 GND.n11014 GND.n270 16.7229
R23203 GND.n7256 GND.n270 16.7229
R23204 GND.n7256 GND.n278 16.7229
R23205 GND.n11008 GND.n278 16.7229
R23206 GND.n11008 GND.n281 16.7229
R23207 GND.n7250 GND.n281 16.7229
R23208 GND.n7250 GND.n288 16.7229
R23209 GND.n11002 GND.n288 16.7229
R23210 GND.n11002 GND.n291 16.7229
R23211 GND.n7244 GND.n291 16.7229
R23212 GND.n7244 GND.n299 16.7229
R23213 GND.n10996 GND.n299 16.7229
R23214 GND.n10996 GND.n302 16.7229
R23215 GND.n7238 GND.n302 16.7229
R23216 GND.n7238 GND.n309 16.7229
R23217 GND.n10990 GND.n309 16.7229
R23218 GND.n10990 GND.n312 16.7229
R23219 GND.n7232 GND.n312 16.7229
R23220 GND.n7232 GND.n320 16.7229
R23221 GND.n10984 GND.n320 16.7229
R23222 GND.n10984 GND.n323 16.7229
R23223 GND.n7226 GND.n330 16.7229
R23224 GND.n10978 GND.n330 16.7229
R23225 GND.n10978 GND.n333 16.7229
R23226 GND.n7220 GND.n333 16.7229
R23227 GND.n7220 GND.n341 16.7229
R23228 GND.n10972 GND.n341 16.7229
R23229 GND.n10972 GND.n344 16.7229
R23230 GND.n7214 GND.n344 16.7229
R23231 GND.n7214 GND.n351 16.7229
R23232 GND.n10966 GND.n351 16.7229
R23233 GND.n10966 GND.n354 16.7229
R23234 GND.n7208 GND.n354 16.7229
R23235 GND.n7208 GND.n362 16.7229
R23236 GND.n10960 GND.n362 16.7229
R23237 GND.n10960 GND.n365 16.7229
R23238 GND.n7202 GND.n365 16.7229
R23239 GND.n7202 GND.n372 16.7229
R23240 GND.n10954 GND.n372 16.7229
R23241 GND.n10954 GND.n375 16.7229
R23242 GND.n7196 GND.n375 16.7229
R23243 GND.n7196 GND.n383 16.7229
R23244 GND.n10948 GND.n383 16.7229
R23245 GND.n10948 GND.n386 16.7229
R23246 GND.n7190 GND.n386 16.7229
R23247 GND.n7190 GND.n393 16.7229
R23248 GND.n10942 GND.n393 16.7229
R23249 GND.n10942 GND.n396 16.7229
R23250 GND.n7184 GND.n396 16.7229
R23251 GND.n7184 GND.n404 16.7229
R23252 GND.n10936 GND.n404 16.7229
R23253 GND.n10936 GND.n407 16.7229
R23254 GND.n7178 GND.n414 16.7229
R23255 GND.n10930 GND.n414 16.7229
R23256 GND.n10930 GND.n417 16.7229
R23257 GND.n7172 GND.n417 16.7229
R23258 GND.n7172 GND.n425 16.7229
R23259 GND.n10924 GND.n425 16.7229
R23260 GND.n10924 GND.n428 16.7229
R23261 GND.n7166 GND.n428 16.7229
R23262 GND.n7166 GND.n435 16.7229
R23263 GND.n10918 GND.n435 16.7229
R23264 GND.n10918 GND.n438 16.7229
R23265 GND.n10905 GND.n438 16.7229
R23266 GND.n10905 GND.n445 16.7229
R23267 GND.n10912 GND.n445 16.7229
R23268 GND.n10912 GND.n448 16.7229
R23269 GND.n3065 GND.t159 16.3885
R23270 GND.t175 GND.n2484 16.3885
R23271 GND.t4 GND.n6241 16.3885
R23272 GND.n7311 GND.t17 16.3885
R23273 GND.n8085 GND.n8084 16.054
R23274 GND.n5250 GND.n3824 16.054
R23275 GND.n5343 GND.n3924 16.054
R23276 GND.n7975 GND.n3934 16.054
R23277 GND.n7933 GND.n4006 16.054
R23278 GND.n4968 GND.n4016 16.054
R23279 GND.n7878 GND.n4111 16.054
R23280 GND.n4937 GND.n4121 16.054
R23281 GND.n7823 GND.n4215 16.054
R23282 GND.n4905 GND.n4225 16.054
R23283 GND.n7768 GND.n4318 16.054
R23284 GND.n4872 GND.n4328 16.054
R23285 GND.n7711 GND.n4406 16.054
R23286 GND.n7704 GND.n4416 16.054
R23287 GND.t41 GND.n2715 15.7196
R23288 GND.t25 GND.n2431 15.7196
R23289 GND.n8056 GND.n3861 15.7196
R23290 GND.n7732 GND.n4376 15.7196
R23291 GND.n6488 GND.t157 15.7196
R23292 GND.t38 GND.n187 15.7196
R23293 GND.t0 GND.n2773 15.0507
R23294 GND.n2606 GND.t191 15.0507
R23295 GND.n5412 GND.t35 15.0507
R23296 GND.n5752 GND.t206 15.0507
R23297 GND.t27 GND.n6106 15.0507
R23298 GND.n7269 GND.t29 15.0507
R23299 GND.n8091 GND.n3806 14.7162
R23300 GND.n8070 GND.n3834 14.7162
R23301 GND.n5332 GND.n3914 14.7162
R23302 GND.n7969 GND.n3944 14.7162
R23303 GND.n7939 GND.n3996 14.7162
R23304 GND.n7884 GND.n4088 14.7162
R23305 GND.n4932 GND.n4131 14.7162
R23306 GND.n5631 GND.n4235 14.7162
R23307 GND.n7774 GND.n4295 14.7162
R23308 GND.n5801 GND.n4338 14.7162
R23309 GND.n7719 GND.n7718 14.7162
R23310 GND.n4486 GND.n4424 14.7162
R23311 GND.n2947 GND.n2946 14.546
R23312 GND.n10665 GND.n458 14.546
R23313 GND.n5889 GND.n5888 14.546
R23314 GND.n8461 GND.n8460 14.546
R23315 GND.t171 GND.n2832 14.3818
R23316 GND.n8178 GND.t22 14.3818
R23317 GND.n6514 GND.t2 14.3818
R23318 GND.t20 GND.n323 14.3818
R23319 GND.n5397 GND.t11 14.0473
R23320 GND.n7805 GND.t186 14.0473
R23321 GND.n5079 GND.n3767 13.7371
R23322 GND.n4728 GND.n4649 13.7371
R23323 GND.n8336 GND.n8331 13.3823
R23324 GND.n8412 GND.n8411 13.3823
R23325 GND.n7624 GND.n7623 13.3823
R23326 GND.n7539 GND.n4827 13.3823
R23327 GND.n10788 GND.n10783 13.3823
R23328 GND.n10876 GND.n10875 13.3823
R23329 GND.n8793 GND.n8792 13.3823
R23330 GND.n8706 GND.n1793 13.3823
R23331 GND.n8099 GND.n8098 13.3784
R23332 GND.n5035 GND.n3842 13.3784
R23333 GND.n5324 GND.n5323 13.3784
R23334 GND.n7963 GND.n3954 13.3784
R23335 GND.n7945 GND.n3986 13.3784
R23336 GND.n5504 GND.n4036 13.3784
R23337 GND.n7890 GND.n4074 13.3784
R23338 GND.n5607 GND.n4141 13.3784
R23339 GND.n7835 GND.n4179 13.3784
R23340 GND.n5710 GND.n4893 13.3784
R23341 GND.n7780 GND.n4281 13.3784
R23342 GND.n5794 GND.n5793 13.3784
R23343 GND.n7725 GND.n4384 13.3784
R23344 GND.n7690 GND.n4434 13.3784
R23345 GND.n7664 GND.n4516 13.3784
R23346 GND.n3766 GND.n3754 13.1884
R23347 GND.n4639 GND.n4638 13.1049
R23348 GND.n5490 GND.t208 13.044
R23349 GND.t8 GND.n4191 13.044
R23350 GND.n4722 GND.t108 12.7095
R23351 GND.n8336 GND.n2196 12.6066
R23352 GND.n8413 GND.n8412 12.6066
R23353 GND.n7623 GND.n7622 12.6066
R23354 GND.n7542 GND.n7539 12.6066
R23355 GND.n10791 GND.n10788 12.6066
R23356 GND.n10875 GND.n10731 12.6066
R23357 GND.n8792 GND.n8791 12.6066
R23358 GND.n8709 GND.n8706 12.6066
R23359 GND.n4648 GND.n4637 12.4126
R23360 GND.n8113 GND.n3780 12.0406
R23361 GND.n8105 GND.n3788 12.0406
R23362 GND.n3881 GND.n3861 12.0406
R23363 GND.n5024 GND.n3893 12.0406
R23364 GND.n7957 GND.n3964 12.0406
R23365 GND.n7951 GND.n3976 12.0406
R23366 GND.n4953 GND.n4046 12.0406
R23367 GND.n7897 GND.n4064 12.0406
R23368 GND.n4922 GND.n4151 12.0406
R23369 GND.n7842 GND.n4169 12.0406
R23370 GND.n4888 GND.n4253 12.0406
R23371 GND.n7787 GND.n4271 12.0406
R23372 GND.n5809 GND.n4357 12.0406
R23373 GND.n7732 GND.n4375 12.0406
R23374 GND.n4498 GND.n4497 12.0406
R23375 GND.n2949 GND.n2947 11.4429
R23376 GND.n10899 GND.n458 11.4429
R23377 GND.n5211 GND.t90 11.3717
R23378 GND.n7993 GND.t114 11.0373
R23379 GND.n7750 GND.t146 11.0373
R23380 GND.t150 GND.n8119 10.7028
R23381 GND.n8113 GND.n8112 10.7028
R23382 GND.n8106 GND.n8105 10.7028
R23383 GND.n3882 GND.n3881 10.7028
R23384 GND.n5024 GND.n3884 10.7028
R23385 GND.n7957 GND.n3966 10.7028
R23386 GND.n7951 GND.n3974 10.7028
R23387 GND.n4953 GND.n4054 10.7028
R23388 GND.n4064 GND.n4057 10.7028
R23389 GND.n4922 GND.n4159 10.7028
R23390 GND.n4169 GND.n4162 10.7028
R23391 GND.n4888 GND.n4261 10.7028
R23392 GND.n4271 GND.n4264 10.7028
R23393 GND.n5809 GND.n4365 10.7028
R23394 GND.n4375 GND.n4368 10.7028
R23395 GND.n4497 GND.n4449 10.7028
R23396 GND.n4504 GND.n4451 10.7028
R23397 GND.n7 GND.t221 10.6171
R23398 GND.n7 GND.t211 10.6171
R23399 GND.n9 GND.t227 10.6171
R23400 GND.n9 GND.t176 10.6171
R23401 GND.n11 GND.t24 10.6171
R23402 GND.n11 GND.t166 10.6171
R23403 GND.n14 GND.t215 10.6171
R23404 GND.n14 GND.t192 10.6171
R23405 GND.n16 GND.t201 10.6171
R23406 GND.n16 GND.t181 10.6171
R23407 GND.n18 GND.t37 10.6171
R23408 GND.n18 GND.t174 10.6171
R23409 GND.n22 GND.t229 10.6171
R23410 GND.n22 GND.t212 10.6171
R23411 GND.n24 GND.t160 10.6171
R23412 GND.n24 GND.t177 10.6171
R23413 GND.n26 GND.t1 10.6171
R23414 GND.n26 GND.t167 10.6171
R23415 GND.n30 GND.t26 10.6171
R23416 GND.n30 GND.t226 10.6171
R23417 GND.n32 GND.t162 10.6171
R23418 GND.n32 GND.t187 10.6171
R23419 GND.n34 GND.t190 10.6171
R23420 GND.n34 GND.t42 10.6171
R23421 GND.n0 GND.t31 10.6171
R23422 GND.n0 GND.t196 10.6171
R23423 GND.n2 GND.t179 10.6171
R23424 GND.n2 GND.t195 10.6171
R23425 GND.n4 GND.t178 10.6171
R23426 GND.n4 GND.t165 10.6171
R23427 GND.n51 GND.t39 10.6171
R23428 GND.n51 GND.t43 10.6171
R23429 GND.n49 GND.t222 10.6171
R23430 GND.n49 GND.t228 10.6171
R23431 GND.n47 GND.t230 10.6171
R23432 GND.n47 GND.t203 10.6171
R23433 GND.n58 GND.t232 10.6171
R23434 GND.n58 GND.t188 10.6171
R23435 GND.n56 GND.t182 10.6171
R23436 GND.n56 GND.t220 10.6171
R23437 GND.n54 GND.t28 10.6171
R23438 GND.n54 GND.t158 10.6171
R23439 GND.n66 GND.t40 10.6171
R23440 GND.n66 GND.t183 10.6171
R23441 GND.n64 GND.t223 10.6171
R23442 GND.n64 GND.t164 10.6171
R23443 GND.n62 GND.t170 10.6171
R23444 GND.n62 GND.t204 10.6171
R23445 GND.n74 GND.t189 10.6171
R23446 GND.n74 GND.t218 10.6171
R23447 GND.n72 GND.t19 10.6171
R23448 GND.n72 GND.t18 10.6171
R23449 GND.n70 GND.t216 10.6171
R23450 GND.n70 GND.t193 10.6171
R23451 GND.n82 GND.t233 10.6171
R23452 GND.n82 GND.t30 10.6171
R23453 GND.n80 GND.t5 10.6171
R23454 GND.n80 GND.t185 10.6171
R23455 GND.n78 GND.t217 10.6171
R23456 GND.n78 GND.t224 10.6171
R23457 GND.n4659 GND.n4634 10.6151
R23458 GND.n4660 GND.n4659 10.6151
R23459 GND.n4663 GND.n4660 10.6151
R23460 GND.n4668 GND.n4665 10.6151
R23461 GND.n4669 GND.n4668 10.6151
R23462 GND.n4672 GND.n4669 10.6151
R23463 GND.n4673 GND.n4672 10.6151
R23464 GND.n4676 GND.n4673 10.6151
R23465 GND.n4677 GND.n4676 10.6151
R23466 GND.n4680 GND.n4677 10.6151
R23467 GND.n4681 GND.n4680 10.6151
R23468 GND.n4684 GND.n4681 10.6151
R23469 GND.n4685 GND.n4684 10.6151
R23470 GND.n4688 GND.n4685 10.6151
R23471 GND.n4689 GND.n4688 10.6151
R23472 GND.n4692 GND.n4689 10.6151
R23473 GND.n4693 GND.n4692 10.6151
R23474 GND.n4696 GND.n4693 10.6151
R23475 GND.n4697 GND.n4696 10.6151
R23476 GND.n4700 GND.n4697 10.6151
R23477 GND.n4701 GND.n4700 10.6151
R23478 GND.n4704 GND.n4701 10.6151
R23479 GND.n4705 GND.n4704 10.6151
R23480 GND.n4708 GND.n4705 10.6151
R23481 GND.n4709 GND.n4708 10.6151
R23482 GND.n4712 GND.n4709 10.6151
R23483 GND.n4713 GND.n4712 10.6151
R23484 GND.n4716 GND.n4713 10.6151
R23485 GND.n4718 GND.n4716 10.6151
R23486 GND.n5207 GND.n5205 10.6151
R23487 GND.n5208 GND.n5207 10.6151
R23488 GND.n5209 GND.n5208 10.6151
R23489 GND.n5209 GND.n5041 10.6151
R23490 GND.n5217 GND.n5041 10.6151
R23491 GND.n5218 GND.n5217 10.6151
R23492 GND.n5220 GND.n5218 10.6151
R23493 GND.n5221 GND.n5220 10.6151
R23494 GND.n5222 GND.n5221 10.6151
R23495 GND.n5222 GND.n5040 10.6151
R23496 GND.n5230 GND.n5040 10.6151
R23497 GND.n5231 GND.n5230 10.6151
R23498 GND.n5233 GND.n5231 10.6151
R23499 GND.n5234 GND.n5233 10.6151
R23500 GND.n5235 GND.n5234 10.6151
R23501 GND.n5235 GND.n5039 10.6151
R23502 GND.n5243 GND.n5039 10.6151
R23503 GND.n5244 GND.n5243 10.6151
R23504 GND.n5246 GND.n5244 10.6151
R23505 GND.n5247 GND.n5246 10.6151
R23506 GND.n5248 GND.n5247 10.6151
R23507 GND.n5248 GND.n5038 10.6151
R23508 GND.n5256 GND.n5038 10.6151
R23509 GND.n5257 GND.n5256 10.6151
R23510 GND.n5259 GND.n5257 10.6151
R23511 GND.n5260 GND.n5259 10.6151
R23512 GND.n5261 GND.n5260 10.6151
R23513 GND.n5303 GND.n5261 10.6151
R23514 GND.n5303 GND.n5302 10.6151
R23515 GND.n5302 GND.n5301 10.6151
R23516 GND.n5301 GND.n5298 10.6151
R23517 GND.n5298 GND.n5297 10.6151
R23518 GND.n5297 GND.n5296 10.6151
R23519 GND.n5296 GND.n5262 10.6151
R23520 GND.n5292 GND.n5262 10.6151
R23521 GND.n5292 GND.n5291 10.6151
R23522 GND.n5291 GND.n5290 10.6151
R23523 GND.n5290 GND.n5289 10.6151
R23524 GND.n5289 GND.n5287 10.6151
R23525 GND.n5287 GND.n5286 10.6151
R23526 GND.n5286 GND.n5283 10.6151
R23527 GND.n5283 GND.n5282 10.6151
R23528 GND.n5282 GND.n5281 10.6151
R23529 GND.n5281 GND.n5278 10.6151
R23530 GND.n5278 GND.n5277 10.6151
R23531 GND.n5277 GND.n5276 10.6151
R23532 GND.n5276 GND.n5273 10.6151
R23533 GND.n5273 GND.n5272 10.6151
R23534 GND.n5272 GND.n5271 10.6151
R23535 GND.n5271 GND.n5268 10.6151
R23536 GND.n5268 GND.n5267 10.6151
R23537 GND.n5267 GND.n5266 10.6151
R23538 GND.n5266 GND.n5264 10.6151
R23539 GND.n5264 GND.n4995 10.6151
R23540 GND.n5424 GND.n4995 10.6151
R23541 GND.n5425 GND.n5424 10.6151
R23542 GND.n5428 GND.n5425 10.6151
R23543 GND.n5428 GND.n5427 10.6151
R23544 GND.n5427 GND.n5426 10.6151
R23545 GND.n5426 GND.n4985 10.6151
R23546 GND.n5442 GND.n4985 10.6151
R23547 GND.n5443 GND.n5442 10.6151
R23548 GND.n5446 GND.n5443 10.6151
R23549 GND.n5446 GND.n5445 10.6151
R23550 GND.n5445 GND.n5444 10.6151
R23551 GND.n5444 GND.n4976 10.6151
R23552 GND.n5460 GND.n4976 10.6151
R23553 GND.n5461 GND.n5460 10.6151
R23554 GND.n5464 GND.n5461 10.6151
R23555 GND.n5464 GND.n5463 10.6151
R23556 GND.n5463 GND.n5462 10.6151
R23557 GND.n5462 GND.n4966 10.6151
R23558 GND.n5478 GND.n4966 10.6151
R23559 GND.n5479 GND.n5478 10.6151
R23560 GND.n5488 GND.n5479 10.6151
R23561 GND.n5488 GND.n5487 10.6151
R23562 GND.n5487 GND.n5486 10.6151
R23563 GND.n5486 GND.n5484 10.6151
R23564 GND.n5484 GND.n5483 10.6151
R23565 GND.n5483 GND.n5480 10.6151
R23566 GND.n5480 GND.n4061 10.6151
R23567 GND.n7901 GND.n4061 10.6151
R23568 GND.n7901 GND.n7900 10.6151
R23569 GND.n7900 GND.n7899 10.6151
R23570 GND.n7899 GND.n4062 10.6151
R23571 GND.n5545 GND.n4062 10.6151
R23572 GND.n5546 GND.n5545 10.6151
R23573 GND.n5549 GND.n5546 10.6151
R23574 GND.n5549 GND.n5548 10.6151
R23575 GND.n5548 GND.n5547 10.6151
R23576 GND.n5547 GND.n4945 10.6151
R23577 GND.n5563 GND.n4945 10.6151
R23578 GND.n5564 GND.n5563 10.6151
R23579 GND.n5567 GND.n5564 10.6151
R23580 GND.n5567 GND.n5566 10.6151
R23581 GND.n5566 GND.n5565 10.6151
R23582 GND.n5565 GND.n4935 10.6151
R23583 GND.n5581 GND.n4935 10.6151
R23584 GND.n5582 GND.n5581 10.6151
R23585 GND.n5591 GND.n5582 10.6151
R23586 GND.n5591 GND.n5590 10.6151
R23587 GND.n5590 GND.n5589 10.6151
R23588 GND.n5589 GND.n5587 10.6151
R23589 GND.n5587 GND.n5586 10.6151
R23590 GND.n5586 GND.n5583 10.6151
R23591 GND.n5583 GND.n4166 10.6151
R23592 GND.n7846 GND.n4166 10.6151
R23593 GND.n7846 GND.n7845 10.6151
R23594 GND.n7845 GND.n7844 10.6151
R23595 GND.n7844 GND.n4167 10.6151
R23596 GND.n5649 GND.n4167 10.6151
R23597 GND.n5650 GND.n5649 10.6151
R23598 GND.n5653 GND.n5650 10.6151
R23599 GND.n5653 GND.n5652 10.6151
R23600 GND.n5652 GND.n5651 10.6151
R23601 GND.n5651 GND.n4913 10.6151
R23602 GND.n5667 GND.n4913 10.6151
R23603 GND.n5668 GND.n5667 10.6151
R23604 GND.n5671 GND.n5668 10.6151
R23605 GND.n5671 GND.n5670 10.6151
R23606 GND.n5670 GND.n5669 10.6151
R23607 GND.n5669 GND.n4904 10.6151
R23608 GND.n4904 GND.n4902 10.6151
R23609 GND.n5687 GND.n4902 10.6151
R23610 GND.n5688 GND.n5687 10.6151
R23611 GND.n5695 GND.n5688 10.6151
R23612 GND.n5695 GND.n5694 10.6151
R23613 GND.n5694 GND.n5693 10.6151
R23614 GND.n5693 GND.n5692 10.6151
R23615 GND.n5692 GND.n5689 10.6151
R23616 GND.n5689 GND.n4268 10.6151
R23617 GND.n7791 GND.n4268 10.6151
R23618 GND.n7791 GND.n7790 10.6151
R23619 GND.n7790 GND.n7789 10.6151
R23620 GND.n7789 GND.n4269 10.6151
R23621 GND.n5746 GND.n4269 10.6151
R23622 GND.n5747 GND.n5746 10.6151
R23623 GND.n5750 GND.n5747 10.6151
R23624 GND.n5750 GND.n5749 10.6151
R23625 GND.n5749 GND.n5748 10.6151
R23626 GND.n5748 GND.n4880 10.6151
R23627 GND.n5764 GND.n4880 10.6151
R23628 GND.n5765 GND.n5764 10.6151
R23629 GND.n5768 GND.n5765 10.6151
R23630 GND.n5768 GND.n5767 10.6151
R23631 GND.n5767 GND.n5766 10.6151
R23632 GND.n5766 GND.n4871 10.6151
R23633 GND.n4871 GND.n4869 10.6151
R23634 GND.n5782 GND.n4869 10.6151
R23635 GND.n5783 GND.n5782 10.6151
R23636 GND.n5785 GND.n5783 10.6151
R23637 GND.n5786 GND.n5785 10.6151
R23638 GND.n5790 GND.n5786 10.6151
R23639 GND.n5790 GND.n5789 10.6151
R23640 GND.n5789 GND.n5788 10.6151
R23641 GND.n5788 GND.n4372 10.6151
R23642 GND.n7736 GND.n4372 10.6151
R23643 GND.n7736 GND.n7735 10.6151
R23644 GND.n7735 GND.n7734 10.6151
R23645 GND.n7734 GND.n4373 10.6151
R23646 GND.n4457 GND.n4373 10.6151
R23647 GND.n4458 GND.n4457 10.6151
R23648 GND.n4458 GND.n4456 10.6151
R23649 GND.n4466 GND.n4456 10.6151
R23650 GND.n4467 GND.n4466 10.6151
R23651 GND.n4469 GND.n4467 10.6151
R23652 GND.n4470 GND.n4469 10.6151
R23653 GND.n4471 GND.n4470 10.6151
R23654 GND.n4471 GND.n4455 10.6151
R23655 GND.n4479 GND.n4455 10.6151
R23656 GND.n4480 GND.n4479 10.6151
R23657 GND.n4482 GND.n4480 10.6151
R23658 GND.n4483 GND.n4482 10.6151
R23659 GND.n4484 GND.n4483 10.6151
R23660 GND.n4484 GND.n4454 10.6151
R23661 GND.n4492 GND.n4454 10.6151
R23662 GND.n4493 GND.n4492 10.6151
R23663 GND.n4495 GND.n4493 10.6151
R23664 GND.n4496 GND.n4495 10.6151
R23665 GND.n4500 GND.n4496 10.6151
R23666 GND.n4501 GND.n4500 10.6151
R23667 GND.n7675 GND.n4501 10.6151
R23668 GND.n7675 GND.n7674 10.6151
R23669 GND.n7674 GND.n7673 10.6151
R23670 GND.n7673 GND.n4502 10.6151
R23671 GND.n4653 GND.n4502 10.6151
R23672 GND.n4654 GND.n4653 10.6151
R23673 GND.n4720 GND.n4654 10.6151
R23674 GND.n4720 GND.n4719 10.6151
R23675 GND.n5142 GND.n5058 10.6151
R23676 GND.n5148 GND.n5058 10.6151
R23677 GND.n5149 GND.n5148 10.6151
R23678 GND.n5151 GND.n5054 10.6151
R23679 GND.n5157 GND.n5054 10.6151
R23680 GND.n5158 GND.n5157 10.6151
R23681 GND.n5159 GND.n5158 10.6151
R23682 GND.n5159 GND.n5052 10.6151
R23683 GND.n5165 GND.n5052 10.6151
R23684 GND.n5166 GND.n5165 10.6151
R23685 GND.n5167 GND.n5166 10.6151
R23686 GND.n5167 GND.n5050 10.6151
R23687 GND.n5173 GND.n5050 10.6151
R23688 GND.n5174 GND.n5173 10.6151
R23689 GND.n5175 GND.n5174 10.6151
R23690 GND.n5175 GND.n5048 10.6151
R23691 GND.n5181 GND.n5048 10.6151
R23692 GND.n5182 GND.n5181 10.6151
R23693 GND.n5183 GND.n5182 10.6151
R23694 GND.n5183 GND.n5046 10.6151
R23695 GND.n5189 GND.n5046 10.6151
R23696 GND.n5190 GND.n5189 10.6151
R23697 GND.n5191 GND.n5190 10.6151
R23698 GND.n5191 GND.n5044 10.6151
R23699 GND.n5197 GND.n5044 10.6151
R23700 GND.n5198 GND.n5197 10.6151
R23701 GND.n5199 GND.n5198 10.6151
R23702 GND.n5199 GND.n5042 10.6151
R23703 GND.n5204 GND.n5042 10.6151
R23704 GND.n5082 GND.n5079 10.6151
R23705 GND.n5083 GND.n5082 10.6151
R23706 GND.n5084 GND.n5083 10.6151
R23707 GND.n5084 GND.n5077 10.6151
R23708 GND.n5090 GND.n5077 10.6151
R23709 GND.n5091 GND.n5090 10.6151
R23710 GND.n5092 GND.n5091 10.6151
R23711 GND.n5092 GND.n5075 10.6151
R23712 GND.n5098 GND.n5075 10.6151
R23713 GND.n5099 GND.n5098 10.6151
R23714 GND.n5100 GND.n5099 10.6151
R23715 GND.n5100 GND.n5073 10.6151
R23716 GND.n5106 GND.n5073 10.6151
R23717 GND.n5107 GND.n5106 10.6151
R23718 GND.n5108 GND.n5107 10.6151
R23719 GND.n5108 GND.n5071 10.6151
R23720 GND.n5114 GND.n5071 10.6151
R23721 GND.n5115 GND.n5114 10.6151
R23722 GND.n5116 GND.n5115 10.6151
R23723 GND.n5116 GND.n5069 10.6151
R23724 GND.n5122 GND.n5069 10.6151
R23725 GND.n5123 GND.n5122 10.6151
R23726 GND.n5124 GND.n5123 10.6151
R23727 GND.n5124 GND.n5067 10.6151
R23728 GND.n5130 GND.n5067 10.6151
R23729 GND.n5131 GND.n5130 10.6151
R23730 GND.n5133 GND.n5063 10.6151
R23731 GND.n5063 GND.n5062 10.6151
R23732 GND.n5140 GND.n5062 10.6151
R23733 GND.n4729 GND.n4728 10.6151
R23734 GND.n4732 GND.n4729 10.6151
R23735 GND.n4733 GND.n4732 10.6151
R23736 GND.n4736 GND.n4733 10.6151
R23737 GND.n4737 GND.n4736 10.6151
R23738 GND.n4740 GND.n4737 10.6151
R23739 GND.n4741 GND.n4740 10.6151
R23740 GND.n4744 GND.n4741 10.6151
R23741 GND.n4745 GND.n4744 10.6151
R23742 GND.n4748 GND.n4745 10.6151
R23743 GND.n4749 GND.n4748 10.6151
R23744 GND.n4752 GND.n4749 10.6151
R23745 GND.n4753 GND.n4752 10.6151
R23746 GND.n4756 GND.n4753 10.6151
R23747 GND.n4757 GND.n4756 10.6151
R23748 GND.n4760 GND.n4757 10.6151
R23749 GND.n4761 GND.n4760 10.6151
R23750 GND.n4764 GND.n4761 10.6151
R23751 GND.n4765 GND.n4764 10.6151
R23752 GND.n4768 GND.n4765 10.6151
R23753 GND.n4769 GND.n4768 10.6151
R23754 GND.n4772 GND.n4769 10.6151
R23755 GND.n4773 GND.n4772 10.6151
R23756 GND.n4776 GND.n4773 10.6151
R23757 GND.n4777 GND.n4776 10.6151
R23758 GND.n4780 GND.n4777 10.6151
R23759 GND.n4785 GND.n4782 10.6151
R23760 GND.n4786 GND.n4785 10.6151
R23761 GND.n4789 GND.n4786 10.6151
R23762 GND.n8124 GND.n8123 10.6151
R23763 GND.n8123 GND.n8122 10.6151
R23764 GND.n8122 GND.n3768 10.6151
R23765 GND.n5212 GND.n3768 10.6151
R23766 GND.n5212 GND.n3784 10.6151
R23767 GND.n8110 GND.n3784 10.6151
R23768 GND.n8110 GND.n8109 10.6151
R23769 GND.n8109 GND.n8108 10.6151
R23770 GND.n8108 GND.n3785 10.6151
R23771 GND.n5225 GND.n3785 10.6151
R23772 GND.n5225 GND.n3801 10.6151
R23773 GND.n8096 GND.n3801 10.6151
R23774 GND.n8096 GND.n8095 10.6151
R23775 GND.n8095 GND.n8094 10.6151
R23776 GND.n8094 GND.n3802 10.6151
R23777 GND.n5238 GND.n3802 10.6151
R23778 GND.n5238 GND.n3819 10.6151
R23779 GND.n8082 GND.n3819 10.6151
R23780 GND.n8082 GND.n8081 10.6151
R23781 GND.n8081 GND.n8080 10.6151
R23782 GND.n8080 GND.n3820 10.6151
R23783 GND.n5251 GND.n3820 10.6151
R23784 GND.n5251 GND.n3837 10.6151
R23785 GND.n8068 GND.n3837 10.6151
R23786 GND.n8068 GND.n8067 10.6151
R23787 GND.n8067 GND.n8066 10.6151
R23788 GND.n8066 GND.n3838 10.6151
R23789 GND.n5307 GND.n3838 10.6151
R23790 GND.n5308 GND.n5307 10.6151
R23791 GND.n5308 GND.n5034 10.6151
R23792 GND.n5312 GND.n5034 10.6151
R23793 GND.n5313 GND.n5312 10.6151
R23794 GND.n5314 GND.n5313 10.6151
R23795 GND.n5314 GND.n5033 10.6151
R23796 GND.n5318 GND.n5033 10.6151
R23797 GND.n5319 GND.n5318 10.6151
R23798 GND.n5321 GND.n5319 10.6151
R23799 GND.n5321 GND.n5320 10.6151
R23800 GND.n5320 GND.n5018 10.6151
R23801 GND.n5336 GND.n5018 10.6151
R23802 GND.n5337 GND.n5336 10.6151
R23803 GND.n5340 GND.n5337 10.6151
R23804 GND.n5340 GND.n5339 10.6151
R23805 GND.n5339 GND.n5338 10.6151
R23806 GND.n5338 GND.n5009 10.6151
R23807 GND.n5355 GND.n5009 10.6151
R23808 GND.n5356 GND.n5355 10.6151
R23809 GND.n5359 GND.n5356 10.6151
R23810 GND.n5359 GND.n5358 10.6151
R23811 GND.n5358 GND.n5357 10.6151
R23812 GND.n5357 GND.n5000 10.6151
R23813 GND.n5415 GND.n5000 10.6151
R23814 GND.n5416 GND.n5415 10.6151
R23815 GND.n5419 GND.n5416 10.6151
R23816 GND.n5419 GND.n5418 10.6151
R23817 GND.n5418 GND.n5417 10.6151
R23818 GND.n5417 GND.n4990 10.6151
R23819 GND.n5433 GND.n4990 10.6151
R23820 GND.n5434 GND.n5433 10.6151
R23821 GND.n5437 GND.n5434 10.6151
R23822 GND.n5437 GND.n5436 10.6151
R23823 GND.n5436 GND.n5435 10.6151
R23824 GND.n5435 GND.n4981 10.6151
R23825 GND.n5451 GND.n4981 10.6151
R23826 GND.n5452 GND.n5451 10.6151
R23827 GND.n5455 GND.n5452 10.6151
R23828 GND.n5455 GND.n5454 10.6151
R23829 GND.n5454 GND.n5453 10.6151
R23830 GND.n5453 GND.n4971 10.6151
R23831 GND.n5469 GND.n4971 10.6151
R23832 GND.n5470 GND.n5469 10.6151
R23833 GND.n5473 GND.n5470 10.6151
R23834 GND.n5473 GND.n5472 10.6151
R23835 GND.n5472 GND.n5471 10.6151
R23836 GND.n5471 GND.n4961 10.6151
R23837 GND.n5493 GND.n4961 10.6151
R23838 GND.n5494 GND.n5493 10.6151
R23839 GND.n5501 GND.n5494 10.6151
R23840 GND.n5501 GND.n5500 10.6151
R23841 GND.n5500 GND.n5499 10.6151
R23842 GND.n5499 GND.n5496 10.6151
R23843 GND.n5496 GND.n5495 10.6151
R23844 GND.n5495 GND.n4068 10.6151
R23845 GND.n7895 GND.n4068 10.6151
R23846 GND.n7895 GND.n7894 10.6151
R23847 GND.n7894 GND.n7893 10.6151
R23848 GND.n7893 GND.n4069 10.6151
R23849 GND.n4950 GND.n4069 10.6151
R23850 GND.n5554 GND.n4950 10.6151
R23851 GND.n5555 GND.n5554 10.6151
R23852 GND.n5558 GND.n5555 10.6151
R23853 GND.n5558 GND.n5557 10.6151
R23854 GND.n5557 GND.n5556 10.6151
R23855 GND.n5556 GND.n4940 10.6151
R23856 GND.n5572 GND.n4940 10.6151
R23857 GND.n5573 GND.n5572 10.6151
R23858 GND.n5576 GND.n5573 10.6151
R23859 GND.n5576 GND.n5575 10.6151
R23860 GND.n5575 GND.n5574 10.6151
R23861 GND.n5574 GND.n4930 10.6151
R23862 GND.n5596 GND.n4930 10.6151
R23863 GND.n5597 GND.n5596 10.6151
R23864 GND.n5604 GND.n5597 10.6151
R23865 GND.n5604 GND.n5603 10.6151
R23866 GND.n5603 GND.n5602 10.6151
R23867 GND.n5602 GND.n5599 10.6151
R23868 GND.n5599 GND.n5598 10.6151
R23869 GND.n5598 GND.n4173 10.6151
R23870 GND.n7840 GND.n4173 10.6151
R23871 GND.n7840 GND.n7839 10.6151
R23872 GND.n7839 GND.n7838 10.6151
R23873 GND.n7838 GND.n4174 10.6151
R23874 GND.n4919 GND.n4174 10.6151
R23875 GND.n5658 GND.n4919 10.6151
R23876 GND.n5659 GND.n5658 10.6151
R23877 GND.n5662 GND.n5659 10.6151
R23878 GND.n5662 GND.n5661 10.6151
R23879 GND.n5661 GND.n5660 10.6151
R23880 GND.n5660 GND.n4908 10.6151
R23881 GND.n5676 GND.n4908 10.6151
R23882 GND.n5677 GND.n5676 10.6151
R23883 GND.n5681 GND.n5677 10.6151
R23884 GND.n5681 GND.n5680 10.6151
R23885 GND.n5680 GND.n5679 10.6151
R23886 GND.n5679 GND.n4897 10.6151
R23887 GND.n5699 GND.n4897 10.6151
R23888 GND.n5700 GND.n5699 10.6151
R23889 GND.n5707 GND.n5700 10.6151
R23890 GND.n5707 GND.n5706 10.6151
R23891 GND.n5706 GND.n5705 10.6151
R23892 GND.n5705 GND.n5702 10.6151
R23893 GND.n5702 GND.n5701 10.6151
R23894 GND.n5701 GND.n4275 10.6151
R23895 GND.n7785 GND.n4275 10.6151
R23896 GND.n7785 GND.n7784 10.6151
R23897 GND.n7784 GND.n7783 10.6151
R23898 GND.n7783 GND.n4276 10.6151
R23899 GND.n4885 GND.n4276 10.6151
R23900 GND.n5755 GND.n4885 10.6151
R23901 GND.n5756 GND.n5755 10.6151
R23902 GND.n5759 GND.n5756 10.6151
R23903 GND.n5759 GND.n5758 10.6151
R23904 GND.n5758 GND.n5757 10.6151
R23905 GND.n5757 GND.n4875 10.6151
R23906 GND.n5773 GND.n4875 10.6151
R23907 GND.n5774 GND.n5773 10.6151
R23908 GND.n5776 GND.n5774 10.6151
R23909 GND.n5776 GND.n5775 10.6151
R23910 GND.n5775 GND.n4856 10.6151
R23911 GND.n5798 GND.n4856 10.6151
R23912 GND.n5798 GND.n5797 10.6151
R23913 GND.n5797 GND.n5796 10.6151
R23914 GND.n5796 GND.n4857 10.6151
R23915 GND.n4863 GND.n4857 10.6151
R23916 GND.n4863 GND.n4862 10.6151
R23917 GND.n4862 GND.n4861 10.6151
R23918 GND.n4861 GND.n4859 10.6151
R23919 GND.n4859 GND.n4379 10.6151
R23920 GND.n7730 GND.n4379 10.6151
R23921 GND.n7730 GND.n7729 10.6151
R23922 GND.n7729 GND.n7728 10.6151
R23923 GND.n7728 GND.n4380 10.6151
R23924 GND.n4461 GND.n4380 10.6151
R23925 GND.n4461 GND.n4401 10.6151
R23926 GND.n7716 GND.n4401 10.6151
R23927 GND.n7716 GND.n7715 10.6151
R23928 GND.n7715 GND.n7714 10.6151
R23929 GND.n7714 GND.n4402 10.6151
R23930 GND.n4474 GND.n4402 10.6151
R23931 GND.n4474 GND.n4419 10.6151
R23932 GND.n7702 GND.n4419 10.6151
R23933 GND.n7702 GND.n7701 10.6151
R23934 GND.n7701 GND.n7700 10.6151
R23935 GND.n7700 GND.n4420 10.6151
R23936 GND.n4487 GND.n4420 10.6151
R23937 GND.n4487 GND.n4437 10.6151
R23938 GND.n7688 GND.n4437 10.6151
R23939 GND.n7688 GND.n7687 10.6151
R23940 GND.n7687 GND.n7686 10.6151
R23941 GND.n7686 GND.n4438 10.6151
R23942 GND.n4509 GND.n4438 10.6151
R23943 GND.n4510 GND.n4509 10.6151
R23944 GND.n4511 GND.n4510 10.6151
R23945 GND.n7669 GND.n4511 10.6151
R23946 GND.n7669 GND.n7668 10.6151
R23947 GND.n7668 GND.n7667 10.6151
R23948 GND.n7667 GND.n4512 10.6151
R23949 GND.n4724 GND.n4512 10.6151
R23950 GND.n4725 GND.n4724 10.6151
R23951 GND.t90 GND.n3780 10.0339
R23952 GND.t108 GND.n4527 10.0339
R23953 GND.t208 GND.n4034 9.6995
R23954 GND.n5655 GND.t8 9.6995
R23955 GND.n4665 GND.n4664 9.36635
R23956 GND.n5151 GND.n5150 9.36635
R23957 GND.n5132 GND.n5131 9.36635
R23958 GND.n4781 GND.n4780 9.36635
R23959 GND.n8119 GND.n3772 9.36505
R23960 GND.n8099 GND.n3796 9.36505
R23961 GND.n5305 GND.n5035 9.36505
R23962 GND.n5324 GND.n5030 9.36505
R23963 GND.n7963 GND.n3956 9.36505
R23964 GND.n7945 GND.n3984 9.36505
R23965 GND.n5504 GND.n5503 9.36505
R23966 GND.n7836 GND.n7835 9.36505
R23967 GND.n5710 GND.n5709 9.36505
R23968 GND.n7781 GND.n7780 9.36505
R23969 GND.n5793 GND.n5792 9.36505
R23970 GND.n7726 GND.n7725 9.36505
R23971 GND.n4440 GND.n4434 9.36505
R23972 GND.n3446 GND.n2653 9.3005
R23973 GND.n3448 GND.n3447 9.3005
R23974 GND.n3449 GND.n2652 9.3005
R23975 GND.n3451 GND.n3450 9.3005
R23976 GND.n2481 GND.n2480 9.3005
R23977 GND.n3503 GND.n3502 9.3005
R23978 GND.n3504 GND.n2479 9.3005
R23979 GND.n3508 GND.n3505 9.3005
R23980 GND.n3507 GND.n3506 9.3005
R23981 GND.n2459 GND.n2458 9.3005
R23982 GND.n3529 GND.n3528 9.3005
R23983 GND.n3530 GND.n2457 9.3005
R23984 GND.n3534 GND.n3531 9.3005
R23985 GND.n3533 GND.n3532 9.3005
R23986 GND.n2438 GND.n2437 9.3005
R23987 GND.n3555 GND.n3554 9.3005
R23988 GND.n3556 GND.n2436 9.3005
R23989 GND.n3560 GND.n3557 9.3005
R23990 GND.n3559 GND.n3558 9.3005
R23991 GND.n2417 GND.n2416 9.3005
R23992 GND.n3581 GND.n3580 9.3005
R23993 GND.n3582 GND.n2415 9.3005
R23994 GND.n3586 GND.n3583 9.3005
R23995 GND.n3585 GND.n3584 9.3005
R23996 GND.n2394 GND.n2393 9.3005
R23997 GND.n3606 GND.n3605 9.3005
R23998 GND.n3607 GND.n2392 9.3005
R23999 GND.n3611 GND.n3608 9.3005
R24000 GND.n3610 GND.n3609 9.3005
R24001 GND.n2374 GND.n2373 9.3005
R24002 GND.n3632 GND.n3631 9.3005
R24003 GND.n3633 GND.n2372 9.3005
R24004 GND.n3637 GND.n3634 9.3005
R24005 GND.n3636 GND.n3635 9.3005
R24006 GND.n2354 GND.n2353 9.3005
R24007 GND.n3658 GND.n3657 9.3005
R24008 GND.n3659 GND.n2352 9.3005
R24009 GND.n3663 GND.n3660 9.3005
R24010 GND.n3662 GND.n3661 9.3005
R24011 GND.n2332 GND.n2331 9.3005
R24012 GND.n3684 GND.n3683 9.3005
R24013 GND.n3685 GND.n2330 9.3005
R24014 GND.n3689 GND.n3686 9.3005
R24015 GND.n3688 GND.n3687 9.3005
R24016 GND.n2305 GND.n2304 9.3005
R24017 GND.n8195 GND.n8194 9.3005
R24018 GND.n8196 GND.n2303 9.3005
R24019 GND.n8200 GND.n8197 9.3005
R24020 GND.n8199 GND.n8198 9.3005
R24021 GND.n2283 GND.n2282 9.3005
R24022 GND.n8221 GND.n8220 9.3005
R24023 GND.n8222 GND.n2281 9.3005
R24024 GND.n8226 GND.n8223 9.3005
R24025 GND.n8225 GND.n8224 9.3005
R24026 GND.n2262 GND.n2261 9.3005
R24027 GND.n8247 GND.n8246 9.3005
R24028 GND.n8248 GND.n2260 9.3005
R24029 GND.n8252 GND.n8249 9.3005
R24030 GND.n8251 GND.n8250 9.3005
R24031 GND.n2241 GND.n2240 9.3005
R24032 GND.n8273 GND.n8272 9.3005
R24033 GND.n8274 GND.n2239 9.3005
R24034 GND.n8278 GND.n8275 9.3005
R24035 GND.n8277 GND.n8276 9.3005
R24036 GND.n2218 GND.n2217 9.3005
R24037 GND.n8297 GND.n8296 9.3005
R24038 GND.n8298 GND.n2216 9.3005
R24039 GND.n8302 GND.n8299 9.3005
R24040 GND.n8301 GND.n8300 9.3005
R24041 GND.n9050 GND.n9049 9.3005
R24042 GND.n1459 GND.n1458 9.3005
R24043 GND.n9057 GND.n9056 9.3005
R24044 GND.n9058 GND.n1457 9.3005
R24045 GND.n9060 GND.n9059 9.3005
R24046 GND.n1453 GND.n1452 9.3005
R24047 GND.n9067 GND.n9066 9.3005
R24048 GND.n9068 GND.n1451 9.3005
R24049 GND.n9070 GND.n9069 9.3005
R24050 GND.n1447 GND.n1446 9.3005
R24051 GND.n9077 GND.n9076 9.3005
R24052 GND.n9078 GND.n1445 9.3005
R24053 GND.n9080 GND.n9079 9.3005
R24054 GND.n1441 GND.n1440 9.3005
R24055 GND.n9087 GND.n9086 9.3005
R24056 GND.n9088 GND.n1439 9.3005
R24057 GND.n9090 GND.n9089 9.3005
R24058 GND.n1435 GND.n1434 9.3005
R24059 GND.n9097 GND.n9096 9.3005
R24060 GND.n9098 GND.n1433 9.3005
R24061 GND.n9100 GND.n9099 9.3005
R24062 GND.n1429 GND.n1428 9.3005
R24063 GND.n9107 GND.n9106 9.3005
R24064 GND.n9108 GND.n1427 9.3005
R24065 GND.n9110 GND.n9109 9.3005
R24066 GND.n1423 GND.n1422 9.3005
R24067 GND.n9117 GND.n9116 9.3005
R24068 GND.n9118 GND.n1421 9.3005
R24069 GND.n9120 GND.n9119 9.3005
R24070 GND.n1417 GND.n1416 9.3005
R24071 GND.n9127 GND.n9126 9.3005
R24072 GND.n9128 GND.n1415 9.3005
R24073 GND.n9130 GND.n9129 9.3005
R24074 GND.n1411 GND.n1410 9.3005
R24075 GND.n9137 GND.n9136 9.3005
R24076 GND.n9138 GND.n1409 9.3005
R24077 GND.n9140 GND.n9139 9.3005
R24078 GND.n1405 GND.n1404 9.3005
R24079 GND.n9147 GND.n9146 9.3005
R24080 GND.n9148 GND.n1403 9.3005
R24081 GND.n9150 GND.n9149 9.3005
R24082 GND.n1399 GND.n1398 9.3005
R24083 GND.n9157 GND.n9156 9.3005
R24084 GND.n9158 GND.n1397 9.3005
R24085 GND.n9160 GND.n9159 9.3005
R24086 GND.n1393 GND.n1392 9.3005
R24087 GND.n9167 GND.n9166 9.3005
R24088 GND.n9168 GND.n1391 9.3005
R24089 GND.n9170 GND.n9169 9.3005
R24090 GND.n1387 GND.n1386 9.3005
R24091 GND.n9177 GND.n9176 9.3005
R24092 GND.n9178 GND.n1385 9.3005
R24093 GND.n9180 GND.n9179 9.3005
R24094 GND.n1381 GND.n1380 9.3005
R24095 GND.n9187 GND.n9186 9.3005
R24096 GND.n9188 GND.n1379 9.3005
R24097 GND.n9190 GND.n9189 9.3005
R24098 GND.n1375 GND.n1374 9.3005
R24099 GND.n9197 GND.n9196 9.3005
R24100 GND.n9198 GND.n1373 9.3005
R24101 GND.n9200 GND.n9199 9.3005
R24102 GND.n1369 GND.n1368 9.3005
R24103 GND.n9207 GND.n9206 9.3005
R24104 GND.n9208 GND.n1367 9.3005
R24105 GND.n9210 GND.n9209 9.3005
R24106 GND.n1363 GND.n1362 9.3005
R24107 GND.n9217 GND.n9216 9.3005
R24108 GND.n9218 GND.n1361 9.3005
R24109 GND.n9220 GND.n9219 9.3005
R24110 GND.n1357 GND.n1356 9.3005
R24111 GND.n9227 GND.n9226 9.3005
R24112 GND.n9228 GND.n1355 9.3005
R24113 GND.n9230 GND.n9229 9.3005
R24114 GND.n1351 GND.n1350 9.3005
R24115 GND.n9237 GND.n9236 9.3005
R24116 GND.n9238 GND.n1349 9.3005
R24117 GND.n9240 GND.n9239 9.3005
R24118 GND.n1345 GND.n1344 9.3005
R24119 GND.n9247 GND.n9246 9.3005
R24120 GND.n9248 GND.n1343 9.3005
R24121 GND.n9250 GND.n9249 9.3005
R24122 GND.n1339 GND.n1338 9.3005
R24123 GND.n9257 GND.n9256 9.3005
R24124 GND.n9258 GND.n1337 9.3005
R24125 GND.n9260 GND.n9259 9.3005
R24126 GND.n1333 GND.n1332 9.3005
R24127 GND.n9267 GND.n9266 9.3005
R24128 GND.n9268 GND.n1331 9.3005
R24129 GND.n9270 GND.n9269 9.3005
R24130 GND.n1327 GND.n1326 9.3005
R24131 GND.n9277 GND.n9276 9.3005
R24132 GND.n9278 GND.n1325 9.3005
R24133 GND.n9280 GND.n9279 9.3005
R24134 GND.n1321 GND.n1320 9.3005
R24135 GND.n9287 GND.n9286 9.3005
R24136 GND.n9288 GND.n1319 9.3005
R24137 GND.n9290 GND.n9289 9.3005
R24138 GND.n1315 GND.n1314 9.3005
R24139 GND.n9297 GND.n9296 9.3005
R24140 GND.n9298 GND.n1313 9.3005
R24141 GND.n9300 GND.n9299 9.3005
R24142 GND.n1309 GND.n1308 9.3005
R24143 GND.n9307 GND.n9306 9.3005
R24144 GND.n9308 GND.n1307 9.3005
R24145 GND.n9310 GND.n9309 9.3005
R24146 GND.n1303 GND.n1302 9.3005
R24147 GND.n9317 GND.n9316 9.3005
R24148 GND.n9318 GND.n1301 9.3005
R24149 GND.n9320 GND.n9319 9.3005
R24150 GND.n1297 GND.n1296 9.3005
R24151 GND.n9327 GND.n9326 9.3005
R24152 GND.n9328 GND.n1295 9.3005
R24153 GND.n9330 GND.n9329 9.3005
R24154 GND.n1291 GND.n1290 9.3005
R24155 GND.n9337 GND.n9336 9.3005
R24156 GND.n9338 GND.n1289 9.3005
R24157 GND.n9340 GND.n9339 9.3005
R24158 GND.n1285 GND.n1284 9.3005
R24159 GND.n9347 GND.n9346 9.3005
R24160 GND.n9348 GND.n1283 9.3005
R24161 GND.n9350 GND.n9349 9.3005
R24162 GND.n1279 GND.n1278 9.3005
R24163 GND.n9357 GND.n9356 9.3005
R24164 GND.n9358 GND.n1277 9.3005
R24165 GND.n9360 GND.n9359 9.3005
R24166 GND.n1273 GND.n1272 9.3005
R24167 GND.n9367 GND.n9366 9.3005
R24168 GND.n9368 GND.n1271 9.3005
R24169 GND.n9370 GND.n9369 9.3005
R24170 GND.n1267 GND.n1266 9.3005
R24171 GND.n9377 GND.n9376 9.3005
R24172 GND.n9378 GND.n1265 9.3005
R24173 GND.n9380 GND.n9379 9.3005
R24174 GND.n1261 GND.n1260 9.3005
R24175 GND.n9387 GND.n9386 9.3005
R24176 GND.n9388 GND.n1259 9.3005
R24177 GND.n9390 GND.n9389 9.3005
R24178 GND.n1255 GND.n1254 9.3005
R24179 GND.n9397 GND.n9396 9.3005
R24180 GND.n9398 GND.n1253 9.3005
R24181 GND.n9400 GND.n9399 9.3005
R24182 GND.n1249 GND.n1248 9.3005
R24183 GND.n9407 GND.n9406 9.3005
R24184 GND.n9408 GND.n1247 9.3005
R24185 GND.n9410 GND.n9409 9.3005
R24186 GND.n1243 GND.n1242 9.3005
R24187 GND.n9417 GND.n9416 9.3005
R24188 GND.n9418 GND.n1241 9.3005
R24189 GND.n9420 GND.n9419 9.3005
R24190 GND.n1237 GND.n1236 9.3005
R24191 GND.n9427 GND.n9426 9.3005
R24192 GND.n9428 GND.n1235 9.3005
R24193 GND.n9430 GND.n9429 9.3005
R24194 GND.n1231 GND.n1230 9.3005
R24195 GND.n9437 GND.n9436 9.3005
R24196 GND.n9438 GND.n1229 9.3005
R24197 GND.n9440 GND.n9439 9.3005
R24198 GND.n1225 GND.n1224 9.3005
R24199 GND.n9447 GND.n9446 9.3005
R24200 GND.n9448 GND.n1223 9.3005
R24201 GND.n9450 GND.n9449 9.3005
R24202 GND.n1219 GND.n1218 9.3005
R24203 GND.n9457 GND.n9456 9.3005
R24204 GND.n9458 GND.n1217 9.3005
R24205 GND.n9460 GND.n9459 9.3005
R24206 GND.n1213 GND.n1212 9.3005
R24207 GND.n9467 GND.n9466 9.3005
R24208 GND.n9468 GND.n1211 9.3005
R24209 GND.n9470 GND.n9469 9.3005
R24210 GND.n1207 GND.n1206 9.3005
R24211 GND.n9477 GND.n9476 9.3005
R24212 GND.n9478 GND.n1205 9.3005
R24213 GND.n9480 GND.n9479 9.3005
R24214 GND.n1201 GND.n1200 9.3005
R24215 GND.n9487 GND.n9486 9.3005
R24216 GND.n9488 GND.n1199 9.3005
R24217 GND.n9490 GND.n9489 9.3005
R24218 GND.n1195 GND.n1194 9.3005
R24219 GND.n9497 GND.n9496 9.3005
R24220 GND.n9498 GND.n1193 9.3005
R24221 GND.n9500 GND.n9499 9.3005
R24222 GND.n1189 GND.n1188 9.3005
R24223 GND.n9507 GND.n9506 9.3005
R24224 GND.n9508 GND.n1187 9.3005
R24225 GND.n9510 GND.n9509 9.3005
R24226 GND.n1183 GND.n1182 9.3005
R24227 GND.n9517 GND.n9516 9.3005
R24228 GND.n9518 GND.n1181 9.3005
R24229 GND.n9520 GND.n9519 9.3005
R24230 GND.n1177 GND.n1176 9.3005
R24231 GND.n9527 GND.n9526 9.3005
R24232 GND.n9528 GND.n1175 9.3005
R24233 GND.n9530 GND.n9529 9.3005
R24234 GND.n1171 GND.n1170 9.3005
R24235 GND.n9537 GND.n9536 9.3005
R24236 GND.n9538 GND.n1169 9.3005
R24237 GND.n9540 GND.n9539 9.3005
R24238 GND.n1165 GND.n1164 9.3005
R24239 GND.n9547 GND.n9546 9.3005
R24240 GND.n9548 GND.n1163 9.3005
R24241 GND.n9550 GND.n9549 9.3005
R24242 GND.n1159 GND.n1158 9.3005
R24243 GND.n9557 GND.n9556 9.3005
R24244 GND.n9558 GND.n1157 9.3005
R24245 GND.n9560 GND.n9559 9.3005
R24246 GND.n1153 GND.n1152 9.3005
R24247 GND.n9567 GND.n9566 9.3005
R24248 GND.n9568 GND.n1151 9.3005
R24249 GND.n9570 GND.n9569 9.3005
R24250 GND.n1147 GND.n1146 9.3005
R24251 GND.n9577 GND.n9576 9.3005
R24252 GND.n9578 GND.n1145 9.3005
R24253 GND.n9580 GND.n9579 9.3005
R24254 GND.n1141 GND.n1140 9.3005
R24255 GND.n9587 GND.n9586 9.3005
R24256 GND.n9588 GND.n1139 9.3005
R24257 GND.n9590 GND.n9589 9.3005
R24258 GND.n1135 GND.n1134 9.3005
R24259 GND.n9597 GND.n9596 9.3005
R24260 GND.n9598 GND.n1133 9.3005
R24261 GND.n9600 GND.n9599 9.3005
R24262 GND.n1129 GND.n1128 9.3005
R24263 GND.n9607 GND.n9606 9.3005
R24264 GND.n9608 GND.n1127 9.3005
R24265 GND.n9610 GND.n9609 9.3005
R24266 GND.n1123 GND.n1122 9.3005
R24267 GND.n9617 GND.n9616 9.3005
R24268 GND.n9618 GND.n1121 9.3005
R24269 GND.n9620 GND.n9619 9.3005
R24270 GND.n1117 GND.n1116 9.3005
R24271 GND.n9627 GND.n9626 9.3005
R24272 GND.n9628 GND.n1115 9.3005
R24273 GND.n9630 GND.n9629 9.3005
R24274 GND.n1111 GND.n1110 9.3005
R24275 GND.n9637 GND.n9636 9.3005
R24276 GND.n9638 GND.n1109 9.3005
R24277 GND.n9640 GND.n9639 9.3005
R24278 GND.n1105 GND.n1104 9.3005
R24279 GND.n9647 GND.n9646 9.3005
R24280 GND.n9648 GND.n1103 9.3005
R24281 GND.n9650 GND.n9649 9.3005
R24282 GND.n1099 GND.n1098 9.3005
R24283 GND.n9657 GND.n9656 9.3005
R24284 GND.n9658 GND.n1097 9.3005
R24285 GND.n9660 GND.n9659 9.3005
R24286 GND.n1093 GND.n1092 9.3005
R24287 GND.n9667 GND.n9666 9.3005
R24288 GND.n9668 GND.n1091 9.3005
R24289 GND.n9670 GND.n9669 9.3005
R24290 GND.n1087 GND.n1086 9.3005
R24291 GND.n9677 GND.n9676 9.3005
R24292 GND.n9678 GND.n1085 9.3005
R24293 GND.n9680 GND.n9679 9.3005
R24294 GND.n1081 GND.n1080 9.3005
R24295 GND.n9687 GND.n9686 9.3005
R24296 GND.n9688 GND.n1079 9.3005
R24297 GND.n9690 GND.n9689 9.3005
R24298 GND.n1075 GND.n1074 9.3005
R24299 GND.n9697 GND.n9696 9.3005
R24300 GND.n9698 GND.n1073 9.3005
R24301 GND.n9700 GND.n9699 9.3005
R24302 GND.n1069 GND.n1068 9.3005
R24303 GND.n9707 GND.n9706 9.3005
R24304 GND.n9708 GND.n1067 9.3005
R24305 GND.n9710 GND.n9709 9.3005
R24306 GND.n1063 GND.n1062 9.3005
R24307 GND.n9717 GND.n9716 9.3005
R24308 GND.n9718 GND.n1061 9.3005
R24309 GND.n9720 GND.n9719 9.3005
R24310 GND.n1057 GND.n1056 9.3005
R24311 GND.n9727 GND.n9726 9.3005
R24312 GND.n9728 GND.n1055 9.3005
R24313 GND.n9730 GND.n9729 9.3005
R24314 GND.n1051 GND.n1050 9.3005
R24315 GND.n9737 GND.n9736 9.3005
R24316 GND.n9738 GND.n1049 9.3005
R24317 GND.n9740 GND.n9739 9.3005
R24318 GND.n1045 GND.n1044 9.3005
R24319 GND.n9747 GND.n9746 9.3005
R24320 GND.n9748 GND.n1043 9.3005
R24321 GND.n9750 GND.n9749 9.3005
R24322 GND.n1039 GND.n1038 9.3005
R24323 GND.n9757 GND.n9756 9.3005
R24324 GND.n9758 GND.n1037 9.3005
R24325 GND.n9760 GND.n9759 9.3005
R24326 GND.n1033 GND.n1032 9.3005
R24327 GND.n9767 GND.n9766 9.3005
R24328 GND.n9768 GND.n1031 9.3005
R24329 GND.n9770 GND.n9769 9.3005
R24330 GND.n1027 GND.n1026 9.3005
R24331 GND.n9777 GND.n9776 9.3005
R24332 GND.n9778 GND.n1025 9.3005
R24333 GND.n9780 GND.n9779 9.3005
R24334 GND.n1021 GND.n1020 9.3005
R24335 GND.n9787 GND.n9786 9.3005
R24336 GND.n9788 GND.n1019 9.3005
R24337 GND.n9790 GND.n9789 9.3005
R24338 GND.n1015 GND.n1014 9.3005
R24339 GND.n9797 GND.n9796 9.3005
R24340 GND.n9798 GND.n1013 9.3005
R24341 GND.n9800 GND.n9799 9.3005
R24342 GND.n1009 GND.n1008 9.3005
R24343 GND.n9807 GND.n9806 9.3005
R24344 GND.n9808 GND.n1007 9.3005
R24345 GND.n9810 GND.n9809 9.3005
R24346 GND.n1003 GND.n1002 9.3005
R24347 GND.n9817 GND.n9816 9.3005
R24348 GND.n9818 GND.n1001 9.3005
R24349 GND.n9820 GND.n9819 9.3005
R24350 GND.n997 GND.n996 9.3005
R24351 GND.n9827 GND.n9826 9.3005
R24352 GND.n9828 GND.n995 9.3005
R24353 GND.n9830 GND.n9829 9.3005
R24354 GND.n991 GND.n990 9.3005
R24355 GND.n9837 GND.n9836 9.3005
R24356 GND.n9838 GND.n989 9.3005
R24357 GND.n9840 GND.n9839 9.3005
R24358 GND.n985 GND.n984 9.3005
R24359 GND.n9847 GND.n9846 9.3005
R24360 GND.n9848 GND.n983 9.3005
R24361 GND.n9850 GND.n9849 9.3005
R24362 GND.n979 GND.n978 9.3005
R24363 GND.n9857 GND.n9856 9.3005
R24364 GND.n9858 GND.n977 9.3005
R24365 GND.n9860 GND.n9859 9.3005
R24366 GND.n973 GND.n972 9.3005
R24367 GND.n9867 GND.n9866 9.3005
R24368 GND.n9868 GND.n971 9.3005
R24369 GND.n9870 GND.n9869 9.3005
R24370 GND.n967 GND.n966 9.3005
R24371 GND.n9877 GND.n9876 9.3005
R24372 GND.n9878 GND.n965 9.3005
R24373 GND.n9880 GND.n9879 9.3005
R24374 GND.n961 GND.n960 9.3005
R24375 GND.n9887 GND.n9886 9.3005
R24376 GND.n9888 GND.n959 9.3005
R24377 GND.n9890 GND.n9889 9.3005
R24378 GND.n955 GND.n954 9.3005
R24379 GND.n9897 GND.n9896 9.3005
R24380 GND.n9898 GND.n953 9.3005
R24381 GND.n9900 GND.n9899 9.3005
R24382 GND.n949 GND.n948 9.3005
R24383 GND.n9907 GND.n9906 9.3005
R24384 GND.n9908 GND.n947 9.3005
R24385 GND.n9910 GND.n9909 9.3005
R24386 GND.n943 GND.n942 9.3005
R24387 GND.n9917 GND.n9916 9.3005
R24388 GND.n9918 GND.n941 9.3005
R24389 GND.n9920 GND.n9919 9.3005
R24390 GND.n937 GND.n936 9.3005
R24391 GND.n9927 GND.n9926 9.3005
R24392 GND.n9928 GND.n935 9.3005
R24393 GND.n9930 GND.n9929 9.3005
R24394 GND.n931 GND.n930 9.3005
R24395 GND.n9937 GND.n9936 9.3005
R24396 GND.n9938 GND.n929 9.3005
R24397 GND.n9940 GND.n9939 9.3005
R24398 GND.n925 GND.n924 9.3005
R24399 GND.n9947 GND.n9946 9.3005
R24400 GND.n9948 GND.n923 9.3005
R24401 GND.n9950 GND.n9949 9.3005
R24402 GND.n919 GND.n918 9.3005
R24403 GND.n9957 GND.n9956 9.3005
R24404 GND.n9958 GND.n917 9.3005
R24405 GND.n9960 GND.n9959 9.3005
R24406 GND.n913 GND.n912 9.3005
R24407 GND.n9967 GND.n9966 9.3005
R24408 GND.n9968 GND.n911 9.3005
R24409 GND.n9970 GND.n9969 9.3005
R24410 GND.n907 GND.n906 9.3005
R24411 GND.n9977 GND.n9976 9.3005
R24412 GND.n9978 GND.n905 9.3005
R24413 GND.n9980 GND.n9979 9.3005
R24414 GND.n901 GND.n900 9.3005
R24415 GND.n9987 GND.n9986 9.3005
R24416 GND.n9988 GND.n899 9.3005
R24417 GND.n9990 GND.n9989 9.3005
R24418 GND.n895 GND.n894 9.3005
R24419 GND.n9997 GND.n9996 9.3005
R24420 GND.n9998 GND.n893 9.3005
R24421 GND.n10000 GND.n9999 9.3005
R24422 GND.n889 GND.n888 9.3005
R24423 GND.n10007 GND.n10006 9.3005
R24424 GND.n10008 GND.n887 9.3005
R24425 GND.n10010 GND.n10009 9.3005
R24426 GND.n883 GND.n882 9.3005
R24427 GND.n10017 GND.n10016 9.3005
R24428 GND.n10018 GND.n881 9.3005
R24429 GND.n10020 GND.n10019 9.3005
R24430 GND.n877 GND.n876 9.3005
R24431 GND.n10027 GND.n10026 9.3005
R24432 GND.n10028 GND.n875 9.3005
R24433 GND.n10030 GND.n10029 9.3005
R24434 GND.n871 GND.n870 9.3005
R24435 GND.n10037 GND.n10036 9.3005
R24436 GND.n10038 GND.n869 9.3005
R24437 GND.n10040 GND.n10039 9.3005
R24438 GND.n865 GND.n864 9.3005
R24439 GND.n10047 GND.n10046 9.3005
R24440 GND.n10048 GND.n863 9.3005
R24441 GND.n10050 GND.n10049 9.3005
R24442 GND.n859 GND.n858 9.3005
R24443 GND.n10057 GND.n10056 9.3005
R24444 GND.n10058 GND.n857 9.3005
R24445 GND.n10060 GND.n10059 9.3005
R24446 GND.n853 GND.n852 9.3005
R24447 GND.n10067 GND.n10066 9.3005
R24448 GND.n10068 GND.n851 9.3005
R24449 GND.n10070 GND.n10069 9.3005
R24450 GND.n847 GND.n846 9.3005
R24451 GND.n10077 GND.n10076 9.3005
R24452 GND.n10078 GND.n845 9.3005
R24453 GND.n10080 GND.n10079 9.3005
R24454 GND.n841 GND.n840 9.3005
R24455 GND.n10087 GND.n10086 9.3005
R24456 GND.n10088 GND.n839 9.3005
R24457 GND.n10090 GND.n10089 9.3005
R24458 GND.n835 GND.n834 9.3005
R24459 GND.n10097 GND.n10096 9.3005
R24460 GND.n10098 GND.n833 9.3005
R24461 GND.n10100 GND.n10099 9.3005
R24462 GND.n829 GND.n828 9.3005
R24463 GND.n10107 GND.n10106 9.3005
R24464 GND.n10108 GND.n827 9.3005
R24465 GND.n10110 GND.n10109 9.3005
R24466 GND.n823 GND.n822 9.3005
R24467 GND.n10117 GND.n10116 9.3005
R24468 GND.n10118 GND.n821 9.3005
R24469 GND.n10120 GND.n10119 9.3005
R24470 GND.n817 GND.n816 9.3005
R24471 GND.n10127 GND.n10126 9.3005
R24472 GND.n10128 GND.n815 9.3005
R24473 GND.n10130 GND.n10129 9.3005
R24474 GND.n811 GND.n810 9.3005
R24475 GND.n10137 GND.n10136 9.3005
R24476 GND.n10138 GND.n809 9.3005
R24477 GND.n10140 GND.n10139 9.3005
R24478 GND.n805 GND.n804 9.3005
R24479 GND.n10147 GND.n10146 9.3005
R24480 GND.n10148 GND.n803 9.3005
R24481 GND.n10150 GND.n10149 9.3005
R24482 GND.n799 GND.n798 9.3005
R24483 GND.n10157 GND.n10156 9.3005
R24484 GND.n10158 GND.n797 9.3005
R24485 GND.n10160 GND.n10159 9.3005
R24486 GND.n793 GND.n792 9.3005
R24487 GND.n10167 GND.n10166 9.3005
R24488 GND.n10168 GND.n791 9.3005
R24489 GND.n10170 GND.n10169 9.3005
R24490 GND.n787 GND.n786 9.3005
R24491 GND.n10177 GND.n10176 9.3005
R24492 GND.n10178 GND.n785 9.3005
R24493 GND.n10180 GND.n10179 9.3005
R24494 GND.n781 GND.n780 9.3005
R24495 GND.n10187 GND.n10186 9.3005
R24496 GND.n10188 GND.n779 9.3005
R24497 GND.n10190 GND.n10189 9.3005
R24498 GND.n775 GND.n774 9.3005
R24499 GND.n10197 GND.n10196 9.3005
R24500 GND.n10198 GND.n773 9.3005
R24501 GND.n10200 GND.n10199 9.3005
R24502 GND.n769 GND.n768 9.3005
R24503 GND.n10207 GND.n10206 9.3005
R24504 GND.n10208 GND.n767 9.3005
R24505 GND.n10210 GND.n10209 9.3005
R24506 GND.n763 GND.n762 9.3005
R24507 GND.n10217 GND.n10216 9.3005
R24508 GND.n10218 GND.n761 9.3005
R24509 GND.n10220 GND.n10219 9.3005
R24510 GND.n757 GND.n756 9.3005
R24511 GND.n10227 GND.n10226 9.3005
R24512 GND.n10228 GND.n755 9.3005
R24513 GND.n10230 GND.n10229 9.3005
R24514 GND.n751 GND.n750 9.3005
R24515 GND.n10237 GND.n10236 9.3005
R24516 GND.n10238 GND.n749 9.3005
R24517 GND.n10240 GND.n10239 9.3005
R24518 GND.n745 GND.n744 9.3005
R24519 GND.n10247 GND.n10246 9.3005
R24520 GND.n10248 GND.n743 9.3005
R24521 GND.n10250 GND.n10249 9.3005
R24522 GND.n739 GND.n738 9.3005
R24523 GND.n10257 GND.n10256 9.3005
R24524 GND.n10258 GND.n737 9.3005
R24525 GND.n10260 GND.n10259 9.3005
R24526 GND.n733 GND.n732 9.3005
R24527 GND.n10267 GND.n10266 9.3005
R24528 GND.n10268 GND.n731 9.3005
R24529 GND.n10270 GND.n10269 9.3005
R24530 GND.n727 GND.n726 9.3005
R24531 GND.n10277 GND.n10276 9.3005
R24532 GND.n10278 GND.n725 9.3005
R24533 GND.n10280 GND.n10279 9.3005
R24534 GND.n721 GND.n720 9.3005
R24535 GND.n10287 GND.n10286 9.3005
R24536 GND.n10288 GND.n719 9.3005
R24537 GND.n10290 GND.n10289 9.3005
R24538 GND.n715 GND.n714 9.3005
R24539 GND.n10297 GND.n10296 9.3005
R24540 GND.n10298 GND.n713 9.3005
R24541 GND.n10300 GND.n10299 9.3005
R24542 GND.n709 GND.n708 9.3005
R24543 GND.n10307 GND.n10306 9.3005
R24544 GND.n10308 GND.n707 9.3005
R24545 GND.n10310 GND.n10309 9.3005
R24546 GND.n703 GND.n702 9.3005
R24547 GND.n10317 GND.n10316 9.3005
R24548 GND.n10318 GND.n701 9.3005
R24549 GND.n10320 GND.n10319 9.3005
R24550 GND.n697 GND.n696 9.3005
R24551 GND.n10327 GND.n10326 9.3005
R24552 GND.n10328 GND.n695 9.3005
R24553 GND.n10330 GND.n10329 9.3005
R24554 GND.n691 GND.n690 9.3005
R24555 GND.n10337 GND.n10336 9.3005
R24556 GND.n10338 GND.n689 9.3005
R24557 GND.n10340 GND.n10339 9.3005
R24558 GND.n685 GND.n684 9.3005
R24559 GND.n10347 GND.n10346 9.3005
R24560 GND.n10348 GND.n683 9.3005
R24561 GND.n10350 GND.n10349 9.3005
R24562 GND.n679 GND.n678 9.3005
R24563 GND.n10357 GND.n10356 9.3005
R24564 GND.n10358 GND.n677 9.3005
R24565 GND.n10360 GND.n10359 9.3005
R24566 GND.n673 GND.n672 9.3005
R24567 GND.n10367 GND.n10366 9.3005
R24568 GND.n10368 GND.n671 9.3005
R24569 GND.n10370 GND.n10369 9.3005
R24570 GND.n667 GND.n666 9.3005
R24571 GND.n10377 GND.n10376 9.3005
R24572 GND.n10378 GND.n665 9.3005
R24573 GND.n10381 GND.n10379 9.3005
R24574 GND.n10380 GND.n661 9.3005
R24575 GND.n10389 GND.n660 9.3005
R24576 GND.n10391 GND.n10390 9.3005
R24577 GND.n656 GND.n655 9.3005
R24578 GND.n10398 GND.n10397 9.3005
R24579 GND.n10399 GND.n654 9.3005
R24580 GND.n10401 GND.n10400 9.3005
R24581 GND.n650 GND.n649 9.3005
R24582 GND.n10408 GND.n10407 9.3005
R24583 GND.n10409 GND.n648 9.3005
R24584 GND.n10411 GND.n10410 9.3005
R24585 GND.n644 GND.n643 9.3005
R24586 GND.n10418 GND.n10417 9.3005
R24587 GND.n10419 GND.n642 9.3005
R24588 GND.n10421 GND.n10420 9.3005
R24589 GND.n638 GND.n637 9.3005
R24590 GND.n10428 GND.n10427 9.3005
R24591 GND.n10429 GND.n636 9.3005
R24592 GND.n10431 GND.n10430 9.3005
R24593 GND.n632 GND.n631 9.3005
R24594 GND.n10438 GND.n10437 9.3005
R24595 GND.n10439 GND.n630 9.3005
R24596 GND.n10441 GND.n10440 9.3005
R24597 GND.n626 GND.n625 9.3005
R24598 GND.n10448 GND.n10447 9.3005
R24599 GND.n10449 GND.n624 9.3005
R24600 GND.n10451 GND.n10450 9.3005
R24601 GND.n620 GND.n619 9.3005
R24602 GND.n10458 GND.n10457 9.3005
R24603 GND.n10459 GND.n618 9.3005
R24604 GND.n10461 GND.n10460 9.3005
R24605 GND.n614 GND.n613 9.3005
R24606 GND.n10468 GND.n10467 9.3005
R24607 GND.n10469 GND.n612 9.3005
R24608 GND.n10471 GND.n10470 9.3005
R24609 GND.n608 GND.n607 9.3005
R24610 GND.n10478 GND.n10477 9.3005
R24611 GND.n10479 GND.n606 9.3005
R24612 GND.n10481 GND.n10480 9.3005
R24613 GND.n602 GND.n601 9.3005
R24614 GND.n10488 GND.n10487 9.3005
R24615 GND.n10489 GND.n600 9.3005
R24616 GND.n10491 GND.n10490 9.3005
R24617 GND.n596 GND.n595 9.3005
R24618 GND.n10498 GND.n10497 9.3005
R24619 GND.n10499 GND.n594 9.3005
R24620 GND.n10501 GND.n10500 9.3005
R24621 GND.n590 GND.n589 9.3005
R24622 GND.n10508 GND.n10507 9.3005
R24623 GND.n10509 GND.n588 9.3005
R24624 GND.n10511 GND.n10510 9.3005
R24625 GND.n584 GND.n583 9.3005
R24626 GND.n10518 GND.n10517 9.3005
R24627 GND.n10519 GND.n582 9.3005
R24628 GND.n10521 GND.n10520 9.3005
R24629 GND.n578 GND.n577 9.3005
R24630 GND.n10528 GND.n10527 9.3005
R24631 GND.n10529 GND.n576 9.3005
R24632 GND.n10532 GND.n10531 9.3005
R24633 GND.n10388 GND.n10387 9.3005
R24634 GND.n5028 GND.n5027 9.3005
R24635 GND.n5029 GND.n5022 9.3005
R24636 GND.n5327 GND.n5326 9.3005
R24637 GND.n5328 GND.n5021 9.3005
R24638 GND.n5330 GND.n5329 9.3005
R24639 GND.n5014 GND.n5013 9.3005
R24640 GND.n5346 GND.n5345 9.3005
R24641 GND.n5347 GND.n5012 9.3005
R24642 GND.n5349 GND.n5348 9.3005
R24643 GND.n5005 GND.n5004 9.3005
R24644 GND.n5365 GND.n5364 9.3005
R24645 GND.n5366 GND.n5003 9.3005
R24646 GND.n5409 GND.n5367 9.3005
R24647 GND.n5408 GND.n5368 9.3005
R24648 GND.n5407 GND.n5369 9.3005
R24649 GND.n5405 GND.n5370 9.3005
R24650 GND.n5404 GND.n5371 9.3005
R24651 GND.n5403 GND.n5372 9.3005
R24652 GND.n5402 GND.n5373 9.3005
R24653 GND.n5400 GND.n5374 9.3005
R24654 GND.n5399 GND.n5375 9.3005
R24655 GND.n5396 GND.n5376 9.3005
R24656 GND.n5395 GND.n5377 9.3005
R24657 GND.n5393 GND.n5378 9.3005
R24658 GND.n5392 GND.n5379 9.3005
R24659 GND.n5390 GND.n5380 9.3005
R24660 GND.n5389 GND.n5381 9.3005
R24661 GND.n5387 GND.n5382 9.3005
R24662 GND.n5386 GND.n5384 9.3005
R24663 GND.n5383 GND.n4957 9.3005
R24664 GND.n5506 GND.n4956 9.3005
R24665 GND.n5508 GND.n5507 9.3005
R24666 GND.n5509 GND.n4955 9.3005
R24667 GND.n5511 GND.n5510 9.3005
R24668 GND.n5512 GND.n4952 9.3005
R24669 GND.n5516 GND.n5515 9.3005
R24670 GND.n5517 GND.n4951 9.3005
R24671 GND.n5540 GND.n5518 9.3005
R24672 GND.n5539 GND.n5519 9.3005
R24673 GND.n5538 GND.n5520 9.3005
R24674 GND.n5536 GND.n5521 9.3005
R24675 GND.n5535 GND.n5522 9.3005
R24676 GND.n5533 GND.n5523 9.3005
R24677 GND.n5532 GND.n5524 9.3005
R24678 GND.n5530 GND.n5525 9.3005
R24679 GND.n5529 GND.n5527 9.3005
R24680 GND.n5526 GND.n4926 9.3005
R24681 GND.n5609 GND.n4925 9.3005
R24682 GND.n5611 GND.n5610 9.3005
R24683 GND.n5612 GND.n4924 9.3005
R24684 GND.n5614 GND.n5613 9.3005
R24685 GND.n5615 GND.n4921 9.3005
R24686 GND.n5619 GND.n5618 9.3005
R24687 GND.n5620 GND.n4920 9.3005
R24688 GND.n5644 GND.n5621 9.3005
R24689 GND.n5643 GND.n5622 9.3005
R24690 GND.n5642 GND.n5623 9.3005
R24691 GND.n5640 GND.n5624 9.3005
R24692 GND.n5639 GND.n5625 9.3005
R24693 GND.n5637 GND.n5626 9.3005
R24694 GND.n5636 GND.n5627 9.3005
R24695 GND.n5634 GND.n5628 9.3005
R24696 GND.n5633 GND.n5630 9.3005
R24697 GND.n5629 GND.n4892 9.3005
R24698 GND.n5712 GND.n4891 9.3005
R24699 GND.n5714 GND.n5713 9.3005
R24700 GND.n5715 GND.n4890 9.3005
R24701 GND.n5717 GND.n5716 9.3005
R24702 GND.n5718 GND.n4887 9.3005
R24703 GND.n5722 GND.n5721 9.3005
R24704 GND.n5723 GND.n4886 9.3005
R24705 GND.n5741 GND.n5724 9.3005
R24706 GND.n5740 GND.n5725 9.3005
R24707 GND.n5739 GND.n5726 9.3005
R24708 GND.n5737 GND.n5727 9.3005
R24709 GND.n5736 GND.n5728 9.3005
R24710 GND.n5734 GND.n5729 9.3005
R24711 GND.n5733 GND.n5731 9.3005
R24712 GND.n5730 GND.n4852 9.3005
R24713 GND.n5803 GND.n4851 9.3005
R24714 GND.n5805 GND.n5804 9.3005
R24715 GND.n5806 GND.n4850 9.3005
R24716 GND.n5808 GND.n5807 9.3005
R24717 GND.n5811 GND.n4849 9.3005
R24718 GND.n5813 GND.n5812 9.3005
R24719 GND.n5026 GND.n5023 9.3005
R24720 GND.n8045 GND.n3870 9.3005
R24721 GND.n8048 GND.n3869 9.3005
R24722 GND.n8050 GND.n3868 9.3005
R24723 GND.n8051 GND.n3867 9.3005
R24724 GND.n8052 GND.n3866 9.3005
R24725 GND.n8053 GND.n3865 9.3005
R24726 GND.n8008 GND.n3874 9.3005
R24727 GND.n3899 GND.n3897 9.3005
R24728 GND.n7997 GND.n3900 9.3005
R24729 GND.n7996 GND.n3901 9.3005
R24730 GND.n7995 GND.n3902 9.3005
R24731 GND.n3918 GND.n3903 9.3005
R24732 GND.n7985 GND.n3919 9.3005
R24733 GND.n7984 GND.n3920 9.3005
R24734 GND.n7983 GND.n3921 9.3005
R24735 GND.n3938 GND.n3922 9.3005
R24736 GND.n7973 GND.n3939 9.3005
R24737 GND.n7972 GND.n3940 9.3005
R24738 GND.n7971 GND.n3941 9.3005
R24739 GND.n3958 GND.n3942 9.3005
R24740 GND.n7961 GND.n3959 9.3005
R24741 GND.n7960 GND.n3960 9.3005
R24742 GND.n7959 GND.n3961 9.3005
R24743 GND.n3978 GND.n3962 9.3005
R24744 GND.n7949 GND.n3979 9.3005
R24745 GND.n7948 GND.n3980 9.3005
R24746 GND.n7947 GND.n3981 9.3005
R24747 GND.n3998 GND.n3982 9.3005
R24748 GND.n7937 GND.n3999 9.3005
R24749 GND.n7936 GND.n4000 9.3005
R24750 GND.n7935 GND.n4001 9.3005
R24751 GND.n4018 GND.n4002 9.3005
R24752 GND.n7925 GND.n4019 9.3005
R24753 GND.n7924 GND.n4020 9.3005
R24754 GND.n7923 GND.n4021 9.3005
R24755 GND.n4038 GND.n4022 9.3005
R24756 GND.n7913 GND.n4039 9.3005
R24757 GND.n7912 GND.n4040 9.3005
R24758 GND.n7911 GND.n4041 9.3005
R24759 GND.n4094 GND.n4042 9.3005
R24760 GND.n4095 GND.n4093 9.3005
R24761 GND.n4097 GND.n4096 9.3005
R24762 GND.n4100 GND.n4092 9.3005
R24763 GND.n4102 GND.n4101 9.3005
R24764 GND.n4103 GND.n4091 9.3005
R24765 GND.n7882 GND.n4104 9.3005
R24766 GND.n7881 GND.n4105 9.3005
R24767 GND.n7880 GND.n4106 9.3005
R24768 GND.n4123 GND.n4107 9.3005
R24769 GND.n7870 GND.n4124 9.3005
R24770 GND.n7869 GND.n4125 9.3005
R24771 GND.n7868 GND.n4126 9.3005
R24772 GND.n4143 GND.n4127 9.3005
R24773 GND.n7858 GND.n4144 9.3005
R24774 GND.n7857 GND.n4145 9.3005
R24775 GND.n7856 GND.n4146 9.3005
R24776 GND.n4198 GND.n4147 9.3005
R24777 GND.n4199 GND.n4197 9.3005
R24778 GND.n4201 GND.n4200 9.3005
R24779 GND.n4204 GND.n4196 9.3005
R24780 GND.n4206 GND.n4205 9.3005
R24781 GND.n4207 GND.n4195 9.3005
R24782 GND.n7827 GND.n4208 9.3005
R24783 GND.n7826 GND.n4209 9.3005
R24784 GND.n7825 GND.n4210 9.3005
R24785 GND.n4227 GND.n4211 9.3005
R24786 GND.n7815 GND.n4228 9.3005
R24787 GND.n7814 GND.n4229 9.3005
R24788 GND.n7813 GND.n4230 9.3005
R24789 GND.n4245 GND.n4231 9.3005
R24790 GND.n7803 GND.n4246 9.3005
R24791 GND.n7802 GND.n4247 9.3005
R24792 GND.n7801 GND.n4248 9.3005
R24793 GND.n4301 GND.n4249 9.3005
R24794 GND.n4302 GND.n4300 9.3005
R24795 GND.n4304 GND.n4303 9.3005
R24796 GND.n4307 GND.n4299 9.3005
R24797 GND.n4309 GND.n4308 9.3005
R24798 GND.n4310 GND.n4298 9.3005
R24799 GND.n7772 GND.n4311 9.3005
R24800 GND.n7771 GND.n4312 9.3005
R24801 GND.n7770 GND.n4313 9.3005
R24802 GND.n4330 GND.n4314 9.3005
R24803 GND.n7760 GND.n4331 9.3005
R24804 GND.n7759 GND.n4332 9.3005
R24805 GND.n7758 GND.n4333 9.3005
R24806 GND.n4349 GND.n4334 9.3005
R24807 GND.n7748 GND.n4350 9.3005
R24808 GND.n7747 GND.n4351 9.3005
R24809 GND.n7746 GND.n4352 9.3005
R24810 GND.n4831 GND.n4353 9.3005
R24811 GND.n4833 GND.n4832 9.3005
R24812 GND.n3898 GND.n3880 9.3005
R24813 GND.n4844 GND.n4834 9.3005
R24814 GND.n5820 GND.n5819 9.3005
R24815 GND.n5821 GND.n4848 9.3005
R24816 GND.n5824 GND.n5823 9.3005
R24817 GND.n5822 GND.n4846 9.3005
R24818 GND.n5829 GND.n4830 9.3005
R24819 GND.n5815 GND.n5814 9.3005
R24820 GND.n5872 GND.n4841 9.3005
R24821 GND.n5872 GND.n5871 9.3005
R24822 GND.n6741 GND.n6738 9.3005
R24823 GND.n6748 GND.n6747 9.3005
R24824 GND.n6749 GND.n6737 9.3005
R24825 GND.n6751 GND.n6750 9.3005
R24826 GND.n6735 GND.n6734 9.3005
R24827 GND.n6763 GND.n6762 9.3005
R24828 GND.n6764 GND.n6733 9.3005
R24829 GND.n6766 GND.n6765 9.3005
R24830 GND.n6529 GND.n6528 9.3005
R24831 GND.n6778 GND.n6777 9.3005
R24832 GND.n6779 GND.n6527 9.3005
R24833 GND.n6781 GND.n6780 9.3005
R24834 GND.n6525 GND.n6524 9.3005
R24835 GND.n6793 GND.n6792 9.3005
R24836 GND.n6794 GND.n6523 9.3005
R24837 GND.n6796 GND.n6795 9.3005
R24838 GND.n6521 GND.n6520 9.3005
R24839 GND.n6808 GND.n6807 9.3005
R24840 GND.n6809 GND.n6519 9.3005
R24841 GND.n6811 GND.n6810 9.3005
R24842 GND.n6517 GND.n6516 9.3005
R24843 GND.n6823 GND.n6822 9.3005
R24844 GND.n6824 GND.n6515 9.3005
R24845 GND.n6826 GND.n6825 9.3005
R24846 GND.n6512 GND.n6511 9.3005
R24847 GND.n6838 GND.n6837 9.3005
R24848 GND.n6839 GND.n6510 9.3005
R24849 GND.n6841 GND.n6840 9.3005
R24850 GND.n6508 GND.n6507 9.3005
R24851 GND.n6853 GND.n6852 9.3005
R24852 GND.n6854 GND.n6506 9.3005
R24853 GND.n6856 GND.n6855 9.3005
R24854 GND.n6504 GND.n6503 9.3005
R24855 GND.n6868 GND.n6867 9.3005
R24856 GND.n6869 GND.n6502 9.3005
R24857 GND.n6871 GND.n6870 9.3005
R24858 GND.n6500 GND.n6499 9.3005
R24859 GND.n6883 GND.n6882 9.3005
R24860 GND.n6884 GND.n6498 9.3005
R24861 GND.n6886 GND.n6885 9.3005
R24862 GND.n6496 GND.n6495 9.3005
R24863 GND.n6898 GND.n6897 9.3005
R24864 GND.n6899 GND.n6494 9.3005
R24865 GND.n6901 GND.n6900 9.3005
R24866 GND.n6492 GND.n6491 9.3005
R24867 GND.n6913 GND.n6912 9.3005
R24868 GND.n6914 GND.n6490 9.3005
R24869 GND.n6916 GND.n6915 9.3005
R24870 GND.n6487 GND.n6486 9.3005
R24871 GND.n6928 GND.n6927 9.3005
R24872 GND.n6929 GND.n6485 9.3005
R24873 GND.n6931 GND.n6930 9.3005
R24874 GND.n6483 GND.n6482 9.3005
R24875 GND.n6943 GND.n6942 9.3005
R24876 GND.n6944 GND.n6481 9.3005
R24877 GND.n6946 GND.n6945 9.3005
R24878 GND.n6479 GND.n6478 9.3005
R24879 GND.n6958 GND.n6957 9.3005
R24880 GND.n6959 GND.n6477 9.3005
R24881 GND.n6961 GND.n6960 9.3005
R24882 GND.n6475 GND.n6474 9.3005
R24883 GND.n6973 GND.n6972 9.3005
R24884 GND.n6974 GND.n6473 9.3005
R24885 GND.n6983 GND.n6975 9.3005
R24886 GND.n6982 GND.n6976 9.3005
R24887 GND.n6981 GND.n6977 9.3005
R24888 GND.n6980 GND.n6978 9.3005
R24889 GND.n88 GND.n86 9.3005
R24890 GND.n6740 GND.n6739 9.3005
R24891 GND.n11114 GND.n11113 9.3005
R24892 GND.n89 GND.n87 9.3005
R24893 GND.n6273 GND.n6272 9.3005
R24894 GND.n7316 GND.n6274 9.3005
R24895 GND.n7315 GND.n6275 9.3005
R24896 GND.n7314 GND.n6276 9.3005
R24897 GND.n6462 GND.n6277 9.3005
R24898 GND.n7020 GND.n7019 9.3005
R24899 GND.n7021 GND.n6461 9.3005
R24900 GND.n7023 GND.n7022 9.3005
R24901 GND.n6459 GND.n6458 9.3005
R24902 GND.n7035 GND.n7034 9.3005
R24903 GND.n7036 GND.n6457 9.3005
R24904 GND.n7038 GND.n7037 9.3005
R24905 GND.n6455 GND.n6454 9.3005
R24906 GND.n7050 GND.n7049 9.3005
R24907 GND.n7051 GND.n6453 9.3005
R24908 GND.n7053 GND.n7052 9.3005
R24909 GND.n6451 GND.n6450 9.3005
R24910 GND.n7065 GND.n7064 9.3005
R24911 GND.n7066 GND.n6449 9.3005
R24912 GND.n7068 GND.n7067 9.3005
R24913 GND.n6447 GND.n6446 9.3005
R24914 GND.n7080 GND.n7079 9.3005
R24915 GND.n7081 GND.n6445 9.3005
R24916 GND.n7083 GND.n7082 9.3005
R24917 GND.n6443 GND.n6442 9.3005
R24918 GND.n7095 GND.n7094 9.3005
R24919 GND.n7096 GND.n6441 9.3005
R24920 GND.n7099 GND.n7098 9.3005
R24921 GND.n7097 GND.n6435 9.3005
R24922 GND.n7266 GND.n6436 9.3005
R24923 GND.n7265 GND.n6437 9.3005
R24924 GND.n7264 GND.n6438 9.3005
R24925 GND.n7110 GND.n6439 9.3005
R24926 GND.n7254 GND.n7111 9.3005
R24927 GND.n7253 GND.n7112 9.3005
R24928 GND.n7252 GND.n7113 9.3005
R24929 GND.n7117 GND.n7114 9.3005
R24930 GND.n7242 GND.n7118 9.3005
R24931 GND.n7241 GND.n7119 9.3005
R24932 GND.n7240 GND.n7120 9.3005
R24933 GND.n7124 GND.n7121 9.3005
R24934 GND.n7230 GND.n7125 9.3005
R24935 GND.n7229 GND.n7126 9.3005
R24936 GND.n7228 GND.n7127 9.3005
R24937 GND.n7131 GND.n7128 9.3005
R24938 GND.n7218 GND.n7132 9.3005
R24939 GND.n7217 GND.n7133 9.3005
R24940 GND.n7216 GND.n7134 9.3005
R24941 GND.n7138 GND.n7135 9.3005
R24942 GND.n7206 GND.n7139 9.3005
R24943 GND.n7205 GND.n7140 9.3005
R24944 GND.n7204 GND.n7141 9.3005
R24945 GND.n7145 GND.n7142 9.3005
R24946 GND.n7194 GND.n7146 9.3005
R24947 GND.n7193 GND.n7147 9.3005
R24948 GND.n7192 GND.n7148 9.3005
R24949 GND.n7152 GND.n7149 9.3005
R24950 GND.n7182 GND.n7153 9.3005
R24951 GND.n7181 GND.n7154 9.3005
R24952 GND.n7180 GND.n7155 9.3005
R24953 GND.n7159 GND.n7156 9.3005
R24954 GND.n7170 GND.n7160 9.3005
R24955 GND.n7169 GND.n7161 9.3005
R24956 GND.n7168 GND.n7163 9.3005
R24957 GND.n7162 GND.n453 9.3005
R24958 GND.n10903 GND.n454 9.3005
R24959 GND.n10902 GND.n10901 9.3005
R24960 GND.n10685 GND.n10684 9.3005
R24961 GND.n10683 GND.n10654 9.3005
R24962 GND.n10682 GND.n10681 9.3005
R24963 GND.n10678 GND.n10656 9.3005
R24964 GND.n10677 GND.n10657 9.3005
R24965 GND.n10674 GND.n10658 9.3005
R24966 GND.n10673 GND.n10659 9.3005
R24967 GND.n10670 GND.n10660 9.3005
R24968 GND.n10669 GND.n10661 9.3005
R24969 GND.n10666 GND.n10662 9.3005
R24970 GND.n10665 GND.n10663 9.3005
R24971 GND.n458 GND.n455 9.3005
R24972 GND.n10900 GND.n10899 9.3005
R24973 GND.n10655 GND.n10653 9.3005
R24974 GND.n10720 GND.n10717 9.3005
R24975 GND.n10893 GND.n10721 9.3005
R24976 GND.n10892 GND.n10722 9.3005
R24977 GND.n10891 GND.n10723 9.3005
R24978 GND.n10888 GND.n10724 9.3005
R24979 GND.n10887 GND.n10725 9.3005
R24980 GND.n10884 GND.n10726 9.3005
R24981 GND.n10883 GND.n10727 9.3005
R24982 GND.n10880 GND.n10728 9.3005
R24983 GND.n10879 GND.n10729 9.3005
R24984 GND.n10876 GND.n10730 9.3005
R24985 GND.n10875 GND.n10874 9.3005
R24986 GND.n10873 GND.n10731 9.3005
R24987 GND.n10872 GND.n10871 9.3005
R24988 GND.n10868 GND.n10736 9.3005
R24989 GND.n10867 GND.n10737 9.3005
R24990 GND.n10864 GND.n10738 9.3005
R24991 GND.n10863 GND.n10739 9.3005
R24992 GND.n10860 GND.n10740 9.3005
R24993 GND.n10859 GND.n10741 9.3005
R24994 GND.n10856 GND.n10742 9.3005
R24995 GND.n10855 GND.n10743 9.3005
R24996 GND.n10852 GND.n10744 9.3005
R24997 GND.n10851 GND.n10745 9.3005
R24998 GND.n10848 GND.n10746 9.3005
R24999 GND.n10847 GND.n10747 9.3005
R25000 GND.n10844 GND.n10751 9.3005
R25001 GND.n10843 GND.n10752 9.3005
R25002 GND.n10840 GND.n10753 9.3005
R25003 GND.n10839 GND.n10754 9.3005
R25004 GND.n10836 GND.n10755 9.3005
R25005 GND.n10835 GND.n10756 9.3005
R25006 GND.n10832 GND.n10757 9.3005
R25007 GND.n10831 GND.n10758 9.3005
R25008 GND.n10828 GND.n10759 9.3005
R25009 GND.n10827 GND.n10760 9.3005
R25010 GND.n10824 GND.n10761 9.3005
R25011 GND.n10823 GND.n10762 9.3005
R25012 GND.n10820 GND.n10763 9.3005
R25013 GND.n10819 GND.n10764 9.3005
R25014 GND.n10816 GND.n10768 9.3005
R25015 GND.n10815 GND.n10769 9.3005
R25016 GND.n10812 GND.n10770 9.3005
R25017 GND.n10811 GND.n10771 9.3005
R25018 GND.n10808 GND.n10772 9.3005
R25019 GND.n10807 GND.n10773 9.3005
R25020 GND.n10804 GND.n10774 9.3005
R25021 GND.n10803 GND.n10775 9.3005
R25022 GND.n10800 GND.n10776 9.3005
R25023 GND.n10799 GND.n10777 9.3005
R25024 GND.n10796 GND.n10778 9.3005
R25025 GND.n10795 GND.n10779 9.3005
R25026 GND.n10792 GND.n10780 9.3005
R25027 GND.n10791 GND.n10781 9.3005
R25028 GND.n10788 GND.n10787 9.3005
R25029 GND.n10786 GND.n10783 9.3005
R25030 GND.n10719 GND.n10718 9.3005
R25031 GND.n5918 GND.n5875 9.3005
R25032 GND.n6742 GND.n5934 9.3005
R25033 GND.n7521 GND.n5935 9.3005
R25034 GND.n7520 GND.n5936 9.3005
R25035 GND.n7519 GND.n5937 9.3005
R25036 GND.n6757 GND.n5938 9.3005
R25037 GND.n7509 GND.n5955 9.3005
R25038 GND.n7508 GND.n5956 9.3005
R25039 GND.n7507 GND.n5957 9.3005
R25040 GND.n6772 GND.n5958 9.3005
R25041 GND.n7497 GND.n5976 9.3005
R25042 GND.n7496 GND.n5977 9.3005
R25043 GND.n7495 GND.n5978 9.3005
R25044 GND.n6787 GND.n5979 9.3005
R25045 GND.n7485 GND.n5997 9.3005
R25046 GND.n7484 GND.n5998 9.3005
R25047 GND.n7483 GND.n5999 9.3005
R25048 GND.n6802 GND.n6000 9.3005
R25049 GND.n7473 GND.n6018 9.3005
R25050 GND.n7472 GND.n6019 9.3005
R25051 GND.n7471 GND.n6020 9.3005
R25052 GND.n6817 GND.n6021 9.3005
R25053 GND.n7461 GND.n6038 9.3005
R25054 GND.n7460 GND.n6039 9.3005
R25055 GND.n7459 GND.n6040 9.3005
R25056 GND.n6832 GND.n6041 9.3005
R25057 GND.n7449 GND.n6059 9.3005
R25058 GND.n7448 GND.n6060 9.3005
R25059 GND.n7447 GND.n6061 9.3005
R25060 GND.n6847 GND.n6062 9.3005
R25061 GND.n7437 GND.n6080 9.3005
R25062 GND.n7436 GND.n6081 9.3005
R25063 GND.n7435 GND.n6082 9.3005
R25064 GND.n6862 GND.n6083 9.3005
R25065 GND.n7425 GND.n6101 9.3005
R25066 GND.n7424 GND.n6102 9.3005
R25067 GND.n7423 GND.n6103 9.3005
R25068 GND.n6877 GND.n6104 9.3005
R25069 GND.n7413 GND.n6122 9.3005
R25070 GND.n7412 GND.n6123 9.3005
R25071 GND.n7411 GND.n6124 9.3005
R25072 GND.n6892 GND.n6125 9.3005
R25073 GND.n7401 GND.n6143 9.3005
R25074 GND.n7400 GND.n6144 9.3005
R25075 GND.n7399 GND.n6145 9.3005
R25076 GND.n6907 GND.n6146 9.3005
R25077 GND.n7389 GND.n6164 9.3005
R25078 GND.n7388 GND.n6165 9.3005
R25079 GND.n7387 GND.n6166 9.3005
R25080 GND.n6922 GND.n6167 9.3005
R25081 GND.n7377 GND.n6184 9.3005
R25082 GND.n7376 GND.n6185 9.3005
R25083 GND.n7375 GND.n6186 9.3005
R25084 GND.n6937 GND.n6187 9.3005
R25085 GND.n7365 GND.n6205 9.3005
R25086 GND.n7364 GND.n6206 9.3005
R25087 GND.n7363 GND.n6207 9.3005
R25088 GND.n6952 GND.n6208 9.3005
R25089 GND.n7353 GND.n6226 9.3005
R25090 GND.n7352 GND.n6227 9.3005
R25091 GND.n7351 GND.n6228 9.3005
R25092 GND.n6967 GND.n6229 9.3005
R25093 GND.n7341 GND.n6246 9.3005
R25094 GND.n7340 GND.n6247 9.3005
R25095 GND.n7339 GND.n6248 9.3005
R25096 GND.n6990 GND.n6249 9.3005
R25097 GND.n6991 GND.n6469 9.3005
R25098 GND.n6997 GND.n6468 9.3005
R25099 GND.n6999 GND.n6998 9.3005
R25100 GND.n6465 GND.n6464 9.3005
R25101 GND.n7008 GND.n7007 9.3005
R25102 GND.n7009 GND.n117 9.3005
R25103 GND.n11102 GND.n118 9.3005
R25104 GND.n11101 GND.n119 9.3005
R25105 GND.n11100 GND.n120 9.3005
R25106 GND.n7014 GND.n121 9.3005
R25107 GND.n11090 GND.n137 9.3005
R25108 GND.n11089 GND.n138 9.3005
R25109 GND.n11088 GND.n139 9.3005
R25110 GND.n7029 GND.n140 9.3005
R25111 GND.n11078 GND.n158 9.3005
R25112 GND.n11077 GND.n159 9.3005
R25113 GND.n11076 GND.n160 9.3005
R25114 GND.n7044 GND.n161 9.3005
R25115 GND.n11066 GND.n179 9.3005
R25116 GND.n11065 GND.n180 9.3005
R25117 GND.n11064 GND.n181 9.3005
R25118 GND.n7059 GND.n182 9.3005
R25119 GND.n11054 GND.n200 9.3005
R25120 GND.n11053 GND.n201 9.3005
R25121 GND.n11052 GND.n202 9.3005
R25122 GND.n7074 GND.n203 9.3005
R25123 GND.n11042 GND.n221 9.3005
R25124 GND.n11041 GND.n222 9.3005
R25125 GND.n11040 GND.n223 9.3005
R25126 GND.n7089 GND.n224 9.3005
R25127 GND.n11030 GND.n242 9.3005
R25128 GND.n11029 GND.n243 9.3005
R25129 GND.n11028 GND.n244 9.3005
R25130 GND.n7105 GND.n245 9.3005
R25131 GND.n11018 GND.n262 9.3005
R25132 GND.n11017 GND.n263 9.3005
R25133 GND.n11016 GND.n264 9.3005
R25134 GND.n7108 GND.n265 9.3005
R25135 GND.n11006 GND.n283 9.3005
R25136 GND.n11005 GND.n284 9.3005
R25137 GND.n11004 GND.n285 9.3005
R25138 GND.n7115 GND.n286 9.3005
R25139 GND.n10994 GND.n304 9.3005
R25140 GND.n10993 GND.n305 9.3005
R25141 GND.n10992 GND.n306 9.3005
R25142 GND.n7122 GND.n307 9.3005
R25143 GND.n10982 GND.n325 9.3005
R25144 GND.n10981 GND.n326 9.3005
R25145 GND.n10980 GND.n327 9.3005
R25146 GND.n7129 GND.n328 9.3005
R25147 GND.n10970 GND.n346 9.3005
R25148 GND.n10969 GND.n347 9.3005
R25149 GND.n10968 GND.n348 9.3005
R25150 GND.n7136 GND.n349 9.3005
R25151 GND.n10958 GND.n367 9.3005
R25152 GND.n10957 GND.n368 9.3005
R25153 GND.n10956 GND.n369 9.3005
R25154 GND.n7143 GND.n370 9.3005
R25155 GND.n10946 GND.n388 9.3005
R25156 GND.n10945 GND.n389 9.3005
R25157 GND.n10944 GND.n390 9.3005
R25158 GND.n7150 GND.n391 9.3005
R25159 GND.n10934 GND.n409 9.3005
R25160 GND.n10933 GND.n410 9.3005
R25161 GND.n10932 GND.n411 9.3005
R25162 GND.n7157 GND.n412 9.3005
R25163 GND.n10922 GND.n430 9.3005
R25164 GND.n10921 GND.n431 9.3005
R25165 GND.n10920 GND.n432 9.3005
R25166 GND.n450 GND.n433 9.3005
R25167 GND.n10910 GND.n10909 9.3005
R25168 GND.n7535 GND.n5874 9.3005
R25169 GND.n5876 GND.n5875 9.3005
R25170 GND.n6743 GND.n6742 9.3005
R25171 GND.n6736 GND.n5935 9.3005
R25172 GND.n6755 GND.n5936 9.3005
R25173 GND.n6756 GND.n5937 9.3005
R25174 GND.n6758 GND.n6757 9.3005
R25175 GND.n6530 GND.n5955 9.3005
R25176 GND.n6770 GND.n5956 9.3005
R25177 GND.n6771 GND.n5957 9.3005
R25178 GND.n6773 GND.n6772 9.3005
R25179 GND.n6526 GND.n5976 9.3005
R25180 GND.n6785 GND.n5977 9.3005
R25181 GND.n6786 GND.n5978 9.3005
R25182 GND.n6788 GND.n6787 9.3005
R25183 GND.n6522 GND.n5997 9.3005
R25184 GND.n6800 GND.n5998 9.3005
R25185 GND.n6801 GND.n5999 9.3005
R25186 GND.n6803 GND.n6802 9.3005
R25187 GND.n6518 GND.n6018 9.3005
R25188 GND.n6815 GND.n6019 9.3005
R25189 GND.n6816 GND.n6020 9.3005
R25190 GND.n6818 GND.n6817 9.3005
R25191 GND.n6513 GND.n6038 9.3005
R25192 GND.n6830 GND.n6039 9.3005
R25193 GND.n6831 GND.n6040 9.3005
R25194 GND.n6833 GND.n6832 9.3005
R25195 GND.n6509 GND.n6059 9.3005
R25196 GND.n6845 GND.n6060 9.3005
R25197 GND.n6846 GND.n6061 9.3005
R25198 GND.n6848 GND.n6847 9.3005
R25199 GND.n6505 GND.n6080 9.3005
R25200 GND.n6860 GND.n6081 9.3005
R25201 GND.n6861 GND.n6082 9.3005
R25202 GND.n6863 GND.n6862 9.3005
R25203 GND.n6501 GND.n6101 9.3005
R25204 GND.n6875 GND.n6102 9.3005
R25205 GND.n6876 GND.n6103 9.3005
R25206 GND.n6878 GND.n6877 9.3005
R25207 GND.n6497 GND.n6122 9.3005
R25208 GND.n6890 GND.n6123 9.3005
R25209 GND.n6891 GND.n6124 9.3005
R25210 GND.n6893 GND.n6892 9.3005
R25211 GND.n6493 GND.n6143 9.3005
R25212 GND.n6905 GND.n6144 9.3005
R25213 GND.n6906 GND.n6145 9.3005
R25214 GND.n6908 GND.n6907 9.3005
R25215 GND.n6489 GND.n6164 9.3005
R25216 GND.n6920 GND.n6165 9.3005
R25217 GND.n6921 GND.n6166 9.3005
R25218 GND.n6923 GND.n6922 9.3005
R25219 GND.n6484 GND.n6184 9.3005
R25220 GND.n6935 GND.n6185 9.3005
R25221 GND.n6936 GND.n6186 9.3005
R25222 GND.n6938 GND.n6937 9.3005
R25223 GND.n6480 GND.n6205 9.3005
R25224 GND.n6950 GND.n6206 9.3005
R25225 GND.n6951 GND.n6207 9.3005
R25226 GND.n6953 GND.n6952 9.3005
R25227 GND.n6476 GND.n6226 9.3005
R25228 GND.n6965 GND.n6227 9.3005
R25229 GND.n6966 GND.n6228 9.3005
R25230 GND.n6968 GND.n6967 9.3005
R25231 GND.n6472 GND.n6246 9.3005
R25232 GND.n6987 GND.n6247 9.3005
R25233 GND.n6988 GND.n6248 9.3005
R25234 GND.n6990 GND.n6989 9.3005
R25235 GND.n6992 GND.n6991 9.3005
R25236 GND.n6468 GND.n6467 9.3005
R25237 GND.n7000 GND.n6999 9.3005
R25238 GND.n7001 GND.n6464 9.3005
R25239 GND.n7008 GND.n6463 9.3005
R25240 GND.n7010 GND.n7009 9.3005
R25241 GND.n7011 GND.n118 9.3005
R25242 GND.n7012 GND.n119 9.3005
R25243 GND.n7013 GND.n120 9.3005
R25244 GND.n7015 GND.n7014 9.3005
R25245 GND.n6460 GND.n137 9.3005
R25246 GND.n7027 GND.n138 9.3005
R25247 GND.n7028 GND.n139 9.3005
R25248 GND.n7030 GND.n7029 9.3005
R25249 GND.n6456 GND.n158 9.3005
R25250 GND.n7042 GND.n159 9.3005
R25251 GND.n7043 GND.n160 9.3005
R25252 GND.n7045 GND.n7044 9.3005
R25253 GND.n6452 GND.n179 9.3005
R25254 GND.n7057 GND.n180 9.3005
R25255 GND.n7058 GND.n181 9.3005
R25256 GND.n7060 GND.n7059 9.3005
R25257 GND.n6448 GND.n200 9.3005
R25258 GND.n7072 GND.n201 9.3005
R25259 GND.n7073 GND.n202 9.3005
R25260 GND.n7075 GND.n7074 9.3005
R25261 GND.n6444 GND.n221 9.3005
R25262 GND.n7087 GND.n222 9.3005
R25263 GND.n7088 GND.n223 9.3005
R25264 GND.n7090 GND.n7089 9.3005
R25265 GND.n6440 GND.n242 9.3005
R25266 GND.n7103 GND.n243 9.3005
R25267 GND.n7104 GND.n244 9.3005
R25268 GND.n7106 GND.n7105 9.3005
R25269 GND.n7107 GND.n262 9.3005
R25270 GND.n7260 GND.n263 9.3005
R25271 GND.n7259 GND.n264 9.3005
R25272 GND.n7258 GND.n7108 9.3005
R25273 GND.n7109 GND.n283 9.3005
R25274 GND.n7248 GND.n284 9.3005
R25275 GND.n7247 GND.n285 9.3005
R25276 GND.n7246 GND.n7115 9.3005
R25277 GND.n7116 GND.n304 9.3005
R25278 GND.n7236 GND.n305 9.3005
R25279 GND.n7235 GND.n306 9.3005
R25280 GND.n7234 GND.n7122 9.3005
R25281 GND.n7123 GND.n325 9.3005
R25282 GND.n7224 GND.n326 9.3005
R25283 GND.n7223 GND.n327 9.3005
R25284 GND.n7222 GND.n7129 9.3005
R25285 GND.n7130 GND.n346 9.3005
R25286 GND.n7212 GND.n347 9.3005
R25287 GND.n7211 GND.n348 9.3005
R25288 GND.n7210 GND.n7136 9.3005
R25289 GND.n7137 GND.n367 9.3005
R25290 GND.n7200 GND.n368 9.3005
R25291 GND.n7199 GND.n369 9.3005
R25292 GND.n7198 GND.n7143 9.3005
R25293 GND.n7144 GND.n388 9.3005
R25294 GND.n7188 GND.n389 9.3005
R25295 GND.n7187 GND.n390 9.3005
R25296 GND.n7186 GND.n7150 9.3005
R25297 GND.n7151 GND.n409 9.3005
R25298 GND.n7176 GND.n410 9.3005
R25299 GND.n7175 GND.n411 9.3005
R25300 GND.n7174 GND.n7157 9.3005
R25301 GND.n7158 GND.n430 9.3005
R25302 GND.n7164 GND.n431 9.3005
R25303 GND.n452 GND.n432 9.3005
R25304 GND.n10907 GND.n450 9.3005
R25305 GND.n10909 GND.n10908 9.3005
R25306 GND.n7535 GND.n7534 9.3005
R25307 GND.n7539 GND.n7538 9.3005
R25308 GND.n7542 GND.n4826 9.3005
R25309 GND.n7543 GND.n4825 9.3005
R25310 GND.n7546 GND.n4824 9.3005
R25311 GND.n7547 GND.n4823 9.3005
R25312 GND.n7550 GND.n4822 9.3005
R25313 GND.n7551 GND.n4821 9.3005
R25314 GND.n7554 GND.n4820 9.3005
R25315 GND.n7555 GND.n4819 9.3005
R25316 GND.n7558 GND.n4818 9.3005
R25317 GND.n7559 GND.n4817 9.3005
R25318 GND.n7562 GND.n4816 9.3005
R25319 GND.n7563 GND.n4815 9.3005
R25320 GND.n7566 GND.n4814 9.3005
R25321 GND.n7567 GND.n4813 9.3005
R25322 GND.n7570 GND.n4809 9.3005
R25323 GND.n7571 GND.n4808 9.3005
R25324 GND.n7574 GND.n4807 9.3005
R25325 GND.n7575 GND.n4806 9.3005
R25326 GND.n7578 GND.n4805 9.3005
R25327 GND.n7579 GND.n4804 9.3005
R25328 GND.n7582 GND.n4803 9.3005
R25329 GND.n7583 GND.n4802 9.3005
R25330 GND.n7586 GND.n4801 9.3005
R25331 GND.n7587 GND.n4800 9.3005
R25332 GND.n7590 GND.n4799 9.3005
R25333 GND.n7591 GND.n4798 9.3005
R25334 GND.n7594 GND.n4797 9.3005
R25335 GND.n7596 GND.n4796 9.3005
R25336 GND.n7600 GND.n4633 9.3005
R25337 GND.n7601 GND.n4632 9.3005
R25338 GND.n7604 GND.n4631 9.3005
R25339 GND.n7605 GND.n4630 9.3005
R25340 GND.n7608 GND.n4629 9.3005
R25341 GND.n7609 GND.n4628 9.3005
R25342 GND.n7612 GND.n4627 9.3005
R25343 GND.n7613 GND.n4626 9.3005
R25344 GND.n7616 GND.n4625 9.3005
R25345 GND.n7617 GND.n4624 9.3005
R25346 GND.n7620 GND.n4623 9.3005
R25347 GND.n7622 GND.n4622 9.3005
R25348 GND.n7624 GND.n4617 9.3005
R25349 GND.n7627 GND.n4616 9.3005
R25350 GND.n7628 GND.n4615 9.3005
R25351 GND.n7631 GND.n4614 9.3005
R25352 GND.n7632 GND.n4613 9.3005
R25353 GND.n7635 GND.n4612 9.3005
R25354 GND.n7636 GND.n4611 9.3005
R25355 GND.n7639 GND.n4610 9.3005
R25356 GND.n7641 GND.n4609 9.3005
R25357 GND.n7642 GND.n4608 9.3005
R25358 GND.n7643 GND.n4607 9.3005
R25359 GND.n7644 GND.n4606 9.3005
R25360 GND.n7623 GND.n4619 9.3005
R25361 GND.n7537 GND.n4827 9.3005
R25362 GND.n7527 GND.n5924 9.3005
R25363 GND.n7526 GND.n5925 9.3005
R25364 GND.n7525 GND.n5926 9.3005
R25365 GND.n5945 GND.n5927 9.3005
R25366 GND.n7515 GND.n5946 9.3005
R25367 GND.n7514 GND.n5947 9.3005
R25368 GND.n7513 GND.n5948 9.3005
R25369 GND.n5965 GND.n5949 9.3005
R25370 GND.n7503 GND.n5966 9.3005
R25371 GND.n7502 GND.n5967 9.3005
R25372 GND.n7501 GND.n5968 9.3005
R25373 GND.n5986 GND.n5969 9.3005
R25374 GND.n7491 GND.n5987 9.3005
R25375 GND.n7490 GND.n5988 9.3005
R25376 GND.n7489 GND.n5989 9.3005
R25377 GND.n6007 GND.n5990 9.3005
R25378 GND.n7479 GND.n6008 9.3005
R25379 GND.n7478 GND.n6009 9.3005
R25380 GND.n7477 GND.n6010 9.3005
R25381 GND.n6028 GND.n6011 9.3005
R25382 GND.n7467 GND.n6029 9.3005
R25383 GND.n7466 GND.n6030 9.3005
R25384 GND.n7465 GND.n6031 9.3005
R25385 GND.n6048 GND.n6032 9.3005
R25386 GND.n7455 GND.n6049 9.3005
R25387 GND.n7454 GND.n6050 9.3005
R25388 GND.n7453 GND.n6051 9.3005
R25389 GND.n6069 GND.n6052 9.3005
R25390 GND.n7443 GND.n6070 9.3005
R25391 GND.n7442 GND.n6071 9.3005
R25392 GND.n7441 GND.n6072 9.3005
R25393 GND.n6090 GND.n6073 9.3005
R25394 GND.n7431 GND.n6091 9.3005
R25395 GND.n7430 GND.n6092 9.3005
R25396 GND.n7429 GND.n6093 9.3005
R25397 GND.n6111 GND.n6094 9.3005
R25398 GND.n7419 GND.n6112 9.3005
R25399 GND.n7418 GND.n6113 9.3005
R25400 GND.n7417 GND.n6114 9.3005
R25401 GND.n6132 GND.n6115 9.3005
R25402 GND.n7407 GND.n6133 9.3005
R25403 GND.n7406 GND.n6134 9.3005
R25404 GND.n7405 GND.n6135 9.3005
R25405 GND.n6153 GND.n6136 9.3005
R25406 GND.n7395 GND.n6154 9.3005
R25407 GND.n7394 GND.n6155 9.3005
R25408 GND.n7393 GND.n6156 9.3005
R25409 GND.n6173 GND.n6157 9.3005
R25410 GND.n7383 GND.n6174 9.3005
R25411 GND.n7382 GND.n6175 9.3005
R25412 GND.n7381 GND.n6176 9.3005
R25413 GND.n6194 GND.n6177 9.3005
R25414 GND.n7371 GND.n6195 9.3005
R25415 GND.n7370 GND.n6196 9.3005
R25416 GND.n7369 GND.n6197 9.3005
R25417 GND.n6215 GND.n6198 9.3005
R25418 GND.n7359 GND.n6216 9.3005
R25419 GND.n7358 GND.n6217 9.3005
R25420 GND.n7357 GND.n6218 9.3005
R25421 GND.n6236 GND.n6219 9.3005
R25422 GND.n7347 GND.n6237 9.3005
R25423 GND.n7346 GND.n6238 9.3005
R25424 GND.n7345 GND.n101 9.3005
R25425 GND.n108 GND.n100 9.3005
R25426 GND.n11096 GND.n127 9.3005
R25427 GND.n11095 GND.n128 9.3005
R25428 GND.n11094 GND.n129 9.3005
R25429 GND.n147 GND.n130 9.3005
R25430 GND.n11084 GND.n148 9.3005
R25431 GND.n11083 GND.n149 9.3005
R25432 GND.n11082 GND.n150 9.3005
R25433 GND.n168 GND.n151 9.3005
R25434 GND.n11072 GND.n169 9.3005
R25435 GND.n11071 GND.n170 9.3005
R25436 GND.n11070 GND.n171 9.3005
R25437 GND.n189 GND.n172 9.3005
R25438 GND.n11060 GND.n190 9.3005
R25439 GND.n11059 GND.n191 9.3005
R25440 GND.n11058 GND.n192 9.3005
R25441 GND.n210 GND.n193 9.3005
R25442 GND.n11048 GND.n211 9.3005
R25443 GND.n11047 GND.n212 9.3005
R25444 GND.n11046 GND.n213 9.3005
R25445 GND.n231 GND.n214 9.3005
R25446 GND.n11036 GND.n232 9.3005
R25447 GND.n11035 GND.n233 9.3005
R25448 GND.n11034 GND.n234 9.3005
R25449 GND.n252 GND.n235 9.3005
R25450 GND.n11024 GND.n253 9.3005
R25451 GND.n11023 GND.n254 9.3005
R25452 GND.n11022 GND.n255 9.3005
R25453 GND.n272 GND.n256 9.3005
R25454 GND.n11012 GND.n273 9.3005
R25455 GND.n11011 GND.n274 9.3005
R25456 GND.n11010 GND.n275 9.3005
R25457 GND.n293 GND.n276 9.3005
R25458 GND.n11000 GND.n294 9.3005
R25459 GND.n10999 GND.n295 9.3005
R25460 GND.n10998 GND.n296 9.3005
R25461 GND.n314 GND.n297 9.3005
R25462 GND.n10988 GND.n315 9.3005
R25463 GND.n10987 GND.n316 9.3005
R25464 GND.n10986 GND.n317 9.3005
R25465 GND.n335 GND.n318 9.3005
R25466 GND.n10976 GND.n336 9.3005
R25467 GND.n10975 GND.n337 9.3005
R25468 GND.n10974 GND.n338 9.3005
R25469 GND.n356 GND.n339 9.3005
R25470 GND.n10964 GND.n357 9.3005
R25471 GND.n10963 GND.n358 9.3005
R25472 GND.n10962 GND.n359 9.3005
R25473 GND.n377 GND.n360 9.3005
R25474 GND.n10952 GND.n378 9.3005
R25475 GND.n10951 GND.n379 9.3005
R25476 GND.n10950 GND.n380 9.3005
R25477 GND.n398 GND.n381 9.3005
R25478 GND.n10940 GND.n399 9.3005
R25479 GND.n10939 GND.n400 9.3005
R25480 GND.n10938 GND.n401 9.3005
R25481 GND.n419 GND.n402 9.3005
R25482 GND.n10928 GND.n420 9.3005
R25483 GND.n10927 GND.n421 9.3005
R25484 GND.n10926 GND.n422 9.3005
R25485 GND.n440 GND.n423 9.3005
R25486 GND.n10916 GND.n441 9.3005
R25487 GND.n10915 GND.n442 9.3005
R25488 GND.n10914 GND.n443 9.3005
R25489 GND.n5923 GND.n5922 9.3005
R25490 GND.n11107 GND.n105 9.3005
R25491 GND.n11107 GND.n11106 9.3005
R25492 GND.n8706 GND.n8705 9.3005
R25493 GND.n8709 GND.n1792 9.3005
R25494 GND.n8710 GND.n1791 9.3005
R25495 GND.n8713 GND.n1790 9.3005
R25496 GND.n8714 GND.n1789 9.3005
R25497 GND.n8717 GND.n1788 9.3005
R25498 GND.n8718 GND.n1787 9.3005
R25499 GND.n8721 GND.n1786 9.3005
R25500 GND.n8722 GND.n1785 9.3005
R25501 GND.n8725 GND.n1784 9.3005
R25502 GND.n8726 GND.n1783 9.3005
R25503 GND.n8729 GND.n1782 9.3005
R25504 GND.n8730 GND.n1781 9.3005
R25505 GND.n8733 GND.n1780 9.3005
R25506 GND.n8734 GND.n1779 9.3005
R25507 GND.n8737 GND.n1775 9.3005
R25508 GND.n8738 GND.n1774 9.3005
R25509 GND.n8741 GND.n1773 9.3005
R25510 GND.n8742 GND.n1772 9.3005
R25511 GND.n8745 GND.n1771 9.3005
R25512 GND.n8746 GND.n1770 9.3005
R25513 GND.n8749 GND.n1769 9.3005
R25514 GND.n8750 GND.n1768 9.3005
R25515 GND.n8753 GND.n1767 9.3005
R25516 GND.n8754 GND.n1766 9.3005
R25517 GND.n8757 GND.n1765 9.3005
R25518 GND.n8758 GND.n1764 9.3005
R25519 GND.n8761 GND.n1763 9.3005
R25520 GND.n8762 GND.n1762 9.3005
R25521 GND.n8766 GND.n1757 9.3005
R25522 GND.n8769 GND.n1756 9.3005
R25523 GND.n8770 GND.n1755 9.3005
R25524 GND.n8773 GND.n1754 9.3005
R25525 GND.n8774 GND.n1753 9.3005
R25526 GND.n8777 GND.n1752 9.3005
R25527 GND.n8778 GND.n1751 9.3005
R25528 GND.n8781 GND.n1750 9.3005
R25529 GND.n8782 GND.n1749 9.3005
R25530 GND.n8785 GND.n1748 9.3005
R25531 GND.n8786 GND.n1747 9.3005
R25532 GND.n8789 GND.n1746 9.3005
R25533 GND.n8791 GND.n1745 9.3005
R25534 GND.n8793 GND.n1740 9.3005
R25535 GND.n8796 GND.n1739 9.3005
R25536 GND.n8797 GND.n1738 9.3005
R25537 GND.n8800 GND.n1737 9.3005
R25538 GND.n8801 GND.n1736 9.3005
R25539 GND.n8804 GND.n1735 9.3005
R25540 GND.n8805 GND.n1734 9.3005
R25541 GND.n8808 GND.n1733 9.3005
R25542 GND.n8810 GND.n1732 9.3005
R25543 GND.n8811 GND.n1731 9.3005
R25544 GND.n8812 GND.n1730 9.3005
R25545 GND.n8813 GND.n1729 9.3005
R25546 GND.n8792 GND.n1742 9.3005
R25547 GND.n8765 GND.n1758 9.3005
R25548 GND.n8704 GND.n1793 9.3005
R25549 GND.n1829 GND.n1828 9.3005
R25550 GND.n1830 GND.n1824 9.3005
R25551 GND.n8688 GND.n1831 9.3005
R25552 GND.n8687 GND.n1832 9.3005
R25553 GND.n8686 GND.n1833 9.3005
R25554 GND.n3154 GND.n1834 9.3005
R25555 GND.n3158 GND.n3155 9.3005
R25556 GND.n3157 GND.n3156 9.3005
R25557 GND.n2895 GND.n2894 9.3005
R25558 GND.n3178 GND.n3177 9.3005
R25559 GND.n3179 GND.n2893 9.3005
R25560 GND.n3183 GND.n3180 9.3005
R25561 GND.n3182 GND.n3181 9.3005
R25562 GND.n2872 GND.n2871 9.3005
R25563 GND.n3203 GND.n3202 9.3005
R25564 GND.n3204 GND.n2870 9.3005
R25565 GND.n3208 GND.n3205 9.3005
R25566 GND.n3207 GND.n3206 9.3005
R25567 GND.n2849 GND.n2848 9.3005
R25568 GND.n3227 GND.n3226 9.3005
R25569 GND.n3228 GND.n2847 9.3005
R25570 GND.n3232 GND.n3229 9.3005
R25571 GND.n3231 GND.n3230 9.3005
R25572 GND.n2826 GND.n2825 9.3005
R25573 GND.n3252 GND.n3251 9.3005
R25574 GND.n3253 GND.n2824 9.3005
R25575 GND.n3257 GND.n3254 9.3005
R25576 GND.n3256 GND.n3255 9.3005
R25577 GND.n2804 GND.n2803 9.3005
R25578 GND.n3277 GND.n3276 9.3005
R25579 GND.n3278 GND.n2802 9.3005
R25580 GND.n3282 GND.n3279 9.3005
R25581 GND.n3281 GND.n3280 9.3005
R25582 GND.n2781 GND.n2780 9.3005
R25583 GND.n3302 GND.n3301 9.3005
R25584 GND.n3303 GND.n2779 9.3005
R25585 GND.n3307 GND.n3304 9.3005
R25586 GND.n3306 GND.n3305 9.3005
R25587 GND.n2758 GND.n2757 9.3005
R25588 GND.n3326 GND.n3325 9.3005
R25589 GND.n3327 GND.n2756 9.3005
R25590 GND.n3331 GND.n3328 9.3005
R25591 GND.n3330 GND.n3329 9.3005
R25592 GND.n2735 GND.n2734 9.3005
R25593 GND.n3351 GND.n3350 9.3005
R25594 GND.n3352 GND.n2733 9.3005
R25595 GND.n3356 GND.n3353 9.3005
R25596 GND.n3355 GND.n3354 9.3005
R25597 GND.n2713 GND.n2712 9.3005
R25598 GND.n3376 GND.n3375 9.3005
R25599 GND.n3377 GND.n2711 9.3005
R25600 GND.n3381 GND.n3378 9.3005
R25601 GND.n3380 GND.n3379 9.3005
R25602 GND.n2690 GND.n2689 9.3005
R25603 GND.n3401 GND.n3400 9.3005
R25604 GND.n3402 GND.n2688 9.3005
R25605 GND.n3406 GND.n3403 9.3005
R25606 GND.n3405 GND.n3404 9.3005
R25607 GND.n2667 GND.n2666 9.3005
R25608 GND.n3425 GND.n3424 9.3005
R25609 GND.n3426 GND.n2665 9.3005
R25610 GND.n3428 GND.n3427 9.3005
R25611 GND.n2498 GND.n2491 9.3005
R25612 GND.n3498 GND.n3495 9.3005
R25613 GND.n3497 GND.n3496 9.3005
R25614 GND.n2470 GND.n2469 9.3005
R25615 GND.n3519 GND.n3518 9.3005
R25616 GND.n3520 GND.n2468 9.3005
R25617 GND.n3524 GND.n3521 9.3005
R25618 GND.n3523 GND.n3522 9.3005
R25619 GND.n2449 GND.n2448 9.3005
R25620 GND.n3545 GND.n3544 9.3005
R25621 GND.n3546 GND.n2447 9.3005
R25622 GND.n3550 GND.n3547 9.3005
R25623 GND.n3549 GND.n3548 9.3005
R25624 GND.n2427 GND.n2426 9.3005
R25625 GND.n3571 GND.n3570 9.3005
R25626 GND.n3572 GND.n2425 9.3005
R25627 GND.n3576 GND.n3573 9.3005
R25628 GND.n3575 GND.n3574 9.3005
R25629 GND.n2405 GND.n2404 9.3005
R25630 GND.n3596 GND.n3595 9.3005
R25631 GND.n3597 GND.n2403 9.3005
R25632 GND.n3601 GND.n3598 9.3005
R25633 GND.n3600 GND.n3599 9.3005
R25634 GND.n2383 GND.n2382 9.3005
R25635 GND.n3622 GND.n3621 9.3005
R25636 GND.n3623 GND.n2381 9.3005
R25637 GND.n3627 GND.n3624 9.3005
R25638 GND.n3626 GND.n3625 9.3005
R25639 GND.n2365 GND.n2364 9.3005
R25640 GND.n3648 GND.n3647 9.3005
R25641 GND.n3649 GND.n2363 9.3005
R25642 GND.n3653 GND.n3650 9.3005
R25643 GND.n3652 GND.n3651 9.3005
R25644 GND.n2343 GND.n2342 9.3005
R25645 GND.n3674 GND.n3673 9.3005
R25646 GND.n3675 GND.n2341 9.3005
R25647 GND.n3679 GND.n3676 9.3005
R25648 GND.n3678 GND.n3677 9.3005
R25649 GND.n2315 GND.n2314 9.3005
R25650 GND.n8185 GND.n8184 9.3005
R25651 GND.n8186 GND.n2313 9.3005
R25652 GND.n8190 GND.n8187 9.3005
R25653 GND.n8189 GND.n8188 9.3005
R25654 GND.n2294 GND.n2293 9.3005
R25655 GND.n8211 GND.n8210 9.3005
R25656 GND.n8212 GND.n2292 9.3005
R25657 GND.n8216 GND.n8213 9.3005
R25658 GND.n8215 GND.n8214 9.3005
R25659 GND.n2273 GND.n2272 9.3005
R25660 GND.n8237 GND.n8236 9.3005
R25661 GND.n8238 GND.n2271 9.3005
R25662 GND.n8242 GND.n8239 9.3005
R25663 GND.n8241 GND.n8240 9.3005
R25664 GND.n2251 GND.n2250 9.3005
R25665 GND.n8263 GND.n8262 9.3005
R25666 GND.n8264 GND.n2249 9.3005
R25667 GND.n8268 GND.n8265 9.3005
R25668 GND.n8267 GND.n8266 9.3005
R25669 GND.n2229 GND.n2228 9.3005
R25670 GND.n8288 GND.n8287 9.3005
R25671 GND.n8289 GND.n2227 9.3005
R25672 GND.n8292 GND.n8291 9.3005
R25673 GND.n8290 GND.n2212 9.3005
R25674 GND.n8306 GND.n2211 9.3005
R25675 GND.n8308 GND.n8307 9.3005
R25676 GND.n1826 GND.n1825 9.3005
R25677 GND.n3494 GND.n2496 9.3005
R25678 GND.n3494 GND.n2490 9.3005
R25679 GND.n3484 GND.n2492 9.3005
R25680 GND.n2646 GND.n2538 9.3005
R25681 GND.n2645 GND.n2539 9.3005
R25682 GND.n2542 GND.n2540 9.3005
R25683 GND.n2641 GND.n2543 9.3005
R25684 GND.n2640 GND.n2544 9.3005
R25685 GND.n2639 GND.n2545 9.3005
R25686 GND.n2548 GND.n2546 9.3005
R25687 GND.n2635 GND.n2549 9.3005
R25688 GND.n2634 GND.n2550 9.3005
R25689 GND.n2633 GND.n2551 9.3005
R25690 GND.n2554 GND.n2552 9.3005
R25691 GND.n2629 GND.n2555 9.3005
R25692 GND.n2628 GND.n2556 9.3005
R25693 GND.n2627 GND.n2557 9.3005
R25694 GND.n2560 GND.n2558 9.3005
R25695 GND.n2623 GND.n2561 9.3005
R25696 GND.n2622 GND.n2562 9.3005
R25697 GND.n2621 GND.n2563 9.3005
R25698 GND.n2566 GND.n2564 9.3005
R25699 GND.n2617 GND.n2567 9.3005
R25700 GND.n2616 GND.n2568 9.3005
R25701 GND.n2615 GND.n2569 9.3005
R25702 GND.n2572 GND.n2570 9.3005
R25703 GND.n2611 GND.n2573 9.3005
R25704 GND.n2610 GND.n2574 9.3005
R25705 GND.n2609 GND.n2575 9.3005
R25706 GND.n2578 GND.n2576 9.3005
R25707 GND.n2602 GND.n2579 9.3005
R25708 GND.n2601 GND.n2580 9.3005
R25709 GND.n2600 GND.n2581 9.3005
R25710 GND.n2584 GND.n2582 9.3005
R25711 GND.n2596 GND.n2585 9.3005
R25712 GND.n2595 GND.n2586 9.3005
R25713 GND.n2594 GND.n2587 9.3005
R25714 GND.n2591 GND.n2588 9.3005
R25715 GND.n2590 GND.n2589 9.3005
R25716 GND.n2326 GND.n2325 9.3005
R25717 GND.n3696 GND.n3695 9.3005
R25718 GND.n3697 GND.n2324 9.3005
R25719 GND.n8176 GND.n3698 9.3005
R25720 GND.n8175 GND.n3699 9.3005
R25721 GND.n8174 GND.n3700 9.3005
R25722 GND.n3703 GND.n3701 9.3005
R25723 GND.n8170 GND.n3704 9.3005
R25724 GND.n8169 GND.n3705 9.3005
R25725 GND.n8168 GND.n3706 9.3005
R25726 GND.n3709 GND.n3707 9.3005
R25727 GND.n8164 GND.n3710 9.3005
R25728 GND.n8163 GND.n3711 9.3005
R25729 GND.n8162 GND.n3712 9.3005
R25730 GND.n3715 GND.n3713 9.3005
R25731 GND.n8158 GND.n3716 9.3005
R25732 GND.n8157 GND.n3717 9.3005
R25733 GND.n8156 GND.n3718 9.3005
R25734 GND.n3721 GND.n3719 9.3005
R25735 GND.n8152 GND.n3722 9.3005
R25736 GND.n8151 GND.n3723 9.3005
R25737 GND.n8150 GND.n3724 9.3005
R25738 GND.n3727 GND.n3725 9.3005
R25739 GND.n8146 GND.n3728 9.3005
R25740 GND.n8145 GND.n3729 9.3005
R25741 GND.n8144 GND.n3730 9.3005
R25742 GND.n3733 GND.n3731 9.3005
R25743 GND.n8140 GND.n3734 9.3005
R25744 GND.n8139 GND.n3735 9.3005
R25745 GND.n8138 GND.n3736 9.3005
R25746 GND.n3742 GND.n3737 9.3005
R25747 GND.n3743 GND.n3741 9.3005
R25748 GND.n8131 GND.n3744 9.3005
R25749 GND.n8130 GND.n3745 9.3005
R25750 GND.n8129 GND.n3746 9.3005
R25751 GND.n3774 GND.n3747 9.3005
R25752 GND.n8117 GND.n3775 9.3005
R25753 GND.n8116 GND.n3776 9.3005
R25754 GND.n8115 GND.n3777 9.3005
R25755 GND.n3790 GND.n3778 9.3005
R25756 GND.n8103 GND.n3791 9.3005
R25757 GND.n8102 GND.n3792 9.3005
R25758 GND.n8101 GND.n3793 9.3005
R25759 GND.n3808 GND.n3794 9.3005
R25760 GND.n8089 GND.n3809 9.3005
R25761 GND.n8088 GND.n3810 9.3005
R25762 GND.n8087 GND.n3811 9.3005
R25763 GND.n3826 GND.n3812 9.3005
R25764 GND.n8075 GND.n3827 9.3005
R25765 GND.n8074 GND.n3828 9.3005
R25766 GND.n8073 GND.n3829 9.3005
R25767 GND.n3844 GND.n3830 9.3005
R25768 GND.n8061 GND.n3845 9.3005
R25769 GND.n8060 GND.n3846 9.3005
R25770 GND.n8059 GND.n3847 9.3005
R25771 GND.n3887 GND.n3848 9.3005
R25772 GND.n8003 GND.n3888 9.3005
R25773 GND.n8002 GND.n3889 9.3005
R25774 GND.n8001 GND.n3890 9.3005
R25775 GND.n3908 GND.n3891 9.3005
R25776 GND.n7991 GND.n3909 9.3005
R25777 GND.n7990 GND.n3910 9.3005
R25778 GND.n7989 GND.n3911 9.3005
R25779 GND.n3928 GND.n3912 9.3005
R25780 GND.n7979 GND.n3929 9.3005
R25781 GND.n7978 GND.n3930 9.3005
R25782 GND.n7977 GND.n3931 9.3005
R25783 GND.n3948 GND.n3932 9.3005
R25784 GND.n7967 GND.n3949 9.3005
R25785 GND.n7966 GND.n3950 9.3005
R25786 GND.n7965 GND.n3951 9.3005
R25787 GND.n3968 GND.n3952 9.3005
R25788 GND.n7955 GND.n3969 9.3005
R25789 GND.n7954 GND.n3970 9.3005
R25790 GND.n7953 GND.n3971 9.3005
R25791 GND.n3988 GND.n3972 9.3005
R25792 GND.n7943 GND.n3989 9.3005
R25793 GND.n7942 GND.n3990 9.3005
R25794 GND.n7941 GND.n3991 9.3005
R25795 GND.n4008 GND.n3992 9.3005
R25796 GND.n7931 GND.n4009 9.3005
R25797 GND.n7930 GND.n4010 9.3005
R25798 GND.n7929 GND.n4011 9.3005
R25799 GND.n4028 GND.n4012 9.3005
R25800 GND.n7919 GND.n4029 9.3005
R25801 GND.n7918 GND.n4030 9.3005
R25802 GND.n7917 GND.n4031 9.3005
R25803 GND.n4048 GND.n4032 9.3005
R25804 GND.n7907 GND.n4049 9.3005
R25805 GND.n7906 GND.n4050 9.3005
R25806 GND.n7905 GND.n4051 9.3005
R25807 GND.n4079 GND.n4052 9.3005
R25808 GND.n4080 GND.n4078 9.3005
R25809 GND.n7888 GND.n4081 9.3005
R25810 GND.n7887 GND.n4082 9.3005
R25811 GND.n7886 GND.n4083 9.3005
R25812 GND.n4113 GND.n4084 9.3005
R25813 GND.n7876 GND.n4114 9.3005
R25814 GND.n7875 GND.n4115 9.3005
R25815 GND.n7874 GND.n4116 9.3005
R25816 GND.n4133 GND.n4117 9.3005
R25817 GND.n7864 GND.n4134 9.3005
R25818 GND.n7863 GND.n4135 9.3005
R25819 GND.n7862 GND.n4136 9.3005
R25820 GND.n4153 GND.n4137 9.3005
R25821 GND.n7852 GND.n4154 9.3005
R25822 GND.n7851 GND.n4155 9.3005
R25823 GND.n7850 GND.n4156 9.3005
R25824 GND.n4184 GND.n4157 9.3005
R25825 GND.n4185 GND.n4183 9.3005
R25826 GND.n7833 GND.n4186 9.3005
R25827 GND.n7832 GND.n4187 9.3005
R25828 GND.n7831 GND.n4188 9.3005
R25829 GND.n4217 GND.n4189 9.3005
R25830 GND.n7821 GND.n4218 9.3005
R25831 GND.n7820 GND.n4219 9.3005
R25832 GND.n7819 GND.n4220 9.3005
R25833 GND.n4237 GND.n4221 9.3005
R25834 GND.n7809 GND.n4238 9.3005
R25835 GND.n7808 GND.n4239 9.3005
R25836 GND.n7807 GND.n4240 9.3005
R25837 GND.n4255 GND.n4241 9.3005
R25838 GND.n7797 GND.n4256 9.3005
R25839 GND.n7796 GND.n4257 9.3005
R25840 GND.n7795 GND.n4258 9.3005
R25841 GND.n4286 GND.n4259 9.3005
R25842 GND.n4287 GND.n4285 9.3005
R25843 GND.n7778 GND.n4288 9.3005
R25844 GND.n7777 GND.n4289 9.3005
R25845 GND.n7776 GND.n4290 9.3005
R25846 GND.n4320 GND.n4291 9.3005
R25847 GND.n7766 GND.n4321 9.3005
R25848 GND.n7765 GND.n4322 9.3005
R25849 GND.n7764 GND.n4323 9.3005
R25850 GND.n4340 GND.n4324 9.3005
R25851 GND.n7754 GND.n4341 9.3005
R25852 GND.n7753 GND.n4342 9.3005
R25853 GND.n7752 GND.n4343 9.3005
R25854 GND.n4359 GND.n4344 9.3005
R25855 GND.n7742 GND.n4360 9.3005
R25856 GND.n7741 GND.n4361 9.3005
R25857 GND.n7740 GND.n4362 9.3005
R25858 GND.n4389 GND.n4363 9.3005
R25859 GND.n4390 GND.n4388 9.3005
R25860 GND.n7723 GND.n4391 9.3005
R25861 GND.n7722 GND.n4392 9.3005
R25862 GND.n7721 GND.n4393 9.3005
R25863 GND.n4408 GND.n4394 9.3005
R25864 GND.n7709 GND.n4409 9.3005
R25865 GND.n7708 GND.n4410 9.3005
R25866 GND.n7707 GND.n4411 9.3005
R25867 GND.n4426 GND.n4412 9.3005
R25868 GND.n7695 GND.n4427 9.3005
R25869 GND.n7694 GND.n4428 9.3005
R25870 GND.n7693 GND.n4429 9.3005
R25871 GND.n4443 GND.n4430 9.3005
R25872 GND.n7681 GND.n4444 9.3005
R25873 GND.n7680 GND.n4445 9.3005
R25874 GND.n7679 GND.n4446 9.3005
R25875 GND.n4520 GND.n4447 9.3005
R25876 GND.n4521 GND.n4519 9.3005
R25877 GND.n7662 GND.n4522 9.3005
R25878 GND.n7661 GND.n4523 9.3005
R25879 GND.n7660 GND.n4524 9.3005
R25880 GND.n4562 GND.n4525 9.3005
R25881 GND.n7653 GND.n4563 9.3005
R25882 GND.n7652 GND.n4564 9.3005
R25883 GND.n7651 GND.n4565 9.3005
R25884 GND.n6542 GND.n4566 9.3005
R25885 GND.n6543 GND.n6541 9.3005
R25886 GND.n6545 GND.n6544 9.3005
R25887 GND.n6539 GND.n6538 9.3005
R25888 GND.n6550 GND.n6549 9.3005
R25889 GND.n6551 GND.n6537 9.3005
R25890 GND.n6553 GND.n6552 9.3005
R25891 GND.n6535 GND.n6534 9.3005
R25892 GND.n6558 GND.n6557 9.3005
R25893 GND.n6559 GND.n6533 9.3005
R25894 GND.n6730 GND.n6560 9.3005
R25895 GND.n6729 GND.n6561 9.3005
R25896 GND.n6728 GND.n6562 9.3005
R25897 GND.n6565 GND.n6563 9.3005
R25898 GND.n6724 GND.n6566 9.3005
R25899 GND.n6723 GND.n6567 9.3005
R25900 GND.n6722 GND.n6568 9.3005
R25901 GND.n6571 GND.n6569 9.3005
R25902 GND.n6718 GND.n6572 9.3005
R25903 GND.n6717 GND.n6573 9.3005
R25904 GND.n6716 GND.n6574 9.3005
R25905 GND.n6577 GND.n6575 9.3005
R25906 GND.n6712 GND.n6578 9.3005
R25907 GND.n6711 GND.n6579 9.3005
R25908 GND.n6710 GND.n6580 9.3005
R25909 GND.n6583 GND.n6581 9.3005
R25910 GND.n6706 GND.n6584 9.3005
R25911 GND.n6705 GND.n6585 9.3005
R25912 GND.n6704 GND.n6586 9.3005
R25913 GND.n6589 GND.n6587 9.3005
R25914 GND.n6700 GND.n6590 9.3005
R25915 GND.n6699 GND.n6591 9.3005
R25916 GND.n6698 GND.n6592 9.3005
R25917 GND.n6595 GND.n6593 9.3005
R25918 GND.n6694 GND.n6596 9.3005
R25919 GND.n6693 GND.n6597 9.3005
R25920 GND.n6692 GND.n6598 9.3005
R25921 GND.n6601 GND.n6599 9.3005
R25922 GND.n6688 GND.n6602 9.3005
R25923 GND.n6687 GND.n6603 9.3005
R25924 GND.n6686 GND.n6604 9.3005
R25925 GND.n6607 GND.n6605 9.3005
R25926 GND.n6682 GND.n6608 9.3005
R25927 GND.n6681 GND.n6609 9.3005
R25928 GND.n6680 GND.n6610 9.3005
R25929 GND.n6613 GND.n6611 9.3005
R25930 GND.n6676 GND.n6614 9.3005
R25931 GND.n6675 GND.n6615 9.3005
R25932 GND.n6674 GND.n6616 9.3005
R25933 GND.n6619 GND.n6617 9.3005
R25934 GND.n6670 GND.n6620 9.3005
R25935 GND.n6669 GND.n6621 9.3005
R25936 GND.n6668 GND.n6622 9.3005
R25937 GND.n6625 GND.n6623 9.3005
R25938 GND.n6664 GND.n6626 9.3005
R25939 GND.n6663 GND.n6627 9.3005
R25940 GND.n6662 GND.n6628 9.3005
R25941 GND.n6631 GND.n6629 9.3005
R25942 GND.n6658 GND.n6632 9.3005
R25943 GND.n6657 GND.n6633 9.3005
R25944 GND.n6656 GND.n6634 9.3005
R25945 GND.n6637 GND.n6635 9.3005
R25946 GND.n6652 GND.n6638 9.3005
R25947 GND.n6651 GND.n6639 9.3005
R25948 GND.n6650 GND.n6640 9.3005
R25949 GND.n6642 GND.n6641 9.3005
R25950 GND.n6646 GND.n102 9.3005
R25951 GND.n7309 GND.n6283 9.3005
R25952 GND.n7308 GND.n6284 9.3005
R25953 GND.n7307 GND.n6285 9.3005
R25954 GND.n6288 GND.n6286 9.3005
R25955 GND.n7303 GND.n6289 9.3005
R25956 GND.n7302 GND.n6290 9.3005
R25957 GND.n7301 GND.n6291 9.3005
R25958 GND.n6294 GND.n6292 9.3005
R25959 GND.n7297 GND.n6295 9.3005
R25960 GND.n7296 GND.n6296 9.3005
R25961 GND.n7295 GND.n6297 9.3005
R25962 GND.n6300 GND.n6298 9.3005
R25963 GND.n7291 GND.n6301 9.3005
R25964 GND.n7290 GND.n6302 9.3005
R25965 GND.n7289 GND.n6303 9.3005
R25966 GND.n6306 GND.n6304 9.3005
R25967 GND.n7285 GND.n6307 9.3005
R25968 GND.n7284 GND.n6308 9.3005
R25969 GND.n7283 GND.n6309 9.3005
R25970 GND.n6312 GND.n6310 9.3005
R25971 GND.n7279 GND.n6313 9.3005
R25972 GND.n7278 GND.n6314 9.3005
R25973 GND.n7277 GND.n6315 9.3005
R25974 GND.n6318 GND.n6316 9.3005
R25975 GND.n7273 GND.n6319 9.3005
R25976 GND.n7272 GND.n6320 9.3005
R25977 GND.n7271 GND.n6321 9.3005
R25978 GND.n6324 GND.n6322 9.3005
R25979 GND.n6431 GND.n6325 9.3005
R25980 GND.n6430 GND.n6326 9.3005
R25981 GND.n6429 GND.n6327 9.3005
R25982 GND.n6330 GND.n6328 9.3005
R25983 GND.n6425 GND.n6331 9.3005
R25984 GND.n6424 GND.n6332 9.3005
R25985 GND.n6423 GND.n6333 9.3005
R25986 GND.n6336 GND.n6334 9.3005
R25987 GND.n6419 GND.n6337 9.3005
R25988 GND.n6418 GND.n6338 9.3005
R25989 GND.n6417 GND.n6339 9.3005
R25990 GND.n6342 GND.n6340 9.3005
R25991 GND.n6413 GND.n6343 9.3005
R25992 GND.n6412 GND.n6344 9.3005
R25993 GND.n6411 GND.n6345 9.3005
R25994 GND.n6348 GND.n6346 9.3005
R25995 GND.n6407 GND.n6349 9.3005
R25996 GND.n6406 GND.n6350 9.3005
R25997 GND.n6405 GND.n6351 9.3005
R25998 GND.n6354 GND.n6352 9.3005
R25999 GND.n6401 GND.n6355 9.3005
R26000 GND.n6400 GND.n6356 9.3005
R26001 GND.n6399 GND.n6357 9.3005
R26002 GND.n6360 GND.n6358 9.3005
R26003 GND.n6395 GND.n6361 9.3005
R26004 GND.n6394 GND.n6362 9.3005
R26005 GND.n6393 GND.n6363 9.3005
R26006 GND.n6366 GND.n6364 9.3005
R26007 GND.n6389 GND.n6367 9.3005
R26008 GND.n6388 GND.n6368 9.3005
R26009 GND.n6387 GND.n6369 9.3005
R26010 GND.n6372 GND.n6370 9.3005
R26011 GND.n6383 GND.n6373 9.3005
R26012 GND.n6382 GND.n6374 9.3005
R26013 GND.n6381 GND.n6375 9.3005
R26014 GND.n6378 GND.n6377 9.3005
R26015 GND.n6376 GND.n464 9.3005
R26016 GND.n10644 GND.n465 9.3005
R26017 GND.n10643 GND.n466 9.3005
R26018 GND.n10642 GND.n467 9.3005
R26019 GND.n472 GND.n468 9.3005
R26020 GND.n10636 GND.n473 9.3005
R26021 GND.n10635 GND.n474 9.3005
R26022 GND.n10634 GND.n475 9.3005
R26023 GND.n480 GND.n476 9.3005
R26024 GND.n10628 GND.n481 9.3005
R26025 GND.n10627 GND.n482 9.3005
R26026 GND.n10626 GND.n483 9.3005
R26027 GND.n488 GND.n484 9.3005
R26028 GND.n10620 GND.n489 9.3005
R26029 GND.n10619 GND.n490 9.3005
R26030 GND.n10618 GND.n491 9.3005
R26031 GND.n496 GND.n492 9.3005
R26032 GND.n10612 GND.n497 9.3005
R26033 GND.n10611 GND.n498 9.3005
R26034 GND.n10610 GND.n499 9.3005
R26035 GND.n504 GND.n500 9.3005
R26036 GND.n10604 GND.n505 9.3005
R26037 GND.n10603 GND.n506 9.3005
R26038 GND.n10602 GND.n507 9.3005
R26039 GND.n512 GND.n508 9.3005
R26040 GND.n10596 GND.n513 9.3005
R26041 GND.n10595 GND.n514 9.3005
R26042 GND.n10594 GND.n515 9.3005
R26043 GND.n520 GND.n516 9.3005
R26044 GND.n10588 GND.n521 9.3005
R26045 GND.n10587 GND.n522 9.3005
R26046 GND.n10586 GND.n523 9.3005
R26047 GND.n528 GND.n524 9.3005
R26048 GND.n10580 GND.n529 9.3005
R26049 GND.n10579 GND.n530 9.3005
R26050 GND.n10578 GND.n531 9.3005
R26051 GND.n536 GND.n532 9.3005
R26052 GND.n10572 GND.n537 9.3005
R26053 GND.n10571 GND.n538 9.3005
R26054 GND.n10570 GND.n539 9.3005
R26055 GND.n544 GND.n540 9.3005
R26056 GND.n10564 GND.n545 9.3005
R26057 GND.n10563 GND.n546 9.3005
R26058 GND.n10562 GND.n547 9.3005
R26059 GND.n552 GND.n548 9.3005
R26060 GND.n10556 GND.n553 9.3005
R26061 GND.n10555 GND.n554 9.3005
R26062 GND.n10554 GND.n555 9.3005
R26063 GND.n560 GND.n556 9.3005
R26064 GND.n10548 GND.n561 9.3005
R26065 GND.n10547 GND.n562 9.3005
R26066 GND.n10546 GND.n563 9.3005
R26067 GND.n568 GND.n564 9.3005
R26068 GND.n10540 GND.n569 9.3005
R26069 GND.n10539 GND.n570 9.3005
R26070 GND.n10538 GND.n571 9.3005
R26071 GND.n10530 GND.n572 9.3005
R26072 GND.n8927 GND.n8926 9.3005
R26073 GND.n8925 GND.n1582 9.3005
R26074 GND.n8924 GND.n8923 9.3005
R26075 GND.n1584 GND.n1583 9.3005
R26076 GND.n8917 GND.n1590 9.3005
R26077 GND.n8916 GND.n1591 9.3005
R26078 GND.n8915 GND.n1592 9.3005
R26079 GND.n1597 GND.n1593 9.3005
R26080 GND.n8909 GND.n1598 9.3005
R26081 GND.n8908 GND.n1599 9.3005
R26082 GND.n8907 GND.n1600 9.3005
R26083 GND.n1605 GND.n1601 9.3005
R26084 GND.n8901 GND.n1606 9.3005
R26085 GND.n8900 GND.n1607 9.3005
R26086 GND.n8899 GND.n1608 9.3005
R26087 GND.n1613 GND.n1609 9.3005
R26088 GND.n8893 GND.n1614 9.3005
R26089 GND.n8892 GND.n1615 9.3005
R26090 GND.n8891 GND.n1616 9.3005
R26091 GND.n1621 GND.n1617 9.3005
R26092 GND.n8885 GND.n1622 9.3005
R26093 GND.n8884 GND.n1623 9.3005
R26094 GND.n8883 GND.n1624 9.3005
R26095 GND.n1629 GND.n1625 9.3005
R26096 GND.n8877 GND.n1630 9.3005
R26097 GND.n8876 GND.n1631 9.3005
R26098 GND.n8875 GND.n1632 9.3005
R26099 GND.n1637 GND.n1633 9.3005
R26100 GND.n8869 GND.n1638 9.3005
R26101 GND.n8868 GND.n1639 9.3005
R26102 GND.n8867 GND.n1640 9.3005
R26103 GND.n1645 GND.n1641 9.3005
R26104 GND.n8861 GND.n1646 9.3005
R26105 GND.n8860 GND.n1647 9.3005
R26106 GND.n8859 GND.n1648 9.3005
R26107 GND.n1653 GND.n1649 9.3005
R26108 GND.n8853 GND.n1654 9.3005
R26109 GND.n8852 GND.n1655 9.3005
R26110 GND.n8851 GND.n1656 9.3005
R26111 GND.n1661 GND.n1657 9.3005
R26112 GND.n8845 GND.n1662 9.3005
R26113 GND.n8844 GND.n1663 9.3005
R26114 GND.n8843 GND.n1664 9.3005
R26115 GND.n1669 GND.n1665 9.3005
R26116 GND.n8837 GND.n1670 9.3005
R26117 GND.n8836 GND.n1671 9.3005
R26118 GND.n8835 GND.n1672 9.3005
R26119 GND.n1677 GND.n1673 9.3005
R26120 GND.n8829 GND.n1678 9.3005
R26121 GND.n8828 GND.n1679 9.3005
R26122 GND.n8827 GND.n1680 9.3005
R26123 GND.n1685 GND.n1681 9.3005
R26124 GND.n8821 GND.n1686 9.3005
R26125 GND.n8820 GND.n1687 9.3005
R26126 GND.n8819 GND.n1688 9.3005
R26127 GND.n1809 GND.n1689 9.3005
R26128 GND.n1810 GND.n1808 9.3005
R26129 GND.n8695 GND.n1811 9.3005
R26130 GND.n8694 GND.n1812 9.3005
R26131 GND.n8693 GND.n1813 9.3005
R26132 GND.n2970 GND.n1814 9.3005
R26133 GND.n2972 GND.n2971 9.3005
R26134 GND.n2976 GND.n2975 9.3005
R26135 GND.n2977 GND.n2969 9.3005
R26136 GND.n3148 GND.n2978 9.3005
R26137 GND.n3147 GND.n2979 9.3005
R26138 GND.n3146 GND.n2980 9.3005
R26139 GND.n2983 GND.n2981 9.3005
R26140 GND.n3142 GND.n2984 9.3005
R26141 GND.n3141 GND.n2985 9.3005
R26142 GND.n3140 GND.n2986 9.3005
R26143 GND.n2989 GND.n2987 9.3005
R26144 GND.n3136 GND.n2990 9.3005
R26145 GND.n3135 GND.n2991 9.3005
R26146 GND.n3134 GND.n2992 9.3005
R26147 GND.n2995 GND.n2993 9.3005
R26148 GND.n3130 GND.n2996 9.3005
R26149 GND.n3129 GND.n2997 9.3005
R26150 GND.n3128 GND.n2998 9.3005
R26151 GND.n3001 GND.n2999 9.3005
R26152 GND.n3124 GND.n3002 9.3005
R26153 GND.n3123 GND.n3003 9.3005
R26154 GND.n3122 GND.n3004 9.3005
R26155 GND.n3007 GND.n3005 9.3005
R26156 GND.n3118 GND.n3008 9.3005
R26157 GND.n3117 GND.n3009 9.3005
R26158 GND.n3116 GND.n3010 9.3005
R26159 GND.n3013 GND.n3011 9.3005
R26160 GND.n3112 GND.n3014 9.3005
R26161 GND.n3111 GND.n3015 9.3005
R26162 GND.n3110 GND.n3016 9.3005
R26163 GND.n3019 GND.n3017 9.3005
R26164 GND.n3106 GND.n3020 9.3005
R26165 GND.n3105 GND.n3021 9.3005
R26166 GND.n3104 GND.n3022 9.3005
R26167 GND.n3025 GND.n3023 9.3005
R26168 GND.n3100 GND.n3026 9.3005
R26169 GND.n3099 GND.n3027 9.3005
R26170 GND.n3098 GND.n3028 9.3005
R26171 GND.n3031 GND.n3029 9.3005
R26172 GND.n3094 GND.n3032 9.3005
R26173 GND.n3093 GND.n3033 9.3005
R26174 GND.n3092 GND.n3034 9.3005
R26175 GND.n3037 GND.n3035 9.3005
R26176 GND.n3088 GND.n3038 9.3005
R26177 GND.n3087 GND.n3039 9.3005
R26178 GND.n3086 GND.n3040 9.3005
R26179 GND.n3043 GND.n3041 9.3005
R26180 GND.n3082 GND.n3044 9.3005
R26181 GND.n3081 GND.n3045 9.3005
R26182 GND.n3080 GND.n3046 9.3005
R26183 GND.n3049 GND.n3047 9.3005
R26184 GND.n3076 GND.n3050 9.3005
R26185 GND.n3075 GND.n3051 9.3005
R26186 GND.n3074 GND.n3052 9.3005
R26187 GND.n3055 GND.n3053 9.3005
R26188 GND.n3070 GND.n3056 9.3005
R26189 GND.n3069 GND.n3057 9.3005
R26190 GND.n3068 GND.n3058 9.3005
R26191 GND.n3060 GND.n3059 9.3005
R26192 GND.n8928 GND.n1581 9.3005
R26193 GND.n8934 GND.n1575 9.3005
R26194 GND.n8935 GND.n1574 9.3005
R26195 GND.n8936 GND.n1573 9.3005
R26196 GND.n1572 GND.n1568 9.3005
R26197 GND.n8942 GND.n1567 9.3005
R26198 GND.n8943 GND.n1566 9.3005
R26199 GND.n8944 GND.n1565 9.3005
R26200 GND.n1564 GND.n1560 9.3005
R26201 GND.n8950 GND.n1559 9.3005
R26202 GND.n8951 GND.n1558 9.3005
R26203 GND.n8952 GND.n1557 9.3005
R26204 GND.n1556 GND.n1552 9.3005
R26205 GND.n8958 GND.n1551 9.3005
R26206 GND.n8959 GND.n1550 9.3005
R26207 GND.n8960 GND.n1549 9.3005
R26208 GND.n1548 GND.n1544 9.3005
R26209 GND.n8966 GND.n1543 9.3005
R26210 GND.n8967 GND.n1542 9.3005
R26211 GND.n8968 GND.n1541 9.3005
R26212 GND.n1540 GND.n1536 9.3005
R26213 GND.n8974 GND.n1535 9.3005
R26214 GND.n8975 GND.n1534 9.3005
R26215 GND.n8976 GND.n1533 9.3005
R26216 GND.n1532 GND.n1528 9.3005
R26217 GND.n8982 GND.n1527 9.3005
R26218 GND.n8983 GND.n1526 9.3005
R26219 GND.n8984 GND.n1525 9.3005
R26220 GND.n1524 GND.n1520 9.3005
R26221 GND.n8990 GND.n1519 9.3005
R26222 GND.n8991 GND.n1518 9.3005
R26223 GND.n8992 GND.n1517 9.3005
R26224 GND.n1516 GND.n1512 9.3005
R26225 GND.n8998 GND.n1511 9.3005
R26226 GND.n8999 GND.n1510 9.3005
R26227 GND.n9000 GND.n1509 9.3005
R26228 GND.n1508 GND.n1504 9.3005
R26229 GND.n9006 GND.n1503 9.3005
R26230 GND.n9007 GND.n1502 9.3005
R26231 GND.n9008 GND.n1501 9.3005
R26232 GND.n1500 GND.n1496 9.3005
R26233 GND.n9014 GND.n1495 9.3005
R26234 GND.n9015 GND.n1494 9.3005
R26235 GND.n9016 GND.n1493 9.3005
R26236 GND.n1492 GND.n1488 9.3005
R26237 GND.n9022 GND.n1487 9.3005
R26238 GND.n9023 GND.n1486 9.3005
R26239 GND.n9024 GND.n1485 9.3005
R26240 GND.n1484 GND.n1480 9.3005
R26241 GND.n9030 GND.n1479 9.3005
R26242 GND.n9031 GND.n1478 9.3005
R26243 GND.n9032 GND.n1477 9.3005
R26244 GND.n1476 GND.n1472 9.3005
R26245 GND.n9038 GND.n1471 9.3005
R26246 GND.n9039 GND.n1470 9.3005
R26247 GND.n9040 GND.n1469 9.3005
R26248 GND.n1468 GND.n1464 9.3005
R26249 GND.n9046 GND.n1463 9.3005
R26250 GND.n9048 GND.n9047 9.3005
R26251 GND.n1580 GND.n1576 9.3005
R26252 GND.n8043 GND.n3875 9.3005
R26253 GND.n8044 GND.n8043 9.3005
R26254 GND.n8361 GND.n8360 9.3005
R26255 GND.n8357 GND.n2187 9.3005
R26256 GND.n8356 GND.n8355 9.3005
R26257 GND.n8354 GND.n2188 9.3005
R26258 GND.n8353 GND.n8352 9.3005
R26259 GND.n8349 GND.n2191 9.3005
R26260 GND.n8348 GND.n8347 9.3005
R26261 GND.n8346 GND.n2192 9.3005
R26262 GND.n8345 GND.n8344 9.3005
R26263 GND.n8341 GND.n2195 9.3005
R26264 GND.n8340 GND.n8339 9.3005
R26265 GND.n8338 GND.n2196 9.3005
R26266 GND.n8337 GND.n8336 9.3005
R26267 GND.n8331 GND.n2199 9.3005
R26268 GND.n8330 GND.n8329 9.3005
R26269 GND.n8328 GND.n2200 9.3005
R26270 GND.n8327 GND.n8326 9.3005
R26271 GND.n8323 GND.n2203 9.3005
R26272 GND.n8322 GND.n8321 9.3005
R26273 GND.n8320 GND.n2204 9.3005
R26274 GND.n8319 GND.n8318 9.3005
R26275 GND.n8315 GND.n2207 9.3005
R26276 GND.n8314 GND.n8313 9.3005
R26277 GND.n8312 GND.n2208 9.3005
R26278 GND.n8311 GND.n8310 9.3005
R26279 GND.n8454 GND.n8453 9.3005
R26280 GND.n8452 GND.n2186 9.3005
R26281 GND.n8451 GND.n8450 9.3005
R26282 GND.n8449 GND.n8363 9.3005
R26283 GND.n8448 GND.n8447 9.3005
R26284 GND.n8446 GND.n8368 9.3005
R26285 GND.n8445 GND.n8444 9.3005
R26286 GND.n8443 GND.n8369 9.3005
R26287 GND.n8442 GND.n8441 9.3005
R26288 GND.n8440 GND.n8374 9.3005
R26289 GND.n8439 GND.n8438 9.3005
R26290 GND.n8437 GND.n8375 9.3005
R26291 GND.n8436 GND.n8435 9.3005
R26292 GND.n8434 GND.n8380 9.3005
R26293 GND.n8433 GND.n8432 9.3005
R26294 GND.n8431 GND.n8381 9.3005
R26295 GND.n8430 GND.n8429 9.3005
R26296 GND.n8428 GND.n8389 9.3005
R26297 GND.n8427 GND.n8426 9.3005
R26298 GND.n8425 GND.n8390 9.3005
R26299 GND.n8424 GND.n8423 9.3005
R26300 GND.n8422 GND.n8395 9.3005
R26301 GND.n8421 GND.n8420 9.3005
R26302 GND.n8419 GND.n8396 9.3005
R26303 GND.n8418 GND.n8417 9.3005
R26304 GND.n8416 GND.n8401 9.3005
R26305 GND.n8415 GND.n8414 9.3005
R26306 GND.n8413 GND.n8402 9.3005
R26307 GND.n8412 GND.n8408 9.3005
R26308 GND.n8411 GND.n8410 9.3005
R26309 GND.n1853 GND.n1852 9.3005
R26310 GND.n1855 GND.n1847 9.3005
R26311 GND.n1857 GND.n1856 9.3005
R26312 GND.n1844 GND.n1842 9.3005
R26313 GND.n8682 GND.n8681 9.3005
R26314 GND.n1845 GND.n1843 9.3005
R26315 GND.n8677 GND.n1863 9.3005
R26316 GND.n8676 GND.n1864 9.3005
R26317 GND.n8675 GND.n1865 9.3005
R26318 GND.n3173 GND.n1866 9.3005
R26319 GND.n8671 GND.n1871 9.3005
R26320 GND.n8670 GND.n1872 9.3005
R26321 GND.n8669 GND.n1873 9.3005
R26322 GND.n2878 GND.n1874 9.3005
R26323 GND.n8665 GND.n1879 9.3005
R26324 GND.n8664 GND.n1880 9.3005
R26325 GND.n8663 GND.n1881 9.3005
R26326 GND.n2855 GND.n1882 9.3005
R26327 GND.n8659 GND.n1887 9.3005
R26328 GND.n8658 GND.n1888 9.3005
R26329 GND.n8657 GND.n1889 9.3005
R26330 GND.n2842 GND.n1890 9.3005
R26331 GND.n8653 GND.n1895 9.3005
R26332 GND.n8652 GND.n1896 9.3005
R26333 GND.n8651 GND.n1897 9.3005
R26334 GND.n3245 GND.n1898 9.3005
R26335 GND.n8647 GND.n1903 9.3005
R26336 GND.n8646 GND.n1904 9.3005
R26337 GND.n8645 GND.n1905 9.3005
R26338 GND.n3272 GND.n1906 9.3005
R26339 GND.n8641 GND.n1911 9.3005
R26340 GND.n8640 GND.n1912 9.3005
R26341 GND.n8639 GND.n1913 9.3005
R26342 GND.n2787 GND.n1914 9.3005
R26343 GND.n8635 GND.n1919 9.3005
R26344 GND.n8634 GND.n1920 9.3005
R26345 GND.n8633 GND.n1921 9.3005
R26346 GND.n2764 GND.n1922 9.3005
R26347 GND.n8629 GND.n1927 9.3005
R26348 GND.n8628 GND.n1928 9.3005
R26349 GND.n8627 GND.n1929 9.3005
R26350 GND.n2751 GND.n1930 9.3005
R26351 GND.n8623 GND.n1935 9.3005
R26352 GND.n8622 GND.n1936 9.3005
R26353 GND.n8621 GND.n1937 9.3005
R26354 GND.n3344 GND.n1938 9.3005
R26355 GND.n8617 GND.n1943 9.3005
R26356 GND.n8616 GND.n1944 9.3005
R26357 GND.n8615 GND.n1945 9.3005
R26358 GND.n3371 GND.n1946 9.3005
R26359 GND.n8611 GND.n1951 9.3005
R26360 GND.n8610 GND.n1952 9.3005
R26361 GND.n8609 GND.n1953 9.3005
R26362 GND.n2696 GND.n1954 9.3005
R26363 GND.n8605 GND.n1959 9.3005
R26364 GND.n8604 GND.n1960 9.3005
R26365 GND.n8603 GND.n1961 9.3005
R26366 GND.n2673 GND.n1962 9.3005
R26367 GND.n8599 GND.n1967 9.3005
R26368 GND.n8598 GND.n1968 9.3005
R26369 GND.n8597 GND.n1969 9.3005
R26370 GND.n2662 GND.n1970 9.3005
R26371 GND.n8593 GND.n1975 9.3005
R26372 GND.n8592 GND.n1976 9.3005
R26373 GND.n8591 GND.n1977 9.3005
R26374 GND.n2506 GND.n1978 9.3005
R26375 GND.n8587 GND.n1983 9.3005
R26376 GND.n8586 GND.n1984 9.3005
R26377 GND.n8585 GND.n1985 9.3005
R26378 GND.n2529 GND.n1986 9.3005
R26379 GND.n8581 GND.n1991 9.3005
R26380 GND.n8580 GND.n1992 9.3005
R26381 GND.n8579 GND.n1993 9.3005
R26382 GND.n2485 GND.n1994 9.3005
R26383 GND.n8575 GND.n1999 9.3005
R26384 GND.n8574 GND.n2000 9.3005
R26385 GND.n8573 GND.n2001 9.3005
R26386 GND.n3512 GND.n2002 9.3005
R26387 GND.n8569 GND.n2007 9.3005
R26388 GND.n8568 GND.n2008 9.3005
R26389 GND.n8567 GND.n2009 9.3005
R26390 GND.n3540 GND.n2010 9.3005
R26391 GND.n8563 GND.n2015 9.3005
R26392 GND.n8562 GND.n2016 9.3005
R26393 GND.n8561 GND.n2017 9.3005
R26394 GND.n2433 GND.n2018 9.3005
R26395 GND.n8557 GND.n2023 9.3005
R26396 GND.n8556 GND.n2024 9.3005
R26397 GND.n8555 GND.n2025 9.3005
R26398 GND.n2411 GND.n2026 9.3005
R26399 GND.n8551 GND.n2031 9.3005
R26400 GND.n8550 GND.n2032 9.3005
R26401 GND.n8549 GND.n2033 9.3005
R26402 GND.n2398 GND.n2034 9.3005
R26403 GND.n8545 GND.n2039 9.3005
R26404 GND.n8544 GND.n2040 9.3005
R26405 GND.n8543 GND.n2041 9.3005
R26406 GND.n3615 GND.n2042 9.3005
R26407 GND.n8539 GND.n2047 9.3005
R26408 GND.n8538 GND.n2048 9.3005
R26409 GND.n8537 GND.n2049 9.3005
R26410 GND.n3643 GND.n2050 9.3005
R26411 GND.n8533 GND.n2055 9.3005
R26412 GND.n8532 GND.n2056 9.3005
R26413 GND.n8531 GND.n2057 9.3005
R26414 GND.n2349 GND.n2058 9.3005
R26415 GND.n8527 GND.n2063 9.3005
R26416 GND.n8526 GND.n2064 9.3005
R26417 GND.n8525 GND.n2065 9.3005
R26418 GND.n2336 GND.n2066 9.3005
R26419 GND.n8521 GND.n2071 9.3005
R26420 GND.n8520 GND.n2072 9.3005
R26421 GND.n8519 GND.n2073 9.3005
R26422 GND.n2308 GND.n2074 9.3005
R26423 GND.n8515 GND.n2079 9.3005
R26424 GND.n8514 GND.n2080 9.3005
R26425 GND.n8513 GND.n2081 9.3005
R26426 GND.n8204 GND.n2082 9.3005
R26427 GND.n8509 GND.n2087 9.3005
R26428 GND.n8508 GND.n2088 9.3005
R26429 GND.n8507 GND.n2089 9.3005
R26430 GND.n8232 GND.n2090 9.3005
R26431 GND.n8503 GND.n2095 9.3005
R26432 GND.n8502 GND.n2096 9.3005
R26433 GND.n8501 GND.n2097 9.3005
R26434 GND.n2257 GND.n2098 9.3005
R26435 GND.n8497 GND.n2103 9.3005
R26436 GND.n8496 GND.n2104 9.3005
R26437 GND.n8495 GND.n2105 9.3005
R26438 GND.n2235 GND.n2106 9.3005
R26439 GND.n8491 GND.n2111 9.3005
R26440 GND.n8490 GND.n2112 9.3005
R26441 GND.n8489 GND.n2113 9.3005
R26442 GND.n2224 GND.n2114 9.3005
R26443 GND.n8485 GND.n2119 9.3005
R26444 GND.n8484 GND.n2120 9.3005
R26445 GND.n8483 GND.n2121 9.3005
R26446 GND.n1800 GND.n1796 9.3005
R26447 GND.n1852 GND.n1851 9.3005
R26448 GND.n1847 GND.n1846 9.3005
R26449 GND.n1858 GND.n1857 9.3005
R26450 GND.n1859 GND.n1844 9.3005
R26451 GND.n8681 GND.n8680 9.3005
R26452 GND.n8679 GND.n1845 9.3005
R26453 GND.n8678 GND.n8677 9.3005
R26454 GND.n8676 GND.n1862 9.3005
R26455 GND.n8675 GND.n8674 9.3005
R26456 GND.n8673 GND.n1866 9.3005
R26457 GND.n8672 GND.n8671 9.3005
R26458 GND.n8670 GND.n1870 9.3005
R26459 GND.n8669 GND.n8668 9.3005
R26460 GND.n8667 GND.n1874 9.3005
R26461 GND.n8666 GND.n8665 9.3005
R26462 GND.n8664 GND.n1878 9.3005
R26463 GND.n8663 GND.n8662 9.3005
R26464 GND.n8661 GND.n1882 9.3005
R26465 GND.n8660 GND.n8659 9.3005
R26466 GND.n8658 GND.n1886 9.3005
R26467 GND.n8657 GND.n8656 9.3005
R26468 GND.n8655 GND.n1890 9.3005
R26469 GND.n8654 GND.n8653 9.3005
R26470 GND.n8652 GND.n1894 9.3005
R26471 GND.n8651 GND.n8650 9.3005
R26472 GND.n8649 GND.n1898 9.3005
R26473 GND.n8648 GND.n8647 9.3005
R26474 GND.n8646 GND.n1902 9.3005
R26475 GND.n8645 GND.n8644 9.3005
R26476 GND.n8643 GND.n1906 9.3005
R26477 GND.n8642 GND.n8641 9.3005
R26478 GND.n8640 GND.n1910 9.3005
R26479 GND.n8639 GND.n8638 9.3005
R26480 GND.n8637 GND.n1914 9.3005
R26481 GND.n8636 GND.n8635 9.3005
R26482 GND.n8634 GND.n1918 9.3005
R26483 GND.n8633 GND.n8632 9.3005
R26484 GND.n8631 GND.n1922 9.3005
R26485 GND.n8630 GND.n8629 9.3005
R26486 GND.n8628 GND.n1926 9.3005
R26487 GND.n8627 GND.n8626 9.3005
R26488 GND.n8625 GND.n1930 9.3005
R26489 GND.n8624 GND.n8623 9.3005
R26490 GND.n8622 GND.n1934 9.3005
R26491 GND.n8621 GND.n8620 9.3005
R26492 GND.n8619 GND.n1938 9.3005
R26493 GND.n8618 GND.n8617 9.3005
R26494 GND.n8616 GND.n1942 9.3005
R26495 GND.n8615 GND.n8614 9.3005
R26496 GND.n8613 GND.n1946 9.3005
R26497 GND.n8612 GND.n8611 9.3005
R26498 GND.n8610 GND.n1950 9.3005
R26499 GND.n8609 GND.n8608 9.3005
R26500 GND.n8607 GND.n1954 9.3005
R26501 GND.n8606 GND.n8605 9.3005
R26502 GND.n8604 GND.n1958 9.3005
R26503 GND.n8603 GND.n8602 9.3005
R26504 GND.n8601 GND.n1962 9.3005
R26505 GND.n8600 GND.n8599 9.3005
R26506 GND.n8598 GND.n1966 9.3005
R26507 GND.n8597 GND.n8596 9.3005
R26508 GND.n8595 GND.n1970 9.3005
R26509 GND.n8594 GND.n8593 9.3005
R26510 GND.n8592 GND.n1974 9.3005
R26511 GND.n8591 GND.n8590 9.3005
R26512 GND.n8589 GND.n1978 9.3005
R26513 GND.n8588 GND.n8587 9.3005
R26514 GND.n8586 GND.n1982 9.3005
R26515 GND.n8585 GND.n8584 9.3005
R26516 GND.n8583 GND.n1986 9.3005
R26517 GND.n8582 GND.n8581 9.3005
R26518 GND.n8580 GND.n1990 9.3005
R26519 GND.n8579 GND.n8578 9.3005
R26520 GND.n8577 GND.n1994 9.3005
R26521 GND.n8576 GND.n8575 9.3005
R26522 GND.n8574 GND.n1998 9.3005
R26523 GND.n8573 GND.n8572 9.3005
R26524 GND.n8571 GND.n2002 9.3005
R26525 GND.n8570 GND.n8569 9.3005
R26526 GND.n8568 GND.n2006 9.3005
R26527 GND.n8567 GND.n8566 9.3005
R26528 GND.n8565 GND.n2010 9.3005
R26529 GND.n8564 GND.n8563 9.3005
R26530 GND.n8562 GND.n2014 9.3005
R26531 GND.n8561 GND.n8560 9.3005
R26532 GND.n8559 GND.n2018 9.3005
R26533 GND.n8558 GND.n8557 9.3005
R26534 GND.n8556 GND.n2022 9.3005
R26535 GND.n8555 GND.n8554 9.3005
R26536 GND.n8553 GND.n2026 9.3005
R26537 GND.n8552 GND.n8551 9.3005
R26538 GND.n8550 GND.n2030 9.3005
R26539 GND.n8549 GND.n8548 9.3005
R26540 GND.n8547 GND.n2034 9.3005
R26541 GND.n8546 GND.n8545 9.3005
R26542 GND.n8544 GND.n2038 9.3005
R26543 GND.n8543 GND.n8542 9.3005
R26544 GND.n8541 GND.n2042 9.3005
R26545 GND.n8540 GND.n8539 9.3005
R26546 GND.n8538 GND.n2046 9.3005
R26547 GND.n8537 GND.n8536 9.3005
R26548 GND.n8535 GND.n2050 9.3005
R26549 GND.n8534 GND.n8533 9.3005
R26550 GND.n8532 GND.n2054 9.3005
R26551 GND.n8531 GND.n8530 9.3005
R26552 GND.n8529 GND.n2058 9.3005
R26553 GND.n8528 GND.n8527 9.3005
R26554 GND.n8526 GND.n2062 9.3005
R26555 GND.n8525 GND.n8524 9.3005
R26556 GND.n8523 GND.n2066 9.3005
R26557 GND.n8522 GND.n8521 9.3005
R26558 GND.n8520 GND.n2070 9.3005
R26559 GND.n8519 GND.n8518 9.3005
R26560 GND.n8517 GND.n2074 9.3005
R26561 GND.n8516 GND.n8515 9.3005
R26562 GND.n8514 GND.n2078 9.3005
R26563 GND.n8513 GND.n8512 9.3005
R26564 GND.n8511 GND.n2082 9.3005
R26565 GND.n8510 GND.n8509 9.3005
R26566 GND.n8508 GND.n2086 9.3005
R26567 GND.n8507 GND.n8506 9.3005
R26568 GND.n8505 GND.n2090 9.3005
R26569 GND.n8504 GND.n8503 9.3005
R26570 GND.n8502 GND.n2094 9.3005
R26571 GND.n8501 GND.n8500 9.3005
R26572 GND.n8499 GND.n2098 9.3005
R26573 GND.n8498 GND.n8497 9.3005
R26574 GND.n8496 GND.n2102 9.3005
R26575 GND.n8495 GND.n8494 9.3005
R26576 GND.n8493 GND.n2106 9.3005
R26577 GND.n8492 GND.n8491 9.3005
R26578 GND.n8490 GND.n2110 9.3005
R26579 GND.n8489 GND.n8488 9.3005
R26580 GND.n8487 GND.n2114 9.3005
R26581 GND.n8486 GND.n8485 9.3005
R26582 GND.n8484 GND.n2118 9.3005
R26583 GND.n8483 GND.n8482 9.3005
R26584 GND.n1848 GND.n1796 9.3005
R26585 GND.n2946 GND.n2945 9.3005
R26586 GND.n2944 GND.n2916 9.3005
R26587 GND.n2943 GND.n2942 9.3005
R26588 GND.n2939 GND.n2918 9.3005
R26589 GND.n2936 GND.n2935 9.3005
R26590 GND.n2934 GND.n2919 9.3005
R26591 GND.n2933 GND.n2932 9.3005
R26592 GND.n2929 GND.n2920 9.3005
R26593 GND.n2926 GND.n2925 9.3005
R26594 GND.n2924 GND.n2923 9.3005
R26595 GND.n1798 GND.n1797 9.3005
R26596 GND.n8702 GND.n8701 9.3005
R26597 GND.n2947 GND.n2912 9.3005
R26598 GND.n2950 GND.n2949 9.3005
R26599 GND.n2953 GND.n2952 9.3005
R26600 GND.n2956 GND.n2910 9.3005
R26601 GND.n2958 GND.n2957 9.3005
R26602 GND.n2959 GND.n2909 9.3005
R26603 GND.n2961 GND.n2960 9.3005
R26604 GND.n2962 GND.n2905 9.3005
R26605 GND.n3163 GND.n3162 9.3005
R26606 GND.n3164 GND.n2903 9.3005
R26607 GND.n3167 GND.n3166 9.3005
R26608 GND.n3165 GND.n2904 9.3005
R26609 GND.n2884 GND.n2883 9.3005
R26610 GND.n3188 GND.n3187 9.3005
R26611 GND.n3189 GND.n2881 9.3005
R26612 GND.n3192 GND.n3191 9.3005
R26613 GND.n3190 GND.n2882 9.3005
R26614 GND.n2862 GND.n2861 9.3005
R26615 GND.n3213 GND.n3212 9.3005
R26616 GND.n3214 GND.n2859 9.3005
R26617 GND.n3217 GND.n3216 9.3005
R26618 GND.n3215 GND.n2860 9.3005
R26619 GND.n2838 GND.n2837 9.3005
R26620 GND.n3237 GND.n3236 9.3005
R26621 GND.n3238 GND.n2835 9.3005
R26622 GND.n3241 GND.n3240 9.3005
R26623 GND.n3239 GND.n2836 9.3005
R26624 GND.n2815 GND.n2814 9.3005
R26625 GND.n3262 GND.n3261 9.3005
R26626 GND.n3263 GND.n2812 9.3005
R26627 GND.n3266 GND.n3265 9.3005
R26628 GND.n3264 GND.n2813 9.3005
R26629 GND.n2793 GND.n2792 9.3005
R26630 GND.n3287 GND.n3286 9.3005
R26631 GND.n3288 GND.n2790 9.3005
R26632 GND.n3291 GND.n3290 9.3005
R26633 GND.n3289 GND.n2791 9.3005
R26634 GND.n2771 GND.n2770 9.3005
R26635 GND.n3312 GND.n3311 9.3005
R26636 GND.n3313 GND.n2768 9.3005
R26637 GND.n3316 GND.n3315 9.3005
R26638 GND.n3314 GND.n2769 9.3005
R26639 GND.n2747 GND.n2746 9.3005
R26640 GND.n3336 GND.n3335 9.3005
R26641 GND.n3337 GND.n2744 9.3005
R26642 GND.n3340 GND.n3339 9.3005
R26643 GND.n3338 GND.n2745 9.3005
R26644 GND.n2724 GND.n2723 9.3005
R26645 GND.n3361 GND.n3360 9.3005
R26646 GND.n3362 GND.n2721 9.3005
R26647 GND.n3365 GND.n3364 9.3005
R26648 GND.n3363 GND.n2722 9.3005
R26649 GND.n2702 GND.n2701 9.3005
R26650 GND.n3386 GND.n3385 9.3005
R26651 GND.n3387 GND.n2699 9.3005
R26652 GND.n3390 GND.n3389 9.3005
R26653 GND.n3388 GND.n2700 9.3005
R26654 GND.n2680 GND.n2679 9.3005
R26655 GND.n3411 GND.n3410 9.3005
R26656 GND.n3412 GND.n2677 9.3005
R26657 GND.n3415 GND.n3414 9.3005
R26658 GND.n3413 GND.n2678 9.3005
R26659 GND.n2658 GND.n2657 9.3005
R26660 GND.n3433 GND.n3432 9.3005
R26661 GND.n3434 GND.n2656 9.3005
R26662 GND.n3436 GND.n3435 9.3005
R26663 GND.n3437 GND.n2655 9.3005
R26664 GND.n3441 GND.n3440 9.3005
R26665 GND.n3442 GND.n2654 9.3005
R26666 GND.n3445 GND.n3444 9.3005
R26667 GND.n2951 GND.n2911 9.3005
R26668 GND.n5323 GND.t114 9.0306
R26669 GND.n5794 GND.t146 9.0306
R26670 GND.n7891 GND.t168 8.69615
R26671 GND.t210 GND.n5606 8.69615
R26672 GND.n8816 GND.n1725 8.3617
R26673 GND.n3160 GND.t70 8.3617
R26674 GND.n3150 GND.t70 8.3617
R26675 GND.t46 GND.n2244 8.3617
R26676 GND.n2247 GND.t46 8.3617
R26677 GND.n8457 GND.n2147 8.3617
R26678 GND.n7647 GND.n4602 8.3617
R26679 GND.n7511 GND.t54 8.3617
R26680 GND.n6732 GND.t54 8.3617
R26681 GND.t74 GND.n407 8.3617
R26682 GND.n7178 GND.t74 8.3617
R26683 GND.n10896 GND.n460 8.3617
R26684 GND.n11116 GND.n11115 8.13519
R26685 GND.n3443 GND.n39 8.13519
R26686 GND.n8092 GND.n8091 8.02726
R26687 GND.n3840 GND.n3834 8.02726
R26688 GND.n5333 GND.n5332 8.02726
R26689 GND.n7969 GND.n3946 8.02726
R26690 GND.n7939 GND.n3994 8.02726
R26691 GND.n5490 GND.n4963 8.02726
R26692 GND.n7884 GND.n4086 8.02726
R26693 GND.n5593 GND.n4932 8.02726
R26694 GND.n7829 GND.n4191 8.02726
R26695 GND.n5631 GND.n4899 8.02726
R26696 GND.n7774 GND.n4293 8.02726
R26697 GND.n5801 GND.n5800 8.02726
R26698 GND.n7719 GND.n4396 8.02726
R26699 GND.n4489 GND.n4486 8.02726
R26700 GND.n7658 GND.n4527 8.02726
R26701 GND.t111 GND.n8126 7.35836
R26702 GND.t32 GND.n4026 7.35836
R26703 GND.n4963 GND.t32 7.35836
R26704 GND.n7829 GND.t199 7.35836
R26705 GND.n4916 GND.t199 7.35836
R26706 GND.n7671 GND.t87 7.35836
R26707 GND.n8085 GND.n3814 6.68946
R26708 GND.n5253 GND.n5250 6.68946
R26709 GND.n5343 GND.n5342 6.68946
R26710 GND.n7975 GND.n3936 6.68946
R26711 GND.n7933 GND.n4004 6.68946
R26712 GND.n5475 GND.n4968 6.68946
R26713 GND.n7878 GND.n4109 6.68946
R26714 GND.n5578 GND.n4937 6.68946
R26715 GND.n7823 GND.n4213 6.68946
R26716 GND.n5683 GND.n4905 6.68946
R26717 GND.n7768 GND.n4316 6.68946
R26718 GND.n5778 GND.n4872 6.68946
R26719 GND.n7712 GND.n7711 6.68946
R26720 GND.n4422 GND.n4416 6.68946
R26721 GND.t153 GND.n7664 6.68946
R26722 GND.n8384 GND.n8380 6.4005
R26723 GND.n7570 GND.n4812 6.4005
R26724 GND.n10844 GND.n10750 6.4005
R26725 GND.n10819 GND.n10767 6.4005
R26726 GND.n8762 GND.n1761 6.4005
R26727 GND.n8737 GND.n1778 6.4005
R26728 GND.t11 GND.n3986 6.02057
R26729 GND.n4893 GND.t186 6.02057
R26730 GND.n8057 GND.n8056 5.68612
R26731 GND.n4385 GND.n4376 5.68612
R26732 GND.n21 GND.n13 5.66717
R26733 GND.n61 GND.n53 5.66717
R26734 GND.n8016 GND.n8015 5.62474
R26735 GND.n5863 GND.n5862 5.62474
R26736 GND.n39 GND.n38 5.46258
R26737 GND.n11116 GND.n85 5.46258
R26738 GND.n3822 GND.n3816 5.35167
R26739 GND.n8078 GND.n8077 5.35167
R26740 GND.n7981 GND.n3926 5.35167
R26741 GND.n5352 GND.n5351 5.35167
R26742 GND.n5466 GND.n4973 5.35167
R26743 GND.n7927 GND.n4014 5.35167
R26744 GND.n5569 GND.n4942 5.35167
R26745 GND.n7872 GND.n4119 5.35167
R26746 GND.n5673 GND.n4910 5.35167
R26747 GND.n7817 GND.n4223 5.35167
R26748 GND.n5770 GND.n4877 5.35167
R26749 GND.n7762 GND.n4326 5.35167
R26750 GND.n4476 GND.n4473 5.35167
R26751 GND.n7705 GND.n4414 5.35167
R26752 GND.n8042 GND.n8041 4.74817
R26753 GND.n8037 GND.n8036 4.74817
R26754 GND.n8032 GND.n8031 4.74817
R26755 GND.n8027 GND.n8026 4.74817
R26756 GND.n8022 GND.n8021 4.74817
R26757 GND.n8017 GND.n8016 4.74817
R26758 GND.n8010 GND.n8009 4.74817
R26759 GND.n4843 GND.n4835 4.74817
R26760 GND.n5830 GND.n4842 4.74817
R26761 GND.n5840 GND.n4840 4.74817
R26762 GND.n5845 GND.n4839 4.74817
R26763 GND.n5850 GND.n4838 4.74817
R26764 GND.n5855 GND.n4837 4.74817
R26765 GND.n5862 GND.n4836 4.74817
R26766 GND.n5911 GND.n5910 4.74817
R26767 GND.n5906 GND.n5905 4.74817
R26768 GND.n5901 GND.n5900 4.74817
R26769 GND.n5896 GND.n5895 4.74817
R26770 GND.n5890 GND.n5889 4.74817
R26771 GND.n5891 GND.n5890 4.74817
R26772 GND.n5895 GND.n5894 4.74817
R26773 GND.n5900 GND.n5899 4.74817
R26774 GND.n5905 GND.n5904 4.74817
R26775 GND.n5910 GND.n5909 4.74817
R26776 GND.n5915 GND.n5914 4.74817
R26777 GND.n5832 GND.n4842 4.74817
R26778 GND.n5836 GND.n4840 4.74817
R26779 GND.n5841 GND.n4839 4.74817
R26780 GND.n5846 GND.n4838 4.74817
R26781 GND.n5851 GND.n4837 4.74817
R26782 GND.n5856 GND.n4836 4.74817
R26783 GND.n5864 GND.n4835 4.74817
R26784 GND.n6239 GND.n106 4.74817
R26785 GND.n104 GND.n98 4.74817
R26786 GND.n11108 GND.n99 4.74817
R26787 GND.n107 GND.n103 4.74817
R26788 GND.n7335 GND.n106 4.74817
R26789 GND.n6255 GND.n104 4.74817
R26790 GND.n11109 GND.n11108 4.74817
R26791 GND.n6267 GND.n103 4.74817
R26792 GND.n3493 GND.n3492 4.74817
R26793 GND.n3476 GND.n2495 4.74817
R26794 GND.n3453 GND.n2494 4.74817
R26795 GND.n3456 GND.n2493 4.74817
R26796 GND.n3493 GND.n2497 4.74817
R26797 GND.n2523 GND.n2495 4.74817
R26798 GND.n3475 GND.n2494 4.74817
R26799 GND.n3454 GND.n2493 4.74817
R26800 GND.n3062 GND.n3061 4.74817
R26801 GND.n3482 GND.n3481 4.74817
R26802 GND.n2535 GND.n2534 4.74817
R26803 GND.n3466 GND.n3465 4.74817
R26804 GND.n2647 GND.n2536 4.74817
R26805 GND.n6644 GND.n6262 4.74817
R26806 GND.n7329 GND.n7328 4.74817
R26807 GND.n7324 GND.n6263 4.74817
R26808 GND.n7322 GND.n7321 4.74817
R26809 GND.n6282 GND.n6281 4.74817
R26810 GND.n3061 GND.n2512 4.74817
R26811 GND.n3483 GND.n3482 4.74817
R26812 GND.n2534 GND.n2513 4.74817
R26813 GND.n3467 GND.n3466 4.74817
R26814 GND.n3464 GND.n2536 4.74817
R26815 GND.n6645 GND.n6644 4.74817
R26816 GND.n7330 GND.n7329 4.74817
R26817 GND.n7327 GND.n6263 4.74817
R26818 GND.n7323 GND.n7322 4.74817
R26819 GND.n6281 GND.n6265 4.74817
R26820 GND.n8477 GND.n8476 4.74817
R26821 GND.n8475 GND.n8474 4.74817
R26822 GND.n8472 GND.n8471 4.74817
R26823 GND.n8469 GND.n8468 4.74817
R26824 GND.n8466 GND.n8465 4.74817
R26825 GND.n8463 GND.n8462 4.74817
R26826 GND.n8474 GND.n8473 4.74817
R26827 GND.n8471 GND.n8470 4.74817
R26828 GND.n8468 GND.n8467 4.74817
R26829 GND.n8465 GND.n8464 4.74817
R26830 GND.n8462 GND.n8461 4.74817
R26831 GND.n8010 GND.n3876 4.74817
R26832 GND.n8020 GND.n8017 4.74817
R26833 GND.n8025 GND.n8022 4.74817
R26834 GND.n8030 GND.n8027 4.74817
R26835 GND.n8035 GND.n8032 4.74817
R26836 GND.n8040 GND.n8037 4.74817
R26837 GND.n8042 GND.n3873 4.74817
R26838 GND.n38 GND.n6 4.70093
R26839 GND.n85 GND.n84 4.70093
R26840 GND.t16 GND.n3946 4.68277
R26841 GND.t14 GND.n4293 4.68277
R26842 GND.t87 GND.n4504 4.68277
R26843 GND.n21 GND.n20 4.63843
R26844 GND.n29 GND.n28 4.63843
R26845 GND.n37 GND.n36 4.63843
R26846 GND.n61 GND.n60 4.63843
R26847 GND.n69 GND.n68 4.63843
R26848 GND.n77 GND.n76 4.63843
R26849 GND.n7597 GND.n4793 4.6132
R26850 GND.n8362 GND.n2185 4.6132
R26851 GND.n5551 GND.t197 4.34833
R26852 GND.t12 GND.n4139 4.34833
R26853 GND.n46 GND.n42 4.05608
R26854 GND.n5240 GND.n5237 4.01388
R26855 GND.n8071 GND.n3832 4.01388
R26856 GND.n7987 GND.n3916 4.01388
R26857 GND.n5362 GND.n5361 4.01388
R26858 GND.n5457 GND.n4978 4.01388
R26859 GND.n7921 GND.n4024 4.01388
R26860 GND.n5560 GND.n4947 4.01388
R26861 GND.n7866 GND.n4129 4.01388
R26862 GND.n5664 GND.n4915 4.01388
R26863 GND.n7811 GND.n4233 4.01388
R26864 GND.n5761 GND.n4882 4.01388
R26865 GND.n7756 GND.n4336 4.01388
R26866 GND.n4404 GND.n4398 4.01388
R26867 GND.n7698 GND.n7697 4.01388
R26868 GND.n7656 GND.t58 4.01388
R26869 GND.n5888 GND.n5884 3.54314
R26870 GND.n8460 GND.n2145 3.54314
R26871 GND.n46 GND.n45 3.53792
R26872 GND.t155 GND.n3906 3.34498
R26873 GND.t15 GND.n4346 3.34498
R26874 GND.t35 GND.t16 3.01053
R26875 GND.t206 GND.t14 3.01053
R26876 GND.n5884 GND.n5873 2.87993
R26877 GND.n2145 GND.n2131 2.87993
R26878 GND.n3770 GND.n3751 2.67609
R26879 GND.n8120 GND.t150 2.67609
R26880 GND.n3804 GND.n3798 2.67609
R26881 GND.n7993 GND.n3906 2.67609
R26882 GND.n5412 GND.n5411 2.67609
R26883 GND.n7915 GND.n4034 2.67609
R26884 GND.n5551 GND.n5542 2.67609
R26885 GND.n7860 GND.n4139 2.67609
R26886 GND.n5655 GND.n5646 2.67609
R26887 GND.n5752 GND.n5743 2.67609
R26888 GND.n7750 GND.n4346 2.67609
R26889 GND.n7691 GND.n4432 2.67609
R26890 GND.n7665 GND.t153 2.67609
R26891 GND.n4722 GND.n4650 2.67609
R26892 GND.n2845 GND.t171 2.34164
R26893 GND.n8192 GND.t22 2.34164
R26894 GND.n7463 GND.t2 2.34164
R26895 GND.n7226 GND.t20 2.34164
R26896 GND.n5890 GND.n5873 2.27742
R26897 GND.n5895 GND.n5873 2.27742
R26898 GND.n5900 GND.n5873 2.27742
R26899 GND.n5905 GND.n5873 2.27742
R26900 GND.n5910 GND.n5873 2.27742
R26901 GND.n5915 GND.n5873 2.27742
R26902 GND.n5872 GND.n4842 2.27742
R26903 GND.n5872 GND.n4840 2.27742
R26904 GND.n5872 GND.n4839 2.27742
R26905 GND.n5872 GND.n4838 2.27742
R26906 GND.n5872 GND.n4837 2.27742
R26907 GND.n5872 GND.n4836 2.27742
R26908 GND.n5872 GND.n4835 2.27742
R26909 GND.n11107 GND.n106 2.27742
R26910 GND.n11107 GND.n104 2.27742
R26911 GND.n11108 GND.n11107 2.27742
R26912 GND.n11107 GND.n103 2.27742
R26913 GND.n3494 GND.n3493 2.27742
R26914 GND.n3494 GND.n2495 2.27742
R26915 GND.n3494 GND.n2494 2.27742
R26916 GND.n3494 GND.n2493 2.27742
R26917 GND.n3482 GND.n2492 2.27742
R26918 GND.n2534 GND.n2492 2.27742
R26919 GND.n3466 GND.n2492 2.27742
R26920 GND.n2536 GND.n2492 2.27742
R26921 GND.n6644 GND.n102 2.27742
R26922 GND.n7329 GND.n102 2.27742
R26923 GND.n6263 GND.n102 2.27742
R26924 GND.n7322 GND.n102 2.27742
R26925 GND.n6281 GND.n102 2.27742
R26926 GND.n3061 GND.n2492 2.27742
R26927 GND.n8477 GND.n2131 2.27742
R26928 GND.n8474 GND.n2131 2.27742
R26929 GND.n8471 GND.n2131 2.27742
R26930 GND.n8468 GND.n2131 2.27742
R26931 GND.n8465 GND.n2131 2.27742
R26932 GND.n8462 GND.n2131 2.27742
R26933 GND.n8043 GND.n8010 2.27742
R26934 GND.n8043 GND.n8017 2.27742
R26935 GND.n8043 GND.n8022 2.27742
R26936 GND.n8043 GND.n8027 2.27742
R26937 GND.n8043 GND.n8032 2.27742
R26938 GND.n8043 GND.n8037 2.27742
R26939 GND.n8043 GND.n8042 2.27742
R26940 GND GND.n39 2.17817
R26941 GND.n5224 GND.t130 2.00719
R26942 GND.n8064 GND.t10 2.00719
R26943 GND.n4463 GND.t156 2.00719
R26944 GND.n7683 GND.t50 2.00719
R26945 GND.n13 GND.n12 1.86544
R26946 GND.n12 GND.n10 1.86544
R26947 GND.n10 GND.n8 1.86544
R26948 GND.n20 GND.n19 1.86544
R26949 GND.n19 GND.n17 1.86544
R26950 GND.n17 GND.n15 1.86544
R26951 GND.n28 GND.n27 1.86544
R26952 GND.n27 GND.n25 1.86544
R26953 GND.n25 GND.n23 1.86544
R26954 GND.n36 GND.n35 1.86544
R26955 GND.n35 GND.n33 1.86544
R26956 GND.n33 GND.n31 1.86544
R26957 GND.n6 GND.n5 1.86544
R26958 GND.n5 GND.n3 1.86544
R26959 GND.n3 GND.n1 1.86544
R26960 GND.n50 GND.n48 1.86544
R26961 GND.n52 GND.n50 1.86544
R26962 GND.n53 GND.n52 1.86544
R26963 GND.n57 GND.n55 1.86544
R26964 GND.n59 GND.n57 1.86544
R26965 GND.n60 GND.n59 1.86544
R26966 GND.n65 GND.n63 1.86544
R26967 GND.n67 GND.n65 1.86544
R26968 GND.n68 GND.n67 1.86544
R26969 GND.n73 GND.n71 1.86544
R26970 GND.n75 GND.n73 1.86544
R26971 GND.n76 GND.n75 1.86544
R26972 GND.n81 GND.n79 1.86544
R26973 GND.n83 GND.n81 1.86544
R26974 GND.n84 GND.n83 1.86544
R26975 GND.n3296 GND.t0 1.67274
R26976 GND.n3639 GND.t191 1.67274
R26977 GND.n5397 GND.t6 1.67274
R26978 GND.n7805 GND.t33 1.67274
R26979 GND.n6873 GND.t27 1.67274
R26980 GND.n11020 GND.t29 1.67274
R26981 GND.n11117 GND.n11116 1.63939
R26982 GND.n38 GND.n37 1.36832
R26983 GND.n85 GND.n77 1.36832
R26984 GND.n5214 GND.n5211 1.33829
R26985 GND.n5227 GND.n5224 1.33829
R26986 GND.n8057 GND.n3850 1.33829
R26987 GND.n7999 GND.n3895 1.33829
R26988 GND.n5421 GND.n4997 1.33829
R26989 GND.n5439 GND.n4987 1.33829
R26990 GND.n7909 GND.n4044 1.33829
R26991 GND.n4071 GND.n4065 1.33829
R26992 GND.n7854 GND.n4149 1.33829
R26993 GND.n4176 GND.n4170 1.33829
R26994 GND.n7799 GND.n4251 1.33829
R26995 GND.n4278 GND.n4272 1.33829
R26996 GND.n7744 GND.n4355 1.33829
R26997 GND.n4385 GND.n4382 1.33829
R26998 GND.n7684 GND.n7683 1.33829
R26999 GND.n4514 GND.n4505 1.33829
R27000 GND.n4664 GND.n4663 1.24928
R27001 GND.n5150 GND.n5149 1.24928
R27002 GND.n5133 GND.n5132 1.24928
R27003 GND.n4782 GND.n4781 1.24928
R27004 GND.n29 GND.n21 1.02924
R27005 GND.n37 GND.n29 1.02924
R27006 GND.n69 GND.n61 1.02924
R27007 GND.n77 GND.n69 1.02924
R27008 GND.n3367 GND.t41 1.00384
R27009 GND.n3565 GND.t25 1.00384
R27010 GND.n3749 GND.n3739 1.00384
R27011 GND.n5448 GND.t6 1.00384
R27012 GND.n5697 GND.t33 1.00384
R27013 GND.n7657 GND.n7656 1.00384
R27014 GND.n7385 GND.t157 1.00384
R27015 GND.n7062 GND.t38 1.00384
R27016 GND.n8454 GND.n2185 0.970197
R27017 GND.n7597 GND.n7596 0.970197
R27018 GND.n8015 GND.n3875 0.970197
R27019 GND.n5864 GND.n5863 0.970197
R27020 GND.n41 GND.n40 0.831895
R27021 GND.n42 GND.n41 0.831895
R27022 GND.n44 GND.n43 0.831895
R27023 GND.n45 GND.n44 0.831895
R27024 GND.n4643 GND.n4637 0.776258
R27025 GND.n8127 GND.t111 0.669396
R27026 GND.t10 GND.n8063 0.669396
R27027 GND.t168 GND.n7890 0.669396
R27028 GND.n5607 GND.t210 0.669396
R27029 GND.t156 GND.n4460 0.669396
R27030 GND.n9049 GND.n9048 0.495927
R27031 GND.n10388 GND.n661 0.495927
R27032 GND.n10531 GND.n10530 0.495927
R27033 GND.n1581 GND.n1580 0.495927
R27034 GND.n5814 GND.n5813 0.492878
R27035 GND.n5026 GND.n3865 0.492878
R27036 GND.n3898 GND.n3874 0.492878
R27037 GND.n4834 GND.n4833 0.492878
R27038 GND.n10719 GND.n443 0.477634
R27039 GND.n5923 GND.n4606 0.477634
R27040 GND.n8311 GND.n8308 0.477634
R27041 GND.n1825 GND.n1729 0.477634
R27042 GND.n10901 GND.n10900 0.468488
R27043 GND.n2951 GND.n2950 0.468488
R27044 GND.n11107 GND.n102 0.429375
R27045 GND.n3494 GND.n2492 0.429375
R27046 GND.n3430 GND.t159 0.334948
R27047 GND.n2488 GND.t175 0.334948
R27048 GND.n6970 GND.t4 0.334948
R27049 GND.n11098 GND.t17 0.334948
R27050 GND.n4791 GND.n4634 0.312695
R27051 GND.n5142 GND.n5141 0.312695
R27052 GND.n5141 GND.n5140 0.312695
R27053 GND.n4791 GND.n4789 0.312695
R27054 GND.n10786 GND.n451 0.273366
R27055 GND.n7537 GND.n7536 0.273366
R27056 GND.n8704 GND.n8703 0.273366
R27057 GND.n8410 GND.n2122 0.273366
R27058 GND GND.n11117 0.271847
R27059 GND.n8300 GND.n2131 0.267268
R27060 GND.n6739 GND.n5873 0.267268
R27061 GND.n10655 GND.n451 0.264219
R27062 GND.n8703 GND.n8702 0.264219
R27063 GND.n11117 GND.n46 0.232523
R27064 GND.n4793 GND.n4633 0.229039
R27065 GND.n4796 GND.n4793 0.229039
R27066 GND.n8362 GND.n8361 0.229039
R27067 GND.n8453 GND.n8362 0.229039
R27068 GND.n5873 GND.n5872 0.207661
R27069 GND.n8043 GND.n2131 0.207661
R27070 GND.n8432 GND.n8384 0.194439
R27071 GND.n7567 GND.n4812 0.194439
R27072 GND.n10816 GND.n10767 0.194439
R27073 GND.n10847 GND.n10750 0.194439
R27074 GND.n8765 GND.n1761 0.194439
R27075 GND.n8734 GND.n1778 0.194439
R27076 GND.n3448 GND.n2653 0.152939
R27077 GND.n3449 GND.n3448 0.152939
R27078 GND.n3450 GND.n3449 0.152939
R27079 GND.n3450 GND.n2480 0.152939
R27080 GND.n3503 GND.n2480 0.152939
R27081 GND.n3504 GND.n3503 0.152939
R27082 GND.n3505 GND.n3504 0.152939
R27083 GND.n3506 GND.n3505 0.152939
R27084 GND.n3506 GND.n2458 0.152939
R27085 GND.n3529 GND.n2458 0.152939
R27086 GND.n3530 GND.n3529 0.152939
R27087 GND.n3531 GND.n3530 0.152939
R27088 GND.n3532 GND.n3531 0.152939
R27089 GND.n3532 GND.n2437 0.152939
R27090 GND.n3555 GND.n2437 0.152939
R27091 GND.n3556 GND.n3555 0.152939
R27092 GND.n3557 GND.n3556 0.152939
R27093 GND.n3558 GND.n3557 0.152939
R27094 GND.n3558 GND.n2416 0.152939
R27095 GND.n3581 GND.n2416 0.152939
R27096 GND.n3582 GND.n3581 0.152939
R27097 GND.n3583 GND.n3582 0.152939
R27098 GND.n3584 GND.n3583 0.152939
R27099 GND.n3584 GND.n2393 0.152939
R27100 GND.n3606 GND.n2393 0.152939
R27101 GND.n3607 GND.n3606 0.152939
R27102 GND.n3608 GND.n3607 0.152939
R27103 GND.n3609 GND.n3608 0.152939
R27104 GND.n3609 GND.n2373 0.152939
R27105 GND.n3632 GND.n2373 0.152939
R27106 GND.n3633 GND.n3632 0.152939
R27107 GND.n3634 GND.n3633 0.152939
R27108 GND.n3635 GND.n3634 0.152939
R27109 GND.n3635 GND.n2353 0.152939
R27110 GND.n3658 GND.n2353 0.152939
R27111 GND.n3659 GND.n3658 0.152939
R27112 GND.n3660 GND.n3659 0.152939
R27113 GND.n3661 GND.n3660 0.152939
R27114 GND.n3661 GND.n2331 0.152939
R27115 GND.n3684 GND.n2331 0.152939
R27116 GND.n3685 GND.n3684 0.152939
R27117 GND.n3686 GND.n3685 0.152939
R27118 GND.n3687 GND.n3686 0.152939
R27119 GND.n3687 GND.n2304 0.152939
R27120 GND.n8195 GND.n2304 0.152939
R27121 GND.n8196 GND.n8195 0.152939
R27122 GND.n8197 GND.n8196 0.152939
R27123 GND.n8198 GND.n8197 0.152939
R27124 GND.n8198 GND.n2282 0.152939
R27125 GND.n8221 GND.n2282 0.152939
R27126 GND.n8222 GND.n8221 0.152939
R27127 GND.n8223 GND.n8222 0.152939
R27128 GND.n8224 GND.n8223 0.152939
R27129 GND.n8224 GND.n2261 0.152939
R27130 GND.n8247 GND.n2261 0.152939
R27131 GND.n8248 GND.n8247 0.152939
R27132 GND.n8249 GND.n8248 0.152939
R27133 GND.n8250 GND.n8249 0.152939
R27134 GND.n8250 GND.n2240 0.152939
R27135 GND.n8273 GND.n2240 0.152939
R27136 GND.n8274 GND.n8273 0.152939
R27137 GND.n8275 GND.n8274 0.152939
R27138 GND.n8276 GND.n8275 0.152939
R27139 GND.n8276 GND.n2217 0.152939
R27140 GND.n8297 GND.n2217 0.152939
R27141 GND.n8298 GND.n8297 0.152939
R27142 GND.n8299 GND.n8298 0.152939
R27143 GND.n8300 GND.n8299 0.152939
R27144 GND.n9049 GND.n1458 0.152939
R27145 GND.n9057 GND.n1458 0.152939
R27146 GND.n9058 GND.n9057 0.152939
R27147 GND.n9059 GND.n9058 0.152939
R27148 GND.n9059 GND.n1452 0.152939
R27149 GND.n9067 GND.n1452 0.152939
R27150 GND.n9068 GND.n9067 0.152939
R27151 GND.n9069 GND.n9068 0.152939
R27152 GND.n9069 GND.n1446 0.152939
R27153 GND.n9077 GND.n1446 0.152939
R27154 GND.n9078 GND.n9077 0.152939
R27155 GND.n9079 GND.n9078 0.152939
R27156 GND.n9079 GND.n1440 0.152939
R27157 GND.n9087 GND.n1440 0.152939
R27158 GND.n9088 GND.n9087 0.152939
R27159 GND.n9089 GND.n9088 0.152939
R27160 GND.n9089 GND.n1434 0.152939
R27161 GND.n9097 GND.n1434 0.152939
R27162 GND.n9098 GND.n9097 0.152939
R27163 GND.n9099 GND.n9098 0.152939
R27164 GND.n9099 GND.n1428 0.152939
R27165 GND.n9107 GND.n1428 0.152939
R27166 GND.n9108 GND.n9107 0.152939
R27167 GND.n9109 GND.n9108 0.152939
R27168 GND.n9109 GND.n1422 0.152939
R27169 GND.n9117 GND.n1422 0.152939
R27170 GND.n9118 GND.n9117 0.152939
R27171 GND.n9119 GND.n9118 0.152939
R27172 GND.n9119 GND.n1416 0.152939
R27173 GND.n9127 GND.n1416 0.152939
R27174 GND.n9128 GND.n9127 0.152939
R27175 GND.n9129 GND.n9128 0.152939
R27176 GND.n9129 GND.n1410 0.152939
R27177 GND.n9137 GND.n1410 0.152939
R27178 GND.n9138 GND.n9137 0.152939
R27179 GND.n9139 GND.n9138 0.152939
R27180 GND.n9139 GND.n1404 0.152939
R27181 GND.n9147 GND.n1404 0.152939
R27182 GND.n9148 GND.n9147 0.152939
R27183 GND.n9149 GND.n9148 0.152939
R27184 GND.n9149 GND.n1398 0.152939
R27185 GND.n9157 GND.n1398 0.152939
R27186 GND.n9158 GND.n9157 0.152939
R27187 GND.n9159 GND.n9158 0.152939
R27188 GND.n9159 GND.n1392 0.152939
R27189 GND.n9167 GND.n1392 0.152939
R27190 GND.n9168 GND.n9167 0.152939
R27191 GND.n9169 GND.n9168 0.152939
R27192 GND.n9169 GND.n1386 0.152939
R27193 GND.n9177 GND.n1386 0.152939
R27194 GND.n9178 GND.n9177 0.152939
R27195 GND.n9179 GND.n9178 0.152939
R27196 GND.n9179 GND.n1380 0.152939
R27197 GND.n9187 GND.n1380 0.152939
R27198 GND.n9188 GND.n9187 0.152939
R27199 GND.n9189 GND.n9188 0.152939
R27200 GND.n9189 GND.n1374 0.152939
R27201 GND.n9197 GND.n1374 0.152939
R27202 GND.n9198 GND.n9197 0.152939
R27203 GND.n9199 GND.n9198 0.152939
R27204 GND.n9199 GND.n1368 0.152939
R27205 GND.n9207 GND.n1368 0.152939
R27206 GND.n9208 GND.n9207 0.152939
R27207 GND.n9209 GND.n9208 0.152939
R27208 GND.n9209 GND.n1362 0.152939
R27209 GND.n9217 GND.n1362 0.152939
R27210 GND.n9218 GND.n9217 0.152939
R27211 GND.n9219 GND.n9218 0.152939
R27212 GND.n9219 GND.n1356 0.152939
R27213 GND.n9227 GND.n1356 0.152939
R27214 GND.n9228 GND.n9227 0.152939
R27215 GND.n9229 GND.n9228 0.152939
R27216 GND.n9229 GND.n1350 0.152939
R27217 GND.n9237 GND.n1350 0.152939
R27218 GND.n9238 GND.n9237 0.152939
R27219 GND.n9239 GND.n9238 0.152939
R27220 GND.n9239 GND.n1344 0.152939
R27221 GND.n9247 GND.n1344 0.152939
R27222 GND.n9248 GND.n9247 0.152939
R27223 GND.n9249 GND.n9248 0.152939
R27224 GND.n9249 GND.n1338 0.152939
R27225 GND.n9257 GND.n1338 0.152939
R27226 GND.n9258 GND.n9257 0.152939
R27227 GND.n9259 GND.n9258 0.152939
R27228 GND.n9259 GND.n1332 0.152939
R27229 GND.n9267 GND.n1332 0.152939
R27230 GND.n9268 GND.n9267 0.152939
R27231 GND.n9269 GND.n9268 0.152939
R27232 GND.n9269 GND.n1326 0.152939
R27233 GND.n9277 GND.n1326 0.152939
R27234 GND.n9278 GND.n9277 0.152939
R27235 GND.n9279 GND.n9278 0.152939
R27236 GND.n9279 GND.n1320 0.152939
R27237 GND.n9287 GND.n1320 0.152939
R27238 GND.n9288 GND.n9287 0.152939
R27239 GND.n9289 GND.n9288 0.152939
R27240 GND.n9289 GND.n1314 0.152939
R27241 GND.n9297 GND.n1314 0.152939
R27242 GND.n9298 GND.n9297 0.152939
R27243 GND.n9299 GND.n9298 0.152939
R27244 GND.n9299 GND.n1308 0.152939
R27245 GND.n9307 GND.n1308 0.152939
R27246 GND.n9308 GND.n9307 0.152939
R27247 GND.n9309 GND.n9308 0.152939
R27248 GND.n9309 GND.n1302 0.152939
R27249 GND.n9317 GND.n1302 0.152939
R27250 GND.n9318 GND.n9317 0.152939
R27251 GND.n9319 GND.n9318 0.152939
R27252 GND.n9319 GND.n1296 0.152939
R27253 GND.n9327 GND.n1296 0.152939
R27254 GND.n9328 GND.n9327 0.152939
R27255 GND.n9329 GND.n9328 0.152939
R27256 GND.n9329 GND.n1290 0.152939
R27257 GND.n9337 GND.n1290 0.152939
R27258 GND.n9338 GND.n9337 0.152939
R27259 GND.n9339 GND.n9338 0.152939
R27260 GND.n9339 GND.n1284 0.152939
R27261 GND.n9347 GND.n1284 0.152939
R27262 GND.n9348 GND.n9347 0.152939
R27263 GND.n9349 GND.n9348 0.152939
R27264 GND.n9349 GND.n1278 0.152939
R27265 GND.n9357 GND.n1278 0.152939
R27266 GND.n9358 GND.n9357 0.152939
R27267 GND.n9359 GND.n9358 0.152939
R27268 GND.n9359 GND.n1272 0.152939
R27269 GND.n9367 GND.n1272 0.152939
R27270 GND.n9368 GND.n9367 0.152939
R27271 GND.n9369 GND.n9368 0.152939
R27272 GND.n9369 GND.n1266 0.152939
R27273 GND.n9377 GND.n1266 0.152939
R27274 GND.n9378 GND.n9377 0.152939
R27275 GND.n9379 GND.n9378 0.152939
R27276 GND.n9379 GND.n1260 0.152939
R27277 GND.n9387 GND.n1260 0.152939
R27278 GND.n9388 GND.n9387 0.152939
R27279 GND.n9389 GND.n9388 0.152939
R27280 GND.n9389 GND.n1254 0.152939
R27281 GND.n9397 GND.n1254 0.152939
R27282 GND.n9398 GND.n9397 0.152939
R27283 GND.n9399 GND.n9398 0.152939
R27284 GND.n9399 GND.n1248 0.152939
R27285 GND.n9407 GND.n1248 0.152939
R27286 GND.n9408 GND.n9407 0.152939
R27287 GND.n9409 GND.n9408 0.152939
R27288 GND.n9409 GND.n1242 0.152939
R27289 GND.n9417 GND.n1242 0.152939
R27290 GND.n9418 GND.n9417 0.152939
R27291 GND.n9419 GND.n9418 0.152939
R27292 GND.n9419 GND.n1236 0.152939
R27293 GND.n9427 GND.n1236 0.152939
R27294 GND.n9428 GND.n9427 0.152939
R27295 GND.n9429 GND.n9428 0.152939
R27296 GND.n9429 GND.n1230 0.152939
R27297 GND.n9437 GND.n1230 0.152939
R27298 GND.n9438 GND.n9437 0.152939
R27299 GND.n9439 GND.n9438 0.152939
R27300 GND.n9439 GND.n1224 0.152939
R27301 GND.n9447 GND.n1224 0.152939
R27302 GND.n9448 GND.n9447 0.152939
R27303 GND.n9449 GND.n9448 0.152939
R27304 GND.n9449 GND.n1218 0.152939
R27305 GND.n9457 GND.n1218 0.152939
R27306 GND.n9458 GND.n9457 0.152939
R27307 GND.n9459 GND.n9458 0.152939
R27308 GND.n9459 GND.n1212 0.152939
R27309 GND.n9467 GND.n1212 0.152939
R27310 GND.n9468 GND.n9467 0.152939
R27311 GND.n9469 GND.n9468 0.152939
R27312 GND.n9469 GND.n1206 0.152939
R27313 GND.n9477 GND.n1206 0.152939
R27314 GND.n9478 GND.n9477 0.152939
R27315 GND.n9479 GND.n9478 0.152939
R27316 GND.n9479 GND.n1200 0.152939
R27317 GND.n9487 GND.n1200 0.152939
R27318 GND.n9488 GND.n9487 0.152939
R27319 GND.n9489 GND.n9488 0.152939
R27320 GND.n9489 GND.n1194 0.152939
R27321 GND.n9497 GND.n1194 0.152939
R27322 GND.n9498 GND.n9497 0.152939
R27323 GND.n9499 GND.n9498 0.152939
R27324 GND.n9499 GND.n1188 0.152939
R27325 GND.n9507 GND.n1188 0.152939
R27326 GND.n9508 GND.n9507 0.152939
R27327 GND.n9509 GND.n9508 0.152939
R27328 GND.n9509 GND.n1182 0.152939
R27329 GND.n9517 GND.n1182 0.152939
R27330 GND.n9518 GND.n9517 0.152939
R27331 GND.n9519 GND.n9518 0.152939
R27332 GND.n9519 GND.n1176 0.152939
R27333 GND.n9527 GND.n1176 0.152939
R27334 GND.n9528 GND.n9527 0.152939
R27335 GND.n9529 GND.n9528 0.152939
R27336 GND.n9529 GND.n1170 0.152939
R27337 GND.n9537 GND.n1170 0.152939
R27338 GND.n9538 GND.n9537 0.152939
R27339 GND.n9539 GND.n9538 0.152939
R27340 GND.n9539 GND.n1164 0.152939
R27341 GND.n9547 GND.n1164 0.152939
R27342 GND.n9548 GND.n9547 0.152939
R27343 GND.n9549 GND.n9548 0.152939
R27344 GND.n9549 GND.n1158 0.152939
R27345 GND.n9557 GND.n1158 0.152939
R27346 GND.n9558 GND.n9557 0.152939
R27347 GND.n9559 GND.n9558 0.152939
R27348 GND.n9559 GND.n1152 0.152939
R27349 GND.n9567 GND.n1152 0.152939
R27350 GND.n9568 GND.n9567 0.152939
R27351 GND.n9569 GND.n9568 0.152939
R27352 GND.n9569 GND.n1146 0.152939
R27353 GND.n9577 GND.n1146 0.152939
R27354 GND.n9578 GND.n9577 0.152939
R27355 GND.n9579 GND.n9578 0.152939
R27356 GND.n9579 GND.n1140 0.152939
R27357 GND.n9587 GND.n1140 0.152939
R27358 GND.n9588 GND.n9587 0.152939
R27359 GND.n9589 GND.n9588 0.152939
R27360 GND.n9589 GND.n1134 0.152939
R27361 GND.n9597 GND.n1134 0.152939
R27362 GND.n9598 GND.n9597 0.152939
R27363 GND.n9599 GND.n9598 0.152939
R27364 GND.n9599 GND.n1128 0.152939
R27365 GND.n9607 GND.n1128 0.152939
R27366 GND.n9608 GND.n9607 0.152939
R27367 GND.n9609 GND.n9608 0.152939
R27368 GND.n9609 GND.n1122 0.152939
R27369 GND.n9617 GND.n1122 0.152939
R27370 GND.n9618 GND.n9617 0.152939
R27371 GND.n9619 GND.n9618 0.152939
R27372 GND.n9619 GND.n1116 0.152939
R27373 GND.n9627 GND.n1116 0.152939
R27374 GND.n9628 GND.n9627 0.152939
R27375 GND.n9629 GND.n9628 0.152939
R27376 GND.n9629 GND.n1110 0.152939
R27377 GND.n9637 GND.n1110 0.152939
R27378 GND.n9638 GND.n9637 0.152939
R27379 GND.n9639 GND.n9638 0.152939
R27380 GND.n9639 GND.n1104 0.152939
R27381 GND.n9647 GND.n1104 0.152939
R27382 GND.n9648 GND.n9647 0.152939
R27383 GND.n9649 GND.n9648 0.152939
R27384 GND.n9649 GND.n1098 0.152939
R27385 GND.n9657 GND.n1098 0.152939
R27386 GND.n9658 GND.n9657 0.152939
R27387 GND.n9659 GND.n9658 0.152939
R27388 GND.n9659 GND.n1092 0.152939
R27389 GND.n9667 GND.n1092 0.152939
R27390 GND.n9668 GND.n9667 0.152939
R27391 GND.n9669 GND.n9668 0.152939
R27392 GND.n9669 GND.n1086 0.152939
R27393 GND.n9677 GND.n1086 0.152939
R27394 GND.n9678 GND.n9677 0.152939
R27395 GND.n9679 GND.n9678 0.152939
R27396 GND.n9679 GND.n1080 0.152939
R27397 GND.n9687 GND.n1080 0.152939
R27398 GND.n9688 GND.n9687 0.152939
R27399 GND.n9689 GND.n9688 0.152939
R27400 GND.n9689 GND.n1074 0.152939
R27401 GND.n9697 GND.n1074 0.152939
R27402 GND.n9698 GND.n9697 0.152939
R27403 GND.n9699 GND.n9698 0.152939
R27404 GND.n9699 GND.n1068 0.152939
R27405 GND.n9707 GND.n1068 0.152939
R27406 GND.n9708 GND.n9707 0.152939
R27407 GND.n9709 GND.n9708 0.152939
R27408 GND.n9709 GND.n1062 0.152939
R27409 GND.n9717 GND.n1062 0.152939
R27410 GND.n9718 GND.n9717 0.152939
R27411 GND.n9719 GND.n9718 0.152939
R27412 GND.n9719 GND.n1056 0.152939
R27413 GND.n9727 GND.n1056 0.152939
R27414 GND.n9728 GND.n9727 0.152939
R27415 GND.n9729 GND.n9728 0.152939
R27416 GND.n9729 GND.n1050 0.152939
R27417 GND.n9737 GND.n1050 0.152939
R27418 GND.n9738 GND.n9737 0.152939
R27419 GND.n9739 GND.n9738 0.152939
R27420 GND.n9739 GND.n1044 0.152939
R27421 GND.n9747 GND.n1044 0.152939
R27422 GND.n9748 GND.n9747 0.152939
R27423 GND.n9749 GND.n9748 0.152939
R27424 GND.n9749 GND.n1038 0.152939
R27425 GND.n9757 GND.n1038 0.152939
R27426 GND.n9758 GND.n9757 0.152939
R27427 GND.n9759 GND.n9758 0.152939
R27428 GND.n9759 GND.n1032 0.152939
R27429 GND.n9767 GND.n1032 0.152939
R27430 GND.n9768 GND.n9767 0.152939
R27431 GND.n9769 GND.n9768 0.152939
R27432 GND.n9769 GND.n1026 0.152939
R27433 GND.n9777 GND.n1026 0.152939
R27434 GND.n9778 GND.n9777 0.152939
R27435 GND.n9779 GND.n9778 0.152939
R27436 GND.n9779 GND.n1020 0.152939
R27437 GND.n9787 GND.n1020 0.152939
R27438 GND.n9788 GND.n9787 0.152939
R27439 GND.n9789 GND.n9788 0.152939
R27440 GND.n9789 GND.n1014 0.152939
R27441 GND.n9797 GND.n1014 0.152939
R27442 GND.n9798 GND.n9797 0.152939
R27443 GND.n9799 GND.n9798 0.152939
R27444 GND.n9799 GND.n1008 0.152939
R27445 GND.n9807 GND.n1008 0.152939
R27446 GND.n9808 GND.n9807 0.152939
R27447 GND.n9809 GND.n9808 0.152939
R27448 GND.n9809 GND.n1002 0.152939
R27449 GND.n9817 GND.n1002 0.152939
R27450 GND.n9818 GND.n9817 0.152939
R27451 GND.n9819 GND.n9818 0.152939
R27452 GND.n9819 GND.n996 0.152939
R27453 GND.n9827 GND.n996 0.152939
R27454 GND.n9828 GND.n9827 0.152939
R27455 GND.n9829 GND.n9828 0.152939
R27456 GND.n9829 GND.n990 0.152939
R27457 GND.n9837 GND.n990 0.152939
R27458 GND.n9838 GND.n9837 0.152939
R27459 GND.n9839 GND.n9838 0.152939
R27460 GND.n9839 GND.n984 0.152939
R27461 GND.n9847 GND.n984 0.152939
R27462 GND.n9848 GND.n9847 0.152939
R27463 GND.n9849 GND.n9848 0.152939
R27464 GND.n9849 GND.n978 0.152939
R27465 GND.n9857 GND.n978 0.152939
R27466 GND.n9858 GND.n9857 0.152939
R27467 GND.n9859 GND.n9858 0.152939
R27468 GND.n9859 GND.n972 0.152939
R27469 GND.n9867 GND.n972 0.152939
R27470 GND.n9868 GND.n9867 0.152939
R27471 GND.n9869 GND.n9868 0.152939
R27472 GND.n9869 GND.n966 0.152939
R27473 GND.n9877 GND.n966 0.152939
R27474 GND.n9878 GND.n9877 0.152939
R27475 GND.n9879 GND.n9878 0.152939
R27476 GND.n9879 GND.n960 0.152939
R27477 GND.n9887 GND.n960 0.152939
R27478 GND.n9888 GND.n9887 0.152939
R27479 GND.n9889 GND.n9888 0.152939
R27480 GND.n9889 GND.n954 0.152939
R27481 GND.n9897 GND.n954 0.152939
R27482 GND.n9898 GND.n9897 0.152939
R27483 GND.n9899 GND.n9898 0.152939
R27484 GND.n9899 GND.n948 0.152939
R27485 GND.n9907 GND.n948 0.152939
R27486 GND.n9908 GND.n9907 0.152939
R27487 GND.n9909 GND.n9908 0.152939
R27488 GND.n9909 GND.n942 0.152939
R27489 GND.n9917 GND.n942 0.152939
R27490 GND.n9918 GND.n9917 0.152939
R27491 GND.n9919 GND.n9918 0.152939
R27492 GND.n9919 GND.n936 0.152939
R27493 GND.n9927 GND.n936 0.152939
R27494 GND.n9928 GND.n9927 0.152939
R27495 GND.n9929 GND.n9928 0.152939
R27496 GND.n9929 GND.n930 0.152939
R27497 GND.n9937 GND.n930 0.152939
R27498 GND.n9938 GND.n9937 0.152939
R27499 GND.n9939 GND.n9938 0.152939
R27500 GND.n9939 GND.n924 0.152939
R27501 GND.n9947 GND.n924 0.152939
R27502 GND.n9948 GND.n9947 0.152939
R27503 GND.n9949 GND.n9948 0.152939
R27504 GND.n9949 GND.n918 0.152939
R27505 GND.n9957 GND.n918 0.152939
R27506 GND.n9958 GND.n9957 0.152939
R27507 GND.n9959 GND.n9958 0.152939
R27508 GND.n9959 GND.n912 0.152939
R27509 GND.n9967 GND.n912 0.152939
R27510 GND.n9968 GND.n9967 0.152939
R27511 GND.n9969 GND.n9968 0.152939
R27512 GND.n9969 GND.n906 0.152939
R27513 GND.n9977 GND.n906 0.152939
R27514 GND.n9978 GND.n9977 0.152939
R27515 GND.n9979 GND.n9978 0.152939
R27516 GND.n9979 GND.n900 0.152939
R27517 GND.n9987 GND.n900 0.152939
R27518 GND.n9988 GND.n9987 0.152939
R27519 GND.n9989 GND.n9988 0.152939
R27520 GND.n9989 GND.n894 0.152939
R27521 GND.n9997 GND.n894 0.152939
R27522 GND.n9998 GND.n9997 0.152939
R27523 GND.n9999 GND.n9998 0.152939
R27524 GND.n9999 GND.n888 0.152939
R27525 GND.n10007 GND.n888 0.152939
R27526 GND.n10008 GND.n10007 0.152939
R27527 GND.n10009 GND.n10008 0.152939
R27528 GND.n10009 GND.n882 0.152939
R27529 GND.n10017 GND.n882 0.152939
R27530 GND.n10018 GND.n10017 0.152939
R27531 GND.n10019 GND.n10018 0.152939
R27532 GND.n10019 GND.n876 0.152939
R27533 GND.n10027 GND.n876 0.152939
R27534 GND.n10028 GND.n10027 0.152939
R27535 GND.n10029 GND.n10028 0.152939
R27536 GND.n10029 GND.n870 0.152939
R27537 GND.n10037 GND.n870 0.152939
R27538 GND.n10038 GND.n10037 0.152939
R27539 GND.n10039 GND.n10038 0.152939
R27540 GND.n10039 GND.n864 0.152939
R27541 GND.n10047 GND.n864 0.152939
R27542 GND.n10048 GND.n10047 0.152939
R27543 GND.n10049 GND.n10048 0.152939
R27544 GND.n10049 GND.n858 0.152939
R27545 GND.n10057 GND.n858 0.152939
R27546 GND.n10058 GND.n10057 0.152939
R27547 GND.n10059 GND.n10058 0.152939
R27548 GND.n10059 GND.n852 0.152939
R27549 GND.n10067 GND.n852 0.152939
R27550 GND.n10068 GND.n10067 0.152939
R27551 GND.n10069 GND.n10068 0.152939
R27552 GND.n10069 GND.n846 0.152939
R27553 GND.n10077 GND.n846 0.152939
R27554 GND.n10078 GND.n10077 0.152939
R27555 GND.n10079 GND.n10078 0.152939
R27556 GND.n10079 GND.n840 0.152939
R27557 GND.n10087 GND.n840 0.152939
R27558 GND.n10088 GND.n10087 0.152939
R27559 GND.n10089 GND.n10088 0.152939
R27560 GND.n10089 GND.n834 0.152939
R27561 GND.n10097 GND.n834 0.152939
R27562 GND.n10098 GND.n10097 0.152939
R27563 GND.n10099 GND.n10098 0.152939
R27564 GND.n10099 GND.n828 0.152939
R27565 GND.n10107 GND.n828 0.152939
R27566 GND.n10108 GND.n10107 0.152939
R27567 GND.n10109 GND.n10108 0.152939
R27568 GND.n10109 GND.n822 0.152939
R27569 GND.n10117 GND.n822 0.152939
R27570 GND.n10118 GND.n10117 0.152939
R27571 GND.n10119 GND.n10118 0.152939
R27572 GND.n10119 GND.n816 0.152939
R27573 GND.n10127 GND.n816 0.152939
R27574 GND.n10128 GND.n10127 0.152939
R27575 GND.n10129 GND.n10128 0.152939
R27576 GND.n10129 GND.n810 0.152939
R27577 GND.n10137 GND.n810 0.152939
R27578 GND.n10138 GND.n10137 0.152939
R27579 GND.n10139 GND.n10138 0.152939
R27580 GND.n10139 GND.n804 0.152939
R27581 GND.n10147 GND.n804 0.152939
R27582 GND.n10148 GND.n10147 0.152939
R27583 GND.n10149 GND.n10148 0.152939
R27584 GND.n10149 GND.n798 0.152939
R27585 GND.n10157 GND.n798 0.152939
R27586 GND.n10158 GND.n10157 0.152939
R27587 GND.n10159 GND.n10158 0.152939
R27588 GND.n10159 GND.n792 0.152939
R27589 GND.n10167 GND.n792 0.152939
R27590 GND.n10168 GND.n10167 0.152939
R27591 GND.n10169 GND.n10168 0.152939
R27592 GND.n10169 GND.n786 0.152939
R27593 GND.n10177 GND.n786 0.152939
R27594 GND.n10178 GND.n10177 0.152939
R27595 GND.n10179 GND.n10178 0.152939
R27596 GND.n10179 GND.n780 0.152939
R27597 GND.n10187 GND.n780 0.152939
R27598 GND.n10188 GND.n10187 0.152939
R27599 GND.n10189 GND.n10188 0.152939
R27600 GND.n10189 GND.n774 0.152939
R27601 GND.n10197 GND.n774 0.152939
R27602 GND.n10198 GND.n10197 0.152939
R27603 GND.n10199 GND.n10198 0.152939
R27604 GND.n10199 GND.n768 0.152939
R27605 GND.n10207 GND.n768 0.152939
R27606 GND.n10208 GND.n10207 0.152939
R27607 GND.n10209 GND.n10208 0.152939
R27608 GND.n10209 GND.n762 0.152939
R27609 GND.n10217 GND.n762 0.152939
R27610 GND.n10218 GND.n10217 0.152939
R27611 GND.n10219 GND.n10218 0.152939
R27612 GND.n10219 GND.n756 0.152939
R27613 GND.n10227 GND.n756 0.152939
R27614 GND.n10228 GND.n10227 0.152939
R27615 GND.n10229 GND.n10228 0.152939
R27616 GND.n10229 GND.n750 0.152939
R27617 GND.n10237 GND.n750 0.152939
R27618 GND.n10238 GND.n10237 0.152939
R27619 GND.n10239 GND.n10238 0.152939
R27620 GND.n10239 GND.n744 0.152939
R27621 GND.n10247 GND.n744 0.152939
R27622 GND.n10248 GND.n10247 0.152939
R27623 GND.n10249 GND.n10248 0.152939
R27624 GND.n10249 GND.n738 0.152939
R27625 GND.n10257 GND.n738 0.152939
R27626 GND.n10258 GND.n10257 0.152939
R27627 GND.n10259 GND.n10258 0.152939
R27628 GND.n10259 GND.n732 0.152939
R27629 GND.n10267 GND.n732 0.152939
R27630 GND.n10268 GND.n10267 0.152939
R27631 GND.n10269 GND.n10268 0.152939
R27632 GND.n10269 GND.n726 0.152939
R27633 GND.n10277 GND.n726 0.152939
R27634 GND.n10278 GND.n10277 0.152939
R27635 GND.n10279 GND.n10278 0.152939
R27636 GND.n10279 GND.n720 0.152939
R27637 GND.n10287 GND.n720 0.152939
R27638 GND.n10288 GND.n10287 0.152939
R27639 GND.n10289 GND.n10288 0.152939
R27640 GND.n10289 GND.n714 0.152939
R27641 GND.n10297 GND.n714 0.152939
R27642 GND.n10298 GND.n10297 0.152939
R27643 GND.n10299 GND.n10298 0.152939
R27644 GND.n10299 GND.n708 0.152939
R27645 GND.n10307 GND.n708 0.152939
R27646 GND.n10308 GND.n10307 0.152939
R27647 GND.n10309 GND.n10308 0.152939
R27648 GND.n10309 GND.n702 0.152939
R27649 GND.n10317 GND.n702 0.152939
R27650 GND.n10318 GND.n10317 0.152939
R27651 GND.n10319 GND.n10318 0.152939
R27652 GND.n10319 GND.n696 0.152939
R27653 GND.n10327 GND.n696 0.152939
R27654 GND.n10328 GND.n10327 0.152939
R27655 GND.n10329 GND.n10328 0.152939
R27656 GND.n10329 GND.n690 0.152939
R27657 GND.n10337 GND.n690 0.152939
R27658 GND.n10338 GND.n10337 0.152939
R27659 GND.n10339 GND.n10338 0.152939
R27660 GND.n10339 GND.n684 0.152939
R27661 GND.n10347 GND.n684 0.152939
R27662 GND.n10348 GND.n10347 0.152939
R27663 GND.n10349 GND.n10348 0.152939
R27664 GND.n10349 GND.n678 0.152939
R27665 GND.n10357 GND.n678 0.152939
R27666 GND.n10358 GND.n10357 0.152939
R27667 GND.n10359 GND.n10358 0.152939
R27668 GND.n10359 GND.n672 0.152939
R27669 GND.n10367 GND.n672 0.152939
R27670 GND.n10368 GND.n10367 0.152939
R27671 GND.n10369 GND.n10368 0.152939
R27672 GND.n10369 GND.n666 0.152939
R27673 GND.n10377 GND.n666 0.152939
R27674 GND.n10378 GND.n10377 0.152939
R27675 GND.n10379 GND.n10378 0.152939
R27676 GND.n10379 GND.n661 0.152939
R27677 GND.n10389 GND.n10388 0.152939
R27678 GND.n10390 GND.n10389 0.152939
R27679 GND.n10390 GND.n655 0.152939
R27680 GND.n10398 GND.n655 0.152939
R27681 GND.n10399 GND.n10398 0.152939
R27682 GND.n10400 GND.n10399 0.152939
R27683 GND.n10400 GND.n649 0.152939
R27684 GND.n10408 GND.n649 0.152939
R27685 GND.n10409 GND.n10408 0.152939
R27686 GND.n10410 GND.n10409 0.152939
R27687 GND.n10410 GND.n643 0.152939
R27688 GND.n10418 GND.n643 0.152939
R27689 GND.n10419 GND.n10418 0.152939
R27690 GND.n10420 GND.n10419 0.152939
R27691 GND.n10420 GND.n637 0.152939
R27692 GND.n10428 GND.n637 0.152939
R27693 GND.n10429 GND.n10428 0.152939
R27694 GND.n10430 GND.n10429 0.152939
R27695 GND.n10430 GND.n631 0.152939
R27696 GND.n10438 GND.n631 0.152939
R27697 GND.n10439 GND.n10438 0.152939
R27698 GND.n10440 GND.n10439 0.152939
R27699 GND.n10440 GND.n625 0.152939
R27700 GND.n10448 GND.n625 0.152939
R27701 GND.n10449 GND.n10448 0.152939
R27702 GND.n10450 GND.n10449 0.152939
R27703 GND.n10450 GND.n619 0.152939
R27704 GND.n10458 GND.n619 0.152939
R27705 GND.n10459 GND.n10458 0.152939
R27706 GND.n10460 GND.n10459 0.152939
R27707 GND.n10460 GND.n613 0.152939
R27708 GND.n10468 GND.n613 0.152939
R27709 GND.n10469 GND.n10468 0.152939
R27710 GND.n10470 GND.n10469 0.152939
R27711 GND.n10470 GND.n607 0.152939
R27712 GND.n10478 GND.n607 0.152939
R27713 GND.n10479 GND.n10478 0.152939
R27714 GND.n10480 GND.n10479 0.152939
R27715 GND.n10480 GND.n601 0.152939
R27716 GND.n10488 GND.n601 0.152939
R27717 GND.n10489 GND.n10488 0.152939
R27718 GND.n10490 GND.n10489 0.152939
R27719 GND.n10490 GND.n595 0.152939
R27720 GND.n10498 GND.n595 0.152939
R27721 GND.n10499 GND.n10498 0.152939
R27722 GND.n10500 GND.n10499 0.152939
R27723 GND.n10500 GND.n589 0.152939
R27724 GND.n10508 GND.n589 0.152939
R27725 GND.n10509 GND.n10508 0.152939
R27726 GND.n10510 GND.n10509 0.152939
R27727 GND.n10510 GND.n583 0.152939
R27728 GND.n10518 GND.n583 0.152939
R27729 GND.n10519 GND.n10518 0.152939
R27730 GND.n10520 GND.n10519 0.152939
R27731 GND.n10520 GND.n577 0.152939
R27732 GND.n10528 GND.n577 0.152939
R27733 GND.n10529 GND.n10528 0.152939
R27734 GND.n10531 GND.n10529 0.152939
R27735 GND.n6283 GND.n102 0.152939
R27736 GND.n6284 GND.n6283 0.152939
R27737 GND.n6285 GND.n6284 0.152939
R27738 GND.n6288 GND.n6285 0.152939
R27739 GND.n6289 GND.n6288 0.152939
R27740 GND.n6290 GND.n6289 0.152939
R27741 GND.n6291 GND.n6290 0.152939
R27742 GND.n6294 GND.n6291 0.152939
R27743 GND.n6295 GND.n6294 0.152939
R27744 GND.n6296 GND.n6295 0.152939
R27745 GND.n6297 GND.n6296 0.152939
R27746 GND.n6300 GND.n6297 0.152939
R27747 GND.n6301 GND.n6300 0.152939
R27748 GND.n6302 GND.n6301 0.152939
R27749 GND.n6303 GND.n6302 0.152939
R27750 GND.n6306 GND.n6303 0.152939
R27751 GND.n6307 GND.n6306 0.152939
R27752 GND.n6308 GND.n6307 0.152939
R27753 GND.n6309 GND.n6308 0.152939
R27754 GND.n6312 GND.n6309 0.152939
R27755 GND.n6313 GND.n6312 0.152939
R27756 GND.n6314 GND.n6313 0.152939
R27757 GND.n6315 GND.n6314 0.152939
R27758 GND.n6318 GND.n6315 0.152939
R27759 GND.n6319 GND.n6318 0.152939
R27760 GND.n6320 GND.n6319 0.152939
R27761 GND.n6321 GND.n6320 0.152939
R27762 GND.n6324 GND.n6321 0.152939
R27763 GND.n6325 GND.n6324 0.152939
R27764 GND.n6326 GND.n6325 0.152939
R27765 GND.n6327 GND.n6326 0.152939
R27766 GND.n6330 GND.n6327 0.152939
R27767 GND.n6331 GND.n6330 0.152939
R27768 GND.n6332 GND.n6331 0.152939
R27769 GND.n6333 GND.n6332 0.152939
R27770 GND.n6336 GND.n6333 0.152939
R27771 GND.n6337 GND.n6336 0.152939
R27772 GND.n6338 GND.n6337 0.152939
R27773 GND.n6339 GND.n6338 0.152939
R27774 GND.n6342 GND.n6339 0.152939
R27775 GND.n6343 GND.n6342 0.152939
R27776 GND.n6344 GND.n6343 0.152939
R27777 GND.n6345 GND.n6344 0.152939
R27778 GND.n6348 GND.n6345 0.152939
R27779 GND.n6349 GND.n6348 0.152939
R27780 GND.n6350 GND.n6349 0.152939
R27781 GND.n6351 GND.n6350 0.152939
R27782 GND.n6354 GND.n6351 0.152939
R27783 GND.n6355 GND.n6354 0.152939
R27784 GND.n6356 GND.n6355 0.152939
R27785 GND.n6357 GND.n6356 0.152939
R27786 GND.n6360 GND.n6357 0.152939
R27787 GND.n6361 GND.n6360 0.152939
R27788 GND.n6362 GND.n6361 0.152939
R27789 GND.n6363 GND.n6362 0.152939
R27790 GND.n6366 GND.n6363 0.152939
R27791 GND.n6367 GND.n6366 0.152939
R27792 GND.n6368 GND.n6367 0.152939
R27793 GND.n6369 GND.n6368 0.152939
R27794 GND.n6372 GND.n6369 0.152939
R27795 GND.n6373 GND.n6372 0.152939
R27796 GND.n6374 GND.n6373 0.152939
R27797 GND.n6375 GND.n6374 0.152939
R27798 GND.n6377 GND.n6375 0.152939
R27799 GND.n6377 GND.n6376 0.152939
R27800 GND.n6376 GND.n465 0.152939
R27801 GND.n466 GND.n465 0.152939
R27802 GND.n467 GND.n466 0.152939
R27803 GND.n472 GND.n467 0.152939
R27804 GND.n473 GND.n472 0.152939
R27805 GND.n474 GND.n473 0.152939
R27806 GND.n475 GND.n474 0.152939
R27807 GND.n480 GND.n475 0.152939
R27808 GND.n481 GND.n480 0.152939
R27809 GND.n482 GND.n481 0.152939
R27810 GND.n483 GND.n482 0.152939
R27811 GND.n488 GND.n483 0.152939
R27812 GND.n489 GND.n488 0.152939
R27813 GND.n490 GND.n489 0.152939
R27814 GND.n491 GND.n490 0.152939
R27815 GND.n496 GND.n491 0.152939
R27816 GND.n497 GND.n496 0.152939
R27817 GND.n498 GND.n497 0.152939
R27818 GND.n499 GND.n498 0.152939
R27819 GND.n504 GND.n499 0.152939
R27820 GND.n505 GND.n504 0.152939
R27821 GND.n506 GND.n505 0.152939
R27822 GND.n507 GND.n506 0.152939
R27823 GND.n512 GND.n507 0.152939
R27824 GND.n513 GND.n512 0.152939
R27825 GND.n514 GND.n513 0.152939
R27826 GND.n515 GND.n514 0.152939
R27827 GND.n520 GND.n515 0.152939
R27828 GND.n521 GND.n520 0.152939
R27829 GND.n522 GND.n521 0.152939
R27830 GND.n523 GND.n522 0.152939
R27831 GND.n528 GND.n523 0.152939
R27832 GND.n529 GND.n528 0.152939
R27833 GND.n530 GND.n529 0.152939
R27834 GND.n531 GND.n530 0.152939
R27835 GND.n536 GND.n531 0.152939
R27836 GND.n537 GND.n536 0.152939
R27837 GND.n538 GND.n537 0.152939
R27838 GND.n539 GND.n538 0.152939
R27839 GND.n544 GND.n539 0.152939
R27840 GND.n545 GND.n544 0.152939
R27841 GND.n546 GND.n545 0.152939
R27842 GND.n547 GND.n546 0.152939
R27843 GND.n552 GND.n547 0.152939
R27844 GND.n553 GND.n552 0.152939
R27845 GND.n554 GND.n553 0.152939
R27846 GND.n555 GND.n554 0.152939
R27847 GND.n560 GND.n555 0.152939
R27848 GND.n561 GND.n560 0.152939
R27849 GND.n562 GND.n561 0.152939
R27850 GND.n563 GND.n562 0.152939
R27851 GND.n568 GND.n563 0.152939
R27852 GND.n569 GND.n568 0.152939
R27853 GND.n570 GND.n569 0.152939
R27854 GND.n571 GND.n570 0.152939
R27855 GND.n10530 GND.n571 0.152939
R27856 GND.n127 GND.n100 0.152939
R27857 GND.n128 GND.n127 0.152939
R27858 GND.n129 GND.n128 0.152939
R27859 GND.n147 GND.n129 0.152939
R27860 GND.n148 GND.n147 0.152939
R27861 GND.n149 GND.n148 0.152939
R27862 GND.n150 GND.n149 0.152939
R27863 GND.n168 GND.n150 0.152939
R27864 GND.n169 GND.n168 0.152939
R27865 GND.n170 GND.n169 0.152939
R27866 GND.n171 GND.n170 0.152939
R27867 GND.n189 GND.n171 0.152939
R27868 GND.n190 GND.n189 0.152939
R27869 GND.n191 GND.n190 0.152939
R27870 GND.n192 GND.n191 0.152939
R27871 GND.n210 GND.n192 0.152939
R27872 GND.n211 GND.n210 0.152939
R27873 GND.n212 GND.n211 0.152939
R27874 GND.n213 GND.n212 0.152939
R27875 GND.n231 GND.n213 0.152939
R27876 GND.n232 GND.n231 0.152939
R27877 GND.n233 GND.n232 0.152939
R27878 GND.n234 GND.n233 0.152939
R27879 GND.n252 GND.n234 0.152939
R27880 GND.n253 GND.n252 0.152939
R27881 GND.n254 GND.n253 0.152939
R27882 GND.n255 GND.n254 0.152939
R27883 GND.n272 GND.n255 0.152939
R27884 GND.n273 GND.n272 0.152939
R27885 GND.n274 GND.n273 0.152939
R27886 GND.n275 GND.n274 0.152939
R27887 GND.n293 GND.n275 0.152939
R27888 GND.n294 GND.n293 0.152939
R27889 GND.n295 GND.n294 0.152939
R27890 GND.n296 GND.n295 0.152939
R27891 GND.n314 GND.n296 0.152939
R27892 GND.n315 GND.n314 0.152939
R27893 GND.n316 GND.n315 0.152939
R27894 GND.n317 GND.n316 0.152939
R27895 GND.n335 GND.n317 0.152939
R27896 GND.n336 GND.n335 0.152939
R27897 GND.n337 GND.n336 0.152939
R27898 GND.n338 GND.n337 0.152939
R27899 GND.n356 GND.n338 0.152939
R27900 GND.n357 GND.n356 0.152939
R27901 GND.n358 GND.n357 0.152939
R27902 GND.n359 GND.n358 0.152939
R27903 GND.n377 GND.n359 0.152939
R27904 GND.n378 GND.n377 0.152939
R27905 GND.n379 GND.n378 0.152939
R27906 GND.n380 GND.n379 0.152939
R27907 GND.n398 GND.n380 0.152939
R27908 GND.n399 GND.n398 0.152939
R27909 GND.n400 GND.n399 0.152939
R27910 GND.n401 GND.n400 0.152939
R27911 GND.n419 GND.n401 0.152939
R27912 GND.n420 GND.n419 0.152939
R27913 GND.n421 GND.n420 0.152939
R27914 GND.n422 GND.n421 0.152939
R27915 GND.n440 GND.n422 0.152939
R27916 GND.n441 GND.n440 0.152939
R27917 GND.n442 GND.n441 0.152939
R27918 GND.n443 GND.n442 0.152939
R27919 GND.n5820 GND.n5814 0.152939
R27920 GND.n5821 GND.n5820 0.152939
R27921 GND.n5823 GND.n5821 0.152939
R27922 GND.n5823 GND.n5822 0.152939
R27923 GND.n5822 GND.n4830 0.152939
R27924 GND.n5027 GND.n5026 0.152939
R27925 GND.n5027 GND.n5022 0.152939
R27926 GND.n5327 GND.n5022 0.152939
R27927 GND.n5328 GND.n5327 0.152939
R27928 GND.n5329 GND.n5328 0.152939
R27929 GND.n5329 GND.n5013 0.152939
R27930 GND.n5346 GND.n5013 0.152939
R27931 GND.n5347 GND.n5346 0.152939
R27932 GND.n5348 GND.n5347 0.152939
R27933 GND.n5348 GND.n5004 0.152939
R27934 GND.n5365 GND.n5004 0.152939
R27935 GND.n5366 GND.n5365 0.152939
R27936 GND.n5367 GND.n5366 0.152939
R27937 GND.n5368 GND.n5367 0.152939
R27938 GND.n5369 GND.n5368 0.152939
R27939 GND.n5370 GND.n5369 0.152939
R27940 GND.n5371 GND.n5370 0.152939
R27941 GND.n5372 GND.n5371 0.152939
R27942 GND.n5373 GND.n5372 0.152939
R27943 GND.n5374 GND.n5373 0.152939
R27944 GND.n5375 GND.n5374 0.152939
R27945 GND.n5376 GND.n5375 0.152939
R27946 GND.n5377 GND.n5376 0.152939
R27947 GND.n5378 GND.n5377 0.152939
R27948 GND.n5379 GND.n5378 0.152939
R27949 GND.n5380 GND.n5379 0.152939
R27950 GND.n5381 GND.n5380 0.152939
R27951 GND.n5382 GND.n5381 0.152939
R27952 GND.n5384 GND.n5382 0.152939
R27953 GND.n5384 GND.n5383 0.152939
R27954 GND.n5383 GND.n4956 0.152939
R27955 GND.n5508 GND.n4956 0.152939
R27956 GND.n5509 GND.n5508 0.152939
R27957 GND.n5510 GND.n5509 0.152939
R27958 GND.n5510 GND.n4952 0.152939
R27959 GND.n5516 GND.n4952 0.152939
R27960 GND.n5517 GND.n5516 0.152939
R27961 GND.n5518 GND.n5517 0.152939
R27962 GND.n5519 GND.n5518 0.152939
R27963 GND.n5520 GND.n5519 0.152939
R27964 GND.n5521 GND.n5520 0.152939
R27965 GND.n5522 GND.n5521 0.152939
R27966 GND.n5523 GND.n5522 0.152939
R27967 GND.n5524 GND.n5523 0.152939
R27968 GND.n5525 GND.n5524 0.152939
R27969 GND.n5527 GND.n5525 0.152939
R27970 GND.n5527 GND.n5526 0.152939
R27971 GND.n5526 GND.n4925 0.152939
R27972 GND.n5611 GND.n4925 0.152939
R27973 GND.n5612 GND.n5611 0.152939
R27974 GND.n5613 GND.n5612 0.152939
R27975 GND.n5613 GND.n4921 0.152939
R27976 GND.n5619 GND.n4921 0.152939
R27977 GND.n5620 GND.n5619 0.152939
R27978 GND.n5621 GND.n5620 0.152939
R27979 GND.n5622 GND.n5621 0.152939
R27980 GND.n5623 GND.n5622 0.152939
R27981 GND.n5624 GND.n5623 0.152939
R27982 GND.n5625 GND.n5624 0.152939
R27983 GND.n5626 GND.n5625 0.152939
R27984 GND.n5627 GND.n5626 0.152939
R27985 GND.n5628 GND.n5627 0.152939
R27986 GND.n5630 GND.n5628 0.152939
R27987 GND.n5630 GND.n5629 0.152939
R27988 GND.n5629 GND.n4891 0.152939
R27989 GND.n5714 GND.n4891 0.152939
R27990 GND.n5715 GND.n5714 0.152939
R27991 GND.n5716 GND.n5715 0.152939
R27992 GND.n5716 GND.n4887 0.152939
R27993 GND.n5722 GND.n4887 0.152939
R27994 GND.n5723 GND.n5722 0.152939
R27995 GND.n5724 GND.n5723 0.152939
R27996 GND.n5725 GND.n5724 0.152939
R27997 GND.n5726 GND.n5725 0.152939
R27998 GND.n5727 GND.n5726 0.152939
R27999 GND.n5728 GND.n5727 0.152939
R28000 GND.n5729 GND.n5728 0.152939
R28001 GND.n5731 GND.n5729 0.152939
R28002 GND.n5731 GND.n5730 0.152939
R28003 GND.n5730 GND.n4851 0.152939
R28004 GND.n5805 GND.n4851 0.152939
R28005 GND.n5806 GND.n5805 0.152939
R28006 GND.n5807 GND.n5806 0.152939
R28007 GND.n5807 GND.n4849 0.152939
R28008 GND.n5813 GND.n4849 0.152939
R28009 GND.n3866 GND.n3865 0.152939
R28010 GND.n3867 GND.n3866 0.152939
R28011 GND.n3868 GND.n3867 0.152939
R28012 GND.n3869 GND.n3868 0.152939
R28013 GND.n3870 GND.n3869 0.152939
R28014 GND.n3899 GND.n3898 0.152939
R28015 GND.n3900 GND.n3899 0.152939
R28016 GND.n3901 GND.n3900 0.152939
R28017 GND.n3902 GND.n3901 0.152939
R28018 GND.n3918 GND.n3902 0.152939
R28019 GND.n3919 GND.n3918 0.152939
R28020 GND.n3920 GND.n3919 0.152939
R28021 GND.n3921 GND.n3920 0.152939
R28022 GND.n3938 GND.n3921 0.152939
R28023 GND.n3939 GND.n3938 0.152939
R28024 GND.n3940 GND.n3939 0.152939
R28025 GND.n3941 GND.n3940 0.152939
R28026 GND.n3958 GND.n3941 0.152939
R28027 GND.n3959 GND.n3958 0.152939
R28028 GND.n3960 GND.n3959 0.152939
R28029 GND.n3961 GND.n3960 0.152939
R28030 GND.n3978 GND.n3961 0.152939
R28031 GND.n3979 GND.n3978 0.152939
R28032 GND.n3980 GND.n3979 0.152939
R28033 GND.n3981 GND.n3980 0.152939
R28034 GND.n3998 GND.n3981 0.152939
R28035 GND.n3999 GND.n3998 0.152939
R28036 GND.n4000 GND.n3999 0.152939
R28037 GND.n4001 GND.n4000 0.152939
R28038 GND.n4018 GND.n4001 0.152939
R28039 GND.n4019 GND.n4018 0.152939
R28040 GND.n4020 GND.n4019 0.152939
R28041 GND.n4021 GND.n4020 0.152939
R28042 GND.n4038 GND.n4021 0.152939
R28043 GND.n4039 GND.n4038 0.152939
R28044 GND.n4040 GND.n4039 0.152939
R28045 GND.n4041 GND.n4040 0.152939
R28046 GND.n4094 GND.n4041 0.152939
R28047 GND.n4095 GND.n4094 0.152939
R28048 GND.n4096 GND.n4095 0.152939
R28049 GND.n4096 GND.n4092 0.152939
R28050 GND.n4102 GND.n4092 0.152939
R28051 GND.n4103 GND.n4102 0.152939
R28052 GND.n4104 GND.n4103 0.152939
R28053 GND.n4105 GND.n4104 0.152939
R28054 GND.n4106 GND.n4105 0.152939
R28055 GND.n4123 GND.n4106 0.152939
R28056 GND.n4124 GND.n4123 0.152939
R28057 GND.n4125 GND.n4124 0.152939
R28058 GND.n4126 GND.n4125 0.152939
R28059 GND.n4143 GND.n4126 0.152939
R28060 GND.n4144 GND.n4143 0.152939
R28061 GND.n4145 GND.n4144 0.152939
R28062 GND.n4146 GND.n4145 0.152939
R28063 GND.n4198 GND.n4146 0.152939
R28064 GND.n4199 GND.n4198 0.152939
R28065 GND.n4200 GND.n4199 0.152939
R28066 GND.n4200 GND.n4196 0.152939
R28067 GND.n4206 GND.n4196 0.152939
R28068 GND.n4207 GND.n4206 0.152939
R28069 GND.n4208 GND.n4207 0.152939
R28070 GND.n4209 GND.n4208 0.152939
R28071 GND.n4210 GND.n4209 0.152939
R28072 GND.n4227 GND.n4210 0.152939
R28073 GND.n4228 GND.n4227 0.152939
R28074 GND.n4229 GND.n4228 0.152939
R28075 GND.n4230 GND.n4229 0.152939
R28076 GND.n4245 GND.n4230 0.152939
R28077 GND.n4246 GND.n4245 0.152939
R28078 GND.n4247 GND.n4246 0.152939
R28079 GND.n4248 GND.n4247 0.152939
R28080 GND.n4301 GND.n4248 0.152939
R28081 GND.n4302 GND.n4301 0.152939
R28082 GND.n4303 GND.n4302 0.152939
R28083 GND.n4303 GND.n4299 0.152939
R28084 GND.n4309 GND.n4299 0.152939
R28085 GND.n4310 GND.n4309 0.152939
R28086 GND.n4311 GND.n4310 0.152939
R28087 GND.n4312 GND.n4311 0.152939
R28088 GND.n4313 GND.n4312 0.152939
R28089 GND.n4330 GND.n4313 0.152939
R28090 GND.n4331 GND.n4330 0.152939
R28091 GND.n4332 GND.n4331 0.152939
R28092 GND.n4333 GND.n4332 0.152939
R28093 GND.n4349 GND.n4333 0.152939
R28094 GND.n4350 GND.n4349 0.152939
R28095 GND.n4351 GND.n4350 0.152939
R28096 GND.n4352 GND.n4351 0.152939
R28097 GND.n4831 GND.n4352 0.152939
R28098 GND.n4833 GND.n4831 0.152939
R28099 GND.n6739 GND.n6738 0.152939
R28100 GND.n6748 GND.n6738 0.152939
R28101 GND.n6749 GND.n6748 0.152939
R28102 GND.n6750 GND.n6749 0.152939
R28103 GND.n6750 GND.n6734 0.152939
R28104 GND.n6763 GND.n6734 0.152939
R28105 GND.n6764 GND.n6763 0.152939
R28106 GND.n6765 GND.n6764 0.152939
R28107 GND.n6765 GND.n6528 0.152939
R28108 GND.n6778 GND.n6528 0.152939
R28109 GND.n6779 GND.n6778 0.152939
R28110 GND.n6780 GND.n6779 0.152939
R28111 GND.n6780 GND.n6524 0.152939
R28112 GND.n6793 GND.n6524 0.152939
R28113 GND.n6794 GND.n6793 0.152939
R28114 GND.n6795 GND.n6794 0.152939
R28115 GND.n6795 GND.n6520 0.152939
R28116 GND.n6808 GND.n6520 0.152939
R28117 GND.n6809 GND.n6808 0.152939
R28118 GND.n6810 GND.n6809 0.152939
R28119 GND.n6810 GND.n6516 0.152939
R28120 GND.n6823 GND.n6516 0.152939
R28121 GND.n6824 GND.n6823 0.152939
R28122 GND.n6825 GND.n6824 0.152939
R28123 GND.n6825 GND.n6511 0.152939
R28124 GND.n6838 GND.n6511 0.152939
R28125 GND.n6839 GND.n6838 0.152939
R28126 GND.n6840 GND.n6839 0.152939
R28127 GND.n6840 GND.n6507 0.152939
R28128 GND.n6853 GND.n6507 0.152939
R28129 GND.n6854 GND.n6853 0.152939
R28130 GND.n6855 GND.n6854 0.152939
R28131 GND.n6855 GND.n6503 0.152939
R28132 GND.n6868 GND.n6503 0.152939
R28133 GND.n6869 GND.n6868 0.152939
R28134 GND.n6870 GND.n6869 0.152939
R28135 GND.n6870 GND.n6499 0.152939
R28136 GND.n6883 GND.n6499 0.152939
R28137 GND.n6884 GND.n6883 0.152939
R28138 GND.n6885 GND.n6884 0.152939
R28139 GND.n6885 GND.n6495 0.152939
R28140 GND.n6898 GND.n6495 0.152939
R28141 GND.n6899 GND.n6898 0.152939
R28142 GND.n6900 GND.n6899 0.152939
R28143 GND.n6900 GND.n6491 0.152939
R28144 GND.n6913 GND.n6491 0.152939
R28145 GND.n6914 GND.n6913 0.152939
R28146 GND.n6915 GND.n6914 0.152939
R28147 GND.n6915 GND.n6486 0.152939
R28148 GND.n6928 GND.n6486 0.152939
R28149 GND.n6929 GND.n6928 0.152939
R28150 GND.n6930 GND.n6929 0.152939
R28151 GND.n6930 GND.n6482 0.152939
R28152 GND.n6943 GND.n6482 0.152939
R28153 GND.n6944 GND.n6943 0.152939
R28154 GND.n6945 GND.n6944 0.152939
R28155 GND.n6945 GND.n6478 0.152939
R28156 GND.n6958 GND.n6478 0.152939
R28157 GND.n6959 GND.n6958 0.152939
R28158 GND.n6960 GND.n6959 0.152939
R28159 GND.n6960 GND.n6474 0.152939
R28160 GND.n6973 GND.n6474 0.152939
R28161 GND.n6974 GND.n6973 0.152939
R28162 GND.n6975 GND.n6974 0.152939
R28163 GND.n6976 GND.n6975 0.152939
R28164 GND.n6977 GND.n6976 0.152939
R28165 GND.n6978 GND.n6977 0.152939
R28166 GND.n6978 GND.n86 0.152939
R28167 GND.n11114 GND.n87 0.152939
R28168 GND.n6273 GND.n87 0.152939
R28169 GND.n6274 GND.n6273 0.152939
R28170 GND.n6275 GND.n6274 0.152939
R28171 GND.n6276 GND.n6275 0.152939
R28172 GND.n6462 GND.n6276 0.152939
R28173 GND.n7020 GND.n6462 0.152939
R28174 GND.n7021 GND.n7020 0.152939
R28175 GND.n7022 GND.n7021 0.152939
R28176 GND.n7022 GND.n6458 0.152939
R28177 GND.n7035 GND.n6458 0.152939
R28178 GND.n7036 GND.n7035 0.152939
R28179 GND.n7037 GND.n7036 0.152939
R28180 GND.n7037 GND.n6454 0.152939
R28181 GND.n7050 GND.n6454 0.152939
R28182 GND.n7051 GND.n7050 0.152939
R28183 GND.n7052 GND.n7051 0.152939
R28184 GND.n7052 GND.n6450 0.152939
R28185 GND.n7065 GND.n6450 0.152939
R28186 GND.n7066 GND.n7065 0.152939
R28187 GND.n7067 GND.n7066 0.152939
R28188 GND.n7067 GND.n6446 0.152939
R28189 GND.n7080 GND.n6446 0.152939
R28190 GND.n7081 GND.n7080 0.152939
R28191 GND.n7082 GND.n7081 0.152939
R28192 GND.n7082 GND.n6442 0.152939
R28193 GND.n7095 GND.n6442 0.152939
R28194 GND.n7096 GND.n7095 0.152939
R28195 GND.n7098 GND.n7096 0.152939
R28196 GND.n7098 GND.n7097 0.152939
R28197 GND.n7097 GND.n6436 0.152939
R28198 GND.n6437 GND.n6436 0.152939
R28199 GND.n6438 GND.n6437 0.152939
R28200 GND.n7110 GND.n6438 0.152939
R28201 GND.n7111 GND.n7110 0.152939
R28202 GND.n7112 GND.n7111 0.152939
R28203 GND.n7113 GND.n7112 0.152939
R28204 GND.n7117 GND.n7113 0.152939
R28205 GND.n7118 GND.n7117 0.152939
R28206 GND.n7119 GND.n7118 0.152939
R28207 GND.n7120 GND.n7119 0.152939
R28208 GND.n7124 GND.n7120 0.152939
R28209 GND.n7125 GND.n7124 0.152939
R28210 GND.n7126 GND.n7125 0.152939
R28211 GND.n7127 GND.n7126 0.152939
R28212 GND.n7131 GND.n7127 0.152939
R28213 GND.n7132 GND.n7131 0.152939
R28214 GND.n7133 GND.n7132 0.152939
R28215 GND.n7134 GND.n7133 0.152939
R28216 GND.n7138 GND.n7134 0.152939
R28217 GND.n7139 GND.n7138 0.152939
R28218 GND.n7140 GND.n7139 0.152939
R28219 GND.n7141 GND.n7140 0.152939
R28220 GND.n7145 GND.n7141 0.152939
R28221 GND.n7146 GND.n7145 0.152939
R28222 GND.n7147 GND.n7146 0.152939
R28223 GND.n7148 GND.n7147 0.152939
R28224 GND.n7152 GND.n7148 0.152939
R28225 GND.n7153 GND.n7152 0.152939
R28226 GND.n7154 GND.n7153 0.152939
R28227 GND.n7155 GND.n7154 0.152939
R28228 GND.n7159 GND.n7155 0.152939
R28229 GND.n7160 GND.n7159 0.152939
R28230 GND.n7161 GND.n7160 0.152939
R28231 GND.n7163 GND.n7161 0.152939
R28232 GND.n7163 GND.n7162 0.152939
R28233 GND.n7162 GND.n454 0.152939
R28234 GND.n10901 GND.n454 0.152939
R28235 GND.n10684 GND.n10655 0.152939
R28236 GND.n10684 GND.n10683 0.152939
R28237 GND.n10683 GND.n10682 0.152939
R28238 GND.n10682 GND.n10656 0.152939
R28239 GND.n10657 GND.n10656 0.152939
R28240 GND.n10658 GND.n10657 0.152939
R28241 GND.n10659 GND.n10658 0.152939
R28242 GND.n10660 GND.n10659 0.152939
R28243 GND.n10661 GND.n10660 0.152939
R28244 GND.n10662 GND.n10661 0.152939
R28245 GND.n10663 GND.n10662 0.152939
R28246 GND.n10663 GND.n455 0.152939
R28247 GND.n10900 GND.n455 0.152939
R28248 GND.n10720 GND.n10719 0.152939
R28249 GND.n10721 GND.n10720 0.152939
R28250 GND.n10722 GND.n10721 0.152939
R28251 GND.n10723 GND.n10722 0.152939
R28252 GND.n10724 GND.n10723 0.152939
R28253 GND.n10725 GND.n10724 0.152939
R28254 GND.n10726 GND.n10725 0.152939
R28255 GND.n10727 GND.n10726 0.152939
R28256 GND.n10728 GND.n10727 0.152939
R28257 GND.n10729 GND.n10728 0.152939
R28258 GND.n10730 GND.n10729 0.152939
R28259 GND.n10874 GND.n10730 0.152939
R28260 GND.n10874 GND.n10873 0.152939
R28261 GND.n10873 GND.n10872 0.152939
R28262 GND.n10872 GND.n10736 0.152939
R28263 GND.n10737 GND.n10736 0.152939
R28264 GND.n10738 GND.n10737 0.152939
R28265 GND.n10739 GND.n10738 0.152939
R28266 GND.n10740 GND.n10739 0.152939
R28267 GND.n10741 GND.n10740 0.152939
R28268 GND.n10742 GND.n10741 0.152939
R28269 GND.n10743 GND.n10742 0.152939
R28270 GND.n10744 GND.n10743 0.152939
R28271 GND.n10745 GND.n10744 0.152939
R28272 GND.n10746 GND.n10745 0.152939
R28273 GND.n10747 GND.n10746 0.152939
R28274 GND.n10751 GND.n10747 0.152939
R28275 GND.n10752 GND.n10751 0.152939
R28276 GND.n10753 GND.n10752 0.152939
R28277 GND.n10754 GND.n10753 0.152939
R28278 GND.n10755 GND.n10754 0.152939
R28279 GND.n10756 GND.n10755 0.152939
R28280 GND.n10757 GND.n10756 0.152939
R28281 GND.n10758 GND.n10757 0.152939
R28282 GND.n10759 GND.n10758 0.152939
R28283 GND.n10760 GND.n10759 0.152939
R28284 GND.n10761 GND.n10760 0.152939
R28285 GND.n10762 GND.n10761 0.152939
R28286 GND.n10763 GND.n10762 0.152939
R28287 GND.n10764 GND.n10763 0.152939
R28288 GND.n10768 GND.n10764 0.152939
R28289 GND.n10769 GND.n10768 0.152939
R28290 GND.n10770 GND.n10769 0.152939
R28291 GND.n10771 GND.n10770 0.152939
R28292 GND.n10772 GND.n10771 0.152939
R28293 GND.n10773 GND.n10772 0.152939
R28294 GND.n10774 GND.n10773 0.152939
R28295 GND.n10775 GND.n10774 0.152939
R28296 GND.n10776 GND.n10775 0.152939
R28297 GND.n10777 GND.n10776 0.152939
R28298 GND.n10778 GND.n10777 0.152939
R28299 GND.n10779 GND.n10778 0.152939
R28300 GND.n10780 GND.n10779 0.152939
R28301 GND.n10781 GND.n10780 0.152939
R28302 GND.n10787 GND.n10781 0.152939
R28303 GND.n10787 GND.n10786 0.152939
R28304 GND.n4607 GND.n4606 0.152939
R28305 GND.n4608 GND.n4607 0.152939
R28306 GND.n4609 GND.n4608 0.152939
R28307 GND.n4610 GND.n4609 0.152939
R28308 GND.n4611 GND.n4610 0.152939
R28309 GND.n4612 GND.n4611 0.152939
R28310 GND.n4613 GND.n4612 0.152939
R28311 GND.n4614 GND.n4613 0.152939
R28312 GND.n4615 GND.n4614 0.152939
R28313 GND.n4616 GND.n4615 0.152939
R28314 GND.n4617 GND.n4616 0.152939
R28315 GND.n4619 GND.n4617 0.152939
R28316 GND.n4622 GND.n4619 0.152939
R28317 GND.n4623 GND.n4622 0.152939
R28318 GND.n4624 GND.n4623 0.152939
R28319 GND.n4625 GND.n4624 0.152939
R28320 GND.n4626 GND.n4625 0.152939
R28321 GND.n4627 GND.n4626 0.152939
R28322 GND.n4628 GND.n4627 0.152939
R28323 GND.n4629 GND.n4628 0.152939
R28324 GND.n4630 GND.n4629 0.152939
R28325 GND.n4631 GND.n4630 0.152939
R28326 GND.n4632 GND.n4631 0.152939
R28327 GND.n4633 GND.n4632 0.152939
R28328 GND.n4797 GND.n4796 0.152939
R28329 GND.n4798 GND.n4797 0.152939
R28330 GND.n4799 GND.n4798 0.152939
R28331 GND.n4800 GND.n4799 0.152939
R28332 GND.n4801 GND.n4800 0.152939
R28333 GND.n4802 GND.n4801 0.152939
R28334 GND.n4803 GND.n4802 0.152939
R28335 GND.n4804 GND.n4803 0.152939
R28336 GND.n4805 GND.n4804 0.152939
R28337 GND.n4806 GND.n4805 0.152939
R28338 GND.n4807 GND.n4806 0.152939
R28339 GND.n4808 GND.n4807 0.152939
R28340 GND.n4809 GND.n4808 0.152939
R28341 GND.n4813 GND.n4809 0.152939
R28342 GND.n4814 GND.n4813 0.152939
R28343 GND.n4815 GND.n4814 0.152939
R28344 GND.n4816 GND.n4815 0.152939
R28345 GND.n4817 GND.n4816 0.152939
R28346 GND.n4818 GND.n4817 0.152939
R28347 GND.n4819 GND.n4818 0.152939
R28348 GND.n4820 GND.n4819 0.152939
R28349 GND.n4821 GND.n4820 0.152939
R28350 GND.n4822 GND.n4821 0.152939
R28351 GND.n4823 GND.n4822 0.152939
R28352 GND.n4824 GND.n4823 0.152939
R28353 GND.n4825 GND.n4824 0.152939
R28354 GND.n4826 GND.n4825 0.152939
R28355 GND.n7538 GND.n4826 0.152939
R28356 GND.n7538 GND.n7537 0.152939
R28357 GND.n5924 GND.n5923 0.152939
R28358 GND.n5925 GND.n5924 0.152939
R28359 GND.n5926 GND.n5925 0.152939
R28360 GND.n5945 GND.n5926 0.152939
R28361 GND.n5946 GND.n5945 0.152939
R28362 GND.n5947 GND.n5946 0.152939
R28363 GND.n5948 GND.n5947 0.152939
R28364 GND.n5965 GND.n5948 0.152939
R28365 GND.n5966 GND.n5965 0.152939
R28366 GND.n5967 GND.n5966 0.152939
R28367 GND.n5968 GND.n5967 0.152939
R28368 GND.n5986 GND.n5968 0.152939
R28369 GND.n5987 GND.n5986 0.152939
R28370 GND.n5988 GND.n5987 0.152939
R28371 GND.n5989 GND.n5988 0.152939
R28372 GND.n6007 GND.n5989 0.152939
R28373 GND.n6008 GND.n6007 0.152939
R28374 GND.n6009 GND.n6008 0.152939
R28375 GND.n6010 GND.n6009 0.152939
R28376 GND.n6028 GND.n6010 0.152939
R28377 GND.n6029 GND.n6028 0.152939
R28378 GND.n6030 GND.n6029 0.152939
R28379 GND.n6031 GND.n6030 0.152939
R28380 GND.n6048 GND.n6031 0.152939
R28381 GND.n6049 GND.n6048 0.152939
R28382 GND.n6050 GND.n6049 0.152939
R28383 GND.n6051 GND.n6050 0.152939
R28384 GND.n6069 GND.n6051 0.152939
R28385 GND.n6070 GND.n6069 0.152939
R28386 GND.n6071 GND.n6070 0.152939
R28387 GND.n6072 GND.n6071 0.152939
R28388 GND.n6090 GND.n6072 0.152939
R28389 GND.n6091 GND.n6090 0.152939
R28390 GND.n6092 GND.n6091 0.152939
R28391 GND.n6093 GND.n6092 0.152939
R28392 GND.n6111 GND.n6093 0.152939
R28393 GND.n6112 GND.n6111 0.152939
R28394 GND.n6113 GND.n6112 0.152939
R28395 GND.n6114 GND.n6113 0.152939
R28396 GND.n6132 GND.n6114 0.152939
R28397 GND.n6133 GND.n6132 0.152939
R28398 GND.n6134 GND.n6133 0.152939
R28399 GND.n6135 GND.n6134 0.152939
R28400 GND.n6153 GND.n6135 0.152939
R28401 GND.n6154 GND.n6153 0.152939
R28402 GND.n6155 GND.n6154 0.152939
R28403 GND.n6156 GND.n6155 0.152939
R28404 GND.n6173 GND.n6156 0.152939
R28405 GND.n6174 GND.n6173 0.152939
R28406 GND.n6175 GND.n6174 0.152939
R28407 GND.n6176 GND.n6175 0.152939
R28408 GND.n6194 GND.n6176 0.152939
R28409 GND.n6195 GND.n6194 0.152939
R28410 GND.n6196 GND.n6195 0.152939
R28411 GND.n6197 GND.n6196 0.152939
R28412 GND.n6215 GND.n6197 0.152939
R28413 GND.n6216 GND.n6215 0.152939
R28414 GND.n6217 GND.n6216 0.152939
R28415 GND.n6218 GND.n6217 0.152939
R28416 GND.n6236 GND.n6218 0.152939
R28417 GND.n6237 GND.n6236 0.152939
R28418 GND.n6238 GND.n6237 0.152939
R28419 GND.n6238 GND.n101 0.152939
R28420 GND.n2538 GND.n2492 0.152939
R28421 GND.n2539 GND.n2538 0.152939
R28422 GND.n2542 GND.n2539 0.152939
R28423 GND.n2543 GND.n2542 0.152939
R28424 GND.n2544 GND.n2543 0.152939
R28425 GND.n2545 GND.n2544 0.152939
R28426 GND.n2548 GND.n2545 0.152939
R28427 GND.n2549 GND.n2548 0.152939
R28428 GND.n2550 GND.n2549 0.152939
R28429 GND.n2551 GND.n2550 0.152939
R28430 GND.n2554 GND.n2551 0.152939
R28431 GND.n2555 GND.n2554 0.152939
R28432 GND.n2556 GND.n2555 0.152939
R28433 GND.n2557 GND.n2556 0.152939
R28434 GND.n2560 GND.n2557 0.152939
R28435 GND.n2561 GND.n2560 0.152939
R28436 GND.n2562 GND.n2561 0.152939
R28437 GND.n2563 GND.n2562 0.152939
R28438 GND.n2566 GND.n2563 0.152939
R28439 GND.n2567 GND.n2566 0.152939
R28440 GND.n2568 GND.n2567 0.152939
R28441 GND.n2569 GND.n2568 0.152939
R28442 GND.n2572 GND.n2569 0.152939
R28443 GND.n2573 GND.n2572 0.152939
R28444 GND.n2574 GND.n2573 0.152939
R28445 GND.n2575 GND.n2574 0.152939
R28446 GND.n2578 GND.n2575 0.152939
R28447 GND.n2579 GND.n2578 0.152939
R28448 GND.n2580 GND.n2579 0.152939
R28449 GND.n2581 GND.n2580 0.152939
R28450 GND.n2584 GND.n2581 0.152939
R28451 GND.n2585 GND.n2584 0.152939
R28452 GND.n2586 GND.n2585 0.152939
R28453 GND.n2587 GND.n2586 0.152939
R28454 GND.n2588 GND.n2587 0.152939
R28455 GND.n2589 GND.n2588 0.152939
R28456 GND.n2589 GND.n2325 0.152939
R28457 GND.n3696 GND.n2325 0.152939
R28458 GND.n3697 GND.n3696 0.152939
R28459 GND.n3698 GND.n3697 0.152939
R28460 GND.n3699 GND.n3698 0.152939
R28461 GND.n3700 GND.n3699 0.152939
R28462 GND.n3703 GND.n3700 0.152939
R28463 GND.n3704 GND.n3703 0.152939
R28464 GND.n3705 GND.n3704 0.152939
R28465 GND.n3706 GND.n3705 0.152939
R28466 GND.n3709 GND.n3706 0.152939
R28467 GND.n3710 GND.n3709 0.152939
R28468 GND.n3711 GND.n3710 0.152939
R28469 GND.n3712 GND.n3711 0.152939
R28470 GND.n3715 GND.n3712 0.152939
R28471 GND.n3716 GND.n3715 0.152939
R28472 GND.n3717 GND.n3716 0.152939
R28473 GND.n3718 GND.n3717 0.152939
R28474 GND.n3721 GND.n3718 0.152939
R28475 GND.n3722 GND.n3721 0.152939
R28476 GND.n3723 GND.n3722 0.152939
R28477 GND.n3724 GND.n3723 0.152939
R28478 GND.n3727 GND.n3724 0.152939
R28479 GND.n3728 GND.n3727 0.152939
R28480 GND.n3729 GND.n3728 0.152939
R28481 GND.n3730 GND.n3729 0.152939
R28482 GND.n3733 GND.n3730 0.152939
R28483 GND.n3734 GND.n3733 0.152939
R28484 GND.n3735 GND.n3734 0.152939
R28485 GND.n3736 GND.n3735 0.152939
R28486 GND.n3742 GND.n3736 0.152939
R28487 GND.n3743 GND.n3742 0.152939
R28488 GND.n3744 GND.n3743 0.152939
R28489 GND.n3745 GND.n3744 0.152939
R28490 GND.n3746 GND.n3745 0.152939
R28491 GND.n3774 GND.n3746 0.152939
R28492 GND.n3775 GND.n3774 0.152939
R28493 GND.n3776 GND.n3775 0.152939
R28494 GND.n3777 GND.n3776 0.152939
R28495 GND.n3790 GND.n3777 0.152939
R28496 GND.n3791 GND.n3790 0.152939
R28497 GND.n3792 GND.n3791 0.152939
R28498 GND.n3793 GND.n3792 0.152939
R28499 GND.n3808 GND.n3793 0.152939
R28500 GND.n3809 GND.n3808 0.152939
R28501 GND.n3810 GND.n3809 0.152939
R28502 GND.n3811 GND.n3810 0.152939
R28503 GND.n3826 GND.n3811 0.152939
R28504 GND.n3827 GND.n3826 0.152939
R28505 GND.n3828 GND.n3827 0.152939
R28506 GND.n3829 GND.n3828 0.152939
R28507 GND.n3844 GND.n3829 0.152939
R28508 GND.n3845 GND.n3844 0.152939
R28509 GND.n3846 GND.n3845 0.152939
R28510 GND.n3847 GND.n3846 0.152939
R28511 GND.n3887 GND.n3847 0.152939
R28512 GND.n3888 GND.n3887 0.152939
R28513 GND.n3889 GND.n3888 0.152939
R28514 GND.n3890 GND.n3889 0.152939
R28515 GND.n3908 GND.n3890 0.152939
R28516 GND.n3909 GND.n3908 0.152939
R28517 GND.n3910 GND.n3909 0.152939
R28518 GND.n3911 GND.n3910 0.152939
R28519 GND.n3928 GND.n3911 0.152939
R28520 GND.n3929 GND.n3928 0.152939
R28521 GND.n3930 GND.n3929 0.152939
R28522 GND.n3931 GND.n3930 0.152939
R28523 GND.n3948 GND.n3931 0.152939
R28524 GND.n3949 GND.n3948 0.152939
R28525 GND.n3950 GND.n3949 0.152939
R28526 GND.n3951 GND.n3950 0.152939
R28527 GND.n3968 GND.n3951 0.152939
R28528 GND.n3969 GND.n3968 0.152939
R28529 GND.n3970 GND.n3969 0.152939
R28530 GND.n3971 GND.n3970 0.152939
R28531 GND.n3988 GND.n3971 0.152939
R28532 GND.n3989 GND.n3988 0.152939
R28533 GND.n3990 GND.n3989 0.152939
R28534 GND.n3991 GND.n3990 0.152939
R28535 GND.n4008 GND.n3991 0.152939
R28536 GND.n4009 GND.n4008 0.152939
R28537 GND.n4010 GND.n4009 0.152939
R28538 GND.n4011 GND.n4010 0.152939
R28539 GND.n4028 GND.n4011 0.152939
R28540 GND.n4029 GND.n4028 0.152939
R28541 GND.n4030 GND.n4029 0.152939
R28542 GND.n4031 GND.n4030 0.152939
R28543 GND.n4048 GND.n4031 0.152939
R28544 GND.n4049 GND.n4048 0.152939
R28545 GND.n4050 GND.n4049 0.152939
R28546 GND.n4051 GND.n4050 0.152939
R28547 GND.n4079 GND.n4051 0.152939
R28548 GND.n4080 GND.n4079 0.152939
R28549 GND.n4081 GND.n4080 0.152939
R28550 GND.n4082 GND.n4081 0.152939
R28551 GND.n4083 GND.n4082 0.152939
R28552 GND.n4113 GND.n4083 0.152939
R28553 GND.n4114 GND.n4113 0.152939
R28554 GND.n4115 GND.n4114 0.152939
R28555 GND.n4116 GND.n4115 0.152939
R28556 GND.n4133 GND.n4116 0.152939
R28557 GND.n4134 GND.n4133 0.152939
R28558 GND.n4135 GND.n4134 0.152939
R28559 GND.n4136 GND.n4135 0.152939
R28560 GND.n4153 GND.n4136 0.152939
R28561 GND.n4154 GND.n4153 0.152939
R28562 GND.n4155 GND.n4154 0.152939
R28563 GND.n4156 GND.n4155 0.152939
R28564 GND.n4184 GND.n4156 0.152939
R28565 GND.n4185 GND.n4184 0.152939
R28566 GND.n4186 GND.n4185 0.152939
R28567 GND.n4187 GND.n4186 0.152939
R28568 GND.n4188 GND.n4187 0.152939
R28569 GND.n4217 GND.n4188 0.152939
R28570 GND.n4218 GND.n4217 0.152939
R28571 GND.n4219 GND.n4218 0.152939
R28572 GND.n4220 GND.n4219 0.152939
R28573 GND.n4237 GND.n4220 0.152939
R28574 GND.n4238 GND.n4237 0.152939
R28575 GND.n4239 GND.n4238 0.152939
R28576 GND.n4240 GND.n4239 0.152939
R28577 GND.n4255 GND.n4240 0.152939
R28578 GND.n4256 GND.n4255 0.152939
R28579 GND.n4257 GND.n4256 0.152939
R28580 GND.n4258 GND.n4257 0.152939
R28581 GND.n4286 GND.n4258 0.152939
R28582 GND.n4287 GND.n4286 0.152939
R28583 GND.n4288 GND.n4287 0.152939
R28584 GND.n4289 GND.n4288 0.152939
R28585 GND.n4290 GND.n4289 0.152939
R28586 GND.n4320 GND.n4290 0.152939
R28587 GND.n4321 GND.n4320 0.152939
R28588 GND.n4322 GND.n4321 0.152939
R28589 GND.n4323 GND.n4322 0.152939
R28590 GND.n4340 GND.n4323 0.152939
R28591 GND.n4341 GND.n4340 0.152939
R28592 GND.n4342 GND.n4341 0.152939
R28593 GND.n4343 GND.n4342 0.152939
R28594 GND.n4359 GND.n4343 0.152939
R28595 GND.n4360 GND.n4359 0.152939
R28596 GND.n4361 GND.n4360 0.152939
R28597 GND.n4362 GND.n4361 0.152939
R28598 GND.n4389 GND.n4362 0.152939
R28599 GND.n4390 GND.n4389 0.152939
R28600 GND.n4391 GND.n4390 0.152939
R28601 GND.n4392 GND.n4391 0.152939
R28602 GND.n4393 GND.n4392 0.152939
R28603 GND.n4408 GND.n4393 0.152939
R28604 GND.n4409 GND.n4408 0.152939
R28605 GND.n4410 GND.n4409 0.152939
R28606 GND.n4411 GND.n4410 0.152939
R28607 GND.n4426 GND.n4411 0.152939
R28608 GND.n4427 GND.n4426 0.152939
R28609 GND.n4428 GND.n4427 0.152939
R28610 GND.n4429 GND.n4428 0.152939
R28611 GND.n4443 GND.n4429 0.152939
R28612 GND.n4444 GND.n4443 0.152939
R28613 GND.n4445 GND.n4444 0.152939
R28614 GND.n4446 GND.n4445 0.152939
R28615 GND.n4520 GND.n4446 0.152939
R28616 GND.n4521 GND.n4520 0.152939
R28617 GND.n4522 GND.n4521 0.152939
R28618 GND.n4523 GND.n4522 0.152939
R28619 GND.n4524 GND.n4523 0.152939
R28620 GND.n4562 GND.n4524 0.152939
R28621 GND.n4563 GND.n4562 0.152939
R28622 GND.n4564 GND.n4563 0.152939
R28623 GND.n4565 GND.n4564 0.152939
R28624 GND.n6542 GND.n4565 0.152939
R28625 GND.n6543 GND.n6542 0.152939
R28626 GND.n6544 GND.n6543 0.152939
R28627 GND.n6544 GND.n6538 0.152939
R28628 GND.n6550 GND.n6538 0.152939
R28629 GND.n6551 GND.n6550 0.152939
R28630 GND.n6552 GND.n6551 0.152939
R28631 GND.n6552 GND.n6534 0.152939
R28632 GND.n6558 GND.n6534 0.152939
R28633 GND.n6559 GND.n6558 0.152939
R28634 GND.n6560 GND.n6559 0.152939
R28635 GND.n6561 GND.n6560 0.152939
R28636 GND.n6562 GND.n6561 0.152939
R28637 GND.n6565 GND.n6562 0.152939
R28638 GND.n6566 GND.n6565 0.152939
R28639 GND.n6567 GND.n6566 0.152939
R28640 GND.n6568 GND.n6567 0.152939
R28641 GND.n6571 GND.n6568 0.152939
R28642 GND.n6572 GND.n6571 0.152939
R28643 GND.n6573 GND.n6572 0.152939
R28644 GND.n6574 GND.n6573 0.152939
R28645 GND.n6577 GND.n6574 0.152939
R28646 GND.n6578 GND.n6577 0.152939
R28647 GND.n6579 GND.n6578 0.152939
R28648 GND.n6580 GND.n6579 0.152939
R28649 GND.n6583 GND.n6580 0.152939
R28650 GND.n6584 GND.n6583 0.152939
R28651 GND.n6585 GND.n6584 0.152939
R28652 GND.n6586 GND.n6585 0.152939
R28653 GND.n6589 GND.n6586 0.152939
R28654 GND.n6590 GND.n6589 0.152939
R28655 GND.n6591 GND.n6590 0.152939
R28656 GND.n6592 GND.n6591 0.152939
R28657 GND.n6595 GND.n6592 0.152939
R28658 GND.n6596 GND.n6595 0.152939
R28659 GND.n6597 GND.n6596 0.152939
R28660 GND.n6598 GND.n6597 0.152939
R28661 GND.n6601 GND.n6598 0.152939
R28662 GND.n6602 GND.n6601 0.152939
R28663 GND.n6603 GND.n6602 0.152939
R28664 GND.n6604 GND.n6603 0.152939
R28665 GND.n6607 GND.n6604 0.152939
R28666 GND.n6608 GND.n6607 0.152939
R28667 GND.n6609 GND.n6608 0.152939
R28668 GND.n6610 GND.n6609 0.152939
R28669 GND.n6613 GND.n6610 0.152939
R28670 GND.n6614 GND.n6613 0.152939
R28671 GND.n6615 GND.n6614 0.152939
R28672 GND.n6616 GND.n6615 0.152939
R28673 GND.n6619 GND.n6616 0.152939
R28674 GND.n6620 GND.n6619 0.152939
R28675 GND.n6621 GND.n6620 0.152939
R28676 GND.n6622 GND.n6621 0.152939
R28677 GND.n6625 GND.n6622 0.152939
R28678 GND.n6626 GND.n6625 0.152939
R28679 GND.n6627 GND.n6626 0.152939
R28680 GND.n6628 GND.n6627 0.152939
R28681 GND.n6631 GND.n6628 0.152939
R28682 GND.n6632 GND.n6631 0.152939
R28683 GND.n6633 GND.n6632 0.152939
R28684 GND.n6634 GND.n6633 0.152939
R28685 GND.n6637 GND.n6634 0.152939
R28686 GND.n6638 GND.n6637 0.152939
R28687 GND.n6639 GND.n6638 0.152939
R28688 GND.n6640 GND.n6639 0.152939
R28689 GND.n6641 GND.n6640 0.152939
R28690 GND.n6641 GND.n102 0.152939
R28691 GND.n3496 GND.n3495 0.152939
R28692 GND.n3496 GND.n2469 0.152939
R28693 GND.n3519 GND.n2469 0.152939
R28694 GND.n3520 GND.n3519 0.152939
R28695 GND.n3521 GND.n3520 0.152939
R28696 GND.n3522 GND.n3521 0.152939
R28697 GND.n3522 GND.n2448 0.152939
R28698 GND.n3545 GND.n2448 0.152939
R28699 GND.n3546 GND.n3545 0.152939
R28700 GND.n3547 GND.n3546 0.152939
R28701 GND.n3548 GND.n3547 0.152939
R28702 GND.n3548 GND.n2426 0.152939
R28703 GND.n3571 GND.n2426 0.152939
R28704 GND.n3572 GND.n3571 0.152939
R28705 GND.n3573 GND.n3572 0.152939
R28706 GND.n3574 GND.n3573 0.152939
R28707 GND.n3574 GND.n2404 0.152939
R28708 GND.n3596 GND.n2404 0.152939
R28709 GND.n3597 GND.n3596 0.152939
R28710 GND.n3598 GND.n3597 0.152939
R28711 GND.n3599 GND.n3598 0.152939
R28712 GND.n3599 GND.n2382 0.152939
R28713 GND.n3622 GND.n2382 0.152939
R28714 GND.n3623 GND.n3622 0.152939
R28715 GND.n3624 GND.n3623 0.152939
R28716 GND.n3625 GND.n3624 0.152939
R28717 GND.n3625 GND.n2364 0.152939
R28718 GND.n3648 GND.n2364 0.152939
R28719 GND.n3649 GND.n3648 0.152939
R28720 GND.n3650 GND.n3649 0.152939
R28721 GND.n3651 GND.n3650 0.152939
R28722 GND.n3651 GND.n2342 0.152939
R28723 GND.n3674 GND.n2342 0.152939
R28724 GND.n3675 GND.n3674 0.152939
R28725 GND.n3676 GND.n3675 0.152939
R28726 GND.n3677 GND.n3676 0.152939
R28727 GND.n3677 GND.n2314 0.152939
R28728 GND.n8185 GND.n2314 0.152939
R28729 GND.n8186 GND.n8185 0.152939
R28730 GND.n8187 GND.n8186 0.152939
R28731 GND.n8188 GND.n8187 0.152939
R28732 GND.n8188 GND.n2293 0.152939
R28733 GND.n8211 GND.n2293 0.152939
R28734 GND.n8212 GND.n8211 0.152939
R28735 GND.n8213 GND.n8212 0.152939
R28736 GND.n8214 GND.n8213 0.152939
R28737 GND.n8214 GND.n2272 0.152939
R28738 GND.n8237 GND.n2272 0.152939
R28739 GND.n8238 GND.n8237 0.152939
R28740 GND.n8239 GND.n8238 0.152939
R28741 GND.n8240 GND.n8239 0.152939
R28742 GND.n8240 GND.n2250 0.152939
R28743 GND.n8263 GND.n2250 0.152939
R28744 GND.n8264 GND.n8263 0.152939
R28745 GND.n8265 GND.n8264 0.152939
R28746 GND.n8266 GND.n8265 0.152939
R28747 GND.n8266 GND.n2228 0.152939
R28748 GND.n8288 GND.n2228 0.152939
R28749 GND.n8289 GND.n8288 0.152939
R28750 GND.n8291 GND.n8289 0.152939
R28751 GND.n8291 GND.n8290 0.152939
R28752 GND.n8290 GND.n2211 0.152939
R28753 GND.n8308 GND.n2211 0.152939
R28754 GND.n1730 GND.n1729 0.152939
R28755 GND.n1731 GND.n1730 0.152939
R28756 GND.n1732 GND.n1731 0.152939
R28757 GND.n1733 GND.n1732 0.152939
R28758 GND.n1734 GND.n1733 0.152939
R28759 GND.n1735 GND.n1734 0.152939
R28760 GND.n1736 GND.n1735 0.152939
R28761 GND.n1737 GND.n1736 0.152939
R28762 GND.n1738 GND.n1737 0.152939
R28763 GND.n1739 GND.n1738 0.152939
R28764 GND.n1740 GND.n1739 0.152939
R28765 GND.n1742 GND.n1740 0.152939
R28766 GND.n1745 GND.n1742 0.152939
R28767 GND.n1746 GND.n1745 0.152939
R28768 GND.n1747 GND.n1746 0.152939
R28769 GND.n1748 GND.n1747 0.152939
R28770 GND.n1749 GND.n1748 0.152939
R28771 GND.n1750 GND.n1749 0.152939
R28772 GND.n1751 GND.n1750 0.152939
R28773 GND.n1752 GND.n1751 0.152939
R28774 GND.n1753 GND.n1752 0.152939
R28775 GND.n1754 GND.n1753 0.152939
R28776 GND.n1755 GND.n1754 0.152939
R28777 GND.n1756 GND.n1755 0.152939
R28778 GND.n1757 GND.n1756 0.152939
R28779 GND.n1758 GND.n1757 0.152939
R28780 GND.n1762 GND.n1758 0.152939
R28781 GND.n1763 GND.n1762 0.152939
R28782 GND.n1764 GND.n1763 0.152939
R28783 GND.n1765 GND.n1764 0.152939
R28784 GND.n1766 GND.n1765 0.152939
R28785 GND.n1767 GND.n1766 0.152939
R28786 GND.n1768 GND.n1767 0.152939
R28787 GND.n1769 GND.n1768 0.152939
R28788 GND.n1770 GND.n1769 0.152939
R28789 GND.n1771 GND.n1770 0.152939
R28790 GND.n1772 GND.n1771 0.152939
R28791 GND.n1773 GND.n1772 0.152939
R28792 GND.n1774 GND.n1773 0.152939
R28793 GND.n1775 GND.n1774 0.152939
R28794 GND.n1779 GND.n1775 0.152939
R28795 GND.n1780 GND.n1779 0.152939
R28796 GND.n1781 GND.n1780 0.152939
R28797 GND.n1782 GND.n1781 0.152939
R28798 GND.n1783 GND.n1782 0.152939
R28799 GND.n1784 GND.n1783 0.152939
R28800 GND.n1785 GND.n1784 0.152939
R28801 GND.n1786 GND.n1785 0.152939
R28802 GND.n1787 GND.n1786 0.152939
R28803 GND.n1788 GND.n1787 0.152939
R28804 GND.n1789 GND.n1788 0.152939
R28805 GND.n1790 GND.n1789 0.152939
R28806 GND.n1791 GND.n1790 0.152939
R28807 GND.n1792 GND.n1791 0.152939
R28808 GND.n8705 GND.n1792 0.152939
R28809 GND.n8705 GND.n8704 0.152939
R28810 GND.n1829 GND.n1825 0.152939
R28811 GND.n1830 GND.n1829 0.152939
R28812 GND.n1831 GND.n1830 0.152939
R28813 GND.n1832 GND.n1831 0.152939
R28814 GND.n1833 GND.n1832 0.152939
R28815 GND.n3154 GND.n1833 0.152939
R28816 GND.n3155 GND.n3154 0.152939
R28817 GND.n3156 GND.n3155 0.152939
R28818 GND.n3156 GND.n2894 0.152939
R28819 GND.n3178 GND.n2894 0.152939
R28820 GND.n3179 GND.n3178 0.152939
R28821 GND.n3180 GND.n3179 0.152939
R28822 GND.n3181 GND.n3180 0.152939
R28823 GND.n3181 GND.n2871 0.152939
R28824 GND.n3203 GND.n2871 0.152939
R28825 GND.n3204 GND.n3203 0.152939
R28826 GND.n3205 GND.n3204 0.152939
R28827 GND.n3206 GND.n3205 0.152939
R28828 GND.n3206 GND.n2848 0.152939
R28829 GND.n3227 GND.n2848 0.152939
R28830 GND.n3228 GND.n3227 0.152939
R28831 GND.n3229 GND.n3228 0.152939
R28832 GND.n3230 GND.n3229 0.152939
R28833 GND.n3230 GND.n2825 0.152939
R28834 GND.n3252 GND.n2825 0.152939
R28835 GND.n3253 GND.n3252 0.152939
R28836 GND.n3254 GND.n3253 0.152939
R28837 GND.n3255 GND.n3254 0.152939
R28838 GND.n3255 GND.n2803 0.152939
R28839 GND.n3277 GND.n2803 0.152939
R28840 GND.n3278 GND.n3277 0.152939
R28841 GND.n3279 GND.n3278 0.152939
R28842 GND.n3280 GND.n3279 0.152939
R28843 GND.n3280 GND.n2780 0.152939
R28844 GND.n3302 GND.n2780 0.152939
R28845 GND.n3303 GND.n3302 0.152939
R28846 GND.n3304 GND.n3303 0.152939
R28847 GND.n3305 GND.n3304 0.152939
R28848 GND.n3305 GND.n2757 0.152939
R28849 GND.n3326 GND.n2757 0.152939
R28850 GND.n3327 GND.n3326 0.152939
R28851 GND.n3328 GND.n3327 0.152939
R28852 GND.n3329 GND.n3328 0.152939
R28853 GND.n3329 GND.n2734 0.152939
R28854 GND.n3351 GND.n2734 0.152939
R28855 GND.n3352 GND.n3351 0.152939
R28856 GND.n3353 GND.n3352 0.152939
R28857 GND.n3354 GND.n3353 0.152939
R28858 GND.n3354 GND.n2712 0.152939
R28859 GND.n3376 GND.n2712 0.152939
R28860 GND.n3377 GND.n3376 0.152939
R28861 GND.n3378 GND.n3377 0.152939
R28862 GND.n3379 GND.n3378 0.152939
R28863 GND.n3379 GND.n2689 0.152939
R28864 GND.n3401 GND.n2689 0.152939
R28865 GND.n3402 GND.n3401 0.152939
R28866 GND.n3403 GND.n3402 0.152939
R28867 GND.n3404 GND.n3403 0.152939
R28868 GND.n3404 GND.n2666 0.152939
R28869 GND.n3425 GND.n2666 0.152939
R28870 GND.n3426 GND.n3425 0.152939
R28871 GND.n3427 GND.n3426 0.152939
R28872 GND.n3427 GND.n2491 0.152939
R28873 GND.n8926 GND.n1581 0.152939
R28874 GND.n8926 GND.n8925 0.152939
R28875 GND.n8925 GND.n8924 0.152939
R28876 GND.n8924 GND.n1583 0.152939
R28877 GND.n1590 GND.n1583 0.152939
R28878 GND.n1591 GND.n1590 0.152939
R28879 GND.n1592 GND.n1591 0.152939
R28880 GND.n1597 GND.n1592 0.152939
R28881 GND.n1598 GND.n1597 0.152939
R28882 GND.n1599 GND.n1598 0.152939
R28883 GND.n1600 GND.n1599 0.152939
R28884 GND.n1605 GND.n1600 0.152939
R28885 GND.n1606 GND.n1605 0.152939
R28886 GND.n1607 GND.n1606 0.152939
R28887 GND.n1608 GND.n1607 0.152939
R28888 GND.n1613 GND.n1608 0.152939
R28889 GND.n1614 GND.n1613 0.152939
R28890 GND.n1615 GND.n1614 0.152939
R28891 GND.n1616 GND.n1615 0.152939
R28892 GND.n1621 GND.n1616 0.152939
R28893 GND.n1622 GND.n1621 0.152939
R28894 GND.n1623 GND.n1622 0.152939
R28895 GND.n1624 GND.n1623 0.152939
R28896 GND.n1629 GND.n1624 0.152939
R28897 GND.n1630 GND.n1629 0.152939
R28898 GND.n1631 GND.n1630 0.152939
R28899 GND.n1632 GND.n1631 0.152939
R28900 GND.n1637 GND.n1632 0.152939
R28901 GND.n1638 GND.n1637 0.152939
R28902 GND.n1639 GND.n1638 0.152939
R28903 GND.n1640 GND.n1639 0.152939
R28904 GND.n1645 GND.n1640 0.152939
R28905 GND.n1646 GND.n1645 0.152939
R28906 GND.n1647 GND.n1646 0.152939
R28907 GND.n1648 GND.n1647 0.152939
R28908 GND.n1653 GND.n1648 0.152939
R28909 GND.n1654 GND.n1653 0.152939
R28910 GND.n1655 GND.n1654 0.152939
R28911 GND.n1656 GND.n1655 0.152939
R28912 GND.n1661 GND.n1656 0.152939
R28913 GND.n1662 GND.n1661 0.152939
R28914 GND.n1663 GND.n1662 0.152939
R28915 GND.n1664 GND.n1663 0.152939
R28916 GND.n1669 GND.n1664 0.152939
R28917 GND.n1670 GND.n1669 0.152939
R28918 GND.n1671 GND.n1670 0.152939
R28919 GND.n1672 GND.n1671 0.152939
R28920 GND.n1677 GND.n1672 0.152939
R28921 GND.n1678 GND.n1677 0.152939
R28922 GND.n1679 GND.n1678 0.152939
R28923 GND.n1680 GND.n1679 0.152939
R28924 GND.n1685 GND.n1680 0.152939
R28925 GND.n1686 GND.n1685 0.152939
R28926 GND.n1687 GND.n1686 0.152939
R28927 GND.n1688 GND.n1687 0.152939
R28928 GND.n1809 GND.n1688 0.152939
R28929 GND.n1810 GND.n1809 0.152939
R28930 GND.n1811 GND.n1810 0.152939
R28931 GND.n1812 GND.n1811 0.152939
R28932 GND.n1813 GND.n1812 0.152939
R28933 GND.n2970 GND.n1813 0.152939
R28934 GND.n2971 GND.n2970 0.152939
R28935 GND.n2976 GND.n2971 0.152939
R28936 GND.n2977 GND.n2976 0.152939
R28937 GND.n2978 GND.n2977 0.152939
R28938 GND.n2979 GND.n2978 0.152939
R28939 GND.n2980 GND.n2979 0.152939
R28940 GND.n2983 GND.n2980 0.152939
R28941 GND.n2984 GND.n2983 0.152939
R28942 GND.n2985 GND.n2984 0.152939
R28943 GND.n2986 GND.n2985 0.152939
R28944 GND.n2989 GND.n2986 0.152939
R28945 GND.n2990 GND.n2989 0.152939
R28946 GND.n2991 GND.n2990 0.152939
R28947 GND.n2992 GND.n2991 0.152939
R28948 GND.n2995 GND.n2992 0.152939
R28949 GND.n2996 GND.n2995 0.152939
R28950 GND.n2997 GND.n2996 0.152939
R28951 GND.n2998 GND.n2997 0.152939
R28952 GND.n3001 GND.n2998 0.152939
R28953 GND.n3002 GND.n3001 0.152939
R28954 GND.n3003 GND.n3002 0.152939
R28955 GND.n3004 GND.n3003 0.152939
R28956 GND.n3007 GND.n3004 0.152939
R28957 GND.n3008 GND.n3007 0.152939
R28958 GND.n3009 GND.n3008 0.152939
R28959 GND.n3010 GND.n3009 0.152939
R28960 GND.n3013 GND.n3010 0.152939
R28961 GND.n3014 GND.n3013 0.152939
R28962 GND.n3015 GND.n3014 0.152939
R28963 GND.n3016 GND.n3015 0.152939
R28964 GND.n3019 GND.n3016 0.152939
R28965 GND.n3020 GND.n3019 0.152939
R28966 GND.n3021 GND.n3020 0.152939
R28967 GND.n3022 GND.n3021 0.152939
R28968 GND.n3025 GND.n3022 0.152939
R28969 GND.n3026 GND.n3025 0.152939
R28970 GND.n3027 GND.n3026 0.152939
R28971 GND.n3028 GND.n3027 0.152939
R28972 GND.n3031 GND.n3028 0.152939
R28973 GND.n3032 GND.n3031 0.152939
R28974 GND.n3033 GND.n3032 0.152939
R28975 GND.n3034 GND.n3033 0.152939
R28976 GND.n3037 GND.n3034 0.152939
R28977 GND.n3038 GND.n3037 0.152939
R28978 GND.n3039 GND.n3038 0.152939
R28979 GND.n3040 GND.n3039 0.152939
R28980 GND.n3043 GND.n3040 0.152939
R28981 GND.n3044 GND.n3043 0.152939
R28982 GND.n3045 GND.n3044 0.152939
R28983 GND.n3046 GND.n3045 0.152939
R28984 GND.n3049 GND.n3046 0.152939
R28985 GND.n3050 GND.n3049 0.152939
R28986 GND.n3051 GND.n3050 0.152939
R28987 GND.n3052 GND.n3051 0.152939
R28988 GND.n3055 GND.n3052 0.152939
R28989 GND.n3056 GND.n3055 0.152939
R28990 GND.n3057 GND.n3056 0.152939
R28991 GND.n3058 GND.n3057 0.152939
R28992 GND.n3059 GND.n3058 0.152939
R28993 GND.n3059 GND.n2492 0.152939
R28994 GND.n9048 GND.n1463 0.152939
R28995 GND.n1468 GND.n1463 0.152939
R28996 GND.n1469 GND.n1468 0.152939
R28997 GND.n1470 GND.n1469 0.152939
R28998 GND.n1471 GND.n1470 0.152939
R28999 GND.n1476 GND.n1471 0.152939
R29000 GND.n1477 GND.n1476 0.152939
R29001 GND.n1478 GND.n1477 0.152939
R29002 GND.n1479 GND.n1478 0.152939
R29003 GND.n1484 GND.n1479 0.152939
R29004 GND.n1485 GND.n1484 0.152939
R29005 GND.n1486 GND.n1485 0.152939
R29006 GND.n1487 GND.n1486 0.152939
R29007 GND.n1492 GND.n1487 0.152939
R29008 GND.n1493 GND.n1492 0.152939
R29009 GND.n1494 GND.n1493 0.152939
R29010 GND.n1495 GND.n1494 0.152939
R29011 GND.n1500 GND.n1495 0.152939
R29012 GND.n1501 GND.n1500 0.152939
R29013 GND.n1502 GND.n1501 0.152939
R29014 GND.n1503 GND.n1502 0.152939
R29015 GND.n1508 GND.n1503 0.152939
R29016 GND.n1509 GND.n1508 0.152939
R29017 GND.n1510 GND.n1509 0.152939
R29018 GND.n1511 GND.n1510 0.152939
R29019 GND.n1516 GND.n1511 0.152939
R29020 GND.n1517 GND.n1516 0.152939
R29021 GND.n1518 GND.n1517 0.152939
R29022 GND.n1519 GND.n1518 0.152939
R29023 GND.n1524 GND.n1519 0.152939
R29024 GND.n1525 GND.n1524 0.152939
R29025 GND.n1526 GND.n1525 0.152939
R29026 GND.n1527 GND.n1526 0.152939
R29027 GND.n1532 GND.n1527 0.152939
R29028 GND.n1533 GND.n1532 0.152939
R29029 GND.n1534 GND.n1533 0.152939
R29030 GND.n1535 GND.n1534 0.152939
R29031 GND.n1540 GND.n1535 0.152939
R29032 GND.n1541 GND.n1540 0.152939
R29033 GND.n1542 GND.n1541 0.152939
R29034 GND.n1543 GND.n1542 0.152939
R29035 GND.n1548 GND.n1543 0.152939
R29036 GND.n1549 GND.n1548 0.152939
R29037 GND.n1550 GND.n1549 0.152939
R29038 GND.n1551 GND.n1550 0.152939
R29039 GND.n1556 GND.n1551 0.152939
R29040 GND.n1557 GND.n1556 0.152939
R29041 GND.n1558 GND.n1557 0.152939
R29042 GND.n1559 GND.n1558 0.152939
R29043 GND.n1564 GND.n1559 0.152939
R29044 GND.n1565 GND.n1564 0.152939
R29045 GND.n1566 GND.n1565 0.152939
R29046 GND.n1567 GND.n1566 0.152939
R29047 GND.n1572 GND.n1567 0.152939
R29048 GND.n1573 GND.n1572 0.152939
R29049 GND.n1574 GND.n1573 0.152939
R29050 GND.n1575 GND.n1574 0.152939
R29051 GND.n1580 GND.n1575 0.152939
R29052 GND.n8312 GND.n8311 0.152939
R29053 GND.n8313 GND.n8312 0.152939
R29054 GND.n8313 GND.n2207 0.152939
R29055 GND.n8319 GND.n2207 0.152939
R29056 GND.n8320 GND.n8319 0.152939
R29057 GND.n8321 GND.n8320 0.152939
R29058 GND.n8321 GND.n2203 0.152939
R29059 GND.n8327 GND.n2203 0.152939
R29060 GND.n8328 GND.n8327 0.152939
R29061 GND.n8329 GND.n8328 0.152939
R29062 GND.n8329 GND.n2199 0.152939
R29063 GND.n8337 GND.n2199 0.152939
R29064 GND.n8338 GND.n8337 0.152939
R29065 GND.n8339 GND.n8338 0.152939
R29066 GND.n8339 GND.n2195 0.152939
R29067 GND.n8345 GND.n2195 0.152939
R29068 GND.n8346 GND.n8345 0.152939
R29069 GND.n8347 GND.n8346 0.152939
R29070 GND.n8347 GND.n2191 0.152939
R29071 GND.n8353 GND.n2191 0.152939
R29072 GND.n8354 GND.n8353 0.152939
R29073 GND.n8355 GND.n8354 0.152939
R29074 GND.n8355 GND.n2187 0.152939
R29075 GND.n8361 GND.n2187 0.152939
R29076 GND.n8453 GND.n8452 0.152939
R29077 GND.n8452 GND.n8451 0.152939
R29078 GND.n8451 GND.n8363 0.152939
R29079 GND.n8447 GND.n8363 0.152939
R29080 GND.n8447 GND.n8446 0.152939
R29081 GND.n8446 GND.n8445 0.152939
R29082 GND.n8445 GND.n8369 0.152939
R29083 GND.n8441 GND.n8369 0.152939
R29084 GND.n8441 GND.n8440 0.152939
R29085 GND.n8440 GND.n8439 0.152939
R29086 GND.n8439 GND.n8375 0.152939
R29087 GND.n8435 GND.n8375 0.152939
R29088 GND.n8435 GND.n8434 0.152939
R29089 GND.n8434 GND.n8433 0.152939
R29090 GND.n8433 GND.n8381 0.152939
R29091 GND.n8429 GND.n8381 0.152939
R29092 GND.n8429 GND.n8428 0.152939
R29093 GND.n8428 GND.n8427 0.152939
R29094 GND.n8427 GND.n8390 0.152939
R29095 GND.n8423 GND.n8390 0.152939
R29096 GND.n8423 GND.n8422 0.152939
R29097 GND.n8422 GND.n8421 0.152939
R29098 GND.n8421 GND.n8396 0.152939
R29099 GND.n8417 GND.n8396 0.152939
R29100 GND.n8417 GND.n8416 0.152939
R29101 GND.n8416 GND.n8415 0.152939
R29102 GND.n8415 GND.n8402 0.152939
R29103 GND.n8408 GND.n8402 0.152939
R29104 GND.n8410 GND.n8408 0.152939
R29105 GND.n8702 GND.n1797 0.152939
R29106 GND.n2924 GND.n1797 0.152939
R29107 GND.n2925 GND.n2924 0.152939
R29108 GND.n2925 GND.n2920 0.152939
R29109 GND.n2933 GND.n2920 0.152939
R29110 GND.n2934 GND.n2933 0.152939
R29111 GND.n2935 GND.n2934 0.152939
R29112 GND.n2935 GND.n2918 0.152939
R29113 GND.n2943 GND.n2918 0.152939
R29114 GND.n2944 GND.n2943 0.152939
R29115 GND.n2945 GND.n2944 0.152939
R29116 GND.n2945 GND.n2912 0.152939
R29117 GND.n2950 GND.n2912 0.152939
R29118 GND.n2952 GND.n2951 0.152939
R29119 GND.n2952 GND.n2910 0.152939
R29120 GND.n2958 GND.n2910 0.152939
R29121 GND.n2959 GND.n2958 0.152939
R29122 GND.n2960 GND.n2959 0.152939
R29123 GND.n2960 GND.n2905 0.152939
R29124 GND.n3163 GND.n2905 0.152939
R29125 GND.n3164 GND.n3163 0.152939
R29126 GND.n3166 GND.n3164 0.152939
R29127 GND.n3166 GND.n3165 0.152939
R29128 GND.n3165 GND.n2883 0.152939
R29129 GND.n3188 GND.n2883 0.152939
R29130 GND.n3189 GND.n3188 0.152939
R29131 GND.n3191 GND.n3189 0.152939
R29132 GND.n3191 GND.n3190 0.152939
R29133 GND.n3190 GND.n2861 0.152939
R29134 GND.n3213 GND.n2861 0.152939
R29135 GND.n3214 GND.n3213 0.152939
R29136 GND.n3216 GND.n3214 0.152939
R29137 GND.n3216 GND.n3215 0.152939
R29138 GND.n3215 GND.n2837 0.152939
R29139 GND.n3237 GND.n2837 0.152939
R29140 GND.n3238 GND.n3237 0.152939
R29141 GND.n3240 GND.n3238 0.152939
R29142 GND.n3240 GND.n3239 0.152939
R29143 GND.n3239 GND.n2814 0.152939
R29144 GND.n3262 GND.n2814 0.152939
R29145 GND.n3263 GND.n3262 0.152939
R29146 GND.n3265 GND.n3263 0.152939
R29147 GND.n3265 GND.n3264 0.152939
R29148 GND.n3264 GND.n2792 0.152939
R29149 GND.n3287 GND.n2792 0.152939
R29150 GND.n3288 GND.n3287 0.152939
R29151 GND.n3290 GND.n3288 0.152939
R29152 GND.n3290 GND.n3289 0.152939
R29153 GND.n3289 GND.n2770 0.152939
R29154 GND.n3312 GND.n2770 0.152939
R29155 GND.n3313 GND.n3312 0.152939
R29156 GND.n3315 GND.n3313 0.152939
R29157 GND.n3315 GND.n3314 0.152939
R29158 GND.n3314 GND.n2746 0.152939
R29159 GND.n3336 GND.n2746 0.152939
R29160 GND.n3337 GND.n3336 0.152939
R29161 GND.n3339 GND.n3337 0.152939
R29162 GND.n3339 GND.n3338 0.152939
R29163 GND.n3338 GND.n2723 0.152939
R29164 GND.n3361 GND.n2723 0.152939
R29165 GND.n3362 GND.n3361 0.152939
R29166 GND.n3364 GND.n3362 0.152939
R29167 GND.n3364 GND.n3363 0.152939
R29168 GND.n3363 GND.n2701 0.152939
R29169 GND.n3386 GND.n2701 0.152939
R29170 GND.n3387 GND.n3386 0.152939
R29171 GND.n3389 GND.n3387 0.152939
R29172 GND.n3389 GND.n3388 0.152939
R29173 GND.n3388 GND.n2679 0.152939
R29174 GND.n3411 GND.n2679 0.152939
R29175 GND.n3412 GND.n3411 0.152939
R29176 GND.n3414 GND.n3412 0.152939
R29177 GND.n3414 GND.n3413 0.152939
R29178 GND.n3413 GND.n2657 0.152939
R29179 GND.n3433 GND.n2657 0.152939
R29180 GND.n3434 GND.n3433 0.152939
R29181 GND.n3435 GND.n3434 0.152939
R29182 GND.n3435 GND.n2655 0.152939
R29183 GND.n3441 GND.n2655 0.152939
R29184 GND.n3442 GND.n3441 0.152939
R29185 GND.n3444 GND.n3442 0.152939
R29186 GND.n8043 GND.n3874 0.131598
R29187 GND.n5872 GND.n4834 0.131598
R29188 GND.n11107 GND.n100 0.0767195
R29189 GND.n5872 GND.n4830 0.0767195
R29190 GND.n8043 GND.n3870 0.0767195
R29191 GND.n11107 GND.n101 0.0767195
R29192 GND.n3495 GND.n3494 0.0767195
R29193 GND.n3494 GND.n2491 0.0767195
R29194 GND.n3443 GND.n2653 0.0695946
R29195 GND.n11115 GND.n86 0.0695946
R29196 GND.n11115 GND.n11114 0.0695946
R29197 GND.n3444 GND.n3443 0.0695946
R29198 GND.n7536 GND.n5873 0.063
R29199 GND.n2131 GND.n2122 0.063
R29200 GND.n7536 GND.n7535 0.0460163
R29201 GND.n10909 GND.n451 0.0460163
R29202 GND.n8703 GND.n1796 0.0460163
R29203 GND.n8483 GND.n2122 0.0460163
R29204 GND.n7535 GND.n5875 0.0344674
R29205 GND.n6742 GND.n5875 0.0344674
R29206 GND.n6742 GND.n5935 0.0344674
R29207 GND.n5936 GND.n5935 0.0344674
R29208 GND.n5937 GND.n5936 0.0344674
R29209 GND.n6757 GND.n5937 0.0344674
R29210 GND.n6757 GND.n5955 0.0344674
R29211 GND.n5956 GND.n5955 0.0344674
R29212 GND.n5957 GND.n5956 0.0344674
R29213 GND.n6772 GND.n5957 0.0344674
R29214 GND.n6772 GND.n5976 0.0344674
R29215 GND.n5977 GND.n5976 0.0344674
R29216 GND.n5978 GND.n5977 0.0344674
R29217 GND.n6787 GND.n5978 0.0344674
R29218 GND.n6787 GND.n5997 0.0344674
R29219 GND.n5998 GND.n5997 0.0344674
R29220 GND.n5999 GND.n5998 0.0344674
R29221 GND.n6802 GND.n5999 0.0344674
R29222 GND.n6802 GND.n6018 0.0344674
R29223 GND.n6019 GND.n6018 0.0344674
R29224 GND.n6020 GND.n6019 0.0344674
R29225 GND.n6817 GND.n6020 0.0344674
R29226 GND.n6817 GND.n6038 0.0344674
R29227 GND.n6039 GND.n6038 0.0344674
R29228 GND.n6040 GND.n6039 0.0344674
R29229 GND.n6832 GND.n6040 0.0344674
R29230 GND.n6832 GND.n6059 0.0344674
R29231 GND.n6060 GND.n6059 0.0344674
R29232 GND.n6061 GND.n6060 0.0344674
R29233 GND.n6847 GND.n6061 0.0344674
R29234 GND.n6847 GND.n6080 0.0344674
R29235 GND.n6081 GND.n6080 0.0344674
R29236 GND.n6082 GND.n6081 0.0344674
R29237 GND.n6862 GND.n6082 0.0344674
R29238 GND.n6862 GND.n6101 0.0344674
R29239 GND.n6102 GND.n6101 0.0344674
R29240 GND.n6103 GND.n6102 0.0344674
R29241 GND.n6877 GND.n6103 0.0344674
R29242 GND.n6877 GND.n6122 0.0344674
R29243 GND.n6123 GND.n6122 0.0344674
R29244 GND.n6124 GND.n6123 0.0344674
R29245 GND.n6892 GND.n6124 0.0344674
R29246 GND.n6892 GND.n6143 0.0344674
R29247 GND.n6144 GND.n6143 0.0344674
R29248 GND.n6145 GND.n6144 0.0344674
R29249 GND.n6907 GND.n6145 0.0344674
R29250 GND.n6907 GND.n6164 0.0344674
R29251 GND.n6165 GND.n6164 0.0344674
R29252 GND.n6166 GND.n6165 0.0344674
R29253 GND.n6922 GND.n6166 0.0344674
R29254 GND.n6922 GND.n6184 0.0344674
R29255 GND.n6185 GND.n6184 0.0344674
R29256 GND.n6186 GND.n6185 0.0344674
R29257 GND.n6937 GND.n6186 0.0344674
R29258 GND.n6937 GND.n6205 0.0344674
R29259 GND.n6206 GND.n6205 0.0344674
R29260 GND.n6207 GND.n6206 0.0344674
R29261 GND.n6952 GND.n6207 0.0344674
R29262 GND.n6952 GND.n6226 0.0344674
R29263 GND.n6227 GND.n6226 0.0344674
R29264 GND.n6228 GND.n6227 0.0344674
R29265 GND.n6967 GND.n6228 0.0344674
R29266 GND.n6967 GND.n6246 0.0344674
R29267 GND.n6247 GND.n6246 0.0344674
R29268 GND.n6248 GND.n6247 0.0344674
R29269 GND.n6990 GND.n6248 0.0344674
R29270 GND.n6991 GND.n6990 0.0344674
R29271 GND.n6991 GND.n6468 0.0344674
R29272 GND.n6999 GND.n6468 0.0344674
R29273 GND.n6999 GND.n6464 0.0344674
R29274 GND.n7008 GND.n6464 0.0344674
R29275 GND.n7009 GND.n7008 0.0344674
R29276 GND.n7009 GND.n118 0.0344674
R29277 GND.n119 GND.n118 0.0344674
R29278 GND.n120 GND.n119 0.0344674
R29279 GND.n7014 GND.n120 0.0344674
R29280 GND.n7014 GND.n137 0.0344674
R29281 GND.n138 GND.n137 0.0344674
R29282 GND.n139 GND.n138 0.0344674
R29283 GND.n7029 GND.n139 0.0344674
R29284 GND.n7029 GND.n158 0.0344674
R29285 GND.n159 GND.n158 0.0344674
R29286 GND.n160 GND.n159 0.0344674
R29287 GND.n7044 GND.n160 0.0344674
R29288 GND.n7044 GND.n179 0.0344674
R29289 GND.n180 GND.n179 0.0344674
R29290 GND.n181 GND.n180 0.0344674
R29291 GND.n7059 GND.n181 0.0344674
R29292 GND.n7059 GND.n200 0.0344674
R29293 GND.n201 GND.n200 0.0344674
R29294 GND.n202 GND.n201 0.0344674
R29295 GND.n7074 GND.n202 0.0344674
R29296 GND.n7074 GND.n221 0.0344674
R29297 GND.n222 GND.n221 0.0344674
R29298 GND.n223 GND.n222 0.0344674
R29299 GND.n7089 GND.n223 0.0344674
R29300 GND.n7089 GND.n242 0.0344674
R29301 GND.n243 GND.n242 0.0344674
R29302 GND.n244 GND.n243 0.0344674
R29303 GND.n7105 GND.n244 0.0344674
R29304 GND.n7105 GND.n262 0.0344674
R29305 GND.n263 GND.n262 0.0344674
R29306 GND.n264 GND.n263 0.0344674
R29307 GND.n7108 GND.n264 0.0344674
R29308 GND.n7108 GND.n283 0.0344674
R29309 GND.n284 GND.n283 0.0344674
R29310 GND.n285 GND.n284 0.0344674
R29311 GND.n7115 GND.n285 0.0344674
R29312 GND.n7115 GND.n304 0.0344674
R29313 GND.n305 GND.n304 0.0344674
R29314 GND.n306 GND.n305 0.0344674
R29315 GND.n7122 GND.n306 0.0344674
R29316 GND.n7122 GND.n325 0.0344674
R29317 GND.n326 GND.n325 0.0344674
R29318 GND.n327 GND.n326 0.0344674
R29319 GND.n7129 GND.n327 0.0344674
R29320 GND.n7129 GND.n346 0.0344674
R29321 GND.n347 GND.n346 0.0344674
R29322 GND.n348 GND.n347 0.0344674
R29323 GND.n7136 GND.n348 0.0344674
R29324 GND.n7136 GND.n367 0.0344674
R29325 GND.n368 GND.n367 0.0344674
R29326 GND.n369 GND.n368 0.0344674
R29327 GND.n7143 GND.n369 0.0344674
R29328 GND.n7143 GND.n388 0.0344674
R29329 GND.n389 GND.n388 0.0344674
R29330 GND.n390 GND.n389 0.0344674
R29331 GND.n7150 GND.n390 0.0344674
R29332 GND.n7150 GND.n409 0.0344674
R29333 GND.n410 GND.n409 0.0344674
R29334 GND.n411 GND.n410 0.0344674
R29335 GND.n7157 GND.n411 0.0344674
R29336 GND.n7157 GND.n430 0.0344674
R29337 GND.n431 GND.n430 0.0344674
R29338 GND.n432 GND.n431 0.0344674
R29339 GND.n450 GND.n432 0.0344674
R29340 GND.n10909 GND.n450 0.0344674
R29341 GND.n1852 GND.n1796 0.0344674
R29342 GND.n1852 GND.n1847 0.0344674
R29343 GND.n1857 GND.n1847 0.0344674
R29344 GND.n1857 GND.n1844 0.0344674
R29345 GND.n8681 GND.n1844 0.0344674
R29346 GND.n8681 GND.n1845 0.0344674
R29347 GND.n8677 GND.n1845 0.0344674
R29348 GND.n8677 GND.n8676 0.0344674
R29349 GND.n8676 GND.n8675 0.0344674
R29350 GND.n8675 GND.n1866 0.0344674
R29351 GND.n8671 GND.n1866 0.0344674
R29352 GND.n8671 GND.n8670 0.0344674
R29353 GND.n8670 GND.n8669 0.0344674
R29354 GND.n8669 GND.n1874 0.0344674
R29355 GND.n8665 GND.n1874 0.0344674
R29356 GND.n8665 GND.n8664 0.0344674
R29357 GND.n8664 GND.n8663 0.0344674
R29358 GND.n8663 GND.n1882 0.0344674
R29359 GND.n8659 GND.n1882 0.0344674
R29360 GND.n8659 GND.n8658 0.0344674
R29361 GND.n8658 GND.n8657 0.0344674
R29362 GND.n8657 GND.n1890 0.0344674
R29363 GND.n8653 GND.n1890 0.0344674
R29364 GND.n8653 GND.n8652 0.0344674
R29365 GND.n8652 GND.n8651 0.0344674
R29366 GND.n8651 GND.n1898 0.0344674
R29367 GND.n8647 GND.n1898 0.0344674
R29368 GND.n8647 GND.n8646 0.0344674
R29369 GND.n8646 GND.n8645 0.0344674
R29370 GND.n8645 GND.n1906 0.0344674
R29371 GND.n8641 GND.n1906 0.0344674
R29372 GND.n8641 GND.n8640 0.0344674
R29373 GND.n8640 GND.n8639 0.0344674
R29374 GND.n8639 GND.n1914 0.0344674
R29375 GND.n8635 GND.n1914 0.0344674
R29376 GND.n8635 GND.n8634 0.0344674
R29377 GND.n8634 GND.n8633 0.0344674
R29378 GND.n8633 GND.n1922 0.0344674
R29379 GND.n8629 GND.n1922 0.0344674
R29380 GND.n8629 GND.n8628 0.0344674
R29381 GND.n8628 GND.n8627 0.0344674
R29382 GND.n8627 GND.n1930 0.0344674
R29383 GND.n8623 GND.n1930 0.0344674
R29384 GND.n8623 GND.n8622 0.0344674
R29385 GND.n8622 GND.n8621 0.0344674
R29386 GND.n8621 GND.n1938 0.0344674
R29387 GND.n8617 GND.n1938 0.0344674
R29388 GND.n8617 GND.n8616 0.0344674
R29389 GND.n8616 GND.n8615 0.0344674
R29390 GND.n8615 GND.n1946 0.0344674
R29391 GND.n8611 GND.n1946 0.0344674
R29392 GND.n8611 GND.n8610 0.0344674
R29393 GND.n8610 GND.n8609 0.0344674
R29394 GND.n8609 GND.n1954 0.0344674
R29395 GND.n8605 GND.n1954 0.0344674
R29396 GND.n8605 GND.n8604 0.0344674
R29397 GND.n8604 GND.n8603 0.0344674
R29398 GND.n8603 GND.n1962 0.0344674
R29399 GND.n8599 GND.n1962 0.0344674
R29400 GND.n8599 GND.n8598 0.0344674
R29401 GND.n8598 GND.n8597 0.0344674
R29402 GND.n8597 GND.n1970 0.0344674
R29403 GND.n8593 GND.n1970 0.0344674
R29404 GND.n8593 GND.n8592 0.0344674
R29405 GND.n8592 GND.n8591 0.0344674
R29406 GND.n8591 GND.n1978 0.0344674
R29407 GND.n8587 GND.n1978 0.0344674
R29408 GND.n8587 GND.n8586 0.0344674
R29409 GND.n8586 GND.n8585 0.0344674
R29410 GND.n8585 GND.n1986 0.0344674
R29411 GND.n8581 GND.n1986 0.0344674
R29412 GND.n8581 GND.n8580 0.0344674
R29413 GND.n8580 GND.n8579 0.0344674
R29414 GND.n8579 GND.n1994 0.0344674
R29415 GND.n8575 GND.n1994 0.0344674
R29416 GND.n8575 GND.n8574 0.0344674
R29417 GND.n8574 GND.n8573 0.0344674
R29418 GND.n8573 GND.n2002 0.0344674
R29419 GND.n8569 GND.n2002 0.0344674
R29420 GND.n8569 GND.n8568 0.0344674
R29421 GND.n8568 GND.n8567 0.0344674
R29422 GND.n8567 GND.n2010 0.0344674
R29423 GND.n8563 GND.n2010 0.0344674
R29424 GND.n8563 GND.n8562 0.0344674
R29425 GND.n8562 GND.n8561 0.0344674
R29426 GND.n8561 GND.n2018 0.0344674
R29427 GND.n8557 GND.n2018 0.0344674
R29428 GND.n8557 GND.n8556 0.0344674
R29429 GND.n8556 GND.n8555 0.0344674
R29430 GND.n8555 GND.n2026 0.0344674
R29431 GND.n8551 GND.n2026 0.0344674
R29432 GND.n8551 GND.n8550 0.0344674
R29433 GND.n8550 GND.n8549 0.0344674
R29434 GND.n8549 GND.n2034 0.0344674
R29435 GND.n8545 GND.n2034 0.0344674
R29436 GND.n8545 GND.n8544 0.0344674
R29437 GND.n8544 GND.n8543 0.0344674
R29438 GND.n8543 GND.n2042 0.0344674
R29439 GND.n8539 GND.n2042 0.0344674
R29440 GND.n8539 GND.n8538 0.0344674
R29441 GND.n8538 GND.n8537 0.0344674
R29442 GND.n8537 GND.n2050 0.0344674
R29443 GND.n8533 GND.n2050 0.0344674
R29444 GND.n8533 GND.n8532 0.0344674
R29445 GND.n8532 GND.n8531 0.0344674
R29446 GND.n8531 GND.n2058 0.0344674
R29447 GND.n8527 GND.n2058 0.0344674
R29448 GND.n8527 GND.n8526 0.0344674
R29449 GND.n8526 GND.n8525 0.0344674
R29450 GND.n8525 GND.n2066 0.0344674
R29451 GND.n8521 GND.n2066 0.0344674
R29452 GND.n8521 GND.n8520 0.0344674
R29453 GND.n8520 GND.n8519 0.0344674
R29454 GND.n8519 GND.n2074 0.0344674
R29455 GND.n8515 GND.n2074 0.0344674
R29456 GND.n8515 GND.n8514 0.0344674
R29457 GND.n8514 GND.n8513 0.0344674
R29458 GND.n8513 GND.n2082 0.0344674
R29459 GND.n8509 GND.n2082 0.0344674
R29460 GND.n8509 GND.n8508 0.0344674
R29461 GND.n8508 GND.n8507 0.0344674
R29462 GND.n8507 GND.n2090 0.0344674
R29463 GND.n8503 GND.n2090 0.0344674
R29464 GND.n8503 GND.n8502 0.0344674
R29465 GND.n8502 GND.n8501 0.0344674
R29466 GND.n8501 GND.n2098 0.0344674
R29467 GND.n8497 GND.n2098 0.0344674
R29468 GND.n8497 GND.n8496 0.0344674
R29469 GND.n8496 GND.n8495 0.0344674
R29470 GND.n8495 GND.n2106 0.0344674
R29471 GND.n8491 GND.n2106 0.0344674
R29472 GND.n8491 GND.n8490 0.0344674
R29473 GND.n8490 GND.n8489 0.0344674
R29474 GND.n8489 GND.n2114 0.0344674
R29475 GND.n8485 GND.n2114 0.0344674
R29476 GND.n8485 GND.n8484 0.0344674
R29477 GND.n8484 GND.n8483 0.0344674
R29478 VP.n148 VP.t1 243.97
R29479 VP.n149 VP.t0 243.255
R29480 VP.n148 VP.n147 223.454
R29481 VP.n95 VP.n94 161.3
R29482 VP.n96 VP.n91 161.3
R29483 VP.n98 VP.n97 161.3
R29484 VP.n99 VP.n90 161.3
R29485 VP.n101 VP.n100 161.3
R29486 VP.n102 VP.n89 161.3
R29487 VP.n104 VP.n103 161.3
R29488 VP.n105 VP.n88 161.3
R29489 VP.n108 VP.n107 161.3
R29490 VP.n109 VP.n87 161.3
R29491 VP.n111 VP.n110 161.3
R29492 VP.n112 VP.n86 161.3
R29493 VP.n114 VP.n113 161.3
R29494 VP.n115 VP.n85 161.3
R29495 VP.n117 VP.n116 161.3
R29496 VP.n118 VP.n83 161.3
R29497 VP.n120 VP.n119 161.3
R29498 VP.n121 VP.n82 161.3
R29499 VP.n123 VP.n122 161.3
R29500 VP.n124 VP.n81 161.3
R29501 VP.n126 VP.n125 161.3
R29502 VP.n127 VP.n80 161.3
R29503 VP.n129 VP.n128 161.3
R29504 VP.n130 VP.n78 161.3
R29505 VP.n132 VP.n131 161.3
R29506 VP.n133 VP.n77 161.3
R29507 VP.n135 VP.n134 161.3
R29508 VP.n136 VP.n76 161.3
R29509 VP.n138 VP.n137 161.3
R29510 VP.n139 VP.n75 161.3
R29511 VP.n141 VP.n140 161.3
R29512 VP.n142 VP.n74 161.3
R29513 VP.n144 VP.n143 161.3
R29514 VP.n71 VP.n70 161.3
R29515 VP.n69 VP.n1 161.3
R29516 VP.n68 VP.n67 161.3
R29517 VP.n66 VP.n2 161.3
R29518 VP.n65 VP.n64 161.3
R29519 VP.n63 VP.n3 161.3
R29520 VP.n62 VP.n61 161.3
R29521 VP.n60 VP.n4 161.3
R29522 VP.n59 VP.n58 161.3
R29523 VP.n56 VP.n5 161.3
R29524 VP.n55 VP.n54 161.3
R29525 VP.n53 VP.n6 161.3
R29526 VP.n52 VP.n51 161.3
R29527 VP.n50 VP.n7 161.3
R29528 VP.n49 VP.n48 161.3
R29529 VP.n47 VP.n8 161.3
R29530 VP.n46 VP.n45 161.3
R29531 VP.n43 VP.n9 161.3
R29532 VP.n42 VP.n41 161.3
R29533 VP.n40 VP.n10 161.3
R29534 VP.n39 VP.n38 161.3
R29535 VP.n37 VP.n11 161.3
R29536 VP.n36 VP.n35 161.3
R29537 VP.n34 VP.n12 161.3
R29538 VP.n33 VP.n32 161.3
R29539 VP.n30 VP.n13 161.3
R29540 VP.n29 VP.n28 161.3
R29541 VP.n27 VP.n14 161.3
R29542 VP.n26 VP.n25 161.3
R29543 VP.n24 VP.n15 161.3
R29544 VP.n23 VP.n22 161.3
R29545 VP.n21 VP.n16 161.3
R29546 VP.n20 VP.n19 161.3
R29547 VP.n145 VP.n73 77.9496
R29548 VP.n72 VP.n0 77.9496
R29549 VP.n17 VP.t9 76.2399
R29550 VP.n92 VP.t5 76.2397
R29551 VP.n137 VP.n75 73.0308
R29552 VP.n64 VP.n2 73.0308
R29553 VP.n93 VP.n92 69.3319
R29554 VP.n18 VP.n17 69.3319
R29555 VP.n125 VP.n80 66.2494
R29556 VP.n100 VP.n99 66.2494
R29557 VP.n25 VP.n24 66.2494
R29558 VP.n51 VP.n6 66.2494
R29559 VP.n113 VP.n85 56.5617
R29560 VP.n113 VP.n112 56.5617
R29561 VP.n38 VP.n37 56.5617
R29562 VP.n38 VP.n10 56.5617
R29563 VP.n146 VP.n145 46.9281
R29564 VP.n125 VP.n124 46.874
R29565 VP.n100 VP.n89 46.874
R29566 VP.n25 VP.n14 46.874
R29567 VP.n51 VP.n50 46.874
R29568 VP.n73 VP.t6 41.7552
R29569 VP.n79 VP.t12 41.7552
R29570 VP.n84 VP.t15 41.7552
R29571 VP.n106 VP.t4 41.7552
R29572 VP.n93 VP.t10 41.7552
R29573 VP.n18 VP.t14 41.7552
R29574 VP.n31 VP.t11 41.7552
R29575 VP.n44 VP.t8 41.7552
R29576 VP.n57 VP.t7 41.7552
R29577 VP.n0 VP.t13 41.7552
R29578 VP.n137 VP.n136 37.1863
R29579 VP.n64 VP.n63 37.1863
R29580 VP.n141 VP.n75 27.4986
R29581 VP.n68 VP.n2 27.4986
R29582 VP.n143 VP.n142 24.5923
R29583 VP.n142 VP.n141 24.5923
R29584 VP.n136 VP.n135 24.5923
R29585 VP.n135 VP.n77 24.5923
R29586 VP.n131 VP.n130 24.5923
R29587 VP.n130 VP.n129 24.5923
R29588 VP.n129 VP.n80 24.5923
R29589 VP.n124 VP.n123 24.5923
R29590 VP.n123 VP.n82 24.5923
R29591 VP.n119 VP.n118 24.5923
R29592 VP.n118 VP.n117 24.5923
R29593 VP.n117 VP.n85 24.5923
R29594 VP.n112 VP.n111 24.5923
R29595 VP.n111 VP.n87 24.5923
R29596 VP.n107 VP.n87 24.5923
R29597 VP.n105 VP.n104 24.5923
R29598 VP.n104 VP.n89 24.5923
R29599 VP.n99 VP.n98 24.5923
R29600 VP.n98 VP.n91 24.5923
R29601 VP.n94 VP.n91 24.5923
R29602 VP.n19 VP.n16 24.5923
R29603 VP.n23 VP.n16 24.5923
R29604 VP.n24 VP.n23 24.5923
R29605 VP.n29 VP.n14 24.5923
R29606 VP.n30 VP.n29 24.5923
R29607 VP.n32 VP.n12 24.5923
R29608 VP.n36 VP.n12 24.5923
R29609 VP.n37 VP.n36 24.5923
R29610 VP.n42 VP.n10 24.5923
R29611 VP.n43 VP.n42 24.5923
R29612 VP.n45 VP.n43 24.5923
R29613 VP.n49 VP.n8 24.5923
R29614 VP.n50 VP.n49 24.5923
R29615 VP.n55 VP.n6 24.5923
R29616 VP.n56 VP.n55 24.5923
R29617 VP.n58 VP.n56 24.5923
R29618 VP.n62 VP.n4 24.5923
R29619 VP.n63 VP.n62 24.5923
R29620 VP.n69 VP.n68 24.5923
R29621 VP.n70 VP.n69 24.5923
R29622 VP.n84 VP.n82 22.1332
R29623 VP.n106 VP.n105 22.1332
R29624 VP.n31 VP.n30 22.1332
R29625 VP.n44 VP.n8 22.1332
R29626 VP.n147 VP.t3 19.8005
R29627 VP.n147 VP.t2 19.8005
R29628 VP.n79 VP.n77 17.2148
R29629 VP.n57 VP.n4 17.2148
R29630 VP VP.n150 15.589
R29631 VP.n146 VP.n72 13.5303
R29632 VP.n143 VP.n73 12.2964
R29633 VP.n70 VP.n0 12.2964
R29634 VP.n131 VP.n79 7.37805
R29635 VP.n94 VP.n93 7.37805
R29636 VP.n19 VP.n18 7.37805
R29637 VP.n58 VP.n57 7.37805
R29638 VP.n150 VP.n149 4.80222
R29639 VP.n20 VP.n17 2.61275
R29640 VP.n95 VP.n92 2.61274
R29641 VP.n119 VP.n84 2.45968
R29642 VP.n107 VP.n106 2.45968
R29643 VP.n32 VP.n31 2.45968
R29644 VP.n45 VP.n44 2.45968
R29645 VP.n150 VP.n146 0.972091
R29646 VP.n149 VP.n148 0.716017
R29647 VP.n145 VP.n144 0.354861
R29648 VP.n72 VP.n71 0.354861
R29649 VP.n144 VP.n74 0.189894
R29650 VP.n140 VP.n74 0.189894
R29651 VP.n140 VP.n139 0.189894
R29652 VP.n139 VP.n138 0.189894
R29653 VP.n138 VP.n76 0.189894
R29654 VP.n134 VP.n76 0.189894
R29655 VP.n134 VP.n133 0.189894
R29656 VP.n133 VP.n132 0.189894
R29657 VP.n132 VP.n78 0.189894
R29658 VP.n128 VP.n78 0.189894
R29659 VP.n128 VP.n127 0.189894
R29660 VP.n127 VP.n126 0.189894
R29661 VP.n126 VP.n81 0.189894
R29662 VP.n122 VP.n81 0.189894
R29663 VP.n122 VP.n121 0.189894
R29664 VP.n121 VP.n120 0.189894
R29665 VP.n120 VP.n83 0.189894
R29666 VP.n116 VP.n83 0.189894
R29667 VP.n116 VP.n115 0.189894
R29668 VP.n115 VP.n114 0.189894
R29669 VP.n114 VP.n86 0.189894
R29670 VP.n110 VP.n86 0.189894
R29671 VP.n110 VP.n109 0.189894
R29672 VP.n109 VP.n108 0.189894
R29673 VP.n108 VP.n88 0.189894
R29674 VP.n103 VP.n88 0.189894
R29675 VP.n103 VP.n102 0.189894
R29676 VP.n102 VP.n101 0.189894
R29677 VP.n101 VP.n90 0.189894
R29678 VP.n97 VP.n90 0.189894
R29679 VP.n97 VP.n96 0.189894
R29680 VP.n96 VP.n95 0.189894
R29681 VP.n21 VP.n20 0.189894
R29682 VP.n22 VP.n21 0.189894
R29683 VP.n22 VP.n15 0.189894
R29684 VP.n26 VP.n15 0.189894
R29685 VP.n27 VP.n26 0.189894
R29686 VP.n28 VP.n27 0.189894
R29687 VP.n28 VP.n13 0.189894
R29688 VP.n33 VP.n13 0.189894
R29689 VP.n34 VP.n33 0.189894
R29690 VP.n35 VP.n34 0.189894
R29691 VP.n35 VP.n11 0.189894
R29692 VP.n39 VP.n11 0.189894
R29693 VP.n40 VP.n39 0.189894
R29694 VP.n41 VP.n40 0.189894
R29695 VP.n41 VP.n9 0.189894
R29696 VP.n46 VP.n9 0.189894
R29697 VP.n47 VP.n46 0.189894
R29698 VP.n48 VP.n47 0.189894
R29699 VP.n48 VP.n7 0.189894
R29700 VP.n52 VP.n7 0.189894
R29701 VP.n53 VP.n52 0.189894
R29702 VP.n54 VP.n53 0.189894
R29703 VP.n54 VP.n5 0.189894
R29704 VP.n59 VP.n5 0.189894
R29705 VP.n60 VP.n59 0.189894
R29706 VP.n61 VP.n60 0.189894
R29707 VP.n61 VP.n3 0.189894
R29708 VP.n65 VP.n3 0.189894
R29709 VP.n66 VP.n65 0.189894
R29710 VP.n67 VP.n66 0.189894
R29711 VP.n67 VP.n1 0.189894
R29712 VP.n71 VP.n1 0.189894
R29713 VN.n148 VN.t0 243.97
R29714 VN.n149 VN.t2 243.255
R29715 VN.n148 VN.n147 223.454
R29716 VN.n144 VN.n143 161.3
R29717 VN.n142 VN.n74 161.3
R29718 VN.n141 VN.n140 161.3
R29719 VN.n139 VN.n75 161.3
R29720 VN.n138 VN.n137 161.3
R29721 VN.n136 VN.n76 161.3
R29722 VN.n135 VN.n134 161.3
R29723 VN.n133 VN.n77 161.3
R29724 VN.n132 VN.n131 161.3
R29725 VN.n129 VN.n78 161.3
R29726 VN.n128 VN.n127 161.3
R29727 VN.n126 VN.n79 161.3
R29728 VN.n125 VN.n124 161.3
R29729 VN.n123 VN.n80 161.3
R29730 VN.n122 VN.n121 161.3
R29731 VN.n120 VN.n81 161.3
R29732 VN.n119 VN.n118 161.3
R29733 VN.n116 VN.n82 161.3
R29734 VN.n115 VN.n114 161.3
R29735 VN.n113 VN.n83 161.3
R29736 VN.n112 VN.n111 161.3
R29737 VN.n110 VN.n84 161.3
R29738 VN.n109 VN.n108 161.3
R29739 VN.n107 VN.n85 161.3
R29740 VN.n106 VN.n105 161.3
R29741 VN.n103 VN.n86 161.3
R29742 VN.n102 VN.n101 161.3
R29743 VN.n100 VN.n87 161.3
R29744 VN.n99 VN.n98 161.3
R29745 VN.n97 VN.n88 161.3
R29746 VN.n96 VN.n95 161.3
R29747 VN.n94 VN.n89 161.3
R29748 VN.n93 VN.n92 161.3
R29749 VN.n22 VN.n21 161.3
R29750 VN.n23 VN.n18 161.3
R29751 VN.n25 VN.n24 161.3
R29752 VN.n26 VN.n17 161.3
R29753 VN.n28 VN.n27 161.3
R29754 VN.n29 VN.n16 161.3
R29755 VN.n31 VN.n30 161.3
R29756 VN.n32 VN.n15 161.3
R29757 VN.n35 VN.n34 161.3
R29758 VN.n36 VN.n14 161.3
R29759 VN.n38 VN.n37 161.3
R29760 VN.n39 VN.n13 161.3
R29761 VN.n41 VN.n40 161.3
R29762 VN.n42 VN.n12 161.3
R29763 VN.n44 VN.n43 161.3
R29764 VN.n45 VN.n10 161.3
R29765 VN.n47 VN.n46 161.3
R29766 VN.n48 VN.n9 161.3
R29767 VN.n50 VN.n49 161.3
R29768 VN.n51 VN.n8 161.3
R29769 VN.n53 VN.n52 161.3
R29770 VN.n54 VN.n7 161.3
R29771 VN.n56 VN.n55 161.3
R29772 VN.n57 VN.n5 161.3
R29773 VN.n59 VN.n58 161.3
R29774 VN.n60 VN.n4 161.3
R29775 VN.n62 VN.n61 161.3
R29776 VN.n63 VN.n3 161.3
R29777 VN.n65 VN.n64 161.3
R29778 VN.n66 VN.n2 161.3
R29779 VN.n68 VN.n67 161.3
R29780 VN.n69 VN.n1 161.3
R29781 VN.n71 VN.n70 161.3
R29782 VN.n145 VN.n73 77.9496
R29783 VN.n72 VN.n0 77.9496
R29784 VN.n90 VN.t12 76.2399
R29785 VN.n19 VN.t6 76.2397
R29786 VN.n137 VN.n75 73.0308
R29787 VN.n64 VN.n2 73.0308
R29788 VN.n20 VN.n19 69.3319
R29789 VN.n91 VN.n90 69.3319
R29790 VN.n98 VN.n97 66.2494
R29791 VN.n124 VN.n79 66.2494
R29792 VN.n52 VN.n7 66.2494
R29793 VN.n27 VN.n26 66.2494
R29794 VN.n111 VN.n110 56.5617
R29795 VN.n111 VN.n83 56.5617
R29796 VN.n40 VN.n12 56.5617
R29797 VN.n40 VN.n39 56.5617
R29798 VN.n98 VN.n87 46.874
R29799 VN.n124 VN.n123 46.874
R29800 VN.n52 VN.n51 46.874
R29801 VN.n27 VN.n16 46.874
R29802 VN.n146 VN.n145 46.7121
R29803 VN.n91 VN.t4 41.7552
R29804 VN.n104 VN.t13 41.7552
R29805 VN.n117 VN.t10 41.7552
R29806 VN.n130 VN.t8 41.7552
R29807 VN.n73 VN.t15 41.7552
R29808 VN.n0 VN.t7 41.7552
R29809 VN.n6 VN.t11 41.7552
R29810 VN.n11 VN.t14 41.7552
R29811 VN.n33 VN.t5 41.7552
R29812 VN.n20 VN.t9 41.7552
R29813 VN.n137 VN.n136 37.1863
R29814 VN.n64 VN.n63 37.1863
R29815 VN.n141 VN.n75 27.4986
R29816 VN.n68 VN.n2 27.4986
R29817 VN.n92 VN.n89 24.5923
R29818 VN.n96 VN.n89 24.5923
R29819 VN.n97 VN.n96 24.5923
R29820 VN.n102 VN.n87 24.5923
R29821 VN.n103 VN.n102 24.5923
R29822 VN.n105 VN.n85 24.5923
R29823 VN.n109 VN.n85 24.5923
R29824 VN.n110 VN.n109 24.5923
R29825 VN.n115 VN.n83 24.5923
R29826 VN.n116 VN.n115 24.5923
R29827 VN.n118 VN.n116 24.5923
R29828 VN.n122 VN.n81 24.5923
R29829 VN.n123 VN.n122 24.5923
R29830 VN.n128 VN.n79 24.5923
R29831 VN.n129 VN.n128 24.5923
R29832 VN.n131 VN.n129 24.5923
R29833 VN.n135 VN.n77 24.5923
R29834 VN.n136 VN.n135 24.5923
R29835 VN.n142 VN.n141 24.5923
R29836 VN.n143 VN.n142 24.5923
R29837 VN.n70 VN.n69 24.5923
R29838 VN.n69 VN.n68 24.5923
R29839 VN.n63 VN.n62 24.5923
R29840 VN.n62 VN.n4 24.5923
R29841 VN.n58 VN.n57 24.5923
R29842 VN.n57 VN.n56 24.5923
R29843 VN.n56 VN.n7 24.5923
R29844 VN.n51 VN.n50 24.5923
R29845 VN.n50 VN.n9 24.5923
R29846 VN.n46 VN.n45 24.5923
R29847 VN.n45 VN.n44 24.5923
R29848 VN.n44 VN.n12 24.5923
R29849 VN.n39 VN.n38 24.5923
R29850 VN.n38 VN.n14 24.5923
R29851 VN.n34 VN.n14 24.5923
R29852 VN.n32 VN.n31 24.5923
R29853 VN.n31 VN.n16 24.5923
R29854 VN.n26 VN.n25 24.5923
R29855 VN.n25 VN.n18 24.5923
R29856 VN.n21 VN.n18 24.5923
R29857 VN.n104 VN.n103 22.1332
R29858 VN.n117 VN.n81 22.1332
R29859 VN.n11 VN.n9 22.1332
R29860 VN.n33 VN.n32 22.1332
R29861 VN VN.n150 20.7475
R29862 VN.n147 VN.t3 19.8005
R29863 VN.n147 VN.t1 19.8005
R29864 VN.n130 VN.n77 17.2148
R29865 VN.n6 VN.n4 17.2148
R29866 VN.n146 VN.n72 13.3144
R29867 VN.n143 VN.n73 12.2964
R29868 VN.n70 VN.n0 12.2964
R29869 VN.n92 VN.n91 7.37805
R29870 VN.n131 VN.n130 7.37805
R29871 VN.n58 VN.n6 7.37805
R29872 VN.n21 VN.n20 7.37805
R29873 VN.n150 VN.n149 5.04791
R29874 VN.n93 VN.n90 2.61275
R29875 VN.n22 VN.n19 2.61274
R29876 VN.n105 VN.n104 2.45968
R29877 VN.n118 VN.n117 2.45968
R29878 VN.n46 VN.n11 2.45968
R29879 VN.n34 VN.n33 2.45968
R29880 VN.n150 VN.n146 1.188
R29881 VN.n149 VN.n148 0.716017
R29882 VN.n145 VN.n144 0.354861
R29883 VN.n72 VN.n71 0.354861
R29884 VN.n94 VN.n93 0.189894
R29885 VN.n95 VN.n94 0.189894
R29886 VN.n95 VN.n88 0.189894
R29887 VN.n99 VN.n88 0.189894
R29888 VN.n100 VN.n99 0.189894
R29889 VN.n101 VN.n100 0.189894
R29890 VN.n101 VN.n86 0.189894
R29891 VN.n106 VN.n86 0.189894
R29892 VN.n107 VN.n106 0.189894
R29893 VN.n108 VN.n107 0.189894
R29894 VN.n108 VN.n84 0.189894
R29895 VN.n112 VN.n84 0.189894
R29896 VN.n113 VN.n112 0.189894
R29897 VN.n114 VN.n113 0.189894
R29898 VN.n114 VN.n82 0.189894
R29899 VN.n119 VN.n82 0.189894
R29900 VN.n120 VN.n119 0.189894
R29901 VN.n121 VN.n120 0.189894
R29902 VN.n121 VN.n80 0.189894
R29903 VN.n125 VN.n80 0.189894
R29904 VN.n126 VN.n125 0.189894
R29905 VN.n127 VN.n126 0.189894
R29906 VN.n127 VN.n78 0.189894
R29907 VN.n132 VN.n78 0.189894
R29908 VN.n133 VN.n132 0.189894
R29909 VN.n134 VN.n133 0.189894
R29910 VN.n134 VN.n76 0.189894
R29911 VN.n138 VN.n76 0.189894
R29912 VN.n139 VN.n138 0.189894
R29913 VN.n140 VN.n139 0.189894
R29914 VN.n140 VN.n74 0.189894
R29915 VN.n144 VN.n74 0.189894
R29916 VN.n71 VN.n1 0.189894
R29917 VN.n67 VN.n1 0.189894
R29918 VN.n67 VN.n66 0.189894
R29919 VN.n66 VN.n65 0.189894
R29920 VN.n65 VN.n3 0.189894
R29921 VN.n61 VN.n3 0.189894
R29922 VN.n61 VN.n60 0.189894
R29923 VN.n60 VN.n59 0.189894
R29924 VN.n59 VN.n5 0.189894
R29925 VN.n55 VN.n5 0.189894
R29926 VN.n55 VN.n54 0.189894
R29927 VN.n54 VN.n53 0.189894
R29928 VN.n53 VN.n8 0.189894
R29929 VN.n49 VN.n8 0.189894
R29930 VN.n49 VN.n48 0.189894
R29931 VN.n48 VN.n47 0.189894
R29932 VN.n47 VN.n10 0.189894
R29933 VN.n43 VN.n10 0.189894
R29934 VN.n43 VN.n42 0.189894
R29935 VN.n42 VN.n41 0.189894
R29936 VN.n41 VN.n13 0.189894
R29937 VN.n37 VN.n13 0.189894
R29938 VN.n37 VN.n36 0.189894
R29939 VN.n36 VN.n35 0.189894
R29940 VN.n35 VN.n15 0.189894
R29941 VN.n30 VN.n15 0.189894
R29942 VN.n30 VN.n29 0.189894
R29943 VN.n29 VN.n28 0.189894
R29944 VN.n28 VN.n17 0.189894
R29945 VN.n24 VN.n17 0.189894
R29946 VN.n24 VN.n23 0.189894
R29947 VN.n23 VN.n22 0.189894
R29948 CS_BIAS.n823 CS_BIAS.n663 161.3
R29949 CS_BIAS.n822 CS_BIAS.n821 161.3
R29950 CS_BIAS.n820 CS_BIAS.n664 161.3
R29951 CS_BIAS.n819 CS_BIAS.n818 161.3
R29952 CS_BIAS.n817 CS_BIAS.n665 161.3
R29953 CS_BIAS.n816 CS_BIAS.n815 161.3
R29954 CS_BIAS.n814 CS_BIAS.n666 161.3
R29955 CS_BIAS.n813 CS_BIAS.n812 161.3
R29956 CS_BIAS.n811 CS_BIAS.n667 161.3
R29957 CS_BIAS.n810 CS_BIAS.n809 161.3
R29958 CS_BIAS.n808 CS_BIAS.n668 161.3
R29959 CS_BIAS.n807 CS_BIAS.n806 161.3
R29960 CS_BIAS.n805 CS_BIAS.n669 161.3
R29961 CS_BIAS.n803 CS_BIAS.n802 161.3
R29962 CS_BIAS.n801 CS_BIAS.n670 161.3
R29963 CS_BIAS.n800 CS_BIAS.n799 161.3
R29964 CS_BIAS.n798 CS_BIAS.n671 161.3
R29965 CS_BIAS.n797 CS_BIAS.n796 161.3
R29966 CS_BIAS.n795 CS_BIAS.n672 161.3
R29967 CS_BIAS.n794 CS_BIAS.n793 161.3
R29968 CS_BIAS.n792 CS_BIAS.n673 161.3
R29969 CS_BIAS.n791 CS_BIAS.n790 161.3
R29970 CS_BIAS.n789 CS_BIAS.n674 161.3
R29971 CS_BIAS.n788 CS_BIAS.n787 161.3
R29972 CS_BIAS.n786 CS_BIAS.n675 161.3
R29973 CS_BIAS.n785 CS_BIAS.n784 161.3
R29974 CS_BIAS.n783 CS_BIAS.n782 161.3
R29975 CS_BIAS.n781 CS_BIAS.n677 161.3
R29976 CS_BIAS.n780 CS_BIAS.n779 161.3
R29977 CS_BIAS.n778 CS_BIAS.n678 161.3
R29978 CS_BIAS.n777 CS_BIAS.n776 161.3
R29979 CS_BIAS.n775 CS_BIAS.n679 161.3
R29980 CS_BIAS.n774 CS_BIAS.n773 161.3
R29981 CS_BIAS.n772 CS_BIAS.n680 161.3
R29982 CS_BIAS.n771 CS_BIAS.n770 161.3
R29983 CS_BIAS.n769 CS_BIAS.n681 161.3
R29984 CS_BIAS.n768 CS_BIAS.n767 161.3
R29985 CS_BIAS.n766 CS_BIAS.n682 161.3
R29986 CS_BIAS.n765 CS_BIAS.n764 161.3
R29987 CS_BIAS.n762 CS_BIAS.n683 161.3
R29988 CS_BIAS.n761 CS_BIAS.n760 161.3
R29989 CS_BIAS.n759 CS_BIAS.n684 161.3
R29990 CS_BIAS.n758 CS_BIAS.n757 161.3
R29991 CS_BIAS.n756 CS_BIAS.n685 161.3
R29992 CS_BIAS.n755 CS_BIAS.n754 161.3
R29993 CS_BIAS.n753 CS_BIAS.n686 161.3
R29994 CS_BIAS.n752 CS_BIAS.n751 161.3
R29995 CS_BIAS.n750 CS_BIAS.n687 161.3
R29996 CS_BIAS.n749 CS_BIAS.n748 161.3
R29997 CS_BIAS.n747 CS_BIAS.n688 161.3
R29998 CS_BIAS.n746 CS_BIAS.n745 161.3
R29999 CS_BIAS.n743 CS_BIAS.n689 161.3
R30000 CS_BIAS.n742 CS_BIAS.n741 161.3
R30001 CS_BIAS.n740 CS_BIAS.n690 161.3
R30002 CS_BIAS.n739 CS_BIAS.n738 161.3
R30003 CS_BIAS.n737 CS_BIAS.n691 161.3
R30004 CS_BIAS.n736 CS_BIAS.n735 161.3
R30005 CS_BIAS.n734 CS_BIAS.n692 161.3
R30006 CS_BIAS.n733 CS_BIAS.n732 161.3
R30007 CS_BIAS.n731 CS_BIAS.n693 161.3
R30008 CS_BIAS.n730 CS_BIAS.n729 161.3
R30009 CS_BIAS.n728 CS_BIAS.n694 161.3
R30010 CS_BIAS.n727 CS_BIAS.n726 161.3
R30011 CS_BIAS.n725 CS_BIAS.n695 161.3
R30012 CS_BIAS.n723 CS_BIAS.n722 161.3
R30013 CS_BIAS.n721 CS_BIAS.n696 161.3
R30014 CS_BIAS.n720 CS_BIAS.n719 161.3
R30015 CS_BIAS.n718 CS_BIAS.n697 161.3
R30016 CS_BIAS.n717 CS_BIAS.n716 161.3
R30017 CS_BIAS.n715 CS_BIAS.n698 161.3
R30018 CS_BIAS.n714 CS_BIAS.n713 161.3
R30019 CS_BIAS.n712 CS_BIAS.n699 161.3
R30020 CS_BIAS.n711 CS_BIAS.n710 161.3
R30021 CS_BIAS.n709 CS_BIAS.n700 161.3
R30022 CS_BIAS.n708 CS_BIAS.n707 161.3
R30023 CS_BIAS.n706 CS_BIAS.n701 161.3
R30024 CS_BIAS.n705 CS_BIAS.n704 161.3
R30025 CS_BIAS.n541 CS_BIAS.n540 161.3
R30026 CS_BIAS.n542 CS_BIAS.n537 161.3
R30027 CS_BIAS.n544 CS_BIAS.n543 161.3
R30028 CS_BIAS.n545 CS_BIAS.n536 161.3
R30029 CS_BIAS.n547 CS_BIAS.n546 161.3
R30030 CS_BIAS.n548 CS_BIAS.n535 161.3
R30031 CS_BIAS.n550 CS_BIAS.n549 161.3
R30032 CS_BIAS.n551 CS_BIAS.n534 161.3
R30033 CS_BIAS.n553 CS_BIAS.n552 161.3
R30034 CS_BIAS.n554 CS_BIAS.n533 161.3
R30035 CS_BIAS.n556 CS_BIAS.n555 161.3
R30036 CS_BIAS.n557 CS_BIAS.n532 161.3
R30037 CS_BIAS.n559 CS_BIAS.n558 161.3
R30038 CS_BIAS.n561 CS_BIAS.n531 161.3
R30039 CS_BIAS.n563 CS_BIAS.n562 161.3
R30040 CS_BIAS.n564 CS_BIAS.n530 161.3
R30041 CS_BIAS.n566 CS_BIAS.n565 161.3
R30042 CS_BIAS.n567 CS_BIAS.n529 161.3
R30043 CS_BIAS.n569 CS_BIAS.n568 161.3
R30044 CS_BIAS.n570 CS_BIAS.n528 161.3
R30045 CS_BIAS.n572 CS_BIAS.n571 161.3
R30046 CS_BIAS.n573 CS_BIAS.n527 161.3
R30047 CS_BIAS.n575 CS_BIAS.n574 161.3
R30048 CS_BIAS.n576 CS_BIAS.n526 161.3
R30049 CS_BIAS.n578 CS_BIAS.n577 161.3
R30050 CS_BIAS.n579 CS_BIAS.n525 161.3
R30051 CS_BIAS.n582 CS_BIAS.n581 161.3
R30052 CS_BIAS.n583 CS_BIAS.n524 161.3
R30053 CS_BIAS.n585 CS_BIAS.n584 161.3
R30054 CS_BIAS.n586 CS_BIAS.n523 161.3
R30055 CS_BIAS.n588 CS_BIAS.n587 161.3
R30056 CS_BIAS.n589 CS_BIAS.n522 161.3
R30057 CS_BIAS.n591 CS_BIAS.n590 161.3
R30058 CS_BIAS.n592 CS_BIAS.n521 161.3
R30059 CS_BIAS.n594 CS_BIAS.n593 161.3
R30060 CS_BIAS.n595 CS_BIAS.n520 161.3
R30061 CS_BIAS.n597 CS_BIAS.n596 161.3
R30062 CS_BIAS.n598 CS_BIAS.n519 161.3
R30063 CS_BIAS.n601 CS_BIAS.n600 161.3
R30064 CS_BIAS.n602 CS_BIAS.n518 161.3
R30065 CS_BIAS.n604 CS_BIAS.n603 161.3
R30066 CS_BIAS.n605 CS_BIAS.n517 161.3
R30067 CS_BIAS.n607 CS_BIAS.n606 161.3
R30068 CS_BIAS.n608 CS_BIAS.n516 161.3
R30069 CS_BIAS.n610 CS_BIAS.n609 161.3
R30070 CS_BIAS.n611 CS_BIAS.n515 161.3
R30071 CS_BIAS.n613 CS_BIAS.n612 161.3
R30072 CS_BIAS.n614 CS_BIAS.n514 161.3
R30073 CS_BIAS.n616 CS_BIAS.n615 161.3
R30074 CS_BIAS.n617 CS_BIAS.n513 161.3
R30075 CS_BIAS.n619 CS_BIAS.n618 161.3
R30076 CS_BIAS.n621 CS_BIAS.n620 161.3
R30077 CS_BIAS.n622 CS_BIAS.n511 161.3
R30078 CS_BIAS.n624 CS_BIAS.n623 161.3
R30079 CS_BIAS.n625 CS_BIAS.n510 161.3
R30080 CS_BIAS.n627 CS_BIAS.n626 161.3
R30081 CS_BIAS.n628 CS_BIAS.n509 161.3
R30082 CS_BIAS.n630 CS_BIAS.n629 161.3
R30083 CS_BIAS.n631 CS_BIAS.n508 161.3
R30084 CS_BIAS.n633 CS_BIAS.n632 161.3
R30085 CS_BIAS.n634 CS_BIAS.n507 161.3
R30086 CS_BIAS.n636 CS_BIAS.n635 161.3
R30087 CS_BIAS.n637 CS_BIAS.n506 161.3
R30088 CS_BIAS.n639 CS_BIAS.n638 161.3
R30089 CS_BIAS.n641 CS_BIAS.n505 161.3
R30090 CS_BIAS.n643 CS_BIAS.n642 161.3
R30091 CS_BIAS.n644 CS_BIAS.n504 161.3
R30092 CS_BIAS.n646 CS_BIAS.n645 161.3
R30093 CS_BIAS.n647 CS_BIAS.n503 161.3
R30094 CS_BIAS.n649 CS_BIAS.n648 161.3
R30095 CS_BIAS.n650 CS_BIAS.n502 161.3
R30096 CS_BIAS.n652 CS_BIAS.n651 161.3
R30097 CS_BIAS.n653 CS_BIAS.n501 161.3
R30098 CS_BIAS.n655 CS_BIAS.n654 161.3
R30099 CS_BIAS.n656 CS_BIAS.n500 161.3
R30100 CS_BIAS.n658 CS_BIAS.n657 161.3
R30101 CS_BIAS.n659 CS_BIAS.n499 161.3
R30102 CS_BIAS.n377 CS_BIAS.n376 161.3
R30103 CS_BIAS.n378 CS_BIAS.n373 161.3
R30104 CS_BIAS.n380 CS_BIAS.n379 161.3
R30105 CS_BIAS.n381 CS_BIAS.n372 161.3
R30106 CS_BIAS.n383 CS_BIAS.n382 161.3
R30107 CS_BIAS.n384 CS_BIAS.n371 161.3
R30108 CS_BIAS.n386 CS_BIAS.n385 161.3
R30109 CS_BIAS.n387 CS_BIAS.n370 161.3
R30110 CS_BIAS.n389 CS_BIAS.n388 161.3
R30111 CS_BIAS.n390 CS_BIAS.n369 161.3
R30112 CS_BIAS.n392 CS_BIAS.n391 161.3
R30113 CS_BIAS.n393 CS_BIAS.n368 161.3
R30114 CS_BIAS.n395 CS_BIAS.n394 161.3
R30115 CS_BIAS.n397 CS_BIAS.n367 161.3
R30116 CS_BIAS.n399 CS_BIAS.n398 161.3
R30117 CS_BIAS.n400 CS_BIAS.n366 161.3
R30118 CS_BIAS.n402 CS_BIAS.n401 161.3
R30119 CS_BIAS.n403 CS_BIAS.n365 161.3
R30120 CS_BIAS.n405 CS_BIAS.n404 161.3
R30121 CS_BIAS.n406 CS_BIAS.n364 161.3
R30122 CS_BIAS.n408 CS_BIAS.n407 161.3
R30123 CS_BIAS.n409 CS_BIAS.n363 161.3
R30124 CS_BIAS.n411 CS_BIAS.n410 161.3
R30125 CS_BIAS.n412 CS_BIAS.n362 161.3
R30126 CS_BIAS.n414 CS_BIAS.n413 161.3
R30127 CS_BIAS.n415 CS_BIAS.n361 161.3
R30128 CS_BIAS.n418 CS_BIAS.n417 161.3
R30129 CS_BIAS.n419 CS_BIAS.n360 161.3
R30130 CS_BIAS.n421 CS_BIAS.n420 161.3
R30131 CS_BIAS.n422 CS_BIAS.n359 161.3
R30132 CS_BIAS.n424 CS_BIAS.n423 161.3
R30133 CS_BIAS.n425 CS_BIAS.n358 161.3
R30134 CS_BIAS.n427 CS_BIAS.n426 161.3
R30135 CS_BIAS.n428 CS_BIAS.n357 161.3
R30136 CS_BIAS.n430 CS_BIAS.n429 161.3
R30137 CS_BIAS.n431 CS_BIAS.n356 161.3
R30138 CS_BIAS.n433 CS_BIAS.n432 161.3
R30139 CS_BIAS.n434 CS_BIAS.n355 161.3
R30140 CS_BIAS.n437 CS_BIAS.n436 161.3
R30141 CS_BIAS.n438 CS_BIAS.n354 161.3
R30142 CS_BIAS.n440 CS_BIAS.n439 161.3
R30143 CS_BIAS.n441 CS_BIAS.n353 161.3
R30144 CS_BIAS.n443 CS_BIAS.n442 161.3
R30145 CS_BIAS.n444 CS_BIAS.n352 161.3
R30146 CS_BIAS.n446 CS_BIAS.n445 161.3
R30147 CS_BIAS.n447 CS_BIAS.n351 161.3
R30148 CS_BIAS.n449 CS_BIAS.n448 161.3
R30149 CS_BIAS.n450 CS_BIAS.n350 161.3
R30150 CS_BIAS.n452 CS_BIAS.n451 161.3
R30151 CS_BIAS.n453 CS_BIAS.n349 161.3
R30152 CS_BIAS.n455 CS_BIAS.n454 161.3
R30153 CS_BIAS.n457 CS_BIAS.n456 161.3
R30154 CS_BIAS.n458 CS_BIAS.n347 161.3
R30155 CS_BIAS.n460 CS_BIAS.n459 161.3
R30156 CS_BIAS.n461 CS_BIAS.n346 161.3
R30157 CS_BIAS.n463 CS_BIAS.n462 161.3
R30158 CS_BIAS.n464 CS_BIAS.n345 161.3
R30159 CS_BIAS.n466 CS_BIAS.n465 161.3
R30160 CS_BIAS.n467 CS_BIAS.n344 161.3
R30161 CS_BIAS.n469 CS_BIAS.n468 161.3
R30162 CS_BIAS.n470 CS_BIAS.n343 161.3
R30163 CS_BIAS.n472 CS_BIAS.n471 161.3
R30164 CS_BIAS.n473 CS_BIAS.n342 161.3
R30165 CS_BIAS.n475 CS_BIAS.n474 161.3
R30166 CS_BIAS.n477 CS_BIAS.n341 161.3
R30167 CS_BIAS.n479 CS_BIAS.n478 161.3
R30168 CS_BIAS.n480 CS_BIAS.n340 161.3
R30169 CS_BIAS.n482 CS_BIAS.n481 161.3
R30170 CS_BIAS.n483 CS_BIAS.n339 161.3
R30171 CS_BIAS.n485 CS_BIAS.n484 161.3
R30172 CS_BIAS.n486 CS_BIAS.n338 161.3
R30173 CS_BIAS.n488 CS_BIAS.n487 161.3
R30174 CS_BIAS.n489 CS_BIAS.n337 161.3
R30175 CS_BIAS.n491 CS_BIAS.n490 161.3
R30176 CS_BIAS.n492 CS_BIAS.n336 161.3
R30177 CS_BIAS.n494 CS_BIAS.n493 161.3
R30178 CS_BIAS.n495 CS_BIAS.n335 161.3
R30179 CS_BIAS.n133 CS_BIAS.n132 161.3
R30180 CS_BIAS.n134 CS_BIAS.n129 161.3
R30181 CS_BIAS.n136 CS_BIAS.n135 161.3
R30182 CS_BIAS.n137 CS_BIAS.n128 161.3
R30183 CS_BIAS.n139 CS_BIAS.n138 161.3
R30184 CS_BIAS.n140 CS_BIAS.n127 161.3
R30185 CS_BIAS.n142 CS_BIAS.n141 161.3
R30186 CS_BIAS.n143 CS_BIAS.n126 161.3
R30187 CS_BIAS.n145 CS_BIAS.n144 161.3
R30188 CS_BIAS.n146 CS_BIAS.n125 161.3
R30189 CS_BIAS.n148 CS_BIAS.n147 161.3
R30190 CS_BIAS.n149 CS_BIAS.n124 161.3
R30191 CS_BIAS.n151 CS_BIAS.n150 161.3
R30192 CS_BIAS.n153 CS_BIAS.n123 161.3
R30193 CS_BIAS.n155 CS_BIAS.n154 161.3
R30194 CS_BIAS.n156 CS_BIAS.n122 161.3
R30195 CS_BIAS.n158 CS_BIAS.n157 161.3
R30196 CS_BIAS.n159 CS_BIAS.n121 161.3
R30197 CS_BIAS.n161 CS_BIAS.n160 161.3
R30198 CS_BIAS.n162 CS_BIAS.n120 161.3
R30199 CS_BIAS.n164 CS_BIAS.n163 161.3
R30200 CS_BIAS.n165 CS_BIAS.n119 161.3
R30201 CS_BIAS.n167 CS_BIAS.n166 161.3
R30202 CS_BIAS.n168 CS_BIAS.n118 161.3
R30203 CS_BIAS.n170 CS_BIAS.n169 161.3
R30204 CS_BIAS.n171 CS_BIAS.n117 161.3
R30205 CS_BIAS.n174 CS_BIAS.n173 161.3
R30206 CS_BIAS.n175 CS_BIAS.n116 161.3
R30207 CS_BIAS.n177 CS_BIAS.n176 161.3
R30208 CS_BIAS.n178 CS_BIAS.n115 161.3
R30209 CS_BIAS.n180 CS_BIAS.n179 161.3
R30210 CS_BIAS.n181 CS_BIAS.n114 161.3
R30211 CS_BIAS.n183 CS_BIAS.n182 161.3
R30212 CS_BIAS.n184 CS_BIAS.n113 161.3
R30213 CS_BIAS.n186 CS_BIAS.n185 161.3
R30214 CS_BIAS.n187 CS_BIAS.n112 161.3
R30215 CS_BIAS.n189 CS_BIAS.n188 161.3
R30216 CS_BIAS.n190 CS_BIAS.n111 161.3
R30217 CS_BIAS.n193 CS_BIAS.n192 161.3
R30218 CS_BIAS.n194 CS_BIAS.n110 161.3
R30219 CS_BIAS.n196 CS_BIAS.n195 161.3
R30220 CS_BIAS.n197 CS_BIAS.n109 161.3
R30221 CS_BIAS.n199 CS_BIAS.n198 161.3
R30222 CS_BIAS.n200 CS_BIAS.n108 161.3
R30223 CS_BIAS.n202 CS_BIAS.n201 161.3
R30224 CS_BIAS.n203 CS_BIAS.n107 161.3
R30225 CS_BIAS.n205 CS_BIAS.n204 161.3
R30226 CS_BIAS.n206 CS_BIAS.n106 161.3
R30227 CS_BIAS.n208 CS_BIAS.n207 161.3
R30228 CS_BIAS.n209 CS_BIAS.n105 161.3
R30229 CS_BIAS.n211 CS_BIAS.n210 161.3
R30230 CS_BIAS.n213 CS_BIAS.n212 161.3
R30231 CS_BIAS.n214 CS_BIAS.n103 161.3
R30232 CS_BIAS.n216 CS_BIAS.n215 161.3
R30233 CS_BIAS.n217 CS_BIAS.n102 161.3
R30234 CS_BIAS.n219 CS_BIAS.n218 161.3
R30235 CS_BIAS.n220 CS_BIAS.n101 161.3
R30236 CS_BIAS.n222 CS_BIAS.n221 161.3
R30237 CS_BIAS.n223 CS_BIAS.n100 161.3
R30238 CS_BIAS.n225 CS_BIAS.n224 161.3
R30239 CS_BIAS.n226 CS_BIAS.n99 161.3
R30240 CS_BIAS.n228 CS_BIAS.n227 161.3
R30241 CS_BIAS.n229 CS_BIAS.n98 161.3
R30242 CS_BIAS.n231 CS_BIAS.n230 161.3
R30243 CS_BIAS.n233 CS_BIAS.n97 161.3
R30244 CS_BIAS.n235 CS_BIAS.n234 161.3
R30245 CS_BIAS.n236 CS_BIAS.n96 161.3
R30246 CS_BIAS.n238 CS_BIAS.n237 161.3
R30247 CS_BIAS.n239 CS_BIAS.n95 161.3
R30248 CS_BIAS.n241 CS_BIAS.n240 161.3
R30249 CS_BIAS.n242 CS_BIAS.n94 161.3
R30250 CS_BIAS.n244 CS_BIAS.n243 161.3
R30251 CS_BIAS.n245 CS_BIAS.n93 161.3
R30252 CS_BIAS.n247 CS_BIAS.n246 161.3
R30253 CS_BIAS.n248 CS_BIAS.n92 161.3
R30254 CS_BIAS.n250 CS_BIAS.n249 161.3
R30255 CS_BIAS.n251 CS_BIAS.n91 161.3
R30256 CS_BIAS.n42 CS_BIAS.n41 161.3
R30257 CS_BIAS.n43 CS_BIAS.n38 161.3
R30258 CS_BIAS.n45 CS_BIAS.n44 161.3
R30259 CS_BIAS.n46 CS_BIAS.n37 161.3
R30260 CS_BIAS.n48 CS_BIAS.n47 161.3
R30261 CS_BIAS.n49 CS_BIAS.n36 161.3
R30262 CS_BIAS.n51 CS_BIAS.n50 161.3
R30263 CS_BIAS.n52 CS_BIAS.n35 161.3
R30264 CS_BIAS.n54 CS_BIAS.n53 161.3
R30265 CS_BIAS.n55 CS_BIAS.n34 161.3
R30266 CS_BIAS.n57 CS_BIAS.n56 161.3
R30267 CS_BIAS.n58 CS_BIAS.n33 161.3
R30268 CS_BIAS.n60 CS_BIAS.n59 161.3
R30269 CS_BIAS.n62 CS_BIAS.n32 161.3
R30270 CS_BIAS.n64 CS_BIAS.n63 161.3
R30271 CS_BIAS.n65 CS_BIAS.n31 161.3
R30272 CS_BIAS.n67 CS_BIAS.n66 161.3
R30273 CS_BIAS.n68 CS_BIAS.n30 161.3
R30274 CS_BIAS.n70 CS_BIAS.n69 161.3
R30275 CS_BIAS.n71 CS_BIAS.n29 161.3
R30276 CS_BIAS.n73 CS_BIAS.n72 161.3
R30277 CS_BIAS.n74 CS_BIAS.n28 161.3
R30278 CS_BIAS.n76 CS_BIAS.n75 161.3
R30279 CS_BIAS.n77 CS_BIAS.n27 161.3
R30280 CS_BIAS.n79 CS_BIAS.n78 161.3
R30281 CS_BIAS.n80 CS_BIAS.n26 161.3
R30282 CS_BIAS.n83 CS_BIAS.n82 161.3
R30283 CS_BIAS.n84 CS_BIAS.n25 161.3
R30284 CS_BIAS.n86 CS_BIAS.n85 161.3
R30285 CS_BIAS.n87 CS_BIAS.n24 161.3
R30286 CS_BIAS.n89 CS_BIAS.n88 161.3
R30287 CS_BIAS.n90 CS_BIAS.n23 161.3
R30288 CS_BIAS.n264 CS_BIAS.n263 161.3
R30289 CS_BIAS.n265 CS_BIAS.n22 161.3
R30290 CS_BIAS.n267 CS_BIAS.n266 161.3
R30291 CS_BIAS.n268 CS_BIAS.n21 161.3
R30292 CS_BIAS.n270 CS_BIAS.n269 161.3
R30293 CS_BIAS.n271 CS_BIAS.n20 161.3
R30294 CS_BIAS.n274 CS_BIAS.n273 161.3
R30295 CS_BIAS.n275 CS_BIAS.n19 161.3
R30296 CS_BIAS.n277 CS_BIAS.n276 161.3
R30297 CS_BIAS.n278 CS_BIAS.n18 161.3
R30298 CS_BIAS.n280 CS_BIAS.n279 161.3
R30299 CS_BIAS.n281 CS_BIAS.n17 161.3
R30300 CS_BIAS.n283 CS_BIAS.n282 161.3
R30301 CS_BIAS.n284 CS_BIAS.n16 161.3
R30302 CS_BIAS.n286 CS_BIAS.n285 161.3
R30303 CS_BIAS.n287 CS_BIAS.n15 161.3
R30304 CS_BIAS.n289 CS_BIAS.n288 161.3
R30305 CS_BIAS.n290 CS_BIAS.n14 161.3
R30306 CS_BIAS.n292 CS_BIAS.n291 161.3
R30307 CS_BIAS.n294 CS_BIAS.n293 161.3
R30308 CS_BIAS.n295 CS_BIAS.n12 161.3
R30309 CS_BIAS.n297 CS_BIAS.n296 161.3
R30310 CS_BIAS.n298 CS_BIAS.n11 161.3
R30311 CS_BIAS.n300 CS_BIAS.n299 161.3
R30312 CS_BIAS.n301 CS_BIAS.n10 161.3
R30313 CS_BIAS.n303 CS_BIAS.n302 161.3
R30314 CS_BIAS.n304 CS_BIAS.n9 161.3
R30315 CS_BIAS.n306 CS_BIAS.n305 161.3
R30316 CS_BIAS.n307 CS_BIAS.n8 161.3
R30317 CS_BIAS.n309 CS_BIAS.n308 161.3
R30318 CS_BIAS.n310 CS_BIAS.n7 161.3
R30319 CS_BIAS.n312 CS_BIAS.n311 161.3
R30320 CS_BIAS.n314 CS_BIAS.n6 161.3
R30321 CS_BIAS.n316 CS_BIAS.n315 161.3
R30322 CS_BIAS.n317 CS_BIAS.n5 161.3
R30323 CS_BIAS.n319 CS_BIAS.n318 161.3
R30324 CS_BIAS.n320 CS_BIAS.n4 161.3
R30325 CS_BIAS.n322 CS_BIAS.n321 161.3
R30326 CS_BIAS.n323 CS_BIAS.n3 161.3
R30327 CS_BIAS.n325 CS_BIAS.n324 161.3
R30328 CS_BIAS.n326 CS_BIAS.n2 161.3
R30329 CS_BIAS.n328 CS_BIAS.n327 161.3
R30330 CS_BIAS.n329 CS_BIAS.n1 161.3
R30331 CS_BIAS.n331 CS_BIAS.n330 161.3
R30332 CS_BIAS.n332 CS_BIAS.n0 161.3
R30333 CS_BIAS.n1650 CS_BIAS.n1490 161.3
R30334 CS_BIAS.n1649 CS_BIAS.n1648 161.3
R30335 CS_BIAS.n1647 CS_BIAS.n1491 161.3
R30336 CS_BIAS.n1646 CS_BIAS.n1645 161.3
R30337 CS_BIAS.n1644 CS_BIAS.n1492 161.3
R30338 CS_BIAS.n1643 CS_BIAS.n1642 161.3
R30339 CS_BIAS.n1641 CS_BIAS.n1493 161.3
R30340 CS_BIAS.n1640 CS_BIAS.n1639 161.3
R30341 CS_BIAS.n1638 CS_BIAS.n1494 161.3
R30342 CS_BIAS.n1637 CS_BIAS.n1636 161.3
R30343 CS_BIAS.n1635 CS_BIAS.n1495 161.3
R30344 CS_BIAS.n1634 CS_BIAS.n1633 161.3
R30345 CS_BIAS.n1632 CS_BIAS.n1496 161.3
R30346 CS_BIAS.n1630 CS_BIAS.n1629 161.3
R30347 CS_BIAS.n1628 CS_BIAS.n1497 161.3
R30348 CS_BIAS.n1627 CS_BIAS.n1626 161.3
R30349 CS_BIAS.n1625 CS_BIAS.n1498 161.3
R30350 CS_BIAS.n1624 CS_BIAS.n1623 161.3
R30351 CS_BIAS.n1622 CS_BIAS.n1499 161.3
R30352 CS_BIAS.n1621 CS_BIAS.n1620 161.3
R30353 CS_BIAS.n1619 CS_BIAS.n1500 161.3
R30354 CS_BIAS.n1618 CS_BIAS.n1617 161.3
R30355 CS_BIAS.n1616 CS_BIAS.n1501 161.3
R30356 CS_BIAS.n1615 CS_BIAS.n1614 161.3
R30357 CS_BIAS.n1613 CS_BIAS.n1502 161.3
R30358 CS_BIAS.n1612 CS_BIAS.n1611 161.3
R30359 CS_BIAS.n1610 CS_BIAS.n1609 161.3
R30360 CS_BIAS.n1608 CS_BIAS.n1504 161.3
R30361 CS_BIAS.n1607 CS_BIAS.n1606 161.3
R30362 CS_BIAS.n1605 CS_BIAS.n1505 161.3
R30363 CS_BIAS.n1604 CS_BIAS.n1603 161.3
R30364 CS_BIAS.n1602 CS_BIAS.n1506 161.3
R30365 CS_BIAS.n1601 CS_BIAS.n1600 161.3
R30366 CS_BIAS.n1599 CS_BIAS.n1507 161.3
R30367 CS_BIAS.n1598 CS_BIAS.n1597 161.3
R30368 CS_BIAS.n1596 CS_BIAS.n1508 161.3
R30369 CS_BIAS.n1595 CS_BIAS.n1594 161.3
R30370 CS_BIAS.n1593 CS_BIAS.n1509 161.3
R30371 CS_BIAS.n1592 CS_BIAS.n1591 161.3
R30372 CS_BIAS.n1589 CS_BIAS.n1510 161.3
R30373 CS_BIAS.n1588 CS_BIAS.n1587 161.3
R30374 CS_BIAS.n1586 CS_BIAS.n1511 161.3
R30375 CS_BIAS.n1585 CS_BIAS.n1584 161.3
R30376 CS_BIAS.n1583 CS_BIAS.n1512 161.3
R30377 CS_BIAS.n1582 CS_BIAS.n1581 161.3
R30378 CS_BIAS.n1580 CS_BIAS.n1513 161.3
R30379 CS_BIAS.n1579 CS_BIAS.n1578 161.3
R30380 CS_BIAS.n1577 CS_BIAS.n1514 161.3
R30381 CS_BIAS.n1576 CS_BIAS.n1575 161.3
R30382 CS_BIAS.n1574 CS_BIAS.n1515 161.3
R30383 CS_BIAS.n1573 CS_BIAS.n1572 161.3
R30384 CS_BIAS.n1570 CS_BIAS.n1516 161.3
R30385 CS_BIAS.n1569 CS_BIAS.n1568 161.3
R30386 CS_BIAS.n1567 CS_BIAS.n1517 161.3
R30387 CS_BIAS.n1566 CS_BIAS.n1565 161.3
R30388 CS_BIAS.n1564 CS_BIAS.n1518 161.3
R30389 CS_BIAS.n1563 CS_BIAS.n1562 161.3
R30390 CS_BIAS.n1561 CS_BIAS.n1519 161.3
R30391 CS_BIAS.n1560 CS_BIAS.n1559 161.3
R30392 CS_BIAS.n1558 CS_BIAS.n1520 161.3
R30393 CS_BIAS.n1557 CS_BIAS.n1556 161.3
R30394 CS_BIAS.n1555 CS_BIAS.n1521 161.3
R30395 CS_BIAS.n1554 CS_BIAS.n1553 161.3
R30396 CS_BIAS.n1552 CS_BIAS.n1522 161.3
R30397 CS_BIAS.n1550 CS_BIAS.n1549 161.3
R30398 CS_BIAS.n1548 CS_BIAS.n1523 161.3
R30399 CS_BIAS.n1547 CS_BIAS.n1546 161.3
R30400 CS_BIAS.n1545 CS_BIAS.n1524 161.3
R30401 CS_BIAS.n1544 CS_BIAS.n1543 161.3
R30402 CS_BIAS.n1542 CS_BIAS.n1525 161.3
R30403 CS_BIAS.n1541 CS_BIAS.n1540 161.3
R30404 CS_BIAS.n1539 CS_BIAS.n1526 161.3
R30405 CS_BIAS.n1538 CS_BIAS.n1537 161.3
R30406 CS_BIAS.n1536 CS_BIAS.n1527 161.3
R30407 CS_BIAS.n1535 CS_BIAS.n1534 161.3
R30408 CS_BIAS.n1533 CS_BIAS.n1528 161.3
R30409 CS_BIAS.n1532 CS_BIAS.n1531 161.3
R30410 CS_BIAS.n1486 CS_BIAS.n1326 161.3
R30411 CS_BIAS.n1485 CS_BIAS.n1484 161.3
R30412 CS_BIAS.n1483 CS_BIAS.n1327 161.3
R30413 CS_BIAS.n1482 CS_BIAS.n1481 161.3
R30414 CS_BIAS.n1480 CS_BIAS.n1328 161.3
R30415 CS_BIAS.n1479 CS_BIAS.n1478 161.3
R30416 CS_BIAS.n1477 CS_BIAS.n1329 161.3
R30417 CS_BIAS.n1476 CS_BIAS.n1475 161.3
R30418 CS_BIAS.n1474 CS_BIAS.n1330 161.3
R30419 CS_BIAS.n1473 CS_BIAS.n1472 161.3
R30420 CS_BIAS.n1471 CS_BIAS.n1331 161.3
R30421 CS_BIAS.n1470 CS_BIAS.n1469 161.3
R30422 CS_BIAS.n1468 CS_BIAS.n1332 161.3
R30423 CS_BIAS.n1466 CS_BIAS.n1465 161.3
R30424 CS_BIAS.n1464 CS_BIAS.n1333 161.3
R30425 CS_BIAS.n1463 CS_BIAS.n1462 161.3
R30426 CS_BIAS.n1461 CS_BIAS.n1334 161.3
R30427 CS_BIAS.n1460 CS_BIAS.n1459 161.3
R30428 CS_BIAS.n1458 CS_BIAS.n1335 161.3
R30429 CS_BIAS.n1457 CS_BIAS.n1456 161.3
R30430 CS_BIAS.n1455 CS_BIAS.n1336 161.3
R30431 CS_BIAS.n1454 CS_BIAS.n1453 161.3
R30432 CS_BIAS.n1452 CS_BIAS.n1337 161.3
R30433 CS_BIAS.n1451 CS_BIAS.n1450 161.3
R30434 CS_BIAS.n1449 CS_BIAS.n1338 161.3
R30435 CS_BIAS.n1448 CS_BIAS.n1447 161.3
R30436 CS_BIAS.n1446 CS_BIAS.n1445 161.3
R30437 CS_BIAS.n1444 CS_BIAS.n1340 161.3
R30438 CS_BIAS.n1443 CS_BIAS.n1442 161.3
R30439 CS_BIAS.n1441 CS_BIAS.n1341 161.3
R30440 CS_BIAS.n1440 CS_BIAS.n1439 161.3
R30441 CS_BIAS.n1438 CS_BIAS.n1342 161.3
R30442 CS_BIAS.n1437 CS_BIAS.n1436 161.3
R30443 CS_BIAS.n1435 CS_BIAS.n1343 161.3
R30444 CS_BIAS.n1434 CS_BIAS.n1433 161.3
R30445 CS_BIAS.n1432 CS_BIAS.n1344 161.3
R30446 CS_BIAS.n1431 CS_BIAS.n1430 161.3
R30447 CS_BIAS.n1429 CS_BIAS.n1345 161.3
R30448 CS_BIAS.n1428 CS_BIAS.n1427 161.3
R30449 CS_BIAS.n1425 CS_BIAS.n1346 161.3
R30450 CS_BIAS.n1424 CS_BIAS.n1423 161.3
R30451 CS_BIAS.n1422 CS_BIAS.n1347 161.3
R30452 CS_BIAS.n1421 CS_BIAS.n1420 161.3
R30453 CS_BIAS.n1419 CS_BIAS.n1348 161.3
R30454 CS_BIAS.n1418 CS_BIAS.n1417 161.3
R30455 CS_BIAS.n1416 CS_BIAS.n1349 161.3
R30456 CS_BIAS.n1415 CS_BIAS.n1414 161.3
R30457 CS_BIAS.n1413 CS_BIAS.n1350 161.3
R30458 CS_BIAS.n1412 CS_BIAS.n1411 161.3
R30459 CS_BIAS.n1410 CS_BIAS.n1351 161.3
R30460 CS_BIAS.n1409 CS_BIAS.n1408 161.3
R30461 CS_BIAS.n1406 CS_BIAS.n1352 161.3
R30462 CS_BIAS.n1405 CS_BIAS.n1404 161.3
R30463 CS_BIAS.n1403 CS_BIAS.n1353 161.3
R30464 CS_BIAS.n1402 CS_BIAS.n1401 161.3
R30465 CS_BIAS.n1400 CS_BIAS.n1354 161.3
R30466 CS_BIAS.n1399 CS_BIAS.n1398 161.3
R30467 CS_BIAS.n1397 CS_BIAS.n1355 161.3
R30468 CS_BIAS.n1396 CS_BIAS.n1395 161.3
R30469 CS_BIAS.n1394 CS_BIAS.n1356 161.3
R30470 CS_BIAS.n1393 CS_BIAS.n1392 161.3
R30471 CS_BIAS.n1391 CS_BIAS.n1357 161.3
R30472 CS_BIAS.n1390 CS_BIAS.n1389 161.3
R30473 CS_BIAS.n1388 CS_BIAS.n1358 161.3
R30474 CS_BIAS.n1386 CS_BIAS.n1385 161.3
R30475 CS_BIAS.n1384 CS_BIAS.n1359 161.3
R30476 CS_BIAS.n1383 CS_BIAS.n1382 161.3
R30477 CS_BIAS.n1381 CS_BIAS.n1360 161.3
R30478 CS_BIAS.n1380 CS_BIAS.n1379 161.3
R30479 CS_BIAS.n1378 CS_BIAS.n1361 161.3
R30480 CS_BIAS.n1377 CS_BIAS.n1376 161.3
R30481 CS_BIAS.n1375 CS_BIAS.n1362 161.3
R30482 CS_BIAS.n1374 CS_BIAS.n1373 161.3
R30483 CS_BIAS.n1372 CS_BIAS.n1363 161.3
R30484 CS_BIAS.n1371 CS_BIAS.n1370 161.3
R30485 CS_BIAS.n1369 CS_BIAS.n1364 161.3
R30486 CS_BIAS.n1368 CS_BIAS.n1367 161.3
R30487 CS_BIAS.n1322 CS_BIAS.n1162 161.3
R30488 CS_BIAS.n1321 CS_BIAS.n1320 161.3
R30489 CS_BIAS.n1319 CS_BIAS.n1163 161.3
R30490 CS_BIAS.n1318 CS_BIAS.n1317 161.3
R30491 CS_BIAS.n1316 CS_BIAS.n1164 161.3
R30492 CS_BIAS.n1315 CS_BIAS.n1314 161.3
R30493 CS_BIAS.n1313 CS_BIAS.n1165 161.3
R30494 CS_BIAS.n1312 CS_BIAS.n1311 161.3
R30495 CS_BIAS.n1310 CS_BIAS.n1166 161.3
R30496 CS_BIAS.n1309 CS_BIAS.n1308 161.3
R30497 CS_BIAS.n1307 CS_BIAS.n1167 161.3
R30498 CS_BIAS.n1306 CS_BIAS.n1305 161.3
R30499 CS_BIAS.n1304 CS_BIAS.n1168 161.3
R30500 CS_BIAS.n1302 CS_BIAS.n1301 161.3
R30501 CS_BIAS.n1300 CS_BIAS.n1169 161.3
R30502 CS_BIAS.n1299 CS_BIAS.n1298 161.3
R30503 CS_BIAS.n1297 CS_BIAS.n1170 161.3
R30504 CS_BIAS.n1296 CS_BIAS.n1295 161.3
R30505 CS_BIAS.n1294 CS_BIAS.n1171 161.3
R30506 CS_BIAS.n1293 CS_BIAS.n1292 161.3
R30507 CS_BIAS.n1291 CS_BIAS.n1172 161.3
R30508 CS_BIAS.n1290 CS_BIAS.n1289 161.3
R30509 CS_BIAS.n1288 CS_BIAS.n1173 161.3
R30510 CS_BIAS.n1287 CS_BIAS.n1286 161.3
R30511 CS_BIAS.n1285 CS_BIAS.n1174 161.3
R30512 CS_BIAS.n1284 CS_BIAS.n1283 161.3
R30513 CS_BIAS.n1282 CS_BIAS.n1281 161.3
R30514 CS_BIAS.n1280 CS_BIAS.n1176 161.3
R30515 CS_BIAS.n1279 CS_BIAS.n1278 161.3
R30516 CS_BIAS.n1277 CS_BIAS.n1177 161.3
R30517 CS_BIAS.n1276 CS_BIAS.n1275 161.3
R30518 CS_BIAS.n1274 CS_BIAS.n1178 161.3
R30519 CS_BIAS.n1273 CS_BIAS.n1272 161.3
R30520 CS_BIAS.n1271 CS_BIAS.n1179 161.3
R30521 CS_BIAS.n1270 CS_BIAS.n1269 161.3
R30522 CS_BIAS.n1268 CS_BIAS.n1180 161.3
R30523 CS_BIAS.n1267 CS_BIAS.n1266 161.3
R30524 CS_BIAS.n1265 CS_BIAS.n1181 161.3
R30525 CS_BIAS.n1264 CS_BIAS.n1263 161.3
R30526 CS_BIAS.n1261 CS_BIAS.n1182 161.3
R30527 CS_BIAS.n1260 CS_BIAS.n1259 161.3
R30528 CS_BIAS.n1258 CS_BIAS.n1183 161.3
R30529 CS_BIAS.n1257 CS_BIAS.n1256 161.3
R30530 CS_BIAS.n1255 CS_BIAS.n1184 161.3
R30531 CS_BIAS.n1254 CS_BIAS.n1253 161.3
R30532 CS_BIAS.n1252 CS_BIAS.n1185 161.3
R30533 CS_BIAS.n1251 CS_BIAS.n1250 161.3
R30534 CS_BIAS.n1249 CS_BIAS.n1186 161.3
R30535 CS_BIAS.n1248 CS_BIAS.n1247 161.3
R30536 CS_BIAS.n1246 CS_BIAS.n1187 161.3
R30537 CS_BIAS.n1245 CS_BIAS.n1244 161.3
R30538 CS_BIAS.n1242 CS_BIAS.n1188 161.3
R30539 CS_BIAS.n1241 CS_BIAS.n1240 161.3
R30540 CS_BIAS.n1239 CS_BIAS.n1189 161.3
R30541 CS_BIAS.n1238 CS_BIAS.n1237 161.3
R30542 CS_BIAS.n1236 CS_BIAS.n1190 161.3
R30543 CS_BIAS.n1235 CS_BIAS.n1234 161.3
R30544 CS_BIAS.n1233 CS_BIAS.n1191 161.3
R30545 CS_BIAS.n1232 CS_BIAS.n1231 161.3
R30546 CS_BIAS.n1230 CS_BIAS.n1192 161.3
R30547 CS_BIAS.n1229 CS_BIAS.n1228 161.3
R30548 CS_BIAS.n1227 CS_BIAS.n1193 161.3
R30549 CS_BIAS.n1226 CS_BIAS.n1225 161.3
R30550 CS_BIAS.n1224 CS_BIAS.n1194 161.3
R30551 CS_BIAS.n1222 CS_BIAS.n1221 161.3
R30552 CS_BIAS.n1220 CS_BIAS.n1195 161.3
R30553 CS_BIAS.n1219 CS_BIAS.n1218 161.3
R30554 CS_BIAS.n1217 CS_BIAS.n1196 161.3
R30555 CS_BIAS.n1216 CS_BIAS.n1215 161.3
R30556 CS_BIAS.n1214 CS_BIAS.n1197 161.3
R30557 CS_BIAS.n1213 CS_BIAS.n1212 161.3
R30558 CS_BIAS.n1211 CS_BIAS.n1198 161.3
R30559 CS_BIAS.n1210 CS_BIAS.n1209 161.3
R30560 CS_BIAS.n1208 CS_BIAS.n1199 161.3
R30561 CS_BIAS.n1207 CS_BIAS.n1206 161.3
R30562 CS_BIAS.n1205 CS_BIAS.n1200 161.3
R30563 CS_BIAS.n1204 CS_BIAS.n1203 161.3
R30564 CS_BIAS.n1081 CS_BIAS.n921 161.3
R30565 CS_BIAS.n1080 CS_BIAS.n1079 161.3
R30566 CS_BIAS.n1078 CS_BIAS.n922 161.3
R30567 CS_BIAS.n1077 CS_BIAS.n1076 161.3
R30568 CS_BIAS.n1075 CS_BIAS.n923 161.3
R30569 CS_BIAS.n1074 CS_BIAS.n1073 161.3
R30570 CS_BIAS.n1072 CS_BIAS.n924 161.3
R30571 CS_BIAS.n1071 CS_BIAS.n1070 161.3
R30572 CS_BIAS.n1069 CS_BIAS.n925 161.3
R30573 CS_BIAS.n1068 CS_BIAS.n1067 161.3
R30574 CS_BIAS.n1066 CS_BIAS.n926 161.3
R30575 CS_BIAS.n1065 CS_BIAS.n1064 161.3
R30576 CS_BIAS.n1063 CS_BIAS.n927 161.3
R30577 CS_BIAS.n1061 CS_BIAS.n1060 161.3
R30578 CS_BIAS.n1059 CS_BIAS.n928 161.3
R30579 CS_BIAS.n1058 CS_BIAS.n1057 161.3
R30580 CS_BIAS.n1056 CS_BIAS.n929 161.3
R30581 CS_BIAS.n1055 CS_BIAS.n1054 161.3
R30582 CS_BIAS.n1053 CS_BIAS.n930 161.3
R30583 CS_BIAS.n1052 CS_BIAS.n1051 161.3
R30584 CS_BIAS.n1050 CS_BIAS.n931 161.3
R30585 CS_BIAS.n1049 CS_BIAS.n1048 161.3
R30586 CS_BIAS.n1047 CS_BIAS.n932 161.3
R30587 CS_BIAS.n1046 CS_BIAS.n1045 161.3
R30588 CS_BIAS.n1044 CS_BIAS.n933 161.3
R30589 CS_BIAS.n1043 CS_BIAS.n1042 161.3
R30590 CS_BIAS.n1041 CS_BIAS.n1040 161.3
R30591 CS_BIAS.n1039 CS_BIAS.n935 161.3
R30592 CS_BIAS.n1038 CS_BIAS.n1037 161.3
R30593 CS_BIAS.n1036 CS_BIAS.n936 161.3
R30594 CS_BIAS.n1035 CS_BIAS.n1034 161.3
R30595 CS_BIAS.n1033 CS_BIAS.n937 161.3
R30596 CS_BIAS.n1032 CS_BIAS.n1031 161.3
R30597 CS_BIAS.n1030 CS_BIAS.n938 161.3
R30598 CS_BIAS.n1029 CS_BIAS.n1028 161.3
R30599 CS_BIAS.n1027 CS_BIAS.n939 161.3
R30600 CS_BIAS.n1026 CS_BIAS.n1025 161.3
R30601 CS_BIAS.n1024 CS_BIAS.n940 161.3
R30602 CS_BIAS.n1023 CS_BIAS.n1022 161.3
R30603 CS_BIAS.n1020 CS_BIAS.n941 161.3
R30604 CS_BIAS.n1019 CS_BIAS.n1018 161.3
R30605 CS_BIAS.n1017 CS_BIAS.n942 161.3
R30606 CS_BIAS.n1016 CS_BIAS.n1015 161.3
R30607 CS_BIAS.n1014 CS_BIAS.n943 161.3
R30608 CS_BIAS.n1013 CS_BIAS.n1012 161.3
R30609 CS_BIAS.n1011 CS_BIAS.n944 161.3
R30610 CS_BIAS.n1010 CS_BIAS.n1009 161.3
R30611 CS_BIAS.n1008 CS_BIAS.n945 161.3
R30612 CS_BIAS.n1007 CS_BIAS.n1006 161.3
R30613 CS_BIAS.n1005 CS_BIAS.n946 161.3
R30614 CS_BIAS.n1004 CS_BIAS.n1003 161.3
R30615 CS_BIAS.n1001 CS_BIAS.n947 161.3
R30616 CS_BIAS.n1000 CS_BIAS.n999 161.3
R30617 CS_BIAS.n998 CS_BIAS.n948 161.3
R30618 CS_BIAS.n997 CS_BIAS.n996 161.3
R30619 CS_BIAS.n995 CS_BIAS.n949 161.3
R30620 CS_BIAS.n994 CS_BIAS.n993 161.3
R30621 CS_BIAS.n992 CS_BIAS.n950 161.3
R30622 CS_BIAS.n991 CS_BIAS.n990 161.3
R30623 CS_BIAS.n989 CS_BIAS.n951 161.3
R30624 CS_BIAS.n988 CS_BIAS.n987 161.3
R30625 CS_BIAS.n986 CS_BIAS.n952 161.3
R30626 CS_BIAS.n985 CS_BIAS.n984 161.3
R30627 CS_BIAS.n983 CS_BIAS.n953 161.3
R30628 CS_BIAS.n981 CS_BIAS.n980 161.3
R30629 CS_BIAS.n979 CS_BIAS.n954 161.3
R30630 CS_BIAS.n978 CS_BIAS.n977 161.3
R30631 CS_BIAS.n976 CS_BIAS.n955 161.3
R30632 CS_BIAS.n975 CS_BIAS.n974 161.3
R30633 CS_BIAS.n973 CS_BIAS.n956 161.3
R30634 CS_BIAS.n972 CS_BIAS.n971 161.3
R30635 CS_BIAS.n970 CS_BIAS.n957 161.3
R30636 CS_BIAS.n969 CS_BIAS.n968 161.3
R30637 CS_BIAS.n967 CS_BIAS.n958 161.3
R30638 CS_BIAS.n966 CS_BIAS.n965 161.3
R30639 CS_BIAS.n964 CS_BIAS.n959 161.3
R30640 CS_BIAS.n963 CS_BIAS.n962 161.3
R30641 CS_BIAS.n917 CS_BIAS.n850 161.3
R30642 CS_BIAS.n916 CS_BIAS.n915 161.3
R30643 CS_BIAS.n914 CS_BIAS.n851 161.3
R30644 CS_BIAS.n913 CS_BIAS.n912 161.3
R30645 CS_BIAS.n911 CS_BIAS.n852 161.3
R30646 CS_BIAS.n910 CS_BIAS.n909 161.3
R30647 CS_BIAS.n907 CS_BIAS.n853 161.3
R30648 CS_BIAS.n906 CS_BIAS.n905 161.3
R30649 CS_BIAS.n904 CS_BIAS.n854 161.3
R30650 CS_BIAS.n903 CS_BIAS.n902 161.3
R30651 CS_BIAS.n901 CS_BIAS.n855 161.3
R30652 CS_BIAS.n900 CS_BIAS.n899 161.3
R30653 CS_BIAS.n898 CS_BIAS.n856 161.3
R30654 CS_BIAS.n897 CS_BIAS.n896 161.3
R30655 CS_BIAS.n895 CS_BIAS.n857 161.3
R30656 CS_BIAS.n894 CS_BIAS.n893 161.3
R30657 CS_BIAS.n892 CS_BIAS.n858 161.3
R30658 CS_BIAS.n891 CS_BIAS.n890 161.3
R30659 CS_BIAS.n889 CS_BIAS.n859 161.3
R30660 CS_BIAS.n887 CS_BIAS.n886 161.3
R30661 CS_BIAS.n885 CS_BIAS.n860 161.3
R30662 CS_BIAS.n884 CS_BIAS.n883 161.3
R30663 CS_BIAS.n882 CS_BIAS.n861 161.3
R30664 CS_BIAS.n881 CS_BIAS.n880 161.3
R30665 CS_BIAS.n879 CS_BIAS.n862 161.3
R30666 CS_BIAS.n878 CS_BIAS.n877 161.3
R30667 CS_BIAS.n876 CS_BIAS.n863 161.3
R30668 CS_BIAS.n875 CS_BIAS.n874 161.3
R30669 CS_BIAS.n873 CS_BIAS.n864 161.3
R30670 CS_BIAS.n872 CS_BIAS.n871 161.3
R30671 CS_BIAS.n870 CS_BIAS.n865 161.3
R30672 CS_BIAS.n869 CS_BIAS.n868 161.3
R30673 CS_BIAS.n1159 CS_BIAS.n827 161.3
R30674 CS_BIAS.n1158 CS_BIAS.n1157 161.3
R30675 CS_BIAS.n1156 CS_BIAS.n828 161.3
R30676 CS_BIAS.n1155 CS_BIAS.n1154 161.3
R30677 CS_BIAS.n1153 CS_BIAS.n829 161.3
R30678 CS_BIAS.n1152 CS_BIAS.n1151 161.3
R30679 CS_BIAS.n1150 CS_BIAS.n830 161.3
R30680 CS_BIAS.n1149 CS_BIAS.n1148 161.3
R30681 CS_BIAS.n1147 CS_BIAS.n831 161.3
R30682 CS_BIAS.n1146 CS_BIAS.n1145 161.3
R30683 CS_BIAS.n1144 CS_BIAS.n832 161.3
R30684 CS_BIAS.n1143 CS_BIAS.n1142 161.3
R30685 CS_BIAS.n1141 CS_BIAS.n833 161.3
R30686 CS_BIAS.n1139 CS_BIAS.n1138 161.3
R30687 CS_BIAS.n1137 CS_BIAS.n834 161.3
R30688 CS_BIAS.n1136 CS_BIAS.n1135 161.3
R30689 CS_BIAS.n1134 CS_BIAS.n835 161.3
R30690 CS_BIAS.n1133 CS_BIAS.n1132 161.3
R30691 CS_BIAS.n1131 CS_BIAS.n836 161.3
R30692 CS_BIAS.n1130 CS_BIAS.n1129 161.3
R30693 CS_BIAS.n1128 CS_BIAS.n837 161.3
R30694 CS_BIAS.n1127 CS_BIAS.n1126 161.3
R30695 CS_BIAS.n1125 CS_BIAS.n838 161.3
R30696 CS_BIAS.n1124 CS_BIAS.n1123 161.3
R30697 CS_BIAS.n1122 CS_BIAS.n839 161.3
R30698 CS_BIAS.n1121 CS_BIAS.n1120 161.3
R30699 CS_BIAS.n1119 CS_BIAS.n1118 161.3
R30700 CS_BIAS.n1117 CS_BIAS.n841 161.3
R30701 CS_BIAS.n1116 CS_BIAS.n1115 161.3
R30702 CS_BIAS.n1114 CS_BIAS.n842 161.3
R30703 CS_BIAS.n1113 CS_BIAS.n1112 161.3
R30704 CS_BIAS.n1111 CS_BIAS.n843 161.3
R30705 CS_BIAS.n1110 CS_BIAS.n1109 161.3
R30706 CS_BIAS.n1108 CS_BIAS.n844 161.3
R30707 CS_BIAS.n1107 CS_BIAS.n1106 161.3
R30708 CS_BIAS.n1105 CS_BIAS.n845 161.3
R30709 CS_BIAS.n1104 CS_BIAS.n1103 161.3
R30710 CS_BIAS.n1102 CS_BIAS.n846 161.3
R30711 CS_BIAS.n1101 CS_BIAS.n1100 161.3
R30712 CS_BIAS.n1098 CS_BIAS.n847 161.3
R30713 CS_BIAS.n1097 CS_BIAS.n1096 161.3
R30714 CS_BIAS.n1095 CS_BIAS.n848 161.3
R30715 CS_BIAS.n1094 CS_BIAS.n1093 161.3
R30716 CS_BIAS.n1092 CS_BIAS.n849 161.3
R30717 CS_BIAS.n1091 CS_BIAS.n1090 161.3
R30718 CS_BIAS.n713 CS_BIAS.n712 73.0308
R30719 CS_BIAS.n732 CS_BIAS.n692 73.0308
R30720 CS_BIAS.n755 CS_BIAS.n686 73.0308
R30721 CS_BIAS.n775 CS_BIAS.n774 73.0308
R30722 CS_BIAS.n793 CS_BIAS.n672 73.0308
R30723 CS_BIAS.n816 CS_BIAS.n666 73.0308
R30724 CS_BIAS.n652 CS_BIAS.n502 73.0308
R30725 CS_BIAS.n629 CS_BIAS.n508 73.0308
R30726 CS_BIAS.n611 CS_BIAS.n610 73.0308
R30727 CS_BIAS.n591 CS_BIAS.n522 73.0308
R30728 CS_BIAS.n568 CS_BIAS.n528 73.0308
R30729 CS_BIAS.n549 CS_BIAS.n548 73.0308
R30730 CS_BIAS.n488 CS_BIAS.n338 73.0308
R30731 CS_BIAS.n465 CS_BIAS.n344 73.0308
R30732 CS_BIAS.n447 CS_BIAS.n446 73.0308
R30733 CS_BIAS.n427 CS_BIAS.n358 73.0308
R30734 CS_BIAS.n404 CS_BIAS.n364 73.0308
R30735 CS_BIAS.n385 CS_BIAS.n384 73.0308
R30736 CS_BIAS.n244 CS_BIAS.n94 73.0308
R30737 CS_BIAS.n221 CS_BIAS.n100 73.0308
R30738 CS_BIAS.n203 CS_BIAS.n202 73.0308
R30739 CS_BIAS.n183 CS_BIAS.n114 73.0308
R30740 CS_BIAS.n160 CS_BIAS.n120 73.0308
R30741 CS_BIAS.n141 CS_BIAS.n140 73.0308
R30742 CS_BIAS.n325 CS_BIAS.n3 73.0308
R30743 CS_BIAS.n302 CS_BIAS.n9 73.0308
R30744 CS_BIAS.n284 CS_BIAS.n283 73.0308
R30745 CS_BIAS.n264 CS_BIAS.n23 73.0308
R30746 CS_BIAS.n69 CS_BIAS.n29 73.0308
R30747 CS_BIAS.n50 CS_BIAS.n49 73.0308
R30748 CS_BIAS.n1540 CS_BIAS.n1539 73.0308
R30749 CS_BIAS.n1559 CS_BIAS.n1519 73.0308
R30750 CS_BIAS.n1582 CS_BIAS.n1513 73.0308
R30751 CS_BIAS.n1602 CS_BIAS.n1601 73.0308
R30752 CS_BIAS.n1620 CS_BIAS.n1499 73.0308
R30753 CS_BIAS.n1643 CS_BIAS.n1493 73.0308
R30754 CS_BIAS.n1376 CS_BIAS.n1375 73.0308
R30755 CS_BIAS.n1395 CS_BIAS.n1355 73.0308
R30756 CS_BIAS.n1418 CS_BIAS.n1349 73.0308
R30757 CS_BIAS.n1438 CS_BIAS.n1437 73.0308
R30758 CS_BIAS.n1456 CS_BIAS.n1335 73.0308
R30759 CS_BIAS.n1479 CS_BIAS.n1329 73.0308
R30760 CS_BIAS.n1212 CS_BIAS.n1211 73.0308
R30761 CS_BIAS.n1231 CS_BIAS.n1191 73.0308
R30762 CS_BIAS.n1254 CS_BIAS.n1185 73.0308
R30763 CS_BIAS.n1274 CS_BIAS.n1273 73.0308
R30764 CS_BIAS.n1292 CS_BIAS.n1171 73.0308
R30765 CS_BIAS.n1315 CS_BIAS.n1165 73.0308
R30766 CS_BIAS.n971 CS_BIAS.n970 73.0308
R30767 CS_BIAS.n990 CS_BIAS.n950 73.0308
R30768 CS_BIAS.n1013 CS_BIAS.n944 73.0308
R30769 CS_BIAS.n1033 CS_BIAS.n1032 73.0308
R30770 CS_BIAS.n1051 CS_BIAS.n930 73.0308
R30771 CS_BIAS.n1074 CS_BIAS.n924 73.0308
R30772 CS_BIAS.n1152 CS_BIAS.n830 73.0308
R30773 CS_BIAS.n1129 CS_BIAS.n836 73.0308
R30774 CS_BIAS.n1111 CS_BIAS.n1110 73.0308
R30775 CS_BIAS.n877 CS_BIAS.n876 73.0308
R30776 CS_BIAS.n896 CS_BIAS.n856 73.0308
R30777 CS_BIAS.n1091 CS_BIAS.n850 73.0308
R30778 CS_BIAS.n260 CS_BIAS.n258 72.7259
R30779 CS_BIAS.n920 CS_BIAS.n918 72.7259
R30780 CS_BIAS.n260 CS_BIAS.n259 70.8609
R30781 CS_BIAS.n257 CS_BIAS.n256 70.8609
R30782 CS_BIAS.n255 CS_BIAS.n254 70.8609
R30783 CS_BIAS.n1085 CS_BIAS.n1084 70.8609
R30784 CS_BIAS.n1087 CS_BIAS.n1086 70.8609
R30785 CS_BIAS.n920 CS_BIAS.n919 70.8609
R30786 CS_BIAS.n825 CS_BIAS.n824 54.5572
R30787 CS_BIAS.n661 CS_BIAS.n660 54.5572
R30788 CS_BIAS.n497 CS_BIAS.n496 54.5572
R30789 CS_BIAS.n253 CS_BIAS.n252 54.5572
R30790 CS_BIAS.n334 CS_BIAS.n333 54.5572
R30791 CS_BIAS.n1652 CS_BIAS.n1651 54.5572
R30792 CS_BIAS.n1488 CS_BIAS.n1487 54.5572
R30793 CS_BIAS.n1324 CS_BIAS.n1323 54.5572
R30794 CS_BIAS.n1083 CS_BIAS.n1082 54.5572
R30795 CS_BIAS.n1161 CS_BIAS.n1160 54.5572
R30796 CS_BIAS.n703 CS_BIAS.n702 52.78
R30797 CS_BIAS.n539 CS_BIAS.n538 52.78
R30798 CS_BIAS.n375 CS_BIAS.n374 52.78
R30799 CS_BIAS.n131 CS_BIAS.n130 52.78
R30800 CS_BIAS.n40 CS_BIAS.n39 52.78
R30801 CS_BIAS.n1530 CS_BIAS.n1529 52.78
R30802 CS_BIAS.n1366 CS_BIAS.n1365 52.78
R30803 CS_BIAS.n1202 CS_BIAS.n1201 52.78
R30804 CS_BIAS.n961 CS_BIAS.n960 52.78
R30805 CS_BIAS.n867 CS_BIAS.n866 52.78
R30806 CS_BIAS.n703 CS_BIAS.t51 48.5512
R30807 CS_BIAS.n1530 CS_BIAS.t64 48.5512
R30808 CS_BIAS.n1366 CS_BIAS.t32 48.5512
R30809 CS_BIAS.n1202 CS_BIAS.t65 48.5512
R30810 CS_BIAS.n961 CS_BIAS.t22 48.5512
R30811 CS_BIAS.n867 CS_BIAS.t77 48.5512
R30812 CS_BIAS.n539 CS_BIAS.t81 48.5508
R30813 CS_BIAS.n375 CS_BIAS.t52 48.5508
R30814 CS_BIAS.n131 CS_BIAS.t6 48.5508
R30815 CS_BIAS.n40 CS_BIAS.t94 48.5508
R30816 CS_BIAS.n812 CS_BIAS.n666 35.1514
R30817 CS_BIAS.n648 CS_BIAS.n502 35.1514
R30818 CS_BIAS.n484 CS_BIAS.n338 35.1514
R30819 CS_BIAS.n240 CS_BIAS.n94 35.1514
R30820 CS_BIAS.n321 CS_BIAS.n3 35.1514
R30821 CS_BIAS.n1639 CS_BIAS.n1493 35.1514
R30822 CS_BIAS.n1475 CS_BIAS.n1329 35.1514
R30823 CS_BIAS.n1311 CS_BIAS.n1165 35.1514
R30824 CS_BIAS.n1070 CS_BIAS.n924 35.1514
R30825 CS_BIAS.n1148 CS_BIAS.n830 35.1514
R30826 CS_BIAS.n713 CS_BIAS.n698 34.1802
R30827 CS_BIAS.n793 CS_BIAS.n792 34.1802
R30828 CS_BIAS.n629 CS_BIAS.n628 34.1802
R30829 CS_BIAS.n549 CS_BIAS.n534 34.1802
R30830 CS_BIAS.n465 CS_BIAS.n464 34.1802
R30831 CS_BIAS.n385 CS_BIAS.n370 34.1802
R30832 CS_BIAS.n221 CS_BIAS.n220 34.1802
R30833 CS_BIAS.n141 CS_BIAS.n126 34.1802
R30834 CS_BIAS.n302 CS_BIAS.n301 34.1802
R30835 CS_BIAS.n50 CS_BIAS.n35 34.1802
R30836 CS_BIAS.n1540 CS_BIAS.n1525 34.1802
R30837 CS_BIAS.n1620 CS_BIAS.n1619 34.1802
R30838 CS_BIAS.n1376 CS_BIAS.n1361 34.1802
R30839 CS_BIAS.n1456 CS_BIAS.n1455 34.1802
R30840 CS_BIAS.n1212 CS_BIAS.n1197 34.1802
R30841 CS_BIAS.n1292 CS_BIAS.n1291 34.1802
R30842 CS_BIAS.n971 CS_BIAS.n956 34.1802
R30843 CS_BIAS.n1051 CS_BIAS.n1050 34.1802
R30844 CS_BIAS.n1129 CS_BIAS.n1128 34.1802
R30845 CS_BIAS.n877 CS_BIAS.n862 34.1802
R30846 CS_BIAS.n736 CS_BIAS.n692 33.2089
R30847 CS_BIAS.n774 CS_BIAS.n680 33.2089
R30848 CS_BIAS.n610 CS_BIAS.n516 33.2089
R30849 CS_BIAS.n572 CS_BIAS.n528 33.2089
R30850 CS_BIAS.n446 CS_BIAS.n352 33.2089
R30851 CS_BIAS.n408 CS_BIAS.n364 33.2089
R30852 CS_BIAS.n202 CS_BIAS.n108 33.2089
R30853 CS_BIAS.n164 CS_BIAS.n120 33.2089
R30854 CS_BIAS.n283 CS_BIAS.n17 33.2089
R30855 CS_BIAS.n73 CS_BIAS.n29 33.2089
R30856 CS_BIAS.n1563 CS_BIAS.n1519 33.2089
R30857 CS_BIAS.n1601 CS_BIAS.n1507 33.2089
R30858 CS_BIAS.n1399 CS_BIAS.n1355 33.2089
R30859 CS_BIAS.n1437 CS_BIAS.n1343 33.2089
R30860 CS_BIAS.n1235 CS_BIAS.n1191 33.2089
R30861 CS_BIAS.n1273 CS_BIAS.n1179 33.2089
R30862 CS_BIAS.n994 CS_BIAS.n950 33.2089
R30863 CS_BIAS.n1032 CS_BIAS.n938 33.2089
R30864 CS_BIAS.n1110 CS_BIAS.n844 33.2089
R30865 CS_BIAS.n900 CS_BIAS.n856 33.2089
R30866 CS_BIAS.n751 CS_BIAS.n686 32.2376
R30867 CS_BIAS.n756 CS_BIAS.n755 32.2376
R30868 CS_BIAS.n592 CS_BIAS.n591 32.2376
R30869 CS_BIAS.n587 CS_BIAS.n522 32.2376
R30870 CS_BIAS.n428 CS_BIAS.n427 32.2376
R30871 CS_BIAS.n423 CS_BIAS.n358 32.2376
R30872 CS_BIAS.n184 CS_BIAS.n183 32.2376
R30873 CS_BIAS.n179 CS_BIAS.n114 32.2376
R30874 CS_BIAS.n265 CS_BIAS.n264 32.2376
R30875 CS_BIAS.n88 CS_BIAS.n23 32.2376
R30876 CS_BIAS.n1578 CS_BIAS.n1513 32.2376
R30877 CS_BIAS.n1583 CS_BIAS.n1582 32.2376
R30878 CS_BIAS.n1414 CS_BIAS.n1349 32.2376
R30879 CS_BIAS.n1419 CS_BIAS.n1418 32.2376
R30880 CS_BIAS.n1250 CS_BIAS.n1185 32.2376
R30881 CS_BIAS.n1255 CS_BIAS.n1254 32.2376
R30882 CS_BIAS.n1009 CS_BIAS.n944 32.2376
R30883 CS_BIAS.n1014 CS_BIAS.n1013 32.2376
R30884 CS_BIAS.n1092 CS_BIAS.n1091 32.2376
R30885 CS_BIAS.n915 CS_BIAS.n850 32.2376
R30886 CS_BIAS.n732 CS_BIAS.n731 31.2664
R30887 CS_BIAS.n776 CS_BIAS.n775 31.2664
R30888 CS_BIAS.n612 CS_BIAS.n611 31.2664
R30889 CS_BIAS.n568 CS_BIAS.n567 31.2664
R30890 CS_BIAS.n448 CS_BIAS.n447 31.2664
R30891 CS_BIAS.n404 CS_BIAS.n403 31.2664
R30892 CS_BIAS.n204 CS_BIAS.n203 31.2664
R30893 CS_BIAS.n160 CS_BIAS.n159 31.2664
R30894 CS_BIAS.n285 CS_BIAS.n284 31.2664
R30895 CS_BIAS.n69 CS_BIAS.n68 31.2664
R30896 CS_BIAS.n1559 CS_BIAS.n1558 31.2664
R30897 CS_BIAS.n1603 CS_BIAS.n1602 31.2664
R30898 CS_BIAS.n1395 CS_BIAS.n1394 31.2664
R30899 CS_BIAS.n1439 CS_BIAS.n1438 31.2664
R30900 CS_BIAS.n1231 CS_BIAS.n1230 31.2664
R30901 CS_BIAS.n1275 CS_BIAS.n1274 31.2664
R30902 CS_BIAS.n990 CS_BIAS.n989 31.2664
R30903 CS_BIAS.n1034 CS_BIAS.n1033 31.2664
R30904 CS_BIAS.n1112 CS_BIAS.n1111 31.2664
R30905 CS_BIAS.n896 CS_BIAS.n895 31.2664
R30906 CS_BIAS.n712 CS_BIAS.n711 30.2951
R30907 CS_BIAS.n797 CS_BIAS.n672 30.2951
R30908 CS_BIAS.n633 CS_BIAS.n508 30.2951
R30909 CS_BIAS.n548 CS_BIAS.n547 30.2951
R30910 CS_BIAS.n469 CS_BIAS.n344 30.2951
R30911 CS_BIAS.n384 CS_BIAS.n383 30.2951
R30912 CS_BIAS.n225 CS_BIAS.n100 30.2951
R30913 CS_BIAS.n140 CS_BIAS.n139 30.2951
R30914 CS_BIAS.n306 CS_BIAS.n9 30.2951
R30915 CS_BIAS.n49 CS_BIAS.n48 30.2951
R30916 CS_BIAS.n1539 CS_BIAS.n1538 30.2951
R30917 CS_BIAS.n1624 CS_BIAS.n1499 30.2951
R30918 CS_BIAS.n1375 CS_BIAS.n1374 30.2951
R30919 CS_BIAS.n1460 CS_BIAS.n1335 30.2951
R30920 CS_BIAS.n1211 CS_BIAS.n1210 30.2951
R30921 CS_BIAS.n1296 CS_BIAS.n1171 30.2951
R30922 CS_BIAS.n970 CS_BIAS.n969 30.2951
R30923 CS_BIAS.n1055 CS_BIAS.n930 30.2951
R30924 CS_BIAS.n1133 CS_BIAS.n836 30.2951
R30925 CS_BIAS.n876 CS_BIAS.n875 30.2951
R30926 CS_BIAS.n817 CS_BIAS.n816 29.3238
R30927 CS_BIAS.n653 CS_BIAS.n652 29.3238
R30928 CS_BIAS.n489 CS_BIAS.n488 29.3238
R30929 CS_BIAS.n245 CS_BIAS.n244 29.3238
R30930 CS_BIAS.n326 CS_BIAS.n325 29.3238
R30931 CS_BIAS.n1644 CS_BIAS.n1643 29.3238
R30932 CS_BIAS.n1480 CS_BIAS.n1479 29.3238
R30933 CS_BIAS.n1316 CS_BIAS.n1315 29.3238
R30934 CS_BIAS.n1075 CS_BIAS.n1074 29.3238
R30935 CS_BIAS.n1153 CS_BIAS.n1152 29.3238
R30936 CS_BIAS.n711 CS_BIAS.n700 24.4675
R30937 CS_BIAS.n707 CS_BIAS.n700 24.4675
R30938 CS_BIAS.n707 CS_BIAS.n706 24.4675
R30939 CS_BIAS.n706 CS_BIAS.n705 24.4675
R30940 CS_BIAS.n731 CS_BIAS.n730 24.4675
R30941 CS_BIAS.n730 CS_BIAS.n694 24.4675
R30942 CS_BIAS.n726 CS_BIAS.n694 24.4675
R30943 CS_BIAS.n726 CS_BIAS.n725 24.4675
R30944 CS_BIAS.n723 CS_BIAS.n696 24.4675
R30945 CS_BIAS.n719 CS_BIAS.n696 24.4675
R30946 CS_BIAS.n719 CS_BIAS.n718 24.4675
R30947 CS_BIAS.n718 CS_BIAS.n717 24.4675
R30948 CS_BIAS.n717 CS_BIAS.n698 24.4675
R30949 CS_BIAS.n751 CS_BIAS.n750 24.4675
R30950 CS_BIAS.n750 CS_BIAS.n749 24.4675
R30951 CS_BIAS.n749 CS_BIAS.n688 24.4675
R30952 CS_BIAS.n745 CS_BIAS.n688 24.4675
R30953 CS_BIAS.n743 CS_BIAS.n742 24.4675
R30954 CS_BIAS.n742 CS_BIAS.n690 24.4675
R30955 CS_BIAS.n738 CS_BIAS.n690 24.4675
R30956 CS_BIAS.n738 CS_BIAS.n737 24.4675
R30957 CS_BIAS.n737 CS_BIAS.n736 24.4675
R30958 CS_BIAS.n770 CS_BIAS.n680 24.4675
R30959 CS_BIAS.n770 CS_BIAS.n769 24.4675
R30960 CS_BIAS.n769 CS_BIAS.n768 24.4675
R30961 CS_BIAS.n768 CS_BIAS.n682 24.4675
R30962 CS_BIAS.n764 CS_BIAS.n682 24.4675
R30963 CS_BIAS.n762 CS_BIAS.n761 24.4675
R30964 CS_BIAS.n761 CS_BIAS.n684 24.4675
R30965 CS_BIAS.n757 CS_BIAS.n684 24.4675
R30966 CS_BIAS.n757 CS_BIAS.n756 24.4675
R30967 CS_BIAS.n792 CS_BIAS.n791 24.4675
R30968 CS_BIAS.n791 CS_BIAS.n674 24.4675
R30969 CS_BIAS.n787 CS_BIAS.n674 24.4675
R30970 CS_BIAS.n787 CS_BIAS.n786 24.4675
R30971 CS_BIAS.n786 CS_BIAS.n785 24.4675
R30972 CS_BIAS.n782 CS_BIAS.n781 24.4675
R30973 CS_BIAS.n781 CS_BIAS.n780 24.4675
R30974 CS_BIAS.n780 CS_BIAS.n678 24.4675
R30975 CS_BIAS.n776 CS_BIAS.n678 24.4675
R30976 CS_BIAS.n812 CS_BIAS.n811 24.4675
R30977 CS_BIAS.n811 CS_BIAS.n810 24.4675
R30978 CS_BIAS.n810 CS_BIAS.n668 24.4675
R30979 CS_BIAS.n806 CS_BIAS.n668 24.4675
R30980 CS_BIAS.n806 CS_BIAS.n805 24.4675
R30981 CS_BIAS.n803 CS_BIAS.n670 24.4675
R30982 CS_BIAS.n799 CS_BIAS.n670 24.4675
R30983 CS_BIAS.n799 CS_BIAS.n798 24.4675
R30984 CS_BIAS.n798 CS_BIAS.n797 24.4675
R30985 CS_BIAS.n823 CS_BIAS.n822 24.4675
R30986 CS_BIAS.n822 CS_BIAS.n664 24.4675
R30987 CS_BIAS.n818 CS_BIAS.n664 24.4675
R30988 CS_BIAS.n818 CS_BIAS.n817 24.4675
R30989 CS_BIAS.n659 CS_BIAS.n658 24.4675
R30990 CS_BIAS.n658 CS_BIAS.n500 24.4675
R30991 CS_BIAS.n654 CS_BIAS.n500 24.4675
R30992 CS_BIAS.n654 CS_BIAS.n653 24.4675
R30993 CS_BIAS.n648 CS_BIAS.n647 24.4675
R30994 CS_BIAS.n647 CS_BIAS.n646 24.4675
R30995 CS_BIAS.n646 CS_BIAS.n504 24.4675
R30996 CS_BIAS.n642 CS_BIAS.n504 24.4675
R30997 CS_BIAS.n642 CS_BIAS.n641 24.4675
R30998 CS_BIAS.n639 CS_BIAS.n506 24.4675
R30999 CS_BIAS.n635 CS_BIAS.n506 24.4675
R31000 CS_BIAS.n635 CS_BIAS.n634 24.4675
R31001 CS_BIAS.n634 CS_BIAS.n633 24.4675
R31002 CS_BIAS.n628 CS_BIAS.n627 24.4675
R31003 CS_BIAS.n627 CS_BIAS.n510 24.4675
R31004 CS_BIAS.n623 CS_BIAS.n510 24.4675
R31005 CS_BIAS.n623 CS_BIAS.n622 24.4675
R31006 CS_BIAS.n622 CS_BIAS.n621 24.4675
R31007 CS_BIAS.n618 CS_BIAS.n617 24.4675
R31008 CS_BIAS.n617 CS_BIAS.n616 24.4675
R31009 CS_BIAS.n616 CS_BIAS.n514 24.4675
R31010 CS_BIAS.n612 CS_BIAS.n514 24.4675
R31011 CS_BIAS.n606 CS_BIAS.n516 24.4675
R31012 CS_BIAS.n606 CS_BIAS.n605 24.4675
R31013 CS_BIAS.n605 CS_BIAS.n604 24.4675
R31014 CS_BIAS.n604 CS_BIAS.n518 24.4675
R31015 CS_BIAS.n600 CS_BIAS.n518 24.4675
R31016 CS_BIAS.n598 CS_BIAS.n597 24.4675
R31017 CS_BIAS.n597 CS_BIAS.n520 24.4675
R31018 CS_BIAS.n593 CS_BIAS.n520 24.4675
R31019 CS_BIAS.n593 CS_BIAS.n592 24.4675
R31020 CS_BIAS.n587 CS_BIAS.n586 24.4675
R31021 CS_BIAS.n586 CS_BIAS.n585 24.4675
R31022 CS_BIAS.n585 CS_BIAS.n524 24.4675
R31023 CS_BIAS.n581 CS_BIAS.n524 24.4675
R31024 CS_BIAS.n579 CS_BIAS.n578 24.4675
R31025 CS_BIAS.n578 CS_BIAS.n526 24.4675
R31026 CS_BIAS.n574 CS_BIAS.n526 24.4675
R31027 CS_BIAS.n574 CS_BIAS.n573 24.4675
R31028 CS_BIAS.n573 CS_BIAS.n572 24.4675
R31029 CS_BIAS.n567 CS_BIAS.n566 24.4675
R31030 CS_BIAS.n566 CS_BIAS.n530 24.4675
R31031 CS_BIAS.n562 CS_BIAS.n530 24.4675
R31032 CS_BIAS.n562 CS_BIAS.n561 24.4675
R31033 CS_BIAS.n559 CS_BIAS.n532 24.4675
R31034 CS_BIAS.n555 CS_BIAS.n532 24.4675
R31035 CS_BIAS.n555 CS_BIAS.n554 24.4675
R31036 CS_BIAS.n554 CS_BIAS.n553 24.4675
R31037 CS_BIAS.n553 CS_BIAS.n534 24.4675
R31038 CS_BIAS.n547 CS_BIAS.n536 24.4675
R31039 CS_BIAS.n543 CS_BIAS.n536 24.4675
R31040 CS_BIAS.n543 CS_BIAS.n542 24.4675
R31041 CS_BIAS.n542 CS_BIAS.n541 24.4675
R31042 CS_BIAS.n495 CS_BIAS.n494 24.4675
R31043 CS_BIAS.n494 CS_BIAS.n336 24.4675
R31044 CS_BIAS.n490 CS_BIAS.n336 24.4675
R31045 CS_BIAS.n490 CS_BIAS.n489 24.4675
R31046 CS_BIAS.n484 CS_BIAS.n483 24.4675
R31047 CS_BIAS.n483 CS_BIAS.n482 24.4675
R31048 CS_BIAS.n482 CS_BIAS.n340 24.4675
R31049 CS_BIAS.n478 CS_BIAS.n340 24.4675
R31050 CS_BIAS.n478 CS_BIAS.n477 24.4675
R31051 CS_BIAS.n475 CS_BIAS.n342 24.4675
R31052 CS_BIAS.n471 CS_BIAS.n342 24.4675
R31053 CS_BIAS.n471 CS_BIAS.n470 24.4675
R31054 CS_BIAS.n470 CS_BIAS.n469 24.4675
R31055 CS_BIAS.n464 CS_BIAS.n463 24.4675
R31056 CS_BIAS.n463 CS_BIAS.n346 24.4675
R31057 CS_BIAS.n459 CS_BIAS.n346 24.4675
R31058 CS_BIAS.n459 CS_BIAS.n458 24.4675
R31059 CS_BIAS.n458 CS_BIAS.n457 24.4675
R31060 CS_BIAS.n454 CS_BIAS.n453 24.4675
R31061 CS_BIAS.n453 CS_BIAS.n452 24.4675
R31062 CS_BIAS.n452 CS_BIAS.n350 24.4675
R31063 CS_BIAS.n448 CS_BIAS.n350 24.4675
R31064 CS_BIAS.n442 CS_BIAS.n352 24.4675
R31065 CS_BIAS.n442 CS_BIAS.n441 24.4675
R31066 CS_BIAS.n441 CS_BIAS.n440 24.4675
R31067 CS_BIAS.n440 CS_BIAS.n354 24.4675
R31068 CS_BIAS.n436 CS_BIAS.n354 24.4675
R31069 CS_BIAS.n434 CS_BIAS.n433 24.4675
R31070 CS_BIAS.n433 CS_BIAS.n356 24.4675
R31071 CS_BIAS.n429 CS_BIAS.n356 24.4675
R31072 CS_BIAS.n429 CS_BIAS.n428 24.4675
R31073 CS_BIAS.n423 CS_BIAS.n422 24.4675
R31074 CS_BIAS.n422 CS_BIAS.n421 24.4675
R31075 CS_BIAS.n421 CS_BIAS.n360 24.4675
R31076 CS_BIAS.n417 CS_BIAS.n360 24.4675
R31077 CS_BIAS.n415 CS_BIAS.n414 24.4675
R31078 CS_BIAS.n414 CS_BIAS.n362 24.4675
R31079 CS_BIAS.n410 CS_BIAS.n362 24.4675
R31080 CS_BIAS.n410 CS_BIAS.n409 24.4675
R31081 CS_BIAS.n409 CS_BIAS.n408 24.4675
R31082 CS_BIAS.n403 CS_BIAS.n402 24.4675
R31083 CS_BIAS.n402 CS_BIAS.n366 24.4675
R31084 CS_BIAS.n398 CS_BIAS.n366 24.4675
R31085 CS_BIAS.n398 CS_BIAS.n397 24.4675
R31086 CS_BIAS.n395 CS_BIAS.n368 24.4675
R31087 CS_BIAS.n391 CS_BIAS.n368 24.4675
R31088 CS_BIAS.n391 CS_BIAS.n390 24.4675
R31089 CS_BIAS.n390 CS_BIAS.n389 24.4675
R31090 CS_BIAS.n389 CS_BIAS.n370 24.4675
R31091 CS_BIAS.n383 CS_BIAS.n372 24.4675
R31092 CS_BIAS.n379 CS_BIAS.n372 24.4675
R31093 CS_BIAS.n379 CS_BIAS.n378 24.4675
R31094 CS_BIAS.n378 CS_BIAS.n377 24.4675
R31095 CS_BIAS.n251 CS_BIAS.n250 24.4675
R31096 CS_BIAS.n250 CS_BIAS.n92 24.4675
R31097 CS_BIAS.n246 CS_BIAS.n92 24.4675
R31098 CS_BIAS.n246 CS_BIAS.n245 24.4675
R31099 CS_BIAS.n240 CS_BIAS.n239 24.4675
R31100 CS_BIAS.n239 CS_BIAS.n238 24.4675
R31101 CS_BIAS.n238 CS_BIAS.n96 24.4675
R31102 CS_BIAS.n234 CS_BIAS.n96 24.4675
R31103 CS_BIAS.n234 CS_BIAS.n233 24.4675
R31104 CS_BIAS.n231 CS_BIAS.n98 24.4675
R31105 CS_BIAS.n227 CS_BIAS.n98 24.4675
R31106 CS_BIAS.n227 CS_BIAS.n226 24.4675
R31107 CS_BIAS.n226 CS_BIAS.n225 24.4675
R31108 CS_BIAS.n220 CS_BIAS.n219 24.4675
R31109 CS_BIAS.n219 CS_BIAS.n102 24.4675
R31110 CS_BIAS.n215 CS_BIAS.n102 24.4675
R31111 CS_BIAS.n215 CS_BIAS.n214 24.4675
R31112 CS_BIAS.n214 CS_BIAS.n213 24.4675
R31113 CS_BIAS.n210 CS_BIAS.n209 24.4675
R31114 CS_BIAS.n209 CS_BIAS.n208 24.4675
R31115 CS_BIAS.n208 CS_BIAS.n106 24.4675
R31116 CS_BIAS.n204 CS_BIAS.n106 24.4675
R31117 CS_BIAS.n198 CS_BIAS.n108 24.4675
R31118 CS_BIAS.n198 CS_BIAS.n197 24.4675
R31119 CS_BIAS.n197 CS_BIAS.n196 24.4675
R31120 CS_BIAS.n196 CS_BIAS.n110 24.4675
R31121 CS_BIAS.n192 CS_BIAS.n110 24.4675
R31122 CS_BIAS.n190 CS_BIAS.n189 24.4675
R31123 CS_BIAS.n189 CS_BIAS.n112 24.4675
R31124 CS_BIAS.n185 CS_BIAS.n112 24.4675
R31125 CS_BIAS.n185 CS_BIAS.n184 24.4675
R31126 CS_BIAS.n179 CS_BIAS.n178 24.4675
R31127 CS_BIAS.n178 CS_BIAS.n177 24.4675
R31128 CS_BIAS.n177 CS_BIAS.n116 24.4675
R31129 CS_BIAS.n173 CS_BIAS.n116 24.4675
R31130 CS_BIAS.n171 CS_BIAS.n170 24.4675
R31131 CS_BIAS.n170 CS_BIAS.n118 24.4675
R31132 CS_BIAS.n166 CS_BIAS.n118 24.4675
R31133 CS_BIAS.n166 CS_BIAS.n165 24.4675
R31134 CS_BIAS.n165 CS_BIAS.n164 24.4675
R31135 CS_BIAS.n159 CS_BIAS.n158 24.4675
R31136 CS_BIAS.n158 CS_BIAS.n122 24.4675
R31137 CS_BIAS.n154 CS_BIAS.n122 24.4675
R31138 CS_BIAS.n154 CS_BIAS.n153 24.4675
R31139 CS_BIAS.n151 CS_BIAS.n124 24.4675
R31140 CS_BIAS.n147 CS_BIAS.n124 24.4675
R31141 CS_BIAS.n147 CS_BIAS.n146 24.4675
R31142 CS_BIAS.n146 CS_BIAS.n145 24.4675
R31143 CS_BIAS.n145 CS_BIAS.n126 24.4675
R31144 CS_BIAS.n139 CS_BIAS.n128 24.4675
R31145 CS_BIAS.n135 CS_BIAS.n128 24.4675
R31146 CS_BIAS.n135 CS_BIAS.n134 24.4675
R31147 CS_BIAS.n134 CS_BIAS.n133 24.4675
R31148 CS_BIAS.n332 CS_BIAS.n331 24.4675
R31149 CS_BIAS.n331 CS_BIAS.n1 24.4675
R31150 CS_BIAS.n327 CS_BIAS.n1 24.4675
R31151 CS_BIAS.n327 CS_BIAS.n326 24.4675
R31152 CS_BIAS.n321 CS_BIAS.n320 24.4675
R31153 CS_BIAS.n320 CS_BIAS.n319 24.4675
R31154 CS_BIAS.n319 CS_BIAS.n5 24.4675
R31155 CS_BIAS.n315 CS_BIAS.n5 24.4675
R31156 CS_BIAS.n315 CS_BIAS.n314 24.4675
R31157 CS_BIAS.n312 CS_BIAS.n7 24.4675
R31158 CS_BIAS.n308 CS_BIAS.n7 24.4675
R31159 CS_BIAS.n308 CS_BIAS.n307 24.4675
R31160 CS_BIAS.n307 CS_BIAS.n306 24.4675
R31161 CS_BIAS.n301 CS_BIAS.n300 24.4675
R31162 CS_BIAS.n300 CS_BIAS.n11 24.4675
R31163 CS_BIAS.n296 CS_BIAS.n11 24.4675
R31164 CS_BIAS.n296 CS_BIAS.n295 24.4675
R31165 CS_BIAS.n295 CS_BIAS.n294 24.4675
R31166 CS_BIAS.n291 CS_BIAS.n290 24.4675
R31167 CS_BIAS.n290 CS_BIAS.n289 24.4675
R31168 CS_BIAS.n289 CS_BIAS.n15 24.4675
R31169 CS_BIAS.n285 CS_BIAS.n15 24.4675
R31170 CS_BIAS.n279 CS_BIAS.n17 24.4675
R31171 CS_BIAS.n279 CS_BIAS.n278 24.4675
R31172 CS_BIAS.n278 CS_BIAS.n277 24.4675
R31173 CS_BIAS.n277 CS_BIAS.n19 24.4675
R31174 CS_BIAS.n273 CS_BIAS.n19 24.4675
R31175 CS_BIAS.n271 CS_BIAS.n270 24.4675
R31176 CS_BIAS.n270 CS_BIAS.n21 24.4675
R31177 CS_BIAS.n266 CS_BIAS.n21 24.4675
R31178 CS_BIAS.n266 CS_BIAS.n265 24.4675
R31179 CS_BIAS.n88 CS_BIAS.n87 24.4675
R31180 CS_BIAS.n87 CS_BIAS.n86 24.4675
R31181 CS_BIAS.n86 CS_BIAS.n25 24.4675
R31182 CS_BIAS.n82 CS_BIAS.n25 24.4675
R31183 CS_BIAS.n80 CS_BIAS.n79 24.4675
R31184 CS_BIAS.n79 CS_BIAS.n27 24.4675
R31185 CS_BIAS.n75 CS_BIAS.n27 24.4675
R31186 CS_BIAS.n75 CS_BIAS.n74 24.4675
R31187 CS_BIAS.n74 CS_BIAS.n73 24.4675
R31188 CS_BIAS.n68 CS_BIAS.n67 24.4675
R31189 CS_BIAS.n67 CS_BIAS.n31 24.4675
R31190 CS_BIAS.n63 CS_BIAS.n31 24.4675
R31191 CS_BIAS.n63 CS_BIAS.n62 24.4675
R31192 CS_BIAS.n60 CS_BIAS.n33 24.4675
R31193 CS_BIAS.n56 CS_BIAS.n33 24.4675
R31194 CS_BIAS.n56 CS_BIAS.n55 24.4675
R31195 CS_BIAS.n55 CS_BIAS.n54 24.4675
R31196 CS_BIAS.n54 CS_BIAS.n35 24.4675
R31197 CS_BIAS.n48 CS_BIAS.n37 24.4675
R31198 CS_BIAS.n44 CS_BIAS.n37 24.4675
R31199 CS_BIAS.n44 CS_BIAS.n43 24.4675
R31200 CS_BIAS.n43 CS_BIAS.n42 24.4675
R31201 CS_BIAS.n1533 CS_BIAS.n1532 24.4675
R31202 CS_BIAS.n1534 CS_BIAS.n1533 24.4675
R31203 CS_BIAS.n1534 CS_BIAS.n1527 24.4675
R31204 CS_BIAS.n1538 CS_BIAS.n1527 24.4675
R31205 CS_BIAS.n1544 CS_BIAS.n1525 24.4675
R31206 CS_BIAS.n1545 CS_BIAS.n1544 24.4675
R31207 CS_BIAS.n1546 CS_BIAS.n1545 24.4675
R31208 CS_BIAS.n1546 CS_BIAS.n1523 24.4675
R31209 CS_BIAS.n1550 CS_BIAS.n1523 24.4675
R31210 CS_BIAS.n1553 CS_BIAS.n1552 24.4675
R31211 CS_BIAS.n1553 CS_BIAS.n1521 24.4675
R31212 CS_BIAS.n1557 CS_BIAS.n1521 24.4675
R31213 CS_BIAS.n1558 CS_BIAS.n1557 24.4675
R31214 CS_BIAS.n1564 CS_BIAS.n1563 24.4675
R31215 CS_BIAS.n1565 CS_BIAS.n1564 24.4675
R31216 CS_BIAS.n1565 CS_BIAS.n1517 24.4675
R31217 CS_BIAS.n1569 CS_BIAS.n1517 24.4675
R31218 CS_BIAS.n1570 CS_BIAS.n1569 24.4675
R31219 CS_BIAS.n1572 CS_BIAS.n1515 24.4675
R31220 CS_BIAS.n1576 CS_BIAS.n1515 24.4675
R31221 CS_BIAS.n1577 CS_BIAS.n1576 24.4675
R31222 CS_BIAS.n1578 CS_BIAS.n1577 24.4675
R31223 CS_BIAS.n1584 CS_BIAS.n1583 24.4675
R31224 CS_BIAS.n1584 CS_BIAS.n1511 24.4675
R31225 CS_BIAS.n1588 CS_BIAS.n1511 24.4675
R31226 CS_BIAS.n1589 CS_BIAS.n1588 24.4675
R31227 CS_BIAS.n1591 CS_BIAS.n1509 24.4675
R31228 CS_BIAS.n1595 CS_BIAS.n1509 24.4675
R31229 CS_BIAS.n1596 CS_BIAS.n1595 24.4675
R31230 CS_BIAS.n1597 CS_BIAS.n1596 24.4675
R31231 CS_BIAS.n1597 CS_BIAS.n1507 24.4675
R31232 CS_BIAS.n1603 CS_BIAS.n1505 24.4675
R31233 CS_BIAS.n1607 CS_BIAS.n1505 24.4675
R31234 CS_BIAS.n1608 CS_BIAS.n1607 24.4675
R31235 CS_BIAS.n1609 CS_BIAS.n1608 24.4675
R31236 CS_BIAS.n1613 CS_BIAS.n1612 24.4675
R31237 CS_BIAS.n1614 CS_BIAS.n1613 24.4675
R31238 CS_BIAS.n1614 CS_BIAS.n1501 24.4675
R31239 CS_BIAS.n1618 CS_BIAS.n1501 24.4675
R31240 CS_BIAS.n1619 CS_BIAS.n1618 24.4675
R31241 CS_BIAS.n1625 CS_BIAS.n1624 24.4675
R31242 CS_BIAS.n1626 CS_BIAS.n1625 24.4675
R31243 CS_BIAS.n1626 CS_BIAS.n1497 24.4675
R31244 CS_BIAS.n1630 CS_BIAS.n1497 24.4675
R31245 CS_BIAS.n1633 CS_BIAS.n1632 24.4675
R31246 CS_BIAS.n1633 CS_BIAS.n1495 24.4675
R31247 CS_BIAS.n1637 CS_BIAS.n1495 24.4675
R31248 CS_BIAS.n1638 CS_BIAS.n1637 24.4675
R31249 CS_BIAS.n1639 CS_BIAS.n1638 24.4675
R31250 CS_BIAS.n1645 CS_BIAS.n1644 24.4675
R31251 CS_BIAS.n1645 CS_BIAS.n1491 24.4675
R31252 CS_BIAS.n1649 CS_BIAS.n1491 24.4675
R31253 CS_BIAS.n1650 CS_BIAS.n1649 24.4675
R31254 CS_BIAS.n1369 CS_BIAS.n1368 24.4675
R31255 CS_BIAS.n1370 CS_BIAS.n1369 24.4675
R31256 CS_BIAS.n1370 CS_BIAS.n1363 24.4675
R31257 CS_BIAS.n1374 CS_BIAS.n1363 24.4675
R31258 CS_BIAS.n1380 CS_BIAS.n1361 24.4675
R31259 CS_BIAS.n1381 CS_BIAS.n1380 24.4675
R31260 CS_BIAS.n1382 CS_BIAS.n1381 24.4675
R31261 CS_BIAS.n1382 CS_BIAS.n1359 24.4675
R31262 CS_BIAS.n1386 CS_BIAS.n1359 24.4675
R31263 CS_BIAS.n1389 CS_BIAS.n1388 24.4675
R31264 CS_BIAS.n1389 CS_BIAS.n1357 24.4675
R31265 CS_BIAS.n1393 CS_BIAS.n1357 24.4675
R31266 CS_BIAS.n1394 CS_BIAS.n1393 24.4675
R31267 CS_BIAS.n1400 CS_BIAS.n1399 24.4675
R31268 CS_BIAS.n1401 CS_BIAS.n1400 24.4675
R31269 CS_BIAS.n1401 CS_BIAS.n1353 24.4675
R31270 CS_BIAS.n1405 CS_BIAS.n1353 24.4675
R31271 CS_BIAS.n1406 CS_BIAS.n1405 24.4675
R31272 CS_BIAS.n1408 CS_BIAS.n1351 24.4675
R31273 CS_BIAS.n1412 CS_BIAS.n1351 24.4675
R31274 CS_BIAS.n1413 CS_BIAS.n1412 24.4675
R31275 CS_BIAS.n1414 CS_BIAS.n1413 24.4675
R31276 CS_BIAS.n1420 CS_BIAS.n1419 24.4675
R31277 CS_BIAS.n1420 CS_BIAS.n1347 24.4675
R31278 CS_BIAS.n1424 CS_BIAS.n1347 24.4675
R31279 CS_BIAS.n1425 CS_BIAS.n1424 24.4675
R31280 CS_BIAS.n1427 CS_BIAS.n1345 24.4675
R31281 CS_BIAS.n1431 CS_BIAS.n1345 24.4675
R31282 CS_BIAS.n1432 CS_BIAS.n1431 24.4675
R31283 CS_BIAS.n1433 CS_BIAS.n1432 24.4675
R31284 CS_BIAS.n1433 CS_BIAS.n1343 24.4675
R31285 CS_BIAS.n1439 CS_BIAS.n1341 24.4675
R31286 CS_BIAS.n1443 CS_BIAS.n1341 24.4675
R31287 CS_BIAS.n1444 CS_BIAS.n1443 24.4675
R31288 CS_BIAS.n1445 CS_BIAS.n1444 24.4675
R31289 CS_BIAS.n1449 CS_BIAS.n1448 24.4675
R31290 CS_BIAS.n1450 CS_BIAS.n1449 24.4675
R31291 CS_BIAS.n1450 CS_BIAS.n1337 24.4675
R31292 CS_BIAS.n1454 CS_BIAS.n1337 24.4675
R31293 CS_BIAS.n1455 CS_BIAS.n1454 24.4675
R31294 CS_BIAS.n1461 CS_BIAS.n1460 24.4675
R31295 CS_BIAS.n1462 CS_BIAS.n1461 24.4675
R31296 CS_BIAS.n1462 CS_BIAS.n1333 24.4675
R31297 CS_BIAS.n1466 CS_BIAS.n1333 24.4675
R31298 CS_BIAS.n1469 CS_BIAS.n1468 24.4675
R31299 CS_BIAS.n1469 CS_BIAS.n1331 24.4675
R31300 CS_BIAS.n1473 CS_BIAS.n1331 24.4675
R31301 CS_BIAS.n1474 CS_BIAS.n1473 24.4675
R31302 CS_BIAS.n1475 CS_BIAS.n1474 24.4675
R31303 CS_BIAS.n1481 CS_BIAS.n1480 24.4675
R31304 CS_BIAS.n1481 CS_BIAS.n1327 24.4675
R31305 CS_BIAS.n1485 CS_BIAS.n1327 24.4675
R31306 CS_BIAS.n1486 CS_BIAS.n1485 24.4675
R31307 CS_BIAS.n1205 CS_BIAS.n1204 24.4675
R31308 CS_BIAS.n1206 CS_BIAS.n1205 24.4675
R31309 CS_BIAS.n1206 CS_BIAS.n1199 24.4675
R31310 CS_BIAS.n1210 CS_BIAS.n1199 24.4675
R31311 CS_BIAS.n1216 CS_BIAS.n1197 24.4675
R31312 CS_BIAS.n1217 CS_BIAS.n1216 24.4675
R31313 CS_BIAS.n1218 CS_BIAS.n1217 24.4675
R31314 CS_BIAS.n1218 CS_BIAS.n1195 24.4675
R31315 CS_BIAS.n1222 CS_BIAS.n1195 24.4675
R31316 CS_BIAS.n1225 CS_BIAS.n1224 24.4675
R31317 CS_BIAS.n1225 CS_BIAS.n1193 24.4675
R31318 CS_BIAS.n1229 CS_BIAS.n1193 24.4675
R31319 CS_BIAS.n1230 CS_BIAS.n1229 24.4675
R31320 CS_BIAS.n1236 CS_BIAS.n1235 24.4675
R31321 CS_BIAS.n1237 CS_BIAS.n1236 24.4675
R31322 CS_BIAS.n1237 CS_BIAS.n1189 24.4675
R31323 CS_BIAS.n1241 CS_BIAS.n1189 24.4675
R31324 CS_BIAS.n1242 CS_BIAS.n1241 24.4675
R31325 CS_BIAS.n1244 CS_BIAS.n1187 24.4675
R31326 CS_BIAS.n1248 CS_BIAS.n1187 24.4675
R31327 CS_BIAS.n1249 CS_BIAS.n1248 24.4675
R31328 CS_BIAS.n1250 CS_BIAS.n1249 24.4675
R31329 CS_BIAS.n1256 CS_BIAS.n1255 24.4675
R31330 CS_BIAS.n1256 CS_BIAS.n1183 24.4675
R31331 CS_BIAS.n1260 CS_BIAS.n1183 24.4675
R31332 CS_BIAS.n1261 CS_BIAS.n1260 24.4675
R31333 CS_BIAS.n1263 CS_BIAS.n1181 24.4675
R31334 CS_BIAS.n1267 CS_BIAS.n1181 24.4675
R31335 CS_BIAS.n1268 CS_BIAS.n1267 24.4675
R31336 CS_BIAS.n1269 CS_BIAS.n1268 24.4675
R31337 CS_BIAS.n1269 CS_BIAS.n1179 24.4675
R31338 CS_BIAS.n1275 CS_BIAS.n1177 24.4675
R31339 CS_BIAS.n1279 CS_BIAS.n1177 24.4675
R31340 CS_BIAS.n1280 CS_BIAS.n1279 24.4675
R31341 CS_BIAS.n1281 CS_BIAS.n1280 24.4675
R31342 CS_BIAS.n1285 CS_BIAS.n1284 24.4675
R31343 CS_BIAS.n1286 CS_BIAS.n1285 24.4675
R31344 CS_BIAS.n1286 CS_BIAS.n1173 24.4675
R31345 CS_BIAS.n1290 CS_BIAS.n1173 24.4675
R31346 CS_BIAS.n1291 CS_BIAS.n1290 24.4675
R31347 CS_BIAS.n1297 CS_BIAS.n1296 24.4675
R31348 CS_BIAS.n1298 CS_BIAS.n1297 24.4675
R31349 CS_BIAS.n1298 CS_BIAS.n1169 24.4675
R31350 CS_BIAS.n1302 CS_BIAS.n1169 24.4675
R31351 CS_BIAS.n1305 CS_BIAS.n1304 24.4675
R31352 CS_BIAS.n1305 CS_BIAS.n1167 24.4675
R31353 CS_BIAS.n1309 CS_BIAS.n1167 24.4675
R31354 CS_BIAS.n1310 CS_BIAS.n1309 24.4675
R31355 CS_BIAS.n1311 CS_BIAS.n1310 24.4675
R31356 CS_BIAS.n1317 CS_BIAS.n1316 24.4675
R31357 CS_BIAS.n1317 CS_BIAS.n1163 24.4675
R31358 CS_BIAS.n1321 CS_BIAS.n1163 24.4675
R31359 CS_BIAS.n1322 CS_BIAS.n1321 24.4675
R31360 CS_BIAS.n964 CS_BIAS.n963 24.4675
R31361 CS_BIAS.n965 CS_BIAS.n964 24.4675
R31362 CS_BIAS.n965 CS_BIAS.n958 24.4675
R31363 CS_BIAS.n969 CS_BIAS.n958 24.4675
R31364 CS_BIAS.n975 CS_BIAS.n956 24.4675
R31365 CS_BIAS.n976 CS_BIAS.n975 24.4675
R31366 CS_BIAS.n977 CS_BIAS.n976 24.4675
R31367 CS_BIAS.n977 CS_BIAS.n954 24.4675
R31368 CS_BIAS.n981 CS_BIAS.n954 24.4675
R31369 CS_BIAS.n984 CS_BIAS.n983 24.4675
R31370 CS_BIAS.n984 CS_BIAS.n952 24.4675
R31371 CS_BIAS.n988 CS_BIAS.n952 24.4675
R31372 CS_BIAS.n989 CS_BIAS.n988 24.4675
R31373 CS_BIAS.n995 CS_BIAS.n994 24.4675
R31374 CS_BIAS.n996 CS_BIAS.n995 24.4675
R31375 CS_BIAS.n996 CS_BIAS.n948 24.4675
R31376 CS_BIAS.n1000 CS_BIAS.n948 24.4675
R31377 CS_BIAS.n1001 CS_BIAS.n1000 24.4675
R31378 CS_BIAS.n1003 CS_BIAS.n946 24.4675
R31379 CS_BIAS.n1007 CS_BIAS.n946 24.4675
R31380 CS_BIAS.n1008 CS_BIAS.n1007 24.4675
R31381 CS_BIAS.n1009 CS_BIAS.n1008 24.4675
R31382 CS_BIAS.n1015 CS_BIAS.n1014 24.4675
R31383 CS_BIAS.n1015 CS_BIAS.n942 24.4675
R31384 CS_BIAS.n1019 CS_BIAS.n942 24.4675
R31385 CS_BIAS.n1020 CS_BIAS.n1019 24.4675
R31386 CS_BIAS.n1022 CS_BIAS.n940 24.4675
R31387 CS_BIAS.n1026 CS_BIAS.n940 24.4675
R31388 CS_BIAS.n1027 CS_BIAS.n1026 24.4675
R31389 CS_BIAS.n1028 CS_BIAS.n1027 24.4675
R31390 CS_BIAS.n1028 CS_BIAS.n938 24.4675
R31391 CS_BIAS.n1034 CS_BIAS.n936 24.4675
R31392 CS_BIAS.n1038 CS_BIAS.n936 24.4675
R31393 CS_BIAS.n1039 CS_BIAS.n1038 24.4675
R31394 CS_BIAS.n1040 CS_BIAS.n1039 24.4675
R31395 CS_BIAS.n1044 CS_BIAS.n1043 24.4675
R31396 CS_BIAS.n1045 CS_BIAS.n1044 24.4675
R31397 CS_BIAS.n1045 CS_BIAS.n932 24.4675
R31398 CS_BIAS.n1049 CS_BIAS.n932 24.4675
R31399 CS_BIAS.n1050 CS_BIAS.n1049 24.4675
R31400 CS_BIAS.n1056 CS_BIAS.n1055 24.4675
R31401 CS_BIAS.n1057 CS_BIAS.n1056 24.4675
R31402 CS_BIAS.n1057 CS_BIAS.n928 24.4675
R31403 CS_BIAS.n1061 CS_BIAS.n928 24.4675
R31404 CS_BIAS.n1064 CS_BIAS.n1063 24.4675
R31405 CS_BIAS.n1064 CS_BIAS.n926 24.4675
R31406 CS_BIAS.n1068 CS_BIAS.n926 24.4675
R31407 CS_BIAS.n1069 CS_BIAS.n1068 24.4675
R31408 CS_BIAS.n1070 CS_BIAS.n1069 24.4675
R31409 CS_BIAS.n1076 CS_BIAS.n1075 24.4675
R31410 CS_BIAS.n1076 CS_BIAS.n922 24.4675
R31411 CS_BIAS.n1080 CS_BIAS.n922 24.4675
R31412 CS_BIAS.n1081 CS_BIAS.n1080 24.4675
R31413 CS_BIAS.n1154 CS_BIAS.n1153 24.4675
R31414 CS_BIAS.n1154 CS_BIAS.n828 24.4675
R31415 CS_BIAS.n1158 CS_BIAS.n828 24.4675
R31416 CS_BIAS.n1159 CS_BIAS.n1158 24.4675
R31417 CS_BIAS.n1134 CS_BIAS.n1133 24.4675
R31418 CS_BIAS.n1135 CS_BIAS.n1134 24.4675
R31419 CS_BIAS.n1135 CS_BIAS.n834 24.4675
R31420 CS_BIAS.n1139 CS_BIAS.n834 24.4675
R31421 CS_BIAS.n1142 CS_BIAS.n1141 24.4675
R31422 CS_BIAS.n1142 CS_BIAS.n832 24.4675
R31423 CS_BIAS.n1146 CS_BIAS.n832 24.4675
R31424 CS_BIAS.n1147 CS_BIAS.n1146 24.4675
R31425 CS_BIAS.n1148 CS_BIAS.n1147 24.4675
R31426 CS_BIAS.n1112 CS_BIAS.n842 24.4675
R31427 CS_BIAS.n1116 CS_BIAS.n842 24.4675
R31428 CS_BIAS.n1117 CS_BIAS.n1116 24.4675
R31429 CS_BIAS.n1118 CS_BIAS.n1117 24.4675
R31430 CS_BIAS.n1122 CS_BIAS.n1121 24.4675
R31431 CS_BIAS.n1123 CS_BIAS.n1122 24.4675
R31432 CS_BIAS.n1123 CS_BIAS.n838 24.4675
R31433 CS_BIAS.n1127 CS_BIAS.n838 24.4675
R31434 CS_BIAS.n1128 CS_BIAS.n1127 24.4675
R31435 CS_BIAS.n1093 CS_BIAS.n1092 24.4675
R31436 CS_BIAS.n1093 CS_BIAS.n848 24.4675
R31437 CS_BIAS.n1097 CS_BIAS.n848 24.4675
R31438 CS_BIAS.n1098 CS_BIAS.n1097 24.4675
R31439 CS_BIAS.n1100 CS_BIAS.n846 24.4675
R31440 CS_BIAS.n1104 CS_BIAS.n846 24.4675
R31441 CS_BIAS.n1105 CS_BIAS.n1104 24.4675
R31442 CS_BIAS.n1106 CS_BIAS.n1105 24.4675
R31443 CS_BIAS.n1106 CS_BIAS.n844 24.4675
R31444 CS_BIAS.n870 CS_BIAS.n869 24.4675
R31445 CS_BIAS.n871 CS_BIAS.n870 24.4675
R31446 CS_BIAS.n871 CS_BIAS.n864 24.4675
R31447 CS_BIAS.n875 CS_BIAS.n864 24.4675
R31448 CS_BIAS.n881 CS_BIAS.n862 24.4675
R31449 CS_BIAS.n882 CS_BIAS.n881 24.4675
R31450 CS_BIAS.n883 CS_BIAS.n882 24.4675
R31451 CS_BIAS.n883 CS_BIAS.n860 24.4675
R31452 CS_BIAS.n887 CS_BIAS.n860 24.4675
R31453 CS_BIAS.n890 CS_BIAS.n889 24.4675
R31454 CS_BIAS.n890 CS_BIAS.n858 24.4675
R31455 CS_BIAS.n894 CS_BIAS.n858 24.4675
R31456 CS_BIAS.n895 CS_BIAS.n894 24.4675
R31457 CS_BIAS.n901 CS_BIAS.n900 24.4675
R31458 CS_BIAS.n902 CS_BIAS.n901 24.4675
R31459 CS_BIAS.n902 CS_BIAS.n854 24.4675
R31460 CS_BIAS.n906 CS_BIAS.n854 24.4675
R31461 CS_BIAS.n907 CS_BIAS.n906 24.4675
R31462 CS_BIAS.n909 CS_BIAS.n852 24.4675
R31463 CS_BIAS.n913 CS_BIAS.n852 24.4675
R31464 CS_BIAS.n914 CS_BIAS.n913 24.4675
R31465 CS_BIAS.n915 CS_BIAS.n914 24.4675
R31466 CS_BIAS.n745 CS_BIAS.n744 24.2228
R31467 CS_BIAS.n763 CS_BIAS.n762 24.2228
R31468 CS_BIAS.n599 CS_BIAS.n598 24.2228
R31469 CS_BIAS.n581 CS_BIAS.n580 24.2228
R31470 CS_BIAS.n435 CS_BIAS.n434 24.2228
R31471 CS_BIAS.n417 CS_BIAS.n416 24.2228
R31472 CS_BIAS.n191 CS_BIAS.n190 24.2228
R31473 CS_BIAS.n173 CS_BIAS.n172 24.2228
R31474 CS_BIAS.n272 CS_BIAS.n271 24.2228
R31475 CS_BIAS.n82 CS_BIAS.n81 24.2228
R31476 CS_BIAS.n1572 CS_BIAS.n1571 24.2228
R31477 CS_BIAS.n1590 CS_BIAS.n1589 24.2228
R31478 CS_BIAS.n1408 CS_BIAS.n1407 24.2228
R31479 CS_BIAS.n1426 CS_BIAS.n1425 24.2228
R31480 CS_BIAS.n1244 CS_BIAS.n1243 24.2228
R31481 CS_BIAS.n1262 CS_BIAS.n1261 24.2228
R31482 CS_BIAS.n1003 CS_BIAS.n1002 24.2228
R31483 CS_BIAS.n1021 CS_BIAS.n1020 24.2228
R31484 CS_BIAS.n1099 CS_BIAS.n1098 24.2228
R31485 CS_BIAS.n909 CS_BIAS.n908 24.2228
R31486 CS_BIAS.n725 CS_BIAS.n724 23.7335
R31487 CS_BIAS.n782 CS_BIAS.n676 23.7335
R31488 CS_BIAS.n618 CS_BIAS.n512 23.7335
R31489 CS_BIAS.n561 CS_BIAS.n560 23.7335
R31490 CS_BIAS.n454 CS_BIAS.n348 23.7335
R31491 CS_BIAS.n397 CS_BIAS.n396 23.7335
R31492 CS_BIAS.n210 CS_BIAS.n104 23.7335
R31493 CS_BIAS.n153 CS_BIAS.n152 23.7335
R31494 CS_BIAS.n291 CS_BIAS.n13 23.7335
R31495 CS_BIAS.n62 CS_BIAS.n61 23.7335
R31496 CS_BIAS.n1552 CS_BIAS.n1551 23.7335
R31497 CS_BIAS.n1609 CS_BIAS.n1503 23.7335
R31498 CS_BIAS.n1388 CS_BIAS.n1387 23.7335
R31499 CS_BIAS.n1445 CS_BIAS.n1339 23.7335
R31500 CS_BIAS.n1224 CS_BIAS.n1223 23.7335
R31501 CS_BIAS.n1281 CS_BIAS.n1175 23.7335
R31502 CS_BIAS.n983 CS_BIAS.n982 23.7335
R31503 CS_BIAS.n1040 CS_BIAS.n934 23.7335
R31504 CS_BIAS.n1118 CS_BIAS.n840 23.7335
R31505 CS_BIAS.n889 CS_BIAS.n888 23.7335
R31506 CS_BIAS.n705 CS_BIAS.n702 23.2442
R31507 CS_BIAS.n804 CS_BIAS.n803 23.2442
R31508 CS_BIAS.n640 CS_BIAS.n639 23.2442
R31509 CS_BIAS.n541 CS_BIAS.n538 23.2442
R31510 CS_BIAS.n476 CS_BIAS.n475 23.2442
R31511 CS_BIAS.n377 CS_BIAS.n374 23.2442
R31512 CS_BIAS.n232 CS_BIAS.n231 23.2442
R31513 CS_BIAS.n133 CS_BIAS.n130 23.2442
R31514 CS_BIAS.n313 CS_BIAS.n312 23.2442
R31515 CS_BIAS.n42 CS_BIAS.n39 23.2442
R31516 CS_BIAS.n1532 CS_BIAS.n1529 23.2442
R31517 CS_BIAS.n1631 CS_BIAS.n1630 23.2442
R31518 CS_BIAS.n1368 CS_BIAS.n1365 23.2442
R31519 CS_BIAS.n1467 CS_BIAS.n1466 23.2442
R31520 CS_BIAS.n1204 CS_BIAS.n1201 23.2442
R31521 CS_BIAS.n1303 CS_BIAS.n1302 23.2442
R31522 CS_BIAS.n963 CS_BIAS.n960 23.2442
R31523 CS_BIAS.n1062 CS_BIAS.n1061 23.2442
R31524 CS_BIAS.n1140 CS_BIAS.n1139 23.2442
R31525 CS_BIAS.n869 CS_BIAS.n866 23.2442
R31526 CS_BIAS.n824 CS_BIAS.n823 22.7548
R31527 CS_BIAS.n660 CS_BIAS.n659 22.7548
R31528 CS_BIAS.n496 CS_BIAS.n495 22.7548
R31529 CS_BIAS.n252 CS_BIAS.n251 22.7548
R31530 CS_BIAS.n333 CS_BIAS.n332 22.7548
R31531 CS_BIAS.n1651 CS_BIAS.n1650 22.7548
R31532 CS_BIAS.n1487 CS_BIAS.n1486 22.7548
R31533 CS_BIAS.n1323 CS_BIAS.n1322 22.7548
R31534 CS_BIAS.n1082 CS_BIAS.n1081 22.7548
R31535 CS_BIAS.n1160 CS_BIAS.n1159 22.7548
R31536 CS_BIAS.n702 CS_BIAS.t49 15.4195
R31537 CS_BIAS.n724 CS_BIAS.t66 15.4195
R31538 CS_BIAS.n744 CS_BIAS.t39 15.4195
R31539 CS_BIAS.n763 CS_BIAS.t36 15.4195
R31540 CS_BIAS.n676 CS_BIAS.t54 15.4195
R31541 CS_BIAS.n804 CS_BIAS.t75 15.4195
R31542 CS_BIAS.n824 CS_BIAS.t93 15.4195
R31543 CS_BIAS.n660 CS_BIAS.t61 15.4195
R31544 CS_BIAS.n640 CS_BIAS.t47 15.4195
R31545 CS_BIAS.n512 CS_BIAS.t87 15.4195
R31546 CS_BIAS.n599 CS_BIAS.t69 15.4195
R31547 CS_BIAS.n580 CS_BIAS.t72 15.4195
R31548 CS_BIAS.n560 CS_BIAS.t33 15.4195
R31549 CS_BIAS.n538 CS_BIAS.t79 15.4195
R31550 CS_BIAS.n496 CS_BIAS.t95 15.4195
R31551 CS_BIAS.n476 CS_BIAS.t76 15.4195
R31552 CS_BIAS.n348 CS_BIAS.t55 15.4195
R31553 CS_BIAS.n435 CS_BIAS.t37 15.4195
R31554 CS_BIAS.n416 CS_BIAS.t43 15.4195
R31555 CS_BIAS.n396 CS_BIAS.t67 15.4195
R31556 CS_BIAS.n374 CS_BIAS.t50 15.4195
R31557 CS_BIAS.n252 CS_BIAS.t12 15.4195
R31558 CS_BIAS.n232 CS_BIAS.t2 15.4195
R31559 CS_BIAS.n104 CS_BIAS.t30 15.4195
R31560 CS_BIAS.n191 CS_BIAS.t18 15.4195
R31561 CS_BIAS.n172 CS_BIAS.t8 15.4195
R31562 CS_BIAS.n152 CS_BIAS.t24 15.4195
R31563 CS_BIAS.n130 CS_BIAS.t16 15.4195
R31564 CS_BIAS.n333 CS_BIAS.t85 15.4195
R31565 CS_BIAS.n313 CS_BIAS.t45 15.4195
R31566 CS_BIAS.n13 CS_BIAS.t57 15.4195
R31567 CS_BIAS.n272 CS_BIAS.t80 15.4195
R31568 CS_BIAS.n81 CS_BIAS.t91 15.4195
R31569 CS_BIAS.n61 CS_BIAS.t62 15.4195
R31570 CS_BIAS.n39 CS_BIAS.t84 15.4195
R31571 CS_BIAS.n1529 CS_BIAS.t59 15.4195
R31572 CS_BIAS.n1551 CS_BIAS.t82 15.4195
R31573 CS_BIAS.n1571 CS_BIAS.t38 15.4195
R31574 CS_BIAS.n1590 CS_BIAS.t34 15.4195
R31575 CS_BIAS.n1503 CS_BIAS.t73 15.4195
R31576 CS_BIAS.n1631 CS_BIAS.t90 15.4195
R31577 CS_BIAS.n1651 CS_BIAS.t42 15.4195
R31578 CS_BIAS.n1365 CS_BIAS.t92 15.4195
R31579 CS_BIAS.n1387 CS_BIAS.t53 15.4195
R31580 CS_BIAS.n1407 CS_BIAS.t70 15.4195
R31581 CS_BIAS.n1426 CS_BIAS.t68 15.4195
R31582 CS_BIAS.n1339 CS_BIAS.t44 15.4195
R31583 CS_BIAS.n1467 CS_BIAS.t56 15.4195
R31584 CS_BIAS.n1487 CS_BIAS.t71 15.4195
R31585 CS_BIAS.n1201 CS_BIAS.t60 15.4195
R31586 CS_BIAS.n1223 CS_BIAS.t83 15.4195
R31587 CS_BIAS.n1243 CS_BIAS.t40 15.4195
R31588 CS_BIAS.n1262 CS_BIAS.t35 15.4195
R31589 CS_BIAS.n1175 CS_BIAS.t74 15.4195
R31590 CS_BIAS.n1303 CS_BIAS.t89 15.4195
R31591 CS_BIAS.n1323 CS_BIAS.t41 15.4195
R31592 CS_BIAS.n960 CS_BIAS.t26 15.4195
R31593 CS_BIAS.n982 CS_BIAS.t0 15.4195
R31594 CS_BIAS.n1002 CS_BIAS.t10 15.4195
R31595 CS_BIAS.n1021 CS_BIAS.t20 15.4195
R31596 CS_BIAS.n934 CS_BIAS.t4 15.4195
R31597 CS_BIAS.n1062 CS_BIAS.t14 15.4195
R31598 CS_BIAS.n1082 CS_BIAS.t28 15.4195
R31599 CS_BIAS.n1160 CS_BIAS.t58 15.4195
R31600 CS_BIAS.n1140 CS_BIAS.t86 15.4195
R31601 CS_BIAS.n840 CS_BIAS.t46 15.4195
R31602 CS_BIAS.n1099 CS_BIAS.t78 15.4195
R31603 CS_BIAS.n866 CS_BIAS.t63 15.4195
R31604 CS_BIAS.n888 CS_BIAS.t48 15.4195
R31605 CS_BIAS.n908 CS_BIAS.t88 15.4195
R31606 CS_BIAS.n255 CS_BIAS.n253 13.1385
R31607 CS_BIAS.n1085 CS_BIAS.n1083 13.1385
R31608 CS_BIAS.n258 CS_BIAS.t17 10.6171
R31609 CS_BIAS.n258 CS_BIAS.t7 10.6171
R31610 CS_BIAS.n259 CS_BIAS.t9 10.6171
R31611 CS_BIAS.n259 CS_BIAS.t25 10.6171
R31612 CS_BIAS.n256 CS_BIAS.t31 10.6171
R31613 CS_BIAS.n256 CS_BIAS.t19 10.6171
R31614 CS_BIAS.n254 CS_BIAS.t13 10.6171
R31615 CS_BIAS.n254 CS_BIAS.t3 10.6171
R31616 CS_BIAS.n1084 CS_BIAS.t15 10.6171
R31617 CS_BIAS.n1084 CS_BIAS.t29 10.6171
R31618 CS_BIAS.n1086 CS_BIAS.t21 10.6171
R31619 CS_BIAS.n1086 CS_BIAS.t5 10.6171
R31620 CS_BIAS.n919 CS_BIAS.t1 10.6171
R31621 CS_BIAS.n919 CS_BIAS.t11 10.6171
R31622 CS_BIAS.n918 CS_BIAS.t23 10.6171
R31623 CS_BIAS.n918 CS_BIAS.t27 10.6171
R31624 CS_BIAS.n1654 CS_BIAS.n826 10.2112
R31625 CS_BIAS.n262 CS_BIAS.n261 9.503
R31626 CS_BIAS.n1089 CS_BIAS.n1088 9.503
R31627 CS_BIAS.n498 CS_BIAS.n334 8.2452
R31628 CS_BIAS.n1325 CS_BIAS.n1161 8.2452
R31629 CS_BIAS.n1654 CS_BIAS.n1653 7.42944
R31630 CS_BIAS CS_BIAS.n1654 5.99958
R31631 CS_BIAS.n826 CS_BIAS.n825 5.57095
R31632 CS_BIAS.n662 CS_BIAS.n661 5.57095
R31633 CS_BIAS.n498 CS_BIAS.n497 5.57095
R31634 CS_BIAS.n1653 CS_BIAS.n1652 5.57095
R31635 CS_BIAS.n1489 CS_BIAS.n1488 5.57095
R31636 CS_BIAS.n1325 CS_BIAS.n1324 5.57095
R31637 CS_BIAS.n662 CS_BIAS.n498 2.67474
R31638 CS_BIAS.n826 CS_BIAS.n662 2.67474
R31639 CS_BIAS.n1489 CS_BIAS.n1325 2.67474
R31640 CS_BIAS.n1653 CS_BIAS.n1489 2.67474
R31641 CS_BIAS.n257 CS_BIAS.n255 1.86544
R31642 CS_BIAS.n1087 CS_BIAS.n1085 1.86544
R31643 CS_BIAS.n805 CS_BIAS.n804 1.22385
R31644 CS_BIAS.n641 CS_BIAS.n640 1.22385
R31645 CS_BIAS.n477 CS_BIAS.n476 1.22385
R31646 CS_BIAS.n233 CS_BIAS.n232 1.22385
R31647 CS_BIAS.n314 CS_BIAS.n313 1.22385
R31648 CS_BIAS.n1632 CS_BIAS.n1631 1.22385
R31649 CS_BIAS.n1468 CS_BIAS.n1467 1.22385
R31650 CS_BIAS.n1304 CS_BIAS.n1303 1.22385
R31651 CS_BIAS.n1063 CS_BIAS.n1062 1.22385
R31652 CS_BIAS.n1141 CS_BIAS.n1140 1.22385
R31653 CS_BIAS.n261 CS_BIAS.n257 0.932971
R31654 CS_BIAS.n261 CS_BIAS.n260 0.932971
R31655 CS_BIAS.n1088 CS_BIAS.n920 0.932971
R31656 CS_BIAS.n1088 CS_BIAS.n1087 0.932971
R31657 CS_BIAS.n704 CS_BIAS.n703 0.794726
R31658 CS_BIAS.n1531 CS_BIAS.n1530 0.794726
R31659 CS_BIAS.n1367 CS_BIAS.n1366 0.794726
R31660 CS_BIAS.n1203 CS_BIAS.n1202 0.794726
R31661 CS_BIAS.n962 CS_BIAS.n961 0.794726
R31662 CS_BIAS.n868 CS_BIAS.n867 0.794726
R31663 CS_BIAS.n540 CS_BIAS.n539 0.794723
R31664 CS_BIAS.n376 CS_BIAS.n375 0.794723
R31665 CS_BIAS.n132 CS_BIAS.n131 0.794723
R31666 CS_BIAS.n41 CS_BIAS.n40 0.794723
R31667 CS_BIAS.n724 CS_BIAS.n723 0.73451
R31668 CS_BIAS.n785 CS_BIAS.n676 0.73451
R31669 CS_BIAS.n621 CS_BIAS.n512 0.73451
R31670 CS_BIAS.n560 CS_BIAS.n559 0.73451
R31671 CS_BIAS.n457 CS_BIAS.n348 0.73451
R31672 CS_BIAS.n396 CS_BIAS.n395 0.73451
R31673 CS_BIAS.n213 CS_BIAS.n104 0.73451
R31674 CS_BIAS.n152 CS_BIAS.n151 0.73451
R31675 CS_BIAS.n294 CS_BIAS.n13 0.73451
R31676 CS_BIAS.n61 CS_BIAS.n60 0.73451
R31677 CS_BIAS.n1551 CS_BIAS.n1550 0.73451
R31678 CS_BIAS.n1612 CS_BIAS.n1503 0.73451
R31679 CS_BIAS.n1387 CS_BIAS.n1386 0.73451
R31680 CS_BIAS.n1448 CS_BIAS.n1339 0.73451
R31681 CS_BIAS.n1223 CS_BIAS.n1222 0.73451
R31682 CS_BIAS.n1284 CS_BIAS.n1175 0.73451
R31683 CS_BIAS.n982 CS_BIAS.n981 0.73451
R31684 CS_BIAS.n1043 CS_BIAS.n934 0.73451
R31685 CS_BIAS.n1121 CS_BIAS.n840 0.73451
R31686 CS_BIAS.n888 CS_BIAS.n887 0.73451
R31687 CS_BIAS.n825 CS_BIAS.n663 0.502622
R31688 CS_BIAS.n661 CS_BIAS.n499 0.502622
R31689 CS_BIAS.n497 CS_BIAS.n335 0.502622
R31690 CS_BIAS.n253 CS_BIAS.n91 0.502622
R31691 CS_BIAS.n334 CS_BIAS.n0 0.502622
R31692 CS_BIAS.n1652 CS_BIAS.n1490 0.502622
R31693 CS_BIAS.n1488 CS_BIAS.n1326 0.502622
R31694 CS_BIAS.n1324 CS_BIAS.n1162 0.502622
R31695 CS_BIAS.n1083 CS_BIAS.n921 0.502622
R31696 CS_BIAS.n1161 CS_BIAS.n827 0.502622
R31697 CS_BIAS.n744 CS_BIAS.n743 0.24517
R31698 CS_BIAS.n764 CS_BIAS.n763 0.24517
R31699 CS_BIAS.n600 CS_BIAS.n599 0.24517
R31700 CS_BIAS.n580 CS_BIAS.n579 0.24517
R31701 CS_BIAS.n436 CS_BIAS.n435 0.24517
R31702 CS_BIAS.n416 CS_BIAS.n415 0.24517
R31703 CS_BIAS.n192 CS_BIAS.n191 0.24517
R31704 CS_BIAS.n172 CS_BIAS.n171 0.24517
R31705 CS_BIAS.n273 CS_BIAS.n272 0.24517
R31706 CS_BIAS.n81 CS_BIAS.n80 0.24517
R31707 CS_BIAS.n1571 CS_BIAS.n1570 0.24517
R31708 CS_BIAS.n1591 CS_BIAS.n1590 0.24517
R31709 CS_BIAS.n1407 CS_BIAS.n1406 0.24517
R31710 CS_BIAS.n1427 CS_BIAS.n1426 0.24517
R31711 CS_BIAS.n1243 CS_BIAS.n1242 0.24517
R31712 CS_BIAS.n1263 CS_BIAS.n1262 0.24517
R31713 CS_BIAS.n1002 CS_BIAS.n1001 0.24517
R31714 CS_BIAS.n1022 CS_BIAS.n1021 0.24517
R31715 CS_BIAS.n1100 CS_BIAS.n1099 0.24517
R31716 CS_BIAS.n908 CS_BIAS.n907 0.24517
R31717 CS_BIAS.n821 CS_BIAS.n663 0.189894
R31718 CS_BIAS.n821 CS_BIAS.n820 0.189894
R31719 CS_BIAS.n820 CS_BIAS.n819 0.189894
R31720 CS_BIAS.n819 CS_BIAS.n665 0.189894
R31721 CS_BIAS.n815 CS_BIAS.n665 0.189894
R31722 CS_BIAS.n815 CS_BIAS.n814 0.189894
R31723 CS_BIAS.n814 CS_BIAS.n813 0.189894
R31724 CS_BIAS.n813 CS_BIAS.n667 0.189894
R31725 CS_BIAS.n809 CS_BIAS.n667 0.189894
R31726 CS_BIAS.n809 CS_BIAS.n808 0.189894
R31727 CS_BIAS.n808 CS_BIAS.n807 0.189894
R31728 CS_BIAS.n807 CS_BIAS.n669 0.189894
R31729 CS_BIAS.n802 CS_BIAS.n669 0.189894
R31730 CS_BIAS.n802 CS_BIAS.n801 0.189894
R31731 CS_BIAS.n801 CS_BIAS.n800 0.189894
R31732 CS_BIAS.n800 CS_BIAS.n671 0.189894
R31733 CS_BIAS.n796 CS_BIAS.n671 0.189894
R31734 CS_BIAS.n796 CS_BIAS.n795 0.189894
R31735 CS_BIAS.n795 CS_BIAS.n794 0.189894
R31736 CS_BIAS.n794 CS_BIAS.n673 0.189894
R31737 CS_BIAS.n790 CS_BIAS.n673 0.189894
R31738 CS_BIAS.n790 CS_BIAS.n789 0.189894
R31739 CS_BIAS.n789 CS_BIAS.n788 0.189894
R31740 CS_BIAS.n788 CS_BIAS.n675 0.189894
R31741 CS_BIAS.n784 CS_BIAS.n675 0.189894
R31742 CS_BIAS.n784 CS_BIAS.n783 0.189894
R31743 CS_BIAS.n783 CS_BIAS.n677 0.189894
R31744 CS_BIAS.n779 CS_BIAS.n677 0.189894
R31745 CS_BIAS.n779 CS_BIAS.n778 0.189894
R31746 CS_BIAS.n778 CS_BIAS.n777 0.189894
R31747 CS_BIAS.n777 CS_BIAS.n679 0.189894
R31748 CS_BIAS.n773 CS_BIAS.n679 0.189894
R31749 CS_BIAS.n773 CS_BIAS.n772 0.189894
R31750 CS_BIAS.n772 CS_BIAS.n771 0.189894
R31751 CS_BIAS.n771 CS_BIAS.n681 0.189894
R31752 CS_BIAS.n767 CS_BIAS.n681 0.189894
R31753 CS_BIAS.n767 CS_BIAS.n766 0.189894
R31754 CS_BIAS.n766 CS_BIAS.n765 0.189894
R31755 CS_BIAS.n765 CS_BIAS.n683 0.189894
R31756 CS_BIAS.n760 CS_BIAS.n683 0.189894
R31757 CS_BIAS.n760 CS_BIAS.n759 0.189894
R31758 CS_BIAS.n759 CS_BIAS.n758 0.189894
R31759 CS_BIAS.n758 CS_BIAS.n685 0.189894
R31760 CS_BIAS.n754 CS_BIAS.n685 0.189894
R31761 CS_BIAS.n754 CS_BIAS.n753 0.189894
R31762 CS_BIAS.n753 CS_BIAS.n752 0.189894
R31763 CS_BIAS.n752 CS_BIAS.n687 0.189894
R31764 CS_BIAS.n748 CS_BIAS.n687 0.189894
R31765 CS_BIAS.n748 CS_BIAS.n747 0.189894
R31766 CS_BIAS.n747 CS_BIAS.n746 0.189894
R31767 CS_BIAS.n746 CS_BIAS.n689 0.189894
R31768 CS_BIAS.n741 CS_BIAS.n689 0.189894
R31769 CS_BIAS.n741 CS_BIAS.n740 0.189894
R31770 CS_BIAS.n740 CS_BIAS.n739 0.189894
R31771 CS_BIAS.n739 CS_BIAS.n691 0.189894
R31772 CS_BIAS.n735 CS_BIAS.n691 0.189894
R31773 CS_BIAS.n735 CS_BIAS.n734 0.189894
R31774 CS_BIAS.n734 CS_BIAS.n733 0.189894
R31775 CS_BIAS.n733 CS_BIAS.n693 0.189894
R31776 CS_BIAS.n729 CS_BIAS.n693 0.189894
R31777 CS_BIAS.n729 CS_BIAS.n728 0.189894
R31778 CS_BIAS.n728 CS_BIAS.n727 0.189894
R31779 CS_BIAS.n727 CS_BIAS.n695 0.189894
R31780 CS_BIAS.n722 CS_BIAS.n695 0.189894
R31781 CS_BIAS.n722 CS_BIAS.n721 0.189894
R31782 CS_BIAS.n721 CS_BIAS.n720 0.189894
R31783 CS_BIAS.n720 CS_BIAS.n697 0.189894
R31784 CS_BIAS.n716 CS_BIAS.n697 0.189894
R31785 CS_BIAS.n716 CS_BIAS.n715 0.189894
R31786 CS_BIAS.n715 CS_BIAS.n714 0.189894
R31787 CS_BIAS.n714 CS_BIAS.n699 0.189894
R31788 CS_BIAS.n710 CS_BIAS.n699 0.189894
R31789 CS_BIAS.n710 CS_BIAS.n709 0.189894
R31790 CS_BIAS.n709 CS_BIAS.n708 0.189894
R31791 CS_BIAS.n708 CS_BIAS.n701 0.189894
R31792 CS_BIAS.n704 CS_BIAS.n701 0.189894
R31793 CS_BIAS.n657 CS_BIAS.n499 0.189894
R31794 CS_BIAS.n657 CS_BIAS.n656 0.189894
R31795 CS_BIAS.n656 CS_BIAS.n655 0.189894
R31796 CS_BIAS.n655 CS_BIAS.n501 0.189894
R31797 CS_BIAS.n651 CS_BIAS.n501 0.189894
R31798 CS_BIAS.n651 CS_BIAS.n650 0.189894
R31799 CS_BIAS.n650 CS_BIAS.n649 0.189894
R31800 CS_BIAS.n649 CS_BIAS.n503 0.189894
R31801 CS_BIAS.n645 CS_BIAS.n503 0.189894
R31802 CS_BIAS.n645 CS_BIAS.n644 0.189894
R31803 CS_BIAS.n644 CS_BIAS.n643 0.189894
R31804 CS_BIAS.n643 CS_BIAS.n505 0.189894
R31805 CS_BIAS.n638 CS_BIAS.n505 0.189894
R31806 CS_BIAS.n638 CS_BIAS.n637 0.189894
R31807 CS_BIAS.n637 CS_BIAS.n636 0.189894
R31808 CS_BIAS.n636 CS_BIAS.n507 0.189894
R31809 CS_BIAS.n632 CS_BIAS.n507 0.189894
R31810 CS_BIAS.n632 CS_BIAS.n631 0.189894
R31811 CS_BIAS.n631 CS_BIAS.n630 0.189894
R31812 CS_BIAS.n630 CS_BIAS.n509 0.189894
R31813 CS_BIAS.n626 CS_BIAS.n509 0.189894
R31814 CS_BIAS.n626 CS_BIAS.n625 0.189894
R31815 CS_BIAS.n625 CS_BIAS.n624 0.189894
R31816 CS_BIAS.n624 CS_BIAS.n511 0.189894
R31817 CS_BIAS.n620 CS_BIAS.n511 0.189894
R31818 CS_BIAS.n620 CS_BIAS.n619 0.189894
R31819 CS_BIAS.n619 CS_BIAS.n513 0.189894
R31820 CS_BIAS.n615 CS_BIAS.n513 0.189894
R31821 CS_BIAS.n615 CS_BIAS.n614 0.189894
R31822 CS_BIAS.n614 CS_BIAS.n613 0.189894
R31823 CS_BIAS.n613 CS_BIAS.n515 0.189894
R31824 CS_BIAS.n609 CS_BIAS.n515 0.189894
R31825 CS_BIAS.n609 CS_BIAS.n608 0.189894
R31826 CS_BIAS.n608 CS_BIAS.n607 0.189894
R31827 CS_BIAS.n607 CS_BIAS.n517 0.189894
R31828 CS_BIAS.n603 CS_BIAS.n517 0.189894
R31829 CS_BIAS.n603 CS_BIAS.n602 0.189894
R31830 CS_BIAS.n602 CS_BIAS.n601 0.189894
R31831 CS_BIAS.n601 CS_BIAS.n519 0.189894
R31832 CS_BIAS.n596 CS_BIAS.n519 0.189894
R31833 CS_BIAS.n596 CS_BIAS.n595 0.189894
R31834 CS_BIAS.n595 CS_BIAS.n594 0.189894
R31835 CS_BIAS.n594 CS_BIAS.n521 0.189894
R31836 CS_BIAS.n590 CS_BIAS.n521 0.189894
R31837 CS_BIAS.n590 CS_BIAS.n589 0.189894
R31838 CS_BIAS.n589 CS_BIAS.n588 0.189894
R31839 CS_BIAS.n588 CS_BIAS.n523 0.189894
R31840 CS_BIAS.n584 CS_BIAS.n523 0.189894
R31841 CS_BIAS.n584 CS_BIAS.n583 0.189894
R31842 CS_BIAS.n583 CS_BIAS.n582 0.189894
R31843 CS_BIAS.n582 CS_BIAS.n525 0.189894
R31844 CS_BIAS.n577 CS_BIAS.n525 0.189894
R31845 CS_BIAS.n577 CS_BIAS.n576 0.189894
R31846 CS_BIAS.n576 CS_BIAS.n575 0.189894
R31847 CS_BIAS.n575 CS_BIAS.n527 0.189894
R31848 CS_BIAS.n571 CS_BIAS.n527 0.189894
R31849 CS_BIAS.n571 CS_BIAS.n570 0.189894
R31850 CS_BIAS.n570 CS_BIAS.n569 0.189894
R31851 CS_BIAS.n569 CS_BIAS.n529 0.189894
R31852 CS_BIAS.n565 CS_BIAS.n529 0.189894
R31853 CS_BIAS.n565 CS_BIAS.n564 0.189894
R31854 CS_BIAS.n564 CS_BIAS.n563 0.189894
R31855 CS_BIAS.n563 CS_BIAS.n531 0.189894
R31856 CS_BIAS.n558 CS_BIAS.n531 0.189894
R31857 CS_BIAS.n558 CS_BIAS.n557 0.189894
R31858 CS_BIAS.n557 CS_BIAS.n556 0.189894
R31859 CS_BIAS.n556 CS_BIAS.n533 0.189894
R31860 CS_BIAS.n552 CS_BIAS.n533 0.189894
R31861 CS_BIAS.n552 CS_BIAS.n551 0.189894
R31862 CS_BIAS.n551 CS_BIAS.n550 0.189894
R31863 CS_BIAS.n550 CS_BIAS.n535 0.189894
R31864 CS_BIAS.n546 CS_BIAS.n535 0.189894
R31865 CS_BIAS.n546 CS_BIAS.n545 0.189894
R31866 CS_BIAS.n545 CS_BIAS.n544 0.189894
R31867 CS_BIAS.n544 CS_BIAS.n537 0.189894
R31868 CS_BIAS.n540 CS_BIAS.n537 0.189894
R31869 CS_BIAS.n493 CS_BIAS.n335 0.189894
R31870 CS_BIAS.n493 CS_BIAS.n492 0.189894
R31871 CS_BIAS.n492 CS_BIAS.n491 0.189894
R31872 CS_BIAS.n491 CS_BIAS.n337 0.189894
R31873 CS_BIAS.n487 CS_BIAS.n337 0.189894
R31874 CS_BIAS.n487 CS_BIAS.n486 0.189894
R31875 CS_BIAS.n486 CS_BIAS.n485 0.189894
R31876 CS_BIAS.n485 CS_BIAS.n339 0.189894
R31877 CS_BIAS.n481 CS_BIAS.n339 0.189894
R31878 CS_BIAS.n481 CS_BIAS.n480 0.189894
R31879 CS_BIAS.n480 CS_BIAS.n479 0.189894
R31880 CS_BIAS.n479 CS_BIAS.n341 0.189894
R31881 CS_BIAS.n474 CS_BIAS.n341 0.189894
R31882 CS_BIAS.n474 CS_BIAS.n473 0.189894
R31883 CS_BIAS.n473 CS_BIAS.n472 0.189894
R31884 CS_BIAS.n472 CS_BIAS.n343 0.189894
R31885 CS_BIAS.n468 CS_BIAS.n343 0.189894
R31886 CS_BIAS.n468 CS_BIAS.n467 0.189894
R31887 CS_BIAS.n467 CS_BIAS.n466 0.189894
R31888 CS_BIAS.n466 CS_BIAS.n345 0.189894
R31889 CS_BIAS.n462 CS_BIAS.n345 0.189894
R31890 CS_BIAS.n462 CS_BIAS.n461 0.189894
R31891 CS_BIAS.n461 CS_BIAS.n460 0.189894
R31892 CS_BIAS.n460 CS_BIAS.n347 0.189894
R31893 CS_BIAS.n456 CS_BIAS.n347 0.189894
R31894 CS_BIAS.n456 CS_BIAS.n455 0.189894
R31895 CS_BIAS.n455 CS_BIAS.n349 0.189894
R31896 CS_BIAS.n451 CS_BIAS.n349 0.189894
R31897 CS_BIAS.n451 CS_BIAS.n450 0.189894
R31898 CS_BIAS.n450 CS_BIAS.n449 0.189894
R31899 CS_BIAS.n449 CS_BIAS.n351 0.189894
R31900 CS_BIAS.n445 CS_BIAS.n351 0.189894
R31901 CS_BIAS.n445 CS_BIAS.n444 0.189894
R31902 CS_BIAS.n444 CS_BIAS.n443 0.189894
R31903 CS_BIAS.n443 CS_BIAS.n353 0.189894
R31904 CS_BIAS.n439 CS_BIAS.n353 0.189894
R31905 CS_BIAS.n439 CS_BIAS.n438 0.189894
R31906 CS_BIAS.n438 CS_BIAS.n437 0.189894
R31907 CS_BIAS.n437 CS_BIAS.n355 0.189894
R31908 CS_BIAS.n432 CS_BIAS.n355 0.189894
R31909 CS_BIAS.n432 CS_BIAS.n431 0.189894
R31910 CS_BIAS.n431 CS_BIAS.n430 0.189894
R31911 CS_BIAS.n430 CS_BIAS.n357 0.189894
R31912 CS_BIAS.n426 CS_BIAS.n357 0.189894
R31913 CS_BIAS.n426 CS_BIAS.n425 0.189894
R31914 CS_BIAS.n425 CS_BIAS.n424 0.189894
R31915 CS_BIAS.n424 CS_BIAS.n359 0.189894
R31916 CS_BIAS.n420 CS_BIAS.n359 0.189894
R31917 CS_BIAS.n420 CS_BIAS.n419 0.189894
R31918 CS_BIAS.n419 CS_BIAS.n418 0.189894
R31919 CS_BIAS.n418 CS_BIAS.n361 0.189894
R31920 CS_BIAS.n413 CS_BIAS.n361 0.189894
R31921 CS_BIAS.n413 CS_BIAS.n412 0.189894
R31922 CS_BIAS.n412 CS_BIAS.n411 0.189894
R31923 CS_BIAS.n411 CS_BIAS.n363 0.189894
R31924 CS_BIAS.n407 CS_BIAS.n363 0.189894
R31925 CS_BIAS.n407 CS_BIAS.n406 0.189894
R31926 CS_BIAS.n406 CS_BIAS.n405 0.189894
R31927 CS_BIAS.n405 CS_BIAS.n365 0.189894
R31928 CS_BIAS.n401 CS_BIAS.n365 0.189894
R31929 CS_BIAS.n401 CS_BIAS.n400 0.189894
R31930 CS_BIAS.n400 CS_BIAS.n399 0.189894
R31931 CS_BIAS.n399 CS_BIAS.n367 0.189894
R31932 CS_BIAS.n394 CS_BIAS.n367 0.189894
R31933 CS_BIAS.n394 CS_BIAS.n393 0.189894
R31934 CS_BIAS.n393 CS_BIAS.n392 0.189894
R31935 CS_BIAS.n392 CS_BIAS.n369 0.189894
R31936 CS_BIAS.n388 CS_BIAS.n369 0.189894
R31937 CS_BIAS.n388 CS_BIAS.n387 0.189894
R31938 CS_BIAS.n387 CS_BIAS.n386 0.189894
R31939 CS_BIAS.n386 CS_BIAS.n371 0.189894
R31940 CS_BIAS.n382 CS_BIAS.n371 0.189894
R31941 CS_BIAS.n382 CS_BIAS.n381 0.189894
R31942 CS_BIAS.n381 CS_BIAS.n380 0.189894
R31943 CS_BIAS.n380 CS_BIAS.n373 0.189894
R31944 CS_BIAS.n376 CS_BIAS.n373 0.189894
R31945 CS_BIAS.n249 CS_BIAS.n91 0.189894
R31946 CS_BIAS.n249 CS_BIAS.n248 0.189894
R31947 CS_BIAS.n248 CS_BIAS.n247 0.189894
R31948 CS_BIAS.n247 CS_BIAS.n93 0.189894
R31949 CS_BIAS.n243 CS_BIAS.n93 0.189894
R31950 CS_BIAS.n243 CS_BIAS.n242 0.189894
R31951 CS_BIAS.n242 CS_BIAS.n241 0.189894
R31952 CS_BIAS.n241 CS_BIAS.n95 0.189894
R31953 CS_BIAS.n237 CS_BIAS.n95 0.189894
R31954 CS_BIAS.n237 CS_BIAS.n236 0.189894
R31955 CS_BIAS.n236 CS_BIAS.n235 0.189894
R31956 CS_BIAS.n235 CS_BIAS.n97 0.189894
R31957 CS_BIAS.n230 CS_BIAS.n97 0.189894
R31958 CS_BIAS.n230 CS_BIAS.n229 0.189894
R31959 CS_BIAS.n229 CS_BIAS.n228 0.189894
R31960 CS_BIAS.n228 CS_BIAS.n99 0.189894
R31961 CS_BIAS.n224 CS_BIAS.n99 0.189894
R31962 CS_BIAS.n224 CS_BIAS.n223 0.189894
R31963 CS_BIAS.n223 CS_BIAS.n222 0.189894
R31964 CS_BIAS.n222 CS_BIAS.n101 0.189894
R31965 CS_BIAS.n218 CS_BIAS.n101 0.189894
R31966 CS_BIAS.n218 CS_BIAS.n217 0.189894
R31967 CS_BIAS.n217 CS_BIAS.n216 0.189894
R31968 CS_BIAS.n216 CS_BIAS.n103 0.189894
R31969 CS_BIAS.n212 CS_BIAS.n103 0.189894
R31970 CS_BIAS.n212 CS_BIAS.n211 0.189894
R31971 CS_BIAS.n211 CS_BIAS.n105 0.189894
R31972 CS_BIAS.n207 CS_BIAS.n105 0.189894
R31973 CS_BIAS.n207 CS_BIAS.n206 0.189894
R31974 CS_BIAS.n206 CS_BIAS.n205 0.189894
R31975 CS_BIAS.n205 CS_BIAS.n107 0.189894
R31976 CS_BIAS.n201 CS_BIAS.n107 0.189894
R31977 CS_BIAS.n201 CS_BIAS.n200 0.189894
R31978 CS_BIAS.n200 CS_BIAS.n199 0.189894
R31979 CS_BIAS.n199 CS_BIAS.n109 0.189894
R31980 CS_BIAS.n195 CS_BIAS.n109 0.189894
R31981 CS_BIAS.n195 CS_BIAS.n194 0.189894
R31982 CS_BIAS.n194 CS_BIAS.n193 0.189894
R31983 CS_BIAS.n193 CS_BIAS.n111 0.189894
R31984 CS_BIAS.n188 CS_BIAS.n111 0.189894
R31985 CS_BIAS.n188 CS_BIAS.n187 0.189894
R31986 CS_BIAS.n187 CS_BIAS.n186 0.189894
R31987 CS_BIAS.n186 CS_BIAS.n113 0.189894
R31988 CS_BIAS.n182 CS_BIAS.n113 0.189894
R31989 CS_BIAS.n182 CS_BIAS.n181 0.189894
R31990 CS_BIAS.n181 CS_BIAS.n180 0.189894
R31991 CS_BIAS.n180 CS_BIAS.n115 0.189894
R31992 CS_BIAS.n176 CS_BIAS.n115 0.189894
R31993 CS_BIAS.n176 CS_BIAS.n175 0.189894
R31994 CS_BIAS.n175 CS_BIAS.n174 0.189894
R31995 CS_BIAS.n174 CS_BIAS.n117 0.189894
R31996 CS_BIAS.n169 CS_BIAS.n117 0.189894
R31997 CS_BIAS.n169 CS_BIAS.n168 0.189894
R31998 CS_BIAS.n168 CS_BIAS.n167 0.189894
R31999 CS_BIAS.n167 CS_BIAS.n119 0.189894
R32000 CS_BIAS.n163 CS_BIAS.n119 0.189894
R32001 CS_BIAS.n163 CS_BIAS.n162 0.189894
R32002 CS_BIAS.n162 CS_BIAS.n161 0.189894
R32003 CS_BIAS.n161 CS_BIAS.n121 0.189894
R32004 CS_BIAS.n157 CS_BIAS.n121 0.189894
R32005 CS_BIAS.n157 CS_BIAS.n156 0.189894
R32006 CS_BIAS.n156 CS_BIAS.n155 0.189894
R32007 CS_BIAS.n155 CS_BIAS.n123 0.189894
R32008 CS_BIAS.n150 CS_BIAS.n123 0.189894
R32009 CS_BIAS.n150 CS_BIAS.n149 0.189894
R32010 CS_BIAS.n149 CS_BIAS.n148 0.189894
R32011 CS_BIAS.n148 CS_BIAS.n125 0.189894
R32012 CS_BIAS.n144 CS_BIAS.n125 0.189894
R32013 CS_BIAS.n144 CS_BIAS.n143 0.189894
R32014 CS_BIAS.n143 CS_BIAS.n142 0.189894
R32015 CS_BIAS.n142 CS_BIAS.n127 0.189894
R32016 CS_BIAS.n138 CS_BIAS.n127 0.189894
R32017 CS_BIAS.n138 CS_BIAS.n137 0.189894
R32018 CS_BIAS.n137 CS_BIAS.n136 0.189894
R32019 CS_BIAS.n136 CS_BIAS.n129 0.189894
R32020 CS_BIAS.n132 CS_BIAS.n129 0.189894
R32021 CS_BIAS.n90 CS_BIAS.n89 0.189894
R32022 CS_BIAS.n89 CS_BIAS.n24 0.189894
R32023 CS_BIAS.n85 CS_BIAS.n24 0.189894
R32024 CS_BIAS.n85 CS_BIAS.n84 0.189894
R32025 CS_BIAS.n84 CS_BIAS.n83 0.189894
R32026 CS_BIAS.n83 CS_BIAS.n26 0.189894
R32027 CS_BIAS.n78 CS_BIAS.n26 0.189894
R32028 CS_BIAS.n78 CS_BIAS.n77 0.189894
R32029 CS_BIAS.n77 CS_BIAS.n76 0.189894
R32030 CS_BIAS.n76 CS_BIAS.n28 0.189894
R32031 CS_BIAS.n72 CS_BIAS.n28 0.189894
R32032 CS_BIAS.n72 CS_BIAS.n71 0.189894
R32033 CS_BIAS.n71 CS_BIAS.n70 0.189894
R32034 CS_BIAS.n70 CS_BIAS.n30 0.189894
R32035 CS_BIAS.n66 CS_BIAS.n30 0.189894
R32036 CS_BIAS.n66 CS_BIAS.n65 0.189894
R32037 CS_BIAS.n65 CS_BIAS.n64 0.189894
R32038 CS_BIAS.n64 CS_BIAS.n32 0.189894
R32039 CS_BIAS.n59 CS_BIAS.n32 0.189894
R32040 CS_BIAS.n59 CS_BIAS.n58 0.189894
R32041 CS_BIAS.n58 CS_BIAS.n57 0.189894
R32042 CS_BIAS.n57 CS_BIAS.n34 0.189894
R32043 CS_BIAS.n53 CS_BIAS.n34 0.189894
R32044 CS_BIAS.n53 CS_BIAS.n52 0.189894
R32045 CS_BIAS.n52 CS_BIAS.n51 0.189894
R32046 CS_BIAS.n51 CS_BIAS.n36 0.189894
R32047 CS_BIAS.n47 CS_BIAS.n36 0.189894
R32048 CS_BIAS.n47 CS_BIAS.n46 0.189894
R32049 CS_BIAS.n46 CS_BIAS.n45 0.189894
R32050 CS_BIAS.n45 CS_BIAS.n38 0.189894
R32051 CS_BIAS.n41 CS_BIAS.n38 0.189894
R32052 CS_BIAS.n330 CS_BIAS.n0 0.189894
R32053 CS_BIAS.n330 CS_BIAS.n329 0.189894
R32054 CS_BIAS.n329 CS_BIAS.n328 0.189894
R32055 CS_BIAS.n328 CS_BIAS.n2 0.189894
R32056 CS_BIAS.n324 CS_BIAS.n2 0.189894
R32057 CS_BIAS.n324 CS_BIAS.n323 0.189894
R32058 CS_BIAS.n323 CS_BIAS.n322 0.189894
R32059 CS_BIAS.n322 CS_BIAS.n4 0.189894
R32060 CS_BIAS.n318 CS_BIAS.n4 0.189894
R32061 CS_BIAS.n318 CS_BIAS.n317 0.189894
R32062 CS_BIAS.n317 CS_BIAS.n316 0.189894
R32063 CS_BIAS.n316 CS_BIAS.n6 0.189894
R32064 CS_BIAS.n311 CS_BIAS.n6 0.189894
R32065 CS_BIAS.n311 CS_BIAS.n310 0.189894
R32066 CS_BIAS.n310 CS_BIAS.n309 0.189894
R32067 CS_BIAS.n309 CS_BIAS.n8 0.189894
R32068 CS_BIAS.n305 CS_BIAS.n8 0.189894
R32069 CS_BIAS.n305 CS_BIAS.n304 0.189894
R32070 CS_BIAS.n304 CS_BIAS.n303 0.189894
R32071 CS_BIAS.n303 CS_BIAS.n10 0.189894
R32072 CS_BIAS.n299 CS_BIAS.n10 0.189894
R32073 CS_BIAS.n299 CS_BIAS.n298 0.189894
R32074 CS_BIAS.n298 CS_BIAS.n297 0.189894
R32075 CS_BIAS.n297 CS_BIAS.n12 0.189894
R32076 CS_BIAS.n293 CS_BIAS.n12 0.189894
R32077 CS_BIAS.n293 CS_BIAS.n292 0.189894
R32078 CS_BIAS.n292 CS_BIAS.n14 0.189894
R32079 CS_BIAS.n288 CS_BIAS.n14 0.189894
R32080 CS_BIAS.n288 CS_BIAS.n287 0.189894
R32081 CS_BIAS.n287 CS_BIAS.n286 0.189894
R32082 CS_BIAS.n286 CS_BIAS.n16 0.189894
R32083 CS_BIAS.n282 CS_BIAS.n16 0.189894
R32084 CS_BIAS.n282 CS_BIAS.n281 0.189894
R32085 CS_BIAS.n281 CS_BIAS.n280 0.189894
R32086 CS_BIAS.n280 CS_BIAS.n18 0.189894
R32087 CS_BIAS.n276 CS_BIAS.n18 0.189894
R32088 CS_BIAS.n276 CS_BIAS.n275 0.189894
R32089 CS_BIAS.n275 CS_BIAS.n274 0.189894
R32090 CS_BIAS.n274 CS_BIAS.n20 0.189894
R32091 CS_BIAS.n269 CS_BIAS.n20 0.189894
R32092 CS_BIAS.n269 CS_BIAS.n268 0.189894
R32093 CS_BIAS.n268 CS_BIAS.n267 0.189894
R32094 CS_BIAS.n267 CS_BIAS.n22 0.189894
R32095 CS_BIAS.n263 CS_BIAS.n22 0.189894
R32096 CS_BIAS.n1531 CS_BIAS.n1528 0.189894
R32097 CS_BIAS.n1535 CS_BIAS.n1528 0.189894
R32098 CS_BIAS.n1536 CS_BIAS.n1535 0.189894
R32099 CS_BIAS.n1537 CS_BIAS.n1536 0.189894
R32100 CS_BIAS.n1537 CS_BIAS.n1526 0.189894
R32101 CS_BIAS.n1541 CS_BIAS.n1526 0.189894
R32102 CS_BIAS.n1542 CS_BIAS.n1541 0.189894
R32103 CS_BIAS.n1543 CS_BIAS.n1542 0.189894
R32104 CS_BIAS.n1543 CS_BIAS.n1524 0.189894
R32105 CS_BIAS.n1547 CS_BIAS.n1524 0.189894
R32106 CS_BIAS.n1548 CS_BIAS.n1547 0.189894
R32107 CS_BIAS.n1549 CS_BIAS.n1548 0.189894
R32108 CS_BIAS.n1549 CS_BIAS.n1522 0.189894
R32109 CS_BIAS.n1554 CS_BIAS.n1522 0.189894
R32110 CS_BIAS.n1555 CS_BIAS.n1554 0.189894
R32111 CS_BIAS.n1556 CS_BIAS.n1555 0.189894
R32112 CS_BIAS.n1556 CS_BIAS.n1520 0.189894
R32113 CS_BIAS.n1560 CS_BIAS.n1520 0.189894
R32114 CS_BIAS.n1561 CS_BIAS.n1560 0.189894
R32115 CS_BIAS.n1562 CS_BIAS.n1561 0.189894
R32116 CS_BIAS.n1562 CS_BIAS.n1518 0.189894
R32117 CS_BIAS.n1566 CS_BIAS.n1518 0.189894
R32118 CS_BIAS.n1567 CS_BIAS.n1566 0.189894
R32119 CS_BIAS.n1568 CS_BIAS.n1567 0.189894
R32120 CS_BIAS.n1568 CS_BIAS.n1516 0.189894
R32121 CS_BIAS.n1573 CS_BIAS.n1516 0.189894
R32122 CS_BIAS.n1574 CS_BIAS.n1573 0.189894
R32123 CS_BIAS.n1575 CS_BIAS.n1574 0.189894
R32124 CS_BIAS.n1575 CS_BIAS.n1514 0.189894
R32125 CS_BIAS.n1579 CS_BIAS.n1514 0.189894
R32126 CS_BIAS.n1580 CS_BIAS.n1579 0.189894
R32127 CS_BIAS.n1581 CS_BIAS.n1580 0.189894
R32128 CS_BIAS.n1581 CS_BIAS.n1512 0.189894
R32129 CS_BIAS.n1585 CS_BIAS.n1512 0.189894
R32130 CS_BIAS.n1586 CS_BIAS.n1585 0.189894
R32131 CS_BIAS.n1587 CS_BIAS.n1586 0.189894
R32132 CS_BIAS.n1587 CS_BIAS.n1510 0.189894
R32133 CS_BIAS.n1592 CS_BIAS.n1510 0.189894
R32134 CS_BIAS.n1593 CS_BIAS.n1592 0.189894
R32135 CS_BIAS.n1594 CS_BIAS.n1593 0.189894
R32136 CS_BIAS.n1594 CS_BIAS.n1508 0.189894
R32137 CS_BIAS.n1598 CS_BIAS.n1508 0.189894
R32138 CS_BIAS.n1599 CS_BIAS.n1598 0.189894
R32139 CS_BIAS.n1600 CS_BIAS.n1599 0.189894
R32140 CS_BIAS.n1600 CS_BIAS.n1506 0.189894
R32141 CS_BIAS.n1604 CS_BIAS.n1506 0.189894
R32142 CS_BIAS.n1605 CS_BIAS.n1604 0.189894
R32143 CS_BIAS.n1606 CS_BIAS.n1605 0.189894
R32144 CS_BIAS.n1606 CS_BIAS.n1504 0.189894
R32145 CS_BIAS.n1610 CS_BIAS.n1504 0.189894
R32146 CS_BIAS.n1611 CS_BIAS.n1610 0.189894
R32147 CS_BIAS.n1611 CS_BIAS.n1502 0.189894
R32148 CS_BIAS.n1615 CS_BIAS.n1502 0.189894
R32149 CS_BIAS.n1616 CS_BIAS.n1615 0.189894
R32150 CS_BIAS.n1617 CS_BIAS.n1616 0.189894
R32151 CS_BIAS.n1617 CS_BIAS.n1500 0.189894
R32152 CS_BIAS.n1621 CS_BIAS.n1500 0.189894
R32153 CS_BIAS.n1622 CS_BIAS.n1621 0.189894
R32154 CS_BIAS.n1623 CS_BIAS.n1622 0.189894
R32155 CS_BIAS.n1623 CS_BIAS.n1498 0.189894
R32156 CS_BIAS.n1627 CS_BIAS.n1498 0.189894
R32157 CS_BIAS.n1628 CS_BIAS.n1627 0.189894
R32158 CS_BIAS.n1629 CS_BIAS.n1628 0.189894
R32159 CS_BIAS.n1629 CS_BIAS.n1496 0.189894
R32160 CS_BIAS.n1634 CS_BIAS.n1496 0.189894
R32161 CS_BIAS.n1635 CS_BIAS.n1634 0.189894
R32162 CS_BIAS.n1636 CS_BIAS.n1635 0.189894
R32163 CS_BIAS.n1636 CS_BIAS.n1494 0.189894
R32164 CS_BIAS.n1640 CS_BIAS.n1494 0.189894
R32165 CS_BIAS.n1641 CS_BIAS.n1640 0.189894
R32166 CS_BIAS.n1642 CS_BIAS.n1641 0.189894
R32167 CS_BIAS.n1642 CS_BIAS.n1492 0.189894
R32168 CS_BIAS.n1646 CS_BIAS.n1492 0.189894
R32169 CS_BIAS.n1647 CS_BIAS.n1646 0.189894
R32170 CS_BIAS.n1648 CS_BIAS.n1647 0.189894
R32171 CS_BIAS.n1648 CS_BIAS.n1490 0.189894
R32172 CS_BIAS.n1367 CS_BIAS.n1364 0.189894
R32173 CS_BIAS.n1371 CS_BIAS.n1364 0.189894
R32174 CS_BIAS.n1372 CS_BIAS.n1371 0.189894
R32175 CS_BIAS.n1373 CS_BIAS.n1372 0.189894
R32176 CS_BIAS.n1373 CS_BIAS.n1362 0.189894
R32177 CS_BIAS.n1377 CS_BIAS.n1362 0.189894
R32178 CS_BIAS.n1378 CS_BIAS.n1377 0.189894
R32179 CS_BIAS.n1379 CS_BIAS.n1378 0.189894
R32180 CS_BIAS.n1379 CS_BIAS.n1360 0.189894
R32181 CS_BIAS.n1383 CS_BIAS.n1360 0.189894
R32182 CS_BIAS.n1384 CS_BIAS.n1383 0.189894
R32183 CS_BIAS.n1385 CS_BIAS.n1384 0.189894
R32184 CS_BIAS.n1385 CS_BIAS.n1358 0.189894
R32185 CS_BIAS.n1390 CS_BIAS.n1358 0.189894
R32186 CS_BIAS.n1391 CS_BIAS.n1390 0.189894
R32187 CS_BIAS.n1392 CS_BIAS.n1391 0.189894
R32188 CS_BIAS.n1392 CS_BIAS.n1356 0.189894
R32189 CS_BIAS.n1396 CS_BIAS.n1356 0.189894
R32190 CS_BIAS.n1397 CS_BIAS.n1396 0.189894
R32191 CS_BIAS.n1398 CS_BIAS.n1397 0.189894
R32192 CS_BIAS.n1398 CS_BIAS.n1354 0.189894
R32193 CS_BIAS.n1402 CS_BIAS.n1354 0.189894
R32194 CS_BIAS.n1403 CS_BIAS.n1402 0.189894
R32195 CS_BIAS.n1404 CS_BIAS.n1403 0.189894
R32196 CS_BIAS.n1404 CS_BIAS.n1352 0.189894
R32197 CS_BIAS.n1409 CS_BIAS.n1352 0.189894
R32198 CS_BIAS.n1410 CS_BIAS.n1409 0.189894
R32199 CS_BIAS.n1411 CS_BIAS.n1410 0.189894
R32200 CS_BIAS.n1411 CS_BIAS.n1350 0.189894
R32201 CS_BIAS.n1415 CS_BIAS.n1350 0.189894
R32202 CS_BIAS.n1416 CS_BIAS.n1415 0.189894
R32203 CS_BIAS.n1417 CS_BIAS.n1416 0.189894
R32204 CS_BIAS.n1417 CS_BIAS.n1348 0.189894
R32205 CS_BIAS.n1421 CS_BIAS.n1348 0.189894
R32206 CS_BIAS.n1422 CS_BIAS.n1421 0.189894
R32207 CS_BIAS.n1423 CS_BIAS.n1422 0.189894
R32208 CS_BIAS.n1423 CS_BIAS.n1346 0.189894
R32209 CS_BIAS.n1428 CS_BIAS.n1346 0.189894
R32210 CS_BIAS.n1429 CS_BIAS.n1428 0.189894
R32211 CS_BIAS.n1430 CS_BIAS.n1429 0.189894
R32212 CS_BIAS.n1430 CS_BIAS.n1344 0.189894
R32213 CS_BIAS.n1434 CS_BIAS.n1344 0.189894
R32214 CS_BIAS.n1435 CS_BIAS.n1434 0.189894
R32215 CS_BIAS.n1436 CS_BIAS.n1435 0.189894
R32216 CS_BIAS.n1436 CS_BIAS.n1342 0.189894
R32217 CS_BIAS.n1440 CS_BIAS.n1342 0.189894
R32218 CS_BIAS.n1441 CS_BIAS.n1440 0.189894
R32219 CS_BIAS.n1442 CS_BIAS.n1441 0.189894
R32220 CS_BIAS.n1442 CS_BIAS.n1340 0.189894
R32221 CS_BIAS.n1446 CS_BIAS.n1340 0.189894
R32222 CS_BIAS.n1447 CS_BIAS.n1446 0.189894
R32223 CS_BIAS.n1447 CS_BIAS.n1338 0.189894
R32224 CS_BIAS.n1451 CS_BIAS.n1338 0.189894
R32225 CS_BIAS.n1452 CS_BIAS.n1451 0.189894
R32226 CS_BIAS.n1453 CS_BIAS.n1452 0.189894
R32227 CS_BIAS.n1453 CS_BIAS.n1336 0.189894
R32228 CS_BIAS.n1457 CS_BIAS.n1336 0.189894
R32229 CS_BIAS.n1458 CS_BIAS.n1457 0.189894
R32230 CS_BIAS.n1459 CS_BIAS.n1458 0.189894
R32231 CS_BIAS.n1459 CS_BIAS.n1334 0.189894
R32232 CS_BIAS.n1463 CS_BIAS.n1334 0.189894
R32233 CS_BIAS.n1464 CS_BIAS.n1463 0.189894
R32234 CS_BIAS.n1465 CS_BIAS.n1464 0.189894
R32235 CS_BIAS.n1465 CS_BIAS.n1332 0.189894
R32236 CS_BIAS.n1470 CS_BIAS.n1332 0.189894
R32237 CS_BIAS.n1471 CS_BIAS.n1470 0.189894
R32238 CS_BIAS.n1472 CS_BIAS.n1471 0.189894
R32239 CS_BIAS.n1472 CS_BIAS.n1330 0.189894
R32240 CS_BIAS.n1476 CS_BIAS.n1330 0.189894
R32241 CS_BIAS.n1477 CS_BIAS.n1476 0.189894
R32242 CS_BIAS.n1478 CS_BIAS.n1477 0.189894
R32243 CS_BIAS.n1478 CS_BIAS.n1328 0.189894
R32244 CS_BIAS.n1482 CS_BIAS.n1328 0.189894
R32245 CS_BIAS.n1483 CS_BIAS.n1482 0.189894
R32246 CS_BIAS.n1484 CS_BIAS.n1483 0.189894
R32247 CS_BIAS.n1484 CS_BIAS.n1326 0.189894
R32248 CS_BIAS.n1203 CS_BIAS.n1200 0.189894
R32249 CS_BIAS.n1207 CS_BIAS.n1200 0.189894
R32250 CS_BIAS.n1208 CS_BIAS.n1207 0.189894
R32251 CS_BIAS.n1209 CS_BIAS.n1208 0.189894
R32252 CS_BIAS.n1209 CS_BIAS.n1198 0.189894
R32253 CS_BIAS.n1213 CS_BIAS.n1198 0.189894
R32254 CS_BIAS.n1214 CS_BIAS.n1213 0.189894
R32255 CS_BIAS.n1215 CS_BIAS.n1214 0.189894
R32256 CS_BIAS.n1215 CS_BIAS.n1196 0.189894
R32257 CS_BIAS.n1219 CS_BIAS.n1196 0.189894
R32258 CS_BIAS.n1220 CS_BIAS.n1219 0.189894
R32259 CS_BIAS.n1221 CS_BIAS.n1220 0.189894
R32260 CS_BIAS.n1221 CS_BIAS.n1194 0.189894
R32261 CS_BIAS.n1226 CS_BIAS.n1194 0.189894
R32262 CS_BIAS.n1227 CS_BIAS.n1226 0.189894
R32263 CS_BIAS.n1228 CS_BIAS.n1227 0.189894
R32264 CS_BIAS.n1228 CS_BIAS.n1192 0.189894
R32265 CS_BIAS.n1232 CS_BIAS.n1192 0.189894
R32266 CS_BIAS.n1233 CS_BIAS.n1232 0.189894
R32267 CS_BIAS.n1234 CS_BIAS.n1233 0.189894
R32268 CS_BIAS.n1234 CS_BIAS.n1190 0.189894
R32269 CS_BIAS.n1238 CS_BIAS.n1190 0.189894
R32270 CS_BIAS.n1239 CS_BIAS.n1238 0.189894
R32271 CS_BIAS.n1240 CS_BIAS.n1239 0.189894
R32272 CS_BIAS.n1240 CS_BIAS.n1188 0.189894
R32273 CS_BIAS.n1245 CS_BIAS.n1188 0.189894
R32274 CS_BIAS.n1246 CS_BIAS.n1245 0.189894
R32275 CS_BIAS.n1247 CS_BIAS.n1246 0.189894
R32276 CS_BIAS.n1247 CS_BIAS.n1186 0.189894
R32277 CS_BIAS.n1251 CS_BIAS.n1186 0.189894
R32278 CS_BIAS.n1252 CS_BIAS.n1251 0.189894
R32279 CS_BIAS.n1253 CS_BIAS.n1252 0.189894
R32280 CS_BIAS.n1253 CS_BIAS.n1184 0.189894
R32281 CS_BIAS.n1257 CS_BIAS.n1184 0.189894
R32282 CS_BIAS.n1258 CS_BIAS.n1257 0.189894
R32283 CS_BIAS.n1259 CS_BIAS.n1258 0.189894
R32284 CS_BIAS.n1259 CS_BIAS.n1182 0.189894
R32285 CS_BIAS.n1264 CS_BIAS.n1182 0.189894
R32286 CS_BIAS.n1265 CS_BIAS.n1264 0.189894
R32287 CS_BIAS.n1266 CS_BIAS.n1265 0.189894
R32288 CS_BIAS.n1266 CS_BIAS.n1180 0.189894
R32289 CS_BIAS.n1270 CS_BIAS.n1180 0.189894
R32290 CS_BIAS.n1271 CS_BIAS.n1270 0.189894
R32291 CS_BIAS.n1272 CS_BIAS.n1271 0.189894
R32292 CS_BIAS.n1272 CS_BIAS.n1178 0.189894
R32293 CS_BIAS.n1276 CS_BIAS.n1178 0.189894
R32294 CS_BIAS.n1277 CS_BIAS.n1276 0.189894
R32295 CS_BIAS.n1278 CS_BIAS.n1277 0.189894
R32296 CS_BIAS.n1278 CS_BIAS.n1176 0.189894
R32297 CS_BIAS.n1282 CS_BIAS.n1176 0.189894
R32298 CS_BIAS.n1283 CS_BIAS.n1282 0.189894
R32299 CS_BIAS.n1283 CS_BIAS.n1174 0.189894
R32300 CS_BIAS.n1287 CS_BIAS.n1174 0.189894
R32301 CS_BIAS.n1288 CS_BIAS.n1287 0.189894
R32302 CS_BIAS.n1289 CS_BIAS.n1288 0.189894
R32303 CS_BIAS.n1289 CS_BIAS.n1172 0.189894
R32304 CS_BIAS.n1293 CS_BIAS.n1172 0.189894
R32305 CS_BIAS.n1294 CS_BIAS.n1293 0.189894
R32306 CS_BIAS.n1295 CS_BIAS.n1294 0.189894
R32307 CS_BIAS.n1295 CS_BIAS.n1170 0.189894
R32308 CS_BIAS.n1299 CS_BIAS.n1170 0.189894
R32309 CS_BIAS.n1300 CS_BIAS.n1299 0.189894
R32310 CS_BIAS.n1301 CS_BIAS.n1300 0.189894
R32311 CS_BIAS.n1301 CS_BIAS.n1168 0.189894
R32312 CS_BIAS.n1306 CS_BIAS.n1168 0.189894
R32313 CS_BIAS.n1307 CS_BIAS.n1306 0.189894
R32314 CS_BIAS.n1308 CS_BIAS.n1307 0.189894
R32315 CS_BIAS.n1308 CS_BIAS.n1166 0.189894
R32316 CS_BIAS.n1312 CS_BIAS.n1166 0.189894
R32317 CS_BIAS.n1313 CS_BIAS.n1312 0.189894
R32318 CS_BIAS.n1314 CS_BIAS.n1313 0.189894
R32319 CS_BIAS.n1314 CS_BIAS.n1164 0.189894
R32320 CS_BIAS.n1318 CS_BIAS.n1164 0.189894
R32321 CS_BIAS.n1319 CS_BIAS.n1318 0.189894
R32322 CS_BIAS.n1320 CS_BIAS.n1319 0.189894
R32323 CS_BIAS.n1320 CS_BIAS.n1162 0.189894
R32324 CS_BIAS.n962 CS_BIAS.n959 0.189894
R32325 CS_BIAS.n966 CS_BIAS.n959 0.189894
R32326 CS_BIAS.n967 CS_BIAS.n966 0.189894
R32327 CS_BIAS.n968 CS_BIAS.n967 0.189894
R32328 CS_BIAS.n968 CS_BIAS.n957 0.189894
R32329 CS_BIAS.n972 CS_BIAS.n957 0.189894
R32330 CS_BIAS.n973 CS_BIAS.n972 0.189894
R32331 CS_BIAS.n974 CS_BIAS.n973 0.189894
R32332 CS_BIAS.n974 CS_BIAS.n955 0.189894
R32333 CS_BIAS.n978 CS_BIAS.n955 0.189894
R32334 CS_BIAS.n979 CS_BIAS.n978 0.189894
R32335 CS_BIAS.n980 CS_BIAS.n979 0.189894
R32336 CS_BIAS.n980 CS_BIAS.n953 0.189894
R32337 CS_BIAS.n985 CS_BIAS.n953 0.189894
R32338 CS_BIAS.n986 CS_BIAS.n985 0.189894
R32339 CS_BIAS.n987 CS_BIAS.n986 0.189894
R32340 CS_BIAS.n987 CS_BIAS.n951 0.189894
R32341 CS_BIAS.n991 CS_BIAS.n951 0.189894
R32342 CS_BIAS.n992 CS_BIAS.n991 0.189894
R32343 CS_BIAS.n993 CS_BIAS.n992 0.189894
R32344 CS_BIAS.n993 CS_BIAS.n949 0.189894
R32345 CS_BIAS.n997 CS_BIAS.n949 0.189894
R32346 CS_BIAS.n998 CS_BIAS.n997 0.189894
R32347 CS_BIAS.n999 CS_BIAS.n998 0.189894
R32348 CS_BIAS.n999 CS_BIAS.n947 0.189894
R32349 CS_BIAS.n1004 CS_BIAS.n947 0.189894
R32350 CS_BIAS.n1005 CS_BIAS.n1004 0.189894
R32351 CS_BIAS.n1006 CS_BIAS.n1005 0.189894
R32352 CS_BIAS.n1006 CS_BIAS.n945 0.189894
R32353 CS_BIAS.n1010 CS_BIAS.n945 0.189894
R32354 CS_BIAS.n1011 CS_BIAS.n1010 0.189894
R32355 CS_BIAS.n1012 CS_BIAS.n1011 0.189894
R32356 CS_BIAS.n1012 CS_BIAS.n943 0.189894
R32357 CS_BIAS.n1016 CS_BIAS.n943 0.189894
R32358 CS_BIAS.n1017 CS_BIAS.n1016 0.189894
R32359 CS_BIAS.n1018 CS_BIAS.n1017 0.189894
R32360 CS_BIAS.n1018 CS_BIAS.n941 0.189894
R32361 CS_BIAS.n1023 CS_BIAS.n941 0.189894
R32362 CS_BIAS.n1024 CS_BIAS.n1023 0.189894
R32363 CS_BIAS.n1025 CS_BIAS.n1024 0.189894
R32364 CS_BIAS.n1025 CS_BIAS.n939 0.189894
R32365 CS_BIAS.n1029 CS_BIAS.n939 0.189894
R32366 CS_BIAS.n1030 CS_BIAS.n1029 0.189894
R32367 CS_BIAS.n1031 CS_BIAS.n1030 0.189894
R32368 CS_BIAS.n1031 CS_BIAS.n937 0.189894
R32369 CS_BIAS.n1035 CS_BIAS.n937 0.189894
R32370 CS_BIAS.n1036 CS_BIAS.n1035 0.189894
R32371 CS_BIAS.n1037 CS_BIAS.n1036 0.189894
R32372 CS_BIAS.n1037 CS_BIAS.n935 0.189894
R32373 CS_BIAS.n1041 CS_BIAS.n935 0.189894
R32374 CS_BIAS.n1042 CS_BIAS.n1041 0.189894
R32375 CS_BIAS.n1042 CS_BIAS.n933 0.189894
R32376 CS_BIAS.n1046 CS_BIAS.n933 0.189894
R32377 CS_BIAS.n1047 CS_BIAS.n1046 0.189894
R32378 CS_BIAS.n1048 CS_BIAS.n1047 0.189894
R32379 CS_BIAS.n1048 CS_BIAS.n931 0.189894
R32380 CS_BIAS.n1052 CS_BIAS.n931 0.189894
R32381 CS_BIAS.n1053 CS_BIAS.n1052 0.189894
R32382 CS_BIAS.n1054 CS_BIAS.n1053 0.189894
R32383 CS_BIAS.n1054 CS_BIAS.n929 0.189894
R32384 CS_BIAS.n1058 CS_BIAS.n929 0.189894
R32385 CS_BIAS.n1059 CS_BIAS.n1058 0.189894
R32386 CS_BIAS.n1060 CS_BIAS.n1059 0.189894
R32387 CS_BIAS.n1060 CS_BIAS.n927 0.189894
R32388 CS_BIAS.n1065 CS_BIAS.n927 0.189894
R32389 CS_BIAS.n1066 CS_BIAS.n1065 0.189894
R32390 CS_BIAS.n1067 CS_BIAS.n1066 0.189894
R32391 CS_BIAS.n1067 CS_BIAS.n925 0.189894
R32392 CS_BIAS.n1071 CS_BIAS.n925 0.189894
R32393 CS_BIAS.n1072 CS_BIAS.n1071 0.189894
R32394 CS_BIAS.n1073 CS_BIAS.n1072 0.189894
R32395 CS_BIAS.n1073 CS_BIAS.n923 0.189894
R32396 CS_BIAS.n1077 CS_BIAS.n923 0.189894
R32397 CS_BIAS.n1078 CS_BIAS.n1077 0.189894
R32398 CS_BIAS.n1079 CS_BIAS.n1078 0.189894
R32399 CS_BIAS.n1079 CS_BIAS.n921 0.189894
R32400 CS_BIAS.n868 CS_BIAS.n865 0.189894
R32401 CS_BIAS.n872 CS_BIAS.n865 0.189894
R32402 CS_BIAS.n873 CS_BIAS.n872 0.189894
R32403 CS_BIAS.n874 CS_BIAS.n873 0.189894
R32404 CS_BIAS.n874 CS_BIAS.n863 0.189894
R32405 CS_BIAS.n878 CS_BIAS.n863 0.189894
R32406 CS_BIAS.n879 CS_BIAS.n878 0.189894
R32407 CS_BIAS.n880 CS_BIAS.n879 0.189894
R32408 CS_BIAS.n880 CS_BIAS.n861 0.189894
R32409 CS_BIAS.n884 CS_BIAS.n861 0.189894
R32410 CS_BIAS.n885 CS_BIAS.n884 0.189894
R32411 CS_BIAS.n886 CS_BIAS.n885 0.189894
R32412 CS_BIAS.n886 CS_BIAS.n859 0.189894
R32413 CS_BIAS.n891 CS_BIAS.n859 0.189894
R32414 CS_BIAS.n892 CS_BIAS.n891 0.189894
R32415 CS_BIAS.n893 CS_BIAS.n892 0.189894
R32416 CS_BIAS.n893 CS_BIAS.n857 0.189894
R32417 CS_BIAS.n897 CS_BIAS.n857 0.189894
R32418 CS_BIAS.n898 CS_BIAS.n897 0.189894
R32419 CS_BIAS.n899 CS_BIAS.n898 0.189894
R32420 CS_BIAS.n899 CS_BIAS.n855 0.189894
R32421 CS_BIAS.n903 CS_BIAS.n855 0.189894
R32422 CS_BIAS.n904 CS_BIAS.n903 0.189894
R32423 CS_BIAS.n905 CS_BIAS.n904 0.189894
R32424 CS_BIAS.n905 CS_BIAS.n853 0.189894
R32425 CS_BIAS.n910 CS_BIAS.n853 0.189894
R32426 CS_BIAS.n911 CS_BIAS.n910 0.189894
R32427 CS_BIAS.n912 CS_BIAS.n911 0.189894
R32428 CS_BIAS.n912 CS_BIAS.n851 0.189894
R32429 CS_BIAS.n916 CS_BIAS.n851 0.189894
R32430 CS_BIAS.n917 CS_BIAS.n916 0.189894
R32431 CS_BIAS.n1090 CS_BIAS.n849 0.189894
R32432 CS_BIAS.n1094 CS_BIAS.n849 0.189894
R32433 CS_BIAS.n1095 CS_BIAS.n1094 0.189894
R32434 CS_BIAS.n1096 CS_BIAS.n1095 0.189894
R32435 CS_BIAS.n1096 CS_BIAS.n847 0.189894
R32436 CS_BIAS.n1101 CS_BIAS.n847 0.189894
R32437 CS_BIAS.n1102 CS_BIAS.n1101 0.189894
R32438 CS_BIAS.n1103 CS_BIAS.n1102 0.189894
R32439 CS_BIAS.n1103 CS_BIAS.n845 0.189894
R32440 CS_BIAS.n1107 CS_BIAS.n845 0.189894
R32441 CS_BIAS.n1108 CS_BIAS.n1107 0.189894
R32442 CS_BIAS.n1109 CS_BIAS.n1108 0.189894
R32443 CS_BIAS.n1109 CS_BIAS.n843 0.189894
R32444 CS_BIAS.n1113 CS_BIAS.n843 0.189894
R32445 CS_BIAS.n1114 CS_BIAS.n1113 0.189894
R32446 CS_BIAS.n1115 CS_BIAS.n1114 0.189894
R32447 CS_BIAS.n1115 CS_BIAS.n841 0.189894
R32448 CS_BIAS.n1119 CS_BIAS.n841 0.189894
R32449 CS_BIAS.n1120 CS_BIAS.n1119 0.189894
R32450 CS_BIAS.n1120 CS_BIAS.n839 0.189894
R32451 CS_BIAS.n1124 CS_BIAS.n839 0.189894
R32452 CS_BIAS.n1125 CS_BIAS.n1124 0.189894
R32453 CS_BIAS.n1126 CS_BIAS.n1125 0.189894
R32454 CS_BIAS.n1126 CS_BIAS.n837 0.189894
R32455 CS_BIAS.n1130 CS_BIAS.n837 0.189894
R32456 CS_BIAS.n1131 CS_BIAS.n1130 0.189894
R32457 CS_BIAS.n1132 CS_BIAS.n1131 0.189894
R32458 CS_BIAS.n1132 CS_BIAS.n835 0.189894
R32459 CS_BIAS.n1136 CS_BIAS.n835 0.189894
R32460 CS_BIAS.n1137 CS_BIAS.n1136 0.189894
R32461 CS_BIAS.n1138 CS_BIAS.n1137 0.189894
R32462 CS_BIAS.n1138 CS_BIAS.n833 0.189894
R32463 CS_BIAS.n1143 CS_BIAS.n833 0.189894
R32464 CS_BIAS.n1144 CS_BIAS.n1143 0.189894
R32465 CS_BIAS.n1145 CS_BIAS.n1144 0.189894
R32466 CS_BIAS.n1145 CS_BIAS.n831 0.189894
R32467 CS_BIAS.n1149 CS_BIAS.n831 0.189894
R32468 CS_BIAS.n1150 CS_BIAS.n1149 0.189894
R32469 CS_BIAS.n1151 CS_BIAS.n1150 0.189894
R32470 CS_BIAS.n1151 CS_BIAS.n829 0.189894
R32471 CS_BIAS.n1155 CS_BIAS.n829 0.189894
R32472 CS_BIAS.n1156 CS_BIAS.n1155 0.189894
R32473 CS_BIAS.n1157 CS_BIAS.n1156 0.189894
R32474 CS_BIAS.n1157 CS_BIAS.n827 0.189894
R32475 CS_BIAS.n262 CS_BIAS.n90 0.0762576
R32476 CS_BIAS.n263 CS_BIAS.n262 0.0762576
R32477 CS_BIAS.n1089 CS_BIAS.n917 0.0762576
R32478 CS_BIAS.n1090 CS_BIAS.n1089 0.0762576
R32479 a_n11922_9718.n23 a_n11922_9718.t17 108.569
R32480 a_n11922_9718.n21 a_n11922_9718.t21 106.66
R32481 a_n11922_9718.n21 a_n11922_9718.n20 91.5944
R32482 a_n11922_9718.n23 a_n11922_9718.n22 89.6864
R32483 a_n11922_9718.n15 a_n11922_9718.n24 63.7938
R32484 a_n11922_9718.n19 a_n11922_9718.n18 63.7936
R32485 a_n11922_9718.n19 a_n11922_9718.n16 63.7936
R32486 a_n11922_9718.n15 a_n11922_9718.n25 62.6156
R32487 a_n11922_9718.n26 a_n11922_9718.n15 62.6156
R32488 a_n11922_9718.n19 a_n11922_9718.n17 62.6154
R32489 a_n11922_9718.n15 a_n11922_9718.n19 34.5935
R32490 a_n11922_9718.n3 a_n11922_9718.n0 1.94338
R32491 a_n11922_9718.t16 a_n11922_9718.n6 47.2366
R32492 a_n11922_9718.n14 a_n11922_9718.n12 23.5785
R32493 a_n11922_9718.n1 a_n11922_9718.n8 23.1543
R32494 a_n11922_9718.n6 a_n11922_9718.n14 21.5217
R32495 a_n11922_9718.n1 a_n11922_9718.n10 19.6429
R32496 a_n11922_9718.n20 a_n11922_9718.t15 16.9744
R32497 a_n11922_9718.n20 a_n11922_9718.t13 16.9744
R32498 a_n11922_9718.n22 a_n11922_9718.t19 16.9744
R32499 a_n11922_9718.n22 a_n11922_9718.t23 16.9744
R32500 a_n11922_9718.n0 a_n11922_9718.t43 46.8066
R32501 a_n11922_9718.n3 a_n11922_9718.t45 49.5445
R32502 a_n11922_9718.n3 a_n11922_9718.t41 46.2442
R32503 a_n11922_9718.n0 a_n11922_9718.t28 48.8027
R32504 a_n11922_9718.n0 a_n11922_9718.t32 46.8066
R32505 a_n11922_9718.n4 a_n11922_9718.t29 49.3716
R32506 a_n11922_9718.n4 a_n11922_9718.t25 46.3259
R32507 a_n11922_9718.n0 a_n11922_9718.t38 48.8027
R32508 a_n11922_9718.n0 a_n11922_9718.t27 46.8066
R32509 a_n11922_9718.n2 a_n11922_9718.t31 49.5445
R32510 a_n11922_9718.n2 a_n11922_9718.t37 46.2442
R32511 a_n11922_9718.n0 a_n11922_9718.t30 48.8027
R32512 a_n11922_9718.n0 a_n11922_9718.t34 46.8066
R32513 a_n11922_9718.n5 a_n11922_9718.t26 49.3716
R32514 a_n11922_9718.n5 a_n11922_9718.t35 46.3259
R32515 a_n11922_9718.n0 a_n11922_9718.t33 48.8027
R32516 a_n11922_9718.n11 a_n11922_9718.t14 48.9611
R32517 a_n11922_9718.n11 a_n11922_9718.t12 46.8708
R32518 a_n11922_9718.n10 a_n11922_9718.t20 47.2225
R32519 a_n11922_9718.n13 a_n11922_9718.t36 48.9611
R32520 a_n11922_9718.n13 a_n11922_9718.t39 46.8708
R32521 a_n11922_9718.n12 a_n11922_9718.t42 47.2225
R32522 a_n11922_9718.n9 a_n11922_9718.t24 48.9611
R32523 a_n11922_9718.n9 a_n11922_9718.t44 46.8708
R32524 a_n11922_9718.n8 a_n11922_9718.t40 47.2225
R32525 a_n11922_9718.n7 a_n11922_9718.t18 48.9465
R32526 a_n11922_9718.n7 a_n11922_9718.t22 46.9107
R32527 a_n11922_9718.n10 a_n11922_9718.n11 2.06013
R32528 a_n11922_9718.n12 a_n11922_9718.n13 2.06013
R32529 a_n11922_9718.n8 a_n11922_9718.n9 2.06013
R32530 a_n11922_9718.n6 a_n11922_9718.n7 2.08332
R32531 a_n11922_9718.n1 a_n11922_9718.n21 11.7984
R32532 a_n11922_9718.n14 a_n11922_9718.n23 10.8619
R32533 a_n11922_9718.n10 a_n11922_9718.n12 10.1679
R32534 a_n11922_9718.n6 a_n11922_9718.n8 9.83592
R32535 a_n11922_9718.n15 a_n11922_9718.n6 25.0777
R32536 a_n11922_9718.n0 a_n11922_9718.n1 12.624
R32537 a_n11922_9718.n14 a_n11922_9718.n0 10.321
R32538 a_n11922_9718.n24 a_n11922_9718.t9 6.6448
R32539 a_n11922_9718.n24 a_n11922_9718.t8 6.6448
R32540 a_n11922_9718.n25 a_n11922_9718.t2 6.6448
R32541 a_n11922_9718.n25 a_n11922_9718.t10 6.6448
R32542 a_n11922_9718.n18 a_n11922_9718.t5 6.6448
R32543 a_n11922_9718.n18 a_n11922_9718.t6 6.6448
R32544 a_n11922_9718.n17 a_n11922_9718.t3 6.6448
R32545 a_n11922_9718.n17 a_n11922_9718.t4 6.6448
R32546 a_n11922_9718.n16 a_n11922_9718.t11 6.6448
R32547 a_n11922_9718.n16 a_n11922_9718.t1 6.6448
R32548 a_n11922_9718.n26 a_n11922_9718.t7 6.6448
R32549 a_n11922_9718.t0 a_n11922_9718.n26 6.6448
R32550 a_n11922_9718.n2 a_n11922_9718.n0 6.5502
R32551 a_n11922_9718.n4 a_n11922_9718.n0 5.58784
R32552 a_n11922_9718.n5 a_n11922_9718.n0 5.58784
R32553 a_n6268_8041.n4 a_n6268_8041.t6 108.569
R32554 a_n6268_8041.n2 a_n6268_8041.t11 108.569
R32555 a_n6268_8041.n10 a_n6268_8041.t10 108.569
R32556 a_n6268_8041.n0 a_n6268_8041.t7 106.66
R32557 a_n6268_8041.n0 a_n6268_8041.t4 106.66
R32558 a_n6268_8041.n7 a_n6268_8041.t3 106.66
R32559 a_n6268_8041.n10 a_n6268_8041.n9 89.6864
R32560 a_n6268_8041.n4 a_n6268_8041.n3 89.6864
R32561 a_n6268_8041.n6 a_n6268_8041.n5 89.6864
R32562 a_n6268_8041.n2 a_n6268_8041.n1 89.6864
R32563 a_n6268_8041.n8 a_n6268_8041.n2 28.7911
R32564 a_n6268_8041.n9 a_n6268_8041.t13 16.9744
R32565 a_n6268_8041.n9 a_n6268_8041.t12 16.9744
R32566 a_n6268_8041.n3 a_n6268_8041.t5 16.9744
R32567 a_n6268_8041.n3 a_n6268_8041.t1 16.9744
R32568 a_n6268_8041.n5 a_n6268_8041.t8 16.9744
R32569 a_n6268_8041.n5 a_n6268_8041.t2 16.9744
R32570 a_n6268_8041.n1 a_n6268_8041.t14 16.9744
R32571 a_n6268_8041.n1 a_n6268_8041.t9 16.9744
R32572 a_n6268_8041.t0 a_n6268_8041.n11 12.8477
R32573 a_n6268_8041.n11 a_n6268_8041.n10 10.9811
R32574 a_n6268_8041.n8 a_n6268_8041.n7 5.86185
R32575 a_n6268_8041.n11 a_n6268_8041.n8 3.93611
R32576 a_n6268_8041.n6 a_n6268_8041.n0 2.36832
R32577 a_n6268_8041.n7 a_n6268_8041.n6 1.90855
R32578 a_n6268_8041.n0 a_n6268_8041.n4 1.90855
R32579 a_n6268_8041.n12 a_n6268_8041.t0 1.46436
R32580 a_n5140_n467.n4 a_n5140_n467.t25 185.928
R32581 a_n5140_n467.n6 a_n5140_n467.t12 185.928
R32582 a_n5140_n467.n7 a_n5140_n467.t27 185.928
R32583 a_n5140_n467.n8 a_n5140_n467.t26 185.928
R32584 a_n5140_n467.n1 a_n5140_n467.t16 49.672
R32585 a_n5140_n467.n1 a_n5140_n467.t10 49.672
R32586 a_n5140_n467.n5 a_n5140_n467.t9 49.672
R32587 a_n5140_n467.n21 a_n5140_n467.t13 49.6719
R32588 a_n5140_n467.n19 a_n5140_n467.t2 49.6719
R32589 a_n5140_n467.n0 a_n5140_n467.t6 49.6719
R32590 a_n5140_n467.n0 a_n5140_n467.t22 49.6719
R32591 a_n5140_n467.n10 a_n5140_n467.t21 49.6719
R32592 a_n5140_n467.n23 a_n5140_n467.n22 43.0277
R32593 a_n5140_n467.n25 a_n5140_n467.n24 43.0277
R32594 a_n5140_n467.n3 a_n5140_n467.n2 43.0277
R32595 a_n5140_n467.n27 a_n5140_n467.n26 43.0277
R32596 a_n5140_n467.n18 a_n5140_n467.n17 43.0276
R32597 a_n5140_n467.n16 a_n5140_n467.n15 43.0276
R32598 a_n5140_n467.n14 a_n5140_n467.n13 43.0276
R32599 a_n5140_n467.n12 a_n5140_n467.n11 43.0276
R32600 a_n5140_n467.n9 a_n5140_n467.n5 11.7167
R32601 a_n5140_n467.n21 a_n5140_n467.n20 11.7167
R32602 a_n5140_n467.n22 a_n5140_n467.t18 6.6448
R32603 a_n5140_n467.n22 a_n5140_n467.t20 6.6448
R32604 a_n5140_n467.n24 a_n5140_n467.t24 6.6448
R32605 a_n5140_n467.n24 a_n5140_n467.t15 6.6448
R32606 a_n5140_n467.n2 a_n5140_n467.t3 6.6448
R32607 a_n5140_n467.n2 a_n5140_n467.t0 6.6448
R32608 a_n5140_n467.n17 a_n5140_n467.t7 6.6448
R32609 a_n5140_n467.n17 a_n5140_n467.t8 6.6448
R32610 a_n5140_n467.n15 a_n5140_n467.t1 6.6448
R32611 a_n5140_n467.n15 a_n5140_n467.t4 6.6448
R32612 a_n5140_n467.n13 a_n5140_n467.t23 6.6448
R32613 a_n5140_n467.n13 a_n5140_n467.t19 6.6448
R32614 a_n5140_n467.n11 a_n5140_n467.t17 6.6448
R32615 a_n5140_n467.n11 a_n5140_n467.t14 6.6448
R32616 a_n5140_n467.t11 a_n5140_n467.n27 6.6448
R32617 a_n5140_n467.n27 a_n5140_n467.t5 6.6448
R32618 a_n5140_n467.n10 a_n5140_n467.n9 5.42507
R32619 a_n5140_n467.n20 a_n5140_n467.n19 5.42507
R32620 a_n5140_n467.n20 a_n5140_n467.n4 4.57943
R32621 a_n5140_n467.n9 a_n5140_n467.n8 3.87497
R32622 a_n5140_n467.n26 a_n5140_n467.n1 1.38268
R32623 a_n5140_n467.n16 a_n5140_n467.n0 1.38268
R32624 a_n5140_n467.n12 a_n5140_n467.n10 1.17866
R32625 a_n5140_n467.n14 a_n5140_n467.n12 1.17866
R32626 a_n5140_n467.n0 a_n5140_n467.n14 1.17866
R32627 a_n5140_n467.n18 a_n5140_n467.n16 1.17866
R32628 a_n5140_n467.n19 a_n5140_n467.n18 1.17866
R32629 a_n5140_n467.n5 a_n5140_n467.n3 1.17866
R32630 a_n5140_n467.n26 a_n5140_n467.n3 1.17866
R32631 a_n5140_n467.n1 a_n5140_n467.n25 1.17866
R32632 a_n5140_n467.n25 a_n5140_n467.n23 1.17866
R32633 a_n5140_n467.n23 a_n5140_n467.n21 1.17866
R32634 a_n5140_n467.n8 a_n5140_n467.n7 0.831895
R32635 a_n5140_n467.n7 a_n5140_n467.n6 0.831895
R32636 a_n5140_n467.n6 a_n5140_n467.n4 0.831895
R32637 a_n12066_9915.n3 a_n12066_9915.t11 128.156
R32638 a_n12066_9915.n5 a_n12066_9915.t9 127.079
R32639 a_n12066_9915.n5 a_n12066_9915.n4 109.275
R32640 a_n12066_9915.n3 a_n12066_9915.n2 109.275
R32641 a_n12066_9915.n8 a_n12066_9915.t4 108.569
R32642 a_n12066_9915.n0 a_n12066_9915.t6 106.66
R32643 a_n12066_9915.n1 a_n12066_9915.t1 106.66
R32644 a_n12066_9915.n1 a_n12066_9915.t3 106.66
R32645 a_n12066_9915.n0 a_n12066_9915.n7 89.6864
R32646 a_n12066_9915.n9 a_n12066_9915.n8 89.6864
R32647 a_n12066_9915.n6 a_n12066_9915.n5 19.1816
R32648 a_n12066_9915.n7 a_n12066_9915.t0 16.9744
R32649 a_n12066_9915.n7 a_n12066_9915.t2 16.9744
R32650 a_n12066_9915.n2 a_n12066_9915.t13 16.9744
R32651 a_n12066_9915.n2 a_n12066_9915.t8 16.9744
R32652 a_n12066_9915.n4 a_n12066_9915.t12 16.9744
R32653 a_n12066_9915.n4 a_n12066_9915.t10 16.9744
R32654 a_n12066_9915.n9 a_n12066_9915.t5 16.9744
R32655 a_n12066_9915.t7 a_n12066_9915.n9 16.9744
R32656 a_n12066_9915.n6 a_n12066_9915.n3 15.1326
R32657 a_n12066_9915.n0 a_n12066_9915.n6 5.86185
R32658 a_n12066_9915.n1 a_n12066_9915.n0 3.81659
R32659 a_n12066_9915.n8 a_n12066_9915.n1 2.36832
R32660 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t11 126.561
R32661 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.t9 124.064
R32662 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.t10 124.064
R32663 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t8 124.064
R32664 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.t5 119.267
R32665 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.t1 118.436
R32666 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.t7 118.436
R32667 DIFFPAIR_BIAS.n3 DIFFPAIR_BIAS.t3 118.436
R32668 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.t4 86.6992
R32669 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.t0 84.2033
R32670 DIFFPAIR_BIAS.n5 DIFFPAIR_BIAS.t6 84.2033
R32671 DIFFPAIR_BIAS.n6 DIFFPAIR_BIAS.t2 84.2033
R32672 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.n6 5.54086
R32673 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.n7 4.33105
R32674 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.n3 4.16522
R32675 DIFFPAIR_BIAS.n6 DIFFPAIR_BIAS.n5 2.49637
R32676 DIFFPAIR_BIAS.n5 DIFFPAIR_BIAS.n4 2.49637
R32677 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.n8 2.49634
R32678 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.n9 1.72645
R32679 DIFFPAIR_BIAS.n3 DIFFPAIR_BIAS.n2 0.831895
R32680 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.n1 0.831895
R32681 DIFFPAIR_BIAS DIFFPAIR_BIAS.n10 0.68425
R32682 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.n0 0.479693
C0 VDD VOUT 74.776f
C1 VDD VN 0.275623f
C2 VOUT VP 6.11438f
C3 a_n13678_9915# VDD 1.99126f
C4 VOUT VN 1.30726f
C5 VOUT CS_BIAS 59.749397f
C6 VP VN 18.1159f
C7 VP CS_BIAS 0.401285f
C8 VP DIFFPAIR_BIAS 8.87e-20
C9 VN CS_BIAS 0.322825f
C10 VN DIFFPAIR_BIAS 1.8e-19
C11 a_12194_9915# VDD 1.99126f
C12 DIFFPAIR_BIAS GND 33.2168f
C13 CS_BIAS GND 0.32141p
C14 VN GND 57.894295f
C15 VP GND 49.199295f
C16 VOUT GND 0.144872p
C17 VDD GND 0.96675p
C18 a_12194_9915# GND 0.765022f
C19 a_n13678_9915# GND 0.765022f
C20 a_n12066_9915.n0 GND 5.8585f
C21 a_n12066_9915.n1 GND 3.98191f
C22 a_n12066_9915.t5 GND 0.120101f
C23 a_n12066_9915.t4 GND 0.701196f
C24 a_n12066_9915.t11 GND 0.811695f
C25 a_n12066_9915.t13 GND 0.120101f
C26 a_n12066_9915.t8 GND 0.120101f
C27 a_n12066_9915.n2 GND 0.604937f
C28 a_n12066_9915.n3 GND 9.34875f
C29 a_n12066_9915.t9 GND 0.806486f
C30 a_n12066_9915.t12 GND 0.120101f
C31 a_n12066_9915.t10 GND 0.120101f
C32 a_n12066_9915.n4 GND 0.604939f
C33 a_n12066_9915.n5 GND 17.8399f
C34 a_n12066_9915.n6 GND 7.14843f
C35 a_n12066_9915.t6 GND 0.670434f
C36 a_n12066_9915.t0 GND 0.120101f
C37 a_n12066_9915.t2 GND 0.120101f
C38 a_n12066_9915.n7 GND 0.490715f
C39 a_n12066_9915.t1 GND 0.670434f
C40 a_n12066_9915.t3 GND 0.670434f
C41 a_n12066_9915.n8 GND 4.43974f
C42 a_n12066_9915.n9 GND 0.490715f
C43 a_n12066_9915.t7 GND 0.120101f
C44 a_n5140_n467.n0 GND 1.37753f
C45 a_n5140_n467.n1 GND 1.37753f
C46 a_n5140_n467.t3 GND 0.096026f
C47 a_n5140_n467.t0 GND 0.096026f
C48 a_n5140_n467.n2 GND 0.606254f
C49 a_n5140_n467.n3 GND 0.878141f
C50 a_n5140_n467.t25 GND 0.485143f
C51 a_n5140_n467.n4 GND 3.09336f
C52 a_n5140_n467.t9 GND 0.734613f
C53 a_n5140_n467.n5 GND 1.31694f
C54 a_n5140_n467.t12 GND 0.485143f
C55 a_n5140_n467.n6 GND 1.40935f
C56 a_n5140_n467.t27 GND 0.485143f
C57 a_n5140_n467.n7 GND 1.40935f
C58 a_n5140_n467.t26 GND 0.485143f
C59 a_n5140_n467.n8 GND 2.49879f
C60 a_n5140_n467.n9 GND 0.981318f
C61 a_n5140_n467.t21 GND 0.734609f
C62 a_n5140_n467.n10 GND 1.14368f
C63 a_n5140_n467.t17 GND 0.096026f
C64 a_n5140_n467.t14 GND 0.096026f
C65 a_n5140_n467.n11 GND 0.60625f
C66 a_n5140_n467.n12 GND 0.878145f
C67 a_n5140_n467.t23 GND 0.096026f
C68 a_n5140_n467.t19 GND 0.096026f
C69 a_n5140_n467.n13 GND 0.60625f
C70 a_n5140_n467.n14 GND 0.878145f
C71 a_n5140_n467.t22 GND 0.734609f
C72 a_n5140_n467.t6 GND 0.734609f
C73 a_n5140_n467.t1 GND 0.096026f
C74 a_n5140_n467.t4 GND 0.096026f
C75 a_n5140_n467.n15 GND 0.60625f
C76 a_n5140_n467.n16 GND 0.878145f
C77 a_n5140_n467.t7 GND 0.096026f
C78 a_n5140_n467.t8 GND 0.096026f
C79 a_n5140_n467.n17 GND 0.60625f
C80 a_n5140_n467.n18 GND 0.878145f
C81 a_n5140_n467.t2 GND 0.734609f
C82 a_n5140_n467.n19 GND 1.14368f
C83 a_n5140_n467.n20 GND 1.30251f
C84 a_n5140_n467.t13 GND 0.734609f
C85 a_n5140_n467.n21 GND 1.31694f
C86 a_n5140_n467.t18 GND 0.096026f
C87 a_n5140_n467.t20 GND 0.096026f
C88 a_n5140_n467.n22 GND 0.606254f
C89 a_n5140_n467.n23 GND 0.878141f
C90 a_n5140_n467.t24 GND 0.096026f
C91 a_n5140_n467.t15 GND 0.096026f
C92 a_n5140_n467.n24 GND 0.606254f
C93 a_n5140_n467.n25 GND 0.878141f
C94 a_n5140_n467.t16 GND 0.734613f
C95 a_n5140_n467.t10 GND 0.734613f
C96 a_n5140_n467.n26 GND 0.878141f
C97 a_n5140_n467.t5 GND 0.096026f
C98 a_n5140_n467.n27 GND 0.606254f
C99 a_n5140_n467.t11 GND 0.096026f
C100 a_n6268_8041.n0 GND 2.66103f
C101 a_n6268_8041.t11 GND 0.468594f
C102 a_n6268_8041.t14 GND 0.080261f
C103 a_n6268_8041.t9 GND 0.080261f
C104 a_n6268_8041.n1 GND 0.327934f
C105 a_n6268_8041.n2 GND 7.32054f
C106 a_n6268_8041.t6 GND 0.468594f
C107 a_n6268_8041.t5 GND 0.080261f
C108 a_n6268_8041.t1 GND 0.080261f
C109 a_n6268_8041.n3 GND 0.327934f
C110 a_n6268_8041.n4 GND 2.96699f
C111 a_n6268_8041.t7 GND 0.448036f
C112 a_n6268_8041.t4 GND 0.448036f
C113 a_n6268_8041.t8 GND 0.080261f
C114 a_n6268_8041.t2 GND 0.080261f
C115 a_n6268_8041.n5 GND 0.327934f
C116 a_n6268_8041.n6 GND 1.8178f
C117 a_n6268_8041.t3 GND 0.448036f
C118 a_n6268_8041.n7 GND 2.09731f
C119 a_n6268_8041.n8 GND 5.65683f
C120 a_n6268_8041.t10 GND 0.468593f
C121 a_n6268_8041.t13 GND 0.080261f
C122 a_n6268_8041.t12 GND 0.080261f
C123 a_n6268_8041.n9 GND 0.327934f
C124 a_n6268_8041.n10 GND 5.75618f
C125 a_n6268_8041.n11 GND 8.40054f
C126 a_n6268_8041.t0 GND 0.108936p
C127 a_n6268_8041.n12 GND -65.716995f
C128 a_n11922_9718.n0 GND 16.6437f
C129 a_n11922_9718.n1 GND 3.37004f
C130 a_n11922_9718.n2 GND 1.13834f
C131 a_n11922_9718.n3 GND 1.13834f
C132 a_n11922_9718.n4 GND 1.14046f
C133 a_n11922_9718.n5 GND 1.14046f
C134 a_n11922_9718.n6 GND 5.8577f
C135 a_n11922_9718.n7 GND 1.13944f
C136 a_n11922_9718.n8 GND 4.15045f
C137 a_n11922_9718.n9 GND 1.14076f
C138 a_n11922_9718.n10 GND 4.04311f
C139 a_n11922_9718.n11 GND 1.14076f
C140 a_n11922_9718.n12 GND 4.19402f
C141 a_n11922_9718.n13 GND 1.14076f
C142 a_n11922_9718.n14 GND 3.58271f
C143 a_n11922_9718.n15 GND 8.51669f
C144 a_n11922_9718.t7 GND 0.127164f
C145 a_n11922_9718.t11 GND 0.127164f
C146 a_n11922_9718.t1 GND 0.127164f
C147 a_n11922_9718.n16 GND 0.923597f
C148 a_n11922_9718.t3 GND 0.127164f
C149 a_n11922_9718.t4 GND 0.127164f
C150 a_n11922_9718.n17 GND 0.902059f
C151 a_n11922_9718.t5 GND 0.127164f
C152 a_n11922_9718.t6 GND 0.127164f
C153 a_n11922_9718.n18 GND 0.923597f
C154 a_n11922_9718.n19 GND 7.09561f
C155 a_n11922_9718.t22 GND 2.74546f
C156 a_n11922_9718.t18 GND 2.77601f
C157 a_n11922_9718.t34 GND 2.74329f
C158 a_n11922_9718.t26 GND 2.77876f
C159 a_n11922_9718.t35 GND 2.73332f
C160 a_n11922_9718.t27 GND 2.74329f
C161 a_n11922_9718.t31 GND 2.78151f
C162 a_n11922_9718.t37 GND 2.7327f
C163 a_n11922_9718.t32 GND 2.74329f
C164 a_n11922_9718.t29 GND 2.77876f
C165 a_n11922_9718.t25 GND 2.73332f
C166 a_n11922_9718.t43 GND 2.74329f
C167 a_n11922_9718.t45 GND 2.78151f
C168 a_n11922_9718.t41 GND 2.7327f
C169 a_n11922_9718.t15 GND 0.081718f
C170 a_n11922_9718.t13 GND 0.081718f
C171 a_n11922_9718.n20 GND 0.372783f
C172 a_n11922_9718.t21 GND 0.456169f
C173 a_n11922_9718.n21 GND 6.2935f
C174 a_n11922_9718.t20 GND 2.74352f
C175 a_n11922_9718.t12 GND 2.74423f
C176 a_n11922_9718.t14 GND 2.77592f
C177 a_n11922_9718.t42 GND 2.74352f
C178 a_n11922_9718.t39 GND 2.74423f
C179 a_n11922_9718.t36 GND 2.77592f
C180 a_n11922_9718.t40 GND 2.74352f
C181 a_n11922_9718.t44 GND 2.74423f
C182 a_n11922_9718.t24 GND 2.77592f
C183 a_n11922_9718.t28 GND 2.77012f
C184 a_n11922_9718.t38 GND 2.77012f
C185 a_n11922_9718.t30 GND 2.77012f
C186 a_n11922_9718.t33 GND 2.77012f
C187 a_n11922_9718.t17 GND 0.477101f
C188 a_n11922_9718.t19 GND 0.081718f
C189 a_n11922_9718.t23 GND 0.081718f
C190 a_n11922_9718.n22 GND 0.333888f
C191 a_n11922_9718.n23 GND 5.80111f
C192 a_n11922_9718.t16 GND 2.74364f
C193 a_n11922_9718.t9 GND 0.127164f
C194 a_n11922_9718.t8 GND 0.127164f
C195 a_n11922_9718.n24 GND 0.9236f
C196 a_n11922_9718.t2 GND 0.127164f
C197 a_n11922_9718.t10 GND 0.127164f
C198 a_n11922_9718.n25 GND 0.902062f
C199 a_n11922_9718.n26 GND 0.902062f
C200 a_n11922_9718.t0 GND 0.127164f
C201 CS_BIAS.n0 GND 0.012472f
C202 CS_BIAS.t85 GND 0.298599f
C203 CS_BIAS.n1 GND 0.010028f
C204 CS_BIAS.n2 GND 0.005381f
C205 CS_BIAS.n3 GND 0.004445f
C206 CS_BIAS.n4 GND 0.005381f
C207 CS_BIAS.n5 GND 0.010028f
C208 CS_BIAS.n6 GND 0.005381f
C209 CS_BIAS.t45 GND 0.298599f
C210 CS_BIAS.n7 GND 0.010028f
C211 CS_BIAS.n8 GND 0.005381f
C212 CS_BIAS.n9 GND 0.005222f
C213 CS_BIAS.n10 GND 0.005381f
C214 CS_BIAS.n11 GND 0.010028f
C215 CS_BIAS.n12 GND 0.005381f
C216 CS_BIAS.t57 GND 0.298599f
C217 CS_BIAS.n13 GND 0.114251f
C218 CS_BIAS.n14 GND 0.005381f
C219 CS_BIAS.n15 GND 0.010028f
C220 CS_BIAS.n16 GND 0.005381f
C221 CS_BIAS.n17 GND 0.010862f
C222 CS_BIAS.n18 GND 0.005381f
C223 CS_BIAS.n19 GND 0.010028f
C224 CS_BIAS.n20 GND 0.005381f
C225 CS_BIAS.t80 GND 0.298599f
C226 CS_BIAS.n21 GND 0.010028f
C227 CS_BIAS.n22 GND 0.005381f
C228 CS_BIAS.n23 GND 0.004871f
C229 CS_BIAS.n24 GND 0.005381f
C230 CS_BIAS.n25 GND 0.010028f
C231 CS_BIAS.n26 GND 0.005381f
C232 CS_BIAS.t91 GND 0.298599f
C233 CS_BIAS.n27 GND 0.010028f
C234 CS_BIAS.n28 GND 0.005381f
C235 CS_BIAS.n29 GND 0.004717f
C236 CS_BIAS.n30 GND 0.005381f
C237 CS_BIAS.n31 GND 0.010028f
C238 CS_BIAS.n32 GND 0.005381f
C239 CS_BIAS.t62 GND 0.298599f
C240 CS_BIAS.n33 GND 0.010028f
C241 CS_BIAS.n34 GND 0.005381f
C242 CS_BIAS.n35 GND 0.010872f
C243 CS_BIAS.n36 GND 0.005381f
C244 CS_BIAS.n37 GND 0.010028f
C245 CS_BIAS.n38 GND 0.005381f
C246 CS_BIAS.t84 GND 0.298599f
C247 CS_BIAS.n39 GND 0.138803f
C248 CS_BIAS.t94 GND 0.412732f
C249 CS_BIAS.n40 GND 0.207254f
C250 CS_BIAS.n41 GND 0.051546f
C251 CS_BIAS.n42 GND 0.00978f
C252 CS_BIAS.n43 GND 0.010028f
C253 CS_BIAS.n44 GND 0.010028f
C254 CS_BIAS.n45 GND 0.005381f
C255 CS_BIAS.n46 GND 0.005381f
C256 CS_BIAS.n47 GND 0.005381f
C257 CS_BIAS.n48 GND 0.010752f
C258 CS_BIAS.n49 GND 0.005222f
C259 CS_BIAS.n50 GND 0.004575f
C260 CS_BIAS.n51 GND 0.005381f
C261 CS_BIAS.n52 GND 0.005381f
C262 CS_BIAS.n53 GND 0.005381f
C263 CS_BIAS.n54 GND 0.010028f
C264 CS_BIAS.n55 GND 0.010028f
C265 CS_BIAS.n56 GND 0.010028f
C266 CS_BIAS.n57 GND 0.005381f
C267 CS_BIAS.n58 GND 0.005381f
C268 CS_BIAS.n59 GND 0.005381f
C269 CS_BIAS.n60 GND 0.005225f
C270 CS_BIAS.n61 GND 0.114251f
C271 CS_BIAS.n62 GND 0.009879f
C272 CS_BIAS.n63 GND 0.010028f
C273 CS_BIAS.n64 GND 0.005381f
C274 CS_BIAS.n65 GND 0.005381f
C275 CS_BIAS.n66 GND 0.005381f
C276 CS_BIAS.n67 GND 0.010028f
C277 CS_BIAS.n68 GND 0.010803f
C278 CS_BIAS.n69 GND 0.005039f
C279 CS_BIAS.n70 GND 0.005381f
C280 CS_BIAS.n71 GND 0.005381f
C281 CS_BIAS.n72 GND 0.005381f
C282 CS_BIAS.n73 GND 0.010862f
C283 CS_BIAS.n74 GND 0.010028f
C284 CS_BIAS.n75 GND 0.010028f
C285 CS_BIAS.n76 GND 0.005381f
C286 CS_BIAS.n77 GND 0.005381f
C287 CS_BIAS.n78 GND 0.005381f
C288 CS_BIAS.n79 GND 0.010028f
C289 CS_BIAS.n80 GND 0.005126f
C290 CS_BIAS.n81 GND 0.114251f
C291 CS_BIAS.n82 GND 0.009978f
C292 CS_BIAS.n83 GND 0.005381f
C293 CS_BIAS.n84 GND 0.005381f
C294 CS_BIAS.n85 GND 0.005381f
C295 CS_BIAS.n86 GND 0.010028f
C296 CS_BIAS.n87 GND 0.010028f
C297 CS_BIAS.n88 GND 0.010839f
C298 CS_BIAS.n89 GND 0.005381f
C299 CS_BIAS.n90 GND 0.004701f
C300 CS_BIAS.n91 GND 0.012472f
C301 CS_BIAS.t12 GND 0.298599f
C302 CS_BIAS.n92 GND 0.010028f
C303 CS_BIAS.n93 GND 0.005381f
C304 CS_BIAS.n94 GND 0.004445f
C305 CS_BIAS.n95 GND 0.005381f
C306 CS_BIAS.n96 GND 0.010028f
C307 CS_BIAS.n97 GND 0.005381f
C308 CS_BIAS.t2 GND 0.298599f
C309 CS_BIAS.n98 GND 0.010028f
C310 CS_BIAS.n99 GND 0.005381f
C311 CS_BIAS.n100 GND 0.005222f
C312 CS_BIAS.n101 GND 0.005381f
C313 CS_BIAS.n102 GND 0.010028f
C314 CS_BIAS.n103 GND 0.005381f
C315 CS_BIAS.t30 GND 0.298599f
C316 CS_BIAS.n104 GND 0.114251f
C317 CS_BIAS.n105 GND 0.005381f
C318 CS_BIAS.n106 GND 0.010028f
C319 CS_BIAS.n107 GND 0.005381f
C320 CS_BIAS.n108 GND 0.010862f
C321 CS_BIAS.n109 GND 0.005381f
C322 CS_BIAS.n110 GND 0.010028f
C323 CS_BIAS.n111 GND 0.005381f
C324 CS_BIAS.t18 GND 0.298599f
C325 CS_BIAS.n112 GND 0.010028f
C326 CS_BIAS.n113 GND 0.005381f
C327 CS_BIAS.n114 GND 0.004871f
C328 CS_BIAS.n115 GND 0.005381f
C329 CS_BIAS.n116 GND 0.010028f
C330 CS_BIAS.n117 GND 0.005381f
C331 CS_BIAS.t8 GND 0.298599f
C332 CS_BIAS.n118 GND 0.010028f
C333 CS_BIAS.n119 GND 0.005381f
C334 CS_BIAS.n120 GND 0.004717f
C335 CS_BIAS.n121 GND 0.005381f
C336 CS_BIAS.n122 GND 0.010028f
C337 CS_BIAS.n123 GND 0.005381f
C338 CS_BIAS.t24 GND 0.298599f
C339 CS_BIAS.n124 GND 0.010028f
C340 CS_BIAS.n125 GND 0.005381f
C341 CS_BIAS.n126 GND 0.010872f
C342 CS_BIAS.n127 GND 0.005381f
C343 CS_BIAS.n128 GND 0.010028f
C344 CS_BIAS.n129 GND 0.005381f
C345 CS_BIAS.t16 GND 0.298599f
C346 CS_BIAS.n130 GND 0.138803f
C347 CS_BIAS.t6 GND 0.412732f
C348 CS_BIAS.n131 GND 0.207254f
C349 CS_BIAS.n132 GND 0.051546f
C350 CS_BIAS.n133 GND 0.00978f
C351 CS_BIAS.n134 GND 0.010028f
C352 CS_BIAS.n135 GND 0.010028f
C353 CS_BIAS.n136 GND 0.005381f
C354 CS_BIAS.n137 GND 0.005381f
C355 CS_BIAS.n138 GND 0.005381f
C356 CS_BIAS.n139 GND 0.010752f
C357 CS_BIAS.n140 GND 0.005222f
C358 CS_BIAS.n141 GND 0.004575f
C359 CS_BIAS.n142 GND 0.005381f
C360 CS_BIAS.n143 GND 0.005381f
C361 CS_BIAS.n144 GND 0.005381f
C362 CS_BIAS.n145 GND 0.010028f
C363 CS_BIAS.n146 GND 0.010028f
C364 CS_BIAS.n147 GND 0.010028f
C365 CS_BIAS.n148 GND 0.005381f
C366 CS_BIAS.n149 GND 0.005381f
C367 CS_BIAS.n150 GND 0.005381f
C368 CS_BIAS.n151 GND 0.005225f
C369 CS_BIAS.n152 GND 0.114251f
C370 CS_BIAS.n153 GND 0.009879f
C371 CS_BIAS.n154 GND 0.010028f
C372 CS_BIAS.n155 GND 0.005381f
C373 CS_BIAS.n156 GND 0.005381f
C374 CS_BIAS.n157 GND 0.005381f
C375 CS_BIAS.n158 GND 0.010028f
C376 CS_BIAS.n159 GND 0.010803f
C377 CS_BIAS.n160 GND 0.005039f
C378 CS_BIAS.n161 GND 0.005381f
C379 CS_BIAS.n162 GND 0.005381f
C380 CS_BIAS.n163 GND 0.005381f
C381 CS_BIAS.n164 GND 0.010862f
C382 CS_BIAS.n165 GND 0.010028f
C383 CS_BIAS.n166 GND 0.010028f
C384 CS_BIAS.n167 GND 0.005381f
C385 CS_BIAS.n168 GND 0.005381f
C386 CS_BIAS.n169 GND 0.005381f
C387 CS_BIAS.n170 GND 0.010028f
C388 CS_BIAS.n171 GND 0.005126f
C389 CS_BIAS.n172 GND 0.114251f
C390 CS_BIAS.n173 GND 0.009978f
C391 CS_BIAS.n174 GND 0.005381f
C392 CS_BIAS.n175 GND 0.005381f
C393 CS_BIAS.n176 GND 0.005381f
C394 CS_BIAS.n177 GND 0.010028f
C395 CS_BIAS.n178 GND 0.010028f
C396 CS_BIAS.n179 GND 0.010839f
C397 CS_BIAS.n180 GND 0.005381f
C398 CS_BIAS.n181 GND 0.005381f
C399 CS_BIAS.n182 GND 0.005381f
C400 CS_BIAS.n183 GND 0.004871f
C401 CS_BIAS.n184 GND 0.010839f
C402 CS_BIAS.n185 GND 0.010028f
C403 CS_BIAS.n186 GND 0.005381f
C404 CS_BIAS.n187 GND 0.005381f
C405 CS_BIAS.n188 GND 0.005381f
C406 CS_BIAS.n189 GND 0.010028f
C407 CS_BIAS.n190 GND 0.009978f
C408 CS_BIAS.n191 GND 0.114251f
C409 CS_BIAS.n192 GND 0.005126f
C410 CS_BIAS.n193 GND 0.005381f
C411 CS_BIAS.n194 GND 0.005381f
C412 CS_BIAS.n195 GND 0.005381f
C413 CS_BIAS.n196 GND 0.010028f
C414 CS_BIAS.n197 GND 0.010028f
C415 CS_BIAS.n198 GND 0.010028f
C416 CS_BIAS.n199 GND 0.005381f
C417 CS_BIAS.n200 GND 0.005381f
C418 CS_BIAS.n201 GND 0.005381f
C419 CS_BIAS.n202 GND 0.004717f
C420 CS_BIAS.n203 GND 0.005039f
C421 CS_BIAS.n204 GND 0.010803f
C422 CS_BIAS.n205 GND 0.005381f
C423 CS_BIAS.n206 GND 0.005381f
C424 CS_BIAS.n207 GND 0.005381f
C425 CS_BIAS.n208 GND 0.010028f
C426 CS_BIAS.n209 GND 0.010028f
C427 CS_BIAS.n210 GND 0.009879f
C428 CS_BIAS.n211 GND 0.005381f
C429 CS_BIAS.n212 GND 0.005381f
C430 CS_BIAS.n213 GND 0.005225f
C431 CS_BIAS.n214 GND 0.010028f
C432 CS_BIAS.n215 GND 0.010028f
C433 CS_BIAS.n216 GND 0.005381f
C434 CS_BIAS.n217 GND 0.005381f
C435 CS_BIAS.n218 GND 0.005381f
C436 CS_BIAS.n219 GND 0.010028f
C437 CS_BIAS.n220 GND 0.010872f
C438 CS_BIAS.n221 GND 0.004575f
C439 CS_BIAS.n222 GND 0.005381f
C440 CS_BIAS.n223 GND 0.005381f
C441 CS_BIAS.n224 GND 0.005381f
C442 CS_BIAS.n225 GND 0.010752f
C443 CS_BIAS.n226 GND 0.010028f
C444 CS_BIAS.n227 GND 0.010028f
C445 CS_BIAS.n228 GND 0.005381f
C446 CS_BIAS.n229 GND 0.005381f
C447 CS_BIAS.n230 GND 0.005381f
C448 CS_BIAS.n231 GND 0.00978f
C449 CS_BIAS.n232 GND 0.114251f
C450 CS_BIAS.n233 GND 0.005324f
C451 CS_BIAS.n234 GND 0.010028f
C452 CS_BIAS.n235 GND 0.005381f
C453 CS_BIAS.n236 GND 0.005381f
C454 CS_BIAS.n237 GND 0.005381f
C455 CS_BIAS.n238 GND 0.010028f
C456 CS_BIAS.n239 GND 0.010028f
C457 CS_BIAS.n240 GND 0.010871f
C458 CS_BIAS.n241 GND 0.005381f
C459 CS_BIAS.n242 GND 0.005381f
C460 CS_BIAS.n243 GND 0.005381f
C461 CS_BIAS.n244 GND 0.005421f
C462 CS_BIAS.n245 GND 0.010684f
C463 CS_BIAS.n246 GND 0.010028f
C464 CS_BIAS.n247 GND 0.005381f
C465 CS_BIAS.n248 GND 0.005381f
C466 CS_BIAS.n249 GND 0.005381f
C467 CS_BIAS.n250 GND 0.010028f
C468 CS_BIAS.n251 GND 0.009681f
C469 CS_BIAS.n252 GND 0.139914f
C470 CS_BIAS.n253 GND 0.103802f
C471 CS_BIAS.t13 GND 0.012374f
C472 CS_BIAS.t3 GND 0.012374f
C473 CS_BIAS.n254 GND 0.082189f
C474 CS_BIAS.n255 GND 0.297682f
C475 CS_BIAS.t31 GND 0.012374f
C476 CS_BIAS.t19 GND 0.012374f
C477 CS_BIAS.n256 GND 0.082189f
C478 CS_BIAS.n257 GND 0.206306f
C479 CS_BIAS.t17 GND 0.012374f
C480 CS_BIAS.t7 GND 0.012374f
C481 CS_BIAS.n258 GND 0.089f
C482 CS_BIAS.t9 GND 0.012374f
C483 CS_BIAS.t25 GND 0.012374f
C484 CS_BIAS.n259 GND 0.082189f
C485 CS_BIAS.n260 GND 0.465097f
C486 CS_BIAS.n261 GND 0.145635f
C487 CS_BIAS.n262 GND 0.034773f
C488 CS_BIAS.n263 GND 0.004701f
C489 CS_BIAS.n264 GND 0.004871f
C490 CS_BIAS.n265 GND 0.010839f
C491 CS_BIAS.n266 GND 0.010028f
C492 CS_BIAS.n267 GND 0.005381f
C493 CS_BIAS.n268 GND 0.005381f
C494 CS_BIAS.n269 GND 0.005381f
C495 CS_BIAS.n270 GND 0.010028f
C496 CS_BIAS.n271 GND 0.009978f
C497 CS_BIAS.n272 GND 0.114251f
C498 CS_BIAS.n273 GND 0.005126f
C499 CS_BIAS.n274 GND 0.005381f
C500 CS_BIAS.n275 GND 0.005381f
C501 CS_BIAS.n276 GND 0.005381f
C502 CS_BIAS.n277 GND 0.010028f
C503 CS_BIAS.n278 GND 0.010028f
C504 CS_BIAS.n279 GND 0.010028f
C505 CS_BIAS.n280 GND 0.005381f
C506 CS_BIAS.n281 GND 0.005381f
C507 CS_BIAS.n282 GND 0.005381f
C508 CS_BIAS.n283 GND 0.004717f
C509 CS_BIAS.n284 GND 0.005039f
C510 CS_BIAS.n285 GND 0.010803f
C511 CS_BIAS.n286 GND 0.005381f
C512 CS_BIAS.n287 GND 0.005381f
C513 CS_BIAS.n288 GND 0.005381f
C514 CS_BIAS.n289 GND 0.010028f
C515 CS_BIAS.n290 GND 0.010028f
C516 CS_BIAS.n291 GND 0.009879f
C517 CS_BIAS.n292 GND 0.005381f
C518 CS_BIAS.n293 GND 0.005381f
C519 CS_BIAS.n294 GND 0.005225f
C520 CS_BIAS.n295 GND 0.010028f
C521 CS_BIAS.n296 GND 0.010028f
C522 CS_BIAS.n297 GND 0.005381f
C523 CS_BIAS.n298 GND 0.005381f
C524 CS_BIAS.n299 GND 0.005381f
C525 CS_BIAS.n300 GND 0.010028f
C526 CS_BIAS.n301 GND 0.010872f
C527 CS_BIAS.n302 GND 0.004575f
C528 CS_BIAS.n303 GND 0.005381f
C529 CS_BIAS.n304 GND 0.005381f
C530 CS_BIAS.n305 GND 0.005381f
C531 CS_BIAS.n306 GND 0.010752f
C532 CS_BIAS.n307 GND 0.010028f
C533 CS_BIAS.n308 GND 0.010028f
C534 CS_BIAS.n309 GND 0.005381f
C535 CS_BIAS.n310 GND 0.005381f
C536 CS_BIAS.n311 GND 0.005381f
C537 CS_BIAS.n312 GND 0.00978f
C538 CS_BIAS.n313 GND 0.114251f
C539 CS_BIAS.n314 GND 0.005324f
C540 CS_BIAS.n315 GND 0.010028f
C541 CS_BIAS.n316 GND 0.005381f
C542 CS_BIAS.n317 GND 0.005381f
C543 CS_BIAS.n318 GND 0.005381f
C544 CS_BIAS.n319 GND 0.010028f
C545 CS_BIAS.n320 GND 0.010028f
C546 CS_BIAS.n321 GND 0.010871f
C547 CS_BIAS.n322 GND 0.005381f
C548 CS_BIAS.n323 GND 0.005381f
C549 CS_BIAS.n324 GND 0.005381f
C550 CS_BIAS.n325 GND 0.005421f
C551 CS_BIAS.n326 GND 0.010684f
C552 CS_BIAS.n327 GND 0.010028f
C553 CS_BIAS.n328 GND 0.005381f
C554 CS_BIAS.n329 GND 0.005381f
C555 CS_BIAS.n330 GND 0.005381f
C556 CS_BIAS.n331 GND 0.010028f
C557 CS_BIAS.n332 GND 0.009681f
C558 CS_BIAS.n333 GND 0.139914f
C559 CS_BIAS.n334 GND 0.071334f
C560 CS_BIAS.n335 GND 0.012472f
C561 CS_BIAS.t95 GND 0.298599f
C562 CS_BIAS.n336 GND 0.010028f
C563 CS_BIAS.n337 GND 0.005381f
C564 CS_BIAS.n338 GND 0.004445f
C565 CS_BIAS.n339 GND 0.005381f
C566 CS_BIAS.n340 GND 0.010028f
C567 CS_BIAS.n341 GND 0.005381f
C568 CS_BIAS.t76 GND 0.298599f
C569 CS_BIAS.n342 GND 0.010028f
C570 CS_BIAS.n343 GND 0.005381f
C571 CS_BIAS.n344 GND 0.005222f
C572 CS_BIAS.n345 GND 0.005381f
C573 CS_BIAS.n346 GND 0.010028f
C574 CS_BIAS.n347 GND 0.005381f
C575 CS_BIAS.t55 GND 0.298599f
C576 CS_BIAS.n348 GND 0.114251f
C577 CS_BIAS.n349 GND 0.005381f
C578 CS_BIAS.n350 GND 0.010028f
C579 CS_BIAS.n351 GND 0.005381f
C580 CS_BIAS.n352 GND 0.010862f
C581 CS_BIAS.n353 GND 0.005381f
C582 CS_BIAS.n354 GND 0.010028f
C583 CS_BIAS.n355 GND 0.005381f
C584 CS_BIAS.t37 GND 0.298599f
C585 CS_BIAS.n356 GND 0.010028f
C586 CS_BIAS.n357 GND 0.005381f
C587 CS_BIAS.n358 GND 0.004871f
C588 CS_BIAS.n359 GND 0.005381f
C589 CS_BIAS.n360 GND 0.010028f
C590 CS_BIAS.n361 GND 0.005381f
C591 CS_BIAS.t43 GND 0.298599f
C592 CS_BIAS.n362 GND 0.010028f
C593 CS_BIAS.n363 GND 0.005381f
C594 CS_BIAS.n364 GND 0.004717f
C595 CS_BIAS.n365 GND 0.005381f
C596 CS_BIAS.n366 GND 0.010028f
C597 CS_BIAS.n367 GND 0.005381f
C598 CS_BIAS.t67 GND 0.298599f
C599 CS_BIAS.n368 GND 0.010028f
C600 CS_BIAS.n369 GND 0.005381f
C601 CS_BIAS.n370 GND 0.010872f
C602 CS_BIAS.n371 GND 0.005381f
C603 CS_BIAS.n372 GND 0.010028f
C604 CS_BIAS.n373 GND 0.005381f
C605 CS_BIAS.t50 GND 0.298599f
C606 CS_BIAS.n374 GND 0.138803f
C607 CS_BIAS.t52 GND 0.412732f
C608 CS_BIAS.n375 GND 0.207254f
C609 CS_BIAS.n376 GND 0.051546f
C610 CS_BIAS.n377 GND 0.00978f
C611 CS_BIAS.n378 GND 0.010028f
C612 CS_BIAS.n379 GND 0.010028f
C613 CS_BIAS.n380 GND 0.005381f
C614 CS_BIAS.n381 GND 0.005381f
C615 CS_BIAS.n382 GND 0.005381f
C616 CS_BIAS.n383 GND 0.010752f
C617 CS_BIAS.n384 GND 0.005222f
C618 CS_BIAS.n385 GND 0.004575f
C619 CS_BIAS.n386 GND 0.005381f
C620 CS_BIAS.n387 GND 0.005381f
C621 CS_BIAS.n388 GND 0.005381f
C622 CS_BIAS.n389 GND 0.010028f
C623 CS_BIAS.n390 GND 0.010028f
C624 CS_BIAS.n391 GND 0.010028f
C625 CS_BIAS.n392 GND 0.005381f
C626 CS_BIAS.n393 GND 0.005381f
C627 CS_BIAS.n394 GND 0.005381f
C628 CS_BIAS.n395 GND 0.005225f
C629 CS_BIAS.n396 GND 0.114251f
C630 CS_BIAS.n397 GND 0.009879f
C631 CS_BIAS.n398 GND 0.010028f
C632 CS_BIAS.n399 GND 0.005381f
C633 CS_BIAS.n400 GND 0.005381f
C634 CS_BIAS.n401 GND 0.005381f
C635 CS_BIAS.n402 GND 0.010028f
C636 CS_BIAS.n403 GND 0.010803f
C637 CS_BIAS.n404 GND 0.005039f
C638 CS_BIAS.n405 GND 0.005381f
C639 CS_BIAS.n406 GND 0.005381f
C640 CS_BIAS.n407 GND 0.005381f
C641 CS_BIAS.n408 GND 0.010862f
C642 CS_BIAS.n409 GND 0.010028f
C643 CS_BIAS.n410 GND 0.010028f
C644 CS_BIAS.n411 GND 0.005381f
C645 CS_BIAS.n412 GND 0.005381f
C646 CS_BIAS.n413 GND 0.005381f
C647 CS_BIAS.n414 GND 0.010028f
C648 CS_BIAS.n415 GND 0.005126f
C649 CS_BIAS.n416 GND 0.114251f
C650 CS_BIAS.n417 GND 0.009978f
C651 CS_BIAS.n418 GND 0.005381f
C652 CS_BIAS.n419 GND 0.005381f
C653 CS_BIAS.n420 GND 0.005381f
C654 CS_BIAS.n421 GND 0.010028f
C655 CS_BIAS.n422 GND 0.010028f
C656 CS_BIAS.n423 GND 0.010839f
C657 CS_BIAS.n424 GND 0.005381f
C658 CS_BIAS.n425 GND 0.005381f
C659 CS_BIAS.n426 GND 0.005381f
C660 CS_BIAS.n427 GND 0.004871f
C661 CS_BIAS.n428 GND 0.010839f
C662 CS_BIAS.n429 GND 0.010028f
C663 CS_BIAS.n430 GND 0.005381f
C664 CS_BIAS.n431 GND 0.005381f
C665 CS_BIAS.n432 GND 0.005381f
C666 CS_BIAS.n433 GND 0.010028f
C667 CS_BIAS.n434 GND 0.009978f
C668 CS_BIAS.n435 GND 0.114251f
C669 CS_BIAS.n436 GND 0.005126f
C670 CS_BIAS.n437 GND 0.005381f
C671 CS_BIAS.n438 GND 0.005381f
C672 CS_BIAS.n439 GND 0.005381f
C673 CS_BIAS.n440 GND 0.010028f
C674 CS_BIAS.n441 GND 0.010028f
C675 CS_BIAS.n442 GND 0.010028f
C676 CS_BIAS.n443 GND 0.005381f
C677 CS_BIAS.n444 GND 0.005381f
C678 CS_BIAS.n445 GND 0.005381f
C679 CS_BIAS.n446 GND 0.004717f
C680 CS_BIAS.n447 GND 0.005039f
C681 CS_BIAS.n448 GND 0.010803f
C682 CS_BIAS.n449 GND 0.005381f
C683 CS_BIAS.n450 GND 0.005381f
C684 CS_BIAS.n451 GND 0.005381f
C685 CS_BIAS.n452 GND 0.010028f
C686 CS_BIAS.n453 GND 0.010028f
C687 CS_BIAS.n454 GND 0.009879f
C688 CS_BIAS.n455 GND 0.005381f
C689 CS_BIAS.n456 GND 0.005381f
C690 CS_BIAS.n457 GND 0.005225f
C691 CS_BIAS.n458 GND 0.010028f
C692 CS_BIAS.n459 GND 0.010028f
C693 CS_BIAS.n460 GND 0.005381f
C694 CS_BIAS.n461 GND 0.005381f
C695 CS_BIAS.n462 GND 0.005381f
C696 CS_BIAS.n463 GND 0.010028f
C697 CS_BIAS.n464 GND 0.010872f
C698 CS_BIAS.n465 GND 0.004575f
C699 CS_BIAS.n466 GND 0.005381f
C700 CS_BIAS.n467 GND 0.005381f
C701 CS_BIAS.n468 GND 0.005381f
C702 CS_BIAS.n469 GND 0.010752f
C703 CS_BIAS.n470 GND 0.010028f
C704 CS_BIAS.n471 GND 0.010028f
C705 CS_BIAS.n472 GND 0.005381f
C706 CS_BIAS.n473 GND 0.005381f
C707 CS_BIAS.n474 GND 0.005381f
C708 CS_BIAS.n475 GND 0.00978f
C709 CS_BIAS.n476 GND 0.114251f
C710 CS_BIAS.n477 GND 0.005324f
C711 CS_BIAS.n478 GND 0.010028f
C712 CS_BIAS.n479 GND 0.005381f
C713 CS_BIAS.n480 GND 0.005381f
C714 CS_BIAS.n481 GND 0.005381f
C715 CS_BIAS.n482 GND 0.010028f
C716 CS_BIAS.n483 GND 0.010028f
C717 CS_BIAS.n484 GND 0.010871f
C718 CS_BIAS.n485 GND 0.005381f
C719 CS_BIAS.n486 GND 0.005381f
C720 CS_BIAS.n487 GND 0.005381f
C721 CS_BIAS.n488 GND 0.005421f
C722 CS_BIAS.n489 GND 0.010684f
C723 CS_BIAS.n490 GND 0.010028f
C724 CS_BIAS.n491 GND 0.005381f
C725 CS_BIAS.n492 GND 0.005381f
C726 CS_BIAS.n493 GND 0.005381f
C727 CS_BIAS.n494 GND 0.010028f
C728 CS_BIAS.n495 GND 0.009681f
C729 CS_BIAS.n496 GND 0.139914f
C730 CS_BIAS.n497 GND 0.061282f
C731 CS_BIAS.n498 GND 0.074252f
C732 CS_BIAS.n499 GND 0.012472f
C733 CS_BIAS.t61 GND 0.298599f
C734 CS_BIAS.n500 GND 0.010028f
C735 CS_BIAS.n501 GND 0.005381f
C736 CS_BIAS.n502 GND 0.004445f
C737 CS_BIAS.n503 GND 0.005381f
C738 CS_BIAS.n504 GND 0.010028f
C739 CS_BIAS.n505 GND 0.005381f
C740 CS_BIAS.t47 GND 0.298599f
C741 CS_BIAS.n506 GND 0.010028f
C742 CS_BIAS.n507 GND 0.005381f
C743 CS_BIAS.n508 GND 0.005222f
C744 CS_BIAS.n509 GND 0.005381f
C745 CS_BIAS.n510 GND 0.010028f
C746 CS_BIAS.n511 GND 0.005381f
C747 CS_BIAS.t87 GND 0.298599f
C748 CS_BIAS.n512 GND 0.114251f
C749 CS_BIAS.n513 GND 0.005381f
C750 CS_BIAS.n514 GND 0.010028f
C751 CS_BIAS.n515 GND 0.005381f
C752 CS_BIAS.n516 GND 0.010862f
C753 CS_BIAS.n517 GND 0.005381f
C754 CS_BIAS.n518 GND 0.010028f
C755 CS_BIAS.n519 GND 0.005381f
C756 CS_BIAS.t69 GND 0.298599f
C757 CS_BIAS.n520 GND 0.010028f
C758 CS_BIAS.n521 GND 0.005381f
C759 CS_BIAS.n522 GND 0.004871f
C760 CS_BIAS.n523 GND 0.005381f
C761 CS_BIAS.n524 GND 0.010028f
C762 CS_BIAS.n525 GND 0.005381f
C763 CS_BIAS.t72 GND 0.298599f
C764 CS_BIAS.n526 GND 0.010028f
C765 CS_BIAS.n527 GND 0.005381f
C766 CS_BIAS.n528 GND 0.004717f
C767 CS_BIAS.n529 GND 0.005381f
C768 CS_BIAS.n530 GND 0.010028f
C769 CS_BIAS.n531 GND 0.005381f
C770 CS_BIAS.t33 GND 0.298599f
C771 CS_BIAS.n532 GND 0.010028f
C772 CS_BIAS.n533 GND 0.005381f
C773 CS_BIAS.n534 GND 0.010872f
C774 CS_BIAS.n535 GND 0.005381f
C775 CS_BIAS.n536 GND 0.010028f
C776 CS_BIAS.n537 GND 0.005381f
C777 CS_BIAS.t79 GND 0.298599f
C778 CS_BIAS.n538 GND 0.138803f
C779 CS_BIAS.t81 GND 0.412732f
C780 CS_BIAS.n539 GND 0.207254f
C781 CS_BIAS.n540 GND 0.051546f
C782 CS_BIAS.n541 GND 0.00978f
C783 CS_BIAS.n542 GND 0.010028f
C784 CS_BIAS.n543 GND 0.010028f
C785 CS_BIAS.n544 GND 0.005381f
C786 CS_BIAS.n545 GND 0.005381f
C787 CS_BIAS.n546 GND 0.005381f
C788 CS_BIAS.n547 GND 0.010752f
C789 CS_BIAS.n548 GND 0.005222f
C790 CS_BIAS.n549 GND 0.004575f
C791 CS_BIAS.n550 GND 0.005381f
C792 CS_BIAS.n551 GND 0.005381f
C793 CS_BIAS.n552 GND 0.005381f
C794 CS_BIAS.n553 GND 0.010028f
C795 CS_BIAS.n554 GND 0.010028f
C796 CS_BIAS.n555 GND 0.010028f
C797 CS_BIAS.n556 GND 0.005381f
C798 CS_BIAS.n557 GND 0.005381f
C799 CS_BIAS.n558 GND 0.005381f
C800 CS_BIAS.n559 GND 0.005225f
C801 CS_BIAS.n560 GND 0.114251f
C802 CS_BIAS.n561 GND 0.009879f
C803 CS_BIAS.n562 GND 0.010028f
C804 CS_BIAS.n563 GND 0.005381f
C805 CS_BIAS.n564 GND 0.005381f
C806 CS_BIAS.n565 GND 0.005381f
C807 CS_BIAS.n566 GND 0.010028f
C808 CS_BIAS.n567 GND 0.010803f
C809 CS_BIAS.n568 GND 0.005039f
C810 CS_BIAS.n569 GND 0.005381f
C811 CS_BIAS.n570 GND 0.005381f
C812 CS_BIAS.n571 GND 0.005381f
C813 CS_BIAS.n572 GND 0.010862f
C814 CS_BIAS.n573 GND 0.010028f
C815 CS_BIAS.n574 GND 0.010028f
C816 CS_BIAS.n575 GND 0.005381f
C817 CS_BIAS.n576 GND 0.005381f
C818 CS_BIAS.n577 GND 0.005381f
C819 CS_BIAS.n578 GND 0.010028f
C820 CS_BIAS.n579 GND 0.005126f
C821 CS_BIAS.n580 GND 0.114251f
C822 CS_BIAS.n581 GND 0.009978f
C823 CS_BIAS.n582 GND 0.005381f
C824 CS_BIAS.n583 GND 0.005381f
C825 CS_BIAS.n584 GND 0.005381f
C826 CS_BIAS.n585 GND 0.010028f
C827 CS_BIAS.n586 GND 0.010028f
C828 CS_BIAS.n587 GND 0.010839f
C829 CS_BIAS.n588 GND 0.005381f
C830 CS_BIAS.n589 GND 0.005381f
C831 CS_BIAS.n590 GND 0.005381f
C832 CS_BIAS.n591 GND 0.004871f
C833 CS_BIAS.n592 GND 0.010839f
C834 CS_BIAS.n593 GND 0.010028f
C835 CS_BIAS.n594 GND 0.005381f
C836 CS_BIAS.n595 GND 0.005381f
C837 CS_BIAS.n596 GND 0.005381f
C838 CS_BIAS.n597 GND 0.010028f
C839 CS_BIAS.n598 GND 0.009978f
C840 CS_BIAS.n599 GND 0.114251f
C841 CS_BIAS.n600 GND 0.005126f
C842 CS_BIAS.n601 GND 0.005381f
C843 CS_BIAS.n602 GND 0.005381f
C844 CS_BIAS.n603 GND 0.005381f
C845 CS_BIAS.n604 GND 0.010028f
C846 CS_BIAS.n605 GND 0.010028f
C847 CS_BIAS.n606 GND 0.010028f
C848 CS_BIAS.n607 GND 0.005381f
C849 CS_BIAS.n608 GND 0.005381f
C850 CS_BIAS.n609 GND 0.005381f
C851 CS_BIAS.n610 GND 0.004717f
C852 CS_BIAS.n611 GND 0.005039f
C853 CS_BIAS.n612 GND 0.010803f
C854 CS_BIAS.n613 GND 0.005381f
C855 CS_BIAS.n614 GND 0.005381f
C856 CS_BIAS.n615 GND 0.005381f
C857 CS_BIAS.n616 GND 0.010028f
C858 CS_BIAS.n617 GND 0.010028f
C859 CS_BIAS.n618 GND 0.009879f
C860 CS_BIAS.n619 GND 0.005381f
C861 CS_BIAS.n620 GND 0.005381f
C862 CS_BIAS.n621 GND 0.005225f
C863 CS_BIAS.n622 GND 0.010028f
C864 CS_BIAS.n623 GND 0.010028f
C865 CS_BIAS.n624 GND 0.005381f
C866 CS_BIAS.n625 GND 0.005381f
C867 CS_BIAS.n626 GND 0.005381f
C868 CS_BIAS.n627 GND 0.010028f
C869 CS_BIAS.n628 GND 0.010872f
C870 CS_BIAS.n629 GND 0.004575f
C871 CS_BIAS.n630 GND 0.005381f
C872 CS_BIAS.n631 GND 0.005381f
C873 CS_BIAS.n632 GND 0.005381f
C874 CS_BIAS.n633 GND 0.010752f
C875 CS_BIAS.n634 GND 0.010028f
C876 CS_BIAS.n635 GND 0.010028f
C877 CS_BIAS.n636 GND 0.005381f
C878 CS_BIAS.n637 GND 0.005381f
C879 CS_BIAS.n638 GND 0.005381f
C880 CS_BIAS.n639 GND 0.00978f
C881 CS_BIAS.n640 GND 0.114251f
C882 CS_BIAS.n641 GND 0.005324f
C883 CS_BIAS.n642 GND 0.010028f
C884 CS_BIAS.n643 GND 0.005381f
C885 CS_BIAS.n644 GND 0.005381f
C886 CS_BIAS.n645 GND 0.005381f
C887 CS_BIAS.n646 GND 0.010028f
C888 CS_BIAS.n647 GND 0.010028f
C889 CS_BIAS.n648 GND 0.010871f
C890 CS_BIAS.n649 GND 0.005381f
C891 CS_BIAS.n650 GND 0.005381f
C892 CS_BIAS.n651 GND 0.005381f
C893 CS_BIAS.n652 GND 0.005421f
C894 CS_BIAS.n653 GND 0.010684f
C895 CS_BIAS.n654 GND 0.010028f
C896 CS_BIAS.n655 GND 0.005381f
C897 CS_BIAS.n656 GND 0.005381f
C898 CS_BIAS.n657 GND 0.005381f
C899 CS_BIAS.n658 GND 0.010028f
C900 CS_BIAS.n659 GND 0.009681f
C901 CS_BIAS.n660 GND 0.139914f
C902 CS_BIAS.n661 GND 0.061282f
C903 CS_BIAS.n662 GND 0.053315f
C904 CS_BIAS.n663 GND 0.012472f
C905 CS_BIAS.t93 GND 0.298599f
C906 CS_BIAS.n664 GND 0.010028f
C907 CS_BIAS.n665 GND 0.005381f
C908 CS_BIAS.n666 GND 0.004445f
C909 CS_BIAS.n667 GND 0.005381f
C910 CS_BIAS.n668 GND 0.010028f
C911 CS_BIAS.n669 GND 0.005381f
C912 CS_BIAS.t75 GND 0.298599f
C913 CS_BIAS.n670 GND 0.010028f
C914 CS_BIAS.n671 GND 0.005381f
C915 CS_BIAS.n672 GND 0.005222f
C916 CS_BIAS.n673 GND 0.005381f
C917 CS_BIAS.n674 GND 0.010028f
C918 CS_BIAS.n675 GND 0.005381f
C919 CS_BIAS.t54 GND 0.298599f
C920 CS_BIAS.n676 GND 0.114251f
C921 CS_BIAS.n677 GND 0.005381f
C922 CS_BIAS.n678 GND 0.010028f
C923 CS_BIAS.n679 GND 0.005381f
C924 CS_BIAS.n680 GND 0.010862f
C925 CS_BIAS.n681 GND 0.005381f
C926 CS_BIAS.n682 GND 0.010028f
C927 CS_BIAS.n683 GND 0.005381f
C928 CS_BIAS.t36 GND 0.298599f
C929 CS_BIAS.n684 GND 0.010028f
C930 CS_BIAS.n685 GND 0.005381f
C931 CS_BIAS.n686 GND 0.004871f
C932 CS_BIAS.n687 GND 0.005381f
C933 CS_BIAS.n688 GND 0.010028f
C934 CS_BIAS.n689 GND 0.005381f
C935 CS_BIAS.t39 GND 0.298599f
C936 CS_BIAS.n690 GND 0.010028f
C937 CS_BIAS.n691 GND 0.005381f
C938 CS_BIAS.n692 GND 0.004717f
C939 CS_BIAS.n693 GND 0.005381f
C940 CS_BIAS.n694 GND 0.010028f
C941 CS_BIAS.n695 GND 0.005381f
C942 CS_BIAS.t66 GND 0.298599f
C943 CS_BIAS.n696 GND 0.010028f
C944 CS_BIAS.n697 GND 0.005381f
C945 CS_BIAS.n698 GND 0.010872f
C946 CS_BIAS.n699 GND 0.005381f
C947 CS_BIAS.n700 GND 0.010028f
C948 CS_BIAS.n701 GND 0.005381f
C949 CS_BIAS.t49 GND 0.298599f
C950 CS_BIAS.n702 GND 0.138803f
C951 CS_BIAS.t51 GND 0.412733f
C952 CS_BIAS.n703 GND 0.207253f
C953 CS_BIAS.n704 GND 0.051546f
C954 CS_BIAS.n705 GND 0.00978f
C955 CS_BIAS.n706 GND 0.010028f
C956 CS_BIAS.n707 GND 0.010028f
C957 CS_BIAS.n708 GND 0.005381f
C958 CS_BIAS.n709 GND 0.005381f
C959 CS_BIAS.n710 GND 0.005381f
C960 CS_BIAS.n711 GND 0.010752f
C961 CS_BIAS.n712 GND 0.005222f
C962 CS_BIAS.n713 GND 0.004575f
C963 CS_BIAS.n714 GND 0.005381f
C964 CS_BIAS.n715 GND 0.005381f
C965 CS_BIAS.n716 GND 0.005381f
C966 CS_BIAS.n717 GND 0.010028f
C967 CS_BIAS.n718 GND 0.010028f
C968 CS_BIAS.n719 GND 0.010028f
C969 CS_BIAS.n720 GND 0.005381f
C970 CS_BIAS.n721 GND 0.005381f
C971 CS_BIAS.n722 GND 0.005381f
C972 CS_BIAS.n723 GND 0.005225f
C973 CS_BIAS.n724 GND 0.114251f
C974 CS_BIAS.n725 GND 0.009879f
C975 CS_BIAS.n726 GND 0.010028f
C976 CS_BIAS.n727 GND 0.005381f
C977 CS_BIAS.n728 GND 0.005381f
C978 CS_BIAS.n729 GND 0.005381f
C979 CS_BIAS.n730 GND 0.010028f
C980 CS_BIAS.n731 GND 0.010803f
C981 CS_BIAS.n732 GND 0.005039f
C982 CS_BIAS.n733 GND 0.005381f
C983 CS_BIAS.n734 GND 0.005381f
C984 CS_BIAS.n735 GND 0.005381f
C985 CS_BIAS.n736 GND 0.010862f
C986 CS_BIAS.n737 GND 0.010028f
C987 CS_BIAS.n738 GND 0.010028f
C988 CS_BIAS.n739 GND 0.005381f
C989 CS_BIAS.n740 GND 0.005381f
C990 CS_BIAS.n741 GND 0.005381f
C991 CS_BIAS.n742 GND 0.010028f
C992 CS_BIAS.n743 GND 0.005126f
C993 CS_BIAS.n744 GND 0.114251f
C994 CS_BIAS.n745 GND 0.009978f
C995 CS_BIAS.n746 GND 0.005381f
C996 CS_BIAS.n747 GND 0.005381f
C997 CS_BIAS.n748 GND 0.005381f
C998 CS_BIAS.n749 GND 0.010028f
C999 CS_BIAS.n750 GND 0.010028f
C1000 CS_BIAS.n751 GND 0.010839f
C1001 CS_BIAS.n752 GND 0.005381f
C1002 CS_BIAS.n753 GND 0.005381f
C1003 CS_BIAS.n754 GND 0.005381f
C1004 CS_BIAS.n755 GND 0.004871f
C1005 CS_BIAS.n756 GND 0.010839f
C1006 CS_BIAS.n757 GND 0.010028f
C1007 CS_BIAS.n758 GND 0.005381f
C1008 CS_BIAS.n759 GND 0.005381f
C1009 CS_BIAS.n760 GND 0.005381f
C1010 CS_BIAS.n761 GND 0.010028f
C1011 CS_BIAS.n762 GND 0.009978f
C1012 CS_BIAS.n763 GND 0.114251f
C1013 CS_BIAS.n764 GND 0.005126f
C1014 CS_BIAS.n765 GND 0.005381f
C1015 CS_BIAS.n766 GND 0.005381f
C1016 CS_BIAS.n767 GND 0.005381f
C1017 CS_BIAS.n768 GND 0.010028f
C1018 CS_BIAS.n769 GND 0.010028f
C1019 CS_BIAS.n770 GND 0.010028f
C1020 CS_BIAS.n771 GND 0.005381f
C1021 CS_BIAS.n772 GND 0.005381f
C1022 CS_BIAS.n773 GND 0.005381f
C1023 CS_BIAS.n774 GND 0.004717f
C1024 CS_BIAS.n775 GND 0.005039f
C1025 CS_BIAS.n776 GND 0.010803f
C1026 CS_BIAS.n777 GND 0.005381f
C1027 CS_BIAS.n778 GND 0.005381f
C1028 CS_BIAS.n779 GND 0.005381f
C1029 CS_BIAS.n780 GND 0.010028f
C1030 CS_BIAS.n781 GND 0.010028f
C1031 CS_BIAS.n782 GND 0.009879f
C1032 CS_BIAS.n783 GND 0.005381f
C1033 CS_BIAS.n784 GND 0.005381f
C1034 CS_BIAS.n785 GND 0.005225f
C1035 CS_BIAS.n786 GND 0.010028f
C1036 CS_BIAS.n787 GND 0.010028f
C1037 CS_BIAS.n788 GND 0.005381f
C1038 CS_BIAS.n789 GND 0.005381f
C1039 CS_BIAS.n790 GND 0.005381f
C1040 CS_BIAS.n791 GND 0.010028f
C1041 CS_BIAS.n792 GND 0.010872f
C1042 CS_BIAS.n793 GND 0.004575f
C1043 CS_BIAS.n794 GND 0.005381f
C1044 CS_BIAS.n795 GND 0.005381f
C1045 CS_BIAS.n796 GND 0.005381f
C1046 CS_BIAS.n797 GND 0.010752f
C1047 CS_BIAS.n798 GND 0.010028f
C1048 CS_BIAS.n799 GND 0.010028f
C1049 CS_BIAS.n800 GND 0.005381f
C1050 CS_BIAS.n801 GND 0.005381f
C1051 CS_BIAS.n802 GND 0.005381f
C1052 CS_BIAS.n803 GND 0.00978f
C1053 CS_BIAS.n804 GND 0.114251f
C1054 CS_BIAS.n805 GND 0.005324f
C1055 CS_BIAS.n806 GND 0.010028f
C1056 CS_BIAS.n807 GND 0.005381f
C1057 CS_BIAS.n808 GND 0.005381f
C1058 CS_BIAS.n809 GND 0.005381f
C1059 CS_BIAS.n810 GND 0.010028f
C1060 CS_BIAS.n811 GND 0.010028f
C1061 CS_BIAS.n812 GND 0.010871f
C1062 CS_BIAS.n813 GND 0.005381f
C1063 CS_BIAS.n814 GND 0.005381f
C1064 CS_BIAS.n815 GND 0.005381f
C1065 CS_BIAS.n816 GND 0.005421f
C1066 CS_BIAS.n817 GND 0.010684f
C1067 CS_BIAS.n818 GND 0.010028f
C1068 CS_BIAS.n819 GND 0.005381f
C1069 CS_BIAS.n820 GND 0.005381f
C1070 CS_BIAS.n821 GND 0.005381f
C1071 CS_BIAS.n822 GND 0.010028f
C1072 CS_BIAS.n823 GND 0.009681f
C1073 CS_BIAS.n824 GND 0.139914f
C1074 CS_BIAS.n825 GND 0.061282f
C1075 CS_BIAS.n826 GND 0.484139f
C1076 CS_BIAS.n827 GND 0.012472f
C1077 CS_BIAS.t58 GND 0.298599f
C1078 CS_BIAS.n828 GND 0.010028f
C1079 CS_BIAS.n829 GND 0.005381f
C1080 CS_BIAS.n830 GND 0.004445f
C1081 CS_BIAS.n831 GND 0.005381f
C1082 CS_BIAS.n832 GND 0.010028f
C1083 CS_BIAS.n833 GND 0.005381f
C1084 CS_BIAS.t86 GND 0.298599f
C1085 CS_BIAS.n834 GND 0.010028f
C1086 CS_BIAS.n835 GND 0.005381f
C1087 CS_BIAS.n836 GND 0.005222f
C1088 CS_BIAS.n837 GND 0.005381f
C1089 CS_BIAS.n838 GND 0.010028f
C1090 CS_BIAS.n839 GND 0.005381f
C1091 CS_BIAS.t46 GND 0.298599f
C1092 CS_BIAS.n840 GND 0.114251f
C1093 CS_BIAS.n841 GND 0.005381f
C1094 CS_BIAS.n842 GND 0.010028f
C1095 CS_BIAS.n843 GND 0.005381f
C1096 CS_BIAS.n844 GND 0.010862f
C1097 CS_BIAS.n845 GND 0.005381f
C1098 CS_BIAS.n846 GND 0.010028f
C1099 CS_BIAS.n847 GND 0.005381f
C1100 CS_BIAS.t78 GND 0.298599f
C1101 CS_BIAS.n848 GND 0.010028f
C1102 CS_BIAS.n849 GND 0.005381f
C1103 CS_BIAS.n850 GND 0.004871f
C1104 CS_BIAS.n851 GND 0.005381f
C1105 CS_BIAS.n852 GND 0.010028f
C1106 CS_BIAS.n853 GND 0.005381f
C1107 CS_BIAS.t88 GND 0.298599f
C1108 CS_BIAS.n854 GND 0.010028f
C1109 CS_BIAS.n855 GND 0.005381f
C1110 CS_BIAS.n856 GND 0.004717f
C1111 CS_BIAS.n857 GND 0.005381f
C1112 CS_BIAS.n858 GND 0.010028f
C1113 CS_BIAS.n859 GND 0.005381f
C1114 CS_BIAS.t48 GND 0.298599f
C1115 CS_BIAS.n860 GND 0.010028f
C1116 CS_BIAS.n861 GND 0.005381f
C1117 CS_BIAS.n862 GND 0.010872f
C1118 CS_BIAS.n863 GND 0.005381f
C1119 CS_BIAS.n864 GND 0.010028f
C1120 CS_BIAS.n865 GND 0.005381f
C1121 CS_BIAS.t63 GND 0.298599f
C1122 CS_BIAS.n866 GND 0.138803f
C1123 CS_BIAS.t77 GND 0.412733f
C1124 CS_BIAS.n867 GND 0.207253f
C1125 CS_BIAS.n868 GND 0.051546f
C1126 CS_BIAS.n869 GND 0.00978f
C1127 CS_BIAS.n870 GND 0.010028f
C1128 CS_BIAS.n871 GND 0.010028f
C1129 CS_BIAS.n872 GND 0.005381f
C1130 CS_BIAS.n873 GND 0.005381f
C1131 CS_BIAS.n874 GND 0.005381f
C1132 CS_BIAS.n875 GND 0.010752f
C1133 CS_BIAS.n876 GND 0.005222f
C1134 CS_BIAS.n877 GND 0.004575f
C1135 CS_BIAS.n878 GND 0.005381f
C1136 CS_BIAS.n879 GND 0.005381f
C1137 CS_BIAS.n880 GND 0.005381f
C1138 CS_BIAS.n881 GND 0.010028f
C1139 CS_BIAS.n882 GND 0.010028f
C1140 CS_BIAS.n883 GND 0.010028f
C1141 CS_BIAS.n884 GND 0.005381f
C1142 CS_BIAS.n885 GND 0.005381f
C1143 CS_BIAS.n886 GND 0.005381f
C1144 CS_BIAS.n887 GND 0.005225f
C1145 CS_BIAS.n888 GND 0.114251f
C1146 CS_BIAS.n889 GND 0.009879f
C1147 CS_BIAS.n890 GND 0.010028f
C1148 CS_BIAS.n891 GND 0.005381f
C1149 CS_BIAS.n892 GND 0.005381f
C1150 CS_BIAS.n893 GND 0.005381f
C1151 CS_BIAS.n894 GND 0.010028f
C1152 CS_BIAS.n895 GND 0.010803f
C1153 CS_BIAS.n896 GND 0.005039f
C1154 CS_BIAS.n897 GND 0.005381f
C1155 CS_BIAS.n898 GND 0.005381f
C1156 CS_BIAS.n899 GND 0.005381f
C1157 CS_BIAS.n900 GND 0.010862f
C1158 CS_BIAS.n901 GND 0.010028f
C1159 CS_BIAS.n902 GND 0.010028f
C1160 CS_BIAS.n903 GND 0.005381f
C1161 CS_BIAS.n904 GND 0.005381f
C1162 CS_BIAS.n905 GND 0.005381f
C1163 CS_BIAS.n906 GND 0.010028f
C1164 CS_BIAS.n907 GND 0.005126f
C1165 CS_BIAS.n908 GND 0.114251f
C1166 CS_BIAS.n909 GND 0.009978f
C1167 CS_BIAS.n910 GND 0.005381f
C1168 CS_BIAS.n911 GND 0.005381f
C1169 CS_BIAS.n912 GND 0.005381f
C1170 CS_BIAS.n913 GND 0.010028f
C1171 CS_BIAS.n914 GND 0.010028f
C1172 CS_BIAS.n915 GND 0.010839f
C1173 CS_BIAS.n916 GND 0.005381f
C1174 CS_BIAS.n917 GND 0.004701f
C1175 CS_BIAS.t23 GND 0.012374f
C1176 CS_BIAS.t27 GND 0.012374f
C1177 CS_BIAS.n918 GND 0.089f
C1178 CS_BIAS.t1 GND 0.012374f
C1179 CS_BIAS.t11 GND 0.012374f
C1180 CS_BIAS.n919 GND 0.082189f
C1181 CS_BIAS.n920 GND 0.465097f
C1182 CS_BIAS.n921 GND 0.012472f
C1183 CS_BIAS.t28 GND 0.298599f
C1184 CS_BIAS.n922 GND 0.010028f
C1185 CS_BIAS.n923 GND 0.005381f
C1186 CS_BIAS.n924 GND 0.004445f
C1187 CS_BIAS.n925 GND 0.005381f
C1188 CS_BIAS.n926 GND 0.010028f
C1189 CS_BIAS.n927 GND 0.005381f
C1190 CS_BIAS.t14 GND 0.298599f
C1191 CS_BIAS.n928 GND 0.010028f
C1192 CS_BIAS.n929 GND 0.005381f
C1193 CS_BIAS.n930 GND 0.005222f
C1194 CS_BIAS.n931 GND 0.005381f
C1195 CS_BIAS.n932 GND 0.010028f
C1196 CS_BIAS.n933 GND 0.005381f
C1197 CS_BIAS.t4 GND 0.298599f
C1198 CS_BIAS.n934 GND 0.114251f
C1199 CS_BIAS.n935 GND 0.005381f
C1200 CS_BIAS.n936 GND 0.010028f
C1201 CS_BIAS.n937 GND 0.005381f
C1202 CS_BIAS.n938 GND 0.010862f
C1203 CS_BIAS.n939 GND 0.005381f
C1204 CS_BIAS.n940 GND 0.010028f
C1205 CS_BIAS.n941 GND 0.005381f
C1206 CS_BIAS.t20 GND 0.298599f
C1207 CS_BIAS.n942 GND 0.010028f
C1208 CS_BIAS.n943 GND 0.005381f
C1209 CS_BIAS.n944 GND 0.004871f
C1210 CS_BIAS.n945 GND 0.005381f
C1211 CS_BIAS.n946 GND 0.010028f
C1212 CS_BIAS.n947 GND 0.005381f
C1213 CS_BIAS.t10 GND 0.298599f
C1214 CS_BIAS.n948 GND 0.010028f
C1215 CS_BIAS.n949 GND 0.005381f
C1216 CS_BIAS.n950 GND 0.004717f
C1217 CS_BIAS.n951 GND 0.005381f
C1218 CS_BIAS.n952 GND 0.010028f
C1219 CS_BIAS.n953 GND 0.005381f
C1220 CS_BIAS.t0 GND 0.298599f
C1221 CS_BIAS.n954 GND 0.010028f
C1222 CS_BIAS.n955 GND 0.005381f
C1223 CS_BIAS.n956 GND 0.010872f
C1224 CS_BIAS.n957 GND 0.005381f
C1225 CS_BIAS.n958 GND 0.010028f
C1226 CS_BIAS.n959 GND 0.005381f
C1227 CS_BIAS.t26 GND 0.298599f
C1228 CS_BIAS.n960 GND 0.138803f
C1229 CS_BIAS.t22 GND 0.412733f
C1230 CS_BIAS.n961 GND 0.207253f
C1231 CS_BIAS.n962 GND 0.051546f
C1232 CS_BIAS.n963 GND 0.00978f
C1233 CS_BIAS.n964 GND 0.010028f
C1234 CS_BIAS.n965 GND 0.010028f
C1235 CS_BIAS.n966 GND 0.005381f
C1236 CS_BIAS.n967 GND 0.005381f
C1237 CS_BIAS.n968 GND 0.005381f
C1238 CS_BIAS.n969 GND 0.010752f
C1239 CS_BIAS.n970 GND 0.005222f
C1240 CS_BIAS.n971 GND 0.004575f
C1241 CS_BIAS.n972 GND 0.005381f
C1242 CS_BIAS.n973 GND 0.005381f
C1243 CS_BIAS.n974 GND 0.005381f
C1244 CS_BIAS.n975 GND 0.010028f
C1245 CS_BIAS.n976 GND 0.010028f
C1246 CS_BIAS.n977 GND 0.010028f
C1247 CS_BIAS.n978 GND 0.005381f
C1248 CS_BIAS.n979 GND 0.005381f
C1249 CS_BIAS.n980 GND 0.005381f
C1250 CS_BIAS.n981 GND 0.005225f
C1251 CS_BIAS.n982 GND 0.114251f
C1252 CS_BIAS.n983 GND 0.009879f
C1253 CS_BIAS.n984 GND 0.010028f
C1254 CS_BIAS.n985 GND 0.005381f
C1255 CS_BIAS.n986 GND 0.005381f
C1256 CS_BIAS.n987 GND 0.005381f
C1257 CS_BIAS.n988 GND 0.010028f
C1258 CS_BIAS.n989 GND 0.010803f
C1259 CS_BIAS.n990 GND 0.005039f
C1260 CS_BIAS.n991 GND 0.005381f
C1261 CS_BIAS.n992 GND 0.005381f
C1262 CS_BIAS.n993 GND 0.005381f
C1263 CS_BIAS.n994 GND 0.010862f
C1264 CS_BIAS.n995 GND 0.010028f
C1265 CS_BIAS.n996 GND 0.010028f
C1266 CS_BIAS.n997 GND 0.005381f
C1267 CS_BIAS.n998 GND 0.005381f
C1268 CS_BIAS.n999 GND 0.005381f
C1269 CS_BIAS.n1000 GND 0.010028f
C1270 CS_BIAS.n1001 GND 0.005126f
C1271 CS_BIAS.n1002 GND 0.114251f
C1272 CS_BIAS.n1003 GND 0.009978f
C1273 CS_BIAS.n1004 GND 0.005381f
C1274 CS_BIAS.n1005 GND 0.005381f
C1275 CS_BIAS.n1006 GND 0.005381f
C1276 CS_BIAS.n1007 GND 0.010028f
C1277 CS_BIAS.n1008 GND 0.010028f
C1278 CS_BIAS.n1009 GND 0.010839f
C1279 CS_BIAS.n1010 GND 0.005381f
C1280 CS_BIAS.n1011 GND 0.005381f
C1281 CS_BIAS.n1012 GND 0.005381f
C1282 CS_BIAS.n1013 GND 0.004871f
C1283 CS_BIAS.n1014 GND 0.010839f
C1284 CS_BIAS.n1015 GND 0.010028f
C1285 CS_BIAS.n1016 GND 0.005381f
C1286 CS_BIAS.n1017 GND 0.005381f
C1287 CS_BIAS.n1018 GND 0.005381f
C1288 CS_BIAS.n1019 GND 0.010028f
C1289 CS_BIAS.n1020 GND 0.009978f
C1290 CS_BIAS.n1021 GND 0.114251f
C1291 CS_BIAS.n1022 GND 0.005126f
C1292 CS_BIAS.n1023 GND 0.005381f
C1293 CS_BIAS.n1024 GND 0.005381f
C1294 CS_BIAS.n1025 GND 0.005381f
C1295 CS_BIAS.n1026 GND 0.010028f
C1296 CS_BIAS.n1027 GND 0.010028f
C1297 CS_BIAS.n1028 GND 0.010028f
C1298 CS_BIAS.n1029 GND 0.005381f
C1299 CS_BIAS.n1030 GND 0.005381f
C1300 CS_BIAS.n1031 GND 0.005381f
C1301 CS_BIAS.n1032 GND 0.004717f
C1302 CS_BIAS.n1033 GND 0.005039f
C1303 CS_BIAS.n1034 GND 0.010803f
C1304 CS_BIAS.n1035 GND 0.005381f
C1305 CS_BIAS.n1036 GND 0.005381f
C1306 CS_BIAS.n1037 GND 0.005381f
C1307 CS_BIAS.n1038 GND 0.010028f
C1308 CS_BIAS.n1039 GND 0.010028f
C1309 CS_BIAS.n1040 GND 0.009879f
C1310 CS_BIAS.n1041 GND 0.005381f
C1311 CS_BIAS.n1042 GND 0.005381f
C1312 CS_BIAS.n1043 GND 0.005225f
C1313 CS_BIAS.n1044 GND 0.010028f
C1314 CS_BIAS.n1045 GND 0.010028f
C1315 CS_BIAS.n1046 GND 0.005381f
C1316 CS_BIAS.n1047 GND 0.005381f
C1317 CS_BIAS.n1048 GND 0.005381f
C1318 CS_BIAS.n1049 GND 0.010028f
C1319 CS_BIAS.n1050 GND 0.010872f
C1320 CS_BIAS.n1051 GND 0.004575f
C1321 CS_BIAS.n1052 GND 0.005381f
C1322 CS_BIAS.n1053 GND 0.005381f
C1323 CS_BIAS.n1054 GND 0.005381f
C1324 CS_BIAS.n1055 GND 0.010752f
C1325 CS_BIAS.n1056 GND 0.010028f
C1326 CS_BIAS.n1057 GND 0.010028f
C1327 CS_BIAS.n1058 GND 0.005381f
C1328 CS_BIAS.n1059 GND 0.005381f
C1329 CS_BIAS.n1060 GND 0.005381f
C1330 CS_BIAS.n1061 GND 0.00978f
C1331 CS_BIAS.n1062 GND 0.114251f
C1332 CS_BIAS.n1063 GND 0.005324f
C1333 CS_BIAS.n1064 GND 0.010028f
C1334 CS_BIAS.n1065 GND 0.005381f
C1335 CS_BIAS.n1066 GND 0.005381f
C1336 CS_BIAS.n1067 GND 0.005381f
C1337 CS_BIAS.n1068 GND 0.010028f
C1338 CS_BIAS.n1069 GND 0.010028f
C1339 CS_BIAS.n1070 GND 0.010871f
C1340 CS_BIAS.n1071 GND 0.005381f
C1341 CS_BIAS.n1072 GND 0.005381f
C1342 CS_BIAS.n1073 GND 0.005381f
C1343 CS_BIAS.n1074 GND 0.005421f
C1344 CS_BIAS.n1075 GND 0.010684f
C1345 CS_BIAS.n1076 GND 0.010028f
C1346 CS_BIAS.n1077 GND 0.005381f
C1347 CS_BIAS.n1078 GND 0.005381f
C1348 CS_BIAS.n1079 GND 0.005381f
C1349 CS_BIAS.n1080 GND 0.010028f
C1350 CS_BIAS.n1081 GND 0.009681f
C1351 CS_BIAS.n1082 GND 0.139914f
C1352 CS_BIAS.n1083 GND 0.103802f
C1353 CS_BIAS.t15 GND 0.012374f
C1354 CS_BIAS.t29 GND 0.012374f
C1355 CS_BIAS.n1084 GND 0.082189f
C1356 CS_BIAS.n1085 GND 0.297682f
C1357 CS_BIAS.t21 GND 0.012374f
C1358 CS_BIAS.t5 GND 0.012374f
C1359 CS_BIAS.n1086 GND 0.082189f
C1360 CS_BIAS.n1087 GND 0.206306f
C1361 CS_BIAS.n1088 GND 0.145635f
C1362 CS_BIAS.n1089 GND 0.034773f
C1363 CS_BIAS.n1090 GND 0.004701f
C1364 CS_BIAS.n1091 GND 0.004871f
C1365 CS_BIAS.n1092 GND 0.010839f
C1366 CS_BIAS.n1093 GND 0.010028f
C1367 CS_BIAS.n1094 GND 0.005381f
C1368 CS_BIAS.n1095 GND 0.005381f
C1369 CS_BIAS.n1096 GND 0.005381f
C1370 CS_BIAS.n1097 GND 0.010028f
C1371 CS_BIAS.n1098 GND 0.009978f
C1372 CS_BIAS.n1099 GND 0.114251f
C1373 CS_BIAS.n1100 GND 0.005126f
C1374 CS_BIAS.n1101 GND 0.005381f
C1375 CS_BIAS.n1102 GND 0.005381f
C1376 CS_BIAS.n1103 GND 0.005381f
C1377 CS_BIAS.n1104 GND 0.010028f
C1378 CS_BIAS.n1105 GND 0.010028f
C1379 CS_BIAS.n1106 GND 0.010028f
C1380 CS_BIAS.n1107 GND 0.005381f
C1381 CS_BIAS.n1108 GND 0.005381f
C1382 CS_BIAS.n1109 GND 0.005381f
C1383 CS_BIAS.n1110 GND 0.004717f
C1384 CS_BIAS.n1111 GND 0.005039f
C1385 CS_BIAS.n1112 GND 0.010803f
C1386 CS_BIAS.n1113 GND 0.005381f
C1387 CS_BIAS.n1114 GND 0.005381f
C1388 CS_BIAS.n1115 GND 0.005381f
C1389 CS_BIAS.n1116 GND 0.010028f
C1390 CS_BIAS.n1117 GND 0.010028f
C1391 CS_BIAS.n1118 GND 0.009879f
C1392 CS_BIAS.n1119 GND 0.005381f
C1393 CS_BIAS.n1120 GND 0.005381f
C1394 CS_BIAS.n1121 GND 0.005225f
C1395 CS_BIAS.n1122 GND 0.010028f
C1396 CS_BIAS.n1123 GND 0.010028f
C1397 CS_BIAS.n1124 GND 0.005381f
C1398 CS_BIAS.n1125 GND 0.005381f
C1399 CS_BIAS.n1126 GND 0.005381f
C1400 CS_BIAS.n1127 GND 0.010028f
C1401 CS_BIAS.n1128 GND 0.010872f
C1402 CS_BIAS.n1129 GND 0.004575f
C1403 CS_BIAS.n1130 GND 0.005381f
C1404 CS_BIAS.n1131 GND 0.005381f
C1405 CS_BIAS.n1132 GND 0.005381f
C1406 CS_BIAS.n1133 GND 0.010752f
C1407 CS_BIAS.n1134 GND 0.010028f
C1408 CS_BIAS.n1135 GND 0.010028f
C1409 CS_BIAS.n1136 GND 0.005381f
C1410 CS_BIAS.n1137 GND 0.005381f
C1411 CS_BIAS.n1138 GND 0.005381f
C1412 CS_BIAS.n1139 GND 0.00978f
C1413 CS_BIAS.n1140 GND 0.114251f
C1414 CS_BIAS.n1141 GND 0.005324f
C1415 CS_BIAS.n1142 GND 0.010028f
C1416 CS_BIAS.n1143 GND 0.005381f
C1417 CS_BIAS.n1144 GND 0.005381f
C1418 CS_BIAS.n1145 GND 0.005381f
C1419 CS_BIAS.n1146 GND 0.010028f
C1420 CS_BIAS.n1147 GND 0.010028f
C1421 CS_BIAS.n1148 GND 0.010871f
C1422 CS_BIAS.n1149 GND 0.005381f
C1423 CS_BIAS.n1150 GND 0.005381f
C1424 CS_BIAS.n1151 GND 0.005381f
C1425 CS_BIAS.n1152 GND 0.005421f
C1426 CS_BIAS.n1153 GND 0.010684f
C1427 CS_BIAS.n1154 GND 0.010028f
C1428 CS_BIAS.n1155 GND 0.005381f
C1429 CS_BIAS.n1156 GND 0.005381f
C1430 CS_BIAS.n1157 GND 0.005381f
C1431 CS_BIAS.n1158 GND 0.010028f
C1432 CS_BIAS.n1159 GND 0.009681f
C1433 CS_BIAS.n1160 GND 0.139914f
C1434 CS_BIAS.n1161 GND 0.071334f
C1435 CS_BIAS.n1162 GND 0.012472f
C1436 CS_BIAS.t41 GND 0.298599f
C1437 CS_BIAS.n1163 GND 0.010028f
C1438 CS_BIAS.n1164 GND 0.005381f
C1439 CS_BIAS.n1165 GND 0.004445f
C1440 CS_BIAS.n1166 GND 0.005381f
C1441 CS_BIAS.n1167 GND 0.010028f
C1442 CS_BIAS.n1168 GND 0.005381f
C1443 CS_BIAS.t89 GND 0.298599f
C1444 CS_BIAS.n1169 GND 0.010028f
C1445 CS_BIAS.n1170 GND 0.005381f
C1446 CS_BIAS.n1171 GND 0.005222f
C1447 CS_BIAS.n1172 GND 0.005381f
C1448 CS_BIAS.n1173 GND 0.010028f
C1449 CS_BIAS.n1174 GND 0.005381f
C1450 CS_BIAS.t74 GND 0.298599f
C1451 CS_BIAS.n1175 GND 0.114251f
C1452 CS_BIAS.n1176 GND 0.005381f
C1453 CS_BIAS.n1177 GND 0.010028f
C1454 CS_BIAS.n1178 GND 0.005381f
C1455 CS_BIAS.n1179 GND 0.010862f
C1456 CS_BIAS.n1180 GND 0.005381f
C1457 CS_BIAS.n1181 GND 0.010028f
C1458 CS_BIAS.n1182 GND 0.005381f
C1459 CS_BIAS.t35 GND 0.298599f
C1460 CS_BIAS.n1183 GND 0.010028f
C1461 CS_BIAS.n1184 GND 0.005381f
C1462 CS_BIAS.n1185 GND 0.004871f
C1463 CS_BIAS.n1186 GND 0.005381f
C1464 CS_BIAS.n1187 GND 0.010028f
C1465 CS_BIAS.n1188 GND 0.005381f
C1466 CS_BIAS.t40 GND 0.298599f
C1467 CS_BIAS.n1189 GND 0.010028f
C1468 CS_BIAS.n1190 GND 0.005381f
C1469 CS_BIAS.n1191 GND 0.004717f
C1470 CS_BIAS.n1192 GND 0.005381f
C1471 CS_BIAS.n1193 GND 0.010028f
C1472 CS_BIAS.n1194 GND 0.005381f
C1473 CS_BIAS.t83 GND 0.298599f
C1474 CS_BIAS.n1195 GND 0.010028f
C1475 CS_BIAS.n1196 GND 0.005381f
C1476 CS_BIAS.n1197 GND 0.010872f
C1477 CS_BIAS.n1198 GND 0.005381f
C1478 CS_BIAS.n1199 GND 0.010028f
C1479 CS_BIAS.n1200 GND 0.005381f
C1480 CS_BIAS.t60 GND 0.298599f
C1481 CS_BIAS.n1201 GND 0.138803f
C1482 CS_BIAS.t65 GND 0.412733f
C1483 CS_BIAS.n1202 GND 0.207253f
C1484 CS_BIAS.n1203 GND 0.051546f
C1485 CS_BIAS.n1204 GND 0.00978f
C1486 CS_BIAS.n1205 GND 0.010028f
C1487 CS_BIAS.n1206 GND 0.010028f
C1488 CS_BIAS.n1207 GND 0.005381f
C1489 CS_BIAS.n1208 GND 0.005381f
C1490 CS_BIAS.n1209 GND 0.005381f
C1491 CS_BIAS.n1210 GND 0.010752f
C1492 CS_BIAS.n1211 GND 0.005222f
C1493 CS_BIAS.n1212 GND 0.004575f
C1494 CS_BIAS.n1213 GND 0.005381f
C1495 CS_BIAS.n1214 GND 0.005381f
C1496 CS_BIAS.n1215 GND 0.005381f
C1497 CS_BIAS.n1216 GND 0.010028f
C1498 CS_BIAS.n1217 GND 0.010028f
C1499 CS_BIAS.n1218 GND 0.010028f
C1500 CS_BIAS.n1219 GND 0.005381f
C1501 CS_BIAS.n1220 GND 0.005381f
C1502 CS_BIAS.n1221 GND 0.005381f
C1503 CS_BIAS.n1222 GND 0.005225f
C1504 CS_BIAS.n1223 GND 0.114251f
C1505 CS_BIAS.n1224 GND 0.009879f
C1506 CS_BIAS.n1225 GND 0.010028f
C1507 CS_BIAS.n1226 GND 0.005381f
C1508 CS_BIAS.n1227 GND 0.005381f
C1509 CS_BIAS.n1228 GND 0.005381f
C1510 CS_BIAS.n1229 GND 0.010028f
C1511 CS_BIAS.n1230 GND 0.010803f
C1512 CS_BIAS.n1231 GND 0.005039f
C1513 CS_BIAS.n1232 GND 0.005381f
C1514 CS_BIAS.n1233 GND 0.005381f
C1515 CS_BIAS.n1234 GND 0.005381f
C1516 CS_BIAS.n1235 GND 0.010862f
C1517 CS_BIAS.n1236 GND 0.010028f
C1518 CS_BIAS.n1237 GND 0.010028f
C1519 CS_BIAS.n1238 GND 0.005381f
C1520 CS_BIAS.n1239 GND 0.005381f
C1521 CS_BIAS.n1240 GND 0.005381f
C1522 CS_BIAS.n1241 GND 0.010028f
C1523 CS_BIAS.n1242 GND 0.005126f
C1524 CS_BIAS.n1243 GND 0.114251f
C1525 CS_BIAS.n1244 GND 0.009978f
C1526 CS_BIAS.n1245 GND 0.005381f
C1527 CS_BIAS.n1246 GND 0.005381f
C1528 CS_BIAS.n1247 GND 0.005381f
C1529 CS_BIAS.n1248 GND 0.010028f
C1530 CS_BIAS.n1249 GND 0.010028f
C1531 CS_BIAS.n1250 GND 0.010839f
C1532 CS_BIAS.n1251 GND 0.005381f
C1533 CS_BIAS.n1252 GND 0.005381f
C1534 CS_BIAS.n1253 GND 0.005381f
C1535 CS_BIAS.n1254 GND 0.004871f
C1536 CS_BIAS.n1255 GND 0.010839f
C1537 CS_BIAS.n1256 GND 0.010028f
C1538 CS_BIAS.n1257 GND 0.005381f
C1539 CS_BIAS.n1258 GND 0.005381f
C1540 CS_BIAS.n1259 GND 0.005381f
C1541 CS_BIAS.n1260 GND 0.010028f
C1542 CS_BIAS.n1261 GND 0.009978f
C1543 CS_BIAS.n1262 GND 0.114251f
C1544 CS_BIAS.n1263 GND 0.005126f
C1545 CS_BIAS.n1264 GND 0.005381f
C1546 CS_BIAS.n1265 GND 0.005381f
C1547 CS_BIAS.n1266 GND 0.005381f
C1548 CS_BIAS.n1267 GND 0.010028f
C1549 CS_BIAS.n1268 GND 0.010028f
C1550 CS_BIAS.n1269 GND 0.010028f
C1551 CS_BIAS.n1270 GND 0.005381f
C1552 CS_BIAS.n1271 GND 0.005381f
C1553 CS_BIAS.n1272 GND 0.005381f
C1554 CS_BIAS.n1273 GND 0.004717f
C1555 CS_BIAS.n1274 GND 0.005039f
C1556 CS_BIAS.n1275 GND 0.010803f
C1557 CS_BIAS.n1276 GND 0.005381f
C1558 CS_BIAS.n1277 GND 0.005381f
C1559 CS_BIAS.n1278 GND 0.005381f
C1560 CS_BIAS.n1279 GND 0.010028f
C1561 CS_BIAS.n1280 GND 0.010028f
C1562 CS_BIAS.n1281 GND 0.009879f
C1563 CS_BIAS.n1282 GND 0.005381f
C1564 CS_BIAS.n1283 GND 0.005381f
C1565 CS_BIAS.n1284 GND 0.005225f
C1566 CS_BIAS.n1285 GND 0.010028f
C1567 CS_BIAS.n1286 GND 0.010028f
C1568 CS_BIAS.n1287 GND 0.005381f
C1569 CS_BIAS.n1288 GND 0.005381f
C1570 CS_BIAS.n1289 GND 0.005381f
C1571 CS_BIAS.n1290 GND 0.010028f
C1572 CS_BIAS.n1291 GND 0.010872f
C1573 CS_BIAS.n1292 GND 0.004575f
C1574 CS_BIAS.n1293 GND 0.005381f
C1575 CS_BIAS.n1294 GND 0.005381f
C1576 CS_BIAS.n1295 GND 0.005381f
C1577 CS_BIAS.n1296 GND 0.010752f
C1578 CS_BIAS.n1297 GND 0.010028f
C1579 CS_BIAS.n1298 GND 0.010028f
C1580 CS_BIAS.n1299 GND 0.005381f
C1581 CS_BIAS.n1300 GND 0.005381f
C1582 CS_BIAS.n1301 GND 0.005381f
C1583 CS_BIAS.n1302 GND 0.00978f
C1584 CS_BIAS.n1303 GND 0.114251f
C1585 CS_BIAS.n1304 GND 0.005324f
C1586 CS_BIAS.n1305 GND 0.010028f
C1587 CS_BIAS.n1306 GND 0.005381f
C1588 CS_BIAS.n1307 GND 0.005381f
C1589 CS_BIAS.n1308 GND 0.005381f
C1590 CS_BIAS.n1309 GND 0.010028f
C1591 CS_BIAS.n1310 GND 0.010028f
C1592 CS_BIAS.n1311 GND 0.010871f
C1593 CS_BIAS.n1312 GND 0.005381f
C1594 CS_BIAS.n1313 GND 0.005381f
C1595 CS_BIAS.n1314 GND 0.005381f
C1596 CS_BIAS.n1315 GND 0.005421f
C1597 CS_BIAS.n1316 GND 0.010684f
C1598 CS_BIAS.n1317 GND 0.010028f
C1599 CS_BIAS.n1318 GND 0.005381f
C1600 CS_BIAS.n1319 GND 0.005381f
C1601 CS_BIAS.n1320 GND 0.005381f
C1602 CS_BIAS.n1321 GND 0.010028f
C1603 CS_BIAS.n1322 GND 0.009681f
C1604 CS_BIAS.n1323 GND 0.139914f
C1605 CS_BIAS.n1324 GND 0.061282f
C1606 CS_BIAS.n1325 GND 0.074252f
C1607 CS_BIAS.n1326 GND 0.012472f
C1608 CS_BIAS.t71 GND 0.298599f
C1609 CS_BIAS.n1327 GND 0.010028f
C1610 CS_BIAS.n1328 GND 0.005381f
C1611 CS_BIAS.n1329 GND 0.004445f
C1612 CS_BIAS.n1330 GND 0.005381f
C1613 CS_BIAS.n1331 GND 0.010028f
C1614 CS_BIAS.n1332 GND 0.005381f
C1615 CS_BIAS.t56 GND 0.298599f
C1616 CS_BIAS.n1333 GND 0.010028f
C1617 CS_BIAS.n1334 GND 0.005381f
C1618 CS_BIAS.n1335 GND 0.005222f
C1619 CS_BIAS.n1336 GND 0.005381f
C1620 CS_BIAS.n1337 GND 0.010028f
C1621 CS_BIAS.n1338 GND 0.005381f
C1622 CS_BIAS.t44 GND 0.298599f
C1623 CS_BIAS.n1339 GND 0.114251f
C1624 CS_BIAS.n1340 GND 0.005381f
C1625 CS_BIAS.n1341 GND 0.010028f
C1626 CS_BIAS.n1342 GND 0.005381f
C1627 CS_BIAS.n1343 GND 0.010862f
C1628 CS_BIAS.n1344 GND 0.005381f
C1629 CS_BIAS.n1345 GND 0.010028f
C1630 CS_BIAS.n1346 GND 0.005381f
C1631 CS_BIAS.t68 GND 0.298599f
C1632 CS_BIAS.n1347 GND 0.010028f
C1633 CS_BIAS.n1348 GND 0.005381f
C1634 CS_BIAS.n1349 GND 0.004871f
C1635 CS_BIAS.n1350 GND 0.005381f
C1636 CS_BIAS.n1351 GND 0.010028f
C1637 CS_BIAS.n1352 GND 0.005381f
C1638 CS_BIAS.t70 GND 0.298599f
C1639 CS_BIAS.n1353 GND 0.010028f
C1640 CS_BIAS.n1354 GND 0.005381f
C1641 CS_BIAS.n1355 GND 0.004717f
C1642 CS_BIAS.n1356 GND 0.005381f
C1643 CS_BIAS.n1357 GND 0.010028f
C1644 CS_BIAS.n1358 GND 0.005381f
C1645 CS_BIAS.t53 GND 0.298599f
C1646 CS_BIAS.n1359 GND 0.010028f
C1647 CS_BIAS.n1360 GND 0.005381f
C1648 CS_BIAS.n1361 GND 0.010872f
C1649 CS_BIAS.n1362 GND 0.005381f
C1650 CS_BIAS.n1363 GND 0.010028f
C1651 CS_BIAS.n1364 GND 0.005381f
C1652 CS_BIAS.t92 GND 0.298599f
C1653 CS_BIAS.n1365 GND 0.138803f
C1654 CS_BIAS.t32 GND 0.412733f
C1655 CS_BIAS.n1366 GND 0.207253f
C1656 CS_BIAS.n1367 GND 0.051546f
C1657 CS_BIAS.n1368 GND 0.00978f
C1658 CS_BIAS.n1369 GND 0.010028f
C1659 CS_BIAS.n1370 GND 0.010028f
C1660 CS_BIAS.n1371 GND 0.005381f
C1661 CS_BIAS.n1372 GND 0.005381f
C1662 CS_BIAS.n1373 GND 0.005381f
C1663 CS_BIAS.n1374 GND 0.010752f
C1664 CS_BIAS.n1375 GND 0.005222f
C1665 CS_BIAS.n1376 GND 0.004575f
C1666 CS_BIAS.n1377 GND 0.005381f
C1667 CS_BIAS.n1378 GND 0.005381f
C1668 CS_BIAS.n1379 GND 0.005381f
C1669 CS_BIAS.n1380 GND 0.010028f
C1670 CS_BIAS.n1381 GND 0.010028f
C1671 CS_BIAS.n1382 GND 0.010028f
C1672 CS_BIAS.n1383 GND 0.005381f
C1673 CS_BIAS.n1384 GND 0.005381f
C1674 CS_BIAS.n1385 GND 0.005381f
C1675 CS_BIAS.n1386 GND 0.005225f
C1676 CS_BIAS.n1387 GND 0.114251f
C1677 CS_BIAS.n1388 GND 0.009879f
C1678 CS_BIAS.n1389 GND 0.010028f
C1679 CS_BIAS.n1390 GND 0.005381f
C1680 CS_BIAS.n1391 GND 0.005381f
C1681 CS_BIAS.n1392 GND 0.005381f
C1682 CS_BIAS.n1393 GND 0.010028f
C1683 CS_BIAS.n1394 GND 0.010803f
C1684 CS_BIAS.n1395 GND 0.005039f
C1685 CS_BIAS.n1396 GND 0.005381f
C1686 CS_BIAS.n1397 GND 0.005381f
C1687 CS_BIAS.n1398 GND 0.005381f
C1688 CS_BIAS.n1399 GND 0.010862f
C1689 CS_BIAS.n1400 GND 0.010028f
C1690 CS_BIAS.n1401 GND 0.010028f
C1691 CS_BIAS.n1402 GND 0.005381f
C1692 CS_BIAS.n1403 GND 0.005381f
C1693 CS_BIAS.n1404 GND 0.005381f
C1694 CS_BIAS.n1405 GND 0.010028f
C1695 CS_BIAS.n1406 GND 0.005126f
C1696 CS_BIAS.n1407 GND 0.114251f
C1697 CS_BIAS.n1408 GND 0.009978f
C1698 CS_BIAS.n1409 GND 0.005381f
C1699 CS_BIAS.n1410 GND 0.005381f
C1700 CS_BIAS.n1411 GND 0.005381f
C1701 CS_BIAS.n1412 GND 0.010028f
C1702 CS_BIAS.n1413 GND 0.010028f
C1703 CS_BIAS.n1414 GND 0.010839f
C1704 CS_BIAS.n1415 GND 0.005381f
C1705 CS_BIAS.n1416 GND 0.005381f
C1706 CS_BIAS.n1417 GND 0.005381f
C1707 CS_BIAS.n1418 GND 0.004871f
C1708 CS_BIAS.n1419 GND 0.010839f
C1709 CS_BIAS.n1420 GND 0.010028f
C1710 CS_BIAS.n1421 GND 0.005381f
C1711 CS_BIAS.n1422 GND 0.005381f
C1712 CS_BIAS.n1423 GND 0.005381f
C1713 CS_BIAS.n1424 GND 0.010028f
C1714 CS_BIAS.n1425 GND 0.009978f
C1715 CS_BIAS.n1426 GND 0.114251f
C1716 CS_BIAS.n1427 GND 0.005126f
C1717 CS_BIAS.n1428 GND 0.005381f
C1718 CS_BIAS.n1429 GND 0.005381f
C1719 CS_BIAS.n1430 GND 0.005381f
C1720 CS_BIAS.n1431 GND 0.010028f
C1721 CS_BIAS.n1432 GND 0.010028f
C1722 CS_BIAS.n1433 GND 0.010028f
C1723 CS_BIAS.n1434 GND 0.005381f
C1724 CS_BIAS.n1435 GND 0.005381f
C1725 CS_BIAS.n1436 GND 0.005381f
C1726 CS_BIAS.n1437 GND 0.004717f
C1727 CS_BIAS.n1438 GND 0.005039f
C1728 CS_BIAS.n1439 GND 0.010803f
C1729 CS_BIAS.n1440 GND 0.005381f
C1730 CS_BIAS.n1441 GND 0.005381f
C1731 CS_BIAS.n1442 GND 0.005381f
C1732 CS_BIAS.n1443 GND 0.010028f
C1733 CS_BIAS.n1444 GND 0.010028f
C1734 CS_BIAS.n1445 GND 0.009879f
C1735 CS_BIAS.n1446 GND 0.005381f
C1736 CS_BIAS.n1447 GND 0.005381f
C1737 CS_BIAS.n1448 GND 0.005225f
C1738 CS_BIAS.n1449 GND 0.010028f
C1739 CS_BIAS.n1450 GND 0.010028f
C1740 CS_BIAS.n1451 GND 0.005381f
C1741 CS_BIAS.n1452 GND 0.005381f
C1742 CS_BIAS.n1453 GND 0.005381f
C1743 CS_BIAS.n1454 GND 0.010028f
C1744 CS_BIAS.n1455 GND 0.010872f
C1745 CS_BIAS.n1456 GND 0.004575f
C1746 CS_BIAS.n1457 GND 0.005381f
C1747 CS_BIAS.n1458 GND 0.005381f
C1748 CS_BIAS.n1459 GND 0.005381f
C1749 CS_BIAS.n1460 GND 0.010752f
C1750 CS_BIAS.n1461 GND 0.010028f
C1751 CS_BIAS.n1462 GND 0.010028f
C1752 CS_BIAS.n1463 GND 0.005381f
C1753 CS_BIAS.n1464 GND 0.005381f
C1754 CS_BIAS.n1465 GND 0.005381f
C1755 CS_BIAS.n1466 GND 0.00978f
C1756 CS_BIAS.n1467 GND 0.114251f
C1757 CS_BIAS.n1468 GND 0.005324f
C1758 CS_BIAS.n1469 GND 0.010028f
C1759 CS_BIAS.n1470 GND 0.005381f
C1760 CS_BIAS.n1471 GND 0.005381f
C1761 CS_BIAS.n1472 GND 0.005381f
C1762 CS_BIAS.n1473 GND 0.010028f
C1763 CS_BIAS.n1474 GND 0.010028f
C1764 CS_BIAS.n1475 GND 0.010871f
C1765 CS_BIAS.n1476 GND 0.005381f
C1766 CS_BIAS.n1477 GND 0.005381f
C1767 CS_BIAS.n1478 GND 0.005381f
C1768 CS_BIAS.n1479 GND 0.005421f
C1769 CS_BIAS.n1480 GND 0.010684f
C1770 CS_BIAS.n1481 GND 0.010028f
C1771 CS_BIAS.n1482 GND 0.005381f
C1772 CS_BIAS.n1483 GND 0.005381f
C1773 CS_BIAS.n1484 GND 0.005381f
C1774 CS_BIAS.n1485 GND 0.010028f
C1775 CS_BIAS.n1486 GND 0.009681f
C1776 CS_BIAS.n1487 GND 0.139914f
C1777 CS_BIAS.n1488 GND 0.061282f
C1778 CS_BIAS.n1489 GND 0.053315f
C1779 CS_BIAS.n1490 GND 0.012472f
C1780 CS_BIAS.t42 GND 0.298599f
C1781 CS_BIAS.n1491 GND 0.010028f
C1782 CS_BIAS.n1492 GND 0.005381f
C1783 CS_BIAS.n1493 GND 0.004445f
C1784 CS_BIAS.n1494 GND 0.005381f
C1785 CS_BIAS.n1495 GND 0.010028f
C1786 CS_BIAS.n1496 GND 0.005381f
C1787 CS_BIAS.t90 GND 0.298599f
C1788 CS_BIAS.n1497 GND 0.010028f
C1789 CS_BIAS.n1498 GND 0.005381f
C1790 CS_BIAS.n1499 GND 0.005222f
C1791 CS_BIAS.n1500 GND 0.005381f
C1792 CS_BIAS.n1501 GND 0.010028f
C1793 CS_BIAS.n1502 GND 0.005381f
C1794 CS_BIAS.t73 GND 0.298599f
C1795 CS_BIAS.n1503 GND 0.114251f
C1796 CS_BIAS.n1504 GND 0.005381f
C1797 CS_BIAS.n1505 GND 0.010028f
C1798 CS_BIAS.n1506 GND 0.005381f
C1799 CS_BIAS.n1507 GND 0.010862f
C1800 CS_BIAS.n1508 GND 0.005381f
C1801 CS_BIAS.n1509 GND 0.010028f
C1802 CS_BIAS.n1510 GND 0.005381f
C1803 CS_BIAS.t34 GND 0.298599f
C1804 CS_BIAS.n1511 GND 0.010028f
C1805 CS_BIAS.n1512 GND 0.005381f
C1806 CS_BIAS.n1513 GND 0.004871f
C1807 CS_BIAS.n1514 GND 0.005381f
C1808 CS_BIAS.n1515 GND 0.010028f
C1809 CS_BIAS.n1516 GND 0.005381f
C1810 CS_BIAS.t38 GND 0.298599f
C1811 CS_BIAS.n1517 GND 0.010028f
C1812 CS_BIAS.n1518 GND 0.005381f
C1813 CS_BIAS.n1519 GND 0.004717f
C1814 CS_BIAS.n1520 GND 0.005381f
C1815 CS_BIAS.n1521 GND 0.010028f
C1816 CS_BIAS.n1522 GND 0.005381f
C1817 CS_BIAS.t82 GND 0.298599f
C1818 CS_BIAS.n1523 GND 0.010028f
C1819 CS_BIAS.n1524 GND 0.005381f
C1820 CS_BIAS.n1525 GND 0.010872f
C1821 CS_BIAS.n1526 GND 0.005381f
C1822 CS_BIAS.n1527 GND 0.010028f
C1823 CS_BIAS.n1528 GND 0.005381f
C1824 CS_BIAS.t59 GND 0.298599f
C1825 CS_BIAS.n1529 GND 0.138803f
C1826 CS_BIAS.t64 GND 0.412733f
C1827 CS_BIAS.n1530 GND 0.207253f
C1828 CS_BIAS.n1531 GND 0.051546f
C1829 CS_BIAS.n1532 GND 0.00978f
C1830 CS_BIAS.n1533 GND 0.010028f
C1831 CS_BIAS.n1534 GND 0.010028f
C1832 CS_BIAS.n1535 GND 0.005381f
C1833 CS_BIAS.n1536 GND 0.005381f
C1834 CS_BIAS.n1537 GND 0.005381f
C1835 CS_BIAS.n1538 GND 0.010752f
C1836 CS_BIAS.n1539 GND 0.005222f
C1837 CS_BIAS.n1540 GND 0.004575f
C1838 CS_BIAS.n1541 GND 0.005381f
C1839 CS_BIAS.n1542 GND 0.005381f
C1840 CS_BIAS.n1543 GND 0.005381f
C1841 CS_BIAS.n1544 GND 0.010028f
C1842 CS_BIAS.n1545 GND 0.010028f
C1843 CS_BIAS.n1546 GND 0.010028f
C1844 CS_BIAS.n1547 GND 0.005381f
C1845 CS_BIAS.n1548 GND 0.005381f
C1846 CS_BIAS.n1549 GND 0.005381f
C1847 CS_BIAS.n1550 GND 0.005225f
C1848 CS_BIAS.n1551 GND 0.114251f
C1849 CS_BIAS.n1552 GND 0.009879f
C1850 CS_BIAS.n1553 GND 0.010028f
C1851 CS_BIAS.n1554 GND 0.005381f
C1852 CS_BIAS.n1555 GND 0.005381f
C1853 CS_BIAS.n1556 GND 0.005381f
C1854 CS_BIAS.n1557 GND 0.010028f
C1855 CS_BIAS.n1558 GND 0.010803f
C1856 CS_BIAS.n1559 GND 0.005039f
C1857 CS_BIAS.n1560 GND 0.005381f
C1858 CS_BIAS.n1561 GND 0.005381f
C1859 CS_BIAS.n1562 GND 0.005381f
C1860 CS_BIAS.n1563 GND 0.010862f
C1861 CS_BIAS.n1564 GND 0.010028f
C1862 CS_BIAS.n1565 GND 0.010028f
C1863 CS_BIAS.n1566 GND 0.005381f
C1864 CS_BIAS.n1567 GND 0.005381f
C1865 CS_BIAS.n1568 GND 0.005381f
C1866 CS_BIAS.n1569 GND 0.010028f
C1867 CS_BIAS.n1570 GND 0.005126f
C1868 CS_BIAS.n1571 GND 0.114251f
C1869 CS_BIAS.n1572 GND 0.009978f
C1870 CS_BIAS.n1573 GND 0.005381f
C1871 CS_BIAS.n1574 GND 0.005381f
C1872 CS_BIAS.n1575 GND 0.005381f
C1873 CS_BIAS.n1576 GND 0.010028f
C1874 CS_BIAS.n1577 GND 0.010028f
C1875 CS_BIAS.n1578 GND 0.010839f
C1876 CS_BIAS.n1579 GND 0.005381f
C1877 CS_BIAS.n1580 GND 0.005381f
C1878 CS_BIAS.n1581 GND 0.005381f
C1879 CS_BIAS.n1582 GND 0.004871f
C1880 CS_BIAS.n1583 GND 0.010839f
C1881 CS_BIAS.n1584 GND 0.010028f
C1882 CS_BIAS.n1585 GND 0.005381f
C1883 CS_BIAS.n1586 GND 0.005381f
C1884 CS_BIAS.n1587 GND 0.005381f
C1885 CS_BIAS.n1588 GND 0.010028f
C1886 CS_BIAS.n1589 GND 0.009978f
C1887 CS_BIAS.n1590 GND 0.114251f
C1888 CS_BIAS.n1591 GND 0.005126f
C1889 CS_BIAS.n1592 GND 0.005381f
C1890 CS_BIAS.n1593 GND 0.005381f
C1891 CS_BIAS.n1594 GND 0.005381f
C1892 CS_BIAS.n1595 GND 0.010028f
C1893 CS_BIAS.n1596 GND 0.010028f
C1894 CS_BIAS.n1597 GND 0.010028f
C1895 CS_BIAS.n1598 GND 0.005381f
C1896 CS_BIAS.n1599 GND 0.005381f
C1897 CS_BIAS.n1600 GND 0.005381f
C1898 CS_BIAS.n1601 GND 0.004717f
C1899 CS_BIAS.n1602 GND 0.005039f
C1900 CS_BIAS.n1603 GND 0.010803f
C1901 CS_BIAS.n1604 GND 0.005381f
C1902 CS_BIAS.n1605 GND 0.005381f
C1903 CS_BIAS.n1606 GND 0.005381f
C1904 CS_BIAS.n1607 GND 0.010028f
C1905 CS_BIAS.n1608 GND 0.010028f
C1906 CS_BIAS.n1609 GND 0.009879f
C1907 CS_BIAS.n1610 GND 0.005381f
C1908 CS_BIAS.n1611 GND 0.005381f
C1909 CS_BIAS.n1612 GND 0.005225f
C1910 CS_BIAS.n1613 GND 0.010028f
C1911 CS_BIAS.n1614 GND 0.010028f
C1912 CS_BIAS.n1615 GND 0.005381f
C1913 CS_BIAS.n1616 GND 0.005381f
C1914 CS_BIAS.n1617 GND 0.005381f
C1915 CS_BIAS.n1618 GND 0.010028f
C1916 CS_BIAS.n1619 GND 0.010872f
C1917 CS_BIAS.n1620 GND 0.004575f
C1918 CS_BIAS.n1621 GND 0.005381f
C1919 CS_BIAS.n1622 GND 0.005381f
C1920 CS_BIAS.n1623 GND 0.005381f
C1921 CS_BIAS.n1624 GND 0.010752f
C1922 CS_BIAS.n1625 GND 0.010028f
C1923 CS_BIAS.n1626 GND 0.010028f
C1924 CS_BIAS.n1627 GND 0.005381f
C1925 CS_BIAS.n1628 GND 0.005381f
C1926 CS_BIAS.n1629 GND 0.005381f
C1927 CS_BIAS.n1630 GND 0.00978f
C1928 CS_BIAS.n1631 GND 0.114251f
C1929 CS_BIAS.n1632 GND 0.005324f
C1930 CS_BIAS.n1633 GND 0.010028f
C1931 CS_BIAS.n1634 GND 0.005381f
C1932 CS_BIAS.n1635 GND 0.005381f
C1933 CS_BIAS.n1636 GND 0.005381f
C1934 CS_BIAS.n1637 GND 0.010028f
C1935 CS_BIAS.n1638 GND 0.010028f
C1936 CS_BIAS.n1639 GND 0.010871f
C1937 CS_BIAS.n1640 GND 0.005381f
C1938 CS_BIAS.n1641 GND 0.005381f
C1939 CS_BIAS.n1642 GND 0.005381f
C1940 CS_BIAS.n1643 GND 0.005421f
C1941 CS_BIAS.n1644 GND 0.010684f
C1942 CS_BIAS.n1645 GND 0.010028f
C1943 CS_BIAS.n1646 GND 0.005381f
C1944 CS_BIAS.n1647 GND 0.005381f
C1945 CS_BIAS.n1648 GND 0.005381f
C1946 CS_BIAS.n1649 GND 0.010028f
C1947 CS_BIAS.n1650 GND 0.009681f
C1948 CS_BIAS.n1651 GND 0.139914f
C1949 CS_BIAS.n1652 GND 0.061282f
C1950 CS_BIAS.n1653 GND 0.101596f
C1951 CS_BIAS.n1654 GND 4.8467f
C1952 VN.t7 GND 0.738633f
C1953 VN.n0 GND 0.326436f
C1954 VN.n1 GND 0.013617f
C1955 VN.n2 GND 0.014832f
C1956 VN.n3 GND 0.013617f
C1957 VN.n4 GND 0.021512f
C1958 VN.n5 GND 0.013617f
C1959 VN.t11 GND 0.738633f
C1960 VN.n6 GND 0.273263f
C1961 VN.n7 GND 0.019608f
C1962 VN.n8 GND 0.013617f
C1963 VN.n9 GND 0.024005f
C1964 VN.n10 GND 0.013617f
C1965 VN.t14 GND 0.738633f
C1966 VN.n11 GND 0.273263f
C1967 VN.n12 GND 0.022997f
C1968 VN.n13 GND 0.013617f
C1969 VN.n14 GND 0.025251f
C1970 VN.n15 GND 0.013617f
C1971 VN.t5 GND 0.738633f
C1972 VN.n16 GND 0.025725f
C1973 VN.n17 GND 0.013617f
C1974 VN.n18 GND 0.025251f
C1975 VN.t6 GND 0.908144f
C1976 VN.n19 GND 0.314076f
C1977 VN.t9 GND 0.738633f
C1978 VN.n20 GND 0.3178f
C1979 VN.n21 GND 0.016525f
C1980 VN.n22 GND 0.162936f
C1981 VN.n23 GND 0.013617f
C1982 VN.n24 GND 0.013617f
C1983 VN.n25 GND 0.025251f
C1984 VN.n26 GND 0.019608f
C1985 VN.n27 GND 0.008593f
C1986 VN.n28 GND 0.013617f
C1987 VN.n29 GND 0.013617f
C1988 VN.n30 GND 0.013617f
C1989 VN.n31 GND 0.025251f
C1990 VN.n32 GND 0.024005f
C1991 VN.n33 GND 0.273263f
C1992 VN.n34 GND 0.014032f
C1993 VN.n35 GND 0.013617f
C1994 VN.n36 GND 0.013617f
C1995 VN.n37 GND 0.013617f
C1996 VN.n38 GND 0.025251f
C1997 VN.n39 GND 0.022997f
C1998 VN.n40 GND 0.007933f
C1999 VN.n41 GND 0.013617f
C2000 VN.n42 GND 0.013617f
C2001 VN.n43 GND 0.013617f
C2002 VN.n44 GND 0.025251f
C2003 VN.n45 GND 0.025251f
C2004 VN.n46 GND 0.014032f
C2005 VN.n47 GND 0.013617f
C2006 VN.n48 GND 0.013617f
C2007 VN.n49 GND 0.013617f
C2008 VN.n50 GND 0.025251f
C2009 VN.n51 GND 0.025725f
C2010 VN.n52 GND 0.008593f
C2011 VN.n53 GND 0.013617f
C2012 VN.n54 GND 0.013617f
C2013 VN.n55 GND 0.013617f
C2014 VN.n56 GND 0.025251f
C2015 VN.n57 GND 0.025251f
C2016 VN.n58 GND 0.016525f
C2017 VN.n59 GND 0.013617f
C2018 VN.n60 GND 0.013617f
C2019 VN.n61 GND 0.013617f
C2020 VN.n62 GND 0.025251f
C2021 VN.n63 GND 0.027278f
C2022 VN.n64 GND 0.010657f
C2023 VN.n65 GND 0.013617f
C2024 VN.n66 GND 0.013617f
C2025 VN.n67 GND 0.013617f
C2026 VN.n68 GND 0.026411f
C2027 VN.n69 GND 0.025251f
C2028 VN.n70 GND 0.019018f
C2029 VN.n71 GND 0.021974f
C2030 VN.n72 GND 0.23762f
C2031 VN.t15 GND 0.738633f
C2032 VN.n73 GND 0.326436f
C2033 VN.n74 GND 0.013617f
C2034 VN.n75 GND 0.014832f
C2035 VN.n76 GND 0.013617f
C2036 VN.n77 GND 0.021512f
C2037 VN.n78 GND 0.013617f
C2038 VN.n79 GND 0.019608f
C2039 VN.n80 GND 0.013617f
C2040 VN.n81 GND 0.024005f
C2041 VN.n82 GND 0.013617f
C2042 VN.n83 GND 0.022997f
C2043 VN.n84 GND 0.013617f
C2044 VN.n85 GND 0.025251f
C2045 VN.n86 GND 0.013617f
C2046 VN.t13 GND 0.738633f
C2047 VN.n87 GND 0.025725f
C2048 VN.n88 GND 0.013617f
C2049 VN.n89 GND 0.025251f
C2050 VN.t12 GND 0.908144f
C2051 VN.n90 GND 0.314076f
C2052 VN.t4 GND 0.738633f
C2053 VN.n91 GND 0.3178f
C2054 VN.n92 GND 0.016525f
C2055 VN.n93 GND 0.162936f
C2056 VN.n94 GND 0.013617f
C2057 VN.n95 GND 0.013617f
C2058 VN.n96 GND 0.025251f
C2059 VN.n97 GND 0.019608f
C2060 VN.n98 GND 0.008593f
C2061 VN.n99 GND 0.013617f
C2062 VN.n100 GND 0.013617f
C2063 VN.n101 GND 0.013617f
C2064 VN.n102 GND 0.025251f
C2065 VN.n103 GND 0.024005f
C2066 VN.n104 GND 0.273263f
C2067 VN.n105 GND 0.014032f
C2068 VN.n106 GND 0.013617f
C2069 VN.n107 GND 0.013617f
C2070 VN.n108 GND 0.013617f
C2071 VN.n109 GND 0.025251f
C2072 VN.n110 GND 0.022997f
C2073 VN.n111 GND 0.007933f
C2074 VN.n112 GND 0.013617f
C2075 VN.n113 GND 0.013617f
C2076 VN.n114 GND 0.013617f
C2077 VN.n115 GND 0.025251f
C2078 VN.n116 GND 0.025251f
C2079 VN.t10 GND 0.738633f
C2080 VN.n117 GND 0.273263f
C2081 VN.n118 GND 0.014032f
C2082 VN.n119 GND 0.013617f
C2083 VN.n120 GND 0.013617f
C2084 VN.n121 GND 0.013617f
C2085 VN.n122 GND 0.025251f
C2086 VN.n123 GND 0.025725f
C2087 VN.n124 GND 0.008593f
C2088 VN.n125 GND 0.013617f
C2089 VN.n126 GND 0.013617f
C2090 VN.n127 GND 0.013617f
C2091 VN.n128 GND 0.025251f
C2092 VN.n129 GND 0.025251f
C2093 VN.t8 GND 0.738633f
C2094 VN.n130 GND 0.273263f
C2095 VN.n131 GND 0.016525f
C2096 VN.n132 GND 0.013617f
C2097 VN.n133 GND 0.013617f
C2098 VN.n134 GND 0.013617f
C2099 VN.n135 GND 0.025251f
C2100 VN.n136 GND 0.027278f
C2101 VN.n137 GND 0.010657f
C2102 VN.n138 GND 0.013617f
C2103 VN.n139 GND 0.013617f
C2104 VN.n140 GND 0.013617f
C2105 VN.n141 GND 0.026411f
C2106 VN.n142 GND 0.025251f
C2107 VN.n143 GND 0.019018f
C2108 VN.n144 GND 0.021974f
C2109 VN.n145 GND 0.774716f
C2110 VN.n146 GND 1.00387f
C2111 VN.t0 GND 0.023507f
C2112 VN.t3 GND 0.004198f
C2113 VN.t1 GND 0.004198f
C2114 VN.n147 GND 0.013614f
C2115 VN.n148 GND 0.105685f
C2116 VN.t2 GND 0.023364f
C2117 VN.n149 GND 0.070789f
C2118 VN.n150 GND 4.91094f
C2119 VP.t13 GND 1.03154f
C2120 VP.n0 GND 0.455883f
C2121 VP.n1 GND 0.019017f
C2122 VP.n2 GND 0.020713f
C2123 VP.n3 GND 0.019017f
C2124 VP.n4 GND 0.030042f
C2125 VP.n5 GND 0.019017f
C2126 VP.n6 GND 0.027383f
C2127 VP.n7 GND 0.019017f
C2128 VP.n8 GND 0.033524f
C2129 VP.n9 GND 0.019017f
C2130 VP.n10 GND 0.032116f
C2131 VP.n11 GND 0.019017f
C2132 VP.n12 GND 0.035265f
C2133 VP.n13 GND 0.019017f
C2134 VP.t11 GND 1.03154f
C2135 VP.n14 GND 0.035927f
C2136 VP.n15 GND 0.019017f
C2137 VP.n16 GND 0.035265f
C2138 VP.t9 GND 1.26827f
C2139 VP.n17 GND 0.438622f
C2140 VP.t14 GND 1.03154f
C2141 VP.n18 GND 0.443823f
C2142 VP.n19 GND 0.023078f
C2143 VP.n20 GND 0.227548f
C2144 VP.n21 GND 0.019017f
C2145 VP.n22 GND 0.019017f
C2146 VP.n23 GND 0.035265f
C2147 VP.n24 GND 0.027383f
C2148 VP.n25 GND 0.012f
C2149 VP.n26 GND 0.019017f
C2150 VP.n27 GND 0.019017f
C2151 VP.n28 GND 0.019017f
C2152 VP.n29 GND 0.035265f
C2153 VP.n30 GND 0.033524f
C2154 VP.n31 GND 0.381625f
C2155 VP.n32 GND 0.019596f
C2156 VP.n33 GND 0.019017f
C2157 VP.n34 GND 0.019017f
C2158 VP.n35 GND 0.019017f
C2159 VP.n36 GND 0.035265f
C2160 VP.n37 GND 0.032116f
C2161 VP.n38 GND 0.011078f
C2162 VP.n39 GND 0.019017f
C2163 VP.n40 GND 0.019017f
C2164 VP.n41 GND 0.019017f
C2165 VP.n42 GND 0.035265f
C2166 VP.n43 GND 0.035265f
C2167 VP.t8 GND 1.03154f
C2168 VP.n44 GND 0.381625f
C2169 VP.n45 GND 0.019596f
C2170 VP.n46 GND 0.019017f
C2171 VP.n47 GND 0.019017f
C2172 VP.n48 GND 0.019017f
C2173 VP.n49 GND 0.035265f
C2174 VP.n50 GND 0.035927f
C2175 VP.n51 GND 0.012f
C2176 VP.n52 GND 0.019017f
C2177 VP.n53 GND 0.019017f
C2178 VP.n54 GND 0.019017f
C2179 VP.n55 GND 0.035265f
C2180 VP.n56 GND 0.035265f
C2181 VP.t7 GND 1.03154f
C2182 VP.n57 GND 0.381625f
C2183 VP.n58 GND 0.023078f
C2184 VP.n59 GND 0.019017f
C2185 VP.n60 GND 0.019017f
C2186 VP.n61 GND 0.019017f
C2187 VP.n62 GND 0.035265f
C2188 VP.n63 GND 0.038095f
C2189 VP.n64 GND 0.014883f
C2190 VP.n65 GND 0.019017f
C2191 VP.n66 GND 0.019017f
C2192 VP.n67 GND 0.019017f
C2193 VP.n68 GND 0.036884f
C2194 VP.n69 GND 0.035265f
C2195 VP.n70 GND 0.02656f
C2196 VP.n71 GND 0.030688f
C2197 VP.n72 GND 0.336603f
C2198 VP.t6 GND 1.03154f
C2199 VP.n73 GND 0.455883f
C2200 VP.n74 GND 0.019017f
C2201 VP.n75 GND 0.020713f
C2202 VP.n76 GND 0.019017f
C2203 VP.n77 GND 0.030042f
C2204 VP.n78 GND 0.019017f
C2205 VP.t12 GND 1.03154f
C2206 VP.n79 GND 0.381625f
C2207 VP.n80 GND 0.027383f
C2208 VP.n81 GND 0.019017f
C2209 VP.n82 GND 0.033524f
C2210 VP.n83 GND 0.019017f
C2211 VP.t15 GND 1.03154f
C2212 VP.n84 GND 0.381625f
C2213 VP.n85 GND 0.032116f
C2214 VP.n86 GND 0.019017f
C2215 VP.n87 GND 0.035265f
C2216 VP.n88 GND 0.019017f
C2217 VP.t4 GND 1.03154f
C2218 VP.n89 GND 0.035927f
C2219 VP.n90 GND 0.019017f
C2220 VP.n91 GND 0.035265f
C2221 VP.t5 GND 1.26827f
C2222 VP.n92 GND 0.438623f
C2223 VP.t10 GND 1.03154f
C2224 VP.n93 GND 0.443823f
C2225 VP.n94 GND 0.023078f
C2226 VP.n95 GND 0.227548f
C2227 VP.n96 GND 0.019017f
C2228 VP.n97 GND 0.019017f
C2229 VP.n98 GND 0.035265f
C2230 VP.n99 GND 0.027383f
C2231 VP.n100 GND 0.012f
C2232 VP.n101 GND 0.019017f
C2233 VP.n102 GND 0.019017f
C2234 VP.n103 GND 0.019017f
C2235 VP.n104 GND 0.035265f
C2236 VP.n105 GND 0.033524f
C2237 VP.n106 GND 0.381625f
C2238 VP.n107 GND 0.019596f
C2239 VP.n108 GND 0.019017f
C2240 VP.n109 GND 0.019017f
C2241 VP.n110 GND 0.019017f
C2242 VP.n111 GND 0.035265f
C2243 VP.n112 GND 0.032116f
C2244 VP.n113 GND 0.011078f
C2245 VP.n114 GND 0.019017f
C2246 VP.n115 GND 0.019017f
C2247 VP.n116 GND 0.019017f
C2248 VP.n117 GND 0.035265f
C2249 VP.n118 GND 0.035265f
C2250 VP.n119 GND 0.019596f
C2251 VP.n120 GND 0.019017f
C2252 VP.n121 GND 0.019017f
C2253 VP.n122 GND 0.019017f
C2254 VP.n123 GND 0.035265f
C2255 VP.n124 GND 0.035927f
C2256 VP.n125 GND 0.012f
C2257 VP.n126 GND 0.019017f
C2258 VP.n127 GND 0.019017f
C2259 VP.n128 GND 0.019017f
C2260 VP.n129 GND 0.035265f
C2261 VP.n130 GND 0.035265f
C2262 VP.n131 GND 0.023078f
C2263 VP.n132 GND 0.019017f
C2264 VP.n133 GND 0.019017f
C2265 VP.n134 GND 0.019017f
C2266 VP.n135 GND 0.035265f
C2267 VP.n136 GND 0.038095f
C2268 VP.n137 GND 0.014883f
C2269 VP.n138 GND 0.019017f
C2270 VP.n139 GND 0.019017f
C2271 VP.n140 GND 0.019017f
C2272 VP.n141 GND 0.036884f
C2273 VP.n142 GND 0.035265f
C2274 VP.n143 GND 0.02656f
C2275 VP.n144 GND 0.030688f
C2276 VP.n145 GND 1.08936f
C2277 VP.n146 GND 1.40982f
C2278 VP.t1 GND 0.032828f
C2279 VP.t3 GND 0.005862f
C2280 VP.t2 GND 0.005862f
C2281 VP.n147 GND 0.019012f
C2282 VP.n148 GND 0.147595f
C2283 VP.t0 GND 0.032629f
C2284 VP.n149 GND 0.088545f
C2285 VP.n150 GND 3.60978f
C2286 VDD.t79 GND 0.020633f
C2287 VDD.t75 GND 0.020633f
C2288 VDD.n0 GND 0.112055f
C2289 VDD.t90 GND 0.020633f
C2290 VDD.t161 GND 0.020633f
C2291 VDD.n1 GND 0.103927f
C2292 VDD.n2 GND 0.980344f
C2293 VDD.t95 GND 0.020633f
C2294 VDD.t97 GND 0.020633f
C2295 VDD.n3 GND 0.103927f
C2296 VDD.n4 GND 0.514901f
C2297 VDD.t101 GND 0.020633f
C2298 VDD.t86 GND 0.020633f
C2299 VDD.n5 GND 0.103927f
C2300 VDD.n6 GND 0.42656f
C2301 VDD.t88 GND 0.020633f
C2302 VDD.t163 GND 0.020633f
C2303 VDD.n7 GND 0.112055f
C2304 VDD.t159 GND 0.020633f
C2305 VDD.t1 GND 0.020633f
C2306 VDD.n8 GND 0.103927f
C2307 VDD.n9 GND 0.980344f
C2308 VDD.t83 GND 0.020633f
C2309 VDD.t93 GND 0.020633f
C2310 VDD.n10 GND 0.103927f
C2311 VDD.n11 GND 0.514901f
C2312 VDD.t77 GND 0.020633f
C2313 VDD.t99 GND 0.020633f
C2314 VDD.n12 GND 0.103927f
C2315 VDD.n13 GND 0.42656f
C2316 VDD.n14 GND 0.31257f
C2317 VDD.n15 GND 3.32598f
C2318 VDD.t154 GND 0.016539f
C2319 VDD.t143 GND 0.016539f
C2320 VDD.n16 GND 0.069944f
C2321 VDD.t109 GND 0.016539f
C2322 VDD.t125 GND 0.016539f
C2323 VDD.n17 GND 0.062673f
C2324 VDD.n18 GND 0.855534f
C2325 VDD.t147 GND 0.016539f
C2326 VDD.t140 GND 0.016539f
C2327 VDD.n19 GND 0.062673f
C2328 VDD.n20 GND 0.429343f
C2329 VDD.t106 GND 0.087299f
C2330 VDD.n21 GND 0.318501f
C2331 VDD.t149 GND 0.016539f
C2332 VDD.t142 GND 0.016539f
C2333 VDD.n22 GND 0.069944f
C2334 VDD.t108 GND 0.016539f
C2335 VDD.t123 GND 0.016539f
C2336 VDD.n23 GND 0.062673f
C2337 VDD.n24 GND 0.855534f
C2338 VDD.t145 GND 0.016539f
C2339 VDD.t139 GND 0.016539f
C2340 VDD.n25 GND 0.062673f
C2341 VDD.n26 GND 0.429343f
C2342 VDD.t105 GND 0.087299f
C2343 VDD.n27 GND 0.301905f
C2344 VDD.n28 GND 0.267638f
C2345 VDD.t119 GND 0.016539f
C2346 VDD.t151 GND 0.016539f
C2347 VDD.n29 GND 0.069944f
C2348 VDD.t146 GND 0.016539f
C2349 VDD.t135 GND 0.016539f
C2350 VDD.n30 GND 0.062673f
C2351 VDD.n31 GND 0.855534f
C2352 VDD.t129 GND 0.016539f
C2353 VDD.t157 GND 0.016539f
C2354 VDD.n32 GND 0.062673f
C2355 VDD.n33 GND 0.429343f
C2356 VDD.t152 GND 0.087299f
C2357 VDD.n34 GND 0.301905f
C2358 VDD.n35 GND 0.423499f
C2359 VDD.n36 GND 0.005144f
C2360 VDD.n37 GND 0.006693f
C2361 VDD.n38 GND 0.005387f
C2362 VDD.n39 GND 0.006693f
C2363 VDD.n40 GND 0.005387f
C2364 VDD.n41 GND 0.006693f
C2365 VDD.n42 GND 0.358495f
C2366 VDD.n43 GND 0.006693f
C2367 VDD.n44 GND 0.006693f
C2368 VDD.n45 GND 0.006693f
C2369 VDD.n46 GND 0.477993f
C2370 VDD.n47 GND 0.006693f
C2371 VDD.n48 GND 0.006693f
C2372 VDD.n49 GND 0.006693f
C2373 VDD.n50 GND 0.006693f
C2374 VDD.n51 GND 0.006693f
C2375 VDD.n52 GND 0.005387f
C2376 VDD.n53 GND 0.006693f
C2377 VDD.n54 GND 0.006693f
C2378 VDD.n55 GND 0.006693f
C2379 VDD.n56 GND 0.006693f
C2380 VDD.n57 GND 0.477993f
C2381 VDD.n58 GND 0.006693f
C2382 VDD.n59 GND 0.006693f
C2383 VDD.n60 GND 0.006693f
C2384 VDD.n61 GND 0.006693f
C2385 VDD.n62 GND 0.006693f
C2386 VDD.n63 GND 0.005387f
C2387 VDD.n64 GND 0.006693f
C2388 VDD.n65 GND 0.006693f
C2389 VDD.n66 GND 0.006693f
C2390 VDD.n67 GND 0.006693f
C2391 VDD.t128 GND 0.238997f
C2392 VDD.n68 GND 0.006693f
C2393 VDD.n69 GND 0.006693f
C2394 VDD.n70 GND 0.006693f
C2395 VDD.n71 GND 0.006693f
C2396 VDD.n72 GND 0.006693f
C2397 VDD.n73 GND 0.005387f
C2398 VDD.n74 GND 0.006693f
C2399 VDD.n75 GND 0.286796f
C2400 VDD.n76 GND 0.006693f
C2401 VDD.n77 GND 0.006693f
C2402 VDD.n78 GND 0.006693f
C2403 VDD.n79 GND 0.477993f
C2404 VDD.n80 GND 0.006693f
C2405 VDD.n81 GND 0.006693f
C2406 VDD.n82 GND 0.006693f
C2407 VDD.n83 GND 0.006693f
C2408 VDD.n84 GND 0.006693f
C2409 VDD.n85 GND 0.005387f
C2410 VDD.n86 GND 0.006693f
C2411 VDD.n87 GND 0.006693f
C2412 VDD.n88 GND 0.006693f
C2413 VDD.n89 GND 0.006693f
C2414 VDD.n90 GND 0.477993f
C2415 VDD.n91 GND 0.006693f
C2416 VDD.n92 GND 0.006693f
C2417 VDD.n93 GND 0.006693f
C2418 VDD.n94 GND 0.006693f
C2419 VDD.n95 GND 0.006693f
C2420 VDD.n96 GND 0.005387f
C2421 VDD.n97 GND 0.006693f
C2422 VDD.n98 GND 0.006693f
C2423 VDD.n99 GND 0.006693f
C2424 VDD.n100 GND 0.006693f
C2425 VDD.n101 GND 0.262896f
C2426 VDD.n102 GND 0.006693f
C2427 VDD.n103 GND 0.006693f
C2428 VDD.n104 GND 0.006693f
C2429 VDD.n105 GND 0.006693f
C2430 VDD.n106 GND 0.006693f
C2431 VDD.n107 GND 0.005387f
C2432 VDD.n108 GND 0.006693f
C2433 VDD.t138 GND 0.238997f
C2434 VDD.n109 GND 0.006693f
C2435 VDD.n110 GND 0.006693f
C2436 VDD.n111 GND 0.006693f
C2437 VDD.n112 GND 0.477993f
C2438 VDD.n113 GND 0.006693f
C2439 VDD.n114 GND 0.006693f
C2440 VDD.n115 GND 0.006693f
C2441 VDD.n116 GND 0.006693f
C2442 VDD.n117 GND 0.006693f
C2443 VDD.n118 GND 0.005387f
C2444 VDD.n119 GND 0.006693f
C2445 VDD.n120 GND 0.006693f
C2446 VDD.n121 GND 0.006693f
C2447 VDD.n122 GND 0.006693f
C2448 VDD.n123 GND 0.477993f
C2449 VDD.n124 GND 0.006693f
C2450 VDD.n125 GND 0.006693f
C2451 VDD.n126 GND 0.006693f
C2452 VDD.n127 GND 0.006693f
C2453 VDD.n128 GND 0.006693f
C2454 VDD.n129 GND 0.005387f
C2455 VDD.n130 GND 0.006693f
C2456 VDD.n131 GND 0.006693f
C2457 VDD.n132 GND 0.006693f
C2458 VDD.n133 GND 0.006693f
C2459 VDD.n134 GND 0.334595f
C2460 VDD.n135 GND 0.006693f
C2461 VDD.n136 GND 0.006693f
C2462 VDD.n137 GND 0.006693f
C2463 VDD.n138 GND 0.006693f
C2464 VDD.n139 GND 0.006693f
C2465 VDD.n140 GND 0.005387f
C2466 VDD.n141 GND 0.006693f
C2467 VDD.t104 GND 0.238997f
C2468 VDD.n142 GND 0.006693f
C2469 VDD.n143 GND 0.006693f
C2470 VDD.n144 GND 0.006693f
C2471 VDD.n145 GND 0.477993f
C2472 VDD.n146 GND 0.006693f
C2473 VDD.n147 GND 0.006693f
C2474 VDD.n148 GND 0.006693f
C2475 VDD.n149 GND 0.006693f
C2476 VDD.n150 GND 0.006693f
C2477 VDD.n151 GND 0.005387f
C2478 VDD.n152 GND 0.006693f
C2479 VDD.n153 GND 0.006693f
C2480 VDD.n154 GND 0.006693f
C2481 VDD.n155 GND 0.006693f
C2482 VDD.n156 GND 0.477993f
C2483 VDD.n157 GND 0.006693f
C2484 VDD.n158 GND 0.006693f
C2485 VDD.n159 GND 0.006693f
C2486 VDD.n160 GND 0.006693f
C2487 VDD.n161 GND 0.006693f
C2488 VDD.n162 GND 0.005387f
C2489 VDD.n163 GND 0.006693f
C2490 VDD.n164 GND 0.006693f
C2491 VDD.n165 GND 0.006693f
C2492 VDD.n166 GND 0.006693f
C2493 VDD.n167 GND 0.477993f
C2494 VDD.n168 GND 0.006693f
C2495 VDD.n169 GND 0.006693f
C2496 VDD.n170 GND 0.006693f
C2497 VDD.n171 GND 0.006693f
C2498 VDD.n172 GND 0.006693f
C2499 VDD.n173 GND 0.005387f
C2500 VDD.n174 GND 0.006693f
C2501 VDD.n175 GND 0.006693f
C2502 VDD.n176 GND 0.006693f
C2503 VDD.n177 GND 0.006693f
C2504 VDD.t9 GND 0.238997f
C2505 VDD.n178 GND 0.006693f
C2506 VDD.n179 GND 0.006693f
C2507 VDD.n180 GND 0.006693f
C2508 VDD.n181 GND 0.006693f
C2509 VDD.n182 GND 0.006693f
C2510 VDD.n183 GND 0.005387f
C2511 VDD.n184 GND 0.006693f
C2512 VDD.n185 GND 0.348935f
C2513 VDD.n186 GND 0.006693f
C2514 VDD.n187 GND 0.006693f
C2515 VDD.n188 GND 0.006693f
C2516 VDD.n189 GND 0.477993f
C2517 VDD.n190 GND 0.006693f
C2518 VDD.n191 GND 0.006693f
C2519 VDD.n192 GND 0.006693f
C2520 VDD.n193 GND 0.006693f
C2521 VDD.n194 GND 0.006693f
C2522 VDD.n195 GND 0.004471f
C2523 VDD.n196 GND 0.01598f
C2524 VDD.n197 GND 0.006693f
C2525 VDD.n198 GND 0.01598f
C2526 VDD.n217 GND 0.006693f
C2527 VDD.t13 GND 0.118593f
C2528 VDD.t12 GND 0.540868f
C2529 VDD.n218 GND 0.08957f
C2530 VDD.t14 GND 0.077791f
C2531 VDD.n219 GND 0.092102f
C2532 VDD.n220 GND 0.007407f
C2533 VDD.n221 GND 0.006693f
C2534 VDD.n222 GND 0.005387f
C2535 VDD.n223 GND 0.006693f
C2536 VDD.n224 GND 0.005387f
C2537 VDD.n225 GND 0.006693f
C2538 VDD.n226 GND 0.005387f
C2539 VDD.n227 GND 0.006693f
C2540 VDD.t10 GND 0.118593f
C2541 VDD.t8 GND 0.540868f
C2542 VDD.n228 GND 0.08957f
C2543 VDD.t11 GND 0.077791f
C2544 VDD.n229 GND 0.092102f
C2545 VDD.n230 GND 0.007407f
C2546 VDD.n231 GND 0.005387f
C2547 VDD.n232 GND 0.006693f
C2548 VDD.n233 GND 0.005387f
C2549 VDD.n234 GND 0.006693f
C2550 VDD.n235 GND 0.005387f
C2551 VDD.n236 GND 0.006693f
C2552 VDD.t19 GND 0.118593f
C2553 VDD.t18 GND 0.540868f
C2554 VDD.n237 GND 0.08957f
C2555 VDD.t20 GND 0.077791f
C2556 VDD.n238 GND 0.092102f
C2557 VDD.n239 GND 0.005387f
C2558 VDD.n240 GND 0.006693f
C2559 VDD.n241 GND 0.005387f
C2560 VDD.n242 GND 0.006693f
C2561 VDD.n243 GND 0.005387f
C2562 VDD.n244 GND 0.01598f
C2563 VDD.n245 GND 0.016349f
C2564 VDD.n246 GND 0.004471f
C2565 VDD.n247 GND 0.016349f
C2566 VDD.n248 GND 0.006693f
C2567 VDD.n249 GND 0.006693f
C2568 VDD.n250 GND 0.006693f
C2569 VDD.n251 GND 0.006693f
C2570 VDD.n252 GND 0.005387f
C2571 VDD.n253 GND 0.005387f
C2572 VDD.n254 GND 0.006693f
C2573 VDD.n255 GND 0.006693f
C2574 VDD.n256 GND 0.005387f
C2575 VDD.n257 GND 0.006693f
C2576 VDD.n258 GND 0.006693f
C2577 VDD.n259 GND 0.006693f
C2578 VDD.n260 GND 0.006693f
C2579 VDD.n261 GND 0.006693f
C2580 VDD.n262 GND 0.005387f
C2581 VDD.n263 GND 0.005387f
C2582 VDD.n264 GND 0.006693f
C2583 VDD.n265 GND 0.006693f
C2584 VDD.n266 GND 0.005387f
C2585 VDD.n267 GND 0.006693f
C2586 VDD.n268 GND 0.006693f
C2587 VDD.n269 GND 0.006693f
C2588 VDD.n270 GND 0.006693f
C2589 VDD.n271 GND 0.006693f
C2590 VDD.n272 GND 0.002721f
C2591 VDD.n273 GND 0.007407f
C2592 VDD.n274 GND 0.003582f
C2593 VDD.n275 GND 0.006693f
C2594 VDD.n276 GND 0.006693f
C2595 VDD.n277 GND 0.005387f
C2596 VDD.n278 GND 0.006693f
C2597 VDD.n279 GND 0.006693f
C2598 VDD.n280 GND 0.006693f
C2599 VDD.n281 GND 0.006693f
C2600 VDD.n282 GND 0.006693f
C2601 VDD.n283 GND 0.005387f
C2602 VDD.n284 GND 0.005387f
C2603 VDD.n285 GND 0.006693f
C2604 VDD.n286 GND 0.006693f
C2605 VDD.n287 GND 0.005387f
C2606 VDD.n288 GND 0.006693f
C2607 VDD.n289 GND 0.006693f
C2608 VDD.n290 GND 0.006693f
C2609 VDD.n291 GND 0.006693f
C2610 VDD.n292 GND 0.006693f
C2611 VDD.n293 GND 0.005387f
C2612 VDD.n294 GND 0.005387f
C2613 VDD.n295 GND 0.006693f
C2614 VDD.n296 GND 0.006693f
C2615 VDD.n297 GND 0.005387f
C2616 VDD.n298 GND 0.006693f
C2617 VDD.n299 GND 0.006693f
C2618 VDD.n300 GND 0.006693f
C2619 VDD.n301 GND 0.006693f
C2620 VDD.n302 GND 0.006693f
C2621 VDD.n303 GND 0.005387f
C2622 VDD.n304 GND 0.002721f
C2623 VDD.n305 GND 0.006693f
C2624 VDD.n306 GND 0.006693f
C2625 VDD.n307 GND 0.003582f
C2626 VDD.n308 GND 0.006693f
C2627 VDD.n309 GND 0.006693f
C2628 VDD.n310 GND 0.006693f
C2629 VDD.n311 GND 0.006693f
C2630 VDD.n312 GND 0.006693f
C2631 VDD.n313 GND 0.005387f
C2632 VDD.n314 GND 0.005387f
C2633 VDD.n315 GND 0.006693f
C2634 VDD.n316 GND 0.006693f
C2635 VDD.n317 GND 0.005387f
C2636 VDD.n318 GND 0.006693f
C2637 VDD.n319 GND 0.006693f
C2638 VDD.n320 GND 0.006693f
C2639 VDD.n321 GND 0.006693f
C2640 VDD.n322 GND 0.006693f
C2641 VDD.n323 GND 0.005387f
C2642 VDD.n324 GND 0.005387f
C2643 VDD.n325 GND 0.006693f
C2644 VDD.n326 GND 0.006693f
C2645 VDD.n327 GND 0.005387f
C2646 VDD.n328 GND 0.006693f
C2647 VDD.n329 GND 0.006693f
C2648 VDD.n330 GND 0.006693f
C2649 VDD.n331 GND 0.006693f
C2650 VDD.n332 GND 0.006693f
C2651 VDD.n333 GND 0.005387f
C2652 VDD.n334 GND 0.006693f
C2653 VDD.n335 GND 0.005387f
C2654 VDD.n336 GND 0.002721f
C2655 VDD.n337 GND 0.006693f
C2656 VDD.n338 GND 0.006693f
C2657 VDD.n339 GND 0.005387f
C2658 VDD.n340 GND 0.006693f
C2659 VDD.n341 GND 0.005387f
C2660 VDD.n342 GND 0.006693f
C2661 VDD.n343 GND 0.005387f
C2662 VDD.n344 GND 0.006693f
C2663 VDD.n345 GND 0.005387f
C2664 VDD.n346 GND 0.006693f
C2665 VDD.n347 GND 0.005387f
C2666 VDD.n348 GND 0.006693f
C2667 VDD.n349 GND 0.005387f
C2668 VDD.n350 GND 0.006693f
C2669 VDD.n351 GND 0.005387f
C2670 VDD.n352 GND 0.006693f
C2671 VDD.n353 GND 0.005387f
C2672 VDD.n354 GND 0.006693f
C2673 VDD.n355 GND 0.005387f
C2674 VDD.n356 GND 0.006693f
C2675 VDD.n357 GND 0.005387f
C2676 VDD.n358 GND 0.006693f
C2677 VDD.n359 GND 0.005387f
C2678 VDD.n360 GND 0.006693f
C2679 VDD.n361 GND 0.005387f
C2680 VDD.n362 GND 0.006693f
C2681 VDD.n363 GND 0.005387f
C2682 VDD.n364 GND 0.006693f
C2683 VDD.n365 GND 0.005387f
C2684 VDD.n366 GND 0.006693f
C2685 VDD.n367 GND 0.005387f
C2686 VDD.n368 GND 0.006693f
C2687 VDD.n369 GND 0.006693f
C2688 VDD.n370 GND 0.477993f
C2689 VDD.t122 GND 0.238997f
C2690 VDD.n371 GND 0.006693f
C2691 VDD.n372 GND 0.005387f
C2692 VDD.n373 GND 0.006693f
C2693 VDD.n374 GND 0.005387f
C2694 VDD.n375 GND 0.006693f
C2695 VDD.n376 GND 0.477993f
C2696 VDD.n377 GND 0.006693f
C2697 VDD.n378 GND 0.005387f
C2698 VDD.n379 GND 0.006693f
C2699 VDD.n380 GND 0.005387f
C2700 VDD.n381 GND 0.006693f
C2701 VDD.n382 GND 0.477993f
C2702 VDD.n383 GND 0.006693f
C2703 VDD.n384 GND 0.005387f
C2704 VDD.n385 GND 0.006693f
C2705 VDD.n386 GND 0.005387f
C2706 VDD.n387 GND 0.006693f
C2707 VDD.n388 GND 0.477993f
C2708 VDD.n389 GND 0.006693f
C2709 VDD.n390 GND 0.005387f
C2710 VDD.n391 GND 0.006693f
C2711 VDD.n392 GND 0.005387f
C2712 VDD.n393 GND 0.006693f
C2713 VDD.n394 GND 0.477993f
C2714 VDD.n395 GND 0.006693f
C2715 VDD.n396 GND 0.005387f
C2716 VDD.n397 GND 0.006693f
C2717 VDD.n398 GND 0.005387f
C2718 VDD.n399 GND 0.006693f
C2719 VDD.t107 GND 0.238997f
C2720 VDD.n400 GND 0.006693f
C2721 VDD.n401 GND 0.005387f
C2722 VDD.n402 GND 0.006693f
C2723 VDD.n403 GND 0.005387f
C2724 VDD.n404 GND 0.006693f
C2725 VDD.n405 GND 0.477993f
C2726 VDD.n406 GND 0.286796f
C2727 VDD.n407 GND 0.006693f
C2728 VDD.n408 GND 0.005387f
C2729 VDD.n409 GND 0.006693f
C2730 VDD.n410 GND 0.005387f
C2731 VDD.n411 GND 0.006693f
C2732 VDD.n412 GND 0.477993f
C2733 VDD.n413 GND 0.006693f
C2734 VDD.n414 GND 0.005387f
C2735 VDD.n415 GND 0.006693f
C2736 VDD.n416 GND 0.005387f
C2737 VDD.n417 GND 0.006693f
C2738 VDD.n418 GND 0.477993f
C2739 VDD.n419 GND 0.006693f
C2740 VDD.n420 GND 0.005387f
C2741 VDD.n421 GND 0.006693f
C2742 VDD.n422 GND 0.005387f
C2743 VDD.n423 GND 0.006693f
C2744 VDD.n424 GND 0.477993f
C2745 VDD.n425 GND 0.006693f
C2746 VDD.n426 GND 0.005387f
C2747 VDD.n427 GND 0.006693f
C2748 VDD.n428 GND 0.005387f
C2749 VDD.n429 GND 0.006693f
C2750 VDD.n430 GND 0.477993f
C2751 VDD.n431 GND 0.006693f
C2752 VDD.n432 GND 0.005387f
C2753 VDD.n433 GND 0.006693f
C2754 VDD.n434 GND 0.005387f
C2755 VDD.n435 GND 0.006693f
C2756 VDD.n436 GND 0.262896f
C2757 VDD.n437 GND 0.006693f
C2758 VDD.n438 GND 0.005387f
C2759 VDD.n439 GND 0.006693f
C2760 VDD.n440 GND 0.005387f
C2761 VDD.n441 GND 0.006693f
C2762 VDD.n442 GND 0.477993f
C2763 VDD.t141 GND 0.238997f
C2764 VDD.n443 GND 0.006693f
C2765 VDD.n444 GND 0.005387f
C2766 VDD.n445 GND 0.006693f
C2767 VDD.n446 GND 0.005387f
C2768 VDD.n447 GND 0.006693f
C2769 VDD.n448 GND 0.477993f
C2770 VDD.n449 GND 0.006693f
C2771 VDD.n450 GND 0.005387f
C2772 VDD.n451 GND 0.006693f
C2773 VDD.n452 GND 0.005387f
C2774 VDD.n453 GND 0.006693f
C2775 VDD.n454 GND 0.477993f
C2776 VDD.n455 GND 0.006693f
C2777 VDD.n456 GND 0.005387f
C2778 VDD.n457 GND 0.006693f
C2779 VDD.n458 GND 0.005387f
C2780 VDD.n459 GND 0.006693f
C2781 VDD.n460 GND 0.477993f
C2782 VDD.n461 GND 0.006693f
C2783 VDD.n462 GND 0.005387f
C2784 VDD.n463 GND 0.006693f
C2785 VDD.n464 GND 0.005387f
C2786 VDD.n465 GND 0.006693f
C2787 VDD.n466 GND 0.477993f
C2788 VDD.n467 GND 0.006693f
C2789 VDD.n468 GND 0.005387f
C2790 VDD.n469 GND 0.006693f
C2791 VDD.n470 GND 0.005387f
C2792 VDD.n471 GND 0.006693f
C2793 VDD.n472 GND 0.334595f
C2794 VDD.n473 GND 0.006693f
C2795 VDD.n474 GND 0.005387f
C2796 VDD.n475 GND 0.006693f
C2797 VDD.n476 GND 0.005387f
C2798 VDD.n477 GND 0.006693f
C2799 VDD.n478 GND 0.477993f
C2800 VDD.t118 GND 0.238997f
C2801 VDD.n479 GND 0.006693f
C2802 VDD.n480 GND 0.005387f
C2803 VDD.n481 GND 0.006693f
C2804 VDD.n482 GND 0.005387f
C2805 VDD.n483 GND 0.006693f
C2806 VDD.n484 GND 0.477993f
C2807 VDD.n485 GND 0.006693f
C2808 VDD.n486 GND 0.005387f
C2809 VDD.n487 GND 0.006693f
C2810 VDD.n488 GND 0.005387f
C2811 VDD.n489 GND 0.006693f
C2812 VDD.n490 GND 0.477993f
C2813 VDD.n491 GND 0.006693f
C2814 VDD.n492 GND 0.005387f
C2815 VDD.n493 GND 0.006693f
C2816 VDD.n494 GND 0.005387f
C2817 VDD.n495 GND 0.006693f
C2818 VDD.n496 GND 0.477993f
C2819 VDD.n497 GND 0.006693f
C2820 VDD.n498 GND 0.005387f
C2821 VDD.n499 GND 0.006693f
C2822 VDD.n500 GND 0.005387f
C2823 VDD.n501 GND 0.006693f
C2824 VDD.n502 GND 0.477993f
C2825 VDD.n503 GND 0.006693f
C2826 VDD.n504 GND 0.005387f
C2827 VDD.n505 GND 0.006693f
C2828 VDD.n506 GND 0.005387f
C2829 VDD.n507 GND 0.006693f
C2830 VDD.n508 GND 0.477993f
C2831 VDD.n509 GND 0.006693f
C2832 VDD.n510 GND 0.005387f
C2833 VDD.n511 GND 0.006693f
C2834 VDD.n512 GND 0.005387f
C2835 VDD.n513 GND 0.006693f
C2836 VDD.n514 GND 0.477993f
C2837 VDD.n515 GND 0.006693f
C2838 VDD.n516 GND 0.005387f
C2839 VDD.n517 GND 0.006693f
C2840 VDD.n518 GND 0.005387f
C2841 VDD.n519 GND 0.006693f
C2842 VDD.t29 GND 0.238997f
C2843 VDD.n520 GND 0.006693f
C2844 VDD.n521 GND 0.005387f
C2845 VDD.n522 GND 0.006693f
C2846 VDD.n523 GND 0.005387f
C2847 VDD.n524 GND 0.006693f
C2848 VDD.n525 GND 0.477993f
C2849 VDD.n526 GND 0.348935f
C2850 VDD.n527 GND 0.006693f
C2851 VDD.n528 GND 0.005387f
C2852 VDD.n529 GND 0.006693f
C2853 VDD.n530 GND 0.005387f
C2854 VDD.n531 GND 0.006693f
C2855 VDD.n532 GND 0.477993f
C2856 VDD.n533 GND 0.006693f
C2857 VDD.n534 GND 0.005387f
C2858 VDD.n535 GND 0.013326f
C2859 VDD.n536 GND 0.004471f
C2860 VDD.n537 GND 0.01598f
C2861 VDD.n538 GND 0.70265f
C2862 VDD.n539 GND 0.01598f
C2863 VDD.n540 GND 0.004471f
C2864 VDD.n541 GND 0.066999f
C2865 VDD.n542 GND 1.90429f
C2866 VDD.n543 GND 0.016349f
C2867 VDD.n544 GND 0.002108f
C2868 VDD.n545 GND 0.005387f
C2869 VDD.n546 GND 0.006693f
C2870 VDD.t80 GND 7.53078f
C2871 VDD.n564 GND 0.006693f
C2872 VDD.t55 GND 0.118593f
C2873 VDD.t53 GND 0.540868f
C2874 VDD.n565 GND 0.08957f
C2875 VDD.t54 GND 0.077791f
C2876 VDD.n566 GND 0.092102f
C2877 VDD.n567 GND 0.007407f
C2878 VDD.n568 GND 0.003347f
C2879 VDD.n569 GND 0.005387f
C2880 VDD.n570 GND 0.003347f
C2881 VDD.n571 GND 0.005387f
C2882 VDD.n572 GND 0.003347f
C2883 VDD.n573 GND 0.005387f
C2884 VDD.n574 GND 0.003347f
C2885 VDD.t52 GND 0.118593f
C2886 VDD.t50 GND 0.540868f
C2887 VDD.n575 GND 0.08957f
C2888 VDD.t51 GND 0.077791f
C2889 VDD.n576 GND 0.092102f
C2890 VDD.n577 GND 0.005387f
C2891 VDD.n578 GND 0.00251f
C2892 VDD.n579 GND 0.005387f
C2893 VDD.n580 GND 0.003347f
C2894 VDD.n581 GND 0.005387f
C2895 VDD.n582 GND 0.003347f
C2896 VDD.t31 GND 0.118593f
C2897 VDD.t28 GND 0.540868f
C2898 VDD.n583 GND 0.08957f
C2899 VDD.t30 GND 0.077791f
C2900 VDD.n584 GND 0.092102f
C2901 VDD.n585 GND 0.007407f
C2902 VDD.n586 GND 0.005387f
C2903 VDD.n587 GND 0.003347f
C2904 VDD.n588 GND 0.005387f
C2905 VDD.n589 GND 0.003347f
C2906 VDD.n590 GND 0.003347f
C2907 VDD.n591 GND 0.006693f
C2908 VDD.n592 GND 0.005387f
C2909 VDD.n593 GND 0.006693f
C2910 VDD.n594 GND 0.006693f
C2911 VDD.n595 GND 0.005387f
C2912 VDD.n596 GND 0.003347f
C2913 VDD.n597 GND 0.003347f
C2914 VDD.n598 GND 0.003347f
C2915 VDD.n599 GND 0.005387f
C2916 VDD.n600 GND 0.006693f
C2917 VDD.n601 GND 0.006693f
C2918 VDD.n602 GND 0.005387f
C2919 VDD.n603 GND 0.006693f
C2920 VDD.n604 GND 0.006693f
C2921 VDD.n605 GND 0.005387f
C2922 VDD.n606 GND 0.003347f
C2923 VDD.n607 GND 0.003347f
C2924 VDD.n608 GND 0.003347f
C2925 VDD.n609 GND 0.002721f
C2926 VDD.n610 GND 0.006693f
C2927 VDD.n611 GND 0.006693f
C2928 VDD.n612 GND 0.003582f
C2929 VDD.n613 GND 0.006693f
C2930 VDD.n614 GND 0.006693f
C2931 VDD.n615 GND 0.005387f
C2932 VDD.n616 GND 0.003347f
C2933 VDD.n617 GND 0.003347f
C2934 VDD.n618 GND 0.003347f
C2935 VDD.n619 GND 0.005387f
C2936 VDD.n620 GND 0.006693f
C2937 VDD.n621 GND 0.006693f
C2938 VDD.n622 GND 0.005387f
C2939 VDD.n623 GND 0.006693f
C2940 VDD.n624 GND 0.006693f
C2941 VDD.n625 GND 0.005387f
C2942 VDD.n626 GND 0.003347f
C2943 VDD.n627 GND 0.003347f
C2944 VDD.n628 GND 0.00251f
C2945 VDD.n629 GND 0.005387f
C2946 VDD.n630 GND 0.006693f
C2947 VDD.n631 GND 0.006693f
C2948 VDD.n632 GND 0.005387f
C2949 VDD.n633 GND 0.006693f
C2950 VDD.n634 GND 0.006693f
C2951 VDD.n635 GND 0.005387f
C2952 VDD.n636 GND 0.003347f
C2953 VDD.n637 GND 0.003347f
C2954 VDD.n638 GND 0.003347f
C2955 VDD.n639 GND 0.005387f
C2956 VDD.n640 GND 0.006693f
C2957 VDD.n641 GND 0.006693f
C2958 VDD.n642 GND 0.002721f
C2959 VDD.n643 GND 0.007407f
C2960 VDD.n644 GND 0.006693f
C2961 VDD.n645 GND 0.006693f
C2962 VDD.n646 GND 0.003582f
C2963 VDD.n647 GND 0.003347f
C2964 VDD.n648 GND 0.003347f
C2965 VDD.n649 GND 0.003347f
C2966 VDD.n650 GND 0.005387f
C2967 VDD.n651 GND 0.006693f
C2968 VDD.n652 GND 0.006693f
C2969 VDD.n653 GND 0.005387f
C2970 VDD.n654 GND 0.006693f
C2971 VDD.n655 GND 0.006693f
C2972 VDD.n656 GND 0.005387f
C2973 VDD.n657 GND 0.003347f
C2974 VDD.n658 GND 0.003347f
C2975 VDD.n659 GND 0.003347f
C2976 VDD.n660 GND 0.005387f
C2977 VDD.n661 GND 0.006693f
C2978 VDD.n662 GND 0.006693f
C2979 VDD.n663 GND 0.005387f
C2980 VDD.n664 GND 0.006693f
C2981 VDD.n665 GND 0.006693f
C2982 VDD.n666 GND 0.005387f
C2983 VDD.n667 GND 0.003347f
C2984 VDD.n668 GND 0.003347f
C2985 VDD.n669 GND 0.003347f
C2986 VDD.n670 GND 0.005387f
C2987 VDD.n671 GND 0.006693f
C2988 VDD.n672 GND 0.006693f
C2989 VDD.n673 GND 0.005387f
C2990 VDD.n674 GND 0.002721f
C2991 VDD.n675 GND 0.002108f
C2992 VDD.n676 GND 0.004551f
C2993 VDD.n677 GND 0.004551f
C2994 VDD.t162 GND 7.0265f
C2995 VDD.t87 GND 6.34775f
C2996 VDD.t0 GND 4.6915f
C2997 VDD.n679 GND 1.82593f
C2998 VDD.n680 GND 0.004551f
C2999 VDD.n681 GND 0.004551f
C3000 VDD.n683 GND 0.004551f
C3001 VDD.t48 GND 0.154197f
C3002 VDD.t47 GND 0.733149f
C3003 VDD.n684 GND 0.09739f
C3004 VDD.t49 GND 0.103896f
C3005 VDD.n685 GND 0.100617f
C3006 VDD.n686 GND 0.004551f
C3007 VDD.n688 GND 0.010814f
C3008 VDD.n689 GND 0.004551f
C3009 VDD.n690 GND 0.004551f
C3010 VDD.n691 GND 0.325035f
C3011 VDD.n692 GND 0.004551f
C3012 VDD.n693 GND 0.470823f
C3013 VDD.n694 GND 0.004551f
C3014 VDD.n695 GND 0.004551f
C3015 VDD.n696 GND 0.010814f
C3016 VDD.n697 GND 0.004551f
C3017 VDD.n698 GND 0.004551f
C3018 VDD.n699 GND 0.004551f
C3019 VDD.n700 GND 0.004551f
C3020 VDD.n702 GND 0.004551f
C3021 VDD.n703 GND 0.004551f
C3022 VDD.n705 GND 0.004551f
C3023 VDD.n706 GND 0.004551f
C3024 VDD.n708 GND 0.004551f
C3025 VDD.t41 GND 0.154197f
C3026 VDD.t39 GND 0.733149f
C3027 VDD.n709 GND 0.09739f
C3028 VDD.t42 GND 0.103896f
C3029 VDD.n710 GND 0.100617f
C3030 VDD.n711 GND 0.005616f
C3031 VDD.n713 GND 0.00261f
C3032 VDD.n714 GND 0.004551f
C3033 VDD.n715 GND 0.004551f
C3034 VDD.n716 GND 0.004551f
C3035 VDD.n717 GND 0.325035f
C3036 VDD.n718 GND 0.004551f
C3037 VDD.n719 GND 0.004551f
C3038 VDD.n720 GND 0.004551f
C3039 VDD.n721 GND 0.004551f
C3040 VDD.n722 GND 0.004551f
C3041 VDD.n723 GND 0.325035f
C3042 VDD.n724 GND 0.004551f
C3043 VDD.n725 GND 0.004551f
C3044 VDD.n726 GND 0.004551f
C3045 VDD.n727 GND 0.004551f
C3046 VDD.n728 GND 0.004551f
C3047 VDD.n729 GND 0.004551f
C3048 VDD.n730 GND 0.210317f
C3049 VDD.n731 GND 0.004551f
C3050 VDD.n732 GND 0.004551f
C3051 VDD.n733 GND 0.004551f
C3052 VDD.n734 GND 0.004551f
C3053 VDD.n735 GND 0.004551f
C3054 VDD.n736 GND 0.325035f
C3055 VDD.n737 GND 0.004551f
C3056 VDD.n738 GND 0.004551f
C3057 VDD.t158 GND 0.162518f
C3058 VDD.n739 GND 0.004551f
C3059 VDD.n740 GND 0.004551f
C3060 VDD.n741 GND 0.004551f
C3061 VDD.t40 GND 0.162518f
C3062 VDD.n742 GND 0.004551f
C3063 VDD.n743 GND 0.004551f
C3064 VDD.n744 GND 0.004551f
C3065 VDD.n745 GND 0.004551f
C3066 VDD.n746 GND 0.004551f
C3067 VDD.n747 GND 0.325035f
C3068 VDD.n748 GND 0.004551f
C3069 VDD.n749 GND 0.004551f
C3070 VDD.n750 GND 0.282016f
C3071 VDD.n751 GND 0.004551f
C3072 VDD.n752 GND 0.004551f
C3073 VDD.n753 GND 0.004551f
C3074 VDD.n754 GND 0.325035f
C3075 VDD.n755 GND 0.004551f
C3076 VDD.n756 GND 0.004551f
C3077 VDD.n757 GND 0.004551f
C3078 VDD.n758 GND 0.004551f
C3079 VDD.n759 GND 0.004551f
C3080 VDD.n760 GND 0.325035f
C3081 VDD.n761 GND 0.004551f
C3082 VDD.n762 GND 0.004551f
C3083 VDD.n763 GND 0.004551f
C3084 VDD.n764 GND 0.004551f
C3085 VDD.n765 GND 0.004551f
C3086 VDD.n766 GND 0.325035f
C3087 VDD.n767 GND 0.004551f
C3088 VDD.n768 GND 0.004551f
C3089 VDD.n769 GND 0.004551f
C3090 VDD.n770 GND 0.004551f
C3091 VDD.n771 GND 0.004551f
C3092 VDD.n772 GND 0.325035f
C3093 VDD.n773 GND 0.004551f
C3094 VDD.n774 GND 0.004551f
C3095 VDD.n775 GND 0.004551f
C3096 VDD.n776 GND 0.004551f
C3097 VDD.n777 GND 0.004551f
C3098 VDD.n778 GND 0.325035f
C3099 VDD.n779 GND 0.004551f
C3100 VDD.n780 GND 0.004551f
C3101 VDD.n781 GND 0.004551f
C3102 VDD.n782 GND 0.004551f
C3103 VDD.n783 GND 0.004551f
C3104 VDD.n784 GND 0.325035f
C3105 VDD.n785 GND 0.004551f
C3106 VDD.n786 GND 0.004551f
C3107 VDD.n787 GND 0.004551f
C3108 VDD.n788 GND 0.004551f
C3109 VDD.n789 GND 0.004551f
C3110 VDD.n790 GND 0.325035f
C3111 VDD.n791 GND 0.004551f
C3112 VDD.n792 GND 0.004551f
C3113 VDD.n793 GND 0.004551f
C3114 VDD.n794 GND 0.004551f
C3115 VDD.n795 GND 0.004551f
C3116 VDD.n796 GND 0.325035f
C3117 VDD.n797 GND 0.004551f
C3118 VDD.n798 GND 0.004551f
C3119 VDD.n799 GND 0.004551f
C3120 VDD.n800 GND 0.004551f
C3121 VDD.n801 GND 0.004551f
C3122 VDD.n802 GND 0.325035f
C3123 VDD.n803 GND 0.004551f
C3124 VDD.n804 GND 0.004551f
C3125 VDD.n805 GND 0.004551f
C3126 VDD.n806 GND 0.004551f
C3127 VDD.n807 GND 0.004551f
C3128 VDD.n808 GND 0.320255f
C3129 VDD.n809 GND 0.004551f
C3130 VDD.n810 GND 0.004551f
C3131 VDD.n811 GND 0.004551f
C3132 VDD.n812 GND 0.004551f
C3133 VDD.n813 GND 0.004551f
C3134 VDD.n814 GND 0.325035f
C3135 VDD.n815 GND 0.004551f
C3136 VDD.n816 GND 0.004551f
C3137 VDD.t81 GND 0.162518f
C3138 VDD.n817 GND 0.004551f
C3139 VDD.n818 GND 0.004551f
C3140 VDD.n819 GND 0.004551f
C3141 VDD.t92 GND 0.162518f
C3142 VDD.n820 GND 0.004551f
C3143 VDD.n821 GND 0.004551f
C3144 VDD.n822 GND 0.004551f
C3145 VDD.n823 GND 0.004551f
C3146 VDD.n824 GND 0.004551f
C3147 VDD.n825 GND 0.325035f
C3148 VDD.n826 GND 0.004551f
C3149 VDD.n827 GND 0.004551f
C3150 VDD.n828 GND 0.286796f
C3151 VDD.n829 GND 0.004551f
C3152 VDD.n830 GND 0.004551f
C3153 VDD.n831 GND 0.004551f
C3154 VDD.n832 GND 0.325035f
C3155 VDD.n833 GND 0.004551f
C3156 VDD.n834 GND 0.004551f
C3157 VDD.n835 GND 0.004551f
C3158 VDD.n836 GND 0.004551f
C3159 VDD.n837 GND 0.004551f
C3160 VDD.n838 GND 0.325035f
C3161 VDD.n839 GND 0.004551f
C3162 VDD.n840 GND 0.004551f
C3163 VDD.n841 GND 0.004551f
C3164 VDD.n842 GND 0.004551f
C3165 VDD.n843 GND 0.004551f
C3166 VDD.n844 GND 0.325035f
C3167 VDD.n845 GND 0.004551f
C3168 VDD.n846 GND 0.004551f
C3169 VDD.n847 GND 0.004551f
C3170 VDD.n848 GND 0.004551f
C3171 VDD.n849 GND 0.004551f
C3172 VDD.n850 GND 0.325035f
C3173 VDD.n851 GND 0.004551f
C3174 VDD.n852 GND 0.004551f
C3175 VDD.n853 GND 0.004551f
C3176 VDD.n854 GND 0.004551f
C3177 VDD.n855 GND 0.004551f
C3178 VDD.n856 GND 0.325035f
C3179 VDD.n857 GND 0.004551f
C3180 VDD.n858 GND 0.004551f
C3181 VDD.n859 GND 0.004551f
C3182 VDD.n860 GND 0.004551f
C3183 VDD.n861 GND 0.004551f
C3184 VDD.n862 GND 0.325035f
C3185 VDD.n863 GND 0.004551f
C3186 VDD.n864 GND 0.004551f
C3187 VDD.n865 GND 0.004551f
C3188 VDD.n866 GND 0.004551f
C3189 VDD.n867 GND 0.004551f
C3190 VDD.n868 GND 0.243776f
C3191 VDD.n869 GND 0.004551f
C3192 VDD.n870 GND 0.004551f
C3193 VDD.n871 GND 0.004551f
C3194 VDD.n872 GND 0.004551f
C3195 VDD.n873 GND 0.004551f
C3196 VDD.n874 GND 0.286796f
C3197 VDD.n875 GND 0.004551f
C3198 VDD.n876 GND 0.004551f
C3199 VDD.t72 GND 0.162518f
C3200 VDD.n877 GND 0.004551f
C3201 VDD.n878 GND 0.004551f
C3202 VDD.n879 GND 0.004551f
C3203 VDD.n880 GND 0.325035f
C3204 VDD.n881 GND 0.004551f
C3205 VDD.n882 GND 0.004551f
C3206 VDD.t82 GND 0.162518f
C3207 VDD.n883 GND 0.004551f
C3208 VDD.n884 GND 0.004551f
C3209 VDD.n885 GND 0.004551f
C3210 VDD.n886 GND 0.325035f
C3211 VDD.n887 GND 0.004551f
C3212 VDD.n888 GND 0.004551f
C3213 VDD.n889 GND 0.004551f
C3214 VDD.n890 GND 0.004551f
C3215 VDD.n891 GND 0.004551f
C3216 VDD.n892 GND 0.325035f
C3217 VDD.n893 GND 0.004551f
C3218 VDD.n894 GND 0.004551f
C3219 VDD.n895 GND 0.004551f
C3220 VDD.n896 GND 0.004551f
C3221 VDD.n897 GND 0.004551f
C3222 VDD.n898 GND 0.325035f
C3223 VDD.n899 GND 0.004551f
C3224 VDD.n900 GND 0.004551f
C3225 VDD.n901 GND 0.004551f
C3226 VDD.n902 GND 0.004551f
C3227 VDD.n903 GND 0.004551f
C3228 VDD.n904 GND 0.325035f
C3229 VDD.n905 GND 0.004551f
C3230 VDD.n906 GND 0.004551f
C3231 VDD.n907 GND 0.004551f
C3232 VDD.n908 GND 0.004551f
C3233 VDD.n909 GND 0.004551f
C3234 VDD.n910 GND 0.325035f
C3235 VDD.n911 GND 0.004551f
C3236 VDD.n912 GND 0.004551f
C3237 VDD.n913 GND 0.004551f
C3238 VDD.n914 GND 0.004551f
C3239 VDD.n915 GND 0.004551f
C3240 VDD.n916 GND 0.325035f
C3241 VDD.n917 GND 0.004551f
C3242 VDD.n918 GND 0.004551f
C3243 VDD.n919 GND 0.004551f
C3244 VDD.n920 GND 0.004551f
C3245 VDD.n921 GND 0.004551f
C3246 VDD.n922 GND 0.325035f
C3247 VDD.n923 GND 0.004551f
C3248 VDD.n924 GND 0.004551f
C3249 VDD.n925 GND 0.004551f
C3250 VDD.n926 GND 0.004551f
C3251 VDD.n927 GND 0.004551f
C3252 VDD.n928 GND 0.167298f
C3253 VDD.n929 GND 0.004551f
C3254 VDD.n930 GND 0.004551f
C3255 VDD.n931 GND 0.004551f
C3256 VDD.n932 GND 0.004551f
C3257 VDD.n933 GND 0.004551f
C3258 VDD.n934 GND 0.210317f
C3259 VDD.n935 GND 0.004551f
C3260 VDD.n936 GND 0.004551f
C3261 VDD.t91 GND 0.162518f
C3262 VDD.n937 GND 0.004551f
C3263 VDD.n938 GND 0.004551f
C3264 VDD.n939 GND 0.004551f
C3265 VDD.n940 GND 0.325035f
C3266 VDD.n941 GND 0.004551f
C3267 VDD.n942 GND 0.004551f
C3268 VDD.t98 GND 0.162518f
C3269 VDD.n943 GND 0.004551f
C3270 VDD.n944 GND 0.004551f
C3271 VDD.n945 GND 0.004551f
C3272 VDD.n946 GND 0.325035f
C3273 VDD.n947 GND 0.004551f
C3274 VDD.n948 GND 0.004551f
C3275 VDD.n949 GND 0.004551f
C3276 VDD.n950 GND 0.004551f
C3277 VDD.n951 GND 0.004551f
C3278 VDD.n952 GND 0.325035f
C3279 VDD.n953 GND 0.004551f
C3280 VDD.n954 GND 0.004551f
C3281 VDD.n955 GND 0.004551f
C3282 VDD.n956 GND 0.004551f
C3283 VDD.n957 GND 0.004551f
C3284 VDD.n958 GND 0.325035f
C3285 VDD.n959 GND 0.004551f
C3286 VDD.n960 GND 0.004551f
C3287 VDD.n961 GND 0.004551f
C3288 VDD.n962 GND 0.004551f
C3289 VDD.n963 GND 0.004551f
C3290 VDD.n964 GND 0.325035f
C3291 VDD.n965 GND 0.004551f
C3292 VDD.n966 GND 0.004551f
C3293 VDD.n967 GND 0.004551f
C3294 VDD.n968 GND 0.004551f
C3295 VDD.n969 GND 0.004551f
C3296 VDD.n970 GND 0.325035f
C3297 VDD.n971 GND 0.004551f
C3298 VDD.n972 GND 0.004551f
C3299 VDD.n973 GND 0.004551f
C3300 VDD.n974 GND 0.004551f
C3301 VDD.n975 GND 0.004551f
C3302 VDD.n976 GND 0.325035f
C3303 VDD.n977 GND 0.004551f
C3304 VDD.n978 GND 0.004551f
C3305 VDD.n979 GND 0.004551f
C3306 VDD.n980 GND 0.004551f
C3307 VDD.n981 GND 0.004551f
C3308 VDD.n982 GND 0.325035f
C3309 VDD.n983 GND 0.004551f
C3310 VDD.n984 GND 0.004551f
C3311 VDD.n985 GND 0.004551f
C3312 VDD.n986 GND 0.004551f
C3313 VDD.n987 GND 0.004551f
C3314 VDD.n988 GND 0.325035f
C3315 VDD.n989 GND 0.004551f
C3316 VDD.n990 GND 0.004551f
C3317 VDD.n991 GND 0.004551f
C3318 VDD.n992 GND 0.004551f
C3319 VDD.n993 GND 0.004551f
C3320 VDD.t76 GND 0.162518f
C3321 VDD.n994 GND 0.004551f
C3322 VDD.n995 GND 0.004551f
C3323 VDD.n996 GND 0.004551f
C3324 VDD.n997 GND 0.004551f
C3325 VDD.n998 GND 0.004551f
C3326 VDD.t63 GND 0.162518f
C3327 VDD.n999 GND 0.004551f
C3328 VDD.n1000 GND 0.004551f
C3329 VDD.n1001 GND 0.191197f
C3330 VDD.n1002 GND 0.004551f
C3331 VDD.n1003 GND 0.004551f
C3332 VDD.n1004 GND 0.004551f
C3333 VDD.n1005 GND 0.325035f
C3334 VDD.n1006 GND 0.004551f
C3335 VDD.n1007 GND 0.004551f
C3336 VDD.n1008 GND 0.205537f
C3337 VDD.n1009 GND 0.004551f
C3338 VDD.n1010 GND 0.004551f
C3339 VDD.n1011 GND 0.004551f
C3340 VDD.n1012 GND 0.325035f
C3341 VDD.n1013 GND 0.004551f
C3342 VDD.n1014 GND 0.004551f
C3343 VDD.n1015 GND 0.004551f
C3344 VDD.n1016 GND 0.004551f
C3345 VDD.n1017 GND 0.004551f
C3346 VDD.n1018 GND 0.325035f
C3347 VDD.n1019 GND 0.004551f
C3348 VDD.n1020 GND 0.004551f
C3349 VDD.n1021 GND 0.004551f
C3350 VDD.n1022 GND 0.004551f
C3351 VDD.n1023 GND 0.004551f
C3352 VDD.n1024 GND 0.325035f
C3353 VDD.n1025 GND 0.004551f
C3354 VDD.n1026 GND 0.004551f
C3355 VDD.n1027 GND 0.004551f
C3356 VDD.n1028 GND 0.004551f
C3357 VDD.n1029 GND 0.004551f
C3358 VDD.n1030 GND 0.325035f
C3359 VDD.n1031 GND 0.004551f
C3360 VDD.n1032 GND 0.004551f
C3361 VDD.n1033 GND 0.004551f
C3362 VDD.n1034 GND 0.011274f
C3363 VDD.n1035 GND 0.011274f
C3364 VDD.n1036 GND 0.470823f
C3365 VDD.n1037 GND 0.011274f
C3366 VDD.n1058 GND 0.010814f
C3367 VDD.n1059 GND 0.004551f
C3368 VDD.n1060 GND 0.010814f
C3369 VDD.t45 GND 0.154197f
C3370 VDD.t43 GND 0.733149f
C3371 VDD.n1061 GND 0.09739f
C3372 VDD.t46 GND 0.103896f
C3373 VDD.n1062 GND 0.100617f
C3374 VDD.n1063 GND 0.005616f
C3375 VDD.n1064 GND 0.011323f
C3376 VDD.n1065 GND 0.004551f
C3377 VDD.n1066 GND 0.004551f
C3378 VDD.n1067 GND 0.325035f
C3379 VDD.n1068 GND 0.004551f
C3380 VDD.n1069 GND 0.004551f
C3381 VDD.n1070 GND 0.004551f
C3382 VDD.n1071 GND 0.004551f
C3383 VDD.n1072 GND 0.004551f
C3384 VDD.n1073 GND 0.325035f
C3385 VDD.n1074 GND 0.004551f
C3386 VDD.n1075 GND 0.004551f
C3387 VDD.n1076 GND 0.004551f
C3388 VDD.n1077 GND 0.004551f
C3389 VDD.n1078 GND 0.004551f
C3390 VDD.t70 GND 0.154197f
C3391 VDD.t69 GND 0.733149f
C3392 VDD.n1079 GND 0.09739f
C3393 VDD.t71 GND 0.103896f
C3394 VDD.n1080 GND 0.100617f
C3395 VDD.n1081 GND 0.005616f
C3396 VDD.n1082 GND 0.004551f
C3397 VDD.n1083 GND 0.004551f
C3398 VDD.n1084 GND 0.325035f
C3399 VDD.n1085 GND 0.004551f
C3400 VDD.n1086 GND 0.004551f
C3401 VDD.n1087 GND 0.004551f
C3402 VDD.n1088 GND 0.004551f
C3403 VDD.n1089 GND 0.004551f
C3404 VDD.n1090 GND 0.325035f
C3405 VDD.n1091 GND 0.004551f
C3406 VDD.n1092 GND 0.004551f
C3407 VDD.n1093 GND 0.004551f
C3408 VDD.n1094 GND 0.004551f
C3409 VDD.n1095 GND 0.004551f
C3410 VDD.n1096 GND 0.004551f
C3411 VDD.n1097 GND 0.325035f
C3412 VDD.n1098 GND 0.004551f
C3413 VDD.n1099 GND 0.004551f
C3414 VDD.n1100 GND 0.004551f
C3415 VDD.n1101 GND 0.004551f
C3416 VDD.n1102 GND 0.004551f
C3417 VDD.t44 GND 0.162518f
C3418 VDD.n1103 GND 0.004551f
C3419 VDD.n1104 GND 0.004551f
C3420 VDD.n1105 GND 0.004551f
C3421 VDD.n1106 GND 0.004551f
C3422 VDD.n1107 GND 0.004551f
C3423 VDD.t85 GND 0.162518f
C3424 VDD.n1108 GND 0.004551f
C3425 VDD.n1109 GND 0.004551f
C3426 VDD.n1110 GND 0.282016f
C3427 VDD.n1111 GND 0.004551f
C3428 VDD.n1112 GND 0.004551f
C3429 VDD.n1113 GND 0.004551f
C3430 VDD.n1114 GND 0.325035f
C3431 VDD.n1115 GND 0.004551f
C3432 VDD.n1116 GND 0.004551f
C3433 VDD.n1117 GND 0.296356f
C3434 VDD.n1118 GND 0.004551f
C3435 VDD.n1119 GND 0.004551f
C3436 VDD.n1120 GND 0.004551f
C3437 VDD.n1121 GND 0.325035f
C3438 VDD.n1122 GND 0.004551f
C3439 VDD.n1123 GND 0.004551f
C3440 VDD.n1124 GND 0.004551f
C3441 VDD.n1125 GND 0.004551f
C3442 VDD.n1126 GND 0.004551f
C3443 VDD.n1127 GND 0.325035f
C3444 VDD.n1128 GND 0.004551f
C3445 VDD.n1129 GND 0.004551f
C3446 VDD.n1130 GND 0.004551f
C3447 VDD.n1131 GND 0.004551f
C3448 VDD.n1132 GND 0.004551f
C3449 VDD.n1133 GND 0.325035f
C3450 VDD.n1134 GND 0.004551f
C3451 VDD.n1135 GND 0.004551f
C3452 VDD.n1136 GND 0.004551f
C3453 VDD.n1137 GND 0.004551f
C3454 VDD.n1138 GND 0.004551f
C3455 VDD.n1139 GND 0.325035f
C3456 VDD.n1140 GND 0.004551f
C3457 VDD.n1141 GND 0.004551f
C3458 VDD.n1142 GND 0.004551f
C3459 VDD.n1143 GND 0.004551f
C3460 VDD.n1144 GND 0.004551f
C3461 VDD.n1145 GND 0.325035f
C3462 VDD.n1146 GND 0.004551f
C3463 VDD.n1147 GND 0.004551f
C3464 VDD.n1148 GND 0.004551f
C3465 VDD.n1149 GND 0.004551f
C3466 VDD.n1150 GND 0.004551f
C3467 VDD.n1151 GND 0.325035f
C3468 VDD.n1152 GND 0.004551f
C3469 VDD.n1153 GND 0.004551f
C3470 VDD.n1154 GND 0.004551f
C3471 VDD.n1155 GND 0.004551f
C3472 VDD.n1156 GND 0.004551f
C3473 VDD.n1157 GND 0.325035f
C3474 VDD.n1158 GND 0.004551f
C3475 VDD.n1159 GND 0.004551f
C3476 VDD.n1160 GND 0.004551f
C3477 VDD.n1161 GND 0.004551f
C3478 VDD.n1162 GND 0.004551f
C3479 VDD.n1163 GND 0.277236f
C3480 VDD.n1164 GND 0.004551f
C3481 VDD.n1165 GND 0.004551f
C3482 VDD.n1166 GND 0.004551f
C3483 VDD.n1167 GND 0.004551f
C3484 VDD.n1168 GND 0.004551f
C3485 VDD.n1169 GND 0.320255f
C3486 VDD.n1170 GND 0.004551f
C3487 VDD.n1171 GND 0.004551f
C3488 VDD.t100 GND 0.162518f
C3489 VDD.n1172 GND 0.004551f
C3490 VDD.n1173 GND 0.004551f
C3491 VDD.n1174 GND 0.004551f
C3492 VDD.n1175 GND 0.325035f
C3493 VDD.n1176 GND 0.004551f
C3494 VDD.n1177 GND 0.004551f
C3495 VDD.t3 GND 0.162518f
C3496 VDD.n1178 GND 0.004551f
C3497 VDD.n1179 GND 0.004551f
C3498 VDD.n1180 GND 0.004551f
C3499 VDD.n1181 GND 0.325035f
C3500 VDD.n1182 GND 0.004551f
C3501 VDD.n1183 GND 0.004551f
C3502 VDD.n1184 GND 0.004551f
C3503 VDD.n1185 GND 0.004551f
C3504 VDD.n1186 GND 0.004551f
C3505 VDD.n1187 GND 0.325035f
C3506 VDD.n1188 GND 0.004551f
C3507 VDD.n1189 GND 0.004551f
C3508 VDD.n1190 GND 0.004551f
C3509 VDD.n1191 GND 0.004551f
C3510 VDD.n1192 GND 0.004551f
C3511 VDD.n1193 GND 0.325035f
C3512 VDD.n1194 GND 0.004551f
C3513 VDD.n1195 GND 0.004551f
C3514 VDD.n1196 GND 0.004551f
C3515 VDD.n1197 GND 0.004551f
C3516 VDD.n1198 GND 0.004551f
C3517 VDD.n1199 GND 0.325035f
C3518 VDD.n1200 GND 0.004551f
C3519 VDD.n1201 GND 0.004551f
C3520 VDD.n1202 GND 0.004551f
C3521 VDD.n1203 GND 0.004551f
C3522 VDD.n1204 GND 0.004551f
C3523 VDD.n1205 GND 0.325035f
C3524 VDD.n1206 GND 0.004551f
C3525 VDD.n1207 GND 0.004551f
C3526 VDD.n1208 GND 0.004551f
C3527 VDD.n1209 GND 0.004551f
C3528 VDD.n1210 GND 0.004551f
C3529 VDD.n1211 GND 0.325035f
C3530 VDD.n1212 GND 0.004551f
C3531 VDD.n1213 GND 0.004551f
C3532 VDD.n1214 GND 0.004551f
C3533 VDD.n1215 GND 0.004551f
C3534 VDD.n1216 GND 0.004551f
C3535 VDD.n1217 GND 0.325035f
C3536 VDD.n1218 GND 0.004551f
C3537 VDD.n1219 GND 0.004551f
C3538 VDD.n1220 GND 0.004551f
C3539 VDD.n1221 GND 0.004551f
C3540 VDD.n1222 GND 0.004551f
C3541 VDD.n1223 GND 0.200757f
C3542 VDD.n1224 GND 0.004551f
C3543 VDD.n1225 GND 0.004551f
C3544 VDD.n1226 GND 0.004551f
C3545 VDD.n1227 GND 0.004551f
C3546 VDD.n1228 GND 0.004551f
C3547 VDD.n1229 GND 0.243776f
C3548 VDD.n1230 GND 0.004551f
C3549 VDD.n1231 GND 0.004551f
C3550 VDD.t96 GND 0.162518f
C3551 VDD.n1232 GND 0.004551f
C3552 VDD.n1233 GND 0.004551f
C3553 VDD.n1234 GND 0.004551f
C3554 VDD.n1235 GND 0.325035f
C3555 VDD.n1236 GND 0.004551f
C3556 VDD.n1237 GND 0.004551f
C3557 VDD.t2 GND 0.162518f
C3558 VDD.n1238 GND 0.004551f
C3559 VDD.n1239 GND 0.004551f
C3560 VDD.n1240 GND 0.004551f
C3561 VDD.n1241 GND 0.325035f
C3562 VDD.n1242 GND 0.004551f
C3563 VDD.n1243 GND 0.004551f
C3564 VDD.n1244 GND 0.004551f
C3565 VDD.n1245 GND 0.004551f
C3566 VDD.n1246 GND 0.004551f
C3567 VDD.n1247 GND 0.325035f
C3568 VDD.n1248 GND 0.004551f
C3569 VDD.n1249 GND 0.004551f
C3570 VDD.n1250 GND 0.004551f
C3571 VDD.n1251 GND 0.004551f
C3572 VDD.n1252 GND 0.004551f
C3573 VDD.n1253 GND 0.325035f
C3574 VDD.n1254 GND 0.004551f
C3575 VDD.n1255 GND 0.004551f
C3576 VDD.n1256 GND 0.004551f
C3577 VDD.n1257 GND 0.004551f
C3578 VDD.n1258 GND 0.004551f
C3579 VDD.n1259 GND 0.325035f
C3580 VDD.n1260 GND 0.004551f
C3581 VDD.n1261 GND 0.004551f
C3582 VDD.n1262 GND 0.004551f
C3583 VDD.n1263 GND 0.004551f
C3584 VDD.n1264 GND 0.004551f
C3585 VDD.n1265 GND 0.325035f
C3586 VDD.n1266 GND 0.004551f
C3587 VDD.n1267 GND 0.004551f
C3588 VDD.n1268 GND 0.004551f
C3589 VDD.n1269 GND 0.004551f
C3590 VDD.n1270 GND 0.004551f
C3591 VDD.n1271 GND 0.325035f
C3592 VDD.n1272 GND 0.004551f
C3593 VDD.n1273 GND 0.004551f
C3594 VDD.n1274 GND 0.004551f
C3595 VDD.n1275 GND 0.004551f
C3596 VDD.n1276 GND 0.004551f
C3597 VDD.n1277 GND 0.325035f
C3598 VDD.n1278 GND 0.004551f
C3599 VDD.n1279 GND 0.004551f
C3600 VDD.n1280 GND 0.004551f
C3601 VDD.n1281 GND 0.004551f
C3602 VDD.n1282 GND 0.004551f
C3603 VDD.t94 GND 0.162518f
C3604 VDD.n1283 GND 0.004551f
C3605 VDD.n1284 GND 0.004551f
C3606 VDD.n1285 GND 0.004551f
C3607 VDD.n1286 GND 0.004551f
C3608 VDD.n1287 GND 0.004551f
C3609 VDD.n1288 GND 0.167298f
C3610 VDD.n1289 GND 0.004551f
C3611 VDD.n1290 GND 0.004551f
C3612 VDD.n1291 GND 0.200757f
C3613 VDD.n1292 GND 0.004551f
C3614 VDD.n1293 GND 0.004551f
C3615 VDD.n1294 GND 0.004551f
C3616 VDD.n1295 GND 0.325035f
C3617 VDD.n1296 GND 0.004551f
C3618 VDD.n1297 GND 0.004551f
C3619 VDD.t84 GND 0.162518f
C3620 VDD.n1298 GND 0.004551f
C3621 VDD.n1299 GND 0.004551f
C3622 VDD.n1300 GND 0.004551f
C3623 VDD.n1301 GND 0.325035f
C3624 VDD.n1302 GND 0.004551f
C3625 VDD.n1303 GND 0.004551f
C3626 VDD.n1304 GND 0.004551f
C3627 VDD.n1305 GND 0.004551f
C3628 VDD.n1306 GND 0.004551f
C3629 VDD.n1307 GND 0.325035f
C3630 VDD.n1308 GND 0.004551f
C3631 VDD.n1309 GND 0.004551f
C3632 VDD.n1310 GND 0.004551f
C3633 VDD.n1311 GND 0.004551f
C3634 VDD.n1312 GND 0.004551f
C3635 VDD.n1313 GND 0.325035f
C3636 VDD.n1314 GND 0.004551f
C3637 VDD.n1315 GND 0.004551f
C3638 VDD.n1316 GND 0.004551f
C3639 VDD.n1317 GND 0.004551f
C3640 VDD.n1318 GND 0.004551f
C3641 VDD.n1319 GND 0.325035f
C3642 VDD.n1320 GND 0.004551f
C3643 VDD.n1321 GND 0.004551f
C3644 VDD.n1322 GND 0.004551f
C3645 VDD.n1323 GND 0.004551f
C3646 VDD.n1324 GND 0.004551f
C3647 VDD.n1325 GND 0.325035f
C3648 VDD.n1326 GND 0.004551f
C3649 VDD.n1327 GND 0.004551f
C3650 VDD.n1328 GND 0.004551f
C3651 VDD.n1329 GND 0.004551f
C3652 VDD.n1330 GND 0.004551f
C3653 VDD.n1331 GND 0.325035f
C3654 VDD.n1332 GND 0.004551f
C3655 VDD.n1333 GND 0.004551f
C3656 VDD.n1334 GND 0.004551f
C3657 VDD.n1335 GND 0.004551f
C3658 VDD.n1336 GND 0.004551f
C3659 VDD.n1337 GND 0.325035f
C3660 VDD.n1338 GND 0.004551f
C3661 VDD.n1339 GND 0.004551f
C3662 VDD.n1340 GND 0.004551f
C3663 VDD.n1341 GND 0.004551f
C3664 VDD.n1342 GND 0.004551f
C3665 VDD.n1343 GND 0.325035f
C3666 VDD.n1344 GND 0.004551f
C3667 VDD.n1345 GND 0.004551f
C3668 VDD.n1346 GND 0.004551f
C3669 VDD.n1347 GND 0.004551f
C3670 VDD.n1348 GND 0.004551f
C3671 VDD.n1349 GND 0.325035f
C3672 VDD.n1350 GND 0.004551f
C3673 VDD.n1351 GND 0.004551f
C3674 VDD.n1352 GND 0.004551f
C3675 VDD.n1353 GND 0.004551f
C3676 VDD.n1354 GND 0.004551f
C3677 VDD.n1355 GND 0.325035f
C3678 VDD.n1356 GND 0.004551f
C3679 VDD.n1357 GND 0.004551f
C3680 VDD.n1358 GND 0.004551f
C3681 VDD.n1359 GND 0.004551f
C3682 VDD.n1360 GND 0.004551f
C3683 VDD.t5 GND 0.162518f
C3684 VDD.n1361 GND 0.004551f
C3685 VDD.n1362 GND 0.004551f
C3686 VDD.n1363 GND 0.004551f
C3687 VDD.n1364 GND 0.004551f
C3688 VDD.n1365 GND 0.004551f
C3689 VDD.n1366 GND 0.277236f
C3690 VDD.n1367 GND 0.004551f
C3691 VDD.n1368 GND 0.004551f
C3692 VDD.n1369 GND 0.205537f
C3693 VDD.n1370 GND 0.004551f
C3694 VDD.n1371 GND 0.004551f
C3695 VDD.n1372 GND 0.004551f
C3696 VDD.n1373 GND 0.325035f
C3697 VDD.n1374 GND 0.004551f
C3698 VDD.n1375 GND 0.004551f
C3699 VDD.t160 GND 0.162518f
C3700 VDD.n1376 GND 0.004551f
C3701 VDD.n1377 GND 0.004551f
C3702 VDD.n1378 GND 0.004551f
C3703 VDD.n1379 GND 0.325035f
C3704 VDD.n1380 GND 0.004551f
C3705 VDD.n1381 GND 0.004551f
C3706 VDD.n1382 GND 0.004551f
C3707 VDD.n1383 GND 0.004551f
C3708 VDD.n1384 GND 0.004551f
C3709 VDD.n1385 GND 0.325035f
C3710 VDD.n1386 GND 0.004551f
C3711 VDD.n1387 GND 0.004551f
C3712 VDD.n1388 GND 0.004551f
C3713 VDD.n1389 GND 0.004551f
C3714 VDD.n1390 GND 0.004551f
C3715 VDD.n1391 GND 0.325035f
C3716 VDD.n1392 GND 0.004551f
C3717 VDD.n1393 GND 0.004551f
C3718 VDD.n1394 GND 0.004551f
C3719 VDD.n1395 GND 0.011274f
C3720 VDD.n1396 GND 0.011274f
C3721 VDD.n1397 GND 1.82593f
C3722 VDD.n1398 GND 0.010814f
C3723 VDD.n1399 GND 0.010814f
C3724 VDD.n1400 GND 0.011274f
C3725 VDD.n1401 GND 0.004551f
C3726 VDD.n1403 GND 0.004551f
C3727 VDD.n1404 GND 0.004551f
C3728 VDD.n1405 GND 0.004551f
C3729 VDD.n1406 GND 0.004551f
C3730 VDD.n1407 GND 0.004551f
C3731 VDD.n1408 GND 0.004551f
C3732 VDD.t17 GND 0.154197f
C3733 VDD.t15 GND 0.733149f
C3734 VDD.n1409 GND 0.09739f
C3735 VDD.t16 GND 0.103896f
C3736 VDD.n1410 GND 0.100617f
C3737 VDD.n1411 GND 0.005616f
C3738 VDD.n1413 GND 0.004551f
C3739 VDD.n1414 GND 0.004551f
C3740 VDD.n1415 GND 0.004551f
C3741 VDD.n1416 GND 0.004551f
C3742 VDD.n1417 GND 0.004551f
C3743 VDD.n1418 GND 0.004551f
C3744 VDD.n1419 GND 0.004551f
C3745 VDD.n1420 GND 0.004551f
C3746 VDD.n1421 GND 0.004551f
C3747 VDD.n1422 GND 0.004551f
C3748 VDD.n1423 GND 0.004551f
C3749 VDD.n1424 GND 0.004551f
C3750 VDD.n1425 GND 0.004551f
C3751 VDD.n1426 GND 0.004551f
C3752 VDD.n1427 GND 0.004551f
C3753 VDD.n1428 GND 0.004551f
C3754 VDD.n1429 GND 0.004551f
C3755 VDD.n1430 GND 0.004551f
C3756 VDD.n1431 GND 0.004551f
C3757 VDD.n1432 GND 0.004551f
C3758 VDD.n1433 GND 0.004551f
C3759 VDD.n1434 GND 0.004551f
C3760 VDD.n1435 GND 0.004551f
C3761 VDD.n1436 GND 0.004551f
C3762 VDD.n1437 GND 0.004551f
C3763 VDD.n1438 GND 0.004551f
C3764 VDD.n1439 GND 0.004551f
C3765 VDD.n1440 GND 0.004551f
C3766 VDD.n1441 GND 0.004551f
C3767 VDD.n1442 GND 0.004551f
C3768 VDD.n1443 GND 0.004551f
C3769 VDD.n1444 GND 0.004551f
C3770 VDD.n1445 GND 0.004551f
C3771 VDD.n1446 GND 0.004551f
C3772 VDD.n1447 GND 0.004551f
C3773 VDD.n1448 GND 0.004551f
C3774 VDD.n1449 GND 0.004551f
C3775 VDD.n1450 GND 0.004551f
C3776 VDD.n1451 GND 0.004551f
C3777 VDD.n1452 GND 0.004551f
C3778 VDD.n1453 GND 0.004551f
C3779 VDD.n1454 GND 0.004551f
C3780 VDD.n1455 GND 0.004551f
C3781 VDD.n1456 GND 0.004551f
C3782 VDD.n1457 GND 0.004551f
C3783 VDD.n1458 GND 0.004551f
C3784 VDD.n1459 GND 0.004551f
C3785 VDD.n1460 GND 0.004551f
C3786 VDD.n1461 GND 0.004551f
C3787 VDD.n1462 GND 0.004551f
C3788 VDD.n1463 GND 0.004551f
C3789 VDD.n1464 GND 0.004551f
C3790 VDD.n1465 GND 0.004551f
C3791 VDD.n1466 GND 0.004551f
C3792 VDD.n1467 GND 0.004551f
C3793 VDD.n1468 GND 0.004551f
C3794 VDD.n1469 GND 0.004551f
C3795 VDD.n1470 GND 0.004551f
C3796 VDD.n1471 GND 0.004551f
C3797 VDD.n1472 GND 0.004551f
C3798 VDD.n1473 GND 0.004551f
C3799 VDD.n1474 GND 0.004551f
C3800 VDD.n1475 GND 0.004551f
C3801 VDD.n1476 GND 0.004551f
C3802 VDD.n1477 GND 0.004551f
C3803 VDD.n1478 GND 0.004551f
C3804 VDD.n1479 GND 0.004551f
C3805 VDD.n1480 GND 0.004551f
C3806 VDD.n1481 GND 0.004551f
C3807 VDD.n1482 GND 0.004551f
C3808 VDD.n1483 GND 0.004551f
C3809 VDD.n1484 GND 0.004551f
C3810 VDD.n1485 GND 0.004551f
C3811 VDD.n1486 GND 0.004551f
C3812 VDD.n1487 GND 0.004551f
C3813 VDD.n1488 GND 0.004551f
C3814 VDD.n1489 GND 0.004551f
C3815 VDD.n1490 GND 0.004551f
C3816 VDD.n1491 GND 0.004551f
C3817 VDD.n1492 GND 0.004551f
C3818 VDD.n1493 GND 0.004551f
C3819 VDD.n1494 GND 0.004551f
C3820 VDD.n1495 GND 0.004551f
C3821 VDD.n1496 GND 0.004551f
C3822 VDD.n1497 GND 0.004551f
C3823 VDD.n1498 GND 0.004551f
C3824 VDD.n1499 GND 0.004551f
C3825 VDD.n1500 GND 0.004551f
C3826 VDD.n1501 GND 0.004551f
C3827 VDD.n1502 GND 0.004551f
C3828 VDD.n1503 GND 0.004551f
C3829 VDD.n1504 GND 0.004551f
C3830 VDD.n1505 GND 0.004551f
C3831 VDD.n1506 GND 0.004551f
C3832 VDD.n1507 GND 0.004551f
C3833 VDD.n1508 GND 0.004551f
C3834 VDD.n1509 GND 0.004551f
C3835 VDD.n1510 GND 0.004551f
C3836 VDD.n1511 GND 0.004551f
C3837 VDD.n1512 GND 0.004551f
C3838 VDD.n1513 GND 0.004551f
C3839 VDD.n1514 GND 0.004551f
C3840 VDD.n1515 GND 0.004551f
C3841 VDD.n1516 GND 0.004551f
C3842 VDD.n1517 GND 0.004551f
C3843 VDD.n1518 GND 0.004551f
C3844 VDD.n1519 GND 0.004551f
C3845 VDD.n1520 GND 0.004551f
C3846 VDD.n1521 GND 0.004551f
C3847 VDD.n1522 GND 0.004551f
C3848 VDD.n1523 GND 0.004551f
C3849 VDD.n1524 GND 0.004551f
C3850 VDD.n1525 GND 0.004551f
C3851 VDD.n1526 GND 0.004551f
C3852 VDD.n1527 GND 0.004551f
C3853 VDD.n1528 GND 0.004551f
C3854 VDD.n1529 GND 0.004551f
C3855 VDD.n1530 GND 0.004551f
C3856 VDD.n1531 GND 0.004551f
C3857 VDD.n1532 GND 0.004551f
C3858 VDD.n1533 GND 0.004551f
C3859 VDD.n1534 GND 0.004551f
C3860 VDD.n1535 GND 0.004551f
C3861 VDD.n1536 GND 0.004551f
C3862 VDD.n1537 GND 0.004551f
C3863 VDD.n1538 GND 0.004551f
C3864 VDD.n1539 GND 0.004551f
C3865 VDD.n1540 GND 0.004551f
C3866 VDD.n1541 GND 0.004551f
C3867 VDD.n1542 GND 0.004551f
C3868 VDD.n1543 GND 0.004551f
C3869 VDD.n1544 GND 0.004551f
C3870 VDD.n1545 GND 0.004551f
C3871 VDD.n1546 GND 0.004551f
C3872 VDD.n1547 GND 0.004551f
C3873 VDD.n1548 GND 0.004551f
C3874 VDD.n1549 GND 0.004551f
C3875 VDD.n1550 GND 0.004551f
C3876 VDD.n1551 GND 0.004551f
C3877 VDD.n1552 GND 0.004551f
C3878 VDD.n1553 GND 0.004551f
C3879 VDD.n1554 GND 0.004551f
C3880 VDD.n1555 GND 0.004551f
C3881 VDD.n1556 GND 0.004551f
C3882 VDD.n1557 GND 0.004551f
C3883 VDD.n1558 GND 0.004551f
C3884 VDD.n1559 GND 0.004551f
C3885 VDD.n1560 GND 0.004551f
C3886 VDD.n1561 GND 0.004551f
C3887 VDD.n1562 GND 0.004551f
C3888 VDD.n1563 GND 0.004551f
C3889 VDD.n1564 GND 0.004551f
C3890 VDD.n1565 GND 0.004551f
C3891 VDD.n1566 GND 0.004551f
C3892 VDD.n1567 GND 0.004551f
C3893 VDD.n1568 GND 0.004551f
C3894 VDD.n1569 GND 0.004551f
C3895 VDD.n1570 GND 0.004551f
C3896 VDD.n1571 GND 0.004551f
C3897 VDD.n1572 GND 0.004551f
C3898 VDD.n1573 GND 0.004551f
C3899 VDD.n1574 GND 0.010814f
C3900 VDD.n1575 GND 0.011274f
C3901 VDD.n1576 GND 0.011274f
C3902 VDD.n1578 GND 0.004551f
C3903 VDD.n1579 GND 0.004551f
C3904 VDD.n1580 GND 0.004551f
C3905 VDD.n1581 GND 0.00261f
C3906 VDD.n1582 GND 0.004551f
C3907 VDD.n1584 GND 0.004551f
C3908 VDD.n1585 GND 0.004217f
C3909 VDD.n1586 GND 0.004551f
C3910 VDD.n1587 GND 0.004551f
C3911 VDD.n1588 GND 0.004551f
C3912 VDD.n1590 GND 0.004551f
C3913 VDD.n1592 GND 0.004551f
C3914 VDD.n1593 GND 0.004551f
C3915 VDD.n1594 GND 0.004551f
C3916 VDD.n1595 GND 0.009997f
C3917 VDD.n1596 GND 0.004551f
C3918 VDD.n1597 GND 0.004551f
C3919 VDD.n1598 GND 0.004551f
C3920 VDD.n1599 GND 0.004551f
C3921 VDD.n1600 GND 0.004551f
C3922 VDD.n1601 GND 0.004551f
C3923 VDD.n1603 GND 0.004551f
C3924 VDD.n1605 GND 0.004551f
C3925 VDD.n1606 GND 0.004551f
C3926 VDD.n1607 GND 0.004551f
C3927 VDD.n1608 GND 0.004551f
C3928 VDD.n1609 GND 0.004551f
C3929 VDD.n1611 GND 0.004551f
C3930 VDD.n1613 GND 0.004551f
C3931 VDD.n1614 GND 0.004551f
C3932 VDD.n1615 GND 0.004551f
C3933 VDD.n1616 GND 0.004551f
C3934 VDD.n1617 GND 0.004551f
C3935 VDD.n1619 GND 0.004551f
C3936 VDD.n1621 GND 0.004551f
C3937 VDD.n1622 GND 0.004551f
C3938 VDD.t7 GND 0.154197f
C3939 VDD.t4 GND 0.733149f
C3940 VDD.n1623 GND 0.09739f
C3941 VDD.t6 GND 0.103896f
C3942 VDD.n1624 GND 0.100617f
C3943 VDD.n1625 GND 0.004551f
C3944 VDD.n1626 GND 0.011274f
C3945 VDD.n1627 GND 0.004551f
C3946 VDD.n1628 GND 0.004551f
C3947 VDD.n1629 GND 0.004551f
C3948 VDD.n1630 GND 0.004551f
C3949 VDD.n1631 GND 0.004551f
C3950 VDD.n1632 GND 0.004551f
C3951 VDD.n1633 GND 0.004551f
C3952 VDD.n1634 GND 0.004551f
C3953 VDD.n1635 GND 0.004551f
C3954 VDD.n1636 GND 0.004551f
C3955 VDD.n1637 GND 0.004551f
C3956 VDD.n1638 GND 0.004551f
C3957 VDD.n1639 GND 0.004551f
C3958 VDD.n1640 GND 0.004551f
C3959 VDD.n1641 GND 0.004551f
C3960 VDD.n1642 GND 0.004551f
C3961 VDD.n1643 GND 0.004551f
C3962 VDD.n1644 GND 0.004551f
C3963 VDD.n1645 GND 0.004551f
C3964 VDD.n1646 GND 0.004551f
C3965 VDD.n1647 GND 0.004551f
C3966 VDD.n1648 GND 0.004551f
C3967 VDD.n1649 GND 0.004551f
C3968 VDD.n1650 GND 0.004551f
C3969 VDD.n1651 GND 0.004551f
C3970 VDD.n1652 GND 0.004551f
C3971 VDD.n1653 GND 0.004551f
C3972 VDD.n1654 GND 0.004551f
C3973 VDD.n1655 GND 0.004551f
C3974 VDD.n1656 GND 0.004551f
C3975 VDD.n1657 GND 0.004551f
C3976 VDD.n1658 GND 0.004551f
C3977 VDD.n1659 GND 0.004551f
C3978 VDD.n1660 GND 0.004551f
C3979 VDD.n1661 GND 0.004551f
C3980 VDD.n1662 GND 0.004551f
C3981 VDD.n1663 GND 0.004551f
C3982 VDD.n1664 GND 0.004551f
C3983 VDD.n1665 GND 0.004551f
C3984 VDD.n1666 GND 0.004551f
C3985 VDD.n1667 GND 0.004551f
C3986 VDD.n1668 GND 0.004551f
C3987 VDD.n1669 GND 0.004551f
C3988 VDD.n1670 GND 0.004551f
C3989 VDD.n1671 GND 0.004551f
C3990 VDD.n1672 GND 0.004551f
C3991 VDD.n1673 GND 0.004551f
C3992 VDD.n1674 GND 0.004551f
C3993 VDD.n1675 GND 0.004551f
C3994 VDD.n1676 GND 0.004551f
C3995 VDD.n1677 GND 0.004551f
C3996 VDD.n1678 GND 0.004551f
C3997 VDD.n1679 GND 0.004551f
C3998 VDD.n1680 GND 0.004551f
C3999 VDD.n1681 GND 0.004551f
C4000 VDD.n1682 GND 0.004551f
C4001 VDD.n1683 GND 0.004551f
C4002 VDD.n1684 GND 0.004551f
C4003 VDD.n1685 GND 0.004551f
C4004 VDD.n1686 GND 0.004551f
C4005 VDD.n1687 GND 0.004551f
C4006 VDD.n1688 GND 0.004551f
C4007 VDD.n1689 GND 0.004551f
C4008 VDD.n1690 GND 0.004551f
C4009 VDD.n1691 GND 0.004551f
C4010 VDD.n1692 GND 0.004551f
C4011 VDD.n1693 GND 0.004551f
C4012 VDD.n1694 GND 0.004551f
C4013 VDD.n1695 GND 0.004551f
C4014 VDD.n1696 GND 0.004551f
C4015 VDD.n1697 GND 0.004551f
C4016 VDD.n1698 GND 0.004551f
C4017 VDD.n1699 GND 0.004551f
C4018 VDD.n1700 GND 0.004551f
C4019 VDD.n1701 GND 0.004551f
C4020 VDD.n1702 GND 0.004551f
C4021 VDD.n1703 GND 0.004551f
C4022 VDD.n1704 GND 0.004551f
C4023 VDD.n1705 GND 0.004551f
C4024 VDD.n1706 GND 0.004551f
C4025 VDD.n1707 GND 0.004551f
C4026 VDD.n1708 GND 0.004551f
C4027 VDD.n1709 GND 0.004551f
C4028 VDD.n1710 GND 0.004551f
C4029 VDD.n1711 GND 0.004551f
C4030 VDD.n1712 GND 0.004551f
C4031 VDD.n1713 GND 0.004551f
C4032 VDD.n1714 GND 0.004551f
C4033 VDD.n1715 GND 0.004551f
C4034 VDD.n1716 GND 0.004551f
C4035 VDD.n1717 GND 0.004551f
C4036 VDD.n1718 GND 0.004551f
C4037 VDD.n1719 GND 0.004551f
C4038 VDD.n1720 GND 0.004551f
C4039 VDD.n1721 GND 0.004551f
C4040 VDD.n1722 GND 0.004551f
C4041 VDD.n1723 GND 0.004551f
C4042 VDD.n1724 GND 0.004551f
C4043 VDD.n1725 GND 0.004551f
C4044 VDD.n1726 GND 0.004551f
C4045 VDD.n1727 GND 0.004551f
C4046 VDD.n1728 GND 0.004551f
C4047 VDD.n1729 GND 0.004551f
C4048 VDD.n1730 GND 0.004551f
C4049 VDD.n1731 GND 0.004551f
C4050 VDD.n1732 GND 0.004551f
C4051 VDD.n1733 GND 0.004551f
C4052 VDD.n1734 GND 0.004551f
C4053 VDD.n1735 GND 0.004551f
C4054 VDD.n1736 GND 0.004551f
C4055 VDD.n1737 GND 0.004551f
C4056 VDD.n1738 GND 0.004551f
C4057 VDD.n1739 GND 0.004551f
C4058 VDD.n1740 GND 0.004551f
C4059 VDD.n1741 GND 0.004551f
C4060 VDD.n1742 GND 0.004551f
C4061 VDD.n1743 GND 0.004551f
C4062 VDD.n1744 GND 0.004551f
C4063 VDD.n1745 GND 0.004551f
C4064 VDD.n1746 GND 0.004551f
C4065 VDD.n1747 GND 0.004551f
C4066 VDD.n1748 GND 0.004551f
C4067 VDD.n1749 GND 0.004551f
C4068 VDD.n1750 GND 0.004551f
C4069 VDD.n1751 GND 0.004551f
C4070 VDD.n1752 GND 0.004551f
C4071 VDD.n1753 GND 0.004551f
C4072 VDD.n1754 GND 0.004551f
C4073 VDD.n1755 GND 0.004551f
C4074 VDD.n1756 GND 0.004551f
C4075 VDD.n1757 GND 0.004551f
C4076 VDD.n1758 GND 0.004551f
C4077 VDD.n1759 GND 0.004551f
C4078 VDD.n1760 GND 0.004551f
C4079 VDD.n1761 GND 0.004551f
C4080 VDD.n1762 GND 0.004551f
C4081 VDD.n1763 GND 0.004551f
C4082 VDD.n1764 GND 0.004551f
C4083 VDD.n1765 GND 0.004551f
C4084 VDD.n1766 GND 0.004551f
C4085 VDD.n1767 GND 0.004551f
C4086 VDD.n1768 GND 0.004551f
C4087 VDD.n1769 GND 0.004551f
C4088 VDD.n1770 GND 0.004551f
C4089 VDD.n1771 GND 0.004551f
C4090 VDD.n1772 GND 0.004551f
C4091 VDD.n1773 GND 0.004551f
C4092 VDD.n1774 GND 0.004551f
C4093 VDD.n1775 GND 0.004551f
C4094 VDD.n1776 GND 0.004551f
C4095 VDD.n1777 GND 0.004551f
C4096 VDD.n1778 GND 0.004551f
C4097 VDD.n1779 GND 0.004551f
C4098 VDD.n1780 GND 0.004551f
C4099 VDD.n1781 GND 0.010814f
C4100 VDD.n1782 GND 0.011274f
C4101 VDD.n1783 GND 0.004551f
C4102 VDD.n1784 GND 0.004551f
C4103 VDD.n1786 GND 0.004551f
C4104 VDD.n1788 GND 0.004551f
C4105 VDD.n1789 GND 0.00261f
C4106 VDD.n1790 GND 0.005616f
C4107 VDD.n1791 GND 0.004217f
C4108 VDD.n1792 GND 0.004551f
C4109 VDD.n1793 GND 0.004551f
C4110 VDD.n1795 GND 0.004551f
C4111 VDD.n1796 GND 0.004551f
C4112 VDD.n1797 GND 0.004551f
C4113 VDD.n1798 GND 0.004551f
C4114 VDD.n1799 GND 0.004551f
C4115 VDD.n1800 GND 0.004551f
C4116 VDD.n1802 GND 0.004551f
C4117 VDD.n1803 GND 0.189549f
C4118 VDD.n1804 GND 1.93121f
C4119 VDD.n1805 GND 0.00251f
C4120 VDD.n1806 GND 0.003347f
C4121 VDD.n1807 GND 0.005387f
C4122 VDD.n1808 GND 0.006693f
C4123 VDD.n1809 GND 0.006693f
C4124 VDD.n1810 GND 0.006693f
C4125 VDD.n1811 GND 0.005387f
C4126 VDD.n1812 GND 0.003347f
C4127 VDD.n1813 GND 0.006693f
C4128 VDD.t23 GND 0.118593f
C4129 VDD.t21 GND 0.540868f
C4130 VDD.n1814 GND 0.08957f
C4131 VDD.t24 GND 0.077791f
C4132 VDD.n1815 GND 0.092102f
C4133 VDD.n1816 GND 0.006693f
C4134 VDD.n1817 GND 0.006693f
C4135 VDD.n1818 GND 0.005387f
C4136 VDD.n1819 GND 0.003347f
C4137 VDD.n1820 GND 0.006693f
C4138 VDD.n1821 GND 0.006693f
C4139 VDD.n1822 GND 0.006693f
C4140 VDD.n1823 GND 0.005387f
C4141 VDD.n1824 GND 0.003347f
C4142 VDD.n1825 GND 0.006693f
C4143 VDD.n1826 GND 0.006693f
C4144 VDD.n1827 GND 0.006693f
C4145 VDD.n1828 GND 0.005387f
C4146 VDD.n1829 GND 0.003347f
C4147 VDD.n1830 GND 0.006693f
C4148 VDD.n1831 GND 0.006693f
C4149 VDD.t26 GND 0.118593f
C4150 VDD.t25 GND 0.540868f
C4151 VDD.n1832 GND 0.08957f
C4152 VDD.t27 GND 0.077791f
C4153 VDD.n1833 GND 0.092102f
C4154 VDD.n1834 GND 0.003782f
C4155 VDD.n1835 GND 0.01598f
C4156 VDD.n1836 GND 0.70265f
C4157 VDD.n1846 GND 0.005387f
C4158 VDD.n1847 GND 0.003347f
C4159 VDD.n1848 GND 0.005387f
C4160 VDD.n1849 GND 0.003347f
C4161 VDD.n1850 GND 0.005387f
C4162 VDD.n1851 GND 0.003347f
C4163 VDD.n1852 GND 0.005387f
C4164 VDD.n1853 GND 0.003347f
C4165 VDD.n1854 GND 0.006693f
C4166 VDD.n1855 GND 0.005387f
C4167 VDD.n1856 GND 0.006693f
C4168 VDD.n1857 GND 0.005387f
C4169 VDD.n1858 GND 0.006693f
C4170 VDD.n1859 GND 0.477993f
C4171 VDD.n1860 GND 0.006693f
C4172 VDD.n1861 GND 0.005387f
C4173 VDD.n1862 GND 0.004471f
C4174 VDD.n1863 GND 0.006693f
C4175 VDD.n1864 GND 0.005387f
C4176 VDD.n1865 GND 0.006693f
C4177 VDD.n1866 GND 0.477993f
C4178 VDD.n1867 GND 0.006693f
C4179 VDD.n1868 GND 0.005387f
C4180 VDD.n1869 GND 0.006693f
C4181 VDD.n1870 GND 0.005387f
C4182 VDD.n1871 GND 0.006693f
C4183 VDD.t22 GND 0.238997f
C4184 VDD.n1872 GND 0.006693f
C4185 VDD.n1873 GND 0.005387f
C4186 VDD.n1874 GND 0.005387f
C4187 VDD.n1875 GND 0.006693f
C4188 VDD.n1876 GND 0.005387f
C4189 VDD.n1877 GND 0.006693f
C4190 VDD.n1878 GND 0.477993f
C4191 VDD.n1879 GND 0.368055f
C4192 VDD.n1880 GND 0.006693f
C4193 VDD.n1881 GND 0.005387f
C4194 VDD.n1882 GND 0.006693f
C4195 VDD.n1883 GND 0.005387f
C4196 VDD.n1884 GND 0.006693f
C4197 VDD.n1885 GND 0.477993f
C4198 VDD.n1886 GND 0.006693f
C4199 VDD.n1887 GND 0.005387f
C4200 VDD.n1888 GND 0.006693f
C4201 VDD.n1889 GND 0.005387f
C4202 VDD.n1890 GND 0.006693f
C4203 VDD.n1891 GND 0.477993f
C4204 VDD.n1892 GND 0.006693f
C4205 VDD.n1893 GND 0.005387f
C4206 VDD.n1894 GND 0.006693f
C4207 VDD.n1895 GND 0.005387f
C4208 VDD.n1896 GND 0.006693f
C4209 VDD.n1897 GND 0.477993f
C4210 VDD.n1898 GND 0.006693f
C4211 VDD.n1899 GND 0.005387f
C4212 VDD.n1900 GND 0.006693f
C4213 VDD.n1901 GND 0.005387f
C4214 VDD.n1902 GND 0.006693f
C4215 VDD.n1903 GND 0.477993f
C4216 VDD.n1904 GND 0.006693f
C4217 VDD.n1905 GND 0.005387f
C4218 VDD.n1906 GND 0.006693f
C4219 VDD.n1907 GND 0.005387f
C4220 VDD.n1908 GND 0.006693f
C4221 VDD.n1909 GND 0.477993f
C4222 VDD.n1910 GND 0.006693f
C4223 VDD.n1911 GND 0.005387f
C4224 VDD.n1912 GND 0.006693f
C4225 VDD.n1913 GND 0.005387f
C4226 VDD.n1914 GND 0.006693f
C4227 VDD.n1915 GND 0.382394f
C4228 VDD.n1916 GND 0.006693f
C4229 VDD.n1917 GND 0.005387f
C4230 VDD.n1918 GND 0.006693f
C4231 VDD.n1919 GND 0.005387f
C4232 VDD.n1920 GND 0.006693f
C4233 VDD.n1921 GND 0.477993f
C4234 VDD.n1922 GND 0.006693f
C4235 VDD.n1923 GND 0.005387f
C4236 VDD.n1924 GND 0.006693f
C4237 VDD.n1925 GND 0.005387f
C4238 VDD.n1926 GND 0.006693f
C4239 VDD.n1927 GND 0.477993f
C4240 VDD.n1928 GND 0.006693f
C4241 VDD.n1929 GND 0.005387f
C4242 VDD.n1930 GND 0.006693f
C4243 VDD.n1931 GND 0.005387f
C4244 VDD.n1932 GND 0.006693f
C4245 VDD.n1933 GND 0.477993f
C4246 VDD.n1934 GND 0.006693f
C4247 VDD.n1935 GND 0.005387f
C4248 VDD.n1936 GND 0.006693f
C4249 VDD.n1937 GND 0.005387f
C4250 VDD.n1938 GND 0.006693f
C4251 VDD.n1939 GND 0.477993f
C4252 VDD.n1940 GND 0.006693f
C4253 VDD.n1941 GND 0.005387f
C4254 VDD.n1942 GND 0.006693f
C4255 VDD.n1943 GND 0.005387f
C4256 VDD.n1944 GND 0.006693f
C4257 VDD.n1945 GND 0.477993f
C4258 VDD.n1946 GND 0.006693f
C4259 VDD.n1947 GND 0.005387f
C4260 VDD.n1948 GND 0.006693f
C4261 VDD.n1949 GND 0.005387f
C4262 VDD.n1950 GND 0.006693f
C4263 VDD.n1951 GND 0.454093f
C4264 VDD.n1952 GND 0.006693f
C4265 VDD.n1953 GND 0.005387f
C4266 VDD.n1954 GND 0.006693f
C4267 VDD.n1955 GND 0.005387f
C4268 VDD.n1956 GND 0.006693f
C4269 VDD.n1957 GND 0.477993f
C4270 VDD.n1958 GND 0.006693f
C4271 VDD.n1959 GND 0.005387f
C4272 VDD.n1960 GND 0.006693f
C4273 VDD.n1961 GND 0.005387f
C4274 VDD.n1962 GND 0.006693f
C4275 VDD.n1963 GND 0.477993f
C4276 VDD.n1964 GND 0.006693f
C4277 VDD.n1965 GND 0.005387f
C4278 VDD.n1966 GND 0.006693f
C4279 VDD.n1967 GND 0.005387f
C4280 VDD.n1968 GND 0.006693f
C4281 VDD.n1969 GND 0.477993f
C4282 VDD.n1970 GND 0.006693f
C4283 VDD.n1971 GND 0.005387f
C4284 VDD.n1972 GND 0.006693f
C4285 VDD.n1973 GND 0.005387f
C4286 VDD.n1974 GND 0.006693f
C4287 VDD.n1975 GND 0.477993f
C4288 VDD.n1976 GND 0.006693f
C4289 VDD.n1977 GND 0.005387f
C4290 VDD.n1978 GND 0.006693f
C4291 VDD.n1979 GND 0.005387f
C4292 VDD.n1980 GND 0.006693f
C4293 VDD.n1981 GND 0.477993f
C4294 VDD.n1982 GND 0.006693f
C4295 VDD.n1983 GND 0.005387f
C4296 VDD.n1984 GND 0.006693f
C4297 VDD.n1985 GND 0.005387f
C4298 VDD.n1986 GND 0.006693f
C4299 VDD.n1987 GND 0.477993f
C4300 VDD.n1988 GND 0.006693f
C4301 VDD.n1989 GND 0.005387f
C4302 VDD.n1990 GND 0.006693f
C4303 VDD.n1991 GND 0.005387f
C4304 VDD.n1992 GND 0.006693f
C4305 VDD.t114 GND 0.238997f
C4306 VDD.n1993 GND 0.006693f
C4307 VDD.n1994 GND 0.005387f
C4308 VDD.n1995 GND 0.006693f
C4309 VDD.n1996 GND 0.005387f
C4310 VDD.n1997 GND 0.006693f
C4311 VDD.n1998 GND 0.477993f
C4312 VDD.n1999 GND 0.430194f
C4313 VDD.n2000 GND 0.006693f
C4314 VDD.n2001 GND 0.005387f
C4315 VDD.n2002 GND 0.006693f
C4316 VDD.n2003 GND 0.005387f
C4317 VDD.n2004 GND 0.006693f
C4318 VDD.n2005 GND 0.477993f
C4319 VDD.n2006 GND 0.006693f
C4320 VDD.n2007 GND 0.005387f
C4321 VDD.n2008 GND 0.006693f
C4322 VDD.n2009 GND 0.005387f
C4323 VDD.n2010 GND 0.006693f
C4324 VDD.n2011 GND 0.477993f
C4325 VDD.n2012 GND 0.006693f
C4326 VDD.n2013 GND 0.005387f
C4327 VDD.n2014 GND 0.006693f
C4328 VDD.n2015 GND 0.005387f
C4329 VDD.n2016 GND 0.006693f
C4330 VDD.n2017 GND 0.477993f
C4331 VDD.n2018 GND 0.006693f
C4332 VDD.n2019 GND 0.005387f
C4333 VDD.n2020 GND 0.006693f
C4334 VDD.n2021 GND 0.005387f
C4335 VDD.n2022 GND 0.006693f
C4336 VDD.n2023 GND 0.477993f
C4337 VDD.n2024 GND 0.006693f
C4338 VDD.n2025 GND 0.005387f
C4339 VDD.t116 GND 0.091115f
C4340 VDD.t137 GND 0.016539f
C4341 VDD.t103 GND 0.016539f
C4342 VDD.n2026 GND 0.062673f
C4343 VDD.n2027 GND 0.698762f
C4344 VDD.t134 GND 0.016539f
C4345 VDD.t155 GND 0.016539f
C4346 VDD.n2028 GND 0.062673f
C4347 VDD.n2029 GND 0.429343f
C4348 VDD.t130 GND 0.016539f
C4349 VDD.t153 GND 0.016539f
C4350 VDD.n2030 GND 0.062673f
C4351 VDD.n2031 GND 0.460012f
C4352 VDD.t113 GND 0.091115f
C4353 VDD.t133 GND 0.016539f
C4354 VDD.t156 GND 0.016539f
C4355 VDD.n2032 GND 0.062673f
C4356 VDD.n2033 GND 0.698762f
C4357 VDD.t132 GND 0.016539f
C4358 VDD.t150 GND 0.016539f
C4359 VDD.n2034 GND 0.062673f
C4360 VDD.n2035 GND 0.429343f
C4361 VDD.t124 GND 0.016539f
C4362 VDD.t148 GND 0.016539f
C4363 VDD.n2036 GND 0.062673f
C4364 VDD.n2037 GND 0.442907f
C4365 VDD.n2038 GND 0.305579f
C4366 VDD.t144 GND 0.091115f
C4367 VDD.t115 GND 0.016539f
C4368 VDD.t117 GND 0.016539f
C4369 VDD.n2039 GND 0.062673f
C4370 VDD.n2040 GND 0.698762f
C4371 VDD.t136 GND 0.016539f
C4372 VDD.t111 GND 0.016539f
C4373 VDD.n2041 GND 0.062673f
C4374 VDD.n2042 GND 0.429343f
C4375 VDD.t121 GND 0.016539f
C4376 VDD.t127 GND 0.016539f
C4377 VDD.n2043 GND 0.062673f
C4378 VDD.n2044 GND 0.442907f
C4379 VDD.n2045 GND 0.442725f
C4380 VDD.n2046 GND 4.10157f
C4381 VDD.n2047 GND 0.409661f
C4382 VDD.n2048 GND 0.005387f
C4383 VDD.n2049 GND 0.006693f
C4384 VDD.t110 GND 0.238997f
C4385 VDD.n2050 GND 0.006693f
C4386 VDD.n2051 GND 0.005387f
C4387 VDD.n2052 GND 0.006693f
C4388 VDD.n2053 GND 0.005387f
C4389 VDD.n2054 GND 0.006693f
C4390 VDD.n2055 GND 0.477993f
C4391 VDD.n2056 GND 0.358495f
C4392 VDD.n2057 GND 0.006693f
C4393 VDD.n2058 GND 0.005387f
C4394 VDD.n2059 GND 0.006693f
C4395 VDD.n2060 GND 0.005387f
C4396 VDD.n2061 GND 0.006693f
C4397 VDD.n2062 GND 0.477993f
C4398 VDD.n2063 GND 0.006693f
C4399 VDD.n2064 GND 0.005387f
C4400 VDD.n2065 GND 0.006693f
C4401 VDD.n2066 GND 0.005387f
C4402 VDD.n2067 GND 0.006693f
C4403 VDD.n2068 GND 0.477993f
C4404 VDD.n2069 GND 0.006693f
C4405 VDD.n2070 GND 0.005387f
C4406 VDD.n2071 GND 0.006693f
C4407 VDD.n2072 GND 0.005387f
C4408 VDD.n2073 GND 0.006693f
C4409 VDD.n2074 GND 0.477993f
C4410 VDD.n2075 GND 0.006693f
C4411 VDD.n2076 GND 0.005387f
C4412 VDD.n2077 GND 0.006693f
C4413 VDD.n2078 GND 0.005387f
C4414 VDD.n2079 GND 0.006693f
C4415 VDD.n2080 GND 0.477993f
C4416 VDD.n2081 GND 0.006693f
C4417 VDD.n2082 GND 0.005387f
C4418 VDD.n2083 GND 0.006693f
C4419 VDD.n2084 GND 0.005387f
C4420 VDD.n2085 GND 0.006693f
C4421 VDD.t131 GND 0.238997f
C4422 VDD.n2086 GND 0.006693f
C4423 VDD.n2087 GND 0.005387f
C4424 VDD.n2088 GND 0.006693f
C4425 VDD.n2089 GND 0.005387f
C4426 VDD.n2090 GND 0.006693f
C4427 VDD.n2091 GND 0.477993f
C4428 VDD.n2092 GND 0.286796f
C4429 VDD.n2093 GND 0.006693f
C4430 VDD.n2094 GND 0.005387f
C4431 VDD.n2095 GND 0.006693f
C4432 VDD.n2096 GND 0.005387f
C4433 VDD.n2097 GND 0.006693f
C4434 VDD.n2098 GND 0.477993f
C4435 VDD.n2099 GND 0.006693f
C4436 VDD.n2100 GND 0.005387f
C4437 VDD.n2101 GND 0.006693f
C4438 VDD.n2102 GND 0.005387f
C4439 VDD.n2103 GND 0.006693f
C4440 VDD.n2104 GND 0.477993f
C4441 VDD.n2105 GND 0.006693f
C4442 VDD.n2106 GND 0.005387f
C4443 VDD.n2107 GND 0.006693f
C4444 VDD.n2108 GND 0.005387f
C4445 VDD.n2109 GND 0.006693f
C4446 VDD.n2110 GND 0.477993f
C4447 VDD.n2111 GND 0.006693f
C4448 VDD.n2112 GND 0.005387f
C4449 VDD.n2113 GND 0.006693f
C4450 VDD.n2114 GND 0.005387f
C4451 VDD.n2115 GND 0.006693f
C4452 VDD.n2116 GND 0.477993f
C4453 VDD.n2117 GND 0.006693f
C4454 VDD.n2118 GND 0.005387f
C4455 VDD.n2119 GND 0.006693f
C4456 VDD.n2120 GND 0.005387f
C4457 VDD.n2121 GND 0.006693f
C4458 VDD.n2122 GND 0.262896f
C4459 VDD.n2123 GND 0.006693f
C4460 VDD.n2124 GND 0.005387f
C4461 VDD.n2125 GND 0.006693f
C4462 VDD.n2126 GND 0.005387f
C4463 VDD.n2127 GND 0.006693f
C4464 VDD.n2128 GND 0.477993f
C4465 VDD.t126 GND 0.238997f
C4466 VDD.n2129 GND 0.006693f
C4467 VDD.n2130 GND 0.005387f
C4468 VDD.n2131 GND 0.006693f
C4469 VDD.n2132 GND 0.005387f
C4470 VDD.n2133 GND 0.006693f
C4471 VDD.n2134 GND 0.477993f
C4472 VDD.n2135 GND 0.006693f
C4473 VDD.n2136 GND 0.005387f
C4474 VDD.n2137 GND 0.006693f
C4475 VDD.n2138 GND 0.005387f
C4476 VDD.n2139 GND 0.006693f
C4477 VDD.n2140 GND 0.477993f
C4478 VDD.n2141 GND 0.006693f
C4479 VDD.n2142 GND 0.005387f
C4480 VDD.n2143 GND 0.006693f
C4481 VDD.n2144 GND 0.005387f
C4482 VDD.n2145 GND 0.006693f
C4483 VDD.n2146 GND 0.477993f
C4484 VDD.n2147 GND 0.006693f
C4485 VDD.n2148 GND 0.005387f
C4486 VDD.n2149 GND 0.006693f
C4487 VDD.n2150 GND 0.005387f
C4488 VDD.n2151 GND 0.006693f
C4489 VDD.n2152 GND 0.477993f
C4490 VDD.n2153 GND 0.006693f
C4491 VDD.n2154 GND 0.005387f
C4492 VDD.n2155 GND 0.006693f
C4493 VDD.n2156 GND 0.005387f
C4494 VDD.n2157 GND 0.006693f
C4495 VDD.n2158 GND 0.334595f
C4496 VDD.n2159 GND 0.006693f
C4497 VDD.n2160 GND 0.005387f
C4498 VDD.n2161 GND 0.006693f
C4499 VDD.n2162 GND 0.005387f
C4500 VDD.n2163 GND 0.006693f
C4501 VDD.n2164 GND 0.477993f
C4502 VDD.t120 GND 0.238997f
C4503 VDD.n2165 GND 0.006693f
C4504 VDD.n2166 GND 0.005387f
C4505 VDD.n2167 GND 0.006693f
C4506 VDD.n2168 GND 0.005387f
C4507 VDD.n2169 GND 0.006693f
C4508 VDD.n2170 GND 0.477993f
C4509 VDD.n2171 GND 0.006693f
C4510 VDD.n2172 GND 0.005387f
C4511 VDD.n2173 GND 0.006693f
C4512 VDD.n2174 GND 0.005387f
C4513 VDD.n2175 GND 0.006693f
C4514 VDD.n2176 GND 0.477993f
C4515 VDD.n2177 GND 0.006693f
C4516 VDD.n2178 GND 0.005387f
C4517 VDD.n2179 GND 0.006693f
C4518 VDD.n2180 GND 0.005387f
C4519 VDD.n2181 GND 0.006693f
C4520 VDD.n2182 GND 0.477993f
C4521 VDD.n2183 GND 0.006693f
C4522 VDD.n2184 GND 0.005387f
C4523 VDD.n2185 GND 0.006693f
C4524 VDD.n2186 GND 0.005387f
C4525 VDD.n2187 GND 0.006693f
C4526 VDD.n2188 GND 0.477993f
C4527 VDD.n2189 GND 0.006693f
C4528 VDD.n2190 GND 0.005387f
C4529 VDD.n2191 GND 0.006693f
C4530 VDD.n2192 GND 0.005387f
C4531 VDD.n2193 GND 0.006693f
C4532 VDD.n2194 GND 0.477993f
C4533 VDD.n2195 GND 0.006693f
C4534 VDD.n2196 GND 0.005387f
C4535 VDD.n2197 GND 0.006693f
C4536 VDD.n2198 GND 0.005387f
C4537 VDD.n2199 GND 0.006693f
C4538 VDD.n2200 GND 0.477993f
C4539 VDD.n2201 GND 0.006693f
C4540 VDD.n2202 GND 0.005387f
C4541 VDD.n2203 GND 0.006693f
C4542 VDD.n2204 GND 0.005387f
C4543 VDD.n2205 GND 0.006693f
C4544 VDD.t33 GND 0.238997f
C4545 VDD.n2206 GND 0.006693f
C4546 VDD.n2207 GND 0.005387f
C4547 VDD.n2208 GND 0.006693f
C4548 VDD.n2209 GND 0.005387f
C4549 VDD.n2210 GND 0.006693f
C4550 VDD.n2211 GND 0.477993f
C4551 VDD.n2212 GND 0.348935f
C4552 VDD.n2213 GND 0.006693f
C4553 VDD.n2214 GND 0.005387f
C4554 VDD.n2215 GND 0.006693f
C4555 VDD.n2216 GND 0.005387f
C4556 VDD.n2217 GND 0.006693f
C4557 VDD.n2218 GND 0.477993f
C4558 VDD.n2219 GND 0.006693f
C4559 VDD.n2220 GND 0.005387f
C4560 VDD.n2221 GND 0.01598f
C4561 VDD.n2222 GND 0.004471f
C4562 VDD.n2223 GND 0.01598f
C4563 VDD.n2224 GND 0.70265f
C4564 VDD.n2225 GND 0.01598f
C4565 VDD.n2226 GND 0.004471f
C4566 VDD.n2227 GND 0.006693f
C4567 VDD.n2228 GND 0.005387f
C4568 VDD.n2229 GND 0.006693f
C4569 VDD.n2247 GND 0.016349f
C4570 VDD.n2248 GND 0.006693f
C4571 VDD.n2249 GND 0.005387f
C4572 VDD.n2250 GND 0.006693f
C4573 VDD.n2251 GND 0.006693f
C4574 VDD.n2252 GND 0.006693f
C4575 VDD.n2253 GND 0.006693f
C4576 VDD.n2254 GND 0.006693f
C4577 VDD.n2255 GND 0.005387f
C4578 VDD.n2256 GND 0.006693f
C4579 VDD.n2257 GND 0.006693f
C4580 VDD.n2258 GND 0.006693f
C4581 VDD.n2259 GND 0.006693f
C4582 VDD.t35 GND 0.118593f
C4583 VDD.t32 GND 0.540868f
C4584 VDD.n2260 GND 0.08957f
C4585 VDD.t34 GND 0.077791f
C4586 VDD.n2261 GND 0.092102f
C4587 VDD.n2262 GND 0.007407f
C4588 VDD.n2263 GND 0.006693f
C4589 VDD.n2264 GND 0.006693f
C4590 VDD.n2265 GND 0.006693f
C4591 VDD.n2266 GND 0.006693f
C4592 VDD.n2267 GND 0.005387f
C4593 VDD.n2268 GND 0.006693f
C4594 VDD.n2269 GND 0.006693f
C4595 VDD.n2270 GND 0.006693f
C4596 VDD.n2271 GND 0.006693f
C4597 VDD.n2272 GND 0.006693f
C4598 VDD.n2273 GND 0.005387f
C4599 VDD.n2274 GND 0.006693f
C4600 VDD.n2275 GND 0.006693f
C4601 VDD.n2276 GND 0.006693f
C4602 VDD.n2277 GND 0.006693f
C4603 VDD.n2278 GND 0.006693f
C4604 VDD.n2279 GND 0.005387f
C4605 VDD.n2280 GND 0.006693f
C4606 VDD.n2281 GND 0.006693f
C4607 VDD.n2282 GND 0.006693f
C4608 VDD.n2283 GND 0.006693f
C4609 VDD.n2284 GND 0.006693f
C4610 VDD.n2285 GND 0.005387f
C4611 VDD.n2286 GND 0.006693f
C4612 VDD.n2287 GND 0.006693f
C4613 VDD.n2288 GND 0.006693f
C4614 VDD.n2289 GND 0.006693f
C4615 VDD.n2290 GND 0.006693f
C4616 VDD.n2291 GND 0.005387f
C4617 VDD.n2292 GND 0.006693f
C4618 VDD.n2293 GND 0.006693f
C4619 VDD.n2294 GND 0.006693f
C4620 VDD.n2295 GND 0.006693f
C4621 VDD.n2296 GND 0.006693f
C4622 VDD.n2297 GND 0.005387f
C4623 VDD.n2298 GND 0.006693f
C4624 VDD.n2299 GND 0.006693f
C4625 VDD.n2300 GND 0.006693f
C4626 VDD.n2301 GND 0.006693f
C4627 VDD.n2302 GND 0.016349f
C4628 VDD.n2303 GND 0.002667f
C4629 VDD.t61 GND 0.118593f
C4630 VDD.t59 GND 0.540868f
C4631 VDD.n2304 GND 0.08957f
C4632 VDD.t60 GND 0.077791f
C4633 VDD.n2305 GND 0.092102f
C4634 VDD.n2306 GND 0.007407f
C4635 VDD.n2307 GND 0.002721f
C4636 VDD.n2308 GND 0.005387f
C4637 VDD.n2309 GND 0.006693f
C4638 VDD.n2310 GND 0.006693f
C4639 VDD.n2311 GND 0.006693f
C4640 VDD.n2312 GND 0.005387f
C4641 VDD.n2313 GND 0.005387f
C4642 VDD.n2314 GND 0.005387f
C4643 VDD.n2315 GND 0.006693f
C4644 VDD.n2316 GND 0.006693f
C4645 VDD.n2317 GND 0.006693f
C4646 VDD.n2318 GND 0.005387f
C4647 VDD.n2319 GND 0.005387f
C4648 VDD.n2320 GND 0.005387f
C4649 VDD.n2321 GND 0.006693f
C4650 VDD.n2322 GND 0.006693f
C4651 VDD.n2323 GND 0.006693f
C4652 VDD.n2324 GND 0.005387f
C4653 VDD.n2325 GND 0.003582f
C4654 VDD.t58 GND 0.118593f
C4655 VDD.t56 GND 0.540868f
C4656 VDD.n2326 GND 0.08957f
C4657 VDD.t57 GND 0.077791f
C4658 VDD.n2327 GND 0.092102f
C4659 VDD.n2328 GND 0.007407f
C4660 VDD.n2329 GND 0.002721f
C4661 VDD.n2330 GND 0.006693f
C4662 VDD.n2331 GND 0.006693f
C4663 VDD.n2332 GND 0.006693f
C4664 VDD.n2333 GND 0.005387f
C4665 VDD.n2334 GND 0.005387f
C4666 VDD.n2335 GND 0.005387f
C4667 VDD.n2336 GND 0.006693f
C4668 VDD.n2337 GND 0.006693f
C4669 VDD.n2338 GND 0.006693f
C4670 VDD.n2339 GND 0.005387f
C4671 VDD.n2340 GND 0.005387f
C4672 VDD.n2341 GND 0.005387f
C4673 VDD.n2342 GND 0.006693f
C4674 VDD.n2343 GND 0.006693f
C4675 VDD.n2344 GND 0.006693f
C4676 VDD.n2345 GND 0.005387f
C4677 VDD.n2346 GND 0.005387f
C4678 VDD.n2347 GND 0.003582f
C4679 VDD.n2348 GND 0.006693f
C4680 VDD.n2349 GND 0.006693f
C4681 VDD.n2350 GND 0.002721f
C4682 VDD.n2351 GND 0.005387f
C4683 VDD.n2352 GND 0.005387f
C4684 VDD.n2353 GND 0.006693f
C4685 VDD.n2354 GND 0.006693f
C4686 VDD.n2355 GND 0.006693f
C4687 VDD.n2356 GND 0.005387f
C4688 VDD.n2357 GND 0.005387f
C4689 VDD.n2358 GND 0.005387f
C4690 VDD.n2359 GND 0.006693f
C4691 VDD.n2360 GND 0.006693f
C4692 VDD.n2361 GND 0.006693f
C4693 VDD.n2362 GND 0.005387f
C4694 VDD.n2363 GND 0.006693f
C4695 VDD.n2364 GND 1.13762f
C4696 VDD.n2366 GND 0.016349f
C4697 VDD.n2367 GND 0.004471f
C4698 VDD.n2368 GND 0.016349f
C4699 VDD.n2369 GND 0.01598f
C4700 VDD.n2370 GND 0.006693f
C4701 VDD.n2371 GND 0.005387f
C4702 VDD.n2372 GND 0.006693f
C4703 VDD.n2373 GND 0.477993f
C4704 VDD.n2374 GND 0.006693f
C4705 VDD.n2375 GND 0.005387f
C4706 VDD.n2376 GND 0.006693f
C4707 VDD.n2377 GND 0.006693f
C4708 VDD.n2378 GND 0.006693f
C4709 VDD.n2379 GND 0.005387f
C4710 VDD.n2380 GND 0.006693f
C4711 VDD.n2381 GND 0.477993f
C4712 VDD.n2382 GND 0.006693f
C4713 VDD.n2383 GND 0.005387f
C4714 VDD.n2384 GND 0.006693f
C4715 VDD.n2385 GND 0.006693f
C4716 VDD.n2386 GND 0.006693f
C4717 VDD.n2387 GND 0.005387f
C4718 VDD.n2388 GND 0.006693f
C4719 VDD.n2389 GND 0.477993f
C4720 VDD.n2390 GND 0.006693f
C4721 VDD.n2391 GND 0.005387f
C4722 VDD.n2392 GND 0.006693f
C4723 VDD.n2393 GND 0.006693f
C4724 VDD.n2394 GND 0.006693f
C4725 VDD.n2395 GND 0.005387f
C4726 VDD.n2396 GND 0.006693f
C4727 VDD.n2397 GND 0.368055f
C4728 VDD.n2398 GND 0.006693f
C4729 VDD.n2399 GND 0.005387f
C4730 VDD.n2400 GND 0.006693f
C4731 VDD.n2401 GND 0.006693f
C4732 VDD.n2402 GND 0.006693f
C4733 VDD.n2403 GND 0.005387f
C4734 VDD.n2404 GND 0.006693f
C4735 VDD.n2405 GND 0.477993f
C4736 VDD.n2406 GND 0.006693f
C4737 VDD.n2407 GND 0.005387f
C4738 VDD.n2408 GND 0.006693f
C4739 VDD.n2409 GND 0.006693f
C4740 VDD.n2410 GND 0.006693f
C4741 VDD.n2411 GND 0.005387f
C4742 VDD.n2412 GND 0.006693f
C4743 VDD.n2413 GND 0.477993f
C4744 VDD.n2414 GND 0.006693f
C4745 VDD.n2415 GND 0.005387f
C4746 VDD.n2416 GND 0.006693f
C4747 VDD.n2417 GND 0.006693f
C4748 VDD.n2418 GND 0.006693f
C4749 VDD.n2419 GND 0.005387f
C4750 VDD.n2420 GND 0.006693f
C4751 VDD.n2421 GND 0.477993f
C4752 VDD.n2422 GND 0.006693f
C4753 VDD.n2423 GND 0.005387f
C4754 VDD.n2424 GND 0.006693f
C4755 VDD.n2425 GND 0.006693f
C4756 VDD.n2426 GND 0.006693f
C4757 VDD.n2427 GND 0.005387f
C4758 VDD.n2428 GND 0.006693f
C4759 VDD.n2429 GND 0.477993f
C4760 VDD.n2430 GND 0.006693f
C4761 VDD.n2431 GND 0.005387f
C4762 VDD.n2432 GND 0.006693f
C4763 VDD.n2433 GND 0.006693f
C4764 VDD.n2434 GND 0.006693f
C4765 VDD.n2435 GND 0.005387f
C4766 VDD.n2436 GND 0.006693f
C4767 VDD.n2437 GND 0.477993f
C4768 VDD.n2438 GND 0.006693f
C4769 VDD.n2439 GND 0.005387f
C4770 VDD.n2440 GND 0.006693f
C4771 VDD.n2441 GND 0.006693f
C4772 VDD.n2442 GND 0.006693f
C4773 VDD.n2443 GND 0.005387f
C4774 VDD.n2444 GND 0.006693f
C4775 VDD.n2445 GND 0.477993f
C4776 VDD.n2446 GND 0.006693f
C4777 VDD.n2447 GND 0.005387f
C4778 VDD.n2448 GND 0.006693f
C4779 VDD.n2449 GND 0.006693f
C4780 VDD.n2450 GND 0.006693f
C4781 VDD.n2451 GND 0.005387f
C4782 VDD.n2452 GND 0.006693f
C4783 VDD.n2453 GND 0.382394f
C4784 VDD.n2454 GND 0.006693f
C4785 VDD.n2455 GND 0.005387f
C4786 VDD.n2456 GND 0.006693f
C4787 VDD.n2457 GND 0.006693f
C4788 VDD.n2458 GND 0.006693f
C4789 VDD.n2459 GND 0.005387f
C4790 VDD.n2460 GND 0.006693f
C4791 VDD.n2461 GND 0.477993f
C4792 VDD.n2462 GND 0.006693f
C4793 VDD.n2463 GND 0.005387f
C4794 VDD.n2464 GND 0.006693f
C4795 VDD.n2465 GND 0.006693f
C4796 VDD.n2466 GND 0.006693f
C4797 VDD.n2467 GND 0.005387f
C4798 VDD.n2468 GND 0.006693f
C4799 VDD.n2469 GND 0.477993f
C4800 VDD.n2470 GND 0.006693f
C4801 VDD.n2471 GND 0.005387f
C4802 VDD.n2472 GND 0.006693f
C4803 VDD.n2473 GND 0.006693f
C4804 VDD.n2474 GND 0.006693f
C4805 VDD.n2475 GND 0.005387f
C4806 VDD.n2476 GND 0.006693f
C4807 VDD.n2477 GND 0.477993f
C4808 VDD.n2478 GND 0.006693f
C4809 VDD.n2479 GND 0.005387f
C4810 VDD.n2480 GND 0.006693f
C4811 VDD.n2481 GND 0.006693f
C4812 VDD.n2482 GND 0.006693f
C4813 VDD.n2483 GND 0.005387f
C4814 VDD.n2484 GND 0.006693f
C4815 VDD.n2485 GND 0.477993f
C4816 VDD.n2486 GND 0.006693f
C4817 VDD.n2487 GND 0.005387f
C4818 VDD.n2488 GND 0.006693f
C4819 VDD.n2489 GND 0.006693f
C4820 VDD.n2490 GND 0.006693f
C4821 VDD.n2491 GND 0.005387f
C4822 VDD.n2492 GND 0.006693f
C4823 VDD.n2493 GND 0.477993f
C4824 VDD.n2494 GND 0.006693f
C4825 VDD.n2495 GND 0.005387f
C4826 VDD.n2496 GND 0.006693f
C4827 VDD.n2497 GND 0.006693f
C4828 VDD.n2498 GND 0.006693f
C4829 VDD.n2499 GND 0.005387f
C4830 VDD.n2500 GND 0.006693f
C4831 VDD.n2501 GND 0.454093f
C4832 VDD.n2502 GND 0.006693f
C4833 VDD.n2503 GND 0.005387f
C4834 VDD.n2504 GND 0.006693f
C4835 VDD.n2505 GND 0.006693f
C4836 VDD.n2506 GND 0.006693f
C4837 VDD.n2507 GND 0.005387f
C4838 VDD.n2508 GND 0.006693f
C4839 VDD.n2509 GND 0.477993f
C4840 VDD.n2510 GND 0.006693f
C4841 VDD.n2511 GND 0.005387f
C4842 VDD.n2512 GND 0.006693f
C4843 VDD.n2513 GND 0.006693f
C4844 VDD.n2514 GND 0.006693f
C4845 VDD.n2515 GND 0.005387f
C4846 VDD.n2516 GND 0.006693f
C4847 VDD.n2517 GND 0.477993f
C4848 VDD.n2518 GND 0.006693f
C4849 VDD.n2519 GND 0.005387f
C4850 VDD.n2520 GND 0.006693f
C4851 VDD.n2521 GND 0.006693f
C4852 VDD.n2522 GND 0.006693f
C4853 VDD.n2523 GND 0.005387f
C4854 VDD.n2524 GND 0.006693f
C4855 VDD.n2525 GND 0.477993f
C4856 VDD.n2526 GND 0.006693f
C4857 VDD.n2527 GND 0.005387f
C4858 VDD.n2528 GND 0.006693f
C4859 VDD.n2529 GND 0.006693f
C4860 VDD.n2530 GND 0.006693f
C4861 VDD.n2531 GND 0.005387f
C4862 VDD.n2532 GND 0.006693f
C4863 VDD.n2533 GND 0.477993f
C4864 VDD.n2534 GND 0.006693f
C4865 VDD.n2535 GND 0.005387f
C4866 VDD.n2536 GND 0.006693f
C4867 VDD.n2537 GND 0.006693f
C4868 VDD.n2538 GND 0.006693f
C4869 VDD.n2539 GND 0.005387f
C4870 VDD.n2540 GND 0.006693f
C4871 VDD.n2541 GND 0.477993f
C4872 VDD.n2542 GND 0.006693f
C4873 VDD.n2543 GND 0.005387f
C4874 VDD.n2544 GND 0.006693f
C4875 VDD.n2545 GND 0.006693f
C4876 VDD.n2546 GND 0.006693f
C4877 VDD.n2547 GND 0.005387f
C4878 VDD.n2548 GND 0.006693f
C4879 VDD.n2549 GND 0.477993f
C4880 VDD.n2550 GND 0.006693f
C4881 VDD.n2551 GND 0.005387f
C4882 VDD.n2552 GND 0.006693f
C4883 VDD.n2553 GND 0.006693f
C4884 VDD.n2554 GND 0.006693f
C4885 VDD.n2555 GND 0.005387f
C4886 VDD.n2556 GND 0.006693f
C4887 VDD.n2557 GND 0.430194f
C4888 VDD.n2558 GND 0.006693f
C4889 VDD.n2559 GND 0.005387f
C4890 VDD.n2560 GND 0.006693f
C4891 VDD.n2561 GND 0.006693f
C4892 VDD.n2562 GND 0.006693f
C4893 VDD.n2563 GND 0.005387f
C4894 VDD.n2564 GND 0.006693f
C4895 VDD.n2565 GND 0.477993f
C4896 VDD.n2566 GND 0.006693f
C4897 VDD.n2567 GND 0.005387f
C4898 VDD.n2568 GND 0.006693f
C4899 VDD.n2569 GND 0.006693f
C4900 VDD.n2570 GND 0.006693f
C4901 VDD.n2571 GND 0.005387f
C4902 VDD.n2572 GND 0.006693f
C4903 VDD.n2573 GND 0.477993f
C4904 VDD.n2574 GND 0.006693f
C4905 VDD.n2575 GND 0.005387f
C4906 VDD.n2576 GND 0.006693f
C4907 VDD.n2577 GND 0.006693f
C4908 VDD.n2578 GND 0.006693f
C4909 VDD.n2579 GND 0.005387f
C4910 VDD.n2580 GND 0.006693f
C4911 VDD.n2581 GND 0.477993f
C4912 VDD.n2582 GND 0.006693f
C4913 VDD.n2583 GND 0.005387f
C4914 VDD.n2584 GND 0.006693f
C4915 VDD.n2585 GND 0.006693f
C4916 VDD.n2586 GND 0.006693f
C4917 VDD.n2587 GND 0.005387f
C4918 VDD.n2588 GND 0.006693f
C4919 VDD.n2589 GND 0.477993f
C4920 VDD.n2590 GND 0.006693f
C4921 VDD.n2591 GND 0.005387f
C4922 VDD.n2592 GND 0.006693f
C4923 VDD.n2593 GND 0.006693f
C4924 VDD.n2594 GND 0.005144f
C4925 VDD.n2595 GND 0.006693f
C4926 VDD.n2596 GND 0.005387f
C4927 VDD.n2597 GND 0.006693f
C4928 VDD.n2598 GND 0.477993f
C4929 VDD.n2599 GND 0.006693f
C4930 VDD.n2600 GND 0.005387f
C4931 VDD.n2601 GND 0.006693f
C4932 VDD.n2602 GND 0.006693f
C4933 VDD.n2603 GND 0.006693f
C4934 VDD.n2604 GND 0.005387f
C4935 VDD.n2605 GND 0.006693f
C4936 VDD.n2606 GND 0.358495f
C4937 VDD.n2607 GND 0.006693f
C4938 VDD.n2608 GND 0.005387f
C4939 VDD.n2609 GND 0.005144f
C4940 VDD.n2610 GND 0.006693f
C4941 VDD.n2611 GND 0.006693f
C4942 VDD.n2612 GND 0.005387f
C4943 VDD.n2613 GND 0.006693f
C4944 VDD.n2614 GND 0.477993f
C4945 VDD.n2615 GND 0.006693f
C4946 VDD.n2616 GND 0.005387f
C4947 VDD.n2617 GND 0.006693f
C4948 VDD.n2618 GND 0.006693f
C4949 VDD.n2619 GND 0.006693f
C4950 VDD.n2620 GND 0.005387f
C4951 VDD.n2621 GND 0.006693f
C4952 VDD.n2622 GND 0.477993f
C4953 VDD.n2623 GND 0.006693f
C4954 VDD.n2624 GND 0.005387f
C4955 VDD.n2625 GND 0.006693f
C4956 VDD.n2626 GND 0.006693f
C4957 VDD.n2627 GND 0.006693f
C4958 VDD.n2628 GND 0.005387f
C4959 VDD.n2629 GND 0.006693f
C4960 VDD.n2630 GND 0.477993f
C4961 VDD.n2631 GND 0.006693f
C4962 VDD.n2632 GND 0.005387f
C4963 VDD.n2633 GND 0.006693f
C4964 VDD.n2634 GND 0.006693f
C4965 VDD.n2635 GND 0.006693f
C4966 VDD.n2636 GND 0.005387f
C4967 VDD.n2637 GND 0.006693f
C4968 VDD.n2638 GND 0.477993f
C4969 VDD.n2639 GND 0.006693f
C4970 VDD.n2640 GND 0.005387f
C4971 VDD.n2641 GND 0.006693f
C4972 VDD.n2642 GND 0.006693f
C4973 VDD.n2643 GND 0.006693f
C4974 VDD.n2644 GND 0.005387f
C4975 VDD.n2645 GND 0.006693f
C4976 VDD.n2646 GND 0.477993f
C4977 VDD.n2647 GND 0.006693f
C4978 VDD.n2648 GND 0.005387f
C4979 VDD.n2649 GND 0.006693f
C4980 VDD.n2650 GND 0.006693f
C4981 VDD.n2651 GND 0.006693f
C4982 VDD.n2652 GND 0.005387f
C4983 VDD.n2653 GND 0.006693f
C4984 VDD.n2654 GND 0.286796f
C4985 VDD.n2655 GND 0.006693f
C4986 VDD.n2656 GND 0.005387f
C4987 VDD.n2657 GND 0.006693f
C4988 VDD.n2658 GND 0.006693f
C4989 VDD.n2659 GND 0.006693f
C4990 VDD.n2660 GND 0.005387f
C4991 VDD.n2661 GND 0.006693f
C4992 VDD.n2662 GND 0.477993f
C4993 VDD.n2663 GND 0.006693f
C4994 VDD.n2664 GND 0.005387f
C4995 VDD.n2665 GND 0.006693f
C4996 VDD.n2666 GND 0.006693f
C4997 VDD.n2667 GND 0.006693f
C4998 VDD.n2668 GND 0.005387f
C4999 VDD.n2669 GND 0.006693f
C5000 VDD.n2670 GND 0.477993f
C5001 VDD.n2671 GND 0.006693f
C5002 VDD.n2672 GND 0.005387f
C5003 VDD.n2673 GND 0.006693f
C5004 VDD.n2674 GND 0.006693f
C5005 VDD.n2675 GND 0.006693f
C5006 VDD.n2676 GND 0.005387f
C5007 VDD.n2677 GND 0.006693f
C5008 VDD.n2678 GND 0.477993f
C5009 VDD.n2679 GND 0.006693f
C5010 VDD.n2680 GND 0.005387f
C5011 VDD.n2681 GND 0.006693f
C5012 VDD.n2682 GND 0.006693f
C5013 VDD.n2683 GND 0.006693f
C5014 VDD.n2684 GND 0.005387f
C5015 VDD.n2685 GND 0.006693f
C5016 VDD.n2686 GND 0.477993f
C5017 VDD.n2687 GND 0.006693f
C5018 VDD.n2688 GND 0.005387f
C5019 VDD.n2689 GND 0.006693f
C5020 VDD.n2690 GND 0.006693f
C5021 VDD.n2691 GND 0.006693f
C5022 VDD.n2692 GND 0.005387f
C5023 VDD.n2693 GND 0.006693f
C5024 VDD.n2694 GND 0.477993f
C5025 VDD.n2695 GND 0.006693f
C5026 VDD.n2696 GND 0.005387f
C5027 VDD.n2697 GND 0.006693f
C5028 VDD.n2698 GND 0.006693f
C5029 VDD.n2699 GND 0.006693f
C5030 VDD.n2700 GND 0.005387f
C5031 VDD.n2701 GND 0.006693f
C5032 VDD.t102 GND 0.238997f
C5033 VDD.n2702 GND 0.262896f
C5034 VDD.n2703 GND 0.006693f
C5035 VDD.n2704 GND 0.005387f
C5036 VDD.n2705 GND 0.006693f
C5037 VDD.n2706 GND 0.006693f
C5038 VDD.n2707 GND 0.006693f
C5039 VDD.n2708 GND 0.005387f
C5040 VDD.n2709 GND 0.006693f
C5041 VDD.n2710 GND 0.477993f
C5042 VDD.n2711 GND 0.006693f
C5043 VDD.n2712 GND 0.005387f
C5044 VDD.n2713 GND 0.006693f
C5045 VDD.n2714 GND 0.006693f
C5046 VDD.n2715 GND 0.006693f
C5047 VDD.n2716 GND 0.005387f
C5048 VDD.n2717 GND 0.006693f
C5049 VDD.n2718 GND 0.477993f
C5050 VDD.n2719 GND 0.006693f
C5051 VDD.n2720 GND 0.005387f
C5052 VDD.n2721 GND 0.006693f
C5053 VDD.n2722 GND 0.006693f
C5054 VDD.n2723 GND 0.006693f
C5055 VDD.n2724 GND 0.005387f
C5056 VDD.n2725 GND 0.006693f
C5057 VDD.n2726 GND 0.477993f
C5058 VDD.n2727 GND 0.006693f
C5059 VDD.n2728 GND 0.005387f
C5060 VDD.n2729 GND 0.006693f
C5061 VDD.n2730 GND 0.006693f
C5062 VDD.n2731 GND 0.006693f
C5063 VDD.n2732 GND 0.005387f
C5064 VDD.n2733 GND 0.006693f
C5065 VDD.n2734 GND 0.477993f
C5066 VDD.n2735 GND 0.006693f
C5067 VDD.n2736 GND 0.005387f
C5068 VDD.n2737 GND 0.006693f
C5069 VDD.n2738 GND 0.006693f
C5070 VDD.n2739 GND 0.006693f
C5071 VDD.n2740 GND 0.005387f
C5072 VDD.n2741 GND 0.006693f
C5073 VDD.n2742 GND 0.477993f
C5074 VDD.n2743 GND 0.006693f
C5075 VDD.n2744 GND 0.005387f
C5076 VDD.n2745 GND 0.006693f
C5077 VDD.n2746 GND 0.006693f
C5078 VDD.n2747 GND 0.006693f
C5079 VDD.n2748 GND 0.005387f
C5080 VDD.n2749 GND 0.006693f
C5081 VDD.t112 GND 0.238997f
C5082 VDD.n2750 GND 0.334595f
C5083 VDD.n2751 GND 0.006693f
C5084 VDD.n2752 GND 0.005387f
C5085 VDD.n2753 GND 0.006693f
C5086 VDD.n2754 GND 0.006693f
C5087 VDD.n2755 GND 0.006693f
C5088 VDD.n2756 GND 0.005387f
C5089 VDD.n2757 GND 0.006693f
C5090 VDD.n2758 GND 0.477993f
C5091 VDD.n2759 GND 0.006693f
C5092 VDD.n2760 GND 0.005387f
C5093 VDD.n2761 GND 0.006693f
C5094 VDD.n2762 GND 0.006693f
C5095 VDD.n2763 GND 0.006693f
C5096 VDD.n2764 GND 0.005387f
C5097 VDD.n2765 GND 0.006693f
C5098 VDD.n2766 GND 0.477993f
C5099 VDD.n2767 GND 0.006693f
C5100 VDD.n2768 GND 0.005387f
C5101 VDD.n2769 GND 0.006693f
C5102 VDD.n2770 GND 0.006693f
C5103 VDD.n2771 GND 0.006693f
C5104 VDD.n2772 GND 0.005387f
C5105 VDD.n2773 GND 0.006693f
C5106 VDD.n2774 GND 0.477993f
C5107 VDD.n2775 GND 0.006693f
C5108 VDD.n2776 GND 0.005387f
C5109 VDD.n2777 GND 0.006693f
C5110 VDD.n2778 GND 0.006693f
C5111 VDD.n2779 GND 0.006693f
C5112 VDD.n2780 GND 0.005387f
C5113 VDD.n2781 GND 0.006693f
C5114 VDD.n2782 GND 0.477993f
C5115 VDD.n2783 GND 0.006693f
C5116 VDD.n2784 GND 0.005387f
C5117 VDD.n2785 GND 0.006693f
C5118 VDD.n2786 GND 0.006693f
C5119 VDD.n2787 GND 0.006693f
C5120 VDD.n2788 GND 0.005387f
C5121 VDD.n2789 GND 0.006693f
C5122 VDD.n2790 GND 0.477993f
C5123 VDD.n2791 GND 0.006693f
C5124 VDD.n2792 GND 0.005387f
C5125 VDD.n2793 GND 0.006693f
C5126 VDD.n2794 GND 0.006693f
C5127 VDD.n2795 GND 0.006693f
C5128 VDD.n2796 GND 0.005387f
C5129 VDD.n2797 GND 0.006693f
C5130 VDD.n2798 GND 0.477993f
C5131 VDD.n2799 GND 0.006693f
C5132 VDD.n2800 GND 0.005387f
C5133 VDD.n2801 GND 0.006693f
C5134 VDD.n2802 GND 0.006693f
C5135 VDD.n2803 GND 0.006693f
C5136 VDD.n2804 GND 0.005387f
C5137 VDD.n2805 GND 0.006693f
C5138 VDD.n2806 GND 0.477993f
C5139 VDD.n2807 GND 0.006693f
C5140 VDD.n2808 GND 0.005387f
C5141 VDD.n2809 GND 0.006693f
C5142 VDD.n2810 GND 0.006693f
C5143 VDD.n2811 GND 0.006693f
C5144 VDD.n2812 GND 0.006693f
C5145 VDD.n2813 GND 0.005387f
C5146 VDD.n2814 GND 0.006693f
C5147 VDD.n2815 GND 0.348935f
C5148 VDD.n2816 GND 0.006693f
C5149 VDD.n2817 GND 0.005387f
C5150 VDD.n2818 GND 0.006693f
C5151 VDD.n2819 GND 0.006693f
C5152 VDD.n2820 GND 0.006693f
C5153 VDD.n2821 GND 0.005387f
C5154 VDD.n2822 GND 0.006693f
C5155 VDD.n2823 GND 0.477993f
C5156 VDD.n2824 GND 0.006693f
C5157 VDD.n2825 GND 0.006693f
C5158 VDD.n2826 GND 0.005387f
C5159 VDD.n2827 GND 0.006693f
C5160 VDD.n2828 GND 0.006693f
C5161 VDD.n2829 GND 0.01249f
C5162 VDD.n2830 GND 0.013326f
C5163 VDD.n2831 GND 0.006693f
C5164 VDD.n2832 GND 0.005387f
C5165 VDD.n2833 GND 0.006693f
C5166 VDD.n2834 GND 0.477993f
C5167 VDD.n2835 GND 0.477993f
C5168 VDD.n2836 GND 0.006693f
C5169 VDD.n2837 GND 0.005387f
C5170 VDD.n2838 GND 0.006693f
C5171 VDD.n2839 GND 0.006693f
C5172 VDD.n2840 GND 0.01341f
C5173 VDD.n2841 GND 0.004471f
C5174 VDD.n2842 GND 0.01598f
C5175 VDD.n2843 GND 0.016349f
C5176 VDD.n2844 GND 0.004471f
C5177 VDD.n2845 GND 0.002978f
C5178 VDD.n2846 GND 0.003347f
C5179 VDD.n2847 GND 0.005387f
C5180 VDD.n2848 GND 0.006693f
C5181 VDD.n2849 GND 0.006693f
C5182 VDD.n2850 GND 0.005387f
C5183 VDD.n2851 GND 0.006693f
C5184 VDD.n2852 GND 0.006693f
C5185 VDD.n2853 GND 0.005387f
C5186 VDD.n2854 GND 0.003347f
C5187 VDD.n2855 GND 0.003347f
C5188 VDD.n2856 GND 0.003347f
C5189 VDD.n2857 GND 0.005387f
C5190 VDD.n2858 GND 0.006693f
C5191 VDD.n2859 GND 0.006693f
C5192 VDD.n2860 GND 0.005387f
C5193 VDD.n2861 GND 0.006693f
C5194 VDD.n2862 GND 0.006693f
C5195 VDD.n2863 GND 0.005387f
C5196 VDD.n2864 GND 0.003347f
C5197 VDD.n2865 GND 0.003347f
C5198 VDD.n2866 GND 0.003347f
C5199 VDD.n2867 GND 0.005387f
C5200 VDD.n2868 GND 0.006693f
C5201 VDD.n2869 GND 0.006693f
C5202 VDD.n2870 GND 0.002721f
C5203 VDD.t37 GND 0.118593f
C5204 VDD.t36 GND 0.540868f
C5205 VDD.n2871 GND 0.08957f
C5206 VDD.t38 GND 0.077791f
C5207 VDD.n2872 GND 0.092102f
C5208 VDD.n2873 GND 0.007407f
C5209 VDD.n2874 GND 0.006693f
C5210 VDD.n2875 GND 0.006693f
C5211 VDD.n2876 GND 0.003582f
C5212 VDD.n2877 GND 0.003347f
C5213 VDD.n2878 GND 0.003347f
C5214 VDD.n2879 GND 0.003347f
C5215 VDD.n2880 GND 0.005387f
C5216 VDD.n2881 GND 0.006693f
C5217 VDD.n2882 GND 0.006693f
C5218 VDD.n2883 GND 0.005387f
C5219 VDD.n2884 GND 0.006693f
C5220 VDD.n2885 GND 0.006693f
C5221 VDD.n2886 GND 0.005387f
C5222 VDD.n2887 GND 0.003347f
C5223 VDD.n2888 GND 0.003347f
C5224 VDD.n2889 GND 0.003347f
C5225 VDD.n2890 GND 0.005387f
C5226 VDD.n2891 GND 0.006693f
C5227 VDD.n2892 GND 0.006693f
C5228 VDD.n2895 GND 0.006693f
C5229 VDD.n2898 GND 0.006693f
C5230 VDD.n2901 GND 0.006693f
C5231 VDD.n2904 GND 0.006693f
C5232 VDD.t89 GND 4.6915f
C5233 VDD.t74 GND 6.34775f
C5234 VDD.t78 GND 7.0265f
C5235 VDD.t73 GND 7.53078f
C5236 VDD.n2906 GND 4.14181f
C5237 VDD.n2908 GND 0.016349f
C5238 VDD.n2909 GND 0.002667f
C5239 VDD.n2910 GND 0.007407f
C5240 VDD.n2911 GND 0.002721f
C5241 VDD.n2912 GND 0.005387f
C5242 VDD.n2913 GND 0.003347f
C5243 VDD.n2914 GND 0.003347f
C5244 VDD.n2915 GND 0.003347f
C5245 VDD.n2916 GND 0.005387f
C5246 VDD.n2917 GND 0.005387f
C5247 VDD.n2918 GND 0.005387f
C5248 VDD.n2919 GND 0.003347f
C5249 VDD.n2920 GND 0.003347f
C5250 VDD.n2921 GND 0.003347f
C5251 VDD.n2922 GND 0.005387f
C5252 VDD.n2923 GND 0.005387f
C5253 VDD.n2924 GND 0.005387f
C5254 VDD.n2925 GND 0.003347f
C5255 VDD.n2926 GND 0.003347f
C5256 VDD.n2927 GND 0.003347f
C5257 VDD.n2928 GND 0.005387f
C5258 VDD.n2929 GND 0.003582f
C5259 VDD.n2930 GND 0.007407f
C5260 VDD.n2931 GND 0.002721f
C5261 VDD.n2932 GND 0.003347f
C5262 VDD.n2933 GND 0.003347f
C5263 VDD.n2934 GND 0.003347f
C5264 VDD.n2935 GND 0.005387f
C5265 VDD.n2936 GND 0.005387f
C5266 VDD.n2937 GND 0.005387f
C5267 VDD.n2938 GND 0.00251f
C5268 VDD.n2939 GND 0.061109f
C5269 VDD.n2940 GND 1.93121f
C5270 VDD.n2941 GND 0.189549f
C5271 VDD.n2942 GND 0.004551f
C5272 VDD.n2944 GND 0.004551f
C5273 VDD.n2946 GND 0.004551f
C5274 VDD.n2947 GND 0.004551f
C5275 VDD.n2948 GND 0.004551f
C5276 VDD.n2949 GND 0.004551f
C5277 VDD.n2950 GND 0.004551f
C5278 VDD.n2952 GND 0.004551f
C5279 VDD.n2953 GND 0.004551f
C5280 VDD.n2954 GND 0.004551f
C5281 VDD.n2955 GND 0.004551f
C5282 VDD.n2956 GND 0.004551f
C5283 VDD.n2957 GND 0.004551f
C5284 VDD.n2959 GND 0.004551f
C5285 VDD.n2960 GND 0.004551f
C5286 VDD.n2961 GND 0.011274f
C5287 VDD.n2962 GND 0.010814f
C5288 VDD.n2963 GND 0.010814f
C5289 VDD.n2964 GND 0.470823f
C5290 VDD.n2965 GND 0.010814f
C5291 VDD.n2966 GND 0.010814f
C5292 VDD.n2967 GND 0.004551f
C5293 VDD.n2968 GND 0.004551f
C5294 VDD.n2969 GND 0.004551f
C5295 VDD.n2970 GND 0.325035f
C5296 VDD.n2971 GND 0.004551f
C5297 VDD.n2972 GND 0.004551f
C5298 VDD.n2973 GND 0.004551f
C5299 VDD.n2974 GND 0.004551f
C5300 VDD.n2975 GND 0.004551f
C5301 VDD.n2976 GND 0.325035f
C5302 VDD.n2977 GND 0.004551f
C5303 VDD.n2978 GND 0.004551f
C5304 VDD.n2979 GND 0.004551f
C5305 VDD.n2980 GND 0.004551f
C5306 VDD.n2981 GND 0.004551f
C5307 VDD.n2982 GND 0.325035f
C5308 VDD.n2983 GND 0.004551f
C5309 VDD.n2984 GND 0.004551f
C5310 VDD.n2985 GND 0.004551f
C5311 VDD.n2986 GND 0.004551f
C5312 VDD.n2987 GND 0.004551f
C5313 VDD.n2988 GND 0.210317f
C5314 VDD.n2989 GND 0.004551f
C5315 VDD.n2990 GND 0.004551f
C5316 VDD.n2991 GND 0.004551f
C5317 VDD.n2992 GND 0.004551f
C5318 VDD.n2993 GND 0.004551f
C5319 VDD.n2994 GND 0.325035f
C5320 VDD.n2995 GND 0.004551f
C5321 VDD.n2996 GND 0.004551f
C5322 VDD.n2997 GND 0.004551f
C5323 VDD.n2998 GND 0.004551f
C5324 VDD.n2999 GND 0.004551f
C5325 VDD.n3000 GND 0.282016f
C5326 VDD.n3001 GND 0.004551f
C5327 VDD.n3002 GND 0.004551f
C5328 VDD.n3003 GND 0.004551f
C5329 VDD.n3004 GND 0.004551f
C5330 VDD.n3005 GND 0.004551f
C5331 VDD.n3006 GND 0.325035f
C5332 VDD.n3007 GND 0.004551f
C5333 VDD.n3008 GND 0.004551f
C5334 VDD.n3009 GND 0.004551f
C5335 VDD.n3010 GND 0.004551f
C5336 VDD.n3011 GND 0.004551f
C5337 VDD.n3012 GND 0.325035f
C5338 VDD.n3013 GND 0.004551f
C5339 VDD.n3014 GND 0.004551f
C5340 VDD.n3015 GND 0.004551f
C5341 VDD.n3016 GND 0.004551f
C5342 VDD.n3017 GND 0.004551f
C5343 VDD.n3018 GND 0.325035f
C5344 VDD.n3019 GND 0.004551f
C5345 VDD.n3020 GND 0.004551f
C5346 VDD.n3021 GND 0.004551f
C5347 VDD.n3022 GND 0.004551f
C5348 VDD.n3023 GND 0.004551f
C5349 VDD.n3024 GND 0.325035f
C5350 VDD.n3025 GND 0.004551f
C5351 VDD.n3026 GND 0.004551f
C5352 VDD.n3027 GND 0.004551f
C5353 VDD.n3028 GND 0.004551f
C5354 VDD.n3029 GND 0.004551f
C5355 VDD.n3030 GND 0.325035f
C5356 VDD.n3031 GND 0.004551f
C5357 VDD.n3032 GND 0.004551f
C5358 VDD.n3033 GND 0.004551f
C5359 VDD.n3034 GND 0.004551f
C5360 VDD.n3035 GND 0.004551f
C5361 VDD.n3036 GND 0.325035f
C5362 VDD.n3037 GND 0.004551f
C5363 VDD.n3038 GND 0.004551f
C5364 VDD.n3039 GND 0.004551f
C5365 VDD.n3040 GND 0.004551f
C5366 VDD.n3041 GND 0.004551f
C5367 VDD.n3042 GND 0.325035f
C5368 VDD.n3043 GND 0.004551f
C5369 VDD.n3044 GND 0.004551f
C5370 VDD.n3045 GND 0.004551f
C5371 VDD.n3046 GND 0.004551f
C5372 VDD.n3047 GND 0.004551f
C5373 VDD.n3048 GND 0.325035f
C5374 VDD.n3049 GND 0.004551f
C5375 VDD.n3050 GND 0.004551f
C5376 VDD.n3051 GND 0.004551f
C5377 VDD.n3052 GND 0.004551f
C5378 VDD.n3053 GND 0.004551f
C5379 VDD.n3054 GND 0.325035f
C5380 VDD.n3055 GND 0.004551f
C5381 VDD.n3056 GND 0.004551f
C5382 VDD.n3057 GND 0.004551f
C5383 VDD.n3058 GND 0.004551f
C5384 VDD.n3059 GND 0.004551f
C5385 VDD.n3060 GND 0.325035f
C5386 VDD.n3061 GND 0.004551f
C5387 VDD.n3062 GND 0.004551f
C5388 VDD.n3063 GND 0.004551f
C5389 VDD.n3064 GND 0.004551f
C5390 VDD.n3065 GND 0.004551f
C5391 VDD.n3066 GND 0.320255f
C5392 VDD.n3067 GND 0.004551f
C5393 VDD.n3068 GND 0.004551f
C5394 VDD.n3069 GND 0.004551f
C5395 VDD.n3070 GND 0.004551f
C5396 VDD.n3071 GND 0.004551f
C5397 VDD.n3072 GND 0.325035f
C5398 VDD.n3073 GND 0.004551f
C5399 VDD.n3074 GND 0.004551f
C5400 VDD.n3075 GND 0.004551f
C5401 VDD.n3076 GND 0.004551f
C5402 VDD.n3077 GND 0.004551f
C5403 VDD.n3078 GND 0.286796f
C5404 VDD.n3079 GND 0.004551f
C5405 VDD.n3080 GND 0.004551f
C5406 VDD.n3081 GND 0.004551f
C5407 VDD.n3082 GND 0.004551f
C5408 VDD.n3083 GND 0.004551f
C5409 VDD.n3084 GND 0.325035f
C5410 VDD.n3085 GND 0.004551f
C5411 VDD.n3086 GND 0.004551f
C5412 VDD.n3087 GND 0.004551f
C5413 VDD.n3088 GND 0.004551f
C5414 VDD.n3089 GND 0.004551f
C5415 VDD.n3090 GND 0.325035f
C5416 VDD.n3091 GND 0.004551f
C5417 VDD.n3092 GND 0.004551f
C5418 VDD.n3093 GND 0.004551f
C5419 VDD.n3094 GND 0.004551f
C5420 VDD.n3095 GND 0.004551f
C5421 VDD.n3096 GND 0.325035f
C5422 VDD.n3097 GND 0.004551f
C5423 VDD.n3098 GND 0.004551f
C5424 VDD.n3099 GND 0.004551f
C5425 VDD.n3100 GND 0.004551f
C5426 VDD.n3101 GND 0.004551f
C5427 VDD.n3102 GND 0.325035f
C5428 VDD.n3103 GND 0.004551f
C5429 VDD.n3104 GND 0.004551f
C5430 VDD.n3105 GND 0.004551f
C5431 VDD.n3106 GND 0.004551f
C5432 VDD.n3107 GND 0.004551f
C5433 VDD.n3108 GND 0.325035f
C5434 VDD.n3109 GND 0.004551f
C5435 VDD.n3110 GND 0.004551f
C5436 VDD.n3111 GND 0.004551f
C5437 VDD.n3112 GND 0.004551f
C5438 VDD.n3113 GND 0.004551f
C5439 VDD.n3114 GND 0.325035f
C5440 VDD.n3115 GND 0.004551f
C5441 VDD.n3116 GND 0.004551f
C5442 VDD.n3117 GND 0.004551f
C5443 VDD.n3118 GND 0.004551f
C5444 VDD.n3119 GND 0.004551f
C5445 VDD.n3120 GND 0.325035f
C5446 VDD.n3121 GND 0.004551f
C5447 VDD.n3122 GND 0.004551f
C5448 VDD.n3123 GND 0.004551f
C5449 VDD.n3124 GND 0.004551f
C5450 VDD.n3125 GND 0.004551f
C5451 VDD.n3126 GND 0.243776f
C5452 VDD.n3127 GND 0.004551f
C5453 VDD.n3128 GND 0.004551f
C5454 VDD.n3129 GND 0.004551f
C5455 VDD.n3130 GND 0.004551f
C5456 VDD.n3131 GND 0.004551f
C5457 VDD.n3132 GND 0.286796f
C5458 VDD.n3133 GND 0.004551f
C5459 VDD.n3134 GND 0.004551f
C5460 VDD.n3135 GND 0.004551f
C5461 VDD.n3136 GND 0.004551f
C5462 VDD.n3137 GND 0.004551f
C5463 VDD.n3138 GND 0.325035f
C5464 VDD.n3139 GND 0.004551f
C5465 VDD.n3140 GND 0.004551f
C5466 VDD.n3141 GND 0.004551f
C5467 VDD.n3142 GND 0.004551f
C5468 VDD.n3143 GND 0.004551f
C5469 VDD.n3144 GND 0.325035f
C5470 VDD.n3145 GND 0.004551f
C5471 VDD.n3146 GND 0.004551f
C5472 VDD.n3147 GND 0.004551f
C5473 VDD.n3148 GND 0.004551f
C5474 VDD.n3149 GND 0.004551f
C5475 VDD.n3150 GND 0.325035f
C5476 VDD.n3151 GND 0.004551f
C5477 VDD.n3152 GND 0.004551f
C5478 VDD.n3153 GND 0.004551f
C5479 VDD.n3154 GND 0.004551f
C5480 VDD.n3155 GND 0.004551f
C5481 VDD.n3156 GND 0.325035f
C5482 VDD.n3157 GND 0.004551f
C5483 VDD.n3158 GND 0.004551f
C5484 VDD.n3159 GND 0.004551f
C5485 VDD.n3160 GND 0.004551f
C5486 VDD.n3161 GND 0.004551f
C5487 VDD.n3162 GND 0.325035f
C5488 VDD.n3163 GND 0.004551f
C5489 VDD.n3164 GND 0.004551f
C5490 VDD.n3165 GND 0.004551f
C5491 VDD.n3166 GND 0.004551f
C5492 VDD.n3167 GND 0.004551f
C5493 VDD.n3168 GND 0.325035f
C5494 VDD.n3169 GND 0.004551f
C5495 VDD.n3170 GND 0.004551f
C5496 VDD.n3171 GND 0.004551f
C5497 VDD.n3172 GND 0.004551f
C5498 VDD.n3173 GND 0.004551f
C5499 VDD.n3174 GND 0.325035f
C5500 VDD.n3175 GND 0.004551f
C5501 VDD.n3176 GND 0.004551f
C5502 VDD.n3177 GND 0.004551f
C5503 VDD.n3178 GND 0.004551f
C5504 VDD.n3179 GND 0.004551f
C5505 VDD.n3180 GND 0.325035f
C5506 VDD.n3181 GND 0.004551f
C5507 VDD.n3182 GND 0.004551f
C5508 VDD.n3183 GND 0.004551f
C5509 VDD.n3184 GND 0.004551f
C5510 VDD.n3185 GND 0.004551f
C5511 VDD.n3186 GND 0.167298f
C5512 VDD.n3187 GND 0.004551f
C5513 VDD.n3188 GND 0.004551f
C5514 VDD.n3189 GND 0.004551f
C5515 VDD.n3190 GND 0.004551f
C5516 VDD.n3191 GND 0.004551f
C5517 VDD.n3192 GND 0.210317f
C5518 VDD.n3193 GND 0.004551f
C5519 VDD.n3194 GND 0.004551f
C5520 VDD.n3195 GND 0.004551f
C5521 VDD.n3196 GND 0.004551f
C5522 VDD.n3197 GND 0.004551f
C5523 VDD.n3198 GND 0.325035f
C5524 VDD.n3199 GND 0.004551f
C5525 VDD.n3200 GND 0.004551f
C5526 VDD.n3201 GND 0.004551f
C5527 VDD.n3202 GND 0.004551f
C5528 VDD.n3203 GND 0.004551f
C5529 VDD.n3204 GND 0.325035f
C5530 VDD.n3205 GND 0.004551f
C5531 VDD.n3206 GND 0.004551f
C5532 VDD.n3207 GND 0.004551f
C5533 VDD.n3208 GND 0.004551f
C5534 VDD.n3209 GND 0.004551f
C5535 VDD.n3210 GND 0.325035f
C5536 VDD.n3211 GND 0.004551f
C5537 VDD.n3212 GND 0.004551f
C5538 VDD.n3213 GND 0.004551f
C5539 VDD.n3214 GND 0.004551f
C5540 VDD.n3215 GND 0.004551f
C5541 VDD.n3216 GND 0.325035f
C5542 VDD.n3217 GND 0.004551f
C5543 VDD.n3218 GND 0.004551f
C5544 VDD.n3219 GND 0.004551f
C5545 VDD.n3220 GND 0.004551f
C5546 VDD.n3221 GND 0.004551f
C5547 VDD.n3222 GND 0.325035f
C5548 VDD.n3223 GND 0.004551f
C5549 VDD.n3224 GND 0.004551f
C5550 VDD.n3225 GND 0.004551f
C5551 VDD.n3226 GND 0.004551f
C5552 VDD.n3227 GND 0.004551f
C5553 VDD.n3228 GND 0.325035f
C5554 VDD.n3229 GND 0.004551f
C5555 VDD.n3230 GND 0.004551f
C5556 VDD.n3231 GND 0.004551f
C5557 VDD.n3232 GND 0.004551f
C5558 VDD.n3233 GND 0.004551f
C5559 VDD.n3234 GND 0.325035f
C5560 VDD.n3235 GND 0.004551f
C5561 VDD.n3236 GND 0.004551f
C5562 VDD.n3237 GND 0.004551f
C5563 VDD.n3238 GND 0.004551f
C5564 VDD.n3239 GND 0.004551f
C5565 VDD.n3240 GND 0.325035f
C5566 VDD.n3241 GND 0.004551f
C5567 VDD.n3242 GND 0.004551f
C5568 VDD.n3243 GND 0.004551f
C5569 VDD.n3244 GND 0.004551f
C5570 VDD.n3245 GND 0.004551f
C5571 VDD.n3246 GND 0.325035f
C5572 VDD.n3247 GND 0.004551f
C5573 VDD.n3248 GND 0.004551f
C5574 VDD.n3249 GND 0.004551f
C5575 VDD.n3250 GND 0.004551f
C5576 VDD.n3251 GND 0.004551f
C5577 VDD.n3252 GND 0.191197f
C5578 VDD.n3253 GND 0.004551f
C5579 VDD.n3254 GND 0.004551f
C5580 VDD.n3255 GND 0.004551f
C5581 VDD.n3256 GND 0.004551f
C5582 VDD.n3257 GND 0.004551f
C5583 VDD.n3258 GND 0.205537f
C5584 VDD.n3259 GND 0.004551f
C5585 VDD.n3260 GND 0.004551f
C5586 VDD.n3261 GND 0.004551f
C5587 VDD.n3262 GND 0.004551f
C5588 VDD.n3263 GND 0.004551f
C5589 VDD.n3264 GND 0.325035f
C5590 VDD.n3265 GND 0.004551f
C5591 VDD.n3266 GND 0.004551f
C5592 VDD.n3267 GND 0.004551f
C5593 VDD.n3268 GND 0.004551f
C5594 VDD.n3269 GND 0.004551f
C5595 VDD.n3270 GND 0.004551f
C5596 VDD.n3271 GND 0.004551f
C5597 VDD.n3272 GND 0.325035f
C5598 VDD.n3273 GND 0.004551f
C5599 VDD.n3274 GND 0.004551f
C5600 VDD.n3275 GND 0.004551f
C5601 VDD.n3276 GND 0.004551f
C5602 VDD.n3277 GND 0.004551f
C5603 VDD.n3278 GND 0.325035f
C5604 VDD.n3279 GND 0.004551f
C5605 VDD.n3280 GND 0.004551f
C5606 VDD.n3281 GND 0.004551f
C5607 VDD.n3282 GND 0.004551f
C5608 VDD.n3283 GND 0.004551f
C5609 VDD.n3284 GND 0.004551f
C5610 VDD.n3285 GND 0.004551f
C5611 VDD.n3286 GND 0.011323f
C5612 VDD.n3287 GND 0.010814f
C5613 VDD.n3288 GND 0.011274f
C5614 VDD.n3289 GND 0.010764f
C5615 VDD.n3290 GND 0.004551f
C5616 VDD.n3291 GND 0.004551f
C5617 VDD.n3292 GND 0.004551f
C5618 VDD.n3293 GND 0.004551f
C5619 VDD.n3294 GND 0.00261f
C5620 VDD.n3295 GND 0.004551f
C5621 VDD.n3296 GND 0.004551f
C5622 VDD.n3297 GND 0.004217f
C5623 VDD.n3298 GND 0.004551f
C5624 VDD.n3299 GND 0.004551f
C5625 VDD.n3300 GND 0.004551f
C5626 VDD.n3301 GND 0.004551f
C5627 VDD.n3302 GND 0.004551f
C5628 VDD.n3303 GND 0.004551f
C5629 VDD.n3304 GND 0.004551f
C5630 VDD.n3305 GND 0.004551f
C5631 VDD.n3306 GND 0.004551f
C5632 VDD.n3307 GND 0.004551f
C5633 VDD.n3308 GND 0.004551f
C5634 VDD.n3309 GND 0.004551f
C5635 VDD.n3310 GND 0.004551f
C5636 VDD.n3311 GND 0.004551f
C5637 VDD.n3312 GND 0.004551f
C5638 VDD.n3313 GND 0.004551f
C5639 VDD.n3314 GND 0.004551f
C5640 VDD.n3315 GND 0.004551f
C5641 VDD.n3316 GND 0.004551f
C5642 VDD.n3317 GND 0.004551f
C5643 VDD.n3318 GND 0.004551f
C5644 VDD.n3319 GND 0.004551f
C5645 VDD.n3320 GND 0.004551f
C5646 VDD.n3321 GND 0.004551f
C5647 VDD.n3322 GND 0.004551f
C5648 VDD.n3323 GND 0.004551f
C5649 VDD.n3324 GND 0.004551f
C5650 VDD.n3325 GND 0.004551f
C5651 VDD.n3326 GND 0.004551f
C5652 VDD.n3327 GND 0.004551f
C5653 VDD.n3328 GND 0.011274f
C5654 VDD.n3329 GND 0.010814f
C5655 VDD.n3330 GND 0.010814f
C5656 VDD.n3331 GND 0.004551f
C5657 VDD.n3332 GND 0.004551f
C5658 VDD.n3333 GND 0.004551f
C5659 VDD.n3334 GND 0.004551f
C5660 VDD.n3335 GND 0.325035f
C5661 VDD.n3336 GND 0.004551f
C5662 VDD.n3337 GND 0.004551f
C5663 VDD.n3338 GND 0.004551f
C5664 VDD.n3339 GND 0.004551f
C5665 VDD.n3340 GND 0.004551f
C5666 VDD.n3341 GND 0.325035f
C5667 VDD.n3342 GND 0.004551f
C5668 VDD.n3343 GND 0.010814f
C5669 VDD.n3344 GND 0.011274f
C5670 VDD.n3345 GND 0.010764f
C5671 VDD.n3346 GND 0.004551f
C5672 VDD.n3347 GND 0.004551f
C5673 VDD.n3348 GND 0.004551f
C5674 VDD.n3349 GND 0.004551f
C5675 VDD.n3350 GND 0.00261f
C5676 VDD.n3351 GND 0.004551f
C5677 VDD.n3352 GND 0.004551f
C5678 VDD.n3353 GND 0.004217f
C5679 VDD.n3354 GND 0.004551f
C5680 VDD.n3355 GND 0.004551f
C5681 VDD.n3356 GND 0.004551f
C5682 VDD.n3357 GND 0.004551f
C5683 VDD.n3358 GND 0.004551f
C5684 VDD.n3359 GND 0.004551f
C5685 VDD.n3360 GND 0.004551f
C5686 VDD.n3361 GND 0.004551f
C5687 VDD.n3362 GND 0.004551f
C5688 VDD.n3363 GND 0.004551f
C5689 VDD.n3364 GND 0.004551f
C5690 VDD.n3365 GND 0.004551f
C5691 VDD.n3366 GND 0.004551f
C5692 VDD.n3367 GND 0.004551f
C5693 VDD.n3368 GND 0.004551f
C5694 VDD.n3369 GND 0.004551f
C5695 VDD.n3370 GND 0.004551f
C5696 VDD.n3371 GND 0.004551f
C5697 VDD.n3372 GND 0.004551f
C5698 VDD.n3373 GND 0.004551f
C5699 VDD.n3374 GND 0.004551f
C5700 VDD.n3375 GND 0.004551f
C5701 VDD.n3376 GND 0.004551f
C5702 VDD.n3377 GND 0.004551f
C5703 VDD.n3378 GND 0.004551f
C5704 VDD.n3379 GND 0.004551f
C5705 VDD.n3380 GND 0.004551f
C5706 VDD.n3381 GND 0.004551f
C5707 VDD.n3382 GND 0.004551f
C5708 VDD.n3383 GND 0.011274f
C5709 VDD.n3384 GND 0.011274f
C5710 VDD.n3385 GND 2.04342f
C5711 VDD.n3386 GND 2.04342f
C5712 VDD.n3387 GND 0.011274f
C5713 VDD.n3388 GND 0.004551f
C5714 VDD.n3389 GND 0.004551f
C5715 VDD.n3390 GND 0.004551f
C5716 VDD.t68 GND 0.154197f
C5717 VDD.t66 GND 0.733149f
C5718 VDD.n3391 GND 0.09739f
C5719 VDD.t67 GND 0.103896f
C5720 VDD.n3392 GND 0.100617f
C5721 VDD.n3393 GND 0.004551f
C5722 VDD.n3394 GND 0.004551f
C5723 VDD.n3395 GND 0.004551f
C5724 VDD.n3396 GND 0.004551f
C5725 VDD.n3397 GND 0.004551f
C5726 VDD.n3398 GND 0.004551f
C5727 VDD.n3399 GND 0.004551f
C5728 VDD.n3400 GND 0.004551f
C5729 VDD.n3402 GND 0.004551f
C5730 VDD.n3403 GND 0.004551f
C5731 VDD.n3405 GND 0.004551f
C5732 VDD.n3406 GND 0.004551f
C5733 VDD.n3407 GND 0.004551f
C5734 VDD.n3408 GND 0.004551f
C5735 VDD.n3409 GND 0.004551f
C5736 VDD.n3411 GND 0.004551f
C5737 VDD.n3413 GND 0.004551f
C5738 VDD.n3414 GND 0.004551f
C5739 VDD.n3415 GND 0.004551f
C5740 VDD.n3416 GND 0.004551f
C5741 VDD.n3417 GND 0.004551f
C5742 VDD.n3419 GND 0.004551f
C5743 VDD.n3421 GND 0.004551f
C5744 VDD.n3422 GND 0.004551f
C5745 VDD.n3423 GND 0.004551f
C5746 VDD.n3424 GND 0.004551f
C5747 VDD.n3425 GND 0.004551f
C5748 VDD.n3427 GND 0.004551f
C5749 VDD.n3429 GND 0.004551f
C5750 VDD.n3430 GND 0.004551f
C5751 VDD.n3431 GND 0.004217f
C5752 VDD.n3432 GND 0.005616f
C5753 VDD.n3433 GND 0.00261f
C5754 VDD.n3434 GND 0.004551f
C5755 VDD.n3436 GND 0.004551f
C5756 VDD.n3438 GND 0.004551f
C5757 VDD.n3439 GND 0.004551f
C5758 VDD.n3440 GND 0.011274f
C5759 VDD.n3441 GND 0.004551f
C5760 VDD.n3442 GND 0.004551f
C5761 VDD.n3443 GND 0.004551f
C5762 VDD.n3444 GND 0.004551f
C5763 VDD.n3445 GND 0.004551f
C5764 VDD.n3446 GND 0.004551f
C5765 VDD.n3447 GND 0.004551f
C5766 VDD.n3448 GND 0.004551f
C5767 VDD.n3449 GND 0.004551f
C5768 VDD.n3450 GND 0.004551f
C5769 VDD.n3451 GND 0.004551f
C5770 VDD.n3452 GND 0.004551f
C5771 VDD.n3453 GND 0.004551f
C5772 VDD.n3454 GND 0.004551f
C5773 VDD.n3455 GND 0.004551f
C5774 VDD.n3456 GND 0.004551f
C5775 VDD.n3457 GND 0.004551f
C5776 VDD.n3458 GND 0.004551f
C5777 VDD.n3459 GND 0.004551f
C5778 VDD.n3460 GND 0.004551f
C5779 VDD.n3461 GND 0.004551f
C5780 VDD.n3462 GND 0.004551f
C5781 VDD.n3463 GND 0.004551f
C5782 VDD.n3464 GND 0.004551f
C5783 VDD.n3465 GND 0.004551f
C5784 VDD.n3466 GND 0.004551f
C5785 VDD.n3467 GND 0.004551f
C5786 VDD.n3468 GND 0.004551f
C5787 VDD.n3469 GND 0.004551f
C5788 VDD.n3470 GND 0.004551f
C5789 VDD.n3471 GND 0.004551f
C5790 VDD.n3472 GND 0.004551f
C5791 VDD.n3473 GND 0.004551f
C5792 VDD.n3474 GND 0.004551f
C5793 VDD.n3475 GND 0.004551f
C5794 VDD.n3476 GND 0.004551f
C5795 VDD.n3477 GND 0.004551f
C5796 VDD.n3478 GND 0.004551f
C5797 VDD.n3479 GND 0.004551f
C5798 VDD.n3480 GND 0.004551f
C5799 VDD.n3481 GND 0.004551f
C5800 VDD.n3482 GND 0.004551f
C5801 VDD.n3483 GND 0.004551f
C5802 VDD.n3484 GND 0.004551f
C5803 VDD.n3485 GND 0.004551f
C5804 VDD.n3486 GND 0.004551f
C5805 VDD.n3487 GND 0.004551f
C5806 VDD.n3488 GND 0.004551f
C5807 VDD.n3489 GND 0.004551f
C5808 VDD.n3490 GND 0.004551f
C5809 VDD.n3491 GND 0.004551f
C5810 VDD.n3492 GND 0.004551f
C5811 VDD.n3493 GND 0.004551f
C5812 VDD.n3494 GND 0.004551f
C5813 VDD.n3495 GND 0.004551f
C5814 VDD.n3496 GND 0.004551f
C5815 VDD.n3497 GND 0.004551f
C5816 VDD.n3498 GND 0.004551f
C5817 VDD.n3499 GND 0.004551f
C5818 VDD.n3500 GND 0.004551f
C5819 VDD.n3501 GND 0.004551f
C5820 VDD.n3502 GND 0.004551f
C5821 VDD.n3503 GND 0.004551f
C5822 VDD.n3504 GND 0.004551f
C5823 VDD.n3505 GND 0.004551f
C5824 VDD.n3506 GND 0.004551f
C5825 VDD.n3507 GND 0.004551f
C5826 VDD.n3508 GND 0.004551f
C5827 VDD.n3509 GND 0.004551f
C5828 VDD.n3510 GND 0.004551f
C5829 VDD.n3511 GND 0.004551f
C5830 VDD.n3512 GND 0.004551f
C5831 VDD.n3513 GND 0.004551f
C5832 VDD.n3514 GND 0.004551f
C5833 VDD.n3515 GND 0.004551f
C5834 VDD.n3516 GND 0.004551f
C5835 VDD.n3517 GND 0.004551f
C5836 VDD.n3518 GND 0.004551f
C5837 VDD.n3519 GND 0.004551f
C5838 VDD.n3520 GND 0.004551f
C5839 VDD.n3521 GND 0.004551f
C5840 VDD.n3522 GND 0.004551f
C5841 VDD.n3523 GND 0.004551f
C5842 VDD.n3524 GND 0.004551f
C5843 VDD.n3525 GND 0.004551f
C5844 VDD.n3526 GND 0.004551f
C5845 VDD.n3527 GND 0.004551f
C5846 VDD.n3528 GND 0.004551f
C5847 VDD.n3529 GND 0.004551f
C5848 VDD.n3530 GND 0.004551f
C5849 VDD.n3531 GND 0.004551f
C5850 VDD.n3532 GND 0.004551f
C5851 VDD.n3533 GND 0.004551f
C5852 VDD.n3534 GND 0.004551f
C5853 VDD.n3535 GND 0.004551f
C5854 VDD.n3536 GND 0.004551f
C5855 VDD.n3537 GND 0.004551f
C5856 VDD.n3538 GND 0.004551f
C5857 VDD.n3539 GND 0.004551f
C5858 VDD.n3540 GND 0.004551f
C5859 VDD.n3541 GND 0.004551f
C5860 VDD.n3542 GND 0.004551f
C5861 VDD.n3543 GND 0.004551f
C5862 VDD.n3544 GND 0.004551f
C5863 VDD.n3545 GND 0.004551f
C5864 VDD.n3546 GND 0.004551f
C5865 VDD.n3547 GND 0.004551f
C5866 VDD.n3548 GND 0.004551f
C5867 VDD.n3549 GND 0.004551f
C5868 VDD.n3550 GND 0.004551f
C5869 VDD.n3551 GND 0.004551f
C5870 VDD.n3552 GND 0.004551f
C5871 VDD.n3553 GND 0.004551f
C5872 VDD.n3554 GND 0.004551f
C5873 VDD.n3555 GND 0.004551f
C5874 VDD.n3556 GND 0.004551f
C5875 VDD.n3557 GND 0.004551f
C5876 VDD.n3558 GND 0.004551f
C5877 VDD.n3559 GND 0.004551f
C5878 VDD.n3560 GND 0.004551f
C5879 VDD.n3561 GND 0.004551f
C5880 VDD.n3562 GND 0.004551f
C5881 VDD.n3563 GND 0.004551f
C5882 VDD.n3564 GND 0.004551f
C5883 VDD.n3565 GND 0.004551f
C5884 VDD.n3566 GND 0.004551f
C5885 VDD.n3567 GND 0.004551f
C5886 VDD.n3568 GND 0.004551f
C5887 VDD.n3569 GND 0.004551f
C5888 VDD.n3570 GND 0.004551f
C5889 VDD.n3571 GND 0.004551f
C5890 VDD.n3572 GND 0.004551f
C5891 VDD.n3573 GND 0.004551f
C5892 VDD.n3574 GND 0.004551f
C5893 VDD.n3575 GND 0.004551f
C5894 VDD.n3576 GND 0.004551f
C5895 VDD.n3577 GND 0.004551f
C5896 VDD.n3578 GND 0.004551f
C5897 VDD.n3579 GND 0.004551f
C5898 VDD.n3580 GND 0.004551f
C5899 VDD.n3581 GND 0.004551f
C5900 VDD.n3582 GND 0.004551f
C5901 VDD.n3583 GND 0.004551f
C5902 VDD.n3584 GND 0.004551f
C5903 VDD.n3585 GND 0.004551f
C5904 VDD.n3586 GND 0.004551f
C5905 VDD.n3587 GND 0.004551f
C5906 VDD.n3588 GND 0.004551f
C5907 VDD.n3589 GND 0.004551f
C5908 VDD.n3590 GND 0.004551f
C5909 VDD.n3591 GND 0.004551f
C5910 VDD.n3592 GND 0.004551f
C5911 VDD.n3593 GND 0.004551f
C5912 VDD.n3594 GND 0.004551f
C5913 VDD.n3595 GND 0.004551f
C5914 VDD.n3596 GND 0.004551f
C5915 VDD.n3597 GND 0.010814f
C5916 VDD.n3598 GND 0.010814f
C5917 VDD.n3599 GND 0.010814f
C5918 VDD.n3600 GND 0.011274f
C5919 VDD.n3601 GND 0.004551f
C5920 VDD.n3602 GND 0.004551f
C5921 VDD.n3603 GND 0.004551f
C5922 VDD.n3604 GND 0.004551f
C5923 VDD.n3605 GND 0.004551f
C5924 VDD.n3606 GND 0.004551f
C5925 VDD.n3607 GND 0.004551f
C5926 VDD.n3608 GND 0.004551f
C5927 VDD.t65 GND 0.154197f
C5928 VDD.t62 GND 0.733149f
C5929 VDD.n3609 GND 0.09739f
C5930 VDD.t64 GND 0.103896f
C5931 VDD.n3610 GND 0.100617f
C5932 VDD.n3611 GND 0.004551f
C5933 VDD.n3612 GND 0.011274f
C5934 VDD.n3613 GND 0.004551f
C5935 VDD.n3614 GND 0.004551f
C5936 VDD.n3615 GND 0.004551f
C5937 VDD.n3616 GND 0.004551f
C5938 VDD.n3617 GND 0.004551f
C5939 VDD.n3618 GND 0.004551f
C5940 VDD.n3619 GND 0.004551f
C5941 VDD.n3620 GND 0.004551f
C5942 VDD.n3621 GND 0.004551f
C5943 VDD.n3622 GND 0.004551f
C5944 VDD.n3623 GND 0.004551f
C5945 VDD.n3624 GND 0.004551f
C5946 VDD.n3625 GND 0.004551f
C5947 VDD.n3626 GND 0.004551f
C5948 VDD.n3627 GND 0.004551f
C5949 VDD.n3628 GND 0.004551f
C5950 VDD.n3629 GND 0.004551f
C5951 VDD.n3630 GND 0.004551f
C5952 VDD.n3631 GND 0.004551f
C5953 VDD.n3632 GND 0.004551f
C5954 VDD.n3633 GND 0.004551f
C5955 VDD.n3634 GND 0.004551f
C5956 VDD.n3635 GND 0.004551f
C5957 VDD.n3636 GND 0.004551f
C5958 VDD.n3637 GND 0.004551f
C5959 VDD.n3638 GND 0.004551f
C5960 VDD.n3639 GND 0.004551f
C5961 VDD.n3640 GND 0.004551f
C5962 VDD.n3641 GND 0.004551f
C5963 VDD.n3642 GND 0.004551f
C5964 VDD.n3643 GND 0.004551f
C5965 VDD.n3644 GND 0.004551f
C5966 VDD.n3645 GND 0.004551f
C5967 VDD.n3646 GND 0.004551f
C5968 VDD.n3647 GND 0.004551f
C5969 VDD.n3648 GND 0.004551f
C5970 VDD.n3649 GND 0.004551f
C5971 VDD.n3650 GND 0.004551f
C5972 VDD.n3651 GND 0.004551f
C5973 VDD.n3652 GND 0.004551f
C5974 VDD.n3653 GND 0.004551f
C5975 VDD.n3654 GND 0.004551f
C5976 VDD.n3655 GND 0.004551f
C5977 VDD.n3656 GND 0.004551f
C5978 VDD.n3657 GND 0.004551f
C5979 VDD.n3658 GND 0.004551f
C5980 VDD.n3659 GND 0.004551f
C5981 VDD.n3660 GND 0.004551f
C5982 VDD.n3661 GND 0.004551f
C5983 VDD.n3662 GND 0.004551f
C5984 VDD.n3663 GND 0.004551f
C5985 VDD.n3664 GND 0.004551f
C5986 VDD.n3665 GND 0.004551f
C5987 VDD.n3666 GND 0.004551f
C5988 VDD.n3667 GND 0.004551f
C5989 VDD.n3668 GND 0.004551f
C5990 VDD.n3669 GND 0.004551f
C5991 VDD.n3670 GND 0.004551f
C5992 VDD.n3671 GND 0.004551f
C5993 VDD.n3672 GND 0.004551f
C5994 VDD.n3673 GND 0.004551f
C5995 VDD.n3674 GND 0.004551f
C5996 VDD.n3675 GND 0.004551f
C5997 VDD.n3676 GND 0.004551f
C5998 VDD.n3677 GND 0.004551f
C5999 VDD.n3678 GND 0.004551f
C6000 VDD.n3679 GND 0.004551f
C6001 VDD.n3680 GND 0.004551f
C6002 VDD.n3681 GND 0.004551f
C6003 VDD.n3682 GND 0.004551f
C6004 VDD.n3683 GND 0.004551f
C6005 VDD.n3684 GND 0.004551f
C6006 VDD.n3685 GND 0.004551f
C6007 VDD.n3686 GND 0.004551f
C6008 VDD.n3687 GND 0.004551f
C6009 VDD.n3688 GND 0.004551f
C6010 VDD.n3689 GND 0.004551f
C6011 VDD.n3690 GND 0.004551f
C6012 VDD.n3691 GND 0.004551f
C6013 VDD.n3692 GND 0.004551f
C6014 VDD.n3693 GND 0.004551f
C6015 VDD.n3694 GND 0.004551f
C6016 VDD.n3695 GND 0.004551f
C6017 VDD.n3696 GND 0.004551f
C6018 VDD.n3697 GND 0.004551f
C6019 VDD.n3698 GND 0.004551f
C6020 VDD.n3699 GND 0.004551f
C6021 VDD.n3700 GND 0.004551f
C6022 VDD.n3701 GND 0.004551f
C6023 VDD.n3702 GND 0.004551f
C6024 VDD.n3703 GND 0.004551f
C6025 VDD.n3704 GND 0.004551f
C6026 VDD.n3705 GND 0.004551f
C6027 VDD.n3706 GND 0.004551f
C6028 VDD.n3707 GND 0.004551f
C6029 VDD.n3708 GND 0.004551f
C6030 VDD.n3709 GND 0.004551f
C6031 VDD.n3710 GND 0.004551f
C6032 VDD.n3711 GND 0.004551f
C6033 VDD.n3712 GND 0.004551f
C6034 VDD.n3713 GND 0.004551f
C6035 VDD.n3714 GND 0.004551f
C6036 VDD.n3715 GND 0.004551f
C6037 VDD.n3716 GND 0.004551f
C6038 VDD.n3717 GND 0.004551f
C6039 VDD.n3718 GND 0.004551f
C6040 VDD.n3719 GND 0.004551f
C6041 VDD.n3720 GND 0.004551f
C6042 VDD.n3721 GND 0.004551f
C6043 VDD.n3722 GND 0.004551f
C6044 VDD.n3723 GND 0.004551f
C6045 VDD.n3724 GND 0.004551f
C6046 VDD.n3725 GND 0.004551f
C6047 VDD.n3726 GND 0.004551f
C6048 VDD.n3727 GND 0.004551f
C6049 VDD.n3728 GND 0.004551f
C6050 VDD.n3729 GND 0.004551f
C6051 VDD.n3730 GND 0.004551f
C6052 VDD.n3731 GND 0.004551f
C6053 VDD.n3732 GND 0.004551f
C6054 VDD.n3733 GND 0.004551f
C6055 VDD.n3734 GND 0.004551f
C6056 VDD.n3735 GND 0.004551f
C6057 VDD.n3736 GND 0.004551f
C6058 VDD.n3737 GND 0.004551f
C6059 VDD.n3738 GND 0.004551f
C6060 VDD.n3739 GND 0.004551f
C6061 VDD.n3740 GND 0.004551f
C6062 VDD.n3741 GND 0.004551f
C6063 VDD.n3742 GND 0.004551f
C6064 VDD.n3743 GND 0.004551f
C6065 VDD.n3744 GND 0.004551f
C6066 VDD.n3745 GND 0.004551f
C6067 VDD.n3746 GND 0.004551f
C6068 VDD.n3747 GND 0.004551f
C6069 VDD.n3748 GND 0.004551f
C6070 VDD.n3749 GND 0.004551f
C6071 VDD.n3750 GND 0.004551f
C6072 VDD.n3751 GND 0.004551f
C6073 VDD.n3752 GND 0.004551f
C6074 VDD.n3753 GND 0.004551f
C6075 VDD.n3754 GND 0.004551f
C6076 VDD.n3755 GND 0.004551f
C6077 VDD.n3756 GND 0.004551f
C6078 VDD.n3757 GND 0.004551f
C6079 VDD.n3758 GND 0.004551f
C6080 VDD.n3759 GND 0.004551f
C6081 VDD.n3760 GND 0.004551f
C6082 VDD.n3761 GND 0.004551f
C6083 VDD.n3762 GND 0.004551f
C6084 VDD.n3763 GND 0.004551f
C6085 VDD.n3764 GND 0.004551f
C6086 VDD.n3765 GND 0.004551f
C6087 VDD.n3766 GND 0.004551f
C6088 VDD.n3767 GND 0.004551f
C6089 VDD.n3768 GND 0.004551f
C6090 VDD.n3769 GND 0.004551f
C6091 VDD.n3770 GND 0.004551f
C6092 VDD.n3771 GND 0.004551f
C6093 VDD.n3772 GND 0.010814f
C6094 VDD.n3773 GND 0.011274f
C6095 VDD.n3774 GND 0.004551f
C6096 VDD.n3775 GND 0.004551f
C6097 VDD.n3777 GND 0.004551f
C6098 VDD.n3779 GND 0.004551f
C6099 VDD.n3780 GND 0.00261f
C6100 VDD.n3781 GND 0.005616f
C6101 VDD.n3782 GND 0.004217f
C6102 VDD.n3783 GND 0.004551f
C6103 VDD.n3784 GND 0.004551f
C6104 VDD.n3786 GND 0.004551f
C6105 VDD.n3788 GND 0.004551f
C6106 VDD.n3789 GND 0.004551f
C6107 VDD.n3790 GND 0.004551f
C6108 VDD.n3791 GND 0.004551f
C6109 VDD.n3792 GND 0.004551f
C6110 VDD.n3794 GND 0.004551f
C6111 VDD.n3796 GND 0.004551f
C6112 VDD.n3797 GND 0.004551f
C6113 VDD.n3798 GND 0.004551f
C6114 VDD.n3799 GND 0.004551f
C6115 VDD.n3800 GND 0.004551f
C6116 VDD.n3802 GND 0.004551f
C6117 VDD.n3804 GND 0.004551f
C6118 VDD.n3805 GND 0.004551f
C6119 VDD.n3806 GND 0.004551f
C6120 VDD.n3807 GND 0.004551f
C6121 VDD.n3808 GND 0.004551f
C6122 VDD.n3810 GND 0.004551f
C6123 VDD.n3812 GND 0.004551f
C6124 VDD.n3813 GND 0.004551f
C6125 VDD.n3814 GND 0.011274f
C6126 VDD.n3815 GND 0.010814f
C6127 VDD.n3816 GND 0.010814f
C6128 VDD.n3817 GND 0.470823f
C6129 VDD.n3818 GND 0.010814f
C6130 VDD.n3819 GND 0.010814f
C6131 VDD.n3820 GND 0.004551f
C6132 VDD.n3821 GND 0.004551f
C6133 VDD.n3822 GND 0.004551f
C6134 VDD.n3823 GND 0.325035f
C6135 VDD.n3824 GND 0.004551f
C6136 VDD.n3825 GND 0.004551f
C6137 VDD.n3826 GND 0.004551f
C6138 VDD.n3827 GND 0.004551f
C6139 VDD.n3828 GND 0.004551f
C6140 VDD.n3829 GND 0.325035f
C6141 VDD.n3830 GND 0.004551f
C6142 VDD.n3831 GND 0.004551f
C6143 VDD.n3832 GND 0.004551f
C6144 VDD.n3833 GND 0.004551f
C6145 VDD.n3834 GND 0.004551f
C6146 VDD.n3835 GND 0.325035f
C6147 VDD.n3836 GND 0.004551f
C6148 VDD.n3837 GND 0.004551f
C6149 VDD.n3838 GND 0.004551f
C6150 VDD.n3839 GND 0.004551f
C6151 VDD.n3840 GND 0.004551f
C6152 VDD.n3841 GND 0.325035f
C6153 VDD.n3842 GND 0.004551f
C6154 VDD.n3843 GND 0.004551f
C6155 VDD.n3844 GND 0.004551f
C6156 VDD.n3845 GND 0.004551f
C6157 VDD.n3846 GND 0.004551f
C6158 VDD.n3847 GND 0.325035f
C6159 VDD.n3848 GND 0.004551f
C6160 VDD.n3849 GND 0.004551f
C6161 VDD.n3850 GND 0.004551f
C6162 VDD.n3851 GND 0.004551f
C6163 VDD.n3852 GND 0.004551f
C6164 VDD.n3853 GND 0.282016f
C6165 VDD.n3854 GND 0.004551f
C6166 VDD.n3855 GND 0.004551f
C6167 VDD.n3856 GND 0.004551f
C6168 VDD.n3857 GND 0.004551f
C6169 VDD.n3858 GND 0.004551f
C6170 VDD.n3859 GND 0.296356f
C6171 VDD.n3860 GND 0.004551f
C6172 VDD.n3861 GND 0.004551f
C6173 VDD.n3862 GND 0.004551f
C6174 VDD.n3863 GND 0.004551f
C6175 VDD.n3864 GND 0.004551f
C6176 VDD.n3865 GND 0.325035f
C6177 VDD.n3866 GND 0.004551f
C6178 VDD.n3867 GND 0.004551f
C6179 VDD.n3868 GND 0.004551f
C6180 VDD.n3869 GND 0.004551f
C6181 VDD.n3870 GND 0.004551f
C6182 VDD.n3871 GND 0.325035f
C6183 VDD.n3872 GND 0.004551f
C6184 VDD.n3873 GND 0.004551f
C6185 VDD.n3874 GND 0.004551f
C6186 VDD.n3875 GND 0.004551f
C6187 VDD.n3876 GND 0.004551f
C6188 VDD.n3877 GND 0.325035f
C6189 VDD.n3878 GND 0.004551f
C6190 VDD.n3879 GND 0.004551f
C6191 VDD.n3880 GND 0.004551f
C6192 VDD.n3881 GND 0.004551f
C6193 VDD.n3882 GND 0.004551f
C6194 VDD.n3883 GND 0.325035f
C6195 VDD.n3884 GND 0.004551f
C6196 VDD.n3885 GND 0.004551f
C6197 VDD.n3886 GND 0.004551f
C6198 VDD.n3887 GND 0.004551f
C6199 VDD.n3888 GND 0.004551f
C6200 VDD.n3889 GND 0.325035f
C6201 VDD.n3890 GND 0.004551f
C6202 VDD.n3891 GND 0.004551f
C6203 VDD.n3892 GND 0.004551f
C6204 VDD.n3893 GND 0.004551f
C6205 VDD.n3894 GND 0.004551f
C6206 VDD.n3895 GND 0.325035f
C6207 VDD.n3896 GND 0.004551f
C6208 VDD.n3897 GND 0.004551f
C6209 VDD.n3898 GND 0.004551f
C6210 VDD.n3899 GND 0.004551f
C6211 VDD.n3900 GND 0.004551f
C6212 VDD.n3901 GND 0.325035f
C6213 VDD.n3902 GND 0.004551f
C6214 VDD.n3903 GND 0.004551f
C6215 VDD.n3904 GND 0.004551f
C6216 VDD.n3905 GND 0.004551f
C6217 VDD.n3906 GND 0.004551f
C6218 VDD.n3907 GND 0.325035f
C6219 VDD.n3908 GND 0.004551f
C6220 VDD.n3909 GND 0.004551f
C6221 VDD.n3910 GND 0.004551f
C6222 VDD.n3911 GND 0.004551f
C6223 VDD.n3912 GND 0.004551f
C6224 VDD.n3913 GND 0.277236f
C6225 VDD.n3914 GND 0.004551f
C6226 VDD.n3915 GND 0.004551f
C6227 VDD.n3916 GND 0.004551f
C6228 VDD.n3917 GND 0.004551f
C6229 VDD.n3918 GND 0.004551f
C6230 VDD.n3919 GND 0.320255f
C6231 VDD.n3920 GND 0.004551f
C6232 VDD.n3921 GND 0.004551f
C6233 VDD.n3922 GND 0.004551f
C6234 VDD.n3923 GND 0.004551f
C6235 VDD.n3924 GND 0.004551f
C6236 VDD.n3925 GND 0.325035f
C6237 VDD.n3926 GND 0.004551f
C6238 VDD.n3927 GND 0.004551f
C6239 VDD.n3928 GND 0.004551f
C6240 VDD.n3929 GND 0.004551f
C6241 VDD.n3930 GND 0.004551f
C6242 VDD.n3931 GND 0.325035f
C6243 VDD.n3932 GND 0.004551f
C6244 VDD.n3933 GND 0.004551f
C6245 VDD.n3934 GND 0.004551f
C6246 VDD.n3935 GND 0.004551f
C6247 VDD.n3936 GND 0.004551f
C6248 VDD.n3937 GND 0.325035f
C6249 VDD.n3938 GND 0.004551f
C6250 VDD.n3939 GND 0.004551f
C6251 VDD.n3940 GND 0.004551f
C6252 VDD.n3941 GND 0.004551f
C6253 VDD.n3942 GND 0.004551f
C6254 VDD.n3943 GND 0.325035f
C6255 VDD.n3944 GND 0.004551f
C6256 VDD.n3945 GND 0.004551f
C6257 VDD.n3946 GND 0.004551f
C6258 VDD.n3947 GND 0.004551f
C6259 VDD.n3948 GND 0.004551f
C6260 VDD.n3949 GND 0.325035f
C6261 VDD.n3950 GND 0.004551f
C6262 VDD.n3951 GND 0.004551f
C6263 VDD.n3952 GND 0.004551f
C6264 VDD.n3953 GND 0.004551f
C6265 VDD.n3954 GND 0.004551f
C6266 VDD.n3955 GND 0.325035f
C6267 VDD.n3956 GND 0.004551f
C6268 VDD.n3957 GND 0.004551f
C6269 VDD.n3958 GND 0.004551f
C6270 VDD.n3959 GND 0.004551f
C6271 VDD.n3960 GND 0.004551f
C6272 VDD.n3961 GND 0.325035f
C6273 VDD.n3962 GND 0.004551f
C6274 VDD.n3963 GND 0.004551f
C6275 VDD.n3964 GND 0.004551f
C6276 VDD.n3965 GND 0.004551f
C6277 VDD.n3966 GND 0.004551f
C6278 VDD.n3967 GND 0.325035f
C6279 VDD.n3968 GND 0.004551f
C6280 VDD.n3969 GND 0.004551f
C6281 VDD.n3970 GND 0.004551f
C6282 VDD.n3971 GND 0.004551f
C6283 VDD.n3972 GND 0.004551f
C6284 VDD.n3973 GND 0.200757f
C6285 VDD.n3974 GND 0.004551f
C6286 VDD.n3975 GND 0.004551f
C6287 VDD.n3976 GND 0.004551f
C6288 VDD.n3977 GND 0.004551f
C6289 VDD.n3978 GND 0.004551f
C6290 VDD.n3979 GND 0.243776f
C6291 VDD.n3980 GND 0.004551f
C6292 VDD.n3981 GND 0.004551f
C6293 VDD.n3982 GND 0.004551f
C6294 VDD.n3983 GND 0.004551f
C6295 VDD.n3984 GND 0.004551f
C6296 VDD.n3985 GND 0.325035f
C6297 VDD.n3986 GND 0.004551f
C6298 VDD.n3987 GND 0.004551f
C6299 VDD.n3988 GND 0.004551f
C6300 VDD.n3989 GND 0.004551f
C6301 VDD.n3990 GND 0.004551f
C6302 VDD.n3991 GND 0.325035f
C6303 VDD.n3992 GND 0.004551f
C6304 VDD.n3993 GND 0.004551f
C6305 VDD.n3994 GND 0.004551f
C6306 VDD.n3995 GND 0.004551f
C6307 VDD.n3996 GND 0.004551f
C6308 VDD.n3997 GND 0.325035f
C6309 VDD.n3998 GND 0.004551f
C6310 VDD.n3999 GND 0.004551f
C6311 VDD.n4000 GND 0.004551f
C6312 VDD.n4001 GND 0.004551f
C6313 VDD.n4002 GND 0.004551f
C6314 VDD.n4003 GND 0.325035f
C6315 VDD.n4004 GND 0.004551f
C6316 VDD.n4005 GND 0.004551f
C6317 VDD.n4006 GND 0.004551f
C6318 VDD.n4007 GND 0.004551f
C6319 VDD.n4008 GND 0.004551f
C6320 VDD.n4009 GND 0.325035f
C6321 VDD.n4010 GND 0.004551f
C6322 VDD.n4011 GND 0.004551f
C6323 VDD.n4012 GND 0.004551f
C6324 VDD.n4013 GND 0.004551f
C6325 VDD.n4014 GND 0.004551f
C6326 VDD.n4015 GND 0.325035f
C6327 VDD.n4016 GND 0.004551f
C6328 VDD.n4017 GND 0.004551f
C6329 VDD.n4018 GND 0.004551f
C6330 VDD.n4019 GND 0.004551f
C6331 VDD.n4020 GND 0.004551f
C6332 VDD.n4021 GND 0.325035f
C6333 VDD.n4022 GND 0.004551f
C6334 VDD.n4023 GND 0.004551f
C6335 VDD.n4024 GND 0.004551f
C6336 VDD.n4025 GND 0.004551f
C6337 VDD.n4026 GND 0.004551f
C6338 VDD.n4027 GND 0.325035f
C6339 VDD.n4028 GND 0.004551f
C6340 VDD.n4029 GND 0.004551f
C6341 VDD.n4030 GND 0.004551f
C6342 VDD.n4031 GND 0.004551f
C6343 VDD.n4032 GND 0.004551f
C6344 VDD.n4033 GND 0.200757f
C6345 VDD.n4034 GND 0.004551f
C6346 VDD.n4035 GND 0.004551f
C6347 VDD.n4036 GND 0.004551f
C6348 VDD.n4037 GND 0.004551f
C6349 VDD.n4038 GND 0.004551f
C6350 VDD.n4039 GND 0.167298f
C6351 VDD.n4040 GND 0.004551f
C6352 VDD.n4041 GND 0.004551f
C6353 VDD.n4042 GND 0.004551f
C6354 VDD.n4043 GND 0.004551f
C6355 VDD.n4044 GND 0.004551f
C6356 VDD.n4045 GND 0.325035f
C6357 VDD.n4046 GND 0.004551f
C6358 VDD.n4047 GND 0.004551f
C6359 VDD.n4048 GND 0.004551f
C6360 VDD.n4049 GND 0.004551f
C6361 VDD.n4050 GND 0.004551f
C6362 VDD.n4051 GND 0.325035f
C6363 VDD.n4052 GND 0.004551f
C6364 VDD.n4053 GND 0.004551f
C6365 VDD.n4054 GND 0.004551f
C6366 VDD.n4055 GND 0.004551f
C6367 VDD.n4056 GND 0.004551f
C6368 VDD.n4057 GND 0.325035f
C6369 VDD.n4058 GND 0.004551f
C6370 VDD.n4059 GND 0.004551f
C6371 VDD.n4060 GND 0.004551f
C6372 VDD.n4061 GND 0.004551f
C6373 VDD.n4062 GND 0.004551f
C6374 VDD.n4063 GND 0.325035f
C6375 VDD.n4064 GND 0.004551f
C6376 VDD.n4065 GND 0.004551f
C6377 VDD.n4066 GND 0.004551f
C6378 VDD.n4067 GND 0.004551f
C6379 VDD.n4068 GND 0.004551f
C6380 VDD.n4069 GND 0.325035f
C6381 VDD.n4070 GND 0.004551f
C6382 VDD.n4071 GND 0.004551f
C6383 VDD.n4072 GND 0.004551f
C6384 VDD.n4073 GND 0.004551f
C6385 VDD.n4074 GND 0.004551f
C6386 VDD.n4075 GND 0.325035f
C6387 VDD.n4076 GND 0.004551f
C6388 VDD.n4077 GND 0.004551f
C6389 VDD.n4078 GND 0.004551f
C6390 VDD.n4079 GND 0.004551f
C6391 VDD.n4080 GND 0.004551f
C6392 VDD.n4081 GND 0.325035f
C6393 VDD.n4082 GND 0.004551f
C6394 VDD.n4083 GND 0.004551f
C6395 VDD.n4084 GND 0.004551f
C6396 VDD.n4085 GND 0.004551f
C6397 VDD.n4086 GND 0.004551f
C6398 VDD.n4087 GND 0.325035f
C6399 VDD.n4088 GND 0.004551f
C6400 VDD.n4089 GND 0.004551f
C6401 VDD.n4090 GND 0.004551f
C6402 VDD.n4091 GND 0.004551f
C6403 VDD.n4092 GND 0.004551f
C6404 VDD.n4093 GND 0.325035f
C6405 VDD.n4094 GND 0.004551f
C6406 VDD.n4095 GND 0.004551f
C6407 VDD.n4096 GND 0.004551f
C6408 VDD.n4097 GND 0.004551f
C6409 VDD.n4098 GND 0.004551f
C6410 VDD.n4099 GND 0.325035f
C6411 VDD.n4100 GND 0.004551f
C6412 VDD.n4101 GND 0.004551f
C6413 VDD.n4102 GND 0.004551f
C6414 VDD.n4103 GND 0.004551f
C6415 VDD.n4104 GND 0.004551f
C6416 VDD.n4105 GND 0.325035f
C6417 VDD.n4106 GND 0.004551f
C6418 VDD.n4107 GND 0.004551f
C6419 VDD.n4108 GND 0.004551f
C6420 VDD.n4109 GND 0.004551f
C6421 VDD.n4110 GND 0.004551f
C6422 VDD.n4111 GND 0.205537f
C6423 VDD.n4112 GND 0.004551f
C6424 VDD.n4113 GND 0.004551f
C6425 VDD.n4114 GND 0.004551f
C6426 VDD.n4115 GND 0.004551f
C6427 VDD.n4116 GND 0.004551f
C6428 VDD.n4117 GND 0.277236f
C6429 VDD.n4118 GND 0.004551f
C6430 VDD.n4119 GND 0.004551f
C6431 VDD.n4120 GND 0.004551f
C6432 VDD.n4121 GND 0.004551f
C6433 VDD.n4122 GND 0.004551f
C6434 VDD.n4123 GND 0.325035f
C6435 VDD.n4124 GND 0.004551f
C6436 VDD.n4125 GND 0.004551f
C6437 VDD.n4126 GND 0.004551f
C6438 VDD.n4127 GND 0.011274f
C6439 VDD.n4128 GND 0.004551f
C6440 VDD.n4129 GND 0.004551f
C6441 VDD.n4130 GND 0.004551f
C6442 VDD.n4132 GND 0.004551f
C6443 VDD.n4134 GND 0.004551f
C6444 VDD.n4135 GND 0.004551f
C6445 VDD.n4136 GND 0.004551f
C6446 VDD.n4137 GND 0.004551f
C6447 VDD.n4138 GND 0.004551f
C6448 VDD.n4139 GND 0.004551f
C6449 VDD.n4141 GND 0.004551f
C6450 VDD.n4142 GND 0.004551f
C6451 VDD.n4143 GND 0.004551f
C6452 VDD.n4144 GND 0.004551f
C6453 VDD.n4145 GND 0.004551f
C6454 VDD.n4146 GND 0.004551f
C6455 VDD.n4148 GND 0.004551f
C6456 VDD.n4149 GND 0.011274f
C6457 VDD.n4150 GND 0.010814f
C6458 VDD.n4151 GND 0.010814f
C6459 VDD.n4152 GND 0.004551f
C6460 VDD.n4153 GND 0.004551f
C6461 VDD.n4154 GND 0.004551f
C6462 VDD.n4155 GND 0.004551f
C6463 VDD.n4156 GND 0.004551f
C6464 VDD.n4157 GND 0.004551f
C6465 VDD.n4158 GND 0.004551f
C6466 VDD.n4159 GND 0.325035f
C6467 VDD.n4160 GND 0.004551f
C6468 VDD.n4161 GND 0.004551f
C6469 VDD.n4162 GND 0.004551f
C6470 VDD.n4163 GND 0.004551f
C6471 VDD.n4164 GND 0.004551f
C6472 VDD.n4165 GND 0.325035f
C6473 VDD.n4166 GND 0.004551f
C6474 VDD.n4167 GND 0.004551f
C6475 VDD.n4168 GND 0.004551f
C6476 VDD.n4169 GND 0.004551f
C6477 VDD.n4170 GND 0.011323f
C6478 VDD.n4172 GND 0.010814f
C6479 VDD.n4173 GND 0.011274f
C6480 VDD.n4174 GND 0.010764f
C6481 VDD.n4175 GND 0.004551f
C6482 VDD.n4176 GND 0.004551f
C6483 VDD.n4177 GND 0.004551f
C6484 VDD.n4179 GND 0.004551f
C6485 VDD.n4180 GND 0.004551f
C6486 VDD.n4181 GND 0.004217f
C6487 VDD.n4182 GND 0.004551f
C6488 VDD.n4183 GND 0.004551f
C6489 VDD.n4184 GND 0.004551f
C6490 VDD.n4186 GND 0.004551f
C6491 VDD.n4187 GND 0.004551f
C6492 VDD.n4188 GND 0.004551f
C6493 VDD.n4189 GND 0.004551f
C6494 VDD.n4190 GND 0.18734f
C6495 VDD.n4191 GND 0.004551f
C6496 VDD.n4193 GND 0.004551f
C6497 VDD.n4194 GND 0.004551f
C6498 VDD.n4195 GND 0.004551f
C6499 VDD.n4196 GND 0.004551f
C6500 VDD.n4197 GND 0.004551f
C6501 VDD.n4198 GND 0.004551f
C6502 VDD.n4200 GND 0.004551f
C6503 VDD.n4201 GND 0.004551f
C6504 VDD.n4202 GND 0.004551f
C6505 VDD.n4203 GND 0.004551f
C6506 VDD.n4204 GND 0.004551f
C6507 VDD.n4205 GND 0.004551f
C6508 VDD.n4207 GND 0.004551f
C6509 VDD.n4208 GND 0.011274f
C6510 VDD.n4209 GND 0.011274f
C6511 VDD.n4210 GND 0.010814f
C6512 VDD.n4211 GND 0.004551f
C6513 VDD.n4212 GND 0.004551f
C6514 VDD.n4213 GND 0.325035f
C6515 VDD.n4214 GND 0.004551f
C6516 VDD.n4215 GND 0.004551f
C6517 VDD.n4216 GND 0.011323f
C6518 VDD.n4217 GND 0.010764f
C6519 VDD.n4218 GND 0.011274f
C6520 VDD.n4220 GND 0.004551f
C6521 VDD.n4221 GND 0.004551f
C6522 VDD.n4222 GND 0.004551f
C6523 VDD.n4223 GND 0.00261f
C6524 VDD.n4224 GND 0.005616f
C6525 VDD.n4225 GND 0.004217f
C6526 VDD.n4226 GND 0.004551f
C6527 VDD.n4228 GND 0.004551f
C6528 VDD.n4229 GND 0.004551f
C6529 VDD.n4230 GND 0.004551f
C6530 VDD.n4231 GND 0.004551f
C6531 VDD.n4232 GND 0.004551f
C6532 VDD.n4233 GND 0.004551f
C6533 VDD.n4235 GND 0.004551f
C6534 VDD.n4236 GND 0.004551f
C6535 VDD.n4237 GND 0.18734f
C6536 VDD.n4238 GND 1.90429f
C6537 VDD.n4239 GND 0.043283f
C6538 VDD.n4240 GND 0.002667f
C6539 VDD.n4241 GND 0.016349f
C6540 VDD.n4242 GND 4.14181f
C6541 VDD.n4244 GND 0.006693f
C6542 VDD.n4245 GND 0.005387f
C6543 VDD.n4246 GND 0.004471f
C6544 VDD.n4247 GND 0.04079f
C6545 VDD.n4248 GND 0.01341f
C6546 VDD.n4249 GND 0.006693f
C6547 VDD.n4250 GND 0.005387f
C6548 VDD.n4251 GND 0.006693f
C6549 VDD.n4252 GND 0.477993f
C6550 VDD.n4253 GND 0.006693f
C6551 VDD.n4254 GND 0.005387f
C6552 VDD.n4255 GND 0.006693f
C6553 VDD.n4256 GND 0.006693f
C6554 VDD.n4257 GND 0.006693f
C6555 VDD.n4258 GND 0.005387f
C6556 VDD.n4259 GND 0.006693f
C6557 VDD.n4260 GND 0.477993f
C6558 VDD.n4261 GND 0.006693f
C6559 VDD.n4262 GND 0.005387f
C6560 VDD.n4263 GND 0.006693f
C6561 VDD.n4264 GND 0.006693f
C6562 VDD.n4265 GND 0.006693f
C6563 VDD.n4266 GND 0.005387f
C6564 VDD.n4267 GND 0.006693f
C6565 VDD.n4268 GND 0.477993f
C6566 VDD.n4269 GND 0.006693f
C6567 VDD.n4270 GND 0.005387f
C6568 VDD.n4271 GND 0.006693f
C6569 VDD.n4272 GND 0.006693f
C6570 VDD.n4273 GND 0.006693f
C6571 VDD.n4274 GND 0.005387f
C6572 VDD.n4275 GND 0.006693f
C6573 VDD.n4276 GND 0.368055f
C6574 VDD.n4277 GND 0.006693f
C6575 VDD.n4278 GND 0.005387f
C6576 VDD.n4279 GND 0.006693f
C6577 VDD.n4280 GND 0.006693f
C6578 VDD.n4281 GND 0.006693f
C6579 VDD.n4282 GND 0.005387f
C6580 VDD.n4283 GND 0.006693f
C6581 VDD.n4284 GND 0.477993f
C6582 VDD.n4285 GND 0.006693f
C6583 VDD.n4286 GND 0.005387f
C6584 VDD.n4287 GND 0.006693f
C6585 VDD.n4288 GND 0.006693f
C6586 VDD.n4289 GND 0.006693f
C6587 VDD.n4290 GND 0.005387f
C6588 VDD.n4291 GND 0.006693f
C6589 VDD.n4292 GND 0.477993f
C6590 VDD.n4293 GND 0.006693f
C6591 VDD.n4294 GND 0.005387f
C6592 VDD.n4295 GND 0.006693f
C6593 VDD.n4296 GND 0.006693f
C6594 VDD.n4297 GND 0.006693f
C6595 VDD.n4298 GND 0.005387f
C6596 VDD.n4299 GND 0.006693f
C6597 VDD.n4300 GND 0.477993f
C6598 VDD.n4301 GND 0.006693f
C6599 VDD.n4302 GND 0.005387f
C6600 VDD.n4303 GND 0.006693f
C6601 VDD.n4304 GND 0.006693f
C6602 VDD.n4305 GND 0.006693f
C6603 VDD.n4306 GND 0.005387f
C6604 VDD.n4307 GND 0.006693f
C6605 VDD.n4308 GND 0.477993f
C6606 VDD.n4309 GND 0.006693f
C6607 VDD.n4310 GND 0.005387f
C6608 VDD.n4311 GND 0.006693f
C6609 VDD.n4312 GND 0.006693f
C6610 VDD.n4313 GND 0.006693f
C6611 VDD.n4314 GND 0.005387f
C6612 VDD.n4315 GND 0.006693f
C6613 VDD.n4316 GND 0.477993f
C6614 VDD.n4317 GND 0.006693f
C6615 VDD.n4318 GND 0.005387f
C6616 VDD.n4319 GND 0.006693f
C6617 VDD.n4320 GND 0.006693f
C6618 VDD.n4321 GND 0.006693f
C6619 VDD.n4322 GND 0.005387f
C6620 VDD.n4323 GND 0.006693f
C6621 VDD.n4324 GND 0.477993f
C6622 VDD.n4325 GND 0.006693f
C6623 VDD.n4326 GND 0.005387f
C6624 VDD.n4327 GND 0.006693f
C6625 VDD.n4328 GND 0.006693f
C6626 VDD.n4329 GND 0.006693f
C6627 VDD.n4330 GND 0.005387f
C6628 VDD.n4331 GND 0.006693f
C6629 VDD.n4332 GND 0.382394f
C6630 VDD.n4333 GND 0.006693f
C6631 VDD.n4334 GND 0.005387f
C6632 VDD.n4335 GND 0.006693f
C6633 VDD.n4336 GND 0.006693f
C6634 VDD.n4337 GND 0.006693f
C6635 VDD.n4338 GND 0.005387f
C6636 VDD.n4339 GND 0.006693f
C6637 VDD.n4340 GND 0.477993f
C6638 VDD.n4341 GND 0.006693f
C6639 VDD.n4342 GND 0.005387f
C6640 VDD.n4343 GND 0.006693f
C6641 VDD.n4344 GND 0.006693f
C6642 VDD.n4345 GND 0.006693f
C6643 VDD.n4346 GND 0.005387f
C6644 VDD.n4347 GND 0.006693f
C6645 VDD.n4348 GND 0.477993f
C6646 VDD.n4349 GND 0.006693f
C6647 VDD.n4350 GND 0.005387f
C6648 VDD.n4351 GND 0.006693f
C6649 VDD.n4352 GND 0.006693f
C6650 VDD.n4353 GND 0.006693f
C6651 VDD.n4354 GND 0.005387f
C6652 VDD.n4355 GND 0.006693f
C6653 VDD.n4356 GND 0.477993f
C6654 VDD.n4357 GND 0.006693f
C6655 VDD.n4358 GND 0.005387f
C6656 VDD.n4359 GND 0.006693f
C6657 VDD.n4360 GND 0.006693f
C6658 VDD.n4361 GND 0.006693f
C6659 VDD.n4362 GND 0.005387f
C6660 VDD.n4363 GND 0.006693f
C6661 VDD.n4364 GND 0.477993f
C6662 VDD.n4365 GND 0.006693f
C6663 VDD.n4366 GND 0.005387f
C6664 VDD.n4367 GND 0.006693f
C6665 VDD.n4368 GND 0.006693f
C6666 VDD.n4369 GND 0.006693f
C6667 VDD.n4370 GND 0.005387f
C6668 VDD.n4371 GND 0.006693f
C6669 VDD.n4372 GND 0.477993f
C6670 VDD.n4373 GND 0.006693f
C6671 VDD.n4374 GND 0.005387f
C6672 VDD.n4375 GND 0.006693f
C6673 VDD.n4376 GND 0.006693f
C6674 VDD.n4377 GND 0.006693f
C6675 VDD.n4378 GND 0.005387f
C6676 VDD.n4379 GND 0.006693f
C6677 VDD.n4380 GND 0.454093f
C6678 VDD.n4381 GND 0.006693f
C6679 VDD.n4382 GND 0.005387f
C6680 VDD.n4383 GND 0.006693f
C6681 VDD.n4384 GND 0.006693f
C6682 VDD.n4385 GND 0.006693f
C6683 VDD.n4386 GND 0.005387f
C6684 VDD.n4387 GND 0.006693f
C6685 VDD.n4388 GND 0.477993f
C6686 VDD.n4389 GND 0.006693f
C6687 VDD.n4390 GND 0.005387f
C6688 VDD.n4391 GND 0.006693f
C6689 VDD.n4392 GND 0.006693f
C6690 VDD.n4393 GND 0.006693f
C6691 VDD.n4394 GND 0.005387f
C6692 VDD.n4395 GND 0.006693f
C6693 VDD.n4396 GND 0.477993f
C6694 VDD.n4397 GND 0.006693f
C6695 VDD.n4398 GND 0.005387f
C6696 VDD.n4399 GND 0.006693f
C6697 VDD.n4400 GND 0.006693f
C6698 VDD.n4401 GND 0.006693f
C6699 VDD.n4402 GND 0.005387f
C6700 VDD.n4403 GND 0.006693f
C6701 VDD.n4404 GND 0.477993f
C6702 VDD.n4405 GND 0.006693f
C6703 VDD.n4406 GND 0.005387f
C6704 VDD.n4407 GND 0.006693f
C6705 VDD.n4408 GND 0.006693f
C6706 VDD.n4409 GND 0.006693f
C6707 VDD.n4410 GND 0.005387f
C6708 VDD.n4411 GND 0.006693f
C6709 VDD.n4412 GND 0.477993f
C6710 VDD.n4413 GND 0.006693f
C6711 VDD.n4414 GND 0.005387f
C6712 VDD.n4415 GND 0.006693f
C6713 VDD.n4416 GND 0.006693f
C6714 VDD.n4417 GND 0.006693f
C6715 VDD.n4418 GND 0.005387f
C6716 VDD.n4419 GND 0.006693f
C6717 VDD.n4420 GND 0.477993f
C6718 VDD.n4421 GND 0.006693f
C6719 VDD.n4422 GND 0.005387f
C6720 VDD.n4423 GND 0.006693f
C6721 VDD.n4424 GND 0.006693f
C6722 VDD.n4425 GND 0.006693f
C6723 VDD.n4426 GND 0.005387f
C6724 VDD.n4427 GND 0.006693f
C6725 VDD.n4428 GND 0.477993f
C6726 VDD.n4429 GND 0.006693f
C6727 VDD.n4430 GND 0.005387f
C6728 VDD.n4431 GND 0.006693f
C6729 VDD.n4432 GND 0.006693f
C6730 VDD.n4433 GND 0.006693f
C6731 VDD.n4434 GND 0.005387f
C6732 VDD.n4435 GND 0.006693f
C6733 VDD.n4436 GND 0.430194f
C6734 VDD.n4437 GND 0.006693f
C6735 VDD.n4438 GND 0.005387f
C6736 VDD.n4439 GND 0.006693f
C6737 VDD.n4440 GND 0.006693f
C6738 VDD.n4441 GND 0.006693f
C6739 VDD.n4442 GND 0.005387f
C6740 VDD.n4443 GND 0.006693f
C6741 VDD.n4444 GND 0.477993f
C6742 VDD.n4445 GND 0.006693f
C6743 VDD.n4446 GND 0.005387f
C6744 VDD.n4447 GND 0.006693f
C6745 VDD.n4448 GND 0.006693f
C6746 VDD.n4449 GND 0.006693f
C6747 VDD.n4450 GND 0.006693f
C6748 VDD.n4451 GND 0.005387f
C6749 VDD.n4452 GND 0.005387f
C6750 VDD.n4453 GND 0.006693f
C6751 VDD.n4454 GND 0.477993f
C6752 VDD.n4455 GND 0.006693f
C6753 VDD.n4456 GND 0.005387f
C6754 VDD.n4457 GND 0.006693f
C6755 VDD.n4458 GND 0.006693f
C6756 VDD.n4459 GND 0.006693f
C6757 VDD.n4460 GND 0.005387f
C6758 VDD.n4461 GND 0.006693f
C6759 VDD.n4462 GND 0.477993f
C6760 VDD.n4463 GND 0.006693f
C6761 VDD.n4464 GND 0.006693f
C6762 VDD.n4465 GND 0.005387f
C6763 VDD.n4466 GND 0.006693f
C6764 VDD.n4467 GND 0.006693f
C6765 VDD.n4468 GND 0.006693f
C6766 VDD.n4469 GND 0.006693f
C6767 VDD.n4470 GND 0.006693f
C6768 VDD.n4471 GND 0.005387f
C6769 VDD.n4472 GND 0.005387f
C6770 VDD.n4473 GND 0.006693f
C6771 VDD.n4474 GND 0.477993f
C6772 VDD.n4475 GND 0.477993f
C6773 VDD.n4476 GND 0.006693f
C6774 VDD.n4477 GND 0.005387f
C6775 VDD.n4478 GND 0.006693f
C6776 VDD.n4479 GND 0.006693f
C6777 VDD.n4480 GND 0.006693f
C6778 VDD.n4481 GND 0.005387f
C6779 VDD.n4482 GND 0.006693f
C6780 VDD.n4483 GND 0.006693f
C6781 VDD.n4484 GND 0.358495f
C6782 VDD.n4485 GND 0.006693f
C6783 VDD.n4486 GND 0.006693f
C6784 VDD.n4487 GND 0.005387f
C6785 VDD.n4488 GND 0.005387f
C6786 VDD.n4489 GND 0.005387f
C6787 VDD.n4490 GND 0.006693f
C6788 VDD.n4491 GND 0.006693f
C6789 VDD.n4492 GND 0.006693f
C6790 VDD.n4493 GND 0.006693f
C6791 VDD.n4494 GND 0.005387f
C6792 VDD.n4495 GND 0.005387f
C6793 VDD.n4496 GND 0.005387f
C6794 VDD.n4497 GND 0.006693f
C6795 VDD.n4498 GND 0.006693f
C6796 VDD.n4499 GND 0.006693f
C6797 VDD.n4500 GND 0.006693f
C6798 VDD.n4501 GND 0.005387f
C6799 VDD.n4502 GND 0.005387f
C6800 VDD.n4503 GND 0.005387f
C6801 VDD.n4504 GND 0.006693f
C6802 VDD.n4505 GND 0.006693f
C6803 VDD.n4506 GND 0.006693f
C6804 VDD.n4507 GND 0.006693f
C6805 VDD.n4508 GND 0.005387f
C6806 VDD.n4509 GND 0.005387f
C6807 VDD.n4510 GND 0.005387f
C6808 VDD.n4511 GND 0.006693f
C6809 VDD.n4512 GND 0.006693f
C6810 VDD.n4513 GND 0.006693f
C6811 VDD.n4514 GND 0.006693f
C6812 VDD.n4515 GND 0.005387f
C6813 VDD.n4516 GND 0.005387f
C6814 VDD.n4517 GND 0.005387f
C6815 VDD.n4518 GND 0.006693f
C6816 VDD.n4519 GND 0.006693f
C6817 VDD.n4520 GND 0.006693f
C6818 VDD.n4521 GND 0.006693f
C6819 VDD.n4522 GND 0.005387f
C6820 VDD.n4523 GND 0.005387f
C6821 VDD.n4524 GND 0.005387f
C6822 VDD.n4525 GND 0.006693f
C6823 VDD.n4526 GND 0.006693f
C6824 VDD.n4527 GND 0.006693f
C6825 VDD.n4528 GND 0.006693f
C6826 VDD.n4529 GND 0.005387f
C6827 VDD.n4530 GND 0.005387f
C6828 VDD.n4531 GND 0.005387f
C6829 VDD.n4532 GND 0.006693f
C6830 VDD.n4533 GND 0.006693f
C6831 VDD.n4534 GND 0.006693f
C6832 VDD.n4535 GND 0.006693f
C6833 VDD.n4536 GND 0.005387f
C6834 VDD.n4537 GND 0.005387f
C6835 VDD.n4538 GND 0.005387f
C6836 VDD.n4539 GND 0.006693f
C6837 VDD.n4540 GND 0.006693f
C6838 VDD.n4541 GND 0.006693f
C6839 VDD.n4542 GND 0.006693f
C6840 VDD.n4543 GND 0.005387f
C6841 VDD.n4544 GND 0.005387f
C6842 VDD.n4545 GND 0.005387f
C6843 VDD.n4546 GND 0.006693f
C6844 VDD.n4547 GND 0.006693f
C6845 VDD.n4548 GND 0.006693f
C6846 VDD.n4549 GND 0.006693f
C6847 VDD.n4550 GND 0.005387f
C6848 VDD.n4551 GND 0.005387f
C6849 VDD.n4552 GND 0.005387f
C6850 VDD.n4553 GND 0.006693f
C6851 VDD.n4554 GND 0.006693f
C6852 VDD.n4555 GND 0.006693f
C6853 VDD.n4556 GND 0.006693f
C6854 VDD.n4557 GND 0.005387f
C6855 VDD.n4558 GND 0.005387f
C6856 VDD.n4559 GND 0.005387f
C6857 VDD.n4560 GND 0.006693f
C6858 VDD.n4561 GND 0.006693f
C6859 VDD.n4562 GND 0.006693f
C6860 VDD.n4563 GND 0.006693f
C6861 VDD.n4564 GND 0.005387f
C6862 VDD.n4565 GND 0.005387f
C6863 VDD.n4566 GND 0.005387f
C6864 VDD.n4567 GND 0.006693f
C6865 VDD.n4568 GND 0.006693f
C6866 VDD.n4569 GND 0.006693f
C6867 VDD.n4570 GND 0.006693f
C6868 VDD.n4571 GND 0.005387f
C6869 VDD.n4572 GND 0.005387f
C6870 VDD.n4573 GND 0.005387f
C6871 VDD.n4574 GND 0.006693f
C6872 VDD.n4575 GND 0.006693f
C6873 VDD.n4576 GND 0.006693f
C6874 VDD.n4577 GND 0.006693f
C6875 VDD.n4578 GND 0.005387f
C6876 VDD.n4579 GND 0.005387f
C6877 VDD.n4580 GND 0.005387f
C6878 VDD.n4581 GND 0.006693f
C6879 VDD.n4582 GND 0.006693f
C6880 VDD.n4583 GND 0.006693f
C6881 VDD.n4584 GND 0.006693f
C6882 VDD.n4585 GND 0.005387f
C6883 VDD.n4586 GND 0.005387f
C6884 VDD.n4587 GND 0.004471f
C6885 VDD.n4588 GND 0.01598f
C6886 VDD.n4589 GND 0.016349f
C6887 VDD.n4590 GND 0.002667f
C6888 VDD.n4591 GND 0.016349f
C6889 VDD.n4593 GND 1.13762f
C6890 VDD.n4594 GND 0.70265f
C6891 VDD.n4595 GND 0.477993f
C6892 VDD.n4596 GND 0.006693f
C6893 VDD.n4597 GND 0.005387f
C6894 VDD.n4598 GND 0.005387f
C6895 VDD.n4599 GND 0.005387f
C6896 VDD.n4600 GND 0.006693f
C6897 VDD.n4601 GND 0.477993f
C6898 VDD.n4602 GND 0.477993f
C6899 VDD.n4603 GND 0.477993f
C6900 VDD.n4604 GND 0.006693f
C6901 VDD.n4605 GND 0.005387f
C6902 VDD.n4606 GND 0.005387f
C6903 VDD.n4607 GND 0.005387f
C6904 VDD.n4608 GND 0.006693f
C6905 VDD.n4609 GND 0.368055f
C6906 VDD.n4610 GND 0.477993f
C6907 VDD.n4611 GND 0.477993f
C6908 VDD.n4612 GND 0.006693f
C6909 VDD.n4613 GND 0.005387f
C6910 VDD.n4614 GND 0.005387f
C6911 VDD.n4615 GND 0.005387f
C6912 VDD.n4616 GND 0.006693f
C6913 VDD.n4617 GND 0.477993f
C6914 VDD.n4618 GND 0.477993f
C6915 VDD.n4619 GND 0.477993f
C6916 VDD.n4620 GND 0.006693f
C6917 VDD.n4621 GND 0.005387f
C6918 VDD.n4622 GND 0.005387f
C6919 VDD.n4623 GND 0.005387f
C6920 VDD.n4624 GND 0.006693f
C6921 VDD.n4625 GND 0.477993f
C6922 VDD.n4626 GND 0.477993f
C6923 VDD.n4627 GND 0.477993f
C6924 VDD.n4628 GND 0.006693f
C6925 VDD.n4629 GND 0.005387f
C6926 VDD.n4630 GND 0.005387f
C6927 VDD.n4631 GND 0.005387f
C6928 VDD.n4632 GND 0.006693f
C6929 VDD.n4633 GND 0.477993f
C6930 VDD.n4634 GND 0.477993f
C6931 VDD.n4635 GND 0.382394f
C6932 VDD.n4636 GND 0.006693f
C6933 VDD.n4637 GND 0.005387f
C6934 VDD.n4638 GND 0.005387f
C6935 VDD.n4639 GND 0.005387f
C6936 VDD.n4640 GND 0.006693f
C6937 VDD.n4641 GND 0.477993f
C6938 VDD.n4642 GND 0.477993f
C6939 VDD.n4643 GND 0.477993f
C6940 VDD.n4644 GND 0.006693f
C6941 VDD.n4645 GND 0.005387f
C6942 VDD.n4646 GND 0.005387f
C6943 VDD.n4647 GND 0.005387f
C6944 VDD.n4648 GND 0.006693f
C6945 VDD.n4649 GND 0.477993f
C6946 VDD.n4650 GND 0.477993f
C6947 VDD.n4651 GND 0.477993f
C6948 VDD.n4652 GND 0.006693f
C6949 VDD.n4653 GND 0.005387f
C6950 VDD.n4654 GND 0.005387f
C6951 VDD.n4655 GND 0.005387f
C6952 VDD.n4656 GND 0.006693f
C6953 VDD.n4657 GND 0.477993f
C6954 VDD.n4658 GND 0.477993f
C6955 VDD.n4659 GND 0.454093f
C6956 VDD.n4660 GND 0.006693f
C6957 VDD.n4661 GND 0.005387f
C6958 VDD.n4662 GND 0.005387f
C6959 VDD.n4663 GND 0.005387f
C6960 VDD.n4664 GND 0.006693f
C6961 VDD.n4665 GND 0.477993f
C6962 VDD.n4666 GND 0.477993f
C6963 VDD.n4667 GND 0.477993f
C6964 VDD.n4668 GND 0.006693f
C6965 VDD.n4669 GND 0.005387f
C6966 VDD.n4670 GND 0.005387f
C6967 VDD.n4671 GND 0.005387f
C6968 VDD.n4672 GND 0.006693f
C6969 VDD.n4673 GND 0.477993f
C6970 VDD.n4674 GND 0.477993f
C6971 VDD.n4675 GND 0.477993f
C6972 VDD.n4676 GND 0.006693f
C6973 VDD.n4677 GND 0.005387f
C6974 VDD.n4678 GND 0.005387f
C6975 VDD.n4679 GND 0.005387f
C6976 VDD.n4680 GND 0.006693f
C6977 VDD.n4681 GND 0.477993f
C6978 VDD.n4682 GND 0.477993f
C6979 VDD.n4683 GND 0.477993f
C6980 VDD.n4684 GND 0.006693f
C6981 VDD.n4685 GND 0.005387f
C6982 VDD.n4686 GND 0.005387f
C6983 VDD.n4687 GND 0.005387f
C6984 VDD.n4688 GND 0.006693f
C6985 VDD.n4689 GND 0.430194f
C6986 VDD.n4690 GND 0.477993f
C6987 VDD.n4691 GND 0.477993f
C6988 VDD.n4692 GND 0.006693f
C6989 VDD.n4693 GND 0.005387f
C6990 VDD.n4694 GND 0.005387f
C6991 VDD.n4695 GND 0.005387f
C6992 VDD.n4696 GND 0.006693f
C6993 VDD.n4697 GND 0.477993f
C6994 VDD.n4698 GND 0.477993f
C6995 VDD.n4699 GND 0.477993f
C6996 VDD.n4700 GND 0.006693f
C6997 VDD.n4701 GND 0.005387f
C6998 VDD.n4702 GND 0.005387f
C6999 VDD.n4703 GND 0.005387f
C7000 VDD.n4704 GND 0.006693f
C7001 VDD.n4705 GND 0.477993f
C7002 VDD.n4706 GND 0.477993f
C7003 VDD.n4707 GND 0.477993f
C7004 VDD.n4708 GND 0.006693f
C7005 VDD.n4709 GND 0.005387f
C7006 VDD.n4710 GND 0.005387f
C7007 VDD.n4711 GND 0.005144f
C7008 VDD.n4712 GND 0.409661f
C7009 VDD.n4713 GND 4.09504f
C7010 VOUT.t45 GND 0.038152f
C7011 VOUT.t58 GND 0.038152f
C7012 VOUT.n0 GND 0.19536f
C7013 VOUT.t53 GND 0.038152f
C7014 VOUT.t72 GND 0.038152f
C7015 VOUT.n1 GND 0.181021f
C7016 VOUT.n2 GND 2.00355f
C7017 VOUT.t51 GND 0.038152f
C7018 VOUT.t48 GND 0.038152f
C7019 VOUT.n3 GND 0.181021f
C7020 VOUT.n4 GND 1.00419f
C7021 VOUT.t65 GND 0.237011f
C7022 VOUT.n5 GND 0.823346f
C7023 VOUT.t77 GND 0.038152f
C7024 VOUT.t76 GND 0.038152f
C7025 VOUT.n6 GND 0.19536f
C7026 VOUT.t85 GND 0.038152f
C7027 VOUT.t47 GND 0.038152f
C7028 VOUT.n7 GND 0.181021f
C7029 VOUT.n8 GND 2.00355f
C7030 VOUT.t83 GND 0.038152f
C7031 VOUT.t46 GND 0.038152f
C7032 VOUT.n9 GND 0.181021f
C7033 VOUT.n10 GND 1.00419f
C7034 VOUT.t61 GND 0.237011f
C7035 VOUT.n11 GND 0.785542f
C7036 VOUT.n12 GND 0.626119f
C7037 VOUT.t59 GND 0.038152f
C7038 VOUT.t79 GND 0.038152f
C7039 VOUT.n13 GND 0.19536f
C7040 VOUT.t75 GND 0.038152f
C7041 VOUT.t57 GND 0.038152f
C7042 VOUT.n14 GND 0.181021f
C7043 VOUT.n15 GND 2.00355f
C7044 VOUT.t63 GND 0.038152f
C7045 VOUT.t71 GND 0.038152f
C7046 VOUT.n16 GND 0.181021f
C7047 VOUT.n17 GND 1.00419f
C7048 VOUT.t67 GND 0.237011f
C7049 VOUT.n18 GND 0.785542f
C7050 VOUT.n19 GND 0.902685f
C7051 VOUT.n20 GND 16.455198f
C7052 VOUT.t106 GND 4.38863f
C7053 VOUT.n21 GND 3.67036f
C7054 VOUT.t109 GND 4.4039f
C7055 VOUT.t107 GND 4.41445f
C7056 VOUT.n22 GND 4.18692f
C7057 VOUT.n23 GND 4.1863f
C7058 VOUT.t108 GND 4.38863f
C7059 VOUT.n24 GND 1.63019f
C7060 VOUT.n25 GND 5.51987f
C7061 VOUT.n26 GND 2.23526f
C7062 VOUT.t52 GND 0.244811f
C7063 VOUT.t56 GND 0.038152f
C7064 VOUT.t74 GND 0.038152f
C7065 VOUT.n27 GND 0.181021f
C7066 VOUT.n28 GND 1.64128f
C7067 VOUT.t62 GND 0.038152f
C7068 VOUT.t82 GND 0.038152f
C7069 VOUT.n29 GND 0.181021f
C7070 VOUT.n30 GND 1.00419f
C7071 VOUT.t54 GND 0.038152f
C7072 VOUT.t69 GND 0.038152f
C7073 VOUT.n31 GND 0.181021f
C7074 VOUT.n32 GND 1.14023f
C7075 VOUT.t84 GND 0.244811f
C7076 VOUT.t55 GND 0.038152f
C7077 VOUT.t70 GND 0.038152f
C7078 VOUT.n33 GND 0.181021f
C7079 VOUT.n34 GND 1.64128f
C7080 VOUT.t60 GND 0.038152f
C7081 VOUT.t80 GND 0.038152f
C7082 VOUT.n35 GND 0.181021f
C7083 VOUT.n36 GND 1.00419f
C7084 VOUT.t73 GND 0.038152f
C7085 VOUT.t68 GND 0.038152f
C7086 VOUT.n37 GND 0.181021f
C7087 VOUT.n38 GND 1.09977f
C7088 VOUT.n39 GND 0.73261f
C7089 VOUT.t66 GND 0.244811f
C7090 VOUT.t86 GND 0.038152f
C7091 VOUT.t81 GND 0.038152f
C7092 VOUT.n40 GND 0.181021f
C7093 VOUT.n41 GND 1.64128f
C7094 VOUT.t49 GND 0.038152f
C7095 VOUT.t64 GND 0.038152f
C7096 VOUT.n42 GND 0.181021f
C7097 VOUT.n43 GND 1.00419f
C7098 VOUT.t78 GND 0.038152f
C7099 VOUT.t50 GND 0.038152f
C7100 VOUT.n44 GND 0.18102f
C7101 VOUT.n45 GND 1.09977f
C7102 VOUT.n46 GND 0.957255f
C7103 VOUT.n47 GND 19.839401f
C7104 VOUT.t94 GND 0.046354f
C7105 VOUT.t92 GND 0.046354f
C7106 VOUT.n48 GND 0.333413f
C7107 VOUT.t39 GND 0.046354f
C7108 VOUT.t3 GND 0.046354f
C7109 VOUT.n49 GND 0.307898f
C7110 VOUT.n50 GND 1.95499f
C7111 VOUT.t2 GND 0.046354f
C7112 VOUT.t36 GND 0.046354f
C7113 VOUT.n51 GND 0.307898f
C7114 VOUT.n52 GND 0.985501f
C7115 VOUT.t93 GND 0.046354f
C7116 VOUT.t22 GND 0.046354f
C7117 VOUT.n53 GND 0.307898f
C7118 VOUT.n54 GND 1.12431f
C7119 VOUT.t40 GND 0.046354f
C7120 VOUT.t23 GND 0.046354f
C7121 VOUT.n55 GND 0.333413f
C7122 VOUT.t44 GND 0.046354f
C7123 VOUT.t98 GND 0.046354f
C7124 VOUT.n56 GND 0.307898f
C7125 VOUT.n57 GND 1.95499f
C7126 VOUT.t19 GND 0.046354f
C7127 VOUT.t11 GND 0.046354f
C7128 VOUT.n58 GND 0.307898f
C7129 VOUT.n59 GND 0.985501f
C7130 VOUT.t32 GND 0.046354f
C7131 VOUT.t25 GND 0.046354f
C7132 VOUT.n60 GND 0.307898f
C7133 VOUT.n61 GND 1.07675f
C7134 VOUT.n62 GND 0.799047f
C7135 VOUT.t1 GND 0.046354f
C7136 VOUT.t8 GND 0.046354f
C7137 VOUT.n63 GND 0.333413f
C7138 VOUT.t14 GND 0.046354f
C7139 VOUT.t31 GND 0.046354f
C7140 VOUT.n64 GND 0.307898f
C7141 VOUT.n65 GND 1.95499f
C7142 VOUT.t95 GND 0.046354f
C7143 VOUT.t105 GND 0.046354f
C7144 VOUT.n66 GND 0.307898f
C7145 VOUT.n67 GND 0.985501f
C7146 VOUT.t35 GND 0.046354f
C7147 VOUT.t4 GND 0.046354f
C7148 VOUT.n68 GND 0.307898f
C7149 VOUT.n69 GND 1.07675f
C7150 VOUT.n70 GND 0.533552f
C7151 VOUT.t29 GND 0.046354f
C7152 VOUT.t103 GND 0.046354f
C7153 VOUT.n71 GND 0.333413f
C7154 VOUT.t43 GND 0.046354f
C7155 VOUT.t97 GND 0.046354f
C7156 VOUT.n72 GND 0.307898f
C7157 VOUT.n73 GND 1.95499f
C7158 VOUT.t101 GND 0.046354f
C7159 VOUT.t10 GND 0.046354f
C7160 VOUT.n74 GND 0.307898f
C7161 VOUT.n75 GND 0.985501f
C7162 VOUT.t13 GND 0.046354f
C7163 VOUT.t33 GND 0.046354f
C7164 VOUT.n76 GND 0.307898f
C7165 VOUT.n77 GND 1.07675f
C7166 VOUT.n78 GND 0.836986f
C7167 VOUT.n79 GND 18.5728f
C7168 VOUT.t99 GND 0.046354f
C7169 VOUT.t5 GND 0.046354f
C7170 VOUT.n80 GND 0.333413f
C7171 VOUT.t34 GND 0.046354f
C7172 VOUT.t7 GND 0.046354f
C7173 VOUT.n81 GND 0.307898f
C7174 VOUT.n82 GND 1.95499f
C7175 VOUT.t12 GND 0.046354f
C7176 VOUT.t17 GND 0.046354f
C7177 VOUT.n83 GND 0.307898f
C7178 VOUT.n84 GND 0.985501f
C7179 VOUT.t24 GND 0.046354f
C7180 VOUT.t37 GND 0.046354f
C7181 VOUT.n85 GND 0.307898f
C7182 VOUT.n86 GND 1.12431f
C7183 VOUT.t88 GND 0.046354f
C7184 VOUT.t16 GND 0.046354f
C7185 VOUT.n87 GND 0.333413f
C7186 VOUT.t28 GND 0.046354f
C7187 VOUT.t102 GND 0.046354f
C7188 VOUT.n88 GND 0.307898f
C7189 VOUT.n89 GND 1.95499f
C7190 VOUT.t21 GND 0.046354f
C7191 VOUT.t15 GND 0.046354f
C7192 VOUT.n90 GND 0.307898f
C7193 VOUT.n91 GND 0.985501f
C7194 VOUT.t90 GND 0.046354f
C7195 VOUT.t0 GND 0.046354f
C7196 VOUT.n92 GND 0.307898f
C7197 VOUT.n93 GND 1.07675f
C7198 VOUT.n94 GND 0.799047f
C7199 VOUT.t38 GND 0.046354f
C7200 VOUT.t42 GND 0.046354f
C7201 VOUT.n95 GND 0.333413f
C7202 VOUT.t30 GND 0.046354f
C7203 VOUT.t91 GND 0.046354f
C7204 VOUT.n96 GND 0.307898f
C7205 VOUT.n97 GND 1.95499f
C7206 VOUT.t26 GND 0.046354f
C7207 VOUT.t41 GND 0.046354f
C7208 VOUT.n98 GND 0.307898f
C7209 VOUT.n99 GND 0.985501f
C7210 VOUT.t104 GND 0.046354f
C7211 VOUT.t9 GND 0.046354f
C7212 VOUT.n100 GND 0.307898f
C7213 VOUT.n101 GND 1.07675f
C7214 VOUT.n102 GND 0.533552f
C7215 VOUT.t87 GND 0.046354f
C7216 VOUT.t18 GND 0.046354f
C7217 VOUT.n103 GND 0.333413f
C7218 VOUT.t27 GND 0.046354f
C7219 VOUT.t96 GND 0.046354f
C7220 VOUT.n104 GND 0.307898f
C7221 VOUT.n105 GND 1.95499f
C7222 VOUT.t20 GND 0.046354f
C7223 VOUT.t100 GND 0.046354f
C7224 VOUT.n106 GND 0.307898f
C7225 VOUT.n107 GND 0.985501f
C7226 VOUT.t89 GND 0.046354f
C7227 VOUT.t6 GND 0.046354f
C7228 VOUT.n108 GND 0.307898f
C7229 VOUT.n109 GND 1.07675f
C7230 VOUT.n110 GND 0.836986f
C7231 VOUT.n111 GND 15.079099f
C7232 VOUT.n112 GND 7.00493f
C7233 a_n24758_8502.n0 GND 4.48003f
C7234 a_n24758_8502.n1 GND 0.837436f
C7235 a_n24758_8502.n2 GND 4.48003f
C7236 a_n24758_8502.n3 GND 0.837436f
C7237 a_n24758_8502.n4 GND 4.53025f
C7238 a_n24758_8502.n5 GND 0.837436f
C7239 a_n24758_8502.n6 GND 5.40161f
C7240 a_n24758_8502.n7 GND 0.84157f
C7241 a_n24758_8502.n8 GND 5.35139f
C7242 a_n24758_8502.n9 GND 0.84157f
C7243 a_n24758_8502.n10 GND 5.35139f
C7244 a_n24758_8502.n11 GND 0.84157f
C7245 a_n24758_8502.n12 GND 0.837192f
C7246 a_n24758_8502.n13 GND 0.854804f
C7247 a_n24758_8502.n14 GND 0.837192f
C7248 a_n24758_8502.n15 GND 0.854804f
C7249 a_n24758_8502.n16 GND 0.837192f
C7250 a_n24758_8502.n17 GND 0.854804f
C7251 a_n24758_8502.n18 GND 0.854812f
C7252 a_n24758_8502.n19 GND 0.854812f
C7253 a_n24758_8502.n20 GND 0.854812f
C7254 a_n24758_8502.n21 GND 2.55434f
C7255 a_n24758_8502.n22 GND 3.74769f
C7256 a_n24758_8502.n23 GND 6.57511f
C7257 a_n24758_8502.t3 GND 0.117868f
C7258 a_n24758_8502.t13 GND 0.075744f
C7259 a_n24758_8502.t14 GND 0.075744f
C7260 a_n24758_8502.n24 GND 0.411352f
C7261 a_n24758_8502.t17 GND 0.495368f
C7262 a_n24758_8502.n25 GND 8.691099f
C7263 a_n24758_8502.t12 GND 0.511913f
C7264 a_n24758_8502.t7 GND 0.075744f
C7265 a_n24758_8502.t9 GND 0.075744f
C7266 a_n24758_8502.n26 GND 0.381518f
C7267 a_n24758_8502.n27 GND 7.45765f
C7268 a_n24758_8502.n28 GND 14.1683f
C7269 a_n24758_8502.t31 GND 1.91462f
C7270 a_n24758_8502.t52 GND 1.92976f
C7271 a_n24758_8502.t54 GND 1.91286f
C7272 a_n24758_8502.t37 GND 1.91301f
C7273 a_n24758_8502.t44 GND 1.9048f
C7274 a_n24758_8502.t48 GND 1.9455f
C7275 a_n24758_8502.t50 GND 1.91283f
C7276 a_n24758_8502.t53 GND 1.91462f
C7277 a_n24758_8502.t40 GND 1.92976f
C7278 a_n24758_8502.t25 GND 1.91286f
C7279 a_n24758_8502.t41 GND 1.91301f
C7280 a_n24758_8502.t27 GND 1.9048f
C7281 a_n24758_8502.t46 GND 1.9455f
C7282 a_n24758_8502.t19 GND 1.91283f
C7283 a_n24758_8502.t51 GND 1.91462f
C7284 a_n24758_8502.t36 GND 1.92976f
C7285 a_n24758_8502.t20 GND 1.91286f
C7286 a_n24758_8502.t39 GND 1.91301f
C7287 a_n24758_8502.t22 GND 1.9048f
C7288 a_n24758_8502.t42 GND 1.9455f
C7289 a_n24758_8502.t59 GND 1.91283f
C7290 a_n24758_8502.t49 GND 1.95081f
C7291 a_n24758_8502.t24 GND 1.90475f
C7292 a_n24758_8502.t29 GND 1.91145f
C7293 a_n24758_8502.t38 GND 1.91282f
C7294 a_n24758_8502.t43 GND 1.89945f
C7295 a_n24758_8502.t18 GND 1.94692f
C7296 a_n24758_8502.t23 GND 1.9455f
C7297 a_n24758_8502.t26 GND 1.95081f
C7298 a_n24758_8502.t33 GND 1.90475f
C7299 a_n24758_8502.t56 GND 1.91145f
C7300 a_n24758_8502.t47 GND 1.91282f
C7301 a_n24758_8502.t30 GND 1.89945f
C7302 a_n24758_8502.t35 GND 1.94692f
C7303 a_n24758_8502.t58 GND 1.9455f
C7304 a_n24758_8502.t21 GND 1.95081f
C7305 a_n24758_8502.t32 GND 1.90475f
C7306 a_n24758_8502.t55 GND 1.91145f
C7307 a_n24758_8502.t45 GND 1.91282f
C7308 a_n24758_8502.t28 GND 1.89945f
C7309 a_n24758_8502.t34 GND 1.94692f
C7310 a_n24758_8502.t57 GND 1.9455f
C7311 a_n24758_8502.n29 GND 24.9052f
C7312 a_n24758_8502.n30 GND 2.7169f
C7313 a_n24758_8502.t15 GND 0.117868f
C7314 a_n24758_8502.t10 GND 0.117868f
C7315 a_n24758_8502.n31 GND 0.856084f
C7316 a_n24758_8502.t8 GND 0.117868f
C7317 a_n24758_8502.t1 GND 0.117868f
C7318 a_n24758_8502.n32 GND 0.836121f
C7319 a_n24758_8502.t2 GND 0.117868f
C7320 a_n24758_8502.t5 GND 0.117868f
C7321 a_n24758_8502.n33 GND 0.836121f
C7322 a_n24758_8502.t6 GND 0.117868f
C7323 a_n24758_8502.t4 GND 0.117868f
C7324 a_n24758_8502.n34 GND 0.856081f
C7325 a_n24758_8502.t16 GND 0.117868f
C7326 a_n24758_8502.t11 GND 0.117868f
C7327 a_n24758_8502.n35 GND 0.856081f
C7328 a_n24758_8502.n36 GND 6.60253f
C7329 a_n24758_8502.n37 GND 0.836117f
C7330 a_n24758_8502.t0 GND 0.117868f
.ends

