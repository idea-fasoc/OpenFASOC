* NGSPICE file created from diff_pair_sample_0977.ext - technology: sky130A

.subckt diff_pair_sample_0977 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t7 w_n2296_n2514# sky130_fd_pr__pfet_01v8 ad=1.27545 pd=8.06 as=3.0147 ps=16.24 w=7.73 l=1.88
X1 VTAIL.t2 VN.t0 VDD2.t3 w_n2296_n2514# sky130_fd_pr__pfet_01v8 ad=3.0147 pd=16.24 as=1.27545 ps=8.06 w=7.73 l=1.88
X2 VDD2.t2 VN.t1 VTAIL.t3 w_n2296_n2514# sky130_fd_pr__pfet_01v8 ad=1.27545 pd=8.06 as=3.0147 ps=16.24 w=7.73 l=1.88
X3 VDD1.t2 VP.t1 VTAIL.t4 w_n2296_n2514# sky130_fd_pr__pfet_01v8 ad=1.27545 pd=8.06 as=3.0147 ps=16.24 w=7.73 l=1.88
X4 VTAIL.t5 VP.t2 VDD1.t1 w_n2296_n2514# sky130_fd_pr__pfet_01v8 ad=3.0147 pd=16.24 as=1.27545 ps=8.06 w=7.73 l=1.88
X5 VDD2.t1 VN.t2 VTAIL.t1 w_n2296_n2514# sky130_fd_pr__pfet_01v8 ad=1.27545 pd=8.06 as=3.0147 ps=16.24 w=7.73 l=1.88
X6 B.t11 B.t9 B.t10 w_n2296_n2514# sky130_fd_pr__pfet_01v8 ad=3.0147 pd=16.24 as=0 ps=0 w=7.73 l=1.88
X7 B.t8 B.t6 B.t7 w_n2296_n2514# sky130_fd_pr__pfet_01v8 ad=3.0147 pd=16.24 as=0 ps=0 w=7.73 l=1.88
X8 VTAIL.t0 VN.t3 VDD2.t0 w_n2296_n2514# sky130_fd_pr__pfet_01v8 ad=3.0147 pd=16.24 as=1.27545 ps=8.06 w=7.73 l=1.88
X9 B.t5 B.t3 B.t4 w_n2296_n2514# sky130_fd_pr__pfet_01v8 ad=3.0147 pd=16.24 as=0 ps=0 w=7.73 l=1.88
X10 B.t2 B.t0 B.t1 w_n2296_n2514# sky130_fd_pr__pfet_01v8 ad=3.0147 pd=16.24 as=0 ps=0 w=7.73 l=1.88
X11 VTAIL.t6 VP.t3 VDD1.t0 w_n2296_n2514# sky130_fd_pr__pfet_01v8 ad=3.0147 pd=16.24 as=1.27545 ps=8.06 w=7.73 l=1.88
R0 VP.n5 VP.n4 180.63
R1 VP.n14 VP.n13 180.63
R2 VP.n12 VP.n0 161.3
R3 VP.n11 VP.n10 161.3
R4 VP.n9 VP.n1 161.3
R5 VP.n8 VP.n7 161.3
R6 VP.n6 VP.n2 161.3
R7 VP.n3 VP.t3 136.806
R8 VP.n3 VP.t0 136.369
R9 VP.n5 VP.t2 99.0925
R10 VP.n13 VP.t1 99.0925
R11 VP.n4 VP.n3 49.959
R12 VP.n7 VP.n1 40.4934
R13 VP.n11 VP.n1 40.4934
R14 VP.n7 VP.n6 24.4675
R15 VP.n12 VP.n11 24.4675
R16 VP.n6 VP.n5 5.13857
R17 VP.n13 VP.n12 5.13857
R18 VP.n4 VP.n2 0.189894
R19 VP.n8 VP.n2 0.189894
R20 VP.n9 VP.n8 0.189894
R21 VP.n10 VP.n9 0.189894
R22 VP.n10 VP.n0 0.189894
R23 VP.n14 VP.n0 0.189894
R24 VP VP.n14 0.0516364
R25 VTAIL.n6 VTAIL.t7 70.1508
R26 VTAIL.n5 VTAIL.t6 70.1507
R27 VTAIL.n4 VTAIL.t1 70.1507
R28 VTAIL.n3 VTAIL.t0 70.1507
R29 VTAIL.n7 VTAIL.t3 70.1506
R30 VTAIL.n0 VTAIL.t2 70.1506
R31 VTAIL.n1 VTAIL.t4 70.1506
R32 VTAIL.n2 VTAIL.t5 70.1506
R33 VTAIL.n7 VTAIL.n6 20.9358
R34 VTAIL.n3 VTAIL.n2 20.9358
R35 VTAIL.n4 VTAIL.n3 1.90567
R36 VTAIL.n6 VTAIL.n5 1.90567
R37 VTAIL.n2 VTAIL.n1 1.90567
R38 VTAIL VTAIL.n0 1.01128
R39 VTAIL VTAIL.n7 0.894897
R40 VTAIL.n5 VTAIL.n4 0.470328
R41 VTAIL.n1 VTAIL.n0 0.470328
R42 VDD1 VDD1.n1 119.243
R43 VDD1 VDD1.n0 82.6827
R44 VDD1.n0 VDD1.t0 4.20555
R45 VDD1.n0 VDD1.t3 4.20555
R46 VDD1.n1 VDD1.t1 4.20555
R47 VDD1.n1 VDD1.t2 4.20555
R48 VN.n0 VN.t0 136.806
R49 VN.n1 VN.t2 136.806
R50 VN.n0 VN.t1 136.369
R51 VN.n1 VN.t3 136.369
R52 VN VN.n1 50.3397
R53 VN VN.n0 9.12382
R54 VDD2.n2 VDD2.n0 118.719
R55 VDD2.n2 VDD2.n1 82.6245
R56 VDD2.n1 VDD2.t0 4.20555
R57 VDD2.n1 VDD2.t1 4.20555
R58 VDD2.n0 VDD2.t3 4.20555
R59 VDD2.n0 VDD2.t2 4.20555
R60 VDD2 VDD2.n2 0.0586897
R61 B.n275 B.n82 585
R62 B.n274 B.n273 585
R63 B.n272 B.n83 585
R64 B.n271 B.n270 585
R65 B.n269 B.n84 585
R66 B.n268 B.n267 585
R67 B.n266 B.n85 585
R68 B.n265 B.n264 585
R69 B.n263 B.n86 585
R70 B.n262 B.n261 585
R71 B.n260 B.n87 585
R72 B.n259 B.n258 585
R73 B.n257 B.n88 585
R74 B.n256 B.n255 585
R75 B.n254 B.n89 585
R76 B.n253 B.n252 585
R77 B.n251 B.n90 585
R78 B.n250 B.n249 585
R79 B.n248 B.n91 585
R80 B.n247 B.n246 585
R81 B.n245 B.n92 585
R82 B.n244 B.n243 585
R83 B.n242 B.n93 585
R84 B.n241 B.n240 585
R85 B.n239 B.n94 585
R86 B.n238 B.n237 585
R87 B.n236 B.n95 585
R88 B.n235 B.n234 585
R89 B.n233 B.n96 585
R90 B.n232 B.n231 585
R91 B.n227 B.n97 585
R92 B.n226 B.n225 585
R93 B.n224 B.n98 585
R94 B.n223 B.n222 585
R95 B.n221 B.n99 585
R96 B.n220 B.n219 585
R97 B.n218 B.n100 585
R98 B.n217 B.n216 585
R99 B.n215 B.n101 585
R100 B.n213 B.n212 585
R101 B.n211 B.n104 585
R102 B.n210 B.n209 585
R103 B.n208 B.n105 585
R104 B.n207 B.n206 585
R105 B.n205 B.n106 585
R106 B.n204 B.n203 585
R107 B.n202 B.n107 585
R108 B.n201 B.n200 585
R109 B.n199 B.n108 585
R110 B.n198 B.n197 585
R111 B.n196 B.n109 585
R112 B.n195 B.n194 585
R113 B.n193 B.n110 585
R114 B.n192 B.n191 585
R115 B.n190 B.n111 585
R116 B.n189 B.n188 585
R117 B.n187 B.n112 585
R118 B.n186 B.n185 585
R119 B.n184 B.n113 585
R120 B.n183 B.n182 585
R121 B.n181 B.n114 585
R122 B.n180 B.n179 585
R123 B.n178 B.n115 585
R124 B.n177 B.n176 585
R125 B.n175 B.n116 585
R126 B.n174 B.n173 585
R127 B.n172 B.n117 585
R128 B.n171 B.n170 585
R129 B.n277 B.n276 585
R130 B.n278 B.n81 585
R131 B.n280 B.n279 585
R132 B.n281 B.n80 585
R133 B.n283 B.n282 585
R134 B.n284 B.n79 585
R135 B.n286 B.n285 585
R136 B.n287 B.n78 585
R137 B.n289 B.n288 585
R138 B.n290 B.n77 585
R139 B.n292 B.n291 585
R140 B.n293 B.n76 585
R141 B.n295 B.n294 585
R142 B.n296 B.n75 585
R143 B.n298 B.n297 585
R144 B.n299 B.n74 585
R145 B.n301 B.n300 585
R146 B.n302 B.n73 585
R147 B.n304 B.n303 585
R148 B.n305 B.n72 585
R149 B.n307 B.n306 585
R150 B.n308 B.n71 585
R151 B.n310 B.n309 585
R152 B.n311 B.n70 585
R153 B.n313 B.n312 585
R154 B.n314 B.n69 585
R155 B.n316 B.n315 585
R156 B.n317 B.n68 585
R157 B.n319 B.n318 585
R158 B.n320 B.n67 585
R159 B.n322 B.n321 585
R160 B.n323 B.n66 585
R161 B.n325 B.n324 585
R162 B.n326 B.n65 585
R163 B.n328 B.n327 585
R164 B.n329 B.n64 585
R165 B.n331 B.n330 585
R166 B.n332 B.n63 585
R167 B.n334 B.n333 585
R168 B.n335 B.n62 585
R169 B.n337 B.n336 585
R170 B.n338 B.n61 585
R171 B.n340 B.n339 585
R172 B.n341 B.n60 585
R173 B.n343 B.n342 585
R174 B.n344 B.n59 585
R175 B.n346 B.n345 585
R176 B.n347 B.n58 585
R177 B.n349 B.n348 585
R178 B.n350 B.n57 585
R179 B.n352 B.n351 585
R180 B.n353 B.n56 585
R181 B.n355 B.n354 585
R182 B.n356 B.n55 585
R183 B.n358 B.n357 585
R184 B.n359 B.n54 585
R185 B.n463 B.n462 585
R186 B.n461 B.n16 585
R187 B.n460 B.n459 585
R188 B.n458 B.n17 585
R189 B.n457 B.n456 585
R190 B.n455 B.n18 585
R191 B.n454 B.n453 585
R192 B.n452 B.n19 585
R193 B.n451 B.n450 585
R194 B.n449 B.n20 585
R195 B.n448 B.n447 585
R196 B.n446 B.n21 585
R197 B.n445 B.n444 585
R198 B.n443 B.n22 585
R199 B.n442 B.n441 585
R200 B.n440 B.n23 585
R201 B.n439 B.n438 585
R202 B.n437 B.n24 585
R203 B.n436 B.n435 585
R204 B.n434 B.n25 585
R205 B.n433 B.n432 585
R206 B.n431 B.n26 585
R207 B.n430 B.n429 585
R208 B.n428 B.n27 585
R209 B.n427 B.n426 585
R210 B.n425 B.n28 585
R211 B.n424 B.n423 585
R212 B.n422 B.n29 585
R213 B.n421 B.n420 585
R214 B.n419 B.n418 585
R215 B.n417 B.n33 585
R216 B.n416 B.n415 585
R217 B.n414 B.n34 585
R218 B.n413 B.n412 585
R219 B.n411 B.n35 585
R220 B.n410 B.n409 585
R221 B.n408 B.n36 585
R222 B.n407 B.n406 585
R223 B.n405 B.n37 585
R224 B.n403 B.n402 585
R225 B.n401 B.n40 585
R226 B.n400 B.n399 585
R227 B.n398 B.n41 585
R228 B.n397 B.n396 585
R229 B.n395 B.n42 585
R230 B.n394 B.n393 585
R231 B.n392 B.n43 585
R232 B.n391 B.n390 585
R233 B.n389 B.n44 585
R234 B.n388 B.n387 585
R235 B.n386 B.n45 585
R236 B.n385 B.n384 585
R237 B.n383 B.n46 585
R238 B.n382 B.n381 585
R239 B.n380 B.n47 585
R240 B.n379 B.n378 585
R241 B.n377 B.n48 585
R242 B.n376 B.n375 585
R243 B.n374 B.n49 585
R244 B.n373 B.n372 585
R245 B.n371 B.n50 585
R246 B.n370 B.n369 585
R247 B.n368 B.n51 585
R248 B.n367 B.n366 585
R249 B.n365 B.n52 585
R250 B.n364 B.n363 585
R251 B.n362 B.n53 585
R252 B.n361 B.n360 585
R253 B.n464 B.n15 585
R254 B.n466 B.n465 585
R255 B.n467 B.n14 585
R256 B.n469 B.n468 585
R257 B.n470 B.n13 585
R258 B.n472 B.n471 585
R259 B.n473 B.n12 585
R260 B.n475 B.n474 585
R261 B.n476 B.n11 585
R262 B.n478 B.n477 585
R263 B.n479 B.n10 585
R264 B.n481 B.n480 585
R265 B.n482 B.n9 585
R266 B.n484 B.n483 585
R267 B.n485 B.n8 585
R268 B.n487 B.n486 585
R269 B.n488 B.n7 585
R270 B.n490 B.n489 585
R271 B.n491 B.n6 585
R272 B.n493 B.n492 585
R273 B.n494 B.n5 585
R274 B.n496 B.n495 585
R275 B.n497 B.n4 585
R276 B.n499 B.n498 585
R277 B.n500 B.n3 585
R278 B.n502 B.n501 585
R279 B.n503 B.n0 585
R280 B.n2 B.n1 585
R281 B.n132 B.n131 585
R282 B.n133 B.n130 585
R283 B.n135 B.n134 585
R284 B.n136 B.n129 585
R285 B.n138 B.n137 585
R286 B.n139 B.n128 585
R287 B.n141 B.n140 585
R288 B.n142 B.n127 585
R289 B.n144 B.n143 585
R290 B.n145 B.n126 585
R291 B.n147 B.n146 585
R292 B.n148 B.n125 585
R293 B.n150 B.n149 585
R294 B.n151 B.n124 585
R295 B.n153 B.n152 585
R296 B.n154 B.n123 585
R297 B.n156 B.n155 585
R298 B.n157 B.n122 585
R299 B.n159 B.n158 585
R300 B.n160 B.n121 585
R301 B.n162 B.n161 585
R302 B.n163 B.n120 585
R303 B.n165 B.n164 585
R304 B.n166 B.n119 585
R305 B.n168 B.n167 585
R306 B.n169 B.n118 585
R307 B.n170 B.n169 492.5
R308 B.n276 B.n275 492.5
R309 B.n360 B.n359 492.5
R310 B.n462 B.n15 492.5
R311 B.n102 B.t0 305.714
R312 B.n228 B.t6 305.714
R313 B.n38 B.t9 305.714
R314 B.n30 B.t3 305.714
R315 B.n505 B.n504 256.663
R316 B.n504 B.n503 235.042
R317 B.n504 B.n2 235.042
R318 B.n170 B.n117 163.367
R319 B.n174 B.n117 163.367
R320 B.n175 B.n174 163.367
R321 B.n176 B.n175 163.367
R322 B.n176 B.n115 163.367
R323 B.n180 B.n115 163.367
R324 B.n181 B.n180 163.367
R325 B.n182 B.n181 163.367
R326 B.n182 B.n113 163.367
R327 B.n186 B.n113 163.367
R328 B.n187 B.n186 163.367
R329 B.n188 B.n187 163.367
R330 B.n188 B.n111 163.367
R331 B.n192 B.n111 163.367
R332 B.n193 B.n192 163.367
R333 B.n194 B.n193 163.367
R334 B.n194 B.n109 163.367
R335 B.n198 B.n109 163.367
R336 B.n199 B.n198 163.367
R337 B.n200 B.n199 163.367
R338 B.n200 B.n107 163.367
R339 B.n204 B.n107 163.367
R340 B.n205 B.n204 163.367
R341 B.n206 B.n205 163.367
R342 B.n206 B.n105 163.367
R343 B.n210 B.n105 163.367
R344 B.n211 B.n210 163.367
R345 B.n212 B.n211 163.367
R346 B.n212 B.n101 163.367
R347 B.n217 B.n101 163.367
R348 B.n218 B.n217 163.367
R349 B.n219 B.n218 163.367
R350 B.n219 B.n99 163.367
R351 B.n223 B.n99 163.367
R352 B.n224 B.n223 163.367
R353 B.n225 B.n224 163.367
R354 B.n225 B.n97 163.367
R355 B.n232 B.n97 163.367
R356 B.n233 B.n232 163.367
R357 B.n234 B.n233 163.367
R358 B.n234 B.n95 163.367
R359 B.n238 B.n95 163.367
R360 B.n239 B.n238 163.367
R361 B.n240 B.n239 163.367
R362 B.n240 B.n93 163.367
R363 B.n244 B.n93 163.367
R364 B.n245 B.n244 163.367
R365 B.n246 B.n245 163.367
R366 B.n246 B.n91 163.367
R367 B.n250 B.n91 163.367
R368 B.n251 B.n250 163.367
R369 B.n252 B.n251 163.367
R370 B.n252 B.n89 163.367
R371 B.n256 B.n89 163.367
R372 B.n257 B.n256 163.367
R373 B.n258 B.n257 163.367
R374 B.n258 B.n87 163.367
R375 B.n262 B.n87 163.367
R376 B.n263 B.n262 163.367
R377 B.n264 B.n263 163.367
R378 B.n264 B.n85 163.367
R379 B.n268 B.n85 163.367
R380 B.n269 B.n268 163.367
R381 B.n270 B.n269 163.367
R382 B.n270 B.n83 163.367
R383 B.n274 B.n83 163.367
R384 B.n275 B.n274 163.367
R385 B.n359 B.n358 163.367
R386 B.n358 B.n55 163.367
R387 B.n354 B.n55 163.367
R388 B.n354 B.n353 163.367
R389 B.n353 B.n352 163.367
R390 B.n352 B.n57 163.367
R391 B.n348 B.n57 163.367
R392 B.n348 B.n347 163.367
R393 B.n347 B.n346 163.367
R394 B.n346 B.n59 163.367
R395 B.n342 B.n59 163.367
R396 B.n342 B.n341 163.367
R397 B.n341 B.n340 163.367
R398 B.n340 B.n61 163.367
R399 B.n336 B.n61 163.367
R400 B.n336 B.n335 163.367
R401 B.n335 B.n334 163.367
R402 B.n334 B.n63 163.367
R403 B.n330 B.n63 163.367
R404 B.n330 B.n329 163.367
R405 B.n329 B.n328 163.367
R406 B.n328 B.n65 163.367
R407 B.n324 B.n65 163.367
R408 B.n324 B.n323 163.367
R409 B.n323 B.n322 163.367
R410 B.n322 B.n67 163.367
R411 B.n318 B.n67 163.367
R412 B.n318 B.n317 163.367
R413 B.n317 B.n316 163.367
R414 B.n316 B.n69 163.367
R415 B.n312 B.n69 163.367
R416 B.n312 B.n311 163.367
R417 B.n311 B.n310 163.367
R418 B.n310 B.n71 163.367
R419 B.n306 B.n71 163.367
R420 B.n306 B.n305 163.367
R421 B.n305 B.n304 163.367
R422 B.n304 B.n73 163.367
R423 B.n300 B.n73 163.367
R424 B.n300 B.n299 163.367
R425 B.n299 B.n298 163.367
R426 B.n298 B.n75 163.367
R427 B.n294 B.n75 163.367
R428 B.n294 B.n293 163.367
R429 B.n293 B.n292 163.367
R430 B.n292 B.n77 163.367
R431 B.n288 B.n77 163.367
R432 B.n288 B.n287 163.367
R433 B.n287 B.n286 163.367
R434 B.n286 B.n79 163.367
R435 B.n282 B.n79 163.367
R436 B.n282 B.n281 163.367
R437 B.n281 B.n280 163.367
R438 B.n280 B.n81 163.367
R439 B.n276 B.n81 163.367
R440 B.n462 B.n461 163.367
R441 B.n461 B.n460 163.367
R442 B.n460 B.n17 163.367
R443 B.n456 B.n17 163.367
R444 B.n456 B.n455 163.367
R445 B.n455 B.n454 163.367
R446 B.n454 B.n19 163.367
R447 B.n450 B.n19 163.367
R448 B.n450 B.n449 163.367
R449 B.n449 B.n448 163.367
R450 B.n448 B.n21 163.367
R451 B.n444 B.n21 163.367
R452 B.n444 B.n443 163.367
R453 B.n443 B.n442 163.367
R454 B.n442 B.n23 163.367
R455 B.n438 B.n23 163.367
R456 B.n438 B.n437 163.367
R457 B.n437 B.n436 163.367
R458 B.n436 B.n25 163.367
R459 B.n432 B.n25 163.367
R460 B.n432 B.n431 163.367
R461 B.n431 B.n430 163.367
R462 B.n430 B.n27 163.367
R463 B.n426 B.n27 163.367
R464 B.n426 B.n425 163.367
R465 B.n425 B.n424 163.367
R466 B.n424 B.n29 163.367
R467 B.n420 B.n29 163.367
R468 B.n420 B.n419 163.367
R469 B.n419 B.n33 163.367
R470 B.n415 B.n33 163.367
R471 B.n415 B.n414 163.367
R472 B.n414 B.n413 163.367
R473 B.n413 B.n35 163.367
R474 B.n409 B.n35 163.367
R475 B.n409 B.n408 163.367
R476 B.n408 B.n407 163.367
R477 B.n407 B.n37 163.367
R478 B.n402 B.n37 163.367
R479 B.n402 B.n401 163.367
R480 B.n401 B.n400 163.367
R481 B.n400 B.n41 163.367
R482 B.n396 B.n41 163.367
R483 B.n396 B.n395 163.367
R484 B.n395 B.n394 163.367
R485 B.n394 B.n43 163.367
R486 B.n390 B.n43 163.367
R487 B.n390 B.n389 163.367
R488 B.n389 B.n388 163.367
R489 B.n388 B.n45 163.367
R490 B.n384 B.n45 163.367
R491 B.n384 B.n383 163.367
R492 B.n383 B.n382 163.367
R493 B.n382 B.n47 163.367
R494 B.n378 B.n47 163.367
R495 B.n378 B.n377 163.367
R496 B.n377 B.n376 163.367
R497 B.n376 B.n49 163.367
R498 B.n372 B.n49 163.367
R499 B.n372 B.n371 163.367
R500 B.n371 B.n370 163.367
R501 B.n370 B.n51 163.367
R502 B.n366 B.n51 163.367
R503 B.n366 B.n365 163.367
R504 B.n365 B.n364 163.367
R505 B.n364 B.n53 163.367
R506 B.n360 B.n53 163.367
R507 B.n466 B.n15 163.367
R508 B.n467 B.n466 163.367
R509 B.n468 B.n467 163.367
R510 B.n468 B.n13 163.367
R511 B.n472 B.n13 163.367
R512 B.n473 B.n472 163.367
R513 B.n474 B.n473 163.367
R514 B.n474 B.n11 163.367
R515 B.n478 B.n11 163.367
R516 B.n479 B.n478 163.367
R517 B.n480 B.n479 163.367
R518 B.n480 B.n9 163.367
R519 B.n484 B.n9 163.367
R520 B.n485 B.n484 163.367
R521 B.n486 B.n485 163.367
R522 B.n486 B.n7 163.367
R523 B.n490 B.n7 163.367
R524 B.n491 B.n490 163.367
R525 B.n492 B.n491 163.367
R526 B.n492 B.n5 163.367
R527 B.n496 B.n5 163.367
R528 B.n497 B.n496 163.367
R529 B.n498 B.n497 163.367
R530 B.n498 B.n3 163.367
R531 B.n502 B.n3 163.367
R532 B.n503 B.n502 163.367
R533 B.n132 B.n2 163.367
R534 B.n133 B.n132 163.367
R535 B.n134 B.n133 163.367
R536 B.n134 B.n129 163.367
R537 B.n138 B.n129 163.367
R538 B.n139 B.n138 163.367
R539 B.n140 B.n139 163.367
R540 B.n140 B.n127 163.367
R541 B.n144 B.n127 163.367
R542 B.n145 B.n144 163.367
R543 B.n146 B.n145 163.367
R544 B.n146 B.n125 163.367
R545 B.n150 B.n125 163.367
R546 B.n151 B.n150 163.367
R547 B.n152 B.n151 163.367
R548 B.n152 B.n123 163.367
R549 B.n156 B.n123 163.367
R550 B.n157 B.n156 163.367
R551 B.n158 B.n157 163.367
R552 B.n158 B.n121 163.367
R553 B.n162 B.n121 163.367
R554 B.n163 B.n162 163.367
R555 B.n164 B.n163 163.367
R556 B.n164 B.n119 163.367
R557 B.n168 B.n119 163.367
R558 B.n169 B.n168 163.367
R559 B.n228 B.t7 156.621
R560 B.n38 B.t11 156.621
R561 B.n102 B.t1 156.613
R562 B.n30 B.t5 156.613
R563 B.n229 B.t8 113.76
R564 B.n39 B.t10 113.76
R565 B.n103 B.t2 113.752
R566 B.n31 B.t4 113.752
R567 B.n214 B.n103 59.5399
R568 B.n230 B.n229 59.5399
R569 B.n404 B.n39 59.5399
R570 B.n32 B.n31 59.5399
R571 B.n103 B.n102 42.8611
R572 B.n229 B.n228 42.8611
R573 B.n39 B.n38 42.8611
R574 B.n31 B.n30 42.8611
R575 B.n464 B.n463 32.0005
R576 B.n361 B.n54 32.0005
R577 B.n277 B.n82 32.0005
R578 B.n171 B.n118 32.0005
R579 B B.n505 18.0485
R580 B.n465 B.n464 10.6151
R581 B.n465 B.n14 10.6151
R582 B.n469 B.n14 10.6151
R583 B.n470 B.n469 10.6151
R584 B.n471 B.n470 10.6151
R585 B.n471 B.n12 10.6151
R586 B.n475 B.n12 10.6151
R587 B.n476 B.n475 10.6151
R588 B.n477 B.n476 10.6151
R589 B.n477 B.n10 10.6151
R590 B.n481 B.n10 10.6151
R591 B.n482 B.n481 10.6151
R592 B.n483 B.n482 10.6151
R593 B.n483 B.n8 10.6151
R594 B.n487 B.n8 10.6151
R595 B.n488 B.n487 10.6151
R596 B.n489 B.n488 10.6151
R597 B.n489 B.n6 10.6151
R598 B.n493 B.n6 10.6151
R599 B.n494 B.n493 10.6151
R600 B.n495 B.n494 10.6151
R601 B.n495 B.n4 10.6151
R602 B.n499 B.n4 10.6151
R603 B.n500 B.n499 10.6151
R604 B.n501 B.n500 10.6151
R605 B.n501 B.n0 10.6151
R606 B.n463 B.n16 10.6151
R607 B.n459 B.n16 10.6151
R608 B.n459 B.n458 10.6151
R609 B.n458 B.n457 10.6151
R610 B.n457 B.n18 10.6151
R611 B.n453 B.n18 10.6151
R612 B.n453 B.n452 10.6151
R613 B.n452 B.n451 10.6151
R614 B.n451 B.n20 10.6151
R615 B.n447 B.n20 10.6151
R616 B.n447 B.n446 10.6151
R617 B.n446 B.n445 10.6151
R618 B.n445 B.n22 10.6151
R619 B.n441 B.n22 10.6151
R620 B.n441 B.n440 10.6151
R621 B.n440 B.n439 10.6151
R622 B.n439 B.n24 10.6151
R623 B.n435 B.n24 10.6151
R624 B.n435 B.n434 10.6151
R625 B.n434 B.n433 10.6151
R626 B.n433 B.n26 10.6151
R627 B.n429 B.n26 10.6151
R628 B.n429 B.n428 10.6151
R629 B.n428 B.n427 10.6151
R630 B.n427 B.n28 10.6151
R631 B.n423 B.n28 10.6151
R632 B.n423 B.n422 10.6151
R633 B.n422 B.n421 10.6151
R634 B.n418 B.n417 10.6151
R635 B.n417 B.n416 10.6151
R636 B.n416 B.n34 10.6151
R637 B.n412 B.n34 10.6151
R638 B.n412 B.n411 10.6151
R639 B.n411 B.n410 10.6151
R640 B.n410 B.n36 10.6151
R641 B.n406 B.n36 10.6151
R642 B.n406 B.n405 10.6151
R643 B.n403 B.n40 10.6151
R644 B.n399 B.n40 10.6151
R645 B.n399 B.n398 10.6151
R646 B.n398 B.n397 10.6151
R647 B.n397 B.n42 10.6151
R648 B.n393 B.n42 10.6151
R649 B.n393 B.n392 10.6151
R650 B.n392 B.n391 10.6151
R651 B.n391 B.n44 10.6151
R652 B.n387 B.n44 10.6151
R653 B.n387 B.n386 10.6151
R654 B.n386 B.n385 10.6151
R655 B.n385 B.n46 10.6151
R656 B.n381 B.n46 10.6151
R657 B.n381 B.n380 10.6151
R658 B.n380 B.n379 10.6151
R659 B.n379 B.n48 10.6151
R660 B.n375 B.n48 10.6151
R661 B.n375 B.n374 10.6151
R662 B.n374 B.n373 10.6151
R663 B.n373 B.n50 10.6151
R664 B.n369 B.n50 10.6151
R665 B.n369 B.n368 10.6151
R666 B.n368 B.n367 10.6151
R667 B.n367 B.n52 10.6151
R668 B.n363 B.n52 10.6151
R669 B.n363 B.n362 10.6151
R670 B.n362 B.n361 10.6151
R671 B.n357 B.n54 10.6151
R672 B.n357 B.n356 10.6151
R673 B.n356 B.n355 10.6151
R674 B.n355 B.n56 10.6151
R675 B.n351 B.n56 10.6151
R676 B.n351 B.n350 10.6151
R677 B.n350 B.n349 10.6151
R678 B.n349 B.n58 10.6151
R679 B.n345 B.n58 10.6151
R680 B.n345 B.n344 10.6151
R681 B.n344 B.n343 10.6151
R682 B.n343 B.n60 10.6151
R683 B.n339 B.n60 10.6151
R684 B.n339 B.n338 10.6151
R685 B.n338 B.n337 10.6151
R686 B.n337 B.n62 10.6151
R687 B.n333 B.n62 10.6151
R688 B.n333 B.n332 10.6151
R689 B.n332 B.n331 10.6151
R690 B.n331 B.n64 10.6151
R691 B.n327 B.n64 10.6151
R692 B.n327 B.n326 10.6151
R693 B.n326 B.n325 10.6151
R694 B.n325 B.n66 10.6151
R695 B.n321 B.n66 10.6151
R696 B.n321 B.n320 10.6151
R697 B.n320 B.n319 10.6151
R698 B.n319 B.n68 10.6151
R699 B.n315 B.n68 10.6151
R700 B.n315 B.n314 10.6151
R701 B.n314 B.n313 10.6151
R702 B.n313 B.n70 10.6151
R703 B.n309 B.n70 10.6151
R704 B.n309 B.n308 10.6151
R705 B.n308 B.n307 10.6151
R706 B.n307 B.n72 10.6151
R707 B.n303 B.n72 10.6151
R708 B.n303 B.n302 10.6151
R709 B.n302 B.n301 10.6151
R710 B.n301 B.n74 10.6151
R711 B.n297 B.n74 10.6151
R712 B.n297 B.n296 10.6151
R713 B.n296 B.n295 10.6151
R714 B.n295 B.n76 10.6151
R715 B.n291 B.n76 10.6151
R716 B.n291 B.n290 10.6151
R717 B.n290 B.n289 10.6151
R718 B.n289 B.n78 10.6151
R719 B.n285 B.n78 10.6151
R720 B.n285 B.n284 10.6151
R721 B.n284 B.n283 10.6151
R722 B.n283 B.n80 10.6151
R723 B.n279 B.n80 10.6151
R724 B.n279 B.n278 10.6151
R725 B.n278 B.n277 10.6151
R726 B.n131 B.n1 10.6151
R727 B.n131 B.n130 10.6151
R728 B.n135 B.n130 10.6151
R729 B.n136 B.n135 10.6151
R730 B.n137 B.n136 10.6151
R731 B.n137 B.n128 10.6151
R732 B.n141 B.n128 10.6151
R733 B.n142 B.n141 10.6151
R734 B.n143 B.n142 10.6151
R735 B.n143 B.n126 10.6151
R736 B.n147 B.n126 10.6151
R737 B.n148 B.n147 10.6151
R738 B.n149 B.n148 10.6151
R739 B.n149 B.n124 10.6151
R740 B.n153 B.n124 10.6151
R741 B.n154 B.n153 10.6151
R742 B.n155 B.n154 10.6151
R743 B.n155 B.n122 10.6151
R744 B.n159 B.n122 10.6151
R745 B.n160 B.n159 10.6151
R746 B.n161 B.n160 10.6151
R747 B.n161 B.n120 10.6151
R748 B.n165 B.n120 10.6151
R749 B.n166 B.n165 10.6151
R750 B.n167 B.n166 10.6151
R751 B.n167 B.n118 10.6151
R752 B.n172 B.n171 10.6151
R753 B.n173 B.n172 10.6151
R754 B.n173 B.n116 10.6151
R755 B.n177 B.n116 10.6151
R756 B.n178 B.n177 10.6151
R757 B.n179 B.n178 10.6151
R758 B.n179 B.n114 10.6151
R759 B.n183 B.n114 10.6151
R760 B.n184 B.n183 10.6151
R761 B.n185 B.n184 10.6151
R762 B.n185 B.n112 10.6151
R763 B.n189 B.n112 10.6151
R764 B.n190 B.n189 10.6151
R765 B.n191 B.n190 10.6151
R766 B.n191 B.n110 10.6151
R767 B.n195 B.n110 10.6151
R768 B.n196 B.n195 10.6151
R769 B.n197 B.n196 10.6151
R770 B.n197 B.n108 10.6151
R771 B.n201 B.n108 10.6151
R772 B.n202 B.n201 10.6151
R773 B.n203 B.n202 10.6151
R774 B.n203 B.n106 10.6151
R775 B.n207 B.n106 10.6151
R776 B.n208 B.n207 10.6151
R777 B.n209 B.n208 10.6151
R778 B.n209 B.n104 10.6151
R779 B.n213 B.n104 10.6151
R780 B.n216 B.n215 10.6151
R781 B.n216 B.n100 10.6151
R782 B.n220 B.n100 10.6151
R783 B.n221 B.n220 10.6151
R784 B.n222 B.n221 10.6151
R785 B.n222 B.n98 10.6151
R786 B.n226 B.n98 10.6151
R787 B.n227 B.n226 10.6151
R788 B.n231 B.n227 10.6151
R789 B.n235 B.n96 10.6151
R790 B.n236 B.n235 10.6151
R791 B.n237 B.n236 10.6151
R792 B.n237 B.n94 10.6151
R793 B.n241 B.n94 10.6151
R794 B.n242 B.n241 10.6151
R795 B.n243 B.n242 10.6151
R796 B.n243 B.n92 10.6151
R797 B.n247 B.n92 10.6151
R798 B.n248 B.n247 10.6151
R799 B.n249 B.n248 10.6151
R800 B.n249 B.n90 10.6151
R801 B.n253 B.n90 10.6151
R802 B.n254 B.n253 10.6151
R803 B.n255 B.n254 10.6151
R804 B.n255 B.n88 10.6151
R805 B.n259 B.n88 10.6151
R806 B.n260 B.n259 10.6151
R807 B.n261 B.n260 10.6151
R808 B.n261 B.n86 10.6151
R809 B.n265 B.n86 10.6151
R810 B.n266 B.n265 10.6151
R811 B.n267 B.n266 10.6151
R812 B.n267 B.n84 10.6151
R813 B.n271 B.n84 10.6151
R814 B.n272 B.n271 10.6151
R815 B.n273 B.n272 10.6151
R816 B.n273 B.n82 10.6151
R817 B.n421 B.n32 9.36635
R818 B.n404 B.n403 9.36635
R819 B.n214 B.n213 9.36635
R820 B.n230 B.n96 9.36635
R821 B.n505 B.n0 8.11757
R822 B.n505 B.n1 8.11757
R823 B.n418 B.n32 1.24928
R824 B.n405 B.n404 1.24928
R825 B.n215 B.n214 1.24928
R826 B.n231 B.n230 1.24928
C0 w_n2296_n2514# VDD2 1.23504f
C1 VP VDD1 3.17232f
C2 VTAIL VP 2.97322f
C3 B VDD1 1.02054f
C4 VN VDD2 2.97273f
C5 VTAIL B 3.2602f
C6 w_n2296_n2514# VP 3.96355f
C7 VTAIL VDD1 4.23787f
C8 w_n2296_n2514# B 7.16271f
C9 w_n2296_n2514# VDD1 1.19502f
C10 VN VP 4.87826f
C11 VP VDD2 0.348313f
C12 VTAIL w_n2296_n2514# 2.98727f
C13 VN B 0.921985f
C14 B VDD2 1.06091f
C15 VN VDD1 0.148172f
C16 VDD2 VDD1 0.851707f
C17 VN VTAIL 2.95911f
C18 VTAIL VDD2 4.28725f
C19 VN w_n2296_n2514# 3.67021f
C20 B VP 1.40542f
C21 VDD2 VSUBS 0.730094f
C22 VDD1 VSUBS 4.761006f
C23 VTAIL VSUBS 0.920597f
C24 VN VSUBS 5.07781f
C25 VP VSUBS 1.736259f
C26 B VSUBS 3.291262f
C27 w_n2296_n2514# VSUBS 71.662704f
C28 B.n0 VSUBS 0.007127f
C29 B.n1 VSUBS 0.007127f
C30 B.n2 VSUBS 0.01054f
C31 B.n3 VSUBS 0.008077f
C32 B.n4 VSUBS 0.008077f
C33 B.n5 VSUBS 0.008077f
C34 B.n6 VSUBS 0.008077f
C35 B.n7 VSUBS 0.008077f
C36 B.n8 VSUBS 0.008077f
C37 B.n9 VSUBS 0.008077f
C38 B.n10 VSUBS 0.008077f
C39 B.n11 VSUBS 0.008077f
C40 B.n12 VSUBS 0.008077f
C41 B.n13 VSUBS 0.008077f
C42 B.n14 VSUBS 0.008077f
C43 B.n15 VSUBS 0.017971f
C44 B.n16 VSUBS 0.008077f
C45 B.n17 VSUBS 0.008077f
C46 B.n18 VSUBS 0.008077f
C47 B.n19 VSUBS 0.008077f
C48 B.n20 VSUBS 0.008077f
C49 B.n21 VSUBS 0.008077f
C50 B.n22 VSUBS 0.008077f
C51 B.n23 VSUBS 0.008077f
C52 B.n24 VSUBS 0.008077f
C53 B.n25 VSUBS 0.008077f
C54 B.n26 VSUBS 0.008077f
C55 B.n27 VSUBS 0.008077f
C56 B.n28 VSUBS 0.008077f
C57 B.n29 VSUBS 0.008077f
C58 B.t4 VSUBS 0.273549f
C59 B.t5 VSUBS 0.292f
C60 B.t3 VSUBS 0.767767f
C61 B.n30 VSUBS 0.150641f
C62 B.n31 VSUBS 0.078939f
C63 B.n32 VSUBS 0.018713f
C64 B.n33 VSUBS 0.008077f
C65 B.n34 VSUBS 0.008077f
C66 B.n35 VSUBS 0.008077f
C67 B.n36 VSUBS 0.008077f
C68 B.n37 VSUBS 0.008077f
C69 B.t10 VSUBS 0.273547f
C70 B.t11 VSUBS 0.291998f
C71 B.t9 VSUBS 0.767767f
C72 B.n38 VSUBS 0.150644f
C73 B.n39 VSUBS 0.07894f
C74 B.n40 VSUBS 0.008077f
C75 B.n41 VSUBS 0.008077f
C76 B.n42 VSUBS 0.008077f
C77 B.n43 VSUBS 0.008077f
C78 B.n44 VSUBS 0.008077f
C79 B.n45 VSUBS 0.008077f
C80 B.n46 VSUBS 0.008077f
C81 B.n47 VSUBS 0.008077f
C82 B.n48 VSUBS 0.008077f
C83 B.n49 VSUBS 0.008077f
C84 B.n50 VSUBS 0.008077f
C85 B.n51 VSUBS 0.008077f
C86 B.n52 VSUBS 0.008077f
C87 B.n53 VSUBS 0.008077f
C88 B.n54 VSUBS 0.017971f
C89 B.n55 VSUBS 0.008077f
C90 B.n56 VSUBS 0.008077f
C91 B.n57 VSUBS 0.008077f
C92 B.n58 VSUBS 0.008077f
C93 B.n59 VSUBS 0.008077f
C94 B.n60 VSUBS 0.008077f
C95 B.n61 VSUBS 0.008077f
C96 B.n62 VSUBS 0.008077f
C97 B.n63 VSUBS 0.008077f
C98 B.n64 VSUBS 0.008077f
C99 B.n65 VSUBS 0.008077f
C100 B.n66 VSUBS 0.008077f
C101 B.n67 VSUBS 0.008077f
C102 B.n68 VSUBS 0.008077f
C103 B.n69 VSUBS 0.008077f
C104 B.n70 VSUBS 0.008077f
C105 B.n71 VSUBS 0.008077f
C106 B.n72 VSUBS 0.008077f
C107 B.n73 VSUBS 0.008077f
C108 B.n74 VSUBS 0.008077f
C109 B.n75 VSUBS 0.008077f
C110 B.n76 VSUBS 0.008077f
C111 B.n77 VSUBS 0.008077f
C112 B.n78 VSUBS 0.008077f
C113 B.n79 VSUBS 0.008077f
C114 B.n80 VSUBS 0.008077f
C115 B.n81 VSUBS 0.008077f
C116 B.n82 VSUBS 0.018351f
C117 B.n83 VSUBS 0.008077f
C118 B.n84 VSUBS 0.008077f
C119 B.n85 VSUBS 0.008077f
C120 B.n86 VSUBS 0.008077f
C121 B.n87 VSUBS 0.008077f
C122 B.n88 VSUBS 0.008077f
C123 B.n89 VSUBS 0.008077f
C124 B.n90 VSUBS 0.008077f
C125 B.n91 VSUBS 0.008077f
C126 B.n92 VSUBS 0.008077f
C127 B.n93 VSUBS 0.008077f
C128 B.n94 VSUBS 0.008077f
C129 B.n95 VSUBS 0.008077f
C130 B.n96 VSUBS 0.007602f
C131 B.n97 VSUBS 0.008077f
C132 B.n98 VSUBS 0.008077f
C133 B.n99 VSUBS 0.008077f
C134 B.n100 VSUBS 0.008077f
C135 B.n101 VSUBS 0.008077f
C136 B.t2 VSUBS 0.273549f
C137 B.t1 VSUBS 0.292f
C138 B.t0 VSUBS 0.767767f
C139 B.n102 VSUBS 0.150641f
C140 B.n103 VSUBS 0.078939f
C141 B.n104 VSUBS 0.008077f
C142 B.n105 VSUBS 0.008077f
C143 B.n106 VSUBS 0.008077f
C144 B.n107 VSUBS 0.008077f
C145 B.n108 VSUBS 0.008077f
C146 B.n109 VSUBS 0.008077f
C147 B.n110 VSUBS 0.008077f
C148 B.n111 VSUBS 0.008077f
C149 B.n112 VSUBS 0.008077f
C150 B.n113 VSUBS 0.008077f
C151 B.n114 VSUBS 0.008077f
C152 B.n115 VSUBS 0.008077f
C153 B.n116 VSUBS 0.008077f
C154 B.n117 VSUBS 0.008077f
C155 B.n118 VSUBS 0.017971f
C156 B.n119 VSUBS 0.008077f
C157 B.n120 VSUBS 0.008077f
C158 B.n121 VSUBS 0.008077f
C159 B.n122 VSUBS 0.008077f
C160 B.n123 VSUBS 0.008077f
C161 B.n124 VSUBS 0.008077f
C162 B.n125 VSUBS 0.008077f
C163 B.n126 VSUBS 0.008077f
C164 B.n127 VSUBS 0.008077f
C165 B.n128 VSUBS 0.008077f
C166 B.n129 VSUBS 0.008077f
C167 B.n130 VSUBS 0.008077f
C168 B.n131 VSUBS 0.008077f
C169 B.n132 VSUBS 0.008077f
C170 B.n133 VSUBS 0.008077f
C171 B.n134 VSUBS 0.008077f
C172 B.n135 VSUBS 0.008077f
C173 B.n136 VSUBS 0.008077f
C174 B.n137 VSUBS 0.008077f
C175 B.n138 VSUBS 0.008077f
C176 B.n139 VSUBS 0.008077f
C177 B.n140 VSUBS 0.008077f
C178 B.n141 VSUBS 0.008077f
C179 B.n142 VSUBS 0.008077f
C180 B.n143 VSUBS 0.008077f
C181 B.n144 VSUBS 0.008077f
C182 B.n145 VSUBS 0.008077f
C183 B.n146 VSUBS 0.008077f
C184 B.n147 VSUBS 0.008077f
C185 B.n148 VSUBS 0.008077f
C186 B.n149 VSUBS 0.008077f
C187 B.n150 VSUBS 0.008077f
C188 B.n151 VSUBS 0.008077f
C189 B.n152 VSUBS 0.008077f
C190 B.n153 VSUBS 0.008077f
C191 B.n154 VSUBS 0.008077f
C192 B.n155 VSUBS 0.008077f
C193 B.n156 VSUBS 0.008077f
C194 B.n157 VSUBS 0.008077f
C195 B.n158 VSUBS 0.008077f
C196 B.n159 VSUBS 0.008077f
C197 B.n160 VSUBS 0.008077f
C198 B.n161 VSUBS 0.008077f
C199 B.n162 VSUBS 0.008077f
C200 B.n163 VSUBS 0.008077f
C201 B.n164 VSUBS 0.008077f
C202 B.n165 VSUBS 0.008077f
C203 B.n166 VSUBS 0.008077f
C204 B.n167 VSUBS 0.008077f
C205 B.n168 VSUBS 0.008077f
C206 B.n169 VSUBS 0.017971f
C207 B.n170 VSUBS 0.019325f
C208 B.n171 VSUBS 0.019325f
C209 B.n172 VSUBS 0.008077f
C210 B.n173 VSUBS 0.008077f
C211 B.n174 VSUBS 0.008077f
C212 B.n175 VSUBS 0.008077f
C213 B.n176 VSUBS 0.008077f
C214 B.n177 VSUBS 0.008077f
C215 B.n178 VSUBS 0.008077f
C216 B.n179 VSUBS 0.008077f
C217 B.n180 VSUBS 0.008077f
C218 B.n181 VSUBS 0.008077f
C219 B.n182 VSUBS 0.008077f
C220 B.n183 VSUBS 0.008077f
C221 B.n184 VSUBS 0.008077f
C222 B.n185 VSUBS 0.008077f
C223 B.n186 VSUBS 0.008077f
C224 B.n187 VSUBS 0.008077f
C225 B.n188 VSUBS 0.008077f
C226 B.n189 VSUBS 0.008077f
C227 B.n190 VSUBS 0.008077f
C228 B.n191 VSUBS 0.008077f
C229 B.n192 VSUBS 0.008077f
C230 B.n193 VSUBS 0.008077f
C231 B.n194 VSUBS 0.008077f
C232 B.n195 VSUBS 0.008077f
C233 B.n196 VSUBS 0.008077f
C234 B.n197 VSUBS 0.008077f
C235 B.n198 VSUBS 0.008077f
C236 B.n199 VSUBS 0.008077f
C237 B.n200 VSUBS 0.008077f
C238 B.n201 VSUBS 0.008077f
C239 B.n202 VSUBS 0.008077f
C240 B.n203 VSUBS 0.008077f
C241 B.n204 VSUBS 0.008077f
C242 B.n205 VSUBS 0.008077f
C243 B.n206 VSUBS 0.008077f
C244 B.n207 VSUBS 0.008077f
C245 B.n208 VSUBS 0.008077f
C246 B.n209 VSUBS 0.008077f
C247 B.n210 VSUBS 0.008077f
C248 B.n211 VSUBS 0.008077f
C249 B.n212 VSUBS 0.008077f
C250 B.n213 VSUBS 0.007602f
C251 B.n214 VSUBS 0.018713f
C252 B.n215 VSUBS 0.004514f
C253 B.n216 VSUBS 0.008077f
C254 B.n217 VSUBS 0.008077f
C255 B.n218 VSUBS 0.008077f
C256 B.n219 VSUBS 0.008077f
C257 B.n220 VSUBS 0.008077f
C258 B.n221 VSUBS 0.008077f
C259 B.n222 VSUBS 0.008077f
C260 B.n223 VSUBS 0.008077f
C261 B.n224 VSUBS 0.008077f
C262 B.n225 VSUBS 0.008077f
C263 B.n226 VSUBS 0.008077f
C264 B.n227 VSUBS 0.008077f
C265 B.t8 VSUBS 0.273547f
C266 B.t7 VSUBS 0.291998f
C267 B.t6 VSUBS 0.767767f
C268 B.n228 VSUBS 0.150644f
C269 B.n229 VSUBS 0.07894f
C270 B.n230 VSUBS 0.018713f
C271 B.n231 VSUBS 0.004514f
C272 B.n232 VSUBS 0.008077f
C273 B.n233 VSUBS 0.008077f
C274 B.n234 VSUBS 0.008077f
C275 B.n235 VSUBS 0.008077f
C276 B.n236 VSUBS 0.008077f
C277 B.n237 VSUBS 0.008077f
C278 B.n238 VSUBS 0.008077f
C279 B.n239 VSUBS 0.008077f
C280 B.n240 VSUBS 0.008077f
C281 B.n241 VSUBS 0.008077f
C282 B.n242 VSUBS 0.008077f
C283 B.n243 VSUBS 0.008077f
C284 B.n244 VSUBS 0.008077f
C285 B.n245 VSUBS 0.008077f
C286 B.n246 VSUBS 0.008077f
C287 B.n247 VSUBS 0.008077f
C288 B.n248 VSUBS 0.008077f
C289 B.n249 VSUBS 0.008077f
C290 B.n250 VSUBS 0.008077f
C291 B.n251 VSUBS 0.008077f
C292 B.n252 VSUBS 0.008077f
C293 B.n253 VSUBS 0.008077f
C294 B.n254 VSUBS 0.008077f
C295 B.n255 VSUBS 0.008077f
C296 B.n256 VSUBS 0.008077f
C297 B.n257 VSUBS 0.008077f
C298 B.n258 VSUBS 0.008077f
C299 B.n259 VSUBS 0.008077f
C300 B.n260 VSUBS 0.008077f
C301 B.n261 VSUBS 0.008077f
C302 B.n262 VSUBS 0.008077f
C303 B.n263 VSUBS 0.008077f
C304 B.n264 VSUBS 0.008077f
C305 B.n265 VSUBS 0.008077f
C306 B.n266 VSUBS 0.008077f
C307 B.n267 VSUBS 0.008077f
C308 B.n268 VSUBS 0.008077f
C309 B.n269 VSUBS 0.008077f
C310 B.n270 VSUBS 0.008077f
C311 B.n271 VSUBS 0.008077f
C312 B.n272 VSUBS 0.008077f
C313 B.n273 VSUBS 0.008077f
C314 B.n274 VSUBS 0.008077f
C315 B.n275 VSUBS 0.019325f
C316 B.n276 VSUBS 0.017971f
C317 B.n277 VSUBS 0.018945f
C318 B.n278 VSUBS 0.008077f
C319 B.n279 VSUBS 0.008077f
C320 B.n280 VSUBS 0.008077f
C321 B.n281 VSUBS 0.008077f
C322 B.n282 VSUBS 0.008077f
C323 B.n283 VSUBS 0.008077f
C324 B.n284 VSUBS 0.008077f
C325 B.n285 VSUBS 0.008077f
C326 B.n286 VSUBS 0.008077f
C327 B.n287 VSUBS 0.008077f
C328 B.n288 VSUBS 0.008077f
C329 B.n289 VSUBS 0.008077f
C330 B.n290 VSUBS 0.008077f
C331 B.n291 VSUBS 0.008077f
C332 B.n292 VSUBS 0.008077f
C333 B.n293 VSUBS 0.008077f
C334 B.n294 VSUBS 0.008077f
C335 B.n295 VSUBS 0.008077f
C336 B.n296 VSUBS 0.008077f
C337 B.n297 VSUBS 0.008077f
C338 B.n298 VSUBS 0.008077f
C339 B.n299 VSUBS 0.008077f
C340 B.n300 VSUBS 0.008077f
C341 B.n301 VSUBS 0.008077f
C342 B.n302 VSUBS 0.008077f
C343 B.n303 VSUBS 0.008077f
C344 B.n304 VSUBS 0.008077f
C345 B.n305 VSUBS 0.008077f
C346 B.n306 VSUBS 0.008077f
C347 B.n307 VSUBS 0.008077f
C348 B.n308 VSUBS 0.008077f
C349 B.n309 VSUBS 0.008077f
C350 B.n310 VSUBS 0.008077f
C351 B.n311 VSUBS 0.008077f
C352 B.n312 VSUBS 0.008077f
C353 B.n313 VSUBS 0.008077f
C354 B.n314 VSUBS 0.008077f
C355 B.n315 VSUBS 0.008077f
C356 B.n316 VSUBS 0.008077f
C357 B.n317 VSUBS 0.008077f
C358 B.n318 VSUBS 0.008077f
C359 B.n319 VSUBS 0.008077f
C360 B.n320 VSUBS 0.008077f
C361 B.n321 VSUBS 0.008077f
C362 B.n322 VSUBS 0.008077f
C363 B.n323 VSUBS 0.008077f
C364 B.n324 VSUBS 0.008077f
C365 B.n325 VSUBS 0.008077f
C366 B.n326 VSUBS 0.008077f
C367 B.n327 VSUBS 0.008077f
C368 B.n328 VSUBS 0.008077f
C369 B.n329 VSUBS 0.008077f
C370 B.n330 VSUBS 0.008077f
C371 B.n331 VSUBS 0.008077f
C372 B.n332 VSUBS 0.008077f
C373 B.n333 VSUBS 0.008077f
C374 B.n334 VSUBS 0.008077f
C375 B.n335 VSUBS 0.008077f
C376 B.n336 VSUBS 0.008077f
C377 B.n337 VSUBS 0.008077f
C378 B.n338 VSUBS 0.008077f
C379 B.n339 VSUBS 0.008077f
C380 B.n340 VSUBS 0.008077f
C381 B.n341 VSUBS 0.008077f
C382 B.n342 VSUBS 0.008077f
C383 B.n343 VSUBS 0.008077f
C384 B.n344 VSUBS 0.008077f
C385 B.n345 VSUBS 0.008077f
C386 B.n346 VSUBS 0.008077f
C387 B.n347 VSUBS 0.008077f
C388 B.n348 VSUBS 0.008077f
C389 B.n349 VSUBS 0.008077f
C390 B.n350 VSUBS 0.008077f
C391 B.n351 VSUBS 0.008077f
C392 B.n352 VSUBS 0.008077f
C393 B.n353 VSUBS 0.008077f
C394 B.n354 VSUBS 0.008077f
C395 B.n355 VSUBS 0.008077f
C396 B.n356 VSUBS 0.008077f
C397 B.n357 VSUBS 0.008077f
C398 B.n358 VSUBS 0.008077f
C399 B.n359 VSUBS 0.017971f
C400 B.n360 VSUBS 0.019325f
C401 B.n361 VSUBS 0.019325f
C402 B.n362 VSUBS 0.008077f
C403 B.n363 VSUBS 0.008077f
C404 B.n364 VSUBS 0.008077f
C405 B.n365 VSUBS 0.008077f
C406 B.n366 VSUBS 0.008077f
C407 B.n367 VSUBS 0.008077f
C408 B.n368 VSUBS 0.008077f
C409 B.n369 VSUBS 0.008077f
C410 B.n370 VSUBS 0.008077f
C411 B.n371 VSUBS 0.008077f
C412 B.n372 VSUBS 0.008077f
C413 B.n373 VSUBS 0.008077f
C414 B.n374 VSUBS 0.008077f
C415 B.n375 VSUBS 0.008077f
C416 B.n376 VSUBS 0.008077f
C417 B.n377 VSUBS 0.008077f
C418 B.n378 VSUBS 0.008077f
C419 B.n379 VSUBS 0.008077f
C420 B.n380 VSUBS 0.008077f
C421 B.n381 VSUBS 0.008077f
C422 B.n382 VSUBS 0.008077f
C423 B.n383 VSUBS 0.008077f
C424 B.n384 VSUBS 0.008077f
C425 B.n385 VSUBS 0.008077f
C426 B.n386 VSUBS 0.008077f
C427 B.n387 VSUBS 0.008077f
C428 B.n388 VSUBS 0.008077f
C429 B.n389 VSUBS 0.008077f
C430 B.n390 VSUBS 0.008077f
C431 B.n391 VSUBS 0.008077f
C432 B.n392 VSUBS 0.008077f
C433 B.n393 VSUBS 0.008077f
C434 B.n394 VSUBS 0.008077f
C435 B.n395 VSUBS 0.008077f
C436 B.n396 VSUBS 0.008077f
C437 B.n397 VSUBS 0.008077f
C438 B.n398 VSUBS 0.008077f
C439 B.n399 VSUBS 0.008077f
C440 B.n400 VSUBS 0.008077f
C441 B.n401 VSUBS 0.008077f
C442 B.n402 VSUBS 0.008077f
C443 B.n403 VSUBS 0.007602f
C444 B.n404 VSUBS 0.018713f
C445 B.n405 VSUBS 0.004514f
C446 B.n406 VSUBS 0.008077f
C447 B.n407 VSUBS 0.008077f
C448 B.n408 VSUBS 0.008077f
C449 B.n409 VSUBS 0.008077f
C450 B.n410 VSUBS 0.008077f
C451 B.n411 VSUBS 0.008077f
C452 B.n412 VSUBS 0.008077f
C453 B.n413 VSUBS 0.008077f
C454 B.n414 VSUBS 0.008077f
C455 B.n415 VSUBS 0.008077f
C456 B.n416 VSUBS 0.008077f
C457 B.n417 VSUBS 0.008077f
C458 B.n418 VSUBS 0.004514f
C459 B.n419 VSUBS 0.008077f
C460 B.n420 VSUBS 0.008077f
C461 B.n421 VSUBS 0.007602f
C462 B.n422 VSUBS 0.008077f
C463 B.n423 VSUBS 0.008077f
C464 B.n424 VSUBS 0.008077f
C465 B.n425 VSUBS 0.008077f
C466 B.n426 VSUBS 0.008077f
C467 B.n427 VSUBS 0.008077f
C468 B.n428 VSUBS 0.008077f
C469 B.n429 VSUBS 0.008077f
C470 B.n430 VSUBS 0.008077f
C471 B.n431 VSUBS 0.008077f
C472 B.n432 VSUBS 0.008077f
C473 B.n433 VSUBS 0.008077f
C474 B.n434 VSUBS 0.008077f
C475 B.n435 VSUBS 0.008077f
C476 B.n436 VSUBS 0.008077f
C477 B.n437 VSUBS 0.008077f
C478 B.n438 VSUBS 0.008077f
C479 B.n439 VSUBS 0.008077f
C480 B.n440 VSUBS 0.008077f
C481 B.n441 VSUBS 0.008077f
C482 B.n442 VSUBS 0.008077f
C483 B.n443 VSUBS 0.008077f
C484 B.n444 VSUBS 0.008077f
C485 B.n445 VSUBS 0.008077f
C486 B.n446 VSUBS 0.008077f
C487 B.n447 VSUBS 0.008077f
C488 B.n448 VSUBS 0.008077f
C489 B.n449 VSUBS 0.008077f
C490 B.n450 VSUBS 0.008077f
C491 B.n451 VSUBS 0.008077f
C492 B.n452 VSUBS 0.008077f
C493 B.n453 VSUBS 0.008077f
C494 B.n454 VSUBS 0.008077f
C495 B.n455 VSUBS 0.008077f
C496 B.n456 VSUBS 0.008077f
C497 B.n457 VSUBS 0.008077f
C498 B.n458 VSUBS 0.008077f
C499 B.n459 VSUBS 0.008077f
C500 B.n460 VSUBS 0.008077f
C501 B.n461 VSUBS 0.008077f
C502 B.n462 VSUBS 0.019325f
C503 B.n463 VSUBS 0.019325f
C504 B.n464 VSUBS 0.017971f
C505 B.n465 VSUBS 0.008077f
C506 B.n466 VSUBS 0.008077f
C507 B.n467 VSUBS 0.008077f
C508 B.n468 VSUBS 0.008077f
C509 B.n469 VSUBS 0.008077f
C510 B.n470 VSUBS 0.008077f
C511 B.n471 VSUBS 0.008077f
C512 B.n472 VSUBS 0.008077f
C513 B.n473 VSUBS 0.008077f
C514 B.n474 VSUBS 0.008077f
C515 B.n475 VSUBS 0.008077f
C516 B.n476 VSUBS 0.008077f
C517 B.n477 VSUBS 0.008077f
C518 B.n478 VSUBS 0.008077f
C519 B.n479 VSUBS 0.008077f
C520 B.n480 VSUBS 0.008077f
C521 B.n481 VSUBS 0.008077f
C522 B.n482 VSUBS 0.008077f
C523 B.n483 VSUBS 0.008077f
C524 B.n484 VSUBS 0.008077f
C525 B.n485 VSUBS 0.008077f
C526 B.n486 VSUBS 0.008077f
C527 B.n487 VSUBS 0.008077f
C528 B.n488 VSUBS 0.008077f
C529 B.n489 VSUBS 0.008077f
C530 B.n490 VSUBS 0.008077f
C531 B.n491 VSUBS 0.008077f
C532 B.n492 VSUBS 0.008077f
C533 B.n493 VSUBS 0.008077f
C534 B.n494 VSUBS 0.008077f
C535 B.n495 VSUBS 0.008077f
C536 B.n496 VSUBS 0.008077f
C537 B.n497 VSUBS 0.008077f
C538 B.n498 VSUBS 0.008077f
C539 B.n499 VSUBS 0.008077f
C540 B.n500 VSUBS 0.008077f
C541 B.n501 VSUBS 0.008077f
C542 B.n502 VSUBS 0.008077f
C543 B.n503 VSUBS 0.01054f
C544 B.n504 VSUBS 0.011228f
C545 B.n505 VSUBS 0.022327f
C546 VDD2.t3 VSUBS 0.165729f
C547 VDD2.t2 VSUBS 0.165729f
C548 VDD2.n0 VSUBS 1.65944f
C549 VDD2.t0 VSUBS 0.165729f
C550 VDD2.t1 VSUBS 0.165729f
C551 VDD2.n1 VSUBS 1.16901f
C552 VDD2.n2 VSUBS 3.63624f
C553 VN.t0 VSUBS 1.94554f
C554 VN.t1 VSUBS 1.94283f
C555 VN.n0 VSUBS 1.33742f
C556 VN.t2 VSUBS 1.94554f
C557 VN.t3 VSUBS 1.94283f
C558 VN.n1 VSUBS 3.02005f
C559 VDD1.t0 VSUBS 0.165724f
C560 VDD1.t3 VSUBS 0.165724f
C561 VDD1.n0 VSUBS 1.16944f
C562 VDD1.t1 VSUBS 0.165724f
C563 VDD1.t2 VSUBS 0.165724f
C564 VDD1.n1 VSUBS 1.68117f
C565 VTAIL.t2 VSUBS 1.31675f
C566 VTAIL.n0 VSUBS 0.712234f
C567 VTAIL.t4 VSUBS 1.31675f
C568 VTAIL.n1 VSUBS 0.784658f
C569 VTAIL.t5 VSUBS 1.31675f
C570 VTAIL.n2 VSUBS 1.78185f
C571 VTAIL.t0 VSUBS 1.31675f
C572 VTAIL.n3 VSUBS 1.78184f
C573 VTAIL.t1 VSUBS 1.31675f
C574 VTAIL.n4 VSUBS 0.78465f
C575 VTAIL.t6 VSUBS 1.31675f
C576 VTAIL.n5 VSUBS 0.78465f
C577 VTAIL.t7 VSUBS 1.31675f
C578 VTAIL.n6 VSUBS 1.78184f
C579 VTAIL.t3 VSUBS 1.31675f
C580 VTAIL.n7 VSUBS 1.7f
C581 VP.n0 VSUBS 0.045548f
C582 VP.t1 VSUBS 1.77503f
C583 VP.n1 VSUBS 0.036822f
C584 VP.n2 VSUBS 0.045548f
C585 VP.t2 VSUBS 1.77503f
C586 VP.t3 VSUBS 2.0207f
C587 VP.t0 VSUBS 2.01788f
C588 VP.n3 VSUBS 3.10928f
C589 VP.n4 VSUBS 2.23263f
C590 VP.n5 VSUBS 0.772357f
C591 VP.n6 VSUBS 0.051779f
C592 VP.n7 VSUBS 0.090527f
C593 VP.n8 VSUBS 0.045548f
C594 VP.n9 VSUBS 0.045548f
C595 VP.n10 VSUBS 0.045548f
C596 VP.n11 VSUBS 0.090527f
C597 VP.n12 VSUBS 0.051779f
C598 VP.n13 VSUBS 0.772357f
C599 VP.n14 VSUBS 0.048732f
.ends

