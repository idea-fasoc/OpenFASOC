* NGSPICE file created from diff_pair_sample_0585.ext - technology: sky130A

.subckt diff_pair_sample_0585 VTAIL VN VP B VDD2 VDD1
X0 B.t18 B.t16 B.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=5.3625 pd=28.28 as=0 ps=0 w=13.75 l=0.32
X1 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=5.3625 pd=28.28 as=0 ps=0 w=13.75 l=0.32
X2 VDD2.t5 VN.t0 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=5.3625 pd=28.28 as=2.26875 ps=14.08 w=13.75 l=0.32
X3 VDD1.t5 VP.t0 VTAIL.t5 B.t19 sky130_fd_pr__nfet_01v8 ad=2.26875 pd=14.08 as=5.3625 ps=28.28 w=13.75 l=0.32
X4 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=5.3625 pd=28.28 as=0 ps=0 w=13.75 l=0.32
X5 VTAIL.t8 VN.t1 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.26875 pd=14.08 as=2.26875 ps=14.08 w=13.75 l=0.32
X6 VTAIL.t4 VP.t1 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.26875 pd=14.08 as=2.26875 ps=14.08 w=13.75 l=0.32
X7 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=5.3625 pd=28.28 as=0 ps=0 w=13.75 l=0.32
X8 VDD2.t3 VN.t2 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.26875 pd=14.08 as=5.3625 ps=28.28 w=13.75 l=0.32
X9 VTAIL.t9 VN.t3 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.26875 pd=14.08 as=2.26875 ps=14.08 w=13.75 l=0.32
X10 VDD2.t1 VN.t4 VTAIL.t10 B.t19 sky130_fd_pr__nfet_01v8 ad=2.26875 pd=14.08 as=5.3625 ps=28.28 w=13.75 l=0.32
X11 VDD2.t0 VN.t5 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=5.3625 pd=28.28 as=2.26875 ps=14.08 w=13.75 l=0.32
X12 VDD1.t3 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.26875 pd=14.08 as=5.3625 ps=28.28 w=13.75 l=0.32
X13 VTAIL.t0 VP.t3 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.26875 pd=14.08 as=2.26875 ps=14.08 w=13.75 l=0.32
X14 VDD1.t1 VP.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=5.3625 pd=28.28 as=2.26875 ps=14.08 w=13.75 l=0.32
X15 VDD1.t0 VP.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.3625 pd=28.28 as=2.26875 ps=14.08 w=13.75 l=0.32
R0 B.n87 B.t5 1249.3
R1 B.n84 B.t16 1249.3
R2 B.n371 B.t13 1249.3
R3 B.n368 B.t9 1249.3
R4 B.n647 B.n646 585
R5 B.n648 B.n647 585
R6 B.n288 B.n82 585
R7 B.n287 B.n286 585
R8 B.n285 B.n284 585
R9 B.n283 B.n282 585
R10 B.n281 B.n280 585
R11 B.n279 B.n278 585
R12 B.n277 B.n276 585
R13 B.n275 B.n274 585
R14 B.n273 B.n272 585
R15 B.n271 B.n270 585
R16 B.n269 B.n268 585
R17 B.n267 B.n266 585
R18 B.n265 B.n264 585
R19 B.n263 B.n262 585
R20 B.n261 B.n260 585
R21 B.n259 B.n258 585
R22 B.n257 B.n256 585
R23 B.n255 B.n254 585
R24 B.n253 B.n252 585
R25 B.n251 B.n250 585
R26 B.n249 B.n248 585
R27 B.n247 B.n246 585
R28 B.n245 B.n244 585
R29 B.n243 B.n242 585
R30 B.n241 B.n240 585
R31 B.n239 B.n238 585
R32 B.n237 B.n236 585
R33 B.n235 B.n234 585
R34 B.n233 B.n232 585
R35 B.n231 B.n230 585
R36 B.n229 B.n228 585
R37 B.n227 B.n226 585
R38 B.n225 B.n224 585
R39 B.n223 B.n222 585
R40 B.n221 B.n220 585
R41 B.n219 B.n218 585
R42 B.n217 B.n216 585
R43 B.n215 B.n214 585
R44 B.n213 B.n212 585
R45 B.n211 B.n210 585
R46 B.n209 B.n208 585
R47 B.n207 B.n206 585
R48 B.n205 B.n204 585
R49 B.n203 B.n202 585
R50 B.n201 B.n200 585
R51 B.n199 B.n198 585
R52 B.n197 B.n196 585
R53 B.n195 B.n194 585
R54 B.n193 B.n192 585
R55 B.n191 B.n190 585
R56 B.n189 B.n188 585
R57 B.n187 B.n186 585
R58 B.n185 B.n184 585
R59 B.n183 B.n182 585
R60 B.n181 B.n180 585
R61 B.n178 B.n177 585
R62 B.n176 B.n175 585
R63 B.n174 B.n173 585
R64 B.n172 B.n171 585
R65 B.n170 B.n169 585
R66 B.n168 B.n167 585
R67 B.n166 B.n165 585
R68 B.n164 B.n163 585
R69 B.n162 B.n161 585
R70 B.n160 B.n159 585
R71 B.n158 B.n157 585
R72 B.n156 B.n155 585
R73 B.n154 B.n153 585
R74 B.n152 B.n151 585
R75 B.n150 B.n149 585
R76 B.n148 B.n147 585
R77 B.n146 B.n145 585
R78 B.n144 B.n143 585
R79 B.n142 B.n141 585
R80 B.n140 B.n139 585
R81 B.n138 B.n137 585
R82 B.n136 B.n135 585
R83 B.n134 B.n133 585
R84 B.n132 B.n131 585
R85 B.n130 B.n129 585
R86 B.n128 B.n127 585
R87 B.n126 B.n125 585
R88 B.n124 B.n123 585
R89 B.n122 B.n121 585
R90 B.n120 B.n119 585
R91 B.n118 B.n117 585
R92 B.n116 B.n115 585
R93 B.n114 B.n113 585
R94 B.n112 B.n111 585
R95 B.n110 B.n109 585
R96 B.n108 B.n107 585
R97 B.n106 B.n105 585
R98 B.n104 B.n103 585
R99 B.n102 B.n101 585
R100 B.n100 B.n99 585
R101 B.n98 B.n97 585
R102 B.n96 B.n95 585
R103 B.n94 B.n93 585
R104 B.n92 B.n91 585
R105 B.n90 B.n89 585
R106 B.n31 B.n30 585
R107 B.n651 B.n650 585
R108 B.n645 B.n83 585
R109 B.n83 B.n28 585
R110 B.n644 B.n27 585
R111 B.n655 B.n27 585
R112 B.n643 B.n26 585
R113 B.n656 B.n26 585
R114 B.n642 B.n25 585
R115 B.n657 B.n25 585
R116 B.n641 B.n640 585
R117 B.n640 B.t6 585
R118 B.n639 B.n21 585
R119 B.n663 B.n21 585
R120 B.n638 B.n20 585
R121 B.n664 B.n20 585
R122 B.n637 B.n19 585
R123 B.n665 B.n19 585
R124 B.n636 B.n635 585
R125 B.n635 B.n15 585
R126 B.n634 B.n14 585
R127 B.n671 B.n14 585
R128 B.n633 B.n13 585
R129 B.n672 B.n13 585
R130 B.n632 B.n12 585
R131 B.n673 B.n12 585
R132 B.n631 B.n630 585
R133 B.n630 B.n629 585
R134 B.n628 B.n627 585
R135 B.n628 B.n8 585
R136 B.n626 B.n7 585
R137 B.n680 B.n7 585
R138 B.n625 B.n6 585
R139 B.n681 B.n6 585
R140 B.n624 B.n5 585
R141 B.n682 B.n5 585
R142 B.n623 B.n622 585
R143 B.n622 B.n4 585
R144 B.n621 B.n289 585
R145 B.n621 B.n620 585
R146 B.n610 B.n290 585
R147 B.n613 B.n290 585
R148 B.n612 B.n611 585
R149 B.n614 B.n612 585
R150 B.n609 B.n295 585
R151 B.n295 B.n294 585
R152 B.n608 B.n607 585
R153 B.n607 B.n606 585
R154 B.n297 B.n296 585
R155 B.n298 B.n297 585
R156 B.n599 B.n598 585
R157 B.n600 B.n599 585
R158 B.n597 B.n303 585
R159 B.n303 B.n302 585
R160 B.n596 B.n595 585
R161 B.n595 B.n594 585
R162 B.n305 B.n304 585
R163 B.t10 B.n305 585
R164 B.n587 B.n586 585
R165 B.n588 B.n587 585
R166 B.n585 B.n310 585
R167 B.n310 B.n309 585
R168 B.n584 B.n583 585
R169 B.n583 B.n582 585
R170 B.n312 B.n311 585
R171 B.n313 B.n312 585
R172 B.n578 B.n577 585
R173 B.n316 B.n315 585
R174 B.n574 B.n573 585
R175 B.n575 B.n574 585
R176 B.n572 B.n367 585
R177 B.n571 B.n570 585
R178 B.n569 B.n568 585
R179 B.n567 B.n566 585
R180 B.n565 B.n564 585
R181 B.n563 B.n562 585
R182 B.n561 B.n560 585
R183 B.n559 B.n558 585
R184 B.n557 B.n556 585
R185 B.n555 B.n554 585
R186 B.n553 B.n552 585
R187 B.n551 B.n550 585
R188 B.n549 B.n548 585
R189 B.n547 B.n546 585
R190 B.n545 B.n544 585
R191 B.n543 B.n542 585
R192 B.n541 B.n540 585
R193 B.n539 B.n538 585
R194 B.n537 B.n536 585
R195 B.n535 B.n534 585
R196 B.n533 B.n532 585
R197 B.n531 B.n530 585
R198 B.n529 B.n528 585
R199 B.n527 B.n526 585
R200 B.n525 B.n524 585
R201 B.n523 B.n522 585
R202 B.n521 B.n520 585
R203 B.n519 B.n518 585
R204 B.n517 B.n516 585
R205 B.n515 B.n514 585
R206 B.n513 B.n512 585
R207 B.n511 B.n510 585
R208 B.n509 B.n508 585
R209 B.n507 B.n506 585
R210 B.n505 B.n504 585
R211 B.n503 B.n502 585
R212 B.n501 B.n500 585
R213 B.n499 B.n498 585
R214 B.n497 B.n496 585
R215 B.n495 B.n494 585
R216 B.n493 B.n492 585
R217 B.n491 B.n490 585
R218 B.n489 B.n488 585
R219 B.n487 B.n486 585
R220 B.n485 B.n484 585
R221 B.n483 B.n482 585
R222 B.n481 B.n480 585
R223 B.n479 B.n478 585
R224 B.n477 B.n476 585
R225 B.n475 B.n474 585
R226 B.n473 B.n472 585
R227 B.n471 B.n470 585
R228 B.n469 B.n468 585
R229 B.n466 B.n465 585
R230 B.n464 B.n463 585
R231 B.n462 B.n461 585
R232 B.n460 B.n459 585
R233 B.n458 B.n457 585
R234 B.n456 B.n455 585
R235 B.n454 B.n453 585
R236 B.n452 B.n451 585
R237 B.n450 B.n449 585
R238 B.n448 B.n447 585
R239 B.n446 B.n445 585
R240 B.n444 B.n443 585
R241 B.n442 B.n441 585
R242 B.n440 B.n439 585
R243 B.n438 B.n437 585
R244 B.n436 B.n435 585
R245 B.n434 B.n433 585
R246 B.n432 B.n431 585
R247 B.n430 B.n429 585
R248 B.n428 B.n427 585
R249 B.n426 B.n425 585
R250 B.n424 B.n423 585
R251 B.n422 B.n421 585
R252 B.n420 B.n419 585
R253 B.n418 B.n417 585
R254 B.n416 B.n415 585
R255 B.n414 B.n413 585
R256 B.n412 B.n411 585
R257 B.n410 B.n409 585
R258 B.n408 B.n407 585
R259 B.n406 B.n405 585
R260 B.n404 B.n403 585
R261 B.n402 B.n401 585
R262 B.n400 B.n399 585
R263 B.n398 B.n397 585
R264 B.n396 B.n395 585
R265 B.n394 B.n393 585
R266 B.n392 B.n391 585
R267 B.n390 B.n389 585
R268 B.n388 B.n387 585
R269 B.n386 B.n385 585
R270 B.n384 B.n383 585
R271 B.n382 B.n381 585
R272 B.n380 B.n379 585
R273 B.n378 B.n377 585
R274 B.n376 B.n375 585
R275 B.n374 B.n373 585
R276 B.n579 B.n314 585
R277 B.n314 B.n313 585
R278 B.n581 B.n580 585
R279 B.n582 B.n581 585
R280 B.n308 B.n307 585
R281 B.n309 B.n308 585
R282 B.n590 B.n589 585
R283 B.n589 B.n588 585
R284 B.n591 B.n306 585
R285 B.n306 B.t10 585
R286 B.n593 B.n592 585
R287 B.n594 B.n593 585
R288 B.n301 B.n300 585
R289 B.n302 B.n301 585
R290 B.n602 B.n601 585
R291 B.n601 B.n600 585
R292 B.n603 B.n299 585
R293 B.n299 B.n298 585
R294 B.n605 B.n604 585
R295 B.n606 B.n605 585
R296 B.n293 B.n292 585
R297 B.n294 B.n293 585
R298 B.n616 B.n615 585
R299 B.n615 B.n614 585
R300 B.n617 B.n291 585
R301 B.n613 B.n291 585
R302 B.n619 B.n618 585
R303 B.n620 B.n619 585
R304 B.n3 B.n0 585
R305 B.n4 B.n3 585
R306 B.n679 B.n1 585
R307 B.n680 B.n679 585
R308 B.n678 B.n677 585
R309 B.n678 B.n8 585
R310 B.n676 B.n9 585
R311 B.n629 B.n9 585
R312 B.n675 B.n674 585
R313 B.n674 B.n673 585
R314 B.n11 B.n10 585
R315 B.n672 B.n11 585
R316 B.n670 B.n669 585
R317 B.n671 B.n670 585
R318 B.n668 B.n16 585
R319 B.n16 B.n15 585
R320 B.n667 B.n666 585
R321 B.n666 B.n665 585
R322 B.n18 B.n17 585
R323 B.n664 B.n18 585
R324 B.n662 B.n661 585
R325 B.n663 B.n662 585
R326 B.n660 B.n22 585
R327 B.n22 B.t6 585
R328 B.n659 B.n658 585
R329 B.n658 B.n657 585
R330 B.n24 B.n23 585
R331 B.n656 B.n24 585
R332 B.n654 B.n653 585
R333 B.n655 B.n654 585
R334 B.n652 B.n29 585
R335 B.n29 B.n28 585
R336 B.n683 B.n682 585
R337 B.n681 B.n2 585
R338 B.n650 B.n29 550.159
R339 B.n647 B.n83 550.159
R340 B.n373 B.n312 550.159
R341 B.n577 B.n314 550.159
R342 B.n648 B.n81 256.663
R343 B.n648 B.n80 256.663
R344 B.n648 B.n79 256.663
R345 B.n648 B.n78 256.663
R346 B.n648 B.n77 256.663
R347 B.n648 B.n76 256.663
R348 B.n648 B.n75 256.663
R349 B.n648 B.n74 256.663
R350 B.n648 B.n73 256.663
R351 B.n648 B.n72 256.663
R352 B.n648 B.n71 256.663
R353 B.n648 B.n70 256.663
R354 B.n648 B.n69 256.663
R355 B.n648 B.n68 256.663
R356 B.n648 B.n67 256.663
R357 B.n648 B.n66 256.663
R358 B.n648 B.n65 256.663
R359 B.n648 B.n64 256.663
R360 B.n648 B.n63 256.663
R361 B.n648 B.n62 256.663
R362 B.n648 B.n61 256.663
R363 B.n648 B.n60 256.663
R364 B.n648 B.n59 256.663
R365 B.n648 B.n58 256.663
R366 B.n648 B.n57 256.663
R367 B.n648 B.n56 256.663
R368 B.n648 B.n55 256.663
R369 B.n648 B.n54 256.663
R370 B.n648 B.n53 256.663
R371 B.n648 B.n52 256.663
R372 B.n648 B.n51 256.663
R373 B.n648 B.n50 256.663
R374 B.n648 B.n49 256.663
R375 B.n648 B.n48 256.663
R376 B.n648 B.n47 256.663
R377 B.n648 B.n46 256.663
R378 B.n648 B.n45 256.663
R379 B.n648 B.n44 256.663
R380 B.n648 B.n43 256.663
R381 B.n648 B.n42 256.663
R382 B.n648 B.n41 256.663
R383 B.n648 B.n40 256.663
R384 B.n648 B.n39 256.663
R385 B.n648 B.n38 256.663
R386 B.n648 B.n37 256.663
R387 B.n648 B.n36 256.663
R388 B.n648 B.n35 256.663
R389 B.n648 B.n34 256.663
R390 B.n648 B.n33 256.663
R391 B.n648 B.n32 256.663
R392 B.n649 B.n648 256.663
R393 B.n576 B.n575 256.663
R394 B.n575 B.n317 256.663
R395 B.n575 B.n318 256.663
R396 B.n575 B.n319 256.663
R397 B.n575 B.n320 256.663
R398 B.n575 B.n321 256.663
R399 B.n575 B.n322 256.663
R400 B.n575 B.n323 256.663
R401 B.n575 B.n324 256.663
R402 B.n575 B.n325 256.663
R403 B.n575 B.n326 256.663
R404 B.n575 B.n327 256.663
R405 B.n575 B.n328 256.663
R406 B.n575 B.n329 256.663
R407 B.n575 B.n330 256.663
R408 B.n575 B.n331 256.663
R409 B.n575 B.n332 256.663
R410 B.n575 B.n333 256.663
R411 B.n575 B.n334 256.663
R412 B.n575 B.n335 256.663
R413 B.n575 B.n336 256.663
R414 B.n575 B.n337 256.663
R415 B.n575 B.n338 256.663
R416 B.n575 B.n339 256.663
R417 B.n575 B.n340 256.663
R418 B.n575 B.n341 256.663
R419 B.n575 B.n342 256.663
R420 B.n575 B.n343 256.663
R421 B.n575 B.n344 256.663
R422 B.n575 B.n345 256.663
R423 B.n575 B.n346 256.663
R424 B.n575 B.n347 256.663
R425 B.n575 B.n348 256.663
R426 B.n575 B.n349 256.663
R427 B.n575 B.n350 256.663
R428 B.n575 B.n351 256.663
R429 B.n575 B.n352 256.663
R430 B.n575 B.n353 256.663
R431 B.n575 B.n354 256.663
R432 B.n575 B.n355 256.663
R433 B.n575 B.n356 256.663
R434 B.n575 B.n357 256.663
R435 B.n575 B.n358 256.663
R436 B.n575 B.n359 256.663
R437 B.n575 B.n360 256.663
R438 B.n575 B.n361 256.663
R439 B.n575 B.n362 256.663
R440 B.n575 B.n363 256.663
R441 B.n575 B.n364 256.663
R442 B.n575 B.n365 256.663
R443 B.n575 B.n366 256.663
R444 B.n685 B.n684 256.663
R445 B.n89 B.n31 163.367
R446 B.n93 B.n92 163.367
R447 B.n97 B.n96 163.367
R448 B.n101 B.n100 163.367
R449 B.n105 B.n104 163.367
R450 B.n109 B.n108 163.367
R451 B.n113 B.n112 163.367
R452 B.n117 B.n116 163.367
R453 B.n121 B.n120 163.367
R454 B.n125 B.n124 163.367
R455 B.n129 B.n128 163.367
R456 B.n133 B.n132 163.367
R457 B.n137 B.n136 163.367
R458 B.n141 B.n140 163.367
R459 B.n145 B.n144 163.367
R460 B.n149 B.n148 163.367
R461 B.n153 B.n152 163.367
R462 B.n157 B.n156 163.367
R463 B.n161 B.n160 163.367
R464 B.n165 B.n164 163.367
R465 B.n169 B.n168 163.367
R466 B.n173 B.n172 163.367
R467 B.n177 B.n176 163.367
R468 B.n182 B.n181 163.367
R469 B.n186 B.n185 163.367
R470 B.n190 B.n189 163.367
R471 B.n194 B.n193 163.367
R472 B.n198 B.n197 163.367
R473 B.n202 B.n201 163.367
R474 B.n206 B.n205 163.367
R475 B.n210 B.n209 163.367
R476 B.n214 B.n213 163.367
R477 B.n218 B.n217 163.367
R478 B.n222 B.n221 163.367
R479 B.n226 B.n225 163.367
R480 B.n230 B.n229 163.367
R481 B.n234 B.n233 163.367
R482 B.n238 B.n237 163.367
R483 B.n242 B.n241 163.367
R484 B.n246 B.n245 163.367
R485 B.n250 B.n249 163.367
R486 B.n254 B.n253 163.367
R487 B.n258 B.n257 163.367
R488 B.n262 B.n261 163.367
R489 B.n266 B.n265 163.367
R490 B.n270 B.n269 163.367
R491 B.n274 B.n273 163.367
R492 B.n278 B.n277 163.367
R493 B.n282 B.n281 163.367
R494 B.n286 B.n285 163.367
R495 B.n647 B.n82 163.367
R496 B.n583 B.n312 163.367
R497 B.n583 B.n310 163.367
R498 B.n587 B.n310 163.367
R499 B.n587 B.n305 163.367
R500 B.n595 B.n305 163.367
R501 B.n595 B.n303 163.367
R502 B.n599 B.n303 163.367
R503 B.n599 B.n297 163.367
R504 B.n607 B.n297 163.367
R505 B.n607 B.n295 163.367
R506 B.n612 B.n295 163.367
R507 B.n612 B.n290 163.367
R508 B.n621 B.n290 163.367
R509 B.n622 B.n621 163.367
R510 B.n622 B.n5 163.367
R511 B.n6 B.n5 163.367
R512 B.n7 B.n6 163.367
R513 B.n628 B.n7 163.367
R514 B.n630 B.n628 163.367
R515 B.n630 B.n12 163.367
R516 B.n13 B.n12 163.367
R517 B.n14 B.n13 163.367
R518 B.n635 B.n14 163.367
R519 B.n635 B.n19 163.367
R520 B.n20 B.n19 163.367
R521 B.n21 B.n20 163.367
R522 B.n640 B.n21 163.367
R523 B.n640 B.n25 163.367
R524 B.n26 B.n25 163.367
R525 B.n27 B.n26 163.367
R526 B.n83 B.n27 163.367
R527 B.n574 B.n316 163.367
R528 B.n574 B.n367 163.367
R529 B.n570 B.n569 163.367
R530 B.n566 B.n565 163.367
R531 B.n562 B.n561 163.367
R532 B.n558 B.n557 163.367
R533 B.n554 B.n553 163.367
R534 B.n550 B.n549 163.367
R535 B.n546 B.n545 163.367
R536 B.n542 B.n541 163.367
R537 B.n538 B.n537 163.367
R538 B.n534 B.n533 163.367
R539 B.n530 B.n529 163.367
R540 B.n526 B.n525 163.367
R541 B.n522 B.n521 163.367
R542 B.n518 B.n517 163.367
R543 B.n514 B.n513 163.367
R544 B.n510 B.n509 163.367
R545 B.n506 B.n505 163.367
R546 B.n502 B.n501 163.367
R547 B.n498 B.n497 163.367
R548 B.n494 B.n493 163.367
R549 B.n490 B.n489 163.367
R550 B.n486 B.n485 163.367
R551 B.n482 B.n481 163.367
R552 B.n478 B.n477 163.367
R553 B.n474 B.n473 163.367
R554 B.n470 B.n469 163.367
R555 B.n465 B.n464 163.367
R556 B.n461 B.n460 163.367
R557 B.n457 B.n456 163.367
R558 B.n453 B.n452 163.367
R559 B.n449 B.n448 163.367
R560 B.n445 B.n444 163.367
R561 B.n441 B.n440 163.367
R562 B.n437 B.n436 163.367
R563 B.n433 B.n432 163.367
R564 B.n429 B.n428 163.367
R565 B.n425 B.n424 163.367
R566 B.n421 B.n420 163.367
R567 B.n417 B.n416 163.367
R568 B.n413 B.n412 163.367
R569 B.n409 B.n408 163.367
R570 B.n405 B.n404 163.367
R571 B.n401 B.n400 163.367
R572 B.n397 B.n396 163.367
R573 B.n393 B.n392 163.367
R574 B.n389 B.n388 163.367
R575 B.n385 B.n384 163.367
R576 B.n381 B.n380 163.367
R577 B.n377 B.n376 163.367
R578 B.n581 B.n314 163.367
R579 B.n581 B.n308 163.367
R580 B.n589 B.n308 163.367
R581 B.n589 B.n306 163.367
R582 B.n593 B.n306 163.367
R583 B.n593 B.n301 163.367
R584 B.n601 B.n301 163.367
R585 B.n601 B.n299 163.367
R586 B.n605 B.n299 163.367
R587 B.n605 B.n293 163.367
R588 B.n615 B.n293 163.367
R589 B.n615 B.n291 163.367
R590 B.n619 B.n291 163.367
R591 B.n619 B.n3 163.367
R592 B.n683 B.n3 163.367
R593 B.n679 B.n2 163.367
R594 B.n679 B.n678 163.367
R595 B.n678 B.n9 163.367
R596 B.n674 B.n9 163.367
R597 B.n674 B.n11 163.367
R598 B.n670 B.n11 163.367
R599 B.n670 B.n16 163.367
R600 B.n666 B.n16 163.367
R601 B.n666 B.n18 163.367
R602 B.n662 B.n18 163.367
R603 B.n662 B.n22 163.367
R604 B.n658 B.n22 163.367
R605 B.n658 B.n24 163.367
R606 B.n654 B.n24 163.367
R607 B.n654 B.n29 163.367
R608 B.n84 B.t17 83.0975
R609 B.n371 B.t15 83.0975
R610 B.n87 B.t7 83.0798
R611 B.n368 B.t12 83.0798
R612 B.n575 B.n313 81.5248
R613 B.n648 B.n28 81.5248
R614 B.n650 B.n649 71.676
R615 B.n89 B.n32 71.676
R616 B.n93 B.n33 71.676
R617 B.n97 B.n34 71.676
R618 B.n101 B.n35 71.676
R619 B.n105 B.n36 71.676
R620 B.n109 B.n37 71.676
R621 B.n113 B.n38 71.676
R622 B.n117 B.n39 71.676
R623 B.n121 B.n40 71.676
R624 B.n125 B.n41 71.676
R625 B.n129 B.n42 71.676
R626 B.n133 B.n43 71.676
R627 B.n137 B.n44 71.676
R628 B.n141 B.n45 71.676
R629 B.n145 B.n46 71.676
R630 B.n149 B.n47 71.676
R631 B.n153 B.n48 71.676
R632 B.n157 B.n49 71.676
R633 B.n161 B.n50 71.676
R634 B.n165 B.n51 71.676
R635 B.n169 B.n52 71.676
R636 B.n173 B.n53 71.676
R637 B.n177 B.n54 71.676
R638 B.n182 B.n55 71.676
R639 B.n186 B.n56 71.676
R640 B.n190 B.n57 71.676
R641 B.n194 B.n58 71.676
R642 B.n198 B.n59 71.676
R643 B.n202 B.n60 71.676
R644 B.n206 B.n61 71.676
R645 B.n210 B.n62 71.676
R646 B.n214 B.n63 71.676
R647 B.n218 B.n64 71.676
R648 B.n222 B.n65 71.676
R649 B.n226 B.n66 71.676
R650 B.n230 B.n67 71.676
R651 B.n234 B.n68 71.676
R652 B.n238 B.n69 71.676
R653 B.n242 B.n70 71.676
R654 B.n246 B.n71 71.676
R655 B.n250 B.n72 71.676
R656 B.n254 B.n73 71.676
R657 B.n258 B.n74 71.676
R658 B.n262 B.n75 71.676
R659 B.n266 B.n76 71.676
R660 B.n270 B.n77 71.676
R661 B.n274 B.n78 71.676
R662 B.n278 B.n79 71.676
R663 B.n282 B.n80 71.676
R664 B.n286 B.n81 71.676
R665 B.n82 B.n81 71.676
R666 B.n285 B.n80 71.676
R667 B.n281 B.n79 71.676
R668 B.n277 B.n78 71.676
R669 B.n273 B.n77 71.676
R670 B.n269 B.n76 71.676
R671 B.n265 B.n75 71.676
R672 B.n261 B.n74 71.676
R673 B.n257 B.n73 71.676
R674 B.n253 B.n72 71.676
R675 B.n249 B.n71 71.676
R676 B.n245 B.n70 71.676
R677 B.n241 B.n69 71.676
R678 B.n237 B.n68 71.676
R679 B.n233 B.n67 71.676
R680 B.n229 B.n66 71.676
R681 B.n225 B.n65 71.676
R682 B.n221 B.n64 71.676
R683 B.n217 B.n63 71.676
R684 B.n213 B.n62 71.676
R685 B.n209 B.n61 71.676
R686 B.n205 B.n60 71.676
R687 B.n201 B.n59 71.676
R688 B.n197 B.n58 71.676
R689 B.n193 B.n57 71.676
R690 B.n189 B.n56 71.676
R691 B.n185 B.n55 71.676
R692 B.n181 B.n54 71.676
R693 B.n176 B.n53 71.676
R694 B.n172 B.n52 71.676
R695 B.n168 B.n51 71.676
R696 B.n164 B.n50 71.676
R697 B.n160 B.n49 71.676
R698 B.n156 B.n48 71.676
R699 B.n152 B.n47 71.676
R700 B.n148 B.n46 71.676
R701 B.n144 B.n45 71.676
R702 B.n140 B.n44 71.676
R703 B.n136 B.n43 71.676
R704 B.n132 B.n42 71.676
R705 B.n128 B.n41 71.676
R706 B.n124 B.n40 71.676
R707 B.n120 B.n39 71.676
R708 B.n116 B.n38 71.676
R709 B.n112 B.n37 71.676
R710 B.n108 B.n36 71.676
R711 B.n104 B.n35 71.676
R712 B.n100 B.n34 71.676
R713 B.n96 B.n33 71.676
R714 B.n92 B.n32 71.676
R715 B.n649 B.n31 71.676
R716 B.n577 B.n576 71.676
R717 B.n367 B.n317 71.676
R718 B.n569 B.n318 71.676
R719 B.n565 B.n319 71.676
R720 B.n561 B.n320 71.676
R721 B.n557 B.n321 71.676
R722 B.n553 B.n322 71.676
R723 B.n549 B.n323 71.676
R724 B.n545 B.n324 71.676
R725 B.n541 B.n325 71.676
R726 B.n537 B.n326 71.676
R727 B.n533 B.n327 71.676
R728 B.n529 B.n328 71.676
R729 B.n525 B.n329 71.676
R730 B.n521 B.n330 71.676
R731 B.n517 B.n331 71.676
R732 B.n513 B.n332 71.676
R733 B.n509 B.n333 71.676
R734 B.n505 B.n334 71.676
R735 B.n501 B.n335 71.676
R736 B.n497 B.n336 71.676
R737 B.n493 B.n337 71.676
R738 B.n489 B.n338 71.676
R739 B.n485 B.n339 71.676
R740 B.n481 B.n340 71.676
R741 B.n477 B.n341 71.676
R742 B.n473 B.n342 71.676
R743 B.n469 B.n343 71.676
R744 B.n464 B.n344 71.676
R745 B.n460 B.n345 71.676
R746 B.n456 B.n346 71.676
R747 B.n452 B.n347 71.676
R748 B.n448 B.n348 71.676
R749 B.n444 B.n349 71.676
R750 B.n440 B.n350 71.676
R751 B.n436 B.n351 71.676
R752 B.n432 B.n352 71.676
R753 B.n428 B.n353 71.676
R754 B.n424 B.n354 71.676
R755 B.n420 B.n355 71.676
R756 B.n416 B.n356 71.676
R757 B.n412 B.n357 71.676
R758 B.n408 B.n358 71.676
R759 B.n404 B.n359 71.676
R760 B.n400 B.n360 71.676
R761 B.n396 B.n361 71.676
R762 B.n392 B.n362 71.676
R763 B.n388 B.n363 71.676
R764 B.n384 B.n364 71.676
R765 B.n380 B.n365 71.676
R766 B.n376 B.n366 71.676
R767 B.n576 B.n316 71.676
R768 B.n570 B.n317 71.676
R769 B.n566 B.n318 71.676
R770 B.n562 B.n319 71.676
R771 B.n558 B.n320 71.676
R772 B.n554 B.n321 71.676
R773 B.n550 B.n322 71.676
R774 B.n546 B.n323 71.676
R775 B.n542 B.n324 71.676
R776 B.n538 B.n325 71.676
R777 B.n534 B.n326 71.676
R778 B.n530 B.n327 71.676
R779 B.n526 B.n328 71.676
R780 B.n522 B.n329 71.676
R781 B.n518 B.n330 71.676
R782 B.n514 B.n331 71.676
R783 B.n510 B.n332 71.676
R784 B.n506 B.n333 71.676
R785 B.n502 B.n334 71.676
R786 B.n498 B.n335 71.676
R787 B.n494 B.n336 71.676
R788 B.n490 B.n337 71.676
R789 B.n486 B.n338 71.676
R790 B.n482 B.n339 71.676
R791 B.n478 B.n340 71.676
R792 B.n474 B.n341 71.676
R793 B.n470 B.n342 71.676
R794 B.n465 B.n343 71.676
R795 B.n461 B.n344 71.676
R796 B.n457 B.n345 71.676
R797 B.n453 B.n346 71.676
R798 B.n449 B.n347 71.676
R799 B.n445 B.n348 71.676
R800 B.n441 B.n349 71.676
R801 B.n437 B.n350 71.676
R802 B.n433 B.n351 71.676
R803 B.n429 B.n352 71.676
R804 B.n425 B.n353 71.676
R805 B.n421 B.n354 71.676
R806 B.n417 B.n355 71.676
R807 B.n413 B.n356 71.676
R808 B.n409 B.n357 71.676
R809 B.n405 B.n358 71.676
R810 B.n401 B.n359 71.676
R811 B.n397 B.n360 71.676
R812 B.n393 B.n361 71.676
R813 B.n389 B.n362 71.676
R814 B.n385 B.n363 71.676
R815 B.n381 B.n364 71.676
R816 B.n377 B.n365 71.676
R817 B.n373 B.n366 71.676
R818 B.n684 B.n683 71.676
R819 B.n684 B.n2 71.676
R820 B.n85 B.t18 70.4915
R821 B.n372 B.t14 70.4915
R822 B.n88 B.t8 70.4738
R823 B.n369 B.t11 70.4738
R824 B.n179 B.n88 59.5399
R825 B.n86 B.n85 59.5399
R826 B.n467 B.n372 59.5399
R827 B.n370 B.n369 59.5399
R828 B.n582 B.n313 39.3172
R829 B.n582 B.n309 39.3172
R830 B.n588 B.n309 39.3172
R831 B.n588 B.t10 39.3172
R832 B.n594 B.t10 39.3172
R833 B.n594 B.n302 39.3172
R834 B.n600 B.n302 39.3172
R835 B.n600 B.n298 39.3172
R836 B.n606 B.n298 39.3172
R837 B.n614 B.n294 39.3172
R838 B.n620 B.n4 39.3172
R839 B.n682 B.n4 39.3172
R840 B.n682 B.n681 39.3172
R841 B.n681 B.n680 39.3172
R842 B.n680 B.n8 39.3172
R843 B.n673 B.n672 39.3172
R844 B.n671 B.n15 39.3172
R845 B.n665 B.n15 39.3172
R846 B.n665 B.n664 39.3172
R847 B.n664 B.n663 39.3172
R848 B.n663 B.t6 39.3172
R849 B.n657 B.t6 39.3172
R850 B.n657 B.n656 39.3172
R851 B.n656 B.n655 39.3172
R852 B.n655 B.n28 39.3172
R853 B.t4 B.n613 38.1608
R854 B.n629 B.t0 38.1608
R855 B.n613 B.t19 37.0044
R856 B.n629 B.t1 37.0044
R857 B.n646 B.n645 35.7468
R858 B.n579 B.n578 35.7468
R859 B.n374 B.n311 35.7468
R860 B.n652 B.n651 35.7468
R861 B.t2 B.n294 34.6917
R862 B.n672 B.t3 34.6917
R863 B B.n685 18.0485
R864 B.n88 B.n87 12.6066
R865 B.n85 B.n84 12.6066
R866 B.n372 B.n371 12.6066
R867 B.n369 B.n368 12.6066
R868 B.n580 B.n579 10.6151
R869 B.n580 B.n307 10.6151
R870 B.n590 B.n307 10.6151
R871 B.n591 B.n590 10.6151
R872 B.n592 B.n591 10.6151
R873 B.n592 B.n300 10.6151
R874 B.n602 B.n300 10.6151
R875 B.n603 B.n602 10.6151
R876 B.n604 B.n603 10.6151
R877 B.n604 B.n292 10.6151
R878 B.n616 B.n292 10.6151
R879 B.n617 B.n616 10.6151
R880 B.n618 B.n617 10.6151
R881 B.n618 B.n0 10.6151
R882 B.n578 B.n315 10.6151
R883 B.n573 B.n315 10.6151
R884 B.n573 B.n572 10.6151
R885 B.n572 B.n571 10.6151
R886 B.n571 B.n568 10.6151
R887 B.n568 B.n567 10.6151
R888 B.n567 B.n564 10.6151
R889 B.n564 B.n563 10.6151
R890 B.n563 B.n560 10.6151
R891 B.n560 B.n559 10.6151
R892 B.n559 B.n556 10.6151
R893 B.n556 B.n555 10.6151
R894 B.n555 B.n552 10.6151
R895 B.n552 B.n551 10.6151
R896 B.n551 B.n548 10.6151
R897 B.n548 B.n547 10.6151
R898 B.n547 B.n544 10.6151
R899 B.n544 B.n543 10.6151
R900 B.n543 B.n540 10.6151
R901 B.n540 B.n539 10.6151
R902 B.n539 B.n536 10.6151
R903 B.n536 B.n535 10.6151
R904 B.n535 B.n532 10.6151
R905 B.n532 B.n531 10.6151
R906 B.n531 B.n528 10.6151
R907 B.n528 B.n527 10.6151
R908 B.n527 B.n524 10.6151
R909 B.n524 B.n523 10.6151
R910 B.n523 B.n520 10.6151
R911 B.n520 B.n519 10.6151
R912 B.n519 B.n516 10.6151
R913 B.n516 B.n515 10.6151
R914 B.n515 B.n512 10.6151
R915 B.n512 B.n511 10.6151
R916 B.n511 B.n508 10.6151
R917 B.n508 B.n507 10.6151
R918 B.n507 B.n504 10.6151
R919 B.n504 B.n503 10.6151
R920 B.n503 B.n500 10.6151
R921 B.n500 B.n499 10.6151
R922 B.n499 B.n496 10.6151
R923 B.n496 B.n495 10.6151
R924 B.n495 B.n492 10.6151
R925 B.n492 B.n491 10.6151
R926 B.n491 B.n488 10.6151
R927 B.n488 B.n487 10.6151
R928 B.n484 B.n483 10.6151
R929 B.n483 B.n480 10.6151
R930 B.n480 B.n479 10.6151
R931 B.n479 B.n476 10.6151
R932 B.n476 B.n475 10.6151
R933 B.n475 B.n472 10.6151
R934 B.n472 B.n471 10.6151
R935 B.n471 B.n468 10.6151
R936 B.n466 B.n463 10.6151
R937 B.n463 B.n462 10.6151
R938 B.n462 B.n459 10.6151
R939 B.n459 B.n458 10.6151
R940 B.n458 B.n455 10.6151
R941 B.n455 B.n454 10.6151
R942 B.n454 B.n451 10.6151
R943 B.n451 B.n450 10.6151
R944 B.n450 B.n447 10.6151
R945 B.n447 B.n446 10.6151
R946 B.n446 B.n443 10.6151
R947 B.n443 B.n442 10.6151
R948 B.n442 B.n439 10.6151
R949 B.n439 B.n438 10.6151
R950 B.n438 B.n435 10.6151
R951 B.n435 B.n434 10.6151
R952 B.n434 B.n431 10.6151
R953 B.n431 B.n430 10.6151
R954 B.n430 B.n427 10.6151
R955 B.n427 B.n426 10.6151
R956 B.n426 B.n423 10.6151
R957 B.n423 B.n422 10.6151
R958 B.n422 B.n419 10.6151
R959 B.n419 B.n418 10.6151
R960 B.n418 B.n415 10.6151
R961 B.n415 B.n414 10.6151
R962 B.n414 B.n411 10.6151
R963 B.n411 B.n410 10.6151
R964 B.n410 B.n407 10.6151
R965 B.n407 B.n406 10.6151
R966 B.n406 B.n403 10.6151
R967 B.n403 B.n402 10.6151
R968 B.n402 B.n399 10.6151
R969 B.n399 B.n398 10.6151
R970 B.n398 B.n395 10.6151
R971 B.n395 B.n394 10.6151
R972 B.n394 B.n391 10.6151
R973 B.n391 B.n390 10.6151
R974 B.n390 B.n387 10.6151
R975 B.n387 B.n386 10.6151
R976 B.n386 B.n383 10.6151
R977 B.n383 B.n382 10.6151
R978 B.n382 B.n379 10.6151
R979 B.n379 B.n378 10.6151
R980 B.n378 B.n375 10.6151
R981 B.n375 B.n374 10.6151
R982 B.n584 B.n311 10.6151
R983 B.n585 B.n584 10.6151
R984 B.n586 B.n585 10.6151
R985 B.n586 B.n304 10.6151
R986 B.n596 B.n304 10.6151
R987 B.n597 B.n596 10.6151
R988 B.n598 B.n597 10.6151
R989 B.n598 B.n296 10.6151
R990 B.n608 B.n296 10.6151
R991 B.n609 B.n608 10.6151
R992 B.n611 B.n609 10.6151
R993 B.n611 B.n610 10.6151
R994 B.n610 B.n289 10.6151
R995 B.n623 B.n289 10.6151
R996 B.n624 B.n623 10.6151
R997 B.n625 B.n624 10.6151
R998 B.n626 B.n625 10.6151
R999 B.n627 B.n626 10.6151
R1000 B.n631 B.n627 10.6151
R1001 B.n632 B.n631 10.6151
R1002 B.n633 B.n632 10.6151
R1003 B.n634 B.n633 10.6151
R1004 B.n636 B.n634 10.6151
R1005 B.n637 B.n636 10.6151
R1006 B.n638 B.n637 10.6151
R1007 B.n639 B.n638 10.6151
R1008 B.n641 B.n639 10.6151
R1009 B.n642 B.n641 10.6151
R1010 B.n643 B.n642 10.6151
R1011 B.n644 B.n643 10.6151
R1012 B.n645 B.n644 10.6151
R1013 B.n677 B.n1 10.6151
R1014 B.n677 B.n676 10.6151
R1015 B.n676 B.n675 10.6151
R1016 B.n675 B.n10 10.6151
R1017 B.n669 B.n10 10.6151
R1018 B.n669 B.n668 10.6151
R1019 B.n668 B.n667 10.6151
R1020 B.n667 B.n17 10.6151
R1021 B.n661 B.n17 10.6151
R1022 B.n661 B.n660 10.6151
R1023 B.n660 B.n659 10.6151
R1024 B.n659 B.n23 10.6151
R1025 B.n653 B.n23 10.6151
R1026 B.n653 B.n652 10.6151
R1027 B.n651 B.n30 10.6151
R1028 B.n90 B.n30 10.6151
R1029 B.n91 B.n90 10.6151
R1030 B.n94 B.n91 10.6151
R1031 B.n95 B.n94 10.6151
R1032 B.n98 B.n95 10.6151
R1033 B.n99 B.n98 10.6151
R1034 B.n102 B.n99 10.6151
R1035 B.n103 B.n102 10.6151
R1036 B.n106 B.n103 10.6151
R1037 B.n107 B.n106 10.6151
R1038 B.n110 B.n107 10.6151
R1039 B.n111 B.n110 10.6151
R1040 B.n114 B.n111 10.6151
R1041 B.n115 B.n114 10.6151
R1042 B.n118 B.n115 10.6151
R1043 B.n119 B.n118 10.6151
R1044 B.n122 B.n119 10.6151
R1045 B.n123 B.n122 10.6151
R1046 B.n126 B.n123 10.6151
R1047 B.n127 B.n126 10.6151
R1048 B.n130 B.n127 10.6151
R1049 B.n131 B.n130 10.6151
R1050 B.n134 B.n131 10.6151
R1051 B.n135 B.n134 10.6151
R1052 B.n138 B.n135 10.6151
R1053 B.n139 B.n138 10.6151
R1054 B.n142 B.n139 10.6151
R1055 B.n143 B.n142 10.6151
R1056 B.n146 B.n143 10.6151
R1057 B.n147 B.n146 10.6151
R1058 B.n150 B.n147 10.6151
R1059 B.n151 B.n150 10.6151
R1060 B.n154 B.n151 10.6151
R1061 B.n155 B.n154 10.6151
R1062 B.n158 B.n155 10.6151
R1063 B.n159 B.n158 10.6151
R1064 B.n162 B.n159 10.6151
R1065 B.n163 B.n162 10.6151
R1066 B.n166 B.n163 10.6151
R1067 B.n167 B.n166 10.6151
R1068 B.n170 B.n167 10.6151
R1069 B.n171 B.n170 10.6151
R1070 B.n174 B.n171 10.6151
R1071 B.n175 B.n174 10.6151
R1072 B.n178 B.n175 10.6151
R1073 B.n183 B.n180 10.6151
R1074 B.n184 B.n183 10.6151
R1075 B.n187 B.n184 10.6151
R1076 B.n188 B.n187 10.6151
R1077 B.n191 B.n188 10.6151
R1078 B.n192 B.n191 10.6151
R1079 B.n195 B.n192 10.6151
R1080 B.n196 B.n195 10.6151
R1081 B.n200 B.n199 10.6151
R1082 B.n203 B.n200 10.6151
R1083 B.n204 B.n203 10.6151
R1084 B.n207 B.n204 10.6151
R1085 B.n208 B.n207 10.6151
R1086 B.n211 B.n208 10.6151
R1087 B.n212 B.n211 10.6151
R1088 B.n215 B.n212 10.6151
R1089 B.n216 B.n215 10.6151
R1090 B.n219 B.n216 10.6151
R1091 B.n220 B.n219 10.6151
R1092 B.n223 B.n220 10.6151
R1093 B.n224 B.n223 10.6151
R1094 B.n227 B.n224 10.6151
R1095 B.n228 B.n227 10.6151
R1096 B.n231 B.n228 10.6151
R1097 B.n232 B.n231 10.6151
R1098 B.n235 B.n232 10.6151
R1099 B.n236 B.n235 10.6151
R1100 B.n239 B.n236 10.6151
R1101 B.n240 B.n239 10.6151
R1102 B.n243 B.n240 10.6151
R1103 B.n244 B.n243 10.6151
R1104 B.n247 B.n244 10.6151
R1105 B.n248 B.n247 10.6151
R1106 B.n251 B.n248 10.6151
R1107 B.n252 B.n251 10.6151
R1108 B.n255 B.n252 10.6151
R1109 B.n256 B.n255 10.6151
R1110 B.n259 B.n256 10.6151
R1111 B.n260 B.n259 10.6151
R1112 B.n263 B.n260 10.6151
R1113 B.n264 B.n263 10.6151
R1114 B.n267 B.n264 10.6151
R1115 B.n268 B.n267 10.6151
R1116 B.n271 B.n268 10.6151
R1117 B.n272 B.n271 10.6151
R1118 B.n275 B.n272 10.6151
R1119 B.n276 B.n275 10.6151
R1120 B.n279 B.n276 10.6151
R1121 B.n280 B.n279 10.6151
R1122 B.n283 B.n280 10.6151
R1123 B.n284 B.n283 10.6151
R1124 B.n287 B.n284 10.6151
R1125 B.n288 B.n287 10.6151
R1126 B.n646 B.n288 10.6151
R1127 B.n685 B.n0 8.11757
R1128 B.n685 B.n1 8.11757
R1129 B.n484 B.n370 6.5566
R1130 B.n468 B.n467 6.5566
R1131 B.n180 B.n179 6.5566
R1132 B.n196 B.n86 6.5566
R1133 B.n606 B.t2 4.62599
R1134 B.t3 B.n671 4.62599
R1135 B.n487 B.n370 4.05904
R1136 B.n467 B.n466 4.05904
R1137 B.n179 B.n178 4.05904
R1138 B.n199 B.n86 4.05904
R1139 B.n620 B.t19 2.31325
R1140 B.t1 B.n8 2.31325
R1141 B.n614 B.t4 1.15687
R1142 B.n673 B.t0 1.15687
R1143 VN.n0 VN.t0 1185.91
R1144 VN.n4 VN.t4 1185.91
R1145 VN.n2 VN.t2 1156.12
R1146 VN.n6 VN.t5 1156.12
R1147 VN.n1 VN.t1 1134.21
R1148 VN.n5 VN.t3 1134.21
R1149 VN.n3 VN.n2 161.3
R1150 VN.n7 VN.n6 161.3
R1151 VN.n2 VN.n1 73.0308
R1152 VN.n6 VN.n5 73.0308
R1153 VN.n7 VN.n4 65.9987
R1154 VN.n3 VN.n0 65.9987
R1155 VN VN.n7 41.4153
R1156 VN.n5 VN.n4 29.7615
R1157 VN.n1 VN.n0 29.7615
R1158 VN VN.n3 0.0516364
R1159 VTAIL.n7 VTAIL.t10 49.5132
R1160 VTAIL.n11 VTAIL.t7 49.513
R1161 VTAIL.n2 VTAIL.t5 49.513
R1162 VTAIL.n10 VTAIL.t3 49.513
R1163 VTAIL.n9 VTAIL.n8 48.0732
R1164 VTAIL.n6 VTAIL.n5 48.0732
R1165 VTAIL.n1 VTAIL.n0 48.073
R1166 VTAIL.n4 VTAIL.n3 48.073
R1167 VTAIL.n6 VTAIL.n4 25.341
R1168 VTAIL.n11 VTAIL.n10 24.7807
R1169 VTAIL.n0 VTAIL.t6 1.4405
R1170 VTAIL.n0 VTAIL.t8 1.4405
R1171 VTAIL.n3 VTAIL.t2 1.4405
R1172 VTAIL.n3 VTAIL.t4 1.4405
R1173 VTAIL.n8 VTAIL.t1 1.4405
R1174 VTAIL.n8 VTAIL.t0 1.4405
R1175 VTAIL.n5 VTAIL.t11 1.4405
R1176 VTAIL.n5 VTAIL.t9 1.4405
R1177 VTAIL.n9 VTAIL.n7 0.7505
R1178 VTAIL.n2 VTAIL.n1 0.7505
R1179 VTAIL.n7 VTAIL.n6 0.560845
R1180 VTAIL.n10 VTAIL.n9 0.560845
R1181 VTAIL.n4 VTAIL.n2 0.560845
R1182 VTAIL VTAIL.n11 0.362569
R1183 VTAIL VTAIL.n1 0.198776
R1184 VDD2.n1 VDD2.t5 66.5567
R1185 VDD2.n2 VDD2.t0 66.192
R1186 VDD2.n1 VDD2.n0 64.8365
R1187 VDD2 VDD2.n3 64.8337
R1188 VDD2.n2 VDD2.n1 37.3899
R1189 VDD2.n3 VDD2.t2 1.4405
R1190 VDD2.n3 VDD2.t1 1.4405
R1191 VDD2.n0 VDD2.t4 1.4405
R1192 VDD2.n0 VDD2.t3 1.4405
R1193 VDD2 VDD2.n2 0.478948
R1194 VP.n1 VP.t5 1185.91
R1195 VP.n8 VP.t0 1156.12
R1196 VP.n6 VP.t4 1156.12
R1197 VP.n3 VP.t2 1156.12
R1198 VP.n7 VP.t1 1134.21
R1199 VP.n2 VP.t3 1134.21
R1200 VP.n9 VP.n8 161.3
R1201 VP.n4 VP.n3 161.3
R1202 VP.n7 VP.n0 161.3
R1203 VP.n6 VP.n5 161.3
R1204 VP.n7 VP.n6 73.0308
R1205 VP.n8 VP.n7 73.0308
R1206 VP.n3 VP.n2 73.0308
R1207 VP.n4 VP.n1 65.9987
R1208 VP.n5 VP.n4 41.0346
R1209 VP.n2 VP.n1 29.7615
R1210 VP.n5 VP.n0 0.189894
R1211 VP.n9 VP.n0 0.189894
R1212 VP VP.n9 0.0516364
R1213 VDD1 VDD1.t0 66.6704
R1214 VDD1.n1 VDD1.t1 66.5567
R1215 VDD1.n1 VDD1.n0 64.8365
R1216 VDD1.n3 VDD1.n2 64.7518
R1217 VDD1.n3 VDD1.n1 38.253
R1218 VDD1.n2 VDD1.t2 1.4405
R1219 VDD1.n2 VDD1.t3 1.4405
R1220 VDD1.n0 VDD1.t4 1.4405
R1221 VDD1.n0 VDD1.t5 1.4405
R1222 VDD1 VDD1.n3 0.0823966
C0 VP VDD2 0.265992f
C1 VN VP 5.03887f
C2 VDD1 VDD2 0.578316f
C3 VDD1 VN 0.147675f
C4 VDD1 VP 3.29277f
C5 VTAIL VDD2 15.350301f
C6 VN VTAIL 2.64907f
C7 VP VTAIL 2.66392f
C8 VDD1 VTAIL 15.321699f
C9 VN VDD2 3.18024f
C10 VDD2 B 4.527487f
C11 VDD1 B 4.732125f
C12 VTAIL B 6.645839f
C13 VN B 7.106019f
C14 VP B 4.736352f
C15 VDD1.t0 B 3.43299f
C16 VDD1.t1 B 3.43237f
C17 VDD1.t4 B 0.298088f
C18 VDD1.t5 B 0.298088f
C19 VDD1.n0 B 2.68762f
C20 VDD1.n1 B 2.28132f
C21 VDD1.t2 B 0.298088f
C22 VDD1.t3 B 0.298088f
C23 VDD1.n2 B 2.68723f
C24 VDD1.n3 B 2.49711f
C25 VP.n0 B 0.057863f
C26 VP.t1 B 0.718866f
C27 VP.t4 B 0.72412f
C28 VP.t5 B 0.731573f
C29 VP.n1 B 0.289518f
C30 VP.t3 B 0.718866f
C31 VP.n2 B 0.297526f
C32 VP.t2 B 0.72412f
C33 VP.n3 B 0.296553f
C34 VP.n4 B 2.4165f
C35 VP.n5 B 2.3476f
C36 VP.n6 B 0.296553f
C37 VP.n7 B 0.297526f
C38 VP.t0 B 0.72412f
C39 VP.n8 B 0.296553f
C40 VP.n9 B 0.044842f
C41 VDD2.t5 B 3.45117f
C42 VDD2.t4 B 0.29972f
C43 VDD2.t3 B 0.29972f
C44 VDD2.n0 B 2.70234f
C45 VDD2.n1 B 2.21796f
C46 VDD2.t0 B 3.44933f
C47 VDD2.n2 B 2.54024f
C48 VDD2.t2 B 0.29972f
C49 VDD2.t1 B 0.29972f
C50 VDD2.n3 B 2.70232f
C51 VTAIL.t6 B 0.304619f
C52 VTAIL.t8 B 0.304619f
C53 VTAIL.n0 B 2.67035f
C54 VTAIL.n1 B 0.347044f
C55 VTAIL.t5 B 3.40816f
C56 VTAIL.n2 B 0.472717f
C57 VTAIL.t2 B 0.304619f
C58 VTAIL.t4 B 0.304619f
C59 VTAIL.n3 B 2.67035f
C60 VTAIL.n4 B 1.86484f
C61 VTAIL.t11 B 0.304619f
C62 VTAIL.t9 B 0.304619f
C63 VTAIL.n5 B 2.67035f
C64 VTAIL.n6 B 1.86484f
C65 VTAIL.t10 B 3.40817f
C66 VTAIL.n7 B 0.472714f
C67 VTAIL.t1 B 0.304619f
C68 VTAIL.t0 B 0.304619f
C69 VTAIL.n8 B 2.67035f
C70 VTAIL.n9 B 0.379748f
C71 VTAIL.t3 B 3.40816f
C72 VTAIL.n10 B 1.90719f
C73 VTAIL.t7 B 3.40816f
C74 VTAIL.n11 B 1.88928f
C75 VN.t0 B 0.712999f
C76 VN.n0 B 0.282167f
C77 VN.t1 B 0.700615f
C78 VN.n1 B 0.289973f
C79 VN.t2 B 0.705736f
C80 VN.n2 B 0.289024f
C81 VN.n3 B 0.160258f
C82 VN.t4 B 0.712999f
C83 VN.n4 B 0.282167f
C84 VN.t5 B 0.705736f
C85 VN.t3 B 0.700615f
C86 VN.n5 B 0.289973f
C87 VN.n6 B 0.289024f
C88 VN.n7 B 2.39222f
.ends

