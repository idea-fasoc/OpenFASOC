* NGSPICE file created from diff_pair_sample_0517.ext - technology: sky130A

.subckt diff_pair_sample_0517 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=2.5707 pd=15.91 as=2.5707 ps=15.91 w=15.58 l=0.87
X1 VTAIL.t14 VN.t1 VDD2.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=6.0762 pd=31.94 as=2.5707 ps=15.91 w=15.58 l=0.87
X2 VDD2.t1 VN.t2 VTAIL.t13 B.t2 sky130_fd_pr__nfet_01v8 ad=2.5707 pd=15.91 as=2.5707 ps=15.91 w=15.58 l=0.87
X3 VDD2.t0 VN.t3 VTAIL.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5707 pd=15.91 as=6.0762 ps=31.94 w=15.58 l=0.87
X4 VTAIL.t5 VP.t0 VDD1.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5707 pd=15.91 as=2.5707 ps=15.91 w=15.58 l=0.87
X5 VTAIL.t11 VN.t4 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=6.0762 pd=31.94 as=2.5707 ps=15.91 w=15.58 l=0.87
X6 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=6.0762 pd=31.94 as=0 ps=0 w=15.58 l=0.87
X7 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=6.0762 pd=31.94 as=0 ps=0 w=15.58 l=0.87
X8 VTAIL.t4 VP.t1 VDD1.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=6.0762 pd=31.94 as=2.5707 ps=15.91 w=15.58 l=0.87
X9 VTAIL.t6 VP.t2 VDD1.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=2.5707 pd=15.91 as=2.5707 ps=15.91 w=15.58 l=0.87
X10 VTAIL.t3 VP.t3 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.0762 pd=31.94 as=2.5707 ps=15.91 w=15.58 l=0.87
X11 VDD1.t3 VP.t4 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.5707 pd=15.91 as=6.0762 ps=31.94 w=15.58 l=0.87
X12 VDD1.t2 VP.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.5707 pd=15.91 as=2.5707 ps=15.91 w=15.58 l=0.87
X13 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=6.0762 pd=31.94 as=0 ps=0 w=15.58 l=0.87
X14 VDD2.t2 VN.t5 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=2.5707 pd=15.91 as=6.0762 ps=31.94 w=15.58 l=0.87
X15 VDD2.t5 VN.t6 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=2.5707 pd=15.91 as=2.5707 ps=15.91 w=15.58 l=0.87
X16 VDD1.t1 VP.t6 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5707 pd=15.91 as=6.0762 ps=31.94 w=15.58 l=0.87
X17 VDD1.t0 VP.t7 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.5707 pd=15.91 as=2.5707 ps=15.91 w=15.58 l=0.87
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.0762 pd=31.94 as=0 ps=0 w=15.58 l=0.87
X19 VTAIL.t8 VN.t7 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5707 pd=15.91 as=2.5707 ps=15.91 w=15.58 l=0.87
R0 VN.n3 VN.t4 498.808
R1 VN.n16 VN.t5 498.808
R2 VN.n11 VN.t3 476.738
R3 VN.n24 VN.t1 476.738
R4 VN.n4 VN.t2 431.584
R5 VN.n1 VN.t7 431.584
R6 VN.n17 VN.t0 431.584
R7 VN.n14 VN.t6 431.584
R8 VN.n12 VN.n11 161.3
R9 VN.n25 VN.n24 161.3
R10 VN.n23 VN.n13 161.3
R11 VN.n22 VN.n21 161.3
R12 VN.n20 VN.n19 161.3
R13 VN.n18 VN.n15 161.3
R14 VN.n10 VN.n0 161.3
R15 VN.n9 VN.n8 161.3
R16 VN.n7 VN.n6 161.3
R17 VN.n5 VN.n2 161.3
R18 VN.n6 VN.n5 56.5617
R19 VN.n19 VN.n18 56.5617
R20 VN VN.n25 45.9266
R21 VN.n10 VN.n9 45.4209
R22 VN.n23 VN.n22 45.4209
R23 VN.n16 VN.n15 42.7264
R24 VN.n3 VN.n2 42.7264
R25 VN.n4 VN.n3 36.9171
R26 VN.n17 VN.n16 36.9171
R27 VN.n5 VN.n4 17.2148
R28 VN.n6 VN.n1 17.2148
R29 VN.n18 VN.n17 17.2148
R30 VN.n19 VN.n14 17.2148
R31 VN.n11 VN.n10 16.7975
R32 VN.n24 VN.n23 16.7975
R33 VN.n9 VN.n1 7.37805
R34 VN.n22 VN.n14 7.37805
R35 VN.n25 VN.n13 0.189894
R36 VN.n21 VN.n13 0.189894
R37 VN.n21 VN.n20 0.189894
R38 VN.n20 VN.n15 0.189894
R39 VN.n7 VN.n2 0.189894
R40 VN.n8 VN.n7 0.189894
R41 VN.n8 VN.n0 0.189894
R42 VN.n12 VN.n0 0.189894
R43 VN VN.n12 0.0516364
R44 VDD2.n2 VDD2.n1 65.571
R45 VDD2.n2 VDD2.n0 65.571
R46 VDD2 VDD2.n5 65.5681
R47 VDD2.n4 VDD2.n3 65.1092
R48 VDD2.n4 VDD2.n2 41.8015
R49 VDD2.n5 VDD2.t7 1.27136
R50 VDD2.n5 VDD2.t2 1.27136
R51 VDD2.n3 VDD2.t6 1.27136
R52 VDD2.n3 VDD2.t5 1.27136
R53 VDD2.n1 VDD2.t4 1.27136
R54 VDD2.n1 VDD2.t0 1.27136
R55 VDD2.n0 VDD2.t3 1.27136
R56 VDD2.n0 VDD2.t1 1.27136
R57 VDD2 VDD2.n4 0.575931
R58 VTAIL.n690 VTAIL.n610 289.615
R59 VTAIL.n82 VTAIL.n2 289.615
R60 VTAIL.n168 VTAIL.n88 289.615
R61 VTAIL.n256 VTAIL.n176 289.615
R62 VTAIL.n604 VTAIL.n524 289.615
R63 VTAIL.n516 VTAIL.n436 289.615
R64 VTAIL.n430 VTAIL.n350 289.615
R65 VTAIL.n342 VTAIL.n262 289.615
R66 VTAIL.n639 VTAIL.n638 185
R67 VTAIL.n641 VTAIL.n640 185
R68 VTAIL.n634 VTAIL.n633 185
R69 VTAIL.n647 VTAIL.n646 185
R70 VTAIL.n649 VTAIL.n648 185
R71 VTAIL.n630 VTAIL.n629 185
R72 VTAIL.n655 VTAIL.n654 185
R73 VTAIL.n657 VTAIL.n656 185
R74 VTAIL.n626 VTAIL.n625 185
R75 VTAIL.n663 VTAIL.n662 185
R76 VTAIL.n665 VTAIL.n664 185
R77 VTAIL.n622 VTAIL.n621 185
R78 VTAIL.n671 VTAIL.n670 185
R79 VTAIL.n673 VTAIL.n672 185
R80 VTAIL.n618 VTAIL.n617 185
R81 VTAIL.n680 VTAIL.n679 185
R82 VTAIL.n681 VTAIL.n616 185
R83 VTAIL.n683 VTAIL.n682 185
R84 VTAIL.n614 VTAIL.n613 185
R85 VTAIL.n689 VTAIL.n688 185
R86 VTAIL.n691 VTAIL.n690 185
R87 VTAIL.n31 VTAIL.n30 185
R88 VTAIL.n33 VTAIL.n32 185
R89 VTAIL.n26 VTAIL.n25 185
R90 VTAIL.n39 VTAIL.n38 185
R91 VTAIL.n41 VTAIL.n40 185
R92 VTAIL.n22 VTAIL.n21 185
R93 VTAIL.n47 VTAIL.n46 185
R94 VTAIL.n49 VTAIL.n48 185
R95 VTAIL.n18 VTAIL.n17 185
R96 VTAIL.n55 VTAIL.n54 185
R97 VTAIL.n57 VTAIL.n56 185
R98 VTAIL.n14 VTAIL.n13 185
R99 VTAIL.n63 VTAIL.n62 185
R100 VTAIL.n65 VTAIL.n64 185
R101 VTAIL.n10 VTAIL.n9 185
R102 VTAIL.n72 VTAIL.n71 185
R103 VTAIL.n73 VTAIL.n8 185
R104 VTAIL.n75 VTAIL.n74 185
R105 VTAIL.n6 VTAIL.n5 185
R106 VTAIL.n81 VTAIL.n80 185
R107 VTAIL.n83 VTAIL.n82 185
R108 VTAIL.n117 VTAIL.n116 185
R109 VTAIL.n119 VTAIL.n118 185
R110 VTAIL.n112 VTAIL.n111 185
R111 VTAIL.n125 VTAIL.n124 185
R112 VTAIL.n127 VTAIL.n126 185
R113 VTAIL.n108 VTAIL.n107 185
R114 VTAIL.n133 VTAIL.n132 185
R115 VTAIL.n135 VTAIL.n134 185
R116 VTAIL.n104 VTAIL.n103 185
R117 VTAIL.n141 VTAIL.n140 185
R118 VTAIL.n143 VTAIL.n142 185
R119 VTAIL.n100 VTAIL.n99 185
R120 VTAIL.n149 VTAIL.n148 185
R121 VTAIL.n151 VTAIL.n150 185
R122 VTAIL.n96 VTAIL.n95 185
R123 VTAIL.n158 VTAIL.n157 185
R124 VTAIL.n159 VTAIL.n94 185
R125 VTAIL.n161 VTAIL.n160 185
R126 VTAIL.n92 VTAIL.n91 185
R127 VTAIL.n167 VTAIL.n166 185
R128 VTAIL.n169 VTAIL.n168 185
R129 VTAIL.n205 VTAIL.n204 185
R130 VTAIL.n207 VTAIL.n206 185
R131 VTAIL.n200 VTAIL.n199 185
R132 VTAIL.n213 VTAIL.n212 185
R133 VTAIL.n215 VTAIL.n214 185
R134 VTAIL.n196 VTAIL.n195 185
R135 VTAIL.n221 VTAIL.n220 185
R136 VTAIL.n223 VTAIL.n222 185
R137 VTAIL.n192 VTAIL.n191 185
R138 VTAIL.n229 VTAIL.n228 185
R139 VTAIL.n231 VTAIL.n230 185
R140 VTAIL.n188 VTAIL.n187 185
R141 VTAIL.n237 VTAIL.n236 185
R142 VTAIL.n239 VTAIL.n238 185
R143 VTAIL.n184 VTAIL.n183 185
R144 VTAIL.n246 VTAIL.n245 185
R145 VTAIL.n247 VTAIL.n182 185
R146 VTAIL.n249 VTAIL.n248 185
R147 VTAIL.n180 VTAIL.n179 185
R148 VTAIL.n255 VTAIL.n254 185
R149 VTAIL.n257 VTAIL.n256 185
R150 VTAIL.n605 VTAIL.n604 185
R151 VTAIL.n603 VTAIL.n602 185
R152 VTAIL.n528 VTAIL.n527 185
R153 VTAIL.n532 VTAIL.n530 185
R154 VTAIL.n597 VTAIL.n596 185
R155 VTAIL.n595 VTAIL.n594 185
R156 VTAIL.n534 VTAIL.n533 185
R157 VTAIL.n589 VTAIL.n588 185
R158 VTAIL.n587 VTAIL.n586 185
R159 VTAIL.n538 VTAIL.n537 185
R160 VTAIL.n581 VTAIL.n580 185
R161 VTAIL.n579 VTAIL.n578 185
R162 VTAIL.n542 VTAIL.n541 185
R163 VTAIL.n573 VTAIL.n572 185
R164 VTAIL.n571 VTAIL.n570 185
R165 VTAIL.n546 VTAIL.n545 185
R166 VTAIL.n565 VTAIL.n564 185
R167 VTAIL.n563 VTAIL.n562 185
R168 VTAIL.n550 VTAIL.n549 185
R169 VTAIL.n557 VTAIL.n556 185
R170 VTAIL.n555 VTAIL.n554 185
R171 VTAIL.n517 VTAIL.n516 185
R172 VTAIL.n515 VTAIL.n514 185
R173 VTAIL.n440 VTAIL.n439 185
R174 VTAIL.n444 VTAIL.n442 185
R175 VTAIL.n509 VTAIL.n508 185
R176 VTAIL.n507 VTAIL.n506 185
R177 VTAIL.n446 VTAIL.n445 185
R178 VTAIL.n501 VTAIL.n500 185
R179 VTAIL.n499 VTAIL.n498 185
R180 VTAIL.n450 VTAIL.n449 185
R181 VTAIL.n493 VTAIL.n492 185
R182 VTAIL.n491 VTAIL.n490 185
R183 VTAIL.n454 VTAIL.n453 185
R184 VTAIL.n485 VTAIL.n484 185
R185 VTAIL.n483 VTAIL.n482 185
R186 VTAIL.n458 VTAIL.n457 185
R187 VTAIL.n477 VTAIL.n476 185
R188 VTAIL.n475 VTAIL.n474 185
R189 VTAIL.n462 VTAIL.n461 185
R190 VTAIL.n469 VTAIL.n468 185
R191 VTAIL.n467 VTAIL.n466 185
R192 VTAIL.n431 VTAIL.n430 185
R193 VTAIL.n429 VTAIL.n428 185
R194 VTAIL.n354 VTAIL.n353 185
R195 VTAIL.n358 VTAIL.n356 185
R196 VTAIL.n423 VTAIL.n422 185
R197 VTAIL.n421 VTAIL.n420 185
R198 VTAIL.n360 VTAIL.n359 185
R199 VTAIL.n415 VTAIL.n414 185
R200 VTAIL.n413 VTAIL.n412 185
R201 VTAIL.n364 VTAIL.n363 185
R202 VTAIL.n407 VTAIL.n406 185
R203 VTAIL.n405 VTAIL.n404 185
R204 VTAIL.n368 VTAIL.n367 185
R205 VTAIL.n399 VTAIL.n398 185
R206 VTAIL.n397 VTAIL.n396 185
R207 VTAIL.n372 VTAIL.n371 185
R208 VTAIL.n391 VTAIL.n390 185
R209 VTAIL.n389 VTAIL.n388 185
R210 VTAIL.n376 VTAIL.n375 185
R211 VTAIL.n383 VTAIL.n382 185
R212 VTAIL.n381 VTAIL.n380 185
R213 VTAIL.n343 VTAIL.n342 185
R214 VTAIL.n341 VTAIL.n340 185
R215 VTAIL.n266 VTAIL.n265 185
R216 VTAIL.n270 VTAIL.n268 185
R217 VTAIL.n335 VTAIL.n334 185
R218 VTAIL.n333 VTAIL.n332 185
R219 VTAIL.n272 VTAIL.n271 185
R220 VTAIL.n327 VTAIL.n326 185
R221 VTAIL.n325 VTAIL.n324 185
R222 VTAIL.n276 VTAIL.n275 185
R223 VTAIL.n319 VTAIL.n318 185
R224 VTAIL.n317 VTAIL.n316 185
R225 VTAIL.n280 VTAIL.n279 185
R226 VTAIL.n311 VTAIL.n310 185
R227 VTAIL.n309 VTAIL.n308 185
R228 VTAIL.n284 VTAIL.n283 185
R229 VTAIL.n303 VTAIL.n302 185
R230 VTAIL.n301 VTAIL.n300 185
R231 VTAIL.n288 VTAIL.n287 185
R232 VTAIL.n295 VTAIL.n294 185
R233 VTAIL.n293 VTAIL.n292 185
R234 VTAIL.n637 VTAIL.t12 147.659
R235 VTAIL.n29 VTAIL.t11 147.659
R236 VTAIL.n115 VTAIL.t7 147.659
R237 VTAIL.n203 VTAIL.t3 147.659
R238 VTAIL.n553 VTAIL.t1 147.659
R239 VTAIL.n465 VTAIL.t4 147.659
R240 VTAIL.n379 VTAIL.t10 147.659
R241 VTAIL.n291 VTAIL.t14 147.659
R242 VTAIL.n640 VTAIL.n639 104.615
R243 VTAIL.n640 VTAIL.n633 104.615
R244 VTAIL.n647 VTAIL.n633 104.615
R245 VTAIL.n648 VTAIL.n647 104.615
R246 VTAIL.n648 VTAIL.n629 104.615
R247 VTAIL.n655 VTAIL.n629 104.615
R248 VTAIL.n656 VTAIL.n655 104.615
R249 VTAIL.n656 VTAIL.n625 104.615
R250 VTAIL.n663 VTAIL.n625 104.615
R251 VTAIL.n664 VTAIL.n663 104.615
R252 VTAIL.n664 VTAIL.n621 104.615
R253 VTAIL.n671 VTAIL.n621 104.615
R254 VTAIL.n672 VTAIL.n671 104.615
R255 VTAIL.n672 VTAIL.n617 104.615
R256 VTAIL.n680 VTAIL.n617 104.615
R257 VTAIL.n681 VTAIL.n680 104.615
R258 VTAIL.n682 VTAIL.n681 104.615
R259 VTAIL.n682 VTAIL.n613 104.615
R260 VTAIL.n689 VTAIL.n613 104.615
R261 VTAIL.n690 VTAIL.n689 104.615
R262 VTAIL.n32 VTAIL.n31 104.615
R263 VTAIL.n32 VTAIL.n25 104.615
R264 VTAIL.n39 VTAIL.n25 104.615
R265 VTAIL.n40 VTAIL.n39 104.615
R266 VTAIL.n40 VTAIL.n21 104.615
R267 VTAIL.n47 VTAIL.n21 104.615
R268 VTAIL.n48 VTAIL.n47 104.615
R269 VTAIL.n48 VTAIL.n17 104.615
R270 VTAIL.n55 VTAIL.n17 104.615
R271 VTAIL.n56 VTAIL.n55 104.615
R272 VTAIL.n56 VTAIL.n13 104.615
R273 VTAIL.n63 VTAIL.n13 104.615
R274 VTAIL.n64 VTAIL.n63 104.615
R275 VTAIL.n64 VTAIL.n9 104.615
R276 VTAIL.n72 VTAIL.n9 104.615
R277 VTAIL.n73 VTAIL.n72 104.615
R278 VTAIL.n74 VTAIL.n73 104.615
R279 VTAIL.n74 VTAIL.n5 104.615
R280 VTAIL.n81 VTAIL.n5 104.615
R281 VTAIL.n82 VTAIL.n81 104.615
R282 VTAIL.n118 VTAIL.n117 104.615
R283 VTAIL.n118 VTAIL.n111 104.615
R284 VTAIL.n125 VTAIL.n111 104.615
R285 VTAIL.n126 VTAIL.n125 104.615
R286 VTAIL.n126 VTAIL.n107 104.615
R287 VTAIL.n133 VTAIL.n107 104.615
R288 VTAIL.n134 VTAIL.n133 104.615
R289 VTAIL.n134 VTAIL.n103 104.615
R290 VTAIL.n141 VTAIL.n103 104.615
R291 VTAIL.n142 VTAIL.n141 104.615
R292 VTAIL.n142 VTAIL.n99 104.615
R293 VTAIL.n149 VTAIL.n99 104.615
R294 VTAIL.n150 VTAIL.n149 104.615
R295 VTAIL.n150 VTAIL.n95 104.615
R296 VTAIL.n158 VTAIL.n95 104.615
R297 VTAIL.n159 VTAIL.n158 104.615
R298 VTAIL.n160 VTAIL.n159 104.615
R299 VTAIL.n160 VTAIL.n91 104.615
R300 VTAIL.n167 VTAIL.n91 104.615
R301 VTAIL.n168 VTAIL.n167 104.615
R302 VTAIL.n206 VTAIL.n205 104.615
R303 VTAIL.n206 VTAIL.n199 104.615
R304 VTAIL.n213 VTAIL.n199 104.615
R305 VTAIL.n214 VTAIL.n213 104.615
R306 VTAIL.n214 VTAIL.n195 104.615
R307 VTAIL.n221 VTAIL.n195 104.615
R308 VTAIL.n222 VTAIL.n221 104.615
R309 VTAIL.n222 VTAIL.n191 104.615
R310 VTAIL.n229 VTAIL.n191 104.615
R311 VTAIL.n230 VTAIL.n229 104.615
R312 VTAIL.n230 VTAIL.n187 104.615
R313 VTAIL.n237 VTAIL.n187 104.615
R314 VTAIL.n238 VTAIL.n237 104.615
R315 VTAIL.n238 VTAIL.n183 104.615
R316 VTAIL.n246 VTAIL.n183 104.615
R317 VTAIL.n247 VTAIL.n246 104.615
R318 VTAIL.n248 VTAIL.n247 104.615
R319 VTAIL.n248 VTAIL.n179 104.615
R320 VTAIL.n255 VTAIL.n179 104.615
R321 VTAIL.n256 VTAIL.n255 104.615
R322 VTAIL.n604 VTAIL.n603 104.615
R323 VTAIL.n603 VTAIL.n527 104.615
R324 VTAIL.n532 VTAIL.n527 104.615
R325 VTAIL.n596 VTAIL.n532 104.615
R326 VTAIL.n596 VTAIL.n595 104.615
R327 VTAIL.n595 VTAIL.n533 104.615
R328 VTAIL.n588 VTAIL.n533 104.615
R329 VTAIL.n588 VTAIL.n587 104.615
R330 VTAIL.n587 VTAIL.n537 104.615
R331 VTAIL.n580 VTAIL.n537 104.615
R332 VTAIL.n580 VTAIL.n579 104.615
R333 VTAIL.n579 VTAIL.n541 104.615
R334 VTAIL.n572 VTAIL.n541 104.615
R335 VTAIL.n572 VTAIL.n571 104.615
R336 VTAIL.n571 VTAIL.n545 104.615
R337 VTAIL.n564 VTAIL.n545 104.615
R338 VTAIL.n564 VTAIL.n563 104.615
R339 VTAIL.n563 VTAIL.n549 104.615
R340 VTAIL.n556 VTAIL.n549 104.615
R341 VTAIL.n556 VTAIL.n555 104.615
R342 VTAIL.n516 VTAIL.n515 104.615
R343 VTAIL.n515 VTAIL.n439 104.615
R344 VTAIL.n444 VTAIL.n439 104.615
R345 VTAIL.n508 VTAIL.n444 104.615
R346 VTAIL.n508 VTAIL.n507 104.615
R347 VTAIL.n507 VTAIL.n445 104.615
R348 VTAIL.n500 VTAIL.n445 104.615
R349 VTAIL.n500 VTAIL.n499 104.615
R350 VTAIL.n499 VTAIL.n449 104.615
R351 VTAIL.n492 VTAIL.n449 104.615
R352 VTAIL.n492 VTAIL.n491 104.615
R353 VTAIL.n491 VTAIL.n453 104.615
R354 VTAIL.n484 VTAIL.n453 104.615
R355 VTAIL.n484 VTAIL.n483 104.615
R356 VTAIL.n483 VTAIL.n457 104.615
R357 VTAIL.n476 VTAIL.n457 104.615
R358 VTAIL.n476 VTAIL.n475 104.615
R359 VTAIL.n475 VTAIL.n461 104.615
R360 VTAIL.n468 VTAIL.n461 104.615
R361 VTAIL.n468 VTAIL.n467 104.615
R362 VTAIL.n430 VTAIL.n429 104.615
R363 VTAIL.n429 VTAIL.n353 104.615
R364 VTAIL.n358 VTAIL.n353 104.615
R365 VTAIL.n422 VTAIL.n358 104.615
R366 VTAIL.n422 VTAIL.n421 104.615
R367 VTAIL.n421 VTAIL.n359 104.615
R368 VTAIL.n414 VTAIL.n359 104.615
R369 VTAIL.n414 VTAIL.n413 104.615
R370 VTAIL.n413 VTAIL.n363 104.615
R371 VTAIL.n406 VTAIL.n363 104.615
R372 VTAIL.n406 VTAIL.n405 104.615
R373 VTAIL.n405 VTAIL.n367 104.615
R374 VTAIL.n398 VTAIL.n367 104.615
R375 VTAIL.n398 VTAIL.n397 104.615
R376 VTAIL.n397 VTAIL.n371 104.615
R377 VTAIL.n390 VTAIL.n371 104.615
R378 VTAIL.n390 VTAIL.n389 104.615
R379 VTAIL.n389 VTAIL.n375 104.615
R380 VTAIL.n382 VTAIL.n375 104.615
R381 VTAIL.n382 VTAIL.n381 104.615
R382 VTAIL.n342 VTAIL.n341 104.615
R383 VTAIL.n341 VTAIL.n265 104.615
R384 VTAIL.n270 VTAIL.n265 104.615
R385 VTAIL.n334 VTAIL.n270 104.615
R386 VTAIL.n334 VTAIL.n333 104.615
R387 VTAIL.n333 VTAIL.n271 104.615
R388 VTAIL.n326 VTAIL.n271 104.615
R389 VTAIL.n326 VTAIL.n325 104.615
R390 VTAIL.n325 VTAIL.n275 104.615
R391 VTAIL.n318 VTAIL.n275 104.615
R392 VTAIL.n318 VTAIL.n317 104.615
R393 VTAIL.n317 VTAIL.n279 104.615
R394 VTAIL.n310 VTAIL.n279 104.615
R395 VTAIL.n310 VTAIL.n309 104.615
R396 VTAIL.n309 VTAIL.n283 104.615
R397 VTAIL.n302 VTAIL.n283 104.615
R398 VTAIL.n302 VTAIL.n301 104.615
R399 VTAIL.n301 VTAIL.n287 104.615
R400 VTAIL.n294 VTAIL.n287 104.615
R401 VTAIL.n294 VTAIL.n293 104.615
R402 VTAIL.n639 VTAIL.t12 52.3082
R403 VTAIL.n31 VTAIL.t11 52.3082
R404 VTAIL.n117 VTAIL.t7 52.3082
R405 VTAIL.n205 VTAIL.t3 52.3082
R406 VTAIL.n555 VTAIL.t1 52.3082
R407 VTAIL.n467 VTAIL.t4 52.3082
R408 VTAIL.n381 VTAIL.t10 52.3082
R409 VTAIL.n293 VTAIL.t14 52.3082
R410 VTAIL.n523 VTAIL.n522 48.4305
R411 VTAIL.n349 VTAIL.n348 48.4305
R412 VTAIL.n1 VTAIL.n0 48.4303
R413 VTAIL.n175 VTAIL.n174 48.4303
R414 VTAIL.n695 VTAIL.n694 36.452
R415 VTAIL.n87 VTAIL.n86 36.452
R416 VTAIL.n173 VTAIL.n172 36.452
R417 VTAIL.n261 VTAIL.n260 36.452
R418 VTAIL.n609 VTAIL.n608 36.452
R419 VTAIL.n521 VTAIL.n520 36.452
R420 VTAIL.n435 VTAIL.n434 36.452
R421 VTAIL.n347 VTAIL.n346 36.452
R422 VTAIL.n695 VTAIL.n609 26.8324
R423 VTAIL.n347 VTAIL.n261 26.8324
R424 VTAIL.n638 VTAIL.n637 15.6677
R425 VTAIL.n30 VTAIL.n29 15.6677
R426 VTAIL.n116 VTAIL.n115 15.6677
R427 VTAIL.n204 VTAIL.n203 15.6677
R428 VTAIL.n554 VTAIL.n553 15.6677
R429 VTAIL.n466 VTAIL.n465 15.6677
R430 VTAIL.n380 VTAIL.n379 15.6677
R431 VTAIL.n292 VTAIL.n291 15.6677
R432 VTAIL.n683 VTAIL.n614 13.1884
R433 VTAIL.n75 VTAIL.n6 13.1884
R434 VTAIL.n161 VTAIL.n92 13.1884
R435 VTAIL.n249 VTAIL.n180 13.1884
R436 VTAIL.n530 VTAIL.n528 13.1884
R437 VTAIL.n442 VTAIL.n440 13.1884
R438 VTAIL.n356 VTAIL.n354 13.1884
R439 VTAIL.n268 VTAIL.n266 13.1884
R440 VTAIL.n641 VTAIL.n636 12.8005
R441 VTAIL.n684 VTAIL.n616 12.8005
R442 VTAIL.n688 VTAIL.n687 12.8005
R443 VTAIL.n33 VTAIL.n28 12.8005
R444 VTAIL.n76 VTAIL.n8 12.8005
R445 VTAIL.n80 VTAIL.n79 12.8005
R446 VTAIL.n119 VTAIL.n114 12.8005
R447 VTAIL.n162 VTAIL.n94 12.8005
R448 VTAIL.n166 VTAIL.n165 12.8005
R449 VTAIL.n207 VTAIL.n202 12.8005
R450 VTAIL.n250 VTAIL.n182 12.8005
R451 VTAIL.n254 VTAIL.n253 12.8005
R452 VTAIL.n602 VTAIL.n601 12.8005
R453 VTAIL.n598 VTAIL.n597 12.8005
R454 VTAIL.n557 VTAIL.n552 12.8005
R455 VTAIL.n514 VTAIL.n513 12.8005
R456 VTAIL.n510 VTAIL.n509 12.8005
R457 VTAIL.n469 VTAIL.n464 12.8005
R458 VTAIL.n428 VTAIL.n427 12.8005
R459 VTAIL.n424 VTAIL.n423 12.8005
R460 VTAIL.n383 VTAIL.n378 12.8005
R461 VTAIL.n340 VTAIL.n339 12.8005
R462 VTAIL.n336 VTAIL.n335 12.8005
R463 VTAIL.n295 VTAIL.n290 12.8005
R464 VTAIL.n642 VTAIL.n634 12.0247
R465 VTAIL.n679 VTAIL.n678 12.0247
R466 VTAIL.n691 VTAIL.n612 12.0247
R467 VTAIL.n34 VTAIL.n26 12.0247
R468 VTAIL.n71 VTAIL.n70 12.0247
R469 VTAIL.n83 VTAIL.n4 12.0247
R470 VTAIL.n120 VTAIL.n112 12.0247
R471 VTAIL.n157 VTAIL.n156 12.0247
R472 VTAIL.n169 VTAIL.n90 12.0247
R473 VTAIL.n208 VTAIL.n200 12.0247
R474 VTAIL.n245 VTAIL.n244 12.0247
R475 VTAIL.n257 VTAIL.n178 12.0247
R476 VTAIL.n605 VTAIL.n526 12.0247
R477 VTAIL.n594 VTAIL.n531 12.0247
R478 VTAIL.n558 VTAIL.n550 12.0247
R479 VTAIL.n517 VTAIL.n438 12.0247
R480 VTAIL.n506 VTAIL.n443 12.0247
R481 VTAIL.n470 VTAIL.n462 12.0247
R482 VTAIL.n431 VTAIL.n352 12.0247
R483 VTAIL.n420 VTAIL.n357 12.0247
R484 VTAIL.n384 VTAIL.n376 12.0247
R485 VTAIL.n343 VTAIL.n264 12.0247
R486 VTAIL.n332 VTAIL.n269 12.0247
R487 VTAIL.n296 VTAIL.n288 12.0247
R488 VTAIL.n646 VTAIL.n645 11.249
R489 VTAIL.n677 VTAIL.n618 11.249
R490 VTAIL.n692 VTAIL.n610 11.249
R491 VTAIL.n38 VTAIL.n37 11.249
R492 VTAIL.n69 VTAIL.n10 11.249
R493 VTAIL.n84 VTAIL.n2 11.249
R494 VTAIL.n124 VTAIL.n123 11.249
R495 VTAIL.n155 VTAIL.n96 11.249
R496 VTAIL.n170 VTAIL.n88 11.249
R497 VTAIL.n212 VTAIL.n211 11.249
R498 VTAIL.n243 VTAIL.n184 11.249
R499 VTAIL.n258 VTAIL.n176 11.249
R500 VTAIL.n606 VTAIL.n524 11.249
R501 VTAIL.n593 VTAIL.n534 11.249
R502 VTAIL.n562 VTAIL.n561 11.249
R503 VTAIL.n518 VTAIL.n436 11.249
R504 VTAIL.n505 VTAIL.n446 11.249
R505 VTAIL.n474 VTAIL.n473 11.249
R506 VTAIL.n432 VTAIL.n350 11.249
R507 VTAIL.n419 VTAIL.n360 11.249
R508 VTAIL.n388 VTAIL.n387 11.249
R509 VTAIL.n344 VTAIL.n262 11.249
R510 VTAIL.n331 VTAIL.n272 11.249
R511 VTAIL.n300 VTAIL.n299 11.249
R512 VTAIL.n649 VTAIL.n632 10.4732
R513 VTAIL.n674 VTAIL.n673 10.4732
R514 VTAIL.n41 VTAIL.n24 10.4732
R515 VTAIL.n66 VTAIL.n65 10.4732
R516 VTAIL.n127 VTAIL.n110 10.4732
R517 VTAIL.n152 VTAIL.n151 10.4732
R518 VTAIL.n215 VTAIL.n198 10.4732
R519 VTAIL.n240 VTAIL.n239 10.4732
R520 VTAIL.n590 VTAIL.n589 10.4732
R521 VTAIL.n565 VTAIL.n548 10.4732
R522 VTAIL.n502 VTAIL.n501 10.4732
R523 VTAIL.n477 VTAIL.n460 10.4732
R524 VTAIL.n416 VTAIL.n415 10.4732
R525 VTAIL.n391 VTAIL.n374 10.4732
R526 VTAIL.n328 VTAIL.n327 10.4732
R527 VTAIL.n303 VTAIL.n286 10.4732
R528 VTAIL.n650 VTAIL.n630 9.69747
R529 VTAIL.n670 VTAIL.n620 9.69747
R530 VTAIL.n42 VTAIL.n22 9.69747
R531 VTAIL.n62 VTAIL.n12 9.69747
R532 VTAIL.n128 VTAIL.n108 9.69747
R533 VTAIL.n148 VTAIL.n98 9.69747
R534 VTAIL.n216 VTAIL.n196 9.69747
R535 VTAIL.n236 VTAIL.n186 9.69747
R536 VTAIL.n586 VTAIL.n536 9.69747
R537 VTAIL.n566 VTAIL.n546 9.69747
R538 VTAIL.n498 VTAIL.n448 9.69747
R539 VTAIL.n478 VTAIL.n458 9.69747
R540 VTAIL.n412 VTAIL.n362 9.69747
R541 VTAIL.n392 VTAIL.n372 9.69747
R542 VTAIL.n324 VTAIL.n274 9.69747
R543 VTAIL.n304 VTAIL.n284 9.69747
R544 VTAIL.n694 VTAIL.n693 9.45567
R545 VTAIL.n86 VTAIL.n85 9.45567
R546 VTAIL.n172 VTAIL.n171 9.45567
R547 VTAIL.n260 VTAIL.n259 9.45567
R548 VTAIL.n608 VTAIL.n607 9.45567
R549 VTAIL.n520 VTAIL.n519 9.45567
R550 VTAIL.n434 VTAIL.n433 9.45567
R551 VTAIL.n346 VTAIL.n345 9.45567
R552 VTAIL.n693 VTAIL.n692 9.3005
R553 VTAIL.n612 VTAIL.n611 9.3005
R554 VTAIL.n687 VTAIL.n686 9.3005
R555 VTAIL.n659 VTAIL.n658 9.3005
R556 VTAIL.n628 VTAIL.n627 9.3005
R557 VTAIL.n653 VTAIL.n652 9.3005
R558 VTAIL.n651 VTAIL.n650 9.3005
R559 VTAIL.n632 VTAIL.n631 9.3005
R560 VTAIL.n645 VTAIL.n644 9.3005
R561 VTAIL.n643 VTAIL.n642 9.3005
R562 VTAIL.n636 VTAIL.n635 9.3005
R563 VTAIL.n661 VTAIL.n660 9.3005
R564 VTAIL.n624 VTAIL.n623 9.3005
R565 VTAIL.n667 VTAIL.n666 9.3005
R566 VTAIL.n669 VTAIL.n668 9.3005
R567 VTAIL.n620 VTAIL.n619 9.3005
R568 VTAIL.n675 VTAIL.n674 9.3005
R569 VTAIL.n677 VTAIL.n676 9.3005
R570 VTAIL.n678 VTAIL.n615 9.3005
R571 VTAIL.n685 VTAIL.n684 9.3005
R572 VTAIL.n85 VTAIL.n84 9.3005
R573 VTAIL.n4 VTAIL.n3 9.3005
R574 VTAIL.n79 VTAIL.n78 9.3005
R575 VTAIL.n51 VTAIL.n50 9.3005
R576 VTAIL.n20 VTAIL.n19 9.3005
R577 VTAIL.n45 VTAIL.n44 9.3005
R578 VTAIL.n43 VTAIL.n42 9.3005
R579 VTAIL.n24 VTAIL.n23 9.3005
R580 VTAIL.n37 VTAIL.n36 9.3005
R581 VTAIL.n35 VTAIL.n34 9.3005
R582 VTAIL.n28 VTAIL.n27 9.3005
R583 VTAIL.n53 VTAIL.n52 9.3005
R584 VTAIL.n16 VTAIL.n15 9.3005
R585 VTAIL.n59 VTAIL.n58 9.3005
R586 VTAIL.n61 VTAIL.n60 9.3005
R587 VTAIL.n12 VTAIL.n11 9.3005
R588 VTAIL.n67 VTAIL.n66 9.3005
R589 VTAIL.n69 VTAIL.n68 9.3005
R590 VTAIL.n70 VTAIL.n7 9.3005
R591 VTAIL.n77 VTAIL.n76 9.3005
R592 VTAIL.n171 VTAIL.n170 9.3005
R593 VTAIL.n90 VTAIL.n89 9.3005
R594 VTAIL.n165 VTAIL.n164 9.3005
R595 VTAIL.n137 VTAIL.n136 9.3005
R596 VTAIL.n106 VTAIL.n105 9.3005
R597 VTAIL.n131 VTAIL.n130 9.3005
R598 VTAIL.n129 VTAIL.n128 9.3005
R599 VTAIL.n110 VTAIL.n109 9.3005
R600 VTAIL.n123 VTAIL.n122 9.3005
R601 VTAIL.n121 VTAIL.n120 9.3005
R602 VTAIL.n114 VTAIL.n113 9.3005
R603 VTAIL.n139 VTAIL.n138 9.3005
R604 VTAIL.n102 VTAIL.n101 9.3005
R605 VTAIL.n145 VTAIL.n144 9.3005
R606 VTAIL.n147 VTAIL.n146 9.3005
R607 VTAIL.n98 VTAIL.n97 9.3005
R608 VTAIL.n153 VTAIL.n152 9.3005
R609 VTAIL.n155 VTAIL.n154 9.3005
R610 VTAIL.n156 VTAIL.n93 9.3005
R611 VTAIL.n163 VTAIL.n162 9.3005
R612 VTAIL.n259 VTAIL.n258 9.3005
R613 VTAIL.n178 VTAIL.n177 9.3005
R614 VTAIL.n253 VTAIL.n252 9.3005
R615 VTAIL.n225 VTAIL.n224 9.3005
R616 VTAIL.n194 VTAIL.n193 9.3005
R617 VTAIL.n219 VTAIL.n218 9.3005
R618 VTAIL.n217 VTAIL.n216 9.3005
R619 VTAIL.n198 VTAIL.n197 9.3005
R620 VTAIL.n211 VTAIL.n210 9.3005
R621 VTAIL.n209 VTAIL.n208 9.3005
R622 VTAIL.n202 VTAIL.n201 9.3005
R623 VTAIL.n227 VTAIL.n226 9.3005
R624 VTAIL.n190 VTAIL.n189 9.3005
R625 VTAIL.n233 VTAIL.n232 9.3005
R626 VTAIL.n235 VTAIL.n234 9.3005
R627 VTAIL.n186 VTAIL.n185 9.3005
R628 VTAIL.n241 VTAIL.n240 9.3005
R629 VTAIL.n243 VTAIL.n242 9.3005
R630 VTAIL.n244 VTAIL.n181 9.3005
R631 VTAIL.n251 VTAIL.n250 9.3005
R632 VTAIL.n540 VTAIL.n539 9.3005
R633 VTAIL.n583 VTAIL.n582 9.3005
R634 VTAIL.n585 VTAIL.n584 9.3005
R635 VTAIL.n536 VTAIL.n535 9.3005
R636 VTAIL.n591 VTAIL.n590 9.3005
R637 VTAIL.n593 VTAIL.n592 9.3005
R638 VTAIL.n531 VTAIL.n529 9.3005
R639 VTAIL.n599 VTAIL.n598 9.3005
R640 VTAIL.n607 VTAIL.n606 9.3005
R641 VTAIL.n526 VTAIL.n525 9.3005
R642 VTAIL.n601 VTAIL.n600 9.3005
R643 VTAIL.n577 VTAIL.n576 9.3005
R644 VTAIL.n575 VTAIL.n574 9.3005
R645 VTAIL.n544 VTAIL.n543 9.3005
R646 VTAIL.n569 VTAIL.n568 9.3005
R647 VTAIL.n567 VTAIL.n566 9.3005
R648 VTAIL.n548 VTAIL.n547 9.3005
R649 VTAIL.n561 VTAIL.n560 9.3005
R650 VTAIL.n559 VTAIL.n558 9.3005
R651 VTAIL.n552 VTAIL.n551 9.3005
R652 VTAIL.n452 VTAIL.n451 9.3005
R653 VTAIL.n495 VTAIL.n494 9.3005
R654 VTAIL.n497 VTAIL.n496 9.3005
R655 VTAIL.n448 VTAIL.n447 9.3005
R656 VTAIL.n503 VTAIL.n502 9.3005
R657 VTAIL.n505 VTAIL.n504 9.3005
R658 VTAIL.n443 VTAIL.n441 9.3005
R659 VTAIL.n511 VTAIL.n510 9.3005
R660 VTAIL.n519 VTAIL.n518 9.3005
R661 VTAIL.n438 VTAIL.n437 9.3005
R662 VTAIL.n513 VTAIL.n512 9.3005
R663 VTAIL.n489 VTAIL.n488 9.3005
R664 VTAIL.n487 VTAIL.n486 9.3005
R665 VTAIL.n456 VTAIL.n455 9.3005
R666 VTAIL.n481 VTAIL.n480 9.3005
R667 VTAIL.n479 VTAIL.n478 9.3005
R668 VTAIL.n460 VTAIL.n459 9.3005
R669 VTAIL.n473 VTAIL.n472 9.3005
R670 VTAIL.n471 VTAIL.n470 9.3005
R671 VTAIL.n464 VTAIL.n463 9.3005
R672 VTAIL.n366 VTAIL.n365 9.3005
R673 VTAIL.n409 VTAIL.n408 9.3005
R674 VTAIL.n411 VTAIL.n410 9.3005
R675 VTAIL.n362 VTAIL.n361 9.3005
R676 VTAIL.n417 VTAIL.n416 9.3005
R677 VTAIL.n419 VTAIL.n418 9.3005
R678 VTAIL.n357 VTAIL.n355 9.3005
R679 VTAIL.n425 VTAIL.n424 9.3005
R680 VTAIL.n433 VTAIL.n432 9.3005
R681 VTAIL.n352 VTAIL.n351 9.3005
R682 VTAIL.n427 VTAIL.n426 9.3005
R683 VTAIL.n403 VTAIL.n402 9.3005
R684 VTAIL.n401 VTAIL.n400 9.3005
R685 VTAIL.n370 VTAIL.n369 9.3005
R686 VTAIL.n395 VTAIL.n394 9.3005
R687 VTAIL.n393 VTAIL.n392 9.3005
R688 VTAIL.n374 VTAIL.n373 9.3005
R689 VTAIL.n387 VTAIL.n386 9.3005
R690 VTAIL.n385 VTAIL.n384 9.3005
R691 VTAIL.n378 VTAIL.n377 9.3005
R692 VTAIL.n278 VTAIL.n277 9.3005
R693 VTAIL.n321 VTAIL.n320 9.3005
R694 VTAIL.n323 VTAIL.n322 9.3005
R695 VTAIL.n274 VTAIL.n273 9.3005
R696 VTAIL.n329 VTAIL.n328 9.3005
R697 VTAIL.n331 VTAIL.n330 9.3005
R698 VTAIL.n269 VTAIL.n267 9.3005
R699 VTAIL.n337 VTAIL.n336 9.3005
R700 VTAIL.n345 VTAIL.n344 9.3005
R701 VTAIL.n264 VTAIL.n263 9.3005
R702 VTAIL.n339 VTAIL.n338 9.3005
R703 VTAIL.n315 VTAIL.n314 9.3005
R704 VTAIL.n313 VTAIL.n312 9.3005
R705 VTAIL.n282 VTAIL.n281 9.3005
R706 VTAIL.n307 VTAIL.n306 9.3005
R707 VTAIL.n305 VTAIL.n304 9.3005
R708 VTAIL.n286 VTAIL.n285 9.3005
R709 VTAIL.n299 VTAIL.n298 9.3005
R710 VTAIL.n297 VTAIL.n296 9.3005
R711 VTAIL.n290 VTAIL.n289 9.3005
R712 VTAIL.n654 VTAIL.n653 8.92171
R713 VTAIL.n669 VTAIL.n622 8.92171
R714 VTAIL.n46 VTAIL.n45 8.92171
R715 VTAIL.n61 VTAIL.n14 8.92171
R716 VTAIL.n132 VTAIL.n131 8.92171
R717 VTAIL.n147 VTAIL.n100 8.92171
R718 VTAIL.n220 VTAIL.n219 8.92171
R719 VTAIL.n235 VTAIL.n188 8.92171
R720 VTAIL.n585 VTAIL.n538 8.92171
R721 VTAIL.n570 VTAIL.n569 8.92171
R722 VTAIL.n497 VTAIL.n450 8.92171
R723 VTAIL.n482 VTAIL.n481 8.92171
R724 VTAIL.n411 VTAIL.n364 8.92171
R725 VTAIL.n396 VTAIL.n395 8.92171
R726 VTAIL.n323 VTAIL.n276 8.92171
R727 VTAIL.n308 VTAIL.n307 8.92171
R728 VTAIL.n657 VTAIL.n628 8.14595
R729 VTAIL.n666 VTAIL.n665 8.14595
R730 VTAIL.n49 VTAIL.n20 8.14595
R731 VTAIL.n58 VTAIL.n57 8.14595
R732 VTAIL.n135 VTAIL.n106 8.14595
R733 VTAIL.n144 VTAIL.n143 8.14595
R734 VTAIL.n223 VTAIL.n194 8.14595
R735 VTAIL.n232 VTAIL.n231 8.14595
R736 VTAIL.n582 VTAIL.n581 8.14595
R737 VTAIL.n573 VTAIL.n544 8.14595
R738 VTAIL.n494 VTAIL.n493 8.14595
R739 VTAIL.n485 VTAIL.n456 8.14595
R740 VTAIL.n408 VTAIL.n407 8.14595
R741 VTAIL.n399 VTAIL.n370 8.14595
R742 VTAIL.n320 VTAIL.n319 8.14595
R743 VTAIL.n311 VTAIL.n282 8.14595
R744 VTAIL.n658 VTAIL.n626 7.3702
R745 VTAIL.n662 VTAIL.n624 7.3702
R746 VTAIL.n50 VTAIL.n18 7.3702
R747 VTAIL.n54 VTAIL.n16 7.3702
R748 VTAIL.n136 VTAIL.n104 7.3702
R749 VTAIL.n140 VTAIL.n102 7.3702
R750 VTAIL.n224 VTAIL.n192 7.3702
R751 VTAIL.n228 VTAIL.n190 7.3702
R752 VTAIL.n578 VTAIL.n540 7.3702
R753 VTAIL.n574 VTAIL.n542 7.3702
R754 VTAIL.n490 VTAIL.n452 7.3702
R755 VTAIL.n486 VTAIL.n454 7.3702
R756 VTAIL.n404 VTAIL.n366 7.3702
R757 VTAIL.n400 VTAIL.n368 7.3702
R758 VTAIL.n316 VTAIL.n278 7.3702
R759 VTAIL.n312 VTAIL.n280 7.3702
R760 VTAIL.n661 VTAIL.n626 6.59444
R761 VTAIL.n662 VTAIL.n661 6.59444
R762 VTAIL.n53 VTAIL.n18 6.59444
R763 VTAIL.n54 VTAIL.n53 6.59444
R764 VTAIL.n139 VTAIL.n104 6.59444
R765 VTAIL.n140 VTAIL.n139 6.59444
R766 VTAIL.n227 VTAIL.n192 6.59444
R767 VTAIL.n228 VTAIL.n227 6.59444
R768 VTAIL.n578 VTAIL.n577 6.59444
R769 VTAIL.n577 VTAIL.n542 6.59444
R770 VTAIL.n490 VTAIL.n489 6.59444
R771 VTAIL.n489 VTAIL.n454 6.59444
R772 VTAIL.n404 VTAIL.n403 6.59444
R773 VTAIL.n403 VTAIL.n368 6.59444
R774 VTAIL.n316 VTAIL.n315 6.59444
R775 VTAIL.n315 VTAIL.n280 6.59444
R776 VTAIL.n658 VTAIL.n657 5.81868
R777 VTAIL.n665 VTAIL.n624 5.81868
R778 VTAIL.n50 VTAIL.n49 5.81868
R779 VTAIL.n57 VTAIL.n16 5.81868
R780 VTAIL.n136 VTAIL.n135 5.81868
R781 VTAIL.n143 VTAIL.n102 5.81868
R782 VTAIL.n224 VTAIL.n223 5.81868
R783 VTAIL.n231 VTAIL.n190 5.81868
R784 VTAIL.n581 VTAIL.n540 5.81868
R785 VTAIL.n574 VTAIL.n573 5.81868
R786 VTAIL.n493 VTAIL.n452 5.81868
R787 VTAIL.n486 VTAIL.n485 5.81868
R788 VTAIL.n407 VTAIL.n366 5.81868
R789 VTAIL.n400 VTAIL.n399 5.81868
R790 VTAIL.n319 VTAIL.n278 5.81868
R791 VTAIL.n312 VTAIL.n311 5.81868
R792 VTAIL.n654 VTAIL.n628 5.04292
R793 VTAIL.n666 VTAIL.n622 5.04292
R794 VTAIL.n46 VTAIL.n20 5.04292
R795 VTAIL.n58 VTAIL.n14 5.04292
R796 VTAIL.n132 VTAIL.n106 5.04292
R797 VTAIL.n144 VTAIL.n100 5.04292
R798 VTAIL.n220 VTAIL.n194 5.04292
R799 VTAIL.n232 VTAIL.n188 5.04292
R800 VTAIL.n582 VTAIL.n538 5.04292
R801 VTAIL.n570 VTAIL.n544 5.04292
R802 VTAIL.n494 VTAIL.n450 5.04292
R803 VTAIL.n482 VTAIL.n456 5.04292
R804 VTAIL.n408 VTAIL.n364 5.04292
R805 VTAIL.n396 VTAIL.n370 5.04292
R806 VTAIL.n320 VTAIL.n276 5.04292
R807 VTAIL.n308 VTAIL.n282 5.04292
R808 VTAIL.n637 VTAIL.n635 4.38563
R809 VTAIL.n29 VTAIL.n27 4.38563
R810 VTAIL.n115 VTAIL.n113 4.38563
R811 VTAIL.n203 VTAIL.n201 4.38563
R812 VTAIL.n553 VTAIL.n551 4.38563
R813 VTAIL.n465 VTAIL.n463 4.38563
R814 VTAIL.n379 VTAIL.n377 4.38563
R815 VTAIL.n291 VTAIL.n289 4.38563
R816 VTAIL.n653 VTAIL.n630 4.26717
R817 VTAIL.n670 VTAIL.n669 4.26717
R818 VTAIL.n45 VTAIL.n22 4.26717
R819 VTAIL.n62 VTAIL.n61 4.26717
R820 VTAIL.n131 VTAIL.n108 4.26717
R821 VTAIL.n148 VTAIL.n147 4.26717
R822 VTAIL.n219 VTAIL.n196 4.26717
R823 VTAIL.n236 VTAIL.n235 4.26717
R824 VTAIL.n586 VTAIL.n585 4.26717
R825 VTAIL.n569 VTAIL.n546 4.26717
R826 VTAIL.n498 VTAIL.n497 4.26717
R827 VTAIL.n481 VTAIL.n458 4.26717
R828 VTAIL.n412 VTAIL.n411 4.26717
R829 VTAIL.n395 VTAIL.n372 4.26717
R830 VTAIL.n324 VTAIL.n323 4.26717
R831 VTAIL.n307 VTAIL.n284 4.26717
R832 VTAIL.n650 VTAIL.n649 3.49141
R833 VTAIL.n673 VTAIL.n620 3.49141
R834 VTAIL.n42 VTAIL.n41 3.49141
R835 VTAIL.n65 VTAIL.n12 3.49141
R836 VTAIL.n128 VTAIL.n127 3.49141
R837 VTAIL.n151 VTAIL.n98 3.49141
R838 VTAIL.n216 VTAIL.n215 3.49141
R839 VTAIL.n239 VTAIL.n186 3.49141
R840 VTAIL.n589 VTAIL.n536 3.49141
R841 VTAIL.n566 VTAIL.n565 3.49141
R842 VTAIL.n501 VTAIL.n448 3.49141
R843 VTAIL.n478 VTAIL.n477 3.49141
R844 VTAIL.n415 VTAIL.n362 3.49141
R845 VTAIL.n392 VTAIL.n391 3.49141
R846 VTAIL.n327 VTAIL.n274 3.49141
R847 VTAIL.n304 VTAIL.n303 3.49141
R848 VTAIL.n646 VTAIL.n632 2.71565
R849 VTAIL.n674 VTAIL.n618 2.71565
R850 VTAIL.n694 VTAIL.n610 2.71565
R851 VTAIL.n38 VTAIL.n24 2.71565
R852 VTAIL.n66 VTAIL.n10 2.71565
R853 VTAIL.n86 VTAIL.n2 2.71565
R854 VTAIL.n124 VTAIL.n110 2.71565
R855 VTAIL.n152 VTAIL.n96 2.71565
R856 VTAIL.n172 VTAIL.n88 2.71565
R857 VTAIL.n212 VTAIL.n198 2.71565
R858 VTAIL.n240 VTAIL.n184 2.71565
R859 VTAIL.n260 VTAIL.n176 2.71565
R860 VTAIL.n608 VTAIL.n524 2.71565
R861 VTAIL.n590 VTAIL.n534 2.71565
R862 VTAIL.n562 VTAIL.n548 2.71565
R863 VTAIL.n520 VTAIL.n436 2.71565
R864 VTAIL.n502 VTAIL.n446 2.71565
R865 VTAIL.n474 VTAIL.n460 2.71565
R866 VTAIL.n434 VTAIL.n350 2.71565
R867 VTAIL.n416 VTAIL.n360 2.71565
R868 VTAIL.n388 VTAIL.n374 2.71565
R869 VTAIL.n346 VTAIL.n262 2.71565
R870 VTAIL.n328 VTAIL.n272 2.71565
R871 VTAIL.n300 VTAIL.n286 2.71565
R872 VTAIL.n645 VTAIL.n634 1.93989
R873 VTAIL.n679 VTAIL.n677 1.93989
R874 VTAIL.n692 VTAIL.n691 1.93989
R875 VTAIL.n37 VTAIL.n26 1.93989
R876 VTAIL.n71 VTAIL.n69 1.93989
R877 VTAIL.n84 VTAIL.n83 1.93989
R878 VTAIL.n123 VTAIL.n112 1.93989
R879 VTAIL.n157 VTAIL.n155 1.93989
R880 VTAIL.n170 VTAIL.n169 1.93989
R881 VTAIL.n211 VTAIL.n200 1.93989
R882 VTAIL.n245 VTAIL.n243 1.93989
R883 VTAIL.n258 VTAIL.n257 1.93989
R884 VTAIL.n606 VTAIL.n605 1.93989
R885 VTAIL.n594 VTAIL.n593 1.93989
R886 VTAIL.n561 VTAIL.n550 1.93989
R887 VTAIL.n518 VTAIL.n517 1.93989
R888 VTAIL.n506 VTAIL.n505 1.93989
R889 VTAIL.n473 VTAIL.n462 1.93989
R890 VTAIL.n432 VTAIL.n431 1.93989
R891 VTAIL.n420 VTAIL.n419 1.93989
R892 VTAIL.n387 VTAIL.n376 1.93989
R893 VTAIL.n344 VTAIL.n343 1.93989
R894 VTAIL.n332 VTAIL.n331 1.93989
R895 VTAIL.n299 VTAIL.n288 1.93989
R896 VTAIL.n0 VTAIL.t13 1.27136
R897 VTAIL.n0 VTAIL.t8 1.27136
R898 VTAIL.n174 VTAIL.t0 1.27136
R899 VTAIL.n174 VTAIL.t6 1.27136
R900 VTAIL.n522 VTAIL.t2 1.27136
R901 VTAIL.n522 VTAIL.t5 1.27136
R902 VTAIL.n348 VTAIL.t9 1.27136
R903 VTAIL.n348 VTAIL.t15 1.27136
R904 VTAIL.n642 VTAIL.n641 1.16414
R905 VTAIL.n678 VTAIL.n616 1.16414
R906 VTAIL.n688 VTAIL.n612 1.16414
R907 VTAIL.n34 VTAIL.n33 1.16414
R908 VTAIL.n70 VTAIL.n8 1.16414
R909 VTAIL.n80 VTAIL.n4 1.16414
R910 VTAIL.n120 VTAIL.n119 1.16414
R911 VTAIL.n156 VTAIL.n94 1.16414
R912 VTAIL.n166 VTAIL.n90 1.16414
R913 VTAIL.n208 VTAIL.n207 1.16414
R914 VTAIL.n244 VTAIL.n182 1.16414
R915 VTAIL.n254 VTAIL.n178 1.16414
R916 VTAIL.n602 VTAIL.n526 1.16414
R917 VTAIL.n597 VTAIL.n531 1.16414
R918 VTAIL.n558 VTAIL.n557 1.16414
R919 VTAIL.n514 VTAIL.n438 1.16414
R920 VTAIL.n509 VTAIL.n443 1.16414
R921 VTAIL.n470 VTAIL.n469 1.16414
R922 VTAIL.n428 VTAIL.n352 1.16414
R923 VTAIL.n423 VTAIL.n357 1.16414
R924 VTAIL.n384 VTAIL.n383 1.16414
R925 VTAIL.n340 VTAIL.n264 1.16414
R926 VTAIL.n335 VTAIL.n269 1.16414
R927 VTAIL.n296 VTAIL.n295 1.16414
R928 VTAIL.n349 VTAIL.n347 1.03498
R929 VTAIL.n435 VTAIL.n349 1.03498
R930 VTAIL.n523 VTAIL.n521 1.03498
R931 VTAIL.n609 VTAIL.n523 1.03498
R932 VTAIL.n261 VTAIL.n175 1.03498
R933 VTAIL.n175 VTAIL.n173 1.03498
R934 VTAIL.n87 VTAIL.n1 1.03498
R935 VTAIL VTAIL.n695 0.976793
R936 VTAIL.n521 VTAIL.n435 0.470328
R937 VTAIL.n173 VTAIL.n87 0.470328
R938 VTAIL.n638 VTAIL.n636 0.388379
R939 VTAIL.n684 VTAIL.n683 0.388379
R940 VTAIL.n687 VTAIL.n614 0.388379
R941 VTAIL.n30 VTAIL.n28 0.388379
R942 VTAIL.n76 VTAIL.n75 0.388379
R943 VTAIL.n79 VTAIL.n6 0.388379
R944 VTAIL.n116 VTAIL.n114 0.388379
R945 VTAIL.n162 VTAIL.n161 0.388379
R946 VTAIL.n165 VTAIL.n92 0.388379
R947 VTAIL.n204 VTAIL.n202 0.388379
R948 VTAIL.n250 VTAIL.n249 0.388379
R949 VTAIL.n253 VTAIL.n180 0.388379
R950 VTAIL.n601 VTAIL.n528 0.388379
R951 VTAIL.n598 VTAIL.n530 0.388379
R952 VTAIL.n554 VTAIL.n552 0.388379
R953 VTAIL.n513 VTAIL.n440 0.388379
R954 VTAIL.n510 VTAIL.n442 0.388379
R955 VTAIL.n466 VTAIL.n464 0.388379
R956 VTAIL.n427 VTAIL.n354 0.388379
R957 VTAIL.n424 VTAIL.n356 0.388379
R958 VTAIL.n380 VTAIL.n378 0.388379
R959 VTAIL.n339 VTAIL.n266 0.388379
R960 VTAIL.n336 VTAIL.n268 0.388379
R961 VTAIL.n292 VTAIL.n290 0.388379
R962 VTAIL.n643 VTAIL.n635 0.155672
R963 VTAIL.n644 VTAIL.n643 0.155672
R964 VTAIL.n644 VTAIL.n631 0.155672
R965 VTAIL.n651 VTAIL.n631 0.155672
R966 VTAIL.n652 VTAIL.n651 0.155672
R967 VTAIL.n652 VTAIL.n627 0.155672
R968 VTAIL.n659 VTAIL.n627 0.155672
R969 VTAIL.n660 VTAIL.n659 0.155672
R970 VTAIL.n660 VTAIL.n623 0.155672
R971 VTAIL.n667 VTAIL.n623 0.155672
R972 VTAIL.n668 VTAIL.n667 0.155672
R973 VTAIL.n668 VTAIL.n619 0.155672
R974 VTAIL.n675 VTAIL.n619 0.155672
R975 VTAIL.n676 VTAIL.n675 0.155672
R976 VTAIL.n676 VTAIL.n615 0.155672
R977 VTAIL.n685 VTAIL.n615 0.155672
R978 VTAIL.n686 VTAIL.n685 0.155672
R979 VTAIL.n686 VTAIL.n611 0.155672
R980 VTAIL.n693 VTAIL.n611 0.155672
R981 VTAIL.n35 VTAIL.n27 0.155672
R982 VTAIL.n36 VTAIL.n35 0.155672
R983 VTAIL.n36 VTAIL.n23 0.155672
R984 VTAIL.n43 VTAIL.n23 0.155672
R985 VTAIL.n44 VTAIL.n43 0.155672
R986 VTAIL.n44 VTAIL.n19 0.155672
R987 VTAIL.n51 VTAIL.n19 0.155672
R988 VTAIL.n52 VTAIL.n51 0.155672
R989 VTAIL.n52 VTAIL.n15 0.155672
R990 VTAIL.n59 VTAIL.n15 0.155672
R991 VTAIL.n60 VTAIL.n59 0.155672
R992 VTAIL.n60 VTAIL.n11 0.155672
R993 VTAIL.n67 VTAIL.n11 0.155672
R994 VTAIL.n68 VTAIL.n67 0.155672
R995 VTAIL.n68 VTAIL.n7 0.155672
R996 VTAIL.n77 VTAIL.n7 0.155672
R997 VTAIL.n78 VTAIL.n77 0.155672
R998 VTAIL.n78 VTAIL.n3 0.155672
R999 VTAIL.n85 VTAIL.n3 0.155672
R1000 VTAIL.n121 VTAIL.n113 0.155672
R1001 VTAIL.n122 VTAIL.n121 0.155672
R1002 VTAIL.n122 VTAIL.n109 0.155672
R1003 VTAIL.n129 VTAIL.n109 0.155672
R1004 VTAIL.n130 VTAIL.n129 0.155672
R1005 VTAIL.n130 VTAIL.n105 0.155672
R1006 VTAIL.n137 VTAIL.n105 0.155672
R1007 VTAIL.n138 VTAIL.n137 0.155672
R1008 VTAIL.n138 VTAIL.n101 0.155672
R1009 VTAIL.n145 VTAIL.n101 0.155672
R1010 VTAIL.n146 VTAIL.n145 0.155672
R1011 VTAIL.n146 VTAIL.n97 0.155672
R1012 VTAIL.n153 VTAIL.n97 0.155672
R1013 VTAIL.n154 VTAIL.n153 0.155672
R1014 VTAIL.n154 VTAIL.n93 0.155672
R1015 VTAIL.n163 VTAIL.n93 0.155672
R1016 VTAIL.n164 VTAIL.n163 0.155672
R1017 VTAIL.n164 VTAIL.n89 0.155672
R1018 VTAIL.n171 VTAIL.n89 0.155672
R1019 VTAIL.n209 VTAIL.n201 0.155672
R1020 VTAIL.n210 VTAIL.n209 0.155672
R1021 VTAIL.n210 VTAIL.n197 0.155672
R1022 VTAIL.n217 VTAIL.n197 0.155672
R1023 VTAIL.n218 VTAIL.n217 0.155672
R1024 VTAIL.n218 VTAIL.n193 0.155672
R1025 VTAIL.n225 VTAIL.n193 0.155672
R1026 VTAIL.n226 VTAIL.n225 0.155672
R1027 VTAIL.n226 VTAIL.n189 0.155672
R1028 VTAIL.n233 VTAIL.n189 0.155672
R1029 VTAIL.n234 VTAIL.n233 0.155672
R1030 VTAIL.n234 VTAIL.n185 0.155672
R1031 VTAIL.n241 VTAIL.n185 0.155672
R1032 VTAIL.n242 VTAIL.n241 0.155672
R1033 VTAIL.n242 VTAIL.n181 0.155672
R1034 VTAIL.n251 VTAIL.n181 0.155672
R1035 VTAIL.n252 VTAIL.n251 0.155672
R1036 VTAIL.n252 VTAIL.n177 0.155672
R1037 VTAIL.n259 VTAIL.n177 0.155672
R1038 VTAIL.n607 VTAIL.n525 0.155672
R1039 VTAIL.n600 VTAIL.n525 0.155672
R1040 VTAIL.n600 VTAIL.n599 0.155672
R1041 VTAIL.n599 VTAIL.n529 0.155672
R1042 VTAIL.n592 VTAIL.n529 0.155672
R1043 VTAIL.n592 VTAIL.n591 0.155672
R1044 VTAIL.n591 VTAIL.n535 0.155672
R1045 VTAIL.n584 VTAIL.n535 0.155672
R1046 VTAIL.n584 VTAIL.n583 0.155672
R1047 VTAIL.n583 VTAIL.n539 0.155672
R1048 VTAIL.n576 VTAIL.n539 0.155672
R1049 VTAIL.n576 VTAIL.n575 0.155672
R1050 VTAIL.n575 VTAIL.n543 0.155672
R1051 VTAIL.n568 VTAIL.n543 0.155672
R1052 VTAIL.n568 VTAIL.n567 0.155672
R1053 VTAIL.n567 VTAIL.n547 0.155672
R1054 VTAIL.n560 VTAIL.n547 0.155672
R1055 VTAIL.n560 VTAIL.n559 0.155672
R1056 VTAIL.n559 VTAIL.n551 0.155672
R1057 VTAIL.n519 VTAIL.n437 0.155672
R1058 VTAIL.n512 VTAIL.n437 0.155672
R1059 VTAIL.n512 VTAIL.n511 0.155672
R1060 VTAIL.n511 VTAIL.n441 0.155672
R1061 VTAIL.n504 VTAIL.n441 0.155672
R1062 VTAIL.n504 VTAIL.n503 0.155672
R1063 VTAIL.n503 VTAIL.n447 0.155672
R1064 VTAIL.n496 VTAIL.n447 0.155672
R1065 VTAIL.n496 VTAIL.n495 0.155672
R1066 VTAIL.n495 VTAIL.n451 0.155672
R1067 VTAIL.n488 VTAIL.n451 0.155672
R1068 VTAIL.n488 VTAIL.n487 0.155672
R1069 VTAIL.n487 VTAIL.n455 0.155672
R1070 VTAIL.n480 VTAIL.n455 0.155672
R1071 VTAIL.n480 VTAIL.n479 0.155672
R1072 VTAIL.n479 VTAIL.n459 0.155672
R1073 VTAIL.n472 VTAIL.n459 0.155672
R1074 VTAIL.n472 VTAIL.n471 0.155672
R1075 VTAIL.n471 VTAIL.n463 0.155672
R1076 VTAIL.n433 VTAIL.n351 0.155672
R1077 VTAIL.n426 VTAIL.n351 0.155672
R1078 VTAIL.n426 VTAIL.n425 0.155672
R1079 VTAIL.n425 VTAIL.n355 0.155672
R1080 VTAIL.n418 VTAIL.n355 0.155672
R1081 VTAIL.n418 VTAIL.n417 0.155672
R1082 VTAIL.n417 VTAIL.n361 0.155672
R1083 VTAIL.n410 VTAIL.n361 0.155672
R1084 VTAIL.n410 VTAIL.n409 0.155672
R1085 VTAIL.n409 VTAIL.n365 0.155672
R1086 VTAIL.n402 VTAIL.n365 0.155672
R1087 VTAIL.n402 VTAIL.n401 0.155672
R1088 VTAIL.n401 VTAIL.n369 0.155672
R1089 VTAIL.n394 VTAIL.n369 0.155672
R1090 VTAIL.n394 VTAIL.n393 0.155672
R1091 VTAIL.n393 VTAIL.n373 0.155672
R1092 VTAIL.n386 VTAIL.n373 0.155672
R1093 VTAIL.n386 VTAIL.n385 0.155672
R1094 VTAIL.n385 VTAIL.n377 0.155672
R1095 VTAIL.n345 VTAIL.n263 0.155672
R1096 VTAIL.n338 VTAIL.n263 0.155672
R1097 VTAIL.n338 VTAIL.n337 0.155672
R1098 VTAIL.n337 VTAIL.n267 0.155672
R1099 VTAIL.n330 VTAIL.n267 0.155672
R1100 VTAIL.n330 VTAIL.n329 0.155672
R1101 VTAIL.n329 VTAIL.n273 0.155672
R1102 VTAIL.n322 VTAIL.n273 0.155672
R1103 VTAIL.n322 VTAIL.n321 0.155672
R1104 VTAIL.n321 VTAIL.n277 0.155672
R1105 VTAIL.n314 VTAIL.n277 0.155672
R1106 VTAIL.n314 VTAIL.n313 0.155672
R1107 VTAIL.n313 VTAIL.n281 0.155672
R1108 VTAIL.n306 VTAIL.n281 0.155672
R1109 VTAIL.n306 VTAIL.n305 0.155672
R1110 VTAIL.n305 VTAIL.n285 0.155672
R1111 VTAIL.n298 VTAIL.n285 0.155672
R1112 VTAIL.n298 VTAIL.n297 0.155672
R1113 VTAIL.n297 VTAIL.n289 0.155672
R1114 VTAIL VTAIL.n1 0.0586897
R1115 B.n110 B.t12 633.54
R1116 B.n107 B.t8 633.54
R1117 B.n445 B.t15 633.54
R1118 B.n443 B.t19 633.54
R1119 B.n786 B.n785 585
R1120 B.n337 B.n106 585
R1121 B.n336 B.n335 585
R1122 B.n334 B.n333 585
R1123 B.n332 B.n331 585
R1124 B.n330 B.n329 585
R1125 B.n328 B.n327 585
R1126 B.n326 B.n325 585
R1127 B.n324 B.n323 585
R1128 B.n322 B.n321 585
R1129 B.n320 B.n319 585
R1130 B.n318 B.n317 585
R1131 B.n316 B.n315 585
R1132 B.n314 B.n313 585
R1133 B.n312 B.n311 585
R1134 B.n310 B.n309 585
R1135 B.n308 B.n307 585
R1136 B.n306 B.n305 585
R1137 B.n304 B.n303 585
R1138 B.n302 B.n301 585
R1139 B.n300 B.n299 585
R1140 B.n298 B.n297 585
R1141 B.n296 B.n295 585
R1142 B.n294 B.n293 585
R1143 B.n292 B.n291 585
R1144 B.n290 B.n289 585
R1145 B.n288 B.n287 585
R1146 B.n286 B.n285 585
R1147 B.n284 B.n283 585
R1148 B.n282 B.n281 585
R1149 B.n280 B.n279 585
R1150 B.n278 B.n277 585
R1151 B.n276 B.n275 585
R1152 B.n274 B.n273 585
R1153 B.n272 B.n271 585
R1154 B.n270 B.n269 585
R1155 B.n268 B.n267 585
R1156 B.n266 B.n265 585
R1157 B.n264 B.n263 585
R1158 B.n262 B.n261 585
R1159 B.n260 B.n259 585
R1160 B.n258 B.n257 585
R1161 B.n256 B.n255 585
R1162 B.n254 B.n253 585
R1163 B.n252 B.n251 585
R1164 B.n250 B.n249 585
R1165 B.n248 B.n247 585
R1166 B.n246 B.n245 585
R1167 B.n244 B.n243 585
R1168 B.n242 B.n241 585
R1169 B.n240 B.n239 585
R1170 B.n238 B.n237 585
R1171 B.n236 B.n235 585
R1172 B.n234 B.n233 585
R1173 B.n232 B.n231 585
R1174 B.n230 B.n229 585
R1175 B.n228 B.n227 585
R1176 B.n226 B.n225 585
R1177 B.n224 B.n223 585
R1178 B.n222 B.n221 585
R1179 B.n220 B.n219 585
R1180 B.n218 B.n217 585
R1181 B.n216 B.n215 585
R1182 B.n214 B.n213 585
R1183 B.n212 B.n211 585
R1184 B.n210 B.n209 585
R1185 B.n208 B.n207 585
R1186 B.n206 B.n205 585
R1187 B.n204 B.n203 585
R1188 B.n202 B.n201 585
R1189 B.n200 B.n199 585
R1190 B.n198 B.n197 585
R1191 B.n196 B.n195 585
R1192 B.n194 B.n193 585
R1193 B.n192 B.n191 585
R1194 B.n190 B.n189 585
R1195 B.n188 B.n187 585
R1196 B.n186 B.n185 585
R1197 B.n184 B.n183 585
R1198 B.n182 B.n181 585
R1199 B.n180 B.n179 585
R1200 B.n178 B.n177 585
R1201 B.n176 B.n175 585
R1202 B.n174 B.n173 585
R1203 B.n172 B.n171 585
R1204 B.n170 B.n169 585
R1205 B.n168 B.n167 585
R1206 B.n166 B.n165 585
R1207 B.n164 B.n163 585
R1208 B.n162 B.n161 585
R1209 B.n160 B.n159 585
R1210 B.n158 B.n157 585
R1211 B.n156 B.n155 585
R1212 B.n154 B.n153 585
R1213 B.n152 B.n151 585
R1214 B.n150 B.n149 585
R1215 B.n148 B.n147 585
R1216 B.n146 B.n145 585
R1217 B.n144 B.n143 585
R1218 B.n142 B.n141 585
R1219 B.n140 B.n139 585
R1220 B.n138 B.n137 585
R1221 B.n136 B.n135 585
R1222 B.n134 B.n133 585
R1223 B.n132 B.n131 585
R1224 B.n130 B.n129 585
R1225 B.n128 B.n127 585
R1226 B.n126 B.n125 585
R1227 B.n124 B.n123 585
R1228 B.n122 B.n121 585
R1229 B.n120 B.n119 585
R1230 B.n118 B.n117 585
R1231 B.n116 B.n115 585
R1232 B.n114 B.n113 585
R1233 B.n784 B.n49 585
R1234 B.n789 B.n49 585
R1235 B.n783 B.n48 585
R1236 B.n790 B.n48 585
R1237 B.n782 B.n781 585
R1238 B.n781 B.n44 585
R1239 B.n780 B.n43 585
R1240 B.n796 B.n43 585
R1241 B.n779 B.n42 585
R1242 B.n797 B.n42 585
R1243 B.n778 B.n41 585
R1244 B.n798 B.n41 585
R1245 B.n777 B.n776 585
R1246 B.n776 B.n37 585
R1247 B.n775 B.n36 585
R1248 B.n804 B.n36 585
R1249 B.n774 B.n35 585
R1250 B.n805 B.n35 585
R1251 B.n773 B.n34 585
R1252 B.n806 B.n34 585
R1253 B.n772 B.n771 585
R1254 B.n771 B.n30 585
R1255 B.n770 B.n29 585
R1256 B.n812 B.n29 585
R1257 B.n769 B.n28 585
R1258 B.n813 B.n28 585
R1259 B.n768 B.n27 585
R1260 B.n814 B.n27 585
R1261 B.n767 B.n766 585
R1262 B.n766 B.n23 585
R1263 B.n765 B.n22 585
R1264 B.n820 B.n22 585
R1265 B.n764 B.n21 585
R1266 B.n821 B.n21 585
R1267 B.n763 B.n20 585
R1268 B.n822 B.n20 585
R1269 B.n762 B.n761 585
R1270 B.n761 B.n19 585
R1271 B.n760 B.n15 585
R1272 B.n828 B.n15 585
R1273 B.n759 B.n14 585
R1274 B.n829 B.n14 585
R1275 B.n758 B.n13 585
R1276 B.n830 B.n13 585
R1277 B.n757 B.n756 585
R1278 B.n756 B.n12 585
R1279 B.n755 B.n754 585
R1280 B.n755 B.n8 585
R1281 B.n753 B.n7 585
R1282 B.n837 B.n7 585
R1283 B.n752 B.n6 585
R1284 B.n838 B.n6 585
R1285 B.n751 B.n5 585
R1286 B.n839 B.n5 585
R1287 B.n750 B.n749 585
R1288 B.n749 B.n4 585
R1289 B.n748 B.n338 585
R1290 B.n748 B.n747 585
R1291 B.n737 B.n339 585
R1292 B.n740 B.n339 585
R1293 B.n739 B.n738 585
R1294 B.n741 B.n739 585
R1295 B.n736 B.n344 585
R1296 B.n344 B.n343 585
R1297 B.n735 B.n734 585
R1298 B.n734 B.n733 585
R1299 B.n346 B.n345 585
R1300 B.n726 B.n346 585
R1301 B.n725 B.n724 585
R1302 B.n727 B.n725 585
R1303 B.n723 B.n351 585
R1304 B.n351 B.n350 585
R1305 B.n722 B.n721 585
R1306 B.n721 B.n720 585
R1307 B.n353 B.n352 585
R1308 B.n354 B.n353 585
R1309 B.n713 B.n712 585
R1310 B.n714 B.n713 585
R1311 B.n711 B.n359 585
R1312 B.n359 B.n358 585
R1313 B.n710 B.n709 585
R1314 B.n709 B.n708 585
R1315 B.n361 B.n360 585
R1316 B.n362 B.n361 585
R1317 B.n701 B.n700 585
R1318 B.n702 B.n701 585
R1319 B.n699 B.n367 585
R1320 B.n367 B.n366 585
R1321 B.n698 B.n697 585
R1322 B.n697 B.n696 585
R1323 B.n369 B.n368 585
R1324 B.n370 B.n369 585
R1325 B.n689 B.n688 585
R1326 B.n690 B.n689 585
R1327 B.n687 B.n374 585
R1328 B.n378 B.n374 585
R1329 B.n686 B.n685 585
R1330 B.n685 B.n684 585
R1331 B.n376 B.n375 585
R1332 B.n377 B.n376 585
R1333 B.n677 B.n676 585
R1334 B.n678 B.n677 585
R1335 B.n675 B.n383 585
R1336 B.n383 B.n382 585
R1337 B.n670 B.n669 585
R1338 B.n668 B.n442 585
R1339 B.n667 B.n441 585
R1340 B.n672 B.n441 585
R1341 B.n666 B.n665 585
R1342 B.n664 B.n663 585
R1343 B.n662 B.n661 585
R1344 B.n660 B.n659 585
R1345 B.n658 B.n657 585
R1346 B.n656 B.n655 585
R1347 B.n654 B.n653 585
R1348 B.n652 B.n651 585
R1349 B.n650 B.n649 585
R1350 B.n648 B.n647 585
R1351 B.n646 B.n645 585
R1352 B.n644 B.n643 585
R1353 B.n642 B.n641 585
R1354 B.n640 B.n639 585
R1355 B.n638 B.n637 585
R1356 B.n636 B.n635 585
R1357 B.n634 B.n633 585
R1358 B.n632 B.n631 585
R1359 B.n630 B.n629 585
R1360 B.n628 B.n627 585
R1361 B.n626 B.n625 585
R1362 B.n624 B.n623 585
R1363 B.n622 B.n621 585
R1364 B.n620 B.n619 585
R1365 B.n618 B.n617 585
R1366 B.n616 B.n615 585
R1367 B.n614 B.n613 585
R1368 B.n612 B.n611 585
R1369 B.n610 B.n609 585
R1370 B.n608 B.n607 585
R1371 B.n606 B.n605 585
R1372 B.n604 B.n603 585
R1373 B.n602 B.n601 585
R1374 B.n600 B.n599 585
R1375 B.n598 B.n597 585
R1376 B.n596 B.n595 585
R1377 B.n594 B.n593 585
R1378 B.n592 B.n591 585
R1379 B.n590 B.n589 585
R1380 B.n588 B.n587 585
R1381 B.n586 B.n585 585
R1382 B.n584 B.n583 585
R1383 B.n582 B.n581 585
R1384 B.n580 B.n579 585
R1385 B.n578 B.n577 585
R1386 B.n576 B.n575 585
R1387 B.n574 B.n573 585
R1388 B.n572 B.n571 585
R1389 B.n570 B.n569 585
R1390 B.n567 B.n566 585
R1391 B.n565 B.n564 585
R1392 B.n563 B.n562 585
R1393 B.n561 B.n560 585
R1394 B.n559 B.n558 585
R1395 B.n557 B.n556 585
R1396 B.n555 B.n554 585
R1397 B.n553 B.n552 585
R1398 B.n551 B.n550 585
R1399 B.n549 B.n548 585
R1400 B.n546 B.n545 585
R1401 B.n544 B.n543 585
R1402 B.n542 B.n541 585
R1403 B.n540 B.n539 585
R1404 B.n538 B.n537 585
R1405 B.n536 B.n535 585
R1406 B.n534 B.n533 585
R1407 B.n532 B.n531 585
R1408 B.n530 B.n529 585
R1409 B.n528 B.n527 585
R1410 B.n526 B.n525 585
R1411 B.n524 B.n523 585
R1412 B.n522 B.n521 585
R1413 B.n520 B.n519 585
R1414 B.n518 B.n517 585
R1415 B.n516 B.n515 585
R1416 B.n514 B.n513 585
R1417 B.n512 B.n511 585
R1418 B.n510 B.n509 585
R1419 B.n508 B.n507 585
R1420 B.n506 B.n505 585
R1421 B.n504 B.n503 585
R1422 B.n502 B.n501 585
R1423 B.n500 B.n499 585
R1424 B.n498 B.n497 585
R1425 B.n496 B.n495 585
R1426 B.n494 B.n493 585
R1427 B.n492 B.n491 585
R1428 B.n490 B.n489 585
R1429 B.n488 B.n487 585
R1430 B.n486 B.n485 585
R1431 B.n484 B.n483 585
R1432 B.n482 B.n481 585
R1433 B.n480 B.n479 585
R1434 B.n478 B.n477 585
R1435 B.n476 B.n475 585
R1436 B.n474 B.n473 585
R1437 B.n472 B.n471 585
R1438 B.n470 B.n469 585
R1439 B.n468 B.n467 585
R1440 B.n466 B.n465 585
R1441 B.n464 B.n463 585
R1442 B.n462 B.n461 585
R1443 B.n460 B.n459 585
R1444 B.n458 B.n457 585
R1445 B.n456 B.n455 585
R1446 B.n454 B.n453 585
R1447 B.n452 B.n451 585
R1448 B.n450 B.n449 585
R1449 B.n448 B.n447 585
R1450 B.n385 B.n384 585
R1451 B.n674 B.n673 585
R1452 B.n673 B.n672 585
R1453 B.n381 B.n380 585
R1454 B.n382 B.n381 585
R1455 B.n680 B.n679 585
R1456 B.n679 B.n678 585
R1457 B.n681 B.n379 585
R1458 B.n379 B.n377 585
R1459 B.n683 B.n682 585
R1460 B.n684 B.n683 585
R1461 B.n373 B.n372 585
R1462 B.n378 B.n373 585
R1463 B.n692 B.n691 585
R1464 B.n691 B.n690 585
R1465 B.n693 B.n371 585
R1466 B.n371 B.n370 585
R1467 B.n695 B.n694 585
R1468 B.n696 B.n695 585
R1469 B.n365 B.n364 585
R1470 B.n366 B.n365 585
R1471 B.n704 B.n703 585
R1472 B.n703 B.n702 585
R1473 B.n705 B.n363 585
R1474 B.n363 B.n362 585
R1475 B.n707 B.n706 585
R1476 B.n708 B.n707 585
R1477 B.n357 B.n356 585
R1478 B.n358 B.n357 585
R1479 B.n716 B.n715 585
R1480 B.n715 B.n714 585
R1481 B.n717 B.n355 585
R1482 B.n355 B.n354 585
R1483 B.n719 B.n718 585
R1484 B.n720 B.n719 585
R1485 B.n349 B.n348 585
R1486 B.n350 B.n349 585
R1487 B.n729 B.n728 585
R1488 B.n728 B.n727 585
R1489 B.n730 B.n347 585
R1490 B.n726 B.n347 585
R1491 B.n732 B.n731 585
R1492 B.n733 B.n732 585
R1493 B.n342 B.n341 585
R1494 B.n343 B.n342 585
R1495 B.n743 B.n742 585
R1496 B.n742 B.n741 585
R1497 B.n744 B.n340 585
R1498 B.n740 B.n340 585
R1499 B.n746 B.n745 585
R1500 B.n747 B.n746 585
R1501 B.n3 B.n0 585
R1502 B.n4 B.n3 585
R1503 B.n836 B.n1 585
R1504 B.n837 B.n836 585
R1505 B.n835 B.n834 585
R1506 B.n835 B.n8 585
R1507 B.n833 B.n9 585
R1508 B.n12 B.n9 585
R1509 B.n832 B.n831 585
R1510 B.n831 B.n830 585
R1511 B.n11 B.n10 585
R1512 B.n829 B.n11 585
R1513 B.n827 B.n826 585
R1514 B.n828 B.n827 585
R1515 B.n825 B.n16 585
R1516 B.n19 B.n16 585
R1517 B.n824 B.n823 585
R1518 B.n823 B.n822 585
R1519 B.n18 B.n17 585
R1520 B.n821 B.n18 585
R1521 B.n819 B.n818 585
R1522 B.n820 B.n819 585
R1523 B.n817 B.n24 585
R1524 B.n24 B.n23 585
R1525 B.n816 B.n815 585
R1526 B.n815 B.n814 585
R1527 B.n26 B.n25 585
R1528 B.n813 B.n26 585
R1529 B.n811 B.n810 585
R1530 B.n812 B.n811 585
R1531 B.n809 B.n31 585
R1532 B.n31 B.n30 585
R1533 B.n808 B.n807 585
R1534 B.n807 B.n806 585
R1535 B.n33 B.n32 585
R1536 B.n805 B.n33 585
R1537 B.n803 B.n802 585
R1538 B.n804 B.n803 585
R1539 B.n801 B.n38 585
R1540 B.n38 B.n37 585
R1541 B.n800 B.n799 585
R1542 B.n799 B.n798 585
R1543 B.n40 B.n39 585
R1544 B.n797 B.n40 585
R1545 B.n795 B.n794 585
R1546 B.n796 B.n795 585
R1547 B.n793 B.n45 585
R1548 B.n45 B.n44 585
R1549 B.n792 B.n791 585
R1550 B.n791 B.n790 585
R1551 B.n47 B.n46 585
R1552 B.n789 B.n47 585
R1553 B.n840 B.n839 585
R1554 B.n838 B.n2 585
R1555 B.n113 B.n47 530.939
R1556 B.n786 B.n49 530.939
R1557 B.n673 B.n383 530.939
R1558 B.n670 B.n381 530.939
R1559 B.n107 B.t10 367.334
R1560 B.n445 B.t18 367.334
R1561 B.n110 B.t13 367.334
R1562 B.n443 B.t21 367.334
R1563 B.n108 B.t11 344.062
R1564 B.n446 B.t17 344.062
R1565 B.n111 B.t14 344.062
R1566 B.n444 B.t20 344.062
R1567 B.n788 B.n787 256.663
R1568 B.n788 B.n105 256.663
R1569 B.n788 B.n104 256.663
R1570 B.n788 B.n103 256.663
R1571 B.n788 B.n102 256.663
R1572 B.n788 B.n101 256.663
R1573 B.n788 B.n100 256.663
R1574 B.n788 B.n99 256.663
R1575 B.n788 B.n98 256.663
R1576 B.n788 B.n97 256.663
R1577 B.n788 B.n96 256.663
R1578 B.n788 B.n95 256.663
R1579 B.n788 B.n94 256.663
R1580 B.n788 B.n93 256.663
R1581 B.n788 B.n92 256.663
R1582 B.n788 B.n91 256.663
R1583 B.n788 B.n90 256.663
R1584 B.n788 B.n89 256.663
R1585 B.n788 B.n88 256.663
R1586 B.n788 B.n87 256.663
R1587 B.n788 B.n86 256.663
R1588 B.n788 B.n85 256.663
R1589 B.n788 B.n84 256.663
R1590 B.n788 B.n83 256.663
R1591 B.n788 B.n82 256.663
R1592 B.n788 B.n81 256.663
R1593 B.n788 B.n80 256.663
R1594 B.n788 B.n79 256.663
R1595 B.n788 B.n78 256.663
R1596 B.n788 B.n77 256.663
R1597 B.n788 B.n76 256.663
R1598 B.n788 B.n75 256.663
R1599 B.n788 B.n74 256.663
R1600 B.n788 B.n73 256.663
R1601 B.n788 B.n72 256.663
R1602 B.n788 B.n71 256.663
R1603 B.n788 B.n70 256.663
R1604 B.n788 B.n69 256.663
R1605 B.n788 B.n68 256.663
R1606 B.n788 B.n67 256.663
R1607 B.n788 B.n66 256.663
R1608 B.n788 B.n65 256.663
R1609 B.n788 B.n64 256.663
R1610 B.n788 B.n63 256.663
R1611 B.n788 B.n62 256.663
R1612 B.n788 B.n61 256.663
R1613 B.n788 B.n60 256.663
R1614 B.n788 B.n59 256.663
R1615 B.n788 B.n58 256.663
R1616 B.n788 B.n57 256.663
R1617 B.n788 B.n56 256.663
R1618 B.n788 B.n55 256.663
R1619 B.n788 B.n54 256.663
R1620 B.n788 B.n53 256.663
R1621 B.n788 B.n52 256.663
R1622 B.n788 B.n51 256.663
R1623 B.n788 B.n50 256.663
R1624 B.n672 B.n671 256.663
R1625 B.n672 B.n386 256.663
R1626 B.n672 B.n387 256.663
R1627 B.n672 B.n388 256.663
R1628 B.n672 B.n389 256.663
R1629 B.n672 B.n390 256.663
R1630 B.n672 B.n391 256.663
R1631 B.n672 B.n392 256.663
R1632 B.n672 B.n393 256.663
R1633 B.n672 B.n394 256.663
R1634 B.n672 B.n395 256.663
R1635 B.n672 B.n396 256.663
R1636 B.n672 B.n397 256.663
R1637 B.n672 B.n398 256.663
R1638 B.n672 B.n399 256.663
R1639 B.n672 B.n400 256.663
R1640 B.n672 B.n401 256.663
R1641 B.n672 B.n402 256.663
R1642 B.n672 B.n403 256.663
R1643 B.n672 B.n404 256.663
R1644 B.n672 B.n405 256.663
R1645 B.n672 B.n406 256.663
R1646 B.n672 B.n407 256.663
R1647 B.n672 B.n408 256.663
R1648 B.n672 B.n409 256.663
R1649 B.n672 B.n410 256.663
R1650 B.n672 B.n411 256.663
R1651 B.n672 B.n412 256.663
R1652 B.n672 B.n413 256.663
R1653 B.n672 B.n414 256.663
R1654 B.n672 B.n415 256.663
R1655 B.n672 B.n416 256.663
R1656 B.n672 B.n417 256.663
R1657 B.n672 B.n418 256.663
R1658 B.n672 B.n419 256.663
R1659 B.n672 B.n420 256.663
R1660 B.n672 B.n421 256.663
R1661 B.n672 B.n422 256.663
R1662 B.n672 B.n423 256.663
R1663 B.n672 B.n424 256.663
R1664 B.n672 B.n425 256.663
R1665 B.n672 B.n426 256.663
R1666 B.n672 B.n427 256.663
R1667 B.n672 B.n428 256.663
R1668 B.n672 B.n429 256.663
R1669 B.n672 B.n430 256.663
R1670 B.n672 B.n431 256.663
R1671 B.n672 B.n432 256.663
R1672 B.n672 B.n433 256.663
R1673 B.n672 B.n434 256.663
R1674 B.n672 B.n435 256.663
R1675 B.n672 B.n436 256.663
R1676 B.n672 B.n437 256.663
R1677 B.n672 B.n438 256.663
R1678 B.n672 B.n439 256.663
R1679 B.n672 B.n440 256.663
R1680 B.n842 B.n841 256.663
R1681 B.n117 B.n116 163.367
R1682 B.n121 B.n120 163.367
R1683 B.n125 B.n124 163.367
R1684 B.n129 B.n128 163.367
R1685 B.n133 B.n132 163.367
R1686 B.n137 B.n136 163.367
R1687 B.n141 B.n140 163.367
R1688 B.n145 B.n144 163.367
R1689 B.n149 B.n148 163.367
R1690 B.n153 B.n152 163.367
R1691 B.n157 B.n156 163.367
R1692 B.n161 B.n160 163.367
R1693 B.n165 B.n164 163.367
R1694 B.n169 B.n168 163.367
R1695 B.n173 B.n172 163.367
R1696 B.n177 B.n176 163.367
R1697 B.n181 B.n180 163.367
R1698 B.n185 B.n184 163.367
R1699 B.n189 B.n188 163.367
R1700 B.n193 B.n192 163.367
R1701 B.n197 B.n196 163.367
R1702 B.n201 B.n200 163.367
R1703 B.n205 B.n204 163.367
R1704 B.n209 B.n208 163.367
R1705 B.n213 B.n212 163.367
R1706 B.n217 B.n216 163.367
R1707 B.n221 B.n220 163.367
R1708 B.n225 B.n224 163.367
R1709 B.n229 B.n228 163.367
R1710 B.n233 B.n232 163.367
R1711 B.n237 B.n236 163.367
R1712 B.n241 B.n240 163.367
R1713 B.n245 B.n244 163.367
R1714 B.n249 B.n248 163.367
R1715 B.n253 B.n252 163.367
R1716 B.n257 B.n256 163.367
R1717 B.n261 B.n260 163.367
R1718 B.n265 B.n264 163.367
R1719 B.n269 B.n268 163.367
R1720 B.n273 B.n272 163.367
R1721 B.n277 B.n276 163.367
R1722 B.n281 B.n280 163.367
R1723 B.n285 B.n284 163.367
R1724 B.n289 B.n288 163.367
R1725 B.n293 B.n292 163.367
R1726 B.n297 B.n296 163.367
R1727 B.n301 B.n300 163.367
R1728 B.n305 B.n304 163.367
R1729 B.n309 B.n308 163.367
R1730 B.n313 B.n312 163.367
R1731 B.n317 B.n316 163.367
R1732 B.n321 B.n320 163.367
R1733 B.n325 B.n324 163.367
R1734 B.n329 B.n328 163.367
R1735 B.n333 B.n332 163.367
R1736 B.n335 B.n106 163.367
R1737 B.n677 B.n383 163.367
R1738 B.n677 B.n376 163.367
R1739 B.n685 B.n376 163.367
R1740 B.n685 B.n374 163.367
R1741 B.n689 B.n374 163.367
R1742 B.n689 B.n369 163.367
R1743 B.n697 B.n369 163.367
R1744 B.n697 B.n367 163.367
R1745 B.n701 B.n367 163.367
R1746 B.n701 B.n361 163.367
R1747 B.n709 B.n361 163.367
R1748 B.n709 B.n359 163.367
R1749 B.n713 B.n359 163.367
R1750 B.n713 B.n353 163.367
R1751 B.n721 B.n353 163.367
R1752 B.n721 B.n351 163.367
R1753 B.n725 B.n351 163.367
R1754 B.n725 B.n346 163.367
R1755 B.n734 B.n346 163.367
R1756 B.n734 B.n344 163.367
R1757 B.n739 B.n344 163.367
R1758 B.n739 B.n339 163.367
R1759 B.n748 B.n339 163.367
R1760 B.n749 B.n748 163.367
R1761 B.n749 B.n5 163.367
R1762 B.n6 B.n5 163.367
R1763 B.n7 B.n6 163.367
R1764 B.n755 B.n7 163.367
R1765 B.n756 B.n755 163.367
R1766 B.n756 B.n13 163.367
R1767 B.n14 B.n13 163.367
R1768 B.n15 B.n14 163.367
R1769 B.n761 B.n15 163.367
R1770 B.n761 B.n20 163.367
R1771 B.n21 B.n20 163.367
R1772 B.n22 B.n21 163.367
R1773 B.n766 B.n22 163.367
R1774 B.n766 B.n27 163.367
R1775 B.n28 B.n27 163.367
R1776 B.n29 B.n28 163.367
R1777 B.n771 B.n29 163.367
R1778 B.n771 B.n34 163.367
R1779 B.n35 B.n34 163.367
R1780 B.n36 B.n35 163.367
R1781 B.n776 B.n36 163.367
R1782 B.n776 B.n41 163.367
R1783 B.n42 B.n41 163.367
R1784 B.n43 B.n42 163.367
R1785 B.n781 B.n43 163.367
R1786 B.n781 B.n48 163.367
R1787 B.n49 B.n48 163.367
R1788 B.n442 B.n441 163.367
R1789 B.n665 B.n441 163.367
R1790 B.n663 B.n662 163.367
R1791 B.n659 B.n658 163.367
R1792 B.n655 B.n654 163.367
R1793 B.n651 B.n650 163.367
R1794 B.n647 B.n646 163.367
R1795 B.n643 B.n642 163.367
R1796 B.n639 B.n638 163.367
R1797 B.n635 B.n634 163.367
R1798 B.n631 B.n630 163.367
R1799 B.n627 B.n626 163.367
R1800 B.n623 B.n622 163.367
R1801 B.n619 B.n618 163.367
R1802 B.n615 B.n614 163.367
R1803 B.n611 B.n610 163.367
R1804 B.n607 B.n606 163.367
R1805 B.n603 B.n602 163.367
R1806 B.n599 B.n598 163.367
R1807 B.n595 B.n594 163.367
R1808 B.n591 B.n590 163.367
R1809 B.n587 B.n586 163.367
R1810 B.n583 B.n582 163.367
R1811 B.n579 B.n578 163.367
R1812 B.n575 B.n574 163.367
R1813 B.n571 B.n570 163.367
R1814 B.n566 B.n565 163.367
R1815 B.n562 B.n561 163.367
R1816 B.n558 B.n557 163.367
R1817 B.n554 B.n553 163.367
R1818 B.n550 B.n549 163.367
R1819 B.n545 B.n544 163.367
R1820 B.n541 B.n540 163.367
R1821 B.n537 B.n536 163.367
R1822 B.n533 B.n532 163.367
R1823 B.n529 B.n528 163.367
R1824 B.n525 B.n524 163.367
R1825 B.n521 B.n520 163.367
R1826 B.n517 B.n516 163.367
R1827 B.n513 B.n512 163.367
R1828 B.n509 B.n508 163.367
R1829 B.n505 B.n504 163.367
R1830 B.n501 B.n500 163.367
R1831 B.n497 B.n496 163.367
R1832 B.n493 B.n492 163.367
R1833 B.n489 B.n488 163.367
R1834 B.n485 B.n484 163.367
R1835 B.n481 B.n480 163.367
R1836 B.n477 B.n476 163.367
R1837 B.n473 B.n472 163.367
R1838 B.n469 B.n468 163.367
R1839 B.n465 B.n464 163.367
R1840 B.n461 B.n460 163.367
R1841 B.n457 B.n456 163.367
R1842 B.n453 B.n452 163.367
R1843 B.n449 B.n448 163.367
R1844 B.n673 B.n385 163.367
R1845 B.n679 B.n381 163.367
R1846 B.n679 B.n379 163.367
R1847 B.n683 B.n379 163.367
R1848 B.n683 B.n373 163.367
R1849 B.n691 B.n373 163.367
R1850 B.n691 B.n371 163.367
R1851 B.n695 B.n371 163.367
R1852 B.n695 B.n365 163.367
R1853 B.n703 B.n365 163.367
R1854 B.n703 B.n363 163.367
R1855 B.n707 B.n363 163.367
R1856 B.n707 B.n357 163.367
R1857 B.n715 B.n357 163.367
R1858 B.n715 B.n355 163.367
R1859 B.n719 B.n355 163.367
R1860 B.n719 B.n349 163.367
R1861 B.n728 B.n349 163.367
R1862 B.n728 B.n347 163.367
R1863 B.n732 B.n347 163.367
R1864 B.n732 B.n342 163.367
R1865 B.n742 B.n342 163.367
R1866 B.n742 B.n340 163.367
R1867 B.n746 B.n340 163.367
R1868 B.n746 B.n3 163.367
R1869 B.n840 B.n3 163.367
R1870 B.n836 B.n2 163.367
R1871 B.n836 B.n835 163.367
R1872 B.n835 B.n9 163.367
R1873 B.n831 B.n9 163.367
R1874 B.n831 B.n11 163.367
R1875 B.n827 B.n11 163.367
R1876 B.n827 B.n16 163.367
R1877 B.n823 B.n16 163.367
R1878 B.n823 B.n18 163.367
R1879 B.n819 B.n18 163.367
R1880 B.n819 B.n24 163.367
R1881 B.n815 B.n24 163.367
R1882 B.n815 B.n26 163.367
R1883 B.n811 B.n26 163.367
R1884 B.n811 B.n31 163.367
R1885 B.n807 B.n31 163.367
R1886 B.n807 B.n33 163.367
R1887 B.n803 B.n33 163.367
R1888 B.n803 B.n38 163.367
R1889 B.n799 B.n38 163.367
R1890 B.n799 B.n40 163.367
R1891 B.n795 B.n40 163.367
R1892 B.n795 B.n45 163.367
R1893 B.n791 B.n45 163.367
R1894 B.n791 B.n47 163.367
R1895 B.n672 B.n382 74.3712
R1896 B.n789 B.n788 74.3712
R1897 B.n113 B.n50 71.676
R1898 B.n117 B.n51 71.676
R1899 B.n121 B.n52 71.676
R1900 B.n125 B.n53 71.676
R1901 B.n129 B.n54 71.676
R1902 B.n133 B.n55 71.676
R1903 B.n137 B.n56 71.676
R1904 B.n141 B.n57 71.676
R1905 B.n145 B.n58 71.676
R1906 B.n149 B.n59 71.676
R1907 B.n153 B.n60 71.676
R1908 B.n157 B.n61 71.676
R1909 B.n161 B.n62 71.676
R1910 B.n165 B.n63 71.676
R1911 B.n169 B.n64 71.676
R1912 B.n173 B.n65 71.676
R1913 B.n177 B.n66 71.676
R1914 B.n181 B.n67 71.676
R1915 B.n185 B.n68 71.676
R1916 B.n189 B.n69 71.676
R1917 B.n193 B.n70 71.676
R1918 B.n197 B.n71 71.676
R1919 B.n201 B.n72 71.676
R1920 B.n205 B.n73 71.676
R1921 B.n209 B.n74 71.676
R1922 B.n213 B.n75 71.676
R1923 B.n217 B.n76 71.676
R1924 B.n221 B.n77 71.676
R1925 B.n225 B.n78 71.676
R1926 B.n229 B.n79 71.676
R1927 B.n233 B.n80 71.676
R1928 B.n237 B.n81 71.676
R1929 B.n241 B.n82 71.676
R1930 B.n245 B.n83 71.676
R1931 B.n249 B.n84 71.676
R1932 B.n253 B.n85 71.676
R1933 B.n257 B.n86 71.676
R1934 B.n261 B.n87 71.676
R1935 B.n265 B.n88 71.676
R1936 B.n269 B.n89 71.676
R1937 B.n273 B.n90 71.676
R1938 B.n277 B.n91 71.676
R1939 B.n281 B.n92 71.676
R1940 B.n285 B.n93 71.676
R1941 B.n289 B.n94 71.676
R1942 B.n293 B.n95 71.676
R1943 B.n297 B.n96 71.676
R1944 B.n301 B.n97 71.676
R1945 B.n305 B.n98 71.676
R1946 B.n309 B.n99 71.676
R1947 B.n313 B.n100 71.676
R1948 B.n317 B.n101 71.676
R1949 B.n321 B.n102 71.676
R1950 B.n325 B.n103 71.676
R1951 B.n329 B.n104 71.676
R1952 B.n333 B.n105 71.676
R1953 B.n787 B.n106 71.676
R1954 B.n787 B.n786 71.676
R1955 B.n335 B.n105 71.676
R1956 B.n332 B.n104 71.676
R1957 B.n328 B.n103 71.676
R1958 B.n324 B.n102 71.676
R1959 B.n320 B.n101 71.676
R1960 B.n316 B.n100 71.676
R1961 B.n312 B.n99 71.676
R1962 B.n308 B.n98 71.676
R1963 B.n304 B.n97 71.676
R1964 B.n300 B.n96 71.676
R1965 B.n296 B.n95 71.676
R1966 B.n292 B.n94 71.676
R1967 B.n288 B.n93 71.676
R1968 B.n284 B.n92 71.676
R1969 B.n280 B.n91 71.676
R1970 B.n276 B.n90 71.676
R1971 B.n272 B.n89 71.676
R1972 B.n268 B.n88 71.676
R1973 B.n264 B.n87 71.676
R1974 B.n260 B.n86 71.676
R1975 B.n256 B.n85 71.676
R1976 B.n252 B.n84 71.676
R1977 B.n248 B.n83 71.676
R1978 B.n244 B.n82 71.676
R1979 B.n240 B.n81 71.676
R1980 B.n236 B.n80 71.676
R1981 B.n232 B.n79 71.676
R1982 B.n228 B.n78 71.676
R1983 B.n224 B.n77 71.676
R1984 B.n220 B.n76 71.676
R1985 B.n216 B.n75 71.676
R1986 B.n212 B.n74 71.676
R1987 B.n208 B.n73 71.676
R1988 B.n204 B.n72 71.676
R1989 B.n200 B.n71 71.676
R1990 B.n196 B.n70 71.676
R1991 B.n192 B.n69 71.676
R1992 B.n188 B.n68 71.676
R1993 B.n184 B.n67 71.676
R1994 B.n180 B.n66 71.676
R1995 B.n176 B.n65 71.676
R1996 B.n172 B.n64 71.676
R1997 B.n168 B.n63 71.676
R1998 B.n164 B.n62 71.676
R1999 B.n160 B.n61 71.676
R2000 B.n156 B.n60 71.676
R2001 B.n152 B.n59 71.676
R2002 B.n148 B.n58 71.676
R2003 B.n144 B.n57 71.676
R2004 B.n140 B.n56 71.676
R2005 B.n136 B.n55 71.676
R2006 B.n132 B.n54 71.676
R2007 B.n128 B.n53 71.676
R2008 B.n124 B.n52 71.676
R2009 B.n120 B.n51 71.676
R2010 B.n116 B.n50 71.676
R2011 B.n671 B.n670 71.676
R2012 B.n665 B.n386 71.676
R2013 B.n662 B.n387 71.676
R2014 B.n658 B.n388 71.676
R2015 B.n654 B.n389 71.676
R2016 B.n650 B.n390 71.676
R2017 B.n646 B.n391 71.676
R2018 B.n642 B.n392 71.676
R2019 B.n638 B.n393 71.676
R2020 B.n634 B.n394 71.676
R2021 B.n630 B.n395 71.676
R2022 B.n626 B.n396 71.676
R2023 B.n622 B.n397 71.676
R2024 B.n618 B.n398 71.676
R2025 B.n614 B.n399 71.676
R2026 B.n610 B.n400 71.676
R2027 B.n606 B.n401 71.676
R2028 B.n602 B.n402 71.676
R2029 B.n598 B.n403 71.676
R2030 B.n594 B.n404 71.676
R2031 B.n590 B.n405 71.676
R2032 B.n586 B.n406 71.676
R2033 B.n582 B.n407 71.676
R2034 B.n578 B.n408 71.676
R2035 B.n574 B.n409 71.676
R2036 B.n570 B.n410 71.676
R2037 B.n565 B.n411 71.676
R2038 B.n561 B.n412 71.676
R2039 B.n557 B.n413 71.676
R2040 B.n553 B.n414 71.676
R2041 B.n549 B.n415 71.676
R2042 B.n544 B.n416 71.676
R2043 B.n540 B.n417 71.676
R2044 B.n536 B.n418 71.676
R2045 B.n532 B.n419 71.676
R2046 B.n528 B.n420 71.676
R2047 B.n524 B.n421 71.676
R2048 B.n520 B.n422 71.676
R2049 B.n516 B.n423 71.676
R2050 B.n512 B.n424 71.676
R2051 B.n508 B.n425 71.676
R2052 B.n504 B.n426 71.676
R2053 B.n500 B.n427 71.676
R2054 B.n496 B.n428 71.676
R2055 B.n492 B.n429 71.676
R2056 B.n488 B.n430 71.676
R2057 B.n484 B.n431 71.676
R2058 B.n480 B.n432 71.676
R2059 B.n476 B.n433 71.676
R2060 B.n472 B.n434 71.676
R2061 B.n468 B.n435 71.676
R2062 B.n464 B.n436 71.676
R2063 B.n460 B.n437 71.676
R2064 B.n456 B.n438 71.676
R2065 B.n452 B.n439 71.676
R2066 B.n448 B.n440 71.676
R2067 B.n671 B.n442 71.676
R2068 B.n663 B.n386 71.676
R2069 B.n659 B.n387 71.676
R2070 B.n655 B.n388 71.676
R2071 B.n651 B.n389 71.676
R2072 B.n647 B.n390 71.676
R2073 B.n643 B.n391 71.676
R2074 B.n639 B.n392 71.676
R2075 B.n635 B.n393 71.676
R2076 B.n631 B.n394 71.676
R2077 B.n627 B.n395 71.676
R2078 B.n623 B.n396 71.676
R2079 B.n619 B.n397 71.676
R2080 B.n615 B.n398 71.676
R2081 B.n611 B.n399 71.676
R2082 B.n607 B.n400 71.676
R2083 B.n603 B.n401 71.676
R2084 B.n599 B.n402 71.676
R2085 B.n595 B.n403 71.676
R2086 B.n591 B.n404 71.676
R2087 B.n587 B.n405 71.676
R2088 B.n583 B.n406 71.676
R2089 B.n579 B.n407 71.676
R2090 B.n575 B.n408 71.676
R2091 B.n571 B.n409 71.676
R2092 B.n566 B.n410 71.676
R2093 B.n562 B.n411 71.676
R2094 B.n558 B.n412 71.676
R2095 B.n554 B.n413 71.676
R2096 B.n550 B.n414 71.676
R2097 B.n545 B.n415 71.676
R2098 B.n541 B.n416 71.676
R2099 B.n537 B.n417 71.676
R2100 B.n533 B.n418 71.676
R2101 B.n529 B.n419 71.676
R2102 B.n525 B.n420 71.676
R2103 B.n521 B.n421 71.676
R2104 B.n517 B.n422 71.676
R2105 B.n513 B.n423 71.676
R2106 B.n509 B.n424 71.676
R2107 B.n505 B.n425 71.676
R2108 B.n501 B.n426 71.676
R2109 B.n497 B.n427 71.676
R2110 B.n493 B.n428 71.676
R2111 B.n489 B.n429 71.676
R2112 B.n485 B.n430 71.676
R2113 B.n481 B.n431 71.676
R2114 B.n477 B.n432 71.676
R2115 B.n473 B.n433 71.676
R2116 B.n469 B.n434 71.676
R2117 B.n465 B.n435 71.676
R2118 B.n461 B.n436 71.676
R2119 B.n457 B.n437 71.676
R2120 B.n453 B.n438 71.676
R2121 B.n449 B.n439 71.676
R2122 B.n440 B.n385 71.676
R2123 B.n841 B.n840 71.676
R2124 B.n841 B.n2 71.676
R2125 B.n112 B.n111 59.5399
R2126 B.n109 B.n108 59.5399
R2127 B.n547 B.n446 59.5399
R2128 B.n568 B.n444 59.5399
R2129 B.n678 B.n382 35.8672
R2130 B.n678 B.n377 35.8672
R2131 B.n684 B.n377 35.8672
R2132 B.n684 B.n378 35.8672
R2133 B.n690 B.n370 35.8672
R2134 B.n696 B.n370 35.8672
R2135 B.n696 B.n366 35.8672
R2136 B.n702 B.n366 35.8672
R2137 B.n702 B.n362 35.8672
R2138 B.n708 B.n362 35.8672
R2139 B.n714 B.n358 35.8672
R2140 B.n714 B.n354 35.8672
R2141 B.n720 B.n354 35.8672
R2142 B.n727 B.n350 35.8672
R2143 B.n727 B.n726 35.8672
R2144 B.n733 B.n343 35.8672
R2145 B.n741 B.n343 35.8672
R2146 B.n741 B.n740 35.8672
R2147 B.n747 B.n4 35.8672
R2148 B.n839 B.n4 35.8672
R2149 B.n839 B.n838 35.8672
R2150 B.n838 B.n837 35.8672
R2151 B.n837 B.n8 35.8672
R2152 B.n830 B.n12 35.8672
R2153 B.n830 B.n829 35.8672
R2154 B.n829 B.n828 35.8672
R2155 B.n822 B.n19 35.8672
R2156 B.n822 B.n821 35.8672
R2157 B.n820 B.n23 35.8672
R2158 B.n814 B.n23 35.8672
R2159 B.n814 B.n813 35.8672
R2160 B.n812 B.n30 35.8672
R2161 B.n806 B.n30 35.8672
R2162 B.n806 B.n805 35.8672
R2163 B.n805 B.n804 35.8672
R2164 B.n804 B.n37 35.8672
R2165 B.n798 B.n37 35.8672
R2166 B.n797 B.n796 35.8672
R2167 B.n796 B.n44 35.8672
R2168 B.n790 B.n44 35.8672
R2169 B.n790 B.n789 35.8672
R2170 B.n669 B.n380 34.4981
R2171 B.n675 B.n674 34.4981
R2172 B.n785 B.n784 34.4981
R2173 B.n114 B.n46 34.4981
R2174 B.t0 B.n350 33.2299
R2175 B.n821 B.t5 33.2299
R2176 B.n747 B.t7 31.1201
R2177 B.t4 B.n8 31.1201
R2178 B.n378 B.t16 29.0103
R2179 B.t9 B.n797 29.0103
R2180 B.n111 B.n110 23.2732
R2181 B.n108 B.n107 23.2732
R2182 B.n446 B.n445 23.2732
R2183 B.n444 B.n443 23.2732
R2184 B.n726 B.t6 21.626
R2185 B.n19 B.t2 21.626
R2186 B.n708 B.t3 19.5162
R2187 B.t1 B.n812 19.5162
R2188 B B.n842 18.0485
R2189 B.t3 B.n358 16.3515
R2190 B.n813 B.t1 16.3515
R2191 B.n733 B.t6 14.2417
R2192 B.n828 B.t2 14.2417
R2193 B.n680 B.n380 10.6151
R2194 B.n681 B.n680 10.6151
R2195 B.n682 B.n681 10.6151
R2196 B.n682 B.n372 10.6151
R2197 B.n692 B.n372 10.6151
R2198 B.n693 B.n692 10.6151
R2199 B.n694 B.n693 10.6151
R2200 B.n694 B.n364 10.6151
R2201 B.n704 B.n364 10.6151
R2202 B.n705 B.n704 10.6151
R2203 B.n706 B.n705 10.6151
R2204 B.n706 B.n356 10.6151
R2205 B.n716 B.n356 10.6151
R2206 B.n717 B.n716 10.6151
R2207 B.n718 B.n717 10.6151
R2208 B.n718 B.n348 10.6151
R2209 B.n729 B.n348 10.6151
R2210 B.n730 B.n729 10.6151
R2211 B.n731 B.n730 10.6151
R2212 B.n731 B.n341 10.6151
R2213 B.n743 B.n341 10.6151
R2214 B.n744 B.n743 10.6151
R2215 B.n745 B.n744 10.6151
R2216 B.n745 B.n0 10.6151
R2217 B.n669 B.n668 10.6151
R2218 B.n668 B.n667 10.6151
R2219 B.n667 B.n666 10.6151
R2220 B.n666 B.n664 10.6151
R2221 B.n664 B.n661 10.6151
R2222 B.n661 B.n660 10.6151
R2223 B.n660 B.n657 10.6151
R2224 B.n657 B.n656 10.6151
R2225 B.n656 B.n653 10.6151
R2226 B.n653 B.n652 10.6151
R2227 B.n652 B.n649 10.6151
R2228 B.n649 B.n648 10.6151
R2229 B.n648 B.n645 10.6151
R2230 B.n645 B.n644 10.6151
R2231 B.n644 B.n641 10.6151
R2232 B.n641 B.n640 10.6151
R2233 B.n640 B.n637 10.6151
R2234 B.n637 B.n636 10.6151
R2235 B.n636 B.n633 10.6151
R2236 B.n633 B.n632 10.6151
R2237 B.n632 B.n629 10.6151
R2238 B.n629 B.n628 10.6151
R2239 B.n628 B.n625 10.6151
R2240 B.n625 B.n624 10.6151
R2241 B.n624 B.n621 10.6151
R2242 B.n621 B.n620 10.6151
R2243 B.n620 B.n617 10.6151
R2244 B.n617 B.n616 10.6151
R2245 B.n616 B.n613 10.6151
R2246 B.n613 B.n612 10.6151
R2247 B.n612 B.n609 10.6151
R2248 B.n609 B.n608 10.6151
R2249 B.n608 B.n605 10.6151
R2250 B.n605 B.n604 10.6151
R2251 B.n604 B.n601 10.6151
R2252 B.n601 B.n600 10.6151
R2253 B.n600 B.n597 10.6151
R2254 B.n597 B.n596 10.6151
R2255 B.n596 B.n593 10.6151
R2256 B.n593 B.n592 10.6151
R2257 B.n592 B.n589 10.6151
R2258 B.n589 B.n588 10.6151
R2259 B.n588 B.n585 10.6151
R2260 B.n585 B.n584 10.6151
R2261 B.n584 B.n581 10.6151
R2262 B.n581 B.n580 10.6151
R2263 B.n580 B.n577 10.6151
R2264 B.n577 B.n576 10.6151
R2265 B.n576 B.n573 10.6151
R2266 B.n573 B.n572 10.6151
R2267 B.n572 B.n569 10.6151
R2268 B.n567 B.n564 10.6151
R2269 B.n564 B.n563 10.6151
R2270 B.n563 B.n560 10.6151
R2271 B.n560 B.n559 10.6151
R2272 B.n559 B.n556 10.6151
R2273 B.n556 B.n555 10.6151
R2274 B.n555 B.n552 10.6151
R2275 B.n552 B.n551 10.6151
R2276 B.n551 B.n548 10.6151
R2277 B.n546 B.n543 10.6151
R2278 B.n543 B.n542 10.6151
R2279 B.n542 B.n539 10.6151
R2280 B.n539 B.n538 10.6151
R2281 B.n538 B.n535 10.6151
R2282 B.n535 B.n534 10.6151
R2283 B.n534 B.n531 10.6151
R2284 B.n531 B.n530 10.6151
R2285 B.n530 B.n527 10.6151
R2286 B.n527 B.n526 10.6151
R2287 B.n526 B.n523 10.6151
R2288 B.n523 B.n522 10.6151
R2289 B.n522 B.n519 10.6151
R2290 B.n519 B.n518 10.6151
R2291 B.n518 B.n515 10.6151
R2292 B.n515 B.n514 10.6151
R2293 B.n514 B.n511 10.6151
R2294 B.n511 B.n510 10.6151
R2295 B.n510 B.n507 10.6151
R2296 B.n507 B.n506 10.6151
R2297 B.n506 B.n503 10.6151
R2298 B.n503 B.n502 10.6151
R2299 B.n502 B.n499 10.6151
R2300 B.n499 B.n498 10.6151
R2301 B.n498 B.n495 10.6151
R2302 B.n495 B.n494 10.6151
R2303 B.n494 B.n491 10.6151
R2304 B.n491 B.n490 10.6151
R2305 B.n490 B.n487 10.6151
R2306 B.n487 B.n486 10.6151
R2307 B.n486 B.n483 10.6151
R2308 B.n483 B.n482 10.6151
R2309 B.n482 B.n479 10.6151
R2310 B.n479 B.n478 10.6151
R2311 B.n478 B.n475 10.6151
R2312 B.n475 B.n474 10.6151
R2313 B.n474 B.n471 10.6151
R2314 B.n471 B.n470 10.6151
R2315 B.n470 B.n467 10.6151
R2316 B.n467 B.n466 10.6151
R2317 B.n466 B.n463 10.6151
R2318 B.n463 B.n462 10.6151
R2319 B.n462 B.n459 10.6151
R2320 B.n459 B.n458 10.6151
R2321 B.n458 B.n455 10.6151
R2322 B.n455 B.n454 10.6151
R2323 B.n454 B.n451 10.6151
R2324 B.n451 B.n450 10.6151
R2325 B.n450 B.n447 10.6151
R2326 B.n447 B.n384 10.6151
R2327 B.n674 B.n384 10.6151
R2328 B.n676 B.n675 10.6151
R2329 B.n676 B.n375 10.6151
R2330 B.n686 B.n375 10.6151
R2331 B.n687 B.n686 10.6151
R2332 B.n688 B.n687 10.6151
R2333 B.n688 B.n368 10.6151
R2334 B.n698 B.n368 10.6151
R2335 B.n699 B.n698 10.6151
R2336 B.n700 B.n699 10.6151
R2337 B.n700 B.n360 10.6151
R2338 B.n710 B.n360 10.6151
R2339 B.n711 B.n710 10.6151
R2340 B.n712 B.n711 10.6151
R2341 B.n712 B.n352 10.6151
R2342 B.n722 B.n352 10.6151
R2343 B.n723 B.n722 10.6151
R2344 B.n724 B.n723 10.6151
R2345 B.n724 B.n345 10.6151
R2346 B.n735 B.n345 10.6151
R2347 B.n736 B.n735 10.6151
R2348 B.n738 B.n736 10.6151
R2349 B.n738 B.n737 10.6151
R2350 B.n737 B.n338 10.6151
R2351 B.n750 B.n338 10.6151
R2352 B.n751 B.n750 10.6151
R2353 B.n752 B.n751 10.6151
R2354 B.n753 B.n752 10.6151
R2355 B.n754 B.n753 10.6151
R2356 B.n757 B.n754 10.6151
R2357 B.n758 B.n757 10.6151
R2358 B.n759 B.n758 10.6151
R2359 B.n760 B.n759 10.6151
R2360 B.n762 B.n760 10.6151
R2361 B.n763 B.n762 10.6151
R2362 B.n764 B.n763 10.6151
R2363 B.n765 B.n764 10.6151
R2364 B.n767 B.n765 10.6151
R2365 B.n768 B.n767 10.6151
R2366 B.n769 B.n768 10.6151
R2367 B.n770 B.n769 10.6151
R2368 B.n772 B.n770 10.6151
R2369 B.n773 B.n772 10.6151
R2370 B.n774 B.n773 10.6151
R2371 B.n775 B.n774 10.6151
R2372 B.n777 B.n775 10.6151
R2373 B.n778 B.n777 10.6151
R2374 B.n779 B.n778 10.6151
R2375 B.n780 B.n779 10.6151
R2376 B.n782 B.n780 10.6151
R2377 B.n783 B.n782 10.6151
R2378 B.n784 B.n783 10.6151
R2379 B.n834 B.n1 10.6151
R2380 B.n834 B.n833 10.6151
R2381 B.n833 B.n832 10.6151
R2382 B.n832 B.n10 10.6151
R2383 B.n826 B.n10 10.6151
R2384 B.n826 B.n825 10.6151
R2385 B.n825 B.n824 10.6151
R2386 B.n824 B.n17 10.6151
R2387 B.n818 B.n17 10.6151
R2388 B.n818 B.n817 10.6151
R2389 B.n817 B.n816 10.6151
R2390 B.n816 B.n25 10.6151
R2391 B.n810 B.n25 10.6151
R2392 B.n810 B.n809 10.6151
R2393 B.n809 B.n808 10.6151
R2394 B.n808 B.n32 10.6151
R2395 B.n802 B.n32 10.6151
R2396 B.n802 B.n801 10.6151
R2397 B.n801 B.n800 10.6151
R2398 B.n800 B.n39 10.6151
R2399 B.n794 B.n39 10.6151
R2400 B.n794 B.n793 10.6151
R2401 B.n793 B.n792 10.6151
R2402 B.n792 B.n46 10.6151
R2403 B.n115 B.n114 10.6151
R2404 B.n118 B.n115 10.6151
R2405 B.n119 B.n118 10.6151
R2406 B.n122 B.n119 10.6151
R2407 B.n123 B.n122 10.6151
R2408 B.n126 B.n123 10.6151
R2409 B.n127 B.n126 10.6151
R2410 B.n130 B.n127 10.6151
R2411 B.n131 B.n130 10.6151
R2412 B.n134 B.n131 10.6151
R2413 B.n135 B.n134 10.6151
R2414 B.n138 B.n135 10.6151
R2415 B.n139 B.n138 10.6151
R2416 B.n142 B.n139 10.6151
R2417 B.n143 B.n142 10.6151
R2418 B.n146 B.n143 10.6151
R2419 B.n147 B.n146 10.6151
R2420 B.n150 B.n147 10.6151
R2421 B.n151 B.n150 10.6151
R2422 B.n154 B.n151 10.6151
R2423 B.n155 B.n154 10.6151
R2424 B.n158 B.n155 10.6151
R2425 B.n159 B.n158 10.6151
R2426 B.n162 B.n159 10.6151
R2427 B.n163 B.n162 10.6151
R2428 B.n166 B.n163 10.6151
R2429 B.n167 B.n166 10.6151
R2430 B.n170 B.n167 10.6151
R2431 B.n171 B.n170 10.6151
R2432 B.n174 B.n171 10.6151
R2433 B.n175 B.n174 10.6151
R2434 B.n178 B.n175 10.6151
R2435 B.n179 B.n178 10.6151
R2436 B.n182 B.n179 10.6151
R2437 B.n183 B.n182 10.6151
R2438 B.n186 B.n183 10.6151
R2439 B.n187 B.n186 10.6151
R2440 B.n190 B.n187 10.6151
R2441 B.n191 B.n190 10.6151
R2442 B.n194 B.n191 10.6151
R2443 B.n195 B.n194 10.6151
R2444 B.n198 B.n195 10.6151
R2445 B.n199 B.n198 10.6151
R2446 B.n202 B.n199 10.6151
R2447 B.n203 B.n202 10.6151
R2448 B.n206 B.n203 10.6151
R2449 B.n207 B.n206 10.6151
R2450 B.n210 B.n207 10.6151
R2451 B.n211 B.n210 10.6151
R2452 B.n214 B.n211 10.6151
R2453 B.n215 B.n214 10.6151
R2454 B.n219 B.n218 10.6151
R2455 B.n222 B.n219 10.6151
R2456 B.n223 B.n222 10.6151
R2457 B.n226 B.n223 10.6151
R2458 B.n227 B.n226 10.6151
R2459 B.n230 B.n227 10.6151
R2460 B.n231 B.n230 10.6151
R2461 B.n234 B.n231 10.6151
R2462 B.n235 B.n234 10.6151
R2463 B.n239 B.n238 10.6151
R2464 B.n242 B.n239 10.6151
R2465 B.n243 B.n242 10.6151
R2466 B.n246 B.n243 10.6151
R2467 B.n247 B.n246 10.6151
R2468 B.n250 B.n247 10.6151
R2469 B.n251 B.n250 10.6151
R2470 B.n254 B.n251 10.6151
R2471 B.n255 B.n254 10.6151
R2472 B.n258 B.n255 10.6151
R2473 B.n259 B.n258 10.6151
R2474 B.n262 B.n259 10.6151
R2475 B.n263 B.n262 10.6151
R2476 B.n266 B.n263 10.6151
R2477 B.n267 B.n266 10.6151
R2478 B.n270 B.n267 10.6151
R2479 B.n271 B.n270 10.6151
R2480 B.n274 B.n271 10.6151
R2481 B.n275 B.n274 10.6151
R2482 B.n278 B.n275 10.6151
R2483 B.n279 B.n278 10.6151
R2484 B.n282 B.n279 10.6151
R2485 B.n283 B.n282 10.6151
R2486 B.n286 B.n283 10.6151
R2487 B.n287 B.n286 10.6151
R2488 B.n290 B.n287 10.6151
R2489 B.n291 B.n290 10.6151
R2490 B.n294 B.n291 10.6151
R2491 B.n295 B.n294 10.6151
R2492 B.n298 B.n295 10.6151
R2493 B.n299 B.n298 10.6151
R2494 B.n302 B.n299 10.6151
R2495 B.n303 B.n302 10.6151
R2496 B.n306 B.n303 10.6151
R2497 B.n307 B.n306 10.6151
R2498 B.n310 B.n307 10.6151
R2499 B.n311 B.n310 10.6151
R2500 B.n314 B.n311 10.6151
R2501 B.n315 B.n314 10.6151
R2502 B.n318 B.n315 10.6151
R2503 B.n319 B.n318 10.6151
R2504 B.n322 B.n319 10.6151
R2505 B.n323 B.n322 10.6151
R2506 B.n326 B.n323 10.6151
R2507 B.n327 B.n326 10.6151
R2508 B.n330 B.n327 10.6151
R2509 B.n331 B.n330 10.6151
R2510 B.n334 B.n331 10.6151
R2511 B.n336 B.n334 10.6151
R2512 B.n337 B.n336 10.6151
R2513 B.n785 B.n337 10.6151
R2514 B.n569 B.n568 9.36635
R2515 B.n547 B.n546 9.36635
R2516 B.n215 B.n112 9.36635
R2517 B.n238 B.n109 9.36635
R2518 B.n842 B.n0 8.11757
R2519 B.n842 B.n1 8.11757
R2520 B.n690 B.t16 6.85737
R2521 B.n798 B.t9 6.85737
R2522 B.n740 B.t7 4.74756
R2523 B.n12 B.t4 4.74756
R2524 B.n720 B.t0 2.63776
R2525 B.t5 B.n820 2.63776
R2526 B.n568 B.n567 1.24928
R2527 B.n548 B.n547 1.24928
R2528 B.n218 B.n112 1.24928
R2529 B.n235 B.n109 1.24928
R2530 VP.n7 VP.t1 498.808
R2531 VP.n17 VP.t3 476.738
R2532 VP.n29 VP.t4 476.738
R2533 VP.n15 VP.t6 476.738
R2534 VP.n22 VP.t5 431.584
R2535 VP.n1 VP.t2 431.584
R2536 VP.n5 VP.t0 431.584
R2537 VP.n8 VP.t7 431.584
R2538 VP.n30 VP.n29 161.3
R2539 VP.n9 VP.n6 161.3
R2540 VP.n11 VP.n10 161.3
R2541 VP.n13 VP.n12 161.3
R2542 VP.n14 VP.n4 161.3
R2543 VP.n16 VP.n15 161.3
R2544 VP.n28 VP.n0 161.3
R2545 VP.n27 VP.n26 161.3
R2546 VP.n25 VP.n24 161.3
R2547 VP.n23 VP.n2 161.3
R2548 VP.n21 VP.n20 161.3
R2549 VP.n19 VP.n3 161.3
R2550 VP.n18 VP.n17 161.3
R2551 VP.n24 VP.n23 56.5617
R2552 VP.n10 VP.n9 56.5617
R2553 VP.n18 VP.n16 45.546
R2554 VP.n21 VP.n3 45.4209
R2555 VP.n28 VP.n27 45.4209
R2556 VP.n14 VP.n13 45.4209
R2557 VP.n7 VP.n6 42.7264
R2558 VP.n8 VP.n7 36.9171
R2559 VP.n23 VP.n22 17.2148
R2560 VP.n24 VP.n1 17.2148
R2561 VP.n10 VP.n5 17.2148
R2562 VP.n9 VP.n8 17.2148
R2563 VP.n17 VP.n3 16.7975
R2564 VP.n29 VP.n28 16.7975
R2565 VP.n15 VP.n14 16.7975
R2566 VP.n22 VP.n21 7.37805
R2567 VP.n27 VP.n1 7.37805
R2568 VP.n13 VP.n5 7.37805
R2569 VP.n11 VP.n6 0.189894
R2570 VP.n12 VP.n11 0.189894
R2571 VP.n12 VP.n4 0.189894
R2572 VP.n16 VP.n4 0.189894
R2573 VP.n19 VP.n18 0.189894
R2574 VP.n20 VP.n19 0.189894
R2575 VP.n20 VP.n2 0.189894
R2576 VP.n25 VP.n2 0.189894
R2577 VP.n26 VP.n25 0.189894
R2578 VP.n26 VP.n0 0.189894
R2579 VP.n30 VP.n0 0.189894
R2580 VP VP.n30 0.0516364
R2581 VDD1 VDD1.n0 65.6847
R2582 VDD1.n3 VDD1.n2 65.571
R2583 VDD1.n3 VDD1.n1 65.571
R2584 VDD1.n5 VDD1.n4 65.1091
R2585 VDD1.n5 VDD1.n3 42.3845
R2586 VDD1.n4 VDD1.t7 1.27136
R2587 VDD1.n4 VDD1.t1 1.27136
R2588 VDD1.n0 VDD1.t6 1.27136
R2589 VDD1.n0 VDD1.t0 1.27136
R2590 VDD1.n2 VDD1.t5 1.27136
R2591 VDD1.n2 VDD1.t3 1.27136
R2592 VDD1.n1 VDD1.t4 1.27136
R2593 VDD1.n1 VDD1.t2 1.27136
R2594 VDD1 VDD1.n5 0.459552
C0 VP VN 6.20469f
C1 VN VTAIL 7.52595f
C2 VP VTAIL 7.540061f
C3 VN VDD1 0.148557f
C4 VP VDD1 8.029181f
C5 VN VDD2 7.842721f
C6 VP VDD2 0.335538f
C7 VTAIL VDD1 12.431299f
C8 VTAIL VDD2 12.474099f
C9 VDD1 VDD2 0.908091f
C10 VDD2 B 3.921554f
C11 VDD1 B 4.172734f
C12 VTAIL B 11.116419f
C13 VN B 9.54934f
C14 VP B 7.535652f
C15 VDD1.t6 B 0.326298f
C16 VDD1.t0 B 0.326298f
C17 VDD1.n0 B 2.9624f
C18 VDD1.t4 B 0.326298f
C19 VDD1.t2 B 0.326298f
C20 VDD1.n1 B 2.96171f
C21 VDD1.t5 B 0.326298f
C22 VDD1.t3 B 0.326298f
C23 VDD1.n2 B 2.96171f
C24 VDD1.n3 B 2.68903f
C25 VDD1.t7 B 0.326298f
C26 VDD1.t1 B 0.326298f
C27 VDD1.n4 B 2.95922f
C28 VDD1.n5 B 2.80924f
C29 VP.n0 B 0.040446f
C30 VP.t2 B 1.50351f
C31 VP.n1 B 0.549155f
C32 VP.n2 B 0.040446f
C33 VP.t5 B 1.50351f
C34 VP.n3 B 0.017346f
C35 VP.n4 B 0.040446f
C36 VP.t6 B 1.55709f
C37 VP.t0 B 1.50351f
C38 VP.n5 B 0.549155f
C39 VP.n6 B 0.172625f
C40 VP.t7 B 1.50351f
C41 VP.t1 B 1.58368f
C42 VP.n7 B 0.591067f
C43 VP.n8 B 0.592405f
C44 VP.n9 B 0.047686f
C45 VP.n10 B 0.047686f
C46 VP.n11 B 0.040446f
C47 VP.n12 B 0.040446f
C48 VP.n13 B 0.051461f
C49 VP.n14 B 0.017346f
C50 VP.n15 B 0.591219f
C51 VP.n16 B 1.90421f
C52 VP.t3 B 1.55709f
C53 VP.n17 B 0.591219f
C54 VP.n18 B 1.93623f
C55 VP.n19 B 0.040446f
C56 VP.n20 B 0.040446f
C57 VP.n21 B 0.051461f
C58 VP.n22 B 0.549155f
C59 VP.n23 B 0.047686f
C60 VP.n24 B 0.047686f
C61 VP.n25 B 0.040446f
C62 VP.n26 B 0.040446f
C63 VP.n27 B 0.051461f
C64 VP.n28 B 0.017346f
C65 VP.t4 B 1.55709f
C66 VP.n29 B 0.591219f
C67 VP.n30 B 0.031344f
C68 VTAIL.t13 B 0.235348f
C69 VTAIL.t8 B 0.235348f
C70 VTAIL.n0 B 2.08274f
C71 VTAIL.n1 B 0.246593f
C72 VTAIL.n2 B 0.027643f
C73 VTAIL.n3 B 0.019116f
C74 VTAIL.n4 B 0.010272f
C75 VTAIL.n5 B 0.024279f
C76 VTAIL.n6 B 0.010574f
C77 VTAIL.n7 B 0.019116f
C78 VTAIL.n8 B 0.010876f
C79 VTAIL.n9 B 0.024279f
C80 VTAIL.n10 B 0.010876f
C81 VTAIL.n11 B 0.019116f
C82 VTAIL.n12 B 0.010272f
C83 VTAIL.n13 B 0.024279f
C84 VTAIL.n14 B 0.010876f
C85 VTAIL.n15 B 0.019116f
C86 VTAIL.n16 B 0.010272f
C87 VTAIL.n17 B 0.024279f
C88 VTAIL.n18 B 0.010876f
C89 VTAIL.n19 B 0.019116f
C90 VTAIL.n20 B 0.010272f
C91 VTAIL.n21 B 0.024279f
C92 VTAIL.n22 B 0.010876f
C93 VTAIL.n23 B 0.019116f
C94 VTAIL.n24 B 0.010272f
C95 VTAIL.n25 B 0.024279f
C96 VTAIL.n26 B 0.010876f
C97 VTAIL.n27 B 1.29451f
C98 VTAIL.n28 B 0.010272f
C99 VTAIL.t11 B 0.040071f
C100 VTAIL.n29 B 0.127456f
C101 VTAIL.n30 B 0.014342f
C102 VTAIL.n31 B 0.018209f
C103 VTAIL.n32 B 0.024279f
C104 VTAIL.n33 B 0.010876f
C105 VTAIL.n34 B 0.010272f
C106 VTAIL.n35 B 0.019116f
C107 VTAIL.n36 B 0.019116f
C108 VTAIL.n37 B 0.010272f
C109 VTAIL.n38 B 0.010876f
C110 VTAIL.n39 B 0.024279f
C111 VTAIL.n40 B 0.024279f
C112 VTAIL.n41 B 0.010876f
C113 VTAIL.n42 B 0.010272f
C114 VTAIL.n43 B 0.019116f
C115 VTAIL.n44 B 0.019116f
C116 VTAIL.n45 B 0.010272f
C117 VTAIL.n46 B 0.010876f
C118 VTAIL.n47 B 0.024279f
C119 VTAIL.n48 B 0.024279f
C120 VTAIL.n49 B 0.010876f
C121 VTAIL.n50 B 0.010272f
C122 VTAIL.n51 B 0.019116f
C123 VTAIL.n52 B 0.019116f
C124 VTAIL.n53 B 0.010272f
C125 VTAIL.n54 B 0.010876f
C126 VTAIL.n55 B 0.024279f
C127 VTAIL.n56 B 0.024279f
C128 VTAIL.n57 B 0.010876f
C129 VTAIL.n58 B 0.010272f
C130 VTAIL.n59 B 0.019116f
C131 VTAIL.n60 B 0.019116f
C132 VTAIL.n61 B 0.010272f
C133 VTAIL.n62 B 0.010876f
C134 VTAIL.n63 B 0.024279f
C135 VTAIL.n64 B 0.024279f
C136 VTAIL.n65 B 0.010876f
C137 VTAIL.n66 B 0.010272f
C138 VTAIL.n67 B 0.019116f
C139 VTAIL.n68 B 0.019116f
C140 VTAIL.n69 B 0.010272f
C141 VTAIL.n70 B 0.010272f
C142 VTAIL.n71 B 0.010876f
C143 VTAIL.n72 B 0.024279f
C144 VTAIL.n73 B 0.024279f
C145 VTAIL.n74 B 0.024279f
C146 VTAIL.n75 B 0.010574f
C147 VTAIL.n76 B 0.010272f
C148 VTAIL.n77 B 0.019116f
C149 VTAIL.n78 B 0.019116f
C150 VTAIL.n79 B 0.010272f
C151 VTAIL.n80 B 0.010876f
C152 VTAIL.n81 B 0.024279f
C153 VTAIL.n82 B 0.053929f
C154 VTAIL.n83 B 0.010876f
C155 VTAIL.n84 B 0.010272f
C156 VTAIL.n85 B 0.04993f
C157 VTAIL.n86 B 0.030483f
C158 VTAIL.n87 B 0.112236f
C159 VTAIL.n88 B 0.027643f
C160 VTAIL.n89 B 0.019116f
C161 VTAIL.n90 B 0.010272f
C162 VTAIL.n91 B 0.024279f
C163 VTAIL.n92 B 0.010574f
C164 VTAIL.n93 B 0.019116f
C165 VTAIL.n94 B 0.010876f
C166 VTAIL.n95 B 0.024279f
C167 VTAIL.n96 B 0.010876f
C168 VTAIL.n97 B 0.019116f
C169 VTAIL.n98 B 0.010272f
C170 VTAIL.n99 B 0.024279f
C171 VTAIL.n100 B 0.010876f
C172 VTAIL.n101 B 0.019116f
C173 VTAIL.n102 B 0.010272f
C174 VTAIL.n103 B 0.024279f
C175 VTAIL.n104 B 0.010876f
C176 VTAIL.n105 B 0.019116f
C177 VTAIL.n106 B 0.010272f
C178 VTAIL.n107 B 0.024279f
C179 VTAIL.n108 B 0.010876f
C180 VTAIL.n109 B 0.019116f
C181 VTAIL.n110 B 0.010272f
C182 VTAIL.n111 B 0.024279f
C183 VTAIL.n112 B 0.010876f
C184 VTAIL.n113 B 1.29451f
C185 VTAIL.n114 B 0.010272f
C186 VTAIL.t7 B 0.040071f
C187 VTAIL.n115 B 0.127456f
C188 VTAIL.n116 B 0.014342f
C189 VTAIL.n117 B 0.018209f
C190 VTAIL.n118 B 0.024279f
C191 VTAIL.n119 B 0.010876f
C192 VTAIL.n120 B 0.010272f
C193 VTAIL.n121 B 0.019116f
C194 VTAIL.n122 B 0.019116f
C195 VTAIL.n123 B 0.010272f
C196 VTAIL.n124 B 0.010876f
C197 VTAIL.n125 B 0.024279f
C198 VTAIL.n126 B 0.024279f
C199 VTAIL.n127 B 0.010876f
C200 VTAIL.n128 B 0.010272f
C201 VTAIL.n129 B 0.019116f
C202 VTAIL.n130 B 0.019116f
C203 VTAIL.n131 B 0.010272f
C204 VTAIL.n132 B 0.010876f
C205 VTAIL.n133 B 0.024279f
C206 VTAIL.n134 B 0.024279f
C207 VTAIL.n135 B 0.010876f
C208 VTAIL.n136 B 0.010272f
C209 VTAIL.n137 B 0.019116f
C210 VTAIL.n138 B 0.019116f
C211 VTAIL.n139 B 0.010272f
C212 VTAIL.n140 B 0.010876f
C213 VTAIL.n141 B 0.024279f
C214 VTAIL.n142 B 0.024279f
C215 VTAIL.n143 B 0.010876f
C216 VTAIL.n144 B 0.010272f
C217 VTAIL.n145 B 0.019116f
C218 VTAIL.n146 B 0.019116f
C219 VTAIL.n147 B 0.010272f
C220 VTAIL.n148 B 0.010876f
C221 VTAIL.n149 B 0.024279f
C222 VTAIL.n150 B 0.024279f
C223 VTAIL.n151 B 0.010876f
C224 VTAIL.n152 B 0.010272f
C225 VTAIL.n153 B 0.019116f
C226 VTAIL.n154 B 0.019116f
C227 VTAIL.n155 B 0.010272f
C228 VTAIL.n156 B 0.010272f
C229 VTAIL.n157 B 0.010876f
C230 VTAIL.n158 B 0.024279f
C231 VTAIL.n159 B 0.024279f
C232 VTAIL.n160 B 0.024279f
C233 VTAIL.n161 B 0.010574f
C234 VTAIL.n162 B 0.010272f
C235 VTAIL.n163 B 0.019116f
C236 VTAIL.n164 B 0.019116f
C237 VTAIL.n165 B 0.010272f
C238 VTAIL.n166 B 0.010876f
C239 VTAIL.n167 B 0.024279f
C240 VTAIL.n168 B 0.053929f
C241 VTAIL.n169 B 0.010876f
C242 VTAIL.n170 B 0.010272f
C243 VTAIL.n171 B 0.04993f
C244 VTAIL.n172 B 0.030483f
C245 VTAIL.n173 B 0.112236f
C246 VTAIL.t0 B 0.235348f
C247 VTAIL.t6 B 0.235348f
C248 VTAIL.n174 B 2.08274f
C249 VTAIL.n175 B 0.306728f
C250 VTAIL.n176 B 0.027643f
C251 VTAIL.n177 B 0.019116f
C252 VTAIL.n178 B 0.010272f
C253 VTAIL.n179 B 0.024279f
C254 VTAIL.n180 B 0.010574f
C255 VTAIL.n181 B 0.019116f
C256 VTAIL.n182 B 0.010876f
C257 VTAIL.n183 B 0.024279f
C258 VTAIL.n184 B 0.010876f
C259 VTAIL.n185 B 0.019116f
C260 VTAIL.n186 B 0.010272f
C261 VTAIL.n187 B 0.024279f
C262 VTAIL.n188 B 0.010876f
C263 VTAIL.n189 B 0.019116f
C264 VTAIL.n190 B 0.010272f
C265 VTAIL.n191 B 0.024279f
C266 VTAIL.n192 B 0.010876f
C267 VTAIL.n193 B 0.019116f
C268 VTAIL.n194 B 0.010272f
C269 VTAIL.n195 B 0.024279f
C270 VTAIL.n196 B 0.010876f
C271 VTAIL.n197 B 0.019116f
C272 VTAIL.n198 B 0.010272f
C273 VTAIL.n199 B 0.024279f
C274 VTAIL.n200 B 0.010876f
C275 VTAIL.n201 B 1.29451f
C276 VTAIL.n202 B 0.010272f
C277 VTAIL.t3 B 0.040071f
C278 VTAIL.n203 B 0.127456f
C279 VTAIL.n204 B 0.014342f
C280 VTAIL.n205 B 0.018209f
C281 VTAIL.n206 B 0.024279f
C282 VTAIL.n207 B 0.010876f
C283 VTAIL.n208 B 0.010272f
C284 VTAIL.n209 B 0.019116f
C285 VTAIL.n210 B 0.019116f
C286 VTAIL.n211 B 0.010272f
C287 VTAIL.n212 B 0.010876f
C288 VTAIL.n213 B 0.024279f
C289 VTAIL.n214 B 0.024279f
C290 VTAIL.n215 B 0.010876f
C291 VTAIL.n216 B 0.010272f
C292 VTAIL.n217 B 0.019116f
C293 VTAIL.n218 B 0.019116f
C294 VTAIL.n219 B 0.010272f
C295 VTAIL.n220 B 0.010876f
C296 VTAIL.n221 B 0.024279f
C297 VTAIL.n222 B 0.024279f
C298 VTAIL.n223 B 0.010876f
C299 VTAIL.n224 B 0.010272f
C300 VTAIL.n225 B 0.019116f
C301 VTAIL.n226 B 0.019116f
C302 VTAIL.n227 B 0.010272f
C303 VTAIL.n228 B 0.010876f
C304 VTAIL.n229 B 0.024279f
C305 VTAIL.n230 B 0.024279f
C306 VTAIL.n231 B 0.010876f
C307 VTAIL.n232 B 0.010272f
C308 VTAIL.n233 B 0.019116f
C309 VTAIL.n234 B 0.019116f
C310 VTAIL.n235 B 0.010272f
C311 VTAIL.n236 B 0.010876f
C312 VTAIL.n237 B 0.024279f
C313 VTAIL.n238 B 0.024279f
C314 VTAIL.n239 B 0.010876f
C315 VTAIL.n240 B 0.010272f
C316 VTAIL.n241 B 0.019116f
C317 VTAIL.n242 B 0.019116f
C318 VTAIL.n243 B 0.010272f
C319 VTAIL.n244 B 0.010272f
C320 VTAIL.n245 B 0.010876f
C321 VTAIL.n246 B 0.024279f
C322 VTAIL.n247 B 0.024279f
C323 VTAIL.n248 B 0.024279f
C324 VTAIL.n249 B 0.010574f
C325 VTAIL.n250 B 0.010272f
C326 VTAIL.n251 B 0.019116f
C327 VTAIL.n252 B 0.019116f
C328 VTAIL.n253 B 0.010272f
C329 VTAIL.n254 B 0.010876f
C330 VTAIL.n255 B 0.024279f
C331 VTAIL.n256 B 0.053929f
C332 VTAIL.n257 B 0.010876f
C333 VTAIL.n258 B 0.010272f
C334 VTAIL.n259 B 0.04993f
C335 VTAIL.n260 B 0.030483f
C336 VTAIL.n261 B 1.23397f
C337 VTAIL.n262 B 0.027643f
C338 VTAIL.n263 B 0.019116f
C339 VTAIL.n264 B 0.010272f
C340 VTAIL.n265 B 0.024279f
C341 VTAIL.n266 B 0.010574f
C342 VTAIL.n267 B 0.019116f
C343 VTAIL.n268 B 0.010574f
C344 VTAIL.n269 B 0.010272f
C345 VTAIL.n270 B 0.024279f
C346 VTAIL.n271 B 0.024279f
C347 VTAIL.n272 B 0.010876f
C348 VTAIL.n273 B 0.019116f
C349 VTAIL.n274 B 0.010272f
C350 VTAIL.n275 B 0.024279f
C351 VTAIL.n276 B 0.010876f
C352 VTAIL.n277 B 0.019116f
C353 VTAIL.n278 B 0.010272f
C354 VTAIL.n279 B 0.024279f
C355 VTAIL.n280 B 0.010876f
C356 VTAIL.n281 B 0.019116f
C357 VTAIL.n282 B 0.010272f
C358 VTAIL.n283 B 0.024279f
C359 VTAIL.n284 B 0.010876f
C360 VTAIL.n285 B 0.019116f
C361 VTAIL.n286 B 0.010272f
C362 VTAIL.n287 B 0.024279f
C363 VTAIL.n288 B 0.010876f
C364 VTAIL.n289 B 1.29451f
C365 VTAIL.n290 B 0.010272f
C366 VTAIL.t14 B 0.040071f
C367 VTAIL.n291 B 0.127456f
C368 VTAIL.n292 B 0.014342f
C369 VTAIL.n293 B 0.018209f
C370 VTAIL.n294 B 0.024279f
C371 VTAIL.n295 B 0.010876f
C372 VTAIL.n296 B 0.010272f
C373 VTAIL.n297 B 0.019116f
C374 VTAIL.n298 B 0.019116f
C375 VTAIL.n299 B 0.010272f
C376 VTAIL.n300 B 0.010876f
C377 VTAIL.n301 B 0.024279f
C378 VTAIL.n302 B 0.024279f
C379 VTAIL.n303 B 0.010876f
C380 VTAIL.n304 B 0.010272f
C381 VTAIL.n305 B 0.019116f
C382 VTAIL.n306 B 0.019116f
C383 VTAIL.n307 B 0.010272f
C384 VTAIL.n308 B 0.010876f
C385 VTAIL.n309 B 0.024279f
C386 VTAIL.n310 B 0.024279f
C387 VTAIL.n311 B 0.010876f
C388 VTAIL.n312 B 0.010272f
C389 VTAIL.n313 B 0.019116f
C390 VTAIL.n314 B 0.019116f
C391 VTAIL.n315 B 0.010272f
C392 VTAIL.n316 B 0.010876f
C393 VTAIL.n317 B 0.024279f
C394 VTAIL.n318 B 0.024279f
C395 VTAIL.n319 B 0.010876f
C396 VTAIL.n320 B 0.010272f
C397 VTAIL.n321 B 0.019116f
C398 VTAIL.n322 B 0.019116f
C399 VTAIL.n323 B 0.010272f
C400 VTAIL.n324 B 0.010876f
C401 VTAIL.n325 B 0.024279f
C402 VTAIL.n326 B 0.024279f
C403 VTAIL.n327 B 0.010876f
C404 VTAIL.n328 B 0.010272f
C405 VTAIL.n329 B 0.019116f
C406 VTAIL.n330 B 0.019116f
C407 VTAIL.n331 B 0.010272f
C408 VTAIL.n332 B 0.010876f
C409 VTAIL.n333 B 0.024279f
C410 VTAIL.n334 B 0.024279f
C411 VTAIL.n335 B 0.010876f
C412 VTAIL.n336 B 0.010272f
C413 VTAIL.n337 B 0.019116f
C414 VTAIL.n338 B 0.019116f
C415 VTAIL.n339 B 0.010272f
C416 VTAIL.n340 B 0.010876f
C417 VTAIL.n341 B 0.024279f
C418 VTAIL.n342 B 0.053929f
C419 VTAIL.n343 B 0.010876f
C420 VTAIL.n344 B 0.010272f
C421 VTAIL.n345 B 0.04993f
C422 VTAIL.n346 B 0.030483f
C423 VTAIL.n347 B 1.23397f
C424 VTAIL.t9 B 0.235348f
C425 VTAIL.t15 B 0.235348f
C426 VTAIL.n348 B 2.08275f
C427 VTAIL.n349 B 0.306719f
C428 VTAIL.n350 B 0.027643f
C429 VTAIL.n351 B 0.019116f
C430 VTAIL.n352 B 0.010272f
C431 VTAIL.n353 B 0.024279f
C432 VTAIL.n354 B 0.010574f
C433 VTAIL.n355 B 0.019116f
C434 VTAIL.n356 B 0.010574f
C435 VTAIL.n357 B 0.010272f
C436 VTAIL.n358 B 0.024279f
C437 VTAIL.n359 B 0.024279f
C438 VTAIL.n360 B 0.010876f
C439 VTAIL.n361 B 0.019116f
C440 VTAIL.n362 B 0.010272f
C441 VTAIL.n363 B 0.024279f
C442 VTAIL.n364 B 0.010876f
C443 VTAIL.n365 B 0.019116f
C444 VTAIL.n366 B 0.010272f
C445 VTAIL.n367 B 0.024279f
C446 VTAIL.n368 B 0.010876f
C447 VTAIL.n369 B 0.019116f
C448 VTAIL.n370 B 0.010272f
C449 VTAIL.n371 B 0.024279f
C450 VTAIL.n372 B 0.010876f
C451 VTAIL.n373 B 0.019116f
C452 VTAIL.n374 B 0.010272f
C453 VTAIL.n375 B 0.024279f
C454 VTAIL.n376 B 0.010876f
C455 VTAIL.n377 B 1.29451f
C456 VTAIL.n378 B 0.010272f
C457 VTAIL.t10 B 0.040071f
C458 VTAIL.n379 B 0.127456f
C459 VTAIL.n380 B 0.014342f
C460 VTAIL.n381 B 0.018209f
C461 VTAIL.n382 B 0.024279f
C462 VTAIL.n383 B 0.010876f
C463 VTAIL.n384 B 0.010272f
C464 VTAIL.n385 B 0.019116f
C465 VTAIL.n386 B 0.019116f
C466 VTAIL.n387 B 0.010272f
C467 VTAIL.n388 B 0.010876f
C468 VTAIL.n389 B 0.024279f
C469 VTAIL.n390 B 0.024279f
C470 VTAIL.n391 B 0.010876f
C471 VTAIL.n392 B 0.010272f
C472 VTAIL.n393 B 0.019116f
C473 VTAIL.n394 B 0.019116f
C474 VTAIL.n395 B 0.010272f
C475 VTAIL.n396 B 0.010876f
C476 VTAIL.n397 B 0.024279f
C477 VTAIL.n398 B 0.024279f
C478 VTAIL.n399 B 0.010876f
C479 VTAIL.n400 B 0.010272f
C480 VTAIL.n401 B 0.019116f
C481 VTAIL.n402 B 0.019116f
C482 VTAIL.n403 B 0.010272f
C483 VTAIL.n404 B 0.010876f
C484 VTAIL.n405 B 0.024279f
C485 VTAIL.n406 B 0.024279f
C486 VTAIL.n407 B 0.010876f
C487 VTAIL.n408 B 0.010272f
C488 VTAIL.n409 B 0.019116f
C489 VTAIL.n410 B 0.019116f
C490 VTAIL.n411 B 0.010272f
C491 VTAIL.n412 B 0.010876f
C492 VTAIL.n413 B 0.024279f
C493 VTAIL.n414 B 0.024279f
C494 VTAIL.n415 B 0.010876f
C495 VTAIL.n416 B 0.010272f
C496 VTAIL.n417 B 0.019116f
C497 VTAIL.n418 B 0.019116f
C498 VTAIL.n419 B 0.010272f
C499 VTAIL.n420 B 0.010876f
C500 VTAIL.n421 B 0.024279f
C501 VTAIL.n422 B 0.024279f
C502 VTAIL.n423 B 0.010876f
C503 VTAIL.n424 B 0.010272f
C504 VTAIL.n425 B 0.019116f
C505 VTAIL.n426 B 0.019116f
C506 VTAIL.n427 B 0.010272f
C507 VTAIL.n428 B 0.010876f
C508 VTAIL.n429 B 0.024279f
C509 VTAIL.n430 B 0.053929f
C510 VTAIL.n431 B 0.010876f
C511 VTAIL.n432 B 0.010272f
C512 VTAIL.n433 B 0.04993f
C513 VTAIL.n434 B 0.030483f
C514 VTAIL.n435 B 0.112236f
C515 VTAIL.n436 B 0.027643f
C516 VTAIL.n437 B 0.019116f
C517 VTAIL.n438 B 0.010272f
C518 VTAIL.n439 B 0.024279f
C519 VTAIL.n440 B 0.010574f
C520 VTAIL.n441 B 0.019116f
C521 VTAIL.n442 B 0.010574f
C522 VTAIL.n443 B 0.010272f
C523 VTAIL.n444 B 0.024279f
C524 VTAIL.n445 B 0.024279f
C525 VTAIL.n446 B 0.010876f
C526 VTAIL.n447 B 0.019116f
C527 VTAIL.n448 B 0.010272f
C528 VTAIL.n449 B 0.024279f
C529 VTAIL.n450 B 0.010876f
C530 VTAIL.n451 B 0.019116f
C531 VTAIL.n452 B 0.010272f
C532 VTAIL.n453 B 0.024279f
C533 VTAIL.n454 B 0.010876f
C534 VTAIL.n455 B 0.019116f
C535 VTAIL.n456 B 0.010272f
C536 VTAIL.n457 B 0.024279f
C537 VTAIL.n458 B 0.010876f
C538 VTAIL.n459 B 0.019116f
C539 VTAIL.n460 B 0.010272f
C540 VTAIL.n461 B 0.024279f
C541 VTAIL.n462 B 0.010876f
C542 VTAIL.n463 B 1.29451f
C543 VTAIL.n464 B 0.010272f
C544 VTAIL.t4 B 0.040071f
C545 VTAIL.n465 B 0.127456f
C546 VTAIL.n466 B 0.014342f
C547 VTAIL.n467 B 0.018209f
C548 VTAIL.n468 B 0.024279f
C549 VTAIL.n469 B 0.010876f
C550 VTAIL.n470 B 0.010272f
C551 VTAIL.n471 B 0.019116f
C552 VTAIL.n472 B 0.019116f
C553 VTAIL.n473 B 0.010272f
C554 VTAIL.n474 B 0.010876f
C555 VTAIL.n475 B 0.024279f
C556 VTAIL.n476 B 0.024279f
C557 VTAIL.n477 B 0.010876f
C558 VTAIL.n478 B 0.010272f
C559 VTAIL.n479 B 0.019116f
C560 VTAIL.n480 B 0.019116f
C561 VTAIL.n481 B 0.010272f
C562 VTAIL.n482 B 0.010876f
C563 VTAIL.n483 B 0.024279f
C564 VTAIL.n484 B 0.024279f
C565 VTAIL.n485 B 0.010876f
C566 VTAIL.n486 B 0.010272f
C567 VTAIL.n487 B 0.019116f
C568 VTAIL.n488 B 0.019116f
C569 VTAIL.n489 B 0.010272f
C570 VTAIL.n490 B 0.010876f
C571 VTAIL.n491 B 0.024279f
C572 VTAIL.n492 B 0.024279f
C573 VTAIL.n493 B 0.010876f
C574 VTAIL.n494 B 0.010272f
C575 VTAIL.n495 B 0.019116f
C576 VTAIL.n496 B 0.019116f
C577 VTAIL.n497 B 0.010272f
C578 VTAIL.n498 B 0.010876f
C579 VTAIL.n499 B 0.024279f
C580 VTAIL.n500 B 0.024279f
C581 VTAIL.n501 B 0.010876f
C582 VTAIL.n502 B 0.010272f
C583 VTAIL.n503 B 0.019116f
C584 VTAIL.n504 B 0.019116f
C585 VTAIL.n505 B 0.010272f
C586 VTAIL.n506 B 0.010876f
C587 VTAIL.n507 B 0.024279f
C588 VTAIL.n508 B 0.024279f
C589 VTAIL.n509 B 0.010876f
C590 VTAIL.n510 B 0.010272f
C591 VTAIL.n511 B 0.019116f
C592 VTAIL.n512 B 0.019116f
C593 VTAIL.n513 B 0.010272f
C594 VTAIL.n514 B 0.010876f
C595 VTAIL.n515 B 0.024279f
C596 VTAIL.n516 B 0.053929f
C597 VTAIL.n517 B 0.010876f
C598 VTAIL.n518 B 0.010272f
C599 VTAIL.n519 B 0.04993f
C600 VTAIL.n520 B 0.030483f
C601 VTAIL.n521 B 0.112236f
C602 VTAIL.t2 B 0.235348f
C603 VTAIL.t5 B 0.235348f
C604 VTAIL.n522 B 2.08275f
C605 VTAIL.n523 B 0.306719f
C606 VTAIL.n524 B 0.027643f
C607 VTAIL.n525 B 0.019116f
C608 VTAIL.n526 B 0.010272f
C609 VTAIL.n527 B 0.024279f
C610 VTAIL.n528 B 0.010574f
C611 VTAIL.n529 B 0.019116f
C612 VTAIL.n530 B 0.010574f
C613 VTAIL.n531 B 0.010272f
C614 VTAIL.n532 B 0.024279f
C615 VTAIL.n533 B 0.024279f
C616 VTAIL.n534 B 0.010876f
C617 VTAIL.n535 B 0.019116f
C618 VTAIL.n536 B 0.010272f
C619 VTAIL.n537 B 0.024279f
C620 VTAIL.n538 B 0.010876f
C621 VTAIL.n539 B 0.019116f
C622 VTAIL.n540 B 0.010272f
C623 VTAIL.n541 B 0.024279f
C624 VTAIL.n542 B 0.010876f
C625 VTAIL.n543 B 0.019116f
C626 VTAIL.n544 B 0.010272f
C627 VTAIL.n545 B 0.024279f
C628 VTAIL.n546 B 0.010876f
C629 VTAIL.n547 B 0.019116f
C630 VTAIL.n548 B 0.010272f
C631 VTAIL.n549 B 0.024279f
C632 VTAIL.n550 B 0.010876f
C633 VTAIL.n551 B 1.29451f
C634 VTAIL.n552 B 0.010272f
C635 VTAIL.t1 B 0.040071f
C636 VTAIL.n553 B 0.127456f
C637 VTAIL.n554 B 0.014342f
C638 VTAIL.n555 B 0.018209f
C639 VTAIL.n556 B 0.024279f
C640 VTAIL.n557 B 0.010876f
C641 VTAIL.n558 B 0.010272f
C642 VTAIL.n559 B 0.019116f
C643 VTAIL.n560 B 0.019116f
C644 VTAIL.n561 B 0.010272f
C645 VTAIL.n562 B 0.010876f
C646 VTAIL.n563 B 0.024279f
C647 VTAIL.n564 B 0.024279f
C648 VTAIL.n565 B 0.010876f
C649 VTAIL.n566 B 0.010272f
C650 VTAIL.n567 B 0.019116f
C651 VTAIL.n568 B 0.019116f
C652 VTAIL.n569 B 0.010272f
C653 VTAIL.n570 B 0.010876f
C654 VTAIL.n571 B 0.024279f
C655 VTAIL.n572 B 0.024279f
C656 VTAIL.n573 B 0.010876f
C657 VTAIL.n574 B 0.010272f
C658 VTAIL.n575 B 0.019116f
C659 VTAIL.n576 B 0.019116f
C660 VTAIL.n577 B 0.010272f
C661 VTAIL.n578 B 0.010876f
C662 VTAIL.n579 B 0.024279f
C663 VTAIL.n580 B 0.024279f
C664 VTAIL.n581 B 0.010876f
C665 VTAIL.n582 B 0.010272f
C666 VTAIL.n583 B 0.019116f
C667 VTAIL.n584 B 0.019116f
C668 VTAIL.n585 B 0.010272f
C669 VTAIL.n586 B 0.010876f
C670 VTAIL.n587 B 0.024279f
C671 VTAIL.n588 B 0.024279f
C672 VTAIL.n589 B 0.010876f
C673 VTAIL.n590 B 0.010272f
C674 VTAIL.n591 B 0.019116f
C675 VTAIL.n592 B 0.019116f
C676 VTAIL.n593 B 0.010272f
C677 VTAIL.n594 B 0.010876f
C678 VTAIL.n595 B 0.024279f
C679 VTAIL.n596 B 0.024279f
C680 VTAIL.n597 B 0.010876f
C681 VTAIL.n598 B 0.010272f
C682 VTAIL.n599 B 0.019116f
C683 VTAIL.n600 B 0.019116f
C684 VTAIL.n601 B 0.010272f
C685 VTAIL.n602 B 0.010876f
C686 VTAIL.n603 B 0.024279f
C687 VTAIL.n604 B 0.053929f
C688 VTAIL.n605 B 0.010876f
C689 VTAIL.n606 B 0.010272f
C690 VTAIL.n607 B 0.04993f
C691 VTAIL.n608 B 0.030483f
C692 VTAIL.n609 B 1.23397f
C693 VTAIL.n610 B 0.027643f
C694 VTAIL.n611 B 0.019116f
C695 VTAIL.n612 B 0.010272f
C696 VTAIL.n613 B 0.024279f
C697 VTAIL.n614 B 0.010574f
C698 VTAIL.n615 B 0.019116f
C699 VTAIL.n616 B 0.010876f
C700 VTAIL.n617 B 0.024279f
C701 VTAIL.n618 B 0.010876f
C702 VTAIL.n619 B 0.019116f
C703 VTAIL.n620 B 0.010272f
C704 VTAIL.n621 B 0.024279f
C705 VTAIL.n622 B 0.010876f
C706 VTAIL.n623 B 0.019116f
C707 VTAIL.n624 B 0.010272f
C708 VTAIL.n625 B 0.024279f
C709 VTAIL.n626 B 0.010876f
C710 VTAIL.n627 B 0.019116f
C711 VTAIL.n628 B 0.010272f
C712 VTAIL.n629 B 0.024279f
C713 VTAIL.n630 B 0.010876f
C714 VTAIL.n631 B 0.019116f
C715 VTAIL.n632 B 0.010272f
C716 VTAIL.n633 B 0.024279f
C717 VTAIL.n634 B 0.010876f
C718 VTAIL.n635 B 1.29451f
C719 VTAIL.n636 B 0.010272f
C720 VTAIL.t12 B 0.040071f
C721 VTAIL.n637 B 0.127456f
C722 VTAIL.n638 B 0.014342f
C723 VTAIL.n639 B 0.018209f
C724 VTAIL.n640 B 0.024279f
C725 VTAIL.n641 B 0.010876f
C726 VTAIL.n642 B 0.010272f
C727 VTAIL.n643 B 0.019116f
C728 VTAIL.n644 B 0.019116f
C729 VTAIL.n645 B 0.010272f
C730 VTAIL.n646 B 0.010876f
C731 VTAIL.n647 B 0.024279f
C732 VTAIL.n648 B 0.024279f
C733 VTAIL.n649 B 0.010876f
C734 VTAIL.n650 B 0.010272f
C735 VTAIL.n651 B 0.019116f
C736 VTAIL.n652 B 0.019116f
C737 VTAIL.n653 B 0.010272f
C738 VTAIL.n654 B 0.010876f
C739 VTAIL.n655 B 0.024279f
C740 VTAIL.n656 B 0.024279f
C741 VTAIL.n657 B 0.010876f
C742 VTAIL.n658 B 0.010272f
C743 VTAIL.n659 B 0.019116f
C744 VTAIL.n660 B 0.019116f
C745 VTAIL.n661 B 0.010272f
C746 VTAIL.n662 B 0.010876f
C747 VTAIL.n663 B 0.024279f
C748 VTAIL.n664 B 0.024279f
C749 VTAIL.n665 B 0.010876f
C750 VTAIL.n666 B 0.010272f
C751 VTAIL.n667 B 0.019116f
C752 VTAIL.n668 B 0.019116f
C753 VTAIL.n669 B 0.010272f
C754 VTAIL.n670 B 0.010876f
C755 VTAIL.n671 B 0.024279f
C756 VTAIL.n672 B 0.024279f
C757 VTAIL.n673 B 0.010876f
C758 VTAIL.n674 B 0.010272f
C759 VTAIL.n675 B 0.019116f
C760 VTAIL.n676 B 0.019116f
C761 VTAIL.n677 B 0.010272f
C762 VTAIL.n678 B 0.010272f
C763 VTAIL.n679 B 0.010876f
C764 VTAIL.n680 B 0.024279f
C765 VTAIL.n681 B 0.024279f
C766 VTAIL.n682 B 0.024279f
C767 VTAIL.n683 B 0.010574f
C768 VTAIL.n684 B 0.010272f
C769 VTAIL.n685 B 0.019116f
C770 VTAIL.n686 B 0.019116f
C771 VTAIL.n687 B 0.010272f
C772 VTAIL.n688 B 0.010876f
C773 VTAIL.n689 B 0.024279f
C774 VTAIL.n690 B 0.053929f
C775 VTAIL.n691 B 0.010876f
C776 VTAIL.n692 B 0.010272f
C777 VTAIL.n693 B 0.04993f
C778 VTAIL.n694 B 0.030483f
C779 VTAIL.n695 B 1.23038f
C780 VDD2.t3 B 0.326264f
C781 VDD2.t1 B 0.326264f
C782 VDD2.n0 B 2.9614f
C783 VDD2.t4 B 0.326264f
C784 VDD2.t0 B 0.326264f
C785 VDD2.n1 B 2.9614f
C786 VDD2.n2 B 2.63256f
C787 VDD2.t6 B 0.326264f
C788 VDD2.t5 B 0.326264f
C789 VDD2.n3 B 2.95892f
C790 VDD2.n4 B 2.77719f
C791 VDD2.t7 B 0.326264f
C792 VDD2.t2 B 0.326264f
C793 VDD2.n5 B 2.96137f
C794 VN.n0 B 0.039968f
C795 VN.t7 B 1.48576f
C796 VN.n1 B 0.542672f
C797 VN.n2 B 0.170587f
C798 VN.t2 B 1.48576f
C799 VN.t4 B 1.56498f
C800 VN.n3 B 0.584089f
C801 VN.n4 B 0.585412f
C802 VN.n5 B 0.047123f
C803 VN.n6 B 0.047123f
C804 VN.n7 B 0.039968f
C805 VN.n8 B 0.039968f
C806 VN.n9 B 0.050853f
C807 VN.n10 B 0.017141f
C808 VN.t3 B 1.53871f
C809 VN.n11 B 0.584239f
C810 VN.n12 B 0.030974f
C811 VN.n13 B 0.039968f
C812 VN.t6 B 1.48576f
C813 VN.n14 B 0.542672f
C814 VN.n15 B 0.170587f
C815 VN.t0 B 1.48576f
C816 VN.t5 B 1.56498f
C817 VN.n16 B 0.584089f
C818 VN.n17 B 0.585412f
C819 VN.n18 B 0.047123f
C820 VN.n19 B 0.047123f
C821 VN.n20 B 0.039968f
C822 VN.n21 B 0.039968f
C823 VN.n22 B 0.050853f
C824 VN.n23 B 0.017141f
C825 VN.t1 B 1.53871f
C826 VN.n24 B 0.584239f
C827 VN.n25 B 1.90785f
.ends

