* NGSPICE file created from diff_pair_sample_1064.ext - technology: sky130A

.subckt diff_pair_sample_1064 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t16 VP.t0 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.5511 pd=3.67 as=0.5511 ps=3.67 w=3.34 l=0.3
X1 VDD2.t9 VN.t0 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.5511 pd=3.67 as=0.5511 ps=3.67 w=3.34 l=0.3
X2 VTAIL.t2 VN.t1 VDD2.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5511 pd=3.67 as=0.5511 ps=3.67 w=3.34 l=0.3
X3 VTAIL.t3 VN.t2 VDD2.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.5511 pd=3.67 as=0.5511 ps=3.67 w=3.34 l=0.3
X4 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=1.3026 pd=7.46 as=0 ps=0 w=3.34 l=0.3
X5 VDD1.t9 VP.t1 VTAIL.t15 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3026 pd=7.46 as=0.5511 ps=3.67 w=3.34 l=0.3
X6 VDD1.t1 VP.t2 VTAIL.t14 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5511 pd=3.67 as=1.3026 ps=7.46 w=3.34 l=0.3
X7 VDD1.t5 VP.t3 VTAIL.t13 B.t6 sky130_fd_pr__nfet_01v8 ad=0.5511 pd=3.67 as=0.5511 ps=3.67 w=3.34 l=0.3
X8 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=1.3026 pd=7.46 as=0 ps=0 w=3.34 l=0.3
X9 VDD1.t3 VP.t4 VTAIL.t12 B.t9 sky130_fd_pr__nfet_01v8 ad=0.5511 pd=3.67 as=1.3026 ps=7.46 w=3.34 l=0.3
X10 VDD2.t6 VN.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.5511 pd=3.67 as=0.5511 ps=3.67 w=3.34 l=0.3
X11 VDD2.t5 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3026 pd=7.46 as=0.5511 ps=3.67 w=3.34 l=0.3
X12 VTAIL.t11 VP.t5 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.5511 pd=3.67 as=0.5511 ps=3.67 w=3.34 l=0.3
X13 VTAIL.t1 VN.t5 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.5511 pd=3.67 as=0.5511 ps=3.67 w=3.34 l=0.3
X14 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=1.3026 pd=7.46 as=0 ps=0 w=3.34 l=0.3
X15 VDD2.t3 VN.t6 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5511 pd=3.67 as=1.3026 ps=7.46 w=3.34 l=0.3
X16 VDD1.t8 VP.t6 VTAIL.t10 B.t8 sky130_fd_pr__nfet_01v8 ad=1.3026 pd=7.46 as=0.5511 ps=3.67 w=3.34 l=0.3
X17 VDD1.t6 VP.t7 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=0.5511 pd=3.67 as=0.5511 ps=3.67 w=3.34 l=0.3
X18 VDD2.t2 VN.t7 VTAIL.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=0.5511 pd=3.67 as=1.3026 ps=7.46 w=3.34 l=0.3
X19 VDD2.t1 VN.t8 VTAIL.t18 B.t8 sky130_fd_pr__nfet_01v8 ad=1.3026 pd=7.46 as=0.5511 ps=3.67 w=3.34 l=0.3
X20 VTAIL.t19 VN.t9 VDD2.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=0.5511 pd=3.67 as=0.5511 ps=3.67 w=3.34 l=0.3
X21 VTAIL.t8 VP.t8 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=0.5511 pd=3.67 as=0.5511 ps=3.67 w=3.34 l=0.3
X22 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.3026 pd=7.46 as=0 ps=0 w=3.34 l=0.3
X23 VTAIL.t7 VP.t9 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5511 pd=3.67 as=0.5511 ps=3.67 w=3.34 l=0.3
R0 VP.n21 VP.t2 410.723
R1 VP.n14 VP.t6 410.723
R2 VP.n5 VP.t1 410.723
R3 VP.n11 VP.t4 410.723
R4 VP.n18 VP.t3 372.748
R5 VP.n20 VP.t8 372.748
R6 VP.n13 VP.t0 372.748
R7 VP.n8 VP.t7 372.748
R8 VP.n4 VP.t5 372.748
R9 VP.n10 VP.t9 372.748
R10 VP.n6 VP.n5 161.489
R11 VP.n22 VP.n21 161.3
R12 VP.n6 VP.n3 161.3
R13 VP.n8 VP.n7 161.3
R14 VP.n9 VP.n2 161.3
R15 VP.n12 VP.n11 161.3
R16 VP.n19 VP.n0 161.3
R17 VP.n18 VP.n17 161.3
R18 VP.n16 VP.n1 161.3
R19 VP.n15 VP.n14 161.3
R20 VP.n18 VP.n1 73.0308
R21 VP.n19 VP.n18 73.0308
R22 VP.n8 VP.n3 73.0308
R23 VP.n9 VP.n8 73.0308
R24 VP.n14 VP.n13 54.0429
R25 VP.n21 VP.n20 54.0429
R26 VP.n5 VP.n4 54.0429
R27 VP.n11 VP.n10 54.0429
R28 VP.n15 VP.n12 34.1028
R29 VP.n13 VP.n1 18.9884
R30 VP.n20 VP.n19 18.9884
R31 VP.n4 VP.n3 18.9884
R32 VP.n10 VP.n9 18.9884
R33 VP.n7 VP.n6 0.189894
R34 VP.n7 VP.n2 0.189894
R35 VP.n12 VP.n2 0.189894
R36 VP.n16 VP.n15 0.189894
R37 VP.n17 VP.n16 0.189894
R38 VP.n17 VP.n0 0.189894
R39 VP.n22 VP.n0 0.189894
R40 VP VP.n22 0.0516364
R41 VDD1.n10 VDD1.n0 289.615
R42 VDD1.n27 VDD1.n17 289.615
R43 VDD1.n11 VDD1.n10 185
R44 VDD1.n9 VDD1.n8 185
R45 VDD1.n4 VDD1.n3 185
R46 VDD1.n21 VDD1.n20 185
R47 VDD1.n26 VDD1.n25 185
R48 VDD1.n28 VDD1.n27 185
R49 VDD1.n5 VDD1.t9 148.606
R50 VDD1.n22 VDD1.t8 148.606
R51 VDD1.n10 VDD1.n9 104.615
R52 VDD1.n9 VDD1.n3 104.615
R53 VDD1.n26 VDD1.n20 104.615
R54 VDD1.n27 VDD1.n26 104.615
R55 VDD1.n35 VDD1.n34 82.3677
R56 VDD1.n16 VDD1.n15 82.0159
R57 VDD1.n37 VDD1.n36 82.0157
R58 VDD1.n33 VDD1.n32 82.0157
R59 VDD1.n16 VDD1.n14 53.6739
R60 VDD1.n33 VDD1.n31 53.6739
R61 VDD1.t9 VDD1.n3 52.3082
R62 VDD1.t8 VDD1.n20 52.3082
R63 VDD1.n37 VDD1.n35 30.0289
R64 VDD1.n5 VDD1.n4 15.5966
R65 VDD1.n22 VDD1.n21 15.5966
R66 VDD1.n8 VDD1.n7 12.8005
R67 VDD1.n25 VDD1.n24 12.8005
R68 VDD1.n11 VDD1.n2 12.0247
R69 VDD1.n28 VDD1.n19 12.0247
R70 VDD1.n12 VDD1.n0 11.249
R71 VDD1.n29 VDD1.n17 11.249
R72 VDD1.n14 VDD1.n13 9.45567
R73 VDD1.n31 VDD1.n30 9.45567
R74 VDD1.n13 VDD1.n12 9.3005
R75 VDD1.n2 VDD1.n1 9.3005
R76 VDD1.n7 VDD1.n6 9.3005
R77 VDD1.n30 VDD1.n29 9.3005
R78 VDD1.n19 VDD1.n18 9.3005
R79 VDD1.n24 VDD1.n23 9.3005
R80 VDD1.n36 VDD1.t2 5.92864
R81 VDD1.n36 VDD1.t3 5.92864
R82 VDD1.n15 VDD1.t7 5.92864
R83 VDD1.n15 VDD1.t6 5.92864
R84 VDD1.n34 VDD1.t4 5.92864
R85 VDD1.n34 VDD1.t1 5.92864
R86 VDD1.n32 VDD1.t0 5.92864
R87 VDD1.n32 VDD1.t5 5.92864
R88 VDD1.n6 VDD1.n5 4.46457
R89 VDD1.n23 VDD1.n22 4.46457
R90 VDD1.n14 VDD1.n0 2.71565
R91 VDD1.n31 VDD1.n17 2.71565
R92 VDD1.n12 VDD1.n11 1.93989
R93 VDD1.n29 VDD1.n28 1.93989
R94 VDD1.n8 VDD1.n2 1.16414
R95 VDD1.n25 VDD1.n19 1.16414
R96 VDD1.n7 VDD1.n4 0.388379
R97 VDD1.n24 VDD1.n21 0.388379
R98 VDD1 VDD1.n37 0.349638
R99 VDD1 VDD1.n16 0.194466
R100 VDD1.n13 VDD1.n1 0.155672
R101 VDD1.n6 VDD1.n1 0.155672
R102 VDD1.n23 VDD1.n18 0.155672
R103 VDD1.n30 VDD1.n18 0.155672
R104 VDD1.n35 VDD1.n33 0.0809298
R105 VTAIL.n72 VTAIL.n62 289.615
R106 VTAIL.n12 VTAIL.n2 289.615
R107 VTAIL.n56 VTAIL.n46 289.615
R108 VTAIL.n36 VTAIL.n26 289.615
R109 VTAIL.n66 VTAIL.n65 185
R110 VTAIL.n71 VTAIL.n70 185
R111 VTAIL.n73 VTAIL.n72 185
R112 VTAIL.n6 VTAIL.n5 185
R113 VTAIL.n11 VTAIL.n10 185
R114 VTAIL.n13 VTAIL.n12 185
R115 VTAIL.n57 VTAIL.n56 185
R116 VTAIL.n55 VTAIL.n54 185
R117 VTAIL.n50 VTAIL.n49 185
R118 VTAIL.n37 VTAIL.n36 185
R119 VTAIL.n35 VTAIL.n34 185
R120 VTAIL.n30 VTAIL.n29 185
R121 VTAIL.n67 VTAIL.t17 148.606
R122 VTAIL.n7 VTAIL.t14 148.606
R123 VTAIL.n51 VTAIL.t12 148.606
R124 VTAIL.n31 VTAIL.t5 148.606
R125 VTAIL.n71 VTAIL.n65 104.615
R126 VTAIL.n72 VTAIL.n71 104.615
R127 VTAIL.n11 VTAIL.n5 104.615
R128 VTAIL.n12 VTAIL.n11 104.615
R129 VTAIL.n56 VTAIL.n55 104.615
R130 VTAIL.n55 VTAIL.n49 104.615
R131 VTAIL.n36 VTAIL.n35 104.615
R132 VTAIL.n35 VTAIL.n29 104.615
R133 VTAIL.n45 VTAIL.n44 65.3371
R134 VTAIL.n43 VTAIL.n42 65.3371
R135 VTAIL.n25 VTAIL.n24 65.3371
R136 VTAIL.n23 VTAIL.n22 65.3371
R137 VTAIL.n79 VTAIL.n78 65.337
R138 VTAIL.n1 VTAIL.n0 65.337
R139 VTAIL.n19 VTAIL.n18 65.337
R140 VTAIL.n21 VTAIL.n20 65.337
R141 VTAIL.t17 VTAIL.n65 52.3082
R142 VTAIL.t14 VTAIL.n5 52.3082
R143 VTAIL.t12 VTAIL.n49 52.3082
R144 VTAIL.t5 VTAIL.n29 52.3082
R145 VTAIL.n77 VTAIL.n76 36.452
R146 VTAIL.n17 VTAIL.n16 36.452
R147 VTAIL.n61 VTAIL.n60 36.452
R148 VTAIL.n41 VTAIL.n40 36.452
R149 VTAIL.n23 VTAIL.n21 16.3324
R150 VTAIL.n77 VTAIL.n61 15.7893
R151 VTAIL.n67 VTAIL.n66 15.5966
R152 VTAIL.n7 VTAIL.n6 15.5966
R153 VTAIL.n51 VTAIL.n50 15.5966
R154 VTAIL.n31 VTAIL.n30 15.5966
R155 VTAIL.n70 VTAIL.n69 12.8005
R156 VTAIL.n10 VTAIL.n9 12.8005
R157 VTAIL.n54 VTAIL.n53 12.8005
R158 VTAIL.n34 VTAIL.n33 12.8005
R159 VTAIL.n73 VTAIL.n64 12.0247
R160 VTAIL.n13 VTAIL.n4 12.0247
R161 VTAIL.n57 VTAIL.n48 12.0247
R162 VTAIL.n37 VTAIL.n28 12.0247
R163 VTAIL.n74 VTAIL.n62 11.249
R164 VTAIL.n14 VTAIL.n2 11.249
R165 VTAIL.n58 VTAIL.n46 11.249
R166 VTAIL.n38 VTAIL.n26 11.249
R167 VTAIL.n76 VTAIL.n75 9.45567
R168 VTAIL.n16 VTAIL.n15 9.45567
R169 VTAIL.n60 VTAIL.n59 9.45567
R170 VTAIL.n40 VTAIL.n39 9.45567
R171 VTAIL.n75 VTAIL.n74 9.3005
R172 VTAIL.n64 VTAIL.n63 9.3005
R173 VTAIL.n69 VTAIL.n68 9.3005
R174 VTAIL.n15 VTAIL.n14 9.3005
R175 VTAIL.n4 VTAIL.n3 9.3005
R176 VTAIL.n9 VTAIL.n8 9.3005
R177 VTAIL.n59 VTAIL.n58 9.3005
R178 VTAIL.n48 VTAIL.n47 9.3005
R179 VTAIL.n53 VTAIL.n52 9.3005
R180 VTAIL.n39 VTAIL.n38 9.3005
R181 VTAIL.n28 VTAIL.n27 9.3005
R182 VTAIL.n33 VTAIL.n32 9.3005
R183 VTAIL.n78 VTAIL.t4 5.92864
R184 VTAIL.n78 VTAIL.t2 5.92864
R185 VTAIL.n0 VTAIL.t0 5.92864
R186 VTAIL.n0 VTAIL.t3 5.92864
R187 VTAIL.n18 VTAIL.t13 5.92864
R188 VTAIL.n18 VTAIL.t8 5.92864
R189 VTAIL.n20 VTAIL.t10 5.92864
R190 VTAIL.n20 VTAIL.t16 5.92864
R191 VTAIL.n44 VTAIL.t9 5.92864
R192 VTAIL.n44 VTAIL.t7 5.92864
R193 VTAIL.n42 VTAIL.t15 5.92864
R194 VTAIL.n42 VTAIL.t11 5.92864
R195 VTAIL.n24 VTAIL.t6 5.92864
R196 VTAIL.n24 VTAIL.t19 5.92864
R197 VTAIL.n22 VTAIL.t18 5.92864
R198 VTAIL.n22 VTAIL.t1 5.92864
R199 VTAIL.n68 VTAIL.n67 4.46457
R200 VTAIL.n8 VTAIL.n7 4.46457
R201 VTAIL.n52 VTAIL.n51 4.46457
R202 VTAIL.n32 VTAIL.n31 4.46457
R203 VTAIL.n76 VTAIL.n62 2.71565
R204 VTAIL.n16 VTAIL.n2 2.71565
R205 VTAIL.n60 VTAIL.n46 2.71565
R206 VTAIL.n40 VTAIL.n26 2.71565
R207 VTAIL.n74 VTAIL.n73 1.93989
R208 VTAIL.n14 VTAIL.n13 1.93989
R209 VTAIL.n58 VTAIL.n57 1.93989
R210 VTAIL.n38 VTAIL.n37 1.93989
R211 VTAIL.n70 VTAIL.n64 1.16414
R212 VTAIL.n10 VTAIL.n4 1.16414
R213 VTAIL.n54 VTAIL.n48 1.16414
R214 VTAIL.n34 VTAIL.n28 1.16414
R215 VTAIL.n43 VTAIL.n41 0.741879
R216 VTAIL.n17 VTAIL.n1 0.741879
R217 VTAIL.n25 VTAIL.n23 0.543603
R218 VTAIL.n41 VTAIL.n25 0.543603
R219 VTAIL.n45 VTAIL.n43 0.543603
R220 VTAIL.n61 VTAIL.n45 0.543603
R221 VTAIL.n21 VTAIL.n19 0.543603
R222 VTAIL.n19 VTAIL.n17 0.543603
R223 VTAIL.n79 VTAIL.n77 0.543603
R224 VTAIL VTAIL.n1 0.466017
R225 VTAIL.n69 VTAIL.n66 0.388379
R226 VTAIL.n9 VTAIL.n6 0.388379
R227 VTAIL.n53 VTAIL.n50 0.388379
R228 VTAIL.n33 VTAIL.n30 0.388379
R229 VTAIL.n68 VTAIL.n63 0.155672
R230 VTAIL.n75 VTAIL.n63 0.155672
R231 VTAIL.n8 VTAIL.n3 0.155672
R232 VTAIL.n15 VTAIL.n3 0.155672
R233 VTAIL.n59 VTAIL.n47 0.155672
R234 VTAIL.n52 VTAIL.n47 0.155672
R235 VTAIL.n39 VTAIL.n27 0.155672
R236 VTAIL.n32 VTAIL.n27 0.155672
R237 VTAIL VTAIL.n79 0.0780862
R238 B.n370 B.n369 585
R239 B.n142 B.n58 585
R240 B.n141 B.n140 585
R241 B.n139 B.n138 585
R242 B.n137 B.n136 585
R243 B.n135 B.n134 585
R244 B.n133 B.n132 585
R245 B.n131 B.n130 585
R246 B.n129 B.n128 585
R247 B.n127 B.n126 585
R248 B.n125 B.n124 585
R249 B.n123 B.n122 585
R250 B.n121 B.n120 585
R251 B.n119 B.n118 585
R252 B.n117 B.n116 585
R253 B.n115 B.n114 585
R254 B.n113 B.n112 585
R255 B.n111 B.n110 585
R256 B.n109 B.n108 585
R257 B.n107 B.n106 585
R258 B.n105 B.n104 585
R259 B.n103 B.n102 585
R260 B.n101 B.n100 585
R261 B.n99 B.n98 585
R262 B.n97 B.n96 585
R263 B.n95 B.n94 585
R264 B.n93 B.n92 585
R265 B.n91 B.n90 585
R266 B.n89 B.n88 585
R267 B.n87 B.n86 585
R268 B.n85 B.n84 585
R269 B.n83 B.n82 585
R270 B.n81 B.n80 585
R271 B.n79 B.n78 585
R272 B.n77 B.n76 585
R273 B.n75 B.n74 585
R274 B.n73 B.n72 585
R275 B.n71 B.n70 585
R276 B.n69 B.n68 585
R277 B.n67 B.n66 585
R278 B.n38 B.n37 585
R279 B.n375 B.n374 585
R280 B.n368 B.n59 585
R281 B.n59 B.n35 585
R282 B.n367 B.n34 585
R283 B.n379 B.n34 585
R284 B.n366 B.n33 585
R285 B.n380 B.n33 585
R286 B.n365 B.n32 585
R287 B.n381 B.n32 585
R288 B.n364 B.n363 585
R289 B.n363 B.t18 585
R290 B.n362 B.n28 585
R291 B.n387 B.n28 585
R292 B.n361 B.n27 585
R293 B.n388 B.n27 585
R294 B.n360 B.n26 585
R295 B.n389 B.n26 585
R296 B.n359 B.n358 585
R297 B.n358 B.n22 585
R298 B.n357 B.n21 585
R299 B.n395 B.n21 585
R300 B.n356 B.n20 585
R301 B.n396 B.n20 585
R302 B.n355 B.n19 585
R303 B.n397 B.n19 585
R304 B.n354 B.n353 585
R305 B.n353 B.n18 585
R306 B.n352 B.n14 585
R307 B.n403 B.n14 585
R308 B.n351 B.n13 585
R309 B.n404 B.n13 585
R310 B.n350 B.n12 585
R311 B.n405 B.n12 585
R312 B.n349 B.n348 585
R313 B.n348 B.n11 585
R314 B.n347 B.n7 585
R315 B.n411 B.n7 585
R316 B.n346 B.n6 585
R317 B.n412 B.n6 585
R318 B.n345 B.n5 585
R319 B.n413 B.n5 585
R320 B.n344 B.n343 585
R321 B.n343 B.n4 585
R322 B.n342 B.n143 585
R323 B.n342 B.n341 585
R324 B.n331 B.n144 585
R325 B.n334 B.n144 585
R326 B.n333 B.n332 585
R327 B.n335 B.n333 585
R328 B.n330 B.n148 585
R329 B.n151 B.n148 585
R330 B.n329 B.n328 585
R331 B.n328 B.n327 585
R332 B.n150 B.n149 585
R333 B.n320 B.n150 585
R334 B.n319 B.n318 585
R335 B.n321 B.n319 585
R336 B.n317 B.n155 585
R337 B.n159 B.n155 585
R338 B.n316 B.n315 585
R339 B.n315 B.n314 585
R340 B.n157 B.n156 585
R341 B.n158 B.n157 585
R342 B.n307 B.n306 585
R343 B.n308 B.n307 585
R344 B.n305 B.n164 585
R345 B.n164 B.n163 585
R346 B.n304 B.n303 585
R347 B.n303 B.n302 585
R348 B.n166 B.n165 585
R349 B.t11 B.n166 585
R350 B.n295 B.n294 585
R351 B.n296 B.n295 585
R352 B.n293 B.n171 585
R353 B.n171 B.n170 585
R354 B.n292 B.n291 585
R355 B.n291 B.n290 585
R356 B.n173 B.n172 585
R357 B.n174 B.n173 585
R358 B.n286 B.n285 585
R359 B.n177 B.n176 585
R360 B.n282 B.n281 585
R361 B.n283 B.n282 585
R362 B.n280 B.n198 585
R363 B.n279 B.n278 585
R364 B.n277 B.n276 585
R365 B.n275 B.n274 585
R366 B.n273 B.n272 585
R367 B.n271 B.n270 585
R368 B.n269 B.n268 585
R369 B.n267 B.n266 585
R370 B.n265 B.n264 585
R371 B.n263 B.n262 585
R372 B.n261 B.n260 585
R373 B.n259 B.n258 585
R374 B.n257 B.n256 585
R375 B.n254 B.n253 585
R376 B.n252 B.n251 585
R377 B.n250 B.n249 585
R378 B.n248 B.n247 585
R379 B.n246 B.n245 585
R380 B.n244 B.n243 585
R381 B.n242 B.n241 585
R382 B.n240 B.n239 585
R383 B.n238 B.n237 585
R384 B.n236 B.n235 585
R385 B.n233 B.n232 585
R386 B.n231 B.n230 585
R387 B.n229 B.n228 585
R388 B.n227 B.n226 585
R389 B.n225 B.n224 585
R390 B.n223 B.n222 585
R391 B.n221 B.n220 585
R392 B.n219 B.n218 585
R393 B.n217 B.n216 585
R394 B.n215 B.n214 585
R395 B.n213 B.n212 585
R396 B.n211 B.n210 585
R397 B.n209 B.n208 585
R398 B.n207 B.n206 585
R399 B.n205 B.n204 585
R400 B.n203 B.n197 585
R401 B.n283 B.n197 585
R402 B.n287 B.n175 585
R403 B.n175 B.n174 585
R404 B.n289 B.n288 585
R405 B.n290 B.n289 585
R406 B.n169 B.n168 585
R407 B.n170 B.n169 585
R408 B.n298 B.n297 585
R409 B.n297 B.n296 585
R410 B.n299 B.n167 585
R411 B.n167 B.t11 585
R412 B.n301 B.n300 585
R413 B.n302 B.n301 585
R414 B.n162 B.n161 585
R415 B.n163 B.n162 585
R416 B.n310 B.n309 585
R417 B.n309 B.n308 585
R418 B.n311 B.n160 585
R419 B.n160 B.n158 585
R420 B.n313 B.n312 585
R421 B.n314 B.n313 585
R422 B.n154 B.n153 585
R423 B.n159 B.n154 585
R424 B.n323 B.n322 585
R425 B.n322 B.n321 585
R426 B.n324 B.n152 585
R427 B.n320 B.n152 585
R428 B.n326 B.n325 585
R429 B.n327 B.n326 585
R430 B.n147 B.n146 585
R431 B.n151 B.n147 585
R432 B.n337 B.n336 585
R433 B.n336 B.n335 585
R434 B.n338 B.n145 585
R435 B.n334 B.n145 585
R436 B.n340 B.n339 585
R437 B.n341 B.n340 585
R438 B.n2 B.n0 585
R439 B.n4 B.n2 585
R440 B.n3 B.n1 585
R441 B.n412 B.n3 585
R442 B.n410 B.n409 585
R443 B.n411 B.n410 585
R444 B.n408 B.n8 585
R445 B.n11 B.n8 585
R446 B.n407 B.n406 585
R447 B.n406 B.n405 585
R448 B.n10 B.n9 585
R449 B.n404 B.n10 585
R450 B.n402 B.n401 585
R451 B.n403 B.n402 585
R452 B.n400 B.n15 585
R453 B.n18 B.n15 585
R454 B.n399 B.n398 585
R455 B.n398 B.n397 585
R456 B.n17 B.n16 585
R457 B.n396 B.n17 585
R458 B.n394 B.n393 585
R459 B.n395 B.n394 585
R460 B.n392 B.n23 585
R461 B.n23 B.n22 585
R462 B.n391 B.n390 585
R463 B.n390 B.n389 585
R464 B.n25 B.n24 585
R465 B.n388 B.n25 585
R466 B.n386 B.n385 585
R467 B.n387 B.n386 585
R468 B.n384 B.n29 585
R469 B.n29 B.t18 585
R470 B.n383 B.n382 585
R471 B.n382 B.n381 585
R472 B.n31 B.n30 585
R473 B.n380 B.n31 585
R474 B.n378 B.n377 585
R475 B.n379 B.n378 585
R476 B.n376 B.n36 585
R477 B.n36 B.n35 585
R478 B.n415 B.n414 585
R479 B.n414 B.n413 585
R480 B.n285 B.n175 526.135
R481 B.n374 B.n36 526.135
R482 B.n197 B.n173 526.135
R483 B.n370 B.n59 526.135
R484 B.n201 B.t10 484.58
R485 B.n199 B.t14 484.58
R486 B.n63 B.t21 484.58
R487 B.n60 B.t17 484.58
R488 B.n372 B.n371 256.663
R489 B.n372 B.n57 256.663
R490 B.n372 B.n56 256.663
R491 B.n372 B.n55 256.663
R492 B.n372 B.n54 256.663
R493 B.n372 B.n53 256.663
R494 B.n372 B.n52 256.663
R495 B.n372 B.n51 256.663
R496 B.n372 B.n50 256.663
R497 B.n372 B.n49 256.663
R498 B.n372 B.n48 256.663
R499 B.n372 B.n47 256.663
R500 B.n372 B.n46 256.663
R501 B.n372 B.n45 256.663
R502 B.n372 B.n44 256.663
R503 B.n372 B.n43 256.663
R504 B.n372 B.n42 256.663
R505 B.n372 B.n41 256.663
R506 B.n372 B.n40 256.663
R507 B.n372 B.n39 256.663
R508 B.n373 B.n372 256.663
R509 B.n284 B.n283 256.663
R510 B.n283 B.n178 256.663
R511 B.n283 B.n179 256.663
R512 B.n283 B.n180 256.663
R513 B.n283 B.n181 256.663
R514 B.n283 B.n182 256.663
R515 B.n283 B.n183 256.663
R516 B.n283 B.n184 256.663
R517 B.n283 B.n185 256.663
R518 B.n283 B.n186 256.663
R519 B.n283 B.n187 256.663
R520 B.n283 B.n188 256.663
R521 B.n283 B.n189 256.663
R522 B.n283 B.n190 256.663
R523 B.n283 B.n191 256.663
R524 B.n283 B.n192 256.663
R525 B.n283 B.n193 256.663
R526 B.n283 B.n194 256.663
R527 B.n283 B.n195 256.663
R528 B.n283 B.n196 256.663
R529 B.n283 B.n174 177.482
R530 B.n372 B.n35 177.482
R531 B.n289 B.n175 163.367
R532 B.n289 B.n169 163.367
R533 B.n297 B.n169 163.367
R534 B.n297 B.n167 163.367
R535 B.n301 B.n167 163.367
R536 B.n301 B.n162 163.367
R537 B.n309 B.n162 163.367
R538 B.n309 B.n160 163.367
R539 B.n313 B.n160 163.367
R540 B.n313 B.n154 163.367
R541 B.n322 B.n154 163.367
R542 B.n322 B.n152 163.367
R543 B.n326 B.n152 163.367
R544 B.n326 B.n147 163.367
R545 B.n336 B.n147 163.367
R546 B.n336 B.n145 163.367
R547 B.n340 B.n145 163.367
R548 B.n340 B.n2 163.367
R549 B.n414 B.n2 163.367
R550 B.n414 B.n3 163.367
R551 B.n410 B.n3 163.367
R552 B.n410 B.n8 163.367
R553 B.n406 B.n8 163.367
R554 B.n406 B.n10 163.367
R555 B.n402 B.n10 163.367
R556 B.n402 B.n15 163.367
R557 B.n398 B.n15 163.367
R558 B.n398 B.n17 163.367
R559 B.n394 B.n17 163.367
R560 B.n394 B.n23 163.367
R561 B.n390 B.n23 163.367
R562 B.n390 B.n25 163.367
R563 B.n386 B.n25 163.367
R564 B.n386 B.n29 163.367
R565 B.n382 B.n29 163.367
R566 B.n382 B.n31 163.367
R567 B.n378 B.n31 163.367
R568 B.n378 B.n36 163.367
R569 B.n282 B.n177 163.367
R570 B.n282 B.n198 163.367
R571 B.n278 B.n277 163.367
R572 B.n274 B.n273 163.367
R573 B.n270 B.n269 163.367
R574 B.n266 B.n265 163.367
R575 B.n262 B.n261 163.367
R576 B.n258 B.n257 163.367
R577 B.n253 B.n252 163.367
R578 B.n249 B.n248 163.367
R579 B.n245 B.n244 163.367
R580 B.n241 B.n240 163.367
R581 B.n237 B.n236 163.367
R582 B.n232 B.n231 163.367
R583 B.n228 B.n227 163.367
R584 B.n224 B.n223 163.367
R585 B.n220 B.n219 163.367
R586 B.n216 B.n215 163.367
R587 B.n212 B.n211 163.367
R588 B.n208 B.n207 163.367
R589 B.n204 B.n197 163.367
R590 B.n291 B.n173 163.367
R591 B.n291 B.n171 163.367
R592 B.n295 B.n171 163.367
R593 B.n295 B.n166 163.367
R594 B.n303 B.n166 163.367
R595 B.n303 B.n164 163.367
R596 B.n307 B.n164 163.367
R597 B.n307 B.n157 163.367
R598 B.n315 B.n157 163.367
R599 B.n315 B.n155 163.367
R600 B.n319 B.n155 163.367
R601 B.n319 B.n150 163.367
R602 B.n328 B.n150 163.367
R603 B.n328 B.n148 163.367
R604 B.n333 B.n148 163.367
R605 B.n333 B.n144 163.367
R606 B.n342 B.n144 163.367
R607 B.n343 B.n342 163.367
R608 B.n343 B.n5 163.367
R609 B.n6 B.n5 163.367
R610 B.n7 B.n6 163.367
R611 B.n348 B.n7 163.367
R612 B.n348 B.n12 163.367
R613 B.n13 B.n12 163.367
R614 B.n14 B.n13 163.367
R615 B.n353 B.n14 163.367
R616 B.n353 B.n19 163.367
R617 B.n20 B.n19 163.367
R618 B.n21 B.n20 163.367
R619 B.n358 B.n21 163.367
R620 B.n358 B.n26 163.367
R621 B.n27 B.n26 163.367
R622 B.n28 B.n27 163.367
R623 B.n363 B.n28 163.367
R624 B.n363 B.n32 163.367
R625 B.n33 B.n32 163.367
R626 B.n34 B.n33 163.367
R627 B.n59 B.n34 163.367
R628 B.n66 B.n38 163.367
R629 B.n70 B.n69 163.367
R630 B.n74 B.n73 163.367
R631 B.n78 B.n77 163.367
R632 B.n82 B.n81 163.367
R633 B.n86 B.n85 163.367
R634 B.n90 B.n89 163.367
R635 B.n94 B.n93 163.367
R636 B.n98 B.n97 163.367
R637 B.n102 B.n101 163.367
R638 B.n106 B.n105 163.367
R639 B.n110 B.n109 163.367
R640 B.n114 B.n113 163.367
R641 B.n118 B.n117 163.367
R642 B.n122 B.n121 163.367
R643 B.n126 B.n125 163.367
R644 B.n130 B.n129 163.367
R645 B.n134 B.n133 163.367
R646 B.n138 B.n137 163.367
R647 B.n140 B.n58 163.367
R648 B.n201 B.t13 147.113
R649 B.n60 B.t19 147.113
R650 B.n199 B.t16 147.113
R651 B.n63 B.t22 147.113
R652 B.n202 B.t12 134.894
R653 B.n61 B.t20 134.894
R654 B.n200 B.t15 134.894
R655 B.n64 B.t23 134.894
R656 B.n290 B.n174 86.8258
R657 B.n290 B.n170 86.8258
R658 B.n296 B.n170 86.8258
R659 B.n296 B.t11 86.8258
R660 B.n302 B.t11 86.8258
R661 B.n302 B.n163 86.8258
R662 B.n308 B.n163 86.8258
R663 B.n308 B.n158 86.8258
R664 B.n314 B.n158 86.8258
R665 B.n321 B.n320 86.8258
R666 B.n327 B.n151 86.8258
R667 B.n335 B.n334 86.8258
R668 B.n341 B.n4 86.8258
R669 B.n413 B.n4 86.8258
R670 B.n413 B.n412 86.8258
R671 B.n412 B.n411 86.8258
R672 B.n405 B.n11 86.8258
R673 B.n404 B.n403 86.8258
R674 B.n397 B.n18 86.8258
R675 B.n395 B.n22 86.8258
R676 B.n389 B.n22 86.8258
R677 B.n389 B.n388 86.8258
R678 B.n388 B.n387 86.8258
R679 B.n387 B.t18 86.8258
R680 B.n381 B.t18 86.8258
R681 B.n381 B.n380 86.8258
R682 B.n380 B.n379 86.8258
R683 B.n379 B.n35 86.8258
R684 B.t8 B.n159 81.7184
R685 B.n396 B.t9 81.7184
R686 B.n159 B.t1 79.1648
R687 B.t2 B.n396 79.1648
R688 B.n285 B.n284 71.676
R689 B.n198 B.n178 71.676
R690 B.n277 B.n179 71.676
R691 B.n273 B.n180 71.676
R692 B.n269 B.n181 71.676
R693 B.n265 B.n182 71.676
R694 B.n261 B.n183 71.676
R695 B.n257 B.n184 71.676
R696 B.n252 B.n185 71.676
R697 B.n248 B.n186 71.676
R698 B.n244 B.n187 71.676
R699 B.n240 B.n188 71.676
R700 B.n236 B.n189 71.676
R701 B.n231 B.n190 71.676
R702 B.n227 B.n191 71.676
R703 B.n223 B.n192 71.676
R704 B.n219 B.n193 71.676
R705 B.n215 B.n194 71.676
R706 B.n211 B.n195 71.676
R707 B.n207 B.n196 71.676
R708 B.n374 B.n373 71.676
R709 B.n66 B.n39 71.676
R710 B.n70 B.n40 71.676
R711 B.n74 B.n41 71.676
R712 B.n78 B.n42 71.676
R713 B.n82 B.n43 71.676
R714 B.n86 B.n44 71.676
R715 B.n90 B.n45 71.676
R716 B.n94 B.n46 71.676
R717 B.n98 B.n47 71.676
R718 B.n102 B.n48 71.676
R719 B.n106 B.n49 71.676
R720 B.n110 B.n50 71.676
R721 B.n114 B.n51 71.676
R722 B.n118 B.n52 71.676
R723 B.n122 B.n53 71.676
R724 B.n126 B.n54 71.676
R725 B.n130 B.n55 71.676
R726 B.n134 B.n56 71.676
R727 B.n138 B.n57 71.676
R728 B.n371 B.n58 71.676
R729 B.n371 B.n370 71.676
R730 B.n140 B.n57 71.676
R731 B.n137 B.n56 71.676
R732 B.n133 B.n55 71.676
R733 B.n129 B.n54 71.676
R734 B.n125 B.n53 71.676
R735 B.n121 B.n52 71.676
R736 B.n117 B.n51 71.676
R737 B.n113 B.n50 71.676
R738 B.n109 B.n49 71.676
R739 B.n105 B.n48 71.676
R740 B.n101 B.n47 71.676
R741 B.n97 B.n46 71.676
R742 B.n93 B.n45 71.676
R743 B.n89 B.n44 71.676
R744 B.n85 B.n43 71.676
R745 B.n81 B.n42 71.676
R746 B.n77 B.n41 71.676
R747 B.n73 B.n40 71.676
R748 B.n69 B.n39 71.676
R749 B.n373 B.n38 71.676
R750 B.n284 B.n177 71.676
R751 B.n278 B.n178 71.676
R752 B.n274 B.n179 71.676
R753 B.n270 B.n180 71.676
R754 B.n266 B.n181 71.676
R755 B.n262 B.n182 71.676
R756 B.n258 B.n183 71.676
R757 B.n253 B.n184 71.676
R758 B.n249 B.n185 71.676
R759 B.n245 B.n186 71.676
R760 B.n241 B.n187 71.676
R761 B.n237 B.n188 71.676
R762 B.n232 B.n189 71.676
R763 B.n228 B.n190 71.676
R764 B.n224 B.n191 71.676
R765 B.n220 B.n192 71.676
R766 B.n216 B.n193 71.676
R767 B.n212 B.n194 71.676
R768 B.n208 B.n195 71.676
R769 B.n204 B.n196 71.676
R770 B.n320 B.t6 66.3963
R771 B.n18 B.t4 66.3963
R772 B.n234 B.n202 59.5399
R773 B.n255 B.n200 59.5399
R774 B.n65 B.n64 59.5399
R775 B.n62 B.n61 59.5399
R776 B.n151 B.t7 53.6279
R777 B.t3 B.n404 53.6279
R778 B.n341 B.t5 45.9668
R779 B.n411 B.t0 45.9668
R780 B.n334 B.t5 40.8595
R781 B.n11 B.t0 40.8595
R782 B.n376 B.n375 34.1859
R783 B.n369 B.n368 34.1859
R784 B.n203 B.n172 34.1859
R785 B.n287 B.n286 34.1859
R786 B.n335 B.t7 33.1984
R787 B.n405 B.t3 33.1984
R788 B.n327 B.t6 20.43
R789 B.n403 B.t4 20.43
R790 B B.n415 18.0485
R791 B.n202 B.n201 12.2187
R792 B.n200 B.n199 12.2187
R793 B.n64 B.n63 12.2187
R794 B.n61 B.n60 12.2187
R795 B.n375 B.n37 10.6151
R796 B.n67 B.n37 10.6151
R797 B.n68 B.n67 10.6151
R798 B.n71 B.n68 10.6151
R799 B.n72 B.n71 10.6151
R800 B.n75 B.n72 10.6151
R801 B.n76 B.n75 10.6151
R802 B.n79 B.n76 10.6151
R803 B.n80 B.n79 10.6151
R804 B.n83 B.n80 10.6151
R805 B.n84 B.n83 10.6151
R806 B.n87 B.n84 10.6151
R807 B.n88 B.n87 10.6151
R808 B.n91 B.n88 10.6151
R809 B.n92 B.n91 10.6151
R810 B.n96 B.n95 10.6151
R811 B.n99 B.n96 10.6151
R812 B.n100 B.n99 10.6151
R813 B.n103 B.n100 10.6151
R814 B.n104 B.n103 10.6151
R815 B.n107 B.n104 10.6151
R816 B.n108 B.n107 10.6151
R817 B.n111 B.n108 10.6151
R818 B.n112 B.n111 10.6151
R819 B.n116 B.n115 10.6151
R820 B.n119 B.n116 10.6151
R821 B.n120 B.n119 10.6151
R822 B.n123 B.n120 10.6151
R823 B.n124 B.n123 10.6151
R824 B.n127 B.n124 10.6151
R825 B.n128 B.n127 10.6151
R826 B.n131 B.n128 10.6151
R827 B.n132 B.n131 10.6151
R828 B.n135 B.n132 10.6151
R829 B.n136 B.n135 10.6151
R830 B.n139 B.n136 10.6151
R831 B.n141 B.n139 10.6151
R832 B.n142 B.n141 10.6151
R833 B.n369 B.n142 10.6151
R834 B.n292 B.n172 10.6151
R835 B.n293 B.n292 10.6151
R836 B.n294 B.n293 10.6151
R837 B.n294 B.n165 10.6151
R838 B.n304 B.n165 10.6151
R839 B.n305 B.n304 10.6151
R840 B.n306 B.n305 10.6151
R841 B.n306 B.n156 10.6151
R842 B.n316 B.n156 10.6151
R843 B.n317 B.n316 10.6151
R844 B.n318 B.n317 10.6151
R845 B.n318 B.n149 10.6151
R846 B.n329 B.n149 10.6151
R847 B.n330 B.n329 10.6151
R848 B.n332 B.n330 10.6151
R849 B.n332 B.n331 10.6151
R850 B.n331 B.n143 10.6151
R851 B.n344 B.n143 10.6151
R852 B.n345 B.n344 10.6151
R853 B.n346 B.n345 10.6151
R854 B.n347 B.n346 10.6151
R855 B.n349 B.n347 10.6151
R856 B.n350 B.n349 10.6151
R857 B.n351 B.n350 10.6151
R858 B.n352 B.n351 10.6151
R859 B.n354 B.n352 10.6151
R860 B.n355 B.n354 10.6151
R861 B.n356 B.n355 10.6151
R862 B.n357 B.n356 10.6151
R863 B.n359 B.n357 10.6151
R864 B.n360 B.n359 10.6151
R865 B.n361 B.n360 10.6151
R866 B.n362 B.n361 10.6151
R867 B.n364 B.n362 10.6151
R868 B.n365 B.n364 10.6151
R869 B.n366 B.n365 10.6151
R870 B.n367 B.n366 10.6151
R871 B.n368 B.n367 10.6151
R872 B.n286 B.n176 10.6151
R873 B.n281 B.n176 10.6151
R874 B.n281 B.n280 10.6151
R875 B.n280 B.n279 10.6151
R876 B.n279 B.n276 10.6151
R877 B.n276 B.n275 10.6151
R878 B.n275 B.n272 10.6151
R879 B.n272 B.n271 10.6151
R880 B.n271 B.n268 10.6151
R881 B.n268 B.n267 10.6151
R882 B.n267 B.n264 10.6151
R883 B.n264 B.n263 10.6151
R884 B.n263 B.n260 10.6151
R885 B.n260 B.n259 10.6151
R886 B.n259 B.n256 10.6151
R887 B.n254 B.n251 10.6151
R888 B.n251 B.n250 10.6151
R889 B.n250 B.n247 10.6151
R890 B.n247 B.n246 10.6151
R891 B.n246 B.n243 10.6151
R892 B.n243 B.n242 10.6151
R893 B.n242 B.n239 10.6151
R894 B.n239 B.n238 10.6151
R895 B.n238 B.n235 10.6151
R896 B.n233 B.n230 10.6151
R897 B.n230 B.n229 10.6151
R898 B.n229 B.n226 10.6151
R899 B.n226 B.n225 10.6151
R900 B.n225 B.n222 10.6151
R901 B.n222 B.n221 10.6151
R902 B.n221 B.n218 10.6151
R903 B.n218 B.n217 10.6151
R904 B.n217 B.n214 10.6151
R905 B.n214 B.n213 10.6151
R906 B.n213 B.n210 10.6151
R907 B.n210 B.n209 10.6151
R908 B.n209 B.n206 10.6151
R909 B.n206 B.n205 10.6151
R910 B.n205 B.n203 10.6151
R911 B.n288 B.n287 10.6151
R912 B.n288 B.n168 10.6151
R913 B.n298 B.n168 10.6151
R914 B.n299 B.n298 10.6151
R915 B.n300 B.n299 10.6151
R916 B.n300 B.n161 10.6151
R917 B.n310 B.n161 10.6151
R918 B.n311 B.n310 10.6151
R919 B.n312 B.n311 10.6151
R920 B.n312 B.n153 10.6151
R921 B.n323 B.n153 10.6151
R922 B.n324 B.n323 10.6151
R923 B.n325 B.n324 10.6151
R924 B.n325 B.n146 10.6151
R925 B.n337 B.n146 10.6151
R926 B.n338 B.n337 10.6151
R927 B.n339 B.n338 10.6151
R928 B.n339 B.n0 10.6151
R929 B.n409 B.n1 10.6151
R930 B.n409 B.n408 10.6151
R931 B.n408 B.n407 10.6151
R932 B.n407 B.n9 10.6151
R933 B.n401 B.n9 10.6151
R934 B.n401 B.n400 10.6151
R935 B.n400 B.n399 10.6151
R936 B.n399 B.n16 10.6151
R937 B.n393 B.n16 10.6151
R938 B.n393 B.n392 10.6151
R939 B.n392 B.n391 10.6151
R940 B.n391 B.n24 10.6151
R941 B.n385 B.n24 10.6151
R942 B.n385 B.n384 10.6151
R943 B.n384 B.n383 10.6151
R944 B.n383 B.n30 10.6151
R945 B.n377 B.n30 10.6151
R946 B.n377 B.n376 10.6151
R947 B.n92 B.n65 9.36635
R948 B.n115 B.n62 9.36635
R949 B.n256 B.n255 9.36635
R950 B.n234 B.n233 9.36635
R951 B.n321 B.t1 7.66156
R952 B.n397 B.t2 7.66156
R953 B.n314 B.t8 5.10787
R954 B.t9 B.n395 5.10787
R955 B.n415 B.n0 2.81026
R956 B.n415 B.n1 2.81026
R957 B.n95 B.n65 1.24928
R958 B.n112 B.n62 1.24928
R959 B.n255 B.n254 1.24928
R960 B.n235 B.n234 1.24928
R961 VN.n9 VN.t7 410.723
R962 VN.n3 VN.t4 410.723
R963 VN.n20 VN.t8 410.723
R964 VN.n14 VN.t6 410.723
R965 VN.n6 VN.t3 372.748
R966 VN.n8 VN.t1 372.748
R967 VN.n2 VN.t2 372.748
R968 VN.n17 VN.t0 372.748
R969 VN.n19 VN.t5 372.748
R970 VN.n13 VN.t9 372.748
R971 VN.n15 VN.n14 161.489
R972 VN.n4 VN.n3 161.489
R973 VN.n10 VN.n9 161.3
R974 VN.n21 VN.n20 161.3
R975 VN.n18 VN.n11 161.3
R976 VN.n17 VN.n16 161.3
R977 VN.n15 VN.n12 161.3
R978 VN.n7 VN.n0 161.3
R979 VN.n6 VN.n5 161.3
R980 VN.n4 VN.n1 161.3
R981 VN.n6 VN.n1 73.0308
R982 VN.n7 VN.n6 73.0308
R983 VN.n18 VN.n17 73.0308
R984 VN.n17 VN.n12 73.0308
R985 VN.n3 VN.n2 54.0429
R986 VN.n9 VN.n8 54.0429
R987 VN.n20 VN.n19 54.0429
R988 VN.n14 VN.n13 54.0429
R989 VN VN.n21 34.4835
R990 VN.n2 VN.n1 18.9884
R991 VN.n8 VN.n7 18.9884
R992 VN.n19 VN.n18 18.9884
R993 VN.n13 VN.n12 18.9884
R994 VN.n21 VN.n11 0.189894
R995 VN.n16 VN.n11 0.189894
R996 VN.n16 VN.n15 0.189894
R997 VN.n5 VN.n4 0.189894
R998 VN.n5 VN.n0 0.189894
R999 VN.n10 VN.n0 0.189894
R1000 VN VN.n10 0.0516364
R1001 VDD2.n29 VDD2.n19 289.615
R1002 VDD2.n10 VDD2.n0 289.615
R1003 VDD2.n30 VDD2.n29 185
R1004 VDD2.n28 VDD2.n27 185
R1005 VDD2.n23 VDD2.n22 185
R1006 VDD2.n4 VDD2.n3 185
R1007 VDD2.n9 VDD2.n8 185
R1008 VDD2.n11 VDD2.n10 185
R1009 VDD2.n24 VDD2.t1 148.606
R1010 VDD2.n5 VDD2.t5 148.606
R1011 VDD2.n29 VDD2.n28 104.615
R1012 VDD2.n28 VDD2.n22 104.615
R1013 VDD2.n9 VDD2.n3 104.615
R1014 VDD2.n10 VDD2.n9 104.615
R1015 VDD2.n18 VDD2.n17 82.3677
R1016 VDD2 VDD2.n37 82.3649
R1017 VDD2.n36 VDD2.n35 82.0159
R1018 VDD2.n16 VDD2.n15 82.0157
R1019 VDD2.n16 VDD2.n14 53.6739
R1020 VDD2.n34 VDD2.n33 53.1308
R1021 VDD2.t1 VDD2.n22 52.3082
R1022 VDD2.t5 VDD2.n3 52.3082
R1023 VDD2.n34 VDD2.n18 29.1743
R1024 VDD2.n24 VDD2.n23 15.5966
R1025 VDD2.n5 VDD2.n4 15.5966
R1026 VDD2.n27 VDD2.n26 12.8005
R1027 VDD2.n8 VDD2.n7 12.8005
R1028 VDD2.n30 VDD2.n21 12.0247
R1029 VDD2.n11 VDD2.n2 12.0247
R1030 VDD2.n31 VDD2.n19 11.249
R1031 VDD2.n12 VDD2.n0 11.249
R1032 VDD2.n33 VDD2.n32 9.45567
R1033 VDD2.n14 VDD2.n13 9.45567
R1034 VDD2.n32 VDD2.n31 9.3005
R1035 VDD2.n21 VDD2.n20 9.3005
R1036 VDD2.n26 VDD2.n25 9.3005
R1037 VDD2.n13 VDD2.n12 9.3005
R1038 VDD2.n2 VDD2.n1 9.3005
R1039 VDD2.n7 VDD2.n6 9.3005
R1040 VDD2.n37 VDD2.t0 5.92864
R1041 VDD2.n37 VDD2.t3 5.92864
R1042 VDD2.n35 VDD2.t4 5.92864
R1043 VDD2.n35 VDD2.t9 5.92864
R1044 VDD2.n17 VDD2.t8 5.92864
R1045 VDD2.n17 VDD2.t2 5.92864
R1046 VDD2.n15 VDD2.t7 5.92864
R1047 VDD2.n15 VDD2.t6 5.92864
R1048 VDD2.n25 VDD2.n24 4.46457
R1049 VDD2.n6 VDD2.n5 4.46457
R1050 VDD2.n33 VDD2.n19 2.71565
R1051 VDD2.n14 VDD2.n0 2.71565
R1052 VDD2.n31 VDD2.n30 1.93989
R1053 VDD2.n12 VDD2.n11 1.93989
R1054 VDD2.n27 VDD2.n21 1.16414
R1055 VDD2.n8 VDD2.n2 1.16414
R1056 VDD2.n36 VDD2.n34 0.543603
R1057 VDD2.n26 VDD2.n23 0.388379
R1058 VDD2.n7 VDD2.n4 0.388379
R1059 VDD2 VDD2.n36 0.194466
R1060 VDD2.n32 VDD2.n20 0.155672
R1061 VDD2.n25 VDD2.n20 0.155672
R1062 VDD2.n6 VDD2.n1 0.155672
R1063 VDD2.n13 VDD2.n1 0.155672
R1064 VDD2.n18 VDD2.n16 0.0809298
C0 VTAIL VN 1.42649f
C1 VDD1 VP 1.52939f
C2 VN VP 3.40791f
C3 VDD1 VDD2 0.722519f
C4 VN VDD2 1.38987f
C5 VTAIL VP 1.44078f
C6 VTAIL VDD2 7.36558f
C7 VDD2 VP 0.29474f
C8 VN VDD1 0.153199f
C9 VTAIL VDD1 7.32972f
C10 VDD2 B 2.901836f
C11 VDD1 B 2.833891f
C12 VTAIL B 2.914506f
C13 VN B 5.834501f
C14 VP B 4.869313f
C15 VDD2.n0 B 0.035314f
C16 VDD2.n1 B 0.024421f
C17 VDD2.n2 B 0.013123f
C18 VDD2.n3 B 0.023263f
C19 VDD2.n4 B 0.018086f
C20 VDD2.t5 B 0.053007f
C21 VDD2.n5 B 0.09255f
C22 VDD2.n6 B 0.276584f
C23 VDD2.n7 B 0.013123f
C24 VDD2.n8 B 0.013895f
C25 VDD2.n9 B 0.031017f
C26 VDD2.n10 B 0.068895f
C27 VDD2.n11 B 0.013895f
C28 VDD2.n12 B 0.013123f
C29 VDD2.n13 B 0.063786f
C30 VDD2.n14 B 0.056705f
C31 VDD2.t7 B 0.064455f
C32 VDD2.t6 B 0.064455f
C33 VDD2.n15 B 0.487579f
C34 VDD2.n16 B 0.336977f
C35 VDD2.t8 B 0.064455f
C36 VDD2.t2 B 0.064455f
C37 VDD2.n17 B 0.488731f
C38 VDD2.n18 B 1.14136f
C39 VDD2.n19 B 0.035314f
C40 VDD2.n20 B 0.024421f
C41 VDD2.n21 B 0.013123f
C42 VDD2.n22 B 0.023263f
C43 VDD2.n23 B 0.018086f
C44 VDD2.t1 B 0.053007f
C45 VDD2.n24 B 0.09255f
C46 VDD2.n25 B 0.276584f
C47 VDD2.n26 B 0.013123f
C48 VDD2.n27 B 0.013895f
C49 VDD2.n28 B 0.031017f
C50 VDD2.n29 B 0.068895f
C51 VDD2.n30 B 0.013895f
C52 VDD2.n31 B 0.013123f
C53 VDD2.n32 B 0.063786f
C54 VDD2.n33 B 0.055754f
C55 VDD2.n34 B 1.27744f
C56 VDD2.t4 B 0.064455f
C57 VDD2.t9 B 0.064455f
C58 VDD2.n35 B 0.487581f
C59 VDD2.n36 B 0.245857f
C60 VDD2.t0 B 0.064455f
C61 VDD2.t3 B 0.064455f
C62 VDD2.n37 B 0.488714f
C63 VN.n0 B 0.029156f
C64 VN.t1 B 0.084322f
C65 VN.t3 B 0.084322f
C66 VN.n1 B 0.012009f
C67 VN.t4 B 0.088758f
C68 VN.t2 B 0.084322f
C69 VN.n2 B 0.0469f
C70 VN.n3 B 0.055592f
C71 VN.n4 B 0.064022f
C72 VN.n5 B 0.029156f
C73 VN.n6 B 0.056572f
C74 VN.n7 B 0.012009f
C75 VN.n8 B 0.0469f
C76 VN.t7 B 0.088758f
C77 VN.n9 B 0.055551f
C78 VN.n10 B 0.022594f
C79 VN.n11 B 0.029156f
C80 VN.t8 B 0.088758f
C81 VN.t5 B 0.084322f
C82 VN.t0 B 0.084322f
C83 VN.n12 B 0.012009f
C84 VN.t9 B 0.084322f
C85 VN.n13 B 0.0469f
C86 VN.t6 B 0.088758f
C87 VN.n14 B 0.055592f
C88 VN.n15 B 0.064022f
C89 VN.n16 B 0.029156f
C90 VN.n17 B 0.056572f
C91 VN.n18 B 0.012009f
C92 VN.n19 B 0.0469f
C93 VN.n20 B 0.055551f
C94 VN.n21 B 0.845167f
C95 VTAIL.t0 B 0.073745f
C96 VTAIL.t3 B 0.073745f
C97 VTAIL.n0 B 0.504347f
C98 VTAIL.n1 B 0.339129f
C99 VTAIL.n2 B 0.040404f
C100 VTAIL.n3 B 0.027941f
C101 VTAIL.n4 B 0.015014f
C102 VTAIL.n5 B 0.026616f
C103 VTAIL.n6 B 0.020693f
C104 VTAIL.t14 B 0.060647f
C105 VTAIL.n7 B 0.105889f
C106 VTAIL.n8 B 0.31645f
C107 VTAIL.n9 B 0.015014f
C108 VTAIL.n10 B 0.015897f
C109 VTAIL.n11 B 0.035488f
C110 VTAIL.n12 B 0.078825f
C111 VTAIL.n13 B 0.015897f
C112 VTAIL.n14 B 0.015014f
C113 VTAIL.n15 B 0.072981f
C114 VTAIL.n16 B 0.044556f
C115 VTAIL.n17 B 0.144259f
C116 VTAIL.t13 B 0.073745f
C117 VTAIL.t8 B 0.073745f
C118 VTAIL.n18 B 0.504347f
C119 VTAIL.n19 B 0.328263f
C120 VTAIL.t10 B 0.073745f
C121 VTAIL.t16 B 0.073745f
C122 VTAIL.n20 B 0.504347f
C123 VTAIL.n21 B 1.01592f
C124 VTAIL.t18 B 0.073745f
C125 VTAIL.t1 B 0.073745f
C126 VTAIL.n22 B 0.50435f
C127 VTAIL.n23 B 1.01592f
C128 VTAIL.t6 B 0.073745f
C129 VTAIL.t19 B 0.073745f
C130 VTAIL.n24 B 0.50435f
C131 VTAIL.n25 B 0.32826f
C132 VTAIL.n26 B 0.040404f
C133 VTAIL.n27 B 0.027941f
C134 VTAIL.n28 B 0.015014f
C135 VTAIL.n29 B 0.026616f
C136 VTAIL.n30 B 0.020693f
C137 VTAIL.t5 B 0.060647f
C138 VTAIL.n31 B 0.105889f
C139 VTAIL.n32 B 0.31645f
C140 VTAIL.n33 B 0.015014f
C141 VTAIL.n34 B 0.015897f
C142 VTAIL.n35 B 0.035488f
C143 VTAIL.n36 B 0.078825f
C144 VTAIL.n37 B 0.015897f
C145 VTAIL.n38 B 0.015014f
C146 VTAIL.n39 B 0.072981f
C147 VTAIL.n40 B 0.044556f
C148 VTAIL.n41 B 0.144259f
C149 VTAIL.t15 B 0.073745f
C150 VTAIL.t11 B 0.073745f
C151 VTAIL.n42 B 0.50435f
C152 VTAIL.n43 B 0.346111f
C153 VTAIL.t9 B 0.073745f
C154 VTAIL.t7 B 0.073745f
C155 VTAIL.n44 B 0.50435f
C156 VTAIL.n45 B 0.32826f
C157 VTAIL.n46 B 0.040404f
C158 VTAIL.n47 B 0.027941f
C159 VTAIL.n48 B 0.015014f
C160 VTAIL.n49 B 0.026616f
C161 VTAIL.n50 B 0.020693f
C162 VTAIL.t12 B 0.060647f
C163 VTAIL.n51 B 0.105889f
C164 VTAIL.n52 B 0.31645f
C165 VTAIL.n53 B 0.015014f
C166 VTAIL.n54 B 0.015897f
C167 VTAIL.n55 B 0.035488f
C168 VTAIL.n56 B 0.078825f
C169 VTAIL.n57 B 0.015897f
C170 VTAIL.n58 B 0.015014f
C171 VTAIL.n59 B 0.072981f
C172 VTAIL.n60 B 0.044556f
C173 VTAIL.n61 B 0.765174f
C174 VTAIL.n62 B 0.040404f
C175 VTAIL.n63 B 0.027941f
C176 VTAIL.n64 B 0.015014f
C177 VTAIL.n65 B 0.026616f
C178 VTAIL.n66 B 0.020693f
C179 VTAIL.t17 B 0.060647f
C180 VTAIL.n67 B 0.105889f
C181 VTAIL.n68 B 0.31645f
C182 VTAIL.n69 B 0.015014f
C183 VTAIL.n70 B 0.015897f
C184 VTAIL.n71 B 0.035488f
C185 VTAIL.n72 B 0.078825f
C186 VTAIL.n73 B 0.015897f
C187 VTAIL.n74 B 0.015014f
C188 VTAIL.n75 B 0.072981f
C189 VTAIL.n76 B 0.044556f
C190 VTAIL.n77 B 0.765174f
C191 VTAIL.t4 B 0.073745f
C192 VTAIL.t2 B 0.073745f
C193 VTAIL.n78 B 0.504347f
C194 VTAIL.n79 B 0.286352f
C195 VDD1.n0 B 0.034417f
C196 VDD1.n1 B 0.023801f
C197 VDD1.n2 B 0.012789f
C198 VDD1.n3 B 0.022672f
C199 VDD1.n4 B 0.017627f
C200 VDD1.t9 B 0.051661f
C201 VDD1.n5 B 0.090199f
C202 VDD1.n6 B 0.269561f
C203 VDD1.n7 B 0.012789f
C204 VDD1.n8 B 0.013542f
C205 VDD1.n9 B 0.030229f
C206 VDD1.n10 B 0.067145f
C207 VDD1.n11 B 0.013542f
C208 VDD1.n12 B 0.012789f
C209 VDD1.n13 B 0.062167f
C210 VDD1.n14 B 0.055265f
C211 VDD1.t7 B 0.062818f
C212 VDD1.t6 B 0.062818f
C213 VDD1.n15 B 0.4752f
C214 VDD1.n16 B 0.330265f
C215 VDD1.n17 B 0.034417f
C216 VDD1.n18 B 0.023801f
C217 VDD1.n19 B 0.012789f
C218 VDD1.n20 B 0.022672f
C219 VDD1.n21 B 0.017627f
C220 VDD1.t8 B 0.051661f
C221 VDD1.n22 B 0.090199f
C222 VDD1.n23 B 0.269561f
C223 VDD1.n24 B 0.012789f
C224 VDD1.n25 B 0.013542f
C225 VDD1.n26 B 0.030229f
C226 VDD1.n27 B 0.067145f
C227 VDD1.n28 B 0.013542f
C228 VDD1.n29 B 0.012789f
C229 VDD1.n30 B 0.062167f
C230 VDD1.n31 B 0.055265f
C231 VDD1.t0 B 0.062818f
C232 VDD1.t5 B 0.062818f
C233 VDD1.n32 B 0.475198f
C234 VDD1.n33 B 0.32842f
C235 VDD1.t4 B 0.062818f
C236 VDD1.t1 B 0.062818f
C237 VDD1.n34 B 0.476321f
C238 VDD1.n35 B 1.17448f
C239 VDD1.t2 B 0.062818f
C240 VDD1.t3 B 0.062818f
C241 VDD1.n36 B 0.475198f
C242 VDD1.n37 B 1.44033f
C243 VP.n0 B 0.029511f
C244 VP.t8 B 0.085351f
C245 VP.t3 B 0.085351f
C246 VP.n1 B 0.012155f
C247 VP.n2 B 0.029511f
C248 VP.t9 B 0.085351f
C249 VP.t7 B 0.085351f
C250 VP.n3 B 0.012155f
C251 VP.t1 B 0.089841f
C252 VP.t5 B 0.085351f
C253 VP.n4 B 0.047472f
C254 VP.n5 B 0.05627f
C255 VP.n6 B 0.064803f
C256 VP.n7 B 0.029511f
C257 VP.n8 B 0.057262f
C258 VP.n9 B 0.012155f
C259 VP.n10 B 0.047472f
C260 VP.t4 B 0.089841f
C261 VP.n11 B 0.056229f
C262 VP.n12 B 0.835824f
C263 VP.t6 B 0.089841f
C264 VP.t0 B 0.085351f
C265 VP.n13 B 0.047472f
C266 VP.n14 B 0.056229f
C267 VP.n15 B 0.86702f
C268 VP.n16 B 0.029511f
C269 VP.n17 B 0.029511f
C270 VP.n18 B 0.057262f
C271 VP.n19 B 0.012155f
C272 VP.n20 B 0.047472f
C273 VP.t2 B 0.089841f
C274 VP.n21 B 0.056229f
C275 VP.n22 B 0.02287f
.ends

