* NGSPICE file created from diff_pair_sample_1027.ext - technology: sky130A

.subckt diff_pair_sample_1027 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1408_n3386# sky130_fd_pr__pfet_01v8 ad=4.7151 pd=24.96 as=0 ps=0 w=12.09 l=0.4
X1 VDD1.t3 VP.t0 VTAIL.t7 w_n1408_n3386# sky130_fd_pr__pfet_01v8 ad=1.99485 pd=12.42 as=4.7151 ps=24.96 w=12.09 l=0.4
X2 VTAIL.t0 VN.t0 VDD2.t3 w_n1408_n3386# sky130_fd_pr__pfet_01v8 ad=4.7151 pd=24.96 as=1.99485 ps=12.42 w=12.09 l=0.4
X3 VTAIL.t6 VP.t1 VDD1.t2 w_n1408_n3386# sky130_fd_pr__pfet_01v8 ad=4.7151 pd=24.96 as=1.99485 ps=12.42 w=12.09 l=0.4
X4 VDD1.t1 VP.t2 VTAIL.t5 w_n1408_n3386# sky130_fd_pr__pfet_01v8 ad=1.99485 pd=12.42 as=4.7151 ps=24.96 w=12.09 l=0.4
X5 VDD2.t2 VN.t1 VTAIL.t1 w_n1408_n3386# sky130_fd_pr__pfet_01v8 ad=1.99485 pd=12.42 as=4.7151 ps=24.96 w=12.09 l=0.4
X6 B.t8 B.t6 B.t7 w_n1408_n3386# sky130_fd_pr__pfet_01v8 ad=4.7151 pd=24.96 as=0 ps=0 w=12.09 l=0.4
X7 VTAIL.t4 VP.t3 VDD1.t0 w_n1408_n3386# sky130_fd_pr__pfet_01v8 ad=4.7151 pd=24.96 as=1.99485 ps=12.42 w=12.09 l=0.4
X8 B.t5 B.t3 B.t4 w_n1408_n3386# sky130_fd_pr__pfet_01v8 ad=4.7151 pd=24.96 as=0 ps=0 w=12.09 l=0.4
X9 B.t2 B.t0 B.t1 w_n1408_n3386# sky130_fd_pr__pfet_01v8 ad=4.7151 pd=24.96 as=0 ps=0 w=12.09 l=0.4
X10 VTAIL.t2 VN.t2 VDD2.t1 w_n1408_n3386# sky130_fd_pr__pfet_01v8 ad=4.7151 pd=24.96 as=1.99485 ps=12.42 w=12.09 l=0.4
X11 VDD2.t0 VN.t3 VTAIL.t3 w_n1408_n3386# sky130_fd_pr__pfet_01v8 ad=1.99485 pd=12.42 as=4.7151 ps=24.96 w=12.09 l=0.4
R0 B.n104 B.t0 937.843
R1 B.n96 B.t9 937.843
R2 B.n38 B.t6 937.843
R3 B.n30 B.t3 937.843
R4 B.n292 B.n75 585
R5 B.n291 B.n290 585
R6 B.n289 B.n76 585
R7 B.n288 B.n287 585
R8 B.n286 B.n77 585
R9 B.n285 B.n284 585
R10 B.n283 B.n78 585
R11 B.n282 B.n281 585
R12 B.n280 B.n79 585
R13 B.n279 B.n278 585
R14 B.n277 B.n80 585
R15 B.n276 B.n275 585
R16 B.n274 B.n81 585
R17 B.n273 B.n272 585
R18 B.n271 B.n82 585
R19 B.n270 B.n269 585
R20 B.n268 B.n83 585
R21 B.n267 B.n266 585
R22 B.n265 B.n84 585
R23 B.n264 B.n263 585
R24 B.n262 B.n85 585
R25 B.n261 B.n260 585
R26 B.n259 B.n86 585
R27 B.n258 B.n257 585
R28 B.n256 B.n87 585
R29 B.n255 B.n254 585
R30 B.n253 B.n88 585
R31 B.n252 B.n251 585
R32 B.n250 B.n89 585
R33 B.n249 B.n248 585
R34 B.n247 B.n90 585
R35 B.n246 B.n245 585
R36 B.n244 B.n91 585
R37 B.n243 B.n242 585
R38 B.n241 B.n92 585
R39 B.n240 B.n239 585
R40 B.n238 B.n93 585
R41 B.n237 B.n236 585
R42 B.n235 B.n94 585
R43 B.n234 B.n233 585
R44 B.n232 B.n95 585
R45 B.n231 B.n230 585
R46 B.n229 B.n228 585
R47 B.n227 B.n99 585
R48 B.n226 B.n225 585
R49 B.n224 B.n100 585
R50 B.n223 B.n222 585
R51 B.n221 B.n101 585
R52 B.n220 B.n219 585
R53 B.n218 B.n102 585
R54 B.n217 B.n216 585
R55 B.n214 B.n103 585
R56 B.n213 B.n212 585
R57 B.n211 B.n106 585
R58 B.n210 B.n209 585
R59 B.n208 B.n107 585
R60 B.n207 B.n206 585
R61 B.n205 B.n108 585
R62 B.n204 B.n203 585
R63 B.n202 B.n109 585
R64 B.n201 B.n200 585
R65 B.n199 B.n110 585
R66 B.n198 B.n197 585
R67 B.n196 B.n111 585
R68 B.n195 B.n194 585
R69 B.n193 B.n112 585
R70 B.n192 B.n191 585
R71 B.n190 B.n113 585
R72 B.n189 B.n188 585
R73 B.n187 B.n114 585
R74 B.n186 B.n185 585
R75 B.n184 B.n115 585
R76 B.n183 B.n182 585
R77 B.n181 B.n116 585
R78 B.n180 B.n179 585
R79 B.n178 B.n117 585
R80 B.n177 B.n176 585
R81 B.n175 B.n118 585
R82 B.n174 B.n173 585
R83 B.n172 B.n119 585
R84 B.n171 B.n170 585
R85 B.n169 B.n120 585
R86 B.n168 B.n167 585
R87 B.n166 B.n121 585
R88 B.n165 B.n164 585
R89 B.n163 B.n122 585
R90 B.n162 B.n161 585
R91 B.n160 B.n123 585
R92 B.n159 B.n158 585
R93 B.n157 B.n124 585
R94 B.n156 B.n155 585
R95 B.n154 B.n125 585
R96 B.n153 B.n152 585
R97 B.n294 B.n293 585
R98 B.n295 B.n74 585
R99 B.n297 B.n296 585
R100 B.n298 B.n73 585
R101 B.n300 B.n299 585
R102 B.n301 B.n72 585
R103 B.n303 B.n302 585
R104 B.n304 B.n71 585
R105 B.n306 B.n305 585
R106 B.n307 B.n70 585
R107 B.n309 B.n308 585
R108 B.n310 B.n69 585
R109 B.n312 B.n311 585
R110 B.n313 B.n68 585
R111 B.n315 B.n314 585
R112 B.n316 B.n67 585
R113 B.n318 B.n317 585
R114 B.n319 B.n66 585
R115 B.n321 B.n320 585
R116 B.n322 B.n65 585
R117 B.n324 B.n323 585
R118 B.n325 B.n64 585
R119 B.n327 B.n326 585
R120 B.n328 B.n63 585
R121 B.n330 B.n329 585
R122 B.n331 B.n62 585
R123 B.n333 B.n332 585
R124 B.n334 B.n61 585
R125 B.n336 B.n335 585
R126 B.n337 B.n60 585
R127 B.n478 B.n9 585
R128 B.n477 B.n476 585
R129 B.n475 B.n10 585
R130 B.n474 B.n473 585
R131 B.n472 B.n11 585
R132 B.n471 B.n470 585
R133 B.n469 B.n12 585
R134 B.n468 B.n467 585
R135 B.n466 B.n13 585
R136 B.n465 B.n464 585
R137 B.n463 B.n14 585
R138 B.n462 B.n461 585
R139 B.n460 B.n15 585
R140 B.n459 B.n458 585
R141 B.n457 B.n16 585
R142 B.n456 B.n455 585
R143 B.n454 B.n17 585
R144 B.n453 B.n452 585
R145 B.n451 B.n18 585
R146 B.n450 B.n449 585
R147 B.n448 B.n19 585
R148 B.n447 B.n446 585
R149 B.n445 B.n20 585
R150 B.n444 B.n443 585
R151 B.n442 B.n21 585
R152 B.n441 B.n440 585
R153 B.n439 B.n22 585
R154 B.n438 B.n437 585
R155 B.n436 B.n23 585
R156 B.n435 B.n434 585
R157 B.n433 B.n24 585
R158 B.n432 B.n431 585
R159 B.n430 B.n25 585
R160 B.n429 B.n428 585
R161 B.n427 B.n26 585
R162 B.n426 B.n425 585
R163 B.n424 B.n27 585
R164 B.n423 B.n422 585
R165 B.n421 B.n28 585
R166 B.n420 B.n419 585
R167 B.n418 B.n29 585
R168 B.n417 B.n416 585
R169 B.n415 B.n414 585
R170 B.n413 B.n33 585
R171 B.n412 B.n411 585
R172 B.n410 B.n34 585
R173 B.n409 B.n408 585
R174 B.n407 B.n35 585
R175 B.n406 B.n405 585
R176 B.n404 B.n36 585
R177 B.n403 B.n402 585
R178 B.n400 B.n37 585
R179 B.n399 B.n398 585
R180 B.n397 B.n40 585
R181 B.n396 B.n395 585
R182 B.n394 B.n41 585
R183 B.n393 B.n392 585
R184 B.n391 B.n42 585
R185 B.n390 B.n389 585
R186 B.n388 B.n43 585
R187 B.n387 B.n386 585
R188 B.n385 B.n44 585
R189 B.n384 B.n383 585
R190 B.n382 B.n45 585
R191 B.n381 B.n380 585
R192 B.n379 B.n46 585
R193 B.n378 B.n377 585
R194 B.n376 B.n47 585
R195 B.n375 B.n374 585
R196 B.n373 B.n48 585
R197 B.n372 B.n371 585
R198 B.n370 B.n49 585
R199 B.n369 B.n368 585
R200 B.n367 B.n50 585
R201 B.n366 B.n365 585
R202 B.n364 B.n51 585
R203 B.n363 B.n362 585
R204 B.n361 B.n52 585
R205 B.n360 B.n359 585
R206 B.n358 B.n53 585
R207 B.n357 B.n356 585
R208 B.n355 B.n54 585
R209 B.n354 B.n353 585
R210 B.n352 B.n55 585
R211 B.n351 B.n350 585
R212 B.n349 B.n56 585
R213 B.n348 B.n347 585
R214 B.n346 B.n57 585
R215 B.n345 B.n344 585
R216 B.n343 B.n58 585
R217 B.n342 B.n341 585
R218 B.n340 B.n59 585
R219 B.n339 B.n338 585
R220 B.n480 B.n479 585
R221 B.n481 B.n8 585
R222 B.n483 B.n482 585
R223 B.n484 B.n7 585
R224 B.n486 B.n485 585
R225 B.n487 B.n6 585
R226 B.n489 B.n488 585
R227 B.n490 B.n5 585
R228 B.n492 B.n491 585
R229 B.n493 B.n4 585
R230 B.n495 B.n494 585
R231 B.n496 B.n3 585
R232 B.n498 B.n497 585
R233 B.n499 B.n0 585
R234 B.n2 B.n1 585
R235 B.n133 B.n132 585
R236 B.n135 B.n134 585
R237 B.n136 B.n131 585
R238 B.n138 B.n137 585
R239 B.n139 B.n130 585
R240 B.n141 B.n140 585
R241 B.n142 B.n129 585
R242 B.n144 B.n143 585
R243 B.n145 B.n128 585
R244 B.n147 B.n146 585
R245 B.n148 B.n127 585
R246 B.n150 B.n149 585
R247 B.n151 B.n126 585
R248 B.n152 B.n151 535.745
R249 B.n294 B.n75 535.745
R250 B.n338 B.n337 535.745
R251 B.n480 B.n9 535.745
R252 B.n96 B.t10 391.433
R253 B.n38 B.t8 391.433
R254 B.n104 B.t1 391.433
R255 B.n30 B.t5 391.433
R256 B.n97 B.t11 377.276
R257 B.n39 B.t7 377.276
R258 B.n105 B.t2 377.276
R259 B.n31 B.t4 377.276
R260 B.n501 B.n500 256.663
R261 B.n500 B.n499 235.042
R262 B.n500 B.n2 235.042
R263 B.n152 B.n125 163.367
R264 B.n156 B.n125 163.367
R265 B.n157 B.n156 163.367
R266 B.n158 B.n157 163.367
R267 B.n158 B.n123 163.367
R268 B.n162 B.n123 163.367
R269 B.n163 B.n162 163.367
R270 B.n164 B.n163 163.367
R271 B.n164 B.n121 163.367
R272 B.n168 B.n121 163.367
R273 B.n169 B.n168 163.367
R274 B.n170 B.n169 163.367
R275 B.n170 B.n119 163.367
R276 B.n174 B.n119 163.367
R277 B.n175 B.n174 163.367
R278 B.n176 B.n175 163.367
R279 B.n176 B.n117 163.367
R280 B.n180 B.n117 163.367
R281 B.n181 B.n180 163.367
R282 B.n182 B.n181 163.367
R283 B.n182 B.n115 163.367
R284 B.n186 B.n115 163.367
R285 B.n187 B.n186 163.367
R286 B.n188 B.n187 163.367
R287 B.n188 B.n113 163.367
R288 B.n192 B.n113 163.367
R289 B.n193 B.n192 163.367
R290 B.n194 B.n193 163.367
R291 B.n194 B.n111 163.367
R292 B.n198 B.n111 163.367
R293 B.n199 B.n198 163.367
R294 B.n200 B.n199 163.367
R295 B.n200 B.n109 163.367
R296 B.n204 B.n109 163.367
R297 B.n205 B.n204 163.367
R298 B.n206 B.n205 163.367
R299 B.n206 B.n107 163.367
R300 B.n210 B.n107 163.367
R301 B.n211 B.n210 163.367
R302 B.n212 B.n211 163.367
R303 B.n212 B.n103 163.367
R304 B.n217 B.n103 163.367
R305 B.n218 B.n217 163.367
R306 B.n219 B.n218 163.367
R307 B.n219 B.n101 163.367
R308 B.n223 B.n101 163.367
R309 B.n224 B.n223 163.367
R310 B.n225 B.n224 163.367
R311 B.n225 B.n99 163.367
R312 B.n229 B.n99 163.367
R313 B.n230 B.n229 163.367
R314 B.n230 B.n95 163.367
R315 B.n234 B.n95 163.367
R316 B.n235 B.n234 163.367
R317 B.n236 B.n235 163.367
R318 B.n236 B.n93 163.367
R319 B.n240 B.n93 163.367
R320 B.n241 B.n240 163.367
R321 B.n242 B.n241 163.367
R322 B.n242 B.n91 163.367
R323 B.n246 B.n91 163.367
R324 B.n247 B.n246 163.367
R325 B.n248 B.n247 163.367
R326 B.n248 B.n89 163.367
R327 B.n252 B.n89 163.367
R328 B.n253 B.n252 163.367
R329 B.n254 B.n253 163.367
R330 B.n254 B.n87 163.367
R331 B.n258 B.n87 163.367
R332 B.n259 B.n258 163.367
R333 B.n260 B.n259 163.367
R334 B.n260 B.n85 163.367
R335 B.n264 B.n85 163.367
R336 B.n265 B.n264 163.367
R337 B.n266 B.n265 163.367
R338 B.n266 B.n83 163.367
R339 B.n270 B.n83 163.367
R340 B.n271 B.n270 163.367
R341 B.n272 B.n271 163.367
R342 B.n272 B.n81 163.367
R343 B.n276 B.n81 163.367
R344 B.n277 B.n276 163.367
R345 B.n278 B.n277 163.367
R346 B.n278 B.n79 163.367
R347 B.n282 B.n79 163.367
R348 B.n283 B.n282 163.367
R349 B.n284 B.n283 163.367
R350 B.n284 B.n77 163.367
R351 B.n288 B.n77 163.367
R352 B.n289 B.n288 163.367
R353 B.n290 B.n289 163.367
R354 B.n290 B.n75 163.367
R355 B.n337 B.n336 163.367
R356 B.n336 B.n61 163.367
R357 B.n332 B.n61 163.367
R358 B.n332 B.n331 163.367
R359 B.n331 B.n330 163.367
R360 B.n330 B.n63 163.367
R361 B.n326 B.n63 163.367
R362 B.n326 B.n325 163.367
R363 B.n325 B.n324 163.367
R364 B.n324 B.n65 163.367
R365 B.n320 B.n65 163.367
R366 B.n320 B.n319 163.367
R367 B.n319 B.n318 163.367
R368 B.n318 B.n67 163.367
R369 B.n314 B.n67 163.367
R370 B.n314 B.n313 163.367
R371 B.n313 B.n312 163.367
R372 B.n312 B.n69 163.367
R373 B.n308 B.n69 163.367
R374 B.n308 B.n307 163.367
R375 B.n307 B.n306 163.367
R376 B.n306 B.n71 163.367
R377 B.n302 B.n71 163.367
R378 B.n302 B.n301 163.367
R379 B.n301 B.n300 163.367
R380 B.n300 B.n73 163.367
R381 B.n296 B.n73 163.367
R382 B.n296 B.n295 163.367
R383 B.n295 B.n294 163.367
R384 B.n476 B.n9 163.367
R385 B.n476 B.n475 163.367
R386 B.n475 B.n474 163.367
R387 B.n474 B.n11 163.367
R388 B.n470 B.n11 163.367
R389 B.n470 B.n469 163.367
R390 B.n469 B.n468 163.367
R391 B.n468 B.n13 163.367
R392 B.n464 B.n13 163.367
R393 B.n464 B.n463 163.367
R394 B.n463 B.n462 163.367
R395 B.n462 B.n15 163.367
R396 B.n458 B.n15 163.367
R397 B.n458 B.n457 163.367
R398 B.n457 B.n456 163.367
R399 B.n456 B.n17 163.367
R400 B.n452 B.n17 163.367
R401 B.n452 B.n451 163.367
R402 B.n451 B.n450 163.367
R403 B.n450 B.n19 163.367
R404 B.n446 B.n19 163.367
R405 B.n446 B.n445 163.367
R406 B.n445 B.n444 163.367
R407 B.n444 B.n21 163.367
R408 B.n440 B.n21 163.367
R409 B.n440 B.n439 163.367
R410 B.n439 B.n438 163.367
R411 B.n438 B.n23 163.367
R412 B.n434 B.n23 163.367
R413 B.n434 B.n433 163.367
R414 B.n433 B.n432 163.367
R415 B.n432 B.n25 163.367
R416 B.n428 B.n25 163.367
R417 B.n428 B.n427 163.367
R418 B.n427 B.n426 163.367
R419 B.n426 B.n27 163.367
R420 B.n422 B.n27 163.367
R421 B.n422 B.n421 163.367
R422 B.n421 B.n420 163.367
R423 B.n420 B.n29 163.367
R424 B.n416 B.n29 163.367
R425 B.n416 B.n415 163.367
R426 B.n415 B.n33 163.367
R427 B.n411 B.n33 163.367
R428 B.n411 B.n410 163.367
R429 B.n410 B.n409 163.367
R430 B.n409 B.n35 163.367
R431 B.n405 B.n35 163.367
R432 B.n405 B.n404 163.367
R433 B.n404 B.n403 163.367
R434 B.n403 B.n37 163.367
R435 B.n398 B.n37 163.367
R436 B.n398 B.n397 163.367
R437 B.n397 B.n396 163.367
R438 B.n396 B.n41 163.367
R439 B.n392 B.n41 163.367
R440 B.n392 B.n391 163.367
R441 B.n391 B.n390 163.367
R442 B.n390 B.n43 163.367
R443 B.n386 B.n43 163.367
R444 B.n386 B.n385 163.367
R445 B.n385 B.n384 163.367
R446 B.n384 B.n45 163.367
R447 B.n380 B.n45 163.367
R448 B.n380 B.n379 163.367
R449 B.n379 B.n378 163.367
R450 B.n378 B.n47 163.367
R451 B.n374 B.n47 163.367
R452 B.n374 B.n373 163.367
R453 B.n373 B.n372 163.367
R454 B.n372 B.n49 163.367
R455 B.n368 B.n49 163.367
R456 B.n368 B.n367 163.367
R457 B.n367 B.n366 163.367
R458 B.n366 B.n51 163.367
R459 B.n362 B.n51 163.367
R460 B.n362 B.n361 163.367
R461 B.n361 B.n360 163.367
R462 B.n360 B.n53 163.367
R463 B.n356 B.n53 163.367
R464 B.n356 B.n355 163.367
R465 B.n355 B.n354 163.367
R466 B.n354 B.n55 163.367
R467 B.n350 B.n55 163.367
R468 B.n350 B.n349 163.367
R469 B.n349 B.n348 163.367
R470 B.n348 B.n57 163.367
R471 B.n344 B.n57 163.367
R472 B.n344 B.n343 163.367
R473 B.n343 B.n342 163.367
R474 B.n342 B.n59 163.367
R475 B.n338 B.n59 163.367
R476 B.n481 B.n480 163.367
R477 B.n482 B.n481 163.367
R478 B.n482 B.n7 163.367
R479 B.n486 B.n7 163.367
R480 B.n487 B.n486 163.367
R481 B.n488 B.n487 163.367
R482 B.n488 B.n5 163.367
R483 B.n492 B.n5 163.367
R484 B.n493 B.n492 163.367
R485 B.n494 B.n493 163.367
R486 B.n494 B.n3 163.367
R487 B.n498 B.n3 163.367
R488 B.n499 B.n498 163.367
R489 B.n133 B.n2 163.367
R490 B.n134 B.n133 163.367
R491 B.n134 B.n131 163.367
R492 B.n138 B.n131 163.367
R493 B.n139 B.n138 163.367
R494 B.n140 B.n139 163.367
R495 B.n140 B.n129 163.367
R496 B.n144 B.n129 163.367
R497 B.n145 B.n144 163.367
R498 B.n146 B.n145 163.367
R499 B.n146 B.n127 163.367
R500 B.n150 B.n127 163.367
R501 B.n151 B.n150 163.367
R502 B.n215 B.n105 59.5399
R503 B.n98 B.n97 59.5399
R504 B.n401 B.n39 59.5399
R505 B.n32 B.n31 59.5399
R506 B.n479 B.n478 34.8103
R507 B.n339 B.n60 34.8103
R508 B.n293 B.n292 34.8103
R509 B.n153 B.n126 34.8103
R510 B B.n501 18.0485
R511 B.n105 B.n104 14.1581
R512 B.n97 B.n96 14.1581
R513 B.n39 B.n38 14.1581
R514 B.n31 B.n30 14.1581
R515 B.n479 B.n8 10.6151
R516 B.n483 B.n8 10.6151
R517 B.n484 B.n483 10.6151
R518 B.n485 B.n484 10.6151
R519 B.n485 B.n6 10.6151
R520 B.n489 B.n6 10.6151
R521 B.n490 B.n489 10.6151
R522 B.n491 B.n490 10.6151
R523 B.n491 B.n4 10.6151
R524 B.n495 B.n4 10.6151
R525 B.n496 B.n495 10.6151
R526 B.n497 B.n496 10.6151
R527 B.n497 B.n0 10.6151
R528 B.n478 B.n477 10.6151
R529 B.n477 B.n10 10.6151
R530 B.n473 B.n10 10.6151
R531 B.n473 B.n472 10.6151
R532 B.n472 B.n471 10.6151
R533 B.n471 B.n12 10.6151
R534 B.n467 B.n12 10.6151
R535 B.n467 B.n466 10.6151
R536 B.n466 B.n465 10.6151
R537 B.n465 B.n14 10.6151
R538 B.n461 B.n14 10.6151
R539 B.n461 B.n460 10.6151
R540 B.n460 B.n459 10.6151
R541 B.n459 B.n16 10.6151
R542 B.n455 B.n16 10.6151
R543 B.n455 B.n454 10.6151
R544 B.n454 B.n453 10.6151
R545 B.n453 B.n18 10.6151
R546 B.n449 B.n18 10.6151
R547 B.n449 B.n448 10.6151
R548 B.n448 B.n447 10.6151
R549 B.n447 B.n20 10.6151
R550 B.n443 B.n20 10.6151
R551 B.n443 B.n442 10.6151
R552 B.n442 B.n441 10.6151
R553 B.n441 B.n22 10.6151
R554 B.n437 B.n22 10.6151
R555 B.n437 B.n436 10.6151
R556 B.n436 B.n435 10.6151
R557 B.n435 B.n24 10.6151
R558 B.n431 B.n24 10.6151
R559 B.n431 B.n430 10.6151
R560 B.n430 B.n429 10.6151
R561 B.n429 B.n26 10.6151
R562 B.n425 B.n26 10.6151
R563 B.n425 B.n424 10.6151
R564 B.n424 B.n423 10.6151
R565 B.n423 B.n28 10.6151
R566 B.n419 B.n28 10.6151
R567 B.n419 B.n418 10.6151
R568 B.n418 B.n417 10.6151
R569 B.n414 B.n413 10.6151
R570 B.n413 B.n412 10.6151
R571 B.n412 B.n34 10.6151
R572 B.n408 B.n34 10.6151
R573 B.n408 B.n407 10.6151
R574 B.n407 B.n406 10.6151
R575 B.n406 B.n36 10.6151
R576 B.n402 B.n36 10.6151
R577 B.n400 B.n399 10.6151
R578 B.n399 B.n40 10.6151
R579 B.n395 B.n40 10.6151
R580 B.n395 B.n394 10.6151
R581 B.n394 B.n393 10.6151
R582 B.n393 B.n42 10.6151
R583 B.n389 B.n42 10.6151
R584 B.n389 B.n388 10.6151
R585 B.n388 B.n387 10.6151
R586 B.n387 B.n44 10.6151
R587 B.n383 B.n44 10.6151
R588 B.n383 B.n382 10.6151
R589 B.n382 B.n381 10.6151
R590 B.n381 B.n46 10.6151
R591 B.n377 B.n46 10.6151
R592 B.n377 B.n376 10.6151
R593 B.n376 B.n375 10.6151
R594 B.n375 B.n48 10.6151
R595 B.n371 B.n48 10.6151
R596 B.n371 B.n370 10.6151
R597 B.n370 B.n369 10.6151
R598 B.n369 B.n50 10.6151
R599 B.n365 B.n50 10.6151
R600 B.n365 B.n364 10.6151
R601 B.n364 B.n363 10.6151
R602 B.n363 B.n52 10.6151
R603 B.n359 B.n52 10.6151
R604 B.n359 B.n358 10.6151
R605 B.n358 B.n357 10.6151
R606 B.n357 B.n54 10.6151
R607 B.n353 B.n54 10.6151
R608 B.n353 B.n352 10.6151
R609 B.n352 B.n351 10.6151
R610 B.n351 B.n56 10.6151
R611 B.n347 B.n56 10.6151
R612 B.n347 B.n346 10.6151
R613 B.n346 B.n345 10.6151
R614 B.n345 B.n58 10.6151
R615 B.n341 B.n58 10.6151
R616 B.n341 B.n340 10.6151
R617 B.n340 B.n339 10.6151
R618 B.n335 B.n60 10.6151
R619 B.n335 B.n334 10.6151
R620 B.n334 B.n333 10.6151
R621 B.n333 B.n62 10.6151
R622 B.n329 B.n62 10.6151
R623 B.n329 B.n328 10.6151
R624 B.n328 B.n327 10.6151
R625 B.n327 B.n64 10.6151
R626 B.n323 B.n64 10.6151
R627 B.n323 B.n322 10.6151
R628 B.n322 B.n321 10.6151
R629 B.n321 B.n66 10.6151
R630 B.n317 B.n66 10.6151
R631 B.n317 B.n316 10.6151
R632 B.n316 B.n315 10.6151
R633 B.n315 B.n68 10.6151
R634 B.n311 B.n68 10.6151
R635 B.n311 B.n310 10.6151
R636 B.n310 B.n309 10.6151
R637 B.n309 B.n70 10.6151
R638 B.n305 B.n70 10.6151
R639 B.n305 B.n304 10.6151
R640 B.n304 B.n303 10.6151
R641 B.n303 B.n72 10.6151
R642 B.n299 B.n72 10.6151
R643 B.n299 B.n298 10.6151
R644 B.n298 B.n297 10.6151
R645 B.n297 B.n74 10.6151
R646 B.n293 B.n74 10.6151
R647 B.n132 B.n1 10.6151
R648 B.n135 B.n132 10.6151
R649 B.n136 B.n135 10.6151
R650 B.n137 B.n136 10.6151
R651 B.n137 B.n130 10.6151
R652 B.n141 B.n130 10.6151
R653 B.n142 B.n141 10.6151
R654 B.n143 B.n142 10.6151
R655 B.n143 B.n128 10.6151
R656 B.n147 B.n128 10.6151
R657 B.n148 B.n147 10.6151
R658 B.n149 B.n148 10.6151
R659 B.n149 B.n126 10.6151
R660 B.n154 B.n153 10.6151
R661 B.n155 B.n154 10.6151
R662 B.n155 B.n124 10.6151
R663 B.n159 B.n124 10.6151
R664 B.n160 B.n159 10.6151
R665 B.n161 B.n160 10.6151
R666 B.n161 B.n122 10.6151
R667 B.n165 B.n122 10.6151
R668 B.n166 B.n165 10.6151
R669 B.n167 B.n166 10.6151
R670 B.n167 B.n120 10.6151
R671 B.n171 B.n120 10.6151
R672 B.n172 B.n171 10.6151
R673 B.n173 B.n172 10.6151
R674 B.n173 B.n118 10.6151
R675 B.n177 B.n118 10.6151
R676 B.n178 B.n177 10.6151
R677 B.n179 B.n178 10.6151
R678 B.n179 B.n116 10.6151
R679 B.n183 B.n116 10.6151
R680 B.n184 B.n183 10.6151
R681 B.n185 B.n184 10.6151
R682 B.n185 B.n114 10.6151
R683 B.n189 B.n114 10.6151
R684 B.n190 B.n189 10.6151
R685 B.n191 B.n190 10.6151
R686 B.n191 B.n112 10.6151
R687 B.n195 B.n112 10.6151
R688 B.n196 B.n195 10.6151
R689 B.n197 B.n196 10.6151
R690 B.n197 B.n110 10.6151
R691 B.n201 B.n110 10.6151
R692 B.n202 B.n201 10.6151
R693 B.n203 B.n202 10.6151
R694 B.n203 B.n108 10.6151
R695 B.n207 B.n108 10.6151
R696 B.n208 B.n207 10.6151
R697 B.n209 B.n208 10.6151
R698 B.n209 B.n106 10.6151
R699 B.n213 B.n106 10.6151
R700 B.n214 B.n213 10.6151
R701 B.n216 B.n102 10.6151
R702 B.n220 B.n102 10.6151
R703 B.n221 B.n220 10.6151
R704 B.n222 B.n221 10.6151
R705 B.n222 B.n100 10.6151
R706 B.n226 B.n100 10.6151
R707 B.n227 B.n226 10.6151
R708 B.n228 B.n227 10.6151
R709 B.n232 B.n231 10.6151
R710 B.n233 B.n232 10.6151
R711 B.n233 B.n94 10.6151
R712 B.n237 B.n94 10.6151
R713 B.n238 B.n237 10.6151
R714 B.n239 B.n238 10.6151
R715 B.n239 B.n92 10.6151
R716 B.n243 B.n92 10.6151
R717 B.n244 B.n243 10.6151
R718 B.n245 B.n244 10.6151
R719 B.n245 B.n90 10.6151
R720 B.n249 B.n90 10.6151
R721 B.n250 B.n249 10.6151
R722 B.n251 B.n250 10.6151
R723 B.n251 B.n88 10.6151
R724 B.n255 B.n88 10.6151
R725 B.n256 B.n255 10.6151
R726 B.n257 B.n256 10.6151
R727 B.n257 B.n86 10.6151
R728 B.n261 B.n86 10.6151
R729 B.n262 B.n261 10.6151
R730 B.n263 B.n262 10.6151
R731 B.n263 B.n84 10.6151
R732 B.n267 B.n84 10.6151
R733 B.n268 B.n267 10.6151
R734 B.n269 B.n268 10.6151
R735 B.n269 B.n82 10.6151
R736 B.n273 B.n82 10.6151
R737 B.n274 B.n273 10.6151
R738 B.n275 B.n274 10.6151
R739 B.n275 B.n80 10.6151
R740 B.n279 B.n80 10.6151
R741 B.n280 B.n279 10.6151
R742 B.n281 B.n280 10.6151
R743 B.n281 B.n78 10.6151
R744 B.n285 B.n78 10.6151
R745 B.n286 B.n285 10.6151
R746 B.n287 B.n286 10.6151
R747 B.n287 B.n76 10.6151
R748 B.n291 B.n76 10.6151
R749 B.n292 B.n291 10.6151
R750 B.n501 B.n0 8.11757
R751 B.n501 B.n1 8.11757
R752 B.n414 B.n32 6.5566
R753 B.n402 B.n401 6.5566
R754 B.n216 B.n215 6.5566
R755 B.n228 B.n98 6.5566
R756 B.n417 B.n32 4.05904
R757 B.n401 B.n400 4.05904
R758 B.n215 B.n214 4.05904
R759 B.n231 B.n98 4.05904
R760 VP.n0 VP.t3 848.215
R761 VP.n0 VP.t2 848.191
R762 VP.n2 VP.t1 827.232
R763 VP.n3 VP.t0 827.232
R764 VP.n4 VP.n3 161.3
R765 VP.n2 VP.n1 161.3
R766 VP.n1 VP.n0 109.745
R767 VP.n3 VP.n2 48.2005
R768 VP.n4 VP.n1 0.189894
R769 VP VP.n4 0.0516364
R770 VTAIL.n522 VTAIL.n462 756.745
R771 VTAIL.n60 VTAIL.n0 756.745
R772 VTAIL.n126 VTAIL.n66 756.745
R773 VTAIL.n192 VTAIL.n132 756.745
R774 VTAIL.n456 VTAIL.n396 756.745
R775 VTAIL.n390 VTAIL.n330 756.745
R776 VTAIL.n324 VTAIL.n264 756.745
R777 VTAIL.n258 VTAIL.n198 756.745
R778 VTAIL.n482 VTAIL.n481 585
R779 VTAIL.n487 VTAIL.n486 585
R780 VTAIL.n489 VTAIL.n488 585
R781 VTAIL.n478 VTAIL.n477 585
R782 VTAIL.n495 VTAIL.n494 585
R783 VTAIL.n497 VTAIL.n496 585
R784 VTAIL.n474 VTAIL.n473 585
R785 VTAIL.n504 VTAIL.n503 585
R786 VTAIL.n505 VTAIL.n472 585
R787 VTAIL.n507 VTAIL.n506 585
R788 VTAIL.n470 VTAIL.n469 585
R789 VTAIL.n513 VTAIL.n512 585
R790 VTAIL.n515 VTAIL.n514 585
R791 VTAIL.n466 VTAIL.n465 585
R792 VTAIL.n521 VTAIL.n520 585
R793 VTAIL.n523 VTAIL.n522 585
R794 VTAIL.n20 VTAIL.n19 585
R795 VTAIL.n25 VTAIL.n24 585
R796 VTAIL.n27 VTAIL.n26 585
R797 VTAIL.n16 VTAIL.n15 585
R798 VTAIL.n33 VTAIL.n32 585
R799 VTAIL.n35 VTAIL.n34 585
R800 VTAIL.n12 VTAIL.n11 585
R801 VTAIL.n42 VTAIL.n41 585
R802 VTAIL.n43 VTAIL.n10 585
R803 VTAIL.n45 VTAIL.n44 585
R804 VTAIL.n8 VTAIL.n7 585
R805 VTAIL.n51 VTAIL.n50 585
R806 VTAIL.n53 VTAIL.n52 585
R807 VTAIL.n4 VTAIL.n3 585
R808 VTAIL.n59 VTAIL.n58 585
R809 VTAIL.n61 VTAIL.n60 585
R810 VTAIL.n86 VTAIL.n85 585
R811 VTAIL.n91 VTAIL.n90 585
R812 VTAIL.n93 VTAIL.n92 585
R813 VTAIL.n82 VTAIL.n81 585
R814 VTAIL.n99 VTAIL.n98 585
R815 VTAIL.n101 VTAIL.n100 585
R816 VTAIL.n78 VTAIL.n77 585
R817 VTAIL.n108 VTAIL.n107 585
R818 VTAIL.n109 VTAIL.n76 585
R819 VTAIL.n111 VTAIL.n110 585
R820 VTAIL.n74 VTAIL.n73 585
R821 VTAIL.n117 VTAIL.n116 585
R822 VTAIL.n119 VTAIL.n118 585
R823 VTAIL.n70 VTAIL.n69 585
R824 VTAIL.n125 VTAIL.n124 585
R825 VTAIL.n127 VTAIL.n126 585
R826 VTAIL.n152 VTAIL.n151 585
R827 VTAIL.n157 VTAIL.n156 585
R828 VTAIL.n159 VTAIL.n158 585
R829 VTAIL.n148 VTAIL.n147 585
R830 VTAIL.n165 VTAIL.n164 585
R831 VTAIL.n167 VTAIL.n166 585
R832 VTAIL.n144 VTAIL.n143 585
R833 VTAIL.n174 VTAIL.n173 585
R834 VTAIL.n175 VTAIL.n142 585
R835 VTAIL.n177 VTAIL.n176 585
R836 VTAIL.n140 VTAIL.n139 585
R837 VTAIL.n183 VTAIL.n182 585
R838 VTAIL.n185 VTAIL.n184 585
R839 VTAIL.n136 VTAIL.n135 585
R840 VTAIL.n191 VTAIL.n190 585
R841 VTAIL.n193 VTAIL.n192 585
R842 VTAIL.n457 VTAIL.n456 585
R843 VTAIL.n455 VTAIL.n454 585
R844 VTAIL.n400 VTAIL.n399 585
R845 VTAIL.n449 VTAIL.n448 585
R846 VTAIL.n447 VTAIL.n446 585
R847 VTAIL.n404 VTAIL.n403 585
R848 VTAIL.n441 VTAIL.n440 585
R849 VTAIL.n439 VTAIL.n406 585
R850 VTAIL.n438 VTAIL.n437 585
R851 VTAIL.n409 VTAIL.n407 585
R852 VTAIL.n432 VTAIL.n431 585
R853 VTAIL.n430 VTAIL.n429 585
R854 VTAIL.n413 VTAIL.n412 585
R855 VTAIL.n424 VTAIL.n423 585
R856 VTAIL.n422 VTAIL.n421 585
R857 VTAIL.n417 VTAIL.n416 585
R858 VTAIL.n391 VTAIL.n390 585
R859 VTAIL.n389 VTAIL.n388 585
R860 VTAIL.n334 VTAIL.n333 585
R861 VTAIL.n383 VTAIL.n382 585
R862 VTAIL.n381 VTAIL.n380 585
R863 VTAIL.n338 VTAIL.n337 585
R864 VTAIL.n375 VTAIL.n374 585
R865 VTAIL.n373 VTAIL.n340 585
R866 VTAIL.n372 VTAIL.n371 585
R867 VTAIL.n343 VTAIL.n341 585
R868 VTAIL.n366 VTAIL.n365 585
R869 VTAIL.n364 VTAIL.n363 585
R870 VTAIL.n347 VTAIL.n346 585
R871 VTAIL.n358 VTAIL.n357 585
R872 VTAIL.n356 VTAIL.n355 585
R873 VTAIL.n351 VTAIL.n350 585
R874 VTAIL.n325 VTAIL.n324 585
R875 VTAIL.n323 VTAIL.n322 585
R876 VTAIL.n268 VTAIL.n267 585
R877 VTAIL.n317 VTAIL.n316 585
R878 VTAIL.n315 VTAIL.n314 585
R879 VTAIL.n272 VTAIL.n271 585
R880 VTAIL.n309 VTAIL.n308 585
R881 VTAIL.n307 VTAIL.n274 585
R882 VTAIL.n306 VTAIL.n305 585
R883 VTAIL.n277 VTAIL.n275 585
R884 VTAIL.n300 VTAIL.n299 585
R885 VTAIL.n298 VTAIL.n297 585
R886 VTAIL.n281 VTAIL.n280 585
R887 VTAIL.n292 VTAIL.n291 585
R888 VTAIL.n290 VTAIL.n289 585
R889 VTAIL.n285 VTAIL.n284 585
R890 VTAIL.n259 VTAIL.n258 585
R891 VTAIL.n257 VTAIL.n256 585
R892 VTAIL.n202 VTAIL.n201 585
R893 VTAIL.n251 VTAIL.n250 585
R894 VTAIL.n249 VTAIL.n248 585
R895 VTAIL.n206 VTAIL.n205 585
R896 VTAIL.n243 VTAIL.n242 585
R897 VTAIL.n241 VTAIL.n208 585
R898 VTAIL.n240 VTAIL.n239 585
R899 VTAIL.n211 VTAIL.n209 585
R900 VTAIL.n234 VTAIL.n233 585
R901 VTAIL.n232 VTAIL.n231 585
R902 VTAIL.n215 VTAIL.n214 585
R903 VTAIL.n226 VTAIL.n225 585
R904 VTAIL.n224 VTAIL.n223 585
R905 VTAIL.n219 VTAIL.n218 585
R906 VTAIL.n483 VTAIL.t3 329.036
R907 VTAIL.n21 VTAIL.t2 329.036
R908 VTAIL.n87 VTAIL.t7 329.036
R909 VTAIL.n153 VTAIL.t6 329.036
R910 VTAIL.n418 VTAIL.t5 329.036
R911 VTAIL.n352 VTAIL.t4 329.036
R912 VTAIL.n286 VTAIL.t1 329.036
R913 VTAIL.n220 VTAIL.t0 329.036
R914 VTAIL.n487 VTAIL.n481 171.744
R915 VTAIL.n488 VTAIL.n487 171.744
R916 VTAIL.n488 VTAIL.n477 171.744
R917 VTAIL.n495 VTAIL.n477 171.744
R918 VTAIL.n496 VTAIL.n495 171.744
R919 VTAIL.n496 VTAIL.n473 171.744
R920 VTAIL.n504 VTAIL.n473 171.744
R921 VTAIL.n505 VTAIL.n504 171.744
R922 VTAIL.n506 VTAIL.n505 171.744
R923 VTAIL.n506 VTAIL.n469 171.744
R924 VTAIL.n513 VTAIL.n469 171.744
R925 VTAIL.n514 VTAIL.n513 171.744
R926 VTAIL.n514 VTAIL.n465 171.744
R927 VTAIL.n521 VTAIL.n465 171.744
R928 VTAIL.n522 VTAIL.n521 171.744
R929 VTAIL.n25 VTAIL.n19 171.744
R930 VTAIL.n26 VTAIL.n25 171.744
R931 VTAIL.n26 VTAIL.n15 171.744
R932 VTAIL.n33 VTAIL.n15 171.744
R933 VTAIL.n34 VTAIL.n33 171.744
R934 VTAIL.n34 VTAIL.n11 171.744
R935 VTAIL.n42 VTAIL.n11 171.744
R936 VTAIL.n43 VTAIL.n42 171.744
R937 VTAIL.n44 VTAIL.n43 171.744
R938 VTAIL.n44 VTAIL.n7 171.744
R939 VTAIL.n51 VTAIL.n7 171.744
R940 VTAIL.n52 VTAIL.n51 171.744
R941 VTAIL.n52 VTAIL.n3 171.744
R942 VTAIL.n59 VTAIL.n3 171.744
R943 VTAIL.n60 VTAIL.n59 171.744
R944 VTAIL.n91 VTAIL.n85 171.744
R945 VTAIL.n92 VTAIL.n91 171.744
R946 VTAIL.n92 VTAIL.n81 171.744
R947 VTAIL.n99 VTAIL.n81 171.744
R948 VTAIL.n100 VTAIL.n99 171.744
R949 VTAIL.n100 VTAIL.n77 171.744
R950 VTAIL.n108 VTAIL.n77 171.744
R951 VTAIL.n109 VTAIL.n108 171.744
R952 VTAIL.n110 VTAIL.n109 171.744
R953 VTAIL.n110 VTAIL.n73 171.744
R954 VTAIL.n117 VTAIL.n73 171.744
R955 VTAIL.n118 VTAIL.n117 171.744
R956 VTAIL.n118 VTAIL.n69 171.744
R957 VTAIL.n125 VTAIL.n69 171.744
R958 VTAIL.n126 VTAIL.n125 171.744
R959 VTAIL.n157 VTAIL.n151 171.744
R960 VTAIL.n158 VTAIL.n157 171.744
R961 VTAIL.n158 VTAIL.n147 171.744
R962 VTAIL.n165 VTAIL.n147 171.744
R963 VTAIL.n166 VTAIL.n165 171.744
R964 VTAIL.n166 VTAIL.n143 171.744
R965 VTAIL.n174 VTAIL.n143 171.744
R966 VTAIL.n175 VTAIL.n174 171.744
R967 VTAIL.n176 VTAIL.n175 171.744
R968 VTAIL.n176 VTAIL.n139 171.744
R969 VTAIL.n183 VTAIL.n139 171.744
R970 VTAIL.n184 VTAIL.n183 171.744
R971 VTAIL.n184 VTAIL.n135 171.744
R972 VTAIL.n191 VTAIL.n135 171.744
R973 VTAIL.n192 VTAIL.n191 171.744
R974 VTAIL.n456 VTAIL.n455 171.744
R975 VTAIL.n455 VTAIL.n399 171.744
R976 VTAIL.n448 VTAIL.n399 171.744
R977 VTAIL.n448 VTAIL.n447 171.744
R978 VTAIL.n447 VTAIL.n403 171.744
R979 VTAIL.n440 VTAIL.n403 171.744
R980 VTAIL.n440 VTAIL.n439 171.744
R981 VTAIL.n439 VTAIL.n438 171.744
R982 VTAIL.n438 VTAIL.n407 171.744
R983 VTAIL.n431 VTAIL.n407 171.744
R984 VTAIL.n431 VTAIL.n430 171.744
R985 VTAIL.n430 VTAIL.n412 171.744
R986 VTAIL.n423 VTAIL.n412 171.744
R987 VTAIL.n423 VTAIL.n422 171.744
R988 VTAIL.n422 VTAIL.n416 171.744
R989 VTAIL.n390 VTAIL.n389 171.744
R990 VTAIL.n389 VTAIL.n333 171.744
R991 VTAIL.n382 VTAIL.n333 171.744
R992 VTAIL.n382 VTAIL.n381 171.744
R993 VTAIL.n381 VTAIL.n337 171.744
R994 VTAIL.n374 VTAIL.n337 171.744
R995 VTAIL.n374 VTAIL.n373 171.744
R996 VTAIL.n373 VTAIL.n372 171.744
R997 VTAIL.n372 VTAIL.n341 171.744
R998 VTAIL.n365 VTAIL.n341 171.744
R999 VTAIL.n365 VTAIL.n364 171.744
R1000 VTAIL.n364 VTAIL.n346 171.744
R1001 VTAIL.n357 VTAIL.n346 171.744
R1002 VTAIL.n357 VTAIL.n356 171.744
R1003 VTAIL.n356 VTAIL.n350 171.744
R1004 VTAIL.n324 VTAIL.n323 171.744
R1005 VTAIL.n323 VTAIL.n267 171.744
R1006 VTAIL.n316 VTAIL.n267 171.744
R1007 VTAIL.n316 VTAIL.n315 171.744
R1008 VTAIL.n315 VTAIL.n271 171.744
R1009 VTAIL.n308 VTAIL.n271 171.744
R1010 VTAIL.n308 VTAIL.n307 171.744
R1011 VTAIL.n307 VTAIL.n306 171.744
R1012 VTAIL.n306 VTAIL.n275 171.744
R1013 VTAIL.n299 VTAIL.n275 171.744
R1014 VTAIL.n299 VTAIL.n298 171.744
R1015 VTAIL.n298 VTAIL.n280 171.744
R1016 VTAIL.n291 VTAIL.n280 171.744
R1017 VTAIL.n291 VTAIL.n290 171.744
R1018 VTAIL.n290 VTAIL.n284 171.744
R1019 VTAIL.n258 VTAIL.n257 171.744
R1020 VTAIL.n257 VTAIL.n201 171.744
R1021 VTAIL.n250 VTAIL.n201 171.744
R1022 VTAIL.n250 VTAIL.n249 171.744
R1023 VTAIL.n249 VTAIL.n205 171.744
R1024 VTAIL.n242 VTAIL.n205 171.744
R1025 VTAIL.n242 VTAIL.n241 171.744
R1026 VTAIL.n241 VTAIL.n240 171.744
R1027 VTAIL.n240 VTAIL.n209 171.744
R1028 VTAIL.n233 VTAIL.n209 171.744
R1029 VTAIL.n233 VTAIL.n232 171.744
R1030 VTAIL.n232 VTAIL.n214 171.744
R1031 VTAIL.n225 VTAIL.n214 171.744
R1032 VTAIL.n225 VTAIL.n224 171.744
R1033 VTAIL.n224 VTAIL.n218 171.744
R1034 VTAIL.t3 VTAIL.n481 85.8723
R1035 VTAIL.t2 VTAIL.n19 85.8723
R1036 VTAIL.t7 VTAIL.n85 85.8723
R1037 VTAIL.t6 VTAIL.n151 85.8723
R1038 VTAIL.t5 VTAIL.n416 85.8723
R1039 VTAIL.t4 VTAIL.n350 85.8723
R1040 VTAIL.t1 VTAIL.n284 85.8723
R1041 VTAIL.t0 VTAIL.n218 85.8723
R1042 VTAIL.n527 VTAIL.n526 31.6035
R1043 VTAIL.n65 VTAIL.n64 31.6035
R1044 VTAIL.n131 VTAIL.n130 31.6035
R1045 VTAIL.n197 VTAIL.n196 31.6035
R1046 VTAIL.n461 VTAIL.n460 31.6035
R1047 VTAIL.n395 VTAIL.n394 31.6035
R1048 VTAIL.n329 VTAIL.n328 31.6035
R1049 VTAIL.n263 VTAIL.n262 31.6035
R1050 VTAIL.n527 VTAIL.n461 23.4186
R1051 VTAIL.n263 VTAIL.n197 23.4186
R1052 VTAIL.n507 VTAIL.n472 13.1884
R1053 VTAIL.n45 VTAIL.n10 13.1884
R1054 VTAIL.n111 VTAIL.n76 13.1884
R1055 VTAIL.n177 VTAIL.n142 13.1884
R1056 VTAIL.n441 VTAIL.n406 13.1884
R1057 VTAIL.n375 VTAIL.n340 13.1884
R1058 VTAIL.n309 VTAIL.n274 13.1884
R1059 VTAIL.n243 VTAIL.n208 13.1884
R1060 VTAIL.n503 VTAIL.n502 12.8005
R1061 VTAIL.n508 VTAIL.n470 12.8005
R1062 VTAIL.n41 VTAIL.n40 12.8005
R1063 VTAIL.n46 VTAIL.n8 12.8005
R1064 VTAIL.n107 VTAIL.n106 12.8005
R1065 VTAIL.n112 VTAIL.n74 12.8005
R1066 VTAIL.n173 VTAIL.n172 12.8005
R1067 VTAIL.n178 VTAIL.n140 12.8005
R1068 VTAIL.n442 VTAIL.n404 12.8005
R1069 VTAIL.n437 VTAIL.n408 12.8005
R1070 VTAIL.n376 VTAIL.n338 12.8005
R1071 VTAIL.n371 VTAIL.n342 12.8005
R1072 VTAIL.n310 VTAIL.n272 12.8005
R1073 VTAIL.n305 VTAIL.n276 12.8005
R1074 VTAIL.n244 VTAIL.n206 12.8005
R1075 VTAIL.n239 VTAIL.n210 12.8005
R1076 VTAIL.n501 VTAIL.n474 12.0247
R1077 VTAIL.n512 VTAIL.n511 12.0247
R1078 VTAIL.n39 VTAIL.n12 12.0247
R1079 VTAIL.n50 VTAIL.n49 12.0247
R1080 VTAIL.n105 VTAIL.n78 12.0247
R1081 VTAIL.n116 VTAIL.n115 12.0247
R1082 VTAIL.n171 VTAIL.n144 12.0247
R1083 VTAIL.n182 VTAIL.n181 12.0247
R1084 VTAIL.n446 VTAIL.n445 12.0247
R1085 VTAIL.n436 VTAIL.n409 12.0247
R1086 VTAIL.n380 VTAIL.n379 12.0247
R1087 VTAIL.n370 VTAIL.n343 12.0247
R1088 VTAIL.n314 VTAIL.n313 12.0247
R1089 VTAIL.n304 VTAIL.n277 12.0247
R1090 VTAIL.n248 VTAIL.n247 12.0247
R1091 VTAIL.n238 VTAIL.n211 12.0247
R1092 VTAIL.n498 VTAIL.n497 11.249
R1093 VTAIL.n515 VTAIL.n468 11.249
R1094 VTAIL.n36 VTAIL.n35 11.249
R1095 VTAIL.n53 VTAIL.n6 11.249
R1096 VTAIL.n102 VTAIL.n101 11.249
R1097 VTAIL.n119 VTAIL.n72 11.249
R1098 VTAIL.n168 VTAIL.n167 11.249
R1099 VTAIL.n185 VTAIL.n138 11.249
R1100 VTAIL.n449 VTAIL.n402 11.249
R1101 VTAIL.n433 VTAIL.n432 11.249
R1102 VTAIL.n383 VTAIL.n336 11.249
R1103 VTAIL.n367 VTAIL.n366 11.249
R1104 VTAIL.n317 VTAIL.n270 11.249
R1105 VTAIL.n301 VTAIL.n300 11.249
R1106 VTAIL.n251 VTAIL.n204 11.249
R1107 VTAIL.n235 VTAIL.n234 11.249
R1108 VTAIL.n483 VTAIL.n482 10.7239
R1109 VTAIL.n21 VTAIL.n20 10.7239
R1110 VTAIL.n87 VTAIL.n86 10.7239
R1111 VTAIL.n153 VTAIL.n152 10.7239
R1112 VTAIL.n418 VTAIL.n417 10.7239
R1113 VTAIL.n352 VTAIL.n351 10.7239
R1114 VTAIL.n286 VTAIL.n285 10.7239
R1115 VTAIL.n220 VTAIL.n219 10.7239
R1116 VTAIL.n494 VTAIL.n476 10.4732
R1117 VTAIL.n516 VTAIL.n466 10.4732
R1118 VTAIL.n32 VTAIL.n14 10.4732
R1119 VTAIL.n54 VTAIL.n4 10.4732
R1120 VTAIL.n98 VTAIL.n80 10.4732
R1121 VTAIL.n120 VTAIL.n70 10.4732
R1122 VTAIL.n164 VTAIL.n146 10.4732
R1123 VTAIL.n186 VTAIL.n136 10.4732
R1124 VTAIL.n450 VTAIL.n400 10.4732
R1125 VTAIL.n429 VTAIL.n411 10.4732
R1126 VTAIL.n384 VTAIL.n334 10.4732
R1127 VTAIL.n363 VTAIL.n345 10.4732
R1128 VTAIL.n318 VTAIL.n268 10.4732
R1129 VTAIL.n297 VTAIL.n279 10.4732
R1130 VTAIL.n252 VTAIL.n202 10.4732
R1131 VTAIL.n231 VTAIL.n213 10.4732
R1132 VTAIL.n493 VTAIL.n478 9.69747
R1133 VTAIL.n520 VTAIL.n519 9.69747
R1134 VTAIL.n31 VTAIL.n16 9.69747
R1135 VTAIL.n58 VTAIL.n57 9.69747
R1136 VTAIL.n97 VTAIL.n82 9.69747
R1137 VTAIL.n124 VTAIL.n123 9.69747
R1138 VTAIL.n163 VTAIL.n148 9.69747
R1139 VTAIL.n190 VTAIL.n189 9.69747
R1140 VTAIL.n454 VTAIL.n453 9.69747
R1141 VTAIL.n428 VTAIL.n413 9.69747
R1142 VTAIL.n388 VTAIL.n387 9.69747
R1143 VTAIL.n362 VTAIL.n347 9.69747
R1144 VTAIL.n322 VTAIL.n321 9.69747
R1145 VTAIL.n296 VTAIL.n281 9.69747
R1146 VTAIL.n256 VTAIL.n255 9.69747
R1147 VTAIL.n230 VTAIL.n215 9.69747
R1148 VTAIL.n526 VTAIL.n525 9.45567
R1149 VTAIL.n64 VTAIL.n63 9.45567
R1150 VTAIL.n130 VTAIL.n129 9.45567
R1151 VTAIL.n196 VTAIL.n195 9.45567
R1152 VTAIL.n460 VTAIL.n459 9.45567
R1153 VTAIL.n394 VTAIL.n393 9.45567
R1154 VTAIL.n328 VTAIL.n327 9.45567
R1155 VTAIL.n262 VTAIL.n261 9.45567
R1156 VTAIL.n525 VTAIL.n524 9.3005
R1157 VTAIL.n464 VTAIL.n463 9.3005
R1158 VTAIL.n519 VTAIL.n518 9.3005
R1159 VTAIL.n517 VTAIL.n516 9.3005
R1160 VTAIL.n468 VTAIL.n467 9.3005
R1161 VTAIL.n511 VTAIL.n510 9.3005
R1162 VTAIL.n509 VTAIL.n508 9.3005
R1163 VTAIL.n485 VTAIL.n484 9.3005
R1164 VTAIL.n480 VTAIL.n479 9.3005
R1165 VTAIL.n491 VTAIL.n490 9.3005
R1166 VTAIL.n493 VTAIL.n492 9.3005
R1167 VTAIL.n476 VTAIL.n475 9.3005
R1168 VTAIL.n499 VTAIL.n498 9.3005
R1169 VTAIL.n501 VTAIL.n500 9.3005
R1170 VTAIL.n502 VTAIL.n471 9.3005
R1171 VTAIL.n63 VTAIL.n62 9.3005
R1172 VTAIL.n2 VTAIL.n1 9.3005
R1173 VTAIL.n57 VTAIL.n56 9.3005
R1174 VTAIL.n55 VTAIL.n54 9.3005
R1175 VTAIL.n6 VTAIL.n5 9.3005
R1176 VTAIL.n49 VTAIL.n48 9.3005
R1177 VTAIL.n47 VTAIL.n46 9.3005
R1178 VTAIL.n23 VTAIL.n22 9.3005
R1179 VTAIL.n18 VTAIL.n17 9.3005
R1180 VTAIL.n29 VTAIL.n28 9.3005
R1181 VTAIL.n31 VTAIL.n30 9.3005
R1182 VTAIL.n14 VTAIL.n13 9.3005
R1183 VTAIL.n37 VTAIL.n36 9.3005
R1184 VTAIL.n39 VTAIL.n38 9.3005
R1185 VTAIL.n40 VTAIL.n9 9.3005
R1186 VTAIL.n129 VTAIL.n128 9.3005
R1187 VTAIL.n68 VTAIL.n67 9.3005
R1188 VTAIL.n123 VTAIL.n122 9.3005
R1189 VTAIL.n121 VTAIL.n120 9.3005
R1190 VTAIL.n72 VTAIL.n71 9.3005
R1191 VTAIL.n115 VTAIL.n114 9.3005
R1192 VTAIL.n113 VTAIL.n112 9.3005
R1193 VTAIL.n89 VTAIL.n88 9.3005
R1194 VTAIL.n84 VTAIL.n83 9.3005
R1195 VTAIL.n95 VTAIL.n94 9.3005
R1196 VTAIL.n97 VTAIL.n96 9.3005
R1197 VTAIL.n80 VTAIL.n79 9.3005
R1198 VTAIL.n103 VTAIL.n102 9.3005
R1199 VTAIL.n105 VTAIL.n104 9.3005
R1200 VTAIL.n106 VTAIL.n75 9.3005
R1201 VTAIL.n195 VTAIL.n194 9.3005
R1202 VTAIL.n134 VTAIL.n133 9.3005
R1203 VTAIL.n189 VTAIL.n188 9.3005
R1204 VTAIL.n187 VTAIL.n186 9.3005
R1205 VTAIL.n138 VTAIL.n137 9.3005
R1206 VTAIL.n181 VTAIL.n180 9.3005
R1207 VTAIL.n179 VTAIL.n178 9.3005
R1208 VTAIL.n155 VTAIL.n154 9.3005
R1209 VTAIL.n150 VTAIL.n149 9.3005
R1210 VTAIL.n161 VTAIL.n160 9.3005
R1211 VTAIL.n163 VTAIL.n162 9.3005
R1212 VTAIL.n146 VTAIL.n145 9.3005
R1213 VTAIL.n169 VTAIL.n168 9.3005
R1214 VTAIL.n171 VTAIL.n170 9.3005
R1215 VTAIL.n172 VTAIL.n141 9.3005
R1216 VTAIL.n420 VTAIL.n419 9.3005
R1217 VTAIL.n415 VTAIL.n414 9.3005
R1218 VTAIL.n426 VTAIL.n425 9.3005
R1219 VTAIL.n428 VTAIL.n427 9.3005
R1220 VTAIL.n411 VTAIL.n410 9.3005
R1221 VTAIL.n434 VTAIL.n433 9.3005
R1222 VTAIL.n436 VTAIL.n435 9.3005
R1223 VTAIL.n408 VTAIL.n405 9.3005
R1224 VTAIL.n459 VTAIL.n458 9.3005
R1225 VTAIL.n398 VTAIL.n397 9.3005
R1226 VTAIL.n453 VTAIL.n452 9.3005
R1227 VTAIL.n451 VTAIL.n450 9.3005
R1228 VTAIL.n402 VTAIL.n401 9.3005
R1229 VTAIL.n445 VTAIL.n444 9.3005
R1230 VTAIL.n443 VTAIL.n442 9.3005
R1231 VTAIL.n354 VTAIL.n353 9.3005
R1232 VTAIL.n349 VTAIL.n348 9.3005
R1233 VTAIL.n360 VTAIL.n359 9.3005
R1234 VTAIL.n362 VTAIL.n361 9.3005
R1235 VTAIL.n345 VTAIL.n344 9.3005
R1236 VTAIL.n368 VTAIL.n367 9.3005
R1237 VTAIL.n370 VTAIL.n369 9.3005
R1238 VTAIL.n342 VTAIL.n339 9.3005
R1239 VTAIL.n393 VTAIL.n392 9.3005
R1240 VTAIL.n332 VTAIL.n331 9.3005
R1241 VTAIL.n387 VTAIL.n386 9.3005
R1242 VTAIL.n385 VTAIL.n384 9.3005
R1243 VTAIL.n336 VTAIL.n335 9.3005
R1244 VTAIL.n379 VTAIL.n378 9.3005
R1245 VTAIL.n377 VTAIL.n376 9.3005
R1246 VTAIL.n288 VTAIL.n287 9.3005
R1247 VTAIL.n283 VTAIL.n282 9.3005
R1248 VTAIL.n294 VTAIL.n293 9.3005
R1249 VTAIL.n296 VTAIL.n295 9.3005
R1250 VTAIL.n279 VTAIL.n278 9.3005
R1251 VTAIL.n302 VTAIL.n301 9.3005
R1252 VTAIL.n304 VTAIL.n303 9.3005
R1253 VTAIL.n276 VTAIL.n273 9.3005
R1254 VTAIL.n327 VTAIL.n326 9.3005
R1255 VTAIL.n266 VTAIL.n265 9.3005
R1256 VTAIL.n321 VTAIL.n320 9.3005
R1257 VTAIL.n319 VTAIL.n318 9.3005
R1258 VTAIL.n270 VTAIL.n269 9.3005
R1259 VTAIL.n313 VTAIL.n312 9.3005
R1260 VTAIL.n311 VTAIL.n310 9.3005
R1261 VTAIL.n222 VTAIL.n221 9.3005
R1262 VTAIL.n217 VTAIL.n216 9.3005
R1263 VTAIL.n228 VTAIL.n227 9.3005
R1264 VTAIL.n230 VTAIL.n229 9.3005
R1265 VTAIL.n213 VTAIL.n212 9.3005
R1266 VTAIL.n236 VTAIL.n235 9.3005
R1267 VTAIL.n238 VTAIL.n237 9.3005
R1268 VTAIL.n210 VTAIL.n207 9.3005
R1269 VTAIL.n261 VTAIL.n260 9.3005
R1270 VTAIL.n200 VTAIL.n199 9.3005
R1271 VTAIL.n255 VTAIL.n254 9.3005
R1272 VTAIL.n253 VTAIL.n252 9.3005
R1273 VTAIL.n204 VTAIL.n203 9.3005
R1274 VTAIL.n247 VTAIL.n246 9.3005
R1275 VTAIL.n245 VTAIL.n244 9.3005
R1276 VTAIL.n490 VTAIL.n489 8.92171
R1277 VTAIL.n523 VTAIL.n464 8.92171
R1278 VTAIL.n28 VTAIL.n27 8.92171
R1279 VTAIL.n61 VTAIL.n2 8.92171
R1280 VTAIL.n94 VTAIL.n93 8.92171
R1281 VTAIL.n127 VTAIL.n68 8.92171
R1282 VTAIL.n160 VTAIL.n159 8.92171
R1283 VTAIL.n193 VTAIL.n134 8.92171
R1284 VTAIL.n457 VTAIL.n398 8.92171
R1285 VTAIL.n425 VTAIL.n424 8.92171
R1286 VTAIL.n391 VTAIL.n332 8.92171
R1287 VTAIL.n359 VTAIL.n358 8.92171
R1288 VTAIL.n325 VTAIL.n266 8.92171
R1289 VTAIL.n293 VTAIL.n292 8.92171
R1290 VTAIL.n259 VTAIL.n200 8.92171
R1291 VTAIL.n227 VTAIL.n226 8.92171
R1292 VTAIL.n486 VTAIL.n480 8.14595
R1293 VTAIL.n524 VTAIL.n462 8.14595
R1294 VTAIL.n24 VTAIL.n18 8.14595
R1295 VTAIL.n62 VTAIL.n0 8.14595
R1296 VTAIL.n90 VTAIL.n84 8.14595
R1297 VTAIL.n128 VTAIL.n66 8.14595
R1298 VTAIL.n156 VTAIL.n150 8.14595
R1299 VTAIL.n194 VTAIL.n132 8.14595
R1300 VTAIL.n458 VTAIL.n396 8.14595
R1301 VTAIL.n421 VTAIL.n415 8.14595
R1302 VTAIL.n392 VTAIL.n330 8.14595
R1303 VTAIL.n355 VTAIL.n349 8.14595
R1304 VTAIL.n326 VTAIL.n264 8.14595
R1305 VTAIL.n289 VTAIL.n283 8.14595
R1306 VTAIL.n260 VTAIL.n198 8.14595
R1307 VTAIL.n223 VTAIL.n217 8.14595
R1308 VTAIL.n485 VTAIL.n482 7.3702
R1309 VTAIL.n23 VTAIL.n20 7.3702
R1310 VTAIL.n89 VTAIL.n86 7.3702
R1311 VTAIL.n155 VTAIL.n152 7.3702
R1312 VTAIL.n420 VTAIL.n417 7.3702
R1313 VTAIL.n354 VTAIL.n351 7.3702
R1314 VTAIL.n288 VTAIL.n285 7.3702
R1315 VTAIL.n222 VTAIL.n219 7.3702
R1316 VTAIL.n486 VTAIL.n485 5.81868
R1317 VTAIL.n526 VTAIL.n462 5.81868
R1318 VTAIL.n24 VTAIL.n23 5.81868
R1319 VTAIL.n64 VTAIL.n0 5.81868
R1320 VTAIL.n90 VTAIL.n89 5.81868
R1321 VTAIL.n130 VTAIL.n66 5.81868
R1322 VTAIL.n156 VTAIL.n155 5.81868
R1323 VTAIL.n196 VTAIL.n132 5.81868
R1324 VTAIL.n460 VTAIL.n396 5.81868
R1325 VTAIL.n421 VTAIL.n420 5.81868
R1326 VTAIL.n394 VTAIL.n330 5.81868
R1327 VTAIL.n355 VTAIL.n354 5.81868
R1328 VTAIL.n328 VTAIL.n264 5.81868
R1329 VTAIL.n289 VTAIL.n288 5.81868
R1330 VTAIL.n262 VTAIL.n198 5.81868
R1331 VTAIL.n223 VTAIL.n222 5.81868
R1332 VTAIL.n489 VTAIL.n480 5.04292
R1333 VTAIL.n524 VTAIL.n523 5.04292
R1334 VTAIL.n27 VTAIL.n18 5.04292
R1335 VTAIL.n62 VTAIL.n61 5.04292
R1336 VTAIL.n93 VTAIL.n84 5.04292
R1337 VTAIL.n128 VTAIL.n127 5.04292
R1338 VTAIL.n159 VTAIL.n150 5.04292
R1339 VTAIL.n194 VTAIL.n193 5.04292
R1340 VTAIL.n458 VTAIL.n457 5.04292
R1341 VTAIL.n424 VTAIL.n415 5.04292
R1342 VTAIL.n392 VTAIL.n391 5.04292
R1343 VTAIL.n358 VTAIL.n349 5.04292
R1344 VTAIL.n326 VTAIL.n325 5.04292
R1345 VTAIL.n292 VTAIL.n283 5.04292
R1346 VTAIL.n260 VTAIL.n259 5.04292
R1347 VTAIL.n226 VTAIL.n217 5.04292
R1348 VTAIL.n490 VTAIL.n478 4.26717
R1349 VTAIL.n520 VTAIL.n464 4.26717
R1350 VTAIL.n28 VTAIL.n16 4.26717
R1351 VTAIL.n58 VTAIL.n2 4.26717
R1352 VTAIL.n94 VTAIL.n82 4.26717
R1353 VTAIL.n124 VTAIL.n68 4.26717
R1354 VTAIL.n160 VTAIL.n148 4.26717
R1355 VTAIL.n190 VTAIL.n134 4.26717
R1356 VTAIL.n454 VTAIL.n398 4.26717
R1357 VTAIL.n425 VTAIL.n413 4.26717
R1358 VTAIL.n388 VTAIL.n332 4.26717
R1359 VTAIL.n359 VTAIL.n347 4.26717
R1360 VTAIL.n322 VTAIL.n266 4.26717
R1361 VTAIL.n293 VTAIL.n281 4.26717
R1362 VTAIL.n256 VTAIL.n200 4.26717
R1363 VTAIL.n227 VTAIL.n215 4.26717
R1364 VTAIL.n494 VTAIL.n493 3.49141
R1365 VTAIL.n519 VTAIL.n466 3.49141
R1366 VTAIL.n32 VTAIL.n31 3.49141
R1367 VTAIL.n57 VTAIL.n4 3.49141
R1368 VTAIL.n98 VTAIL.n97 3.49141
R1369 VTAIL.n123 VTAIL.n70 3.49141
R1370 VTAIL.n164 VTAIL.n163 3.49141
R1371 VTAIL.n189 VTAIL.n136 3.49141
R1372 VTAIL.n453 VTAIL.n400 3.49141
R1373 VTAIL.n429 VTAIL.n428 3.49141
R1374 VTAIL.n387 VTAIL.n334 3.49141
R1375 VTAIL.n363 VTAIL.n362 3.49141
R1376 VTAIL.n321 VTAIL.n268 3.49141
R1377 VTAIL.n297 VTAIL.n296 3.49141
R1378 VTAIL.n255 VTAIL.n202 3.49141
R1379 VTAIL.n231 VTAIL.n230 3.49141
R1380 VTAIL.n497 VTAIL.n476 2.71565
R1381 VTAIL.n516 VTAIL.n515 2.71565
R1382 VTAIL.n35 VTAIL.n14 2.71565
R1383 VTAIL.n54 VTAIL.n53 2.71565
R1384 VTAIL.n101 VTAIL.n80 2.71565
R1385 VTAIL.n120 VTAIL.n119 2.71565
R1386 VTAIL.n167 VTAIL.n146 2.71565
R1387 VTAIL.n186 VTAIL.n185 2.71565
R1388 VTAIL.n450 VTAIL.n449 2.71565
R1389 VTAIL.n432 VTAIL.n411 2.71565
R1390 VTAIL.n384 VTAIL.n383 2.71565
R1391 VTAIL.n366 VTAIL.n345 2.71565
R1392 VTAIL.n318 VTAIL.n317 2.71565
R1393 VTAIL.n300 VTAIL.n279 2.71565
R1394 VTAIL.n252 VTAIL.n251 2.71565
R1395 VTAIL.n234 VTAIL.n213 2.71565
R1396 VTAIL.n419 VTAIL.n418 2.41282
R1397 VTAIL.n353 VTAIL.n352 2.41282
R1398 VTAIL.n287 VTAIL.n286 2.41282
R1399 VTAIL.n221 VTAIL.n220 2.41282
R1400 VTAIL.n484 VTAIL.n483 2.41282
R1401 VTAIL.n22 VTAIL.n21 2.41282
R1402 VTAIL.n88 VTAIL.n87 2.41282
R1403 VTAIL.n154 VTAIL.n153 2.41282
R1404 VTAIL.n498 VTAIL.n474 1.93989
R1405 VTAIL.n512 VTAIL.n468 1.93989
R1406 VTAIL.n36 VTAIL.n12 1.93989
R1407 VTAIL.n50 VTAIL.n6 1.93989
R1408 VTAIL.n102 VTAIL.n78 1.93989
R1409 VTAIL.n116 VTAIL.n72 1.93989
R1410 VTAIL.n168 VTAIL.n144 1.93989
R1411 VTAIL.n182 VTAIL.n138 1.93989
R1412 VTAIL.n446 VTAIL.n402 1.93989
R1413 VTAIL.n433 VTAIL.n409 1.93989
R1414 VTAIL.n380 VTAIL.n336 1.93989
R1415 VTAIL.n367 VTAIL.n343 1.93989
R1416 VTAIL.n314 VTAIL.n270 1.93989
R1417 VTAIL.n301 VTAIL.n277 1.93989
R1418 VTAIL.n248 VTAIL.n204 1.93989
R1419 VTAIL.n235 VTAIL.n211 1.93989
R1420 VTAIL.n503 VTAIL.n501 1.16414
R1421 VTAIL.n511 VTAIL.n470 1.16414
R1422 VTAIL.n41 VTAIL.n39 1.16414
R1423 VTAIL.n49 VTAIL.n8 1.16414
R1424 VTAIL.n107 VTAIL.n105 1.16414
R1425 VTAIL.n115 VTAIL.n74 1.16414
R1426 VTAIL.n173 VTAIL.n171 1.16414
R1427 VTAIL.n181 VTAIL.n140 1.16414
R1428 VTAIL.n445 VTAIL.n404 1.16414
R1429 VTAIL.n437 VTAIL.n436 1.16414
R1430 VTAIL.n379 VTAIL.n338 1.16414
R1431 VTAIL.n371 VTAIL.n370 1.16414
R1432 VTAIL.n313 VTAIL.n272 1.16414
R1433 VTAIL.n305 VTAIL.n304 1.16414
R1434 VTAIL.n247 VTAIL.n206 1.16414
R1435 VTAIL.n239 VTAIL.n238 1.16414
R1436 VTAIL.n329 VTAIL.n263 0.62981
R1437 VTAIL.n461 VTAIL.n395 0.62981
R1438 VTAIL.n197 VTAIL.n131 0.62981
R1439 VTAIL.n395 VTAIL.n329 0.470328
R1440 VTAIL.n131 VTAIL.n65 0.470328
R1441 VTAIL.n502 VTAIL.n472 0.388379
R1442 VTAIL.n508 VTAIL.n507 0.388379
R1443 VTAIL.n40 VTAIL.n10 0.388379
R1444 VTAIL.n46 VTAIL.n45 0.388379
R1445 VTAIL.n106 VTAIL.n76 0.388379
R1446 VTAIL.n112 VTAIL.n111 0.388379
R1447 VTAIL.n172 VTAIL.n142 0.388379
R1448 VTAIL.n178 VTAIL.n177 0.388379
R1449 VTAIL.n442 VTAIL.n441 0.388379
R1450 VTAIL.n408 VTAIL.n406 0.388379
R1451 VTAIL.n376 VTAIL.n375 0.388379
R1452 VTAIL.n342 VTAIL.n340 0.388379
R1453 VTAIL.n310 VTAIL.n309 0.388379
R1454 VTAIL.n276 VTAIL.n274 0.388379
R1455 VTAIL.n244 VTAIL.n243 0.388379
R1456 VTAIL.n210 VTAIL.n208 0.388379
R1457 VTAIL VTAIL.n65 0.373345
R1458 VTAIL VTAIL.n527 0.256966
R1459 VTAIL.n484 VTAIL.n479 0.155672
R1460 VTAIL.n491 VTAIL.n479 0.155672
R1461 VTAIL.n492 VTAIL.n491 0.155672
R1462 VTAIL.n492 VTAIL.n475 0.155672
R1463 VTAIL.n499 VTAIL.n475 0.155672
R1464 VTAIL.n500 VTAIL.n499 0.155672
R1465 VTAIL.n500 VTAIL.n471 0.155672
R1466 VTAIL.n509 VTAIL.n471 0.155672
R1467 VTAIL.n510 VTAIL.n509 0.155672
R1468 VTAIL.n510 VTAIL.n467 0.155672
R1469 VTAIL.n517 VTAIL.n467 0.155672
R1470 VTAIL.n518 VTAIL.n517 0.155672
R1471 VTAIL.n518 VTAIL.n463 0.155672
R1472 VTAIL.n525 VTAIL.n463 0.155672
R1473 VTAIL.n22 VTAIL.n17 0.155672
R1474 VTAIL.n29 VTAIL.n17 0.155672
R1475 VTAIL.n30 VTAIL.n29 0.155672
R1476 VTAIL.n30 VTAIL.n13 0.155672
R1477 VTAIL.n37 VTAIL.n13 0.155672
R1478 VTAIL.n38 VTAIL.n37 0.155672
R1479 VTAIL.n38 VTAIL.n9 0.155672
R1480 VTAIL.n47 VTAIL.n9 0.155672
R1481 VTAIL.n48 VTAIL.n47 0.155672
R1482 VTAIL.n48 VTAIL.n5 0.155672
R1483 VTAIL.n55 VTAIL.n5 0.155672
R1484 VTAIL.n56 VTAIL.n55 0.155672
R1485 VTAIL.n56 VTAIL.n1 0.155672
R1486 VTAIL.n63 VTAIL.n1 0.155672
R1487 VTAIL.n88 VTAIL.n83 0.155672
R1488 VTAIL.n95 VTAIL.n83 0.155672
R1489 VTAIL.n96 VTAIL.n95 0.155672
R1490 VTAIL.n96 VTAIL.n79 0.155672
R1491 VTAIL.n103 VTAIL.n79 0.155672
R1492 VTAIL.n104 VTAIL.n103 0.155672
R1493 VTAIL.n104 VTAIL.n75 0.155672
R1494 VTAIL.n113 VTAIL.n75 0.155672
R1495 VTAIL.n114 VTAIL.n113 0.155672
R1496 VTAIL.n114 VTAIL.n71 0.155672
R1497 VTAIL.n121 VTAIL.n71 0.155672
R1498 VTAIL.n122 VTAIL.n121 0.155672
R1499 VTAIL.n122 VTAIL.n67 0.155672
R1500 VTAIL.n129 VTAIL.n67 0.155672
R1501 VTAIL.n154 VTAIL.n149 0.155672
R1502 VTAIL.n161 VTAIL.n149 0.155672
R1503 VTAIL.n162 VTAIL.n161 0.155672
R1504 VTAIL.n162 VTAIL.n145 0.155672
R1505 VTAIL.n169 VTAIL.n145 0.155672
R1506 VTAIL.n170 VTAIL.n169 0.155672
R1507 VTAIL.n170 VTAIL.n141 0.155672
R1508 VTAIL.n179 VTAIL.n141 0.155672
R1509 VTAIL.n180 VTAIL.n179 0.155672
R1510 VTAIL.n180 VTAIL.n137 0.155672
R1511 VTAIL.n187 VTAIL.n137 0.155672
R1512 VTAIL.n188 VTAIL.n187 0.155672
R1513 VTAIL.n188 VTAIL.n133 0.155672
R1514 VTAIL.n195 VTAIL.n133 0.155672
R1515 VTAIL.n459 VTAIL.n397 0.155672
R1516 VTAIL.n452 VTAIL.n397 0.155672
R1517 VTAIL.n452 VTAIL.n451 0.155672
R1518 VTAIL.n451 VTAIL.n401 0.155672
R1519 VTAIL.n444 VTAIL.n401 0.155672
R1520 VTAIL.n444 VTAIL.n443 0.155672
R1521 VTAIL.n443 VTAIL.n405 0.155672
R1522 VTAIL.n435 VTAIL.n405 0.155672
R1523 VTAIL.n435 VTAIL.n434 0.155672
R1524 VTAIL.n434 VTAIL.n410 0.155672
R1525 VTAIL.n427 VTAIL.n410 0.155672
R1526 VTAIL.n427 VTAIL.n426 0.155672
R1527 VTAIL.n426 VTAIL.n414 0.155672
R1528 VTAIL.n419 VTAIL.n414 0.155672
R1529 VTAIL.n393 VTAIL.n331 0.155672
R1530 VTAIL.n386 VTAIL.n331 0.155672
R1531 VTAIL.n386 VTAIL.n385 0.155672
R1532 VTAIL.n385 VTAIL.n335 0.155672
R1533 VTAIL.n378 VTAIL.n335 0.155672
R1534 VTAIL.n378 VTAIL.n377 0.155672
R1535 VTAIL.n377 VTAIL.n339 0.155672
R1536 VTAIL.n369 VTAIL.n339 0.155672
R1537 VTAIL.n369 VTAIL.n368 0.155672
R1538 VTAIL.n368 VTAIL.n344 0.155672
R1539 VTAIL.n361 VTAIL.n344 0.155672
R1540 VTAIL.n361 VTAIL.n360 0.155672
R1541 VTAIL.n360 VTAIL.n348 0.155672
R1542 VTAIL.n353 VTAIL.n348 0.155672
R1543 VTAIL.n327 VTAIL.n265 0.155672
R1544 VTAIL.n320 VTAIL.n265 0.155672
R1545 VTAIL.n320 VTAIL.n319 0.155672
R1546 VTAIL.n319 VTAIL.n269 0.155672
R1547 VTAIL.n312 VTAIL.n269 0.155672
R1548 VTAIL.n312 VTAIL.n311 0.155672
R1549 VTAIL.n311 VTAIL.n273 0.155672
R1550 VTAIL.n303 VTAIL.n273 0.155672
R1551 VTAIL.n303 VTAIL.n302 0.155672
R1552 VTAIL.n302 VTAIL.n278 0.155672
R1553 VTAIL.n295 VTAIL.n278 0.155672
R1554 VTAIL.n295 VTAIL.n294 0.155672
R1555 VTAIL.n294 VTAIL.n282 0.155672
R1556 VTAIL.n287 VTAIL.n282 0.155672
R1557 VTAIL.n261 VTAIL.n199 0.155672
R1558 VTAIL.n254 VTAIL.n199 0.155672
R1559 VTAIL.n254 VTAIL.n253 0.155672
R1560 VTAIL.n253 VTAIL.n203 0.155672
R1561 VTAIL.n246 VTAIL.n203 0.155672
R1562 VTAIL.n246 VTAIL.n245 0.155672
R1563 VTAIL.n245 VTAIL.n207 0.155672
R1564 VTAIL.n237 VTAIL.n207 0.155672
R1565 VTAIL.n237 VTAIL.n236 0.155672
R1566 VTAIL.n236 VTAIL.n212 0.155672
R1567 VTAIL.n229 VTAIL.n212 0.155672
R1568 VTAIL.n229 VTAIL.n228 0.155672
R1569 VTAIL.n228 VTAIL.n216 0.155672
R1570 VTAIL.n221 VTAIL.n216 0.155672
R1571 VDD1 VDD1.n1 109.808
R1572 VDD1 VDD1.n0 73.3154
R1573 VDD1.n0 VDD1.t0 2.68909
R1574 VDD1.n0 VDD1.t1 2.68909
R1575 VDD1.n1 VDD1.t2 2.68909
R1576 VDD1.n1 VDD1.t3 2.68909
R1577 VN.n0 VN.t2 848.215
R1578 VN.n1 VN.t1 848.215
R1579 VN.n0 VN.t3 848.191
R1580 VN.n1 VN.t0 848.191
R1581 VN VN.n1 110.124
R1582 VN VN.n0 70.265
R1583 VDD2.n2 VDD2.n0 109.282
R1584 VDD2.n2 VDD2.n1 73.2572
R1585 VDD2.n1 VDD2.t3 2.68909
R1586 VDD2.n1 VDD2.t2 2.68909
R1587 VDD2.n0 VDD2.t1 2.68909
R1588 VDD2.n0 VDD2.t0 2.68909
R1589 VDD2 VDD2.n2 0.0586897
C0 VTAIL VDD2 8.51091f
C1 VTAIL B 3.61238f
C2 w_n1408_n3386# VN 1.98676f
C3 VP w_n1408_n3386# 2.1622f
C4 VDD1 w_n1408_n3386# 0.998938f
C5 VTAIL VN 1.93125f
C6 VTAIL VP 1.94536f
C7 VTAIL VDD1 8.47145f
C8 VDD2 B 0.892242f
C9 VTAIL w_n1408_n3386# 4.24969f
C10 VDD2 VN 2.41681f
C11 VN B 0.688444f
C12 VDD2 VP 0.254419f
C13 VDD1 VDD2 0.50175f
C14 VP B 0.96934f
C15 VDD1 B 0.874892f
C16 VP VN 4.62597f
C17 VDD1 VN 0.147115f
C18 VDD2 w_n1408_n3386# 1.00768f
C19 VDD1 VP 2.52393f
C20 w_n1408_n3386# B 6.56425f
C21 VDD2 VSUBS 0.643003f
C22 VDD1 VSUBS 5.228796f
C23 VTAIL VSUBS 0.771475f
C24 VN VSUBS 4.57095f
C25 VP VSUBS 1.136628f
C26 B VSUBS 2.370393f
C27 w_n1408_n3386# VSUBS 58.6798f
C28 VDD2.t1 VSUBS 0.295777f
C29 VDD2.t0 VSUBS 0.295777f
C30 VDD2.n0 VSUBS 3.00057f
C31 VDD2.t3 VSUBS 0.295777f
C32 VDD2.t2 VSUBS 0.295777f
C33 VDD2.n1 VSUBS 2.30778f
C34 VDD2.n2 VSUBS 4.3391f
C35 VN.t2 VSUBS 0.623008f
C36 VN.t3 VSUBS 0.622999f
C37 VN.n0 VSUBS 0.488966f
C38 VN.t1 VSUBS 0.623008f
C39 VN.t0 VSUBS 0.622999f
C40 VN.n1 VSUBS 1.12052f
C41 VDD1.t0 VSUBS 0.295392f
C42 VDD1.t1 VSUBS 0.295392f
C43 VDD1.n0 VSUBS 2.30531f
C44 VDD1.t2 VSUBS 0.295392f
C45 VDD1.t3 VSUBS 0.295392f
C46 VDD1.n1 VSUBS 3.02433f
C47 VTAIL.n0 VSUBS 0.023046f
C48 VTAIL.n1 VSUBS 0.021301f
C49 VTAIL.n2 VSUBS 0.011446f
C50 VTAIL.n3 VSUBS 0.027055f
C51 VTAIL.n4 VSUBS 0.01212f
C52 VTAIL.n5 VSUBS 0.021301f
C53 VTAIL.n6 VSUBS 0.011446f
C54 VTAIL.n7 VSUBS 0.027055f
C55 VTAIL.n8 VSUBS 0.01212f
C56 VTAIL.n9 VSUBS 0.021301f
C57 VTAIL.n10 VSUBS 0.011783f
C58 VTAIL.n11 VSUBS 0.027055f
C59 VTAIL.n12 VSUBS 0.01212f
C60 VTAIL.n13 VSUBS 0.021301f
C61 VTAIL.n14 VSUBS 0.011446f
C62 VTAIL.n15 VSUBS 0.027055f
C63 VTAIL.n16 VSUBS 0.01212f
C64 VTAIL.n17 VSUBS 0.021301f
C65 VTAIL.n18 VSUBS 0.011446f
C66 VTAIL.n19 VSUBS 0.020291f
C67 VTAIL.n20 VSUBS 0.020352f
C68 VTAIL.t2 VSUBS 0.058307f
C69 VTAIL.n21 VSUBS 0.168628f
C70 VTAIL.n22 VSUBS 1.05501f
C71 VTAIL.n23 VSUBS 0.011446f
C72 VTAIL.n24 VSUBS 0.01212f
C73 VTAIL.n25 VSUBS 0.027055f
C74 VTAIL.n26 VSUBS 0.027055f
C75 VTAIL.n27 VSUBS 0.01212f
C76 VTAIL.n28 VSUBS 0.011446f
C77 VTAIL.n29 VSUBS 0.021301f
C78 VTAIL.n30 VSUBS 0.021301f
C79 VTAIL.n31 VSUBS 0.011446f
C80 VTAIL.n32 VSUBS 0.01212f
C81 VTAIL.n33 VSUBS 0.027055f
C82 VTAIL.n34 VSUBS 0.027055f
C83 VTAIL.n35 VSUBS 0.01212f
C84 VTAIL.n36 VSUBS 0.011446f
C85 VTAIL.n37 VSUBS 0.021301f
C86 VTAIL.n38 VSUBS 0.021301f
C87 VTAIL.n39 VSUBS 0.011446f
C88 VTAIL.n40 VSUBS 0.011446f
C89 VTAIL.n41 VSUBS 0.01212f
C90 VTAIL.n42 VSUBS 0.027055f
C91 VTAIL.n43 VSUBS 0.027055f
C92 VTAIL.n44 VSUBS 0.027055f
C93 VTAIL.n45 VSUBS 0.011783f
C94 VTAIL.n46 VSUBS 0.011446f
C95 VTAIL.n47 VSUBS 0.021301f
C96 VTAIL.n48 VSUBS 0.021301f
C97 VTAIL.n49 VSUBS 0.011446f
C98 VTAIL.n50 VSUBS 0.01212f
C99 VTAIL.n51 VSUBS 0.027055f
C100 VTAIL.n52 VSUBS 0.027055f
C101 VTAIL.n53 VSUBS 0.01212f
C102 VTAIL.n54 VSUBS 0.011446f
C103 VTAIL.n55 VSUBS 0.021301f
C104 VTAIL.n56 VSUBS 0.021301f
C105 VTAIL.n57 VSUBS 0.011446f
C106 VTAIL.n58 VSUBS 0.01212f
C107 VTAIL.n59 VSUBS 0.027055f
C108 VTAIL.n60 VSUBS 0.064272f
C109 VTAIL.n61 VSUBS 0.01212f
C110 VTAIL.n62 VSUBS 0.011446f
C111 VTAIL.n63 VSUBS 0.048364f
C112 VTAIL.n64 VSUBS 0.03224f
C113 VTAIL.n65 VSUBS 0.07554f
C114 VTAIL.n66 VSUBS 0.023046f
C115 VTAIL.n67 VSUBS 0.021301f
C116 VTAIL.n68 VSUBS 0.011446f
C117 VTAIL.n69 VSUBS 0.027055f
C118 VTAIL.n70 VSUBS 0.01212f
C119 VTAIL.n71 VSUBS 0.021301f
C120 VTAIL.n72 VSUBS 0.011446f
C121 VTAIL.n73 VSUBS 0.027055f
C122 VTAIL.n74 VSUBS 0.01212f
C123 VTAIL.n75 VSUBS 0.021301f
C124 VTAIL.n76 VSUBS 0.011783f
C125 VTAIL.n77 VSUBS 0.027055f
C126 VTAIL.n78 VSUBS 0.01212f
C127 VTAIL.n79 VSUBS 0.021301f
C128 VTAIL.n80 VSUBS 0.011446f
C129 VTAIL.n81 VSUBS 0.027055f
C130 VTAIL.n82 VSUBS 0.01212f
C131 VTAIL.n83 VSUBS 0.021301f
C132 VTAIL.n84 VSUBS 0.011446f
C133 VTAIL.n85 VSUBS 0.020291f
C134 VTAIL.n86 VSUBS 0.020352f
C135 VTAIL.t7 VSUBS 0.058307f
C136 VTAIL.n87 VSUBS 0.168628f
C137 VTAIL.n88 VSUBS 1.05501f
C138 VTAIL.n89 VSUBS 0.011446f
C139 VTAIL.n90 VSUBS 0.01212f
C140 VTAIL.n91 VSUBS 0.027055f
C141 VTAIL.n92 VSUBS 0.027055f
C142 VTAIL.n93 VSUBS 0.01212f
C143 VTAIL.n94 VSUBS 0.011446f
C144 VTAIL.n95 VSUBS 0.021301f
C145 VTAIL.n96 VSUBS 0.021301f
C146 VTAIL.n97 VSUBS 0.011446f
C147 VTAIL.n98 VSUBS 0.01212f
C148 VTAIL.n99 VSUBS 0.027055f
C149 VTAIL.n100 VSUBS 0.027055f
C150 VTAIL.n101 VSUBS 0.01212f
C151 VTAIL.n102 VSUBS 0.011446f
C152 VTAIL.n103 VSUBS 0.021301f
C153 VTAIL.n104 VSUBS 0.021301f
C154 VTAIL.n105 VSUBS 0.011446f
C155 VTAIL.n106 VSUBS 0.011446f
C156 VTAIL.n107 VSUBS 0.01212f
C157 VTAIL.n108 VSUBS 0.027055f
C158 VTAIL.n109 VSUBS 0.027055f
C159 VTAIL.n110 VSUBS 0.027055f
C160 VTAIL.n111 VSUBS 0.011783f
C161 VTAIL.n112 VSUBS 0.011446f
C162 VTAIL.n113 VSUBS 0.021301f
C163 VTAIL.n114 VSUBS 0.021301f
C164 VTAIL.n115 VSUBS 0.011446f
C165 VTAIL.n116 VSUBS 0.01212f
C166 VTAIL.n117 VSUBS 0.027055f
C167 VTAIL.n118 VSUBS 0.027055f
C168 VTAIL.n119 VSUBS 0.01212f
C169 VTAIL.n120 VSUBS 0.011446f
C170 VTAIL.n121 VSUBS 0.021301f
C171 VTAIL.n122 VSUBS 0.021301f
C172 VTAIL.n123 VSUBS 0.011446f
C173 VTAIL.n124 VSUBS 0.01212f
C174 VTAIL.n125 VSUBS 0.027055f
C175 VTAIL.n126 VSUBS 0.064272f
C176 VTAIL.n127 VSUBS 0.01212f
C177 VTAIL.n128 VSUBS 0.011446f
C178 VTAIL.n129 VSUBS 0.048364f
C179 VTAIL.n130 VSUBS 0.03224f
C180 VTAIL.n131 VSUBS 0.093143f
C181 VTAIL.n132 VSUBS 0.023046f
C182 VTAIL.n133 VSUBS 0.021301f
C183 VTAIL.n134 VSUBS 0.011446f
C184 VTAIL.n135 VSUBS 0.027055f
C185 VTAIL.n136 VSUBS 0.01212f
C186 VTAIL.n137 VSUBS 0.021301f
C187 VTAIL.n138 VSUBS 0.011446f
C188 VTAIL.n139 VSUBS 0.027055f
C189 VTAIL.n140 VSUBS 0.01212f
C190 VTAIL.n141 VSUBS 0.021301f
C191 VTAIL.n142 VSUBS 0.011783f
C192 VTAIL.n143 VSUBS 0.027055f
C193 VTAIL.n144 VSUBS 0.01212f
C194 VTAIL.n145 VSUBS 0.021301f
C195 VTAIL.n146 VSUBS 0.011446f
C196 VTAIL.n147 VSUBS 0.027055f
C197 VTAIL.n148 VSUBS 0.01212f
C198 VTAIL.n149 VSUBS 0.021301f
C199 VTAIL.n150 VSUBS 0.011446f
C200 VTAIL.n151 VSUBS 0.020291f
C201 VTAIL.n152 VSUBS 0.020352f
C202 VTAIL.t6 VSUBS 0.058307f
C203 VTAIL.n153 VSUBS 0.168628f
C204 VTAIL.n154 VSUBS 1.05501f
C205 VTAIL.n155 VSUBS 0.011446f
C206 VTAIL.n156 VSUBS 0.01212f
C207 VTAIL.n157 VSUBS 0.027055f
C208 VTAIL.n158 VSUBS 0.027055f
C209 VTAIL.n159 VSUBS 0.01212f
C210 VTAIL.n160 VSUBS 0.011446f
C211 VTAIL.n161 VSUBS 0.021301f
C212 VTAIL.n162 VSUBS 0.021301f
C213 VTAIL.n163 VSUBS 0.011446f
C214 VTAIL.n164 VSUBS 0.01212f
C215 VTAIL.n165 VSUBS 0.027055f
C216 VTAIL.n166 VSUBS 0.027055f
C217 VTAIL.n167 VSUBS 0.01212f
C218 VTAIL.n168 VSUBS 0.011446f
C219 VTAIL.n169 VSUBS 0.021301f
C220 VTAIL.n170 VSUBS 0.021301f
C221 VTAIL.n171 VSUBS 0.011446f
C222 VTAIL.n172 VSUBS 0.011446f
C223 VTAIL.n173 VSUBS 0.01212f
C224 VTAIL.n174 VSUBS 0.027055f
C225 VTAIL.n175 VSUBS 0.027055f
C226 VTAIL.n176 VSUBS 0.027055f
C227 VTAIL.n177 VSUBS 0.011783f
C228 VTAIL.n178 VSUBS 0.011446f
C229 VTAIL.n179 VSUBS 0.021301f
C230 VTAIL.n180 VSUBS 0.021301f
C231 VTAIL.n181 VSUBS 0.011446f
C232 VTAIL.n182 VSUBS 0.01212f
C233 VTAIL.n183 VSUBS 0.027055f
C234 VTAIL.n184 VSUBS 0.027055f
C235 VTAIL.n185 VSUBS 0.01212f
C236 VTAIL.n186 VSUBS 0.011446f
C237 VTAIL.n187 VSUBS 0.021301f
C238 VTAIL.n188 VSUBS 0.021301f
C239 VTAIL.n189 VSUBS 0.011446f
C240 VTAIL.n190 VSUBS 0.01212f
C241 VTAIL.n191 VSUBS 0.027055f
C242 VTAIL.n192 VSUBS 0.064272f
C243 VTAIL.n193 VSUBS 0.01212f
C244 VTAIL.n194 VSUBS 0.011446f
C245 VTAIL.n195 VSUBS 0.048364f
C246 VTAIL.n196 VSUBS 0.03224f
C247 VTAIL.n197 VSUBS 1.10882f
C248 VTAIL.n198 VSUBS 0.023046f
C249 VTAIL.n199 VSUBS 0.021301f
C250 VTAIL.n200 VSUBS 0.011446f
C251 VTAIL.n201 VSUBS 0.027055f
C252 VTAIL.n202 VSUBS 0.01212f
C253 VTAIL.n203 VSUBS 0.021301f
C254 VTAIL.n204 VSUBS 0.011446f
C255 VTAIL.n205 VSUBS 0.027055f
C256 VTAIL.n206 VSUBS 0.01212f
C257 VTAIL.n207 VSUBS 0.021301f
C258 VTAIL.n208 VSUBS 0.011783f
C259 VTAIL.n209 VSUBS 0.027055f
C260 VTAIL.n210 VSUBS 0.011446f
C261 VTAIL.n211 VSUBS 0.01212f
C262 VTAIL.n212 VSUBS 0.021301f
C263 VTAIL.n213 VSUBS 0.011446f
C264 VTAIL.n214 VSUBS 0.027055f
C265 VTAIL.n215 VSUBS 0.01212f
C266 VTAIL.n216 VSUBS 0.021301f
C267 VTAIL.n217 VSUBS 0.011446f
C268 VTAIL.n218 VSUBS 0.020291f
C269 VTAIL.n219 VSUBS 0.020352f
C270 VTAIL.t0 VSUBS 0.058307f
C271 VTAIL.n220 VSUBS 0.168628f
C272 VTAIL.n221 VSUBS 1.05501f
C273 VTAIL.n222 VSUBS 0.011446f
C274 VTAIL.n223 VSUBS 0.01212f
C275 VTAIL.n224 VSUBS 0.027055f
C276 VTAIL.n225 VSUBS 0.027055f
C277 VTAIL.n226 VSUBS 0.01212f
C278 VTAIL.n227 VSUBS 0.011446f
C279 VTAIL.n228 VSUBS 0.021301f
C280 VTAIL.n229 VSUBS 0.021301f
C281 VTAIL.n230 VSUBS 0.011446f
C282 VTAIL.n231 VSUBS 0.01212f
C283 VTAIL.n232 VSUBS 0.027055f
C284 VTAIL.n233 VSUBS 0.027055f
C285 VTAIL.n234 VSUBS 0.01212f
C286 VTAIL.n235 VSUBS 0.011446f
C287 VTAIL.n236 VSUBS 0.021301f
C288 VTAIL.n237 VSUBS 0.021301f
C289 VTAIL.n238 VSUBS 0.011446f
C290 VTAIL.n239 VSUBS 0.01212f
C291 VTAIL.n240 VSUBS 0.027055f
C292 VTAIL.n241 VSUBS 0.027055f
C293 VTAIL.n242 VSUBS 0.027055f
C294 VTAIL.n243 VSUBS 0.011783f
C295 VTAIL.n244 VSUBS 0.011446f
C296 VTAIL.n245 VSUBS 0.021301f
C297 VTAIL.n246 VSUBS 0.021301f
C298 VTAIL.n247 VSUBS 0.011446f
C299 VTAIL.n248 VSUBS 0.01212f
C300 VTAIL.n249 VSUBS 0.027055f
C301 VTAIL.n250 VSUBS 0.027055f
C302 VTAIL.n251 VSUBS 0.01212f
C303 VTAIL.n252 VSUBS 0.011446f
C304 VTAIL.n253 VSUBS 0.021301f
C305 VTAIL.n254 VSUBS 0.021301f
C306 VTAIL.n255 VSUBS 0.011446f
C307 VTAIL.n256 VSUBS 0.01212f
C308 VTAIL.n257 VSUBS 0.027055f
C309 VTAIL.n258 VSUBS 0.064272f
C310 VTAIL.n259 VSUBS 0.01212f
C311 VTAIL.n260 VSUBS 0.011446f
C312 VTAIL.n261 VSUBS 0.048364f
C313 VTAIL.n262 VSUBS 0.03224f
C314 VTAIL.n263 VSUBS 1.10882f
C315 VTAIL.n264 VSUBS 0.023046f
C316 VTAIL.n265 VSUBS 0.021301f
C317 VTAIL.n266 VSUBS 0.011446f
C318 VTAIL.n267 VSUBS 0.027055f
C319 VTAIL.n268 VSUBS 0.01212f
C320 VTAIL.n269 VSUBS 0.021301f
C321 VTAIL.n270 VSUBS 0.011446f
C322 VTAIL.n271 VSUBS 0.027055f
C323 VTAIL.n272 VSUBS 0.01212f
C324 VTAIL.n273 VSUBS 0.021301f
C325 VTAIL.n274 VSUBS 0.011783f
C326 VTAIL.n275 VSUBS 0.027055f
C327 VTAIL.n276 VSUBS 0.011446f
C328 VTAIL.n277 VSUBS 0.01212f
C329 VTAIL.n278 VSUBS 0.021301f
C330 VTAIL.n279 VSUBS 0.011446f
C331 VTAIL.n280 VSUBS 0.027055f
C332 VTAIL.n281 VSUBS 0.01212f
C333 VTAIL.n282 VSUBS 0.021301f
C334 VTAIL.n283 VSUBS 0.011446f
C335 VTAIL.n284 VSUBS 0.020291f
C336 VTAIL.n285 VSUBS 0.020352f
C337 VTAIL.t1 VSUBS 0.058307f
C338 VTAIL.n286 VSUBS 0.168628f
C339 VTAIL.n287 VSUBS 1.05501f
C340 VTAIL.n288 VSUBS 0.011446f
C341 VTAIL.n289 VSUBS 0.01212f
C342 VTAIL.n290 VSUBS 0.027055f
C343 VTAIL.n291 VSUBS 0.027055f
C344 VTAIL.n292 VSUBS 0.01212f
C345 VTAIL.n293 VSUBS 0.011446f
C346 VTAIL.n294 VSUBS 0.021301f
C347 VTAIL.n295 VSUBS 0.021301f
C348 VTAIL.n296 VSUBS 0.011446f
C349 VTAIL.n297 VSUBS 0.01212f
C350 VTAIL.n298 VSUBS 0.027055f
C351 VTAIL.n299 VSUBS 0.027055f
C352 VTAIL.n300 VSUBS 0.01212f
C353 VTAIL.n301 VSUBS 0.011446f
C354 VTAIL.n302 VSUBS 0.021301f
C355 VTAIL.n303 VSUBS 0.021301f
C356 VTAIL.n304 VSUBS 0.011446f
C357 VTAIL.n305 VSUBS 0.01212f
C358 VTAIL.n306 VSUBS 0.027055f
C359 VTAIL.n307 VSUBS 0.027055f
C360 VTAIL.n308 VSUBS 0.027055f
C361 VTAIL.n309 VSUBS 0.011783f
C362 VTAIL.n310 VSUBS 0.011446f
C363 VTAIL.n311 VSUBS 0.021301f
C364 VTAIL.n312 VSUBS 0.021301f
C365 VTAIL.n313 VSUBS 0.011446f
C366 VTAIL.n314 VSUBS 0.01212f
C367 VTAIL.n315 VSUBS 0.027055f
C368 VTAIL.n316 VSUBS 0.027055f
C369 VTAIL.n317 VSUBS 0.01212f
C370 VTAIL.n318 VSUBS 0.011446f
C371 VTAIL.n319 VSUBS 0.021301f
C372 VTAIL.n320 VSUBS 0.021301f
C373 VTAIL.n321 VSUBS 0.011446f
C374 VTAIL.n322 VSUBS 0.01212f
C375 VTAIL.n323 VSUBS 0.027055f
C376 VTAIL.n324 VSUBS 0.064272f
C377 VTAIL.n325 VSUBS 0.01212f
C378 VTAIL.n326 VSUBS 0.011446f
C379 VTAIL.n327 VSUBS 0.048364f
C380 VTAIL.n328 VSUBS 0.03224f
C381 VTAIL.n329 VSUBS 0.093143f
C382 VTAIL.n330 VSUBS 0.023046f
C383 VTAIL.n331 VSUBS 0.021301f
C384 VTAIL.n332 VSUBS 0.011446f
C385 VTAIL.n333 VSUBS 0.027055f
C386 VTAIL.n334 VSUBS 0.01212f
C387 VTAIL.n335 VSUBS 0.021301f
C388 VTAIL.n336 VSUBS 0.011446f
C389 VTAIL.n337 VSUBS 0.027055f
C390 VTAIL.n338 VSUBS 0.01212f
C391 VTAIL.n339 VSUBS 0.021301f
C392 VTAIL.n340 VSUBS 0.011783f
C393 VTAIL.n341 VSUBS 0.027055f
C394 VTAIL.n342 VSUBS 0.011446f
C395 VTAIL.n343 VSUBS 0.01212f
C396 VTAIL.n344 VSUBS 0.021301f
C397 VTAIL.n345 VSUBS 0.011446f
C398 VTAIL.n346 VSUBS 0.027055f
C399 VTAIL.n347 VSUBS 0.01212f
C400 VTAIL.n348 VSUBS 0.021301f
C401 VTAIL.n349 VSUBS 0.011446f
C402 VTAIL.n350 VSUBS 0.020291f
C403 VTAIL.n351 VSUBS 0.020352f
C404 VTAIL.t4 VSUBS 0.058307f
C405 VTAIL.n352 VSUBS 0.168628f
C406 VTAIL.n353 VSUBS 1.05501f
C407 VTAIL.n354 VSUBS 0.011446f
C408 VTAIL.n355 VSUBS 0.01212f
C409 VTAIL.n356 VSUBS 0.027055f
C410 VTAIL.n357 VSUBS 0.027055f
C411 VTAIL.n358 VSUBS 0.01212f
C412 VTAIL.n359 VSUBS 0.011446f
C413 VTAIL.n360 VSUBS 0.021301f
C414 VTAIL.n361 VSUBS 0.021301f
C415 VTAIL.n362 VSUBS 0.011446f
C416 VTAIL.n363 VSUBS 0.01212f
C417 VTAIL.n364 VSUBS 0.027055f
C418 VTAIL.n365 VSUBS 0.027055f
C419 VTAIL.n366 VSUBS 0.01212f
C420 VTAIL.n367 VSUBS 0.011446f
C421 VTAIL.n368 VSUBS 0.021301f
C422 VTAIL.n369 VSUBS 0.021301f
C423 VTAIL.n370 VSUBS 0.011446f
C424 VTAIL.n371 VSUBS 0.01212f
C425 VTAIL.n372 VSUBS 0.027055f
C426 VTAIL.n373 VSUBS 0.027055f
C427 VTAIL.n374 VSUBS 0.027055f
C428 VTAIL.n375 VSUBS 0.011783f
C429 VTAIL.n376 VSUBS 0.011446f
C430 VTAIL.n377 VSUBS 0.021301f
C431 VTAIL.n378 VSUBS 0.021301f
C432 VTAIL.n379 VSUBS 0.011446f
C433 VTAIL.n380 VSUBS 0.01212f
C434 VTAIL.n381 VSUBS 0.027055f
C435 VTAIL.n382 VSUBS 0.027055f
C436 VTAIL.n383 VSUBS 0.01212f
C437 VTAIL.n384 VSUBS 0.011446f
C438 VTAIL.n385 VSUBS 0.021301f
C439 VTAIL.n386 VSUBS 0.021301f
C440 VTAIL.n387 VSUBS 0.011446f
C441 VTAIL.n388 VSUBS 0.01212f
C442 VTAIL.n389 VSUBS 0.027055f
C443 VTAIL.n390 VSUBS 0.064272f
C444 VTAIL.n391 VSUBS 0.01212f
C445 VTAIL.n392 VSUBS 0.011446f
C446 VTAIL.n393 VSUBS 0.048364f
C447 VTAIL.n394 VSUBS 0.03224f
C448 VTAIL.n395 VSUBS 0.093143f
C449 VTAIL.n396 VSUBS 0.023046f
C450 VTAIL.n397 VSUBS 0.021301f
C451 VTAIL.n398 VSUBS 0.011446f
C452 VTAIL.n399 VSUBS 0.027055f
C453 VTAIL.n400 VSUBS 0.01212f
C454 VTAIL.n401 VSUBS 0.021301f
C455 VTAIL.n402 VSUBS 0.011446f
C456 VTAIL.n403 VSUBS 0.027055f
C457 VTAIL.n404 VSUBS 0.01212f
C458 VTAIL.n405 VSUBS 0.021301f
C459 VTAIL.n406 VSUBS 0.011783f
C460 VTAIL.n407 VSUBS 0.027055f
C461 VTAIL.n408 VSUBS 0.011446f
C462 VTAIL.n409 VSUBS 0.01212f
C463 VTAIL.n410 VSUBS 0.021301f
C464 VTAIL.n411 VSUBS 0.011446f
C465 VTAIL.n412 VSUBS 0.027055f
C466 VTAIL.n413 VSUBS 0.01212f
C467 VTAIL.n414 VSUBS 0.021301f
C468 VTAIL.n415 VSUBS 0.011446f
C469 VTAIL.n416 VSUBS 0.020291f
C470 VTAIL.n417 VSUBS 0.020352f
C471 VTAIL.t5 VSUBS 0.058307f
C472 VTAIL.n418 VSUBS 0.168628f
C473 VTAIL.n419 VSUBS 1.05501f
C474 VTAIL.n420 VSUBS 0.011446f
C475 VTAIL.n421 VSUBS 0.01212f
C476 VTAIL.n422 VSUBS 0.027055f
C477 VTAIL.n423 VSUBS 0.027055f
C478 VTAIL.n424 VSUBS 0.01212f
C479 VTAIL.n425 VSUBS 0.011446f
C480 VTAIL.n426 VSUBS 0.021301f
C481 VTAIL.n427 VSUBS 0.021301f
C482 VTAIL.n428 VSUBS 0.011446f
C483 VTAIL.n429 VSUBS 0.01212f
C484 VTAIL.n430 VSUBS 0.027055f
C485 VTAIL.n431 VSUBS 0.027055f
C486 VTAIL.n432 VSUBS 0.01212f
C487 VTAIL.n433 VSUBS 0.011446f
C488 VTAIL.n434 VSUBS 0.021301f
C489 VTAIL.n435 VSUBS 0.021301f
C490 VTAIL.n436 VSUBS 0.011446f
C491 VTAIL.n437 VSUBS 0.01212f
C492 VTAIL.n438 VSUBS 0.027055f
C493 VTAIL.n439 VSUBS 0.027055f
C494 VTAIL.n440 VSUBS 0.027055f
C495 VTAIL.n441 VSUBS 0.011783f
C496 VTAIL.n442 VSUBS 0.011446f
C497 VTAIL.n443 VSUBS 0.021301f
C498 VTAIL.n444 VSUBS 0.021301f
C499 VTAIL.n445 VSUBS 0.011446f
C500 VTAIL.n446 VSUBS 0.01212f
C501 VTAIL.n447 VSUBS 0.027055f
C502 VTAIL.n448 VSUBS 0.027055f
C503 VTAIL.n449 VSUBS 0.01212f
C504 VTAIL.n450 VSUBS 0.011446f
C505 VTAIL.n451 VSUBS 0.021301f
C506 VTAIL.n452 VSUBS 0.021301f
C507 VTAIL.n453 VSUBS 0.011446f
C508 VTAIL.n454 VSUBS 0.01212f
C509 VTAIL.n455 VSUBS 0.027055f
C510 VTAIL.n456 VSUBS 0.064272f
C511 VTAIL.n457 VSUBS 0.01212f
C512 VTAIL.n458 VSUBS 0.011446f
C513 VTAIL.n459 VSUBS 0.048364f
C514 VTAIL.n460 VSUBS 0.03224f
C515 VTAIL.n461 VSUBS 1.10882f
C516 VTAIL.n462 VSUBS 0.023046f
C517 VTAIL.n463 VSUBS 0.021301f
C518 VTAIL.n464 VSUBS 0.011446f
C519 VTAIL.n465 VSUBS 0.027055f
C520 VTAIL.n466 VSUBS 0.01212f
C521 VTAIL.n467 VSUBS 0.021301f
C522 VTAIL.n468 VSUBS 0.011446f
C523 VTAIL.n469 VSUBS 0.027055f
C524 VTAIL.n470 VSUBS 0.01212f
C525 VTAIL.n471 VSUBS 0.021301f
C526 VTAIL.n472 VSUBS 0.011783f
C527 VTAIL.n473 VSUBS 0.027055f
C528 VTAIL.n474 VSUBS 0.01212f
C529 VTAIL.n475 VSUBS 0.021301f
C530 VTAIL.n476 VSUBS 0.011446f
C531 VTAIL.n477 VSUBS 0.027055f
C532 VTAIL.n478 VSUBS 0.01212f
C533 VTAIL.n479 VSUBS 0.021301f
C534 VTAIL.n480 VSUBS 0.011446f
C535 VTAIL.n481 VSUBS 0.020291f
C536 VTAIL.n482 VSUBS 0.020352f
C537 VTAIL.t3 VSUBS 0.058307f
C538 VTAIL.n483 VSUBS 0.168628f
C539 VTAIL.n484 VSUBS 1.05501f
C540 VTAIL.n485 VSUBS 0.011446f
C541 VTAIL.n486 VSUBS 0.01212f
C542 VTAIL.n487 VSUBS 0.027055f
C543 VTAIL.n488 VSUBS 0.027055f
C544 VTAIL.n489 VSUBS 0.01212f
C545 VTAIL.n490 VSUBS 0.011446f
C546 VTAIL.n491 VSUBS 0.021301f
C547 VTAIL.n492 VSUBS 0.021301f
C548 VTAIL.n493 VSUBS 0.011446f
C549 VTAIL.n494 VSUBS 0.01212f
C550 VTAIL.n495 VSUBS 0.027055f
C551 VTAIL.n496 VSUBS 0.027055f
C552 VTAIL.n497 VSUBS 0.01212f
C553 VTAIL.n498 VSUBS 0.011446f
C554 VTAIL.n499 VSUBS 0.021301f
C555 VTAIL.n500 VSUBS 0.021301f
C556 VTAIL.n501 VSUBS 0.011446f
C557 VTAIL.n502 VSUBS 0.011446f
C558 VTAIL.n503 VSUBS 0.01212f
C559 VTAIL.n504 VSUBS 0.027055f
C560 VTAIL.n505 VSUBS 0.027055f
C561 VTAIL.n506 VSUBS 0.027055f
C562 VTAIL.n507 VSUBS 0.011783f
C563 VTAIL.n508 VSUBS 0.011446f
C564 VTAIL.n509 VSUBS 0.021301f
C565 VTAIL.n510 VSUBS 0.021301f
C566 VTAIL.n511 VSUBS 0.011446f
C567 VTAIL.n512 VSUBS 0.01212f
C568 VTAIL.n513 VSUBS 0.027055f
C569 VTAIL.n514 VSUBS 0.027055f
C570 VTAIL.n515 VSUBS 0.01212f
C571 VTAIL.n516 VSUBS 0.011446f
C572 VTAIL.n517 VSUBS 0.021301f
C573 VTAIL.n518 VSUBS 0.021301f
C574 VTAIL.n519 VSUBS 0.011446f
C575 VTAIL.n520 VSUBS 0.01212f
C576 VTAIL.n521 VSUBS 0.027055f
C577 VTAIL.n522 VSUBS 0.064272f
C578 VTAIL.n523 VSUBS 0.01212f
C579 VTAIL.n524 VSUBS 0.011446f
C580 VTAIL.n525 VSUBS 0.048364f
C581 VTAIL.n526 VSUBS 0.03224f
C582 VTAIL.n527 VSUBS 1.08323f
C583 VP.t2 VSUBS 0.8352f
C584 VP.t3 VSUBS 0.835212f
C585 VP.n0 VSUBS 1.48279f
C586 VP.n1 VSUBS 3.75627f
C587 VP.t1 VSUBS 0.826899f
C588 VP.n2 VSUBS 0.335986f
C589 VP.t0 VSUBS 0.826899f
C590 VP.n3 VSUBS 0.335986f
C591 VP.n4 VSUBS 0.046463f
C592 B.n0 VSUBS 0.007588f
C593 B.n1 VSUBS 0.007588f
C594 B.n2 VSUBS 0.011223f
C595 B.n3 VSUBS 0.0086f
C596 B.n4 VSUBS 0.0086f
C597 B.n5 VSUBS 0.0086f
C598 B.n6 VSUBS 0.0086f
C599 B.n7 VSUBS 0.0086f
C600 B.n8 VSUBS 0.0086f
C601 B.n9 VSUBS 0.021355f
C602 B.n10 VSUBS 0.0086f
C603 B.n11 VSUBS 0.0086f
C604 B.n12 VSUBS 0.0086f
C605 B.n13 VSUBS 0.0086f
C606 B.n14 VSUBS 0.0086f
C607 B.n15 VSUBS 0.0086f
C608 B.n16 VSUBS 0.0086f
C609 B.n17 VSUBS 0.0086f
C610 B.n18 VSUBS 0.0086f
C611 B.n19 VSUBS 0.0086f
C612 B.n20 VSUBS 0.0086f
C613 B.n21 VSUBS 0.0086f
C614 B.n22 VSUBS 0.0086f
C615 B.n23 VSUBS 0.0086f
C616 B.n24 VSUBS 0.0086f
C617 B.n25 VSUBS 0.0086f
C618 B.n26 VSUBS 0.0086f
C619 B.n27 VSUBS 0.0086f
C620 B.n28 VSUBS 0.0086f
C621 B.n29 VSUBS 0.0086f
C622 B.t4 VSUBS 0.261751f
C623 B.t5 VSUBS 0.272147f
C624 B.t3 VSUBS 0.236657f
C625 B.n30 VSUBS 0.352881f
C626 B.n31 VSUBS 0.299706f
C627 B.n32 VSUBS 0.019925f
C628 B.n33 VSUBS 0.0086f
C629 B.n34 VSUBS 0.0086f
C630 B.n35 VSUBS 0.0086f
C631 B.n36 VSUBS 0.0086f
C632 B.n37 VSUBS 0.0086f
C633 B.t7 VSUBS 0.261754f
C634 B.t8 VSUBS 0.27215f
C635 B.t6 VSUBS 0.236657f
C636 B.n38 VSUBS 0.352877f
C637 B.n39 VSUBS 0.299702f
C638 B.n40 VSUBS 0.0086f
C639 B.n41 VSUBS 0.0086f
C640 B.n42 VSUBS 0.0086f
C641 B.n43 VSUBS 0.0086f
C642 B.n44 VSUBS 0.0086f
C643 B.n45 VSUBS 0.0086f
C644 B.n46 VSUBS 0.0086f
C645 B.n47 VSUBS 0.0086f
C646 B.n48 VSUBS 0.0086f
C647 B.n49 VSUBS 0.0086f
C648 B.n50 VSUBS 0.0086f
C649 B.n51 VSUBS 0.0086f
C650 B.n52 VSUBS 0.0086f
C651 B.n53 VSUBS 0.0086f
C652 B.n54 VSUBS 0.0086f
C653 B.n55 VSUBS 0.0086f
C654 B.n56 VSUBS 0.0086f
C655 B.n57 VSUBS 0.0086f
C656 B.n58 VSUBS 0.0086f
C657 B.n59 VSUBS 0.0086f
C658 B.n60 VSUBS 0.020634f
C659 B.n61 VSUBS 0.0086f
C660 B.n62 VSUBS 0.0086f
C661 B.n63 VSUBS 0.0086f
C662 B.n64 VSUBS 0.0086f
C663 B.n65 VSUBS 0.0086f
C664 B.n66 VSUBS 0.0086f
C665 B.n67 VSUBS 0.0086f
C666 B.n68 VSUBS 0.0086f
C667 B.n69 VSUBS 0.0086f
C668 B.n70 VSUBS 0.0086f
C669 B.n71 VSUBS 0.0086f
C670 B.n72 VSUBS 0.0086f
C671 B.n73 VSUBS 0.0086f
C672 B.n74 VSUBS 0.0086f
C673 B.n75 VSUBS 0.021355f
C674 B.n76 VSUBS 0.0086f
C675 B.n77 VSUBS 0.0086f
C676 B.n78 VSUBS 0.0086f
C677 B.n79 VSUBS 0.0086f
C678 B.n80 VSUBS 0.0086f
C679 B.n81 VSUBS 0.0086f
C680 B.n82 VSUBS 0.0086f
C681 B.n83 VSUBS 0.0086f
C682 B.n84 VSUBS 0.0086f
C683 B.n85 VSUBS 0.0086f
C684 B.n86 VSUBS 0.0086f
C685 B.n87 VSUBS 0.0086f
C686 B.n88 VSUBS 0.0086f
C687 B.n89 VSUBS 0.0086f
C688 B.n90 VSUBS 0.0086f
C689 B.n91 VSUBS 0.0086f
C690 B.n92 VSUBS 0.0086f
C691 B.n93 VSUBS 0.0086f
C692 B.n94 VSUBS 0.0086f
C693 B.n95 VSUBS 0.0086f
C694 B.t11 VSUBS 0.261754f
C695 B.t10 VSUBS 0.27215f
C696 B.t9 VSUBS 0.236657f
C697 B.n96 VSUBS 0.352877f
C698 B.n97 VSUBS 0.299702f
C699 B.n98 VSUBS 0.019925f
C700 B.n99 VSUBS 0.0086f
C701 B.n100 VSUBS 0.0086f
C702 B.n101 VSUBS 0.0086f
C703 B.n102 VSUBS 0.0086f
C704 B.n103 VSUBS 0.0086f
C705 B.t2 VSUBS 0.261751f
C706 B.t1 VSUBS 0.272147f
C707 B.t0 VSUBS 0.236657f
C708 B.n104 VSUBS 0.352881f
C709 B.n105 VSUBS 0.299706f
C710 B.n106 VSUBS 0.0086f
C711 B.n107 VSUBS 0.0086f
C712 B.n108 VSUBS 0.0086f
C713 B.n109 VSUBS 0.0086f
C714 B.n110 VSUBS 0.0086f
C715 B.n111 VSUBS 0.0086f
C716 B.n112 VSUBS 0.0086f
C717 B.n113 VSUBS 0.0086f
C718 B.n114 VSUBS 0.0086f
C719 B.n115 VSUBS 0.0086f
C720 B.n116 VSUBS 0.0086f
C721 B.n117 VSUBS 0.0086f
C722 B.n118 VSUBS 0.0086f
C723 B.n119 VSUBS 0.0086f
C724 B.n120 VSUBS 0.0086f
C725 B.n121 VSUBS 0.0086f
C726 B.n122 VSUBS 0.0086f
C727 B.n123 VSUBS 0.0086f
C728 B.n124 VSUBS 0.0086f
C729 B.n125 VSUBS 0.0086f
C730 B.n126 VSUBS 0.020634f
C731 B.n127 VSUBS 0.0086f
C732 B.n128 VSUBS 0.0086f
C733 B.n129 VSUBS 0.0086f
C734 B.n130 VSUBS 0.0086f
C735 B.n131 VSUBS 0.0086f
C736 B.n132 VSUBS 0.0086f
C737 B.n133 VSUBS 0.0086f
C738 B.n134 VSUBS 0.0086f
C739 B.n135 VSUBS 0.0086f
C740 B.n136 VSUBS 0.0086f
C741 B.n137 VSUBS 0.0086f
C742 B.n138 VSUBS 0.0086f
C743 B.n139 VSUBS 0.0086f
C744 B.n140 VSUBS 0.0086f
C745 B.n141 VSUBS 0.0086f
C746 B.n142 VSUBS 0.0086f
C747 B.n143 VSUBS 0.0086f
C748 B.n144 VSUBS 0.0086f
C749 B.n145 VSUBS 0.0086f
C750 B.n146 VSUBS 0.0086f
C751 B.n147 VSUBS 0.0086f
C752 B.n148 VSUBS 0.0086f
C753 B.n149 VSUBS 0.0086f
C754 B.n150 VSUBS 0.0086f
C755 B.n151 VSUBS 0.020634f
C756 B.n152 VSUBS 0.021355f
C757 B.n153 VSUBS 0.021355f
C758 B.n154 VSUBS 0.0086f
C759 B.n155 VSUBS 0.0086f
C760 B.n156 VSUBS 0.0086f
C761 B.n157 VSUBS 0.0086f
C762 B.n158 VSUBS 0.0086f
C763 B.n159 VSUBS 0.0086f
C764 B.n160 VSUBS 0.0086f
C765 B.n161 VSUBS 0.0086f
C766 B.n162 VSUBS 0.0086f
C767 B.n163 VSUBS 0.0086f
C768 B.n164 VSUBS 0.0086f
C769 B.n165 VSUBS 0.0086f
C770 B.n166 VSUBS 0.0086f
C771 B.n167 VSUBS 0.0086f
C772 B.n168 VSUBS 0.0086f
C773 B.n169 VSUBS 0.0086f
C774 B.n170 VSUBS 0.0086f
C775 B.n171 VSUBS 0.0086f
C776 B.n172 VSUBS 0.0086f
C777 B.n173 VSUBS 0.0086f
C778 B.n174 VSUBS 0.0086f
C779 B.n175 VSUBS 0.0086f
C780 B.n176 VSUBS 0.0086f
C781 B.n177 VSUBS 0.0086f
C782 B.n178 VSUBS 0.0086f
C783 B.n179 VSUBS 0.0086f
C784 B.n180 VSUBS 0.0086f
C785 B.n181 VSUBS 0.0086f
C786 B.n182 VSUBS 0.0086f
C787 B.n183 VSUBS 0.0086f
C788 B.n184 VSUBS 0.0086f
C789 B.n185 VSUBS 0.0086f
C790 B.n186 VSUBS 0.0086f
C791 B.n187 VSUBS 0.0086f
C792 B.n188 VSUBS 0.0086f
C793 B.n189 VSUBS 0.0086f
C794 B.n190 VSUBS 0.0086f
C795 B.n191 VSUBS 0.0086f
C796 B.n192 VSUBS 0.0086f
C797 B.n193 VSUBS 0.0086f
C798 B.n194 VSUBS 0.0086f
C799 B.n195 VSUBS 0.0086f
C800 B.n196 VSUBS 0.0086f
C801 B.n197 VSUBS 0.0086f
C802 B.n198 VSUBS 0.0086f
C803 B.n199 VSUBS 0.0086f
C804 B.n200 VSUBS 0.0086f
C805 B.n201 VSUBS 0.0086f
C806 B.n202 VSUBS 0.0086f
C807 B.n203 VSUBS 0.0086f
C808 B.n204 VSUBS 0.0086f
C809 B.n205 VSUBS 0.0086f
C810 B.n206 VSUBS 0.0086f
C811 B.n207 VSUBS 0.0086f
C812 B.n208 VSUBS 0.0086f
C813 B.n209 VSUBS 0.0086f
C814 B.n210 VSUBS 0.0086f
C815 B.n211 VSUBS 0.0086f
C816 B.n212 VSUBS 0.0086f
C817 B.n213 VSUBS 0.0086f
C818 B.n214 VSUBS 0.005944f
C819 B.n215 VSUBS 0.019925f
C820 B.n216 VSUBS 0.006956f
C821 B.n217 VSUBS 0.0086f
C822 B.n218 VSUBS 0.0086f
C823 B.n219 VSUBS 0.0086f
C824 B.n220 VSUBS 0.0086f
C825 B.n221 VSUBS 0.0086f
C826 B.n222 VSUBS 0.0086f
C827 B.n223 VSUBS 0.0086f
C828 B.n224 VSUBS 0.0086f
C829 B.n225 VSUBS 0.0086f
C830 B.n226 VSUBS 0.0086f
C831 B.n227 VSUBS 0.0086f
C832 B.n228 VSUBS 0.006956f
C833 B.n229 VSUBS 0.0086f
C834 B.n230 VSUBS 0.0086f
C835 B.n231 VSUBS 0.005944f
C836 B.n232 VSUBS 0.0086f
C837 B.n233 VSUBS 0.0086f
C838 B.n234 VSUBS 0.0086f
C839 B.n235 VSUBS 0.0086f
C840 B.n236 VSUBS 0.0086f
C841 B.n237 VSUBS 0.0086f
C842 B.n238 VSUBS 0.0086f
C843 B.n239 VSUBS 0.0086f
C844 B.n240 VSUBS 0.0086f
C845 B.n241 VSUBS 0.0086f
C846 B.n242 VSUBS 0.0086f
C847 B.n243 VSUBS 0.0086f
C848 B.n244 VSUBS 0.0086f
C849 B.n245 VSUBS 0.0086f
C850 B.n246 VSUBS 0.0086f
C851 B.n247 VSUBS 0.0086f
C852 B.n248 VSUBS 0.0086f
C853 B.n249 VSUBS 0.0086f
C854 B.n250 VSUBS 0.0086f
C855 B.n251 VSUBS 0.0086f
C856 B.n252 VSUBS 0.0086f
C857 B.n253 VSUBS 0.0086f
C858 B.n254 VSUBS 0.0086f
C859 B.n255 VSUBS 0.0086f
C860 B.n256 VSUBS 0.0086f
C861 B.n257 VSUBS 0.0086f
C862 B.n258 VSUBS 0.0086f
C863 B.n259 VSUBS 0.0086f
C864 B.n260 VSUBS 0.0086f
C865 B.n261 VSUBS 0.0086f
C866 B.n262 VSUBS 0.0086f
C867 B.n263 VSUBS 0.0086f
C868 B.n264 VSUBS 0.0086f
C869 B.n265 VSUBS 0.0086f
C870 B.n266 VSUBS 0.0086f
C871 B.n267 VSUBS 0.0086f
C872 B.n268 VSUBS 0.0086f
C873 B.n269 VSUBS 0.0086f
C874 B.n270 VSUBS 0.0086f
C875 B.n271 VSUBS 0.0086f
C876 B.n272 VSUBS 0.0086f
C877 B.n273 VSUBS 0.0086f
C878 B.n274 VSUBS 0.0086f
C879 B.n275 VSUBS 0.0086f
C880 B.n276 VSUBS 0.0086f
C881 B.n277 VSUBS 0.0086f
C882 B.n278 VSUBS 0.0086f
C883 B.n279 VSUBS 0.0086f
C884 B.n280 VSUBS 0.0086f
C885 B.n281 VSUBS 0.0086f
C886 B.n282 VSUBS 0.0086f
C887 B.n283 VSUBS 0.0086f
C888 B.n284 VSUBS 0.0086f
C889 B.n285 VSUBS 0.0086f
C890 B.n286 VSUBS 0.0086f
C891 B.n287 VSUBS 0.0086f
C892 B.n288 VSUBS 0.0086f
C893 B.n289 VSUBS 0.0086f
C894 B.n290 VSUBS 0.0086f
C895 B.n291 VSUBS 0.0086f
C896 B.n292 VSUBS 0.020401f
C897 B.n293 VSUBS 0.021587f
C898 B.n294 VSUBS 0.020634f
C899 B.n295 VSUBS 0.0086f
C900 B.n296 VSUBS 0.0086f
C901 B.n297 VSUBS 0.0086f
C902 B.n298 VSUBS 0.0086f
C903 B.n299 VSUBS 0.0086f
C904 B.n300 VSUBS 0.0086f
C905 B.n301 VSUBS 0.0086f
C906 B.n302 VSUBS 0.0086f
C907 B.n303 VSUBS 0.0086f
C908 B.n304 VSUBS 0.0086f
C909 B.n305 VSUBS 0.0086f
C910 B.n306 VSUBS 0.0086f
C911 B.n307 VSUBS 0.0086f
C912 B.n308 VSUBS 0.0086f
C913 B.n309 VSUBS 0.0086f
C914 B.n310 VSUBS 0.0086f
C915 B.n311 VSUBS 0.0086f
C916 B.n312 VSUBS 0.0086f
C917 B.n313 VSUBS 0.0086f
C918 B.n314 VSUBS 0.0086f
C919 B.n315 VSUBS 0.0086f
C920 B.n316 VSUBS 0.0086f
C921 B.n317 VSUBS 0.0086f
C922 B.n318 VSUBS 0.0086f
C923 B.n319 VSUBS 0.0086f
C924 B.n320 VSUBS 0.0086f
C925 B.n321 VSUBS 0.0086f
C926 B.n322 VSUBS 0.0086f
C927 B.n323 VSUBS 0.0086f
C928 B.n324 VSUBS 0.0086f
C929 B.n325 VSUBS 0.0086f
C930 B.n326 VSUBS 0.0086f
C931 B.n327 VSUBS 0.0086f
C932 B.n328 VSUBS 0.0086f
C933 B.n329 VSUBS 0.0086f
C934 B.n330 VSUBS 0.0086f
C935 B.n331 VSUBS 0.0086f
C936 B.n332 VSUBS 0.0086f
C937 B.n333 VSUBS 0.0086f
C938 B.n334 VSUBS 0.0086f
C939 B.n335 VSUBS 0.0086f
C940 B.n336 VSUBS 0.0086f
C941 B.n337 VSUBS 0.020634f
C942 B.n338 VSUBS 0.021355f
C943 B.n339 VSUBS 0.021355f
C944 B.n340 VSUBS 0.0086f
C945 B.n341 VSUBS 0.0086f
C946 B.n342 VSUBS 0.0086f
C947 B.n343 VSUBS 0.0086f
C948 B.n344 VSUBS 0.0086f
C949 B.n345 VSUBS 0.0086f
C950 B.n346 VSUBS 0.0086f
C951 B.n347 VSUBS 0.0086f
C952 B.n348 VSUBS 0.0086f
C953 B.n349 VSUBS 0.0086f
C954 B.n350 VSUBS 0.0086f
C955 B.n351 VSUBS 0.0086f
C956 B.n352 VSUBS 0.0086f
C957 B.n353 VSUBS 0.0086f
C958 B.n354 VSUBS 0.0086f
C959 B.n355 VSUBS 0.0086f
C960 B.n356 VSUBS 0.0086f
C961 B.n357 VSUBS 0.0086f
C962 B.n358 VSUBS 0.0086f
C963 B.n359 VSUBS 0.0086f
C964 B.n360 VSUBS 0.0086f
C965 B.n361 VSUBS 0.0086f
C966 B.n362 VSUBS 0.0086f
C967 B.n363 VSUBS 0.0086f
C968 B.n364 VSUBS 0.0086f
C969 B.n365 VSUBS 0.0086f
C970 B.n366 VSUBS 0.0086f
C971 B.n367 VSUBS 0.0086f
C972 B.n368 VSUBS 0.0086f
C973 B.n369 VSUBS 0.0086f
C974 B.n370 VSUBS 0.0086f
C975 B.n371 VSUBS 0.0086f
C976 B.n372 VSUBS 0.0086f
C977 B.n373 VSUBS 0.0086f
C978 B.n374 VSUBS 0.0086f
C979 B.n375 VSUBS 0.0086f
C980 B.n376 VSUBS 0.0086f
C981 B.n377 VSUBS 0.0086f
C982 B.n378 VSUBS 0.0086f
C983 B.n379 VSUBS 0.0086f
C984 B.n380 VSUBS 0.0086f
C985 B.n381 VSUBS 0.0086f
C986 B.n382 VSUBS 0.0086f
C987 B.n383 VSUBS 0.0086f
C988 B.n384 VSUBS 0.0086f
C989 B.n385 VSUBS 0.0086f
C990 B.n386 VSUBS 0.0086f
C991 B.n387 VSUBS 0.0086f
C992 B.n388 VSUBS 0.0086f
C993 B.n389 VSUBS 0.0086f
C994 B.n390 VSUBS 0.0086f
C995 B.n391 VSUBS 0.0086f
C996 B.n392 VSUBS 0.0086f
C997 B.n393 VSUBS 0.0086f
C998 B.n394 VSUBS 0.0086f
C999 B.n395 VSUBS 0.0086f
C1000 B.n396 VSUBS 0.0086f
C1001 B.n397 VSUBS 0.0086f
C1002 B.n398 VSUBS 0.0086f
C1003 B.n399 VSUBS 0.0086f
C1004 B.n400 VSUBS 0.005944f
C1005 B.n401 VSUBS 0.019925f
C1006 B.n402 VSUBS 0.006956f
C1007 B.n403 VSUBS 0.0086f
C1008 B.n404 VSUBS 0.0086f
C1009 B.n405 VSUBS 0.0086f
C1010 B.n406 VSUBS 0.0086f
C1011 B.n407 VSUBS 0.0086f
C1012 B.n408 VSUBS 0.0086f
C1013 B.n409 VSUBS 0.0086f
C1014 B.n410 VSUBS 0.0086f
C1015 B.n411 VSUBS 0.0086f
C1016 B.n412 VSUBS 0.0086f
C1017 B.n413 VSUBS 0.0086f
C1018 B.n414 VSUBS 0.006956f
C1019 B.n415 VSUBS 0.0086f
C1020 B.n416 VSUBS 0.0086f
C1021 B.n417 VSUBS 0.005944f
C1022 B.n418 VSUBS 0.0086f
C1023 B.n419 VSUBS 0.0086f
C1024 B.n420 VSUBS 0.0086f
C1025 B.n421 VSUBS 0.0086f
C1026 B.n422 VSUBS 0.0086f
C1027 B.n423 VSUBS 0.0086f
C1028 B.n424 VSUBS 0.0086f
C1029 B.n425 VSUBS 0.0086f
C1030 B.n426 VSUBS 0.0086f
C1031 B.n427 VSUBS 0.0086f
C1032 B.n428 VSUBS 0.0086f
C1033 B.n429 VSUBS 0.0086f
C1034 B.n430 VSUBS 0.0086f
C1035 B.n431 VSUBS 0.0086f
C1036 B.n432 VSUBS 0.0086f
C1037 B.n433 VSUBS 0.0086f
C1038 B.n434 VSUBS 0.0086f
C1039 B.n435 VSUBS 0.0086f
C1040 B.n436 VSUBS 0.0086f
C1041 B.n437 VSUBS 0.0086f
C1042 B.n438 VSUBS 0.0086f
C1043 B.n439 VSUBS 0.0086f
C1044 B.n440 VSUBS 0.0086f
C1045 B.n441 VSUBS 0.0086f
C1046 B.n442 VSUBS 0.0086f
C1047 B.n443 VSUBS 0.0086f
C1048 B.n444 VSUBS 0.0086f
C1049 B.n445 VSUBS 0.0086f
C1050 B.n446 VSUBS 0.0086f
C1051 B.n447 VSUBS 0.0086f
C1052 B.n448 VSUBS 0.0086f
C1053 B.n449 VSUBS 0.0086f
C1054 B.n450 VSUBS 0.0086f
C1055 B.n451 VSUBS 0.0086f
C1056 B.n452 VSUBS 0.0086f
C1057 B.n453 VSUBS 0.0086f
C1058 B.n454 VSUBS 0.0086f
C1059 B.n455 VSUBS 0.0086f
C1060 B.n456 VSUBS 0.0086f
C1061 B.n457 VSUBS 0.0086f
C1062 B.n458 VSUBS 0.0086f
C1063 B.n459 VSUBS 0.0086f
C1064 B.n460 VSUBS 0.0086f
C1065 B.n461 VSUBS 0.0086f
C1066 B.n462 VSUBS 0.0086f
C1067 B.n463 VSUBS 0.0086f
C1068 B.n464 VSUBS 0.0086f
C1069 B.n465 VSUBS 0.0086f
C1070 B.n466 VSUBS 0.0086f
C1071 B.n467 VSUBS 0.0086f
C1072 B.n468 VSUBS 0.0086f
C1073 B.n469 VSUBS 0.0086f
C1074 B.n470 VSUBS 0.0086f
C1075 B.n471 VSUBS 0.0086f
C1076 B.n472 VSUBS 0.0086f
C1077 B.n473 VSUBS 0.0086f
C1078 B.n474 VSUBS 0.0086f
C1079 B.n475 VSUBS 0.0086f
C1080 B.n476 VSUBS 0.0086f
C1081 B.n477 VSUBS 0.0086f
C1082 B.n478 VSUBS 0.021355f
C1083 B.n479 VSUBS 0.020634f
C1084 B.n480 VSUBS 0.020634f
C1085 B.n481 VSUBS 0.0086f
C1086 B.n482 VSUBS 0.0086f
C1087 B.n483 VSUBS 0.0086f
C1088 B.n484 VSUBS 0.0086f
C1089 B.n485 VSUBS 0.0086f
C1090 B.n486 VSUBS 0.0086f
C1091 B.n487 VSUBS 0.0086f
C1092 B.n488 VSUBS 0.0086f
C1093 B.n489 VSUBS 0.0086f
C1094 B.n490 VSUBS 0.0086f
C1095 B.n491 VSUBS 0.0086f
C1096 B.n492 VSUBS 0.0086f
C1097 B.n493 VSUBS 0.0086f
C1098 B.n494 VSUBS 0.0086f
C1099 B.n495 VSUBS 0.0086f
C1100 B.n496 VSUBS 0.0086f
C1101 B.n497 VSUBS 0.0086f
C1102 B.n498 VSUBS 0.0086f
C1103 B.n499 VSUBS 0.011223f
C1104 B.n500 VSUBS 0.011955f
C1105 B.n501 VSUBS 0.023773f
.ends

