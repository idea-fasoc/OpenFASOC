* NGSPICE file created from diff_pair_sample_0024.ext - technology: sky130A

.subckt diff_pair_sample_0024 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t12 w_n4190_n3512# sky130_fd_pr__pfet_01v8 ad=2.0988 pd=13.05 as=2.0988 ps=13.05 w=12.72 l=2.89
X1 VTAIL.t0 VN.t0 VDD2.t7 w_n4190_n3512# sky130_fd_pr__pfet_01v8 ad=2.0988 pd=13.05 as=2.0988 ps=13.05 w=12.72 l=2.89
X2 VTAIL.t3 VN.t1 VDD2.t6 w_n4190_n3512# sky130_fd_pr__pfet_01v8 ad=4.9608 pd=26.22 as=2.0988 ps=13.05 w=12.72 l=2.89
X3 VDD2.t5 VN.t2 VTAIL.t1 w_n4190_n3512# sky130_fd_pr__pfet_01v8 ad=2.0988 pd=13.05 as=4.9608 ps=26.22 w=12.72 l=2.89
X4 VTAIL.t8 VP.t1 VDD1.t6 w_n4190_n3512# sky130_fd_pr__pfet_01v8 ad=4.9608 pd=26.22 as=2.0988 ps=13.05 w=12.72 l=2.89
X5 VDD1.t5 VP.t2 VTAIL.t11 w_n4190_n3512# sky130_fd_pr__pfet_01v8 ad=2.0988 pd=13.05 as=4.9608 ps=26.22 w=12.72 l=2.89
X6 VTAIL.t6 VN.t3 VDD2.t4 w_n4190_n3512# sky130_fd_pr__pfet_01v8 ad=2.0988 pd=13.05 as=2.0988 ps=13.05 w=12.72 l=2.89
X7 VTAIL.t15 VP.t3 VDD1.t4 w_n4190_n3512# sky130_fd_pr__pfet_01v8 ad=2.0988 pd=13.05 as=2.0988 ps=13.05 w=12.72 l=2.89
X8 VDD2.t3 VN.t4 VTAIL.t2 w_n4190_n3512# sky130_fd_pr__pfet_01v8 ad=2.0988 pd=13.05 as=4.9608 ps=26.22 w=12.72 l=2.89
X9 VDD1.t3 VP.t4 VTAIL.t14 w_n4190_n3512# sky130_fd_pr__pfet_01v8 ad=2.0988 pd=13.05 as=2.0988 ps=13.05 w=12.72 l=2.89
X10 VDD2.t2 VN.t5 VTAIL.t4 w_n4190_n3512# sky130_fd_pr__pfet_01v8 ad=2.0988 pd=13.05 as=2.0988 ps=13.05 w=12.72 l=2.89
X11 VDD1.t2 VP.t5 VTAIL.t10 w_n4190_n3512# sky130_fd_pr__pfet_01v8 ad=2.0988 pd=13.05 as=4.9608 ps=26.22 w=12.72 l=2.89
X12 B.t11 B.t9 B.t10 w_n4190_n3512# sky130_fd_pr__pfet_01v8 ad=4.9608 pd=26.22 as=0 ps=0 w=12.72 l=2.89
X13 VDD2.t1 VN.t6 VTAIL.t7 w_n4190_n3512# sky130_fd_pr__pfet_01v8 ad=2.0988 pd=13.05 as=2.0988 ps=13.05 w=12.72 l=2.89
X14 VTAIL.t5 VN.t7 VDD2.t0 w_n4190_n3512# sky130_fd_pr__pfet_01v8 ad=4.9608 pd=26.22 as=2.0988 ps=13.05 w=12.72 l=2.89
X15 B.t8 B.t6 B.t7 w_n4190_n3512# sky130_fd_pr__pfet_01v8 ad=4.9608 pd=26.22 as=0 ps=0 w=12.72 l=2.89
X16 VTAIL.t9 VP.t6 VDD1.t1 w_n4190_n3512# sky130_fd_pr__pfet_01v8 ad=4.9608 pd=26.22 as=2.0988 ps=13.05 w=12.72 l=2.89
X17 B.t5 B.t3 B.t4 w_n4190_n3512# sky130_fd_pr__pfet_01v8 ad=4.9608 pd=26.22 as=0 ps=0 w=12.72 l=2.89
X18 VTAIL.t13 VP.t7 VDD1.t0 w_n4190_n3512# sky130_fd_pr__pfet_01v8 ad=2.0988 pd=13.05 as=2.0988 ps=13.05 w=12.72 l=2.89
X19 B.t2 B.t0 B.t1 w_n4190_n3512# sky130_fd_pr__pfet_01v8 ad=4.9608 pd=26.22 as=0 ps=0 w=12.72 l=2.89
R0 VP.n19 VP.n16 161.3
R1 VP.n21 VP.n20 161.3
R2 VP.n22 VP.n15 161.3
R3 VP.n24 VP.n23 161.3
R4 VP.n25 VP.n14 161.3
R5 VP.n28 VP.n27 161.3
R6 VP.n29 VP.n13 161.3
R7 VP.n31 VP.n30 161.3
R8 VP.n32 VP.n12 161.3
R9 VP.n34 VP.n33 161.3
R10 VP.n35 VP.n11 161.3
R11 VP.n37 VP.n36 161.3
R12 VP.n38 VP.n10 161.3
R13 VP.n74 VP.n0 161.3
R14 VP.n73 VP.n72 161.3
R15 VP.n71 VP.n1 161.3
R16 VP.n70 VP.n69 161.3
R17 VP.n68 VP.n2 161.3
R18 VP.n67 VP.n66 161.3
R19 VP.n65 VP.n3 161.3
R20 VP.n64 VP.n63 161.3
R21 VP.n61 VP.n4 161.3
R22 VP.n60 VP.n59 161.3
R23 VP.n58 VP.n5 161.3
R24 VP.n57 VP.n56 161.3
R25 VP.n55 VP.n6 161.3
R26 VP.n53 VP.n52 161.3
R27 VP.n51 VP.n7 161.3
R28 VP.n50 VP.n49 161.3
R29 VP.n48 VP.n8 161.3
R30 VP.n47 VP.n46 161.3
R31 VP.n45 VP.n9 161.3
R32 VP.n44 VP.n43 161.3
R33 VP.n17 VP.t6 139.519
R34 VP.n42 VP.n41 106.712
R35 VP.n76 VP.n75 106.712
R36 VP.n40 VP.n39 106.712
R37 VP.n42 VP.t1 106.073
R38 VP.n54 VP.t0 106.073
R39 VP.n62 VP.t7 106.073
R40 VP.n75 VP.t5 106.073
R41 VP.n39 VP.t2 106.073
R42 VP.n26 VP.t3 106.073
R43 VP.n18 VP.t4 106.073
R44 VP.n60 VP.n5 56.4773
R45 VP.n24 VP.n15 56.4773
R46 VP.n18 VP.n17 55.9247
R47 VP.n41 VP.n40 52.795
R48 VP.n49 VP.n48 43.3318
R49 VP.n69 VP.n68 43.3318
R50 VP.n33 VP.n32 43.3318
R51 VP.n48 VP.n47 37.4894
R52 VP.n69 VP.n1 37.4894
R53 VP.n33 VP.n11 37.4894
R54 VP.n43 VP.n9 24.3439
R55 VP.n47 VP.n9 24.3439
R56 VP.n49 VP.n7 24.3439
R57 VP.n53 VP.n7 24.3439
R58 VP.n56 VP.n55 24.3439
R59 VP.n56 VP.n5 24.3439
R60 VP.n61 VP.n60 24.3439
R61 VP.n63 VP.n61 24.3439
R62 VP.n67 VP.n3 24.3439
R63 VP.n68 VP.n67 24.3439
R64 VP.n73 VP.n1 24.3439
R65 VP.n74 VP.n73 24.3439
R66 VP.n37 VP.n11 24.3439
R67 VP.n38 VP.n37 24.3439
R68 VP.n25 VP.n24 24.3439
R69 VP.n27 VP.n25 24.3439
R70 VP.n31 VP.n13 24.3439
R71 VP.n32 VP.n31 24.3439
R72 VP.n20 VP.n19 24.3439
R73 VP.n20 VP.n15 24.3439
R74 VP.n55 VP.n54 17.5278
R75 VP.n63 VP.n62 17.5278
R76 VP.n27 VP.n26 17.5278
R77 VP.n19 VP.n18 17.5278
R78 VP.n54 VP.n53 6.81666
R79 VP.n62 VP.n3 6.81666
R80 VP.n26 VP.n13 6.81666
R81 VP.n17 VP.n16 5.04473
R82 VP.n43 VP.n42 3.89545
R83 VP.n75 VP.n74 3.89545
R84 VP.n39 VP.n38 3.89545
R85 VP.n40 VP.n10 0.278398
R86 VP.n44 VP.n41 0.278398
R87 VP.n76 VP.n0 0.278398
R88 VP.n21 VP.n16 0.189894
R89 VP.n22 VP.n21 0.189894
R90 VP.n23 VP.n22 0.189894
R91 VP.n23 VP.n14 0.189894
R92 VP.n28 VP.n14 0.189894
R93 VP.n29 VP.n28 0.189894
R94 VP.n30 VP.n29 0.189894
R95 VP.n30 VP.n12 0.189894
R96 VP.n34 VP.n12 0.189894
R97 VP.n35 VP.n34 0.189894
R98 VP.n36 VP.n35 0.189894
R99 VP.n36 VP.n10 0.189894
R100 VP.n45 VP.n44 0.189894
R101 VP.n46 VP.n45 0.189894
R102 VP.n46 VP.n8 0.189894
R103 VP.n50 VP.n8 0.189894
R104 VP.n51 VP.n50 0.189894
R105 VP.n52 VP.n51 0.189894
R106 VP.n52 VP.n6 0.189894
R107 VP.n57 VP.n6 0.189894
R108 VP.n58 VP.n57 0.189894
R109 VP.n59 VP.n58 0.189894
R110 VP.n59 VP.n4 0.189894
R111 VP.n64 VP.n4 0.189894
R112 VP.n65 VP.n64 0.189894
R113 VP.n66 VP.n65 0.189894
R114 VP.n66 VP.n2 0.189894
R115 VP.n70 VP.n2 0.189894
R116 VP.n71 VP.n70 0.189894
R117 VP.n72 VP.n71 0.189894
R118 VP.n72 VP.n0 0.189894
R119 VP VP.n76 0.153422
R120 VTAIL.n562 VTAIL.n498 756.745
R121 VTAIL.n66 VTAIL.n2 756.745
R122 VTAIL.n136 VTAIL.n72 756.745
R123 VTAIL.n208 VTAIL.n144 756.745
R124 VTAIL.n492 VTAIL.n428 756.745
R125 VTAIL.n420 VTAIL.n356 756.745
R126 VTAIL.n350 VTAIL.n286 756.745
R127 VTAIL.n278 VTAIL.n214 756.745
R128 VTAIL.n521 VTAIL.n520 585
R129 VTAIL.n518 VTAIL.n517 585
R130 VTAIL.n527 VTAIL.n526 585
R131 VTAIL.n529 VTAIL.n528 585
R132 VTAIL.n514 VTAIL.n513 585
R133 VTAIL.n535 VTAIL.n534 585
R134 VTAIL.n538 VTAIL.n537 585
R135 VTAIL.n536 VTAIL.n510 585
R136 VTAIL.n543 VTAIL.n509 585
R137 VTAIL.n545 VTAIL.n544 585
R138 VTAIL.n547 VTAIL.n546 585
R139 VTAIL.n506 VTAIL.n505 585
R140 VTAIL.n553 VTAIL.n552 585
R141 VTAIL.n555 VTAIL.n554 585
R142 VTAIL.n502 VTAIL.n501 585
R143 VTAIL.n561 VTAIL.n560 585
R144 VTAIL.n563 VTAIL.n562 585
R145 VTAIL.n25 VTAIL.n24 585
R146 VTAIL.n22 VTAIL.n21 585
R147 VTAIL.n31 VTAIL.n30 585
R148 VTAIL.n33 VTAIL.n32 585
R149 VTAIL.n18 VTAIL.n17 585
R150 VTAIL.n39 VTAIL.n38 585
R151 VTAIL.n42 VTAIL.n41 585
R152 VTAIL.n40 VTAIL.n14 585
R153 VTAIL.n47 VTAIL.n13 585
R154 VTAIL.n49 VTAIL.n48 585
R155 VTAIL.n51 VTAIL.n50 585
R156 VTAIL.n10 VTAIL.n9 585
R157 VTAIL.n57 VTAIL.n56 585
R158 VTAIL.n59 VTAIL.n58 585
R159 VTAIL.n6 VTAIL.n5 585
R160 VTAIL.n65 VTAIL.n64 585
R161 VTAIL.n67 VTAIL.n66 585
R162 VTAIL.n95 VTAIL.n94 585
R163 VTAIL.n92 VTAIL.n91 585
R164 VTAIL.n101 VTAIL.n100 585
R165 VTAIL.n103 VTAIL.n102 585
R166 VTAIL.n88 VTAIL.n87 585
R167 VTAIL.n109 VTAIL.n108 585
R168 VTAIL.n112 VTAIL.n111 585
R169 VTAIL.n110 VTAIL.n84 585
R170 VTAIL.n117 VTAIL.n83 585
R171 VTAIL.n119 VTAIL.n118 585
R172 VTAIL.n121 VTAIL.n120 585
R173 VTAIL.n80 VTAIL.n79 585
R174 VTAIL.n127 VTAIL.n126 585
R175 VTAIL.n129 VTAIL.n128 585
R176 VTAIL.n76 VTAIL.n75 585
R177 VTAIL.n135 VTAIL.n134 585
R178 VTAIL.n137 VTAIL.n136 585
R179 VTAIL.n167 VTAIL.n166 585
R180 VTAIL.n164 VTAIL.n163 585
R181 VTAIL.n173 VTAIL.n172 585
R182 VTAIL.n175 VTAIL.n174 585
R183 VTAIL.n160 VTAIL.n159 585
R184 VTAIL.n181 VTAIL.n180 585
R185 VTAIL.n184 VTAIL.n183 585
R186 VTAIL.n182 VTAIL.n156 585
R187 VTAIL.n189 VTAIL.n155 585
R188 VTAIL.n191 VTAIL.n190 585
R189 VTAIL.n193 VTAIL.n192 585
R190 VTAIL.n152 VTAIL.n151 585
R191 VTAIL.n199 VTAIL.n198 585
R192 VTAIL.n201 VTAIL.n200 585
R193 VTAIL.n148 VTAIL.n147 585
R194 VTAIL.n207 VTAIL.n206 585
R195 VTAIL.n209 VTAIL.n208 585
R196 VTAIL.n493 VTAIL.n492 585
R197 VTAIL.n491 VTAIL.n490 585
R198 VTAIL.n432 VTAIL.n431 585
R199 VTAIL.n485 VTAIL.n484 585
R200 VTAIL.n483 VTAIL.n482 585
R201 VTAIL.n436 VTAIL.n435 585
R202 VTAIL.n477 VTAIL.n476 585
R203 VTAIL.n475 VTAIL.n474 585
R204 VTAIL.n473 VTAIL.n439 585
R205 VTAIL.n443 VTAIL.n440 585
R206 VTAIL.n468 VTAIL.n467 585
R207 VTAIL.n466 VTAIL.n465 585
R208 VTAIL.n445 VTAIL.n444 585
R209 VTAIL.n460 VTAIL.n459 585
R210 VTAIL.n458 VTAIL.n457 585
R211 VTAIL.n449 VTAIL.n448 585
R212 VTAIL.n452 VTAIL.n451 585
R213 VTAIL.n421 VTAIL.n420 585
R214 VTAIL.n419 VTAIL.n418 585
R215 VTAIL.n360 VTAIL.n359 585
R216 VTAIL.n413 VTAIL.n412 585
R217 VTAIL.n411 VTAIL.n410 585
R218 VTAIL.n364 VTAIL.n363 585
R219 VTAIL.n405 VTAIL.n404 585
R220 VTAIL.n403 VTAIL.n402 585
R221 VTAIL.n401 VTAIL.n367 585
R222 VTAIL.n371 VTAIL.n368 585
R223 VTAIL.n396 VTAIL.n395 585
R224 VTAIL.n394 VTAIL.n393 585
R225 VTAIL.n373 VTAIL.n372 585
R226 VTAIL.n388 VTAIL.n387 585
R227 VTAIL.n386 VTAIL.n385 585
R228 VTAIL.n377 VTAIL.n376 585
R229 VTAIL.n380 VTAIL.n379 585
R230 VTAIL.n351 VTAIL.n350 585
R231 VTAIL.n349 VTAIL.n348 585
R232 VTAIL.n290 VTAIL.n289 585
R233 VTAIL.n343 VTAIL.n342 585
R234 VTAIL.n341 VTAIL.n340 585
R235 VTAIL.n294 VTAIL.n293 585
R236 VTAIL.n335 VTAIL.n334 585
R237 VTAIL.n333 VTAIL.n332 585
R238 VTAIL.n331 VTAIL.n297 585
R239 VTAIL.n301 VTAIL.n298 585
R240 VTAIL.n326 VTAIL.n325 585
R241 VTAIL.n324 VTAIL.n323 585
R242 VTAIL.n303 VTAIL.n302 585
R243 VTAIL.n318 VTAIL.n317 585
R244 VTAIL.n316 VTAIL.n315 585
R245 VTAIL.n307 VTAIL.n306 585
R246 VTAIL.n310 VTAIL.n309 585
R247 VTAIL.n279 VTAIL.n278 585
R248 VTAIL.n277 VTAIL.n276 585
R249 VTAIL.n218 VTAIL.n217 585
R250 VTAIL.n271 VTAIL.n270 585
R251 VTAIL.n269 VTAIL.n268 585
R252 VTAIL.n222 VTAIL.n221 585
R253 VTAIL.n263 VTAIL.n262 585
R254 VTAIL.n261 VTAIL.n260 585
R255 VTAIL.n259 VTAIL.n225 585
R256 VTAIL.n229 VTAIL.n226 585
R257 VTAIL.n254 VTAIL.n253 585
R258 VTAIL.n252 VTAIL.n251 585
R259 VTAIL.n231 VTAIL.n230 585
R260 VTAIL.n246 VTAIL.n245 585
R261 VTAIL.n244 VTAIL.n243 585
R262 VTAIL.n235 VTAIL.n234 585
R263 VTAIL.n238 VTAIL.n237 585
R264 VTAIL.t1 VTAIL.n519 329.036
R265 VTAIL.t5 VTAIL.n23 329.036
R266 VTAIL.t10 VTAIL.n93 329.036
R267 VTAIL.t8 VTAIL.n165 329.036
R268 VTAIL.t11 VTAIL.n450 329.036
R269 VTAIL.t9 VTAIL.n378 329.036
R270 VTAIL.t2 VTAIL.n308 329.036
R271 VTAIL.t3 VTAIL.n236 329.036
R272 VTAIL.n520 VTAIL.n517 171.744
R273 VTAIL.n527 VTAIL.n517 171.744
R274 VTAIL.n528 VTAIL.n527 171.744
R275 VTAIL.n528 VTAIL.n513 171.744
R276 VTAIL.n535 VTAIL.n513 171.744
R277 VTAIL.n537 VTAIL.n535 171.744
R278 VTAIL.n537 VTAIL.n536 171.744
R279 VTAIL.n536 VTAIL.n509 171.744
R280 VTAIL.n545 VTAIL.n509 171.744
R281 VTAIL.n546 VTAIL.n545 171.744
R282 VTAIL.n546 VTAIL.n505 171.744
R283 VTAIL.n553 VTAIL.n505 171.744
R284 VTAIL.n554 VTAIL.n553 171.744
R285 VTAIL.n554 VTAIL.n501 171.744
R286 VTAIL.n561 VTAIL.n501 171.744
R287 VTAIL.n562 VTAIL.n561 171.744
R288 VTAIL.n24 VTAIL.n21 171.744
R289 VTAIL.n31 VTAIL.n21 171.744
R290 VTAIL.n32 VTAIL.n31 171.744
R291 VTAIL.n32 VTAIL.n17 171.744
R292 VTAIL.n39 VTAIL.n17 171.744
R293 VTAIL.n41 VTAIL.n39 171.744
R294 VTAIL.n41 VTAIL.n40 171.744
R295 VTAIL.n40 VTAIL.n13 171.744
R296 VTAIL.n49 VTAIL.n13 171.744
R297 VTAIL.n50 VTAIL.n49 171.744
R298 VTAIL.n50 VTAIL.n9 171.744
R299 VTAIL.n57 VTAIL.n9 171.744
R300 VTAIL.n58 VTAIL.n57 171.744
R301 VTAIL.n58 VTAIL.n5 171.744
R302 VTAIL.n65 VTAIL.n5 171.744
R303 VTAIL.n66 VTAIL.n65 171.744
R304 VTAIL.n94 VTAIL.n91 171.744
R305 VTAIL.n101 VTAIL.n91 171.744
R306 VTAIL.n102 VTAIL.n101 171.744
R307 VTAIL.n102 VTAIL.n87 171.744
R308 VTAIL.n109 VTAIL.n87 171.744
R309 VTAIL.n111 VTAIL.n109 171.744
R310 VTAIL.n111 VTAIL.n110 171.744
R311 VTAIL.n110 VTAIL.n83 171.744
R312 VTAIL.n119 VTAIL.n83 171.744
R313 VTAIL.n120 VTAIL.n119 171.744
R314 VTAIL.n120 VTAIL.n79 171.744
R315 VTAIL.n127 VTAIL.n79 171.744
R316 VTAIL.n128 VTAIL.n127 171.744
R317 VTAIL.n128 VTAIL.n75 171.744
R318 VTAIL.n135 VTAIL.n75 171.744
R319 VTAIL.n136 VTAIL.n135 171.744
R320 VTAIL.n166 VTAIL.n163 171.744
R321 VTAIL.n173 VTAIL.n163 171.744
R322 VTAIL.n174 VTAIL.n173 171.744
R323 VTAIL.n174 VTAIL.n159 171.744
R324 VTAIL.n181 VTAIL.n159 171.744
R325 VTAIL.n183 VTAIL.n181 171.744
R326 VTAIL.n183 VTAIL.n182 171.744
R327 VTAIL.n182 VTAIL.n155 171.744
R328 VTAIL.n191 VTAIL.n155 171.744
R329 VTAIL.n192 VTAIL.n191 171.744
R330 VTAIL.n192 VTAIL.n151 171.744
R331 VTAIL.n199 VTAIL.n151 171.744
R332 VTAIL.n200 VTAIL.n199 171.744
R333 VTAIL.n200 VTAIL.n147 171.744
R334 VTAIL.n207 VTAIL.n147 171.744
R335 VTAIL.n208 VTAIL.n207 171.744
R336 VTAIL.n492 VTAIL.n491 171.744
R337 VTAIL.n491 VTAIL.n431 171.744
R338 VTAIL.n484 VTAIL.n431 171.744
R339 VTAIL.n484 VTAIL.n483 171.744
R340 VTAIL.n483 VTAIL.n435 171.744
R341 VTAIL.n476 VTAIL.n435 171.744
R342 VTAIL.n476 VTAIL.n475 171.744
R343 VTAIL.n475 VTAIL.n439 171.744
R344 VTAIL.n443 VTAIL.n439 171.744
R345 VTAIL.n467 VTAIL.n443 171.744
R346 VTAIL.n467 VTAIL.n466 171.744
R347 VTAIL.n466 VTAIL.n444 171.744
R348 VTAIL.n459 VTAIL.n444 171.744
R349 VTAIL.n459 VTAIL.n458 171.744
R350 VTAIL.n458 VTAIL.n448 171.744
R351 VTAIL.n451 VTAIL.n448 171.744
R352 VTAIL.n420 VTAIL.n419 171.744
R353 VTAIL.n419 VTAIL.n359 171.744
R354 VTAIL.n412 VTAIL.n359 171.744
R355 VTAIL.n412 VTAIL.n411 171.744
R356 VTAIL.n411 VTAIL.n363 171.744
R357 VTAIL.n404 VTAIL.n363 171.744
R358 VTAIL.n404 VTAIL.n403 171.744
R359 VTAIL.n403 VTAIL.n367 171.744
R360 VTAIL.n371 VTAIL.n367 171.744
R361 VTAIL.n395 VTAIL.n371 171.744
R362 VTAIL.n395 VTAIL.n394 171.744
R363 VTAIL.n394 VTAIL.n372 171.744
R364 VTAIL.n387 VTAIL.n372 171.744
R365 VTAIL.n387 VTAIL.n386 171.744
R366 VTAIL.n386 VTAIL.n376 171.744
R367 VTAIL.n379 VTAIL.n376 171.744
R368 VTAIL.n350 VTAIL.n349 171.744
R369 VTAIL.n349 VTAIL.n289 171.744
R370 VTAIL.n342 VTAIL.n289 171.744
R371 VTAIL.n342 VTAIL.n341 171.744
R372 VTAIL.n341 VTAIL.n293 171.744
R373 VTAIL.n334 VTAIL.n293 171.744
R374 VTAIL.n334 VTAIL.n333 171.744
R375 VTAIL.n333 VTAIL.n297 171.744
R376 VTAIL.n301 VTAIL.n297 171.744
R377 VTAIL.n325 VTAIL.n301 171.744
R378 VTAIL.n325 VTAIL.n324 171.744
R379 VTAIL.n324 VTAIL.n302 171.744
R380 VTAIL.n317 VTAIL.n302 171.744
R381 VTAIL.n317 VTAIL.n316 171.744
R382 VTAIL.n316 VTAIL.n306 171.744
R383 VTAIL.n309 VTAIL.n306 171.744
R384 VTAIL.n278 VTAIL.n277 171.744
R385 VTAIL.n277 VTAIL.n217 171.744
R386 VTAIL.n270 VTAIL.n217 171.744
R387 VTAIL.n270 VTAIL.n269 171.744
R388 VTAIL.n269 VTAIL.n221 171.744
R389 VTAIL.n262 VTAIL.n221 171.744
R390 VTAIL.n262 VTAIL.n261 171.744
R391 VTAIL.n261 VTAIL.n225 171.744
R392 VTAIL.n229 VTAIL.n225 171.744
R393 VTAIL.n253 VTAIL.n229 171.744
R394 VTAIL.n253 VTAIL.n252 171.744
R395 VTAIL.n252 VTAIL.n230 171.744
R396 VTAIL.n245 VTAIL.n230 171.744
R397 VTAIL.n245 VTAIL.n244 171.744
R398 VTAIL.n244 VTAIL.n234 171.744
R399 VTAIL.n237 VTAIL.n234 171.744
R400 VTAIL.n520 VTAIL.t1 85.8723
R401 VTAIL.n24 VTAIL.t5 85.8723
R402 VTAIL.n94 VTAIL.t10 85.8723
R403 VTAIL.n166 VTAIL.t8 85.8723
R404 VTAIL.n451 VTAIL.t11 85.8723
R405 VTAIL.n379 VTAIL.t9 85.8723
R406 VTAIL.n309 VTAIL.t2 85.8723
R407 VTAIL.n237 VTAIL.t3 85.8723
R408 VTAIL.n1 VTAIL.n0 54.0053
R409 VTAIL.n143 VTAIL.n142 54.0053
R410 VTAIL.n427 VTAIL.n426 54.0053
R411 VTAIL.n285 VTAIL.n284 54.0053
R412 VTAIL.n567 VTAIL.n566 29.8581
R413 VTAIL.n71 VTAIL.n70 29.8581
R414 VTAIL.n141 VTAIL.n140 29.8581
R415 VTAIL.n213 VTAIL.n212 29.8581
R416 VTAIL.n497 VTAIL.n496 29.8581
R417 VTAIL.n425 VTAIL.n424 29.8581
R418 VTAIL.n355 VTAIL.n354 29.8581
R419 VTAIL.n283 VTAIL.n282 29.8581
R420 VTAIL.n567 VTAIL.n497 26.1083
R421 VTAIL.n283 VTAIL.n213 26.1083
R422 VTAIL.n544 VTAIL.n543 13.1884
R423 VTAIL.n48 VTAIL.n47 13.1884
R424 VTAIL.n118 VTAIL.n117 13.1884
R425 VTAIL.n190 VTAIL.n189 13.1884
R426 VTAIL.n474 VTAIL.n473 13.1884
R427 VTAIL.n402 VTAIL.n401 13.1884
R428 VTAIL.n332 VTAIL.n331 13.1884
R429 VTAIL.n260 VTAIL.n259 13.1884
R430 VTAIL.n542 VTAIL.n510 12.8005
R431 VTAIL.n547 VTAIL.n508 12.8005
R432 VTAIL.n46 VTAIL.n14 12.8005
R433 VTAIL.n51 VTAIL.n12 12.8005
R434 VTAIL.n116 VTAIL.n84 12.8005
R435 VTAIL.n121 VTAIL.n82 12.8005
R436 VTAIL.n188 VTAIL.n156 12.8005
R437 VTAIL.n193 VTAIL.n154 12.8005
R438 VTAIL.n477 VTAIL.n438 12.8005
R439 VTAIL.n472 VTAIL.n440 12.8005
R440 VTAIL.n405 VTAIL.n366 12.8005
R441 VTAIL.n400 VTAIL.n368 12.8005
R442 VTAIL.n335 VTAIL.n296 12.8005
R443 VTAIL.n330 VTAIL.n298 12.8005
R444 VTAIL.n263 VTAIL.n224 12.8005
R445 VTAIL.n258 VTAIL.n226 12.8005
R446 VTAIL.n539 VTAIL.n538 12.0247
R447 VTAIL.n548 VTAIL.n506 12.0247
R448 VTAIL.n43 VTAIL.n42 12.0247
R449 VTAIL.n52 VTAIL.n10 12.0247
R450 VTAIL.n113 VTAIL.n112 12.0247
R451 VTAIL.n122 VTAIL.n80 12.0247
R452 VTAIL.n185 VTAIL.n184 12.0247
R453 VTAIL.n194 VTAIL.n152 12.0247
R454 VTAIL.n478 VTAIL.n436 12.0247
R455 VTAIL.n469 VTAIL.n468 12.0247
R456 VTAIL.n406 VTAIL.n364 12.0247
R457 VTAIL.n397 VTAIL.n396 12.0247
R458 VTAIL.n336 VTAIL.n294 12.0247
R459 VTAIL.n327 VTAIL.n326 12.0247
R460 VTAIL.n264 VTAIL.n222 12.0247
R461 VTAIL.n255 VTAIL.n254 12.0247
R462 VTAIL.n534 VTAIL.n512 11.249
R463 VTAIL.n552 VTAIL.n551 11.249
R464 VTAIL.n38 VTAIL.n16 11.249
R465 VTAIL.n56 VTAIL.n55 11.249
R466 VTAIL.n108 VTAIL.n86 11.249
R467 VTAIL.n126 VTAIL.n125 11.249
R468 VTAIL.n180 VTAIL.n158 11.249
R469 VTAIL.n198 VTAIL.n197 11.249
R470 VTAIL.n482 VTAIL.n481 11.249
R471 VTAIL.n465 VTAIL.n442 11.249
R472 VTAIL.n410 VTAIL.n409 11.249
R473 VTAIL.n393 VTAIL.n370 11.249
R474 VTAIL.n340 VTAIL.n339 11.249
R475 VTAIL.n323 VTAIL.n300 11.249
R476 VTAIL.n268 VTAIL.n267 11.249
R477 VTAIL.n251 VTAIL.n228 11.249
R478 VTAIL.n521 VTAIL.n519 10.7239
R479 VTAIL.n25 VTAIL.n23 10.7239
R480 VTAIL.n95 VTAIL.n93 10.7239
R481 VTAIL.n167 VTAIL.n165 10.7239
R482 VTAIL.n452 VTAIL.n450 10.7239
R483 VTAIL.n380 VTAIL.n378 10.7239
R484 VTAIL.n310 VTAIL.n308 10.7239
R485 VTAIL.n238 VTAIL.n236 10.7239
R486 VTAIL.n533 VTAIL.n514 10.4732
R487 VTAIL.n555 VTAIL.n504 10.4732
R488 VTAIL.n37 VTAIL.n18 10.4732
R489 VTAIL.n59 VTAIL.n8 10.4732
R490 VTAIL.n107 VTAIL.n88 10.4732
R491 VTAIL.n129 VTAIL.n78 10.4732
R492 VTAIL.n179 VTAIL.n160 10.4732
R493 VTAIL.n201 VTAIL.n150 10.4732
R494 VTAIL.n485 VTAIL.n434 10.4732
R495 VTAIL.n464 VTAIL.n445 10.4732
R496 VTAIL.n413 VTAIL.n362 10.4732
R497 VTAIL.n392 VTAIL.n373 10.4732
R498 VTAIL.n343 VTAIL.n292 10.4732
R499 VTAIL.n322 VTAIL.n303 10.4732
R500 VTAIL.n271 VTAIL.n220 10.4732
R501 VTAIL.n250 VTAIL.n231 10.4732
R502 VTAIL.n530 VTAIL.n529 9.69747
R503 VTAIL.n556 VTAIL.n502 9.69747
R504 VTAIL.n34 VTAIL.n33 9.69747
R505 VTAIL.n60 VTAIL.n6 9.69747
R506 VTAIL.n104 VTAIL.n103 9.69747
R507 VTAIL.n130 VTAIL.n76 9.69747
R508 VTAIL.n176 VTAIL.n175 9.69747
R509 VTAIL.n202 VTAIL.n148 9.69747
R510 VTAIL.n486 VTAIL.n432 9.69747
R511 VTAIL.n461 VTAIL.n460 9.69747
R512 VTAIL.n414 VTAIL.n360 9.69747
R513 VTAIL.n389 VTAIL.n388 9.69747
R514 VTAIL.n344 VTAIL.n290 9.69747
R515 VTAIL.n319 VTAIL.n318 9.69747
R516 VTAIL.n272 VTAIL.n218 9.69747
R517 VTAIL.n247 VTAIL.n246 9.69747
R518 VTAIL.n566 VTAIL.n565 9.45567
R519 VTAIL.n70 VTAIL.n69 9.45567
R520 VTAIL.n140 VTAIL.n139 9.45567
R521 VTAIL.n212 VTAIL.n211 9.45567
R522 VTAIL.n496 VTAIL.n495 9.45567
R523 VTAIL.n424 VTAIL.n423 9.45567
R524 VTAIL.n354 VTAIL.n353 9.45567
R525 VTAIL.n282 VTAIL.n281 9.45567
R526 VTAIL.n500 VTAIL.n499 9.3005
R527 VTAIL.n559 VTAIL.n558 9.3005
R528 VTAIL.n557 VTAIL.n556 9.3005
R529 VTAIL.n504 VTAIL.n503 9.3005
R530 VTAIL.n551 VTAIL.n550 9.3005
R531 VTAIL.n549 VTAIL.n548 9.3005
R532 VTAIL.n508 VTAIL.n507 9.3005
R533 VTAIL.n523 VTAIL.n522 9.3005
R534 VTAIL.n525 VTAIL.n524 9.3005
R535 VTAIL.n516 VTAIL.n515 9.3005
R536 VTAIL.n531 VTAIL.n530 9.3005
R537 VTAIL.n533 VTAIL.n532 9.3005
R538 VTAIL.n512 VTAIL.n511 9.3005
R539 VTAIL.n540 VTAIL.n539 9.3005
R540 VTAIL.n542 VTAIL.n541 9.3005
R541 VTAIL.n565 VTAIL.n564 9.3005
R542 VTAIL.n4 VTAIL.n3 9.3005
R543 VTAIL.n63 VTAIL.n62 9.3005
R544 VTAIL.n61 VTAIL.n60 9.3005
R545 VTAIL.n8 VTAIL.n7 9.3005
R546 VTAIL.n55 VTAIL.n54 9.3005
R547 VTAIL.n53 VTAIL.n52 9.3005
R548 VTAIL.n12 VTAIL.n11 9.3005
R549 VTAIL.n27 VTAIL.n26 9.3005
R550 VTAIL.n29 VTAIL.n28 9.3005
R551 VTAIL.n20 VTAIL.n19 9.3005
R552 VTAIL.n35 VTAIL.n34 9.3005
R553 VTAIL.n37 VTAIL.n36 9.3005
R554 VTAIL.n16 VTAIL.n15 9.3005
R555 VTAIL.n44 VTAIL.n43 9.3005
R556 VTAIL.n46 VTAIL.n45 9.3005
R557 VTAIL.n69 VTAIL.n68 9.3005
R558 VTAIL.n74 VTAIL.n73 9.3005
R559 VTAIL.n133 VTAIL.n132 9.3005
R560 VTAIL.n131 VTAIL.n130 9.3005
R561 VTAIL.n78 VTAIL.n77 9.3005
R562 VTAIL.n125 VTAIL.n124 9.3005
R563 VTAIL.n123 VTAIL.n122 9.3005
R564 VTAIL.n82 VTAIL.n81 9.3005
R565 VTAIL.n97 VTAIL.n96 9.3005
R566 VTAIL.n99 VTAIL.n98 9.3005
R567 VTAIL.n90 VTAIL.n89 9.3005
R568 VTAIL.n105 VTAIL.n104 9.3005
R569 VTAIL.n107 VTAIL.n106 9.3005
R570 VTAIL.n86 VTAIL.n85 9.3005
R571 VTAIL.n114 VTAIL.n113 9.3005
R572 VTAIL.n116 VTAIL.n115 9.3005
R573 VTAIL.n139 VTAIL.n138 9.3005
R574 VTAIL.n146 VTAIL.n145 9.3005
R575 VTAIL.n205 VTAIL.n204 9.3005
R576 VTAIL.n203 VTAIL.n202 9.3005
R577 VTAIL.n150 VTAIL.n149 9.3005
R578 VTAIL.n197 VTAIL.n196 9.3005
R579 VTAIL.n195 VTAIL.n194 9.3005
R580 VTAIL.n154 VTAIL.n153 9.3005
R581 VTAIL.n169 VTAIL.n168 9.3005
R582 VTAIL.n171 VTAIL.n170 9.3005
R583 VTAIL.n162 VTAIL.n161 9.3005
R584 VTAIL.n177 VTAIL.n176 9.3005
R585 VTAIL.n179 VTAIL.n178 9.3005
R586 VTAIL.n158 VTAIL.n157 9.3005
R587 VTAIL.n186 VTAIL.n185 9.3005
R588 VTAIL.n188 VTAIL.n187 9.3005
R589 VTAIL.n211 VTAIL.n210 9.3005
R590 VTAIL.n454 VTAIL.n453 9.3005
R591 VTAIL.n456 VTAIL.n455 9.3005
R592 VTAIL.n447 VTAIL.n446 9.3005
R593 VTAIL.n462 VTAIL.n461 9.3005
R594 VTAIL.n464 VTAIL.n463 9.3005
R595 VTAIL.n442 VTAIL.n441 9.3005
R596 VTAIL.n470 VTAIL.n469 9.3005
R597 VTAIL.n472 VTAIL.n471 9.3005
R598 VTAIL.n495 VTAIL.n494 9.3005
R599 VTAIL.n430 VTAIL.n429 9.3005
R600 VTAIL.n489 VTAIL.n488 9.3005
R601 VTAIL.n487 VTAIL.n486 9.3005
R602 VTAIL.n434 VTAIL.n433 9.3005
R603 VTAIL.n481 VTAIL.n480 9.3005
R604 VTAIL.n479 VTAIL.n478 9.3005
R605 VTAIL.n438 VTAIL.n437 9.3005
R606 VTAIL.n382 VTAIL.n381 9.3005
R607 VTAIL.n384 VTAIL.n383 9.3005
R608 VTAIL.n375 VTAIL.n374 9.3005
R609 VTAIL.n390 VTAIL.n389 9.3005
R610 VTAIL.n392 VTAIL.n391 9.3005
R611 VTAIL.n370 VTAIL.n369 9.3005
R612 VTAIL.n398 VTAIL.n397 9.3005
R613 VTAIL.n400 VTAIL.n399 9.3005
R614 VTAIL.n423 VTAIL.n422 9.3005
R615 VTAIL.n358 VTAIL.n357 9.3005
R616 VTAIL.n417 VTAIL.n416 9.3005
R617 VTAIL.n415 VTAIL.n414 9.3005
R618 VTAIL.n362 VTAIL.n361 9.3005
R619 VTAIL.n409 VTAIL.n408 9.3005
R620 VTAIL.n407 VTAIL.n406 9.3005
R621 VTAIL.n366 VTAIL.n365 9.3005
R622 VTAIL.n312 VTAIL.n311 9.3005
R623 VTAIL.n314 VTAIL.n313 9.3005
R624 VTAIL.n305 VTAIL.n304 9.3005
R625 VTAIL.n320 VTAIL.n319 9.3005
R626 VTAIL.n322 VTAIL.n321 9.3005
R627 VTAIL.n300 VTAIL.n299 9.3005
R628 VTAIL.n328 VTAIL.n327 9.3005
R629 VTAIL.n330 VTAIL.n329 9.3005
R630 VTAIL.n353 VTAIL.n352 9.3005
R631 VTAIL.n288 VTAIL.n287 9.3005
R632 VTAIL.n347 VTAIL.n346 9.3005
R633 VTAIL.n345 VTAIL.n344 9.3005
R634 VTAIL.n292 VTAIL.n291 9.3005
R635 VTAIL.n339 VTAIL.n338 9.3005
R636 VTAIL.n337 VTAIL.n336 9.3005
R637 VTAIL.n296 VTAIL.n295 9.3005
R638 VTAIL.n240 VTAIL.n239 9.3005
R639 VTAIL.n242 VTAIL.n241 9.3005
R640 VTAIL.n233 VTAIL.n232 9.3005
R641 VTAIL.n248 VTAIL.n247 9.3005
R642 VTAIL.n250 VTAIL.n249 9.3005
R643 VTAIL.n228 VTAIL.n227 9.3005
R644 VTAIL.n256 VTAIL.n255 9.3005
R645 VTAIL.n258 VTAIL.n257 9.3005
R646 VTAIL.n281 VTAIL.n280 9.3005
R647 VTAIL.n216 VTAIL.n215 9.3005
R648 VTAIL.n275 VTAIL.n274 9.3005
R649 VTAIL.n273 VTAIL.n272 9.3005
R650 VTAIL.n220 VTAIL.n219 9.3005
R651 VTAIL.n267 VTAIL.n266 9.3005
R652 VTAIL.n265 VTAIL.n264 9.3005
R653 VTAIL.n224 VTAIL.n223 9.3005
R654 VTAIL.n526 VTAIL.n516 8.92171
R655 VTAIL.n560 VTAIL.n559 8.92171
R656 VTAIL.n30 VTAIL.n20 8.92171
R657 VTAIL.n64 VTAIL.n63 8.92171
R658 VTAIL.n100 VTAIL.n90 8.92171
R659 VTAIL.n134 VTAIL.n133 8.92171
R660 VTAIL.n172 VTAIL.n162 8.92171
R661 VTAIL.n206 VTAIL.n205 8.92171
R662 VTAIL.n490 VTAIL.n489 8.92171
R663 VTAIL.n457 VTAIL.n447 8.92171
R664 VTAIL.n418 VTAIL.n417 8.92171
R665 VTAIL.n385 VTAIL.n375 8.92171
R666 VTAIL.n348 VTAIL.n347 8.92171
R667 VTAIL.n315 VTAIL.n305 8.92171
R668 VTAIL.n276 VTAIL.n275 8.92171
R669 VTAIL.n243 VTAIL.n233 8.92171
R670 VTAIL.n525 VTAIL.n518 8.14595
R671 VTAIL.n563 VTAIL.n500 8.14595
R672 VTAIL.n29 VTAIL.n22 8.14595
R673 VTAIL.n67 VTAIL.n4 8.14595
R674 VTAIL.n99 VTAIL.n92 8.14595
R675 VTAIL.n137 VTAIL.n74 8.14595
R676 VTAIL.n171 VTAIL.n164 8.14595
R677 VTAIL.n209 VTAIL.n146 8.14595
R678 VTAIL.n493 VTAIL.n430 8.14595
R679 VTAIL.n456 VTAIL.n449 8.14595
R680 VTAIL.n421 VTAIL.n358 8.14595
R681 VTAIL.n384 VTAIL.n377 8.14595
R682 VTAIL.n351 VTAIL.n288 8.14595
R683 VTAIL.n314 VTAIL.n307 8.14595
R684 VTAIL.n279 VTAIL.n216 8.14595
R685 VTAIL.n242 VTAIL.n235 8.14595
R686 VTAIL.n522 VTAIL.n521 7.3702
R687 VTAIL.n564 VTAIL.n498 7.3702
R688 VTAIL.n26 VTAIL.n25 7.3702
R689 VTAIL.n68 VTAIL.n2 7.3702
R690 VTAIL.n96 VTAIL.n95 7.3702
R691 VTAIL.n138 VTAIL.n72 7.3702
R692 VTAIL.n168 VTAIL.n167 7.3702
R693 VTAIL.n210 VTAIL.n144 7.3702
R694 VTAIL.n494 VTAIL.n428 7.3702
R695 VTAIL.n453 VTAIL.n452 7.3702
R696 VTAIL.n422 VTAIL.n356 7.3702
R697 VTAIL.n381 VTAIL.n380 7.3702
R698 VTAIL.n352 VTAIL.n286 7.3702
R699 VTAIL.n311 VTAIL.n310 7.3702
R700 VTAIL.n280 VTAIL.n214 7.3702
R701 VTAIL.n239 VTAIL.n238 7.3702
R702 VTAIL.n566 VTAIL.n498 6.59444
R703 VTAIL.n70 VTAIL.n2 6.59444
R704 VTAIL.n140 VTAIL.n72 6.59444
R705 VTAIL.n212 VTAIL.n144 6.59444
R706 VTAIL.n496 VTAIL.n428 6.59444
R707 VTAIL.n424 VTAIL.n356 6.59444
R708 VTAIL.n354 VTAIL.n286 6.59444
R709 VTAIL.n282 VTAIL.n214 6.59444
R710 VTAIL.n522 VTAIL.n518 5.81868
R711 VTAIL.n564 VTAIL.n563 5.81868
R712 VTAIL.n26 VTAIL.n22 5.81868
R713 VTAIL.n68 VTAIL.n67 5.81868
R714 VTAIL.n96 VTAIL.n92 5.81868
R715 VTAIL.n138 VTAIL.n137 5.81868
R716 VTAIL.n168 VTAIL.n164 5.81868
R717 VTAIL.n210 VTAIL.n209 5.81868
R718 VTAIL.n494 VTAIL.n493 5.81868
R719 VTAIL.n453 VTAIL.n449 5.81868
R720 VTAIL.n422 VTAIL.n421 5.81868
R721 VTAIL.n381 VTAIL.n377 5.81868
R722 VTAIL.n352 VTAIL.n351 5.81868
R723 VTAIL.n311 VTAIL.n307 5.81868
R724 VTAIL.n280 VTAIL.n279 5.81868
R725 VTAIL.n239 VTAIL.n235 5.81868
R726 VTAIL.n526 VTAIL.n525 5.04292
R727 VTAIL.n560 VTAIL.n500 5.04292
R728 VTAIL.n30 VTAIL.n29 5.04292
R729 VTAIL.n64 VTAIL.n4 5.04292
R730 VTAIL.n100 VTAIL.n99 5.04292
R731 VTAIL.n134 VTAIL.n74 5.04292
R732 VTAIL.n172 VTAIL.n171 5.04292
R733 VTAIL.n206 VTAIL.n146 5.04292
R734 VTAIL.n490 VTAIL.n430 5.04292
R735 VTAIL.n457 VTAIL.n456 5.04292
R736 VTAIL.n418 VTAIL.n358 5.04292
R737 VTAIL.n385 VTAIL.n384 5.04292
R738 VTAIL.n348 VTAIL.n288 5.04292
R739 VTAIL.n315 VTAIL.n314 5.04292
R740 VTAIL.n276 VTAIL.n216 5.04292
R741 VTAIL.n243 VTAIL.n242 5.04292
R742 VTAIL.n529 VTAIL.n516 4.26717
R743 VTAIL.n559 VTAIL.n502 4.26717
R744 VTAIL.n33 VTAIL.n20 4.26717
R745 VTAIL.n63 VTAIL.n6 4.26717
R746 VTAIL.n103 VTAIL.n90 4.26717
R747 VTAIL.n133 VTAIL.n76 4.26717
R748 VTAIL.n175 VTAIL.n162 4.26717
R749 VTAIL.n205 VTAIL.n148 4.26717
R750 VTAIL.n489 VTAIL.n432 4.26717
R751 VTAIL.n460 VTAIL.n447 4.26717
R752 VTAIL.n417 VTAIL.n360 4.26717
R753 VTAIL.n388 VTAIL.n375 4.26717
R754 VTAIL.n347 VTAIL.n290 4.26717
R755 VTAIL.n318 VTAIL.n305 4.26717
R756 VTAIL.n275 VTAIL.n218 4.26717
R757 VTAIL.n246 VTAIL.n233 4.26717
R758 VTAIL.n530 VTAIL.n514 3.49141
R759 VTAIL.n556 VTAIL.n555 3.49141
R760 VTAIL.n34 VTAIL.n18 3.49141
R761 VTAIL.n60 VTAIL.n59 3.49141
R762 VTAIL.n104 VTAIL.n88 3.49141
R763 VTAIL.n130 VTAIL.n129 3.49141
R764 VTAIL.n176 VTAIL.n160 3.49141
R765 VTAIL.n202 VTAIL.n201 3.49141
R766 VTAIL.n486 VTAIL.n485 3.49141
R767 VTAIL.n461 VTAIL.n445 3.49141
R768 VTAIL.n414 VTAIL.n413 3.49141
R769 VTAIL.n389 VTAIL.n373 3.49141
R770 VTAIL.n344 VTAIL.n343 3.49141
R771 VTAIL.n319 VTAIL.n303 3.49141
R772 VTAIL.n272 VTAIL.n271 3.49141
R773 VTAIL.n247 VTAIL.n231 3.49141
R774 VTAIL.n285 VTAIL.n283 2.77636
R775 VTAIL.n355 VTAIL.n285 2.77636
R776 VTAIL.n427 VTAIL.n425 2.77636
R777 VTAIL.n497 VTAIL.n427 2.77636
R778 VTAIL.n213 VTAIL.n143 2.77636
R779 VTAIL.n143 VTAIL.n141 2.77636
R780 VTAIL.n71 VTAIL.n1 2.77636
R781 VTAIL VTAIL.n567 2.71817
R782 VTAIL.n534 VTAIL.n533 2.71565
R783 VTAIL.n552 VTAIL.n504 2.71565
R784 VTAIL.n38 VTAIL.n37 2.71565
R785 VTAIL.n56 VTAIL.n8 2.71565
R786 VTAIL.n108 VTAIL.n107 2.71565
R787 VTAIL.n126 VTAIL.n78 2.71565
R788 VTAIL.n180 VTAIL.n179 2.71565
R789 VTAIL.n198 VTAIL.n150 2.71565
R790 VTAIL.n482 VTAIL.n434 2.71565
R791 VTAIL.n465 VTAIL.n464 2.71565
R792 VTAIL.n410 VTAIL.n362 2.71565
R793 VTAIL.n393 VTAIL.n392 2.71565
R794 VTAIL.n340 VTAIL.n292 2.71565
R795 VTAIL.n323 VTAIL.n322 2.71565
R796 VTAIL.n268 VTAIL.n220 2.71565
R797 VTAIL.n251 VTAIL.n250 2.71565
R798 VTAIL.n0 VTAIL.t7 2.55592
R799 VTAIL.n0 VTAIL.t0 2.55592
R800 VTAIL.n142 VTAIL.t12 2.55592
R801 VTAIL.n142 VTAIL.t13 2.55592
R802 VTAIL.n426 VTAIL.t14 2.55592
R803 VTAIL.n426 VTAIL.t15 2.55592
R804 VTAIL.n284 VTAIL.t4 2.55592
R805 VTAIL.n284 VTAIL.t6 2.55592
R806 VTAIL.n523 VTAIL.n519 2.41282
R807 VTAIL.n27 VTAIL.n23 2.41282
R808 VTAIL.n97 VTAIL.n93 2.41282
R809 VTAIL.n169 VTAIL.n165 2.41282
R810 VTAIL.n454 VTAIL.n450 2.41282
R811 VTAIL.n382 VTAIL.n378 2.41282
R812 VTAIL.n312 VTAIL.n308 2.41282
R813 VTAIL.n240 VTAIL.n236 2.41282
R814 VTAIL.n538 VTAIL.n512 1.93989
R815 VTAIL.n551 VTAIL.n506 1.93989
R816 VTAIL.n42 VTAIL.n16 1.93989
R817 VTAIL.n55 VTAIL.n10 1.93989
R818 VTAIL.n112 VTAIL.n86 1.93989
R819 VTAIL.n125 VTAIL.n80 1.93989
R820 VTAIL.n184 VTAIL.n158 1.93989
R821 VTAIL.n197 VTAIL.n152 1.93989
R822 VTAIL.n481 VTAIL.n436 1.93989
R823 VTAIL.n468 VTAIL.n442 1.93989
R824 VTAIL.n409 VTAIL.n364 1.93989
R825 VTAIL.n396 VTAIL.n370 1.93989
R826 VTAIL.n339 VTAIL.n294 1.93989
R827 VTAIL.n326 VTAIL.n300 1.93989
R828 VTAIL.n267 VTAIL.n222 1.93989
R829 VTAIL.n254 VTAIL.n228 1.93989
R830 VTAIL.n539 VTAIL.n510 1.16414
R831 VTAIL.n548 VTAIL.n547 1.16414
R832 VTAIL.n43 VTAIL.n14 1.16414
R833 VTAIL.n52 VTAIL.n51 1.16414
R834 VTAIL.n113 VTAIL.n84 1.16414
R835 VTAIL.n122 VTAIL.n121 1.16414
R836 VTAIL.n185 VTAIL.n156 1.16414
R837 VTAIL.n194 VTAIL.n193 1.16414
R838 VTAIL.n478 VTAIL.n477 1.16414
R839 VTAIL.n469 VTAIL.n440 1.16414
R840 VTAIL.n406 VTAIL.n405 1.16414
R841 VTAIL.n397 VTAIL.n368 1.16414
R842 VTAIL.n336 VTAIL.n335 1.16414
R843 VTAIL.n327 VTAIL.n298 1.16414
R844 VTAIL.n264 VTAIL.n263 1.16414
R845 VTAIL.n255 VTAIL.n226 1.16414
R846 VTAIL.n425 VTAIL.n355 0.470328
R847 VTAIL.n141 VTAIL.n71 0.470328
R848 VTAIL.n543 VTAIL.n542 0.388379
R849 VTAIL.n544 VTAIL.n508 0.388379
R850 VTAIL.n47 VTAIL.n46 0.388379
R851 VTAIL.n48 VTAIL.n12 0.388379
R852 VTAIL.n117 VTAIL.n116 0.388379
R853 VTAIL.n118 VTAIL.n82 0.388379
R854 VTAIL.n189 VTAIL.n188 0.388379
R855 VTAIL.n190 VTAIL.n154 0.388379
R856 VTAIL.n474 VTAIL.n438 0.388379
R857 VTAIL.n473 VTAIL.n472 0.388379
R858 VTAIL.n402 VTAIL.n366 0.388379
R859 VTAIL.n401 VTAIL.n400 0.388379
R860 VTAIL.n332 VTAIL.n296 0.388379
R861 VTAIL.n331 VTAIL.n330 0.388379
R862 VTAIL.n260 VTAIL.n224 0.388379
R863 VTAIL.n259 VTAIL.n258 0.388379
R864 VTAIL.n524 VTAIL.n523 0.155672
R865 VTAIL.n524 VTAIL.n515 0.155672
R866 VTAIL.n531 VTAIL.n515 0.155672
R867 VTAIL.n532 VTAIL.n531 0.155672
R868 VTAIL.n532 VTAIL.n511 0.155672
R869 VTAIL.n540 VTAIL.n511 0.155672
R870 VTAIL.n541 VTAIL.n540 0.155672
R871 VTAIL.n541 VTAIL.n507 0.155672
R872 VTAIL.n549 VTAIL.n507 0.155672
R873 VTAIL.n550 VTAIL.n549 0.155672
R874 VTAIL.n550 VTAIL.n503 0.155672
R875 VTAIL.n557 VTAIL.n503 0.155672
R876 VTAIL.n558 VTAIL.n557 0.155672
R877 VTAIL.n558 VTAIL.n499 0.155672
R878 VTAIL.n565 VTAIL.n499 0.155672
R879 VTAIL.n28 VTAIL.n27 0.155672
R880 VTAIL.n28 VTAIL.n19 0.155672
R881 VTAIL.n35 VTAIL.n19 0.155672
R882 VTAIL.n36 VTAIL.n35 0.155672
R883 VTAIL.n36 VTAIL.n15 0.155672
R884 VTAIL.n44 VTAIL.n15 0.155672
R885 VTAIL.n45 VTAIL.n44 0.155672
R886 VTAIL.n45 VTAIL.n11 0.155672
R887 VTAIL.n53 VTAIL.n11 0.155672
R888 VTAIL.n54 VTAIL.n53 0.155672
R889 VTAIL.n54 VTAIL.n7 0.155672
R890 VTAIL.n61 VTAIL.n7 0.155672
R891 VTAIL.n62 VTAIL.n61 0.155672
R892 VTAIL.n62 VTAIL.n3 0.155672
R893 VTAIL.n69 VTAIL.n3 0.155672
R894 VTAIL.n98 VTAIL.n97 0.155672
R895 VTAIL.n98 VTAIL.n89 0.155672
R896 VTAIL.n105 VTAIL.n89 0.155672
R897 VTAIL.n106 VTAIL.n105 0.155672
R898 VTAIL.n106 VTAIL.n85 0.155672
R899 VTAIL.n114 VTAIL.n85 0.155672
R900 VTAIL.n115 VTAIL.n114 0.155672
R901 VTAIL.n115 VTAIL.n81 0.155672
R902 VTAIL.n123 VTAIL.n81 0.155672
R903 VTAIL.n124 VTAIL.n123 0.155672
R904 VTAIL.n124 VTAIL.n77 0.155672
R905 VTAIL.n131 VTAIL.n77 0.155672
R906 VTAIL.n132 VTAIL.n131 0.155672
R907 VTAIL.n132 VTAIL.n73 0.155672
R908 VTAIL.n139 VTAIL.n73 0.155672
R909 VTAIL.n170 VTAIL.n169 0.155672
R910 VTAIL.n170 VTAIL.n161 0.155672
R911 VTAIL.n177 VTAIL.n161 0.155672
R912 VTAIL.n178 VTAIL.n177 0.155672
R913 VTAIL.n178 VTAIL.n157 0.155672
R914 VTAIL.n186 VTAIL.n157 0.155672
R915 VTAIL.n187 VTAIL.n186 0.155672
R916 VTAIL.n187 VTAIL.n153 0.155672
R917 VTAIL.n195 VTAIL.n153 0.155672
R918 VTAIL.n196 VTAIL.n195 0.155672
R919 VTAIL.n196 VTAIL.n149 0.155672
R920 VTAIL.n203 VTAIL.n149 0.155672
R921 VTAIL.n204 VTAIL.n203 0.155672
R922 VTAIL.n204 VTAIL.n145 0.155672
R923 VTAIL.n211 VTAIL.n145 0.155672
R924 VTAIL.n495 VTAIL.n429 0.155672
R925 VTAIL.n488 VTAIL.n429 0.155672
R926 VTAIL.n488 VTAIL.n487 0.155672
R927 VTAIL.n487 VTAIL.n433 0.155672
R928 VTAIL.n480 VTAIL.n433 0.155672
R929 VTAIL.n480 VTAIL.n479 0.155672
R930 VTAIL.n479 VTAIL.n437 0.155672
R931 VTAIL.n471 VTAIL.n437 0.155672
R932 VTAIL.n471 VTAIL.n470 0.155672
R933 VTAIL.n470 VTAIL.n441 0.155672
R934 VTAIL.n463 VTAIL.n441 0.155672
R935 VTAIL.n463 VTAIL.n462 0.155672
R936 VTAIL.n462 VTAIL.n446 0.155672
R937 VTAIL.n455 VTAIL.n446 0.155672
R938 VTAIL.n455 VTAIL.n454 0.155672
R939 VTAIL.n423 VTAIL.n357 0.155672
R940 VTAIL.n416 VTAIL.n357 0.155672
R941 VTAIL.n416 VTAIL.n415 0.155672
R942 VTAIL.n415 VTAIL.n361 0.155672
R943 VTAIL.n408 VTAIL.n361 0.155672
R944 VTAIL.n408 VTAIL.n407 0.155672
R945 VTAIL.n407 VTAIL.n365 0.155672
R946 VTAIL.n399 VTAIL.n365 0.155672
R947 VTAIL.n399 VTAIL.n398 0.155672
R948 VTAIL.n398 VTAIL.n369 0.155672
R949 VTAIL.n391 VTAIL.n369 0.155672
R950 VTAIL.n391 VTAIL.n390 0.155672
R951 VTAIL.n390 VTAIL.n374 0.155672
R952 VTAIL.n383 VTAIL.n374 0.155672
R953 VTAIL.n383 VTAIL.n382 0.155672
R954 VTAIL.n353 VTAIL.n287 0.155672
R955 VTAIL.n346 VTAIL.n287 0.155672
R956 VTAIL.n346 VTAIL.n345 0.155672
R957 VTAIL.n345 VTAIL.n291 0.155672
R958 VTAIL.n338 VTAIL.n291 0.155672
R959 VTAIL.n338 VTAIL.n337 0.155672
R960 VTAIL.n337 VTAIL.n295 0.155672
R961 VTAIL.n329 VTAIL.n295 0.155672
R962 VTAIL.n329 VTAIL.n328 0.155672
R963 VTAIL.n328 VTAIL.n299 0.155672
R964 VTAIL.n321 VTAIL.n299 0.155672
R965 VTAIL.n321 VTAIL.n320 0.155672
R966 VTAIL.n320 VTAIL.n304 0.155672
R967 VTAIL.n313 VTAIL.n304 0.155672
R968 VTAIL.n313 VTAIL.n312 0.155672
R969 VTAIL.n281 VTAIL.n215 0.155672
R970 VTAIL.n274 VTAIL.n215 0.155672
R971 VTAIL.n274 VTAIL.n273 0.155672
R972 VTAIL.n273 VTAIL.n219 0.155672
R973 VTAIL.n266 VTAIL.n219 0.155672
R974 VTAIL.n266 VTAIL.n265 0.155672
R975 VTAIL.n265 VTAIL.n223 0.155672
R976 VTAIL.n257 VTAIL.n223 0.155672
R977 VTAIL.n257 VTAIL.n256 0.155672
R978 VTAIL.n256 VTAIL.n227 0.155672
R979 VTAIL.n249 VTAIL.n227 0.155672
R980 VTAIL.n249 VTAIL.n248 0.155672
R981 VTAIL.n248 VTAIL.n232 0.155672
R982 VTAIL.n241 VTAIL.n232 0.155672
R983 VTAIL.n241 VTAIL.n240 0.155672
R984 VTAIL VTAIL.n1 0.0586897
R985 VDD1 VDD1.n0 72.1302
R986 VDD1.n3 VDD1.n2 72.0167
R987 VDD1.n3 VDD1.n1 72.0167
R988 VDD1.n5 VDD1.n4 70.6839
R989 VDD1.n5 VDD1.n3 47.7552
R990 VDD1.n4 VDD1.t4 2.55592
R991 VDD1.n4 VDD1.t5 2.55592
R992 VDD1.n0 VDD1.t1 2.55592
R993 VDD1.n0 VDD1.t3 2.55592
R994 VDD1.n2 VDD1.t0 2.55592
R995 VDD1.n2 VDD1.t2 2.55592
R996 VDD1.n1 VDD1.t6 2.55592
R997 VDD1.n1 VDD1.t7 2.55592
R998 VDD1 VDD1.n5 1.33024
R999 VN.n59 VN.n31 161.3
R1000 VN.n58 VN.n57 161.3
R1001 VN.n56 VN.n32 161.3
R1002 VN.n55 VN.n54 161.3
R1003 VN.n53 VN.n33 161.3
R1004 VN.n52 VN.n51 161.3
R1005 VN.n50 VN.n34 161.3
R1006 VN.n49 VN.n48 161.3
R1007 VN.n47 VN.n35 161.3
R1008 VN.n46 VN.n45 161.3
R1009 VN.n44 VN.n37 161.3
R1010 VN.n43 VN.n42 161.3
R1011 VN.n41 VN.n38 161.3
R1012 VN.n28 VN.n0 161.3
R1013 VN.n27 VN.n26 161.3
R1014 VN.n25 VN.n1 161.3
R1015 VN.n24 VN.n23 161.3
R1016 VN.n22 VN.n2 161.3
R1017 VN.n21 VN.n20 161.3
R1018 VN.n19 VN.n3 161.3
R1019 VN.n18 VN.n17 161.3
R1020 VN.n15 VN.n4 161.3
R1021 VN.n14 VN.n13 161.3
R1022 VN.n12 VN.n5 161.3
R1023 VN.n11 VN.n10 161.3
R1024 VN.n9 VN.n6 161.3
R1025 VN.n7 VN.t7 139.519
R1026 VN.n39 VN.t4 139.519
R1027 VN.n30 VN.n29 106.712
R1028 VN.n61 VN.n60 106.712
R1029 VN.n8 VN.t6 106.073
R1030 VN.n16 VN.t0 106.073
R1031 VN.n29 VN.t2 106.073
R1032 VN.n40 VN.t3 106.073
R1033 VN.n36 VN.t5 106.073
R1034 VN.n60 VN.t1 106.073
R1035 VN.n14 VN.n5 56.4773
R1036 VN.n46 VN.n37 56.4773
R1037 VN.n8 VN.n7 55.9247
R1038 VN.n40 VN.n39 55.9247
R1039 VN VN.n61 53.0739
R1040 VN.n23 VN.n22 43.3318
R1041 VN.n54 VN.n53 43.3318
R1042 VN.n23 VN.n1 37.4894
R1043 VN.n54 VN.n32 37.4894
R1044 VN.n10 VN.n9 24.3439
R1045 VN.n10 VN.n5 24.3439
R1046 VN.n15 VN.n14 24.3439
R1047 VN.n17 VN.n15 24.3439
R1048 VN.n21 VN.n3 24.3439
R1049 VN.n22 VN.n21 24.3439
R1050 VN.n27 VN.n1 24.3439
R1051 VN.n28 VN.n27 24.3439
R1052 VN.n42 VN.n37 24.3439
R1053 VN.n42 VN.n41 24.3439
R1054 VN.n53 VN.n52 24.3439
R1055 VN.n52 VN.n34 24.3439
R1056 VN.n48 VN.n47 24.3439
R1057 VN.n47 VN.n46 24.3439
R1058 VN.n59 VN.n58 24.3439
R1059 VN.n58 VN.n32 24.3439
R1060 VN.n9 VN.n8 17.5278
R1061 VN.n17 VN.n16 17.5278
R1062 VN.n41 VN.n40 17.5278
R1063 VN.n48 VN.n36 17.5278
R1064 VN.n16 VN.n3 6.81666
R1065 VN.n36 VN.n34 6.81666
R1066 VN.n39 VN.n38 5.04473
R1067 VN.n7 VN.n6 5.04473
R1068 VN.n29 VN.n28 3.89545
R1069 VN.n60 VN.n59 3.89545
R1070 VN.n61 VN.n31 0.278398
R1071 VN.n30 VN.n0 0.278398
R1072 VN.n57 VN.n31 0.189894
R1073 VN.n57 VN.n56 0.189894
R1074 VN.n56 VN.n55 0.189894
R1075 VN.n55 VN.n33 0.189894
R1076 VN.n51 VN.n33 0.189894
R1077 VN.n51 VN.n50 0.189894
R1078 VN.n50 VN.n49 0.189894
R1079 VN.n49 VN.n35 0.189894
R1080 VN.n45 VN.n35 0.189894
R1081 VN.n45 VN.n44 0.189894
R1082 VN.n44 VN.n43 0.189894
R1083 VN.n43 VN.n38 0.189894
R1084 VN.n11 VN.n6 0.189894
R1085 VN.n12 VN.n11 0.189894
R1086 VN.n13 VN.n12 0.189894
R1087 VN.n13 VN.n4 0.189894
R1088 VN.n18 VN.n4 0.189894
R1089 VN.n19 VN.n18 0.189894
R1090 VN.n20 VN.n19 0.189894
R1091 VN.n20 VN.n2 0.189894
R1092 VN.n24 VN.n2 0.189894
R1093 VN.n25 VN.n24 0.189894
R1094 VN.n26 VN.n25 0.189894
R1095 VN.n26 VN.n0 0.189894
R1096 VN VN.n30 0.153422
R1097 VDD2.n2 VDD2.n1 72.0167
R1098 VDD2.n2 VDD2.n0 72.0167
R1099 VDD2 VDD2.n5 72.0136
R1100 VDD2.n4 VDD2.n3 70.6841
R1101 VDD2.n4 VDD2.n2 47.1722
R1102 VDD2.n5 VDD2.t4 2.55592
R1103 VDD2.n5 VDD2.t3 2.55592
R1104 VDD2.n3 VDD2.t6 2.55592
R1105 VDD2.n3 VDD2.t2 2.55592
R1106 VDD2.n1 VDD2.t7 2.55592
R1107 VDD2.n1 VDD2.t5 2.55592
R1108 VDD2.n0 VDD2.t0 2.55592
R1109 VDD2.n0 VDD2.t1 2.55592
R1110 VDD2 VDD2.n4 1.44662
R1111 B.n446 B.n445 585
R1112 B.n444 B.n139 585
R1113 B.n443 B.n442 585
R1114 B.n441 B.n140 585
R1115 B.n440 B.n439 585
R1116 B.n438 B.n141 585
R1117 B.n437 B.n436 585
R1118 B.n435 B.n142 585
R1119 B.n434 B.n433 585
R1120 B.n432 B.n143 585
R1121 B.n431 B.n430 585
R1122 B.n429 B.n144 585
R1123 B.n428 B.n427 585
R1124 B.n426 B.n145 585
R1125 B.n425 B.n424 585
R1126 B.n423 B.n146 585
R1127 B.n422 B.n421 585
R1128 B.n420 B.n147 585
R1129 B.n419 B.n418 585
R1130 B.n417 B.n148 585
R1131 B.n416 B.n415 585
R1132 B.n414 B.n149 585
R1133 B.n413 B.n412 585
R1134 B.n411 B.n150 585
R1135 B.n410 B.n409 585
R1136 B.n408 B.n151 585
R1137 B.n407 B.n406 585
R1138 B.n405 B.n152 585
R1139 B.n404 B.n403 585
R1140 B.n402 B.n153 585
R1141 B.n401 B.n400 585
R1142 B.n399 B.n154 585
R1143 B.n398 B.n397 585
R1144 B.n396 B.n155 585
R1145 B.n395 B.n394 585
R1146 B.n393 B.n156 585
R1147 B.n392 B.n391 585
R1148 B.n390 B.n157 585
R1149 B.n389 B.n388 585
R1150 B.n387 B.n158 585
R1151 B.n386 B.n385 585
R1152 B.n384 B.n159 585
R1153 B.n383 B.n382 585
R1154 B.n381 B.n160 585
R1155 B.n380 B.n379 585
R1156 B.n375 B.n161 585
R1157 B.n374 B.n373 585
R1158 B.n372 B.n162 585
R1159 B.n371 B.n370 585
R1160 B.n369 B.n163 585
R1161 B.n368 B.n367 585
R1162 B.n366 B.n164 585
R1163 B.n365 B.n364 585
R1164 B.n362 B.n165 585
R1165 B.n361 B.n360 585
R1166 B.n359 B.n168 585
R1167 B.n358 B.n357 585
R1168 B.n356 B.n169 585
R1169 B.n355 B.n354 585
R1170 B.n353 B.n170 585
R1171 B.n352 B.n351 585
R1172 B.n350 B.n171 585
R1173 B.n349 B.n348 585
R1174 B.n347 B.n172 585
R1175 B.n346 B.n345 585
R1176 B.n344 B.n173 585
R1177 B.n343 B.n342 585
R1178 B.n341 B.n174 585
R1179 B.n340 B.n339 585
R1180 B.n338 B.n175 585
R1181 B.n337 B.n336 585
R1182 B.n335 B.n176 585
R1183 B.n334 B.n333 585
R1184 B.n332 B.n177 585
R1185 B.n331 B.n330 585
R1186 B.n329 B.n178 585
R1187 B.n328 B.n327 585
R1188 B.n326 B.n179 585
R1189 B.n325 B.n324 585
R1190 B.n323 B.n180 585
R1191 B.n322 B.n321 585
R1192 B.n320 B.n181 585
R1193 B.n319 B.n318 585
R1194 B.n317 B.n182 585
R1195 B.n316 B.n315 585
R1196 B.n314 B.n183 585
R1197 B.n313 B.n312 585
R1198 B.n311 B.n184 585
R1199 B.n310 B.n309 585
R1200 B.n308 B.n185 585
R1201 B.n307 B.n306 585
R1202 B.n305 B.n186 585
R1203 B.n304 B.n303 585
R1204 B.n302 B.n187 585
R1205 B.n301 B.n300 585
R1206 B.n299 B.n188 585
R1207 B.n298 B.n297 585
R1208 B.n447 B.n138 585
R1209 B.n449 B.n448 585
R1210 B.n450 B.n137 585
R1211 B.n452 B.n451 585
R1212 B.n453 B.n136 585
R1213 B.n455 B.n454 585
R1214 B.n456 B.n135 585
R1215 B.n458 B.n457 585
R1216 B.n459 B.n134 585
R1217 B.n461 B.n460 585
R1218 B.n462 B.n133 585
R1219 B.n464 B.n463 585
R1220 B.n465 B.n132 585
R1221 B.n467 B.n466 585
R1222 B.n468 B.n131 585
R1223 B.n470 B.n469 585
R1224 B.n471 B.n130 585
R1225 B.n473 B.n472 585
R1226 B.n474 B.n129 585
R1227 B.n476 B.n475 585
R1228 B.n477 B.n128 585
R1229 B.n479 B.n478 585
R1230 B.n480 B.n127 585
R1231 B.n482 B.n481 585
R1232 B.n483 B.n126 585
R1233 B.n485 B.n484 585
R1234 B.n486 B.n125 585
R1235 B.n488 B.n487 585
R1236 B.n489 B.n124 585
R1237 B.n491 B.n490 585
R1238 B.n492 B.n123 585
R1239 B.n494 B.n493 585
R1240 B.n495 B.n122 585
R1241 B.n497 B.n496 585
R1242 B.n498 B.n121 585
R1243 B.n500 B.n499 585
R1244 B.n501 B.n120 585
R1245 B.n503 B.n502 585
R1246 B.n504 B.n119 585
R1247 B.n506 B.n505 585
R1248 B.n507 B.n118 585
R1249 B.n509 B.n508 585
R1250 B.n510 B.n117 585
R1251 B.n512 B.n511 585
R1252 B.n513 B.n116 585
R1253 B.n515 B.n514 585
R1254 B.n516 B.n115 585
R1255 B.n518 B.n517 585
R1256 B.n519 B.n114 585
R1257 B.n521 B.n520 585
R1258 B.n522 B.n113 585
R1259 B.n524 B.n523 585
R1260 B.n525 B.n112 585
R1261 B.n527 B.n526 585
R1262 B.n528 B.n111 585
R1263 B.n530 B.n529 585
R1264 B.n531 B.n110 585
R1265 B.n533 B.n532 585
R1266 B.n534 B.n109 585
R1267 B.n536 B.n535 585
R1268 B.n537 B.n108 585
R1269 B.n539 B.n538 585
R1270 B.n540 B.n107 585
R1271 B.n542 B.n541 585
R1272 B.n543 B.n106 585
R1273 B.n545 B.n544 585
R1274 B.n546 B.n105 585
R1275 B.n548 B.n547 585
R1276 B.n549 B.n104 585
R1277 B.n551 B.n550 585
R1278 B.n552 B.n103 585
R1279 B.n554 B.n553 585
R1280 B.n555 B.n102 585
R1281 B.n557 B.n556 585
R1282 B.n558 B.n101 585
R1283 B.n560 B.n559 585
R1284 B.n561 B.n100 585
R1285 B.n563 B.n562 585
R1286 B.n564 B.n99 585
R1287 B.n566 B.n565 585
R1288 B.n567 B.n98 585
R1289 B.n569 B.n568 585
R1290 B.n570 B.n97 585
R1291 B.n572 B.n571 585
R1292 B.n573 B.n96 585
R1293 B.n575 B.n574 585
R1294 B.n576 B.n95 585
R1295 B.n578 B.n577 585
R1296 B.n579 B.n94 585
R1297 B.n581 B.n580 585
R1298 B.n582 B.n93 585
R1299 B.n584 B.n583 585
R1300 B.n585 B.n92 585
R1301 B.n587 B.n586 585
R1302 B.n588 B.n91 585
R1303 B.n590 B.n589 585
R1304 B.n591 B.n90 585
R1305 B.n593 B.n592 585
R1306 B.n594 B.n89 585
R1307 B.n596 B.n595 585
R1308 B.n597 B.n88 585
R1309 B.n599 B.n598 585
R1310 B.n600 B.n87 585
R1311 B.n602 B.n601 585
R1312 B.n603 B.n86 585
R1313 B.n605 B.n604 585
R1314 B.n606 B.n85 585
R1315 B.n608 B.n607 585
R1316 B.n609 B.n84 585
R1317 B.n611 B.n610 585
R1318 B.n612 B.n83 585
R1319 B.n614 B.n613 585
R1320 B.n761 B.n760 585
R1321 B.n759 B.n30 585
R1322 B.n758 B.n757 585
R1323 B.n756 B.n31 585
R1324 B.n755 B.n754 585
R1325 B.n753 B.n32 585
R1326 B.n752 B.n751 585
R1327 B.n750 B.n33 585
R1328 B.n749 B.n748 585
R1329 B.n747 B.n34 585
R1330 B.n746 B.n745 585
R1331 B.n744 B.n35 585
R1332 B.n743 B.n742 585
R1333 B.n741 B.n36 585
R1334 B.n740 B.n739 585
R1335 B.n738 B.n37 585
R1336 B.n737 B.n736 585
R1337 B.n735 B.n38 585
R1338 B.n734 B.n733 585
R1339 B.n732 B.n39 585
R1340 B.n731 B.n730 585
R1341 B.n729 B.n40 585
R1342 B.n728 B.n727 585
R1343 B.n726 B.n41 585
R1344 B.n725 B.n724 585
R1345 B.n723 B.n42 585
R1346 B.n722 B.n721 585
R1347 B.n720 B.n43 585
R1348 B.n719 B.n718 585
R1349 B.n717 B.n44 585
R1350 B.n716 B.n715 585
R1351 B.n714 B.n45 585
R1352 B.n713 B.n712 585
R1353 B.n711 B.n46 585
R1354 B.n710 B.n709 585
R1355 B.n708 B.n47 585
R1356 B.n707 B.n706 585
R1357 B.n705 B.n48 585
R1358 B.n704 B.n703 585
R1359 B.n702 B.n49 585
R1360 B.n701 B.n700 585
R1361 B.n699 B.n50 585
R1362 B.n698 B.n697 585
R1363 B.n696 B.n51 585
R1364 B.n694 B.n693 585
R1365 B.n692 B.n54 585
R1366 B.n691 B.n690 585
R1367 B.n689 B.n55 585
R1368 B.n688 B.n687 585
R1369 B.n686 B.n56 585
R1370 B.n685 B.n684 585
R1371 B.n683 B.n57 585
R1372 B.n682 B.n681 585
R1373 B.n680 B.n679 585
R1374 B.n678 B.n61 585
R1375 B.n677 B.n676 585
R1376 B.n675 B.n62 585
R1377 B.n674 B.n673 585
R1378 B.n672 B.n63 585
R1379 B.n671 B.n670 585
R1380 B.n669 B.n64 585
R1381 B.n668 B.n667 585
R1382 B.n666 B.n65 585
R1383 B.n665 B.n664 585
R1384 B.n663 B.n66 585
R1385 B.n662 B.n661 585
R1386 B.n660 B.n67 585
R1387 B.n659 B.n658 585
R1388 B.n657 B.n68 585
R1389 B.n656 B.n655 585
R1390 B.n654 B.n69 585
R1391 B.n653 B.n652 585
R1392 B.n651 B.n70 585
R1393 B.n650 B.n649 585
R1394 B.n648 B.n71 585
R1395 B.n647 B.n646 585
R1396 B.n645 B.n72 585
R1397 B.n644 B.n643 585
R1398 B.n642 B.n73 585
R1399 B.n641 B.n640 585
R1400 B.n639 B.n74 585
R1401 B.n638 B.n637 585
R1402 B.n636 B.n75 585
R1403 B.n635 B.n634 585
R1404 B.n633 B.n76 585
R1405 B.n632 B.n631 585
R1406 B.n630 B.n77 585
R1407 B.n629 B.n628 585
R1408 B.n627 B.n78 585
R1409 B.n626 B.n625 585
R1410 B.n624 B.n79 585
R1411 B.n623 B.n622 585
R1412 B.n621 B.n80 585
R1413 B.n620 B.n619 585
R1414 B.n618 B.n81 585
R1415 B.n617 B.n616 585
R1416 B.n615 B.n82 585
R1417 B.n762 B.n29 585
R1418 B.n764 B.n763 585
R1419 B.n765 B.n28 585
R1420 B.n767 B.n766 585
R1421 B.n768 B.n27 585
R1422 B.n770 B.n769 585
R1423 B.n771 B.n26 585
R1424 B.n773 B.n772 585
R1425 B.n774 B.n25 585
R1426 B.n776 B.n775 585
R1427 B.n777 B.n24 585
R1428 B.n779 B.n778 585
R1429 B.n780 B.n23 585
R1430 B.n782 B.n781 585
R1431 B.n783 B.n22 585
R1432 B.n785 B.n784 585
R1433 B.n786 B.n21 585
R1434 B.n788 B.n787 585
R1435 B.n789 B.n20 585
R1436 B.n791 B.n790 585
R1437 B.n792 B.n19 585
R1438 B.n794 B.n793 585
R1439 B.n795 B.n18 585
R1440 B.n797 B.n796 585
R1441 B.n798 B.n17 585
R1442 B.n800 B.n799 585
R1443 B.n801 B.n16 585
R1444 B.n803 B.n802 585
R1445 B.n804 B.n15 585
R1446 B.n806 B.n805 585
R1447 B.n807 B.n14 585
R1448 B.n809 B.n808 585
R1449 B.n810 B.n13 585
R1450 B.n812 B.n811 585
R1451 B.n813 B.n12 585
R1452 B.n815 B.n814 585
R1453 B.n816 B.n11 585
R1454 B.n818 B.n817 585
R1455 B.n819 B.n10 585
R1456 B.n821 B.n820 585
R1457 B.n822 B.n9 585
R1458 B.n824 B.n823 585
R1459 B.n825 B.n8 585
R1460 B.n827 B.n826 585
R1461 B.n828 B.n7 585
R1462 B.n830 B.n829 585
R1463 B.n831 B.n6 585
R1464 B.n833 B.n832 585
R1465 B.n834 B.n5 585
R1466 B.n836 B.n835 585
R1467 B.n837 B.n4 585
R1468 B.n839 B.n838 585
R1469 B.n840 B.n3 585
R1470 B.n842 B.n841 585
R1471 B.n843 B.n0 585
R1472 B.n2 B.n1 585
R1473 B.n217 B.n216 585
R1474 B.n218 B.n215 585
R1475 B.n220 B.n219 585
R1476 B.n221 B.n214 585
R1477 B.n223 B.n222 585
R1478 B.n224 B.n213 585
R1479 B.n226 B.n225 585
R1480 B.n227 B.n212 585
R1481 B.n229 B.n228 585
R1482 B.n230 B.n211 585
R1483 B.n232 B.n231 585
R1484 B.n233 B.n210 585
R1485 B.n235 B.n234 585
R1486 B.n236 B.n209 585
R1487 B.n238 B.n237 585
R1488 B.n239 B.n208 585
R1489 B.n241 B.n240 585
R1490 B.n242 B.n207 585
R1491 B.n244 B.n243 585
R1492 B.n245 B.n206 585
R1493 B.n247 B.n246 585
R1494 B.n248 B.n205 585
R1495 B.n250 B.n249 585
R1496 B.n251 B.n204 585
R1497 B.n253 B.n252 585
R1498 B.n254 B.n203 585
R1499 B.n256 B.n255 585
R1500 B.n257 B.n202 585
R1501 B.n259 B.n258 585
R1502 B.n260 B.n201 585
R1503 B.n262 B.n261 585
R1504 B.n263 B.n200 585
R1505 B.n265 B.n264 585
R1506 B.n266 B.n199 585
R1507 B.n268 B.n267 585
R1508 B.n269 B.n198 585
R1509 B.n271 B.n270 585
R1510 B.n272 B.n197 585
R1511 B.n274 B.n273 585
R1512 B.n275 B.n196 585
R1513 B.n277 B.n276 585
R1514 B.n278 B.n195 585
R1515 B.n280 B.n279 585
R1516 B.n281 B.n194 585
R1517 B.n283 B.n282 585
R1518 B.n284 B.n193 585
R1519 B.n286 B.n285 585
R1520 B.n287 B.n192 585
R1521 B.n289 B.n288 585
R1522 B.n290 B.n191 585
R1523 B.n292 B.n291 585
R1524 B.n293 B.n190 585
R1525 B.n295 B.n294 585
R1526 B.n296 B.n189 585
R1527 B.n298 B.n189 497.305
R1528 B.n447 B.n446 497.305
R1529 B.n615 B.n614 497.305
R1530 B.n760 B.n29 497.305
R1531 B.n376 B.t10 451.002
R1532 B.n58 B.t5 451.002
R1533 B.n166 B.t7 451
R1534 B.n52 B.t2 451
R1535 B.n377 B.t11 388.553
R1536 B.n59 B.t4 388.553
R1537 B.n167 B.t8 388.553
R1538 B.n53 B.t1 388.553
R1539 B.n166 B.t6 314.519
R1540 B.n376 B.t9 314.519
R1541 B.n58 B.t3 314.519
R1542 B.n52 B.t0 314.519
R1543 B.n845 B.n844 256.663
R1544 B.n844 B.n843 235.042
R1545 B.n844 B.n2 235.042
R1546 B.n299 B.n298 163.367
R1547 B.n300 B.n299 163.367
R1548 B.n300 B.n187 163.367
R1549 B.n304 B.n187 163.367
R1550 B.n305 B.n304 163.367
R1551 B.n306 B.n305 163.367
R1552 B.n306 B.n185 163.367
R1553 B.n310 B.n185 163.367
R1554 B.n311 B.n310 163.367
R1555 B.n312 B.n311 163.367
R1556 B.n312 B.n183 163.367
R1557 B.n316 B.n183 163.367
R1558 B.n317 B.n316 163.367
R1559 B.n318 B.n317 163.367
R1560 B.n318 B.n181 163.367
R1561 B.n322 B.n181 163.367
R1562 B.n323 B.n322 163.367
R1563 B.n324 B.n323 163.367
R1564 B.n324 B.n179 163.367
R1565 B.n328 B.n179 163.367
R1566 B.n329 B.n328 163.367
R1567 B.n330 B.n329 163.367
R1568 B.n330 B.n177 163.367
R1569 B.n334 B.n177 163.367
R1570 B.n335 B.n334 163.367
R1571 B.n336 B.n335 163.367
R1572 B.n336 B.n175 163.367
R1573 B.n340 B.n175 163.367
R1574 B.n341 B.n340 163.367
R1575 B.n342 B.n341 163.367
R1576 B.n342 B.n173 163.367
R1577 B.n346 B.n173 163.367
R1578 B.n347 B.n346 163.367
R1579 B.n348 B.n347 163.367
R1580 B.n348 B.n171 163.367
R1581 B.n352 B.n171 163.367
R1582 B.n353 B.n352 163.367
R1583 B.n354 B.n353 163.367
R1584 B.n354 B.n169 163.367
R1585 B.n358 B.n169 163.367
R1586 B.n359 B.n358 163.367
R1587 B.n360 B.n359 163.367
R1588 B.n360 B.n165 163.367
R1589 B.n365 B.n165 163.367
R1590 B.n366 B.n365 163.367
R1591 B.n367 B.n366 163.367
R1592 B.n367 B.n163 163.367
R1593 B.n371 B.n163 163.367
R1594 B.n372 B.n371 163.367
R1595 B.n373 B.n372 163.367
R1596 B.n373 B.n161 163.367
R1597 B.n380 B.n161 163.367
R1598 B.n381 B.n380 163.367
R1599 B.n382 B.n381 163.367
R1600 B.n382 B.n159 163.367
R1601 B.n386 B.n159 163.367
R1602 B.n387 B.n386 163.367
R1603 B.n388 B.n387 163.367
R1604 B.n388 B.n157 163.367
R1605 B.n392 B.n157 163.367
R1606 B.n393 B.n392 163.367
R1607 B.n394 B.n393 163.367
R1608 B.n394 B.n155 163.367
R1609 B.n398 B.n155 163.367
R1610 B.n399 B.n398 163.367
R1611 B.n400 B.n399 163.367
R1612 B.n400 B.n153 163.367
R1613 B.n404 B.n153 163.367
R1614 B.n405 B.n404 163.367
R1615 B.n406 B.n405 163.367
R1616 B.n406 B.n151 163.367
R1617 B.n410 B.n151 163.367
R1618 B.n411 B.n410 163.367
R1619 B.n412 B.n411 163.367
R1620 B.n412 B.n149 163.367
R1621 B.n416 B.n149 163.367
R1622 B.n417 B.n416 163.367
R1623 B.n418 B.n417 163.367
R1624 B.n418 B.n147 163.367
R1625 B.n422 B.n147 163.367
R1626 B.n423 B.n422 163.367
R1627 B.n424 B.n423 163.367
R1628 B.n424 B.n145 163.367
R1629 B.n428 B.n145 163.367
R1630 B.n429 B.n428 163.367
R1631 B.n430 B.n429 163.367
R1632 B.n430 B.n143 163.367
R1633 B.n434 B.n143 163.367
R1634 B.n435 B.n434 163.367
R1635 B.n436 B.n435 163.367
R1636 B.n436 B.n141 163.367
R1637 B.n440 B.n141 163.367
R1638 B.n441 B.n440 163.367
R1639 B.n442 B.n441 163.367
R1640 B.n442 B.n139 163.367
R1641 B.n446 B.n139 163.367
R1642 B.n614 B.n83 163.367
R1643 B.n610 B.n83 163.367
R1644 B.n610 B.n609 163.367
R1645 B.n609 B.n608 163.367
R1646 B.n608 B.n85 163.367
R1647 B.n604 B.n85 163.367
R1648 B.n604 B.n603 163.367
R1649 B.n603 B.n602 163.367
R1650 B.n602 B.n87 163.367
R1651 B.n598 B.n87 163.367
R1652 B.n598 B.n597 163.367
R1653 B.n597 B.n596 163.367
R1654 B.n596 B.n89 163.367
R1655 B.n592 B.n89 163.367
R1656 B.n592 B.n591 163.367
R1657 B.n591 B.n590 163.367
R1658 B.n590 B.n91 163.367
R1659 B.n586 B.n91 163.367
R1660 B.n586 B.n585 163.367
R1661 B.n585 B.n584 163.367
R1662 B.n584 B.n93 163.367
R1663 B.n580 B.n93 163.367
R1664 B.n580 B.n579 163.367
R1665 B.n579 B.n578 163.367
R1666 B.n578 B.n95 163.367
R1667 B.n574 B.n95 163.367
R1668 B.n574 B.n573 163.367
R1669 B.n573 B.n572 163.367
R1670 B.n572 B.n97 163.367
R1671 B.n568 B.n97 163.367
R1672 B.n568 B.n567 163.367
R1673 B.n567 B.n566 163.367
R1674 B.n566 B.n99 163.367
R1675 B.n562 B.n99 163.367
R1676 B.n562 B.n561 163.367
R1677 B.n561 B.n560 163.367
R1678 B.n560 B.n101 163.367
R1679 B.n556 B.n101 163.367
R1680 B.n556 B.n555 163.367
R1681 B.n555 B.n554 163.367
R1682 B.n554 B.n103 163.367
R1683 B.n550 B.n103 163.367
R1684 B.n550 B.n549 163.367
R1685 B.n549 B.n548 163.367
R1686 B.n548 B.n105 163.367
R1687 B.n544 B.n105 163.367
R1688 B.n544 B.n543 163.367
R1689 B.n543 B.n542 163.367
R1690 B.n542 B.n107 163.367
R1691 B.n538 B.n107 163.367
R1692 B.n538 B.n537 163.367
R1693 B.n537 B.n536 163.367
R1694 B.n536 B.n109 163.367
R1695 B.n532 B.n109 163.367
R1696 B.n532 B.n531 163.367
R1697 B.n531 B.n530 163.367
R1698 B.n530 B.n111 163.367
R1699 B.n526 B.n111 163.367
R1700 B.n526 B.n525 163.367
R1701 B.n525 B.n524 163.367
R1702 B.n524 B.n113 163.367
R1703 B.n520 B.n113 163.367
R1704 B.n520 B.n519 163.367
R1705 B.n519 B.n518 163.367
R1706 B.n518 B.n115 163.367
R1707 B.n514 B.n115 163.367
R1708 B.n514 B.n513 163.367
R1709 B.n513 B.n512 163.367
R1710 B.n512 B.n117 163.367
R1711 B.n508 B.n117 163.367
R1712 B.n508 B.n507 163.367
R1713 B.n507 B.n506 163.367
R1714 B.n506 B.n119 163.367
R1715 B.n502 B.n119 163.367
R1716 B.n502 B.n501 163.367
R1717 B.n501 B.n500 163.367
R1718 B.n500 B.n121 163.367
R1719 B.n496 B.n121 163.367
R1720 B.n496 B.n495 163.367
R1721 B.n495 B.n494 163.367
R1722 B.n494 B.n123 163.367
R1723 B.n490 B.n123 163.367
R1724 B.n490 B.n489 163.367
R1725 B.n489 B.n488 163.367
R1726 B.n488 B.n125 163.367
R1727 B.n484 B.n125 163.367
R1728 B.n484 B.n483 163.367
R1729 B.n483 B.n482 163.367
R1730 B.n482 B.n127 163.367
R1731 B.n478 B.n127 163.367
R1732 B.n478 B.n477 163.367
R1733 B.n477 B.n476 163.367
R1734 B.n476 B.n129 163.367
R1735 B.n472 B.n129 163.367
R1736 B.n472 B.n471 163.367
R1737 B.n471 B.n470 163.367
R1738 B.n470 B.n131 163.367
R1739 B.n466 B.n131 163.367
R1740 B.n466 B.n465 163.367
R1741 B.n465 B.n464 163.367
R1742 B.n464 B.n133 163.367
R1743 B.n460 B.n133 163.367
R1744 B.n460 B.n459 163.367
R1745 B.n459 B.n458 163.367
R1746 B.n458 B.n135 163.367
R1747 B.n454 B.n135 163.367
R1748 B.n454 B.n453 163.367
R1749 B.n453 B.n452 163.367
R1750 B.n452 B.n137 163.367
R1751 B.n448 B.n137 163.367
R1752 B.n448 B.n447 163.367
R1753 B.n760 B.n759 163.367
R1754 B.n759 B.n758 163.367
R1755 B.n758 B.n31 163.367
R1756 B.n754 B.n31 163.367
R1757 B.n754 B.n753 163.367
R1758 B.n753 B.n752 163.367
R1759 B.n752 B.n33 163.367
R1760 B.n748 B.n33 163.367
R1761 B.n748 B.n747 163.367
R1762 B.n747 B.n746 163.367
R1763 B.n746 B.n35 163.367
R1764 B.n742 B.n35 163.367
R1765 B.n742 B.n741 163.367
R1766 B.n741 B.n740 163.367
R1767 B.n740 B.n37 163.367
R1768 B.n736 B.n37 163.367
R1769 B.n736 B.n735 163.367
R1770 B.n735 B.n734 163.367
R1771 B.n734 B.n39 163.367
R1772 B.n730 B.n39 163.367
R1773 B.n730 B.n729 163.367
R1774 B.n729 B.n728 163.367
R1775 B.n728 B.n41 163.367
R1776 B.n724 B.n41 163.367
R1777 B.n724 B.n723 163.367
R1778 B.n723 B.n722 163.367
R1779 B.n722 B.n43 163.367
R1780 B.n718 B.n43 163.367
R1781 B.n718 B.n717 163.367
R1782 B.n717 B.n716 163.367
R1783 B.n716 B.n45 163.367
R1784 B.n712 B.n45 163.367
R1785 B.n712 B.n711 163.367
R1786 B.n711 B.n710 163.367
R1787 B.n710 B.n47 163.367
R1788 B.n706 B.n47 163.367
R1789 B.n706 B.n705 163.367
R1790 B.n705 B.n704 163.367
R1791 B.n704 B.n49 163.367
R1792 B.n700 B.n49 163.367
R1793 B.n700 B.n699 163.367
R1794 B.n699 B.n698 163.367
R1795 B.n698 B.n51 163.367
R1796 B.n693 B.n51 163.367
R1797 B.n693 B.n692 163.367
R1798 B.n692 B.n691 163.367
R1799 B.n691 B.n55 163.367
R1800 B.n687 B.n55 163.367
R1801 B.n687 B.n686 163.367
R1802 B.n686 B.n685 163.367
R1803 B.n685 B.n57 163.367
R1804 B.n681 B.n57 163.367
R1805 B.n681 B.n680 163.367
R1806 B.n680 B.n61 163.367
R1807 B.n676 B.n61 163.367
R1808 B.n676 B.n675 163.367
R1809 B.n675 B.n674 163.367
R1810 B.n674 B.n63 163.367
R1811 B.n670 B.n63 163.367
R1812 B.n670 B.n669 163.367
R1813 B.n669 B.n668 163.367
R1814 B.n668 B.n65 163.367
R1815 B.n664 B.n65 163.367
R1816 B.n664 B.n663 163.367
R1817 B.n663 B.n662 163.367
R1818 B.n662 B.n67 163.367
R1819 B.n658 B.n67 163.367
R1820 B.n658 B.n657 163.367
R1821 B.n657 B.n656 163.367
R1822 B.n656 B.n69 163.367
R1823 B.n652 B.n69 163.367
R1824 B.n652 B.n651 163.367
R1825 B.n651 B.n650 163.367
R1826 B.n650 B.n71 163.367
R1827 B.n646 B.n71 163.367
R1828 B.n646 B.n645 163.367
R1829 B.n645 B.n644 163.367
R1830 B.n644 B.n73 163.367
R1831 B.n640 B.n73 163.367
R1832 B.n640 B.n639 163.367
R1833 B.n639 B.n638 163.367
R1834 B.n638 B.n75 163.367
R1835 B.n634 B.n75 163.367
R1836 B.n634 B.n633 163.367
R1837 B.n633 B.n632 163.367
R1838 B.n632 B.n77 163.367
R1839 B.n628 B.n77 163.367
R1840 B.n628 B.n627 163.367
R1841 B.n627 B.n626 163.367
R1842 B.n626 B.n79 163.367
R1843 B.n622 B.n79 163.367
R1844 B.n622 B.n621 163.367
R1845 B.n621 B.n620 163.367
R1846 B.n620 B.n81 163.367
R1847 B.n616 B.n81 163.367
R1848 B.n616 B.n615 163.367
R1849 B.n764 B.n29 163.367
R1850 B.n765 B.n764 163.367
R1851 B.n766 B.n765 163.367
R1852 B.n766 B.n27 163.367
R1853 B.n770 B.n27 163.367
R1854 B.n771 B.n770 163.367
R1855 B.n772 B.n771 163.367
R1856 B.n772 B.n25 163.367
R1857 B.n776 B.n25 163.367
R1858 B.n777 B.n776 163.367
R1859 B.n778 B.n777 163.367
R1860 B.n778 B.n23 163.367
R1861 B.n782 B.n23 163.367
R1862 B.n783 B.n782 163.367
R1863 B.n784 B.n783 163.367
R1864 B.n784 B.n21 163.367
R1865 B.n788 B.n21 163.367
R1866 B.n789 B.n788 163.367
R1867 B.n790 B.n789 163.367
R1868 B.n790 B.n19 163.367
R1869 B.n794 B.n19 163.367
R1870 B.n795 B.n794 163.367
R1871 B.n796 B.n795 163.367
R1872 B.n796 B.n17 163.367
R1873 B.n800 B.n17 163.367
R1874 B.n801 B.n800 163.367
R1875 B.n802 B.n801 163.367
R1876 B.n802 B.n15 163.367
R1877 B.n806 B.n15 163.367
R1878 B.n807 B.n806 163.367
R1879 B.n808 B.n807 163.367
R1880 B.n808 B.n13 163.367
R1881 B.n812 B.n13 163.367
R1882 B.n813 B.n812 163.367
R1883 B.n814 B.n813 163.367
R1884 B.n814 B.n11 163.367
R1885 B.n818 B.n11 163.367
R1886 B.n819 B.n818 163.367
R1887 B.n820 B.n819 163.367
R1888 B.n820 B.n9 163.367
R1889 B.n824 B.n9 163.367
R1890 B.n825 B.n824 163.367
R1891 B.n826 B.n825 163.367
R1892 B.n826 B.n7 163.367
R1893 B.n830 B.n7 163.367
R1894 B.n831 B.n830 163.367
R1895 B.n832 B.n831 163.367
R1896 B.n832 B.n5 163.367
R1897 B.n836 B.n5 163.367
R1898 B.n837 B.n836 163.367
R1899 B.n838 B.n837 163.367
R1900 B.n838 B.n3 163.367
R1901 B.n842 B.n3 163.367
R1902 B.n843 B.n842 163.367
R1903 B.n216 B.n2 163.367
R1904 B.n216 B.n215 163.367
R1905 B.n220 B.n215 163.367
R1906 B.n221 B.n220 163.367
R1907 B.n222 B.n221 163.367
R1908 B.n222 B.n213 163.367
R1909 B.n226 B.n213 163.367
R1910 B.n227 B.n226 163.367
R1911 B.n228 B.n227 163.367
R1912 B.n228 B.n211 163.367
R1913 B.n232 B.n211 163.367
R1914 B.n233 B.n232 163.367
R1915 B.n234 B.n233 163.367
R1916 B.n234 B.n209 163.367
R1917 B.n238 B.n209 163.367
R1918 B.n239 B.n238 163.367
R1919 B.n240 B.n239 163.367
R1920 B.n240 B.n207 163.367
R1921 B.n244 B.n207 163.367
R1922 B.n245 B.n244 163.367
R1923 B.n246 B.n245 163.367
R1924 B.n246 B.n205 163.367
R1925 B.n250 B.n205 163.367
R1926 B.n251 B.n250 163.367
R1927 B.n252 B.n251 163.367
R1928 B.n252 B.n203 163.367
R1929 B.n256 B.n203 163.367
R1930 B.n257 B.n256 163.367
R1931 B.n258 B.n257 163.367
R1932 B.n258 B.n201 163.367
R1933 B.n262 B.n201 163.367
R1934 B.n263 B.n262 163.367
R1935 B.n264 B.n263 163.367
R1936 B.n264 B.n199 163.367
R1937 B.n268 B.n199 163.367
R1938 B.n269 B.n268 163.367
R1939 B.n270 B.n269 163.367
R1940 B.n270 B.n197 163.367
R1941 B.n274 B.n197 163.367
R1942 B.n275 B.n274 163.367
R1943 B.n276 B.n275 163.367
R1944 B.n276 B.n195 163.367
R1945 B.n280 B.n195 163.367
R1946 B.n281 B.n280 163.367
R1947 B.n282 B.n281 163.367
R1948 B.n282 B.n193 163.367
R1949 B.n286 B.n193 163.367
R1950 B.n287 B.n286 163.367
R1951 B.n288 B.n287 163.367
R1952 B.n288 B.n191 163.367
R1953 B.n292 B.n191 163.367
R1954 B.n293 B.n292 163.367
R1955 B.n294 B.n293 163.367
R1956 B.n294 B.n189 163.367
R1957 B.n167 B.n166 62.449
R1958 B.n377 B.n376 62.449
R1959 B.n59 B.n58 62.449
R1960 B.n53 B.n52 62.449
R1961 B.n363 B.n167 59.5399
R1962 B.n378 B.n377 59.5399
R1963 B.n60 B.n59 59.5399
R1964 B.n695 B.n53 59.5399
R1965 B.n762 B.n761 32.3127
R1966 B.n613 B.n82 32.3127
R1967 B.n445 B.n138 32.3127
R1968 B.n297 B.n296 32.3127
R1969 B B.n845 18.0485
R1970 B.n763 B.n762 10.6151
R1971 B.n763 B.n28 10.6151
R1972 B.n767 B.n28 10.6151
R1973 B.n768 B.n767 10.6151
R1974 B.n769 B.n768 10.6151
R1975 B.n769 B.n26 10.6151
R1976 B.n773 B.n26 10.6151
R1977 B.n774 B.n773 10.6151
R1978 B.n775 B.n774 10.6151
R1979 B.n775 B.n24 10.6151
R1980 B.n779 B.n24 10.6151
R1981 B.n780 B.n779 10.6151
R1982 B.n781 B.n780 10.6151
R1983 B.n781 B.n22 10.6151
R1984 B.n785 B.n22 10.6151
R1985 B.n786 B.n785 10.6151
R1986 B.n787 B.n786 10.6151
R1987 B.n787 B.n20 10.6151
R1988 B.n791 B.n20 10.6151
R1989 B.n792 B.n791 10.6151
R1990 B.n793 B.n792 10.6151
R1991 B.n793 B.n18 10.6151
R1992 B.n797 B.n18 10.6151
R1993 B.n798 B.n797 10.6151
R1994 B.n799 B.n798 10.6151
R1995 B.n799 B.n16 10.6151
R1996 B.n803 B.n16 10.6151
R1997 B.n804 B.n803 10.6151
R1998 B.n805 B.n804 10.6151
R1999 B.n805 B.n14 10.6151
R2000 B.n809 B.n14 10.6151
R2001 B.n810 B.n809 10.6151
R2002 B.n811 B.n810 10.6151
R2003 B.n811 B.n12 10.6151
R2004 B.n815 B.n12 10.6151
R2005 B.n816 B.n815 10.6151
R2006 B.n817 B.n816 10.6151
R2007 B.n817 B.n10 10.6151
R2008 B.n821 B.n10 10.6151
R2009 B.n822 B.n821 10.6151
R2010 B.n823 B.n822 10.6151
R2011 B.n823 B.n8 10.6151
R2012 B.n827 B.n8 10.6151
R2013 B.n828 B.n827 10.6151
R2014 B.n829 B.n828 10.6151
R2015 B.n829 B.n6 10.6151
R2016 B.n833 B.n6 10.6151
R2017 B.n834 B.n833 10.6151
R2018 B.n835 B.n834 10.6151
R2019 B.n835 B.n4 10.6151
R2020 B.n839 B.n4 10.6151
R2021 B.n840 B.n839 10.6151
R2022 B.n841 B.n840 10.6151
R2023 B.n841 B.n0 10.6151
R2024 B.n761 B.n30 10.6151
R2025 B.n757 B.n30 10.6151
R2026 B.n757 B.n756 10.6151
R2027 B.n756 B.n755 10.6151
R2028 B.n755 B.n32 10.6151
R2029 B.n751 B.n32 10.6151
R2030 B.n751 B.n750 10.6151
R2031 B.n750 B.n749 10.6151
R2032 B.n749 B.n34 10.6151
R2033 B.n745 B.n34 10.6151
R2034 B.n745 B.n744 10.6151
R2035 B.n744 B.n743 10.6151
R2036 B.n743 B.n36 10.6151
R2037 B.n739 B.n36 10.6151
R2038 B.n739 B.n738 10.6151
R2039 B.n738 B.n737 10.6151
R2040 B.n737 B.n38 10.6151
R2041 B.n733 B.n38 10.6151
R2042 B.n733 B.n732 10.6151
R2043 B.n732 B.n731 10.6151
R2044 B.n731 B.n40 10.6151
R2045 B.n727 B.n40 10.6151
R2046 B.n727 B.n726 10.6151
R2047 B.n726 B.n725 10.6151
R2048 B.n725 B.n42 10.6151
R2049 B.n721 B.n42 10.6151
R2050 B.n721 B.n720 10.6151
R2051 B.n720 B.n719 10.6151
R2052 B.n719 B.n44 10.6151
R2053 B.n715 B.n44 10.6151
R2054 B.n715 B.n714 10.6151
R2055 B.n714 B.n713 10.6151
R2056 B.n713 B.n46 10.6151
R2057 B.n709 B.n46 10.6151
R2058 B.n709 B.n708 10.6151
R2059 B.n708 B.n707 10.6151
R2060 B.n707 B.n48 10.6151
R2061 B.n703 B.n48 10.6151
R2062 B.n703 B.n702 10.6151
R2063 B.n702 B.n701 10.6151
R2064 B.n701 B.n50 10.6151
R2065 B.n697 B.n50 10.6151
R2066 B.n697 B.n696 10.6151
R2067 B.n694 B.n54 10.6151
R2068 B.n690 B.n54 10.6151
R2069 B.n690 B.n689 10.6151
R2070 B.n689 B.n688 10.6151
R2071 B.n688 B.n56 10.6151
R2072 B.n684 B.n56 10.6151
R2073 B.n684 B.n683 10.6151
R2074 B.n683 B.n682 10.6151
R2075 B.n679 B.n678 10.6151
R2076 B.n678 B.n677 10.6151
R2077 B.n677 B.n62 10.6151
R2078 B.n673 B.n62 10.6151
R2079 B.n673 B.n672 10.6151
R2080 B.n672 B.n671 10.6151
R2081 B.n671 B.n64 10.6151
R2082 B.n667 B.n64 10.6151
R2083 B.n667 B.n666 10.6151
R2084 B.n666 B.n665 10.6151
R2085 B.n665 B.n66 10.6151
R2086 B.n661 B.n66 10.6151
R2087 B.n661 B.n660 10.6151
R2088 B.n660 B.n659 10.6151
R2089 B.n659 B.n68 10.6151
R2090 B.n655 B.n68 10.6151
R2091 B.n655 B.n654 10.6151
R2092 B.n654 B.n653 10.6151
R2093 B.n653 B.n70 10.6151
R2094 B.n649 B.n70 10.6151
R2095 B.n649 B.n648 10.6151
R2096 B.n648 B.n647 10.6151
R2097 B.n647 B.n72 10.6151
R2098 B.n643 B.n72 10.6151
R2099 B.n643 B.n642 10.6151
R2100 B.n642 B.n641 10.6151
R2101 B.n641 B.n74 10.6151
R2102 B.n637 B.n74 10.6151
R2103 B.n637 B.n636 10.6151
R2104 B.n636 B.n635 10.6151
R2105 B.n635 B.n76 10.6151
R2106 B.n631 B.n76 10.6151
R2107 B.n631 B.n630 10.6151
R2108 B.n630 B.n629 10.6151
R2109 B.n629 B.n78 10.6151
R2110 B.n625 B.n78 10.6151
R2111 B.n625 B.n624 10.6151
R2112 B.n624 B.n623 10.6151
R2113 B.n623 B.n80 10.6151
R2114 B.n619 B.n80 10.6151
R2115 B.n619 B.n618 10.6151
R2116 B.n618 B.n617 10.6151
R2117 B.n617 B.n82 10.6151
R2118 B.n613 B.n612 10.6151
R2119 B.n612 B.n611 10.6151
R2120 B.n611 B.n84 10.6151
R2121 B.n607 B.n84 10.6151
R2122 B.n607 B.n606 10.6151
R2123 B.n606 B.n605 10.6151
R2124 B.n605 B.n86 10.6151
R2125 B.n601 B.n86 10.6151
R2126 B.n601 B.n600 10.6151
R2127 B.n600 B.n599 10.6151
R2128 B.n599 B.n88 10.6151
R2129 B.n595 B.n88 10.6151
R2130 B.n595 B.n594 10.6151
R2131 B.n594 B.n593 10.6151
R2132 B.n593 B.n90 10.6151
R2133 B.n589 B.n90 10.6151
R2134 B.n589 B.n588 10.6151
R2135 B.n588 B.n587 10.6151
R2136 B.n587 B.n92 10.6151
R2137 B.n583 B.n92 10.6151
R2138 B.n583 B.n582 10.6151
R2139 B.n582 B.n581 10.6151
R2140 B.n581 B.n94 10.6151
R2141 B.n577 B.n94 10.6151
R2142 B.n577 B.n576 10.6151
R2143 B.n576 B.n575 10.6151
R2144 B.n575 B.n96 10.6151
R2145 B.n571 B.n96 10.6151
R2146 B.n571 B.n570 10.6151
R2147 B.n570 B.n569 10.6151
R2148 B.n569 B.n98 10.6151
R2149 B.n565 B.n98 10.6151
R2150 B.n565 B.n564 10.6151
R2151 B.n564 B.n563 10.6151
R2152 B.n563 B.n100 10.6151
R2153 B.n559 B.n100 10.6151
R2154 B.n559 B.n558 10.6151
R2155 B.n558 B.n557 10.6151
R2156 B.n557 B.n102 10.6151
R2157 B.n553 B.n102 10.6151
R2158 B.n553 B.n552 10.6151
R2159 B.n552 B.n551 10.6151
R2160 B.n551 B.n104 10.6151
R2161 B.n547 B.n104 10.6151
R2162 B.n547 B.n546 10.6151
R2163 B.n546 B.n545 10.6151
R2164 B.n545 B.n106 10.6151
R2165 B.n541 B.n106 10.6151
R2166 B.n541 B.n540 10.6151
R2167 B.n540 B.n539 10.6151
R2168 B.n539 B.n108 10.6151
R2169 B.n535 B.n108 10.6151
R2170 B.n535 B.n534 10.6151
R2171 B.n534 B.n533 10.6151
R2172 B.n533 B.n110 10.6151
R2173 B.n529 B.n110 10.6151
R2174 B.n529 B.n528 10.6151
R2175 B.n528 B.n527 10.6151
R2176 B.n527 B.n112 10.6151
R2177 B.n523 B.n112 10.6151
R2178 B.n523 B.n522 10.6151
R2179 B.n522 B.n521 10.6151
R2180 B.n521 B.n114 10.6151
R2181 B.n517 B.n114 10.6151
R2182 B.n517 B.n516 10.6151
R2183 B.n516 B.n515 10.6151
R2184 B.n515 B.n116 10.6151
R2185 B.n511 B.n116 10.6151
R2186 B.n511 B.n510 10.6151
R2187 B.n510 B.n509 10.6151
R2188 B.n509 B.n118 10.6151
R2189 B.n505 B.n118 10.6151
R2190 B.n505 B.n504 10.6151
R2191 B.n504 B.n503 10.6151
R2192 B.n503 B.n120 10.6151
R2193 B.n499 B.n120 10.6151
R2194 B.n499 B.n498 10.6151
R2195 B.n498 B.n497 10.6151
R2196 B.n497 B.n122 10.6151
R2197 B.n493 B.n122 10.6151
R2198 B.n493 B.n492 10.6151
R2199 B.n492 B.n491 10.6151
R2200 B.n491 B.n124 10.6151
R2201 B.n487 B.n124 10.6151
R2202 B.n487 B.n486 10.6151
R2203 B.n486 B.n485 10.6151
R2204 B.n485 B.n126 10.6151
R2205 B.n481 B.n126 10.6151
R2206 B.n481 B.n480 10.6151
R2207 B.n480 B.n479 10.6151
R2208 B.n479 B.n128 10.6151
R2209 B.n475 B.n128 10.6151
R2210 B.n475 B.n474 10.6151
R2211 B.n474 B.n473 10.6151
R2212 B.n473 B.n130 10.6151
R2213 B.n469 B.n130 10.6151
R2214 B.n469 B.n468 10.6151
R2215 B.n468 B.n467 10.6151
R2216 B.n467 B.n132 10.6151
R2217 B.n463 B.n132 10.6151
R2218 B.n463 B.n462 10.6151
R2219 B.n462 B.n461 10.6151
R2220 B.n461 B.n134 10.6151
R2221 B.n457 B.n134 10.6151
R2222 B.n457 B.n456 10.6151
R2223 B.n456 B.n455 10.6151
R2224 B.n455 B.n136 10.6151
R2225 B.n451 B.n136 10.6151
R2226 B.n451 B.n450 10.6151
R2227 B.n450 B.n449 10.6151
R2228 B.n449 B.n138 10.6151
R2229 B.n217 B.n1 10.6151
R2230 B.n218 B.n217 10.6151
R2231 B.n219 B.n218 10.6151
R2232 B.n219 B.n214 10.6151
R2233 B.n223 B.n214 10.6151
R2234 B.n224 B.n223 10.6151
R2235 B.n225 B.n224 10.6151
R2236 B.n225 B.n212 10.6151
R2237 B.n229 B.n212 10.6151
R2238 B.n230 B.n229 10.6151
R2239 B.n231 B.n230 10.6151
R2240 B.n231 B.n210 10.6151
R2241 B.n235 B.n210 10.6151
R2242 B.n236 B.n235 10.6151
R2243 B.n237 B.n236 10.6151
R2244 B.n237 B.n208 10.6151
R2245 B.n241 B.n208 10.6151
R2246 B.n242 B.n241 10.6151
R2247 B.n243 B.n242 10.6151
R2248 B.n243 B.n206 10.6151
R2249 B.n247 B.n206 10.6151
R2250 B.n248 B.n247 10.6151
R2251 B.n249 B.n248 10.6151
R2252 B.n249 B.n204 10.6151
R2253 B.n253 B.n204 10.6151
R2254 B.n254 B.n253 10.6151
R2255 B.n255 B.n254 10.6151
R2256 B.n255 B.n202 10.6151
R2257 B.n259 B.n202 10.6151
R2258 B.n260 B.n259 10.6151
R2259 B.n261 B.n260 10.6151
R2260 B.n261 B.n200 10.6151
R2261 B.n265 B.n200 10.6151
R2262 B.n266 B.n265 10.6151
R2263 B.n267 B.n266 10.6151
R2264 B.n267 B.n198 10.6151
R2265 B.n271 B.n198 10.6151
R2266 B.n272 B.n271 10.6151
R2267 B.n273 B.n272 10.6151
R2268 B.n273 B.n196 10.6151
R2269 B.n277 B.n196 10.6151
R2270 B.n278 B.n277 10.6151
R2271 B.n279 B.n278 10.6151
R2272 B.n279 B.n194 10.6151
R2273 B.n283 B.n194 10.6151
R2274 B.n284 B.n283 10.6151
R2275 B.n285 B.n284 10.6151
R2276 B.n285 B.n192 10.6151
R2277 B.n289 B.n192 10.6151
R2278 B.n290 B.n289 10.6151
R2279 B.n291 B.n290 10.6151
R2280 B.n291 B.n190 10.6151
R2281 B.n295 B.n190 10.6151
R2282 B.n296 B.n295 10.6151
R2283 B.n297 B.n188 10.6151
R2284 B.n301 B.n188 10.6151
R2285 B.n302 B.n301 10.6151
R2286 B.n303 B.n302 10.6151
R2287 B.n303 B.n186 10.6151
R2288 B.n307 B.n186 10.6151
R2289 B.n308 B.n307 10.6151
R2290 B.n309 B.n308 10.6151
R2291 B.n309 B.n184 10.6151
R2292 B.n313 B.n184 10.6151
R2293 B.n314 B.n313 10.6151
R2294 B.n315 B.n314 10.6151
R2295 B.n315 B.n182 10.6151
R2296 B.n319 B.n182 10.6151
R2297 B.n320 B.n319 10.6151
R2298 B.n321 B.n320 10.6151
R2299 B.n321 B.n180 10.6151
R2300 B.n325 B.n180 10.6151
R2301 B.n326 B.n325 10.6151
R2302 B.n327 B.n326 10.6151
R2303 B.n327 B.n178 10.6151
R2304 B.n331 B.n178 10.6151
R2305 B.n332 B.n331 10.6151
R2306 B.n333 B.n332 10.6151
R2307 B.n333 B.n176 10.6151
R2308 B.n337 B.n176 10.6151
R2309 B.n338 B.n337 10.6151
R2310 B.n339 B.n338 10.6151
R2311 B.n339 B.n174 10.6151
R2312 B.n343 B.n174 10.6151
R2313 B.n344 B.n343 10.6151
R2314 B.n345 B.n344 10.6151
R2315 B.n345 B.n172 10.6151
R2316 B.n349 B.n172 10.6151
R2317 B.n350 B.n349 10.6151
R2318 B.n351 B.n350 10.6151
R2319 B.n351 B.n170 10.6151
R2320 B.n355 B.n170 10.6151
R2321 B.n356 B.n355 10.6151
R2322 B.n357 B.n356 10.6151
R2323 B.n357 B.n168 10.6151
R2324 B.n361 B.n168 10.6151
R2325 B.n362 B.n361 10.6151
R2326 B.n364 B.n164 10.6151
R2327 B.n368 B.n164 10.6151
R2328 B.n369 B.n368 10.6151
R2329 B.n370 B.n369 10.6151
R2330 B.n370 B.n162 10.6151
R2331 B.n374 B.n162 10.6151
R2332 B.n375 B.n374 10.6151
R2333 B.n379 B.n375 10.6151
R2334 B.n383 B.n160 10.6151
R2335 B.n384 B.n383 10.6151
R2336 B.n385 B.n384 10.6151
R2337 B.n385 B.n158 10.6151
R2338 B.n389 B.n158 10.6151
R2339 B.n390 B.n389 10.6151
R2340 B.n391 B.n390 10.6151
R2341 B.n391 B.n156 10.6151
R2342 B.n395 B.n156 10.6151
R2343 B.n396 B.n395 10.6151
R2344 B.n397 B.n396 10.6151
R2345 B.n397 B.n154 10.6151
R2346 B.n401 B.n154 10.6151
R2347 B.n402 B.n401 10.6151
R2348 B.n403 B.n402 10.6151
R2349 B.n403 B.n152 10.6151
R2350 B.n407 B.n152 10.6151
R2351 B.n408 B.n407 10.6151
R2352 B.n409 B.n408 10.6151
R2353 B.n409 B.n150 10.6151
R2354 B.n413 B.n150 10.6151
R2355 B.n414 B.n413 10.6151
R2356 B.n415 B.n414 10.6151
R2357 B.n415 B.n148 10.6151
R2358 B.n419 B.n148 10.6151
R2359 B.n420 B.n419 10.6151
R2360 B.n421 B.n420 10.6151
R2361 B.n421 B.n146 10.6151
R2362 B.n425 B.n146 10.6151
R2363 B.n426 B.n425 10.6151
R2364 B.n427 B.n426 10.6151
R2365 B.n427 B.n144 10.6151
R2366 B.n431 B.n144 10.6151
R2367 B.n432 B.n431 10.6151
R2368 B.n433 B.n432 10.6151
R2369 B.n433 B.n142 10.6151
R2370 B.n437 B.n142 10.6151
R2371 B.n438 B.n437 10.6151
R2372 B.n439 B.n438 10.6151
R2373 B.n439 B.n140 10.6151
R2374 B.n443 B.n140 10.6151
R2375 B.n444 B.n443 10.6151
R2376 B.n445 B.n444 10.6151
R2377 B.n845 B.n0 8.11757
R2378 B.n845 B.n1 8.11757
R2379 B.n695 B.n694 6.5566
R2380 B.n682 B.n60 6.5566
R2381 B.n364 B.n363 6.5566
R2382 B.n379 B.n378 6.5566
R2383 B.n696 B.n695 4.05904
R2384 B.n679 B.n60 4.05904
R2385 B.n363 B.n362 4.05904
R2386 B.n378 B.n160 4.05904
C0 VP VDD2 0.549816f
C1 VP VN 8.15529f
C2 VP w_n4190_n3512# 9.17418f
C3 B VP 2.21195f
C4 VTAIL VDD1 8.38212f
C5 VTAIL VDD2 8.43848f
C6 VDD1 VDD2 1.92577f
C7 VN VTAIL 9.83145f
C8 VN VDD1 0.151539f
C9 w_n4190_n3512# VTAIL 4.39778f
C10 w_n4190_n3512# VDD1 2.06227f
C11 VN VDD2 9.379f
C12 w_n4190_n3512# VDD2 2.18914f
C13 w_n4190_n3512# VN 8.62938f
C14 B VTAIL 5.35206f
C15 B VDD1 1.75651f
C16 VP VTAIL 9.845559f
C17 VP VDD1 9.77573f
C18 B VDD2 1.86166f
C19 B VN 1.29712f
C20 B w_n4190_n3512# 10.7616f
C21 VDD2 VSUBS 2.009299f
C22 VDD1 VSUBS 2.71114f
C23 VTAIL VSUBS 1.419305f
C24 VN VSUBS 7.13379f
C25 VP VSUBS 3.902028f
C26 B VSUBS 5.389269f
C27 w_n4190_n3512# VSUBS 0.180958p
C28 B.n0 VSUBS 0.00651f
C29 B.n1 VSUBS 0.00651f
C30 B.n2 VSUBS 0.009628f
C31 B.n3 VSUBS 0.007378f
C32 B.n4 VSUBS 0.007378f
C33 B.n5 VSUBS 0.007378f
C34 B.n6 VSUBS 0.007378f
C35 B.n7 VSUBS 0.007378f
C36 B.n8 VSUBS 0.007378f
C37 B.n9 VSUBS 0.007378f
C38 B.n10 VSUBS 0.007378f
C39 B.n11 VSUBS 0.007378f
C40 B.n12 VSUBS 0.007378f
C41 B.n13 VSUBS 0.007378f
C42 B.n14 VSUBS 0.007378f
C43 B.n15 VSUBS 0.007378f
C44 B.n16 VSUBS 0.007378f
C45 B.n17 VSUBS 0.007378f
C46 B.n18 VSUBS 0.007378f
C47 B.n19 VSUBS 0.007378f
C48 B.n20 VSUBS 0.007378f
C49 B.n21 VSUBS 0.007378f
C50 B.n22 VSUBS 0.007378f
C51 B.n23 VSUBS 0.007378f
C52 B.n24 VSUBS 0.007378f
C53 B.n25 VSUBS 0.007378f
C54 B.n26 VSUBS 0.007378f
C55 B.n27 VSUBS 0.007378f
C56 B.n28 VSUBS 0.007378f
C57 B.n29 VSUBS 0.016767f
C58 B.n30 VSUBS 0.007378f
C59 B.n31 VSUBS 0.007378f
C60 B.n32 VSUBS 0.007378f
C61 B.n33 VSUBS 0.007378f
C62 B.n34 VSUBS 0.007378f
C63 B.n35 VSUBS 0.007378f
C64 B.n36 VSUBS 0.007378f
C65 B.n37 VSUBS 0.007378f
C66 B.n38 VSUBS 0.007378f
C67 B.n39 VSUBS 0.007378f
C68 B.n40 VSUBS 0.007378f
C69 B.n41 VSUBS 0.007378f
C70 B.n42 VSUBS 0.007378f
C71 B.n43 VSUBS 0.007378f
C72 B.n44 VSUBS 0.007378f
C73 B.n45 VSUBS 0.007378f
C74 B.n46 VSUBS 0.007378f
C75 B.n47 VSUBS 0.007378f
C76 B.n48 VSUBS 0.007378f
C77 B.n49 VSUBS 0.007378f
C78 B.n50 VSUBS 0.007378f
C79 B.n51 VSUBS 0.007378f
C80 B.t1 VSUBS 0.23938f
C81 B.t2 VSUBS 0.276304f
C82 B.t0 VSUBS 1.77104f
C83 B.n52 VSUBS 0.438265f
C84 B.n53 VSUBS 0.27719f
C85 B.n54 VSUBS 0.007378f
C86 B.n55 VSUBS 0.007378f
C87 B.n56 VSUBS 0.007378f
C88 B.n57 VSUBS 0.007378f
C89 B.t4 VSUBS 0.239383f
C90 B.t5 VSUBS 0.276307f
C91 B.t3 VSUBS 1.77104f
C92 B.n58 VSUBS 0.438262f
C93 B.n59 VSUBS 0.277187f
C94 B.n60 VSUBS 0.017095f
C95 B.n61 VSUBS 0.007378f
C96 B.n62 VSUBS 0.007378f
C97 B.n63 VSUBS 0.007378f
C98 B.n64 VSUBS 0.007378f
C99 B.n65 VSUBS 0.007378f
C100 B.n66 VSUBS 0.007378f
C101 B.n67 VSUBS 0.007378f
C102 B.n68 VSUBS 0.007378f
C103 B.n69 VSUBS 0.007378f
C104 B.n70 VSUBS 0.007378f
C105 B.n71 VSUBS 0.007378f
C106 B.n72 VSUBS 0.007378f
C107 B.n73 VSUBS 0.007378f
C108 B.n74 VSUBS 0.007378f
C109 B.n75 VSUBS 0.007378f
C110 B.n76 VSUBS 0.007378f
C111 B.n77 VSUBS 0.007378f
C112 B.n78 VSUBS 0.007378f
C113 B.n79 VSUBS 0.007378f
C114 B.n80 VSUBS 0.007378f
C115 B.n81 VSUBS 0.007378f
C116 B.n82 VSUBS 0.01752f
C117 B.n83 VSUBS 0.007378f
C118 B.n84 VSUBS 0.007378f
C119 B.n85 VSUBS 0.007378f
C120 B.n86 VSUBS 0.007378f
C121 B.n87 VSUBS 0.007378f
C122 B.n88 VSUBS 0.007378f
C123 B.n89 VSUBS 0.007378f
C124 B.n90 VSUBS 0.007378f
C125 B.n91 VSUBS 0.007378f
C126 B.n92 VSUBS 0.007378f
C127 B.n93 VSUBS 0.007378f
C128 B.n94 VSUBS 0.007378f
C129 B.n95 VSUBS 0.007378f
C130 B.n96 VSUBS 0.007378f
C131 B.n97 VSUBS 0.007378f
C132 B.n98 VSUBS 0.007378f
C133 B.n99 VSUBS 0.007378f
C134 B.n100 VSUBS 0.007378f
C135 B.n101 VSUBS 0.007378f
C136 B.n102 VSUBS 0.007378f
C137 B.n103 VSUBS 0.007378f
C138 B.n104 VSUBS 0.007378f
C139 B.n105 VSUBS 0.007378f
C140 B.n106 VSUBS 0.007378f
C141 B.n107 VSUBS 0.007378f
C142 B.n108 VSUBS 0.007378f
C143 B.n109 VSUBS 0.007378f
C144 B.n110 VSUBS 0.007378f
C145 B.n111 VSUBS 0.007378f
C146 B.n112 VSUBS 0.007378f
C147 B.n113 VSUBS 0.007378f
C148 B.n114 VSUBS 0.007378f
C149 B.n115 VSUBS 0.007378f
C150 B.n116 VSUBS 0.007378f
C151 B.n117 VSUBS 0.007378f
C152 B.n118 VSUBS 0.007378f
C153 B.n119 VSUBS 0.007378f
C154 B.n120 VSUBS 0.007378f
C155 B.n121 VSUBS 0.007378f
C156 B.n122 VSUBS 0.007378f
C157 B.n123 VSUBS 0.007378f
C158 B.n124 VSUBS 0.007378f
C159 B.n125 VSUBS 0.007378f
C160 B.n126 VSUBS 0.007378f
C161 B.n127 VSUBS 0.007378f
C162 B.n128 VSUBS 0.007378f
C163 B.n129 VSUBS 0.007378f
C164 B.n130 VSUBS 0.007378f
C165 B.n131 VSUBS 0.007378f
C166 B.n132 VSUBS 0.007378f
C167 B.n133 VSUBS 0.007378f
C168 B.n134 VSUBS 0.007378f
C169 B.n135 VSUBS 0.007378f
C170 B.n136 VSUBS 0.007378f
C171 B.n137 VSUBS 0.007378f
C172 B.n138 VSUBS 0.017649f
C173 B.n139 VSUBS 0.007378f
C174 B.n140 VSUBS 0.007378f
C175 B.n141 VSUBS 0.007378f
C176 B.n142 VSUBS 0.007378f
C177 B.n143 VSUBS 0.007378f
C178 B.n144 VSUBS 0.007378f
C179 B.n145 VSUBS 0.007378f
C180 B.n146 VSUBS 0.007378f
C181 B.n147 VSUBS 0.007378f
C182 B.n148 VSUBS 0.007378f
C183 B.n149 VSUBS 0.007378f
C184 B.n150 VSUBS 0.007378f
C185 B.n151 VSUBS 0.007378f
C186 B.n152 VSUBS 0.007378f
C187 B.n153 VSUBS 0.007378f
C188 B.n154 VSUBS 0.007378f
C189 B.n155 VSUBS 0.007378f
C190 B.n156 VSUBS 0.007378f
C191 B.n157 VSUBS 0.007378f
C192 B.n158 VSUBS 0.007378f
C193 B.n159 VSUBS 0.007378f
C194 B.n160 VSUBS 0.0051f
C195 B.n161 VSUBS 0.007378f
C196 B.n162 VSUBS 0.007378f
C197 B.n163 VSUBS 0.007378f
C198 B.n164 VSUBS 0.007378f
C199 B.n165 VSUBS 0.007378f
C200 B.t8 VSUBS 0.23938f
C201 B.t7 VSUBS 0.276304f
C202 B.t6 VSUBS 1.77104f
C203 B.n166 VSUBS 0.438265f
C204 B.n167 VSUBS 0.27719f
C205 B.n168 VSUBS 0.007378f
C206 B.n169 VSUBS 0.007378f
C207 B.n170 VSUBS 0.007378f
C208 B.n171 VSUBS 0.007378f
C209 B.n172 VSUBS 0.007378f
C210 B.n173 VSUBS 0.007378f
C211 B.n174 VSUBS 0.007378f
C212 B.n175 VSUBS 0.007378f
C213 B.n176 VSUBS 0.007378f
C214 B.n177 VSUBS 0.007378f
C215 B.n178 VSUBS 0.007378f
C216 B.n179 VSUBS 0.007378f
C217 B.n180 VSUBS 0.007378f
C218 B.n181 VSUBS 0.007378f
C219 B.n182 VSUBS 0.007378f
C220 B.n183 VSUBS 0.007378f
C221 B.n184 VSUBS 0.007378f
C222 B.n185 VSUBS 0.007378f
C223 B.n186 VSUBS 0.007378f
C224 B.n187 VSUBS 0.007378f
C225 B.n188 VSUBS 0.007378f
C226 B.n189 VSUBS 0.016767f
C227 B.n190 VSUBS 0.007378f
C228 B.n191 VSUBS 0.007378f
C229 B.n192 VSUBS 0.007378f
C230 B.n193 VSUBS 0.007378f
C231 B.n194 VSUBS 0.007378f
C232 B.n195 VSUBS 0.007378f
C233 B.n196 VSUBS 0.007378f
C234 B.n197 VSUBS 0.007378f
C235 B.n198 VSUBS 0.007378f
C236 B.n199 VSUBS 0.007378f
C237 B.n200 VSUBS 0.007378f
C238 B.n201 VSUBS 0.007378f
C239 B.n202 VSUBS 0.007378f
C240 B.n203 VSUBS 0.007378f
C241 B.n204 VSUBS 0.007378f
C242 B.n205 VSUBS 0.007378f
C243 B.n206 VSUBS 0.007378f
C244 B.n207 VSUBS 0.007378f
C245 B.n208 VSUBS 0.007378f
C246 B.n209 VSUBS 0.007378f
C247 B.n210 VSUBS 0.007378f
C248 B.n211 VSUBS 0.007378f
C249 B.n212 VSUBS 0.007378f
C250 B.n213 VSUBS 0.007378f
C251 B.n214 VSUBS 0.007378f
C252 B.n215 VSUBS 0.007378f
C253 B.n216 VSUBS 0.007378f
C254 B.n217 VSUBS 0.007378f
C255 B.n218 VSUBS 0.007378f
C256 B.n219 VSUBS 0.007378f
C257 B.n220 VSUBS 0.007378f
C258 B.n221 VSUBS 0.007378f
C259 B.n222 VSUBS 0.007378f
C260 B.n223 VSUBS 0.007378f
C261 B.n224 VSUBS 0.007378f
C262 B.n225 VSUBS 0.007378f
C263 B.n226 VSUBS 0.007378f
C264 B.n227 VSUBS 0.007378f
C265 B.n228 VSUBS 0.007378f
C266 B.n229 VSUBS 0.007378f
C267 B.n230 VSUBS 0.007378f
C268 B.n231 VSUBS 0.007378f
C269 B.n232 VSUBS 0.007378f
C270 B.n233 VSUBS 0.007378f
C271 B.n234 VSUBS 0.007378f
C272 B.n235 VSUBS 0.007378f
C273 B.n236 VSUBS 0.007378f
C274 B.n237 VSUBS 0.007378f
C275 B.n238 VSUBS 0.007378f
C276 B.n239 VSUBS 0.007378f
C277 B.n240 VSUBS 0.007378f
C278 B.n241 VSUBS 0.007378f
C279 B.n242 VSUBS 0.007378f
C280 B.n243 VSUBS 0.007378f
C281 B.n244 VSUBS 0.007378f
C282 B.n245 VSUBS 0.007378f
C283 B.n246 VSUBS 0.007378f
C284 B.n247 VSUBS 0.007378f
C285 B.n248 VSUBS 0.007378f
C286 B.n249 VSUBS 0.007378f
C287 B.n250 VSUBS 0.007378f
C288 B.n251 VSUBS 0.007378f
C289 B.n252 VSUBS 0.007378f
C290 B.n253 VSUBS 0.007378f
C291 B.n254 VSUBS 0.007378f
C292 B.n255 VSUBS 0.007378f
C293 B.n256 VSUBS 0.007378f
C294 B.n257 VSUBS 0.007378f
C295 B.n258 VSUBS 0.007378f
C296 B.n259 VSUBS 0.007378f
C297 B.n260 VSUBS 0.007378f
C298 B.n261 VSUBS 0.007378f
C299 B.n262 VSUBS 0.007378f
C300 B.n263 VSUBS 0.007378f
C301 B.n264 VSUBS 0.007378f
C302 B.n265 VSUBS 0.007378f
C303 B.n266 VSUBS 0.007378f
C304 B.n267 VSUBS 0.007378f
C305 B.n268 VSUBS 0.007378f
C306 B.n269 VSUBS 0.007378f
C307 B.n270 VSUBS 0.007378f
C308 B.n271 VSUBS 0.007378f
C309 B.n272 VSUBS 0.007378f
C310 B.n273 VSUBS 0.007378f
C311 B.n274 VSUBS 0.007378f
C312 B.n275 VSUBS 0.007378f
C313 B.n276 VSUBS 0.007378f
C314 B.n277 VSUBS 0.007378f
C315 B.n278 VSUBS 0.007378f
C316 B.n279 VSUBS 0.007378f
C317 B.n280 VSUBS 0.007378f
C318 B.n281 VSUBS 0.007378f
C319 B.n282 VSUBS 0.007378f
C320 B.n283 VSUBS 0.007378f
C321 B.n284 VSUBS 0.007378f
C322 B.n285 VSUBS 0.007378f
C323 B.n286 VSUBS 0.007378f
C324 B.n287 VSUBS 0.007378f
C325 B.n288 VSUBS 0.007378f
C326 B.n289 VSUBS 0.007378f
C327 B.n290 VSUBS 0.007378f
C328 B.n291 VSUBS 0.007378f
C329 B.n292 VSUBS 0.007378f
C330 B.n293 VSUBS 0.007378f
C331 B.n294 VSUBS 0.007378f
C332 B.n295 VSUBS 0.007378f
C333 B.n296 VSUBS 0.016767f
C334 B.n297 VSUBS 0.01752f
C335 B.n298 VSUBS 0.01752f
C336 B.n299 VSUBS 0.007378f
C337 B.n300 VSUBS 0.007378f
C338 B.n301 VSUBS 0.007378f
C339 B.n302 VSUBS 0.007378f
C340 B.n303 VSUBS 0.007378f
C341 B.n304 VSUBS 0.007378f
C342 B.n305 VSUBS 0.007378f
C343 B.n306 VSUBS 0.007378f
C344 B.n307 VSUBS 0.007378f
C345 B.n308 VSUBS 0.007378f
C346 B.n309 VSUBS 0.007378f
C347 B.n310 VSUBS 0.007378f
C348 B.n311 VSUBS 0.007378f
C349 B.n312 VSUBS 0.007378f
C350 B.n313 VSUBS 0.007378f
C351 B.n314 VSUBS 0.007378f
C352 B.n315 VSUBS 0.007378f
C353 B.n316 VSUBS 0.007378f
C354 B.n317 VSUBS 0.007378f
C355 B.n318 VSUBS 0.007378f
C356 B.n319 VSUBS 0.007378f
C357 B.n320 VSUBS 0.007378f
C358 B.n321 VSUBS 0.007378f
C359 B.n322 VSUBS 0.007378f
C360 B.n323 VSUBS 0.007378f
C361 B.n324 VSUBS 0.007378f
C362 B.n325 VSUBS 0.007378f
C363 B.n326 VSUBS 0.007378f
C364 B.n327 VSUBS 0.007378f
C365 B.n328 VSUBS 0.007378f
C366 B.n329 VSUBS 0.007378f
C367 B.n330 VSUBS 0.007378f
C368 B.n331 VSUBS 0.007378f
C369 B.n332 VSUBS 0.007378f
C370 B.n333 VSUBS 0.007378f
C371 B.n334 VSUBS 0.007378f
C372 B.n335 VSUBS 0.007378f
C373 B.n336 VSUBS 0.007378f
C374 B.n337 VSUBS 0.007378f
C375 B.n338 VSUBS 0.007378f
C376 B.n339 VSUBS 0.007378f
C377 B.n340 VSUBS 0.007378f
C378 B.n341 VSUBS 0.007378f
C379 B.n342 VSUBS 0.007378f
C380 B.n343 VSUBS 0.007378f
C381 B.n344 VSUBS 0.007378f
C382 B.n345 VSUBS 0.007378f
C383 B.n346 VSUBS 0.007378f
C384 B.n347 VSUBS 0.007378f
C385 B.n348 VSUBS 0.007378f
C386 B.n349 VSUBS 0.007378f
C387 B.n350 VSUBS 0.007378f
C388 B.n351 VSUBS 0.007378f
C389 B.n352 VSUBS 0.007378f
C390 B.n353 VSUBS 0.007378f
C391 B.n354 VSUBS 0.007378f
C392 B.n355 VSUBS 0.007378f
C393 B.n356 VSUBS 0.007378f
C394 B.n357 VSUBS 0.007378f
C395 B.n358 VSUBS 0.007378f
C396 B.n359 VSUBS 0.007378f
C397 B.n360 VSUBS 0.007378f
C398 B.n361 VSUBS 0.007378f
C399 B.n362 VSUBS 0.0051f
C400 B.n363 VSUBS 0.017095f
C401 B.n364 VSUBS 0.005968f
C402 B.n365 VSUBS 0.007378f
C403 B.n366 VSUBS 0.007378f
C404 B.n367 VSUBS 0.007378f
C405 B.n368 VSUBS 0.007378f
C406 B.n369 VSUBS 0.007378f
C407 B.n370 VSUBS 0.007378f
C408 B.n371 VSUBS 0.007378f
C409 B.n372 VSUBS 0.007378f
C410 B.n373 VSUBS 0.007378f
C411 B.n374 VSUBS 0.007378f
C412 B.n375 VSUBS 0.007378f
C413 B.t11 VSUBS 0.239383f
C414 B.t10 VSUBS 0.276307f
C415 B.t9 VSUBS 1.77104f
C416 B.n376 VSUBS 0.438262f
C417 B.n377 VSUBS 0.277187f
C418 B.n378 VSUBS 0.017095f
C419 B.n379 VSUBS 0.005968f
C420 B.n380 VSUBS 0.007378f
C421 B.n381 VSUBS 0.007378f
C422 B.n382 VSUBS 0.007378f
C423 B.n383 VSUBS 0.007378f
C424 B.n384 VSUBS 0.007378f
C425 B.n385 VSUBS 0.007378f
C426 B.n386 VSUBS 0.007378f
C427 B.n387 VSUBS 0.007378f
C428 B.n388 VSUBS 0.007378f
C429 B.n389 VSUBS 0.007378f
C430 B.n390 VSUBS 0.007378f
C431 B.n391 VSUBS 0.007378f
C432 B.n392 VSUBS 0.007378f
C433 B.n393 VSUBS 0.007378f
C434 B.n394 VSUBS 0.007378f
C435 B.n395 VSUBS 0.007378f
C436 B.n396 VSUBS 0.007378f
C437 B.n397 VSUBS 0.007378f
C438 B.n398 VSUBS 0.007378f
C439 B.n399 VSUBS 0.007378f
C440 B.n400 VSUBS 0.007378f
C441 B.n401 VSUBS 0.007378f
C442 B.n402 VSUBS 0.007378f
C443 B.n403 VSUBS 0.007378f
C444 B.n404 VSUBS 0.007378f
C445 B.n405 VSUBS 0.007378f
C446 B.n406 VSUBS 0.007378f
C447 B.n407 VSUBS 0.007378f
C448 B.n408 VSUBS 0.007378f
C449 B.n409 VSUBS 0.007378f
C450 B.n410 VSUBS 0.007378f
C451 B.n411 VSUBS 0.007378f
C452 B.n412 VSUBS 0.007378f
C453 B.n413 VSUBS 0.007378f
C454 B.n414 VSUBS 0.007378f
C455 B.n415 VSUBS 0.007378f
C456 B.n416 VSUBS 0.007378f
C457 B.n417 VSUBS 0.007378f
C458 B.n418 VSUBS 0.007378f
C459 B.n419 VSUBS 0.007378f
C460 B.n420 VSUBS 0.007378f
C461 B.n421 VSUBS 0.007378f
C462 B.n422 VSUBS 0.007378f
C463 B.n423 VSUBS 0.007378f
C464 B.n424 VSUBS 0.007378f
C465 B.n425 VSUBS 0.007378f
C466 B.n426 VSUBS 0.007378f
C467 B.n427 VSUBS 0.007378f
C468 B.n428 VSUBS 0.007378f
C469 B.n429 VSUBS 0.007378f
C470 B.n430 VSUBS 0.007378f
C471 B.n431 VSUBS 0.007378f
C472 B.n432 VSUBS 0.007378f
C473 B.n433 VSUBS 0.007378f
C474 B.n434 VSUBS 0.007378f
C475 B.n435 VSUBS 0.007378f
C476 B.n436 VSUBS 0.007378f
C477 B.n437 VSUBS 0.007378f
C478 B.n438 VSUBS 0.007378f
C479 B.n439 VSUBS 0.007378f
C480 B.n440 VSUBS 0.007378f
C481 B.n441 VSUBS 0.007378f
C482 B.n442 VSUBS 0.007378f
C483 B.n443 VSUBS 0.007378f
C484 B.n444 VSUBS 0.007378f
C485 B.n445 VSUBS 0.016638f
C486 B.n446 VSUBS 0.01752f
C487 B.n447 VSUBS 0.016767f
C488 B.n448 VSUBS 0.007378f
C489 B.n449 VSUBS 0.007378f
C490 B.n450 VSUBS 0.007378f
C491 B.n451 VSUBS 0.007378f
C492 B.n452 VSUBS 0.007378f
C493 B.n453 VSUBS 0.007378f
C494 B.n454 VSUBS 0.007378f
C495 B.n455 VSUBS 0.007378f
C496 B.n456 VSUBS 0.007378f
C497 B.n457 VSUBS 0.007378f
C498 B.n458 VSUBS 0.007378f
C499 B.n459 VSUBS 0.007378f
C500 B.n460 VSUBS 0.007378f
C501 B.n461 VSUBS 0.007378f
C502 B.n462 VSUBS 0.007378f
C503 B.n463 VSUBS 0.007378f
C504 B.n464 VSUBS 0.007378f
C505 B.n465 VSUBS 0.007378f
C506 B.n466 VSUBS 0.007378f
C507 B.n467 VSUBS 0.007378f
C508 B.n468 VSUBS 0.007378f
C509 B.n469 VSUBS 0.007378f
C510 B.n470 VSUBS 0.007378f
C511 B.n471 VSUBS 0.007378f
C512 B.n472 VSUBS 0.007378f
C513 B.n473 VSUBS 0.007378f
C514 B.n474 VSUBS 0.007378f
C515 B.n475 VSUBS 0.007378f
C516 B.n476 VSUBS 0.007378f
C517 B.n477 VSUBS 0.007378f
C518 B.n478 VSUBS 0.007378f
C519 B.n479 VSUBS 0.007378f
C520 B.n480 VSUBS 0.007378f
C521 B.n481 VSUBS 0.007378f
C522 B.n482 VSUBS 0.007378f
C523 B.n483 VSUBS 0.007378f
C524 B.n484 VSUBS 0.007378f
C525 B.n485 VSUBS 0.007378f
C526 B.n486 VSUBS 0.007378f
C527 B.n487 VSUBS 0.007378f
C528 B.n488 VSUBS 0.007378f
C529 B.n489 VSUBS 0.007378f
C530 B.n490 VSUBS 0.007378f
C531 B.n491 VSUBS 0.007378f
C532 B.n492 VSUBS 0.007378f
C533 B.n493 VSUBS 0.007378f
C534 B.n494 VSUBS 0.007378f
C535 B.n495 VSUBS 0.007378f
C536 B.n496 VSUBS 0.007378f
C537 B.n497 VSUBS 0.007378f
C538 B.n498 VSUBS 0.007378f
C539 B.n499 VSUBS 0.007378f
C540 B.n500 VSUBS 0.007378f
C541 B.n501 VSUBS 0.007378f
C542 B.n502 VSUBS 0.007378f
C543 B.n503 VSUBS 0.007378f
C544 B.n504 VSUBS 0.007378f
C545 B.n505 VSUBS 0.007378f
C546 B.n506 VSUBS 0.007378f
C547 B.n507 VSUBS 0.007378f
C548 B.n508 VSUBS 0.007378f
C549 B.n509 VSUBS 0.007378f
C550 B.n510 VSUBS 0.007378f
C551 B.n511 VSUBS 0.007378f
C552 B.n512 VSUBS 0.007378f
C553 B.n513 VSUBS 0.007378f
C554 B.n514 VSUBS 0.007378f
C555 B.n515 VSUBS 0.007378f
C556 B.n516 VSUBS 0.007378f
C557 B.n517 VSUBS 0.007378f
C558 B.n518 VSUBS 0.007378f
C559 B.n519 VSUBS 0.007378f
C560 B.n520 VSUBS 0.007378f
C561 B.n521 VSUBS 0.007378f
C562 B.n522 VSUBS 0.007378f
C563 B.n523 VSUBS 0.007378f
C564 B.n524 VSUBS 0.007378f
C565 B.n525 VSUBS 0.007378f
C566 B.n526 VSUBS 0.007378f
C567 B.n527 VSUBS 0.007378f
C568 B.n528 VSUBS 0.007378f
C569 B.n529 VSUBS 0.007378f
C570 B.n530 VSUBS 0.007378f
C571 B.n531 VSUBS 0.007378f
C572 B.n532 VSUBS 0.007378f
C573 B.n533 VSUBS 0.007378f
C574 B.n534 VSUBS 0.007378f
C575 B.n535 VSUBS 0.007378f
C576 B.n536 VSUBS 0.007378f
C577 B.n537 VSUBS 0.007378f
C578 B.n538 VSUBS 0.007378f
C579 B.n539 VSUBS 0.007378f
C580 B.n540 VSUBS 0.007378f
C581 B.n541 VSUBS 0.007378f
C582 B.n542 VSUBS 0.007378f
C583 B.n543 VSUBS 0.007378f
C584 B.n544 VSUBS 0.007378f
C585 B.n545 VSUBS 0.007378f
C586 B.n546 VSUBS 0.007378f
C587 B.n547 VSUBS 0.007378f
C588 B.n548 VSUBS 0.007378f
C589 B.n549 VSUBS 0.007378f
C590 B.n550 VSUBS 0.007378f
C591 B.n551 VSUBS 0.007378f
C592 B.n552 VSUBS 0.007378f
C593 B.n553 VSUBS 0.007378f
C594 B.n554 VSUBS 0.007378f
C595 B.n555 VSUBS 0.007378f
C596 B.n556 VSUBS 0.007378f
C597 B.n557 VSUBS 0.007378f
C598 B.n558 VSUBS 0.007378f
C599 B.n559 VSUBS 0.007378f
C600 B.n560 VSUBS 0.007378f
C601 B.n561 VSUBS 0.007378f
C602 B.n562 VSUBS 0.007378f
C603 B.n563 VSUBS 0.007378f
C604 B.n564 VSUBS 0.007378f
C605 B.n565 VSUBS 0.007378f
C606 B.n566 VSUBS 0.007378f
C607 B.n567 VSUBS 0.007378f
C608 B.n568 VSUBS 0.007378f
C609 B.n569 VSUBS 0.007378f
C610 B.n570 VSUBS 0.007378f
C611 B.n571 VSUBS 0.007378f
C612 B.n572 VSUBS 0.007378f
C613 B.n573 VSUBS 0.007378f
C614 B.n574 VSUBS 0.007378f
C615 B.n575 VSUBS 0.007378f
C616 B.n576 VSUBS 0.007378f
C617 B.n577 VSUBS 0.007378f
C618 B.n578 VSUBS 0.007378f
C619 B.n579 VSUBS 0.007378f
C620 B.n580 VSUBS 0.007378f
C621 B.n581 VSUBS 0.007378f
C622 B.n582 VSUBS 0.007378f
C623 B.n583 VSUBS 0.007378f
C624 B.n584 VSUBS 0.007378f
C625 B.n585 VSUBS 0.007378f
C626 B.n586 VSUBS 0.007378f
C627 B.n587 VSUBS 0.007378f
C628 B.n588 VSUBS 0.007378f
C629 B.n589 VSUBS 0.007378f
C630 B.n590 VSUBS 0.007378f
C631 B.n591 VSUBS 0.007378f
C632 B.n592 VSUBS 0.007378f
C633 B.n593 VSUBS 0.007378f
C634 B.n594 VSUBS 0.007378f
C635 B.n595 VSUBS 0.007378f
C636 B.n596 VSUBS 0.007378f
C637 B.n597 VSUBS 0.007378f
C638 B.n598 VSUBS 0.007378f
C639 B.n599 VSUBS 0.007378f
C640 B.n600 VSUBS 0.007378f
C641 B.n601 VSUBS 0.007378f
C642 B.n602 VSUBS 0.007378f
C643 B.n603 VSUBS 0.007378f
C644 B.n604 VSUBS 0.007378f
C645 B.n605 VSUBS 0.007378f
C646 B.n606 VSUBS 0.007378f
C647 B.n607 VSUBS 0.007378f
C648 B.n608 VSUBS 0.007378f
C649 B.n609 VSUBS 0.007378f
C650 B.n610 VSUBS 0.007378f
C651 B.n611 VSUBS 0.007378f
C652 B.n612 VSUBS 0.007378f
C653 B.n613 VSUBS 0.016767f
C654 B.n614 VSUBS 0.016767f
C655 B.n615 VSUBS 0.01752f
C656 B.n616 VSUBS 0.007378f
C657 B.n617 VSUBS 0.007378f
C658 B.n618 VSUBS 0.007378f
C659 B.n619 VSUBS 0.007378f
C660 B.n620 VSUBS 0.007378f
C661 B.n621 VSUBS 0.007378f
C662 B.n622 VSUBS 0.007378f
C663 B.n623 VSUBS 0.007378f
C664 B.n624 VSUBS 0.007378f
C665 B.n625 VSUBS 0.007378f
C666 B.n626 VSUBS 0.007378f
C667 B.n627 VSUBS 0.007378f
C668 B.n628 VSUBS 0.007378f
C669 B.n629 VSUBS 0.007378f
C670 B.n630 VSUBS 0.007378f
C671 B.n631 VSUBS 0.007378f
C672 B.n632 VSUBS 0.007378f
C673 B.n633 VSUBS 0.007378f
C674 B.n634 VSUBS 0.007378f
C675 B.n635 VSUBS 0.007378f
C676 B.n636 VSUBS 0.007378f
C677 B.n637 VSUBS 0.007378f
C678 B.n638 VSUBS 0.007378f
C679 B.n639 VSUBS 0.007378f
C680 B.n640 VSUBS 0.007378f
C681 B.n641 VSUBS 0.007378f
C682 B.n642 VSUBS 0.007378f
C683 B.n643 VSUBS 0.007378f
C684 B.n644 VSUBS 0.007378f
C685 B.n645 VSUBS 0.007378f
C686 B.n646 VSUBS 0.007378f
C687 B.n647 VSUBS 0.007378f
C688 B.n648 VSUBS 0.007378f
C689 B.n649 VSUBS 0.007378f
C690 B.n650 VSUBS 0.007378f
C691 B.n651 VSUBS 0.007378f
C692 B.n652 VSUBS 0.007378f
C693 B.n653 VSUBS 0.007378f
C694 B.n654 VSUBS 0.007378f
C695 B.n655 VSUBS 0.007378f
C696 B.n656 VSUBS 0.007378f
C697 B.n657 VSUBS 0.007378f
C698 B.n658 VSUBS 0.007378f
C699 B.n659 VSUBS 0.007378f
C700 B.n660 VSUBS 0.007378f
C701 B.n661 VSUBS 0.007378f
C702 B.n662 VSUBS 0.007378f
C703 B.n663 VSUBS 0.007378f
C704 B.n664 VSUBS 0.007378f
C705 B.n665 VSUBS 0.007378f
C706 B.n666 VSUBS 0.007378f
C707 B.n667 VSUBS 0.007378f
C708 B.n668 VSUBS 0.007378f
C709 B.n669 VSUBS 0.007378f
C710 B.n670 VSUBS 0.007378f
C711 B.n671 VSUBS 0.007378f
C712 B.n672 VSUBS 0.007378f
C713 B.n673 VSUBS 0.007378f
C714 B.n674 VSUBS 0.007378f
C715 B.n675 VSUBS 0.007378f
C716 B.n676 VSUBS 0.007378f
C717 B.n677 VSUBS 0.007378f
C718 B.n678 VSUBS 0.007378f
C719 B.n679 VSUBS 0.0051f
C720 B.n680 VSUBS 0.007378f
C721 B.n681 VSUBS 0.007378f
C722 B.n682 VSUBS 0.005968f
C723 B.n683 VSUBS 0.007378f
C724 B.n684 VSUBS 0.007378f
C725 B.n685 VSUBS 0.007378f
C726 B.n686 VSUBS 0.007378f
C727 B.n687 VSUBS 0.007378f
C728 B.n688 VSUBS 0.007378f
C729 B.n689 VSUBS 0.007378f
C730 B.n690 VSUBS 0.007378f
C731 B.n691 VSUBS 0.007378f
C732 B.n692 VSUBS 0.007378f
C733 B.n693 VSUBS 0.007378f
C734 B.n694 VSUBS 0.005968f
C735 B.n695 VSUBS 0.017095f
C736 B.n696 VSUBS 0.0051f
C737 B.n697 VSUBS 0.007378f
C738 B.n698 VSUBS 0.007378f
C739 B.n699 VSUBS 0.007378f
C740 B.n700 VSUBS 0.007378f
C741 B.n701 VSUBS 0.007378f
C742 B.n702 VSUBS 0.007378f
C743 B.n703 VSUBS 0.007378f
C744 B.n704 VSUBS 0.007378f
C745 B.n705 VSUBS 0.007378f
C746 B.n706 VSUBS 0.007378f
C747 B.n707 VSUBS 0.007378f
C748 B.n708 VSUBS 0.007378f
C749 B.n709 VSUBS 0.007378f
C750 B.n710 VSUBS 0.007378f
C751 B.n711 VSUBS 0.007378f
C752 B.n712 VSUBS 0.007378f
C753 B.n713 VSUBS 0.007378f
C754 B.n714 VSUBS 0.007378f
C755 B.n715 VSUBS 0.007378f
C756 B.n716 VSUBS 0.007378f
C757 B.n717 VSUBS 0.007378f
C758 B.n718 VSUBS 0.007378f
C759 B.n719 VSUBS 0.007378f
C760 B.n720 VSUBS 0.007378f
C761 B.n721 VSUBS 0.007378f
C762 B.n722 VSUBS 0.007378f
C763 B.n723 VSUBS 0.007378f
C764 B.n724 VSUBS 0.007378f
C765 B.n725 VSUBS 0.007378f
C766 B.n726 VSUBS 0.007378f
C767 B.n727 VSUBS 0.007378f
C768 B.n728 VSUBS 0.007378f
C769 B.n729 VSUBS 0.007378f
C770 B.n730 VSUBS 0.007378f
C771 B.n731 VSUBS 0.007378f
C772 B.n732 VSUBS 0.007378f
C773 B.n733 VSUBS 0.007378f
C774 B.n734 VSUBS 0.007378f
C775 B.n735 VSUBS 0.007378f
C776 B.n736 VSUBS 0.007378f
C777 B.n737 VSUBS 0.007378f
C778 B.n738 VSUBS 0.007378f
C779 B.n739 VSUBS 0.007378f
C780 B.n740 VSUBS 0.007378f
C781 B.n741 VSUBS 0.007378f
C782 B.n742 VSUBS 0.007378f
C783 B.n743 VSUBS 0.007378f
C784 B.n744 VSUBS 0.007378f
C785 B.n745 VSUBS 0.007378f
C786 B.n746 VSUBS 0.007378f
C787 B.n747 VSUBS 0.007378f
C788 B.n748 VSUBS 0.007378f
C789 B.n749 VSUBS 0.007378f
C790 B.n750 VSUBS 0.007378f
C791 B.n751 VSUBS 0.007378f
C792 B.n752 VSUBS 0.007378f
C793 B.n753 VSUBS 0.007378f
C794 B.n754 VSUBS 0.007378f
C795 B.n755 VSUBS 0.007378f
C796 B.n756 VSUBS 0.007378f
C797 B.n757 VSUBS 0.007378f
C798 B.n758 VSUBS 0.007378f
C799 B.n759 VSUBS 0.007378f
C800 B.n760 VSUBS 0.01752f
C801 B.n761 VSUBS 0.01752f
C802 B.n762 VSUBS 0.016767f
C803 B.n763 VSUBS 0.007378f
C804 B.n764 VSUBS 0.007378f
C805 B.n765 VSUBS 0.007378f
C806 B.n766 VSUBS 0.007378f
C807 B.n767 VSUBS 0.007378f
C808 B.n768 VSUBS 0.007378f
C809 B.n769 VSUBS 0.007378f
C810 B.n770 VSUBS 0.007378f
C811 B.n771 VSUBS 0.007378f
C812 B.n772 VSUBS 0.007378f
C813 B.n773 VSUBS 0.007378f
C814 B.n774 VSUBS 0.007378f
C815 B.n775 VSUBS 0.007378f
C816 B.n776 VSUBS 0.007378f
C817 B.n777 VSUBS 0.007378f
C818 B.n778 VSUBS 0.007378f
C819 B.n779 VSUBS 0.007378f
C820 B.n780 VSUBS 0.007378f
C821 B.n781 VSUBS 0.007378f
C822 B.n782 VSUBS 0.007378f
C823 B.n783 VSUBS 0.007378f
C824 B.n784 VSUBS 0.007378f
C825 B.n785 VSUBS 0.007378f
C826 B.n786 VSUBS 0.007378f
C827 B.n787 VSUBS 0.007378f
C828 B.n788 VSUBS 0.007378f
C829 B.n789 VSUBS 0.007378f
C830 B.n790 VSUBS 0.007378f
C831 B.n791 VSUBS 0.007378f
C832 B.n792 VSUBS 0.007378f
C833 B.n793 VSUBS 0.007378f
C834 B.n794 VSUBS 0.007378f
C835 B.n795 VSUBS 0.007378f
C836 B.n796 VSUBS 0.007378f
C837 B.n797 VSUBS 0.007378f
C838 B.n798 VSUBS 0.007378f
C839 B.n799 VSUBS 0.007378f
C840 B.n800 VSUBS 0.007378f
C841 B.n801 VSUBS 0.007378f
C842 B.n802 VSUBS 0.007378f
C843 B.n803 VSUBS 0.007378f
C844 B.n804 VSUBS 0.007378f
C845 B.n805 VSUBS 0.007378f
C846 B.n806 VSUBS 0.007378f
C847 B.n807 VSUBS 0.007378f
C848 B.n808 VSUBS 0.007378f
C849 B.n809 VSUBS 0.007378f
C850 B.n810 VSUBS 0.007378f
C851 B.n811 VSUBS 0.007378f
C852 B.n812 VSUBS 0.007378f
C853 B.n813 VSUBS 0.007378f
C854 B.n814 VSUBS 0.007378f
C855 B.n815 VSUBS 0.007378f
C856 B.n816 VSUBS 0.007378f
C857 B.n817 VSUBS 0.007378f
C858 B.n818 VSUBS 0.007378f
C859 B.n819 VSUBS 0.007378f
C860 B.n820 VSUBS 0.007378f
C861 B.n821 VSUBS 0.007378f
C862 B.n822 VSUBS 0.007378f
C863 B.n823 VSUBS 0.007378f
C864 B.n824 VSUBS 0.007378f
C865 B.n825 VSUBS 0.007378f
C866 B.n826 VSUBS 0.007378f
C867 B.n827 VSUBS 0.007378f
C868 B.n828 VSUBS 0.007378f
C869 B.n829 VSUBS 0.007378f
C870 B.n830 VSUBS 0.007378f
C871 B.n831 VSUBS 0.007378f
C872 B.n832 VSUBS 0.007378f
C873 B.n833 VSUBS 0.007378f
C874 B.n834 VSUBS 0.007378f
C875 B.n835 VSUBS 0.007378f
C876 B.n836 VSUBS 0.007378f
C877 B.n837 VSUBS 0.007378f
C878 B.n838 VSUBS 0.007378f
C879 B.n839 VSUBS 0.007378f
C880 B.n840 VSUBS 0.007378f
C881 B.n841 VSUBS 0.007378f
C882 B.n842 VSUBS 0.007378f
C883 B.n843 VSUBS 0.009628f
C884 B.n844 VSUBS 0.010256f
C885 B.n845 VSUBS 0.020396f
C886 VDD2.t0 VSUBS 0.27321f
C887 VDD2.t1 VSUBS 0.27321f
C888 VDD2.n0 VSUBS 2.15886f
C889 VDD2.t7 VSUBS 0.27321f
C890 VDD2.t5 VSUBS 0.27321f
C891 VDD2.n1 VSUBS 2.15886f
C892 VDD2.n2 VSUBS 4.39272f
C893 VDD2.t6 VSUBS 0.27321f
C894 VDD2.t2 VSUBS 0.27321f
C895 VDD2.n3 VSUBS 2.14225f
C896 VDD2.n4 VSUBS 3.6792f
C897 VDD2.t4 VSUBS 0.27321f
C898 VDD2.t3 VSUBS 0.27321f
C899 VDD2.n5 VSUBS 2.15881f
C900 VN.n0 VSUBS 0.035625f
C901 VN.t2 VSUBS 2.71065f
C902 VN.n1 VSUBS 0.054641f
C903 VN.n2 VSUBS 0.02702f
C904 VN.n3 VSUBS 0.032619f
C905 VN.n4 VSUBS 0.02702f
C906 VN.n5 VSUBS 0.039616f
C907 VN.n6 VSUBS 0.286386f
C908 VN.t6 VSUBS 2.71065f
C909 VN.t7 VSUBS 2.98352f
C910 VN.n7 VSUBS 1.00067f
C911 VN.n8 VSUBS 1.04316f
C912 VN.n9 VSUBS 0.043614f
C913 VN.n10 VSUBS 0.05061f
C914 VN.n11 VSUBS 0.02702f
C915 VN.n12 VSUBS 0.02702f
C916 VN.n13 VSUBS 0.02702f
C917 VN.n14 VSUBS 0.039616f
C918 VN.n15 VSUBS 0.05061f
C919 VN.t0 VSUBS 2.71065f
C920 VN.n16 VSUBS 0.952855f
C921 VN.n17 VSUBS 0.043614f
C922 VN.n18 VSUBS 0.02702f
C923 VN.n19 VSUBS 0.02702f
C924 VN.n20 VSUBS 0.02702f
C925 VN.n21 VSUBS 0.05061f
C926 VN.n22 VSUBS 0.053019f
C927 VN.n23 VSUBS 0.022181f
C928 VN.n24 VSUBS 0.02702f
C929 VN.n25 VSUBS 0.02702f
C930 VN.n26 VSUBS 0.02702f
C931 VN.n27 VSUBS 0.05061f
C932 VN.n28 VSUBS 0.02962f
C933 VN.n29 VSUBS 1.04539f
C934 VN.n30 VSUBS 0.050776f
C935 VN.n31 VSUBS 0.035625f
C936 VN.t1 VSUBS 2.71065f
C937 VN.n32 VSUBS 0.054641f
C938 VN.n33 VSUBS 0.02702f
C939 VN.n34 VSUBS 0.032619f
C940 VN.n35 VSUBS 0.02702f
C941 VN.t5 VSUBS 2.71065f
C942 VN.n36 VSUBS 0.952855f
C943 VN.n37 VSUBS 0.039616f
C944 VN.n38 VSUBS 0.286386f
C945 VN.t3 VSUBS 2.71065f
C946 VN.t4 VSUBS 2.98352f
C947 VN.n39 VSUBS 1.00067f
C948 VN.n40 VSUBS 1.04316f
C949 VN.n41 VSUBS 0.043614f
C950 VN.n42 VSUBS 0.05061f
C951 VN.n43 VSUBS 0.02702f
C952 VN.n44 VSUBS 0.02702f
C953 VN.n45 VSUBS 0.02702f
C954 VN.n46 VSUBS 0.039616f
C955 VN.n47 VSUBS 0.05061f
C956 VN.n48 VSUBS 0.043614f
C957 VN.n49 VSUBS 0.02702f
C958 VN.n50 VSUBS 0.02702f
C959 VN.n51 VSUBS 0.02702f
C960 VN.n52 VSUBS 0.05061f
C961 VN.n53 VSUBS 0.053019f
C962 VN.n54 VSUBS 0.022181f
C963 VN.n55 VSUBS 0.02702f
C964 VN.n56 VSUBS 0.02702f
C965 VN.n57 VSUBS 0.02702f
C966 VN.n58 VSUBS 0.05061f
C967 VN.n59 VSUBS 0.02962f
C968 VN.n60 VSUBS 1.04539f
C969 VN.n61 VSUBS 1.64847f
C970 VDD1.t1 VSUBS 0.275923f
C971 VDD1.t3 VSUBS 0.275923f
C972 VDD1.n0 VSUBS 2.1819f
C973 VDD1.t6 VSUBS 0.275923f
C974 VDD1.t7 VSUBS 0.275923f
C975 VDD1.n1 VSUBS 2.1803f
C976 VDD1.t0 VSUBS 0.275923f
C977 VDD1.t2 VSUBS 0.275923f
C978 VDD1.n2 VSUBS 2.1803f
C979 VDD1.n3 VSUBS 4.49331f
C980 VDD1.t4 VSUBS 0.275923f
C981 VDD1.t5 VSUBS 0.275923f
C982 VDD1.n4 VSUBS 2.16352f
C983 VDD1.n5 VSUBS 3.74987f
C984 VTAIL.t7 VSUBS 0.252073f
C985 VTAIL.t0 VSUBS 0.252073f
C986 VTAIL.n0 VSUBS 1.82794f
C987 VTAIL.n1 VSUBS 0.829298f
C988 VTAIL.n2 VSUBS 0.0266f
C989 VTAIL.n3 VSUBS 0.025077f
C990 VTAIL.n4 VSUBS 0.013476f
C991 VTAIL.n5 VSUBS 0.031851f
C992 VTAIL.n6 VSUBS 0.014268f
C993 VTAIL.n7 VSUBS 0.025077f
C994 VTAIL.n8 VSUBS 0.013476f
C995 VTAIL.n9 VSUBS 0.031851f
C996 VTAIL.n10 VSUBS 0.014268f
C997 VTAIL.n11 VSUBS 0.025077f
C998 VTAIL.n12 VSUBS 0.013476f
C999 VTAIL.n13 VSUBS 0.031851f
C1000 VTAIL.n14 VSUBS 0.014268f
C1001 VTAIL.n15 VSUBS 0.025077f
C1002 VTAIL.n16 VSUBS 0.013476f
C1003 VTAIL.n17 VSUBS 0.031851f
C1004 VTAIL.n18 VSUBS 0.014268f
C1005 VTAIL.n19 VSUBS 0.025077f
C1006 VTAIL.n20 VSUBS 0.013476f
C1007 VTAIL.n21 VSUBS 0.031851f
C1008 VTAIL.n22 VSUBS 0.014268f
C1009 VTAIL.n23 VSUBS 0.205662f
C1010 VTAIL.t5 VSUBS 0.068695f
C1011 VTAIL.n24 VSUBS 0.023889f
C1012 VTAIL.n25 VSUBS 0.02396f
C1013 VTAIL.n26 VSUBS 0.013476f
C1014 VTAIL.n27 VSUBS 1.31126f
C1015 VTAIL.n28 VSUBS 0.025077f
C1016 VTAIL.n29 VSUBS 0.013476f
C1017 VTAIL.n30 VSUBS 0.014268f
C1018 VTAIL.n31 VSUBS 0.031851f
C1019 VTAIL.n32 VSUBS 0.031851f
C1020 VTAIL.n33 VSUBS 0.014268f
C1021 VTAIL.n34 VSUBS 0.013476f
C1022 VTAIL.n35 VSUBS 0.025077f
C1023 VTAIL.n36 VSUBS 0.025077f
C1024 VTAIL.n37 VSUBS 0.013476f
C1025 VTAIL.n38 VSUBS 0.014268f
C1026 VTAIL.n39 VSUBS 0.031851f
C1027 VTAIL.n40 VSUBS 0.031851f
C1028 VTAIL.n41 VSUBS 0.031851f
C1029 VTAIL.n42 VSUBS 0.014268f
C1030 VTAIL.n43 VSUBS 0.013476f
C1031 VTAIL.n44 VSUBS 0.025077f
C1032 VTAIL.n45 VSUBS 0.025077f
C1033 VTAIL.n46 VSUBS 0.013476f
C1034 VTAIL.n47 VSUBS 0.013872f
C1035 VTAIL.n48 VSUBS 0.013872f
C1036 VTAIL.n49 VSUBS 0.031851f
C1037 VTAIL.n50 VSUBS 0.031851f
C1038 VTAIL.n51 VSUBS 0.014268f
C1039 VTAIL.n52 VSUBS 0.013476f
C1040 VTAIL.n53 VSUBS 0.025077f
C1041 VTAIL.n54 VSUBS 0.025077f
C1042 VTAIL.n55 VSUBS 0.013476f
C1043 VTAIL.n56 VSUBS 0.014268f
C1044 VTAIL.n57 VSUBS 0.031851f
C1045 VTAIL.n58 VSUBS 0.031851f
C1046 VTAIL.n59 VSUBS 0.014268f
C1047 VTAIL.n60 VSUBS 0.013476f
C1048 VTAIL.n61 VSUBS 0.025077f
C1049 VTAIL.n62 VSUBS 0.025077f
C1050 VTAIL.n63 VSUBS 0.013476f
C1051 VTAIL.n64 VSUBS 0.014268f
C1052 VTAIL.n65 VSUBS 0.031851f
C1053 VTAIL.n66 VSUBS 0.073855f
C1054 VTAIL.n67 VSUBS 0.014268f
C1055 VTAIL.n68 VSUBS 0.013476f
C1056 VTAIL.n69 VSUBS 0.053854f
C1057 VTAIL.n70 VSUBS 0.036866f
C1058 VTAIL.n71 VSUBS 0.281372f
C1059 VTAIL.n72 VSUBS 0.0266f
C1060 VTAIL.n73 VSUBS 0.025077f
C1061 VTAIL.n74 VSUBS 0.013476f
C1062 VTAIL.n75 VSUBS 0.031851f
C1063 VTAIL.n76 VSUBS 0.014268f
C1064 VTAIL.n77 VSUBS 0.025077f
C1065 VTAIL.n78 VSUBS 0.013476f
C1066 VTAIL.n79 VSUBS 0.031851f
C1067 VTAIL.n80 VSUBS 0.014268f
C1068 VTAIL.n81 VSUBS 0.025077f
C1069 VTAIL.n82 VSUBS 0.013476f
C1070 VTAIL.n83 VSUBS 0.031851f
C1071 VTAIL.n84 VSUBS 0.014268f
C1072 VTAIL.n85 VSUBS 0.025077f
C1073 VTAIL.n86 VSUBS 0.013476f
C1074 VTAIL.n87 VSUBS 0.031851f
C1075 VTAIL.n88 VSUBS 0.014268f
C1076 VTAIL.n89 VSUBS 0.025077f
C1077 VTAIL.n90 VSUBS 0.013476f
C1078 VTAIL.n91 VSUBS 0.031851f
C1079 VTAIL.n92 VSUBS 0.014268f
C1080 VTAIL.n93 VSUBS 0.205662f
C1081 VTAIL.t10 VSUBS 0.068695f
C1082 VTAIL.n94 VSUBS 0.023889f
C1083 VTAIL.n95 VSUBS 0.02396f
C1084 VTAIL.n96 VSUBS 0.013476f
C1085 VTAIL.n97 VSUBS 1.31126f
C1086 VTAIL.n98 VSUBS 0.025077f
C1087 VTAIL.n99 VSUBS 0.013476f
C1088 VTAIL.n100 VSUBS 0.014268f
C1089 VTAIL.n101 VSUBS 0.031851f
C1090 VTAIL.n102 VSUBS 0.031851f
C1091 VTAIL.n103 VSUBS 0.014268f
C1092 VTAIL.n104 VSUBS 0.013476f
C1093 VTAIL.n105 VSUBS 0.025077f
C1094 VTAIL.n106 VSUBS 0.025077f
C1095 VTAIL.n107 VSUBS 0.013476f
C1096 VTAIL.n108 VSUBS 0.014268f
C1097 VTAIL.n109 VSUBS 0.031851f
C1098 VTAIL.n110 VSUBS 0.031851f
C1099 VTAIL.n111 VSUBS 0.031851f
C1100 VTAIL.n112 VSUBS 0.014268f
C1101 VTAIL.n113 VSUBS 0.013476f
C1102 VTAIL.n114 VSUBS 0.025077f
C1103 VTAIL.n115 VSUBS 0.025077f
C1104 VTAIL.n116 VSUBS 0.013476f
C1105 VTAIL.n117 VSUBS 0.013872f
C1106 VTAIL.n118 VSUBS 0.013872f
C1107 VTAIL.n119 VSUBS 0.031851f
C1108 VTAIL.n120 VSUBS 0.031851f
C1109 VTAIL.n121 VSUBS 0.014268f
C1110 VTAIL.n122 VSUBS 0.013476f
C1111 VTAIL.n123 VSUBS 0.025077f
C1112 VTAIL.n124 VSUBS 0.025077f
C1113 VTAIL.n125 VSUBS 0.013476f
C1114 VTAIL.n126 VSUBS 0.014268f
C1115 VTAIL.n127 VSUBS 0.031851f
C1116 VTAIL.n128 VSUBS 0.031851f
C1117 VTAIL.n129 VSUBS 0.014268f
C1118 VTAIL.n130 VSUBS 0.013476f
C1119 VTAIL.n131 VSUBS 0.025077f
C1120 VTAIL.n132 VSUBS 0.025077f
C1121 VTAIL.n133 VSUBS 0.013476f
C1122 VTAIL.n134 VSUBS 0.014268f
C1123 VTAIL.n135 VSUBS 0.031851f
C1124 VTAIL.n136 VSUBS 0.073855f
C1125 VTAIL.n137 VSUBS 0.014268f
C1126 VTAIL.n138 VSUBS 0.013476f
C1127 VTAIL.n139 VSUBS 0.053854f
C1128 VTAIL.n140 VSUBS 0.036866f
C1129 VTAIL.n141 VSUBS 0.281372f
C1130 VTAIL.t12 VSUBS 0.252073f
C1131 VTAIL.t13 VSUBS 0.252073f
C1132 VTAIL.n142 VSUBS 1.82794f
C1133 VTAIL.n143 VSUBS 1.0489f
C1134 VTAIL.n144 VSUBS 0.0266f
C1135 VTAIL.n145 VSUBS 0.025077f
C1136 VTAIL.n146 VSUBS 0.013476f
C1137 VTAIL.n147 VSUBS 0.031851f
C1138 VTAIL.n148 VSUBS 0.014268f
C1139 VTAIL.n149 VSUBS 0.025077f
C1140 VTAIL.n150 VSUBS 0.013476f
C1141 VTAIL.n151 VSUBS 0.031851f
C1142 VTAIL.n152 VSUBS 0.014268f
C1143 VTAIL.n153 VSUBS 0.025077f
C1144 VTAIL.n154 VSUBS 0.013476f
C1145 VTAIL.n155 VSUBS 0.031851f
C1146 VTAIL.n156 VSUBS 0.014268f
C1147 VTAIL.n157 VSUBS 0.025077f
C1148 VTAIL.n158 VSUBS 0.013476f
C1149 VTAIL.n159 VSUBS 0.031851f
C1150 VTAIL.n160 VSUBS 0.014268f
C1151 VTAIL.n161 VSUBS 0.025077f
C1152 VTAIL.n162 VSUBS 0.013476f
C1153 VTAIL.n163 VSUBS 0.031851f
C1154 VTAIL.n164 VSUBS 0.014268f
C1155 VTAIL.n165 VSUBS 0.205662f
C1156 VTAIL.t8 VSUBS 0.068695f
C1157 VTAIL.n166 VSUBS 0.023889f
C1158 VTAIL.n167 VSUBS 0.02396f
C1159 VTAIL.n168 VSUBS 0.013476f
C1160 VTAIL.n169 VSUBS 1.31126f
C1161 VTAIL.n170 VSUBS 0.025077f
C1162 VTAIL.n171 VSUBS 0.013476f
C1163 VTAIL.n172 VSUBS 0.014268f
C1164 VTAIL.n173 VSUBS 0.031851f
C1165 VTAIL.n174 VSUBS 0.031851f
C1166 VTAIL.n175 VSUBS 0.014268f
C1167 VTAIL.n176 VSUBS 0.013476f
C1168 VTAIL.n177 VSUBS 0.025077f
C1169 VTAIL.n178 VSUBS 0.025077f
C1170 VTAIL.n179 VSUBS 0.013476f
C1171 VTAIL.n180 VSUBS 0.014268f
C1172 VTAIL.n181 VSUBS 0.031851f
C1173 VTAIL.n182 VSUBS 0.031851f
C1174 VTAIL.n183 VSUBS 0.031851f
C1175 VTAIL.n184 VSUBS 0.014268f
C1176 VTAIL.n185 VSUBS 0.013476f
C1177 VTAIL.n186 VSUBS 0.025077f
C1178 VTAIL.n187 VSUBS 0.025077f
C1179 VTAIL.n188 VSUBS 0.013476f
C1180 VTAIL.n189 VSUBS 0.013872f
C1181 VTAIL.n190 VSUBS 0.013872f
C1182 VTAIL.n191 VSUBS 0.031851f
C1183 VTAIL.n192 VSUBS 0.031851f
C1184 VTAIL.n193 VSUBS 0.014268f
C1185 VTAIL.n194 VSUBS 0.013476f
C1186 VTAIL.n195 VSUBS 0.025077f
C1187 VTAIL.n196 VSUBS 0.025077f
C1188 VTAIL.n197 VSUBS 0.013476f
C1189 VTAIL.n198 VSUBS 0.014268f
C1190 VTAIL.n199 VSUBS 0.031851f
C1191 VTAIL.n200 VSUBS 0.031851f
C1192 VTAIL.n201 VSUBS 0.014268f
C1193 VTAIL.n202 VSUBS 0.013476f
C1194 VTAIL.n203 VSUBS 0.025077f
C1195 VTAIL.n204 VSUBS 0.025077f
C1196 VTAIL.n205 VSUBS 0.013476f
C1197 VTAIL.n206 VSUBS 0.014268f
C1198 VTAIL.n207 VSUBS 0.031851f
C1199 VTAIL.n208 VSUBS 0.073855f
C1200 VTAIL.n209 VSUBS 0.014268f
C1201 VTAIL.n210 VSUBS 0.013476f
C1202 VTAIL.n211 VSUBS 0.053854f
C1203 VTAIL.n212 VSUBS 0.036866f
C1204 VTAIL.n213 VSUBS 1.69443f
C1205 VTAIL.n214 VSUBS 0.0266f
C1206 VTAIL.n215 VSUBS 0.025077f
C1207 VTAIL.n216 VSUBS 0.013476f
C1208 VTAIL.n217 VSUBS 0.031851f
C1209 VTAIL.n218 VSUBS 0.014268f
C1210 VTAIL.n219 VSUBS 0.025077f
C1211 VTAIL.n220 VSUBS 0.013476f
C1212 VTAIL.n221 VSUBS 0.031851f
C1213 VTAIL.n222 VSUBS 0.014268f
C1214 VTAIL.n223 VSUBS 0.025077f
C1215 VTAIL.n224 VSUBS 0.013476f
C1216 VTAIL.n225 VSUBS 0.031851f
C1217 VTAIL.n226 VSUBS 0.014268f
C1218 VTAIL.n227 VSUBS 0.025077f
C1219 VTAIL.n228 VSUBS 0.013476f
C1220 VTAIL.n229 VSUBS 0.031851f
C1221 VTAIL.n230 VSUBS 0.031851f
C1222 VTAIL.n231 VSUBS 0.014268f
C1223 VTAIL.n232 VSUBS 0.025077f
C1224 VTAIL.n233 VSUBS 0.013476f
C1225 VTAIL.n234 VSUBS 0.031851f
C1226 VTAIL.n235 VSUBS 0.014268f
C1227 VTAIL.n236 VSUBS 0.205662f
C1228 VTAIL.t3 VSUBS 0.068695f
C1229 VTAIL.n237 VSUBS 0.023889f
C1230 VTAIL.n238 VSUBS 0.02396f
C1231 VTAIL.n239 VSUBS 0.013476f
C1232 VTAIL.n240 VSUBS 1.31126f
C1233 VTAIL.n241 VSUBS 0.025077f
C1234 VTAIL.n242 VSUBS 0.013476f
C1235 VTAIL.n243 VSUBS 0.014268f
C1236 VTAIL.n244 VSUBS 0.031851f
C1237 VTAIL.n245 VSUBS 0.031851f
C1238 VTAIL.n246 VSUBS 0.014268f
C1239 VTAIL.n247 VSUBS 0.013476f
C1240 VTAIL.n248 VSUBS 0.025077f
C1241 VTAIL.n249 VSUBS 0.025077f
C1242 VTAIL.n250 VSUBS 0.013476f
C1243 VTAIL.n251 VSUBS 0.014268f
C1244 VTAIL.n252 VSUBS 0.031851f
C1245 VTAIL.n253 VSUBS 0.031851f
C1246 VTAIL.n254 VSUBS 0.014268f
C1247 VTAIL.n255 VSUBS 0.013476f
C1248 VTAIL.n256 VSUBS 0.025077f
C1249 VTAIL.n257 VSUBS 0.025077f
C1250 VTAIL.n258 VSUBS 0.013476f
C1251 VTAIL.n259 VSUBS 0.013872f
C1252 VTAIL.n260 VSUBS 0.013872f
C1253 VTAIL.n261 VSUBS 0.031851f
C1254 VTAIL.n262 VSUBS 0.031851f
C1255 VTAIL.n263 VSUBS 0.014268f
C1256 VTAIL.n264 VSUBS 0.013476f
C1257 VTAIL.n265 VSUBS 0.025077f
C1258 VTAIL.n266 VSUBS 0.025077f
C1259 VTAIL.n267 VSUBS 0.013476f
C1260 VTAIL.n268 VSUBS 0.014268f
C1261 VTAIL.n269 VSUBS 0.031851f
C1262 VTAIL.n270 VSUBS 0.031851f
C1263 VTAIL.n271 VSUBS 0.014268f
C1264 VTAIL.n272 VSUBS 0.013476f
C1265 VTAIL.n273 VSUBS 0.025077f
C1266 VTAIL.n274 VSUBS 0.025077f
C1267 VTAIL.n275 VSUBS 0.013476f
C1268 VTAIL.n276 VSUBS 0.014268f
C1269 VTAIL.n277 VSUBS 0.031851f
C1270 VTAIL.n278 VSUBS 0.073855f
C1271 VTAIL.n279 VSUBS 0.014268f
C1272 VTAIL.n280 VSUBS 0.013476f
C1273 VTAIL.n281 VSUBS 0.053854f
C1274 VTAIL.n282 VSUBS 0.036866f
C1275 VTAIL.n283 VSUBS 1.69443f
C1276 VTAIL.t4 VSUBS 0.252073f
C1277 VTAIL.t6 VSUBS 0.252073f
C1278 VTAIL.n284 VSUBS 1.82795f
C1279 VTAIL.n285 VSUBS 1.04889f
C1280 VTAIL.n286 VSUBS 0.0266f
C1281 VTAIL.n287 VSUBS 0.025077f
C1282 VTAIL.n288 VSUBS 0.013476f
C1283 VTAIL.n289 VSUBS 0.031851f
C1284 VTAIL.n290 VSUBS 0.014268f
C1285 VTAIL.n291 VSUBS 0.025077f
C1286 VTAIL.n292 VSUBS 0.013476f
C1287 VTAIL.n293 VSUBS 0.031851f
C1288 VTAIL.n294 VSUBS 0.014268f
C1289 VTAIL.n295 VSUBS 0.025077f
C1290 VTAIL.n296 VSUBS 0.013476f
C1291 VTAIL.n297 VSUBS 0.031851f
C1292 VTAIL.n298 VSUBS 0.014268f
C1293 VTAIL.n299 VSUBS 0.025077f
C1294 VTAIL.n300 VSUBS 0.013476f
C1295 VTAIL.n301 VSUBS 0.031851f
C1296 VTAIL.n302 VSUBS 0.031851f
C1297 VTAIL.n303 VSUBS 0.014268f
C1298 VTAIL.n304 VSUBS 0.025077f
C1299 VTAIL.n305 VSUBS 0.013476f
C1300 VTAIL.n306 VSUBS 0.031851f
C1301 VTAIL.n307 VSUBS 0.014268f
C1302 VTAIL.n308 VSUBS 0.205662f
C1303 VTAIL.t2 VSUBS 0.068695f
C1304 VTAIL.n309 VSUBS 0.023889f
C1305 VTAIL.n310 VSUBS 0.02396f
C1306 VTAIL.n311 VSUBS 0.013476f
C1307 VTAIL.n312 VSUBS 1.31126f
C1308 VTAIL.n313 VSUBS 0.025077f
C1309 VTAIL.n314 VSUBS 0.013476f
C1310 VTAIL.n315 VSUBS 0.014268f
C1311 VTAIL.n316 VSUBS 0.031851f
C1312 VTAIL.n317 VSUBS 0.031851f
C1313 VTAIL.n318 VSUBS 0.014268f
C1314 VTAIL.n319 VSUBS 0.013476f
C1315 VTAIL.n320 VSUBS 0.025077f
C1316 VTAIL.n321 VSUBS 0.025077f
C1317 VTAIL.n322 VSUBS 0.013476f
C1318 VTAIL.n323 VSUBS 0.014268f
C1319 VTAIL.n324 VSUBS 0.031851f
C1320 VTAIL.n325 VSUBS 0.031851f
C1321 VTAIL.n326 VSUBS 0.014268f
C1322 VTAIL.n327 VSUBS 0.013476f
C1323 VTAIL.n328 VSUBS 0.025077f
C1324 VTAIL.n329 VSUBS 0.025077f
C1325 VTAIL.n330 VSUBS 0.013476f
C1326 VTAIL.n331 VSUBS 0.013872f
C1327 VTAIL.n332 VSUBS 0.013872f
C1328 VTAIL.n333 VSUBS 0.031851f
C1329 VTAIL.n334 VSUBS 0.031851f
C1330 VTAIL.n335 VSUBS 0.014268f
C1331 VTAIL.n336 VSUBS 0.013476f
C1332 VTAIL.n337 VSUBS 0.025077f
C1333 VTAIL.n338 VSUBS 0.025077f
C1334 VTAIL.n339 VSUBS 0.013476f
C1335 VTAIL.n340 VSUBS 0.014268f
C1336 VTAIL.n341 VSUBS 0.031851f
C1337 VTAIL.n342 VSUBS 0.031851f
C1338 VTAIL.n343 VSUBS 0.014268f
C1339 VTAIL.n344 VSUBS 0.013476f
C1340 VTAIL.n345 VSUBS 0.025077f
C1341 VTAIL.n346 VSUBS 0.025077f
C1342 VTAIL.n347 VSUBS 0.013476f
C1343 VTAIL.n348 VSUBS 0.014268f
C1344 VTAIL.n349 VSUBS 0.031851f
C1345 VTAIL.n350 VSUBS 0.073855f
C1346 VTAIL.n351 VSUBS 0.014268f
C1347 VTAIL.n352 VSUBS 0.013476f
C1348 VTAIL.n353 VSUBS 0.053854f
C1349 VTAIL.n354 VSUBS 0.036866f
C1350 VTAIL.n355 VSUBS 0.281372f
C1351 VTAIL.n356 VSUBS 0.0266f
C1352 VTAIL.n357 VSUBS 0.025077f
C1353 VTAIL.n358 VSUBS 0.013476f
C1354 VTAIL.n359 VSUBS 0.031851f
C1355 VTAIL.n360 VSUBS 0.014268f
C1356 VTAIL.n361 VSUBS 0.025077f
C1357 VTAIL.n362 VSUBS 0.013476f
C1358 VTAIL.n363 VSUBS 0.031851f
C1359 VTAIL.n364 VSUBS 0.014268f
C1360 VTAIL.n365 VSUBS 0.025077f
C1361 VTAIL.n366 VSUBS 0.013476f
C1362 VTAIL.n367 VSUBS 0.031851f
C1363 VTAIL.n368 VSUBS 0.014268f
C1364 VTAIL.n369 VSUBS 0.025077f
C1365 VTAIL.n370 VSUBS 0.013476f
C1366 VTAIL.n371 VSUBS 0.031851f
C1367 VTAIL.n372 VSUBS 0.031851f
C1368 VTAIL.n373 VSUBS 0.014268f
C1369 VTAIL.n374 VSUBS 0.025077f
C1370 VTAIL.n375 VSUBS 0.013476f
C1371 VTAIL.n376 VSUBS 0.031851f
C1372 VTAIL.n377 VSUBS 0.014268f
C1373 VTAIL.n378 VSUBS 0.205662f
C1374 VTAIL.t9 VSUBS 0.068695f
C1375 VTAIL.n379 VSUBS 0.023889f
C1376 VTAIL.n380 VSUBS 0.02396f
C1377 VTAIL.n381 VSUBS 0.013476f
C1378 VTAIL.n382 VSUBS 1.31126f
C1379 VTAIL.n383 VSUBS 0.025077f
C1380 VTAIL.n384 VSUBS 0.013476f
C1381 VTAIL.n385 VSUBS 0.014268f
C1382 VTAIL.n386 VSUBS 0.031851f
C1383 VTAIL.n387 VSUBS 0.031851f
C1384 VTAIL.n388 VSUBS 0.014268f
C1385 VTAIL.n389 VSUBS 0.013476f
C1386 VTAIL.n390 VSUBS 0.025077f
C1387 VTAIL.n391 VSUBS 0.025077f
C1388 VTAIL.n392 VSUBS 0.013476f
C1389 VTAIL.n393 VSUBS 0.014268f
C1390 VTAIL.n394 VSUBS 0.031851f
C1391 VTAIL.n395 VSUBS 0.031851f
C1392 VTAIL.n396 VSUBS 0.014268f
C1393 VTAIL.n397 VSUBS 0.013476f
C1394 VTAIL.n398 VSUBS 0.025077f
C1395 VTAIL.n399 VSUBS 0.025077f
C1396 VTAIL.n400 VSUBS 0.013476f
C1397 VTAIL.n401 VSUBS 0.013872f
C1398 VTAIL.n402 VSUBS 0.013872f
C1399 VTAIL.n403 VSUBS 0.031851f
C1400 VTAIL.n404 VSUBS 0.031851f
C1401 VTAIL.n405 VSUBS 0.014268f
C1402 VTAIL.n406 VSUBS 0.013476f
C1403 VTAIL.n407 VSUBS 0.025077f
C1404 VTAIL.n408 VSUBS 0.025077f
C1405 VTAIL.n409 VSUBS 0.013476f
C1406 VTAIL.n410 VSUBS 0.014268f
C1407 VTAIL.n411 VSUBS 0.031851f
C1408 VTAIL.n412 VSUBS 0.031851f
C1409 VTAIL.n413 VSUBS 0.014268f
C1410 VTAIL.n414 VSUBS 0.013476f
C1411 VTAIL.n415 VSUBS 0.025077f
C1412 VTAIL.n416 VSUBS 0.025077f
C1413 VTAIL.n417 VSUBS 0.013476f
C1414 VTAIL.n418 VSUBS 0.014268f
C1415 VTAIL.n419 VSUBS 0.031851f
C1416 VTAIL.n420 VSUBS 0.073855f
C1417 VTAIL.n421 VSUBS 0.014268f
C1418 VTAIL.n422 VSUBS 0.013476f
C1419 VTAIL.n423 VSUBS 0.053854f
C1420 VTAIL.n424 VSUBS 0.036866f
C1421 VTAIL.n425 VSUBS 0.281372f
C1422 VTAIL.t14 VSUBS 0.252073f
C1423 VTAIL.t15 VSUBS 0.252073f
C1424 VTAIL.n426 VSUBS 1.82795f
C1425 VTAIL.n427 VSUBS 1.04889f
C1426 VTAIL.n428 VSUBS 0.0266f
C1427 VTAIL.n429 VSUBS 0.025077f
C1428 VTAIL.n430 VSUBS 0.013476f
C1429 VTAIL.n431 VSUBS 0.031851f
C1430 VTAIL.n432 VSUBS 0.014268f
C1431 VTAIL.n433 VSUBS 0.025077f
C1432 VTAIL.n434 VSUBS 0.013476f
C1433 VTAIL.n435 VSUBS 0.031851f
C1434 VTAIL.n436 VSUBS 0.014268f
C1435 VTAIL.n437 VSUBS 0.025077f
C1436 VTAIL.n438 VSUBS 0.013476f
C1437 VTAIL.n439 VSUBS 0.031851f
C1438 VTAIL.n440 VSUBS 0.014268f
C1439 VTAIL.n441 VSUBS 0.025077f
C1440 VTAIL.n442 VSUBS 0.013476f
C1441 VTAIL.n443 VSUBS 0.031851f
C1442 VTAIL.n444 VSUBS 0.031851f
C1443 VTAIL.n445 VSUBS 0.014268f
C1444 VTAIL.n446 VSUBS 0.025077f
C1445 VTAIL.n447 VSUBS 0.013476f
C1446 VTAIL.n448 VSUBS 0.031851f
C1447 VTAIL.n449 VSUBS 0.014268f
C1448 VTAIL.n450 VSUBS 0.205662f
C1449 VTAIL.t11 VSUBS 0.068695f
C1450 VTAIL.n451 VSUBS 0.023889f
C1451 VTAIL.n452 VSUBS 0.02396f
C1452 VTAIL.n453 VSUBS 0.013476f
C1453 VTAIL.n454 VSUBS 1.31126f
C1454 VTAIL.n455 VSUBS 0.025077f
C1455 VTAIL.n456 VSUBS 0.013476f
C1456 VTAIL.n457 VSUBS 0.014268f
C1457 VTAIL.n458 VSUBS 0.031851f
C1458 VTAIL.n459 VSUBS 0.031851f
C1459 VTAIL.n460 VSUBS 0.014268f
C1460 VTAIL.n461 VSUBS 0.013476f
C1461 VTAIL.n462 VSUBS 0.025077f
C1462 VTAIL.n463 VSUBS 0.025077f
C1463 VTAIL.n464 VSUBS 0.013476f
C1464 VTAIL.n465 VSUBS 0.014268f
C1465 VTAIL.n466 VSUBS 0.031851f
C1466 VTAIL.n467 VSUBS 0.031851f
C1467 VTAIL.n468 VSUBS 0.014268f
C1468 VTAIL.n469 VSUBS 0.013476f
C1469 VTAIL.n470 VSUBS 0.025077f
C1470 VTAIL.n471 VSUBS 0.025077f
C1471 VTAIL.n472 VSUBS 0.013476f
C1472 VTAIL.n473 VSUBS 0.013872f
C1473 VTAIL.n474 VSUBS 0.013872f
C1474 VTAIL.n475 VSUBS 0.031851f
C1475 VTAIL.n476 VSUBS 0.031851f
C1476 VTAIL.n477 VSUBS 0.014268f
C1477 VTAIL.n478 VSUBS 0.013476f
C1478 VTAIL.n479 VSUBS 0.025077f
C1479 VTAIL.n480 VSUBS 0.025077f
C1480 VTAIL.n481 VSUBS 0.013476f
C1481 VTAIL.n482 VSUBS 0.014268f
C1482 VTAIL.n483 VSUBS 0.031851f
C1483 VTAIL.n484 VSUBS 0.031851f
C1484 VTAIL.n485 VSUBS 0.014268f
C1485 VTAIL.n486 VSUBS 0.013476f
C1486 VTAIL.n487 VSUBS 0.025077f
C1487 VTAIL.n488 VSUBS 0.025077f
C1488 VTAIL.n489 VSUBS 0.013476f
C1489 VTAIL.n490 VSUBS 0.014268f
C1490 VTAIL.n491 VSUBS 0.031851f
C1491 VTAIL.n492 VSUBS 0.073855f
C1492 VTAIL.n493 VSUBS 0.014268f
C1493 VTAIL.n494 VSUBS 0.013476f
C1494 VTAIL.n495 VSUBS 0.053854f
C1495 VTAIL.n496 VSUBS 0.036866f
C1496 VTAIL.n497 VSUBS 1.69443f
C1497 VTAIL.n498 VSUBS 0.0266f
C1498 VTAIL.n499 VSUBS 0.025077f
C1499 VTAIL.n500 VSUBS 0.013476f
C1500 VTAIL.n501 VSUBS 0.031851f
C1501 VTAIL.n502 VSUBS 0.014268f
C1502 VTAIL.n503 VSUBS 0.025077f
C1503 VTAIL.n504 VSUBS 0.013476f
C1504 VTAIL.n505 VSUBS 0.031851f
C1505 VTAIL.n506 VSUBS 0.014268f
C1506 VTAIL.n507 VSUBS 0.025077f
C1507 VTAIL.n508 VSUBS 0.013476f
C1508 VTAIL.n509 VSUBS 0.031851f
C1509 VTAIL.n510 VSUBS 0.014268f
C1510 VTAIL.n511 VSUBS 0.025077f
C1511 VTAIL.n512 VSUBS 0.013476f
C1512 VTAIL.n513 VSUBS 0.031851f
C1513 VTAIL.n514 VSUBS 0.014268f
C1514 VTAIL.n515 VSUBS 0.025077f
C1515 VTAIL.n516 VSUBS 0.013476f
C1516 VTAIL.n517 VSUBS 0.031851f
C1517 VTAIL.n518 VSUBS 0.014268f
C1518 VTAIL.n519 VSUBS 0.205662f
C1519 VTAIL.t1 VSUBS 0.068695f
C1520 VTAIL.n520 VSUBS 0.023889f
C1521 VTAIL.n521 VSUBS 0.02396f
C1522 VTAIL.n522 VSUBS 0.013476f
C1523 VTAIL.n523 VSUBS 1.31126f
C1524 VTAIL.n524 VSUBS 0.025077f
C1525 VTAIL.n525 VSUBS 0.013476f
C1526 VTAIL.n526 VSUBS 0.014268f
C1527 VTAIL.n527 VSUBS 0.031851f
C1528 VTAIL.n528 VSUBS 0.031851f
C1529 VTAIL.n529 VSUBS 0.014268f
C1530 VTAIL.n530 VSUBS 0.013476f
C1531 VTAIL.n531 VSUBS 0.025077f
C1532 VTAIL.n532 VSUBS 0.025077f
C1533 VTAIL.n533 VSUBS 0.013476f
C1534 VTAIL.n534 VSUBS 0.014268f
C1535 VTAIL.n535 VSUBS 0.031851f
C1536 VTAIL.n536 VSUBS 0.031851f
C1537 VTAIL.n537 VSUBS 0.031851f
C1538 VTAIL.n538 VSUBS 0.014268f
C1539 VTAIL.n539 VSUBS 0.013476f
C1540 VTAIL.n540 VSUBS 0.025077f
C1541 VTAIL.n541 VSUBS 0.025077f
C1542 VTAIL.n542 VSUBS 0.013476f
C1543 VTAIL.n543 VSUBS 0.013872f
C1544 VTAIL.n544 VSUBS 0.013872f
C1545 VTAIL.n545 VSUBS 0.031851f
C1546 VTAIL.n546 VSUBS 0.031851f
C1547 VTAIL.n547 VSUBS 0.014268f
C1548 VTAIL.n548 VSUBS 0.013476f
C1549 VTAIL.n549 VSUBS 0.025077f
C1550 VTAIL.n550 VSUBS 0.025077f
C1551 VTAIL.n551 VSUBS 0.013476f
C1552 VTAIL.n552 VSUBS 0.014268f
C1553 VTAIL.n553 VSUBS 0.031851f
C1554 VTAIL.n554 VSUBS 0.031851f
C1555 VTAIL.n555 VSUBS 0.014268f
C1556 VTAIL.n556 VSUBS 0.013476f
C1557 VTAIL.n557 VSUBS 0.025077f
C1558 VTAIL.n558 VSUBS 0.025077f
C1559 VTAIL.n559 VSUBS 0.013476f
C1560 VTAIL.n560 VSUBS 0.014268f
C1561 VTAIL.n561 VSUBS 0.031851f
C1562 VTAIL.n562 VSUBS 0.073855f
C1563 VTAIL.n563 VSUBS 0.014268f
C1564 VTAIL.n564 VSUBS 0.013476f
C1565 VTAIL.n565 VSUBS 0.053854f
C1566 VTAIL.n566 VSUBS 0.036866f
C1567 VTAIL.n567 VSUBS 1.68973f
C1568 VP.n0 VSUBS 0.038833f
C1569 VP.t5 VSUBS 2.95472f
C1570 VP.n1 VSUBS 0.059561f
C1571 VP.n2 VSUBS 0.029453f
C1572 VP.n3 VSUBS 0.035556f
C1573 VP.n4 VSUBS 0.029453f
C1574 VP.n5 VSUBS 0.043182f
C1575 VP.n6 VSUBS 0.029453f
C1576 VP.t0 VSUBS 2.95472f
C1577 VP.n7 VSUBS 0.055167f
C1578 VP.n8 VSUBS 0.029453f
C1579 VP.n9 VSUBS 0.055167f
C1580 VP.n10 VSUBS 0.038833f
C1581 VP.t2 VSUBS 2.95472f
C1582 VP.n11 VSUBS 0.059561f
C1583 VP.n12 VSUBS 0.029453f
C1584 VP.n13 VSUBS 0.035556f
C1585 VP.n14 VSUBS 0.029453f
C1586 VP.n15 VSUBS 0.043182f
C1587 VP.n16 VSUBS 0.312172f
C1588 VP.t4 VSUBS 2.95472f
C1589 VP.t6 VSUBS 3.25215f
C1590 VP.n17 VSUBS 1.09077f
C1591 VP.n18 VSUBS 1.13708f
C1592 VP.n19 VSUBS 0.047541f
C1593 VP.n20 VSUBS 0.055167f
C1594 VP.n21 VSUBS 0.029453f
C1595 VP.n22 VSUBS 0.029453f
C1596 VP.n23 VSUBS 0.029453f
C1597 VP.n24 VSUBS 0.043182f
C1598 VP.n25 VSUBS 0.055167f
C1599 VP.t3 VSUBS 2.95472f
C1600 VP.n26 VSUBS 1.03865f
C1601 VP.n27 VSUBS 0.047541f
C1602 VP.n28 VSUBS 0.029453f
C1603 VP.n29 VSUBS 0.029453f
C1604 VP.n30 VSUBS 0.029453f
C1605 VP.n31 VSUBS 0.055167f
C1606 VP.n32 VSUBS 0.057793f
C1607 VP.n33 VSUBS 0.024178f
C1608 VP.n34 VSUBS 0.029453f
C1609 VP.n35 VSUBS 0.029453f
C1610 VP.n36 VSUBS 0.029453f
C1611 VP.n37 VSUBS 0.055167f
C1612 VP.n38 VSUBS 0.032287f
C1613 VP.n39 VSUBS 1.13951f
C1614 VP.n40 VSUBS 1.78121f
C1615 VP.n41 VSUBS 1.8012f
C1616 VP.t1 VSUBS 2.95472f
C1617 VP.n42 VSUBS 1.13951f
C1618 VP.n43 VSUBS 0.032287f
C1619 VP.n44 VSUBS 0.038833f
C1620 VP.n45 VSUBS 0.029453f
C1621 VP.n46 VSUBS 0.029453f
C1622 VP.n47 VSUBS 0.059561f
C1623 VP.n48 VSUBS 0.024178f
C1624 VP.n49 VSUBS 0.057793f
C1625 VP.n50 VSUBS 0.029453f
C1626 VP.n51 VSUBS 0.029453f
C1627 VP.n52 VSUBS 0.029453f
C1628 VP.n53 VSUBS 0.035556f
C1629 VP.n54 VSUBS 1.03865f
C1630 VP.n55 VSUBS 0.047541f
C1631 VP.n56 VSUBS 0.055167f
C1632 VP.n57 VSUBS 0.029453f
C1633 VP.n58 VSUBS 0.029453f
C1634 VP.n59 VSUBS 0.029453f
C1635 VP.n60 VSUBS 0.043182f
C1636 VP.n61 VSUBS 0.055167f
C1637 VP.t7 VSUBS 2.95472f
C1638 VP.n62 VSUBS 1.03865f
C1639 VP.n63 VSUBS 0.047541f
C1640 VP.n64 VSUBS 0.029453f
C1641 VP.n65 VSUBS 0.029453f
C1642 VP.n66 VSUBS 0.029453f
C1643 VP.n67 VSUBS 0.055167f
C1644 VP.n68 VSUBS 0.057793f
C1645 VP.n69 VSUBS 0.024178f
C1646 VP.n70 VSUBS 0.029453f
C1647 VP.n71 VSUBS 0.029453f
C1648 VP.n72 VSUBS 0.029453f
C1649 VP.n73 VSUBS 0.055167f
C1650 VP.n74 VSUBS 0.032287f
C1651 VP.n75 VSUBS 1.13951f
C1652 VP.n76 VSUBS 0.055348f
.ends

