* NGSPICE file created from diff_pair_sample_0169.ext - technology: sky130A

.subckt diff_pair_sample_0169 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 w_n4322_n1230# sky130_fd_pr__pfet_01v8 ad=0.5109 pd=3.4 as=0.21615 ps=1.64 w=1.31 l=3.86
X1 VDD1.t4 VP.t1 VTAIL.t7 w_n4322_n1230# sky130_fd_pr__pfet_01v8 ad=0.5109 pd=3.4 as=0.21615 ps=1.64 w=1.31 l=3.86
X2 VTAIL.t6 VP.t2 VDD1.t3 w_n4322_n1230# sky130_fd_pr__pfet_01v8 ad=0.21615 pd=1.64 as=0.21615 ps=1.64 w=1.31 l=3.86
X3 VDD1.t2 VP.t3 VTAIL.t9 w_n4322_n1230# sky130_fd_pr__pfet_01v8 ad=0.21615 pd=1.64 as=0.5109 ps=3.4 w=1.31 l=3.86
X4 VDD2.t5 VN.t0 VTAIL.t5 w_n4322_n1230# sky130_fd_pr__pfet_01v8 ad=0.5109 pd=3.4 as=0.21615 ps=1.64 w=1.31 l=3.86
X5 B.t11 B.t9 B.t10 w_n4322_n1230# sky130_fd_pr__pfet_01v8 ad=0.5109 pd=3.4 as=0 ps=0 w=1.31 l=3.86
X6 B.t8 B.t6 B.t7 w_n4322_n1230# sky130_fd_pr__pfet_01v8 ad=0.5109 pd=3.4 as=0 ps=0 w=1.31 l=3.86
X7 VTAIL.t10 VP.t4 VDD1.t1 w_n4322_n1230# sky130_fd_pr__pfet_01v8 ad=0.21615 pd=1.64 as=0.21615 ps=1.64 w=1.31 l=3.86
X8 VDD2.t4 VN.t1 VTAIL.t1 w_n4322_n1230# sky130_fd_pr__pfet_01v8 ad=0.21615 pd=1.64 as=0.5109 ps=3.4 w=1.31 l=3.86
X9 VDD2.t3 VN.t2 VTAIL.t4 w_n4322_n1230# sky130_fd_pr__pfet_01v8 ad=0.21615 pd=1.64 as=0.5109 ps=3.4 w=1.31 l=3.86
X10 VDD2.t2 VN.t3 VTAIL.t3 w_n4322_n1230# sky130_fd_pr__pfet_01v8 ad=0.5109 pd=3.4 as=0.21615 ps=1.64 w=1.31 l=3.86
X11 VTAIL.t0 VN.t4 VDD2.t1 w_n4322_n1230# sky130_fd_pr__pfet_01v8 ad=0.21615 pd=1.64 as=0.21615 ps=1.64 w=1.31 l=3.86
X12 B.t5 B.t3 B.t4 w_n4322_n1230# sky130_fd_pr__pfet_01v8 ad=0.5109 pd=3.4 as=0 ps=0 w=1.31 l=3.86
X13 VDD1.t0 VP.t5 VTAIL.t11 w_n4322_n1230# sky130_fd_pr__pfet_01v8 ad=0.21615 pd=1.64 as=0.5109 ps=3.4 w=1.31 l=3.86
X14 B.t2 B.t0 B.t1 w_n4322_n1230# sky130_fd_pr__pfet_01v8 ad=0.5109 pd=3.4 as=0 ps=0 w=1.31 l=3.86
X15 VTAIL.t2 VN.t5 VDD2.t0 w_n4322_n1230# sky130_fd_pr__pfet_01v8 ad=0.21615 pd=1.64 as=0.21615 ps=1.64 w=1.31 l=3.86
R0 VP.n15 VP.n14 161.3
R1 VP.n16 VP.n11 161.3
R2 VP.n18 VP.n17 161.3
R3 VP.n19 VP.n10 161.3
R4 VP.n21 VP.n20 161.3
R5 VP.n22 VP.n9 161.3
R6 VP.n24 VP.n23 161.3
R7 VP.n25 VP.n8 161.3
R8 VP.n54 VP.n0 161.3
R9 VP.n53 VP.n52 161.3
R10 VP.n51 VP.n1 161.3
R11 VP.n50 VP.n49 161.3
R12 VP.n48 VP.n2 161.3
R13 VP.n47 VP.n46 161.3
R14 VP.n45 VP.n3 161.3
R15 VP.n44 VP.n43 161.3
R16 VP.n41 VP.n4 161.3
R17 VP.n40 VP.n39 161.3
R18 VP.n38 VP.n5 161.3
R19 VP.n37 VP.n36 161.3
R20 VP.n35 VP.n6 161.3
R21 VP.n34 VP.n33 161.3
R22 VP.n32 VP.n7 161.3
R23 VP.n31 VP.n30 161.3
R24 VP.n13 VP.n12 62.8644
R25 VP.n29 VP.n28 60.6508
R26 VP.n56 VP.n55 60.6508
R27 VP.n27 VP.n26 60.6508
R28 VP.n36 VP.n35 55.548
R29 VP.n49 VP.n48 55.548
R30 VP.n20 VP.n19 55.548
R31 VP.n28 VP.n27 45.7502
R32 VP.n12 VP.t0 40.3864
R33 VP.n35 VP.n34 25.4388
R34 VP.n49 VP.n1 25.4388
R35 VP.n20 VP.n9 25.4388
R36 VP.n30 VP.n7 24.4675
R37 VP.n34 VP.n7 24.4675
R38 VP.n36 VP.n5 24.4675
R39 VP.n40 VP.n5 24.4675
R40 VP.n41 VP.n40 24.4675
R41 VP.n43 VP.n3 24.4675
R42 VP.n47 VP.n3 24.4675
R43 VP.n48 VP.n47 24.4675
R44 VP.n53 VP.n1 24.4675
R45 VP.n54 VP.n53 24.4675
R46 VP.n24 VP.n9 24.4675
R47 VP.n25 VP.n24 24.4675
R48 VP.n14 VP.n11 24.4675
R49 VP.n18 VP.n11 24.4675
R50 VP.n19 VP.n18 24.4675
R51 VP.n30 VP.n29 21.5315
R52 VP.n55 VP.n54 21.5315
R53 VP.n26 VP.n25 21.5315
R54 VP.n42 VP.n41 12.234
R55 VP.n43 VP.n42 12.234
R56 VP.n14 VP.n13 12.234
R57 VP.n29 VP.t1 8.17952
R58 VP.n42 VP.t4 8.17952
R59 VP.n55 VP.t5 8.17952
R60 VP.n26 VP.t3 8.17952
R61 VP.n13 VP.t2 8.17952
R62 VP.n15 VP.n12 2.6395
R63 VP.n27 VP.n8 0.417535
R64 VP.n31 VP.n28 0.417535
R65 VP.n56 VP.n0 0.417535
R66 VP VP.n56 0.394291
R67 VP.n16 VP.n15 0.189894
R68 VP.n17 VP.n16 0.189894
R69 VP.n17 VP.n10 0.189894
R70 VP.n21 VP.n10 0.189894
R71 VP.n22 VP.n21 0.189894
R72 VP.n23 VP.n22 0.189894
R73 VP.n23 VP.n8 0.189894
R74 VP.n32 VP.n31 0.189894
R75 VP.n33 VP.n32 0.189894
R76 VP.n33 VP.n6 0.189894
R77 VP.n37 VP.n6 0.189894
R78 VP.n38 VP.n37 0.189894
R79 VP.n39 VP.n38 0.189894
R80 VP.n39 VP.n4 0.189894
R81 VP.n44 VP.n4 0.189894
R82 VP.n45 VP.n44 0.189894
R83 VP.n46 VP.n45 0.189894
R84 VP.n46 VP.n2 0.189894
R85 VP.n50 VP.n2 0.189894
R86 VP.n51 VP.n50 0.189894
R87 VP.n52 VP.n51 0.189894
R88 VP.n52 VP.n0 0.189894
R89 VTAIL.n7 VTAIL.t1 373.281
R90 VTAIL.n11 VTAIL.t4 373.281
R91 VTAIL.n2 VTAIL.t11 373.281
R92 VTAIL.n10 VTAIL.t9 373.281
R93 VTAIL.n1 VTAIL.n0 330.344
R94 VTAIL.n4 VTAIL.n3 330.344
R95 VTAIL.n9 VTAIL.n8 330.344
R96 VTAIL.n6 VTAIL.n5 330.344
R97 VTAIL.n0 VTAIL.t3 24.8135
R98 VTAIL.n0 VTAIL.t2 24.8135
R99 VTAIL.n3 VTAIL.t7 24.8135
R100 VTAIL.n3 VTAIL.t10 24.8135
R101 VTAIL.n8 VTAIL.t8 24.8135
R102 VTAIL.n8 VTAIL.t6 24.8135
R103 VTAIL.n5 VTAIL.t5 24.8135
R104 VTAIL.n5 VTAIL.t0 24.8135
R105 VTAIL.n6 VTAIL.n4 20.7203
R106 VTAIL.n11 VTAIL.n10 17.1083
R107 VTAIL.n7 VTAIL.n6 3.61257
R108 VTAIL.n10 VTAIL.n9 3.61257
R109 VTAIL.n4 VTAIL.n2 3.61257
R110 VTAIL VTAIL.n11 2.65136
R111 VTAIL.n9 VTAIL.n7 2.27636
R112 VTAIL.n2 VTAIL.n1 2.27636
R113 VTAIL VTAIL.n1 0.961707
R114 VDD1 VDD1.t5 392.728
R115 VDD1.n1 VDD1.t4 392.613
R116 VDD1.n1 VDD1.n0 347.872
R117 VDD1.n3 VDD1.n2 347.024
R118 VDD1.n3 VDD1.n1 38.9729
R119 VDD1.n2 VDD1.t3 24.8135
R120 VDD1.n2 VDD1.t2 24.8135
R121 VDD1.n0 VDD1.t1 24.8135
R122 VDD1.n0 VDD1.t0 24.8135
R123 VDD1 VDD1.n3 0.845328
R124 VN.n37 VN.n20 161.3
R125 VN.n36 VN.n35 161.3
R126 VN.n34 VN.n21 161.3
R127 VN.n33 VN.n32 161.3
R128 VN.n31 VN.n22 161.3
R129 VN.n30 VN.n29 161.3
R130 VN.n28 VN.n23 161.3
R131 VN.n27 VN.n26 161.3
R132 VN.n17 VN.n0 161.3
R133 VN.n16 VN.n15 161.3
R134 VN.n14 VN.n1 161.3
R135 VN.n13 VN.n12 161.3
R136 VN.n11 VN.n2 161.3
R137 VN.n10 VN.n9 161.3
R138 VN.n8 VN.n3 161.3
R139 VN.n7 VN.n6 161.3
R140 VN.n5 VN.n4 62.8644
R141 VN.n25 VN.n24 62.8644
R142 VN.n19 VN.n18 60.6508
R143 VN.n39 VN.n38 60.6508
R144 VN.n12 VN.n11 55.548
R145 VN.n32 VN.n31 55.548
R146 VN VN.n39 45.7882
R147 VN.n4 VN.t3 40.3868
R148 VN.n24 VN.t1 40.3868
R149 VN.n12 VN.n1 25.4388
R150 VN.n32 VN.n21 25.4388
R151 VN.n6 VN.n3 24.4675
R152 VN.n10 VN.n3 24.4675
R153 VN.n11 VN.n10 24.4675
R154 VN.n16 VN.n1 24.4675
R155 VN.n17 VN.n16 24.4675
R156 VN.n31 VN.n30 24.4675
R157 VN.n30 VN.n23 24.4675
R158 VN.n26 VN.n23 24.4675
R159 VN.n37 VN.n36 24.4675
R160 VN.n36 VN.n21 24.4675
R161 VN.n18 VN.n17 21.5315
R162 VN.n38 VN.n37 21.5315
R163 VN.n6 VN.n5 12.234
R164 VN.n26 VN.n25 12.234
R165 VN.n5 VN.t5 8.17952
R166 VN.n18 VN.t2 8.17952
R167 VN.n25 VN.t4 8.17952
R168 VN.n38 VN.t0 8.17952
R169 VN.n27 VN.n24 2.63953
R170 VN.n7 VN.n4 2.63953
R171 VN.n39 VN.n20 0.417535
R172 VN.n19 VN.n0 0.417535
R173 VN VN.n19 0.394291
R174 VN.n35 VN.n20 0.189894
R175 VN.n35 VN.n34 0.189894
R176 VN.n34 VN.n33 0.189894
R177 VN.n33 VN.n22 0.189894
R178 VN.n29 VN.n22 0.189894
R179 VN.n29 VN.n28 0.189894
R180 VN.n28 VN.n27 0.189894
R181 VN.n8 VN.n7 0.189894
R182 VN.n9 VN.n8 0.189894
R183 VN.n9 VN.n2 0.189894
R184 VN.n13 VN.n2 0.189894
R185 VN.n14 VN.n13 0.189894
R186 VN.n15 VN.n14 0.189894
R187 VN.n15 VN.n0 0.189894
R188 VDD2.n1 VDD2.t2 392.613
R189 VDD2.n2 VDD2.t5 389.961
R190 VDD2.n1 VDD2.n0 347.872
R191 VDD2 VDD2.n3 347.868
R192 VDD2.n2 VDD2.n1 36.5838
R193 VDD2.n3 VDD2.t1 24.8135
R194 VDD2.n3 VDD2.t4 24.8135
R195 VDD2.n0 VDD2.t0 24.8135
R196 VDD2.n0 VDD2.t3 24.8135
R197 VDD2 VDD2.n2 2.76774
R198 B.n286 B.n285 585
R199 B.n284 B.n109 585
R200 B.n283 B.n282 585
R201 B.n281 B.n110 585
R202 B.n280 B.n279 585
R203 B.n278 B.n111 585
R204 B.n277 B.n276 585
R205 B.n275 B.n112 585
R206 B.n274 B.n273 585
R207 B.n272 B.n113 585
R208 B.n271 B.n270 585
R209 B.n266 B.n114 585
R210 B.n265 B.n264 585
R211 B.n263 B.n115 585
R212 B.n262 B.n261 585
R213 B.n260 B.n116 585
R214 B.n259 B.n258 585
R215 B.n257 B.n117 585
R216 B.n256 B.n255 585
R217 B.n254 B.n118 585
R218 B.n252 B.n251 585
R219 B.n250 B.n121 585
R220 B.n249 B.n248 585
R221 B.n247 B.n122 585
R222 B.n246 B.n245 585
R223 B.n244 B.n123 585
R224 B.n243 B.n242 585
R225 B.n241 B.n124 585
R226 B.n240 B.n239 585
R227 B.n238 B.n125 585
R228 B.n287 B.n108 585
R229 B.n289 B.n288 585
R230 B.n290 B.n107 585
R231 B.n292 B.n291 585
R232 B.n293 B.n106 585
R233 B.n295 B.n294 585
R234 B.n296 B.n105 585
R235 B.n298 B.n297 585
R236 B.n299 B.n104 585
R237 B.n301 B.n300 585
R238 B.n302 B.n103 585
R239 B.n304 B.n303 585
R240 B.n305 B.n102 585
R241 B.n307 B.n306 585
R242 B.n308 B.n101 585
R243 B.n310 B.n309 585
R244 B.n311 B.n100 585
R245 B.n313 B.n312 585
R246 B.n314 B.n99 585
R247 B.n316 B.n315 585
R248 B.n317 B.n98 585
R249 B.n319 B.n318 585
R250 B.n320 B.n97 585
R251 B.n322 B.n321 585
R252 B.n323 B.n96 585
R253 B.n325 B.n324 585
R254 B.n326 B.n95 585
R255 B.n328 B.n327 585
R256 B.n329 B.n94 585
R257 B.n331 B.n330 585
R258 B.n332 B.n93 585
R259 B.n334 B.n333 585
R260 B.n335 B.n92 585
R261 B.n337 B.n336 585
R262 B.n338 B.n91 585
R263 B.n340 B.n339 585
R264 B.n341 B.n90 585
R265 B.n343 B.n342 585
R266 B.n344 B.n89 585
R267 B.n346 B.n345 585
R268 B.n347 B.n88 585
R269 B.n349 B.n348 585
R270 B.n350 B.n87 585
R271 B.n352 B.n351 585
R272 B.n353 B.n86 585
R273 B.n355 B.n354 585
R274 B.n356 B.n85 585
R275 B.n358 B.n357 585
R276 B.n359 B.n84 585
R277 B.n361 B.n360 585
R278 B.n362 B.n83 585
R279 B.n364 B.n363 585
R280 B.n365 B.n82 585
R281 B.n367 B.n366 585
R282 B.n368 B.n81 585
R283 B.n370 B.n369 585
R284 B.n371 B.n80 585
R285 B.n373 B.n372 585
R286 B.n374 B.n79 585
R287 B.n376 B.n375 585
R288 B.n377 B.n78 585
R289 B.n379 B.n378 585
R290 B.n380 B.n77 585
R291 B.n382 B.n381 585
R292 B.n383 B.n76 585
R293 B.n385 B.n384 585
R294 B.n386 B.n75 585
R295 B.n388 B.n387 585
R296 B.n389 B.n74 585
R297 B.n391 B.n390 585
R298 B.n392 B.n73 585
R299 B.n394 B.n393 585
R300 B.n395 B.n72 585
R301 B.n397 B.n396 585
R302 B.n398 B.n71 585
R303 B.n400 B.n399 585
R304 B.n401 B.n70 585
R305 B.n403 B.n402 585
R306 B.n404 B.n69 585
R307 B.n406 B.n405 585
R308 B.n407 B.n68 585
R309 B.n409 B.n408 585
R310 B.n410 B.n67 585
R311 B.n412 B.n411 585
R312 B.n413 B.n66 585
R313 B.n415 B.n414 585
R314 B.n416 B.n65 585
R315 B.n418 B.n417 585
R316 B.n419 B.n64 585
R317 B.n421 B.n420 585
R318 B.n422 B.n63 585
R319 B.n424 B.n423 585
R320 B.n425 B.n62 585
R321 B.n427 B.n426 585
R322 B.n428 B.n61 585
R323 B.n430 B.n429 585
R324 B.n431 B.n60 585
R325 B.n433 B.n432 585
R326 B.n434 B.n59 585
R327 B.n436 B.n435 585
R328 B.n437 B.n58 585
R329 B.n439 B.n438 585
R330 B.n440 B.n57 585
R331 B.n442 B.n441 585
R332 B.n443 B.n56 585
R333 B.n445 B.n444 585
R334 B.n446 B.n55 585
R335 B.n448 B.n447 585
R336 B.n449 B.n54 585
R337 B.n451 B.n450 585
R338 B.n452 B.n53 585
R339 B.n454 B.n453 585
R340 B.n455 B.n52 585
R341 B.n457 B.n456 585
R342 B.n458 B.n51 585
R343 B.n460 B.n459 585
R344 B.n506 B.n505 585
R345 B.n504 B.n31 585
R346 B.n503 B.n502 585
R347 B.n501 B.n32 585
R348 B.n500 B.n499 585
R349 B.n498 B.n33 585
R350 B.n497 B.n496 585
R351 B.n495 B.n34 585
R352 B.n494 B.n493 585
R353 B.n492 B.n35 585
R354 B.n490 B.n489 585
R355 B.n488 B.n38 585
R356 B.n487 B.n486 585
R357 B.n485 B.n39 585
R358 B.n484 B.n483 585
R359 B.n482 B.n40 585
R360 B.n481 B.n480 585
R361 B.n479 B.n41 585
R362 B.n478 B.n477 585
R363 B.n476 B.n42 585
R364 B.n475 B.n474 585
R365 B.n473 B.n43 585
R366 B.n472 B.n471 585
R367 B.n470 B.n47 585
R368 B.n469 B.n468 585
R369 B.n467 B.n48 585
R370 B.n466 B.n465 585
R371 B.n464 B.n49 585
R372 B.n463 B.n462 585
R373 B.n461 B.n50 585
R374 B.n507 B.n30 585
R375 B.n509 B.n508 585
R376 B.n510 B.n29 585
R377 B.n512 B.n511 585
R378 B.n513 B.n28 585
R379 B.n515 B.n514 585
R380 B.n516 B.n27 585
R381 B.n518 B.n517 585
R382 B.n519 B.n26 585
R383 B.n521 B.n520 585
R384 B.n522 B.n25 585
R385 B.n524 B.n523 585
R386 B.n525 B.n24 585
R387 B.n527 B.n526 585
R388 B.n528 B.n23 585
R389 B.n530 B.n529 585
R390 B.n531 B.n22 585
R391 B.n533 B.n532 585
R392 B.n534 B.n21 585
R393 B.n536 B.n535 585
R394 B.n537 B.n20 585
R395 B.n539 B.n538 585
R396 B.n540 B.n19 585
R397 B.n542 B.n541 585
R398 B.n543 B.n18 585
R399 B.n545 B.n544 585
R400 B.n546 B.n17 585
R401 B.n548 B.n547 585
R402 B.n549 B.n16 585
R403 B.n551 B.n550 585
R404 B.n552 B.n15 585
R405 B.n554 B.n553 585
R406 B.n555 B.n14 585
R407 B.n557 B.n556 585
R408 B.n558 B.n13 585
R409 B.n560 B.n559 585
R410 B.n561 B.n12 585
R411 B.n563 B.n562 585
R412 B.n564 B.n11 585
R413 B.n566 B.n565 585
R414 B.n567 B.n10 585
R415 B.n569 B.n568 585
R416 B.n570 B.n9 585
R417 B.n572 B.n571 585
R418 B.n573 B.n8 585
R419 B.n575 B.n574 585
R420 B.n576 B.n7 585
R421 B.n578 B.n577 585
R422 B.n579 B.n6 585
R423 B.n581 B.n580 585
R424 B.n582 B.n5 585
R425 B.n584 B.n583 585
R426 B.n585 B.n4 585
R427 B.n587 B.n586 585
R428 B.n588 B.n3 585
R429 B.n590 B.n589 585
R430 B.n591 B.n0 585
R431 B.n2 B.n1 585
R432 B.n154 B.n153 585
R433 B.n156 B.n155 585
R434 B.n157 B.n152 585
R435 B.n159 B.n158 585
R436 B.n160 B.n151 585
R437 B.n162 B.n161 585
R438 B.n163 B.n150 585
R439 B.n165 B.n164 585
R440 B.n166 B.n149 585
R441 B.n168 B.n167 585
R442 B.n169 B.n148 585
R443 B.n171 B.n170 585
R444 B.n172 B.n147 585
R445 B.n174 B.n173 585
R446 B.n175 B.n146 585
R447 B.n177 B.n176 585
R448 B.n178 B.n145 585
R449 B.n180 B.n179 585
R450 B.n181 B.n144 585
R451 B.n183 B.n182 585
R452 B.n184 B.n143 585
R453 B.n186 B.n185 585
R454 B.n187 B.n142 585
R455 B.n189 B.n188 585
R456 B.n190 B.n141 585
R457 B.n192 B.n191 585
R458 B.n193 B.n140 585
R459 B.n195 B.n194 585
R460 B.n196 B.n139 585
R461 B.n198 B.n197 585
R462 B.n199 B.n138 585
R463 B.n201 B.n200 585
R464 B.n202 B.n137 585
R465 B.n204 B.n203 585
R466 B.n205 B.n136 585
R467 B.n207 B.n206 585
R468 B.n208 B.n135 585
R469 B.n210 B.n209 585
R470 B.n211 B.n134 585
R471 B.n213 B.n212 585
R472 B.n214 B.n133 585
R473 B.n216 B.n215 585
R474 B.n217 B.n132 585
R475 B.n219 B.n218 585
R476 B.n220 B.n131 585
R477 B.n222 B.n221 585
R478 B.n223 B.n130 585
R479 B.n225 B.n224 585
R480 B.n226 B.n129 585
R481 B.n228 B.n227 585
R482 B.n229 B.n128 585
R483 B.n231 B.n230 585
R484 B.n232 B.n127 585
R485 B.n234 B.n233 585
R486 B.n235 B.n126 585
R487 B.n237 B.n236 585
R488 B.n238 B.n237 478.086
R489 B.n285 B.n108 478.086
R490 B.n459 B.n50 478.086
R491 B.n507 B.n506 478.086
R492 B.n119 B.t1 448.471
R493 B.n267 B.t10 448.471
R494 B.n44 B.t8 448.471
R495 B.n36 B.t5 448.471
R496 B.n120 B.t2 367.212
R497 B.n268 B.t11 367.212
R498 B.n45 B.t7 367.212
R499 B.n37 B.t4 367.212
R500 B.n593 B.n592 256.663
R501 B.n592 B.n591 235.042
R502 B.n592 B.n2 235.042
R503 B.n119 B.t0 209.897
R504 B.n267 B.t9 209.897
R505 B.n44 B.t6 209.897
R506 B.n36 B.t3 209.897
R507 B.n239 B.n238 163.367
R508 B.n239 B.n124 163.367
R509 B.n243 B.n124 163.367
R510 B.n244 B.n243 163.367
R511 B.n245 B.n244 163.367
R512 B.n245 B.n122 163.367
R513 B.n249 B.n122 163.367
R514 B.n250 B.n249 163.367
R515 B.n251 B.n250 163.367
R516 B.n251 B.n118 163.367
R517 B.n256 B.n118 163.367
R518 B.n257 B.n256 163.367
R519 B.n258 B.n257 163.367
R520 B.n258 B.n116 163.367
R521 B.n262 B.n116 163.367
R522 B.n263 B.n262 163.367
R523 B.n264 B.n263 163.367
R524 B.n264 B.n114 163.367
R525 B.n271 B.n114 163.367
R526 B.n272 B.n271 163.367
R527 B.n273 B.n272 163.367
R528 B.n273 B.n112 163.367
R529 B.n277 B.n112 163.367
R530 B.n278 B.n277 163.367
R531 B.n279 B.n278 163.367
R532 B.n279 B.n110 163.367
R533 B.n283 B.n110 163.367
R534 B.n284 B.n283 163.367
R535 B.n285 B.n284 163.367
R536 B.n459 B.n458 163.367
R537 B.n458 B.n457 163.367
R538 B.n457 B.n52 163.367
R539 B.n453 B.n52 163.367
R540 B.n453 B.n452 163.367
R541 B.n452 B.n451 163.367
R542 B.n451 B.n54 163.367
R543 B.n447 B.n54 163.367
R544 B.n447 B.n446 163.367
R545 B.n446 B.n445 163.367
R546 B.n445 B.n56 163.367
R547 B.n441 B.n56 163.367
R548 B.n441 B.n440 163.367
R549 B.n440 B.n439 163.367
R550 B.n439 B.n58 163.367
R551 B.n435 B.n58 163.367
R552 B.n435 B.n434 163.367
R553 B.n434 B.n433 163.367
R554 B.n433 B.n60 163.367
R555 B.n429 B.n60 163.367
R556 B.n429 B.n428 163.367
R557 B.n428 B.n427 163.367
R558 B.n427 B.n62 163.367
R559 B.n423 B.n62 163.367
R560 B.n423 B.n422 163.367
R561 B.n422 B.n421 163.367
R562 B.n421 B.n64 163.367
R563 B.n417 B.n64 163.367
R564 B.n417 B.n416 163.367
R565 B.n416 B.n415 163.367
R566 B.n415 B.n66 163.367
R567 B.n411 B.n66 163.367
R568 B.n411 B.n410 163.367
R569 B.n410 B.n409 163.367
R570 B.n409 B.n68 163.367
R571 B.n405 B.n68 163.367
R572 B.n405 B.n404 163.367
R573 B.n404 B.n403 163.367
R574 B.n403 B.n70 163.367
R575 B.n399 B.n70 163.367
R576 B.n399 B.n398 163.367
R577 B.n398 B.n397 163.367
R578 B.n397 B.n72 163.367
R579 B.n393 B.n72 163.367
R580 B.n393 B.n392 163.367
R581 B.n392 B.n391 163.367
R582 B.n391 B.n74 163.367
R583 B.n387 B.n74 163.367
R584 B.n387 B.n386 163.367
R585 B.n386 B.n385 163.367
R586 B.n385 B.n76 163.367
R587 B.n381 B.n76 163.367
R588 B.n381 B.n380 163.367
R589 B.n380 B.n379 163.367
R590 B.n379 B.n78 163.367
R591 B.n375 B.n78 163.367
R592 B.n375 B.n374 163.367
R593 B.n374 B.n373 163.367
R594 B.n373 B.n80 163.367
R595 B.n369 B.n80 163.367
R596 B.n369 B.n368 163.367
R597 B.n368 B.n367 163.367
R598 B.n367 B.n82 163.367
R599 B.n363 B.n82 163.367
R600 B.n363 B.n362 163.367
R601 B.n362 B.n361 163.367
R602 B.n361 B.n84 163.367
R603 B.n357 B.n84 163.367
R604 B.n357 B.n356 163.367
R605 B.n356 B.n355 163.367
R606 B.n355 B.n86 163.367
R607 B.n351 B.n86 163.367
R608 B.n351 B.n350 163.367
R609 B.n350 B.n349 163.367
R610 B.n349 B.n88 163.367
R611 B.n345 B.n88 163.367
R612 B.n345 B.n344 163.367
R613 B.n344 B.n343 163.367
R614 B.n343 B.n90 163.367
R615 B.n339 B.n90 163.367
R616 B.n339 B.n338 163.367
R617 B.n338 B.n337 163.367
R618 B.n337 B.n92 163.367
R619 B.n333 B.n92 163.367
R620 B.n333 B.n332 163.367
R621 B.n332 B.n331 163.367
R622 B.n331 B.n94 163.367
R623 B.n327 B.n94 163.367
R624 B.n327 B.n326 163.367
R625 B.n326 B.n325 163.367
R626 B.n325 B.n96 163.367
R627 B.n321 B.n96 163.367
R628 B.n321 B.n320 163.367
R629 B.n320 B.n319 163.367
R630 B.n319 B.n98 163.367
R631 B.n315 B.n98 163.367
R632 B.n315 B.n314 163.367
R633 B.n314 B.n313 163.367
R634 B.n313 B.n100 163.367
R635 B.n309 B.n100 163.367
R636 B.n309 B.n308 163.367
R637 B.n308 B.n307 163.367
R638 B.n307 B.n102 163.367
R639 B.n303 B.n102 163.367
R640 B.n303 B.n302 163.367
R641 B.n302 B.n301 163.367
R642 B.n301 B.n104 163.367
R643 B.n297 B.n104 163.367
R644 B.n297 B.n296 163.367
R645 B.n296 B.n295 163.367
R646 B.n295 B.n106 163.367
R647 B.n291 B.n106 163.367
R648 B.n291 B.n290 163.367
R649 B.n290 B.n289 163.367
R650 B.n289 B.n108 163.367
R651 B.n506 B.n31 163.367
R652 B.n502 B.n31 163.367
R653 B.n502 B.n501 163.367
R654 B.n501 B.n500 163.367
R655 B.n500 B.n33 163.367
R656 B.n496 B.n33 163.367
R657 B.n496 B.n495 163.367
R658 B.n495 B.n494 163.367
R659 B.n494 B.n35 163.367
R660 B.n489 B.n35 163.367
R661 B.n489 B.n488 163.367
R662 B.n488 B.n487 163.367
R663 B.n487 B.n39 163.367
R664 B.n483 B.n39 163.367
R665 B.n483 B.n482 163.367
R666 B.n482 B.n481 163.367
R667 B.n481 B.n41 163.367
R668 B.n477 B.n41 163.367
R669 B.n477 B.n476 163.367
R670 B.n476 B.n475 163.367
R671 B.n475 B.n43 163.367
R672 B.n471 B.n43 163.367
R673 B.n471 B.n470 163.367
R674 B.n470 B.n469 163.367
R675 B.n469 B.n48 163.367
R676 B.n465 B.n48 163.367
R677 B.n465 B.n464 163.367
R678 B.n464 B.n463 163.367
R679 B.n463 B.n50 163.367
R680 B.n508 B.n507 163.367
R681 B.n508 B.n29 163.367
R682 B.n512 B.n29 163.367
R683 B.n513 B.n512 163.367
R684 B.n514 B.n513 163.367
R685 B.n514 B.n27 163.367
R686 B.n518 B.n27 163.367
R687 B.n519 B.n518 163.367
R688 B.n520 B.n519 163.367
R689 B.n520 B.n25 163.367
R690 B.n524 B.n25 163.367
R691 B.n525 B.n524 163.367
R692 B.n526 B.n525 163.367
R693 B.n526 B.n23 163.367
R694 B.n530 B.n23 163.367
R695 B.n531 B.n530 163.367
R696 B.n532 B.n531 163.367
R697 B.n532 B.n21 163.367
R698 B.n536 B.n21 163.367
R699 B.n537 B.n536 163.367
R700 B.n538 B.n537 163.367
R701 B.n538 B.n19 163.367
R702 B.n542 B.n19 163.367
R703 B.n543 B.n542 163.367
R704 B.n544 B.n543 163.367
R705 B.n544 B.n17 163.367
R706 B.n548 B.n17 163.367
R707 B.n549 B.n548 163.367
R708 B.n550 B.n549 163.367
R709 B.n550 B.n15 163.367
R710 B.n554 B.n15 163.367
R711 B.n555 B.n554 163.367
R712 B.n556 B.n555 163.367
R713 B.n556 B.n13 163.367
R714 B.n560 B.n13 163.367
R715 B.n561 B.n560 163.367
R716 B.n562 B.n561 163.367
R717 B.n562 B.n11 163.367
R718 B.n566 B.n11 163.367
R719 B.n567 B.n566 163.367
R720 B.n568 B.n567 163.367
R721 B.n568 B.n9 163.367
R722 B.n572 B.n9 163.367
R723 B.n573 B.n572 163.367
R724 B.n574 B.n573 163.367
R725 B.n574 B.n7 163.367
R726 B.n578 B.n7 163.367
R727 B.n579 B.n578 163.367
R728 B.n580 B.n579 163.367
R729 B.n580 B.n5 163.367
R730 B.n584 B.n5 163.367
R731 B.n585 B.n584 163.367
R732 B.n586 B.n585 163.367
R733 B.n586 B.n3 163.367
R734 B.n590 B.n3 163.367
R735 B.n591 B.n590 163.367
R736 B.n154 B.n2 163.367
R737 B.n155 B.n154 163.367
R738 B.n155 B.n152 163.367
R739 B.n159 B.n152 163.367
R740 B.n160 B.n159 163.367
R741 B.n161 B.n160 163.367
R742 B.n161 B.n150 163.367
R743 B.n165 B.n150 163.367
R744 B.n166 B.n165 163.367
R745 B.n167 B.n166 163.367
R746 B.n167 B.n148 163.367
R747 B.n171 B.n148 163.367
R748 B.n172 B.n171 163.367
R749 B.n173 B.n172 163.367
R750 B.n173 B.n146 163.367
R751 B.n177 B.n146 163.367
R752 B.n178 B.n177 163.367
R753 B.n179 B.n178 163.367
R754 B.n179 B.n144 163.367
R755 B.n183 B.n144 163.367
R756 B.n184 B.n183 163.367
R757 B.n185 B.n184 163.367
R758 B.n185 B.n142 163.367
R759 B.n189 B.n142 163.367
R760 B.n190 B.n189 163.367
R761 B.n191 B.n190 163.367
R762 B.n191 B.n140 163.367
R763 B.n195 B.n140 163.367
R764 B.n196 B.n195 163.367
R765 B.n197 B.n196 163.367
R766 B.n197 B.n138 163.367
R767 B.n201 B.n138 163.367
R768 B.n202 B.n201 163.367
R769 B.n203 B.n202 163.367
R770 B.n203 B.n136 163.367
R771 B.n207 B.n136 163.367
R772 B.n208 B.n207 163.367
R773 B.n209 B.n208 163.367
R774 B.n209 B.n134 163.367
R775 B.n213 B.n134 163.367
R776 B.n214 B.n213 163.367
R777 B.n215 B.n214 163.367
R778 B.n215 B.n132 163.367
R779 B.n219 B.n132 163.367
R780 B.n220 B.n219 163.367
R781 B.n221 B.n220 163.367
R782 B.n221 B.n130 163.367
R783 B.n225 B.n130 163.367
R784 B.n226 B.n225 163.367
R785 B.n227 B.n226 163.367
R786 B.n227 B.n128 163.367
R787 B.n231 B.n128 163.367
R788 B.n232 B.n231 163.367
R789 B.n233 B.n232 163.367
R790 B.n233 B.n126 163.367
R791 B.n237 B.n126 163.367
R792 B.n120 B.n119 81.2611
R793 B.n268 B.n267 81.2611
R794 B.n45 B.n44 81.2611
R795 B.n37 B.n36 81.2611
R796 B.n253 B.n120 59.5399
R797 B.n269 B.n268 59.5399
R798 B.n46 B.n45 59.5399
R799 B.n491 B.n37 59.5399
R800 B.n505 B.n30 31.0639
R801 B.n461 B.n460 31.0639
R802 B.n287 B.n286 31.0639
R803 B.n236 B.n125 31.0639
R804 B B.n593 18.0485
R805 B.n509 B.n30 10.6151
R806 B.n510 B.n509 10.6151
R807 B.n511 B.n510 10.6151
R808 B.n511 B.n28 10.6151
R809 B.n515 B.n28 10.6151
R810 B.n516 B.n515 10.6151
R811 B.n517 B.n516 10.6151
R812 B.n517 B.n26 10.6151
R813 B.n521 B.n26 10.6151
R814 B.n522 B.n521 10.6151
R815 B.n523 B.n522 10.6151
R816 B.n523 B.n24 10.6151
R817 B.n527 B.n24 10.6151
R818 B.n528 B.n527 10.6151
R819 B.n529 B.n528 10.6151
R820 B.n529 B.n22 10.6151
R821 B.n533 B.n22 10.6151
R822 B.n534 B.n533 10.6151
R823 B.n535 B.n534 10.6151
R824 B.n535 B.n20 10.6151
R825 B.n539 B.n20 10.6151
R826 B.n540 B.n539 10.6151
R827 B.n541 B.n540 10.6151
R828 B.n541 B.n18 10.6151
R829 B.n545 B.n18 10.6151
R830 B.n546 B.n545 10.6151
R831 B.n547 B.n546 10.6151
R832 B.n547 B.n16 10.6151
R833 B.n551 B.n16 10.6151
R834 B.n552 B.n551 10.6151
R835 B.n553 B.n552 10.6151
R836 B.n553 B.n14 10.6151
R837 B.n557 B.n14 10.6151
R838 B.n558 B.n557 10.6151
R839 B.n559 B.n558 10.6151
R840 B.n559 B.n12 10.6151
R841 B.n563 B.n12 10.6151
R842 B.n564 B.n563 10.6151
R843 B.n565 B.n564 10.6151
R844 B.n565 B.n10 10.6151
R845 B.n569 B.n10 10.6151
R846 B.n570 B.n569 10.6151
R847 B.n571 B.n570 10.6151
R848 B.n571 B.n8 10.6151
R849 B.n575 B.n8 10.6151
R850 B.n576 B.n575 10.6151
R851 B.n577 B.n576 10.6151
R852 B.n577 B.n6 10.6151
R853 B.n581 B.n6 10.6151
R854 B.n582 B.n581 10.6151
R855 B.n583 B.n582 10.6151
R856 B.n583 B.n4 10.6151
R857 B.n587 B.n4 10.6151
R858 B.n588 B.n587 10.6151
R859 B.n589 B.n588 10.6151
R860 B.n589 B.n0 10.6151
R861 B.n505 B.n504 10.6151
R862 B.n504 B.n503 10.6151
R863 B.n503 B.n32 10.6151
R864 B.n499 B.n32 10.6151
R865 B.n499 B.n498 10.6151
R866 B.n498 B.n497 10.6151
R867 B.n497 B.n34 10.6151
R868 B.n493 B.n34 10.6151
R869 B.n493 B.n492 10.6151
R870 B.n490 B.n38 10.6151
R871 B.n486 B.n38 10.6151
R872 B.n486 B.n485 10.6151
R873 B.n485 B.n484 10.6151
R874 B.n484 B.n40 10.6151
R875 B.n480 B.n40 10.6151
R876 B.n480 B.n479 10.6151
R877 B.n479 B.n478 10.6151
R878 B.n478 B.n42 10.6151
R879 B.n474 B.n473 10.6151
R880 B.n473 B.n472 10.6151
R881 B.n472 B.n47 10.6151
R882 B.n468 B.n47 10.6151
R883 B.n468 B.n467 10.6151
R884 B.n467 B.n466 10.6151
R885 B.n466 B.n49 10.6151
R886 B.n462 B.n49 10.6151
R887 B.n462 B.n461 10.6151
R888 B.n460 B.n51 10.6151
R889 B.n456 B.n51 10.6151
R890 B.n456 B.n455 10.6151
R891 B.n455 B.n454 10.6151
R892 B.n454 B.n53 10.6151
R893 B.n450 B.n53 10.6151
R894 B.n450 B.n449 10.6151
R895 B.n449 B.n448 10.6151
R896 B.n448 B.n55 10.6151
R897 B.n444 B.n55 10.6151
R898 B.n444 B.n443 10.6151
R899 B.n443 B.n442 10.6151
R900 B.n442 B.n57 10.6151
R901 B.n438 B.n57 10.6151
R902 B.n438 B.n437 10.6151
R903 B.n437 B.n436 10.6151
R904 B.n436 B.n59 10.6151
R905 B.n432 B.n59 10.6151
R906 B.n432 B.n431 10.6151
R907 B.n431 B.n430 10.6151
R908 B.n430 B.n61 10.6151
R909 B.n426 B.n61 10.6151
R910 B.n426 B.n425 10.6151
R911 B.n425 B.n424 10.6151
R912 B.n424 B.n63 10.6151
R913 B.n420 B.n63 10.6151
R914 B.n420 B.n419 10.6151
R915 B.n419 B.n418 10.6151
R916 B.n418 B.n65 10.6151
R917 B.n414 B.n65 10.6151
R918 B.n414 B.n413 10.6151
R919 B.n413 B.n412 10.6151
R920 B.n412 B.n67 10.6151
R921 B.n408 B.n67 10.6151
R922 B.n408 B.n407 10.6151
R923 B.n407 B.n406 10.6151
R924 B.n406 B.n69 10.6151
R925 B.n402 B.n69 10.6151
R926 B.n402 B.n401 10.6151
R927 B.n401 B.n400 10.6151
R928 B.n400 B.n71 10.6151
R929 B.n396 B.n71 10.6151
R930 B.n396 B.n395 10.6151
R931 B.n395 B.n394 10.6151
R932 B.n394 B.n73 10.6151
R933 B.n390 B.n73 10.6151
R934 B.n390 B.n389 10.6151
R935 B.n389 B.n388 10.6151
R936 B.n388 B.n75 10.6151
R937 B.n384 B.n75 10.6151
R938 B.n384 B.n383 10.6151
R939 B.n383 B.n382 10.6151
R940 B.n382 B.n77 10.6151
R941 B.n378 B.n77 10.6151
R942 B.n378 B.n377 10.6151
R943 B.n377 B.n376 10.6151
R944 B.n376 B.n79 10.6151
R945 B.n372 B.n79 10.6151
R946 B.n372 B.n371 10.6151
R947 B.n371 B.n370 10.6151
R948 B.n370 B.n81 10.6151
R949 B.n366 B.n81 10.6151
R950 B.n366 B.n365 10.6151
R951 B.n365 B.n364 10.6151
R952 B.n364 B.n83 10.6151
R953 B.n360 B.n83 10.6151
R954 B.n360 B.n359 10.6151
R955 B.n359 B.n358 10.6151
R956 B.n358 B.n85 10.6151
R957 B.n354 B.n85 10.6151
R958 B.n354 B.n353 10.6151
R959 B.n353 B.n352 10.6151
R960 B.n352 B.n87 10.6151
R961 B.n348 B.n87 10.6151
R962 B.n348 B.n347 10.6151
R963 B.n347 B.n346 10.6151
R964 B.n346 B.n89 10.6151
R965 B.n342 B.n89 10.6151
R966 B.n342 B.n341 10.6151
R967 B.n341 B.n340 10.6151
R968 B.n340 B.n91 10.6151
R969 B.n336 B.n91 10.6151
R970 B.n336 B.n335 10.6151
R971 B.n335 B.n334 10.6151
R972 B.n334 B.n93 10.6151
R973 B.n330 B.n93 10.6151
R974 B.n330 B.n329 10.6151
R975 B.n329 B.n328 10.6151
R976 B.n328 B.n95 10.6151
R977 B.n324 B.n95 10.6151
R978 B.n324 B.n323 10.6151
R979 B.n323 B.n322 10.6151
R980 B.n322 B.n97 10.6151
R981 B.n318 B.n97 10.6151
R982 B.n318 B.n317 10.6151
R983 B.n317 B.n316 10.6151
R984 B.n316 B.n99 10.6151
R985 B.n312 B.n99 10.6151
R986 B.n312 B.n311 10.6151
R987 B.n311 B.n310 10.6151
R988 B.n310 B.n101 10.6151
R989 B.n306 B.n101 10.6151
R990 B.n306 B.n305 10.6151
R991 B.n305 B.n304 10.6151
R992 B.n304 B.n103 10.6151
R993 B.n300 B.n103 10.6151
R994 B.n300 B.n299 10.6151
R995 B.n299 B.n298 10.6151
R996 B.n298 B.n105 10.6151
R997 B.n294 B.n105 10.6151
R998 B.n294 B.n293 10.6151
R999 B.n293 B.n292 10.6151
R1000 B.n292 B.n107 10.6151
R1001 B.n288 B.n107 10.6151
R1002 B.n288 B.n287 10.6151
R1003 B.n153 B.n1 10.6151
R1004 B.n156 B.n153 10.6151
R1005 B.n157 B.n156 10.6151
R1006 B.n158 B.n157 10.6151
R1007 B.n158 B.n151 10.6151
R1008 B.n162 B.n151 10.6151
R1009 B.n163 B.n162 10.6151
R1010 B.n164 B.n163 10.6151
R1011 B.n164 B.n149 10.6151
R1012 B.n168 B.n149 10.6151
R1013 B.n169 B.n168 10.6151
R1014 B.n170 B.n169 10.6151
R1015 B.n170 B.n147 10.6151
R1016 B.n174 B.n147 10.6151
R1017 B.n175 B.n174 10.6151
R1018 B.n176 B.n175 10.6151
R1019 B.n176 B.n145 10.6151
R1020 B.n180 B.n145 10.6151
R1021 B.n181 B.n180 10.6151
R1022 B.n182 B.n181 10.6151
R1023 B.n182 B.n143 10.6151
R1024 B.n186 B.n143 10.6151
R1025 B.n187 B.n186 10.6151
R1026 B.n188 B.n187 10.6151
R1027 B.n188 B.n141 10.6151
R1028 B.n192 B.n141 10.6151
R1029 B.n193 B.n192 10.6151
R1030 B.n194 B.n193 10.6151
R1031 B.n194 B.n139 10.6151
R1032 B.n198 B.n139 10.6151
R1033 B.n199 B.n198 10.6151
R1034 B.n200 B.n199 10.6151
R1035 B.n200 B.n137 10.6151
R1036 B.n204 B.n137 10.6151
R1037 B.n205 B.n204 10.6151
R1038 B.n206 B.n205 10.6151
R1039 B.n206 B.n135 10.6151
R1040 B.n210 B.n135 10.6151
R1041 B.n211 B.n210 10.6151
R1042 B.n212 B.n211 10.6151
R1043 B.n212 B.n133 10.6151
R1044 B.n216 B.n133 10.6151
R1045 B.n217 B.n216 10.6151
R1046 B.n218 B.n217 10.6151
R1047 B.n218 B.n131 10.6151
R1048 B.n222 B.n131 10.6151
R1049 B.n223 B.n222 10.6151
R1050 B.n224 B.n223 10.6151
R1051 B.n224 B.n129 10.6151
R1052 B.n228 B.n129 10.6151
R1053 B.n229 B.n228 10.6151
R1054 B.n230 B.n229 10.6151
R1055 B.n230 B.n127 10.6151
R1056 B.n234 B.n127 10.6151
R1057 B.n235 B.n234 10.6151
R1058 B.n236 B.n235 10.6151
R1059 B.n240 B.n125 10.6151
R1060 B.n241 B.n240 10.6151
R1061 B.n242 B.n241 10.6151
R1062 B.n242 B.n123 10.6151
R1063 B.n246 B.n123 10.6151
R1064 B.n247 B.n246 10.6151
R1065 B.n248 B.n247 10.6151
R1066 B.n248 B.n121 10.6151
R1067 B.n252 B.n121 10.6151
R1068 B.n255 B.n254 10.6151
R1069 B.n255 B.n117 10.6151
R1070 B.n259 B.n117 10.6151
R1071 B.n260 B.n259 10.6151
R1072 B.n261 B.n260 10.6151
R1073 B.n261 B.n115 10.6151
R1074 B.n265 B.n115 10.6151
R1075 B.n266 B.n265 10.6151
R1076 B.n270 B.n266 10.6151
R1077 B.n274 B.n113 10.6151
R1078 B.n275 B.n274 10.6151
R1079 B.n276 B.n275 10.6151
R1080 B.n276 B.n111 10.6151
R1081 B.n280 B.n111 10.6151
R1082 B.n281 B.n280 10.6151
R1083 B.n282 B.n281 10.6151
R1084 B.n282 B.n109 10.6151
R1085 B.n286 B.n109 10.6151
R1086 B.n492 B.n491 9.36635
R1087 B.n474 B.n46 9.36635
R1088 B.n253 B.n252 9.36635
R1089 B.n269 B.n113 9.36635
R1090 B.n593 B.n0 8.11757
R1091 B.n593 B.n1 8.11757
R1092 B.n491 B.n490 1.24928
R1093 B.n46 B.n42 1.24928
R1094 B.n254 B.n253 1.24928
R1095 B.n270 B.n269 1.24928
C0 VTAIL VN 2.54355f
C1 VTAIL w_n4322_n1230# 1.58749f
C2 VTAIL VDD2 4.86642f
C3 VTAIL B 1.40297f
C4 VDD1 VP 1.55972f
C5 VN w_n4322_n1230# 8.3296f
C6 VDD1 VTAIL 4.80451f
C7 VDD2 VN 1.1498f
C8 B VN 1.26779f
C9 VDD2 w_n4322_n1230# 1.98519f
C10 VTAIL VP 2.55773f
C11 B w_n4322_n1230# 8.52467f
C12 VDD2 B 1.65975f
C13 VDD1 VN 0.159943f
C14 VDD1 w_n4322_n1230# 1.86077f
C15 VP VN 6.18405f
C16 VDD1 VDD2 1.89842f
C17 VP w_n4322_n1230# 8.88516f
C18 VDD1 B 1.55475f
C19 VDD2 VP 0.573728f
C20 VP B 2.21186f
C21 VDD2 VSUBS 1.31372f
C22 VDD1 VSUBS 1.878151f
C23 VTAIL VSUBS 0.685573f
C24 VN VSUBS 7.50148f
C25 VP VSUBS 3.325172f
C26 B VSUBS 4.66896f
C27 w_n4322_n1230# VSUBS 68.3049f
C28 B.n0 VSUBS 0.010866f
C29 B.n1 VSUBS 0.010866f
C30 B.n2 VSUBS 0.01607f
C31 B.n3 VSUBS 0.012315f
C32 B.n4 VSUBS 0.012315f
C33 B.n5 VSUBS 0.012315f
C34 B.n6 VSUBS 0.012315f
C35 B.n7 VSUBS 0.012315f
C36 B.n8 VSUBS 0.012315f
C37 B.n9 VSUBS 0.012315f
C38 B.n10 VSUBS 0.012315f
C39 B.n11 VSUBS 0.012315f
C40 B.n12 VSUBS 0.012315f
C41 B.n13 VSUBS 0.012315f
C42 B.n14 VSUBS 0.012315f
C43 B.n15 VSUBS 0.012315f
C44 B.n16 VSUBS 0.012315f
C45 B.n17 VSUBS 0.012315f
C46 B.n18 VSUBS 0.012315f
C47 B.n19 VSUBS 0.012315f
C48 B.n20 VSUBS 0.012315f
C49 B.n21 VSUBS 0.012315f
C50 B.n22 VSUBS 0.012315f
C51 B.n23 VSUBS 0.012315f
C52 B.n24 VSUBS 0.012315f
C53 B.n25 VSUBS 0.012315f
C54 B.n26 VSUBS 0.012315f
C55 B.n27 VSUBS 0.012315f
C56 B.n28 VSUBS 0.012315f
C57 B.n29 VSUBS 0.012315f
C58 B.n30 VSUBS 0.027236f
C59 B.n31 VSUBS 0.012315f
C60 B.n32 VSUBS 0.012315f
C61 B.n33 VSUBS 0.012315f
C62 B.n34 VSUBS 0.012315f
C63 B.n35 VSUBS 0.012315f
C64 B.t4 VSUBS 0.043579f
C65 B.t5 VSUBS 0.058506f
C66 B.t3 VSUBS 0.446688f
C67 B.n36 VSUBS 0.138159f
C68 B.n37 VSUBS 0.099943f
C69 B.n38 VSUBS 0.012315f
C70 B.n39 VSUBS 0.012315f
C71 B.n40 VSUBS 0.012315f
C72 B.n41 VSUBS 0.012315f
C73 B.n42 VSUBS 0.006882f
C74 B.n43 VSUBS 0.012315f
C75 B.t7 VSUBS 0.043579f
C76 B.t8 VSUBS 0.058506f
C77 B.t6 VSUBS 0.446688f
C78 B.n44 VSUBS 0.138159f
C79 B.n45 VSUBS 0.099943f
C80 B.n46 VSUBS 0.028532f
C81 B.n47 VSUBS 0.012315f
C82 B.n48 VSUBS 0.012315f
C83 B.n49 VSUBS 0.012315f
C84 B.n50 VSUBS 0.028542f
C85 B.n51 VSUBS 0.012315f
C86 B.n52 VSUBS 0.012315f
C87 B.n53 VSUBS 0.012315f
C88 B.n54 VSUBS 0.012315f
C89 B.n55 VSUBS 0.012315f
C90 B.n56 VSUBS 0.012315f
C91 B.n57 VSUBS 0.012315f
C92 B.n58 VSUBS 0.012315f
C93 B.n59 VSUBS 0.012315f
C94 B.n60 VSUBS 0.012315f
C95 B.n61 VSUBS 0.012315f
C96 B.n62 VSUBS 0.012315f
C97 B.n63 VSUBS 0.012315f
C98 B.n64 VSUBS 0.012315f
C99 B.n65 VSUBS 0.012315f
C100 B.n66 VSUBS 0.012315f
C101 B.n67 VSUBS 0.012315f
C102 B.n68 VSUBS 0.012315f
C103 B.n69 VSUBS 0.012315f
C104 B.n70 VSUBS 0.012315f
C105 B.n71 VSUBS 0.012315f
C106 B.n72 VSUBS 0.012315f
C107 B.n73 VSUBS 0.012315f
C108 B.n74 VSUBS 0.012315f
C109 B.n75 VSUBS 0.012315f
C110 B.n76 VSUBS 0.012315f
C111 B.n77 VSUBS 0.012315f
C112 B.n78 VSUBS 0.012315f
C113 B.n79 VSUBS 0.012315f
C114 B.n80 VSUBS 0.012315f
C115 B.n81 VSUBS 0.012315f
C116 B.n82 VSUBS 0.012315f
C117 B.n83 VSUBS 0.012315f
C118 B.n84 VSUBS 0.012315f
C119 B.n85 VSUBS 0.012315f
C120 B.n86 VSUBS 0.012315f
C121 B.n87 VSUBS 0.012315f
C122 B.n88 VSUBS 0.012315f
C123 B.n89 VSUBS 0.012315f
C124 B.n90 VSUBS 0.012315f
C125 B.n91 VSUBS 0.012315f
C126 B.n92 VSUBS 0.012315f
C127 B.n93 VSUBS 0.012315f
C128 B.n94 VSUBS 0.012315f
C129 B.n95 VSUBS 0.012315f
C130 B.n96 VSUBS 0.012315f
C131 B.n97 VSUBS 0.012315f
C132 B.n98 VSUBS 0.012315f
C133 B.n99 VSUBS 0.012315f
C134 B.n100 VSUBS 0.012315f
C135 B.n101 VSUBS 0.012315f
C136 B.n102 VSUBS 0.012315f
C137 B.n103 VSUBS 0.012315f
C138 B.n104 VSUBS 0.012315f
C139 B.n105 VSUBS 0.012315f
C140 B.n106 VSUBS 0.012315f
C141 B.n107 VSUBS 0.012315f
C142 B.n108 VSUBS 0.027236f
C143 B.n109 VSUBS 0.012315f
C144 B.n110 VSUBS 0.012315f
C145 B.n111 VSUBS 0.012315f
C146 B.n112 VSUBS 0.012315f
C147 B.n113 VSUBS 0.01159f
C148 B.n114 VSUBS 0.012315f
C149 B.n115 VSUBS 0.012315f
C150 B.n116 VSUBS 0.012315f
C151 B.n117 VSUBS 0.012315f
C152 B.n118 VSUBS 0.012315f
C153 B.t2 VSUBS 0.043579f
C154 B.t1 VSUBS 0.058506f
C155 B.t0 VSUBS 0.446688f
C156 B.n119 VSUBS 0.138159f
C157 B.n120 VSUBS 0.099943f
C158 B.n121 VSUBS 0.012315f
C159 B.n122 VSUBS 0.012315f
C160 B.n123 VSUBS 0.012315f
C161 B.n124 VSUBS 0.012315f
C162 B.n125 VSUBS 0.028542f
C163 B.n126 VSUBS 0.012315f
C164 B.n127 VSUBS 0.012315f
C165 B.n128 VSUBS 0.012315f
C166 B.n129 VSUBS 0.012315f
C167 B.n130 VSUBS 0.012315f
C168 B.n131 VSUBS 0.012315f
C169 B.n132 VSUBS 0.012315f
C170 B.n133 VSUBS 0.012315f
C171 B.n134 VSUBS 0.012315f
C172 B.n135 VSUBS 0.012315f
C173 B.n136 VSUBS 0.012315f
C174 B.n137 VSUBS 0.012315f
C175 B.n138 VSUBS 0.012315f
C176 B.n139 VSUBS 0.012315f
C177 B.n140 VSUBS 0.012315f
C178 B.n141 VSUBS 0.012315f
C179 B.n142 VSUBS 0.012315f
C180 B.n143 VSUBS 0.012315f
C181 B.n144 VSUBS 0.012315f
C182 B.n145 VSUBS 0.012315f
C183 B.n146 VSUBS 0.012315f
C184 B.n147 VSUBS 0.012315f
C185 B.n148 VSUBS 0.012315f
C186 B.n149 VSUBS 0.012315f
C187 B.n150 VSUBS 0.012315f
C188 B.n151 VSUBS 0.012315f
C189 B.n152 VSUBS 0.012315f
C190 B.n153 VSUBS 0.012315f
C191 B.n154 VSUBS 0.012315f
C192 B.n155 VSUBS 0.012315f
C193 B.n156 VSUBS 0.012315f
C194 B.n157 VSUBS 0.012315f
C195 B.n158 VSUBS 0.012315f
C196 B.n159 VSUBS 0.012315f
C197 B.n160 VSUBS 0.012315f
C198 B.n161 VSUBS 0.012315f
C199 B.n162 VSUBS 0.012315f
C200 B.n163 VSUBS 0.012315f
C201 B.n164 VSUBS 0.012315f
C202 B.n165 VSUBS 0.012315f
C203 B.n166 VSUBS 0.012315f
C204 B.n167 VSUBS 0.012315f
C205 B.n168 VSUBS 0.012315f
C206 B.n169 VSUBS 0.012315f
C207 B.n170 VSUBS 0.012315f
C208 B.n171 VSUBS 0.012315f
C209 B.n172 VSUBS 0.012315f
C210 B.n173 VSUBS 0.012315f
C211 B.n174 VSUBS 0.012315f
C212 B.n175 VSUBS 0.012315f
C213 B.n176 VSUBS 0.012315f
C214 B.n177 VSUBS 0.012315f
C215 B.n178 VSUBS 0.012315f
C216 B.n179 VSUBS 0.012315f
C217 B.n180 VSUBS 0.012315f
C218 B.n181 VSUBS 0.012315f
C219 B.n182 VSUBS 0.012315f
C220 B.n183 VSUBS 0.012315f
C221 B.n184 VSUBS 0.012315f
C222 B.n185 VSUBS 0.012315f
C223 B.n186 VSUBS 0.012315f
C224 B.n187 VSUBS 0.012315f
C225 B.n188 VSUBS 0.012315f
C226 B.n189 VSUBS 0.012315f
C227 B.n190 VSUBS 0.012315f
C228 B.n191 VSUBS 0.012315f
C229 B.n192 VSUBS 0.012315f
C230 B.n193 VSUBS 0.012315f
C231 B.n194 VSUBS 0.012315f
C232 B.n195 VSUBS 0.012315f
C233 B.n196 VSUBS 0.012315f
C234 B.n197 VSUBS 0.012315f
C235 B.n198 VSUBS 0.012315f
C236 B.n199 VSUBS 0.012315f
C237 B.n200 VSUBS 0.012315f
C238 B.n201 VSUBS 0.012315f
C239 B.n202 VSUBS 0.012315f
C240 B.n203 VSUBS 0.012315f
C241 B.n204 VSUBS 0.012315f
C242 B.n205 VSUBS 0.012315f
C243 B.n206 VSUBS 0.012315f
C244 B.n207 VSUBS 0.012315f
C245 B.n208 VSUBS 0.012315f
C246 B.n209 VSUBS 0.012315f
C247 B.n210 VSUBS 0.012315f
C248 B.n211 VSUBS 0.012315f
C249 B.n212 VSUBS 0.012315f
C250 B.n213 VSUBS 0.012315f
C251 B.n214 VSUBS 0.012315f
C252 B.n215 VSUBS 0.012315f
C253 B.n216 VSUBS 0.012315f
C254 B.n217 VSUBS 0.012315f
C255 B.n218 VSUBS 0.012315f
C256 B.n219 VSUBS 0.012315f
C257 B.n220 VSUBS 0.012315f
C258 B.n221 VSUBS 0.012315f
C259 B.n222 VSUBS 0.012315f
C260 B.n223 VSUBS 0.012315f
C261 B.n224 VSUBS 0.012315f
C262 B.n225 VSUBS 0.012315f
C263 B.n226 VSUBS 0.012315f
C264 B.n227 VSUBS 0.012315f
C265 B.n228 VSUBS 0.012315f
C266 B.n229 VSUBS 0.012315f
C267 B.n230 VSUBS 0.012315f
C268 B.n231 VSUBS 0.012315f
C269 B.n232 VSUBS 0.012315f
C270 B.n233 VSUBS 0.012315f
C271 B.n234 VSUBS 0.012315f
C272 B.n235 VSUBS 0.012315f
C273 B.n236 VSUBS 0.027236f
C274 B.n237 VSUBS 0.027236f
C275 B.n238 VSUBS 0.028542f
C276 B.n239 VSUBS 0.012315f
C277 B.n240 VSUBS 0.012315f
C278 B.n241 VSUBS 0.012315f
C279 B.n242 VSUBS 0.012315f
C280 B.n243 VSUBS 0.012315f
C281 B.n244 VSUBS 0.012315f
C282 B.n245 VSUBS 0.012315f
C283 B.n246 VSUBS 0.012315f
C284 B.n247 VSUBS 0.012315f
C285 B.n248 VSUBS 0.012315f
C286 B.n249 VSUBS 0.012315f
C287 B.n250 VSUBS 0.012315f
C288 B.n251 VSUBS 0.012315f
C289 B.n252 VSUBS 0.01159f
C290 B.n253 VSUBS 0.028532f
C291 B.n254 VSUBS 0.006882f
C292 B.n255 VSUBS 0.012315f
C293 B.n256 VSUBS 0.012315f
C294 B.n257 VSUBS 0.012315f
C295 B.n258 VSUBS 0.012315f
C296 B.n259 VSUBS 0.012315f
C297 B.n260 VSUBS 0.012315f
C298 B.n261 VSUBS 0.012315f
C299 B.n262 VSUBS 0.012315f
C300 B.n263 VSUBS 0.012315f
C301 B.n264 VSUBS 0.012315f
C302 B.n265 VSUBS 0.012315f
C303 B.n266 VSUBS 0.012315f
C304 B.t11 VSUBS 0.043579f
C305 B.t10 VSUBS 0.058506f
C306 B.t9 VSUBS 0.446688f
C307 B.n267 VSUBS 0.138159f
C308 B.n268 VSUBS 0.099943f
C309 B.n269 VSUBS 0.028532f
C310 B.n270 VSUBS 0.006882f
C311 B.n271 VSUBS 0.012315f
C312 B.n272 VSUBS 0.012315f
C313 B.n273 VSUBS 0.012315f
C314 B.n274 VSUBS 0.012315f
C315 B.n275 VSUBS 0.012315f
C316 B.n276 VSUBS 0.012315f
C317 B.n277 VSUBS 0.012315f
C318 B.n278 VSUBS 0.012315f
C319 B.n279 VSUBS 0.012315f
C320 B.n280 VSUBS 0.012315f
C321 B.n281 VSUBS 0.012315f
C322 B.n282 VSUBS 0.012315f
C323 B.n283 VSUBS 0.012315f
C324 B.n284 VSUBS 0.012315f
C325 B.n285 VSUBS 0.028542f
C326 B.n286 VSUBS 0.027012f
C327 B.n287 VSUBS 0.028766f
C328 B.n288 VSUBS 0.012315f
C329 B.n289 VSUBS 0.012315f
C330 B.n290 VSUBS 0.012315f
C331 B.n291 VSUBS 0.012315f
C332 B.n292 VSUBS 0.012315f
C333 B.n293 VSUBS 0.012315f
C334 B.n294 VSUBS 0.012315f
C335 B.n295 VSUBS 0.012315f
C336 B.n296 VSUBS 0.012315f
C337 B.n297 VSUBS 0.012315f
C338 B.n298 VSUBS 0.012315f
C339 B.n299 VSUBS 0.012315f
C340 B.n300 VSUBS 0.012315f
C341 B.n301 VSUBS 0.012315f
C342 B.n302 VSUBS 0.012315f
C343 B.n303 VSUBS 0.012315f
C344 B.n304 VSUBS 0.012315f
C345 B.n305 VSUBS 0.012315f
C346 B.n306 VSUBS 0.012315f
C347 B.n307 VSUBS 0.012315f
C348 B.n308 VSUBS 0.012315f
C349 B.n309 VSUBS 0.012315f
C350 B.n310 VSUBS 0.012315f
C351 B.n311 VSUBS 0.012315f
C352 B.n312 VSUBS 0.012315f
C353 B.n313 VSUBS 0.012315f
C354 B.n314 VSUBS 0.012315f
C355 B.n315 VSUBS 0.012315f
C356 B.n316 VSUBS 0.012315f
C357 B.n317 VSUBS 0.012315f
C358 B.n318 VSUBS 0.012315f
C359 B.n319 VSUBS 0.012315f
C360 B.n320 VSUBS 0.012315f
C361 B.n321 VSUBS 0.012315f
C362 B.n322 VSUBS 0.012315f
C363 B.n323 VSUBS 0.012315f
C364 B.n324 VSUBS 0.012315f
C365 B.n325 VSUBS 0.012315f
C366 B.n326 VSUBS 0.012315f
C367 B.n327 VSUBS 0.012315f
C368 B.n328 VSUBS 0.012315f
C369 B.n329 VSUBS 0.012315f
C370 B.n330 VSUBS 0.012315f
C371 B.n331 VSUBS 0.012315f
C372 B.n332 VSUBS 0.012315f
C373 B.n333 VSUBS 0.012315f
C374 B.n334 VSUBS 0.012315f
C375 B.n335 VSUBS 0.012315f
C376 B.n336 VSUBS 0.012315f
C377 B.n337 VSUBS 0.012315f
C378 B.n338 VSUBS 0.012315f
C379 B.n339 VSUBS 0.012315f
C380 B.n340 VSUBS 0.012315f
C381 B.n341 VSUBS 0.012315f
C382 B.n342 VSUBS 0.012315f
C383 B.n343 VSUBS 0.012315f
C384 B.n344 VSUBS 0.012315f
C385 B.n345 VSUBS 0.012315f
C386 B.n346 VSUBS 0.012315f
C387 B.n347 VSUBS 0.012315f
C388 B.n348 VSUBS 0.012315f
C389 B.n349 VSUBS 0.012315f
C390 B.n350 VSUBS 0.012315f
C391 B.n351 VSUBS 0.012315f
C392 B.n352 VSUBS 0.012315f
C393 B.n353 VSUBS 0.012315f
C394 B.n354 VSUBS 0.012315f
C395 B.n355 VSUBS 0.012315f
C396 B.n356 VSUBS 0.012315f
C397 B.n357 VSUBS 0.012315f
C398 B.n358 VSUBS 0.012315f
C399 B.n359 VSUBS 0.012315f
C400 B.n360 VSUBS 0.012315f
C401 B.n361 VSUBS 0.012315f
C402 B.n362 VSUBS 0.012315f
C403 B.n363 VSUBS 0.012315f
C404 B.n364 VSUBS 0.012315f
C405 B.n365 VSUBS 0.012315f
C406 B.n366 VSUBS 0.012315f
C407 B.n367 VSUBS 0.012315f
C408 B.n368 VSUBS 0.012315f
C409 B.n369 VSUBS 0.012315f
C410 B.n370 VSUBS 0.012315f
C411 B.n371 VSUBS 0.012315f
C412 B.n372 VSUBS 0.012315f
C413 B.n373 VSUBS 0.012315f
C414 B.n374 VSUBS 0.012315f
C415 B.n375 VSUBS 0.012315f
C416 B.n376 VSUBS 0.012315f
C417 B.n377 VSUBS 0.012315f
C418 B.n378 VSUBS 0.012315f
C419 B.n379 VSUBS 0.012315f
C420 B.n380 VSUBS 0.012315f
C421 B.n381 VSUBS 0.012315f
C422 B.n382 VSUBS 0.012315f
C423 B.n383 VSUBS 0.012315f
C424 B.n384 VSUBS 0.012315f
C425 B.n385 VSUBS 0.012315f
C426 B.n386 VSUBS 0.012315f
C427 B.n387 VSUBS 0.012315f
C428 B.n388 VSUBS 0.012315f
C429 B.n389 VSUBS 0.012315f
C430 B.n390 VSUBS 0.012315f
C431 B.n391 VSUBS 0.012315f
C432 B.n392 VSUBS 0.012315f
C433 B.n393 VSUBS 0.012315f
C434 B.n394 VSUBS 0.012315f
C435 B.n395 VSUBS 0.012315f
C436 B.n396 VSUBS 0.012315f
C437 B.n397 VSUBS 0.012315f
C438 B.n398 VSUBS 0.012315f
C439 B.n399 VSUBS 0.012315f
C440 B.n400 VSUBS 0.012315f
C441 B.n401 VSUBS 0.012315f
C442 B.n402 VSUBS 0.012315f
C443 B.n403 VSUBS 0.012315f
C444 B.n404 VSUBS 0.012315f
C445 B.n405 VSUBS 0.012315f
C446 B.n406 VSUBS 0.012315f
C447 B.n407 VSUBS 0.012315f
C448 B.n408 VSUBS 0.012315f
C449 B.n409 VSUBS 0.012315f
C450 B.n410 VSUBS 0.012315f
C451 B.n411 VSUBS 0.012315f
C452 B.n412 VSUBS 0.012315f
C453 B.n413 VSUBS 0.012315f
C454 B.n414 VSUBS 0.012315f
C455 B.n415 VSUBS 0.012315f
C456 B.n416 VSUBS 0.012315f
C457 B.n417 VSUBS 0.012315f
C458 B.n418 VSUBS 0.012315f
C459 B.n419 VSUBS 0.012315f
C460 B.n420 VSUBS 0.012315f
C461 B.n421 VSUBS 0.012315f
C462 B.n422 VSUBS 0.012315f
C463 B.n423 VSUBS 0.012315f
C464 B.n424 VSUBS 0.012315f
C465 B.n425 VSUBS 0.012315f
C466 B.n426 VSUBS 0.012315f
C467 B.n427 VSUBS 0.012315f
C468 B.n428 VSUBS 0.012315f
C469 B.n429 VSUBS 0.012315f
C470 B.n430 VSUBS 0.012315f
C471 B.n431 VSUBS 0.012315f
C472 B.n432 VSUBS 0.012315f
C473 B.n433 VSUBS 0.012315f
C474 B.n434 VSUBS 0.012315f
C475 B.n435 VSUBS 0.012315f
C476 B.n436 VSUBS 0.012315f
C477 B.n437 VSUBS 0.012315f
C478 B.n438 VSUBS 0.012315f
C479 B.n439 VSUBS 0.012315f
C480 B.n440 VSUBS 0.012315f
C481 B.n441 VSUBS 0.012315f
C482 B.n442 VSUBS 0.012315f
C483 B.n443 VSUBS 0.012315f
C484 B.n444 VSUBS 0.012315f
C485 B.n445 VSUBS 0.012315f
C486 B.n446 VSUBS 0.012315f
C487 B.n447 VSUBS 0.012315f
C488 B.n448 VSUBS 0.012315f
C489 B.n449 VSUBS 0.012315f
C490 B.n450 VSUBS 0.012315f
C491 B.n451 VSUBS 0.012315f
C492 B.n452 VSUBS 0.012315f
C493 B.n453 VSUBS 0.012315f
C494 B.n454 VSUBS 0.012315f
C495 B.n455 VSUBS 0.012315f
C496 B.n456 VSUBS 0.012315f
C497 B.n457 VSUBS 0.012315f
C498 B.n458 VSUBS 0.012315f
C499 B.n459 VSUBS 0.027236f
C500 B.n460 VSUBS 0.027236f
C501 B.n461 VSUBS 0.028542f
C502 B.n462 VSUBS 0.012315f
C503 B.n463 VSUBS 0.012315f
C504 B.n464 VSUBS 0.012315f
C505 B.n465 VSUBS 0.012315f
C506 B.n466 VSUBS 0.012315f
C507 B.n467 VSUBS 0.012315f
C508 B.n468 VSUBS 0.012315f
C509 B.n469 VSUBS 0.012315f
C510 B.n470 VSUBS 0.012315f
C511 B.n471 VSUBS 0.012315f
C512 B.n472 VSUBS 0.012315f
C513 B.n473 VSUBS 0.012315f
C514 B.n474 VSUBS 0.01159f
C515 B.n475 VSUBS 0.012315f
C516 B.n476 VSUBS 0.012315f
C517 B.n477 VSUBS 0.012315f
C518 B.n478 VSUBS 0.012315f
C519 B.n479 VSUBS 0.012315f
C520 B.n480 VSUBS 0.012315f
C521 B.n481 VSUBS 0.012315f
C522 B.n482 VSUBS 0.012315f
C523 B.n483 VSUBS 0.012315f
C524 B.n484 VSUBS 0.012315f
C525 B.n485 VSUBS 0.012315f
C526 B.n486 VSUBS 0.012315f
C527 B.n487 VSUBS 0.012315f
C528 B.n488 VSUBS 0.012315f
C529 B.n489 VSUBS 0.012315f
C530 B.n490 VSUBS 0.006882f
C531 B.n491 VSUBS 0.028532f
C532 B.n492 VSUBS 0.01159f
C533 B.n493 VSUBS 0.012315f
C534 B.n494 VSUBS 0.012315f
C535 B.n495 VSUBS 0.012315f
C536 B.n496 VSUBS 0.012315f
C537 B.n497 VSUBS 0.012315f
C538 B.n498 VSUBS 0.012315f
C539 B.n499 VSUBS 0.012315f
C540 B.n500 VSUBS 0.012315f
C541 B.n501 VSUBS 0.012315f
C542 B.n502 VSUBS 0.012315f
C543 B.n503 VSUBS 0.012315f
C544 B.n504 VSUBS 0.012315f
C545 B.n505 VSUBS 0.028542f
C546 B.n506 VSUBS 0.028542f
C547 B.n507 VSUBS 0.027236f
C548 B.n508 VSUBS 0.012315f
C549 B.n509 VSUBS 0.012315f
C550 B.n510 VSUBS 0.012315f
C551 B.n511 VSUBS 0.012315f
C552 B.n512 VSUBS 0.012315f
C553 B.n513 VSUBS 0.012315f
C554 B.n514 VSUBS 0.012315f
C555 B.n515 VSUBS 0.012315f
C556 B.n516 VSUBS 0.012315f
C557 B.n517 VSUBS 0.012315f
C558 B.n518 VSUBS 0.012315f
C559 B.n519 VSUBS 0.012315f
C560 B.n520 VSUBS 0.012315f
C561 B.n521 VSUBS 0.012315f
C562 B.n522 VSUBS 0.012315f
C563 B.n523 VSUBS 0.012315f
C564 B.n524 VSUBS 0.012315f
C565 B.n525 VSUBS 0.012315f
C566 B.n526 VSUBS 0.012315f
C567 B.n527 VSUBS 0.012315f
C568 B.n528 VSUBS 0.012315f
C569 B.n529 VSUBS 0.012315f
C570 B.n530 VSUBS 0.012315f
C571 B.n531 VSUBS 0.012315f
C572 B.n532 VSUBS 0.012315f
C573 B.n533 VSUBS 0.012315f
C574 B.n534 VSUBS 0.012315f
C575 B.n535 VSUBS 0.012315f
C576 B.n536 VSUBS 0.012315f
C577 B.n537 VSUBS 0.012315f
C578 B.n538 VSUBS 0.012315f
C579 B.n539 VSUBS 0.012315f
C580 B.n540 VSUBS 0.012315f
C581 B.n541 VSUBS 0.012315f
C582 B.n542 VSUBS 0.012315f
C583 B.n543 VSUBS 0.012315f
C584 B.n544 VSUBS 0.012315f
C585 B.n545 VSUBS 0.012315f
C586 B.n546 VSUBS 0.012315f
C587 B.n547 VSUBS 0.012315f
C588 B.n548 VSUBS 0.012315f
C589 B.n549 VSUBS 0.012315f
C590 B.n550 VSUBS 0.012315f
C591 B.n551 VSUBS 0.012315f
C592 B.n552 VSUBS 0.012315f
C593 B.n553 VSUBS 0.012315f
C594 B.n554 VSUBS 0.012315f
C595 B.n555 VSUBS 0.012315f
C596 B.n556 VSUBS 0.012315f
C597 B.n557 VSUBS 0.012315f
C598 B.n558 VSUBS 0.012315f
C599 B.n559 VSUBS 0.012315f
C600 B.n560 VSUBS 0.012315f
C601 B.n561 VSUBS 0.012315f
C602 B.n562 VSUBS 0.012315f
C603 B.n563 VSUBS 0.012315f
C604 B.n564 VSUBS 0.012315f
C605 B.n565 VSUBS 0.012315f
C606 B.n566 VSUBS 0.012315f
C607 B.n567 VSUBS 0.012315f
C608 B.n568 VSUBS 0.012315f
C609 B.n569 VSUBS 0.012315f
C610 B.n570 VSUBS 0.012315f
C611 B.n571 VSUBS 0.012315f
C612 B.n572 VSUBS 0.012315f
C613 B.n573 VSUBS 0.012315f
C614 B.n574 VSUBS 0.012315f
C615 B.n575 VSUBS 0.012315f
C616 B.n576 VSUBS 0.012315f
C617 B.n577 VSUBS 0.012315f
C618 B.n578 VSUBS 0.012315f
C619 B.n579 VSUBS 0.012315f
C620 B.n580 VSUBS 0.012315f
C621 B.n581 VSUBS 0.012315f
C622 B.n582 VSUBS 0.012315f
C623 B.n583 VSUBS 0.012315f
C624 B.n584 VSUBS 0.012315f
C625 B.n585 VSUBS 0.012315f
C626 B.n586 VSUBS 0.012315f
C627 B.n587 VSUBS 0.012315f
C628 B.n588 VSUBS 0.012315f
C629 B.n589 VSUBS 0.012315f
C630 B.n590 VSUBS 0.012315f
C631 B.n591 VSUBS 0.01607f
C632 B.n592 VSUBS 0.017119f
C633 B.n593 VSUBS 0.034042f
C634 VDD2.t2 VSUBS 0.107493f
C635 VDD2.t0 VSUBS 0.019434f
C636 VDD2.t3 VSUBS 0.019434f
C637 VDD2.n0 VSUBS 0.064755f
C638 VDD2.n1 VSUBS 2.11332f
C639 VDD2.t5 VSUBS 0.105136f
C640 VDD2.n2 VSUBS 1.7032f
C641 VDD2.t1 VSUBS 0.019434f
C642 VDD2.t4 VSUBS 0.019434f
C643 VDD2.n3 VSUBS 0.06475f
C644 VN.n0 VSUBS 0.099673f
C645 VN.t2 VSUBS 0.559842f
C646 VN.n1 VSUBS 0.100547f
C647 VN.n2 VSUBS 0.05299f
C648 VN.n3 VSUBS 0.098759f
C649 VN.t3 VSUBS 1.12958f
C650 VN.n4 VSUBS 0.631022f
C651 VN.t5 VSUBS 0.559842f
C652 VN.n5 VSUBS 0.490348f
C653 VN.n6 VSUBS 0.07438f
C654 VN.n7 VSUBS 0.696304f
C655 VN.n8 VSUBS 0.05299f
C656 VN.n9 VSUBS 0.05299f
C657 VN.n10 VSUBS 0.098759f
C658 VN.n11 VSUBS 0.091121f
C659 VN.n12 VSUBS 0.061813f
C660 VN.n13 VSUBS 0.05299f
C661 VN.n14 VSUBS 0.05299f
C662 VN.n15 VSUBS 0.05299f
C663 VN.n16 VSUBS 0.098759f
C664 VN.n17 VSUBS 0.092909f
C665 VN.n18 VSUBS 0.531266f
C666 VN.n19 VSUBS 0.162424f
C667 VN.n20 VSUBS 0.099673f
C668 VN.t0 VSUBS 0.559842f
C669 VN.n21 VSUBS 0.100547f
C670 VN.n22 VSUBS 0.05299f
C671 VN.n23 VSUBS 0.098759f
C672 VN.t1 VSUBS 1.12958f
C673 VN.n24 VSUBS 0.631022f
C674 VN.t4 VSUBS 0.559842f
C675 VN.n25 VSUBS 0.490348f
C676 VN.n26 VSUBS 0.07438f
C677 VN.n27 VSUBS 0.696304f
C678 VN.n28 VSUBS 0.05299f
C679 VN.n29 VSUBS 0.05299f
C680 VN.n30 VSUBS 0.098759f
C681 VN.n31 VSUBS 0.091121f
C682 VN.n32 VSUBS 0.061813f
C683 VN.n33 VSUBS 0.05299f
C684 VN.n34 VSUBS 0.05299f
C685 VN.n35 VSUBS 0.05299f
C686 VN.n36 VSUBS 0.098759f
C687 VN.n37 VSUBS 0.092909f
C688 VN.n38 VSUBS 0.531266f
C689 VN.n39 VSUBS 2.72393f
C690 VDD1.t5 VSUBS 0.103973f
C691 VDD1.t4 VSUBS 0.10383f
C692 VDD1.t1 VSUBS 0.018772f
C693 VDD1.t0 VSUBS 0.018772f
C694 VDD1.n0 VSUBS 0.062549f
C695 VDD1.n1 VSUBS 2.14578f
C696 VDD1.t3 VSUBS 0.018772f
C697 VDD1.t2 VSUBS 0.018772f
C698 VDD1.n2 VSUBS 0.061497f
C699 VDD1.n3 VSUBS 1.69526f
C700 VTAIL.t3 VSUBS 0.041517f
C701 VTAIL.t2 VSUBS 0.041517f
C702 VTAIL.n0 VSUBS 0.118166f
C703 VTAIL.n1 VSUBS 0.742738f
C704 VTAIL.t11 VSUBS 0.207709f
C705 VTAIL.n2 VSUBS 1.10899f
C706 VTAIL.t7 VSUBS 0.041517f
C707 VTAIL.t10 VSUBS 0.041517f
C708 VTAIL.n3 VSUBS 0.118166f
C709 VTAIL.n4 VSUBS 2.41549f
C710 VTAIL.t5 VSUBS 0.041517f
C711 VTAIL.t0 VSUBS 0.041517f
C712 VTAIL.n5 VSUBS 0.118165f
C713 VTAIL.n6 VSUBS 2.41549f
C714 VTAIL.t1 VSUBS 0.207709f
C715 VTAIL.n7 VSUBS 1.10899f
C716 VTAIL.t8 VSUBS 0.041517f
C717 VTAIL.t6 VSUBS 0.041517f
C718 VTAIL.n8 VSUBS 0.118165f
C719 VTAIL.n9 VSUBS 1.08531f
C720 VTAIL.t9 VSUBS 0.207709f
C721 VTAIL.n10 VSUBS 1.97239f
C722 VTAIL.t4 VSUBS 0.207709f
C723 VTAIL.n11 VSUBS 1.84818f
C724 VP.n0 VSUBS 0.11719f
C725 VP.t5 VSUBS 0.658229f
C726 VP.n1 VSUBS 0.118217f
C727 VP.n2 VSUBS 0.062302f
C728 VP.n3 VSUBS 0.116115f
C729 VP.n4 VSUBS 0.062302f
C730 VP.t4 VSUBS 0.658229f
C731 VP.n5 VSUBS 0.116115f
C732 VP.n6 VSUBS 0.062302f
C733 VP.n7 VSUBS 0.116115f
C734 VP.n8 VSUBS 0.11719f
C735 VP.t3 VSUBS 0.658229f
C736 VP.n9 VSUBS 0.118217f
C737 VP.n10 VSUBS 0.062302f
C738 VP.n11 VSUBS 0.116115f
C739 VP.t0 VSUBS 1.32809f
C740 VP.n12 VSUBS 0.74192f
C741 VP.t2 VSUBS 0.658229f
C742 VP.n13 VSUBS 0.576522f
C743 VP.n14 VSUBS 0.087452f
C744 VP.n15 VSUBS 0.818675f
C745 VP.n16 VSUBS 0.062302f
C746 VP.n17 VSUBS 0.062302f
C747 VP.n18 VSUBS 0.116115f
C748 VP.n19 VSUBS 0.107134f
C749 VP.n20 VSUBS 0.072676f
C750 VP.n21 VSUBS 0.062302f
C751 VP.n22 VSUBS 0.062302f
C752 VP.n23 VSUBS 0.062302f
C753 VP.n24 VSUBS 0.116115f
C754 VP.n25 VSUBS 0.109236f
C755 VP.n26 VSUBS 0.62463f
C756 VP.n27 VSUBS 3.18516f
C757 VP.n28 VSUBS 3.23412f
C758 VP.t1 VSUBS 0.658229f
C759 VP.n29 VSUBS 0.62463f
C760 VP.n30 VSUBS 0.109236f
C761 VP.n31 VSUBS 0.11719f
C762 VP.n32 VSUBS 0.062302f
C763 VP.n33 VSUBS 0.062302f
C764 VP.n34 VSUBS 0.118217f
C765 VP.n35 VSUBS 0.072676f
C766 VP.n36 VSUBS 0.107134f
C767 VP.n37 VSUBS 0.062302f
C768 VP.n38 VSUBS 0.062302f
C769 VP.n39 VSUBS 0.062302f
C770 VP.n40 VSUBS 0.116115f
C771 VP.n41 VSUBS 0.087452f
C772 VP.n42 VSUBS 0.35162f
C773 VP.n43 VSUBS 0.087452f
C774 VP.n44 VSUBS 0.062302f
C775 VP.n45 VSUBS 0.062302f
C776 VP.n46 VSUBS 0.062302f
C777 VP.n47 VSUBS 0.116115f
C778 VP.n48 VSUBS 0.107134f
C779 VP.n49 VSUBS 0.072676f
C780 VP.n50 VSUBS 0.062302f
C781 VP.n51 VSUBS 0.062302f
C782 VP.n52 VSUBS 0.062302f
C783 VP.n53 VSUBS 0.116115f
C784 VP.n54 VSUBS 0.109236f
C785 VP.n55 VSUBS 0.62463f
C786 VP.n56 VSUBS 0.190968f
.ends

