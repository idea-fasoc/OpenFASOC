* NGSPICE file created from diff_pair_sample_0351.ext - technology: sky130A

.subckt diff_pair_sample_0351 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=1.09395 pd=6.96 as=1.09395 ps=6.96 w=6.63 l=0.96
X1 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=2.5857 pd=14.04 as=0 ps=0 w=6.63 l=0.96
X2 VDD1.t6 VP.t1 VTAIL.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=1.09395 pd=6.96 as=1.09395 ps=6.96 w=6.63 l=0.96
X3 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=2.5857 pd=14.04 as=0 ps=0 w=6.63 l=0.96
X4 VDD2.t7 VN.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.09395 pd=6.96 as=2.5857 ps=14.04 w=6.63 l=0.96
X5 VTAIL.t2 VN.t1 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.09395 pd=6.96 as=1.09395 ps=6.96 w=6.63 l=0.96
X6 VDD2.t5 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.09395 pd=6.96 as=1.09395 ps=6.96 w=6.63 l=0.96
X7 VTAIL.t1 VN.t3 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5857 pd=14.04 as=1.09395 ps=6.96 w=6.63 l=0.96
X8 VTAIL.t11 VP.t2 VDD1.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=2.5857 pd=14.04 as=1.09395 ps=6.96 w=6.63 l=0.96
X9 VTAIL.t9 VP.t3 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5857 pd=14.04 as=1.09395 ps=6.96 w=6.63 l=0.96
X10 VDD1.t3 VP.t4 VTAIL.t15 B.t4 sky130_fd_pr__nfet_01v8 ad=1.09395 pd=6.96 as=2.5857 ps=14.04 w=6.63 l=0.96
X11 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=2.5857 pd=14.04 as=0 ps=0 w=6.63 l=0.96
X12 VDD2.t3 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.09395 pd=6.96 as=2.5857 ps=14.04 w=6.63 l=0.96
X13 VTAIL.t7 VN.t5 VDD2.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=2.5857 pd=14.04 as=1.09395 ps=6.96 w=6.63 l=0.96
X14 VDD1.t2 VP.t5 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=1.09395 pd=6.96 as=2.5857 ps=14.04 w=6.63 l=0.96
X15 VTAIL.t13 VP.t6 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=1.09395 pd=6.96 as=1.09395 ps=6.96 w=6.63 l=0.96
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.5857 pd=14.04 as=0 ps=0 w=6.63 l=0.96
X17 VDD2.t1 VN.t6 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.09395 pd=6.96 as=1.09395 ps=6.96 w=6.63 l=0.96
X18 VTAIL.t5 VN.t7 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=1.09395 pd=6.96 as=1.09395 ps=6.96 w=6.63 l=0.96
X19 VTAIL.t12 VP.t7 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.09395 pd=6.96 as=1.09395 ps=6.96 w=6.63 l=0.96
R0 VP.n5 VP.t3 222.43
R1 VP.n17 VP.t2 207.612
R2 VP.n27 VP.t5 207.612
R3 VP.n14 VP.t4 207.612
R4 VP.n19 VP.t1 166.441
R5 VP.n25 VP.t7 166.441
R6 VP.n12 VP.t6 166.441
R7 VP.n6 VP.t0 166.441
R8 VP.n8 VP.n7 161.3
R9 VP.n9 VP.n4 161.3
R10 VP.n11 VP.n10 161.3
R11 VP.n13 VP.n3 161.3
R12 VP.n26 VP.n0 161.3
R13 VP.n24 VP.n23 161.3
R14 VP.n22 VP.n1 161.3
R15 VP.n21 VP.n20 161.3
R16 VP.n18 VP.n2 161.3
R17 VP.n15 VP.n14 80.6037
R18 VP.n28 VP.n27 80.6037
R19 VP.n17 VP.n16 80.6037
R20 VP.n18 VP.n17 54.3172
R21 VP.n27 VP.n26 54.3172
R22 VP.n14 VP.n13 54.3172
R23 VP.n6 VP.n5 46.9212
R24 VP.n8 VP.n5 44.1937
R25 VP.n20 VP.n1 40.4934
R26 VP.n24 VP.n1 40.4934
R27 VP.n11 VP.n4 40.4934
R28 VP.n7 VP.n4 40.4934
R29 VP.n16 VP.n15 39.312
R30 VP.n19 VP.n18 17.3721
R31 VP.n26 VP.n25 17.3721
R32 VP.n13 VP.n12 17.3721
R33 VP.n20 VP.n19 7.09593
R34 VP.n25 VP.n24 7.09593
R35 VP.n12 VP.n11 7.09593
R36 VP.n7 VP.n6 7.09593
R37 VP.n15 VP.n3 0.285035
R38 VP.n16 VP.n2 0.285035
R39 VP.n28 VP.n0 0.285035
R40 VP.n9 VP.n8 0.189894
R41 VP.n10 VP.n9 0.189894
R42 VP.n10 VP.n3 0.189894
R43 VP.n21 VP.n2 0.189894
R44 VP.n22 VP.n21 0.189894
R45 VP.n23 VP.n22 0.189894
R46 VP.n23 VP.n0 0.189894
R47 VP VP.n28 0.146778
R48 VTAIL.n290 VTAIL.n260 289.615
R49 VTAIL.n32 VTAIL.n2 289.615
R50 VTAIL.n68 VTAIL.n38 289.615
R51 VTAIL.n106 VTAIL.n76 289.615
R52 VTAIL.n254 VTAIL.n224 289.615
R53 VTAIL.n216 VTAIL.n186 289.615
R54 VTAIL.n180 VTAIL.n150 289.615
R55 VTAIL.n142 VTAIL.n112 289.615
R56 VTAIL.n273 VTAIL.n272 185
R57 VTAIL.n275 VTAIL.n274 185
R58 VTAIL.n268 VTAIL.n267 185
R59 VTAIL.n281 VTAIL.n280 185
R60 VTAIL.n283 VTAIL.n282 185
R61 VTAIL.n264 VTAIL.n263 185
R62 VTAIL.n289 VTAIL.n288 185
R63 VTAIL.n291 VTAIL.n290 185
R64 VTAIL.n15 VTAIL.n14 185
R65 VTAIL.n17 VTAIL.n16 185
R66 VTAIL.n10 VTAIL.n9 185
R67 VTAIL.n23 VTAIL.n22 185
R68 VTAIL.n25 VTAIL.n24 185
R69 VTAIL.n6 VTAIL.n5 185
R70 VTAIL.n31 VTAIL.n30 185
R71 VTAIL.n33 VTAIL.n32 185
R72 VTAIL.n51 VTAIL.n50 185
R73 VTAIL.n53 VTAIL.n52 185
R74 VTAIL.n46 VTAIL.n45 185
R75 VTAIL.n59 VTAIL.n58 185
R76 VTAIL.n61 VTAIL.n60 185
R77 VTAIL.n42 VTAIL.n41 185
R78 VTAIL.n67 VTAIL.n66 185
R79 VTAIL.n69 VTAIL.n68 185
R80 VTAIL.n89 VTAIL.n88 185
R81 VTAIL.n91 VTAIL.n90 185
R82 VTAIL.n84 VTAIL.n83 185
R83 VTAIL.n97 VTAIL.n96 185
R84 VTAIL.n99 VTAIL.n98 185
R85 VTAIL.n80 VTAIL.n79 185
R86 VTAIL.n105 VTAIL.n104 185
R87 VTAIL.n107 VTAIL.n106 185
R88 VTAIL.n255 VTAIL.n254 185
R89 VTAIL.n253 VTAIL.n252 185
R90 VTAIL.n228 VTAIL.n227 185
R91 VTAIL.n247 VTAIL.n246 185
R92 VTAIL.n245 VTAIL.n244 185
R93 VTAIL.n232 VTAIL.n231 185
R94 VTAIL.n239 VTAIL.n238 185
R95 VTAIL.n237 VTAIL.n236 185
R96 VTAIL.n217 VTAIL.n216 185
R97 VTAIL.n215 VTAIL.n214 185
R98 VTAIL.n190 VTAIL.n189 185
R99 VTAIL.n209 VTAIL.n208 185
R100 VTAIL.n207 VTAIL.n206 185
R101 VTAIL.n194 VTAIL.n193 185
R102 VTAIL.n201 VTAIL.n200 185
R103 VTAIL.n199 VTAIL.n198 185
R104 VTAIL.n181 VTAIL.n180 185
R105 VTAIL.n179 VTAIL.n178 185
R106 VTAIL.n154 VTAIL.n153 185
R107 VTAIL.n173 VTAIL.n172 185
R108 VTAIL.n171 VTAIL.n170 185
R109 VTAIL.n158 VTAIL.n157 185
R110 VTAIL.n165 VTAIL.n164 185
R111 VTAIL.n163 VTAIL.n162 185
R112 VTAIL.n143 VTAIL.n142 185
R113 VTAIL.n141 VTAIL.n140 185
R114 VTAIL.n116 VTAIL.n115 185
R115 VTAIL.n135 VTAIL.n134 185
R116 VTAIL.n133 VTAIL.n132 185
R117 VTAIL.n120 VTAIL.n119 185
R118 VTAIL.n127 VTAIL.n126 185
R119 VTAIL.n125 VTAIL.n124 185
R120 VTAIL.n271 VTAIL.t4 147.659
R121 VTAIL.n13 VTAIL.t1 147.659
R122 VTAIL.n49 VTAIL.t14 147.659
R123 VTAIL.n87 VTAIL.t11 147.659
R124 VTAIL.n235 VTAIL.t15 147.659
R125 VTAIL.n197 VTAIL.t9 147.659
R126 VTAIL.n161 VTAIL.t0 147.659
R127 VTAIL.n123 VTAIL.t7 147.659
R128 VTAIL.n274 VTAIL.n273 104.615
R129 VTAIL.n274 VTAIL.n267 104.615
R130 VTAIL.n281 VTAIL.n267 104.615
R131 VTAIL.n282 VTAIL.n281 104.615
R132 VTAIL.n282 VTAIL.n263 104.615
R133 VTAIL.n289 VTAIL.n263 104.615
R134 VTAIL.n290 VTAIL.n289 104.615
R135 VTAIL.n16 VTAIL.n15 104.615
R136 VTAIL.n16 VTAIL.n9 104.615
R137 VTAIL.n23 VTAIL.n9 104.615
R138 VTAIL.n24 VTAIL.n23 104.615
R139 VTAIL.n24 VTAIL.n5 104.615
R140 VTAIL.n31 VTAIL.n5 104.615
R141 VTAIL.n32 VTAIL.n31 104.615
R142 VTAIL.n52 VTAIL.n51 104.615
R143 VTAIL.n52 VTAIL.n45 104.615
R144 VTAIL.n59 VTAIL.n45 104.615
R145 VTAIL.n60 VTAIL.n59 104.615
R146 VTAIL.n60 VTAIL.n41 104.615
R147 VTAIL.n67 VTAIL.n41 104.615
R148 VTAIL.n68 VTAIL.n67 104.615
R149 VTAIL.n90 VTAIL.n89 104.615
R150 VTAIL.n90 VTAIL.n83 104.615
R151 VTAIL.n97 VTAIL.n83 104.615
R152 VTAIL.n98 VTAIL.n97 104.615
R153 VTAIL.n98 VTAIL.n79 104.615
R154 VTAIL.n105 VTAIL.n79 104.615
R155 VTAIL.n106 VTAIL.n105 104.615
R156 VTAIL.n254 VTAIL.n253 104.615
R157 VTAIL.n253 VTAIL.n227 104.615
R158 VTAIL.n246 VTAIL.n227 104.615
R159 VTAIL.n246 VTAIL.n245 104.615
R160 VTAIL.n245 VTAIL.n231 104.615
R161 VTAIL.n238 VTAIL.n231 104.615
R162 VTAIL.n238 VTAIL.n237 104.615
R163 VTAIL.n216 VTAIL.n215 104.615
R164 VTAIL.n215 VTAIL.n189 104.615
R165 VTAIL.n208 VTAIL.n189 104.615
R166 VTAIL.n208 VTAIL.n207 104.615
R167 VTAIL.n207 VTAIL.n193 104.615
R168 VTAIL.n200 VTAIL.n193 104.615
R169 VTAIL.n200 VTAIL.n199 104.615
R170 VTAIL.n180 VTAIL.n179 104.615
R171 VTAIL.n179 VTAIL.n153 104.615
R172 VTAIL.n172 VTAIL.n153 104.615
R173 VTAIL.n172 VTAIL.n171 104.615
R174 VTAIL.n171 VTAIL.n157 104.615
R175 VTAIL.n164 VTAIL.n157 104.615
R176 VTAIL.n164 VTAIL.n163 104.615
R177 VTAIL.n142 VTAIL.n141 104.615
R178 VTAIL.n141 VTAIL.n115 104.615
R179 VTAIL.n134 VTAIL.n115 104.615
R180 VTAIL.n134 VTAIL.n133 104.615
R181 VTAIL.n133 VTAIL.n119 104.615
R182 VTAIL.n126 VTAIL.n119 104.615
R183 VTAIL.n126 VTAIL.n125 104.615
R184 VTAIL.n273 VTAIL.t4 52.3082
R185 VTAIL.n15 VTAIL.t1 52.3082
R186 VTAIL.n51 VTAIL.t14 52.3082
R187 VTAIL.n89 VTAIL.t11 52.3082
R188 VTAIL.n237 VTAIL.t15 52.3082
R189 VTAIL.n199 VTAIL.t9 52.3082
R190 VTAIL.n163 VTAIL.t0 52.3082
R191 VTAIL.n125 VTAIL.t7 52.3082
R192 VTAIL.n223 VTAIL.n222 47.6499
R193 VTAIL.n149 VTAIL.n148 47.6499
R194 VTAIL.n1 VTAIL.n0 47.6497
R195 VTAIL.n75 VTAIL.n74 47.6497
R196 VTAIL.n295 VTAIL.n294 30.4399
R197 VTAIL.n37 VTAIL.n36 30.4399
R198 VTAIL.n73 VTAIL.n72 30.4399
R199 VTAIL.n111 VTAIL.n110 30.4399
R200 VTAIL.n259 VTAIL.n258 30.4399
R201 VTAIL.n221 VTAIL.n220 30.4399
R202 VTAIL.n185 VTAIL.n184 30.4399
R203 VTAIL.n147 VTAIL.n146 30.4399
R204 VTAIL.n295 VTAIL.n259 19.1945
R205 VTAIL.n147 VTAIL.n111 19.1945
R206 VTAIL.n272 VTAIL.n271 15.6676
R207 VTAIL.n14 VTAIL.n13 15.6676
R208 VTAIL.n50 VTAIL.n49 15.6676
R209 VTAIL.n88 VTAIL.n87 15.6676
R210 VTAIL.n236 VTAIL.n235 15.6676
R211 VTAIL.n198 VTAIL.n197 15.6676
R212 VTAIL.n162 VTAIL.n161 15.6676
R213 VTAIL.n124 VTAIL.n123 15.6676
R214 VTAIL.n275 VTAIL.n270 12.8005
R215 VTAIL.n17 VTAIL.n12 12.8005
R216 VTAIL.n53 VTAIL.n48 12.8005
R217 VTAIL.n91 VTAIL.n86 12.8005
R218 VTAIL.n239 VTAIL.n234 12.8005
R219 VTAIL.n201 VTAIL.n196 12.8005
R220 VTAIL.n165 VTAIL.n160 12.8005
R221 VTAIL.n127 VTAIL.n122 12.8005
R222 VTAIL.n276 VTAIL.n268 12.0247
R223 VTAIL.n18 VTAIL.n10 12.0247
R224 VTAIL.n54 VTAIL.n46 12.0247
R225 VTAIL.n92 VTAIL.n84 12.0247
R226 VTAIL.n240 VTAIL.n232 12.0247
R227 VTAIL.n202 VTAIL.n194 12.0247
R228 VTAIL.n166 VTAIL.n158 12.0247
R229 VTAIL.n128 VTAIL.n120 12.0247
R230 VTAIL.n280 VTAIL.n279 11.249
R231 VTAIL.n22 VTAIL.n21 11.249
R232 VTAIL.n58 VTAIL.n57 11.249
R233 VTAIL.n96 VTAIL.n95 11.249
R234 VTAIL.n244 VTAIL.n243 11.249
R235 VTAIL.n206 VTAIL.n205 11.249
R236 VTAIL.n170 VTAIL.n169 11.249
R237 VTAIL.n132 VTAIL.n131 11.249
R238 VTAIL.n283 VTAIL.n266 10.4732
R239 VTAIL.n25 VTAIL.n8 10.4732
R240 VTAIL.n61 VTAIL.n44 10.4732
R241 VTAIL.n99 VTAIL.n82 10.4732
R242 VTAIL.n247 VTAIL.n230 10.4732
R243 VTAIL.n209 VTAIL.n192 10.4732
R244 VTAIL.n173 VTAIL.n156 10.4732
R245 VTAIL.n135 VTAIL.n118 10.4732
R246 VTAIL.n284 VTAIL.n264 9.69747
R247 VTAIL.n26 VTAIL.n6 9.69747
R248 VTAIL.n62 VTAIL.n42 9.69747
R249 VTAIL.n100 VTAIL.n80 9.69747
R250 VTAIL.n248 VTAIL.n228 9.69747
R251 VTAIL.n210 VTAIL.n190 9.69747
R252 VTAIL.n174 VTAIL.n154 9.69747
R253 VTAIL.n136 VTAIL.n116 9.69747
R254 VTAIL.n294 VTAIL.n293 9.45567
R255 VTAIL.n36 VTAIL.n35 9.45567
R256 VTAIL.n72 VTAIL.n71 9.45567
R257 VTAIL.n110 VTAIL.n109 9.45567
R258 VTAIL.n258 VTAIL.n257 9.45567
R259 VTAIL.n220 VTAIL.n219 9.45567
R260 VTAIL.n184 VTAIL.n183 9.45567
R261 VTAIL.n146 VTAIL.n145 9.45567
R262 VTAIL.n262 VTAIL.n261 9.3005
R263 VTAIL.n287 VTAIL.n286 9.3005
R264 VTAIL.n285 VTAIL.n284 9.3005
R265 VTAIL.n266 VTAIL.n265 9.3005
R266 VTAIL.n279 VTAIL.n278 9.3005
R267 VTAIL.n277 VTAIL.n276 9.3005
R268 VTAIL.n270 VTAIL.n269 9.3005
R269 VTAIL.n293 VTAIL.n292 9.3005
R270 VTAIL.n4 VTAIL.n3 9.3005
R271 VTAIL.n29 VTAIL.n28 9.3005
R272 VTAIL.n27 VTAIL.n26 9.3005
R273 VTAIL.n8 VTAIL.n7 9.3005
R274 VTAIL.n21 VTAIL.n20 9.3005
R275 VTAIL.n19 VTAIL.n18 9.3005
R276 VTAIL.n12 VTAIL.n11 9.3005
R277 VTAIL.n35 VTAIL.n34 9.3005
R278 VTAIL.n40 VTAIL.n39 9.3005
R279 VTAIL.n65 VTAIL.n64 9.3005
R280 VTAIL.n63 VTAIL.n62 9.3005
R281 VTAIL.n44 VTAIL.n43 9.3005
R282 VTAIL.n57 VTAIL.n56 9.3005
R283 VTAIL.n55 VTAIL.n54 9.3005
R284 VTAIL.n48 VTAIL.n47 9.3005
R285 VTAIL.n71 VTAIL.n70 9.3005
R286 VTAIL.n78 VTAIL.n77 9.3005
R287 VTAIL.n103 VTAIL.n102 9.3005
R288 VTAIL.n101 VTAIL.n100 9.3005
R289 VTAIL.n82 VTAIL.n81 9.3005
R290 VTAIL.n95 VTAIL.n94 9.3005
R291 VTAIL.n93 VTAIL.n92 9.3005
R292 VTAIL.n86 VTAIL.n85 9.3005
R293 VTAIL.n109 VTAIL.n108 9.3005
R294 VTAIL.n257 VTAIL.n256 9.3005
R295 VTAIL.n226 VTAIL.n225 9.3005
R296 VTAIL.n251 VTAIL.n250 9.3005
R297 VTAIL.n249 VTAIL.n248 9.3005
R298 VTAIL.n230 VTAIL.n229 9.3005
R299 VTAIL.n243 VTAIL.n242 9.3005
R300 VTAIL.n241 VTAIL.n240 9.3005
R301 VTAIL.n234 VTAIL.n233 9.3005
R302 VTAIL.n219 VTAIL.n218 9.3005
R303 VTAIL.n188 VTAIL.n187 9.3005
R304 VTAIL.n213 VTAIL.n212 9.3005
R305 VTAIL.n211 VTAIL.n210 9.3005
R306 VTAIL.n192 VTAIL.n191 9.3005
R307 VTAIL.n205 VTAIL.n204 9.3005
R308 VTAIL.n203 VTAIL.n202 9.3005
R309 VTAIL.n196 VTAIL.n195 9.3005
R310 VTAIL.n183 VTAIL.n182 9.3005
R311 VTAIL.n152 VTAIL.n151 9.3005
R312 VTAIL.n177 VTAIL.n176 9.3005
R313 VTAIL.n175 VTAIL.n174 9.3005
R314 VTAIL.n156 VTAIL.n155 9.3005
R315 VTAIL.n169 VTAIL.n168 9.3005
R316 VTAIL.n167 VTAIL.n166 9.3005
R317 VTAIL.n160 VTAIL.n159 9.3005
R318 VTAIL.n145 VTAIL.n144 9.3005
R319 VTAIL.n114 VTAIL.n113 9.3005
R320 VTAIL.n139 VTAIL.n138 9.3005
R321 VTAIL.n137 VTAIL.n136 9.3005
R322 VTAIL.n118 VTAIL.n117 9.3005
R323 VTAIL.n131 VTAIL.n130 9.3005
R324 VTAIL.n129 VTAIL.n128 9.3005
R325 VTAIL.n122 VTAIL.n121 9.3005
R326 VTAIL.n288 VTAIL.n287 8.92171
R327 VTAIL.n30 VTAIL.n29 8.92171
R328 VTAIL.n66 VTAIL.n65 8.92171
R329 VTAIL.n104 VTAIL.n103 8.92171
R330 VTAIL.n252 VTAIL.n251 8.92171
R331 VTAIL.n214 VTAIL.n213 8.92171
R332 VTAIL.n178 VTAIL.n177 8.92171
R333 VTAIL.n140 VTAIL.n139 8.92171
R334 VTAIL.n291 VTAIL.n262 8.14595
R335 VTAIL.n33 VTAIL.n4 8.14595
R336 VTAIL.n69 VTAIL.n40 8.14595
R337 VTAIL.n107 VTAIL.n78 8.14595
R338 VTAIL.n255 VTAIL.n226 8.14595
R339 VTAIL.n217 VTAIL.n188 8.14595
R340 VTAIL.n181 VTAIL.n152 8.14595
R341 VTAIL.n143 VTAIL.n114 8.14595
R342 VTAIL.n292 VTAIL.n260 7.3702
R343 VTAIL.n34 VTAIL.n2 7.3702
R344 VTAIL.n70 VTAIL.n38 7.3702
R345 VTAIL.n108 VTAIL.n76 7.3702
R346 VTAIL.n256 VTAIL.n224 7.3702
R347 VTAIL.n218 VTAIL.n186 7.3702
R348 VTAIL.n182 VTAIL.n150 7.3702
R349 VTAIL.n144 VTAIL.n112 7.3702
R350 VTAIL.n294 VTAIL.n260 6.59444
R351 VTAIL.n36 VTAIL.n2 6.59444
R352 VTAIL.n72 VTAIL.n38 6.59444
R353 VTAIL.n110 VTAIL.n76 6.59444
R354 VTAIL.n258 VTAIL.n224 6.59444
R355 VTAIL.n220 VTAIL.n186 6.59444
R356 VTAIL.n184 VTAIL.n150 6.59444
R357 VTAIL.n146 VTAIL.n112 6.59444
R358 VTAIL.n292 VTAIL.n291 5.81868
R359 VTAIL.n34 VTAIL.n33 5.81868
R360 VTAIL.n70 VTAIL.n69 5.81868
R361 VTAIL.n108 VTAIL.n107 5.81868
R362 VTAIL.n256 VTAIL.n255 5.81868
R363 VTAIL.n218 VTAIL.n217 5.81868
R364 VTAIL.n182 VTAIL.n181 5.81868
R365 VTAIL.n144 VTAIL.n143 5.81868
R366 VTAIL.n288 VTAIL.n262 5.04292
R367 VTAIL.n30 VTAIL.n4 5.04292
R368 VTAIL.n66 VTAIL.n40 5.04292
R369 VTAIL.n104 VTAIL.n78 5.04292
R370 VTAIL.n252 VTAIL.n226 5.04292
R371 VTAIL.n214 VTAIL.n188 5.04292
R372 VTAIL.n178 VTAIL.n152 5.04292
R373 VTAIL.n140 VTAIL.n114 5.04292
R374 VTAIL.n271 VTAIL.n269 4.38571
R375 VTAIL.n13 VTAIL.n11 4.38571
R376 VTAIL.n49 VTAIL.n47 4.38571
R377 VTAIL.n87 VTAIL.n85 4.38571
R378 VTAIL.n235 VTAIL.n233 4.38571
R379 VTAIL.n197 VTAIL.n195 4.38571
R380 VTAIL.n161 VTAIL.n159 4.38571
R381 VTAIL.n123 VTAIL.n121 4.38571
R382 VTAIL.n287 VTAIL.n264 4.26717
R383 VTAIL.n29 VTAIL.n6 4.26717
R384 VTAIL.n65 VTAIL.n42 4.26717
R385 VTAIL.n103 VTAIL.n80 4.26717
R386 VTAIL.n251 VTAIL.n228 4.26717
R387 VTAIL.n213 VTAIL.n190 4.26717
R388 VTAIL.n177 VTAIL.n154 4.26717
R389 VTAIL.n139 VTAIL.n116 4.26717
R390 VTAIL.n284 VTAIL.n283 3.49141
R391 VTAIL.n26 VTAIL.n25 3.49141
R392 VTAIL.n62 VTAIL.n61 3.49141
R393 VTAIL.n100 VTAIL.n99 3.49141
R394 VTAIL.n248 VTAIL.n247 3.49141
R395 VTAIL.n210 VTAIL.n209 3.49141
R396 VTAIL.n174 VTAIL.n173 3.49141
R397 VTAIL.n136 VTAIL.n135 3.49141
R398 VTAIL.n0 VTAIL.t3 2.98693
R399 VTAIL.n0 VTAIL.t5 2.98693
R400 VTAIL.n74 VTAIL.t8 2.98693
R401 VTAIL.n74 VTAIL.t12 2.98693
R402 VTAIL.n222 VTAIL.t10 2.98693
R403 VTAIL.n222 VTAIL.t13 2.98693
R404 VTAIL.n148 VTAIL.t6 2.98693
R405 VTAIL.n148 VTAIL.t2 2.98693
R406 VTAIL.n280 VTAIL.n266 2.71565
R407 VTAIL.n22 VTAIL.n8 2.71565
R408 VTAIL.n58 VTAIL.n44 2.71565
R409 VTAIL.n96 VTAIL.n82 2.71565
R410 VTAIL.n244 VTAIL.n230 2.71565
R411 VTAIL.n206 VTAIL.n192 2.71565
R412 VTAIL.n170 VTAIL.n156 2.71565
R413 VTAIL.n132 VTAIL.n118 2.71565
R414 VTAIL.n279 VTAIL.n268 1.93989
R415 VTAIL.n21 VTAIL.n10 1.93989
R416 VTAIL.n57 VTAIL.n46 1.93989
R417 VTAIL.n95 VTAIL.n84 1.93989
R418 VTAIL.n243 VTAIL.n232 1.93989
R419 VTAIL.n205 VTAIL.n194 1.93989
R420 VTAIL.n169 VTAIL.n158 1.93989
R421 VTAIL.n131 VTAIL.n120 1.93989
R422 VTAIL.n276 VTAIL.n275 1.16414
R423 VTAIL.n18 VTAIL.n17 1.16414
R424 VTAIL.n54 VTAIL.n53 1.16414
R425 VTAIL.n92 VTAIL.n91 1.16414
R426 VTAIL.n240 VTAIL.n239 1.16414
R427 VTAIL.n202 VTAIL.n201 1.16414
R428 VTAIL.n166 VTAIL.n165 1.16414
R429 VTAIL.n128 VTAIL.n127 1.16414
R430 VTAIL.n149 VTAIL.n147 1.11257
R431 VTAIL.n185 VTAIL.n149 1.11257
R432 VTAIL.n223 VTAIL.n221 1.11257
R433 VTAIL.n259 VTAIL.n223 1.11257
R434 VTAIL.n111 VTAIL.n75 1.11257
R435 VTAIL.n75 VTAIL.n73 1.11257
R436 VTAIL.n37 VTAIL.n1 1.11257
R437 VTAIL VTAIL.n295 1.05438
R438 VTAIL.n221 VTAIL.n185 0.470328
R439 VTAIL.n73 VTAIL.n37 0.470328
R440 VTAIL.n272 VTAIL.n270 0.388379
R441 VTAIL.n14 VTAIL.n12 0.388379
R442 VTAIL.n50 VTAIL.n48 0.388379
R443 VTAIL.n88 VTAIL.n86 0.388379
R444 VTAIL.n236 VTAIL.n234 0.388379
R445 VTAIL.n198 VTAIL.n196 0.388379
R446 VTAIL.n162 VTAIL.n160 0.388379
R447 VTAIL.n124 VTAIL.n122 0.388379
R448 VTAIL.n277 VTAIL.n269 0.155672
R449 VTAIL.n278 VTAIL.n277 0.155672
R450 VTAIL.n278 VTAIL.n265 0.155672
R451 VTAIL.n285 VTAIL.n265 0.155672
R452 VTAIL.n286 VTAIL.n285 0.155672
R453 VTAIL.n286 VTAIL.n261 0.155672
R454 VTAIL.n293 VTAIL.n261 0.155672
R455 VTAIL.n19 VTAIL.n11 0.155672
R456 VTAIL.n20 VTAIL.n19 0.155672
R457 VTAIL.n20 VTAIL.n7 0.155672
R458 VTAIL.n27 VTAIL.n7 0.155672
R459 VTAIL.n28 VTAIL.n27 0.155672
R460 VTAIL.n28 VTAIL.n3 0.155672
R461 VTAIL.n35 VTAIL.n3 0.155672
R462 VTAIL.n55 VTAIL.n47 0.155672
R463 VTAIL.n56 VTAIL.n55 0.155672
R464 VTAIL.n56 VTAIL.n43 0.155672
R465 VTAIL.n63 VTAIL.n43 0.155672
R466 VTAIL.n64 VTAIL.n63 0.155672
R467 VTAIL.n64 VTAIL.n39 0.155672
R468 VTAIL.n71 VTAIL.n39 0.155672
R469 VTAIL.n93 VTAIL.n85 0.155672
R470 VTAIL.n94 VTAIL.n93 0.155672
R471 VTAIL.n94 VTAIL.n81 0.155672
R472 VTAIL.n101 VTAIL.n81 0.155672
R473 VTAIL.n102 VTAIL.n101 0.155672
R474 VTAIL.n102 VTAIL.n77 0.155672
R475 VTAIL.n109 VTAIL.n77 0.155672
R476 VTAIL.n257 VTAIL.n225 0.155672
R477 VTAIL.n250 VTAIL.n225 0.155672
R478 VTAIL.n250 VTAIL.n249 0.155672
R479 VTAIL.n249 VTAIL.n229 0.155672
R480 VTAIL.n242 VTAIL.n229 0.155672
R481 VTAIL.n242 VTAIL.n241 0.155672
R482 VTAIL.n241 VTAIL.n233 0.155672
R483 VTAIL.n219 VTAIL.n187 0.155672
R484 VTAIL.n212 VTAIL.n187 0.155672
R485 VTAIL.n212 VTAIL.n211 0.155672
R486 VTAIL.n211 VTAIL.n191 0.155672
R487 VTAIL.n204 VTAIL.n191 0.155672
R488 VTAIL.n204 VTAIL.n203 0.155672
R489 VTAIL.n203 VTAIL.n195 0.155672
R490 VTAIL.n183 VTAIL.n151 0.155672
R491 VTAIL.n176 VTAIL.n151 0.155672
R492 VTAIL.n176 VTAIL.n175 0.155672
R493 VTAIL.n175 VTAIL.n155 0.155672
R494 VTAIL.n168 VTAIL.n155 0.155672
R495 VTAIL.n168 VTAIL.n167 0.155672
R496 VTAIL.n167 VTAIL.n159 0.155672
R497 VTAIL.n145 VTAIL.n113 0.155672
R498 VTAIL.n138 VTAIL.n113 0.155672
R499 VTAIL.n138 VTAIL.n137 0.155672
R500 VTAIL.n137 VTAIL.n117 0.155672
R501 VTAIL.n130 VTAIL.n117 0.155672
R502 VTAIL.n130 VTAIL.n129 0.155672
R503 VTAIL.n129 VTAIL.n121 0.155672
R504 VTAIL VTAIL.n1 0.0586897
R505 VDD1 VDD1.n0 64.9429
R506 VDD1.n3 VDD1.n2 64.8292
R507 VDD1.n3 VDD1.n1 64.8292
R508 VDD1.n5 VDD1.n4 64.3285
R509 VDD1.n5 VDD1.n3 35.0181
R510 VDD1.n4 VDD1.t1 2.98693
R511 VDD1.n4 VDD1.t3 2.98693
R512 VDD1.n0 VDD1.t4 2.98693
R513 VDD1.n0 VDD1.t7 2.98693
R514 VDD1.n2 VDD1.t0 2.98693
R515 VDD1.n2 VDD1.t2 2.98693
R516 VDD1.n1 VDD1.t5 2.98693
R517 VDD1.n1 VDD1.t6 2.98693
R518 VDD1 VDD1.n5 0.498345
R519 B.n532 B.n531 585
R520 B.n533 B.n532 585
R521 B.n205 B.n83 585
R522 B.n204 B.n203 585
R523 B.n202 B.n201 585
R524 B.n200 B.n199 585
R525 B.n198 B.n197 585
R526 B.n196 B.n195 585
R527 B.n194 B.n193 585
R528 B.n192 B.n191 585
R529 B.n190 B.n189 585
R530 B.n188 B.n187 585
R531 B.n186 B.n185 585
R532 B.n184 B.n183 585
R533 B.n182 B.n181 585
R534 B.n180 B.n179 585
R535 B.n178 B.n177 585
R536 B.n176 B.n175 585
R537 B.n174 B.n173 585
R538 B.n172 B.n171 585
R539 B.n170 B.n169 585
R540 B.n168 B.n167 585
R541 B.n166 B.n165 585
R542 B.n164 B.n163 585
R543 B.n162 B.n161 585
R544 B.n160 B.n159 585
R545 B.n158 B.n157 585
R546 B.n155 B.n154 585
R547 B.n153 B.n152 585
R548 B.n151 B.n150 585
R549 B.n149 B.n148 585
R550 B.n147 B.n146 585
R551 B.n145 B.n144 585
R552 B.n143 B.n142 585
R553 B.n141 B.n140 585
R554 B.n139 B.n138 585
R555 B.n137 B.n136 585
R556 B.n135 B.n134 585
R557 B.n133 B.n132 585
R558 B.n131 B.n130 585
R559 B.n129 B.n128 585
R560 B.n127 B.n126 585
R561 B.n125 B.n124 585
R562 B.n123 B.n122 585
R563 B.n121 B.n120 585
R564 B.n119 B.n118 585
R565 B.n117 B.n116 585
R566 B.n115 B.n114 585
R567 B.n113 B.n112 585
R568 B.n111 B.n110 585
R569 B.n109 B.n108 585
R570 B.n107 B.n106 585
R571 B.n105 B.n104 585
R572 B.n103 B.n102 585
R573 B.n101 B.n100 585
R574 B.n99 B.n98 585
R575 B.n97 B.n96 585
R576 B.n95 B.n94 585
R577 B.n93 B.n92 585
R578 B.n91 B.n90 585
R579 B.n53 B.n52 585
R580 B.n536 B.n535 585
R581 B.n530 B.n84 585
R582 B.n84 B.n50 585
R583 B.n529 B.n49 585
R584 B.n540 B.n49 585
R585 B.n528 B.n48 585
R586 B.n541 B.n48 585
R587 B.n527 B.n47 585
R588 B.n542 B.n47 585
R589 B.n526 B.n525 585
R590 B.n525 B.n43 585
R591 B.n524 B.n42 585
R592 B.n548 B.n42 585
R593 B.n523 B.n41 585
R594 B.n549 B.n41 585
R595 B.n522 B.n40 585
R596 B.n550 B.n40 585
R597 B.n521 B.n520 585
R598 B.n520 B.n36 585
R599 B.n519 B.n35 585
R600 B.n556 B.n35 585
R601 B.n518 B.n34 585
R602 B.n557 B.n34 585
R603 B.n517 B.n33 585
R604 B.n558 B.n33 585
R605 B.n516 B.n515 585
R606 B.n515 B.n32 585
R607 B.n514 B.n28 585
R608 B.n564 B.n28 585
R609 B.n513 B.n27 585
R610 B.n565 B.n27 585
R611 B.n512 B.n26 585
R612 B.n566 B.n26 585
R613 B.n511 B.n510 585
R614 B.n510 B.n22 585
R615 B.n509 B.n21 585
R616 B.n572 B.n21 585
R617 B.n508 B.n20 585
R618 B.n573 B.n20 585
R619 B.n507 B.n19 585
R620 B.n574 B.n19 585
R621 B.n506 B.n505 585
R622 B.n505 B.n15 585
R623 B.n504 B.n14 585
R624 B.n580 B.n14 585
R625 B.n503 B.n13 585
R626 B.n581 B.n13 585
R627 B.n502 B.n12 585
R628 B.n582 B.n12 585
R629 B.n501 B.n500 585
R630 B.n500 B.n8 585
R631 B.n499 B.n7 585
R632 B.n588 B.n7 585
R633 B.n498 B.n6 585
R634 B.n589 B.n6 585
R635 B.n497 B.n5 585
R636 B.n590 B.n5 585
R637 B.n496 B.n495 585
R638 B.n495 B.n4 585
R639 B.n494 B.n206 585
R640 B.n494 B.n493 585
R641 B.n484 B.n207 585
R642 B.n208 B.n207 585
R643 B.n486 B.n485 585
R644 B.n487 B.n486 585
R645 B.n483 B.n213 585
R646 B.n213 B.n212 585
R647 B.n482 B.n481 585
R648 B.n481 B.n480 585
R649 B.n215 B.n214 585
R650 B.n216 B.n215 585
R651 B.n473 B.n472 585
R652 B.n474 B.n473 585
R653 B.n471 B.n221 585
R654 B.n221 B.n220 585
R655 B.n470 B.n469 585
R656 B.n469 B.n468 585
R657 B.n223 B.n222 585
R658 B.n224 B.n223 585
R659 B.n461 B.n460 585
R660 B.n462 B.n461 585
R661 B.n459 B.n229 585
R662 B.n229 B.n228 585
R663 B.n458 B.n457 585
R664 B.n457 B.n456 585
R665 B.n231 B.n230 585
R666 B.n449 B.n231 585
R667 B.n448 B.n447 585
R668 B.n450 B.n448 585
R669 B.n446 B.n236 585
R670 B.n236 B.n235 585
R671 B.n445 B.n444 585
R672 B.n444 B.n443 585
R673 B.n238 B.n237 585
R674 B.n239 B.n238 585
R675 B.n436 B.n435 585
R676 B.n437 B.n436 585
R677 B.n434 B.n244 585
R678 B.n244 B.n243 585
R679 B.n433 B.n432 585
R680 B.n432 B.n431 585
R681 B.n246 B.n245 585
R682 B.n247 B.n246 585
R683 B.n424 B.n423 585
R684 B.n425 B.n424 585
R685 B.n422 B.n252 585
R686 B.n252 B.n251 585
R687 B.n421 B.n420 585
R688 B.n420 B.n419 585
R689 B.n254 B.n253 585
R690 B.n255 B.n254 585
R691 B.n415 B.n414 585
R692 B.n258 B.n257 585
R693 B.n411 B.n410 585
R694 B.n412 B.n411 585
R695 B.n409 B.n288 585
R696 B.n408 B.n407 585
R697 B.n406 B.n405 585
R698 B.n404 B.n403 585
R699 B.n402 B.n401 585
R700 B.n400 B.n399 585
R701 B.n398 B.n397 585
R702 B.n396 B.n395 585
R703 B.n394 B.n393 585
R704 B.n392 B.n391 585
R705 B.n390 B.n389 585
R706 B.n388 B.n387 585
R707 B.n386 B.n385 585
R708 B.n384 B.n383 585
R709 B.n382 B.n381 585
R710 B.n380 B.n379 585
R711 B.n378 B.n377 585
R712 B.n376 B.n375 585
R713 B.n374 B.n373 585
R714 B.n372 B.n371 585
R715 B.n370 B.n369 585
R716 B.n368 B.n367 585
R717 B.n366 B.n365 585
R718 B.n363 B.n362 585
R719 B.n361 B.n360 585
R720 B.n359 B.n358 585
R721 B.n357 B.n356 585
R722 B.n355 B.n354 585
R723 B.n353 B.n352 585
R724 B.n351 B.n350 585
R725 B.n349 B.n348 585
R726 B.n347 B.n346 585
R727 B.n345 B.n344 585
R728 B.n343 B.n342 585
R729 B.n341 B.n340 585
R730 B.n339 B.n338 585
R731 B.n337 B.n336 585
R732 B.n335 B.n334 585
R733 B.n333 B.n332 585
R734 B.n331 B.n330 585
R735 B.n329 B.n328 585
R736 B.n327 B.n326 585
R737 B.n325 B.n324 585
R738 B.n323 B.n322 585
R739 B.n321 B.n320 585
R740 B.n319 B.n318 585
R741 B.n317 B.n316 585
R742 B.n315 B.n314 585
R743 B.n313 B.n312 585
R744 B.n311 B.n310 585
R745 B.n309 B.n308 585
R746 B.n307 B.n306 585
R747 B.n305 B.n304 585
R748 B.n303 B.n302 585
R749 B.n301 B.n300 585
R750 B.n299 B.n298 585
R751 B.n297 B.n296 585
R752 B.n295 B.n294 585
R753 B.n416 B.n256 585
R754 B.n256 B.n255 585
R755 B.n418 B.n417 585
R756 B.n419 B.n418 585
R757 B.n250 B.n249 585
R758 B.n251 B.n250 585
R759 B.n427 B.n426 585
R760 B.n426 B.n425 585
R761 B.n428 B.n248 585
R762 B.n248 B.n247 585
R763 B.n430 B.n429 585
R764 B.n431 B.n430 585
R765 B.n242 B.n241 585
R766 B.n243 B.n242 585
R767 B.n439 B.n438 585
R768 B.n438 B.n437 585
R769 B.n440 B.n240 585
R770 B.n240 B.n239 585
R771 B.n442 B.n441 585
R772 B.n443 B.n442 585
R773 B.n234 B.n233 585
R774 B.n235 B.n234 585
R775 B.n452 B.n451 585
R776 B.n451 B.n450 585
R777 B.n453 B.n232 585
R778 B.n449 B.n232 585
R779 B.n455 B.n454 585
R780 B.n456 B.n455 585
R781 B.n227 B.n226 585
R782 B.n228 B.n227 585
R783 B.n464 B.n463 585
R784 B.n463 B.n462 585
R785 B.n465 B.n225 585
R786 B.n225 B.n224 585
R787 B.n467 B.n466 585
R788 B.n468 B.n467 585
R789 B.n219 B.n218 585
R790 B.n220 B.n219 585
R791 B.n476 B.n475 585
R792 B.n475 B.n474 585
R793 B.n477 B.n217 585
R794 B.n217 B.n216 585
R795 B.n479 B.n478 585
R796 B.n480 B.n479 585
R797 B.n211 B.n210 585
R798 B.n212 B.n211 585
R799 B.n489 B.n488 585
R800 B.n488 B.n487 585
R801 B.n490 B.n209 585
R802 B.n209 B.n208 585
R803 B.n492 B.n491 585
R804 B.n493 B.n492 585
R805 B.n2 B.n0 585
R806 B.n4 B.n2 585
R807 B.n3 B.n1 585
R808 B.n589 B.n3 585
R809 B.n587 B.n586 585
R810 B.n588 B.n587 585
R811 B.n585 B.n9 585
R812 B.n9 B.n8 585
R813 B.n584 B.n583 585
R814 B.n583 B.n582 585
R815 B.n11 B.n10 585
R816 B.n581 B.n11 585
R817 B.n579 B.n578 585
R818 B.n580 B.n579 585
R819 B.n577 B.n16 585
R820 B.n16 B.n15 585
R821 B.n576 B.n575 585
R822 B.n575 B.n574 585
R823 B.n18 B.n17 585
R824 B.n573 B.n18 585
R825 B.n571 B.n570 585
R826 B.n572 B.n571 585
R827 B.n569 B.n23 585
R828 B.n23 B.n22 585
R829 B.n568 B.n567 585
R830 B.n567 B.n566 585
R831 B.n25 B.n24 585
R832 B.n565 B.n25 585
R833 B.n563 B.n562 585
R834 B.n564 B.n563 585
R835 B.n561 B.n29 585
R836 B.n32 B.n29 585
R837 B.n560 B.n559 585
R838 B.n559 B.n558 585
R839 B.n31 B.n30 585
R840 B.n557 B.n31 585
R841 B.n555 B.n554 585
R842 B.n556 B.n555 585
R843 B.n553 B.n37 585
R844 B.n37 B.n36 585
R845 B.n552 B.n551 585
R846 B.n551 B.n550 585
R847 B.n39 B.n38 585
R848 B.n549 B.n39 585
R849 B.n547 B.n546 585
R850 B.n548 B.n547 585
R851 B.n545 B.n44 585
R852 B.n44 B.n43 585
R853 B.n544 B.n543 585
R854 B.n543 B.n542 585
R855 B.n46 B.n45 585
R856 B.n541 B.n46 585
R857 B.n539 B.n538 585
R858 B.n540 B.n539 585
R859 B.n537 B.n51 585
R860 B.n51 B.n50 585
R861 B.n592 B.n591 585
R862 B.n591 B.n590 585
R863 B.n414 B.n256 530.939
R864 B.n535 B.n51 530.939
R865 B.n294 B.n254 530.939
R866 B.n532 B.n84 530.939
R867 B.n291 B.t16 369.087
R868 B.n289 B.t8 369.087
R869 B.n87 B.t12 369.087
R870 B.n85 B.t19 369.087
R871 B.n533 B.n82 256.663
R872 B.n533 B.n81 256.663
R873 B.n533 B.n80 256.663
R874 B.n533 B.n79 256.663
R875 B.n533 B.n78 256.663
R876 B.n533 B.n77 256.663
R877 B.n533 B.n76 256.663
R878 B.n533 B.n75 256.663
R879 B.n533 B.n74 256.663
R880 B.n533 B.n73 256.663
R881 B.n533 B.n72 256.663
R882 B.n533 B.n71 256.663
R883 B.n533 B.n70 256.663
R884 B.n533 B.n69 256.663
R885 B.n533 B.n68 256.663
R886 B.n533 B.n67 256.663
R887 B.n533 B.n66 256.663
R888 B.n533 B.n65 256.663
R889 B.n533 B.n64 256.663
R890 B.n533 B.n63 256.663
R891 B.n533 B.n62 256.663
R892 B.n533 B.n61 256.663
R893 B.n533 B.n60 256.663
R894 B.n533 B.n59 256.663
R895 B.n533 B.n58 256.663
R896 B.n533 B.n57 256.663
R897 B.n533 B.n56 256.663
R898 B.n533 B.n55 256.663
R899 B.n533 B.n54 256.663
R900 B.n534 B.n533 256.663
R901 B.n413 B.n412 256.663
R902 B.n412 B.n259 256.663
R903 B.n412 B.n260 256.663
R904 B.n412 B.n261 256.663
R905 B.n412 B.n262 256.663
R906 B.n412 B.n263 256.663
R907 B.n412 B.n264 256.663
R908 B.n412 B.n265 256.663
R909 B.n412 B.n266 256.663
R910 B.n412 B.n267 256.663
R911 B.n412 B.n268 256.663
R912 B.n412 B.n269 256.663
R913 B.n412 B.n270 256.663
R914 B.n412 B.n271 256.663
R915 B.n412 B.n272 256.663
R916 B.n412 B.n273 256.663
R917 B.n412 B.n274 256.663
R918 B.n412 B.n275 256.663
R919 B.n412 B.n276 256.663
R920 B.n412 B.n277 256.663
R921 B.n412 B.n278 256.663
R922 B.n412 B.n279 256.663
R923 B.n412 B.n280 256.663
R924 B.n412 B.n281 256.663
R925 B.n412 B.n282 256.663
R926 B.n412 B.n283 256.663
R927 B.n412 B.n284 256.663
R928 B.n412 B.n285 256.663
R929 B.n412 B.n286 256.663
R930 B.n412 B.n287 256.663
R931 B.n291 B.t18 214.714
R932 B.n85 B.t20 214.714
R933 B.n289 B.t11 214.714
R934 B.n87 B.t14 214.714
R935 B.n292 B.t17 189.696
R936 B.n86 B.t21 189.696
R937 B.n290 B.t10 189.696
R938 B.n88 B.t15 189.696
R939 B.n418 B.n256 163.367
R940 B.n418 B.n250 163.367
R941 B.n426 B.n250 163.367
R942 B.n426 B.n248 163.367
R943 B.n430 B.n248 163.367
R944 B.n430 B.n242 163.367
R945 B.n438 B.n242 163.367
R946 B.n438 B.n240 163.367
R947 B.n442 B.n240 163.367
R948 B.n442 B.n234 163.367
R949 B.n451 B.n234 163.367
R950 B.n451 B.n232 163.367
R951 B.n455 B.n232 163.367
R952 B.n455 B.n227 163.367
R953 B.n463 B.n227 163.367
R954 B.n463 B.n225 163.367
R955 B.n467 B.n225 163.367
R956 B.n467 B.n219 163.367
R957 B.n475 B.n219 163.367
R958 B.n475 B.n217 163.367
R959 B.n479 B.n217 163.367
R960 B.n479 B.n211 163.367
R961 B.n488 B.n211 163.367
R962 B.n488 B.n209 163.367
R963 B.n492 B.n209 163.367
R964 B.n492 B.n2 163.367
R965 B.n591 B.n2 163.367
R966 B.n591 B.n3 163.367
R967 B.n587 B.n3 163.367
R968 B.n587 B.n9 163.367
R969 B.n583 B.n9 163.367
R970 B.n583 B.n11 163.367
R971 B.n579 B.n11 163.367
R972 B.n579 B.n16 163.367
R973 B.n575 B.n16 163.367
R974 B.n575 B.n18 163.367
R975 B.n571 B.n18 163.367
R976 B.n571 B.n23 163.367
R977 B.n567 B.n23 163.367
R978 B.n567 B.n25 163.367
R979 B.n563 B.n25 163.367
R980 B.n563 B.n29 163.367
R981 B.n559 B.n29 163.367
R982 B.n559 B.n31 163.367
R983 B.n555 B.n31 163.367
R984 B.n555 B.n37 163.367
R985 B.n551 B.n37 163.367
R986 B.n551 B.n39 163.367
R987 B.n547 B.n39 163.367
R988 B.n547 B.n44 163.367
R989 B.n543 B.n44 163.367
R990 B.n543 B.n46 163.367
R991 B.n539 B.n46 163.367
R992 B.n539 B.n51 163.367
R993 B.n411 B.n258 163.367
R994 B.n411 B.n288 163.367
R995 B.n407 B.n406 163.367
R996 B.n403 B.n402 163.367
R997 B.n399 B.n398 163.367
R998 B.n395 B.n394 163.367
R999 B.n391 B.n390 163.367
R1000 B.n387 B.n386 163.367
R1001 B.n383 B.n382 163.367
R1002 B.n379 B.n378 163.367
R1003 B.n375 B.n374 163.367
R1004 B.n371 B.n370 163.367
R1005 B.n367 B.n366 163.367
R1006 B.n362 B.n361 163.367
R1007 B.n358 B.n357 163.367
R1008 B.n354 B.n353 163.367
R1009 B.n350 B.n349 163.367
R1010 B.n346 B.n345 163.367
R1011 B.n342 B.n341 163.367
R1012 B.n338 B.n337 163.367
R1013 B.n334 B.n333 163.367
R1014 B.n330 B.n329 163.367
R1015 B.n326 B.n325 163.367
R1016 B.n322 B.n321 163.367
R1017 B.n318 B.n317 163.367
R1018 B.n314 B.n313 163.367
R1019 B.n310 B.n309 163.367
R1020 B.n306 B.n305 163.367
R1021 B.n302 B.n301 163.367
R1022 B.n298 B.n297 163.367
R1023 B.n420 B.n254 163.367
R1024 B.n420 B.n252 163.367
R1025 B.n424 B.n252 163.367
R1026 B.n424 B.n246 163.367
R1027 B.n432 B.n246 163.367
R1028 B.n432 B.n244 163.367
R1029 B.n436 B.n244 163.367
R1030 B.n436 B.n238 163.367
R1031 B.n444 B.n238 163.367
R1032 B.n444 B.n236 163.367
R1033 B.n448 B.n236 163.367
R1034 B.n448 B.n231 163.367
R1035 B.n457 B.n231 163.367
R1036 B.n457 B.n229 163.367
R1037 B.n461 B.n229 163.367
R1038 B.n461 B.n223 163.367
R1039 B.n469 B.n223 163.367
R1040 B.n469 B.n221 163.367
R1041 B.n473 B.n221 163.367
R1042 B.n473 B.n215 163.367
R1043 B.n481 B.n215 163.367
R1044 B.n481 B.n213 163.367
R1045 B.n486 B.n213 163.367
R1046 B.n486 B.n207 163.367
R1047 B.n494 B.n207 163.367
R1048 B.n495 B.n494 163.367
R1049 B.n495 B.n5 163.367
R1050 B.n6 B.n5 163.367
R1051 B.n7 B.n6 163.367
R1052 B.n500 B.n7 163.367
R1053 B.n500 B.n12 163.367
R1054 B.n13 B.n12 163.367
R1055 B.n14 B.n13 163.367
R1056 B.n505 B.n14 163.367
R1057 B.n505 B.n19 163.367
R1058 B.n20 B.n19 163.367
R1059 B.n21 B.n20 163.367
R1060 B.n510 B.n21 163.367
R1061 B.n510 B.n26 163.367
R1062 B.n27 B.n26 163.367
R1063 B.n28 B.n27 163.367
R1064 B.n515 B.n28 163.367
R1065 B.n515 B.n33 163.367
R1066 B.n34 B.n33 163.367
R1067 B.n35 B.n34 163.367
R1068 B.n520 B.n35 163.367
R1069 B.n520 B.n40 163.367
R1070 B.n41 B.n40 163.367
R1071 B.n42 B.n41 163.367
R1072 B.n525 B.n42 163.367
R1073 B.n525 B.n47 163.367
R1074 B.n48 B.n47 163.367
R1075 B.n49 B.n48 163.367
R1076 B.n84 B.n49 163.367
R1077 B.n90 B.n53 163.367
R1078 B.n94 B.n93 163.367
R1079 B.n98 B.n97 163.367
R1080 B.n102 B.n101 163.367
R1081 B.n106 B.n105 163.367
R1082 B.n110 B.n109 163.367
R1083 B.n114 B.n113 163.367
R1084 B.n118 B.n117 163.367
R1085 B.n122 B.n121 163.367
R1086 B.n126 B.n125 163.367
R1087 B.n130 B.n129 163.367
R1088 B.n134 B.n133 163.367
R1089 B.n138 B.n137 163.367
R1090 B.n142 B.n141 163.367
R1091 B.n146 B.n145 163.367
R1092 B.n150 B.n149 163.367
R1093 B.n154 B.n153 163.367
R1094 B.n159 B.n158 163.367
R1095 B.n163 B.n162 163.367
R1096 B.n167 B.n166 163.367
R1097 B.n171 B.n170 163.367
R1098 B.n175 B.n174 163.367
R1099 B.n179 B.n178 163.367
R1100 B.n183 B.n182 163.367
R1101 B.n187 B.n186 163.367
R1102 B.n191 B.n190 163.367
R1103 B.n195 B.n194 163.367
R1104 B.n199 B.n198 163.367
R1105 B.n203 B.n202 163.367
R1106 B.n532 B.n83 163.367
R1107 B.n412 B.n255 119.195
R1108 B.n533 B.n50 119.195
R1109 B.n414 B.n413 71.676
R1110 B.n288 B.n259 71.676
R1111 B.n406 B.n260 71.676
R1112 B.n402 B.n261 71.676
R1113 B.n398 B.n262 71.676
R1114 B.n394 B.n263 71.676
R1115 B.n390 B.n264 71.676
R1116 B.n386 B.n265 71.676
R1117 B.n382 B.n266 71.676
R1118 B.n378 B.n267 71.676
R1119 B.n374 B.n268 71.676
R1120 B.n370 B.n269 71.676
R1121 B.n366 B.n270 71.676
R1122 B.n361 B.n271 71.676
R1123 B.n357 B.n272 71.676
R1124 B.n353 B.n273 71.676
R1125 B.n349 B.n274 71.676
R1126 B.n345 B.n275 71.676
R1127 B.n341 B.n276 71.676
R1128 B.n337 B.n277 71.676
R1129 B.n333 B.n278 71.676
R1130 B.n329 B.n279 71.676
R1131 B.n325 B.n280 71.676
R1132 B.n321 B.n281 71.676
R1133 B.n317 B.n282 71.676
R1134 B.n313 B.n283 71.676
R1135 B.n309 B.n284 71.676
R1136 B.n305 B.n285 71.676
R1137 B.n301 B.n286 71.676
R1138 B.n297 B.n287 71.676
R1139 B.n535 B.n534 71.676
R1140 B.n90 B.n54 71.676
R1141 B.n94 B.n55 71.676
R1142 B.n98 B.n56 71.676
R1143 B.n102 B.n57 71.676
R1144 B.n106 B.n58 71.676
R1145 B.n110 B.n59 71.676
R1146 B.n114 B.n60 71.676
R1147 B.n118 B.n61 71.676
R1148 B.n122 B.n62 71.676
R1149 B.n126 B.n63 71.676
R1150 B.n130 B.n64 71.676
R1151 B.n134 B.n65 71.676
R1152 B.n138 B.n66 71.676
R1153 B.n142 B.n67 71.676
R1154 B.n146 B.n68 71.676
R1155 B.n150 B.n69 71.676
R1156 B.n154 B.n70 71.676
R1157 B.n159 B.n71 71.676
R1158 B.n163 B.n72 71.676
R1159 B.n167 B.n73 71.676
R1160 B.n171 B.n74 71.676
R1161 B.n175 B.n75 71.676
R1162 B.n179 B.n76 71.676
R1163 B.n183 B.n77 71.676
R1164 B.n187 B.n78 71.676
R1165 B.n191 B.n79 71.676
R1166 B.n195 B.n80 71.676
R1167 B.n199 B.n81 71.676
R1168 B.n203 B.n82 71.676
R1169 B.n83 B.n82 71.676
R1170 B.n202 B.n81 71.676
R1171 B.n198 B.n80 71.676
R1172 B.n194 B.n79 71.676
R1173 B.n190 B.n78 71.676
R1174 B.n186 B.n77 71.676
R1175 B.n182 B.n76 71.676
R1176 B.n178 B.n75 71.676
R1177 B.n174 B.n74 71.676
R1178 B.n170 B.n73 71.676
R1179 B.n166 B.n72 71.676
R1180 B.n162 B.n71 71.676
R1181 B.n158 B.n70 71.676
R1182 B.n153 B.n69 71.676
R1183 B.n149 B.n68 71.676
R1184 B.n145 B.n67 71.676
R1185 B.n141 B.n66 71.676
R1186 B.n137 B.n65 71.676
R1187 B.n133 B.n64 71.676
R1188 B.n129 B.n63 71.676
R1189 B.n125 B.n62 71.676
R1190 B.n121 B.n61 71.676
R1191 B.n117 B.n60 71.676
R1192 B.n113 B.n59 71.676
R1193 B.n109 B.n58 71.676
R1194 B.n105 B.n57 71.676
R1195 B.n101 B.n56 71.676
R1196 B.n97 B.n55 71.676
R1197 B.n93 B.n54 71.676
R1198 B.n534 B.n53 71.676
R1199 B.n413 B.n258 71.676
R1200 B.n407 B.n259 71.676
R1201 B.n403 B.n260 71.676
R1202 B.n399 B.n261 71.676
R1203 B.n395 B.n262 71.676
R1204 B.n391 B.n263 71.676
R1205 B.n387 B.n264 71.676
R1206 B.n383 B.n265 71.676
R1207 B.n379 B.n266 71.676
R1208 B.n375 B.n267 71.676
R1209 B.n371 B.n268 71.676
R1210 B.n367 B.n269 71.676
R1211 B.n362 B.n270 71.676
R1212 B.n358 B.n271 71.676
R1213 B.n354 B.n272 71.676
R1214 B.n350 B.n273 71.676
R1215 B.n346 B.n274 71.676
R1216 B.n342 B.n275 71.676
R1217 B.n338 B.n276 71.676
R1218 B.n334 B.n277 71.676
R1219 B.n330 B.n278 71.676
R1220 B.n326 B.n279 71.676
R1221 B.n322 B.n280 71.676
R1222 B.n318 B.n281 71.676
R1223 B.n314 B.n282 71.676
R1224 B.n310 B.n283 71.676
R1225 B.n306 B.n284 71.676
R1226 B.n302 B.n285 71.676
R1227 B.n298 B.n286 71.676
R1228 B.n294 B.n287 71.676
R1229 B.n419 B.n255 62.8312
R1230 B.n419 B.n251 62.8312
R1231 B.n425 B.n251 62.8312
R1232 B.n425 B.n247 62.8312
R1233 B.n431 B.n247 62.8312
R1234 B.n437 B.n243 62.8312
R1235 B.n437 B.n239 62.8312
R1236 B.n443 B.n239 62.8312
R1237 B.n443 B.n235 62.8312
R1238 B.n450 B.n235 62.8312
R1239 B.n450 B.n449 62.8312
R1240 B.n456 B.n228 62.8312
R1241 B.n462 B.n228 62.8312
R1242 B.n468 B.n224 62.8312
R1243 B.n468 B.n220 62.8312
R1244 B.n474 B.n220 62.8312
R1245 B.n480 B.n216 62.8312
R1246 B.n480 B.n212 62.8312
R1247 B.n487 B.n212 62.8312
R1248 B.n493 B.n208 62.8312
R1249 B.n493 B.n4 62.8312
R1250 B.n590 B.n4 62.8312
R1251 B.n590 B.n589 62.8312
R1252 B.n589 B.n588 62.8312
R1253 B.n588 B.n8 62.8312
R1254 B.n582 B.n581 62.8312
R1255 B.n581 B.n580 62.8312
R1256 B.n580 B.n15 62.8312
R1257 B.n574 B.n573 62.8312
R1258 B.n573 B.n572 62.8312
R1259 B.n572 B.n22 62.8312
R1260 B.n566 B.n565 62.8312
R1261 B.n565 B.n564 62.8312
R1262 B.n558 B.n32 62.8312
R1263 B.n558 B.n557 62.8312
R1264 B.n557 B.n556 62.8312
R1265 B.n556 B.n36 62.8312
R1266 B.n550 B.n36 62.8312
R1267 B.n550 B.n549 62.8312
R1268 B.n548 B.n43 62.8312
R1269 B.n542 B.n43 62.8312
R1270 B.n542 B.n541 62.8312
R1271 B.n541 B.n540 62.8312
R1272 B.n540 B.n50 62.8312
R1273 B.n293 B.n292 59.5399
R1274 B.n364 B.n290 59.5399
R1275 B.n89 B.n88 59.5399
R1276 B.n156 B.n86 59.5399
R1277 B.n462 B.t6 57.2874
R1278 B.n566 B.t5 57.2874
R1279 B.t9 B.n243 55.4394
R1280 B.n456 B.t7 55.4394
R1281 B.n564 B.t4 55.4394
R1282 B.n549 B.t13 55.4394
R1283 B.n474 B.t2 44.3516
R1284 B.n574 B.t3 44.3516
R1285 B.n537 B.n536 34.4981
R1286 B.n531 B.n530 34.4981
R1287 B.n295 B.n253 34.4981
R1288 B.n416 B.n415 34.4981
R1289 B.n487 B.t0 31.4159
R1290 B.t0 B.n208 31.4159
R1291 B.t1 B.n8 31.4159
R1292 B.n582 B.t1 31.4159
R1293 B.n292 B.n291 25.0187
R1294 B.n290 B.n289 25.0187
R1295 B.n88 B.n87 25.0187
R1296 B.n86 B.n85 25.0187
R1297 B.t2 B.n216 18.4801
R1298 B.t3 B.n15 18.4801
R1299 B B.n592 18.0485
R1300 B.n536 B.n52 10.6151
R1301 B.n91 B.n52 10.6151
R1302 B.n92 B.n91 10.6151
R1303 B.n95 B.n92 10.6151
R1304 B.n96 B.n95 10.6151
R1305 B.n99 B.n96 10.6151
R1306 B.n100 B.n99 10.6151
R1307 B.n103 B.n100 10.6151
R1308 B.n104 B.n103 10.6151
R1309 B.n107 B.n104 10.6151
R1310 B.n108 B.n107 10.6151
R1311 B.n111 B.n108 10.6151
R1312 B.n112 B.n111 10.6151
R1313 B.n115 B.n112 10.6151
R1314 B.n116 B.n115 10.6151
R1315 B.n119 B.n116 10.6151
R1316 B.n120 B.n119 10.6151
R1317 B.n123 B.n120 10.6151
R1318 B.n124 B.n123 10.6151
R1319 B.n127 B.n124 10.6151
R1320 B.n128 B.n127 10.6151
R1321 B.n131 B.n128 10.6151
R1322 B.n132 B.n131 10.6151
R1323 B.n135 B.n132 10.6151
R1324 B.n136 B.n135 10.6151
R1325 B.n140 B.n139 10.6151
R1326 B.n143 B.n140 10.6151
R1327 B.n144 B.n143 10.6151
R1328 B.n147 B.n144 10.6151
R1329 B.n148 B.n147 10.6151
R1330 B.n151 B.n148 10.6151
R1331 B.n152 B.n151 10.6151
R1332 B.n155 B.n152 10.6151
R1333 B.n160 B.n157 10.6151
R1334 B.n161 B.n160 10.6151
R1335 B.n164 B.n161 10.6151
R1336 B.n165 B.n164 10.6151
R1337 B.n168 B.n165 10.6151
R1338 B.n169 B.n168 10.6151
R1339 B.n172 B.n169 10.6151
R1340 B.n173 B.n172 10.6151
R1341 B.n176 B.n173 10.6151
R1342 B.n177 B.n176 10.6151
R1343 B.n180 B.n177 10.6151
R1344 B.n181 B.n180 10.6151
R1345 B.n184 B.n181 10.6151
R1346 B.n185 B.n184 10.6151
R1347 B.n188 B.n185 10.6151
R1348 B.n189 B.n188 10.6151
R1349 B.n192 B.n189 10.6151
R1350 B.n193 B.n192 10.6151
R1351 B.n196 B.n193 10.6151
R1352 B.n197 B.n196 10.6151
R1353 B.n200 B.n197 10.6151
R1354 B.n201 B.n200 10.6151
R1355 B.n204 B.n201 10.6151
R1356 B.n205 B.n204 10.6151
R1357 B.n531 B.n205 10.6151
R1358 B.n421 B.n253 10.6151
R1359 B.n422 B.n421 10.6151
R1360 B.n423 B.n422 10.6151
R1361 B.n423 B.n245 10.6151
R1362 B.n433 B.n245 10.6151
R1363 B.n434 B.n433 10.6151
R1364 B.n435 B.n434 10.6151
R1365 B.n435 B.n237 10.6151
R1366 B.n445 B.n237 10.6151
R1367 B.n446 B.n445 10.6151
R1368 B.n447 B.n446 10.6151
R1369 B.n447 B.n230 10.6151
R1370 B.n458 B.n230 10.6151
R1371 B.n459 B.n458 10.6151
R1372 B.n460 B.n459 10.6151
R1373 B.n460 B.n222 10.6151
R1374 B.n470 B.n222 10.6151
R1375 B.n471 B.n470 10.6151
R1376 B.n472 B.n471 10.6151
R1377 B.n472 B.n214 10.6151
R1378 B.n482 B.n214 10.6151
R1379 B.n483 B.n482 10.6151
R1380 B.n485 B.n483 10.6151
R1381 B.n485 B.n484 10.6151
R1382 B.n484 B.n206 10.6151
R1383 B.n496 B.n206 10.6151
R1384 B.n497 B.n496 10.6151
R1385 B.n498 B.n497 10.6151
R1386 B.n499 B.n498 10.6151
R1387 B.n501 B.n499 10.6151
R1388 B.n502 B.n501 10.6151
R1389 B.n503 B.n502 10.6151
R1390 B.n504 B.n503 10.6151
R1391 B.n506 B.n504 10.6151
R1392 B.n507 B.n506 10.6151
R1393 B.n508 B.n507 10.6151
R1394 B.n509 B.n508 10.6151
R1395 B.n511 B.n509 10.6151
R1396 B.n512 B.n511 10.6151
R1397 B.n513 B.n512 10.6151
R1398 B.n514 B.n513 10.6151
R1399 B.n516 B.n514 10.6151
R1400 B.n517 B.n516 10.6151
R1401 B.n518 B.n517 10.6151
R1402 B.n519 B.n518 10.6151
R1403 B.n521 B.n519 10.6151
R1404 B.n522 B.n521 10.6151
R1405 B.n523 B.n522 10.6151
R1406 B.n524 B.n523 10.6151
R1407 B.n526 B.n524 10.6151
R1408 B.n527 B.n526 10.6151
R1409 B.n528 B.n527 10.6151
R1410 B.n529 B.n528 10.6151
R1411 B.n530 B.n529 10.6151
R1412 B.n415 B.n257 10.6151
R1413 B.n410 B.n257 10.6151
R1414 B.n410 B.n409 10.6151
R1415 B.n409 B.n408 10.6151
R1416 B.n408 B.n405 10.6151
R1417 B.n405 B.n404 10.6151
R1418 B.n404 B.n401 10.6151
R1419 B.n401 B.n400 10.6151
R1420 B.n400 B.n397 10.6151
R1421 B.n397 B.n396 10.6151
R1422 B.n396 B.n393 10.6151
R1423 B.n393 B.n392 10.6151
R1424 B.n392 B.n389 10.6151
R1425 B.n389 B.n388 10.6151
R1426 B.n388 B.n385 10.6151
R1427 B.n385 B.n384 10.6151
R1428 B.n384 B.n381 10.6151
R1429 B.n381 B.n380 10.6151
R1430 B.n380 B.n377 10.6151
R1431 B.n377 B.n376 10.6151
R1432 B.n376 B.n373 10.6151
R1433 B.n373 B.n372 10.6151
R1434 B.n372 B.n369 10.6151
R1435 B.n369 B.n368 10.6151
R1436 B.n368 B.n365 10.6151
R1437 B.n363 B.n360 10.6151
R1438 B.n360 B.n359 10.6151
R1439 B.n359 B.n356 10.6151
R1440 B.n356 B.n355 10.6151
R1441 B.n355 B.n352 10.6151
R1442 B.n352 B.n351 10.6151
R1443 B.n351 B.n348 10.6151
R1444 B.n348 B.n347 10.6151
R1445 B.n344 B.n343 10.6151
R1446 B.n343 B.n340 10.6151
R1447 B.n340 B.n339 10.6151
R1448 B.n339 B.n336 10.6151
R1449 B.n336 B.n335 10.6151
R1450 B.n335 B.n332 10.6151
R1451 B.n332 B.n331 10.6151
R1452 B.n331 B.n328 10.6151
R1453 B.n328 B.n327 10.6151
R1454 B.n327 B.n324 10.6151
R1455 B.n324 B.n323 10.6151
R1456 B.n323 B.n320 10.6151
R1457 B.n320 B.n319 10.6151
R1458 B.n319 B.n316 10.6151
R1459 B.n316 B.n315 10.6151
R1460 B.n315 B.n312 10.6151
R1461 B.n312 B.n311 10.6151
R1462 B.n311 B.n308 10.6151
R1463 B.n308 B.n307 10.6151
R1464 B.n307 B.n304 10.6151
R1465 B.n304 B.n303 10.6151
R1466 B.n303 B.n300 10.6151
R1467 B.n300 B.n299 10.6151
R1468 B.n299 B.n296 10.6151
R1469 B.n296 B.n295 10.6151
R1470 B.n417 B.n416 10.6151
R1471 B.n417 B.n249 10.6151
R1472 B.n427 B.n249 10.6151
R1473 B.n428 B.n427 10.6151
R1474 B.n429 B.n428 10.6151
R1475 B.n429 B.n241 10.6151
R1476 B.n439 B.n241 10.6151
R1477 B.n440 B.n439 10.6151
R1478 B.n441 B.n440 10.6151
R1479 B.n441 B.n233 10.6151
R1480 B.n452 B.n233 10.6151
R1481 B.n453 B.n452 10.6151
R1482 B.n454 B.n453 10.6151
R1483 B.n454 B.n226 10.6151
R1484 B.n464 B.n226 10.6151
R1485 B.n465 B.n464 10.6151
R1486 B.n466 B.n465 10.6151
R1487 B.n466 B.n218 10.6151
R1488 B.n476 B.n218 10.6151
R1489 B.n477 B.n476 10.6151
R1490 B.n478 B.n477 10.6151
R1491 B.n478 B.n210 10.6151
R1492 B.n489 B.n210 10.6151
R1493 B.n490 B.n489 10.6151
R1494 B.n491 B.n490 10.6151
R1495 B.n491 B.n0 10.6151
R1496 B.n586 B.n1 10.6151
R1497 B.n586 B.n585 10.6151
R1498 B.n585 B.n584 10.6151
R1499 B.n584 B.n10 10.6151
R1500 B.n578 B.n10 10.6151
R1501 B.n578 B.n577 10.6151
R1502 B.n577 B.n576 10.6151
R1503 B.n576 B.n17 10.6151
R1504 B.n570 B.n17 10.6151
R1505 B.n570 B.n569 10.6151
R1506 B.n569 B.n568 10.6151
R1507 B.n568 B.n24 10.6151
R1508 B.n562 B.n24 10.6151
R1509 B.n562 B.n561 10.6151
R1510 B.n561 B.n560 10.6151
R1511 B.n560 B.n30 10.6151
R1512 B.n554 B.n30 10.6151
R1513 B.n554 B.n553 10.6151
R1514 B.n553 B.n552 10.6151
R1515 B.n552 B.n38 10.6151
R1516 B.n546 B.n38 10.6151
R1517 B.n546 B.n545 10.6151
R1518 B.n545 B.n544 10.6151
R1519 B.n544 B.n45 10.6151
R1520 B.n538 B.n45 10.6151
R1521 B.n538 B.n537 10.6151
R1522 B.n431 B.t9 7.39235
R1523 B.n449 B.t7 7.39235
R1524 B.n32 B.t4 7.39235
R1525 B.t13 B.n548 7.39235
R1526 B.n139 B.n89 6.5566
R1527 B.n156 B.n155 6.5566
R1528 B.n364 B.n363 6.5566
R1529 B.n347 B.n293 6.5566
R1530 B.t6 B.n224 5.54439
R1531 B.t5 B.n22 5.54439
R1532 B.n136 B.n89 4.05904
R1533 B.n157 B.n156 4.05904
R1534 B.n365 B.n364 4.05904
R1535 B.n344 B.n293 4.05904
R1536 B.n592 B.n0 2.81026
R1537 B.n592 B.n1 2.81026
R1538 VN.n2 VN.t3 222.43
R1539 VN.n15 VN.t4 222.43
R1540 VN.n11 VN.t0 207.612
R1541 VN.n24 VN.t5 207.612
R1542 VN.n3 VN.t2 166.441
R1543 VN.n9 VN.t7 166.441
R1544 VN.n16 VN.t1 166.441
R1545 VN.n22 VN.t6 166.441
R1546 VN.n23 VN.n13 161.3
R1547 VN.n21 VN.n20 161.3
R1548 VN.n19 VN.n14 161.3
R1549 VN.n18 VN.n17 161.3
R1550 VN.n10 VN.n0 161.3
R1551 VN.n8 VN.n7 161.3
R1552 VN.n6 VN.n1 161.3
R1553 VN.n5 VN.n4 161.3
R1554 VN.n25 VN.n24 80.6037
R1555 VN.n12 VN.n11 80.6037
R1556 VN.n11 VN.n10 54.3172
R1557 VN.n24 VN.n23 54.3172
R1558 VN.n3 VN.n2 46.9212
R1559 VN.n16 VN.n15 46.9212
R1560 VN.n18 VN.n15 44.1937
R1561 VN.n5 VN.n2 44.1937
R1562 VN.n4 VN.n1 40.4934
R1563 VN.n8 VN.n1 40.4934
R1564 VN.n17 VN.n14 40.4934
R1565 VN.n21 VN.n14 40.4934
R1566 VN VN.n25 39.5975
R1567 VN.n10 VN.n9 17.3721
R1568 VN.n23 VN.n22 17.3721
R1569 VN.n4 VN.n3 7.09593
R1570 VN.n9 VN.n8 7.09593
R1571 VN.n17 VN.n16 7.09593
R1572 VN.n22 VN.n21 7.09593
R1573 VN.n25 VN.n13 0.285035
R1574 VN.n12 VN.n0 0.285035
R1575 VN.n20 VN.n13 0.189894
R1576 VN.n20 VN.n19 0.189894
R1577 VN.n19 VN.n18 0.189894
R1578 VN.n6 VN.n5 0.189894
R1579 VN.n7 VN.n6 0.189894
R1580 VN.n7 VN.n0 0.189894
R1581 VN VN.n12 0.146778
R1582 VDD2.n2 VDD2.n1 64.8292
R1583 VDD2.n2 VDD2.n0 64.8292
R1584 VDD2 VDD2.n5 64.8264
R1585 VDD2.n4 VDD2.n3 64.3287
R1586 VDD2.n4 VDD2.n2 34.4351
R1587 VDD2.n5 VDD2.t6 2.98693
R1588 VDD2.n5 VDD2.t3 2.98693
R1589 VDD2.n3 VDD2.t2 2.98693
R1590 VDD2.n3 VDD2.t1 2.98693
R1591 VDD2.n1 VDD2.t0 2.98693
R1592 VDD2.n1 VDD2.t7 2.98693
R1593 VDD2.n0 VDD2.t4 2.98693
R1594 VDD2.n0 VDD2.t5 2.98693
R1595 VDD2 VDD2.n4 0.614724
C0 VTAIL VDD2 6.47529f
C1 VDD1 VTAIL 6.43187f
C2 VTAIL VP 3.88118f
C3 VDD2 VN 3.71086f
C4 VDD1 VN 0.148814f
C5 VN VP 4.66309f
C6 VDD1 VDD2 0.95612f
C7 VDD2 VP 0.345209f
C8 VDD1 VP 3.90669f
C9 VTAIL VN 3.86708f
C10 VDD2 B 3.321292f
C11 VDD1 B 3.581624f
C12 VTAIL B 5.939304f
C13 VN B 8.82966f
C14 VP B 7.214141f
C15 VDD2.t4 B 0.135447f
C16 VDD2.t5 B 0.135447f
C17 VDD2.n0 B 1.14459f
C18 VDD2.t0 B 0.135447f
C19 VDD2.t7 B 0.135447f
C20 VDD2.n1 B 1.14459f
C21 VDD2.n2 B 2.06835f
C22 VDD2.t2 B 0.135447f
C23 VDD2.t1 B 0.135447f
C24 VDD2.n3 B 1.14182f
C25 VDD2.n4 B 2.02533f
C26 VDD2.t6 B 0.135447f
C27 VDD2.t3 B 0.135447f
C28 VDD2.n5 B 1.14456f
C29 VN.n0 B 0.053624f
C30 VN.t7 B 0.68078f
C31 VN.n1 B 0.032487f
C32 VN.t3 B 0.762143f
C33 VN.n2 B 0.331622f
C34 VN.t2 B 0.68078f
C35 VN.n3 B 0.308595f
C36 VN.n4 B 0.053615f
C37 VN.n5 B 0.168109f
C38 VN.n6 B 0.040187f
C39 VN.n7 B 0.040187f
C40 VN.n8 B 0.053615f
C41 VN.n9 B 0.275914f
C42 VN.n10 B 0.051895f
C43 VN.t0 B 0.739884f
C44 VN.n11 B 0.333853f
C45 VN.n12 B 0.037637f
C46 VN.n13 B 0.053624f
C47 VN.t6 B 0.68078f
C48 VN.n14 B 0.032487f
C49 VN.t4 B 0.762143f
C50 VN.n15 B 0.331622f
C51 VN.t1 B 0.68078f
C52 VN.n16 B 0.308595f
C53 VN.n17 B 0.053615f
C54 VN.n18 B 0.168109f
C55 VN.n19 B 0.040187f
C56 VN.n20 B 0.040187f
C57 VN.n21 B 0.053615f
C58 VN.n22 B 0.275914f
C59 VN.n23 B 0.051895f
C60 VN.t5 B 0.739884f
C61 VN.n24 B 0.333853f
C62 VN.n25 B 1.51891f
C63 VDD1.t4 B 0.135506f
C64 VDD1.t7 B 0.135506f
C65 VDD1.n0 B 1.1458f
C66 VDD1.t5 B 0.135506f
C67 VDD1.t6 B 0.135506f
C68 VDD1.n1 B 1.14509f
C69 VDD1.t0 B 0.135506f
C70 VDD1.t2 B 0.135506f
C71 VDD1.n2 B 1.14509f
C72 VDD1.n3 B 2.12446f
C73 VDD1.t1 B 0.135506f
C74 VDD1.t3 B 0.135506f
C75 VDD1.n4 B 1.14232f
C76 VDD1.n5 B 2.05685f
C77 VTAIL.t3 B 0.111302f
C78 VTAIL.t5 B 0.111302f
C79 VTAIL.n0 B 0.878489f
C80 VTAIL.n1 B 0.285851f
C81 VTAIL.n2 B 0.029143f
C82 VTAIL.n3 B 0.021244f
C83 VTAIL.n4 B 0.011416f
C84 VTAIL.n5 B 0.026982f
C85 VTAIL.n6 B 0.012087f
C86 VTAIL.n7 B 0.021244f
C87 VTAIL.n8 B 0.011416f
C88 VTAIL.n9 B 0.026982f
C89 VTAIL.n10 B 0.012087f
C90 VTAIL.n11 B 0.567051f
C91 VTAIL.n12 B 0.011416f
C92 VTAIL.t1 B 0.043945f
C93 VTAIL.n13 B 0.094107f
C94 VTAIL.n14 B 0.015939f
C95 VTAIL.n15 B 0.020237f
C96 VTAIL.n16 B 0.026982f
C97 VTAIL.n17 B 0.012087f
C98 VTAIL.n18 B 0.011416f
C99 VTAIL.n19 B 0.021244f
C100 VTAIL.n20 B 0.021244f
C101 VTAIL.n21 B 0.011416f
C102 VTAIL.n22 B 0.012087f
C103 VTAIL.n23 B 0.026982f
C104 VTAIL.n24 B 0.026982f
C105 VTAIL.n25 B 0.012087f
C106 VTAIL.n26 B 0.011416f
C107 VTAIL.n27 B 0.021244f
C108 VTAIL.n28 B 0.021244f
C109 VTAIL.n29 B 0.011416f
C110 VTAIL.n30 B 0.012087f
C111 VTAIL.n31 B 0.026982f
C112 VTAIL.n32 B 0.057145f
C113 VTAIL.n33 B 0.012087f
C114 VTAIL.n34 B 0.011416f
C115 VTAIL.n35 B 0.046492f
C116 VTAIL.n36 B 0.031762f
C117 VTAIL.n37 B 0.124957f
C118 VTAIL.n38 B 0.029143f
C119 VTAIL.n39 B 0.021244f
C120 VTAIL.n40 B 0.011416f
C121 VTAIL.n41 B 0.026982f
C122 VTAIL.n42 B 0.012087f
C123 VTAIL.n43 B 0.021244f
C124 VTAIL.n44 B 0.011416f
C125 VTAIL.n45 B 0.026982f
C126 VTAIL.n46 B 0.012087f
C127 VTAIL.n47 B 0.567051f
C128 VTAIL.n48 B 0.011416f
C129 VTAIL.t14 B 0.043945f
C130 VTAIL.n49 B 0.094107f
C131 VTAIL.n50 B 0.015939f
C132 VTAIL.n51 B 0.020237f
C133 VTAIL.n52 B 0.026982f
C134 VTAIL.n53 B 0.012087f
C135 VTAIL.n54 B 0.011416f
C136 VTAIL.n55 B 0.021244f
C137 VTAIL.n56 B 0.021244f
C138 VTAIL.n57 B 0.011416f
C139 VTAIL.n58 B 0.012087f
C140 VTAIL.n59 B 0.026982f
C141 VTAIL.n60 B 0.026982f
C142 VTAIL.n61 B 0.012087f
C143 VTAIL.n62 B 0.011416f
C144 VTAIL.n63 B 0.021244f
C145 VTAIL.n64 B 0.021244f
C146 VTAIL.n65 B 0.011416f
C147 VTAIL.n66 B 0.012087f
C148 VTAIL.n67 B 0.026982f
C149 VTAIL.n68 B 0.057145f
C150 VTAIL.n69 B 0.012087f
C151 VTAIL.n70 B 0.011416f
C152 VTAIL.n71 B 0.046492f
C153 VTAIL.n72 B 0.031762f
C154 VTAIL.n73 B 0.124957f
C155 VTAIL.t8 B 0.111302f
C156 VTAIL.t12 B 0.111302f
C157 VTAIL.n74 B 0.878489f
C158 VTAIL.n75 B 0.357992f
C159 VTAIL.n76 B 0.029143f
C160 VTAIL.n77 B 0.021244f
C161 VTAIL.n78 B 0.011416f
C162 VTAIL.n79 B 0.026982f
C163 VTAIL.n80 B 0.012087f
C164 VTAIL.n81 B 0.021244f
C165 VTAIL.n82 B 0.011416f
C166 VTAIL.n83 B 0.026982f
C167 VTAIL.n84 B 0.012087f
C168 VTAIL.n85 B 0.567051f
C169 VTAIL.n86 B 0.011416f
C170 VTAIL.t11 B 0.043945f
C171 VTAIL.n87 B 0.094107f
C172 VTAIL.n88 B 0.015939f
C173 VTAIL.n89 B 0.020237f
C174 VTAIL.n90 B 0.026982f
C175 VTAIL.n91 B 0.012087f
C176 VTAIL.n92 B 0.011416f
C177 VTAIL.n93 B 0.021244f
C178 VTAIL.n94 B 0.021244f
C179 VTAIL.n95 B 0.011416f
C180 VTAIL.n96 B 0.012087f
C181 VTAIL.n97 B 0.026982f
C182 VTAIL.n98 B 0.026982f
C183 VTAIL.n99 B 0.012087f
C184 VTAIL.n100 B 0.011416f
C185 VTAIL.n101 B 0.021244f
C186 VTAIL.n102 B 0.021244f
C187 VTAIL.n103 B 0.011416f
C188 VTAIL.n104 B 0.012087f
C189 VTAIL.n105 B 0.026982f
C190 VTAIL.n106 B 0.057145f
C191 VTAIL.n107 B 0.012087f
C192 VTAIL.n108 B 0.011416f
C193 VTAIL.n109 B 0.046492f
C194 VTAIL.n110 B 0.031762f
C195 VTAIL.n111 B 0.848735f
C196 VTAIL.n112 B 0.029143f
C197 VTAIL.n113 B 0.021244f
C198 VTAIL.n114 B 0.011416f
C199 VTAIL.n115 B 0.026982f
C200 VTAIL.n116 B 0.012087f
C201 VTAIL.n117 B 0.021244f
C202 VTAIL.n118 B 0.011416f
C203 VTAIL.n119 B 0.026982f
C204 VTAIL.n120 B 0.012087f
C205 VTAIL.n121 B 0.567051f
C206 VTAIL.n122 B 0.011416f
C207 VTAIL.t7 B 0.043945f
C208 VTAIL.n123 B 0.094107f
C209 VTAIL.n124 B 0.015939f
C210 VTAIL.n125 B 0.020237f
C211 VTAIL.n126 B 0.026982f
C212 VTAIL.n127 B 0.012087f
C213 VTAIL.n128 B 0.011416f
C214 VTAIL.n129 B 0.021244f
C215 VTAIL.n130 B 0.021244f
C216 VTAIL.n131 B 0.011416f
C217 VTAIL.n132 B 0.012087f
C218 VTAIL.n133 B 0.026982f
C219 VTAIL.n134 B 0.026982f
C220 VTAIL.n135 B 0.012087f
C221 VTAIL.n136 B 0.011416f
C222 VTAIL.n137 B 0.021244f
C223 VTAIL.n138 B 0.021244f
C224 VTAIL.n139 B 0.011416f
C225 VTAIL.n140 B 0.012087f
C226 VTAIL.n141 B 0.026982f
C227 VTAIL.n142 B 0.057145f
C228 VTAIL.n143 B 0.012087f
C229 VTAIL.n144 B 0.011416f
C230 VTAIL.n145 B 0.046492f
C231 VTAIL.n146 B 0.031762f
C232 VTAIL.n147 B 0.848735f
C233 VTAIL.t6 B 0.111302f
C234 VTAIL.t2 B 0.111302f
C235 VTAIL.n148 B 0.878495f
C236 VTAIL.n149 B 0.357986f
C237 VTAIL.n150 B 0.029143f
C238 VTAIL.n151 B 0.021244f
C239 VTAIL.n152 B 0.011416f
C240 VTAIL.n153 B 0.026982f
C241 VTAIL.n154 B 0.012087f
C242 VTAIL.n155 B 0.021244f
C243 VTAIL.n156 B 0.011416f
C244 VTAIL.n157 B 0.026982f
C245 VTAIL.n158 B 0.012087f
C246 VTAIL.n159 B 0.567051f
C247 VTAIL.n160 B 0.011416f
C248 VTAIL.t0 B 0.043945f
C249 VTAIL.n161 B 0.094107f
C250 VTAIL.n162 B 0.015939f
C251 VTAIL.n163 B 0.020237f
C252 VTAIL.n164 B 0.026982f
C253 VTAIL.n165 B 0.012087f
C254 VTAIL.n166 B 0.011416f
C255 VTAIL.n167 B 0.021244f
C256 VTAIL.n168 B 0.021244f
C257 VTAIL.n169 B 0.011416f
C258 VTAIL.n170 B 0.012087f
C259 VTAIL.n171 B 0.026982f
C260 VTAIL.n172 B 0.026982f
C261 VTAIL.n173 B 0.012087f
C262 VTAIL.n174 B 0.011416f
C263 VTAIL.n175 B 0.021244f
C264 VTAIL.n176 B 0.021244f
C265 VTAIL.n177 B 0.011416f
C266 VTAIL.n178 B 0.012087f
C267 VTAIL.n179 B 0.026982f
C268 VTAIL.n180 B 0.057145f
C269 VTAIL.n181 B 0.012087f
C270 VTAIL.n182 B 0.011416f
C271 VTAIL.n183 B 0.046492f
C272 VTAIL.n184 B 0.031762f
C273 VTAIL.n185 B 0.124957f
C274 VTAIL.n186 B 0.029143f
C275 VTAIL.n187 B 0.021244f
C276 VTAIL.n188 B 0.011416f
C277 VTAIL.n189 B 0.026982f
C278 VTAIL.n190 B 0.012087f
C279 VTAIL.n191 B 0.021244f
C280 VTAIL.n192 B 0.011416f
C281 VTAIL.n193 B 0.026982f
C282 VTAIL.n194 B 0.012087f
C283 VTAIL.n195 B 0.567051f
C284 VTAIL.n196 B 0.011416f
C285 VTAIL.t9 B 0.043945f
C286 VTAIL.n197 B 0.094107f
C287 VTAIL.n198 B 0.015939f
C288 VTAIL.n199 B 0.020237f
C289 VTAIL.n200 B 0.026982f
C290 VTAIL.n201 B 0.012087f
C291 VTAIL.n202 B 0.011416f
C292 VTAIL.n203 B 0.021244f
C293 VTAIL.n204 B 0.021244f
C294 VTAIL.n205 B 0.011416f
C295 VTAIL.n206 B 0.012087f
C296 VTAIL.n207 B 0.026982f
C297 VTAIL.n208 B 0.026982f
C298 VTAIL.n209 B 0.012087f
C299 VTAIL.n210 B 0.011416f
C300 VTAIL.n211 B 0.021244f
C301 VTAIL.n212 B 0.021244f
C302 VTAIL.n213 B 0.011416f
C303 VTAIL.n214 B 0.012087f
C304 VTAIL.n215 B 0.026982f
C305 VTAIL.n216 B 0.057145f
C306 VTAIL.n217 B 0.012087f
C307 VTAIL.n218 B 0.011416f
C308 VTAIL.n219 B 0.046492f
C309 VTAIL.n220 B 0.031762f
C310 VTAIL.n221 B 0.124957f
C311 VTAIL.t10 B 0.111302f
C312 VTAIL.t13 B 0.111302f
C313 VTAIL.n222 B 0.878495f
C314 VTAIL.n223 B 0.357986f
C315 VTAIL.n224 B 0.029143f
C316 VTAIL.n225 B 0.021244f
C317 VTAIL.n226 B 0.011416f
C318 VTAIL.n227 B 0.026982f
C319 VTAIL.n228 B 0.012087f
C320 VTAIL.n229 B 0.021244f
C321 VTAIL.n230 B 0.011416f
C322 VTAIL.n231 B 0.026982f
C323 VTAIL.n232 B 0.012087f
C324 VTAIL.n233 B 0.567051f
C325 VTAIL.n234 B 0.011416f
C326 VTAIL.t15 B 0.043945f
C327 VTAIL.n235 B 0.094107f
C328 VTAIL.n236 B 0.015939f
C329 VTAIL.n237 B 0.020237f
C330 VTAIL.n238 B 0.026982f
C331 VTAIL.n239 B 0.012087f
C332 VTAIL.n240 B 0.011416f
C333 VTAIL.n241 B 0.021244f
C334 VTAIL.n242 B 0.021244f
C335 VTAIL.n243 B 0.011416f
C336 VTAIL.n244 B 0.012087f
C337 VTAIL.n245 B 0.026982f
C338 VTAIL.n246 B 0.026982f
C339 VTAIL.n247 B 0.012087f
C340 VTAIL.n248 B 0.011416f
C341 VTAIL.n249 B 0.021244f
C342 VTAIL.n250 B 0.021244f
C343 VTAIL.n251 B 0.011416f
C344 VTAIL.n252 B 0.012087f
C345 VTAIL.n253 B 0.026982f
C346 VTAIL.n254 B 0.057145f
C347 VTAIL.n255 B 0.012087f
C348 VTAIL.n256 B 0.011416f
C349 VTAIL.n257 B 0.046492f
C350 VTAIL.n258 B 0.031762f
C351 VTAIL.n259 B 0.848735f
C352 VTAIL.n260 B 0.029143f
C353 VTAIL.n261 B 0.021244f
C354 VTAIL.n262 B 0.011416f
C355 VTAIL.n263 B 0.026982f
C356 VTAIL.n264 B 0.012087f
C357 VTAIL.n265 B 0.021244f
C358 VTAIL.n266 B 0.011416f
C359 VTAIL.n267 B 0.026982f
C360 VTAIL.n268 B 0.012087f
C361 VTAIL.n269 B 0.567051f
C362 VTAIL.n270 B 0.011416f
C363 VTAIL.t4 B 0.043945f
C364 VTAIL.n271 B 0.094107f
C365 VTAIL.n272 B 0.015939f
C366 VTAIL.n273 B 0.020237f
C367 VTAIL.n274 B 0.026982f
C368 VTAIL.n275 B 0.012087f
C369 VTAIL.n276 B 0.011416f
C370 VTAIL.n277 B 0.021244f
C371 VTAIL.n278 B 0.021244f
C372 VTAIL.n279 B 0.011416f
C373 VTAIL.n280 B 0.012087f
C374 VTAIL.n281 B 0.026982f
C375 VTAIL.n282 B 0.026982f
C376 VTAIL.n283 B 0.012087f
C377 VTAIL.n284 B 0.011416f
C378 VTAIL.n285 B 0.021244f
C379 VTAIL.n286 B 0.021244f
C380 VTAIL.n287 B 0.011416f
C381 VTAIL.n288 B 0.012087f
C382 VTAIL.n289 B 0.026982f
C383 VTAIL.n290 B 0.057145f
C384 VTAIL.n291 B 0.012087f
C385 VTAIL.n292 B 0.011416f
C386 VTAIL.n293 B 0.046492f
C387 VTAIL.n294 B 0.031762f
C388 VTAIL.n295 B 0.844752f
C389 VP.n0 B 0.054748f
C390 VP.t7 B 0.695042f
C391 VP.n1 B 0.033168f
C392 VP.n2 B 0.054748f
C393 VP.t1 B 0.695042f
C394 VP.n3 B 0.054748f
C395 VP.t4 B 0.755384f
C396 VP.t6 B 0.695042f
C397 VP.n4 B 0.033168f
C398 VP.t3 B 0.778109f
C399 VP.n5 B 0.338569f
C400 VP.t0 B 0.695042f
C401 VP.n6 B 0.31506f
C402 VP.n7 B 0.054738f
C403 VP.n8 B 0.171631f
C404 VP.n9 B 0.041029f
C405 VP.n10 B 0.041029f
C406 VP.n11 B 0.054738f
C407 VP.n12 B 0.281694f
C408 VP.n13 B 0.052982f
C409 VP.n14 B 0.340847f
C410 VP.n15 B 1.52743f
C411 VP.n16 B 1.56495f
C412 VP.t2 B 0.755384f
C413 VP.n17 B 0.340847f
C414 VP.n18 B 0.052982f
C415 VP.n19 B 0.281694f
C416 VP.n20 B 0.054738f
C417 VP.n21 B 0.041029f
C418 VP.n22 B 0.041029f
C419 VP.n23 B 0.041029f
C420 VP.n24 B 0.054738f
C421 VP.n25 B 0.281694f
C422 VP.n26 B 0.052982f
C423 VP.t5 B 0.755384f
C424 VP.n27 B 0.340847f
C425 VP.n28 B 0.038425f
.ends

