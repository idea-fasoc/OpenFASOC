* NGSPICE file created from diff_pair_sample_1234.ext - technology: sky130A

.subckt diff_pair_sample_1234 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=7.4529 pd=39 as=0 ps=0 w=19.11 l=2.7
X1 VTAIL.t14 VP.t0 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=3.15315 pd=19.44 as=3.15315 ps=19.44 w=19.11 l=2.7
X2 VDD1.t2 VP.t1 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=3.15315 pd=19.44 as=3.15315 ps=19.44 w=19.11 l=2.7
X3 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=7.4529 pd=39 as=0 ps=0 w=19.11 l=2.7
X4 VDD2.t7 VN.t0 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=3.15315 pd=19.44 as=3.15315 ps=19.44 w=19.11 l=2.7
X5 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=7.4529 pd=39 as=0 ps=0 w=19.11 l=2.7
X6 VTAIL.t4 VN.t1 VDD2.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=7.4529 pd=39 as=3.15315 ps=19.44 w=19.11 l=2.7
X7 VDD1.t1 VP.t2 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=3.15315 pd=19.44 as=3.15315 ps=19.44 w=19.11 l=2.7
X8 VTAIL.t15 VN.t2 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=3.15315 pd=19.44 as=3.15315 ps=19.44 w=19.11 l=2.7
X9 VTAIL.t11 VP.t3 VDD1.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=3.15315 pd=19.44 as=3.15315 ps=19.44 w=19.11 l=2.7
X10 VDD1.t5 VP.t4 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=3.15315 pd=19.44 as=7.4529 ps=39 w=19.11 l=2.7
X11 VTAIL.t2 VN.t3 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=7.4529 pd=39 as=3.15315 ps=19.44 w=19.11 l=2.7
X12 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.4529 pd=39 as=0 ps=0 w=19.11 l=2.7
X13 VDD1.t3 VP.t5 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=3.15315 pd=19.44 as=7.4529 ps=39 w=19.11 l=2.7
X14 VDD2.t3 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.15315 pd=19.44 as=7.4529 ps=39 w=19.11 l=2.7
X15 VTAIL.t8 VP.t6 VDD1.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=7.4529 pd=39 as=3.15315 ps=19.44 w=19.11 l=2.7
X16 VTAIL.t1 VN.t5 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=3.15315 pd=19.44 as=3.15315 ps=19.44 w=19.11 l=2.7
X17 VDD2.t1 VN.t6 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=3.15315 pd=19.44 as=7.4529 ps=39 w=19.11 l=2.7
X18 VTAIL.t7 VP.t7 VDD1.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=7.4529 pd=39 as=3.15315 ps=19.44 w=19.11 l=2.7
X19 VDD2.t0 VN.t7 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.15315 pd=19.44 as=3.15315 ps=19.44 w=19.11 l=2.7
R0 B.n1107 B.n1106 585
R1 B.n1108 B.n1107 585
R2 B.n436 B.n165 585
R3 B.n435 B.n434 585
R4 B.n433 B.n432 585
R5 B.n431 B.n430 585
R6 B.n429 B.n428 585
R7 B.n427 B.n426 585
R8 B.n425 B.n424 585
R9 B.n423 B.n422 585
R10 B.n421 B.n420 585
R11 B.n419 B.n418 585
R12 B.n417 B.n416 585
R13 B.n415 B.n414 585
R14 B.n413 B.n412 585
R15 B.n411 B.n410 585
R16 B.n409 B.n408 585
R17 B.n407 B.n406 585
R18 B.n405 B.n404 585
R19 B.n403 B.n402 585
R20 B.n401 B.n400 585
R21 B.n399 B.n398 585
R22 B.n397 B.n396 585
R23 B.n395 B.n394 585
R24 B.n393 B.n392 585
R25 B.n391 B.n390 585
R26 B.n389 B.n388 585
R27 B.n387 B.n386 585
R28 B.n385 B.n384 585
R29 B.n383 B.n382 585
R30 B.n381 B.n380 585
R31 B.n379 B.n378 585
R32 B.n377 B.n376 585
R33 B.n375 B.n374 585
R34 B.n373 B.n372 585
R35 B.n371 B.n370 585
R36 B.n369 B.n368 585
R37 B.n367 B.n366 585
R38 B.n365 B.n364 585
R39 B.n363 B.n362 585
R40 B.n361 B.n360 585
R41 B.n359 B.n358 585
R42 B.n357 B.n356 585
R43 B.n355 B.n354 585
R44 B.n353 B.n352 585
R45 B.n351 B.n350 585
R46 B.n349 B.n348 585
R47 B.n347 B.n346 585
R48 B.n345 B.n344 585
R49 B.n343 B.n342 585
R50 B.n341 B.n340 585
R51 B.n339 B.n338 585
R52 B.n337 B.n336 585
R53 B.n335 B.n334 585
R54 B.n333 B.n332 585
R55 B.n331 B.n330 585
R56 B.n329 B.n328 585
R57 B.n327 B.n326 585
R58 B.n325 B.n324 585
R59 B.n323 B.n322 585
R60 B.n321 B.n320 585
R61 B.n319 B.n318 585
R62 B.n317 B.n316 585
R63 B.n315 B.n314 585
R64 B.n313 B.n312 585
R65 B.n311 B.n310 585
R66 B.n309 B.n308 585
R67 B.n307 B.n306 585
R68 B.n305 B.n304 585
R69 B.n303 B.n302 585
R70 B.n301 B.n300 585
R71 B.n299 B.n298 585
R72 B.n297 B.n296 585
R73 B.n294 B.n293 585
R74 B.n292 B.n291 585
R75 B.n290 B.n289 585
R76 B.n288 B.n287 585
R77 B.n286 B.n285 585
R78 B.n284 B.n283 585
R79 B.n282 B.n281 585
R80 B.n280 B.n279 585
R81 B.n278 B.n277 585
R82 B.n276 B.n275 585
R83 B.n274 B.n273 585
R84 B.n272 B.n271 585
R85 B.n270 B.n269 585
R86 B.n268 B.n267 585
R87 B.n266 B.n265 585
R88 B.n264 B.n263 585
R89 B.n262 B.n261 585
R90 B.n260 B.n259 585
R91 B.n258 B.n257 585
R92 B.n256 B.n255 585
R93 B.n254 B.n253 585
R94 B.n252 B.n251 585
R95 B.n250 B.n249 585
R96 B.n248 B.n247 585
R97 B.n246 B.n245 585
R98 B.n244 B.n243 585
R99 B.n242 B.n241 585
R100 B.n240 B.n239 585
R101 B.n238 B.n237 585
R102 B.n236 B.n235 585
R103 B.n234 B.n233 585
R104 B.n232 B.n231 585
R105 B.n230 B.n229 585
R106 B.n228 B.n227 585
R107 B.n226 B.n225 585
R108 B.n224 B.n223 585
R109 B.n222 B.n221 585
R110 B.n220 B.n219 585
R111 B.n218 B.n217 585
R112 B.n216 B.n215 585
R113 B.n214 B.n213 585
R114 B.n212 B.n211 585
R115 B.n210 B.n209 585
R116 B.n208 B.n207 585
R117 B.n206 B.n205 585
R118 B.n204 B.n203 585
R119 B.n202 B.n201 585
R120 B.n200 B.n199 585
R121 B.n198 B.n197 585
R122 B.n196 B.n195 585
R123 B.n194 B.n193 585
R124 B.n192 B.n191 585
R125 B.n190 B.n189 585
R126 B.n188 B.n187 585
R127 B.n186 B.n185 585
R128 B.n184 B.n183 585
R129 B.n182 B.n181 585
R130 B.n180 B.n179 585
R131 B.n178 B.n177 585
R132 B.n176 B.n175 585
R133 B.n174 B.n173 585
R134 B.n172 B.n171 585
R135 B.n96 B.n95 585
R136 B.n1105 B.n97 585
R137 B.n1109 B.n97 585
R138 B.n1104 B.n1103 585
R139 B.n1103 B.n93 585
R140 B.n1102 B.n92 585
R141 B.n1115 B.n92 585
R142 B.n1101 B.n91 585
R143 B.n1116 B.n91 585
R144 B.n1100 B.n90 585
R145 B.n1117 B.n90 585
R146 B.n1099 B.n1098 585
R147 B.n1098 B.n86 585
R148 B.n1097 B.n85 585
R149 B.n1123 B.n85 585
R150 B.n1096 B.n84 585
R151 B.n1124 B.n84 585
R152 B.n1095 B.n83 585
R153 B.n1125 B.n83 585
R154 B.n1094 B.n1093 585
R155 B.n1093 B.n79 585
R156 B.n1092 B.n78 585
R157 B.n1131 B.n78 585
R158 B.n1091 B.n77 585
R159 B.n1132 B.n77 585
R160 B.n1090 B.n76 585
R161 B.n1133 B.n76 585
R162 B.n1089 B.n1088 585
R163 B.n1088 B.n72 585
R164 B.n1087 B.n71 585
R165 B.n1139 B.n71 585
R166 B.n1086 B.n70 585
R167 B.n1140 B.n70 585
R168 B.n1085 B.n69 585
R169 B.n1141 B.n69 585
R170 B.n1084 B.n1083 585
R171 B.n1083 B.n65 585
R172 B.n1082 B.n64 585
R173 B.n1147 B.n64 585
R174 B.n1081 B.n63 585
R175 B.n1148 B.n63 585
R176 B.n1080 B.n62 585
R177 B.n1149 B.n62 585
R178 B.n1079 B.n1078 585
R179 B.n1078 B.n58 585
R180 B.n1077 B.n57 585
R181 B.n1155 B.n57 585
R182 B.n1076 B.n56 585
R183 B.n1156 B.n56 585
R184 B.n1075 B.n55 585
R185 B.n1157 B.n55 585
R186 B.n1074 B.n1073 585
R187 B.n1073 B.n51 585
R188 B.n1072 B.n50 585
R189 B.n1163 B.n50 585
R190 B.n1071 B.n49 585
R191 B.n1164 B.n49 585
R192 B.n1070 B.n48 585
R193 B.n1165 B.n48 585
R194 B.n1069 B.n1068 585
R195 B.n1068 B.n44 585
R196 B.n1067 B.n43 585
R197 B.n1171 B.n43 585
R198 B.n1066 B.n42 585
R199 B.n1172 B.n42 585
R200 B.n1065 B.n41 585
R201 B.n1173 B.n41 585
R202 B.n1064 B.n1063 585
R203 B.n1063 B.n37 585
R204 B.n1062 B.n36 585
R205 B.n1179 B.n36 585
R206 B.n1061 B.n35 585
R207 B.n1180 B.n35 585
R208 B.n1060 B.n34 585
R209 B.n1181 B.n34 585
R210 B.n1059 B.n1058 585
R211 B.n1058 B.n33 585
R212 B.n1057 B.n29 585
R213 B.n1187 B.n29 585
R214 B.n1056 B.n28 585
R215 B.n1188 B.n28 585
R216 B.n1055 B.n27 585
R217 B.n1189 B.n27 585
R218 B.n1054 B.n1053 585
R219 B.n1053 B.n23 585
R220 B.n1052 B.n22 585
R221 B.n1195 B.n22 585
R222 B.n1051 B.n21 585
R223 B.n1196 B.n21 585
R224 B.n1050 B.n20 585
R225 B.n1197 B.n20 585
R226 B.n1049 B.n1048 585
R227 B.n1048 B.n16 585
R228 B.n1047 B.n15 585
R229 B.n1203 B.n15 585
R230 B.n1046 B.n14 585
R231 B.n1204 B.n14 585
R232 B.n1045 B.n13 585
R233 B.n1205 B.n13 585
R234 B.n1044 B.n1043 585
R235 B.n1043 B.n12 585
R236 B.n1042 B.n1041 585
R237 B.n1042 B.n8 585
R238 B.n1040 B.n7 585
R239 B.n1212 B.n7 585
R240 B.n1039 B.n6 585
R241 B.n1213 B.n6 585
R242 B.n1038 B.n5 585
R243 B.n1214 B.n5 585
R244 B.n1037 B.n1036 585
R245 B.n1036 B.n4 585
R246 B.n1035 B.n437 585
R247 B.n1035 B.n1034 585
R248 B.n1025 B.n438 585
R249 B.n439 B.n438 585
R250 B.n1027 B.n1026 585
R251 B.n1028 B.n1027 585
R252 B.n1024 B.n444 585
R253 B.n444 B.n443 585
R254 B.n1023 B.n1022 585
R255 B.n1022 B.n1021 585
R256 B.n446 B.n445 585
R257 B.n447 B.n446 585
R258 B.n1014 B.n1013 585
R259 B.n1015 B.n1014 585
R260 B.n1012 B.n452 585
R261 B.n452 B.n451 585
R262 B.n1011 B.n1010 585
R263 B.n1010 B.n1009 585
R264 B.n454 B.n453 585
R265 B.n455 B.n454 585
R266 B.n1002 B.n1001 585
R267 B.n1003 B.n1002 585
R268 B.n1000 B.n460 585
R269 B.n460 B.n459 585
R270 B.n999 B.n998 585
R271 B.n998 B.n997 585
R272 B.n462 B.n461 585
R273 B.n990 B.n462 585
R274 B.n989 B.n988 585
R275 B.n991 B.n989 585
R276 B.n987 B.n467 585
R277 B.n467 B.n466 585
R278 B.n986 B.n985 585
R279 B.n985 B.n984 585
R280 B.n469 B.n468 585
R281 B.n470 B.n469 585
R282 B.n977 B.n976 585
R283 B.n978 B.n977 585
R284 B.n975 B.n475 585
R285 B.n475 B.n474 585
R286 B.n974 B.n973 585
R287 B.n973 B.n972 585
R288 B.n477 B.n476 585
R289 B.n478 B.n477 585
R290 B.n965 B.n964 585
R291 B.n966 B.n965 585
R292 B.n963 B.n483 585
R293 B.n483 B.n482 585
R294 B.n962 B.n961 585
R295 B.n961 B.n960 585
R296 B.n485 B.n484 585
R297 B.n486 B.n485 585
R298 B.n953 B.n952 585
R299 B.n954 B.n953 585
R300 B.n951 B.n491 585
R301 B.n491 B.n490 585
R302 B.n950 B.n949 585
R303 B.n949 B.n948 585
R304 B.n493 B.n492 585
R305 B.n494 B.n493 585
R306 B.n941 B.n940 585
R307 B.n942 B.n941 585
R308 B.n939 B.n498 585
R309 B.n502 B.n498 585
R310 B.n938 B.n937 585
R311 B.n937 B.n936 585
R312 B.n500 B.n499 585
R313 B.n501 B.n500 585
R314 B.n929 B.n928 585
R315 B.n930 B.n929 585
R316 B.n927 B.n507 585
R317 B.n507 B.n506 585
R318 B.n926 B.n925 585
R319 B.n925 B.n924 585
R320 B.n509 B.n508 585
R321 B.n510 B.n509 585
R322 B.n917 B.n916 585
R323 B.n918 B.n917 585
R324 B.n915 B.n515 585
R325 B.n515 B.n514 585
R326 B.n914 B.n913 585
R327 B.n913 B.n912 585
R328 B.n517 B.n516 585
R329 B.n518 B.n517 585
R330 B.n905 B.n904 585
R331 B.n906 B.n905 585
R332 B.n903 B.n522 585
R333 B.n526 B.n522 585
R334 B.n902 B.n901 585
R335 B.n901 B.n900 585
R336 B.n524 B.n523 585
R337 B.n525 B.n524 585
R338 B.n893 B.n892 585
R339 B.n894 B.n893 585
R340 B.n891 B.n531 585
R341 B.n531 B.n530 585
R342 B.n890 B.n889 585
R343 B.n889 B.n888 585
R344 B.n533 B.n532 585
R345 B.n534 B.n533 585
R346 B.n881 B.n880 585
R347 B.n882 B.n881 585
R348 B.n537 B.n536 585
R349 B.n610 B.n609 585
R350 B.n611 B.n607 585
R351 B.n607 B.n538 585
R352 B.n613 B.n612 585
R353 B.n615 B.n606 585
R354 B.n618 B.n617 585
R355 B.n619 B.n605 585
R356 B.n621 B.n620 585
R357 B.n623 B.n604 585
R358 B.n626 B.n625 585
R359 B.n627 B.n603 585
R360 B.n629 B.n628 585
R361 B.n631 B.n602 585
R362 B.n634 B.n633 585
R363 B.n635 B.n601 585
R364 B.n637 B.n636 585
R365 B.n639 B.n600 585
R366 B.n642 B.n641 585
R367 B.n643 B.n599 585
R368 B.n645 B.n644 585
R369 B.n647 B.n598 585
R370 B.n650 B.n649 585
R371 B.n651 B.n597 585
R372 B.n653 B.n652 585
R373 B.n655 B.n596 585
R374 B.n658 B.n657 585
R375 B.n659 B.n595 585
R376 B.n661 B.n660 585
R377 B.n663 B.n594 585
R378 B.n666 B.n665 585
R379 B.n667 B.n593 585
R380 B.n669 B.n668 585
R381 B.n671 B.n592 585
R382 B.n674 B.n673 585
R383 B.n675 B.n591 585
R384 B.n677 B.n676 585
R385 B.n679 B.n590 585
R386 B.n682 B.n681 585
R387 B.n683 B.n589 585
R388 B.n685 B.n684 585
R389 B.n687 B.n588 585
R390 B.n690 B.n689 585
R391 B.n691 B.n587 585
R392 B.n693 B.n692 585
R393 B.n695 B.n586 585
R394 B.n698 B.n697 585
R395 B.n699 B.n585 585
R396 B.n701 B.n700 585
R397 B.n703 B.n584 585
R398 B.n706 B.n705 585
R399 B.n707 B.n583 585
R400 B.n709 B.n708 585
R401 B.n711 B.n582 585
R402 B.n714 B.n713 585
R403 B.n715 B.n581 585
R404 B.n717 B.n716 585
R405 B.n719 B.n580 585
R406 B.n722 B.n721 585
R407 B.n723 B.n579 585
R408 B.n725 B.n724 585
R409 B.n727 B.n578 585
R410 B.n730 B.n729 585
R411 B.n731 B.n575 585
R412 B.n734 B.n733 585
R413 B.n736 B.n574 585
R414 B.n739 B.n738 585
R415 B.n740 B.n573 585
R416 B.n742 B.n741 585
R417 B.n744 B.n572 585
R418 B.n747 B.n746 585
R419 B.n748 B.n571 585
R420 B.n753 B.n752 585
R421 B.n755 B.n570 585
R422 B.n758 B.n757 585
R423 B.n759 B.n569 585
R424 B.n761 B.n760 585
R425 B.n763 B.n568 585
R426 B.n766 B.n765 585
R427 B.n767 B.n567 585
R428 B.n769 B.n768 585
R429 B.n771 B.n566 585
R430 B.n774 B.n773 585
R431 B.n775 B.n565 585
R432 B.n777 B.n776 585
R433 B.n779 B.n564 585
R434 B.n782 B.n781 585
R435 B.n783 B.n563 585
R436 B.n785 B.n784 585
R437 B.n787 B.n562 585
R438 B.n790 B.n789 585
R439 B.n791 B.n561 585
R440 B.n793 B.n792 585
R441 B.n795 B.n560 585
R442 B.n798 B.n797 585
R443 B.n799 B.n559 585
R444 B.n801 B.n800 585
R445 B.n803 B.n558 585
R446 B.n806 B.n805 585
R447 B.n807 B.n557 585
R448 B.n809 B.n808 585
R449 B.n811 B.n556 585
R450 B.n814 B.n813 585
R451 B.n815 B.n555 585
R452 B.n817 B.n816 585
R453 B.n819 B.n554 585
R454 B.n822 B.n821 585
R455 B.n823 B.n553 585
R456 B.n825 B.n824 585
R457 B.n827 B.n552 585
R458 B.n830 B.n829 585
R459 B.n831 B.n551 585
R460 B.n833 B.n832 585
R461 B.n835 B.n550 585
R462 B.n838 B.n837 585
R463 B.n839 B.n549 585
R464 B.n841 B.n840 585
R465 B.n843 B.n548 585
R466 B.n846 B.n845 585
R467 B.n847 B.n547 585
R468 B.n849 B.n848 585
R469 B.n851 B.n546 585
R470 B.n854 B.n853 585
R471 B.n855 B.n545 585
R472 B.n857 B.n856 585
R473 B.n859 B.n544 585
R474 B.n862 B.n861 585
R475 B.n863 B.n543 585
R476 B.n865 B.n864 585
R477 B.n867 B.n542 585
R478 B.n870 B.n869 585
R479 B.n871 B.n541 585
R480 B.n873 B.n872 585
R481 B.n875 B.n540 585
R482 B.n878 B.n877 585
R483 B.n879 B.n539 585
R484 B.n884 B.n883 585
R485 B.n883 B.n882 585
R486 B.n885 B.n535 585
R487 B.n535 B.n534 585
R488 B.n887 B.n886 585
R489 B.n888 B.n887 585
R490 B.n529 B.n528 585
R491 B.n530 B.n529 585
R492 B.n896 B.n895 585
R493 B.n895 B.n894 585
R494 B.n897 B.n527 585
R495 B.n527 B.n525 585
R496 B.n899 B.n898 585
R497 B.n900 B.n899 585
R498 B.n521 B.n520 585
R499 B.n526 B.n521 585
R500 B.n908 B.n907 585
R501 B.n907 B.n906 585
R502 B.n909 B.n519 585
R503 B.n519 B.n518 585
R504 B.n911 B.n910 585
R505 B.n912 B.n911 585
R506 B.n513 B.n512 585
R507 B.n514 B.n513 585
R508 B.n920 B.n919 585
R509 B.n919 B.n918 585
R510 B.n921 B.n511 585
R511 B.n511 B.n510 585
R512 B.n923 B.n922 585
R513 B.n924 B.n923 585
R514 B.n505 B.n504 585
R515 B.n506 B.n505 585
R516 B.n932 B.n931 585
R517 B.n931 B.n930 585
R518 B.n933 B.n503 585
R519 B.n503 B.n501 585
R520 B.n935 B.n934 585
R521 B.n936 B.n935 585
R522 B.n497 B.n496 585
R523 B.n502 B.n497 585
R524 B.n944 B.n943 585
R525 B.n943 B.n942 585
R526 B.n945 B.n495 585
R527 B.n495 B.n494 585
R528 B.n947 B.n946 585
R529 B.n948 B.n947 585
R530 B.n489 B.n488 585
R531 B.n490 B.n489 585
R532 B.n956 B.n955 585
R533 B.n955 B.n954 585
R534 B.n957 B.n487 585
R535 B.n487 B.n486 585
R536 B.n959 B.n958 585
R537 B.n960 B.n959 585
R538 B.n481 B.n480 585
R539 B.n482 B.n481 585
R540 B.n968 B.n967 585
R541 B.n967 B.n966 585
R542 B.n969 B.n479 585
R543 B.n479 B.n478 585
R544 B.n971 B.n970 585
R545 B.n972 B.n971 585
R546 B.n473 B.n472 585
R547 B.n474 B.n473 585
R548 B.n980 B.n979 585
R549 B.n979 B.n978 585
R550 B.n981 B.n471 585
R551 B.n471 B.n470 585
R552 B.n983 B.n982 585
R553 B.n984 B.n983 585
R554 B.n465 B.n464 585
R555 B.n466 B.n465 585
R556 B.n993 B.n992 585
R557 B.n992 B.n991 585
R558 B.n994 B.n463 585
R559 B.n990 B.n463 585
R560 B.n996 B.n995 585
R561 B.n997 B.n996 585
R562 B.n458 B.n457 585
R563 B.n459 B.n458 585
R564 B.n1005 B.n1004 585
R565 B.n1004 B.n1003 585
R566 B.n1006 B.n456 585
R567 B.n456 B.n455 585
R568 B.n1008 B.n1007 585
R569 B.n1009 B.n1008 585
R570 B.n450 B.n449 585
R571 B.n451 B.n450 585
R572 B.n1017 B.n1016 585
R573 B.n1016 B.n1015 585
R574 B.n1018 B.n448 585
R575 B.n448 B.n447 585
R576 B.n1020 B.n1019 585
R577 B.n1021 B.n1020 585
R578 B.n442 B.n441 585
R579 B.n443 B.n442 585
R580 B.n1030 B.n1029 585
R581 B.n1029 B.n1028 585
R582 B.n1031 B.n440 585
R583 B.n440 B.n439 585
R584 B.n1033 B.n1032 585
R585 B.n1034 B.n1033 585
R586 B.n3 B.n0 585
R587 B.n4 B.n3 585
R588 B.n1211 B.n1 585
R589 B.n1212 B.n1211 585
R590 B.n1210 B.n1209 585
R591 B.n1210 B.n8 585
R592 B.n1208 B.n9 585
R593 B.n12 B.n9 585
R594 B.n1207 B.n1206 585
R595 B.n1206 B.n1205 585
R596 B.n11 B.n10 585
R597 B.n1204 B.n11 585
R598 B.n1202 B.n1201 585
R599 B.n1203 B.n1202 585
R600 B.n1200 B.n17 585
R601 B.n17 B.n16 585
R602 B.n1199 B.n1198 585
R603 B.n1198 B.n1197 585
R604 B.n19 B.n18 585
R605 B.n1196 B.n19 585
R606 B.n1194 B.n1193 585
R607 B.n1195 B.n1194 585
R608 B.n1192 B.n24 585
R609 B.n24 B.n23 585
R610 B.n1191 B.n1190 585
R611 B.n1190 B.n1189 585
R612 B.n26 B.n25 585
R613 B.n1188 B.n26 585
R614 B.n1186 B.n1185 585
R615 B.n1187 B.n1186 585
R616 B.n1184 B.n30 585
R617 B.n33 B.n30 585
R618 B.n1183 B.n1182 585
R619 B.n1182 B.n1181 585
R620 B.n32 B.n31 585
R621 B.n1180 B.n32 585
R622 B.n1178 B.n1177 585
R623 B.n1179 B.n1178 585
R624 B.n1176 B.n38 585
R625 B.n38 B.n37 585
R626 B.n1175 B.n1174 585
R627 B.n1174 B.n1173 585
R628 B.n40 B.n39 585
R629 B.n1172 B.n40 585
R630 B.n1170 B.n1169 585
R631 B.n1171 B.n1170 585
R632 B.n1168 B.n45 585
R633 B.n45 B.n44 585
R634 B.n1167 B.n1166 585
R635 B.n1166 B.n1165 585
R636 B.n47 B.n46 585
R637 B.n1164 B.n47 585
R638 B.n1162 B.n1161 585
R639 B.n1163 B.n1162 585
R640 B.n1160 B.n52 585
R641 B.n52 B.n51 585
R642 B.n1159 B.n1158 585
R643 B.n1158 B.n1157 585
R644 B.n54 B.n53 585
R645 B.n1156 B.n54 585
R646 B.n1154 B.n1153 585
R647 B.n1155 B.n1154 585
R648 B.n1152 B.n59 585
R649 B.n59 B.n58 585
R650 B.n1151 B.n1150 585
R651 B.n1150 B.n1149 585
R652 B.n61 B.n60 585
R653 B.n1148 B.n61 585
R654 B.n1146 B.n1145 585
R655 B.n1147 B.n1146 585
R656 B.n1144 B.n66 585
R657 B.n66 B.n65 585
R658 B.n1143 B.n1142 585
R659 B.n1142 B.n1141 585
R660 B.n68 B.n67 585
R661 B.n1140 B.n68 585
R662 B.n1138 B.n1137 585
R663 B.n1139 B.n1138 585
R664 B.n1136 B.n73 585
R665 B.n73 B.n72 585
R666 B.n1135 B.n1134 585
R667 B.n1134 B.n1133 585
R668 B.n75 B.n74 585
R669 B.n1132 B.n75 585
R670 B.n1130 B.n1129 585
R671 B.n1131 B.n1130 585
R672 B.n1128 B.n80 585
R673 B.n80 B.n79 585
R674 B.n1127 B.n1126 585
R675 B.n1126 B.n1125 585
R676 B.n82 B.n81 585
R677 B.n1124 B.n82 585
R678 B.n1122 B.n1121 585
R679 B.n1123 B.n1122 585
R680 B.n1120 B.n87 585
R681 B.n87 B.n86 585
R682 B.n1119 B.n1118 585
R683 B.n1118 B.n1117 585
R684 B.n89 B.n88 585
R685 B.n1116 B.n89 585
R686 B.n1114 B.n1113 585
R687 B.n1115 B.n1114 585
R688 B.n1112 B.n94 585
R689 B.n94 B.n93 585
R690 B.n1111 B.n1110 585
R691 B.n1110 B.n1109 585
R692 B.n1215 B.n1214 585
R693 B.n1213 B.n2 585
R694 B.n1110 B.n96 497.305
R695 B.n1107 B.n97 497.305
R696 B.n881 B.n539 497.305
R697 B.n883 B.n537 497.305
R698 B.n169 B.t16 378.767
R699 B.n166 B.t8 378.767
R700 B.n749 B.t12 378.767
R701 B.n576 B.t19 378.767
R702 B.n1108 B.n164 256.663
R703 B.n1108 B.n163 256.663
R704 B.n1108 B.n162 256.663
R705 B.n1108 B.n161 256.663
R706 B.n1108 B.n160 256.663
R707 B.n1108 B.n159 256.663
R708 B.n1108 B.n158 256.663
R709 B.n1108 B.n157 256.663
R710 B.n1108 B.n156 256.663
R711 B.n1108 B.n155 256.663
R712 B.n1108 B.n154 256.663
R713 B.n1108 B.n153 256.663
R714 B.n1108 B.n152 256.663
R715 B.n1108 B.n151 256.663
R716 B.n1108 B.n150 256.663
R717 B.n1108 B.n149 256.663
R718 B.n1108 B.n148 256.663
R719 B.n1108 B.n147 256.663
R720 B.n1108 B.n146 256.663
R721 B.n1108 B.n145 256.663
R722 B.n1108 B.n144 256.663
R723 B.n1108 B.n143 256.663
R724 B.n1108 B.n142 256.663
R725 B.n1108 B.n141 256.663
R726 B.n1108 B.n140 256.663
R727 B.n1108 B.n139 256.663
R728 B.n1108 B.n138 256.663
R729 B.n1108 B.n137 256.663
R730 B.n1108 B.n136 256.663
R731 B.n1108 B.n135 256.663
R732 B.n1108 B.n134 256.663
R733 B.n1108 B.n133 256.663
R734 B.n1108 B.n132 256.663
R735 B.n1108 B.n131 256.663
R736 B.n1108 B.n130 256.663
R737 B.n1108 B.n129 256.663
R738 B.n1108 B.n128 256.663
R739 B.n1108 B.n127 256.663
R740 B.n1108 B.n126 256.663
R741 B.n1108 B.n125 256.663
R742 B.n1108 B.n124 256.663
R743 B.n1108 B.n123 256.663
R744 B.n1108 B.n122 256.663
R745 B.n1108 B.n121 256.663
R746 B.n1108 B.n120 256.663
R747 B.n1108 B.n119 256.663
R748 B.n1108 B.n118 256.663
R749 B.n1108 B.n117 256.663
R750 B.n1108 B.n116 256.663
R751 B.n1108 B.n115 256.663
R752 B.n1108 B.n114 256.663
R753 B.n1108 B.n113 256.663
R754 B.n1108 B.n112 256.663
R755 B.n1108 B.n111 256.663
R756 B.n1108 B.n110 256.663
R757 B.n1108 B.n109 256.663
R758 B.n1108 B.n108 256.663
R759 B.n1108 B.n107 256.663
R760 B.n1108 B.n106 256.663
R761 B.n1108 B.n105 256.663
R762 B.n1108 B.n104 256.663
R763 B.n1108 B.n103 256.663
R764 B.n1108 B.n102 256.663
R765 B.n1108 B.n101 256.663
R766 B.n1108 B.n100 256.663
R767 B.n1108 B.n99 256.663
R768 B.n1108 B.n98 256.663
R769 B.n608 B.n538 256.663
R770 B.n614 B.n538 256.663
R771 B.n616 B.n538 256.663
R772 B.n622 B.n538 256.663
R773 B.n624 B.n538 256.663
R774 B.n630 B.n538 256.663
R775 B.n632 B.n538 256.663
R776 B.n638 B.n538 256.663
R777 B.n640 B.n538 256.663
R778 B.n646 B.n538 256.663
R779 B.n648 B.n538 256.663
R780 B.n654 B.n538 256.663
R781 B.n656 B.n538 256.663
R782 B.n662 B.n538 256.663
R783 B.n664 B.n538 256.663
R784 B.n670 B.n538 256.663
R785 B.n672 B.n538 256.663
R786 B.n678 B.n538 256.663
R787 B.n680 B.n538 256.663
R788 B.n686 B.n538 256.663
R789 B.n688 B.n538 256.663
R790 B.n694 B.n538 256.663
R791 B.n696 B.n538 256.663
R792 B.n702 B.n538 256.663
R793 B.n704 B.n538 256.663
R794 B.n710 B.n538 256.663
R795 B.n712 B.n538 256.663
R796 B.n718 B.n538 256.663
R797 B.n720 B.n538 256.663
R798 B.n726 B.n538 256.663
R799 B.n728 B.n538 256.663
R800 B.n735 B.n538 256.663
R801 B.n737 B.n538 256.663
R802 B.n743 B.n538 256.663
R803 B.n745 B.n538 256.663
R804 B.n754 B.n538 256.663
R805 B.n756 B.n538 256.663
R806 B.n762 B.n538 256.663
R807 B.n764 B.n538 256.663
R808 B.n770 B.n538 256.663
R809 B.n772 B.n538 256.663
R810 B.n778 B.n538 256.663
R811 B.n780 B.n538 256.663
R812 B.n786 B.n538 256.663
R813 B.n788 B.n538 256.663
R814 B.n794 B.n538 256.663
R815 B.n796 B.n538 256.663
R816 B.n802 B.n538 256.663
R817 B.n804 B.n538 256.663
R818 B.n810 B.n538 256.663
R819 B.n812 B.n538 256.663
R820 B.n818 B.n538 256.663
R821 B.n820 B.n538 256.663
R822 B.n826 B.n538 256.663
R823 B.n828 B.n538 256.663
R824 B.n834 B.n538 256.663
R825 B.n836 B.n538 256.663
R826 B.n842 B.n538 256.663
R827 B.n844 B.n538 256.663
R828 B.n850 B.n538 256.663
R829 B.n852 B.n538 256.663
R830 B.n858 B.n538 256.663
R831 B.n860 B.n538 256.663
R832 B.n866 B.n538 256.663
R833 B.n868 B.n538 256.663
R834 B.n874 B.n538 256.663
R835 B.n876 B.n538 256.663
R836 B.n1217 B.n1216 256.663
R837 B.n173 B.n172 163.367
R838 B.n177 B.n176 163.367
R839 B.n181 B.n180 163.367
R840 B.n185 B.n184 163.367
R841 B.n189 B.n188 163.367
R842 B.n193 B.n192 163.367
R843 B.n197 B.n196 163.367
R844 B.n201 B.n200 163.367
R845 B.n205 B.n204 163.367
R846 B.n209 B.n208 163.367
R847 B.n213 B.n212 163.367
R848 B.n217 B.n216 163.367
R849 B.n221 B.n220 163.367
R850 B.n225 B.n224 163.367
R851 B.n229 B.n228 163.367
R852 B.n233 B.n232 163.367
R853 B.n237 B.n236 163.367
R854 B.n241 B.n240 163.367
R855 B.n245 B.n244 163.367
R856 B.n249 B.n248 163.367
R857 B.n253 B.n252 163.367
R858 B.n257 B.n256 163.367
R859 B.n261 B.n260 163.367
R860 B.n265 B.n264 163.367
R861 B.n269 B.n268 163.367
R862 B.n273 B.n272 163.367
R863 B.n277 B.n276 163.367
R864 B.n281 B.n280 163.367
R865 B.n285 B.n284 163.367
R866 B.n289 B.n288 163.367
R867 B.n293 B.n292 163.367
R868 B.n298 B.n297 163.367
R869 B.n302 B.n301 163.367
R870 B.n306 B.n305 163.367
R871 B.n310 B.n309 163.367
R872 B.n314 B.n313 163.367
R873 B.n318 B.n317 163.367
R874 B.n322 B.n321 163.367
R875 B.n326 B.n325 163.367
R876 B.n330 B.n329 163.367
R877 B.n334 B.n333 163.367
R878 B.n338 B.n337 163.367
R879 B.n342 B.n341 163.367
R880 B.n346 B.n345 163.367
R881 B.n350 B.n349 163.367
R882 B.n354 B.n353 163.367
R883 B.n358 B.n357 163.367
R884 B.n362 B.n361 163.367
R885 B.n366 B.n365 163.367
R886 B.n370 B.n369 163.367
R887 B.n374 B.n373 163.367
R888 B.n378 B.n377 163.367
R889 B.n382 B.n381 163.367
R890 B.n386 B.n385 163.367
R891 B.n390 B.n389 163.367
R892 B.n394 B.n393 163.367
R893 B.n398 B.n397 163.367
R894 B.n402 B.n401 163.367
R895 B.n406 B.n405 163.367
R896 B.n410 B.n409 163.367
R897 B.n414 B.n413 163.367
R898 B.n418 B.n417 163.367
R899 B.n422 B.n421 163.367
R900 B.n426 B.n425 163.367
R901 B.n430 B.n429 163.367
R902 B.n434 B.n433 163.367
R903 B.n1107 B.n165 163.367
R904 B.n881 B.n533 163.367
R905 B.n889 B.n533 163.367
R906 B.n889 B.n531 163.367
R907 B.n893 B.n531 163.367
R908 B.n893 B.n524 163.367
R909 B.n901 B.n524 163.367
R910 B.n901 B.n522 163.367
R911 B.n905 B.n522 163.367
R912 B.n905 B.n517 163.367
R913 B.n913 B.n517 163.367
R914 B.n913 B.n515 163.367
R915 B.n917 B.n515 163.367
R916 B.n917 B.n509 163.367
R917 B.n925 B.n509 163.367
R918 B.n925 B.n507 163.367
R919 B.n929 B.n507 163.367
R920 B.n929 B.n500 163.367
R921 B.n937 B.n500 163.367
R922 B.n937 B.n498 163.367
R923 B.n941 B.n498 163.367
R924 B.n941 B.n493 163.367
R925 B.n949 B.n493 163.367
R926 B.n949 B.n491 163.367
R927 B.n953 B.n491 163.367
R928 B.n953 B.n485 163.367
R929 B.n961 B.n485 163.367
R930 B.n961 B.n483 163.367
R931 B.n965 B.n483 163.367
R932 B.n965 B.n477 163.367
R933 B.n973 B.n477 163.367
R934 B.n973 B.n475 163.367
R935 B.n977 B.n475 163.367
R936 B.n977 B.n469 163.367
R937 B.n985 B.n469 163.367
R938 B.n985 B.n467 163.367
R939 B.n989 B.n467 163.367
R940 B.n989 B.n462 163.367
R941 B.n998 B.n462 163.367
R942 B.n998 B.n460 163.367
R943 B.n1002 B.n460 163.367
R944 B.n1002 B.n454 163.367
R945 B.n1010 B.n454 163.367
R946 B.n1010 B.n452 163.367
R947 B.n1014 B.n452 163.367
R948 B.n1014 B.n446 163.367
R949 B.n1022 B.n446 163.367
R950 B.n1022 B.n444 163.367
R951 B.n1027 B.n444 163.367
R952 B.n1027 B.n438 163.367
R953 B.n1035 B.n438 163.367
R954 B.n1036 B.n1035 163.367
R955 B.n1036 B.n5 163.367
R956 B.n6 B.n5 163.367
R957 B.n7 B.n6 163.367
R958 B.n1042 B.n7 163.367
R959 B.n1043 B.n1042 163.367
R960 B.n1043 B.n13 163.367
R961 B.n14 B.n13 163.367
R962 B.n15 B.n14 163.367
R963 B.n1048 B.n15 163.367
R964 B.n1048 B.n20 163.367
R965 B.n21 B.n20 163.367
R966 B.n22 B.n21 163.367
R967 B.n1053 B.n22 163.367
R968 B.n1053 B.n27 163.367
R969 B.n28 B.n27 163.367
R970 B.n29 B.n28 163.367
R971 B.n1058 B.n29 163.367
R972 B.n1058 B.n34 163.367
R973 B.n35 B.n34 163.367
R974 B.n36 B.n35 163.367
R975 B.n1063 B.n36 163.367
R976 B.n1063 B.n41 163.367
R977 B.n42 B.n41 163.367
R978 B.n43 B.n42 163.367
R979 B.n1068 B.n43 163.367
R980 B.n1068 B.n48 163.367
R981 B.n49 B.n48 163.367
R982 B.n50 B.n49 163.367
R983 B.n1073 B.n50 163.367
R984 B.n1073 B.n55 163.367
R985 B.n56 B.n55 163.367
R986 B.n57 B.n56 163.367
R987 B.n1078 B.n57 163.367
R988 B.n1078 B.n62 163.367
R989 B.n63 B.n62 163.367
R990 B.n64 B.n63 163.367
R991 B.n1083 B.n64 163.367
R992 B.n1083 B.n69 163.367
R993 B.n70 B.n69 163.367
R994 B.n71 B.n70 163.367
R995 B.n1088 B.n71 163.367
R996 B.n1088 B.n76 163.367
R997 B.n77 B.n76 163.367
R998 B.n78 B.n77 163.367
R999 B.n1093 B.n78 163.367
R1000 B.n1093 B.n83 163.367
R1001 B.n84 B.n83 163.367
R1002 B.n85 B.n84 163.367
R1003 B.n1098 B.n85 163.367
R1004 B.n1098 B.n90 163.367
R1005 B.n91 B.n90 163.367
R1006 B.n92 B.n91 163.367
R1007 B.n1103 B.n92 163.367
R1008 B.n1103 B.n97 163.367
R1009 B.n609 B.n607 163.367
R1010 B.n613 B.n607 163.367
R1011 B.n617 B.n615 163.367
R1012 B.n621 B.n605 163.367
R1013 B.n625 B.n623 163.367
R1014 B.n629 B.n603 163.367
R1015 B.n633 B.n631 163.367
R1016 B.n637 B.n601 163.367
R1017 B.n641 B.n639 163.367
R1018 B.n645 B.n599 163.367
R1019 B.n649 B.n647 163.367
R1020 B.n653 B.n597 163.367
R1021 B.n657 B.n655 163.367
R1022 B.n661 B.n595 163.367
R1023 B.n665 B.n663 163.367
R1024 B.n669 B.n593 163.367
R1025 B.n673 B.n671 163.367
R1026 B.n677 B.n591 163.367
R1027 B.n681 B.n679 163.367
R1028 B.n685 B.n589 163.367
R1029 B.n689 B.n687 163.367
R1030 B.n693 B.n587 163.367
R1031 B.n697 B.n695 163.367
R1032 B.n701 B.n585 163.367
R1033 B.n705 B.n703 163.367
R1034 B.n709 B.n583 163.367
R1035 B.n713 B.n711 163.367
R1036 B.n717 B.n581 163.367
R1037 B.n721 B.n719 163.367
R1038 B.n725 B.n579 163.367
R1039 B.n729 B.n727 163.367
R1040 B.n734 B.n575 163.367
R1041 B.n738 B.n736 163.367
R1042 B.n742 B.n573 163.367
R1043 B.n746 B.n744 163.367
R1044 B.n753 B.n571 163.367
R1045 B.n757 B.n755 163.367
R1046 B.n761 B.n569 163.367
R1047 B.n765 B.n763 163.367
R1048 B.n769 B.n567 163.367
R1049 B.n773 B.n771 163.367
R1050 B.n777 B.n565 163.367
R1051 B.n781 B.n779 163.367
R1052 B.n785 B.n563 163.367
R1053 B.n789 B.n787 163.367
R1054 B.n793 B.n561 163.367
R1055 B.n797 B.n795 163.367
R1056 B.n801 B.n559 163.367
R1057 B.n805 B.n803 163.367
R1058 B.n809 B.n557 163.367
R1059 B.n813 B.n811 163.367
R1060 B.n817 B.n555 163.367
R1061 B.n821 B.n819 163.367
R1062 B.n825 B.n553 163.367
R1063 B.n829 B.n827 163.367
R1064 B.n833 B.n551 163.367
R1065 B.n837 B.n835 163.367
R1066 B.n841 B.n549 163.367
R1067 B.n845 B.n843 163.367
R1068 B.n849 B.n547 163.367
R1069 B.n853 B.n851 163.367
R1070 B.n857 B.n545 163.367
R1071 B.n861 B.n859 163.367
R1072 B.n865 B.n543 163.367
R1073 B.n869 B.n867 163.367
R1074 B.n873 B.n541 163.367
R1075 B.n877 B.n875 163.367
R1076 B.n883 B.n535 163.367
R1077 B.n887 B.n535 163.367
R1078 B.n887 B.n529 163.367
R1079 B.n895 B.n529 163.367
R1080 B.n895 B.n527 163.367
R1081 B.n899 B.n527 163.367
R1082 B.n899 B.n521 163.367
R1083 B.n907 B.n521 163.367
R1084 B.n907 B.n519 163.367
R1085 B.n911 B.n519 163.367
R1086 B.n911 B.n513 163.367
R1087 B.n919 B.n513 163.367
R1088 B.n919 B.n511 163.367
R1089 B.n923 B.n511 163.367
R1090 B.n923 B.n505 163.367
R1091 B.n931 B.n505 163.367
R1092 B.n931 B.n503 163.367
R1093 B.n935 B.n503 163.367
R1094 B.n935 B.n497 163.367
R1095 B.n943 B.n497 163.367
R1096 B.n943 B.n495 163.367
R1097 B.n947 B.n495 163.367
R1098 B.n947 B.n489 163.367
R1099 B.n955 B.n489 163.367
R1100 B.n955 B.n487 163.367
R1101 B.n959 B.n487 163.367
R1102 B.n959 B.n481 163.367
R1103 B.n967 B.n481 163.367
R1104 B.n967 B.n479 163.367
R1105 B.n971 B.n479 163.367
R1106 B.n971 B.n473 163.367
R1107 B.n979 B.n473 163.367
R1108 B.n979 B.n471 163.367
R1109 B.n983 B.n471 163.367
R1110 B.n983 B.n465 163.367
R1111 B.n992 B.n465 163.367
R1112 B.n992 B.n463 163.367
R1113 B.n996 B.n463 163.367
R1114 B.n996 B.n458 163.367
R1115 B.n1004 B.n458 163.367
R1116 B.n1004 B.n456 163.367
R1117 B.n1008 B.n456 163.367
R1118 B.n1008 B.n450 163.367
R1119 B.n1016 B.n450 163.367
R1120 B.n1016 B.n448 163.367
R1121 B.n1020 B.n448 163.367
R1122 B.n1020 B.n442 163.367
R1123 B.n1029 B.n442 163.367
R1124 B.n1029 B.n440 163.367
R1125 B.n1033 B.n440 163.367
R1126 B.n1033 B.n3 163.367
R1127 B.n1215 B.n3 163.367
R1128 B.n1211 B.n2 163.367
R1129 B.n1211 B.n1210 163.367
R1130 B.n1210 B.n9 163.367
R1131 B.n1206 B.n9 163.367
R1132 B.n1206 B.n11 163.367
R1133 B.n1202 B.n11 163.367
R1134 B.n1202 B.n17 163.367
R1135 B.n1198 B.n17 163.367
R1136 B.n1198 B.n19 163.367
R1137 B.n1194 B.n19 163.367
R1138 B.n1194 B.n24 163.367
R1139 B.n1190 B.n24 163.367
R1140 B.n1190 B.n26 163.367
R1141 B.n1186 B.n26 163.367
R1142 B.n1186 B.n30 163.367
R1143 B.n1182 B.n30 163.367
R1144 B.n1182 B.n32 163.367
R1145 B.n1178 B.n32 163.367
R1146 B.n1178 B.n38 163.367
R1147 B.n1174 B.n38 163.367
R1148 B.n1174 B.n40 163.367
R1149 B.n1170 B.n40 163.367
R1150 B.n1170 B.n45 163.367
R1151 B.n1166 B.n45 163.367
R1152 B.n1166 B.n47 163.367
R1153 B.n1162 B.n47 163.367
R1154 B.n1162 B.n52 163.367
R1155 B.n1158 B.n52 163.367
R1156 B.n1158 B.n54 163.367
R1157 B.n1154 B.n54 163.367
R1158 B.n1154 B.n59 163.367
R1159 B.n1150 B.n59 163.367
R1160 B.n1150 B.n61 163.367
R1161 B.n1146 B.n61 163.367
R1162 B.n1146 B.n66 163.367
R1163 B.n1142 B.n66 163.367
R1164 B.n1142 B.n68 163.367
R1165 B.n1138 B.n68 163.367
R1166 B.n1138 B.n73 163.367
R1167 B.n1134 B.n73 163.367
R1168 B.n1134 B.n75 163.367
R1169 B.n1130 B.n75 163.367
R1170 B.n1130 B.n80 163.367
R1171 B.n1126 B.n80 163.367
R1172 B.n1126 B.n82 163.367
R1173 B.n1122 B.n82 163.367
R1174 B.n1122 B.n87 163.367
R1175 B.n1118 B.n87 163.367
R1176 B.n1118 B.n89 163.367
R1177 B.n1114 B.n89 163.367
R1178 B.n1114 B.n94 163.367
R1179 B.n1110 B.n94 163.367
R1180 B.n166 B.t10 127.308
R1181 B.n749 B.t15 127.308
R1182 B.n169 B.t17 127.281
R1183 B.n576 B.t21 127.281
R1184 B.n98 B.n96 71.676
R1185 B.n173 B.n99 71.676
R1186 B.n177 B.n100 71.676
R1187 B.n181 B.n101 71.676
R1188 B.n185 B.n102 71.676
R1189 B.n189 B.n103 71.676
R1190 B.n193 B.n104 71.676
R1191 B.n197 B.n105 71.676
R1192 B.n201 B.n106 71.676
R1193 B.n205 B.n107 71.676
R1194 B.n209 B.n108 71.676
R1195 B.n213 B.n109 71.676
R1196 B.n217 B.n110 71.676
R1197 B.n221 B.n111 71.676
R1198 B.n225 B.n112 71.676
R1199 B.n229 B.n113 71.676
R1200 B.n233 B.n114 71.676
R1201 B.n237 B.n115 71.676
R1202 B.n241 B.n116 71.676
R1203 B.n245 B.n117 71.676
R1204 B.n249 B.n118 71.676
R1205 B.n253 B.n119 71.676
R1206 B.n257 B.n120 71.676
R1207 B.n261 B.n121 71.676
R1208 B.n265 B.n122 71.676
R1209 B.n269 B.n123 71.676
R1210 B.n273 B.n124 71.676
R1211 B.n277 B.n125 71.676
R1212 B.n281 B.n126 71.676
R1213 B.n285 B.n127 71.676
R1214 B.n289 B.n128 71.676
R1215 B.n293 B.n129 71.676
R1216 B.n298 B.n130 71.676
R1217 B.n302 B.n131 71.676
R1218 B.n306 B.n132 71.676
R1219 B.n310 B.n133 71.676
R1220 B.n314 B.n134 71.676
R1221 B.n318 B.n135 71.676
R1222 B.n322 B.n136 71.676
R1223 B.n326 B.n137 71.676
R1224 B.n330 B.n138 71.676
R1225 B.n334 B.n139 71.676
R1226 B.n338 B.n140 71.676
R1227 B.n342 B.n141 71.676
R1228 B.n346 B.n142 71.676
R1229 B.n350 B.n143 71.676
R1230 B.n354 B.n144 71.676
R1231 B.n358 B.n145 71.676
R1232 B.n362 B.n146 71.676
R1233 B.n366 B.n147 71.676
R1234 B.n370 B.n148 71.676
R1235 B.n374 B.n149 71.676
R1236 B.n378 B.n150 71.676
R1237 B.n382 B.n151 71.676
R1238 B.n386 B.n152 71.676
R1239 B.n390 B.n153 71.676
R1240 B.n394 B.n154 71.676
R1241 B.n398 B.n155 71.676
R1242 B.n402 B.n156 71.676
R1243 B.n406 B.n157 71.676
R1244 B.n410 B.n158 71.676
R1245 B.n414 B.n159 71.676
R1246 B.n418 B.n160 71.676
R1247 B.n422 B.n161 71.676
R1248 B.n426 B.n162 71.676
R1249 B.n430 B.n163 71.676
R1250 B.n434 B.n164 71.676
R1251 B.n165 B.n164 71.676
R1252 B.n433 B.n163 71.676
R1253 B.n429 B.n162 71.676
R1254 B.n425 B.n161 71.676
R1255 B.n421 B.n160 71.676
R1256 B.n417 B.n159 71.676
R1257 B.n413 B.n158 71.676
R1258 B.n409 B.n157 71.676
R1259 B.n405 B.n156 71.676
R1260 B.n401 B.n155 71.676
R1261 B.n397 B.n154 71.676
R1262 B.n393 B.n153 71.676
R1263 B.n389 B.n152 71.676
R1264 B.n385 B.n151 71.676
R1265 B.n381 B.n150 71.676
R1266 B.n377 B.n149 71.676
R1267 B.n373 B.n148 71.676
R1268 B.n369 B.n147 71.676
R1269 B.n365 B.n146 71.676
R1270 B.n361 B.n145 71.676
R1271 B.n357 B.n144 71.676
R1272 B.n353 B.n143 71.676
R1273 B.n349 B.n142 71.676
R1274 B.n345 B.n141 71.676
R1275 B.n341 B.n140 71.676
R1276 B.n337 B.n139 71.676
R1277 B.n333 B.n138 71.676
R1278 B.n329 B.n137 71.676
R1279 B.n325 B.n136 71.676
R1280 B.n321 B.n135 71.676
R1281 B.n317 B.n134 71.676
R1282 B.n313 B.n133 71.676
R1283 B.n309 B.n132 71.676
R1284 B.n305 B.n131 71.676
R1285 B.n301 B.n130 71.676
R1286 B.n297 B.n129 71.676
R1287 B.n292 B.n128 71.676
R1288 B.n288 B.n127 71.676
R1289 B.n284 B.n126 71.676
R1290 B.n280 B.n125 71.676
R1291 B.n276 B.n124 71.676
R1292 B.n272 B.n123 71.676
R1293 B.n268 B.n122 71.676
R1294 B.n264 B.n121 71.676
R1295 B.n260 B.n120 71.676
R1296 B.n256 B.n119 71.676
R1297 B.n252 B.n118 71.676
R1298 B.n248 B.n117 71.676
R1299 B.n244 B.n116 71.676
R1300 B.n240 B.n115 71.676
R1301 B.n236 B.n114 71.676
R1302 B.n232 B.n113 71.676
R1303 B.n228 B.n112 71.676
R1304 B.n224 B.n111 71.676
R1305 B.n220 B.n110 71.676
R1306 B.n216 B.n109 71.676
R1307 B.n212 B.n108 71.676
R1308 B.n208 B.n107 71.676
R1309 B.n204 B.n106 71.676
R1310 B.n200 B.n105 71.676
R1311 B.n196 B.n104 71.676
R1312 B.n192 B.n103 71.676
R1313 B.n188 B.n102 71.676
R1314 B.n184 B.n101 71.676
R1315 B.n180 B.n100 71.676
R1316 B.n176 B.n99 71.676
R1317 B.n172 B.n98 71.676
R1318 B.n608 B.n537 71.676
R1319 B.n614 B.n613 71.676
R1320 B.n617 B.n616 71.676
R1321 B.n622 B.n621 71.676
R1322 B.n625 B.n624 71.676
R1323 B.n630 B.n629 71.676
R1324 B.n633 B.n632 71.676
R1325 B.n638 B.n637 71.676
R1326 B.n641 B.n640 71.676
R1327 B.n646 B.n645 71.676
R1328 B.n649 B.n648 71.676
R1329 B.n654 B.n653 71.676
R1330 B.n657 B.n656 71.676
R1331 B.n662 B.n661 71.676
R1332 B.n665 B.n664 71.676
R1333 B.n670 B.n669 71.676
R1334 B.n673 B.n672 71.676
R1335 B.n678 B.n677 71.676
R1336 B.n681 B.n680 71.676
R1337 B.n686 B.n685 71.676
R1338 B.n689 B.n688 71.676
R1339 B.n694 B.n693 71.676
R1340 B.n697 B.n696 71.676
R1341 B.n702 B.n701 71.676
R1342 B.n705 B.n704 71.676
R1343 B.n710 B.n709 71.676
R1344 B.n713 B.n712 71.676
R1345 B.n718 B.n717 71.676
R1346 B.n721 B.n720 71.676
R1347 B.n726 B.n725 71.676
R1348 B.n729 B.n728 71.676
R1349 B.n735 B.n734 71.676
R1350 B.n738 B.n737 71.676
R1351 B.n743 B.n742 71.676
R1352 B.n746 B.n745 71.676
R1353 B.n754 B.n753 71.676
R1354 B.n757 B.n756 71.676
R1355 B.n762 B.n761 71.676
R1356 B.n765 B.n764 71.676
R1357 B.n770 B.n769 71.676
R1358 B.n773 B.n772 71.676
R1359 B.n778 B.n777 71.676
R1360 B.n781 B.n780 71.676
R1361 B.n786 B.n785 71.676
R1362 B.n789 B.n788 71.676
R1363 B.n794 B.n793 71.676
R1364 B.n797 B.n796 71.676
R1365 B.n802 B.n801 71.676
R1366 B.n805 B.n804 71.676
R1367 B.n810 B.n809 71.676
R1368 B.n813 B.n812 71.676
R1369 B.n818 B.n817 71.676
R1370 B.n821 B.n820 71.676
R1371 B.n826 B.n825 71.676
R1372 B.n829 B.n828 71.676
R1373 B.n834 B.n833 71.676
R1374 B.n837 B.n836 71.676
R1375 B.n842 B.n841 71.676
R1376 B.n845 B.n844 71.676
R1377 B.n850 B.n849 71.676
R1378 B.n853 B.n852 71.676
R1379 B.n858 B.n857 71.676
R1380 B.n861 B.n860 71.676
R1381 B.n866 B.n865 71.676
R1382 B.n869 B.n868 71.676
R1383 B.n874 B.n873 71.676
R1384 B.n877 B.n876 71.676
R1385 B.n609 B.n608 71.676
R1386 B.n615 B.n614 71.676
R1387 B.n616 B.n605 71.676
R1388 B.n623 B.n622 71.676
R1389 B.n624 B.n603 71.676
R1390 B.n631 B.n630 71.676
R1391 B.n632 B.n601 71.676
R1392 B.n639 B.n638 71.676
R1393 B.n640 B.n599 71.676
R1394 B.n647 B.n646 71.676
R1395 B.n648 B.n597 71.676
R1396 B.n655 B.n654 71.676
R1397 B.n656 B.n595 71.676
R1398 B.n663 B.n662 71.676
R1399 B.n664 B.n593 71.676
R1400 B.n671 B.n670 71.676
R1401 B.n672 B.n591 71.676
R1402 B.n679 B.n678 71.676
R1403 B.n680 B.n589 71.676
R1404 B.n687 B.n686 71.676
R1405 B.n688 B.n587 71.676
R1406 B.n695 B.n694 71.676
R1407 B.n696 B.n585 71.676
R1408 B.n703 B.n702 71.676
R1409 B.n704 B.n583 71.676
R1410 B.n711 B.n710 71.676
R1411 B.n712 B.n581 71.676
R1412 B.n719 B.n718 71.676
R1413 B.n720 B.n579 71.676
R1414 B.n727 B.n726 71.676
R1415 B.n728 B.n575 71.676
R1416 B.n736 B.n735 71.676
R1417 B.n737 B.n573 71.676
R1418 B.n744 B.n743 71.676
R1419 B.n745 B.n571 71.676
R1420 B.n755 B.n754 71.676
R1421 B.n756 B.n569 71.676
R1422 B.n763 B.n762 71.676
R1423 B.n764 B.n567 71.676
R1424 B.n771 B.n770 71.676
R1425 B.n772 B.n565 71.676
R1426 B.n779 B.n778 71.676
R1427 B.n780 B.n563 71.676
R1428 B.n787 B.n786 71.676
R1429 B.n788 B.n561 71.676
R1430 B.n795 B.n794 71.676
R1431 B.n796 B.n559 71.676
R1432 B.n803 B.n802 71.676
R1433 B.n804 B.n557 71.676
R1434 B.n811 B.n810 71.676
R1435 B.n812 B.n555 71.676
R1436 B.n819 B.n818 71.676
R1437 B.n820 B.n553 71.676
R1438 B.n827 B.n826 71.676
R1439 B.n828 B.n551 71.676
R1440 B.n835 B.n834 71.676
R1441 B.n836 B.n549 71.676
R1442 B.n843 B.n842 71.676
R1443 B.n844 B.n547 71.676
R1444 B.n851 B.n850 71.676
R1445 B.n852 B.n545 71.676
R1446 B.n859 B.n858 71.676
R1447 B.n860 B.n543 71.676
R1448 B.n867 B.n866 71.676
R1449 B.n868 B.n541 71.676
R1450 B.n875 B.n874 71.676
R1451 B.n876 B.n539 71.676
R1452 B.n1216 B.n1215 71.676
R1453 B.n1216 B.n2 71.676
R1454 B.n167 B.t11 68.5441
R1455 B.n750 B.t14 68.5441
R1456 B.n170 B.t18 68.5183
R1457 B.n577 B.t20 68.5183
R1458 B.n882 B.n538 60.8986
R1459 B.n1109 B.n1108 60.8986
R1460 B.n295 B.n170 59.5399
R1461 B.n168 B.n167 59.5399
R1462 B.n751 B.n750 59.5399
R1463 B.n732 B.n577 59.5399
R1464 B.n170 B.n169 58.7641
R1465 B.n167 B.n166 58.7641
R1466 B.n750 B.n749 58.7641
R1467 B.n577 B.n576 58.7641
R1468 B.n884 B.n536 32.3127
R1469 B.n880 B.n879 32.3127
R1470 B.n1106 B.n1105 32.3127
R1471 B.n1111 B.n95 32.3127
R1472 B.n882 B.n534 30.6751
R1473 B.n888 B.n534 30.6751
R1474 B.n888 B.n530 30.6751
R1475 B.n894 B.n530 30.6751
R1476 B.n894 B.n525 30.6751
R1477 B.n900 B.n525 30.6751
R1478 B.n900 B.n526 30.6751
R1479 B.n906 B.n518 30.6751
R1480 B.n912 B.n518 30.6751
R1481 B.n912 B.n514 30.6751
R1482 B.n918 B.n514 30.6751
R1483 B.n918 B.n510 30.6751
R1484 B.n924 B.n510 30.6751
R1485 B.n924 B.n506 30.6751
R1486 B.n930 B.n506 30.6751
R1487 B.n930 B.n501 30.6751
R1488 B.n936 B.n501 30.6751
R1489 B.n936 B.n502 30.6751
R1490 B.n942 B.n494 30.6751
R1491 B.n948 B.n494 30.6751
R1492 B.n948 B.n490 30.6751
R1493 B.n954 B.n490 30.6751
R1494 B.n954 B.n486 30.6751
R1495 B.n960 B.n486 30.6751
R1496 B.n960 B.n482 30.6751
R1497 B.n966 B.n482 30.6751
R1498 B.n972 B.n478 30.6751
R1499 B.n972 B.n474 30.6751
R1500 B.n978 B.n474 30.6751
R1501 B.n978 B.n470 30.6751
R1502 B.n984 B.n470 30.6751
R1503 B.n984 B.n466 30.6751
R1504 B.n991 B.n466 30.6751
R1505 B.n991 B.n990 30.6751
R1506 B.n997 B.n459 30.6751
R1507 B.n1003 B.n459 30.6751
R1508 B.n1003 B.n455 30.6751
R1509 B.n1009 B.n455 30.6751
R1510 B.n1009 B.n451 30.6751
R1511 B.n1015 B.n451 30.6751
R1512 B.n1015 B.n447 30.6751
R1513 B.n1021 B.n447 30.6751
R1514 B.n1028 B.n443 30.6751
R1515 B.n1028 B.n439 30.6751
R1516 B.n1034 B.n439 30.6751
R1517 B.n1034 B.n4 30.6751
R1518 B.n1214 B.n4 30.6751
R1519 B.n1214 B.n1213 30.6751
R1520 B.n1213 B.n1212 30.6751
R1521 B.n1212 B.n8 30.6751
R1522 B.n12 B.n8 30.6751
R1523 B.n1205 B.n12 30.6751
R1524 B.n1205 B.n1204 30.6751
R1525 B.n1203 B.n16 30.6751
R1526 B.n1197 B.n16 30.6751
R1527 B.n1197 B.n1196 30.6751
R1528 B.n1196 B.n1195 30.6751
R1529 B.n1195 B.n23 30.6751
R1530 B.n1189 B.n23 30.6751
R1531 B.n1189 B.n1188 30.6751
R1532 B.n1188 B.n1187 30.6751
R1533 B.n1181 B.n33 30.6751
R1534 B.n1181 B.n1180 30.6751
R1535 B.n1180 B.n1179 30.6751
R1536 B.n1179 B.n37 30.6751
R1537 B.n1173 B.n37 30.6751
R1538 B.n1173 B.n1172 30.6751
R1539 B.n1172 B.n1171 30.6751
R1540 B.n1171 B.n44 30.6751
R1541 B.n1165 B.n1164 30.6751
R1542 B.n1164 B.n1163 30.6751
R1543 B.n1163 B.n51 30.6751
R1544 B.n1157 B.n51 30.6751
R1545 B.n1157 B.n1156 30.6751
R1546 B.n1156 B.n1155 30.6751
R1547 B.n1155 B.n58 30.6751
R1548 B.n1149 B.n58 30.6751
R1549 B.n1148 B.n1147 30.6751
R1550 B.n1147 B.n65 30.6751
R1551 B.n1141 B.n65 30.6751
R1552 B.n1141 B.n1140 30.6751
R1553 B.n1140 B.n1139 30.6751
R1554 B.n1139 B.n72 30.6751
R1555 B.n1133 B.n72 30.6751
R1556 B.n1133 B.n1132 30.6751
R1557 B.n1132 B.n1131 30.6751
R1558 B.n1131 B.n79 30.6751
R1559 B.n1125 B.n79 30.6751
R1560 B.n1124 B.n1123 30.6751
R1561 B.n1123 B.n86 30.6751
R1562 B.n1117 B.n86 30.6751
R1563 B.n1117 B.n1116 30.6751
R1564 B.n1116 B.n1115 30.6751
R1565 B.n1115 B.n93 30.6751
R1566 B.n1109 B.n93 30.6751
R1567 B.n502 B.t2 21.6532
R1568 B.t6 B.n1148 21.6532
R1569 B.n966 B.t5 18.9466
R1570 B.n1165 B.t7 18.9466
R1571 B B.n1217 18.0485
R1572 B.n526 B.t13 18.0444
R1573 B.t9 B.n1124 18.0444
R1574 B.t0 B.n443 17.1422
R1575 B.n1204 B.t4 17.1422
R1576 B.n990 B.t1 16.24
R1577 B.n33 B.t3 16.24
R1578 B.n997 B.t1 14.4356
R1579 B.n1187 B.t3 14.4356
R1580 B.n1021 B.t0 13.5334
R1581 B.t4 B.n1203 13.5334
R1582 B.n906 B.t13 12.6312
R1583 B.n1125 B.t9 12.6312
R1584 B.t5 B.n478 11.729
R1585 B.t7 B.n44 11.729
R1586 B.n885 B.n884 10.6151
R1587 B.n886 B.n885 10.6151
R1588 B.n886 B.n528 10.6151
R1589 B.n896 B.n528 10.6151
R1590 B.n897 B.n896 10.6151
R1591 B.n898 B.n897 10.6151
R1592 B.n898 B.n520 10.6151
R1593 B.n908 B.n520 10.6151
R1594 B.n909 B.n908 10.6151
R1595 B.n910 B.n909 10.6151
R1596 B.n910 B.n512 10.6151
R1597 B.n920 B.n512 10.6151
R1598 B.n921 B.n920 10.6151
R1599 B.n922 B.n921 10.6151
R1600 B.n922 B.n504 10.6151
R1601 B.n932 B.n504 10.6151
R1602 B.n933 B.n932 10.6151
R1603 B.n934 B.n933 10.6151
R1604 B.n934 B.n496 10.6151
R1605 B.n944 B.n496 10.6151
R1606 B.n945 B.n944 10.6151
R1607 B.n946 B.n945 10.6151
R1608 B.n946 B.n488 10.6151
R1609 B.n956 B.n488 10.6151
R1610 B.n957 B.n956 10.6151
R1611 B.n958 B.n957 10.6151
R1612 B.n958 B.n480 10.6151
R1613 B.n968 B.n480 10.6151
R1614 B.n969 B.n968 10.6151
R1615 B.n970 B.n969 10.6151
R1616 B.n970 B.n472 10.6151
R1617 B.n980 B.n472 10.6151
R1618 B.n981 B.n980 10.6151
R1619 B.n982 B.n981 10.6151
R1620 B.n982 B.n464 10.6151
R1621 B.n993 B.n464 10.6151
R1622 B.n994 B.n993 10.6151
R1623 B.n995 B.n994 10.6151
R1624 B.n995 B.n457 10.6151
R1625 B.n1005 B.n457 10.6151
R1626 B.n1006 B.n1005 10.6151
R1627 B.n1007 B.n1006 10.6151
R1628 B.n1007 B.n449 10.6151
R1629 B.n1017 B.n449 10.6151
R1630 B.n1018 B.n1017 10.6151
R1631 B.n1019 B.n1018 10.6151
R1632 B.n1019 B.n441 10.6151
R1633 B.n1030 B.n441 10.6151
R1634 B.n1031 B.n1030 10.6151
R1635 B.n1032 B.n1031 10.6151
R1636 B.n1032 B.n0 10.6151
R1637 B.n610 B.n536 10.6151
R1638 B.n611 B.n610 10.6151
R1639 B.n612 B.n611 10.6151
R1640 B.n612 B.n606 10.6151
R1641 B.n618 B.n606 10.6151
R1642 B.n619 B.n618 10.6151
R1643 B.n620 B.n619 10.6151
R1644 B.n620 B.n604 10.6151
R1645 B.n626 B.n604 10.6151
R1646 B.n627 B.n626 10.6151
R1647 B.n628 B.n627 10.6151
R1648 B.n628 B.n602 10.6151
R1649 B.n634 B.n602 10.6151
R1650 B.n635 B.n634 10.6151
R1651 B.n636 B.n635 10.6151
R1652 B.n636 B.n600 10.6151
R1653 B.n642 B.n600 10.6151
R1654 B.n643 B.n642 10.6151
R1655 B.n644 B.n643 10.6151
R1656 B.n644 B.n598 10.6151
R1657 B.n650 B.n598 10.6151
R1658 B.n651 B.n650 10.6151
R1659 B.n652 B.n651 10.6151
R1660 B.n652 B.n596 10.6151
R1661 B.n658 B.n596 10.6151
R1662 B.n659 B.n658 10.6151
R1663 B.n660 B.n659 10.6151
R1664 B.n660 B.n594 10.6151
R1665 B.n666 B.n594 10.6151
R1666 B.n667 B.n666 10.6151
R1667 B.n668 B.n667 10.6151
R1668 B.n668 B.n592 10.6151
R1669 B.n674 B.n592 10.6151
R1670 B.n675 B.n674 10.6151
R1671 B.n676 B.n675 10.6151
R1672 B.n676 B.n590 10.6151
R1673 B.n682 B.n590 10.6151
R1674 B.n683 B.n682 10.6151
R1675 B.n684 B.n683 10.6151
R1676 B.n684 B.n588 10.6151
R1677 B.n690 B.n588 10.6151
R1678 B.n691 B.n690 10.6151
R1679 B.n692 B.n691 10.6151
R1680 B.n692 B.n586 10.6151
R1681 B.n698 B.n586 10.6151
R1682 B.n699 B.n698 10.6151
R1683 B.n700 B.n699 10.6151
R1684 B.n700 B.n584 10.6151
R1685 B.n706 B.n584 10.6151
R1686 B.n707 B.n706 10.6151
R1687 B.n708 B.n707 10.6151
R1688 B.n708 B.n582 10.6151
R1689 B.n714 B.n582 10.6151
R1690 B.n715 B.n714 10.6151
R1691 B.n716 B.n715 10.6151
R1692 B.n716 B.n580 10.6151
R1693 B.n722 B.n580 10.6151
R1694 B.n723 B.n722 10.6151
R1695 B.n724 B.n723 10.6151
R1696 B.n724 B.n578 10.6151
R1697 B.n730 B.n578 10.6151
R1698 B.n731 B.n730 10.6151
R1699 B.n733 B.n574 10.6151
R1700 B.n739 B.n574 10.6151
R1701 B.n740 B.n739 10.6151
R1702 B.n741 B.n740 10.6151
R1703 B.n741 B.n572 10.6151
R1704 B.n747 B.n572 10.6151
R1705 B.n748 B.n747 10.6151
R1706 B.n752 B.n748 10.6151
R1707 B.n758 B.n570 10.6151
R1708 B.n759 B.n758 10.6151
R1709 B.n760 B.n759 10.6151
R1710 B.n760 B.n568 10.6151
R1711 B.n766 B.n568 10.6151
R1712 B.n767 B.n766 10.6151
R1713 B.n768 B.n767 10.6151
R1714 B.n768 B.n566 10.6151
R1715 B.n774 B.n566 10.6151
R1716 B.n775 B.n774 10.6151
R1717 B.n776 B.n775 10.6151
R1718 B.n776 B.n564 10.6151
R1719 B.n782 B.n564 10.6151
R1720 B.n783 B.n782 10.6151
R1721 B.n784 B.n783 10.6151
R1722 B.n784 B.n562 10.6151
R1723 B.n790 B.n562 10.6151
R1724 B.n791 B.n790 10.6151
R1725 B.n792 B.n791 10.6151
R1726 B.n792 B.n560 10.6151
R1727 B.n798 B.n560 10.6151
R1728 B.n799 B.n798 10.6151
R1729 B.n800 B.n799 10.6151
R1730 B.n800 B.n558 10.6151
R1731 B.n806 B.n558 10.6151
R1732 B.n807 B.n806 10.6151
R1733 B.n808 B.n807 10.6151
R1734 B.n808 B.n556 10.6151
R1735 B.n814 B.n556 10.6151
R1736 B.n815 B.n814 10.6151
R1737 B.n816 B.n815 10.6151
R1738 B.n816 B.n554 10.6151
R1739 B.n822 B.n554 10.6151
R1740 B.n823 B.n822 10.6151
R1741 B.n824 B.n823 10.6151
R1742 B.n824 B.n552 10.6151
R1743 B.n830 B.n552 10.6151
R1744 B.n831 B.n830 10.6151
R1745 B.n832 B.n831 10.6151
R1746 B.n832 B.n550 10.6151
R1747 B.n838 B.n550 10.6151
R1748 B.n839 B.n838 10.6151
R1749 B.n840 B.n839 10.6151
R1750 B.n840 B.n548 10.6151
R1751 B.n846 B.n548 10.6151
R1752 B.n847 B.n846 10.6151
R1753 B.n848 B.n847 10.6151
R1754 B.n848 B.n546 10.6151
R1755 B.n854 B.n546 10.6151
R1756 B.n855 B.n854 10.6151
R1757 B.n856 B.n855 10.6151
R1758 B.n856 B.n544 10.6151
R1759 B.n862 B.n544 10.6151
R1760 B.n863 B.n862 10.6151
R1761 B.n864 B.n863 10.6151
R1762 B.n864 B.n542 10.6151
R1763 B.n870 B.n542 10.6151
R1764 B.n871 B.n870 10.6151
R1765 B.n872 B.n871 10.6151
R1766 B.n872 B.n540 10.6151
R1767 B.n878 B.n540 10.6151
R1768 B.n879 B.n878 10.6151
R1769 B.n880 B.n532 10.6151
R1770 B.n890 B.n532 10.6151
R1771 B.n891 B.n890 10.6151
R1772 B.n892 B.n891 10.6151
R1773 B.n892 B.n523 10.6151
R1774 B.n902 B.n523 10.6151
R1775 B.n903 B.n902 10.6151
R1776 B.n904 B.n903 10.6151
R1777 B.n904 B.n516 10.6151
R1778 B.n914 B.n516 10.6151
R1779 B.n915 B.n914 10.6151
R1780 B.n916 B.n915 10.6151
R1781 B.n916 B.n508 10.6151
R1782 B.n926 B.n508 10.6151
R1783 B.n927 B.n926 10.6151
R1784 B.n928 B.n927 10.6151
R1785 B.n928 B.n499 10.6151
R1786 B.n938 B.n499 10.6151
R1787 B.n939 B.n938 10.6151
R1788 B.n940 B.n939 10.6151
R1789 B.n940 B.n492 10.6151
R1790 B.n950 B.n492 10.6151
R1791 B.n951 B.n950 10.6151
R1792 B.n952 B.n951 10.6151
R1793 B.n952 B.n484 10.6151
R1794 B.n962 B.n484 10.6151
R1795 B.n963 B.n962 10.6151
R1796 B.n964 B.n963 10.6151
R1797 B.n964 B.n476 10.6151
R1798 B.n974 B.n476 10.6151
R1799 B.n975 B.n974 10.6151
R1800 B.n976 B.n975 10.6151
R1801 B.n976 B.n468 10.6151
R1802 B.n986 B.n468 10.6151
R1803 B.n987 B.n986 10.6151
R1804 B.n988 B.n987 10.6151
R1805 B.n988 B.n461 10.6151
R1806 B.n999 B.n461 10.6151
R1807 B.n1000 B.n999 10.6151
R1808 B.n1001 B.n1000 10.6151
R1809 B.n1001 B.n453 10.6151
R1810 B.n1011 B.n453 10.6151
R1811 B.n1012 B.n1011 10.6151
R1812 B.n1013 B.n1012 10.6151
R1813 B.n1013 B.n445 10.6151
R1814 B.n1023 B.n445 10.6151
R1815 B.n1024 B.n1023 10.6151
R1816 B.n1026 B.n1024 10.6151
R1817 B.n1026 B.n1025 10.6151
R1818 B.n1025 B.n437 10.6151
R1819 B.n1037 B.n437 10.6151
R1820 B.n1038 B.n1037 10.6151
R1821 B.n1039 B.n1038 10.6151
R1822 B.n1040 B.n1039 10.6151
R1823 B.n1041 B.n1040 10.6151
R1824 B.n1044 B.n1041 10.6151
R1825 B.n1045 B.n1044 10.6151
R1826 B.n1046 B.n1045 10.6151
R1827 B.n1047 B.n1046 10.6151
R1828 B.n1049 B.n1047 10.6151
R1829 B.n1050 B.n1049 10.6151
R1830 B.n1051 B.n1050 10.6151
R1831 B.n1052 B.n1051 10.6151
R1832 B.n1054 B.n1052 10.6151
R1833 B.n1055 B.n1054 10.6151
R1834 B.n1056 B.n1055 10.6151
R1835 B.n1057 B.n1056 10.6151
R1836 B.n1059 B.n1057 10.6151
R1837 B.n1060 B.n1059 10.6151
R1838 B.n1061 B.n1060 10.6151
R1839 B.n1062 B.n1061 10.6151
R1840 B.n1064 B.n1062 10.6151
R1841 B.n1065 B.n1064 10.6151
R1842 B.n1066 B.n1065 10.6151
R1843 B.n1067 B.n1066 10.6151
R1844 B.n1069 B.n1067 10.6151
R1845 B.n1070 B.n1069 10.6151
R1846 B.n1071 B.n1070 10.6151
R1847 B.n1072 B.n1071 10.6151
R1848 B.n1074 B.n1072 10.6151
R1849 B.n1075 B.n1074 10.6151
R1850 B.n1076 B.n1075 10.6151
R1851 B.n1077 B.n1076 10.6151
R1852 B.n1079 B.n1077 10.6151
R1853 B.n1080 B.n1079 10.6151
R1854 B.n1081 B.n1080 10.6151
R1855 B.n1082 B.n1081 10.6151
R1856 B.n1084 B.n1082 10.6151
R1857 B.n1085 B.n1084 10.6151
R1858 B.n1086 B.n1085 10.6151
R1859 B.n1087 B.n1086 10.6151
R1860 B.n1089 B.n1087 10.6151
R1861 B.n1090 B.n1089 10.6151
R1862 B.n1091 B.n1090 10.6151
R1863 B.n1092 B.n1091 10.6151
R1864 B.n1094 B.n1092 10.6151
R1865 B.n1095 B.n1094 10.6151
R1866 B.n1096 B.n1095 10.6151
R1867 B.n1097 B.n1096 10.6151
R1868 B.n1099 B.n1097 10.6151
R1869 B.n1100 B.n1099 10.6151
R1870 B.n1101 B.n1100 10.6151
R1871 B.n1102 B.n1101 10.6151
R1872 B.n1104 B.n1102 10.6151
R1873 B.n1105 B.n1104 10.6151
R1874 B.n1209 B.n1 10.6151
R1875 B.n1209 B.n1208 10.6151
R1876 B.n1208 B.n1207 10.6151
R1877 B.n1207 B.n10 10.6151
R1878 B.n1201 B.n10 10.6151
R1879 B.n1201 B.n1200 10.6151
R1880 B.n1200 B.n1199 10.6151
R1881 B.n1199 B.n18 10.6151
R1882 B.n1193 B.n18 10.6151
R1883 B.n1193 B.n1192 10.6151
R1884 B.n1192 B.n1191 10.6151
R1885 B.n1191 B.n25 10.6151
R1886 B.n1185 B.n25 10.6151
R1887 B.n1185 B.n1184 10.6151
R1888 B.n1184 B.n1183 10.6151
R1889 B.n1183 B.n31 10.6151
R1890 B.n1177 B.n31 10.6151
R1891 B.n1177 B.n1176 10.6151
R1892 B.n1176 B.n1175 10.6151
R1893 B.n1175 B.n39 10.6151
R1894 B.n1169 B.n39 10.6151
R1895 B.n1169 B.n1168 10.6151
R1896 B.n1168 B.n1167 10.6151
R1897 B.n1167 B.n46 10.6151
R1898 B.n1161 B.n46 10.6151
R1899 B.n1161 B.n1160 10.6151
R1900 B.n1160 B.n1159 10.6151
R1901 B.n1159 B.n53 10.6151
R1902 B.n1153 B.n53 10.6151
R1903 B.n1153 B.n1152 10.6151
R1904 B.n1152 B.n1151 10.6151
R1905 B.n1151 B.n60 10.6151
R1906 B.n1145 B.n60 10.6151
R1907 B.n1145 B.n1144 10.6151
R1908 B.n1144 B.n1143 10.6151
R1909 B.n1143 B.n67 10.6151
R1910 B.n1137 B.n67 10.6151
R1911 B.n1137 B.n1136 10.6151
R1912 B.n1136 B.n1135 10.6151
R1913 B.n1135 B.n74 10.6151
R1914 B.n1129 B.n74 10.6151
R1915 B.n1129 B.n1128 10.6151
R1916 B.n1128 B.n1127 10.6151
R1917 B.n1127 B.n81 10.6151
R1918 B.n1121 B.n81 10.6151
R1919 B.n1121 B.n1120 10.6151
R1920 B.n1120 B.n1119 10.6151
R1921 B.n1119 B.n88 10.6151
R1922 B.n1113 B.n88 10.6151
R1923 B.n1113 B.n1112 10.6151
R1924 B.n1112 B.n1111 10.6151
R1925 B.n171 B.n95 10.6151
R1926 B.n174 B.n171 10.6151
R1927 B.n175 B.n174 10.6151
R1928 B.n178 B.n175 10.6151
R1929 B.n179 B.n178 10.6151
R1930 B.n182 B.n179 10.6151
R1931 B.n183 B.n182 10.6151
R1932 B.n186 B.n183 10.6151
R1933 B.n187 B.n186 10.6151
R1934 B.n190 B.n187 10.6151
R1935 B.n191 B.n190 10.6151
R1936 B.n194 B.n191 10.6151
R1937 B.n195 B.n194 10.6151
R1938 B.n198 B.n195 10.6151
R1939 B.n199 B.n198 10.6151
R1940 B.n202 B.n199 10.6151
R1941 B.n203 B.n202 10.6151
R1942 B.n206 B.n203 10.6151
R1943 B.n207 B.n206 10.6151
R1944 B.n210 B.n207 10.6151
R1945 B.n211 B.n210 10.6151
R1946 B.n214 B.n211 10.6151
R1947 B.n215 B.n214 10.6151
R1948 B.n218 B.n215 10.6151
R1949 B.n219 B.n218 10.6151
R1950 B.n222 B.n219 10.6151
R1951 B.n223 B.n222 10.6151
R1952 B.n226 B.n223 10.6151
R1953 B.n227 B.n226 10.6151
R1954 B.n230 B.n227 10.6151
R1955 B.n231 B.n230 10.6151
R1956 B.n234 B.n231 10.6151
R1957 B.n235 B.n234 10.6151
R1958 B.n238 B.n235 10.6151
R1959 B.n239 B.n238 10.6151
R1960 B.n242 B.n239 10.6151
R1961 B.n243 B.n242 10.6151
R1962 B.n246 B.n243 10.6151
R1963 B.n247 B.n246 10.6151
R1964 B.n250 B.n247 10.6151
R1965 B.n251 B.n250 10.6151
R1966 B.n254 B.n251 10.6151
R1967 B.n255 B.n254 10.6151
R1968 B.n258 B.n255 10.6151
R1969 B.n259 B.n258 10.6151
R1970 B.n262 B.n259 10.6151
R1971 B.n263 B.n262 10.6151
R1972 B.n266 B.n263 10.6151
R1973 B.n267 B.n266 10.6151
R1974 B.n270 B.n267 10.6151
R1975 B.n271 B.n270 10.6151
R1976 B.n274 B.n271 10.6151
R1977 B.n275 B.n274 10.6151
R1978 B.n278 B.n275 10.6151
R1979 B.n279 B.n278 10.6151
R1980 B.n282 B.n279 10.6151
R1981 B.n283 B.n282 10.6151
R1982 B.n286 B.n283 10.6151
R1983 B.n287 B.n286 10.6151
R1984 B.n290 B.n287 10.6151
R1985 B.n291 B.n290 10.6151
R1986 B.n294 B.n291 10.6151
R1987 B.n299 B.n296 10.6151
R1988 B.n300 B.n299 10.6151
R1989 B.n303 B.n300 10.6151
R1990 B.n304 B.n303 10.6151
R1991 B.n307 B.n304 10.6151
R1992 B.n308 B.n307 10.6151
R1993 B.n311 B.n308 10.6151
R1994 B.n312 B.n311 10.6151
R1995 B.n316 B.n315 10.6151
R1996 B.n319 B.n316 10.6151
R1997 B.n320 B.n319 10.6151
R1998 B.n323 B.n320 10.6151
R1999 B.n324 B.n323 10.6151
R2000 B.n327 B.n324 10.6151
R2001 B.n328 B.n327 10.6151
R2002 B.n331 B.n328 10.6151
R2003 B.n332 B.n331 10.6151
R2004 B.n335 B.n332 10.6151
R2005 B.n336 B.n335 10.6151
R2006 B.n339 B.n336 10.6151
R2007 B.n340 B.n339 10.6151
R2008 B.n343 B.n340 10.6151
R2009 B.n344 B.n343 10.6151
R2010 B.n347 B.n344 10.6151
R2011 B.n348 B.n347 10.6151
R2012 B.n351 B.n348 10.6151
R2013 B.n352 B.n351 10.6151
R2014 B.n355 B.n352 10.6151
R2015 B.n356 B.n355 10.6151
R2016 B.n359 B.n356 10.6151
R2017 B.n360 B.n359 10.6151
R2018 B.n363 B.n360 10.6151
R2019 B.n364 B.n363 10.6151
R2020 B.n367 B.n364 10.6151
R2021 B.n368 B.n367 10.6151
R2022 B.n371 B.n368 10.6151
R2023 B.n372 B.n371 10.6151
R2024 B.n375 B.n372 10.6151
R2025 B.n376 B.n375 10.6151
R2026 B.n379 B.n376 10.6151
R2027 B.n380 B.n379 10.6151
R2028 B.n383 B.n380 10.6151
R2029 B.n384 B.n383 10.6151
R2030 B.n387 B.n384 10.6151
R2031 B.n388 B.n387 10.6151
R2032 B.n391 B.n388 10.6151
R2033 B.n392 B.n391 10.6151
R2034 B.n395 B.n392 10.6151
R2035 B.n396 B.n395 10.6151
R2036 B.n399 B.n396 10.6151
R2037 B.n400 B.n399 10.6151
R2038 B.n403 B.n400 10.6151
R2039 B.n404 B.n403 10.6151
R2040 B.n407 B.n404 10.6151
R2041 B.n408 B.n407 10.6151
R2042 B.n411 B.n408 10.6151
R2043 B.n412 B.n411 10.6151
R2044 B.n415 B.n412 10.6151
R2045 B.n416 B.n415 10.6151
R2046 B.n419 B.n416 10.6151
R2047 B.n420 B.n419 10.6151
R2048 B.n423 B.n420 10.6151
R2049 B.n424 B.n423 10.6151
R2050 B.n427 B.n424 10.6151
R2051 B.n428 B.n427 10.6151
R2052 B.n431 B.n428 10.6151
R2053 B.n432 B.n431 10.6151
R2054 B.n435 B.n432 10.6151
R2055 B.n436 B.n435 10.6151
R2056 B.n1106 B.n436 10.6151
R2057 B.n942 B.t2 9.02244
R2058 B.n1149 B.t6 9.02244
R2059 B.n1217 B.n0 8.11757
R2060 B.n1217 B.n1 8.11757
R2061 B.n733 B.n732 6.5566
R2062 B.n752 B.n751 6.5566
R2063 B.n296 B.n295 6.5566
R2064 B.n312 B.n168 6.5566
R2065 B.n732 B.n731 4.05904
R2066 B.n751 B.n570 4.05904
R2067 B.n295 B.n294 4.05904
R2068 B.n315 B.n168 4.05904
R2069 VP.n19 VP.t7 201.38
R2070 VP.n43 VP.t6 170.575
R2071 VP.n7 VP.t2 170.575
R2072 VP.n3 VP.t0 170.575
R2073 VP.n73 VP.t5 170.575
R2074 VP.n40 VP.t4 170.575
R2075 VP.n14 VP.t3 170.575
R2076 VP.n18 VP.t1 170.575
R2077 VP.n21 VP.n20 161.3
R2078 VP.n22 VP.n17 161.3
R2079 VP.n24 VP.n23 161.3
R2080 VP.n25 VP.n16 161.3
R2081 VP.n27 VP.n26 161.3
R2082 VP.n28 VP.n15 161.3
R2083 VP.n30 VP.n29 161.3
R2084 VP.n32 VP.n31 161.3
R2085 VP.n33 VP.n13 161.3
R2086 VP.n35 VP.n34 161.3
R2087 VP.n36 VP.n12 161.3
R2088 VP.n38 VP.n37 161.3
R2089 VP.n39 VP.n11 161.3
R2090 VP.n72 VP.n0 161.3
R2091 VP.n71 VP.n70 161.3
R2092 VP.n69 VP.n1 161.3
R2093 VP.n68 VP.n67 161.3
R2094 VP.n66 VP.n2 161.3
R2095 VP.n65 VP.n64 161.3
R2096 VP.n63 VP.n62 161.3
R2097 VP.n61 VP.n4 161.3
R2098 VP.n60 VP.n59 161.3
R2099 VP.n58 VP.n5 161.3
R2100 VP.n57 VP.n56 161.3
R2101 VP.n55 VP.n6 161.3
R2102 VP.n54 VP.n53 161.3
R2103 VP.n52 VP.n51 161.3
R2104 VP.n50 VP.n8 161.3
R2105 VP.n49 VP.n48 161.3
R2106 VP.n47 VP.n9 161.3
R2107 VP.n46 VP.n45 161.3
R2108 VP.n44 VP.n10 161.3
R2109 VP.n43 VP.n42 108.555
R2110 VP.n74 VP.n73 108.555
R2111 VP.n41 VP.n40 108.555
R2112 VP.n19 VP.n18 72.6301
R2113 VP.n42 VP.n41 56.6738
R2114 VP.n49 VP.n9 43.4072
R2115 VP.n67 VP.n1 43.4072
R2116 VP.n34 VP.n12 43.4072
R2117 VP.n56 VP.n5 40.4934
R2118 VP.n60 VP.n5 40.4934
R2119 VP.n27 VP.n16 40.4934
R2120 VP.n23 VP.n16 40.4934
R2121 VP.n50 VP.n49 37.5796
R2122 VP.n67 VP.n66 37.5796
R2123 VP.n34 VP.n33 37.5796
R2124 VP.n45 VP.n44 24.4675
R2125 VP.n45 VP.n9 24.4675
R2126 VP.n51 VP.n50 24.4675
R2127 VP.n55 VP.n54 24.4675
R2128 VP.n56 VP.n55 24.4675
R2129 VP.n61 VP.n60 24.4675
R2130 VP.n62 VP.n61 24.4675
R2131 VP.n66 VP.n65 24.4675
R2132 VP.n71 VP.n1 24.4675
R2133 VP.n72 VP.n71 24.4675
R2134 VP.n38 VP.n12 24.4675
R2135 VP.n39 VP.n38 24.4675
R2136 VP.n28 VP.n27 24.4675
R2137 VP.n29 VP.n28 24.4675
R2138 VP.n33 VP.n32 24.4675
R2139 VP.n22 VP.n21 24.4675
R2140 VP.n23 VP.n22 24.4675
R2141 VP.n51 VP.n7 23.7335
R2142 VP.n65 VP.n3 23.7335
R2143 VP.n32 VP.n14 23.7335
R2144 VP.n20 VP.n19 7.35942
R2145 VP.n44 VP.n43 2.20253
R2146 VP.n73 VP.n72 2.20253
R2147 VP.n40 VP.n39 2.20253
R2148 VP.n54 VP.n7 0.73451
R2149 VP.n62 VP.n3 0.73451
R2150 VP.n29 VP.n14 0.73451
R2151 VP.n21 VP.n18 0.73451
R2152 VP.n41 VP.n11 0.278367
R2153 VP.n42 VP.n10 0.278367
R2154 VP.n74 VP.n0 0.278367
R2155 VP.n20 VP.n17 0.189894
R2156 VP.n24 VP.n17 0.189894
R2157 VP.n25 VP.n24 0.189894
R2158 VP.n26 VP.n25 0.189894
R2159 VP.n26 VP.n15 0.189894
R2160 VP.n30 VP.n15 0.189894
R2161 VP.n31 VP.n30 0.189894
R2162 VP.n31 VP.n13 0.189894
R2163 VP.n35 VP.n13 0.189894
R2164 VP.n36 VP.n35 0.189894
R2165 VP.n37 VP.n36 0.189894
R2166 VP.n37 VP.n11 0.189894
R2167 VP.n46 VP.n10 0.189894
R2168 VP.n47 VP.n46 0.189894
R2169 VP.n48 VP.n47 0.189894
R2170 VP.n48 VP.n8 0.189894
R2171 VP.n52 VP.n8 0.189894
R2172 VP.n53 VP.n52 0.189894
R2173 VP.n53 VP.n6 0.189894
R2174 VP.n57 VP.n6 0.189894
R2175 VP.n58 VP.n57 0.189894
R2176 VP.n59 VP.n58 0.189894
R2177 VP.n59 VP.n4 0.189894
R2178 VP.n63 VP.n4 0.189894
R2179 VP.n64 VP.n63 0.189894
R2180 VP.n64 VP.n2 0.189894
R2181 VP.n68 VP.n2 0.189894
R2182 VP.n69 VP.n68 0.189894
R2183 VP.n70 VP.n69 0.189894
R2184 VP.n70 VP.n0 0.189894
R2185 VP VP.n74 0.153454
R2186 VDD1 VDD1.n0 64.4729
R2187 VDD1.n3 VDD1.n2 64.3581
R2188 VDD1.n3 VDD1.n1 64.3581
R2189 VDD1.n5 VDD1.n4 63.1085
R2190 VDD1.n5 VDD1.n3 52.5268
R2191 VDD1 VDD1.n5 1.24834
R2192 VDD1.n4 VDD1.t0 1.03661
R2193 VDD1.n4 VDD1.t5 1.03661
R2194 VDD1.n0 VDD1.t6 1.03661
R2195 VDD1.n0 VDD1.t2 1.03661
R2196 VDD1.n2 VDD1.t4 1.03661
R2197 VDD1.n2 VDD1.t3 1.03661
R2198 VDD1.n1 VDD1.t7 1.03661
R2199 VDD1.n1 VDD1.t1 1.03661
R2200 VTAIL.n11 VTAIL.t7 47.4659
R2201 VTAIL.n10 VTAIL.t0 47.4659
R2202 VTAIL.n7 VTAIL.t2 47.4659
R2203 VTAIL.n15 VTAIL.t6 47.4658
R2204 VTAIL.n2 VTAIL.t4 47.4658
R2205 VTAIL.n3 VTAIL.t9 47.4658
R2206 VTAIL.n6 VTAIL.t8 47.4658
R2207 VTAIL.n14 VTAIL.t10 47.4658
R2208 VTAIL.n13 VTAIL.n12 46.4298
R2209 VTAIL.n9 VTAIL.n8 46.4298
R2210 VTAIL.n1 VTAIL.n0 46.4287
R2211 VTAIL.n5 VTAIL.n4 46.4287
R2212 VTAIL.n15 VTAIL.n14 31.4531
R2213 VTAIL.n7 VTAIL.n6 31.4531
R2214 VTAIL.n9 VTAIL.n7 2.61257
R2215 VTAIL.n10 VTAIL.n9 2.61257
R2216 VTAIL.n13 VTAIL.n11 2.61257
R2217 VTAIL.n14 VTAIL.n13 2.61257
R2218 VTAIL.n6 VTAIL.n5 2.61257
R2219 VTAIL.n5 VTAIL.n3 2.61257
R2220 VTAIL.n2 VTAIL.n1 2.61257
R2221 VTAIL VTAIL.n15 2.55438
R2222 VTAIL.n0 VTAIL.t3 1.03661
R2223 VTAIL.n0 VTAIL.t15 1.03661
R2224 VTAIL.n4 VTAIL.t12 1.03661
R2225 VTAIL.n4 VTAIL.t14 1.03661
R2226 VTAIL.n12 VTAIL.t13 1.03661
R2227 VTAIL.n12 VTAIL.t11 1.03661
R2228 VTAIL.n8 VTAIL.t5 1.03661
R2229 VTAIL.n8 VTAIL.t1 1.03661
R2230 VTAIL.n11 VTAIL.n10 0.470328
R2231 VTAIL.n3 VTAIL.n2 0.470328
R2232 VTAIL VTAIL.n1 0.0586897
R2233 VN.n8 VN.t1 201.38
R2234 VN.n39 VN.t4 201.38
R2235 VN.n7 VN.t7 170.575
R2236 VN.n3 VN.t2 170.575
R2237 VN.n29 VN.t6 170.575
R2238 VN.n38 VN.t5 170.575
R2239 VN.n34 VN.t0 170.575
R2240 VN.n60 VN.t3 170.575
R2241 VN.n59 VN.n31 161.3
R2242 VN.n58 VN.n57 161.3
R2243 VN.n56 VN.n32 161.3
R2244 VN.n55 VN.n54 161.3
R2245 VN.n53 VN.n33 161.3
R2246 VN.n52 VN.n51 161.3
R2247 VN.n50 VN.n49 161.3
R2248 VN.n48 VN.n35 161.3
R2249 VN.n47 VN.n46 161.3
R2250 VN.n45 VN.n36 161.3
R2251 VN.n44 VN.n43 161.3
R2252 VN.n42 VN.n37 161.3
R2253 VN.n41 VN.n40 161.3
R2254 VN.n28 VN.n0 161.3
R2255 VN.n27 VN.n26 161.3
R2256 VN.n25 VN.n1 161.3
R2257 VN.n24 VN.n23 161.3
R2258 VN.n22 VN.n2 161.3
R2259 VN.n21 VN.n20 161.3
R2260 VN.n19 VN.n18 161.3
R2261 VN.n17 VN.n4 161.3
R2262 VN.n16 VN.n15 161.3
R2263 VN.n14 VN.n5 161.3
R2264 VN.n13 VN.n12 161.3
R2265 VN.n11 VN.n6 161.3
R2266 VN.n10 VN.n9 161.3
R2267 VN.n30 VN.n29 108.555
R2268 VN.n61 VN.n60 108.555
R2269 VN.n8 VN.n7 72.6301
R2270 VN.n39 VN.n38 72.6301
R2271 VN VN.n61 56.9527
R2272 VN.n23 VN.n1 43.4072
R2273 VN.n54 VN.n32 43.4072
R2274 VN.n12 VN.n5 40.4934
R2275 VN.n16 VN.n5 40.4934
R2276 VN.n43 VN.n36 40.4934
R2277 VN.n47 VN.n36 40.4934
R2278 VN.n23 VN.n22 37.5796
R2279 VN.n54 VN.n53 37.5796
R2280 VN.n11 VN.n10 24.4675
R2281 VN.n12 VN.n11 24.4675
R2282 VN.n17 VN.n16 24.4675
R2283 VN.n18 VN.n17 24.4675
R2284 VN.n22 VN.n21 24.4675
R2285 VN.n27 VN.n1 24.4675
R2286 VN.n28 VN.n27 24.4675
R2287 VN.n43 VN.n42 24.4675
R2288 VN.n42 VN.n41 24.4675
R2289 VN.n53 VN.n52 24.4675
R2290 VN.n49 VN.n48 24.4675
R2291 VN.n48 VN.n47 24.4675
R2292 VN.n59 VN.n58 24.4675
R2293 VN.n58 VN.n32 24.4675
R2294 VN.n21 VN.n3 23.7335
R2295 VN.n52 VN.n34 23.7335
R2296 VN.n40 VN.n39 7.35942
R2297 VN.n9 VN.n8 7.35942
R2298 VN.n29 VN.n28 2.20253
R2299 VN.n60 VN.n59 2.20253
R2300 VN.n10 VN.n7 0.73451
R2301 VN.n18 VN.n3 0.73451
R2302 VN.n41 VN.n38 0.73451
R2303 VN.n49 VN.n34 0.73451
R2304 VN.n61 VN.n31 0.278367
R2305 VN.n30 VN.n0 0.278367
R2306 VN.n57 VN.n31 0.189894
R2307 VN.n57 VN.n56 0.189894
R2308 VN.n56 VN.n55 0.189894
R2309 VN.n55 VN.n33 0.189894
R2310 VN.n51 VN.n33 0.189894
R2311 VN.n51 VN.n50 0.189894
R2312 VN.n50 VN.n35 0.189894
R2313 VN.n46 VN.n35 0.189894
R2314 VN.n46 VN.n45 0.189894
R2315 VN.n45 VN.n44 0.189894
R2316 VN.n44 VN.n37 0.189894
R2317 VN.n40 VN.n37 0.189894
R2318 VN.n9 VN.n6 0.189894
R2319 VN.n13 VN.n6 0.189894
R2320 VN.n14 VN.n13 0.189894
R2321 VN.n15 VN.n14 0.189894
R2322 VN.n15 VN.n4 0.189894
R2323 VN.n19 VN.n4 0.189894
R2324 VN.n20 VN.n19 0.189894
R2325 VN.n20 VN.n2 0.189894
R2326 VN.n24 VN.n2 0.189894
R2327 VN.n25 VN.n24 0.189894
R2328 VN.n26 VN.n25 0.189894
R2329 VN.n26 VN.n0 0.189894
R2330 VN VN.n30 0.153454
R2331 VDD2.n2 VDD2.n1 64.3581
R2332 VDD2.n2 VDD2.n0 64.3581
R2333 VDD2 VDD2.n5 64.3563
R2334 VDD2.n4 VDD2.n3 63.1086
R2335 VDD2.n4 VDD2.n2 51.9437
R2336 VDD2 VDD2.n4 1.36472
R2337 VDD2.n5 VDD2.t2 1.03661
R2338 VDD2.n5 VDD2.t3 1.03661
R2339 VDD2.n3 VDD2.t4 1.03661
R2340 VDD2.n3 VDD2.t7 1.03661
R2341 VDD2.n1 VDD2.t5 1.03661
R2342 VDD2.n1 VDD2.t1 1.03661
R2343 VDD2.n0 VDD2.t6 1.03661
R2344 VDD2.n0 VDD2.t0 1.03661
C0 VP VDD1 14.064599f
C1 VTAIL VDD2 10.498099f
C2 VDD2 VN 13.687599f
C3 VTAIL VN 13.793f
C4 VDD2 VDD1 1.82674f
C5 VP VDD2 0.529926f
C6 VTAIL VDD1 10.443f
C7 VTAIL VP 13.807099f
C8 VDD1 VN 0.151523f
C9 VP VN 9.10405f
C10 VDD2 B 5.978796f
C11 VDD1 B 6.423375f
C12 VTAIL B 14.81352f
C13 VN B 16.48973f
C14 VP B 14.968886f
C15 VDD2.t6 B 0.367116f
C16 VDD2.t0 B 0.367116f
C17 VDD2.n0 B 3.37016f
C18 VDD2.t5 B 0.367116f
C19 VDD2.t1 B 0.367116f
C20 VDD2.n1 B 3.37016f
C21 VDD2.n2 B 3.67166f
C22 VDD2.t4 B 0.367116f
C23 VDD2.t7 B 0.367116f
C24 VDD2.n3 B 3.3603f
C25 VDD2.n4 B 3.41902f
C26 VDD2.t2 B 0.367116f
C27 VDD2.t3 B 0.367116f
C28 VDD2.n5 B 3.37011f
C29 VN.n0 B 0.027086f
C30 VN.t6 B 2.91888f
C31 VN.n1 B 0.040103f
C32 VN.n2 B 0.020544f
C33 VN.t2 B 2.91888f
C34 VN.n3 B 1.00913f
C35 VN.n4 B 0.020544f
C36 VN.n5 B 0.016608f
C37 VN.n6 B 0.020544f
C38 VN.t7 B 2.91888f
C39 VN.n7 B 1.06263f
C40 VN.t1 B 3.09279f
C41 VN.n8 B 1.05119f
C42 VN.n9 B 0.20032f
C43 VN.n10 B 0.019952f
C44 VN.n11 B 0.03829f
C45 VN.n12 B 0.040832f
C46 VN.n13 B 0.020544f
C47 VN.n14 B 0.020544f
C48 VN.n15 B 0.020544f
C49 VN.n16 B 0.040832f
C50 VN.n17 B 0.03829f
C51 VN.n18 B 0.019952f
C52 VN.n19 B 0.020544f
C53 VN.n20 B 0.020544f
C54 VN.n21 B 0.037721f
C55 VN.n22 B 0.041322f
C56 VN.n23 B 0.016847f
C57 VN.n24 B 0.020544f
C58 VN.n25 B 0.020544f
C59 VN.n26 B 0.020544f
C60 VN.n27 B 0.03829f
C61 VN.n28 B 0.021086f
C62 VN.n29 B 1.07221f
C63 VN.n30 B 0.037771f
C64 VN.n31 B 0.027086f
C65 VN.t3 B 2.91888f
C66 VN.n32 B 0.040103f
C67 VN.n33 B 0.020544f
C68 VN.t0 B 2.91888f
C69 VN.n34 B 1.00913f
C70 VN.n35 B 0.020544f
C71 VN.n36 B 0.016608f
C72 VN.n37 B 0.020544f
C73 VN.t5 B 2.91888f
C74 VN.n38 B 1.06263f
C75 VN.t4 B 3.09279f
C76 VN.n39 B 1.05119f
C77 VN.n40 B 0.20032f
C78 VN.n41 B 0.019952f
C79 VN.n42 B 0.03829f
C80 VN.n43 B 0.040832f
C81 VN.n44 B 0.020544f
C82 VN.n45 B 0.020544f
C83 VN.n46 B 0.020544f
C84 VN.n47 B 0.040832f
C85 VN.n48 B 0.03829f
C86 VN.n49 B 0.019952f
C87 VN.n50 B 0.020544f
C88 VN.n51 B 0.020544f
C89 VN.n52 B 0.037721f
C90 VN.n53 B 0.041322f
C91 VN.n54 B 0.016847f
C92 VN.n55 B 0.020544f
C93 VN.n56 B 0.020544f
C94 VN.n57 B 0.020544f
C95 VN.n58 B 0.03829f
C96 VN.n59 B 0.021086f
C97 VN.n60 B 1.07221f
C98 VN.n61 B 1.38176f
C99 VTAIL.t3 B 0.278498f
C100 VTAIL.t15 B 0.278498f
C101 VTAIL.n0 B 2.49735f
C102 VTAIL.n1 B 0.333143f
C103 VTAIL.t4 B 3.19186f
C104 VTAIL.n2 B 0.42263f
C105 VTAIL.t9 B 3.19186f
C106 VTAIL.n3 B 0.42263f
C107 VTAIL.t12 B 0.278498f
C108 VTAIL.t14 B 0.278498f
C109 VTAIL.n4 B 2.49735f
C110 VTAIL.n5 B 0.484905f
C111 VTAIL.t8 B 3.19186f
C112 VTAIL.n6 B 1.77941f
C113 VTAIL.t2 B 3.19188f
C114 VTAIL.n7 B 1.77938f
C115 VTAIL.t5 B 0.278498f
C116 VTAIL.t1 B 0.278498f
C117 VTAIL.n8 B 2.49735f
C118 VTAIL.n9 B 0.484898f
C119 VTAIL.t0 B 3.19188f
C120 VTAIL.n10 B 0.422607f
C121 VTAIL.t7 B 3.19188f
C122 VTAIL.n11 B 0.422607f
C123 VTAIL.t13 B 0.278498f
C124 VTAIL.t11 B 0.278498f
C125 VTAIL.n12 B 2.49735f
C126 VTAIL.n13 B 0.484898f
C127 VTAIL.t10 B 3.19186f
C128 VTAIL.n14 B 1.77941f
C129 VTAIL.t6 B 3.19186f
C130 VTAIL.n15 B 1.77595f
C131 VDD1.t6 B 0.370293f
C132 VDD1.t2 B 0.370293f
C133 VDD1.n0 B 3.40039f
C134 VDD1.t7 B 0.370293f
C135 VDD1.t1 B 0.370293f
C136 VDD1.n1 B 3.39932f
C137 VDD1.t4 B 0.370293f
C138 VDD1.t3 B 0.370293f
C139 VDD1.n2 B 3.39932f
C140 VDD1.n3 B 3.75416f
C141 VDD1.t0 B 0.370293f
C142 VDD1.t5 B 0.370293f
C143 VDD1.n4 B 3.38936f
C144 VDD1.n5 B 3.47927f
C145 VP.n0 B 0.027403f
C146 VP.t5 B 2.95311f
C147 VP.n1 B 0.040573f
C148 VP.n2 B 0.020785f
C149 VP.t0 B 2.95311f
C150 VP.n3 B 1.02097f
C151 VP.n4 B 0.020785f
C152 VP.n5 B 0.016803f
C153 VP.n6 B 0.020785f
C154 VP.t2 B 2.95311f
C155 VP.n7 B 1.02097f
C156 VP.n8 B 0.020785f
C157 VP.n9 B 0.040573f
C158 VP.n10 B 0.027403f
C159 VP.t6 B 2.95311f
C160 VP.n11 B 0.027403f
C161 VP.t4 B 2.95311f
C162 VP.n12 B 0.040573f
C163 VP.n13 B 0.020785f
C164 VP.t3 B 2.95311f
C165 VP.n14 B 1.02097f
C166 VP.n15 B 0.020785f
C167 VP.n16 B 0.016803f
C168 VP.n17 B 0.020785f
C169 VP.t1 B 2.95311f
C170 VP.n18 B 1.07509f
C171 VP.t7 B 3.12906f
C172 VP.n19 B 1.06351f
C173 VP.n20 B 0.202669f
C174 VP.n21 B 0.020186f
C175 VP.n22 B 0.038739f
C176 VP.n23 B 0.041311f
C177 VP.n24 B 0.020785f
C178 VP.n25 B 0.020785f
C179 VP.n26 B 0.020785f
C180 VP.n27 B 0.041311f
C181 VP.n28 B 0.038739f
C182 VP.n29 B 0.020186f
C183 VP.n30 B 0.020785f
C184 VP.n31 B 0.020785f
C185 VP.n32 B 0.038164f
C186 VP.n33 B 0.041807f
C187 VP.n34 B 0.017044f
C188 VP.n35 B 0.020785f
C189 VP.n36 B 0.020785f
C190 VP.n37 B 0.020785f
C191 VP.n38 B 0.038739f
C192 VP.n39 B 0.021333f
C193 VP.n40 B 1.08479f
C194 VP.n41 B 1.38701f
C195 VP.n42 B 1.40019f
C196 VP.n43 B 1.08479f
C197 VP.n44 B 0.021333f
C198 VP.n45 B 0.038739f
C199 VP.n46 B 0.020785f
C200 VP.n47 B 0.020785f
C201 VP.n48 B 0.020785f
C202 VP.n49 B 0.017044f
C203 VP.n50 B 0.041807f
C204 VP.n51 B 0.038164f
C205 VP.n52 B 0.020785f
C206 VP.n53 B 0.020785f
C207 VP.n54 B 0.020186f
C208 VP.n55 B 0.038739f
C209 VP.n56 B 0.041311f
C210 VP.n57 B 0.020785f
C211 VP.n58 B 0.020785f
C212 VP.n59 B 0.020785f
C213 VP.n60 B 0.041311f
C214 VP.n61 B 0.038739f
C215 VP.n62 B 0.020186f
C216 VP.n63 B 0.020785f
C217 VP.n64 B 0.020785f
C218 VP.n65 B 0.038164f
C219 VP.n66 B 0.041807f
C220 VP.n67 B 0.017044f
C221 VP.n68 B 0.020785f
C222 VP.n69 B 0.020785f
C223 VP.n70 B 0.020785f
C224 VP.n71 B 0.038739f
C225 VP.n72 B 0.021333f
C226 VP.n73 B 1.08479f
C227 VP.n74 B 0.038214f
.ends

