* NGSPICE file created from diff_pair_sample_1250.ext - technology: sky130A

.subckt diff_pair_sample_1250 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=2.4024 pd=13.1 as=0 ps=0 w=6.16 l=0.51
X1 VDD2.t1 VN.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=2.4024 pd=13.1 as=2.4024 ps=13.1 w=6.16 l=0.51
X2 VDD2.t0 VN.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.4024 pd=13.1 as=2.4024 ps=13.1 w=6.16 l=0.51
X3 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=2.4024 pd=13.1 as=0 ps=0 w=6.16 l=0.51
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.4024 pd=13.1 as=0 ps=0 w=6.16 l=0.51
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.4024 pd=13.1 as=0 ps=0 w=6.16 l=0.51
X6 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.4024 pd=13.1 as=2.4024 ps=13.1 w=6.16 l=0.51
X7 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.4024 pd=13.1 as=2.4024 ps=13.1 w=6.16 l=0.51
R0 B.n413 B.n412 585
R1 B.n414 B.n413 585
R2 B.n178 B.n57 585
R3 B.n177 B.n176 585
R4 B.n175 B.n174 585
R5 B.n173 B.n172 585
R6 B.n171 B.n170 585
R7 B.n169 B.n168 585
R8 B.n167 B.n166 585
R9 B.n165 B.n164 585
R10 B.n163 B.n162 585
R11 B.n161 B.n160 585
R12 B.n159 B.n158 585
R13 B.n157 B.n156 585
R14 B.n155 B.n154 585
R15 B.n153 B.n152 585
R16 B.n151 B.n150 585
R17 B.n149 B.n148 585
R18 B.n147 B.n146 585
R19 B.n145 B.n144 585
R20 B.n143 B.n142 585
R21 B.n141 B.n140 585
R22 B.n139 B.n138 585
R23 B.n137 B.n136 585
R24 B.n135 B.n134 585
R25 B.n133 B.n132 585
R26 B.n131 B.n130 585
R27 B.n129 B.n128 585
R28 B.n127 B.n126 585
R29 B.n125 B.n124 585
R30 B.n123 B.n122 585
R31 B.n121 B.n120 585
R32 B.n119 B.n118 585
R33 B.n117 B.n116 585
R34 B.n115 B.n114 585
R35 B.n112 B.n111 585
R36 B.n110 B.n109 585
R37 B.n108 B.n107 585
R38 B.n106 B.n105 585
R39 B.n104 B.n103 585
R40 B.n102 B.n101 585
R41 B.n100 B.n99 585
R42 B.n98 B.n97 585
R43 B.n96 B.n95 585
R44 B.n94 B.n93 585
R45 B.n92 B.n91 585
R46 B.n90 B.n89 585
R47 B.n88 B.n87 585
R48 B.n86 B.n85 585
R49 B.n84 B.n83 585
R50 B.n82 B.n81 585
R51 B.n80 B.n79 585
R52 B.n78 B.n77 585
R53 B.n76 B.n75 585
R54 B.n74 B.n73 585
R55 B.n72 B.n71 585
R56 B.n70 B.n69 585
R57 B.n68 B.n67 585
R58 B.n66 B.n65 585
R59 B.n64 B.n63 585
R60 B.n411 B.n27 585
R61 B.n415 B.n27 585
R62 B.n410 B.n26 585
R63 B.n416 B.n26 585
R64 B.n409 B.n408 585
R65 B.n408 B.n22 585
R66 B.n407 B.n21 585
R67 B.n422 B.n21 585
R68 B.n406 B.n20 585
R69 B.n423 B.n20 585
R70 B.n405 B.n19 585
R71 B.n424 B.n19 585
R72 B.n404 B.n403 585
R73 B.n403 B.n15 585
R74 B.n402 B.n14 585
R75 B.n430 B.n14 585
R76 B.n401 B.n13 585
R77 B.n431 B.n13 585
R78 B.n400 B.n12 585
R79 B.n432 B.n12 585
R80 B.n399 B.n398 585
R81 B.n398 B.n11 585
R82 B.n397 B.n7 585
R83 B.n438 B.n7 585
R84 B.n396 B.n6 585
R85 B.n439 B.n6 585
R86 B.n395 B.n5 585
R87 B.n440 B.n5 585
R88 B.n394 B.n393 585
R89 B.n393 B.n4 585
R90 B.n392 B.n179 585
R91 B.n392 B.n391 585
R92 B.n381 B.n180 585
R93 B.n384 B.n180 585
R94 B.n383 B.n382 585
R95 B.n385 B.n383 585
R96 B.n380 B.n185 585
R97 B.n185 B.n184 585
R98 B.n379 B.n378 585
R99 B.n378 B.n377 585
R100 B.n187 B.n186 585
R101 B.n188 B.n187 585
R102 B.n370 B.n369 585
R103 B.n371 B.n370 585
R104 B.n368 B.n192 585
R105 B.n196 B.n192 585
R106 B.n367 B.n366 585
R107 B.n366 B.n365 585
R108 B.n194 B.n193 585
R109 B.n195 B.n194 585
R110 B.n358 B.n357 585
R111 B.n359 B.n358 585
R112 B.n356 B.n201 585
R113 B.n201 B.n200 585
R114 B.n350 B.n349 585
R115 B.n348 B.n232 585
R116 B.n347 B.n231 585
R117 B.n352 B.n231 585
R118 B.n346 B.n345 585
R119 B.n344 B.n343 585
R120 B.n342 B.n341 585
R121 B.n340 B.n339 585
R122 B.n338 B.n337 585
R123 B.n336 B.n335 585
R124 B.n334 B.n333 585
R125 B.n332 B.n331 585
R126 B.n330 B.n329 585
R127 B.n328 B.n327 585
R128 B.n326 B.n325 585
R129 B.n324 B.n323 585
R130 B.n322 B.n321 585
R131 B.n320 B.n319 585
R132 B.n318 B.n317 585
R133 B.n316 B.n315 585
R134 B.n314 B.n313 585
R135 B.n312 B.n311 585
R136 B.n310 B.n309 585
R137 B.n308 B.n307 585
R138 B.n306 B.n305 585
R139 B.n304 B.n303 585
R140 B.n302 B.n301 585
R141 B.n300 B.n299 585
R142 B.n298 B.n297 585
R143 B.n296 B.n295 585
R144 B.n294 B.n293 585
R145 B.n292 B.n291 585
R146 B.n290 B.n289 585
R147 B.n288 B.n287 585
R148 B.n286 B.n285 585
R149 B.n283 B.n282 585
R150 B.n281 B.n280 585
R151 B.n279 B.n278 585
R152 B.n277 B.n276 585
R153 B.n275 B.n274 585
R154 B.n273 B.n272 585
R155 B.n271 B.n270 585
R156 B.n269 B.n268 585
R157 B.n267 B.n266 585
R158 B.n265 B.n264 585
R159 B.n263 B.n262 585
R160 B.n261 B.n260 585
R161 B.n259 B.n258 585
R162 B.n257 B.n256 585
R163 B.n255 B.n254 585
R164 B.n253 B.n252 585
R165 B.n251 B.n250 585
R166 B.n249 B.n248 585
R167 B.n247 B.n246 585
R168 B.n245 B.n244 585
R169 B.n243 B.n242 585
R170 B.n241 B.n240 585
R171 B.n239 B.n238 585
R172 B.n203 B.n202 585
R173 B.n355 B.n354 585
R174 B.n199 B.n198 585
R175 B.n200 B.n199 585
R176 B.n361 B.n360 585
R177 B.n360 B.n359 585
R178 B.n362 B.n197 585
R179 B.n197 B.n195 585
R180 B.n364 B.n363 585
R181 B.n365 B.n364 585
R182 B.n191 B.n190 585
R183 B.n196 B.n191 585
R184 B.n373 B.n372 585
R185 B.n372 B.n371 585
R186 B.n374 B.n189 585
R187 B.n189 B.n188 585
R188 B.n376 B.n375 585
R189 B.n377 B.n376 585
R190 B.n183 B.n182 585
R191 B.n184 B.n183 585
R192 B.n387 B.n386 585
R193 B.n386 B.n385 585
R194 B.n388 B.n181 585
R195 B.n384 B.n181 585
R196 B.n390 B.n389 585
R197 B.n391 B.n390 585
R198 B.n2 B.n0 585
R199 B.n4 B.n2 585
R200 B.n3 B.n1 585
R201 B.n439 B.n3 585
R202 B.n437 B.n436 585
R203 B.n438 B.n437 585
R204 B.n435 B.n8 585
R205 B.n11 B.n8 585
R206 B.n434 B.n433 585
R207 B.n433 B.n432 585
R208 B.n10 B.n9 585
R209 B.n431 B.n10 585
R210 B.n429 B.n428 585
R211 B.n430 B.n429 585
R212 B.n427 B.n16 585
R213 B.n16 B.n15 585
R214 B.n426 B.n425 585
R215 B.n425 B.n424 585
R216 B.n18 B.n17 585
R217 B.n423 B.n18 585
R218 B.n421 B.n420 585
R219 B.n422 B.n421 585
R220 B.n419 B.n23 585
R221 B.n23 B.n22 585
R222 B.n418 B.n417 585
R223 B.n417 B.n416 585
R224 B.n25 B.n24 585
R225 B.n415 B.n25 585
R226 B.n442 B.n441 585
R227 B.n441 B.n440 585
R228 B.n236 B.t13 497.262
R229 B.n233 B.t6 497.262
R230 B.n61 B.t10 497.262
R231 B.n58 B.t2 497.262
R232 B.n350 B.n199 473.281
R233 B.n63 B.n25 473.281
R234 B.n354 B.n201 473.281
R235 B.n413 B.n27 473.281
R236 B.n414 B.n56 256.663
R237 B.n414 B.n55 256.663
R238 B.n414 B.n54 256.663
R239 B.n414 B.n53 256.663
R240 B.n414 B.n52 256.663
R241 B.n414 B.n51 256.663
R242 B.n414 B.n50 256.663
R243 B.n414 B.n49 256.663
R244 B.n414 B.n48 256.663
R245 B.n414 B.n47 256.663
R246 B.n414 B.n46 256.663
R247 B.n414 B.n45 256.663
R248 B.n414 B.n44 256.663
R249 B.n414 B.n43 256.663
R250 B.n414 B.n42 256.663
R251 B.n414 B.n41 256.663
R252 B.n414 B.n40 256.663
R253 B.n414 B.n39 256.663
R254 B.n414 B.n38 256.663
R255 B.n414 B.n37 256.663
R256 B.n414 B.n36 256.663
R257 B.n414 B.n35 256.663
R258 B.n414 B.n34 256.663
R259 B.n414 B.n33 256.663
R260 B.n414 B.n32 256.663
R261 B.n414 B.n31 256.663
R262 B.n414 B.n30 256.663
R263 B.n414 B.n29 256.663
R264 B.n414 B.n28 256.663
R265 B.n352 B.n351 256.663
R266 B.n352 B.n204 256.663
R267 B.n352 B.n205 256.663
R268 B.n352 B.n206 256.663
R269 B.n352 B.n207 256.663
R270 B.n352 B.n208 256.663
R271 B.n352 B.n209 256.663
R272 B.n352 B.n210 256.663
R273 B.n352 B.n211 256.663
R274 B.n352 B.n212 256.663
R275 B.n352 B.n213 256.663
R276 B.n352 B.n214 256.663
R277 B.n352 B.n215 256.663
R278 B.n352 B.n216 256.663
R279 B.n352 B.n217 256.663
R280 B.n352 B.n218 256.663
R281 B.n352 B.n219 256.663
R282 B.n352 B.n220 256.663
R283 B.n352 B.n221 256.663
R284 B.n352 B.n222 256.663
R285 B.n352 B.n223 256.663
R286 B.n352 B.n224 256.663
R287 B.n352 B.n225 256.663
R288 B.n352 B.n226 256.663
R289 B.n352 B.n227 256.663
R290 B.n352 B.n228 256.663
R291 B.n352 B.n229 256.663
R292 B.n352 B.n230 256.663
R293 B.n353 B.n352 256.663
R294 B.n360 B.n199 163.367
R295 B.n360 B.n197 163.367
R296 B.n364 B.n197 163.367
R297 B.n364 B.n191 163.367
R298 B.n372 B.n191 163.367
R299 B.n372 B.n189 163.367
R300 B.n376 B.n189 163.367
R301 B.n376 B.n183 163.367
R302 B.n386 B.n183 163.367
R303 B.n386 B.n181 163.367
R304 B.n390 B.n181 163.367
R305 B.n390 B.n2 163.367
R306 B.n441 B.n2 163.367
R307 B.n441 B.n3 163.367
R308 B.n437 B.n3 163.367
R309 B.n437 B.n8 163.367
R310 B.n433 B.n8 163.367
R311 B.n433 B.n10 163.367
R312 B.n429 B.n10 163.367
R313 B.n429 B.n16 163.367
R314 B.n425 B.n16 163.367
R315 B.n425 B.n18 163.367
R316 B.n421 B.n18 163.367
R317 B.n421 B.n23 163.367
R318 B.n417 B.n23 163.367
R319 B.n417 B.n25 163.367
R320 B.n232 B.n231 163.367
R321 B.n345 B.n231 163.367
R322 B.n343 B.n342 163.367
R323 B.n339 B.n338 163.367
R324 B.n335 B.n334 163.367
R325 B.n331 B.n330 163.367
R326 B.n327 B.n326 163.367
R327 B.n323 B.n322 163.367
R328 B.n319 B.n318 163.367
R329 B.n315 B.n314 163.367
R330 B.n311 B.n310 163.367
R331 B.n307 B.n306 163.367
R332 B.n303 B.n302 163.367
R333 B.n299 B.n298 163.367
R334 B.n295 B.n294 163.367
R335 B.n291 B.n290 163.367
R336 B.n287 B.n286 163.367
R337 B.n282 B.n281 163.367
R338 B.n278 B.n277 163.367
R339 B.n274 B.n273 163.367
R340 B.n270 B.n269 163.367
R341 B.n266 B.n265 163.367
R342 B.n262 B.n261 163.367
R343 B.n258 B.n257 163.367
R344 B.n254 B.n253 163.367
R345 B.n250 B.n249 163.367
R346 B.n246 B.n245 163.367
R347 B.n242 B.n241 163.367
R348 B.n238 B.n203 163.367
R349 B.n358 B.n201 163.367
R350 B.n358 B.n194 163.367
R351 B.n366 B.n194 163.367
R352 B.n366 B.n192 163.367
R353 B.n370 B.n192 163.367
R354 B.n370 B.n187 163.367
R355 B.n378 B.n187 163.367
R356 B.n378 B.n185 163.367
R357 B.n383 B.n185 163.367
R358 B.n383 B.n180 163.367
R359 B.n392 B.n180 163.367
R360 B.n393 B.n392 163.367
R361 B.n393 B.n5 163.367
R362 B.n6 B.n5 163.367
R363 B.n7 B.n6 163.367
R364 B.n398 B.n7 163.367
R365 B.n398 B.n12 163.367
R366 B.n13 B.n12 163.367
R367 B.n14 B.n13 163.367
R368 B.n403 B.n14 163.367
R369 B.n403 B.n19 163.367
R370 B.n20 B.n19 163.367
R371 B.n21 B.n20 163.367
R372 B.n408 B.n21 163.367
R373 B.n408 B.n26 163.367
R374 B.n27 B.n26 163.367
R375 B.n67 B.n66 163.367
R376 B.n71 B.n70 163.367
R377 B.n75 B.n74 163.367
R378 B.n79 B.n78 163.367
R379 B.n83 B.n82 163.367
R380 B.n87 B.n86 163.367
R381 B.n91 B.n90 163.367
R382 B.n95 B.n94 163.367
R383 B.n99 B.n98 163.367
R384 B.n103 B.n102 163.367
R385 B.n107 B.n106 163.367
R386 B.n111 B.n110 163.367
R387 B.n116 B.n115 163.367
R388 B.n120 B.n119 163.367
R389 B.n124 B.n123 163.367
R390 B.n128 B.n127 163.367
R391 B.n132 B.n131 163.367
R392 B.n136 B.n135 163.367
R393 B.n140 B.n139 163.367
R394 B.n144 B.n143 163.367
R395 B.n148 B.n147 163.367
R396 B.n152 B.n151 163.367
R397 B.n156 B.n155 163.367
R398 B.n160 B.n159 163.367
R399 B.n164 B.n163 163.367
R400 B.n168 B.n167 163.367
R401 B.n172 B.n171 163.367
R402 B.n176 B.n175 163.367
R403 B.n413 B.n57 163.367
R404 B.n352 B.n200 121.956
R405 B.n415 B.n414 121.956
R406 B.n236 B.t15 86.4241
R407 B.n58 B.t4 86.4241
R408 B.n233 B.t9 86.4173
R409 B.n61 B.t11 86.4173
R410 B.n351 B.n350 71.676
R411 B.n345 B.n204 71.676
R412 B.n342 B.n205 71.676
R413 B.n338 B.n206 71.676
R414 B.n334 B.n207 71.676
R415 B.n330 B.n208 71.676
R416 B.n326 B.n209 71.676
R417 B.n322 B.n210 71.676
R418 B.n318 B.n211 71.676
R419 B.n314 B.n212 71.676
R420 B.n310 B.n213 71.676
R421 B.n306 B.n214 71.676
R422 B.n302 B.n215 71.676
R423 B.n298 B.n216 71.676
R424 B.n294 B.n217 71.676
R425 B.n290 B.n218 71.676
R426 B.n286 B.n219 71.676
R427 B.n281 B.n220 71.676
R428 B.n277 B.n221 71.676
R429 B.n273 B.n222 71.676
R430 B.n269 B.n223 71.676
R431 B.n265 B.n224 71.676
R432 B.n261 B.n225 71.676
R433 B.n257 B.n226 71.676
R434 B.n253 B.n227 71.676
R435 B.n249 B.n228 71.676
R436 B.n245 B.n229 71.676
R437 B.n241 B.n230 71.676
R438 B.n353 B.n203 71.676
R439 B.n63 B.n28 71.676
R440 B.n67 B.n29 71.676
R441 B.n71 B.n30 71.676
R442 B.n75 B.n31 71.676
R443 B.n79 B.n32 71.676
R444 B.n83 B.n33 71.676
R445 B.n87 B.n34 71.676
R446 B.n91 B.n35 71.676
R447 B.n95 B.n36 71.676
R448 B.n99 B.n37 71.676
R449 B.n103 B.n38 71.676
R450 B.n107 B.n39 71.676
R451 B.n111 B.n40 71.676
R452 B.n116 B.n41 71.676
R453 B.n120 B.n42 71.676
R454 B.n124 B.n43 71.676
R455 B.n128 B.n44 71.676
R456 B.n132 B.n45 71.676
R457 B.n136 B.n46 71.676
R458 B.n140 B.n47 71.676
R459 B.n144 B.n48 71.676
R460 B.n148 B.n49 71.676
R461 B.n152 B.n50 71.676
R462 B.n156 B.n51 71.676
R463 B.n160 B.n52 71.676
R464 B.n164 B.n53 71.676
R465 B.n168 B.n54 71.676
R466 B.n172 B.n55 71.676
R467 B.n176 B.n56 71.676
R468 B.n57 B.n56 71.676
R469 B.n175 B.n55 71.676
R470 B.n171 B.n54 71.676
R471 B.n167 B.n53 71.676
R472 B.n163 B.n52 71.676
R473 B.n159 B.n51 71.676
R474 B.n155 B.n50 71.676
R475 B.n151 B.n49 71.676
R476 B.n147 B.n48 71.676
R477 B.n143 B.n47 71.676
R478 B.n139 B.n46 71.676
R479 B.n135 B.n45 71.676
R480 B.n131 B.n44 71.676
R481 B.n127 B.n43 71.676
R482 B.n123 B.n42 71.676
R483 B.n119 B.n41 71.676
R484 B.n115 B.n40 71.676
R485 B.n110 B.n39 71.676
R486 B.n106 B.n38 71.676
R487 B.n102 B.n37 71.676
R488 B.n98 B.n36 71.676
R489 B.n94 B.n35 71.676
R490 B.n90 B.n34 71.676
R491 B.n86 B.n33 71.676
R492 B.n82 B.n32 71.676
R493 B.n78 B.n31 71.676
R494 B.n74 B.n30 71.676
R495 B.n70 B.n29 71.676
R496 B.n66 B.n28 71.676
R497 B.n351 B.n232 71.676
R498 B.n343 B.n204 71.676
R499 B.n339 B.n205 71.676
R500 B.n335 B.n206 71.676
R501 B.n331 B.n207 71.676
R502 B.n327 B.n208 71.676
R503 B.n323 B.n209 71.676
R504 B.n319 B.n210 71.676
R505 B.n315 B.n211 71.676
R506 B.n311 B.n212 71.676
R507 B.n307 B.n213 71.676
R508 B.n303 B.n214 71.676
R509 B.n299 B.n215 71.676
R510 B.n295 B.n216 71.676
R511 B.n291 B.n217 71.676
R512 B.n287 B.n218 71.676
R513 B.n282 B.n219 71.676
R514 B.n278 B.n220 71.676
R515 B.n274 B.n221 71.676
R516 B.n270 B.n222 71.676
R517 B.n266 B.n223 71.676
R518 B.n262 B.n224 71.676
R519 B.n258 B.n225 71.676
R520 B.n254 B.n226 71.676
R521 B.n250 B.n227 71.676
R522 B.n246 B.n228 71.676
R523 B.n242 B.n229 71.676
R524 B.n238 B.n230 71.676
R525 B.n354 B.n353 71.676
R526 B.n237 B.t14 70.1332
R527 B.n59 B.t5 70.1332
R528 B.n234 B.t8 70.1264
R529 B.n62 B.t12 70.1264
R530 B.n359 B.n200 65.2995
R531 B.n359 B.n195 65.2995
R532 B.n365 B.n195 65.2995
R533 B.n365 B.n196 65.2995
R534 B.n371 B.n188 65.2995
R535 B.n377 B.n188 65.2995
R536 B.n377 B.n184 65.2995
R537 B.n385 B.n184 65.2995
R538 B.n385 B.n384 65.2995
R539 B.n391 B.n4 65.2995
R540 B.n440 B.n4 65.2995
R541 B.n440 B.n439 65.2995
R542 B.n439 B.n438 65.2995
R543 B.n432 B.n11 65.2995
R544 B.n432 B.n431 65.2995
R545 B.n431 B.n430 65.2995
R546 B.n430 B.n15 65.2995
R547 B.n424 B.n15 65.2995
R548 B.n423 B.n422 65.2995
R549 B.n422 B.n22 65.2995
R550 B.n416 B.n22 65.2995
R551 B.n416 B.n415 65.2995
R552 B.n284 B.n237 59.5399
R553 B.n235 B.n234 59.5399
R554 B.n113 B.n62 59.5399
R555 B.n60 B.n59 59.5399
R556 B.n391 B.t0 54.7364
R557 B.n438 B.t1 54.7364
R558 B.n371 B.t7 33.6103
R559 B.n424 B.t3 33.6103
R560 B.n196 B.t7 31.6897
R561 B.t3 B.n423 31.6897
R562 B.n412 B.n411 30.7517
R563 B.n64 B.n24 30.7517
R564 B.n356 B.n355 30.7517
R565 B.n349 B.n198 30.7517
R566 B B.n442 18.0485
R567 B.n237 B.n236 16.2914
R568 B.n234 B.n233 16.2914
R569 B.n62 B.n61 16.2914
R570 B.n59 B.n58 16.2914
R571 B.n65 B.n64 10.6151
R572 B.n68 B.n65 10.6151
R573 B.n69 B.n68 10.6151
R574 B.n72 B.n69 10.6151
R575 B.n73 B.n72 10.6151
R576 B.n76 B.n73 10.6151
R577 B.n77 B.n76 10.6151
R578 B.n80 B.n77 10.6151
R579 B.n81 B.n80 10.6151
R580 B.n84 B.n81 10.6151
R581 B.n85 B.n84 10.6151
R582 B.n88 B.n85 10.6151
R583 B.n89 B.n88 10.6151
R584 B.n92 B.n89 10.6151
R585 B.n93 B.n92 10.6151
R586 B.n96 B.n93 10.6151
R587 B.n97 B.n96 10.6151
R588 B.n100 B.n97 10.6151
R589 B.n101 B.n100 10.6151
R590 B.n104 B.n101 10.6151
R591 B.n105 B.n104 10.6151
R592 B.n108 B.n105 10.6151
R593 B.n109 B.n108 10.6151
R594 B.n112 B.n109 10.6151
R595 B.n117 B.n114 10.6151
R596 B.n118 B.n117 10.6151
R597 B.n121 B.n118 10.6151
R598 B.n122 B.n121 10.6151
R599 B.n125 B.n122 10.6151
R600 B.n126 B.n125 10.6151
R601 B.n129 B.n126 10.6151
R602 B.n130 B.n129 10.6151
R603 B.n134 B.n133 10.6151
R604 B.n137 B.n134 10.6151
R605 B.n138 B.n137 10.6151
R606 B.n141 B.n138 10.6151
R607 B.n142 B.n141 10.6151
R608 B.n145 B.n142 10.6151
R609 B.n146 B.n145 10.6151
R610 B.n149 B.n146 10.6151
R611 B.n150 B.n149 10.6151
R612 B.n153 B.n150 10.6151
R613 B.n154 B.n153 10.6151
R614 B.n157 B.n154 10.6151
R615 B.n158 B.n157 10.6151
R616 B.n161 B.n158 10.6151
R617 B.n162 B.n161 10.6151
R618 B.n165 B.n162 10.6151
R619 B.n166 B.n165 10.6151
R620 B.n169 B.n166 10.6151
R621 B.n170 B.n169 10.6151
R622 B.n173 B.n170 10.6151
R623 B.n174 B.n173 10.6151
R624 B.n177 B.n174 10.6151
R625 B.n178 B.n177 10.6151
R626 B.n412 B.n178 10.6151
R627 B.n357 B.n356 10.6151
R628 B.n357 B.n193 10.6151
R629 B.n367 B.n193 10.6151
R630 B.n368 B.n367 10.6151
R631 B.n369 B.n368 10.6151
R632 B.n369 B.n186 10.6151
R633 B.n379 B.n186 10.6151
R634 B.n380 B.n379 10.6151
R635 B.n382 B.n380 10.6151
R636 B.n382 B.n381 10.6151
R637 B.n381 B.n179 10.6151
R638 B.n394 B.n179 10.6151
R639 B.n395 B.n394 10.6151
R640 B.n396 B.n395 10.6151
R641 B.n397 B.n396 10.6151
R642 B.n399 B.n397 10.6151
R643 B.n400 B.n399 10.6151
R644 B.n401 B.n400 10.6151
R645 B.n402 B.n401 10.6151
R646 B.n404 B.n402 10.6151
R647 B.n405 B.n404 10.6151
R648 B.n406 B.n405 10.6151
R649 B.n407 B.n406 10.6151
R650 B.n409 B.n407 10.6151
R651 B.n410 B.n409 10.6151
R652 B.n411 B.n410 10.6151
R653 B.n349 B.n348 10.6151
R654 B.n348 B.n347 10.6151
R655 B.n347 B.n346 10.6151
R656 B.n346 B.n344 10.6151
R657 B.n344 B.n341 10.6151
R658 B.n341 B.n340 10.6151
R659 B.n340 B.n337 10.6151
R660 B.n337 B.n336 10.6151
R661 B.n336 B.n333 10.6151
R662 B.n333 B.n332 10.6151
R663 B.n332 B.n329 10.6151
R664 B.n329 B.n328 10.6151
R665 B.n328 B.n325 10.6151
R666 B.n325 B.n324 10.6151
R667 B.n324 B.n321 10.6151
R668 B.n321 B.n320 10.6151
R669 B.n320 B.n317 10.6151
R670 B.n317 B.n316 10.6151
R671 B.n316 B.n313 10.6151
R672 B.n313 B.n312 10.6151
R673 B.n312 B.n309 10.6151
R674 B.n309 B.n308 10.6151
R675 B.n308 B.n305 10.6151
R676 B.n305 B.n304 10.6151
R677 B.n301 B.n300 10.6151
R678 B.n300 B.n297 10.6151
R679 B.n297 B.n296 10.6151
R680 B.n296 B.n293 10.6151
R681 B.n293 B.n292 10.6151
R682 B.n292 B.n289 10.6151
R683 B.n289 B.n288 10.6151
R684 B.n288 B.n285 10.6151
R685 B.n283 B.n280 10.6151
R686 B.n280 B.n279 10.6151
R687 B.n279 B.n276 10.6151
R688 B.n276 B.n275 10.6151
R689 B.n275 B.n272 10.6151
R690 B.n272 B.n271 10.6151
R691 B.n271 B.n268 10.6151
R692 B.n268 B.n267 10.6151
R693 B.n267 B.n264 10.6151
R694 B.n264 B.n263 10.6151
R695 B.n263 B.n260 10.6151
R696 B.n260 B.n259 10.6151
R697 B.n259 B.n256 10.6151
R698 B.n256 B.n255 10.6151
R699 B.n255 B.n252 10.6151
R700 B.n252 B.n251 10.6151
R701 B.n251 B.n248 10.6151
R702 B.n248 B.n247 10.6151
R703 B.n247 B.n244 10.6151
R704 B.n244 B.n243 10.6151
R705 B.n243 B.n240 10.6151
R706 B.n240 B.n239 10.6151
R707 B.n239 B.n202 10.6151
R708 B.n355 B.n202 10.6151
R709 B.n361 B.n198 10.6151
R710 B.n362 B.n361 10.6151
R711 B.n363 B.n362 10.6151
R712 B.n363 B.n190 10.6151
R713 B.n373 B.n190 10.6151
R714 B.n374 B.n373 10.6151
R715 B.n375 B.n374 10.6151
R716 B.n375 B.n182 10.6151
R717 B.n387 B.n182 10.6151
R718 B.n388 B.n387 10.6151
R719 B.n389 B.n388 10.6151
R720 B.n389 B.n0 10.6151
R721 B.n436 B.n1 10.6151
R722 B.n436 B.n435 10.6151
R723 B.n435 B.n434 10.6151
R724 B.n434 B.n9 10.6151
R725 B.n428 B.n9 10.6151
R726 B.n428 B.n427 10.6151
R727 B.n427 B.n426 10.6151
R728 B.n426 B.n17 10.6151
R729 B.n420 B.n17 10.6151
R730 B.n420 B.n419 10.6151
R731 B.n419 B.n418 10.6151
R732 B.n418 B.n24 10.6151
R733 B.n384 B.t0 10.5636
R734 B.n11 B.t1 10.5636
R735 B.n114 B.n113 7.18099
R736 B.n130 B.n60 7.18099
R737 B.n301 B.n235 7.18099
R738 B.n285 B.n284 7.18099
R739 B.n113 B.n112 3.43465
R740 B.n133 B.n60 3.43465
R741 B.n304 B.n235 3.43465
R742 B.n284 B.n283 3.43465
R743 B.n442 B.n0 2.81026
R744 B.n442 B.n1 2.81026
R745 VN VN.t0 564.501
R746 VN VN.t1 529.467
R747 VTAIL.n1 VTAIL.t3 55.5006
R748 VTAIL.n2 VTAIL.t1 55.4996
R749 VTAIL.n3 VTAIL.t2 55.4996
R750 VTAIL.n0 VTAIL.t0 55.4996
R751 VTAIL.n1 VTAIL.n0 19.1427
R752 VTAIL.n3 VTAIL.n2 18.4186
R753 VTAIL.n2 VTAIL.n1 0.832397
R754 VTAIL VTAIL.n0 0.709552
R755 VTAIL VTAIL.n3 0.123345
R756 VDD2.n0 VDD2.t0 102.614
R757 VDD2.n0 VDD2.t1 72.1784
R758 VDD2 VDD2.n0 0.239724
R759 VP.n0 VP.t1 564.12
R760 VP.n0 VP.t0 529.417
R761 VP VP.n0 0.0516364
R762 VDD1 VDD1.t1 103.32
R763 VDD1 VDD1.t0 72.4176
C0 VDD2 VP 0.246492f
C1 VDD2 VDD1 0.44274f
C2 VP VN 3.39233f
C3 VDD1 VN 0.148835f
C4 VTAIL VP 0.798692f
C5 VDD1 VTAIL 3.68715f
C6 VDD2 VN 1.02075f
C7 VDD1 VP 1.11592f
C8 VDD2 VTAIL 3.72255f
C9 VTAIL VN 0.784295f
C10 VDD2 B 2.620238f
C11 VDD1 B 4.4254f
C12 VTAIL B 3.696132f
C13 VN B 5.95784f
C14 VP B 3.356203f
C15 VDD1.t0 B 0.870596f
C16 VDD1.t1 B 1.11607f
C17 VP.t1 B 0.486958f
C18 VP.t0 B 0.408802f
C19 VP.n0 B 2.4951f
C20 VDD2.t0 B 1.11895f
C21 VDD2.t1 B 0.8847f
C22 VDD2.n0 B 1.66305f
C23 VTAIL.t0 B 0.933263f
C24 VTAIL.n0 B 0.931332f
C25 VTAIL.t3 B 0.933263f
C26 VTAIL.n1 B 0.938826f
C27 VTAIL.t1 B 0.933259f
C28 VTAIL.n2 B 0.894652f
C29 VTAIL.t2 B 0.933263f
C30 VTAIL.n3 B 0.85139f
C31 VN.t1 B 0.40224f
C32 VN.t0 B 0.481525f
.ends

