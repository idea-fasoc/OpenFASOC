* NGSPICE file created from diff_pair_sample_1394.ext - technology: sky130A

.subckt diff_pair_sample_1394 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9617 pd=10.84 as=0.82995 ps=5.36 w=5.03 l=1.93
X1 VTAIL.t11 VP.t1 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=0.82995 pd=5.36 as=0.82995 ps=5.36 w=5.03 l=1.93
X2 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=1.9617 pd=10.84 as=0 ps=0 w=5.03 l=1.93
X3 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=1.9617 pd=10.84 as=0 ps=0 w=5.03 l=1.93
X4 VDD1.t3 VP.t2 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=0.82995 pd=5.36 as=1.9617 ps=10.84 w=5.03 l=1.93
X5 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.9617 pd=10.84 as=0 ps=0 w=5.03 l=1.93
X6 VTAIL.t5 VN.t0 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.82995 pd=5.36 as=0.82995 ps=5.36 w=5.03 l=1.93
X7 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.9617 pd=10.84 as=0 ps=0 w=5.03 l=1.93
X8 VDD2.t4 VN.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.82995 pd=5.36 as=1.9617 ps=10.84 w=5.03 l=1.93
X9 VDD2.t3 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.82995 pd=5.36 as=1.9617 ps=10.84 w=5.03 l=1.93
X10 VTAIL.t2 VN.t3 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.82995 pd=5.36 as=0.82995 ps=5.36 w=5.03 l=1.93
X11 VDD2.t1 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9617 pd=10.84 as=0.82995 ps=5.36 w=5.03 l=1.93
X12 VDD1.t2 VP.t3 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=0.82995 pd=5.36 as=1.9617 ps=10.84 w=5.03 l=1.93
X13 VTAIL.t7 VP.t4 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.82995 pd=5.36 as=0.82995 ps=5.36 w=5.03 l=1.93
X14 VDD2.t0 VN.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9617 pd=10.84 as=0.82995 ps=5.36 w=5.03 l=1.93
X15 VDD1.t0 VP.t5 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9617 pd=10.84 as=0.82995 ps=5.36 w=5.03 l=1.93
R0 VP.n20 VP.n5 185.279
R1 VP.n38 VP.n37 185.279
R2 VP.n19 VP.n18 185.279
R3 VP.n11 VP.n8 161.3
R4 VP.n13 VP.n12 161.3
R5 VP.n14 VP.n7 161.3
R6 VP.n16 VP.n15 161.3
R7 VP.n17 VP.n6 161.3
R8 VP.n36 VP.n0 161.3
R9 VP.n35 VP.n34 161.3
R10 VP.n33 VP.n1 161.3
R11 VP.n32 VP.n31 161.3
R12 VP.n30 VP.n2 161.3
R13 VP.n28 VP.n27 161.3
R14 VP.n26 VP.n3 161.3
R15 VP.n25 VP.n24 161.3
R16 VP.n23 VP.n4 161.3
R17 VP.n22 VP.n21 161.3
R18 VP.n9 VP.t5 94.5642
R19 VP.n5 VP.t0 62.8103
R20 VP.n29 VP.t1 62.8103
R21 VP.n37 VP.t2 62.8103
R22 VP.n18 VP.t3 62.8103
R23 VP.n10 VP.t4 62.8103
R24 VP.n10 VP.n9 57.9196
R25 VP.n24 VP.n3 52.1486
R26 VP.n31 VP.n1 52.1486
R27 VP.n12 VP.n7 52.1486
R28 VP.n20 VP.n19 40.652
R29 VP.n24 VP.n23 28.8382
R30 VP.n35 VP.n1 28.8382
R31 VP.n16 VP.n7 28.8382
R32 VP.n23 VP.n22 24.4675
R33 VP.n28 VP.n3 24.4675
R34 VP.n31 VP.n30 24.4675
R35 VP.n36 VP.n35 24.4675
R36 VP.n17 VP.n16 24.4675
R37 VP.n12 VP.n11 24.4675
R38 VP.n9 VP.n8 12.5909
R39 VP.n29 VP.n28 12.234
R40 VP.n30 VP.n29 12.234
R41 VP.n11 VP.n10 12.234
R42 VP.n22 VP.n5 0.48984
R43 VP.n37 VP.n36 0.48984
R44 VP.n18 VP.n17 0.48984
R45 VP.n13 VP.n8 0.189894
R46 VP.n14 VP.n13 0.189894
R47 VP.n15 VP.n14 0.189894
R48 VP.n15 VP.n6 0.189894
R49 VP.n19 VP.n6 0.189894
R50 VP.n21 VP.n20 0.189894
R51 VP.n21 VP.n4 0.189894
R52 VP.n25 VP.n4 0.189894
R53 VP.n26 VP.n25 0.189894
R54 VP.n27 VP.n26 0.189894
R55 VP.n27 VP.n2 0.189894
R56 VP.n32 VP.n2 0.189894
R57 VP.n33 VP.n32 0.189894
R58 VP.n34 VP.n33 0.189894
R59 VP.n34 VP.n0 0.189894
R60 VP.n38 VP.n0 0.189894
R61 VP VP.n38 0.0516364
R62 VTAIL.n7 VTAIL.t3 58.9579
R63 VTAIL.n11 VTAIL.t4 58.9579
R64 VTAIL.n2 VTAIL.t9 58.9579
R65 VTAIL.n10 VTAIL.t10 58.9579
R66 VTAIL.n9 VTAIL.n8 55.0216
R67 VTAIL.n6 VTAIL.n5 55.0216
R68 VTAIL.n1 VTAIL.n0 55.0214
R69 VTAIL.n4 VTAIL.n3 55.0214
R70 VTAIL.n6 VTAIL.n4 20.5996
R71 VTAIL.n11 VTAIL.n10 18.6514
R72 VTAIL.n0 VTAIL.t1 3.93688
R73 VTAIL.n0 VTAIL.t2 3.93688
R74 VTAIL.n3 VTAIL.t8 3.93688
R75 VTAIL.n3 VTAIL.t11 3.93688
R76 VTAIL.n8 VTAIL.t6 3.93688
R77 VTAIL.n8 VTAIL.t7 3.93688
R78 VTAIL.n5 VTAIL.t0 3.93688
R79 VTAIL.n5 VTAIL.t5 3.93688
R80 VTAIL.n7 VTAIL.n6 1.94878
R81 VTAIL.n10 VTAIL.n9 1.94878
R82 VTAIL.n4 VTAIL.n2 1.94878
R83 VTAIL.n9 VTAIL.n7 1.44447
R84 VTAIL.n2 VTAIL.n1 1.44447
R85 VTAIL VTAIL.n11 1.40352
R86 VTAIL VTAIL.n1 0.545759
R87 VDD1 VDD1.t0 77.1561
R88 VDD1.n1 VDD1.t5 77.0425
R89 VDD1.n1 VDD1.n0 72.1319
R90 VDD1.n3 VDD1.n2 71.7003
R91 VDD1.n3 VDD1.n1 35.9405
R92 VDD1.n2 VDD1.t1 3.93688
R93 VDD1.n2 VDD1.t2 3.93688
R94 VDD1.n0 VDD1.t4 3.93688
R95 VDD1.n0 VDD1.t3 3.93688
R96 VDD1 VDD1.n3 0.429379
R97 B.n446 B.n445 585
R98 B.n448 B.n96 585
R99 B.n451 B.n450 585
R100 B.n452 B.n95 585
R101 B.n454 B.n453 585
R102 B.n456 B.n94 585
R103 B.n459 B.n458 585
R104 B.n460 B.n93 585
R105 B.n462 B.n461 585
R106 B.n464 B.n92 585
R107 B.n467 B.n466 585
R108 B.n468 B.n91 585
R109 B.n470 B.n469 585
R110 B.n472 B.n90 585
R111 B.n475 B.n474 585
R112 B.n476 B.n89 585
R113 B.n478 B.n477 585
R114 B.n480 B.n88 585
R115 B.n483 B.n482 585
R116 B.n484 B.n84 585
R117 B.n486 B.n485 585
R118 B.n488 B.n83 585
R119 B.n491 B.n490 585
R120 B.n492 B.n82 585
R121 B.n494 B.n493 585
R122 B.n496 B.n81 585
R123 B.n499 B.n498 585
R124 B.n500 B.n80 585
R125 B.n502 B.n501 585
R126 B.n504 B.n79 585
R127 B.n507 B.n506 585
R128 B.n509 B.n76 585
R129 B.n511 B.n510 585
R130 B.n513 B.n75 585
R131 B.n516 B.n515 585
R132 B.n517 B.n74 585
R133 B.n519 B.n518 585
R134 B.n521 B.n73 585
R135 B.n524 B.n523 585
R136 B.n525 B.n72 585
R137 B.n527 B.n526 585
R138 B.n529 B.n71 585
R139 B.n532 B.n531 585
R140 B.n533 B.n70 585
R141 B.n535 B.n534 585
R142 B.n537 B.n69 585
R143 B.n540 B.n539 585
R144 B.n541 B.n68 585
R145 B.n543 B.n542 585
R146 B.n545 B.n67 585
R147 B.n548 B.n547 585
R148 B.n549 B.n66 585
R149 B.n444 B.n64 585
R150 B.n552 B.n64 585
R151 B.n443 B.n63 585
R152 B.n553 B.n63 585
R153 B.n442 B.n62 585
R154 B.n554 B.n62 585
R155 B.n441 B.n440 585
R156 B.n440 B.n58 585
R157 B.n439 B.n57 585
R158 B.n560 B.n57 585
R159 B.n438 B.n56 585
R160 B.n561 B.n56 585
R161 B.n437 B.n55 585
R162 B.n562 B.n55 585
R163 B.n436 B.n435 585
R164 B.n435 B.n51 585
R165 B.n434 B.n50 585
R166 B.n568 B.n50 585
R167 B.n433 B.n49 585
R168 B.n569 B.n49 585
R169 B.n432 B.n48 585
R170 B.n570 B.n48 585
R171 B.n431 B.n430 585
R172 B.n430 B.n44 585
R173 B.n429 B.n43 585
R174 B.n576 B.n43 585
R175 B.n428 B.n42 585
R176 B.n577 B.n42 585
R177 B.n427 B.n41 585
R178 B.n578 B.n41 585
R179 B.n426 B.n425 585
R180 B.n425 B.n37 585
R181 B.n424 B.n36 585
R182 B.n584 B.n36 585
R183 B.n423 B.n35 585
R184 B.n585 B.n35 585
R185 B.n422 B.n34 585
R186 B.n586 B.n34 585
R187 B.n421 B.n420 585
R188 B.n420 B.n30 585
R189 B.n419 B.n29 585
R190 B.n592 B.n29 585
R191 B.n418 B.n28 585
R192 B.n593 B.n28 585
R193 B.n417 B.n27 585
R194 B.n594 B.n27 585
R195 B.n416 B.n415 585
R196 B.n415 B.n23 585
R197 B.n414 B.n22 585
R198 B.n600 B.n22 585
R199 B.n413 B.n21 585
R200 B.n601 B.n21 585
R201 B.n412 B.n20 585
R202 B.n602 B.n20 585
R203 B.n411 B.n410 585
R204 B.n410 B.n16 585
R205 B.n409 B.n15 585
R206 B.n608 B.n15 585
R207 B.n408 B.n14 585
R208 B.n609 B.n14 585
R209 B.n407 B.n13 585
R210 B.n610 B.n13 585
R211 B.n406 B.n405 585
R212 B.n405 B.n12 585
R213 B.n404 B.n403 585
R214 B.n404 B.n8 585
R215 B.n402 B.n7 585
R216 B.n617 B.n7 585
R217 B.n401 B.n6 585
R218 B.n618 B.n6 585
R219 B.n400 B.n5 585
R220 B.n619 B.n5 585
R221 B.n399 B.n398 585
R222 B.n398 B.n4 585
R223 B.n397 B.n97 585
R224 B.n397 B.n396 585
R225 B.n387 B.n98 585
R226 B.n99 B.n98 585
R227 B.n389 B.n388 585
R228 B.n390 B.n389 585
R229 B.n386 B.n103 585
R230 B.n107 B.n103 585
R231 B.n385 B.n384 585
R232 B.n384 B.n383 585
R233 B.n105 B.n104 585
R234 B.n106 B.n105 585
R235 B.n376 B.n375 585
R236 B.n377 B.n376 585
R237 B.n374 B.n112 585
R238 B.n112 B.n111 585
R239 B.n373 B.n372 585
R240 B.n372 B.n371 585
R241 B.n114 B.n113 585
R242 B.n115 B.n114 585
R243 B.n364 B.n363 585
R244 B.n365 B.n364 585
R245 B.n362 B.n120 585
R246 B.n120 B.n119 585
R247 B.n361 B.n360 585
R248 B.n360 B.n359 585
R249 B.n122 B.n121 585
R250 B.n123 B.n122 585
R251 B.n352 B.n351 585
R252 B.n353 B.n352 585
R253 B.n350 B.n128 585
R254 B.n128 B.n127 585
R255 B.n349 B.n348 585
R256 B.n348 B.n347 585
R257 B.n130 B.n129 585
R258 B.n131 B.n130 585
R259 B.n340 B.n339 585
R260 B.n341 B.n340 585
R261 B.n338 B.n136 585
R262 B.n136 B.n135 585
R263 B.n337 B.n336 585
R264 B.n336 B.n335 585
R265 B.n138 B.n137 585
R266 B.n139 B.n138 585
R267 B.n328 B.n327 585
R268 B.n329 B.n328 585
R269 B.n326 B.n144 585
R270 B.n144 B.n143 585
R271 B.n325 B.n324 585
R272 B.n324 B.n323 585
R273 B.n146 B.n145 585
R274 B.n147 B.n146 585
R275 B.n316 B.n315 585
R276 B.n317 B.n316 585
R277 B.n314 B.n152 585
R278 B.n152 B.n151 585
R279 B.n313 B.n312 585
R280 B.n312 B.n311 585
R281 B.n154 B.n153 585
R282 B.n155 B.n154 585
R283 B.n304 B.n303 585
R284 B.n305 B.n304 585
R285 B.n302 B.n160 585
R286 B.n160 B.n159 585
R287 B.n301 B.n300 585
R288 B.n300 B.n299 585
R289 B.n296 B.n164 585
R290 B.n295 B.n294 585
R291 B.n292 B.n165 585
R292 B.n292 B.n163 585
R293 B.n291 B.n290 585
R294 B.n289 B.n288 585
R295 B.n287 B.n167 585
R296 B.n285 B.n284 585
R297 B.n283 B.n168 585
R298 B.n282 B.n281 585
R299 B.n279 B.n169 585
R300 B.n277 B.n276 585
R301 B.n275 B.n170 585
R302 B.n274 B.n273 585
R303 B.n271 B.n171 585
R304 B.n269 B.n268 585
R305 B.n267 B.n172 585
R306 B.n266 B.n265 585
R307 B.n263 B.n173 585
R308 B.n261 B.n260 585
R309 B.n259 B.n174 585
R310 B.n258 B.n257 585
R311 B.n255 B.n254 585
R312 B.n253 B.n252 585
R313 B.n251 B.n179 585
R314 B.n249 B.n248 585
R315 B.n247 B.n180 585
R316 B.n246 B.n245 585
R317 B.n243 B.n181 585
R318 B.n241 B.n240 585
R319 B.n239 B.n182 585
R320 B.n238 B.n237 585
R321 B.n235 B.n234 585
R322 B.n233 B.n232 585
R323 B.n231 B.n187 585
R324 B.n229 B.n228 585
R325 B.n227 B.n188 585
R326 B.n226 B.n225 585
R327 B.n223 B.n189 585
R328 B.n221 B.n220 585
R329 B.n219 B.n190 585
R330 B.n218 B.n217 585
R331 B.n215 B.n191 585
R332 B.n213 B.n212 585
R333 B.n211 B.n192 585
R334 B.n210 B.n209 585
R335 B.n207 B.n193 585
R336 B.n205 B.n204 585
R337 B.n203 B.n194 585
R338 B.n202 B.n201 585
R339 B.n199 B.n195 585
R340 B.n197 B.n196 585
R341 B.n162 B.n161 585
R342 B.n163 B.n162 585
R343 B.n298 B.n297 585
R344 B.n299 B.n298 585
R345 B.n158 B.n157 585
R346 B.n159 B.n158 585
R347 B.n307 B.n306 585
R348 B.n306 B.n305 585
R349 B.n308 B.n156 585
R350 B.n156 B.n155 585
R351 B.n310 B.n309 585
R352 B.n311 B.n310 585
R353 B.n150 B.n149 585
R354 B.n151 B.n150 585
R355 B.n319 B.n318 585
R356 B.n318 B.n317 585
R357 B.n320 B.n148 585
R358 B.n148 B.n147 585
R359 B.n322 B.n321 585
R360 B.n323 B.n322 585
R361 B.n142 B.n141 585
R362 B.n143 B.n142 585
R363 B.n331 B.n330 585
R364 B.n330 B.n329 585
R365 B.n332 B.n140 585
R366 B.n140 B.n139 585
R367 B.n334 B.n333 585
R368 B.n335 B.n334 585
R369 B.n134 B.n133 585
R370 B.n135 B.n134 585
R371 B.n343 B.n342 585
R372 B.n342 B.n341 585
R373 B.n344 B.n132 585
R374 B.n132 B.n131 585
R375 B.n346 B.n345 585
R376 B.n347 B.n346 585
R377 B.n126 B.n125 585
R378 B.n127 B.n126 585
R379 B.n355 B.n354 585
R380 B.n354 B.n353 585
R381 B.n356 B.n124 585
R382 B.n124 B.n123 585
R383 B.n358 B.n357 585
R384 B.n359 B.n358 585
R385 B.n118 B.n117 585
R386 B.n119 B.n118 585
R387 B.n367 B.n366 585
R388 B.n366 B.n365 585
R389 B.n368 B.n116 585
R390 B.n116 B.n115 585
R391 B.n370 B.n369 585
R392 B.n371 B.n370 585
R393 B.n110 B.n109 585
R394 B.n111 B.n110 585
R395 B.n379 B.n378 585
R396 B.n378 B.n377 585
R397 B.n380 B.n108 585
R398 B.n108 B.n106 585
R399 B.n382 B.n381 585
R400 B.n383 B.n382 585
R401 B.n102 B.n101 585
R402 B.n107 B.n102 585
R403 B.n392 B.n391 585
R404 B.n391 B.n390 585
R405 B.n393 B.n100 585
R406 B.n100 B.n99 585
R407 B.n395 B.n394 585
R408 B.n396 B.n395 585
R409 B.n3 B.n0 585
R410 B.n4 B.n3 585
R411 B.n616 B.n1 585
R412 B.n617 B.n616 585
R413 B.n615 B.n614 585
R414 B.n615 B.n8 585
R415 B.n613 B.n9 585
R416 B.n12 B.n9 585
R417 B.n612 B.n611 585
R418 B.n611 B.n610 585
R419 B.n11 B.n10 585
R420 B.n609 B.n11 585
R421 B.n607 B.n606 585
R422 B.n608 B.n607 585
R423 B.n605 B.n17 585
R424 B.n17 B.n16 585
R425 B.n604 B.n603 585
R426 B.n603 B.n602 585
R427 B.n19 B.n18 585
R428 B.n601 B.n19 585
R429 B.n599 B.n598 585
R430 B.n600 B.n599 585
R431 B.n597 B.n24 585
R432 B.n24 B.n23 585
R433 B.n596 B.n595 585
R434 B.n595 B.n594 585
R435 B.n26 B.n25 585
R436 B.n593 B.n26 585
R437 B.n591 B.n590 585
R438 B.n592 B.n591 585
R439 B.n589 B.n31 585
R440 B.n31 B.n30 585
R441 B.n588 B.n587 585
R442 B.n587 B.n586 585
R443 B.n33 B.n32 585
R444 B.n585 B.n33 585
R445 B.n583 B.n582 585
R446 B.n584 B.n583 585
R447 B.n581 B.n38 585
R448 B.n38 B.n37 585
R449 B.n580 B.n579 585
R450 B.n579 B.n578 585
R451 B.n40 B.n39 585
R452 B.n577 B.n40 585
R453 B.n575 B.n574 585
R454 B.n576 B.n575 585
R455 B.n573 B.n45 585
R456 B.n45 B.n44 585
R457 B.n572 B.n571 585
R458 B.n571 B.n570 585
R459 B.n47 B.n46 585
R460 B.n569 B.n47 585
R461 B.n567 B.n566 585
R462 B.n568 B.n567 585
R463 B.n565 B.n52 585
R464 B.n52 B.n51 585
R465 B.n564 B.n563 585
R466 B.n563 B.n562 585
R467 B.n54 B.n53 585
R468 B.n561 B.n54 585
R469 B.n559 B.n558 585
R470 B.n560 B.n559 585
R471 B.n557 B.n59 585
R472 B.n59 B.n58 585
R473 B.n556 B.n555 585
R474 B.n555 B.n554 585
R475 B.n61 B.n60 585
R476 B.n553 B.n61 585
R477 B.n551 B.n550 585
R478 B.n552 B.n551 585
R479 B.n620 B.n619 585
R480 B.n618 B.n2 585
R481 B.n551 B.n66 516.524
R482 B.n446 B.n64 516.524
R483 B.n300 B.n162 516.524
R484 B.n298 B.n164 516.524
R485 B.n77 B.t14 269.558
R486 B.n85 B.t6 269.558
R487 B.n183 B.t17 269.558
R488 B.n175 B.t10 269.558
R489 B.n447 B.n65 256.663
R490 B.n449 B.n65 256.663
R491 B.n455 B.n65 256.663
R492 B.n457 B.n65 256.663
R493 B.n463 B.n65 256.663
R494 B.n465 B.n65 256.663
R495 B.n471 B.n65 256.663
R496 B.n473 B.n65 256.663
R497 B.n479 B.n65 256.663
R498 B.n481 B.n65 256.663
R499 B.n487 B.n65 256.663
R500 B.n489 B.n65 256.663
R501 B.n495 B.n65 256.663
R502 B.n497 B.n65 256.663
R503 B.n503 B.n65 256.663
R504 B.n505 B.n65 256.663
R505 B.n512 B.n65 256.663
R506 B.n514 B.n65 256.663
R507 B.n520 B.n65 256.663
R508 B.n522 B.n65 256.663
R509 B.n528 B.n65 256.663
R510 B.n530 B.n65 256.663
R511 B.n536 B.n65 256.663
R512 B.n538 B.n65 256.663
R513 B.n544 B.n65 256.663
R514 B.n546 B.n65 256.663
R515 B.n293 B.n163 256.663
R516 B.n166 B.n163 256.663
R517 B.n286 B.n163 256.663
R518 B.n280 B.n163 256.663
R519 B.n278 B.n163 256.663
R520 B.n272 B.n163 256.663
R521 B.n270 B.n163 256.663
R522 B.n264 B.n163 256.663
R523 B.n262 B.n163 256.663
R524 B.n256 B.n163 256.663
R525 B.n178 B.n163 256.663
R526 B.n250 B.n163 256.663
R527 B.n244 B.n163 256.663
R528 B.n242 B.n163 256.663
R529 B.n236 B.n163 256.663
R530 B.n186 B.n163 256.663
R531 B.n230 B.n163 256.663
R532 B.n224 B.n163 256.663
R533 B.n222 B.n163 256.663
R534 B.n216 B.n163 256.663
R535 B.n214 B.n163 256.663
R536 B.n208 B.n163 256.663
R537 B.n206 B.n163 256.663
R538 B.n200 B.n163 256.663
R539 B.n198 B.n163 256.663
R540 B.n622 B.n621 256.663
R541 B.n547 B.n545 163.367
R542 B.n543 B.n68 163.367
R543 B.n539 B.n537 163.367
R544 B.n535 B.n70 163.367
R545 B.n531 B.n529 163.367
R546 B.n527 B.n72 163.367
R547 B.n523 B.n521 163.367
R548 B.n519 B.n74 163.367
R549 B.n515 B.n513 163.367
R550 B.n511 B.n76 163.367
R551 B.n506 B.n504 163.367
R552 B.n502 B.n80 163.367
R553 B.n498 B.n496 163.367
R554 B.n494 B.n82 163.367
R555 B.n490 B.n488 163.367
R556 B.n486 B.n84 163.367
R557 B.n482 B.n480 163.367
R558 B.n478 B.n89 163.367
R559 B.n474 B.n472 163.367
R560 B.n470 B.n91 163.367
R561 B.n466 B.n464 163.367
R562 B.n462 B.n93 163.367
R563 B.n458 B.n456 163.367
R564 B.n454 B.n95 163.367
R565 B.n450 B.n448 163.367
R566 B.n300 B.n160 163.367
R567 B.n304 B.n160 163.367
R568 B.n304 B.n154 163.367
R569 B.n312 B.n154 163.367
R570 B.n312 B.n152 163.367
R571 B.n316 B.n152 163.367
R572 B.n316 B.n146 163.367
R573 B.n324 B.n146 163.367
R574 B.n324 B.n144 163.367
R575 B.n328 B.n144 163.367
R576 B.n328 B.n138 163.367
R577 B.n336 B.n138 163.367
R578 B.n336 B.n136 163.367
R579 B.n340 B.n136 163.367
R580 B.n340 B.n130 163.367
R581 B.n348 B.n130 163.367
R582 B.n348 B.n128 163.367
R583 B.n352 B.n128 163.367
R584 B.n352 B.n122 163.367
R585 B.n360 B.n122 163.367
R586 B.n360 B.n120 163.367
R587 B.n364 B.n120 163.367
R588 B.n364 B.n114 163.367
R589 B.n372 B.n114 163.367
R590 B.n372 B.n112 163.367
R591 B.n376 B.n112 163.367
R592 B.n376 B.n105 163.367
R593 B.n384 B.n105 163.367
R594 B.n384 B.n103 163.367
R595 B.n389 B.n103 163.367
R596 B.n389 B.n98 163.367
R597 B.n397 B.n98 163.367
R598 B.n398 B.n397 163.367
R599 B.n398 B.n5 163.367
R600 B.n6 B.n5 163.367
R601 B.n7 B.n6 163.367
R602 B.n404 B.n7 163.367
R603 B.n405 B.n404 163.367
R604 B.n405 B.n13 163.367
R605 B.n14 B.n13 163.367
R606 B.n15 B.n14 163.367
R607 B.n410 B.n15 163.367
R608 B.n410 B.n20 163.367
R609 B.n21 B.n20 163.367
R610 B.n22 B.n21 163.367
R611 B.n415 B.n22 163.367
R612 B.n415 B.n27 163.367
R613 B.n28 B.n27 163.367
R614 B.n29 B.n28 163.367
R615 B.n420 B.n29 163.367
R616 B.n420 B.n34 163.367
R617 B.n35 B.n34 163.367
R618 B.n36 B.n35 163.367
R619 B.n425 B.n36 163.367
R620 B.n425 B.n41 163.367
R621 B.n42 B.n41 163.367
R622 B.n43 B.n42 163.367
R623 B.n430 B.n43 163.367
R624 B.n430 B.n48 163.367
R625 B.n49 B.n48 163.367
R626 B.n50 B.n49 163.367
R627 B.n435 B.n50 163.367
R628 B.n435 B.n55 163.367
R629 B.n56 B.n55 163.367
R630 B.n57 B.n56 163.367
R631 B.n440 B.n57 163.367
R632 B.n440 B.n62 163.367
R633 B.n63 B.n62 163.367
R634 B.n64 B.n63 163.367
R635 B.n294 B.n292 163.367
R636 B.n292 B.n291 163.367
R637 B.n288 B.n287 163.367
R638 B.n285 B.n168 163.367
R639 B.n281 B.n279 163.367
R640 B.n277 B.n170 163.367
R641 B.n273 B.n271 163.367
R642 B.n269 B.n172 163.367
R643 B.n265 B.n263 163.367
R644 B.n261 B.n174 163.367
R645 B.n257 B.n255 163.367
R646 B.n252 B.n251 163.367
R647 B.n249 B.n180 163.367
R648 B.n245 B.n243 163.367
R649 B.n241 B.n182 163.367
R650 B.n237 B.n235 163.367
R651 B.n232 B.n231 163.367
R652 B.n229 B.n188 163.367
R653 B.n225 B.n223 163.367
R654 B.n221 B.n190 163.367
R655 B.n217 B.n215 163.367
R656 B.n213 B.n192 163.367
R657 B.n209 B.n207 163.367
R658 B.n205 B.n194 163.367
R659 B.n201 B.n199 163.367
R660 B.n197 B.n162 163.367
R661 B.n298 B.n158 163.367
R662 B.n306 B.n158 163.367
R663 B.n306 B.n156 163.367
R664 B.n310 B.n156 163.367
R665 B.n310 B.n150 163.367
R666 B.n318 B.n150 163.367
R667 B.n318 B.n148 163.367
R668 B.n322 B.n148 163.367
R669 B.n322 B.n142 163.367
R670 B.n330 B.n142 163.367
R671 B.n330 B.n140 163.367
R672 B.n334 B.n140 163.367
R673 B.n334 B.n134 163.367
R674 B.n342 B.n134 163.367
R675 B.n342 B.n132 163.367
R676 B.n346 B.n132 163.367
R677 B.n346 B.n126 163.367
R678 B.n354 B.n126 163.367
R679 B.n354 B.n124 163.367
R680 B.n358 B.n124 163.367
R681 B.n358 B.n118 163.367
R682 B.n366 B.n118 163.367
R683 B.n366 B.n116 163.367
R684 B.n370 B.n116 163.367
R685 B.n370 B.n110 163.367
R686 B.n378 B.n110 163.367
R687 B.n378 B.n108 163.367
R688 B.n382 B.n108 163.367
R689 B.n382 B.n102 163.367
R690 B.n391 B.n102 163.367
R691 B.n391 B.n100 163.367
R692 B.n395 B.n100 163.367
R693 B.n395 B.n3 163.367
R694 B.n620 B.n3 163.367
R695 B.n616 B.n2 163.367
R696 B.n616 B.n615 163.367
R697 B.n615 B.n9 163.367
R698 B.n611 B.n9 163.367
R699 B.n611 B.n11 163.367
R700 B.n607 B.n11 163.367
R701 B.n607 B.n17 163.367
R702 B.n603 B.n17 163.367
R703 B.n603 B.n19 163.367
R704 B.n599 B.n19 163.367
R705 B.n599 B.n24 163.367
R706 B.n595 B.n24 163.367
R707 B.n595 B.n26 163.367
R708 B.n591 B.n26 163.367
R709 B.n591 B.n31 163.367
R710 B.n587 B.n31 163.367
R711 B.n587 B.n33 163.367
R712 B.n583 B.n33 163.367
R713 B.n583 B.n38 163.367
R714 B.n579 B.n38 163.367
R715 B.n579 B.n40 163.367
R716 B.n575 B.n40 163.367
R717 B.n575 B.n45 163.367
R718 B.n571 B.n45 163.367
R719 B.n571 B.n47 163.367
R720 B.n567 B.n47 163.367
R721 B.n567 B.n52 163.367
R722 B.n563 B.n52 163.367
R723 B.n563 B.n54 163.367
R724 B.n559 B.n54 163.367
R725 B.n559 B.n59 163.367
R726 B.n555 B.n59 163.367
R727 B.n555 B.n61 163.367
R728 B.n551 B.n61 163.367
R729 B.n299 B.n163 146.24
R730 B.n552 B.n65 146.24
R731 B.n85 B.t8 119.231
R732 B.n183 B.t19 119.231
R733 B.n77 B.t15 119.227
R734 B.n175 B.t13 119.227
R735 B.n86 B.t9 75.4007
R736 B.n184 B.t18 75.4007
R737 B.n78 B.t16 75.3958
R738 B.n176 B.t12 75.3958
R739 B.n299 B.n159 72.5866
R740 B.n305 B.n159 72.5866
R741 B.n305 B.n155 72.5866
R742 B.n311 B.n155 72.5866
R743 B.n311 B.n151 72.5866
R744 B.n317 B.n151 72.5866
R745 B.n323 B.n147 72.5866
R746 B.n323 B.n143 72.5866
R747 B.n329 B.n143 72.5866
R748 B.n329 B.n139 72.5866
R749 B.n335 B.n139 72.5866
R750 B.n335 B.n135 72.5866
R751 B.n341 B.n135 72.5866
R752 B.n341 B.n131 72.5866
R753 B.n347 B.n131 72.5866
R754 B.n353 B.n127 72.5866
R755 B.n353 B.n123 72.5866
R756 B.n359 B.n123 72.5866
R757 B.n359 B.n119 72.5866
R758 B.n365 B.n119 72.5866
R759 B.n371 B.n115 72.5866
R760 B.n371 B.n111 72.5866
R761 B.n377 B.n111 72.5866
R762 B.n377 B.n106 72.5866
R763 B.n383 B.n106 72.5866
R764 B.n383 B.n107 72.5866
R765 B.n390 B.n99 72.5866
R766 B.n396 B.n99 72.5866
R767 B.n396 B.n4 72.5866
R768 B.n619 B.n4 72.5866
R769 B.n619 B.n618 72.5866
R770 B.n618 B.n617 72.5866
R771 B.n617 B.n8 72.5866
R772 B.n12 B.n8 72.5866
R773 B.n610 B.n12 72.5866
R774 B.n609 B.n608 72.5866
R775 B.n608 B.n16 72.5866
R776 B.n602 B.n16 72.5866
R777 B.n602 B.n601 72.5866
R778 B.n601 B.n600 72.5866
R779 B.n600 B.n23 72.5866
R780 B.n594 B.n593 72.5866
R781 B.n593 B.n592 72.5866
R782 B.n592 B.n30 72.5866
R783 B.n586 B.n30 72.5866
R784 B.n586 B.n585 72.5866
R785 B.n584 B.n37 72.5866
R786 B.n578 B.n37 72.5866
R787 B.n578 B.n577 72.5866
R788 B.n577 B.n576 72.5866
R789 B.n576 B.n44 72.5866
R790 B.n570 B.n44 72.5866
R791 B.n570 B.n569 72.5866
R792 B.n569 B.n568 72.5866
R793 B.n568 B.n51 72.5866
R794 B.n562 B.n561 72.5866
R795 B.n561 B.n560 72.5866
R796 B.n560 B.n58 72.5866
R797 B.n554 B.n58 72.5866
R798 B.n554 B.n553 72.5866
R799 B.n553 B.n552 72.5866
R800 B.n546 B.n66 71.676
R801 B.n545 B.n544 71.676
R802 B.n538 B.n68 71.676
R803 B.n537 B.n536 71.676
R804 B.n530 B.n70 71.676
R805 B.n529 B.n528 71.676
R806 B.n522 B.n72 71.676
R807 B.n521 B.n520 71.676
R808 B.n514 B.n74 71.676
R809 B.n513 B.n512 71.676
R810 B.n505 B.n76 71.676
R811 B.n504 B.n503 71.676
R812 B.n497 B.n80 71.676
R813 B.n496 B.n495 71.676
R814 B.n489 B.n82 71.676
R815 B.n488 B.n487 71.676
R816 B.n481 B.n84 71.676
R817 B.n480 B.n479 71.676
R818 B.n473 B.n89 71.676
R819 B.n472 B.n471 71.676
R820 B.n465 B.n91 71.676
R821 B.n464 B.n463 71.676
R822 B.n457 B.n93 71.676
R823 B.n456 B.n455 71.676
R824 B.n449 B.n95 71.676
R825 B.n448 B.n447 71.676
R826 B.n447 B.n446 71.676
R827 B.n450 B.n449 71.676
R828 B.n455 B.n454 71.676
R829 B.n458 B.n457 71.676
R830 B.n463 B.n462 71.676
R831 B.n466 B.n465 71.676
R832 B.n471 B.n470 71.676
R833 B.n474 B.n473 71.676
R834 B.n479 B.n478 71.676
R835 B.n482 B.n481 71.676
R836 B.n487 B.n486 71.676
R837 B.n490 B.n489 71.676
R838 B.n495 B.n494 71.676
R839 B.n498 B.n497 71.676
R840 B.n503 B.n502 71.676
R841 B.n506 B.n505 71.676
R842 B.n512 B.n511 71.676
R843 B.n515 B.n514 71.676
R844 B.n520 B.n519 71.676
R845 B.n523 B.n522 71.676
R846 B.n528 B.n527 71.676
R847 B.n531 B.n530 71.676
R848 B.n536 B.n535 71.676
R849 B.n539 B.n538 71.676
R850 B.n544 B.n543 71.676
R851 B.n547 B.n546 71.676
R852 B.n293 B.n164 71.676
R853 B.n291 B.n166 71.676
R854 B.n287 B.n286 71.676
R855 B.n280 B.n168 71.676
R856 B.n279 B.n278 71.676
R857 B.n272 B.n170 71.676
R858 B.n271 B.n270 71.676
R859 B.n264 B.n172 71.676
R860 B.n263 B.n262 71.676
R861 B.n256 B.n174 71.676
R862 B.n255 B.n178 71.676
R863 B.n251 B.n250 71.676
R864 B.n244 B.n180 71.676
R865 B.n243 B.n242 71.676
R866 B.n236 B.n182 71.676
R867 B.n235 B.n186 71.676
R868 B.n231 B.n230 71.676
R869 B.n224 B.n188 71.676
R870 B.n223 B.n222 71.676
R871 B.n216 B.n190 71.676
R872 B.n215 B.n214 71.676
R873 B.n208 B.n192 71.676
R874 B.n207 B.n206 71.676
R875 B.n200 B.n194 71.676
R876 B.n199 B.n198 71.676
R877 B.n294 B.n293 71.676
R878 B.n288 B.n166 71.676
R879 B.n286 B.n285 71.676
R880 B.n281 B.n280 71.676
R881 B.n278 B.n277 71.676
R882 B.n273 B.n272 71.676
R883 B.n270 B.n269 71.676
R884 B.n265 B.n264 71.676
R885 B.n262 B.n261 71.676
R886 B.n257 B.n256 71.676
R887 B.n252 B.n178 71.676
R888 B.n250 B.n249 71.676
R889 B.n245 B.n244 71.676
R890 B.n242 B.n241 71.676
R891 B.n237 B.n236 71.676
R892 B.n232 B.n186 71.676
R893 B.n230 B.n229 71.676
R894 B.n225 B.n224 71.676
R895 B.n222 B.n221 71.676
R896 B.n217 B.n216 71.676
R897 B.n214 B.n213 71.676
R898 B.n209 B.n208 71.676
R899 B.n206 B.n205 71.676
R900 B.n201 B.n200 71.676
R901 B.n198 B.n197 71.676
R902 B.n621 B.n620 71.676
R903 B.n621 B.n2 71.676
R904 B.n365 B.t5 67.2494
R905 B.n594 B.t2 67.2494
R906 B.n508 B.n78 59.5399
R907 B.n87 B.n86 59.5399
R908 B.n185 B.n184 59.5399
R909 B.n177 B.n176 59.5399
R910 B.t0 B.n127 52.3052
R911 B.n585 B.t4 52.3052
R912 B.n78 B.n77 43.8308
R913 B.n86 B.n85 43.8308
R914 B.n184 B.n183 43.8308
R915 B.n176 B.n175 43.8308
R916 B.t11 B.n147 41.6308
R917 B.n107 B.t3 41.6308
R918 B.t1 B.n609 41.6308
R919 B.t7 B.n51 41.6308
R920 B.n297 B.n296 33.5615
R921 B.n301 B.n161 33.5615
R922 B.n445 B.n444 33.5615
R923 B.n550 B.n549 33.5615
R924 B.n317 B.t11 30.9563
R925 B.n390 B.t3 30.9563
R926 B.n610 B.t1 30.9563
R927 B.n562 B.t7 30.9563
R928 B.n347 B.t0 20.2819
R929 B.t4 B.n584 20.2819
R930 B B.n622 18.0485
R931 B.n297 B.n157 10.6151
R932 B.n307 B.n157 10.6151
R933 B.n308 B.n307 10.6151
R934 B.n309 B.n308 10.6151
R935 B.n309 B.n149 10.6151
R936 B.n319 B.n149 10.6151
R937 B.n320 B.n319 10.6151
R938 B.n321 B.n320 10.6151
R939 B.n321 B.n141 10.6151
R940 B.n331 B.n141 10.6151
R941 B.n332 B.n331 10.6151
R942 B.n333 B.n332 10.6151
R943 B.n333 B.n133 10.6151
R944 B.n343 B.n133 10.6151
R945 B.n344 B.n343 10.6151
R946 B.n345 B.n344 10.6151
R947 B.n345 B.n125 10.6151
R948 B.n355 B.n125 10.6151
R949 B.n356 B.n355 10.6151
R950 B.n357 B.n356 10.6151
R951 B.n357 B.n117 10.6151
R952 B.n367 B.n117 10.6151
R953 B.n368 B.n367 10.6151
R954 B.n369 B.n368 10.6151
R955 B.n369 B.n109 10.6151
R956 B.n379 B.n109 10.6151
R957 B.n380 B.n379 10.6151
R958 B.n381 B.n380 10.6151
R959 B.n381 B.n101 10.6151
R960 B.n392 B.n101 10.6151
R961 B.n393 B.n392 10.6151
R962 B.n394 B.n393 10.6151
R963 B.n394 B.n0 10.6151
R964 B.n296 B.n295 10.6151
R965 B.n295 B.n165 10.6151
R966 B.n290 B.n165 10.6151
R967 B.n290 B.n289 10.6151
R968 B.n289 B.n167 10.6151
R969 B.n284 B.n167 10.6151
R970 B.n284 B.n283 10.6151
R971 B.n283 B.n282 10.6151
R972 B.n282 B.n169 10.6151
R973 B.n276 B.n169 10.6151
R974 B.n276 B.n275 10.6151
R975 B.n275 B.n274 10.6151
R976 B.n274 B.n171 10.6151
R977 B.n268 B.n171 10.6151
R978 B.n268 B.n267 10.6151
R979 B.n267 B.n266 10.6151
R980 B.n266 B.n173 10.6151
R981 B.n260 B.n173 10.6151
R982 B.n260 B.n259 10.6151
R983 B.n259 B.n258 10.6151
R984 B.n254 B.n253 10.6151
R985 B.n253 B.n179 10.6151
R986 B.n248 B.n179 10.6151
R987 B.n248 B.n247 10.6151
R988 B.n247 B.n246 10.6151
R989 B.n246 B.n181 10.6151
R990 B.n240 B.n181 10.6151
R991 B.n240 B.n239 10.6151
R992 B.n239 B.n238 10.6151
R993 B.n234 B.n233 10.6151
R994 B.n233 B.n187 10.6151
R995 B.n228 B.n187 10.6151
R996 B.n228 B.n227 10.6151
R997 B.n227 B.n226 10.6151
R998 B.n226 B.n189 10.6151
R999 B.n220 B.n189 10.6151
R1000 B.n220 B.n219 10.6151
R1001 B.n219 B.n218 10.6151
R1002 B.n218 B.n191 10.6151
R1003 B.n212 B.n191 10.6151
R1004 B.n212 B.n211 10.6151
R1005 B.n211 B.n210 10.6151
R1006 B.n210 B.n193 10.6151
R1007 B.n204 B.n193 10.6151
R1008 B.n204 B.n203 10.6151
R1009 B.n203 B.n202 10.6151
R1010 B.n202 B.n195 10.6151
R1011 B.n196 B.n195 10.6151
R1012 B.n196 B.n161 10.6151
R1013 B.n302 B.n301 10.6151
R1014 B.n303 B.n302 10.6151
R1015 B.n303 B.n153 10.6151
R1016 B.n313 B.n153 10.6151
R1017 B.n314 B.n313 10.6151
R1018 B.n315 B.n314 10.6151
R1019 B.n315 B.n145 10.6151
R1020 B.n325 B.n145 10.6151
R1021 B.n326 B.n325 10.6151
R1022 B.n327 B.n326 10.6151
R1023 B.n327 B.n137 10.6151
R1024 B.n337 B.n137 10.6151
R1025 B.n338 B.n337 10.6151
R1026 B.n339 B.n338 10.6151
R1027 B.n339 B.n129 10.6151
R1028 B.n349 B.n129 10.6151
R1029 B.n350 B.n349 10.6151
R1030 B.n351 B.n350 10.6151
R1031 B.n351 B.n121 10.6151
R1032 B.n361 B.n121 10.6151
R1033 B.n362 B.n361 10.6151
R1034 B.n363 B.n362 10.6151
R1035 B.n363 B.n113 10.6151
R1036 B.n373 B.n113 10.6151
R1037 B.n374 B.n373 10.6151
R1038 B.n375 B.n374 10.6151
R1039 B.n375 B.n104 10.6151
R1040 B.n385 B.n104 10.6151
R1041 B.n386 B.n385 10.6151
R1042 B.n388 B.n386 10.6151
R1043 B.n388 B.n387 10.6151
R1044 B.n387 B.n97 10.6151
R1045 B.n399 B.n97 10.6151
R1046 B.n400 B.n399 10.6151
R1047 B.n401 B.n400 10.6151
R1048 B.n402 B.n401 10.6151
R1049 B.n403 B.n402 10.6151
R1050 B.n406 B.n403 10.6151
R1051 B.n407 B.n406 10.6151
R1052 B.n408 B.n407 10.6151
R1053 B.n409 B.n408 10.6151
R1054 B.n411 B.n409 10.6151
R1055 B.n412 B.n411 10.6151
R1056 B.n413 B.n412 10.6151
R1057 B.n414 B.n413 10.6151
R1058 B.n416 B.n414 10.6151
R1059 B.n417 B.n416 10.6151
R1060 B.n418 B.n417 10.6151
R1061 B.n419 B.n418 10.6151
R1062 B.n421 B.n419 10.6151
R1063 B.n422 B.n421 10.6151
R1064 B.n423 B.n422 10.6151
R1065 B.n424 B.n423 10.6151
R1066 B.n426 B.n424 10.6151
R1067 B.n427 B.n426 10.6151
R1068 B.n428 B.n427 10.6151
R1069 B.n429 B.n428 10.6151
R1070 B.n431 B.n429 10.6151
R1071 B.n432 B.n431 10.6151
R1072 B.n433 B.n432 10.6151
R1073 B.n434 B.n433 10.6151
R1074 B.n436 B.n434 10.6151
R1075 B.n437 B.n436 10.6151
R1076 B.n438 B.n437 10.6151
R1077 B.n439 B.n438 10.6151
R1078 B.n441 B.n439 10.6151
R1079 B.n442 B.n441 10.6151
R1080 B.n443 B.n442 10.6151
R1081 B.n444 B.n443 10.6151
R1082 B.n614 B.n1 10.6151
R1083 B.n614 B.n613 10.6151
R1084 B.n613 B.n612 10.6151
R1085 B.n612 B.n10 10.6151
R1086 B.n606 B.n10 10.6151
R1087 B.n606 B.n605 10.6151
R1088 B.n605 B.n604 10.6151
R1089 B.n604 B.n18 10.6151
R1090 B.n598 B.n18 10.6151
R1091 B.n598 B.n597 10.6151
R1092 B.n597 B.n596 10.6151
R1093 B.n596 B.n25 10.6151
R1094 B.n590 B.n25 10.6151
R1095 B.n590 B.n589 10.6151
R1096 B.n589 B.n588 10.6151
R1097 B.n588 B.n32 10.6151
R1098 B.n582 B.n32 10.6151
R1099 B.n582 B.n581 10.6151
R1100 B.n581 B.n580 10.6151
R1101 B.n580 B.n39 10.6151
R1102 B.n574 B.n39 10.6151
R1103 B.n574 B.n573 10.6151
R1104 B.n573 B.n572 10.6151
R1105 B.n572 B.n46 10.6151
R1106 B.n566 B.n46 10.6151
R1107 B.n566 B.n565 10.6151
R1108 B.n565 B.n564 10.6151
R1109 B.n564 B.n53 10.6151
R1110 B.n558 B.n53 10.6151
R1111 B.n558 B.n557 10.6151
R1112 B.n557 B.n556 10.6151
R1113 B.n556 B.n60 10.6151
R1114 B.n550 B.n60 10.6151
R1115 B.n549 B.n548 10.6151
R1116 B.n548 B.n67 10.6151
R1117 B.n542 B.n67 10.6151
R1118 B.n542 B.n541 10.6151
R1119 B.n541 B.n540 10.6151
R1120 B.n540 B.n69 10.6151
R1121 B.n534 B.n69 10.6151
R1122 B.n534 B.n533 10.6151
R1123 B.n533 B.n532 10.6151
R1124 B.n532 B.n71 10.6151
R1125 B.n526 B.n71 10.6151
R1126 B.n526 B.n525 10.6151
R1127 B.n525 B.n524 10.6151
R1128 B.n524 B.n73 10.6151
R1129 B.n518 B.n73 10.6151
R1130 B.n518 B.n517 10.6151
R1131 B.n517 B.n516 10.6151
R1132 B.n516 B.n75 10.6151
R1133 B.n510 B.n75 10.6151
R1134 B.n510 B.n509 10.6151
R1135 B.n507 B.n79 10.6151
R1136 B.n501 B.n79 10.6151
R1137 B.n501 B.n500 10.6151
R1138 B.n500 B.n499 10.6151
R1139 B.n499 B.n81 10.6151
R1140 B.n493 B.n81 10.6151
R1141 B.n493 B.n492 10.6151
R1142 B.n492 B.n491 10.6151
R1143 B.n491 B.n83 10.6151
R1144 B.n485 B.n484 10.6151
R1145 B.n484 B.n483 10.6151
R1146 B.n483 B.n88 10.6151
R1147 B.n477 B.n88 10.6151
R1148 B.n477 B.n476 10.6151
R1149 B.n476 B.n475 10.6151
R1150 B.n475 B.n90 10.6151
R1151 B.n469 B.n90 10.6151
R1152 B.n469 B.n468 10.6151
R1153 B.n468 B.n467 10.6151
R1154 B.n467 B.n92 10.6151
R1155 B.n461 B.n92 10.6151
R1156 B.n461 B.n460 10.6151
R1157 B.n460 B.n459 10.6151
R1158 B.n459 B.n94 10.6151
R1159 B.n453 B.n94 10.6151
R1160 B.n453 B.n452 10.6151
R1161 B.n452 B.n451 10.6151
R1162 B.n451 B.n96 10.6151
R1163 B.n445 B.n96 10.6151
R1164 B.n258 B.n177 9.36635
R1165 B.n234 B.n185 9.36635
R1166 B.n509 B.n508 9.36635
R1167 B.n485 B.n87 9.36635
R1168 B.n622 B.n0 8.11757
R1169 B.n622 B.n1 8.11757
R1170 B.t5 B.n115 5.33771
R1171 B.t2 B.n23 5.33771
R1172 B.n254 B.n177 1.24928
R1173 B.n238 B.n185 1.24928
R1174 B.n508 B.n507 1.24928
R1175 B.n87 B.n83 1.24928
R1176 VN.n13 VN.n12 185.279
R1177 VN.n27 VN.n26 185.279
R1178 VN.n25 VN.n14 161.3
R1179 VN.n24 VN.n23 161.3
R1180 VN.n22 VN.n15 161.3
R1181 VN.n21 VN.n20 161.3
R1182 VN.n19 VN.n16 161.3
R1183 VN.n11 VN.n0 161.3
R1184 VN.n10 VN.n9 161.3
R1185 VN.n8 VN.n1 161.3
R1186 VN.n7 VN.n6 161.3
R1187 VN.n5 VN.n2 161.3
R1188 VN.n3 VN.t5 94.5642
R1189 VN.n17 VN.t2 94.5642
R1190 VN.n4 VN.t3 62.8103
R1191 VN.n12 VN.t1 62.8103
R1192 VN.n18 VN.t0 62.8103
R1193 VN.n26 VN.t4 62.8103
R1194 VN.n4 VN.n3 57.9196
R1195 VN.n18 VN.n17 57.9196
R1196 VN.n6 VN.n1 52.1486
R1197 VN.n20 VN.n15 52.1486
R1198 VN VN.n27 41.0327
R1199 VN.n10 VN.n1 28.8382
R1200 VN.n24 VN.n15 28.8382
R1201 VN.n6 VN.n5 24.4675
R1202 VN.n11 VN.n10 24.4675
R1203 VN.n20 VN.n19 24.4675
R1204 VN.n25 VN.n24 24.4675
R1205 VN.n17 VN.n16 12.5909
R1206 VN.n3 VN.n2 12.5909
R1207 VN.n5 VN.n4 12.234
R1208 VN.n19 VN.n18 12.234
R1209 VN.n12 VN.n11 0.48984
R1210 VN.n26 VN.n25 0.48984
R1211 VN.n27 VN.n14 0.189894
R1212 VN.n23 VN.n14 0.189894
R1213 VN.n23 VN.n22 0.189894
R1214 VN.n22 VN.n21 0.189894
R1215 VN.n21 VN.n16 0.189894
R1216 VN.n7 VN.n2 0.189894
R1217 VN.n8 VN.n7 0.189894
R1218 VN.n9 VN.n8 0.189894
R1219 VN.n9 VN.n0 0.189894
R1220 VN.n13 VN.n0 0.189894
R1221 VN VN.n13 0.0516364
R1222 VDD2.n1 VDD2.t0 77.0425
R1223 VDD2.n2 VDD2.t1 75.6367
R1224 VDD2.n1 VDD2.n0 72.1319
R1225 VDD2 VDD2.n3 72.1291
R1226 VDD2.n2 VDD2.n1 34.3834
R1227 VDD2.n3 VDD2.t5 3.93688
R1228 VDD2.n3 VDD2.t3 3.93688
R1229 VDD2.n0 VDD2.t2 3.93688
R1230 VDD2.n0 VDD2.t4 3.93688
R1231 VDD2 VDD2.n2 1.5199
C0 VN VDD2 2.85856f
C1 VP VDD1 3.10762f
C2 VTAIL VDD2 4.94506f
C3 VN VTAIL 3.27873f
C4 VP VDD2 0.405001f
C5 VDD1 VDD2 1.16894f
C6 VP VN 4.98421f
C7 VP VTAIL 3.29294f
C8 VN VDD1 0.149807f
C9 VTAIL VDD1 4.89748f
C10 VDD2 B 4.195135f
C11 VDD1 B 4.48169f
C12 VTAIL B 4.365514f
C13 VN B 10.244649f
C14 VP B 8.854128f
C15 VDD2.t0 B 0.912828f
C16 VDD2.t2 B 0.087497f
C17 VDD2.t4 B 0.087497f
C18 VDD2.n0 B 0.715291f
C19 VDD2.n1 B 1.91408f
C20 VDD2.t1 B 0.906822f
C21 VDD2.n2 B 1.79676f
C22 VDD2.t5 B 0.087497f
C23 VDD2.t3 B 0.087497f
C24 VDD2.n3 B 0.715268f
C25 VN.n0 B 0.031583f
C26 VN.t1 B 0.802301f
C27 VN.n1 B 0.0319f
C28 VN.n2 B 0.234447f
C29 VN.t3 B 0.802301f
C30 VN.t5 B 0.960767f
C31 VN.n3 B 0.388797f
C32 VN.n4 B 0.389303f
C33 VN.n5 B 0.044332f
C34 VN.n6 B 0.0567f
C35 VN.n7 B 0.031583f
C36 VN.n8 B 0.031583f
C37 VN.n9 B 0.031583f
C38 VN.n10 B 0.062472f
C39 VN.n11 B 0.030383f
C40 VN.n12 B 0.388983f
C41 VN.n13 B 0.035403f
C42 VN.n14 B 0.031583f
C43 VN.t4 B 0.802301f
C44 VN.n15 B 0.0319f
C45 VN.n16 B 0.234447f
C46 VN.t0 B 0.802301f
C47 VN.t2 B 0.960767f
C48 VN.n17 B 0.388797f
C49 VN.n18 B 0.389303f
C50 VN.n19 B 0.044332f
C51 VN.n20 B 0.0567f
C52 VN.n21 B 0.031583f
C53 VN.n22 B 0.031583f
C54 VN.n23 B 0.031583f
C55 VN.n24 B 0.062472f
C56 VN.n25 B 0.030383f
C57 VN.n26 B 0.388983f
C58 VN.n27 B 1.2656f
C59 VDD1.t0 B 0.927216f
C60 VDD1.t5 B 0.926576f
C61 VDD1.t4 B 0.088815f
C62 VDD1.t3 B 0.088815f
C63 VDD1.n0 B 0.726064f
C64 VDD1.n1 B 2.0334f
C65 VDD1.t1 B 0.088815f
C66 VDD1.t2 B 0.088815f
C67 VDD1.n2 B 0.723911f
C68 VDD1.n3 B 1.83195f
C69 VTAIL.t1 B 0.107938f
C70 VTAIL.t2 B 0.107938f
C71 VTAIL.n0 B 0.815751f
C72 VTAIL.n1 B 0.417535f
C73 VTAIL.t9 B 1.04321f
C74 VTAIL.n2 B 0.607213f
C75 VTAIL.t8 B 0.107938f
C76 VTAIL.t11 B 0.107938f
C77 VTAIL.n3 B 0.815751f
C78 VTAIL.n4 B 1.50319f
C79 VTAIL.t0 B 0.107938f
C80 VTAIL.t5 B 0.107938f
C81 VTAIL.n5 B 0.815755f
C82 VTAIL.n6 B 1.50318f
C83 VTAIL.t3 B 1.04322f
C84 VTAIL.n7 B 0.607206f
C85 VTAIL.t6 B 0.107938f
C86 VTAIL.t7 B 0.107938f
C87 VTAIL.n8 B 0.815755f
C88 VTAIL.n9 B 0.540295f
C89 VTAIL.t10 B 1.04321f
C90 VTAIL.n10 B 1.39963f
C91 VTAIL.t4 B 1.04321f
C92 VTAIL.n11 B 1.35192f
C93 VP.n0 B 0.032275f
C94 VP.t2 B 0.819878f
C95 VP.n1 B 0.032599f
C96 VP.n2 B 0.032275f
C97 VP.t1 B 0.819878f
C98 VP.n3 B 0.057942f
C99 VP.n4 B 0.032275f
C100 VP.t0 B 0.819878f
C101 VP.n5 B 0.397505f
C102 VP.n6 B 0.032275f
C103 VP.t3 B 0.819878f
C104 VP.n7 B 0.032599f
C105 VP.n8 B 0.239584f
C106 VP.t4 B 0.819878f
C107 VP.t5 B 0.981815f
C108 VP.n9 B 0.397315f
C109 VP.n10 B 0.397832f
C110 VP.n11 B 0.045303f
C111 VP.n12 B 0.057942f
C112 VP.n13 B 0.032275f
C113 VP.n14 B 0.032275f
C114 VP.n15 B 0.032275f
C115 VP.n16 B 0.063841f
C116 VP.n17 B 0.031048f
C117 VP.n18 B 0.397505f
C118 VP.n19 B 1.27209f
C119 VP.n20 B 1.30063f
C120 VP.n21 B 0.032275f
C121 VP.n22 B 0.031048f
C122 VP.n23 B 0.063841f
C123 VP.n24 B 0.032599f
C124 VP.n25 B 0.032275f
C125 VP.n26 B 0.032275f
C126 VP.n27 B 0.032275f
C127 VP.n28 B 0.045303f
C128 VP.n29 B 0.322386f
C129 VP.n30 B 0.045303f
C130 VP.n31 B 0.057942f
C131 VP.n32 B 0.032275f
C132 VP.n33 B 0.032275f
C133 VP.n34 B 0.032275f
C134 VP.n35 B 0.063841f
C135 VP.n36 B 0.031048f
C136 VP.n37 B 0.397505f
C137 VP.n38 B 0.036178f
.ends

