* NGSPICE file created from diff_pair_sample_0658.ext - technology: sky130A

.subckt diff_pair_sample_0658 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2034_n1242# sky130_fd_pr__pfet_01v8 ad=0.5343 pd=3.52 as=0 ps=0 w=1.37 l=2.33
X1 B.t8 B.t6 B.t7 w_n2034_n1242# sky130_fd_pr__pfet_01v8 ad=0.5343 pd=3.52 as=0 ps=0 w=1.37 l=2.33
X2 VDD2.t1 VN.t0 VTAIL.t3 w_n2034_n1242# sky130_fd_pr__pfet_01v8 ad=0.5343 pd=3.52 as=0.5343 ps=3.52 w=1.37 l=2.33
X3 VDD2.t0 VN.t1 VTAIL.t2 w_n2034_n1242# sky130_fd_pr__pfet_01v8 ad=0.5343 pd=3.52 as=0.5343 ps=3.52 w=1.37 l=2.33
X4 B.t5 B.t3 B.t4 w_n2034_n1242# sky130_fd_pr__pfet_01v8 ad=0.5343 pd=3.52 as=0 ps=0 w=1.37 l=2.33
X5 B.t2 B.t0 B.t1 w_n2034_n1242# sky130_fd_pr__pfet_01v8 ad=0.5343 pd=3.52 as=0 ps=0 w=1.37 l=2.33
X6 VDD1.t1 VP.t0 VTAIL.t1 w_n2034_n1242# sky130_fd_pr__pfet_01v8 ad=0.5343 pd=3.52 as=0.5343 ps=3.52 w=1.37 l=2.33
X7 VDD1.t0 VP.t1 VTAIL.t0 w_n2034_n1242# sky130_fd_pr__pfet_01v8 ad=0.5343 pd=3.52 as=0.5343 ps=3.52 w=1.37 l=2.33
R0 B.n167 B.n166 585
R1 B.n165 B.n58 585
R2 B.n164 B.n163 585
R3 B.n162 B.n59 585
R4 B.n161 B.n160 585
R5 B.n159 B.n60 585
R6 B.n158 B.n157 585
R7 B.n156 B.n61 585
R8 B.n155 B.n154 585
R9 B.n153 B.n62 585
R10 B.n151 B.n150 585
R11 B.n149 B.n65 585
R12 B.n148 B.n147 585
R13 B.n146 B.n66 585
R14 B.n145 B.n144 585
R15 B.n143 B.n67 585
R16 B.n142 B.n141 585
R17 B.n140 B.n68 585
R18 B.n139 B.n138 585
R19 B.n137 B.n69 585
R20 B.n136 B.n135 585
R21 B.n131 B.n70 585
R22 B.n130 B.n129 585
R23 B.n128 B.n71 585
R24 B.n127 B.n126 585
R25 B.n125 B.n72 585
R26 B.n124 B.n123 585
R27 B.n122 B.n73 585
R28 B.n121 B.n120 585
R29 B.n119 B.n74 585
R30 B.n168 B.n57 585
R31 B.n170 B.n169 585
R32 B.n171 B.n56 585
R33 B.n173 B.n172 585
R34 B.n174 B.n55 585
R35 B.n176 B.n175 585
R36 B.n177 B.n54 585
R37 B.n179 B.n178 585
R38 B.n180 B.n53 585
R39 B.n182 B.n181 585
R40 B.n183 B.n52 585
R41 B.n185 B.n184 585
R42 B.n186 B.n51 585
R43 B.n188 B.n187 585
R44 B.n189 B.n50 585
R45 B.n191 B.n190 585
R46 B.n192 B.n49 585
R47 B.n194 B.n193 585
R48 B.n195 B.n48 585
R49 B.n197 B.n196 585
R50 B.n198 B.n47 585
R51 B.n200 B.n199 585
R52 B.n201 B.n46 585
R53 B.n203 B.n202 585
R54 B.n204 B.n45 585
R55 B.n206 B.n205 585
R56 B.n207 B.n44 585
R57 B.n209 B.n208 585
R58 B.n210 B.n43 585
R59 B.n212 B.n211 585
R60 B.n213 B.n42 585
R61 B.n215 B.n214 585
R62 B.n216 B.n41 585
R63 B.n218 B.n217 585
R64 B.n219 B.n40 585
R65 B.n221 B.n220 585
R66 B.n222 B.n39 585
R67 B.n224 B.n223 585
R68 B.n225 B.n38 585
R69 B.n227 B.n226 585
R70 B.n228 B.n37 585
R71 B.n230 B.n229 585
R72 B.n231 B.n36 585
R73 B.n233 B.n232 585
R74 B.n234 B.n35 585
R75 B.n236 B.n235 585
R76 B.n237 B.n34 585
R77 B.n239 B.n238 585
R78 B.n285 B.n284 585
R79 B.n283 B.n14 585
R80 B.n282 B.n281 585
R81 B.n280 B.n15 585
R82 B.n279 B.n278 585
R83 B.n277 B.n16 585
R84 B.n276 B.n275 585
R85 B.n274 B.n17 585
R86 B.n273 B.n272 585
R87 B.n271 B.n18 585
R88 B.n270 B.n269 585
R89 B.n268 B.n19 585
R90 B.n267 B.n266 585
R91 B.n265 B.n23 585
R92 B.n264 B.n263 585
R93 B.n262 B.n24 585
R94 B.n261 B.n260 585
R95 B.n259 B.n25 585
R96 B.n258 B.n257 585
R97 B.n256 B.n26 585
R98 B.n254 B.n253 585
R99 B.n252 B.n29 585
R100 B.n251 B.n250 585
R101 B.n249 B.n30 585
R102 B.n248 B.n247 585
R103 B.n246 B.n31 585
R104 B.n245 B.n244 585
R105 B.n243 B.n32 585
R106 B.n242 B.n241 585
R107 B.n240 B.n33 585
R108 B.n286 B.n13 585
R109 B.n288 B.n287 585
R110 B.n289 B.n12 585
R111 B.n291 B.n290 585
R112 B.n292 B.n11 585
R113 B.n294 B.n293 585
R114 B.n295 B.n10 585
R115 B.n297 B.n296 585
R116 B.n298 B.n9 585
R117 B.n300 B.n299 585
R118 B.n301 B.n8 585
R119 B.n303 B.n302 585
R120 B.n304 B.n7 585
R121 B.n306 B.n305 585
R122 B.n307 B.n6 585
R123 B.n309 B.n308 585
R124 B.n310 B.n5 585
R125 B.n312 B.n311 585
R126 B.n313 B.n4 585
R127 B.n315 B.n314 585
R128 B.n316 B.n3 585
R129 B.n318 B.n317 585
R130 B.n319 B.n0 585
R131 B.n2 B.n1 585
R132 B.n86 B.n85 585
R133 B.n88 B.n87 585
R134 B.n89 B.n84 585
R135 B.n91 B.n90 585
R136 B.n92 B.n83 585
R137 B.n94 B.n93 585
R138 B.n95 B.n82 585
R139 B.n97 B.n96 585
R140 B.n98 B.n81 585
R141 B.n100 B.n99 585
R142 B.n101 B.n80 585
R143 B.n103 B.n102 585
R144 B.n104 B.n79 585
R145 B.n106 B.n105 585
R146 B.n107 B.n78 585
R147 B.n109 B.n108 585
R148 B.n110 B.n77 585
R149 B.n112 B.n111 585
R150 B.n113 B.n76 585
R151 B.n115 B.n114 585
R152 B.n116 B.n75 585
R153 B.n118 B.n117 585
R154 B.n117 B.n74 564.573
R155 B.n168 B.n167 564.573
R156 B.n240 B.n239 564.573
R157 B.n284 B.n13 564.573
R158 B.n63 B.t7 300.57
R159 B.n27 B.t5 300.57
R160 B.n132 B.t1 300.57
R161 B.n20 B.t11 300.57
R162 B.n321 B.n320 256.663
R163 B.n64 B.t8 248.982
R164 B.n28 B.t4 248.982
R165 B.n133 B.t2 248.982
R166 B.n21 B.t10 248.982
R167 B.n320 B.n319 235.042
R168 B.n320 B.n2 235.042
R169 B.n132 B.t0 221.77
R170 B.n63 B.t6 221.77
R171 B.n27 B.t3 221.77
R172 B.n20 B.t9 221.77
R173 B.n121 B.n74 163.367
R174 B.n122 B.n121 163.367
R175 B.n123 B.n122 163.367
R176 B.n123 B.n72 163.367
R177 B.n127 B.n72 163.367
R178 B.n128 B.n127 163.367
R179 B.n129 B.n128 163.367
R180 B.n129 B.n70 163.367
R181 B.n136 B.n70 163.367
R182 B.n137 B.n136 163.367
R183 B.n138 B.n137 163.367
R184 B.n138 B.n68 163.367
R185 B.n142 B.n68 163.367
R186 B.n143 B.n142 163.367
R187 B.n144 B.n143 163.367
R188 B.n144 B.n66 163.367
R189 B.n148 B.n66 163.367
R190 B.n149 B.n148 163.367
R191 B.n150 B.n149 163.367
R192 B.n150 B.n62 163.367
R193 B.n155 B.n62 163.367
R194 B.n156 B.n155 163.367
R195 B.n157 B.n156 163.367
R196 B.n157 B.n60 163.367
R197 B.n161 B.n60 163.367
R198 B.n162 B.n161 163.367
R199 B.n163 B.n162 163.367
R200 B.n163 B.n58 163.367
R201 B.n167 B.n58 163.367
R202 B.n239 B.n34 163.367
R203 B.n235 B.n34 163.367
R204 B.n235 B.n234 163.367
R205 B.n234 B.n233 163.367
R206 B.n233 B.n36 163.367
R207 B.n229 B.n36 163.367
R208 B.n229 B.n228 163.367
R209 B.n228 B.n227 163.367
R210 B.n227 B.n38 163.367
R211 B.n223 B.n38 163.367
R212 B.n223 B.n222 163.367
R213 B.n222 B.n221 163.367
R214 B.n221 B.n40 163.367
R215 B.n217 B.n40 163.367
R216 B.n217 B.n216 163.367
R217 B.n216 B.n215 163.367
R218 B.n215 B.n42 163.367
R219 B.n211 B.n42 163.367
R220 B.n211 B.n210 163.367
R221 B.n210 B.n209 163.367
R222 B.n209 B.n44 163.367
R223 B.n205 B.n44 163.367
R224 B.n205 B.n204 163.367
R225 B.n204 B.n203 163.367
R226 B.n203 B.n46 163.367
R227 B.n199 B.n46 163.367
R228 B.n199 B.n198 163.367
R229 B.n198 B.n197 163.367
R230 B.n197 B.n48 163.367
R231 B.n193 B.n48 163.367
R232 B.n193 B.n192 163.367
R233 B.n192 B.n191 163.367
R234 B.n191 B.n50 163.367
R235 B.n187 B.n50 163.367
R236 B.n187 B.n186 163.367
R237 B.n186 B.n185 163.367
R238 B.n185 B.n52 163.367
R239 B.n181 B.n52 163.367
R240 B.n181 B.n180 163.367
R241 B.n180 B.n179 163.367
R242 B.n179 B.n54 163.367
R243 B.n175 B.n54 163.367
R244 B.n175 B.n174 163.367
R245 B.n174 B.n173 163.367
R246 B.n173 B.n56 163.367
R247 B.n169 B.n56 163.367
R248 B.n169 B.n168 163.367
R249 B.n284 B.n283 163.367
R250 B.n283 B.n282 163.367
R251 B.n282 B.n15 163.367
R252 B.n278 B.n15 163.367
R253 B.n278 B.n277 163.367
R254 B.n277 B.n276 163.367
R255 B.n276 B.n17 163.367
R256 B.n272 B.n17 163.367
R257 B.n272 B.n271 163.367
R258 B.n271 B.n270 163.367
R259 B.n270 B.n19 163.367
R260 B.n266 B.n19 163.367
R261 B.n266 B.n265 163.367
R262 B.n265 B.n264 163.367
R263 B.n264 B.n24 163.367
R264 B.n260 B.n24 163.367
R265 B.n260 B.n259 163.367
R266 B.n259 B.n258 163.367
R267 B.n258 B.n26 163.367
R268 B.n253 B.n26 163.367
R269 B.n253 B.n252 163.367
R270 B.n252 B.n251 163.367
R271 B.n251 B.n30 163.367
R272 B.n247 B.n30 163.367
R273 B.n247 B.n246 163.367
R274 B.n246 B.n245 163.367
R275 B.n245 B.n32 163.367
R276 B.n241 B.n32 163.367
R277 B.n241 B.n240 163.367
R278 B.n288 B.n13 163.367
R279 B.n289 B.n288 163.367
R280 B.n290 B.n289 163.367
R281 B.n290 B.n11 163.367
R282 B.n294 B.n11 163.367
R283 B.n295 B.n294 163.367
R284 B.n296 B.n295 163.367
R285 B.n296 B.n9 163.367
R286 B.n300 B.n9 163.367
R287 B.n301 B.n300 163.367
R288 B.n302 B.n301 163.367
R289 B.n302 B.n7 163.367
R290 B.n306 B.n7 163.367
R291 B.n307 B.n306 163.367
R292 B.n308 B.n307 163.367
R293 B.n308 B.n5 163.367
R294 B.n312 B.n5 163.367
R295 B.n313 B.n312 163.367
R296 B.n314 B.n313 163.367
R297 B.n314 B.n3 163.367
R298 B.n318 B.n3 163.367
R299 B.n319 B.n318 163.367
R300 B.n86 B.n2 163.367
R301 B.n87 B.n86 163.367
R302 B.n87 B.n84 163.367
R303 B.n91 B.n84 163.367
R304 B.n92 B.n91 163.367
R305 B.n93 B.n92 163.367
R306 B.n93 B.n82 163.367
R307 B.n97 B.n82 163.367
R308 B.n98 B.n97 163.367
R309 B.n99 B.n98 163.367
R310 B.n99 B.n80 163.367
R311 B.n103 B.n80 163.367
R312 B.n104 B.n103 163.367
R313 B.n105 B.n104 163.367
R314 B.n105 B.n78 163.367
R315 B.n109 B.n78 163.367
R316 B.n110 B.n109 163.367
R317 B.n111 B.n110 163.367
R318 B.n111 B.n76 163.367
R319 B.n115 B.n76 163.367
R320 B.n116 B.n115 163.367
R321 B.n117 B.n116 163.367
R322 B.n134 B.n133 59.5399
R323 B.n152 B.n64 59.5399
R324 B.n255 B.n28 59.5399
R325 B.n22 B.n21 59.5399
R326 B.n133 B.n132 51.5884
R327 B.n64 B.n63 51.5884
R328 B.n28 B.n27 51.5884
R329 B.n21 B.n20 51.5884
R330 B.n286 B.n285 36.6834
R331 B.n238 B.n33 36.6834
R332 B.n166 B.n57 36.6834
R333 B.n119 B.n118 36.6834
R334 B B.n321 18.0485
R335 B.n287 B.n286 10.6151
R336 B.n287 B.n12 10.6151
R337 B.n291 B.n12 10.6151
R338 B.n292 B.n291 10.6151
R339 B.n293 B.n292 10.6151
R340 B.n293 B.n10 10.6151
R341 B.n297 B.n10 10.6151
R342 B.n298 B.n297 10.6151
R343 B.n299 B.n298 10.6151
R344 B.n299 B.n8 10.6151
R345 B.n303 B.n8 10.6151
R346 B.n304 B.n303 10.6151
R347 B.n305 B.n304 10.6151
R348 B.n305 B.n6 10.6151
R349 B.n309 B.n6 10.6151
R350 B.n310 B.n309 10.6151
R351 B.n311 B.n310 10.6151
R352 B.n311 B.n4 10.6151
R353 B.n315 B.n4 10.6151
R354 B.n316 B.n315 10.6151
R355 B.n317 B.n316 10.6151
R356 B.n317 B.n0 10.6151
R357 B.n285 B.n14 10.6151
R358 B.n281 B.n14 10.6151
R359 B.n281 B.n280 10.6151
R360 B.n280 B.n279 10.6151
R361 B.n279 B.n16 10.6151
R362 B.n275 B.n16 10.6151
R363 B.n275 B.n274 10.6151
R364 B.n274 B.n273 10.6151
R365 B.n273 B.n18 10.6151
R366 B.n269 B.n268 10.6151
R367 B.n268 B.n267 10.6151
R368 B.n267 B.n23 10.6151
R369 B.n263 B.n23 10.6151
R370 B.n263 B.n262 10.6151
R371 B.n262 B.n261 10.6151
R372 B.n261 B.n25 10.6151
R373 B.n257 B.n25 10.6151
R374 B.n257 B.n256 10.6151
R375 B.n254 B.n29 10.6151
R376 B.n250 B.n29 10.6151
R377 B.n250 B.n249 10.6151
R378 B.n249 B.n248 10.6151
R379 B.n248 B.n31 10.6151
R380 B.n244 B.n31 10.6151
R381 B.n244 B.n243 10.6151
R382 B.n243 B.n242 10.6151
R383 B.n242 B.n33 10.6151
R384 B.n238 B.n237 10.6151
R385 B.n237 B.n236 10.6151
R386 B.n236 B.n35 10.6151
R387 B.n232 B.n35 10.6151
R388 B.n232 B.n231 10.6151
R389 B.n231 B.n230 10.6151
R390 B.n230 B.n37 10.6151
R391 B.n226 B.n37 10.6151
R392 B.n226 B.n225 10.6151
R393 B.n225 B.n224 10.6151
R394 B.n224 B.n39 10.6151
R395 B.n220 B.n39 10.6151
R396 B.n220 B.n219 10.6151
R397 B.n219 B.n218 10.6151
R398 B.n218 B.n41 10.6151
R399 B.n214 B.n41 10.6151
R400 B.n214 B.n213 10.6151
R401 B.n213 B.n212 10.6151
R402 B.n212 B.n43 10.6151
R403 B.n208 B.n43 10.6151
R404 B.n208 B.n207 10.6151
R405 B.n207 B.n206 10.6151
R406 B.n206 B.n45 10.6151
R407 B.n202 B.n45 10.6151
R408 B.n202 B.n201 10.6151
R409 B.n201 B.n200 10.6151
R410 B.n200 B.n47 10.6151
R411 B.n196 B.n47 10.6151
R412 B.n196 B.n195 10.6151
R413 B.n195 B.n194 10.6151
R414 B.n194 B.n49 10.6151
R415 B.n190 B.n49 10.6151
R416 B.n190 B.n189 10.6151
R417 B.n189 B.n188 10.6151
R418 B.n188 B.n51 10.6151
R419 B.n184 B.n51 10.6151
R420 B.n184 B.n183 10.6151
R421 B.n183 B.n182 10.6151
R422 B.n182 B.n53 10.6151
R423 B.n178 B.n53 10.6151
R424 B.n178 B.n177 10.6151
R425 B.n177 B.n176 10.6151
R426 B.n176 B.n55 10.6151
R427 B.n172 B.n55 10.6151
R428 B.n172 B.n171 10.6151
R429 B.n171 B.n170 10.6151
R430 B.n170 B.n57 10.6151
R431 B.n85 B.n1 10.6151
R432 B.n88 B.n85 10.6151
R433 B.n89 B.n88 10.6151
R434 B.n90 B.n89 10.6151
R435 B.n90 B.n83 10.6151
R436 B.n94 B.n83 10.6151
R437 B.n95 B.n94 10.6151
R438 B.n96 B.n95 10.6151
R439 B.n96 B.n81 10.6151
R440 B.n100 B.n81 10.6151
R441 B.n101 B.n100 10.6151
R442 B.n102 B.n101 10.6151
R443 B.n102 B.n79 10.6151
R444 B.n106 B.n79 10.6151
R445 B.n107 B.n106 10.6151
R446 B.n108 B.n107 10.6151
R447 B.n108 B.n77 10.6151
R448 B.n112 B.n77 10.6151
R449 B.n113 B.n112 10.6151
R450 B.n114 B.n113 10.6151
R451 B.n114 B.n75 10.6151
R452 B.n118 B.n75 10.6151
R453 B.n120 B.n119 10.6151
R454 B.n120 B.n73 10.6151
R455 B.n124 B.n73 10.6151
R456 B.n125 B.n124 10.6151
R457 B.n126 B.n125 10.6151
R458 B.n126 B.n71 10.6151
R459 B.n130 B.n71 10.6151
R460 B.n131 B.n130 10.6151
R461 B.n135 B.n131 10.6151
R462 B.n139 B.n69 10.6151
R463 B.n140 B.n139 10.6151
R464 B.n141 B.n140 10.6151
R465 B.n141 B.n67 10.6151
R466 B.n145 B.n67 10.6151
R467 B.n146 B.n145 10.6151
R468 B.n147 B.n146 10.6151
R469 B.n147 B.n65 10.6151
R470 B.n151 B.n65 10.6151
R471 B.n154 B.n153 10.6151
R472 B.n154 B.n61 10.6151
R473 B.n158 B.n61 10.6151
R474 B.n159 B.n158 10.6151
R475 B.n160 B.n159 10.6151
R476 B.n160 B.n59 10.6151
R477 B.n164 B.n59 10.6151
R478 B.n165 B.n164 10.6151
R479 B.n166 B.n165 10.6151
R480 B.n22 B.n18 9.36635
R481 B.n255 B.n254 9.36635
R482 B.n135 B.n134 9.36635
R483 B.n153 B.n152 9.36635
R484 B.n321 B.n0 8.11757
R485 B.n321 B.n1 8.11757
R486 B.n269 B.n22 1.24928
R487 B.n256 B.n255 1.24928
R488 B.n134 B.n69 1.24928
R489 B.n152 B.n151 1.24928
R490 VN VN.t1 99.3252
R491 VN VN.t0 63.6775
R492 VTAIL.n1 VTAIL.t2 255.478
R493 VTAIL.n3 VTAIL.t3 255.478
R494 VTAIL.n0 VTAIL.t1 255.478
R495 VTAIL.n2 VTAIL.t0 255.478
R496 VTAIL.n1 VTAIL.n0 18.1341
R497 VTAIL.n3 VTAIL.n2 15.841
R498 VTAIL.n2 VTAIL.n1 1.61688
R499 VTAIL VTAIL.n0 1.10179
R500 VTAIL VTAIL.n3 0.515586
R501 VDD2.n0 VDD2.t1 301.584
R502 VDD2.n0 VDD2.t0 272.158
R503 VDD2 VDD2.n0 0.631965
R504 VP.n0 VP.t1 99.2287
R505 VP.n0 VP.t0 63.3412
R506 VP VP.n0 0.336784
R507 VDD1 VDD1.t1 302.683
R508 VDD1 VDD1.t0 272.788
C0 w_n2034_n1242# VTAIL 1.17682f
C1 B VDD2 0.86207f
C2 VDD1 VTAIL 2.16733f
C3 VDD2 VN 0.537578f
C4 w_n2034_n1242# VP 2.80536f
C5 VP VDD1 0.709646f
C6 B w_n2034_n1242# 5.56832f
C7 VP VTAIL 0.868498f
C8 w_n2034_n1242# VN 2.55339f
C9 B VDD1 0.833923f
C10 VDD1 VN 0.155238f
C11 B VTAIL 1.08819f
C12 VN VTAIL 0.854368f
C13 B VP 1.25225f
C14 VP VN 3.36953f
C15 B VN 0.829363f
C16 w_n2034_n1242# VDD2 1.02177f
C17 VDD1 VDD2 0.640957f
C18 VDD2 VTAIL 2.21856f
C19 VP VDD2 0.32903f
C20 w_n2034_n1242# VDD1 1.00005f
C21 VDD2 VSUBS 0.509233f
C22 VDD1 VSUBS 2.539893f
C23 VTAIL VSUBS 0.33132f
C24 VN VSUBS 5.38271f
C25 VP VSUBS 1.121862f
C26 B VSUBS 2.661599f
C27 w_n2034_n1242# VSUBS 32.4382f
C28 VDD1.t0 VSUBS 0.115115f
C29 VDD1.t1 VSUBS 0.195855f
C30 VP.t1 VSUBS 1.66219f
C31 VP.t0 VSUBS 0.8643f
C32 VP.n0 VSUBS 3.54662f
C33 VDD2.t1 VSUBS 0.19379f
C34 VDD2.t0 VSUBS 0.118118f
C35 VDD2.n0 VSUBS 1.78404f
C36 VTAIL.t1 VSUBS 0.135858f
C37 VTAIL.n0 VSUBS 1.01065f
C38 VTAIL.t2 VSUBS 0.135858f
C39 VTAIL.n1 VSUBS 1.04859f
C40 VTAIL.t0 VSUBS 0.135858f
C41 VTAIL.n2 VSUBS 0.879689f
C42 VTAIL.t3 VSUBS 0.135858f
C43 VTAIL.n3 VSUBS 0.79857f
C44 VN.t0 VSUBS 0.827165f
C45 VN.t1 VSUBS 1.59679f
C46 B.n0 VSUBS 0.009225f
C47 B.n1 VSUBS 0.009225f
C48 B.n2 VSUBS 0.013644f
C49 B.n3 VSUBS 0.010455f
C50 B.n4 VSUBS 0.010455f
C51 B.n5 VSUBS 0.010455f
C52 B.n6 VSUBS 0.010455f
C53 B.n7 VSUBS 0.010455f
C54 B.n8 VSUBS 0.010455f
C55 B.n9 VSUBS 0.010455f
C56 B.n10 VSUBS 0.010455f
C57 B.n11 VSUBS 0.010455f
C58 B.n12 VSUBS 0.010455f
C59 B.n13 VSUBS 0.025815f
C60 B.n14 VSUBS 0.010455f
C61 B.n15 VSUBS 0.010455f
C62 B.n16 VSUBS 0.010455f
C63 B.n17 VSUBS 0.010455f
C64 B.n18 VSUBS 0.00984f
C65 B.n19 VSUBS 0.010455f
C66 B.t10 VSUBS 0.041049f
C67 B.t11 VSUBS 0.051289f
C68 B.t9 VSUBS 0.237654f
C69 B.n20 VSUBS 0.09227f
C70 B.n21 VSUBS 0.074576f
C71 B.n22 VSUBS 0.024224f
C72 B.n23 VSUBS 0.010455f
C73 B.n24 VSUBS 0.010455f
C74 B.n25 VSUBS 0.010455f
C75 B.n26 VSUBS 0.010455f
C76 B.t4 VSUBS 0.041049f
C77 B.t5 VSUBS 0.051289f
C78 B.t3 VSUBS 0.237654f
C79 B.n27 VSUBS 0.09227f
C80 B.n28 VSUBS 0.074576f
C81 B.n29 VSUBS 0.010455f
C82 B.n30 VSUBS 0.010455f
C83 B.n31 VSUBS 0.010455f
C84 B.n32 VSUBS 0.010455f
C85 B.n33 VSUBS 0.027076f
C86 B.n34 VSUBS 0.010455f
C87 B.n35 VSUBS 0.010455f
C88 B.n36 VSUBS 0.010455f
C89 B.n37 VSUBS 0.010455f
C90 B.n38 VSUBS 0.010455f
C91 B.n39 VSUBS 0.010455f
C92 B.n40 VSUBS 0.010455f
C93 B.n41 VSUBS 0.010455f
C94 B.n42 VSUBS 0.010455f
C95 B.n43 VSUBS 0.010455f
C96 B.n44 VSUBS 0.010455f
C97 B.n45 VSUBS 0.010455f
C98 B.n46 VSUBS 0.010455f
C99 B.n47 VSUBS 0.010455f
C100 B.n48 VSUBS 0.010455f
C101 B.n49 VSUBS 0.010455f
C102 B.n50 VSUBS 0.010455f
C103 B.n51 VSUBS 0.010455f
C104 B.n52 VSUBS 0.010455f
C105 B.n53 VSUBS 0.010455f
C106 B.n54 VSUBS 0.010455f
C107 B.n55 VSUBS 0.010455f
C108 B.n56 VSUBS 0.010455f
C109 B.n57 VSUBS 0.026915f
C110 B.n58 VSUBS 0.010455f
C111 B.n59 VSUBS 0.010455f
C112 B.n60 VSUBS 0.010455f
C113 B.n61 VSUBS 0.010455f
C114 B.n62 VSUBS 0.010455f
C115 B.t8 VSUBS 0.041049f
C116 B.t7 VSUBS 0.051289f
C117 B.t6 VSUBS 0.237654f
C118 B.n63 VSUBS 0.09227f
C119 B.n64 VSUBS 0.074576f
C120 B.n65 VSUBS 0.010455f
C121 B.n66 VSUBS 0.010455f
C122 B.n67 VSUBS 0.010455f
C123 B.n68 VSUBS 0.010455f
C124 B.n69 VSUBS 0.005843f
C125 B.n70 VSUBS 0.010455f
C126 B.n71 VSUBS 0.010455f
C127 B.n72 VSUBS 0.010455f
C128 B.n73 VSUBS 0.010455f
C129 B.n74 VSUBS 0.027076f
C130 B.n75 VSUBS 0.010455f
C131 B.n76 VSUBS 0.010455f
C132 B.n77 VSUBS 0.010455f
C133 B.n78 VSUBS 0.010455f
C134 B.n79 VSUBS 0.010455f
C135 B.n80 VSUBS 0.010455f
C136 B.n81 VSUBS 0.010455f
C137 B.n82 VSUBS 0.010455f
C138 B.n83 VSUBS 0.010455f
C139 B.n84 VSUBS 0.010455f
C140 B.n85 VSUBS 0.010455f
C141 B.n86 VSUBS 0.010455f
C142 B.n87 VSUBS 0.010455f
C143 B.n88 VSUBS 0.010455f
C144 B.n89 VSUBS 0.010455f
C145 B.n90 VSUBS 0.010455f
C146 B.n91 VSUBS 0.010455f
C147 B.n92 VSUBS 0.010455f
C148 B.n93 VSUBS 0.010455f
C149 B.n94 VSUBS 0.010455f
C150 B.n95 VSUBS 0.010455f
C151 B.n96 VSUBS 0.010455f
C152 B.n97 VSUBS 0.010455f
C153 B.n98 VSUBS 0.010455f
C154 B.n99 VSUBS 0.010455f
C155 B.n100 VSUBS 0.010455f
C156 B.n101 VSUBS 0.010455f
C157 B.n102 VSUBS 0.010455f
C158 B.n103 VSUBS 0.010455f
C159 B.n104 VSUBS 0.010455f
C160 B.n105 VSUBS 0.010455f
C161 B.n106 VSUBS 0.010455f
C162 B.n107 VSUBS 0.010455f
C163 B.n108 VSUBS 0.010455f
C164 B.n109 VSUBS 0.010455f
C165 B.n110 VSUBS 0.010455f
C166 B.n111 VSUBS 0.010455f
C167 B.n112 VSUBS 0.010455f
C168 B.n113 VSUBS 0.010455f
C169 B.n114 VSUBS 0.010455f
C170 B.n115 VSUBS 0.010455f
C171 B.n116 VSUBS 0.010455f
C172 B.n117 VSUBS 0.025815f
C173 B.n118 VSUBS 0.025815f
C174 B.n119 VSUBS 0.027076f
C175 B.n120 VSUBS 0.010455f
C176 B.n121 VSUBS 0.010455f
C177 B.n122 VSUBS 0.010455f
C178 B.n123 VSUBS 0.010455f
C179 B.n124 VSUBS 0.010455f
C180 B.n125 VSUBS 0.010455f
C181 B.n126 VSUBS 0.010455f
C182 B.n127 VSUBS 0.010455f
C183 B.n128 VSUBS 0.010455f
C184 B.n129 VSUBS 0.010455f
C185 B.n130 VSUBS 0.010455f
C186 B.n131 VSUBS 0.010455f
C187 B.t2 VSUBS 0.041049f
C188 B.t1 VSUBS 0.051289f
C189 B.t0 VSUBS 0.237654f
C190 B.n132 VSUBS 0.09227f
C191 B.n133 VSUBS 0.074576f
C192 B.n134 VSUBS 0.024224f
C193 B.n135 VSUBS 0.00984f
C194 B.n136 VSUBS 0.010455f
C195 B.n137 VSUBS 0.010455f
C196 B.n138 VSUBS 0.010455f
C197 B.n139 VSUBS 0.010455f
C198 B.n140 VSUBS 0.010455f
C199 B.n141 VSUBS 0.010455f
C200 B.n142 VSUBS 0.010455f
C201 B.n143 VSUBS 0.010455f
C202 B.n144 VSUBS 0.010455f
C203 B.n145 VSUBS 0.010455f
C204 B.n146 VSUBS 0.010455f
C205 B.n147 VSUBS 0.010455f
C206 B.n148 VSUBS 0.010455f
C207 B.n149 VSUBS 0.010455f
C208 B.n150 VSUBS 0.010455f
C209 B.n151 VSUBS 0.005843f
C210 B.n152 VSUBS 0.024224f
C211 B.n153 VSUBS 0.00984f
C212 B.n154 VSUBS 0.010455f
C213 B.n155 VSUBS 0.010455f
C214 B.n156 VSUBS 0.010455f
C215 B.n157 VSUBS 0.010455f
C216 B.n158 VSUBS 0.010455f
C217 B.n159 VSUBS 0.010455f
C218 B.n160 VSUBS 0.010455f
C219 B.n161 VSUBS 0.010455f
C220 B.n162 VSUBS 0.010455f
C221 B.n163 VSUBS 0.010455f
C222 B.n164 VSUBS 0.010455f
C223 B.n165 VSUBS 0.010455f
C224 B.n166 VSUBS 0.025976f
C225 B.n167 VSUBS 0.027076f
C226 B.n168 VSUBS 0.025815f
C227 B.n169 VSUBS 0.010455f
C228 B.n170 VSUBS 0.010455f
C229 B.n171 VSUBS 0.010455f
C230 B.n172 VSUBS 0.010455f
C231 B.n173 VSUBS 0.010455f
C232 B.n174 VSUBS 0.010455f
C233 B.n175 VSUBS 0.010455f
C234 B.n176 VSUBS 0.010455f
C235 B.n177 VSUBS 0.010455f
C236 B.n178 VSUBS 0.010455f
C237 B.n179 VSUBS 0.010455f
C238 B.n180 VSUBS 0.010455f
C239 B.n181 VSUBS 0.010455f
C240 B.n182 VSUBS 0.010455f
C241 B.n183 VSUBS 0.010455f
C242 B.n184 VSUBS 0.010455f
C243 B.n185 VSUBS 0.010455f
C244 B.n186 VSUBS 0.010455f
C245 B.n187 VSUBS 0.010455f
C246 B.n188 VSUBS 0.010455f
C247 B.n189 VSUBS 0.010455f
C248 B.n190 VSUBS 0.010455f
C249 B.n191 VSUBS 0.010455f
C250 B.n192 VSUBS 0.010455f
C251 B.n193 VSUBS 0.010455f
C252 B.n194 VSUBS 0.010455f
C253 B.n195 VSUBS 0.010455f
C254 B.n196 VSUBS 0.010455f
C255 B.n197 VSUBS 0.010455f
C256 B.n198 VSUBS 0.010455f
C257 B.n199 VSUBS 0.010455f
C258 B.n200 VSUBS 0.010455f
C259 B.n201 VSUBS 0.010455f
C260 B.n202 VSUBS 0.010455f
C261 B.n203 VSUBS 0.010455f
C262 B.n204 VSUBS 0.010455f
C263 B.n205 VSUBS 0.010455f
C264 B.n206 VSUBS 0.010455f
C265 B.n207 VSUBS 0.010455f
C266 B.n208 VSUBS 0.010455f
C267 B.n209 VSUBS 0.010455f
C268 B.n210 VSUBS 0.010455f
C269 B.n211 VSUBS 0.010455f
C270 B.n212 VSUBS 0.010455f
C271 B.n213 VSUBS 0.010455f
C272 B.n214 VSUBS 0.010455f
C273 B.n215 VSUBS 0.010455f
C274 B.n216 VSUBS 0.010455f
C275 B.n217 VSUBS 0.010455f
C276 B.n218 VSUBS 0.010455f
C277 B.n219 VSUBS 0.010455f
C278 B.n220 VSUBS 0.010455f
C279 B.n221 VSUBS 0.010455f
C280 B.n222 VSUBS 0.010455f
C281 B.n223 VSUBS 0.010455f
C282 B.n224 VSUBS 0.010455f
C283 B.n225 VSUBS 0.010455f
C284 B.n226 VSUBS 0.010455f
C285 B.n227 VSUBS 0.010455f
C286 B.n228 VSUBS 0.010455f
C287 B.n229 VSUBS 0.010455f
C288 B.n230 VSUBS 0.010455f
C289 B.n231 VSUBS 0.010455f
C290 B.n232 VSUBS 0.010455f
C291 B.n233 VSUBS 0.010455f
C292 B.n234 VSUBS 0.010455f
C293 B.n235 VSUBS 0.010455f
C294 B.n236 VSUBS 0.010455f
C295 B.n237 VSUBS 0.010455f
C296 B.n238 VSUBS 0.025815f
C297 B.n239 VSUBS 0.025815f
C298 B.n240 VSUBS 0.027076f
C299 B.n241 VSUBS 0.010455f
C300 B.n242 VSUBS 0.010455f
C301 B.n243 VSUBS 0.010455f
C302 B.n244 VSUBS 0.010455f
C303 B.n245 VSUBS 0.010455f
C304 B.n246 VSUBS 0.010455f
C305 B.n247 VSUBS 0.010455f
C306 B.n248 VSUBS 0.010455f
C307 B.n249 VSUBS 0.010455f
C308 B.n250 VSUBS 0.010455f
C309 B.n251 VSUBS 0.010455f
C310 B.n252 VSUBS 0.010455f
C311 B.n253 VSUBS 0.010455f
C312 B.n254 VSUBS 0.00984f
C313 B.n255 VSUBS 0.024224f
C314 B.n256 VSUBS 0.005843f
C315 B.n257 VSUBS 0.010455f
C316 B.n258 VSUBS 0.010455f
C317 B.n259 VSUBS 0.010455f
C318 B.n260 VSUBS 0.010455f
C319 B.n261 VSUBS 0.010455f
C320 B.n262 VSUBS 0.010455f
C321 B.n263 VSUBS 0.010455f
C322 B.n264 VSUBS 0.010455f
C323 B.n265 VSUBS 0.010455f
C324 B.n266 VSUBS 0.010455f
C325 B.n267 VSUBS 0.010455f
C326 B.n268 VSUBS 0.010455f
C327 B.n269 VSUBS 0.005843f
C328 B.n270 VSUBS 0.010455f
C329 B.n271 VSUBS 0.010455f
C330 B.n272 VSUBS 0.010455f
C331 B.n273 VSUBS 0.010455f
C332 B.n274 VSUBS 0.010455f
C333 B.n275 VSUBS 0.010455f
C334 B.n276 VSUBS 0.010455f
C335 B.n277 VSUBS 0.010455f
C336 B.n278 VSUBS 0.010455f
C337 B.n279 VSUBS 0.010455f
C338 B.n280 VSUBS 0.010455f
C339 B.n281 VSUBS 0.010455f
C340 B.n282 VSUBS 0.010455f
C341 B.n283 VSUBS 0.010455f
C342 B.n284 VSUBS 0.027076f
C343 B.n285 VSUBS 0.027076f
C344 B.n286 VSUBS 0.025815f
C345 B.n287 VSUBS 0.010455f
C346 B.n288 VSUBS 0.010455f
C347 B.n289 VSUBS 0.010455f
C348 B.n290 VSUBS 0.010455f
C349 B.n291 VSUBS 0.010455f
C350 B.n292 VSUBS 0.010455f
C351 B.n293 VSUBS 0.010455f
C352 B.n294 VSUBS 0.010455f
C353 B.n295 VSUBS 0.010455f
C354 B.n296 VSUBS 0.010455f
C355 B.n297 VSUBS 0.010455f
C356 B.n298 VSUBS 0.010455f
C357 B.n299 VSUBS 0.010455f
C358 B.n300 VSUBS 0.010455f
C359 B.n301 VSUBS 0.010455f
C360 B.n302 VSUBS 0.010455f
C361 B.n303 VSUBS 0.010455f
C362 B.n304 VSUBS 0.010455f
C363 B.n305 VSUBS 0.010455f
C364 B.n306 VSUBS 0.010455f
C365 B.n307 VSUBS 0.010455f
C366 B.n308 VSUBS 0.010455f
C367 B.n309 VSUBS 0.010455f
C368 B.n310 VSUBS 0.010455f
C369 B.n311 VSUBS 0.010455f
C370 B.n312 VSUBS 0.010455f
C371 B.n313 VSUBS 0.010455f
C372 B.n314 VSUBS 0.010455f
C373 B.n315 VSUBS 0.010455f
C374 B.n316 VSUBS 0.010455f
C375 B.n317 VSUBS 0.010455f
C376 B.n318 VSUBS 0.010455f
C377 B.n319 VSUBS 0.013644f
C378 B.n320 VSUBS 0.014534f
C379 B.n321 VSUBS 0.028902f
.ends

