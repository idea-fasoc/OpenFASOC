* NGSPICE file created from diff_pair_sample_1089.ext - technology: sky130A

.subckt diff_pair_sample_1089 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=7.0356 pd=36.86 as=0 ps=0 w=18.04 l=0.56
X1 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=7.0356 pd=36.86 as=0 ps=0 w=18.04 l=0.56
X2 VDD1.t3 VP.t0 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.9766 pd=18.37 as=7.0356 ps=36.86 w=18.04 l=0.56
X3 VTAIL.t0 VN.t0 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=7.0356 pd=36.86 as=2.9766 ps=18.37 w=18.04 l=0.56
X4 VDD2.t2 VN.t1 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9766 pd=18.37 as=7.0356 ps=36.86 w=18.04 l=0.56
X5 VTAIL.t6 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=7.0356 pd=36.86 as=2.9766 ps=18.37 w=18.04 l=0.56
X6 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.0356 pd=36.86 as=0 ps=0 w=18.04 l=0.56
X7 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.0356 pd=36.86 as=0 ps=0 w=18.04 l=0.56
X8 VTAIL.t2 VN.t2 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=7.0356 pd=36.86 as=2.9766 ps=18.37 w=18.04 l=0.56
X9 VDD2.t0 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.9766 pd=18.37 as=7.0356 ps=36.86 w=18.04 l=0.56
X10 VDD1.t1 VP.t2 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9766 pd=18.37 as=7.0356 ps=36.86 w=18.04 l=0.56
X11 VTAIL.t4 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=7.0356 pd=36.86 as=2.9766 ps=18.37 w=18.04 l=0.56
R0 B.n415 B.t12 981.481
R1 B.n424 B.t8 981.481
R2 B.n100 B.t15 981.481
R3 B.n98 B.t4 981.481
R4 B.n780 B.n779 585
R5 B.n354 B.n97 585
R6 B.n353 B.n352 585
R7 B.n351 B.n350 585
R8 B.n349 B.n348 585
R9 B.n347 B.n346 585
R10 B.n345 B.n344 585
R11 B.n343 B.n342 585
R12 B.n341 B.n340 585
R13 B.n339 B.n338 585
R14 B.n337 B.n336 585
R15 B.n335 B.n334 585
R16 B.n333 B.n332 585
R17 B.n331 B.n330 585
R18 B.n329 B.n328 585
R19 B.n327 B.n326 585
R20 B.n325 B.n324 585
R21 B.n323 B.n322 585
R22 B.n321 B.n320 585
R23 B.n319 B.n318 585
R24 B.n317 B.n316 585
R25 B.n315 B.n314 585
R26 B.n313 B.n312 585
R27 B.n311 B.n310 585
R28 B.n309 B.n308 585
R29 B.n307 B.n306 585
R30 B.n305 B.n304 585
R31 B.n303 B.n302 585
R32 B.n301 B.n300 585
R33 B.n299 B.n298 585
R34 B.n297 B.n296 585
R35 B.n295 B.n294 585
R36 B.n293 B.n292 585
R37 B.n291 B.n290 585
R38 B.n289 B.n288 585
R39 B.n287 B.n286 585
R40 B.n285 B.n284 585
R41 B.n283 B.n282 585
R42 B.n281 B.n280 585
R43 B.n279 B.n278 585
R44 B.n277 B.n276 585
R45 B.n275 B.n274 585
R46 B.n273 B.n272 585
R47 B.n271 B.n270 585
R48 B.n269 B.n268 585
R49 B.n267 B.n266 585
R50 B.n265 B.n264 585
R51 B.n263 B.n262 585
R52 B.n261 B.n260 585
R53 B.n259 B.n258 585
R54 B.n257 B.n256 585
R55 B.n255 B.n254 585
R56 B.n253 B.n252 585
R57 B.n251 B.n250 585
R58 B.n249 B.n248 585
R59 B.n247 B.n246 585
R60 B.n245 B.n244 585
R61 B.n243 B.n242 585
R62 B.n241 B.n240 585
R63 B.n238 B.n237 585
R64 B.n236 B.n235 585
R65 B.n234 B.n233 585
R66 B.n232 B.n231 585
R67 B.n230 B.n229 585
R68 B.n228 B.n227 585
R69 B.n226 B.n225 585
R70 B.n224 B.n223 585
R71 B.n222 B.n221 585
R72 B.n220 B.n219 585
R73 B.n217 B.n216 585
R74 B.n215 B.n214 585
R75 B.n213 B.n212 585
R76 B.n211 B.n210 585
R77 B.n209 B.n208 585
R78 B.n207 B.n206 585
R79 B.n205 B.n204 585
R80 B.n203 B.n202 585
R81 B.n201 B.n200 585
R82 B.n199 B.n198 585
R83 B.n197 B.n196 585
R84 B.n195 B.n194 585
R85 B.n193 B.n192 585
R86 B.n191 B.n190 585
R87 B.n189 B.n188 585
R88 B.n187 B.n186 585
R89 B.n185 B.n184 585
R90 B.n183 B.n182 585
R91 B.n181 B.n180 585
R92 B.n179 B.n178 585
R93 B.n177 B.n176 585
R94 B.n175 B.n174 585
R95 B.n173 B.n172 585
R96 B.n171 B.n170 585
R97 B.n169 B.n168 585
R98 B.n167 B.n166 585
R99 B.n165 B.n164 585
R100 B.n163 B.n162 585
R101 B.n161 B.n160 585
R102 B.n159 B.n158 585
R103 B.n157 B.n156 585
R104 B.n155 B.n154 585
R105 B.n153 B.n152 585
R106 B.n151 B.n150 585
R107 B.n149 B.n148 585
R108 B.n147 B.n146 585
R109 B.n145 B.n144 585
R110 B.n143 B.n142 585
R111 B.n141 B.n140 585
R112 B.n139 B.n138 585
R113 B.n137 B.n136 585
R114 B.n135 B.n134 585
R115 B.n133 B.n132 585
R116 B.n131 B.n130 585
R117 B.n129 B.n128 585
R118 B.n127 B.n126 585
R119 B.n125 B.n124 585
R120 B.n123 B.n122 585
R121 B.n121 B.n120 585
R122 B.n119 B.n118 585
R123 B.n117 B.n116 585
R124 B.n115 B.n114 585
R125 B.n113 B.n112 585
R126 B.n111 B.n110 585
R127 B.n109 B.n108 585
R128 B.n107 B.n106 585
R129 B.n105 B.n104 585
R130 B.n103 B.n102 585
R131 B.n32 B.n31 585
R132 B.n778 B.n33 585
R133 B.n783 B.n33 585
R134 B.n777 B.n776 585
R135 B.n776 B.n29 585
R136 B.n775 B.n28 585
R137 B.n789 B.n28 585
R138 B.n774 B.n27 585
R139 B.n790 B.n27 585
R140 B.n773 B.n26 585
R141 B.n791 B.n26 585
R142 B.n772 B.n771 585
R143 B.n771 B.n22 585
R144 B.n770 B.n21 585
R145 B.n797 B.n21 585
R146 B.n769 B.n20 585
R147 B.n798 B.n20 585
R148 B.n768 B.n19 585
R149 B.n799 B.n19 585
R150 B.n767 B.n766 585
R151 B.n766 B.n15 585
R152 B.n765 B.n14 585
R153 B.n805 B.n14 585
R154 B.n764 B.n13 585
R155 B.n806 B.n13 585
R156 B.n763 B.n12 585
R157 B.n807 B.n12 585
R158 B.n762 B.n761 585
R159 B.n761 B.n11 585
R160 B.n760 B.n7 585
R161 B.n813 B.n7 585
R162 B.n759 B.n6 585
R163 B.n814 B.n6 585
R164 B.n758 B.n5 585
R165 B.n815 B.n5 585
R166 B.n757 B.n756 585
R167 B.n756 B.n4 585
R168 B.n755 B.n355 585
R169 B.n755 B.n754 585
R170 B.n744 B.n356 585
R171 B.n747 B.n356 585
R172 B.n746 B.n745 585
R173 B.n748 B.n746 585
R174 B.n743 B.n361 585
R175 B.n361 B.n360 585
R176 B.n742 B.n741 585
R177 B.n741 B.n740 585
R178 B.n363 B.n362 585
R179 B.n364 B.n363 585
R180 B.n733 B.n732 585
R181 B.n734 B.n733 585
R182 B.n731 B.n369 585
R183 B.n369 B.n368 585
R184 B.n730 B.n729 585
R185 B.n729 B.n728 585
R186 B.n371 B.n370 585
R187 B.n372 B.n371 585
R188 B.n721 B.n720 585
R189 B.n722 B.n721 585
R190 B.n719 B.n377 585
R191 B.n377 B.n376 585
R192 B.n718 B.n717 585
R193 B.n717 B.n716 585
R194 B.n379 B.n378 585
R195 B.n380 B.n379 585
R196 B.n709 B.n708 585
R197 B.n710 B.n709 585
R198 B.n383 B.n382 585
R199 B.n456 B.n455 585
R200 B.n457 B.n453 585
R201 B.n453 B.n384 585
R202 B.n459 B.n458 585
R203 B.n461 B.n452 585
R204 B.n464 B.n463 585
R205 B.n465 B.n451 585
R206 B.n467 B.n466 585
R207 B.n469 B.n450 585
R208 B.n472 B.n471 585
R209 B.n473 B.n449 585
R210 B.n475 B.n474 585
R211 B.n477 B.n448 585
R212 B.n480 B.n479 585
R213 B.n481 B.n447 585
R214 B.n483 B.n482 585
R215 B.n485 B.n446 585
R216 B.n488 B.n487 585
R217 B.n489 B.n445 585
R218 B.n491 B.n490 585
R219 B.n493 B.n444 585
R220 B.n496 B.n495 585
R221 B.n497 B.n443 585
R222 B.n499 B.n498 585
R223 B.n501 B.n442 585
R224 B.n504 B.n503 585
R225 B.n505 B.n441 585
R226 B.n507 B.n506 585
R227 B.n509 B.n440 585
R228 B.n512 B.n511 585
R229 B.n513 B.n439 585
R230 B.n515 B.n514 585
R231 B.n517 B.n438 585
R232 B.n520 B.n519 585
R233 B.n521 B.n437 585
R234 B.n523 B.n522 585
R235 B.n525 B.n436 585
R236 B.n528 B.n527 585
R237 B.n529 B.n435 585
R238 B.n531 B.n530 585
R239 B.n533 B.n434 585
R240 B.n536 B.n535 585
R241 B.n537 B.n433 585
R242 B.n539 B.n538 585
R243 B.n541 B.n432 585
R244 B.n544 B.n543 585
R245 B.n545 B.n431 585
R246 B.n547 B.n546 585
R247 B.n549 B.n430 585
R248 B.n552 B.n551 585
R249 B.n553 B.n429 585
R250 B.n555 B.n554 585
R251 B.n557 B.n428 585
R252 B.n560 B.n559 585
R253 B.n561 B.n427 585
R254 B.n563 B.n562 585
R255 B.n565 B.n426 585
R256 B.n568 B.n567 585
R257 B.n569 B.n423 585
R258 B.n572 B.n571 585
R259 B.n574 B.n422 585
R260 B.n577 B.n576 585
R261 B.n578 B.n421 585
R262 B.n580 B.n579 585
R263 B.n582 B.n420 585
R264 B.n585 B.n584 585
R265 B.n586 B.n419 585
R266 B.n588 B.n587 585
R267 B.n590 B.n418 585
R268 B.n593 B.n592 585
R269 B.n594 B.n414 585
R270 B.n596 B.n595 585
R271 B.n598 B.n413 585
R272 B.n601 B.n600 585
R273 B.n602 B.n412 585
R274 B.n604 B.n603 585
R275 B.n606 B.n411 585
R276 B.n609 B.n608 585
R277 B.n610 B.n410 585
R278 B.n612 B.n611 585
R279 B.n614 B.n409 585
R280 B.n617 B.n616 585
R281 B.n618 B.n408 585
R282 B.n620 B.n619 585
R283 B.n622 B.n407 585
R284 B.n625 B.n624 585
R285 B.n626 B.n406 585
R286 B.n628 B.n627 585
R287 B.n630 B.n405 585
R288 B.n633 B.n632 585
R289 B.n634 B.n404 585
R290 B.n636 B.n635 585
R291 B.n638 B.n403 585
R292 B.n641 B.n640 585
R293 B.n642 B.n402 585
R294 B.n644 B.n643 585
R295 B.n646 B.n401 585
R296 B.n649 B.n648 585
R297 B.n650 B.n400 585
R298 B.n652 B.n651 585
R299 B.n654 B.n399 585
R300 B.n657 B.n656 585
R301 B.n658 B.n398 585
R302 B.n660 B.n659 585
R303 B.n662 B.n397 585
R304 B.n665 B.n664 585
R305 B.n666 B.n396 585
R306 B.n668 B.n667 585
R307 B.n670 B.n395 585
R308 B.n673 B.n672 585
R309 B.n674 B.n394 585
R310 B.n676 B.n675 585
R311 B.n678 B.n393 585
R312 B.n681 B.n680 585
R313 B.n682 B.n392 585
R314 B.n684 B.n683 585
R315 B.n686 B.n391 585
R316 B.n689 B.n688 585
R317 B.n690 B.n390 585
R318 B.n692 B.n691 585
R319 B.n694 B.n389 585
R320 B.n697 B.n696 585
R321 B.n698 B.n388 585
R322 B.n700 B.n699 585
R323 B.n702 B.n387 585
R324 B.n703 B.n386 585
R325 B.n706 B.n705 585
R326 B.n707 B.n385 585
R327 B.n385 B.n384 585
R328 B.n712 B.n711 585
R329 B.n711 B.n710 585
R330 B.n713 B.n381 585
R331 B.n381 B.n380 585
R332 B.n715 B.n714 585
R333 B.n716 B.n715 585
R334 B.n375 B.n374 585
R335 B.n376 B.n375 585
R336 B.n724 B.n723 585
R337 B.n723 B.n722 585
R338 B.n725 B.n373 585
R339 B.n373 B.n372 585
R340 B.n727 B.n726 585
R341 B.n728 B.n727 585
R342 B.n367 B.n366 585
R343 B.n368 B.n367 585
R344 B.n736 B.n735 585
R345 B.n735 B.n734 585
R346 B.n737 B.n365 585
R347 B.n365 B.n364 585
R348 B.n739 B.n738 585
R349 B.n740 B.n739 585
R350 B.n359 B.n358 585
R351 B.n360 B.n359 585
R352 B.n750 B.n749 585
R353 B.n749 B.n748 585
R354 B.n751 B.n357 585
R355 B.n747 B.n357 585
R356 B.n753 B.n752 585
R357 B.n754 B.n753 585
R358 B.n2 B.n0 585
R359 B.n4 B.n2 585
R360 B.n3 B.n1 585
R361 B.n814 B.n3 585
R362 B.n812 B.n811 585
R363 B.n813 B.n812 585
R364 B.n810 B.n8 585
R365 B.n11 B.n8 585
R366 B.n809 B.n808 585
R367 B.n808 B.n807 585
R368 B.n10 B.n9 585
R369 B.n806 B.n10 585
R370 B.n804 B.n803 585
R371 B.n805 B.n804 585
R372 B.n802 B.n16 585
R373 B.n16 B.n15 585
R374 B.n801 B.n800 585
R375 B.n800 B.n799 585
R376 B.n18 B.n17 585
R377 B.n798 B.n18 585
R378 B.n796 B.n795 585
R379 B.n797 B.n796 585
R380 B.n794 B.n23 585
R381 B.n23 B.n22 585
R382 B.n793 B.n792 585
R383 B.n792 B.n791 585
R384 B.n25 B.n24 585
R385 B.n790 B.n25 585
R386 B.n788 B.n787 585
R387 B.n789 B.n788 585
R388 B.n786 B.n30 585
R389 B.n30 B.n29 585
R390 B.n785 B.n784 585
R391 B.n784 B.n783 585
R392 B.n817 B.n816 585
R393 B.n816 B.n815 585
R394 B.n711 B.n383 521.33
R395 B.n784 B.n32 521.33
R396 B.n709 B.n385 521.33
R397 B.n780 B.n33 521.33
R398 B.n415 B.t14 403.128
R399 B.n98 B.t6 403.128
R400 B.n424 B.t11 403.128
R401 B.n100 B.t16 403.128
R402 B.n416 B.t13 385.868
R403 B.n99 B.t7 385.868
R404 B.n425 B.t10 385.868
R405 B.n101 B.t17 385.868
R406 B.n782 B.n781 256.663
R407 B.n782 B.n96 256.663
R408 B.n782 B.n95 256.663
R409 B.n782 B.n94 256.663
R410 B.n782 B.n93 256.663
R411 B.n782 B.n92 256.663
R412 B.n782 B.n91 256.663
R413 B.n782 B.n90 256.663
R414 B.n782 B.n89 256.663
R415 B.n782 B.n88 256.663
R416 B.n782 B.n87 256.663
R417 B.n782 B.n86 256.663
R418 B.n782 B.n85 256.663
R419 B.n782 B.n84 256.663
R420 B.n782 B.n83 256.663
R421 B.n782 B.n82 256.663
R422 B.n782 B.n81 256.663
R423 B.n782 B.n80 256.663
R424 B.n782 B.n79 256.663
R425 B.n782 B.n78 256.663
R426 B.n782 B.n77 256.663
R427 B.n782 B.n76 256.663
R428 B.n782 B.n75 256.663
R429 B.n782 B.n74 256.663
R430 B.n782 B.n73 256.663
R431 B.n782 B.n72 256.663
R432 B.n782 B.n71 256.663
R433 B.n782 B.n70 256.663
R434 B.n782 B.n69 256.663
R435 B.n782 B.n68 256.663
R436 B.n782 B.n67 256.663
R437 B.n782 B.n66 256.663
R438 B.n782 B.n65 256.663
R439 B.n782 B.n64 256.663
R440 B.n782 B.n63 256.663
R441 B.n782 B.n62 256.663
R442 B.n782 B.n61 256.663
R443 B.n782 B.n60 256.663
R444 B.n782 B.n59 256.663
R445 B.n782 B.n58 256.663
R446 B.n782 B.n57 256.663
R447 B.n782 B.n56 256.663
R448 B.n782 B.n55 256.663
R449 B.n782 B.n54 256.663
R450 B.n782 B.n53 256.663
R451 B.n782 B.n52 256.663
R452 B.n782 B.n51 256.663
R453 B.n782 B.n50 256.663
R454 B.n782 B.n49 256.663
R455 B.n782 B.n48 256.663
R456 B.n782 B.n47 256.663
R457 B.n782 B.n46 256.663
R458 B.n782 B.n45 256.663
R459 B.n782 B.n44 256.663
R460 B.n782 B.n43 256.663
R461 B.n782 B.n42 256.663
R462 B.n782 B.n41 256.663
R463 B.n782 B.n40 256.663
R464 B.n782 B.n39 256.663
R465 B.n782 B.n38 256.663
R466 B.n782 B.n37 256.663
R467 B.n782 B.n36 256.663
R468 B.n782 B.n35 256.663
R469 B.n782 B.n34 256.663
R470 B.n454 B.n384 256.663
R471 B.n460 B.n384 256.663
R472 B.n462 B.n384 256.663
R473 B.n468 B.n384 256.663
R474 B.n470 B.n384 256.663
R475 B.n476 B.n384 256.663
R476 B.n478 B.n384 256.663
R477 B.n484 B.n384 256.663
R478 B.n486 B.n384 256.663
R479 B.n492 B.n384 256.663
R480 B.n494 B.n384 256.663
R481 B.n500 B.n384 256.663
R482 B.n502 B.n384 256.663
R483 B.n508 B.n384 256.663
R484 B.n510 B.n384 256.663
R485 B.n516 B.n384 256.663
R486 B.n518 B.n384 256.663
R487 B.n524 B.n384 256.663
R488 B.n526 B.n384 256.663
R489 B.n532 B.n384 256.663
R490 B.n534 B.n384 256.663
R491 B.n540 B.n384 256.663
R492 B.n542 B.n384 256.663
R493 B.n548 B.n384 256.663
R494 B.n550 B.n384 256.663
R495 B.n556 B.n384 256.663
R496 B.n558 B.n384 256.663
R497 B.n564 B.n384 256.663
R498 B.n566 B.n384 256.663
R499 B.n573 B.n384 256.663
R500 B.n575 B.n384 256.663
R501 B.n581 B.n384 256.663
R502 B.n583 B.n384 256.663
R503 B.n589 B.n384 256.663
R504 B.n591 B.n384 256.663
R505 B.n597 B.n384 256.663
R506 B.n599 B.n384 256.663
R507 B.n605 B.n384 256.663
R508 B.n607 B.n384 256.663
R509 B.n613 B.n384 256.663
R510 B.n615 B.n384 256.663
R511 B.n621 B.n384 256.663
R512 B.n623 B.n384 256.663
R513 B.n629 B.n384 256.663
R514 B.n631 B.n384 256.663
R515 B.n637 B.n384 256.663
R516 B.n639 B.n384 256.663
R517 B.n645 B.n384 256.663
R518 B.n647 B.n384 256.663
R519 B.n653 B.n384 256.663
R520 B.n655 B.n384 256.663
R521 B.n661 B.n384 256.663
R522 B.n663 B.n384 256.663
R523 B.n669 B.n384 256.663
R524 B.n671 B.n384 256.663
R525 B.n677 B.n384 256.663
R526 B.n679 B.n384 256.663
R527 B.n685 B.n384 256.663
R528 B.n687 B.n384 256.663
R529 B.n693 B.n384 256.663
R530 B.n695 B.n384 256.663
R531 B.n701 B.n384 256.663
R532 B.n704 B.n384 256.663
R533 B.n711 B.n381 163.367
R534 B.n715 B.n381 163.367
R535 B.n715 B.n375 163.367
R536 B.n723 B.n375 163.367
R537 B.n723 B.n373 163.367
R538 B.n727 B.n373 163.367
R539 B.n727 B.n367 163.367
R540 B.n735 B.n367 163.367
R541 B.n735 B.n365 163.367
R542 B.n739 B.n365 163.367
R543 B.n739 B.n359 163.367
R544 B.n749 B.n359 163.367
R545 B.n749 B.n357 163.367
R546 B.n753 B.n357 163.367
R547 B.n753 B.n2 163.367
R548 B.n816 B.n2 163.367
R549 B.n816 B.n3 163.367
R550 B.n812 B.n3 163.367
R551 B.n812 B.n8 163.367
R552 B.n808 B.n8 163.367
R553 B.n808 B.n10 163.367
R554 B.n804 B.n10 163.367
R555 B.n804 B.n16 163.367
R556 B.n800 B.n16 163.367
R557 B.n800 B.n18 163.367
R558 B.n796 B.n18 163.367
R559 B.n796 B.n23 163.367
R560 B.n792 B.n23 163.367
R561 B.n792 B.n25 163.367
R562 B.n788 B.n25 163.367
R563 B.n788 B.n30 163.367
R564 B.n784 B.n30 163.367
R565 B.n455 B.n453 163.367
R566 B.n459 B.n453 163.367
R567 B.n463 B.n461 163.367
R568 B.n467 B.n451 163.367
R569 B.n471 B.n469 163.367
R570 B.n475 B.n449 163.367
R571 B.n479 B.n477 163.367
R572 B.n483 B.n447 163.367
R573 B.n487 B.n485 163.367
R574 B.n491 B.n445 163.367
R575 B.n495 B.n493 163.367
R576 B.n499 B.n443 163.367
R577 B.n503 B.n501 163.367
R578 B.n507 B.n441 163.367
R579 B.n511 B.n509 163.367
R580 B.n515 B.n439 163.367
R581 B.n519 B.n517 163.367
R582 B.n523 B.n437 163.367
R583 B.n527 B.n525 163.367
R584 B.n531 B.n435 163.367
R585 B.n535 B.n533 163.367
R586 B.n539 B.n433 163.367
R587 B.n543 B.n541 163.367
R588 B.n547 B.n431 163.367
R589 B.n551 B.n549 163.367
R590 B.n555 B.n429 163.367
R591 B.n559 B.n557 163.367
R592 B.n563 B.n427 163.367
R593 B.n567 B.n565 163.367
R594 B.n572 B.n423 163.367
R595 B.n576 B.n574 163.367
R596 B.n580 B.n421 163.367
R597 B.n584 B.n582 163.367
R598 B.n588 B.n419 163.367
R599 B.n592 B.n590 163.367
R600 B.n596 B.n414 163.367
R601 B.n600 B.n598 163.367
R602 B.n604 B.n412 163.367
R603 B.n608 B.n606 163.367
R604 B.n612 B.n410 163.367
R605 B.n616 B.n614 163.367
R606 B.n620 B.n408 163.367
R607 B.n624 B.n622 163.367
R608 B.n628 B.n406 163.367
R609 B.n632 B.n630 163.367
R610 B.n636 B.n404 163.367
R611 B.n640 B.n638 163.367
R612 B.n644 B.n402 163.367
R613 B.n648 B.n646 163.367
R614 B.n652 B.n400 163.367
R615 B.n656 B.n654 163.367
R616 B.n660 B.n398 163.367
R617 B.n664 B.n662 163.367
R618 B.n668 B.n396 163.367
R619 B.n672 B.n670 163.367
R620 B.n676 B.n394 163.367
R621 B.n680 B.n678 163.367
R622 B.n684 B.n392 163.367
R623 B.n688 B.n686 163.367
R624 B.n692 B.n390 163.367
R625 B.n696 B.n694 163.367
R626 B.n700 B.n388 163.367
R627 B.n703 B.n702 163.367
R628 B.n705 B.n385 163.367
R629 B.n709 B.n379 163.367
R630 B.n717 B.n379 163.367
R631 B.n717 B.n377 163.367
R632 B.n721 B.n377 163.367
R633 B.n721 B.n371 163.367
R634 B.n729 B.n371 163.367
R635 B.n729 B.n369 163.367
R636 B.n733 B.n369 163.367
R637 B.n733 B.n363 163.367
R638 B.n741 B.n363 163.367
R639 B.n741 B.n361 163.367
R640 B.n746 B.n361 163.367
R641 B.n746 B.n356 163.367
R642 B.n755 B.n356 163.367
R643 B.n756 B.n755 163.367
R644 B.n756 B.n5 163.367
R645 B.n6 B.n5 163.367
R646 B.n7 B.n6 163.367
R647 B.n761 B.n7 163.367
R648 B.n761 B.n12 163.367
R649 B.n13 B.n12 163.367
R650 B.n14 B.n13 163.367
R651 B.n766 B.n14 163.367
R652 B.n766 B.n19 163.367
R653 B.n20 B.n19 163.367
R654 B.n21 B.n20 163.367
R655 B.n771 B.n21 163.367
R656 B.n771 B.n26 163.367
R657 B.n27 B.n26 163.367
R658 B.n28 B.n27 163.367
R659 B.n776 B.n28 163.367
R660 B.n776 B.n33 163.367
R661 B.n104 B.n103 163.367
R662 B.n108 B.n107 163.367
R663 B.n112 B.n111 163.367
R664 B.n116 B.n115 163.367
R665 B.n120 B.n119 163.367
R666 B.n124 B.n123 163.367
R667 B.n128 B.n127 163.367
R668 B.n132 B.n131 163.367
R669 B.n136 B.n135 163.367
R670 B.n140 B.n139 163.367
R671 B.n144 B.n143 163.367
R672 B.n148 B.n147 163.367
R673 B.n152 B.n151 163.367
R674 B.n156 B.n155 163.367
R675 B.n160 B.n159 163.367
R676 B.n164 B.n163 163.367
R677 B.n168 B.n167 163.367
R678 B.n172 B.n171 163.367
R679 B.n176 B.n175 163.367
R680 B.n180 B.n179 163.367
R681 B.n184 B.n183 163.367
R682 B.n188 B.n187 163.367
R683 B.n192 B.n191 163.367
R684 B.n196 B.n195 163.367
R685 B.n200 B.n199 163.367
R686 B.n204 B.n203 163.367
R687 B.n208 B.n207 163.367
R688 B.n212 B.n211 163.367
R689 B.n216 B.n215 163.367
R690 B.n221 B.n220 163.367
R691 B.n225 B.n224 163.367
R692 B.n229 B.n228 163.367
R693 B.n233 B.n232 163.367
R694 B.n237 B.n236 163.367
R695 B.n242 B.n241 163.367
R696 B.n246 B.n245 163.367
R697 B.n250 B.n249 163.367
R698 B.n254 B.n253 163.367
R699 B.n258 B.n257 163.367
R700 B.n262 B.n261 163.367
R701 B.n266 B.n265 163.367
R702 B.n270 B.n269 163.367
R703 B.n274 B.n273 163.367
R704 B.n278 B.n277 163.367
R705 B.n282 B.n281 163.367
R706 B.n286 B.n285 163.367
R707 B.n290 B.n289 163.367
R708 B.n294 B.n293 163.367
R709 B.n298 B.n297 163.367
R710 B.n302 B.n301 163.367
R711 B.n306 B.n305 163.367
R712 B.n310 B.n309 163.367
R713 B.n314 B.n313 163.367
R714 B.n318 B.n317 163.367
R715 B.n322 B.n321 163.367
R716 B.n326 B.n325 163.367
R717 B.n330 B.n329 163.367
R718 B.n334 B.n333 163.367
R719 B.n338 B.n337 163.367
R720 B.n342 B.n341 163.367
R721 B.n346 B.n345 163.367
R722 B.n350 B.n349 163.367
R723 B.n352 B.n97 163.367
R724 B.n454 B.n383 71.676
R725 B.n460 B.n459 71.676
R726 B.n463 B.n462 71.676
R727 B.n468 B.n467 71.676
R728 B.n471 B.n470 71.676
R729 B.n476 B.n475 71.676
R730 B.n479 B.n478 71.676
R731 B.n484 B.n483 71.676
R732 B.n487 B.n486 71.676
R733 B.n492 B.n491 71.676
R734 B.n495 B.n494 71.676
R735 B.n500 B.n499 71.676
R736 B.n503 B.n502 71.676
R737 B.n508 B.n507 71.676
R738 B.n511 B.n510 71.676
R739 B.n516 B.n515 71.676
R740 B.n519 B.n518 71.676
R741 B.n524 B.n523 71.676
R742 B.n527 B.n526 71.676
R743 B.n532 B.n531 71.676
R744 B.n535 B.n534 71.676
R745 B.n540 B.n539 71.676
R746 B.n543 B.n542 71.676
R747 B.n548 B.n547 71.676
R748 B.n551 B.n550 71.676
R749 B.n556 B.n555 71.676
R750 B.n559 B.n558 71.676
R751 B.n564 B.n563 71.676
R752 B.n567 B.n566 71.676
R753 B.n573 B.n572 71.676
R754 B.n576 B.n575 71.676
R755 B.n581 B.n580 71.676
R756 B.n584 B.n583 71.676
R757 B.n589 B.n588 71.676
R758 B.n592 B.n591 71.676
R759 B.n597 B.n596 71.676
R760 B.n600 B.n599 71.676
R761 B.n605 B.n604 71.676
R762 B.n608 B.n607 71.676
R763 B.n613 B.n612 71.676
R764 B.n616 B.n615 71.676
R765 B.n621 B.n620 71.676
R766 B.n624 B.n623 71.676
R767 B.n629 B.n628 71.676
R768 B.n632 B.n631 71.676
R769 B.n637 B.n636 71.676
R770 B.n640 B.n639 71.676
R771 B.n645 B.n644 71.676
R772 B.n648 B.n647 71.676
R773 B.n653 B.n652 71.676
R774 B.n656 B.n655 71.676
R775 B.n661 B.n660 71.676
R776 B.n664 B.n663 71.676
R777 B.n669 B.n668 71.676
R778 B.n672 B.n671 71.676
R779 B.n677 B.n676 71.676
R780 B.n680 B.n679 71.676
R781 B.n685 B.n684 71.676
R782 B.n688 B.n687 71.676
R783 B.n693 B.n692 71.676
R784 B.n696 B.n695 71.676
R785 B.n701 B.n700 71.676
R786 B.n704 B.n703 71.676
R787 B.n34 B.n32 71.676
R788 B.n104 B.n35 71.676
R789 B.n108 B.n36 71.676
R790 B.n112 B.n37 71.676
R791 B.n116 B.n38 71.676
R792 B.n120 B.n39 71.676
R793 B.n124 B.n40 71.676
R794 B.n128 B.n41 71.676
R795 B.n132 B.n42 71.676
R796 B.n136 B.n43 71.676
R797 B.n140 B.n44 71.676
R798 B.n144 B.n45 71.676
R799 B.n148 B.n46 71.676
R800 B.n152 B.n47 71.676
R801 B.n156 B.n48 71.676
R802 B.n160 B.n49 71.676
R803 B.n164 B.n50 71.676
R804 B.n168 B.n51 71.676
R805 B.n172 B.n52 71.676
R806 B.n176 B.n53 71.676
R807 B.n180 B.n54 71.676
R808 B.n184 B.n55 71.676
R809 B.n188 B.n56 71.676
R810 B.n192 B.n57 71.676
R811 B.n196 B.n58 71.676
R812 B.n200 B.n59 71.676
R813 B.n204 B.n60 71.676
R814 B.n208 B.n61 71.676
R815 B.n212 B.n62 71.676
R816 B.n216 B.n63 71.676
R817 B.n221 B.n64 71.676
R818 B.n225 B.n65 71.676
R819 B.n229 B.n66 71.676
R820 B.n233 B.n67 71.676
R821 B.n237 B.n68 71.676
R822 B.n242 B.n69 71.676
R823 B.n246 B.n70 71.676
R824 B.n250 B.n71 71.676
R825 B.n254 B.n72 71.676
R826 B.n258 B.n73 71.676
R827 B.n262 B.n74 71.676
R828 B.n266 B.n75 71.676
R829 B.n270 B.n76 71.676
R830 B.n274 B.n77 71.676
R831 B.n278 B.n78 71.676
R832 B.n282 B.n79 71.676
R833 B.n286 B.n80 71.676
R834 B.n290 B.n81 71.676
R835 B.n294 B.n82 71.676
R836 B.n298 B.n83 71.676
R837 B.n302 B.n84 71.676
R838 B.n306 B.n85 71.676
R839 B.n310 B.n86 71.676
R840 B.n314 B.n87 71.676
R841 B.n318 B.n88 71.676
R842 B.n322 B.n89 71.676
R843 B.n326 B.n90 71.676
R844 B.n330 B.n91 71.676
R845 B.n334 B.n92 71.676
R846 B.n338 B.n93 71.676
R847 B.n342 B.n94 71.676
R848 B.n346 B.n95 71.676
R849 B.n350 B.n96 71.676
R850 B.n781 B.n97 71.676
R851 B.n781 B.n780 71.676
R852 B.n352 B.n96 71.676
R853 B.n349 B.n95 71.676
R854 B.n345 B.n94 71.676
R855 B.n341 B.n93 71.676
R856 B.n337 B.n92 71.676
R857 B.n333 B.n91 71.676
R858 B.n329 B.n90 71.676
R859 B.n325 B.n89 71.676
R860 B.n321 B.n88 71.676
R861 B.n317 B.n87 71.676
R862 B.n313 B.n86 71.676
R863 B.n309 B.n85 71.676
R864 B.n305 B.n84 71.676
R865 B.n301 B.n83 71.676
R866 B.n297 B.n82 71.676
R867 B.n293 B.n81 71.676
R868 B.n289 B.n80 71.676
R869 B.n285 B.n79 71.676
R870 B.n281 B.n78 71.676
R871 B.n277 B.n77 71.676
R872 B.n273 B.n76 71.676
R873 B.n269 B.n75 71.676
R874 B.n265 B.n74 71.676
R875 B.n261 B.n73 71.676
R876 B.n257 B.n72 71.676
R877 B.n253 B.n71 71.676
R878 B.n249 B.n70 71.676
R879 B.n245 B.n69 71.676
R880 B.n241 B.n68 71.676
R881 B.n236 B.n67 71.676
R882 B.n232 B.n66 71.676
R883 B.n228 B.n65 71.676
R884 B.n224 B.n64 71.676
R885 B.n220 B.n63 71.676
R886 B.n215 B.n62 71.676
R887 B.n211 B.n61 71.676
R888 B.n207 B.n60 71.676
R889 B.n203 B.n59 71.676
R890 B.n199 B.n58 71.676
R891 B.n195 B.n57 71.676
R892 B.n191 B.n56 71.676
R893 B.n187 B.n55 71.676
R894 B.n183 B.n54 71.676
R895 B.n179 B.n53 71.676
R896 B.n175 B.n52 71.676
R897 B.n171 B.n51 71.676
R898 B.n167 B.n50 71.676
R899 B.n163 B.n49 71.676
R900 B.n159 B.n48 71.676
R901 B.n155 B.n47 71.676
R902 B.n151 B.n46 71.676
R903 B.n147 B.n45 71.676
R904 B.n143 B.n44 71.676
R905 B.n139 B.n43 71.676
R906 B.n135 B.n42 71.676
R907 B.n131 B.n41 71.676
R908 B.n127 B.n40 71.676
R909 B.n123 B.n39 71.676
R910 B.n119 B.n38 71.676
R911 B.n115 B.n37 71.676
R912 B.n111 B.n36 71.676
R913 B.n107 B.n35 71.676
R914 B.n103 B.n34 71.676
R915 B.n455 B.n454 71.676
R916 B.n461 B.n460 71.676
R917 B.n462 B.n451 71.676
R918 B.n469 B.n468 71.676
R919 B.n470 B.n449 71.676
R920 B.n477 B.n476 71.676
R921 B.n478 B.n447 71.676
R922 B.n485 B.n484 71.676
R923 B.n486 B.n445 71.676
R924 B.n493 B.n492 71.676
R925 B.n494 B.n443 71.676
R926 B.n501 B.n500 71.676
R927 B.n502 B.n441 71.676
R928 B.n509 B.n508 71.676
R929 B.n510 B.n439 71.676
R930 B.n517 B.n516 71.676
R931 B.n518 B.n437 71.676
R932 B.n525 B.n524 71.676
R933 B.n526 B.n435 71.676
R934 B.n533 B.n532 71.676
R935 B.n534 B.n433 71.676
R936 B.n541 B.n540 71.676
R937 B.n542 B.n431 71.676
R938 B.n549 B.n548 71.676
R939 B.n550 B.n429 71.676
R940 B.n557 B.n556 71.676
R941 B.n558 B.n427 71.676
R942 B.n565 B.n564 71.676
R943 B.n566 B.n423 71.676
R944 B.n574 B.n573 71.676
R945 B.n575 B.n421 71.676
R946 B.n582 B.n581 71.676
R947 B.n583 B.n419 71.676
R948 B.n590 B.n589 71.676
R949 B.n591 B.n414 71.676
R950 B.n598 B.n597 71.676
R951 B.n599 B.n412 71.676
R952 B.n606 B.n605 71.676
R953 B.n607 B.n410 71.676
R954 B.n614 B.n613 71.676
R955 B.n615 B.n408 71.676
R956 B.n622 B.n621 71.676
R957 B.n623 B.n406 71.676
R958 B.n630 B.n629 71.676
R959 B.n631 B.n404 71.676
R960 B.n638 B.n637 71.676
R961 B.n639 B.n402 71.676
R962 B.n646 B.n645 71.676
R963 B.n647 B.n400 71.676
R964 B.n654 B.n653 71.676
R965 B.n655 B.n398 71.676
R966 B.n662 B.n661 71.676
R967 B.n663 B.n396 71.676
R968 B.n670 B.n669 71.676
R969 B.n671 B.n394 71.676
R970 B.n678 B.n677 71.676
R971 B.n679 B.n392 71.676
R972 B.n686 B.n685 71.676
R973 B.n687 B.n390 71.676
R974 B.n694 B.n693 71.676
R975 B.n695 B.n388 71.676
R976 B.n702 B.n701 71.676
R977 B.n705 B.n704 71.676
R978 B.n417 B.n416 59.5399
R979 B.n570 B.n425 59.5399
R980 B.n218 B.n101 59.5399
R981 B.n239 B.n99 59.5399
R982 B.n710 B.n384 57.0882
R983 B.n783 B.n782 57.0882
R984 B.n785 B.n31 33.8737
R985 B.n779 B.n778 33.8737
R986 B.n708 B.n707 33.8737
R987 B.n712 B.n382 33.8737
R988 B.n710 B.n380 32.0828
R989 B.n716 B.n380 32.0828
R990 B.n716 B.n376 32.0828
R991 B.n722 B.n376 32.0828
R992 B.n728 B.n372 32.0828
R993 B.n728 B.n368 32.0828
R994 B.n734 B.n368 32.0828
R995 B.n734 B.n364 32.0828
R996 B.n740 B.n364 32.0828
R997 B.n748 B.n360 32.0828
R998 B.n748 B.n747 32.0828
R999 B.n754 B.n4 32.0828
R1000 B.n815 B.n4 32.0828
R1001 B.n815 B.n814 32.0828
R1002 B.n814 B.n813 32.0828
R1003 B.n807 B.n11 32.0828
R1004 B.n807 B.n806 32.0828
R1005 B.n805 B.n15 32.0828
R1006 B.n799 B.n15 32.0828
R1007 B.n799 B.n798 32.0828
R1008 B.n798 B.n797 32.0828
R1009 B.n797 B.n22 32.0828
R1010 B.n791 B.n790 32.0828
R1011 B.n790 B.n789 32.0828
R1012 B.n789 B.n29 32.0828
R1013 B.n783 B.n29 32.0828
R1014 B.n754 B.t3 29.2521
R1015 B.n813 B.t2 29.2521
R1016 B.n722 B.t9 20.7597
R1017 B.n791 B.t5 20.7597
R1018 B B.n817 18.0485
R1019 B.n416 B.n415 17.2611
R1020 B.n425 B.n424 17.2611
R1021 B.n101 B.n100 17.2611
R1022 B.n99 B.n98 17.2611
R1023 B.t1 B.n360 16.9853
R1024 B.n806 B.t0 16.9853
R1025 B.n740 B.t1 15.0981
R1026 B.t0 B.n805 15.0981
R1027 B.t9 B.n372 11.3237
R1028 B.t5 B.n22 11.3237
R1029 B.n102 B.n31 10.6151
R1030 B.n105 B.n102 10.6151
R1031 B.n106 B.n105 10.6151
R1032 B.n109 B.n106 10.6151
R1033 B.n110 B.n109 10.6151
R1034 B.n113 B.n110 10.6151
R1035 B.n114 B.n113 10.6151
R1036 B.n117 B.n114 10.6151
R1037 B.n118 B.n117 10.6151
R1038 B.n121 B.n118 10.6151
R1039 B.n122 B.n121 10.6151
R1040 B.n125 B.n122 10.6151
R1041 B.n126 B.n125 10.6151
R1042 B.n129 B.n126 10.6151
R1043 B.n130 B.n129 10.6151
R1044 B.n133 B.n130 10.6151
R1045 B.n134 B.n133 10.6151
R1046 B.n137 B.n134 10.6151
R1047 B.n138 B.n137 10.6151
R1048 B.n141 B.n138 10.6151
R1049 B.n142 B.n141 10.6151
R1050 B.n145 B.n142 10.6151
R1051 B.n146 B.n145 10.6151
R1052 B.n149 B.n146 10.6151
R1053 B.n150 B.n149 10.6151
R1054 B.n153 B.n150 10.6151
R1055 B.n154 B.n153 10.6151
R1056 B.n157 B.n154 10.6151
R1057 B.n158 B.n157 10.6151
R1058 B.n161 B.n158 10.6151
R1059 B.n162 B.n161 10.6151
R1060 B.n165 B.n162 10.6151
R1061 B.n166 B.n165 10.6151
R1062 B.n169 B.n166 10.6151
R1063 B.n170 B.n169 10.6151
R1064 B.n173 B.n170 10.6151
R1065 B.n174 B.n173 10.6151
R1066 B.n177 B.n174 10.6151
R1067 B.n178 B.n177 10.6151
R1068 B.n181 B.n178 10.6151
R1069 B.n182 B.n181 10.6151
R1070 B.n185 B.n182 10.6151
R1071 B.n186 B.n185 10.6151
R1072 B.n189 B.n186 10.6151
R1073 B.n190 B.n189 10.6151
R1074 B.n193 B.n190 10.6151
R1075 B.n194 B.n193 10.6151
R1076 B.n197 B.n194 10.6151
R1077 B.n198 B.n197 10.6151
R1078 B.n201 B.n198 10.6151
R1079 B.n202 B.n201 10.6151
R1080 B.n205 B.n202 10.6151
R1081 B.n206 B.n205 10.6151
R1082 B.n209 B.n206 10.6151
R1083 B.n210 B.n209 10.6151
R1084 B.n213 B.n210 10.6151
R1085 B.n214 B.n213 10.6151
R1086 B.n217 B.n214 10.6151
R1087 B.n222 B.n219 10.6151
R1088 B.n223 B.n222 10.6151
R1089 B.n226 B.n223 10.6151
R1090 B.n227 B.n226 10.6151
R1091 B.n230 B.n227 10.6151
R1092 B.n231 B.n230 10.6151
R1093 B.n234 B.n231 10.6151
R1094 B.n235 B.n234 10.6151
R1095 B.n238 B.n235 10.6151
R1096 B.n243 B.n240 10.6151
R1097 B.n244 B.n243 10.6151
R1098 B.n247 B.n244 10.6151
R1099 B.n248 B.n247 10.6151
R1100 B.n251 B.n248 10.6151
R1101 B.n252 B.n251 10.6151
R1102 B.n255 B.n252 10.6151
R1103 B.n256 B.n255 10.6151
R1104 B.n259 B.n256 10.6151
R1105 B.n260 B.n259 10.6151
R1106 B.n263 B.n260 10.6151
R1107 B.n264 B.n263 10.6151
R1108 B.n267 B.n264 10.6151
R1109 B.n268 B.n267 10.6151
R1110 B.n271 B.n268 10.6151
R1111 B.n272 B.n271 10.6151
R1112 B.n275 B.n272 10.6151
R1113 B.n276 B.n275 10.6151
R1114 B.n279 B.n276 10.6151
R1115 B.n280 B.n279 10.6151
R1116 B.n283 B.n280 10.6151
R1117 B.n284 B.n283 10.6151
R1118 B.n287 B.n284 10.6151
R1119 B.n288 B.n287 10.6151
R1120 B.n291 B.n288 10.6151
R1121 B.n292 B.n291 10.6151
R1122 B.n295 B.n292 10.6151
R1123 B.n296 B.n295 10.6151
R1124 B.n299 B.n296 10.6151
R1125 B.n300 B.n299 10.6151
R1126 B.n303 B.n300 10.6151
R1127 B.n304 B.n303 10.6151
R1128 B.n307 B.n304 10.6151
R1129 B.n308 B.n307 10.6151
R1130 B.n311 B.n308 10.6151
R1131 B.n312 B.n311 10.6151
R1132 B.n315 B.n312 10.6151
R1133 B.n316 B.n315 10.6151
R1134 B.n319 B.n316 10.6151
R1135 B.n320 B.n319 10.6151
R1136 B.n323 B.n320 10.6151
R1137 B.n324 B.n323 10.6151
R1138 B.n327 B.n324 10.6151
R1139 B.n328 B.n327 10.6151
R1140 B.n331 B.n328 10.6151
R1141 B.n332 B.n331 10.6151
R1142 B.n335 B.n332 10.6151
R1143 B.n336 B.n335 10.6151
R1144 B.n339 B.n336 10.6151
R1145 B.n340 B.n339 10.6151
R1146 B.n343 B.n340 10.6151
R1147 B.n344 B.n343 10.6151
R1148 B.n347 B.n344 10.6151
R1149 B.n348 B.n347 10.6151
R1150 B.n351 B.n348 10.6151
R1151 B.n353 B.n351 10.6151
R1152 B.n354 B.n353 10.6151
R1153 B.n779 B.n354 10.6151
R1154 B.n708 B.n378 10.6151
R1155 B.n718 B.n378 10.6151
R1156 B.n719 B.n718 10.6151
R1157 B.n720 B.n719 10.6151
R1158 B.n720 B.n370 10.6151
R1159 B.n730 B.n370 10.6151
R1160 B.n731 B.n730 10.6151
R1161 B.n732 B.n731 10.6151
R1162 B.n732 B.n362 10.6151
R1163 B.n742 B.n362 10.6151
R1164 B.n743 B.n742 10.6151
R1165 B.n745 B.n743 10.6151
R1166 B.n745 B.n744 10.6151
R1167 B.n744 B.n355 10.6151
R1168 B.n757 B.n355 10.6151
R1169 B.n758 B.n757 10.6151
R1170 B.n759 B.n758 10.6151
R1171 B.n760 B.n759 10.6151
R1172 B.n762 B.n760 10.6151
R1173 B.n763 B.n762 10.6151
R1174 B.n764 B.n763 10.6151
R1175 B.n765 B.n764 10.6151
R1176 B.n767 B.n765 10.6151
R1177 B.n768 B.n767 10.6151
R1178 B.n769 B.n768 10.6151
R1179 B.n770 B.n769 10.6151
R1180 B.n772 B.n770 10.6151
R1181 B.n773 B.n772 10.6151
R1182 B.n774 B.n773 10.6151
R1183 B.n775 B.n774 10.6151
R1184 B.n777 B.n775 10.6151
R1185 B.n778 B.n777 10.6151
R1186 B.n456 B.n382 10.6151
R1187 B.n457 B.n456 10.6151
R1188 B.n458 B.n457 10.6151
R1189 B.n458 B.n452 10.6151
R1190 B.n464 B.n452 10.6151
R1191 B.n465 B.n464 10.6151
R1192 B.n466 B.n465 10.6151
R1193 B.n466 B.n450 10.6151
R1194 B.n472 B.n450 10.6151
R1195 B.n473 B.n472 10.6151
R1196 B.n474 B.n473 10.6151
R1197 B.n474 B.n448 10.6151
R1198 B.n480 B.n448 10.6151
R1199 B.n481 B.n480 10.6151
R1200 B.n482 B.n481 10.6151
R1201 B.n482 B.n446 10.6151
R1202 B.n488 B.n446 10.6151
R1203 B.n489 B.n488 10.6151
R1204 B.n490 B.n489 10.6151
R1205 B.n490 B.n444 10.6151
R1206 B.n496 B.n444 10.6151
R1207 B.n497 B.n496 10.6151
R1208 B.n498 B.n497 10.6151
R1209 B.n498 B.n442 10.6151
R1210 B.n504 B.n442 10.6151
R1211 B.n505 B.n504 10.6151
R1212 B.n506 B.n505 10.6151
R1213 B.n506 B.n440 10.6151
R1214 B.n512 B.n440 10.6151
R1215 B.n513 B.n512 10.6151
R1216 B.n514 B.n513 10.6151
R1217 B.n514 B.n438 10.6151
R1218 B.n520 B.n438 10.6151
R1219 B.n521 B.n520 10.6151
R1220 B.n522 B.n521 10.6151
R1221 B.n522 B.n436 10.6151
R1222 B.n528 B.n436 10.6151
R1223 B.n529 B.n528 10.6151
R1224 B.n530 B.n529 10.6151
R1225 B.n530 B.n434 10.6151
R1226 B.n536 B.n434 10.6151
R1227 B.n537 B.n536 10.6151
R1228 B.n538 B.n537 10.6151
R1229 B.n538 B.n432 10.6151
R1230 B.n544 B.n432 10.6151
R1231 B.n545 B.n544 10.6151
R1232 B.n546 B.n545 10.6151
R1233 B.n546 B.n430 10.6151
R1234 B.n552 B.n430 10.6151
R1235 B.n553 B.n552 10.6151
R1236 B.n554 B.n553 10.6151
R1237 B.n554 B.n428 10.6151
R1238 B.n560 B.n428 10.6151
R1239 B.n561 B.n560 10.6151
R1240 B.n562 B.n561 10.6151
R1241 B.n562 B.n426 10.6151
R1242 B.n568 B.n426 10.6151
R1243 B.n569 B.n568 10.6151
R1244 B.n571 B.n422 10.6151
R1245 B.n577 B.n422 10.6151
R1246 B.n578 B.n577 10.6151
R1247 B.n579 B.n578 10.6151
R1248 B.n579 B.n420 10.6151
R1249 B.n585 B.n420 10.6151
R1250 B.n586 B.n585 10.6151
R1251 B.n587 B.n586 10.6151
R1252 B.n587 B.n418 10.6151
R1253 B.n594 B.n593 10.6151
R1254 B.n595 B.n594 10.6151
R1255 B.n595 B.n413 10.6151
R1256 B.n601 B.n413 10.6151
R1257 B.n602 B.n601 10.6151
R1258 B.n603 B.n602 10.6151
R1259 B.n603 B.n411 10.6151
R1260 B.n609 B.n411 10.6151
R1261 B.n610 B.n609 10.6151
R1262 B.n611 B.n610 10.6151
R1263 B.n611 B.n409 10.6151
R1264 B.n617 B.n409 10.6151
R1265 B.n618 B.n617 10.6151
R1266 B.n619 B.n618 10.6151
R1267 B.n619 B.n407 10.6151
R1268 B.n625 B.n407 10.6151
R1269 B.n626 B.n625 10.6151
R1270 B.n627 B.n626 10.6151
R1271 B.n627 B.n405 10.6151
R1272 B.n633 B.n405 10.6151
R1273 B.n634 B.n633 10.6151
R1274 B.n635 B.n634 10.6151
R1275 B.n635 B.n403 10.6151
R1276 B.n641 B.n403 10.6151
R1277 B.n642 B.n641 10.6151
R1278 B.n643 B.n642 10.6151
R1279 B.n643 B.n401 10.6151
R1280 B.n649 B.n401 10.6151
R1281 B.n650 B.n649 10.6151
R1282 B.n651 B.n650 10.6151
R1283 B.n651 B.n399 10.6151
R1284 B.n657 B.n399 10.6151
R1285 B.n658 B.n657 10.6151
R1286 B.n659 B.n658 10.6151
R1287 B.n659 B.n397 10.6151
R1288 B.n665 B.n397 10.6151
R1289 B.n666 B.n665 10.6151
R1290 B.n667 B.n666 10.6151
R1291 B.n667 B.n395 10.6151
R1292 B.n673 B.n395 10.6151
R1293 B.n674 B.n673 10.6151
R1294 B.n675 B.n674 10.6151
R1295 B.n675 B.n393 10.6151
R1296 B.n681 B.n393 10.6151
R1297 B.n682 B.n681 10.6151
R1298 B.n683 B.n682 10.6151
R1299 B.n683 B.n391 10.6151
R1300 B.n689 B.n391 10.6151
R1301 B.n690 B.n689 10.6151
R1302 B.n691 B.n690 10.6151
R1303 B.n691 B.n389 10.6151
R1304 B.n697 B.n389 10.6151
R1305 B.n698 B.n697 10.6151
R1306 B.n699 B.n698 10.6151
R1307 B.n699 B.n387 10.6151
R1308 B.n387 B.n386 10.6151
R1309 B.n706 B.n386 10.6151
R1310 B.n707 B.n706 10.6151
R1311 B.n713 B.n712 10.6151
R1312 B.n714 B.n713 10.6151
R1313 B.n714 B.n374 10.6151
R1314 B.n724 B.n374 10.6151
R1315 B.n725 B.n724 10.6151
R1316 B.n726 B.n725 10.6151
R1317 B.n726 B.n366 10.6151
R1318 B.n736 B.n366 10.6151
R1319 B.n737 B.n736 10.6151
R1320 B.n738 B.n737 10.6151
R1321 B.n738 B.n358 10.6151
R1322 B.n750 B.n358 10.6151
R1323 B.n751 B.n750 10.6151
R1324 B.n752 B.n751 10.6151
R1325 B.n752 B.n0 10.6151
R1326 B.n811 B.n1 10.6151
R1327 B.n811 B.n810 10.6151
R1328 B.n810 B.n809 10.6151
R1329 B.n809 B.n9 10.6151
R1330 B.n803 B.n9 10.6151
R1331 B.n803 B.n802 10.6151
R1332 B.n802 B.n801 10.6151
R1333 B.n801 B.n17 10.6151
R1334 B.n795 B.n17 10.6151
R1335 B.n795 B.n794 10.6151
R1336 B.n794 B.n793 10.6151
R1337 B.n793 B.n24 10.6151
R1338 B.n787 B.n24 10.6151
R1339 B.n787 B.n786 10.6151
R1340 B.n786 B.n785 10.6151
R1341 B.n218 B.n217 9.36635
R1342 B.n240 B.n239 9.36635
R1343 B.n570 B.n569 9.36635
R1344 B.n593 B.n417 9.36635
R1345 B.n747 B.t3 2.8313
R1346 B.n11 B.t2 2.8313
R1347 B.n817 B.n0 2.81026
R1348 B.n817 B.n1 2.81026
R1349 B.n219 B.n218 1.24928
R1350 B.n239 B.n238 1.24928
R1351 B.n571 B.n570 1.24928
R1352 B.n418 B.n417 1.24928
R1353 VP.n0 VP.t1 867.495
R1354 VP.n0 VP.t2 867.471
R1355 VP.n2 VP.t3 846.514
R1356 VP.n3 VP.t0 846.514
R1357 VP.n4 VP.n3 161.3
R1358 VP.n2 VP.n1 161.3
R1359 VP.n1 VP.n0 114.858
R1360 VP.n3 VP.n2 48.2005
R1361 VP.n4 VP.n1 0.189894
R1362 VP VP.n4 0.0516364
R1363 VTAIL.n798 VTAIL.n797 289.615
R1364 VTAIL.n98 VTAIL.n97 289.615
R1365 VTAIL.n198 VTAIL.n197 289.615
R1366 VTAIL.n298 VTAIL.n297 289.615
R1367 VTAIL.n698 VTAIL.n697 289.615
R1368 VTAIL.n598 VTAIL.n597 289.615
R1369 VTAIL.n498 VTAIL.n497 289.615
R1370 VTAIL.n398 VTAIL.n397 289.615
R1371 VTAIL.n733 VTAIL.n732 185
R1372 VTAIL.n730 VTAIL.n729 185
R1373 VTAIL.n739 VTAIL.n738 185
R1374 VTAIL.n741 VTAIL.n740 185
R1375 VTAIL.n726 VTAIL.n725 185
R1376 VTAIL.n747 VTAIL.n746 185
R1377 VTAIL.n750 VTAIL.n749 185
R1378 VTAIL.n748 VTAIL.n722 185
R1379 VTAIL.n755 VTAIL.n721 185
R1380 VTAIL.n757 VTAIL.n756 185
R1381 VTAIL.n759 VTAIL.n758 185
R1382 VTAIL.n718 VTAIL.n717 185
R1383 VTAIL.n765 VTAIL.n764 185
R1384 VTAIL.n767 VTAIL.n766 185
R1385 VTAIL.n714 VTAIL.n713 185
R1386 VTAIL.n773 VTAIL.n772 185
R1387 VTAIL.n775 VTAIL.n774 185
R1388 VTAIL.n710 VTAIL.n709 185
R1389 VTAIL.n781 VTAIL.n780 185
R1390 VTAIL.n783 VTAIL.n782 185
R1391 VTAIL.n706 VTAIL.n705 185
R1392 VTAIL.n789 VTAIL.n788 185
R1393 VTAIL.n791 VTAIL.n790 185
R1394 VTAIL.n702 VTAIL.n701 185
R1395 VTAIL.n797 VTAIL.n796 185
R1396 VTAIL.n33 VTAIL.n32 185
R1397 VTAIL.n30 VTAIL.n29 185
R1398 VTAIL.n39 VTAIL.n38 185
R1399 VTAIL.n41 VTAIL.n40 185
R1400 VTAIL.n26 VTAIL.n25 185
R1401 VTAIL.n47 VTAIL.n46 185
R1402 VTAIL.n50 VTAIL.n49 185
R1403 VTAIL.n48 VTAIL.n22 185
R1404 VTAIL.n55 VTAIL.n21 185
R1405 VTAIL.n57 VTAIL.n56 185
R1406 VTAIL.n59 VTAIL.n58 185
R1407 VTAIL.n18 VTAIL.n17 185
R1408 VTAIL.n65 VTAIL.n64 185
R1409 VTAIL.n67 VTAIL.n66 185
R1410 VTAIL.n14 VTAIL.n13 185
R1411 VTAIL.n73 VTAIL.n72 185
R1412 VTAIL.n75 VTAIL.n74 185
R1413 VTAIL.n10 VTAIL.n9 185
R1414 VTAIL.n81 VTAIL.n80 185
R1415 VTAIL.n83 VTAIL.n82 185
R1416 VTAIL.n6 VTAIL.n5 185
R1417 VTAIL.n89 VTAIL.n88 185
R1418 VTAIL.n91 VTAIL.n90 185
R1419 VTAIL.n2 VTAIL.n1 185
R1420 VTAIL.n97 VTAIL.n96 185
R1421 VTAIL.n133 VTAIL.n132 185
R1422 VTAIL.n130 VTAIL.n129 185
R1423 VTAIL.n139 VTAIL.n138 185
R1424 VTAIL.n141 VTAIL.n140 185
R1425 VTAIL.n126 VTAIL.n125 185
R1426 VTAIL.n147 VTAIL.n146 185
R1427 VTAIL.n150 VTAIL.n149 185
R1428 VTAIL.n148 VTAIL.n122 185
R1429 VTAIL.n155 VTAIL.n121 185
R1430 VTAIL.n157 VTAIL.n156 185
R1431 VTAIL.n159 VTAIL.n158 185
R1432 VTAIL.n118 VTAIL.n117 185
R1433 VTAIL.n165 VTAIL.n164 185
R1434 VTAIL.n167 VTAIL.n166 185
R1435 VTAIL.n114 VTAIL.n113 185
R1436 VTAIL.n173 VTAIL.n172 185
R1437 VTAIL.n175 VTAIL.n174 185
R1438 VTAIL.n110 VTAIL.n109 185
R1439 VTAIL.n181 VTAIL.n180 185
R1440 VTAIL.n183 VTAIL.n182 185
R1441 VTAIL.n106 VTAIL.n105 185
R1442 VTAIL.n189 VTAIL.n188 185
R1443 VTAIL.n191 VTAIL.n190 185
R1444 VTAIL.n102 VTAIL.n101 185
R1445 VTAIL.n197 VTAIL.n196 185
R1446 VTAIL.n233 VTAIL.n232 185
R1447 VTAIL.n230 VTAIL.n229 185
R1448 VTAIL.n239 VTAIL.n238 185
R1449 VTAIL.n241 VTAIL.n240 185
R1450 VTAIL.n226 VTAIL.n225 185
R1451 VTAIL.n247 VTAIL.n246 185
R1452 VTAIL.n250 VTAIL.n249 185
R1453 VTAIL.n248 VTAIL.n222 185
R1454 VTAIL.n255 VTAIL.n221 185
R1455 VTAIL.n257 VTAIL.n256 185
R1456 VTAIL.n259 VTAIL.n258 185
R1457 VTAIL.n218 VTAIL.n217 185
R1458 VTAIL.n265 VTAIL.n264 185
R1459 VTAIL.n267 VTAIL.n266 185
R1460 VTAIL.n214 VTAIL.n213 185
R1461 VTAIL.n273 VTAIL.n272 185
R1462 VTAIL.n275 VTAIL.n274 185
R1463 VTAIL.n210 VTAIL.n209 185
R1464 VTAIL.n281 VTAIL.n280 185
R1465 VTAIL.n283 VTAIL.n282 185
R1466 VTAIL.n206 VTAIL.n205 185
R1467 VTAIL.n289 VTAIL.n288 185
R1468 VTAIL.n291 VTAIL.n290 185
R1469 VTAIL.n202 VTAIL.n201 185
R1470 VTAIL.n297 VTAIL.n296 185
R1471 VTAIL.n697 VTAIL.n696 185
R1472 VTAIL.n602 VTAIL.n601 185
R1473 VTAIL.n691 VTAIL.n690 185
R1474 VTAIL.n689 VTAIL.n688 185
R1475 VTAIL.n606 VTAIL.n605 185
R1476 VTAIL.n683 VTAIL.n682 185
R1477 VTAIL.n681 VTAIL.n680 185
R1478 VTAIL.n610 VTAIL.n609 185
R1479 VTAIL.n675 VTAIL.n674 185
R1480 VTAIL.n673 VTAIL.n672 185
R1481 VTAIL.n614 VTAIL.n613 185
R1482 VTAIL.n667 VTAIL.n666 185
R1483 VTAIL.n665 VTAIL.n664 185
R1484 VTAIL.n618 VTAIL.n617 185
R1485 VTAIL.n659 VTAIL.n658 185
R1486 VTAIL.n657 VTAIL.n656 185
R1487 VTAIL.n655 VTAIL.n621 185
R1488 VTAIL.n625 VTAIL.n622 185
R1489 VTAIL.n650 VTAIL.n649 185
R1490 VTAIL.n648 VTAIL.n647 185
R1491 VTAIL.n627 VTAIL.n626 185
R1492 VTAIL.n642 VTAIL.n641 185
R1493 VTAIL.n640 VTAIL.n639 185
R1494 VTAIL.n631 VTAIL.n630 185
R1495 VTAIL.n634 VTAIL.n633 185
R1496 VTAIL.n597 VTAIL.n596 185
R1497 VTAIL.n502 VTAIL.n501 185
R1498 VTAIL.n591 VTAIL.n590 185
R1499 VTAIL.n589 VTAIL.n588 185
R1500 VTAIL.n506 VTAIL.n505 185
R1501 VTAIL.n583 VTAIL.n582 185
R1502 VTAIL.n581 VTAIL.n580 185
R1503 VTAIL.n510 VTAIL.n509 185
R1504 VTAIL.n575 VTAIL.n574 185
R1505 VTAIL.n573 VTAIL.n572 185
R1506 VTAIL.n514 VTAIL.n513 185
R1507 VTAIL.n567 VTAIL.n566 185
R1508 VTAIL.n565 VTAIL.n564 185
R1509 VTAIL.n518 VTAIL.n517 185
R1510 VTAIL.n559 VTAIL.n558 185
R1511 VTAIL.n557 VTAIL.n556 185
R1512 VTAIL.n555 VTAIL.n521 185
R1513 VTAIL.n525 VTAIL.n522 185
R1514 VTAIL.n550 VTAIL.n549 185
R1515 VTAIL.n548 VTAIL.n547 185
R1516 VTAIL.n527 VTAIL.n526 185
R1517 VTAIL.n542 VTAIL.n541 185
R1518 VTAIL.n540 VTAIL.n539 185
R1519 VTAIL.n531 VTAIL.n530 185
R1520 VTAIL.n534 VTAIL.n533 185
R1521 VTAIL.n497 VTAIL.n496 185
R1522 VTAIL.n402 VTAIL.n401 185
R1523 VTAIL.n491 VTAIL.n490 185
R1524 VTAIL.n489 VTAIL.n488 185
R1525 VTAIL.n406 VTAIL.n405 185
R1526 VTAIL.n483 VTAIL.n482 185
R1527 VTAIL.n481 VTAIL.n480 185
R1528 VTAIL.n410 VTAIL.n409 185
R1529 VTAIL.n475 VTAIL.n474 185
R1530 VTAIL.n473 VTAIL.n472 185
R1531 VTAIL.n414 VTAIL.n413 185
R1532 VTAIL.n467 VTAIL.n466 185
R1533 VTAIL.n465 VTAIL.n464 185
R1534 VTAIL.n418 VTAIL.n417 185
R1535 VTAIL.n459 VTAIL.n458 185
R1536 VTAIL.n457 VTAIL.n456 185
R1537 VTAIL.n455 VTAIL.n421 185
R1538 VTAIL.n425 VTAIL.n422 185
R1539 VTAIL.n450 VTAIL.n449 185
R1540 VTAIL.n448 VTAIL.n447 185
R1541 VTAIL.n427 VTAIL.n426 185
R1542 VTAIL.n442 VTAIL.n441 185
R1543 VTAIL.n440 VTAIL.n439 185
R1544 VTAIL.n431 VTAIL.n430 185
R1545 VTAIL.n434 VTAIL.n433 185
R1546 VTAIL.n397 VTAIL.n396 185
R1547 VTAIL.n302 VTAIL.n301 185
R1548 VTAIL.n391 VTAIL.n390 185
R1549 VTAIL.n389 VTAIL.n388 185
R1550 VTAIL.n306 VTAIL.n305 185
R1551 VTAIL.n383 VTAIL.n382 185
R1552 VTAIL.n381 VTAIL.n380 185
R1553 VTAIL.n310 VTAIL.n309 185
R1554 VTAIL.n375 VTAIL.n374 185
R1555 VTAIL.n373 VTAIL.n372 185
R1556 VTAIL.n314 VTAIL.n313 185
R1557 VTAIL.n367 VTAIL.n366 185
R1558 VTAIL.n365 VTAIL.n364 185
R1559 VTAIL.n318 VTAIL.n317 185
R1560 VTAIL.n359 VTAIL.n358 185
R1561 VTAIL.n357 VTAIL.n356 185
R1562 VTAIL.n355 VTAIL.n321 185
R1563 VTAIL.n325 VTAIL.n322 185
R1564 VTAIL.n350 VTAIL.n349 185
R1565 VTAIL.n348 VTAIL.n347 185
R1566 VTAIL.n327 VTAIL.n326 185
R1567 VTAIL.n342 VTAIL.n341 185
R1568 VTAIL.n340 VTAIL.n339 185
R1569 VTAIL.n331 VTAIL.n330 185
R1570 VTAIL.n334 VTAIL.n333 185
R1571 VTAIL.t1 VTAIL.n731 149.524
R1572 VTAIL.t2 VTAIL.n31 149.524
R1573 VTAIL.t7 VTAIL.n131 149.524
R1574 VTAIL.t4 VTAIL.n231 149.524
R1575 VTAIL.t5 VTAIL.n632 149.524
R1576 VTAIL.t6 VTAIL.n532 149.524
R1577 VTAIL.t3 VTAIL.n432 149.524
R1578 VTAIL.t0 VTAIL.n332 149.524
R1579 VTAIL.n732 VTAIL.n729 104.615
R1580 VTAIL.n739 VTAIL.n729 104.615
R1581 VTAIL.n740 VTAIL.n739 104.615
R1582 VTAIL.n740 VTAIL.n725 104.615
R1583 VTAIL.n747 VTAIL.n725 104.615
R1584 VTAIL.n749 VTAIL.n747 104.615
R1585 VTAIL.n749 VTAIL.n748 104.615
R1586 VTAIL.n748 VTAIL.n721 104.615
R1587 VTAIL.n757 VTAIL.n721 104.615
R1588 VTAIL.n758 VTAIL.n757 104.615
R1589 VTAIL.n758 VTAIL.n717 104.615
R1590 VTAIL.n765 VTAIL.n717 104.615
R1591 VTAIL.n766 VTAIL.n765 104.615
R1592 VTAIL.n766 VTAIL.n713 104.615
R1593 VTAIL.n773 VTAIL.n713 104.615
R1594 VTAIL.n774 VTAIL.n773 104.615
R1595 VTAIL.n774 VTAIL.n709 104.615
R1596 VTAIL.n781 VTAIL.n709 104.615
R1597 VTAIL.n782 VTAIL.n781 104.615
R1598 VTAIL.n782 VTAIL.n705 104.615
R1599 VTAIL.n789 VTAIL.n705 104.615
R1600 VTAIL.n790 VTAIL.n789 104.615
R1601 VTAIL.n790 VTAIL.n701 104.615
R1602 VTAIL.n797 VTAIL.n701 104.615
R1603 VTAIL.n32 VTAIL.n29 104.615
R1604 VTAIL.n39 VTAIL.n29 104.615
R1605 VTAIL.n40 VTAIL.n39 104.615
R1606 VTAIL.n40 VTAIL.n25 104.615
R1607 VTAIL.n47 VTAIL.n25 104.615
R1608 VTAIL.n49 VTAIL.n47 104.615
R1609 VTAIL.n49 VTAIL.n48 104.615
R1610 VTAIL.n48 VTAIL.n21 104.615
R1611 VTAIL.n57 VTAIL.n21 104.615
R1612 VTAIL.n58 VTAIL.n57 104.615
R1613 VTAIL.n58 VTAIL.n17 104.615
R1614 VTAIL.n65 VTAIL.n17 104.615
R1615 VTAIL.n66 VTAIL.n65 104.615
R1616 VTAIL.n66 VTAIL.n13 104.615
R1617 VTAIL.n73 VTAIL.n13 104.615
R1618 VTAIL.n74 VTAIL.n73 104.615
R1619 VTAIL.n74 VTAIL.n9 104.615
R1620 VTAIL.n81 VTAIL.n9 104.615
R1621 VTAIL.n82 VTAIL.n81 104.615
R1622 VTAIL.n82 VTAIL.n5 104.615
R1623 VTAIL.n89 VTAIL.n5 104.615
R1624 VTAIL.n90 VTAIL.n89 104.615
R1625 VTAIL.n90 VTAIL.n1 104.615
R1626 VTAIL.n97 VTAIL.n1 104.615
R1627 VTAIL.n132 VTAIL.n129 104.615
R1628 VTAIL.n139 VTAIL.n129 104.615
R1629 VTAIL.n140 VTAIL.n139 104.615
R1630 VTAIL.n140 VTAIL.n125 104.615
R1631 VTAIL.n147 VTAIL.n125 104.615
R1632 VTAIL.n149 VTAIL.n147 104.615
R1633 VTAIL.n149 VTAIL.n148 104.615
R1634 VTAIL.n148 VTAIL.n121 104.615
R1635 VTAIL.n157 VTAIL.n121 104.615
R1636 VTAIL.n158 VTAIL.n157 104.615
R1637 VTAIL.n158 VTAIL.n117 104.615
R1638 VTAIL.n165 VTAIL.n117 104.615
R1639 VTAIL.n166 VTAIL.n165 104.615
R1640 VTAIL.n166 VTAIL.n113 104.615
R1641 VTAIL.n173 VTAIL.n113 104.615
R1642 VTAIL.n174 VTAIL.n173 104.615
R1643 VTAIL.n174 VTAIL.n109 104.615
R1644 VTAIL.n181 VTAIL.n109 104.615
R1645 VTAIL.n182 VTAIL.n181 104.615
R1646 VTAIL.n182 VTAIL.n105 104.615
R1647 VTAIL.n189 VTAIL.n105 104.615
R1648 VTAIL.n190 VTAIL.n189 104.615
R1649 VTAIL.n190 VTAIL.n101 104.615
R1650 VTAIL.n197 VTAIL.n101 104.615
R1651 VTAIL.n232 VTAIL.n229 104.615
R1652 VTAIL.n239 VTAIL.n229 104.615
R1653 VTAIL.n240 VTAIL.n239 104.615
R1654 VTAIL.n240 VTAIL.n225 104.615
R1655 VTAIL.n247 VTAIL.n225 104.615
R1656 VTAIL.n249 VTAIL.n247 104.615
R1657 VTAIL.n249 VTAIL.n248 104.615
R1658 VTAIL.n248 VTAIL.n221 104.615
R1659 VTAIL.n257 VTAIL.n221 104.615
R1660 VTAIL.n258 VTAIL.n257 104.615
R1661 VTAIL.n258 VTAIL.n217 104.615
R1662 VTAIL.n265 VTAIL.n217 104.615
R1663 VTAIL.n266 VTAIL.n265 104.615
R1664 VTAIL.n266 VTAIL.n213 104.615
R1665 VTAIL.n273 VTAIL.n213 104.615
R1666 VTAIL.n274 VTAIL.n273 104.615
R1667 VTAIL.n274 VTAIL.n209 104.615
R1668 VTAIL.n281 VTAIL.n209 104.615
R1669 VTAIL.n282 VTAIL.n281 104.615
R1670 VTAIL.n282 VTAIL.n205 104.615
R1671 VTAIL.n289 VTAIL.n205 104.615
R1672 VTAIL.n290 VTAIL.n289 104.615
R1673 VTAIL.n290 VTAIL.n201 104.615
R1674 VTAIL.n297 VTAIL.n201 104.615
R1675 VTAIL.n697 VTAIL.n601 104.615
R1676 VTAIL.n690 VTAIL.n601 104.615
R1677 VTAIL.n690 VTAIL.n689 104.615
R1678 VTAIL.n689 VTAIL.n605 104.615
R1679 VTAIL.n682 VTAIL.n605 104.615
R1680 VTAIL.n682 VTAIL.n681 104.615
R1681 VTAIL.n681 VTAIL.n609 104.615
R1682 VTAIL.n674 VTAIL.n609 104.615
R1683 VTAIL.n674 VTAIL.n673 104.615
R1684 VTAIL.n673 VTAIL.n613 104.615
R1685 VTAIL.n666 VTAIL.n613 104.615
R1686 VTAIL.n666 VTAIL.n665 104.615
R1687 VTAIL.n665 VTAIL.n617 104.615
R1688 VTAIL.n658 VTAIL.n617 104.615
R1689 VTAIL.n658 VTAIL.n657 104.615
R1690 VTAIL.n657 VTAIL.n621 104.615
R1691 VTAIL.n625 VTAIL.n621 104.615
R1692 VTAIL.n649 VTAIL.n625 104.615
R1693 VTAIL.n649 VTAIL.n648 104.615
R1694 VTAIL.n648 VTAIL.n626 104.615
R1695 VTAIL.n641 VTAIL.n626 104.615
R1696 VTAIL.n641 VTAIL.n640 104.615
R1697 VTAIL.n640 VTAIL.n630 104.615
R1698 VTAIL.n633 VTAIL.n630 104.615
R1699 VTAIL.n597 VTAIL.n501 104.615
R1700 VTAIL.n590 VTAIL.n501 104.615
R1701 VTAIL.n590 VTAIL.n589 104.615
R1702 VTAIL.n589 VTAIL.n505 104.615
R1703 VTAIL.n582 VTAIL.n505 104.615
R1704 VTAIL.n582 VTAIL.n581 104.615
R1705 VTAIL.n581 VTAIL.n509 104.615
R1706 VTAIL.n574 VTAIL.n509 104.615
R1707 VTAIL.n574 VTAIL.n573 104.615
R1708 VTAIL.n573 VTAIL.n513 104.615
R1709 VTAIL.n566 VTAIL.n513 104.615
R1710 VTAIL.n566 VTAIL.n565 104.615
R1711 VTAIL.n565 VTAIL.n517 104.615
R1712 VTAIL.n558 VTAIL.n517 104.615
R1713 VTAIL.n558 VTAIL.n557 104.615
R1714 VTAIL.n557 VTAIL.n521 104.615
R1715 VTAIL.n525 VTAIL.n521 104.615
R1716 VTAIL.n549 VTAIL.n525 104.615
R1717 VTAIL.n549 VTAIL.n548 104.615
R1718 VTAIL.n548 VTAIL.n526 104.615
R1719 VTAIL.n541 VTAIL.n526 104.615
R1720 VTAIL.n541 VTAIL.n540 104.615
R1721 VTAIL.n540 VTAIL.n530 104.615
R1722 VTAIL.n533 VTAIL.n530 104.615
R1723 VTAIL.n497 VTAIL.n401 104.615
R1724 VTAIL.n490 VTAIL.n401 104.615
R1725 VTAIL.n490 VTAIL.n489 104.615
R1726 VTAIL.n489 VTAIL.n405 104.615
R1727 VTAIL.n482 VTAIL.n405 104.615
R1728 VTAIL.n482 VTAIL.n481 104.615
R1729 VTAIL.n481 VTAIL.n409 104.615
R1730 VTAIL.n474 VTAIL.n409 104.615
R1731 VTAIL.n474 VTAIL.n473 104.615
R1732 VTAIL.n473 VTAIL.n413 104.615
R1733 VTAIL.n466 VTAIL.n413 104.615
R1734 VTAIL.n466 VTAIL.n465 104.615
R1735 VTAIL.n465 VTAIL.n417 104.615
R1736 VTAIL.n458 VTAIL.n417 104.615
R1737 VTAIL.n458 VTAIL.n457 104.615
R1738 VTAIL.n457 VTAIL.n421 104.615
R1739 VTAIL.n425 VTAIL.n421 104.615
R1740 VTAIL.n449 VTAIL.n425 104.615
R1741 VTAIL.n449 VTAIL.n448 104.615
R1742 VTAIL.n448 VTAIL.n426 104.615
R1743 VTAIL.n441 VTAIL.n426 104.615
R1744 VTAIL.n441 VTAIL.n440 104.615
R1745 VTAIL.n440 VTAIL.n430 104.615
R1746 VTAIL.n433 VTAIL.n430 104.615
R1747 VTAIL.n397 VTAIL.n301 104.615
R1748 VTAIL.n390 VTAIL.n301 104.615
R1749 VTAIL.n390 VTAIL.n389 104.615
R1750 VTAIL.n389 VTAIL.n305 104.615
R1751 VTAIL.n382 VTAIL.n305 104.615
R1752 VTAIL.n382 VTAIL.n381 104.615
R1753 VTAIL.n381 VTAIL.n309 104.615
R1754 VTAIL.n374 VTAIL.n309 104.615
R1755 VTAIL.n374 VTAIL.n373 104.615
R1756 VTAIL.n373 VTAIL.n313 104.615
R1757 VTAIL.n366 VTAIL.n313 104.615
R1758 VTAIL.n366 VTAIL.n365 104.615
R1759 VTAIL.n365 VTAIL.n317 104.615
R1760 VTAIL.n358 VTAIL.n317 104.615
R1761 VTAIL.n358 VTAIL.n357 104.615
R1762 VTAIL.n357 VTAIL.n321 104.615
R1763 VTAIL.n325 VTAIL.n321 104.615
R1764 VTAIL.n349 VTAIL.n325 104.615
R1765 VTAIL.n349 VTAIL.n348 104.615
R1766 VTAIL.n348 VTAIL.n326 104.615
R1767 VTAIL.n341 VTAIL.n326 104.615
R1768 VTAIL.n341 VTAIL.n340 104.615
R1769 VTAIL.n340 VTAIL.n330 104.615
R1770 VTAIL.n333 VTAIL.n330 104.615
R1771 VTAIL.n732 VTAIL.t1 52.3082
R1772 VTAIL.n32 VTAIL.t2 52.3082
R1773 VTAIL.n132 VTAIL.t7 52.3082
R1774 VTAIL.n232 VTAIL.t4 52.3082
R1775 VTAIL.n633 VTAIL.t5 52.3082
R1776 VTAIL.n533 VTAIL.t6 52.3082
R1777 VTAIL.n433 VTAIL.t3 52.3082
R1778 VTAIL.n333 VTAIL.t0 52.3082
R1779 VTAIL.n799 VTAIL.n798 34.1247
R1780 VTAIL.n99 VTAIL.n98 34.1247
R1781 VTAIL.n199 VTAIL.n198 34.1247
R1782 VTAIL.n299 VTAIL.n298 34.1247
R1783 VTAIL.n699 VTAIL.n698 34.1247
R1784 VTAIL.n599 VTAIL.n598 34.1247
R1785 VTAIL.n499 VTAIL.n498 34.1247
R1786 VTAIL.n399 VTAIL.n398 34.1247
R1787 VTAIL.n799 VTAIL.n699 28.6858
R1788 VTAIL.n399 VTAIL.n299 28.6858
R1789 VTAIL.n756 VTAIL.n755 13.1884
R1790 VTAIL.n56 VTAIL.n55 13.1884
R1791 VTAIL.n156 VTAIL.n155 13.1884
R1792 VTAIL.n256 VTAIL.n255 13.1884
R1793 VTAIL.n656 VTAIL.n655 13.1884
R1794 VTAIL.n556 VTAIL.n555 13.1884
R1795 VTAIL.n456 VTAIL.n455 13.1884
R1796 VTAIL.n356 VTAIL.n355 13.1884
R1797 VTAIL.n754 VTAIL.n722 12.8005
R1798 VTAIL.n759 VTAIL.n720 12.8005
R1799 VTAIL.n54 VTAIL.n22 12.8005
R1800 VTAIL.n59 VTAIL.n20 12.8005
R1801 VTAIL.n154 VTAIL.n122 12.8005
R1802 VTAIL.n159 VTAIL.n120 12.8005
R1803 VTAIL.n254 VTAIL.n222 12.8005
R1804 VTAIL.n259 VTAIL.n220 12.8005
R1805 VTAIL.n659 VTAIL.n620 12.8005
R1806 VTAIL.n654 VTAIL.n622 12.8005
R1807 VTAIL.n559 VTAIL.n520 12.8005
R1808 VTAIL.n554 VTAIL.n522 12.8005
R1809 VTAIL.n459 VTAIL.n420 12.8005
R1810 VTAIL.n454 VTAIL.n422 12.8005
R1811 VTAIL.n359 VTAIL.n320 12.8005
R1812 VTAIL.n354 VTAIL.n322 12.8005
R1813 VTAIL.n751 VTAIL.n750 12.0247
R1814 VTAIL.n760 VTAIL.n718 12.0247
R1815 VTAIL.n796 VTAIL.n700 12.0247
R1816 VTAIL.n51 VTAIL.n50 12.0247
R1817 VTAIL.n60 VTAIL.n18 12.0247
R1818 VTAIL.n96 VTAIL.n0 12.0247
R1819 VTAIL.n151 VTAIL.n150 12.0247
R1820 VTAIL.n160 VTAIL.n118 12.0247
R1821 VTAIL.n196 VTAIL.n100 12.0247
R1822 VTAIL.n251 VTAIL.n250 12.0247
R1823 VTAIL.n260 VTAIL.n218 12.0247
R1824 VTAIL.n296 VTAIL.n200 12.0247
R1825 VTAIL.n696 VTAIL.n600 12.0247
R1826 VTAIL.n660 VTAIL.n618 12.0247
R1827 VTAIL.n651 VTAIL.n650 12.0247
R1828 VTAIL.n596 VTAIL.n500 12.0247
R1829 VTAIL.n560 VTAIL.n518 12.0247
R1830 VTAIL.n551 VTAIL.n550 12.0247
R1831 VTAIL.n496 VTAIL.n400 12.0247
R1832 VTAIL.n460 VTAIL.n418 12.0247
R1833 VTAIL.n451 VTAIL.n450 12.0247
R1834 VTAIL.n396 VTAIL.n300 12.0247
R1835 VTAIL.n360 VTAIL.n318 12.0247
R1836 VTAIL.n351 VTAIL.n350 12.0247
R1837 VTAIL.n746 VTAIL.n724 11.249
R1838 VTAIL.n764 VTAIL.n763 11.249
R1839 VTAIL.n795 VTAIL.n702 11.249
R1840 VTAIL.n46 VTAIL.n24 11.249
R1841 VTAIL.n64 VTAIL.n63 11.249
R1842 VTAIL.n95 VTAIL.n2 11.249
R1843 VTAIL.n146 VTAIL.n124 11.249
R1844 VTAIL.n164 VTAIL.n163 11.249
R1845 VTAIL.n195 VTAIL.n102 11.249
R1846 VTAIL.n246 VTAIL.n224 11.249
R1847 VTAIL.n264 VTAIL.n263 11.249
R1848 VTAIL.n295 VTAIL.n202 11.249
R1849 VTAIL.n695 VTAIL.n602 11.249
R1850 VTAIL.n664 VTAIL.n663 11.249
R1851 VTAIL.n647 VTAIL.n624 11.249
R1852 VTAIL.n595 VTAIL.n502 11.249
R1853 VTAIL.n564 VTAIL.n563 11.249
R1854 VTAIL.n547 VTAIL.n524 11.249
R1855 VTAIL.n495 VTAIL.n402 11.249
R1856 VTAIL.n464 VTAIL.n463 11.249
R1857 VTAIL.n447 VTAIL.n424 11.249
R1858 VTAIL.n395 VTAIL.n302 11.249
R1859 VTAIL.n364 VTAIL.n363 11.249
R1860 VTAIL.n347 VTAIL.n324 11.249
R1861 VTAIL.n745 VTAIL.n726 10.4732
R1862 VTAIL.n767 VTAIL.n716 10.4732
R1863 VTAIL.n792 VTAIL.n791 10.4732
R1864 VTAIL.n45 VTAIL.n26 10.4732
R1865 VTAIL.n67 VTAIL.n16 10.4732
R1866 VTAIL.n92 VTAIL.n91 10.4732
R1867 VTAIL.n145 VTAIL.n126 10.4732
R1868 VTAIL.n167 VTAIL.n116 10.4732
R1869 VTAIL.n192 VTAIL.n191 10.4732
R1870 VTAIL.n245 VTAIL.n226 10.4732
R1871 VTAIL.n267 VTAIL.n216 10.4732
R1872 VTAIL.n292 VTAIL.n291 10.4732
R1873 VTAIL.n692 VTAIL.n691 10.4732
R1874 VTAIL.n667 VTAIL.n616 10.4732
R1875 VTAIL.n646 VTAIL.n627 10.4732
R1876 VTAIL.n592 VTAIL.n591 10.4732
R1877 VTAIL.n567 VTAIL.n516 10.4732
R1878 VTAIL.n546 VTAIL.n527 10.4732
R1879 VTAIL.n492 VTAIL.n491 10.4732
R1880 VTAIL.n467 VTAIL.n416 10.4732
R1881 VTAIL.n446 VTAIL.n427 10.4732
R1882 VTAIL.n392 VTAIL.n391 10.4732
R1883 VTAIL.n367 VTAIL.n316 10.4732
R1884 VTAIL.n346 VTAIL.n327 10.4732
R1885 VTAIL.n733 VTAIL.n731 10.2747
R1886 VTAIL.n33 VTAIL.n31 10.2747
R1887 VTAIL.n133 VTAIL.n131 10.2747
R1888 VTAIL.n233 VTAIL.n231 10.2747
R1889 VTAIL.n634 VTAIL.n632 10.2747
R1890 VTAIL.n534 VTAIL.n532 10.2747
R1891 VTAIL.n434 VTAIL.n432 10.2747
R1892 VTAIL.n334 VTAIL.n332 10.2747
R1893 VTAIL.n742 VTAIL.n741 9.69747
R1894 VTAIL.n768 VTAIL.n714 9.69747
R1895 VTAIL.n788 VTAIL.n704 9.69747
R1896 VTAIL.n42 VTAIL.n41 9.69747
R1897 VTAIL.n68 VTAIL.n14 9.69747
R1898 VTAIL.n88 VTAIL.n4 9.69747
R1899 VTAIL.n142 VTAIL.n141 9.69747
R1900 VTAIL.n168 VTAIL.n114 9.69747
R1901 VTAIL.n188 VTAIL.n104 9.69747
R1902 VTAIL.n242 VTAIL.n241 9.69747
R1903 VTAIL.n268 VTAIL.n214 9.69747
R1904 VTAIL.n288 VTAIL.n204 9.69747
R1905 VTAIL.n688 VTAIL.n604 9.69747
R1906 VTAIL.n668 VTAIL.n614 9.69747
R1907 VTAIL.n643 VTAIL.n642 9.69747
R1908 VTAIL.n588 VTAIL.n504 9.69747
R1909 VTAIL.n568 VTAIL.n514 9.69747
R1910 VTAIL.n543 VTAIL.n542 9.69747
R1911 VTAIL.n488 VTAIL.n404 9.69747
R1912 VTAIL.n468 VTAIL.n414 9.69747
R1913 VTAIL.n443 VTAIL.n442 9.69747
R1914 VTAIL.n388 VTAIL.n304 9.69747
R1915 VTAIL.n368 VTAIL.n314 9.69747
R1916 VTAIL.n343 VTAIL.n342 9.69747
R1917 VTAIL.n794 VTAIL.n700 9.45567
R1918 VTAIL.n94 VTAIL.n0 9.45567
R1919 VTAIL.n194 VTAIL.n100 9.45567
R1920 VTAIL.n294 VTAIL.n200 9.45567
R1921 VTAIL.n694 VTAIL.n600 9.45567
R1922 VTAIL.n594 VTAIL.n500 9.45567
R1923 VTAIL.n494 VTAIL.n400 9.45567
R1924 VTAIL.n394 VTAIL.n300 9.45567
R1925 VTAIL.n779 VTAIL.n778 9.3005
R1926 VTAIL.n708 VTAIL.n707 9.3005
R1927 VTAIL.n785 VTAIL.n784 9.3005
R1928 VTAIL.n787 VTAIL.n786 9.3005
R1929 VTAIL.n704 VTAIL.n703 9.3005
R1930 VTAIL.n793 VTAIL.n792 9.3005
R1931 VTAIL.n795 VTAIL.n794 9.3005
R1932 VTAIL.n712 VTAIL.n711 9.3005
R1933 VTAIL.n771 VTAIL.n770 9.3005
R1934 VTAIL.n769 VTAIL.n768 9.3005
R1935 VTAIL.n716 VTAIL.n715 9.3005
R1936 VTAIL.n763 VTAIL.n762 9.3005
R1937 VTAIL.n761 VTAIL.n760 9.3005
R1938 VTAIL.n720 VTAIL.n719 9.3005
R1939 VTAIL.n735 VTAIL.n734 9.3005
R1940 VTAIL.n737 VTAIL.n736 9.3005
R1941 VTAIL.n728 VTAIL.n727 9.3005
R1942 VTAIL.n743 VTAIL.n742 9.3005
R1943 VTAIL.n745 VTAIL.n744 9.3005
R1944 VTAIL.n724 VTAIL.n723 9.3005
R1945 VTAIL.n752 VTAIL.n751 9.3005
R1946 VTAIL.n754 VTAIL.n753 9.3005
R1947 VTAIL.n777 VTAIL.n776 9.3005
R1948 VTAIL.n79 VTAIL.n78 9.3005
R1949 VTAIL.n8 VTAIL.n7 9.3005
R1950 VTAIL.n85 VTAIL.n84 9.3005
R1951 VTAIL.n87 VTAIL.n86 9.3005
R1952 VTAIL.n4 VTAIL.n3 9.3005
R1953 VTAIL.n93 VTAIL.n92 9.3005
R1954 VTAIL.n95 VTAIL.n94 9.3005
R1955 VTAIL.n12 VTAIL.n11 9.3005
R1956 VTAIL.n71 VTAIL.n70 9.3005
R1957 VTAIL.n69 VTAIL.n68 9.3005
R1958 VTAIL.n16 VTAIL.n15 9.3005
R1959 VTAIL.n63 VTAIL.n62 9.3005
R1960 VTAIL.n61 VTAIL.n60 9.3005
R1961 VTAIL.n20 VTAIL.n19 9.3005
R1962 VTAIL.n35 VTAIL.n34 9.3005
R1963 VTAIL.n37 VTAIL.n36 9.3005
R1964 VTAIL.n28 VTAIL.n27 9.3005
R1965 VTAIL.n43 VTAIL.n42 9.3005
R1966 VTAIL.n45 VTAIL.n44 9.3005
R1967 VTAIL.n24 VTAIL.n23 9.3005
R1968 VTAIL.n52 VTAIL.n51 9.3005
R1969 VTAIL.n54 VTAIL.n53 9.3005
R1970 VTAIL.n77 VTAIL.n76 9.3005
R1971 VTAIL.n179 VTAIL.n178 9.3005
R1972 VTAIL.n108 VTAIL.n107 9.3005
R1973 VTAIL.n185 VTAIL.n184 9.3005
R1974 VTAIL.n187 VTAIL.n186 9.3005
R1975 VTAIL.n104 VTAIL.n103 9.3005
R1976 VTAIL.n193 VTAIL.n192 9.3005
R1977 VTAIL.n195 VTAIL.n194 9.3005
R1978 VTAIL.n112 VTAIL.n111 9.3005
R1979 VTAIL.n171 VTAIL.n170 9.3005
R1980 VTAIL.n169 VTAIL.n168 9.3005
R1981 VTAIL.n116 VTAIL.n115 9.3005
R1982 VTAIL.n163 VTAIL.n162 9.3005
R1983 VTAIL.n161 VTAIL.n160 9.3005
R1984 VTAIL.n120 VTAIL.n119 9.3005
R1985 VTAIL.n135 VTAIL.n134 9.3005
R1986 VTAIL.n137 VTAIL.n136 9.3005
R1987 VTAIL.n128 VTAIL.n127 9.3005
R1988 VTAIL.n143 VTAIL.n142 9.3005
R1989 VTAIL.n145 VTAIL.n144 9.3005
R1990 VTAIL.n124 VTAIL.n123 9.3005
R1991 VTAIL.n152 VTAIL.n151 9.3005
R1992 VTAIL.n154 VTAIL.n153 9.3005
R1993 VTAIL.n177 VTAIL.n176 9.3005
R1994 VTAIL.n279 VTAIL.n278 9.3005
R1995 VTAIL.n208 VTAIL.n207 9.3005
R1996 VTAIL.n285 VTAIL.n284 9.3005
R1997 VTAIL.n287 VTAIL.n286 9.3005
R1998 VTAIL.n204 VTAIL.n203 9.3005
R1999 VTAIL.n293 VTAIL.n292 9.3005
R2000 VTAIL.n295 VTAIL.n294 9.3005
R2001 VTAIL.n212 VTAIL.n211 9.3005
R2002 VTAIL.n271 VTAIL.n270 9.3005
R2003 VTAIL.n269 VTAIL.n268 9.3005
R2004 VTAIL.n216 VTAIL.n215 9.3005
R2005 VTAIL.n263 VTAIL.n262 9.3005
R2006 VTAIL.n261 VTAIL.n260 9.3005
R2007 VTAIL.n220 VTAIL.n219 9.3005
R2008 VTAIL.n235 VTAIL.n234 9.3005
R2009 VTAIL.n237 VTAIL.n236 9.3005
R2010 VTAIL.n228 VTAIL.n227 9.3005
R2011 VTAIL.n243 VTAIL.n242 9.3005
R2012 VTAIL.n245 VTAIL.n244 9.3005
R2013 VTAIL.n224 VTAIL.n223 9.3005
R2014 VTAIL.n252 VTAIL.n251 9.3005
R2015 VTAIL.n254 VTAIL.n253 9.3005
R2016 VTAIL.n277 VTAIL.n276 9.3005
R2017 VTAIL.n695 VTAIL.n694 9.3005
R2018 VTAIL.n693 VTAIL.n692 9.3005
R2019 VTAIL.n604 VTAIL.n603 9.3005
R2020 VTAIL.n687 VTAIL.n686 9.3005
R2021 VTAIL.n685 VTAIL.n684 9.3005
R2022 VTAIL.n608 VTAIL.n607 9.3005
R2023 VTAIL.n679 VTAIL.n678 9.3005
R2024 VTAIL.n677 VTAIL.n676 9.3005
R2025 VTAIL.n612 VTAIL.n611 9.3005
R2026 VTAIL.n671 VTAIL.n670 9.3005
R2027 VTAIL.n669 VTAIL.n668 9.3005
R2028 VTAIL.n616 VTAIL.n615 9.3005
R2029 VTAIL.n663 VTAIL.n662 9.3005
R2030 VTAIL.n661 VTAIL.n660 9.3005
R2031 VTAIL.n620 VTAIL.n619 9.3005
R2032 VTAIL.n654 VTAIL.n653 9.3005
R2033 VTAIL.n652 VTAIL.n651 9.3005
R2034 VTAIL.n624 VTAIL.n623 9.3005
R2035 VTAIL.n646 VTAIL.n645 9.3005
R2036 VTAIL.n644 VTAIL.n643 9.3005
R2037 VTAIL.n629 VTAIL.n628 9.3005
R2038 VTAIL.n638 VTAIL.n637 9.3005
R2039 VTAIL.n636 VTAIL.n635 9.3005
R2040 VTAIL.n536 VTAIL.n535 9.3005
R2041 VTAIL.n538 VTAIL.n537 9.3005
R2042 VTAIL.n529 VTAIL.n528 9.3005
R2043 VTAIL.n544 VTAIL.n543 9.3005
R2044 VTAIL.n546 VTAIL.n545 9.3005
R2045 VTAIL.n524 VTAIL.n523 9.3005
R2046 VTAIL.n552 VTAIL.n551 9.3005
R2047 VTAIL.n554 VTAIL.n553 9.3005
R2048 VTAIL.n508 VTAIL.n507 9.3005
R2049 VTAIL.n585 VTAIL.n584 9.3005
R2050 VTAIL.n587 VTAIL.n586 9.3005
R2051 VTAIL.n504 VTAIL.n503 9.3005
R2052 VTAIL.n593 VTAIL.n592 9.3005
R2053 VTAIL.n595 VTAIL.n594 9.3005
R2054 VTAIL.n579 VTAIL.n578 9.3005
R2055 VTAIL.n577 VTAIL.n576 9.3005
R2056 VTAIL.n512 VTAIL.n511 9.3005
R2057 VTAIL.n571 VTAIL.n570 9.3005
R2058 VTAIL.n569 VTAIL.n568 9.3005
R2059 VTAIL.n516 VTAIL.n515 9.3005
R2060 VTAIL.n563 VTAIL.n562 9.3005
R2061 VTAIL.n561 VTAIL.n560 9.3005
R2062 VTAIL.n520 VTAIL.n519 9.3005
R2063 VTAIL.n436 VTAIL.n435 9.3005
R2064 VTAIL.n438 VTAIL.n437 9.3005
R2065 VTAIL.n429 VTAIL.n428 9.3005
R2066 VTAIL.n444 VTAIL.n443 9.3005
R2067 VTAIL.n446 VTAIL.n445 9.3005
R2068 VTAIL.n424 VTAIL.n423 9.3005
R2069 VTAIL.n452 VTAIL.n451 9.3005
R2070 VTAIL.n454 VTAIL.n453 9.3005
R2071 VTAIL.n408 VTAIL.n407 9.3005
R2072 VTAIL.n485 VTAIL.n484 9.3005
R2073 VTAIL.n487 VTAIL.n486 9.3005
R2074 VTAIL.n404 VTAIL.n403 9.3005
R2075 VTAIL.n493 VTAIL.n492 9.3005
R2076 VTAIL.n495 VTAIL.n494 9.3005
R2077 VTAIL.n479 VTAIL.n478 9.3005
R2078 VTAIL.n477 VTAIL.n476 9.3005
R2079 VTAIL.n412 VTAIL.n411 9.3005
R2080 VTAIL.n471 VTAIL.n470 9.3005
R2081 VTAIL.n469 VTAIL.n468 9.3005
R2082 VTAIL.n416 VTAIL.n415 9.3005
R2083 VTAIL.n463 VTAIL.n462 9.3005
R2084 VTAIL.n461 VTAIL.n460 9.3005
R2085 VTAIL.n420 VTAIL.n419 9.3005
R2086 VTAIL.n336 VTAIL.n335 9.3005
R2087 VTAIL.n338 VTAIL.n337 9.3005
R2088 VTAIL.n329 VTAIL.n328 9.3005
R2089 VTAIL.n344 VTAIL.n343 9.3005
R2090 VTAIL.n346 VTAIL.n345 9.3005
R2091 VTAIL.n324 VTAIL.n323 9.3005
R2092 VTAIL.n352 VTAIL.n351 9.3005
R2093 VTAIL.n354 VTAIL.n353 9.3005
R2094 VTAIL.n308 VTAIL.n307 9.3005
R2095 VTAIL.n385 VTAIL.n384 9.3005
R2096 VTAIL.n387 VTAIL.n386 9.3005
R2097 VTAIL.n304 VTAIL.n303 9.3005
R2098 VTAIL.n393 VTAIL.n392 9.3005
R2099 VTAIL.n395 VTAIL.n394 9.3005
R2100 VTAIL.n379 VTAIL.n378 9.3005
R2101 VTAIL.n377 VTAIL.n376 9.3005
R2102 VTAIL.n312 VTAIL.n311 9.3005
R2103 VTAIL.n371 VTAIL.n370 9.3005
R2104 VTAIL.n369 VTAIL.n368 9.3005
R2105 VTAIL.n316 VTAIL.n315 9.3005
R2106 VTAIL.n363 VTAIL.n362 9.3005
R2107 VTAIL.n361 VTAIL.n360 9.3005
R2108 VTAIL.n320 VTAIL.n319 9.3005
R2109 VTAIL.n738 VTAIL.n728 8.92171
R2110 VTAIL.n772 VTAIL.n771 8.92171
R2111 VTAIL.n787 VTAIL.n706 8.92171
R2112 VTAIL.n38 VTAIL.n28 8.92171
R2113 VTAIL.n72 VTAIL.n71 8.92171
R2114 VTAIL.n87 VTAIL.n6 8.92171
R2115 VTAIL.n138 VTAIL.n128 8.92171
R2116 VTAIL.n172 VTAIL.n171 8.92171
R2117 VTAIL.n187 VTAIL.n106 8.92171
R2118 VTAIL.n238 VTAIL.n228 8.92171
R2119 VTAIL.n272 VTAIL.n271 8.92171
R2120 VTAIL.n287 VTAIL.n206 8.92171
R2121 VTAIL.n687 VTAIL.n606 8.92171
R2122 VTAIL.n672 VTAIL.n671 8.92171
R2123 VTAIL.n639 VTAIL.n629 8.92171
R2124 VTAIL.n587 VTAIL.n506 8.92171
R2125 VTAIL.n572 VTAIL.n571 8.92171
R2126 VTAIL.n539 VTAIL.n529 8.92171
R2127 VTAIL.n487 VTAIL.n406 8.92171
R2128 VTAIL.n472 VTAIL.n471 8.92171
R2129 VTAIL.n439 VTAIL.n429 8.92171
R2130 VTAIL.n387 VTAIL.n306 8.92171
R2131 VTAIL.n372 VTAIL.n371 8.92171
R2132 VTAIL.n339 VTAIL.n329 8.92171
R2133 VTAIL.n737 VTAIL.n730 8.14595
R2134 VTAIL.n775 VTAIL.n712 8.14595
R2135 VTAIL.n784 VTAIL.n783 8.14595
R2136 VTAIL.n37 VTAIL.n30 8.14595
R2137 VTAIL.n75 VTAIL.n12 8.14595
R2138 VTAIL.n84 VTAIL.n83 8.14595
R2139 VTAIL.n137 VTAIL.n130 8.14595
R2140 VTAIL.n175 VTAIL.n112 8.14595
R2141 VTAIL.n184 VTAIL.n183 8.14595
R2142 VTAIL.n237 VTAIL.n230 8.14595
R2143 VTAIL.n275 VTAIL.n212 8.14595
R2144 VTAIL.n284 VTAIL.n283 8.14595
R2145 VTAIL.n684 VTAIL.n683 8.14595
R2146 VTAIL.n675 VTAIL.n612 8.14595
R2147 VTAIL.n638 VTAIL.n631 8.14595
R2148 VTAIL.n584 VTAIL.n583 8.14595
R2149 VTAIL.n575 VTAIL.n512 8.14595
R2150 VTAIL.n538 VTAIL.n531 8.14595
R2151 VTAIL.n484 VTAIL.n483 8.14595
R2152 VTAIL.n475 VTAIL.n412 8.14595
R2153 VTAIL.n438 VTAIL.n431 8.14595
R2154 VTAIL.n384 VTAIL.n383 8.14595
R2155 VTAIL.n375 VTAIL.n312 8.14595
R2156 VTAIL.n338 VTAIL.n331 8.14595
R2157 VTAIL.n734 VTAIL.n733 7.3702
R2158 VTAIL.n776 VTAIL.n710 7.3702
R2159 VTAIL.n780 VTAIL.n708 7.3702
R2160 VTAIL.n34 VTAIL.n33 7.3702
R2161 VTAIL.n76 VTAIL.n10 7.3702
R2162 VTAIL.n80 VTAIL.n8 7.3702
R2163 VTAIL.n134 VTAIL.n133 7.3702
R2164 VTAIL.n176 VTAIL.n110 7.3702
R2165 VTAIL.n180 VTAIL.n108 7.3702
R2166 VTAIL.n234 VTAIL.n233 7.3702
R2167 VTAIL.n276 VTAIL.n210 7.3702
R2168 VTAIL.n280 VTAIL.n208 7.3702
R2169 VTAIL.n680 VTAIL.n608 7.3702
R2170 VTAIL.n676 VTAIL.n610 7.3702
R2171 VTAIL.n635 VTAIL.n634 7.3702
R2172 VTAIL.n580 VTAIL.n508 7.3702
R2173 VTAIL.n576 VTAIL.n510 7.3702
R2174 VTAIL.n535 VTAIL.n534 7.3702
R2175 VTAIL.n480 VTAIL.n408 7.3702
R2176 VTAIL.n476 VTAIL.n410 7.3702
R2177 VTAIL.n435 VTAIL.n434 7.3702
R2178 VTAIL.n380 VTAIL.n308 7.3702
R2179 VTAIL.n376 VTAIL.n310 7.3702
R2180 VTAIL.n335 VTAIL.n334 7.3702
R2181 VTAIL.n779 VTAIL.n710 6.59444
R2182 VTAIL.n780 VTAIL.n779 6.59444
R2183 VTAIL.n79 VTAIL.n10 6.59444
R2184 VTAIL.n80 VTAIL.n79 6.59444
R2185 VTAIL.n179 VTAIL.n110 6.59444
R2186 VTAIL.n180 VTAIL.n179 6.59444
R2187 VTAIL.n279 VTAIL.n210 6.59444
R2188 VTAIL.n280 VTAIL.n279 6.59444
R2189 VTAIL.n680 VTAIL.n679 6.59444
R2190 VTAIL.n679 VTAIL.n610 6.59444
R2191 VTAIL.n580 VTAIL.n579 6.59444
R2192 VTAIL.n579 VTAIL.n510 6.59444
R2193 VTAIL.n480 VTAIL.n479 6.59444
R2194 VTAIL.n479 VTAIL.n410 6.59444
R2195 VTAIL.n380 VTAIL.n379 6.59444
R2196 VTAIL.n379 VTAIL.n310 6.59444
R2197 VTAIL.n734 VTAIL.n730 5.81868
R2198 VTAIL.n776 VTAIL.n775 5.81868
R2199 VTAIL.n783 VTAIL.n708 5.81868
R2200 VTAIL.n34 VTAIL.n30 5.81868
R2201 VTAIL.n76 VTAIL.n75 5.81868
R2202 VTAIL.n83 VTAIL.n8 5.81868
R2203 VTAIL.n134 VTAIL.n130 5.81868
R2204 VTAIL.n176 VTAIL.n175 5.81868
R2205 VTAIL.n183 VTAIL.n108 5.81868
R2206 VTAIL.n234 VTAIL.n230 5.81868
R2207 VTAIL.n276 VTAIL.n275 5.81868
R2208 VTAIL.n283 VTAIL.n208 5.81868
R2209 VTAIL.n683 VTAIL.n608 5.81868
R2210 VTAIL.n676 VTAIL.n675 5.81868
R2211 VTAIL.n635 VTAIL.n631 5.81868
R2212 VTAIL.n583 VTAIL.n508 5.81868
R2213 VTAIL.n576 VTAIL.n575 5.81868
R2214 VTAIL.n535 VTAIL.n531 5.81868
R2215 VTAIL.n483 VTAIL.n408 5.81868
R2216 VTAIL.n476 VTAIL.n475 5.81868
R2217 VTAIL.n435 VTAIL.n431 5.81868
R2218 VTAIL.n383 VTAIL.n308 5.81868
R2219 VTAIL.n376 VTAIL.n375 5.81868
R2220 VTAIL.n335 VTAIL.n331 5.81868
R2221 VTAIL.n738 VTAIL.n737 5.04292
R2222 VTAIL.n772 VTAIL.n712 5.04292
R2223 VTAIL.n784 VTAIL.n706 5.04292
R2224 VTAIL.n38 VTAIL.n37 5.04292
R2225 VTAIL.n72 VTAIL.n12 5.04292
R2226 VTAIL.n84 VTAIL.n6 5.04292
R2227 VTAIL.n138 VTAIL.n137 5.04292
R2228 VTAIL.n172 VTAIL.n112 5.04292
R2229 VTAIL.n184 VTAIL.n106 5.04292
R2230 VTAIL.n238 VTAIL.n237 5.04292
R2231 VTAIL.n272 VTAIL.n212 5.04292
R2232 VTAIL.n284 VTAIL.n206 5.04292
R2233 VTAIL.n684 VTAIL.n606 5.04292
R2234 VTAIL.n672 VTAIL.n612 5.04292
R2235 VTAIL.n639 VTAIL.n638 5.04292
R2236 VTAIL.n584 VTAIL.n506 5.04292
R2237 VTAIL.n572 VTAIL.n512 5.04292
R2238 VTAIL.n539 VTAIL.n538 5.04292
R2239 VTAIL.n484 VTAIL.n406 5.04292
R2240 VTAIL.n472 VTAIL.n412 5.04292
R2241 VTAIL.n439 VTAIL.n438 5.04292
R2242 VTAIL.n384 VTAIL.n306 5.04292
R2243 VTAIL.n372 VTAIL.n312 5.04292
R2244 VTAIL.n339 VTAIL.n338 5.04292
R2245 VTAIL.n741 VTAIL.n728 4.26717
R2246 VTAIL.n771 VTAIL.n714 4.26717
R2247 VTAIL.n788 VTAIL.n787 4.26717
R2248 VTAIL.n41 VTAIL.n28 4.26717
R2249 VTAIL.n71 VTAIL.n14 4.26717
R2250 VTAIL.n88 VTAIL.n87 4.26717
R2251 VTAIL.n141 VTAIL.n128 4.26717
R2252 VTAIL.n171 VTAIL.n114 4.26717
R2253 VTAIL.n188 VTAIL.n187 4.26717
R2254 VTAIL.n241 VTAIL.n228 4.26717
R2255 VTAIL.n271 VTAIL.n214 4.26717
R2256 VTAIL.n288 VTAIL.n287 4.26717
R2257 VTAIL.n688 VTAIL.n687 4.26717
R2258 VTAIL.n671 VTAIL.n614 4.26717
R2259 VTAIL.n642 VTAIL.n629 4.26717
R2260 VTAIL.n588 VTAIL.n587 4.26717
R2261 VTAIL.n571 VTAIL.n514 4.26717
R2262 VTAIL.n542 VTAIL.n529 4.26717
R2263 VTAIL.n488 VTAIL.n487 4.26717
R2264 VTAIL.n471 VTAIL.n414 4.26717
R2265 VTAIL.n442 VTAIL.n429 4.26717
R2266 VTAIL.n388 VTAIL.n387 4.26717
R2267 VTAIL.n371 VTAIL.n314 4.26717
R2268 VTAIL.n342 VTAIL.n329 4.26717
R2269 VTAIL.n742 VTAIL.n726 3.49141
R2270 VTAIL.n768 VTAIL.n767 3.49141
R2271 VTAIL.n791 VTAIL.n704 3.49141
R2272 VTAIL.n42 VTAIL.n26 3.49141
R2273 VTAIL.n68 VTAIL.n67 3.49141
R2274 VTAIL.n91 VTAIL.n4 3.49141
R2275 VTAIL.n142 VTAIL.n126 3.49141
R2276 VTAIL.n168 VTAIL.n167 3.49141
R2277 VTAIL.n191 VTAIL.n104 3.49141
R2278 VTAIL.n242 VTAIL.n226 3.49141
R2279 VTAIL.n268 VTAIL.n267 3.49141
R2280 VTAIL.n291 VTAIL.n204 3.49141
R2281 VTAIL.n691 VTAIL.n604 3.49141
R2282 VTAIL.n668 VTAIL.n667 3.49141
R2283 VTAIL.n643 VTAIL.n627 3.49141
R2284 VTAIL.n591 VTAIL.n504 3.49141
R2285 VTAIL.n568 VTAIL.n567 3.49141
R2286 VTAIL.n543 VTAIL.n527 3.49141
R2287 VTAIL.n491 VTAIL.n404 3.49141
R2288 VTAIL.n468 VTAIL.n467 3.49141
R2289 VTAIL.n443 VTAIL.n427 3.49141
R2290 VTAIL.n391 VTAIL.n304 3.49141
R2291 VTAIL.n368 VTAIL.n367 3.49141
R2292 VTAIL.n343 VTAIL.n327 3.49141
R2293 VTAIL.n536 VTAIL.n532 2.84303
R2294 VTAIL.n436 VTAIL.n432 2.84303
R2295 VTAIL.n336 VTAIL.n332 2.84303
R2296 VTAIL.n735 VTAIL.n731 2.84303
R2297 VTAIL.n35 VTAIL.n31 2.84303
R2298 VTAIL.n135 VTAIL.n131 2.84303
R2299 VTAIL.n235 VTAIL.n231 2.84303
R2300 VTAIL.n636 VTAIL.n632 2.84303
R2301 VTAIL.n746 VTAIL.n745 2.71565
R2302 VTAIL.n764 VTAIL.n716 2.71565
R2303 VTAIL.n792 VTAIL.n702 2.71565
R2304 VTAIL.n46 VTAIL.n45 2.71565
R2305 VTAIL.n64 VTAIL.n16 2.71565
R2306 VTAIL.n92 VTAIL.n2 2.71565
R2307 VTAIL.n146 VTAIL.n145 2.71565
R2308 VTAIL.n164 VTAIL.n116 2.71565
R2309 VTAIL.n192 VTAIL.n102 2.71565
R2310 VTAIL.n246 VTAIL.n245 2.71565
R2311 VTAIL.n264 VTAIL.n216 2.71565
R2312 VTAIL.n292 VTAIL.n202 2.71565
R2313 VTAIL.n692 VTAIL.n602 2.71565
R2314 VTAIL.n664 VTAIL.n616 2.71565
R2315 VTAIL.n647 VTAIL.n646 2.71565
R2316 VTAIL.n592 VTAIL.n502 2.71565
R2317 VTAIL.n564 VTAIL.n516 2.71565
R2318 VTAIL.n547 VTAIL.n546 2.71565
R2319 VTAIL.n492 VTAIL.n402 2.71565
R2320 VTAIL.n464 VTAIL.n416 2.71565
R2321 VTAIL.n447 VTAIL.n446 2.71565
R2322 VTAIL.n392 VTAIL.n302 2.71565
R2323 VTAIL.n364 VTAIL.n316 2.71565
R2324 VTAIL.n347 VTAIL.n346 2.71565
R2325 VTAIL.n750 VTAIL.n724 1.93989
R2326 VTAIL.n763 VTAIL.n718 1.93989
R2327 VTAIL.n796 VTAIL.n795 1.93989
R2328 VTAIL.n50 VTAIL.n24 1.93989
R2329 VTAIL.n63 VTAIL.n18 1.93989
R2330 VTAIL.n96 VTAIL.n95 1.93989
R2331 VTAIL.n150 VTAIL.n124 1.93989
R2332 VTAIL.n163 VTAIL.n118 1.93989
R2333 VTAIL.n196 VTAIL.n195 1.93989
R2334 VTAIL.n250 VTAIL.n224 1.93989
R2335 VTAIL.n263 VTAIL.n218 1.93989
R2336 VTAIL.n296 VTAIL.n295 1.93989
R2337 VTAIL.n696 VTAIL.n695 1.93989
R2338 VTAIL.n663 VTAIL.n618 1.93989
R2339 VTAIL.n650 VTAIL.n624 1.93989
R2340 VTAIL.n596 VTAIL.n595 1.93989
R2341 VTAIL.n563 VTAIL.n518 1.93989
R2342 VTAIL.n550 VTAIL.n524 1.93989
R2343 VTAIL.n496 VTAIL.n495 1.93989
R2344 VTAIL.n463 VTAIL.n418 1.93989
R2345 VTAIL.n450 VTAIL.n424 1.93989
R2346 VTAIL.n396 VTAIL.n395 1.93989
R2347 VTAIL.n363 VTAIL.n318 1.93989
R2348 VTAIL.n350 VTAIL.n324 1.93989
R2349 VTAIL.n751 VTAIL.n722 1.16414
R2350 VTAIL.n760 VTAIL.n759 1.16414
R2351 VTAIL.n798 VTAIL.n700 1.16414
R2352 VTAIL.n51 VTAIL.n22 1.16414
R2353 VTAIL.n60 VTAIL.n59 1.16414
R2354 VTAIL.n98 VTAIL.n0 1.16414
R2355 VTAIL.n151 VTAIL.n122 1.16414
R2356 VTAIL.n160 VTAIL.n159 1.16414
R2357 VTAIL.n198 VTAIL.n100 1.16414
R2358 VTAIL.n251 VTAIL.n222 1.16414
R2359 VTAIL.n260 VTAIL.n259 1.16414
R2360 VTAIL.n298 VTAIL.n200 1.16414
R2361 VTAIL.n698 VTAIL.n600 1.16414
R2362 VTAIL.n660 VTAIL.n659 1.16414
R2363 VTAIL.n651 VTAIL.n622 1.16414
R2364 VTAIL.n598 VTAIL.n500 1.16414
R2365 VTAIL.n560 VTAIL.n559 1.16414
R2366 VTAIL.n551 VTAIL.n522 1.16414
R2367 VTAIL.n498 VTAIL.n400 1.16414
R2368 VTAIL.n460 VTAIL.n459 1.16414
R2369 VTAIL.n451 VTAIL.n422 1.16414
R2370 VTAIL.n398 VTAIL.n300 1.16414
R2371 VTAIL.n360 VTAIL.n359 1.16414
R2372 VTAIL.n351 VTAIL.n322 1.16414
R2373 VTAIL.n499 VTAIL.n399 0.767741
R2374 VTAIL.n699 VTAIL.n599 0.767741
R2375 VTAIL.n299 VTAIL.n199 0.767741
R2376 VTAIL.n599 VTAIL.n499 0.470328
R2377 VTAIL.n199 VTAIL.n99 0.470328
R2378 VTAIL VTAIL.n99 0.44231
R2379 VTAIL.n755 VTAIL.n754 0.388379
R2380 VTAIL.n756 VTAIL.n720 0.388379
R2381 VTAIL.n55 VTAIL.n54 0.388379
R2382 VTAIL.n56 VTAIL.n20 0.388379
R2383 VTAIL.n155 VTAIL.n154 0.388379
R2384 VTAIL.n156 VTAIL.n120 0.388379
R2385 VTAIL.n255 VTAIL.n254 0.388379
R2386 VTAIL.n256 VTAIL.n220 0.388379
R2387 VTAIL.n656 VTAIL.n620 0.388379
R2388 VTAIL.n655 VTAIL.n654 0.388379
R2389 VTAIL.n556 VTAIL.n520 0.388379
R2390 VTAIL.n555 VTAIL.n554 0.388379
R2391 VTAIL.n456 VTAIL.n420 0.388379
R2392 VTAIL.n455 VTAIL.n454 0.388379
R2393 VTAIL.n356 VTAIL.n320 0.388379
R2394 VTAIL.n355 VTAIL.n354 0.388379
R2395 VTAIL VTAIL.n799 0.325931
R2396 VTAIL.n736 VTAIL.n735 0.155672
R2397 VTAIL.n736 VTAIL.n727 0.155672
R2398 VTAIL.n743 VTAIL.n727 0.155672
R2399 VTAIL.n744 VTAIL.n743 0.155672
R2400 VTAIL.n744 VTAIL.n723 0.155672
R2401 VTAIL.n752 VTAIL.n723 0.155672
R2402 VTAIL.n753 VTAIL.n752 0.155672
R2403 VTAIL.n753 VTAIL.n719 0.155672
R2404 VTAIL.n761 VTAIL.n719 0.155672
R2405 VTAIL.n762 VTAIL.n761 0.155672
R2406 VTAIL.n762 VTAIL.n715 0.155672
R2407 VTAIL.n769 VTAIL.n715 0.155672
R2408 VTAIL.n770 VTAIL.n769 0.155672
R2409 VTAIL.n770 VTAIL.n711 0.155672
R2410 VTAIL.n777 VTAIL.n711 0.155672
R2411 VTAIL.n778 VTAIL.n777 0.155672
R2412 VTAIL.n778 VTAIL.n707 0.155672
R2413 VTAIL.n785 VTAIL.n707 0.155672
R2414 VTAIL.n786 VTAIL.n785 0.155672
R2415 VTAIL.n786 VTAIL.n703 0.155672
R2416 VTAIL.n793 VTAIL.n703 0.155672
R2417 VTAIL.n794 VTAIL.n793 0.155672
R2418 VTAIL.n36 VTAIL.n35 0.155672
R2419 VTAIL.n36 VTAIL.n27 0.155672
R2420 VTAIL.n43 VTAIL.n27 0.155672
R2421 VTAIL.n44 VTAIL.n43 0.155672
R2422 VTAIL.n44 VTAIL.n23 0.155672
R2423 VTAIL.n52 VTAIL.n23 0.155672
R2424 VTAIL.n53 VTAIL.n52 0.155672
R2425 VTAIL.n53 VTAIL.n19 0.155672
R2426 VTAIL.n61 VTAIL.n19 0.155672
R2427 VTAIL.n62 VTAIL.n61 0.155672
R2428 VTAIL.n62 VTAIL.n15 0.155672
R2429 VTAIL.n69 VTAIL.n15 0.155672
R2430 VTAIL.n70 VTAIL.n69 0.155672
R2431 VTAIL.n70 VTAIL.n11 0.155672
R2432 VTAIL.n77 VTAIL.n11 0.155672
R2433 VTAIL.n78 VTAIL.n77 0.155672
R2434 VTAIL.n78 VTAIL.n7 0.155672
R2435 VTAIL.n85 VTAIL.n7 0.155672
R2436 VTAIL.n86 VTAIL.n85 0.155672
R2437 VTAIL.n86 VTAIL.n3 0.155672
R2438 VTAIL.n93 VTAIL.n3 0.155672
R2439 VTAIL.n94 VTAIL.n93 0.155672
R2440 VTAIL.n136 VTAIL.n135 0.155672
R2441 VTAIL.n136 VTAIL.n127 0.155672
R2442 VTAIL.n143 VTAIL.n127 0.155672
R2443 VTAIL.n144 VTAIL.n143 0.155672
R2444 VTAIL.n144 VTAIL.n123 0.155672
R2445 VTAIL.n152 VTAIL.n123 0.155672
R2446 VTAIL.n153 VTAIL.n152 0.155672
R2447 VTAIL.n153 VTAIL.n119 0.155672
R2448 VTAIL.n161 VTAIL.n119 0.155672
R2449 VTAIL.n162 VTAIL.n161 0.155672
R2450 VTAIL.n162 VTAIL.n115 0.155672
R2451 VTAIL.n169 VTAIL.n115 0.155672
R2452 VTAIL.n170 VTAIL.n169 0.155672
R2453 VTAIL.n170 VTAIL.n111 0.155672
R2454 VTAIL.n177 VTAIL.n111 0.155672
R2455 VTAIL.n178 VTAIL.n177 0.155672
R2456 VTAIL.n178 VTAIL.n107 0.155672
R2457 VTAIL.n185 VTAIL.n107 0.155672
R2458 VTAIL.n186 VTAIL.n185 0.155672
R2459 VTAIL.n186 VTAIL.n103 0.155672
R2460 VTAIL.n193 VTAIL.n103 0.155672
R2461 VTAIL.n194 VTAIL.n193 0.155672
R2462 VTAIL.n236 VTAIL.n235 0.155672
R2463 VTAIL.n236 VTAIL.n227 0.155672
R2464 VTAIL.n243 VTAIL.n227 0.155672
R2465 VTAIL.n244 VTAIL.n243 0.155672
R2466 VTAIL.n244 VTAIL.n223 0.155672
R2467 VTAIL.n252 VTAIL.n223 0.155672
R2468 VTAIL.n253 VTAIL.n252 0.155672
R2469 VTAIL.n253 VTAIL.n219 0.155672
R2470 VTAIL.n261 VTAIL.n219 0.155672
R2471 VTAIL.n262 VTAIL.n261 0.155672
R2472 VTAIL.n262 VTAIL.n215 0.155672
R2473 VTAIL.n269 VTAIL.n215 0.155672
R2474 VTAIL.n270 VTAIL.n269 0.155672
R2475 VTAIL.n270 VTAIL.n211 0.155672
R2476 VTAIL.n277 VTAIL.n211 0.155672
R2477 VTAIL.n278 VTAIL.n277 0.155672
R2478 VTAIL.n278 VTAIL.n207 0.155672
R2479 VTAIL.n285 VTAIL.n207 0.155672
R2480 VTAIL.n286 VTAIL.n285 0.155672
R2481 VTAIL.n286 VTAIL.n203 0.155672
R2482 VTAIL.n293 VTAIL.n203 0.155672
R2483 VTAIL.n294 VTAIL.n293 0.155672
R2484 VTAIL.n694 VTAIL.n693 0.155672
R2485 VTAIL.n693 VTAIL.n603 0.155672
R2486 VTAIL.n686 VTAIL.n603 0.155672
R2487 VTAIL.n686 VTAIL.n685 0.155672
R2488 VTAIL.n685 VTAIL.n607 0.155672
R2489 VTAIL.n678 VTAIL.n607 0.155672
R2490 VTAIL.n678 VTAIL.n677 0.155672
R2491 VTAIL.n677 VTAIL.n611 0.155672
R2492 VTAIL.n670 VTAIL.n611 0.155672
R2493 VTAIL.n670 VTAIL.n669 0.155672
R2494 VTAIL.n669 VTAIL.n615 0.155672
R2495 VTAIL.n662 VTAIL.n615 0.155672
R2496 VTAIL.n662 VTAIL.n661 0.155672
R2497 VTAIL.n661 VTAIL.n619 0.155672
R2498 VTAIL.n653 VTAIL.n619 0.155672
R2499 VTAIL.n653 VTAIL.n652 0.155672
R2500 VTAIL.n652 VTAIL.n623 0.155672
R2501 VTAIL.n645 VTAIL.n623 0.155672
R2502 VTAIL.n645 VTAIL.n644 0.155672
R2503 VTAIL.n644 VTAIL.n628 0.155672
R2504 VTAIL.n637 VTAIL.n628 0.155672
R2505 VTAIL.n637 VTAIL.n636 0.155672
R2506 VTAIL.n594 VTAIL.n593 0.155672
R2507 VTAIL.n593 VTAIL.n503 0.155672
R2508 VTAIL.n586 VTAIL.n503 0.155672
R2509 VTAIL.n586 VTAIL.n585 0.155672
R2510 VTAIL.n585 VTAIL.n507 0.155672
R2511 VTAIL.n578 VTAIL.n507 0.155672
R2512 VTAIL.n578 VTAIL.n577 0.155672
R2513 VTAIL.n577 VTAIL.n511 0.155672
R2514 VTAIL.n570 VTAIL.n511 0.155672
R2515 VTAIL.n570 VTAIL.n569 0.155672
R2516 VTAIL.n569 VTAIL.n515 0.155672
R2517 VTAIL.n562 VTAIL.n515 0.155672
R2518 VTAIL.n562 VTAIL.n561 0.155672
R2519 VTAIL.n561 VTAIL.n519 0.155672
R2520 VTAIL.n553 VTAIL.n519 0.155672
R2521 VTAIL.n553 VTAIL.n552 0.155672
R2522 VTAIL.n552 VTAIL.n523 0.155672
R2523 VTAIL.n545 VTAIL.n523 0.155672
R2524 VTAIL.n545 VTAIL.n544 0.155672
R2525 VTAIL.n544 VTAIL.n528 0.155672
R2526 VTAIL.n537 VTAIL.n528 0.155672
R2527 VTAIL.n537 VTAIL.n536 0.155672
R2528 VTAIL.n494 VTAIL.n493 0.155672
R2529 VTAIL.n493 VTAIL.n403 0.155672
R2530 VTAIL.n486 VTAIL.n403 0.155672
R2531 VTAIL.n486 VTAIL.n485 0.155672
R2532 VTAIL.n485 VTAIL.n407 0.155672
R2533 VTAIL.n478 VTAIL.n407 0.155672
R2534 VTAIL.n478 VTAIL.n477 0.155672
R2535 VTAIL.n477 VTAIL.n411 0.155672
R2536 VTAIL.n470 VTAIL.n411 0.155672
R2537 VTAIL.n470 VTAIL.n469 0.155672
R2538 VTAIL.n469 VTAIL.n415 0.155672
R2539 VTAIL.n462 VTAIL.n415 0.155672
R2540 VTAIL.n462 VTAIL.n461 0.155672
R2541 VTAIL.n461 VTAIL.n419 0.155672
R2542 VTAIL.n453 VTAIL.n419 0.155672
R2543 VTAIL.n453 VTAIL.n452 0.155672
R2544 VTAIL.n452 VTAIL.n423 0.155672
R2545 VTAIL.n445 VTAIL.n423 0.155672
R2546 VTAIL.n445 VTAIL.n444 0.155672
R2547 VTAIL.n444 VTAIL.n428 0.155672
R2548 VTAIL.n437 VTAIL.n428 0.155672
R2549 VTAIL.n437 VTAIL.n436 0.155672
R2550 VTAIL.n394 VTAIL.n393 0.155672
R2551 VTAIL.n393 VTAIL.n303 0.155672
R2552 VTAIL.n386 VTAIL.n303 0.155672
R2553 VTAIL.n386 VTAIL.n385 0.155672
R2554 VTAIL.n385 VTAIL.n307 0.155672
R2555 VTAIL.n378 VTAIL.n307 0.155672
R2556 VTAIL.n378 VTAIL.n377 0.155672
R2557 VTAIL.n377 VTAIL.n311 0.155672
R2558 VTAIL.n370 VTAIL.n311 0.155672
R2559 VTAIL.n370 VTAIL.n369 0.155672
R2560 VTAIL.n369 VTAIL.n315 0.155672
R2561 VTAIL.n362 VTAIL.n315 0.155672
R2562 VTAIL.n362 VTAIL.n361 0.155672
R2563 VTAIL.n361 VTAIL.n319 0.155672
R2564 VTAIL.n353 VTAIL.n319 0.155672
R2565 VTAIL.n353 VTAIL.n352 0.155672
R2566 VTAIL.n352 VTAIL.n323 0.155672
R2567 VTAIL.n345 VTAIL.n323 0.155672
R2568 VTAIL.n345 VTAIL.n344 0.155672
R2569 VTAIL.n344 VTAIL.n328 0.155672
R2570 VTAIL.n337 VTAIL.n328 0.155672
R2571 VTAIL.n337 VTAIL.n336 0.155672
R2572 VDD1 VDD1.n1 105.302
R2573 VDD1 VDD1.n0 63.267
R2574 VDD1.n0 VDD1.t2 1.09806
R2575 VDD1.n0 VDD1.t1 1.09806
R2576 VDD1.n1 VDD1.t0 1.09806
R2577 VDD1.n1 VDD1.t3 1.09806
R2578 VN.n0 VN.t2 867.495
R2579 VN.n1 VN.t3 867.495
R2580 VN.n0 VN.t1 867.471
R2581 VN.n1 VN.t0 867.471
R2582 VN VN.n1 115.239
R2583 VN VN.n0 70.265
R2584 VDD2.n2 VDD2.n0 104.778
R2585 VDD2.n2 VDD2.n1 63.2088
R2586 VDD2.n1 VDD2.t3 1.09806
R2587 VDD2.n1 VDD2.t0 1.09806
R2588 VDD2.n0 VDD2.t1 1.09806
R2589 VDD2.n0 VDD2.t2 1.09806
R2590 VDD2 VDD2.n2 0.0586897
C0 VP VTAIL 3.47074f
C1 VP VN 5.83561f
C2 VN VTAIL 3.45663f
C3 VDD1 VDD2 0.536834f
C4 VP VDD1 4.25268f
C5 VDD1 VTAIL 10.3857f
C6 VP VDD2 0.264935f
C7 VDD2 VTAIL 10.426201f
C8 VDD1 VN 0.147594f
C9 VDD2 VN 4.13556f
C10 VDD2 B 3.097583f
C11 VDD1 B 7.648991f
C12 VTAIL B 12.07692f
C13 VN B 9.1631f
C14 VP B 5.005805f
C15 VDD2.t1 B 0.41705f
C16 VDD2.t2 B 0.41705f
C17 VDD2.n0 B 4.64693f
C18 VDD2.t3 B 0.41705f
C19 VDD2.t0 B 0.41705f
C20 VDD2.n1 B 3.81042f
C21 VDD2.n2 B 4.29583f
C22 VN.t2 B 1.5249f
C23 VN.t1 B 1.52488f
C24 VN.n0 B 1.11857f
C25 VN.t3 B 1.5249f
C26 VN.t0 B 1.52488f
C27 VN.n1 B 2.09833f
C28 VDD1.t2 B 0.419675f
C29 VDD1.t1 B 0.419675f
C30 VDD1.n0 B 3.8347f
C31 VDD1.t0 B 0.419675f
C32 VDD1.t3 B 0.419675f
C33 VDD1.n1 B 4.70613f
C34 VTAIL.n0 B 0.009226f
C35 VTAIL.n1 B 0.020817f
C36 VTAIL.n2 B 0.009325f
C37 VTAIL.n3 B 0.01639f
C38 VTAIL.n4 B 0.008807f
C39 VTAIL.n5 B 0.020817f
C40 VTAIL.n6 B 0.009325f
C41 VTAIL.n7 B 0.01639f
C42 VTAIL.n8 B 0.008807f
C43 VTAIL.n9 B 0.020817f
C44 VTAIL.n10 B 0.009325f
C45 VTAIL.n11 B 0.01639f
C46 VTAIL.n12 B 0.008807f
C47 VTAIL.n13 B 0.020817f
C48 VTAIL.n14 B 0.009325f
C49 VTAIL.n15 B 0.01639f
C50 VTAIL.n16 B 0.008807f
C51 VTAIL.n17 B 0.020817f
C52 VTAIL.n18 B 0.009325f
C53 VTAIL.n19 B 0.01639f
C54 VTAIL.n20 B 0.008807f
C55 VTAIL.n21 B 0.020817f
C56 VTAIL.n22 B 0.009325f
C57 VTAIL.n23 B 0.01639f
C58 VTAIL.n24 B 0.008807f
C59 VTAIL.n25 B 0.020817f
C60 VTAIL.n26 B 0.009325f
C61 VTAIL.n27 B 0.01639f
C62 VTAIL.n28 B 0.008807f
C63 VTAIL.n29 B 0.020817f
C64 VTAIL.n30 B 0.009325f
C65 VTAIL.n31 B 0.156174f
C66 VTAIL.t2 B 0.035691f
C67 VTAIL.n32 B 0.015613f
C68 VTAIL.n33 B 0.014716f
C69 VTAIL.n34 B 0.008807f
C70 VTAIL.n35 B 1.26715f
C71 VTAIL.n36 B 0.01639f
C72 VTAIL.n37 B 0.008807f
C73 VTAIL.n38 B 0.009325f
C74 VTAIL.n39 B 0.020817f
C75 VTAIL.n40 B 0.020817f
C76 VTAIL.n41 B 0.009325f
C77 VTAIL.n42 B 0.008807f
C78 VTAIL.n43 B 0.01639f
C79 VTAIL.n44 B 0.01639f
C80 VTAIL.n45 B 0.008807f
C81 VTAIL.n46 B 0.009325f
C82 VTAIL.n47 B 0.020817f
C83 VTAIL.n48 B 0.020817f
C84 VTAIL.n49 B 0.020817f
C85 VTAIL.n50 B 0.009325f
C86 VTAIL.n51 B 0.008807f
C87 VTAIL.n52 B 0.01639f
C88 VTAIL.n53 B 0.01639f
C89 VTAIL.n54 B 0.008807f
C90 VTAIL.n55 B 0.009066f
C91 VTAIL.n56 B 0.009066f
C92 VTAIL.n57 B 0.020817f
C93 VTAIL.n58 B 0.020817f
C94 VTAIL.n59 B 0.009325f
C95 VTAIL.n60 B 0.008807f
C96 VTAIL.n61 B 0.01639f
C97 VTAIL.n62 B 0.01639f
C98 VTAIL.n63 B 0.008807f
C99 VTAIL.n64 B 0.009325f
C100 VTAIL.n65 B 0.020817f
C101 VTAIL.n66 B 0.020817f
C102 VTAIL.n67 B 0.009325f
C103 VTAIL.n68 B 0.008807f
C104 VTAIL.n69 B 0.01639f
C105 VTAIL.n70 B 0.01639f
C106 VTAIL.n71 B 0.008807f
C107 VTAIL.n72 B 0.009325f
C108 VTAIL.n73 B 0.020817f
C109 VTAIL.n74 B 0.020817f
C110 VTAIL.n75 B 0.009325f
C111 VTAIL.n76 B 0.008807f
C112 VTAIL.n77 B 0.01639f
C113 VTAIL.n78 B 0.01639f
C114 VTAIL.n79 B 0.008807f
C115 VTAIL.n80 B 0.009325f
C116 VTAIL.n81 B 0.020817f
C117 VTAIL.n82 B 0.020817f
C118 VTAIL.n83 B 0.009325f
C119 VTAIL.n84 B 0.008807f
C120 VTAIL.n85 B 0.01639f
C121 VTAIL.n86 B 0.01639f
C122 VTAIL.n87 B 0.008807f
C123 VTAIL.n88 B 0.009325f
C124 VTAIL.n89 B 0.020817f
C125 VTAIL.n90 B 0.020817f
C126 VTAIL.n91 B 0.009325f
C127 VTAIL.n92 B 0.008807f
C128 VTAIL.n93 B 0.01639f
C129 VTAIL.n94 B 0.041466f
C130 VTAIL.n95 B 0.008807f
C131 VTAIL.n96 B 0.009325f
C132 VTAIL.n97 B 0.041154f
C133 VTAIL.n98 B 0.034574f
C134 VTAIL.n99 B 0.063408f
C135 VTAIL.n100 B 0.009226f
C136 VTAIL.n101 B 0.020817f
C137 VTAIL.n102 B 0.009325f
C138 VTAIL.n103 B 0.01639f
C139 VTAIL.n104 B 0.008807f
C140 VTAIL.n105 B 0.020817f
C141 VTAIL.n106 B 0.009325f
C142 VTAIL.n107 B 0.01639f
C143 VTAIL.n108 B 0.008807f
C144 VTAIL.n109 B 0.020817f
C145 VTAIL.n110 B 0.009325f
C146 VTAIL.n111 B 0.01639f
C147 VTAIL.n112 B 0.008807f
C148 VTAIL.n113 B 0.020817f
C149 VTAIL.n114 B 0.009325f
C150 VTAIL.n115 B 0.01639f
C151 VTAIL.n116 B 0.008807f
C152 VTAIL.n117 B 0.020817f
C153 VTAIL.n118 B 0.009325f
C154 VTAIL.n119 B 0.01639f
C155 VTAIL.n120 B 0.008807f
C156 VTAIL.n121 B 0.020817f
C157 VTAIL.n122 B 0.009325f
C158 VTAIL.n123 B 0.01639f
C159 VTAIL.n124 B 0.008807f
C160 VTAIL.n125 B 0.020817f
C161 VTAIL.n126 B 0.009325f
C162 VTAIL.n127 B 0.01639f
C163 VTAIL.n128 B 0.008807f
C164 VTAIL.n129 B 0.020817f
C165 VTAIL.n130 B 0.009325f
C166 VTAIL.n131 B 0.156174f
C167 VTAIL.t7 B 0.035691f
C168 VTAIL.n132 B 0.015613f
C169 VTAIL.n133 B 0.014716f
C170 VTAIL.n134 B 0.008807f
C171 VTAIL.n135 B 1.26715f
C172 VTAIL.n136 B 0.01639f
C173 VTAIL.n137 B 0.008807f
C174 VTAIL.n138 B 0.009325f
C175 VTAIL.n139 B 0.020817f
C176 VTAIL.n140 B 0.020817f
C177 VTAIL.n141 B 0.009325f
C178 VTAIL.n142 B 0.008807f
C179 VTAIL.n143 B 0.01639f
C180 VTAIL.n144 B 0.01639f
C181 VTAIL.n145 B 0.008807f
C182 VTAIL.n146 B 0.009325f
C183 VTAIL.n147 B 0.020817f
C184 VTAIL.n148 B 0.020817f
C185 VTAIL.n149 B 0.020817f
C186 VTAIL.n150 B 0.009325f
C187 VTAIL.n151 B 0.008807f
C188 VTAIL.n152 B 0.01639f
C189 VTAIL.n153 B 0.01639f
C190 VTAIL.n154 B 0.008807f
C191 VTAIL.n155 B 0.009066f
C192 VTAIL.n156 B 0.009066f
C193 VTAIL.n157 B 0.020817f
C194 VTAIL.n158 B 0.020817f
C195 VTAIL.n159 B 0.009325f
C196 VTAIL.n160 B 0.008807f
C197 VTAIL.n161 B 0.01639f
C198 VTAIL.n162 B 0.01639f
C199 VTAIL.n163 B 0.008807f
C200 VTAIL.n164 B 0.009325f
C201 VTAIL.n165 B 0.020817f
C202 VTAIL.n166 B 0.020817f
C203 VTAIL.n167 B 0.009325f
C204 VTAIL.n168 B 0.008807f
C205 VTAIL.n169 B 0.01639f
C206 VTAIL.n170 B 0.01639f
C207 VTAIL.n171 B 0.008807f
C208 VTAIL.n172 B 0.009325f
C209 VTAIL.n173 B 0.020817f
C210 VTAIL.n174 B 0.020817f
C211 VTAIL.n175 B 0.009325f
C212 VTAIL.n176 B 0.008807f
C213 VTAIL.n177 B 0.01639f
C214 VTAIL.n178 B 0.01639f
C215 VTAIL.n179 B 0.008807f
C216 VTAIL.n180 B 0.009325f
C217 VTAIL.n181 B 0.020817f
C218 VTAIL.n182 B 0.020817f
C219 VTAIL.n183 B 0.009325f
C220 VTAIL.n184 B 0.008807f
C221 VTAIL.n185 B 0.01639f
C222 VTAIL.n186 B 0.01639f
C223 VTAIL.n187 B 0.008807f
C224 VTAIL.n188 B 0.009325f
C225 VTAIL.n189 B 0.020817f
C226 VTAIL.n190 B 0.020817f
C227 VTAIL.n191 B 0.009325f
C228 VTAIL.n192 B 0.008807f
C229 VTAIL.n193 B 0.01639f
C230 VTAIL.n194 B 0.041466f
C231 VTAIL.n195 B 0.008807f
C232 VTAIL.n196 B 0.009325f
C233 VTAIL.n197 B 0.041154f
C234 VTAIL.n198 B 0.034574f
C235 VTAIL.n199 B 0.080595f
C236 VTAIL.n200 B 0.009226f
C237 VTAIL.n201 B 0.020817f
C238 VTAIL.n202 B 0.009325f
C239 VTAIL.n203 B 0.01639f
C240 VTAIL.n204 B 0.008807f
C241 VTAIL.n205 B 0.020817f
C242 VTAIL.n206 B 0.009325f
C243 VTAIL.n207 B 0.01639f
C244 VTAIL.n208 B 0.008807f
C245 VTAIL.n209 B 0.020817f
C246 VTAIL.n210 B 0.009325f
C247 VTAIL.n211 B 0.01639f
C248 VTAIL.n212 B 0.008807f
C249 VTAIL.n213 B 0.020817f
C250 VTAIL.n214 B 0.009325f
C251 VTAIL.n215 B 0.01639f
C252 VTAIL.n216 B 0.008807f
C253 VTAIL.n217 B 0.020817f
C254 VTAIL.n218 B 0.009325f
C255 VTAIL.n219 B 0.01639f
C256 VTAIL.n220 B 0.008807f
C257 VTAIL.n221 B 0.020817f
C258 VTAIL.n222 B 0.009325f
C259 VTAIL.n223 B 0.01639f
C260 VTAIL.n224 B 0.008807f
C261 VTAIL.n225 B 0.020817f
C262 VTAIL.n226 B 0.009325f
C263 VTAIL.n227 B 0.01639f
C264 VTAIL.n228 B 0.008807f
C265 VTAIL.n229 B 0.020817f
C266 VTAIL.n230 B 0.009325f
C267 VTAIL.n231 B 0.156174f
C268 VTAIL.t4 B 0.035691f
C269 VTAIL.n232 B 0.015613f
C270 VTAIL.n233 B 0.014716f
C271 VTAIL.n234 B 0.008807f
C272 VTAIL.n235 B 1.26715f
C273 VTAIL.n236 B 0.01639f
C274 VTAIL.n237 B 0.008807f
C275 VTAIL.n238 B 0.009325f
C276 VTAIL.n239 B 0.020817f
C277 VTAIL.n240 B 0.020817f
C278 VTAIL.n241 B 0.009325f
C279 VTAIL.n242 B 0.008807f
C280 VTAIL.n243 B 0.01639f
C281 VTAIL.n244 B 0.01639f
C282 VTAIL.n245 B 0.008807f
C283 VTAIL.n246 B 0.009325f
C284 VTAIL.n247 B 0.020817f
C285 VTAIL.n248 B 0.020817f
C286 VTAIL.n249 B 0.020817f
C287 VTAIL.n250 B 0.009325f
C288 VTAIL.n251 B 0.008807f
C289 VTAIL.n252 B 0.01639f
C290 VTAIL.n253 B 0.01639f
C291 VTAIL.n254 B 0.008807f
C292 VTAIL.n255 B 0.009066f
C293 VTAIL.n256 B 0.009066f
C294 VTAIL.n257 B 0.020817f
C295 VTAIL.n258 B 0.020817f
C296 VTAIL.n259 B 0.009325f
C297 VTAIL.n260 B 0.008807f
C298 VTAIL.n261 B 0.01639f
C299 VTAIL.n262 B 0.01639f
C300 VTAIL.n263 B 0.008807f
C301 VTAIL.n264 B 0.009325f
C302 VTAIL.n265 B 0.020817f
C303 VTAIL.n266 B 0.020817f
C304 VTAIL.n267 B 0.009325f
C305 VTAIL.n268 B 0.008807f
C306 VTAIL.n269 B 0.01639f
C307 VTAIL.n270 B 0.01639f
C308 VTAIL.n271 B 0.008807f
C309 VTAIL.n272 B 0.009325f
C310 VTAIL.n273 B 0.020817f
C311 VTAIL.n274 B 0.020817f
C312 VTAIL.n275 B 0.009325f
C313 VTAIL.n276 B 0.008807f
C314 VTAIL.n277 B 0.01639f
C315 VTAIL.n278 B 0.01639f
C316 VTAIL.n279 B 0.008807f
C317 VTAIL.n280 B 0.009325f
C318 VTAIL.n281 B 0.020817f
C319 VTAIL.n282 B 0.020817f
C320 VTAIL.n283 B 0.009325f
C321 VTAIL.n284 B 0.008807f
C322 VTAIL.n285 B 0.01639f
C323 VTAIL.n286 B 0.01639f
C324 VTAIL.n287 B 0.008807f
C325 VTAIL.n288 B 0.009325f
C326 VTAIL.n289 B 0.020817f
C327 VTAIL.n290 B 0.020817f
C328 VTAIL.n291 B 0.009325f
C329 VTAIL.n292 B 0.008807f
C330 VTAIL.n293 B 0.01639f
C331 VTAIL.n294 B 0.041466f
C332 VTAIL.n295 B 0.008807f
C333 VTAIL.n296 B 0.009325f
C334 VTAIL.n297 B 0.041154f
C335 VTAIL.n298 B 0.034574f
C336 VTAIL.n299 B 1.14024f
C337 VTAIL.n300 B 0.009226f
C338 VTAIL.n301 B 0.020817f
C339 VTAIL.n302 B 0.009325f
C340 VTAIL.n303 B 0.01639f
C341 VTAIL.n304 B 0.008807f
C342 VTAIL.n305 B 0.020817f
C343 VTAIL.n306 B 0.009325f
C344 VTAIL.n307 B 0.01639f
C345 VTAIL.n308 B 0.008807f
C346 VTAIL.n309 B 0.020817f
C347 VTAIL.n310 B 0.009325f
C348 VTAIL.n311 B 0.01639f
C349 VTAIL.n312 B 0.008807f
C350 VTAIL.n313 B 0.020817f
C351 VTAIL.n314 B 0.009325f
C352 VTAIL.n315 B 0.01639f
C353 VTAIL.n316 B 0.008807f
C354 VTAIL.n317 B 0.020817f
C355 VTAIL.n318 B 0.009325f
C356 VTAIL.n319 B 0.01639f
C357 VTAIL.n320 B 0.008807f
C358 VTAIL.n321 B 0.020817f
C359 VTAIL.n322 B 0.009325f
C360 VTAIL.n323 B 0.01639f
C361 VTAIL.n324 B 0.008807f
C362 VTAIL.n325 B 0.020817f
C363 VTAIL.n326 B 0.020817f
C364 VTAIL.n327 B 0.009325f
C365 VTAIL.n328 B 0.01639f
C366 VTAIL.n329 B 0.008807f
C367 VTAIL.n330 B 0.020817f
C368 VTAIL.n331 B 0.009325f
C369 VTAIL.n332 B 0.156174f
C370 VTAIL.t0 B 0.035691f
C371 VTAIL.n333 B 0.015613f
C372 VTAIL.n334 B 0.014716f
C373 VTAIL.n335 B 0.008807f
C374 VTAIL.n336 B 1.26715f
C375 VTAIL.n337 B 0.01639f
C376 VTAIL.n338 B 0.008807f
C377 VTAIL.n339 B 0.009325f
C378 VTAIL.n340 B 0.020817f
C379 VTAIL.n341 B 0.020817f
C380 VTAIL.n342 B 0.009325f
C381 VTAIL.n343 B 0.008807f
C382 VTAIL.n344 B 0.01639f
C383 VTAIL.n345 B 0.01639f
C384 VTAIL.n346 B 0.008807f
C385 VTAIL.n347 B 0.009325f
C386 VTAIL.n348 B 0.020817f
C387 VTAIL.n349 B 0.020817f
C388 VTAIL.n350 B 0.009325f
C389 VTAIL.n351 B 0.008807f
C390 VTAIL.n352 B 0.01639f
C391 VTAIL.n353 B 0.01639f
C392 VTAIL.n354 B 0.008807f
C393 VTAIL.n355 B 0.009066f
C394 VTAIL.n356 B 0.009066f
C395 VTAIL.n357 B 0.020817f
C396 VTAIL.n358 B 0.020817f
C397 VTAIL.n359 B 0.009325f
C398 VTAIL.n360 B 0.008807f
C399 VTAIL.n361 B 0.01639f
C400 VTAIL.n362 B 0.01639f
C401 VTAIL.n363 B 0.008807f
C402 VTAIL.n364 B 0.009325f
C403 VTAIL.n365 B 0.020817f
C404 VTAIL.n366 B 0.020817f
C405 VTAIL.n367 B 0.009325f
C406 VTAIL.n368 B 0.008807f
C407 VTAIL.n369 B 0.01639f
C408 VTAIL.n370 B 0.01639f
C409 VTAIL.n371 B 0.008807f
C410 VTAIL.n372 B 0.009325f
C411 VTAIL.n373 B 0.020817f
C412 VTAIL.n374 B 0.020817f
C413 VTAIL.n375 B 0.009325f
C414 VTAIL.n376 B 0.008807f
C415 VTAIL.n377 B 0.01639f
C416 VTAIL.n378 B 0.01639f
C417 VTAIL.n379 B 0.008807f
C418 VTAIL.n380 B 0.009325f
C419 VTAIL.n381 B 0.020817f
C420 VTAIL.n382 B 0.020817f
C421 VTAIL.n383 B 0.009325f
C422 VTAIL.n384 B 0.008807f
C423 VTAIL.n385 B 0.01639f
C424 VTAIL.n386 B 0.01639f
C425 VTAIL.n387 B 0.008807f
C426 VTAIL.n388 B 0.009325f
C427 VTAIL.n389 B 0.020817f
C428 VTAIL.n390 B 0.020817f
C429 VTAIL.n391 B 0.009325f
C430 VTAIL.n392 B 0.008807f
C431 VTAIL.n393 B 0.01639f
C432 VTAIL.n394 B 0.041466f
C433 VTAIL.n395 B 0.008807f
C434 VTAIL.n396 B 0.009325f
C435 VTAIL.n397 B 0.041154f
C436 VTAIL.n398 B 0.034574f
C437 VTAIL.n399 B 1.14024f
C438 VTAIL.n400 B 0.009226f
C439 VTAIL.n401 B 0.020817f
C440 VTAIL.n402 B 0.009325f
C441 VTAIL.n403 B 0.01639f
C442 VTAIL.n404 B 0.008807f
C443 VTAIL.n405 B 0.020817f
C444 VTAIL.n406 B 0.009325f
C445 VTAIL.n407 B 0.01639f
C446 VTAIL.n408 B 0.008807f
C447 VTAIL.n409 B 0.020817f
C448 VTAIL.n410 B 0.009325f
C449 VTAIL.n411 B 0.01639f
C450 VTAIL.n412 B 0.008807f
C451 VTAIL.n413 B 0.020817f
C452 VTAIL.n414 B 0.009325f
C453 VTAIL.n415 B 0.01639f
C454 VTAIL.n416 B 0.008807f
C455 VTAIL.n417 B 0.020817f
C456 VTAIL.n418 B 0.009325f
C457 VTAIL.n419 B 0.01639f
C458 VTAIL.n420 B 0.008807f
C459 VTAIL.n421 B 0.020817f
C460 VTAIL.n422 B 0.009325f
C461 VTAIL.n423 B 0.01639f
C462 VTAIL.n424 B 0.008807f
C463 VTAIL.n425 B 0.020817f
C464 VTAIL.n426 B 0.020817f
C465 VTAIL.n427 B 0.009325f
C466 VTAIL.n428 B 0.01639f
C467 VTAIL.n429 B 0.008807f
C468 VTAIL.n430 B 0.020817f
C469 VTAIL.n431 B 0.009325f
C470 VTAIL.n432 B 0.156174f
C471 VTAIL.t3 B 0.035691f
C472 VTAIL.n433 B 0.015613f
C473 VTAIL.n434 B 0.014716f
C474 VTAIL.n435 B 0.008807f
C475 VTAIL.n436 B 1.26715f
C476 VTAIL.n437 B 0.01639f
C477 VTAIL.n438 B 0.008807f
C478 VTAIL.n439 B 0.009325f
C479 VTAIL.n440 B 0.020817f
C480 VTAIL.n441 B 0.020817f
C481 VTAIL.n442 B 0.009325f
C482 VTAIL.n443 B 0.008807f
C483 VTAIL.n444 B 0.01639f
C484 VTAIL.n445 B 0.01639f
C485 VTAIL.n446 B 0.008807f
C486 VTAIL.n447 B 0.009325f
C487 VTAIL.n448 B 0.020817f
C488 VTAIL.n449 B 0.020817f
C489 VTAIL.n450 B 0.009325f
C490 VTAIL.n451 B 0.008807f
C491 VTAIL.n452 B 0.01639f
C492 VTAIL.n453 B 0.01639f
C493 VTAIL.n454 B 0.008807f
C494 VTAIL.n455 B 0.009066f
C495 VTAIL.n456 B 0.009066f
C496 VTAIL.n457 B 0.020817f
C497 VTAIL.n458 B 0.020817f
C498 VTAIL.n459 B 0.009325f
C499 VTAIL.n460 B 0.008807f
C500 VTAIL.n461 B 0.01639f
C501 VTAIL.n462 B 0.01639f
C502 VTAIL.n463 B 0.008807f
C503 VTAIL.n464 B 0.009325f
C504 VTAIL.n465 B 0.020817f
C505 VTAIL.n466 B 0.020817f
C506 VTAIL.n467 B 0.009325f
C507 VTAIL.n468 B 0.008807f
C508 VTAIL.n469 B 0.01639f
C509 VTAIL.n470 B 0.01639f
C510 VTAIL.n471 B 0.008807f
C511 VTAIL.n472 B 0.009325f
C512 VTAIL.n473 B 0.020817f
C513 VTAIL.n474 B 0.020817f
C514 VTAIL.n475 B 0.009325f
C515 VTAIL.n476 B 0.008807f
C516 VTAIL.n477 B 0.01639f
C517 VTAIL.n478 B 0.01639f
C518 VTAIL.n479 B 0.008807f
C519 VTAIL.n480 B 0.009325f
C520 VTAIL.n481 B 0.020817f
C521 VTAIL.n482 B 0.020817f
C522 VTAIL.n483 B 0.009325f
C523 VTAIL.n484 B 0.008807f
C524 VTAIL.n485 B 0.01639f
C525 VTAIL.n486 B 0.01639f
C526 VTAIL.n487 B 0.008807f
C527 VTAIL.n488 B 0.009325f
C528 VTAIL.n489 B 0.020817f
C529 VTAIL.n490 B 0.020817f
C530 VTAIL.n491 B 0.009325f
C531 VTAIL.n492 B 0.008807f
C532 VTAIL.n493 B 0.01639f
C533 VTAIL.n494 B 0.041466f
C534 VTAIL.n495 B 0.008807f
C535 VTAIL.n496 B 0.009325f
C536 VTAIL.n497 B 0.041154f
C537 VTAIL.n498 B 0.034574f
C538 VTAIL.n499 B 0.080595f
C539 VTAIL.n500 B 0.009226f
C540 VTAIL.n501 B 0.020817f
C541 VTAIL.n502 B 0.009325f
C542 VTAIL.n503 B 0.01639f
C543 VTAIL.n504 B 0.008807f
C544 VTAIL.n505 B 0.020817f
C545 VTAIL.n506 B 0.009325f
C546 VTAIL.n507 B 0.01639f
C547 VTAIL.n508 B 0.008807f
C548 VTAIL.n509 B 0.020817f
C549 VTAIL.n510 B 0.009325f
C550 VTAIL.n511 B 0.01639f
C551 VTAIL.n512 B 0.008807f
C552 VTAIL.n513 B 0.020817f
C553 VTAIL.n514 B 0.009325f
C554 VTAIL.n515 B 0.01639f
C555 VTAIL.n516 B 0.008807f
C556 VTAIL.n517 B 0.020817f
C557 VTAIL.n518 B 0.009325f
C558 VTAIL.n519 B 0.01639f
C559 VTAIL.n520 B 0.008807f
C560 VTAIL.n521 B 0.020817f
C561 VTAIL.n522 B 0.009325f
C562 VTAIL.n523 B 0.01639f
C563 VTAIL.n524 B 0.008807f
C564 VTAIL.n525 B 0.020817f
C565 VTAIL.n526 B 0.020817f
C566 VTAIL.n527 B 0.009325f
C567 VTAIL.n528 B 0.01639f
C568 VTAIL.n529 B 0.008807f
C569 VTAIL.n530 B 0.020817f
C570 VTAIL.n531 B 0.009325f
C571 VTAIL.n532 B 0.156174f
C572 VTAIL.t6 B 0.035691f
C573 VTAIL.n533 B 0.015613f
C574 VTAIL.n534 B 0.014716f
C575 VTAIL.n535 B 0.008807f
C576 VTAIL.n536 B 1.26715f
C577 VTAIL.n537 B 0.01639f
C578 VTAIL.n538 B 0.008807f
C579 VTAIL.n539 B 0.009325f
C580 VTAIL.n540 B 0.020817f
C581 VTAIL.n541 B 0.020817f
C582 VTAIL.n542 B 0.009325f
C583 VTAIL.n543 B 0.008807f
C584 VTAIL.n544 B 0.01639f
C585 VTAIL.n545 B 0.01639f
C586 VTAIL.n546 B 0.008807f
C587 VTAIL.n547 B 0.009325f
C588 VTAIL.n548 B 0.020817f
C589 VTAIL.n549 B 0.020817f
C590 VTAIL.n550 B 0.009325f
C591 VTAIL.n551 B 0.008807f
C592 VTAIL.n552 B 0.01639f
C593 VTAIL.n553 B 0.01639f
C594 VTAIL.n554 B 0.008807f
C595 VTAIL.n555 B 0.009066f
C596 VTAIL.n556 B 0.009066f
C597 VTAIL.n557 B 0.020817f
C598 VTAIL.n558 B 0.020817f
C599 VTAIL.n559 B 0.009325f
C600 VTAIL.n560 B 0.008807f
C601 VTAIL.n561 B 0.01639f
C602 VTAIL.n562 B 0.01639f
C603 VTAIL.n563 B 0.008807f
C604 VTAIL.n564 B 0.009325f
C605 VTAIL.n565 B 0.020817f
C606 VTAIL.n566 B 0.020817f
C607 VTAIL.n567 B 0.009325f
C608 VTAIL.n568 B 0.008807f
C609 VTAIL.n569 B 0.01639f
C610 VTAIL.n570 B 0.01639f
C611 VTAIL.n571 B 0.008807f
C612 VTAIL.n572 B 0.009325f
C613 VTAIL.n573 B 0.020817f
C614 VTAIL.n574 B 0.020817f
C615 VTAIL.n575 B 0.009325f
C616 VTAIL.n576 B 0.008807f
C617 VTAIL.n577 B 0.01639f
C618 VTAIL.n578 B 0.01639f
C619 VTAIL.n579 B 0.008807f
C620 VTAIL.n580 B 0.009325f
C621 VTAIL.n581 B 0.020817f
C622 VTAIL.n582 B 0.020817f
C623 VTAIL.n583 B 0.009325f
C624 VTAIL.n584 B 0.008807f
C625 VTAIL.n585 B 0.01639f
C626 VTAIL.n586 B 0.01639f
C627 VTAIL.n587 B 0.008807f
C628 VTAIL.n588 B 0.009325f
C629 VTAIL.n589 B 0.020817f
C630 VTAIL.n590 B 0.020817f
C631 VTAIL.n591 B 0.009325f
C632 VTAIL.n592 B 0.008807f
C633 VTAIL.n593 B 0.01639f
C634 VTAIL.n594 B 0.041466f
C635 VTAIL.n595 B 0.008807f
C636 VTAIL.n596 B 0.009325f
C637 VTAIL.n597 B 0.041154f
C638 VTAIL.n598 B 0.034574f
C639 VTAIL.n599 B 0.080595f
C640 VTAIL.n600 B 0.009226f
C641 VTAIL.n601 B 0.020817f
C642 VTAIL.n602 B 0.009325f
C643 VTAIL.n603 B 0.01639f
C644 VTAIL.n604 B 0.008807f
C645 VTAIL.n605 B 0.020817f
C646 VTAIL.n606 B 0.009325f
C647 VTAIL.n607 B 0.01639f
C648 VTAIL.n608 B 0.008807f
C649 VTAIL.n609 B 0.020817f
C650 VTAIL.n610 B 0.009325f
C651 VTAIL.n611 B 0.01639f
C652 VTAIL.n612 B 0.008807f
C653 VTAIL.n613 B 0.020817f
C654 VTAIL.n614 B 0.009325f
C655 VTAIL.n615 B 0.01639f
C656 VTAIL.n616 B 0.008807f
C657 VTAIL.n617 B 0.020817f
C658 VTAIL.n618 B 0.009325f
C659 VTAIL.n619 B 0.01639f
C660 VTAIL.n620 B 0.008807f
C661 VTAIL.n621 B 0.020817f
C662 VTAIL.n622 B 0.009325f
C663 VTAIL.n623 B 0.01639f
C664 VTAIL.n624 B 0.008807f
C665 VTAIL.n625 B 0.020817f
C666 VTAIL.n626 B 0.020817f
C667 VTAIL.n627 B 0.009325f
C668 VTAIL.n628 B 0.01639f
C669 VTAIL.n629 B 0.008807f
C670 VTAIL.n630 B 0.020817f
C671 VTAIL.n631 B 0.009325f
C672 VTAIL.n632 B 0.156174f
C673 VTAIL.t5 B 0.035691f
C674 VTAIL.n633 B 0.015613f
C675 VTAIL.n634 B 0.014716f
C676 VTAIL.n635 B 0.008807f
C677 VTAIL.n636 B 1.26715f
C678 VTAIL.n637 B 0.01639f
C679 VTAIL.n638 B 0.008807f
C680 VTAIL.n639 B 0.009325f
C681 VTAIL.n640 B 0.020817f
C682 VTAIL.n641 B 0.020817f
C683 VTAIL.n642 B 0.009325f
C684 VTAIL.n643 B 0.008807f
C685 VTAIL.n644 B 0.01639f
C686 VTAIL.n645 B 0.01639f
C687 VTAIL.n646 B 0.008807f
C688 VTAIL.n647 B 0.009325f
C689 VTAIL.n648 B 0.020817f
C690 VTAIL.n649 B 0.020817f
C691 VTAIL.n650 B 0.009325f
C692 VTAIL.n651 B 0.008807f
C693 VTAIL.n652 B 0.01639f
C694 VTAIL.n653 B 0.01639f
C695 VTAIL.n654 B 0.008807f
C696 VTAIL.n655 B 0.009066f
C697 VTAIL.n656 B 0.009066f
C698 VTAIL.n657 B 0.020817f
C699 VTAIL.n658 B 0.020817f
C700 VTAIL.n659 B 0.009325f
C701 VTAIL.n660 B 0.008807f
C702 VTAIL.n661 B 0.01639f
C703 VTAIL.n662 B 0.01639f
C704 VTAIL.n663 B 0.008807f
C705 VTAIL.n664 B 0.009325f
C706 VTAIL.n665 B 0.020817f
C707 VTAIL.n666 B 0.020817f
C708 VTAIL.n667 B 0.009325f
C709 VTAIL.n668 B 0.008807f
C710 VTAIL.n669 B 0.01639f
C711 VTAIL.n670 B 0.01639f
C712 VTAIL.n671 B 0.008807f
C713 VTAIL.n672 B 0.009325f
C714 VTAIL.n673 B 0.020817f
C715 VTAIL.n674 B 0.020817f
C716 VTAIL.n675 B 0.009325f
C717 VTAIL.n676 B 0.008807f
C718 VTAIL.n677 B 0.01639f
C719 VTAIL.n678 B 0.01639f
C720 VTAIL.n679 B 0.008807f
C721 VTAIL.n680 B 0.009325f
C722 VTAIL.n681 B 0.020817f
C723 VTAIL.n682 B 0.020817f
C724 VTAIL.n683 B 0.009325f
C725 VTAIL.n684 B 0.008807f
C726 VTAIL.n685 B 0.01639f
C727 VTAIL.n686 B 0.01639f
C728 VTAIL.n687 B 0.008807f
C729 VTAIL.n688 B 0.009325f
C730 VTAIL.n689 B 0.020817f
C731 VTAIL.n690 B 0.020817f
C732 VTAIL.n691 B 0.009325f
C733 VTAIL.n692 B 0.008807f
C734 VTAIL.n693 B 0.01639f
C735 VTAIL.n694 B 0.041466f
C736 VTAIL.n695 B 0.008807f
C737 VTAIL.n696 B 0.009325f
C738 VTAIL.n697 B 0.041154f
C739 VTAIL.n698 B 0.034574f
C740 VTAIL.n699 B 1.14024f
C741 VTAIL.n700 B 0.009226f
C742 VTAIL.n701 B 0.020817f
C743 VTAIL.n702 B 0.009325f
C744 VTAIL.n703 B 0.01639f
C745 VTAIL.n704 B 0.008807f
C746 VTAIL.n705 B 0.020817f
C747 VTAIL.n706 B 0.009325f
C748 VTAIL.n707 B 0.01639f
C749 VTAIL.n708 B 0.008807f
C750 VTAIL.n709 B 0.020817f
C751 VTAIL.n710 B 0.009325f
C752 VTAIL.n711 B 0.01639f
C753 VTAIL.n712 B 0.008807f
C754 VTAIL.n713 B 0.020817f
C755 VTAIL.n714 B 0.009325f
C756 VTAIL.n715 B 0.01639f
C757 VTAIL.n716 B 0.008807f
C758 VTAIL.n717 B 0.020817f
C759 VTAIL.n718 B 0.009325f
C760 VTAIL.n719 B 0.01639f
C761 VTAIL.n720 B 0.008807f
C762 VTAIL.n721 B 0.020817f
C763 VTAIL.n722 B 0.009325f
C764 VTAIL.n723 B 0.01639f
C765 VTAIL.n724 B 0.008807f
C766 VTAIL.n725 B 0.020817f
C767 VTAIL.n726 B 0.009325f
C768 VTAIL.n727 B 0.01639f
C769 VTAIL.n728 B 0.008807f
C770 VTAIL.n729 B 0.020817f
C771 VTAIL.n730 B 0.009325f
C772 VTAIL.n731 B 0.156174f
C773 VTAIL.t1 B 0.035691f
C774 VTAIL.n732 B 0.015613f
C775 VTAIL.n733 B 0.014716f
C776 VTAIL.n734 B 0.008807f
C777 VTAIL.n735 B 1.26715f
C778 VTAIL.n736 B 0.01639f
C779 VTAIL.n737 B 0.008807f
C780 VTAIL.n738 B 0.009325f
C781 VTAIL.n739 B 0.020817f
C782 VTAIL.n740 B 0.020817f
C783 VTAIL.n741 B 0.009325f
C784 VTAIL.n742 B 0.008807f
C785 VTAIL.n743 B 0.01639f
C786 VTAIL.n744 B 0.01639f
C787 VTAIL.n745 B 0.008807f
C788 VTAIL.n746 B 0.009325f
C789 VTAIL.n747 B 0.020817f
C790 VTAIL.n748 B 0.020817f
C791 VTAIL.n749 B 0.020817f
C792 VTAIL.n750 B 0.009325f
C793 VTAIL.n751 B 0.008807f
C794 VTAIL.n752 B 0.01639f
C795 VTAIL.n753 B 0.01639f
C796 VTAIL.n754 B 0.008807f
C797 VTAIL.n755 B 0.009066f
C798 VTAIL.n756 B 0.009066f
C799 VTAIL.n757 B 0.020817f
C800 VTAIL.n758 B 0.020817f
C801 VTAIL.n759 B 0.009325f
C802 VTAIL.n760 B 0.008807f
C803 VTAIL.n761 B 0.01639f
C804 VTAIL.n762 B 0.01639f
C805 VTAIL.n763 B 0.008807f
C806 VTAIL.n764 B 0.009325f
C807 VTAIL.n765 B 0.020817f
C808 VTAIL.n766 B 0.020817f
C809 VTAIL.n767 B 0.009325f
C810 VTAIL.n768 B 0.008807f
C811 VTAIL.n769 B 0.01639f
C812 VTAIL.n770 B 0.01639f
C813 VTAIL.n771 B 0.008807f
C814 VTAIL.n772 B 0.009325f
C815 VTAIL.n773 B 0.020817f
C816 VTAIL.n774 B 0.020817f
C817 VTAIL.n775 B 0.009325f
C818 VTAIL.n776 B 0.008807f
C819 VTAIL.n777 B 0.01639f
C820 VTAIL.n778 B 0.01639f
C821 VTAIL.n779 B 0.008807f
C822 VTAIL.n780 B 0.009325f
C823 VTAIL.n781 B 0.020817f
C824 VTAIL.n782 B 0.020817f
C825 VTAIL.n783 B 0.009325f
C826 VTAIL.n784 B 0.008807f
C827 VTAIL.n785 B 0.01639f
C828 VTAIL.n786 B 0.01639f
C829 VTAIL.n787 B 0.008807f
C830 VTAIL.n788 B 0.009325f
C831 VTAIL.n789 B 0.020817f
C832 VTAIL.n790 B 0.020817f
C833 VTAIL.n791 B 0.009325f
C834 VTAIL.n792 B 0.008807f
C835 VTAIL.n793 B 0.01639f
C836 VTAIL.n794 B 0.041466f
C837 VTAIL.n795 B 0.008807f
C838 VTAIL.n796 B 0.009325f
C839 VTAIL.n797 B 0.041154f
C840 VTAIL.n798 B 0.034574f
C841 VTAIL.n799 B 1.11691f
C842 VP.t2 B 1.55626f
C843 VP.t1 B 1.55628f
C844 VP.n0 B 2.12264f
C845 VP.n1 B 4.04209f
C846 VP.t3 B 1.54213f
C847 VP.n2 B 0.584847f
C848 VP.t0 B 1.54213f
C849 VP.n3 B 0.584847f
C850 VP.n4 B 0.041726f
.ends

