* NGSPICE file created from diff_pair_sample_1533.ext - technology: sky130A

.subckt diff_pair_sample_1533 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=4.6137 pd=24.44 as=1.95195 ps=12.16 w=11.83 l=2.64
X1 VDD2.t4 VN.t1 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=1.95195 pd=12.16 as=4.6137 ps=24.44 w=11.83 l=2.64
X2 VDD1.t5 VP.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.95195 pd=12.16 as=4.6137 ps=24.44 w=11.83 l=2.64
X3 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=4.6137 pd=24.44 as=0 ps=0 w=11.83 l=2.64
X4 VDD2.t3 VN.t2 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=4.6137 pd=24.44 as=1.95195 ps=12.16 w=11.83 l=2.64
X5 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=4.6137 pd=24.44 as=0 ps=0 w=11.83 l=2.64
X6 VDD1.t4 VP.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.95195 pd=12.16 as=4.6137 ps=24.44 w=11.83 l=2.64
X7 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.6137 pd=24.44 as=0 ps=0 w=11.83 l=2.64
X8 VTAIL.t11 VN.t3 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.95195 pd=12.16 as=1.95195 ps=12.16 w=11.83 l=2.64
X9 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.6137 pd=24.44 as=0 ps=0 w=11.83 l=2.64
X10 VDD2.t1 VN.t4 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.95195 pd=12.16 as=4.6137 ps=24.44 w=11.83 l=2.64
X11 VTAIL.t9 VN.t5 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=1.95195 pd=12.16 as=1.95195 ps=12.16 w=11.83 l=2.64
X12 VDD1.t3 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.6137 pd=24.44 as=1.95195 ps=12.16 w=11.83 l=2.64
X13 VTAIL.t5 VP.t3 VDD1.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=1.95195 pd=12.16 as=1.95195 ps=12.16 w=11.83 l=2.64
X14 VTAIL.t2 VP.t4 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.95195 pd=12.16 as=1.95195 ps=12.16 w=11.83 l=2.64
X15 VDD1.t0 VP.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.6137 pd=24.44 as=1.95195 ps=12.16 w=11.83 l=2.64
R0 VN.n29 VN.n16 161.3
R1 VN.n28 VN.n27 161.3
R2 VN.n26 VN.n17 161.3
R3 VN.n25 VN.n24 161.3
R4 VN.n23 VN.n18 161.3
R5 VN.n22 VN.n21 161.3
R6 VN.n13 VN.n0 161.3
R7 VN.n12 VN.n11 161.3
R8 VN.n10 VN.n1 161.3
R9 VN.n9 VN.n8 161.3
R10 VN.n7 VN.n2 161.3
R11 VN.n6 VN.n5 161.3
R12 VN.n4 VN.t2 141.812
R13 VN.n20 VN.t4 141.812
R14 VN.n3 VN.t3 107.995
R15 VN.n14 VN.t1 107.995
R16 VN.n19 VN.t5 107.995
R17 VN.n30 VN.t0 107.995
R18 VN.n15 VN.n14 99.991
R19 VN.n31 VN.n30 99.991
R20 VN.n4 VN.n3 60.2677
R21 VN.n20 VN.n19 60.2677
R22 VN.n8 VN.n1 56.5193
R23 VN.n24 VN.n17 56.5193
R24 VN VN.n31 49.0247
R25 VN.n7 VN.n6 24.4675
R26 VN.n8 VN.n7 24.4675
R27 VN.n12 VN.n1 24.4675
R28 VN.n13 VN.n12 24.4675
R29 VN.n24 VN.n23 24.4675
R30 VN.n23 VN.n22 24.4675
R31 VN.n29 VN.n28 24.4675
R32 VN.n28 VN.n17 24.4675
R33 VN.n6 VN.n3 12.234
R34 VN.n22 VN.n19 12.234
R35 VN.n14 VN.n13 10.766
R36 VN.n30 VN.n29 10.766
R37 VN.n21 VN.n20 6.80183
R38 VN.n5 VN.n4 6.80183
R39 VN.n31 VN.n16 0.278367
R40 VN.n15 VN.n0 0.278367
R41 VN.n27 VN.n16 0.189894
R42 VN.n27 VN.n26 0.189894
R43 VN.n26 VN.n25 0.189894
R44 VN.n25 VN.n18 0.189894
R45 VN.n21 VN.n18 0.189894
R46 VN.n5 VN.n2 0.189894
R47 VN.n9 VN.n2 0.189894
R48 VN.n10 VN.n9 0.189894
R49 VN.n11 VN.n10 0.189894
R50 VN.n11 VN.n0 0.189894
R51 VN VN.n15 0.153454
R52 VTAIL.n7 VTAIL.t6 48.3325
R53 VTAIL.n11 VTAIL.t8 48.3323
R54 VTAIL.n2 VTAIL.t3 48.3323
R55 VTAIL.n10 VTAIL.t4 48.3323
R56 VTAIL.n9 VTAIL.n8 46.6588
R57 VTAIL.n6 VTAIL.n5 46.6588
R58 VTAIL.n1 VTAIL.n0 46.6586
R59 VTAIL.n4 VTAIL.n3 46.6586
R60 VTAIL.n6 VTAIL.n4 27.6858
R61 VTAIL.n11 VTAIL.n10 25.1255
R62 VTAIL.n7 VTAIL.n6 2.56084
R63 VTAIL.n10 VTAIL.n9 2.56084
R64 VTAIL.n4 VTAIL.n2 2.56084
R65 VTAIL VTAIL.n11 1.86257
R66 VTAIL.n9 VTAIL.n7 1.7505
R67 VTAIL.n2 VTAIL.n1 1.7505
R68 VTAIL.n0 VTAIL.t10 1.67421
R69 VTAIL.n0 VTAIL.t11 1.67421
R70 VTAIL.n3 VTAIL.t0 1.67421
R71 VTAIL.n3 VTAIL.t5 1.67421
R72 VTAIL.n8 VTAIL.t1 1.67421
R73 VTAIL.n8 VTAIL.t2 1.67421
R74 VTAIL.n5 VTAIL.t7 1.67421
R75 VTAIL.n5 VTAIL.t9 1.67421
R76 VTAIL VTAIL.n1 0.698776
R77 VDD2.n1 VDD2.t3 66.876
R78 VDD2.n2 VDD2.t5 65.0113
R79 VDD2.n1 VDD2.n0 63.9221
R80 VDD2 VDD2.n3 63.9193
R81 VDD2.n2 VDD2.n1 42.2347
R82 VDD2 VDD2.n2 1.97895
R83 VDD2.n3 VDD2.t0 1.67421
R84 VDD2.n3 VDD2.t1 1.67421
R85 VDD2.n0 VDD2.t2 1.67421
R86 VDD2.n0 VDD2.t4 1.67421
R87 B.n814 B.n813 585
R88 B.n310 B.n126 585
R89 B.n309 B.n308 585
R90 B.n307 B.n306 585
R91 B.n305 B.n304 585
R92 B.n303 B.n302 585
R93 B.n301 B.n300 585
R94 B.n299 B.n298 585
R95 B.n297 B.n296 585
R96 B.n295 B.n294 585
R97 B.n293 B.n292 585
R98 B.n291 B.n290 585
R99 B.n289 B.n288 585
R100 B.n287 B.n286 585
R101 B.n285 B.n284 585
R102 B.n283 B.n282 585
R103 B.n281 B.n280 585
R104 B.n279 B.n278 585
R105 B.n277 B.n276 585
R106 B.n275 B.n274 585
R107 B.n273 B.n272 585
R108 B.n271 B.n270 585
R109 B.n269 B.n268 585
R110 B.n267 B.n266 585
R111 B.n265 B.n264 585
R112 B.n263 B.n262 585
R113 B.n261 B.n260 585
R114 B.n259 B.n258 585
R115 B.n257 B.n256 585
R116 B.n255 B.n254 585
R117 B.n253 B.n252 585
R118 B.n251 B.n250 585
R119 B.n249 B.n248 585
R120 B.n247 B.n246 585
R121 B.n245 B.n244 585
R122 B.n243 B.n242 585
R123 B.n241 B.n240 585
R124 B.n239 B.n238 585
R125 B.n237 B.n236 585
R126 B.n235 B.n234 585
R127 B.n233 B.n232 585
R128 B.n230 B.n229 585
R129 B.n228 B.n227 585
R130 B.n226 B.n225 585
R131 B.n224 B.n223 585
R132 B.n222 B.n221 585
R133 B.n220 B.n219 585
R134 B.n218 B.n217 585
R135 B.n216 B.n215 585
R136 B.n214 B.n213 585
R137 B.n212 B.n211 585
R138 B.n209 B.n208 585
R139 B.n207 B.n206 585
R140 B.n205 B.n204 585
R141 B.n203 B.n202 585
R142 B.n201 B.n200 585
R143 B.n199 B.n198 585
R144 B.n197 B.n196 585
R145 B.n195 B.n194 585
R146 B.n193 B.n192 585
R147 B.n191 B.n190 585
R148 B.n189 B.n188 585
R149 B.n187 B.n186 585
R150 B.n185 B.n184 585
R151 B.n183 B.n182 585
R152 B.n181 B.n180 585
R153 B.n179 B.n178 585
R154 B.n177 B.n176 585
R155 B.n175 B.n174 585
R156 B.n173 B.n172 585
R157 B.n171 B.n170 585
R158 B.n169 B.n168 585
R159 B.n167 B.n166 585
R160 B.n165 B.n164 585
R161 B.n163 B.n162 585
R162 B.n161 B.n160 585
R163 B.n159 B.n158 585
R164 B.n157 B.n156 585
R165 B.n155 B.n154 585
R166 B.n153 B.n152 585
R167 B.n151 B.n150 585
R168 B.n149 B.n148 585
R169 B.n147 B.n146 585
R170 B.n145 B.n144 585
R171 B.n143 B.n142 585
R172 B.n141 B.n140 585
R173 B.n139 B.n138 585
R174 B.n137 B.n136 585
R175 B.n135 B.n134 585
R176 B.n133 B.n132 585
R177 B.n81 B.n80 585
R178 B.n819 B.n818 585
R179 B.n812 B.n127 585
R180 B.n127 B.n78 585
R181 B.n811 B.n77 585
R182 B.n823 B.n77 585
R183 B.n810 B.n76 585
R184 B.n824 B.n76 585
R185 B.n809 B.n75 585
R186 B.n825 B.n75 585
R187 B.n808 B.n807 585
R188 B.n807 B.n71 585
R189 B.n806 B.n70 585
R190 B.n831 B.n70 585
R191 B.n805 B.n69 585
R192 B.n832 B.n69 585
R193 B.n804 B.n68 585
R194 B.n833 B.n68 585
R195 B.n803 B.n802 585
R196 B.n802 B.n64 585
R197 B.n801 B.n63 585
R198 B.n839 B.n63 585
R199 B.n800 B.n62 585
R200 B.n840 B.n62 585
R201 B.n799 B.n61 585
R202 B.n841 B.n61 585
R203 B.n798 B.n797 585
R204 B.n797 B.n57 585
R205 B.n796 B.n56 585
R206 B.n847 B.n56 585
R207 B.n795 B.n55 585
R208 B.n848 B.n55 585
R209 B.n794 B.n54 585
R210 B.n849 B.n54 585
R211 B.n793 B.n792 585
R212 B.n792 B.n50 585
R213 B.n791 B.n49 585
R214 B.n855 B.n49 585
R215 B.n790 B.n48 585
R216 B.n856 B.n48 585
R217 B.n789 B.n47 585
R218 B.n857 B.n47 585
R219 B.n788 B.n787 585
R220 B.n787 B.n43 585
R221 B.n786 B.n42 585
R222 B.n863 B.n42 585
R223 B.n785 B.n41 585
R224 B.n864 B.n41 585
R225 B.n784 B.n40 585
R226 B.n865 B.n40 585
R227 B.n783 B.n782 585
R228 B.n782 B.n36 585
R229 B.n781 B.n35 585
R230 B.n871 B.n35 585
R231 B.n780 B.n34 585
R232 B.n872 B.n34 585
R233 B.n779 B.n33 585
R234 B.n873 B.n33 585
R235 B.n778 B.n777 585
R236 B.n777 B.n32 585
R237 B.n776 B.n28 585
R238 B.n879 B.n28 585
R239 B.n775 B.n27 585
R240 B.n880 B.n27 585
R241 B.n774 B.n26 585
R242 B.n881 B.n26 585
R243 B.n773 B.n772 585
R244 B.n772 B.n22 585
R245 B.n771 B.n21 585
R246 B.n887 B.n21 585
R247 B.n770 B.n20 585
R248 B.n888 B.n20 585
R249 B.n769 B.n19 585
R250 B.n889 B.n19 585
R251 B.n768 B.n767 585
R252 B.n767 B.n15 585
R253 B.n766 B.n14 585
R254 B.n895 B.n14 585
R255 B.n765 B.n13 585
R256 B.n896 B.n13 585
R257 B.n764 B.n12 585
R258 B.n897 B.n12 585
R259 B.n763 B.n762 585
R260 B.n762 B.n8 585
R261 B.n761 B.n7 585
R262 B.n903 B.n7 585
R263 B.n760 B.n6 585
R264 B.n904 B.n6 585
R265 B.n759 B.n5 585
R266 B.n905 B.n5 585
R267 B.n758 B.n757 585
R268 B.n757 B.n4 585
R269 B.n756 B.n311 585
R270 B.n756 B.n755 585
R271 B.n746 B.n312 585
R272 B.n313 B.n312 585
R273 B.n748 B.n747 585
R274 B.n749 B.n748 585
R275 B.n745 B.n318 585
R276 B.n318 B.n317 585
R277 B.n744 B.n743 585
R278 B.n743 B.n742 585
R279 B.n320 B.n319 585
R280 B.n321 B.n320 585
R281 B.n735 B.n734 585
R282 B.n736 B.n735 585
R283 B.n733 B.n326 585
R284 B.n326 B.n325 585
R285 B.n732 B.n731 585
R286 B.n731 B.n730 585
R287 B.n328 B.n327 585
R288 B.n329 B.n328 585
R289 B.n723 B.n722 585
R290 B.n724 B.n723 585
R291 B.n721 B.n334 585
R292 B.n334 B.n333 585
R293 B.n720 B.n719 585
R294 B.n719 B.n718 585
R295 B.n336 B.n335 585
R296 B.n711 B.n336 585
R297 B.n710 B.n709 585
R298 B.n712 B.n710 585
R299 B.n708 B.n341 585
R300 B.n341 B.n340 585
R301 B.n707 B.n706 585
R302 B.n706 B.n705 585
R303 B.n343 B.n342 585
R304 B.n344 B.n343 585
R305 B.n698 B.n697 585
R306 B.n699 B.n698 585
R307 B.n696 B.n349 585
R308 B.n349 B.n348 585
R309 B.n695 B.n694 585
R310 B.n694 B.n693 585
R311 B.n351 B.n350 585
R312 B.n352 B.n351 585
R313 B.n686 B.n685 585
R314 B.n687 B.n686 585
R315 B.n684 B.n357 585
R316 B.n357 B.n356 585
R317 B.n683 B.n682 585
R318 B.n682 B.n681 585
R319 B.n359 B.n358 585
R320 B.n360 B.n359 585
R321 B.n674 B.n673 585
R322 B.n675 B.n674 585
R323 B.n672 B.n365 585
R324 B.n365 B.n364 585
R325 B.n671 B.n670 585
R326 B.n670 B.n669 585
R327 B.n367 B.n366 585
R328 B.n368 B.n367 585
R329 B.n662 B.n661 585
R330 B.n663 B.n662 585
R331 B.n660 B.n373 585
R332 B.n373 B.n372 585
R333 B.n659 B.n658 585
R334 B.n658 B.n657 585
R335 B.n375 B.n374 585
R336 B.n376 B.n375 585
R337 B.n650 B.n649 585
R338 B.n651 B.n650 585
R339 B.n648 B.n381 585
R340 B.n381 B.n380 585
R341 B.n647 B.n646 585
R342 B.n646 B.n645 585
R343 B.n383 B.n382 585
R344 B.n384 B.n383 585
R345 B.n638 B.n637 585
R346 B.n639 B.n638 585
R347 B.n636 B.n389 585
R348 B.n389 B.n388 585
R349 B.n635 B.n634 585
R350 B.n634 B.n633 585
R351 B.n391 B.n390 585
R352 B.n392 B.n391 585
R353 B.n629 B.n628 585
R354 B.n395 B.n394 585
R355 B.n625 B.n624 585
R356 B.n626 B.n625 585
R357 B.n623 B.n441 585
R358 B.n622 B.n621 585
R359 B.n620 B.n619 585
R360 B.n618 B.n617 585
R361 B.n616 B.n615 585
R362 B.n614 B.n613 585
R363 B.n612 B.n611 585
R364 B.n610 B.n609 585
R365 B.n608 B.n607 585
R366 B.n606 B.n605 585
R367 B.n604 B.n603 585
R368 B.n602 B.n601 585
R369 B.n600 B.n599 585
R370 B.n598 B.n597 585
R371 B.n596 B.n595 585
R372 B.n594 B.n593 585
R373 B.n592 B.n591 585
R374 B.n590 B.n589 585
R375 B.n588 B.n587 585
R376 B.n586 B.n585 585
R377 B.n584 B.n583 585
R378 B.n582 B.n581 585
R379 B.n580 B.n579 585
R380 B.n578 B.n577 585
R381 B.n576 B.n575 585
R382 B.n574 B.n573 585
R383 B.n572 B.n571 585
R384 B.n570 B.n569 585
R385 B.n568 B.n567 585
R386 B.n566 B.n565 585
R387 B.n564 B.n563 585
R388 B.n562 B.n561 585
R389 B.n560 B.n559 585
R390 B.n558 B.n557 585
R391 B.n556 B.n555 585
R392 B.n554 B.n553 585
R393 B.n552 B.n551 585
R394 B.n550 B.n549 585
R395 B.n548 B.n547 585
R396 B.n546 B.n545 585
R397 B.n544 B.n543 585
R398 B.n542 B.n541 585
R399 B.n540 B.n539 585
R400 B.n538 B.n537 585
R401 B.n536 B.n535 585
R402 B.n534 B.n533 585
R403 B.n532 B.n531 585
R404 B.n530 B.n529 585
R405 B.n528 B.n527 585
R406 B.n526 B.n525 585
R407 B.n524 B.n523 585
R408 B.n522 B.n521 585
R409 B.n520 B.n519 585
R410 B.n518 B.n517 585
R411 B.n516 B.n515 585
R412 B.n514 B.n513 585
R413 B.n512 B.n511 585
R414 B.n510 B.n509 585
R415 B.n508 B.n507 585
R416 B.n506 B.n505 585
R417 B.n504 B.n503 585
R418 B.n502 B.n501 585
R419 B.n500 B.n499 585
R420 B.n498 B.n497 585
R421 B.n496 B.n495 585
R422 B.n494 B.n493 585
R423 B.n492 B.n491 585
R424 B.n490 B.n489 585
R425 B.n488 B.n487 585
R426 B.n486 B.n485 585
R427 B.n484 B.n483 585
R428 B.n482 B.n481 585
R429 B.n480 B.n479 585
R430 B.n478 B.n477 585
R431 B.n476 B.n475 585
R432 B.n474 B.n473 585
R433 B.n472 B.n471 585
R434 B.n470 B.n469 585
R435 B.n468 B.n467 585
R436 B.n466 B.n465 585
R437 B.n464 B.n463 585
R438 B.n462 B.n461 585
R439 B.n460 B.n459 585
R440 B.n458 B.n457 585
R441 B.n456 B.n455 585
R442 B.n454 B.n453 585
R443 B.n452 B.n451 585
R444 B.n450 B.n449 585
R445 B.n448 B.n440 585
R446 B.n626 B.n440 585
R447 B.n630 B.n393 585
R448 B.n393 B.n392 585
R449 B.n632 B.n631 585
R450 B.n633 B.n632 585
R451 B.n387 B.n386 585
R452 B.n388 B.n387 585
R453 B.n641 B.n640 585
R454 B.n640 B.n639 585
R455 B.n642 B.n385 585
R456 B.n385 B.n384 585
R457 B.n644 B.n643 585
R458 B.n645 B.n644 585
R459 B.n379 B.n378 585
R460 B.n380 B.n379 585
R461 B.n653 B.n652 585
R462 B.n652 B.n651 585
R463 B.n654 B.n377 585
R464 B.n377 B.n376 585
R465 B.n656 B.n655 585
R466 B.n657 B.n656 585
R467 B.n371 B.n370 585
R468 B.n372 B.n371 585
R469 B.n665 B.n664 585
R470 B.n664 B.n663 585
R471 B.n666 B.n369 585
R472 B.n369 B.n368 585
R473 B.n668 B.n667 585
R474 B.n669 B.n668 585
R475 B.n363 B.n362 585
R476 B.n364 B.n363 585
R477 B.n677 B.n676 585
R478 B.n676 B.n675 585
R479 B.n678 B.n361 585
R480 B.n361 B.n360 585
R481 B.n680 B.n679 585
R482 B.n681 B.n680 585
R483 B.n355 B.n354 585
R484 B.n356 B.n355 585
R485 B.n689 B.n688 585
R486 B.n688 B.n687 585
R487 B.n690 B.n353 585
R488 B.n353 B.n352 585
R489 B.n692 B.n691 585
R490 B.n693 B.n692 585
R491 B.n347 B.n346 585
R492 B.n348 B.n347 585
R493 B.n701 B.n700 585
R494 B.n700 B.n699 585
R495 B.n702 B.n345 585
R496 B.n345 B.n344 585
R497 B.n704 B.n703 585
R498 B.n705 B.n704 585
R499 B.n339 B.n338 585
R500 B.n340 B.n339 585
R501 B.n714 B.n713 585
R502 B.n713 B.n712 585
R503 B.n715 B.n337 585
R504 B.n711 B.n337 585
R505 B.n717 B.n716 585
R506 B.n718 B.n717 585
R507 B.n332 B.n331 585
R508 B.n333 B.n332 585
R509 B.n726 B.n725 585
R510 B.n725 B.n724 585
R511 B.n727 B.n330 585
R512 B.n330 B.n329 585
R513 B.n729 B.n728 585
R514 B.n730 B.n729 585
R515 B.n324 B.n323 585
R516 B.n325 B.n324 585
R517 B.n738 B.n737 585
R518 B.n737 B.n736 585
R519 B.n739 B.n322 585
R520 B.n322 B.n321 585
R521 B.n741 B.n740 585
R522 B.n742 B.n741 585
R523 B.n316 B.n315 585
R524 B.n317 B.n316 585
R525 B.n751 B.n750 585
R526 B.n750 B.n749 585
R527 B.n752 B.n314 585
R528 B.n314 B.n313 585
R529 B.n754 B.n753 585
R530 B.n755 B.n754 585
R531 B.n2 B.n0 585
R532 B.n4 B.n2 585
R533 B.n3 B.n1 585
R534 B.n904 B.n3 585
R535 B.n902 B.n901 585
R536 B.n903 B.n902 585
R537 B.n900 B.n9 585
R538 B.n9 B.n8 585
R539 B.n899 B.n898 585
R540 B.n898 B.n897 585
R541 B.n11 B.n10 585
R542 B.n896 B.n11 585
R543 B.n894 B.n893 585
R544 B.n895 B.n894 585
R545 B.n892 B.n16 585
R546 B.n16 B.n15 585
R547 B.n891 B.n890 585
R548 B.n890 B.n889 585
R549 B.n18 B.n17 585
R550 B.n888 B.n18 585
R551 B.n886 B.n885 585
R552 B.n887 B.n886 585
R553 B.n884 B.n23 585
R554 B.n23 B.n22 585
R555 B.n883 B.n882 585
R556 B.n882 B.n881 585
R557 B.n25 B.n24 585
R558 B.n880 B.n25 585
R559 B.n878 B.n877 585
R560 B.n879 B.n878 585
R561 B.n876 B.n29 585
R562 B.n32 B.n29 585
R563 B.n875 B.n874 585
R564 B.n874 B.n873 585
R565 B.n31 B.n30 585
R566 B.n872 B.n31 585
R567 B.n870 B.n869 585
R568 B.n871 B.n870 585
R569 B.n868 B.n37 585
R570 B.n37 B.n36 585
R571 B.n867 B.n866 585
R572 B.n866 B.n865 585
R573 B.n39 B.n38 585
R574 B.n864 B.n39 585
R575 B.n862 B.n861 585
R576 B.n863 B.n862 585
R577 B.n860 B.n44 585
R578 B.n44 B.n43 585
R579 B.n859 B.n858 585
R580 B.n858 B.n857 585
R581 B.n46 B.n45 585
R582 B.n856 B.n46 585
R583 B.n854 B.n853 585
R584 B.n855 B.n854 585
R585 B.n852 B.n51 585
R586 B.n51 B.n50 585
R587 B.n851 B.n850 585
R588 B.n850 B.n849 585
R589 B.n53 B.n52 585
R590 B.n848 B.n53 585
R591 B.n846 B.n845 585
R592 B.n847 B.n846 585
R593 B.n844 B.n58 585
R594 B.n58 B.n57 585
R595 B.n843 B.n842 585
R596 B.n842 B.n841 585
R597 B.n60 B.n59 585
R598 B.n840 B.n60 585
R599 B.n838 B.n837 585
R600 B.n839 B.n838 585
R601 B.n836 B.n65 585
R602 B.n65 B.n64 585
R603 B.n835 B.n834 585
R604 B.n834 B.n833 585
R605 B.n67 B.n66 585
R606 B.n832 B.n67 585
R607 B.n830 B.n829 585
R608 B.n831 B.n830 585
R609 B.n828 B.n72 585
R610 B.n72 B.n71 585
R611 B.n827 B.n826 585
R612 B.n826 B.n825 585
R613 B.n74 B.n73 585
R614 B.n824 B.n74 585
R615 B.n822 B.n821 585
R616 B.n823 B.n822 585
R617 B.n820 B.n79 585
R618 B.n79 B.n78 585
R619 B.n907 B.n906 585
R620 B.n906 B.n905 585
R621 B.n628 B.n393 492.5
R622 B.n818 B.n79 492.5
R623 B.n440 B.n391 492.5
R624 B.n814 B.n127 492.5
R625 B.n445 B.t17 316.101
R626 B.n442 B.t10 316.101
R627 B.n130 B.t6 316.101
R628 B.n128 B.t14 316.101
R629 B.n816 B.n815 256.663
R630 B.n816 B.n125 256.663
R631 B.n816 B.n124 256.663
R632 B.n816 B.n123 256.663
R633 B.n816 B.n122 256.663
R634 B.n816 B.n121 256.663
R635 B.n816 B.n120 256.663
R636 B.n816 B.n119 256.663
R637 B.n816 B.n118 256.663
R638 B.n816 B.n117 256.663
R639 B.n816 B.n116 256.663
R640 B.n816 B.n115 256.663
R641 B.n816 B.n114 256.663
R642 B.n816 B.n113 256.663
R643 B.n816 B.n112 256.663
R644 B.n816 B.n111 256.663
R645 B.n816 B.n110 256.663
R646 B.n816 B.n109 256.663
R647 B.n816 B.n108 256.663
R648 B.n816 B.n107 256.663
R649 B.n816 B.n106 256.663
R650 B.n816 B.n105 256.663
R651 B.n816 B.n104 256.663
R652 B.n816 B.n103 256.663
R653 B.n816 B.n102 256.663
R654 B.n816 B.n101 256.663
R655 B.n816 B.n100 256.663
R656 B.n816 B.n99 256.663
R657 B.n816 B.n98 256.663
R658 B.n816 B.n97 256.663
R659 B.n816 B.n96 256.663
R660 B.n816 B.n95 256.663
R661 B.n816 B.n94 256.663
R662 B.n816 B.n93 256.663
R663 B.n816 B.n92 256.663
R664 B.n816 B.n91 256.663
R665 B.n816 B.n90 256.663
R666 B.n816 B.n89 256.663
R667 B.n816 B.n88 256.663
R668 B.n816 B.n87 256.663
R669 B.n816 B.n86 256.663
R670 B.n816 B.n85 256.663
R671 B.n816 B.n84 256.663
R672 B.n816 B.n83 256.663
R673 B.n816 B.n82 256.663
R674 B.n817 B.n816 256.663
R675 B.n627 B.n626 256.663
R676 B.n626 B.n396 256.663
R677 B.n626 B.n397 256.663
R678 B.n626 B.n398 256.663
R679 B.n626 B.n399 256.663
R680 B.n626 B.n400 256.663
R681 B.n626 B.n401 256.663
R682 B.n626 B.n402 256.663
R683 B.n626 B.n403 256.663
R684 B.n626 B.n404 256.663
R685 B.n626 B.n405 256.663
R686 B.n626 B.n406 256.663
R687 B.n626 B.n407 256.663
R688 B.n626 B.n408 256.663
R689 B.n626 B.n409 256.663
R690 B.n626 B.n410 256.663
R691 B.n626 B.n411 256.663
R692 B.n626 B.n412 256.663
R693 B.n626 B.n413 256.663
R694 B.n626 B.n414 256.663
R695 B.n626 B.n415 256.663
R696 B.n626 B.n416 256.663
R697 B.n626 B.n417 256.663
R698 B.n626 B.n418 256.663
R699 B.n626 B.n419 256.663
R700 B.n626 B.n420 256.663
R701 B.n626 B.n421 256.663
R702 B.n626 B.n422 256.663
R703 B.n626 B.n423 256.663
R704 B.n626 B.n424 256.663
R705 B.n626 B.n425 256.663
R706 B.n626 B.n426 256.663
R707 B.n626 B.n427 256.663
R708 B.n626 B.n428 256.663
R709 B.n626 B.n429 256.663
R710 B.n626 B.n430 256.663
R711 B.n626 B.n431 256.663
R712 B.n626 B.n432 256.663
R713 B.n626 B.n433 256.663
R714 B.n626 B.n434 256.663
R715 B.n626 B.n435 256.663
R716 B.n626 B.n436 256.663
R717 B.n626 B.n437 256.663
R718 B.n626 B.n438 256.663
R719 B.n626 B.n439 256.663
R720 B.n632 B.n393 163.367
R721 B.n632 B.n387 163.367
R722 B.n640 B.n387 163.367
R723 B.n640 B.n385 163.367
R724 B.n644 B.n385 163.367
R725 B.n644 B.n379 163.367
R726 B.n652 B.n379 163.367
R727 B.n652 B.n377 163.367
R728 B.n656 B.n377 163.367
R729 B.n656 B.n371 163.367
R730 B.n664 B.n371 163.367
R731 B.n664 B.n369 163.367
R732 B.n668 B.n369 163.367
R733 B.n668 B.n363 163.367
R734 B.n676 B.n363 163.367
R735 B.n676 B.n361 163.367
R736 B.n680 B.n361 163.367
R737 B.n680 B.n355 163.367
R738 B.n688 B.n355 163.367
R739 B.n688 B.n353 163.367
R740 B.n692 B.n353 163.367
R741 B.n692 B.n347 163.367
R742 B.n700 B.n347 163.367
R743 B.n700 B.n345 163.367
R744 B.n704 B.n345 163.367
R745 B.n704 B.n339 163.367
R746 B.n713 B.n339 163.367
R747 B.n713 B.n337 163.367
R748 B.n717 B.n337 163.367
R749 B.n717 B.n332 163.367
R750 B.n725 B.n332 163.367
R751 B.n725 B.n330 163.367
R752 B.n729 B.n330 163.367
R753 B.n729 B.n324 163.367
R754 B.n737 B.n324 163.367
R755 B.n737 B.n322 163.367
R756 B.n741 B.n322 163.367
R757 B.n741 B.n316 163.367
R758 B.n750 B.n316 163.367
R759 B.n750 B.n314 163.367
R760 B.n754 B.n314 163.367
R761 B.n754 B.n2 163.367
R762 B.n906 B.n2 163.367
R763 B.n906 B.n3 163.367
R764 B.n902 B.n3 163.367
R765 B.n902 B.n9 163.367
R766 B.n898 B.n9 163.367
R767 B.n898 B.n11 163.367
R768 B.n894 B.n11 163.367
R769 B.n894 B.n16 163.367
R770 B.n890 B.n16 163.367
R771 B.n890 B.n18 163.367
R772 B.n886 B.n18 163.367
R773 B.n886 B.n23 163.367
R774 B.n882 B.n23 163.367
R775 B.n882 B.n25 163.367
R776 B.n878 B.n25 163.367
R777 B.n878 B.n29 163.367
R778 B.n874 B.n29 163.367
R779 B.n874 B.n31 163.367
R780 B.n870 B.n31 163.367
R781 B.n870 B.n37 163.367
R782 B.n866 B.n37 163.367
R783 B.n866 B.n39 163.367
R784 B.n862 B.n39 163.367
R785 B.n862 B.n44 163.367
R786 B.n858 B.n44 163.367
R787 B.n858 B.n46 163.367
R788 B.n854 B.n46 163.367
R789 B.n854 B.n51 163.367
R790 B.n850 B.n51 163.367
R791 B.n850 B.n53 163.367
R792 B.n846 B.n53 163.367
R793 B.n846 B.n58 163.367
R794 B.n842 B.n58 163.367
R795 B.n842 B.n60 163.367
R796 B.n838 B.n60 163.367
R797 B.n838 B.n65 163.367
R798 B.n834 B.n65 163.367
R799 B.n834 B.n67 163.367
R800 B.n830 B.n67 163.367
R801 B.n830 B.n72 163.367
R802 B.n826 B.n72 163.367
R803 B.n826 B.n74 163.367
R804 B.n822 B.n74 163.367
R805 B.n822 B.n79 163.367
R806 B.n625 B.n395 163.367
R807 B.n625 B.n441 163.367
R808 B.n621 B.n620 163.367
R809 B.n617 B.n616 163.367
R810 B.n613 B.n612 163.367
R811 B.n609 B.n608 163.367
R812 B.n605 B.n604 163.367
R813 B.n601 B.n600 163.367
R814 B.n597 B.n596 163.367
R815 B.n593 B.n592 163.367
R816 B.n589 B.n588 163.367
R817 B.n585 B.n584 163.367
R818 B.n581 B.n580 163.367
R819 B.n577 B.n576 163.367
R820 B.n573 B.n572 163.367
R821 B.n569 B.n568 163.367
R822 B.n565 B.n564 163.367
R823 B.n561 B.n560 163.367
R824 B.n557 B.n556 163.367
R825 B.n553 B.n552 163.367
R826 B.n549 B.n548 163.367
R827 B.n545 B.n544 163.367
R828 B.n541 B.n540 163.367
R829 B.n537 B.n536 163.367
R830 B.n533 B.n532 163.367
R831 B.n529 B.n528 163.367
R832 B.n525 B.n524 163.367
R833 B.n521 B.n520 163.367
R834 B.n517 B.n516 163.367
R835 B.n513 B.n512 163.367
R836 B.n509 B.n508 163.367
R837 B.n505 B.n504 163.367
R838 B.n501 B.n500 163.367
R839 B.n497 B.n496 163.367
R840 B.n493 B.n492 163.367
R841 B.n489 B.n488 163.367
R842 B.n485 B.n484 163.367
R843 B.n481 B.n480 163.367
R844 B.n477 B.n476 163.367
R845 B.n473 B.n472 163.367
R846 B.n469 B.n468 163.367
R847 B.n465 B.n464 163.367
R848 B.n461 B.n460 163.367
R849 B.n457 B.n456 163.367
R850 B.n453 B.n452 163.367
R851 B.n449 B.n440 163.367
R852 B.n634 B.n391 163.367
R853 B.n634 B.n389 163.367
R854 B.n638 B.n389 163.367
R855 B.n638 B.n383 163.367
R856 B.n646 B.n383 163.367
R857 B.n646 B.n381 163.367
R858 B.n650 B.n381 163.367
R859 B.n650 B.n375 163.367
R860 B.n658 B.n375 163.367
R861 B.n658 B.n373 163.367
R862 B.n662 B.n373 163.367
R863 B.n662 B.n367 163.367
R864 B.n670 B.n367 163.367
R865 B.n670 B.n365 163.367
R866 B.n674 B.n365 163.367
R867 B.n674 B.n359 163.367
R868 B.n682 B.n359 163.367
R869 B.n682 B.n357 163.367
R870 B.n686 B.n357 163.367
R871 B.n686 B.n351 163.367
R872 B.n694 B.n351 163.367
R873 B.n694 B.n349 163.367
R874 B.n698 B.n349 163.367
R875 B.n698 B.n343 163.367
R876 B.n706 B.n343 163.367
R877 B.n706 B.n341 163.367
R878 B.n710 B.n341 163.367
R879 B.n710 B.n336 163.367
R880 B.n719 B.n336 163.367
R881 B.n719 B.n334 163.367
R882 B.n723 B.n334 163.367
R883 B.n723 B.n328 163.367
R884 B.n731 B.n328 163.367
R885 B.n731 B.n326 163.367
R886 B.n735 B.n326 163.367
R887 B.n735 B.n320 163.367
R888 B.n743 B.n320 163.367
R889 B.n743 B.n318 163.367
R890 B.n748 B.n318 163.367
R891 B.n748 B.n312 163.367
R892 B.n756 B.n312 163.367
R893 B.n757 B.n756 163.367
R894 B.n757 B.n5 163.367
R895 B.n6 B.n5 163.367
R896 B.n7 B.n6 163.367
R897 B.n762 B.n7 163.367
R898 B.n762 B.n12 163.367
R899 B.n13 B.n12 163.367
R900 B.n14 B.n13 163.367
R901 B.n767 B.n14 163.367
R902 B.n767 B.n19 163.367
R903 B.n20 B.n19 163.367
R904 B.n21 B.n20 163.367
R905 B.n772 B.n21 163.367
R906 B.n772 B.n26 163.367
R907 B.n27 B.n26 163.367
R908 B.n28 B.n27 163.367
R909 B.n777 B.n28 163.367
R910 B.n777 B.n33 163.367
R911 B.n34 B.n33 163.367
R912 B.n35 B.n34 163.367
R913 B.n782 B.n35 163.367
R914 B.n782 B.n40 163.367
R915 B.n41 B.n40 163.367
R916 B.n42 B.n41 163.367
R917 B.n787 B.n42 163.367
R918 B.n787 B.n47 163.367
R919 B.n48 B.n47 163.367
R920 B.n49 B.n48 163.367
R921 B.n792 B.n49 163.367
R922 B.n792 B.n54 163.367
R923 B.n55 B.n54 163.367
R924 B.n56 B.n55 163.367
R925 B.n797 B.n56 163.367
R926 B.n797 B.n61 163.367
R927 B.n62 B.n61 163.367
R928 B.n63 B.n62 163.367
R929 B.n802 B.n63 163.367
R930 B.n802 B.n68 163.367
R931 B.n69 B.n68 163.367
R932 B.n70 B.n69 163.367
R933 B.n807 B.n70 163.367
R934 B.n807 B.n75 163.367
R935 B.n76 B.n75 163.367
R936 B.n77 B.n76 163.367
R937 B.n127 B.n77 163.367
R938 B.n132 B.n81 163.367
R939 B.n136 B.n135 163.367
R940 B.n140 B.n139 163.367
R941 B.n144 B.n143 163.367
R942 B.n148 B.n147 163.367
R943 B.n152 B.n151 163.367
R944 B.n156 B.n155 163.367
R945 B.n160 B.n159 163.367
R946 B.n164 B.n163 163.367
R947 B.n168 B.n167 163.367
R948 B.n172 B.n171 163.367
R949 B.n176 B.n175 163.367
R950 B.n180 B.n179 163.367
R951 B.n184 B.n183 163.367
R952 B.n188 B.n187 163.367
R953 B.n192 B.n191 163.367
R954 B.n196 B.n195 163.367
R955 B.n200 B.n199 163.367
R956 B.n204 B.n203 163.367
R957 B.n208 B.n207 163.367
R958 B.n213 B.n212 163.367
R959 B.n217 B.n216 163.367
R960 B.n221 B.n220 163.367
R961 B.n225 B.n224 163.367
R962 B.n229 B.n228 163.367
R963 B.n234 B.n233 163.367
R964 B.n238 B.n237 163.367
R965 B.n242 B.n241 163.367
R966 B.n246 B.n245 163.367
R967 B.n250 B.n249 163.367
R968 B.n254 B.n253 163.367
R969 B.n258 B.n257 163.367
R970 B.n262 B.n261 163.367
R971 B.n266 B.n265 163.367
R972 B.n270 B.n269 163.367
R973 B.n274 B.n273 163.367
R974 B.n278 B.n277 163.367
R975 B.n282 B.n281 163.367
R976 B.n286 B.n285 163.367
R977 B.n290 B.n289 163.367
R978 B.n294 B.n293 163.367
R979 B.n298 B.n297 163.367
R980 B.n302 B.n301 163.367
R981 B.n306 B.n305 163.367
R982 B.n308 B.n126 163.367
R983 B.n445 B.t19 130.649
R984 B.n128 B.t15 130.649
R985 B.n442 B.t13 130.635
R986 B.n130 B.t8 130.635
R987 B.n626 B.n392 81.6725
R988 B.n816 B.n78 81.6725
R989 B.n446 B.t18 73.0495
R990 B.n129 B.t16 73.0495
R991 B.n443 B.t12 73.0347
R992 B.n131 B.t9 73.0347
R993 B.n628 B.n627 71.676
R994 B.n441 B.n396 71.676
R995 B.n620 B.n397 71.676
R996 B.n616 B.n398 71.676
R997 B.n612 B.n399 71.676
R998 B.n608 B.n400 71.676
R999 B.n604 B.n401 71.676
R1000 B.n600 B.n402 71.676
R1001 B.n596 B.n403 71.676
R1002 B.n592 B.n404 71.676
R1003 B.n588 B.n405 71.676
R1004 B.n584 B.n406 71.676
R1005 B.n580 B.n407 71.676
R1006 B.n576 B.n408 71.676
R1007 B.n572 B.n409 71.676
R1008 B.n568 B.n410 71.676
R1009 B.n564 B.n411 71.676
R1010 B.n560 B.n412 71.676
R1011 B.n556 B.n413 71.676
R1012 B.n552 B.n414 71.676
R1013 B.n548 B.n415 71.676
R1014 B.n544 B.n416 71.676
R1015 B.n540 B.n417 71.676
R1016 B.n536 B.n418 71.676
R1017 B.n532 B.n419 71.676
R1018 B.n528 B.n420 71.676
R1019 B.n524 B.n421 71.676
R1020 B.n520 B.n422 71.676
R1021 B.n516 B.n423 71.676
R1022 B.n512 B.n424 71.676
R1023 B.n508 B.n425 71.676
R1024 B.n504 B.n426 71.676
R1025 B.n500 B.n427 71.676
R1026 B.n496 B.n428 71.676
R1027 B.n492 B.n429 71.676
R1028 B.n488 B.n430 71.676
R1029 B.n484 B.n431 71.676
R1030 B.n480 B.n432 71.676
R1031 B.n476 B.n433 71.676
R1032 B.n472 B.n434 71.676
R1033 B.n468 B.n435 71.676
R1034 B.n464 B.n436 71.676
R1035 B.n460 B.n437 71.676
R1036 B.n456 B.n438 71.676
R1037 B.n452 B.n439 71.676
R1038 B.n818 B.n817 71.676
R1039 B.n132 B.n82 71.676
R1040 B.n136 B.n83 71.676
R1041 B.n140 B.n84 71.676
R1042 B.n144 B.n85 71.676
R1043 B.n148 B.n86 71.676
R1044 B.n152 B.n87 71.676
R1045 B.n156 B.n88 71.676
R1046 B.n160 B.n89 71.676
R1047 B.n164 B.n90 71.676
R1048 B.n168 B.n91 71.676
R1049 B.n172 B.n92 71.676
R1050 B.n176 B.n93 71.676
R1051 B.n180 B.n94 71.676
R1052 B.n184 B.n95 71.676
R1053 B.n188 B.n96 71.676
R1054 B.n192 B.n97 71.676
R1055 B.n196 B.n98 71.676
R1056 B.n200 B.n99 71.676
R1057 B.n204 B.n100 71.676
R1058 B.n208 B.n101 71.676
R1059 B.n213 B.n102 71.676
R1060 B.n217 B.n103 71.676
R1061 B.n221 B.n104 71.676
R1062 B.n225 B.n105 71.676
R1063 B.n229 B.n106 71.676
R1064 B.n234 B.n107 71.676
R1065 B.n238 B.n108 71.676
R1066 B.n242 B.n109 71.676
R1067 B.n246 B.n110 71.676
R1068 B.n250 B.n111 71.676
R1069 B.n254 B.n112 71.676
R1070 B.n258 B.n113 71.676
R1071 B.n262 B.n114 71.676
R1072 B.n266 B.n115 71.676
R1073 B.n270 B.n116 71.676
R1074 B.n274 B.n117 71.676
R1075 B.n278 B.n118 71.676
R1076 B.n282 B.n119 71.676
R1077 B.n286 B.n120 71.676
R1078 B.n290 B.n121 71.676
R1079 B.n294 B.n122 71.676
R1080 B.n298 B.n123 71.676
R1081 B.n302 B.n124 71.676
R1082 B.n306 B.n125 71.676
R1083 B.n815 B.n126 71.676
R1084 B.n815 B.n814 71.676
R1085 B.n308 B.n125 71.676
R1086 B.n305 B.n124 71.676
R1087 B.n301 B.n123 71.676
R1088 B.n297 B.n122 71.676
R1089 B.n293 B.n121 71.676
R1090 B.n289 B.n120 71.676
R1091 B.n285 B.n119 71.676
R1092 B.n281 B.n118 71.676
R1093 B.n277 B.n117 71.676
R1094 B.n273 B.n116 71.676
R1095 B.n269 B.n115 71.676
R1096 B.n265 B.n114 71.676
R1097 B.n261 B.n113 71.676
R1098 B.n257 B.n112 71.676
R1099 B.n253 B.n111 71.676
R1100 B.n249 B.n110 71.676
R1101 B.n245 B.n109 71.676
R1102 B.n241 B.n108 71.676
R1103 B.n237 B.n107 71.676
R1104 B.n233 B.n106 71.676
R1105 B.n228 B.n105 71.676
R1106 B.n224 B.n104 71.676
R1107 B.n220 B.n103 71.676
R1108 B.n216 B.n102 71.676
R1109 B.n212 B.n101 71.676
R1110 B.n207 B.n100 71.676
R1111 B.n203 B.n99 71.676
R1112 B.n199 B.n98 71.676
R1113 B.n195 B.n97 71.676
R1114 B.n191 B.n96 71.676
R1115 B.n187 B.n95 71.676
R1116 B.n183 B.n94 71.676
R1117 B.n179 B.n93 71.676
R1118 B.n175 B.n92 71.676
R1119 B.n171 B.n91 71.676
R1120 B.n167 B.n90 71.676
R1121 B.n163 B.n89 71.676
R1122 B.n159 B.n88 71.676
R1123 B.n155 B.n87 71.676
R1124 B.n151 B.n86 71.676
R1125 B.n147 B.n85 71.676
R1126 B.n143 B.n84 71.676
R1127 B.n139 B.n83 71.676
R1128 B.n135 B.n82 71.676
R1129 B.n817 B.n81 71.676
R1130 B.n627 B.n395 71.676
R1131 B.n621 B.n396 71.676
R1132 B.n617 B.n397 71.676
R1133 B.n613 B.n398 71.676
R1134 B.n609 B.n399 71.676
R1135 B.n605 B.n400 71.676
R1136 B.n601 B.n401 71.676
R1137 B.n597 B.n402 71.676
R1138 B.n593 B.n403 71.676
R1139 B.n589 B.n404 71.676
R1140 B.n585 B.n405 71.676
R1141 B.n581 B.n406 71.676
R1142 B.n577 B.n407 71.676
R1143 B.n573 B.n408 71.676
R1144 B.n569 B.n409 71.676
R1145 B.n565 B.n410 71.676
R1146 B.n561 B.n411 71.676
R1147 B.n557 B.n412 71.676
R1148 B.n553 B.n413 71.676
R1149 B.n549 B.n414 71.676
R1150 B.n545 B.n415 71.676
R1151 B.n541 B.n416 71.676
R1152 B.n537 B.n417 71.676
R1153 B.n533 B.n418 71.676
R1154 B.n529 B.n419 71.676
R1155 B.n525 B.n420 71.676
R1156 B.n521 B.n421 71.676
R1157 B.n517 B.n422 71.676
R1158 B.n513 B.n423 71.676
R1159 B.n509 B.n424 71.676
R1160 B.n505 B.n425 71.676
R1161 B.n501 B.n426 71.676
R1162 B.n497 B.n427 71.676
R1163 B.n493 B.n428 71.676
R1164 B.n489 B.n429 71.676
R1165 B.n485 B.n430 71.676
R1166 B.n481 B.n431 71.676
R1167 B.n477 B.n432 71.676
R1168 B.n473 B.n433 71.676
R1169 B.n469 B.n434 71.676
R1170 B.n465 B.n435 71.676
R1171 B.n461 B.n436 71.676
R1172 B.n457 B.n437 71.676
R1173 B.n453 B.n438 71.676
R1174 B.n449 B.n439 71.676
R1175 B.n447 B.n446 59.5399
R1176 B.n444 B.n443 59.5399
R1177 B.n210 B.n131 59.5399
R1178 B.n231 B.n129 59.5399
R1179 B.n446 B.n445 57.6005
R1180 B.n443 B.n442 57.6005
R1181 B.n131 B.n130 57.6005
R1182 B.n129 B.n128 57.6005
R1183 B.n633 B.n392 43.7304
R1184 B.n633 B.n388 43.7304
R1185 B.n639 B.n388 43.7304
R1186 B.n639 B.n384 43.7304
R1187 B.n645 B.n384 43.7304
R1188 B.n645 B.n380 43.7304
R1189 B.n651 B.n380 43.7304
R1190 B.n657 B.n376 43.7304
R1191 B.n657 B.n372 43.7304
R1192 B.n663 B.n372 43.7304
R1193 B.n663 B.n368 43.7304
R1194 B.n669 B.n368 43.7304
R1195 B.n669 B.n364 43.7304
R1196 B.n675 B.n364 43.7304
R1197 B.n675 B.n360 43.7304
R1198 B.n681 B.n360 43.7304
R1199 B.n681 B.n356 43.7304
R1200 B.n687 B.n356 43.7304
R1201 B.n693 B.n352 43.7304
R1202 B.n693 B.n348 43.7304
R1203 B.n699 B.n348 43.7304
R1204 B.n699 B.n344 43.7304
R1205 B.n705 B.n344 43.7304
R1206 B.n705 B.n340 43.7304
R1207 B.n712 B.n340 43.7304
R1208 B.n712 B.n711 43.7304
R1209 B.n718 B.n333 43.7304
R1210 B.n724 B.n333 43.7304
R1211 B.n724 B.n329 43.7304
R1212 B.n730 B.n329 43.7304
R1213 B.n730 B.n325 43.7304
R1214 B.n736 B.n325 43.7304
R1215 B.n736 B.n321 43.7304
R1216 B.n742 B.n321 43.7304
R1217 B.n749 B.n317 43.7304
R1218 B.n749 B.n313 43.7304
R1219 B.n755 B.n313 43.7304
R1220 B.n755 B.n4 43.7304
R1221 B.n905 B.n4 43.7304
R1222 B.n905 B.n904 43.7304
R1223 B.n904 B.n903 43.7304
R1224 B.n903 B.n8 43.7304
R1225 B.n897 B.n8 43.7304
R1226 B.n897 B.n896 43.7304
R1227 B.n895 B.n15 43.7304
R1228 B.n889 B.n15 43.7304
R1229 B.n889 B.n888 43.7304
R1230 B.n888 B.n887 43.7304
R1231 B.n887 B.n22 43.7304
R1232 B.n881 B.n22 43.7304
R1233 B.n881 B.n880 43.7304
R1234 B.n880 B.n879 43.7304
R1235 B.n873 B.n32 43.7304
R1236 B.n873 B.n872 43.7304
R1237 B.n872 B.n871 43.7304
R1238 B.n871 B.n36 43.7304
R1239 B.n865 B.n36 43.7304
R1240 B.n865 B.n864 43.7304
R1241 B.n864 B.n863 43.7304
R1242 B.n863 B.n43 43.7304
R1243 B.n857 B.n856 43.7304
R1244 B.n856 B.n855 43.7304
R1245 B.n855 B.n50 43.7304
R1246 B.n849 B.n50 43.7304
R1247 B.n849 B.n848 43.7304
R1248 B.n848 B.n847 43.7304
R1249 B.n847 B.n57 43.7304
R1250 B.n841 B.n57 43.7304
R1251 B.n841 B.n840 43.7304
R1252 B.n840 B.n839 43.7304
R1253 B.n839 B.n64 43.7304
R1254 B.n833 B.n832 43.7304
R1255 B.n832 B.n831 43.7304
R1256 B.n831 B.n71 43.7304
R1257 B.n825 B.n71 43.7304
R1258 B.n825 B.n824 43.7304
R1259 B.n824 B.n823 43.7304
R1260 B.n823 B.n78 43.7304
R1261 B.t3 B.n317 42.4442
R1262 B.n896 B.t1 42.4442
R1263 B.n820 B.n819 32.0005
R1264 B.n813 B.n812 32.0005
R1265 B.n448 B.n390 32.0005
R1266 B.n630 B.n629 32.0005
R1267 B.n718 B.t5 30.8687
R1268 B.n879 B.t2 30.8687
R1269 B.n651 B.t11 27.0101
R1270 B.n833 B.t7 27.0101
R1271 B.n687 B.t0 24.4378
R1272 B.n857 B.t4 24.4378
R1273 B.t0 B.n352 19.2931
R1274 B.t4 B.n43 19.2931
R1275 B B.n907 18.0485
R1276 B.t11 B.n376 16.7208
R1277 B.t7 B.n64 16.7208
R1278 B.n711 B.t5 12.8622
R1279 B.n32 B.t2 12.8622
R1280 B.n819 B.n80 10.6151
R1281 B.n133 B.n80 10.6151
R1282 B.n134 B.n133 10.6151
R1283 B.n137 B.n134 10.6151
R1284 B.n138 B.n137 10.6151
R1285 B.n141 B.n138 10.6151
R1286 B.n142 B.n141 10.6151
R1287 B.n145 B.n142 10.6151
R1288 B.n146 B.n145 10.6151
R1289 B.n149 B.n146 10.6151
R1290 B.n150 B.n149 10.6151
R1291 B.n153 B.n150 10.6151
R1292 B.n154 B.n153 10.6151
R1293 B.n157 B.n154 10.6151
R1294 B.n158 B.n157 10.6151
R1295 B.n161 B.n158 10.6151
R1296 B.n162 B.n161 10.6151
R1297 B.n165 B.n162 10.6151
R1298 B.n166 B.n165 10.6151
R1299 B.n169 B.n166 10.6151
R1300 B.n170 B.n169 10.6151
R1301 B.n173 B.n170 10.6151
R1302 B.n174 B.n173 10.6151
R1303 B.n177 B.n174 10.6151
R1304 B.n178 B.n177 10.6151
R1305 B.n181 B.n178 10.6151
R1306 B.n182 B.n181 10.6151
R1307 B.n185 B.n182 10.6151
R1308 B.n186 B.n185 10.6151
R1309 B.n189 B.n186 10.6151
R1310 B.n190 B.n189 10.6151
R1311 B.n193 B.n190 10.6151
R1312 B.n194 B.n193 10.6151
R1313 B.n197 B.n194 10.6151
R1314 B.n198 B.n197 10.6151
R1315 B.n201 B.n198 10.6151
R1316 B.n202 B.n201 10.6151
R1317 B.n205 B.n202 10.6151
R1318 B.n206 B.n205 10.6151
R1319 B.n209 B.n206 10.6151
R1320 B.n214 B.n211 10.6151
R1321 B.n215 B.n214 10.6151
R1322 B.n218 B.n215 10.6151
R1323 B.n219 B.n218 10.6151
R1324 B.n222 B.n219 10.6151
R1325 B.n223 B.n222 10.6151
R1326 B.n226 B.n223 10.6151
R1327 B.n227 B.n226 10.6151
R1328 B.n230 B.n227 10.6151
R1329 B.n235 B.n232 10.6151
R1330 B.n236 B.n235 10.6151
R1331 B.n239 B.n236 10.6151
R1332 B.n240 B.n239 10.6151
R1333 B.n243 B.n240 10.6151
R1334 B.n244 B.n243 10.6151
R1335 B.n247 B.n244 10.6151
R1336 B.n248 B.n247 10.6151
R1337 B.n251 B.n248 10.6151
R1338 B.n252 B.n251 10.6151
R1339 B.n255 B.n252 10.6151
R1340 B.n256 B.n255 10.6151
R1341 B.n259 B.n256 10.6151
R1342 B.n260 B.n259 10.6151
R1343 B.n263 B.n260 10.6151
R1344 B.n264 B.n263 10.6151
R1345 B.n267 B.n264 10.6151
R1346 B.n268 B.n267 10.6151
R1347 B.n271 B.n268 10.6151
R1348 B.n272 B.n271 10.6151
R1349 B.n275 B.n272 10.6151
R1350 B.n276 B.n275 10.6151
R1351 B.n279 B.n276 10.6151
R1352 B.n280 B.n279 10.6151
R1353 B.n283 B.n280 10.6151
R1354 B.n284 B.n283 10.6151
R1355 B.n287 B.n284 10.6151
R1356 B.n288 B.n287 10.6151
R1357 B.n291 B.n288 10.6151
R1358 B.n292 B.n291 10.6151
R1359 B.n295 B.n292 10.6151
R1360 B.n296 B.n295 10.6151
R1361 B.n299 B.n296 10.6151
R1362 B.n300 B.n299 10.6151
R1363 B.n303 B.n300 10.6151
R1364 B.n304 B.n303 10.6151
R1365 B.n307 B.n304 10.6151
R1366 B.n309 B.n307 10.6151
R1367 B.n310 B.n309 10.6151
R1368 B.n813 B.n310 10.6151
R1369 B.n635 B.n390 10.6151
R1370 B.n636 B.n635 10.6151
R1371 B.n637 B.n636 10.6151
R1372 B.n637 B.n382 10.6151
R1373 B.n647 B.n382 10.6151
R1374 B.n648 B.n647 10.6151
R1375 B.n649 B.n648 10.6151
R1376 B.n649 B.n374 10.6151
R1377 B.n659 B.n374 10.6151
R1378 B.n660 B.n659 10.6151
R1379 B.n661 B.n660 10.6151
R1380 B.n661 B.n366 10.6151
R1381 B.n671 B.n366 10.6151
R1382 B.n672 B.n671 10.6151
R1383 B.n673 B.n672 10.6151
R1384 B.n673 B.n358 10.6151
R1385 B.n683 B.n358 10.6151
R1386 B.n684 B.n683 10.6151
R1387 B.n685 B.n684 10.6151
R1388 B.n685 B.n350 10.6151
R1389 B.n695 B.n350 10.6151
R1390 B.n696 B.n695 10.6151
R1391 B.n697 B.n696 10.6151
R1392 B.n697 B.n342 10.6151
R1393 B.n707 B.n342 10.6151
R1394 B.n708 B.n707 10.6151
R1395 B.n709 B.n708 10.6151
R1396 B.n709 B.n335 10.6151
R1397 B.n720 B.n335 10.6151
R1398 B.n721 B.n720 10.6151
R1399 B.n722 B.n721 10.6151
R1400 B.n722 B.n327 10.6151
R1401 B.n732 B.n327 10.6151
R1402 B.n733 B.n732 10.6151
R1403 B.n734 B.n733 10.6151
R1404 B.n734 B.n319 10.6151
R1405 B.n744 B.n319 10.6151
R1406 B.n745 B.n744 10.6151
R1407 B.n747 B.n745 10.6151
R1408 B.n747 B.n746 10.6151
R1409 B.n746 B.n311 10.6151
R1410 B.n758 B.n311 10.6151
R1411 B.n759 B.n758 10.6151
R1412 B.n760 B.n759 10.6151
R1413 B.n761 B.n760 10.6151
R1414 B.n763 B.n761 10.6151
R1415 B.n764 B.n763 10.6151
R1416 B.n765 B.n764 10.6151
R1417 B.n766 B.n765 10.6151
R1418 B.n768 B.n766 10.6151
R1419 B.n769 B.n768 10.6151
R1420 B.n770 B.n769 10.6151
R1421 B.n771 B.n770 10.6151
R1422 B.n773 B.n771 10.6151
R1423 B.n774 B.n773 10.6151
R1424 B.n775 B.n774 10.6151
R1425 B.n776 B.n775 10.6151
R1426 B.n778 B.n776 10.6151
R1427 B.n779 B.n778 10.6151
R1428 B.n780 B.n779 10.6151
R1429 B.n781 B.n780 10.6151
R1430 B.n783 B.n781 10.6151
R1431 B.n784 B.n783 10.6151
R1432 B.n785 B.n784 10.6151
R1433 B.n786 B.n785 10.6151
R1434 B.n788 B.n786 10.6151
R1435 B.n789 B.n788 10.6151
R1436 B.n790 B.n789 10.6151
R1437 B.n791 B.n790 10.6151
R1438 B.n793 B.n791 10.6151
R1439 B.n794 B.n793 10.6151
R1440 B.n795 B.n794 10.6151
R1441 B.n796 B.n795 10.6151
R1442 B.n798 B.n796 10.6151
R1443 B.n799 B.n798 10.6151
R1444 B.n800 B.n799 10.6151
R1445 B.n801 B.n800 10.6151
R1446 B.n803 B.n801 10.6151
R1447 B.n804 B.n803 10.6151
R1448 B.n805 B.n804 10.6151
R1449 B.n806 B.n805 10.6151
R1450 B.n808 B.n806 10.6151
R1451 B.n809 B.n808 10.6151
R1452 B.n810 B.n809 10.6151
R1453 B.n811 B.n810 10.6151
R1454 B.n812 B.n811 10.6151
R1455 B.n629 B.n394 10.6151
R1456 B.n624 B.n394 10.6151
R1457 B.n624 B.n623 10.6151
R1458 B.n623 B.n622 10.6151
R1459 B.n622 B.n619 10.6151
R1460 B.n619 B.n618 10.6151
R1461 B.n618 B.n615 10.6151
R1462 B.n615 B.n614 10.6151
R1463 B.n614 B.n611 10.6151
R1464 B.n611 B.n610 10.6151
R1465 B.n610 B.n607 10.6151
R1466 B.n607 B.n606 10.6151
R1467 B.n606 B.n603 10.6151
R1468 B.n603 B.n602 10.6151
R1469 B.n602 B.n599 10.6151
R1470 B.n599 B.n598 10.6151
R1471 B.n598 B.n595 10.6151
R1472 B.n595 B.n594 10.6151
R1473 B.n594 B.n591 10.6151
R1474 B.n591 B.n590 10.6151
R1475 B.n590 B.n587 10.6151
R1476 B.n587 B.n586 10.6151
R1477 B.n586 B.n583 10.6151
R1478 B.n583 B.n582 10.6151
R1479 B.n582 B.n579 10.6151
R1480 B.n579 B.n578 10.6151
R1481 B.n578 B.n575 10.6151
R1482 B.n575 B.n574 10.6151
R1483 B.n574 B.n571 10.6151
R1484 B.n571 B.n570 10.6151
R1485 B.n570 B.n567 10.6151
R1486 B.n567 B.n566 10.6151
R1487 B.n566 B.n563 10.6151
R1488 B.n563 B.n562 10.6151
R1489 B.n562 B.n559 10.6151
R1490 B.n559 B.n558 10.6151
R1491 B.n558 B.n555 10.6151
R1492 B.n555 B.n554 10.6151
R1493 B.n554 B.n551 10.6151
R1494 B.n551 B.n550 10.6151
R1495 B.n547 B.n546 10.6151
R1496 B.n546 B.n543 10.6151
R1497 B.n543 B.n542 10.6151
R1498 B.n542 B.n539 10.6151
R1499 B.n539 B.n538 10.6151
R1500 B.n538 B.n535 10.6151
R1501 B.n535 B.n534 10.6151
R1502 B.n534 B.n531 10.6151
R1503 B.n531 B.n530 10.6151
R1504 B.n527 B.n526 10.6151
R1505 B.n526 B.n523 10.6151
R1506 B.n523 B.n522 10.6151
R1507 B.n522 B.n519 10.6151
R1508 B.n519 B.n518 10.6151
R1509 B.n518 B.n515 10.6151
R1510 B.n515 B.n514 10.6151
R1511 B.n514 B.n511 10.6151
R1512 B.n511 B.n510 10.6151
R1513 B.n510 B.n507 10.6151
R1514 B.n507 B.n506 10.6151
R1515 B.n506 B.n503 10.6151
R1516 B.n503 B.n502 10.6151
R1517 B.n502 B.n499 10.6151
R1518 B.n499 B.n498 10.6151
R1519 B.n498 B.n495 10.6151
R1520 B.n495 B.n494 10.6151
R1521 B.n494 B.n491 10.6151
R1522 B.n491 B.n490 10.6151
R1523 B.n490 B.n487 10.6151
R1524 B.n487 B.n486 10.6151
R1525 B.n486 B.n483 10.6151
R1526 B.n483 B.n482 10.6151
R1527 B.n482 B.n479 10.6151
R1528 B.n479 B.n478 10.6151
R1529 B.n478 B.n475 10.6151
R1530 B.n475 B.n474 10.6151
R1531 B.n474 B.n471 10.6151
R1532 B.n471 B.n470 10.6151
R1533 B.n470 B.n467 10.6151
R1534 B.n467 B.n466 10.6151
R1535 B.n466 B.n463 10.6151
R1536 B.n463 B.n462 10.6151
R1537 B.n462 B.n459 10.6151
R1538 B.n459 B.n458 10.6151
R1539 B.n458 B.n455 10.6151
R1540 B.n455 B.n454 10.6151
R1541 B.n454 B.n451 10.6151
R1542 B.n451 B.n450 10.6151
R1543 B.n450 B.n448 10.6151
R1544 B.n631 B.n630 10.6151
R1545 B.n631 B.n386 10.6151
R1546 B.n641 B.n386 10.6151
R1547 B.n642 B.n641 10.6151
R1548 B.n643 B.n642 10.6151
R1549 B.n643 B.n378 10.6151
R1550 B.n653 B.n378 10.6151
R1551 B.n654 B.n653 10.6151
R1552 B.n655 B.n654 10.6151
R1553 B.n655 B.n370 10.6151
R1554 B.n665 B.n370 10.6151
R1555 B.n666 B.n665 10.6151
R1556 B.n667 B.n666 10.6151
R1557 B.n667 B.n362 10.6151
R1558 B.n677 B.n362 10.6151
R1559 B.n678 B.n677 10.6151
R1560 B.n679 B.n678 10.6151
R1561 B.n679 B.n354 10.6151
R1562 B.n689 B.n354 10.6151
R1563 B.n690 B.n689 10.6151
R1564 B.n691 B.n690 10.6151
R1565 B.n691 B.n346 10.6151
R1566 B.n701 B.n346 10.6151
R1567 B.n702 B.n701 10.6151
R1568 B.n703 B.n702 10.6151
R1569 B.n703 B.n338 10.6151
R1570 B.n714 B.n338 10.6151
R1571 B.n715 B.n714 10.6151
R1572 B.n716 B.n715 10.6151
R1573 B.n716 B.n331 10.6151
R1574 B.n726 B.n331 10.6151
R1575 B.n727 B.n726 10.6151
R1576 B.n728 B.n727 10.6151
R1577 B.n728 B.n323 10.6151
R1578 B.n738 B.n323 10.6151
R1579 B.n739 B.n738 10.6151
R1580 B.n740 B.n739 10.6151
R1581 B.n740 B.n315 10.6151
R1582 B.n751 B.n315 10.6151
R1583 B.n752 B.n751 10.6151
R1584 B.n753 B.n752 10.6151
R1585 B.n753 B.n0 10.6151
R1586 B.n901 B.n1 10.6151
R1587 B.n901 B.n900 10.6151
R1588 B.n900 B.n899 10.6151
R1589 B.n899 B.n10 10.6151
R1590 B.n893 B.n10 10.6151
R1591 B.n893 B.n892 10.6151
R1592 B.n892 B.n891 10.6151
R1593 B.n891 B.n17 10.6151
R1594 B.n885 B.n17 10.6151
R1595 B.n885 B.n884 10.6151
R1596 B.n884 B.n883 10.6151
R1597 B.n883 B.n24 10.6151
R1598 B.n877 B.n24 10.6151
R1599 B.n877 B.n876 10.6151
R1600 B.n876 B.n875 10.6151
R1601 B.n875 B.n30 10.6151
R1602 B.n869 B.n30 10.6151
R1603 B.n869 B.n868 10.6151
R1604 B.n868 B.n867 10.6151
R1605 B.n867 B.n38 10.6151
R1606 B.n861 B.n38 10.6151
R1607 B.n861 B.n860 10.6151
R1608 B.n860 B.n859 10.6151
R1609 B.n859 B.n45 10.6151
R1610 B.n853 B.n45 10.6151
R1611 B.n853 B.n852 10.6151
R1612 B.n852 B.n851 10.6151
R1613 B.n851 B.n52 10.6151
R1614 B.n845 B.n52 10.6151
R1615 B.n845 B.n844 10.6151
R1616 B.n844 B.n843 10.6151
R1617 B.n843 B.n59 10.6151
R1618 B.n837 B.n59 10.6151
R1619 B.n837 B.n836 10.6151
R1620 B.n836 B.n835 10.6151
R1621 B.n835 B.n66 10.6151
R1622 B.n829 B.n66 10.6151
R1623 B.n829 B.n828 10.6151
R1624 B.n828 B.n827 10.6151
R1625 B.n827 B.n73 10.6151
R1626 B.n821 B.n73 10.6151
R1627 B.n821 B.n820 10.6151
R1628 B.n210 B.n209 9.36635
R1629 B.n232 B.n231 9.36635
R1630 B.n550 B.n444 9.36635
R1631 B.n527 B.n447 9.36635
R1632 B.n907 B.n0 2.81026
R1633 B.n907 B.n1 2.81026
R1634 B.n742 B.t3 1.28667
R1635 B.t1 B.n895 1.28667
R1636 B.n211 B.n210 1.24928
R1637 B.n231 B.n230 1.24928
R1638 B.n547 B.n444 1.24928
R1639 B.n530 B.n447 1.24928
R1640 VP.n13 VP.n12 161.3
R1641 VP.n14 VP.n9 161.3
R1642 VP.n16 VP.n15 161.3
R1643 VP.n17 VP.n8 161.3
R1644 VP.n19 VP.n18 161.3
R1645 VP.n20 VP.n7 161.3
R1646 VP.n42 VP.n0 161.3
R1647 VP.n41 VP.n40 161.3
R1648 VP.n39 VP.n1 161.3
R1649 VP.n38 VP.n37 161.3
R1650 VP.n36 VP.n2 161.3
R1651 VP.n35 VP.n34 161.3
R1652 VP.n33 VP.n32 161.3
R1653 VP.n31 VP.n4 161.3
R1654 VP.n30 VP.n29 161.3
R1655 VP.n28 VP.n5 161.3
R1656 VP.n27 VP.n26 161.3
R1657 VP.n25 VP.n6 161.3
R1658 VP.n11 VP.t2 141.812
R1659 VP.n24 VP.t5 107.995
R1660 VP.n3 VP.t3 107.995
R1661 VP.n43 VP.t1 107.995
R1662 VP.n21 VP.t0 107.995
R1663 VP.n10 VP.t4 107.995
R1664 VP.n24 VP.n23 99.991
R1665 VP.n44 VP.n43 99.991
R1666 VP.n22 VP.n21 99.991
R1667 VP.n11 VP.n10 60.2677
R1668 VP.n30 VP.n5 56.5193
R1669 VP.n37 VP.n1 56.5193
R1670 VP.n15 VP.n8 56.5193
R1671 VP.n23 VP.n22 48.7458
R1672 VP.n26 VP.n25 24.4675
R1673 VP.n26 VP.n5 24.4675
R1674 VP.n31 VP.n30 24.4675
R1675 VP.n32 VP.n31 24.4675
R1676 VP.n36 VP.n35 24.4675
R1677 VP.n37 VP.n36 24.4675
R1678 VP.n41 VP.n1 24.4675
R1679 VP.n42 VP.n41 24.4675
R1680 VP.n19 VP.n8 24.4675
R1681 VP.n20 VP.n19 24.4675
R1682 VP.n14 VP.n13 24.4675
R1683 VP.n15 VP.n14 24.4675
R1684 VP.n32 VP.n3 12.234
R1685 VP.n35 VP.n3 12.234
R1686 VP.n13 VP.n10 12.234
R1687 VP.n25 VP.n24 10.766
R1688 VP.n43 VP.n42 10.766
R1689 VP.n21 VP.n20 10.766
R1690 VP.n12 VP.n11 6.80183
R1691 VP.n22 VP.n7 0.278367
R1692 VP.n23 VP.n6 0.278367
R1693 VP.n44 VP.n0 0.278367
R1694 VP.n12 VP.n9 0.189894
R1695 VP.n16 VP.n9 0.189894
R1696 VP.n17 VP.n16 0.189894
R1697 VP.n18 VP.n17 0.189894
R1698 VP.n18 VP.n7 0.189894
R1699 VP.n27 VP.n6 0.189894
R1700 VP.n28 VP.n27 0.189894
R1701 VP.n29 VP.n28 0.189894
R1702 VP.n29 VP.n4 0.189894
R1703 VP.n33 VP.n4 0.189894
R1704 VP.n34 VP.n33 0.189894
R1705 VP.n34 VP.n2 0.189894
R1706 VP.n38 VP.n2 0.189894
R1707 VP.n39 VP.n38 0.189894
R1708 VP.n40 VP.n39 0.189894
R1709 VP.n40 VP.n0 0.189894
R1710 VP VP.n44 0.153454
R1711 VDD1 VDD1.t3 66.9898
R1712 VDD1.n1 VDD1.t0 66.876
R1713 VDD1.n1 VDD1.n0 63.9221
R1714 VDD1.n3 VDD1.n2 63.3374
R1715 VDD1.n3 VDD1.n1 44.0979
R1716 VDD1.n2 VDD1.t1 1.67421
R1717 VDD1.n2 VDD1.t5 1.67421
R1718 VDD1.n0 VDD1.t2 1.67421
R1719 VDD1.n0 VDD1.t4 1.67421
R1720 VDD1 VDD1.n3 0.582397
C0 VDD2 VN 6.65067f
C1 VDD1 VTAIL 7.67555f
C2 VP VTAIL 6.83827f
C3 VTAIL VN 6.82399f
C4 VP VDD1 6.95842f
C5 VDD1 VN 0.150876f
C6 VDD2 VTAIL 7.72673f
C7 VP VN 6.93172f
C8 VDD2 VDD1 1.42313f
C9 VP VDD2 0.46178f
C10 VDD2 B 5.990422f
C11 VDD1 B 6.316774f
C12 VTAIL B 7.772713f
C13 VN B 12.978339f
C14 VP B 11.612831f
C15 VDD1.t3 B 2.32166f
C16 VDD1.t0 B 2.32081f
C17 VDD1.t2 B 0.20335f
C18 VDD1.t4 B 0.20335f
C19 VDD1.n0 B 1.81521f
C20 VDD1.n1 B 2.64186f
C21 VDD1.t1 B 0.20335f
C22 VDD1.t5 B 0.20335f
C23 VDD1.n2 B 1.81146f
C24 VDD1.n3 B 2.42552f
C25 VP.n0 B 0.03096f
C26 VP.t1 B 1.9974f
C27 VP.n1 B 0.035264f
C28 VP.n2 B 0.023483f
C29 VP.t3 B 1.9974f
C30 VP.n3 B 0.706712f
C31 VP.n4 B 0.023483f
C32 VP.n5 B 0.035264f
C33 VP.n6 B 0.03096f
C34 VP.t5 B 1.9974f
C35 VP.n7 B 0.03096f
C36 VP.t0 B 1.9974f
C37 VP.n8 B 0.035264f
C38 VP.n9 B 0.023483f
C39 VP.t4 B 1.9974f
C40 VP.n10 B 0.775016f
C41 VP.t2 B 2.20118f
C42 VP.n11 B 0.750259f
C43 VP.n12 B 0.227927f
C44 VP.n13 B 0.032962f
C45 VP.n14 B 0.043766f
C46 VP.n15 B 0.033301f
C47 VP.n16 B 0.023483f
C48 VP.n17 B 0.023483f
C49 VP.n18 B 0.023483f
C50 VP.n19 B 0.043766f
C51 VP.n20 B 0.031666f
C52 VP.n21 B 0.787851f
C53 VP.n22 B 1.2587f
C54 VP.n23 B 1.27601f
C55 VP.n24 B 0.787851f
C56 VP.n25 B 0.031666f
C57 VP.n26 B 0.043766f
C58 VP.n27 B 0.023483f
C59 VP.n28 B 0.023483f
C60 VP.n29 B 0.023483f
C61 VP.n30 B 0.033301f
C62 VP.n31 B 0.043766f
C63 VP.n32 B 0.032962f
C64 VP.n33 B 0.023483f
C65 VP.n34 B 0.023483f
C66 VP.n35 B 0.032962f
C67 VP.n36 B 0.043766f
C68 VP.n37 B 0.033301f
C69 VP.n38 B 0.023483f
C70 VP.n39 B 0.023483f
C71 VP.n40 B 0.023483f
C72 VP.n41 B 0.043766f
C73 VP.n42 B 0.031666f
C74 VP.n43 B 0.787851f
C75 VP.n44 B 0.038005f
C76 VDD2.t3 B 2.28594f
C77 VDD2.t2 B 0.200295f
C78 VDD2.t4 B 0.200295f
C79 VDD2.n0 B 1.78793f
C80 VDD2.n1 B 2.49502f
C81 VDD2.t5 B 2.27567f
C82 VDD2.n2 B 2.39159f
C83 VDD2.t0 B 0.200295f
C84 VDD2.t1 B 0.200295f
C85 VDD2.n3 B 1.7879f
C86 VTAIL.t10 B 0.221907f
C87 VTAIL.t11 B 0.221907f
C88 VTAIL.n0 B 1.90865f
C89 VTAIL.n1 B 0.418229f
C90 VTAIL.t3 B 2.43448f
C91 VTAIL.n2 B 0.640023f
C92 VTAIL.t0 B 0.221907f
C93 VTAIL.t5 B 0.221907f
C94 VTAIL.n3 B 1.90865f
C95 VTAIL.n4 B 1.92095f
C96 VTAIL.t7 B 0.221907f
C97 VTAIL.t9 B 0.221907f
C98 VTAIL.n5 B 1.90865f
C99 VTAIL.n6 B 1.92094f
C100 VTAIL.t6 B 2.43449f
C101 VTAIL.n7 B 0.640017f
C102 VTAIL.t1 B 0.221907f
C103 VTAIL.t2 B 0.221907f
C104 VTAIL.n8 B 1.90865f
C105 VTAIL.n9 B 0.560648f
C106 VTAIL.t4 B 2.43448f
C107 VTAIL.n10 B 1.80449f
C108 VTAIL.t8 B 2.43448f
C109 VTAIL.n11 B 1.75108f
C110 VN.n0 B 0.030462f
C111 VN.t1 B 1.96532f
C112 VN.n1 B 0.034698f
C113 VN.n2 B 0.023105f
C114 VN.t3 B 1.96532f
C115 VN.n3 B 0.762568f
C116 VN.t2 B 2.16582f
C117 VN.n4 B 0.738209f
C118 VN.n5 B 0.224266f
C119 VN.n6 B 0.032433f
C120 VN.n7 B 0.043063f
C121 VN.n8 B 0.032766f
C122 VN.n9 B 0.023105f
C123 VN.n10 B 0.023105f
C124 VN.n11 B 0.023105f
C125 VN.n12 B 0.043063f
C126 VN.n13 B 0.031157f
C127 VN.n14 B 0.775197f
C128 VN.n15 B 0.037394f
C129 VN.n16 B 0.030462f
C130 VN.t0 B 1.96532f
C131 VN.n17 B 0.034698f
C132 VN.n18 B 0.023105f
C133 VN.t5 B 1.96532f
C134 VN.n19 B 0.762568f
C135 VN.t4 B 2.16582f
C136 VN.n20 B 0.738209f
C137 VN.n21 B 0.224266f
C138 VN.n22 B 0.032433f
C139 VN.n23 B 0.043063f
C140 VN.n24 B 0.032766f
C141 VN.n25 B 0.023105f
C142 VN.n26 B 0.023105f
C143 VN.n27 B 0.023105f
C144 VN.n28 B 0.043063f
C145 VN.n29 B 0.031157f
C146 VN.n30 B 0.775197f
C147 VN.n31 B 1.25094f
.ends

