* NGSPICE file created from diff_pair_sample_1351.ext - technology: sky130A

.subckt diff_pair_sample_1351 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t10 VP.t0 VDD1.t2 w_n1674_n2146# sky130_fd_pr__pfet_01v8 ad=0.97185 pd=6.22 as=0.97185 ps=6.22 w=5.89 l=0.55
X1 VTAIL.t9 VP.t1 VDD1.t4 w_n1674_n2146# sky130_fd_pr__pfet_01v8 ad=0.97185 pd=6.22 as=0.97185 ps=6.22 w=5.89 l=0.55
X2 VDD1.t0 VP.t2 VTAIL.t8 w_n1674_n2146# sky130_fd_pr__pfet_01v8 ad=2.2971 pd=12.56 as=0.97185 ps=6.22 w=5.89 l=0.55
X3 VDD1.t3 VP.t3 VTAIL.t7 w_n1674_n2146# sky130_fd_pr__pfet_01v8 ad=0.97185 pd=6.22 as=2.2971 ps=12.56 w=5.89 l=0.55
X4 VDD2.t5 VN.t0 VTAIL.t0 w_n1674_n2146# sky130_fd_pr__pfet_01v8 ad=2.2971 pd=12.56 as=0.97185 ps=6.22 w=5.89 l=0.55
X5 VDD1.t1 VP.t4 VTAIL.t6 w_n1674_n2146# sky130_fd_pr__pfet_01v8 ad=0.97185 pd=6.22 as=2.2971 ps=12.56 w=5.89 l=0.55
X6 B.t11 B.t9 B.t10 w_n1674_n2146# sky130_fd_pr__pfet_01v8 ad=2.2971 pd=12.56 as=0 ps=0 w=5.89 l=0.55
X7 VDD2.t4 VN.t1 VTAIL.t4 w_n1674_n2146# sky130_fd_pr__pfet_01v8 ad=0.97185 pd=6.22 as=2.2971 ps=12.56 w=5.89 l=0.55
X8 VDD2.t3 VN.t2 VTAIL.t1 w_n1674_n2146# sky130_fd_pr__pfet_01v8 ad=0.97185 pd=6.22 as=2.2971 ps=12.56 w=5.89 l=0.55
X9 VDD2.t2 VN.t3 VTAIL.t3 w_n1674_n2146# sky130_fd_pr__pfet_01v8 ad=2.2971 pd=12.56 as=0.97185 ps=6.22 w=5.89 l=0.55
X10 VTAIL.t2 VN.t4 VDD2.t1 w_n1674_n2146# sky130_fd_pr__pfet_01v8 ad=0.97185 pd=6.22 as=0.97185 ps=6.22 w=5.89 l=0.55
X11 B.t8 B.t6 B.t7 w_n1674_n2146# sky130_fd_pr__pfet_01v8 ad=2.2971 pd=12.56 as=0 ps=0 w=5.89 l=0.55
X12 VDD1.t5 VP.t5 VTAIL.t5 w_n1674_n2146# sky130_fd_pr__pfet_01v8 ad=2.2971 pd=12.56 as=0.97185 ps=6.22 w=5.89 l=0.55
X13 B.t5 B.t3 B.t4 w_n1674_n2146# sky130_fd_pr__pfet_01v8 ad=2.2971 pd=12.56 as=0 ps=0 w=5.89 l=0.55
X14 B.t2 B.t0 B.t1 w_n1674_n2146# sky130_fd_pr__pfet_01v8 ad=2.2971 pd=12.56 as=0 ps=0 w=5.89 l=0.55
X15 VTAIL.t11 VN.t5 VDD2.t0 w_n1674_n2146# sky130_fd_pr__pfet_01v8 ad=0.97185 pd=6.22 as=0.97185 ps=6.22 w=5.89 l=0.55
R0 VP.n1 VP.t5 356.772
R1 VP.n6 VP.t2 329.952
R2 VP.n7 VP.t1 329.952
R3 VP.n8 VP.t4 329.952
R4 VP.n3 VP.t3 329.952
R5 VP.n2 VP.t0 329.952
R6 VP.n9 VP.n8 161.3
R7 VP.n4 VP.n3 161.3
R8 VP.n6 VP.n5 161.3
R9 VP.n7 VP.n0 80.6037
R10 VP.n7 VP.n6 48.2005
R11 VP.n8 VP.n7 48.2005
R12 VP.n3 VP.n2 48.2005
R13 VP.n4 VP.n1 45.1367
R14 VP.n5 VP.n4 36.0232
R15 VP.n2 VP.n1 13.3799
R16 VP.n5 VP.n0 0.285035
R17 VP.n9 VP.n0 0.285035
R18 VP VP.n9 0.0516364
R19 VDD1.n26 VDD1.n0 756.745
R20 VDD1.n57 VDD1.n31 756.745
R21 VDD1.n27 VDD1.n26 585
R22 VDD1.n25 VDD1.n24 585
R23 VDD1.n4 VDD1.n3 585
R24 VDD1.n19 VDD1.n18 585
R25 VDD1.n17 VDD1.n16 585
R26 VDD1.n8 VDD1.n7 585
R27 VDD1.n11 VDD1.n10 585
R28 VDD1.n42 VDD1.n41 585
R29 VDD1.n39 VDD1.n38 585
R30 VDD1.n48 VDD1.n47 585
R31 VDD1.n50 VDD1.n49 585
R32 VDD1.n35 VDD1.n34 585
R33 VDD1.n56 VDD1.n55 585
R34 VDD1.n58 VDD1.n57 585
R35 VDD1.t5 VDD1.n9 327.601
R36 VDD1.t0 VDD1.n40 327.601
R37 VDD1.n26 VDD1.n25 171.744
R38 VDD1.n25 VDD1.n3 171.744
R39 VDD1.n18 VDD1.n3 171.744
R40 VDD1.n18 VDD1.n17 171.744
R41 VDD1.n17 VDD1.n7 171.744
R42 VDD1.n10 VDD1.n7 171.744
R43 VDD1.n41 VDD1.n38 171.744
R44 VDD1.n48 VDD1.n38 171.744
R45 VDD1.n49 VDD1.n48 171.744
R46 VDD1.n49 VDD1.n34 171.744
R47 VDD1.n56 VDD1.n34 171.744
R48 VDD1.n57 VDD1.n56 171.744
R49 VDD1.n63 VDD1.n62 90.2951
R50 VDD1.n65 VDD1.n64 90.1608
R51 VDD1.n10 VDD1.t5 85.8723
R52 VDD1.n41 VDD1.t0 85.8723
R53 VDD1 VDD1.n30 47.358
R54 VDD1.n63 VDD1.n61 47.2444
R55 VDD1.n65 VDD1.n63 32.2207
R56 VDD1.n11 VDD1.n9 16.3865
R57 VDD1.n42 VDD1.n40 16.3865
R58 VDD1.n12 VDD1.n8 12.8005
R59 VDD1.n43 VDD1.n39 12.8005
R60 VDD1.n16 VDD1.n15 12.0247
R61 VDD1.n47 VDD1.n46 12.0247
R62 VDD1.n19 VDD1.n6 11.249
R63 VDD1.n50 VDD1.n37 11.249
R64 VDD1.n20 VDD1.n4 10.4732
R65 VDD1.n51 VDD1.n35 10.4732
R66 VDD1.n24 VDD1.n23 9.69747
R67 VDD1.n55 VDD1.n54 9.69747
R68 VDD1.n30 VDD1.n29 9.45567
R69 VDD1.n61 VDD1.n60 9.45567
R70 VDD1.n29 VDD1.n28 9.3005
R71 VDD1.n2 VDD1.n1 9.3005
R72 VDD1.n23 VDD1.n22 9.3005
R73 VDD1.n21 VDD1.n20 9.3005
R74 VDD1.n6 VDD1.n5 9.3005
R75 VDD1.n15 VDD1.n14 9.3005
R76 VDD1.n13 VDD1.n12 9.3005
R77 VDD1.n60 VDD1.n59 9.3005
R78 VDD1.n33 VDD1.n32 9.3005
R79 VDD1.n54 VDD1.n53 9.3005
R80 VDD1.n52 VDD1.n51 9.3005
R81 VDD1.n37 VDD1.n36 9.3005
R82 VDD1.n46 VDD1.n45 9.3005
R83 VDD1.n44 VDD1.n43 9.3005
R84 VDD1.n27 VDD1.n2 8.92171
R85 VDD1.n58 VDD1.n33 8.92171
R86 VDD1.n28 VDD1.n0 8.14595
R87 VDD1.n59 VDD1.n31 8.14595
R88 VDD1.n30 VDD1.n0 5.81868
R89 VDD1.n61 VDD1.n31 5.81868
R90 VDD1.n64 VDD1.t2 5.51918
R91 VDD1.n64 VDD1.t3 5.51918
R92 VDD1.n62 VDD1.t4 5.51918
R93 VDD1.n62 VDD1.t1 5.51918
R94 VDD1.n28 VDD1.n27 5.04292
R95 VDD1.n59 VDD1.n58 5.04292
R96 VDD1.n24 VDD1.n2 4.26717
R97 VDD1.n55 VDD1.n33 4.26717
R98 VDD1.n13 VDD1.n9 3.71286
R99 VDD1.n44 VDD1.n40 3.71286
R100 VDD1.n23 VDD1.n4 3.49141
R101 VDD1.n54 VDD1.n35 3.49141
R102 VDD1.n20 VDD1.n19 2.71565
R103 VDD1.n51 VDD1.n50 2.71565
R104 VDD1.n16 VDD1.n6 1.93989
R105 VDD1.n47 VDD1.n37 1.93989
R106 VDD1.n15 VDD1.n8 1.16414
R107 VDD1.n46 VDD1.n39 1.16414
R108 VDD1.n12 VDD1.n11 0.388379
R109 VDD1.n43 VDD1.n42 0.388379
R110 VDD1.n29 VDD1.n1 0.155672
R111 VDD1.n22 VDD1.n1 0.155672
R112 VDD1.n22 VDD1.n21 0.155672
R113 VDD1.n21 VDD1.n5 0.155672
R114 VDD1.n14 VDD1.n5 0.155672
R115 VDD1.n14 VDD1.n13 0.155672
R116 VDD1.n45 VDD1.n44 0.155672
R117 VDD1.n45 VDD1.n36 0.155672
R118 VDD1.n52 VDD1.n36 0.155672
R119 VDD1.n53 VDD1.n52 0.155672
R120 VDD1.n53 VDD1.n32 0.155672
R121 VDD1.n60 VDD1.n32 0.155672
R122 VDD1 VDD1.n65 0.131966
R123 VTAIL.n130 VTAIL.n104 756.745
R124 VTAIL.n28 VTAIL.n2 756.745
R125 VTAIL.n98 VTAIL.n72 756.745
R126 VTAIL.n64 VTAIL.n38 756.745
R127 VTAIL.n115 VTAIL.n114 585
R128 VTAIL.n112 VTAIL.n111 585
R129 VTAIL.n121 VTAIL.n120 585
R130 VTAIL.n123 VTAIL.n122 585
R131 VTAIL.n108 VTAIL.n107 585
R132 VTAIL.n129 VTAIL.n128 585
R133 VTAIL.n131 VTAIL.n130 585
R134 VTAIL.n13 VTAIL.n12 585
R135 VTAIL.n10 VTAIL.n9 585
R136 VTAIL.n19 VTAIL.n18 585
R137 VTAIL.n21 VTAIL.n20 585
R138 VTAIL.n6 VTAIL.n5 585
R139 VTAIL.n27 VTAIL.n26 585
R140 VTAIL.n29 VTAIL.n28 585
R141 VTAIL.n99 VTAIL.n98 585
R142 VTAIL.n97 VTAIL.n96 585
R143 VTAIL.n76 VTAIL.n75 585
R144 VTAIL.n91 VTAIL.n90 585
R145 VTAIL.n89 VTAIL.n88 585
R146 VTAIL.n80 VTAIL.n79 585
R147 VTAIL.n83 VTAIL.n82 585
R148 VTAIL.n65 VTAIL.n64 585
R149 VTAIL.n63 VTAIL.n62 585
R150 VTAIL.n42 VTAIL.n41 585
R151 VTAIL.n57 VTAIL.n56 585
R152 VTAIL.n55 VTAIL.n54 585
R153 VTAIL.n46 VTAIL.n45 585
R154 VTAIL.n49 VTAIL.n48 585
R155 VTAIL.t1 VTAIL.n113 327.601
R156 VTAIL.t6 VTAIL.n11 327.601
R157 VTAIL.t7 VTAIL.n81 327.601
R158 VTAIL.t4 VTAIL.n47 327.601
R159 VTAIL.n114 VTAIL.n111 171.744
R160 VTAIL.n121 VTAIL.n111 171.744
R161 VTAIL.n122 VTAIL.n121 171.744
R162 VTAIL.n122 VTAIL.n107 171.744
R163 VTAIL.n129 VTAIL.n107 171.744
R164 VTAIL.n130 VTAIL.n129 171.744
R165 VTAIL.n12 VTAIL.n9 171.744
R166 VTAIL.n19 VTAIL.n9 171.744
R167 VTAIL.n20 VTAIL.n19 171.744
R168 VTAIL.n20 VTAIL.n5 171.744
R169 VTAIL.n27 VTAIL.n5 171.744
R170 VTAIL.n28 VTAIL.n27 171.744
R171 VTAIL.n98 VTAIL.n97 171.744
R172 VTAIL.n97 VTAIL.n75 171.744
R173 VTAIL.n90 VTAIL.n75 171.744
R174 VTAIL.n90 VTAIL.n89 171.744
R175 VTAIL.n89 VTAIL.n79 171.744
R176 VTAIL.n82 VTAIL.n79 171.744
R177 VTAIL.n64 VTAIL.n63 171.744
R178 VTAIL.n63 VTAIL.n41 171.744
R179 VTAIL.n56 VTAIL.n41 171.744
R180 VTAIL.n56 VTAIL.n55 171.744
R181 VTAIL.n55 VTAIL.n45 171.744
R182 VTAIL.n48 VTAIL.n45 171.744
R183 VTAIL.n114 VTAIL.t1 85.8723
R184 VTAIL.n12 VTAIL.t6 85.8723
R185 VTAIL.n82 VTAIL.t7 85.8723
R186 VTAIL.n48 VTAIL.t4 85.8723
R187 VTAIL.n71 VTAIL.n70 73.4821
R188 VTAIL.n37 VTAIL.n36 73.4821
R189 VTAIL.n1 VTAIL.n0 73.482
R190 VTAIL.n35 VTAIL.n34 73.482
R191 VTAIL.n135 VTAIL.n134 30.052
R192 VTAIL.n33 VTAIL.n32 30.052
R193 VTAIL.n103 VTAIL.n102 30.052
R194 VTAIL.n69 VTAIL.n68 30.052
R195 VTAIL.n37 VTAIL.n35 18.9617
R196 VTAIL.n135 VTAIL.n103 18.2031
R197 VTAIL.n115 VTAIL.n113 16.3865
R198 VTAIL.n13 VTAIL.n11 16.3865
R199 VTAIL.n83 VTAIL.n81 16.3865
R200 VTAIL.n49 VTAIL.n47 16.3865
R201 VTAIL.n116 VTAIL.n112 12.8005
R202 VTAIL.n14 VTAIL.n10 12.8005
R203 VTAIL.n84 VTAIL.n80 12.8005
R204 VTAIL.n50 VTAIL.n46 12.8005
R205 VTAIL.n120 VTAIL.n119 12.0247
R206 VTAIL.n18 VTAIL.n17 12.0247
R207 VTAIL.n88 VTAIL.n87 12.0247
R208 VTAIL.n54 VTAIL.n53 12.0247
R209 VTAIL.n123 VTAIL.n110 11.249
R210 VTAIL.n21 VTAIL.n8 11.249
R211 VTAIL.n91 VTAIL.n78 11.249
R212 VTAIL.n57 VTAIL.n44 11.249
R213 VTAIL.n124 VTAIL.n108 10.4732
R214 VTAIL.n22 VTAIL.n6 10.4732
R215 VTAIL.n92 VTAIL.n76 10.4732
R216 VTAIL.n58 VTAIL.n42 10.4732
R217 VTAIL.n128 VTAIL.n127 9.69747
R218 VTAIL.n26 VTAIL.n25 9.69747
R219 VTAIL.n96 VTAIL.n95 9.69747
R220 VTAIL.n62 VTAIL.n61 9.69747
R221 VTAIL.n134 VTAIL.n133 9.45567
R222 VTAIL.n32 VTAIL.n31 9.45567
R223 VTAIL.n102 VTAIL.n101 9.45567
R224 VTAIL.n68 VTAIL.n67 9.45567
R225 VTAIL.n133 VTAIL.n132 9.3005
R226 VTAIL.n106 VTAIL.n105 9.3005
R227 VTAIL.n127 VTAIL.n126 9.3005
R228 VTAIL.n125 VTAIL.n124 9.3005
R229 VTAIL.n110 VTAIL.n109 9.3005
R230 VTAIL.n119 VTAIL.n118 9.3005
R231 VTAIL.n117 VTAIL.n116 9.3005
R232 VTAIL.n31 VTAIL.n30 9.3005
R233 VTAIL.n4 VTAIL.n3 9.3005
R234 VTAIL.n25 VTAIL.n24 9.3005
R235 VTAIL.n23 VTAIL.n22 9.3005
R236 VTAIL.n8 VTAIL.n7 9.3005
R237 VTAIL.n17 VTAIL.n16 9.3005
R238 VTAIL.n15 VTAIL.n14 9.3005
R239 VTAIL.n101 VTAIL.n100 9.3005
R240 VTAIL.n74 VTAIL.n73 9.3005
R241 VTAIL.n95 VTAIL.n94 9.3005
R242 VTAIL.n93 VTAIL.n92 9.3005
R243 VTAIL.n78 VTAIL.n77 9.3005
R244 VTAIL.n87 VTAIL.n86 9.3005
R245 VTAIL.n85 VTAIL.n84 9.3005
R246 VTAIL.n67 VTAIL.n66 9.3005
R247 VTAIL.n40 VTAIL.n39 9.3005
R248 VTAIL.n61 VTAIL.n60 9.3005
R249 VTAIL.n59 VTAIL.n58 9.3005
R250 VTAIL.n44 VTAIL.n43 9.3005
R251 VTAIL.n53 VTAIL.n52 9.3005
R252 VTAIL.n51 VTAIL.n50 9.3005
R253 VTAIL.n131 VTAIL.n106 8.92171
R254 VTAIL.n29 VTAIL.n4 8.92171
R255 VTAIL.n99 VTAIL.n74 8.92171
R256 VTAIL.n65 VTAIL.n40 8.92171
R257 VTAIL.n132 VTAIL.n104 8.14595
R258 VTAIL.n30 VTAIL.n2 8.14595
R259 VTAIL.n100 VTAIL.n72 8.14595
R260 VTAIL.n66 VTAIL.n38 8.14595
R261 VTAIL.n134 VTAIL.n104 5.81868
R262 VTAIL.n32 VTAIL.n2 5.81868
R263 VTAIL.n102 VTAIL.n72 5.81868
R264 VTAIL.n68 VTAIL.n38 5.81868
R265 VTAIL.n0 VTAIL.t0 5.51918
R266 VTAIL.n0 VTAIL.t11 5.51918
R267 VTAIL.n34 VTAIL.t8 5.51918
R268 VTAIL.n34 VTAIL.t9 5.51918
R269 VTAIL.n70 VTAIL.t5 5.51918
R270 VTAIL.n70 VTAIL.t10 5.51918
R271 VTAIL.n36 VTAIL.t3 5.51918
R272 VTAIL.n36 VTAIL.t2 5.51918
R273 VTAIL.n132 VTAIL.n131 5.04292
R274 VTAIL.n30 VTAIL.n29 5.04292
R275 VTAIL.n100 VTAIL.n99 5.04292
R276 VTAIL.n66 VTAIL.n65 5.04292
R277 VTAIL.n128 VTAIL.n106 4.26717
R278 VTAIL.n26 VTAIL.n4 4.26717
R279 VTAIL.n96 VTAIL.n74 4.26717
R280 VTAIL.n62 VTAIL.n40 4.26717
R281 VTAIL.n85 VTAIL.n81 3.71286
R282 VTAIL.n51 VTAIL.n47 3.71286
R283 VTAIL.n117 VTAIL.n113 3.71286
R284 VTAIL.n15 VTAIL.n11 3.71286
R285 VTAIL.n127 VTAIL.n108 3.49141
R286 VTAIL.n25 VTAIL.n6 3.49141
R287 VTAIL.n95 VTAIL.n76 3.49141
R288 VTAIL.n61 VTAIL.n42 3.49141
R289 VTAIL.n124 VTAIL.n123 2.71565
R290 VTAIL.n22 VTAIL.n21 2.71565
R291 VTAIL.n92 VTAIL.n91 2.71565
R292 VTAIL.n58 VTAIL.n57 2.71565
R293 VTAIL.n120 VTAIL.n110 1.93989
R294 VTAIL.n18 VTAIL.n8 1.93989
R295 VTAIL.n88 VTAIL.n78 1.93989
R296 VTAIL.n54 VTAIL.n44 1.93989
R297 VTAIL.n119 VTAIL.n112 1.16414
R298 VTAIL.n17 VTAIL.n10 1.16414
R299 VTAIL.n87 VTAIL.n80 1.16414
R300 VTAIL.n53 VTAIL.n46 1.16414
R301 VTAIL.n71 VTAIL.n69 0.849638
R302 VTAIL.n33 VTAIL.n1 0.849638
R303 VTAIL.n69 VTAIL.n37 0.759121
R304 VTAIL.n103 VTAIL.n71 0.759121
R305 VTAIL.n35 VTAIL.n33 0.759121
R306 VTAIL VTAIL.n135 0.511276
R307 VTAIL.n116 VTAIL.n115 0.388379
R308 VTAIL.n14 VTAIL.n13 0.388379
R309 VTAIL.n84 VTAIL.n83 0.388379
R310 VTAIL.n50 VTAIL.n49 0.388379
R311 VTAIL VTAIL.n1 0.248345
R312 VTAIL.n118 VTAIL.n117 0.155672
R313 VTAIL.n118 VTAIL.n109 0.155672
R314 VTAIL.n125 VTAIL.n109 0.155672
R315 VTAIL.n126 VTAIL.n125 0.155672
R316 VTAIL.n126 VTAIL.n105 0.155672
R317 VTAIL.n133 VTAIL.n105 0.155672
R318 VTAIL.n16 VTAIL.n15 0.155672
R319 VTAIL.n16 VTAIL.n7 0.155672
R320 VTAIL.n23 VTAIL.n7 0.155672
R321 VTAIL.n24 VTAIL.n23 0.155672
R322 VTAIL.n24 VTAIL.n3 0.155672
R323 VTAIL.n31 VTAIL.n3 0.155672
R324 VTAIL.n101 VTAIL.n73 0.155672
R325 VTAIL.n94 VTAIL.n73 0.155672
R326 VTAIL.n94 VTAIL.n93 0.155672
R327 VTAIL.n93 VTAIL.n77 0.155672
R328 VTAIL.n86 VTAIL.n77 0.155672
R329 VTAIL.n86 VTAIL.n85 0.155672
R330 VTAIL.n67 VTAIL.n39 0.155672
R331 VTAIL.n60 VTAIL.n39 0.155672
R332 VTAIL.n60 VTAIL.n59 0.155672
R333 VTAIL.n59 VTAIL.n43 0.155672
R334 VTAIL.n52 VTAIL.n43 0.155672
R335 VTAIL.n52 VTAIL.n51 0.155672
R336 VN.n0 VN.t0 356.772
R337 VN.n4 VN.t1 356.772
R338 VN.n1 VN.t5 329.952
R339 VN.n2 VN.t2 329.952
R340 VN.n5 VN.t4 329.952
R341 VN.n6 VN.t3 329.952
R342 VN.n3 VN.n2 161.3
R343 VN.n7 VN.n6 161.3
R344 VN.n2 VN.n1 48.2005
R345 VN.n6 VN.n5 48.2005
R346 VN.n7 VN.n4 45.1367
R347 VN.n3 VN.n0 45.1367
R348 VN VN.n7 36.4039
R349 VN.n5 VN.n4 13.3799
R350 VN.n1 VN.n0 13.3799
R351 VN VN.n3 0.0516364
R352 VDD2.n59 VDD2.n33 756.745
R353 VDD2.n26 VDD2.n0 756.745
R354 VDD2.n60 VDD2.n59 585
R355 VDD2.n58 VDD2.n57 585
R356 VDD2.n37 VDD2.n36 585
R357 VDD2.n52 VDD2.n51 585
R358 VDD2.n50 VDD2.n49 585
R359 VDD2.n41 VDD2.n40 585
R360 VDD2.n44 VDD2.n43 585
R361 VDD2.n11 VDD2.n10 585
R362 VDD2.n8 VDD2.n7 585
R363 VDD2.n17 VDD2.n16 585
R364 VDD2.n19 VDD2.n18 585
R365 VDD2.n4 VDD2.n3 585
R366 VDD2.n25 VDD2.n24 585
R367 VDD2.n27 VDD2.n26 585
R368 VDD2.t2 VDD2.n42 327.601
R369 VDD2.t5 VDD2.n9 327.601
R370 VDD2.n59 VDD2.n58 171.744
R371 VDD2.n58 VDD2.n36 171.744
R372 VDD2.n51 VDD2.n36 171.744
R373 VDD2.n51 VDD2.n50 171.744
R374 VDD2.n50 VDD2.n40 171.744
R375 VDD2.n43 VDD2.n40 171.744
R376 VDD2.n10 VDD2.n7 171.744
R377 VDD2.n17 VDD2.n7 171.744
R378 VDD2.n18 VDD2.n17 171.744
R379 VDD2.n18 VDD2.n3 171.744
R380 VDD2.n25 VDD2.n3 171.744
R381 VDD2.n26 VDD2.n25 171.744
R382 VDD2.n32 VDD2.n31 90.2951
R383 VDD2 VDD2.n65 90.2922
R384 VDD2.n43 VDD2.t2 85.8723
R385 VDD2.n10 VDD2.t5 85.8723
R386 VDD2.n32 VDD2.n30 47.2444
R387 VDD2.n64 VDD2.n63 46.7308
R388 VDD2.n64 VDD2.n32 31.2584
R389 VDD2.n44 VDD2.n42 16.3865
R390 VDD2.n11 VDD2.n9 16.3865
R391 VDD2.n45 VDD2.n41 12.8005
R392 VDD2.n12 VDD2.n8 12.8005
R393 VDD2.n49 VDD2.n48 12.0247
R394 VDD2.n16 VDD2.n15 12.0247
R395 VDD2.n52 VDD2.n39 11.249
R396 VDD2.n19 VDD2.n6 11.249
R397 VDD2.n53 VDD2.n37 10.4732
R398 VDD2.n20 VDD2.n4 10.4732
R399 VDD2.n57 VDD2.n56 9.69747
R400 VDD2.n24 VDD2.n23 9.69747
R401 VDD2.n63 VDD2.n62 9.45567
R402 VDD2.n30 VDD2.n29 9.45567
R403 VDD2.n62 VDD2.n61 9.3005
R404 VDD2.n35 VDD2.n34 9.3005
R405 VDD2.n56 VDD2.n55 9.3005
R406 VDD2.n54 VDD2.n53 9.3005
R407 VDD2.n39 VDD2.n38 9.3005
R408 VDD2.n48 VDD2.n47 9.3005
R409 VDD2.n46 VDD2.n45 9.3005
R410 VDD2.n29 VDD2.n28 9.3005
R411 VDD2.n2 VDD2.n1 9.3005
R412 VDD2.n23 VDD2.n22 9.3005
R413 VDD2.n21 VDD2.n20 9.3005
R414 VDD2.n6 VDD2.n5 9.3005
R415 VDD2.n15 VDD2.n14 9.3005
R416 VDD2.n13 VDD2.n12 9.3005
R417 VDD2.n60 VDD2.n35 8.92171
R418 VDD2.n27 VDD2.n2 8.92171
R419 VDD2.n61 VDD2.n33 8.14595
R420 VDD2.n28 VDD2.n0 8.14595
R421 VDD2.n63 VDD2.n33 5.81868
R422 VDD2.n30 VDD2.n0 5.81868
R423 VDD2.n65 VDD2.t1 5.51918
R424 VDD2.n65 VDD2.t4 5.51918
R425 VDD2.n31 VDD2.t0 5.51918
R426 VDD2.n31 VDD2.t3 5.51918
R427 VDD2.n61 VDD2.n60 5.04292
R428 VDD2.n28 VDD2.n27 5.04292
R429 VDD2.n57 VDD2.n35 4.26717
R430 VDD2.n24 VDD2.n2 4.26717
R431 VDD2.n46 VDD2.n42 3.71286
R432 VDD2.n13 VDD2.n9 3.71286
R433 VDD2.n56 VDD2.n37 3.49141
R434 VDD2.n23 VDD2.n4 3.49141
R435 VDD2.n53 VDD2.n52 2.71565
R436 VDD2.n20 VDD2.n19 2.71565
R437 VDD2.n49 VDD2.n39 1.93989
R438 VDD2.n16 VDD2.n6 1.93989
R439 VDD2.n48 VDD2.n41 1.16414
R440 VDD2.n15 VDD2.n8 1.16414
R441 VDD2 VDD2.n64 0.627655
R442 VDD2.n45 VDD2.n44 0.388379
R443 VDD2.n12 VDD2.n11 0.388379
R444 VDD2.n62 VDD2.n34 0.155672
R445 VDD2.n55 VDD2.n34 0.155672
R446 VDD2.n55 VDD2.n54 0.155672
R447 VDD2.n54 VDD2.n38 0.155672
R448 VDD2.n47 VDD2.n38 0.155672
R449 VDD2.n47 VDD2.n46 0.155672
R450 VDD2.n14 VDD2.n13 0.155672
R451 VDD2.n14 VDD2.n5 0.155672
R452 VDD2.n21 VDD2.n5 0.155672
R453 VDD2.n22 VDD2.n21 0.155672
R454 VDD2.n22 VDD2.n1 0.155672
R455 VDD2.n29 VDD2.n1 0.155672
R456 B.n216 B.n215 585
R457 B.n214 B.n63 585
R458 B.n213 B.n212 585
R459 B.n211 B.n64 585
R460 B.n210 B.n209 585
R461 B.n208 B.n65 585
R462 B.n207 B.n206 585
R463 B.n205 B.n66 585
R464 B.n204 B.n203 585
R465 B.n202 B.n67 585
R466 B.n201 B.n200 585
R467 B.n199 B.n68 585
R468 B.n198 B.n197 585
R469 B.n196 B.n69 585
R470 B.n195 B.n194 585
R471 B.n193 B.n70 585
R472 B.n192 B.n191 585
R473 B.n190 B.n71 585
R474 B.n189 B.n188 585
R475 B.n187 B.n72 585
R476 B.n186 B.n185 585
R477 B.n184 B.n73 585
R478 B.n183 B.n182 585
R479 B.n181 B.n74 585
R480 B.n180 B.n179 585
R481 B.n175 B.n75 585
R482 B.n174 B.n173 585
R483 B.n172 B.n76 585
R484 B.n171 B.n170 585
R485 B.n169 B.n77 585
R486 B.n168 B.n167 585
R487 B.n166 B.n78 585
R488 B.n165 B.n164 585
R489 B.n162 B.n79 585
R490 B.n161 B.n160 585
R491 B.n159 B.n82 585
R492 B.n158 B.n157 585
R493 B.n156 B.n83 585
R494 B.n155 B.n154 585
R495 B.n153 B.n84 585
R496 B.n152 B.n151 585
R497 B.n150 B.n85 585
R498 B.n149 B.n148 585
R499 B.n147 B.n86 585
R500 B.n146 B.n145 585
R501 B.n144 B.n87 585
R502 B.n143 B.n142 585
R503 B.n141 B.n88 585
R504 B.n140 B.n139 585
R505 B.n138 B.n89 585
R506 B.n137 B.n136 585
R507 B.n135 B.n90 585
R508 B.n134 B.n133 585
R509 B.n132 B.n91 585
R510 B.n131 B.n130 585
R511 B.n129 B.n92 585
R512 B.n128 B.n127 585
R513 B.n217 B.n62 585
R514 B.n219 B.n218 585
R515 B.n220 B.n61 585
R516 B.n222 B.n221 585
R517 B.n223 B.n60 585
R518 B.n225 B.n224 585
R519 B.n226 B.n59 585
R520 B.n228 B.n227 585
R521 B.n229 B.n58 585
R522 B.n231 B.n230 585
R523 B.n232 B.n57 585
R524 B.n234 B.n233 585
R525 B.n235 B.n56 585
R526 B.n237 B.n236 585
R527 B.n238 B.n55 585
R528 B.n240 B.n239 585
R529 B.n241 B.n54 585
R530 B.n243 B.n242 585
R531 B.n244 B.n53 585
R532 B.n246 B.n245 585
R533 B.n247 B.n52 585
R534 B.n249 B.n248 585
R535 B.n250 B.n51 585
R536 B.n252 B.n251 585
R537 B.n253 B.n50 585
R538 B.n255 B.n254 585
R539 B.n256 B.n49 585
R540 B.n258 B.n257 585
R541 B.n259 B.n48 585
R542 B.n261 B.n260 585
R543 B.n262 B.n47 585
R544 B.n264 B.n263 585
R545 B.n265 B.n46 585
R546 B.n267 B.n266 585
R547 B.n268 B.n45 585
R548 B.n270 B.n269 585
R549 B.n271 B.n44 585
R550 B.n273 B.n272 585
R551 B.n360 B.n11 585
R552 B.n359 B.n358 585
R553 B.n357 B.n12 585
R554 B.n356 B.n355 585
R555 B.n354 B.n13 585
R556 B.n353 B.n352 585
R557 B.n351 B.n14 585
R558 B.n350 B.n349 585
R559 B.n348 B.n15 585
R560 B.n347 B.n346 585
R561 B.n345 B.n16 585
R562 B.n344 B.n343 585
R563 B.n342 B.n17 585
R564 B.n341 B.n340 585
R565 B.n339 B.n18 585
R566 B.n338 B.n337 585
R567 B.n336 B.n19 585
R568 B.n335 B.n334 585
R569 B.n333 B.n20 585
R570 B.n332 B.n331 585
R571 B.n330 B.n21 585
R572 B.n329 B.n328 585
R573 B.n327 B.n22 585
R574 B.n326 B.n325 585
R575 B.n323 B.n23 585
R576 B.n322 B.n321 585
R577 B.n320 B.n26 585
R578 B.n319 B.n318 585
R579 B.n317 B.n27 585
R580 B.n316 B.n315 585
R581 B.n314 B.n28 585
R582 B.n313 B.n312 585
R583 B.n311 B.n29 585
R584 B.n309 B.n308 585
R585 B.n307 B.n32 585
R586 B.n306 B.n305 585
R587 B.n304 B.n33 585
R588 B.n303 B.n302 585
R589 B.n301 B.n34 585
R590 B.n300 B.n299 585
R591 B.n298 B.n35 585
R592 B.n297 B.n296 585
R593 B.n295 B.n36 585
R594 B.n294 B.n293 585
R595 B.n292 B.n37 585
R596 B.n291 B.n290 585
R597 B.n289 B.n38 585
R598 B.n288 B.n287 585
R599 B.n286 B.n39 585
R600 B.n285 B.n284 585
R601 B.n283 B.n40 585
R602 B.n282 B.n281 585
R603 B.n280 B.n41 585
R604 B.n279 B.n278 585
R605 B.n277 B.n42 585
R606 B.n276 B.n275 585
R607 B.n274 B.n43 585
R608 B.n362 B.n361 585
R609 B.n363 B.n10 585
R610 B.n365 B.n364 585
R611 B.n366 B.n9 585
R612 B.n368 B.n367 585
R613 B.n369 B.n8 585
R614 B.n371 B.n370 585
R615 B.n372 B.n7 585
R616 B.n374 B.n373 585
R617 B.n375 B.n6 585
R618 B.n377 B.n376 585
R619 B.n378 B.n5 585
R620 B.n380 B.n379 585
R621 B.n381 B.n4 585
R622 B.n383 B.n382 585
R623 B.n384 B.n3 585
R624 B.n386 B.n385 585
R625 B.n387 B.n0 585
R626 B.n2 B.n1 585
R627 B.n102 B.n101 585
R628 B.n104 B.n103 585
R629 B.n105 B.n100 585
R630 B.n107 B.n106 585
R631 B.n108 B.n99 585
R632 B.n110 B.n109 585
R633 B.n111 B.n98 585
R634 B.n113 B.n112 585
R635 B.n114 B.n97 585
R636 B.n116 B.n115 585
R637 B.n117 B.n96 585
R638 B.n119 B.n118 585
R639 B.n120 B.n95 585
R640 B.n122 B.n121 585
R641 B.n123 B.n94 585
R642 B.n125 B.n124 585
R643 B.n126 B.n93 585
R644 B.n128 B.n93 482.89
R645 B.n217 B.n216 482.89
R646 B.n272 B.n43 482.89
R647 B.n362 B.n11 482.89
R648 B.n80 B.t6 463.401
R649 B.n176 B.t3 463.401
R650 B.n30 B.t0 463.401
R651 B.n24 B.t9 463.401
R652 B.n176 B.t4 283.127
R653 B.n30 B.t2 283.127
R654 B.n80 B.t7 283.127
R655 B.n24 B.t11 283.127
R656 B.n177 B.t5 266.06
R657 B.n31 B.t1 266.06
R658 B.n81 B.t8 266.06
R659 B.n25 B.t10 266.06
R660 B.n389 B.n388 256.663
R661 B.n388 B.n387 235.042
R662 B.n388 B.n2 235.042
R663 B.n129 B.n128 163.367
R664 B.n130 B.n129 163.367
R665 B.n130 B.n91 163.367
R666 B.n134 B.n91 163.367
R667 B.n135 B.n134 163.367
R668 B.n136 B.n135 163.367
R669 B.n136 B.n89 163.367
R670 B.n140 B.n89 163.367
R671 B.n141 B.n140 163.367
R672 B.n142 B.n141 163.367
R673 B.n142 B.n87 163.367
R674 B.n146 B.n87 163.367
R675 B.n147 B.n146 163.367
R676 B.n148 B.n147 163.367
R677 B.n148 B.n85 163.367
R678 B.n152 B.n85 163.367
R679 B.n153 B.n152 163.367
R680 B.n154 B.n153 163.367
R681 B.n154 B.n83 163.367
R682 B.n158 B.n83 163.367
R683 B.n159 B.n158 163.367
R684 B.n160 B.n159 163.367
R685 B.n160 B.n79 163.367
R686 B.n165 B.n79 163.367
R687 B.n166 B.n165 163.367
R688 B.n167 B.n166 163.367
R689 B.n167 B.n77 163.367
R690 B.n171 B.n77 163.367
R691 B.n172 B.n171 163.367
R692 B.n173 B.n172 163.367
R693 B.n173 B.n75 163.367
R694 B.n180 B.n75 163.367
R695 B.n181 B.n180 163.367
R696 B.n182 B.n181 163.367
R697 B.n182 B.n73 163.367
R698 B.n186 B.n73 163.367
R699 B.n187 B.n186 163.367
R700 B.n188 B.n187 163.367
R701 B.n188 B.n71 163.367
R702 B.n192 B.n71 163.367
R703 B.n193 B.n192 163.367
R704 B.n194 B.n193 163.367
R705 B.n194 B.n69 163.367
R706 B.n198 B.n69 163.367
R707 B.n199 B.n198 163.367
R708 B.n200 B.n199 163.367
R709 B.n200 B.n67 163.367
R710 B.n204 B.n67 163.367
R711 B.n205 B.n204 163.367
R712 B.n206 B.n205 163.367
R713 B.n206 B.n65 163.367
R714 B.n210 B.n65 163.367
R715 B.n211 B.n210 163.367
R716 B.n212 B.n211 163.367
R717 B.n212 B.n63 163.367
R718 B.n216 B.n63 163.367
R719 B.n272 B.n271 163.367
R720 B.n271 B.n270 163.367
R721 B.n270 B.n45 163.367
R722 B.n266 B.n45 163.367
R723 B.n266 B.n265 163.367
R724 B.n265 B.n264 163.367
R725 B.n264 B.n47 163.367
R726 B.n260 B.n47 163.367
R727 B.n260 B.n259 163.367
R728 B.n259 B.n258 163.367
R729 B.n258 B.n49 163.367
R730 B.n254 B.n49 163.367
R731 B.n254 B.n253 163.367
R732 B.n253 B.n252 163.367
R733 B.n252 B.n51 163.367
R734 B.n248 B.n51 163.367
R735 B.n248 B.n247 163.367
R736 B.n247 B.n246 163.367
R737 B.n246 B.n53 163.367
R738 B.n242 B.n53 163.367
R739 B.n242 B.n241 163.367
R740 B.n241 B.n240 163.367
R741 B.n240 B.n55 163.367
R742 B.n236 B.n55 163.367
R743 B.n236 B.n235 163.367
R744 B.n235 B.n234 163.367
R745 B.n234 B.n57 163.367
R746 B.n230 B.n57 163.367
R747 B.n230 B.n229 163.367
R748 B.n229 B.n228 163.367
R749 B.n228 B.n59 163.367
R750 B.n224 B.n59 163.367
R751 B.n224 B.n223 163.367
R752 B.n223 B.n222 163.367
R753 B.n222 B.n61 163.367
R754 B.n218 B.n61 163.367
R755 B.n218 B.n217 163.367
R756 B.n358 B.n11 163.367
R757 B.n358 B.n357 163.367
R758 B.n357 B.n356 163.367
R759 B.n356 B.n13 163.367
R760 B.n352 B.n13 163.367
R761 B.n352 B.n351 163.367
R762 B.n351 B.n350 163.367
R763 B.n350 B.n15 163.367
R764 B.n346 B.n15 163.367
R765 B.n346 B.n345 163.367
R766 B.n345 B.n344 163.367
R767 B.n344 B.n17 163.367
R768 B.n340 B.n17 163.367
R769 B.n340 B.n339 163.367
R770 B.n339 B.n338 163.367
R771 B.n338 B.n19 163.367
R772 B.n334 B.n19 163.367
R773 B.n334 B.n333 163.367
R774 B.n333 B.n332 163.367
R775 B.n332 B.n21 163.367
R776 B.n328 B.n21 163.367
R777 B.n328 B.n327 163.367
R778 B.n327 B.n326 163.367
R779 B.n326 B.n23 163.367
R780 B.n321 B.n23 163.367
R781 B.n321 B.n320 163.367
R782 B.n320 B.n319 163.367
R783 B.n319 B.n27 163.367
R784 B.n315 B.n27 163.367
R785 B.n315 B.n314 163.367
R786 B.n314 B.n313 163.367
R787 B.n313 B.n29 163.367
R788 B.n308 B.n29 163.367
R789 B.n308 B.n307 163.367
R790 B.n307 B.n306 163.367
R791 B.n306 B.n33 163.367
R792 B.n302 B.n33 163.367
R793 B.n302 B.n301 163.367
R794 B.n301 B.n300 163.367
R795 B.n300 B.n35 163.367
R796 B.n296 B.n35 163.367
R797 B.n296 B.n295 163.367
R798 B.n295 B.n294 163.367
R799 B.n294 B.n37 163.367
R800 B.n290 B.n37 163.367
R801 B.n290 B.n289 163.367
R802 B.n289 B.n288 163.367
R803 B.n288 B.n39 163.367
R804 B.n284 B.n39 163.367
R805 B.n284 B.n283 163.367
R806 B.n283 B.n282 163.367
R807 B.n282 B.n41 163.367
R808 B.n278 B.n41 163.367
R809 B.n278 B.n277 163.367
R810 B.n277 B.n276 163.367
R811 B.n276 B.n43 163.367
R812 B.n363 B.n362 163.367
R813 B.n364 B.n363 163.367
R814 B.n364 B.n9 163.367
R815 B.n368 B.n9 163.367
R816 B.n369 B.n368 163.367
R817 B.n370 B.n369 163.367
R818 B.n370 B.n7 163.367
R819 B.n374 B.n7 163.367
R820 B.n375 B.n374 163.367
R821 B.n376 B.n375 163.367
R822 B.n376 B.n5 163.367
R823 B.n380 B.n5 163.367
R824 B.n381 B.n380 163.367
R825 B.n382 B.n381 163.367
R826 B.n382 B.n3 163.367
R827 B.n386 B.n3 163.367
R828 B.n387 B.n386 163.367
R829 B.n101 B.n2 163.367
R830 B.n104 B.n101 163.367
R831 B.n105 B.n104 163.367
R832 B.n106 B.n105 163.367
R833 B.n106 B.n99 163.367
R834 B.n110 B.n99 163.367
R835 B.n111 B.n110 163.367
R836 B.n112 B.n111 163.367
R837 B.n112 B.n97 163.367
R838 B.n116 B.n97 163.367
R839 B.n117 B.n116 163.367
R840 B.n118 B.n117 163.367
R841 B.n118 B.n95 163.367
R842 B.n122 B.n95 163.367
R843 B.n123 B.n122 163.367
R844 B.n124 B.n123 163.367
R845 B.n124 B.n93 163.367
R846 B.n163 B.n81 59.5399
R847 B.n178 B.n177 59.5399
R848 B.n310 B.n31 59.5399
R849 B.n324 B.n25 59.5399
R850 B.n361 B.n360 31.3761
R851 B.n274 B.n273 31.3761
R852 B.n215 B.n62 31.3761
R853 B.n127 B.n126 31.3761
R854 B B.n389 18.0485
R855 B.n81 B.n80 17.0672
R856 B.n177 B.n176 17.0672
R857 B.n31 B.n30 17.0672
R858 B.n25 B.n24 17.0672
R859 B.n361 B.n10 10.6151
R860 B.n365 B.n10 10.6151
R861 B.n366 B.n365 10.6151
R862 B.n367 B.n366 10.6151
R863 B.n367 B.n8 10.6151
R864 B.n371 B.n8 10.6151
R865 B.n372 B.n371 10.6151
R866 B.n373 B.n372 10.6151
R867 B.n373 B.n6 10.6151
R868 B.n377 B.n6 10.6151
R869 B.n378 B.n377 10.6151
R870 B.n379 B.n378 10.6151
R871 B.n379 B.n4 10.6151
R872 B.n383 B.n4 10.6151
R873 B.n384 B.n383 10.6151
R874 B.n385 B.n384 10.6151
R875 B.n385 B.n0 10.6151
R876 B.n360 B.n359 10.6151
R877 B.n359 B.n12 10.6151
R878 B.n355 B.n12 10.6151
R879 B.n355 B.n354 10.6151
R880 B.n354 B.n353 10.6151
R881 B.n353 B.n14 10.6151
R882 B.n349 B.n14 10.6151
R883 B.n349 B.n348 10.6151
R884 B.n348 B.n347 10.6151
R885 B.n347 B.n16 10.6151
R886 B.n343 B.n16 10.6151
R887 B.n343 B.n342 10.6151
R888 B.n342 B.n341 10.6151
R889 B.n341 B.n18 10.6151
R890 B.n337 B.n18 10.6151
R891 B.n337 B.n336 10.6151
R892 B.n336 B.n335 10.6151
R893 B.n335 B.n20 10.6151
R894 B.n331 B.n20 10.6151
R895 B.n331 B.n330 10.6151
R896 B.n330 B.n329 10.6151
R897 B.n329 B.n22 10.6151
R898 B.n325 B.n22 10.6151
R899 B.n323 B.n322 10.6151
R900 B.n322 B.n26 10.6151
R901 B.n318 B.n26 10.6151
R902 B.n318 B.n317 10.6151
R903 B.n317 B.n316 10.6151
R904 B.n316 B.n28 10.6151
R905 B.n312 B.n28 10.6151
R906 B.n312 B.n311 10.6151
R907 B.n309 B.n32 10.6151
R908 B.n305 B.n32 10.6151
R909 B.n305 B.n304 10.6151
R910 B.n304 B.n303 10.6151
R911 B.n303 B.n34 10.6151
R912 B.n299 B.n34 10.6151
R913 B.n299 B.n298 10.6151
R914 B.n298 B.n297 10.6151
R915 B.n297 B.n36 10.6151
R916 B.n293 B.n36 10.6151
R917 B.n293 B.n292 10.6151
R918 B.n292 B.n291 10.6151
R919 B.n291 B.n38 10.6151
R920 B.n287 B.n38 10.6151
R921 B.n287 B.n286 10.6151
R922 B.n286 B.n285 10.6151
R923 B.n285 B.n40 10.6151
R924 B.n281 B.n40 10.6151
R925 B.n281 B.n280 10.6151
R926 B.n280 B.n279 10.6151
R927 B.n279 B.n42 10.6151
R928 B.n275 B.n42 10.6151
R929 B.n275 B.n274 10.6151
R930 B.n273 B.n44 10.6151
R931 B.n269 B.n44 10.6151
R932 B.n269 B.n268 10.6151
R933 B.n268 B.n267 10.6151
R934 B.n267 B.n46 10.6151
R935 B.n263 B.n46 10.6151
R936 B.n263 B.n262 10.6151
R937 B.n262 B.n261 10.6151
R938 B.n261 B.n48 10.6151
R939 B.n257 B.n48 10.6151
R940 B.n257 B.n256 10.6151
R941 B.n256 B.n255 10.6151
R942 B.n255 B.n50 10.6151
R943 B.n251 B.n50 10.6151
R944 B.n251 B.n250 10.6151
R945 B.n250 B.n249 10.6151
R946 B.n249 B.n52 10.6151
R947 B.n245 B.n52 10.6151
R948 B.n245 B.n244 10.6151
R949 B.n244 B.n243 10.6151
R950 B.n243 B.n54 10.6151
R951 B.n239 B.n54 10.6151
R952 B.n239 B.n238 10.6151
R953 B.n238 B.n237 10.6151
R954 B.n237 B.n56 10.6151
R955 B.n233 B.n56 10.6151
R956 B.n233 B.n232 10.6151
R957 B.n232 B.n231 10.6151
R958 B.n231 B.n58 10.6151
R959 B.n227 B.n58 10.6151
R960 B.n227 B.n226 10.6151
R961 B.n226 B.n225 10.6151
R962 B.n225 B.n60 10.6151
R963 B.n221 B.n60 10.6151
R964 B.n221 B.n220 10.6151
R965 B.n220 B.n219 10.6151
R966 B.n219 B.n62 10.6151
R967 B.n102 B.n1 10.6151
R968 B.n103 B.n102 10.6151
R969 B.n103 B.n100 10.6151
R970 B.n107 B.n100 10.6151
R971 B.n108 B.n107 10.6151
R972 B.n109 B.n108 10.6151
R973 B.n109 B.n98 10.6151
R974 B.n113 B.n98 10.6151
R975 B.n114 B.n113 10.6151
R976 B.n115 B.n114 10.6151
R977 B.n115 B.n96 10.6151
R978 B.n119 B.n96 10.6151
R979 B.n120 B.n119 10.6151
R980 B.n121 B.n120 10.6151
R981 B.n121 B.n94 10.6151
R982 B.n125 B.n94 10.6151
R983 B.n126 B.n125 10.6151
R984 B.n127 B.n92 10.6151
R985 B.n131 B.n92 10.6151
R986 B.n132 B.n131 10.6151
R987 B.n133 B.n132 10.6151
R988 B.n133 B.n90 10.6151
R989 B.n137 B.n90 10.6151
R990 B.n138 B.n137 10.6151
R991 B.n139 B.n138 10.6151
R992 B.n139 B.n88 10.6151
R993 B.n143 B.n88 10.6151
R994 B.n144 B.n143 10.6151
R995 B.n145 B.n144 10.6151
R996 B.n145 B.n86 10.6151
R997 B.n149 B.n86 10.6151
R998 B.n150 B.n149 10.6151
R999 B.n151 B.n150 10.6151
R1000 B.n151 B.n84 10.6151
R1001 B.n155 B.n84 10.6151
R1002 B.n156 B.n155 10.6151
R1003 B.n157 B.n156 10.6151
R1004 B.n157 B.n82 10.6151
R1005 B.n161 B.n82 10.6151
R1006 B.n162 B.n161 10.6151
R1007 B.n164 B.n78 10.6151
R1008 B.n168 B.n78 10.6151
R1009 B.n169 B.n168 10.6151
R1010 B.n170 B.n169 10.6151
R1011 B.n170 B.n76 10.6151
R1012 B.n174 B.n76 10.6151
R1013 B.n175 B.n174 10.6151
R1014 B.n179 B.n175 10.6151
R1015 B.n183 B.n74 10.6151
R1016 B.n184 B.n183 10.6151
R1017 B.n185 B.n184 10.6151
R1018 B.n185 B.n72 10.6151
R1019 B.n189 B.n72 10.6151
R1020 B.n190 B.n189 10.6151
R1021 B.n191 B.n190 10.6151
R1022 B.n191 B.n70 10.6151
R1023 B.n195 B.n70 10.6151
R1024 B.n196 B.n195 10.6151
R1025 B.n197 B.n196 10.6151
R1026 B.n197 B.n68 10.6151
R1027 B.n201 B.n68 10.6151
R1028 B.n202 B.n201 10.6151
R1029 B.n203 B.n202 10.6151
R1030 B.n203 B.n66 10.6151
R1031 B.n207 B.n66 10.6151
R1032 B.n208 B.n207 10.6151
R1033 B.n209 B.n208 10.6151
R1034 B.n209 B.n64 10.6151
R1035 B.n213 B.n64 10.6151
R1036 B.n214 B.n213 10.6151
R1037 B.n215 B.n214 10.6151
R1038 B.n389 B.n0 8.11757
R1039 B.n389 B.n1 8.11757
R1040 B.n324 B.n323 6.5566
R1041 B.n311 B.n310 6.5566
R1042 B.n164 B.n163 6.5566
R1043 B.n179 B.n178 6.5566
R1044 B.n325 B.n324 4.05904
R1045 B.n310 B.n309 4.05904
R1046 B.n163 B.n162 4.05904
R1047 B.n178 B.n74 4.05904
C0 VTAIL VDD1 6.2486f
C1 VTAIL VN 1.98193f
C2 B VDD2 1.09913f
C3 w_n1674_n2146# VDD2 1.33493f
C4 VDD1 VP 2.17913f
C5 VP VN 3.80386f
C6 VTAIL VDD2 6.28475f
C7 w_n1674_n2146# B 5.13697f
C8 VP VDD2 0.284054f
C9 VDD1 VN 0.147992f
C10 VTAIL B 1.54648f
C11 VTAIL w_n1674_n2146# 1.96521f
C12 VP B 0.999716f
C13 VDD1 VDD2 0.655783f
C14 w_n1674_n2146# VP 2.7686f
C15 VN VDD2 2.04556f
C16 VTAIL VP 1.99631f
C17 VDD1 B 1.07367f
C18 w_n1674_n2146# VDD1 1.31551f
C19 B VN 0.658232f
C20 w_n1674_n2146# VN 2.55788f
C21 VDD2 VSUBS 1.040762f
C22 VDD1 VSUBS 0.894153f
C23 VTAIL VSUBS 0.39338f
C24 VN VSUBS 3.45629f
C25 VP VSUBS 1.066195f
C26 B VSUBS 2.087405f
C27 w_n1674_n2146# VSUBS 44.8565f
C28 B.n0 VSUBS 0.005837f
C29 B.n1 VSUBS 0.005837f
C30 B.n2 VSUBS 0.008633f
C31 B.n3 VSUBS 0.006616f
C32 B.n4 VSUBS 0.006616f
C33 B.n5 VSUBS 0.006616f
C34 B.n6 VSUBS 0.006616f
C35 B.n7 VSUBS 0.006616f
C36 B.n8 VSUBS 0.006616f
C37 B.n9 VSUBS 0.006616f
C38 B.n10 VSUBS 0.006616f
C39 B.n11 VSUBS 0.015487f
C40 B.n12 VSUBS 0.006616f
C41 B.n13 VSUBS 0.006616f
C42 B.n14 VSUBS 0.006616f
C43 B.n15 VSUBS 0.006616f
C44 B.n16 VSUBS 0.006616f
C45 B.n17 VSUBS 0.006616f
C46 B.n18 VSUBS 0.006616f
C47 B.n19 VSUBS 0.006616f
C48 B.n20 VSUBS 0.006616f
C49 B.n21 VSUBS 0.006616f
C50 B.n22 VSUBS 0.006616f
C51 B.n23 VSUBS 0.006616f
C52 B.t10 VSUBS 0.082565f
C53 B.t11 VSUBS 0.09032f
C54 B.t9 VSUBS 0.130311f
C55 B.n24 VSUBS 0.156382f
C56 B.n25 VSUBS 0.13808f
C57 B.n26 VSUBS 0.006616f
C58 B.n27 VSUBS 0.006616f
C59 B.n28 VSUBS 0.006616f
C60 B.n29 VSUBS 0.006616f
C61 B.t1 VSUBS 0.082567f
C62 B.t2 VSUBS 0.090321f
C63 B.t0 VSUBS 0.130311f
C64 B.n30 VSUBS 0.15638f
C65 B.n31 VSUBS 0.138079f
C66 B.n32 VSUBS 0.006616f
C67 B.n33 VSUBS 0.006616f
C68 B.n34 VSUBS 0.006616f
C69 B.n35 VSUBS 0.006616f
C70 B.n36 VSUBS 0.006616f
C71 B.n37 VSUBS 0.006616f
C72 B.n38 VSUBS 0.006616f
C73 B.n39 VSUBS 0.006616f
C74 B.n40 VSUBS 0.006616f
C75 B.n41 VSUBS 0.006616f
C76 B.n42 VSUBS 0.006616f
C77 B.n43 VSUBS 0.015487f
C78 B.n44 VSUBS 0.006616f
C79 B.n45 VSUBS 0.006616f
C80 B.n46 VSUBS 0.006616f
C81 B.n47 VSUBS 0.006616f
C82 B.n48 VSUBS 0.006616f
C83 B.n49 VSUBS 0.006616f
C84 B.n50 VSUBS 0.006616f
C85 B.n51 VSUBS 0.006616f
C86 B.n52 VSUBS 0.006616f
C87 B.n53 VSUBS 0.006616f
C88 B.n54 VSUBS 0.006616f
C89 B.n55 VSUBS 0.006616f
C90 B.n56 VSUBS 0.006616f
C91 B.n57 VSUBS 0.006616f
C92 B.n58 VSUBS 0.006616f
C93 B.n59 VSUBS 0.006616f
C94 B.n60 VSUBS 0.006616f
C95 B.n61 VSUBS 0.006616f
C96 B.n62 VSUBS 0.015487f
C97 B.n63 VSUBS 0.006616f
C98 B.n64 VSUBS 0.006616f
C99 B.n65 VSUBS 0.006616f
C100 B.n66 VSUBS 0.006616f
C101 B.n67 VSUBS 0.006616f
C102 B.n68 VSUBS 0.006616f
C103 B.n69 VSUBS 0.006616f
C104 B.n70 VSUBS 0.006616f
C105 B.n71 VSUBS 0.006616f
C106 B.n72 VSUBS 0.006616f
C107 B.n73 VSUBS 0.006616f
C108 B.n74 VSUBS 0.004573f
C109 B.n75 VSUBS 0.006616f
C110 B.n76 VSUBS 0.006616f
C111 B.n77 VSUBS 0.006616f
C112 B.n78 VSUBS 0.006616f
C113 B.n79 VSUBS 0.006616f
C114 B.t8 VSUBS 0.082565f
C115 B.t7 VSUBS 0.09032f
C116 B.t6 VSUBS 0.130311f
C117 B.n80 VSUBS 0.156382f
C118 B.n81 VSUBS 0.13808f
C119 B.n82 VSUBS 0.006616f
C120 B.n83 VSUBS 0.006616f
C121 B.n84 VSUBS 0.006616f
C122 B.n85 VSUBS 0.006616f
C123 B.n86 VSUBS 0.006616f
C124 B.n87 VSUBS 0.006616f
C125 B.n88 VSUBS 0.006616f
C126 B.n89 VSUBS 0.006616f
C127 B.n90 VSUBS 0.006616f
C128 B.n91 VSUBS 0.006616f
C129 B.n92 VSUBS 0.006616f
C130 B.n93 VSUBS 0.014673f
C131 B.n94 VSUBS 0.006616f
C132 B.n95 VSUBS 0.006616f
C133 B.n96 VSUBS 0.006616f
C134 B.n97 VSUBS 0.006616f
C135 B.n98 VSUBS 0.006616f
C136 B.n99 VSUBS 0.006616f
C137 B.n100 VSUBS 0.006616f
C138 B.n101 VSUBS 0.006616f
C139 B.n102 VSUBS 0.006616f
C140 B.n103 VSUBS 0.006616f
C141 B.n104 VSUBS 0.006616f
C142 B.n105 VSUBS 0.006616f
C143 B.n106 VSUBS 0.006616f
C144 B.n107 VSUBS 0.006616f
C145 B.n108 VSUBS 0.006616f
C146 B.n109 VSUBS 0.006616f
C147 B.n110 VSUBS 0.006616f
C148 B.n111 VSUBS 0.006616f
C149 B.n112 VSUBS 0.006616f
C150 B.n113 VSUBS 0.006616f
C151 B.n114 VSUBS 0.006616f
C152 B.n115 VSUBS 0.006616f
C153 B.n116 VSUBS 0.006616f
C154 B.n117 VSUBS 0.006616f
C155 B.n118 VSUBS 0.006616f
C156 B.n119 VSUBS 0.006616f
C157 B.n120 VSUBS 0.006616f
C158 B.n121 VSUBS 0.006616f
C159 B.n122 VSUBS 0.006616f
C160 B.n123 VSUBS 0.006616f
C161 B.n124 VSUBS 0.006616f
C162 B.n125 VSUBS 0.006616f
C163 B.n126 VSUBS 0.014673f
C164 B.n127 VSUBS 0.015487f
C165 B.n128 VSUBS 0.015487f
C166 B.n129 VSUBS 0.006616f
C167 B.n130 VSUBS 0.006616f
C168 B.n131 VSUBS 0.006616f
C169 B.n132 VSUBS 0.006616f
C170 B.n133 VSUBS 0.006616f
C171 B.n134 VSUBS 0.006616f
C172 B.n135 VSUBS 0.006616f
C173 B.n136 VSUBS 0.006616f
C174 B.n137 VSUBS 0.006616f
C175 B.n138 VSUBS 0.006616f
C176 B.n139 VSUBS 0.006616f
C177 B.n140 VSUBS 0.006616f
C178 B.n141 VSUBS 0.006616f
C179 B.n142 VSUBS 0.006616f
C180 B.n143 VSUBS 0.006616f
C181 B.n144 VSUBS 0.006616f
C182 B.n145 VSUBS 0.006616f
C183 B.n146 VSUBS 0.006616f
C184 B.n147 VSUBS 0.006616f
C185 B.n148 VSUBS 0.006616f
C186 B.n149 VSUBS 0.006616f
C187 B.n150 VSUBS 0.006616f
C188 B.n151 VSUBS 0.006616f
C189 B.n152 VSUBS 0.006616f
C190 B.n153 VSUBS 0.006616f
C191 B.n154 VSUBS 0.006616f
C192 B.n155 VSUBS 0.006616f
C193 B.n156 VSUBS 0.006616f
C194 B.n157 VSUBS 0.006616f
C195 B.n158 VSUBS 0.006616f
C196 B.n159 VSUBS 0.006616f
C197 B.n160 VSUBS 0.006616f
C198 B.n161 VSUBS 0.006616f
C199 B.n162 VSUBS 0.004573f
C200 B.n163 VSUBS 0.015328f
C201 B.n164 VSUBS 0.005351f
C202 B.n165 VSUBS 0.006616f
C203 B.n166 VSUBS 0.006616f
C204 B.n167 VSUBS 0.006616f
C205 B.n168 VSUBS 0.006616f
C206 B.n169 VSUBS 0.006616f
C207 B.n170 VSUBS 0.006616f
C208 B.n171 VSUBS 0.006616f
C209 B.n172 VSUBS 0.006616f
C210 B.n173 VSUBS 0.006616f
C211 B.n174 VSUBS 0.006616f
C212 B.n175 VSUBS 0.006616f
C213 B.t5 VSUBS 0.082567f
C214 B.t4 VSUBS 0.090321f
C215 B.t3 VSUBS 0.130311f
C216 B.n176 VSUBS 0.15638f
C217 B.n177 VSUBS 0.138079f
C218 B.n178 VSUBS 0.015328f
C219 B.n179 VSUBS 0.005351f
C220 B.n180 VSUBS 0.006616f
C221 B.n181 VSUBS 0.006616f
C222 B.n182 VSUBS 0.006616f
C223 B.n183 VSUBS 0.006616f
C224 B.n184 VSUBS 0.006616f
C225 B.n185 VSUBS 0.006616f
C226 B.n186 VSUBS 0.006616f
C227 B.n187 VSUBS 0.006616f
C228 B.n188 VSUBS 0.006616f
C229 B.n189 VSUBS 0.006616f
C230 B.n190 VSUBS 0.006616f
C231 B.n191 VSUBS 0.006616f
C232 B.n192 VSUBS 0.006616f
C233 B.n193 VSUBS 0.006616f
C234 B.n194 VSUBS 0.006616f
C235 B.n195 VSUBS 0.006616f
C236 B.n196 VSUBS 0.006616f
C237 B.n197 VSUBS 0.006616f
C238 B.n198 VSUBS 0.006616f
C239 B.n199 VSUBS 0.006616f
C240 B.n200 VSUBS 0.006616f
C241 B.n201 VSUBS 0.006616f
C242 B.n202 VSUBS 0.006616f
C243 B.n203 VSUBS 0.006616f
C244 B.n204 VSUBS 0.006616f
C245 B.n205 VSUBS 0.006616f
C246 B.n206 VSUBS 0.006616f
C247 B.n207 VSUBS 0.006616f
C248 B.n208 VSUBS 0.006616f
C249 B.n209 VSUBS 0.006616f
C250 B.n210 VSUBS 0.006616f
C251 B.n211 VSUBS 0.006616f
C252 B.n212 VSUBS 0.006616f
C253 B.n213 VSUBS 0.006616f
C254 B.n214 VSUBS 0.006616f
C255 B.n215 VSUBS 0.014673f
C256 B.n216 VSUBS 0.015487f
C257 B.n217 VSUBS 0.014673f
C258 B.n218 VSUBS 0.006616f
C259 B.n219 VSUBS 0.006616f
C260 B.n220 VSUBS 0.006616f
C261 B.n221 VSUBS 0.006616f
C262 B.n222 VSUBS 0.006616f
C263 B.n223 VSUBS 0.006616f
C264 B.n224 VSUBS 0.006616f
C265 B.n225 VSUBS 0.006616f
C266 B.n226 VSUBS 0.006616f
C267 B.n227 VSUBS 0.006616f
C268 B.n228 VSUBS 0.006616f
C269 B.n229 VSUBS 0.006616f
C270 B.n230 VSUBS 0.006616f
C271 B.n231 VSUBS 0.006616f
C272 B.n232 VSUBS 0.006616f
C273 B.n233 VSUBS 0.006616f
C274 B.n234 VSUBS 0.006616f
C275 B.n235 VSUBS 0.006616f
C276 B.n236 VSUBS 0.006616f
C277 B.n237 VSUBS 0.006616f
C278 B.n238 VSUBS 0.006616f
C279 B.n239 VSUBS 0.006616f
C280 B.n240 VSUBS 0.006616f
C281 B.n241 VSUBS 0.006616f
C282 B.n242 VSUBS 0.006616f
C283 B.n243 VSUBS 0.006616f
C284 B.n244 VSUBS 0.006616f
C285 B.n245 VSUBS 0.006616f
C286 B.n246 VSUBS 0.006616f
C287 B.n247 VSUBS 0.006616f
C288 B.n248 VSUBS 0.006616f
C289 B.n249 VSUBS 0.006616f
C290 B.n250 VSUBS 0.006616f
C291 B.n251 VSUBS 0.006616f
C292 B.n252 VSUBS 0.006616f
C293 B.n253 VSUBS 0.006616f
C294 B.n254 VSUBS 0.006616f
C295 B.n255 VSUBS 0.006616f
C296 B.n256 VSUBS 0.006616f
C297 B.n257 VSUBS 0.006616f
C298 B.n258 VSUBS 0.006616f
C299 B.n259 VSUBS 0.006616f
C300 B.n260 VSUBS 0.006616f
C301 B.n261 VSUBS 0.006616f
C302 B.n262 VSUBS 0.006616f
C303 B.n263 VSUBS 0.006616f
C304 B.n264 VSUBS 0.006616f
C305 B.n265 VSUBS 0.006616f
C306 B.n266 VSUBS 0.006616f
C307 B.n267 VSUBS 0.006616f
C308 B.n268 VSUBS 0.006616f
C309 B.n269 VSUBS 0.006616f
C310 B.n270 VSUBS 0.006616f
C311 B.n271 VSUBS 0.006616f
C312 B.n272 VSUBS 0.014673f
C313 B.n273 VSUBS 0.014673f
C314 B.n274 VSUBS 0.015487f
C315 B.n275 VSUBS 0.006616f
C316 B.n276 VSUBS 0.006616f
C317 B.n277 VSUBS 0.006616f
C318 B.n278 VSUBS 0.006616f
C319 B.n279 VSUBS 0.006616f
C320 B.n280 VSUBS 0.006616f
C321 B.n281 VSUBS 0.006616f
C322 B.n282 VSUBS 0.006616f
C323 B.n283 VSUBS 0.006616f
C324 B.n284 VSUBS 0.006616f
C325 B.n285 VSUBS 0.006616f
C326 B.n286 VSUBS 0.006616f
C327 B.n287 VSUBS 0.006616f
C328 B.n288 VSUBS 0.006616f
C329 B.n289 VSUBS 0.006616f
C330 B.n290 VSUBS 0.006616f
C331 B.n291 VSUBS 0.006616f
C332 B.n292 VSUBS 0.006616f
C333 B.n293 VSUBS 0.006616f
C334 B.n294 VSUBS 0.006616f
C335 B.n295 VSUBS 0.006616f
C336 B.n296 VSUBS 0.006616f
C337 B.n297 VSUBS 0.006616f
C338 B.n298 VSUBS 0.006616f
C339 B.n299 VSUBS 0.006616f
C340 B.n300 VSUBS 0.006616f
C341 B.n301 VSUBS 0.006616f
C342 B.n302 VSUBS 0.006616f
C343 B.n303 VSUBS 0.006616f
C344 B.n304 VSUBS 0.006616f
C345 B.n305 VSUBS 0.006616f
C346 B.n306 VSUBS 0.006616f
C347 B.n307 VSUBS 0.006616f
C348 B.n308 VSUBS 0.006616f
C349 B.n309 VSUBS 0.004573f
C350 B.n310 VSUBS 0.015328f
C351 B.n311 VSUBS 0.005351f
C352 B.n312 VSUBS 0.006616f
C353 B.n313 VSUBS 0.006616f
C354 B.n314 VSUBS 0.006616f
C355 B.n315 VSUBS 0.006616f
C356 B.n316 VSUBS 0.006616f
C357 B.n317 VSUBS 0.006616f
C358 B.n318 VSUBS 0.006616f
C359 B.n319 VSUBS 0.006616f
C360 B.n320 VSUBS 0.006616f
C361 B.n321 VSUBS 0.006616f
C362 B.n322 VSUBS 0.006616f
C363 B.n323 VSUBS 0.005351f
C364 B.n324 VSUBS 0.015328f
C365 B.n325 VSUBS 0.004573f
C366 B.n326 VSUBS 0.006616f
C367 B.n327 VSUBS 0.006616f
C368 B.n328 VSUBS 0.006616f
C369 B.n329 VSUBS 0.006616f
C370 B.n330 VSUBS 0.006616f
C371 B.n331 VSUBS 0.006616f
C372 B.n332 VSUBS 0.006616f
C373 B.n333 VSUBS 0.006616f
C374 B.n334 VSUBS 0.006616f
C375 B.n335 VSUBS 0.006616f
C376 B.n336 VSUBS 0.006616f
C377 B.n337 VSUBS 0.006616f
C378 B.n338 VSUBS 0.006616f
C379 B.n339 VSUBS 0.006616f
C380 B.n340 VSUBS 0.006616f
C381 B.n341 VSUBS 0.006616f
C382 B.n342 VSUBS 0.006616f
C383 B.n343 VSUBS 0.006616f
C384 B.n344 VSUBS 0.006616f
C385 B.n345 VSUBS 0.006616f
C386 B.n346 VSUBS 0.006616f
C387 B.n347 VSUBS 0.006616f
C388 B.n348 VSUBS 0.006616f
C389 B.n349 VSUBS 0.006616f
C390 B.n350 VSUBS 0.006616f
C391 B.n351 VSUBS 0.006616f
C392 B.n352 VSUBS 0.006616f
C393 B.n353 VSUBS 0.006616f
C394 B.n354 VSUBS 0.006616f
C395 B.n355 VSUBS 0.006616f
C396 B.n356 VSUBS 0.006616f
C397 B.n357 VSUBS 0.006616f
C398 B.n358 VSUBS 0.006616f
C399 B.n359 VSUBS 0.006616f
C400 B.n360 VSUBS 0.015487f
C401 B.n361 VSUBS 0.014673f
C402 B.n362 VSUBS 0.014673f
C403 B.n363 VSUBS 0.006616f
C404 B.n364 VSUBS 0.006616f
C405 B.n365 VSUBS 0.006616f
C406 B.n366 VSUBS 0.006616f
C407 B.n367 VSUBS 0.006616f
C408 B.n368 VSUBS 0.006616f
C409 B.n369 VSUBS 0.006616f
C410 B.n370 VSUBS 0.006616f
C411 B.n371 VSUBS 0.006616f
C412 B.n372 VSUBS 0.006616f
C413 B.n373 VSUBS 0.006616f
C414 B.n374 VSUBS 0.006616f
C415 B.n375 VSUBS 0.006616f
C416 B.n376 VSUBS 0.006616f
C417 B.n377 VSUBS 0.006616f
C418 B.n378 VSUBS 0.006616f
C419 B.n379 VSUBS 0.006616f
C420 B.n380 VSUBS 0.006616f
C421 B.n381 VSUBS 0.006616f
C422 B.n382 VSUBS 0.006616f
C423 B.n383 VSUBS 0.006616f
C424 B.n384 VSUBS 0.006616f
C425 B.n385 VSUBS 0.006616f
C426 B.n386 VSUBS 0.006616f
C427 B.n387 VSUBS 0.008633f
C428 B.n388 VSUBS 0.009197f
C429 B.n389 VSUBS 0.018288f
C430 VDD2.n0 VSUBS 0.025323f
C431 VDD2.n1 VSUBS 0.024164f
C432 VDD2.n2 VSUBS 0.012984f
C433 VDD2.n3 VSUBS 0.030691f
C434 VDD2.n4 VSUBS 0.013748f
C435 VDD2.n5 VSUBS 0.024164f
C436 VDD2.n6 VSUBS 0.012984f
C437 VDD2.n7 VSUBS 0.030691f
C438 VDD2.n8 VSUBS 0.013748f
C439 VDD2.n9 VSUBS 0.105911f
C440 VDD2.t5 VSUBS 0.065704f
C441 VDD2.n10 VSUBS 0.023018f
C442 VDD2.n11 VSUBS 0.019514f
C443 VDD2.n12 VSUBS 0.012984f
C444 VDD2.n13 VSUBS 0.542515f
C445 VDD2.n14 VSUBS 0.024164f
C446 VDD2.n15 VSUBS 0.012984f
C447 VDD2.n16 VSUBS 0.013748f
C448 VDD2.n17 VSUBS 0.030691f
C449 VDD2.n18 VSUBS 0.030691f
C450 VDD2.n19 VSUBS 0.013748f
C451 VDD2.n20 VSUBS 0.012984f
C452 VDD2.n21 VSUBS 0.024164f
C453 VDD2.n22 VSUBS 0.024164f
C454 VDD2.n23 VSUBS 0.012984f
C455 VDD2.n24 VSUBS 0.013748f
C456 VDD2.n25 VSUBS 0.030691f
C457 VDD2.n26 VSUBS 0.070116f
C458 VDD2.n27 VSUBS 0.013748f
C459 VDD2.n28 VSUBS 0.012984f
C460 VDD2.n29 VSUBS 0.052222f
C461 VDD2.n30 VSUBS 0.052606f
C462 VDD2.t0 VSUBS 0.112468f
C463 VDD2.t3 VSUBS 0.112468f
C464 VDD2.n31 VSUBS 0.738994f
C465 VDD2.n32 VSUBS 1.5695f
C466 VDD2.n33 VSUBS 0.025323f
C467 VDD2.n34 VSUBS 0.024164f
C468 VDD2.n35 VSUBS 0.012984f
C469 VDD2.n36 VSUBS 0.030691f
C470 VDD2.n37 VSUBS 0.013748f
C471 VDD2.n38 VSUBS 0.024164f
C472 VDD2.n39 VSUBS 0.012984f
C473 VDD2.n40 VSUBS 0.030691f
C474 VDD2.n41 VSUBS 0.013748f
C475 VDD2.n42 VSUBS 0.105911f
C476 VDD2.t2 VSUBS 0.065704f
C477 VDD2.n43 VSUBS 0.023018f
C478 VDD2.n44 VSUBS 0.019514f
C479 VDD2.n45 VSUBS 0.012984f
C480 VDD2.n46 VSUBS 0.542515f
C481 VDD2.n47 VSUBS 0.024164f
C482 VDD2.n48 VSUBS 0.012984f
C483 VDD2.n49 VSUBS 0.013748f
C484 VDD2.n50 VSUBS 0.030691f
C485 VDD2.n51 VSUBS 0.030691f
C486 VDD2.n52 VSUBS 0.013748f
C487 VDD2.n53 VSUBS 0.012984f
C488 VDD2.n54 VSUBS 0.024164f
C489 VDD2.n55 VSUBS 0.024164f
C490 VDD2.n56 VSUBS 0.012984f
C491 VDD2.n57 VSUBS 0.013748f
C492 VDD2.n58 VSUBS 0.030691f
C493 VDD2.n59 VSUBS 0.070116f
C494 VDD2.n60 VSUBS 0.013748f
C495 VDD2.n61 VSUBS 0.012984f
C496 VDD2.n62 VSUBS 0.052222f
C497 VDD2.n63 VSUBS 0.051676f
C498 VDD2.n64 VSUBS 1.46367f
C499 VDD2.t1 VSUBS 0.112468f
C500 VDD2.t4 VSUBS 0.112468f
C501 VDD2.n65 VSUBS 0.738973f
C502 VN.t0 VSUBS 0.527055f
C503 VN.n0 VSUBS 0.223023f
C504 VN.t5 VSUBS 0.509005f
C505 VN.n1 VSUBS 0.252232f
C506 VN.t2 VSUBS 0.509005f
C507 VN.n2 VSUBS 0.239954f
C508 VN.n3 VSUBS 0.213474f
C509 VN.t1 VSUBS 0.527055f
C510 VN.n4 VSUBS 0.223023f
C511 VN.t4 VSUBS 0.509005f
C512 VN.n5 VSUBS 0.252232f
C513 VN.t3 VSUBS 0.509005f
C514 VN.n6 VSUBS 0.239954f
C515 VN.n7 VSUBS 1.91059f
C516 VTAIL.t0 VSUBS 0.094335f
C517 VTAIL.t11 VSUBS 0.094335f
C518 VTAIL.n0 VSUBS 0.545242f
C519 VTAIL.n1 VSUBS 0.448038f
C520 VTAIL.n2 VSUBS 0.02124f
C521 VTAIL.n3 VSUBS 0.020268f
C522 VTAIL.n4 VSUBS 0.010891f
C523 VTAIL.n5 VSUBS 0.025742f
C524 VTAIL.n6 VSUBS 0.011532f
C525 VTAIL.n7 VSUBS 0.020268f
C526 VTAIL.n8 VSUBS 0.010891f
C527 VTAIL.n9 VSUBS 0.025742f
C528 VTAIL.n10 VSUBS 0.011532f
C529 VTAIL.n11 VSUBS 0.088836f
C530 VTAIL.t6 VSUBS 0.055111f
C531 VTAIL.n12 VSUBS 0.019307f
C532 VTAIL.n13 VSUBS 0.016367f
C533 VTAIL.n14 VSUBS 0.010891f
C534 VTAIL.n15 VSUBS 0.455047f
C535 VTAIL.n16 VSUBS 0.020268f
C536 VTAIL.n17 VSUBS 0.010891f
C537 VTAIL.n18 VSUBS 0.011532f
C538 VTAIL.n19 VSUBS 0.025742f
C539 VTAIL.n20 VSUBS 0.025742f
C540 VTAIL.n21 VSUBS 0.011532f
C541 VTAIL.n22 VSUBS 0.010891f
C542 VTAIL.n23 VSUBS 0.020268f
C543 VTAIL.n24 VSUBS 0.020268f
C544 VTAIL.n25 VSUBS 0.010891f
C545 VTAIL.n26 VSUBS 0.011532f
C546 VTAIL.n27 VSUBS 0.025742f
C547 VTAIL.n28 VSUBS 0.058812f
C548 VTAIL.n29 VSUBS 0.011532f
C549 VTAIL.n30 VSUBS 0.010891f
C550 VTAIL.n31 VSUBS 0.043802f
C551 VTAIL.n32 VSUBS 0.029323f
C552 VTAIL.n33 VSUBS 0.120592f
C553 VTAIL.t8 VSUBS 0.094335f
C554 VTAIL.t9 VSUBS 0.094335f
C555 VTAIL.n34 VSUBS 0.545242f
C556 VTAIL.n35 VSUBS 1.13194f
C557 VTAIL.t3 VSUBS 0.094335f
C558 VTAIL.t2 VSUBS 0.094335f
C559 VTAIL.n36 VSUBS 0.545246f
C560 VTAIL.n37 VSUBS 1.13194f
C561 VTAIL.n38 VSUBS 0.02124f
C562 VTAIL.n39 VSUBS 0.020268f
C563 VTAIL.n40 VSUBS 0.010891f
C564 VTAIL.n41 VSUBS 0.025742f
C565 VTAIL.n42 VSUBS 0.011532f
C566 VTAIL.n43 VSUBS 0.020268f
C567 VTAIL.n44 VSUBS 0.010891f
C568 VTAIL.n45 VSUBS 0.025742f
C569 VTAIL.n46 VSUBS 0.011532f
C570 VTAIL.n47 VSUBS 0.088836f
C571 VTAIL.t4 VSUBS 0.055111f
C572 VTAIL.n48 VSUBS 0.019307f
C573 VTAIL.n49 VSUBS 0.016367f
C574 VTAIL.n50 VSUBS 0.010891f
C575 VTAIL.n51 VSUBS 0.455047f
C576 VTAIL.n52 VSUBS 0.020268f
C577 VTAIL.n53 VSUBS 0.010891f
C578 VTAIL.n54 VSUBS 0.011532f
C579 VTAIL.n55 VSUBS 0.025742f
C580 VTAIL.n56 VSUBS 0.025742f
C581 VTAIL.n57 VSUBS 0.011532f
C582 VTAIL.n58 VSUBS 0.010891f
C583 VTAIL.n59 VSUBS 0.020268f
C584 VTAIL.n60 VSUBS 0.020268f
C585 VTAIL.n61 VSUBS 0.010891f
C586 VTAIL.n62 VSUBS 0.011532f
C587 VTAIL.n63 VSUBS 0.025742f
C588 VTAIL.n64 VSUBS 0.058812f
C589 VTAIL.n65 VSUBS 0.011532f
C590 VTAIL.n66 VSUBS 0.010891f
C591 VTAIL.n67 VSUBS 0.043802f
C592 VTAIL.n68 VSUBS 0.029323f
C593 VTAIL.n69 VSUBS 0.120592f
C594 VTAIL.t5 VSUBS 0.094335f
C595 VTAIL.t10 VSUBS 0.094335f
C596 VTAIL.n70 VSUBS 0.545246f
C597 VTAIL.n71 VSUBS 0.481392f
C598 VTAIL.n72 VSUBS 0.02124f
C599 VTAIL.n73 VSUBS 0.020268f
C600 VTAIL.n74 VSUBS 0.010891f
C601 VTAIL.n75 VSUBS 0.025742f
C602 VTAIL.n76 VSUBS 0.011532f
C603 VTAIL.n77 VSUBS 0.020268f
C604 VTAIL.n78 VSUBS 0.010891f
C605 VTAIL.n79 VSUBS 0.025742f
C606 VTAIL.n80 VSUBS 0.011532f
C607 VTAIL.n81 VSUBS 0.088836f
C608 VTAIL.t7 VSUBS 0.055111f
C609 VTAIL.n82 VSUBS 0.019307f
C610 VTAIL.n83 VSUBS 0.016367f
C611 VTAIL.n84 VSUBS 0.010891f
C612 VTAIL.n85 VSUBS 0.455047f
C613 VTAIL.n86 VSUBS 0.020268f
C614 VTAIL.n87 VSUBS 0.010891f
C615 VTAIL.n88 VSUBS 0.011532f
C616 VTAIL.n89 VSUBS 0.025742f
C617 VTAIL.n90 VSUBS 0.025742f
C618 VTAIL.n91 VSUBS 0.011532f
C619 VTAIL.n92 VSUBS 0.010891f
C620 VTAIL.n93 VSUBS 0.020268f
C621 VTAIL.n94 VSUBS 0.020268f
C622 VTAIL.n95 VSUBS 0.010891f
C623 VTAIL.n96 VSUBS 0.011532f
C624 VTAIL.n97 VSUBS 0.025742f
C625 VTAIL.n98 VSUBS 0.058812f
C626 VTAIL.n99 VSUBS 0.011532f
C627 VTAIL.n100 VSUBS 0.010891f
C628 VTAIL.n101 VSUBS 0.043802f
C629 VTAIL.n102 VSUBS 0.029323f
C630 VTAIL.n103 VSUBS 0.721597f
C631 VTAIL.n104 VSUBS 0.02124f
C632 VTAIL.n105 VSUBS 0.020268f
C633 VTAIL.n106 VSUBS 0.010891f
C634 VTAIL.n107 VSUBS 0.025742f
C635 VTAIL.n108 VSUBS 0.011532f
C636 VTAIL.n109 VSUBS 0.020268f
C637 VTAIL.n110 VSUBS 0.010891f
C638 VTAIL.n111 VSUBS 0.025742f
C639 VTAIL.n112 VSUBS 0.011532f
C640 VTAIL.n113 VSUBS 0.088836f
C641 VTAIL.t1 VSUBS 0.055111f
C642 VTAIL.n114 VSUBS 0.019307f
C643 VTAIL.n115 VSUBS 0.016367f
C644 VTAIL.n116 VSUBS 0.010891f
C645 VTAIL.n117 VSUBS 0.455047f
C646 VTAIL.n118 VSUBS 0.020268f
C647 VTAIL.n119 VSUBS 0.010891f
C648 VTAIL.n120 VSUBS 0.011532f
C649 VTAIL.n121 VSUBS 0.025742f
C650 VTAIL.n122 VSUBS 0.025742f
C651 VTAIL.n123 VSUBS 0.011532f
C652 VTAIL.n124 VSUBS 0.010891f
C653 VTAIL.n125 VSUBS 0.020268f
C654 VTAIL.n126 VSUBS 0.020268f
C655 VTAIL.n127 VSUBS 0.010891f
C656 VTAIL.n128 VSUBS 0.011532f
C657 VTAIL.n129 VSUBS 0.025742f
C658 VTAIL.n130 VSUBS 0.058812f
C659 VTAIL.n131 VSUBS 0.011532f
C660 VTAIL.n132 VSUBS 0.010891f
C661 VTAIL.n133 VSUBS 0.043802f
C662 VTAIL.n134 VSUBS 0.029323f
C663 VTAIL.n135 VSUBS 0.705411f
C664 VDD1.n0 VSUBS 0.025355f
C665 VDD1.n1 VSUBS 0.024194f
C666 VDD1.n2 VSUBS 0.013001f
C667 VDD1.n3 VSUBS 0.03073f
C668 VDD1.n4 VSUBS 0.013766f
C669 VDD1.n5 VSUBS 0.024194f
C670 VDD1.n6 VSUBS 0.013001f
C671 VDD1.n7 VSUBS 0.03073f
C672 VDD1.n8 VSUBS 0.013766f
C673 VDD1.n9 VSUBS 0.106047f
C674 VDD1.t5 VSUBS 0.065788f
C675 VDD1.n10 VSUBS 0.023047f
C676 VDD1.n11 VSUBS 0.019538f
C677 VDD1.n12 VSUBS 0.013001f
C678 VDD1.n13 VSUBS 0.543211f
C679 VDD1.n14 VSUBS 0.024194f
C680 VDD1.n15 VSUBS 0.013001f
C681 VDD1.n16 VSUBS 0.013766f
C682 VDD1.n17 VSUBS 0.03073f
C683 VDD1.n18 VSUBS 0.03073f
C684 VDD1.n19 VSUBS 0.013766f
C685 VDD1.n20 VSUBS 0.013001f
C686 VDD1.n21 VSUBS 0.024194f
C687 VDD1.n22 VSUBS 0.024194f
C688 VDD1.n23 VSUBS 0.013001f
C689 VDD1.n24 VSUBS 0.013766f
C690 VDD1.n25 VSUBS 0.03073f
C691 VDD1.n26 VSUBS 0.070206f
C692 VDD1.n27 VSUBS 0.013766f
C693 VDD1.n28 VSUBS 0.013001f
C694 VDD1.n29 VSUBS 0.052289f
C695 VDD1.n30 VSUBS 0.052979f
C696 VDD1.n31 VSUBS 0.025355f
C697 VDD1.n32 VSUBS 0.024194f
C698 VDD1.n33 VSUBS 0.013001f
C699 VDD1.n34 VSUBS 0.03073f
C700 VDD1.n35 VSUBS 0.013766f
C701 VDD1.n36 VSUBS 0.024194f
C702 VDD1.n37 VSUBS 0.013001f
C703 VDD1.n38 VSUBS 0.03073f
C704 VDD1.n39 VSUBS 0.013766f
C705 VDD1.n40 VSUBS 0.106047f
C706 VDD1.t0 VSUBS 0.065788f
C707 VDD1.n41 VSUBS 0.023047f
C708 VDD1.n42 VSUBS 0.019538f
C709 VDD1.n43 VSUBS 0.013001f
C710 VDD1.n44 VSUBS 0.543211f
C711 VDD1.n45 VSUBS 0.024194f
C712 VDD1.n46 VSUBS 0.013001f
C713 VDD1.n47 VSUBS 0.013766f
C714 VDD1.n48 VSUBS 0.03073f
C715 VDD1.n49 VSUBS 0.03073f
C716 VDD1.n50 VSUBS 0.013766f
C717 VDD1.n51 VSUBS 0.013001f
C718 VDD1.n52 VSUBS 0.024194f
C719 VDD1.n53 VSUBS 0.024194f
C720 VDD1.n54 VSUBS 0.013001f
C721 VDD1.n55 VSUBS 0.013766f
C722 VDD1.n56 VSUBS 0.03073f
C723 VDD1.n57 VSUBS 0.070206f
C724 VDD1.n58 VSUBS 0.013766f
C725 VDD1.n59 VSUBS 0.013001f
C726 VDD1.n60 VSUBS 0.052289f
C727 VDD1.n61 VSUBS 0.052673f
C728 VDD1.t4 VSUBS 0.112612f
C729 VDD1.t1 VSUBS 0.112612f
C730 VDD1.n62 VSUBS 0.739942f
C731 VDD1.n63 VSUBS 1.64063f
C732 VDD1.t2 VSUBS 0.112612f
C733 VDD1.t3 VSUBS 0.112612f
C734 VDD1.n64 VSUBS 0.739231f
C735 VDD1.n65 VSUBS 1.86538f
C736 VP.n0 VSUBS 0.076149f
C737 VP.t5 VSUBS 0.557198f
C738 VP.n1 VSUBS 0.235778f
C739 VP.t3 VSUBS 0.538116f
C740 VP.t0 VSUBS 0.538116f
C741 VP.n2 VSUBS 0.266658f
C742 VP.n3 VSUBS 0.253678f
C743 VP.n4 VSUBS 1.98192f
C744 VP.n5 VSUBS 1.87677f
C745 VP.t2 VSUBS 0.538116f
C746 VP.n6 VSUBS 0.253678f
C747 VP.t1 VSUBS 0.538116f
C748 VP.n7 VSUBS 0.266658f
C749 VP.t4 VSUBS 0.538116f
C750 VP.n8 VSUBS 0.253678f
C751 VP.n9 VSUBS 0.063455f
.ends

