* NGSPICE file created from diff_pair_sample_0410.ext - technology: sky130A

.subckt diff_pair_sample_0410 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t8 w_n1510_n1244# sky130_fd_pr__pfet_01v8 ad=0.2277 pd=1.71 as=0.5382 ps=3.54 w=1.38 l=0.21
X1 VDD1.t7 VP.t0 VTAIL.t0 w_n1510_n1244# sky130_fd_pr__pfet_01v8 ad=0.2277 pd=1.71 as=0.5382 ps=3.54 w=1.38 l=0.21
X2 VTAIL.t4 VP.t1 VDD1.t6 w_n1510_n1244# sky130_fd_pr__pfet_01v8 ad=0.2277 pd=1.71 as=0.2277 ps=1.71 w=1.38 l=0.21
X3 VDD1.t5 VP.t2 VTAIL.t5 w_n1510_n1244# sky130_fd_pr__pfet_01v8 ad=0.2277 pd=1.71 as=0.5382 ps=3.54 w=1.38 l=0.21
X4 B.t11 B.t9 B.t10 w_n1510_n1244# sky130_fd_pr__pfet_01v8 ad=0.5382 pd=3.54 as=0 ps=0 w=1.38 l=0.21
X5 B.t8 B.t6 B.t7 w_n1510_n1244# sky130_fd_pr__pfet_01v8 ad=0.5382 pd=3.54 as=0 ps=0 w=1.38 l=0.21
X6 VDD2.t6 VN.t1 VTAIL.t9 w_n1510_n1244# sky130_fd_pr__pfet_01v8 ad=0.2277 pd=1.71 as=0.5382 ps=3.54 w=1.38 l=0.21
X7 VTAIL.t14 VN.t2 VDD2.t5 w_n1510_n1244# sky130_fd_pr__pfet_01v8 ad=0.2277 pd=1.71 as=0.2277 ps=1.71 w=1.38 l=0.21
X8 VTAIL.t13 VN.t3 VDD2.t4 w_n1510_n1244# sky130_fd_pr__pfet_01v8 ad=0.2277 pd=1.71 as=0.2277 ps=1.71 w=1.38 l=0.21
X9 B.t5 B.t3 B.t4 w_n1510_n1244# sky130_fd_pr__pfet_01v8 ad=0.5382 pd=3.54 as=0 ps=0 w=1.38 l=0.21
X10 VDD2.t3 VN.t4 VTAIL.t10 w_n1510_n1244# sky130_fd_pr__pfet_01v8 ad=0.2277 pd=1.71 as=0.2277 ps=1.71 w=1.38 l=0.21
X11 VTAIL.t6 VP.t3 VDD1.t4 w_n1510_n1244# sky130_fd_pr__pfet_01v8 ad=0.5382 pd=3.54 as=0.2277 ps=1.71 w=1.38 l=0.21
X12 VDD2.t2 VN.t5 VTAIL.t12 w_n1510_n1244# sky130_fd_pr__pfet_01v8 ad=0.2277 pd=1.71 as=0.2277 ps=1.71 w=1.38 l=0.21
X13 VDD1.t3 VP.t4 VTAIL.t7 w_n1510_n1244# sky130_fd_pr__pfet_01v8 ad=0.2277 pd=1.71 as=0.2277 ps=1.71 w=1.38 l=0.21
X14 VTAIL.t15 VN.t6 VDD2.t1 w_n1510_n1244# sky130_fd_pr__pfet_01v8 ad=0.5382 pd=3.54 as=0.2277 ps=1.71 w=1.38 l=0.21
X15 VTAIL.t11 VN.t7 VDD2.t0 w_n1510_n1244# sky130_fd_pr__pfet_01v8 ad=0.5382 pd=3.54 as=0.2277 ps=1.71 w=1.38 l=0.21
X16 B.t2 B.t0 B.t1 w_n1510_n1244# sky130_fd_pr__pfet_01v8 ad=0.5382 pd=3.54 as=0 ps=0 w=1.38 l=0.21
X17 VTAIL.t1 VP.t5 VDD1.t2 w_n1510_n1244# sky130_fd_pr__pfet_01v8 ad=0.2277 pd=1.71 as=0.2277 ps=1.71 w=1.38 l=0.21
X18 VTAIL.t3 VP.t6 VDD1.t1 w_n1510_n1244# sky130_fd_pr__pfet_01v8 ad=0.5382 pd=3.54 as=0.2277 ps=1.71 w=1.38 l=0.21
X19 VDD1.t0 VP.t7 VTAIL.t2 w_n1510_n1244# sky130_fd_pr__pfet_01v8 ad=0.2277 pd=1.71 as=0.2277 ps=1.71 w=1.38 l=0.21
R0 VN.n5 VN.t0 352.841
R1 VN.n1 VN.t7 352.841
R2 VN.n12 VN.t6 352.841
R3 VN.n8 VN.t1 352.841
R4 VN.n4 VN.t2 307.562
R5 VN.n2 VN.t5 307.562
R6 VN.n11 VN.t4 307.562
R7 VN.n9 VN.t3 307.562
R8 VN.n8 VN.n7 161.489
R9 VN.n1 VN.n0 161.489
R10 VN.n6 VN.n5 161.3
R11 VN.n13 VN.n12 161.3
R12 VN.n10 VN.n7 161.3
R13 VN.n3 VN.n0 161.3
R14 VN.n3 VN.n2 39.4369
R15 VN.n4 VN.n3 39.4369
R16 VN.n11 VN.n10 39.4369
R17 VN.n10 VN.n9 39.4369
R18 VN.n2 VN.n1 33.5944
R19 VN.n5 VN.n4 33.5944
R20 VN.n12 VN.n11 33.5944
R21 VN.n9 VN.n8 33.5944
R22 VN VN.n13 32.116
R23 VN.n13 VN.n7 0.189894
R24 VN.n6 VN.n0 0.189894
R25 VN VN.n6 0.0516364
R26 VTAIL.n11 VTAIL.t6 255.5
R27 VTAIL.n10 VTAIL.t9 255.5
R28 VTAIL.n7 VTAIL.t15 255.5
R29 VTAIL.n15 VTAIL.t8 255.5
R30 VTAIL.n2 VTAIL.t11 255.5
R31 VTAIL.n3 VTAIL.t5 255.5
R32 VTAIL.n6 VTAIL.t3 255.5
R33 VTAIL.n14 VTAIL.t0 255.5
R34 VTAIL.n13 VTAIL.n12 231.946
R35 VTAIL.n9 VTAIL.n8 231.946
R36 VTAIL.n1 VTAIL.n0 231.946
R37 VTAIL.n5 VTAIL.n4 231.946
R38 VTAIL.n0 VTAIL.t12 23.5548
R39 VTAIL.n0 VTAIL.t14 23.5548
R40 VTAIL.n4 VTAIL.t2 23.5548
R41 VTAIL.n4 VTAIL.t4 23.5548
R42 VTAIL.n12 VTAIL.t7 23.5548
R43 VTAIL.n12 VTAIL.t1 23.5548
R44 VTAIL.n8 VTAIL.t10 23.5548
R45 VTAIL.n8 VTAIL.t13 23.5548
R46 VTAIL.n15 VTAIL.n14 14.0221
R47 VTAIL.n7 VTAIL.n6 14.0221
R48 VTAIL.n11 VTAIL.n10 0.470328
R49 VTAIL.n3 VTAIL.n2 0.470328
R50 VTAIL.n9 VTAIL.n7 0.466017
R51 VTAIL.n10 VTAIL.n9 0.466017
R52 VTAIL.n13 VTAIL.n11 0.466017
R53 VTAIL.n14 VTAIL.n13 0.466017
R54 VTAIL.n6 VTAIL.n5 0.466017
R55 VTAIL.n5 VTAIL.n3 0.466017
R56 VTAIL.n2 VTAIL.n1 0.466017
R57 VTAIL VTAIL.n15 0.407828
R58 VTAIL VTAIL.n1 0.0586897
R59 VDD2.n2 VDD2.n1 248.803
R60 VDD2.n2 VDD2.n0 248.803
R61 VDD2 VDD2.n5 248.799
R62 VDD2.n4 VDD2.n3 248.625
R63 VDD2.n4 VDD2.n2 26.9998
R64 VDD2.n5 VDD2.t4 23.5548
R65 VDD2.n5 VDD2.t6 23.5548
R66 VDD2.n3 VDD2.t1 23.5548
R67 VDD2.n3 VDD2.t3 23.5548
R68 VDD2.n1 VDD2.t5 23.5548
R69 VDD2.n1 VDD2.t7 23.5548
R70 VDD2.n0 VDD2.t0 23.5548
R71 VDD2.n0 VDD2.t2 23.5548
R72 VDD2 VDD2.n4 0.291448
R73 VP.n13 VP.t2 352.841
R74 VP.n9 VP.t6 352.841
R75 VP.n2 VP.t3 352.841
R76 VP.n6 VP.t0 352.841
R77 VP.n12 VP.t1 307.562
R78 VP.n10 VP.t7 307.562
R79 VP.n3 VP.t4 307.562
R80 VP.n5 VP.t5 307.562
R81 VP.n2 VP.n1 161.489
R82 VP.n14 VP.n13 161.3
R83 VP.n4 VP.n1 161.3
R84 VP.n7 VP.n6 161.3
R85 VP.n11 VP.n0 161.3
R86 VP.n9 VP.n8 161.3
R87 VP.n11 VP.n10 39.4369
R88 VP.n12 VP.n11 39.4369
R89 VP.n4 VP.n3 39.4369
R90 VP.n5 VP.n4 39.4369
R91 VP.n10 VP.n9 33.5944
R92 VP.n13 VP.n12 33.5944
R93 VP.n3 VP.n2 33.5944
R94 VP.n6 VP.n5 33.5944
R95 VP.n8 VP.n7 31.7353
R96 VP.n7 VP.n1 0.189894
R97 VP.n8 VP.n0 0.189894
R98 VP.n14 VP.n0 0.189894
R99 VP VP.n14 0.0516364
R100 VDD1 VDD1.n0 248.917
R101 VDD1.n3 VDD1.n2 248.803
R102 VDD1.n3 VDD1.n1 248.803
R103 VDD1.n5 VDD1.n4 248.625
R104 VDD1.n5 VDD1.n3 27.5828
R105 VDD1.n4 VDD1.t2 23.5548
R106 VDD1.n4 VDD1.t7 23.5548
R107 VDD1.n0 VDD1.t4 23.5548
R108 VDD1.n0 VDD1.t3 23.5548
R109 VDD1.n2 VDD1.t6 23.5548
R110 VDD1.n2 VDD1.t5 23.5548
R111 VDD1.n1 VDD1.t1 23.5548
R112 VDD1.n1 VDD1.t0 23.5548
R113 VDD1 VDD1.n5 0.175069
R114 B.n192 B.n29 585
R115 B.n194 B.n193 585
R116 B.n195 B.n28 585
R117 B.n197 B.n196 585
R118 B.n198 B.n27 585
R119 B.n200 B.n199 585
R120 B.n201 B.n26 585
R121 B.n203 B.n202 585
R122 B.n204 B.n25 585
R123 B.n206 B.n205 585
R124 B.n208 B.n207 585
R125 B.n209 B.n21 585
R126 B.n211 B.n210 585
R127 B.n212 B.n20 585
R128 B.n214 B.n213 585
R129 B.n215 B.n19 585
R130 B.n217 B.n216 585
R131 B.n218 B.n18 585
R132 B.n220 B.n219 585
R133 B.n221 B.n15 585
R134 B.n224 B.n223 585
R135 B.n225 B.n14 585
R136 B.n227 B.n226 585
R137 B.n228 B.n13 585
R138 B.n230 B.n229 585
R139 B.n231 B.n12 585
R140 B.n233 B.n232 585
R141 B.n234 B.n11 585
R142 B.n236 B.n235 585
R143 B.n237 B.n10 585
R144 B.n191 B.n190 585
R145 B.n189 B.n30 585
R146 B.n188 B.n187 585
R147 B.n186 B.n31 585
R148 B.n185 B.n184 585
R149 B.n183 B.n32 585
R150 B.n182 B.n181 585
R151 B.n180 B.n33 585
R152 B.n179 B.n178 585
R153 B.n177 B.n34 585
R154 B.n176 B.n175 585
R155 B.n174 B.n35 585
R156 B.n173 B.n172 585
R157 B.n171 B.n36 585
R158 B.n170 B.n169 585
R159 B.n168 B.n37 585
R160 B.n167 B.n166 585
R161 B.n165 B.n38 585
R162 B.n164 B.n163 585
R163 B.n162 B.n39 585
R164 B.n161 B.n160 585
R165 B.n159 B.n40 585
R166 B.n158 B.n157 585
R167 B.n156 B.n41 585
R168 B.n155 B.n154 585
R169 B.n153 B.n42 585
R170 B.n152 B.n151 585
R171 B.n150 B.n43 585
R172 B.n149 B.n148 585
R173 B.n147 B.n44 585
R174 B.n146 B.n145 585
R175 B.n144 B.n45 585
R176 B.n143 B.n142 585
R177 B.n96 B.n65 585
R178 B.n98 B.n97 585
R179 B.n99 B.n64 585
R180 B.n101 B.n100 585
R181 B.n102 B.n63 585
R182 B.n104 B.n103 585
R183 B.n105 B.n62 585
R184 B.n107 B.n106 585
R185 B.n108 B.n61 585
R186 B.n110 B.n109 585
R187 B.n112 B.n111 585
R188 B.n113 B.n57 585
R189 B.n115 B.n114 585
R190 B.n116 B.n56 585
R191 B.n118 B.n117 585
R192 B.n119 B.n55 585
R193 B.n121 B.n120 585
R194 B.n122 B.n54 585
R195 B.n124 B.n123 585
R196 B.n125 B.n51 585
R197 B.n128 B.n127 585
R198 B.n129 B.n50 585
R199 B.n131 B.n130 585
R200 B.n132 B.n49 585
R201 B.n134 B.n133 585
R202 B.n135 B.n48 585
R203 B.n137 B.n136 585
R204 B.n138 B.n47 585
R205 B.n140 B.n139 585
R206 B.n141 B.n46 585
R207 B.n95 B.n94 585
R208 B.n93 B.n66 585
R209 B.n92 B.n91 585
R210 B.n90 B.n67 585
R211 B.n89 B.n88 585
R212 B.n87 B.n68 585
R213 B.n86 B.n85 585
R214 B.n84 B.n69 585
R215 B.n83 B.n82 585
R216 B.n81 B.n70 585
R217 B.n80 B.n79 585
R218 B.n78 B.n71 585
R219 B.n77 B.n76 585
R220 B.n75 B.n72 585
R221 B.n74 B.n73 585
R222 B.n2 B.n0 585
R223 B.n261 B.n1 585
R224 B.n260 B.n259 585
R225 B.n258 B.n3 585
R226 B.n257 B.n256 585
R227 B.n255 B.n4 585
R228 B.n254 B.n253 585
R229 B.n252 B.n5 585
R230 B.n251 B.n250 585
R231 B.n249 B.n6 585
R232 B.n248 B.n247 585
R233 B.n246 B.n7 585
R234 B.n245 B.n244 585
R235 B.n243 B.n8 585
R236 B.n242 B.n241 585
R237 B.n240 B.n9 585
R238 B.n239 B.n238 585
R239 B.n263 B.n262 585
R240 B.n94 B.n65 535.745
R241 B.n238 B.n237 535.745
R242 B.n142 B.n141 535.745
R243 B.n190 B.n29 535.745
R244 B.n52 B.t9 391.853
R245 B.n58 B.t6 391.853
R246 B.n16 B.t0 391.853
R247 B.n22 B.t3 391.853
R248 B.n52 B.t11 259.478
R249 B.n22 B.t4 259.478
R250 B.n58 B.t8 259.478
R251 B.n16 B.t1 259.478
R252 B.n53 B.t10 249.005
R253 B.n23 B.t5 249.005
R254 B.n59 B.t7 249.005
R255 B.n17 B.t2 249.005
R256 B.n94 B.n93 163.367
R257 B.n93 B.n92 163.367
R258 B.n92 B.n67 163.367
R259 B.n88 B.n67 163.367
R260 B.n88 B.n87 163.367
R261 B.n87 B.n86 163.367
R262 B.n86 B.n69 163.367
R263 B.n82 B.n69 163.367
R264 B.n82 B.n81 163.367
R265 B.n81 B.n80 163.367
R266 B.n80 B.n71 163.367
R267 B.n76 B.n71 163.367
R268 B.n76 B.n75 163.367
R269 B.n75 B.n74 163.367
R270 B.n74 B.n2 163.367
R271 B.n262 B.n2 163.367
R272 B.n262 B.n261 163.367
R273 B.n261 B.n260 163.367
R274 B.n260 B.n3 163.367
R275 B.n256 B.n3 163.367
R276 B.n256 B.n255 163.367
R277 B.n255 B.n254 163.367
R278 B.n254 B.n5 163.367
R279 B.n250 B.n5 163.367
R280 B.n250 B.n249 163.367
R281 B.n249 B.n248 163.367
R282 B.n248 B.n7 163.367
R283 B.n244 B.n7 163.367
R284 B.n244 B.n243 163.367
R285 B.n243 B.n242 163.367
R286 B.n242 B.n9 163.367
R287 B.n238 B.n9 163.367
R288 B.n98 B.n65 163.367
R289 B.n99 B.n98 163.367
R290 B.n100 B.n99 163.367
R291 B.n100 B.n63 163.367
R292 B.n104 B.n63 163.367
R293 B.n105 B.n104 163.367
R294 B.n106 B.n105 163.367
R295 B.n106 B.n61 163.367
R296 B.n110 B.n61 163.367
R297 B.n111 B.n110 163.367
R298 B.n111 B.n57 163.367
R299 B.n115 B.n57 163.367
R300 B.n116 B.n115 163.367
R301 B.n117 B.n116 163.367
R302 B.n117 B.n55 163.367
R303 B.n121 B.n55 163.367
R304 B.n122 B.n121 163.367
R305 B.n123 B.n122 163.367
R306 B.n123 B.n51 163.367
R307 B.n128 B.n51 163.367
R308 B.n129 B.n128 163.367
R309 B.n130 B.n129 163.367
R310 B.n130 B.n49 163.367
R311 B.n134 B.n49 163.367
R312 B.n135 B.n134 163.367
R313 B.n136 B.n135 163.367
R314 B.n136 B.n47 163.367
R315 B.n140 B.n47 163.367
R316 B.n141 B.n140 163.367
R317 B.n142 B.n45 163.367
R318 B.n146 B.n45 163.367
R319 B.n147 B.n146 163.367
R320 B.n148 B.n147 163.367
R321 B.n148 B.n43 163.367
R322 B.n152 B.n43 163.367
R323 B.n153 B.n152 163.367
R324 B.n154 B.n153 163.367
R325 B.n154 B.n41 163.367
R326 B.n158 B.n41 163.367
R327 B.n159 B.n158 163.367
R328 B.n160 B.n159 163.367
R329 B.n160 B.n39 163.367
R330 B.n164 B.n39 163.367
R331 B.n165 B.n164 163.367
R332 B.n166 B.n165 163.367
R333 B.n166 B.n37 163.367
R334 B.n170 B.n37 163.367
R335 B.n171 B.n170 163.367
R336 B.n172 B.n171 163.367
R337 B.n172 B.n35 163.367
R338 B.n176 B.n35 163.367
R339 B.n177 B.n176 163.367
R340 B.n178 B.n177 163.367
R341 B.n178 B.n33 163.367
R342 B.n182 B.n33 163.367
R343 B.n183 B.n182 163.367
R344 B.n184 B.n183 163.367
R345 B.n184 B.n31 163.367
R346 B.n188 B.n31 163.367
R347 B.n189 B.n188 163.367
R348 B.n190 B.n189 163.367
R349 B.n237 B.n236 163.367
R350 B.n236 B.n11 163.367
R351 B.n232 B.n11 163.367
R352 B.n232 B.n231 163.367
R353 B.n231 B.n230 163.367
R354 B.n230 B.n13 163.367
R355 B.n226 B.n13 163.367
R356 B.n226 B.n225 163.367
R357 B.n225 B.n224 163.367
R358 B.n224 B.n15 163.367
R359 B.n219 B.n15 163.367
R360 B.n219 B.n218 163.367
R361 B.n218 B.n217 163.367
R362 B.n217 B.n19 163.367
R363 B.n213 B.n19 163.367
R364 B.n213 B.n212 163.367
R365 B.n212 B.n211 163.367
R366 B.n211 B.n21 163.367
R367 B.n207 B.n21 163.367
R368 B.n207 B.n206 163.367
R369 B.n206 B.n25 163.367
R370 B.n202 B.n25 163.367
R371 B.n202 B.n201 163.367
R372 B.n201 B.n200 163.367
R373 B.n200 B.n27 163.367
R374 B.n196 B.n27 163.367
R375 B.n196 B.n195 163.367
R376 B.n195 B.n194 163.367
R377 B.n194 B.n29 163.367
R378 B.n126 B.n53 59.5399
R379 B.n60 B.n59 59.5399
R380 B.n222 B.n17 59.5399
R381 B.n24 B.n23 59.5399
R382 B.n239 B.n10 34.8103
R383 B.n192 B.n191 34.8103
R384 B.n143 B.n46 34.8103
R385 B.n96 B.n95 34.8103
R386 B B.n263 18.0485
R387 B.n235 B.n10 10.6151
R388 B.n235 B.n234 10.6151
R389 B.n234 B.n233 10.6151
R390 B.n233 B.n12 10.6151
R391 B.n229 B.n12 10.6151
R392 B.n229 B.n228 10.6151
R393 B.n228 B.n227 10.6151
R394 B.n227 B.n14 10.6151
R395 B.n223 B.n14 10.6151
R396 B.n221 B.n220 10.6151
R397 B.n220 B.n18 10.6151
R398 B.n216 B.n18 10.6151
R399 B.n216 B.n215 10.6151
R400 B.n215 B.n214 10.6151
R401 B.n214 B.n20 10.6151
R402 B.n210 B.n20 10.6151
R403 B.n210 B.n209 10.6151
R404 B.n209 B.n208 10.6151
R405 B.n205 B.n204 10.6151
R406 B.n204 B.n203 10.6151
R407 B.n203 B.n26 10.6151
R408 B.n199 B.n26 10.6151
R409 B.n199 B.n198 10.6151
R410 B.n198 B.n197 10.6151
R411 B.n197 B.n28 10.6151
R412 B.n193 B.n28 10.6151
R413 B.n193 B.n192 10.6151
R414 B.n144 B.n143 10.6151
R415 B.n145 B.n144 10.6151
R416 B.n145 B.n44 10.6151
R417 B.n149 B.n44 10.6151
R418 B.n150 B.n149 10.6151
R419 B.n151 B.n150 10.6151
R420 B.n151 B.n42 10.6151
R421 B.n155 B.n42 10.6151
R422 B.n156 B.n155 10.6151
R423 B.n157 B.n156 10.6151
R424 B.n157 B.n40 10.6151
R425 B.n161 B.n40 10.6151
R426 B.n162 B.n161 10.6151
R427 B.n163 B.n162 10.6151
R428 B.n163 B.n38 10.6151
R429 B.n167 B.n38 10.6151
R430 B.n168 B.n167 10.6151
R431 B.n169 B.n168 10.6151
R432 B.n169 B.n36 10.6151
R433 B.n173 B.n36 10.6151
R434 B.n174 B.n173 10.6151
R435 B.n175 B.n174 10.6151
R436 B.n175 B.n34 10.6151
R437 B.n179 B.n34 10.6151
R438 B.n180 B.n179 10.6151
R439 B.n181 B.n180 10.6151
R440 B.n181 B.n32 10.6151
R441 B.n185 B.n32 10.6151
R442 B.n186 B.n185 10.6151
R443 B.n187 B.n186 10.6151
R444 B.n187 B.n30 10.6151
R445 B.n191 B.n30 10.6151
R446 B.n97 B.n96 10.6151
R447 B.n97 B.n64 10.6151
R448 B.n101 B.n64 10.6151
R449 B.n102 B.n101 10.6151
R450 B.n103 B.n102 10.6151
R451 B.n103 B.n62 10.6151
R452 B.n107 B.n62 10.6151
R453 B.n108 B.n107 10.6151
R454 B.n109 B.n108 10.6151
R455 B.n113 B.n112 10.6151
R456 B.n114 B.n113 10.6151
R457 B.n114 B.n56 10.6151
R458 B.n118 B.n56 10.6151
R459 B.n119 B.n118 10.6151
R460 B.n120 B.n119 10.6151
R461 B.n120 B.n54 10.6151
R462 B.n124 B.n54 10.6151
R463 B.n125 B.n124 10.6151
R464 B.n127 B.n50 10.6151
R465 B.n131 B.n50 10.6151
R466 B.n132 B.n131 10.6151
R467 B.n133 B.n132 10.6151
R468 B.n133 B.n48 10.6151
R469 B.n137 B.n48 10.6151
R470 B.n138 B.n137 10.6151
R471 B.n139 B.n138 10.6151
R472 B.n139 B.n46 10.6151
R473 B.n95 B.n66 10.6151
R474 B.n91 B.n66 10.6151
R475 B.n91 B.n90 10.6151
R476 B.n90 B.n89 10.6151
R477 B.n89 B.n68 10.6151
R478 B.n85 B.n68 10.6151
R479 B.n85 B.n84 10.6151
R480 B.n84 B.n83 10.6151
R481 B.n83 B.n70 10.6151
R482 B.n79 B.n70 10.6151
R483 B.n79 B.n78 10.6151
R484 B.n78 B.n77 10.6151
R485 B.n77 B.n72 10.6151
R486 B.n73 B.n72 10.6151
R487 B.n73 B.n0 10.6151
R488 B.n259 B.n1 10.6151
R489 B.n259 B.n258 10.6151
R490 B.n258 B.n257 10.6151
R491 B.n257 B.n4 10.6151
R492 B.n253 B.n4 10.6151
R493 B.n253 B.n252 10.6151
R494 B.n252 B.n251 10.6151
R495 B.n251 B.n6 10.6151
R496 B.n247 B.n6 10.6151
R497 B.n247 B.n246 10.6151
R498 B.n246 B.n245 10.6151
R499 B.n245 B.n8 10.6151
R500 B.n241 B.n8 10.6151
R501 B.n241 B.n240 10.6151
R502 B.n240 B.n239 10.6151
R503 B.n53 B.n52 10.4732
R504 B.n59 B.n58 10.4732
R505 B.n17 B.n16 10.4732
R506 B.n23 B.n22 10.4732
R507 B.n223 B.n222 9.36635
R508 B.n205 B.n24 9.36635
R509 B.n109 B.n60 9.36635
R510 B.n127 B.n126 9.36635
R511 B.n263 B.n0 2.81026
R512 B.n263 B.n1 2.81026
R513 B.n222 B.n221 1.24928
R514 B.n208 B.n24 1.24928
R515 B.n112 B.n60 1.24928
R516 B.n126 B.n125 1.24928
C0 VN B 0.524249f
C1 w_n1510_n1244# B 3.50419f
C2 VDD2 B 0.654243f
C3 w_n1510_n1244# VN 2.15522f
C4 VDD2 VN 0.616875f
C5 VDD2 w_n1510_n1244# 0.811531f
C6 VTAIL B 0.780376f
C7 VP B 0.827287f
C8 VN VTAIL 0.68762f
C9 w_n1510_n1244# VTAIL 1.4098f
C10 VDD2 VTAIL 3.75581f
C11 VN VP 2.77925f
C12 w_n1510_n1244# VP 2.33768f
C13 VDD2 VP 0.272639f
C14 B VDD1 0.632103f
C15 VTAIL VP 0.701727f
C16 VN VDD1 0.153875f
C17 w_n1510_n1244# VDD1 0.797494f
C18 VDD2 VDD1 0.587463f
C19 VTAIL VDD1 3.71742f
C20 VP VDD1 0.734651f
C21 VDD2 VSUBS 0.670622f
C22 VDD1 VSUBS 0.857061f
C23 VTAIL VSUBS 0.251805f
C24 VN VSUBS 3.04436f
C25 VP VSUBS 0.687723f
C26 B VSUBS 1.372f
C27 w_n1510_n1244# VSUBS 24.117699f
C28 B.n0 VSUBS 0.005961f
C29 B.n1 VSUBS 0.005961f
C30 B.n2 VSUBS 0.009427f
C31 B.n3 VSUBS 0.009427f
C32 B.n4 VSUBS 0.009427f
C33 B.n5 VSUBS 0.009427f
C34 B.n6 VSUBS 0.009427f
C35 B.n7 VSUBS 0.009427f
C36 B.n8 VSUBS 0.009427f
C37 B.n9 VSUBS 0.009427f
C38 B.n10 VSUBS 0.023409f
C39 B.n11 VSUBS 0.009427f
C40 B.n12 VSUBS 0.009427f
C41 B.n13 VSUBS 0.009427f
C42 B.n14 VSUBS 0.009427f
C43 B.n15 VSUBS 0.009427f
C44 B.t2 VSUBS 0.037321f
C45 B.t1 VSUBS 0.039022f
C46 B.t0 VSUBS 0.018894f
C47 B.n16 VSUBS 0.054543f
C48 B.n17 VSUBS 0.055595f
C49 B.n18 VSUBS 0.009427f
C50 B.n19 VSUBS 0.009427f
C51 B.n20 VSUBS 0.009427f
C52 B.n21 VSUBS 0.009427f
C53 B.t5 VSUBS 0.037321f
C54 B.t4 VSUBS 0.039022f
C55 B.t3 VSUBS 0.018894f
C56 B.n22 VSUBS 0.054543f
C57 B.n23 VSUBS 0.055595f
C58 B.n24 VSUBS 0.021842f
C59 B.n25 VSUBS 0.009427f
C60 B.n26 VSUBS 0.009427f
C61 B.n27 VSUBS 0.009427f
C62 B.n28 VSUBS 0.009427f
C63 B.n29 VSUBS 0.023409f
C64 B.n30 VSUBS 0.009427f
C65 B.n31 VSUBS 0.009427f
C66 B.n32 VSUBS 0.009427f
C67 B.n33 VSUBS 0.009427f
C68 B.n34 VSUBS 0.009427f
C69 B.n35 VSUBS 0.009427f
C70 B.n36 VSUBS 0.009427f
C71 B.n37 VSUBS 0.009427f
C72 B.n38 VSUBS 0.009427f
C73 B.n39 VSUBS 0.009427f
C74 B.n40 VSUBS 0.009427f
C75 B.n41 VSUBS 0.009427f
C76 B.n42 VSUBS 0.009427f
C77 B.n43 VSUBS 0.009427f
C78 B.n44 VSUBS 0.009427f
C79 B.n45 VSUBS 0.009427f
C80 B.n46 VSUBS 0.023409f
C81 B.n47 VSUBS 0.009427f
C82 B.n48 VSUBS 0.009427f
C83 B.n49 VSUBS 0.009427f
C84 B.n50 VSUBS 0.009427f
C85 B.n51 VSUBS 0.009427f
C86 B.t10 VSUBS 0.037321f
C87 B.t11 VSUBS 0.039022f
C88 B.t9 VSUBS 0.018894f
C89 B.n52 VSUBS 0.054543f
C90 B.n53 VSUBS 0.055595f
C91 B.n54 VSUBS 0.009427f
C92 B.n55 VSUBS 0.009427f
C93 B.n56 VSUBS 0.009427f
C94 B.n57 VSUBS 0.009427f
C95 B.t7 VSUBS 0.037321f
C96 B.t8 VSUBS 0.039022f
C97 B.t6 VSUBS 0.018894f
C98 B.n58 VSUBS 0.054543f
C99 B.n59 VSUBS 0.055595f
C100 B.n60 VSUBS 0.021842f
C101 B.n61 VSUBS 0.009427f
C102 B.n62 VSUBS 0.009427f
C103 B.n63 VSUBS 0.009427f
C104 B.n64 VSUBS 0.009427f
C105 B.n65 VSUBS 0.023409f
C106 B.n66 VSUBS 0.009427f
C107 B.n67 VSUBS 0.009427f
C108 B.n68 VSUBS 0.009427f
C109 B.n69 VSUBS 0.009427f
C110 B.n70 VSUBS 0.009427f
C111 B.n71 VSUBS 0.009427f
C112 B.n72 VSUBS 0.009427f
C113 B.n73 VSUBS 0.009427f
C114 B.n74 VSUBS 0.009427f
C115 B.n75 VSUBS 0.009427f
C116 B.n76 VSUBS 0.009427f
C117 B.n77 VSUBS 0.009427f
C118 B.n78 VSUBS 0.009427f
C119 B.n79 VSUBS 0.009427f
C120 B.n80 VSUBS 0.009427f
C121 B.n81 VSUBS 0.009427f
C122 B.n82 VSUBS 0.009427f
C123 B.n83 VSUBS 0.009427f
C124 B.n84 VSUBS 0.009427f
C125 B.n85 VSUBS 0.009427f
C126 B.n86 VSUBS 0.009427f
C127 B.n87 VSUBS 0.009427f
C128 B.n88 VSUBS 0.009427f
C129 B.n89 VSUBS 0.009427f
C130 B.n90 VSUBS 0.009427f
C131 B.n91 VSUBS 0.009427f
C132 B.n92 VSUBS 0.009427f
C133 B.n93 VSUBS 0.009427f
C134 B.n94 VSUBS 0.022619f
C135 B.n95 VSUBS 0.022619f
C136 B.n96 VSUBS 0.023409f
C137 B.n97 VSUBS 0.009427f
C138 B.n98 VSUBS 0.009427f
C139 B.n99 VSUBS 0.009427f
C140 B.n100 VSUBS 0.009427f
C141 B.n101 VSUBS 0.009427f
C142 B.n102 VSUBS 0.009427f
C143 B.n103 VSUBS 0.009427f
C144 B.n104 VSUBS 0.009427f
C145 B.n105 VSUBS 0.009427f
C146 B.n106 VSUBS 0.009427f
C147 B.n107 VSUBS 0.009427f
C148 B.n108 VSUBS 0.009427f
C149 B.n109 VSUBS 0.008873f
C150 B.n110 VSUBS 0.009427f
C151 B.n111 VSUBS 0.009427f
C152 B.n112 VSUBS 0.005268f
C153 B.n113 VSUBS 0.009427f
C154 B.n114 VSUBS 0.009427f
C155 B.n115 VSUBS 0.009427f
C156 B.n116 VSUBS 0.009427f
C157 B.n117 VSUBS 0.009427f
C158 B.n118 VSUBS 0.009427f
C159 B.n119 VSUBS 0.009427f
C160 B.n120 VSUBS 0.009427f
C161 B.n121 VSUBS 0.009427f
C162 B.n122 VSUBS 0.009427f
C163 B.n123 VSUBS 0.009427f
C164 B.n124 VSUBS 0.009427f
C165 B.n125 VSUBS 0.005268f
C166 B.n126 VSUBS 0.021842f
C167 B.n127 VSUBS 0.008873f
C168 B.n128 VSUBS 0.009427f
C169 B.n129 VSUBS 0.009427f
C170 B.n130 VSUBS 0.009427f
C171 B.n131 VSUBS 0.009427f
C172 B.n132 VSUBS 0.009427f
C173 B.n133 VSUBS 0.009427f
C174 B.n134 VSUBS 0.009427f
C175 B.n135 VSUBS 0.009427f
C176 B.n136 VSUBS 0.009427f
C177 B.n137 VSUBS 0.009427f
C178 B.n138 VSUBS 0.009427f
C179 B.n139 VSUBS 0.009427f
C180 B.n140 VSUBS 0.009427f
C181 B.n141 VSUBS 0.023409f
C182 B.n142 VSUBS 0.022619f
C183 B.n143 VSUBS 0.022619f
C184 B.n144 VSUBS 0.009427f
C185 B.n145 VSUBS 0.009427f
C186 B.n146 VSUBS 0.009427f
C187 B.n147 VSUBS 0.009427f
C188 B.n148 VSUBS 0.009427f
C189 B.n149 VSUBS 0.009427f
C190 B.n150 VSUBS 0.009427f
C191 B.n151 VSUBS 0.009427f
C192 B.n152 VSUBS 0.009427f
C193 B.n153 VSUBS 0.009427f
C194 B.n154 VSUBS 0.009427f
C195 B.n155 VSUBS 0.009427f
C196 B.n156 VSUBS 0.009427f
C197 B.n157 VSUBS 0.009427f
C198 B.n158 VSUBS 0.009427f
C199 B.n159 VSUBS 0.009427f
C200 B.n160 VSUBS 0.009427f
C201 B.n161 VSUBS 0.009427f
C202 B.n162 VSUBS 0.009427f
C203 B.n163 VSUBS 0.009427f
C204 B.n164 VSUBS 0.009427f
C205 B.n165 VSUBS 0.009427f
C206 B.n166 VSUBS 0.009427f
C207 B.n167 VSUBS 0.009427f
C208 B.n168 VSUBS 0.009427f
C209 B.n169 VSUBS 0.009427f
C210 B.n170 VSUBS 0.009427f
C211 B.n171 VSUBS 0.009427f
C212 B.n172 VSUBS 0.009427f
C213 B.n173 VSUBS 0.009427f
C214 B.n174 VSUBS 0.009427f
C215 B.n175 VSUBS 0.009427f
C216 B.n176 VSUBS 0.009427f
C217 B.n177 VSUBS 0.009427f
C218 B.n178 VSUBS 0.009427f
C219 B.n179 VSUBS 0.009427f
C220 B.n180 VSUBS 0.009427f
C221 B.n181 VSUBS 0.009427f
C222 B.n182 VSUBS 0.009427f
C223 B.n183 VSUBS 0.009427f
C224 B.n184 VSUBS 0.009427f
C225 B.n185 VSUBS 0.009427f
C226 B.n186 VSUBS 0.009427f
C227 B.n187 VSUBS 0.009427f
C228 B.n188 VSUBS 0.009427f
C229 B.n189 VSUBS 0.009427f
C230 B.n190 VSUBS 0.022619f
C231 B.n191 VSUBS 0.023664f
C232 B.n192 VSUBS 0.022364f
C233 B.n193 VSUBS 0.009427f
C234 B.n194 VSUBS 0.009427f
C235 B.n195 VSUBS 0.009427f
C236 B.n196 VSUBS 0.009427f
C237 B.n197 VSUBS 0.009427f
C238 B.n198 VSUBS 0.009427f
C239 B.n199 VSUBS 0.009427f
C240 B.n200 VSUBS 0.009427f
C241 B.n201 VSUBS 0.009427f
C242 B.n202 VSUBS 0.009427f
C243 B.n203 VSUBS 0.009427f
C244 B.n204 VSUBS 0.009427f
C245 B.n205 VSUBS 0.008873f
C246 B.n206 VSUBS 0.009427f
C247 B.n207 VSUBS 0.009427f
C248 B.n208 VSUBS 0.005268f
C249 B.n209 VSUBS 0.009427f
C250 B.n210 VSUBS 0.009427f
C251 B.n211 VSUBS 0.009427f
C252 B.n212 VSUBS 0.009427f
C253 B.n213 VSUBS 0.009427f
C254 B.n214 VSUBS 0.009427f
C255 B.n215 VSUBS 0.009427f
C256 B.n216 VSUBS 0.009427f
C257 B.n217 VSUBS 0.009427f
C258 B.n218 VSUBS 0.009427f
C259 B.n219 VSUBS 0.009427f
C260 B.n220 VSUBS 0.009427f
C261 B.n221 VSUBS 0.005268f
C262 B.n222 VSUBS 0.021842f
C263 B.n223 VSUBS 0.008873f
C264 B.n224 VSUBS 0.009427f
C265 B.n225 VSUBS 0.009427f
C266 B.n226 VSUBS 0.009427f
C267 B.n227 VSUBS 0.009427f
C268 B.n228 VSUBS 0.009427f
C269 B.n229 VSUBS 0.009427f
C270 B.n230 VSUBS 0.009427f
C271 B.n231 VSUBS 0.009427f
C272 B.n232 VSUBS 0.009427f
C273 B.n233 VSUBS 0.009427f
C274 B.n234 VSUBS 0.009427f
C275 B.n235 VSUBS 0.009427f
C276 B.n236 VSUBS 0.009427f
C277 B.n237 VSUBS 0.023409f
C278 B.n238 VSUBS 0.022619f
C279 B.n239 VSUBS 0.022619f
C280 B.n240 VSUBS 0.009427f
C281 B.n241 VSUBS 0.009427f
C282 B.n242 VSUBS 0.009427f
C283 B.n243 VSUBS 0.009427f
C284 B.n244 VSUBS 0.009427f
C285 B.n245 VSUBS 0.009427f
C286 B.n246 VSUBS 0.009427f
C287 B.n247 VSUBS 0.009427f
C288 B.n248 VSUBS 0.009427f
C289 B.n249 VSUBS 0.009427f
C290 B.n250 VSUBS 0.009427f
C291 B.n251 VSUBS 0.009427f
C292 B.n252 VSUBS 0.009427f
C293 B.n253 VSUBS 0.009427f
C294 B.n254 VSUBS 0.009427f
C295 B.n255 VSUBS 0.009427f
C296 B.n256 VSUBS 0.009427f
C297 B.n257 VSUBS 0.009427f
C298 B.n258 VSUBS 0.009427f
C299 B.n259 VSUBS 0.009427f
C300 B.n260 VSUBS 0.009427f
C301 B.n261 VSUBS 0.009427f
C302 B.n262 VSUBS 0.009427f
C303 B.n263 VSUBS 0.021347f
C304 VDD1.t4 VSUBS 0.027895f
C305 VDD1.t3 VSUBS 0.027895f
C306 VDD1.n0 VSUBS 0.106149f
C307 VDD1.t1 VSUBS 0.027895f
C308 VDD1.t0 VSUBS 0.027895f
C309 VDD1.n1 VSUBS 0.106009f
C310 VDD1.t6 VSUBS 0.027895f
C311 VDD1.t5 VSUBS 0.027895f
C312 VDD1.n2 VSUBS 0.106009f
C313 VDD1.n3 VSUBS 1.38557f
C314 VDD1.t2 VSUBS 0.027895f
C315 VDD1.t7 VSUBS 0.027895f
C316 VDD1.n4 VSUBS 0.105802f
C317 VDD1.n5 VSUBS 1.33192f
C318 VP.n0 VSUBS 0.072619f
C319 VP.t1 VSUBS 0.063252f
C320 VP.t7 VSUBS 0.063252f
C321 VP.t6 VSUBS 0.071139f
C322 VP.n1 VSUBS 0.159911f
C323 VP.t5 VSUBS 0.063252f
C324 VP.t4 VSUBS 0.063252f
C325 VP.t3 VSUBS 0.071139f
C326 VP.n2 VSUBS 0.079557f
C327 VP.n3 VSUBS 0.060565f
C328 VP.n4 VSUBS 0.025881f
C329 VP.n5 VSUBS 0.060565f
C330 VP.t0 VSUBS 0.071139f
C331 VP.n6 VSUBS 0.079455f
C332 VP.n7 VSUBS 1.77404f
C333 VP.n8 VSUBS 1.85653f
C334 VP.n9 VSUBS 0.079455f
C335 VP.n10 VSUBS 0.060565f
C336 VP.n11 VSUBS 0.025881f
C337 VP.n12 VSUBS 0.060565f
C338 VP.t2 VSUBS 0.071139f
C339 VP.n13 VSUBS 0.079455f
C340 VP.n14 VSUBS 0.056277f
C341 VDD2.t0 VSUBS 0.029399f
C342 VDD2.t2 VSUBS 0.029399f
C343 VDD2.n0 VSUBS 0.111727f
C344 VDD2.t5 VSUBS 0.029399f
C345 VDD2.t7 VSUBS 0.029399f
C346 VDD2.n1 VSUBS 0.111727f
C347 VDD2.n2 VSUBS 1.40214f
C348 VDD2.t1 VSUBS 0.029399f
C349 VDD2.t3 VSUBS 0.029399f
C350 VDD2.n3 VSUBS 0.111509f
C351 VDD2.n4 VSUBS 1.37246f
C352 VDD2.t4 VSUBS 0.029399f
C353 VDD2.t6 VSUBS 0.029399f
C354 VDD2.n5 VSUBS 0.111721f
C355 VTAIL.t12 VSUBS 0.029528f
C356 VTAIL.t14 VSUBS 0.029528f
C357 VTAIL.n0 VSUBS 0.095264f
C358 VTAIL.n1 VSUBS 0.263494f
C359 VTAIL.t11 VSUBS 0.162312f
C360 VTAIL.n2 VSUBS 0.312893f
C361 VTAIL.t5 VSUBS 0.162312f
C362 VTAIL.n3 VSUBS 0.312893f
C363 VTAIL.t2 VSUBS 0.029528f
C364 VTAIL.t4 VSUBS 0.029528f
C365 VTAIL.n4 VSUBS 0.095264f
C366 VTAIL.n5 VSUBS 0.299033f
C367 VTAIL.t3 VSUBS 0.162312f
C368 VTAIL.n6 VSUBS 0.78413f
C369 VTAIL.t15 VSUBS 0.162312f
C370 VTAIL.n7 VSUBS 0.78413f
C371 VTAIL.t10 VSUBS 0.029528f
C372 VTAIL.t13 VSUBS 0.029528f
C373 VTAIL.n8 VSUBS 0.095264f
C374 VTAIL.n9 VSUBS 0.299033f
C375 VTAIL.t9 VSUBS 0.162312f
C376 VTAIL.n10 VSUBS 0.312893f
C377 VTAIL.t6 VSUBS 0.162312f
C378 VTAIL.n11 VSUBS 0.312893f
C379 VTAIL.t7 VSUBS 0.029528f
C380 VTAIL.t1 VSUBS 0.029528f
C381 VTAIL.n12 VSUBS 0.095264f
C382 VTAIL.n13 VSUBS 0.299033f
C383 VTAIL.t0 VSUBS 0.162312f
C384 VTAIL.n14 VSUBS 0.78413f
C385 VTAIL.t8 VSUBS 0.162312f
C386 VTAIL.n15 VSUBS 0.779053f
C387 VN.n0 VSUBS 0.153699f
C388 VN.t2 VSUBS 0.060795f
C389 VN.t5 VSUBS 0.060795f
C390 VN.t7 VSUBS 0.068375f
C391 VN.n1 VSUBS 0.076467f
C392 VN.n2 VSUBS 0.058213f
C393 VN.n3 VSUBS 0.024876f
C394 VN.n4 VSUBS 0.058213f
C395 VN.t0 VSUBS 0.068375f
C396 VN.n5 VSUBS 0.076368f
C397 VN.n6 VSUBS 0.054091f
C398 VN.n7 VSUBS 0.153699f
C399 VN.t6 VSUBS 0.068375f
C400 VN.t4 VSUBS 0.060795f
C401 VN.t3 VSUBS 0.060795f
C402 VN.t1 VSUBS 0.068375f
C403 VN.n8 VSUBS 0.076467f
C404 VN.n9 VSUBS 0.058213f
C405 VN.n10 VSUBS 0.024876f
C406 VN.n11 VSUBS 0.058213f
C407 VN.n12 VSUBS 0.076368f
C408 VN.n13 VSUBS 1.75188f
.ends

