* NGSPICE file created from diff_pair_sample_1706.ext - technology: sky130A

.subckt diff_pair_sample_1706 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=4.8516 pd=25.66 as=4.8516 ps=25.66 w=12.44 l=0.9
X1 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=4.8516 pd=25.66 as=0 ps=0 w=12.44 l=0.9
X2 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=4.8516 pd=25.66 as=4.8516 ps=25.66 w=12.44 l=0.9
X3 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=4.8516 pd=25.66 as=0 ps=0 w=12.44 l=0.9
X4 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.8516 pd=25.66 as=4.8516 ps=25.66 w=12.44 l=0.9
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.8516 pd=25.66 as=0 ps=0 w=12.44 l=0.9
X6 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.8516 pd=25.66 as=4.8516 ps=25.66 w=12.44 l=0.9
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.8516 pd=25.66 as=0 ps=0 w=12.44 l=0.9
R0 VN VN.t0 578.941
R1 VN VN.t1 538.115
R2 VTAIL.n1 VTAIL.t3 45.9246
R3 VTAIL.n3 VTAIL.t2 45.9245
R4 VTAIL.n0 VTAIL.t1 45.9245
R5 VTAIL.n2 VTAIL.t0 45.9245
R6 VTAIL.n1 VTAIL.n0 25.2289
R7 VTAIL.n3 VTAIL.n2 24.1686
R8 VTAIL.n2 VTAIL.n1 1.0005
R9 VTAIL VTAIL.n0 0.793603
R10 VTAIL VTAIL.n3 0.207397
R11 VDD2.n0 VDD2.t0 99.1248
R12 VDD2.n0 VDD2.t1 62.6032
R13 VDD2 VDD2.n0 0.323776
R14 B.n609 B.n608 585
R15 B.n610 B.n609 585
R16 B.n270 B.n80 585
R17 B.n269 B.n268 585
R18 B.n267 B.n266 585
R19 B.n265 B.n264 585
R20 B.n263 B.n262 585
R21 B.n261 B.n260 585
R22 B.n259 B.n258 585
R23 B.n257 B.n256 585
R24 B.n255 B.n254 585
R25 B.n253 B.n252 585
R26 B.n251 B.n250 585
R27 B.n249 B.n248 585
R28 B.n247 B.n246 585
R29 B.n245 B.n244 585
R30 B.n243 B.n242 585
R31 B.n241 B.n240 585
R32 B.n239 B.n238 585
R33 B.n237 B.n236 585
R34 B.n235 B.n234 585
R35 B.n233 B.n232 585
R36 B.n231 B.n230 585
R37 B.n229 B.n228 585
R38 B.n227 B.n226 585
R39 B.n225 B.n224 585
R40 B.n223 B.n222 585
R41 B.n221 B.n220 585
R42 B.n219 B.n218 585
R43 B.n217 B.n216 585
R44 B.n215 B.n214 585
R45 B.n213 B.n212 585
R46 B.n211 B.n210 585
R47 B.n209 B.n208 585
R48 B.n207 B.n206 585
R49 B.n205 B.n204 585
R50 B.n203 B.n202 585
R51 B.n201 B.n200 585
R52 B.n199 B.n198 585
R53 B.n197 B.n196 585
R54 B.n195 B.n194 585
R55 B.n193 B.n192 585
R56 B.n191 B.n190 585
R57 B.n189 B.n188 585
R58 B.n187 B.n186 585
R59 B.n185 B.n184 585
R60 B.n183 B.n182 585
R61 B.n181 B.n180 585
R62 B.n179 B.n178 585
R63 B.n177 B.n176 585
R64 B.n175 B.n174 585
R65 B.n173 B.n172 585
R66 B.n171 B.n170 585
R67 B.n168 B.n167 585
R68 B.n166 B.n165 585
R69 B.n164 B.n163 585
R70 B.n162 B.n161 585
R71 B.n160 B.n159 585
R72 B.n158 B.n157 585
R73 B.n156 B.n155 585
R74 B.n154 B.n153 585
R75 B.n152 B.n151 585
R76 B.n150 B.n149 585
R77 B.n148 B.n147 585
R78 B.n146 B.n145 585
R79 B.n144 B.n143 585
R80 B.n142 B.n141 585
R81 B.n140 B.n139 585
R82 B.n138 B.n137 585
R83 B.n136 B.n135 585
R84 B.n134 B.n133 585
R85 B.n132 B.n131 585
R86 B.n130 B.n129 585
R87 B.n128 B.n127 585
R88 B.n126 B.n125 585
R89 B.n124 B.n123 585
R90 B.n122 B.n121 585
R91 B.n120 B.n119 585
R92 B.n118 B.n117 585
R93 B.n116 B.n115 585
R94 B.n114 B.n113 585
R95 B.n112 B.n111 585
R96 B.n110 B.n109 585
R97 B.n108 B.n107 585
R98 B.n106 B.n105 585
R99 B.n104 B.n103 585
R100 B.n102 B.n101 585
R101 B.n100 B.n99 585
R102 B.n98 B.n97 585
R103 B.n96 B.n95 585
R104 B.n94 B.n93 585
R105 B.n92 B.n91 585
R106 B.n90 B.n89 585
R107 B.n88 B.n87 585
R108 B.n33 B.n32 585
R109 B.n613 B.n612 585
R110 B.n607 B.n81 585
R111 B.n81 B.n30 585
R112 B.n606 B.n29 585
R113 B.n617 B.n29 585
R114 B.n605 B.n28 585
R115 B.n618 B.n28 585
R116 B.n604 B.n27 585
R117 B.n619 B.n27 585
R118 B.n603 B.n602 585
R119 B.n602 B.n23 585
R120 B.n601 B.n22 585
R121 B.n625 B.n22 585
R122 B.n600 B.n21 585
R123 B.n626 B.n21 585
R124 B.n599 B.n20 585
R125 B.n627 B.n20 585
R126 B.n598 B.n597 585
R127 B.n597 B.n16 585
R128 B.n596 B.n15 585
R129 B.n633 B.n15 585
R130 B.n595 B.n14 585
R131 B.n634 B.n14 585
R132 B.n594 B.n13 585
R133 B.n635 B.n13 585
R134 B.n593 B.n592 585
R135 B.n592 B.n12 585
R136 B.n591 B.n590 585
R137 B.n591 B.n8 585
R138 B.n589 B.n7 585
R139 B.n642 B.n7 585
R140 B.n588 B.n6 585
R141 B.n643 B.n6 585
R142 B.n587 B.n5 585
R143 B.n644 B.n5 585
R144 B.n586 B.n585 585
R145 B.n585 B.n4 585
R146 B.n584 B.n271 585
R147 B.n584 B.n583 585
R148 B.n573 B.n272 585
R149 B.n576 B.n272 585
R150 B.n575 B.n574 585
R151 B.n577 B.n575 585
R152 B.n572 B.n277 585
R153 B.n277 B.n276 585
R154 B.n571 B.n570 585
R155 B.n570 B.n569 585
R156 B.n279 B.n278 585
R157 B.n280 B.n279 585
R158 B.n562 B.n561 585
R159 B.n563 B.n562 585
R160 B.n560 B.n285 585
R161 B.n285 B.n284 585
R162 B.n559 B.n558 585
R163 B.n558 B.n557 585
R164 B.n287 B.n286 585
R165 B.n288 B.n287 585
R166 B.n550 B.n549 585
R167 B.n551 B.n550 585
R168 B.n548 B.n293 585
R169 B.n293 B.n292 585
R170 B.n547 B.n546 585
R171 B.n546 B.n545 585
R172 B.n295 B.n294 585
R173 B.n296 B.n295 585
R174 B.n541 B.n540 585
R175 B.n299 B.n298 585
R176 B.n537 B.n536 585
R177 B.n538 B.n537 585
R178 B.n535 B.n346 585
R179 B.n534 B.n533 585
R180 B.n532 B.n531 585
R181 B.n530 B.n529 585
R182 B.n528 B.n527 585
R183 B.n526 B.n525 585
R184 B.n524 B.n523 585
R185 B.n522 B.n521 585
R186 B.n520 B.n519 585
R187 B.n518 B.n517 585
R188 B.n516 B.n515 585
R189 B.n514 B.n513 585
R190 B.n512 B.n511 585
R191 B.n510 B.n509 585
R192 B.n508 B.n507 585
R193 B.n506 B.n505 585
R194 B.n504 B.n503 585
R195 B.n502 B.n501 585
R196 B.n500 B.n499 585
R197 B.n498 B.n497 585
R198 B.n496 B.n495 585
R199 B.n494 B.n493 585
R200 B.n492 B.n491 585
R201 B.n490 B.n489 585
R202 B.n488 B.n487 585
R203 B.n486 B.n485 585
R204 B.n484 B.n483 585
R205 B.n482 B.n481 585
R206 B.n480 B.n479 585
R207 B.n478 B.n477 585
R208 B.n476 B.n475 585
R209 B.n474 B.n473 585
R210 B.n472 B.n471 585
R211 B.n470 B.n469 585
R212 B.n468 B.n467 585
R213 B.n466 B.n465 585
R214 B.n464 B.n463 585
R215 B.n462 B.n461 585
R216 B.n460 B.n459 585
R217 B.n458 B.n457 585
R218 B.n456 B.n455 585
R219 B.n454 B.n453 585
R220 B.n452 B.n451 585
R221 B.n450 B.n449 585
R222 B.n448 B.n447 585
R223 B.n446 B.n445 585
R224 B.n444 B.n443 585
R225 B.n442 B.n441 585
R226 B.n440 B.n439 585
R227 B.n437 B.n436 585
R228 B.n435 B.n434 585
R229 B.n433 B.n432 585
R230 B.n431 B.n430 585
R231 B.n429 B.n428 585
R232 B.n427 B.n426 585
R233 B.n425 B.n424 585
R234 B.n423 B.n422 585
R235 B.n421 B.n420 585
R236 B.n419 B.n418 585
R237 B.n417 B.n416 585
R238 B.n415 B.n414 585
R239 B.n413 B.n412 585
R240 B.n411 B.n410 585
R241 B.n409 B.n408 585
R242 B.n407 B.n406 585
R243 B.n405 B.n404 585
R244 B.n403 B.n402 585
R245 B.n401 B.n400 585
R246 B.n399 B.n398 585
R247 B.n397 B.n396 585
R248 B.n395 B.n394 585
R249 B.n393 B.n392 585
R250 B.n391 B.n390 585
R251 B.n389 B.n388 585
R252 B.n387 B.n386 585
R253 B.n385 B.n384 585
R254 B.n383 B.n382 585
R255 B.n381 B.n380 585
R256 B.n379 B.n378 585
R257 B.n377 B.n376 585
R258 B.n375 B.n374 585
R259 B.n373 B.n372 585
R260 B.n371 B.n370 585
R261 B.n369 B.n368 585
R262 B.n367 B.n366 585
R263 B.n365 B.n364 585
R264 B.n363 B.n362 585
R265 B.n361 B.n360 585
R266 B.n359 B.n358 585
R267 B.n357 B.n356 585
R268 B.n355 B.n354 585
R269 B.n353 B.n352 585
R270 B.n542 B.n297 585
R271 B.n297 B.n296 585
R272 B.n544 B.n543 585
R273 B.n545 B.n544 585
R274 B.n291 B.n290 585
R275 B.n292 B.n291 585
R276 B.n553 B.n552 585
R277 B.n552 B.n551 585
R278 B.n554 B.n289 585
R279 B.n289 B.n288 585
R280 B.n556 B.n555 585
R281 B.n557 B.n556 585
R282 B.n283 B.n282 585
R283 B.n284 B.n283 585
R284 B.n565 B.n564 585
R285 B.n564 B.n563 585
R286 B.n566 B.n281 585
R287 B.n281 B.n280 585
R288 B.n568 B.n567 585
R289 B.n569 B.n568 585
R290 B.n275 B.n274 585
R291 B.n276 B.n275 585
R292 B.n579 B.n578 585
R293 B.n578 B.n577 585
R294 B.n580 B.n273 585
R295 B.n576 B.n273 585
R296 B.n582 B.n581 585
R297 B.n583 B.n582 585
R298 B.n3 B.n0 585
R299 B.n4 B.n3 585
R300 B.n641 B.n1 585
R301 B.n642 B.n641 585
R302 B.n640 B.n639 585
R303 B.n640 B.n8 585
R304 B.n638 B.n9 585
R305 B.n12 B.n9 585
R306 B.n637 B.n636 585
R307 B.n636 B.n635 585
R308 B.n11 B.n10 585
R309 B.n634 B.n11 585
R310 B.n632 B.n631 585
R311 B.n633 B.n632 585
R312 B.n630 B.n17 585
R313 B.n17 B.n16 585
R314 B.n629 B.n628 585
R315 B.n628 B.n627 585
R316 B.n19 B.n18 585
R317 B.n626 B.n19 585
R318 B.n624 B.n623 585
R319 B.n625 B.n624 585
R320 B.n622 B.n24 585
R321 B.n24 B.n23 585
R322 B.n621 B.n620 585
R323 B.n620 B.n619 585
R324 B.n26 B.n25 585
R325 B.n618 B.n26 585
R326 B.n616 B.n615 585
R327 B.n617 B.n616 585
R328 B.n614 B.n31 585
R329 B.n31 B.n30 585
R330 B.n645 B.n644 585
R331 B.n643 B.n2 585
R332 B.n85 B.t6 535.312
R333 B.n82 B.t13 535.312
R334 B.n350 B.t2 535.312
R335 B.n347 B.t10 535.312
R336 B.n612 B.n31 516.524
R337 B.n609 B.n81 516.524
R338 B.n352 B.n295 516.524
R339 B.n540 B.n297 516.524
R340 B.n610 B.n79 256.663
R341 B.n610 B.n78 256.663
R342 B.n610 B.n77 256.663
R343 B.n610 B.n76 256.663
R344 B.n610 B.n75 256.663
R345 B.n610 B.n74 256.663
R346 B.n610 B.n73 256.663
R347 B.n610 B.n72 256.663
R348 B.n610 B.n71 256.663
R349 B.n610 B.n70 256.663
R350 B.n610 B.n69 256.663
R351 B.n610 B.n68 256.663
R352 B.n610 B.n67 256.663
R353 B.n610 B.n66 256.663
R354 B.n610 B.n65 256.663
R355 B.n610 B.n64 256.663
R356 B.n610 B.n63 256.663
R357 B.n610 B.n62 256.663
R358 B.n610 B.n61 256.663
R359 B.n610 B.n60 256.663
R360 B.n610 B.n59 256.663
R361 B.n610 B.n58 256.663
R362 B.n610 B.n57 256.663
R363 B.n610 B.n56 256.663
R364 B.n610 B.n55 256.663
R365 B.n610 B.n54 256.663
R366 B.n610 B.n53 256.663
R367 B.n610 B.n52 256.663
R368 B.n610 B.n51 256.663
R369 B.n610 B.n50 256.663
R370 B.n610 B.n49 256.663
R371 B.n610 B.n48 256.663
R372 B.n610 B.n47 256.663
R373 B.n610 B.n46 256.663
R374 B.n610 B.n45 256.663
R375 B.n610 B.n44 256.663
R376 B.n610 B.n43 256.663
R377 B.n610 B.n42 256.663
R378 B.n610 B.n41 256.663
R379 B.n610 B.n40 256.663
R380 B.n610 B.n39 256.663
R381 B.n610 B.n38 256.663
R382 B.n610 B.n37 256.663
R383 B.n610 B.n36 256.663
R384 B.n610 B.n35 256.663
R385 B.n610 B.n34 256.663
R386 B.n611 B.n610 256.663
R387 B.n539 B.n538 256.663
R388 B.n538 B.n300 256.663
R389 B.n538 B.n301 256.663
R390 B.n538 B.n302 256.663
R391 B.n538 B.n303 256.663
R392 B.n538 B.n304 256.663
R393 B.n538 B.n305 256.663
R394 B.n538 B.n306 256.663
R395 B.n538 B.n307 256.663
R396 B.n538 B.n308 256.663
R397 B.n538 B.n309 256.663
R398 B.n538 B.n310 256.663
R399 B.n538 B.n311 256.663
R400 B.n538 B.n312 256.663
R401 B.n538 B.n313 256.663
R402 B.n538 B.n314 256.663
R403 B.n538 B.n315 256.663
R404 B.n538 B.n316 256.663
R405 B.n538 B.n317 256.663
R406 B.n538 B.n318 256.663
R407 B.n538 B.n319 256.663
R408 B.n538 B.n320 256.663
R409 B.n538 B.n321 256.663
R410 B.n538 B.n322 256.663
R411 B.n538 B.n323 256.663
R412 B.n538 B.n324 256.663
R413 B.n538 B.n325 256.663
R414 B.n538 B.n326 256.663
R415 B.n538 B.n327 256.663
R416 B.n538 B.n328 256.663
R417 B.n538 B.n329 256.663
R418 B.n538 B.n330 256.663
R419 B.n538 B.n331 256.663
R420 B.n538 B.n332 256.663
R421 B.n538 B.n333 256.663
R422 B.n538 B.n334 256.663
R423 B.n538 B.n335 256.663
R424 B.n538 B.n336 256.663
R425 B.n538 B.n337 256.663
R426 B.n538 B.n338 256.663
R427 B.n538 B.n339 256.663
R428 B.n538 B.n340 256.663
R429 B.n538 B.n341 256.663
R430 B.n538 B.n342 256.663
R431 B.n538 B.n343 256.663
R432 B.n538 B.n344 256.663
R433 B.n538 B.n345 256.663
R434 B.n647 B.n646 256.663
R435 B.n87 B.n33 163.367
R436 B.n91 B.n90 163.367
R437 B.n95 B.n94 163.367
R438 B.n99 B.n98 163.367
R439 B.n103 B.n102 163.367
R440 B.n107 B.n106 163.367
R441 B.n111 B.n110 163.367
R442 B.n115 B.n114 163.367
R443 B.n119 B.n118 163.367
R444 B.n123 B.n122 163.367
R445 B.n127 B.n126 163.367
R446 B.n131 B.n130 163.367
R447 B.n135 B.n134 163.367
R448 B.n139 B.n138 163.367
R449 B.n143 B.n142 163.367
R450 B.n147 B.n146 163.367
R451 B.n151 B.n150 163.367
R452 B.n155 B.n154 163.367
R453 B.n159 B.n158 163.367
R454 B.n163 B.n162 163.367
R455 B.n167 B.n166 163.367
R456 B.n172 B.n171 163.367
R457 B.n176 B.n175 163.367
R458 B.n180 B.n179 163.367
R459 B.n184 B.n183 163.367
R460 B.n188 B.n187 163.367
R461 B.n192 B.n191 163.367
R462 B.n196 B.n195 163.367
R463 B.n200 B.n199 163.367
R464 B.n204 B.n203 163.367
R465 B.n208 B.n207 163.367
R466 B.n212 B.n211 163.367
R467 B.n216 B.n215 163.367
R468 B.n220 B.n219 163.367
R469 B.n224 B.n223 163.367
R470 B.n228 B.n227 163.367
R471 B.n232 B.n231 163.367
R472 B.n236 B.n235 163.367
R473 B.n240 B.n239 163.367
R474 B.n244 B.n243 163.367
R475 B.n248 B.n247 163.367
R476 B.n252 B.n251 163.367
R477 B.n256 B.n255 163.367
R478 B.n260 B.n259 163.367
R479 B.n264 B.n263 163.367
R480 B.n268 B.n267 163.367
R481 B.n609 B.n80 163.367
R482 B.n546 B.n295 163.367
R483 B.n546 B.n293 163.367
R484 B.n550 B.n293 163.367
R485 B.n550 B.n287 163.367
R486 B.n558 B.n287 163.367
R487 B.n558 B.n285 163.367
R488 B.n562 B.n285 163.367
R489 B.n562 B.n279 163.367
R490 B.n570 B.n279 163.367
R491 B.n570 B.n277 163.367
R492 B.n575 B.n277 163.367
R493 B.n575 B.n272 163.367
R494 B.n584 B.n272 163.367
R495 B.n585 B.n584 163.367
R496 B.n585 B.n5 163.367
R497 B.n6 B.n5 163.367
R498 B.n7 B.n6 163.367
R499 B.n591 B.n7 163.367
R500 B.n592 B.n591 163.367
R501 B.n592 B.n13 163.367
R502 B.n14 B.n13 163.367
R503 B.n15 B.n14 163.367
R504 B.n597 B.n15 163.367
R505 B.n597 B.n20 163.367
R506 B.n21 B.n20 163.367
R507 B.n22 B.n21 163.367
R508 B.n602 B.n22 163.367
R509 B.n602 B.n27 163.367
R510 B.n28 B.n27 163.367
R511 B.n29 B.n28 163.367
R512 B.n81 B.n29 163.367
R513 B.n537 B.n299 163.367
R514 B.n537 B.n346 163.367
R515 B.n533 B.n532 163.367
R516 B.n529 B.n528 163.367
R517 B.n525 B.n524 163.367
R518 B.n521 B.n520 163.367
R519 B.n517 B.n516 163.367
R520 B.n513 B.n512 163.367
R521 B.n509 B.n508 163.367
R522 B.n505 B.n504 163.367
R523 B.n501 B.n500 163.367
R524 B.n497 B.n496 163.367
R525 B.n493 B.n492 163.367
R526 B.n489 B.n488 163.367
R527 B.n485 B.n484 163.367
R528 B.n481 B.n480 163.367
R529 B.n477 B.n476 163.367
R530 B.n473 B.n472 163.367
R531 B.n469 B.n468 163.367
R532 B.n465 B.n464 163.367
R533 B.n461 B.n460 163.367
R534 B.n457 B.n456 163.367
R535 B.n453 B.n452 163.367
R536 B.n449 B.n448 163.367
R537 B.n445 B.n444 163.367
R538 B.n441 B.n440 163.367
R539 B.n436 B.n435 163.367
R540 B.n432 B.n431 163.367
R541 B.n428 B.n427 163.367
R542 B.n424 B.n423 163.367
R543 B.n420 B.n419 163.367
R544 B.n416 B.n415 163.367
R545 B.n412 B.n411 163.367
R546 B.n408 B.n407 163.367
R547 B.n404 B.n403 163.367
R548 B.n400 B.n399 163.367
R549 B.n396 B.n395 163.367
R550 B.n392 B.n391 163.367
R551 B.n388 B.n387 163.367
R552 B.n384 B.n383 163.367
R553 B.n380 B.n379 163.367
R554 B.n376 B.n375 163.367
R555 B.n372 B.n371 163.367
R556 B.n368 B.n367 163.367
R557 B.n364 B.n363 163.367
R558 B.n360 B.n359 163.367
R559 B.n356 B.n355 163.367
R560 B.n544 B.n297 163.367
R561 B.n544 B.n291 163.367
R562 B.n552 B.n291 163.367
R563 B.n552 B.n289 163.367
R564 B.n556 B.n289 163.367
R565 B.n556 B.n283 163.367
R566 B.n564 B.n283 163.367
R567 B.n564 B.n281 163.367
R568 B.n568 B.n281 163.367
R569 B.n568 B.n275 163.367
R570 B.n578 B.n275 163.367
R571 B.n578 B.n273 163.367
R572 B.n582 B.n273 163.367
R573 B.n582 B.n3 163.367
R574 B.n645 B.n3 163.367
R575 B.n641 B.n2 163.367
R576 B.n641 B.n640 163.367
R577 B.n640 B.n9 163.367
R578 B.n636 B.n9 163.367
R579 B.n636 B.n11 163.367
R580 B.n632 B.n11 163.367
R581 B.n632 B.n17 163.367
R582 B.n628 B.n17 163.367
R583 B.n628 B.n19 163.367
R584 B.n624 B.n19 163.367
R585 B.n624 B.n24 163.367
R586 B.n620 B.n24 163.367
R587 B.n620 B.n26 163.367
R588 B.n616 B.n26 163.367
R589 B.n616 B.n31 163.367
R590 B.n82 B.t14 95.4654
R591 B.n350 B.t5 95.4654
R592 B.n85 B.t8 95.4496
R593 B.n347 B.t12 95.4496
R594 B.n612 B.n611 71.676
R595 B.n87 B.n34 71.676
R596 B.n91 B.n35 71.676
R597 B.n95 B.n36 71.676
R598 B.n99 B.n37 71.676
R599 B.n103 B.n38 71.676
R600 B.n107 B.n39 71.676
R601 B.n111 B.n40 71.676
R602 B.n115 B.n41 71.676
R603 B.n119 B.n42 71.676
R604 B.n123 B.n43 71.676
R605 B.n127 B.n44 71.676
R606 B.n131 B.n45 71.676
R607 B.n135 B.n46 71.676
R608 B.n139 B.n47 71.676
R609 B.n143 B.n48 71.676
R610 B.n147 B.n49 71.676
R611 B.n151 B.n50 71.676
R612 B.n155 B.n51 71.676
R613 B.n159 B.n52 71.676
R614 B.n163 B.n53 71.676
R615 B.n167 B.n54 71.676
R616 B.n172 B.n55 71.676
R617 B.n176 B.n56 71.676
R618 B.n180 B.n57 71.676
R619 B.n184 B.n58 71.676
R620 B.n188 B.n59 71.676
R621 B.n192 B.n60 71.676
R622 B.n196 B.n61 71.676
R623 B.n200 B.n62 71.676
R624 B.n204 B.n63 71.676
R625 B.n208 B.n64 71.676
R626 B.n212 B.n65 71.676
R627 B.n216 B.n66 71.676
R628 B.n220 B.n67 71.676
R629 B.n224 B.n68 71.676
R630 B.n228 B.n69 71.676
R631 B.n232 B.n70 71.676
R632 B.n236 B.n71 71.676
R633 B.n240 B.n72 71.676
R634 B.n244 B.n73 71.676
R635 B.n248 B.n74 71.676
R636 B.n252 B.n75 71.676
R637 B.n256 B.n76 71.676
R638 B.n260 B.n77 71.676
R639 B.n264 B.n78 71.676
R640 B.n268 B.n79 71.676
R641 B.n80 B.n79 71.676
R642 B.n267 B.n78 71.676
R643 B.n263 B.n77 71.676
R644 B.n259 B.n76 71.676
R645 B.n255 B.n75 71.676
R646 B.n251 B.n74 71.676
R647 B.n247 B.n73 71.676
R648 B.n243 B.n72 71.676
R649 B.n239 B.n71 71.676
R650 B.n235 B.n70 71.676
R651 B.n231 B.n69 71.676
R652 B.n227 B.n68 71.676
R653 B.n223 B.n67 71.676
R654 B.n219 B.n66 71.676
R655 B.n215 B.n65 71.676
R656 B.n211 B.n64 71.676
R657 B.n207 B.n63 71.676
R658 B.n203 B.n62 71.676
R659 B.n199 B.n61 71.676
R660 B.n195 B.n60 71.676
R661 B.n191 B.n59 71.676
R662 B.n187 B.n58 71.676
R663 B.n183 B.n57 71.676
R664 B.n179 B.n56 71.676
R665 B.n175 B.n55 71.676
R666 B.n171 B.n54 71.676
R667 B.n166 B.n53 71.676
R668 B.n162 B.n52 71.676
R669 B.n158 B.n51 71.676
R670 B.n154 B.n50 71.676
R671 B.n150 B.n49 71.676
R672 B.n146 B.n48 71.676
R673 B.n142 B.n47 71.676
R674 B.n138 B.n46 71.676
R675 B.n134 B.n45 71.676
R676 B.n130 B.n44 71.676
R677 B.n126 B.n43 71.676
R678 B.n122 B.n42 71.676
R679 B.n118 B.n41 71.676
R680 B.n114 B.n40 71.676
R681 B.n110 B.n39 71.676
R682 B.n106 B.n38 71.676
R683 B.n102 B.n37 71.676
R684 B.n98 B.n36 71.676
R685 B.n94 B.n35 71.676
R686 B.n90 B.n34 71.676
R687 B.n611 B.n33 71.676
R688 B.n540 B.n539 71.676
R689 B.n346 B.n300 71.676
R690 B.n532 B.n301 71.676
R691 B.n528 B.n302 71.676
R692 B.n524 B.n303 71.676
R693 B.n520 B.n304 71.676
R694 B.n516 B.n305 71.676
R695 B.n512 B.n306 71.676
R696 B.n508 B.n307 71.676
R697 B.n504 B.n308 71.676
R698 B.n500 B.n309 71.676
R699 B.n496 B.n310 71.676
R700 B.n492 B.n311 71.676
R701 B.n488 B.n312 71.676
R702 B.n484 B.n313 71.676
R703 B.n480 B.n314 71.676
R704 B.n476 B.n315 71.676
R705 B.n472 B.n316 71.676
R706 B.n468 B.n317 71.676
R707 B.n464 B.n318 71.676
R708 B.n460 B.n319 71.676
R709 B.n456 B.n320 71.676
R710 B.n452 B.n321 71.676
R711 B.n448 B.n322 71.676
R712 B.n444 B.n323 71.676
R713 B.n440 B.n324 71.676
R714 B.n435 B.n325 71.676
R715 B.n431 B.n326 71.676
R716 B.n427 B.n327 71.676
R717 B.n423 B.n328 71.676
R718 B.n419 B.n329 71.676
R719 B.n415 B.n330 71.676
R720 B.n411 B.n331 71.676
R721 B.n407 B.n332 71.676
R722 B.n403 B.n333 71.676
R723 B.n399 B.n334 71.676
R724 B.n395 B.n335 71.676
R725 B.n391 B.n336 71.676
R726 B.n387 B.n337 71.676
R727 B.n383 B.n338 71.676
R728 B.n379 B.n339 71.676
R729 B.n375 B.n340 71.676
R730 B.n371 B.n341 71.676
R731 B.n367 B.n342 71.676
R732 B.n363 B.n343 71.676
R733 B.n359 B.n344 71.676
R734 B.n355 B.n345 71.676
R735 B.n539 B.n299 71.676
R736 B.n533 B.n300 71.676
R737 B.n529 B.n301 71.676
R738 B.n525 B.n302 71.676
R739 B.n521 B.n303 71.676
R740 B.n517 B.n304 71.676
R741 B.n513 B.n305 71.676
R742 B.n509 B.n306 71.676
R743 B.n505 B.n307 71.676
R744 B.n501 B.n308 71.676
R745 B.n497 B.n309 71.676
R746 B.n493 B.n310 71.676
R747 B.n489 B.n311 71.676
R748 B.n485 B.n312 71.676
R749 B.n481 B.n313 71.676
R750 B.n477 B.n314 71.676
R751 B.n473 B.n315 71.676
R752 B.n469 B.n316 71.676
R753 B.n465 B.n317 71.676
R754 B.n461 B.n318 71.676
R755 B.n457 B.n319 71.676
R756 B.n453 B.n320 71.676
R757 B.n449 B.n321 71.676
R758 B.n445 B.n322 71.676
R759 B.n441 B.n323 71.676
R760 B.n436 B.n324 71.676
R761 B.n432 B.n325 71.676
R762 B.n428 B.n326 71.676
R763 B.n424 B.n327 71.676
R764 B.n420 B.n328 71.676
R765 B.n416 B.n329 71.676
R766 B.n412 B.n330 71.676
R767 B.n408 B.n331 71.676
R768 B.n404 B.n332 71.676
R769 B.n400 B.n333 71.676
R770 B.n396 B.n334 71.676
R771 B.n392 B.n335 71.676
R772 B.n388 B.n336 71.676
R773 B.n384 B.n337 71.676
R774 B.n380 B.n338 71.676
R775 B.n376 B.n339 71.676
R776 B.n372 B.n340 71.676
R777 B.n368 B.n341 71.676
R778 B.n364 B.n342 71.676
R779 B.n360 B.n343 71.676
R780 B.n356 B.n344 71.676
R781 B.n352 B.n345 71.676
R782 B.n646 B.n645 71.676
R783 B.n646 B.n2 71.676
R784 B.n83 B.t15 71.6108
R785 B.n351 B.t4 71.6108
R786 B.n86 B.t9 71.5951
R787 B.n348 B.t11 71.5951
R788 B.n538 B.n296 70.0879
R789 B.n610 B.n30 70.0879
R790 B.n169 B.n86 59.5399
R791 B.n84 B.n83 59.5399
R792 B.n438 B.n351 59.5399
R793 B.n349 B.n348 59.5399
R794 B.n545 B.n296 42.177
R795 B.n545 B.n292 42.177
R796 B.n551 B.n292 42.177
R797 B.n551 B.n288 42.177
R798 B.n557 B.n288 42.177
R799 B.n563 B.n284 42.177
R800 B.n563 B.n280 42.177
R801 B.n569 B.n280 42.177
R802 B.n569 B.n276 42.177
R803 B.n577 B.n276 42.177
R804 B.n577 B.n576 42.177
R805 B.n583 B.n4 42.177
R806 B.n644 B.n4 42.177
R807 B.n644 B.n643 42.177
R808 B.n643 B.n642 42.177
R809 B.n642 B.n8 42.177
R810 B.n635 B.n12 42.177
R811 B.n635 B.n634 42.177
R812 B.n634 B.n633 42.177
R813 B.n633 B.n16 42.177
R814 B.n627 B.n16 42.177
R815 B.n627 B.n626 42.177
R816 B.n625 B.n23 42.177
R817 B.n619 B.n23 42.177
R818 B.n619 B.n618 42.177
R819 B.n618 B.n617 42.177
R820 B.n617 B.n30 42.177
R821 B.n583 B.t1 38.4555
R822 B.t0 B.n8 38.4555
R823 B.n542 B.n541 33.5615
R824 B.n353 B.n294 33.5615
R825 B.n608 B.n607 33.5615
R826 B.n614 B.n613 33.5615
R827 B.t3 B.n284 31.0126
R828 B.n626 B.t7 31.0126
R829 B.n86 B.n85 23.855
R830 B.n83 B.n82 23.855
R831 B.n351 B.n350 23.855
R832 B.n348 B.n347 23.855
R833 B B.n647 18.0485
R834 B.n557 B.t3 11.1649
R835 B.t7 B.n625 11.1649
R836 B.n543 B.n542 10.6151
R837 B.n543 B.n290 10.6151
R838 B.n553 B.n290 10.6151
R839 B.n554 B.n553 10.6151
R840 B.n555 B.n554 10.6151
R841 B.n555 B.n282 10.6151
R842 B.n565 B.n282 10.6151
R843 B.n566 B.n565 10.6151
R844 B.n567 B.n566 10.6151
R845 B.n567 B.n274 10.6151
R846 B.n579 B.n274 10.6151
R847 B.n580 B.n579 10.6151
R848 B.n581 B.n580 10.6151
R849 B.n581 B.n0 10.6151
R850 B.n541 B.n298 10.6151
R851 B.n536 B.n298 10.6151
R852 B.n536 B.n535 10.6151
R853 B.n535 B.n534 10.6151
R854 B.n534 B.n531 10.6151
R855 B.n531 B.n530 10.6151
R856 B.n530 B.n527 10.6151
R857 B.n527 B.n526 10.6151
R858 B.n526 B.n523 10.6151
R859 B.n523 B.n522 10.6151
R860 B.n522 B.n519 10.6151
R861 B.n519 B.n518 10.6151
R862 B.n518 B.n515 10.6151
R863 B.n515 B.n514 10.6151
R864 B.n514 B.n511 10.6151
R865 B.n511 B.n510 10.6151
R866 B.n510 B.n507 10.6151
R867 B.n507 B.n506 10.6151
R868 B.n506 B.n503 10.6151
R869 B.n503 B.n502 10.6151
R870 B.n502 B.n499 10.6151
R871 B.n499 B.n498 10.6151
R872 B.n498 B.n495 10.6151
R873 B.n495 B.n494 10.6151
R874 B.n494 B.n491 10.6151
R875 B.n491 B.n490 10.6151
R876 B.n490 B.n487 10.6151
R877 B.n487 B.n486 10.6151
R878 B.n486 B.n483 10.6151
R879 B.n483 B.n482 10.6151
R880 B.n482 B.n479 10.6151
R881 B.n479 B.n478 10.6151
R882 B.n478 B.n475 10.6151
R883 B.n475 B.n474 10.6151
R884 B.n474 B.n471 10.6151
R885 B.n471 B.n470 10.6151
R886 B.n470 B.n467 10.6151
R887 B.n467 B.n466 10.6151
R888 B.n466 B.n463 10.6151
R889 B.n463 B.n462 10.6151
R890 B.n462 B.n459 10.6151
R891 B.n459 B.n458 10.6151
R892 B.n455 B.n454 10.6151
R893 B.n454 B.n451 10.6151
R894 B.n451 B.n450 10.6151
R895 B.n450 B.n447 10.6151
R896 B.n447 B.n446 10.6151
R897 B.n446 B.n443 10.6151
R898 B.n443 B.n442 10.6151
R899 B.n442 B.n439 10.6151
R900 B.n437 B.n434 10.6151
R901 B.n434 B.n433 10.6151
R902 B.n433 B.n430 10.6151
R903 B.n430 B.n429 10.6151
R904 B.n429 B.n426 10.6151
R905 B.n426 B.n425 10.6151
R906 B.n425 B.n422 10.6151
R907 B.n422 B.n421 10.6151
R908 B.n421 B.n418 10.6151
R909 B.n418 B.n417 10.6151
R910 B.n417 B.n414 10.6151
R911 B.n414 B.n413 10.6151
R912 B.n413 B.n410 10.6151
R913 B.n410 B.n409 10.6151
R914 B.n409 B.n406 10.6151
R915 B.n406 B.n405 10.6151
R916 B.n405 B.n402 10.6151
R917 B.n402 B.n401 10.6151
R918 B.n401 B.n398 10.6151
R919 B.n398 B.n397 10.6151
R920 B.n397 B.n394 10.6151
R921 B.n394 B.n393 10.6151
R922 B.n393 B.n390 10.6151
R923 B.n390 B.n389 10.6151
R924 B.n389 B.n386 10.6151
R925 B.n386 B.n385 10.6151
R926 B.n385 B.n382 10.6151
R927 B.n382 B.n381 10.6151
R928 B.n381 B.n378 10.6151
R929 B.n378 B.n377 10.6151
R930 B.n377 B.n374 10.6151
R931 B.n374 B.n373 10.6151
R932 B.n373 B.n370 10.6151
R933 B.n370 B.n369 10.6151
R934 B.n369 B.n366 10.6151
R935 B.n366 B.n365 10.6151
R936 B.n365 B.n362 10.6151
R937 B.n362 B.n361 10.6151
R938 B.n361 B.n358 10.6151
R939 B.n358 B.n357 10.6151
R940 B.n357 B.n354 10.6151
R941 B.n354 B.n353 10.6151
R942 B.n547 B.n294 10.6151
R943 B.n548 B.n547 10.6151
R944 B.n549 B.n548 10.6151
R945 B.n549 B.n286 10.6151
R946 B.n559 B.n286 10.6151
R947 B.n560 B.n559 10.6151
R948 B.n561 B.n560 10.6151
R949 B.n561 B.n278 10.6151
R950 B.n571 B.n278 10.6151
R951 B.n572 B.n571 10.6151
R952 B.n574 B.n572 10.6151
R953 B.n574 B.n573 10.6151
R954 B.n573 B.n271 10.6151
R955 B.n586 B.n271 10.6151
R956 B.n587 B.n586 10.6151
R957 B.n588 B.n587 10.6151
R958 B.n589 B.n588 10.6151
R959 B.n590 B.n589 10.6151
R960 B.n593 B.n590 10.6151
R961 B.n594 B.n593 10.6151
R962 B.n595 B.n594 10.6151
R963 B.n596 B.n595 10.6151
R964 B.n598 B.n596 10.6151
R965 B.n599 B.n598 10.6151
R966 B.n600 B.n599 10.6151
R967 B.n601 B.n600 10.6151
R968 B.n603 B.n601 10.6151
R969 B.n604 B.n603 10.6151
R970 B.n605 B.n604 10.6151
R971 B.n606 B.n605 10.6151
R972 B.n607 B.n606 10.6151
R973 B.n639 B.n1 10.6151
R974 B.n639 B.n638 10.6151
R975 B.n638 B.n637 10.6151
R976 B.n637 B.n10 10.6151
R977 B.n631 B.n10 10.6151
R978 B.n631 B.n630 10.6151
R979 B.n630 B.n629 10.6151
R980 B.n629 B.n18 10.6151
R981 B.n623 B.n18 10.6151
R982 B.n623 B.n622 10.6151
R983 B.n622 B.n621 10.6151
R984 B.n621 B.n25 10.6151
R985 B.n615 B.n25 10.6151
R986 B.n615 B.n614 10.6151
R987 B.n613 B.n32 10.6151
R988 B.n88 B.n32 10.6151
R989 B.n89 B.n88 10.6151
R990 B.n92 B.n89 10.6151
R991 B.n93 B.n92 10.6151
R992 B.n96 B.n93 10.6151
R993 B.n97 B.n96 10.6151
R994 B.n100 B.n97 10.6151
R995 B.n101 B.n100 10.6151
R996 B.n104 B.n101 10.6151
R997 B.n105 B.n104 10.6151
R998 B.n108 B.n105 10.6151
R999 B.n109 B.n108 10.6151
R1000 B.n112 B.n109 10.6151
R1001 B.n113 B.n112 10.6151
R1002 B.n116 B.n113 10.6151
R1003 B.n117 B.n116 10.6151
R1004 B.n120 B.n117 10.6151
R1005 B.n121 B.n120 10.6151
R1006 B.n124 B.n121 10.6151
R1007 B.n125 B.n124 10.6151
R1008 B.n128 B.n125 10.6151
R1009 B.n129 B.n128 10.6151
R1010 B.n132 B.n129 10.6151
R1011 B.n133 B.n132 10.6151
R1012 B.n136 B.n133 10.6151
R1013 B.n137 B.n136 10.6151
R1014 B.n140 B.n137 10.6151
R1015 B.n141 B.n140 10.6151
R1016 B.n144 B.n141 10.6151
R1017 B.n145 B.n144 10.6151
R1018 B.n148 B.n145 10.6151
R1019 B.n149 B.n148 10.6151
R1020 B.n152 B.n149 10.6151
R1021 B.n153 B.n152 10.6151
R1022 B.n156 B.n153 10.6151
R1023 B.n157 B.n156 10.6151
R1024 B.n160 B.n157 10.6151
R1025 B.n161 B.n160 10.6151
R1026 B.n164 B.n161 10.6151
R1027 B.n165 B.n164 10.6151
R1028 B.n168 B.n165 10.6151
R1029 B.n173 B.n170 10.6151
R1030 B.n174 B.n173 10.6151
R1031 B.n177 B.n174 10.6151
R1032 B.n178 B.n177 10.6151
R1033 B.n181 B.n178 10.6151
R1034 B.n182 B.n181 10.6151
R1035 B.n185 B.n182 10.6151
R1036 B.n186 B.n185 10.6151
R1037 B.n190 B.n189 10.6151
R1038 B.n193 B.n190 10.6151
R1039 B.n194 B.n193 10.6151
R1040 B.n197 B.n194 10.6151
R1041 B.n198 B.n197 10.6151
R1042 B.n201 B.n198 10.6151
R1043 B.n202 B.n201 10.6151
R1044 B.n205 B.n202 10.6151
R1045 B.n206 B.n205 10.6151
R1046 B.n209 B.n206 10.6151
R1047 B.n210 B.n209 10.6151
R1048 B.n213 B.n210 10.6151
R1049 B.n214 B.n213 10.6151
R1050 B.n217 B.n214 10.6151
R1051 B.n218 B.n217 10.6151
R1052 B.n221 B.n218 10.6151
R1053 B.n222 B.n221 10.6151
R1054 B.n225 B.n222 10.6151
R1055 B.n226 B.n225 10.6151
R1056 B.n229 B.n226 10.6151
R1057 B.n230 B.n229 10.6151
R1058 B.n233 B.n230 10.6151
R1059 B.n234 B.n233 10.6151
R1060 B.n237 B.n234 10.6151
R1061 B.n238 B.n237 10.6151
R1062 B.n241 B.n238 10.6151
R1063 B.n242 B.n241 10.6151
R1064 B.n245 B.n242 10.6151
R1065 B.n246 B.n245 10.6151
R1066 B.n249 B.n246 10.6151
R1067 B.n250 B.n249 10.6151
R1068 B.n253 B.n250 10.6151
R1069 B.n254 B.n253 10.6151
R1070 B.n257 B.n254 10.6151
R1071 B.n258 B.n257 10.6151
R1072 B.n261 B.n258 10.6151
R1073 B.n262 B.n261 10.6151
R1074 B.n265 B.n262 10.6151
R1075 B.n266 B.n265 10.6151
R1076 B.n269 B.n266 10.6151
R1077 B.n270 B.n269 10.6151
R1078 B.n608 B.n270 10.6151
R1079 B.n647 B.n0 8.11757
R1080 B.n647 B.n1 8.11757
R1081 B.n455 B.n349 7.18099
R1082 B.n439 B.n438 7.18099
R1083 B.n170 B.n169 7.18099
R1084 B.n186 B.n84 7.18099
R1085 B.n576 B.t1 3.72195
R1086 B.n12 B.t0 3.72195
R1087 B.n458 B.n349 3.43465
R1088 B.n438 B.n437 3.43465
R1089 B.n169 B.n168 3.43465
R1090 B.n189 B.n84 3.43465
R1091 VP.n0 VP.t1 578.561
R1092 VP.n0 VP.t0 538.063
R1093 VP VP.n0 0.0516364
R1094 VDD1 VDD1.t1 99.9147
R1095 VDD1 VDD1.t0 62.9265
C0 VTAIL VP 1.75276f
C1 VN VP 4.73141f
C2 VP VDD1 2.34377f
C3 VDD2 VTAIL 5.5781f
C4 VDD2 VN 2.23326f
C5 VDD2 VDD1 0.481971f
C6 VN VTAIL 1.73819f
C7 VTAIL VDD1 5.5424f
C8 VN VDD1 0.149013f
C9 VDD2 VP 0.263705f
C10 VDD2 B 3.90802f
C11 VDD1 B 6.72601f
C12 VTAIL B 6.642742f
C13 VN B 8.232241f
C14 VP B 4.300385f
C15 VDD1.t0 B 2.27789f
C16 VDD1.t1 B 2.78463f
C17 VP.t1 B 1.62716f
C18 VP.t0 B 1.48762f
C19 VP.n0 B 3.86553f
C20 VDD2.t0 B 2.7853f
C21 VDD2.t1 B 2.29874f
C22 VDD2.n0 B 2.65889f
C23 VTAIL.t1 B 1.68235f
C24 VTAIL.n0 B 1.10888f
C25 VTAIL.t3 B 1.68236f
C26 VTAIL.n1 B 1.11926f
C27 VTAIL.t0 B 1.68235f
C28 VTAIL.n2 B 1.06603f
C29 VTAIL.t2 B 1.68235f
C30 VTAIL.n3 B 1.02621f
C31 VN.t1 B 1.45421f
C32 VN.t0 B 1.59367f
.ends

