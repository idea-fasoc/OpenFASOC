* NGSPICE file created from diff_pair_sample_0050.ext - technology: sky130A

.subckt diff_pair_sample_0050 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=6.1308 pd=32.22 as=2.5938 ps=16.05 w=15.72 l=2.1
X1 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=6.1308 pd=32.22 as=0 ps=0 w=15.72 l=2.1
X2 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=6.1308 pd=32.22 as=0 ps=0 w=15.72 l=2.1
X3 VTAIL.t1 VN.t0 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=6.1308 pd=32.22 as=2.5938 ps=16.05 w=15.72 l=2.1
X4 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.1308 pd=32.22 as=0 ps=0 w=15.72 l=2.1
X5 VDD2.t2 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.5938 pd=16.05 as=6.1308 ps=32.22 w=15.72 l=2.1
X6 VDD2.t1 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.5938 pd=16.05 as=6.1308 ps=32.22 w=15.72 l=2.1
X7 VTAIL.t0 VN.t3 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.1308 pd=32.22 as=2.5938 ps=16.05 w=15.72 l=2.1
X8 VTAIL.t6 VP.t1 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=6.1308 pd=32.22 as=2.5938 ps=16.05 w=15.72 l=2.1
X9 VDD1.t1 VP.t2 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.5938 pd=16.05 as=6.1308 ps=32.22 w=15.72 l=2.1
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.1308 pd=32.22 as=0 ps=0 w=15.72 l=2.1
X11 VDD1.t2 VP.t3 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.5938 pd=16.05 as=6.1308 ps=32.22 w=15.72 l=2.1
R0 VP.n2 VP.t1 216.589
R1 VP.n2 VP.t2 216.041
R2 VP.n4 VP.t0 180.406
R3 VP.n11 VP.t3 180.406
R4 VP.n10 VP.n0 161.3
R5 VP.n9 VP.n8 161.3
R6 VP.n7 VP.n1 161.3
R7 VP.n6 VP.n5 161.3
R8 VP.n4 VP.n3 88.0378
R9 VP.n12 VP.n11 88.0378
R10 VP.n9 VP.n1 56.5617
R11 VP.n3 VP.n2 54.5209
R12 VP.n5 VP.n1 24.5923
R13 VP.n10 VP.n9 24.5923
R14 VP.n5 VP.n4 22.8709
R15 VP.n11 VP.n10 22.8709
R16 VP.n6 VP.n3 0.278335
R17 VP.n12 VP.n0 0.278335
R18 VP.n7 VP.n6 0.189894
R19 VP.n8 VP.n7 0.189894
R20 VP.n8 VP.n0 0.189894
R21 VP VP.n12 0.153485
R22 VDD1 VDD1.n1 104.883
R23 VDD1 VDD1.n0 60.8663
R24 VDD1.n0 VDD1.t0 1.26004
R25 VDD1.n0 VDD1.t1 1.26004
R26 VDD1.n1 VDD1.t3 1.26004
R27 VDD1.n1 VDD1.t2 1.26004
R28 VTAIL.n5 VTAIL.t6 45.389
R29 VTAIL.n4 VTAIL.t3 45.389
R30 VTAIL.n3 VTAIL.t0 45.389
R31 VTAIL.n7 VTAIL.t2 45.3889
R32 VTAIL.n0 VTAIL.t1 45.3889
R33 VTAIL.n1 VTAIL.t4 45.3889
R34 VTAIL.n2 VTAIL.t7 45.3889
R35 VTAIL.n6 VTAIL.t5 45.3889
R36 VTAIL.n7 VTAIL.n6 28.0134
R37 VTAIL.n3 VTAIL.n2 28.0134
R38 VTAIL.n4 VTAIL.n3 2.09533
R39 VTAIL.n6 VTAIL.n5 2.09533
R40 VTAIL.n2 VTAIL.n1 2.09533
R41 VTAIL VTAIL.n0 1.1061
R42 VTAIL VTAIL.n7 0.989724
R43 VTAIL.n5 VTAIL.n4 0.470328
R44 VTAIL.n1 VTAIL.n0 0.470328
R45 B.n824 B.n823 585
R46 B.n825 B.n824 585
R47 B.n347 B.n114 585
R48 B.n346 B.n345 585
R49 B.n344 B.n343 585
R50 B.n342 B.n341 585
R51 B.n340 B.n339 585
R52 B.n338 B.n337 585
R53 B.n336 B.n335 585
R54 B.n334 B.n333 585
R55 B.n332 B.n331 585
R56 B.n330 B.n329 585
R57 B.n328 B.n327 585
R58 B.n326 B.n325 585
R59 B.n324 B.n323 585
R60 B.n322 B.n321 585
R61 B.n320 B.n319 585
R62 B.n318 B.n317 585
R63 B.n316 B.n315 585
R64 B.n314 B.n313 585
R65 B.n312 B.n311 585
R66 B.n310 B.n309 585
R67 B.n308 B.n307 585
R68 B.n306 B.n305 585
R69 B.n304 B.n303 585
R70 B.n302 B.n301 585
R71 B.n300 B.n299 585
R72 B.n298 B.n297 585
R73 B.n296 B.n295 585
R74 B.n294 B.n293 585
R75 B.n292 B.n291 585
R76 B.n290 B.n289 585
R77 B.n288 B.n287 585
R78 B.n286 B.n285 585
R79 B.n284 B.n283 585
R80 B.n282 B.n281 585
R81 B.n280 B.n279 585
R82 B.n278 B.n277 585
R83 B.n276 B.n275 585
R84 B.n274 B.n273 585
R85 B.n272 B.n271 585
R86 B.n270 B.n269 585
R87 B.n268 B.n267 585
R88 B.n266 B.n265 585
R89 B.n264 B.n263 585
R90 B.n262 B.n261 585
R91 B.n260 B.n259 585
R92 B.n258 B.n257 585
R93 B.n256 B.n255 585
R94 B.n254 B.n253 585
R95 B.n252 B.n251 585
R96 B.n250 B.n249 585
R97 B.n248 B.n247 585
R98 B.n246 B.n245 585
R99 B.n244 B.n243 585
R100 B.n242 B.n241 585
R101 B.n240 B.n239 585
R102 B.n238 B.n237 585
R103 B.n236 B.n235 585
R104 B.n234 B.n233 585
R105 B.n232 B.n231 585
R106 B.n230 B.n229 585
R107 B.n228 B.n227 585
R108 B.n225 B.n224 585
R109 B.n223 B.n222 585
R110 B.n221 B.n220 585
R111 B.n219 B.n218 585
R112 B.n217 B.n216 585
R113 B.n215 B.n214 585
R114 B.n213 B.n212 585
R115 B.n211 B.n210 585
R116 B.n209 B.n208 585
R117 B.n207 B.n206 585
R118 B.n205 B.n204 585
R119 B.n203 B.n202 585
R120 B.n201 B.n200 585
R121 B.n199 B.n198 585
R122 B.n197 B.n196 585
R123 B.n195 B.n194 585
R124 B.n193 B.n192 585
R125 B.n191 B.n190 585
R126 B.n189 B.n188 585
R127 B.n187 B.n186 585
R128 B.n185 B.n184 585
R129 B.n183 B.n182 585
R130 B.n181 B.n180 585
R131 B.n179 B.n178 585
R132 B.n177 B.n176 585
R133 B.n175 B.n174 585
R134 B.n173 B.n172 585
R135 B.n171 B.n170 585
R136 B.n169 B.n168 585
R137 B.n167 B.n166 585
R138 B.n165 B.n164 585
R139 B.n163 B.n162 585
R140 B.n161 B.n160 585
R141 B.n159 B.n158 585
R142 B.n157 B.n156 585
R143 B.n155 B.n154 585
R144 B.n153 B.n152 585
R145 B.n151 B.n150 585
R146 B.n149 B.n148 585
R147 B.n147 B.n146 585
R148 B.n145 B.n144 585
R149 B.n143 B.n142 585
R150 B.n141 B.n140 585
R151 B.n139 B.n138 585
R152 B.n137 B.n136 585
R153 B.n135 B.n134 585
R154 B.n133 B.n132 585
R155 B.n131 B.n130 585
R156 B.n129 B.n128 585
R157 B.n127 B.n126 585
R158 B.n125 B.n124 585
R159 B.n123 B.n122 585
R160 B.n121 B.n120 585
R161 B.n822 B.n56 585
R162 B.n826 B.n56 585
R163 B.n821 B.n55 585
R164 B.n827 B.n55 585
R165 B.n820 B.n819 585
R166 B.n819 B.n51 585
R167 B.n818 B.n50 585
R168 B.n833 B.n50 585
R169 B.n817 B.n49 585
R170 B.n834 B.n49 585
R171 B.n816 B.n48 585
R172 B.n835 B.n48 585
R173 B.n815 B.n814 585
R174 B.n814 B.n47 585
R175 B.n813 B.n43 585
R176 B.n841 B.n43 585
R177 B.n812 B.n42 585
R178 B.n842 B.n42 585
R179 B.n811 B.n41 585
R180 B.n843 B.n41 585
R181 B.n810 B.n809 585
R182 B.n809 B.n37 585
R183 B.n808 B.n36 585
R184 B.n849 B.n36 585
R185 B.n807 B.n35 585
R186 B.n850 B.n35 585
R187 B.n806 B.n34 585
R188 B.n851 B.n34 585
R189 B.n805 B.n804 585
R190 B.n804 B.n30 585
R191 B.n803 B.n29 585
R192 B.n857 B.n29 585
R193 B.n802 B.n28 585
R194 B.n858 B.n28 585
R195 B.n801 B.n27 585
R196 B.n859 B.n27 585
R197 B.n800 B.n799 585
R198 B.n799 B.n23 585
R199 B.n798 B.n22 585
R200 B.n865 B.n22 585
R201 B.n797 B.n21 585
R202 B.n866 B.n21 585
R203 B.n796 B.n20 585
R204 B.n867 B.n20 585
R205 B.n795 B.n794 585
R206 B.n794 B.n16 585
R207 B.n793 B.n15 585
R208 B.n873 B.n15 585
R209 B.n792 B.n14 585
R210 B.n874 B.n14 585
R211 B.n791 B.n13 585
R212 B.n875 B.n13 585
R213 B.n790 B.n789 585
R214 B.n789 B.n12 585
R215 B.n788 B.n787 585
R216 B.n788 B.n8 585
R217 B.n786 B.n7 585
R218 B.n882 B.n7 585
R219 B.n785 B.n6 585
R220 B.n883 B.n6 585
R221 B.n784 B.n5 585
R222 B.n884 B.n5 585
R223 B.n783 B.n782 585
R224 B.n782 B.n4 585
R225 B.n781 B.n348 585
R226 B.n781 B.n780 585
R227 B.n771 B.n349 585
R228 B.n350 B.n349 585
R229 B.n773 B.n772 585
R230 B.n774 B.n773 585
R231 B.n770 B.n354 585
R232 B.n358 B.n354 585
R233 B.n769 B.n768 585
R234 B.n768 B.n767 585
R235 B.n356 B.n355 585
R236 B.n357 B.n356 585
R237 B.n760 B.n759 585
R238 B.n761 B.n760 585
R239 B.n758 B.n363 585
R240 B.n363 B.n362 585
R241 B.n757 B.n756 585
R242 B.n756 B.n755 585
R243 B.n365 B.n364 585
R244 B.n366 B.n365 585
R245 B.n748 B.n747 585
R246 B.n749 B.n748 585
R247 B.n746 B.n371 585
R248 B.n371 B.n370 585
R249 B.n745 B.n744 585
R250 B.n744 B.n743 585
R251 B.n373 B.n372 585
R252 B.n374 B.n373 585
R253 B.n736 B.n735 585
R254 B.n737 B.n736 585
R255 B.n734 B.n379 585
R256 B.n379 B.n378 585
R257 B.n733 B.n732 585
R258 B.n732 B.n731 585
R259 B.n381 B.n380 585
R260 B.n382 B.n381 585
R261 B.n724 B.n723 585
R262 B.n725 B.n724 585
R263 B.n722 B.n387 585
R264 B.n387 B.n386 585
R265 B.n721 B.n720 585
R266 B.n720 B.n719 585
R267 B.n389 B.n388 585
R268 B.n712 B.n389 585
R269 B.n711 B.n710 585
R270 B.n713 B.n711 585
R271 B.n709 B.n394 585
R272 B.n394 B.n393 585
R273 B.n708 B.n707 585
R274 B.n707 B.n706 585
R275 B.n396 B.n395 585
R276 B.n397 B.n396 585
R277 B.n699 B.n698 585
R278 B.n700 B.n699 585
R279 B.n697 B.n402 585
R280 B.n402 B.n401 585
R281 B.n691 B.n690 585
R282 B.n689 B.n461 585
R283 B.n688 B.n460 585
R284 B.n693 B.n460 585
R285 B.n687 B.n686 585
R286 B.n685 B.n684 585
R287 B.n683 B.n682 585
R288 B.n681 B.n680 585
R289 B.n679 B.n678 585
R290 B.n677 B.n676 585
R291 B.n675 B.n674 585
R292 B.n673 B.n672 585
R293 B.n671 B.n670 585
R294 B.n669 B.n668 585
R295 B.n667 B.n666 585
R296 B.n665 B.n664 585
R297 B.n663 B.n662 585
R298 B.n661 B.n660 585
R299 B.n659 B.n658 585
R300 B.n657 B.n656 585
R301 B.n655 B.n654 585
R302 B.n653 B.n652 585
R303 B.n651 B.n650 585
R304 B.n649 B.n648 585
R305 B.n647 B.n646 585
R306 B.n645 B.n644 585
R307 B.n643 B.n642 585
R308 B.n641 B.n640 585
R309 B.n639 B.n638 585
R310 B.n637 B.n636 585
R311 B.n635 B.n634 585
R312 B.n633 B.n632 585
R313 B.n631 B.n630 585
R314 B.n629 B.n628 585
R315 B.n627 B.n626 585
R316 B.n625 B.n624 585
R317 B.n623 B.n622 585
R318 B.n621 B.n620 585
R319 B.n619 B.n618 585
R320 B.n617 B.n616 585
R321 B.n615 B.n614 585
R322 B.n613 B.n612 585
R323 B.n611 B.n610 585
R324 B.n609 B.n608 585
R325 B.n607 B.n606 585
R326 B.n605 B.n604 585
R327 B.n603 B.n602 585
R328 B.n601 B.n600 585
R329 B.n599 B.n598 585
R330 B.n597 B.n596 585
R331 B.n595 B.n594 585
R332 B.n593 B.n592 585
R333 B.n591 B.n590 585
R334 B.n589 B.n588 585
R335 B.n587 B.n586 585
R336 B.n585 B.n584 585
R337 B.n583 B.n582 585
R338 B.n581 B.n580 585
R339 B.n579 B.n578 585
R340 B.n577 B.n576 585
R341 B.n575 B.n574 585
R342 B.n573 B.n572 585
R343 B.n571 B.n570 585
R344 B.n568 B.n567 585
R345 B.n566 B.n565 585
R346 B.n564 B.n563 585
R347 B.n562 B.n561 585
R348 B.n560 B.n559 585
R349 B.n558 B.n557 585
R350 B.n556 B.n555 585
R351 B.n554 B.n553 585
R352 B.n552 B.n551 585
R353 B.n550 B.n549 585
R354 B.n548 B.n547 585
R355 B.n546 B.n545 585
R356 B.n544 B.n543 585
R357 B.n542 B.n541 585
R358 B.n540 B.n539 585
R359 B.n538 B.n537 585
R360 B.n536 B.n535 585
R361 B.n534 B.n533 585
R362 B.n532 B.n531 585
R363 B.n530 B.n529 585
R364 B.n528 B.n527 585
R365 B.n526 B.n525 585
R366 B.n524 B.n523 585
R367 B.n522 B.n521 585
R368 B.n520 B.n519 585
R369 B.n518 B.n517 585
R370 B.n516 B.n515 585
R371 B.n514 B.n513 585
R372 B.n512 B.n511 585
R373 B.n510 B.n509 585
R374 B.n508 B.n507 585
R375 B.n506 B.n505 585
R376 B.n504 B.n503 585
R377 B.n502 B.n501 585
R378 B.n500 B.n499 585
R379 B.n498 B.n497 585
R380 B.n496 B.n495 585
R381 B.n494 B.n493 585
R382 B.n492 B.n491 585
R383 B.n490 B.n489 585
R384 B.n488 B.n487 585
R385 B.n486 B.n485 585
R386 B.n484 B.n483 585
R387 B.n482 B.n481 585
R388 B.n480 B.n479 585
R389 B.n478 B.n477 585
R390 B.n476 B.n475 585
R391 B.n474 B.n473 585
R392 B.n472 B.n471 585
R393 B.n470 B.n469 585
R394 B.n468 B.n467 585
R395 B.n404 B.n403 585
R396 B.n696 B.n695 585
R397 B.n400 B.n399 585
R398 B.n401 B.n400 585
R399 B.n702 B.n701 585
R400 B.n701 B.n700 585
R401 B.n703 B.n398 585
R402 B.n398 B.n397 585
R403 B.n705 B.n704 585
R404 B.n706 B.n705 585
R405 B.n392 B.n391 585
R406 B.n393 B.n392 585
R407 B.n715 B.n714 585
R408 B.n714 B.n713 585
R409 B.n716 B.n390 585
R410 B.n712 B.n390 585
R411 B.n718 B.n717 585
R412 B.n719 B.n718 585
R413 B.n385 B.n384 585
R414 B.n386 B.n385 585
R415 B.n727 B.n726 585
R416 B.n726 B.n725 585
R417 B.n728 B.n383 585
R418 B.n383 B.n382 585
R419 B.n730 B.n729 585
R420 B.n731 B.n730 585
R421 B.n377 B.n376 585
R422 B.n378 B.n377 585
R423 B.n739 B.n738 585
R424 B.n738 B.n737 585
R425 B.n740 B.n375 585
R426 B.n375 B.n374 585
R427 B.n742 B.n741 585
R428 B.n743 B.n742 585
R429 B.n369 B.n368 585
R430 B.n370 B.n369 585
R431 B.n751 B.n750 585
R432 B.n750 B.n749 585
R433 B.n752 B.n367 585
R434 B.n367 B.n366 585
R435 B.n754 B.n753 585
R436 B.n755 B.n754 585
R437 B.n361 B.n360 585
R438 B.n362 B.n361 585
R439 B.n763 B.n762 585
R440 B.n762 B.n761 585
R441 B.n764 B.n359 585
R442 B.n359 B.n357 585
R443 B.n766 B.n765 585
R444 B.n767 B.n766 585
R445 B.n353 B.n352 585
R446 B.n358 B.n353 585
R447 B.n776 B.n775 585
R448 B.n775 B.n774 585
R449 B.n777 B.n351 585
R450 B.n351 B.n350 585
R451 B.n779 B.n778 585
R452 B.n780 B.n779 585
R453 B.n3 B.n0 585
R454 B.n4 B.n3 585
R455 B.n881 B.n1 585
R456 B.n882 B.n881 585
R457 B.n880 B.n879 585
R458 B.n880 B.n8 585
R459 B.n878 B.n9 585
R460 B.n12 B.n9 585
R461 B.n877 B.n876 585
R462 B.n876 B.n875 585
R463 B.n11 B.n10 585
R464 B.n874 B.n11 585
R465 B.n872 B.n871 585
R466 B.n873 B.n872 585
R467 B.n870 B.n17 585
R468 B.n17 B.n16 585
R469 B.n869 B.n868 585
R470 B.n868 B.n867 585
R471 B.n19 B.n18 585
R472 B.n866 B.n19 585
R473 B.n864 B.n863 585
R474 B.n865 B.n864 585
R475 B.n862 B.n24 585
R476 B.n24 B.n23 585
R477 B.n861 B.n860 585
R478 B.n860 B.n859 585
R479 B.n26 B.n25 585
R480 B.n858 B.n26 585
R481 B.n856 B.n855 585
R482 B.n857 B.n856 585
R483 B.n854 B.n31 585
R484 B.n31 B.n30 585
R485 B.n853 B.n852 585
R486 B.n852 B.n851 585
R487 B.n33 B.n32 585
R488 B.n850 B.n33 585
R489 B.n848 B.n847 585
R490 B.n849 B.n848 585
R491 B.n846 B.n38 585
R492 B.n38 B.n37 585
R493 B.n845 B.n844 585
R494 B.n844 B.n843 585
R495 B.n40 B.n39 585
R496 B.n842 B.n40 585
R497 B.n840 B.n839 585
R498 B.n841 B.n840 585
R499 B.n838 B.n44 585
R500 B.n47 B.n44 585
R501 B.n837 B.n836 585
R502 B.n836 B.n835 585
R503 B.n46 B.n45 585
R504 B.n834 B.n46 585
R505 B.n832 B.n831 585
R506 B.n833 B.n832 585
R507 B.n830 B.n52 585
R508 B.n52 B.n51 585
R509 B.n829 B.n828 585
R510 B.n828 B.n827 585
R511 B.n54 B.n53 585
R512 B.n826 B.n54 585
R513 B.n885 B.n884 585
R514 B.n883 B.n2 585
R515 B.n120 B.n54 482.89
R516 B.n824 B.n56 482.89
R517 B.n695 B.n402 482.89
R518 B.n691 B.n400 482.89
R519 B.n118 B.t15 387.548
R520 B.n115 B.t8 387.548
R521 B.n465 B.t4 387.548
R522 B.n462 B.t12 387.548
R523 B.n825 B.n113 256.663
R524 B.n825 B.n112 256.663
R525 B.n825 B.n111 256.663
R526 B.n825 B.n110 256.663
R527 B.n825 B.n109 256.663
R528 B.n825 B.n108 256.663
R529 B.n825 B.n107 256.663
R530 B.n825 B.n106 256.663
R531 B.n825 B.n105 256.663
R532 B.n825 B.n104 256.663
R533 B.n825 B.n103 256.663
R534 B.n825 B.n102 256.663
R535 B.n825 B.n101 256.663
R536 B.n825 B.n100 256.663
R537 B.n825 B.n99 256.663
R538 B.n825 B.n98 256.663
R539 B.n825 B.n97 256.663
R540 B.n825 B.n96 256.663
R541 B.n825 B.n95 256.663
R542 B.n825 B.n94 256.663
R543 B.n825 B.n93 256.663
R544 B.n825 B.n92 256.663
R545 B.n825 B.n91 256.663
R546 B.n825 B.n90 256.663
R547 B.n825 B.n89 256.663
R548 B.n825 B.n88 256.663
R549 B.n825 B.n87 256.663
R550 B.n825 B.n86 256.663
R551 B.n825 B.n85 256.663
R552 B.n825 B.n84 256.663
R553 B.n825 B.n83 256.663
R554 B.n825 B.n82 256.663
R555 B.n825 B.n81 256.663
R556 B.n825 B.n80 256.663
R557 B.n825 B.n79 256.663
R558 B.n825 B.n78 256.663
R559 B.n825 B.n77 256.663
R560 B.n825 B.n76 256.663
R561 B.n825 B.n75 256.663
R562 B.n825 B.n74 256.663
R563 B.n825 B.n73 256.663
R564 B.n825 B.n72 256.663
R565 B.n825 B.n71 256.663
R566 B.n825 B.n70 256.663
R567 B.n825 B.n69 256.663
R568 B.n825 B.n68 256.663
R569 B.n825 B.n67 256.663
R570 B.n825 B.n66 256.663
R571 B.n825 B.n65 256.663
R572 B.n825 B.n64 256.663
R573 B.n825 B.n63 256.663
R574 B.n825 B.n62 256.663
R575 B.n825 B.n61 256.663
R576 B.n825 B.n60 256.663
R577 B.n825 B.n59 256.663
R578 B.n825 B.n58 256.663
R579 B.n825 B.n57 256.663
R580 B.n693 B.n692 256.663
R581 B.n693 B.n405 256.663
R582 B.n693 B.n406 256.663
R583 B.n693 B.n407 256.663
R584 B.n693 B.n408 256.663
R585 B.n693 B.n409 256.663
R586 B.n693 B.n410 256.663
R587 B.n693 B.n411 256.663
R588 B.n693 B.n412 256.663
R589 B.n693 B.n413 256.663
R590 B.n693 B.n414 256.663
R591 B.n693 B.n415 256.663
R592 B.n693 B.n416 256.663
R593 B.n693 B.n417 256.663
R594 B.n693 B.n418 256.663
R595 B.n693 B.n419 256.663
R596 B.n693 B.n420 256.663
R597 B.n693 B.n421 256.663
R598 B.n693 B.n422 256.663
R599 B.n693 B.n423 256.663
R600 B.n693 B.n424 256.663
R601 B.n693 B.n425 256.663
R602 B.n693 B.n426 256.663
R603 B.n693 B.n427 256.663
R604 B.n693 B.n428 256.663
R605 B.n693 B.n429 256.663
R606 B.n693 B.n430 256.663
R607 B.n693 B.n431 256.663
R608 B.n693 B.n432 256.663
R609 B.n693 B.n433 256.663
R610 B.n693 B.n434 256.663
R611 B.n693 B.n435 256.663
R612 B.n693 B.n436 256.663
R613 B.n693 B.n437 256.663
R614 B.n693 B.n438 256.663
R615 B.n693 B.n439 256.663
R616 B.n693 B.n440 256.663
R617 B.n693 B.n441 256.663
R618 B.n693 B.n442 256.663
R619 B.n693 B.n443 256.663
R620 B.n693 B.n444 256.663
R621 B.n693 B.n445 256.663
R622 B.n693 B.n446 256.663
R623 B.n693 B.n447 256.663
R624 B.n693 B.n448 256.663
R625 B.n693 B.n449 256.663
R626 B.n693 B.n450 256.663
R627 B.n693 B.n451 256.663
R628 B.n693 B.n452 256.663
R629 B.n693 B.n453 256.663
R630 B.n693 B.n454 256.663
R631 B.n693 B.n455 256.663
R632 B.n693 B.n456 256.663
R633 B.n693 B.n457 256.663
R634 B.n693 B.n458 256.663
R635 B.n693 B.n459 256.663
R636 B.n694 B.n693 256.663
R637 B.n887 B.n886 256.663
R638 B.n124 B.n123 163.367
R639 B.n128 B.n127 163.367
R640 B.n132 B.n131 163.367
R641 B.n136 B.n135 163.367
R642 B.n140 B.n139 163.367
R643 B.n144 B.n143 163.367
R644 B.n148 B.n147 163.367
R645 B.n152 B.n151 163.367
R646 B.n156 B.n155 163.367
R647 B.n160 B.n159 163.367
R648 B.n164 B.n163 163.367
R649 B.n168 B.n167 163.367
R650 B.n172 B.n171 163.367
R651 B.n176 B.n175 163.367
R652 B.n180 B.n179 163.367
R653 B.n184 B.n183 163.367
R654 B.n188 B.n187 163.367
R655 B.n192 B.n191 163.367
R656 B.n196 B.n195 163.367
R657 B.n200 B.n199 163.367
R658 B.n204 B.n203 163.367
R659 B.n208 B.n207 163.367
R660 B.n212 B.n211 163.367
R661 B.n216 B.n215 163.367
R662 B.n220 B.n219 163.367
R663 B.n224 B.n223 163.367
R664 B.n229 B.n228 163.367
R665 B.n233 B.n232 163.367
R666 B.n237 B.n236 163.367
R667 B.n241 B.n240 163.367
R668 B.n245 B.n244 163.367
R669 B.n249 B.n248 163.367
R670 B.n253 B.n252 163.367
R671 B.n257 B.n256 163.367
R672 B.n261 B.n260 163.367
R673 B.n265 B.n264 163.367
R674 B.n269 B.n268 163.367
R675 B.n273 B.n272 163.367
R676 B.n277 B.n276 163.367
R677 B.n281 B.n280 163.367
R678 B.n285 B.n284 163.367
R679 B.n289 B.n288 163.367
R680 B.n293 B.n292 163.367
R681 B.n297 B.n296 163.367
R682 B.n301 B.n300 163.367
R683 B.n305 B.n304 163.367
R684 B.n309 B.n308 163.367
R685 B.n313 B.n312 163.367
R686 B.n317 B.n316 163.367
R687 B.n321 B.n320 163.367
R688 B.n325 B.n324 163.367
R689 B.n329 B.n328 163.367
R690 B.n333 B.n332 163.367
R691 B.n337 B.n336 163.367
R692 B.n341 B.n340 163.367
R693 B.n345 B.n344 163.367
R694 B.n824 B.n114 163.367
R695 B.n699 B.n402 163.367
R696 B.n699 B.n396 163.367
R697 B.n707 B.n396 163.367
R698 B.n707 B.n394 163.367
R699 B.n711 B.n394 163.367
R700 B.n711 B.n389 163.367
R701 B.n720 B.n389 163.367
R702 B.n720 B.n387 163.367
R703 B.n724 B.n387 163.367
R704 B.n724 B.n381 163.367
R705 B.n732 B.n381 163.367
R706 B.n732 B.n379 163.367
R707 B.n736 B.n379 163.367
R708 B.n736 B.n373 163.367
R709 B.n744 B.n373 163.367
R710 B.n744 B.n371 163.367
R711 B.n748 B.n371 163.367
R712 B.n748 B.n365 163.367
R713 B.n756 B.n365 163.367
R714 B.n756 B.n363 163.367
R715 B.n760 B.n363 163.367
R716 B.n760 B.n356 163.367
R717 B.n768 B.n356 163.367
R718 B.n768 B.n354 163.367
R719 B.n773 B.n354 163.367
R720 B.n773 B.n349 163.367
R721 B.n781 B.n349 163.367
R722 B.n782 B.n781 163.367
R723 B.n782 B.n5 163.367
R724 B.n6 B.n5 163.367
R725 B.n7 B.n6 163.367
R726 B.n788 B.n7 163.367
R727 B.n789 B.n788 163.367
R728 B.n789 B.n13 163.367
R729 B.n14 B.n13 163.367
R730 B.n15 B.n14 163.367
R731 B.n794 B.n15 163.367
R732 B.n794 B.n20 163.367
R733 B.n21 B.n20 163.367
R734 B.n22 B.n21 163.367
R735 B.n799 B.n22 163.367
R736 B.n799 B.n27 163.367
R737 B.n28 B.n27 163.367
R738 B.n29 B.n28 163.367
R739 B.n804 B.n29 163.367
R740 B.n804 B.n34 163.367
R741 B.n35 B.n34 163.367
R742 B.n36 B.n35 163.367
R743 B.n809 B.n36 163.367
R744 B.n809 B.n41 163.367
R745 B.n42 B.n41 163.367
R746 B.n43 B.n42 163.367
R747 B.n814 B.n43 163.367
R748 B.n814 B.n48 163.367
R749 B.n49 B.n48 163.367
R750 B.n50 B.n49 163.367
R751 B.n819 B.n50 163.367
R752 B.n819 B.n55 163.367
R753 B.n56 B.n55 163.367
R754 B.n461 B.n460 163.367
R755 B.n686 B.n460 163.367
R756 B.n684 B.n683 163.367
R757 B.n680 B.n679 163.367
R758 B.n676 B.n675 163.367
R759 B.n672 B.n671 163.367
R760 B.n668 B.n667 163.367
R761 B.n664 B.n663 163.367
R762 B.n660 B.n659 163.367
R763 B.n656 B.n655 163.367
R764 B.n652 B.n651 163.367
R765 B.n648 B.n647 163.367
R766 B.n644 B.n643 163.367
R767 B.n640 B.n639 163.367
R768 B.n636 B.n635 163.367
R769 B.n632 B.n631 163.367
R770 B.n628 B.n627 163.367
R771 B.n624 B.n623 163.367
R772 B.n620 B.n619 163.367
R773 B.n616 B.n615 163.367
R774 B.n612 B.n611 163.367
R775 B.n608 B.n607 163.367
R776 B.n604 B.n603 163.367
R777 B.n600 B.n599 163.367
R778 B.n596 B.n595 163.367
R779 B.n592 B.n591 163.367
R780 B.n588 B.n587 163.367
R781 B.n584 B.n583 163.367
R782 B.n580 B.n579 163.367
R783 B.n576 B.n575 163.367
R784 B.n572 B.n571 163.367
R785 B.n567 B.n566 163.367
R786 B.n563 B.n562 163.367
R787 B.n559 B.n558 163.367
R788 B.n555 B.n554 163.367
R789 B.n551 B.n550 163.367
R790 B.n547 B.n546 163.367
R791 B.n543 B.n542 163.367
R792 B.n539 B.n538 163.367
R793 B.n535 B.n534 163.367
R794 B.n531 B.n530 163.367
R795 B.n527 B.n526 163.367
R796 B.n523 B.n522 163.367
R797 B.n519 B.n518 163.367
R798 B.n515 B.n514 163.367
R799 B.n511 B.n510 163.367
R800 B.n507 B.n506 163.367
R801 B.n503 B.n502 163.367
R802 B.n499 B.n498 163.367
R803 B.n495 B.n494 163.367
R804 B.n491 B.n490 163.367
R805 B.n487 B.n486 163.367
R806 B.n483 B.n482 163.367
R807 B.n479 B.n478 163.367
R808 B.n475 B.n474 163.367
R809 B.n471 B.n470 163.367
R810 B.n467 B.n404 163.367
R811 B.n701 B.n400 163.367
R812 B.n701 B.n398 163.367
R813 B.n705 B.n398 163.367
R814 B.n705 B.n392 163.367
R815 B.n714 B.n392 163.367
R816 B.n714 B.n390 163.367
R817 B.n718 B.n390 163.367
R818 B.n718 B.n385 163.367
R819 B.n726 B.n385 163.367
R820 B.n726 B.n383 163.367
R821 B.n730 B.n383 163.367
R822 B.n730 B.n377 163.367
R823 B.n738 B.n377 163.367
R824 B.n738 B.n375 163.367
R825 B.n742 B.n375 163.367
R826 B.n742 B.n369 163.367
R827 B.n750 B.n369 163.367
R828 B.n750 B.n367 163.367
R829 B.n754 B.n367 163.367
R830 B.n754 B.n361 163.367
R831 B.n762 B.n361 163.367
R832 B.n762 B.n359 163.367
R833 B.n766 B.n359 163.367
R834 B.n766 B.n353 163.367
R835 B.n775 B.n353 163.367
R836 B.n775 B.n351 163.367
R837 B.n779 B.n351 163.367
R838 B.n779 B.n3 163.367
R839 B.n885 B.n3 163.367
R840 B.n881 B.n2 163.367
R841 B.n881 B.n880 163.367
R842 B.n880 B.n9 163.367
R843 B.n876 B.n9 163.367
R844 B.n876 B.n11 163.367
R845 B.n872 B.n11 163.367
R846 B.n872 B.n17 163.367
R847 B.n868 B.n17 163.367
R848 B.n868 B.n19 163.367
R849 B.n864 B.n19 163.367
R850 B.n864 B.n24 163.367
R851 B.n860 B.n24 163.367
R852 B.n860 B.n26 163.367
R853 B.n856 B.n26 163.367
R854 B.n856 B.n31 163.367
R855 B.n852 B.n31 163.367
R856 B.n852 B.n33 163.367
R857 B.n848 B.n33 163.367
R858 B.n848 B.n38 163.367
R859 B.n844 B.n38 163.367
R860 B.n844 B.n40 163.367
R861 B.n840 B.n40 163.367
R862 B.n840 B.n44 163.367
R863 B.n836 B.n44 163.367
R864 B.n836 B.n46 163.367
R865 B.n832 B.n46 163.367
R866 B.n832 B.n52 163.367
R867 B.n828 B.n52 163.367
R868 B.n828 B.n54 163.367
R869 B.n115 B.t10 116.084
R870 B.n465 B.t7 116.084
R871 B.n118 B.t16 116.062
R872 B.n462 B.t14 116.062
R873 B.n120 B.n57 71.676
R874 B.n124 B.n58 71.676
R875 B.n128 B.n59 71.676
R876 B.n132 B.n60 71.676
R877 B.n136 B.n61 71.676
R878 B.n140 B.n62 71.676
R879 B.n144 B.n63 71.676
R880 B.n148 B.n64 71.676
R881 B.n152 B.n65 71.676
R882 B.n156 B.n66 71.676
R883 B.n160 B.n67 71.676
R884 B.n164 B.n68 71.676
R885 B.n168 B.n69 71.676
R886 B.n172 B.n70 71.676
R887 B.n176 B.n71 71.676
R888 B.n180 B.n72 71.676
R889 B.n184 B.n73 71.676
R890 B.n188 B.n74 71.676
R891 B.n192 B.n75 71.676
R892 B.n196 B.n76 71.676
R893 B.n200 B.n77 71.676
R894 B.n204 B.n78 71.676
R895 B.n208 B.n79 71.676
R896 B.n212 B.n80 71.676
R897 B.n216 B.n81 71.676
R898 B.n220 B.n82 71.676
R899 B.n224 B.n83 71.676
R900 B.n229 B.n84 71.676
R901 B.n233 B.n85 71.676
R902 B.n237 B.n86 71.676
R903 B.n241 B.n87 71.676
R904 B.n245 B.n88 71.676
R905 B.n249 B.n89 71.676
R906 B.n253 B.n90 71.676
R907 B.n257 B.n91 71.676
R908 B.n261 B.n92 71.676
R909 B.n265 B.n93 71.676
R910 B.n269 B.n94 71.676
R911 B.n273 B.n95 71.676
R912 B.n277 B.n96 71.676
R913 B.n281 B.n97 71.676
R914 B.n285 B.n98 71.676
R915 B.n289 B.n99 71.676
R916 B.n293 B.n100 71.676
R917 B.n297 B.n101 71.676
R918 B.n301 B.n102 71.676
R919 B.n305 B.n103 71.676
R920 B.n309 B.n104 71.676
R921 B.n313 B.n105 71.676
R922 B.n317 B.n106 71.676
R923 B.n321 B.n107 71.676
R924 B.n325 B.n108 71.676
R925 B.n329 B.n109 71.676
R926 B.n333 B.n110 71.676
R927 B.n337 B.n111 71.676
R928 B.n341 B.n112 71.676
R929 B.n345 B.n113 71.676
R930 B.n114 B.n113 71.676
R931 B.n344 B.n112 71.676
R932 B.n340 B.n111 71.676
R933 B.n336 B.n110 71.676
R934 B.n332 B.n109 71.676
R935 B.n328 B.n108 71.676
R936 B.n324 B.n107 71.676
R937 B.n320 B.n106 71.676
R938 B.n316 B.n105 71.676
R939 B.n312 B.n104 71.676
R940 B.n308 B.n103 71.676
R941 B.n304 B.n102 71.676
R942 B.n300 B.n101 71.676
R943 B.n296 B.n100 71.676
R944 B.n292 B.n99 71.676
R945 B.n288 B.n98 71.676
R946 B.n284 B.n97 71.676
R947 B.n280 B.n96 71.676
R948 B.n276 B.n95 71.676
R949 B.n272 B.n94 71.676
R950 B.n268 B.n93 71.676
R951 B.n264 B.n92 71.676
R952 B.n260 B.n91 71.676
R953 B.n256 B.n90 71.676
R954 B.n252 B.n89 71.676
R955 B.n248 B.n88 71.676
R956 B.n244 B.n87 71.676
R957 B.n240 B.n86 71.676
R958 B.n236 B.n85 71.676
R959 B.n232 B.n84 71.676
R960 B.n228 B.n83 71.676
R961 B.n223 B.n82 71.676
R962 B.n219 B.n81 71.676
R963 B.n215 B.n80 71.676
R964 B.n211 B.n79 71.676
R965 B.n207 B.n78 71.676
R966 B.n203 B.n77 71.676
R967 B.n199 B.n76 71.676
R968 B.n195 B.n75 71.676
R969 B.n191 B.n74 71.676
R970 B.n187 B.n73 71.676
R971 B.n183 B.n72 71.676
R972 B.n179 B.n71 71.676
R973 B.n175 B.n70 71.676
R974 B.n171 B.n69 71.676
R975 B.n167 B.n68 71.676
R976 B.n163 B.n67 71.676
R977 B.n159 B.n66 71.676
R978 B.n155 B.n65 71.676
R979 B.n151 B.n64 71.676
R980 B.n147 B.n63 71.676
R981 B.n143 B.n62 71.676
R982 B.n139 B.n61 71.676
R983 B.n135 B.n60 71.676
R984 B.n131 B.n59 71.676
R985 B.n127 B.n58 71.676
R986 B.n123 B.n57 71.676
R987 B.n692 B.n691 71.676
R988 B.n686 B.n405 71.676
R989 B.n683 B.n406 71.676
R990 B.n679 B.n407 71.676
R991 B.n675 B.n408 71.676
R992 B.n671 B.n409 71.676
R993 B.n667 B.n410 71.676
R994 B.n663 B.n411 71.676
R995 B.n659 B.n412 71.676
R996 B.n655 B.n413 71.676
R997 B.n651 B.n414 71.676
R998 B.n647 B.n415 71.676
R999 B.n643 B.n416 71.676
R1000 B.n639 B.n417 71.676
R1001 B.n635 B.n418 71.676
R1002 B.n631 B.n419 71.676
R1003 B.n627 B.n420 71.676
R1004 B.n623 B.n421 71.676
R1005 B.n619 B.n422 71.676
R1006 B.n615 B.n423 71.676
R1007 B.n611 B.n424 71.676
R1008 B.n607 B.n425 71.676
R1009 B.n603 B.n426 71.676
R1010 B.n599 B.n427 71.676
R1011 B.n595 B.n428 71.676
R1012 B.n591 B.n429 71.676
R1013 B.n587 B.n430 71.676
R1014 B.n583 B.n431 71.676
R1015 B.n579 B.n432 71.676
R1016 B.n575 B.n433 71.676
R1017 B.n571 B.n434 71.676
R1018 B.n566 B.n435 71.676
R1019 B.n562 B.n436 71.676
R1020 B.n558 B.n437 71.676
R1021 B.n554 B.n438 71.676
R1022 B.n550 B.n439 71.676
R1023 B.n546 B.n440 71.676
R1024 B.n542 B.n441 71.676
R1025 B.n538 B.n442 71.676
R1026 B.n534 B.n443 71.676
R1027 B.n530 B.n444 71.676
R1028 B.n526 B.n445 71.676
R1029 B.n522 B.n446 71.676
R1030 B.n518 B.n447 71.676
R1031 B.n514 B.n448 71.676
R1032 B.n510 B.n449 71.676
R1033 B.n506 B.n450 71.676
R1034 B.n502 B.n451 71.676
R1035 B.n498 B.n452 71.676
R1036 B.n494 B.n453 71.676
R1037 B.n490 B.n454 71.676
R1038 B.n486 B.n455 71.676
R1039 B.n482 B.n456 71.676
R1040 B.n478 B.n457 71.676
R1041 B.n474 B.n458 71.676
R1042 B.n470 B.n459 71.676
R1043 B.n694 B.n404 71.676
R1044 B.n692 B.n461 71.676
R1045 B.n684 B.n405 71.676
R1046 B.n680 B.n406 71.676
R1047 B.n676 B.n407 71.676
R1048 B.n672 B.n408 71.676
R1049 B.n668 B.n409 71.676
R1050 B.n664 B.n410 71.676
R1051 B.n660 B.n411 71.676
R1052 B.n656 B.n412 71.676
R1053 B.n652 B.n413 71.676
R1054 B.n648 B.n414 71.676
R1055 B.n644 B.n415 71.676
R1056 B.n640 B.n416 71.676
R1057 B.n636 B.n417 71.676
R1058 B.n632 B.n418 71.676
R1059 B.n628 B.n419 71.676
R1060 B.n624 B.n420 71.676
R1061 B.n620 B.n421 71.676
R1062 B.n616 B.n422 71.676
R1063 B.n612 B.n423 71.676
R1064 B.n608 B.n424 71.676
R1065 B.n604 B.n425 71.676
R1066 B.n600 B.n426 71.676
R1067 B.n596 B.n427 71.676
R1068 B.n592 B.n428 71.676
R1069 B.n588 B.n429 71.676
R1070 B.n584 B.n430 71.676
R1071 B.n580 B.n431 71.676
R1072 B.n576 B.n432 71.676
R1073 B.n572 B.n433 71.676
R1074 B.n567 B.n434 71.676
R1075 B.n563 B.n435 71.676
R1076 B.n559 B.n436 71.676
R1077 B.n555 B.n437 71.676
R1078 B.n551 B.n438 71.676
R1079 B.n547 B.n439 71.676
R1080 B.n543 B.n440 71.676
R1081 B.n539 B.n441 71.676
R1082 B.n535 B.n442 71.676
R1083 B.n531 B.n443 71.676
R1084 B.n527 B.n444 71.676
R1085 B.n523 B.n445 71.676
R1086 B.n519 B.n446 71.676
R1087 B.n515 B.n447 71.676
R1088 B.n511 B.n448 71.676
R1089 B.n507 B.n449 71.676
R1090 B.n503 B.n450 71.676
R1091 B.n499 B.n451 71.676
R1092 B.n495 B.n452 71.676
R1093 B.n491 B.n453 71.676
R1094 B.n487 B.n454 71.676
R1095 B.n483 B.n455 71.676
R1096 B.n479 B.n456 71.676
R1097 B.n475 B.n457 71.676
R1098 B.n471 B.n458 71.676
R1099 B.n467 B.n459 71.676
R1100 B.n695 B.n694 71.676
R1101 B.n886 B.n885 71.676
R1102 B.n886 B.n2 71.676
R1103 B.n116 B.t11 68.9564
R1104 B.n466 B.t6 68.9564
R1105 B.n119 B.t17 68.9357
R1106 B.n463 B.t13 68.9357
R1107 B.n693 B.n401 66.5401
R1108 B.n826 B.n825 66.5401
R1109 B.n226 B.n119 59.5399
R1110 B.n117 B.n116 59.5399
R1111 B.n569 B.n466 59.5399
R1112 B.n464 B.n463 59.5399
R1113 B.n119 B.n118 47.1278
R1114 B.n116 B.n115 47.1278
R1115 B.n466 B.n465 47.1278
R1116 B.n463 B.n462 47.1278
R1117 B.n700 B.n401 35.628
R1118 B.n700 B.n397 35.628
R1119 B.n706 B.n397 35.628
R1120 B.n706 B.n393 35.628
R1121 B.n713 B.n393 35.628
R1122 B.n713 B.n712 35.628
R1123 B.n719 B.n386 35.628
R1124 B.n725 B.n386 35.628
R1125 B.n725 B.n382 35.628
R1126 B.n731 B.n382 35.628
R1127 B.n731 B.n378 35.628
R1128 B.n737 B.n378 35.628
R1129 B.n737 B.n374 35.628
R1130 B.n743 B.n374 35.628
R1131 B.n743 B.n370 35.628
R1132 B.n749 B.n370 35.628
R1133 B.n755 B.n366 35.628
R1134 B.n755 B.n362 35.628
R1135 B.n761 B.n362 35.628
R1136 B.n761 B.n357 35.628
R1137 B.n767 B.n357 35.628
R1138 B.n767 B.n358 35.628
R1139 B.n774 B.n350 35.628
R1140 B.n780 B.n350 35.628
R1141 B.n780 B.n4 35.628
R1142 B.n884 B.n4 35.628
R1143 B.n884 B.n883 35.628
R1144 B.n883 B.n882 35.628
R1145 B.n882 B.n8 35.628
R1146 B.n12 B.n8 35.628
R1147 B.n875 B.n12 35.628
R1148 B.n874 B.n873 35.628
R1149 B.n873 B.n16 35.628
R1150 B.n867 B.n16 35.628
R1151 B.n867 B.n866 35.628
R1152 B.n866 B.n865 35.628
R1153 B.n865 B.n23 35.628
R1154 B.n859 B.n858 35.628
R1155 B.n858 B.n857 35.628
R1156 B.n857 B.n30 35.628
R1157 B.n851 B.n30 35.628
R1158 B.n851 B.n850 35.628
R1159 B.n850 B.n849 35.628
R1160 B.n849 B.n37 35.628
R1161 B.n843 B.n37 35.628
R1162 B.n843 B.n842 35.628
R1163 B.n842 B.n841 35.628
R1164 B.n835 B.n47 35.628
R1165 B.n835 B.n834 35.628
R1166 B.n834 B.n833 35.628
R1167 B.n833 B.n51 35.628
R1168 B.n827 B.n51 35.628
R1169 B.n827 B.n826 35.628
R1170 B.n690 B.n399 31.3761
R1171 B.n697 B.n696 31.3761
R1172 B.n823 B.n822 31.3761
R1173 B.n121 B.n53 31.3761
R1174 B.n712 B.t5 29.3408
R1175 B.t0 B.n366 29.3408
R1176 B.t2 B.n23 29.3408
R1177 B.n47 B.t9 29.3408
R1178 B.n774 B.t3 24.1015
R1179 B.n875 B.t1 24.1015
R1180 B B.n887 18.0485
R1181 B.n358 B.t3 11.5271
R1182 B.t1 B.n874 11.5271
R1183 B.n702 B.n399 10.6151
R1184 B.n703 B.n702 10.6151
R1185 B.n704 B.n703 10.6151
R1186 B.n704 B.n391 10.6151
R1187 B.n715 B.n391 10.6151
R1188 B.n716 B.n715 10.6151
R1189 B.n717 B.n716 10.6151
R1190 B.n717 B.n384 10.6151
R1191 B.n727 B.n384 10.6151
R1192 B.n728 B.n727 10.6151
R1193 B.n729 B.n728 10.6151
R1194 B.n729 B.n376 10.6151
R1195 B.n739 B.n376 10.6151
R1196 B.n740 B.n739 10.6151
R1197 B.n741 B.n740 10.6151
R1198 B.n741 B.n368 10.6151
R1199 B.n751 B.n368 10.6151
R1200 B.n752 B.n751 10.6151
R1201 B.n753 B.n752 10.6151
R1202 B.n753 B.n360 10.6151
R1203 B.n763 B.n360 10.6151
R1204 B.n764 B.n763 10.6151
R1205 B.n765 B.n764 10.6151
R1206 B.n765 B.n352 10.6151
R1207 B.n776 B.n352 10.6151
R1208 B.n777 B.n776 10.6151
R1209 B.n778 B.n777 10.6151
R1210 B.n778 B.n0 10.6151
R1211 B.n690 B.n689 10.6151
R1212 B.n689 B.n688 10.6151
R1213 B.n688 B.n687 10.6151
R1214 B.n687 B.n685 10.6151
R1215 B.n685 B.n682 10.6151
R1216 B.n682 B.n681 10.6151
R1217 B.n681 B.n678 10.6151
R1218 B.n678 B.n677 10.6151
R1219 B.n677 B.n674 10.6151
R1220 B.n674 B.n673 10.6151
R1221 B.n673 B.n670 10.6151
R1222 B.n670 B.n669 10.6151
R1223 B.n669 B.n666 10.6151
R1224 B.n666 B.n665 10.6151
R1225 B.n665 B.n662 10.6151
R1226 B.n662 B.n661 10.6151
R1227 B.n661 B.n658 10.6151
R1228 B.n658 B.n657 10.6151
R1229 B.n657 B.n654 10.6151
R1230 B.n654 B.n653 10.6151
R1231 B.n653 B.n650 10.6151
R1232 B.n650 B.n649 10.6151
R1233 B.n649 B.n646 10.6151
R1234 B.n646 B.n645 10.6151
R1235 B.n645 B.n642 10.6151
R1236 B.n642 B.n641 10.6151
R1237 B.n641 B.n638 10.6151
R1238 B.n638 B.n637 10.6151
R1239 B.n637 B.n634 10.6151
R1240 B.n634 B.n633 10.6151
R1241 B.n633 B.n630 10.6151
R1242 B.n630 B.n629 10.6151
R1243 B.n629 B.n626 10.6151
R1244 B.n626 B.n625 10.6151
R1245 B.n625 B.n622 10.6151
R1246 B.n622 B.n621 10.6151
R1247 B.n621 B.n618 10.6151
R1248 B.n618 B.n617 10.6151
R1249 B.n617 B.n614 10.6151
R1250 B.n614 B.n613 10.6151
R1251 B.n613 B.n610 10.6151
R1252 B.n610 B.n609 10.6151
R1253 B.n609 B.n606 10.6151
R1254 B.n606 B.n605 10.6151
R1255 B.n605 B.n602 10.6151
R1256 B.n602 B.n601 10.6151
R1257 B.n601 B.n598 10.6151
R1258 B.n598 B.n597 10.6151
R1259 B.n597 B.n594 10.6151
R1260 B.n594 B.n593 10.6151
R1261 B.n593 B.n590 10.6151
R1262 B.n590 B.n589 10.6151
R1263 B.n586 B.n585 10.6151
R1264 B.n585 B.n582 10.6151
R1265 B.n582 B.n581 10.6151
R1266 B.n581 B.n578 10.6151
R1267 B.n578 B.n577 10.6151
R1268 B.n577 B.n574 10.6151
R1269 B.n574 B.n573 10.6151
R1270 B.n573 B.n570 10.6151
R1271 B.n568 B.n565 10.6151
R1272 B.n565 B.n564 10.6151
R1273 B.n564 B.n561 10.6151
R1274 B.n561 B.n560 10.6151
R1275 B.n560 B.n557 10.6151
R1276 B.n557 B.n556 10.6151
R1277 B.n556 B.n553 10.6151
R1278 B.n553 B.n552 10.6151
R1279 B.n552 B.n549 10.6151
R1280 B.n549 B.n548 10.6151
R1281 B.n548 B.n545 10.6151
R1282 B.n545 B.n544 10.6151
R1283 B.n544 B.n541 10.6151
R1284 B.n541 B.n540 10.6151
R1285 B.n540 B.n537 10.6151
R1286 B.n537 B.n536 10.6151
R1287 B.n536 B.n533 10.6151
R1288 B.n533 B.n532 10.6151
R1289 B.n532 B.n529 10.6151
R1290 B.n529 B.n528 10.6151
R1291 B.n528 B.n525 10.6151
R1292 B.n525 B.n524 10.6151
R1293 B.n524 B.n521 10.6151
R1294 B.n521 B.n520 10.6151
R1295 B.n520 B.n517 10.6151
R1296 B.n517 B.n516 10.6151
R1297 B.n516 B.n513 10.6151
R1298 B.n513 B.n512 10.6151
R1299 B.n512 B.n509 10.6151
R1300 B.n509 B.n508 10.6151
R1301 B.n508 B.n505 10.6151
R1302 B.n505 B.n504 10.6151
R1303 B.n504 B.n501 10.6151
R1304 B.n501 B.n500 10.6151
R1305 B.n500 B.n497 10.6151
R1306 B.n497 B.n496 10.6151
R1307 B.n496 B.n493 10.6151
R1308 B.n493 B.n492 10.6151
R1309 B.n492 B.n489 10.6151
R1310 B.n489 B.n488 10.6151
R1311 B.n488 B.n485 10.6151
R1312 B.n485 B.n484 10.6151
R1313 B.n484 B.n481 10.6151
R1314 B.n481 B.n480 10.6151
R1315 B.n480 B.n477 10.6151
R1316 B.n477 B.n476 10.6151
R1317 B.n476 B.n473 10.6151
R1318 B.n473 B.n472 10.6151
R1319 B.n472 B.n469 10.6151
R1320 B.n469 B.n468 10.6151
R1321 B.n468 B.n403 10.6151
R1322 B.n696 B.n403 10.6151
R1323 B.n698 B.n697 10.6151
R1324 B.n698 B.n395 10.6151
R1325 B.n708 B.n395 10.6151
R1326 B.n709 B.n708 10.6151
R1327 B.n710 B.n709 10.6151
R1328 B.n710 B.n388 10.6151
R1329 B.n721 B.n388 10.6151
R1330 B.n722 B.n721 10.6151
R1331 B.n723 B.n722 10.6151
R1332 B.n723 B.n380 10.6151
R1333 B.n733 B.n380 10.6151
R1334 B.n734 B.n733 10.6151
R1335 B.n735 B.n734 10.6151
R1336 B.n735 B.n372 10.6151
R1337 B.n745 B.n372 10.6151
R1338 B.n746 B.n745 10.6151
R1339 B.n747 B.n746 10.6151
R1340 B.n747 B.n364 10.6151
R1341 B.n757 B.n364 10.6151
R1342 B.n758 B.n757 10.6151
R1343 B.n759 B.n758 10.6151
R1344 B.n759 B.n355 10.6151
R1345 B.n769 B.n355 10.6151
R1346 B.n770 B.n769 10.6151
R1347 B.n772 B.n770 10.6151
R1348 B.n772 B.n771 10.6151
R1349 B.n771 B.n348 10.6151
R1350 B.n783 B.n348 10.6151
R1351 B.n784 B.n783 10.6151
R1352 B.n785 B.n784 10.6151
R1353 B.n786 B.n785 10.6151
R1354 B.n787 B.n786 10.6151
R1355 B.n790 B.n787 10.6151
R1356 B.n791 B.n790 10.6151
R1357 B.n792 B.n791 10.6151
R1358 B.n793 B.n792 10.6151
R1359 B.n795 B.n793 10.6151
R1360 B.n796 B.n795 10.6151
R1361 B.n797 B.n796 10.6151
R1362 B.n798 B.n797 10.6151
R1363 B.n800 B.n798 10.6151
R1364 B.n801 B.n800 10.6151
R1365 B.n802 B.n801 10.6151
R1366 B.n803 B.n802 10.6151
R1367 B.n805 B.n803 10.6151
R1368 B.n806 B.n805 10.6151
R1369 B.n807 B.n806 10.6151
R1370 B.n808 B.n807 10.6151
R1371 B.n810 B.n808 10.6151
R1372 B.n811 B.n810 10.6151
R1373 B.n812 B.n811 10.6151
R1374 B.n813 B.n812 10.6151
R1375 B.n815 B.n813 10.6151
R1376 B.n816 B.n815 10.6151
R1377 B.n817 B.n816 10.6151
R1378 B.n818 B.n817 10.6151
R1379 B.n820 B.n818 10.6151
R1380 B.n821 B.n820 10.6151
R1381 B.n822 B.n821 10.6151
R1382 B.n879 B.n1 10.6151
R1383 B.n879 B.n878 10.6151
R1384 B.n878 B.n877 10.6151
R1385 B.n877 B.n10 10.6151
R1386 B.n871 B.n10 10.6151
R1387 B.n871 B.n870 10.6151
R1388 B.n870 B.n869 10.6151
R1389 B.n869 B.n18 10.6151
R1390 B.n863 B.n18 10.6151
R1391 B.n863 B.n862 10.6151
R1392 B.n862 B.n861 10.6151
R1393 B.n861 B.n25 10.6151
R1394 B.n855 B.n25 10.6151
R1395 B.n855 B.n854 10.6151
R1396 B.n854 B.n853 10.6151
R1397 B.n853 B.n32 10.6151
R1398 B.n847 B.n32 10.6151
R1399 B.n847 B.n846 10.6151
R1400 B.n846 B.n845 10.6151
R1401 B.n845 B.n39 10.6151
R1402 B.n839 B.n39 10.6151
R1403 B.n839 B.n838 10.6151
R1404 B.n838 B.n837 10.6151
R1405 B.n837 B.n45 10.6151
R1406 B.n831 B.n45 10.6151
R1407 B.n831 B.n830 10.6151
R1408 B.n830 B.n829 10.6151
R1409 B.n829 B.n53 10.6151
R1410 B.n122 B.n121 10.6151
R1411 B.n125 B.n122 10.6151
R1412 B.n126 B.n125 10.6151
R1413 B.n129 B.n126 10.6151
R1414 B.n130 B.n129 10.6151
R1415 B.n133 B.n130 10.6151
R1416 B.n134 B.n133 10.6151
R1417 B.n137 B.n134 10.6151
R1418 B.n138 B.n137 10.6151
R1419 B.n141 B.n138 10.6151
R1420 B.n142 B.n141 10.6151
R1421 B.n145 B.n142 10.6151
R1422 B.n146 B.n145 10.6151
R1423 B.n149 B.n146 10.6151
R1424 B.n150 B.n149 10.6151
R1425 B.n153 B.n150 10.6151
R1426 B.n154 B.n153 10.6151
R1427 B.n157 B.n154 10.6151
R1428 B.n158 B.n157 10.6151
R1429 B.n161 B.n158 10.6151
R1430 B.n162 B.n161 10.6151
R1431 B.n165 B.n162 10.6151
R1432 B.n166 B.n165 10.6151
R1433 B.n169 B.n166 10.6151
R1434 B.n170 B.n169 10.6151
R1435 B.n173 B.n170 10.6151
R1436 B.n174 B.n173 10.6151
R1437 B.n177 B.n174 10.6151
R1438 B.n178 B.n177 10.6151
R1439 B.n181 B.n178 10.6151
R1440 B.n182 B.n181 10.6151
R1441 B.n185 B.n182 10.6151
R1442 B.n186 B.n185 10.6151
R1443 B.n189 B.n186 10.6151
R1444 B.n190 B.n189 10.6151
R1445 B.n193 B.n190 10.6151
R1446 B.n194 B.n193 10.6151
R1447 B.n197 B.n194 10.6151
R1448 B.n198 B.n197 10.6151
R1449 B.n201 B.n198 10.6151
R1450 B.n202 B.n201 10.6151
R1451 B.n205 B.n202 10.6151
R1452 B.n206 B.n205 10.6151
R1453 B.n209 B.n206 10.6151
R1454 B.n210 B.n209 10.6151
R1455 B.n213 B.n210 10.6151
R1456 B.n214 B.n213 10.6151
R1457 B.n217 B.n214 10.6151
R1458 B.n218 B.n217 10.6151
R1459 B.n221 B.n218 10.6151
R1460 B.n222 B.n221 10.6151
R1461 B.n225 B.n222 10.6151
R1462 B.n230 B.n227 10.6151
R1463 B.n231 B.n230 10.6151
R1464 B.n234 B.n231 10.6151
R1465 B.n235 B.n234 10.6151
R1466 B.n238 B.n235 10.6151
R1467 B.n239 B.n238 10.6151
R1468 B.n242 B.n239 10.6151
R1469 B.n243 B.n242 10.6151
R1470 B.n247 B.n246 10.6151
R1471 B.n250 B.n247 10.6151
R1472 B.n251 B.n250 10.6151
R1473 B.n254 B.n251 10.6151
R1474 B.n255 B.n254 10.6151
R1475 B.n258 B.n255 10.6151
R1476 B.n259 B.n258 10.6151
R1477 B.n262 B.n259 10.6151
R1478 B.n263 B.n262 10.6151
R1479 B.n266 B.n263 10.6151
R1480 B.n267 B.n266 10.6151
R1481 B.n270 B.n267 10.6151
R1482 B.n271 B.n270 10.6151
R1483 B.n274 B.n271 10.6151
R1484 B.n275 B.n274 10.6151
R1485 B.n278 B.n275 10.6151
R1486 B.n279 B.n278 10.6151
R1487 B.n282 B.n279 10.6151
R1488 B.n283 B.n282 10.6151
R1489 B.n286 B.n283 10.6151
R1490 B.n287 B.n286 10.6151
R1491 B.n290 B.n287 10.6151
R1492 B.n291 B.n290 10.6151
R1493 B.n294 B.n291 10.6151
R1494 B.n295 B.n294 10.6151
R1495 B.n298 B.n295 10.6151
R1496 B.n299 B.n298 10.6151
R1497 B.n302 B.n299 10.6151
R1498 B.n303 B.n302 10.6151
R1499 B.n306 B.n303 10.6151
R1500 B.n307 B.n306 10.6151
R1501 B.n310 B.n307 10.6151
R1502 B.n311 B.n310 10.6151
R1503 B.n314 B.n311 10.6151
R1504 B.n315 B.n314 10.6151
R1505 B.n318 B.n315 10.6151
R1506 B.n319 B.n318 10.6151
R1507 B.n322 B.n319 10.6151
R1508 B.n323 B.n322 10.6151
R1509 B.n326 B.n323 10.6151
R1510 B.n327 B.n326 10.6151
R1511 B.n330 B.n327 10.6151
R1512 B.n331 B.n330 10.6151
R1513 B.n334 B.n331 10.6151
R1514 B.n335 B.n334 10.6151
R1515 B.n338 B.n335 10.6151
R1516 B.n339 B.n338 10.6151
R1517 B.n342 B.n339 10.6151
R1518 B.n343 B.n342 10.6151
R1519 B.n346 B.n343 10.6151
R1520 B.n347 B.n346 10.6151
R1521 B.n823 B.n347 10.6151
R1522 B.n887 B.n0 8.11757
R1523 B.n887 B.n1 8.11757
R1524 B.n586 B.n464 6.5566
R1525 B.n570 B.n569 6.5566
R1526 B.n227 B.n226 6.5566
R1527 B.n243 B.n117 6.5566
R1528 B.n719 B.t5 6.28771
R1529 B.n749 B.t0 6.28771
R1530 B.n859 B.t2 6.28771
R1531 B.n841 B.t9 6.28771
R1532 B.n589 B.n464 4.05904
R1533 B.n569 B.n568 4.05904
R1534 B.n226 B.n225 4.05904
R1535 B.n246 B.n117 4.05904
R1536 VN.n0 VN.t0 216.589
R1537 VN.n1 VN.t2 216.589
R1538 VN.n0 VN.t1 216.041
R1539 VN.n1 VN.t3 216.041
R1540 VN VN.n1 54.7997
R1541 VN VN.n0 6.88683
R1542 VDD2.n2 VDD2.n0 104.359
R1543 VDD2.n2 VDD2.n1 60.8081
R1544 VDD2.n1 VDD2.t0 1.26004
R1545 VDD2.n1 VDD2.t1 1.26004
R1546 VDD2.n0 VDD2.t3 1.26004
R1547 VDD2.n0 VDD2.t2 1.26004
R1548 VDD2 VDD2.n2 0.0586897
C0 VP VDD2 0.36295f
C1 VP VN 6.51397f
C2 VDD2 VDD1 0.908845f
C3 VTAIL VDD2 6.38914f
C4 VN VDD1 0.149009f
C5 VTAIL VN 5.5541f
C6 VP VDD1 6.08014f
C7 VTAIL VP 5.56821f
C8 VTAIL VDD1 6.33828f
C9 VDD2 VN 5.86681f
C10 VDD2 B 3.773211f
C11 VDD1 B 8.10859f
C12 VTAIL B 12.000009f
C13 VN B 10.11609f
C14 VP B 8.123648f
C15 VDD2.t3 B 0.330783f
C16 VDD2.t2 B 0.330783f
C17 VDD2.n0 B 3.7788f
C18 VDD2.t0 B 0.330783f
C19 VDD2.t1 B 0.330783f
C20 VDD2.n1 B 2.99622f
C21 VDD2.n2 B 4.01638f
C22 VN.t0 B 2.74298f
C23 VN.t1 B 2.74033f
C24 VN.n0 B 1.83683f
C25 VN.t2 B 2.74298f
C26 VN.t3 B 2.74033f
C27 VN.n1 B 3.29627f
C28 VTAIL.t1 B 2.16548f
C29 VTAIL.n0 B 0.288428f
C30 VTAIL.t4 B 2.16548f
C31 VTAIL.n1 B 0.337827f
C32 VTAIL.t7 B 2.16548f
C33 VTAIL.n2 B 1.30621f
C34 VTAIL.t0 B 2.1655f
C35 VTAIL.n3 B 1.3062f
C36 VTAIL.t3 B 2.1655f
C37 VTAIL.n4 B 0.337812f
C38 VTAIL.t6 B 2.1655f
C39 VTAIL.n5 B 0.337812f
C40 VTAIL.t5 B 2.16548f
C41 VTAIL.n6 B 1.30621f
C42 VTAIL.t2 B 2.16548f
C43 VTAIL.n7 B 1.251f
C44 VDD1.t0 B 0.330827f
C45 VDD1.t1 B 0.330827f
C46 VDD1.n0 B 2.99701f
C47 VDD1.t3 B 0.330827f
C48 VDD1.t2 B 0.330827f
C49 VDD1.n1 B 3.80697f
C50 VP.n0 B 0.037859f
C51 VP.t3 B 2.60048f
C52 VP.n1 B 0.041745f
C53 VP.t2 B 2.77692f
C54 VP.t1 B 2.77961f
C55 VP.n2 B 3.3256f
C56 VP.n3 B 1.70878f
C57 VP.t0 B 2.60048f
C58 VP.n4 B 1.00915f
C59 VP.n5 B 0.051414f
C60 VP.n6 B 0.037859f
C61 VP.n7 B 0.028718f
C62 VP.n8 B 0.028718f
C63 VP.n9 B 0.041745f
C64 VP.n10 B 0.051414f
C65 VP.n11 B 1.00915f
C66 VP.n12 B 0.032542f
.ends

