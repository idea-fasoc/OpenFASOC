* NGSPICE file created from diff_pair_sample_1606.ext - technology: sky130A

.subckt diff_pair_sample_1606 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=0.1287 pd=1.11 as=0.3042 ps=2.34 w=0.78 l=1.9
X1 VTAIL.t10 VN.t1 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.3042 pd=2.34 as=0.1287 ps=1.11 w=0.78 l=1.9
X2 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=0.3042 pd=2.34 as=0 ps=0 w=0.78 l=1.9
X3 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=0.3042 pd=2.34 as=0 ps=0 w=0.78 l=1.9
X4 VDD1.t7 VP.t0 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.1287 pd=1.11 as=0.3042 ps=2.34 w=0.78 l=1.9
X5 VTAIL.t11 VN.t2 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=0.3042 pd=2.34 as=0.1287 ps=1.11 w=0.78 l=1.9
X6 VTAIL.t15 VN.t3 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=0.1287 pd=1.11 as=0.1287 ps=1.11 w=0.78 l=1.9
X7 VDD2.t3 VN.t4 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=0.1287 pd=1.11 as=0.1287 ps=1.11 w=0.78 l=1.9
X8 VDD1.t6 VP.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.1287 pd=1.11 as=0.3042 ps=2.34 w=0.78 l=1.9
X9 VTAIL.t7 VP.t2 VDD1.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=0.3042 pd=2.34 as=0.1287 ps=1.11 w=0.78 l=1.9
X10 VDD2.t2 VN.t5 VTAIL.t9 B.t6 sky130_fd_pr__nfet_01v8 ad=0.1287 pd=1.11 as=0.3042 ps=2.34 w=0.78 l=1.9
X11 VDD2.t1 VN.t6 VTAIL.t14 B.t4 sky130_fd_pr__nfet_01v8 ad=0.1287 pd=1.11 as=0.1287 ps=1.11 w=0.78 l=1.9
X12 VTAIL.t1 VP.t3 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.1287 pd=1.11 as=0.1287 ps=1.11 w=0.78 l=1.9
X13 VDD1.t3 VP.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.1287 pd=1.11 as=0.1287 ps=1.11 w=0.78 l=1.9
X14 VTAIL.t0 VP.t5 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.1287 pd=1.11 as=0.1287 ps=1.11 w=0.78 l=1.9
X15 VTAIL.t2 VP.t6 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.3042 pd=2.34 as=0.1287 ps=1.11 w=0.78 l=1.9
X16 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=0.3042 pd=2.34 as=0 ps=0 w=0.78 l=1.9
X17 VTAIL.t12 VN.t7 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.1287 pd=1.11 as=0.1287 ps=1.11 w=0.78 l=1.9
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.3042 pd=2.34 as=0 ps=0 w=0.78 l=1.9
X19 VDD1.t0 VP.t7 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.1287 pd=1.11 as=0.1287 ps=1.11 w=0.78 l=1.9
R0 VN.n22 VN.n21 181.22
R1 VN.n45 VN.n44 181.22
R2 VN.n43 VN.n23 161.3
R3 VN.n42 VN.n41 161.3
R4 VN.n40 VN.n24 161.3
R5 VN.n39 VN.n38 161.3
R6 VN.n37 VN.n25 161.3
R7 VN.n35 VN.n34 161.3
R8 VN.n33 VN.n26 161.3
R9 VN.n32 VN.n31 161.3
R10 VN.n30 VN.n27 161.3
R11 VN.n20 VN.n0 161.3
R12 VN.n19 VN.n18 161.3
R13 VN.n17 VN.n1 161.3
R14 VN.n16 VN.n15 161.3
R15 VN.n14 VN.n2 161.3
R16 VN.n12 VN.n11 161.3
R17 VN.n10 VN.n3 161.3
R18 VN.n9 VN.n8 161.3
R19 VN.n7 VN.n4 161.3
R20 VN.n8 VN.n3 56.5617
R21 VN.n31 VN.n26 56.5617
R22 VN.n6 VN.n5 51.8866
R23 VN.n29 VN.n28 51.8866
R24 VN.n5 VN.t1 44.7858
R25 VN.n28 VN.t5 44.7858
R26 VN.n15 VN.n1 42.5146
R27 VN.n38 VN.n24 42.5146
R28 VN VN.n45 39.4418
R29 VN.n19 VN.n1 38.6395
R30 VN.n42 VN.n24 38.6395
R31 VN.n8 VN.n7 24.5923
R32 VN.n12 VN.n3 24.5923
R33 VN.n15 VN.n14 24.5923
R34 VN.n20 VN.n19 24.5923
R35 VN.n31 VN.n30 24.5923
R36 VN.n38 VN.n37 24.5923
R37 VN.n35 VN.n26 24.5923
R38 VN.n43 VN.n42 24.5923
R39 VN.n7 VN.n6 17.9525
R40 VN.n13 VN.n12 17.9525
R41 VN.n30 VN.n29 17.9525
R42 VN.n36 VN.n35 17.9525
R43 VN.n28 VN.n27 12.2198
R44 VN.n5 VN.n4 12.2198
R45 VN.n6 VN.t4 9.89418
R46 VN.n13 VN.t7 9.89418
R47 VN.n21 VN.t0 9.89418
R48 VN.n29 VN.t3 9.89418
R49 VN.n36 VN.t6 9.89418
R50 VN.n44 VN.t2 9.89418
R51 VN.n14 VN.n13 6.6403
R52 VN.n37 VN.n36 6.6403
R53 VN.n21 VN.n20 4.67295
R54 VN.n44 VN.n43 4.67295
R55 VN.n45 VN.n23 0.189894
R56 VN.n41 VN.n23 0.189894
R57 VN.n41 VN.n40 0.189894
R58 VN.n40 VN.n39 0.189894
R59 VN.n39 VN.n25 0.189894
R60 VN.n34 VN.n25 0.189894
R61 VN.n34 VN.n33 0.189894
R62 VN.n33 VN.n32 0.189894
R63 VN.n32 VN.n27 0.189894
R64 VN.n9 VN.n4 0.189894
R65 VN.n10 VN.n9 0.189894
R66 VN.n11 VN.n10 0.189894
R67 VN.n11 VN.n2 0.189894
R68 VN.n16 VN.n2 0.189894
R69 VN.n17 VN.n16 0.189894
R70 VN.n18 VN.n17 0.189894
R71 VN.n18 VN.n0 0.189894
R72 VN.n22 VN.n0 0.189894
R73 VN VN.n22 0.0516364
R74 VTAIL.n15 VTAIL.t13 246.06
R75 VTAIL.n2 VTAIL.t10 246.06
R76 VTAIL.n3 VTAIL.t6 246.06
R77 VTAIL.n6 VTAIL.t7 246.06
R78 VTAIL.n14 VTAIL.t5 246.06
R79 VTAIL.n11 VTAIL.t2 246.06
R80 VTAIL.n10 VTAIL.t9 246.06
R81 VTAIL.n7 VTAIL.t11 246.06
R82 VTAIL.n1 VTAIL.n0 220.677
R83 VTAIL.n5 VTAIL.n4 220.677
R84 VTAIL.n13 VTAIL.n12 220.677
R85 VTAIL.n9 VTAIL.n8 220.677
R86 VTAIL.n0 VTAIL.t8 25.3851
R87 VTAIL.n0 VTAIL.t12 25.3851
R88 VTAIL.n4 VTAIL.t4 25.3851
R89 VTAIL.n4 VTAIL.t0 25.3851
R90 VTAIL.n12 VTAIL.t3 25.3851
R91 VTAIL.n12 VTAIL.t1 25.3851
R92 VTAIL.n8 VTAIL.t14 25.3851
R93 VTAIL.n8 VTAIL.t15 25.3851
R94 VTAIL.n15 VTAIL.n14 14.9617
R95 VTAIL.n7 VTAIL.n6 14.9617
R96 VTAIL.n9 VTAIL.n7 1.92291
R97 VTAIL.n10 VTAIL.n9 1.92291
R98 VTAIL.n13 VTAIL.n11 1.92291
R99 VTAIL.n14 VTAIL.n13 1.92291
R100 VTAIL.n6 VTAIL.n5 1.92291
R101 VTAIL.n5 VTAIL.n3 1.92291
R102 VTAIL.n2 VTAIL.n1 1.92291
R103 VTAIL VTAIL.n15 1.86472
R104 VTAIL.n11 VTAIL.n10 0.470328
R105 VTAIL.n3 VTAIL.n2 0.470328
R106 VTAIL VTAIL.n1 0.0586897
R107 VDD2.n2 VDD2.n1 238.261
R108 VDD2.n2 VDD2.n0 238.261
R109 VDD2 VDD2.n5 238.258
R110 VDD2.n4 VDD2.n3 237.356
R111 VDD2.n4 VDD2.n2 33.0386
R112 VDD2.n5 VDD2.t4 25.3851
R113 VDD2.n5 VDD2.t2 25.3851
R114 VDD2.n3 VDD2.t5 25.3851
R115 VDD2.n3 VDD2.t1 25.3851
R116 VDD2.n1 VDD2.t0 25.3851
R117 VDD2.n1 VDD2.t7 25.3851
R118 VDD2.n0 VDD2.t6 25.3851
R119 VDD2.n0 VDD2.t3 25.3851
R120 VDD2 VDD2.n4 1.0199
R121 B.n476 B.n475 585
R122 B.n477 B.n476 585
R123 B.n147 B.n90 585
R124 B.n146 B.n145 585
R125 B.n144 B.n143 585
R126 B.n142 B.n141 585
R127 B.n140 B.n139 585
R128 B.n138 B.n137 585
R129 B.n136 B.n135 585
R130 B.n134 B.n133 585
R131 B.n132 B.n131 585
R132 B.n130 B.n129 585
R133 B.n128 B.n127 585
R134 B.n126 B.n125 585
R135 B.n124 B.n123 585
R136 B.n122 B.n121 585
R137 B.n120 B.n119 585
R138 B.n118 B.n117 585
R139 B.n116 B.n115 585
R140 B.n113 B.n112 585
R141 B.n111 B.n110 585
R142 B.n109 B.n108 585
R143 B.n107 B.n106 585
R144 B.n105 B.n104 585
R145 B.n103 B.n102 585
R146 B.n101 B.n100 585
R147 B.n99 B.n98 585
R148 B.n97 B.n96 585
R149 B.n474 B.n76 585
R150 B.n478 B.n76 585
R151 B.n473 B.n75 585
R152 B.n479 B.n75 585
R153 B.n472 B.n471 585
R154 B.n471 B.n71 585
R155 B.n470 B.n70 585
R156 B.n485 B.n70 585
R157 B.n469 B.n69 585
R158 B.n486 B.n69 585
R159 B.n468 B.n68 585
R160 B.n487 B.n68 585
R161 B.n467 B.n466 585
R162 B.n466 B.n67 585
R163 B.n465 B.n63 585
R164 B.n493 B.n63 585
R165 B.n464 B.n62 585
R166 B.n494 B.n62 585
R167 B.n463 B.n61 585
R168 B.n495 B.n61 585
R169 B.n462 B.n461 585
R170 B.n461 B.n57 585
R171 B.n460 B.n56 585
R172 B.n501 B.n56 585
R173 B.n459 B.n55 585
R174 B.n502 B.n55 585
R175 B.n458 B.n54 585
R176 B.n503 B.n54 585
R177 B.n457 B.n456 585
R178 B.n456 B.n50 585
R179 B.n455 B.n49 585
R180 B.n509 B.n49 585
R181 B.n454 B.n48 585
R182 B.n510 B.n48 585
R183 B.n453 B.n47 585
R184 B.n511 B.n47 585
R185 B.n452 B.n451 585
R186 B.n451 B.n43 585
R187 B.n450 B.n42 585
R188 B.n517 B.n42 585
R189 B.n449 B.n41 585
R190 B.n518 B.n41 585
R191 B.n448 B.n40 585
R192 B.n519 B.n40 585
R193 B.n447 B.n446 585
R194 B.n446 B.n36 585
R195 B.n445 B.n35 585
R196 B.t1 B.n35 585
R197 B.n444 B.n34 585
R198 B.n525 B.n34 585
R199 B.n443 B.n33 585
R200 B.n526 B.n33 585
R201 B.n442 B.n441 585
R202 B.n441 B.n29 585
R203 B.n440 B.n28 585
R204 B.n532 B.n28 585
R205 B.n439 B.n27 585
R206 B.n533 B.n27 585
R207 B.n438 B.n26 585
R208 B.n534 B.n26 585
R209 B.n437 B.n436 585
R210 B.n436 B.n22 585
R211 B.n435 B.n21 585
R212 B.n540 B.n21 585
R213 B.n434 B.n20 585
R214 B.n541 B.n20 585
R215 B.n433 B.n19 585
R216 B.n542 B.n19 585
R217 B.n432 B.n431 585
R218 B.n431 B.n15 585
R219 B.n430 B.n14 585
R220 B.n548 B.n14 585
R221 B.n429 B.n13 585
R222 B.n549 B.n13 585
R223 B.n428 B.n12 585
R224 B.n550 B.n12 585
R225 B.n427 B.n426 585
R226 B.n426 B.n8 585
R227 B.n425 B.n7 585
R228 B.n556 B.n7 585
R229 B.n424 B.n6 585
R230 B.n557 B.n6 585
R231 B.n423 B.n5 585
R232 B.n558 B.n5 585
R233 B.n422 B.n421 585
R234 B.n421 B.n4 585
R235 B.n420 B.n148 585
R236 B.n420 B.n419 585
R237 B.n410 B.n149 585
R238 B.n150 B.n149 585
R239 B.n412 B.n411 585
R240 B.n413 B.n412 585
R241 B.n409 B.n154 585
R242 B.n158 B.n154 585
R243 B.n408 B.n407 585
R244 B.n407 B.n406 585
R245 B.n156 B.n155 585
R246 B.n157 B.n156 585
R247 B.n399 B.n398 585
R248 B.n400 B.n399 585
R249 B.n397 B.n163 585
R250 B.n163 B.n162 585
R251 B.n396 B.n395 585
R252 B.n395 B.n394 585
R253 B.n165 B.n164 585
R254 B.n166 B.n165 585
R255 B.n387 B.n386 585
R256 B.n388 B.n387 585
R257 B.n385 B.n171 585
R258 B.n171 B.n170 585
R259 B.n384 B.n383 585
R260 B.n383 B.n382 585
R261 B.n173 B.n172 585
R262 B.n174 B.n173 585
R263 B.n375 B.n374 585
R264 B.n376 B.n375 585
R265 B.n373 B.n179 585
R266 B.n179 B.n178 585
R267 B.n372 B.n371 585
R268 B.n371 B.t4 585
R269 B.n181 B.n180 585
R270 B.n182 B.n181 585
R271 B.n364 B.n363 585
R272 B.n365 B.n364 585
R273 B.n362 B.n187 585
R274 B.n187 B.n186 585
R275 B.n361 B.n360 585
R276 B.n360 B.n359 585
R277 B.n189 B.n188 585
R278 B.n190 B.n189 585
R279 B.n352 B.n351 585
R280 B.n353 B.n352 585
R281 B.n350 B.n194 585
R282 B.n198 B.n194 585
R283 B.n349 B.n348 585
R284 B.n348 B.n347 585
R285 B.n196 B.n195 585
R286 B.n197 B.n196 585
R287 B.n340 B.n339 585
R288 B.n341 B.n340 585
R289 B.n338 B.n203 585
R290 B.n203 B.n202 585
R291 B.n337 B.n336 585
R292 B.n336 B.n335 585
R293 B.n205 B.n204 585
R294 B.n206 B.n205 585
R295 B.n328 B.n327 585
R296 B.n329 B.n328 585
R297 B.n326 B.n211 585
R298 B.n211 B.n210 585
R299 B.n325 B.n324 585
R300 B.n324 B.n323 585
R301 B.n213 B.n212 585
R302 B.n316 B.n213 585
R303 B.n315 B.n314 585
R304 B.n317 B.n315 585
R305 B.n313 B.n218 585
R306 B.n218 B.n217 585
R307 B.n312 B.n311 585
R308 B.n311 B.n310 585
R309 B.n220 B.n219 585
R310 B.n221 B.n220 585
R311 B.n303 B.n302 585
R312 B.n304 B.n303 585
R313 B.n301 B.n226 585
R314 B.n226 B.n225 585
R315 B.n295 B.n294 585
R316 B.n293 B.n241 585
R317 B.n292 B.n240 585
R318 B.n297 B.n240 585
R319 B.n291 B.n290 585
R320 B.n289 B.n288 585
R321 B.n287 B.n286 585
R322 B.n285 B.n284 585
R323 B.n283 B.n282 585
R324 B.n281 B.n280 585
R325 B.n279 B.n278 585
R326 B.n277 B.n276 585
R327 B.n275 B.n274 585
R328 B.n273 B.n272 585
R329 B.n271 B.n270 585
R330 B.n269 B.n268 585
R331 B.n267 B.n266 585
R332 B.n265 B.n264 585
R333 B.n263 B.n262 585
R334 B.n260 B.n259 585
R335 B.n258 B.n257 585
R336 B.n256 B.n255 585
R337 B.n254 B.n253 585
R338 B.n252 B.n251 585
R339 B.n250 B.n249 585
R340 B.n248 B.n247 585
R341 B.n228 B.n227 585
R342 B.n300 B.n299 585
R343 B.n224 B.n223 585
R344 B.n225 B.n224 585
R345 B.n306 B.n305 585
R346 B.n305 B.n304 585
R347 B.n307 B.n222 585
R348 B.n222 B.n221 585
R349 B.n309 B.n308 585
R350 B.n310 B.n309 585
R351 B.n216 B.n215 585
R352 B.n217 B.n216 585
R353 B.n319 B.n318 585
R354 B.n318 B.n317 585
R355 B.n320 B.n214 585
R356 B.n316 B.n214 585
R357 B.n322 B.n321 585
R358 B.n323 B.n322 585
R359 B.n209 B.n208 585
R360 B.n210 B.n209 585
R361 B.n331 B.n330 585
R362 B.n330 B.n329 585
R363 B.n332 B.n207 585
R364 B.n207 B.n206 585
R365 B.n334 B.n333 585
R366 B.n335 B.n334 585
R367 B.n201 B.n200 585
R368 B.n202 B.n201 585
R369 B.n343 B.n342 585
R370 B.n342 B.n341 585
R371 B.n344 B.n199 585
R372 B.n199 B.n197 585
R373 B.n346 B.n345 585
R374 B.n347 B.n346 585
R375 B.n193 B.n192 585
R376 B.n198 B.n193 585
R377 B.n355 B.n354 585
R378 B.n354 B.n353 585
R379 B.n356 B.n191 585
R380 B.n191 B.n190 585
R381 B.n358 B.n357 585
R382 B.n359 B.n358 585
R383 B.n185 B.n184 585
R384 B.n186 B.n185 585
R385 B.n367 B.n366 585
R386 B.n366 B.n365 585
R387 B.n368 B.n183 585
R388 B.n183 B.n182 585
R389 B.n370 B.n369 585
R390 B.t4 B.n370 585
R391 B.n177 B.n176 585
R392 B.n178 B.n177 585
R393 B.n378 B.n377 585
R394 B.n377 B.n376 585
R395 B.n379 B.n175 585
R396 B.n175 B.n174 585
R397 B.n381 B.n380 585
R398 B.n382 B.n381 585
R399 B.n169 B.n168 585
R400 B.n170 B.n169 585
R401 B.n390 B.n389 585
R402 B.n389 B.n388 585
R403 B.n391 B.n167 585
R404 B.n167 B.n166 585
R405 B.n393 B.n392 585
R406 B.n394 B.n393 585
R407 B.n161 B.n160 585
R408 B.n162 B.n161 585
R409 B.n402 B.n401 585
R410 B.n401 B.n400 585
R411 B.n403 B.n159 585
R412 B.n159 B.n157 585
R413 B.n405 B.n404 585
R414 B.n406 B.n405 585
R415 B.n153 B.n152 585
R416 B.n158 B.n153 585
R417 B.n415 B.n414 585
R418 B.n414 B.n413 585
R419 B.n416 B.n151 585
R420 B.n151 B.n150 585
R421 B.n418 B.n417 585
R422 B.n419 B.n418 585
R423 B.n2 B.n0 585
R424 B.n4 B.n2 585
R425 B.n3 B.n1 585
R426 B.n557 B.n3 585
R427 B.n555 B.n554 585
R428 B.n556 B.n555 585
R429 B.n553 B.n9 585
R430 B.n9 B.n8 585
R431 B.n552 B.n551 585
R432 B.n551 B.n550 585
R433 B.n11 B.n10 585
R434 B.n549 B.n11 585
R435 B.n547 B.n546 585
R436 B.n548 B.n547 585
R437 B.n545 B.n16 585
R438 B.n16 B.n15 585
R439 B.n544 B.n543 585
R440 B.n543 B.n542 585
R441 B.n18 B.n17 585
R442 B.n541 B.n18 585
R443 B.n539 B.n538 585
R444 B.n540 B.n539 585
R445 B.n537 B.n23 585
R446 B.n23 B.n22 585
R447 B.n536 B.n535 585
R448 B.n535 B.n534 585
R449 B.n25 B.n24 585
R450 B.n533 B.n25 585
R451 B.n531 B.n530 585
R452 B.n532 B.n531 585
R453 B.n529 B.n30 585
R454 B.n30 B.n29 585
R455 B.n528 B.n527 585
R456 B.n527 B.n526 585
R457 B.n32 B.n31 585
R458 B.n525 B.n32 585
R459 B.n524 B.n523 585
R460 B.t1 B.n524 585
R461 B.n522 B.n37 585
R462 B.n37 B.n36 585
R463 B.n521 B.n520 585
R464 B.n520 B.n519 585
R465 B.n39 B.n38 585
R466 B.n518 B.n39 585
R467 B.n516 B.n515 585
R468 B.n517 B.n516 585
R469 B.n514 B.n44 585
R470 B.n44 B.n43 585
R471 B.n513 B.n512 585
R472 B.n512 B.n511 585
R473 B.n46 B.n45 585
R474 B.n510 B.n46 585
R475 B.n508 B.n507 585
R476 B.n509 B.n508 585
R477 B.n506 B.n51 585
R478 B.n51 B.n50 585
R479 B.n505 B.n504 585
R480 B.n504 B.n503 585
R481 B.n53 B.n52 585
R482 B.n502 B.n53 585
R483 B.n500 B.n499 585
R484 B.n501 B.n500 585
R485 B.n498 B.n58 585
R486 B.n58 B.n57 585
R487 B.n497 B.n496 585
R488 B.n496 B.n495 585
R489 B.n60 B.n59 585
R490 B.n494 B.n60 585
R491 B.n492 B.n491 585
R492 B.n493 B.n492 585
R493 B.n490 B.n64 585
R494 B.n67 B.n64 585
R495 B.n489 B.n488 585
R496 B.n488 B.n487 585
R497 B.n66 B.n65 585
R498 B.n486 B.n66 585
R499 B.n484 B.n483 585
R500 B.n485 B.n484 585
R501 B.n482 B.n72 585
R502 B.n72 B.n71 585
R503 B.n481 B.n480 585
R504 B.n480 B.n479 585
R505 B.n74 B.n73 585
R506 B.n478 B.n74 585
R507 B.n560 B.n559 585
R508 B.n559 B.n558 585
R509 B.n295 B.n224 468.476
R510 B.n96 B.n74 468.476
R511 B.n299 B.n226 468.476
R512 B.n476 B.n76 468.476
R513 B.n245 B.t18 278.457
R514 B.n242 B.t15 278.457
R515 B.n94 B.t10 278.457
R516 B.n91 B.t20 278.457
R517 B.n477 B.n89 256.663
R518 B.n477 B.n88 256.663
R519 B.n477 B.n87 256.663
R520 B.n477 B.n86 256.663
R521 B.n477 B.n85 256.663
R522 B.n477 B.n84 256.663
R523 B.n477 B.n83 256.663
R524 B.n477 B.n82 256.663
R525 B.n477 B.n81 256.663
R526 B.n477 B.n80 256.663
R527 B.n477 B.n79 256.663
R528 B.n477 B.n78 256.663
R529 B.n477 B.n77 256.663
R530 B.n297 B.n296 256.663
R531 B.n297 B.n229 256.663
R532 B.n297 B.n230 256.663
R533 B.n297 B.n231 256.663
R534 B.n297 B.n232 256.663
R535 B.n297 B.n233 256.663
R536 B.n297 B.n234 256.663
R537 B.n297 B.n235 256.663
R538 B.n297 B.n236 256.663
R539 B.n297 B.n237 256.663
R540 B.n297 B.n238 256.663
R541 B.n297 B.n239 256.663
R542 B.n298 B.n297 256.663
R543 B.n246 B.t17 235.209
R544 B.n243 B.t14 235.209
R545 B.n95 B.t11 235.209
R546 B.n92 B.t21 235.209
R547 B.n297 B.n225 212.553
R548 B.n478 B.n477 212.553
R549 B.n245 B.t16 208.07
R550 B.n242 B.t12 208.07
R551 B.n94 B.t8 208.07
R552 B.n91 B.t19 208.07
R553 B.n305 B.n224 163.367
R554 B.n305 B.n222 163.367
R555 B.n309 B.n222 163.367
R556 B.n309 B.n216 163.367
R557 B.n318 B.n216 163.367
R558 B.n318 B.n214 163.367
R559 B.n322 B.n214 163.367
R560 B.n322 B.n209 163.367
R561 B.n330 B.n209 163.367
R562 B.n330 B.n207 163.367
R563 B.n334 B.n207 163.367
R564 B.n334 B.n201 163.367
R565 B.n342 B.n201 163.367
R566 B.n342 B.n199 163.367
R567 B.n346 B.n199 163.367
R568 B.n346 B.n193 163.367
R569 B.n354 B.n193 163.367
R570 B.n354 B.n191 163.367
R571 B.n358 B.n191 163.367
R572 B.n358 B.n185 163.367
R573 B.n366 B.n185 163.367
R574 B.n366 B.n183 163.367
R575 B.n370 B.n183 163.367
R576 B.n370 B.n177 163.367
R577 B.n377 B.n177 163.367
R578 B.n377 B.n175 163.367
R579 B.n381 B.n175 163.367
R580 B.n381 B.n169 163.367
R581 B.n389 B.n169 163.367
R582 B.n389 B.n167 163.367
R583 B.n393 B.n167 163.367
R584 B.n393 B.n161 163.367
R585 B.n401 B.n161 163.367
R586 B.n401 B.n159 163.367
R587 B.n405 B.n159 163.367
R588 B.n405 B.n153 163.367
R589 B.n414 B.n153 163.367
R590 B.n414 B.n151 163.367
R591 B.n418 B.n151 163.367
R592 B.n418 B.n2 163.367
R593 B.n559 B.n2 163.367
R594 B.n559 B.n3 163.367
R595 B.n555 B.n3 163.367
R596 B.n555 B.n9 163.367
R597 B.n551 B.n9 163.367
R598 B.n551 B.n11 163.367
R599 B.n547 B.n11 163.367
R600 B.n547 B.n16 163.367
R601 B.n543 B.n16 163.367
R602 B.n543 B.n18 163.367
R603 B.n539 B.n18 163.367
R604 B.n539 B.n23 163.367
R605 B.n535 B.n23 163.367
R606 B.n535 B.n25 163.367
R607 B.n531 B.n25 163.367
R608 B.n531 B.n30 163.367
R609 B.n527 B.n30 163.367
R610 B.n527 B.n32 163.367
R611 B.n524 B.n32 163.367
R612 B.n524 B.n37 163.367
R613 B.n520 B.n37 163.367
R614 B.n520 B.n39 163.367
R615 B.n516 B.n39 163.367
R616 B.n516 B.n44 163.367
R617 B.n512 B.n44 163.367
R618 B.n512 B.n46 163.367
R619 B.n508 B.n46 163.367
R620 B.n508 B.n51 163.367
R621 B.n504 B.n51 163.367
R622 B.n504 B.n53 163.367
R623 B.n500 B.n53 163.367
R624 B.n500 B.n58 163.367
R625 B.n496 B.n58 163.367
R626 B.n496 B.n60 163.367
R627 B.n492 B.n60 163.367
R628 B.n492 B.n64 163.367
R629 B.n488 B.n64 163.367
R630 B.n488 B.n66 163.367
R631 B.n484 B.n66 163.367
R632 B.n484 B.n72 163.367
R633 B.n480 B.n72 163.367
R634 B.n480 B.n74 163.367
R635 B.n241 B.n240 163.367
R636 B.n290 B.n240 163.367
R637 B.n288 B.n287 163.367
R638 B.n284 B.n283 163.367
R639 B.n280 B.n279 163.367
R640 B.n276 B.n275 163.367
R641 B.n272 B.n271 163.367
R642 B.n268 B.n267 163.367
R643 B.n264 B.n263 163.367
R644 B.n259 B.n258 163.367
R645 B.n255 B.n254 163.367
R646 B.n251 B.n250 163.367
R647 B.n247 B.n228 163.367
R648 B.n303 B.n226 163.367
R649 B.n303 B.n220 163.367
R650 B.n311 B.n220 163.367
R651 B.n311 B.n218 163.367
R652 B.n315 B.n218 163.367
R653 B.n315 B.n213 163.367
R654 B.n324 B.n213 163.367
R655 B.n324 B.n211 163.367
R656 B.n328 B.n211 163.367
R657 B.n328 B.n205 163.367
R658 B.n336 B.n205 163.367
R659 B.n336 B.n203 163.367
R660 B.n340 B.n203 163.367
R661 B.n340 B.n196 163.367
R662 B.n348 B.n196 163.367
R663 B.n348 B.n194 163.367
R664 B.n352 B.n194 163.367
R665 B.n352 B.n189 163.367
R666 B.n360 B.n189 163.367
R667 B.n360 B.n187 163.367
R668 B.n364 B.n187 163.367
R669 B.n364 B.n181 163.367
R670 B.n371 B.n181 163.367
R671 B.n371 B.n179 163.367
R672 B.n375 B.n179 163.367
R673 B.n375 B.n173 163.367
R674 B.n383 B.n173 163.367
R675 B.n383 B.n171 163.367
R676 B.n387 B.n171 163.367
R677 B.n387 B.n165 163.367
R678 B.n395 B.n165 163.367
R679 B.n395 B.n163 163.367
R680 B.n399 B.n163 163.367
R681 B.n399 B.n156 163.367
R682 B.n407 B.n156 163.367
R683 B.n407 B.n154 163.367
R684 B.n412 B.n154 163.367
R685 B.n412 B.n149 163.367
R686 B.n420 B.n149 163.367
R687 B.n421 B.n420 163.367
R688 B.n421 B.n5 163.367
R689 B.n6 B.n5 163.367
R690 B.n7 B.n6 163.367
R691 B.n426 B.n7 163.367
R692 B.n426 B.n12 163.367
R693 B.n13 B.n12 163.367
R694 B.n14 B.n13 163.367
R695 B.n431 B.n14 163.367
R696 B.n431 B.n19 163.367
R697 B.n20 B.n19 163.367
R698 B.n21 B.n20 163.367
R699 B.n436 B.n21 163.367
R700 B.n436 B.n26 163.367
R701 B.n27 B.n26 163.367
R702 B.n28 B.n27 163.367
R703 B.n441 B.n28 163.367
R704 B.n441 B.n33 163.367
R705 B.n34 B.n33 163.367
R706 B.n35 B.n34 163.367
R707 B.n446 B.n35 163.367
R708 B.n446 B.n40 163.367
R709 B.n41 B.n40 163.367
R710 B.n42 B.n41 163.367
R711 B.n451 B.n42 163.367
R712 B.n451 B.n47 163.367
R713 B.n48 B.n47 163.367
R714 B.n49 B.n48 163.367
R715 B.n456 B.n49 163.367
R716 B.n456 B.n54 163.367
R717 B.n55 B.n54 163.367
R718 B.n56 B.n55 163.367
R719 B.n461 B.n56 163.367
R720 B.n461 B.n61 163.367
R721 B.n62 B.n61 163.367
R722 B.n63 B.n62 163.367
R723 B.n466 B.n63 163.367
R724 B.n466 B.n68 163.367
R725 B.n69 B.n68 163.367
R726 B.n70 B.n69 163.367
R727 B.n471 B.n70 163.367
R728 B.n471 B.n75 163.367
R729 B.n76 B.n75 163.367
R730 B.n100 B.n99 163.367
R731 B.n104 B.n103 163.367
R732 B.n108 B.n107 163.367
R733 B.n112 B.n111 163.367
R734 B.n117 B.n116 163.367
R735 B.n121 B.n120 163.367
R736 B.n125 B.n124 163.367
R737 B.n129 B.n128 163.367
R738 B.n133 B.n132 163.367
R739 B.n137 B.n136 163.367
R740 B.n141 B.n140 163.367
R741 B.n145 B.n144 163.367
R742 B.n476 B.n90 163.367
R743 B.n304 B.n225 123.534
R744 B.n304 B.n221 123.534
R745 B.n310 B.n221 123.534
R746 B.n310 B.n217 123.534
R747 B.n317 B.n217 123.534
R748 B.n317 B.n316 123.534
R749 B.n323 B.n210 123.534
R750 B.n329 B.n210 123.534
R751 B.n329 B.n206 123.534
R752 B.n335 B.n206 123.534
R753 B.n335 B.n202 123.534
R754 B.n341 B.n202 123.534
R755 B.n341 B.n197 123.534
R756 B.n347 B.n197 123.534
R757 B.n347 B.n198 123.534
R758 B.n353 B.n190 123.534
R759 B.n359 B.n190 123.534
R760 B.n359 B.n186 123.534
R761 B.n365 B.n186 123.534
R762 B.n365 B.n182 123.534
R763 B.t4 B.n182 123.534
R764 B.t4 B.n178 123.534
R765 B.n376 B.n178 123.534
R766 B.n376 B.n174 123.534
R767 B.n382 B.n174 123.534
R768 B.n382 B.n170 123.534
R769 B.n388 B.n170 123.534
R770 B.n394 B.n166 123.534
R771 B.n394 B.n162 123.534
R772 B.n400 B.n162 123.534
R773 B.n400 B.n157 123.534
R774 B.n406 B.n157 123.534
R775 B.n406 B.n158 123.534
R776 B.n413 B.n150 123.534
R777 B.n419 B.n150 123.534
R778 B.n419 B.n4 123.534
R779 B.n558 B.n4 123.534
R780 B.n558 B.n557 123.534
R781 B.n557 B.n556 123.534
R782 B.n556 B.n8 123.534
R783 B.n550 B.n8 123.534
R784 B.n549 B.n548 123.534
R785 B.n548 B.n15 123.534
R786 B.n542 B.n15 123.534
R787 B.n542 B.n541 123.534
R788 B.n541 B.n540 123.534
R789 B.n540 B.n22 123.534
R790 B.n534 B.n533 123.534
R791 B.n533 B.n532 123.534
R792 B.n532 B.n29 123.534
R793 B.n526 B.n29 123.534
R794 B.n526 B.n525 123.534
R795 B.n525 B.t1 123.534
R796 B.t1 B.n36 123.534
R797 B.n519 B.n36 123.534
R798 B.n519 B.n518 123.534
R799 B.n518 B.n517 123.534
R800 B.n517 B.n43 123.534
R801 B.n511 B.n43 123.534
R802 B.n510 B.n509 123.534
R803 B.n509 B.n50 123.534
R804 B.n503 B.n50 123.534
R805 B.n503 B.n502 123.534
R806 B.n502 B.n501 123.534
R807 B.n501 B.n57 123.534
R808 B.n495 B.n57 123.534
R809 B.n495 B.n494 123.534
R810 B.n494 B.n493 123.534
R811 B.n487 B.n67 123.534
R812 B.n487 B.n486 123.534
R813 B.n486 B.n485 123.534
R814 B.n485 B.n71 123.534
R815 B.n479 B.n71 123.534
R816 B.n479 B.n478 123.534
R817 B.n413 B.t6 109.001
R818 B.n550 B.t2 109.001
R819 B.n316 B.t13 83.5678
R820 B.n67 B.t9 83.5678
R821 B.n296 B.n295 71.676
R822 B.n290 B.n229 71.676
R823 B.n287 B.n230 71.676
R824 B.n283 B.n231 71.676
R825 B.n279 B.n232 71.676
R826 B.n275 B.n233 71.676
R827 B.n271 B.n234 71.676
R828 B.n267 B.n235 71.676
R829 B.n263 B.n236 71.676
R830 B.n258 B.n237 71.676
R831 B.n254 B.n238 71.676
R832 B.n250 B.n239 71.676
R833 B.n298 B.n228 71.676
R834 B.n96 B.n77 71.676
R835 B.n100 B.n78 71.676
R836 B.n104 B.n79 71.676
R837 B.n108 B.n80 71.676
R838 B.n112 B.n81 71.676
R839 B.n117 B.n82 71.676
R840 B.n121 B.n83 71.676
R841 B.n125 B.n84 71.676
R842 B.n129 B.n85 71.676
R843 B.n133 B.n86 71.676
R844 B.n137 B.n87 71.676
R845 B.n141 B.n88 71.676
R846 B.n145 B.n89 71.676
R847 B.n90 B.n89 71.676
R848 B.n144 B.n88 71.676
R849 B.n140 B.n87 71.676
R850 B.n136 B.n86 71.676
R851 B.n132 B.n85 71.676
R852 B.n128 B.n84 71.676
R853 B.n124 B.n83 71.676
R854 B.n120 B.n82 71.676
R855 B.n116 B.n81 71.676
R856 B.n111 B.n80 71.676
R857 B.n107 B.n79 71.676
R858 B.n103 B.n78 71.676
R859 B.n99 B.n77 71.676
R860 B.n296 B.n241 71.676
R861 B.n288 B.n229 71.676
R862 B.n284 B.n230 71.676
R863 B.n280 B.n231 71.676
R864 B.n276 B.n232 71.676
R865 B.n272 B.n233 71.676
R866 B.n268 B.n234 71.676
R867 B.n264 B.n235 71.676
R868 B.n259 B.n236 71.676
R869 B.n255 B.n237 71.676
R870 B.n251 B.n238 71.676
R871 B.n247 B.n239 71.676
R872 B.n299 B.n298 71.676
R873 B.n353 B.t7 69.0344
R874 B.n388 B.t0 69.0344
R875 B.n534 B.t3 69.0344
R876 B.n511 B.t5 69.0344
R877 B.n261 B.n246 59.5399
R878 B.n244 B.n243 59.5399
R879 B.n114 B.n95 59.5399
R880 B.n93 B.n92 59.5399
R881 B.n198 B.t7 54.5009
R882 B.t0 B.n166 54.5009
R883 B.t3 B.n22 54.5009
R884 B.t5 B.n510 54.5009
R885 B.n246 B.n245 43.249
R886 B.n243 B.n242 43.249
R887 B.n95 B.n94 43.249
R888 B.n92 B.n91 43.249
R889 B.n323 B.t13 39.9675
R890 B.n493 B.t9 39.9675
R891 B.n97 B.n73 30.4395
R892 B.n475 B.n474 30.4395
R893 B.n301 B.n300 30.4395
R894 B.n294 B.n223 30.4395
R895 B B.n560 18.0485
R896 B.n158 B.t6 14.5339
R897 B.t2 B.n549 14.5339
R898 B.n98 B.n97 10.6151
R899 B.n101 B.n98 10.6151
R900 B.n102 B.n101 10.6151
R901 B.n105 B.n102 10.6151
R902 B.n106 B.n105 10.6151
R903 B.n109 B.n106 10.6151
R904 B.n110 B.n109 10.6151
R905 B.n113 B.n110 10.6151
R906 B.n118 B.n115 10.6151
R907 B.n119 B.n118 10.6151
R908 B.n122 B.n119 10.6151
R909 B.n123 B.n122 10.6151
R910 B.n126 B.n123 10.6151
R911 B.n127 B.n126 10.6151
R912 B.n130 B.n127 10.6151
R913 B.n131 B.n130 10.6151
R914 B.n135 B.n134 10.6151
R915 B.n138 B.n135 10.6151
R916 B.n139 B.n138 10.6151
R917 B.n142 B.n139 10.6151
R918 B.n143 B.n142 10.6151
R919 B.n146 B.n143 10.6151
R920 B.n147 B.n146 10.6151
R921 B.n475 B.n147 10.6151
R922 B.n302 B.n301 10.6151
R923 B.n302 B.n219 10.6151
R924 B.n312 B.n219 10.6151
R925 B.n313 B.n312 10.6151
R926 B.n314 B.n313 10.6151
R927 B.n314 B.n212 10.6151
R928 B.n325 B.n212 10.6151
R929 B.n326 B.n325 10.6151
R930 B.n327 B.n326 10.6151
R931 B.n327 B.n204 10.6151
R932 B.n337 B.n204 10.6151
R933 B.n338 B.n337 10.6151
R934 B.n339 B.n338 10.6151
R935 B.n339 B.n195 10.6151
R936 B.n349 B.n195 10.6151
R937 B.n350 B.n349 10.6151
R938 B.n351 B.n350 10.6151
R939 B.n351 B.n188 10.6151
R940 B.n361 B.n188 10.6151
R941 B.n362 B.n361 10.6151
R942 B.n363 B.n362 10.6151
R943 B.n363 B.n180 10.6151
R944 B.n372 B.n180 10.6151
R945 B.n373 B.n372 10.6151
R946 B.n374 B.n373 10.6151
R947 B.n374 B.n172 10.6151
R948 B.n384 B.n172 10.6151
R949 B.n385 B.n384 10.6151
R950 B.n386 B.n385 10.6151
R951 B.n386 B.n164 10.6151
R952 B.n396 B.n164 10.6151
R953 B.n397 B.n396 10.6151
R954 B.n398 B.n397 10.6151
R955 B.n398 B.n155 10.6151
R956 B.n408 B.n155 10.6151
R957 B.n409 B.n408 10.6151
R958 B.n411 B.n409 10.6151
R959 B.n411 B.n410 10.6151
R960 B.n410 B.n148 10.6151
R961 B.n422 B.n148 10.6151
R962 B.n423 B.n422 10.6151
R963 B.n424 B.n423 10.6151
R964 B.n425 B.n424 10.6151
R965 B.n427 B.n425 10.6151
R966 B.n428 B.n427 10.6151
R967 B.n429 B.n428 10.6151
R968 B.n430 B.n429 10.6151
R969 B.n432 B.n430 10.6151
R970 B.n433 B.n432 10.6151
R971 B.n434 B.n433 10.6151
R972 B.n435 B.n434 10.6151
R973 B.n437 B.n435 10.6151
R974 B.n438 B.n437 10.6151
R975 B.n439 B.n438 10.6151
R976 B.n440 B.n439 10.6151
R977 B.n442 B.n440 10.6151
R978 B.n443 B.n442 10.6151
R979 B.n444 B.n443 10.6151
R980 B.n445 B.n444 10.6151
R981 B.n447 B.n445 10.6151
R982 B.n448 B.n447 10.6151
R983 B.n449 B.n448 10.6151
R984 B.n450 B.n449 10.6151
R985 B.n452 B.n450 10.6151
R986 B.n453 B.n452 10.6151
R987 B.n454 B.n453 10.6151
R988 B.n455 B.n454 10.6151
R989 B.n457 B.n455 10.6151
R990 B.n458 B.n457 10.6151
R991 B.n459 B.n458 10.6151
R992 B.n460 B.n459 10.6151
R993 B.n462 B.n460 10.6151
R994 B.n463 B.n462 10.6151
R995 B.n464 B.n463 10.6151
R996 B.n465 B.n464 10.6151
R997 B.n467 B.n465 10.6151
R998 B.n468 B.n467 10.6151
R999 B.n469 B.n468 10.6151
R1000 B.n470 B.n469 10.6151
R1001 B.n472 B.n470 10.6151
R1002 B.n473 B.n472 10.6151
R1003 B.n474 B.n473 10.6151
R1004 B.n294 B.n293 10.6151
R1005 B.n293 B.n292 10.6151
R1006 B.n292 B.n291 10.6151
R1007 B.n291 B.n289 10.6151
R1008 B.n289 B.n286 10.6151
R1009 B.n286 B.n285 10.6151
R1010 B.n285 B.n282 10.6151
R1011 B.n282 B.n281 10.6151
R1012 B.n278 B.n277 10.6151
R1013 B.n277 B.n274 10.6151
R1014 B.n274 B.n273 10.6151
R1015 B.n273 B.n270 10.6151
R1016 B.n270 B.n269 10.6151
R1017 B.n269 B.n266 10.6151
R1018 B.n266 B.n265 10.6151
R1019 B.n265 B.n262 10.6151
R1020 B.n260 B.n257 10.6151
R1021 B.n257 B.n256 10.6151
R1022 B.n256 B.n253 10.6151
R1023 B.n253 B.n252 10.6151
R1024 B.n252 B.n249 10.6151
R1025 B.n249 B.n248 10.6151
R1026 B.n248 B.n227 10.6151
R1027 B.n300 B.n227 10.6151
R1028 B.n306 B.n223 10.6151
R1029 B.n307 B.n306 10.6151
R1030 B.n308 B.n307 10.6151
R1031 B.n308 B.n215 10.6151
R1032 B.n319 B.n215 10.6151
R1033 B.n320 B.n319 10.6151
R1034 B.n321 B.n320 10.6151
R1035 B.n321 B.n208 10.6151
R1036 B.n331 B.n208 10.6151
R1037 B.n332 B.n331 10.6151
R1038 B.n333 B.n332 10.6151
R1039 B.n333 B.n200 10.6151
R1040 B.n343 B.n200 10.6151
R1041 B.n344 B.n343 10.6151
R1042 B.n345 B.n344 10.6151
R1043 B.n345 B.n192 10.6151
R1044 B.n355 B.n192 10.6151
R1045 B.n356 B.n355 10.6151
R1046 B.n357 B.n356 10.6151
R1047 B.n357 B.n184 10.6151
R1048 B.n367 B.n184 10.6151
R1049 B.n368 B.n367 10.6151
R1050 B.n369 B.n368 10.6151
R1051 B.n369 B.n176 10.6151
R1052 B.n378 B.n176 10.6151
R1053 B.n379 B.n378 10.6151
R1054 B.n380 B.n379 10.6151
R1055 B.n380 B.n168 10.6151
R1056 B.n390 B.n168 10.6151
R1057 B.n391 B.n390 10.6151
R1058 B.n392 B.n391 10.6151
R1059 B.n392 B.n160 10.6151
R1060 B.n402 B.n160 10.6151
R1061 B.n403 B.n402 10.6151
R1062 B.n404 B.n403 10.6151
R1063 B.n404 B.n152 10.6151
R1064 B.n415 B.n152 10.6151
R1065 B.n416 B.n415 10.6151
R1066 B.n417 B.n416 10.6151
R1067 B.n417 B.n0 10.6151
R1068 B.n554 B.n1 10.6151
R1069 B.n554 B.n553 10.6151
R1070 B.n553 B.n552 10.6151
R1071 B.n552 B.n10 10.6151
R1072 B.n546 B.n10 10.6151
R1073 B.n546 B.n545 10.6151
R1074 B.n545 B.n544 10.6151
R1075 B.n544 B.n17 10.6151
R1076 B.n538 B.n17 10.6151
R1077 B.n538 B.n537 10.6151
R1078 B.n537 B.n536 10.6151
R1079 B.n536 B.n24 10.6151
R1080 B.n530 B.n24 10.6151
R1081 B.n530 B.n529 10.6151
R1082 B.n529 B.n528 10.6151
R1083 B.n528 B.n31 10.6151
R1084 B.n523 B.n31 10.6151
R1085 B.n523 B.n522 10.6151
R1086 B.n522 B.n521 10.6151
R1087 B.n521 B.n38 10.6151
R1088 B.n515 B.n38 10.6151
R1089 B.n515 B.n514 10.6151
R1090 B.n514 B.n513 10.6151
R1091 B.n513 B.n45 10.6151
R1092 B.n507 B.n45 10.6151
R1093 B.n507 B.n506 10.6151
R1094 B.n506 B.n505 10.6151
R1095 B.n505 B.n52 10.6151
R1096 B.n499 B.n52 10.6151
R1097 B.n499 B.n498 10.6151
R1098 B.n498 B.n497 10.6151
R1099 B.n497 B.n59 10.6151
R1100 B.n491 B.n59 10.6151
R1101 B.n491 B.n490 10.6151
R1102 B.n490 B.n489 10.6151
R1103 B.n489 B.n65 10.6151
R1104 B.n483 B.n65 10.6151
R1105 B.n483 B.n482 10.6151
R1106 B.n482 B.n481 10.6151
R1107 B.n481 B.n73 10.6151
R1108 B.n115 B.n114 6.5566
R1109 B.n131 B.n93 6.5566
R1110 B.n278 B.n244 6.5566
R1111 B.n262 B.n261 6.5566
R1112 B.n114 B.n113 4.05904
R1113 B.n134 B.n93 4.05904
R1114 B.n281 B.n244 4.05904
R1115 B.n261 B.n260 4.05904
R1116 B.n560 B.n0 2.81026
R1117 B.n560 B.n1 2.81026
R1118 VP.n31 VP.n7 181.22
R1119 VP.n56 VP.n55 181.22
R1120 VP.n30 VP.n29 181.22
R1121 VP.n15 VP.n12 161.3
R1122 VP.n17 VP.n16 161.3
R1123 VP.n18 VP.n11 161.3
R1124 VP.n20 VP.n19 161.3
R1125 VP.n22 VP.n10 161.3
R1126 VP.n24 VP.n23 161.3
R1127 VP.n25 VP.n9 161.3
R1128 VP.n27 VP.n26 161.3
R1129 VP.n28 VP.n8 161.3
R1130 VP.n54 VP.n0 161.3
R1131 VP.n53 VP.n52 161.3
R1132 VP.n51 VP.n1 161.3
R1133 VP.n50 VP.n49 161.3
R1134 VP.n48 VP.n2 161.3
R1135 VP.n46 VP.n45 161.3
R1136 VP.n44 VP.n3 161.3
R1137 VP.n43 VP.n42 161.3
R1138 VP.n41 VP.n4 161.3
R1139 VP.n39 VP.n38 161.3
R1140 VP.n37 VP.n5 161.3
R1141 VP.n36 VP.n35 161.3
R1142 VP.n34 VP.n6 161.3
R1143 VP.n33 VP.n32 161.3
R1144 VP.n42 VP.n3 56.5617
R1145 VP.n16 VP.n11 56.5617
R1146 VP.n14 VP.n13 51.8866
R1147 VP.n13 VP.t6 44.7859
R1148 VP.n35 VP.n5 42.5146
R1149 VP.n49 VP.n1 42.5146
R1150 VP.n23 VP.n9 42.5146
R1151 VP.n31 VP.n30 39.0611
R1152 VP.n35 VP.n34 38.6395
R1153 VP.n53 VP.n1 38.6395
R1154 VP.n27 VP.n9 38.6395
R1155 VP.n34 VP.n33 24.5923
R1156 VP.n39 VP.n5 24.5923
R1157 VP.n42 VP.n41 24.5923
R1158 VP.n46 VP.n3 24.5923
R1159 VP.n49 VP.n48 24.5923
R1160 VP.n54 VP.n53 24.5923
R1161 VP.n28 VP.n27 24.5923
R1162 VP.n20 VP.n11 24.5923
R1163 VP.n23 VP.n22 24.5923
R1164 VP.n16 VP.n15 24.5923
R1165 VP.n41 VP.n40 17.9525
R1166 VP.n47 VP.n46 17.9525
R1167 VP.n21 VP.n20 17.9525
R1168 VP.n15 VP.n14 17.9525
R1169 VP.n13 VP.n12 12.2198
R1170 VP.n7 VP.t2 9.89418
R1171 VP.n40 VP.t7 9.89418
R1172 VP.n47 VP.t5 9.89418
R1173 VP.n55 VP.t0 9.89418
R1174 VP.n29 VP.t1 9.89418
R1175 VP.n21 VP.t3 9.89418
R1176 VP.n14 VP.t4 9.89418
R1177 VP.n40 VP.n39 6.6403
R1178 VP.n48 VP.n47 6.6403
R1179 VP.n22 VP.n21 6.6403
R1180 VP.n33 VP.n7 4.67295
R1181 VP.n55 VP.n54 4.67295
R1182 VP.n29 VP.n28 4.67295
R1183 VP.n17 VP.n12 0.189894
R1184 VP.n18 VP.n17 0.189894
R1185 VP.n19 VP.n18 0.189894
R1186 VP.n19 VP.n10 0.189894
R1187 VP.n24 VP.n10 0.189894
R1188 VP.n25 VP.n24 0.189894
R1189 VP.n26 VP.n25 0.189894
R1190 VP.n26 VP.n8 0.189894
R1191 VP.n30 VP.n8 0.189894
R1192 VP.n32 VP.n31 0.189894
R1193 VP.n32 VP.n6 0.189894
R1194 VP.n36 VP.n6 0.189894
R1195 VP.n37 VP.n36 0.189894
R1196 VP.n38 VP.n37 0.189894
R1197 VP.n38 VP.n4 0.189894
R1198 VP.n43 VP.n4 0.189894
R1199 VP.n44 VP.n43 0.189894
R1200 VP.n45 VP.n44 0.189894
R1201 VP.n45 VP.n2 0.189894
R1202 VP.n50 VP.n2 0.189894
R1203 VP.n51 VP.n50 0.189894
R1204 VP.n52 VP.n51 0.189894
R1205 VP.n52 VP.n0 0.189894
R1206 VP.n56 VP.n0 0.189894
R1207 VP VP.n56 0.0516364
R1208 VDD1 VDD1.n0 238.375
R1209 VDD1.n3 VDD1.n2 238.261
R1210 VDD1.n3 VDD1.n1 238.261
R1211 VDD1.n5 VDD1.n4 237.356
R1212 VDD1.n5 VDD1.n3 33.6216
R1213 VDD1.n4 VDD1.t4 25.3851
R1214 VDD1.n4 VDD1.t6 25.3851
R1215 VDD1.n0 VDD1.t1 25.3851
R1216 VDD1.n0 VDD1.t3 25.3851
R1217 VDD1.n2 VDD1.t2 25.3851
R1218 VDD1.n2 VDD1.t7 25.3851
R1219 VDD1.n1 VDD1.t5 25.3851
R1220 VDD1.n1 VDD1.t0 25.3851
R1221 VDD1 VDD1.n5 0.903517
C0 VP VTAIL 1.93223f
C1 VDD2 VTAIL 3.68278f
C2 VDD1 VTAIL 3.63306f
C3 VN VP 4.73043f
C4 VN VDD2 0.94876f
C5 VN VDD1 0.157844f
C6 VDD2 VP 0.454373f
C7 VDD1 VP 1.24207f
C8 VDD1 VDD2 1.41008f
C9 VN VTAIL 1.91812f
C10 VDD2 B 3.58884f
C11 VDD1 B 3.928842f
C12 VTAIL B 2.881919f
C13 VN B 11.359744f
C14 VP B 10.296801f
C15 VDD1.t1 B 0.012519f
C16 VDD1.t3 B 0.012519f
C17 VDD1.n0 B 0.031405f
C18 VDD1.t5 B 0.012519f
C19 VDD1.t0 B 0.012519f
C20 VDD1.n1 B 0.031259f
C21 VDD1.t2 B 0.012519f
C22 VDD1.t7 B 0.012519f
C23 VDD1.n2 B 0.031259f
C24 VDD1.n3 B 1.60848f
C25 VDD1.t4 B 0.012519f
C26 VDD1.t6 B 0.012519f
C27 VDD1.n4 B 0.030322f
C28 VDD1.n5 B 1.38923f
C29 VP.n0 B 0.024286f
C30 VP.t0 B 0.057761f
C31 VP.n1 B 0.019739f
C32 VP.n2 B 0.024286f
C33 VP.t5 B 0.057761f
C34 VP.n3 B 0.035304f
C35 VP.n4 B 0.024286f
C36 VP.t7 B 0.057761f
C37 VP.n5 B 0.047474f
C38 VP.n6 B 0.024286f
C39 VP.t2 B 0.057761f
C40 VP.n7 B 0.115534f
C41 VP.n8 B 0.024286f
C42 VP.t1 B 0.057761f
C43 VP.n9 B 0.019739f
C44 VP.n10 B 0.024286f
C45 VP.t3 B 0.057761f
C46 VP.n11 B 0.035304f
C47 VP.n12 B 0.181132f
C48 VP.t4 B 0.057761f
C49 VP.t6 B 0.194404f
C50 VP.n13 B 0.094902f
C51 VP.n14 B 0.116398f
C52 VP.n15 B 0.039034f
C53 VP.n16 B 0.035304f
C54 VP.n17 B 0.024286f
C55 VP.n18 B 0.024286f
C56 VP.n19 B 0.024286f
C57 VP.n20 B 0.039034f
C58 VP.n21 B 0.055856f
C59 VP.n22 B 0.028806f
C60 VP.n23 B 0.047474f
C61 VP.n24 B 0.024286f
C62 VP.n25 B 0.024286f
C63 VP.n26 B 0.024286f
C64 VP.n27 B 0.048431f
C65 VP.n28 B 0.027027f
C66 VP.n29 B 0.115534f
C67 VP.n30 B 0.892841f
C68 VP.n31 B 0.915256f
C69 VP.n32 B 0.024286f
C70 VP.n33 B 0.027027f
C71 VP.n34 B 0.048431f
C72 VP.n35 B 0.019739f
C73 VP.n36 B 0.024286f
C74 VP.n37 B 0.024286f
C75 VP.n38 B 0.024286f
C76 VP.n39 B 0.028806f
C77 VP.n40 B 0.055856f
C78 VP.n41 B 0.039034f
C79 VP.n42 B 0.035304f
C80 VP.n43 B 0.024286f
C81 VP.n44 B 0.024286f
C82 VP.n45 B 0.024286f
C83 VP.n46 B 0.039034f
C84 VP.n47 B 0.055856f
C85 VP.n48 B 0.028806f
C86 VP.n49 B 0.047474f
C87 VP.n50 B 0.024286f
C88 VP.n51 B 0.024286f
C89 VP.n52 B 0.024286f
C90 VP.n53 B 0.048431f
C91 VP.n54 B 0.027027f
C92 VP.n55 B 0.115534f
C93 VP.n56 B 0.026191f
C94 VDD2.t6 B 0.01314f
C95 VDD2.t3 B 0.01314f
C96 VDD2.n0 B 0.032811f
C97 VDD2.t0 B 0.01314f
C98 VDD2.t7 B 0.01314f
C99 VDD2.n1 B 0.032811f
C100 VDD2.n2 B 1.64342f
C101 VDD2.t5 B 0.01314f
C102 VDD2.t1 B 0.01314f
C103 VDD2.n3 B 0.031828f
C104 VDD2.n4 B 1.43239f
C105 VDD2.t4 B 0.01314f
C106 VDD2.t2 B 0.01314f
C107 VDD2.n5 B 0.032805f
C108 VTAIL.t8 B 0.018446f
C109 VTAIL.t12 B 0.018446f
C110 VTAIL.n0 B 0.039268f
C111 VTAIL.n1 B 0.233032f
C112 VTAIL.t10 B 0.082238f
C113 VTAIL.n2 B 0.280065f
C114 VTAIL.t6 B 0.082238f
C115 VTAIL.n3 B 0.280065f
C116 VTAIL.t4 B 0.018446f
C117 VTAIL.t0 B 0.018446f
C118 VTAIL.n4 B 0.039268f
C119 VTAIL.n5 B 0.4128f
C120 VTAIL.t7 B 0.082238f
C121 VTAIL.n6 B 0.891499f
C122 VTAIL.t11 B 0.082238f
C123 VTAIL.n7 B 0.891499f
C124 VTAIL.t14 B 0.018446f
C125 VTAIL.t15 B 0.018446f
C126 VTAIL.n8 B 0.039268f
C127 VTAIL.n9 B 0.4128f
C128 VTAIL.t9 B 0.082238f
C129 VTAIL.n10 B 0.280065f
C130 VTAIL.t2 B 0.082238f
C131 VTAIL.n11 B 0.280065f
C132 VTAIL.t3 B 0.018446f
C133 VTAIL.t1 B 0.018446f
C134 VTAIL.n12 B 0.039268f
C135 VTAIL.n13 B 0.4128f
C136 VTAIL.t5 B 0.082238f
C137 VTAIL.n14 B 0.891499f
C138 VTAIL.t13 B 0.082238f
C139 VTAIL.n15 B 0.885888f
C140 VN.n0 B 0.024111f
C141 VN.t0 B 0.057345f
C142 VN.n1 B 0.019597f
C143 VN.n2 B 0.024111f
C144 VN.t7 B 0.057345f
C145 VN.n3 B 0.035049f
C146 VN.n4 B 0.179826f
C147 VN.t4 B 0.057345f
C148 VN.t1 B 0.193002f
C149 VN.n5 B 0.094217f
C150 VN.n6 B 0.115559f
C151 VN.n7 B 0.038752f
C152 VN.n8 B 0.035049f
C153 VN.n9 B 0.024111f
C154 VN.n10 B 0.024111f
C155 VN.n11 B 0.024111f
C156 VN.n12 B 0.038752f
C157 VN.n13 B 0.055453f
C158 VN.n14 B 0.028598f
C159 VN.n15 B 0.047131f
C160 VN.n16 B 0.024111f
C161 VN.n17 B 0.024111f
C162 VN.n18 B 0.024111f
C163 VN.n19 B 0.048082f
C164 VN.n20 B 0.026833f
C165 VN.n21 B 0.1147f
C166 VN.n22 B 0.026002f
C167 VN.n23 B 0.024111f
C168 VN.t2 B 0.057345f
C169 VN.n24 B 0.019597f
C170 VN.n25 B 0.024111f
C171 VN.t6 B 0.057345f
C172 VN.n26 B 0.035049f
C173 VN.n27 B 0.179826f
C174 VN.t3 B 0.057345f
C175 VN.t5 B 0.193002f
C176 VN.n28 B 0.094217f
C177 VN.n29 B 0.115559f
C178 VN.n30 B 0.038752f
C179 VN.n31 B 0.035049f
C180 VN.n32 B 0.024111f
C181 VN.n33 B 0.024111f
C182 VN.n34 B 0.024111f
C183 VN.n35 B 0.038752f
C184 VN.n36 B 0.055453f
C185 VN.n37 B 0.028598f
C186 VN.n38 B 0.047131f
C187 VN.n39 B 0.024111f
C188 VN.n40 B 0.024111f
C189 VN.n41 B 0.024111f
C190 VN.n42 B 0.048082f
C191 VN.n43 B 0.026833f
C192 VN.n44 B 0.1147f
C193 VN.n45 B 0.902305f
.ends

