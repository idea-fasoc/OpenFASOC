* NGSPICE file created from diff_pair_sample_0597.ext - technology: sky130A

.subckt diff_pair_sample_0597 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t1 w_n3670_n4802# sky130_fd_pr__pfet_01v8 ad=3.16305 pd=19.5 as=3.16305 ps=19.5 w=19.17 l=2.37
X1 VTAIL.t5 VN.t0 VDD2.t7 w_n3670_n4802# sky130_fd_pr__pfet_01v8 ad=7.4763 pd=39.12 as=3.16305 ps=19.5 w=19.17 l=2.37
X2 B.t11 B.t9 B.t10 w_n3670_n4802# sky130_fd_pr__pfet_01v8 ad=7.4763 pd=39.12 as=0 ps=0 w=19.17 l=2.37
X3 VDD2.t6 VN.t1 VTAIL.t0 w_n3670_n4802# sky130_fd_pr__pfet_01v8 ad=3.16305 pd=19.5 as=7.4763 ps=39.12 w=19.17 l=2.37
X4 VDD1.t0 VP.t1 VTAIL.t14 w_n3670_n4802# sky130_fd_pr__pfet_01v8 ad=3.16305 pd=19.5 as=3.16305 ps=19.5 w=19.17 l=2.37
X5 VTAIL.t13 VP.t2 VDD1.t3 w_n3670_n4802# sky130_fd_pr__pfet_01v8 ad=7.4763 pd=39.12 as=3.16305 ps=19.5 w=19.17 l=2.37
X6 VTAIL.t3 VN.t2 VDD2.t5 w_n3670_n4802# sky130_fd_pr__pfet_01v8 ad=7.4763 pd=39.12 as=3.16305 ps=19.5 w=19.17 l=2.37
X7 VDD2.t4 VN.t3 VTAIL.t4 w_n3670_n4802# sky130_fd_pr__pfet_01v8 ad=3.16305 pd=19.5 as=7.4763 ps=39.12 w=19.17 l=2.37
X8 VTAIL.t6 VN.t4 VDD2.t3 w_n3670_n4802# sky130_fd_pr__pfet_01v8 ad=3.16305 pd=19.5 as=3.16305 ps=19.5 w=19.17 l=2.37
X9 VTAIL.t12 VP.t3 VDD1.t2 w_n3670_n4802# sky130_fd_pr__pfet_01v8 ad=3.16305 pd=19.5 as=3.16305 ps=19.5 w=19.17 l=2.37
X10 B.t8 B.t6 B.t7 w_n3670_n4802# sky130_fd_pr__pfet_01v8 ad=7.4763 pd=39.12 as=0 ps=0 w=19.17 l=2.37
X11 VDD1.t5 VP.t4 VTAIL.t11 w_n3670_n4802# sky130_fd_pr__pfet_01v8 ad=3.16305 pd=19.5 as=7.4763 ps=39.12 w=19.17 l=2.37
X12 B.t5 B.t3 B.t4 w_n3670_n4802# sky130_fd_pr__pfet_01v8 ad=7.4763 pd=39.12 as=0 ps=0 w=19.17 l=2.37
X13 VDD1.t4 VP.t5 VTAIL.t10 w_n3670_n4802# sky130_fd_pr__pfet_01v8 ad=3.16305 pd=19.5 as=3.16305 ps=19.5 w=19.17 l=2.37
X14 VDD2.t2 VN.t5 VTAIL.t1 w_n3670_n4802# sky130_fd_pr__pfet_01v8 ad=3.16305 pd=19.5 as=3.16305 ps=19.5 w=19.17 l=2.37
X15 B.t2 B.t0 B.t1 w_n3670_n4802# sky130_fd_pr__pfet_01v8 ad=7.4763 pd=39.12 as=0 ps=0 w=19.17 l=2.37
X16 VTAIL.t9 VP.t6 VDD1.t7 w_n3670_n4802# sky130_fd_pr__pfet_01v8 ad=7.4763 pd=39.12 as=3.16305 ps=19.5 w=19.17 l=2.37
X17 VDD2.t1 VN.t6 VTAIL.t7 w_n3670_n4802# sky130_fd_pr__pfet_01v8 ad=3.16305 pd=19.5 as=3.16305 ps=19.5 w=19.17 l=2.37
X18 VTAIL.t2 VN.t7 VDD2.t0 w_n3670_n4802# sky130_fd_pr__pfet_01v8 ad=3.16305 pd=19.5 as=3.16305 ps=19.5 w=19.17 l=2.37
X19 VDD1.t6 VP.t7 VTAIL.t8 w_n3670_n4802# sky130_fd_pr__pfet_01v8 ad=3.16305 pd=19.5 as=7.4763 ps=39.12 w=19.17 l=2.37
R0 VP.n15 VP.t2 227.355
R1 VP.n36 VP.t6 194.935
R2 VP.n43 VP.t1 194.935
R3 VP.n55 VP.t3 194.935
R4 VP.n63 VP.t7 194.935
R5 VP.n33 VP.t4 194.935
R6 VP.n25 VP.t0 194.935
R7 VP.n14 VP.t5 194.935
R8 VP.n16 VP.n13 161.3
R9 VP.n18 VP.n17 161.3
R10 VP.n19 VP.n12 161.3
R11 VP.n21 VP.n20 161.3
R12 VP.n22 VP.n11 161.3
R13 VP.n24 VP.n23 161.3
R14 VP.n26 VP.n10 161.3
R15 VP.n28 VP.n27 161.3
R16 VP.n29 VP.n9 161.3
R17 VP.n31 VP.n30 161.3
R18 VP.n32 VP.n8 161.3
R19 VP.n62 VP.n0 161.3
R20 VP.n61 VP.n60 161.3
R21 VP.n59 VP.n1 161.3
R22 VP.n58 VP.n57 161.3
R23 VP.n56 VP.n2 161.3
R24 VP.n54 VP.n53 161.3
R25 VP.n52 VP.n3 161.3
R26 VP.n51 VP.n50 161.3
R27 VP.n49 VP.n4 161.3
R28 VP.n48 VP.n47 161.3
R29 VP.n46 VP.n5 161.3
R30 VP.n45 VP.n44 161.3
R31 VP.n42 VP.n6 161.3
R32 VP.n41 VP.n40 161.3
R33 VP.n39 VP.n7 161.3
R34 VP.n38 VP.n37 161.3
R35 VP.n36 VP.n35 96.0763
R36 VP.n64 VP.n63 96.0763
R37 VP.n34 VP.n33 96.0763
R38 VP.n15 VP.n14 67.2582
R39 VP.n50 VP.n49 56.5193
R40 VP.n20 VP.n19 56.5193
R41 VP.n35 VP.n34 55.2875
R42 VP.n42 VP.n41 45.3497
R43 VP.n57 VP.n1 45.3497
R44 VP.n27 VP.n9 45.3497
R45 VP.n41 VP.n7 35.6371
R46 VP.n61 VP.n1 35.6371
R47 VP.n31 VP.n9 35.6371
R48 VP.n37 VP.n7 24.4675
R49 VP.n44 VP.n42 24.4675
R50 VP.n48 VP.n5 24.4675
R51 VP.n49 VP.n48 24.4675
R52 VP.n50 VP.n3 24.4675
R53 VP.n54 VP.n3 24.4675
R54 VP.n57 VP.n56 24.4675
R55 VP.n62 VP.n61 24.4675
R56 VP.n32 VP.n31 24.4675
R57 VP.n20 VP.n11 24.4675
R58 VP.n24 VP.n11 24.4675
R59 VP.n27 VP.n26 24.4675
R60 VP.n18 VP.n13 24.4675
R61 VP.n19 VP.n18 24.4675
R62 VP.n44 VP.n43 19.5741
R63 VP.n56 VP.n55 19.5741
R64 VP.n26 VP.n25 19.5741
R65 VP.n37 VP.n36 14.6807
R66 VP.n63 VP.n62 14.6807
R67 VP.n33 VP.n32 14.6807
R68 VP.n16 VP.n15 9.52612
R69 VP.n43 VP.n5 4.8939
R70 VP.n55 VP.n54 4.8939
R71 VP.n25 VP.n24 4.8939
R72 VP.n14 VP.n13 4.8939
R73 VP.n34 VP.n8 0.278367
R74 VP.n38 VP.n35 0.278367
R75 VP.n64 VP.n0 0.278367
R76 VP.n17 VP.n16 0.189894
R77 VP.n17 VP.n12 0.189894
R78 VP.n21 VP.n12 0.189894
R79 VP.n22 VP.n21 0.189894
R80 VP.n23 VP.n22 0.189894
R81 VP.n23 VP.n10 0.189894
R82 VP.n28 VP.n10 0.189894
R83 VP.n29 VP.n28 0.189894
R84 VP.n30 VP.n29 0.189894
R85 VP.n30 VP.n8 0.189894
R86 VP.n39 VP.n38 0.189894
R87 VP.n40 VP.n39 0.189894
R88 VP.n40 VP.n6 0.189894
R89 VP.n45 VP.n6 0.189894
R90 VP.n46 VP.n45 0.189894
R91 VP.n47 VP.n46 0.189894
R92 VP.n47 VP.n4 0.189894
R93 VP.n51 VP.n4 0.189894
R94 VP.n52 VP.n51 0.189894
R95 VP.n53 VP.n52 0.189894
R96 VP.n53 VP.n2 0.189894
R97 VP.n58 VP.n2 0.189894
R98 VP.n59 VP.n58 0.189894
R99 VP.n60 VP.n59 0.189894
R100 VP.n60 VP.n0 0.189894
R101 VP VP.n64 0.153454
R102 VDD1 VDD1.n0 73.2647
R103 VDD1.n3 VDD1.n2 73.1499
R104 VDD1.n3 VDD1.n1 73.1499
R105 VDD1.n5 VDD1.n4 72.0425
R106 VDD1.n5 VDD1.n3 51.2983
R107 VDD1.n4 VDD1.t1 1.69612
R108 VDD1.n4 VDD1.t5 1.69612
R109 VDD1.n0 VDD1.t3 1.69612
R110 VDD1.n0 VDD1.t4 1.69612
R111 VDD1.n2 VDD1.t2 1.69612
R112 VDD1.n2 VDD1.t6 1.69612
R113 VDD1.n1 VDD1.t7 1.69612
R114 VDD1.n1 VDD1.t0 1.69612
R115 VDD1 VDD1.n5 1.1061
R116 VTAIL.n11 VTAIL.t13 57.0595
R117 VTAIL.n10 VTAIL.t4 57.0595
R118 VTAIL.n7 VTAIL.t5 57.0595
R119 VTAIL.n15 VTAIL.t0 57.0594
R120 VTAIL.n2 VTAIL.t3 57.0594
R121 VTAIL.n3 VTAIL.t8 57.0594
R122 VTAIL.n6 VTAIL.t9 57.0594
R123 VTAIL.n14 VTAIL.t11 57.0594
R124 VTAIL.n13 VTAIL.n12 55.3639
R125 VTAIL.n9 VTAIL.n8 55.3639
R126 VTAIL.n1 VTAIL.n0 55.3627
R127 VTAIL.n5 VTAIL.n4 55.3627
R128 VTAIL.n15 VTAIL.n14 31.2203
R129 VTAIL.n7 VTAIL.n6 31.2203
R130 VTAIL.n9 VTAIL.n7 2.32809
R131 VTAIL.n10 VTAIL.n9 2.32809
R132 VTAIL.n13 VTAIL.n11 2.32809
R133 VTAIL.n14 VTAIL.n13 2.32809
R134 VTAIL.n6 VTAIL.n5 2.32809
R135 VTAIL.n5 VTAIL.n3 2.32809
R136 VTAIL.n2 VTAIL.n1 2.32809
R137 VTAIL VTAIL.n15 2.2699
R138 VTAIL.n0 VTAIL.t7 1.69612
R139 VTAIL.n0 VTAIL.t6 1.69612
R140 VTAIL.n4 VTAIL.t14 1.69612
R141 VTAIL.n4 VTAIL.t12 1.69612
R142 VTAIL.n12 VTAIL.t10 1.69612
R143 VTAIL.n12 VTAIL.t15 1.69612
R144 VTAIL.n8 VTAIL.t1 1.69612
R145 VTAIL.n8 VTAIL.t2 1.69612
R146 VTAIL.n11 VTAIL.n10 0.470328
R147 VTAIL.n3 VTAIL.n2 0.470328
R148 VTAIL VTAIL.n1 0.0586897
R149 VN.n7 VN.t2 227.355
R150 VN.n34 VN.t3 227.355
R151 VN.n6 VN.t6 194.935
R152 VN.n17 VN.t4 194.935
R153 VN.n25 VN.t1 194.935
R154 VN.n33 VN.t7 194.935
R155 VN.n44 VN.t5 194.935
R156 VN.n52 VN.t0 194.935
R157 VN.n51 VN.n27 161.3
R158 VN.n50 VN.n49 161.3
R159 VN.n48 VN.n28 161.3
R160 VN.n47 VN.n46 161.3
R161 VN.n45 VN.n29 161.3
R162 VN.n43 VN.n42 161.3
R163 VN.n41 VN.n30 161.3
R164 VN.n40 VN.n39 161.3
R165 VN.n38 VN.n31 161.3
R166 VN.n37 VN.n36 161.3
R167 VN.n35 VN.n32 161.3
R168 VN.n24 VN.n0 161.3
R169 VN.n23 VN.n22 161.3
R170 VN.n21 VN.n1 161.3
R171 VN.n20 VN.n19 161.3
R172 VN.n18 VN.n2 161.3
R173 VN.n16 VN.n15 161.3
R174 VN.n14 VN.n3 161.3
R175 VN.n13 VN.n12 161.3
R176 VN.n11 VN.n4 161.3
R177 VN.n10 VN.n9 161.3
R178 VN.n8 VN.n5 161.3
R179 VN.n26 VN.n25 96.0763
R180 VN.n53 VN.n52 96.0763
R181 VN.n7 VN.n6 67.2582
R182 VN.n34 VN.n33 67.2582
R183 VN.n12 VN.n11 56.5193
R184 VN.n39 VN.n38 56.5193
R185 VN VN.n53 55.5663
R186 VN.n19 VN.n1 45.3497
R187 VN.n46 VN.n28 45.3497
R188 VN.n23 VN.n1 35.6371
R189 VN.n50 VN.n28 35.6371
R190 VN.n10 VN.n5 24.4675
R191 VN.n11 VN.n10 24.4675
R192 VN.n12 VN.n3 24.4675
R193 VN.n16 VN.n3 24.4675
R194 VN.n19 VN.n18 24.4675
R195 VN.n24 VN.n23 24.4675
R196 VN.n38 VN.n37 24.4675
R197 VN.n37 VN.n32 24.4675
R198 VN.n46 VN.n45 24.4675
R199 VN.n43 VN.n30 24.4675
R200 VN.n39 VN.n30 24.4675
R201 VN.n51 VN.n50 24.4675
R202 VN.n18 VN.n17 19.5741
R203 VN.n45 VN.n44 19.5741
R204 VN.n25 VN.n24 14.6807
R205 VN.n52 VN.n51 14.6807
R206 VN.n35 VN.n34 9.52612
R207 VN.n8 VN.n7 9.52612
R208 VN.n6 VN.n5 4.8939
R209 VN.n17 VN.n16 4.8939
R210 VN.n33 VN.n32 4.8939
R211 VN.n44 VN.n43 4.8939
R212 VN.n53 VN.n27 0.278367
R213 VN.n26 VN.n0 0.278367
R214 VN.n49 VN.n27 0.189894
R215 VN.n49 VN.n48 0.189894
R216 VN.n48 VN.n47 0.189894
R217 VN.n47 VN.n29 0.189894
R218 VN.n42 VN.n29 0.189894
R219 VN.n42 VN.n41 0.189894
R220 VN.n41 VN.n40 0.189894
R221 VN.n40 VN.n31 0.189894
R222 VN.n36 VN.n31 0.189894
R223 VN.n36 VN.n35 0.189894
R224 VN.n9 VN.n8 0.189894
R225 VN.n9 VN.n4 0.189894
R226 VN.n13 VN.n4 0.189894
R227 VN.n14 VN.n13 0.189894
R228 VN.n15 VN.n14 0.189894
R229 VN.n15 VN.n2 0.189894
R230 VN.n20 VN.n2 0.189894
R231 VN.n21 VN.n20 0.189894
R232 VN.n22 VN.n21 0.189894
R233 VN.n22 VN.n0 0.189894
R234 VN VN.n26 0.153454
R235 VDD2.n2 VDD2.n1 73.1499
R236 VDD2.n2 VDD2.n0 73.1499
R237 VDD2 VDD2.n5 73.1481
R238 VDD2.n4 VDD2.n3 72.0427
R239 VDD2.n4 VDD2.n2 50.7153
R240 VDD2.n5 VDD2.t0 1.69612
R241 VDD2.n5 VDD2.t4 1.69612
R242 VDD2.n3 VDD2.t7 1.69612
R243 VDD2.n3 VDD2.t2 1.69612
R244 VDD2.n1 VDD2.t3 1.69612
R245 VDD2.n1 VDD2.t6 1.69612
R246 VDD2.n0 VDD2.t5 1.69612
R247 VDD2.n0 VDD2.t1 1.69612
R248 VDD2 VDD2.n4 1.22248
R249 B.n663 B.n662 585
R250 B.n664 B.n97 585
R251 B.n666 B.n665 585
R252 B.n667 B.n96 585
R253 B.n669 B.n668 585
R254 B.n670 B.n95 585
R255 B.n672 B.n671 585
R256 B.n673 B.n94 585
R257 B.n675 B.n674 585
R258 B.n676 B.n93 585
R259 B.n678 B.n677 585
R260 B.n679 B.n92 585
R261 B.n681 B.n680 585
R262 B.n682 B.n91 585
R263 B.n684 B.n683 585
R264 B.n685 B.n90 585
R265 B.n687 B.n686 585
R266 B.n688 B.n89 585
R267 B.n690 B.n689 585
R268 B.n691 B.n88 585
R269 B.n693 B.n692 585
R270 B.n694 B.n87 585
R271 B.n696 B.n695 585
R272 B.n697 B.n86 585
R273 B.n699 B.n698 585
R274 B.n700 B.n85 585
R275 B.n702 B.n701 585
R276 B.n703 B.n84 585
R277 B.n705 B.n704 585
R278 B.n706 B.n83 585
R279 B.n708 B.n707 585
R280 B.n709 B.n82 585
R281 B.n711 B.n710 585
R282 B.n712 B.n81 585
R283 B.n714 B.n713 585
R284 B.n715 B.n80 585
R285 B.n717 B.n716 585
R286 B.n718 B.n79 585
R287 B.n720 B.n719 585
R288 B.n721 B.n78 585
R289 B.n723 B.n722 585
R290 B.n724 B.n77 585
R291 B.n726 B.n725 585
R292 B.n727 B.n76 585
R293 B.n729 B.n728 585
R294 B.n730 B.n75 585
R295 B.n732 B.n731 585
R296 B.n733 B.n74 585
R297 B.n735 B.n734 585
R298 B.n736 B.n73 585
R299 B.n738 B.n737 585
R300 B.n739 B.n72 585
R301 B.n741 B.n740 585
R302 B.n742 B.n71 585
R303 B.n744 B.n743 585
R304 B.n745 B.n70 585
R305 B.n747 B.n746 585
R306 B.n748 B.n69 585
R307 B.n750 B.n749 585
R308 B.n751 B.n68 585
R309 B.n753 B.n752 585
R310 B.n754 B.n67 585
R311 B.n756 B.n755 585
R312 B.n758 B.n757 585
R313 B.n759 B.n63 585
R314 B.n761 B.n760 585
R315 B.n762 B.n62 585
R316 B.n764 B.n763 585
R317 B.n765 B.n61 585
R318 B.n767 B.n766 585
R319 B.n768 B.n60 585
R320 B.n770 B.n769 585
R321 B.n772 B.n57 585
R322 B.n774 B.n773 585
R323 B.n775 B.n56 585
R324 B.n777 B.n776 585
R325 B.n778 B.n55 585
R326 B.n780 B.n779 585
R327 B.n781 B.n54 585
R328 B.n783 B.n782 585
R329 B.n784 B.n53 585
R330 B.n786 B.n785 585
R331 B.n787 B.n52 585
R332 B.n789 B.n788 585
R333 B.n790 B.n51 585
R334 B.n792 B.n791 585
R335 B.n793 B.n50 585
R336 B.n795 B.n794 585
R337 B.n796 B.n49 585
R338 B.n798 B.n797 585
R339 B.n799 B.n48 585
R340 B.n801 B.n800 585
R341 B.n802 B.n47 585
R342 B.n804 B.n803 585
R343 B.n805 B.n46 585
R344 B.n807 B.n806 585
R345 B.n808 B.n45 585
R346 B.n810 B.n809 585
R347 B.n811 B.n44 585
R348 B.n813 B.n812 585
R349 B.n814 B.n43 585
R350 B.n816 B.n815 585
R351 B.n817 B.n42 585
R352 B.n819 B.n818 585
R353 B.n820 B.n41 585
R354 B.n822 B.n821 585
R355 B.n823 B.n40 585
R356 B.n825 B.n824 585
R357 B.n826 B.n39 585
R358 B.n828 B.n827 585
R359 B.n829 B.n38 585
R360 B.n831 B.n830 585
R361 B.n832 B.n37 585
R362 B.n834 B.n833 585
R363 B.n835 B.n36 585
R364 B.n837 B.n836 585
R365 B.n838 B.n35 585
R366 B.n840 B.n839 585
R367 B.n841 B.n34 585
R368 B.n843 B.n842 585
R369 B.n844 B.n33 585
R370 B.n846 B.n845 585
R371 B.n847 B.n32 585
R372 B.n849 B.n848 585
R373 B.n850 B.n31 585
R374 B.n852 B.n851 585
R375 B.n853 B.n30 585
R376 B.n855 B.n854 585
R377 B.n856 B.n29 585
R378 B.n858 B.n857 585
R379 B.n859 B.n28 585
R380 B.n861 B.n860 585
R381 B.n862 B.n27 585
R382 B.n864 B.n863 585
R383 B.n865 B.n26 585
R384 B.n661 B.n98 585
R385 B.n660 B.n659 585
R386 B.n658 B.n99 585
R387 B.n657 B.n656 585
R388 B.n655 B.n100 585
R389 B.n654 B.n653 585
R390 B.n652 B.n101 585
R391 B.n651 B.n650 585
R392 B.n649 B.n102 585
R393 B.n648 B.n647 585
R394 B.n646 B.n103 585
R395 B.n645 B.n644 585
R396 B.n643 B.n104 585
R397 B.n642 B.n641 585
R398 B.n640 B.n105 585
R399 B.n639 B.n638 585
R400 B.n637 B.n106 585
R401 B.n636 B.n635 585
R402 B.n634 B.n107 585
R403 B.n633 B.n632 585
R404 B.n631 B.n108 585
R405 B.n630 B.n629 585
R406 B.n628 B.n109 585
R407 B.n627 B.n626 585
R408 B.n625 B.n110 585
R409 B.n624 B.n623 585
R410 B.n622 B.n111 585
R411 B.n621 B.n620 585
R412 B.n619 B.n112 585
R413 B.n618 B.n617 585
R414 B.n616 B.n113 585
R415 B.n615 B.n614 585
R416 B.n613 B.n114 585
R417 B.n612 B.n611 585
R418 B.n610 B.n115 585
R419 B.n609 B.n608 585
R420 B.n607 B.n116 585
R421 B.n606 B.n605 585
R422 B.n604 B.n117 585
R423 B.n603 B.n602 585
R424 B.n601 B.n118 585
R425 B.n600 B.n599 585
R426 B.n598 B.n119 585
R427 B.n597 B.n596 585
R428 B.n595 B.n120 585
R429 B.n594 B.n593 585
R430 B.n592 B.n121 585
R431 B.n591 B.n590 585
R432 B.n589 B.n122 585
R433 B.n588 B.n587 585
R434 B.n586 B.n123 585
R435 B.n585 B.n584 585
R436 B.n583 B.n124 585
R437 B.n582 B.n581 585
R438 B.n580 B.n125 585
R439 B.n579 B.n578 585
R440 B.n577 B.n126 585
R441 B.n576 B.n575 585
R442 B.n574 B.n127 585
R443 B.n573 B.n572 585
R444 B.n571 B.n128 585
R445 B.n570 B.n569 585
R446 B.n568 B.n129 585
R447 B.n567 B.n566 585
R448 B.n565 B.n130 585
R449 B.n564 B.n563 585
R450 B.n562 B.n131 585
R451 B.n561 B.n560 585
R452 B.n559 B.n132 585
R453 B.n558 B.n557 585
R454 B.n556 B.n133 585
R455 B.n555 B.n554 585
R456 B.n553 B.n134 585
R457 B.n552 B.n551 585
R458 B.n550 B.n135 585
R459 B.n549 B.n548 585
R460 B.n547 B.n136 585
R461 B.n546 B.n545 585
R462 B.n544 B.n137 585
R463 B.n543 B.n542 585
R464 B.n541 B.n138 585
R465 B.n540 B.n539 585
R466 B.n538 B.n139 585
R467 B.n537 B.n536 585
R468 B.n535 B.n140 585
R469 B.n534 B.n533 585
R470 B.n532 B.n141 585
R471 B.n531 B.n530 585
R472 B.n529 B.n142 585
R473 B.n528 B.n527 585
R474 B.n526 B.n143 585
R475 B.n525 B.n524 585
R476 B.n523 B.n144 585
R477 B.n522 B.n521 585
R478 B.n520 B.n145 585
R479 B.n519 B.n518 585
R480 B.n517 B.n146 585
R481 B.n313 B.n218 585
R482 B.n315 B.n314 585
R483 B.n316 B.n217 585
R484 B.n318 B.n317 585
R485 B.n319 B.n216 585
R486 B.n321 B.n320 585
R487 B.n322 B.n215 585
R488 B.n324 B.n323 585
R489 B.n325 B.n214 585
R490 B.n327 B.n326 585
R491 B.n328 B.n213 585
R492 B.n330 B.n329 585
R493 B.n331 B.n212 585
R494 B.n333 B.n332 585
R495 B.n334 B.n211 585
R496 B.n336 B.n335 585
R497 B.n337 B.n210 585
R498 B.n339 B.n338 585
R499 B.n340 B.n209 585
R500 B.n342 B.n341 585
R501 B.n343 B.n208 585
R502 B.n345 B.n344 585
R503 B.n346 B.n207 585
R504 B.n348 B.n347 585
R505 B.n349 B.n206 585
R506 B.n351 B.n350 585
R507 B.n352 B.n205 585
R508 B.n354 B.n353 585
R509 B.n355 B.n204 585
R510 B.n357 B.n356 585
R511 B.n358 B.n203 585
R512 B.n360 B.n359 585
R513 B.n361 B.n202 585
R514 B.n363 B.n362 585
R515 B.n364 B.n201 585
R516 B.n366 B.n365 585
R517 B.n367 B.n200 585
R518 B.n369 B.n368 585
R519 B.n370 B.n199 585
R520 B.n372 B.n371 585
R521 B.n373 B.n198 585
R522 B.n375 B.n374 585
R523 B.n376 B.n197 585
R524 B.n378 B.n377 585
R525 B.n379 B.n196 585
R526 B.n381 B.n380 585
R527 B.n382 B.n195 585
R528 B.n384 B.n383 585
R529 B.n385 B.n194 585
R530 B.n387 B.n386 585
R531 B.n388 B.n193 585
R532 B.n390 B.n389 585
R533 B.n391 B.n192 585
R534 B.n393 B.n392 585
R535 B.n394 B.n191 585
R536 B.n396 B.n395 585
R537 B.n397 B.n190 585
R538 B.n399 B.n398 585
R539 B.n400 B.n189 585
R540 B.n402 B.n401 585
R541 B.n403 B.n188 585
R542 B.n405 B.n404 585
R543 B.n406 B.n185 585
R544 B.n409 B.n408 585
R545 B.n410 B.n184 585
R546 B.n412 B.n411 585
R547 B.n413 B.n183 585
R548 B.n415 B.n414 585
R549 B.n416 B.n182 585
R550 B.n418 B.n417 585
R551 B.n419 B.n181 585
R552 B.n421 B.n420 585
R553 B.n423 B.n422 585
R554 B.n424 B.n177 585
R555 B.n426 B.n425 585
R556 B.n427 B.n176 585
R557 B.n429 B.n428 585
R558 B.n430 B.n175 585
R559 B.n432 B.n431 585
R560 B.n433 B.n174 585
R561 B.n435 B.n434 585
R562 B.n436 B.n173 585
R563 B.n438 B.n437 585
R564 B.n439 B.n172 585
R565 B.n441 B.n440 585
R566 B.n442 B.n171 585
R567 B.n444 B.n443 585
R568 B.n445 B.n170 585
R569 B.n447 B.n446 585
R570 B.n448 B.n169 585
R571 B.n450 B.n449 585
R572 B.n451 B.n168 585
R573 B.n453 B.n452 585
R574 B.n454 B.n167 585
R575 B.n456 B.n455 585
R576 B.n457 B.n166 585
R577 B.n459 B.n458 585
R578 B.n460 B.n165 585
R579 B.n462 B.n461 585
R580 B.n463 B.n164 585
R581 B.n465 B.n464 585
R582 B.n466 B.n163 585
R583 B.n468 B.n467 585
R584 B.n469 B.n162 585
R585 B.n471 B.n470 585
R586 B.n472 B.n161 585
R587 B.n474 B.n473 585
R588 B.n475 B.n160 585
R589 B.n477 B.n476 585
R590 B.n478 B.n159 585
R591 B.n480 B.n479 585
R592 B.n481 B.n158 585
R593 B.n483 B.n482 585
R594 B.n484 B.n157 585
R595 B.n486 B.n485 585
R596 B.n487 B.n156 585
R597 B.n489 B.n488 585
R598 B.n490 B.n155 585
R599 B.n492 B.n491 585
R600 B.n493 B.n154 585
R601 B.n495 B.n494 585
R602 B.n496 B.n153 585
R603 B.n498 B.n497 585
R604 B.n499 B.n152 585
R605 B.n501 B.n500 585
R606 B.n502 B.n151 585
R607 B.n504 B.n503 585
R608 B.n505 B.n150 585
R609 B.n507 B.n506 585
R610 B.n508 B.n149 585
R611 B.n510 B.n509 585
R612 B.n511 B.n148 585
R613 B.n513 B.n512 585
R614 B.n514 B.n147 585
R615 B.n516 B.n515 585
R616 B.n312 B.n311 585
R617 B.n310 B.n219 585
R618 B.n309 B.n308 585
R619 B.n307 B.n220 585
R620 B.n306 B.n305 585
R621 B.n304 B.n221 585
R622 B.n303 B.n302 585
R623 B.n301 B.n222 585
R624 B.n300 B.n299 585
R625 B.n298 B.n223 585
R626 B.n297 B.n296 585
R627 B.n295 B.n224 585
R628 B.n294 B.n293 585
R629 B.n292 B.n225 585
R630 B.n291 B.n290 585
R631 B.n289 B.n226 585
R632 B.n288 B.n287 585
R633 B.n286 B.n227 585
R634 B.n285 B.n284 585
R635 B.n283 B.n228 585
R636 B.n282 B.n281 585
R637 B.n280 B.n229 585
R638 B.n279 B.n278 585
R639 B.n277 B.n230 585
R640 B.n276 B.n275 585
R641 B.n274 B.n231 585
R642 B.n273 B.n272 585
R643 B.n271 B.n232 585
R644 B.n270 B.n269 585
R645 B.n268 B.n233 585
R646 B.n267 B.n266 585
R647 B.n265 B.n234 585
R648 B.n264 B.n263 585
R649 B.n262 B.n235 585
R650 B.n261 B.n260 585
R651 B.n259 B.n236 585
R652 B.n258 B.n257 585
R653 B.n256 B.n237 585
R654 B.n255 B.n254 585
R655 B.n253 B.n238 585
R656 B.n252 B.n251 585
R657 B.n250 B.n239 585
R658 B.n249 B.n248 585
R659 B.n247 B.n240 585
R660 B.n246 B.n245 585
R661 B.n244 B.n241 585
R662 B.n243 B.n242 585
R663 B.n2 B.n0 585
R664 B.n937 B.n1 585
R665 B.n936 B.n935 585
R666 B.n934 B.n3 585
R667 B.n933 B.n932 585
R668 B.n931 B.n4 585
R669 B.n930 B.n929 585
R670 B.n928 B.n5 585
R671 B.n927 B.n926 585
R672 B.n925 B.n6 585
R673 B.n924 B.n923 585
R674 B.n922 B.n7 585
R675 B.n921 B.n920 585
R676 B.n919 B.n8 585
R677 B.n918 B.n917 585
R678 B.n916 B.n9 585
R679 B.n915 B.n914 585
R680 B.n913 B.n10 585
R681 B.n912 B.n911 585
R682 B.n910 B.n11 585
R683 B.n909 B.n908 585
R684 B.n907 B.n12 585
R685 B.n906 B.n905 585
R686 B.n904 B.n13 585
R687 B.n903 B.n902 585
R688 B.n901 B.n14 585
R689 B.n900 B.n899 585
R690 B.n898 B.n15 585
R691 B.n897 B.n896 585
R692 B.n895 B.n16 585
R693 B.n894 B.n893 585
R694 B.n892 B.n17 585
R695 B.n891 B.n890 585
R696 B.n889 B.n18 585
R697 B.n888 B.n887 585
R698 B.n886 B.n19 585
R699 B.n885 B.n884 585
R700 B.n883 B.n20 585
R701 B.n882 B.n881 585
R702 B.n880 B.n21 585
R703 B.n879 B.n878 585
R704 B.n877 B.n22 585
R705 B.n876 B.n875 585
R706 B.n874 B.n23 585
R707 B.n873 B.n872 585
R708 B.n871 B.n24 585
R709 B.n870 B.n869 585
R710 B.n868 B.n25 585
R711 B.n867 B.n866 585
R712 B.n939 B.n938 585
R713 B.n313 B.n312 468.476
R714 B.n866 B.n865 468.476
R715 B.n517 B.n516 468.476
R716 B.n662 B.n661 468.476
R717 B.n178 B.t6 402.608
R718 B.n186 B.t9 402.608
R719 B.n58 B.t3 402.608
R720 B.n64 B.t0 402.608
R721 B.n312 B.n219 163.367
R722 B.n308 B.n219 163.367
R723 B.n308 B.n307 163.367
R724 B.n307 B.n306 163.367
R725 B.n306 B.n221 163.367
R726 B.n302 B.n221 163.367
R727 B.n302 B.n301 163.367
R728 B.n301 B.n300 163.367
R729 B.n300 B.n223 163.367
R730 B.n296 B.n223 163.367
R731 B.n296 B.n295 163.367
R732 B.n295 B.n294 163.367
R733 B.n294 B.n225 163.367
R734 B.n290 B.n225 163.367
R735 B.n290 B.n289 163.367
R736 B.n289 B.n288 163.367
R737 B.n288 B.n227 163.367
R738 B.n284 B.n227 163.367
R739 B.n284 B.n283 163.367
R740 B.n283 B.n282 163.367
R741 B.n282 B.n229 163.367
R742 B.n278 B.n229 163.367
R743 B.n278 B.n277 163.367
R744 B.n277 B.n276 163.367
R745 B.n276 B.n231 163.367
R746 B.n272 B.n231 163.367
R747 B.n272 B.n271 163.367
R748 B.n271 B.n270 163.367
R749 B.n270 B.n233 163.367
R750 B.n266 B.n233 163.367
R751 B.n266 B.n265 163.367
R752 B.n265 B.n264 163.367
R753 B.n264 B.n235 163.367
R754 B.n260 B.n235 163.367
R755 B.n260 B.n259 163.367
R756 B.n259 B.n258 163.367
R757 B.n258 B.n237 163.367
R758 B.n254 B.n237 163.367
R759 B.n254 B.n253 163.367
R760 B.n253 B.n252 163.367
R761 B.n252 B.n239 163.367
R762 B.n248 B.n239 163.367
R763 B.n248 B.n247 163.367
R764 B.n247 B.n246 163.367
R765 B.n246 B.n241 163.367
R766 B.n242 B.n241 163.367
R767 B.n242 B.n2 163.367
R768 B.n938 B.n2 163.367
R769 B.n938 B.n937 163.367
R770 B.n937 B.n936 163.367
R771 B.n936 B.n3 163.367
R772 B.n932 B.n3 163.367
R773 B.n932 B.n931 163.367
R774 B.n931 B.n930 163.367
R775 B.n930 B.n5 163.367
R776 B.n926 B.n5 163.367
R777 B.n926 B.n925 163.367
R778 B.n925 B.n924 163.367
R779 B.n924 B.n7 163.367
R780 B.n920 B.n7 163.367
R781 B.n920 B.n919 163.367
R782 B.n919 B.n918 163.367
R783 B.n918 B.n9 163.367
R784 B.n914 B.n9 163.367
R785 B.n914 B.n913 163.367
R786 B.n913 B.n912 163.367
R787 B.n912 B.n11 163.367
R788 B.n908 B.n11 163.367
R789 B.n908 B.n907 163.367
R790 B.n907 B.n906 163.367
R791 B.n906 B.n13 163.367
R792 B.n902 B.n13 163.367
R793 B.n902 B.n901 163.367
R794 B.n901 B.n900 163.367
R795 B.n900 B.n15 163.367
R796 B.n896 B.n15 163.367
R797 B.n896 B.n895 163.367
R798 B.n895 B.n894 163.367
R799 B.n894 B.n17 163.367
R800 B.n890 B.n17 163.367
R801 B.n890 B.n889 163.367
R802 B.n889 B.n888 163.367
R803 B.n888 B.n19 163.367
R804 B.n884 B.n19 163.367
R805 B.n884 B.n883 163.367
R806 B.n883 B.n882 163.367
R807 B.n882 B.n21 163.367
R808 B.n878 B.n21 163.367
R809 B.n878 B.n877 163.367
R810 B.n877 B.n876 163.367
R811 B.n876 B.n23 163.367
R812 B.n872 B.n23 163.367
R813 B.n872 B.n871 163.367
R814 B.n871 B.n870 163.367
R815 B.n870 B.n25 163.367
R816 B.n866 B.n25 163.367
R817 B.n314 B.n313 163.367
R818 B.n314 B.n217 163.367
R819 B.n318 B.n217 163.367
R820 B.n319 B.n318 163.367
R821 B.n320 B.n319 163.367
R822 B.n320 B.n215 163.367
R823 B.n324 B.n215 163.367
R824 B.n325 B.n324 163.367
R825 B.n326 B.n325 163.367
R826 B.n326 B.n213 163.367
R827 B.n330 B.n213 163.367
R828 B.n331 B.n330 163.367
R829 B.n332 B.n331 163.367
R830 B.n332 B.n211 163.367
R831 B.n336 B.n211 163.367
R832 B.n337 B.n336 163.367
R833 B.n338 B.n337 163.367
R834 B.n338 B.n209 163.367
R835 B.n342 B.n209 163.367
R836 B.n343 B.n342 163.367
R837 B.n344 B.n343 163.367
R838 B.n344 B.n207 163.367
R839 B.n348 B.n207 163.367
R840 B.n349 B.n348 163.367
R841 B.n350 B.n349 163.367
R842 B.n350 B.n205 163.367
R843 B.n354 B.n205 163.367
R844 B.n355 B.n354 163.367
R845 B.n356 B.n355 163.367
R846 B.n356 B.n203 163.367
R847 B.n360 B.n203 163.367
R848 B.n361 B.n360 163.367
R849 B.n362 B.n361 163.367
R850 B.n362 B.n201 163.367
R851 B.n366 B.n201 163.367
R852 B.n367 B.n366 163.367
R853 B.n368 B.n367 163.367
R854 B.n368 B.n199 163.367
R855 B.n372 B.n199 163.367
R856 B.n373 B.n372 163.367
R857 B.n374 B.n373 163.367
R858 B.n374 B.n197 163.367
R859 B.n378 B.n197 163.367
R860 B.n379 B.n378 163.367
R861 B.n380 B.n379 163.367
R862 B.n380 B.n195 163.367
R863 B.n384 B.n195 163.367
R864 B.n385 B.n384 163.367
R865 B.n386 B.n385 163.367
R866 B.n386 B.n193 163.367
R867 B.n390 B.n193 163.367
R868 B.n391 B.n390 163.367
R869 B.n392 B.n391 163.367
R870 B.n392 B.n191 163.367
R871 B.n396 B.n191 163.367
R872 B.n397 B.n396 163.367
R873 B.n398 B.n397 163.367
R874 B.n398 B.n189 163.367
R875 B.n402 B.n189 163.367
R876 B.n403 B.n402 163.367
R877 B.n404 B.n403 163.367
R878 B.n404 B.n185 163.367
R879 B.n409 B.n185 163.367
R880 B.n410 B.n409 163.367
R881 B.n411 B.n410 163.367
R882 B.n411 B.n183 163.367
R883 B.n415 B.n183 163.367
R884 B.n416 B.n415 163.367
R885 B.n417 B.n416 163.367
R886 B.n417 B.n181 163.367
R887 B.n421 B.n181 163.367
R888 B.n422 B.n421 163.367
R889 B.n422 B.n177 163.367
R890 B.n426 B.n177 163.367
R891 B.n427 B.n426 163.367
R892 B.n428 B.n427 163.367
R893 B.n428 B.n175 163.367
R894 B.n432 B.n175 163.367
R895 B.n433 B.n432 163.367
R896 B.n434 B.n433 163.367
R897 B.n434 B.n173 163.367
R898 B.n438 B.n173 163.367
R899 B.n439 B.n438 163.367
R900 B.n440 B.n439 163.367
R901 B.n440 B.n171 163.367
R902 B.n444 B.n171 163.367
R903 B.n445 B.n444 163.367
R904 B.n446 B.n445 163.367
R905 B.n446 B.n169 163.367
R906 B.n450 B.n169 163.367
R907 B.n451 B.n450 163.367
R908 B.n452 B.n451 163.367
R909 B.n452 B.n167 163.367
R910 B.n456 B.n167 163.367
R911 B.n457 B.n456 163.367
R912 B.n458 B.n457 163.367
R913 B.n458 B.n165 163.367
R914 B.n462 B.n165 163.367
R915 B.n463 B.n462 163.367
R916 B.n464 B.n463 163.367
R917 B.n464 B.n163 163.367
R918 B.n468 B.n163 163.367
R919 B.n469 B.n468 163.367
R920 B.n470 B.n469 163.367
R921 B.n470 B.n161 163.367
R922 B.n474 B.n161 163.367
R923 B.n475 B.n474 163.367
R924 B.n476 B.n475 163.367
R925 B.n476 B.n159 163.367
R926 B.n480 B.n159 163.367
R927 B.n481 B.n480 163.367
R928 B.n482 B.n481 163.367
R929 B.n482 B.n157 163.367
R930 B.n486 B.n157 163.367
R931 B.n487 B.n486 163.367
R932 B.n488 B.n487 163.367
R933 B.n488 B.n155 163.367
R934 B.n492 B.n155 163.367
R935 B.n493 B.n492 163.367
R936 B.n494 B.n493 163.367
R937 B.n494 B.n153 163.367
R938 B.n498 B.n153 163.367
R939 B.n499 B.n498 163.367
R940 B.n500 B.n499 163.367
R941 B.n500 B.n151 163.367
R942 B.n504 B.n151 163.367
R943 B.n505 B.n504 163.367
R944 B.n506 B.n505 163.367
R945 B.n506 B.n149 163.367
R946 B.n510 B.n149 163.367
R947 B.n511 B.n510 163.367
R948 B.n512 B.n511 163.367
R949 B.n512 B.n147 163.367
R950 B.n516 B.n147 163.367
R951 B.n518 B.n517 163.367
R952 B.n518 B.n145 163.367
R953 B.n522 B.n145 163.367
R954 B.n523 B.n522 163.367
R955 B.n524 B.n523 163.367
R956 B.n524 B.n143 163.367
R957 B.n528 B.n143 163.367
R958 B.n529 B.n528 163.367
R959 B.n530 B.n529 163.367
R960 B.n530 B.n141 163.367
R961 B.n534 B.n141 163.367
R962 B.n535 B.n534 163.367
R963 B.n536 B.n535 163.367
R964 B.n536 B.n139 163.367
R965 B.n540 B.n139 163.367
R966 B.n541 B.n540 163.367
R967 B.n542 B.n541 163.367
R968 B.n542 B.n137 163.367
R969 B.n546 B.n137 163.367
R970 B.n547 B.n546 163.367
R971 B.n548 B.n547 163.367
R972 B.n548 B.n135 163.367
R973 B.n552 B.n135 163.367
R974 B.n553 B.n552 163.367
R975 B.n554 B.n553 163.367
R976 B.n554 B.n133 163.367
R977 B.n558 B.n133 163.367
R978 B.n559 B.n558 163.367
R979 B.n560 B.n559 163.367
R980 B.n560 B.n131 163.367
R981 B.n564 B.n131 163.367
R982 B.n565 B.n564 163.367
R983 B.n566 B.n565 163.367
R984 B.n566 B.n129 163.367
R985 B.n570 B.n129 163.367
R986 B.n571 B.n570 163.367
R987 B.n572 B.n571 163.367
R988 B.n572 B.n127 163.367
R989 B.n576 B.n127 163.367
R990 B.n577 B.n576 163.367
R991 B.n578 B.n577 163.367
R992 B.n578 B.n125 163.367
R993 B.n582 B.n125 163.367
R994 B.n583 B.n582 163.367
R995 B.n584 B.n583 163.367
R996 B.n584 B.n123 163.367
R997 B.n588 B.n123 163.367
R998 B.n589 B.n588 163.367
R999 B.n590 B.n589 163.367
R1000 B.n590 B.n121 163.367
R1001 B.n594 B.n121 163.367
R1002 B.n595 B.n594 163.367
R1003 B.n596 B.n595 163.367
R1004 B.n596 B.n119 163.367
R1005 B.n600 B.n119 163.367
R1006 B.n601 B.n600 163.367
R1007 B.n602 B.n601 163.367
R1008 B.n602 B.n117 163.367
R1009 B.n606 B.n117 163.367
R1010 B.n607 B.n606 163.367
R1011 B.n608 B.n607 163.367
R1012 B.n608 B.n115 163.367
R1013 B.n612 B.n115 163.367
R1014 B.n613 B.n612 163.367
R1015 B.n614 B.n613 163.367
R1016 B.n614 B.n113 163.367
R1017 B.n618 B.n113 163.367
R1018 B.n619 B.n618 163.367
R1019 B.n620 B.n619 163.367
R1020 B.n620 B.n111 163.367
R1021 B.n624 B.n111 163.367
R1022 B.n625 B.n624 163.367
R1023 B.n626 B.n625 163.367
R1024 B.n626 B.n109 163.367
R1025 B.n630 B.n109 163.367
R1026 B.n631 B.n630 163.367
R1027 B.n632 B.n631 163.367
R1028 B.n632 B.n107 163.367
R1029 B.n636 B.n107 163.367
R1030 B.n637 B.n636 163.367
R1031 B.n638 B.n637 163.367
R1032 B.n638 B.n105 163.367
R1033 B.n642 B.n105 163.367
R1034 B.n643 B.n642 163.367
R1035 B.n644 B.n643 163.367
R1036 B.n644 B.n103 163.367
R1037 B.n648 B.n103 163.367
R1038 B.n649 B.n648 163.367
R1039 B.n650 B.n649 163.367
R1040 B.n650 B.n101 163.367
R1041 B.n654 B.n101 163.367
R1042 B.n655 B.n654 163.367
R1043 B.n656 B.n655 163.367
R1044 B.n656 B.n99 163.367
R1045 B.n660 B.n99 163.367
R1046 B.n661 B.n660 163.367
R1047 B.n865 B.n864 163.367
R1048 B.n864 B.n27 163.367
R1049 B.n860 B.n27 163.367
R1050 B.n860 B.n859 163.367
R1051 B.n859 B.n858 163.367
R1052 B.n858 B.n29 163.367
R1053 B.n854 B.n29 163.367
R1054 B.n854 B.n853 163.367
R1055 B.n853 B.n852 163.367
R1056 B.n852 B.n31 163.367
R1057 B.n848 B.n31 163.367
R1058 B.n848 B.n847 163.367
R1059 B.n847 B.n846 163.367
R1060 B.n846 B.n33 163.367
R1061 B.n842 B.n33 163.367
R1062 B.n842 B.n841 163.367
R1063 B.n841 B.n840 163.367
R1064 B.n840 B.n35 163.367
R1065 B.n836 B.n35 163.367
R1066 B.n836 B.n835 163.367
R1067 B.n835 B.n834 163.367
R1068 B.n834 B.n37 163.367
R1069 B.n830 B.n37 163.367
R1070 B.n830 B.n829 163.367
R1071 B.n829 B.n828 163.367
R1072 B.n828 B.n39 163.367
R1073 B.n824 B.n39 163.367
R1074 B.n824 B.n823 163.367
R1075 B.n823 B.n822 163.367
R1076 B.n822 B.n41 163.367
R1077 B.n818 B.n41 163.367
R1078 B.n818 B.n817 163.367
R1079 B.n817 B.n816 163.367
R1080 B.n816 B.n43 163.367
R1081 B.n812 B.n43 163.367
R1082 B.n812 B.n811 163.367
R1083 B.n811 B.n810 163.367
R1084 B.n810 B.n45 163.367
R1085 B.n806 B.n45 163.367
R1086 B.n806 B.n805 163.367
R1087 B.n805 B.n804 163.367
R1088 B.n804 B.n47 163.367
R1089 B.n800 B.n47 163.367
R1090 B.n800 B.n799 163.367
R1091 B.n799 B.n798 163.367
R1092 B.n798 B.n49 163.367
R1093 B.n794 B.n49 163.367
R1094 B.n794 B.n793 163.367
R1095 B.n793 B.n792 163.367
R1096 B.n792 B.n51 163.367
R1097 B.n788 B.n51 163.367
R1098 B.n788 B.n787 163.367
R1099 B.n787 B.n786 163.367
R1100 B.n786 B.n53 163.367
R1101 B.n782 B.n53 163.367
R1102 B.n782 B.n781 163.367
R1103 B.n781 B.n780 163.367
R1104 B.n780 B.n55 163.367
R1105 B.n776 B.n55 163.367
R1106 B.n776 B.n775 163.367
R1107 B.n775 B.n774 163.367
R1108 B.n774 B.n57 163.367
R1109 B.n769 B.n57 163.367
R1110 B.n769 B.n768 163.367
R1111 B.n768 B.n767 163.367
R1112 B.n767 B.n61 163.367
R1113 B.n763 B.n61 163.367
R1114 B.n763 B.n762 163.367
R1115 B.n762 B.n761 163.367
R1116 B.n761 B.n63 163.367
R1117 B.n757 B.n63 163.367
R1118 B.n757 B.n756 163.367
R1119 B.n756 B.n67 163.367
R1120 B.n752 B.n67 163.367
R1121 B.n752 B.n751 163.367
R1122 B.n751 B.n750 163.367
R1123 B.n750 B.n69 163.367
R1124 B.n746 B.n69 163.367
R1125 B.n746 B.n745 163.367
R1126 B.n745 B.n744 163.367
R1127 B.n744 B.n71 163.367
R1128 B.n740 B.n71 163.367
R1129 B.n740 B.n739 163.367
R1130 B.n739 B.n738 163.367
R1131 B.n738 B.n73 163.367
R1132 B.n734 B.n73 163.367
R1133 B.n734 B.n733 163.367
R1134 B.n733 B.n732 163.367
R1135 B.n732 B.n75 163.367
R1136 B.n728 B.n75 163.367
R1137 B.n728 B.n727 163.367
R1138 B.n727 B.n726 163.367
R1139 B.n726 B.n77 163.367
R1140 B.n722 B.n77 163.367
R1141 B.n722 B.n721 163.367
R1142 B.n721 B.n720 163.367
R1143 B.n720 B.n79 163.367
R1144 B.n716 B.n79 163.367
R1145 B.n716 B.n715 163.367
R1146 B.n715 B.n714 163.367
R1147 B.n714 B.n81 163.367
R1148 B.n710 B.n81 163.367
R1149 B.n710 B.n709 163.367
R1150 B.n709 B.n708 163.367
R1151 B.n708 B.n83 163.367
R1152 B.n704 B.n83 163.367
R1153 B.n704 B.n703 163.367
R1154 B.n703 B.n702 163.367
R1155 B.n702 B.n85 163.367
R1156 B.n698 B.n85 163.367
R1157 B.n698 B.n697 163.367
R1158 B.n697 B.n696 163.367
R1159 B.n696 B.n87 163.367
R1160 B.n692 B.n87 163.367
R1161 B.n692 B.n691 163.367
R1162 B.n691 B.n690 163.367
R1163 B.n690 B.n89 163.367
R1164 B.n686 B.n89 163.367
R1165 B.n686 B.n685 163.367
R1166 B.n685 B.n684 163.367
R1167 B.n684 B.n91 163.367
R1168 B.n680 B.n91 163.367
R1169 B.n680 B.n679 163.367
R1170 B.n679 B.n678 163.367
R1171 B.n678 B.n93 163.367
R1172 B.n674 B.n93 163.367
R1173 B.n674 B.n673 163.367
R1174 B.n673 B.n672 163.367
R1175 B.n672 B.n95 163.367
R1176 B.n668 B.n95 163.367
R1177 B.n668 B.n667 163.367
R1178 B.n667 B.n666 163.367
R1179 B.n666 B.n97 163.367
R1180 B.n662 B.n97 163.367
R1181 B.n178 B.t8 160.981
R1182 B.n64 B.t1 160.981
R1183 B.n186 B.t11 160.956
R1184 B.n58 B.t4 160.956
R1185 B.n179 B.t7 108.617
R1186 B.n65 B.t2 108.617
R1187 B.n187 B.t10 108.591
R1188 B.n59 B.t5 108.591
R1189 B.n180 B.n179 59.5399
R1190 B.n407 B.n187 59.5399
R1191 B.n771 B.n59 59.5399
R1192 B.n66 B.n65 59.5399
R1193 B.n179 B.n178 52.3641
R1194 B.n187 B.n186 52.3641
R1195 B.n59 B.n58 52.3641
R1196 B.n65 B.n64 52.3641
R1197 B.n867 B.n26 30.4395
R1198 B.n515 B.n146 30.4395
R1199 B.n311 B.n218 30.4395
R1200 B.n663 B.n98 30.4395
R1201 B B.n939 18.0485
R1202 B.n863 B.n26 10.6151
R1203 B.n863 B.n862 10.6151
R1204 B.n862 B.n861 10.6151
R1205 B.n861 B.n28 10.6151
R1206 B.n857 B.n28 10.6151
R1207 B.n857 B.n856 10.6151
R1208 B.n856 B.n855 10.6151
R1209 B.n855 B.n30 10.6151
R1210 B.n851 B.n30 10.6151
R1211 B.n851 B.n850 10.6151
R1212 B.n850 B.n849 10.6151
R1213 B.n849 B.n32 10.6151
R1214 B.n845 B.n32 10.6151
R1215 B.n845 B.n844 10.6151
R1216 B.n844 B.n843 10.6151
R1217 B.n843 B.n34 10.6151
R1218 B.n839 B.n34 10.6151
R1219 B.n839 B.n838 10.6151
R1220 B.n838 B.n837 10.6151
R1221 B.n837 B.n36 10.6151
R1222 B.n833 B.n36 10.6151
R1223 B.n833 B.n832 10.6151
R1224 B.n832 B.n831 10.6151
R1225 B.n831 B.n38 10.6151
R1226 B.n827 B.n38 10.6151
R1227 B.n827 B.n826 10.6151
R1228 B.n826 B.n825 10.6151
R1229 B.n825 B.n40 10.6151
R1230 B.n821 B.n40 10.6151
R1231 B.n821 B.n820 10.6151
R1232 B.n820 B.n819 10.6151
R1233 B.n819 B.n42 10.6151
R1234 B.n815 B.n42 10.6151
R1235 B.n815 B.n814 10.6151
R1236 B.n814 B.n813 10.6151
R1237 B.n813 B.n44 10.6151
R1238 B.n809 B.n44 10.6151
R1239 B.n809 B.n808 10.6151
R1240 B.n808 B.n807 10.6151
R1241 B.n807 B.n46 10.6151
R1242 B.n803 B.n46 10.6151
R1243 B.n803 B.n802 10.6151
R1244 B.n802 B.n801 10.6151
R1245 B.n801 B.n48 10.6151
R1246 B.n797 B.n48 10.6151
R1247 B.n797 B.n796 10.6151
R1248 B.n796 B.n795 10.6151
R1249 B.n795 B.n50 10.6151
R1250 B.n791 B.n50 10.6151
R1251 B.n791 B.n790 10.6151
R1252 B.n790 B.n789 10.6151
R1253 B.n789 B.n52 10.6151
R1254 B.n785 B.n52 10.6151
R1255 B.n785 B.n784 10.6151
R1256 B.n784 B.n783 10.6151
R1257 B.n783 B.n54 10.6151
R1258 B.n779 B.n54 10.6151
R1259 B.n779 B.n778 10.6151
R1260 B.n778 B.n777 10.6151
R1261 B.n777 B.n56 10.6151
R1262 B.n773 B.n56 10.6151
R1263 B.n773 B.n772 10.6151
R1264 B.n770 B.n60 10.6151
R1265 B.n766 B.n60 10.6151
R1266 B.n766 B.n765 10.6151
R1267 B.n765 B.n764 10.6151
R1268 B.n764 B.n62 10.6151
R1269 B.n760 B.n62 10.6151
R1270 B.n760 B.n759 10.6151
R1271 B.n759 B.n758 10.6151
R1272 B.n755 B.n754 10.6151
R1273 B.n754 B.n753 10.6151
R1274 B.n753 B.n68 10.6151
R1275 B.n749 B.n68 10.6151
R1276 B.n749 B.n748 10.6151
R1277 B.n748 B.n747 10.6151
R1278 B.n747 B.n70 10.6151
R1279 B.n743 B.n70 10.6151
R1280 B.n743 B.n742 10.6151
R1281 B.n742 B.n741 10.6151
R1282 B.n741 B.n72 10.6151
R1283 B.n737 B.n72 10.6151
R1284 B.n737 B.n736 10.6151
R1285 B.n736 B.n735 10.6151
R1286 B.n735 B.n74 10.6151
R1287 B.n731 B.n74 10.6151
R1288 B.n731 B.n730 10.6151
R1289 B.n730 B.n729 10.6151
R1290 B.n729 B.n76 10.6151
R1291 B.n725 B.n76 10.6151
R1292 B.n725 B.n724 10.6151
R1293 B.n724 B.n723 10.6151
R1294 B.n723 B.n78 10.6151
R1295 B.n719 B.n78 10.6151
R1296 B.n719 B.n718 10.6151
R1297 B.n718 B.n717 10.6151
R1298 B.n717 B.n80 10.6151
R1299 B.n713 B.n80 10.6151
R1300 B.n713 B.n712 10.6151
R1301 B.n712 B.n711 10.6151
R1302 B.n711 B.n82 10.6151
R1303 B.n707 B.n82 10.6151
R1304 B.n707 B.n706 10.6151
R1305 B.n706 B.n705 10.6151
R1306 B.n705 B.n84 10.6151
R1307 B.n701 B.n84 10.6151
R1308 B.n701 B.n700 10.6151
R1309 B.n700 B.n699 10.6151
R1310 B.n699 B.n86 10.6151
R1311 B.n695 B.n86 10.6151
R1312 B.n695 B.n694 10.6151
R1313 B.n694 B.n693 10.6151
R1314 B.n693 B.n88 10.6151
R1315 B.n689 B.n88 10.6151
R1316 B.n689 B.n688 10.6151
R1317 B.n688 B.n687 10.6151
R1318 B.n687 B.n90 10.6151
R1319 B.n683 B.n90 10.6151
R1320 B.n683 B.n682 10.6151
R1321 B.n682 B.n681 10.6151
R1322 B.n681 B.n92 10.6151
R1323 B.n677 B.n92 10.6151
R1324 B.n677 B.n676 10.6151
R1325 B.n676 B.n675 10.6151
R1326 B.n675 B.n94 10.6151
R1327 B.n671 B.n94 10.6151
R1328 B.n671 B.n670 10.6151
R1329 B.n670 B.n669 10.6151
R1330 B.n669 B.n96 10.6151
R1331 B.n665 B.n96 10.6151
R1332 B.n665 B.n664 10.6151
R1333 B.n664 B.n663 10.6151
R1334 B.n519 B.n146 10.6151
R1335 B.n520 B.n519 10.6151
R1336 B.n521 B.n520 10.6151
R1337 B.n521 B.n144 10.6151
R1338 B.n525 B.n144 10.6151
R1339 B.n526 B.n525 10.6151
R1340 B.n527 B.n526 10.6151
R1341 B.n527 B.n142 10.6151
R1342 B.n531 B.n142 10.6151
R1343 B.n532 B.n531 10.6151
R1344 B.n533 B.n532 10.6151
R1345 B.n533 B.n140 10.6151
R1346 B.n537 B.n140 10.6151
R1347 B.n538 B.n537 10.6151
R1348 B.n539 B.n538 10.6151
R1349 B.n539 B.n138 10.6151
R1350 B.n543 B.n138 10.6151
R1351 B.n544 B.n543 10.6151
R1352 B.n545 B.n544 10.6151
R1353 B.n545 B.n136 10.6151
R1354 B.n549 B.n136 10.6151
R1355 B.n550 B.n549 10.6151
R1356 B.n551 B.n550 10.6151
R1357 B.n551 B.n134 10.6151
R1358 B.n555 B.n134 10.6151
R1359 B.n556 B.n555 10.6151
R1360 B.n557 B.n556 10.6151
R1361 B.n557 B.n132 10.6151
R1362 B.n561 B.n132 10.6151
R1363 B.n562 B.n561 10.6151
R1364 B.n563 B.n562 10.6151
R1365 B.n563 B.n130 10.6151
R1366 B.n567 B.n130 10.6151
R1367 B.n568 B.n567 10.6151
R1368 B.n569 B.n568 10.6151
R1369 B.n569 B.n128 10.6151
R1370 B.n573 B.n128 10.6151
R1371 B.n574 B.n573 10.6151
R1372 B.n575 B.n574 10.6151
R1373 B.n575 B.n126 10.6151
R1374 B.n579 B.n126 10.6151
R1375 B.n580 B.n579 10.6151
R1376 B.n581 B.n580 10.6151
R1377 B.n581 B.n124 10.6151
R1378 B.n585 B.n124 10.6151
R1379 B.n586 B.n585 10.6151
R1380 B.n587 B.n586 10.6151
R1381 B.n587 B.n122 10.6151
R1382 B.n591 B.n122 10.6151
R1383 B.n592 B.n591 10.6151
R1384 B.n593 B.n592 10.6151
R1385 B.n593 B.n120 10.6151
R1386 B.n597 B.n120 10.6151
R1387 B.n598 B.n597 10.6151
R1388 B.n599 B.n598 10.6151
R1389 B.n599 B.n118 10.6151
R1390 B.n603 B.n118 10.6151
R1391 B.n604 B.n603 10.6151
R1392 B.n605 B.n604 10.6151
R1393 B.n605 B.n116 10.6151
R1394 B.n609 B.n116 10.6151
R1395 B.n610 B.n609 10.6151
R1396 B.n611 B.n610 10.6151
R1397 B.n611 B.n114 10.6151
R1398 B.n615 B.n114 10.6151
R1399 B.n616 B.n615 10.6151
R1400 B.n617 B.n616 10.6151
R1401 B.n617 B.n112 10.6151
R1402 B.n621 B.n112 10.6151
R1403 B.n622 B.n621 10.6151
R1404 B.n623 B.n622 10.6151
R1405 B.n623 B.n110 10.6151
R1406 B.n627 B.n110 10.6151
R1407 B.n628 B.n627 10.6151
R1408 B.n629 B.n628 10.6151
R1409 B.n629 B.n108 10.6151
R1410 B.n633 B.n108 10.6151
R1411 B.n634 B.n633 10.6151
R1412 B.n635 B.n634 10.6151
R1413 B.n635 B.n106 10.6151
R1414 B.n639 B.n106 10.6151
R1415 B.n640 B.n639 10.6151
R1416 B.n641 B.n640 10.6151
R1417 B.n641 B.n104 10.6151
R1418 B.n645 B.n104 10.6151
R1419 B.n646 B.n645 10.6151
R1420 B.n647 B.n646 10.6151
R1421 B.n647 B.n102 10.6151
R1422 B.n651 B.n102 10.6151
R1423 B.n652 B.n651 10.6151
R1424 B.n653 B.n652 10.6151
R1425 B.n653 B.n100 10.6151
R1426 B.n657 B.n100 10.6151
R1427 B.n658 B.n657 10.6151
R1428 B.n659 B.n658 10.6151
R1429 B.n659 B.n98 10.6151
R1430 B.n315 B.n218 10.6151
R1431 B.n316 B.n315 10.6151
R1432 B.n317 B.n316 10.6151
R1433 B.n317 B.n216 10.6151
R1434 B.n321 B.n216 10.6151
R1435 B.n322 B.n321 10.6151
R1436 B.n323 B.n322 10.6151
R1437 B.n323 B.n214 10.6151
R1438 B.n327 B.n214 10.6151
R1439 B.n328 B.n327 10.6151
R1440 B.n329 B.n328 10.6151
R1441 B.n329 B.n212 10.6151
R1442 B.n333 B.n212 10.6151
R1443 B.n334 B.n333 10.6151
R1444 B.n335 B.n334 10.6151
R1445 B.n335 B.n210 10.6151
R1446 B.n339 B.n210 10.6151
R1447 B.n340 B.n339 10.6151
R1448 B.n341 B.n340 10.6151
R1449 B.n341 B.n208 10.6151
R1450 B.n345 B.n208 10.6151
R1451 B.n346 B.n345 10.6151
R1452 B.n347 B.n346 10.6151
R1453 B.n347 B.n206 10.6151
R1454 B.n351 B.n206 10.6151
R1455 B.n352 B.n351 10.6151
R1456 B.n353 B.n352 10.6151
R1457 B.n353 B.n204 10.6151
R1458 B.n357 B.n204 10.6151
R1459 B.n358 B.n357 10.6151
R1460 B.n359 B.n358 10.6151
R1461 B.n359 B.n202 10.6151
R1462 B.n363 B.n202 10.6151
R1463 B.n364 B.n363 10.6151
R1464 B.n365 B.n364 10.6151
R1465 B.n365 B.n200 10.6151
R1466 B.n369 B.n200 10.6151
R1467 B.n370 B.n369 10.6151
R1468 B.n371 B.n370 10.6151
R1469 B.n371 B.n198 10.6151
R1470 B.n375 B.n198 10.6151
R1471 B.n376 B.n375 10.6151
R1472 B.n377 B.n376 10.6151
R1473 B.n377 B.n196 10.6151
R1474 B.n381 B.n196 10.6151
R1475 B.n382 B.n381 10.6151
R1476 B.n383 B.n382 10.6151
R1477 B.n383 B.n194 10.6151
R1478 B.n387 B.n194 10.6151
R1479 B.n388 B.n387 10.6151
R1480 B.n389 B.n388 10.6151
R1481 B.n389 B.n192 10.6151
R1482 B.n393 B.n192 10.6151
R1483 B.n394 B.n393 10.6151
R1484 B.n395 B.n394 10.6151
R1485 B.n395 B.n190 10.6151
R1486 B.n399 B.n190 10.6151
R1487 B.n400 B.n399 10.6151
R1488 B.n401 B.n400 10.6151
R1489 B.n401 B.n188 10.6151
R1490 B.n405 B.n188 10.6151
R1491 B.n406 B.n405 10.6151
R1492 B.n408 B.n184 10.6151
R1493 B.n412 B.n184 10.6151
R1494 B.n413 B.n412 10.6151
R1495 B.n414 B.n413 10.6151
R1496 B.n414 B.n182 10.6151
R1497 B.n418 B.n182 10.6151
R1498 B.n419 B.n418 10.6151
R1499 B.n420 B.n419 10.6151
R1500 B.n424 B.n423 10.6151
R1501 B.n425 B.n424 10.6151
R1502 B.n425 B.n176 10.6151
R1503 B.n429 B.n176 10.6151
R1504 B.n430 B.n429 10.6151
R1505 B.n431 B.n430 10.6151
R1506 B.n431 B.n174 10.6151
R1507 B.n435 B.n174 10.6151
R1508 B.n436 B.n435 10.6151
R1509 B.n437 B.n436 10.6151
R1510 B.n437 B.n172 10.6151
R1511 B.n441 B.n172 10.6151
R1512 B.n442 B.n441 10.6151
R1513 B.n443 B.n442 10.6151
R1514 B.n443 B.n170 10.6151
R1515 B.n447 B.n170 10.6151
R1516 B.n448 B.n447 10.6151
R1517 B.n449 B.n448 10.6151
R1518 B.n449 B.n168 10.6151
R1519 B.n453 B.n168 10.6151
R1520 B.n454 B.n453 10.6151
R1521 B.n455 B.n454 10.6151
R1522 B.n455 B.n166 10.6151
R1523 B.n459 B.n166 10.6151
R1524 B.n460 B.n459 10.6151
R1525 B.n461 B.n460 10.6151
R1526 B.n461 B.n164 10.6151
R1527 B.n465 B.n164 10.6151
R1528 B.n466 B.n465 10.6151
R1529 B.n467 B.n466 10.6151
R1530 B.n467 B.n162 10.6151
R1531 B.n471 B.n162 10.6151
R1532 B.n472 B.n471 10.6151
R1533 B.n473 B.n472 10.6151
R1534 B.n473 B.n160 10.6151
R1535 B.n477 B.n160 10.6151
R1536 B.n478 B.n477 10.6151
R1537 B.n479 B.n478 10.6151
R1538 B.n479 B.n158 10.6151
R1539 B.n483 B.n158 10.6151
R1540 B.n484 B.n483 10.6151
R1541 B.n485 B.n484 10.6151
R1542 B.n485 B.n156 10.6151
R1543 B.n489 B.n156 10.6151
R1544 B.n490 B.n489 10.6151
R1545 B.n491 B.n490 10.6151
R1546 B.n491 B.n154 10.6151
R1547 B.n495 B.n154 10.6151
R1548 B.n496 B.n495 10.6151
R1549 B.n497 B.n496 10.6151
R1550 B.n497 B.n152 10.6151
R1551 B.n501 B.n152 10.6151
R1552 B.n502 B.n501 10.6151
R1553 B.n503 B.n502 10.6151
R1554 B.n503 B.n150 10.6151
R1555 B.n507 B.n150 10.6151
R1556 B.n508 B.n507 10.6151
R1557 B.n509 B.n508 10.6151
R1558 B.n509 B.n148 10.6151
R1559 B.n513 B.n148 10.6151
R1560 B.n514 B.n513 10.6151
R1561 B.n515 B.n514 10.6151
R1562 B.n311 B.n310 10.6151
R1563 B.n310 B.n309 10.6151
R1564 B.n309 B.n220 10.6151
R1565 B.n305 B.n220 10.6151
R1566 B.n305 B.n304 10.6151
R1567 B.n304 B.n303 10.6151
R1568 B.n303 B.n222 10.6151
R1569 B.n299 B.n222 10.6151
R1570 B.n299 B.n298 10.6151
R1571 B.n298 B.n297 10.6151
R1572 B.n297 B.n224 10.6151
R1573 B.n293 B.n224 10.6151
R1574 B.n293 B.n292 10.6151
R1575 B.n292 B.n291 10.6151
R1576 B.n291 B.n226 10.6151
R1577 B.n287 B.n226 10.6151
R1578 B.n287 B.n286 10.6151
R1579 B.n286 B.n285 10.6151
R1580 B.n285 B.n228 10.6151
R1581 B.n281 B.n228 10.6151
R1582 B.n281 B.n280 10.6151
R1583 B.n280 B.n279 10.6151
R1584 B.n279 B.n230 10.6151
R1585 B.n275 B.n230 10.6151
R1586 B.n275 B.n274 10.6151
R1587 B.n274 B.n273 10.6151
R1588 B.n273 B.n232 10.6151
R1589 B.n269 B.n232 10.6151
R1590 B.n269 B.n268 10.6151
R1591 B.n268 B.n267 10.6151
R1592 B.n267 B.n234 10.6151
R1593 B.n263 B.n234 10.6151
R1594 B.n263 B.n262 10.6151
R1595 B.n262 B.n261 10.6151
R1596 B.n261 B.n236 10.6151
R1597 B.n257 B.n236 10.6151
R1598 B.n257 B.n256 10.6151
R1599 B.n256 B.n255 10.6151
R1600 B.n255 B.n238 10.6151
R1601 B.n251 B.n238 10.6151
R1602 B.n251 B.n250 10.6151
R1603 B.n250 B.n249 10.6151
R1604 B.n249 B.n240 10.6151
R1605 B.n245 B.n240 10.6151
R1606 B.n245 B.n244 10.6151
R1607 B.n244 B.n243 10.6151
R1608 B.n243 B.n0 10.6151
R1609 B.n935 B.n1 10.6151
R1610 B.n935 B.n934 10.6151
R1611 B.n934 B.n933 10.6151
R1612 B.n933 B.n4 10.6151
R1613 B.n929 B.n4 10.6151
R1614 B.n929 B.n928 10.6151
R1615 B.n928 B.n927 10.6151
R1616 B.n927 B.n6 10.6151
R1617 B.n923 B.n6 10.6151
R1618 B.n923 B.n922 10.6151
R1619 B.n922 B.n921 10.6151
R1620 B.n921 B.n8 10.6151
R1621 B.n917 B.n8 10.6151
R1622 B.n917 B.n916 10.6151
R1623 B.n916 B.n915 10.6151
R1624 B.n915 B.n10 10.6151
R1625 B.n911 B.n10 10.6151
R1626 B.n911 B.n910 10.6151
R1627 B.n910 B.n909 10.6151
R1628 B.n909 B.n12 10.6151
R1629 B.n905 B.n12 10.6151
R1630 B.n905 B.n904 10.6151
R1631 B.n904 B.n903 10.6151
R1632 B.n903 B.n14 10.6151
R1633 B.n899 B.n14 10.6151
R1634 B.n899 B.n898 10.6151
R1635 B.n898 B.n897 10.6151
R1636 B.n897 B.n16 10.6151
R1637 B.n893 B.n16 10.6151
R1638 B.n893 B.n892 10.6151
R1639 B.n892 B.n891 10.6151
R1640 B.n891 B.n18 10.6151
R1641 B.n887 B.n18 10.6151
R1642 B.n887 B.n886 10.6151
R1643 B.n886 B.n885 10.6151
R1644 B.n885 B.n20 10.6151
R1645 B.n881 B.n20 10.6151
R1646 B.n881 B.n880 10.6151
R1647 B.n880 B.n879 10.6151
R1648 B.n879 B.n22 10.6151
R1649 B.n875 B.n22 10.6151
R1650 B.n875 B.n874 10.6151
R1651 B.n874 B.n873 10.6151
R1652 B.n873 B.n24 10.6151
R1653 B.n869 B.n24 10.6151
R1654 B.n869 B.n868 10.6151
R1655 B.n868 B.n867 10.6151
R1656 B.n771 B.n770 6.5566
R1657 B.n758 B.n66 6.5566
R1658 B.n408 B.n407 6.5566
R1659 B.n420 B.n180 6.5566
R1660 B.n772 B.n771 4.05904
R1661 B.n755 B.n66 4.05904
R1662 B.n407 B.n406 4.05904
R1663 B.n423 B.n180 4.05904
R1664 B.n939 B.n0 2.81026
R1665 B.n939 B.n1 2.81026
C0 B VDD1 1.77366f
C1 VDD2 w_n3670_n4802# 2.17275f
C2 VDD2 VP 0.49487f
C3 B VN 1.25593f
C4 VDD1 VTAIL 10.589901f
C5 VN VTAIL 13.369201f
C6 B VTAIL 7.19526f
C7 VP w_n3670_n4802# 8.01346f
C8 VDD2 VDD1 1.65542f
C9 VDD2 VN 13.3697f
C10 VDD2 B 1.86245f
C11 VDD2 VTAIL 10.642799f
C12 VDD1 w_n3670_n4802# 2.06769f
C13 VP VDD1 13.712299f
C14 VN w_n3670_n4802# 7.537701f
C15 VN VP 8.70837f
C16 B w_n3670_n4802# 11.7739f
C17 B VP 2.05225f
C18 w_n3670_n4802# VTAIL 5.82224f
C19 VP VTAIL 13.3833f
C20 VN VDD1 0.150986f
C21 VDD2 VSUBS 1.979317f
C22 VDD1 VSUBS 2.58202f
C23 VTAIL VSUBS 1.627493f
C24 VN VSUBS 6.76701f
C25 VP VSUBS 3.614995f
C26 B VSUBS 5.34881f
C27 w_n3670_n4802# VSUBS 0.215312p
C28 B.n0 VSUBS 0.004311f
C29 B.n1 VSUBS 0.004311f
C30 B.n2 VSUBS 0.006818f
C31 B.n3 VSUBS 0.006818f
C32 B.n4 VSUBS 0.006818f
C33 B.n5 VSUBS 0.006818f
C34 B.n6 VSUBS 0.006818f
C35 B.n7 VSUBS 0.006818f
C36 B.n8 VSUBS 0.006818f
C37 B.n9 VSUBS 0.006818f
C38 B.n10 VSUBS 0.006818f
C39 B.n11 VSUBS 0.006818f
C40 B.n12 VSUBS 0.006818f
C41 B.n13 VSUBS 0.006818f
C42 B.n14 VSUBS 0.006818f
C43 B.n15 VSUBS 0.006818f
C44 B.n16 VSUBS 0.006818f
C45 B.n17 VSUBS 0.006818f
C46 B.n18 VSUBS 0.006818f
C47 B.n19 VSUBS 0.006818f
C48 B.n20 VSUBS 0.006818f
C49 B.n21 VSUBS 0.006818f
C50 B.n22 VSUBS 0.006818f
C51 B.n23 VSUBS 0.006818f
C52 B.n24 VSUBS 0.006818f
C53 B.n25 VSUBS 0.006818f
C54 B.n26 VSUBS 0.015524f
C55 B.n27 VSUBS 0.006818f
C56 B.n28 VSUBS 0.006818f
C57 B.n29 VSUBS 0.006818f
C58 B.n30 VSUBS 0.006818f
C59 B.n31 VSUBS 0.006818f
C60 B.n32 VSUBS 0.006818f
C61 B.n33 VSUBS 0.006818f
C62 B.n34 VSUBS 0.006818f
C63 B.n35 VSUBS 0.006818f
C64 B.n36 VSUBS 0.006818f
C65 B.n37 VSUBS 0.006818f
C66 B.n38 VSUBS 0.006818f
C67 B.n39 VSUBS 0.006818f
C68 B.n40 VSUBS 0.006818f
C69 B.n41 VSUBS 0.006818f
C70 B.n42 VSUBS 0.006818f
C71 B.n43 VSUBS 0.006818f
C72 B.n44 VSUBS 0.006818f
C73 B.n45 VSUBS 0.006818f
C74 B.n46 VSUBS 0.006818f
C75 B.n47 VSUBS 0.006818f
C76 B.n48 VSUBS 0.006818f
C77 B.n49 VSUBS 0.006818f
C78 B.n50 VSUBS 0.006818f
C79 B.n51 VSUBS 0.006818f
C80 B.n52 VSUBS 0.006818f
C81 B.n53 VSUBS 0.006818f
C82 B.n54 VSUBS 0.006818f
C83 B.n55 VSUBS 0.006818f
C84 B.n56 VSUBS 0.006818f
C85 B.n57 VSUBS 0.006818f
C86 B.t5 VSUBS 0.633012f
C87 B.t4 VSUBS 0.65241f
C88 B.t3 VSUBS 1.94077f
C89 B.n58 VSUBS 0.348603f
C90 B.n59 VSUBS 0.069352f
C91 B.n60 VSUBS 0.006818f
C92 B.n61 VSUBS 0.006818f
C93 B.n62 VSUBS 0.006818f
C94 B.n63 VSUBS 0.006818f
C95 B.t2 VSUBS 0.632986f
C96 B.t1 VSUBS 0.65239f
C97 B.t0 VSUBS 1.94077f
C98 B.n64 VSUBS 0.348624f
C99 B.n65 VSUBS 0.069378f
C100 B.n66 VSUBS 0.015796f
C101 B.n67 VSUBS 0.006818f
C102 B.n68 VSUBS 0.006818f
C103 B.n69 VSUBS 0.006818f
C104 B.n70 VSUBS 0.006818f
C105 B.n71 VSUBS 0.006818f
C106 B.n72 VSUBS 0.006818f
C107 B.n73 VSUBS 0.006818f
C108 B.n74 VSUBS 0.006818f
C109 B.n75 VSUBS 0.006818f
C110 B.n76 VSUBS 0.006818f
C111 B.n77 VSUBS 0.006818f
C112 B.n78 VSUBS 0.006818f
C113 B.n79 VSUBS 0.006818f
C114 B.n80 VSUBS 0.006818f
C115 B.n81 VSUBS 0.006818f
C116 B.n82 VSUBS 0.006818f
C117 B.n83 VSUBS 0.006818f
C118 B.n84 VSUBS 0.006818f
C119 B.n85 VSUBS 0.006818f
C120 B.n86 VSUBS 0.006818f
C121 B.n87 VSUBS 0.006818f
C122 B.n88 VSUBS 0.006818f
C123 B.n89 VSUBS 0.006818f
C124 B.n90 VSUBS 0.006818f
C125 B.n91 VSUBS 0.006818f
C126 B.n92 VSUBS 0.006818f
C127 B.n93 VSUBS 0.006818f
C128 B.n94 VSUBS 0.006818f
C129 B.n95 VSUBS 0.006818f
C130 B.n96 VSUBS 0.006818f
C131 B.n97 VSUBS 0.006818f
C132 B.n98 VSUBS 0.015819f
C133 B.n99 VSUBS 0.006818f
C134 B.n100 VSUBS 0.006818f
C135 B.n101 VSUBS 0.006818f
C136 B.n102 VSUBS 0.006818f
C137 B.n103 VSUBS 0.006818f
C138 B.n104 VSUBS 0.006818f
C139 B.n105 VSUBS 0.006818f
C140 B.n106 VSUBS 0.006818f
C141 B.n107 VSUBS 0.006818f
C142 B.n108 VSUBS 0.006818f
C143 B.n109 VSUBS 0.006818f
C144 B.n110 VSUBS 0.006818f
C145 B.n111 VSUBS 0.006818f
C146 B.n112 VSUBS 0.006818f
C147 B.n113 VSUBS 0.006818f
C148 B.n114 VSUBS 0.006818f
C149 B.n115 VSUBS 0.006818f
C150 B.n116 VSUBS 0.006818f
C151 B.n117 VSUBS 0.006818f
C152 B.n118 VSUBS 0.006818f
C153 B.n119 VSUBS 0.006818f
C154 B.n120 VSUBS 0.006818f
C155 B.n121 VSUBS 0.006818f
C156 B.n122 VSUBS 0.006818f
C157 B.n123 VSUBS 0.006818f
C158 B.n124 VSUBS 0.006818f
C159 B.n125 VSUBS 0.006818f
C160 B.n126 VSUBS 0.006818f
C161 B.n127 VSUBS 0.006818f
C162 B.n128 VSUBS 0.006818f
C163 B.n129 VSUBS 0.006818f
C164 B.n130 VSUBS 0.006818f
C165 B.n131 VSUBS 0.006818f
C166 B.n132 VSUBS 0.006818f
C167 B.n133 VSUBS 0.006818f
C168 B.n134 VSUBS 0.006818f
C169 B.n135 VSUBS 0.006818f
C170 B.n136 VSUBS 0.006818f
C171 B.n137 VSUBS 0.006818f
C172 B.n138 VSUBS 0.006818f
C173 B.n139 VSUBS 0.006818f
C174 B.n140 VSUBS 0.006818f
C175 B.n141 VSUBS 0.006818f
C176 B.n142 VSUBS 0.006818f
C177 B.n143 VSUBS 0.006818f
C178 B.n144 VSUBS 0.006818f
C179 B.n145 VSUBS 0.006818f
C180 B.n146 VSUBS 0.014955f
C181 B.n147 VSUBS 0.006818f
C182 B.n148 VSUBS 0.006818f
C183 B.n149 VSUBS 0.006818f
C184 B.n150 VSUBS 0.006818f
C185 B.n151 VSUBS 0.006818f
C186 B.n152 VSUBS 0.006818f
C187 B.n153 VSUBS 0.006818f
C188 B.n154 VSUBS 0.006818f
C189 B.n155 VSUBS 0.006818f
C190 B.n156 VSUBS 0.006818f
C191 B.n157 VSUBS 0.006818f
C192 B.n158 VSUBS 0.006818f
C193 B.n159 VSUBS 0.006818f
C194 B.n160 VSUBS 0.006818f
C195 B.n161 VSUBS 0.006818f
C196 B.n162 VSUBS 0.006818f
C197 B.n163 VSUBS 0.006818f
C198 B.n164 VSUBS 0.006818f
C199 B.n165 VSUBS 0.006818f
C200 B.n166 VSUBS 0.006818f
C201 B.n167 VSUBS 0.006818f
C202 B.n168 VSUBS 0.006818f
C203 B.n169 VSUBS 0.006818f
C204 B.n170 VSUBS 0.006818f
C205 B.n171 VSUBS 0.006818f
C206 B.n172 VSUBS 0.006818f
C207 B.n173 VSUBS 0.006818f
C208 B.n174 VSUBS 0.006818f
C209 B.n175 VSUBS 0.006818f
C210 B.n176 VSUBS 0.006818f
C211 B.n177 VSUBS 0.006818f
C212 B.t7 VSUBS 0.632986f
C213 B.t8 VSUBS 0.65239f
C214 B.t6 VSUBS 1.94077f
C215 B.n178 VSUBS 0.348624f
C216 B.n179 VSUBS 0.069378f
C217 B.n180 VSUBS 0.015796f
C218 B.n181 VSUBS 0.006818f
C219 B.n182 VSUBS 0.006818f
C220 B.n183 VSUBS 0.006818f
C221 B.n184 VSUBS 0.006818f
C222 B.n185 VSUBS 0.006818f
C223 B.t10 VSUBS 0.633012f
C224 B.t11 VSUBS 0.65241f
C225 B.t9 VSUBS 1.94077f
C226 B.n186 VSUBS 0.348603f
C227 B.n187 VSUBS 0.069352f
C228 B.n188 VSUBS 0.006818f
C229 B.n189 VSUBS 0.006818f
C230 B.n190 VSUBS 0.006818f
C231 B.n191 VSUBS 0.006818f
C232 B.n192 VSUBS 0.006818f
C233 B.n193 VSUBS 0.006818f
C234 B.n194 VSUBS 0.006818f
C235 B.n195 VSUBS 0.006818f
C236 B.n196 VSUBS 0.006818f
C237 B.n197 VSUBS 0.006818f
C238 B.n198 VSUBS 0.006818f
C239 B.n199 VSUBS 0.006818f
C240 B.n200 VSUBS 0.006818f
C241 B.n201 VSUBS 0.006818f
C242 B.n202 VSUBS 0.006818f
C243 B.n203 VSUBS 0.006818f
C244 B.n204 VSUBS 0.006818f
C245 B.n205 VSUBS 0.006818f
C246 B.n206 VSUBS 0.006818f
C247 B.n207 VSUBS 0.006818f
C248 B.n208 VSUBS 0.006818f
C249 B.n209 VSUBS 0.006818f
C250 B.n210 VSUBS 0.006818f
C251 B.n211 VSUBS 0.006818f
C252 B.n212 VSUBS 0.006818f
C253 B.n213 VSUBS 0.006818f
C254 B.n214 VSUBS 0.006818f
C255 B.n215 VSUBS 0.006818f
C256 B.n216 VSUBS 0.006818f
C257 B.n217 VSUBS 0.006818f
C258 B.n218 VSUBS 0.015524f
C259 B.n219 VSUBS 0.006818f
C260 B.n220 VSUBS 0.006818f
C261 B.n221 VSUBS 0.006818f
C262 B.n222 VSUBS 0.006818f
C263 B.n223 VSUBS 0.006818f
C264 B.n224 VSUBS 0.006818f
C265 B.n225 VSUBS 0.006818f
C266 B.n226 VSUBS 0.006818f
C267 B.n227 VSUBS 0.006818f
C268 B.n228 VSUBS 0.006818f
C269 B.n229 VSUBS 0.006818f
C270 B.n230 VSUBS 0.006818f
C271 B.n231 VSUBS 0.006818f
C272 B.n232 VSUBS 0.006818f
C273 B.n233 VSUBS 0.006818f
C274 B.n234 VSUBS 0.006818f
C275 B.n235 VSUBS 0.006818f
C276 B.n236 VSUBS 0.006818f
C277 B.n237 VSUBS 0.006818f
C278 B.n238 VSUBS 0.006818f
C279 B.n239 VSUBS 0.006818f
C280 B.n240 VSUBS 0.006818f
C281 B.n241 VSUBS 0.006818f
C282 B.n242 VSUBS 0.006818f
C283 B.n243 VSUBS 0.006818f
C284 B.n244 VSUBS 0.006818f
C285 B.n245 VSUBS 0.006818f
C286 B.n246 VSUBS 0.006818f
C287 B.n247 VSUBS 0.006818f
C288 B.n248 VSUBS 0.006818f
C289 B.n249 VSUBS 0.006818f
C290 B.n250 VSUBS 0.006818f
C291 B.n251 VSUBS 0.006818f
C292 B.n252 VSUBS 0.006818f
C293 B.n253 VSUBS 0.006818f
C294 B.n254 VSUBS 0.006818f
C295 B.n255 VSUBS 0.006818f
C296 B.n256 VSUBS 0.006818f
C297 B.n257 VSUBS 0.006818f
C298 B.n258 VSUBS 0.006818f
C299 B.n259 VSUBS 0.006818f
C300 B.n260 VSUBS 0.006818f
C301 B.n261 VSUBS 0.006818f
C302 B.n262 VSUBS 0.006818f
C303 B.n263 VSUBS 0.006818f
C304 B.n264 VSUBS 0.006818f
C305 B.n265 VSUBS 0.006818f
C306 B.n266 VSUBS 0.006818f
C307 B.n267 VSUBS 0.006818f
C308 B.n268 VSUBS 0.006818f
C309 B.n269 VSUBS 0.006818f
C310 B.n270 VSUBS 0.006818f
C311 B.n271 VSUBS 0.006818f
C312 B.n272 VSUBS 0.006818f
C313 B.n273 VSUBS 0.006818f
C314 B.n274 VSUBS 0.006818f
C315 B.n275 VSUBS 0.006818f
C316 B.n276 VSUBS 0.006818f
C317 B.n277 VSUBS 0.006818f
C318 B.n278 VSUBS 0.006818f
C319 B.n279 VSUBS 0.006818f
C320 B.n280 VSUBS 0.006818f
C321 B.n281 VSUBS 0.006818f
C322 B.n282 VSUBS 0.006818f
C323 B.n283 VSUBS 0.006818f
C324 B.n284 VSUBS 0.006818f
C325 B.n285 VSUBS 0.006818f
C326 B.n286 VSUBS 0.006818f
C327 B.n287 VSUBS 0.006818f
C328 B.n288 VSUBS 0.006818f
C329 B.n289 VSUBS 0.006818f
C330 B.n290 VSUBS 0.006818f
C331 B.n291 VSUBS 0.006818f
C332 B.n292 VSUBS 0.006818f
C333 B.n293 VSUBS 0.006818f
C334 B.n294 VSUBS 0.006818f
C335 B.n295 VSUBS 0.006818f
C336 B.n296 VSUBS 0.006818f
C337 B.n297 VSUBS 0.006818f
C338 B.n298 VSUBS 0.006818f
C339 B.n299 VSUBS 0.006818f
C340 B.n300 VSUBS 0.006818f
C341 B.n301 VSUBS 0.006818f
C342 B.n302 VSUBS 0.006818f
C343 B.n303 VSUBS 0.006818f
C344 B.n304 VSUBS 0.006818f
C345 B.n305 VSUBS 0.006818f
C346 B.n306 VSUBS 0.006818f
C347 B.n307 VSUBS 0.006818f
C348 B.n308 VSUBS 0.006818f
C349 B.n309 VSUBS 0.006818f
C350 B.n310 VSUBS 0.006818f
C351 B.n311 VSUBS 0.014955f
C352 B.n312 VSUBS 0.014955f
C353 B.n313 VSUBS 0.015524f
C354 B.n314 VSUBS 0.006818f
C355 B.n315 VSUBS 0.006818f
C356 B.n316 VSUBS 0.006818f
C357 B.n317 VSUBS 0.006818f
C358 B.n318 VSUBS 0.006818f
C359 B.n319 VSUBS 0.006818f
C360 B.n320 VSUBS 0.006818f
C361 B.n321 VSUBS 0.006818f
C362 B.n322 VSUBS 0.006818f
C363 B.n323 VSUBS 0.006818f
C364 B.n324 VSUBS 0.006818f
C365 B.n325 VSUBS 0.006818f
C366 B.n326 VSUBS 0.006818f
C367 B.n327 VSUBS 0.006818f
C368 B.n328 VSUBS 0.006818f
C369 B.n329 VSUBS 0.006818f
C370 B.n330 VSUBS 0.006818f
C371 B.n331 VSUBS 0.006818f
C372 B.n332 VSUBS 0.006818f
C373 B.n333 VSUBS 0.006818f
C374 B.n334 VSUBS 0.006818f
C375 B.n335 VSUBS 0.006818f
C376 B.n336 VSUBS 0.006818f
C377 B.n337 VSUBS 0.006818f
C378 B.n338 VSUBS 0.006818f
C379 B.n339 VSUBS 0.006818f
C380 B.n340 VSUBS 0.006818f
C381 B.n341 VSUBS 0.006818f
C382 B.n342 VSUBS 0.006818f
C383 B.n343 VSUBS 0.006818f
C384 B.n344 VSUBS 0.006818f
C385 B.n345 VSUBS 0.006818f
C386 B.n346 VSUBS 0.006818f
C387 B.n347 VSUBS 0.006818f
C388 B.n348 VSUBS 0.006818f
C389 B.n349 VSUBS 0.006818f
C390 B.n350 VSUBS 0.006818f
C391 B.n351 VSUBS 0.006818f
C392 B.n352 VSUBS 0.006818f
C393 B.n353 VSUBS 0.006818f
C394 B.n354 VSUBS 0.006818f
C395 B.n355 VSUBS 0.006818f
C396 B.n356 VSUBS 0.006818f
C397 B.n357 VSUBS 0.006818f
C398 B.n358 VSUBS 0.006818f
C399 B.n359 VSUBS 0.006818f
C400 B.n360 VSUBS 0.006818f
C401 B.n361 VSUBS 0.006818f
C402 B.n362 VSUBS 0.006818f
C403 B.n363 VSUBS 0.006818f
C404 B.n364 VSUBS 0.006818f
C405 B.n365 VSUBS 0.006818f
C406 B.n366 VSUBS 0.006818f
C407 B.n367 VSUBS 0.006818f
C408 B.n368 VSUBS 0.006818f
C409 B.n369 VSUBS 0.006818f
C410 B.n370 VSUBS 0.006818f
C411 B.n371 VSUBS 0.006818f
C412 B.n372 VSUBS 0.006818f
C413 B.n373 VSUBS 0.006818f
C414 B.n374 VSUBS 0.006818f
C415 B.n375 VSUBS 0.006818f
C416 B.n376 VSUBS 0.006818f
C417 B.n377 VSUBS 0.006818f
C418 B.n378 VSUBS 0.006818f
C419 B.n379 VSUBS 0.006818f
C420 B.n380 VSUBS 0.006818f
C421 B.n381 VSUBS 0.006818f
C422 B.n382 VSUBS 0.006818f
C423 B.n383 VSUBS 0.006818f
C424 B.n384 VSUBS 0.006818f
C425 B.n385 VSUBS 0.006818f
C426 B.n386 VSUBS 0.006818f
C427 B.n387 VSUBS 0.006818f
C428 B.n388 VSUBS 0.006818f
C429 B.n389 VSUBS 0.006818f
C430 B.n390 VSUBS 0.006818f
C431 B.n391 VSUBS 0.006818f
C432 B.n392 VSUBS 0.006818f
C433 B.n393 VSUBS 0.006818f
C434 B.n394 VSUBS 0.006818f
C435 B.n395 VSUBS 0.006818f
C436 B.n396 VSUBS 0.006818f
C437 B.n397 VSUBS 0.006818f
C438 B.n398 VSUBS 0.006818f
C439 B.n399 VSUBS 0.006818f
C440 B.n400 VSUBS 0.006818f
C441 B.n401 VSUBS 0.006818f
C442 B.n402 VSUBS 0.006818f
C443 B.n403 VSUBS 0.006818f
C444 B.n404 VSUBS 0.006818f
C445 B.n405 VSUBS 0.006818f
C446 B.n406 VSUBS 0.004712f
C447 B.n407 VSUBS 0.015796f
C448 B.n408 VSUBS 0.005514f
C449 B.n409 VSUBS 0.006818f
C450 B.n410 VSUBS 0.006818f
C451 B.n411 VSUBS 0.006818f
C452 B.n412 VSUBS 0.006818f
C453 B.n413 VSUBS 0.006818f
C454 B.n414 VSUBS 0.006818f
C455 B.n415 VSUBS 0.006818f
C456 B.n416 VSUBS 0.006818f
C457 B.n417 VSUBS 0.006818f
C458 B.n418 VSUBS 0.006818f
C459 B.n419 VSUBS 0.006818f
C460 B.n420 VSUBS 0.005514f
C461 B.n421 VSUBS 0.006818f
C462 B.n422 VSUBS 0.006818f
C463 B.n423 VSUBS 0.004712f
C464 B.n424 VSUBS 0.006818f
C465 B.n425 VSUBS 0.006818f
C466 B.n426 VSUBS 0.006818f
C467 B.n427 VSUBS 0.006818f
C468 B.n428 VSUBS 0.006818f
C469 B.n429 VSUBS 0.006818f
C470 B.n430 VSUBS 0.006818f
C471 B.n431 VSUBS 0.006818f
C472 B.n432 VSUBS 0.006818f
C473 B.n433 VSUBS 0.006818f
C474 B.n434 VSUBS 0.006818f
C475 B.n435 VSUBS 0.006818f
C476 B.n436 VSUBS 0.006818f
C477 B.n437 VSUBS 0.006818f
C478 B.n438 VSUBS 0.006818f
C479 B.n439 VSUBS 0.006818f
C480 B.n440 VSUBS 0.006818f
C481 B.n441 VSUBS 0.006818f
C482 B.n442 VSUBS 0.006818f
C483 B.n443 VSUBS 0.006818f
C484 B.n444 VSUBS 0.006818f
C485 B.n445 VSUBS 0.006818f
C486 B.n446 VSUBS 0.006818f
C487 B.n447 VSUBS 0.006818f
C488 B.n448 VSUBS 0.006818f
C489 B.n449 VSUBS 0.006818f
C490 B.n450 VSUBS 0.006818f
C491 B.n451 VSUBS 0.006818f
C492 B.n452 VSUBS 0.006818f
C493 B.n453 VSUBS 0.006818f
C494 B.n454 VSUBS 0.006818f
C495 B.n455 VSUBS 0.006818f
C496 B.n456 VSUBS 0.006818f
C497 B.n457 VSUBS 0.006818f
C498 B.n458 VSUBS 0.006818f
C499 B.n459 VSUBS 0.006818f
C500 B.n460 VSUBS 0.006818f
C501 B.n461 VSUBS 0.006818f
C502 B.n462 VSUBS 0.006818f
C503 B.n463 VSUBS 0.006818f
C504 B.n464 VSUBS 0.006818f
C505 B.n465 VSUBS 0.006818f
C506 B.n466 VSUBS 0.006818f
C507 B.n467 VSUBS 0.006818f
C508 B.n468 VSUBS 0.006818f
C509 B.n469 VSUBS 0.006818f
C510 B.n470 VSUBS 0.006818f
C511 B.n471 VSUBS 0.006818f
C512 B.n472 VSUBS 0.006818f
C513 B.n473 VSUBS 0.006818f
C514 B.n474 VSUBS 0.006818f
C515 B.n475 VSUBS 0.006818f
C516 B.n476 VSUBS 0.006818f
C517 B.n477 VSUBS 0.006818f
C518 B.n478 VSUBS 0.006818f
C519 B.n479 VSUBS 0.006818f
C520 B.n480 VSUBS 0.006818f
C521 B.n481 VSUBS 0.006818f
C522 B.n482 VSUBS 0.006818f
C523 B.n483 VSUBS 0.006818f
C524 B.n484 VSUBS 0.006818f
C525 B.n485 VSUBS 0.006818f
C526 B.n486 VSUBS 0.006818f
C527 B.n487 VSUBS 0.006818f
C528 B.n488 VSUBS 0.006818f
C529 B.n489 VSUBS 0.006818f
C530 B.n490 VSUBS 0.006818f
C531 B.n491 VSUBS 0.006818f
C532 B.n492 VSUBS 0.006818f
C533 B.n493 VSUBS 0.006818f
C534 B.n494 VSUBS 0.006818f
C535 B.n495 VSUBS 0.006818f
C536 B.n496 VSUBS 0.006818f
C537 B.n497 VSUBS 0.006818f
C538 B.n498 VSUBS 0.006818f
C539 B.n499 VSUBS 0.006818f
C540 B.n500 VSUBS 0.006818f
C541 B.n501 VSUBS 0.006818f
C542 B.n502 VSUBS 0.006818f
C543 B.n503 VSUBS 0.006818f
C544 B.n504 VSUBS 0.006818f
C545 B.n505 VSUBS 0.006818f
C546 B.n506 VSUBS 0.006818f
C547 B.n507 VSUBS 0.006818f
C548 B.n508 VSUBS 0.006818f
C549 B.n509 VSUBS 0.006818f
C550 B.n510 VSUBS 0.006818f
C551 B.n511 VSUBS 0.006818f
C552 B.n512 VSUBS 0.006818f
C553 B.n513 VSUBS 0.006818f
C554 B.n514 VSUBS 0.006818f
C555 B.n515 VSUBS 0.015524f
C556 B.n516 VSUBS 0.015524f
C557 B.n517 VSUBS 0.014955f
C558 B.n518 VSUBS 0.006818f
C559 B.n519 VSUBS 0.006818f
C560 B.n520 VSUBS 0.006818f
C561 B.n521 VSUBS 0.006818f
C562 B.n522 VSUBS 0.006818f
C563 B.n523 VSUBS 0.006818f
C564 B.n524 VSUBS 0.006818f
C565 B.n525 VSUBS 0.006818f
C566 B.n526 VSUBS 0.006818f
C567 B.n527 VSUBS 0.006818f
C568 B.n528 VSUBS 0.006818f
C569 B.n529 VSUBS 0.006818f
C570 B.n530 VSUBS 0.006818f
C571 B.n531 VSUBS 0.006818f
C572 B.n532 VSUBS 0.006818f
C573 B.n533 VSUBS 0.006818f
C574 B.n534 VSUBS 0.006818f
C575 B.n535 VSUBS 0.006818f
C576 B.n536 VSUBS 0.006818f
C577 B.n537 VSUBS 0.006818f
C578 B.n538 VSUBS 0.006818f
C579 B.n539 VSUBS 0.006818f
C580 B.n540 VSUBS 0.006818f
C581 B.n541 VSUBS 0.006818f
C582 B.n542 VSUBS 0.006818f
C583 B.n543 VSUBS 0.006818f
C584 B.n544 VSUBS 0.006818f
C585 B.n545 VSUBS 0.006818f
C586 B.n546 VSUBS 0.006818f
C587 B.n547 VSUBS 0.006818f
C588 B.n548 VSUBS 0.006818f
C589 B.n549 VSUBS 0.006818f
C590 B.n550 VSUBS 0.006818f
C591 B.n551 VSUBS 0.006818f
C592 B.n552 VSUBS 0.006818f
C593 B.n553 VSUBS 0.006818f
C594 B.n554 VSUBS 0.006818f
C595 B.n555 VSUBS 0.006818f
C596 B.n556 VSUBS 0.006818f
C597 B.n557 VSUBS 0.006818f
C598 B.n558 VSUBS 0.006818f
C599 B.n559 VSUBS 0.006818f
C600 B.n560 VSUBS 0.006818f
C601 B.n561 VSUBS 0.006818f
C602 B.n562 VSUBS 0.006818f
C603 B.n563 VSUBS 0.006818f
C604 B.n564 VSUBS 0.006818f
C605 B.n565 VSUBS 0.006818f
C606 B.n566 VSUBS 0.006818f
C607 B.n567 VSUBS 0.006818f
C608 B.n568 VSUBS 0.006818f
C609 B.n569 VSUBS 0.006818f
C610 B.n570 VSUBS 0.006818f
C611 B.n571 VSUBS 0.006818f
C612 B.n572 VSUBS 0.006818f
C613 B.n573 VSUBS 0.006818f
C614 B.n574 VSUBS 0.006818f
C615 B.n575 VSUBS 0.006818f
C616 B.n576 VSUBS 0.006818f
C617 B.n577 VSUBS 0.006818f
C618 B.n578 VSUBS 0.006818f
C619 B.n579 VSUBS 0.006818f
C620 B.n580 VSUBS 0.006818f
C621 B.n581 VSUBS 0.006818f
C622 B.n582 VSUBS 0.006818f
C623 B.n583 VSUBS 0.006818f
C624 B.n584 VSUBS 0.006818f
C625 B.n585 VSUBS 0.006818f
C626 B.n586 VSUBS 0.006818f
C627 B.n587 VSUBS 0.006818f
C628 B.n588 VSUBS 0.006818f
C629 B.n589 VSUBS 0.006818f
C630 B.n590 VSUBS 0.006818f
C631 B.n591 VSUBS 0.006818f
C632 B.n592 VSUBS 0.006818f
C633 B.n593 VSUBS 0.006818f
C634 B.n594 VSUBS 0.006818f
C635 B.n595 VSUBS 0.006818f
C636 B.n596 VSUBS 0.006818f
C637 B.n597 VSUBS 0.006818f
C638 B.n598 VSUBS 0.006818f
C639 B.n599 VSUBS 0.006818f
C640 B.n600 VSUBS 0.006818f
C641 B.n601 VSUBS 0.006818f
C642 B.n602 VSUBS 0.006818f
C643 B.n603 VSUBS 0.006818f
C644 B.n604 VSUBS 0.006818f
C645 B.n605 VSUBS 0.006818f
C646 B.n606 VSUBS 0.006818f
C647 B.n607 VSUBS 0.006818f
C648 B.n608 VSUBS 0.006818f
C649 B.n609 VSUBS 0.006818f
C650 B.n610 VSUBS 0.006818f
C651 B.n611 VSUBS 0.006818f
C652 B.n612 VSUBS 0.006818f
C653 B.n613 VSUBS 0.006818f
C654 B.n614 VSUBS 0.006818f
C655 B.n615 VSUBS 0.006818f
C656 B.n616 VSUBS 0.006818f
C657 B.n617 VSUBS 0.006818f
C658 B.n618 VSUBS 0.006818f
C659 B.n619 VSUBS 0.006818f
C660 B.n620 VSUBS 0.006818f
C661 B.n621 VSUBS 0.006818f
C662 B.n622 VSUBS 0.006818f
C663 B.n623 VSUBS 0.006818f
C664 B.n624 VSUBS 0.006818f
C665 B.n625 VSUBS 0.006818f
C666 B.n626 VSUBS 0.006818f
C667 B.n627 VSUBS 0.006818f
C668 B.n628 VSUBS 0.006818f
C669 B.n629 VSUBS 0.006818f
C670 B.n630 VSUBS 0.006818f
C671 B.n631 VSUBS 0.006818f
C672 B.n632 VSUBS 0.006818f
C673 B.n633 VSUBS 0.006818f
C674 B.n634 VSUBS 0.006818f
C675 B.n635 VSUBS 0.006818f
C676 B.n636 VSUBS 0.006818f
C677 B.n637 VSUBS 0.006818f
C678 B.n638 VSUBS 0.006818f
C679 B.n639 VSUBS 0.006818f
C680 B.n640 VSUBS 0.006818f
C681 B.n641 VSUBS 0.006818f
C682 B.n642 VSUBS 0.006818f
C683 B.n643 VSUBS 0.006818f
C684 B.n644 VSUBS 0.006818f
C685 B.n645 VSUBS 0.006818f
C686 B.n646 VSUBS 0.006818f
C687 B.n647 VSUBS 0.006818f
C688 B.n648 VSUBS 0.006818f
C689 B.n649 VSUBS 0.006818f
C690 B.n650 VSUBS 0.006818f
C691 B.n651 VSUBS 0.006818f
C692 B.n652 VSUBS 0.006818f
C693 B.n653 VSUBS 0.006818f
C694 B.n654 VSUBS 0.006818f
C695 B.n655 VSUBS 0.006818f
C696 B.n656 VSUBS 0.006818f
C697 B.n657 VSUBS 0.006818f
C698 B.n658 VSUBS 0.006818f
C699 B.n659 VSUBS 0.006818f
C700 B.n660 VSUBS 0.006818f
C701 B.n661 VSUBS 0.014955f
C702 B.n662 VSUBS 0.015524f
C703 B.n663 VSUBS 0.01466f
C704 B.n664 VSUBS 0.006818f
C705 B.n665 VSUBS 0.006818f
C706 B.n666 VSUBS 0.006818f
C707 B.n667 VSUBS 0.006818f
C708 B.n668 VSUBS 0.006818f
C709 B.n669 VSUBS 0.006818f
C710 B.n670 VSUBS 0.006818f
C711 B.n671 VSUBS 0.006818f
C712 B.n672 VSUBS 0.006818f
C713 B.n673 VSUBS 0.006818f
C714 B.n674 VSUBS 0.006818f
C715 B.n675 VSUBS 0.006818f
C716 B.n676 VSUBS 0.006818f
C717 B.n677 VSUBS 0.006818f
C718 B.n678 VSUBS 0.006818f
C719 B.n679 VSUBS 0.006818f
C720 B.n680 VSUBS 0.006818f
C721 B.n681 VSUBS 0.006818f
C722 B.n682 VSUBS 0.006818f
C723 B.n683 VSUBS 0.006818f
C724 B.n684 VSUBS 0.006818f
C725 B.n685 VSUBS 0.006818f
C726 B.n686 VSUBS 0.006818f
C727 B.n687 VSUBS 0.006818f
C728 B.n688 VSUBS 0.006818f
C729 B.n689 VSUBS 0.006818f
C730 B.n690 VSUBS 0.006818f
C731 B.n691 VSUBS 0.006818f
C732 B.n692 VSUBS 0.006818f
C733 B.n693 VSUBS 0.006818f
C734 B.n694 VSUBS 0.006818f
C735 B.n695 VSUBS 0.006818f
C736 B.n696 VSUBS 0.006818f
C737 B.n697 VSUBS 0.006818f
C738 B.n698 VSUBS 0.006818f
C739 B.n699 VSUBS 0.006818f
C740 B.n700 VSUBS 0.006818f
C741 B.n701 VSUBS 0.006818f
C742 B.n702 VSUBS 0.006818f
C743 B.n703 VSUBS 0.006818f
C744 B.n704 VSUBS 0.006818f
C745 B.n705 VSUBS 0.006818f
C746 B.n706 VSUBS 0.006818f
C747 B.n707 VSUBS 0.006818f
C748 B.n708 VSUBS 0.006818f
C749 B.n709 VSUBS 0.006818f
C750 B.n710 VSUBS 0.006818f
C751 B.n711 VSUBS 0.006818f
C752 B.n712 VSUBS 0.006818f
C753 B.n713 VSUBS 0.006818f
C754 B.n714 VSUBS 0.006818f
C755 B.n715 VSUBS 0.006818f
C756 B.n716 VSUBS 0.006818f
C757 B.n717 VSUBS 0.006818f
C758 B.n718 VSUBS 0.006818f
C759 B.n719 VSUBS 0.006818f
C760 B.n720 VSUBS 0.006818f
C761 B.n721 VSUBS 0.006818f
C762 B.n722 VSUBS 0.006818f
C763 B.n723 VSUBS 0.006818f
C764 B.n724 VSUBS 0.006818f
C765 B.n725 VSUBS 0.006818f
C766 B.n726 VSUBS 0.006818f
C767 B.n727 VSUBS 0.006818f
C768 B.n728 VSUBS 0.006818f
C769 B.n729 VSUBS 0.006818f
C770 B.n730 VSUBS 0.006818f
C771 B.n731 VSUBS 0.006818f
C772 B.n732 VSUBS 0.006818f
C773 B.n733 VSUBS 0.006818f
C774 B.n734 VSUBS 0.006818f
C775 B.n735 VSUBS 0.006818f
C776 B.n736 VSUBS 0.006818f
C777 B.n737 VSUBS 0.006818f
C778 B.n738 VSUBS 0.006818f
C779 B.n739 VSUBS 0.006818f
C780 B.n740 VSUBS 0.006818f
C781 B.n741 VSUBS 0.006818f
C782 B.n742 VSUBS 0.006818f
C783 B.n743 VSUBS 0.006818f
C784 B.n744 VSUBS 0.006818f
C785 B.n745 VSUBS 0.006818f
C786 B.n746 VSUBS 0.006818f
C787 B.n747 VSUBS 0.006818f
C788 B.n748 VSUBS 0.006818f
C789 B.n749 VSUBS 0.006818f
C790 B.n750 VSUBS 0.006818f
C791 B.n751 VSUBS 0.006818f
C792 B.n752 VSUBS 0.006818f
C793 B.n753 VSUBS 0.006818f
C794 B.n754 VSUBS 0.006818f
C795 B.n755 VSUBS 0.004712f
C796 B.n756 VSUBS 0.006818f
C797 B.n757 VSUBS 0.006818f
C798 B.n758 VSUBS 0.005514f
C799 B.n759 VSUBS 0.006818f
C800 B.n760 VSUBS 0.006818f
C801 B.n761 VSUBS 0.006818f
C802 B.n762 VSUBS 0.006818f
C803 B.n763 VSUBS 0.006818f
C804 B.n764 VSUBS 0.006818f
C805 B.n765 VSUBS 0.006818f
C806 B.n766 VSUBS 0.006818f
C807 B.n767 VSUBS 0.006818f
C808 B.n768 VSUBS 0.006818f
C809 B.n769 VSUBS 0.006818f
C810 B.n770 VSUBS 0.005514f
C811 B.n771 VSUBS 0.015796f
C812 B.n772 VSUBS 0.004712f
C813 B.n773 VSUBS 0.006818f
C814 B.n774 VSUBS 0.006818f
C815 B.n775 VSUBS 0.006818f
C816 B.n776 VSUBS 0.006818f
C817 B.n777 VSUBS 0.006818f
C818 B.n778 VSUBS 0.006818f
C819 B.n779 VSUBS 0.006818f
C820 B.n780 VSUBS 0.006818f
C821 B.n781 VSUBS 0.006818f
C822 B.n782 VSUBS 0.006818f
C823 B.n783 VSUBS 0.006818f
C824 B.n784 VSUBS 0.006818f
C825 B.n785 VSUBS 0.006818f
C826 B.n786 VSUBS 0.006818f
C827 B.n787 VSUBS 0.006818f
C828 B.n788 VSUBS 0.006818f
C829 B.n789 VSUBS 0.006818f
C830 B.n790 VSUBS 0.006818f
C831 B.n791 VSUBS 0.006818f
C832 B.n792 VSUBS 0.006818f
C833 B.n793 VSUBS 0.006818f
C834 B.n794 VSUBS 0.006818f
C835 B.n795 VSUBS 0.006818f
C836 B.n796 VSUBS 0.006818f
C837 B.n797 VSUBS 0.006818f
C838 B.n798 VSUBS 0.006818f
C839 B.n799 VSUBS 0.006818f
C840 B.n800 VSUBS 0.006818f
C841 B.n801 VSUBS 0.006818f
C842 B.n802 VSUBS 0.006818f
C843 B.n803 VSUBS 0.006818f
C844 B.n804 VSUBS 0.006818f
C845 B.n805 VSUBS 0.006818f
C846 B.n806 VSUBS 0.006818f
C847 B.n807 VSUBS 0.006818f
C848 B.n808 VSUBS 0.006818f
C849 B.n809 VSUBS 0.006818f
C850 B.n810 VSUBS 0.006818f
C851 B.n811 VSUBS 0.006818f
C852 B.n812 VSUBS 0.006818f
C853 B.n813 VSUBS 0.006818f
C854 B.n814 VSUBS 0.006818f
C855 B.n815 VSUBS 0.006818f
C856 B.n816 VSUBS 0.006818f
C857 B.n817 VSUBS 0.006818f
C858 B.n818 VSUBS 0.006818f
C859 B.n819 VSUBS 0.006818f
C860 B.n820 VSUBS 0.006818f
C861 B.n821 VSUBS 0.006818f
C862 B.n822 VSUBS 0.006818f
C863 B.n823 VSUBS 0.006818f
C864 B.n824 VSUBS 0.006818f
C865 B.n825 VSUBS 0.006818f
C866 B.n826 VSUBS 0.006818f
C867 B.n827 VSUBS 0.006818f
C868 B.n828 VSUBS 0.006818f
C869 B.n829 VSUBS 0.006818f
C870 B.n830 VSUBS 0.006818f
C871 B.n831 VSUBS 0.006818f
C872 B.n832 VSUBS 0.006818f
C873 B.n833 VSUBS 0.006818f
C874 B.n834 VSUBS 0.006818f
C875 B.n835 VSUBS 0.006818f
C876 B.n836 VSUBS 0.006818f
C877 B.n837 VSUBS 0.006818f
C878 B.n838 VSUBS 0.006818f
C879 B.n839 VSUBS 0.006818f
C880 B.n840 VSUBS 0.006818f
C881 B.n841 VSUBS 0.006818f
C882 B.n842 VSUBS 0.006818f
C883 B.n843 VSUBS 0.006818f
C884 B.n844 VSUBS 0.006818f
C885 B.n845 VSUBS 0.006818f
C886 B.n846 VSUBS 0.006818f
C887 B.n847 VSUBS 0.006818f
C888 B.n848 VSUBS 0.006818f
C889 B.n849 VSUBS 0.006818f
C890 B.n850 VSUBS 0.006818f
C891 B.n851 VSUBS 0.006818f
C892 B.n852 VSUBS 0.006818f
C893 B.n853 VSUBS 0.006818f
C894 B.n854 VSUBS 0.006818f
C895 B.n855 VSUBS 0.006818f
C896 B.n856 VSUBS 0.006818f
C897 B.n857 VSUBS 0.006818f
C898 B.n858 VSUBS 0.006818f
C899 B.n859 VSUBS 0.006818f
C900 B.n860 VSUBS 0.006818f
C901 B.n861 VSUBS 0.006818f
C902 B.n862 VSUBS 0.006818f
C903 B.n863 VSUBS 0.006818f
C904 B.n864 VSUBS 0.006818f
C905 B.n865 VSUBS 0.015524f
C906 B.n866 VSUBS 0.014955f
C907 B.n867 VSUBS 0.014955f
C908 B.n868 VSUBS 0.006818f
C909 B.n869 VSUBS 0.006818f
C910 B.n870 VSUBS 0.006818f
C911 B.n871 VSUBS 0.006818f
C912 B.n872 VSUBS 0.006818f
C913 B.n873 VSUBS 0.006818f
C914 B.n874 VSUBS 0.006818f
C915 B.n875 VSUBS 0.006818f
C916 B.n876 VSUBS 0.006818f
C917 B.n877 VSUBS 0.006818f
C918 B.n878 VSUBS 0.006818f
C919 B.n879 VSUBS 0.006818f
C920 B.n880 VSUBS 0.006818f
C921 B.n881 VSUBS 0.006818f
C922 B.n882 VSUBS 0.006818f
C923 B.n883 VSUBS 0.006818f
C924 B.n884 VSUBS 0.006818f
C925 B.n885 VSUBS 0.006818f
C926 B.n886 VSUBS 0.006818f
C927 B.n887 VSUBS 0.006818f
C928 B.n888 VSUBS 0.006818f
C929 B.n889 VSUBS 0.006818f
C930 B.n890 VSUBS 0.006818f
C931 B.n891 VSUBS 0.006818f
C932 B.n892 VSUBS 0.006818f
C933 B.n893 VSUBS 0.006818f
C934 B.n894 VSUBS 0.006818f
C935 B.n895 VSUBS 0.006818f
C936 B.n896 VSUBS 0.006818f
C937 B.n897 VSUBS 0.006818f
C938 B.n898 VSUBS 0.006818f
C939 B.n899 VSUBS 0.006818f
C940 B.n900 VSUBS 0.006818f
C941 B.n901 VSUBS 0.006818f
C942 B.n902 VSUBS 0.006818f
C943 B.n903 VSUBS 0.006818f
C944 B.n904 VSUBS 0.006818f
C945 B.n905 VSUBS 0.006818f
C946 B.n906 VSUBS 0.006818f
C947 B.n907 VSUBS 0.006818f
C948 B.n908 VSUBS 0.006818f
C949 B.n909 VSUBS 0.006818f
C950 B.n910 VSUBS 0.006818f
C951 B.n911 VSUBS 0.006818f
C952 B.n912 VSUBS 0.006818f
C953 B.n913 VSUBS 0.006818f
C954 B.n914 VSUBS 0.006818f
C955 B.n915 VSUBS 0.006818f
C956 B.n916 VSUBS 0.006818f
C957 B.n917 VSUBS 0.006818f
C958 B.n918 VSUBS 0.006818f
C959 B.n919 VSUBS 0.006818f
C960 B.n920 VSUBS 0.006818f
C961 B.n921 VSUBS 0.006818f
C962 B.n922 VSUBS 0.006818f
C963 B.n923 VSUBS 0.006818f
C964 B.n924 VSUBS 0.006818f
C965 B.n925 VSUBS 0.006818f
C966 B.n926 VSUBS 0.006818f
C967 B.n927 VSUBS 0.006818f
C968 B.n928 VSUBS 0.006818f
C969 B.n929 VSUBS 0.006818f
C970 B.n930 VSUBS 0.006818f
C971 B.n931 VSUBS 0.006818f
C972 B.n932 VSUBS 0.006818f
C973 B.n933 VSUBS 0.006818f
C974 B.n934 VSUBS 0.006818f
C975 B.n935 VSUBS 0.006818f
C976 B.n936 VSUBS 0.006818f
C977 B.n937 VSUBS 0.006818f
C978 B.n938 VSUBS 0.006818f
C979 B.n939 VSUBS 0.015438f
C980 VDD2.t5 VSUBS 0.40363f
C981 VDD2.t1 VSUBS 0.40363f
C982 VDD2.n0 VSUBS 3.41744f
C983 VDD2.t3 VSUBS 0.40363f
C984 VDD2.t6 VSUBS 0.40363f
C985 VDD2.n1 VSUBS 3.41744f
C986 VDD2.n2 VSUBS 4.39623f
C987 VDD2.t7 VSUBS 0.40363f
C988 VDD2.t2 VSUBS 0.40363f
C989 VDD2.n3 VSUBS 3.40519f
C990 VDD2.n4 VSUBS 3.92093f
C991 VDD2.t0 VSUBS 0.40363f
C992 VDD2.t4 VSUBS 0.40363f
C993 VDD2.n5 VSUBS 3.41739f
C994 VN.n0 VSUBS 0.03589f
C995 VN.t1 VSUBS 3.40584f
C996 VN.n1 VSUBS 0.022894f
C997 VN.n2 VSUBS 0.027223f
C998 VN.t4 VSUBS 3.40584f
C999 VN.n3 VSUBS 0.050736f
C1000 VN.n4 VSUBS 0.027223f
C1001 VN.n5 VSUBS 0.030697f
C1002 VN.t2 VSUBS 3.59619f
C1003 VN.t6 VSUBS 3.40584f
C1004 VN.n6 VSUBS 1.24758f
C1005 VN.n7 VSUBS 1.23887f
C1006 VN.n8 VSUBS 0.23636f
C1007 VN.n9 VSUBS 0.027223f
C1008 VN.n10 VSUBS 0.050736f
C1009 VN.n11 VSUBS 0.03974f
C1010 VN.n12 VSUBS 0.03974f
C1011 VN.n13 VSUBS 0.027223f
C1012 VN.n14 VSUBS 0.027223f
C1013 VN.n15 VSUBS 0.027223f
C1014 VN.n16 VSUBS 0.030697f
C1015 VN.n17 VSUBS 1.18042f
C1016 VN.n18 VSUBS 0.045727f
C1017 VN.n19 VSUBS 0.052349f
C1018 VN.n20 VSUBS 0.027223f
C1019 VN.n21 VSUBS 0.027223f
C1020 VN.n22 VSUBS 0.027223f
C1021 VN.n23 VSUBS 0.054974f
C1022 VN.n24 VSUBS 0.040717f
C1023 VN.n25 VSUBS 1.27042f
C1024 VN.n26 VSUBS 0.039086f
C1025 VN.n27 VSUBS 0.03589f
C1026 VN.t0 VSUBS 3.40584f
C1027 VN.n28 VSUBS 0.022894f
C1028 VN.n29 VSUBS 0.027223f
C1029 VN.t5 VSUBS 3.40584f
C1030 VN.n30 VSUBS 0.050736f
C1031 VN.n31 VSUBS 0.027223f
C1032 VN.n32 VSUBS 0.030697f
C1033 VN.t3 VSUBS 3.59619f
C1034 VN.t7 VSUBS 3.40584f
C1035 VN.n33 VSUBS 1.24758f
C1036 VN.n34 VSUBS 1.23887f
C1037 VN.n35 VSUBS 0.23636f
C1038 VN.n36 VSUBS 0.027223f
C1039 VN.n37 VSUBS 0.050736f
C1040 VN.n38 VSUBS 0.03974f
C1041 VN.n39 VSUBS 0.03974f
C1042 VN.n40 VSUBS 0.027223f
C1043 VN.n41 VSUBS 0.027223f
C1044 VN.n42 VSUBS 0.027223f
C1045 VN.n43 VSUBS 0.030697f
C1046 VN.n44 VSUBS 1.18042f
C1047 VN.n45 VSUBS 0.045727f
C1048 VN.n46 VSUBS 0.052349f
C1049 VN.n47 VSUBS 0.027223f
C1050 VN.n48 VSUBS 0.027223f
C1051 VN.n49 VSUBS 0.027223f
C1052 VN.n50 VSUBS 0.054974f
C1053 VN.n51 VSUBS 0.040717f
C1054 VN.n52 VSUBS 1.27042f
C1055 VN.n53 VSUBS 1.75916f
C1056 VTAIL.t7 VSUBS 0.35283f
C1057 VTAIL.t6 VSUBS 0.35283f
C1058 VTAIL.n0 VSUBS 2.84541f
C1059 VTAIL.n1 VSUBS 0.718472f
C1060 VTAIL.t3 VSUBS 3.705f
C1061 VTAIL.n2 VSUBS 0.852045f
C1062 VTAIL.t8 VSUBS 3.705f
C1063 VTAIL.n3 VSUBS 0.852045f
C1064 VTAIL.t14 VSUBS 0.35283f
C1065 VTAIL.t12 VSUBS 0.35283f
C1066 VTAIL.n4 VSUBS 2.84541f
C1067 VTAIL.n5 VSUBS 0.888788f
C1068 VTAIL.t9 VSUBS 3.705f
C1069 VTAIL.n6 VSUBS 2.5481f
C1070 VTAIL.t5 VSUBS 3.70503f
C1071 VTAIL.n7 VSUBS 2.54807f
C1072 VTAIL.t1 VSUBS 0.35283f
C1073 VTAIL.t2 VSUBS 0.35283f
C1074 VTAIL.n8 VSUBS 2.84543f
C1075 VTAIL.n9 VSUBS 0.888772f
C1076 VTAIL.t4 VSUBS 3.70503f
C1077 VTAIL.n10 VSUBS 0.852011f
C1078 VTAIL.t13 VSUBS 3.70503f
C1079 VTAIL.n11 VSUBS 0.852011f
C1080 VTAIL.t10 VSUBS 0.35283f
C1081 VTAIL.t15 VSUBS 0.35283f
C1082 VTAIL.n12 VSUBS 2.84543f
C1083 VTAIL.n13 VSUBS 0.888772f
C1084 VTAIL.t11 VSUBS 3.705f
C1085 VTAIL.n14 VSUBS 2.5481f
C1086 VTAIL.t0 VSUBS 3.705f
C1087 VTAIL.n15 VSUBS 2.54373f
C1088 VDD1.t3 VSUBS 0.405189f
C1089 VDD1.t4 VSUBS 0.405189f
C1090 VDD1.n0 VSUBS 3.43205f
C1091 VDD1.t7 VSUBS 0.405189f
C1092 VDD1.t0 VSUBS 0.405189f
C1093 VDD1.n1 VSUBS 3.43064f
C1094 VDD1.t2 VSUBS 0.405189f
C1095 VDD1.t6 VSUBS 0.405189f
C1096 VDD1.n2 VSUBS 3.43064f
C1097 VDD1.n3 VSUBS 4.46873f
C1098 VDD1.t1 VSUBS 0.405189f
C1099 VDD1.t5 VSUBS 0.405189f
C1100 VDD1.n4 VSUBS 3.41832f
C1101 VDD1.n5 VSUBS 3.96935f
C1102 VP.n0 VSUBS 0.038345f
C1103 VP.t7 VSUBS 3.63878f
C1104 VP.n1 VSUBS 0.02446f
C1105 VP.n2 VSUBS 0.029084f
C1106 VP.t3 VSUBS 3.63878f
C1107 VP.n3 VSUBS 0.054206f
C1108 VP.n4 VSUBS 0.029084f
C1109 VP.n5 VSUBS 0.032797f
C1110 VP.n6 VSUBS 0.029084f
C1111 VP.n7 VSUBS 0.058734f
C1112 VP.n8 VSUBS 0.038345f
C1113 VP.t4 VSUBS 3.63878f
C1114 VP.n9 VSUBS 0.02446f
C1115 VP.n10 VSUBS 0.029084f
C1116 VP.t0 VSUBS 3.63878f
C1117 VP.n11 VSUBS 0.054206f
C1118 VP.n12 VSUBS 0.029084f
C1119 VP.n13 VSUBS 0.032797f
C1120 VP.t2 VSUBS 3.84214f
C1121 VP.t5 VSUBS 3.63878f
C1122 VP.n14 VSUBS 1.3329f
C1123 VP.n15 VSUBS 1.3236f
C1124 VP.n16 VSUBS 0.252526f
C1125 VP.n17 VSUBS 0.029084f
C1126 VP.n18 VSUBS 0.054206f
C1127 VP.n19 VSUBS 0.042458f
C1128 VP.n20 VSUBS 0.042458f
C1129 VP.n21 VSUBS 0.029084f
C1130 VP.n22 VSUBS 0.029084f
C1131 VP.n23 VSUBS 0.029084f
C1132 VP.n24 VSUBS 0.032797f
C1133 VP.n25 VSUBS 1.26115f
C1134 VP.n26 VSUBS 0.048854f
C1135 VP.n27 VSUBS 0.055929f
C1136 VP.n28 VSUBS 0.029084f
C1137 VP.n29 VSUBS 0.029084f
C1138 VP.n30 VSUBS 0.029084f
C1139 VP.n31 VSUBS 0.058734f
C1140 VP.n32 VSUBS 0.043501f
C1141 VP.n33 VSUBS 1.3573f
C1142 VP.n34 VSUBS 1.86408f
C1143 VP.n35 VSUBS 1.88299f
C1144 VP.t6 VSUBS 3.63878f
C1145 VP.n36 VSUBS 1.3573f
C1146 VP.n37 VSUBS 0.043501f
C1147 VP.n38 VSUBS 0.038345f
C1148 VP.n39 VSUBS 0.029084f
C1149 VP.n40 VSUBS 0.029084f
C1150 VP.n41 VSUBS 0.02446f
C1151 VP.n42 VSUBS 0.055929f
C1152 VP.t1 VSUBS 3.63878f
C1153 VP.n43 VSUBS 1.26115f
C1154 VP.n44 VSUBS 0.048854f
C1155 VP.n45 VSUBS 0.029084f
C1156 VP.n46 VSUBS 0.029084f
C1157 VP.n47 VSUBS 0.029084f
C1158 VP.n48 VSUBS 0.054206f
C1159 VP.n49 VSUBS 0.042458f
C1160 VP.n50 VSUBS 0.042458f
C1161 VP.n51 VSUBS 0.029084f
C1162 VP.n52 VSUBS 0.029084f
C1163 VP.n53 VSUBS 0.029084f
C1164 VP.n54 VSUBS 0.032797f
C1165 VP.n55 VSUBS 1.26115f
C1166 VP.n56 VSUBS 0.048854f
C1167 VP.n57 VSUBS 0.055929f
C1168 VP.n58 VSUBS 0.029084f
C1169 VP.n59 VSUBS 0.029084f
C1170 VP.n60 VSUBS 0.029084f
C1171 VP.n61 VSUBS 0.058734f
C1172 VP.n62 VSUBS 0.043501f
C1173 VP.n63 VSUBS 1.3573f
C1174 VP.n64 VSUBS 0.04176f
.ends

