* NGSPICE file created from diff_pair_sample_0770.ext - technology: sky130A

.subckt diff_pair_sample_0770 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VN.t0 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.8083 pd=17.35 as=2.8083 ps=17.35 w=17.02 l=3.54
X1 VTAIL.t8 VP.t0 VDD1.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=2.8083 pd=17.35 as=2.8083 ps=17.35 w=17.02 l=3.54
X2 VDD1.t8 VP.t1 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.8083 pd=17.35 as=2.8083 ps=17.35 w=17.02 l=3.54
X3 VTAIL.t6 VP.t2 VDD1.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=2.8083 pd=17.35 as=2.8083 ps=17.35 w=17.02 l=3.54
X4 VDD1.t6 VP.t3 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.8083 pd=17.35 as=6.6378 ps=34.82 w=17.02 l=3.54
X5 VDD2.t2 VN.t1 VTAIL.t17 B.t3 sky130_fd_pr__nfet_01v8 ad=6.6378 pd=34.82 as=2.8083 ps=17.35 w=17.02 l=3.54
X6 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=6.6378 pd=34.82 as=0 ps=0 w=17.02 l=3.54
X7 VDD1.t5 VP.t4 VTAIL.t19 B.t9 sky130_fd_pr__nfet_01v8 ad=2.8083 pd=17.35 as=6.6378 ps=34.82 w=17.02 l=3.54
X8 VDD1.t4 VP.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.8083 pd=17.35 as=2.8083 ps=17.35 w=17.02 l=3.54
X9 VDD2.t1 VN.t2 VTAIL.t16 B.t4 sky130_fd_pr__nfet_01v8 ad=2.8083 pd=17.35 as=2.8083 ps=17.35 w=17.02 l=3.54
X10 VTAIL.t15 VN.t3 VDD2.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=2.8083 pd=17.35 as=2.8083 ps=17.35 w=17.02 l=3.54
X11 VDD1.t3 VP.t6 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=6.6378 pd=34.82 as=2.8083 ps=17.35 w=17.02 l=3.54
X12 VDD2.t8 VN.t4 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=6.6378 pd=34.82 as=2.8083 ps=17.35 w=17.02 l=3.54
X13 VDD2.t7 VN.t5 VTAIL.t13 B.t7 sky130_fd_pr__nfet_01v8 ad=2.8083 pd=17.35 as=2.8083 ps=17.35 w=17.02 l=3.54
X14 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=6.6378 pd=34.82 as=0 ps=0 w=17.02 l=3.54
X15 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=6.6378 pd=34.82 as=0 ps=0 w=17.02 l=3.54
X16 VDD2.t6 VN.t6 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=2.8083 pd=17.35 as=6.6378 ps=34.82 w=17.02 l=3.54
X17 VDD2.t5 VN.t7 VTAIL.t11 B.t9 sky130_fd_pr__nfet_01v8 ad=2.8083 pd=17.35 as=6.6378 ps=34.82 w=17.02 l=3.54
X18 VTAIL.t10 VN.t8 VDD2.t4 B.t8 sky130_fd_pr__nfet_01v8 ad=2.8083 pd=17.35 as=2.8083 ps=17.35 w=17.02 l=3.54
X19 VTAIL.t2 VP.t7 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.8083 pd=17.35 as=2.8083 ps=17.35 w=17.02 l=3.54
X20 VTAIL.t1 VP.t8 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.8083 pd=17.35 as=2.8083 ps=17.35 w=17.02 l=3.54
X21 VTAIL.t9 VN.t9 VDD2.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=2.8083 pd=17.35 as=2.8083 ps=17.35 w=17.02 l=3.54
X22 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.6378 pd=34.82 as=0 ps=0 w=17.02 l=3.54
X23 VDD1.t0 VP.t9 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.6378 pd=34.82 as=2.8083 ps=17.35 w=17.02 l=3.54
R0 VN.n100 VN.n99 161.3
R1 VN.n98 VN.n52 161.3
R2 VN.n97 VN.n96 161.3
R3 VN.n95 VN.n53 161.3
R4 VN.n94 VN.n93 161.3
R5 VN.n92 VN.n54 161.3
R6 VN.n91 VN.n90 161.3
R7 VN.n89 VN.n55 161.3
R8 VN.n88 VN.n87 161.3
R9 VN.n86 VN.n56 161.3
R10 VN.n85 VN.n84 161.3
R11 VN.n83 VN.n58 161.3
R12 VN.n82 VN.n81 161.3
R13 VN.n80 VN.n59 161.3
R14 VN.n79 VN.n78 161.3
R15 VN.n77 VN.n60 161.3
R16 VN.n76 VN.n75 161.3
R17 VN.n74 VN.n61 161.3
R18 VN.n73 VN.n72 161.3
R19 VN.n71 VN.n62 161.3
R20 VN.n70 VN.n69 161.3
R21 VN.n68 VN.n63 161.3
R22 VN.n67 VN.n66 161.3
R23 VN.n49 VN.n48 161.3
R24 VN.n47 VN.n1 161.3
R25 VN.n46 VN.n45 161.3
R26 VN.n44 VN.n2 161.3
R27 VN.n43 VN.n42 161.3
R28 VN.n41 VN.n3 161.3
R29 VN.n40 VN.n39 161.3
R30 VN.n38 VN.n4 161.3
R31 VN.n37 VN.n36 161.3
R32 VN.n34 VN.n5 161.3
R33 VN.n33 VN.n32 161.3
R34 VN.n31 VN.n6 161.3
R35 VN.n30 VN.n29 161.3
R36 VN.n28 VN.n7 161.3
R37 VN.n27 VN.n26 161.3
R38 VN.n25 VN.n8 161.3
R39 VN.n24 VN.n23 161.3
R40 VN.n22 VN.n9 161.3
R41 VN.n21 VN.n20 161.3
R42 VN.n19 VN.n10 161.3
R43 VN.n18 VN.n17 161.3
R44 VN.n16 VN.n11 161.3
R45 VN.n15 VN.n14 161.3
R46 VN.n65 VN.t6 149.602
R47 VN.n13 VN.t4 149.602
R48 VN.n8 VN.t2 115.871
R49 VN.n12 VN.t0 115.871
R50 VN.n35 VN.t9 115.871
R51 VN.n0 VN.t7 115.871
R52 VN.n60 VN.t5 115.871
R53 VN.n64 VN.t8 115.871
R54 VN.n57 VN.t3 115.871
R55 VN.n51 VN.t1 115.871
R56 VN.n50 VN.n0 78.4415
R57 VN.n101 VN.n51 78.4415
R58 VN VN.n101 62.3201
R59 VN.n13 VN.n12 56.696
R60 VN.n65 VN.n64 56.696
R61 VN.n42 VN.n2 56.5617
R62 VN.n93 VN.n53 56.5617
R63 VN.n21 VN.n10 46.874
R64 VN.n29 VN.n6 46.874
R65 VN.n73 VN.n62 46.874
R66 VN.n81 VN.n58 46.874
R67 VN.n17 VN.n10 34.28
R68 VN.n33 VN.n6 34.28
R69 VN.n69 VN.n62 34.28
R70 VN.n85 VN.n58 34.28
R71 VN.n16 VN.n15 24.5923
R72 VN.n17 VN.n16 24.5923
R73 VN.n22 VN.n21 24.5923
R74 VN.n23 VN.n22 24.5923
R75 VN.n23 VN.n8 24.5923
R76 VN.n27 VN.n8 24.5923
R77 VN.n28 VN.n27 24.5923
R78 VN.n29 VN.n28 24.5923
R79 VN.n34 VN.n33 24.5923
R80 VN.n36 VN.n34 24.5923
R81 VN.n40 VN.n4 24.5923
R82 VN.n41 VN.n40 24.5923
R83 VN.n42 VN.n41 24.5923
R84 VN.n46 VN.n2 24.5923
R85 VN.n47 VN.n46 24.5923
R86 VN.n48 VN.n47 24.5923
R87 VN.n69 VN.n68 24.5923
R88 VN.n68 VN.n67 24.5923
R89 VN.n81 VN.n80 24.5923
R90 VN.n80 VN.n79 24.5923
R91 VN.n79 VN.n60 24.5923
R92 VN.n75 VN.n60 24.5923
R93 VN.n75 VN.n74 24.5923
R94 VN.n74 VN.n73 24.5923
R95 VN.n93 VN.n92 24.5923
R96 VN.n92 VN.n91 24.5923
R97 VN.n91 VN.n55 24.5923
R98 VN.n87 VN.n86 24.5923
R99 VN.n86 VN.n85 24.5923
R100 VN.n99 VN.n98 24.5923
R101 VN.n98 VN.n97 24.5923
R102 VN.n97 VN.n53 24.5923
R103 VN.n15 VN.n12 18.1985
R104 VN.n36 VN.n35 18.1985
R105 VN.n67 VN.n64 18.1985
R106 VN.n87 VN.n57 18.1985
R107 VN.n48 VN.n0 11.8046
R108 VN.n99 VN.n51 11.8046
R109 VN.n35 VN.n4 6.39438
R110 VN.n57 VN.n55 6.39438
R111 VN.n66 VN.n65 3.08737
R112 VN.n14 VN.n13 3.08737
R113 VN.n101 VN.n100 0.354861
R114 VN.n50 VN.n49 0.354861
R115 VN VN.n50 0.267071
R116 VN.n100 VN.n52 0.189894
R117 VN.n96 VN.n52 0.189894
R118 VN.n96 VN.n95 0.189894
R119 VN.n95 VN.n94 0.189894
R120 VN.n94 VN.n54 0.189894
R121 VN.n90 VN.n54 0.189894
R122 VN.n90 VN.n89 0.189894
R123 VN.n89 VN.n88 0.189894
R124 VN.n88 VN.n56 0.189894
R125 VN.n84 VN.n56 0.189894
R126 VN.n84 VN.n83 0.189894
R127 VN.n83 VN.n82 0.189894
R128 VN.n82 VN.n59 0.189894
R129 VN.n78 VN.n59 0.189894
R130 VN.n78 VN.n77 0.189894
R131 VN.n77 VN.n76 0.189894
R132 VN.n76 VN.n61 0.189894
R133 VN.n72 VN.n61 0.189894
R134 VN.n72 VN.n71 0.189894
R135 VN.n71 VN.n70 0.189894
R136 VN.n70 VN.n63 0.189894
R137 VN.n66 VN.n63 0.189894
R138 VN.n14 VN.n11 0.189894
R139 VN.n18 VN.n11 0.189894
R140 VN.n19 VN.n18 0.189894
R141 VN.n20 VN.n19 0.189894
R142 VN.n20 VN.n9 0.189894
R143 VN.n24 VN.n9 0.189894
R144 VN.n25 VN.n24 0.189894
R145 VN.n26 VN.n25 0.189894
R146 VN.n26 VN.n7 0.189894
R147 VN.n30 VN.n7 0.189894
R148 VN.n31 VN.n30 0.189894
R149 VN.n32 VN.n31 0.189894
R150 VN.n32 VN.n5 0.189894
R151 VN.n37 VN.n5 0.189894
R152 VN.n38 VN.n37 0.189894
R153 VN.n39 VN.n38 0.189894
R154 VN.n39 VN.n3 0.189894
R155 VN.n43 VN.n3 0.189894
R156 VN.n44 VN.n43 0.189894
R157 VN.n45 VN.n44 0.189894
R158 VN.n45 VN.n1 0.189894
R159 VN.n49 VN.n1 0.189894
R160 VDD2.n1 VDD2.t8 68.7814
R161 VDD2.n3 VDD2.n2 66.7286
R162 VDD2 VDD2.n7 66.7258
R163 VDD2.n4 VDD2.t2 65.4462
R164 VDD2.n6 VDD2.n5 64.2828
R165 VDD2.n1 VDD2.n0 64.2818
R166 VDD2.n4 VDD2.n3 54.2347
R167 VDD2.n6 VDD2.n4 3.33671
R168 VDD2.n7 VDD2.t4 1.16384
R169 VDD2.n7 VDD2.t6 1.16384
R170 VDD2.n5 VDD2.t9 1.16384
R171 VDD2.n5 VDD2.t7 1.16384
R172 VDD2.n2 VDD2.t0 1.16384
R173 VDD2.n2 VDD2.t5 1.16384
R174 VDD2.n0 VDD2.t3 1.16384
R175 VDD2.n0 VDD2.t1 1.16384
R176 VDD2 VDD2.n6 0.892741
R177 VDD2.n3 VDD2.n1 0.779206
R178 VTAIL.n11 VTAIL.t12 48.7674
R179 VTAIL.n17 VTAIL.t11 48.7664
R180 VTAIL.n2 VTAIL.t5 48.7664
R181 VTAIL.n16 VTAIL.t19 48.7664
R182 VTAIL.n15 VTAIL.n14 47.6041
R183 VTAIL.n13 VTAIL.n12 47.6041
R184 VTAIL.n10 VTAIL.n9 47.6041
R185 VTAIL.n8 VTAIL.n7 47.6041
R186 VTAIL.n19 VTAIL.n18 47.603
R187 VTAIL.n1 VTAIL.n0 47.603
R188 VTAIL.n4 VTAIL.n3 47.603
R189 VTAIL.n6 VTAIL.n5 47.603
R190 VTAIL.n8 VTAIL.n6 33.7117
R191 VTAIL.n17 VTAIL.n16 30.3755
R192 VTAIL.n10 VTAIL.n8 3.33671
R193 VTAIL.n11 VTAIL.n10 3.33671
R194 VTAIL.n15 VTAIL.n13 3.33671
R195 VTAIL.n16 VTAIL.n15 3.33671
R196 VTAIL.n6 VTAIL.n4 3.33671
R197 VTAIL.n4 VTAIL.n2 3.33671
R198 VTAIL.n19 VTAIL.n17 3.33671
R199 VTAIL VTAIL.n1 2.56084
R200 VTAIL.n13 VTAIL.n11 2.13843
R201 VTAIL.n2 VTAIL.n1 2.13843
R202 VTAIL.n18 VTAIL.t16 1.16384
R203 VTAIL.n18 VTAIL.t9 1.16384
R204 VTAIL.n0 VTAIL.t14 1.16384
R205 VTAIL.n0 VTAIL.t18 1.16384
R206 VTAIL.n3 VTAIL.t7 1.16384
R207 VTAIL.n3 VTAIL.t8 1.16384
R208 VTAIL.n5 VTAIL.t3 1.16384
R209 VTAIL.n5 VTAIL.t2 1.16384
R210 VTAIL.n14 VTAIL.t4 1.16384
R211 VTAIL.n14 VTAIL.t6 1.16384
R212 VTAIL.n12 VTAIL.t0 1.16384
R213 VTAIL.n12 VTAIL.t1 1.16384
R214 VTAIL.n9 VTAIL.t13 1.16384
R215 VTAIL.n9 VTAIL.t10 1.16384
R216 VTAIL.n7 VTAIL.t17 1.16384
R217 VTAIL.n7 VTAIL.t15 1.16384
R218 VTAIL VTAIL.n19 0.776362
R219 B.n1233 B.n1232 585
R220 B.n445 B.n200 585
R221 B.n444 B.n443 585
R222 B.n442 B.n441 585
R223 B.n440 B.n439 585
R224 B.n438 B.n437 585
R225 B.n436 B.n435 585
R226 B.n434 B.n433 585
R227 B.n432 B.n431 585
R228 B.n430 B.n429 585
R229 B.n428 B.n427 585
R230 B.n426 B.n425 585
R231 B.n424 B.n423 585
R232 B.n422 B.n421 585
R233 B.n420 B.n419 585
R234 B.n418 B.n417 585
R235 B.n416 B.n415 585
R236 B.n414 B.n413 585
R237 B.n412 B.n411 585
R238 B.n410 B.n409 585
R239 B.n408 B.n407 585
R240 B.n406 B.n405 585
R241 B.n404 B.n403 585
R242 B.n402 B.n401 585
R243 B.n400 B.n399 585
R244 B.n398 B.n397 585
R245 B.n396 B.n395 585
R246 B.n394 B.n393 585
R247 B.n392 B.n391 585
R248 B.n390 B.n389 585
R249 B.n388 B.n387 585
R250 B.n386 B.n385 585
R251 B.n384 B.n383 585
R252 B.n382 B.n381 585
R253 B.n380 B.n379 585
R254 B.n378 B.n377 585
R255 B.n376 B.n375 585
R256 B.n374 B.n373 585
R257 B.n372 B.n371 585
R258 B.n370 B.n369 585
R259 B.n368 B.n367 585
R260 B.n366 B.n365 585
R261 B.n364 B.n363 585
R262 B.n362 B.n361 585
R263 B.n360 B.n359 585
R264 B.n358 B.n357 585
R265 B.n356 B.n355 585
R266 B.n354 B.n353 585
R267 B.n352 B.n351 585
R268 B.n350 B.n349 585
R269 B.n348 B.n347 585
R270 B.n346 B.n345 585
R271 B.n344 B.n343 585
R272 B.n342 B.n341 585
R273 B.n340 B.n339 585
R274 B.n338 B.n337 585
R275 B.n336 B.n335 585
R276 B.n334 B.n333 585
R277 B.n332 B.n331 585
R278 B.n330 B.n329 585
R279 B.n328 B.n327 585
R280 B.n326 B.n325 585
R281 B.n324 B.n323 585
R282 B.n322 B.n321 585
R283 B.n320 B.n319 585
R284 B.n318 B.n317 585
R285 B.n316 B.n315 585
R286 B.n314 B.n313 585
R287 B.n312 B.n311 585
R288 B.n310 B.n309 585
R289 B.n308 B.n307 585
R290 B.n306 B.n305 585
R291 B.n304 B.n303 585
R292 B.n302 B.n301 585
R293 B.n300 B.n299 585
R294 B.n298 B.n297 585
R295 B.n296 B.n295 585
R296 B.n294 B.n293 585
R297 B.n292 B.n291 585
R298 B.n290 B.n289 585
R299 B.n288 B.n287 585
R300 B.n286 B.n285 585
R301 B.n284 B.n283 585
R302 B.n282 B.n281 585
R303 B.n280 B.n279 585
R304 B.n278 B.n277 585
R305 B.n276 B.n275 585
R306 B.n274 B.n273 585
R307 B.n272 B.n271 585
R308 B.n270 B.n269 585
R309 B.n268 B.n267 585
R310 B.n266 B.n265 585
R311 B.n264 B.n263 585
R312 B.n262 B.n261 585
R313 B.n260 B.n259 585
R314 B.n258 B.n257 585
R315 B.n256 B.n255 585
R316 B.n254 B.n253 585
R317 B.n252 B.n251 585
R318 B.n250 B.n249 585
R319 B.n248 B.n247 585
R320 B.n246 B.n245 585
R321 B.n244 B.n243 585
R322 B.n242 B.n241 585
R323 B.n240 B.n239 585
R324 B.n238 B.n237 585
R325 B.n236 B.n235 585
R326 B.n234 B.n233 585
R327 B.n232 B.n231 585
R328 B.n230 B.n229 585
R329 B.n228 B.n227 585
R330 B.n226 B.n225 585
R331 B.n224 B.n223 585
R332 B.n222 B.n221 585
R333 B.n220 B.n219 585
R334 B.n218 B.n217 585
R335 B.n216 B.n215 585
R336 B.n214 B.n213 585
R337 B.n212 B.n211 585
R338 B.n210 B.n209 585
R339 B.n208 B.n207 585
R340 B.n138 B.n137 585
R341 B.n1231 B.n139 585
R342 B.n1236 B.n139 585
R343 B.n1230 B.n1229 585
R344 B.n1229 B.n135 585
R345 B.n1228 B.n134 585
R346 B.n1242 B.n134 585
R347 B.n1227 B.n133 585
R348 B.n1243 B.n133 585
R349 B.n1226 B.n132 585
R350 B.n1244 B.n132 585
R351 B.n1225 B.n1224 585
R352 B.n1224 B.n128 585
R353 B.n1223 B.n127 585
R354 B.n1250 B.n127 585
R355 B.n1222 B.n126 585
R356 B.n1251 B.n126 585
R357 B.n1221 B.n125 585
R358 B.n1252 B.n125 585
R359 B.n1220 B.n1219 585
R360 B.n1219 B.n124 585
R361 B.n1218 B.n120 585
R362 B.n1258 B.n120 585
R363 B.n1217 B.n119 585
R364 B.n1259 B.n119 585
R365 B.n1216 B.n118 585
R366 B.n1260 B.n118 585
R367 B.n1215 B.n1214 585
R368 B.n1214 B.n114 585
R369 B.n1213 B.n113 585
R370 B.n1266 B.n113 585
R371 B.n1212 B.n112 585
R372 B.n1267 B.n112 585
R373 B.n1211 B.n111 585
R374 B.n1268 B.n111 585
R375 B.n1210 B.n1209 585
R376 B.n1209 B.n107 585
R377 B.n1208 B.n106 585
R378 B.n1274 B.n106 585
R379 B.n1207 B.n105 585
R380 B.n1275 B.n105 585
R381 B.n1206 B.n104 585
R382 B.n1276 B.n104 585
R383 B.n1205 B.n1204 585
R384 B.n1204 B.n100 585
R385 B.n1203 B.n99 585
R386 B.n1282 B.n99 585
R387 B.n1202 B.n98 585
R388 B.n1283 B.n98 585
R389 B.n1201 B.n97 585
R390 B.n1284 B.n97 585
R391 B.n1200 B.n1199 585
R392 B.n1199 B.n93 585
R393 B.n1198 B.n92 585
R394 B.n1290 B.n92 585
R395 B.n1197 B.n91 585
R396 B.n1291 B.n91 585
R397 B.n1196 B.n90 585
R398 B.n1292 B.n90 585
R399 B.n1195 B.n1194 585
R400 B.n1194 B.n86 585
R401 B.n1193 B.n85 585
R402 B.n1298 B.n85 585
R403 B.n1192 B.n84 585
R404 B.n1299 B.n84 585
R405 B.n1191 B.n83 585
R406 B.n1300 B.n83 585
R407 B.n1190 B.n1189 585
R408 B.n1189 B.n79 585
R409 B.n1188 B.n78 585
R410 B.n1306 B.n78 585
R411 B.n1187 B.n77 585
R412 B.n1307 B.n77 585
R413 B.n1186 B.n76 585
R414 B.n1308 B.n76 585
R415 B.n1185 B.n1184 585
R416 B.n1184 B.n72 585
R417 B.n1183 B.n71 585
R418 B.n1314 B.n71 585
R419 B.n1182 B.n70 585
R420 B.n1315 B.n70 585
R421 B.n1181 B.n69 585
R422 B.n1316 B.n69 585
R423 B.n1180 B.n1179 585
R424 B.n1179 B.n65 585
R425 B.n1178 B.n64 585
R426 B.n1322 B.n64 585
R427 B.n1177 B.n63 585
R428 B.n1323 B.n63 585
R429 B.n1176 B.n62 585
R430 B.n1324 B.n62 585
R431 B.n1175 B.n1174 585
R432 B.n1174 B.n58 585
R433 B.n1173 B.n57 585
R434 B.n1330 B.n57 585
R435 B.n1172 B.n56 585
R436 B.n1331 B.n56 585
R437 B.n1171 B.n55 585
R438 B.n1332 B.n55 585
R439 B.n1170 B.n1169 585
R440 B.n1169 B.n51 585
R441 B.n1168 B.n50 585
R442 B.n1338 B.n50 585
R443 B.n1167 B.n49 585
R444 B.n1339 B.n49 585
R445 B.n1166 B.n48 585
R446 B.n1340 B.n48 585
R447 B.n1165 B.n1164 585
R448 B.n1164 B.n44 585
R449 B.n1163 B.n43 585
R450 B.n1346 B.n43 585
R451 B.n1162 B.n42 585
R452 B.n1347 B.n42 585
R453 B.n1161 B.n41 585
R454 B.n1348 B.n41 585
R455 B.n1160 B.n1159 585
R456 B.n1159 B.n40 585
R457 B.n1158 B.n36 585
R458 B.n1354 B.n36 585
R459 B.n1157 B.n35 585
R460 B.n1355 B.n35 585
R461 B.n1156 B.n34 585
R462 B.n1356 B.n34 585
R463 B.n1155 B.n1154 585
R464 B.n1154 B.n30 585
R465 B.n1153 B.n29 585
R466 B.n1362 B.n29 585
R467 B.n1152 B.n28 585
R468 B.n1363 B.n28 585
R469 B.n1151 B.n27 585
R470 B.n1364 B.n27 585
R471 B.n1150 B.n1149 585
R472 B.n1149 B.n23 585
R473 B.n1148 B.n22 585
R474 B.n1370 B.n22 585
R475 B.n1147 B.n21 585
R476 B.n1371 B.n21 585
R477 B.n1146 B.n20 585
R478 B.n1372 B.n20 585
R479 B.n1145 B.n1144 585
R480 B.n1144 B.n19 585
R481 B.n1143 B.n15 585
R482 B.n1378 B.n15 585
R483 B.n1142 B.n14 585
R484 B.n1379 B.n14 585
R485 B.n1141 B.n13 585
R486 B.n1380 B.n13 585
R487 B.n1140 B.n1139 585
R488 B.n1139 B.n12 585
R489 B.n1138 B.n1137 585
R490 B.n1138 B.n8 585
R491 B.n1136 B.n7 585
R492 B.n1387 B.n7 585
R493 B.n1135 B.n6 585
R494 B.n1388 B.n6 585
R495 B.n1134 B.n5 585
R496 B.n1389 B.n5 585
R497 B.n1133 B.n1132 585
R498 B.n1132 B.n4 585
R499 B.n1131 B.n446 585
R500 B.n1131 B.n1130 585
R501 B.n1121 B.n447 585
R502 B.n448 B.n447 585
R503 B.n1123 B.n1122 585
R504 B.n1124 B.n1123 585
R505 B.n1120 B.n453 585
R506 B.n453 B.n452 585
R507 B.n1119 B.n1118 585
R508 B.n1118 B.n1117 585
R509 B.n455 B.n454 585
R510 B.n1110 B.n455 585
R511 B.n1109 B.n1108 585
R512 B.n1111 B.n1109 585
R513 B.n1107 B.n460 585
R514 B.n460 B.n459 585
R515 B.n1106 B.n1105 585
R516 B.n1105 B.n1104 585
R517 B.n462 B.n461 585
R518 B.n463 B.n462 585
R519 B.n1097 B.n1096 585
R520 B.n1098 B.n1097 585
R521 B.n1095 B.n468 585
R522 B.n468 B.n467 585
R523 B.n1094 B.n1093 585
R524 B.n1093 B.n1092 585
R525 B.n470 B.n469 585
R526 B.n471 B.n470 585
R527 B.n1085 B.n1084 585
R528 B.n1086 B.n1085 585
R529 B.n1083 B.n476 585
R530 B.n476 B.n475 585
R531 B.n1082 B.n1081 585
R532 B.n1081 B.n1080 585
R533 B.n478 B.n477 585
R534 B.n1073 B.n478 585
R535 B.n1072 B.n1071 585
R536 B.n1074 B.n1072 585
R537 B.n1070 B.n483 585
R538 B.n483 B.n482 585
R539 B.n1069 B.n1068 585
R540 B.n1068 B.n1067 585
R541 B.n485 B.n484 585
R542 B.n486 B.n485 585
R543 B.n1060 B.n1059 585
R544 B.n1061 B.n1060 585
R545 B.n1058 B.n491 585
R546 B.n491 B.n490 585
R547 B.n1057 B.n1056 585
R548 B.n1056 B.n1055 585
R549 B.n493 B.n492 585
R550 B.n494 B.n493 585
R551 B.n1048 B.n1047 585
R552 B.n1049 B.n1048 585
R553 B.n1046 B.n499 585
R554 B.n499 B.n498 585
R555 B.n1045 B.n1044 585
R556 B.n1044 B.n1043 585
R557 B.n501 B.n500 585
R558 B.n502 B.n501 585
R559 B.n1036 B.n1035 585
R560 B.n1037 B.n1036 585
R561 B.n1034 B.n507 585
R562 B.n507 B.n506 585
R563 B.n1033 B.n1032 585
R564 B.n1032 B.n1031 585
R565 B.n509 B.n508 585
R566 B.n510 B.n509 585
R567 B.n1024 B.n1023 585
R568 B.n1025 B.n1024 585
R569 B.n1022 B.n515 585
R570 B.n515 B.n514 585
R571 B.n1021 B.n1020 585
R572 B.n1020 B.n1019 585
R573 B.n517 B.n516 585
R574 B.n518 B.n517 585
R575 B.n1012 B.n1011 585
R576 B.n1013 B.n1012 585
R577 B.n1010 B.n522 585
R578 B.n526 B.n522 585
R579 B.n1009 B.n1008 585
R580 B.n1008 B.n1007 585
R581 B.n524 B.n523 585
R582 B.n525 B.n524 585
R583 B.n1000 B.n999 585
R584 B.n1001 B.n1000 585
R585 B.n998 B.n531 585
R586 B.n531 B.n530 585
R587 B.n997 B.n996 585
R588 B.n996 B.n995 585
R589 B.n533 B.n532 585
R590 B.n534 B.n533 585
R591 B.n988 B.n987 585
R592 B.n989 B.n988 585
R593 B.n986 B.n539 585
R594 B.n539 B.n538 585
R595 B.n985 B.n984 585
R596 B.n984 B.n983 585
R597 B.n541 B.n540 585
R598 B.n542 B.n541 585
R599 B.n976 B.n975 585
R600 B.n977 B.n976 585
R601 B.n974 B.n546 585
R602 B.n550 B.n546 585
R603 B.n973 B.n972 585
R604 B.n972 B.n971 585
R605 B.n548 B.n547 585
R606 B.n549 B.n548 585
R607 B.n964 B.n963 585
R608 B.n965 B.n964 585
R609 B.n962 B.n555 585
R610 B.n555 B.n554 585
R611 B.n961 B.n960 585
R612 B.n960 B.n959 585
R613 B.n557 B.n556 585
R614 B.n558 B.n557 585
R615 B.n952 B.n951 585
R616 B.n953 B.n952 585
R617 B.n950 B.n563 585
R618 B.n563 B.n562 585
R619 B.n949 B.n948 585
R620 B.n948 B.n947 585
R621 B.n565 B.n564 585
R622 B.n566 B.n565 585
R623 B.n940 B.n939 585
R624 B.n941 B.n940 585
R625 B.n938 B.n571 585
R626 B.n571 B.n570 585
R627 B.n937 B.n936 585
R628 B.n936 B.n935 585
R629 B.n573 B.n572 585
R630 B.n928 B.n573 585
R631 B.n927 B.n926 585
R632 B.n929 B.n927 585
R633 B.n925 B.n578 585
R634 B.n578 B.n577 585
R635 B.n924 B.n923 585
R636 B.n923 B.n922 585
R637 B.n580 B.n579 585
R638 B.n581 B.n580 585
R639 B.n915 B.n914 585
R640 B.n916 B.n915 585
R641 B.n913 B.n586 585
R642 B.n586 B.n585 585
R643 B.n912 B.n911 585
R644 B.n911 B.n910 585
R645 B.n588 B.n587 585
R646 B.n589 B.n588 585
R647 B.n903 B.n902 585
R648 B.n904 B.n903 585
R649 B.n592 B.n591 585
R650 B.n659 B.n657 585
R651 B.n660 B.n656 585
R652 B.n660 B.n593 585
R653 B.n663 B.n662 585
R654 B.n664 B.n655 585
R655 B.n666 B.n665 585
R656 B.n668 B.n654 585
R657 B.n671 B.n670 585
R658 B.n672 B.n653 585
R659 B.n674 B.n673 585
R660 B.n676 B.n652 585
R661 B.n679 B.n678 585
R662 B.n680 B.n651 585
R663 B.n682 B.n681 585
R664 B.n684 B.n650 585
R665 B.n687 B.n686 585
R666 B.n688 B.n649 585
R667 B.n690 B.n689 585
R668 B.n692 B.n648 585
R669 B.n695 B.n694 585
R670 B.n696 B.n647 585
R671 B.n698 B.n697 585
R672 B.n700 B.n646 585
R673 B.n703 B.n702 585
R674 B.n704 B.n645 585
R675 B.n706 B.n705 585
R676 B.n708 B.n644 585
R677 B.n711 B.n710 585
R678 B.n712 B.n643 585
R679 B.n714 B.n713 585
R680 B.n716 B.n642 585
R681 B.n719 B.n718 585
R682 B.n720 B.n641 585
R683 B.n722 B.n721 585
R684 B.n724 B.n640 585
R685 B.n727 B.n726 585
R686 B.n728 B.n639 585
R687 B.n730 B.n729 585
R688 B.n732 B.n638 585
R689 B.n735 B.n734 585
R690 B.n736 B.n637 585
R691 B.n738 B.n737 585
R692 B.n740 B.n636 585
R693 B.n743 B.n742 585
R694 B.n744 B.n635 585
R695 B.n746 B.n745 585
R696 B.n748 B.n634 585
R697 B.n751 B.n750 585
R698 B.n752 B.n633 585
R699 B.n754 B.n753 585
R700 B.n756 B.n632 585
R701 B.n759 B.n758 585
R702 B.n760 B.n631 585
R703 B.n762 B.n761 585
R704 B.n764 B.n630 585
R705 B.n767 B.n766 585
R706 B.n769 B.n627 585
R707 B.n771 B.n770 585
R708 B.n773 B.n626 585
R709 B.n776 B.n775 585
R710 B.n777 B.n625 585
R711 B.n779 B.n778 585
R712 B.n781 B.n624 585
R713 B.n784 B.n783 585
R714 B.n785 B.n623 585
R715 B.n790 B.n789 585
R716 B.n792 B.n622 585
R717 B.n795 B.n794 585
R718 B.n796 B.n621 585
R719 B.n798 B.n797 585
R720 B.n800 B.n620 585
R721 B.n803 B.n802 585
R722 B.n804 B.n619 585
R723 B.n806 B.n805 585
R724 B.n808 B.n618 585
R725 B.n811 B.n810 585
R726 B.n812 B.n617 585
R727 B.n814 B.n813 585
R728 B.n816 B.n616 585
R729 B.n819 B.n818 585
R730 B.n820 B.n615 585
R731 B.n822 B.n821 585
R732 B.n824 B.n614 585
R733 B.n827 B.n826 585
R734 B.n828 B.n613 585
R735 B.n830 B.n829 585
R736 B.n832 B.n612 585
R737 B.n835 B.n834 585
R738 B.n836 B.n611 585
R739 B.n838 B.n837 585
R740 B.n840 B.n610 585
R741 B.n843 B.n842 585
R742 B.n844 B.n609 585
R743 B.n846 B.n845 585
R744 B.n848 B.n608 585
R745 B.n851 B.n850 585
R746 B.n852 B.n607 585
R747 B.n854 B.n853 585
R748 B.n856 B.n606 585
R749 B.n859 B.n858 585
R750 B.n860 B.n605 585
R751 B.n862 B.n861 585
R752 B.n864 B.n604 585
R753 B.n867 B.n866 585
R754 B.n868 B.n603 585
R755 B.n870 B.n869 585
R756 B.n872 B.n602 585
R757 B.n875 B.n874 585
R758 B.n876 B.n601 585
R759 B.n878 B.n877 585
R760 B.n880 B.n600 585
R761 B.n883 B.n882 585
R762 B.n884 B.n599 585
R763 B.n886 B.n885 585
R764 B.n888 B.n598 585
R765 B.n891 B.n890 585
R766 B.n892 B.n597 585
R767 B.n894 B.n893 585
R768 B.n896 B.n596 585
R769 B.n897 B.n595 585
R770 B.n900 B.n899 585
R771 B.n901 B.n594 585
R772 B.n594 B.n593 585
R773 B.n906 B.n905 585
R774 B.n905 B.n904 585
R775 B.n907 B.n590 585
R776 B.n590 B.n589 585
R777 B.n909 B.n908 585
R778 B.n910 B.n909 585
R779 B.n584 B.n583 585
R780 B.n585 B.n584 585
R781 B.n918 B.n917 585
R782 B.n917 B.n916 585
R783 B.n919 B.n582 585
R784 B.n582 B.n581 585
R785 B.n921 B.n920 585
R786 B.n922 B.n921 585
R787 B.n576 B.n575 585
R788 B.n577 B.n576 585
R789 B.n931 B.n930 585
R790 B.n930 B.n929 585
R791 B.n932 B.n574 585
R792 B.n928 B.n574 585
R793 B.n934 B.n933 585
R794 B.n935 B.n934 585
R795 B.n569 B.n568 585
R796 B.n570 B.n569 585
R797 B.n943 B.n942 585
R798 B.n942 B.n941 585
R799 B.n944 B.n567 585
R800 B.n567 B.n566 585
R801 B.n946 B.n945 585
R802 B.n947 B.n946 585
R803 B.n561 B.n560 585
R804 B.n562 B.n561 585
R805 B.n955 B.n954 585
R806 B.n954 B.n953 585
R807 B.n956 B.n559 585
R808 B.n559 B.n558 585
R809 B.n958 B.n957 585
R810 B.n959 B.n958 585
R811 B.n553 B.n552 585
R812 B.n554 B.n553 585
R813 B.n967 B.n966 585
R814 B.n966 B.n965 585
R815 B.n968 B.n551 585
R816 B.n551 B.n549 585
R817 B.n970 B.n969 585
R818 B.n971 B.n970 585
R819 B.n545 B.n544 585
R820 B.n550 B.n545 585
R821 B.n979 B.n978 585
R822 B.n978 B.n977 585
R823 B.n980 B.n543 585
R824 B.n543 B.n542 585
R825 B.n982 B.n981 585
R826 B.n983 B.n982 585
R827 B.n537 B.n536 585
R828 B.n538 B.n537 585
R829 B.n991 B.n990 585
R830 B.n990 B.n989 585
R831 B.n992 B.n535 585
R832 B.n535 B.n534 585
R833 B.n994 B.n993 585
R834 B.n995 B.n994 585
R835 B.n529 B.n528 585
R836 B.n530 B.n529 585
R837 B.n1003 B.n1002 585
R838 B.n1002 B.n1001 585
R839 B.n1004 B.n527 585
R840 B.n527 B.n525 585
R841 B.n1006 B.n1005 585
R842 B.n1007 B.n1006 585
R843 B.n521 B.n520 585
R844 B.n526 B.n521 585
R845 B.n1015 B.n1014 585
R846 B.n1014 B.n1013 585
R847 B.n1016 B.n519 585
R848 B.n519 B.n518 585
R849 B.n1018 B.n1017 585
R850 B.n1019 B.n1018 585
R851 B.n513 B.n512 585
R852 B.n514 B.n513 585
R853 B.n1027 B.n1026 585
R854 B.n1026 B.n1025 585
R855 B.n1028 B.n511 585
R856 B.n511 B.n510 585
R857 B.n1030 B.n1029 585
R858 B.n1031 B.n1030 585
R859 B.n505 B.n504 585
R860 B.n506 B.n505 585
R861 B.n1039 B.n1038 585
R862 B.n1038 B.n1037 585
R863 B.n1040 B.n503 585
R864 B.n503 B.n502 585
R865 B.n1042 B.n1041 585
R866 B.n1043 B.n1042 585
R867 B.n497 B.n496 585
R868 B.n498 B.n497 585
R869 B.n1051 B.n1050 585
R870 B.n1050 B.n1049 585
R871 B.n1052 B.n495 585
R872 B.n495 B.n494 585
R873 B.n1054 B.n1053 585
R874 B.n1055 B.n1054 585
R875 B.n489 B.n488 585
R876 B.n490 B.n489 585
R877 B.n1063 B.n1062 585
R878 B.n1062 B.n1061 585
R879 B.n1064 B.n487 585
R880 B.n487 B.n486 585
R881 B.n1066 B.n1065 585
R882 B.n1067 B.n1066 585
R883 B.n481 B.n480 585
R884 B.n482 B.n481 585
R885 B.n1076 B.n1075 585
R886 B.n1075 B.n1074 585
R887 B.n1077 B.n479 585
R888 B.n1073 B.n479 585
R889 B.n1079 B.n1078 585
R890 B.n1080 B.n1079 585
R891 B.n474 B.n473 585
R892 B.n475 B.n474 585
R893 B.n1088 B.n1087 585
R894 B.n1087 B.n1086 585
R895 B.n1089 B.n472 585
R896 B.n472 B.n471 585
R897 B.n1091 B.n1090 585
R898 B.n1092 B.n1091 585
R899 B.n466 B.n465 585
R900 B.n467 B.n466 585
R901 B.n1100 B.n1099 585
R902 B.n1099 B.n1098 585
R903 B.n1101 B.n464 585
R904 B.n464 B.n463 585
R905 B.n1103 B.n1102 585
R906 B.n1104 B.n1103 585
R907 B.n458 B.n457 585
R908 B.n459 B.n458 585
R909 B.n1113 B.n1112 585
R910 B.n1112 B.n1111 585
R911 B.n1114 B.n456 585
R912 B.n1110 B.n456 585
R913 B.n1116 B.n1115 585
R914 B.n1117 B.n1116 585
R915 B.n451 B.n450 585
R916 B.n452 B.n451 585
R917 B.n1126 B.n1125 585
R918 B.n1125 B.n1124 585
R919 B.n1127 B.n449 585
R920 B.n449 B.n448 585
R921 B.n1129 B.n1128 585
R922 B.n1130 B.n1129 585
R923 B.n3 B.n0 585
R924 B.n4 B.n3 585
R925 B.n1386 B.n1 585
R926 B.n1387 B.n1386 585
R927 B.n1385 B.n1384 585
R928 B.n1385 B.n8 585
R929 B.n1383 B.n9 585
R930 B.n12 B.n9 585
R931 B.n1382 B.n1381 585
R932 B.n1381 B.n1380 585
R933 B.n11 B.n10 585
R934 B.n1379 B.n11 585
R935 B.n1377 B.n1376 585
R936 B.n1378 B.n1377 585
R937 B.n1375 B.n16 585
R938 B.n19 B.n16 585
R939 B.n1374 B.n1373 585
R940 B.n1373 B.n1372 585
R941 B.n18 B.n17 585
R942 B.n1371 B.n18 585
R943 B.n1369 B.n1368 585
R944 B.n1370 B.n1369 585
R945 B.n1367 B.n24 585
R946 B.n24 B.n23 585
R947 B.n1366 B.n1365 585
R948 B.n1365 B.n1364 585
R949 B.n26 B.n25 585
R950 B.n1363 B.n26 585
R951 B.n1361 B.n1360 585
R952 B.n1362 B.n1361 585
R953 B.n1359 B.n31 585
R954 B.n31 B.n30 585
R955 B.n1358 B.n1357 585
R956 B.n1357 B.n1356 585
R957 B.n33 B.n32 585
R958 B.n1355 B.n33 585
R959 B.n1353 B.n1352 585
R960 B.n1354 B.n1353 585
R961 B.n1351 B.n37 585
R962 B.n40 B.n37 585
R963 B.n1350 B.n1349 585
R964 B.n1349 B.n1348 585
R965 B.n39 B.n38 585
R966 B.n1347 B.n39 585
R967 B.n1345 B.n1344 585
R968 B.n1346 B.n1345 585
R969 B.n1343 B.n45 585
R970 B.n45 B.n44 585
R971 B.n1342 B.n1341 585
R972 B.n1341 B.n1340 585
R973 B.n47 B.n46 585
R974 B.n1339 B.n47 585
R975 B.n1337 B.n1336 585
R976 B.n1338 B.n1337 585
R977 B.n1335 B.n52 585
R978 B.n52 B.n51 585
R979 B.n1334 B.n1333 585
R980 B.n1333 B.n1332 585
R981 B.n54 B.n53 585
R982 B.n1331 B.n54 585
R983 B.n1329 B.n1328 585
R984 B.n1330 B.n1329 585
R985 B.n1327 B.n59 585
R986 B.n59 B.n58 585
R987 B.n1326 B.n1325 585
R988 B.n1325 B.n1324 585
R989 B.n61 B.n60 585
R990 B.n1323 B.n61 585
R991 B.n1321 B.n1320 585
R992 B.n1322 B.n1321 585
R993 B.n1319 B.n66 585
R994 B.n66 B.n65 585
R995 B.n1318 B.n1317 585
R996 B.n1317 B.n1316 585
R997 B.n68 B.n67 585
R998 B.n1315 B.n68 585
R999 B.n1313 B.n1312 585
R1000 B.n1314 B.n1313 585
R1001 B.n1311 B.n73 585
R1002 B.n73 B.n72 585
R1003 B.n1310 B.n1309 585
R1004 B.n1309 B.n1308 585
R1005 B.n75 B.n74 585
R1006 B.n1307 B.n75 585
R1007 B.n1305 B.n1304 585
R1008 B.n1306 B.n1305 585
R1009 B.n1303 B.n80 585
R1010 B.n80 B.n79 585
R1011 B.n1302 B.n1301 585
R1012 B.n1301 B.n1300 585
R1013 B.n82 B.n81 585
R1014 B.n1299 B.n82 585
R1015 B.n1297 B.n1296 585
R1016 B.n1298 B.n1297 585
R1017 B.n1295 B.n87 585
R1018 B.n87 B.n86 585
R1019 B.n1294 B.n1293 585
R1020 B.n1293 B.n1292 585
R1021 B.n89 B.n88 585
R1022 B.n1291 B.n89 585
R1023 B.n1289 B.n1288 585
R1024 B.n1290 B.n1289 585
R1025 B.n1287 B.n94 585
R1026 B.n94 B.n93 585
R1027 B.n1286 B.n1285 585
R1028 B.n1285 B.n1284 585
R1029 B.n96 B.n95 585
R1030 B.n1283 B.n96 585
R1031 B.n1281 B.n1280 585
R1032 B.n1282 B.n1281 585
R1033 B.n1279 B.n101 585
R1034 B.n101 B.n100 585
R1035 B.n1278 B.n1277 585
R1036 B.n1277 B.n1276 585
R1037 B.n103 B.n102 585
R1038 B.n1275 B.n103 585
R1039 B.n1273 B.n1272 585
R1040 B.n1274 B.n1273 585
R1041 B.n1271 B.n108 585
R1042 B.n108 B.n107 585
R1043 B.n1270 B.n1269 585
R1044 B.n1269 B.n1268 585
R1045 B.n110 B.n109 585
R1046 B.n1267 B.n110 585
R1047 B.n1265 B.n1264 585
R1048 B.n1266 B.n1265 585
R1049 B.n1263 B.n115 585
R1050 B.n115 B.n114 585
R1051 B.n1262 B.n1261 585
R1052 B.n1261 B.n1260 585
R1053 B.n117 B.n116 585
R1054 B.n1259 B.n117 585
R1055 B.n1257 B.n1256 585
R1056 B.n1258 B.n1257 585
R1057 B.n1255 B.n121 585
R1058 B.n124 B.n121 585
R1059 B.n1254 B.n1253 585
R1060 B.n1253 B.n1252 585
R1061 B.n123 B.n122 585
R1062 B.n1251 B.n123 585
R1063 B.n1249 B.n1248 585
R1064 B.n1250 B.n1249 585
R1065 B.n1247 B.n129 585
R1066 B.n129 B.n128 585
R1067 B.n1246 B.n1245 585
R1068 B.n1245 B.n1244 585
R1069 B.n131 B.n130 585
R1070 B.n1243 B.n131 585
R1071 B.n1241 B.n1240 585
R1072 B.n1242 B.n1241 585
R1073 B.n1239 B.n136 585
R1074 B.n136 B.n135 585
R1075 B.n1238 B.n1237 585
R1076 B.n1237 B.n1236 585
R1077 B.n1390 B.n1389 585
R1078 B.n1388 B.n2 585
R1079 B.n1237 B.n138 511.721
R1080 B.n1233 B.n139 511.721
R1081 B.n903 B.n594 511.721
R1082 B.n905 B.n592 511.721
R1083 B.n204 B.t14 325
R1084 B.n201 B.t21 325
R1085 B.n786 B.t10 325
R1086 B.n628 B.t18 325
R1087 B.n1235 B.n1234 256.663
R1088 B.n1235 B.n199 256.663
R1089 B.n1235 B.n198 256.663
R1090 B.n1235 B.n197 256.663
R1091 B.n1235 B.n196 256.663
R1092 B.n1235 B.n195 256.663
R1093 B.n1235 B.n194 256.663
R1094 B.n1235 B.n193 256.663
R1095 B.n1235 B.n192 256.663
R1096 B.n1235 B.n191 256.663
R1097 B.n1235 B.n190 256.663
R1098 B.n1235 B.n189 256.663
R1099 B.n1235 B.n188 256.663
R1100 B.n1235 B.n187 256.663
R1101 B.n1235 B.n186 256.663
R1102 B.n1235 B.n185 256.663
R1103 B.n1235 B.n184 256.663
R1104 B.n1235 B.n183 256.663
R1105 B.n1235 B.n182 256.663
R1106 B.n1235 B.n181 256.663
R1107 B.n1235 B.n180 256.663
R1108 B.n1235 B.n179 256.663
R1109 B.n1235 B.n178 256.663
R1110 B.n1235 B.n177 256.663
R1111 B.n1235 B.n176 256.663
R1112 B.n1235 B.n175 256.663
R1113 B.n1235 B.n174 256.663
R1114 B.n1235 B.n173 256.663
R1115 B.n1235 B.n172 256.663
R1116 B.n1235 B.n171 256.663
R1117 B.n1235 B.n170 256.663
R1118 B.n1235 B.n169 256.663
R1119 B.n1235 B.n168 256.663
R1120 B.n1235 B.n167 256.663
R1121 B.n1235 B.n166 256.663
R1122 B.n1235 B.n165 256.663
R1123 B.n1235 B.n164 256.663
R1124 B.n1235 B.n163 256.663
R1125 B.n1235 B.n162 256.663
R1126 B.n1235 B.n161 256.663
R1127 B.n1235 B.n160 256.663
R1128 B.n1235 B.n159 256.663
R1129 B.n1235 B.n158 256.663
R1130 B.n1235 B.n157 256.663
R1131 B.n1235 B.n156 256.663
R1132 B.n1235 B.n155 256.663
R1133 B.n1235 B.n154 256.663
R1134 B.n1235 B.n153 256.663
R1135 B.n1235 B.n152 256.663
R1136 B.n1235 B.n151 256.663
R1137 B.n1235 B.n150 256.663
R1138 B.n1235 B.n149 256.663
R1139 B.n1235 B.n148 256.663
R1140 B.n1235 B.n147 256.663
R1141 B.n1235 B.n146 256.663
R1142 B.n1235 B.n145 256.663
R1143 B.n1235 B.n144 256.663
R1144 B.n1235 B.n143 256.663
R1145 B.n1235 B.n142 256.663
R1146 B.n1235 B.n141 256.663
R1147 B.n1235 B.n140 256.663
R1148 B.n658 B.n593 256.663
R1149 B.n661 B.n593 256.663
R1150 B.n667 B.n593 256.663
R1151 B.n669 B.n593 256.663
R1152 B.n675 B.n593 256.663
R1153 B.n677 B.n593 256.663
R1154 B.n683 B.n593 256.663
R1155 B.n685 B.n593 256.663
R1156 B.n691 B.n593 256.663
R1157 B.n693 B.n593 256.663
R1158 B.n699 B.n593 256.663
R1159 B.n701 B.n593 256.663
R1160 B.n707 B.n593 256.663
R1161 B.n709 B.n593 256.663
R1162 B.n715 B.n593 256.663
R1163 B.n717 B.n593 256.663
R1164 B.n723 B.n593 256.663
R1165 B.n725 B.n593 256.663
R1166 B.n731 B.n593 256.663
R1167 B.n733 B.n593 256.663
R1168 B.n739 B.n593 256.663
R1169 B.n741 B.n593 256.663
R1170 B.n747 B.n593 256.663
R1171 B.n749 B.n593 256.663
R1172 B.n755 B.n593 256.663
R1173 B.n757 B.n593 256.663
R1174 B.n763 B.n593 256.663
R1175 B.n765 B.n593 256.663
R1176 B.n772 B.n593 256.663
R1177 B.n774 B.n593 256.663
R1178 B.n780 B.n593 256.663
R1179 B.n782 B.n593 256.663
R1180 B.n791 B.n593 256.663
R1181 B.n793 B.n593 256.663
R1182 B.n799 B.n593 256.663
R1183 B.n801 B.n593 256.663
R1184 B.n807 B.n593 256.663
R1185 B.n809 B.n593 256.663
R1186 B.n815 B.n593 256.663
R1187 B.n817 B.n593 256.663
R1188 B.n823 B.n593 256.663
R1189 B.n825 B.n593 256.663
R1190 B.n831 B.n593 256.663
R1191 B.n833 B.n593 256.663
R1192 B.n839 B.n593 256.663
R1193 B.n841 B.n593 256.663
R1194 B.n847 B.n593 256.663
R1195 B.n849 B.n593 256.663
R1196 B.n855 B.n593 256.663
R1197 B.n857 B.n593 256.663
R1198 B.n863 B.n593 256.663
R1199 B.n865 B.n593 256.663
R1200 B.n871 B.n593 256.663
R1201 B.n873 B.n593 256.663
R1202 B.n879 B.n593 256.663
R1203 B.n881 B.n593 256.663
R1204 B.n887 B.n593 256.663
R1205 B.n889 B.n593 256.663
R1206 B.n895 B.n593 256.663
R1207 B.n898 B.n593 256.663
R1208 B.n1392 B.n1391 256.663
R1209 B.n209 B.n208 163.367
R1210 B.n213 B.n212 163.367
R1211 B.n217 B.n216 163.367
R1212 B.n221 B.n220 163.367
R1213 B.n225 B.n224 163.367
R1214 B.n229 B.n228 163.367
R1215 B.n233 B.n232 163.367
R1216 B.n237 B.n236 163.367
R1217 B.n241 B.n240 163.367
R1218 B.n245 B.n244 163.367
R1219 B.n249 B.n248 163.367
R1220 B.n253 B.n252 163.367
R1221 B.n257 B.n256 163.367
R1222 B.n261 B.n260 163.367
R1223 B.n265 B.n264 163.367
R1224 B.n269 B.n268 163.367
R1225 B.n273 B.n272 163.367
R1226 B.n277 B.n276 163.367
R1227 B.n281 B.n280 163.367
R1228 B.n285 B.n284 163.367
R1229 B.n289 B.n288 163.367
R1230 B.n293 B.n292 163.367
R1231 B.n297 B.n296 163.367
R1232 B.n301 B.n300 163.367
R1233 B.n305 B.n304 163.367
R1234 B.n309 B.n308 163.367
R1235 B.n313 B.n312 163.367
R1236 B.n317 B.n316 163.367
R1237 B.n321 B.n320 163.367
R1238 B.n325 B.n324 163.367
R1239 B.n329 B.n328 163.367
R1240 B.n333 B.n332 163.367
R1241 B.n337 B.n336 163.367
R1242 B.n341 B.n340 163.367
R1243 B.n345 B.n344 163.367
R1244 B.n349 B.n348 163.367
R1245 B.n353 B.n352 163.367
R1246 B.n357 B.n356 163.367
R1247 B.n361 B.n360 163.367
R1248 B.n365 B.n364 163.367
R1249 B.n369 B.n368 163.367
R1250 B.n373 B.n372 163.367
R1251 B.n377 B.n376 163.367
R1252 B.n381 B.n380 163.367
R1253 B.n385 B.n384 163.367
R1254 B.n389 B.n388 163.367
R1255 B.n393 B.n392 163.367
R1256 B.n397 B.n396 163.367
R1257 B.n401 B.n400 163.367
R1258 B.n405 B.n404 163.367
R1259 B.n409 B.n408 163.367
R1260 B.n413 B.n412 163.367
R1261 B.n417 B.n416 163.367
R1262 B.n421 B.n420 163.367
R1263 B.n425 B.n424 163.367
R1264 B.n429 B.n428 163.367
R1265 B.n433 B.n432 163.367
R1266 B.n437 B.n436 163.367
R1267 B.n441 B.n440 163.367
R1268 B.n443 B.n200 163.367
R1269 B.n903 B.n588 163.367
R1270 B.n911 B.n588 163.367
R1271 B.n911 B.n586 163.367
R1272 B.n915 B.n586 163.367
R1273 B.n915 B.n580 163.367
R1274 B.n923 B.n580 163.367
R1275 B.n923 B.n578 163.367
R1276 B.n927 B.n578 163.367
R1277 B.n927 B.n573 163.367
R1278 B.n936 B.n573 163.367
R1279 B.n936 B.n571 163.367
R1280 B.n940 B.n571 163.367
R1281 B.n940 B.n565 163.367
R1282 B.n948 B.n565 163.367
R1283 B.n948 B.n563 163.367
R1284 B.n952 B.n563 163.367
R1285 B.n952 B.n557 163.367
R1286 B.n960 B.n557 163.367
R1287 B.n960 B.n555 163.367
R1288 B.n964 B.n555 163.367
R1289 B.n964 B.n548 163.367
R1290 B.n972 B.n548 163.367
R1291 B.n972 B.n546 163.367
R1292 B.n976 B.n546 163.367
R1293 B.n976 B.n541 163.367
R1294 B.n984 B.n541 163.367
R1295 B.n984 B.n539 163.367
R1296 B.n988 B.n539 163.367
R1297 B.n988 B.n533 163.367
R1298 B.n996 B.n533 163.367
R1299 B.n996 B.n531 163.367
R1300 B.n1000 B.n531 163.367
R1301 B.n1000 B.n524 163.367
R1302 B.n1008 B.n524 163.367
R1303 B.n1008 B.n522 163.367
R1304 B.n1012 B.n522 163.367
R1305 B.n1012 B.n517 163.367
R1306 B.n1020 B.n517 163.367
R1307 B.n1020 B.n515 163.367
R1308 B.n1024 B.n515 163.367
R1309 B.n1024 B.n509 163.367
R1310 B.n1032 B.n509 163.367
R1311 B.n1032 B.n507 163.367
R1312 B.n1036 B.n507 163.367
R1313 B.n1036 B.n501 163.367
R1314 B.n1044 B.n501 163.367
R1315 B.n1044 B.n499 163.367
R1316 B.n1048 B.n499 163.367
R1317 B.n1048 B.n493 163.367
R1318 B.n1056 B.n493 163.367
R1319 B.n1056 B.n491 163.367
R1320 B.n1060 B.n491 163.367
R1321 B.n1060 B.n485 163.367
R1322 B.n1068 B.n485 163.367
R1323 B.n1068 B.n483 163.367
R1324 B.n1072 B.n483 163.367
R1325 B.n1072 B.n478 163.367
R1326 B.n1081 B.n478 163.367
R1327 B.n1081 B.n476 163.367
R1328 B.n1085 B.n476 163.367
R1329 B.n1085 B.n470 163.367
R1330 B.n1093 B.n470 163.367
R1331 B.n1093 B.n468 163.367
R1332 B.n1097 B.n468 163.367
R1333 B.n1097 B.n462 163.367
R1334 B.n1105 B.n462 163.367
R1335 B.n1105 B.n460 163.367
R1336 B.n1109 B.n460 163.367
R1337 B.n1109 B.n455 163.367
R1338 B.n1118 B.n455 163.367
R1339 B.n1118 B.n453 163.367
R1340 B.n1123 B.n453 163.367
R1341 B.n1123 B.n447 163.367
R1342 B.n1131 B.n447 163.367
R1343 B.n1132 B.n1131 163.367
R1344 B.n1132 B.n5 163.367
R1345 B.n6 B.n5 163.367
R1346 B.n7 B.n6 163.367
R1347 B.n1138 B.n7 163.367
R1348 B.n1139 B.n1138 163.367
R1349 B.n1139 B.n13 163.367
R1350 B.n14 B.n13 163.367
R1351 B.n15 B.n14 163.367
R1352 B.n1144 B.n15 163.367
R1353 B.n1144 B.n20 163.367
R1354 B.n21 B.n20 163.367
R1355 B.n22 B.n21 163.367
R1356 B.n1149 B.n22 163.367
R1357 B.n1149 B.n27 163.367
R1358 B.n28 B.n27 163.367
R1359 B.n29 B.n28 163.367
R1360 B.n1154 B.n29 163.367
R1361 B.n1154 B.n34 163.367
R1362 B.n35 B.n34 163.367
R1363 B.n36 B.n35 163.367
R1364 B.n1159 B.n36 163.367
R1365 B.n1159 B.n41 163.367
R1366 B.n42 B.n41 163.367
R1367 B.n43 B.n42 163.367
R1368 B.n1164 B.n43 163.367
R1369 B.n1164 B.n48 163.367
R1370 B.n49 B.n48 163.367
R1371 B.n50 B.n49 163.367
R1372 B.n1169 B.n50 163.367
R1373 B.n1169 B.n55 163.367
R1374 B.n56 B.n55 163.367
R1375 B.n57 B.n56 163.367
R1376 B.n1174 B.n57 163.367
R1377 B.n1174 B.n62 163.367
R1378 B.n63 B.n62 163.367
R1379 B.n64 B.n63 163.367
R1380 B.n1179 B.n64 163.367
R1381 B.n1179 B.n69 163.367
R1382 B.n70 B.n69 163.367
R1383 B.n71 B.n70 163.367
R1384 B.n1184 B.n71 163.367
R1385 B.n1184 B.n76 163.367
R1386 B.n77 B.n76 163.367
R1387 B.n78 B.n77 163.367
R1388 B.n1189 B.n78 163.367
R1389 B.n1189 B.n83 163.367
R1390 B.n84 B.n83 163.367
R1391 B.n85 B.n84 163.367
R1392 B.n1194 B.n85 163.367
R1393 B.n1194 B.n90 163.367
R1394 B.n91 B.n90 163.367
R1395 B.n92 B.n91 163.367
R1396 B.n1199 B.n92 163.367
R1397 B.n1199 B.n97 163.367
R1398 B.n98 B.n97 163.367
R1399 B.n99 B.n98 163.367
R1400 B.n1204 B.n99 163.367
R1401 B.n1204 B.n104 163.367
R1402 B.n105 B.n104 163.367
R1403 B.n106 B.n105 163.367
R1404 B.n1209 B.n106 163.367
R1405 B.n1209 B.n111 163.367
R1406 B.n112 B.n111 163.367
R1407 B.n113 B.n112 163.367
R1408 B.n1214 B.n113 163.367
R1409 B.n1214 B.n118 163.367
R1410 B.n119 B.n118 163.367
R1411 B.n120 B.n119 163.367
R1412 B.n1219 B.n120 163.367
R1413 B.n1219 B.n125 163.367
R1414 B.n126 B.n125 163.367
R1415 B.n127 B.n126 163.367
R1416 B.n1224 B.n127 163.367
R1417 B.n1224 B.n132 163.367
R1418 B.n133 B.n132 163.367
R1419 B.n134 B.n133 163.367
R1420 B.n1229 B.n134 163.367
R1421 B.n1229 B.n139 163.367
R1422 B.n660 B.n659 163.367
R1423 B.n662 B.n660 163.367
R1424 B.n666 B.n655 163.367
R1425 B.n670 B.n668 163.367
R1426 B.n674 B.n653 163.367
R1427 B.n678 B.n676 163.367
R1428 B.n682 B.n651 163.367
R1429 B.n686 B.n684 163.367
R1430 B.n690 B.n649 163.367
R1431 B.n694 B.n692 163.367
R1432 B.n698 B.n647 163.367
R1433 B.n702 B.n700 163.367
R1434 B.n706 B.n645 163.367
R1435 B.n710 B.n708 163.367
R1436 B.n714 B.n643 163.367
R1437 B.n718 B.n716 163.367
R1438 B.n722 B.n641 163.367
R1439 B.n726 B.n724 163.367
R1440 B.n730 B.n639 163.367
R1441 B.n734 B.n732 163.367
R1442 B.n738 B.n637 163.367
R1443 B.n742 B.n740 163.367
R1444 B.n746 B.n635 163.367
R1445 B.n750 B.n748 163.367
R1446 B.n754 B.n633 163.367
R1447 B.n758 B.n756 163.367
R1448 B.n762 B.n631 163.367
R1449 B.n766 B.n764 163.367
R1450 B.n771 B.n627 163.367
R1451 B.n775 B.n773 163.367
R1452 B.n779 B.n625 163.367
R1453 B.n783 B.n781 163.367
R1454 B.n790 B.n623 163.367
R1455 B.n794 B.n792 163.367
R1456 B.n798 B.n621 163.367
R1457 B.n802 B.n800 163.367
R1458 B.n806 B.n619 163.367
R1459 B.n810 B.n808 163.367
R1460 B.n814 B.n617 163.367
R1461 B.n818 B.n816 163.367
R1462 B.n822 B.n615 163.367
R1463 B.n826 B.n824 163.367
R1464 B.n830 B.n613 163.367
R1465 B.n834 B.n832 163.367
R1466 B.n838 B.n611 163.367
R1467 B.n842 B.n840 163.367
R1468 B.n846 B.n609 163.367
R1469 B.n850 B.n848 163.367
R1470 B.n854 B.n607 163.367
R1471 B.n858 B.n856 163.367
R1472 B.n862 B.n605 163.367
R1473 B.n866 B.n864 163.367
R1474 B.n870 B.n603 163.367
R1475 B.n874 B.n872 163.367
R1476 B.n878 B.n601 163.367
R1477 B.n882 B.n880 163.367
R1478 B.n886 B.n599 163.367
R1479 B.n890 B.n888 163.367
R1480 B.n894 B.n597 163.367
R1481 B.n897 B.n896 163.367
R1482 B.n899 B.n594 163.367
R1483 B.n905 B.n590 163.367
R1484 B.n909 B.n590 163.367
R1485 B.n909 B.n584 163.367
R1486 B.n917 B.n584 163.367
R1487 B.n917 B.n582 163.367
R1488 B.n921 B.n582 163.367
R1489 B.n921 B.n576 163.367
R1490 B.n930 B.n576 163.367
R1491 B.n930 B.n574 163.367
R1492 B.n934 B.n574 163.367
R1493 B.n934 B.n569 163.367
R1494 B.n942 B.n569 163.367
R1495 B.n942 B.n567 163.367
R1496 B.n946 B.n567 163.367
R1497 B.n946 B.n561 163.367
R1498 B.n954 B.n561 163.367
R1499 B.n954 B.n559 163.367
R1500 B.n958 B.n559 163.367
R1501 B.n958 B.n553 163.367
R1502 B.n966 B.n553 163.367
R1503 B.n966 B.n551 163.367
R1504 B.n970 B.n551 163.367
R1505 B.n970 B.n545 163.367
R1506 B.n978 B.n545 163.367
R1507 B.n978 B.n543 163.367
R1508 B.n982 B.n543 163.367
R1509 B.n982 B.n537 163.367
R1510 B.n990 B.n537 163.367
R1511 B.n990 B.n535 163.367
R1512 B.n994 B.n535 163.367
R1513 B.n994 B.n529 163.367
R1514 B.n1002 B.n529 163.367
R1515 B.n1002 B.n527 163.367
R1516 B.n1006 B.n527 163.367
R1517 B.n1006 B.n521 163.367
R1518 B.n1014 B.n521 163.367
R1519 B.n1014 B.n519 163.367
R1520 B.n1018 B.n519 163.367
R1521 B.n1018 B.n513 163.367
R1522 B.n1026 B.n513 163.367
R1523 B.n1026 B.n511 163.367
R1524 B.n1030 B.n511 163.367
R1525 B.n1030 B.n505 163.367
R1526 B.n1038 B.n505 163.367
R1527 B.n1038 B.n503 163.367
R1528 B.n1042 B.n503 163.367
R1529 B.n1042 B.n497 163.367
R1530 B.n1050 B.n497 163.367
R1531 B.n1050 B.n495 163.367
R1532 B.n1054 B.n495 163.367
R1533 B.n1054 B.n489 163.367
R1534 B.n1062 B.n489 163.367
R1535 B.n1062 B.n487 163.367
R1536 B.n1066 B.n487 163.367
R1537 B.n1066 B.n481 163.367
R1538 B.n1075 B.n481 163.367
R1539 B.n1075 B.n479 163.367
R1540 B.n1079 B.n479 163.367
R1541 B.n1079 B.n474 163.367
R1542 B.n1087 B.n474 163.367
R1543 B.n1087 B.n472 163.367
R1544 B.n1091 B.n472 163.367
R1545 B.n1091 B.n466 163.367
R1546 B.n1099 B.n466 163.367
R1547 B.n1099 B.n464 163.367
R1548 B.n1103 B.n464 163.367
R1549 B.n1103 B.n458 163.367
R1550 B.n1112 B.n458 163.367
R1551 B.n1112 B.n456 163.367
R1552 B.n1116 B.n456 163.367
R1553 B.n1116 B.n451 163.367
R1554 B.n1125 B.n451 163.367
R1555 B.n1125 B.n449 163.367
R1556 B.n1129 B.n449 163.367
R1557 B.n1129 B.n3 163.367
R1558 B.n1390 B.n3 163.367
R1559 B.n1386 B.n2 163.367
R1560 B.n1386 B.n1385 163.367
R1561 B.n1385 B.n9 163.367
R1562 B.n1381 B.n9 163.367
R1563 B.n1381 B.n11 163.367
R1564 B.n1377 B.n11 163.367
R1565 B.n1377 B.n16 163.367
R1566 B.n1373 B.n16 163.367
R1567 B.n1373 B.n18 163.367
R1568 B.n1369 B.n18 163.367
R1569 B.n1369 B.n24 163.367
R1570 B.n1365 B.n24 163.367
R1571 B.n1365 B.n26 163.367
R1572 B.n1361 B.n26 163.367
R1573 B.n1361 B.n31 163.367
R1574 B.n1357 B.n31 163.367
R1575 B.n1357 B.n33 163.367
R1576 B.n1353 B.n33 163.367
R1577 B.n1353 B.n37 163.367
R1578 B.n1349 B.n37 163.367
R1579 B.n1349 B.n39 163.367
R1580 B.n1345 B.n39 163.367
R1581 B.n1345 B.n45 163.367
R1582 B.n1341 B.n45 163.367
R1583 B.n1341 B.n47 163.367
R1584 B.n1337 B.n47 163.367
R1585 B.n1337 B.n52 163.367
R1586 B.n1333 B.n52 163.367
R1587 B.n1333 B.n54 163.367
R1588 B.n1329 B.n54 163.367
R1589 B.n1329 B.n59 163.367
R1590 B.n1325 B.n59 163.367
R1591 B.n1325 B.n61 163.367
R1592 B.n1321 B.n61 163.367
R1593 B.n1321 B.n66 163.367
R1594 B.n1317 B.n66 163.367
R1595 B.n1317 B.n68 163.367
R1596 B.n1313 B.n68 163.367
R1597 B.n1313 B.n73 163.367
R1598 B.n1309 B.n73 163.367
R1599 B.n1309 B.n75 163.367
R1600 B.n1305 B.n75 163.367
R1601 B.n1305 B.n80 163.367
R1602 B.n1301 B.n80 163.367
R1603 B.n1301 B.n82 163.367
R1604 B.n1297 B.n82 163.367
R1605 B.n1297 B.n87 163.367
R1606 B.n1293 B.n87 163.367
R1607 B.n1293 B.n89 163.367
R1608 B.n1289 B.n89 163.367
R1609 B.n1289 B.n94 163.367
R1610 B.n1285 B.n94 163.367
R1611 B.n1285 B.n96 163.367
R1612 B.n1281 B.n96 163.367
R1613 B.n1281 B.n101 163.367
R1614 B.n1277 B.n101 163.367
R1615 B.n1277 B.n103 163.367
R1616 B.n1273 B.n103 163.367
R1617 B.n1273 B.n108 163.367
R1618 B.n1269 B.n108 163.367
R1619 B.n1269 B.n110 163.367
R1620 B.n1265 B.n110 163.367
R1621 B.n1265 B.n115 163.367
R1622 B.n1261 B.n115 163.367
R1623 B.n1261 B.n117 163.367
R1624 B.n1257 B.n117 163.367
R1625 B.n1257 B.n121 163.367
R1626 B.n1253 B.n121 163.367
R1627 B.n1253 B.n123 163.367
R1628 B.n1249 B.n123 163.367
R1629 B.n1249 B.n129 163.367
R1630 B.n1245 B.n129 163.367
R1631 B.n1245 B.n131 163.367
R1632 B.n1241 B.n131 163.367
R1633 B.n1241 B.n136 163.367
R1634 B.n1237 B.n136 163.367
R1635 B.n201 B.t22 142.754
R1636 B.n786 B.t13 142.754
R1637 B.n204 B.t16 142.731
R1638 B.n628 B.t20 142.731
R1639 B.n205 B.n204 75.0551
R1640 B.n202 B.n201 75.0551
R1641 B.n787 B.n786 75.0551
R1642 B.n629 B.n628 75.0551
R1643 B.n140 B.n138 71.676
R1644 B.n209 B.n141 71.676
R1645 B.n213 B.n142 71.676
R1646 B.n217 B.n143 71.676
R1647 B.n221 B.n144 71.676
R1648 B.n225 B.n145 71.676
R1649 B.n229 B.n146 71.676
R1650 B.n233 B.n147 71.676
R1651 B.n237 B.n148 71.676
R1652 B.n241 B.n149 71.676
R1653 B.n245 B.n150 71.676
R1654 B.n249 B.n151 71.676
R1655 B.n253 B.n152 71.676
R1656 B.n257 B.n153 71.676
R1657 B.n261 B.n154 71.676
R1658 B.n265 B.n155 71.676
R1659 B.n269 B.n156 71.676
R1660 B.n273 B.n157 71.676
R1661 B.n277 B.n158 71.676
R1662 B.n281 B.n159 71.676
R1663 B.n285 B.n160 71.676
R1664 B.n289 B.n161 71.676
R1665 B.n293 B.n162 71.676
R1666 B.n297 B.n163 71.676
R1667 B.n301 B.n164 71.676
R1668 B.n305 B.n165 71.676
R1669 B.n309 B.n166 71.676
R1670 B.n313 B.n167 71.676
R1671 B.n317 B.n168 71.676
R1672 B.n321 B.n169 71.676
R1673 B.n325 B.n170 71.676
R1674 B.n329 B.n171 71.676
R1675 B.n333 B.n172 71.676
R1676 B.n337 B.n173 71.676
R1677 B.n341 B.n174 71.676
R1678 B.n345 B.n175 71.676
R1679 B.n349 B.n176 71.676
R1680 B.n353 B.n177 71.676
R1681 B.n357 B.n178 71.676
R1682 B.n361 B.n179 71.676
R1683 B.n365 B.n180 71.676
R1684 B.n369 B.n181 71.676
R1685 B.n373 B.n182 71.676
R1686 B.n377 B.n183 71.676
R1687 B.n381 B.n184 71.676
R1688 B.n385 B.n185 71.676
R1689 B.n389 B.n186 71.676
R1690 B.n393 B.n187 71.676
R1691 B.n397 B.n188 71.676
R1692 B.n401 B.n189 71.676
R1693 B.n405 B.n190 71.676
R1694 B.n409 B.n191 71.676
R1695 B.n413 B.n192 71.676
R1696 B.n417 B.n193 71.676
R1697 B.n421 B.n194 71.676
R1698 B.n425 B.n195 71.676
R1699 B.n429 B.n196 71.676
R1700 B.n433 B.n197 71.676
R1701 B.n437 B.n198 71.676
R1702 B.n441 B.n199 71.676
R1703 B.n1234 B.n200 71.676
R1704 B.n1234 B.n1233 71.676
R1705 B.n443 B.n199 71.676
R1706 B.n440 B.n198 71.676
R1707 B.n436 B.n197 71.676
R1708 B.n432 B.n196 71.676
R1709 B.n428 B.n195 71.676
R1710 B.n424 B.n194 71.676
R1711 B.n420 B.n193 71.676
R1712 B.n416 B.n192 71.676
R1713 B.n412 B.n191 71.676
R1714 B.n408 B.n190 71.676
R1715 B.n404 B.n189 71.676
R1716 B.n400 B.n188 71.676
R1717 B.n396 B.n187 71.676
R1718 B.n392 B.n186 71.676
R1719 B.n388 B.n185 71.676
R1720 B.n384 B.n184 71.676
R1721 B.n380 B.n183 71.676
R1722 B.n376 B.n182 71.676
R1723 B.n372 B.n181 71.676
R1724 B.n368 B.n180 71.676
R1725 B.n364 B.n179 71.676
R1726 B.n360 B.n178 71.676
R1727 B.n356 B.n177 71.676
R1728 B.n352 B.n176 71.676
R1729 B.n348 B.n175 71.676
R1730 B.n344 B.n174 71.676
R1731 B.n340 B.n173 71.676
R1732 B.n336 B.n172 71.676
R1733 B.n332 B.n171 71.676
R1734 B.n328 B.n170 71.676
R1735 B.n324 B.n169 71.676
R1736 B.n320 B.n168 71.676
R1737 B.n316 B.n167 71.676
R1738 B.n312 B.n166 71.676
R1739 B.n308 B.n165 71.676
R1740 B.n304 B.n164 71.676
R1741 B.n300 B.n163 71.676
R1742 B.n296 B.n162 71.676
R1743 B.n292 B.n161 71.676
R1744 B.n288 B.n160 71.676
R1745 B.n284 B.n159 71.676
R1746 B.n280 B.n158 71.676
R1747 B.n276 B.n157 71.676
R1748 B.n272 B.n156 71.676
R1749 B.n268 B.n155 71.676
R1750 B.n264 B.n154 71.676
R1751 B.n260 B.n153 71.676
R1752 B.n256 B.n152 71.676
R1753 B.n252 B.n151 71.676
R1754 B.n248 B.n150 71.676
R1755 B.n244 B.n149 71.676
R1756 B.n240 B.n148 71.676
R1757 B.n236 B.n147 71.676
R1758 B.n232 B.n146 71.676
R1759 B.n228 B.n145 71.676
R1760 B.n224 B.n144 71.676
R1761 B.n220 B.n143 71.676
R1762 B.n216 B.n142 71.676
R1763 B.n212 B.n141 71.676
R1764 B.n208 B.n140 71.676
R1765 B.n658 B.n592 71.676
R1766 B.n662 B.n661 71.676
R1767 B.n667 B.n666 71.676
R1768 B.n670 B.n669 71.676
R1769 B.n675 B.n674 71.676
R1770 B.n678 B.n677 71.676
R1771 B.n683 B.n682 71.676
R1772 B.n686 B.n685 71.676
R1773 B.n691 B.n690 71.676
R1774 B.n694 B.n693 71.676
R1775 B.n699 B.n698 71.676
R1776 B.n702 B.n701 71.676
R1777 B.n707 B.n706 71.676
R1778 B.n710 B.n709 71.676
R1779 B.n715 B.n714 71.676
R1780 B.n718 B.n717 71.676
R1781 B.n723 B.n722 71.676
R1782 B.n726 B.n725 71.676
R1783 B.n731 B.n730 71.676
R1784 B.n734 B.n733 71.676
R1785 B.n739 B.n738 71.676
R1786 B.n742 B.n741 71.676
R1787 B.n747 B.n746 71.676
R1788 B.n750 B.n749 71.676
R1789 B.n755 B.n754 71.676
R1790 B.n758 B.n757 71.676
R1791 B.n763 B.n762 71.676
R1792 B.n766 B.n765 71.676
R1793 B.n772 B.n771 71.676
R1794 B.n775 B.n774 71.676
R1795 B.n780 B.n779 71.676
R1796 B.n783 B.n782 71.676
R1797 B.n791 B.n790 71.676
R1798 B.n794 B.n793 71.676
R1799 B.n799 B.n798 71.676
R1800 B.n802 B.n801 71.676
R1801 B.n807 B.n806 71.676
R1802 B.n810 B.n809 71.676
R1803 B.n815 B.n814 71.676
R1804 B.n818 B.n817 71.676
R1805 B.n823 B.n822 71.676
R1806 B.n826 B.n825 71.676
R1807 B.n831 B.n830 71.676
R1808 B.n834 B.n833 71.676
R1809 B.n839 B.n838 71.676
R1810 B.n842 B.n841 71.676
R1811 B.n847 B.n846 71.676
R1812 B.n850 B.n849 71.676
R1813 B.n855 B.n854 71.676
R1814 B.n858 B.n857 71.676
R1815 B.n863 B.n862 71.676
R1816 B.n866 B.n865 71.676
R1817 B.n871 B.n870 71.676
R1818 B.n874 B.n873 71.676
R1819 B.n879 B.n878 71.676
R1820 B.n882 B.n881 71.676
R1821 B.n887 B.n886 71.676
R1822 B.n890 B.n889 71.676
R1823 B.n895 B.n894 71.676
R1824 B.n898 B.n897 71.676
R1825 B.n659 B.n658 71.676
R1826 B.n661 B.n655 71.676
R1827 B.n668 B.n667 71.676
R1828 B.n669 B.n653 71.676
R1829 B.n676 B.n675 71.676
R1830 B.n677 B.n651 71.676
R1831 B.n684 B.n683 71.676
R1832 B.n685 B.n649 71.676
R1833 B.n692 B.n691 71.676
R1834 B.n693 B.n647 71.676
R1835 B.n700 B.n699 71.676
R1836 B.n701 B.n645 71.676
R1837 B.n708 B.n707 71.676
R1838 B.n709 B.n643 71.676
R1839 B.n716 B.n715 71.676
R1840 B.n717 B.n641 71.676
R1841 B.n724 B.n723 71.676
R1842 B.n725 B.n639 71.676
R1843 B.n732 B.n731 71.676
R1844 B.n733 B.n637 71.676
R1845 B.n740 B.n739 71.676
R1846 B.n741 B.n635 71.676
R1847 B.n748 B.n747 71.676
R1848 B.n749 B.n633 71.676
R1849 B.n756 B.n755 71.676
R1850 B.n757 B.n631 71.676
R1851 B.n764 B.n763 71.676
R1852 B.n765 B.n627 71.676
R1853 B.n773 B.n772 71.676
R1854 B.n774 B.n625 71.676
R1855 B.n781 B.n780 71.676
R1856 B.n782 B.n623 71.676
R1857 B.n792 B.n791 71.676
R1858 B.n793 B.n621 71.676
R1859 B.n800 B.n799 71.676
R1860 B.n801 B.n619 71.676
R1861 B.n808 B.n807 71.676
R1862 B.n809 B.n617 71.676
R1863 B.n816 B.n815 71.676
R1864 B.n817 B.n615 71.676
R1865 B.n824 B.n823 71.676
R1866 B.n825 B.n613 71.676
R1867 B.n832 B.n831 71.676
R1868 B.n833 B.n611 71.676
R1869 B.n840 B.n839 71.676
R1870 B.n841 B.n609 71.676
R1871 B.n848 B.n847 71.676
R1872 B.n849 B.n607 71.676
R1873 B.n856 B.n855 71.676
R1874 B.n857 B.n605 71.676
R1875 B.n864 B.n863 71.676
R1876 B.n865 B.n603 71.676
R1877 B.n872 B.n871 71.676
R1878 B.n873 B.n601 71.676
R1879 B.n880 B.n879 71.676
R1880 B.n881 B.n599 71.676
R1881 B.n888 B.n887 71.676
R1882 B.n889 B.n597 71.676
R1883 B.n896 B.n895 71.676
R1884 B.n899 B.n898 71.676
R1885 B.n1391 B.n1390 71.676
R1886 B.n1391 B.n2 71.676
R1887 B.n202 B.t23 67.6986
R1888 B.n787 B.t12 67.6986
R1889 B.n205 B.t17 67.6759
R1890 B.n629 B.t19 67.6759
R1891 B.n206 B.n205 59.5399
R1892 B.n203 B.n202 59.5399
R1893 B.n788 B.n787 59.5399
R1894 B.n768 B.n629 59.5399
R1895 B.n904 B.n593 57.7264
R1896 B.n1236 B.n1235 57.7264
R1897 B.n904 B.n589 33.5506
R1898 B.n910 B.n589 33.5506
R1899 B.n910 B.n585 33.5506
R1900 B.n916 B.n585 33.5506
R1901 B.n916 B.n581 33.5506
R1902 B.n922 B.n581 33.5506
R1903 B.n922 B.n577 33.5506
R1904 B.n929 B.n577 33.5506
R1905 B.n929 B.n928 33.5506
R1906 B.n935 B.n570 33.5506
R1907 B.n941 B.n570 33.5506
R1908 B.n941 B.n566 33.5506
R1909 B.n947 B.n566 33.5506
R1910 B.n947 B.n562 33.5506
R1911 B.n953 B.n562 33.5506
R1912 B.n953 B.n558 33.5506
R1913 B.n959 B.n558 33.5506
R1914 B.n959 B.n554 33.5506
R1915 B.n965 B.n554 33.5506
R1916 B.n965 B.n549 33.5506
R1917 B.n971 B.n549 33.5506
R1918 B.n971 B.n550 33.5506
R1919 B.n977 B.n542 33.5506
R1920 B.n983 B.n542 33.5506
R1921 B.n983 B.n538 33.5506
R1922 B.n989 B.n538 33.5506
R1923 B.n989 B.n534 33.5506
R1924 B.n995 B.n534 33.5506
R1925 B.n995 B.n530 33.5506
R1926 B.n1001 B.n530 33.5506
R1927 B.n1001 B.n525 33.5506
R1928 B.n1007 B.n525 33.5506
R1929 B.n1007 B.n526 33.5506
R1930 B.n1013 B.n518 33.5506
R1931 B.n1019 B.n518 33.5506
R1932 B.n1019 B.n514 33.5506
R1933 B.n1025 B.n514 33.5506
R1934 B.n1025 B.n510 33.5506
R1935 B.n1031 B.n510 33.5506
R1936 B.n1031 B.n506 33.5506
R1937 B.n1037 B.n506 33.5506
R1938 B.n1037 B.n502 33.5506
R1939 B.n1043 B.n502 33.5506
R1940 B.n1049 B.n498 33.5506
R1941 B.n1049 B.n494 33.5506
R1942 B.n1055 B.n494 33.5506
R1943 B.n1055 B.n490 33.5506
R1944 B.n1061 B.n490 33.5506
R1945 B.n1061 B.n486 33.5506
R1946 B.n1067 B.n486 33.5506
R1947 B.n1067 B.n482 33.5506
R1948 B.n1074 B.n482 33.5506
R1949 B.n1074 B.n1073 33.5506
R1950 B.n1080 B.n475 33.5506
R1951 B.n1086 B.n475 33.5506
R1952 B.n1086 B.n471 33.5506
R1953 B.n1092 B.n471 33.5506
R1954 B.n1092 B.n467 33.5506
R1955 B.n1098 B.n467 33.5506
R1956 B.n1098 B.n463 33.5506
R1957 B.n1104 B.n463 33.5506
R1958 B.n1104 B.n459 33.5506
R1959 B.n1111 B.n459 33.5506
R1960 B.n1111 B.n1110 33.5506
R1961 B.n1117 B.n452 33.5506
R1962 B.n1124 B.n452 33.5506
R1963 B.n1124 B.n448 33.5506
R1964 B.n1130 B.n448 33.5506
R1965 B.n1130 B.n4 33.5506
R1966 B.n1389 B.n4 33.5506
R1967 B.n1389 B.n1388 33.5506
R1968 B.n1388 B.n1387 33.5506
R1969 B.n1387 B.n8 33.5506
R1970 B.n12 B.n8 33.5506
R1971 B.n1380 B.n12 33.5506
R1972 B.n1380 B.n1379 33.5506
R1973 B.n1379 B.n1378 33.5506
R1974 B.n1372 B.n19 33.5506
R1975 B.n1372 B.n1371 33.5506
R1976 B.n1371 B.n1370 33.5506
R1977 B.n1370 B.n23 33.5506
R1978 B.n1364 B.n23 33.5506
R1979 B.n1364 B.n1363 33.5506
R1980 B.n1363 B.n1362 33.5506
R1981 B.n1362 B.n30 33.5506
R1982 B.n1356 B.n30 33.5506
R1983 B.n1356 B.n1355 33.5506
R1984 B.n1355 B.n1354 33.5506
R1985 B.n1348 B.n40 33.5506
R1986 B.n1348 B.n1347 33.5506
R1987 B.n1347 B.n1346 33.5506
R1988 B.n1346 B.n44 33.5506
R1989 B.n1340 B.n44 33.5506
R1990 B.n1340 B.n1339 33.5506
R1991 B.n1339 B.n1338 33.5506
R1992 B.n1338 B.n51 33.5506
R1993 B.n1332 B.n51 33.5506
R1994 B.n1332 B.n1331 33.5506
R1995 B.n1330 B.n58 33.5506
R1996 B.n1324 B.n58 33.5506
R1997 B.n1324 B.n1323 33.5506
R1998 B.n1323 B.n1322 33.5506
R1999 B.n1322 B.n65 33.5506
R2000 B.n1316 B.n65 33.5506
R2001 B.n1316 B.n1315 33.5506
R2002 B.n1315 B.n1314 33.5506
R2003 B.n1314 B.n72 33.5506
R2004 B.n1308 B.n72 33.5506
R2005 B.n1307 B.n1306 33.5506
R2006 B.n1306 B.n79 33.5506
R2007 B.n1300 B.n79 33.5506
R2008 B.n1300 B.n1299 33.5506
R2009 B.n1299 B.n1298 33.5506
R2010 B.n1298 B.n86 33.5506
R2011 B.n1292 B.n86 33.5506
R2012 B.n1292 B.n1291 33.5506
R2013 B.n1291 B.n1290 33.5506
R2014 B.n1290 B.n93 33.5506
R2015 B.n1284 B.n93 33.5506
R2016 B.n1283 B.n1282 33.5506
R2017 B.n1282 B.n100 33.5506
R2018 B.n1276 B.n100 33.5506
R2019 B.n1276 B.n1275 33.5506
R2020 B.n1275 B.n1274 33.5506
R2021 B.n1274 B.n107 33.5506
R2022 B.n1268 B.n107 33.5506
R2023 B.n1268 B.n1267 33.5506
R2024 B.n1267 B.n1266 33.5506
R2025 B.n1266 B.n114 33.5506
R2026 B.n1260 B.n114 33.5506
R2027 B.n1260 B.n1259 33.5506
R2028 B.n1259 B.n1258 33.5506
R2029 B.n1252 B.n124 33.5506
R2030 B.n1252 B.n1251 33.5506
R2031 B.n1251 B.n1250 33.5506
R2032 B.n1250 B.n128 33.5506
R2033 B.n1244 B.n128 33.5506
R2034 B.n1244 B.n1243 33.5506
R2035 B.n1243 B.n1242 33.5506
R2036 B.n1242 B.n135 33.5506
R2037 B.n1236 B.n135 33.5506
R2038 B.n906 B.n591 33.2493
R2039 B.n902 B.n901 33.2493
R2040 B.n1232 B.n1231 33.2493
R2041 B.n1238 B.n137 33.2493
R2042 B.n1013 B.t2 31.5771
R2043 B.n1308 B.t6 31.5771
R2044 B.n935 B.t11 30.5903
R2045 B.n1258 B.t15 30.5903
R2046 B.n1073 B.t8 27.63
R2047 B.n40 B.t1 27.63
R2048 B.n1117 B.t5 26.6432
R2049 B.n1378 B.t0 26.6432
R2050 B.n550 B.t3 22.6962
R2051 B.t9 B.n1283 22.6962
R2052 B.t7 B.n498 18.7491
R2053 B.n1331 B.t4 18.7491
R2054 B B.n1392 18.0485
R2055 B.n1043 B.t7 14.802
R2056 B.t4 B.n1330 14.802
R2057 B.n977 B.t3 10.855
R2058 B.n1284 B.t9 10.855
R2059 B.n907 B.n906 10.6151
R2060 B.n908 B.n907 10.6151
R2061 B.n908 B.n583 10.6151
R2062 B.n918 B.n583 10.6151
R2063 B.n919 B.n918 10.6151
R2064 B.n920 B.n919 10.6151
R2065 B.n920 B.n575 10.6151
R2066 B.n931 B.n575 10.6151
R2067 B.n932 B.n931 10.6151
R2068 B.n933 B.n932 10.6151
R2069 B.n933 B.n568 10.6151
R2070 B.n943 B.n568 10.6151
R2071 B.n944 B.n943 10.6151
R2072 B.n945 B.n944 10.6151
R2073 B.n945 B.n560 10.6151
R2074 B.n955 B.n560 10.6151
R2075 B.n956 B.n955 10.6151
R2076 B.n957 B.n956 10.6151
R2077 B.n957 B.n552 10.6151
R2078 B.n967 B.n552 10.6151
R2079 B.n968 B.n967 10.6151
R2080 B.n969 B.n968 10.6151
R2081 B.n969 B.n544 10.6151
R2082 B.n979 B.n544 10.6151
R2083 B.n980 B.n979 10.6151
R2084 B.n981 B.n980 10.6151
R2085 B.n981 B.n536 10.6151
R2086 B.n991 B.n536 10.6151
R2087 B.n992 B.n991 10.6151
R2088 B.n993 B.n992 10.6151
R2089 B.n993 B.n528 10.6151
R2090 B.n1003 B.n528 10.6151
R2091 B.n1004 B.n1003 10.6151
R2092 B.n1005 B.n1004 10.6151
R2093 B.n1005 B.n520 10.6151
R2094 B.n1015 B.n520 10.6151
R2095 B.n1016 B.n1015 10.6151
R2096 B.n1017 B.n1016 10.6151
R2097 B.n1017 B.n512 10.6151
R2098 B.n1027 B.n512 10.6151
R2099 B.n1028 B.n1027 10.6151
R2100 B.n1029 B.n1028 10.6151
R2101 B.n1029 B.n504 10.6151
R2102 B.n1039 B.n504 10.6151
R2103 B.n1040 B.n1039 10.6151
R2104 B.n1041 B.n1040 10.6151
R2105 B.n1041 B.n496 10.6151
R2106 B.n1051 B.n496 10.6151
R2107 B.n1052 B.n1051 10.6151
R2108 B.n1053 B.n1052 10.6151
R2109 B.n1053 B.n488 10.6151
R2110 B.n1063 B.n488 10.6151
R2111 B.n1064 B.n1063 10.6151
R2112 B.n1065 B.n1064 10.6151
R2113 B.n1065 B.n480 10.6151
R2114 B.n1076 B.n480 10.6151
R2115 B.n1077 B.n1076 10.6151
R2116 B.n1078 B.n1077 10.6151
R2117 B.n1078 B.n473 10.6151
R2118 B.n1088 B.n473 10.6151
R2119 B.n1089 B.n1088 10.6151
R2120 B.n1090 B.n1089 10.6151
R2121 B.n1090 B.n465 10.6151
R2122 B.n1100 B.n465 10.6151
R2123 B.n1101 B.n1100 10.6151
R2124 B.n1102 B.n1101 10.6151
R2125 B.n1102 B.n457 10.6151
R2126 B.n1113 B.n457 10.6151
R2127 B.n1114 B.n1113 10.6151
R2128 B.n1115 B.n1114 10.6151
R2129 B.n1115 B.n450 10.6151
R2130 B.n1126 B.n450 10.6151
R2131 B.n1127 B.n1126 10.6151
R2132 B.n1128 B.n1127 10.6151
R2133 B.n1128 B.n0 10.6151
R2134 B.n657 B.n591 10.6151
R2135 B.n657 B.n656 10.6151
R2136 B.n663 B.n656 10.6151
R2137 B.n664 B.n663 10.6151
R2138 B.n665 B.n664 10.6151
R2139 B.n665 B.n654 10.6151
R2140 B.n671 B.n654 10.6151
R2141 B.n672 B.n671 10.6151
R2142 B.n673 B.n672 10.6151
R2143 B.n673 B.n652 10.6151
R2144 B.n679 B.n652 10.6151
R2145 B.n680 B.n679 10.6151
R2146 B.n681 B.n680 10.6151
R2147 B.n681 B.n650 10.6151
R2148 B.n687 B.n650 10.6151
R2149 B.n688 B.n687 10.6151
R2150 B.n689 B.n688 10.6151
R2151 B.n689 B.n648 10.6151
R2152 B.n695 B.n648 10.6151
R2153 B.n696 B.n695 10.6151
R2154 B.n697 B.n696 10.6151
R2155 B.n697 B.n646 10.6151
R2156 B.n703 B.n646 10.6151
R2157 B.n704 B.n703 10.6151
R2158 B.n705 B.n704 10.6151
R2159 B.n705 B.n644 10.6151
R2160 B.n711 B.n644 10.6151
R2161 B.n712 B.n711 10.6151
R2162 B.n713 B.n712 10.6151
R2163 B.n713 B.n642 10.6151
R2164 B.n719 B.n642 10.6151
R2165 B.n720 B.n719 10.6151
R2166 B.n721 B.n720 10.6151
R2167 B.n721 B.n640 10.6151
R2168 B.n727 B.n640 10.6151
R2169 B.n728 B.n727 10.6151
R2170 B.n729 B.n728 10.6151
R2171 B.n729 B.n638 10.6151
R2172 B.n735 B.n638 10.6151
R2173 B.n736 B.n735 10.6151
R2174 B.n737 B.n736 10.6151
R2175 B.n737 B.n636 10.6151
R2176 B.n743 B.n636 10.6151
R2177 B.n744 B.n743 10.6151
R2178 B.n745 B.n744 10.6151
R2179 B.n745 B.n634 10.6151
R2180 B.n751 B.n634 10.6151
R2181 B.n752 B.n751 10.6151
R2182 B.n753 B.n752 10.6151
R2183 B.n753 B.n632 10.6151
R2184 B.n759 B.n632 10.6151
R2185 B.n760 B.n759 10.6151
R2186 B.n761 B.n760 10.6151
R2187 B.n761 B.n630 10.6151
R2188 B.n767 B.n630 10.6151
R2189 B.n770 B.n769 10.6151
R2190 B.n770 B.n626 10.6151
R2191 B.n776 B.n626 10.6151
R2192 B.n777 B.n776 10.6151
R2193 B.n778 B.n777 10.6151
R2194 B.n778 B.n624 10.6151
R2195 B.n784 B.n624 10.6151
R2196 B.n785 B.n784 10.6151
R2197 B.n789 B.n785 10.6151
R2198 B.n795 B.n622 10.6151
R2199 B.n796 B.n795 10.6151
R2200 B.n797 B.n796 10.6151
R2201 B.n797 B.n620 10.6151
R2202 B.n803 B.n620 10.6151
R2203 B.n804 B.n803 10.6151
R2204 B.n805 B.n804 10.6151
R2205 B.n805 B.n618 10.6151
R2206 B.n811 B.n618 10.6151
R2207 B.n812 B.n811 10.6151
R2208 B.n813 B.n812 10.6151
R2209 B.n813 B.n616 10.6151
R2210 B.n819 B.n616 10.6151
R2211 B.n820 B.n819 10.6151
R2212 B.n821 B.n820 10.6151
R2213 B.n821 B.n614 10.6151
R2214 B.n827 B.n614 10.6151
R2215 B.n828 B.n827 10.6151
R2216 B.n829 B.n828 10.6151
R2217 B.n829 B.n612 10.6151
R2218 B.n835 B.n612 10.6151
R2219 B.n836 B.n835 10.6151
R2220 B.n837 B.n836 10.6151
R2221 B.n837 B.n610 10.6151
R2222 B.n843 B.n610 10.6151
R2223 B.n844 B.n843 10.6151
R2224 B.n845 B.n844 10.6151
R2225 B.n845 B.n608 10.6151
R2226 B.n851 B.n608 10.6151
R2227 B.n852 B.n851 10.6151
R2228 B.n853 B.n852 10.6151
R2229 B.n853 B.n606 10.6151
R2230 B.n859 B.n606 10.6151
R2231 B.n860 B.n859 10.6151
R2232 B.n861 B.n860 10.6151
R2233 B.n861 B.n604 10.6151
R2234 B.n867 B.n604 10.6151
R2235 B.n868 B.n867 10.6151
R2236 B.n869 B.n868 10.6151
R2237 B.n869 B.n602 10.6151
R2238 B.n875 B.n602 10.6151
R2239 B.n876 B.n875 10.6151
R2240 B.n877 B.n876 10.6151
R2241 B.n877 B.n600 10.6151
R2242 B.n883 B.n600 10.6151
R2243 B.n884 B.n883 10.6151
R2244 B.n885 B.n884 10.6151
R2245 B.n885 B.n598 10.6151
R2246 B.n891 B.n598 10.6151
R2247 B.n892 B.n891 10.6151
R2248 B.n893 B.n892 10.6151
R2249 B.n893 B.n596 10.6151
R2250 B.n596 B.n595 10.6151
R2251 B.n900 B.n595 10.6151
R2252 B.n901 B.n900 10.6151
R2253 B.n902 B.n587 10.6151
R2254 B.n912 B.n587 10.6151
R2255 B.n913 B.n912 10.6151
R2256 B.n914 B.n913 10.6151
R2257 B.n914 B.n579 10.6151
R2258 B.n924 B.n579 10.6151
R2259 B.n925 B.n924 10.6151
R2260 B.n926 B.n925 10.6151
R2261 B.n926 B.n572 10.6151
R2262 B.n937 B.n572 10.6151
R2263 B.n938 B.n937 10.6151
R2264 B.n939 B.n938 10.6151
R2265 B.n939 B.n564 10.6151
R2266 B.n949 B.n564 10.6151
R2267 B.n950 B.n949 10.6151
R2268 B.n951 B.n950 10.6151
R2269 B.n951 B.n556 10.6151
R2270 B.n961 B.n556 10.6151
R2271 B.n962 B.n961 10.6151
R2272 B.n963 B.n962 10.6151
R2273 B.n963 B.n547 10.6151
R2274 B.n973 B.n547 10.6151
R2275 B.n974 B.n973 10.6151
R2276 B.n975 B.n974 10.6151
R2277 B.n975 B.n540 10.6151
R2278 B.n985 B.n540 10.6151
R2279 B.n986 B.n985 10.6151
R2280 B.n987 B.n986 10.6151
R2281 B.n987 B.n532 10.6151
R2282 B.n997 B.n532 10.6151
R2283 B.n998 B.n997 10.6151
R2284 B.n999 B.n998 10.6151
R2285 B.n999 B.n523 10.6151
R2286 B.n1009 B.n523 10.6151
R2287 B.n1010 B.n1009 10.6151
R2288 B.n1011 B.n1010 10.6151
R2289 B.n1011 B.n516 10.6151
R2290 B.n1021 B.n516 10.6151
R2291 B.n1022 B.n1021 10.6151
R2292 B.n1023 B.n1022 10.6151
R2293 B.n1023 B.n508 10.6151
R2294 B.n1033 B.n508 10.6151
R2295 B.n1034 B.n1033 10.6151
R2296 B.n1035 B.n1034 10.6151
R2297 B.n1035 B.n500 10.6151
R2298 B.n1045 B.n500 10.6151
R2299 B.n1046 B.n1045 10.6151
R2300 B.n1047 B.n1046 10.6151
R2301 B.n1047 B.n492 10.6151
R2302 B.n1057 B.n492 10.6151
R2303 B.n1058 B.n1057 10.6151
R2304 B.n1059 B.n1058 10.6151
R2305 B.n1059 B.n484 10.6151
R2306 B.n1069 B.n484 10.6151
R2307 B.n1070 B.n1069 10.6151
R2308 B.n1071 B.n1070 10.6151
R2309 B.n1071 B.n477 10.6151
R2310 B.n1082 B.n477 10.6151
R2311 B.n1083 B.n1082 10.6151
R2312 B.n1084 B.n1083 10.6151
R2313 B.n1084 B.n469 10.6151
R2314 B.n1094 B.n469 10.6151
R2315 B.n1095 B.n1094 10.6151
R2316 B.n1096 B.n1095 10.6151
R2317 B.n1096 B.n461 10.6151
R2318 B.n1106 B.n461 10.6151
R2319 B.n1107 B.n1106 10.6151
R2320 B.n1108 B.n1107 10.6151
R2321 B.n1108 B.n454 10.6151
R2322 B.n1119 B.n454 10.6151
R2323 B.n1120 B.n1119 10.6151
R2324 B.n1122 B.n1120 10.6151
R2325 B.n1122 B.n1121 10.6151
R2326 B.n1121 B.n446 10.6151
R2327 B.n1133 B.n446 10.6151
R2328 B.n1134 B.n1133 10.6151
R2329 B.n1135 B.n1134 10.6151
R2330 B.n1136 B.n1135 10.6151
R2331 B.n1137 B.n1136 10.6151
R2332 B.n1140 B.n1137 10.6151
R2333 B.n1141 B.n1140 10.6151
R2334 B.n1142 B.n1141 10.6151
R2335 B.n1143 B.n1142 10.6151
R2336 B.n1145 B.n1143 10.6151
R2337 B.n1146 B.n1145 10.6151
R2338 B.n1147 B.n1146 10.6151
R2339 B.n1148 B.n1147 10.6151
R2340 B.n1150 B.n1148 10.6151
R2341 B.n1151 B.n1150 10.6151
R2342 B.n1152 B.n1151 10.6151
R2343 B.n1153 B.n1152 10.6151
R2344 B.n1155 B.n1153 10.6151
R2345 B.n1156 B.n1155 10.6151
R2346 B.n1157 B.n1156 10.6151
R2347 B.n1158 B.n1157 10.6151
R2348 B.n1160 B.n1158 10.6151
R2349 B.n1161 B.n1160 10.6151
R2350 B.n1162 B.n1161 10.6151
R2351 B.n1163 B.n1162 10.6151
R2352 B.n1165 B.n1163 10.6151
R2353 B.n1166 B.n1165 10.6151
R2354 B.n1167 B.n1166 10.6151
R2355 B.n1168 B.n1167 10.6151
R2356 B.n1170 B.n1168 10.6151
R2357 B.n1171 B.n1170 10.6151
R2358 B.n1172 B.n1171 10.6151
R2359 B.n1173 B.n1172 10.6151
R2360 B.n1175 B.n1173 10.6151
R2361 B.n1176 B.n1175 10.6151
R2362 B.n1177 B.n1176 10.6151
R2363 B.n1178 B.n1177 10.6151
R2364 B.n1180 B.n1178 10.6151
R2365 B.n1181 B.n1180 10.6151
R2366 B.n1182 B.n1181 10.6151
R2367 B.n1183 B.n1182 10.6151
R2368 B.n1185 B.n1183 10.6151
R2369 B.n1186 B.n1185 10.6151
R2370 B.n1187 B.n1186 10.6151
R2371 B.n1188 B.n1187 10.6151
R2372 B.n1190 B.n1188 10.6151
R2373 B.n1191 B.n1190 10.6151
R2374 B.n1192 B.n1191 10.6151
R2375 B.n1193 B.n1192 10.6151
R2376 B.n1195 B.n1193 10.6151
R2377 B.n1196 B.n1195 10.6151
R2378 B.n1197 B.n1196 10.6151
R2379 B.n1198 B.n1197 10.6151
R2380 B.n1200 B.n1198 10.6151
R2381 B.n1201 B.n1200 10.6151
R2382 B.n1202 B.n1201 10.6151
R2383 B.n1203 B.n1202 10.6151
R2384 B.n1205 B.n1203 10.6151
R2385 B.n1206 B.n1205 10.6151
R2386 B.n1207 B.n1206 10.6151
R2387 B.n1208 B.n1207 10.6151
R2388 B.n1210 B.n1208 10.6151
R2389 B.n1211 B.n1210 10.6151
R2390 B.n1212 B.n1211 10.6151
R2391 B.n1213 B.n1212 10.6151
R2392 B.n1215 B.n1213 10.6151
R2393 B.n1216 B.n1215 10.6151
R2394 B.n1217 B.n1216 10.6151
R2395 B.n1218 B.n1217 10.6151
R2396 B.n1220 B.n1218 10.6151
R2397 B.n1221 B.n1220 10.6151
R2398 B.n1222 B.n1221 10.6151
R2399 B.n1223 B.n1222 10.6151
R2400 B.n1225 B.n1223 10.6151
R2401 B.n1226 B.n1225 10.6151
R2402 B.n1227 B.n1226 10.6151
R2403 B.n1228 B.n1227 10.6151
R2404 B.n1230 B.n1228 10.6151
R2405 B.n1231 B.n1230 10.6151
R2406 B.n1384 B.n1 10.6151
R2407 B.n1384 B.n1383 10.6151
R2408 B.n1383 B.n1382 10.6151
R2409 B.n1382 B.n10 10.6151
R2410 B.n1376 B.n10 10.6151
R2411 B.n1376 B.n1375 10.6151
R2412 B.n1375 B.n1374 10.6151
R2413 B.n1374 B.n17 10.6151
R2414 B.n1368 B.n17 10.6151
R2415 B.n1368 B.n1367 10.6151
R2416 B.n1367 B.n1366 10.6151
R2417 B.n1366 B.n25 10.6151
R2418 B.n1360 B.n25 10.6151
R2419 B.n1360 B.n1359 10.6151
R2420 B.n1359 B.n1358 10.6151
R2421 B.n1358 B.n32 10.6151
R2422 B.n1352 B.n32 10.6151
R2423 B.n1352 B.n1351 10.6151
R2424 B.n1351 B.n1350 10.6151
R2425 B.n1350 B.n38 10.6151
R2426 B.n1344 B.n38 10.6151
R2427 B.n1344 B.n1343 10.6151
R2428 B.n1343 B.n1342 10.6151
R2429 B.n1342 B.n46 10.6151
R2430 B.n1336 B.n46 10.6151
R2431 B.n1336 B.n1335 10.6151
R2432 B.n1335 B.n1334 10.6151
R2433 B.n1334 B.n53 10.6151
R2434 B.n1328 B.n53 10.6151
R2435 B.n1328 B.n1327 10.6151
R2436 B.n1327 B.n1326 10.6151
R2437 B.n1326 B.n60 10.6151
R2438 B.n1320 B.n60 10.6151
R2439 B.n1320 B.n1319 10.6151
R2440 B.n1319 B.n1318 10.6151
R2441 B.n1318 B.n67 10.6151
R2442 B.n1312 B.n67 10.6151
R2443 B.n1312 B.n1311 10.6151
R2444 B.n1311 B.n1310 10.6151
R2445 B.n1310 B.n74 10.6151
R2446 B.n1304 B.n74 10.6151
R2447 B.n1304 B.n1303 10.6151
R2448 B.n1303 B.n1302 10.6151
R2449 B.n1302 B.n81 10.6151
R2450 B.n1296 B.n81 10.6151
R2451 B.n1296 B.n1295 10.6151
R2452 B.n1295 B.n1294 10.6151
R2453 B.n1294 B.n88 10.6151
R2454 B.n1288 B.n88 10.6151
R2455 B.n1288 B.n1287 10.6151
R2456 B.n1287 B.n1286 10.6151
R2457 B.n1286 B.n95 10.6151
R2458 B.n1280 B.n95 10.6151
R2459 B.n1280 B.n1279 10.6151
R2460 B.n1279 B.n1278 10.6151
R2461 B.n1278 B.n102 10.6151
R2462 B.n1272 B.n102 10.6151
R2463 B.n1272 B.n1271 10.6151
R2464 B.n1271 B.n1270 10.6151
R2465 B.n1270 B.n109 10.6151
R2466 B.n1264 B.n109 10.6151
R2467 B.n1264 B.n1263 10.6151
R2468 B.n1263 B.n1262 10.6151
R2469 B.n1262 B.n116 10.6151
R2470 B.n1256 B.n116 10.6151
R2471 B.n1256 B.n1255 10.6151
R2472 B.n1255 B.n1254 10.6151
R2473 B.n1254 B.n122 10.6151
R2474 B.n1248 B.n122 10.6151
R2475 B.n1248 B.n1247 10.6151
R2476 B.n1247 B.n1246 10.6151
R2477 B.n1246 B.n130 10.6151
R2478 B.n1240 B.n130 10.6151
R2479 B.n1240 B.n1239 10.6151
R2480 B.n1239 B.n1238 10.6151
R2481 B.n207 B.n137 10.6151
R2482 B.n210 B.n207 10.6151
R2483 B.n211 B.n210 10.6151
R2484 B.n214 B.n211 10.6151
R2485 B.n215 B.n214 10.6151
R2486 B.n218 B.n215 10.6151
R2487 B.n219 B.n218 10.6151
R2488 B.n222 B.n219 10.6151
R2489 B.n223 B.n222 10.6151
R2490 B.n226 B.n223 10.6151
R2491 B.n227 B.n226 10.6151
R2492 B.n230 B.n227 10.6151
R2493 B.n231 B.n230 10.6151
R2494 B.n234 B.n231 10.6151
R2495 B.n235 B.n234 10.6151
R2496 B.n238 B.n235 10.6151
R2497 B.n239 B.n238 10.6151
R2498 B.n242 B.n239 10.6151
R2499 B.n243 B.n242 10.6151
R2500 B.n246 B.n243 10.6151
R2501 B.n247 B.n246 10.6151
R2502 B.n250 B.n247 10.6151
R2503 B.n251 B.n250 10.6151
R2504 B.n254 B.n251 10.6151
R2505 B.n255 B.n254 10.6151
R2506 B.n258 B.n255 10.6151
R2507 B.n259 B.n258 10.6151
R2508 B.n262 B.n259 10.6151
R2509 B.n263 B.n262 10.6151
R2510 B.n266 B.n263 10.6151
R2511 B.n267 B.n266 10.6151
R2512 B.n270 B.n267 10.6151
R2513 B.n271 B.n270 10.6151
R2514 B.n274 B.n271 10.6151
R2515 B.n275 B.n274 10.6151
R2516 B.n278 B.n275 10.6151
R2517 B.n279 B.n278 10.6151
R2518 B.n282 B.n279 10.6151
R2519 B.n283 B.n282 10.6151
R2520 B.n286 B.n283 10.6151
R2521 B.n287 B.n286 10.6151
R2522 B.n290 B.n287 10.6151
R2523 B.n291 B.n290 10.6151
R2524 B.n294 B.n291 10.6151
R2525 B.n295 B.n294 10.6151
R2526 B.n298 B.n295 10.6151
R2527 B.n299 B.n298 10.6151
R2528 B.n302 B.n299 10.6151
R2529 B.n303 B.n302 10.6151
R2530 B.n306 B.n303 10.6151
R2531 B.n307 B.n306 10.6151
R2532 B.n310 B.n307 10.6151
R2533 B.n311 B.n310 10.6151
R2534 B.n314 B.n311 10.6151
R2535 B.n315 B.n314 10.6151
R2536 B.n319 B.n318 10.6151
R2537 B.n322 B.n319 10.6151
R2538 B.n323 B.n322 10.6151
R2539 B.n326 B.n323 10.6151
R2540 B.n327 B.n326 10.6151
R2541 B.n330 B.n327 10.6151
R2542 B.n331 B.n330 10.6151
R2543 B.n334 B.n331 10.6151
R2544 B.n335 B.n334 10.6151
R2545 B.n339 B.n338 10.6151
R2546 B.n342 B.n339 10.6151
R2547 B.n343 B.n342 10.6151
R2548 B.n346 B.n343 10.6151
R2549 B.n347 B.n346 10.6151
R2550 B.n350 B.n347 10.6151
R2551 B.n351 B.n350 10.6151
R2552 B.n354 B.n351 10.6151
R2553 B.n355 B.n354 10.6151
R2554 B.n358 B.n355 10.6151
R2555 B.n359 B.n358 10.6151
R2556 B.n362 B.n359 10.6151
R2557 B.n363 B.n362 10.6151
R2558 B.n366 B.n363 10.6151
R2559 B.n367 B.n366 10.6151
R2560 B.n370 B.n367 10.6151
R2561 B.n371 B.n370 10.6151
R2562 B.n374 B.n371 10.6151
R2563 B.n375 B.n374 10.6151
R2564 B.n378 B.n375 10.6151
R2565 B.n379 B.n378 10.6151
R2566 B.n382 B.n379 10.6151
R2567 B.n383 B.n382 10.6151
R2568 B.n386 B.n383 10.6151
R2569 B.n387 B.n386 10.6151
R2570 B.n390 B.n387 10.6151
R2571 B.n391 B.n390 10.6151
R2572 B.n394 B.n391 10.6151
R2573 B.n395 B.n394 10.6151
R2574 B.n398 B.n395 10.6151
R2575 B.n399 B.n398 10.6151
R2576 B.n402 B.n399 10.6151
R2577 B.n403 B.n402 10.6151
R2578 B.n406 B.n403 10.6151
R2579 B.n407 B.n406 10.6151
R2580 B.n410 B.n407 10.6151
R2581 B.n411 B.n410 10.6151
R2582 B.n414 B.n411 10.6151
R2583 B.n415 B.n414 10.6151
R2584 B.n418 B.n415 10.6151
R2585 B.n419 B.n418 10.6151
R2586 B.n422 B.n419 10.6151
R2587 B.n423 B.n422 10.6151
R2588 B.n426 B.n423 10.6151
R2589 B.n427 B.n426 10.6151
R2590 B.n430 B.n427 10.6151
R2591 B.n431 B.n430 10.6151
R2592 B.n434 B.n431 10.6151
R2593 B.n435 B.n434 10.6151
R2594 B.n438 B.n435 10.6151
R2595 B.n439 B.n438 10.6151
R2596 B.n442 B.n439 10.6151
R2597 B.n444 B.n442 10.6151
R2598 B.n445 B.n444 10.6151
R2599 B.n1232 B.n445 10.6151
R2600 B.n768 B.n767 9.36635
R2601 B.n788 B.n622 9.36635
R2602 B.n315 B.n206 9.36635
R2603 B.n338 B.n203 9.36635
R2604 B.n1392 B.n0 8.11757
R2605 B.n1392 B.n1 8.11757
R2606 B.n1110 B.t5 6.90788
R2607 B.n19 B.t0 6.90788
R2608 B.n1080 B.t8 5.92111
R2609 B.n1354 B.t1 5.92111
R2610 B.n928 B.t11 2.9608
R2611 B.n124 B.t15 2.9608
R2612 B.n526 B.t2 1.97404
R2613 B.t6 B.n1307 1.97404
R2614 B.n769 B.n768 1.24928
R2615 B.n789 B.n788 1.24928
R2616 B.n318 B.n206 1.24928
R2617 B.n335 B.n203 1.24928
R2618 VP.n32 VP.n31 161.3
R2619 VP.n33 VP.n28 161.3
R2620 VP.n35 VP.n34 161.3
R2621 VP.n36 VP.n27 161.3
R2622 VP.n38 VP.n37 161.3
R2623 VP.n39 VP.n26 161.3
R2624 VP.n41 VP.n40 161.3
R2625 VP.n42 VP.n25 161.3
R2626 VP.n44 VP.n43 161.3
R2627 VP.n45 VP.n24 161.3
R2628 VP.n47 VP.n46 161.3
R2629 VP.n48 VP.n23 161.3
R2630 VP.n50 VP.n49 161.3
R2631 VP.n51 VP.n22 161.3
R2632 VP.n54 VP.n53 161.3
R2633 VP.n55 VP.n21 161.3
R2634 VP.n57 VP.n56 161.3
R2635 VP.n58 VP.n20 161.3
R2636 VP.n60 VP.n59 161.3
R2637 VP.n61 VP.n19 161.3
R2638 VP.n63 VP.n62 161.3
R2639 VP.n64 VP.n18 161.3
R2640 VP.n66 VP.n65 161.3
R2641 VP.n117 VP.n116 161.3
R2642 VP.n115 VP.n1 161.3
R2643 VP.n114 VP.n113 161.3
R2644 VP.n112 VP.n2 161.3
R2645 VP.n111 VP.n110 161.3
R2646 VP.n109 VP.n3 161.3
R2647 VP.n108 VP.n107 161.3
R2648 VP.n106 VP.n4 161.3
R2649 VP.n105 VP.n104 161.3
R2650 VP.n102 VP.n5 161.3
R2651 VP.n101 VP.n100 161.3
R2652 VP.n99 VP.n6 161.3
R2653 VP.n98 VP.n97 161.3
R2654 VP.n96 VP.n7 161.3
R2655 VP.n95 VP.n94 161.3
R2656 VP.n93 VP.n8 161.3
R2657 VP.n92 VP.n91 161.3
R2658 VP.n90 VP.n9 161.3
R2659 VP.n89 VP.n88 161.3
R2660 VP.n87 VP.n10 161.3
R2661 VP.n86 VP.n85 161.3
R2662 VP.n84 VP.n11 161.3
R2663 VP.n83 VP.n82 161.3
R2664 VP.n81 VP.n80 161.3
R2665 VP.n79 VP.n13 161.3
R2666 VP.n78 VP.n77 161.3
R2667 VP.n76 VP.n14 161.3
R2668 VP.n75 VP.n74 161.3
R2669 VP.n73 VP.n15 161.3
R2670 VP.n72 VP.n71 161.3
R2671 VP.n70 VP.n16 161.3
R2672 VP.n30 VP.t9 149.601
R2673 VP.n8 VP.t1 115.871
R2674 VP.n68 VP.t6 115.871
R2675 VP.n12 VP.t7 115.871
R2676 VP.n103 VP.t0 115.871
R2677 VP.n0 VP.t3 115.871
R2678 VP.n25 VP.t5 115.871
R2679 VP.n17 VP.t4 115.871
R2680 VP.n52 VP.t2 115.871
R2681 VP.n29 VP.t8 115.871
R2682 VP.n69 VP.n68 78.4415
R2683 VP.n118 VP.n0 78.4415
R2684 VP.n67 VP.n17 78.4415
R2685 VP.n69 VP.n67 62.1549
R2686 VP.n30 VP.n29 56.6961
R2687 VP.n74 VP.n14 56.5617
R2688 VP.n110 VP.n2 56.5617
R2689 VP.n59 VP.n19 56.5617
R2690 VP.n89 VP.n10 46.874
R2691 VP.n97 VP.n6 46.874
R2692 VP.n46 VP.n23 46.874
R2693 VP.n38 VP.n27 46.874
R2694 VP.n85 VP.n10 34.28
R2695 VP.n101 VP.n6 34.28
R2696 VP.n50 VP.n23 34.28
R2697 VP.n34 VP.n27 34.28
R2698 VP.n72 VP.n16 24.5923
R2699 VP.n73 VP.n72 24.5923
R2700 VP.n74 VP.n73 24.5923
R2701 VP.n78 VP.n14 24.5923
R2702 VP.n79 VP.n78 24.5923
R2703 VP.n80 VP.n79 24.5923
R2704 VP.n84 VP.n83 24.5923
R2705 VP.n85 VP.n84 24.5923
R2706 VP.n90 VP.n89 24.5923
R2707 VP.n91 VP.n90 24.5923
R2708 VP.n91 VP.n8 24.5923
R2709 VP.n95 VP.n8 24.5923
R2710 VP.n96 VP.n95 24.5923
R2711 VP.n97 VP.n96 24.5923
R2712 VP.n102 VP.n101 24.5923
R2713 VP.n104 VP.n102 24.5923
R2714 VP.n108 VP.n4 24.5923
R2715 VP.n109 VP.n108 24.5923
R2716 VP.n110 VP.n109 24.5923
R2717 VP.n114 VP.n2 24.5923
R2718 VP.n115 VP.n114 24.5923
R2719 VP.n116 VP.n115 24.5923
R2720 VP.n63 VP.n19 24.5923
R2721 VP.n64 VP.n63 24.5923
R2722 VP.n65 VP.n64 24.5923
R2723 VP.n51 VP.n50 24.5923
R2724 VP.n53 VP.n51 24.5923
R2725 VP.n57 VP.n21 24.5923
R2726 VP.n58 VP.n57 24.5923
R2727 VP.n59 VP.n58 24.5923
R2728 VP.n39 VP.n38 24.5923
R2729 VP.n40 VP.n39 24.5923
R2730 VP.n40 VP.n25 24.5923
R2731 VP.n44 VP.n25 24.5923
R2732 VP.n45 VP.n44 24.5923
R2733 VP.n46 VP.n45 24.5923
R2734 VP.n33 VP.n32 24.5923
R2735 VP.n34 VP.n33 24.5923
R2736 VP.n83 VP.n12 18.1985
R2737 VP.n104 VP.n103 18.1985
R2738 VP.n53 VP.n52 18.1985
R2739 VP.n32 VP.n29 18.1985
R2740 VP.n68 VP.n16 11.8046
R2741 VP.n116 VP.n0 11.8046
R2742 VP.n65 VP.n17 11.8046
R2743 VP.n80 VP.n12 6.39438
R2744 VP.n103 VP.n4 6.39438
R2745 VP.n52 VP.n21 6.39438
R2746 VP.n31 VP.n30 3.08735
R2747 VP.n67 VP.n66 0.354861
R2748 VP.n70 VP.n69 0.354861
R2749 VP.n118 VP.n117 0.354861
R2750 VP VP.n118 0.267071
R2751 VP.n31 VP.n28 0.189894
R2752 VP.n35 VP.n28 0.189894
R2753 VP.n36 VP.n35 0.189894
R2754 VP.n37 VP.n36 0.189894
R2755 VP.n37 VP.n26 0.189894
R2756 VP.n41 VP.n26 0.189894
R2757 VP.n42 VP.n41 0.189894
R2758 VP.n43 VP.n42 0.189894
R2759 VP.n43 VP.n24 0.189894
R2760 VP.n47 VP.n24 0.189894
R2761 VP.n48 VP.n47 0.189894
R2762 VP.n49 VP.n48 0.189894
R2763 VP.n49 VP.n22 0.189894
R2764 VP.n54 VP.n22 0.189894
R2765 VP.n55 VP.n54 0.189894
R2766 VP.n56 VP.n55 0.189894
R2767 VP.n56 VP.n20 0.189894
R2768 VP.n60 VP.n20 0.189894
R2769 VP.n61 VP.n60 0.189894
R2770 VP.n62 VP.n61 0.189894
R2771 VP.n62 VP.n18 0.189894
R2772 VP.n66 VP.n18 0.189894
R2773 VP.n71 VP.n70 0.189894
R2774 VP.n71 VP.n15 0.189894
R2775 VP.n75 VP.n15 0.189894
R2776 VP.n76 VP.n75 0.189894
R2777 VP.n77 VP.n76 0.189894
R2778 VP.n77 VP.n13 0.189894
R2779 VP.n81 VP.n13 0.189894
R2780 VP.n82 VP.n81 0.189894
R2781 VP.n82 VP.n11 0.189894
R2782 VP.n86 VP.n11 0.189894
R2783 VP.n87 VP.n86 0.189894
R2784 VP.n88 VP.n87 0.189894
R2785 VP.n88 VP.n9 0.189894
R2786 VP.n92 VP.n9 0.189894
R2787 VP.n93 VP.n92 0.189894
R2788 VP.n94 VP.n93 0.189894
R2789 VP.n94 VP.n7 0.189894
R2790 VP.n98 VP.n7 0.189894
R2791 VP.n99 VP.n98 0.189894
R2792 VP.n100 VP.n99 0.189894
R2793 VP.n100 VP.n5 0.189894
R2794 VP.n105 VP.n5 0.189894
R2795 VP.n106 VP.n105 0.189894
R2796 VP.n107 VP.n106 0.189894
R2797 VP.n107 VP.n3 0.189894
R2798 VP.n111 VP.n3 0.189894
R2799 VP.n112 VP.n111 0.189894
R2800 VP.n113 VP.n112 0.189894
R2801 VP.n113 VP.n1 0.189894
R2802 VP.n117 VP.n1 0.189894
R2803 VDD1.n1 VDD1.t0 68.7824
R2804 VDD1.n3 VDD1.t3 68.7814
R2805 VDD1.n5 VDD1.n4 66.7286
R2806 VDD1.n1 VDD1.n0 64.2828
R2807 VDD1.n7 VDD1.n6 64.2818
R2808 VDD1.n3 VDD1.n2 64.2818
R2809 VDD1.n7 VDD1.n5 56.4858
R2810 VDD1 VDD1.n7 2.44447
R2811 VDD1.n6 VDD1.t7 1.16384
R2812 VDD1.n6 VDD1.t5 1.16384
R2813 VDD1.n0 VDD1.t1 1.16384
R2814 VDD1.n0 VDD1.t4 1.16384
R2815 VDD1.n4 VDD1.t9 1.16384
R2816 VDD1.n4 VDD1.t6 1.16384
R2817 VDD1.n2 VDD1.t2 1.16384
R2818 VDD1.n2 VDD1.t8 1.16384
R2819 VDD1 VDD1.n1 0.892741
R2820 VDD1.n5 VDD1.n3 0.779206
C0 VTAIL VP 16.561802f
C1 VDD1 VP 16.283098f
C2 VDD2 VP 0.704153f
C3 VTAIL VN 16.5475f
C4 VDD1 VN 0.155832f
C5 VDD2 VN 15.7394f
C6 VTAIL VDD1 12.833f
C7 VTAIL VDD2 12.8902f
C8 VDD1 VDD2 2.78711f
C9 VP VN 10.7046f
C10 VDD2 B 9.155993f
C11 VDD1 B 9.156056f
C12 VTAIL B 10.955367f
C13 VN B 22.994202f
C14 VP B 21.533428f
C15 VDD1.t0 B 3.81156f
C16 VDD1.t1 B 0.324829f
C17 VDD1.t4 B 0.324829f
C18 VDD1.n0 B 2.96303f
C19 VDD1.n1 B 1.01423f
C20 VDD1.t3 B 3.81157f
C21 VDD1.t2 B 0.324829f
C22 VDD1.t8 B 0.324829f
C23 VDD1.n2 B 2.96304f
C24 VDD1.n3 B 1.00609f
C25 VDD1.t9 B 0.324829f
C26 VDD1.t6 B 0.324829f
C27 VDD1.n4 B 2.98684f
C28 VDD1.n5 B 3.72476f
C29 VDD1.t7 B 0.324829f
C30 VDD1.t5 B 0.324829f
C31 VDD1.n6 B 2.96302f
C32 VDD1.n7 B 3.79761f
C33 VP.t3 B 2.805f
C34 VP.n0 B 1.0366f
C35 VP.n1 B 0.016944f
C36 VP.n2 B 0.022053f
C37 VP.n3 B 0.016944f
C38 VP.n4 B 0.019942f
C39 VP.n5 B 0.016944f
C40 VP.n6 B 0.01462f
C41 VP.n7 B 0.016944f
C42 VP.t1 B 2.805f
C43 VP.n8 B 0.9851f
C44 VP.n9 B 0.016944f
C45 VP.n10 B 0.01462f
C46 VP.n11 B 0.016944f
C47 VP.t7 B 2.805f
C48 VP.n12 B 0.96919f
C49 VP.n13 B 0.016944f
C50 VP.n14 B 0.027209f
C51 VP.n15 B 0.016944f
C52 VP.n16 B 0.023355f
C53 VP.t4 B 2.805f
C54 VP.n17 B 1.0366f
C55 VP.n18 B 0.016944f
C56 VP.n19 B 0.022053f
C57 VP.n20 B 0.016944f
C58 VP.n21 B 0.019942f
C59 VP.n22 B 0.016944f
C60 VP.n23 B 0.01462f
C61 VP.n24 B 0.016944f
C62 VP.t5 B 2.805f
C63 VP.n25 B 0.9851f
C64 VP.n26 B 0.016944f
C65 VP.n27 B 0.01462f
C66 VP.n28 B 0.016944f
C67 VP.t8 B 2.805f
C68 VP.n29 B 1.03143f
C69 VP.t9 B 3.05235f
C70 VP.n30 B 0.980107f
C71 VP.n31 B 0.209455f
C72 VP.n32 B 0.027388f
C73 VP.n33 B 0.031421f
C74 VP.n34 B 0.034052f
C75 VP.n35 B 0.016944f
C76 VP.n36 B 0.016944f
C77 VP.n37 B 0.016944f
C78 VP.n38 B 0.032011f
C79 VP.n39 B 0.031421f
C80 VP.n40 B 0.031421f
C81 VP.n41 B 0.016944f
C82 VP.n42 B 0.016944f
C83 VP.n43 B 0.016944f
C84 VP.n44 B 0.031421f
C85 VP.n45 B 0.031421f
C86 VP.n46 B 0.032011f
C87 VP.n47 B 0.016944f
C88 VP.n48 B 0.016944f
C89 VP.n49 B 0.016944f
C90 VP.n50 B 0.034052f
C91 VP.n51 B 0.031421f
C92 VP.t2 B 2.805f
C93 VP.n52 B 0.96919f
C94 VP.n53 B 0.027388f
C95 VP.n54 B 0.016944f
C96 VP.n55 B 0.016944f
C97 VP.n56 B 0.016944f
C98 VP.n57 B 0.031421f
C99 VP.n58 B 0.031421f
C100 VP.n59 B 0.027209f
C101 VP.n60 B 0.016944f
C102 VP.n61 B 0.016944f
C103 VP.n62 B 0.016944f
C104 VP.n63 B 0.031421f
C105 VP.n64 B 0.031421f
C106 VP.n65 B 0.023355f
C107 VP.n66 B 0.027343f
C108 VP.n67 B 1.30474f
C109 VP.t6 B 2.805f
C110 VP.n68 B 1.0366f
C111 VP.n69 B 1.31457f
C112 VP.n70 B 0.027343f
C113 VP.n71 B 0.016944f
C114 VP.n72 B 0.031421f
C115 VP.n73 B 0.031421f
C116 VP.n74 B 0.022053f
C117 VP.n75 B 0.016944f
C118 VP.n76 B 0.016944f
C119 VP.n77 B 0.016944f
C120 VP.n78 B 0.031421f
C121 VP.n79 B 0.031421f
C122 VP.n80 B 0.019942f
C123 VP.n81 B 0.016944f
C124 VP.n82 B 0.016944f
C125 VP.n83 B 0.027388f
C126 VP.n84 B 0.031421f
C127 VP.n85 B 0.034052f
C128 VP.n86 B 0.016944f
C129 VP.n87 B 0.016944f
C130 VP.n88 B 0.016944f
C131 VP.n89 B 0.032011f
C132 VP.n90 B 0.031421f
C133 VP.n91 B 0.031421f
C134 VP.n92 B 0.016944f
C135 VP.n93 B 0.016944f
C136 VP.n94 B 0.016944f
C137 VP.n95 B 0.031421f
C138 VP.n96 B 0.031421f
C139 VP.n97 B 0.032011f
C140 VP.n98 B 0.016944f
C141 VP.n99 B 0.016944f
C142 VP.n100 B 0.016944f
C143 VP.n101 B 0.034052f
C144 VP.n102 B 0.031421f
C145 VP.t0 B 2.805f
C146 VP.n103 B 0.96919f
C147 VP.n104 B 0.027388f
C148 VP.n105 B 0.016944f
C149 VP.n106 B 0.016944f
C150 VP.n107 B 0.016944f
C151 VP.n108 B 0.031421f
C152 VP.n109 B 0.031421f
C153 VP.n110 B 0.027209f
C154 VP.n111 B 0.016944f
C155 VP.n112 B 0.016944f
C156 VP.n113 B 0.016944f
C157 VP.n114 B 0.031421f
C158 VP.n115 B 0.031421f
C159 VP.n116 B 0.023355f
C160 VP.n117 B 0.027343f
C161 VP.n118 B 0.044673f
C162 VTAIL.t14 B 0.326881f
C163 VTAIL.t18 B 0.326881f
C164 VTAIL.n0 B 2.91667f
C165 VTAIL.n1 B 0.590402f
C166 VTAIL.t5 B 3.72511f
C167 VTAIL.n2 B 0.73421f
C168 VTAIL.t7 B 0.326881f
C169 VTAIL.t8 B 0.326881f
C170 VTAIL.n3 B 2.91667f
C171 VTAIL.n4 B 0.745002f
C172 VTAIL.t3 B 0.326881f
C173 VTAIL.t2 B 0.326881f
C174 VTAIL.n5 B 2.91667f
C175 VTAIL.n6 B 2.48545f
C176 VTAIL.t17 B 0.326881f
C177 VTAIL.t15 B 0.326881f
C178 VTAIL.n7 B 2.91665f
C179 VTAIL.n8 B 2.48546f
C180 VTAIL.t13 B 0.326881f
C181 VTAIL.t10 B 0.326881f
C182 VTAIL.n9 B 2.91665f
C183 VTAIL.n10 B 0.745016f
C184 VTAIL.t12 B 3.7251f
C185 VTAIL.n11 B 0.734222f
C186 VTAIL.t0 B 0.326881f
C187 VTAIL.t1 B 0.326881f
C188 VTAIL.n12 B 2.91665f
C189 VTAIL.n13 B 0.651176f
C190 VTAIL.t4 B 0.326881f
C191 VTAIL.t6 B 0.326881f
C192 VTAIL.n14 B 2.91665f
C193 VTAIL.n15 B 0.745016f
C194 VTAIL.t19 B 3.7251f
C195 VTAIL.n16 B 2.30724f
C196 VTAIL.t11 B 3.72511f
C197 VTAIL.n17 B 2.30723f
C198 VTAIL.t16 B 0.326881f
C199 VTAIL.t9 B 0.326881f
C200 VTAIL.n18 B 2.91667f
C201 VTAIL.n19 B 0.544494f
C202 VDD2.t8 B 3.76235f
C203 VDD2.t3 B 0.320634f
C204 VDD2.t1 B 0.320634f
C205 VDD2.n0 B 2.92477f
C206 VDD2.n1 B 0.993095f
C207 VDD2.t0 B 0.320634f
C208 VDD2.t5 B 0.320634f
C209 VDD2.n2 B 2.94827f
C210 VDD2.n3 B 3.52941f
C211 VDD2.t2 B 3.73739f
C212 VDD2.n4 B 3.68185f
C213 VDD2.t9 B 0.320634f
C214 VDD2.t7 B 0.320634f
C215 VDD2.n5 B 2.92476f
C216 VDD2.n6 B 0.511593f
C217 VDD2.t4 B 0.320634f
C218 VDD2.t6 B 0.320634f
C219 VDD2.n7 B 2.94822f
C220 VN.t7 B 2.75846f
C221 VN.n0 B 1.0194f
C222 VN.n1 B 0.016663f
C223 VN.n2 B 0.021687f
C224 VN.n3 B 0.016663f
C225 VN.n4 B 0.019612f
C226 VN.n5 B 0.016663f
C227 VN.n6 B 0.014378f
C228 VN.n7 B 0.016663f
C229 VN.t2 B 2.75846f
C230 VN.n8 B 0.968755f
C231 VN.n9 B 0.016663f
C232 VN.n10 B 0.014378f
C233 VN.n11 B 0.016663f
C234 VN.t0 B 2.75846f
C235 VN.n12 B 1.01432f
C236 VN.t4 B 3.0017f
C237 VN.n13 B 0.963844f
C238 VN.n14 B 0.205979f
C239 VN.n15 B 0.026934f
C240 VN.n16 B 0.0309f
C241 VN.n17 B 0.033487f
C242 VN.n18 B 0.016663f
C243 VN.n19 B 0.016663f
C244 VN.n20 B 0.016663f
C245 VN.n21 B 0.03148f
C246 VN.n22 B 0.0309f
C247 VN.n23 B 0.0309f
C248 VN.n24 B 0.016663f
C249 VN.n25 B 0.016663f
C250 VN.n26 B 0.016663f
C251 VN.n27 B 0.0309f
C252 VN.n28 B 0.0309f
C253 VN.n29 B 0.03148f
C254 VN.n30 B 0.016663f
C255 VN.n31 B 0.016663f
C256 VN.n32 B 0.016663f
C257 VN.n33 B 0.033487f
C258 VN.n34 B 0.0309f
C259 VN.t9 B 2.75846f
C260 VN.n35 B 0.953109f
C261 VN.n36 B 0.026934f
C262 VN.n37 B 0.016663f
C263 VN.n38 B 0.016663f
C264 VN.n39 B 0.016663f
C265 VN.n40 B 0.0309f
C266 VN.n41 B 0.0309f
C267 VN.n42 B 0.026758f
C268 VN.n43 B 0.016663f
C269 VN.n44 B 0.016663f
C270 VN.n45 B 0.016663f
C271 VN.n46 B 0.0309f
C272 VN.n47 B 0.0309f
C273 VN.n48 B 0.022968f
C274 VN.n49 B 0.026889f
C275 VN.n50 B 0.043932f
C276 VN.t1 B 2.75846f
C277 VN.n51 B 1.0194f
C278 VN.n52 B 0.016663f
C279 VN.n53 B 0.021687f
C280 VN.n54 B 0.016663f
C281 VN.n55 B 0.019612f
C282 VN.n56 B 0.016663f
C283 VN.t3 B 2.75846f
C284 VN.n57 B 0.953109f
C285 VN.n58 B 0.014378f
C286 VN.n59 B 0.016663f
C287 VN.t5 B 2.75846f
C288 VN.n60 B 0.968755f
C289 VN.n61 B 0.016663f
C290 VN.n62 B 0.014378f
C291 VN.n63 B 0.016663f
C292 VN.t8 B 2.75846f
C293 VN.n64 B 1.01432f
C294 VN.t6 B 3.0017f
C295 VN.n65 B 0.963844f
C296 VN.n66 B 0.205979f
C297 VN.n67 B 0.026934f
C298 VN.n68 B 0.0309f
C299 VN.n69 B 0.033487f
C300 VN.n70 B 0.016663f
C301 VN.n71 B 0.016663f
C302 VN.n72 B 0.016663f
C303 VN.n73 B 0.03148f
C304 VN.n74 B 0.0309f
C305 VN.n75 B 0.0309f
C306 VN.n76 B 0.016663f
C307 VN.n77 B 0.016663f
C308 VN.n78 B 0.016663f
C309 VN.n79 B 0.0309f
C310 VN.n80 B 0.0309f
C311 VN.n81 B 0.03148f
C312 VN.n82 B 0.016663f
C313 VN.n83 B 0.016663f
C314 VN.n84 B 0.016663f
C315 VN.n85 B 0.033487f
C316 VN.n86 B 0.0309f
C317 VN.n87 B 0.026934f
C318 VN.n88 B 0.016663f
C319 VN.n89 B 0.016663f
C320 VN.n90 B 0.016663f
C321 VN.n91 B 0.0309f
C322 VN.n92 B 0.0309f
C323 VN.n93 B 0.026758f
C324 VN.n94 B 0.016663f
C325 VN.n95 B 0.016663f
C326 VN.n96 B 0.016663f
C327 VN.n97 B 0.0309f
C328 VN.n98 B 0.0309f
C329 VN.n99 B 0.022968f
C330 VN.n100 B 0.026889f
C331 VN.n101 B 1.28945f
.ends

