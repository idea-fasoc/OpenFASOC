* NGSPICE file created from diff_pair_sample_1385.ext - technology: sky130A

.subckt diff_pair_sample_1385 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 w_n2470_n1796# sky130_fd_pr__pfet_01v8 ad=1.6146 pd=9.06 as=1.6146 ps=9.06 w=4.14 l=3.42
X1 VDD1.t1 VP.t0 VTAIL.t1 w_n2470_n1796# sky130_fd_pr__pfet_01v8 ad=1.6146 pd=9.06 as=1.6146 ps=9.06 w=4.14 l=3.42
X2 B.t11 B.t9 B.t10 w_n2470_n1796# sky130_fd_pr__pfet_01v8 ad=1.6146 pd=9.06 as=0 ps=0 w=4.14 l=3.42
X3 VDD2.t0 VN.t1 VTAIL.t3 w_n2470_n1796# sky130_fd_pr__pfet_01v8 ad=1.6146 pd=9.06 as=1.6146 ps=9.06 w=4.14 l=3.42
X4 B.t8 B.t6 B.t7 w_n2470_n1796# sky130_fd_pr__pfet_01v8 ad=1.6146 pd=9.06 as=0 ps=0 w=4.14 l=3.42
X5 VDD1.t0 VP.t1 VTAIL.t0 w_n2470_n1796# sky130_fd_pr__pfet_01v8 ad=1.6146 pd=9.06 as=1.6146 ps=9.06 w=4.14 l=3.42
X6 B.t5 B.t3 B.t4 w_n2470_n1796# sky130_fd_pr__pfet_01v8 ad=1.6146 pd=9.06 as=0 ps=0 w=4.14 l=3.42
X7 B.t2 B.t0 B.t1 w_n2470_n1796# sky130_fd_pr__pfet_01v8 ad=1.6146 pd=9.06 as=0 ps=0 w=4.14 l=3.42
R0 VN VN.t0 108.803
R1 VN VN.t1 68.5457
R2 VTAIL.n1 VTAIL.t2 98.3957
R3 VTAIL.n3 VTAIL.t3 98.3954
R4 VTAIL.n0 VTAIL.t0 98.3954
R5 VTAIL.n2 VTAIL.t1 98.3954
R6 VTAIL.n1 VTAIL.n0 22.4014
R7 VTAIL.n3 VTAIL.n2 19.1686
R8 VTAIL.n2 VTAIL.n1 2.08671
R9 VTAIL VTAIL.n0 1.33671
R10 VTAIL VTAIL.n3 0.7505
R11 VDD2.n0 VDD2.t0 148.768
R12 VDD2.n0 VDD2.t1 115.075
R13 VDD2 VDD2.n0 0.866879
R14 VP.n0 VP.t0 108.897
R15 VP.n0 VP.t1 68.0198
R16 VP VP.n0 0.526373
R17 VDD1 VDD1.t0 150.101
R18 VDD1 VDD1.t1 115.941
R19 B.n326 B.n45 585
R20 B.n328 B.n327 585
R21 B.n329 B.n44 585
R22 B.n331 B.n330 585
R23 B.n332 B.n43 585
R24 B.n334 B.n333 585
R25 B.n335 B.n42 585
R26 B.n337 B.n336 585
R27 B.n338 B.n41 585
R28 B.n340 B.n339 585
R29 B.n341 B.n40 585
R30 B.n343 B.n342 585
R31 B.n344 B.n39 585
R32 B.n346 B.n345 585
R33 B.n347 B.n38 585
R34 B.n349 B.n348 585
R35 B.n350 B.n37 585
R36 B.n352 B.n351 585
R37 B.n353 B.n34 585
R38 B.n356 B.n355 585
R39 B.n357 B.n33 585
R40 B.n359 B.n358 585
R41 B.n360 B.n32 585
R42 B.n362 B.n361 585
R43 B.n363 B.n31 585
R44 B.n365 B.n364 585
R45 B.n366 B.n27 585
R46 B.n368 B.n367 585
R47 B.n369 B.n26 585
R48 B.n371 B.n370 585
R49 B.n372 B.n25 585
R50 B.n374 B.n373 585
R51 B.n375 B.n24 585
R52 B.n377 B.n376 585
R53 B.n378 B.n23 585
R54 B.n380 B.n379 585
R55 B.n381 B.n22 585
R56 B.n383 B.n382 585
R57 B.n384 B.n21 585
R58 B.n386 B.n385 585
R59 B.n387 B.n20 585
R60 B.n389 B.n388 585
R61 B.n390 B.n19 585
R62 B.n392 B.n391 585
R63 B.n393 B.n18 585
R64 B.n395 B.n394 585
R65 B.n396 B.n17 585
R66 B.n325 B.n324 585
R67 B.n323 B.n46 585
R68 B.n322 B.n321 585
R69 B.n320 B.n47 585
R70 B.n319 B.n318 585
R71 B.n317 B.n48 585
R72 B.n316 B.n315 585
R73 B.n314 B.n49 585
R74 B.n313 B.n312 585
R75 B.n311 B.n50 585
R76 B.n310 B.n309 585
R77 B.n308 B.n51 585
R78 B.n307 B.n306 585
R79 B.n305 B.n52 585
R80 B.n304 B.n303 585
R81 B.n302 B.n53 585
R82 B.n301 B.n300 585
R83 B.n299 B.n54 585
R84 B.n298 B.n297 585
R85 B.n296 B.n55 585
R86 B.n295 B.n294 585
R87 B.n293 B.n56 585
R88 B.n292 B.n291 585
R89 B.n290 B.n57 585
R90 B.n289 B.n288 585
R91 B.n287 B.n58 585
R92 B.n286 B.n285 585
R93 B.n284 B.n59 585
R94 B.n283 B.n282 585
R95 B.n281 B.n60 585
R96 B.n280 B.n279 585
R97 B.n278 B.n61 585
R98 B.n277 B.n276 585
R99 B.n275 B.n62 585
R100 B.n274 B.n273 585
R101 B.n272 B.n63 585
R102 B.n271 B.n270 585
R103 B.n269 B.n64 585
R104 B.n268 B.n267 585
R105 B.n266 B.n65 585
R106 B.n265 B.n264 585
R107 B.n263 B.n66 585
R108 B.n262 B.n261 585
R109 B.n260 B.n67 585
R110 B.n259 B.n258 585
R111 B.n257 B.n68 585
R112 B.n256 B.n255 585
R113 B.n254 B.n69 585
R114 B.n253 B.n252 585
R115 B.n251 B.n70 585
R116 B.n250 B.n249 585
R117 B.n248 B.n71 585
R118 B.n247 B.n246 585
R119 B.n245 B.n72 585
R120 B.n244 B.n243 585
R121 B.n242 B.n73 585
R122 B.n241 B.n240 585
R123 B.n239 B.n74 585
R124 B.n238 B.n237 585
R125 B.n236 B.n75 585
R126 B.n235 B.n234 585
R127 B.n160 B.n101 585
R128 B.n162 B.n161 585
R129 B.n163 B.n100 585
R130 B.n165 B.n164 585
R131 B.n166 B.n99 585
R132 B.n168 B.n167 585
R133 B.n169 B.n98 585
R134 B.n171 B.n170 585
R135 B.n172 B.n97 585
R136 B.n174 B.n173 585
R137 B.n175 B.n96 585
R138 B.n177 B.n176 585
R139 B.n178 B.n95 585
R140 B.n180 B.n179 585
R141 B.n181 B.n94 585
R142 B.n183 B.n182 585
R143 B.n184 B.n93 585
R144 B.n186 B.n185 585
R145 B.n187 B.n90 585
R146 B.n190 B.n189 585
R147 B.n191 B.n89 585
R148 B.n193 B.n192 585
R149 B.n194 B.n88 585
R150 B.n196 B.n195 585
R151 B.n197 B.n87 585
R152 B.n199 B.n198 585
R153 B.n200 B.n86 585
R154 B.n205 B.n204 585
R155 B.n206 B.n85 585
R156 B.n208 B.n207 585
R157 B.n209 B.n84 585
R158 B.n211 B.n210 585
R159 B.n212 B.n83 585
R160 B.n214 B.n213 585
R161 B.n215 B.n82 585
R162 B.n217 B.n216 585
R163 B.n218 B.n81 585
R164 B.n220 B.n219 585
R165 B.n221 B.n80 585
R166 B.n223 B.n222 585
R167 B.n224 B.n79 585
R168 B.n226 B.n225 585
R169 B.n227 B.n78 585
R170 B.n229 B.n228 585
R171 B.n230 B.n77 585
R172 B.n232 B.n231 585
R173 B.n233 B.n76 585
R174 B.n159 B.n158 585
R175 B.n157 B.n102 585
R176 B.n156 B.n155 585
R177 B.n154 B.n103 585
R178 B.n153 B.n152 585
R179 B.n151 B.n104 585
R180 B.n150 B.n149 585
R181 B.n148 B.n105 585
R182 B.n147 B.n146 585
R183 B.n145 B.n106 585
R184 B.n144 B.n143 585
R185 B.n142 B.n107 585
R186 B.n141 B.n140 585
R187 B.n139 B.n108 585
R188 B.n138 B.n137 585
R189 B.n136 B.n109 585
R190 B.n135 B.n134 585
R191 B.n133 B.n110 585
R192 B.n132 B.n131 585
R193 B.n130 B.n111 585
R194 B.n129 B.n128 585
R195 B.n127 B.n112 585
R196 B.n126 B.n125 585
R197 B.n124 B.n113 585
R198 B.n123 B.n122 585
R199 B.n121 B.n114 585
R200 B.n120 B.n119 585
R201 B.n118 B.n115 585
R202 B.n117 B.n116 585
R203 B.n2 B.n0 585
R204 B.n441 B.n1 585
R205 B.n440 B.n439 585
R206 B.n438 B.n3 585
R207 B.n437 B.n436 585
R208 B.n435 B.n4 585
R209 B.n434 B.n433 585
R210 B.n432 B.n5 585
R211 B.n431 B.n430 585
R212 B.n429 B.n6 585
R213 B.n428 B.n427 585
R214 B.n426 B.n7 585
R215 B.n425 B.n424 585
R216 B.n423 B.n8 585
R217 B.n422 B.n421 585
R218 B.n420 B.n9 585
R219 B.n419 B.n418 585
R220 B.n417 B.n10 585
R221 B.n416 B.n415 585
R222 B.n414 B.n11 585
R223 B.n413 B.n412 585
R224 B.n411 B.n12 585
R225 B.n410 B.n409 585
R226 B.n408 B.n13 585
R227 B.n407 B.n406 585
R228 B.n405 B.n14 585
R229 B.n404 B.n403 585
R230 B.n402 B.n15 585
R231 B.n401 B.n400 585
R232 B.n399 B.n16 585
R233 B.n398 B.n397 585
R234 B.n443 B.n442 585
R235 B.n160 B.n159 492.5
R236 B.n398 B.n17 492.5
R237 B.n235 B.n76 492.5
R238 B.n326 B.n325 492.5
R239 B.n201 B.t0 238.195
R240 B.n91 B.t3 238.195
R241 B.n28 B.t9 238.195
R242 B.n35 B.t6 238.195
R243 B.n201 B.t2 192.867
R244 B.n35 B.t7 192.867
R245 B.n91 B.t5 192.863
R246 B.n28 B.t10 192.863
R247 B.n159 B.n102 163.367
R248 B.n155 B.n102 163.367
R249 B.n155 B.n154 163.367
R250 B.n154 B.n153 163.367
R251 B.n153 B.n104 163.367
R252 B.n149 B.n104 163.367
R253 B.n149 B.n148 163.367
R254 B.n148 B.n147 163.367
R255 B.n147 B.n106 163.367
R256 B.n143 B.n106 163.367
R257 B.n143 B.n142 163.367
R258 B.n142 B.n141 163.367
R259 B.n141 B.n108 163.367
R260 B.n137 B.n108 163.367
R261 B.n137 B.n136 163.367
R262 B.n136 B.n135 163.367
R263 B.n135 B.n110 163.367
R264 B.n131 B.n110 163.367
R265 B.n131 B.n130 163.367
R266 B.n130 B.n129 163.367
R267 B.n129 B.n112 163.367
R268 B.n125 B.n112 163.367
R269 B.n125 B.n124 163.367
R270 B.n124 B.n123 163.367
R271 B.n123 B.n114 163.367
R272 B.n119 B.n114 163.367
R273 B.n119 B.n118 163.367
R274 B.n118 B.n117 163.367
R275 B.n117 B.n2 163.367
R276 B.n442 B.n2 163.367
R277 B.n442 B.n441 163.367
R278 B.n441 B.n440 163.367
R279 B.n440 B.n3 163.367
R280 B.n436 B.n3 163.367
R281 B.n436 B.n435 163.367
R282 B.n435 B.n434 163.367
R283 B.n434 B.n5 163.367
R284 B.n430 B.n5 163.367
R285 B.n430 B.n429 163.367
R286 B.n429 B.n428 163.367
R287 B.n428 B.n7 163.367
R288 B.n424 B.n7 163.367
R289 B.n424 B.n423 163.367
R290 B.n423 B.n422 163.367
R291 B.n422 B.n9 163.367
R292 B.n418 B.n9 163.367
R293 B.n418 B.n417 163.367
R294 B.n417 B.n416 163.367
R295 B.n416 B.n11 163.367
R296 B.n412 B.n11 163.367
R297 B.n412 B.n411 163.367
R298 B.n411 B.n410 163.367
R299 B.n410 B.n13 163.367
R300 B.n406 B.n13 163.367
R301 B.n406 B.n405 163.367
R302 B.n405 B.n404 163.367
R303 B.n404 B.n15 163.367
R304 B.n400 B.n15 163.367
R305 B.n400 B.n399 163.367
R306 B.n399 B.n398 163.367
R307 B.n161 B.n160 163.367
R308 B.n161 B.n100 163.367
R309 B.n165 B.n100 163.367
R310 B.n166 B.n165 163.367
R311 B.n167 B.n166 163.367
R312 B.n167 B.n98 163.367
R313 B.n171 B.n98 163.367
R314 B.n172 B.n171 163.367
R315 B.n173 B.n172 163.367
R316 B.n173 B.n96 163.367
R317 B.n177 B.n96 163.367
R318 B.n178 B.n177 163.367
R319 B.n179 B.n178 163.367
R320 B.n179 B.n94 163.367
R321 B.n183 B.n94 163.367
R322 B.n184 B.n183 163.367
R323 B.n185 B.n184 163.367
R324 B.n185 B.n90 163.367
R325 B.n190 B.n90 163.367
R326 B.n191 B.n190 163.367
R327 B.n192 B.n191 163.367
R328 B.n192 B.n88 163.367
R329 B.n196 B.n88 163.367
R330 B.n197 B.n196 163.367
R331 B.n198 B.n197 163.367
R332 B.n198 B.n86 163.367
R333 B.n205 B.n86 163.367
R334 B.n206 B.n205 163.367
R335 B.n207 B.n206 163.367
R336 B.n207 B.n84 163.367
R337 B.n211 B.n84 163.367
R338 B.n212 B.n211 163.367
R339 B.n213 B.n212 163.367
R340 B.n213 B.n82 163.367
R341 B.n217 B.n82 163.367
R342 B.n218 B.n217 163.367
R343 B.n219 B.n218 163.367
R344 B.n219 B.n80 163.367
R345 B.n223 B.n80 163.367
R346 B.n224 B.n223 163.367
R347 B.n225 B.n224 163.367
R348 B.n225 B.n78 163.367
R349 B.n229 B.n78 163.367
R350 B.n230 B.n229 163.367
R351 B.n231 B.n230 163.367
R352 B.n231 B.n76 163.367
R353 B.n236 B.n235 163.367
R354 B.n237 B.n236 163.367
R355 B.n237 B.n74 163.367
R356 B.n241 B.n74 163.367
R357 B.n242 B.n241 163.367
R358 B.n243 B.n242 163.367
R359 B.n243 B.n72 163.367
R360 B.n247 B.n72 163.367
R361 B.n248 B.n247 163.367
R362 B.n249 B.n248 163.367
R363 B.n249 B.n70 163.367
R364 B.n253 B.n70 163.367
R365 B.n254 B.n253 163.367
R366 B.n255 B.n254 163.367
R367 B.n255 B.n68 163.367
R368 B.n259 B.n68 163.367
R369 B.n260 B.n259 163.367
R370 B.n261 B.n260 163.367
R371 B.n261 B.n66 163.367
R372 B.n265 B.n66 163.367
R373 B.n266 B.n265 163.367
R374 B.n267 B.n266 163.367
R375 B.n267 B.n64 163.367
R376 B.n271 B.n64 163.367
R377 B.n272 B.n271 163.367
R378 B.n273 B.n272 163.367
R379 B.n273 B.n62 163.367
R380 B.n277 B.n62 163.367
R381 B.n278 B.n277 163.367
R382 B.n279 B.n278 163.367
R383 B.n279 B.n60 163.367
R384 B.n283 B.n60 163.367
R385 B.n284 B.n283 163.367
R386 B.n285 B.n284 163.367
R387 B.n285 B.n58 163.367
R388 B.n289 B.n58 163.367
R389 B.n290 B.n289 163.367
R390 B.n291 B.n290 163.367
R391 B.n291 B.n56 163.367
R392 B.n295 B.n56 163.367
R393 B.n296 B.n295 163.367
R394 B.n297 B.n296 163.367
R395 B.n297 B.n54 163.367
R396 B.n301 B.n54 163.367
R397 B.n302 B.n301 163.367
R398 B.n303 B.n302 163.367
R399 B.n303 B.n52 163.367
R400 B.n307 B.n52 163.367
R401 B.n308 B.n307 163.367
R402 B.n309 B.n308 163.367
R403 B.n309 B.n50 163.367
R404 B.n313 B.n50 163.367
R405 B.n314 B.n313 163.367
R406 B.n315 B.n314 163.367
R407 B.n315 B.n48 163.367
R408 B.n319 B.n48 163.367
R409 B.n320 B.n319 163.367
R410 B.n321 B.n320 163.367
R411 B.n321 B.n46 163.367
R412 B.n325 B.n46 163.367
R413 B.n394 B.n17 163.367
R414 B.n394 B.n393 163.367
R415 B.n393 B.n392 163.367
R416 B.n392 B.n19 163.367
R417 B.n388 B.n19 163.367
R418 B.n388 B.n387 163.367
R419 B.n387 B.n386 163.367
R420 B.n386 B.n21 163.367
R421 B.n382 B.n21 163.367
R422 B.n382 B.n381 163.367
R423 B.n381 B.n380 163.367
R424 B.n380 B.n23 163.367
R425 B.n376 B.n23 163.367
R426 B.n376 B.n375 163.367
R427 B.n375 B.n374 163.367
R428 B.n374 B.n25 163.367
R429 B.n370 B.n25 163.367
R430 B.n370 B.n369 163.367
R431 B.n369 B.n368 163.367
R432 B.n368 B.n27 163.367
R433 B.n364 B.n27 163.367
R434 B.n364 B.n363 163.367
R435 B.n363 B.n362 163.367
R436 B.n362 B.n32 163.367
R437 B.n358 B.n32 163.367
R438 B.n358 B.n357 163.367
R439 B.n357 B.n356 163.367
R440 B.n356 B.n34 163.367
R441 B.n351 B.n34 163.367
R442 B.n351 B.n350 163.367
R443 B.n350 B.n349 163.367
R444 B.n349 B.n38 163.367
R445 B.n345 B.n38 163.367
R446 B.n345 B.n344 163.367
R447 B.n344 B.n343 163.367
R448 B.n343 B.n40 163.367
R449 B.n339 B.n40 163.367
R450 B.n339 B.n338 163.367
R451 B.n338 B.n337 163.367
R452 B.n337 B.n42 163.367
R453 B.n333 B.n42 163.367
R454 B.n333 B.n332 163.367
R455 B.n332 B.n331 163.367
R456 B.n331 B.n44 163.367
R457 B.n327 B.n44 163.367
R458 B.n327 B.n326 163.367
R459 B.n202 B.t1 120.139
R460 B.n36 B.t8 120.139
R461 B.n92 B.t4 120.135
R462 B.n29 B.t11 120.135
R463 B.n202 B.n201 72.7278
R464 B.n92 B.n91 72.7278
R465 B.n29 B.n28 72.7278
R466 B.n36 B.n35 72.7278
R467 B.n203 B.n202 59.5399
R468 B.n188 B.n92 59.5399
R469 B.n30 B.n29 59.5399
R470 B.n354 B.n36 59.5399
R471 B.n397 B.n396 32.0005
R472 B.n324 B.n45 32.0005
R473 B.n234 B.n233 32.0005
R474 B.n158 B.n101 32.0005
R475 B B.n443 18.0485
R476 B.n396 B.n395 10.6151
R477 B.n395 B.n18 10.6151
R478 B.n391 B.n18 10.6151
R479 B.n391 B.n390 10.6151
R480 B.n390 B.n389 10.6151
R481 B.n389 B.n20 10.6151
R482 B.n385 B.n20 10.6151
R483 B.n385 B.n384 10.6151
R484 B.n384 B.n383 10.6151
R485 B.n383 B.n22 10.6151
R486 B.n379 B.n22 10.6151
R487 B.n379 B.n378 10.6151
R488 B.n378 B.n377 10.6151
R489 B.n377 B.n24 10.6151
R490 B.n373 B.n24 10.6151
R491 B.n373 B.n372 10.6151
R492 B.n372 B.n371 10.6151
R493 B.n371 B.n26 10.6151
R494 B.n367 B.n366 10.6151
R495 B.n366 B.n365 10.6151
R496 B.n365 B.n31 10.6151
R497 B.n361 B.n31 10.6151
R498 B.n361 B.n360 10.6151
R499 B.n360 B.n359 10.6151
R500 B.n359 B.n33 10.6151
R501 B.n355 B.n33 10.6151
R502 B.n353 B.n352 10.6151
R503 B.n352 B.n37 10.6151
R504 B.n348 B.n37 10.6151
R505 B.n348 B.n347 10.6151
R506 B.n347 B.n346 10.6151
R507 B.n346 B.n39 10.6151
R508 B.n342 B.n39 10.6151
R509 B.n342 B.n341 10.6151
R510 B.n341 B.n340 10.6151
R511 B.n340 B.n41 10.6151
R512 B.n336 B.n41 10.6151
R513 B.n336 B.n335 10.6151
R514 B.n335 B.n334 10.6151
R515 B.n334 B.n43 10.6151
R516 B.n330 B.n43 10.6151
R517 B.n330 B.n329 10.6151
R518 B.n329 B.n328 10.6151
R519 B.n328 B.n45 10.6151
R520 B.n234 B.n75 10.6151
R521 B.n238 B.n75 10.6151
R522 B.n239 B.n238 10.6151
R523 B.n240 B.n239 10.6151
R524 B.n240 B.n73 10.6151
R525 B.n244 B.n73 10.6151
R526 B.n245 B.n244 10.6151
R527 B.n246 B.n245 10.6151
R528 B.n246 B.n71 10.6151
R529 B.n250 B.n71 10.6151
R530 B.n251 B.n250 10.6151
R531 B.n252 B.n251 10.6151
R532 B.n252 B.n69 10.6151
R533 B.n256 B.n69 10.6151
R534 B.n257 B.n256 10.6151
R535 B.n258 B.n257 10.6151
R536 B.n258 B.n67 10.6151
R537 B.n262 B.n67 10.6151
R538 B.n263 B.n262 10.6151
R539 B.n264 B.n263 10.6151
R540 B.n264 B.n65 10.6151
R541 B.n268 B.n65 10.6151
R542 B.n269 B.n268 10.6151
R543 B.n270 B.n269 10.6151
R544 B.n270 B.n63 10.6151
R545 B.n274 B.n63 10.6151
R546 B.n275 B.n274 10.6151
R547 B.n276 B.n275 10.6151
R548 B.n276 B.n61 10.6151
R549 B.n280 B.n61 10.6151
R550 B.n281 B.n280 10.6151
R551 B.n282 B.n281 10.6151
R552 B.n282 B.n59 10.6151
R553 B.n286 B.n59 10.6151
R554 B.n287 B.n286 10.6151
R555 B.n288 B.n287 10.6151
R556 B.n288 B.n57 10.6151
R557 B.n292 B.n57 10.6151
R558 B.n293 B.n292 10.6151
R559 B.n294 B.n293 10.6151
R560 B.n294 B.n55 10.6151
R561 B.n298 B.n55 10.6151
R562 B.n299 B.n298 10.6151
R563 B.n300 B.n299 10.6151
R564 B.n300 B.n53 10.6151
R565 B.n304 B.n53 10.6151
R566 B.n305 B.n304 10.6151
R567 B.n306 B.n305 10.6151
R568 B.n306 B.n51 10.6151
R569 B.n310 B.n51 10.6151
R570 B.n311 B.n310 10.6151
R571 B.n312 B.n311 10.6151
R572 B.n312 B.n49 10.6151
R573 B.n316 B.n49 10.6151
R574 B.n317 B.n316 10.6151
R575 B.n318 B.n317 10.6151
R576 B.n318 B.n47 10.6151
R577 B.n322 B.n47 10.6151
R578 B.n323 B.n322 10.6151
R579 B.n324 B.n323 10.6151
R580 B.n162 B.n101 10.6151
R581 B.n163 B.n162 10.6151
R582 B.n164 B.n163 10.6151
R583 B.n164 B.n99 10.6151
R584 B.n168 B.n99 10.6151
R585 B.n169 B.n168 10.6151
R586 B.n170 B.n169 10.6151
R587 B.n170 B.n97 10.6151
R588 B.n174 B.n97 10.6151
R589 B.n175 B.n174 10.6151
R590 B.n176 B.n175 10.6151
R591 B.n176 B.n95 10.6151
R592 B.n180 B.n95 10.6151
R593 B.n181 B.n180 10.6151
R594 B.n182 B.n181 10.6151
R595 B.n182 B.n93 10.6151
R596 B.n186 B.n93 10.6151
R597 B.n187 B.n186 10.6151
R598 B.n189 B.n89 10.6151
R599 B.n193 B.n89 10.6151
R600 B.n194 B.n193 10.6151
R601 B.n195 B.n194 10.6151
R602 B.n195 B.n87 10.6151
R603 B.n199 B.n87 10.6151
R604 B.n200 B.n199 10.6151
R605 B.n204 B.n200 10.6151
R606 B.n208 B.n85 10.6151
R607 B.n209 B.n208 10.6151
R608 B.n210 B.n209 10.6151
R609 B.n210 B.n83 10.6151
R610 B.n214 B.n83 10.6151
R611 B.n215 B.n214 10.6151
R612 B.n216 B.n215 10.6151
R613 B.n216 B.n81 10.6151
R614 B.n220 B.n81 10.6151
R615 B.n221 B.n220 10.6151
R616 B.n222 B.n221 10.6151
R617 B.n222 B.n79 10.6151
R618 B.n226 B.n79 10.6151
R619 B.n227 B.n226 10.6151
R620 B.n228 B.n227 10.6151
R621 B.n228 B.n77 10.6151
R622 B.n232 B.n77 10.6151
R623 B.n233 B.n232 10.6151
R624 B.n158 B.n157 10.6151
R625 B.n157 B.n156 10.6151
R626 B.n156 B.n103 10.6151
R627 B.n152 B.n103 10.6151
R628 B.n152 B.n151 10.6151
R629 B.n151 B.n150 10.6151
R630 B.n150 B.n105 10.6151
R631 B.n146 B.n105 10.6151
R632 B.n146 B.n145 10.6151
R633 B.n145 B.n144 10.6151
R634 B.n144 B.n107 10.6151
R635 B.n140 B.n107 10.6151
R636 B.n140 B.n139 10.6151
R637 B.n139 B.n138 10.6151
R638 B.n138 B.n109 10.6151
R639 B.n134 B.n109 10.6151
R640 B.n134 B.n133 10.6151
R641 B.n133 B.n132 10.6151
R642 B.n132 B.n111 10.6151
R643 B.n128 B.n111 10.6151
R644 B.n128 B.n127 10.6151
R645 B.n127 B.n126 10.6151
R646 B.n126 B.n113 10.6151
R647 B.n122 B.n113 10.6151
R648 B.n122 B.n121 10.6151
R649 B.n121 B.n120 10.6151
R650 B.n120 B.n115 10.6151
R651 B.n116 B.n115 10.6151
R652 B.n116 B.n0 10.6151
R653 B.n439 B.n1 10.6151
R654 B.n439 B.n438 10.6151
R655 B.n438 B.n437 10.6151
R656 B.n437 B.n4 10.6151
R657 B.n433 B.n4 10.6151
R658 B.n433 B.n432 10.6151
R659 B.n432 B.n431 10.6151
R660 B.n431 B.n6 10.6151
R661 B.n427 B.n6 10.6151
R662 B.n427 B.n426 10.6151
R663 B.n426 B.n425 10.6151
R664 B.n425 B.n8 10.6151
R665 B.n421 B.n8 10.6151
R666 B.n421 B.n420 10.6151
R667 B.n420 B.n419 10.6151
R668 B.n419 B.n10 10.6151
R669 B.n415 B.n10 10.6151
R670 B.n415 B.n414 10.6151
R671 B.n414 B.n413 10.6151
R672 B.n413 B.n12 10.6151
R673 B.n409 B.n12 10.6151
R674 B.n409 B.n408 10.6151
R675 B.n408 B.n407 10.6151
R676 B.n407 B.n14 10.6151
R677 B.n403 B.n14 10.6151
R678 B.n403 B.n402 10.6151
R679 B.n402 B.n401 10.6151
R680 B.n401 B.n16 10.6151
R681 B.n397 B.n16 10.6151
R682 B.n367 B.n30 6.5566
R683 B.n355 B.n354 6.5566
R684 B.n189 B.n188 6.5566
R685 B.n204 B.n203 6.5566
R686 B.n30 B.n26 4.05904
R687 B.n354 B.n353 4.05904
R688 B.n188 B.n187 4.05904
R689 B.n203 B.n85 4.05904
R690 B.n443 B.n0 2.81026
R691 B.n443 B.n1 2.81026
C0 VN VTAIL 1.38625f
C1 B VN 1.09261f
C2 VDD1 VDD2 0.774023f
C3 VDD2 VTAIL 3.29292f
C4 B VDD2 1.22035f
C5 VN VDD2 1.16581f
C6 VDD1 VP 1.38317f
C7 VP VTAIL 1.4004f
C8 VP B 1.6159f
C9 VP VN 4.38698f
C10 VP VDD2 0.371904f
C11 VDD1 w_n2470_n1796# 1.33335f
C12 w_n2470_n1796# VTAIL 1.67762f
C13 B w_n2470_n1796# 7.51179f
C14 w_n2470_n1796# VN 3.33417f
C15 w_n2470_n1796# VDD2 1.36906f
C16 VDD1 VTAIL 3.23472f
C17 VDD1 B 1.18278f
C18 B VTAIL 2.07333f
C19 VDD1 VN 0.152997f
C20 VP w_n2470_n1796# 3.64986f
C21 VDD2 VSUBS 0.67124f
C22 VDD1 VSUBS 2.992059f
C23 VTAIL VSUBS 0.503256f
C24 VN VSUBS 5.72858f
C25 VP VSUBS 1.489932f
C26 B VSUBS 3.6478f
C27 w_n2470_n1796# VSUBS 55.812103f
C28 B.n0 VSUBS 0.005561f
C29 B.n1 VSUBS 0.005561f
C30 B.n2 VSUBS 0.008795f
C31 B.n3 VSUBS 0.008795f
C32 B.n4 VSUBS 0.008795f
C33 B.n5 VSUBS 0.008795f
C34 B.n6 VSUBS 0.008795f
C35 B.n7 VSUBS 0.008795f
C36 B.n8 VSUBS 0.008795f
C37 B.n9 VSUBS 0.008795f
C38 B.n10 VSUBS 0.008795f
C39 B.n11 VSUBS 0.008795f
C40 B.n12 VSUBS 0.008795f
C41 B.n13 VSUBS 0.008795f
C42 B.n14 VSUBS 0.008795f
C43 B.n15 VSUBS 0.008795f
C44 B.n16 VSUBS 0.008795f
C45 B.n17 VSUBS 0.021147f
C46 B.n18 VSUBS 0.008795f
C47 B.n19 VSUBS 0.008795f
C48 B.n20 VSUBS 0.008795f
C49 B.n21 VSUBS 0.008795f
C50 B.n22 VSUBS 0.008795f
C51 B.n23 VSUBS 0.008795f
C52 B.n24 VSUBS 0.008795f
C53 B.n25 VSUBS 0.008795f
C54 B.n26 VSUBS 0.006079f
C55 B.n27 VSUBS 0.008795f
C56 B.t11 VSUBS 0.138183f
C57 B.t10 VSUBS 0.16761f
C58 B.t9 VSUBS 0.862802f
C59 B.n28 VSUBS 0.12501f
C60 B.n29 VSUBS 0.090582f
C61 B.n30 VSUBS 0.020377f
C62 B.n31 VSUBS 0.008795f
C63 B.n32 VSUBS 0.008795f
C64 B.n33 VSUBS 0.008795f
C65 B.n34 VSUBS 0.008795f
C66 B.t8 VSUBS 0.138183f
C67 B.t7 VSUBS 0.16761f
C68 B.t6 VSUBS 0.862802f
C69 B.n35 VSUBS 0.12501f
C70 B.n36 VSUBS 0.090582f
C71 B.n37 VSUBS 0.008795f
C72 B.n38 VSUBS 0.008795f
C73 B.n39 VSUBS 0.008795f
C74 B.n40 VSUBS 0.008795f
C75 B.n41 VSUBS 0.008795f
C76 B.n42 VSUBS 0.008795f
C77 B.n43 VSUBS 0.008795f
C78 B.n44 VSUBS 0.008795f
C79 B.n45 VSUBS 0.020086f
C80 B.n46 VSUBS 0.008795f
C81 B.n47 VSUBS 0.008795f
C82 B.n48 VSUBS 0.008795f
C83 B.n49 VSUBS 0.008795f
C84 B.n50 VSUBS 0.008795f
C85 B.n51 VSUBS 0.008795f
C86 B.n52 VSUBS 0.008795f
C87 B.n53 VSUBS 0.008795f
C88 B.n54 VSUBS 0.008795f
C89 B.n55 VSUBS 0.008795f
C90 B.n56 VSUBS 0.008795f
C91 B.n57 VSUBS 0.008795f
C92 B.n58 VSUBS 0.008795f
C93 B.n59 VSUBS 0.008795f
C94 B.n60 VSUBS 0.008795f
C95 B.n61 VSUBS 0.008795f
C96 B.n62 VSUBS 0.008795f
C97 B.n63 VSUBS 0.008795f
C98 B.n64 VSUBS 0.008795f
C99 B.n65 VSUBS 0.008795f
C100 B.n66 VSUBS 0.008795f
C101 B.n67 VSUBS 0.008795f
C102 B.n68 VSUBS 0.008795f
C103 B.n69 VSUBS 0.008795f
C104 B.n70 VSUBS 0.008795f
C105 B.n71 VSUBS 0.008795f
C106 B.n72 VSUBS 0.008795f
C107 B.n73 VSUBS 0.008795f
C108 B.n74 VSUBS 0.008795f
C109 B.n75 VSUBS 0.008795f
C110 B.n76 VSUBS 0.021147f
C111 B.n77 VSUBS 0.008795f
C112 B.n78 VSUBS 0.008795f
C113 B.n79 VSUBS 0.008795f
C114 B.n80 VSUBS 0.008795f
C115 B.n81 VSUBS 0.008795f
C116 B.n82 VSUBS 0.008795f
C117 B.n83 VSUBS 0.008795f
C118 B.n84 VSUBS 0.008795f
C119 B.n85 VSUBS 0.006079f
C120 B.n86 VSUBS 0.008795f
C121 B.n87 VSUBS 0.008795f
C122 B.n88 VSUBS 0.008795f
C123 B.n89 VSUBS 0.008795f
C124 B.n90 VSUBS 0.008795f
C125 B.t4 VSUBS 0.138183f
C126 B.t5 VSUBS 0.16761f
C127 B.t3 VSUBS 0.862802f
C128 B.n91 VSUBS 0.12501f
C129 B.n92 VSUBS 0.090582f
C130 B.n93 VSUBS 0.008795f
C131 B.n94 VSUBS 0.008795f
C132 B.n95 VSUBS 0.008795f
C133 B.n96 VSUBS 0.008795f
C134 B.n97 VSUBS 0.008795f
C135 B.n98 VSUBS 0.008795f
C136 B.n99 VSUBS 0.008795f
C137 B.n100 VSUBS 0.008795f
C138 B.n101 VSUBS 0.021147f
C139 B.n102 VSUBS 0.008795f
C140 B.n103 VSUBS 0.008795f
C141 B.n104 VSUBS 0.008795f
C142 B.n105 VSUBS 0.008795f
C143 B.n106 VSUBS 0.008795f
C144 B.n107 VSUBS 0.008795f
C145 B.n108 VSUBS 0.008795f
C146 B.n109 VSUBS 0.008795f
C147 B.n110 VSUBS 0.008795f
C148 B.n111 VSUBS 0.008795f
C149 B.n112 VSUBS 0.008795f
C150 B.n113 VSUBS 0.008795f
C151 B.n114 VSUBS 0.008795f
C152 B.n115 VSUBS 0.008795f
C153 B.n116 VSUBS 0.008795f
C154 B.n117 VSUBS 0.008795f
C155 B.n118 VSUBS 0.008795f
C156 B.n119 VSUBS 0.008795f
C157 B.n120 VSUBS 0.008795f
C158 B.n121 VSUBS 0.008795f
C159 B.n122 VSUBS 0.008795f
C160 B.n123 VSUBS 0.008795f
C161 B.n124 VSUBS 0.008795f
C162 B.n125 VSUBS 0.008795f
C163 B.n126 VSUBS 0.008795f
C164 B.n127 VSUBS 0.008795f
C165 B.n128 VSUBS 0.008795f
C166 B.n129 VSUBS 0.008795f
C167 B.n130 VSUBS 0.008795f
C168 B.n131 VSUBS 0.008795f
C169 B.n132 VSUBS 0.008795f
C170 B.n133 VSUBS 0.008795f
C171 B.n134 VSUBS 0.008795f
C172 B.n135 VSUBS 0.008795f
C173 B.n136 VSUBS 0.008795f
C174 B.n137 VSUBS 0.008795f
C175 B.n138 VSUBS 0.008795f
C176 B.n139 VSUBS 0.008795f
C177 B.n140 VSUBS 0.008795f
C178 B.n141 VSUBS 0.008795f
C179 B.n142 VSUBS 0.008795f
C180 B.n143 VSUBS 0.008795f
C181 B.n144 VSUBS 0.008795f
C182 B.n145 VSUBS 0.008795f
C183 B.n146 VSUBS 0.008795f
C184 B.n147 VSUBS 0.008795f
C185 B.n148 VSUBS 0.008795f
C186 B.n149 VSUBS 0.008795f
C187 B.n150 VSUBS 0.008795f
C188 B.n151 VSUBS 0.008795f
C189 B.n152 VSUBS 0.008795f
C190 B.n153 VSUBS 0.008795f
C191 B.n154 VSUBS 0.008795f
C192 B.n155 VSUBS 0.008795f
C193 B.n156 VSUBS 0.008795f
C194 B.n157 VSUBS 0.008795f
C195 B.n158 VSUBS 0.019465f
C196 B.n159 VSUBS 0.019465f
C197 B.n160 VSUBS 0.021147f
C198 B.n161 VSUBS 0.008795f
C199 B.n162 VSUBS 0.008795f
C200 B.n163 VSUBS 0.008795f
C201 B.n164 VSUBS 0.008795f
C202 B.n165 VSUBS 0.008795f
C203 B.n166 VSUBS 0.008795f
C204 B.n167 VSUBS 0.008795f
C205 B.n168 VSUBS 0.008795f
C206 B.n169 VSUBS 0.008795f
C207 B.n170 VSUBS 0.008795f
C208 B.n171 VSUBS 0.008795f
C209 B.n172 VSUBS 0.008795f
C210 B.n173 VSUBS 0.008795f
C211 B.n174 VSUBS 0.008795f
C212 B.n175 VSUBS 0.008795f
C213 B.n176 VSUBS 0.008795f
C214 B.n177 VSUBS 0.008795f
C215 B.n178 VSUBS 0.008795f
C216 B.n179 VSUBS 0.008795f
C217 B.n180 VSUBS 0.008795f
C218 B.n181 VSUBS 0.008795f
C219 B.n182 VSUBS 0.008795f
C220 B.n183 VSUBS 0.008795f
C221 B.n184 VSUBS 0.008795f
C222 B.n185 VSUBS 0.008795f
C223 B.n186 VSUBS 0.008795f
C224 B.n187 VSUBS 0.006079f
C225 B.n188 VSUBS 0.020377f
C226 B.n189 VSUBS 0.007114f
C227 B.n190 VSUBS 0.008795f
C228 B.n191 VSUBS 0.008795f
C229 B.n192 VSUBS 0.008795f
C230 B.n193 VSUBS 0.008795f
C231 B.n194 VSUBS 0.008795f
C232 B.n195 VSUBS 0.008795f
C233 B.n196 VSUBS 0.008795f
C234 B.n197 VSUBS 0.008795f
C235 B.n198 VSUBS 0.008795f
C236 B.n199 VSUBS 0.008795f
C237 B.n200 VSUBS 0.008795f
C238 B.t1 VSUBS 0.138183f
C239 B.t2 VSUBS 0.16761f
C240 B.t0 VSUBS 0.862802f
C241 B.n201 VSUBS 0.12501f
C242 B.n202 VSUBS 0.090582f
C243 B.n203 VSUBS 0.020377f
C244 B.n204 VSUBS 0.007114f
C245 B.n205 VSUBS 0.008795f
C246 B.n206 VSUBS 0.008795f
C247 B.n207 VSUBS 0.008795f
C248 B.n208 VSUBS 0.008795f
C249 B.n209 VSUBS 0.008795f
C250 B.n210 VSUBS 0.008795f
C251 B.n211 VSUBS 0.008795f
C252 B.n212 VSUBS 0.008795f
C253 B.n213 VSUBS 0.008795f
C254 B.n214 VSUBS 0.008795f
C255 B.n215 VSUBS 0.008795f
C256 B.n216 VSUBS 0.008795f
C257 B.n217 VSUBS 0.008795f
C258 B.n218 VSUBS 0.008795f
C259 B.n219 VSUBS 0.008795f
C260 B.n220 VSUBS 0.008795f
C261 B.n221 VSUBS 0.008795f
C262 B.n222 VSUBS 0.008795f
C263 B.n223 VSUBS 0.008795f
C264 B.n224 VSUBS 0.008795f
C265 B.n225 VSUBS 0.008795f
C266 B.n226 VSUBS 0.008795f
C267 B.n227 VSUBS 0.008795f
C268 B.n228 VSUBS 0.008795f
C269 B.n229 VSUBS 0.008795f
C270 B.n230 VSUBS 0.008795f
C271 B.n231 VSUBS 0.008795f
C272 B.n232 VSUBS 0.008795f
C273 B.n233 VSUBS 0.021147f
C274 B.n234 VSUBS 0.019465f
C275 B.n235 VSUBS 0.019465f
C276 B.n236 VSUBS 0.008795f
C277 B.n237 VSUBS 0.008795f
C278 B.n238 VSUBS 0.008795f
C279 B.n239 VSUBS 0.008795f
C280 B.n240 VSUBS 0.008795f
C281 B.n241 VSUBS 0.008795f
C282 B.n242 VSUBS 0.008795f
C283 B.n243 VSUBS 0.008795f
C284 B.n244 VSUBS 0.008795f
C285 B.n245 VSUBS 0.008795f
C286 B.n246 VSUBS 0.008795f
C287 B.n247 VSUBS 0.008795f
C288 B.n248 VSUBS 0.008795f
C289 B.n249 VSUBS 0.008795f
C290 B.n250 VSUBS 0.008795f
C291 B.n251 VSUBS 0.008795f
C292 B.n252 VSUBS 0.008795f
C293 B.n253 VSUBS 0.008795f
C294 B.n254 VSUBS 0.008795f
C295 B.n255 VSUBS 0.008795f
C296 B.n256 VSUBS 0.008795f
C297 B.n257 VSUBS 0.008795f
C298 B.n258 VSUBS 0.008795f
C299 B.n259 VSUBS 0.008795f
C300 B.n260 VSUBS 0.008795f
C301 B.n261 VSUBS 0.008795f
C302 B.n262 VSUBS 0.008795f
C303 B.n263 VSUBS 0.008795f
C304 B.n264 VSUBS 0.008795f
C305 B.n265 VSUBS 0.008795f
C306 B.n266 VSUBS 0.008795f
C307 B.n267 VSUBS 0.008795f
C308 B.n268 VSUBS 0.008795f
C309 B.n269 VSUBS 0.008795f
C310 B.n270 VSUBS 0.008795f
C311 B.n271 VSUBS 0.008795f
C312 B.n272 VSUBS 0.008795f
C313 B.n273 VSUBS 0.008795f
C314 B.n274 VSUBS 0.008795f
C315 B.n275 VSUBS 0.008795f
C316 B.n276 VSUBS 0.008795f
C317 B.n277 VSUBS 0.008795f
C318 B.n278 VSUBS 0.008795f
C319 B.n279 VSUBS 0.008795f
C320 B.n280 VSUBS 0.008795f
C321 B.n281 VSUBS 0.008795f
C322 B.n282 VSUBS 0.008795f
C323 B.n283 VSUBS 0.008795f
C324 B.n284 VSUBS 0.008795f
C325 B.n285 VSUBS 0.008795f
C326 B.n286 VSUBS 0.008795f
C327 B.n287 VSUBS 0.008795f
C328 B.n288 VSUBS 0.008795f
C329 B.n289 VSUBS 0.008795f
C330 B.n290 VSUBS 0.008795f
C331 B.n291 VSUBS 0.008795f
C332 B.n292 VSUBS 0.008795f
C333 B.n293 VSUBS 0.008795f
C334 B.n294 VSUBS 0.008795f
C335 B.n295 VSUBS 0.008795f
C336 B.n296 VSUBS 0.008795f
C337 B.n297 VSUBS 0.008795f
C338 B.n298 VSUBS 0.008795f
C339 B.n299 VSUBS 0.008795f
C340 B.n300 VSUBS 0.008795f
C341 B.n301 VSUBS 0.008795f
C342 B.n302 VSUBS 0.008795f
C343 B.n303 VSUBS 0.008795f
C344 B.n304 VSUBS 0.008795f
C345 B.n305 VSUBS 0.008795f
C346 B.n306 VSUBS 0.008795f
C347 B.n307 VSUBS 0.008795f
C348 B.n308 VSUBS 0.008795f
C349 B.n309 VSUBS 0.008795f
C350 B.n310 VSUBS 0.008795f
C351 B.n311 VSUBS 0.008795f
C352 B.n312 VSUBS 0.008795f
C353 B.n313 VSUBS 0.008795f
C354 B.n314 VSUBS 0.008795f
C355 B.n315 VSUBS 0.008795f
C356 B.n316 VSUBS 0.008795f
C357 B.n317 VSUBS 0.008795f
C358 B.n318 VSUBS 0.008795f
C359 B.n319 VSUBS 0.008795f
C360 B.n320 VSUBS 0.008795f
C361 B.n321 VSUBS 0.008795f
C362 B.n322 VSUBS 0.008795f
C363 B.n323 VSUBS 0.008795f
C364 B.n324 VSUBS 0.020526f
C365 B.n325 VSUBS 0.019465f
C366 B.n326 VSUBS 0.021147f
C367 B.n327 VSUBS 0.008795f
C368 B.n328 VSUBS 0.008795f
C369 B.n329 VSUBS 0.008795f
C370 B.n330 VSUBS 0.008795f
C371 B.n331 VSUBS 0.008795f
C372 B.n332 VSUBS 0.008795f
C373 B.n333 VSUBS 0.008795f
C374 B.n334 VSUBS 0.008795f
C375 B.n335 VSUBS 0.008795f
C376 B.n336 VSUBS 0.008795f
C377 B.n337 VSUBS 0.008795f
C378 B.n338 VSUBS 0.008795f
C379 B.n339 VSUBS 0.008795f
C380 B.n340 VSUBS 0.008795f
C381 B.n341 VSUBS 0.008795f
C382 B.n342 VSUBS 0.008795f
C383 B.n343 VSUBS 0.008795f
C384 B.n344 VSUBS 0.008795f
C385 B.n345 VSUBS 0.008795f
C386 B.n346 VSUBS 0.008795f
C387 B.n347 VSUBS 0.008795f
C388 B.n348 VSUBS 0.008795f
C389 B.n349 VSUBS 0.008795f
C390 B.n350 VSUBS 0.008795f
C391 B.n351 VSUBS 0.008795f
C392 B.n352 VSUBS 0.008795f
C393 B.n353 VSUBS 0.006079f
C394 B.n354 VSUBS 0.020377f
C395 B.n355 VSUBS 0.007114f
C396 B.n356 VSUBS 0.008795f
C397 B.n357 VSUBS 0.008795f
C398 B.n358 VSUBS 0.008795f
C399 B.n359 VSUBS 0.008795f
C400 B.n360 VSUBS 0.008795f
C401 B.n361 VSUBS 0.008795f
C402 B.n362 VSUBS 0.008795f
C403 B.n363 VSUBS 0.008795f
C404 B.n364 VSUBS 0.008795f
C405 B.n365 VSUBS 0.008795f
C406 B.n366 VSUBS 0.008795f
C407 B.n367 VSUBS 0.007114f
C408 B.n368 VSUBS 0.008795f
C409 B.n369 VSUBS 0.008795f
C410 B.n370 VSUBS 0.008795f
C411 B.n371 VSUBS 0.008795f
C412 B.n372 VSUBS 0.008795f
C413 B.n373 VSUBS 0.008795f
C414 B.n374 VSUBS 0.008795f
C415 B.n375 VSUBS 0.008795f
C416 B.n376 VSUBS 0.008795f
C417 B.n377 VSUBS 0.008795f
C418 B.n378 VSUBS 0.008795f
C419 B.n379 VSUBS 0.008795f
C420 B.n380 VSUBS 0.008795f
C421 B.n381 VSUBS 0.008795f
C422 B.n382 VSUBS 0.008795f
C423 B.n383 VSUBS 0.008795f
C424 B.n384 VSUBS 0.008795f
C425 B.n385 VSUBS 0.008795f
C426 B.n386 VSUBS 0.008795f
C427 B.n387 VSUBS 0.008795f
C428 B.n388 VSUBS 0.008795f
C429 B.n389 VSUBS 0.008795f
C430 B.n390 VSUBS 0.008795f
C431 B.n391 VSUBS 0.008795f
C432 B.n392 VSUBS 0.008795f
C433 B.n393 VSUBS 0.008795f
C434 B.n394 VSUBS 0.008795f
C435 B.n395 VSUBS 0.008795f
C436 B.n396 VSUBS 0.021147f
C437 B.n397 VSUBS 0.019465f
C438 B.n398 VSUBS 0.019465f
C439 B.n399 VSUBS 0.008795f
C440 B.n400 VSUBS 0.008795f
C441 B.n401 VSUBS 0.008795f
C442 B.n402 VSUBS 0.008795f
C443 B.n403 VSUBS 0.008795f
C444 B.n404 VSUBS 0.008795f
C445 B.n405 VSUBS 0.008795f
C446 B.n406 VSUBS 0.008795f
C447 B.n407 VSUBS 0.008795f
C448 B.n408 VSUBS 0.008795f
C449 B.n409 VSUBS 0.008795f
C450 B.n410 VSUBS 0.008795f
C451 B.n411 VSUBS 0.008795f
C452 B.n412 VSUBS 0.008795f
C453 B.n413 VSUBS 0.008795f
C454 B.n414 VSUBS 0.008795f
C455 B.n415 VSUBS 0.008795f
C456 B.n416 VSUBS 0.008795f
C457 B.n417 VSUBS 0.008795f
C458 B.n418 VSUBS 0.008795f
C459 B.n419 VSUBS 0.008795f
C460 B.n420 VSUBS 0.008795f
C461 B.n421 VSUBS 0.008795f
C462 B.n422 VSUBS 0.008795f
C463 B.n423 VSUBS 0.008795f
C464 B.n424 VSUBS 0.008795f
C465 B.n425 VSUBS 0.008795f
C466 B.n426 VSUBS 0.008795f
C467 B.n427 VSUBS 0.008795f
C468 B.n428 VSUBS 0.008795f
C469 B.n429 VSUBS 0.008795f
C470 B.n430 VSUBS 0.008795f
C471 B.n431 VSUBS 0.008795f
C472 B.n432 VSUBS 0.008795f
C473 B.n433 VSUBS 0.008795f
C474 B.n434 VSUBS 0.008795f
C475 B.n435 VSUBS 0.008795f
C476 B.n436 VSUBS 0.008795f
C477 B.n437 VSUBS 0.008795f
C478 B.n438 VSUBS 0.008795f
C479 B.n439 VSUBS 0.008795f
C480 B.n440 VSUBS 0.008795f
C481 B.n441 VSUBS 0.008795f
C482 B.n442 VSUBS 0.008795f
C483 B.n443 VSUBS 0.019915f
C484 VDD1.t1 VSUBS 0.410615f
C485 VDD1.t0 VSUBS 0.63859f
C486 VP.t0 VSUBS 2.65052f
C487 VP.t1 VSUBS 1.84953f
C488 VP.n0 VSUBS 3.36261f
C489 VDD2.t0 VSUBS 0.650309f
C490 VDD2.t1 VSUBS 0.428778f
C491 VDD2.n0 VSUBS 2.09126f
C492 VTAIL.t0 VSUBS 0.578604f
C493 VTAIL.n0 VSUBS 1.63909f
C494 VTAIL.t2 VSUBS 0.578607f
C495 VTAIL.n1 VSUBS 1.69768f
C496 VTAIL.t1 VSUBS 0.578604f
C497 VTAIL.n2 VSUBS 1.44511f
C498 VTAIL.t3 VSUBS 0.578604f
C499 VTAIL.n3 VSUBS 1.34071f
C500 VN.t1 VSUBS 1.77294f
C501 VN.t0 VSUBS 2.53548f
.ends

