* NGSPICE file created from diff_pair_sample_0255.ext - technology: sky130A

.subckt diff_pair_sample_0255 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7761 pd=4.76 as=0.7761 ps=4.76 w=1.99 l=2.74
X1 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7761 pd=4.76 as=0.7761 ps=4.76 w=1.99 l=2.74
X2 VDD2.t1 VN.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7761 pd=4.76 as=0.7761 ps=4.76 w=1.99 l=2.74
X3 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=0.7761 pd=4.76 as=0 ps=0 w=1.99 l=2.74
X4 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=0.7761 pd=4.76 as=0 ps=0 w=1.99 l=2.74
X5 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7761 pd=4.76 as=0 ps=0 w=1.99 l=2.74
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7761 pd=4.76 as=0 ps=0 w=1.99 l=2.74
X7 VDD2.t0 VN.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7761 pd=4.76 as=0.7761 ps=4.76 w=1.99 l=2.74
R0 VP.n0 VP.t1 96.0443
R1 VP.n0 VP.t0 58.5995
R2 VP VP.n0 0.431811
R3 VTAIL.n26 VTAIL.n24 289.615
R4 VTAIL.n2 VTAIL.n0 289.615
R5 VTAIL.n18 VTAIL.n16 289.615
R6 VTAIL.n10 VTAIL.n8 289.615
R7 VTAIL.n27 VTAIL.n26 185
R8 VTAIL.n3 VTAIL.n2 185
R9 VTAIL.n19 VTAIL.n18 185
R10 VTAIL.n11 VTAIL.n10 185
R11 VTAIL.t3 VTAIL.n25 167.117
R12 VTAIL.t1 VTAIL.n1 167.117
R13 VTAIL.t0 VTAIL.n17 167.117
R14 VTAIL.t2 VTAIL.n9 167.117
R15 VTAIL.n26 VTAIL.t3 52.3082
R16 VTAIL.n2 VTAIL.t1 52.3082
R17 VTAIL.n18 VTAIL.t0 52.3082
R18 VTAIL.n10 VTAIL.t2 52.3082
R19 VTAIL.n31 VTAIL.n30 31.2157
R20 VTAIL.n7 VTAIL.n6 31.2157
R21 VTAIL.n23 VTAIL.n22 31.2157
R22 VTAIL.n15 VTAIL.n14 31.2157
R23 VTAIL.n15 VTAIL.n7 19.3755
R24 VTAIL.n31 VTAIL.n23 16.7289
R25 VTAIL.n27 VTAIL.n25 9.71174
R26 VTAIL.n3 VTAIL.n1 9.71174
R27 VTAIL.n19 VTAIL.n17 9.71174
R28 VTAIL.n11 VTAIL.n9 9.71174
R29 VTAIL.n30 VTAIL.n29 9.45567
R30 VTAIL.n6 VTAIL.n5 9.45567
R31 VTAIL.n22 VTAIL.n21 9.45567
R32 VTAIL.n14 VTAIL.n13 9.45567
R33 VTAIL.n29 VTAIL.n28 9.3005
R34 VTAIL.n5 VTAIL.n4 9.3005
R35 VTAIL.n21 VTAIL.n20 9.3005
R36 VTAIL.n13 VTAIL.n12 9.3005
R37 VTAIL.n30 VTAIL.n24 8.14595
R38 VTAIL.n6 VTAIL.n0 8.14595
R39 VTAIL.n22 VTAIL.n16 8.14595
R40 VTAIL.n14 VTAIL.n8 8.14595
R41 VTAIL.n28 VTAIL.n27 7.3702
R42 VTAIL.n4 VTAIL.n3 7.3702
R43 VTAIL.n20 VTAIL.n19 7.3702
R44 VTAIL.n12 VTAIL.n11 7.3702
R45 VTAIL.n28 VTAIL.n24 5.81868
R46 VTAIL.n4 VTAIL.n0 5.81868
R47 VTAIL.n20 VTAIL.n16 5.81868
R48 VTAIL.n12 VTAIL.n8 5.81868
R49 VTAIL.n29 VTAIL.n25 3.44771
R50 VTAIL.n5 VTAIL.n1 3.44771
R51 VTAIL.n21 VTAIL.n17 3.44771
R52 VTAIL.n13 VTAIL.n9 3.44771
R53 VTAIL.n23 VTAIL.n15 1.7936
R54 VTAIL VTAIL.n7 1.19016
R55 VTAIL VTAIL.n31 0.603948
R56 VDD1.n2 VDD1.n0 289.615
R57 VDD1.n9 VDD1.n7 289.615
R58 VDD1.n3 VDD1.n2 185
R59 VDD1.n10 VDD1.n9 185
R60 VDD1.t0 VDD1.n1 167.117
R61 VDD1.t1 VDD1.n8 167.117
R62 VDD1 VDD1.n13 79.749
R63 VDD1.n2 VDD1.t0 52.3082
R64 VDD1.n9 VDD1.t1 52.3082
R65 VDD1 VDD1.n6 48.6143
R66 VDD1.n3 VDD1.n1 9.71174
R67 VDD1.n10 VDD1.n8 9.71174
R68 VDD1.n6 VDD1.n5 9.45567
R69 VDD1.n13 VDD1.n12 9.45567
R70 VDD1.n5 VDD1.n4 9.3005
R71 VDD1.n12 VDD1.n11 9.3005
R72 VDD1.n6 VDD1.n0 8.14595
R73 VDD1.n13 VDD1.n7 8.14595
R74 VDD1.n4 VDD1.n3 7.3702
R75 VDD1.n11 VDD1.n10 7.3702
R76 VDD1.n4 VDD1.n0 5.81868
R77 VDD1.n11 VDD1.n7 5.81868
R78 VDD1.n5 VDD1.n1 3.44771
R79 VDD1.n12 VDD1.n8 3.44771
R80 B.n325 B.n324 585
R81 B.n327 B.n72 585
R82 B.n330 B.n329 585
R83 B.n331 B.n71 585
R84 B.n333 B.n332 585
R85 B.n335 B.n70 585
R86 B.n338 B.n337 585
R87 B.n339 B.n69 585
R88 B.n341 B.n340 585
R89 B.n343 B.n68 585
R90 B.n345 B.n344 585
R91 B.n347 B.n346 585
R92 B.n350 B.n349 585
R93 B.n351 B.n63 585
R94 B.n353 B.n352 585
R95 B.n355 B.n62 585
R96 B.n358 B.n357 585
R97 B.n359 B.n61 585
R98 B.n361 B.n360 585
R99 B.n363 B.n60 585
R100 B.n366 B.n365 585
R101 B.n367 B.n57 585
R102 B.n370 B.n369 585
R103 B.n372 B.n56 585
R104 B.n375 B.n374 585
R105 B.n376 B.n55 585
R106 B.n378 B.n377 585
R107 B.n380 B.n54 585
R108 B.n383 B.n382 585
R109 B.n384 B.n53 585
R110 B.n386 B.n385 585
R111 B.n388 B.n52 585
R112 B.n391 B.n390 585
R113 B.n392 B.n51 585
R114 B.n323 B.n49 585
R115 B.n395 B.n49 585
R116 B.n322 B.n48 585
R117 B.n396 B.n48 585
R118 B.n321 B.n47 585
R119 B.n397 B.n47 585
R120 B.n320 B.n319 585
R121 B.n319 B.n43 585
R122 B.n318 B.n42 585
R123 B.n403 B.n42 585
R124 B.n317 B.n41 585
R125 B.n404 B.n41 585
R126 B.n316 B.n40 585
R127 B.n405 B.n40 585
R128 B.n315 B.n314 585
R129 B.n314 B.n39 585
R130 B.n313 B.n35 585
R131 B.n411 B.n35 585
R132 B.n312 B.n34 585
R133 B.n412 B.n34 585
R134 B.n311 B.n33 585
R135 B.n413 B.n33 585
R136 B.n310 B.n309 585
R137 B.n309 B.n29 585
R138 B.n308 B.n28 585
R139 B.n419 B.n28 585
R140 B.n307 B.n27 585
R141 B.n420 B.n27 585
R142 B.n306 B.n26 585
R143 B.n421 B.n26 585
R144 B.n305 B.n304 585
R145 B.n304 B.n22 585
R146 B.n303 B.n21 585
R147 B.n427 B.n21 585
R148 B.n302 B.n20 585
R149 B.n428 B.n20 585
R150 B.n301 B.n19 585
R151 B.n429 B.n19 585
R152 B.n300 B.n299 585
R153 B.n299 B.n18 585
R154 B.n298 B.n14 585
R155 B.n435 B.n14 585
R156 B.n297 B.n13 585
R157 B.n436 B.n13 585
R158 B.n296 B.n12 585
R159 B.n437 B.n12 585
R160 B.n295 B.n294 585
R161 B.n294 B.n8 585
R162 B.n293 B.n7 585
R163 B.n443 B.n7 585
R164 B.n292 B.n6 585
R165 B.n444 B.n6 585
R166 B.n291 B.n5 585
R167 B.n445 B.n5 585
R168 B.n290 B.n289 585
R169 B.n289 B.n4 585
R170 B.n288 B.n73 585
R171 B.n288 B.n287 585
R172 B.n278 B.n74 585
R173 B.n75 B.n74 585
R174 B.n280 B.n279 585
R175 B.n281 B.n280 585
R176 B.n277 B.n80 585
R177 B.n80 B.n79 585
R178 B.n276 B.n275 585
R179 B.n275 B.n274 585
R180 B.n82 B.n81 585
R181 B.n267 B.n82 585
R182 B.n266 B.n265 585
R183 B.n268 B.n266 585
R184 B.n264 B.n87 585
R185 B.n87 B.n86 585
R186 B.n263 B.n262 585
R187 B.n262 B.n261 585
R188 B.n89 B.n88 585
R189 B.n90 B.n89 585
R190 B.n254 B.n253 585
R191 B.n255 B.n254 585
R192 B.n252 B.n95 585
R193 B.n95 B.n94 585
R194 B.n251 B.n250 585
R195 B.n250 B.n249 585
R196 B.n97 B.n96 585
R197 B.n98 B.n97 585
R198 B.n242 B.n241 585
R199 B.n243 B.n242 585
R200 B.n240 B.n103 585
R201 B.n103 B.n102 585
R202 B.n239 B.n238 585
R203 B.n238 B.n237 585
R204 B.n105 B.n104 585
R205 B.n230 B.n105 585
R206 B.n229 B.n228 585
R207 B.n231 B.n229 585
R208 B.n227 B.n110 585
R209 B.n110 B.n109 585
R210 B.n226 B.n225 585
R211 B.n225 B.n224 585
R212 B.n112 B.n111 585
R213 B.n113 B.n112 585
R214 B.n217 B.n216 585
R215 B.n218 B.n217 585
R216 B.n215 B.n118 585
R217 B.n118 B.n117 585
R218 B.n214 B.n213 585
R219 B.n213 B.n212 585
R220 B.n209 B.n122 585
R221 B.n208 B.n207 585
R222 B.n205 B.n123 585
R223 B.n205 B.n121 585
R224 B.n204 B.n203 585
R225 B.n202 B.n201 585
R226 B.n200 B.n125 585
R227 B.n198 B.n197 585
R228 B.n196 B.n126 585
R229 B.n195 B.n194 585
R230 B.n192 B.n127 585
R231 B.n190 B.n189 585
R232 B.n188 B.n128 585
R233 B.n186 B.n185 585
R234 B.n183 B.n131 585
R235 B.n181 B.n180 585
R236 B.n179 B.n132 585
R237 B.n178 B.n177 585
R238 B.n175 B.n133 585
R239 B.n173 B.n172 585
R240 B.n171 B.n134 585
R241 B.n170 B.n169 585
R242 B.n167 B.n135 585
R243 B.n165 B.n164 585
R244 B.n163 B.n136 585
R245 B.n162 B.n161 585
R246 B.n159 B.n140 585
R247 B.n157 B.n156 585
R248 B.n155 B.n141 585
R249 B.n154 B.n153 585
R250 B.n151 B.n142 585
R251 B.n149 B.n148 585
R252 B.n147 B.n143 585
R253 B.n146 B.n145 585
R254 B.n120 B.n119 585
R255 B.n121 B.n120 585
R256 B.n211 B.n210 585
R257 B.n212 B.n211 585
R258 B.n116 B.n115 585
R259 B.n117 B.n116 585
R260 B.n220 B.n219 585
R261 B.n219 B.n218 585
R262 B.n221 B.n114 585
R263 B.n114 B.n113 585
R264 B.n223 B.n222 585
R265 B.n224 B.n223 585
R266 B.n108 B.n107 585
R267 B.n109 B.n108 585
R268 B.n233 B.n232 585
R269 B.n232 B.n231 585
R270 B.n234 B.n106 585
R271 B.n230 B.n106 585
R272 B.n236 B.n235 585
R273 B.n237 B.n236 585
R274 B.n101 B.n100 585
R275 B.n102 B.n101 585
R276 B.n245 B.n244 585
R277 B.n244 B.n243 585
R278 B.n246 B.n99 585
R279 B.n99 B.n98 585
R280 B.n248 B.n247 585
R281 B.n249 B.n248 585
R282 B.n93 B.n92 585
R283 B.n94 B.n93 585
R284 B.n257 B.n256 585
R285 B.n256 B.n255 585
R286 B.n258 B.n91 585
R287 B.n91 B.n90 585
R288 B.n260 B.n259 585
R289 B.n261 B.n260 585
R290 B.n85 B.n84 585
R291 B.n86 B.n85 585
R292 B.n270 B.n269 585
R293 B.n269 B.n268 585
R294 B.n271 B.n83 585
R295 B.n267 B.n83 585
R296 B.n273 B.n272 585
R297 B.n274 B.n273 585
R298 B.n78 B.n77 585
R299 B.n79 B.n78 585
R300 B.n283 B.n282 585
R301 B.n282 B.n281 585
R302 B.n284 B.n76 585
R303 B.n76 B.n75 585
R304 B.n286 B.n285 585
R305 B.n287 B.n286 585
R306 B.n2 B.n0 585
R307 B.n4 B.n2 585
R308 B.n3 B.n1 585
R309 B.n444 B.n3 585
R310 B.n442 B.n441 585
R311 B.n443 B.n442 585
R312 B.n440 B.n9 585
R313 B.n9 B.n8 585
R314 B.n439 B.n438 585
R315 B.n438 B.n437 585
R316 B.n11 B.n10 585
R317 B.n436 B.n11 585
R318 B.n434 B.n433 585
R319 B.n435 B.n434 585
R320 B.n432 B.n15 585
R321 B.n18 B.n15 585
R322 B.n431 B.n430 585
R323 B.n430 B.n429 585
R324 B.n17 B.n16 585
R325 B.n428 B.n17 585
R326 B.n426 B.n425 585
R327 B.n427 B.n426 585
R328 B.n424 B.n23 585
R329 B.n23 B.n22 585
R330 B.n423 B.n422 585
R331 B.n422 B.n421 585
R332 B.n25 B.n24 585
R333 B.n420 B.n25 585
R334 B.n418 B.n417 585
R335 B.n419 B.n418 585
R336 B.n416 B.n30 585
R337 B.n30 B.n29 585
R338 B.n415 B.n414 585
R339 B.n414 B.n413 585
R340 B.n32 B.n31 585
R341 B.n412 B.n32 585
R342 B.n410 B.n409 585
R343 B.n411 B.n410 585
R344 B.n408 B.n36 585
R345 B.n39 B.n36 585
R346 B.n407 B.n406 585
R347 B.n406 B.n405 585
R348 B.n38 B.n37 585
R349 B.n404 B.n38 585
R350 B.n402 B.n401 585
R351 B.n403 B.n402 585
R352 B.n400 B.n44 585
R353 B.n44 B.n43 585
R354 B.n399 B.n398 585
R355 B.n398 B.n397 585
R356 B.n46 B.n45 585
R357 B.n396 B.n46 585
R358 B.n394 B.n393 585
R359 B.n395 B.n394 585
R360 B.n447 B.n446 585
R361 B.n446 B.n445 585
R362 B.n211 B.n122 521.33
R363 B.n394 B.n51 521.33
R364 B.n213 B.n120 521.33
R365 B.n325 B.n49 521.33
R366 B.n326 B.n50 256.663
R367 B.n328 B.n50 256.663
R368 B.n334 B.n50 256.663
R369 B.n336 B.n50 256.663
R370 B.n342 B.n50 256.663
R371 B.n67 B.n50 256.663
R372 B.n348 B.n50 256.663
R373 B.n354 B.n50 256.663
R374 B.n356 B.n50 256.663
R375 B.n362 B.n50 256.663
R376 B.n364 B.n50 256.663
R377 B.n371 B.n50 256.663
R378 B.n373 B.n50 256.663
R379 B.n379 B.n50 256.663
R380 B.n381 B.n50 256.663
R381 B.n387 B.n50 256.663
R382 B.n389 B.n50 256.663
R383 B.n206 B.n121 256.663
R384 B.n124 B.n121 256.663
R385 B.n199 B.n121 256.663
R386 B.n193 B.n121 256.663
R387 B.n191 B.n121 256.663
R388 B.n184 B.n121 256.663
R389 B.n182 B.n121 256.663
R390 B.n176 B.n121 256.663
R391 B.n174 B.n121 256.663
R392 B.n168 B.n121 256.663
R393 B.n166 B.n121 256.663
R394 B.n160 B.n121 256.663
R395 B.n158 B.n121 256.663
R396 B.n152 B.n121 256.663
R397 B.n150 B.n121 256.663
R398 B.n144 B.n121 256.663
R399 B.n137 B.t2 225.752
R400 B.n129 B.t6 225.752
R401 B.n58 B.t9 225.752
R402 B.n64 B.t13 225.752
R403 B.n212 B.n121 204.405
R404 B.n395 B.n50 204.405
R405 B.n137 B.t5 182.363
R406 B.n64 B.t14 182.363
R407 B.n129 B.t8 182.363
R408 B.n58 B.t11 182.363
R409 B.n211 B.n116 163.367
R410 B.n219 B.n116 163.367
R411 B.n219 B.n114 163.367
R412 B.n223 B.n114 163.367
R413 B.n223 B.n108 163.367
R414 B.n232 B.n108 163.367
R415 B.n232 B.n106 163.367
R416 B.n236 B.n106 163.367
R417 B.n236 B.n101 163.367
R418 B.n244 B.n101 163.367
R419 B.n244 B.n99 163.367
R420 B.n248 B.n99 163.367
R421 B.n248 B.n93 163.367
R422 B.n256 B.n93 163.367
R423 B.n256 B.n91 163.367
R424 B.n260 B.n91 163.367
R425 B.n260 B.n85 163.367
R426 B.n269 B.n85 163.367
R427 B.n269 B.n83 163.367
R428 B.n273 B.n83 163.367
R429 B.n273 B.n78 163.367
R430 B.n282 B.n78 163.367
R431 B.n282 B.n76 163.367
R432 B.n286 B.n76 163.367
R433 B.n286 B.n2 163.367
R434 B.n446 B.n2 163.367
R435 B.n446 B.n3 163.367
R436 B.n442 B.n3 163.367
R437 B.n442 B.n9 163.367
R438 B.n438 B.n9 163.367
R439 B.n438 B.n11 163.367
R440 B.n434 B.n11 163.367
R441 B.n434 B.n15 163.367
R442 B.n430 B.n15 163.367
R443 B.n430 B.n17 163.367
R444 B.n426 B.n17 163.367
R445 B.n426 B.n23 163.367
R446 B.n422 B.n23 163.367
R447 B.n422 B.n25 163.367
R448 B.n418 B.n25 163.367
R449 B.n418 B.n30 163.367
R450 B.n414 B.n30 163.367
R451 B.n414 B.n32 163.367
R452 B.n410 B.n32 163.367
R453 B.n410 B.n36 163.367
R454 B.n406 B.n36 163.367
R455 B.n406 B.n38 163.367
R456 B.n402 B.n38 163.367
R457 B.n402 B.n44 163.367
R458 B.n398 B.n44 163.367
R459 B.n398 B.n46 163.367
R460 B.n394 B.n46 163.367
R461 B.n207 B.n205 163.367
R462 B.n205 B.n204 163.367
R463 B.n201 B.n200 163.367
R464 B.n198 B.n126 163.367
R465 B.n194 B.n192 163.367
R466 B.n190 B.n128 163.367
R467 B.n185 B.n183 163.367
R468 B.n181 B.n132 163.367
R469 B.n177 B.n175 163.367
R470 B.n173 B.n134 163.367
R471 B.n169 B.n167 163.367
R472 B.n165 B.n136 163.367
R473 B.n161 B.n159 163.367
R474 B.n157 B.n141 163.367
R475 B.n153 B.n151 163.367
R476 B.n149 B.n143 163.367
R477 B.n145 B.n120 163.367
R478 B.n213 B.n118 163.367
R479 B.n217 B.n118 163.367
R480 B.n217 B.n112 163.367
R481 B.n225 B.n112 163.367
R482 B.n225 B.n110 163.367
R483 B.n229 B.n110 163.367
R484 B.n229 B.n105 163.367
R485 B.n238 B.n105 163.367
R486 B.n238 B.n103 163.367
R487 B.n242 B.n103 163.367
R488 B.n242 B.n97 163.367
R489 B.n250 B.n97 163.367
R490 B.n250 B.n95 163.367
R491 B.n254 B.n95 163.367
R492 B.n254 B.n89 163.367
R493 B.n262 B.n89 163.367
R494 B.n262 B.n87 163.367
R495 B.n266 B.n87 163.367
R496 B.n266 B.n82 163.367
R497 B.n275 B.n82 163.367
R498 B.n275 B.n80 163.367
R499 B.n280 B.n80 163.367
R500 B.n280 B.n74 163.367
R501 B.n288 B.n74 163.367
R502 B.n289 B.n288 163.367
R503 B.n289 B.n5 163.367
R504 B.n6 B.n5 163.367
R505 B.n7 B.n6 163.367
R506 B.n294 B.n7 163.367
R507 B.n294 B.n12 163.367
R508 B.n13 B.n12 163.367
R509 B.n14 B.n13 163.367
R510 B.n299 B.n14 163.367
R511 B.n299 B.n19 163.367
R512 B.n20 B.n19 163.367
R513 B.n21 B.n20 163.367
R514 B.n304 B.n21 163.367
R515 B.n304 B.n26 163.367
R516 B.n27 B.n26 163.367
R517 B.n28 B.n27 163.367
R518 B.n309 B.n28 163.367
R519 B.n309 B.n33 163.367
R520 B.n34 B.n33 163.367
R521 B.n35 B.n34 163.367
R522 B.n314 B.n35 163.367
R523 B.n314 B.n40 163.367
R524 B.n41 B.n40 163.367
R525 B.n42 B.n41 163.367
R526 B.n319 B.n42 163.367
R527 B.n319 B.n47 163.367
R528 B.n48 B.n47 163.367
R529 B.n49 B.n48 163.367
R530 B.n390 B.n388 163.367
R531 B.n386 B.n53 163.367
R532 B.n382 B.n380 163.367
R533 B.n378 B.n55 163.367
R534 B.n374 B.n372 163.367
R535 B.n370 B.n57 163.367
R536 B.n365 B.n363 163.367
R537 B.n361 B.n61 163.367
R538 B.n357 B.n355 163.367
R539 B.n353 B.n63 163.367
R540 B.n349 B.n347 163.367
R541 B.n344 B.n343 163.367
R542 B.n341 B.n69 163.367
R543 B.n337 B.n335 163.367
R544 B.n333 B.n71 163.367
R545 B.n329 B.n327 163.367
R546 B.n138 B.t4 122.825
R547 B.n65 B.t15 122.825
R548 B.n130 B.t7 122.825
R549 B.n59 B.t12 122.825
R550 B.n212 B.n117 102.96
R551 B.n218 B.n117 102.96
R552 B.n218 B.n113 102.96
R553 B.n224 B.n113 102.96
R554 B.n224 B.n109 102.96
R555 B.n231 B.n109 102.96
R556 B.n231 B.n230 102.96
R557 B.n237 B.n102 102.96
R558 B.n243 B.n102 102.96
R559 B.n243 B.n98 102.96
R560 B.n249 B.n98 102.96
R561 B.n249 B.n94 102.96
R562 B.n255 B.n94 102.96
R563 B.n255 B.n90 102.96
R564 B.n261 B.n90 102.96
R565 B.n261 B.n86 102.96
R566 B.n268 B.n86 102.96
R567 B.n268 B.n267 102.96
R568 B.n274 B.n79 102.96
R569 B.n281 B.n79 102.96
R570 B.n281 B.n75 102.96
R571 B.n287 B.n75 102.96
R572 B.n287 B.n4 102.96
R573 B.n445 B.n4 102.96
R574 B.n445 B.n444 102.96
R575 B.n444 B.n443 102.96
R576 B.n443 B.n8 102.96
R577 B.n437 B.n8 102.96
R578 B.n437 B.n436 102.96
R579 B.n436 B.n435 102.96
R580 B.n429 B.n18 102.96
R581 B.n429 B.n428 102.96
R582 B.n428 B.n427 102.96
R583 B.n427 B.n22 102.96
R584 B.n421 B.n22 102.96
R585 B.n421 B.n420 102.96
R586 B.n420 B.n419 102.96
R587 B.n419 B.n29 102.96
R588 B.n413 B.n29 102.96
R589 B.n413 B.n412 102.96
R590 B.n412 B.n411 102.96
R591 B.n405 B.n39 102.96
R592 B.n405 B.n404 102.96
R593 B.n404 B.n403 102.96
R594 B.n403 B.n43 102.96
R595 B.n397 B.n43 102.96
R596 B.n397 B.n396 102.96
R597 B.n396 B.n395 102.96
R598 B.n267 B.t1 90.847
R599 B.n18 B.t0 90.847
R600 B.n206 B.n122 71.676
R601 B.n204 B.n124 71.676
R602 B.n200 B.n199 71.676
R603 B.n193 B.n126 71.676
R604 B.n192 B.n191 71.676
R605 B.n184 B.n128 71.676
R606 B.n183 B.n182 71.676
R607 B.n176 B.n132 71.676
R608 B.n175 B.n174 71.676
R609 B.n168 B.n134 71.676
R610 B.n167 B.n166 71.676
R611 B.n160 B.n136 71.676
R612 B.n159 B.n158 71.676
R613 B.n152 B.n141 71.676
R614 B.n151 B.n150 71.676
R615 B.n144 B.n143 71.676
R616 B.n389 B.n51 71.676
R617 B.n388 B.n387 71.676
R618 B.n381 B.n53 71.676
R619 B.n380 B.n379 71.676
R620 B.n373 B.n55 71.676
R621 B.n372 B.n371 71.676
R622 B.n364 B.n57 71.676
R623 B.n363 B.n362 71.676
R624 B.n356 B.n61 71.676
R625 B.n355 B.n354 71.676
R626 B.n348 B.n63 71.676
R627 B.n347 B.n67 71.676
R628 B.n343 B.n342 71.676
R629 B.n336 B.n69 71.676
R630 B.n335 B.n334 71.676
R631 B.n328 B.n71 71.676
R632 B.n327 B.n326 71.676
R633 B.n326 B.n325 71.676
R634 B.n329 B.n328 71.676
R635 B.n334 B.n333 71.676
R636 B.n337 B.n336 71.676
R637 B.n342 B.n341 71.676
R638 B.n344 B.n67 71.676
R639 B.n349 B.n348 71.676
R640 B.n354 B.n353 71.676
R641 B.n357 B.n356 71.676
R642 B.n362 B.n361 71.676
R643 B.n365 B.n364 71.676
R644 B.n371 B.n370 71.676
R645 B.n374 B.n373 71.676
R646 B.n379 B.n378 71.676
R647 B.n382 B.n381 71.676
R648 B.n387 B.n386 71.676
R649 B.n390 B.n389 71.676
R650 B.n207 B.n206 71.676
R651 B.n201 B.n124 71.676
R652 B.n199 B.n198 71.676
R653 B.n194 B.n193 71.676
R654 B.n191 B.n190 71.676
R655 B.n185 B.n184 71.676
R656 B.n182 B.n181 71.676
R657 B.n177 B.n176 71.676
R658 B.n174 B.n173 71.676
R659 B.n169 B.n168 71.676
R660 B.n166 B.n165 71.676
R661 B.n161 B.n160 71.676
R662 B.n158 B.n157 71.676
R663 B.n153 B.n152 71.676
R664 B.n150 B.n149 71.676
R665 B.n145 B.n144 71.676
R666 B.n230 B.t3 66.6213
R667 B.n39 B.t10 66.6213
R668 B.n139 B.n138 59.5399
R669 B.n138 B.n137 59.5399
R670 B.n187 B.n130 59.5399
R671 B.n130 B.n129 59.5399
R672 B.n59 B.n58 59.5399
R673 B.n368 B.n59 59.5399
R674 B.n65 B.n64 59.5399
R675 B.n66 B.n65 59.5399
R676 B.n237 B.t3 36.3391
R677 B.n411 B.t10 36.3391
R678 B.n393 B.n392 33.8737
R679 B.n324 B.n323 33.8737
R680 B.n214 B.n119 33.8737
R681 B.n210 B.n209 33.8737
R682 B B.n447 18.0485
R683 B.n274 B.t1 12.1134
R684 B.n435 B.t0 12.1134
R685 B.n392 B.n391 10.6151
R686 B.n391 B.n52 10.6151
R687 B.n385 B.n52 10.6151
R688 B.n385 B.n384 10.6151
R689 B.n384 B.n383 10.6151
R690 B.n383 B.n54 10.6151
R691 B.n377 B.n54 10.6151
R692 B.n377 B.n376 10.6151
R693 B.n376 B.n375 10.6151
R694 B.n375 B.n56 10.6151
R695 B.n369 B.n56 10.6151
R696 B.n367 B.n366 10.6151
R697 B.n366 B.n60 10.6151
R698 B.n360 B.n60 10.6151
R699 B.n360 B.n359 10.6151
R700 B.n359 B.n358 10.6151
R701 B.n358 B.n62 10.6151
R702 B.n352 B.n62 10.6151
R703 B.n352 B.n351 10.6151
R704 B.n351 B.n350 10.6151
R705 B.n346 B.n345 10.6151
R706 B.n345 B.n68 10.6151
R707 B.n340 B.n68 10.6151
R708 B.n340 B.n339 10.6151
R709 B.n339 B.n338 10.6151
R710 B.n338 B.n70 10.6151
R711 B.n332 B.n70 10.6151
R712 B.n332 B.n331 10.6151
R713 B.n331 B.n330 10.6151
R714 B.n330 B.n72 10.6151
R715 B.n324 B.n72 10.6151
R716 B.n215 B.n214 10.6151
R717 B.n216 B.n215 10.6151
R718 B.n216 B.n111 10.6151
R719 B.n226 B.n111 10.6151
R720 B.n227 B.n226 10.6151
R721 B.n228 B.n227 10.6151
R722 B.n228 B.n104 10.6151
R723 B.n239 B.n104 10.6151
R724 B.n240 B.n239 10.6151
R725 B.n241 B.n240 10.6151
R726 B.n241 B.n96 10.6151
R727 B.n251 B.n96 10.6151
R728 B.n252 B.n251 10.6151
R729 B.n253 B.n252 10.6151
R730 B.n253 B.n88 10.6151
R731 B.n263 B.n88 10.6151
R732 B.n264 B.n263 10.6151
R733 B.n265 B.n264 10.6151
R734 B.n265 B.n81 10.6151
R735 B.n276 B.n81 10.6151
R736 B.n277 B.n276 10.6151
R737 B.n279 B.n277 10.6151
R738 B.n279 B.n278 10.6151
R739 B.n278 B.n73 10.6151
R740 B.n290 B.n73 10.6151
R741 B.n291 B.n290 10.6151
R742 B.n292 B.n291 10.6151
R743 B.n293 B.n292 10.6151
R744 B.n295 B.n293 10.6151
R745 B.n296 B.n295 10.6151
R746 B.n297 B.n296 10.6151
R747 B.n298 B.n297 10.6151
R748 B.n300 B.n298 10.6151
R749 B.n301 B.n300 10.6151
R750 B.n302 B.n301 10.6151
R751 B.n303 B.n302 10.6151
R752 B.n305 B.n303 10.6151
R753 B.n306 B.n305 10.6151
R754 B.n307 B.n306 10.6151
R755 B.n308 B.n307 10.6151
R756 B.n310 B.n308 10.6151
R757 B.n311 B.n310 10.6151
R758 B.n312 B.n311 10.6151
R759 B.n313 B.n312 10.6151
R760 B.n315 B.n313 10.6151
R761 B.n316 B.n315 10.6151
R762 B.n317 B.n316 10.6151
R763 B.n318 B.n317 10.6151
R764 B.n320 B.n318 10.6151
R765 B.n321 B.n320 10.6151
R766 B.n322 B.n321 10.6151
R767 B.n323 B.n322 10.6151
R768 B.n209 B.n208 10.6151
R769 B.n208 B.n123 10.6151
R770 B.n203 B.n123 10.6151
R771 B.n203 B.n202 10.6151
R772 B.n202 B.n125 10.6151
R773 B.n197 B.n125 10.6151
R774 B.n197 B.n196 10.6151
R775 B.n196 B.n195 10.6151
R776 B.n195 B.n127 10.6151
R777 B.n189 B.n127 10.6151
R778 B.n189 B.n188 10.6151
R779 B.n186 B.n131 10.6151
R780 B.n180 B.n131 10.6151
R781 B.n180 B.n179 10.6151
R782 B.n179 B.n178 10.6151
R783 B.n178 B.n133 10.6151
R784 B.n172 B.n133 10.6151
R785 B.n172 B.n171 10.6151
R786 B.n171 B.n170 10.6151
R787 B.n170 B.n135 10.6151
R788 B.n164 B.n163 10.6151
R789 B.n163 B.n162 10.6151
R790 B.n162 B.n140 10.6151
R791 B.n156 B.n140 10.6151
R792 B.n156 B.n155 10.6151
R793 B.n155 B.n154 10.6151
R794 B.n154 B.n142 10.6151
R795 B.n148 B.n142 10.6151
R796 B.n148 B.n147 10.6151
R797 B.n147 B.n146 10.6151
R798 B.n146 B.n119 10.6151
R799 B.n210 B.n115 10.6151
R800 B.n220 B.n115 10.6151
R801 B.n221 B.n220 10.6151
R802 B.n222 B.n221 10.6151
R803 B.n222 B.n107 10.6151
R804 B.n233 B.n107 10.6151
R805 B.n234 B.n233 10.6151
R806 B.n235 B.n234 10.6151
R807 B.n235 B.n100 10.6151
R808 B.n245 B.n100 10.6151
R809 B.n246 B.n245 10.6151
R810 B.n247 B.n246 10.6151
R811 B.n247 B.n92 10.6151
R812 B.n257 B.n92 10.6151
R813 B.n258 B.n257 10.6151
R814 B.n259 B.n258 10.6151
R815 B.n259 B.n84 10.6151
R816 B.n270 B.n84 10.6151
R817 B.n271 B.n270 10.6151
R818 B.n272 B.n271 10.6151
R819 B.n272 B.n77 10.6151
R820 B.n283 B.n77 10.6151
R821 B.n284 B.n283 10.6151
R822 B.n285 B.n284 10.6151
R823 B.n285 B.n0 10.6151
R824 B.n441 B.n1 10.6151
R825 B.n441 B.n440 10.6151
R826 B.n440 B.n439 10.6151
R827 B.n439 B.n10 10.6151
R828 B.n433 B.n10 10.6151
R829 B.n433 B.n432 10.6151
R830 B.n432 B.n431 10.6151
R831 B.n431 B.n16 10.6151
R832 B.n425 B.n16 10.6151
R833 B.n425 B.n424 10.6151
R834 B.n424 B.n423 10.6151
R835 B.n423 B.n24 10.6151
R836 B.n417 B.n24 10.6151
R837 B.n417 B.n416 10.6151
R838 B.n416 B.n415 10.6151
R839 B.n415 B.n31 10.6151
R840 B.n409 B.n31 10.6151
R841 B.n409 B.n408 10.6151
R842 B.n408 B.n407 10.6151
R843 B.n407 B.n37 10.6151
R844 B.n401 B.n37 10.6151
R845 B.n401 B.n400 10.6151
R846 B.n400 B.n399 10.6151
R847 B.n399 B.n45 10.6151
R848 B.n393 B.n45 10.6151
R849 B.n369 B.n368 9.36635
R850 B.n346 B.n66 9.36635
R851 B.n188 B.n187 9.36635
R852 B.n164 B.n139 9.36635
R853 B.n447 B.n0 2.81026
R854 B.n447 B.n1 2.81026
R855 B.n368 B.n367 1.24928
R856 B.n350 B.n66 1.24928
R857 B.n187 B.n186 1.24928
R858 B.n139 B.n135 1.24928
R859 VN VN.t0 96.0459
R860 VN VN.t1 59.0308
R861 VDD2.n9 VDD2.n7 289.615
R862 VDD2.n2 VDD2.n0 289.615
R863 VDD2.n10 VDD2.n9 185
R864 VDD2.n3 VDD2.n2 185
R865 VDD2.t1 VDD2.n8 167.117
R866 VDD2.t0 VDD2.n1 167.117
R867 VDD2.n14 VDD2.n6 78.5625
R868 VDD2.n9 VDD2.t1 52.3082
R869 VDD2.n2 VDD2.t0 52.3082
R870 VDD2.n14 VDD2.n13 47.8944
R871 VDD2.n10 VDD2.n8 9.71174
R872 VDD2.n3 VDD2.n1 9.71174
R873 VDD2.n13 VDD2.n12 9.45567
R874 VDD2.n6 VDD2.n5 9.45567
R875 VDD2.n12 VDD2.n11 9.3005
R876 VDD2.n5 VDD2.n4 9.3005
R877 VDD2.n13 VDD2.n7 8.14595
R878 VDD2.n6 VDD2.n0 8.14595
R879 VDD2.n11 VDD2.n10 7.3702
R880 VDD2.n4 VDD2.n3 7.3702
R881 VDD2.n11 VDD2.n7 5.81868
R882 VDD2.n4 VDD2.n0 5.81868
R883 VDD2.n12 VDD2.n8 3.44771
R884 VDD2.n5 VDD2.n1 3.44771
R885 VDD2 VDD2.n14 0.720328
C0 VN VDD1 0.154498f
C1 VN VTAIL 0.986541f
C2 VDD2 VDD1 0.69041f
C3 VDD2 VTAIL 2.51958f
C4 VDD1 VP 0.868019f
C5 VTAIL VP 1.00068f
C6 VN VDD2 0.678869f
C7 VN VP 3.67764f
C8 VTAIL VDD1 2.46567f
C9 VDD2 VP 0.345259f
C10 VDD2 B 2.646674f
C11 VDD1 B 4.25786f
C12 VTAIL B 3.021838f
C13 VN B 7.76072f
C14 VP B 5.68861f
C15 VDD2.n0 B 0.025525f
C16 VDD2.n1 B 0.056518f
C17 VDD2.t0 B 0.042432f
C18 VDD2.n2 B 0.044197f
C19 VDD2.n3 B 0.014315f
C20 VDD2.n4 B 0.009441f
C21 VDD2.n5 B 0.12435f
C22 VDD2.n6 B 0.302313f
C23 VDD2.n7 B 0.025525f
C24 VDD2.n8 B 0.056518f
C25 VDD2.t1 B 0.042432f
C26 VDD2.n9 B 0.044197f
C27 VDD2.n10 B 0.014315f
C28 VDD2.n11 B 0.009441f
C29 VDD2.n12 B 0.12435f
C30 VDD2.n13 B 0.040106f
C31 VDD2.n14 B 1.40787f
C32 VN.t1 B 0.614259f
C33 VN.t0 B 1.08525f
C34 VDD1.n0 B 0.02488f
C35 VDD1.n1 B 0.055089f
C36 VDD1.t0 B 0.041358f
C37 VDD1.n2 B 0.043079f
C38 VDD1.n3 B 0.013953f
C39 VDD1.n4 B 0.009202f
C40 VDD1.n5 B 0.121204f
C41 VDD1.n6 B 0.040158f
C42 VDD1.n7 B 0.02488f
C43 VDD1.n8 B 0.055089f
C44 VDD1.t1 B 0.041358f
C45 VDD1.n9 B 0.043079f
C46 VDD1.n10 B 0.013953f
C47 VDD1.n11 B 0.009202f
C48 VDD1.n12 B 0.121204f
C49 VDD1.n13 B 0.322421f
C50 VTAIL.n0 B 0.031247f
C51 VTAIL.n1 B 0.069187f
C52 VTAIL.t1 B 0.051943f
C53 VTAIL.n2 B 0.054105f
C54 VTAIL.n3 B 0.017524f
C55 VTAIL.n4 B 0.011557f
C56 VTAIL.n5 B 0.152224f
C57 VTAIL.n6 B 0.034234f
C58 VTAIL.n7 B 0.877865f
C59 VTAIL.n8 B 0.031247f
C60 VTAIL.n9 B 0.069187f
C61 VTAIL.t2 B 0.051943f
C62 VTAIL.n10 B 0.054105f
C63 VTAIL.n11 B 0.017524f
C64 VTAIL.n12 B 0.011557f
C65 VTAIL.n13 B 0.152224f
C66 VTAIL.n14 B 0.034234f
C67 VTAIL.n15 B 0.919686f
C68 VTAIL.n16 B 0.031247f
C69 VTAIL.n17 B 0.069187f
C70 VTAIL.t0 B 0.051943f
C71 VTAIL.n18 B 0.054105f
C72 VTAIL.n19 B 0.017524f
C73 VTAIL.n20 B 0.011557f
C74 VTAIL.n21 B 0.152224f
C75 VTAIL.n22 B 0.034234f
C76 VTAIL.n23 B 0.736272f
C77 VTAIL.n24 B 0.031247f
C78 VTAIL.n25 B 0.069187f
C79 VTAIL.t3 B 0.051943f
C80 VTAIL.n26 B 0.054105f
C81 VTAIL.n27 B 0.017524f
C82 VTAIL.n28 B 0.011557f
C83 VTAIL.n29 B 0.152224f
C84 VTAIL.n30 B 0.034234f
C85 VTAIL.n31 B 0.653825f
C86 VP.t0 B 0.619058f
C87 VP.t1 B 1.09366f
C88 VP.n0 B 1.91049f
.ends

