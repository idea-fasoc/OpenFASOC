* NGSPICE file created from diff_pair_sample_0960.ext - technology: sky130A

.subckt diff_pair_sample_0960 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t3 w_n1414_n1846# sky130_fd_pr__pfet_01v8 ad=0.72435 pd=4.72 as=1.7121 ps=9.56 w=4.39 l=0.41
X1 VTAIL.t0 VN.t0 VDD2.t3 w_n1414_n1846# sky130_fd_pr__pfet_01v8 ad=1.7121 pd=9.56 as=0.72435 ps=4.72 w=4.39 l=0.41
X2 B.t11 B.t9 B.t10 w_n1414_n1846# sky130_fd_pr__pfet_01v8 ad=1.7121 pd=9.56 as=0 ps=0 w=4.39 l=0.41
X3 B.t8 B.t6 B.t7 w_n1414_n1846# sky130_fd_pr__pfet_01v8 ad=1.7121 pd=9.56 as=0 ps=0 w=4.39 l=0.41
X4 B.t5 B.t3 B.t4 w_n1414_n1846# sky130_fd_pr__pfet_01v8 ad=1.7121 pd=9.56 as=0 ps=0 w=4.39 l=0.41
X5 VDD2.t2 VN.t1 VTAIL.t1 w_n1414_n1846# sky130_fd_pr__pfet_01v8 ad=0.72435 pd=4.72 as=1.7121 ps=9.56 w=4.39 l=0.41
X6 VTAIL.t5 VP.t1 VDD1.t2 w_n1414_n1846# sky130_fd_pr__pfet_01v8 ad=1.7121 pd=9.56 as=0.72435 ps=4.72 w=4.39 l=0.41
X7 VTAIL.t2 VN.t2 VDD2.t1 w_n1414_n1846# sky130_fd_pr__pfet_01v8 ad=1.7121 pd=9.56 as=0.72435 ps=4.72 w=4.39 l=0.41
X8 VDD2.t0 VN.t3 VTAIL.t7 w_n1414_n1846# sky130_fd_pr__pfet_01v8 ad=0.72435 pd=4.72 as=1.7121 ps=9.56 w=4.39 l=0.41
X9 B.t2 B.t0 B.t1 w_n1414_n1846# sky130_fd_pr__pfet_01v8 ad=1.7121 pd=9.56 as=0 ps=0 w=4.39 l=0.41
X10 VTAIL.t4 VP.t2 VDD1.t1 w_n1414_n1846# sky130_fd_pr__pfet_01v8 ad=1.7121 pd=9.56 as=0.72435 ps=4.72 w=4.39 l=0.41
X11 VDD1.t0 VP.t3 VTAIL.t6 w_n1414_n1846# sky130_fd_pr__pfet_01v8 ad=0.72435 pd=4.72 as=1.7121 ps=9.56 w=4.39 l=0.41
R0 VP.n0 VP.t2 375.428
R1 VP.n0 VP.t3 375.404
R2 VP.n2 VP.t1 354.447
R3 VP.n3 VP.t0 354.447
R4 VP.n4 VP.n3 161.3
R5 VP.n2 VP.n1 161.3
R6 VP.n1 VP.n0 103.948
R7 VP.n3 VP.n2 48.2005
R8 VP.n4 VP.n1 0.189894
R9 VP VP.n4 0.0516364
R10 VTAIL.n5 VTAIL.t4 102.797
R11 VTAIL.n4 VTAIL.t1 102.797
R12 VTAIL.n3 VTAIL.t2 102.797
R13 VTAIL.n7 VTAIL.t7 102.796
R14 VTAIL.n0 VTAIL.t0 102.796
R15 VTAIL.n1 VTAIL.t3 102.796
R16 VTAIL.n2 VTAIL.t5 102.796
R17 VTAIL.n6 VTAIL.t6 102.796
R18 VTAIL.n7 VTAIL.n6 16.7893
R19 VTAIL.n3 VTAIL.n2 16.7893
R20 VTAIL.n4 VTAIL.n3 0.638431
R21 VTAIL.n6 VTAIL.n5 0.638431
R22 VTAIL.n2 VTAIL.n1 0.638431
R23 VTAIL.n5 VTAIL.n4 0.470328
R24 VTAIL.n1 VTAIL.n0 0.470328
R25 VTAIL VTAIL.n0 0.377655
R26 VTAIL VTAIL.n7 0.261276
R27 VDD1 VDD1.n1 142.01
R28 VDD1 VDD1.n0 112.129
R29 VDD1.n0 VDD1.t1 7.40483
R30 VDD1.n0 VDD1.t0 7.40483
R31 VDD1.n1 VDD1.t2 7.40483
R32 VDD1.n1 VDD1.t3 7.40483
R33 VN.n0 VN.t0 375.428
R34 VN.n1 VN.t1 375.428
R35 VN.n0 VN.t3 375.404
R36 VN.n1 VN.t2 375.404
R37 VN VN.n1 104.329
R38 VN VN.n0 70.265
R39 VDD2.n2 VDD2.n0 141.484
R40 VDD2.n2 VDD2.n1 112.072
R41 VDD2.n1 VDD2.t1 7.40483
R42 VDD2.n1 VDD2.t2 7.40483
R43 VDD2.n0 VDD2.t3 7.40483
R44 VDD2.n0 VDD2.t0 7.40483
R45 VDD2 VDD2.n2 0.0586897
R46 B.n180 B.n53 585
R47 B.n179 B.n178 585
R48 B.n177 B.n54 585
R49 B.n176 B.n175 585
R50 B.n174 B.n55 585
R51 B.n173 B.n172 585
R52 B.n171 B.n56 585
R53 B.n170 B.n169 585
R54 B.n168 B.n57 585
R55 B.n167 B.n166 585
R56 B.n165 B.n58 585
R57 B.n164 B.n163 585
R58 B.n162 B.n59 585
R59 B.n161 B.n160 585
R60 B.n159 B.n60 585
R61 B.n158 B.n157 585
R62 B.n156 B.n61 585
R63 B.n155 B.n154 585
R64 B.n153 B.n62 585
R65 B.n151 B.n150 585
R66 B.n149 B.n65 585
R67 B.n148 B.n147 585
R68 B.n146 B.n66 585
R69 B.n145 B.n144 585
R70 B.n143 B.n67 585
R71 B.n142 B.n141 585
R72 B.n140 B.n68 585
R73 B.n139 B.n138 585
R74 B.n137 B.n69 585
R75 B.n136 B.n135 585
R76 B.n131 B.n70 585
R77 B.n130 B.n129 585
R78 B.n128 B.n71 585
R79 B.n127 B.n126 585
R80 B.n125 B.n72 585
R81 B.n124 B.n123 585
R82 B.n122 B.n73 585
R83 B.n121 B.n120 585
R84 B.n119 B.n74 585
R85 B.n118 B.n117 585
R86 B.n116 B.n75 585
R87 B.n115 B.n114 585
R88 B.n113 B.n76 585
R89 B.n112 B.n111 585
R90 B.n110 B.n77 585
R91 B.n109 B.n108 585
R92 B.n107 B.n78 585
R93 B.n106 B.n105 585
R94 B.n182 B.n181 585
R95 B.n183 B.n52 585
R96 B.n185 B.n184 585
R97 B.n186 B.n51 585
R98 B.n188 B.n187 585
R99 B.n189 B.n50 585
R100 B.n191 B.n190 585
R101 B.n192 B.n49 585
R102 B.n194 B.n193 585
R103 B.n195 B.n48 585
R104 B.n197 B.n196 585
R105 B.n198 B.n47 585
R106 B.n200 B.n199 585
R107 B.n201 B.n46 585
R108 B.n203 B.n202 585
R109 B.n204 B.n45 585
R110 B.n206 B.n205 585
R111 B.n207 B.n44 585
R112 B.n209 B.n208 585
R113 B.n210 B.n43 585
R114 B.n212 B.n211 585
R115 B.n213 B.n42 585
R116 B.n215 B.n214 585
R117 B.n216 B.n41 585
R118 B.n218 B.n217 585
R119 B.n219 B.n40 585
R120 B.n221 B.n220 585
R121 B.n222 B.n39 585
R122 B.n224 B.n223 585
R123 B.n225 B.n38 585
R124 B.n298 B.n9 585
R125 B.n297 B.n296 585
R126 B.n295 B.n10 585
R127 B.n294 B.n293 585
R128 B.n292 B.n11 585
R129 B.n291 B.n290 585
R130 B.n289 B.n12 585
R131 B.n288 B.n287 585
R132 B.n286 B.n13 585
R133 B.n285 B.n284 585
R134 B.n283 B.n14 585
R135 B.n282 B.n281 585
R136 B.n280 B.n15 585
R137 B.n279 B.n278 585
R138 B.n277 B.n16 585
R139 B.n276 B.n275 585
R140 B.n274 B.n17 585
R141 B.n273 B.n272 585
R142 B.n271 B.n18 585
R143 B.n270 B.n269 585
R144 B.n268 B.n19 585
R145 B.n267 B.n266 585
R146 B.n265 B.n23 585
R147 B.n264 B.n263 585
R148 B.n262 B.n24 585
R149 B.n261 B.n260 585
R150 B.n259 B.n25 585
R151 B.n258 B.n257 585
R152 B.n256 B.n26 585
R153 B.n254 B.n253 585
R154 B.n252 B.n29 585
R155 B.n251 B.n250 585
R156 B.n249 B.n30 585
R157 B.n248 B.n247 585
R158 B.n246 B.n31 585
R159 B.n245 B.n244 585
R160 B.n243 B.n32 585
R161 B.n242 B.n241 585
R162 B.n240 B.n33 585
R163 B.n239 B.n238 585
R164 B.n237 B.n34 585
R165 B.n236 B.n235 585
R166 B.n234 B.n35 585
R167 B.n233 B.n232 585
R168 B.n231 B.n36 585
R169 B.n230 B.n229 585
R170 B.n228 B.n37 585
R171 B.n227 B.n226 585
R172 B.n300 B.n299 585
R173 B.n301 B.n8 585
R174 B.n303 B.n302 585
R175 B.n304 B.n7 585
R176 B.n306 B.n305 585
R177 B.n307 B.n6 585
R178 B.n309 B.n308 585
R179 B.n310 B.n5 585
R180 B.n312 B.n311 585
R181 B.n313 B.n4 585
R182 B.n315 B.n314 585
R183 B.n316 B.n3 585
R184 B.n318 B.n317 585
R185 B.n319 B.n0 585
R186 B.n2 B.n1 585
R187 B.n86 B.n85 585
R188 B.n88 B.n87 585
R189 B.n89 B.n84 585
R190 B.n91 B.n90 585
R191 B.n92 B.n83 585
R192 B.n94 B.n93 585
R193 B.n95 B.n82 585
R194 B.n97 B.n96 585
R195 B.n98 B.n81 585
R196 B.n100 B.n99 585
R197 B.n101 B.n80 585
R198 B.n103 B.n102 585
R199 B.n104 B.n79 585
R200 B.n105 B.n104 526.135
R201 B.n181 B.n180 526.135
R202 B.n227 B.n38 526.135
R203 B.n300 B.n9 526.135
R204 B.n132 B.t0 467.099
R205 B.n63 B.t3 467.099
R206 B.n27 B.t9 467.099
R207 B.n20 B.t6 467.099
R208 B.n321 B.n320 256.663
R209 B.n320 B.n319 235.042
R210 B.n320 B.n2 235.042
R211 B.n105 B.n78 163.367
R212 B.n109 B.n78 163.367
R213 B.n110 B.n109 163.367
R214 B.n111 B.n110 163.367
R215 B.n111 B.n76 163.367
R216 B.n115 B.n76 163.367
R217 B.n116 B.n115 163.367
R218 B.n117 B.n116 163.367
R219 B.n117 B.n74 163.367
R220 B.n121 B.n74 163.367
R221 B.n122 B.n121 163.367
R222 B.n123 B.n122 163.367
R223 B.n123 B.n72 163.367
R224 B.n127 B.n72 163.367
R225 B.n128 B.n127 163.367
R226 B.n129 B.n128 163.367
R227 B.n129 B.n70 163.367
R228 B.n136 B.n70 163.367
R229 B.n137 B.n136 163.367
R230 B.n138 B.n137 163.367
R231 B.n138 B.n68 163.367
R232 B.n142 B.n68 163.367
R233 B.n143 B.n142 163.367
R234 B.n144 B.n143 163.367
R235 B.n144 B.n66 163.367
R236 B.n148 B.n66 163.367
R237 B.n149 B.n148 163.367
R238 B.n150 B.n149 163.367
R239 B.n150 B.n62 163.367
R240 B.n155 B.n62 163.367
R241 B.n156 B.n155 163.367
R242 B.n157 B.n156 163.367
R243 B.n157 B.n60 163.367
R244 B.n161 B.n60 163.367
R245 B.n162 B.n161 163.367
R246 B.n163 B.n162 163.367
R247 B.n163 B.n58 163.367
R248 B.n167 B.n58 163.367
R249 B.n168 B.n167 163.367
R250 B.n169 B.n168 163.367
R251 B.n169 B.n56 163.367
R252 B.n173 B.n56 163.367
R253 B.n174 B.n173 163.367
R254 B.n175 B.n174 163.367
R255 B.n175 B.n54 163.367
R256 B.n179 B.n54 163.367
R257 B.n180 B.n179 163.367
R258 B.n223 B.n38 163.367
R259 B.n223 B.n222 163.367
R260 B.n222 B.n221 163.367
R261 B.n221 B.n40 163.367
R262 B.n217 B.n40 163.367
R263 B.n217 B.n216 163.367
R264 B.n216 B.n215 163.367
R265 B.n215 B.n42 163.367
R266 B.n211 B.n42 163.367
R267 B.n211 B.n210 163.367
R268 B.n210 B.n209 163.367
R269 B.n209 B.n44 163.367
R270 B.n205 B.n44 163.367
R271 B.n205 B.n204 163.367
R272 B.n204 B.n203 163.367
R273 B.n203 B.n46 163.367
R274 B.n199 B.n46 163.367
R275 B.n199 B.n198 163.367
R276 B.n198 B.n197 163.367
R277 B.n197 B.n48 163.367
R278 B.n193 B.n48 163.367
R279 B.n193 B.n192 163.367
R280 B.n192 B.n191 163.367
R281 B.n191 B.n50 163.367
R282 B.n187 B.n50 163.367
R283 B.n187 B.n186 163.367
R284 B.n186 B.n185 163.367
R285 B.n185 B.n52 163.367
R286 B.n181 B.n52 163.367
R287 B.n296 B.n9 163.367
R288 B.n296 B.n295 163.367
R289 B.n295 B.n294 163.367
R290 B.n294 B.n11 163.367
R291 B.n290 B.n11 163.367
R292 B.n290 B.n289 163.367
R293 B.n289 B.n288 163.367
R294 B.n288 B.n13 163.367
R295 B.n284 B.n13 163.367
R296 B.n284 B.n283 163.367
R297 B.n283 B.n282 163.367
R298 B.n282 B.n15 163.367
R299 B.n278 B.n15 163.367
R300 B.n278 B.n277 163.367
R301 B.n277 B.n276 163.367
R302 B.n276 B.n17 163.367
R303 B.n272 B.n17 163.367
R304 B.n272 B.n271 163.367
R305 B.n271 B.n270 163.367
R306 B.n270 B.n19 163.367
R307 B.n266 B.n19 163.367
R308 B.n266 B.n265 163.367
R309 B.n265 B.n264 163.367
R310 B.n264 B.n24 163.367
R311 B.n260 B.n24 163.367
R312 B.n260 B.n259 163.367
R313 B.n259 B.n258 163.367
R314 B.n258 B.n26 163.367
R315 B.n253 B.n26 163.367
R316 B.n253 B.n252 163.367
R317 B.n252 B.n251 163.367
R318 B.n251 B.n30 163.367
R319 B.n247 B.n30 163.367
R320 B.n247 B.n246 163.367
R321 B.n246 B.n245 163.367
R322 B.n245 B.n32 163.367
R323 B.n241 B.n32 163.367
R324 B.n241 B.n240 163.367
R325 B.n240 B.n239 163.367
R326 B.n239 B.n34 163.367
R327 B.n235 B.n34 163.367
R328 B.n235 B.n234 163.367
R329 B.n234 B.n233 163.367
R330 B.n233 B.n36 163.367
R331 B.n229 B.n36 163.367
R332 B.n229 B.n228 163.367
R333 B.n228 B.n227 163.367
R334 B.n301 B.n300 163.367
R335 B.n302 B.n301 163.367
R336 B.n302 B.n7 163.367
R337 B.n306 B.n7 163.367
R338 B.n307 B.n306 163.367
R339 B.n308 B.n307 163.367
R340 B.n308 B.n5 163.367
R341 B.n312 B.n5 163.367
R342 B.n313 B.n312 163.367
R343 B.n314 B.n313 163.367
R344 B.n314 B.n3 163.367
R345 B.n318 B.n3 163.367
R346 B.n319 B.n318 163.367
R347 B.n86 B.n2 163.367
R348 B.n87 B.n86 163.367
R349 B.n87 B.n84 163.367
R350 B.n91 B.n84 163.367
R351 B.n92 B.n91 163.367
R352 B.n93 B.n92 163.367
R353 B.n93 B.n82 163.367
R354 B.n97 B.n82 163.367
R355 B.n98 B.n97 163.367
R356 B.n99 B.n98 163.367
R357 B.n99 B.n80 163.367
R358 B.n103 B.n80 163.367
R359 B.n104 B.n103 163.367
R360 B.n63 B.t4 138.893
R361 B.n27 B.t11 138.893
R362 B.n132 B.t1 138.888
R363 B.n20 B.t8 138.888
R364 B.n64 B.t5 124.54
R365 B.n28 B.t10 124.54
R366 B.n133 B.t2 124.537
R367 B.n21 B.t7 124.537
R368 B.n134 B.n133 59.5399
R369 B.n152 B.n64 59.5399
R370 B.n255 B.n28 59.5399
R371 B.n22 B.n21 59.5399
R372 B.n299 B.n298 34.1859
R373 B.n226 B.n225 34.1859
R374 B.n182 B.n53 34.1859
R375 B.n106 B.n79 34.1859
R376 B B.n321 18.0485
R377 B.n133 B.n132 14.352
R378 B.n64 B.n63 14.352
R379 B.n28 B.n27 14.352
R380 B.n21 B.n20 14.352
R381 B.n299 B.n8 10.6151
R382 B.n303 B.n8 10.6151
R383 B.n304 B.n303 10.6151
R384 B.n305 B.n304 10.6151
R385 B.n305 B.n6 10.6151
R386 B.n309 B.n6 10.6151
R387 B.n310 B.n309 10.6151
R388 B.n311 B.n310 10.6151
R389 B.n311 B.n4 10.6151
R390 B.n315 B.n4 10.6151
R391 B.n316 B.n315 10.6151
R392 B.n317 B.n316 10.6151
R393 B.n317 B.n0 10.6151
R394 B.n298 B.n297 10.6151
R395 B.n297 B.n10 10.6151
R396 B.n293 B.n10 10.6151
R397 B.n293 B.n292 10.6151
R398 B.n292 B.n291 10.6151
R399 B.n291 B.n12 10.6151
R400 B.n287 B.n12 10.6151
R401 B.n287 B.n286 10.6151
R402 B.n286 B.n285 10.6151
R403 B.n285 B.n14 10.6151
R404 B.n281 B.n14 10.6151
R405 B.n281 B.n280 10.6151
R406 B.n280 B.n279 10.6151
R407 B.n279 B.n16 10.6151
R408 B.n275 B.n16 10.6151
R409 B.n275 B.n274 10.6151
R410 B.n274 B.n273 10.6151
R411 B.n273 B.n18 10.6151
R412 B.n269 B.n268 10.6151
R413 B.n268 B.n267 10.6151
R414 B.n267 B.n23 10.6151
R415 B.n263 B.n23 10.6151
R416 B.n263 B.n262 10.6151
R417 B.n262 B.n261 10.6151
R418 B.n261 B.n25 10.6151
R419 B.n257 B.n25 10.6151
R420 B.n257 B.n256 10.6151
R421 B.n254 B.n29 10.6151
R422 B.n250 B.n29 10.6151
R423 B.n250 B.n249 10.6151
R424 B.n249 B.n248 10.6151
R425 B.n248 B.n31 10.6151
R426 B.n244 B.n31 10.6151
R427 B.n244 B.n243 10.6151
R428 B.n243 B.n242 10.6151
R429 B.n242 B.n33 10.6151
R430 B.n238 B.n33 10.6151
R431 B.n238 B.n237 10.6151
R432 B.n237 B.n236 10.6151
R433 B.n236 B.n35 10.6151
R434 B.n232 B.n35 10.6151
R435 B.n232 B.n231 10.6151
R436 B.n231 B.n230 10.6151
R437 B.n230 B.n37 10.6151
R438 B.n226 B.n37 10.6151
R439 B.n225 B.n224 10.6151
R440 B.n224 B.n39 10.6151
R441 B.n220 B.n39 10.6151
R442 B.n220 B.n219 10.6151
R443 B.n219 B.n218 10.6151
R444 B.n218 B.n41 10.6151
R445 B.n214 B.n41 10.6151
R446 B.n214 B.n213 10.6151
R447 B.n213 B.n212 10.6151
R448 B.n212 B.n43 10.6151
R449 B.n208 B.n43 10.6151
R450 B.n208 B.n207 10.6151
R451 B.n207 B.n206 10.6151
R452 B.n206 B.n45 10.6151
R453 B.n202 B.n45 10.6151
R454 B.n202 B.n201 10.6151
R455 B.n201 B.n200 10.6151
R456 B.n200 B.n47 10.6151
R457 B.n196 B.n47 10.6151
R458 B.n196 B.n195 10.6151
R459 B.n195 B.n194 10.6151
R460 B.n194 B.n49 10.6151
R461 B.n190 B.n49 10.6151
R462 B.n190 B.n189 10.6151
R463 B.n189 B.n188 10.6151
R464 B.n188 B.n51 10.6151
R465 B.n184 B.n51 10.6151
R466 B.n184 B.n183 10.6151
R467 B.n183 B.n182 10.6151
R468 B.n85 B.n1 10.6151
R469 B.n88 B.n85 10.6151
R470 B.n89 B.n88 10.6151
R471 B.n90 B.n89 10.6151
R472 B.n90 B.n83 10.6151
R473 B.n94 B.n83 10.6151
R474 B.n95 B.n94 10.6151
R475 B.n96 B.n95 10.6151
R476 B.n96 B.n81 10.6151
R477 B.n100 B.n81 10.6151
R478 B.n101 B.n100 10.6151
R479 B.n102 B.n101 10.6151
R480 B.n102 B.n79 10.6151
R481 B.n107 B.n106 10.6151
R482 B.n108 B.n107 10.6151
R483 B.n108 B.n77 10.6151
R484 B.n112 B.n77 10.6151
R485 B.n113 B.n112 10.6151
R486 B.n114 B.n113 10.6151
R487 B.n114 B.n75 10.6151
R488 B.n118 B.n75 10.6151
R489 B.n119 B.n118 10.6151
R490 B.n120 B.n119 10.6151
R491 B.n120 B.n73 10.6151
R492 B.n124 B.n73 10.6151
R493 B.n125 B.n124 10.6151
R494 B.n126 B.n125 10.6151
R495 B.n126 B.n71 10.6151
R496 B.n130 B.n71 10.6151
R497 B.n131 B.n130 10.6151
R498 B.n135 B.n131 10.6151
R499 B.n139 B.n69 10.6151
R500 B.n140 B.n139 10.6151
R501 B.n141 B.n140 10.6151
R502 B.n141 B.n67 10.6151
R503 B.n145 B.n67 10.6151
R504 B.n146 B.n145 10.6151
R505 B.n147 B.n146 10.6151
R506 B.n147 B.n65 10.6151
R507 B.n151 B.n65 10.6151
R508 B.n154 B.n153 10.6151
R509 B.n154 B.n61 10.6151
R510 B.n158 B.n61 10.6151
R511 B.n159 B.n158 10.6151
R512 B.n160 B.n159 10.6151
R513 B.n160 B.n59 10.6151
R514 B.n164 B.n59 10.6151
R515 B.n165 B.n164 10.6151
R516 B.n166 B.n165 10.6151
R517 B.n166 B.n57 10.6151
R518 B.n170 B.n57 10.6151
R519 B.n171 B.n170 10.6151
R520 B.n172 B.n171 10.6151
R521 B.n172 B.n55 10.6151
R522 B.n176 B.n55 10.6151
R523 B.n177 B.n176 10.6151
R524 B.n178 B.n177 10.6151
R525 B.n178 B.n53 10.6151
R526 B.n22 B.n18 9.36635
R527 B.n255 B.n254 9.36635
R528 B.n135 B.n134 9.36635
R529 B.n153 B.n152 9.36635
R530 B.n321 B.n0 8.11757
R531 B.n321 B.n1 8.11757
R532 B.n269 B.n22 1.24928
R533 B.n256 B.n255 1.24928
R534 B.n134 B.n69 1.24928
R535 B.n152 B.n151 1.24928
C0 VDD1 VP 1.17039f
C1 VN w_n1414_n1846# 1.84533f
C2 VDD2 w_n1414_n1846# 0.802243f
C3 VTAIL B 1.62844f
C4 VDD2 VN 1.06265f
C5 VTAIL VP 0.973867f
C6 VDD1 w_n1414_n1846# 0.793645f
C7 VDD1 VN 0.151173f
C8 VDD2 VDD1 0.5039f
C9 VP B 0.881259f
C10 VTAIL w_n1414_n1846# 2.1982f
C11 VTAIL VN 0.959761f
C12 VDD2 VTAIL 3.92439f
C13 w_n1414_n1846# B 4.41371f
C14 VN B 0.59912f
C15 VDD2 B 0.686422f
C16 VP w_n1414_n1846# 2.0212f
C17 VTAIL VDD1 3.88487f
C18 VP VN 3.21226f
C19 VDD2 VP 0.259408f
C20 VDD1 B 0.668893f
C21 VDD2 VSUBS 0.432426f
C22 VDD1 VSUBS 2.964145f
C23 VTAIL VSUBS 0.388424f
C24 VN VSUBS 3.07725f
C25 VP VSUBS 0.77824f
C26 B VSUBS 1.655256f
C27 w_n1414_n1846# VSUBS 32.799103f
C28 B.n0 VSUBS 0.006466f
C29 B.n1 VSUBS 0.006466f
C30 B.n2 VSUBS 0.009563f
C31 B.n3 VSUBS 0.007329f
C32 B.n4 VSUBS 0.007329f
C33 B.n5 VSUBS 0.007329f
C34 B.n6 VSUBS 0.007329f
C35 B.n7 VSUBS 0.007329f
C36 B.n8 VSUBS 0.007329f
C37 B.n9 VSUBS 0.018149f
C38 B.n10 VSUBS 0.007329f
C39 B.n11 VSUBS 0.007329f
C40 B.n12 VSUBS 0.007329f
C41 B.n13 VSUBS 0.007329f
C42 B.n14 VSUBS 0.007329f
C43 B.n15 VSUBS 0.007329f
C44 B.n16 VSUBS 0.007329f
C45 B.n17 VSUBS 0.007329f
C46 B.n18 VSUBS 0.006898f
C47 B.n19 VSUBS 0.007329f
C48 B.t7 VSUBS 0.123637f
C49 B.t8 VSUBS 0.129107f
C50 B.t6 VSUBS 0.080347f
C51 B.n20 VSUBS 0.073896f
C52 B.n21 VSUBS 0.063396f
C53 B.n22 VSUBS 0.01698f
C54 B.n23 VSUBS 0.007329f
C55 B.n24 VSUBS 0.007329f
C56 B.n25 VSUBS 0.007329f
C57 B.n26 VSUBS 0.007329f
C58 B.t10 VSUBS 0.123637f
C59 B.t11 VSUBS 0.129107f
C60 B.t9 VSUBS 0.080347f
C61 B.n27 VSUBS 0.073896f
C62 B.n28 VSUBS 0.063396f
C63 B.n29 VSUBS 0.007329f
C64 B.n30 VSUBS 0.007329f
C65 B.n31 VSUBS 0.007329f
C66 B.n32 VSUBS 0.007329f
C67 B.n33 VSUBS 0.007329f
C68 B.n34 VSUBS 0.007329f
C69 B.n35 VSUBS 0.007329f
C70 B.n36 VSUBS 0.007329f
C71 B.n37 VSUBS 0.007329f
C72 B.n38 VSUBS 0.017201f
C73 B.n39 VSUBS 0.007329f
C74 B.n40 VSUBS 0.007329f
C75 B.n41 VSUBS 0.007329f
C76 B.n42 VSUBS 0.007329f
C77 B.n43 VSUBS 0.007329f
C78 B.n44 VSUBS 0.007329f
C79 B.n45 VSUBS 0.007329f
C80 B.n46 VSUBS 0.007329f
C81 B.n47 VSUBS 0.007329f
C82 B.n48 VSUBS 0.007329f
C83 B.n49 VSUBS 0.007329f
C84 B.n50 VSUBS 0.007329f
C85 B.n51 VSUBS 0.007329f
C86 B.n52 VSUBS 0.007329f
C87 B.n53 VSUBS 0.017322f
C88 B.n54 VSUBS 0.007329f
C89 B.n55 VSUBS 0.007329f
C90 B.n56 VSUBS 0.007329f
C91 B.n57 VSUBS 0.007329f
C92 B.n58 VSUBS 0.007329f
C93 B.n59 VSUBS 0.007329f
C94 B.n60 VSUBS 0.007329f
C95 B.n61 VSUBS 0.007329f
C96 B.n62 VSUBS 0.007329f
C97 B.t5 VSUBS 0.123637f
C98 B.t4 VSUBS 0.129107f
C99 B.t3 VSUBS 0.080347f
C100 B.n63 VSUBS 0.073896f
C101 B.n64 VSUBS 0.063396f
C102 B.n65 VSUBS 0.007329f
C103 B.n66 VSUBS 0.007329f
C104 B.n67 VSUBS 0.007329f
C105 B.n68 VSUBS 0.007329f
C106 B.n69 VSUBS 0.004095f
C107 B.n70 VSUBS 0.007329f
C108 B.n71 VSUBS 0.007329f
C109 B.n72 VSUBS 0.007329f
C110 B.n73 VSUBS 0.007329f
C111 B.n74 VSUBS 0.007329f
C112 B.n75 VSUBS 0.007329f
C113 B.n76 VSUBS 0.007329f
C114 B.n77 VSUBS 0.007329f
C115 B.n78 VSUBS 0.007329f
C116 B.n79 VSUBS 0.017201f
C117 B.n80 VSUBS 0.007329f
C118 B.n81 VSUBS 0.007329f
C119 B.n82 VSUBS 0.007329f
C120 B.n83 VSUBS 0.007329f
C121 B.n84 VSUBS 0.007329f
C122 B.n85 VSUBS 0.007329f
C123 B.n86 VSUBS 0.007329f
C124 B.n87 VSUBS 0.007329f
C125 B.n88 VSUBS 0.007329f
C126 B.n89 VSUBS 0.007329f
C127 B.n90 VSUBS 0.007329f
C128 B.n91 VSUBS 0.007329f
C129 B.n92 VSUBS 0.007329f
C130 B.n93 VSUBS 0.007329f
C131 B.n94 VSUBS 0.007329f
C132 B.n95 VSUBS 0.007329f
C133 B.n96 VSUBS 0.007329f
C134 B.n97 VSUBS 0.007329f
C135 B.n98 VSUBS 0.007329f
C136 B.n99 VSUBS 0.007329f
C137 B.n100 VSUBS 0.007329f
C138 B.n101 VSUBS 0.007329f
C139 B.n102 VSUBS 0.007329f
C140 B.n103 VSUBS 0.007329f
C141 B.n104 VSUBS 0.017201f
C142 B.n105 VSUBS 0.018149f
C143 B.n106 VSUBS 0.018149f
C144 B.n107 VSUBS 0.007329f
C145 B.n108 VSUBS 0.007329f
C146 B.n109 VSUBS 0.007329f
C147 B.n110 VSUBS 0.007329f
C148 B.n111 VSUBS 0.007329f
C149 B.n112 VSUBS 0.007329f
C150 B.n113 VSUBS 0.007329f
C151 B.n114 VSUBS 0.007329f
C152 B.n115 VSUBS 0.007329f
C153 B.n116 VSUBS 0.007329f
C154 B.n117 VSUBS 0.007329f
C155 B.n118 VSUBS 0.007329f
C156 B.n119 VSUBS 0.007329f
C157 B.n120 VSUBS 0.007329f
C158 B.n121 VSUBS 0.007329f
C159 B.n122 VSUBS 0.007329f
C160 B.n123 VSUBS 0.007329f
C161 B.n124 VSUBS 0.007329f
C162 B.n125 VSUBS 0.007329f
C163 B.n126 VSUBS 0.007329f
C164 B.n127 VSUBS 0.007329f
C165 B.n128 VSUBS 0.007329f
C166 B.n129 VSUBS 0.007329f
C167 B.n130 VSUBS 0.007329f
C168 B.n131 VSUBS 0.007329f
C169 B.t2 VSUBS 0.123637f
C170 B.t1 VSUBS 0.129107f
C171 B.t0 VSUBS 0.080347f
C172 B.n132 VSUBS 0.073896f
C173 B.n133 VSUBS 0.063396f
C174 B.n134 VSUBS 0.01698f
C175 B.n135 VSUBS 0.006898f
C176 B.n136 VSUBS 0.007329f
C177 B.n137 VSUBS 0.007329f
C178 B.n138 VSUBS 0.007329f
C179 B.n139 VSUBS 0.007329f
C180 B.n140 VSUBS 0.007329f
C181 B.n141 VSUBS 0.007329f
C182 B.n142 VSUBS 0.007329f
C183 B.n143 VSUBS 0.007329f
C184 B.n144 VSUBS 0.007329f
C185 B.n145 VSUBS 0.007329f
C186 B.n146 VSUBS 0.007329f
C187 B.n147 VSUBS 0.007329f
C188 B.n148 VSUBS 0.007329f
C189 B.n149 VSUBS 0.007329f
C190 B.n150 VSUBS 0.007329f
C191 B.n151 VSUBS 0.004095f
C192 B.n152 VSUBS 0.01698f
C193 B.n153 VSUBS 0.006898f
C194 B.n154 VSUBS 0.007329f
C195 B.n155 VSUBS 0.007329f
C196 B.n156 VSUBS 0.007329f
C197 B.n157 VSUBS 0.007329f
C198 B.n158 VSUBS 0.007329f
C199 B.n159 VSUBS 0.007329f
C200 B.n160 VSUBS 0.007329f
C201 B.n161 VSUBS 0.007329f
C202 B.n162 VSUBS 0.007329f
C203 B.n163 VSUBS 0.007329f
C204 B.n164 VSUBS 0.007329f
C205 B.n165 VSUBS 0.007329f
C206 B.n166 VSUBS 0.007329f
C207 B.n167 VSUBS 0.007329f
C208 B.n168 VSUBS 0.007329f
C209 B.n169 VSUBS 0.007329f
C210 B.n170 VSUBS 0.007329f
C211 B.n171 VSUBS 0.007329f
C212 B.n172 VSUBS 0.007329f
C213 B.n173 VSUBS 0.007329f
C214 B.n174 VSUBS 0.007329f
C215 B.n175 VSUBS 0.007329f
C216 B.n176 VSUBS 0.007329f
C217 B.n177 VSUBS 0.007329f
C218 B.n178 VSUBS 0.007329f
C219 B.n179 VSUBS 0.007329f
C220 B.n180 VSUBS 0.018149f
C221 B.n181 VSUBS 0.017201f
C222 B.n182 VSUBS 0.018028f
C223 B.n183 VSUBS 0.007329f
C224 B.n184 VSUBS 0.007329f
C225 B.n185 VSUBS 0.007329f
C226 B.n186 VSUBS 0.007329f
C227 B.n187 VSUBS 0.007329f
C228 B.n188 VSUBS 0.007329f
C229 B.n189 VSUBS 0.007329f
C230 B.n190 VSUBS 0.007329f
C231 B.n191 VSUBS 0.007329f
C232 B.n192 VSUBS 0.007329f
C233 B.n193 VSUBS 0.007329f
C234 B.n194 VSUBS 0.007329f
C235 B.n195 VSUBS 0.007329f
C236 B.n196 VSUBS 0.007329f
C237 B.n197 VSUBS 0.007329f
C238 B.n198 VSUBS 0.007329f
C239 B.n199 VSUBS 0.007329f
C240 B.n200 VSUBS 0.007329f
C241 B.n201 VSUBS 0.007329f
C242 B.n202 VSUBS 0.007329f
C243 B.n203 VSUBS 0.007329f
C244 B.n204 VSUBS 0.007329f
C245 B.n205 VSUBS 0.007329f
C246 B.n206 VSUBS 0.007329f
C247 B.n207 VSUBS 0.007329f
C248 B.n208 VSUBS 0.007329f
C249 B.n209 VSUBS 0.007329f
C250 B.n210 VSUBS 0.007329f
C251 B.n211 VSUBS 0.007329f
C252 B.n212 VSUBS 0.007329f
C253 B.n213 VSUBS 0.007329f
C254 B.n214 VSUBS 0.007329f
C255 B.n215 VSUBS 0.007329f
C256 B.n216 VSUBS 0.007329f
C257 B.n217 VSUBS 0.007329f
C258 B.n218 VSUBS 0.007329f
C259 B.n219 VSUBS 0.007329f
C260 B.n220 VSUBS 0.007329f
C261 B.n221 VSUBS 0.007329f
C262 B.n222 VSUBS 0.007329f
C263 B.n223 VSUBS 0.007329f
C264 B.n224 VSUBS 0.007329f
C265 B.n225 VSUBS 0.017201f
C266 B.n226 VSUBS 0.018149f
C267 B.n227 VSUBS 0.018149f
C268 B.n228 VSUBS 0.007329f
C269 B.n229 VSUBS 0.007329f
C270 B.n230 VSUBS 0.007329f
C271 B.n231 VSUBS 0.007329f
C272 B.n232 VSUBS 0.007329f
C273 B.n233 VSUBS 0.007329f
C274 B.n234 VSUBS 0.007329f
C275 B.n235 VSUBS 0.007329f
C276 B.n236 VSUBS 0.007329f
C277 B.n237 VSUBS 0.007329f
C278 B.n238 VSUBS 0.007329f
C279 B.n239 VSUBS 0.007329f
C280 B.n240 VSUBS 0.007329f
C281 B.n241 VSUBS 0.007329f
C282 B.n242 VSUBS 0.007329f
C283 B.n243 VSUBS 0.007329f
C284 B.n244 VSUBS 0.007329f
C285 B.n245 VSUBS 0.007329f
C286 B.n246 VSUBS 0.007329f
C287 B.n247 VSUBS 0.007329f
C288 B.n248 VSUBS 0.007329f
C289 B.n249 VSUBS 0.007329f
C290 B.n250 VSUBS 0.007329f
C291 B.n251 VSUBS 0.007329f
C292 B.n252 VSUBS 0.007329f
C293 B.n253 VSUBS 0.007329f
C294 B.n254 VSUBS 0.006898f
C295 B.n255 VSUBS 0.01698f
C296 B.n256 VSUBS 0.004095f
C297 B.n257 VSUBS 0.007329f
C298 B.n258 VSUBS 0.007329f
C299 B.n259 VSUBS 0.007329f
C300 B.n260 VSUBS 0.007329f
C301 B.n261 VSUBS 0.007329f
C302 B.n262 VSUBS 0.007329f
C303 B.n263 VSUBS 0.007329f
C304 B.n264 VSUBS 0.007329f
C305 B.n265 VSUBS 0.007329f
C306 B.n266 VSUBS 0.007329f
C307 B.n267 VSUBS 0.007329f
C308 B.n268 VSUBS 0.007329f
C309 B.n269 VSUBS 0.004095f
C310 B.n270 VSUBS 0.007329f
C311 B.n271 VSUBS 0.007329f
C312 B.n272 VSUBS 0.007329f
C313 B.n273 VSUBS 0.007329f
C314 B.n274 VSUBS 0.007329f
C315 B.n275 VSUBS 0.007329f
C316 B.n276 VSUBS 0.007329f
C317 B.n277 VSUBS 0.007329f
C318 B.n278 VSUBS 0.007329f
C319 B.n279 VSUBS 0.007329f
C320 B.n280 VSUBS 0.007329f
C321 B.n281 VSUBS 0.007329f
C322 B.n282 VSUBS 0.007329f
C323 B.n283 VSUBS 0.007329f
C324 B.n284 VSUBS 0.007329f
C325 B.n285 VSUBS 0.007329f
C326 B.n286 VSUBS 0.007329f
C327 B.n287 VSUBS 0.007329f
C328 B.n288 VSUBS 0.007329f
C329 B.n289 VSUBS 0.007329f
C330 B.n290 VSUBS 0.007329f
C331 B.n291 VSUBS 0.007329f
C332 B.n292 VSUBS 0.007329f
C333 B.n293 VSUBS 0.007329f
C334 B.n294 VSUBS 0.007329f
C335 B.n295 VSUBS 0.007329f
C336 B.n296 VSUBS 0.007329f
C337 B.n297 VSUBS 0.007329f
C338 B.n298 VSUBS 0.018149f
C339 B.n299 VSUBS 0.017201f
C340 B.n300 VSUBS 0.017201f
C341 B.n301 VSUBS 0.007329f
C342 B.n302 VSUBS 0.007329f
C343 B.n303 VSUBS 0.007329f
C344 B.n304 VSUBS 0.007329f
C345 B.n305 VSUBS 0.007329f
C346 B.n306 VSUBS 0.007329f
C347 B.n307 VSUBS 0.007329f
C348 B.n308 VSUBS 0.007329f
C349 B.n309 VSUBS 0.007329f
C350 B.n310 VSUBS 0.007329f
C351 B.n311 VSUBS 0.007329f
C352 B.n312 VSUBS 0.007329f
C353 B.n313 VSUBS 0.007329f
C354 B.n314 VSUBS 0.007329f
C355 B.n315 VSUBS 0.007329f
C356 B.n316 VSUBS 0.007329f
C357 B.n317 VSUBS 0.007329f
C358 B.n318 VSUBS 0.007329f
C359 B.n319 VSUBS 0.009563f
C360 B.n320 VSUBS 0.010188f
C361 B.n321 VSUBS 0.020259f
C362 VDD2.t3 VSUBS 0.079911f
C363 VDD2.t0 VSUBS 0.079911f
C364 VDD2.n0 VSUBS 0.700134f
C365 VDD2.t1 VSUBS 0.079911f
C366 VDD2.t2 VSUBS 0.079911f
C367 VDD2.n1 VSUBS 0.482574f
C368 VDD2.n2 VSUBS 2.34534f
C369 VN.t0 VSUBS 0.188559f
C370 VN.t3 VSUBS 0.188551f
C371 VN.n0 VSUBS 0.182471f
C372 VN.t1 VSUBS 0.188559f
C373 VN.t2 VSUBS 0.188551f
C374 VN.n1 VSUBS 0.516212f
C375 VDD1.t1 VSUBS 0.078205f
C376 VDD1.t0 VSUBS 0.078205f
C377 VDD1.n0 VSUBS 0.472473f
C378 VDD1.t2 VSUBS 0.078205f
C379 VDD1.t3 VSUBS 0.078205f
C380 VDD1.n1 VSUBS 0.698014f
C381 VTAIL.t0 VSUBS 0.540937f
C382 VTAIL.n0 VSUBS 0.419252f
C383 VTAIL.t3 VSUBS 0.540937f
C384 VTAIL.n1 VSUBS 0.436646f
C385 VTAIL.t5 VSUBS 0.540937f
C386 VTAIL.n2 VSUBS 0.981481f
C387 VTAIL.t2 VSUBS 0.540939f
C388 VTAIL.n3 VSUBS 0.981479f
C389 VTAIL.t1 VSUBS 0.540939f
C390 VTAIL.n4 VSUBS 0.436644f
C391 VTAIL.t4 VSUBS 0.540939f
C392 VTAIL.n5 VSUBS 0.436644f
C393 VTAIL.t6 VSUBS 0.540937f
C394 VTAIL.n6 VSUBS 0.981481f
C395 VTAIL.t7 VSUBS 0.540937f
C396 VTAIL.n7 VSUBS 0.956324f
C397 VP.t3 VSUBS 0.311128f
C398 VP.t2 VSUBS 0.311142f
C399 VP.n0 VSUBS 0.83529f
C400 VP.n1 VSUBS 2.7568f
C401 VP.t1 VSUBS 0.30223f
C402 VP.n2 VSUBS 0.159376f
C403 VP.t0 VSUBS 0.30223f
C404 VP.n3 VSUBS 0.159376f
C405 VP.n4 VSUBS 0.044281f
.ends

