* NGSPICE file created from diff_pair_sample_0365.ext - technology: sky130A

.subckt diff_pair_sample_0365 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 w_n1378_n2336# sky130_fd_pr__pfet_01v8 ad=2.6598 pd=14.42 as=2.6598 ps=14.42 w=6.82 l=0.69
X1 VDD1.t1 VP.t0 VTAIL.t0 w_n1378_n2336# sky130_fd_pr__pfet_01v8 ad=2.6598 pd=14.42 as=2.6598 ps=14.42 w=6.82 l=0.69
X2 B.t11 B.t9 B.t10 w_n1378_n2336# sky130_fd_pr__pfet_01v8 ad=2.6598 pd=14.42 as=0 ps=0 w=6.82 l=0.69
X3 B.t8 B.t6 B.t7 w_n1378_n2336# sky130_fd_pr__pfet_01v8 ad=2.6598 pd=14.42 as=0 ps=0 w=6.82 l=0.69
X4 B.t5 B.t3 B.t4 w_n1378_n2336# sky130_fd_pr__pfet_01v8 ad=2.6598 pd=14.42 as=0 ps=0 w=6.82 l=0.69
X5 VDD2.t0 VN.t1 VTAIL.t2 w_n1378_n2336# sky130_fd_pr__pfet_01v8 ad=2.6598 pd=14.42 as=2.6598 ps=14.42 w=6.82 l=0.69
X6 B.t2 B.t0 B.t1 w_n1378_n2336# sky130_fd_pr__pfet_01v8 ad=2.6598 pd=14.42 as=0 ps=0 w=6.82 l=0.69
X7 VDD1.t0 VP.t1 VTAIL.t1 w_n1378_n2336# sky130_fd_pr__pfet_01v8 ad=2.6598 pd=14.42 as=2.6598 ps=14.42 w=6.82 l=0.69
R0 VN VN.t1 493.2
R1 VN VN.t0 457.188
R2 VTAIL.n1 VTAIL.t2 76.306
R3 VTAIL.n3 VTAIL.t3 76.3059
R4 VTAIL.n0 VTAIL.t1 76.3059
R5 VTAIL.n2 VTAIL.t0 76.3059
R6 VTAIL.n1 VTAIL.n0 20.0221
R7 VTAIL.n3 VTAIL.n2 19.1427
R8 VTAIL.n2 VTAIL.n1 0.909983
R9 VTAIL VTAIL.n0 0.748345
R10 VTAIL VTAIL.n3 0.162138
R11 VDD2.n0 VDD2.t1 124.299
R12 VDD2.n0 VDD2.t0 92.9847
R13 VDD2 VDD2.n0 0.278517
R14 VP.n0 VP.t0 492.818
R15 VP.n0 VP.t1 457.137
R16 VP VP.n0 0.0516364
R17 VDD1 VDD1.t0 125.043
R18 VDD1 VDD1.t1 93.2627
R19 B.n259 B.n44 585
R20 B.n261 B.n260 585
R21 B.n262 B.n43 585
R22 B.n264 B.n263 585
R23 B.n265 B.n42 585
R24 B.n267 B.n266 585
R25 B.n268 B.n41 585
R26 B.n270 B.n269 585
R27 B.n271 B.n40 585
R28 B.n273 B.n272 585
R29 B.n274 B.n39 585
R30 B.n276 B.n275 585
R31 B.n277 B.n38 585
R32 B.n279 B.n278 585
R33 B.n280 B.n37 585
R34 B.n282 B.n281 585
R35 B.n283 B.n36 585
R36 B.n285 B.n284 585
R37 B.n286 B.n35 585
R38 B.n288 B.n287 585
R39 B.n289 B.n34 585
R40 B.n291 B.n290 585
R41 B.n292 B.n33 585
R42 B.n294 B.n293 585
R43 B.n295 B.n32 585
R44 B.n297 B.n296 585
R45 B.n299 B.n29 585
R46 B.n301 B.n300 585
R47 B.n302 B.n28 585
R48 B.n304 B.n303 585
R49 B.n305 B.n27 585
R50 B.n307 B.n306 585
R51 B.n308 B.n26 585
R52 B.n310 B.n309 585
R53 B.n311 B.n25 585
R54 B.n313 B.n312 585
R55 B.n315 B.n314 585
R56 B.n316 B.n21 585
R57 B.n318 B.n317 585
R58 B.n319 B.n20 585
R59 B.n321 B.n320 585
R60 B.n322 B.n19 585
R61 B.n324 B.n323 585
R62 B.n325 B.n18 585
R63 B.n327 B.n326 585
R64 B.n328 B.n17 585
R65 B.n330 B.n329 585
R66 B.n331 B.n16 585
R67 B.n333 B.n332 585
R68 B.n334 B.n15 585
R69 B.n336 B.n335 585
R70 B.n337 B.n14 585
R71 B.n339 B.n338 585
R72 B.n340 B.n13 585
R73 B.n342 B.n341 585
R74 B.n343 B.n12 585
R75 B.n345 B.n344 585
R76 B.n346 B.n11 585
R77 B.n348 B.n347 585
R78 B.n349 B.n10 585
R79 B.n351 B.n350 585
R80 B.n352 B.n9 585
R81 B.n258 B.n257 585
R82 B.n256 B.n45 585
R83 B.n255 B.n254 585
R84 B.n253 B.n46 585
R85 B.n252 B.n251 585
R86 B.n250 B.n47 585
R87 B.n249 B.n248 585
R88 B.n247 B.n48 585
R89 B.n246 B.n245 585
R90 B.n244 B.n49 585
R91 B.n243 B.n242 585
R92 B.n241 B.n50 585
R93 B.n240 B.n239 585
R94 B.n238 B.n51 585
R95 B.n237 B.n236 585
R96 B.n235 B.n52 585
R97 B.n234 B.n233 585
R98 B.n232 B.n53 585
R99 B.n231 B.n230 585
R100 B.n229 B.n54 585
R101 B.n228 B.n227 585
R102 B.n226 B.n55 585
R103 B.n225 B.n224 585
R104 B.n223 B.n56 585
R105 B.n222 B.n221 585
R106 B.n220 B.n57 585
R107 B.n219 B.n218 585
R108 B.n217 B.n58 585
R109 B.n216 B.n215 585
R110 B.n121 B.n94 585
R111 B.n123 B.n122 585
R112 B.n124 B.n93 585
R113 B.n126 B.n125 585
R114 B.n127 B.n92 585
R115 B.n129 B.n128 585
R116 B.n130 B.n91 585
R117 B.n132 B.n131 585
R118 B.n133 B.n90 585
R119 B.n135 B.n134 585
R120 B.n136 B.n89 585
R121 B.n138 B.n137 585
R122 B.n139 B.n88 585
R123 B.n141 B.n140 585
R124 B.n142 B.n87 585
R125 B.n144 B.n143 585
R126 B.n145 B.n86 585
R127 B.n147 B.n146 585
R128 B.n148 B.n85 585
R129 B.n150 B.n149 585
R130 B.n151 B.n84 585
R131 B.n153 B.n152 585
R132 B.n154 B.n83 585
R133 B.n156 B.n155 585
R134 B.n157 B.n82 585
R135 B.n159 B.n158 585
R136 B.n161 B.n79 585
R137 B.n163 B.n162 585
R138 B.n164 B.n78 585
R139 B.n166 B.n165 585
R140 B.n167 B.n77 585
R141 B.n169 B.n168 585
R142 B.n170 B.n76 585
R143 B.n172 B.n171 585
R144 B.n173 B.n75 585
R145 B.n175 B.n174 585
R146 B.n177 B.n176 585
R147 B.n178 B.n71 585
R148 B.n180 B.n179 585
R149 B.n181 B.n70 585
R150 B.n183 B.n182 585
R151 B.n184 B.n69 585
R152 B.n186 B.n185 585
R153 B.n187 B.n68 585
R154 B.n189 B.n188 585
R155 B.n190 B.n67 585
R156 B.n192 B.n191 585
R157 B.n193 B.n66 585
R158 B.n195 B.n194 585
R159 B.n196 B.n65 585
R160 B.n198 B.n197 585
R161 B.n199 B.n64 585
R162 B.n201 B.n200 585
R163 B.n202 B.n63 585
R164 B.n204 B.n203 585
R165 B.n205 B.n62 585
R166 B.n207 B.n206 585
R167 B.n208 B.n61 585
R168 B.n210 B.n209 585
R169 B.n211 B.n60 585
R170 B.n213 B.n212 585
R171 B.n214 B.n59 585
R172 B.n120 B.n119 585
R173 B.n118 B.n95 585
R174 B.n117 B.n116 585
R175 B.n115 B.n96 585
R176 B.n114 B.n113 585
R177 B.n112 B.n97 585
R178 B.n111 B.n110 585
R179 B.n109 B.n98 585
R180 B.n108 B.n107 585
R181 B.n106 B.n99 585
R182 B.n105 B.n104 585
R183 B.n103 B.n100 585
R184 B.n102 B.n101 585
R185 B.n2 B.n0 585
R186 B.n373 B.n1 585
R187 B.n372 B.n371 585
R188 B.n370 B.n3 585
R189 B.n369 B.n368 585
R190 B.n367 B.n4 585
R191 B.n366 B.n365 585
R192 B.n364 B.n5 585
R193 B.n363 B.n362 585
R194 B.n361 B.n6 585
R195 B.n360 B.n359 585
R196 B.n358 B.n7 585
R197 B.n357 B.n356 585
R198 B.n355 B.n8 585
R199 B.n354 B.n353 585
R200 B.n375 B.n374 585
R201 B.n121 B.n120 554.963
R202 B.n354 B.n9 554.963
R203 B.n216 B.n59 554.963
R204 B.n259 B.n258 554.963
R205 B.n72 B.t6 441.296
R206 B.n80 B.t9 441.296
R207 B.n22 B.t0 441.296
R208 B.n30 B.t3 441.296
R209 B.n120 B.n95 163.367
R210 B.n116 B.n95 163.367
R211 B.n116 B.n115 163.367
R212 B.n115 B.n114 163.367
R213 B.n114 B.n97 163.367
R214 B.n110 B.n97 163.367
R215 B.n110 B.n109 163.367
R216 B.n109 B.n108 163.367
R217 B.n108 B.n99 163.367
R218 B.n104 B.n99 163.367
R219 B.n104 B.n103 163.367
R220 B.n103 B.n102 163.367
R221 B.n102 B.n2 163.367
R222 B.n374 B.n2 163.367
R223 B.n374 B.n373 163.367
R224 B.n373 B.n372 163.367
R225 B.n372 B.n3 163.367
R226 B.n368 B.n3 163.367
R227 B.n368 B.n367 163.367
R228 B.n367 B.n366 163.367
R229 B.n366 B.n5 163.367
R230 B.n362 B.n5 163.367
R231 B.n362 B.n361 163.367
R232 B.n361 B.n360 163.367
R233 B.n360 B.n7 163.367
R234 B.n356 B.n7 163.367
R235 B.n356 B.n355 163.367
R236 B.n355 B.n354 163.367
R237 B.n122 B.n121 163.367
R238 B.n122 B.n93 163.367
R239 B.n126 B.n93 163.367
R240 B.n127 B.n126 163.367
R241 B.n128 B.n127 163.367
R242 B.n128 B.n91 163.367
R243 B.n132 B.n91 163.367
R244 B.n133 B.n132 163.367
R245 B.n134 B.n133 163.367
R246 B.n134 B.n89 163.367
R247 B.n138 B.n89 163.367
R248 B.n139 B.n138 163.367
R249 B.n140 B.n139 163.367
R250 B.n140 B.n87 163.367
R251 B.n144 B.n87 163.367
R252 B.n145 B.n144 163.367
R253 B.n146 B.n145 163.367
R254 B.n146 B.n85 163.367
R255 B.n150 B.n85 163.367
R256 B.n151 B.n150 163.367
R257 B.n152 B.n151 163.367
R258 B.n152 B.n83 163.367
R259 B.n156 B.n83 163.367
R260 B.n157 B.n156 163.367
R261 B.n158 B.n157 163.367
R262 B.n158 B.n79 163.367
R263 B.n163 B.n79 163.367
R264 B.n164 B.n163 163.367
R265 B.n165 B.n164 163.367
R266 B.n165 B.n77 163.367
R267 B.n169 B.n77 163.367
R268 B.n170 B.n169 163.367
R269 B.n171 B.n170 163.367
R270 B.n171 B.n75 163.367
R271 B.n175 B.n75 163.367
R272 B.n176 B.n175 163.367
R273 B.n176 B.n71 163.367
R274 B.n180 B.n71 163.367
R275 B.n181 B.n180 163.367
R276 B.n182 B.n181 163.367
R277 B.n182 B.n69 163.367
R278 B.n186 B.n69 163.367
R279 B.n187 B.n186 163.367
R280 B.n188 B.n187 163.367
R281 B.n188 B.n67 163.367
R282 B.n192 B.n67 163.367
R283 B.n193 B.n192 163.367
R284 B.n194 B.n193 163.367
R285 B.n194 B.n65 163.367
R286 B.n198 B.n65 163.367
R287 B.n199 B.n198 163.367
R288 B.n200 B.n199 163.367
R289 B.n200 B.n63 163.367
R290 B.n204 B.n63 163.367
R291 B.n205 B.n204 163.367
R292 B.n206 B.n205 163.367
R293 B.n206 B.n61 163.367
R294 B.n210 B.n61 163.367
R295 B.n211 B.n210 163.367
R296 B.n212 B.n211 163.367
R297 B.n212 B.n59 163.367
R298 B.n217 B.n216 163.367
R299 B.n218 B.n217 163.367
R300 B.n218 B.n57 163.367
R301 B.n222 B.n57 163.367
R302 B.n223 B.n222 163.367
R303 B.n224 B.n223 163.367
R304 B.n224 B.n55 163.367
R305 B.n228 B.n55 163.367
R306 B.n229 B.n228 163.367
R307 B.n230 B.n229 163.367
R308 B.n230 B.n53 163.367
R309 B.n234 B.n53 163.367
R310 B.n235 B.n234 163.367
R311 B.n236 B.n235 163.367
R312 B.n236 B.n51 163.367
R313 B.n240 B.n51 163.367
R314 B.n241 B.n240 163.367
R315 B.n242 B.n241 163.367
R316 B.n242 B.n49 163.367
R317 B.n246 B.n49 163.367
R318 B.n247 B.n246 163.367
R319 B.n248 B.n247 163.367
R320 B.n248 B.n47 163.367
R321 B.n252 B.n47 163.367
R322 B.n253 B.n252 163.367
R323 B.n254 B.n253 163.367
R324 B.n254 B.n45 163.367
R325 B.n258 B.n45 163.367
R326 B.n350 B.n9 163.367
R327 B.n350 B.n349 163.367
R328 B.n349 B.n348 163.367
R329 B.n348 B.n11 163.367
R330 B.n344 B.n11 163.367
R331 B.n344 B.n343 163.367
R332 B.n343 B.n342 163.367
R333 B.n342 B.n13 163.367
R334 B.n338 B.n13 163.367
R335 B.n338 B.n337 163.367
R336 B.n337 B.n336 163.367
R337 B.n336 B.n15 163.367
R338 B.n332 B.n15 163.367
R339 B.n332 B.n331 163.367
R340 B.n331 B.n330 163.367
R341 B.n330 B.n17 163.367
R342 B.n326 B.n17 163.367
R343 B.n326 B.n325 163.367
R344 B.n325 B.n324 163.367
R345 B.n324 B.n19 163.367
R346 B.n320 B.n19 163.367
R347 B.n320 B.n319 163.367
R348 B.n319 B.n318 163.367
R349 B.n318 B.n21 163.367
R350 B.n314 B.n21 163.367
R351 B.n314 B.n313 163.367
R352 B.n313 B.n25 163.367
R353 B.n309 B.n25 163.367
R354 B.n309 B.n308 163.367
R355 B.n308 B.n307 163.367
R356 B.n307 B.n27 163.367
R357 B.n303 B.n27 163.367
R358 B.n303 B.n302 163.367
R359 B.n302 B.n301 163.367
R360 B.n301 B.n29 163.367
R361 B.n296 B.n29 163.367
R362 B.n296 B.n295 163.367
R363 B.n295 B.n294 163.367
R364 B.n294 B.n33 163.367
R365 B.n290 B.n33 163.367
R366 B.n290 B.n289 163.367
R367 B.n289 B.n288 163.367
R368 B.n288 B.n35 163.367
R369 B.n284 B.n35 163.367
R370 B.n284 B.n283 163.367
R371 B.n283 B.n282 163.367
R372 B.n282 B.n37 163.367
R373 B.n278 B.n37 163.367
R374 B.n278 B.n277 163.367
R375 B.n277 B.n276 163.367
R376 B.n276 B.n39 163.367
R377 B.n272 B.n39 163.367
R378 B.n272 B.n271 163.367
R379 B.n271 B.n270 163.367
R380 B.n270 B.n41 163.367
R381 B.n266 B.n41 163.367
R382 B.n266 B.n265 163.367
R383 B.n265 B.n264 163.367
R384 B.n264 B.n43 163.367
R385 B.n260 B.n43 163.367
R386 B.n260 B.n259 163.367
R387 B.n72 B.t8 129.91
R388 B.n30 B.t4 129.91
R389 B.n80 B.t11 129.903
R390 B.n22 B.t1 129.903
R391 B.n73 B.t7 110.127
R392 B.n31 B.t5 110.127
R393 B.n81 B.t10 110.121
R394 B.n23 B.t2 110.121
R395 B.n74 B.n73 59.5399
R396 B.n160 B.n81 59.5399
R397 B.n24 B.n23 59.5399
R398 B.n298 B.n31 59.5399
R399 B.n353 B.n352 36.059
R400 B.n215 B.n214 36.059
R401 B.n119 B.n94 36.059
R402 B.n257 B.n44 36.059
R403 B.n73 B.n72 19.7823
R404 B.n81 B.n80 19.7823
R405 B.n23 B.n22 19.7823
R406 B.n31 B.n30 19.7823
R407 B B.n375 18.0485
R408 B.n352 B.n351 10.6151
R409 B.n351 B.n10 10.6151
R410 B.n347 B.n10 10.6151
R411 B.n347 B.n346 10.6151
R412 B.n346 B.n345 10.6151
R413 B.n345 B.n12 10.6151
R414 B.n341 B.n12 10.6151
R415 B.n341 B.n340 10.6151
R416 B.n340 B.n339 10.6151
R417 B.n339 B.n14 10.6151
R418 B.n335 B.n14 10.6151
R419 B.n335 B.n334 10.6151
R420 B.n334 B.n333 10.6151
R421 B.n333 B.n16 10.6151
R422 B.n329 B.n16 10.6151
R423 B.n329 B.n328 10.6151
R424 B.n328 B.n327 10.6151
R425 B.n327 B.n18 10.6151
R426 B.n323 B.n18 10.6151
R427 B.n323 B.n322 10.6151
R428 B.n322 B.n321 10.6151
R429 B.n321 B.n20 10.6151
R430 B.n317 B.n20 10.6151
R431 B.n317 B.n316 10.6151
R432 B.n316 B.n315 10.6151
R433 B.n312 B.n311 10.6151
R434 B.n311 B.n310 10.6151
R435 B.n310 B.n26 10.6151
R436 B.n306 B.n26 10.6151
R437 B.n306 B.n305 10.6151
R438 B.n305 B.n304 10.6151
R439 B.n304 B.n28 10.6151
R440 B.n300 B.n28 10.6151
R441 B.n300 B.n299 10.6151
R442 B.n297 B.n32 10.6151
R443 B.n293 B.n32 10.6151
R444 B.n293 B.n292 10.6151
R445 B.n292 B.n291 10.6151
R446 B.n291 B.n34 10.6151
R447 B.n287 B.n34 10.6151
R448 B.n287 B.n286 10.6151
R449 B.n286 B.n285 10.6151
R450 B.n285 B.n36 10.6151
R451 B.n281 B.n36 10.6151
R452 B.n281 B.n280 10.6151
R453 B.n280 B.n279 10.6151
R454 B.n279 B.n38 10.6151
R455 B.n275 B.n38 10.6151
R456 B.n275 B.n274 10.6151
R457 B.n274 B.n273 10.6151
R458 B.n273 B.n40 10.6151
R459 B.n269 B.n40 10.6151
R460 B.n269 B.n268 10.6151
R461 B.n268 B.n267 10.6151
R462 B.n267 B.n42 10.6151
R463 B.n263 B.n42 10.6151
R464 B.n263 B.n262 10.6151
R465 B.n262 B.n261 10.6151
R466 B.n261 B.n44 10.6151
R467 B.n215 B.n58 10.6151
R468 B.n219 B.n58 10.6151
R469 B.n220 B.n219 10.6151
R470 B.n221 B.n220 10.6151
R471 B.n221 B.n56 10.6151
R472 B.n225 B.n56 10.6151
R473 B.n226 B.n225 10.6151
R474 B.n227 B.n226 10.6151
R475 B.n227 B.n54 10.6151
R476 B.n231 B.n54 10.6151
R477 B.n232 B.n231 10.6151
R478 B.n233 B.n232 10.6151
R479 B.n233 B.n52 10.6151
R480 B.n237 B.n52 10.6151
R481 B.n238 B.n237 10.6151
R482 B.n239 B.n238 10.6151
R483 B.n239 B.n50 10.6151
R484 B.n243 B.n50 10.6151
R485 B.n244 B.n243 10.6151
R486 B.n245 B.n244 10.6151
R487 B.n245 B.n48 10.6151
R488 B.n249 B.n48 10.6151
R489 B.n250 B.n249 10.6151
R490 B.n251 B.n250 10.6151
R491 B.n251 B.n46 10.6151
R492 B.n255 B.n46 10.6151
R493 B.n256 B.n255 10.6151
R494 B.n257 B.n256 10.6151
R495 B.n123 B.n94 10.6151
R496 B.n124 B.n123 10.6151
R497 B.n125 B.n124 10.6151
R498 B.n125 B.n92 10.6151
R499 B.n129 B.n92 10.6151
R500 B.n130 B.n129 10.6151
R501 B.n131 B.n130 10.6151
R502 B.n131 B.n90 10.6151
R503 B.n135 B.n90 10.6151
R504 B.n136 B.n135 10.6151
R505 B.n137 B.n136 10.6151
R506 B.n137 B.n88 10.6151
R507 B.n141 B.n88 10.6151
R508 B.n142 B.n141 10.6151
R509 B.n143 B.n142 10.6151
R510 B.n143 B.n86 10.6151
R511 B.n147 B.n86 10.6151
R512 B.n148 B.n147 10.6151
R513 B.n149 B.n148 10.6151
R514 B.n149 B.n84 10.6151
R515 B.n153 B.n84 10.6151
R516 B.n154 B.n153 10.6151
R517 B.n155 B.n154 10.6151
R518 B.n155 B.n82 10.6151
R519 B.n159 B.n82 10.6151
R520 B.n162 B.n161 10.6151
R521 B.n162 B.n78 10.6151
R522 B.n166 B.n78 10.6151
R523 B.n167 B.n166 10.6151
R524 B.n168 B.n167 10.6151
R525 B.n168 B.n76 10.6151
R526 B.n172 B.n76 10.6151
R527 B.n173 B.n172 10.6151
R528 B.n174 B.n173 10.6151
R529 B.n178 B.n177 10.6151
R530 B.n179 B.n178 10.6151
R531 B.n179 B.n70 10.6151
R532 B.n183 B.n70 10.6151
R533 B.n184 B.n183 10.6151
R534 B.n185 B.n184 10.6151
R535 B.n185 B.n68 10.6151
R536 B.n189 B.n68 10.6151
R537 B.n190 B.n189 10.6151
R538 B.n191 B.n190 10.6151
R539 B.n191 B.n66 10.6151
R540 B.n195 B.n66 10.6151
R541 B.n196 B.n195 10.6151
R542 B.n197 B.n196 10.6151
R543 B.n197 B.n64 10.6151
R544 B.n201 B.n64 10.6151
R545 B.n202 B.n201 10.6151
R546 B.n203 B.n202 10.6151
R547 B.n203 B.n62 10.6151
R548 B.n207 B.n62 10.6151
R549 B.n208 B.n207 10.6151
R550 B.n209 B.n208 10.6151
R551 B.n209 B.n60 10.6151
R552 B.n213 B.n60 10.6151
R553 B.n214 B.n213 10.6151
R554 B.n119 B.n118 10.6151
R555 B.n118 B.n117 10.6151
R556 B.n117 B.n96 10.6151
R557 B.n113 B.n96 10.6151
R558 B.n113 B.n112 10.6151
R559 B.n112 B.n111 10.6151
R560 B.n111 B.n98 10.6151
R561 B.n107 B.n98 10.6151
R562 B.n107 B.n106 10.6151
R563 B.n106 B.n105 10.6151
R564 B.n105 B.n100 10.6151
R565 B.n101 B.n100 10.6151
R566 B.n101 B.n0 10.6151
R567 B.n371 B.n1 10.6151
R568 B.n371 B.n370 10.6151
R569 B.n370 B.n369 10.6151
R570 B.n369 B.n4 10.6151
R571 B.n365 B.n4 10.6151
R572 B.n365 B.n364 10.6151
R573 B.n364 B.n363 10.6151
R574 B.n363 B.n6 10.6151
R575 B.n359 B.n6 10.6151
R576 B.n359 B.n358 10.6151
R577 B.n358 B.n357 10.6151
R578 B.n357 B.n8 10.6151
R579 B.n353 B.n8 10.6151
R580 B.n315 B.n24 8.74196
R581 B.n298 B.n297 8.74196
R582 B.n160 B.n159 8.74196
R583 B.n177 B.n74 8.74196
R584 B.n375 B.n0 2.81026
R585 B.n375 B.n1 2.81026
R586 B.n312 B.n24 1.87367
R587 B.n299 B.n298 1.87367
R588 B.n161 B.n160 1.87367
R589 B.n174 B.n74 1.87367
C0 B VTAIL 1.78795f
C1 VN B 0.662161f
C2 VDD1 B 1.03728f
C3 VP B 0.936308f
C4 B w_n1378_n2336# 5.29788f
C5 VN VTAIL 0.986096f
C6 VDD1 VTAIL 3.75357f
C7 VP VTAIL 1.00049f
C8 VTAIL w_n1378_n2336# 2.05687f
C9 VDD1 VN 0.148251f
C10 VN VP 3.60008f
C11 VDD2 B 1.05172f
C12 VDD1 VP 1.32486f
C13 VN w_n1378_n2336# 1.6452f
C14 VDD1 w_n1378_n2336# 1.18853f
C15 VP w_n1378_n2336# 1.81661f
C16 VDD2 VTAIL 3.79022f
C17 VDD2 VN 1.22222f
C18 VDD1 VDD2 0.459723f
C19 VDD2 VP 0.253459f
C20 VDD2 w_n1378_n2336# 1.19308f
C21 VDD2 VSUBS 0.56298f
C22 VDD1 VSUBS 2.656066f
C23 VTAIL VSUBS 0.476189f
C24 VN VSUBS 3.81195f
C25 VP VSUBS 0.863435f
C26 B VSUBS 2.049735f
C27 w_n1378_n2336# VSUBS 40.066696f
C28 B.n0 VSUBS 0.003989f
C29 B.n1 VSUBS 0.003989f
C30 B.n2 VSUBS 0.006308f
C31 B.n3 VSUBS 0.006308f
C32 B.n4 VSUBS 0.006308f
C33 B.n5 VSUBS 0.006308f
C34 B.n6 VSUBS 0.006308f
C35 B.n7 VSUBS 0.006308f
C36 B.n8 VSUBS 0.006308f
C37 B.n9 VSUBS 0.016025f
C38 B.n10 VSUBS 0.006308f
C39 B.n11 VSUBS 0.006308f
C40 B.n12 VSUBS 0.006308f
C41 B.n13 VSUBS 0.006308f
C42 B.n14 VSUBS 0.006308f
C43 B.n15 VSUBS 0.006308f
C44 B.n16 VSUBS 0.006308f
C45 B.n17 VSUBS 0.006308f
C46 B.n18 VSUBS 0.006308f
C47 B.n19 VSUBS 0.006308f
C48 B.n20 VSUBS 0.006308f
C49 B.n21 VSUBS 0.006308f
C50 B.t2 VSUBS 0.184294f
C51 B.t1 VSUBS 0.191589f
C52 B.t0 VSUBS 0.181595f
C53 B.n22 VSUBS 0.084487f
C54 B.n23 VSUBS 0.056898f
C55 B.n24 VSUBS 0.014614f
C56 B.n25 VSUBS 0.006308f
C57 B.n26 VSUBS 0.006308f
C58 B.n27 VSUBS 0.006308f
C59 B.n28 VSUBS 0.006308f
C60 B.n29 VSUBS 0.006308f
C61 B.t5 VSUBS 0.184293f
C62 B.t4 VSUBS 0.191588f
C63 B.t3 VSUBS 0.181595f
C64 B.n30 VSUBS 0.084489f
C65 B.n31 VSUBS 0.056898f
C66 B.n32 VSUBS 0.006308f
C67 B.n33 VSUBS 0.006308f
C68 B.n34 VSUBS 0.006308f
C69 B.n35 VSUBS 0.006308f
C70 B.n36 VSUBS 0.006308f
C71 B.n37 VSUBS 0.006308f
C72 B.n38 VSUBS 0.006308f
C73 B.n39 VSUBS 0.006308f
C74 B.n40 VSUBS 0.006308f
C75 B.n41 VSUBS 0.006308f
C76 B.n42 VSUBS 0.006308f
C77 B.n43 VSUBS 0.006308f
C78 B.n44 VSUBS 0.015349f
C79 B.n45 VSUBS 0.006308f
C80 B.n46 VSUBS 0.006308f
C81 B.n47 VSUBS 0.006308f
C82 B.n48 VSUBS 0.006308f
C83 B.n49 VSUBS 0.006308f
C84 B.n50 VSUBS 0.006308f
C85 B.n51 VSUBS 0.006308f
C86 B.n52 VSUBS 0.006308f
C87 B.n53 VSUBS 0.006308f
C88 B.n54 VSUBS 0.006308f
C89 B.n55 VSUBS 0.006308f
C90 B.n56 VSUBS 0.006308f
C91 B.n57 VSUBS 0.006308f
C92 B.n58 VSUBS 0.006308f
C93 B.n59 VSUBS 0.016025f
C94 B.n60 VSUBS 0.006308f
C95 B.n61 VSUBS 0.006308f
C96 B.n62 VSUBS 0.006308f
C97 B.n63 VSUBS 0.006308f
C98 B.n64 VSUBS 0.006308f
C99 B.n65 VSUBS 0.006308f
C100 B.n66 VSUBS 0.006308f
C101 B.n67 VSUBS 0.006308f
C102 B.n68 VSUBS 0.006308f
C103 B.n69 VSUBS 0.006308f
C104 B.n70 VSUBS 0.006308f
C105 B.n71 VSUBS 0.006308f
C106 B.t7 VSUBS 0.184293f
C107 B.t8 VSUBS 0.191588f
C108 B.t6 VSUBS 0.181595f
C109 B.n72 VSUBS 0.084489f
C110 B.n73 VSUBS 0.056898f
C111 B.n74 VSUBS 0.014614f
C112 B.n75 VSUBS 0.006308f
C113 B.n76 VSUBS 0.006308f
C114 B.n77 VSUBS 0.006308f
C115 B.n78 VSUBS 0.006308f
C116 B.n79 VSUBS 0.006308f
C117 B.t10 VSUBS 0.184294f
C118 B.t11 VSUBS 0.191589f
C119 B.t9 VSUBS 0.181595f
C120 B.n80 VSUBS 0.084487f
C121 B.n81 VSUBS 0.056898f
C122 B.n82 VSUBS 0.006308f
C123 B.n83 VSUBS 0.006308f
C124 B.n84 VSUBS 0.006308f
C125 B.n85 VSUBS 0.006308f
C126 B.n86 VSUBS 0.006308f
C127 B.n87 VSUBS 0.006308f
C128 B.n88 VSUBS 0.006308f
C129 B.n89 VSUBS 0.006308f
C130 B.n90 VSUBS 0.006308f
C131 B.n91 VSUBS 0.006308f
C132 B.n92 VSUBS 0.006308f
C133 B.n93 VSUBS 0.006308f
C134 B.n94 VSUBS 0.016025f
C135 B.n95 VSUBS 0.006308f
C136 B.n96 VSUBS 0.006308f
C137 B.n97 VSUBS 0.006308f
C138 B.n98 VSUBS 0.006308f
C139 B.n99 VSUBS 0.006308f
C140 B.n100 VSUBS 0.006308f
C141 B.n101 VSUBS 0.006308f
C142 B.n102 VSUBS 0.006308f
C143 B.n103 VSUBS 0.006308f
C144 B.n104 VSUBS 0.006308f
C145 B.n105 VSUBS 0.006308f
C146 B.n106 VSUBS 0.006308f
C147 B.n107 VSUBS 0.006308f
C148 B.n108 VSUBS 0.006308f
C149 B.n109 VSUBS 0.006308f
C150 B.n110 VSUBS 0.006308f
C151 B.n111 VSUBS 0.006308f
C152 B.n112 VSUBS 0.006308f
C153 B.n113 VSUBS 0.006308f
C154 B.n114 VSUBS 0.006308f
C155 B.n115 VSUBS 0.006308f
C156 B.n116 VSUBS 0.006308f
C157 B.n117 VSUBS 0.006308f
C158 B.n118 VSUBS 0.006308f
C159 B.n119 VSUBS 0.015514f
C160 B.n120 VSUBS 0.015514f
C161 B.n121 VSUBS 0.016025f
C162 B.n122 VSUBS 0.006308f
C163 B.n123 VSUBS 0.006308f
C164 B.n124 VSUBS 0.006308f
C165 B.n125 VSUBS 0.006308f
C166 B.n126 VSUBS 0.006308f
C167 B.n127 VSUBS 0.006308f
C168 B.n128 VSUBS 0.006308f
C169 B.n129 VSUBS 0.006308f
C170 B.n130 VSUBS 0.006308f
C171 B.n131 VSUBS 0.006308f
C172 B.n132 VSUBS 0.006308f
C173 B.n133 VSUBS 0.006308f
C174 B.n134 VSUBS 0.006308f
C175 B.n135 VSUBS 0.006308f
C176 B.n136 VSUBS 0.006308f
C177 B.n137 VSUBS 0.006308f
C178 B.n138 VSUBS 0.006308f
C179 B.n139 VSUBS 0.006308f
C180 B.n140 VSUBS 0.006308f
C181 B.n141 VSUBS 0.006308f
C182 B.n142 VSUBS 0.006308f
C183 B.n143 VSUBS 0.006308f
C184 B.n144 VSUBS 0.006308f
C185 B.n145 VSUBS 0.006308f
C186 B.n146 VSUBS 0.006308f
C187 B.n147 VSUBS 0.006308f
C188 B.n148 VSUBS 0.006308f
C189 B.n149 VSUBS 0.006308f
C190 B.n150 VSUBS 0.006308f
C191 B.n151 VSUBS 0.006308f
C192 B.n152 VSUBS 0.006308f
C193 B.n153 VSUBS 0.006308f
C194 B.n154 VSUBS 0.006308f
C195 B.n155 VSUBS 0.006308f
C196 B.n156 VSUBS 0.006308f
C197 B.n157 VSUBS 0.006308f
C198 B.n158 VSUBS 0.006308f
C199 B.n159 VSUBS 0.005751f
C200 B.n160 VSUBS 0.014614f
C201 B.n161 VSUBS 0.00371f
C202 B.n162 VSUBS 0.006308f
C203 B.n163 VSUBS 0.006308f
C204 B.n164 VSUBS 0.006308f
C205 B.n165 VSUBS 0.006308f
C206 B.n166 VSUBS 0.006308f
C207 B.n167 VSUBS 0.006308f
C208 B.n168 VSUBS 0.006308f
C209 B.n169 VSUBS 0.006308f
C210 B.n170 VSUBS 0.006308f
C211 B.n171 VSUBS 0.006308f
C212 B.n172 VSUBS 0.006308f
C213 B.n173 VSUBS 0.006308f
C214 B.n174 VSUBS 0.00371f
C215 B.n175 VSUBS 0.006308f
C216 B.n176 VSUBS 0.006308f
C217 B.n177 VSUBS 0.005751f
C218 B.n178 VSUBS 0.006308f
C219 B.n179 VSUBS 0.006308f
C220 B.n180 VSUBS 0.006308f
C221 B.n181 VSUBS 0.006308f
C222 B.n182 VSUBS 0.006308f
C223 B.n183 VSUBS 0.006308f
C224 B.n184 VSUBS 0.006308f
C225 B.n185 VSUBS 0.006308f
C226 B.n186 VSUBS 0.006308f
C227 B.n187 VSUBS 0.006308f
C228 B.n188 VSUBS 0.006308f
C229 B.n189 VSUBS 0.006308f
C230 B.n190 VSUBS 0.006308f
C231 B.n191 VSUBS 0.006308f
C232 B.n192 VSUBS 0.006308f
C233 B.n193 VSUBS 0.006308f
C234 B.n194 VSUBS 0.006308f
C235 B.n195 VSUBS 0.006308f
C236 B.n196 VSUBS 0.006308f
C237 B.n197 VSUBS 0.006308f
C238 B.n198 VSUBS 0.006308f
C239 B.n199 VSUBS 0.006308f
C240 B.n200 VSUBS 0.006308f
C241 B.n201 VSUBS 0.006308f
C242 B.n202 VSUBS 0.006308f
C243 B.n203 VSUBS 0.006308f
C244 B.n204 VSUBS 0.006308f
C245 B.n205 VSUBS 0.006308f
C246 B.n206 VSUBS 0.006308f
C247 B.n207 VSUBS 0.006308f
C248 B.n208 VSUBS 0.006308f
C249 B.n209 VSUBS 0.006308f
C250 B.n210 VSUBS 0.006308f
C251 B.n211 VSUBS 0.006308f
C252 B.n212 VSUBS 0.006308f
C253 B.n213 VSUBS 0.006308f
C254 B.n214 VSUBS 0.016025f
C255 B.n215 VSUBS 0.015514f
C256 B.n216 VSUBS 0.015514f
C257 B.n217 VSUBS 0.006308f
C258 B.n218 VSUBS 0.006308f
C259 B.n219 VSUBS 0.006308f
C260 B.n220 VSUBS 0.006308f
C261 B.n221 VSUBS 0.006308f
C262 B.n222 VSUBS 0.006308f
C263 B.n223 VSUBS 0.006308f
C264 B.n224 VSUBS 0.006308f
C265 B.n225 VSUBS 0.006308f
C266 B.n226 VSUBS 0.006308f
C267 B.n227 VSUBS 0.006308f
C268 B.n228 VSUBS 0.006308f
C269 B.n229 VSUBS 0.006308f
C270 B.n230 VSUBS 0.006308f
C271 B.n231 VSUBS 0.006308f
C272 B.n232 VSUBS 0.006308f
C273 B.n233 VSUBS 0.006308f
C274 B.n234 VSUBS 0.006308f
C275 B.n235 VSUBS 0.006308f
C276 B.n236 VSUBS 0.006308f
C277 B.n237 VSUBS 0.006308f
C278 B.n238 VSUBS 0.006308f
C279 B.n239 VSUBS 0.006308f
C280 B.n240 VSUBS 0.006308f
C281 B.n241 VSUBS 0.006308f
C282 B.n242 VSUBS 0.006308f
C283 B.n243 VSUBS 0.006308f
C284 B.n244 VSUBS 0.006308f
C285 B.n245 VSUBS 0.006308f
C286 B.n246 VSUBS 0.006308f
C287 B.n247 VSUBS 0.006308f
C288 B.n248 VSUBS 0.006308f
C289 B.n249 VSUBS 0.006308f
C290 B.n250 VSUBS 0.006308f
C291 B.n251 VSUBS 0.006308f
C292 B.n252 VSUBS 0.006308f
C293 B.n253 VSUBS 0.006308f
C294 B.n254 VSUBS 0.006308f
C295 B.n255 VSUBS 0.006308f
C296 B.n256 VSUBS 0.006308f
C297 B.n257 VSUBS 0.016189f
C298 B.n258 VSUBS 0.015514f
C299 B.n259 VSUBS 0.016025f
C300 B.n260 VSUBS 0.006308f
C301 B.n261 VSUBS 0.006308f
C302 B.n262 VSUBS 0.006308f
C303 B.n263 VSUBS 0.006308f
C304 B.n264 VSUBS 0.006308f
C305 B.n265 VSUBS 0.006308f
C306 B.n266 VSUBS 0.006308f
C307 B.n267 VSUBS 0.006308f
C308 B.n268 VSUBS 0.006308f
C309 B.n269 VSUBS 0.006308f
C310 B.n270 VSUBS 0.006308f
C311 B.n271 VSUBS 0.006308f
C312 B.n272 VSUBS 0.006308f
C313 B.n273 VSUBS 0.006308f
C314 B.n274 VSUBS 0.006308f
C315 B.n275 VSUBS 0.006308f
C316 B.n276 VSUBS 0.006308f
C317 B.n277 VSUBS 0.006308f
C318 B.n278 VSUBS 0.006308f
C319 B.n279 VSUBS 0.006308f
C320 B.n280 VSUBS 0.006308f
C321 B.n281 VSUBS 0.006308f
C322 B.n282 VSUBS 0.006308f
C323 B.n283 VSUBS 0.006308f
C324 B.n284 VSUBS 0.006308f
C325 B.n285 VSUBS 0.006308f
C326 B.n286 VSUBS 0.006308f
C327 B.n287 VSUBS 0.006308f
C328 B.n288 VSUBS 0.006308f
C329 B.n289 VSUBS 0.006308f
C330 B.n290 VSUBS 0.006308f
C331 B.n291 VSUBS 0.006308f
C332 B.n292 VSUBS 0.006308f
C333 B.n293 VSUBS 0.006308f
C334 B.n294 VSUBS 0.006308f
C335 B.n295 VSUBS 0.006308f
C336 B.n296 VSUBS 0.006308f
C337 B.n297 VSUBS 0.005751f
C338 B.n298 VSUBS 0.014614f
C339 B.n299 VSUBS 0.00371f
C340 B.n300 VSUBS 0.006308f
C341 B.n301 VSUBS 0.006308f
C342 B.n302 VSUBS 0.006308f
C343 B.n303 VSUBS 0.006308f
C344 B.n304 VSUBS 0.006308f
C345 B.n305 VSUBS 0.006308f
C346 B.n306 VSUBS 0.006308f
C347 B.n307 VSUBS 0.006308f
C348 B.n308 VSUBS 0.006308f
C349 B.n309 VSUBS 0.006308f
C350 B.n310 VSUBS 0.006308f
C351 B.n311 VSUBS 0.006308f
C352 B.n312 VSUBS 0.00371f
C353 B.n313 VSUBS 0.006308f
C354 B.n314 VSUBS 0.006308f
C355 B.n315 VSUBS 0.005751f
C356 B.n316 VSUBS 0.006308f
C357 B.n317 VSUBS 0.006308f
C358 B.n318 VSUBS 0.006308f
C359 B.n319 VSUBS 0.006308f
C360 B.n320 VSUBS 0.006308f
C361 B.n321 VSUBS 0.006308f
C362 B.n322 VSUBS 0.006308f
C363 B.n323 VSUBS 0.006308f
C364 B.n324 VSUBS 0.006308f
C365 B.n325 VSUBS 0.006308f
C366 B.n326 VSUBS 0.006308f
C367 B.n327 VSUBS 0.006308f
C368 B.n328 VSUBS 0.006308f
C369 B.n329 VSUBS 0.006308f
C370 B.n330 VSUBS 0.006308f
C371 B.n331 VSUBS 0.006308f
C372 B.n332 VSUBS 0.006308f
C373 B.n333 VSUBS 0.006308f
C374 B.n334 VSUBS 0.006308f
C375 B.n335 VSUBS 0.006308f
C376 B.n336 VSUBS 0.006308f
C377 B.n337 VSUBS 0.006308f
C378 B.n338 VSUBS 0.006308f
C379 B.n339 VSUBS 0.006308f
C380 B.n340 VSUBS 0.006308f
C381 B.n341 VSUBS 0.006308f
C382 B.n342 VSUBS 0.006308f
C383 B.n343 VSUBS 0.006308f
C384 B.n344 VSUBS 0.006308f
C385 B.n345 VSUBS 0.006308f
C386 B.n346 VSUBS 0.006308f
C387 B.n347 VSUBS 0.006308f
C388 B.n348 VSUBS 0.006308f
C389 B.n349 VSUBS 0.006308f
C390 B.n350 VSUBS 0.006308f
C391 B.n351 VSUBS 0.006308f
C392 B.n352 VSUBS 0.016025f
C393 B.n353 VSUBS 0.015514f
C394 B.n354 VSUBS 0.015514f
C395 B.n355 VSUBS 0.006308f
C396 B.n356 VSUBS 0.006308f
C397 B.n357 VSUBS 0.006308f
C398 B.n358 VSUBS 0.006308f
C399 B.n359 VSUBS 0.006308f
C400 B.n360 VSUBS 0.006308f
C401 B.n361 VSUBS 0.006308f
C402 B.n362 VSUBS 0.006308f
C403 B.n363 VSUBS 0.006308f
C404 B.n364 VSUBS 0.006308f
C405 B.n365 VSUBS 0.006308f
C406 B.n366 VSUBS 0.006308f
C407 B.n367 VSUBS 0.006308f
C408 B.n368 VSUBS 0.006308f
C409 B.n369 VSUBS 0.006308f
C410 B.n370 VSUBS 0.006308f
C411 B.n371 VSUBS 0.006308f
C412 B.n372 VSUBS 0.006308f
C413 B.n373 VSUBS 0.006308f
C414 B.n374 VSUBS 0.006308f
C415 B.n375 VSUBS 0.014283f
C416 VDD1.t1 VSUBS 0.788583f
C417 VDD1.t0 VSUBS 1.03074f
C418 VP.t0 VSUBS 0.642208f
C419 VP.t1 VSUBS 0.553234f
C420 VP.n0 VSUBS 2.39249f
C421 VDD2.t1 VSUBS 1.03256f
C422 VDD2.t0 VSUBS 0.799918f
C423 VDD2.n0 VSUBS 1.93f
C424 VTAIL.t1 VSUBS 1.04038f
C425 VTAIL.n0 VSUBS 1.40493f
C426 VTAIL.t2 VSUBS 1.04039f
C427 VTAIL.n1 VSUBS 1.41674f
C428 VTAIL.t0 VSUBS 1.04038f
C429 VTAIL.n2 VSUBS 1.35249f
C430 VTAIL.t3 VSUBS 1.04038f
C431 VTAIL.n3 VSUBS 1.29784f
C432 VN.t0 VSUBS 0.54574f
C433 VN.t1 VSUBS 0.636042f
.ends

