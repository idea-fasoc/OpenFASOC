* NGSPICE file created from diff_pair_sample_0435.ext - technology: sky130A

.subckt diff_pair_sample_0435 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 w_n1678_n3640# sky130_fd_pr__pfet_01v8 ad=5.2104 pd=27.5 as=5.2104 ps=27.5 w=13.36 l=1.44
X1 VDD1.t0 VP.t1 VTAIL.t2 w_n1678_n3640# sky130_fd_pr__pfet_01v8 ad=5.2104 pd=27.5 as=5.2104 ps=27.5 w=13.36 l=1.44
X2 VDD2.t1 VN.t0 VTAIL.t1 w_n1678_n3640# sky130_fd_pr__pfet_01v8 ad=5.2104 pd=27.5 as=5.2104 ps=27.5 w=13.36 l=1.44
X3 VDD2.t0 VN.t1 VTAIL.t0 w_n1678_n3640# sky130_fd_pr__pfet_01v8 ad=5.2104 pd=27.5 as=5.2104 ps=27.5 w=13.36 l=1.44
X4 B.t11 B.t9 B.t10 w_n1678_n3640# sky130_fd_pr__pfet_01v8 ad=5.2104 pd=27.5 as=0 ps=0 w=13.36 l=1.44
X5 B.t8 B.t6 B.t7 w_n1678_n3640# sky130_fd_pr__pfet_01v8 ad=5.2104 pd=27.5 as=0 ps=0 w=13.36 l=1.44
X6 B.t5 B.t3 B.t4 w_n1678_n3640# sky130_fd_pr__pfet_01v8 ad=5.2104 pd=27.5 as=0 ps=0 w=13.36 l=1.44
X7 B.t2 B.t0 B.t1 w_n1678_n3640# sky130_fd_pr__pfet_01v8 ad=5.2104 pd=27.5 as=0 ps=0 w=13.36 l=1.44
R0 VP.n0 VP.t0 374.089
R1 VP.n0 VP.t1 331.478
R2 VP VP.n0 0.146778
R3 VTAIL.n241 VTAIL.n240 585
R4 VTAIL.n243 VTAIL.n242 585
R5 VTAIL.n236 VTAIL.n235 585
R6 VTAIL.n249 VTAIL.n248 585
R7 VTAIL.n251 VTAIL.n250 585
R8 VTAIL.n232 VTAIL.n231 585
R9 VTAIL.n257 VTAIL.n256 585
R10 VTAIL.n259 VTAIL.n258 585
R11 VTAIL.n228 VTAIL.n227 585
R12 VTAIL.n265 VTAIL.n264 585
R13 VTAIL.n267 VTAIL.n266 585
R14 VTAIL.n224 VTAIL.n223 585
R15 VTAIL.n273 VTAIL.n272 585
R16 VTAIL.n275 VTAIL.n274 585
R17 VTAIL.n220 VTAIL.n219 585
R18 VTAIL.n281 VTAIL.n280 585
R19 VTAIL.n283 VTAIL.n282 585
R20 VTAIL.n25 VTAIL.n24 585
R21 VTAIL.n27 VTAIL.n26 585
R22 VTAIL.n20 VTAIL.n19 585
R23 VTAIL.n33 VTAIL.n32 585
R24 VTAIL.n35 VTAIL.n34 585
R25 VTAIL.n16 VTAIL.n15 585
R26 VTAIL.n41 VTAIL.n40 585
R27 VTAIL.n43 VTAIL.n42 585
R28 VTAIL.n12 VTAIL.n11 585
R29 VTAIL.n49 VTAIL.n48 585
R30 VTAIL.n51 VTAIL.n50 585
R31 VTAIL.n8 VTAIL.n7 585
R32 VTAIL.n57 VTAIL.n56 585
R33 VTAIL.n59 VTAIL.n58 585
R34 VTAIL.n4 VTAIL.n3 585
R35 VTAIL.n65 VTAIL.n64 585
R36 VTAIL.n67 VTAIL.n66 585
R37 VTAIL.n211 VTAIL.n210 585
R38 VTAIL.n209 VTAIL.n208 585
R39 VTAIL.n148 VTAIL.n147 585
R40 VTAIL.n203 VTAIL.n202 585
R41 VTAIL.n201 VTAIL.n200 585
R42 VTAIL.n152 VTAIL.n151 585
R43 VTAIL.n195 VTAIL.n194 585
R44 VTAIL.n193 VTAIL.n192 585
R45 VTAIL.n156 VTAIL.n155 585
R46 VTAIL.n187 VTAIL.n186 585
R47 VTAIL.n185 VTAIL.n184 585
R48 VTAIL.n160 VTAIL.n159 585
R49 VTAIL.n179 VTAIL.n178 585
R50 VTAIL.n177 VTAIL.n176 585
R51 VTAIL.n164 VTAIL.n163 585
R52 VTAIL.n171 VTAIL.n170 585
R53 VTAIL.n169 VTAIL.n168 585
R54 VTAIL.n139 VTAIL.n138 585
R55 VTAIL.n137 VTAIL.n136 585
R56 VTAIL.n76 VTAIL.n75 585
R57 VTAIL.n131 VTAIL.n130 585
R58 VTAIL.n129 VTAIL.n128 585
R59 VTAIL.n80 VTAIL.n79 585
R60 VTAIL.n123 VTAIL.n122 585
R61 VTAIL.n121 VTAIL.n120 585
R62 VTAIL.n84 VTAIL.n83 585
R63 VTAIL.n115 VTAIL.n114 585
R64 VTAIL.n113 VTAIL.n112 585
R65 VTAIL.n88 VTAIL.n87 585
R66 VTAIL.n107 VTAIL.n106 585
R67 VTAIL.n105 VTAIL.n104 585
R68 VTAIL.n92 VTAIL.n91 585
R69 VTAIL.n99 VTAIL.n98 585
R70 VTAIL.n97 VTAIL.n96 585
R71 VTAIL.n282 VTAIL.n216 498.474
R72 VTAIL.n66 VTAIL.n0 498.474
R73 VTAIL.n210 VTAIL.n144 498.474
R74 VTAIL.n138 VTAIL.n72 498.474
R75 VTAIL.n239 VTAIL.t0 327.466
R76 VTAIL.n23 VTAIL.t2 327.466
R77 VTAIL.n167 VTAIL.t3 327.466
R78 VTAIL.n95 VTAIL.t1 327.466
R79 VTAIL.n242 VTAIL.n241 171.744
R80 VTAIL.n242 VTAIL.n235 171.744
R81 VTAIL.n249 VTAIL.n235 171.744
R82 VTAIL.n250 VTAIL.n249 171.744
R83 VTAIL.n250 VTAIL.n231 171.744
R84 VTAIL.n257 VTAIL.n231 171.744
R85 VTAIL.n258 VTAIL.n257 171.744
R86 VTAIL.n258 VTAIL.n227 171.744
R87 VTAIL.n265 VTAIL.n227 171.744
R88 VTAIL.n266 VTAIL.n265 171.744
R89 VTAIL.n266 VTAIL.n223 171.744
R90 VTAIL.n273 VTAIL.n223 171.744
R91 VTAIL.n274 VTAIL.n273 171.744
R92 VTAIL.n274 VTAIL.n219 171.744
R93 VTAIL.n281 VTAIL.n219 171.744
R94 VTAIL.n282 VTAIL.n281 171.744
R95 VTAIL.n26 VTAIL.n25 171.744
R96 VTAIL.n26 VTAIL.n19 171.744
R97 VTAIL.n33 VTAIL.n19 171.744
R98 VTAIL.n34 VTAIL.n33 171.744
R99 VTAIL.n34 VTAIL.n15 171.744
R100 VTAIL.n41 VTAIL.n15 171.744
R101 VTAIL.n42 VTAIL.n41 171.744
R102 VTAIL.n42 VTAIL.n11 171.744
R103 VTAIL.n49 VTAIL.n11 171.744
R104 VTAIL.n50 VTAIL.n49 171.744
R105 VTAIL.n50 VTAIL.n7 171.744
R106 VTAIL.n57 VTAIL.n7 171.744
R107 VTAIL.n58 VTAIL.n57 171.744
R108 VTAIL.n58 VTAIL.n3 171.744
R109 VTAIL.n65 VTAIL.n3 171.744
R110 VTAIL.n66 VTAIL.n65 171.744
R111 VTAIL.n210 VTAIL.n209 171.744
R112 VTAIL.n209 VTAIL.n147 171.744
R113 VTAIL.n202 VTAIL.n147 171.744
R114 VTAIL.n202 VTAIL.n201 171.744
R115 VTAIL.n201 VTAIL.n151 171.744
R116 VTAIL.n194 VTAIL.n151 171.744
R117 VTAIL.n194 VTAIL.n193 171.744
R118 VTAIL.n193 VTAIL.n155 171.744
R119 VTAIL.n186 VTAIL.n155 171.744
R120 VTAIL.n186 VTAIL.n185 171.744
R121 VTAIL.n185 VTAIL.n159 171.744
R122 VTAIL.n178 VTAIL.n159 171.744
R123 VTAIL.n178 VTAIL.n177 171.744
R124 VTAIL.n177 VTAIL.n163 171.744
R125 VTAIL.n170 VTAIL.n163 171.744
R126 VTAIL.n170 VTAIL.n169 171.744
R127 VTAIL.n138 VTAIL.n137 171.744
R128 VTAIL.n137 VTAIL.n75 171.744
R129 VTAIL.n130 VTAIL.n75 171.744
R130 VTAIL.n130 VTAIL.n129 171.744
R131 VTAIL.n129 VTAIL.n79 171.744
R132 VTAIL.n122 VTAIL.n79 171.744
R133 VTAIL.n122 VTAIL.n121 171.744
R134 VTAIL.n121 VTAIL.n83 171.744
R135 VTAIL.n114 VTAIL.n83 171.744
R136 VTAIL.n114 VTAIL.n113 171.744
R137 VTAIL.n113 VTAIL.n87 171.744
R138 VTAIL.n106 VTAIL.n87 171.744
R139 VTAIL.n106 VTAIL.n105 171.744
R140 VTAIL.n105 VTAIL.n91 171.744
R141 VTAIL.n98 VTAIL.n91 171.744
R142 VTAIL.n98 VTAIL.n97 171.744
R143 VTAIL.n241 VTAIL.t0 85.8723
R144 VTAIL.n25 VTAIL.t2 85.8723
R145 VTAIL.n169 VTAIL.t3 85.8723
R146 VTAIL.n97 VTAIL.t1 85.8723
R147 VTAIL.n287 VTAIL.n286 35.2884
R148 VTAIL.n71 VTAIL.n70 35.2884
R149 VTAIL.n215 VTAIL.n214 35.2884
R150 VTAIL.n143 VTAIL.n142 35.2884
R151 VTAIL.n143 VTAIL.n71 26.9358
R152 VTAIL.n287 VTAIL.n215 25.41
R153 VTAIL.n240 VTAIL.n239 16.3895
R154 VTAIL.n24 VTAIL.n23 16.3895
R155 VTAIL.n168 VTAIL.n167 16.3895
R156 VTAIL.n96 VTAIL.n95 16.3895
R157 VTAIL.n243 VTAIL.n238 12.8005
R158 VTAIL.n284 VTAIL.n283 12.8005
R159 VTAIL.n27 VTAIL.n22 12.8005
R160 VTAIL.n68 VTAIL.n67 12.8005
R161 VTAIL.n212 VTAIL.n211 12.8005
R162 VTAIL.n171 VTAIL.n166 12.8005
R163 VTAIL.n140 VTAIL.n139 12.8005
R164 VTAIL.n99 VTAIL.n94 12.8005
R165 VTAIL.n244 VTAIL.n236 12.0247
R166 VTAIL.n280 VTAIL.n218 12.0247
R167 VTAIL.n28 VTAIL.n20 12.0247
R168 VTAIL.n64 VTAIL.n2 12.0247
R169 VTAIL.n208 VTAIL.n146 12.0247
R170 VTAIL.n172 VTAIL.n164 12.0247
R171 VTAIL.n136 VTAIL.n74 12.0247
R172 VTAIL.n100 VTAIL.n92 12.0247
R173 VTAIL.n248 VTAIL.n247 11.249
R174 VTAIL.n279 VTAIL.n220 11.249
R175 VTAIL.n32 VTAIL.n31 11.249
R176 VTAIL.n63 VTAIL.n4 11.249
R177 VTAIL.n207 VTAIL.n148 11.249
R178 VTAIL.n176 VTAIL.n175 11.249
R179 VTAIL.n135 VTAIL.n76 11.249
R180 VTAIL.n104 VTAIL.n103 11.249
R181 VTAIL.n251 VTAIL.n234 10.4732
R182 VTAIL.n276 VTAIL.n275 10.4732
R183 VTAIL.n35 VTAIL.n18 10.4732
R184 VTAIL.n60 VTAIL.n59 10.4732
R185 VTAIL.n204 VTAIL.n203 10.4732
R186 VTAIL.n179 VTAIL.n162 10.4732
R187 VTAIL.n132 VTAIL.n131 10.4732
R188 VTAIL.n107 VTAIL.n90 10.4732
R189 VTAIL.n252 VTAIL.n232 9.69747
R190 VTAIL.n272 VTAIL.n222 9.69747
R191 VTAIL.n36 VTAIL.n16 9.69747
R192 VTAIL.n56 VTAIL.n6 9.69747
R193 VTAIL.n200 VTAIL.n150 9.69747
R194 VTAIL.n180 VTAIL.n160 9.69747
R195 VTAIL.n128 VTAIL.n78 9.69747
R196 VTAIL.n108 VTAIL.n88 9.69747
R197 VTAIL.n286 VTAIL.n285 9.45567
R198 VTAIL.n70 VTAIL.n69 9.45567
R199 VTAIL.n214 VTAIL.n213 9.45567
R200 VTAIL.n142 VTAIL.n141 9.45567
R201 VTAIL.n261 VTAIL.n260 9.3005
R202 VTAIL.n230 VTAIL.n229 9.3005
R203 VTAIL.n255 VTAIL.n254 9.3005
R204 VTAIL.n253 VTAIL.n252 9.3005
R205 VTAIL.n234 VTAIL.n233 9.3005
R206 VTAIL.n247 VTAIL.n246 9.3005
R207 VTAIL.n245 VTAIL.n244 9.3005
R208 VTAIL.n238 VTAIL.n237 9.3005
R209 VTAIL.n263 VTAIL.n262 9.3005
R210 VTAIL.n226 VTAIL.n225 9.3005
R211 VTAIL.n269 VTAIL.n268 9.3005
R212 VTAIL.n271 VTAIL.n270 9.3005
R213 VTAIL.n222 VTAIL.n221 9.3005
R214 VTAIL.n277 VTAIL.n276 9.3005
R215 VTAIL.n279 VTAIL.n278 9.3005
R216 VTAIL.n218 VTAIL.n217 9.3005
R217 VTAIL.n285 VTAIL.n284 9.3005
R218 VTAIL.n45 VTAIL.n44 9.3005
R219 VTAIL.n14 VTAIL.n13 9.3005
R220 VTAIL.n39 VTAIL.n38 9.3005
R221 VTAIL.n37 VTAIL.n36 9.3005
R222 VTAIL.n18 VTAIL.n17 9.3005
R223 VTAIL.n31 VTAIL.n30 9.3005
R224 VTAIL.n29 VTAIL.n28 9.3005
R225 VTAIL.n22 VTAIL.n21 9.3005
R226 VTAIL.n47 VTAIL.n46 9.3005
R227 VTAIL.n10 VTAIL.n9 9.3005
R228 VTAIL.n53 VTAIL.n52 9.3005
R229 VTAIL.n55 VTAIL.n54 9.3005
R230 VTAIL.n6 VTAIL.n5 9.3005
R231 VTAIL.n61 VTAIL.n60 9.3005
R232 VTAIL.n63 VTAIL.n62 9.3005
R233 VTAIL.n2 VTAIL.n1 9.3005
R234 VTAIL.n69 VTAIL.n68 9.3005
R235 VTAIL.n154 VTAIL.n153 9.3005
R236 VTAIL.n197 VTAIL.n196 9.3005
R237 VTAIL.n199 VTAIL.n198 9.3005
R238 VTAIL.n150 VTAIL.n149 9.3005
R239 VTAIL.n205 VTAIL.n204 9.3005
R240 VTAIL.n207 VTAIL.n206 9.3005
R241 VTAIL.n146 VTAIL.n145 9.3005
R242 VTAIL.n213 VTAIL.n212 9.3005
R243 VTAIL.n191 VTAIL.n190 9.3005
R244 VTAIL.n189 VTAIL.n188 9.3005
R245 VTAIL.n158 VTAIL.n157 9.3005
R246 VTAIL.n183 VTAIL.n182 9.3005
R247 VTAIL.n181 VTAIL.n180 9.3005
R248 VTAIL.n162 VTAIL.n161 9.3005
R249 VTAIL.n175 VTAIL.n174 9.3005
R250 VTAIL.n173 VTAIL.n172 9.3005
R251 VTAIL.n166 VTAIL.n165 9.3005
R252 VTAIL.n82 VTAIL.n81 9.3005
R253 VTAIL.n125 VTAIL.n124 9.3005
R254 VTAIL.n127 VTAIL.n126 9.3005
R255 VTAIL.n78 VTAIL.n77 9.3005
R256 VTAIL.n133 VTAIL.n132 9.3005
R257 VTAIL.n135 VTAIL.n134 9.3005
R258 VTAIL.n74 VTAIL.n73 9.3005
R259 VTAIL.n141 VTAIL.n140 9.3005
R260 VTAIL.n119 VTAIL.n118 9.3005
R261 VTAIL.n117 VTAIL.n116 9.3005
R262 VTAIL.n86 VTAIL.n85 9.3005
R263 VTAIL.n111 VTAIL.n110 9.3005
R264 VTAIL.n109 VTAIL.n108 9.3005
R265 VTAIL.n90 VTAIL.n89 9.3005
R266 VTAIL.n103 VTAIL.n102 9.3005
R267 VTAIL.n101 VTAIL.n100 9.3005
R268 VTAIL.n94 VTAIL.n93 9.3005
R269 VTAIL.n256 VTAIL.n255 8.92171
R270 VTAIL.n271 VTAIL.n224 8.92171
R271 VTAIL.n40 VTAIL.n39 8.92171
R272 VTAIL.n55 VTAIL.n8 8.92171
R273 VTAIL.n199 VTAIL.n152 8.92171
R274 VTAIL.n184 VTAIL.n183 8.92171
R275 VTAIL.n127 VTAIL.n80 8.92171
R276 VTAIL.n112 VTAIL.n111 8.92171
R277 VTAIL.n259 VTAIL.n230 8.14595
R278 VTAIL.n268 VTAIL.n267 8.14595
R279 VTAIL.n43 VTAIL.n14 8.14595
R280 VTAIL.n52 VTAIL.n51 8.14595
R281 VTAIL.n196 VTAIL.n195 8.14595
R282 VTAIL.n187 VTAIL.n158 8.14595
R283 VTAIL.n124 VTAIL.n123 8.14595
R284 VTAIL.n115 VTAIL.n86 8.14595
R285 VTAIL.n286 VTAIL.n216 7.75445
R286 VTAIL.n70 VTAIL.n0 7.75445
R287 VTAIL.n214 VTAIL.n144 7.75445
R288 VTAIL.n142 VTAIL.n72 7.75445
R289 VTAIL.n260 VTAIL.n228 7.3702
R290 VTAIL.n264 VTAIL.n226 7.3702
R291 VTAIL.n44 VTAIL.n12 7.3702
R292 VTAIL.n48 VTAIL.n10 7.3702
R293 VTAIL.n192 VTAIL.n154 7.3702
R294 VTAIL.n188 VTAIL.n156 7.3702
R295 VTAIL.n120 VTAIL.n82 7.3702
R296 VTAIL.n116 VTAIL.n84 7.3702
R297 VTAIL.n263 VTAIL.n228 6.59444
R298 VTAIL.n264 VTAIL.n263 6.59444
R299 VTAIL.n47 VTAIL.n12 6.59444
R300 VTAIL.n48 VTAIL.n47 6.59444
R301 VTAIL.n192 VTAIL.n191 6.59444
R302 VTAIL.n191 VTAIL.n156 6.59444
R303 VTAIL.n120 VTAIL.n119 6.59444
R304 VTAIL.n119 VTAIL.n84 6.59444
R305 VTAIL.n284 VTAIL.n216 6.08283
R306 VTAIL.n68 VTAIL.n0 6.08283
R307 VTAIL.n212 VTAIL.n144 6.08283
R308 VTAIL.n140 VTAIL.n72 6.08283
R309 VTAIL.n260 VTAIL.n259 5.81868
R310 VTAIL.n267 VTAIL.n226 5.81868
R311 VTAIL.n44 VTAIL.n43 5.81868
R312 VTAIL.n51 VTAIL.n10 5.81868
R313 VTAIL.n195 VTAIL.n154 5.81868
R314 VTAIL.n188 VTAIL.n187 5.81868
R315 VTAIL.n123 VTAIL.n82 5.81868
R316 VTAIL.n116 VTAIL.n115 5.81868
R317 VTAIL.n256 VTAIL.n230 5.04292
R318 VTAIL.n268 VTAIL.n224 5.04292
R319 VTAIL.n40 VTAIL.n14 5.04292
R320 VTAIL.n52 VTAIL.n8 5.04292
R321 VTAIL.n196 VTAIL.n152 5.04292
R322 VTAIL.n184 VTAIL.n158 5.04292
R323 VTAIL.n124 VTAIL.n80 5.04292
R324 VTAIL.n112 VTAIL.n86 5.04292
R325 VTAIL.n255 VTAIL.n232 4.26717
R326 VTAIL.n272 VTAIL.n271 4.26717
R327 VTAIL.n39 VTAIL.n16 4.26717
R328 VTAIL.n56 VTAIL.n55 4.26717
R329 VTAIL.n200 VTAIL.n199 4.26717
R330 VTAIL.n183 VTAIL.n160 4.26717
R331 VTAIL.n128 VTAIL.n127 4.26717
R332 VTAIL.n111 VTAIL.n88 4.26717
R333 VTAIL.n239 VTAIL.n237 3.70982
R334 VTAIL.n23 VTAIL.n21 3.70982
R335 VTAIL.n167 VTAIL.n165 3.70982
R336 VTAIL.n95 VTAIL.n93 3.70982
R337 VTAIL.n252 VTAIL.n251 3.49141
R338 VTAIL.n275 VTAIL.n222 3.49141
R339 VTAIL.n36 VTAIL.n35 3.49141
R340 VTAIL.n59 VTAIL.n6 3.49141
R341 VTAIL.n203 VTAIL.n150 3.49141
R342 VTAIL.n180 VTAIL.n179 3.49141
R343 VTAIL.n131 VTAIL.n78 3.49141
R344 VTAIL.n108 VTAIL.n107 3.49141
R345 VTAIL.n248 VTAIL.n234 2.71565
R346 VTAIL.n276 VTAIL.n220 2.71565
R347 VTAIL.n32 VTAIL.n18 2.71565
R348 VTAIL.n60 VTAIL.n4 2.71565
R349 VTAIL.n204 VTAIL.n148 2.71565
R350 VTAIL.n176 VTAIL.n162 2.71565
R351 VTAIL.n132 VTAIL.n76 2.71565
R352 VTAIL.n104 VTAIL.n90 2.71565
R353 VTAIL.n247 VTAIL.n236 1.93989
R354 VTAIL.n280 VTAIL.n279 1.93989
R355 VTAIL.n31 VTAIL.n20 1.93989
R356 VTAIL.n64 VTAIL.n63 1.93989
R357 VTAIL.n208 VTAIL.n207 1.93989
R358 VTAIL.n175 VTAIL.n164 1.93989
R359 VTAIL.n136 VTAIL.n135 1.93989
R360 VTAIL.n103 VTAIL.n92 1.93989
R361 VTAIL.n215 VTAIL.n143 1.23326
R362 VTAIL.n244 VTAIL.n243 1.16414
R363 VTAIL.n283 VTAIL.n218 1.16414
R364 VTAIL.n28 VTAIL.n27 1.16414
R365 VTAIL.n67 VTAIL.n2 1.16414
R366 VTAIL.n211 VTAIL.n146 1.16414
R367 VTAIL.n172 VTAIL.n171 1.16414
R368 VTAIL.n139 VTAIL.n74 1.16414
R369 VTAIL.n100 VTAIL.n99 1.16414
R370 VTAIL VTAIL.n71 0.909983
R371 VTAIL.n240 VTAIL.n238 0.388379
R372 VTAIL.n24 VTAIL.n22 0.388379
R373 VTAIL.n168 VTAIL.n166 0.388379
R374 VTAIL.n96 VTAIL.n94 0.388379
R375 VTAIL VTAIL.n287 0.323776
R376 VTAIL.n245 VTAIL.n237 0.155672
R377 VTAIL.n246 VTAIL.n245 0.155672
R378 VTAIL.n246 VTAIL.n233 0.155672
R379 VTAIL.n253 VTAIL.n233 0.155672
R380 VTAIL.n254 VTAIL.n253 0.155672
R381 VTAIL.n254 VTAIL.n229 0.155672
R382 VTAIL.n261 VTAIL.n229 0.155672
R383 VTAIL.n262 VTAIL.n261 0.155672
R384 VTAIL.n262 VTAIL.n225 0.155672
R385 VTAIL.n269 VTAIL.n225 0.155672
R386 VTAIL.n270 VTAIL.n269 0.155672
R387 VTAIL.n270 VTAIL.n221 0.155672
R388 VTAIL.n277 VTAIL.n221 0.155672
R389 VTAIL.n278 VTAIL.n277 0.155672
R390 VTAIL.n278 VTAIL.n217 0.155672
R391 VTAIL.n285 VTAIL.n217 0.155672
R392 VTAIL.n29 VTAIL.n21 0.155672
R393 VTAIL.n30 VTAIL.n29 0.155672
R394 VTAIL.n30 VTAIL.n17 0.155672
R395 VTAIL.n37 VTAIL.n17 0.155672
R396 VTAIL.n38 VTAIL.n37 0.155672
R397 VTAIL.n38 VTAIL.n13 0.155672
R398 VTAIL.n45 VTAIL.n13 0.155672
R399 VTAIL.n46 VTAIL.n45 0.155672
R400 VTAIL.n46 VTAIL.n9 0.155672
R401 VTAIL.n53 VTAIL.n9 0.155672
R402 VTAIL.n54 VTAIL.n53 0.155672
R403 VTAIL.n54 VTAIL.n5 0.155672
R404 VTAIL.n61 VTAIL.n5 0.155672
R405 VTAIL.n62 VTAIL.n61 0.155672
R406 VTAIL.n62 VTAIL.n1 0.155672
R407 VTAIL.n69 VTAIL.n1 0.155672
R408 VTAIL.n213 VTAIL.n145 0.155672
R409 VTAIL.n206 VTAIL.n145 0.155672
R410 VTAIL.n206 VTAIL.n205 0.155672
R411 VTAIL.n205 VTAIL.n149 0.155672
R412 VTAIL.n198 VTAIL.n149 0.155672
R413 VTAIL.n198 VTAIL.n197 0.155672
R414 VTAIL.n197 VTAIL.n153 0.155672
R415 VTAIL.n190 VTAIL.n153 0.155672
R416 VTAIL.n190 VTAIL.n189 0.155672
R417 VTAIL.n189 VTAIL.n157 0.155672
R418 VTAIL.n182 VTAIL.n157 0.155672
R419 VTAIL.n182 VTAIL.n181 0.155672
R420 VTAIL.n181 VTAIL.n161 0.155672
R421 VTAIL.n174 VTAIL.n161 0.155672
R422 VTAIL.n174 VTAIL.n173 0.155672
R423 VTAIL.n173 VTAIL.n165 0.155672
R424 VTAIL.n141 VTAIL.n73 0.155672
R425 VTAIL.n134 VTAIL.n73 0.155672
R426 VTAIL.n134 VTAIL.n133 0.155672
R427 VTAIL.n133 VTAIL.n77 0.155672
R428 VTAIL.n126 VTAIL.n77 0.155672
R429 VTAIL.n126 VTAIL.n125 0.155672
R430 VTAIL.n125 VTAIL.n81 0.155672
R431 VTAIL.n118 VTAIL.n81 0.155672
R432 VTAIL.n118 VTAIL.n117 0.155672
R433 VTAIL.n117 VTAIL.n85 0.155672
R434 VTAIL.n110 VTAIL.n85 0.155672
R435 VTAIL.n110 VTAIL.n109 0.155672
R436 VTAIL.n109 VTAIL.n89 0.155672
R437 VTAIL.n102 VTAIL.n89 0.155672
R438 VTAIL.n102 VTAIL.n101 0.155672
R439 VTAIL.n101 VTAIL.n93 0.155672
R440 VDD1.n67 VDD1.n66 585
R441 VDD1.n65 VDD1.n64 585
R442 VDD1.n4 VDD1.n3 585
R443 VDD1.n59 VDD1.n58 585
R444 VDD1.n57 VDD1.n56 585
R445 VDD1.n8 VDD1.n7 585
R446 VDD1.n51 VDD1.n50 585
R447 VDD1.n49 VDD1.n48 585
R448 VDD1.n12 VDD1.n11 585
R449 VDD1.n43 VDD1.n42 585
R450 VDD1.n41 VDD1.n40 585
R451 VDD1.n16 VDD1.n15 585
R452 VDD1.n35 VDD1.n34 585
R453 VDD1.n33 VDD1.n32 585
R454 VDD1.n20 VDD1.n19 585
R455 VDD1.n27 VDD1.n26 585
R456 VDD1.n25 VDD1.n24 585
R457 VDD1.n96 VDD1.n95 585
R458 VDD1.n98 VDD1.n97 585
R459 VDD1.n91 VDD1.n90 585
R460 VDD1.n104 VDD1.n103 585
R461 VDD1.n106 VDD1.n105 585
R462 VDD1.n87 VDD1.n86 585
R463 VDD1.n112 VDD1.n111 585
R464 VDD1.n114 VDD1.n113 585
R465 VDD1.n83 VDD1.n82 585
R466 VDD1.n120 VDD1.n119 585
R467 VDD1.n122 VDD1.n121 585
R468 VDD1.n79 VDD1.n78 585
R469 VDD1.n128 VDD1.n127 585
R470 VDD1.n130 VDD1.n129 585
R471 VDD1.n75 VDD1.n74 585
R472 VDD1.n136 VDD1.n135 585
R473 VDD1.n138 VDD1.n137 585
R474 VDD1.n66 VDD1.n0 498.474
R475 VDD1.n137 VDD1.n71 498.474
R476 VDD1.n23 VDD1.t1 327.466
R477 VDD1.n94 VDD1.t0 327.466
R478 VDD1.n66 VDD1.n65 171.744
R479 VDD1.n65 VDD1.n3 171.744
R480 VDD1.n58 VDD1.n3 171.744
R481 VDD1.n58 VDD1.n57 171.744
R482 VDD1.n57 VDD1.n7 171.744
R483 VDD1.n50 VDD1.n7 171.744
R484 VDD1.n50 VDD1.n49 171.744
R485 VDD1.n49 VDD1.n11 171.744
R486 VDD1.n42 VDD1.n11 171.744
R487 VDD1.n42 VDD1.n41 171.744
R488 VDD1.n41 VDD1.n15 171.744
R489 VDD1.n34 VDD1.n15 171.744
R490 VDD1.n34 VDD1.n33 171.744
R491 VDD1.n33 VDD1.n19 171.744
R492 VDD1.n26 VDD1.n19 171.744
R493 VDD1.n26 VDD1.n25 171.744
R494 VDD1.n97 VDD1.n96 171.744
R495 VDD1.n97 VDD1.n90 171.744
R496 VDD1.n104 VDD1.n90 171.744
R497 VDD1.n105 VDD1.n104 171.744
R498 VDD1.n105 VDD1.n86 171.744
R499 VDD1.n112 VDD1.n86 171.744
R500 VDD1.n113 VDD1.n112 171.744
R501 VDD1.n113 VDD1.n82 171.744
R502 VDD1.n120 VDD1.n82 171.744
R503 VDD1.n121 VDD1.n120 171.744
R504 VDD1.n121 VDD1.n78 171.744
R505 VDD1.n128 VDD1.n78 171.744
R506 VDD1.n129 VDD1.n128 171.744
R507 VDD1.n129 VDD1.n74 171.744
R508 VDD1.n136 VDD1.n74 171.744
R509 VDD1.n137 VDD1.n136 171.744
R510 VDD1 VDD1.n141 91.1019
R511 VDD1.n25 VDD1.t1 85.8723
R512 VDD1.n96 VDD1.t0 85.8723
R513 VDD1 VDD1.n70 52.4068
R514 VDD1.n24 VDD1.n23 16.3895
R515 VDD1.n95 VDD1.n94 16.3895
R516 VDD1.n68 VDD1.n67 12.8005
R517 VDD1.n27 VDD1.n22 12.8005
R518 VDD1.n98 VDD1.n93 12.8005
R519 VDD1.n139 VDD1.n138 12.8005
R520 VDD1.n64 VDD1.n2 12.0247
R521 VDD1.n28 VDD1.n20 12.0247
R522 VDD1.n99 VDD1.n91 12.0247
R523 VDD1.n135 VDD1.n73 12.0247
R524 VDD1.n63 VDD1.n4 11.249
R525 VDD1.n32 VDD1.n31 11.249
R526 VDD1.n103 VDD1.n102 11.249
R527 VDD1.n134 VDD1.n75 11.249
R528 VDD1.n60 VDD1.n59 10.4732
R529 VDD1.n35 VDD1.n18 10.4732
R530 VDD1.n106 VDD1.n89 10.4732
R531 VDD1.n131 VDD1.n130 10.4732
R532 VDD1.n56 VDD1.n6 9.69747
R533 VDD1.n36 VDD1.n16 9.69747
R534 VDD1.n107 VDD1.n87 9.69747
R535 VDD1.n127 VDD1.n77 9.69747
R536 VDD1.n70 VDD1.n69 9.45567
R537 VDD1.n141 VDD1.n140 9.45567
R538 VDD1.n10 VDD1.n9 9.3005
R539 VDD1.n53 VDD1.n52 9.3005
R540 VDD1.n55 VDD1.n54 9.3005
R541 VDD1.n6 VDD1.n5 9.3005
R542 VDD1.n61 VDD1.n60 9.3005
R543 VDD1.n63 VDD1.n62 9.3005
R544 VDD1.n2 VDD1.n1 9.3005
R545 VDD1.n69 VDD1.n68 9.3005
R546 VDD1.n47 VDD1.n46 9.3005
R547 VDD1.n45 VDD1.n44 9.3005
R548 VDD1.n14 VDD1.n13 9.3005
R549 VDD1.n39 VDD1.n38 9.3005
R550 VDD1.n37 VDD1.n36 9.3005
R551 VDD1.n18 VDD1.n17 9.3005
R552 VDD1.n31 VDD1.n30 9.3005
R553 VDD1.n29 VDD1.n28 9.3005
R554 VDD1.n22 VDD1.n21 9.3005
R555 VDD1.n116 VDD1.n115 9.3005
R556 VDD1.n85 VDD1.n84 9.3005
R557 VDD1.n110 VDD1.n109 9.3005
R558 VDD1.n108 VDD1.n107 9.3005
R559 VDD1.n89 VDD1.n88 9.3005
R560 VDD1.n102 VDD1.n101 9.3005
R561 VDD1.n100 VDD1.n99 9.3005
R562 VDD1.n93 VDD1.n92 9.3005
R563 VDD1.n118 VDD1.n117 9.3005
R564 VDD1.n81 VDD1.n80 9.3005
R565 VDD1.n124 VDD1.n123 9.3005
R566 VDD1.n126 VDD1.n125 9.3005
R567 VDD1.n77 VDD1.n76 9.3005
R568 VDD1.n132 VDD1.n131 9.3005
R569 VDD1.n134 VDD1.n133 9.3005
R570 VDD1.n73 VDD1.n72 9.3005
R571 VDD1.n140 VDD1.n139 9.3005
R572 VDD1.n55 VDD1.n8 8.92171
R573 VDD1.n40 VDD1.n39 8.92171
R574 VDD1.n111 VDD1.n110 8.92171
R575 VDD1.n126 VDD1.n79 8.92171
R576 VDD1.n52 VDD1.n51 8.14595
R577 VDD1.n43 VDD1.n14 8.14595
R578 VDD1.n114 VDD1.n85 8.14595
R579 VDD1.n123 VDD1.n122 8.14595
R580 VDD1.n70 VDD1.n0 7.75445
R581 VDD1.n141 VDD1.n71 7.75445
R582 VDD1.n48 VDD1.n10 7.3702
R583 VDD1.n44 VDD1.n12 7.3702
R584 VDD1.n115 VDD1.n83 7.3702
R585 VDD1.n119 VDD1.n81 7.3702
R586 VDD1.n48 VDD1.n47 6.59444
R587 VDD1.n47 VDD1.n12 6.59444
R588 VDD1.n118 VDD1.n83 6.59444
R589 VDD1.n119 VDD1.n118 6.59444
R590 VDD1.n68 VDD1.n0 6.08283
R591 VDD1.n139 VDD1.n71 6.08283
R592 VDD1.n51 VDD1.n10 5.81868
R593 VDD1.n44 VDD1.n43 5.81868
R594 VDD1.n115 VDD1.n114 5.81868
R595 VDD1.n122 VDD1.n81 5.81868
R596 VDD1.n52 VDD1.n8 5.04292
R597 VDD1.n40 VDD1.n14 5.04292
R598 VDD1.n111 VDD1.n85 5.04292
R599 VDD1.n123 VDD1.n79 5.04292
R600 VDD1.n56 VDD1.n55 4.26717
R601 VDD1.n39 VDD1.n16 4.26717
R602 VDD1.n110 VDD1.n87 4.26717
R603 VDD1.n127 VDD1.n126 4.26717
R604 VDD1.n23 VDD1.n21 3.70982
R605 VDD1.n94 VDD1.n92 3.70982
R606 VDD1.n59 VDD1.n6 3.49141
R607 VDD1.n36 VDD1.n35 3.49141
R608 VDD1.n107 VDD1.n106 3.49141
R609 VDD1.n130 VDD1.n77 3.49141
R610 VDD1.n60 VDD1.n4 2.71565
R611 VDD1.n32 VDD1.n18 2.71565
R612 VDD1.n103 VDD1.n89 2.71565
R613 VDD1.n131 VDD1.n75 2.71565
R614 VDD1.n64 VDD1.n63 1.93989
R615 VDD1.n31 VDD1.n20 1.93989
R616 VDD1.n102 VDD1.n91 1.93989
R617 VDD1.n135 VDD1.n134 1.93989
R618 VDD1.n67 VDD1.n2 1.16414
R619 VDD1.n28 VDD1.n27 1.16414
R620 VDD1.n99 VDD1.n98 1.16414
R621 VDD1.n138 VDD1.n73 1.16414
R622 VDD1.n24 VDD1.n22 0.388379
R623 VDD1.n95 VDD1.n93 0.388379
R624 VDD1.n69 VDD1.n1 0.155672
R625 VDD1.n62 VDD1.n1 0.155672
R626 VDD1.n62 VDD1.n61 0.155672
R627 VDD1.n61 VDD1.n5 0.155672
R628 VDD1.n54 VDD1.n5 0.155672
R629 VDD1.n54 VDD1.n53 0.155672
R630 VDD1.n53 VDD1.n9 0.155672
R631 VDD1.n46 VDD1.n9 0.155672
R632 VDD1.n46 VDD1.n45 0.155672
R633 VDD1.n45 VDD1.n13 0.155672
R634 VDD1.n38 VDD1.n13 0.155672
R635 VDD1.n38 VDD1.n37 0.155672
R636 VDD1.n37 VDD1.n17 0.155672
R637 VDD1.n30 VDD1.n17 0.155672
R638 VDD1.n30 VDD1.n29 0.155672
R639 VDD1.n29 VDD1.n21 0.155672
R640 VDD1.n100 VDD1.n92 0.155672
R641 VDD1.n101 VDD1.n100 0.155672
R642 VDD1.n101 VDD1.n88 0.155672
R643 VDD1.n108 VDD1.n88 0.155672
R644 VDD1.n109 VDD1.n108 0.155672
R645 VDD1.n109 VDD1.n84 0.155672
R646 VDD1.n116 VDD1.n84 0.155672
R647 VDD1.n117 VDD1.n116 0.155672
R648 VDD1.n117 VDD1.n80 0.155672
R649 VDD1.n124 VDD1.n80 0.155672
R650 VDD1.n125 VDD1.n124 0.155672
R651 VDD1.n125 VDD1.n76 0.155672
R652 VDD1.n132 VDD1.n76 0.155672
R653 VDD1.n133 VDD1.n132 0.155672
R654 VDD1.n133 VDD1.n72 0.155672
R655 VDD1.n140 VDD1.n72 0.155672
R656 VN VN.t0 374.375
R657 VN VN.t1 331.625
R658 VDD2.n138 VDD2.n137 585
R659 VDD2.n136 VDD2.n135 585
R660 VDD2.n75 VDD2.n74 585
R661 VDD2.n130 VDD2.n129 585
R662 VDD2.n128 VDD2.n127 585
R663 VDD2.n79 VDD2.n78 585
R664 VDD2.n122 VDD2.n121 585
R665 VDD2.n120 VDD2.n119 585
R666 VDD2.n83 VDD2.n82 585
R667 VDD2.n114 VDD2.n113 585
R668 VDD2.n112 VDD2.n111 585
R669 VDD2.n87 VDD2.n86 585
R670 VDD2.n106 VDD2.n105 585
R671 VDD2.n104 VDD2.n103 585
R672 VDD2.n91 VDD2.n90 585
R673 VDD2.n98 VDD2.n97 585
R674 VDD2.n96 VDD2.n95 585
R675 VDD2.n25 VDD2.n24 585
R676 VDD2.n27 VDD2.n26 585
R677 VDD2.n20 VDD2.n19 585
R678 VDD2.n33 VDD2.n32 585
R679 VDD2.n35 VDD2.n34 585
R680 VDD2.n16 VDD2.n15 585
R681 VDD2.n41 VDD2.n40 585
R682 VDD2.n43 VDD2.n42 585
R683 VDD2.n12 VDD2.n11 585
R684 VDD2.n49 VDD2.n48 585
R685 VDD2.n51 VDD2.n50 585
R686 VDD2.n8 VDD2.n7 585
R687 VDD2.n57 VDD2.n56 585
R688 VDD2.n59 VDD2.n58 585
R689 VDD2.n4 VDD2.n3 585
R690 VDD2.n65 VDD2.n64 585
R691 VDD2.n67 VDD2.n66 585
R692 VDD2.n137 VDD2.n71 498.474
R693 VDD2.n66 VDD2.n0 498.474
R694 VDD2.n94 VDD2.t1 327.466
R695 VDD2.n23 VDD2.t0 327.466
R696 VDD2.n137 VDD2.n136 171.744
R697 VDD2.n136 VDD2.n74 171.744
R698 VDD2.n129 VDD2.n74 171.744
R699 VDD2.n129 VDD2.n128 171.744
R700 VDD2.n128 VDD2.n78 171.744
R701 VDD2.n121 VDD2.n78 171.744
R702 VDD2.n121 VDD2.n120 171.744
R703 VDD2.n120 VDD2.n82 171.744
R704 VDD2.n113 VDD2.n82 171.744
R705 VDD2.n113 VDD2.n112 171.744
R706 VDD2.n112 VDD2.n86 171.744
R707 VDD2.n105 VDD2.n86 171.744
R708 VDD2.n105 VDD2.n104 171.744
R709 VDD2.n104 VDD2.n90 171.744
R710 VDD2.n97 VDD2.n90 171.744
R711 VDD2.n97 VDD2.n96 171.744
R712 VDD2.n26 VDD2.n25 171.744
R713 VDD2.n26 VDD2.n19 171.744
R714 VDD2.n33 VDD2.n19 171.744
R715 VDD2.n34 VDD2.n33 171.744
R716 VDD2.n34 VDD2.n15 171.744
R717 VDD2.n41 VDD2.n15 171.744
R718 VDD2.n42 VDD2.n41 171.744
R719 VDD2.n42 VDD2.n11 171.744
R720 VDD2.n49 VDD2.n11 171.744
R721 VDD2.n50 VDD2.n49 171.744
R722 VDD2.n50 VDD2.n7 171.744
R723 VDD2.n57 VDD2.n7 171.744
R724 VDD2.n58 VDD2.n57 171.744
R725 VDD2.n58 VDD2.n3 171.744
R726 VDD2.n65 VDD2.n3 171.744
R727 VDD2.n66 VDD2.n65 171.744
R728 VDD2.n142 VDD2.n70 90.1956
R729 VDD2.n96 VDD2.t1 85.8723
R730 VDD2.n25 VDD2.t0 85.8723
R731 VDD2.n142 VDD2.n141 51.9672
R732 VDD2.n95 VDD2.n94 16.3895
R733 VDD2.n24 VDD2.n23 16.3895
R734 VDD2.n139 VDD2.n138 12.8005
R735 VDD2.n98 VDD2.n93 12.8005
R736 VDD2.n27 VDD2.n22 12.8005
R737 VDD2.n68 VDD2.n67 12.8005
R738 VDD2.n135 VDD2.n73 12.0247
R739 VDD2.n99 VDD2.n91 12.0247
R740 VDD2.n28 VDD2.n20 12.0247
R741 VDD2.n64 VDD2.n2 12.0247
R742 VDD2.n134 VDD2.n75 11.249
R743 VDD2.n103 VDD2.n102 11.249
R744 VDD2.n32 VDD2.n31 11.249
R745 VDD2.n63 VDD2.n4 11.249
R746 VDD2.n131 VDD2.n130 10.4732
R747 VDD2.n106 VDD2.n89 10.4732
R748 VDD2.n35 VDD2.n18 10.4732
R749 VDD2.n60 VDD2.n59 10.4732
R750 VDD2.n127 VDD2.n77 9.69747
R751 VDD2.n107 VDD2.n87 9.69747
R752 VDD2.n36 VDD2.n16 9.69747
R753 VDD2.n56 VDD2.n6 9.69747
R754 VDD2.n141 VDD2.n140 9.45567
R755 VDD2.n70 VDD2.n69 9.45567
R756 VDD2.n81 VDD2.n80 9.3005
R757 VDD2.n124 VDD2.n123 9.3005
R758 VDD2.n126 VDD2.n125 9.3005
R759 VDD2.n77 VDD2.n76 9.3005
R760 VDD2.n132 VDD2.n131 9.3005
R761 VDD2.n134 VDD2.n133 9.3005
R762 VDD2.n73 VDD2.n72 9.3005
R763 VDD2.n140 VDD2.n139 9.3005
R764 VDD2.n118 VDD2.n117 9.3005
R765 VDD2.n116 VDD2.n115 9.3005
R766 VDD2.n85 VDD2.n84 9.3005
R767 VDD2.n110 VDD2.n109 9.3005
R768 VDD2.n108 VDD2.n107 9.3005
R769 VDD2.n89 VDD2.n88 9.3005
R770 VDD2.n102 VDD2.n101 9.3005
R771 VDD2.n100 VDD2.n99 9.3005
R772 VDD2.n93 VDD2.n92 9.3005
R773 VDD2.n45 VDD2.n44 9.3005
R774 VDD2.n14 VDD2.n13 9.3005
R775 VDD2.n39 VDD2.n38 9.3005
R776 VDD2.n37 VDD2.n36 9.3005
R777 VDD2.n18 VDD2.n17 9.3005
R778 VDD2.n31 VDD2.n30 9.3005
R779 VDD2.n29 VDD2.n28 9.3005
R780 VDD2.n22 VDD2.n21 9.3005
R781 VDD2.n47 VDD2.n46 9.3005
R782 VDD2.n10 VDD2.n9 9.3005
R783 VDD2.n53 VDD2.n52 9.3005
R784 VDD2.n55 VDD2.n54 9.3005
R785 VDD2.n6 VDD2.n5 9.3005
R786 VDD2.n61 VDD2.n60 9.3005
R787 VDD2.n63 VDD2.n62 9.3005
R788 VDD2.n2 VDD2.n1 9.3005
R789 VDD2.n69 VDD2.n68 9.3005
R790 VDD2.n126 VDD2.n79 8.92171
R791 VDD2.n111 VDD2.n110 8.92171
R792 VDD2.n40 VDD2.n39 8.92171
R793 VDD2.n55 VDD2.n8 8.92171
R794 VDD2.n123 VDD2.n122 8.14595
R795 VDD2.n114 VDD2.n85 8.14595
R796 VDD2.n43 VDD2.n14 8.14595
R797 VDD2.n52 VDD2.n51 8.14595
R798 VDD2.n141 VDD2.n71 7.75445
R799 VDD2.n70 VDD2.n0 7.75445
R800 VDD2.n119 VDD2.n81 7.3702
R801 VDD2.n115 VDD2.n83 7.3702
R802 VDD2.n44 VDD2.n12 7.3702
R803 VDD2.n48 VDD2.n10 7.3702
R804 VDD2.n119 VDD2.n118 6.59444
R805 VDD2.n118 VDD2.n83 6.59444
R806 VDD2.n47 VDD2.n12 6.59444
R807 VDD2.n48 VDD2.n47 6.59444
R808 VDD2.n139 VDD2.n71 6.08283
R809 VDD2.n68 VDD2.n0 6.08283
R810 VDD2.n122 VDD2.n81 5.81868
R811 VDD2.n115 VDD2.n114 5.81868
R812 VDD2.n44 VDD2.n43 5.81868
R813 VDD2.n51 VDD2.n10 5.81868
R814 VDD2.n123 VDD2.n79 5.04292
R815 VDD2.n111 VDD2.n85 5.04292
R816 VDD2.n40 VDD2.n14 5.04292
R817 VDD2.n52 VDD2.n8 5.04292
R818 VDD2.n127 VDD2.n126 4.26717
R819 VDD2.n110 VDD2.n87 4.26717
R820 VDD2.n39 VDD2.n16 4.26717
R821 VDD2.n56 VDD2.n55 4.26717
R822 VDD2.n94 VDD2.n92 3.70982
R823 VDD2.n23 VDD2.n21 3.70982
R824 VDD2.n130 VDD2.n77 3.49141
R825 VDD2.n107 VDD2.n106 3.49141
R826 VDD2.n36 VDD2.n35 3.49141
R827 VDD2.n59 VDD2.n6 3.49141
R828 VDD2.n131 VDD2.n75 2.71565
R829 VDD2.n103 VDD2.n89 2.71565
R830 VDD2.n32 VDD2.n18 2.71565
R831 VDD2.n60 VDD2.n4 2.71565
R832 VDD2.n135 VDD2.n134 1.93989
R833 VDD2.n102 VDD2.n91 1.93989
R834 VDD2.n31 VDD2.n20 1.93989
R835 VDD2.n64 VDD2.n63 1.93989
R836 VDD2.n138 VDD2.n73 1.16414
R837 VDD2.n99 VDD2.n98 1.16414
R838 VDD2.n28 VDD2.n27 1.16414
R839 VDD2.n67 VDD2.n2 1.16414
R840 VDD2 VDD2.n142 0.440155
R841 VDD2.n95 VDD2.n93 0.388379
R842 VDD2.n24 VDD2.n22 0.388379
R843 VDD2.n140 VDD2.n72 0.155672
R844 VDD2.n133 VDD2.n72 0.155672
R845 VDD2.n133 VDD2.n132 0.155672
R846 VDD2.n132 VDD2.n76 0.155672
R847 VDD2.n125 VDD2.n76 0.155672
R848 VDD2.n125 VDD2.n124 0.155672
R849 VDD2.n124 VDD2.n80 0.155672
R850 VDD2.n117 VDD2.n80 0.155672
R851 VDD2.n117 VDD2.n116 0.155672
R852 VDD2.n116 VDD2.n84 0.155672
R853 VDD2.n109 VDD2.n84 0.155672
R854 VDD2.n109 VDD2.n108 0.155672
R855 VDD2.n108 VDD2.n88 0.155672
R856 VDD2.n101 VDD2.n88 0.155672
R857 VDD2.n101 VDD2.n100 0.155672
R858 VDD2.n100 VDD2.n92 0.155672
R859 VDD2.n29 VDD2.n21 0.155672
R860 VDD2.n30 VDD2.n29 0.155672
R861 VDD2.n30 VDD2.n17 0.155672
R862 VDD2.n37 VDD2.n17 0.155672
R863 VDD2.n38 VDD2.n37 0.155672
R864 VDD2.n38 VDD2.n13 0.155672
R865 VDD2.n45 VDD2.n13 0.155672
R866 VDD2.n46 VDD2.n45 0.155672
R867 VDD2.n46 VDD2.n9 0.155672
R868 VDD2.n53 VDD2.n9 0.155672
R869 VDD2.n54 VDD2.n53 0.155672
R870 VDD2.n54 VDD2.n5 0.155672
R871 VDD2.n61 VDD2.n5 0.155672
R872 VDD2.n62 VDD2.n61 0.155672
R873 VDD2.n62 VDD2.n1 0.155672
R874 VDD2.n69 VDD2.n1 0.155672
R875 B.n326 B.n85 585
R876 B.n325 B.n324 585
R877 B.n323 B.n86 585
R878 B.n322 B.n321 585
R879 B.n320 B.n87 585
R880 B.n319 B.n318 585
R881 B.n317 B.n88 585
R882 B.n316 B.n315 585
R883 B.n314 B.n89 585
R884 B.n313 B.n312 585
R885 B.n311 B.n90 585
R886 B.n310 B.n309 585
R887 B.n308 B.n91 585
R888 B.n307 B.n306 585
R889 B.n305 B.n92 585
R890 B.n304 B.n303 585
R891 B.n302 B.n93 585
R892 B.n301 B.n300 585
R893 B.n299 B.n94 585
R894 B.n298 B.n297 585
R895 B.n296 B.n95 585
R896 B.n295 B.n294 585
R897 B.n293 B.n96 585
R898 B.n292 B.n291 585
R899 B.n290 B.n97 585
R900 B.n289 B.n288 585
R901 B.n287 B.n98 585
R902 B.n286 B.n285 585
R903 B.n284 B.n99 585
R904 B.n283 B.n282 585
R905 B.n281 B.n100 585
R906 B.n280 B.n279 585
R907 B.n278 B.n101 585
R908 B.n277 B.n276 585
R909 B.n275 B.n102 585
R910 B.n274 B.n273 585
R911 B.n272 B.n103 585
R912 B.n271 B.n270 585
R913 B.n269 B.n104 585
R914 B.n268 B.n267 585
R915 B.n266 B.n105 585
R916 B.n265 B.n264 585
R917 B.n263 B.n106 585
R918 B.n262 B.n261 585
R919 B.n260 B.n107 585
R920 B.n259 B.n258 585
R921 B.n257 B.n256 585
R922 B.n255 B.n111 585
R923 B.n254 B.n253 585
R924 B.n252 B.n112 585
R925 B.n251 B.n250 585
R926 B.n249 B.n113 585
R927 B.n248 B.n247 585
R928 B.n246 B.n114 585
R929 B.n245 B.n244 585
R930 B.n242 B.n115 585
R931 B.n241 B.n240 585
R932 B.n239 B.n118 585
R933 B.n238 B.n237 585
R934 B.n236 B.n119 585
R935 B.n235 B.n234 585
R936 B.n233 B.n120 585
R937 B.n232 B.n231 585
R938 B.n230 B.n121 585
R939 B.n229 B.n228 585
R940 B.n227 B.n122 585
R941 B.n226 B.n225 585
R942 B.n224 B.n123 585
R943 B.n223 B.n222 585
R944 B.n221 B.n124 585
R945 B.n220 B.n219 585
R946 B.n218 B.n125 585
R947 B.n217 B.n216 585
R948 B.n215 B.n126 585
R949 B.n214 B.n213 585
R950 B.n212 B.n127 585
R951 B.n211 B.n210 585
R952 B.n209 B.n128 585
R953 B.n208 B.n207 585
R954 B.n206 B.n129 585
R955 B.n205 B.n204 585
R956 B.n203 B.n130 585
R957 B.n202 B.n201 585
R958 B.n200 B.n131 585
R959 B.n199 B.n198 585
R960 B.n197 B.n132 585
R961 B.n196 B.n195 585
R962 B.n194 B.n133 585
R963 B.n193 B.n192 585
R964 B.n191 B.n134 585
R965 B.n190 B.n189 585
R966 B.n188 B.n135 585
R967 B.n187 B.n186 585
R968 B.n185 B.n136 585
R969 B.n184 B.n183 585
R970 B.n182 B.n137 585
R971 B.n181 B.n180 585
R972 B.n179 B.n138 585
R973 B.n178 B.n177 585
R974 B.n176 B.n139 585
R975 B.n175 B.n174 585
R976 B.n328 B.n327 585
R977 B.n329 B.n84 585
R978 B.n331 B.n330 585
R979 B.n332 B.n83 585
R980 B.n334 B.n333 585
R981 B.n335 B.n82 585
R982 B.n337 B.n336 585
R983 B.n338 B.n81 585
R984 B.n340 B.n339 585
R985 B.n341 B.n80 585
R986 B.n343 B.n342 585
R987 B.n344 B.n79 585
R988 B.n346 B.n345 585
R989 B.n347 B.n78 585
R990 B.n349 B.n348 585
R991 B.n350 B.n77 585
R992 B.n352 B.n351 585
R993 B.n353 B.n76 585
R994 B.n355 B.n354 585
R995 B.n356 B.n75 585
R996 B.n358 B.n357 585
R997 B.n359 B.n74 585
R998 B.n361 B.n360 585
R999 B.n362 B.n73 585
R1000 B.n364 B.n363 585
R1001 B.n365 B.n72 585
R1002 B.n367 B.n366 585
R1003 B.n368 B.n71 585
R1004 B.n370 B.n369 585
R1005 B.n371 B.n70 585
R1006 B.n373 B.n372 585
R1007 B.n374 B.n69 585
R1008 B.n376 B.n375 585
R1009 B.n377 B.n68 585
R1010 B.n379 B.n378 585
R1011 B.n380 B.n67 585
R1012 B.n382 B.n381 585
R1013 B.n383 B.n66 585
R1014 B.n536 B.n11 585
R1015 B.n535 B.n534 585
R1016 B.n533 B.n12 585
R1017 B.n532 B.n531 585
R1018 B.n530 B.n13 585
R1019 B.n529 B.n528 585
R1020 B.n527 B.n14 585
R1021 B.n526 B.n525 585
R1022 B.n524 B.n15 585
R1023 B.n523 B.n522 585
R1024 B.n521 B.n16 585
R1025 B.n520 B.n519 585
R1026 B.n518 B.n17 585
R1027 B.n517 B.n516 585
R1028 B.n515 B.n18 585
R1029 B.n514 B.n513 585
R1030 B.n512 B.n19 585
R1031 B.n511 B.n510 585
R1032 B.n509 B.n20 585
R1033 B.n508 B.n507 585
R1034 B.n506 B.n21 585
R1035 B.n505 B.n504 585
R1036 B.n503 B.n22 585
R1037 B.n502 B.n501 585
R1038 B.n500 B.n23 585
R1039 B.n499 B.n498 585
R1040 B.n497 B.n24 585
R1041 B.n496 B.n495 585
R1042 B.n494 B.n25 585
R1043 B.n493 B.n492 585
R1044 B.n491 B.n26 585
R1045 B.n490 B.n489 585
R1046 B.n488 B.n27 585
R1047 B.n487 B.n486 585
R1048 B.n485 B.n28 585
R1049 B.n484 B.n483 585
R1050 B.n482 B.n29 585
R1051 B.n481 B.n480 585
R1052 B.n479 B.n30 585
R1053 B.n478 B.n477 585
R1054 B.n476 B.n31 585
R1055 B.n475 B.n474 585
R1056 B.n473 B.n32 585
R1057 B.n472 B.n471 585
R1058 B.n470 B.n33 585
R1059 B.n469 B.n468 585
R1060 B.n467 B.n466 585
R1061 B.n465 B.n37 585
R1062 B.n464 B.n463 585
R1063 B.n462 B.n38 585
R1064 B.n461 B.n460 585
R1065 B.n459 B.n39 585
R1066 B.n458 B.n457 585
R1067 B.n456 B.n40 585
R1068 B.n455 B.n454 585
R1069 B.n452 B.n41 585
R1070 B.n451 B.n450 585
R1071 B.n449 B.n44 585
R1072 B.n448 B.n447 585
R1073 B.n446 B.n45 585
R1074 B.n445 B.n444 585
R1075 B.n443 B.n46 585
R1076 B.n442 B.n441 585
R1077 B.n440 B.n47 585
R1078 B.n439 B.n438 585
R1079 B.n437 B.n48 585
R1080 B.n436 B.n435 585
R1081 B.n434 B.n49 585
R1082 B.n433 B.n432 585
R1083 B.n431 B.n50 585
R1084 B.n430 B.n429 585
R1085 B.n428 B.n51 585
R1086 B.n427 B.n426 585
R1087 B.n425 B.n52 585
R1088 B.n424 B.n423 585
R1089 B.n422 B.n53 585
R1090 B.n421 B.n420 585
R1091 B.n419 B.n54 585
R1092 B.n418 B.n417 585
R1093 B.n416 B.n55 585
R1094 B.n415 B.n414 585
R1095 B.n413 B.n56 585
R1096 B.n412 B.n411 585
R1097 B.n410 B.n57 585
R1098 B.n409 B.n408 585
R1099 B.n407 B.n58 585
R1100 B.n406 B.n405 585
R1101 B.n404 B.n59 585
R1102 B.n403 B.n402 585
R1103 B.n401 B.n60 585
R1104 B.n400 B.n399 585
R1105 B.n398 B.n61 585
R1106 B.n397 B.n396 585
R1107 B.n395 B.n62 585
R1108 B.n394 B.n393 585
R1109 B.n392 B.n63 585
R1110 B.n391 B.n390 585
R1111 B.n389 B.n64 585
R1112 B.n388 B.n387 585
R1113 B.n386 B.n65 585
R1114 B.n385 B.n384 585
R1115 B.n538 B.n537 585
R1116 B.n539 B.n10 585
R1117 B.n541 B.n540 585
R1118 B.n542 B.n9 585
R1119 B.n544 B.n543 585
R1120 B.n545 B.n8 585
R1121 B.n547 B.n546 585
R1122 B.n548 B.n7 585
R1123 B.n550 B.n549 585
R1124 B.n551 B.n6 585
R1125 B.n553 B.n552 585
R1126 B.n554 B.n5 585
R1127 B.n556 B.n555 585
R1128 B.n557 B.n4 585
R1129 B.n559 B.n558 585
R1130 B.n560 B.n3 585
R1131 B.n562 B.n561 585
R1132 B.n563 B.n0 585
R1133 B.n2 B.n1 585
R1134 B.n149 B.n148 585
R1135 B.n151 B.n150 585
R1136 B.n152 B.n147 585
R1137 B.n154 B.n153 585
R1138 B.n155 B.n146 585
R1139 B.n157 B.n156 585
R1140 B.n158 B.n145 585
R1141 B.n160 B.n159 585
R1142 B.n161 B.n144 585
R1143 B.n163 B.n162 585
R1144 B.n164 B.n143 585
R1145 B.n166 B.n165 585
R1146 B.n167 B.n142 585
R1147 B.n169 B.n168 585
R1148 B.n170 B.n141 585
R1149 B.n172 B.n171 585
R1150 B.n173 B.n140 585
R1151 B.n174 B.n173 487.695
R1152 B.n328 B.n85 487.695
R1153 B.n384 B.n383 487.695
R1154 B.n538 B.n11 487.695
R1155 B.n108 B.t4 434.351
R1156 B.n42 B.t2 434.351
R1157 B.n116 B.t10 434.351
R1158 B.n34 B.t8 434.351
R1159 B.n116 B.t9 428.803
R1160 B.n108 B.t3 428.803
R1161 B.n42 B.t0 428.803
R1162 B.n34 B.t6 428.803
R1163 B.n109 B.t5 400.024
R1164 B.n43 B.t1 400.024
R1165 B.n117 B.t11 400.024
R1166 B.n35 B.t7 400.024
R1167 B.n565 B.n564 256.663
R1168 B.n564 B.n563 235.042
R1169 B.n564 B.n2 235.042
R1170 B.n174 B.n139 163.367
R1171 B.n178 B.n139 163.367
R1172 B.n179 B.n178 163.367
R1173 B.n180 B.n179 163.367
R1174 B.n180 B.n137 163.367
R1175 B.n184 B.n137 163.367
R1176 B.n185 B.n184 163.367
R1177 B.n186 B.n185 163.367
R1178 B.n186 B.n135 163.367
R1179 B.n190 B.n135 163.367
R1180 B.n191 B.n190 163.367
R1181 B.n192 B.n191 163.367
R1182 B.n192 B.n133 163.367
R1183 B.n196 B.n133 163.367
R1184 B.n197 B.n196 163.367
R1185 B.n198 B.n197 163.367
R1186 B.n198 B.n131 163.367
R1187 B.n202 B.n131 163.367
R1188 B.n203 B.n202 163.367
R1189 B.n204 B.n203 163.367
R1190 B.n204 B.n129 163.367
R1191 B.n208 B.n129 163.367
R1192 B.n209 B.n208 163.367
R1193 B.n210 B.n209 163.367
R1194 B.n210 B.n127 163.367
R1195 B.n214 B.n127 163.367
R1196 B.n215 B.n214 163.367
R1197 B.n216 B.n215 163.367
R1198 B.n216 B.n125 163.367
R1199 B.n220 B.n125 163.367
R1200 B.n221 B.n220 163.367
R1201 B.n222 B.n221 163.367
R1202 B.n222 B.n123 163.367
R1203 B.n226 B.n123 163.367
R1204 B.n227 B.n226 163.367
R1205 B.n228 B.n227 163.367
R1206 B.n228 B.n121 163.367
R1207 B.n232 B.n121 163.367
R1208 B.n233 B.n232 163.367
R1209 B.n234 B.n233 163.367
R1210 B.n234 B.n119 163.367
R1211 B.n238 B.n119 163.367
R1212 B.n239 B.n238 163.367
R1213 B.n240 B.n239 163.367
R1214 B.n240 B.n115 163.367
R1215 B.n245 B.n115 163.367
R1216 B.n246 B.n245 163.367
R1217 B.n247 B.n246 163.367
R1218 B.n247 B.n113 163.367
R1219 B.n251 B.n113 163.367
R1220 B.n252 B.n251 163.367
R1221 B.n253 B.n252 163.367
R1222 B.n253 B.n111 163.367
R1223 B.n257 B.n111 163.367
R1224 B.n258 B.n257 163.367
R1225 B.n258 B.n107 163.367
R1226 B.n262 B.n107 163.367
R1227 B.n263 B.n262 163.367
R1228 B.n264 B.n263 163.367
R1229 B.n264 B.n105 163.367
R1230 B.n268 B.n105 163.367
R1231 B.n269 B.n268 163.367
R1232 B.n270 B.n269 163.367
R1233 B.n270 B.n103 163.367
R1234 B.n274 B.n103 163.367
R1235 B.n275 B.n274 163.367
R1236 B.n276 B.n275 163.367
R1237 B.n276 B.n101 163.367
R1238 B.n280 B.n101 163.367
R1239 B.n281 B.n280 163.367
R1240 B.n282 B.n281 163.367
R1241 B.n282 B.n99 163.367
R1242 B.n286 B.n99 163.367
R1243 B.n287 B.n286 163.367
R1244 B.n288 B.n287 163.367
R1245 B.n288 B.n97 163.367
R1246 B.n292 B.n97 163.367
R1247 B.n293 B.n292 163.367
R1248 B.n294 B.n293 163.367
R1249 B.n294 B.n95 163.367
R1250 B.n298 B.n95 163.367
R1251 B.n299 B.n298 163.367
R1252 B.n300 B.n299 163.367
R1253 B.n300 B.n93 163.367
R1254 B.n304 B.n93 163.367
R1255 B.n305 B.n304 163.367
R1256 B.n306 B.n305 163.367
R1257 B.n306 B.n91 163.367
R1258 B.n310 B.n91 163.367
R1259 B.n311 B.n310 163.367
R1260 B.n312 B.n311 163.367
R1261 B.n312 B.n89 163.367
R1262 B.n316 B.n89 163.367
R1263 B.n317 B.n316 163.367
R1264 B.n318 B.n317 163.367
R1265 B.n318 B.n87 163.367
R1266 B.n322 B.n87 163.367
R1267 B.n323 B.n322 163.367
R1268 B.n324 B.n323 163.367
R1269 B.n324 B.n85 163.367
R1270 B.n383 B.n382 163.367
R1271 B.n382 B.n67 163.367
R1272 B.n378 B.n67 163.367
R1273 B.n378 B.n377 163.367
R1274 B.n377 B.n376 163.367
R1275 B.n376 B.n69 163.367
R1276 B.n372 B.n69 163.367
R1277 B.n372 B.n371 163.367
R1278 B.n371 B.n370 163.367
R1279 B.n370 B.n71 163.367
R1280 B.n366 B.n71 163.367
R1281 B.n366 B.n365 163.367
R1282 B.n365 B.n364 163.367
R1283 B.n364 B.n73 163.367
R1284 B.n360 B.n73 163.367
R1285 B.n360 B.n359 163.367
R1286 B.n359 B.n358 163.367
R1287 B.n358 B.n75 163.367
R1288 B.n354 B.n75 163.367
R1289 B.n354 B.n353 163.367
R1290 B.n353 B.n352 163.367
R1291 B.n352 B.n77 163.367
R1292 B.n348 B.n77 163.367
R1293 B.n348 B.n347 163.367
R1294 B.n347 B.n346 163.367
R1295 B.n346 B.n79 163.367
R1296 B.n342 B.n79 163.367
R1297 B.n342 B.n341 163.367
R1298 B.n341 B.n340 163.367
R1299 B.n340 B.n81 163.367
R1300 B.n336 B.n81 163.367
R1301 B.n336 B.n335 163.367
R1302 B.n335 B.n334 163.367
R1303 B.n334 B.n83 163.367
R1304 B.n330 B.n83 163.367
R1305 B.n330 B.n329 163.367
R1306 B.n329 B.n328 163.367
R1307 B.n534 B.n11 163.367
R1308 B.n534 B.n533 163.367
R1309 B.n533 B.n532 163.367
R1310 B.n532 B.n13 163.367
R1311 B.n528 B.n13 163.367
R1312 B.n528 B.n527 163.367
R1313 B.n527 B.n526 163.367
R1314 B.n526 B.n15 163.367
R1315 B.n522 B.n15 163.367
R1316 B.n522 B.n521 163.367
R1317 B.n521 B.n520 163.367
R1318 B.n520 B.n17 163.367
R1319 B.n516 B.n17 163.367
R1320 B.n516 B.n515 163.367
R1321 B.n515 B.n514 163.367
R1322 B.n514 B.n19 163.367
R1323 B.n510 B.n19 163.367
R1324 B.n510 B.n509 163.367
R1325 B.n509 B.n508 163.367
R1326 B.n508 B.n21 163.367
R1327 B.n504 B.n21 163.367
R1328 B.n504 B.n503 163.367
R1329 B.n503 B.n502 163.367
R1330 B.n502 B.n23 163.367
R1331 B.n498 B.n23 163.367
R1332 B.n498 B.n497 163.367
R1333 B.n497 B.n496 163.367
R1334 B.n496 B.n25 163.367
R1335 B.n492 B.n25 163.367
R1336 B.n492 B.n491 163.367
R1337 B.n491 B.n490 163.367
R1338 B.n490 B.n27 163.367
R1339 B.n486 B.n27 163.367
R1340 B.n486 B.n485 163.367
R1341 B.n485 B.n484 163.367
R1342 B.n484 B.n29 163.367
R1343 B.n480 B.n29 163.367
R1344 B.n480 B.n479 163.367
R1345 B.n479 B.n478 163.367
R1346 B.n478 B.n31 163.367
R1347 B.n474 B.n31 163.367
R1348 B.n474 B.n473 163.367
R1349 B.n473 B.n472 163.367
R1350 B.n472 B.n33 163.367
R1351 B.n468 B.n33 163.367
R1352 B.n468 B.n467 163.367
R1353 B.n467 B.n37 163.367
R1354 B.n463 B.n37 163.367
R1355 B.n463 B.n462 163.367
R1356 B.n462 B.n461 163.367
R1357 B.n461 B.n39 163.367
R1358 B.n457 B.n39 163.367
R1359 B.n457 B.n456 163.367
R1360 B.n456 B.n455 163.367
R1361 B.n455 B.n41 163.367
R1362 B.n450 B.n41 163.367
R1363 B.n450 B.n449 163.367
R1364 B.n449 B.n448 163.367
R1365 B.n448 B.n45 163.367
R1366 B.n444 B.n45 163.367
R1367 B.n444 B.n443 163.367
R1368 B.n443 B.n442 163.367
R1369 B.n442 B.n47 163.367
R1370 B.n438 B.n47 163.367
R1371 B.n438 B.n437 163.367
R1372 B.n437 B.n436 163.367
R1373 B.n436 B.n49 163.367
R1374 B.n432 B.n49 163.367
R1375 B.n432 B.n431 163.367
R1376 B.n431 B.n430 163.367
R1377 B.n430 B.n51 163.367
R1378 B.n426 B.n51 163.367
R1379 B.n426 B.n425 163.367
R1380 B.n425 B.n424 163.367
R1381 B.n424 B.n53 163.367
R1382 B.n420 B.n53 163.367
R1383 B.n420 B.n419 163.367
R1384 B.n419 B.n418 163.367
R1385 B.n418 B.n55 163.367
R1386 B.n414 B.n55 163.367
R1387 B.n414 B.n413 163.367
R1388 B.n413 B.n412 163.367
R1389 B.n412 B.n57 163.367
R1390 B.n408 B.n57 163.367
R1391 B.n408 B.n407 163.367
R1392 B.n407 B.n406 163.367
R1393 B.n406 B.n59 163.367
R1394 B.n402 B.n59 163.367
R1395 B.n402 B.n401 163.367
R1396 B.n401 B.n400 163.367
R1397 B.n400 B.n61 163.367
R1398 B.n396 B.n61 163.367
R1399 B.n396 B.n395 163.367
R1400 B.n395 B.n394 163.367
R1401 B.n394 B.n63 163.367
R1402 B.n390 B.n63 163.367
R1403 B.n390 B.n389 163.367
R1404 B.n389 B.n388 163.367
R1405 B.n388 B.n65 163.367
R1406 B.n384 B.n65 163.367
R1407 B.n539 B.n538 163.367
R1408 B.n540 B.n539 163.367
R1409 B.n540 B.n9 163.367
R1410 B.n544 B.n9 163.367
R1411 B.n545 B.n544 163.367
R1412 B.n546 B.n545 163.367
R1413 B.n546 B.n7 163.367
R1414 B.n550 B.n7 163.367
R1415 B.n551 B.n550 163.367
R1416 B.n552 B.n551 163.367
R1417 B.n552 B.n5 163.367
R1418 B.n556 B.n5 163.367
R1419 B.n557 B.n556 163.367
R1420 B.n558 B.n557 163.367
R1421 B.n558 B.n3 163.367
R1422 B.n562 B.n3 163.367
R1423 B.n563 B.n562 163.367
R1424 B.n149 B.n2 163.367
R1425 B.n150 B.n149 163.367
R1426 B.n150 B.n147 163.367
R1427 B.n154 B.n147 163.367
R1428 B.n155 B.n154 163.367
R1429 B.n156 B.n155 163.367
R1430 B.n156 B.n145 163.367
R1431 B.n160 B.n145 163.367
R1432 B.n161 B.n160 163.367
R1433 B.n162 B.n161 163.367
R1434 B.n162 B.n143 163.367
R1435 B.n166 B.n143 163.367
R1436 B.n167 B.n166 163.367
R1437 B.n168 B.n167 163.367
R1438 B.n168 B.n141 163.367
R1439 B.n172 B.n141 163.367
R1440 B.n173 B.n172 163.367
R1441 B.n243 B.n117 59.5399
R1442 B.n110 B.n109 59.5399
R1443 B.n453 B.n43 59.5399
R1444 B.n36 B.n35 59.5399
R1445 B.n117 B.n116 34.3278
R1446 B.n109 B.n108 34.3278
R1447 B.n43 B.n42 34.3278
R1448 B.n35 B.n34 34.3278
R1449 B.n537 B.n536 31.6883
R1450 B.n385 B.n66 31.6883
R1451 B.n327 B.n326 31.6883
R1452 B.n175 B.n140 31.6883
R1453 B B.n565 18.0485
R1454 B.n537 B.n10 10.6151
R1455 B.n541 B.n10 10.6151
R1456 B.n542 B.n541 10.6151
R1457 B.n543 B.n542 10.6151
R1458 B.n543 B.n8 10.6151
R1459 B.n547 B.n8 10.6151
R1460 B.n548 B.n547 10.6151
R1461 B.n549 B.n548 10.6151
R1462 B.n549 B.n6 10.6151
R1463 B.n553 B.n6 10.6151
R1464 B.n554 B.n553 10.6151
R1465 B.n555 B.n554 10.6151
R1466 B.n555 B.n4 10.6151
R1467 B.n559 B.n4 10.6151
R1468 B.n560 B.n559 10.6151
R1469 B.n561 B.n560 10.6151
R1470 B.n561 B.n0 10.6151
R1471 B.n536 B.n535 10.6151
R1472 B.n535 B.n12 10.6151
R1473 B.n531 B.n12 10.6151
R1474 B.n531 B.n530 10.6151
R1475 B.n530 B.n529 10.6151
R1476 B.n529 B.n14 10.6151
R1477 B.n525 B.n14 10.6151
R1478 B.n525 B.n524 10.6151
R1479 B.n524 B.n523 10.6151
R1480 B.n523 B.n16 10.6151
R1481 B.n519 B.n16 10.6151
R1482 B.n519 B.n518 10.6151
R1483 B.n518 B.n517 10.6151
R1484 B.n517 B.n18 10.6151
R1485 B.n513 B.n18 10.6151
R1486 B.n513 B.n512 10.6151
R1487 B.n512 B.n511 10.6151
R1488 B.n511 B.n20 10.6151
R1489 B.n507 B.n20 10.6151
R1490 B.n507 B.n506 10.6151
R1491 B.n506 B.n505 10.6151
R1492 B.n505 B.n22 10.6151
R1493 B.n501 B.n22 10.6151
R1494 B.n501 B.n500 10.6151
R1495 B.n500 B.n499 10.6151
R1496 B.n499 B.n24 10.6151
R1497 B.n495 B.n24 10.6151
R1498 B.n495 B.n494 10.6151
R1499 B.n494 B.n493 10.6151
R1500 B.n493 B.n26 10.6151
R1501 B.n489 B.n26 10.6151
R1502 B.n489 B.n488 10.6151
R1503 B.n488 B.n487 10.6151
R1504 B.n487 B.n28 10.6151
R1505 B.n483 B.n28 10.6151
R1506 B.n483 B.n482 10.6151
R1507 B.n482 B.n481 10.6151
R1508 B.n481 B.n30 10.6151
R1509 B.n477 B.n30 10.6151
R1510 B.n477 B.n476 10.6151
R1511 B.n476 B.n475 10.6151
R1512 B.n475 B.n32 10.6151
R1513 B.n471 B.n32 10.6151
R1514 B.n471 B.n470 10.6151
R1515 B.n470 B.n469 10.6151
R1516 B.n466 B.n465 10.6151
R1517 B.n465 B.n464 10.6151
R1518 B.n464 B.n38 10.6151
R1519 B.n460 B.n38 10.6151
R1520 B.n460 B.n459 10.6151
R1521 B.n459 B.n458 10.6151
R1522 B.n458 B.n40 10.6151
R1523 B.n454 B.n40 10.6151
R1524 B.n452 B.n451 10.6151
R1525 B.n451 B.n44 10.6151
R1526 B.n447 B.n44 10.6151
R1527 B.n447 B.n446 10.6151
R1528 B.n446 B.n445 10.6151
R1529 B.n445 B.n46 10.6151
R1530 B.n441 B.n46 10.6151
R1531 B.n441 B.n440 10.6151
R1532 B.n440 B.n439 10.6151
R1533 B.n439 B.n48 10.6151
R1534 B.n435 B.n48 10.6151
R1535 B.n435 B.n434 10.6151
R1536 B.n434 B.n433 10.6151
R1537 B.n433 B.n50 10.6151
R1538 B.n429 B.n50 10.6151
R1539 B.n429 B.n428 10.6151
R1540 B.n428 B.n427 10.6151
R1541 B.n427 B.n52 10.6151
R1542 B.n423 B.n52 10.6151
R1543 B.n423 B.n422 10.6151
R1544 B.n422 B.n421 10.6151
R1545 B.n421 B.n54 10.6151
R1546 B.n417 B.n54 10.6151
R1547 B.n417 B.n416 10.6151
R1548 B.n416 B.n415 10.6151
R1549 B.n415 B.n56 10.6151
R1550 B.n411 B.n56 10.6151
R1551 B.n411 B.n410 10.6151
R1552 B.n410 B.n409 10.6151
R1553 B.n409 B.n58 10.6151
R1554 B.n405 B.n58 10.6151
R1555 B.n405 B.n404 10.6151
R1556 B.n404 B.n403 10.6151
R1557 B.n403 B.n60 10.6151
R1558 B.n399 B.n60 10.6151
R1559 B.n399 B.n398 10.6151
R1560 B.n398 B.n397 10.6151
R1561 B.n397 B.n62 10.6151
R1562 B.n393 B.n62 10.6151
R1563 B.n393 B.n392 10.6151
R1564 B.n392 B.n391 10.6151
R1565 B.n391 B.n64 10.6151
R1566 B.n387 B.n64 10.6151
R1567 B.n387 B.n386 10.6151
R1568 B.n386 B.n385 10.6151
R1569 B.n381 B.n66 10.6151
R1570 B.n381 B.n380 10.6151
R1571 B.n380 B.n379 10.6151
R1572 B.n379 B.n68 10.6151
R1573 B.n375 B.n68 10.6151
R1574 B.n375 B.n374 10.6151
R1575 B.n374 B.n373 10.6151
R1576 B.n373 B.n70 10.6151
R1577 B.n369 B.n70 10.6151
R1578 B.n369 B.n368 10.6151
R1579 B.n368 B.n367 10.6151
R1580 B.n367 B.n72 10.6151
R1581 B.n363 B.n72 10.6151
R1582 B.n363 B.n362 10.6151
R1583 B.n362 B.n361 10.6151
R1584 B.n361 B.n74 10.6151
R1585 B.n357 B.n74 10.6151
R1586 B.n357 B.n356 10.6151
R1587 B.n356 B.n355 10.6151
R1588 B.n355 B.n76 10.6151
R1589 B.n351 B.n76 10.6151
R1590 B.n351 B.n350 10.6151
R1591 B.n350 B.n349 10.6151
R1592 B.n349 B.n78 10.6151
R1593 B.n345 B.n78 10.6151
R1594 B.n345 B.n344 10.6151
R1595 B.n344 B.n343 10.6151
R1596 B.n343 B.n80 10.6151
R1597 B.n339 B.n80 10.6151
R1598 B.n339 B.n338 10.6151
R1599 B.n338 B.n337 10.6151
R1600 B.n337 B.n82 10.6151
R1601 B.n333 B.n82 10.6151
R1602 B.n333 B.n332 10.6151
R1603 B.n332 B.n331 10.6151
R1604 B.n331 B.n84 10.6151
R1605 B.n327 B.n84 10.6151
R1606 B.n148 B.n1 10.6151
R1607 B.n151 B.n148 10.6151
R1608 B.n152 B.n151 10.6151
R1609 B.n153 B.n152 10.6151
R1610 B.n153 B.n146 10.6151
R1611 B.n157 B.n146 10.6151
R1612 B.n158 B.n157 10.6151
R1613 B.n159 B.n158 10.6151
R1614 B.n159 B.n144 10.6151
R1615 B.n163 B.n144 10.6151
R1616 B.n164 B.n163 10.6151
R1617 B.n165 B.n164 10.6151
R1618 B.n165 B.n142 10.6151
R1619 B.n169 B.n142 10.6151
R1620 B.n170 B.n169 10.6151
R1621 B.n171 B.n170 10.6151
R1622 B.n171 B.n140 10.6151
R1623 B.n176 B.n175 10.6151
R1624 B.n177 B.n176 10.6151
R1625 B.n177 B.n138 10.6151
R1626 B.n181 B.n138 10.6151
R1627 B.n182 B.n181 10.6151
R1628 B.n183 B.n182 10.6151
R1629 B.n183 B.n136 10.6151
R1630 B.n187 B.n136 10.6151
R1631 B.n188 B.n187 10.6151
R1632 B.n189 B.n188 10.6151
R1633 B.n189 B.n134 10.6151
R1634 B.n193 B.n134 10.6151
R1635 B.n194 B.n193 10.6151
R1636 B.n195 B.n194 10.6151
R1637 B.n195 B.n132 10.6151
R1638 B.n199 B.n132 10.6151
R1639 B.n200 B.n199 10.6151
R1640 B.n201 B.n200 10.6151
R1641 B.n201 B.n130 10.6151
R1642 B.n205 B.n130 10.6151
R1643 B.n206 B.n205 10.6151
R1644 B.n207 B.n206 10.6151
R1645 B.n207 B.n128 10.6151
R1646 B.n211 B.n128 10.6151
R1647 B.n212 B.n211 10.6151
R1648 B.n213 B.n212 10.6151
R1649 B.n213 B.n126 10.6151
R1650 B.n217 B.n126 10.6151
R1651 B.n218 B.n217 10.6151
R1652 B.n219 B.n218 10.6151
R1653 B.n219 B.n124 10.6151
R1654 B.n223 B.n124 10.6151
R1655 B.n224 B.n223 10.6151
R1656 B.n225 B.n224 10.6151
R1657 B.n225 B.n122 10.6151
R1658 B.n229 B.n122 10.6151
R1659 B.n230 B.n229 10.6151
R1660 B.n231 B.n230 10.6151
R1661 B.n231 B.n120 10.6151
R1662 B.n235 B.n120 10.6151
R1663 B.n236 B.n235 10.6151
R1664 B.n237 B.n236 10.6151
R1665 B.n237 B.n118 10.6151
R1666 B.n241 B.n118 10.6151
R1667 B.n242 B.n241 10.6151
R1668 B.n244 B.n114 10.6151
R1669 B.n248 B.n114 10.6151
R1670 B.n249 B.n248 10.6151
R1671 B.n250 B.n249 10.6151
R1672 B.n250 B.n112 10.6151
R1673 B.n254 B.n112 10.6151
R1674 B.n255 B.n254 10.6151
R1675 B.n256 B.n255 10.6151
R1676 B.n260 B.n259 10.6151
R1677 B.n261 B.n260 10.6151
R1678 B.n261 B.n106 10.6151
R1679 B.n265 B.n106 10.6151
R1680 B.n266 B.n265 10.6151
R1681 B.n267 B.n266 10.6151
R1682 B.n267 B.n104 10.6151
R1683 B.n271 B.n104 10.6151
R1684 B.n272 B.n271 10.6151
R1685 B.n273 B.n272 10.6151
R1686 B.n273 B.n102 10.6151
R1687 B.n277 B.n102 10.6151
R1688 B.n278 B.n277 10.6151
R1689 B.n279 B.n278 10.6151
R1690 B.n279 B.n100 10.6151
R1691 B.n283 B.n100 10.6151
R1692 B.n284 B.n283 10.6151
R1693 B.n285 B.n284 10.6151
R1694 B.n285 B.n98 10.6151
R1695 B.n289 B.n98 10.6151
R1696 B.n290 B.n289 10.6151
R1697 B.n291 B.n290 10.6151
R1698 B.n291 B.n96 10.6151
R1699 B.n295 B.n96 10.6151
R1700 B.n296 B.n295 10.6151
R1701 B.n297 B.n296 10.6151
R1702 B.n297 B.n94 10.6151
R1703 B.n301 B.n94 10.6151
R1704 B.n302 B.n301 10.6151
R1705 B.n303 B.n302 10.6151
R1706 B.n303 B.n92 10.6151
R1707 B.n307 B.n92 10.6151
R1708 B.n308 B.n307 10.6151
R1709 B.n309 B.n308 10.6151
R1710 B.n309 B.n90 10.6151
R1711 B.n313 B.n90 10.6151
R1712 B.n314 B.n313 10.6151
R1713 B.n315 B.n314 10.6151
R1714 B.n315 B.n88 10.6151
R1715 B.n319 B.n88 10.6151
R1716 B.n320 B.n319 10.6151
R1717 B.n321 B.n320 10.6151
R1718 B.n321 B.n86 10.6151
R1719 B.n325 B.n86 10.6151
R1720 B.n326 B.n325 10.6151
R1721 B.n565 B.n0 8.11757
R1722 B.n565 B.n1 8.11757
R1723 B.n466 B.n36 6.5566
R1724 B.n454 B.n453 6.5566
R1725 B.n244 B.n243 6.5566
R1726 B.n256 B.n110 6.5566
R1727 B.n469 B.n36 4.05904
R1728 B.n453 B.n452 4.05904
R1729 B.n243 B.n242 4.05904
R1730 B.n259 B.n110 4.05904
C0 VN w_n1678_n3640# 2.23544f
C1 B VDD2 1.66245f
C2 B VP 1.21516f
C3 VDD2 VP 0.284975f
C4 VTAIL B 3.3972f
C5 VTAIL VDD2 5.52858f
C6 VTAIL VP 2.27381f
C7 VDD1 B 1.6425f
C8 VDD1 VDD2 0.539758f
C9 VDD1 VP 2.85988f
C10 VDD1 VTAIL 5.48807f
C11 B w_n1678_n3640# 7.93605f
C12 VDD2 w_n1678_n3640# 1.76129f
C13 VP w_n1678_n3640# 2.44668f
C14 B VN 0.87252f
C15 VTAIL w_n1678_n3640# 3.00153f
C16 VN VDD2 2.72656f
C17 VN VP 5.15913f
C18 VDD1 w_n1678_n3640# 1.74911f
C19 VTAIL VN 2.25934f
C20 VDD1 VN 0.147924f
C21 VDD2 VSUBS 0.842528f
C22 VDD1 VSUBS 3.51002f
C23 VTAIL VSUBS 0.923901f
C24 VN VSUBS 7.86341f
C25 VP VSUBS 1.387786f
C26 B VSUBS 3.151361f
C27 w_n1678_n3640# VSUBS 75.0469f
C28 B.n0 VSUBS 0.005786f
C29 B.n1 VSUBS 0.005786f
C30 B.n2 VSUBS 0.008557f
C31 B.n3 VSUBS 0.006557f
C32 B.n4 VSUBS 0.006557f
C33 B.n5 VSUBS 0.006557f
C34 B.n6 VSUBS 0.006557f
C35 B.n7 VSUBS 0.006557f
C36 B.n8 VSUBS 0.006557f
C37 B.n9 VSUBS 0.006557f
C38 B.n10 VSUBS 0.006557f
C39 B.n11 VSUBS 0.015501f
C40 B.n12 VSUBS 0.006557f
C41 B.n13 VSUBS 0.006557f
C42 B.n14 VSUBS 0.006557f
C43 B.n15 VSUBS 0.006557f
C44 B.n16 VSUBS 0.006557f
C45 B.n17 VSUBS 0.006557f
C46 B.n18 VSUBS 0.006557f
C47 B.n19 VSUBS 0.006557f
C48 B.n20 VSUBS 0.006557f
C49 B.n21 VSUBS 0.006557f
C50 B.n22 VSUBS 0.006557f
C51 B.n23 VSUBS 0.006557f
C52 B.n24 VSUBS 0.006557f
C53 B.n25 VSUBS 0.006557f
C54 B.n26 VSUBS 0.006557f
C55 B.n27 VSUBS 0.006557f
C56 B.n28 VSUBS 0.006557f
C57 B.n29 VSUBS 0.006557f
C58 B.n30 VSUBS 0.006557f
C59 B.n31 VSUBS 0.006557f
C60 B.n32 VSUBS 0.006557f
C61 B.n33 VSUBS 0.006557f
C62 B.t7 VSUBS 0.2263f
C63 B.t8 VSUBS 0.245227f
C64 B.t6 VSUBS 0.779846f
C65 B.n34 VSUBS 0.364531f
C66 B.n35 VSUBS 0.248841f
C67 B.n36 VSUBS 0.015192f
C68 B.n37 VSUBS 0.006557f
C69 B.n38 VSUBS 0.006557f
C70 B.n39 VSUBS 0.006557f
C71 B.n40 VSUBS 0.006557f
C72 B.n41 VSUBS 0.006557f
C73 B.t1 VSUBS 0.226303f
C74 B.t2 VSUBS 0.24523f
C75 B.t0 VSUBS 0.779846f
C76 B.n42 VSUBS 0.364529f
C77 B.n43 VSUBS 0.248838f
C78 B.n44 VSUBS 0.006557f
C79 B.n45 VSUBS 0.006557f
C80 B.n46 VSUBS 0.006557f
C81 B.n47 VSUBS 0.006557f
C82 B.n48 VSUBS 0.006557f
C83 B.n49 VSUBS 0.006557f
C84 B.n50 VSUBS 0.006557f
C85 B.n51 VSUBS 0.006557f
C86 B.n52 VSUBS 0.006557f
C87 B.n53 VSUBS 0.006557f
C88 B.n54 VSUBS 0.006557f
C89 B.n55 VSUBS 0.006557f
C90 B.n56 VSUBS 0.006557f
C91 B.n57 VSUBS 0.006557f
C92 B.n58 VSUBS 0.006557f
C93 B.n59 VSUBS 0.006557f
C94 B.n60 VSUBS 0.006557f
C95 B.n61 VSUBS 0.006557f
C96 B.n62 VSUBS 0.006557f
C97 B.n63 VSUBS 0.006557f
C98 B.n64 VSUBS 0.006557f
C99 B.n65 VSUBS 0.006557f
C100 B.n66 VSUBS 0.014585f
C101 B.n67 VSUBS 0.006557f
C102 B.n68 VSUBS 0.006557f
C103 B.n69 VSUBS 0.006557f
C104 B.n70 VSUBS 0.006557f
C105 B.n71 VSUBS 0.006557f
C106 B.n72 VSUBS 0.006557f
C107 B.n73 VSUBS 0.006557f
C108 B.n74 VSUBS 0.006557f
C109 B.n75 VSUBS 0.006557f
C110 B.n76 VSUBS 0.006557f
C111 B.n77 VSUBS 0.006557f
C112 B.n78 VSUBS 0.006557f
C113 B.n79 VSUBS 0.006557f
C114 B.n80 VSUBS 0.006557f
C115 B.n81 VSUBS 0.006557f
C116 B.n82 VSUBS 0.006557f
C117 B.n83 VSUBS 0.006557f
C118 B.n84 VSUBS 0.006557f
C119 B.n85 VSUBS 0.015501f
C120 B.n86 VSUBS 0.006557f
C121 B.n87 VSUBS 0.006557f
C122 B.n88 VSUBS 0.006557f
C123 B.n89 VSUBS 0.006557f
C124 B.n90 VSUBS 0.006557f
C125 B.n91 VSUBS 0.006557f
C126 B.n92 VSUBS 0.006557f
C127 B.n93 VSUBS 0.006557f
C128 B.n94 VSUBS 0.006557f
C129 B.n95 VSUBS 0.006557f
C130 B.n96 VSUBS 0.006557f
C131 B.n97 VSUBS 0.006557f
C132 B.n98 VSUBS 0.006557f
C133 B.n99 VSUBS 0.006557f
C134 B.n100 VSUBS 0.006557f
C135 B.n101 VSUBS 0.006557f
C136 B.n102 VSUBS 0.006557f
C137 B.n103 VSUBS 0.006557f
C138 B.n104 VSUBS 0.006557f
C139 B.n105 VSUBS 0.006557f
C140 B.n106 VSUBS 0.006557f
C141 B.n107 VSUBS 0.006557f
C142 B.t5 VSUBS 0.226303f
C143 B.t4 VSUBS 0.24523f
C144 B.t3 VSUBS 0.779846f
C145 B.n108 VSUBS 0.364529f
C146 B.n109 VSUBS 0.248838f
C147 B.n110 VSUBS 0.015192f
C148 B.n111 VSUBS 0.006557f
C149 B.n112 VSUBS 0.006557f
C150 B.n113 VSUBS 0.006557f
C151 B.n114 VSUBS 0.006557f
C152 B.n115 VSUBS 0.006557f
C153 B.t11 VSUBS 0.2263f
C154 B.t10 VSUBS 0.245227f
C155 B.t9 VSUBS 0.779846f
C156 B.n116 VSUBS 0.364531f
C157 B.n117 VSUBS 0.248841f
C158 B.n118 VSUBS 0.006557f
C159 B.n119 VSUBS 0.006557f
C160 B.n120 VSUBS 0.006557f
C161 B.n121 VSUBS 0.006557f
C162 B.n122 VSUBS 0.006557f
C163 B.n123 VSUBS 0.006557f
C164 B.n124 VSUBS 0.006557f
C165 B.n125 VSUBS 0.006557f
C166 B.n126 VSUBS 0.006557f
C167 B.n127 VSUBS 0.006557f
C168 B.n128 VSUBS 0.006557f
C169 B.n129 VSUBS 0.006557f
C170 B.n130 VSUBS 0.006557f
C171 B.n131 VSUBS 0.006557f
C172 B.n132 VSUBS 0.006557f
C173 B.n133 VSUBS 0.006557f
C174 B.n134 VSUBS 0.006557f
C175 B.n135 VSUBS 0.006557f
C176 B.n136 VSUBS 0.006557f
C177 B.n137 VSUBS 0.006557f
C178 B.n138 VSUBS 0.006557f
C179 B.n139 VSUBS 0.006557f
C180 B.n140 VSUBS 0.014585f
C181 B.n141 VSUBS 0.006557f
C182 B.n142 VSUBS 0.006557f
C183 B.n143 VSUBS 0.006557f
C184 B.n144 VSUBS 0.006557f
C185 B.n145 VSUBS 0.006557f
C186 B.n146 VSUBS 0.006557f
C187 B.n147 VSUBS 0.006557f
C188 B.n148 VSUBS 0.006557f
C189 B.n149 VSUBS 0.006557f
C190 B.n150 VSUBS 0.006557f
C191 B.n151 VSUBS 0.006557f
C192 B.n152 VSUBS 0.006557f
C193 B.n153 VSUBS 0.006557f
C194 B.n154 VSUBS 0.006557f
C195 B.n155 VSUBS 0.006557f
C196 B.n156 VSUBS 0.006557f
C197 B.n157 VSUBS 0.006557f
C198 B.n158 VSUBS 0.006557f
C199 B.n159 VSUBS 0.006557f
C200 B.n160 VSUBS 0.006557f
C201 B.n161 VSUBS 0.006557f
C202 B.n162 VSUBS 0.006557f
C203 B.n163 VSUBS 0.006557f
C204 B.n164 VSUBS 0.006557f
C205 B.n165 VSUBS 0.006557f
C206 B.n166 VSUBS 0.006557f
C207 B.n167 VSUBS 0.006557f
C208 B.n168 VSUBS 0.006557f
C209 B.n169 VSUBS 0.006557f
C210 B.n170 VSUBS 0.006557f
C211 B.n171 VSUBS 0.006557f
C212 B.n172 VSUBS 0.006557f
C213 B.n173 VSUBS 0.014585f
C214 B.n174 VSUBS 0.015501f
C215 B.n175 VSUBS 0.015501f
C216 B.n176 VSUBS 0.006557f
C217 B.n177 VSUBS 0.006557f
C218 B.n178 VSUBS 0.006557f
C219 B.n179 VSUBS 0.006557f
C220 B.n180 VSUBS 0.006557f
C221 B.n181 VSUBS 0.006557f
C222 B.n182 VSUBS 0.006557f
C223 B.n183 VSUBS 0.006557f
C224 B.n184 VSUBS 0.006557f
C225 B.n185 VSUBS 0.006557f
C226 B.n186 VSUBS 0.006557f
C227 B.n187 VSUBS 0.006557f
C228 B.n188 VSUBS 0.006557f
C229 B.n189 VSUBS 0.006557f
C230 B.n190 VSUBS 0.006557f
C231 B.n191 VSUBS 0.006557f
C232 B.n192 VSUBS 0.006557f
C233 B.n193 VSUBS 0.006557f
C234 B.n194 VSUBS 0.006557f
C235 B.n195 VSUBS 0.006557f
C236 B.n196 VSUBS 0.006557f
C237 B.n197 VSUBS 0.006557f
C238 B.n198 VSUBS 0.006557f
C239 B.n199 VSUBS 0.006557f
C240 B.n200 VSUBS 0.006557f
C241 B.n201 VSUBS 0.006557f
C242 B.n202 VSUBS 0.006557f
C243 B.n203 VSUBS 0.006557f
C244 B.n204 VSUBS 0.006557f
C245 B.n205 VSUBS 0.006557f
C246 B.n206 VSUBS 0.006557f
C247 B.n207 VSUBS 0.006557f
C248 B.n208 VSUBS 0.006557f
C249 B.n209 VSUBS 0.006557f
C250 B.n210 VSUBS 0.006557f
C251 B.n211 VSUBS 0.006557f
C252 B.n212 VSUBS 0.006557f
C253 B.n213 VSUBS 0.006557f
C254 B.n214 VSUBS 0.006557f
C255 B.n215 VSUBS 0.006557f
C256 B.n216 VSUBS 0.006557f
C257 B.n217 VSUBS 0.006557f
C258 B.n218 VSUBS 0.006557f
C259 B.n219 VSUBS 0.006557f
C260 B.n220 VSUBS 0.006557f
C261 B.n221 VSUBS 0.006557f
C262 B.n222 VSUBS 0.006557f
C263 B.n223 VSUBS 0.006557f
C264 B.n224 VSUBS 0.006557f
C265 B.n225 VSUBS 0.006557f
C266 B.n226 VSUBS 0.006557f
C267 B.n227 VSUBS 0.006557f
C268 B.n228 VSUBS 0.006557f
C269 B.n229 VSUBS 0.006557f
C270 B.n230 VSUBS 0.006557f
C271 B.n231 VSUBS 0.006557f
C272 B.n232 VSUBS 0.006557f
C273 B.n233 VSUBS 0.006557f
C274 B.n234 VSUBS 0.006557f
C275 B.n235 VSUBS 0.006557f
C276 B.n236 VSUBS 0.006557f
C277 B.n237 VSUBS 0.006557f
C278 B.n238 VSUBS 0.006557f
C279 B.n239 VSUBS 0.006557f
C280 B.n240 VSUBS 0.006557f
C281 B.n241 VSUBS 0.006557f
C282 B.n242 VSUBS 0.004532f
C283 B.n243 VSUBS 0.015192f
C284 B.n244 VSUBS 0.005304f
C285 B.n245 VSUBS 0.006557f
C286 B.n246 VSUBS 0.006557f
C287 B.n247 VSUBS 0.006557f
C288 B.n248 VSUBS 0.006557f
C289 B.n249 VSUBS 0.006557f
C290 B.n250 VSUBS 0.006557f
C291 B.n251 VSUBS 0.006557f
C292 B.n252 VSUBS 0.006557f
C293 B.n253 VSUBS 0.006557f
C294 B.n254 VSUBS 0.006557f
C295 B.n255 VSUBS 0.006557f
C296 B.n256 VSUBS 0.005304f
C297 B.n257 VSUBS 0.006557f
C298 B.n258 VSUBS 0.006557f
C299 B.n259 VSUBS 0.004532f
C300 B.n260 VSUBS 0.006557f
C301 B.n261 VSUBS 0.006557f
C302 B.n262 VSUBS 0.006557f
C303 B.n263 VSUBS 0.006557f
C304 B.n264 VSUBS 0.006557f
C305 B.n265 VSUBS 0.006557f
C306 B.n266 VSUBS 0.006557f
C307 B.n267 VSUBS 0.006557f
C308 B.n268 VSUBS 0.006557f
C309 B.n269 VSUBS 0.006557f
C310 B.n270 VSUBS 0.006557f
C311 B.n271 VSUBS 0.006557f
C312 B.n272 VSUBS 0.006557f
C313 B.n273 VSUBS 0.006557f
C314 B.n274 VSUBS 0.006557f
C315 B.n275 VSUBS 0.006557f
C316 B.n276 VSUBS 0.006557f
C317 B.n277 VSUBS 0.006557f
C318 B.n278 VSUBS 0.006557f
C319 B.n279 VSUBS 0.006557f
C320 B.n280 VSUBS 0.006557f
C321 B.n281 VSUBS 0.006557f
C322 B.n282 VSUBS 0.006557f
C323 B.n283 VSUBS 0.006557f
C324 B.n284 VSUBS 0.006557f
C325 B.n285 VSUBS 0.006557f
C326 B.n286 VSUBS 0.006557f
C327 B.n287 VSUBS 0.006557f
C328 B.n288 VSUBS 0.006557f
C329 B.n289 VSUBS 0.006557f
C330 B.n290 VSUBS 0.006557f
C331 B.n291 VSUBS 0.006557f
C332 B.n292 VSUBS 0.006557f
C333 B.n293 VSUBS 0.006557f
C334 B.n294 VSUBS 0.006557f
C335 B.n295 VSUBS 0.006557f
C336 B.n296 VSUBS 0.006557f
C337 B.n297 VSUBS 0.006557f
C338 B.n298 VSUBS 0.006557f
C339 B.n299 VSUBS 0.006557f
C340 B.n300 VSUBS 0.006557f
C341 B.n301 VSUBS 0.006557f
C342 B.n302 VSUBS 0.006557f
C343 B.n303 VSUBS 0.006557f
C344 B.n304 VSUBS 0.006557f
C345 B.n305 VSUBS 0.006557f
C346 B.n306 VSUBS 0.006557f
C347 B.n307 VSUBS 0.006557f
C348 B.n308 VSUBS 0.006557f
C349 B.n309 VSUBS 0.006557f
C350 B.n310 VSUBS 0.006557f
C351 B.n311 VSUBS 0.006557f
C352 B.n312 VSUBS 0.006557f
C353 B.n313 VSUBS 0.006557f
C354 B.n314 VSUBS 0.006557f
C355 B.n315 VSUBS 0.006557f
C356 B.n316 VSUBS 0.006557f
C357 B.n317 VSUBS 0.006557f
C358 B.n318 VSUBS 0.006557f
C359 B.n319 VSUBS 0.006557f
C360 B.n320 VSUBS 0.006557f
C361 B.n321 VSUBS 0.006557f
C362 B.n322 VSUBS 0.006557f
C363 B.n323 VSUBS 0.006557f
C364 B.n324 VSUBS 0.006557f
C365 B.n325 VSUBS 0.006557f
C366 B.n326 VSUBS 0.014702f
C367 B.n327 VSUBS 0.015384f
C368 B.n328 VSUBS 0.014585f
C369 B.n329 VSUBS 0.006557f
C370 B.n330 VSUBS 0.006557f
C371 B.n331 VSUBS 0.006557f
C372 B.n332 VSUBS 0.006557f
C373 B.n333 VSUBS 0.006557f
C374 B.n334 VSUBS 0.006557f
C375 B.n335 VSUBS 0.006557f
C376 B.n336 VSUBS 0.006557f
C377 B.n337 VSUBS 0.006557f
C378 B.n338 VSUBS 0.006557f
C379 B.n339 VSUBS 0.006557f
C380 B.n340 VSUBS 0.006557f
C381 B.n341 VSUBS 0.006557f
C382 B.n342 VSUBS 0.006557f
C383 B.n343 VSUBS 0.006557f
C384 B.n344 VSUBS 0.006557f
C385 B.n345 VSUBS 0.006557f
C386 B.n346 VSUBS 0.006557f
C387 B.n347 VSUBS 0.006557f
C388 B.n348 VSUBS 0.006557f
C389 B.n349 VSUBS 0.006557f
C390 B.n350 VSUBS 0.006557f
C391 B.n351 VSUBS 0.006557f
C392 B.n352 VSUBS 0.006557f
C393 B.n353 VSUBS 0.006557f
C394 B.n354 VSUBS 0.006557f
C395 B.n355 VSUBS 0.006557f
C396 B.n356 VSUBS 0.006557f
C397 B.n357 VSUBS 0.006557f
C398 B.n358 VSUBS 0.006557f
C399 B.n359 VSUBS 0.006557f
C400 B.n360 VSUBS 0.006557f
C401 B.n361 VSUBS 0.006557f
C402 B.n362 VSUBS 0.006557f
C403 B.n363 VSUBS 0.006557f
C404 B.n364 VSUBS 0.006557f
C405 B.n365 VSUBS 0.006557f
C406 B.n366 VSUBS 0.006557f
C407 B.n367 VSUBS 0.006557f
C408 B.n368 VSUBS 0.006557f
C409 B.n369 VSUBS 0.006557f
C410 B.n370 VSUBS 0.006557f
C411 B.n371 VSUBS 0.006557f
C412 B.n372 VSUBS 0.006557f
C413 B.n373 VSUBS 0.006557f
C414 B.n374 VSUBS 0.006557f
C415 B.n375 VSUBS 0.006557f
C416 B.n376 VSUBS 0.006557f
C417 B.n377 VSUBS 0.006557f
C418 B.n378 VSUBS 0.006557f
C419 B.n379 VSUBS 0.006557f
C420 B.n380 VSUBS 0.006557f
C421 B.n381 VSUBS 0.006557f
C422 B.n382 VSUBS 0.006557f
C423 B.n383 VSUBS 0.014585f
C424 B.n384 VSUBS 0.015501f
C425 B.n385 VSUBS 0.015501f
C426 B.n386 VSUBS 0.006557f
C427 B.n387 VSUBS 0.006557f
C428 B.n388 VSUBS 0.006557f
C429 B.n389 VSUBS 0.006557f
C430 B.n390 VSUBS 0.006557f
C431 B.n391 VSUBS 0.006557f
C432 B.n392 VSUBS 0.006557f
C433 B.n393 VSUBS 0.006557f
C434 B.n394 VSUBS 0.006557f
C435 B.n395 VSUBS 0.006557f
C436 B.n396 VSUBS 0.006557f
C437 B.n397 VSUBS 0.006557f
C438 B.n398 VSUBS 0.006557f
C439 B.n399 VSUBS 0.006557f
C440 B.n400 VSUBS 0.006557f
C441 B.n401 VSUBS 0.006557f
C442 B.n402 VSUBS 0.006557f
C443 B.n403 VSUBS 0.006557f
C444 B.n404 VSUBS 0.006557f
C445 B.n405 VSUBS 0.006557f
C446 B.n406 VSUBS 0.006557f
C447 B.n407 VSUBS 0.006557f
C448 B.n408 VSUBS 0.006557f
C449 B.n409 VSUBS 0.006557f
C450 B.n410 VSUBS 0.006557f
C451 B.n411 VSUBS 0.006557f
C452 B.n412 VSUBS 0.006557f
C453 B.n413 VSUBS 0.006557f
C454 B.n414 VSUBS 0.006557f
C455 B.n415 VSUBS 0.006557f
C456 B.n416 VSUBS 0.006557f
C457 B.n417 VSUBS 0.006557f
C458 B.n418 VSUBS 0.006557f
C459 B.n419 VSUBS 0.006557f
C460 B.n420 VSUBS 0.006557f
C461 B.n421 VSUBS 0.006557f
C462 B.n422 VSUBS 0.006557f
C463 B.n423 VSUBS 0.006557f
C464 B.n424 VSUBS 0.006557f
C465 B.n425 VSUBS 0.006557f
C466 B.n426 VSUBS 0.006557f
C467 B.n427 VSUBS 0.006557f
C468 B.n428 VSUBS 0.006557f
C469 B.n429 VSUBS 0.006557f
C470 B.n430 VSUBS 0.006557f
C471 B.n431 VSUBS 0.006557f
C472 B.n432 VSUBS 0.006557f
C473 B.n433 VSUBS 0.006557f
C474 B.n434 VSUBS 0.006557f
C475 B.n435 VSUBS 0.006557f
C476 B.n436 VSUBS 0.006557f
C477 B.n437 VSUBS 0.006557f
C478 B.n438 VSUBS 0.006557f
C479 B.n439 VSUBS 0.006557f
C480 B.n440 VSUBS 0.006557f
C481 B.n441 VSUBS 0.006557f
C482 B.n442 VSUBS 0.006557f
C483 B.n443 VSUBS 0.006557f
C484 B.n444 VSUBS 0.006557f
C485 B.n445 VSUBS 0.006557f
C486 B.n446 VSUBS 0.006557f
C487 B.n447 VSUBS 0.006557f
C488 B.n448 VSUBS 0.006557f
C489 B.n449 VSUBS 0.006557f
C490 B.n450 VSUBS 0.006557f
C491 B.n451 VSUBS 0.006557f
C492 B.n452 VSUBS 0.004532f
C493 B.n453 VSUBS 0.015192f
C494 B.n454 VSUBS 0.005304f
C495 B.n455 VSUBS 0.006557f
C496 B.n456 VSUBS 0.006557f
C497 B.n457 VSUBS 0.006557f
C498 B.n458 VSUBS 0.006557f
C499 B.n459 VSUBS 0.006557f
C500 B.n460 VSUBS 0.006557f
C501 B.n461 VSUBS 0.006557f
C502 B.n462 VSUBS 0.006557f
C503 B.n463 VSUBS 0.006557f
C504 B.n464 VSUBS 0.006557f
C505 B.n465 VSUBS 0.006557f
C506 B.n466 VSUBS 0.005304f
C507 B.n467 VSUBS 0.006557f
C508 B.n468 VSUBS 0.006557f
C509 B.n469 VSUBS 0.004532f
C510 B.n470 VSUBS 0.006557f
C511 B.n471 VSUBS 0.006557f
C512 B.n472 VSUBS 0.006557f
C513 B.n473 VSUBS 0.006557f
C514 B.n474 VSUBS 0.006557f
C515 B.n475 VSUBS 0.006557f
C516 B.n476 VSUBS 0.006557f
C517 B.n477 VSUBS 0.006557f
C518 B.n478 VSUBS 0.006557f
C519 B.n479 VSUBS 0.006557f
C520 B.n480 VSUBS 0.006557f
C521 B.n481 VSUBS 0.006557f
C522 B.n482 VSUBS 0.006557f
C523 B.n483 VSUBS 0.006557f
C524 B.n484 VSUBS 0.006557f
C525 B.n485 VSUBS 0.006557f
C526 B.n486 VSUBS 0.006557f
C527 B.n487 VSUBS 0.006557f
C528 B.n488 VSUBS 0.006557f
C529 B.n489 VSUBS 0.006557f
C530 B.n490 VSUBS 0.006557f
C531 B.n491 VSUBS 0.006557f
C532 B.n492 VSUBS 0.006557f
C533 B.n493 VSUBS 0.006557f
C534 B.n494 VSUBS 0.006557f
C535 B.n495 VSUBS 0.006557f
C536 B.n496 VSUBS 0.006557f
C537 B.n497 VSUBS 0.006557f
C538 B.n498 VSUBS 0.006557f
C539 B.n499 VSUBS 0.006557f
C540 B.n500 VSUBS 0.006557f
C541 B.n501 VSUBS 0.006557f
C542 B.n502 VSUBS 0.006557f
C543 B.n503 VSUBS 0.006557f
C544 B.n504 VSUBS 0.006557f
C545 B.n505 VSUBS 0.006557f
C546 B.n506 VSUBS 0.006557f
C547 B.n507 VSUBS 0.006557f
C548 B.n508 VSUBS 0.006557f
C549 B.n509 VSUBS 0.006557f
C550 B.n510 VSUBS 0.006557f
C551 B.n511 VSUBS 0.006557f
C552 B.n512 VSUBS 0.006557f
C553 B.n513 VSUBS 0.006557f
C554 B.n514 VSUBS 0.006557f
C555 B.n515 VSUBS 0.006557f
C556 B.n516 VSUBS 0.006557f
C557 B.n517 VSUBS 0.006557f
C558 B.n518 VSUBS 0.006557f
C559 B.n519 VSUBS 0.006557f
C560 B.n520 VSUBS 0.006557f
C561 B.n521 VSUBS 0.006557f
C562 B.n522 VSUBS 0.006557f
C563 B.n523 VSUBS 0.006557f
C564 B.n524 VSUBS 0.006557f
C565 B.n525 VSUBS 0.006557f
C566 B.n526 VSUBS 0.006557f
C567 B.n527 VSUBS 0.006557f
C568 B.n528 VSUBS 0.006557f
C569 B.n529 VSUBS 0.006557f
C570 B.n530 VSUBS 0.006557f
C571 B.n531 VSUBS 0.006557f
C572 B.n532 VSUBS 0.006557f
C573 B.n533 VSUBS 0.006557f
C574 B.n534 VSUBS 0.006557f
C575 B.n535 VSUBS 0.006557f
C576 B.n536 VSUBS 0.015501f
C577 B.n537 VSUBS 0.014585f
C578 B.n538 VSUBS 0.014585f
C579 B.n539 VSUBS 0.006557f
C580 B.n540 VSUBS 0.006557f
C581 B.n541 VSUBS 0.006557f
C582 B.n542 VSUBS 0.006557f
C583 B.n543 VSUBS 0.006557f
C584 B.n544 VSUBS 0.006557f
C585 B.n545 VSUBS 0.006557f
C586 B.n546 VSUBS 0.006557f
C587 B.n547 VSUBS 0.006557f
C588 B.n548 VSUBS 0.006557f
C589 B.n549 VSUBS 0.006557f
C590 B.n550 VSUBS 0.006557f
C591 B.n551 VSUBS 0.006557f
C592 B.n552 VSUBS 0.006557f
C593 B.n553 VSUBS 0.006557f
C594 B.n554 VSUBS 0.006557f
C595 B.n555 VSUBS 0.006557f
C596 B.n556 VSUBS 0.006557f
C597 B.n557 VSUBS 0.006557f
C598 B.n558 VSUBS 0.006557f
C599 B.n559 VSUBS 0.006557f
C600 B.n560 VSUBS 0.006557f
C601 B.n561 VSUBS 0.006557f
C602 B.n562 VSUBS 0.006557f
C603 B.n563 VSUBS 0.008557f
C604 B.n564 VSUBS 0.009115f
C605 B.n565 VSUBS 0.018126f
C606 VDD2.n0 VSUBS 0.021672f
C607 VDD2.n1 VSUBS 0.020039f
C608 VDD2.n2 VSUBS 0.010768f
C609 VDD2.n3 VSUBS 0.025452f
C610 VDD2.n4 VSUBS 0.011401f
C611 VDD2.n5 VSUBS 0.020039f
C612 VDD2.n6 VSUBS 0.010768f
C613 VDD2.n7 VSUBS 0.025452f
C614 VDD2.n8 VSUBS 0.011401f
C615 VDD2.n9 VSUBS 0.020039f
C616 VDD2.n10 VSUBS 0.010768f
C617 VDD2.n11 VSUBS 0.025452f
C618 VDD2.n12 VSUBS 0.011401f
C619 VDD2.n13 VSUBS 0.020039f
C620 VDD2.n14 VSUBS 0.010768f
C621 VDD2.n15 VSUBS 0.025452f
C622 VDD2.n16 VSUBS 0.011401f
C623 VDD2.n17 VSUBS 0.020039f
C624 VDD2.n18 VSUBS 0.010768f
C625 VDD2.n19 VSUBS 0.025452f
C626 VDD2.n20 VSUBS 0.011401f
C627 VDD2.n21 VSUBS 1.13033f
C628 VDD2.n22 VSUBS 0.010768f
C629 VDD2.t0 VSUBS 0.054406f
C630 VDD2.n23 VSUBS 0.131565f
C631 VDD2.n24 VSUBS 0.016191f
C632 VDD2.n25 VSUBS 0.019089f
C633 VDD2.n26 VSUBS 0.025452f
C634 VDD2.n27 VSUBS 0.011401f
C635 VDD2.n28 VSUBS 0.010768f
C636 VDD2.n29 VSUBS 0.020039f
C637 VDD2.n30 VSUBS 0.020039f
C638 VDD2.n31 VSUBS 0.010768f
C639 VDD2.n32 VSUBS 0.011401f
C640 VDD2.n33 VSUBS 0.025452f
C641 VDD2.n34 VSUBS 0.025452f
C642 VDD2.n35 VSUBS 0.011401f
C643 VDD2.n36 VSUBS 0.010768f
C644 VDD2.n37 VSUBS 0.020039f
C645 VDD2.n38 VSUBS 0.020039f
C646 VDD2.n39 VSUBS 0.010768f
C647 VDD2.n40 VSUBS 0.011401f
C648 VDD2.n41 VSUBS 0.025452f
C649 VDD2.n42 VSUBS 0.025452f
C650 VDD2.n43 VSUBS 0.011401f
C651 VDD2.n44 VSUBS 0.010768f
C652 VDD2.n45 VSUBS 0.020039f
C653 VDD2.n46 VSUBS 0.020039f
C654 VDD2.n47 VSUBS 0.010768f
C655 VDD2.n48 VSUBS 0.011401f
C656 VDD2.n49 VSUBS 0.025452f
C657 VDD2.n50 VSUBS 0.025452f
C658 VDD2.n51 VSUBS 0.011401f
C659 VDD2.n52 VSUBS 0.010768f
C660 VDD2.n53 VSUBS 0.020039f
C661 VDD2.n54 VSUBS 0.020039f
C662 VDD2.n55 VSUBS 0.010768f
C663 VDD2.n56 VSUBS 0.011401f
C664 VDD2.n57 VSUBS 0.025452f
C665 VDD2.n58 VSUBS 0.025452f
C666 VDD2.n59 VSUBS 0.011401f
C667 VDD2.n60 VSUBS 0.010768f
C668 VDD2.n61 VSUBS 0.020039f
C669 VDD2.n62 VSUBS 0.020039f
C670 VDD2.n63 VSUBS 0.010768f
C671 VDD2.n64 VSUBS 0.011401f
C672 VDD2.n65 VSUBS 0.025452f
C673 VDD2.n66 VSUBS 0.063376f
C674 VDD2.n67 VSUBS 0.011401f
C675 VDD2.n68 VSUBS 0.021146f
C676 VDD2.n69 VSUBS 0.050699f
C677 VDD2.n70 VSUBS 0.567823f
C678 VDD2.n71 VSUBS 0.021672f
C679 VDD2.n72 VSUBS 0.020039f
C680 VDD2.n73 VSUBS 0.010768f
C681 VDD2.n74 VSUBS 0.025452f
C682 VDD2.n75 VSUBS 0.011401f
C683 VDD2.n76 VSUBS 0.020039f
C684 VDD2.n77 VSUBS 0.010768f
C685 VDD2.n78 VSUBS 0.025452f
C686 VDD2.n79 VSUBS 0.011401f
C687 VDD2.n80 VSUBS 0.020039f
C688 VDD2.n81 VSUBS 0.010768f
C689 VDD2.n82 VSUBS 0.025452f
C690 VDD2.n83 VSUBS 0.011401f
C691 VDD2.n84 VSUBS 0.020039f
C692 VDD2.n85 VSUBS 0.010768f
C693 VDD2.n86 VSUBS 0.025452f
C694 VDD2.n87 VSUBS 0.011401f
C695 VDD2.n88 VSUBS 0.020039f
C696 VDD2.n89 VSUBS 0.010768f
C697 VDD2.n90 VSUBS 0.025452f
C698 VDD2.n91 VSUBS 0.011401f
C699 VDD2.n92 VSUBS 1.13033f
C700 VDD2.n93 VSUBS 0.010768f
C701 VDD2.t1 VSUBS 0.054406f
C702 VDD2.n94 VSUBS 0.131565f
C703 VDD2.n95 VSUBS 0.016191f
C704 VDD2.n96 VSUBS 0.019089f
C705 VDD2.n97 VSUBS 0.025452f
C706 VDD2.n98 VSUBS 0.011401f
C707 VDD2.n99 VSUBS 0.010768f
C708 VDD2.n100 VSUBS 0.020039f
C709 VDD2.n101 VSUBS 0.020039f
C710 VDD2.n102 VSUBS 0.010768f
C711 VDD2.n103 VSUBS 0.011401f
C712 VDD2.n104 VSUBS 0.025452f
C713 VDD2.n105 VSUBS 0.025452f
C714 VDD2.n106 VSUBS 0.011401f
C715 VDD2.n107 VSUBS 0.010768f
C716 VDD2.n108 VSUBS 0.020039f
C717 VDD2.n109 VSUBS 0.020039f
C718 VDD2.n110 VSUBS 0.010768f
C719 VDD2.n111 VSUBS 0.011401f
C720 VDD2.n112 VSUBS 0.025452f
C721 VDD2.n113 VSUBS 0.025452f
C722 VDD2.n114 VSUBS 0.011401f
C723 VDD2.n115 VSUBS 0.010768f
C724 VDD2.n116 VSUBS 0.020039f
C725 VDD2.n117 VSUBS 0.020039f
C726 VDD2.n118 VSUBS 0.010768f
C727 VDD2.n119 VSUBS 0.011401f
C728 VDD2.n120 VSUBS 0.025452f
C729 VDD2.n121 VSUBS 0.025452f
C730 VDD2.n122 VSUBS 0.011401f
C731 VDD2.n123 VSUBS 0.010768f
C732 VDD2.n124 VSUBS 0.020039f
C733 VDD2.n125 VSUBS 0.020039f
C734 VDD2.n126 VSUBS 0.010768f
C735 VDD2.n127 VSUBS 0.011401f
C736 VDD2.n128 VSUBS 0.025452f
C737 VDD2.n129 VSUBS 0.025452f
C738 VDD2.n130 VSUBS 0.011401f
C739 VDD2.n131 VSUBS 0.010768f
C740 VDD2.n132 VSUBS 0.020039f
C741 VDD2.n133 VSUBS 0.020039f
C742 VDD2.n134 VSUBS 0.010768f
C743 VDD2.n135 VSUBS 0.011401f
C744 VDD2.n136 VSUBS 0.025452f
C745 VDD2.n137 VSUBS 0.063376f
C746 VDD2.n138 VSUBS 0.011401f
C747 VDD2.n139 VSUBS 0.021146f
C748 VDD2.n140 VSUBS 0.050699f
C749 VDD2.n141 VSUBS 0.062433f
C750 VDD2.n142 VSUBS 2.40043f
C751 VN.t1 VSUBS 3.08906f
C752 VN.t0 VSUBS 3.44182f
C753 VDD1.n0 VSUBS 0.022002f
C754 VDD1.n1 VSUBS 0.020344f
C755 VDD1.n2 VSUBS 0.010932f
C756 VDD1.n3 VSUBS 0.025839f
C757 VDD1.n4 VSUBS 0.011575f
C758 VDD1.n5 VSUBS 0.020344f
C759 VDD1.n6 VSUBS 0.010932f
C760 VDD1.n7 VSUBS 0.025839f
C761 VDD1.n8 VSUBS 0.011575f
C762 VDD1.n9 VSUBS 0.020344f
C763 VDD1.n10 VSUBS 0.010932f
C764 VDD1.n11 VSUBS 0.025839f
C765 VDD1.n12 VSUBS 0.011575f
C766 VDD1.n13 VSUBS 0.020344f
C767 VDD1.n14 VSUBS 0.010932f
C768 VDD1.n15 VSUBS 0.025839f
C769 VDD1.n16 VSUBS 0.011575f
C770 VDD1.n17 VSUBS 0.020344f
C771 VDD1.n18 VSUBS 0.010932f
C772 VDD1.n19 VSUBS 0.025839f
C773 VDD1.n20 VSUBS 0.011575f
C774 VDD1.n21 VSUBS 1.14754f
C775 VDD1.n22 VSUBS 0.010932f
C776 VDD1.t1 VSUBS 0.055235f
C777 VDD1.n23 VSUBS 0.133568f
C778 VDD1.n24 VSUBS 0.016438f
C779 VDD1.n25 VSUBS 0.01938f
C780 VDD1.n26 VSUBS 0.025839f
C781 VDD1.n27 VSUBS 0.011575f
C782 VDD1.n28 VSUBS 0.010932f
C783 VDD1.n29 VSUBS 0.020344f
C784 VDD1.n30 VSUBS 0.020344f
C785 VDD1.n31 VSUBS 0.010932f
C786 VDD1.n32 VSUBS 0.011575f
C787 VDD1.n33 VSUBS 0.025839f
C788 VDD1.n34 VSUBS 0.025839f
C789 VDD1.n35 VSUBS 0.011575f
C790 VDD1.n36 VSUBS 0.010932f
C791 VDD1.n37 VSUBS 0.020344f
C792 VDD1.n38 VSUBS 0.020344f
C793 VDD1.n39 VSUBS 0.010932f
C794 VDD1.n40 VSUBS 0.011575f
C795 VDD1.n41 VSUBS 0.025839f
C796 VDD1.n42 VSUBS 0.025839f
C797 VDD1.n43 VSUBS 0.011575f
C798 VDD1.n44 VSUBS 0.010932f
C799 VDD1.n45 VSUBS 0.020344f
C800 VDD1.n46 VSUBS 0.020344f
C801 VDD1.n47 VSUBS 0.010932f
C802 VDD1.n48 VSUBS 0.011575f
C803 VDD1.n49 VSUBS 0.025839f
C804 VDD1.n50 VSUBS 0.025839f
C805 VDD1.n51 VSUBS 0.011575f
C806 VDD1.n52 VSUBS 0.010932f
C807 VDD1.n53 VSUBS 0.020344f
C808 VDD1.n54 VSUBS 0.020344f
C809 VDD1.n55 VSUBS 0.010932f
C810 VDD1.n56 VSUBS 0.011575f
C811 VDD1.n57 VSUBS 0.025839f
C812 VDD1.n58 VSUBS 0.025839f
C813 VDD1.n59 VSUBS 0.011575f
C814 VDD1.n60 VSUBS 0.010932f
C815 VDD1.n61 VSUBS 0.020344f
C816 VDD1.n62 VSUBS 0.020344f
C817 VDD1.n63 VSUBS 0.010932f
C818 VDD1.n64 VSUBS 0.011575f
C819 VDD1.n65 VSUBS 0.025839f
C820 VDD1.n66 VSUBS 0.064341f
C821 VDD1.n67 VSUBS 0.011575f
C822 VDD1.n68 VSUBS 0.021468f
C823 VDD1.n69 VSUBS 0.051471f
C824 VDD1.n70 VSUBS 0.063975f
C825 VDD1.n71 VSUBS 0.022002f
C826 VDD1.n72 VSUBS 0.020344f
C827 VDD1.n73 VSUBS 0.010932f
C828 VDD1.n74 VSUBS 0.025839f
C829 VDD1.n75 VSUBS 0.011575f
C830 VDD1.n76 VSUBS 0.020344f
C831 VDD1.n77 VSUBS 0.010932f
C832 VDD1.n78 VSUBS 0.025839f
C833 VDD1.n79 VSUBS 0.011575f
C834 VDD1.n80 VSUBS 0.020344f
C835 VDD1.n81 VSUBS 0.010932f
C836 VDD1.n82 VSUBS 0.025839f
C837 VDD1.n83 VSUBS 0.011575f
C838 VDD1.n84 VSUBS 0.020344f
C839 VDD1.n85 VSUBS 0.010932f
C840 VDD1.n86 VSUBS 0.025839f
C841 VDD1.n87 VSUBS 0.011575f
C842 VDD1.n88 VSUBS 0.020344f
C843 VDD1.n89 VSUBS 0.010932f
C844 VDD1.n90 VSUBS 0.025839f
C845 VDD1.n91 VSUBS 0.011575f
C846 VDD1.n92 VSUBS 1.14754f
C847 VDD1.n93 VSUBS 0.010932f
C848 VDD1.t0 VSUBS 0.055235f
C849 VDD1.n94 VSUBS 0.133568f
C850 VDD1.n95 VSUBS 0.016438f
C851 VDD1.n96 VSUBS 0.01938f
C852 VDD1.n97 VSUBS 0.025839f
C853 VDD1.n98 VSUBS 0.011575f
C854 VDD1.n99 VSUBS 0.010932f
C855 VDD1.n100 VSUBS 0.020344f
C856 VDD1.n101 VSUBS 0.020344f
C857 VDD1.n102 VSUBS 0.010932f
C858 VDD1.n103 VSUBS 0.011575f
C859 VDD1.n104 VSUBS 0.025839f
C860 VDD1.n105 VSUBS 0.025839f
C861 VDD1.n106 VSUBS 0.011575f
C862 VDD1.n107 VSUBS 0.010932f
C863 VDD1.n108 VSUBS 0.020344f
C864 VDD1.n109 VSUBS 0.020344f
C865 VDD1.n110 VSUBS 0.010932f
C866 VDD1.n111 VSUBS 0.011575f
C867 VDD1.n112 VSUBS 0.025839f
C868 VDD1.n113 VSUBS 0.025839f
C869 VDD1.n114 VSUBS 0.011575f
C870 VDD1.n115 VSUBS 0.010932f
C871 VDD1.n116 VSUBS 0.020344f
C872 VDD1.n117 VSUBS 0.020344f
C873 VDD1.n118 VSUBS 0.010932f
C874 VDD1.n119 VSUBS 0.011575f
C875 VDD1.n120 VSUBS 0.025839f
C876 VDD1.n121 VSUBS 0.025839f
C877 VDD1.n122 VSUBS 0.011575f
C878 VDD1.n123 VSUBS 0.010932f
C879 VDD1.n124 VSUBS 0.020344f
C880 VDD1.n125 VSUBS 0.020344f
C881 VDD1.n126 VSUBS 0.010932f
C882 VDD1.n127 VSUBS 0.011575f
C883 VDD1.n128 VSUBS 0.025839f
C884 VDD1.n129 VSUBS 0.025839f
C885 VDD1.n130 VSUBS 0.011575f
C886 VDD1.n131 VSUBS 0.010932f
C887 VDD1.n132 VSUBS 0.020344f
C888 VDD1.n133 VSUBS 0.020344f
C889 VDD1.n134 VSUBS 0.010932f
C890 VDD1.n135 VSUBS 0.011575f
C891 VDD1.n136 VSUBS 0.025839f
C892 VDD1.n137 VSUBS 0.064341f
C893 VDD1.n138 VSUBS 0.011575f
C894 VDD1.n139 VSUBS 0.021468f
C895 VDD1.n140 VSUBS 0.051471f
C896 VDD1.n141 VSUBS 0.608204f
C897 VTAIL.n0 VSUBS 0.030903f
C898 VTAIL.n1 VSUBS 0.028575f
C899 VTAIL.n2 VSUBS 0.015355f
C900 VTAIL.n3 VSUBS 0.036293f
C901 VTAIL.n4 VSUBS 0.016258f
C902 VTAIL.n5 VSUBS 0.028575f
C903 VTAIL.n6 VSUBS 0.015355f
C904 VTAIL.n7 VSUBS 0.036293f
C905 VTAIL.n8 VSUBS 0.016258f
C906 VTAIL.n9 VSUBS 0.028575f
C907 VTAIL.n10 VSUBS 0.015355f
C908 VTAIL.n11 VSUBS 0.036293f
C909 VTAIL.n12 VSUBS 0.016258f
C910 VTAIL.n13 VSUBS 0.028575f
C911 VTAIL.n14 VSUBS 0.015355f
C912 VTAIL.n15 VSUBS 0.036293f
C913 VTAIL.n16 VSUBS 0.016258f
C914 VTAIL.n17 VSUBS 0.028575f
C915 VTAIL.n18 VSUBS 0.015355f
C916 VTAIL.n19 VSUBS 0.036293f
C917 VTAIL.n20 VSUBS 0.016258f
C918 VTAIL.n21 VSUBS 1.61182f
C919 VTAIL.n22 VSUBS 0.015355f
C920 VTAIL.t2 VSUBS 0.077582f
C921 VTAIL.n23 VSUBS 0.187607f
C922 VTAIL.n24 VSUBS 0.023088f
C923 VTAIL.n25 VSUBS 0.02722f
C924 VTAIL.n26 VSUBS 0.036293f
C925 VTAIL.n27 VSUBS 0.016258f
C926 VTAIL.n28 VSUBS 0.015355f
C927 VTAIL.n29 VSUBS 0.028575f
C928 VTAIL.n30 VSUBS 0.028575f
C929 VTAIL.n31 VSUBS 0.015355f
C930 VTAIL.n32 VSUBS 0.016258f
C931 VTAIL.n33 VSUBS 0.036293f
C932 VTAIL.n34 VSUBS 0.036293f
C933 VTAIL.n35 VSUBS 0.016258f
C934 VTAIL.n36 VSUBS 0.015355f
C935 VTAIL.n37 VSUBS 0.028575f
C936 VTAIL.n38 VSUBS 0.028575f
C937 VTAIL.n39 VSUBS 0.015355f
C938 VTAIL.n40 VSUBS 0.016258f
C939 VTAIL.n41 VSUBS 0.036293f
C940 VTAIL.n42 VSUBS 0.036293f
C941 VTAIL.n43 VSUBS 0.016258f
C942 VTAIL.n44 VSUBS 0.015355f
C943 VTAIL.n45 VSUBS 0.028575f
C944 VTAIL.n46 VSUBS 0.028575f
C945 VTAIL.n47 VSUBS 0.015355f
C946 VTAIL.n48 VSUBS 0.016258f
C947 VTAIL.n49 VSUBS 0.036293f
C948 VTAIL.n50 VSUBS 0.036293f
C949 VTAIL.n51 VSUBS 0.016258f
C950 VTAIL.n52 VSUBS 0.015355f
C951 VTAIL.n53 VSUBS 0.028575f
C952 VTAIL.n54 VSUBS 0.028575f
C953 VTAIL.n55 VSUBS 0.015355f
C954 VTAIL.n56 VSUBS 0.016258f
C955 VTAIL.n57 VSUBS 0.036293f
C956 VTAIL.n58 VSUBS 0.036293f
C957 VTAIL.n59 VSUBS 0.016258f
C958 VTAIL.n60 VSUBS 0.015355f
C959 VTAIL.n61 VSUBS 0.028575f
C960 VTAIL.n62 VSUBS 0.028575f
C961 VTAIL.n63 VSUBS 0.015355f
C962 VTAIL.n64 VSUBS 0.016258f
C963 VTAIL.n65 VSUBS 0.036293f
C964 VTAIL.n66 VSUBS 0.090372f
C965 VTAIL.n67 VSUBS 0.016258f
C966 VTAIL.n68 VSUBS 0.030153f
C967 VTAIL.n69 VSUBS 0.072295f
C968 VTAIL.n70 VSUBS 0.069341f
C969 VTAIL.n71 VSUBS 1.84127f
C970 VTAIL.n72 VSUBS 0.030903f
C971 VTAIL.n73 VSUBS 0.028575f
C972 VTAIL.n74 VSUBS 0.015355f
C973 VTAIL.n75 VSUBS 0.036293f
C974 VTAIL.n76 VSUBS 0.016258f
C975 VTAIL.n77 VSUBS 0.028575f
C976 VTAIL.n78 VSUBS 0.015355f
C977 VTAIL.n79 VSUBS 0.036293f
C978 VTAIL.n80 VSUBS 0.016258f
C979 VTAIL.n81 VSUBS 0.028575f
C980 VTAIL.n82 VSUBS 0.015355f
C981 VTAIL.n83 VSUBS 0.036293f
C982 VTAIL.n84 VSUBS 0.016258f
C983 VTAIL.n85 VSUBS 0.028575f
C984 VTAIL.n86 VSUBS 0.015355f
C985 VTAIL.n87 VSUBS 0.036293f
C986 VTAIL.n88 VSUBS 0.016258f
C987 VTAIL.n89 VSUBS 0.028575f
C988 VTAIL.n90 VSUBS 0.015355f
C989 VTAIL.n91 VSUBS 0.036293f
C990 VTAIL.n92 VSUBS 0.016258f
C991 VTAIL.n93 VSUBS 1.61182f
C992 VTAIL.n94 VSUBS 0.015355f
C993 VTAIL.t1 VSUBS 0.077582f
C994 VTAIL.n95 VSUBS 0.187607f
C995 VTAIL.n96 VSUBS 0.023088f
C996 VTAIL.n97 VSUBS 0.02722f
C997 VTAIL.n98 VSUBS 0.036293f
C998 VTAIL.n99 VSUBS 0.016258f
C999 VTAIL.n100 VSUBS 0.015355f
C1000 VTAIL.n101 VSUBS 0.028575f
C1001 VTAIL.n102 VSUBS 0.028575f
C1002 VTAIL.n103 VSUBS 0.015355f
C1003 VTAIL.n104 VSUBS 0.016258f
C1004 VTAIL.n105 VSUBS 0.036293f
C1005 VTAIL.n106 VSUBS 0.036293f
C1006 VTAIL.n107 VSUBS 0.016258f
C1007 VTAIL.n108 VSUBS 0.015355f
C1008 VTAIL.n109 VSUBS 0.028575f
C1009 VTAIL.n110 VSUBS 0.028575f
C1010 VTAIL.n111 VSUBS 0.015355f
C1011 VTAIL.n112 VSUBS 0.016258f
C1012 VTAIL.n113 VSUBS 0.036293f
C1013 VTAIL.n114 VSUBS 0.036293f
C1014 VTAIL.n115 VSUBS 0.016258f
C1015 VTAIL.n116 VSUBS 0.015355f
C1016 VTAIL.n117 VSUBS 0.028575f
C1017 VTAIL.n118 VSUBS 0.028575f
C1018 VTAIL.n119 VSUBS 0.015355f
C1019 VTAIL.n120 VSUBS 0.016258f
C1020 VTAIL.n121 VSUBS 0.036293f
C1021 VTAIL.n122 VSUBS 0.036293f
C1022 VTAIL.n123 VSUBS 0.016258f
C1023 VTAIL.n124 VSUBS 0.015355f
C1024 VTAIL.n125 VSUBS 0.028575f
C1025 VTAIL.n126 VSUBS 0.028575f
C1026 VTAIL.n127 VSUBS 0.015355f
C1027 VTAIL.n128 VSUBS 0.016258f
C1028 VTAIL.n129 VSUBS 0.036293f
C1029 VTAIL.n130 VSUBS 0.036293f
C1030 VTAIL.n131 VSUBS 0.016258f
C1031 VTAIL.n132 VSUBS 0.015355f
C1032 VTAIL.n133 VSUBS 0.028575f
C1033 VTAIL.n134 VSUBS 0.028575f
C1034 VTAIL.n135 VSUBS 0.015355f
C1035 VTAIL.n136 VSUBS 0.016258f
C1036 VTAIL.n137 VSUBS 0.036293f
C1037 VTAIL.n138 VSUBS 0.090372f
C1038 VTAIL.n139 VSUBS 0.016258f
C1039 VTAIL.n140 VSUBS 0.030153f
C1040 VTAIL.n141 VSUBS 0.072295f
C1041 VTAIL.n142 VSUBS 0.069341f
C1042 VTAIL.n143 VSUBS 1.87103f
C1043 VTAIL.n144 VSUBS 0.030903f
C1044 VTAIL.n145 VSUBS 0.028575f
C1045 VTAIL.n146 VSUBS 0.015355f
C1046 VTAIL.n147 VSUBS 0.036293f
C1047 VTAIL.n148 VSUBS 0.016258f
C1048 VTAIL.n149 VSUBS 0.028575f
C1049 VTAIL.n150 VSUBS 0.015355f
C1050 VTAIL.n151 VSUBS 0.036293f
C1051 VTAIL.n152 VSUBS 0.016258f
C1052 VTAIL.n153 VSUBS 0.028575f
C1053 VTAIL.n154 VSUBS 0.015355f
C1054 VTAIL.n155 VSUBS 0.036293f
C1055 VTAIL.n156 VSUBS 0.016258f
C1056 VTAIL.n157 VSUBS 0.028575f
C1057 VTAIL.n158 VSUBS 0.015355f
C1058 VTAIL.n159 VSUBS 0.036293f
C1059 VTAIL.n160 VSUBS 0.016258f
C1060 VTAIL.n161 VSUBS 0.028575f
C1061 VTAIL.n162 VSUBS 0.015355f
C1062 VTAIL.n163 VSUBS 0.036293f
C1063 VTAIL.n164 VSUBS 0.016258f
C1064 VTAIL.n165 VSUBS 1.61182f
C1065 VTAIL.n166 VSUBS 0.015355f
C1066 VTAIL.t3 VSUBS 0.077582f
C1067 VTAIL.n167 VSUBS 0.187607f
C1068 VTAIL.n168 VSUBS 0.023088f
C1069 VTAIL.n169 VSUBS 0.02722f
C1070 VTAIL.n170 VSUBS 0.036293f
C1071 VTAIL.n171 VSUBS 0.016258f
C1072 VTAIL.n172 VSUBS 0.015355f
C1073 VTAIL.n173 VSUBS 0.028575f
C1074 VTAIL.n174 VSUBS 0.028575f
C1075 VTAIL.n175 VSUBS 0.015355f
C1076 VTAIL.n176 VSUBS 0.016258f
C1077 VTAIL.n177 VSUBS 0.036293f
C1078 VTAIL.n178 VSUBS 0.036293f
C1079 VTAIL.n179 VSUBS 0.016258f
C1080 VTAIL.n180 VSUBS 0.015355f
C1081 VTAIL.n181 VSUBS 0.028575f
C1082 VTAIL.n182 VSUBS 0.028575f
C1083 VTAIL.n183 VSUBS 0.015355f
C1084 VTAIL.n184 VSUBS 0.016258f
C1085 VTAIL.n185 VSUBS 0.036293f
C1086 VTAIL.n186 VSUBS 0.036293f
C1087 VTAIL.n187 VSUBS 0.016258f
C1088 VTAIL.n188 VSUBS 0.015355f
C1089 VTAIL.n189 VSUBS 0.028575f
C1090 VTAIL.n190 VSUBS 0.028575f
C1091 VTAIL.n191 VSUBS 0.015355f
C1092 VTAIL.n192 VSUBS 0.016258f
C1093 VTAIL.n193 VSUBS 0.036293f
C1094 VTAIL.n194 VSUBS 0.036293f
C1095 VTAIL.n195 VSUBS 0.016258f
C1096 VTAIL.n196 VSUBS 0.015355f
C1097 VTAIL.n197 VSUBS 0.028575f
C1098 VTAIL.n198 VSUBS 0.028575f
C1099 VTAIL.n199 VSUBS 0.015355f
C1100 VTAIL.n200 VSUBS 0.016258f
C1101 VTAIL.n201 VSUBS 0.036293f
C1102 VTAIL.n202 VSUBS 0.036293f
C1103 VTAIL.n203 VSUBS 0.016258f
C1104 VTAIL.n204 VSUBS 0.015355f
C1105 VTAIL.n205 VSUBS 0.028575f
C1106 VTAIL.n206 VSUBS 0.028575f
C1107 VTAIL.n207 VSUBS 0.015355f
C1108 VTAIL.n208 VSUBS 0.016258f
C1109 VTAIL.n209 VSUBS 0.036293f
C1110 VTAIL.n210 VSUBS 0.090372f
C1111 VTAIL.n211 VSUBS 0.016258f
C1112 VTAIL.n212 VSUBS 0.030153f
C1113 VTAIL.n213 VSUBS 0.072295f
C1114 VTAIL.n214 VSUBS 0.069341f
C1115 VTAIL.n215 VSUBS 1.73054f
C1116 VTAIL.n216 VSUBS 0.030903f
C1117 VTAIL.n217 VSUBS 0.028575f
C1118 VTAIL.n218 VSUBS 0.015355f
C1119 VTAIL.n219 VSUBS 0.036293f
C1120 VTAIL.n220 VSUBS 0.016258f
C1121 VTAIL.n221 VSUBS 0.028575f
C1122 VTAIL.n222 VSUBS 0.015355f
C1123 VTAIL.n223 VSUBS 0.036293f
C1124 VTAIL.n224 VSUBS 0.016258f
C1125 VTAIL.n225 VSUBS 0.028575f
C1126 VTAIL.n226 VSUBS 0.015355f
C1127 VTAIL.n227 VSUBS 0.036293f
C1128 VTAIL.n228 VSUBS 0.016258f
C1129 VTAIL.n229 VSUBS 0.028575f
C1130 VTAIL.n230 VSUBS 0.015355f
C1131 VTAIL.n231 VSUBS 0.036293f
C1132 VTAIL.n232 VSUBS 0.016258f
C1133 VTAIL.n233 VSUBS 0.028575f
C1134 VTAIL.n234 VSUBS 0.015355f
C1135 VTAIL.n235 VSUBS 0.036293f
C1136 VTAIL.n236 VSUBS 0.016258f
C1137 VTAIL.n237 VSUBS 1.61182f
C1138 VTAIL.n238 VSUBS 0.015355f
C1139 VTAIL.t0 VSUBS 0.077582f
C1140 VTAIL.n239 VSUBS 0.187607f
C1141 VTAIL.n240 VSUBS 0.023088f
C1142 VTAIL.n241 VSUBS 0.02722f
C1143 VTAIL.n242 VSUBS 0.036293f
C1144 VTAIL.n243 VSUBS 0.016258f
C1145 VTAIL.n244 VSUBS 0.015355f
C1146 VTAIL.n245 VSUBS 0.028575f
C1147 VTAIL.n246 VSUBS 0.028575f
C1148 VTAIL.n247 VSUBS 0.015355f
C1149 VTAIL.n248 VSUBS 0.016258f
C1150 VTAIL.n249 VSUBS 0.036293f
C1151 VTAIL.n250 VSUBS 0.036293f
C1152 VTAIL.n251 VSUBS 0.016258f
C1153 VTAIL.n252 VSUBS 0.015355f
C1154 VTAIL.n253 VSUBS 0.028575f
C1155 VTAIL.n254 VSUBS 0.028575f
C1156 VTAIL.n255 VSUBS 0.015355f
C1157 VTAIL.n256 VSUBS 0.016258f
C1158 VTAIL.n257 VSUBS 0.036293f
C1159 VTAIL.n258 VSUBS 0.036293f
C1160 VTAIL.n259 VSUBS 0.016258f
C1161 VTAIL.n260 VSUBS 0.015355f
C1162 VTAIL.n261 VSUBS 0.028575f
C1163 VTAIL.n262 VSUBS 0.028575f
C1164 VTAIL.n263 VSUBS 0.015355f
C1165 VTAIL.n264 VSUBS 0.016258f
C1166 VTAIL.n265 VSUBS 0.036293f
C1167 VTAIL.n266 VSUBS 0.036293f
C1168 VTAIL.n267 VSUBS 0.016258f
C1169 VTAIL.n268 VSUBS 0.015355f
C1170 VTAIL.n269 VSUBS 0.028575f
C1171 VTAIL.n270 VSUBS 0.028575f
C1172 VTAIL.n271 VSUBS 0.015355f
C1173 VTAIL.n272 VSUBS 0.016258f
C1174 VTAIL.n273 VSUBS 0.036293f
C1175 VTAIL.n274 VSUBS 0.036293f
C1176 VTAIL.n275 VSUBS 0.016258f
C1177 VTAIL.n276 VSUBS 0.015355f
C1178 VTAIL.n277 VSUBS 0.028575f
C1179 VTAIL.n278 VSUBS 0.028575f
C1180 VTAIL.n279 VSUBS 0.015355f
C1181 VTAIL.n280 VSUBS 0.016258f
C1182 VTAIL.n281 VSUBS 0.036293f
C1183 VTAIL.n282 VSUBS 0.090372f
C1184 VTAIL.n283 VSUBS 0.016258f
C1185 VTAIL.n284 VSUBS 0.030153f
C1186 VTAIL.n285 VSUBS 0.072295f
C1187 VTAIL.n286 VSUBS 0.069341f
C1188 VTAIL.n287 VSUBS 1.6468f
C1189 VP.t0 VSUBS 3.56816f
C1190 VP.t1 VSUBS 3.20704f
C1191 VP.n0 VSUBS 5.97123f
.ends

