* NGSPICE file created from diff_pair_sample_1276.ext - technology: sky130A

.subckt diff_pair_sample_1276 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t0 w_n1990_n3046# sky130_fd_pr__pfet_01v8 ad=4.0521 pd=21.56 as=1.71435 ps=10.72 w=10.39 l=1.37
X1 B.t11 B.t9 B.t10 w_n1990_n3046# sky130_fd_pr__pfet_01v8 ad=4.0521 pd=21.56 as=0 ps=0 w=10.39 l=1.37
X2 VTAIL.t3 VP.t0 VDD1.t3 w_n1990_n3046# sky130_fd_pr__pfet_01v8 ad=4.0521 pd=21.56 as=1.71435 ps=10.72 w=10.39 l=1.37
X3 VDD2.t3 VN.t1 VTAIL.t6 w_n1990_n3046# sky130_fd_pr__pfet_01v8 ad=1.71435 pd=10.72 as=4.0521 ps=21.56 w=10.39 l=1.37
X4 B.t8 B.t6 B.t7 w_n1990_n3046# sky130_fd_pr__pfet_01v8 ad=4.0521 pd=21.56 as=0 ps=0 w=10.39 l=1.37
X5 VTAIL.t5 VN.t2 VDD2.t2 w_n1990_n3046# sky130_fd_pr__pfet_01v8 ad=4.0521 pd=21.56 as=1.71435 ps=10.72 w=10.39 l=1.37
X6 VDD1.t2 VP.t1 VTAIL.t2 w_n1990_n3046# sky130_fd_pr__pfet_01v8 ad=1.71435 pd=10.72 as=4.0521 ps=21.56 w=10.39 l=1.37
X7 B.t5 B.t3 B.t4 w_n1990_n3046# sky130_fd_pr__pfet_01v8 ad=4.0521 pd=21.56 as=0 ps=0 w=10.39 l=1.37
X8 B.t2 B.t0 B.t1 w_n1990_n3046# sky130_fd_pr__pfet_01v8 ad=4.0521 pd=21.56 as=0 ps=0 w=10.39 l=1.37
X9 VDD2.t1 VN.t3 VTAIL.t4 w_n1990_n3046# sky130_fd_pr__pfet_01v8 ad=1.71435 pd=10.72 as=4.0521 ps=21.56 w=10.39 l=1.37
X10 VTAIL.t1 VP.t2 VDD1.t1 w_n1990_n3046# sky130_fd_pr__pfet_01v8 ad=4.0521 pd=21.56 as=1.71435 ps=10.72 w=10.39 l=1.37
X11 VDD1.t0 VP.t3 VTAIL.t0 w_n1990_n3046# sky130_fd_pr__pfet_01v8 ad=1.71435 pd=10.72 as=4.0521 ps=21.56 w=10.39 l=1.37
R0 VN.n0 VN.t0 221.192
R1 VN.n1 VN.t1 221.192
R2 VN.n0 VN.t3 220.96
R3 VN.n1 VN.t2 220.96
R4 VN VN.n1 59.3171
R5 VN VN.n0 17.6391
R6 VDD2.n2 VDD2.n0 114.894
R7 VDD2.n2 VDD2.n1 77.8261
R8 VDD2.n1 VDD2.t2 3.12899
R9 VDD2.n1 VDD2.t3 3.12899
R10 VDD2.n0 VDD2.t0 3.12899
R11 VDD2.n0 VDD2.t1 3.12899
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t1 64.276
R14 VTAIL.n4 VTAIL.t6 64.276
R15 VTAIL.n3 VTAIL.t5 64.276
R16 VTAIL.n6 VTAIL.t0 64.2757
R17 VTAIL.n7 VTAIL.t4 64.2757
R18 VTAIL.n0 VTAIL.t7 64.2757
R19 VTAIL.n1 VTAIL.t2 64.2757
R20 VTAIL.n2 VTAIL.t3 64.2757
R21 VTAIL.n7 VTAIL.n6 22.7893
R22 VTAIL.n3 VTAIL.n2 22.7893
R23 VTAIL.n4 VTAIL.n3 1.46602
R24 VTAIL.n6 VTAIL.n5 1.46602
R25 VTAIL.n2 VTAIL.n1 1.46602
R26 VTAIL VTAIL.n0 0.791448
R27 VTAIL VTAIL.n7 0.675069
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 B.n370 B.n59 585
R31 B.n372 B.n371 585
R32 B.n373 B.n58 585
R33 B.n375 B.n374 585
R34 B.n376 B.n57 585
R35 B.n378 B.n377 585
R36 B.n379 B.n56 585
R37 B.n381 B.n380 585
R38 B.n382 B.n55 585
R39 B.n384 B.n383 585
R40 B.n385 B.n54 585
R41 B.n387 B.n386 585
R42 B.n388 B.n53 585
R43 B.n390 B.n389 585
R44 B.n391 B.n52 585
R45 B.n393 B.n392 585
R46 B.n394 B.n51 585
R47 B.n396 B.n395 585
R48 B.n397 B.n50 585
R49 B.n399 B.n398 585
R50 B.n400 B.n49 585
R51 B.n402 B.n401 585
R52 B.n403 B.n48 585
R53 B.n405 B.n404 585
R54 B.n406 B.n47 585
R55 B.n408 B.n407 585
R56 B.n409 B.n46 585
R57 B.n411 B.n410 585
R58 B.n412 B.n45 585
R59 B.n414 B.n413 585
R60 B.n415 B.n44 585
R61 B.n417 B.n416 585
R62 B.n418 B.n43 585
R63 B.n420 B.n419 585
R64 B.n421 B.n42 585
R65 B.n423 B.n422 585
R66 B.n424 B.n39 585
R67 B.n427 B.n426 585
R68 B.n428 B.n38 585
R69 B.n430 B.n429 585
R70 B.n431 B.n37 585
R71 B.n433 B.n432 585
R72 B.n434 B.n36 585
R73 B.n436 B.n435 585
R74 B.n437 B.n35 585
R75 B.n439 B.n438 585
R76 B.n441 B.n440 585
R77 B.n442 B.n31 585
R78 B.n444 B.n443 585
R79 B.n445 B.n30 585
R80 B.n447 B.n446 585
R81 B.n448 B.n29 585
R82 B.n450 B.n449 585
R83 B.n451 B.n28 585
R84 B.n453 B.n452 585
R85 B.n454 B.n27 585
R86 B.n456 B.n455 585
R87 B.n457 B.n26 585
R88 B.n459 B.n458 585
R89 B.n460 B.n25 585
R90 B.n462 B.n461 585
R91 B.n463 B.n24 585
R92 B.n465 B.n464 585
R93 B.n466 B.n23 585
R94 B.n468 B.n467 585
R95 B.n469 B.n22 585
R96 B.n471 B.n470 585
R97 B.n472 B.n21 585
R98 B.n474 B.n473 585
R99 B.n475 B.n20 585
R100 B.n477 B.n476 585
R101 B.n478 B.n19 585
R102 B.n480 B.n479 585
R103 B.n481 B.n18 585
R104 B.n483 B.n482 585
R105 B.n484 B.n17 585
R106 B.n486 B.n485 585
R107 B.n487 B.n16 585
R108 B.n489 B.n488 585
R109 B.n490 B.n15 585
R110 B.n492 B.n491 585
R111 B.n493 B.n14 585
R112 B.n495 B.n494 585
R113 B.n369 B.n368 585
R114 B.n367 B.n60 585
R115 B.n366 B.n365 585
R116 B.n364 B.n61 585
R117 B.n363 B.n362 585
R118 B.n361 B.n62 585
R119 B.n360 B.n359 585
R120 B.n358 B.n63 585
R121 B.n357 B.n356 585
R122 B.n355 B.n64 585
R123 B.n354 B.n353 585
R124 B.n352 B.n65 585
R125 B.n351 B.n350 585
R126 B.n349 B.n66 585
R127 B.n348 B.n347 585
R128 B.n346 B.n67 585
R129 B.n345 B.n344 585
R130 B.n343 B.n68 585
R131 B.n342 B.n341 585
R132 B.n340 B.n69 585
R133 B.n339 B.n338 585
R134 B.n337 B.n70 585
R135 B.n336 B.n335 585
R136 B.n334 B.n71 585
R137 B.n333 B.n332 585
R138 B.n331 B.n72 585
R139 B.n330 B.n329 585
R140 B.n328 B.n73 585
R141 B.n327 B.n326 585
R142 B.n325 B.n74 585
R143 B.n324 B.n323 585
R144 B.n322 B.n75 585
R145 B.n321 B.n320 585
R146 B.n319 B.n76 585
R147 B.n318 B.n317 585
R148 B.n316 B.n77 585
R149 B.n315 B.n314 585
R150 B.n313 B.n78 585
R151 B.n312 B.n311 585
R152 B.n310 B.n79 585
R153 B.n309 B.n308 585
R154 B.n307 B.n80 585
R155 B.n306 B.n305 585
R156 B.n304 B.n81 585
R157 B.n303 B.n302 585
R158 B.n301 B.n82 585
R159 B.n300 B.n299 585
R160 B.n174 B.n173 585
R161 B.n175 B.n128 585
R162 B.n177 B.n176 585
R163 B.n178 B.n127 585
R164 B.n180 B.n179 585
R165 B.n181 B.n126 585
R166 B.n183 B.n182 585
R167 B.n184 B.n125 585
R168 B.n186 B.n185 585
R169 B.n187 B.n124 585
R170 B.n189 B.n188 585
R171 B.n190 B.n123 585
R172 B.n192 B.n191 585
R173 B.n193 B.n122 585
R174 B.n195 B.n194 585
R175 B.n196 B.n121 585
R176 B.n198 B.n197 585
R177 B.n199 B.n120 585
R178 B.n201 B.n200 585
R179 B.n202 B.n119 585
R180 B.n204 B.n203 585
R181 B.n205 B.n118 585
R182 B.n207 B.n206 585
R183 B.n208 B.n117 585
R184 B.n210 B.n209 585
R185 B.n211 B.n116 585
R186 B.n213 B.n212 585
R187 B.n214 B.n115 585
R188 B.n216 B.n215 585
R189 B.n217 B.n114 585
R190 B.n219 B.n218 585
R191 B.n220 B.n113 585
R192 B.n222 B.n221 585
R193 B.n223 B.n112 585
R194 B.n225 B.n224 585
R195 B.n226 B.n111 585
R196 B.n228 B.n227 585
R197 B.n230 B.n229 585
R198 B.n231 B.n107 585
R199 B.n233 B.n232 585
R200 B.n234 B.n106 585
R201 B.n236 B.n235 585
R202 B.n237 B.n105 585
R203 B.n239 B.n238 585
R204 B.n240 B.n104 585
R205 B.n242 B.n241 585
R206 B.n244 B.n101 585
R207 B.n246 B.n245 585
R208 B.n247 B.n100 585
R209 B.n249 B.n248 585
R210 B.n250 B.n99 585
R211 B.n252 B.n251 585
R212 B.n253 B.n98 585
R213 B.n255 B.n254 585
R214 B.n256 B.n97 585
R215 B.n258 B.n257 585
R216 B.n259 B.n96 585
R217 B.n261 B.n260 585
R218 B.n262 B.n95 585
R219 B.n264 B.n263 585
R220 B.n265 B.n94 585
R221 B.n267 B.n266 585
R222 B.n268 B.n93 585
R223 B.n270 B.n269 585
R224 B.n271 B.n92 585
R225 B.n273 B.n272 585
R226 B.n274 B.n91 585
R227 B.n276 B.n275 585
R228 B.n277 B.n90 585
R229 B.n279 B.n278 585
R230 B.n280 B.n89 585
R231 B.n282 B.n281 585
R232 B.n283 B.n88 585
R233 B.n285 B.n284 585
R234 B.n286 B.n87 585
R235 B.n288 B.n287 585
R236 B.n289 B.n86 585
R237 B.n291 B.n290 585
R238 B.n292 B.n85 585
R239 B.n294 B.n293 585
R240 B.n295 B.n84 585
R241 B.n297 B.n296 585
R242 B.n298 B.n83 585
R243 B.n172 B.n129 585
R244 B.n171 B.n170 585
R245 B.n169 B.n130 585
R246 B.n168 B.n167 585
R247 B.n166 B.n131 585
R248 B.n165 B.n164 585
R249 B.n163 B.n132 585
R250 B.n162 B.n161 585
R251 B.n160 B.n133 585
R252 B.n159 B.n158 585
R253 B.n157 B.n134 585
R254 B.n156 B.n155 585
R255 B.n154 B.n135 585
R256 B.n153 B.n152 585
R257 B.n151 B.n136 585
R258 B.n150 B.n149 585
R259 B.n148 B.n137 585
R260 B.n147 B.n146 585
R261 B.n145 B.n138 585
R262 B.n144 B.n143 585
R263 B.n142 B.n139 585
R264 B.n141 B.n140 585
R265 B.n2 B.n0 585
R266 B.n529 B.n1 585
R267 B.n528 B.n527 585
R268 B.n526 B.n3 585
R269 B.n525 B.n524 585
R270 B.n523 B.n4 585
R271 B.n522 B.n521 585
R272 B.n520 B.n5 585
R273 B.n519 B.n518 585
R274 B.n517 B.n6 585
R275 B.n516 B.n515 585
R276 B.n514 B.n7 585
R277 B.n513 B.n512 585
R278 B.n511 B.n8 585
R279 B.n510 B.n509 585
R280 B.n508 B.n9 585
R281 B.n507 B.n506 585
R282 B.n505 B.n10 585
R283 B.n504 B.n503 585
R284 B.n502 B.n11 585
R285 B.n501 B.n500 585
R286 B.n499 B.n12 585
R287 B.n498 B.n497 585
R288 B.n496 B.n13 585
R289 B.n531 B.n530 585
R290 B.n174 B.n129 545.355
R291 B.n494 B.n13 545.355
R292 B.n300 B.n83 545.355
R293 B.n368 B.n59 545.355
R294 B.n102 B.t9 387.695
R295 B.n108 B.t6 387.695
R296 B.n32 B.t3 387.695
R297 B.n40 B.t0 387.695
R298 B.n170 B.n129 163.367
R299 B.n170 B.n169 163.367
R300 B.n169 B.n168 163.367
R301 B.n168 B.n131 163.367
R302 B.n164 B.n131 163.367
R303 B.n164 B.n163 163.367
R304 B.n163 B.n162 163.367
R305 B.n162 B.n133 163.367
R306 B.n158 B.n133 163.367
R307 B.n158 B.n157 163.367
R308 B.n157 B.n156 163.367
R309 B.n156 B.n135 163.367
R310 B.n152 B.n135 163.367
R311 B.n152 B.n151 163.367
R312 B.n151 B.n150 163.367
R313 B.n150 B.n137 163.367
R314 B.n146 B.n137 163.367
R315 B.n146 B.n145 163.367
R316 B.n145 B.n144 163.367
R317 B.n144 B.n139 163.367
R318 B.n140 B.n139 163.367
R319 B.n140 B.n2 163.367
R320 B.n530 B.n2 163.367
R321 B.n530 B.n529 163.367
R322 B.n529 B.n528 163.367
R323 B.n528 B.n3 163.367
R324 B.n524 B.n3 163.367
R325 B.n524 B.n523 163.367
R326 B.n523 B.n522 163.367
R327 B.n522 B.n5 163.367
R328 B.n518 B.n5 163.367
R329 B.n518 B.n517 163.367
R330 B.n517 B.n516 163.367
R331 B.n516 B.n7 163.367
R332 B.n512 B.n7 163.367
R333 B.n512 B.n511 163.367
R334 B.n511 B.n510 163.367
R335 B.n510 B.n9 163.367
R336 B.n506 B.n9 163.367
R337 B.n506 B.n505 163.367
R338 B.n505 B.n504 163.367
R339 B.n504 B.n11 163.367
R340 B.n500 B.n11 163.367
R341 B.n500 B.n499 163.367
R342 B.n499 B.n498 163.367
R343 B.n498 B.n13 163.367
R344 B.n175 B.n174 163.367
R345 B.n176 B.n175 163.367
R346 B.n176 B.n127 163.367
R347 B.n180 B.n127 163.367
R348 B.n181 B.n180 163.367
R349 B.n182 B.n181 163.367
R350 B.n182 B.n125 163.367
R351 B.n186 B.n125 163.367
R352 B.n187 B.n186 163.367
R353 B.n188 B.n187 163.367
R354 B.n188 B.n123 163.367
R355 B.n192 B.n123 163.367
R356 B.n193 B.n192 163.367
R357 B.n194 B.n193 163.367
R358 B.n194 B.n121 163.367
R359 B.n198 B.n121 163.367
R360 B.n199 B.n198 163.367
R361 B.n200 B.n199 163.367
R362 B.n200 B.n119 163.367
R363 B.n204 B.n119 163.367
R364 B.n205 B.n204 163.367
R365 B.n206 B.n205 163.367
R366 B.n206 B.n117 163.367
R367 B.n210 B.n117 163.367
R368 B.n211 B.n210 163.367
R369 B.n212 B.n211 163.367
R370 B.n212 B.n115 163.367
R371 B.n216 B.n115 163.367
R372 B.n217 B.n216 163.367
R373 B.n218 B.n217 163.367
R374 B.n218 B.n113 163.367
R375 B.n222 B.n113 163.367
R376 B.n223 B.n222 163.367
R377 B.n224 B.n223 163.367
R378 B.n224 B.n111 163.367
R379 B.n228 B.n111 163.367
R380 B.n229 B.n228 163.367
R381 B.n229 B.n107 163.367
R382 B.n233 B.n107 163.367
R383 B.n234 B.n233 163.367
R384 B.n235 B.n234 163.367
R385 B.n235 B.n105 163.367
R386 B.n239 B.n105 163.367
R387 B.n240 B.n239 163.367
R388 B.n241 B.n240 163.367
R389 B.n241 B.n101 163.367
R390 B.n246 B.n101 163.367
R391 B.n247 B.n246 163.367
R392 B.n248 B.n247 163.367
R393 B.n248 B.n99 163.367
R394 B.n252 B.n99 163.367
R395 B.n253 B.n252 163.367
R396 B.n254 B.n253 163.367
R397 B.n254 B.n97 163.367
R398 B.n258 B.n97 163.367
R399 B.n259 B.n258 163.367
R400 B.n260 B.n259 163.367
R401 B.n260 B.n95 163.367
R402 B.n264 B.n95 163.367
R403 B.n265 B.n264 163.367
R404 B.n266 B.n265 163.367
R405 B.n266 B.n93 163.367
R406 B.n270 B.n93 163.367
R407 B.n271 B.n270 163.367
R408 B.n272 B.n271 163.367
R409 B.n272 B.n91 163.367
R410 B.n276 B.n91 163.367
R411 B.n277 B.n276 163.367
R412 B.n278 B.n277 163.367
R413 B.n278 B.n89 163.367
R414 B.n282 B.n89 163.367
R415 B.n283 B.n282 163.367
R416 B.n284 B.n283 163.367
R417 B.n284 B.n87 163.367
R418 B.n288 B.n87 163.367
R419 B.n289 B.n288 163.367
R420 B.n290 B.n289 163.367
R421 B.n290 B.n85 163.367
R422 B.n294 B.n85 163.367
R423 B.n295 B.n294 163.367
R424 B.n296 B.n295 163.367
R425 B.n296 B.n83 163.367
R426 B.n301 B.n300 163.367
R427 B.n302 B.n301 163.367
R428 B.n302 B.n81 163.367
R429 B.n306 B.n81 163.367
R430 B.n307 B.n306 163.367
R431 B.n308 B.n307 163.367
R432 B.n308 B.n79 163.367
R433 B.n312 B.n79 163.367
R434 B.n313 B.n312 163.367
R435 B.n314 B.n313 163.367
R436 B.n314 B.n77 163.367
R437 B.n318 B.n77 163.367
R438 B.n319 B.n318 163.367
R439 B.n320 B.n319 163.367
R440 B.n320 B.n75 163.367
R441 B.n324 B.n75 163.367
R442 B.n325 B.n324 163.367
R443 B.n326 B.n325 163.367
R444 B.n326 B.n73 163.367
R445 B.n330 B.n73 163.367
R446 B.n331 B.n330 163.367
R447 B.n332 B.n331 163.367
R448 B.n332 B.n71 163.367
R449 B.n336 B.n71 163.367
R450 B.n337 B.n336 163.367
R451 B.n338 B.n337 163.367
R452 B.n338 B.n69 163.367
R453 B.n342 B.n69 163.367
R454 B.n343 B.n342 163.367
R455 B.n344 B.n343 163.367
R456 B.n344 B.n67 163.367
R457 B.n348 B.n67 163.367
R458 B.n349 B.n348 163.367
R459 B.n350 B.n349 163.367
R460 B.n350 B.n65 163.367
R461 B.n354 B.n65 163.367
R462 B.n355 B.n354 163.367
R463 B.n356 B.n355 163.367
R464 B.n356 B.n63 163.367
R465 B.n360 B.n63 163.367
R466 B.n361 B.n360 163.367
R467 B.n362 B.n361 163.367
R468 B.n362 B.n61 163.367
R469 B.n366 B.n61 163.367
R470 B.n367 B.n366 163.367
R471 B.n368 B.n367 163.367
R472 B.n494 B.n493 163.367
R473 B.n493 B.n492 163.367
R474 B.n492 B.n15 163.367
R475 B.n488 B.n15 163.367
R476 B.n488 B.n487 163.367
R477 B.n487 B.n486 163.367
R478 B.n486 B.n17 163.367
R479 B.n482 B.n17 163.367
R480 B.n482 B.n481 163.367
R481 B.n481 B.n480 163.367
R482 B.n480 B.n19 163.367
R483 B.n476 B.n19 163.367
R484 B.n476 B.n475 163.367
R485 B.n475 B.n474 163.367
R486 B.n474 B.n21 163.367
R487 B.n470 B.n21 163.367
R488 B.n470 B.n469 163.367
R489 B.n469 B.n468 163.367
R490 B.n468 B.n23 163.367
R491 B.n464 B.n23 163.367
R492 B.n464 B.n463 163.367
R493 B.n463 B.n462 163.367
R494 B.n462 B.n25 163.367
R495 B.n458 B.n25 163.367
R496 B.n458 B.n457 163.367
R497 B.n457 B.n456 163.367
R498 B.n456 B.n27 163.367
R499 B.n452 B.n27 163.367
R500 B.n452 B.n451 163.367
R501 B.n451 B.n450 163.367
R502 B.n450 B.n29 163.367
R503 B.n446 B.n29 163.367
R504 B.n446 B.n445 163.367
R505 B.n445 B.n444 163.367
R506 B.n444 B.n31 163.367
R507 B.n440 B.n31 163.367
R508 B.n440 B.n439 163.367
R509 B.n439 B.n35 163.367
R510 B.n435 B.n35 163.367
R511 B.n435 B.n434 163.367
R512 B.n434 B.n433 163.367
R513 B.n433 B.n37 163.367
R514 B.n429 B.n37 163.367
R515 B.n429 B.n428 163.367
R516 B.n428 B.n427 163.367
R517 B.n427 B.n39 163.367
R518 B.n422 B.n39 163.367
R519 B.n422 B.n421 163.367
R520 B.n421 B.n420 163.367
R521 B.n420 B.n43 163.367
R522 B.n416 B.n43 163.367
R523 B.n416 B.n415 163.367
R524 B.n415 B.n414 163.367
R525 B.n414 B.n45 163.367
R526 B.n410 B.n45 163.367
R527 B.n410 B.n409 163.367
R528 B.n409 B.n408 163.367
R529 B.n408 B.n47 163.367
R530 B.n404 B.n47 163.367
R531 B.n404 B.n403 163.367
R532 B.n403 B.n402 163.367
R533 B.n402 B.n49 163.367
R534 B.n398 B.n49 163.367
R535 B.n398 B.n397 163.367
R536 B.n397 B.n396 163.367
R537 B.n396 B.n51 163.367
R538 B.n392 B.n51 163.367
R539 B.n392 B.n391 163.367
R540 B.n391 B.n390 163.367
R541 B.n390 B.n53 163.367
R542 B.n386 B.n53 163.367
R543 B.n386 B.n385 163.367
R544 B.n385 B.n384 163.367
R545 B.n384 B.n55 163.367
R546 B.n380 B.n55 163.367
R547 B.n380 B.n379 163.367
R548 B.n379 B.n378 163.367
R549 B.n378 B.n57 163.367
R550 B.n374 B.n57 163.367
R551 B.n374 B.n373 163.367
R552 B.n373 B.n372 163.367
R553 B.n372 B.n59 163.367
R554 B.n102 B.t11 144.2
R555 B.n40 B.t1 144.2
R556 B.n108 B.t8 144.188
R557 B.n32 B.t4 144.188
R558 B.n103 B.t10 111.23
R559 B.n41 B.t2 111.23
R560 B.n109 B.t7 111.218
R561 B.n33 B.t5 111.218
R562 B.n243 B.n103 59.5399
R563 B.n110 B.n109 59.5399
R564 B.n34 B.n33 59.5399
R565 B.n425 B.n41 59.5399
R566 B.n496 B.n495 35.4346
R567 B.n299 B.n298 35.4346
R568 B.n173 B.n172 35.4346
R569 B.n370 B.n369 35.4346
R570 B.n103 B.n102 32.9702
R571 B.n109 B.n108 32.9702
R572 B.n33 B.n32 32.9702
R573 B.n41 B.n40 32.9702
R574 B B.n531 18.0485
R575 B.n495 B.n14 10.6151
R576 B.n491 B.n14 10.6151
R577 B.n491 B.n490 10.6151
R578 B.n490 B.n489 10.6151
R579 B.n489 B.n16 10.6151
R580 B.n485 B.n16 10.6151
R581 B.n485 B.n484 10.6151
R582 B.n484 B.n483 10.6151
R583 B.n483 B.n18 10.6151
R584 B.n479 B.n18 10.6151
R585 B.n479 B.n478 10.6151
R586 B.n478 B.n477 10.6151
R587 B.n477 B.n20 10.6151
R588 B.n473 B.n20 10.6151
R589 B.n473 B.n472 10.6151
R590 B.n472 B.n471 10.6151
R591 B.n471 B.n22 10.6151
R592 B.n467 B.n22 10.6151
R593 B.n467 B.n466 10.6151
R594 B.n466 B.n465 10.6151
R595 B.n465 B.n24 10.6151
R596 B.n461 B.n24 10.6151
R597 B.n461 B.n460 10.6151
R598 B.n460 B.n459 10.6151
R599 B.n459 B.n26 10.6151
R600 B.n455 B.n26 10.6151
R601 B.n455 B.n454 10.6151
R602 B.n454 B.n453 10.6151
R603 B.n453 B.n28 10.6151
R604 B.n449 B.n28 10.6151
R605 B.n449 B.n448 10.6151
R606 B.n448 B.n447 10.6151
R607 B.n447 B.n30 10.6151
R608 B.n443 B.n30 10.6151
R609 B.n443 B.n442 10.6151
R610 B.n442 B.n441 10.6151
R611 B.n438 B.n437 10.6151
R612 B.n437 B.n436 10.6151
R613 B.n436 B.n36 10.6151
R614 B.n432 B.n36 10.6151
R615 B.n432 B.n431 10.6151
R616 B.n431 B.n430 10.6151
R617 B.n430 B.n38 10.6151
R618 B.n426 B.n38 10.6151
R619 B.n424 B.n423 10.6151
R620 B.n423 B.n42 10.6151
R621 B.n419 B.n42 10.6151
R622 B.n419 B.n418 10.6151
R623 B.n418 B.n417 10.6151
R624 B.n417 B.n44 10.6151
R625 B.n413 B.n44 10.6151
R626 B.n413 B.n412 10.6151
R627 B.n412 B.n411 10.6151
R628 B.n411 B.n46 10.6151
R629 B.n407 B.n46 10.6151
R630 B.n407 B.n406 10.6151
R631 B.n406 B.n405 10.6151
R632 B.n405 B.n48 10.6151
R633 B.n401 B.n48 10.6151
R634 B.n401 B.n400 10.6151
R635 B.n400 B.n399 10.6151
R636 B.n399 B.n50 10.6151
R637 B.n395 B.n50 10.6151
R638 B.n395 B.n394 10.6151
R639 B.n394 B.n393 10.6151
R640 B.n393 B.n52 10.6151
R641 B.n389 B.n52 10.6151
R642 B.n389 B.n388 10.6151
R643 B.n388 B.n387 10.6151
R644 B.n387 B.n54 10.6151
R645 B.n383 B.n54 10.6151
R646 B.n383 B.n382 10.6151
R647 B.n382 B.n381 10.6151
R648 B.n381 B.n56 10.6151
R649 B.n377 B.n56 10.6151
R650 B.n377 B.n376 10.6151
R651 B.n376 B.n375 10.6151
R652 B.n375 B.n58 10.6151
R653 B.n371 B.n58 10.6151
R654 B.n371 B.n370 10.6151
R655 B.n299 B.n82 10.6151
R656 B.n303 B.n82 10.6151
R657 B.n304 B.n303 10.6151
R658 B.n305 B.n304 10.6151
R659 B.n305 B.n80 10.6151
R660 B.n309 B.n80 10.6151
R661 B.n310 B.n309 10.6151
R662 B.n311 B.n310 10.6151
R663 B.n311 B.n78 10.6151
R664 B.n315 B.n78 10.6151
R665 B.n316 B.n315 10.6151
R666 B.n317 B.n316 10.6151
R667 B.n317 B.n76 10.6151
R668 B.n321 B.n76 10.6151
R669 B.n322 B.n321 10.6151
R670 B.n323 B.n322 10.6151
R671 B.n323 B.n74 10.6151
R672 B.n327 B.n74 10.6151
R673 B.n328 B.n327 10.6151
R674 B.n329 B.n328 10.6151
R675 B.n329 B.n72 10.6151
R676 B.n333 B.n72 10.6151
R677 B.n334 B.n333 10.6151
R678 B.n335 B.n334 10.6151
R679 B.n335 B.n70 10.6151
R680 B.n339 B.n70 10.6151
R681 B.n340 B.n339 10.6151
R682 B.n341 B.n340 10.6151
R683 B.n341 B.n68 10.6151
R684 B.n345 B.n68 10.6151
R685 B.n346 B.n345 10.6151
R686 B.n347 B.n346 10.6151
R687 B.n347 B.n66 10.6151
R688 B.n351 B.n66 10.6151
R689 B.n352 B.n351 10.6151
R690 B.n353 B.n352 10.6151
R691 B.n353 B.n64 10.6151
R692 B.n357 B.n64 10.6151
R693 B.n358 B.n357 10.6151
R694 B.n359 B.n358 10.6151
R695 B.n359 B.n62 10.6151
R696 B.n363 B.n62 10.6151
R697 B.n364 B.n363 10.6151
R698 B.n365 B.n364 10.6151
R699 B.n365 B.n60 10.6151
R700 B.n369 B.n60 10.6151
R701 B.n173 B.n128 10.6151
R702 B.n177 B.n128 10.6151
R703 B.n178 B.n177 10.6151
R704 B.n179 B.n178 10.6151
R705 B.n179 B.n126 10.6151
R706 B.n183 B.n126 10.6151
R707 B.n184 B.n183 10.6151
R708 B.n185 B.n184 10.6151
R709 B.n185 B.n124 10.6151
R710 B.n189 B.n124 10.6151
R711 B.n190 B.n189 10.6151
R712 B.n191 B.n190 10.6151
R713 B.n191 B.n122 10.6151
R714 B.n195 B.n122 10.6151
R715 B.n196 B.n195 10.6151
R716 B.n197 B.n196 10.6151
R717 B.n197 B.n120 10.6151
R718 B.n201 B.n120 10.6151
R719 B.n202 B.n201 10.6151
R720 B.n203 B.n202 10.6151
R721 B.n203 B.n118 10.6151
R722 B.n207 B.n118 10.6151
R723 B.n208 B.n207 10.6151
R724 B.n209 B.n208 10.6151
R725 B.n209 B.n116 10.6151
R726 B.n213 B.n116 10.6151
R727 B.n214 B.n213 10.6151
R728 B.n215 B.n214 10.6151
R729 B.n215 B.n114 10.6151
R730 B.n219 B.n114 10.6151
R731 B.n220 B.n219 10.6151
R732 B.n221 B.n220 10.6151
R733 B.n221 B.n112 10.6151
R734 B.n225 B.n112 10.6151
R735 B.n226 B.n225 10.6151
R736 B.n227 B.n226 10.6151
R737 B.n231 B.n230 10.6151
R738 B.n232 B.n231 10.6151
R739 B.n232 B.n106 10.6151
R740 B.n236 B.n106 10.6151
R741 B.n237 B.n236 10.6151
R742 B.n238 B.n237 10.6151
R743 B.n238 B.n104 10.6151
R744 B.n242 B.n104 10.6151
R745 B.n245 B.n244 10.6151
R746 B.n245 B.n100 10.6151
R747 B.n249 B.n100 10.6151
R748 B.n250 B.n249 10.6151
R749 B.n251 B.n250 10.6151
R750 B.n251 B.n98 10.6151
R751 B.n255 B.n98 10.6151
R752 B.n256 B.n255 10.6151
R753 B.n257 B.n256 10.6151
R754 B.n257 B.n96 10.6151
R755 B.n261 B.n96 10.6151
R756 B.n262 B.n261 10.6151
R757 B.n263 B.n262 10.6151
R758 B.n263 B.n94 10.6151
R759 B.n267 B.n94 10.6151
R760 B.n268 B.n267 10.6151
R761 B.n269 B.n268 10.6151
R762 B.n269 B.n92 10.6151
R763 B.n273 B.n92 10.6151
R764 B.n274 B.n273 10.6151
R765 B.n275 B.n274 10.6151
R766 B.n275 B.n90 10.6151
R767 B.n279 B.n90 10.6151
R768 B.n280 B.n279 10.6151
R769 B.n281 B.n280 10.6151
R770 B.n281 B.n88 10.6151
R771 B.n285 B.n88 10.6151
R772 B.n286 B.n285 10.6151
R773 B.n287 B.n286 10.6151
R774 B.n287 B.n86 10.6151
R775 B.n291 B.n86 10.6151
R776 B.n292 B.n291 10.6151
R777 B.n293 B.n292 10.6151
R778 B.n293 B.n84 10.6151
R779 B.n297 B.n84 10.6151
R780 B.n298 B.n297 10.6151
R781 B.n172 B.n171 10.6151
R782 B.n171 B.n130 10.6151
R783 B.n167 B.n130 10.6151
R784 B.n167 B.n166 10.6151
R785 B.n166 B.n165 10.6151
R786 B.n165 B.n132 10.6151
R787 B.n161 B.n132 10.6151
R788 B.n161 B.n160 10.6151
R789 B.n160 B.n159 10.6151
R790 B.n159 B.n134 10.6151
R791 B.n155 B.n134 10.6151
R792 B.n155 B.n154 10.6151
R793 B.n154 B.n153 10.6151
R794 B.n153 B.n136 10.6151
R795 B.n149 B.n136 10.6151
R796 B.n149 B.n148 10.6151
R797 B.n148 B.n147 10.6151
R798 B.n147 B.n138 10.6151
R799 B.n143 B.n138 10.6151
R800 B.n143 B.n142 10.6151
R801 B.n142 B.n141 10.6151
R802 B.n141 B.n0 10.6151
R803 B.n527 B.n1 10.6151
R804 B.n527 B.n526 10.6151
R805 B.n526 B.n525 10.6151
R806 B.n525 B.n4 10.6151
R807 B.n521 B.n4 10.6151
R808 B.n521 B.n520 10.6151
R809 B.n520 B.n519 10.6151
R810 B.n519 B.n6 10.6151
R811 B.n515 B.n6 10.6151
R812 B.n515 B.n514 10.6151
R813 B.n514 B.n513 10.6151
R814 B.n513 B.n8 10.6151
R815 B.n509 B.n8 10.6151
R816 B.n509 B.n508 10.6151
R817 B.n508 B.n507 10.6151
R818 B.n507 B.n10 10.6151
R819 B.n503 B.n10 10.6151
R820 B.n503 B.n502 10.6151
R821 B.n502 B.n501 10.6151
R822 B.n501 B.n12 10.6151
R823 B.n497 B.n12 10.6151
R824 B.n497 B.n496 10.6151
R825 B.n438 B.n34 6.5566
R826 B.n426 B.n425 6.5566
R827 B.n230 B.n110 6.5566
R828 B.n243 B.n242 6.5566
R829 B.n441 B.n34 4.05904
R830 B.n425 B.n424 4.05904
R831 B.n227 B.n110 4.05904
R832 B.n244 B.n243 4.05904
R833 B.n531 B.n0 2.81026
R834 B.n531 B.n1 2.81026
R835 VP.n2 VP.t2 221.192
R836 VP.n2 VP.t3 220.96
R837 VP.n3 VP.t0 182.774
R838 VP.n9 VP.t1 182.774
R839 VP.n4 VP.n3 168.641
R840 VP.n10 VP.n9 168.641
R841 VP.n8 VP.n0 161.3
R842 VP.n7 VP.n6 161.3
R843 VP.n5 VP.n1 161.3
R844 VP.n4 VP.n2 58.9364
R845 VP.n7 VP.n1 40.4934
R846 VP.n8 VP.n7 40.4934
R847 VP.n3 VP.n1 17.1274
R848 VP.n9 VP.n8 17.1274
R849 VP.n5 VP.n4 0.189894
R850 VP.n6 VP.n5 0.189894
R851 VP.n6 VP.n0 0.189894
R852 VP.n10 VP.n0 0.189894
R853 VP VP.n10 0.0516364
R854 VDD1 VDD1.n1 115.419
R855 VDD1 VDD1.n0 77.8843
R856 VDD1.n0 VDD1.t1 3.12899
R857 VDD1.n0 VDD1.t0 3.12899
R858 VDD1.n1 VDD1.t3 3.12899
R859 VDD1.n1 VDD1.t2 3.12899
C0 VDD1 VP 3.73983f
C1 VDD2 w_n1990_n3046# 1.19137f
C2 VTAIL w_n1990_n3046# 3.64663f
C3 w_n1990_n3046# VN 3.10764f
C4 VDD2 VTAIL 5.15796f
C5 VDD2 VN 3.57211f
C6 B w_n1990_n3046# 7.28078f
C7 w_n1990_n3046# VP 3.36035f
C8 VDD2 B 1.03371f
C9 VTAIL VN 3.35394f
C10 VDD2 VP 0.315854f
C11 VTAIL B 3.81608f
C12 B VN 0.856233f
C13 VTAIL VP 3.36804f
C14 VDD1 w_n1990_n3046# 1.16262f
C15 VP VN 5.00339f
C16 VDD2 VDD1 0.725731f
C17 B VP 1.26987f
C18 VDD1 VTAIL 5.112f
C19 VDD1 VN 0.147704f
C20 VDD1 B 1.00162f
C21 VDD2 VSUBS 0.724533f
C22 VDD1 VSUBS 4.845682f
C23 VTAIL VSUBS 0.931206f
C24 VN VSUBS 5.14776f
C25 VP VSUBS 1.575664f
C26 B VSUBS 3.077732f
C27 w_n1990_n3046# VSUBS 74.816f
C28 VDD1.t1 VSUBS 0.219703f
C29 VDD1.t0 VSUBS 0.219703f
C30 VDD1.n0 VSUBS 1.67556f
C31 VDD1.t3 VSUBS 0.219703f
C32 VDD1.t2 VSUBS 0.219703f
C33 VDD1.n1 VSUBS 2.26103f
C34 VP.n0 VSUBS 0.048613f
C35 VP.t1 VSUBS 1.87702f
C36 VP.n1 VSUBS 0.083199f
C37 VP.t2 VSUBS 2.02826f
C38 VP.t3 VSUBS 2.02732f
C39 VP.n2 VSUBS 3.02476f
C40 VP.t0 VSUBS 1.87702f
C41 VP.n3 VSUBS 0.796625f
C42 VP.n4 VSUBS 2.65035f
C43 VP.n5 VSUBS 0.048613f
C44 VP.n6 VSUBS 0.048613f
C45 VP.n7 VSUBS 0.039299f
C46 VP.n8 VSUBS 0.083199f
C47 VP.n9 VSUBS 0.796625f
C48 VP.n10 VSUBS 0.042473f
C49 B.n0 VSUBS 0.004932f
C50 B.n1 VSUBS 0.004932f
C51 B.n2 VSUBS 0.0078f
C52 B.n3 VSUBS 0.0078f
C53 B.n4 VSUBS 0.0078f
C54 B.n5 VSUBS 0.0078f
C55 B.n6 VSUBS 0.0078f
C56 B.n7 VSUBS 0.0078f
C57 B.n8 VSUBS 0.0078f
C58 B.n9 VSUBS 0.0078f
C59 B.n10 VSUBS 0.0078f
C60 B.n11 VSUBS 0.0078f
C61 B.n12 VSUBS 0.0078f
C62 B.n13 VSUBS 0.018907f
C63 B.n14 VSUBS 0.0078f
C64 B.n15 VSUBS 0.0078f
C65 B.n16 VSUBS 0.0078f
C66 B.n17 VSUBS 0.0078f
C67 B.n18 VSUBS 0.0078f
C68 B.n19 VSUBS 0.0078f
C69 B.n20 VSUBS 0.0078f
C70 B.n21 VSUBS 0.0078f
C71 B.n22 VSUBS 0.0078f
C72 B.n23 VSUBS 0.0078f
C73 B.n24 VSUBS 0.0078f
C74 B.n25 VSUBS 0.0078f
C75 B.n26 VSUBS 0.0078f
C76 B.n27 VSUBS 0.0078f
C77 B.n28 VSUBS 0.0078f
C78 B.n29 VSUBS 0.0078f
C79 B.n30 VSUBS 0.0078f
C80 B.n31 VSUBS 0.0078f
C81 B.t5 VSUBS 0.371023f
C82 B.t4 VSUBS 0.38544f
C83 B.t3 VSUBS 0.695769f
C84 B.n32 VSUBS 0.171087f
C85 B.n33 VSUBS 0.074175f
C86 B.n34 VSUBS 0.018071f
C87 B.n35 VSUBS 0.0078f
C88 B.n36 VSUBS 0.0078f
C89 B.n37 VSUBS 0.0078f
C90 B.n38 VSUBS 0.0078f
C91 B.n39 VSUBS 0.0078f
C92 B.t2 VSUBS 0.371018f
C93 B.t1 VSUBS 0.385435f
C94 B.t0 VSUBS 0.695769f
C95 B.n40 VSUBS 0.171092f
C96 B.n41 VSUBS 0.07418f
C97 B.n42 VSUBS 0.0078f
C98 B.n43 VSUBS 0.0078f
C99 B.n44 VSUBS 0.0078f
C100 B.n45 VSUBS 0.0078f
C101 B.n46 VSUBS 0.0078f
C102 B.n47 VSUBS 0.0078f
C103 B.n48 VSUBS 0.0078f
C104 B.n49 VSUBS 0.0078f
C105 B.n50 VSUBS 0.0078f
C106 B.n51 VSUBS 0.0078f
C107 B.n52 VSUBS 0.0078f
C108 B.n53 VSUBS 0.0078f
C109 B.n54 VSUBS 0.0078f
C110 B.n55 VSUBS 0.0078f
C111 B.n56 VSUBS 0.0078f
C112 B.n57 VSUBS 0.0078f
C113 B.n58 VSUBS 0.0078f
C114 B.n59 VSUBS 0.019632f
C115 B.n60 VSUBS 0.0078f
C116 B.n61 VSUBS 0.0078f
C117 B.n62 VSUBS 0.0078f
C118 B.n63 VSUBS 0.0078f
C119 B.n64 VSUBS 0.0078f
C120 B.n65 VSUBS 0.0078f
C121 B.n66 VSUBS 0.0078f
C122 B.n67 VSUBS 0.0078f
C123 B.n68 VSUBS 0.0078f
C124 B.n69 VSUBS 0.0078f
C125 B.n70 VSUBS 0.0078f
C126 B.n71 VSUBS 0.0078f
C127 B.n72 VSUBS 0.0078f
C128 B.n73 VSUBS 0.0078f
C129 B.n74 VSUBS 0.0078f
C130 B.n75 VSUBS 0.0078f
C131 B.n76 VSUBS 0.0078f
C132 B.n77 VSUBS 0.0078f
C133 B.n78 VSUBS 0.0078f
C134 B.n79 VSUBS 0.0078f
C135 B.n80 VSUBS 0.0078f
C136 B.n81 VSUBS 0.0078f
C137 B.n82 VSUBS 0.0078f
C138 B.n83 VSUBS 0.019632f
C139 B.n84 VSUBS 0.0078f
C140 B.n85 VSUBS 0.0078f
C141 B.n86 VSUBS 0.0078f
C142 B.n87 VSUBS 0.0078f
C143 B.n88 VSUBS 0.0078f
C144 B.n89 VSUBS 0.0078f
C145 B.n90 VSUBS 0.0078f
C146 B.n91 VSUBS 0.0078f
C147 B.n92 VSUBS 0.0078f
C148 B.n93 VSUBS 0.0078f
C149 B.n94 VSUBS 0.0078f
C150 B.n95 VSUBS 0.0078f
C151 B.n96 VSUBS 0.0078f
C152 B.n97 VSUBS 0.0078f
C153 B.n98 VSUBS 0.0078f
C154 B.n99 VSUBS 0.0078f
C155 B.n100 VSUBS 0.0078f
C156 B.n101 VSUBS 0.0078f
C157 B.t10 VSUBS 0.371018f
C158 B.t11 VSUBS 0.385435f
C159 B.t9 VSUBS 0.695769f
C160 B.n102 VSUBS 0.171092f
C161 B.n103 VSUBS 0.07418f
C162 B.n104 VSUBS 0.0078f
C163 B.n105 VSUBS 0.0078f
C164 B.n106 VSUBS 0.0078f
C165 B.n107 VSUBS 0.0078f
C166 B.t7 VSUBS 0.371023f
C167 B.t8 VSUBS 0.38544f
C168 B.t6 VSUBS 0.695769f
C169 B.n108 VSUBS 0.171087f
C170 B.n109 VSUBS 0.074175f
C171 B.n110 VSUBS 0.018071f
C172 B.n111 VSUBS 0.0078f
C173 B.n112 VSUBS 0.0078f
C174 B.n113 VSUBS 0.0078f
C175 B.n114 VSUBS 0.0078f
C176 B.n115 VSUBS 0.0078f
C177 B.n116 VSUBS 0.0078f
C178 B.n117 VSUBS 0.0078f
C179 B.n118 VSUBS 0.0078f
C180 B.n119 VSUBS 0.0078f
C181 B.n120 VSUBS 0.0078f
C182 B.n121 VSUBS 0.0078f
C183 B.n122 VSUBS 0.0078f
C184 B.n123 VSUBS 0.0078f
C185 B.n124 VSUBS 0.0078f
C186 B.n125 VSUBS 0.0078f
C187 B.n126 VSUBS 0.0078f
C188 B.n127 VSUBS 0.0078f
C189 B.n128 VSUBS 0.0078f
C190 B.n129 VSUBS 0.018907f
C191 B.n130 VSUBS 0.0078f
C192 B.n131 VSUBS 0.0078f
C193 B.n132 VSUBS 0.0078f
C194 B.n133 VSUBS 0.0078f
C195 B.n134 VSUBS 0.0078f
C196 B.n135 VSUBS 0.0078f
C197 B.n136 VSUBS 0.0078f
C198 B.n137 VSUBS 0.0078f
C199 B.n138 VSUBS 0.0078f
C200 B.n139 VSUBS 0.0078f
C201 B.n140 VSUBS 0.0078f
C202 B.n141 VSUBS 0.0078f
C203 B.n142 VSUBS 0.0078f
C204 B.n143 VSUBS 0.0078f
C205 B.n144 VSUBS 0.0078f
C206 B.n145 VSUBS 0.0078f
C207 B.n146 VSUBS 0.0078f
C208 B.n147 VSUBS 0.0078f
C209 B.n148 VSUBS 0.0078f
C210 B.n149 VSUBS 0.0078f
C211 B.n150 VSUBS 0.0078f
C212 B.n151 VSUBS 0.0078f
C213 B.n152 VSUBS 0.0078f
C214 B.n153 VSUBS 0.0078f
C215 B.n154 VSUBS 0.0078f
C216 B.n155 VSUBS 0.0078f
C217 B.n156 VSUBS 0.0078f
C218 B.n157 VSUBS 0.0078f
C219 B.n158 VSUBS 0.0078f
C220 B.n159 VSUBS 0.0078f
C221 B.n160 VSUBS 0.0078f
C222 B.n161 VSUBS 0.0078f
C223 B.n162 VSUBS 0.0078f
C224 B.n163 VSUBS 0.0078f
C225 B.n164 VSUBS 0.0078f
C226 B.n165 VSUBS 0.0078f
C227 B.n166 VSUBS 0.0078f
C228 B.n167 VSUBS 0.0078f
C229 B.n168 VSUBS 0.0078f
C230 B.n169 VSUBS 0.0078f
C231 B.n170 VSUBS 0.0078f
C232 B.n171 VSUBS 0.0078f
C233 B.n172 VSUBS 0.018907f
C234 B.n173 VSUBS 0.019632f
C235 B.n174 VSUBS 0.019632f
C236 B.n175 VSUBS 0.0078f
C237 B.n176 VSUBS 0.0078f
C238 B.n177 VSUBS 0.0078f
C239 B.n178 VSUBS 0.0078f
C240 B.n179 VSUBS 0.0078f
C241 B.n180 VSUBS 0.0078f
C242 B.n181 VSUBS 0.0078f
C243 B.n182 VSUBS 0.0078f
C244 B.n183 VSUBS 0.0078f
C245 B.n184 VSUBS 0.0078f
C246 B.n185 VSUBS 0.0078f
C247 B.n186 VSUBS 0.0078f
C248 B.n187 VSUBS 0.0078f
C249 B.n188 VSUBS 0.0078f
C250 B.n189 VSUBS 0.0078f
C251 B.n190 VSUBS 0.0078f
C252 B.n191 VSUBS 0.0078f
C253 B.n192 VSUBS 0.0078f
C254 B.n193 VSUBS 0.0078f
C255 B.n194 VSUBS 0.0078f
C256 B.n195 VSUBS 0.0078f
C257 B.n196 VSUBS 0.0078f
C258 B.n197 VSUBS 0.0078f
C259 B.n198 VSUBS 0.0078f
C260 B.n199 VSUBS 0.0078f
C261 B.n200 VSUBS 0.0078f
C262 B.n201 VSUBS 0.0078f
C263 B.n202 VSUBS 0.0078f
C264 B.n203 VSUBS 0.0078f
C265 B.n204 VSUBS 0.0078f
C266 B.n205 VSUBS 0.0078f
C267 B.n206 VSUBS 0.0078f
C268 B.n207 VSUBS 0.0078f
C269 B.n208 VSUBS 0.0078f
C270 B.n209 VSUBS 0.0078f
C271 B.n210 VSUBS 0.0078f
C272 B.n211 VSUBS 0.0078f
C273 B.n212 VSUBS 0.0078f
C274 B.n213 VSUBS 0.0078f
C275 B.n214 VSUBS 0.0078f
C276 B.n215 VSUBS 0.0078f
C277 B.n216 VSUBS 0.0078f
C278 B.n217 VSUBS 0.0078f
C279 B.n218 VSUBS 0.0078f
C280 B.n219 VSUBS 0.0078f
C281 B.n220 VSUBS 0.0078f
C282 B.n221 VSUBS 0.0078f
C283 B.n222 VSUBS 0.0078f
C284 B.n223 VSUBS 0.0078f
C285 B.n224 VSUBS 0.0078f
C286 B.n225 VSUBS 0.0078f
C287 B.n226 VSUBS 0.0078f
C288 B.n227 VSUBS 0.005391f
C289 B.n228 VSUBS 0.0078f
C290 B.n229 VSUBS 0.0078f
C291 B.n230 VSUBS 0.006309f
C292 B.n231 VSUBS 0.0078f
C293 B.n232 VSUBS 0.0078f
C294 B.n233 VSUBS 0.0078f
C295 B.n234 VSUBS 0.0078f
C296 B.n235 VSUBS 0.0078f
C297 B.n236 VSUBS 0.0078f
C298 B.n237 VSUBS 0.0078f
C299 B.n238 VSUBS 0.0078f
C300 B.n239 VSUBS 0.0078f
C301 B.n240 VSUBS 0.0078f
C302 B.n241 VSUBS 0.0078f
C303 B.n242 VSUBS 0.006309f
C304 B.n243 VSUBS 0.018071f
C305 B.n244 VSUBS 0.005391f
C306 B.n245 VSUBS 0.0078f
C307 B.n246 VSUBS 0.0078f
C308 B.n247 VSUBS 0.0078f
C309 B.n248 VSUBS 0.0078f
C310 B.n249 VSUBS 0.0078f
C311 B.n250 VSUBS 0.0078f
C312 B.n251 VSUBS 0.0078f
C313 B.n252 VSUBS 0.0078f
C314 B.n253 VSUBS 0.0078f
C315 B.n254 VSUBS 0.0078f
C316 B.n255 VSUBS 0.0078f
C317 B.n256 VSUBS 0.0078f
C318 B.n257 VSUBS 0.0078f
C319 B.n258 VSUBS 0.0078f
C320 B.n259 VSUBS 0.0078f
C321 B.n260 VSUBS 0.0078f
C322 B.n261 VSUBS 0.0078f
C323 B.n262 VSUBS 0.0078f
C324 B.n263 VSUBS 0.0078f
C325 B.n264 VSUBS 0.0078f
C326 B.n265 VSUBS 0.0078f
C327 B.n266 VSUBS 0.0078f
C328 B.n267 VSUBS 0.0078f
C329 B.n268 VSUBS 0.0078f
C330 B.n269 VSUBS 0.0078f
C331 B.n270 VSUBS 0.0078f
C332 B.n271 VSUBS 0.0078f
C333 B.n272 VSUBS 0.0078f
C334 B.n273 VSUBS 0.0078f
C335 B.n274 VSUBS 0.0078f
C336 B.n275 VSUBS 0.0078f
C337 B.n276 VSUBS 0.0078f
C338 B.n277 VSUBS 0.0078f
C339 B.n278 VSUBS 0.0078f
C340 B.n279 VSUBS 0.0078f
C341 B.n280 VSUBS 0.0078f
C342 B.n281 VSUBS 0.0078f
C343 B.n282 VSUBS 0.0078f
C344 B.n283 VSUBS 0.0078f
C345 B.n284 VSUBS 0.0078f
C346 B.n285 VSUBS 0.0078f
C347 B.n286 VSUBS 0.0078f
C348 B.n287 VSUBS 0.0078f
C349 B.n288 VSUBS 0.0078f
C350 B.n289 VSUBS 0.0078f
C351 B.n290 VSUBS 0.0078f
C352 B.n291 VSUBS 0.0078f
C353 B.n292 VSUBS 0.0078f
C354 B.n293 VSUBS 0.0078f
C355 B.n294 VSUBS 0.0078f
C356 B.n295 VSUBS 0.0078f
C357 B.n296 VSUBS 0.0078f
C358 B.n297 VSUBS 0.0078f
C359 B.n298 VSUBS 0.019632f
C360 B.n299 VSUBS 0.018907f
C361 B.n300 VSUBS 0.018907f
C362 B.n301 VSUBS 0.0078f
C363 B.n302 VSUBS 0.0078f
C364 B.n303 VSUBS 0.0078f
C365 B.n304 VSUBS 0.0078f
C366 B.n305 VSUBS 0.0078f
C367 B.n306 VSUBS 0.0078f
C368 B.n307 VSUBS 0.0078f
C369 B.n308 VSUBS 0.0078f
C370 B.n309 VSUBS 0.0078f
C371 B.n310 VSUBS 0.0078f
C372 B.n311 VSUBS 0.0078f
C373 B.n312 VSUBS 0.0078f
C374 B.n313 VSUBS 0.0078f
C375 B.n314 VSUBS 0.0078f
C376 B.n315 VSUBS 0.0078f
C377 B.n316 VSUBS 0.0078f
C378 B.n317 VSUBS 0.0078f
C379 B.n318 VSUBS 0.0078f
C380 B.n319 VSUBS 0.0078f
C381 B.n320 VSUBS 0.0078f
C382 B.n321 VSUBS 0.0078f
C383 B.n322 VSUBS 0.0078f
C384 B.n323 VSUBS 0.0078f
C385 B.n324 VSUBS 0.0078f
C386 B.n325 VSUBS 0.0078f
C387 B.n326 VSUBS 0.0078f
C388 B.n327 VSUBS 0.0078f
C389 B.n328 VSUBS 0.0078f
C390 B.n329 VSUBS 0.0078f
C391 B.n330 VSUBS 0.0078f
C392 B.n331 VSUBS 0.0078f
C393 B.n332 VSUBS 0.0078f
C394 B.n333 VSUBS 0.0078f
C395 B.n334 VSUBS 0.0078f
C396 B.n335 VSUBS 0.0078f
C397 B.n336 VSUBS 0.0078f
C398 B.n337 VSUBS 0.0078f
C399 B.n338 VSUBS 0.0078f
C400 B.n339 VSUBS 0.0078f
C401 B.n340 VSUBS 0.0078f
C402 B.n341 VSUBS 0.0078f
C403 B.n342 VSUBS 0.0078f
C404 B.n343 VSUBS 0.0078f
C405 B.n344 VSUBS 0.0078f
C406 B.n345 VSUBS 0.0078f
C407 B.n346 VSUBS 0.0078f
C408 B.n347 VSUBS 0.0078f
C409 B.n348 VSUBS 0.0078f
C410 B.n349 VSUBS 0.0078f
C411 B.n350 VSUBS 0.0078f
C412 B.n351 VSUBS 0.0078f
C413 B.n352 VSUBS 0.0078f
C414 B.n353 VSUBS 0.0078f
C415 B.n354 VSUBS 0.0078f
C416 B.n355 VSUBS 0.0078f
C417 B.n356 VSUBS 0.0078f
C418 B.n357 VSUBS 0.0078f
C419 B.n358 VSUBS 0.0078f
C420 B.n359 VSUBS 0.0078f
C421 B.n360 VSUBS 0.0078f
C422 B.n361 VSUBS 0.0078f
C423 B.n362 VSUBS 0.0078f
C424 B.n363 VSUBS 0.0078f
C425 B.n364 VSUBS 0.0078f
C426 B.n365 VSUBS 0.0078f
C427 B.n366 VSUBS 0.0078f
C428 B.n367 VSUBS 0.0078f
C429 B.n368 VSUBS 0.018907f
C430 B.n369 VSUBS 0.019757f
C431 B.n370 VSUBS 0.018783f
C432 B.n371 VSUBS 0.0078f
C433 B.n372 VSUBS 0.0078f
C434 B.n373 VSUBS 0.0078f
C435 B.n374 VSUBS 0.0078f
C436 B.n375 VSUBS 0.0078f
C437 B.n376 VSUBS 0.0078f
C438 B.n377 VSUBS 0.0078f
C439 B.n378 VSUBS 0.0078f
C440 B.n379 VSUBS 0.0078f
C441 B.n380 VSUBS 0.0078f
C442 B.n381 VSUBS 0.0078f
C443 B.n382 VSUBS 0.0078f
C444 B.n383 VSUBS 0.0078f
C445 B.n384 VSUBS 0.0078f
C446 B.n385 VSUBS 0.0078f
C447 B.n386 VSUBS 0.0078f
C448 B.n387 VSUBS 0.0078f
C449 B.n388 VSUBS 0.0078f
C450 B.n389 VSUBS 0.0078f
C451 B.n390 VSUBS 0.0078f
C452 B.n391 VSUBS 0.0078f
C453 B.n392 VSUBS 0.0078f
C454 B.n393 VSUBS 0.0078f
C455 B.n394 VSUBS 0.0078f
C456 B.n395 VSUBS 0.0078f
C457 B.n396 VSUBS 0.0078f
C458 B.n397 VSUBS 0.0078f
C459 B.n398 VSUBS 0.0078f
C460 B.n399 VSUBS 0.0078f
C461 B.n400 VSUBS 0.0078f
C462 B.n401 VSUBS 0.0078f
C463 B.n402 VSUBS 0.0078f
C464 B.n403 VSUBS 0.0078f
C465 B.n404 VSUBS 0.0078f
C466 B.n405 VSUBS 0.0078f
C467 B.n406 VSUBS 0.0078f
C468 B.n407 VSUBS 0.0078f
C469 B.n408 VSUBS 0.0078f
C470 B.n409 VSUBS 0.0078f
C471 B.n410 VSUBS 0.0078f
C472 B.n411 VSUBS 0.0078f
C473 B.n412 VSUBS 0.0078f
C474 B.n413 VSUBS 0.0078f
C475 B.n414 VSUBS 0.0078f
C476 B.n415 VSUBS 0.0078f
C477 B.n416 VSUBS 0.0078f
C478 B.n417 VSUBS 0.0078f
C479 B.n418 VSUBS 0.0078f
C480 B.n419 VSUBS 0.0078f
C481 B.n420 VSUBS 0.0078f
C482 B.n421 VSUBS 0.0078f
C483 B.n422 VSUBS 0.0078f
C484 B.n423 VSUBS 0.0078f
C485 B.n424 VSUBS 0.005391f
C486 B.n425 VSUBS 0.018071f
C487 B.n426 VSUBS 0.006309f
C488 B.n427 VSUBS 0.0078f
C489 B.n428 VSUBS 0.0078f
C490 B.n429 VSUBS 0.0078f
C491 B.n430 VSUBS 0.0078f
C492 B.n431 VSUBS 0.0078f
C493 B.n432 VSUBS 0.0078f
C494 B.n433 VSUBS 0.0078f
C495 B.n434 VSUBS 0.0078f
C496 B.n435 VSUBS 0.0078f
C497 B.n436 VSUBS 0.0078f
C498 B.n437 VSUBS 0.0078f
C499 B.n438 VSUBS 0.006309f
C500 B.n439 VSUBS 0.0078f
C501 B.n440 VSUBS 0.0078f
C502 B.n441 VSUBS 0.005391f
C503 B.n442 VSUBS 0.0078f
C504 B.n443 VSUBS 0.0078f
C505 B.n444 VSUBS 0.0078f
C506 B.n445 VSUBS 0.0078f
C507 B.n446 VSUBS 0.0078f
C508 B.n447 VSUBS 0.0078f
C509 B.n448 VSUBS 0.0078f
C510 B.n449 VSUBS 0.0078f
C511 B.n450 VSUBS 0.0078f
C512 B.n451 VSUBS 0.0078f
C513 B.n452 VSUBS 0.0078f
C514 B.n453 VSUBS 0.0078f
C515 B.n454 VSUBS 0.0078f
C516 B.n455 VSUBS 0.0078f
C517 B.n456 VSUBS 0.0078f
C518 B.n457 VSUBS 0.0078f
C519 B.n458 VSUBS 0.0078f
C520 B.n459 VSUBS 0.0078f
C521 B.n460 VSUBS 0.0078f
C522 B.n461 VSUBS 0.0078f
C523 B.n462 VSUBS 0.0078f
C524 B.n463 VSUBS 0.0078f
C525 B.n464 VSUBS 0.0078f
C526 B.n465 VSUBS 0.0078f
C527 B.n466 VSUBS 0.0078f
C528 B.n467 VSUBS 0.0078f
C529 B.n468 VSUBS 0.0078f
C530 B.n469 VSUBS 0.0078f
C531 B.n470 VSUBS 0.0078f
C532 B.n471 VSUBS 0.0078f
C533 B.n472 VSUBS 0.0078f
C534 B.n473 VSUBS 0.0078f
C535 B.n474 VSUBS 0.0078f
C536 B.n475 VSUBS 0.0078f
C537 B.n476 VSUBS 0.0078f
C538 B.n477 VSUBS 0.0078f
C539 B.n478 VSUBS 0.0078f
C540 B.n479 VSUBS 0.0078f
C541 B.n480 VSUBS 0.0078f
C542 B.n481 VSUBS 0.0078f
C543 B.n482 VSUBS 0.0078f
C544 B.n483 VSUBS 0.0078f
C545 B.n484 VSUBS 0.0078f
C546 B.n485 VSUBS 0.0078f
C547 B.n486 VSUBS 0.0078f
C548 B.n487 VSUBS 0.0078f
C549 B.n488 VSUBS 0.0078f
C550 B.n489 VSUBS 0.0078f
C551 B.n490 VSUBS 0.0078f
C552 B.n491 VSUBS 0.0078f
C553 B.n492 VSUBS 0.0078f
C554 B.n493 VSUBS 0.0078f
C555 B.n494 VSUBS 0.019632f
C556 B.n495 VSUBS 0.019632f
C557 B.n496 VSUBS 0.018907f
C558 B.n497 VSUBS 0.0078f
C559 B.n498 VSUBS 0.0078f
C560 B.n499 VSUBS 0.0078f
C561 B.n500 VSUBS 0.0078f
C562 B.n501 VSUBS 0.0078f
C563 B.n502 VSUBS 0.0078f
C564 B.n503 VSUBS 0.0078f
C565 B.n504 VSUBS 0.0078f
C566 B.n505 VSUBS 0.0078f
C567 B.n506 VSUBS 0.0078f
C568 B.n507 VSUBS 0.0078f
C569 B.n508 VSUBS 0.0078f
C570 B.n509 VSUBS 0.0078f
C571 B.n510 VSUBS 0.0078f
C572 B.n511 VSUBS 0.0078f
C573 B.n512 VSUBS 0.0078f
C574 B.n513 VSUBS 0.0078f
C575 B.n514 VSUBS 0.0078f
C576 B.n515 VSUBS 0.0078f
C577 B.n516 VSUBS 0.0078f
C578 B.n517 VSUBS 0.0078f
C579 B.n518 VSUBS 0.0078f
C580 B.n519 VSUBS 0.0078f
C581 B.n520 VSUBS 0.0078f
C582 B.n521 VSUBS 0.0078f
C583 B.n522 VSUBS 0.0078f
C584 B.n523 VSUBS 0.0078f
C585 B.n524 VSUBS 0.0078f
C586 B.n525 VSUBS 0.0078f
C587 B.n526 VSUBS 0.0078f
C588 B.n527 VSUBS 0.0078f
C589 B.n528 VSUBS 0.0078f
C590 B.n529 VSUBS 0.0078f
C591 B.n530 VSUBS 0.0078f
C592 B.n531 VSUBS 0.017661f
C593 VTAIL.t7 VSUBS 1.79433f
C594 VTAIL.n0 VSUBS 0.682666f
C595 VTAIL.t2 VSUBS 1.79433f
C596 VTAIL.n1 VSUBS 0.733572f
C597 VTAIL.t3 VSUBS 1.79433f
C598 VTAIL.n2 VSUBS 1.80277f
C599 VTAIL.t5 VSUBS 1.79433f
C600 VTAIL.n3 VSUBS 1.80277f
C601 VTAIL.t6 VSUBS 1.79433f
C602 VTAIL.n4 VSUBS 0.733567f
C603 VTAIL.t1 VSUBS 1.79433f
C604 VTAIL.n5 VSUBS 0.733567f
C605 VTAIL.t0 VSUBS 1.79433f
C606 VTAIL.n6 VSUBS 1.80277f
C607 VTAIL.t4 VSUBS 1.79433f
C608 VTAIL.n7 VSUBS 1.74308f
C609 VDD2.t0 VSUBS 0.222199f
C610 VDD2.t1 VSUBS 0.222199f
C611 VDD2.n0 VSUBS 2.26346f
C612 VDD2.t2 VSUBS 0.222199f
C613 VDD2.t3 VSUBS 0.222199f
C614 VDD2.n1 VSUBS 1.69412f
C615 VDD2.n2 VSUBS 3.82f
C616 VN.t0 VSUBS 1.96724f
C617 VN.t3 VSUBS 1.96633f
C618 VN.n0 VSUBS 1.45563f
C619 VN.t1 VSUBS 1.96724f
C620 VN.t2 VSUBS 1.96633f
C621 VN.n1 VSUBS 2.9596f
.ends

