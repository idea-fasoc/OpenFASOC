* NGSPICE file created from diff_pair_sample_1633.ext - technology: sky130A

.subckt diff_pair_sample_1633 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t17 VN.t0 VDD2.t6 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=1.18635 pd=7.52 as=1.18635 ps=7.52 w=7.19 l=1.22
X1 B.t11 B.t9 B.t10 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=2.8041 pd=15.16 as=0 ps=0 w=7.19 l=1.22
X2 VTAIL.t4 VP.t0 VDD1.t9 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=1.18635 pd=7.52 as=1.18635 ps=7.52 w=7.19 l=1.22
X3 B.t8 B.t6 B.t7 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=2.8041 pd=15.16 as=0 ps=0 w=7.19 l=1.22
X4 B.t5 B.t3 B.t4 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=2.8041 pd=15.16 as=0 ps=0 w=7.19 l=1.22
X5 VTAIL.t0 VP.t1 VDD1.t8 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=1.18635 pd=7.52 as=1.18635 ps=7.52 w=7.19 l=1.22
X6 VDD2.t3 VN.t1 VTAIL.t16 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=1.18635 pd=7.52 as=1.18635 ps=7.52 w=7.19 l=1.22
X7 VTAIL.t5 VP.t2 VDD1.t7 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=1.18635 pd=7.52 as=1.18635 ps=7.52 w=7.19 l=1.22
X8 VTAIL.t15 VN.t2 VDD2.t9 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=1.18635 pd=7.52 as=1.18635 ps=7.52 w=7.19 l=1.22
X9 VDD1.t6 VP.t3 VTAIL.t18 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=1.18635 pd=7.52 as=1.18635 ps=7.52 w=7.19 l=1.22
X10 VTAIL.t14 VN.t3 VDD2.t5 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=1.18635 pd=7.52 as=1.18635 ps=7.52 w=7.19 l=1.22
X11 VDD1.t5 VP.t4 VTAIL.t3 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=2.8041 pd=15.16 as=1.18635 ps=7.52 w=7.19 l=1.22
X12 VDD1.t4 VP.t5 VTAIL.t6 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=2.8041 pd=15.16 as=1.18635 ps=7.52 w=7.19 l=1.22
X13 VDD2.t0 VN.t4 VTAIL.t13 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=1.18635 pd=7.52 as=2.8041 ps=15.16 w=7.19 l=1.22
X14 VDD2.t1 VN.t5 VTAIL.t12 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=2.8041 pd=15.16 as=1.18635 ps=7.52 w=7.19 l=1.22
X15 VDD1.t3 VP.t6 VTAIL.t7 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=1.18635 pd=7.52 as=1.18635 ps=7.52 w=7.19 l=1.22
X16 B.t2 B.t0 B.t1 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=2.8041 pd=15.16 as=0 ps=0 w=7.19 l=1.22
X17 VDD1.t2 VP.t7 VTAIL.t2 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=1.18635 pd=7.52 as=2.8041 ps=15.16 w=7.19 l=1.22
X18 VDD2.t4 VN.t6 VTAIL.t11 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=1.18635 pd=7.52 as=2.8041 ps=15.16 w=7.19 l=1.22
X19 VDD2.t2 VN.t7 VTAIL.t10 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=1.18635 pd=7.52 as=1.18635 ps=7.52 w=7.19 l=1.22
X20 VTAIL.t1 VP.t8 VDD1.t1 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=1.18635 pd=7.52 as=1.18635 ps=7.52 w=7.19 l=1.22
X21 VDD2.t8 VN.t8 VTAIL.t9 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=2.8041 pd=15.16 as=1.18635 ps=7.52 w=7.19 l=1.22
X22 VDD1.t0 VP.t9 VTAIL.t19 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=1.18635 pd=7.52 as=2.8041 ps=15.16 w=7.19 l=1.22
X23 VTAIL.t8 VN.t9 VDD2.t7 w_n2830_n2406# sky130_fd_pr__pfet_01v8 ad=1.18635 pd=7.52 as=1.18635 ps=7.52 w=7.19 l=1.22
R0 VN.n6 VN.t5 194.32
R1 VN.n28 VN.t4 194.32
R2 VN.n20 VN.t6 174.429
R3 VN.n42 VN.t8 174.429
R4 VN.n41 VN.n22 161.3
R5 VN.n40 VN.n39 161.3
R6 VN.n38 VN.n37 161.3
R7 VN.n36 VN.n24 161.3
R8 VN.n35 VN.n34 161.3
R9 VN.n33 VN.n32 161.3
R10 VN.n31 VN.n26 161.3
R11 VN.n30 VN.n29 161.3
R12 VN.n19 VN.n0 161.3
R13 VN.n18 VN.n17 161.3
R14 VN.n16 VN.n15 161.3
R15 VN.n14 VN.n2 161.3
R16 VN.n13 VN.n12 161.3
R17 VN.n11 VN.n10 161.3
R18 VN.n9 VN.n4 161.3
R19 VN.n8 VN.n7 161.3
R20 VN.n5 VN.t9 142.032
R21 VN.n3 VN.t7 142.032
R22 VN.n1 VN.t2 142.032
R23 VN.n27 VN.t3 142.032
R24 VN.n25 VN.t1 142.032
R25 VN.n23 VN.t0 142.032
R26 VN.n43 VN.n42 80.6037
R27 VN.n21 VN.n20 80.6037
R28 VN.n9 VN.n8 42.9216
R29 VN.n15 VN.n14 42.9216
R30 VN.n31 VN.n30 42.9216
R31 VN.n37 VN.n36 42.9216
R32 VN.n6 VN.n5 42.7694
R33 VN.n28 VN.n27 42.7694
R34 VN VN.n43 42.4119
R35 VN.n10 VN.n9 38.0652
R36 VN.n14 VN.n13 38.0652
R37 VN.n32 VN.n31 38.0652
R38 VN.n36 VN.n35 38.0652
R39 VN.n20 VN.n19 35.055
R40 VN.n42 VN.n41 35.055
R41 VN.n19 VN.n18 33.2089
R42 VN.n41 VN.n40 33.2089
R43 VN.n29 VN.n28 29.263
R44 VN.n7 VN.n6 29.263
R45 VN.n8 VN.n5 14.6807
R46 VN.n15 VN.n1 14.6807
R47 VN.n30 VN.n27 14.6807
R48 VN.n37 VN.n23 14.6807
R49 VN.n10 VN.n3 12.234
R50 VN.n13 VN.n3 12.234
R51 VN.n35 VN.n25 12.234
R52 VN.n32 VN.n25 12.234
R53 VN.n18 VN.n1 9.7873
R54 VN.n40 VN.n23 9.7873
R55 VN.n43 VN.n22 0.285035
R56 VN.n21 VN.n0 0.285035
R57 VN.n39 VN.n22 0.189894
R58 VN.n39 VN.n38 0.189894
R59 VN.n38 VN.n24 0.189894
R60 VN.n34 VN.n24 0.189894
R61 VN.n34 VN.n33 0.189894
R62 VN.n33 VN.n26 0.189894
R63 VN.n29 VN.n26 0.189894
R64 VN.n7 VN.n4 0.189894
R65 VN.n11 VN.n4 0.189894
R66 VN.n12 VN.n11 0.189894
R67 VN.n12 VN.n2 0.189894
R68 VN.n16 VN.n2 0.189894
R69 VN.n17 VN.n16 0.189894
R70 VN.n17 VN.n0 0.189894
R71 VN VN.n21 0.146778
R72 VDD2.n70 VDD2.n69 585
R73 VDD2.n68 VDD2.n67 585
R74 VDD2.n43 VDD2.n42 585
R75 VDD2.n62 VDD2.n61 585
R76 VDD2.n60 VDD2.n59 585
R77 VDD2.n47 VDD2.n46 585
R78 VDD2.n54 VDD2.n53 585
R79 VDD2.n52 VDD2.n51 585
R80 VDD2.n13 VDD2.n12 585
R81 VDD2.n15 VDD2.n14 585
R82 VDD2.n8 VDD2.n7 585
R83 VDD2.n21 VDD2.n20 585
R84 VDD2.n23 VDD2.n22 585
R85 VDD2.n4 VDD2.n3 585
R86 VDD2.n29 VDD2.n28 585
R87 VDD2.n31 VDD2.n30 585
R88 VDD2.n69 VDD2.n39 498.474
R89 VDD2.n30 VDD2.n0 498.474
R90 VDD2.n50 VDD2.t8 329.053
R91 VDD2.n11 VDD2.t1 329.053
R92 VDD2.n69 VDD2.n68 171.744
R93 VDD2.n68 VDD2.n42 171.744
R94 VDD2.n61 VDD2.n42 171.744
R95 VDD2.n61 VDD2.n60 171.744
R96 VDD2.n60 VDD2.n46 171.744
R97 VDD2.n53 VDD2.n46 171.744
R98 VDD2.n53 VDD2.n52 171.744
R99 VDD2.n14 VDD2.n13 171.744
R100 VDD2.n14 VDD2.n7 171.744
R101 VDD2.n21 VDD2.n7 171.744
R102 VDD2.n22 VDD2.n21 171.744
R103 VDD2.n22 VDD2.n3 171.744
R104 VDD2.n29 VDD2.n3 171.744
R105 VDD2.n30 VDD2.n29 171.744
R106 VDD2.n38 VDD2.n37 87.9189
R107 VDD2 VDD2.n77 87.916
R108 VDD2.n76 VDD2.n75 86.9722
R109 VDD2.n36 VDD2.n35 86.972
R110 VDD2.n52 VDD2.t8 85.8723
R111 VDD2.n13 VDD2.t1 85.8723
R112 VDD2.n36 VDD2.n34 52.3337
R113 VDD2.n74 VDD2.n73 50.9975
R114 VDD2.n74 VDD2.n38 36.2606
R115 VDD2.n71 VDD2.n70 12.8005
R116 VDD2.n32 VDD2.n31 12.8005
R117 VDD2.n67 VDD2.n41 12.0247
R118 VDD2.n28 VDD2.n2 12.0247
R119 VDD2.n66 VDD2.n43 11.249
R120 VDD2.n27 VDD2.n4 11.249
R121 VDD2.n51 VDD2.n50 10.7237
R122 VDD2.n12 VDD2.n11 10.7237
R123 VDD2.n63 VDD2.n62 10.4732
R124 VDD2.n24 VDD2.n23 10.4732
R125 VDD2.n59 VDD2.n45 9.69747
R126 VDD2.n20 VDD2.n6 9.69747
R127 VDD2.n73 VDD2.n72 9.45567
R128 VDD2.n34 VDD2.n33 9.45567
R129 VDD2.n49 VDD2.n48 9.3005
R130 VDD2.n56 VDD2.n55 9.3005
R131 VDD2.n58 VDD2.n57 9.3005
R132 VDD2.n45 VDD2.n44 9.3005
R133 VDD2.n64 VDD2.n63 9.3005
R134 VDD2.n66 VDD2.n65 9.3005
R135 VDD2.n41 VDD2.n40 9.3005
R136 VDD2.n72 VDD2.n71 9.3005
R137 VDD2.n10 VDD2.n9 9.3005
R138 VDD2.n17 VDD2.n16 9.3005
R139 VDD2.n19 VDD2.n18 9.3005
R140 VDD2.n6 VDD2.n5 9.3005
R141 VDD2.n25 VDD2.n24 9.3005
R142 VDD2.n27 VDD2.n26 9.3005
R143 VDD2.n2 VDD2.n1 9.3005
R144 VDD2.n33 VDD2.n32 9.3005
R145 VDD2.n58 VDD2.n47 8.92171
R146 VDD2.n19 VDD2.n8 8.92171
R147 VDD2.n55 VDD2.n54 8.14595
R148 VDD2.n16 VDD2.n15 8.14595
R149 VDD2.n73 VDD2.n39 7.75445
R150 VDD2.n34 VDD2.n0 7.75445
R151 VDD2.n51 VDD2.n49 7.3702
R152 VDD2.n12 VDD2.n10 7.3702
R153 VDD2.n71 VDD2.n39 6.08283
R154 VDD2.n32 VDD2.n0 6.08283
R155 VDD2.n54 VDD2.n49 5.81868
R156 VDD2.n15 VDD2.n10 5.81868
R157 VDD2.n55 VDD2.n47 5.04292
R158 VDD2.n16 VDD2.n8 5.04292
R159 VDD2.n77 VDD2.t5 4.52136
R160 VDD2.n77 VDD2.t0 4.52136
R161 VDD2.n75 VDD2.t6 4.52136
R162 VDD2.n75 VDD2.t3 4.52136
R163 VDD2.n37 VDD2.t9 4.52136
R164 VDD2.n37 VDD2.t4 4.52136
R165 VDD2.n35 VDD2.t7 4.52136
R166 VDD2.n35 VDD2.t2 4.52136
R167 VDD2.n59 VDD2.n58 4.26717
R168 VDD2.n20 VDD2.n19 4.26717
R169 VDD2.n62 VDD2.n45 3.49141
R170 VDD2.n23 VDD2.n6 3.49141
R171 VDD2.n63 VDD2.n43 2.71565
R172 VDD2.n24 VDD2.n4 2.71565
R173 VDD2.n50 VDD2.n48 2.41305
R174 VDD2.n11 VDD2.n9 2.41305
R175 VDD2.n67 VDD2.n66 1.93989
R176 VDD2.n28 VDD2.n27 1.93989
R177 VDD2.n76 VDD2.n74 1.33671
R178 VDD2.n70 VDD2.n41 1.16414
R179 VDD2.n31 VDD2.n2 1.16414
R180 VDD2 VDD2.n76 0.392741
R181 VDD2.n38 VDD2.n36 0.279206
R182 VDD2.n72 VDD2.n40 0.155672
R183 VDD2.n65 VDD2.n40 0.155672
R184 VDD2.n65 VDD2.n64 0.155672
R185 VDD2.n64 VDD2.n44 0.155672
R186 VDD2.n57 VDD2.n44 0.155672
R187 VDD2.n57 VDD2.n56 0.155672
R188 VDD2.n56 VDD2.n48 0.155672
R189 VDD2.n17 VDD2.n9 0.155672
R190 VDD2.n18 VDD2.n17 0.155672
R191 VDD2.n18 VDD2.n5 0.155672
R192 VDD2.n25 VDD2.n5 0.155672
R193 VDD2.n26 VDD2.n25 0.155672
R194 VDD2.n26 VDD2.n1 0.155672
R195 VDD2.n33 VDD2.n1 0.155672
R196 VTAIL.n135 VTAIL.n134 585
R197 VTAIL.n137 VTAIL.n136 585
R198 VTAIL.n130 VTAIL.n129 585
R199 VTAIL.n143 VTAIL.n142 585
R200 VTAIL.n145 VTAIL.n144 585
R201 VTAIL.n126 VTAIL.n125 585
R202 VTAIL.n151 VTAIL.n150 585
R203 VTAIL.n153 VTAIL.n152 585
R204 VTAIL.n15 VTAIL.n14 585
R205 VTAIL.n17 VTAIL.n16 585
R206 VTAIL.n10 VTAIL.n9 585
R207 VTAIL.n23 VTAIL.n22 585
R208 VTAIL.n25 VTAIL.n24 585
R209 VTAIL.n6 VTAIL.n5 585
R210 VTAIL.n31 VTAIL.n30 585
R211 VTAIL.n33 VTAIL.n32 585
R212 VTAIL.n117 VTAIL.n116 585
R213 VTAIL.n115 VTAIL.n114 585
R214 VTAIL.n90 VTAIL.n89 585
R215 VTAIL.n109 VTAIL.n108 585
R216 VTAIL.n107 VTAIL.n106 585
R217 VTAIL.n94 VTAIL.n93 585
R218 VTAIL.n101 VTAIL.n100 585
R219 VTAIL.n99 VTAIL.n98 585
R220 VTAIL.n77 VTAIL.n76 585
R221 VTAIL.n75 VTAIL.n74 585
R222 VTAIL.n50 VTAIL.n49 585
R223 VTAIL.n69 VTAIL.n68 585
R224 VTAIL.n67 VTAIL.n66 585
R225 VTAIL.n54 VTAIL.n53 585
R226 VTAIL.n61 VTAIL.n60 585
R227 VTAIL.n59 VTAIL.n58 585
R228 VTAIL.n152 VTAIL.n122 498.474
R229 VTAIL.n32 VTAIL.n2 498.474
R230 VTAIL.n116 VTAIL.n86 498.474
R231 VTAIL.n76 VTAIL.n46 498.474
R232 VTAIL.n133 VTAIL.t11 329.053
R233 VTAIL.n13 VTAIL.t2 329.053
R234 VTAIL.n97 VTAIL.t19 329.053
R235 VTAIL.n57 VTAIL.t13 329.053
R236 VTAIL.n136 VTAIL.n135 171.744
R237 VTAIL.n136 VTAIL.n129 171.744
R238 VTAIL.n143 VTAIL.n129 171.744
R239 VTAIL.n144 VTAIL.n143 171.744
R240 VTAIL.n144 VTAIL.n125 171.744
R241 VTAIL.n151 VTAIL.n125 171.744
R242 VTAIL.n152 VTAIL.n151 171.744
R243 VTAIL.n16 VTAIL.n15 171.744
R244 VTAIL.n16 VTAIL.n9 171.744
R245 VTAIL.n23 VTAIL.n9 171.744
R246 VTAIL.n24 VTAIL.n23 171.744
R247 VTAIL.n24 VTAIL.n5 171.744
R248 VTAIL.n31 VTAIL.n5 171.744
R249 VTAIL.n32 VTAIL.n31 171.744
R250 VTAIL.n116 VTAIL.n115 171.744
R251 VTAIL.n115 VTAIL.n89 171.744
R252 VTAIL.n108 VTAIL.n89 171.744
R253 VTAIL.n108 VTAIL.n107 171.744
R254 VTAIL.n107 VTAIL.n93 171.744
R255 VTAIL.n100 VTAIL.n93 171.744
R256 VTAIL.n100 VTAIL.n99 171.744
R257 VTAIL.n76 VTAIL.n75 171.744
R258 VTAIL.n75 VTAIL.n49 171.744
R259 VTAIL.n68 VTAIL.n49 171.744
R260 VTAIL.n68 VTAIL.n67 171.744
R261 VTAIL.n67 VTAIL.n53 171.744
R262 VTAIL.n60 VTAIL.n53 171.744
R263 VTAIL.n60 VTAIL.n59 171.744
R264 VTAIL.n135 VTAIL.t11 85.8723
R265 VTAIL.n15 VTAIL.t2 85.8723
R266 VTAIL.n99 VTAIL.t19 85.8723
R267 VTAIL.n59 VTAIL.t13 85.8723
R268 VTAIL.n85 VTAIL.n84 70.2934
R269 VTAIL.n83 VTAIL.n82 70.2934
R270 VTAIL.n45 VTAIL.n44 70.2934
R271 VTAIL.n43 VTAIL.n42 70.2934
R272 VTAIL.n159 VTAIL.n158 70.2933
R273 VTAIL.n1 VTAIL.n0 70.2933
R274 VTAIL.n39 VTAIL.n38 70.2933
R275 VTAIL.n41 VTAIL.n40 70.2933
R276 VTAIL.n157 VTAIL.n156 34.3187
R277 VTAIL.n37 VTAIL.n36 34.3187
R278 VTAIL.n121 VTAIL.n120 34.3187
R279 VTAIL.n81 VTAIL.n80 34.3187
R280 VTAIL.n43 VTAIL.n41 21.2376
R281 VTAIL.n157 VTAIL.n121 19.9014
R282 VTAIL.n154 VTAIL.n153 12.8005
R283 VTAIL.n34 VTAIL.n33 12.8005
R284 VTAIL.n118 VTAIL.n117 12.8005
R285 VTAIL.n78 VTAIL.n77 12.8005
R286 VTAIL.n150 VTAIL.n124 12.0247
R287 VTAIL.n30 VTAIL.n4 12.0247
R288 VTAIL.n114 VTAIL.n88 12.0247
R289 VTAIL.n74 VTAIL.n48 12.0247
R290 VTAIL.n149 VTAIL.n126 11.249
R291 VTAIL.n29 VTAIL.n6 11.249
R292 VTAIL.n113 VTAIL.n90 11.249
R293 VTAIL.n73 VTAIL.n50 11.249
R294 VTAIL.n134 VTAIL.n133 10.7237
R295 VTAIL.n14 VTAIL.n13 10.7237
R296 VTAIL.n98 VTAIL.n97 10.7237
R297 VTAIL.n58 VTAIL.n57 10.7237
R298 VTAIL.n146 VTAIL.n145 10.4732
R299 VTAIL.n26 VTAIL.n25 10.4732
R300 VTAIL.n110 VTAIL.n109 10.4732
R301 VTAIL.n70 VTAIL.n69 10.4732
R302 VTAIL.n142 VTAIL.n128 9.69747
R303 VTAIL.n22 VTAIL.n8 9.69747
R304 VTAIL.n106 VTAIL.n92 9.69747
R305 VTAIL.n66 VTAIL.n52 9.69747
R306 VTAIL.n156 VTAIL.n155 9.45567
R307 VTAIL.n36 VTAIL.n35 9.45567
R308 VTAIL.n120 VTAIL.n119 9.45567
R309 VTAIL.n80 VTAIL.n79 9.45567
R310 VTAIL.n132 VTAIL.n131 9.3005
R311 VTAIL.n139 VTAIL.n138 9.3005
R312 VTAIL.n141 VTAIL.n140 9.3005
R313 VTAIL.n128 VTAIL.n127 9.3005
R314 VTAIL.n147 VTAIL.n146 9.3005
R315 VTAIL.n149 VTAIL.n148 9.3005
R316 VTAIL.n124 VTAIL.n123 9.3005
R317 VTAIL.n155 VTAIL.n154 9.3005
R318 VTAIL.n12 VTAIL.n11 9.3005
R319 VTAIL.n19 VTAIL.n18 9.3005
R320 VTAIL.n21 VTAIL.n20 9.3005
R321 VTAIL.n8 VTAIL.n7 9.3005
R322 VTAIL.n27 VTAIL.n26 9.3005
R323 VTAIL.n29 VTAIL.n28 9.3005
R324 VTAIL.n4 VTAIL.n3 9.3005
R325 VTAIL.n35 VTAIL.n34 9.3005
R326 VTAIL.n96 VTAIL.n95 9.3005
R327 VTAIL.n103 VTAIL.n102 9.3005
R328 VTAIL.n105 VTAIL.n104 9.3005
R329 VTAIL.n92 VTAIL.n91 9.3005
R330 VTAIL.n111 VTAIL.n110 9.3005
R331 VTAIL.n113 VTAIL.n112 9.3005
R332 VTAIL.n88 VTAIL.n87 9.3005
R333 VTAIL.n119 VTAIL.n118 9.3005
R334 VTAIL.n56 VTAIL.n55 9.3005
R335 VTAIL.n63 VTAIL.n62 9.3005
R336 VTAIL.n65 VTAIL.n64 9.3005
R337 VTAIL.n52 VTAIL.n51 9.3005
R338 VTAIL.n71 VTAIL.n70 9.3005
R339 VTAIL.n73 VTAIL.n72 9.3005
R340 VTAIL.n48 VTAIL.n47 9.3005
R341 VTAIL.n79 VTAIL.n78 9.3005
R342 VTAIL.n141 VTAIL.n130 8.92171
R343 VTAIL.n21 VTAIL.n10 8.92171
R344 VTAIL.n105 VTAIL.n94 8.92171
R345 VTAIL.n65 VTAIL.n54 8.92171
R346 VTAIL.n138 VTAIL.n137 8.14595
R347 VTAIL.n18 VTAIL.n17 8.14595
R348 VTAIL.n102 VTAIL.n101 8.14595
R349 VTAIL.n62 VTAIL.n61 8.14595
R350 VTAIL.n156 VTAIL.n122 7.75445
R351 VTAIL.n36 VTAIL.n2 7.75445
R352 VTAIL.n120 VTAIL.n86 7.75445
R353 VTAIL.n80 VTAIL.n46 7.75445
R354 VTAIL.n134 VTAIL.n132 7.3702
R355 VTAIL.n14 VTAIL.n12 7.3702
R356 VTAIL.n98 VTAIL.n96 7.3702
R357 VTAIL.n58 VTAIL.n56 7.3702
R358 VTAIL.n154 VTAIL.n122 6.08283
R359 VTAIL.n34 VTAIL.n2 6.08283
R360 VTAIL.n118 VTAIL.n86 6.08283
R361 VTAIL.n78 VTAIL.n46 6.08283
R362 VTAIL.n137 VTAIL.n132 5.81868
R363 VTAIL.n17 VTAIL.n12 5.81868
R364 VTAIL.n101 VTAIL.n96 5.81868
R365 VTAIL.n61 VTAIL.n56 5.81868
R366 VTAIL.n138 VTAIL.n130 5.04292
R367 VTAIL.n18 VTAIL.n10 5.04292
R368 VTAIL.n102 VTAIL.n94 5.04292
R369 VTAIL.n62 VTAIL.n54 5.04292
R370 VTAIL.n158 VTAIL.t10 4.52136
R371 VTAIL.n158 VTAIL.t15 4.52136
R372 VTAIL.n0 VTAIL.t12 4.52136
R373 VTAIL.n0 VTAIL.t8 4.52136
R374 VTAIL.n38 VTAIL.t7 4.52136
R375 VTAIL.n38 VTAIL.t4 4.52136
R376 VTAIL.n40 VTAIL.t3 4.52136
R377 VTAIL.n40 VTAIL.t1 4.52136
R378 VTAIL.n84 VTAIL.t18 4.52136
R379 VTAIL.n84 VTAIL.t0 4.52136
R380 VTAIL.n82 VTAIL.t6 4.52136
R381 VTAIL.n82 VTAIL.t5 4.52136
R382 VTAIL.n44 VTAIL.t16 4.52136
R383 VTAIL.n44 VTAIL.t14 4.52136
R384 VTAIL.n42 VTAIL.t9 4.52136
R385 VTAIL.n42 VTAIL.t17 4.52136
R386 VTAIL.n142 VTAIL.n141 4.26717
R387 VTAIL.n22 VTAIL.n21 4.26717
R388 VTAIL.n106 VTAIL.n105 4.26717
R389 VTAIL.n66 VTAIL.n65 4.26717
R390 VTAIL.n145 VTAIL.n128 3.49141
R391 VTAIL.n25 VTAIL.n8 3.49141
R392 VTAIL.n109 VTAIL.n92 3.49141
R393 VTAIL.n69 VTAIL.n52 3.49141
R394 VTAIL.n146 VTAIL.n126 2.71565
R395 VTAIL.n26 VTAIL.n6 2.71565
R396 VTAIL.n110 VTAIL.n90 2.71565
R397 VTAIL.n70 VTAIL.n50 2.71565
R398 VTAIL.n133 VTAIL.n131 2.41305
R399 VTAIL.n13 VTAIL.n11 2.41305
R400 VTAIL.n97 VTAIL.n95 2.41305
R401 VTAIL.n57 VTAIL.n55 2.41305
R402 VTAIL.n150 VTAIL.n149 1.93989
R403 VTAIL.n30 VTAIL.n29 1.93989
R404 VTAIL.n114 VTAIL.n113 1.93989
R405 VTAIL.n74 VTAIL.n73 1.93989
R406 VTAIL.n45 VTAIL.n43 1.33671
R407 VTAIL.n81 VTAIL.n45 1.33671
R408 VTAIL.n85 VTAIL.n83 1.33671
R409 VTAIL.n121 VTAIL.n85 1.33671
R410 VTAIL.n41 VTAIL.n39 1.33671
R411 VTAIL.n39 VTAIL.n37 1.33671
R412 VTAIL.n159 VTAIL.n157 1.33671
R413 VTAIL.n153 VTAIL.n124 1.16414
R414 VTAIL.n33 VTAIL.n4 1.16414
R415 VTAIL.n117 VTAIL.n88 1.16414
R416 VTAIL.n77 VTAIL.n48 1.16414
R417 VTAIL.n83 VTAIL.n81 1.13843
R418 VTAIL.n37 VTAIL.n1 1.13843
R419 VTAIL VTAIL.n1 1.06084
R420 VTAIL VTAIL.n159 0.276362
R421 VTAIL.n139 VTAIL.n131 0.155672
R422 VTAIL.n140 VTAIL.n139 0.155672
R423 VTAIL.n140 VTAIL.n127 0.155672
R424 VTAIL.n147 VTAIL.n127 0.155672
R425 VTAIL.n148 VTAIL.n147 0.155672
R426 VTAIL.n148 VTAIL.n123 0.155672
R427 VTAIL.n155 VTAIL.n123 0.155672
R428 VTAIL.n19 VTAIL.n11 0.155672
R429 VTAIL.n20 VTAIL.n19 0.155672
R430 VTAIL.n20 VTAIL.n7 0.155672
R431 VTAIL.n27 VTAIL.n7 0.155672
R432 VTAIL.n28 VTAIL.n27 0.155672
R433 VTAIL.n28 VTAIL.n3 0.155672
R434 VTAIL.n35 VTAIL.n3 0.155672
R435 VTAIL.n119 VTAIL.n87 0.155672
R436 VTAIL.n112 VTAIL.n87 0.155672
R437 VTAIL.n112 VTAIL.n111 0.155672
R438 VTAIL.n111 VTAIL.n91 0.155672
R439 VTAIL.n104 VTAIL.n91 0.155672
R440 VTAIL.n104 VTAIL.n103 0.155672
R441 VTAIL.n103 VTAIL.n95 0.155672
R442 VTAIL.n79 VTAIL.n47 0.155672
R443 VTAIL.n72 VTAIL.n47 0.155672
R444 VTAIL.n72 VTAIL.n71 0.155672
R445 VTAIL.n71 VTAIL.n51 0.155672
R446 VTAIL.n64 VTAIL.n51 0.155672
R447 VTAIL.n64 VTAIL.n63 0.155672
R448 VTAIL.n63 VTAIL.n55 0.155672
R449 B.n296 B.n295 585
R450 B.n294 B.n93 585
R451 B.n293 B.n292 585
R452 B.n291 B.n94 585
R453 B.n290 B.n289 585
R454 B.n288 B.n95 585
R455 B.n287 B.n286 585
R456 B.n285 B.n96 585
R457 B.n284 B.n283 585
R458 B.n282 B.n97 585
R459 B.n281 B.n280 585
R460 B.n279 B.n98 585
R461 B.n278 B.n277 585
R462 B.n276 B.n99 585
R463 B.n275 B.n274 585
R464 B.n273 B.n100 585
R465 B.n272 B.n271 585
R466 B.n270 B.n101 585
R467 B.n269 B.n268 585
R468 B.n267 B.n102 585
R469 B.n266 B.n265 585
R470 B.n264 B.n103 585
R471 B.n263 B.n262 585
R472 B.n261 B.n104 585
R473 B.n260 B.n259 585
R474 B.n258 B.n105 585
R475 B.n257 B.n256 585
R476 B.n255 B.n106 585
R477 B.n254 B.n253 585
R478 B.n249 B.n107 585
R479 B.n248 B.n247 585
R480 B.n246 B.n108 585
R481 B.n245 B.n244 585
R482 B.n243 B.n109 585
R483 B.n242 B.n241 585
R484 B.n240 B.n110 585
R485 B.n239 B.n238 585
R486 B.n236 B.n111 585
R487 B.n235 B.n234 585
R488 B.n233 B.n114 585
R489 B.n232 B.n231 585
R490 B.n230 B.n115 585
R491 B.n229 B.n228 585
R492 B.n227 B.n116 585
R493 B.n226 B.n225 585
R494 B.n224 B.n117 585
R495 B.n223 B.n222 585
R496 B.n221 B.n118 585
R497 B.n220 B.n219 585
R498 B.n218 B.n119 585
R499 B.n217 B.n216 585
R500 B.n215 B.n120 585
R501 B.n214 B.n213 585
R502 B.n212 B.n121 585
R503 B.n211 B.n210 585
R504 B.n209 B.n122 585
R505 B.n208 B.n207 585
R506 B.n206 B.n123 585
R507 B.n205 B.n204 585
R508 B.n203 B.n124 585
R509 B.n202 B.n201 585
R510 B.n200 B.n125 585
R511 B.n199 B.n198 585
R512 B.n197 B.n126 585
R513 B.n196 B.n195 585
R514 B.n297 B.n92 585
R515 B.n299 B.n298 585
R516 B.n300 B.n91 585
R517 B.n302 B.n301 585
R518 B.n303 B.n90 585
R519 B.n305 B.n304 585
R520 B.n306 B.n89 585
R521 B.n308 B.n307 585
R522 B.n309 B.n88 585
R523 B.n311 B.n310 585
R524 B.n312 B.n87 585
R525 B.n314 B.n313 585
R526 B.n315 B.n86 585
R527 B.n317 B.n316 585
R528 B.n318 B.n85 585
R529 B.n320 B.n319 585
R530 B.n321 B.n84 585
R531 B.n323 B.n322 585
R532 B.n324 B.n83 585
R533 B.n326 B.n325 585
R534 B.n327 B.n82 585
R535 B.n329 B.n328 585
R536 B.n330 B.n81 585
R537 B.n332 B.n331 585
R538 B.n333 B.n80 585
R539 B.n335 B.n334 585
R540 B.n336 B.n79 585
R541 B.n338 B.n337 585
R542 B.n339 B.n78 585
R543 B.n341 B.n340 585
R544 B.n342 B.n77 585
R545 B.n344 B.n343 585
R546 B.n345 B.n76 585
R547 B.n347 B.n346 585
R548 B.n348 B.n75 585
R549 B.n350 B.n349 585
R550 B.n351 B.n74 585
R551 B.n353 B.n352 585
R552 B.n354 B.n73 585
R553 B.n356 B.n355 585
R554 B.n357 B.n72 585
R555 B.n359 B.n358 585
R556 B.n360 B.n71 585
R557 B.n362 B.n361 585
R558 B.n363 B.n70 585
R559 B.n365 B.n364 585
R560 B.n366 B.n69 585
R561 B.n368 B.n367 585
R562 B.n369 B.n68 585
R563 B.n371 B.n370 585
R564 B.n372 B.n67 585
R565 B.n374 B.n373 585
R566 B.n375 B.n66 585
R567 B.n377 B.n376 585
R568 B.n378 B.n65 585
R569 B.n380 B.n379 585
R570 B.n381 B.n64 585
R571 B.n383 B.n382 585
R572 B.n384 B.n63 585
R573 B.n386 B.n385 585
R574 B.n387 B.n62 585
R575 B.n389 B.n388 585
R576 B.n390 B.n61 585
R577 B.n392 B.n391 585
R578 B.n393 B.n60 585
R579 B.n395 B.n394 585
R580 B.n396 B.n59 585
R581 B.n398 B.n397 585
R582 B.n399 B.n58 585
R583 B.n401 B.n400 585
R584 B.n402 B.n57 585
R585 B.n404 B.n403 585
R586 B.n503 B.n502 585
R587 B.n501 B.n20 585
R588 B.n500 B.n499 585
R589 B.n498 B.n21 585
R590 B.n497 B.n496 585
R591 B.n495 B.n22 585
R592 B.n494 B.n493 585
R593 B.n492 B.n23 585
R594 B.n491 B.n490 585
R595 B.n489 B.n24 585
R596 B.n488 B.n487 585
R597 B.n486 B.n25 585
R598 B.n485 B.n484 585
R599 B.n483 B.n26 585
R600 B.n482 B.n481 585
R601 B.n480 B.n27 585
R602 B.n479 B.n478 585
R603 B.n477 B.n28 585
R604 B.n476 B.n475 585
R605 B.n474 B.n29 585
R606 B.n473 B.n472 585
R607 B.n471 B.n30 585
R608 B.n470 B.n469 585
R609 B.n468 B.n31 585
R610 B.n467 B.n466 585
R611 B.n465 B.n32 585
R612 B.n464 B.n463 585
R613 B.n462 B.n33 585
R614 B.n460 B.n459 585
R615 B.n458 B.n36 585
R616 B.n457 B.n456 585
R617 B.n455 B.n37 585
R618 B.n454 B.n453 585
R619 B.n452 B.n38 585
R620 B.n451 B.n450 585
R621 B.n449 B.n39 585
R622 B.n448 B.n447 585
R623 B.n446 B.n445 585
R624 B.n444 B.n43 585
R625 B.n443 B.n442 585
R626 B.n441 B.n44 585
R627 B.n440 B.n439 585
R628 B.n438 B.n45 585
R629 B.n437 B.n436 585
R630 B.n435 B.n46 585
R631 B.n434 B.n433 585
R632 B.n432 B.n47 585
R633 B.n431 B.n430 585
R634 B.n429 B.n48 585
R635 B.n428 B.n427 585
R636 B.n426 B.n49 585
R637 B.n425 B.n424 585
R638 B.n423 B.n50 585
R639 B.n422 B.n421 585
R640 B.n420 B.n51 585
R641 B.n419 B.n418 585
R642 B.n417 B.n52 585
R643 B.n416 B.n415 585
R644 B.n414 B.n53 585
R645 B.n413 B.n412 585
R646 B.n411 B.n54 585
R647 B.n410 B.n409 585
R648 B.n408 B.n55 585
R649 B.n407 B.n406 585
R650 B.n405 B.n56 585
R651 B.n504 B.n19 585
R652 B.n506 B.n505 585
R653 B.n507 B.n18 585
R654 B.n509 B.n508 585
R655 B.n510 B.n17 585
R656 B.n512 B.n511 585
R657 B.n513 B.n16 585
R658 B.n515 B.n514 585
R659 B.n516 B.n15 585
R660 B.n518 B.n517 585
R661 B.n519 B.n14 585
R662 B.n521 B.n520 585
R663 B.n522 B.n13 585
R664 B.n524 B.n523 585
R665 B.n525 B.n12 585
R666 B.n527 B.n526 585
R667 B.n528 B.n11 585
R668 B.n530 B.n529 585
R669 B.n531 B.n10 585
R670 B.n533 B.n532 585
R671 B.n534 B.n9 585
R672 B.n536 B.n535 585
R673 B.n537 B.n8 585
R674 B.n539 B.n538 585
R675 B.n540 B.n7 585
R676 B.n542 B.n541 585
R677 B.n543 B.n6 585
R678 B.n545 B.n544 585
R679 B.n546 B.n5 585
R680 B.n548 B.n547 585
R681 B.n549 B.n4 585
R682 B.n551 B.n550 585
R683 B.n552 B.n3 585
R684 B.n554 B.n553 585
R685 B.n555 B.n0 585
R686 B.n2 B.n1 585
R687 B.n145 B.n144 585
R688 B.n146 B.n143 585
R689 B.n148 B.n147 585
R690 B.n149 B.n142 585
R691 B.n151 B.n150 585
R692 B.n152 B.n141 585
R693 B.n154 B.n153 585
R694 B.n155 B.n140 585
R695 B.n157 B.n156 585
R696 B.n158 B.n139 585
R697 B.n160 B.n159 585
R698 B.n161 B.n138 585
R699 B.n163 B.n162 585
R700 B.n164 B.n137 585
R701 B.n166 B.n165 585
R702 B.n167 B.n136 585
R703 B.n169 B.n168 585
R704 B.n170 B.n135 585
R705 B.n172 B.n171 585
R706 B.n173 B.n134 585
R707 B.n175 B.n174 585
R708 B.n176 B.n133 585
R709 B.n178 B.n177 585
R710 B.n179 B.n132 585
R711 B.n181 B.n180 585
R712 B.n182 B.n131 585
R713 B.n184 B.n183 585
R714 B.n185 B.n130 585
R715 B.n187 B.n186 585
R716 B.n188 B.n129 585
R717 B.n190 B.n189 585
R718 B.n191 B.n128 585
R719 B.n193 B.n192 585
R720 B.n194 B.n127 585
R721 B.n196 B.n127 454.062
R722 B.n297 B.n296 454.062
R723 B.n405 B.n404 454.062
R724 B.n502 B.n19 454.062
R725 B.n112 B.t3 346.252
R726 B.n250 B.t9 346.252
R727 B.n40 B.t6 346.252
R728 B.n34 B.t0 346.252
R729 B.n250 B.t10 319.06
R730 B.n40 B.t8 319.06
R731 B.n112 B.t4 319.06
R732 B.n34 B.t2 319.06
R733 B.n251 B.t11 288.998
R734 B.n41 B.t7 288.998
R735 B.n113 B.t5 288.998
R736 B.n35 B.t1 288.998
R737 B.n557 B.n556 256.663
R738 B.n556 B.n555 235.042
R739 B.n556 B.n2 235.042
R740 B.n197 B.n196 163.367
R741 B.n198 B.n197 163.367
R742 B.n198 B.n125 163.367
R743 B.n202 B.n125 163.367
R744 B.n203 B.n202 163.367
R745 B.n204 B.n203 163.367
R746 B.n204 B.n123 163.367
R747 B.n208 B.n123 163.367
R748 B.n209 B.n208 163.367
R749 B.n210 B.n209 163.367
R750 B.n210 B.n121 163.367
R751 B.n214 B.n121 163.367
R752 B.n215 B.n214 163.367
R753 B.n216 B.n215 163.367
R754 B.n216 B.n119 163.367
R755 B.n220 B.n119 163.367
R756 B.n221 B.n220 163.367
R757 B.n222 B.n221 163.367
R758 B.n222 B.n117 163.367
R759 B.n226 B.n117 163.367
R760 B.n227 B.n226 163.367
R761 B.n228 B.n227 163.367
R762 B.n228 B.n115 163.367
R763 B.n232 B.n115 163.367
R764 B.n233 B.n232 163.367
R765 B.n234 B.n233 163.367
R766 B.n234 B.n111 163.367
R767 B.n239 B.n111 163.367
R768 B.n240 B.n239 163.367
R769 B.n241 B.n240 163.367
R770 B.n241 B.n109 163.367
R771 B.n245 B.n109 163.367
R772 B.n246 B.n245 163.367
R773 B.n247 B.n246 163.367
R774 B.n247 B.n107 163.367
R775 B.n254 B.n107 163.367
R776 B.n255 B.n254 163.367
R777 B.n256 B.n255 163.367
R778 B.n256 B.n105 163.367
R779 B.n260 B.n105 163.367
R780 B.n261 B.n260 163.367
R781 B.n262 B.n261 163.367
R782 B.n262 B.n103 163.367
R783 B.n266 B.n103 163.367
R784 B.n267 B.n266 163.367
R785 B.n268 B.n267 163.367
R786 B.n268 B.n101 163.367
R787 B.n272 B.n101 163.367
R788 B.n273 B.n272 163.367
R789 B.n274 B.n273 163.367
R790 B.n274 B.n99 163.367
R791 B.n278 B.n99 163.367
R792 B.n279 B.n278 163.367
R793 B.n280 B.n279 163.367
R794 B.n280 B.n97 163.367
R795 B.n284 B.n97 163.367
R796 B.n285 B.n284 163.367
R797 B.n286 B.n285 163.367
R798 B.n286 B.n95 163.367
R799 B.n290 B.n95 163.367
R800 B.n291 B.n290 163.367
R801 B.n292 B.n291 163.367
R802 B.n292 B.n93 163.367
R803 B.n296 B.n93 163.367
R804 B.n404 B.n57 163.367
R805 B.n400 B.n57 163.367
R806 B.n400 B.n399 163.367
R807 B.n399 B.n398 163.367
R808 B.n398 B.n59 163.367
R809 B.n394 B.n59 163.367
R810 B.n394 B.n393 163.367
R811 B.n393 B.n392 163.367
R812 B.n392 B.n61 163.367
R813 B.n388 B.n61 163.367
R814 B.n388 B.n387 163.367
R815 B.n387 B.n386 163.367
R816 B.n386 B.n63 163.367
R817 B.n382 B.n63 163.367
R818 B.n382 B.n381 163.367
R819 B.n381 B.n380 163.367
R820 B.n380 B.n65 163.367
R821 B.n376 B.n65 163.367
R822 B.n376 B.n375 163.367
R823 B.n375 B.n374 163.367
R824 B.n374 B.n67 163.367
R825 B.n370 B.n67 163.367
R826 B.n370 B.n369 163.367
R827 B.n369 B.n368 163.367
R828 B.n368 B.n69 163.367
R829 B.n364 B.n69 163.367
R830 B.n364 B.n363 163.367
R831 B.n363 B.n362 163.367
R832 B.n362 B.n71 163.367
R833 B.n358 B.n71 163.367
R834 B.n358 B.n357 163.367
R835 B.n357 B.n356 163.367
R836 B.n356 B.n73 163.367
R837 B.n352 B.n73 163.367
R838 B.n352 B.n351 163.367
R839 B.n351 B.n350 163.367
R840 B.n350 B.n75 163.367
R841 B.n346 B.n75 163.367
R842 B.n346 B.n345 163.367
R843 B.n345 B.n344 163.367
R844 B.n344 B.n77 163.367
R845 B.n340 B.n77 163.367
R846 B.n340 B.n339 163.367
R847 B.n339 B.n338 163.367
R848 B.n338 B.n79 163.367
R849 B.n334 B.n79 163.367
R850 B.n334 B.n333 163.367
R851 B.n333 B.n332 163.367
R852 B.n332 B.n81 163.367
R853 B.n328 B.n81 163.367
R854 B.n328 B.n327 163.367
R855 B.n327 B.n326 163.367
R856 B.n326 B.n83 163.367
R857 B.n322 B.n83 163.367
R858 B.n322 B.n321 163.367
R859 B.n321 B.n320 163.367
R860 B.n320 B.n85 163.367
R861 B.n316 B.n85 163.367
R862 B.n316 B.n315 163.367
R863 B.n315 B.n314 163.367
R864 B.n314 B.n87 163.367
R865 B.n310 B.n87 163.367
R866 B.n310 B.n309 163.367
R867 B.n309 B.n308 163.367
R868 B.n308 B.n89 163.367
R869 B.n304 B.n89 163.367
R870 B.n304 B.n303 163.367
R871 B.n303 B.n302 163.367
R872 B.n302 B.n91 163.367
R873 B.n298 B.n91 163.367
R874 B.n298 B.n297 163.367
R875 B.n502 B.n501 163.367
R876 B.n501 B.n500 163.367
R877 B.n500 B.n21 163.367
R878 B.n496 B.n21 163.367
R879 B.n496 B.n495 163.367
R880 B.n495 B.n494 163.367
R881 B.n494 B.n23 163.367
R882 B.n490 B.n23 163.367
R883 B.n490 B.n489 163.367
R884 B.n489 B.n488 163.367
R885 B.n488 B.n25 163.367
R886 B.n484 B.n25 163.367
R887 B.n484 B.n483 163.367
R888 B.n483 B.n482 163.367
R889 B.n482 B.n27 163.367
R890 B.n478 B.n27 163.367
R891 B.n478 B.n477 163.367
R892 B.n477 B.n476 163.367
R893 B.n476 B.n29 163.367
R894 B.n472 B.n29 163.367
R895 B.n472 B.n471 163.367
R896 B.n471 B.n470 163.367
R897 B.n470 B.n31 163.367
R898 B.n466 B.n31 163.367
R899 B.n466 B.n465 163.367
R900 B.n465 B.n464 163.367
R901 B.n464 B.n33 163.367
R902 B.n459 B.n33 163.367
R903 B.n459 B.n458 163.367
R904 B.n458 B.n457 163.367
R905 B.n457 B.n37 163.367
R906 B.n453 B.n37 163.367
R907 B.n453 B.n452 163.367
R908 B.n452 B.n451 163.367
R909 B.n451 B.n39 163.367
R910 B.n447 B.n39 163.367
R911 B.n447 B.n446 163.367
R912 B.n446 B.n43 163.367
R913 B.n442 B.n43 163.367
R914 B.n442 B.n441 163.367
R915 B.n441 B.n440 163.367
R916 B.n440 B.n45 163.367
R917 B.n436 B.n45 163.367
R918 B.n436 B.n435 163.367
R919 B.n435 B.n434 163.367
R920 B.n434 B.n47 163.367
R921 B.n430 B.n47 163.367
R922 B.n430 B.n429 163.367
R923 B.n429 B.n428 163.367
R924 B.n428 B.n49 163.367
R925 B.n424 B.n49 163.367
R926 B.n424 B.n423 163.367
R927 B.n423 B.n422 163.367
R928 B.n422 B.n51 163.367
R929 B.n418 B.n51 163.367
R930 B.n418 B.n417 163.367
R931 B.n417 B.n416 163.367
R932 B.n416 B.n53 163.367
R933 B.n412 B.n53 163.367
R934 B.n412 B.n411 163.367
R935 B.n411 B.n410 163.367
R936 B.n410 B.n55 163.367
R937 B.n406 B.n55 163.367
R938 B.n406 B.n405 163.367
R939 B.n506 B.n19 163.367
R940 B.n507 B.n506 163.367
R941 B.n508 B.n507 163.367
R942 B.n508 B.n17 163.367
R943 B.n512 B.n17 163.367
R944 B.n513 B.n512 163.367
R945 B.n514 B.n513 163.367
R946 B.n514 B.n15 163.367
R947 B.n518 B.n15 163.367
R948 B.n519 B.n518 163.367
R949 B.n520 B.n519 163.367
R950 B.n520 B.n13 163.367
R951 B.n524 B.n13 163.367
R952 B.n525 B.n524 163.367
R953 B.n526 B.n525 163.367
R954 B.n526 B.n11 163.367
R955 B.n530 B.n11 163.367
R956 B.n531 B.n530 163.367
R957 B.n532 B.n531 163.367
R958 B.n532 B.n9 163.367
R959 B.n536 B.n9 163.367
R960 B.n537 B.n536 163.367
R961 B.n538 B.n537 163.367
R962 B.n538 B.n7 163.367
R963 B.n542 B.n7 163.367
R964 B.n543 B.n542 163.367
R965 B.n544 B.n543 163.367
R966 B.n544 B.n5 163.367
R967 B.n548 B.n5 163.367
R968 B.n549 B.n548 163.367
R969 B.n550 B.n549 163.367
R970 B.n550 B.n3 163.367
R971 B.n554 B.n3 163.367
R972 B.n555 B.n554 163.367
R973 B.n144 B.n2 163.367
R974 B.n144 B.n143 163.367
R975 B.n148 B.n143 163.367
R976 B.n149 B.n148 163.367
R977 B.n150 B.n149 163.367
R978 B.n150 B.n141 163.367
R979 B.n154 B.n141 163.367
R980 B.n155 B.n154 163.367
R981 B.n156 B.n155 163.367
R982 B.n156 B.n139 163.367
R983 B.n160 B.n139 163.367
R984 B.n161 B.n160 163.367
R985 B.n162 B.n161 163.367
R986 B.n162 B.n137 163.367
R987 B.n166 B.n137 163.367
R988 B.n167 B.n166 163.367
R989 B.n168 B.n167 163.367
R990 B.n168 B.n135 163.367
R991 B.n172 B.n135 163.367
R992 B.n173 B.n172 163.367
R993 B.n174 B.n173 163.367
R994 B.n174 B.n133 163.367
R995 B.n178 B.n133 163.367
R996 B.n179 B.n178 163.367
R997 B.n180 B.n179 163.367
R998 B.n180 B.n131 163.367
R999 B.n184 B.n131 163.367
R1000 B.n185 B.n184 163.367
R1001 B.n186 B.n185 163.367
R1002 B.n186 B.n129 163.367
R1003 B.n190 B.n129 163.367
R1004 B.n191 B.n190 163.367
R1005 B.n192 B.n191 163.367
R1006 B.n192 B.n127 163.367
R1007 B.n237 B.n113 59.5399
R1008 B.n252 B.n251 59.5399
R1009 B.n42 B.n41 59.5399
R1010 B.n461 B.n35 59.5399
R1011 B.n113 B.n112 30.0611
R1012 B.n251 B.n250 30.0611
R1013 B.n41 B.n40 30.0611
R1014 B.n35 B.n34 30.0611
R1015 B.n295 B.n92 29.5029
R1016 B.n504 B.n503 29.5029
R1017 B.n403 B.n56 29.5029
R1018 B.n195 B.n194 29.5029
R1019 B B.n557 18.0485
R1020 B.n505 B.n504 10.6151
R1021 B.n505 B.n18 10.6151
R1022 B.n509 B.n18 10.6151
R1023 B.n510 B.n509 10.6151
R1024 B.n511 B.n510 10.6151
R1025 B.n511 B.n16 10.6151
R1026 B.n515 B.n16 10.6151
R1027 B.n516 B.n515 10.6151
R1028 B.n517 B.n516 10.6151
R1029 B.n517 B.n14 10.6151
R1030 B.n521 B.n14 10.6151
R1031 B.n522 B.n521 10.6151
R1032 B.n523 B.n522 10.6151
R1033 B.n523 B.n12 10.6151
R1034 B.n527 B.n12 10.6151
R1035 B.n528 B.n527 10.6151
R1036 B.n529 B.n528 10.6151
R1037 B.n529 B.n10 10.6151
R1038 B.n533 B.n10 10.6151
R1039 B.n534 B.n533 10.6151
R1040 B.n535 B.n534 10.6151
R1041 B.n535 B.n8 10.6151
R1042 B.n539 B.n8 10.6151
R1043 B.n540 B.n539 10.6151
R1044 B.n541 B.n540 10.6151
R1045 B.n541 B.n6 10.6151
R1046 B.n545 B.n6 10.6151
R1047 B.n546 B.n545 10.6151
R1048 B.n547 B.n546 10.6151
R1049 B.n547 B.n4 10.6151
R1050 B.n551 B.n4 10.6151
R1051 B.n552 B.n551 10.6151
R1052 B.n553 B.n552 10.6151
R1053 B.n553 B.n0 10.6151
R1054 B.n503 B.n20 10.6151
R1055 B.n499 B.n20 10.6151
R1056 B.n499 B.n498 10.6151
R1057 B.n498 B.n497 10.6151
R1058 B.n497 B.n22 10.6151
R1059 B.n493 B.n22 10.6151
R1060 B.n493 B.n492 10.6151
R1061 B.n492 B.n491 10.6151
R1062 B.n491 B.n24 10.6151
R1063 B.n487 B.n24 10.6151
R1064 B.n487 B.n486 10.6151
R1065 B.n486 B.n485 10.6151
R1066 B.n485 B.n26 10.6151
R1067 B.n481 B.n26 10.6151
R1068 B.n481 B.n480 10.6151
R1069 B.n480 B.n479 10.6151
R1070 B.n479 B.n28 10.6151
R1071 B.n475 B.n28 10.6151
R1072 B.n475 B.n474 10.6151
R1073 B.n474 B.n473 10.6151
R1074 B.n473 B.n30 10.6151
R1075 B.n469 B.n30 10.6151
R1076 B.n469 B.n468 10.6151
R1077 B.n468 B.n467 10.6151
R1078 B.n467 B.n32 10.6151
R1079 B.n463 B.n32 10.6151
R1080 B.n463 B.n462 10.6151
R1081 B.n460 B.n36 10.6151
R1082 B.n456 B.n36 10.6151
R1083 B.n456 B.n455 10.6151
R1084 B.n455 B.n454 10.6151
R1085 B.n454 B.n38 10.6151
R1086 B.n450 B.n38 10.6151
R1087 B.n450 B.n449 10.6151
R1088 B.n449 B.n448 10.6151
R1089 B.n445 B.n444 10.6151
R1090 B.n444 B.n443 10.6151
R1091 B.n443 B.n44 10.6151
R1092 B.n439 B.n44 10.6151
R1093 B.n439 B.n438 10.6151
R1094 B.n438 B.n437 10.6151
R1095 B.n437 B.n46 10.6151
R1096 B.n433 B.n46 10.6151
R1097 B.n433 B.n432 10.6151
R1098 B.n432 B.n431 10.6151
R1099 B.n431 B.n48 10.6151
R1100 B.n427 B.n48 10.6151
R1101 B.n427 B.n426 10.6151
R1102 B.n426 B.n425 10.6151
R1103 B.n425 B.n50 10.6151
R1104 B.n421 B.n50 10.6151
R1105 B.n421 B.n420 10.6151
R1106 B.n420 B.n419 10.6151
R1107 B.n419 B.n52 10.6151
R1108 B.n415 B.n52 10.6151
R1109 B.n415 B.n414 10.6151
R1110 B.n414 B.n413 10.6151
R1111 B.n413 B.n54 10.6151
R1112 B.n409 B.n54 10.6151
R1113 B.n409 B.n408 10.6151
R1114 B.n408 B.n407 10.6151
R1115 B.n407 B.n56 10.6151
R1116 B.n403 B.n402 10.6151
R1117 B.n402 B.n401 10.6151
R1118 B.n401 B.n58 10.6151
R1119 B.n397 B.n58 10.6151
R1120 B.n397 B.n396 10.6151
R1121 B.n396 B.n395 10.6151
R1122 B.n395 B.n60 10.6151
R1123 B.n391 B.n60 10.6151
R1124 B.n391 B.n390 10.6151
R1125 B.n390 B.n389 10.6151
R1126 B.n389 B.n62 10.6151
R1127 B.n385 B.n62 10.6151
R1128 B.n385 B.n384 10.6151
R1129 B.n384 B.n383 10.6151
R1130 B.n383 B.n64 10.6151
R1131 B.n379 B.n64 10.6151
R1132 B.n379 B.n378 10.6151
R1133 B.n378 B.n377 10.6151
R1134 B.n377 B.n66 10.6151
R1135 B.n373 B.n66 10.6151
R1136 B.n373 B.n372 10.6151
R1137 B.n372 B.n371 10.6151
R1138 B.n371 B.n68 10.6151
R1139 B.n367 B.n68 10.6151
R1140 B.n367 B.n366 10.6151
R1141 B.n366 B.n365 10.6151
R1142 B.n365 B.n70 10.6151
R1143 B.n361 B.n70 10.6151
R1144 B.n361 B.n360 10.6151
R1145 B.n360 B.n359 10.6151
R1146 B.n359 B.n72 10.6151
R1147 B.n355 B.n72 10.6151
R1148 B.n355 B.n354 10.6151
R1149 B.n354 B.n353 10.6151
R1150 B.n353 B.n74 10.6151
R1151 B.n349 B.n74 10.6151
R1152 B.n349 B.n348 10.6151
R1153 B.n348 B.n347 10.6151
R1154 B.n347 B.n76 10.6151
R1155 B.n343 B.n76 10.6151
R1156 B.n343 B.n342 10.6151
R1157 B.n342 B.n341 10.6151
R1158 B.n341 B.n78 10.6151
R1159 B.n337 B.n78 10.6151
R1160 B.n337 B.n336 10.6151
R1161 B.n336 B.n335 10.6151
R1162 B.n335 B.n80 10.6151
R1163 B.n331 B.n80 10.6151
R1164 B.n331 B.n330 10.6151
R1165 B.n330 B.n329 10.6151
R1166 B.n329 B.n82 10.6151
R1167 B.n325 B.n82 10.6151
R1168 B.n325 B.n324 10.6151
R1169 B.n324 B.n323 10.6151
R1170 B.n323 B.n84 10.6151
R1171 B.n319 B.n84 10.6151
R1172 B.n319 B.n318 10.6151
R1173 B.n318 B.n317 10.6151
R1174 B.n317 B.n86 10.6151
R1175 B.n313 B.n86 10.6151
R1176 B.n313 B.n312 10.6151
R1177 B.n312 B.n311 10.6151
R1178 B.n311 B.n88 10.6151
R1179 B.n307 B.n88 10.6151
R1180 B.n307 B.n306 10.6151
R1181 B.n306 B.n305 10.6151
R1182 B.n305 B.n90 10.6151
R1183 B.n301 B.n90 10.6151
R1184 B.n301 B.n300 10.6151
R1185 B.n300 B.n299 10.6151
R1186 B.n299 B.n92 10.6151
R1187 B.n145 B.n1 10.6151
R1188 B.n146 B.n145 10.6151
R1189 B.n147 B.n146 10.6151
R1190 B.n147 B.n142 10.6151
R1191 B.n151 B.n142 10.6151
R1192 B.n152 B.n151 10.6151
R1193 B.n153 B.n152 10.6151
R1194 B.n153 B.n140 10.6151
R1195 B.n157 B.n140 10.6151
R1196 B.n158 B.n157 10.6151
R1197 B.n159 B.n158 10.6151
R1198 B.n159 B.n138 10.6151
R1199 B.n163 B.n138 10.6151
R1200 B.n164 B.n163 10.6151
R1201 B.n165 B.n164 10.6151
R1202 B.n165 B.n136 10.6151
R1203 B.n169 B.n136 10.6151
R1204 B.n170 B.n169 10.6151
R1205 B.n171 B.n170 10.6151
R1206 B.n171 B.n134 10.6151
R1207 B.n175 B.n134 10.6151
R1208 B.n176 B.n175 10.6151
R1209 B.n177 B.n176 10.6151
R1210 B.n177 B.n132 10.6151
R1211 B.n181 B.n132 10.6151
R1212 B.n182 B.n181 10.6151
R1213 B.n183 B.n182 10.6151
R1214 B.n183 B.n130 10.6151
R1215 B.n187 B.n130 10.6151
R1216 B.n188 B.n187 10.6151
R1217 B.n189 B.n188 10.6151
R1218 B.n189 B.n128 10.6151
R1219 B.n193 B.n128 10.6151
R1220 B.n194 B.n193 10.6151
R1221 B.n195 B.n126 10.6151
R1222 B.n199 B.n126 10.6151
R1223 B.n200 B.n199 10.6151
R1224 B.n201 B.n200 10.6151
R1225 B.n201 B.n124 10.6151
R1226 B.n205 B.n124 10.6151
R1227 B.n206 B.n205 10.6151
R1228 B.n207 B.n206 10.6151
R1229 B.n207 B.n122 10.6151
R1230 B.n211 B.n122 10.6151
R1231 B.n212 B.n211 10.6151
R1232 B.n213 B.n212 10.6151
R1233 B.n213 B.n120 10.6151
R1234 B.n217 B.n120 10.6151
R1235 B.n218 B.n217 10.6151
R1236 B.n219 B.n218 10.6151
R1237 B.n219 B.n118 10.6151
R1238 B.n223 B.n118 10.6151
R1239 B.n224 B.n223 10.6151
R1240 B.n225 B.n224 10.6151
R1241 B.n225 B.n116 10.6151
R1242 B.n229 B.n116 10.6151
R1243 B.n230 B.n229 10.6151
R1244 B.n231 B.n230 10.6151
R1245 B.n231 B.n114 10.6151
R1246 B.n235 B.n114 10.6151
R1247 B.n236 B.n235 10.6151
R1248 B.n238 B.n110 10.6151
R1249 B.n242 B.n110 10.6151
R1250 B.n243 B.n242 10.6151
R1251 B.n244 B.n243 10.6151
R1252 B.n244 B.n108 10.6151
R1253 B.n248 B.n108 10.6151
R1254 B.n249 B.n248 10.6151
R1255 B.n253 B.n249 10.6151
R1256 B.n257 B.n106 10.6151
R1257 B.n258 B.n257 10.6151
R1258 B.n259 B.n258 10.6151
R1259 B.n259 B.n104 10.6151
R1260 B.n263 B.n104 10.6151
R1261 B.n264 B.n263 10.6151
R1262 B.n265 B.n264 10.6151
R1263 B.n265 B.n102 10.6151
R1264 B.n269 B.n102 10.6151
R1265 B.n270 B.n269 10.6151
R1266 B.n271 B.n270 10.6151
R1267 B.n271 B.n100 10.6151
R1268 B.n275 B.n100 10.6151
R1269 B.n276 B.n275 10.6151
R1270 B.n277 B.n276 10.6151
R1271 B.n277 B.n98 10.6151
R1272 B.n281 B.n98 10.6151
R1273 B.n282 B.n281 10.6151
R1274 B.n283 B.n282 10.6151
R1275 B.n283 B.n96 10.6151
R1276 B.n287 B.n96 10.6151
R1277 B.n288 B.n287 10.6151
R1278 B.n289 B.n288 10.6151
R1279 B.n289 B.n94 10.6151
R1280 B.n293 B.n94 10.6151
R1281 B.n294 B.n293 10.6151
R1282 B.n295 B.n294 10.6151
R1283 B.n557 B.n0 8.11757
R1284 B.n557 B.n1 8.11757
R1285 B.n461 B.n460 6.5566
R1286 B.n448 B.n42 6.5566
R1287 B.n238 B.n237 6.5566
R1288 B.n253 B.n252 6.5566
R1289 B.n462 B.n461 4.05904
R1290 B.n445 B.n42 4.05904
R1291 B.n237 B.n236 4.05904
R1292 B.n252 B.n106 4.05904
R1293 VP.n13 VP.t5 194.32
R1294 VP.n30 VP.t4 174.429
R1295 VP.n47 VP.t7 174.429
R1296 VP.n27 VP.t9 174.429
R1297 VP.n15 VP.n14 161.3
R1298 VP.n16 VP.n11 161.3
R1299 VP.n18 VP.n17 161.3
R1300 VP.n20 VP.n19 161.3
R1301 VP.n21 VP.n9 161.3
R1302 VP.n23 VP.n22 161.3
R1303 VP.n25 VP.n24 161.3
R1304 VP.n26 VP.n7 161.3
R1305 VP.n46 VP.n0 161.3
R1306 VP.n45 VP.n44 161.3
R1307 VP.n43 VP.n42 161.3
R1308 VP.n41 VP.n2 161.3
R1309 VP.n40 VP.n39 161.3
R1310 VP.n38 VP.n37 161.3
R1311 VP.n36 VP.n4 161.3
R1312 VP.n35 VP.n34 161.3
R1313 VP.n33 VP.n32 161.3
R1314 VP.n31 VP.n6 161.3
R1315 VP.n5 VP.t8 142.032
R1316 VP.n3 VP.t6 142.032
R1317 VP.n1 VP.t0 142.032
R1318 VP.n8 VP.t1 142.032
R1319 VP.n10 VP.t3 142.032
R1320 VP.n12 VP.t2 142.032
R1321 VP.n28 VP.n27 80.6037
R1322 VP.n48 VP.n47 80.6037
R1323 VP.n30 VP.n29 80.6037
R1324 VP.n36 VP.n35 42.9216
R1325 VP.n42 VP.n41 42.9216
R1326 VP.n22 VP.n21 42.9216
R1327 VP.n16 VP.n15 42.9216
R1328 VP.n13 VP.n12 42.7694
R1329 VP.n29 VP.n28 42.1264
R1330 VP.n37 VP.n36 38.0652
R1331 VP.n41 VP.n40 38.0652
R1332 VP.n21 VP.n20 38.0652
R1333 VP.n17 VP.n16 38.0652
R1334 VP.n31 VP.n30 35.055
R1335 VP.n47 VP.n46 35.055
R1336 VP.n27 VP.n26 35.055
R1337 VP.n32 VP.n31 33.2089
R1338 VP.n46 VP.n45 33.2089
R1339 VP.n26 VP.n25 33.2089
R1340 VP.n14 VP.n13 29.263
R1341 VP.n35 VP.n5 14.6807
R1342 VP.n42 VP.n1 14.6807
R1343 VP.n22 VP.n8 14.6807
R1344 VP.n15 VP.n12 14.6807
R1345 VP.n37 VP.n3 12.234
R1346 VP.n40 VP.n3 12.234
R1347 VP.n17 VP.n10 12.234
R1348 VP.n20 VP.n10 12.234
R1349 VP.n32 VP.n5 9.7873
R1350 VP.n45 VP.n1 9.7873
R1351 VP.n25 VP.n8 9.7873
R1352 VP.n28 VP.n7 0.285035
R1353 VP.n29 VP.n6 0.285035
R1354 VP.n48 VP.n0 0.285035
R1355 VP.n14 VP.n11 0.189894
R1356 VP.n18 VP.n11 0.189894
R1357 VP.n19 VP.n18 0.189894
R1358 VP.n19 VP.n9 0.189894
R1359 VP.n23 VP.n9 0.189894
R1360 VP.n24 VP.n23 0.189894
R1361 VP.n24 VP.n7 0.189894
R1362 VP.n33 VP.n6 0.189894
R1363 VP.n34 VP.n33 0.189894
R1364 VP.n34 VP.n4 0.189894
R1365 VP.n38 VP.n4 0.189894
R1366 VP.n39 VP.n38 0.189894
R1367 VP.n39 VP.n2 0.189894
R1368 VP.n43 VP.n2 0.189894
R1369 VP.n44 VP.n43 0.189894
R1370 VP.n44 VP.n0 0.189894
R1371 VP VP.n48 0.146778
R1372 VDD1.n31 VDD1.n30 585
R1373 VDD1.n29 VDD1.n28 585
R1374 VDD1.n4 VDD1.n3 585
R1375 VDD1.n23 VDD1.n22 585
R1376 VDD1.n21 VDD1.n20 585
R1377 VDD1.n8 VDD1.n7 585
R1378 VDD1.n15 VDD1.n14 585
R1379 VDD1.n13 VDD1.n12 585
R1380 VDD1.n50 VDD1.n49 585
R1381 VDD1.n52 VDD1.n51 585
R1382 VDD1.n45 VDD1.n44 585
R1383 VDD1.n58 VDD1.n57 585
R1384 VDD1.n60 VDD1.n59 585
R1385 VDD1.n41 VDD1.n40 585
R1386 VDD1.n66 VDD1.n65 585
R1387 VDD1.n68 VDD1.n67 585
R1388 VDD1.n30 VDD1.n0 498.474
R1389 VDD1.n67 VDD1.n37 498.474
R1390 VDD1.n11 VDD1.t4 329.053
R1391 VDD1.n48 VDD1.t5 329.053
R1392 VDD1.n30 VDD1.n29 171.744
R1393 VDD1.n29 VDD1.n3 171.744
R1394 VDD1.n22 VDD1.n3 171.744
R1395 VDD1.n22 VDD1.n21 171.744
R1396 VDD1.n21 VDD1.n7 171.744
R1397 VDD1.n14 VDD1.n7 171.744
R1398 VDD1.n14 VDD1.n13 171.744
R1399 VDD1.n51 VDD1.n50 171.744
R1400 VDD1.n51 VDD1.n44 171.744
R1401 VDD1.n58 VDD1.n44 171.744
R1402 VDD1.n59 VDD1.n58 171.744
R1403 VDD1.n59 VDD1.n40 171.744
R1404 VDD1.n66 VDD1.n40 171.744
R1405 VDD1.n67 VDD1.n66 171.744
R1406 VDD1.n75 VDD1.n74 87.9189
R1407 VDD1.n36 VDD1.n35 86.9722
R1408 VDD1.n77 VDD1.n76 86.972
R1409 VDD1.n73 VDD1.n72 86.972
R1410 VDD1.n13 VDD1.t4 85.8723
R1411 VDD1.n50 VDD1.t5 85.8723
R1412 VDD1.n36 VDD1.n34 52.3337
R1413 VDD1.n73 VDD1.n71 52.3337
R1414 VDD1.n77 VDD1.n75 37.5117
R1415 VDD1.n32 VDD1.n31 12.8005
R1416 VDD1.n69 VDD1.n68 12.8005
R1417 VDD1.n28 VDD1.n2 12.0247
R1418 VDD1.n65 VDD1.n39 12.0247
R1419 VDD1.n27 VDD1.n4 11.249
R1420 VDD1.n64 VDD1.n41 11.249
R1421 VDD1.n12 VDD1.n11 10.7237
R1422 VDD1.n49 VDD1.n48 10.7237
R1423 VDD1.n24 VDD1.n23 10.4732
R1424 VDD1.n61 VDD1.n60 10.4732
R1425 VDD1.n20 VDD1.n6 9.69747
R1426 VDD1.n57 VDD1.n43 9.69747
R1427 VDD1.n34 VDD1.n33 9.45567
R1428 VDD1.n71 VDD1.n70 9.45567
R1429 VDD1.n10 VDD1.n9 9.3005
R1430 VDD1.n17 VDD1.n16 9.3005
R1431 VDD1.n19 VDD1.n18 9.3005
R1432 VDD1.n6 VDD1.n5 9.3005
R1433 VDD1.n25 VDD1.n24 9.3005
R1434 VDD1.n27 VDD1.n26 9.3005
R1435 VDD1.n2 VDD1.n1 9.3005
R1436 VDD1.n33 VDD1.n32 9.3005
R1437 VDD1.n47 VDD1.n46 9.3005
R1438 VDD1.n54 VDD1.n53 9.3005
R1439 VDD1.n56 VDD1.n55 9.3005
R1440 VDD1.n43 VDD1.n42 9.3005
R1441 VDD1.n62 VDD1.n61 9.3005
R1442 VDD1.n64 VDD1.n63 9.3005
R1443 VDD1.n39 VDD1.n38 9.3005
R1444 VDD1.n70 VDD1.n69 9.3005
R1445 VDD1.n19 VDD1.n8 8.92171
R1446 VDD1.n56 VDD1.n45 8.92171
R1447 VDD1.n16 VDD1.n15 8.14595
R1448 VDD1.n53 VDD1.n52 8.14595
R1449 VDD1.n34 VDD1.n0 7.75445
R1450 VDD1.n71 VDD1.n37 7.75445
R1451 VDD1.n12 VDD1.n10 7.3702
R1452 VDD1.n49 VDD1.n47 7.3702
R1453 VDD1.n32 VDD1.n0 6.08283
R1454 VDD1.n69 VDD1.n37 6.08283
R1455 VDD1.n15 VDD1.n10 5.81868
R1456 VDD1.n52 VDD1.n47 5.81868
R1457 VDD1.n16 VDD1.n8 5.04292
R1458 VDD1.n53 VDD1.n45 5.04292
R1459 VDD1.n76 VDD1.t8 4.52136
R1460 VDD1.n76 VDD1.t0 4.52136
R1461 VDD1.n35 VDD1.t7 4.52136
R1462 VDD1.n35 VDD1.t6 4.52136
R1463 VDD1.n74 VDD1.t9 4.52136
R1464 VDD1.n74 VDD1.t2 4.52136
R1465 VDD1.n72 VDD1.t1 4.52136
R1466 VDD1.n72 VDD1.t3 4.52136
R1467 VDD1.n20 VDD1.n19 4.26717
R1468 VDD1.n57 VDD1.n56 4.26717
R1469 VDD1.n23 VDD1.n6 3.49141
R1470 VDD1.n60 VDD1.n43 3.49141
R1471 VDD1.n24 VDD1.n4 2.71565
R1472 VDD1.n61 VDD1.n41 2.71565
R1473 VDD1.n11 VDD1.n9 2.41305
R1474 VDD1.n48 VDD1.n46 2.41305
R1475 VDD1.n28 VDD1.n27 1.93989
R1476 VDD1.n65 VDD1.n64 1.93989
R1477 VDD1.n31 VDD1.n2 1.16414
R1478 VDD1.n68 VDD1.n39 1.16414
R1479 VDD1 VDD1.n77 0.944465
R1480 VDD1 VDD1.n36 0.392741
R1481 VDD1.n75 VDD1.n73 0.279206
R1482 VDD1.n33 VDD1.n1 0.155672
R1483 VDD1.n26 VDD1.n1 0.155672
R1484 VDD1.n26 VDD1.n25 0.155672
R1485 VDD1.n25 VDD1.n5 0.155672
R1486 VDD1.n18 VDD1.n5 0.155672
R1487 VDD1.n18 VDD1.n17 0.155672
R1488 VDD1.n17 VDD1.n9 0.155672
R1489 VDD1.n54 VDD1.n46 0.155672
R1490 VDD1.n55 VDD1.n54 0.155672
R1491 VDD1.n55 VDD1.n42 0.155672
R1492 VDD1.n62 VDD1.n42 0.155672
R1493 VDD1.n63 VDD1.n62 0.155672
R1494 VDD1.n63 VDD1.n38 0.155672
R1495 VDD1.n70 VDD1.n38 0.155672
C0 VP w_n2830_n2406# 5.91199f
C1 VN w_n2830_n2406# 5.54779f
C2 VDD1 w_n2830_n2406# 1.90699f
C3 VDD2 w_n2830_n2406# 1.97883f
C4 B VTAIL 2.12063f
C5 B VP 1.48024f
C6 VTAIL VP 5.72292f
C7 VN B 0.87544f
C8 VDD1 B 1.5636f
C9 VN VTAIL 5.7086f
C10 VDD1 VTAIL 8.16852f
C11 VN VP 5.47263f
C12 VDD1 VP 5.60383f
C13 VDD2 B 1.62782f
C14 VDD2 VTAIL 8.209901f
C15 VN VDD1 0.149917f
C16 VDD2 VP 0.40683f
C17 B w_n2830_n2406# 6.87827f
C18 VN VDD2 5.34981f
C19 VTAIL w_n2830_n2406# 2.3257f
C20 VDD2 VDD1 1.28987f
C21 VDD2 VSUBS 1.305503f
C22 VDD1 VSUBS 1.21151f
C23 VTAIL VSUBS 0.554923f
C24 VN VSUBS 5.23218f
C25 VP VSUBS 2.199607f
C26 B VSUBS 3.247451f
C27 w_n2830_n2406# VSUBS 84.6623f
C28 VDD1.n0 VSUBS 0.024582f
C29 VDD1.n1 VSUBS 0.023289f
C30 VDD1.n2 VSUBS 0.012514f
C31 VDD1.n3 VSUBS 0.029579f
C32 VDD1.n4 VSUBS 0.01325f
C33 VDD1.n5 VSUBS 0.023289f
C34 VDD1.n6 VSUBS 0.012514f
C35 VDD1.n7 VSUBS 0.029579f
C36 VDD1.n8 VSUBS 0.01325f
C37 VDD1.n9 VSUBS 0.653135f
C38 VDD1.n10 VSUBS 0.012514f
C39 VDD1.t4 VSUBS 0.063519f
C40 VDD1.n11 VSUBS 0.132891f
C41 VDD1.n12 VSUBS 0.02225f
C42 VDD1.n13 VSUBS 0.022184f
C43 VDD1.n14 VSUBS 0.029579f
C44 VDD1.n15 VSUBS 0.01325f
C45 VDD1.n16 VSUBS 0.012514f
C46 VDD1.n17 VSUBS 0.023289f
C47 VDD1.n18 VSUBS 0.023289f
C48 VDD1.n19 VSUBS 0.012514f
C49 VDD1.n20 VSUBS 0.01325f
C50 VDD1.n21 VSUBS 0.029579f
C51 VDD1.n22 VSUBS 0.029579f
C52 VDD1.n23 VSUBS 0.01325f
C53 VDD1.n24 VSUBS 0.012514f
C54 VDD1.n25 VSUBS 0.023289f
C55 VDD1.n26 VSUBS 0.023289f
C56 VDD1.n27 VSUBS 0.012514f
C57 VDD1.n28 VSUBS 0.01325f
C58 VDD1.n29 VSUBS 0.029579f
C59 VDD1.n30 VSUBS 0.072551f
C60 VDD1.n31 VSUBS 0.01325f
C61 VDD1.n32 VSUBS 0.024575f
C62 VDD1.n33 VSUBS 0.05733f
C63 VDD1.n34 VSUBS 0.074889f
C64 VDD1.t7 VSUBS 0.13232f
C65 VDD1.t6 VSUBS 0.13232f
C66 VDD1.n35 VSUBS 0.935353f
C67 VDD1.n36 VSUBS 0.656017f
C68 VDD1.n37 VSUBS 0.024582f
C69 VDD1.n38 VSUBS 0.023289f
C70 VDD1.n39 VSUBS 0.012514f
C71 VDD1.n40 VSUBS 0.029579f
C72 VDD1.n41 VSUBS 0.01325f
C73 VDD1.n42 VSUBS 0.023289f
C74 VDD1.n43 VSUBS 0.012514f
C75 VDD1.n44 VSUBS 0.029579f
C76 VDD1.n45 VSUBS 0.01325f
C77 VDD1.n46 VSUBS 0.653135f
C78 VDD1.n47 VSUBS 0.012514f
C79 VDD1.t5 VSUBS 0.063519f
C80 VDD1.n48 VSUBS 0.132891f
C81 VDD1.n49 VSUBS 0.02225f
C82 VDD1.n50 VSUBS 0.022184f
C83 VDD1.n51 VSUBS 0.029579f
C84 VDD1.n52 VSUBS 0.01325f
C85 VDD1.n53 VSUBS 0.012514f
C86 VDD1.n54 VSUBS 0.023289f
C87 VDD1.n55 VSUBS 0.023289f
C88 VDD1.n56 VSUBS 0.012514f
C89 VDD1.n57 VSUBS 0.01325f
C90 VDD1.n58 VSUBS 0.029579f
C91 VDD1.n59 VSUBS 0.029579f
C92 VDD1.n60 VSUBS 0.01325f
C93 VDD1.n61 VSUBS 0.012514f
C94 VDD1.n62 VSUBS 0.023289f
C95 VDD1.n63 VSUBS 0.023289f
C96 VDD1.n64 VSUBS 0.012514f
C97 VDD1.n65 VSUBS 0.01325f
C98 VDD1.n66 VSUBS 0.029579f
C99 VDD1.n67 VSUBS 0.072551f
C100 VDD1.n68 VSUBS 0.01325f
C101 VDD1.n69 VSUBS 0.024575f
C102 VDD1.n70 VSUBS 0.05733f
C103 VDD1.n71 VSUBS 0.074889f
C104 VDD1.t1 VSUBS 0.13232f
C105 VDD1.t3 VSUBS 0.13232f
C106 VDD1.n72 VSUBS 0.935348f
C107 VDD1.n73 VSUBS 0.64944f
C108 VDD1.t9 VSUBS 0.13232f
C109 VDD1.t2 VSUBS 0.13232f
C110 VDD1.n74 VSUBS 0.941424f
C111 VDD1.n75 VSUBS 2.03271f
C112 VDD1.t8 VSUBS 0.13232f
C113 VDD1.t0 VSUBS 0.13232f
C114 VDD1.n76 VSUBS 0.935348f
C115 VDD1.n77 VSUBS 2.26459f
C116 VP.n0 VSUBS 0.063781f
C117 VP.t0 VSUBS 1.12055f
C118 VP.n1 VSUBS 0.435656f
C119 VP.n2 VSUBS 0.047799f
C120 VP.t6 VSUBS 1.12055f
C121 VP.n3 VSUBS 0.435656f
C122 VP.n4 VSUBS 0.047799f
C123 VP.t8 VSUBS 1.12055f
C124 VP.n5 VSUBS 0.435656f
C125 VP.n6 VSUBS 0.063781f
C126 VP.n7 VSUBS 0.063781f
C127 VP.t9 VSUBS 1.20989f
C128 VP.t1 VSUBS 1.12055f
C129 VP.n8 VSUBS 0.435656f
C130 VP.n9 VSUBS 0.047799f
C131 VP.t3 VSUBS 1.12055f
C132 VP.n10 VSUBS 0.435656f
C133 VP.n11 VSUBS 0.047799f
C134 VP.t2 VSUBS 1.12055f
C135 VP.n12 VSUBS 0.499765f
C136 VP.t5 VSUBS 1.26487f
C137 VP.n13 VSUBS 0.513786f
C138 VP.n14 VSUBS 0.249114f
C139 VP.n15 VSUBS 0.076031f
C140 VP.n16 VSUBS 0.039028f
C141 VP.n17 VSUBS 0.074007f
C142 VP.n18 VSUBS 0.047799f
C143 VP.n19 VSUBS 0.047799f
C144 VP.n20 VSUBS 0.074007f
C145 VP.n21 VSUBS 0.039028f
C146 VP.n22 VSUBS 0.076031f
C147 VP.n23 VSUBS 0.047799f
C148 VP.n24 VSUBS 0.047799f
C149 VP.n25 VSUBS 0.070105f
C150 VP.n26 VSUBS 0.034238f
C151 VP.n27 VSUBS 0.526282f
C152 VP.n28 VSUBS 1.99989f
C153 VP.n29 VSUBS 2.04068f
C154 VP.t4 VSUBS 1.20989f
C155 VP.n30 VSUBS 0.526282f
C156 VP.n31 VSUBS 0.034238f
C157 VP.n32 VSUBS 0.070105f
C158 VP.n33 VSUBS 0.047799f
C159 VP.n34 VSUBS 0.047799f
C160 VP.n35 VSUBS 0.076031f
C161 VP.n36 VSUBS 0.039028f
C162 VP.n37 VSUBS 0.074007f
C163 VP.n38 VSUBS 0.047799f
C164 VP.n39 VSUBS 0.047799f
C165 VP.n40 VSUBS 0.074007f
C166 VP.n41 VSUBS 0.039028f
C167 VP.n42 VSUBS 0.076031f
C168 VP.n43 VSUBS 0.047799f
C169 VP.n44 VSUBS 0.047799f
C170 VP.n45 VSUBS 0.070105f
C171 VP.n46 VSUBS 0.034238f
C172 VP.t7 VSUBS 1.20989f
C173 VP.n47 VSUBS 0.526282f
C174 VP.n48 VSUBS 0.044765f
C175 B.n0 VSUBS 0.006868f
C176 B.n1 VSUBS 0.006868f
C177 B.n2 VSUBS 0.010157f
C178 B.n3 VSUBS 0.007784f
C179 B.n4 VSUBS 0.007784f
C180 B.n5 VSUBS 0.007784f
C181 B.n6 VSUBS 0.007784f
C182 B.n7 VSUBS 0.007784f
C183 B.n8 VSUBS 0.007784f
C184 B.n9 VSUBS 0.007784f
C185 B.n10 VSUBS 0.007784f
C186 B.n11 VSUBS 0.007784f
C187 B.n12 VSUBS 0.007784f
C188 B.n13 VSUBS 0.007784f
C189 B.n14 VSUBS 0.007784f
C190 B.n15 VSUBS 0.007784f
C191 B.n16 VSUBS 0.007784f
C192 B.n17 VSUBS 0.007784f
C193 B.n18 VSUBS 0.007784f
C194 B.n19 VSUBS 0.016397f
C195 B.n20 VSUBS 0.007784f
C196 B.n21 VSUBS 0.007784f
C197 B.n22 VSUBS 0.007784f
C198 B.n23 VSUBS 0.007784f
C199 B.n24 VSUBS 0.007784f
C200 B.n25 VSUBS 0.007784f
C201 B.n26 VSUBS 0.007784f
C202 B.n27 VSUBS 0.007784f
C203 B.n28 VSUBS 0.007784f
C204 B.n29 VSUBS 0.007784f
C205 B.n30 VSUBS 0.007784f
C206 B.n31 VSUBS 0.007784f
C207 B.n32 VSUBS 0.007784f
C208 B.n33 VSUBS 0.007784f
C209 B.t1 VSUBS 0.123207f
C210 B.t2 VSUBS 0.140226f
C211 B.t0 VSUBS 0.4351f
C212 B.n34 VSUBS 0.238661f
C213 B.n35 VSUBS 0.191735f
C214 B.n36 VSUBS 0.007784f
C215 B.n37 VSUBS 0.007784f
C216 B.n38 VSUBS 0.007784f
C217 B.n39 VSUBS 0.007784f
C218 B.t7 VSUBS 0.12321f
C219 B.t8 VSUBS 0.140228f
C220 B.t6 VSUBS 0.4351f
C221 B.n40 VSUBS 0.238659f
C222 B.n41 VSUBS 0.191733f
C223 B.n42 VSUBS 0.018034f
C224 B.n43 VSUBS 0.007784f
C225 B.n44 VSUBS 0.007784f
C226 B.n45 VSUBS 0.007784f
C227 B.n46 VSUBS 0.007784f
C228 B.n47 VSUBS 0.007784f
C229 B.n48 VSUBS 0.007784f
C230 B.n49 VSUBS 0.007784f
C231 B.n50 VSUBS 0.007784f
C232 B.n51 VSUBS 0.007784f
C233 B.n52 VSUBS 0.007784f
C234 B.n53 VSUBS 0.007784f
C235 B.n54 VSUBS 0.007784f
C236 B.n55 VSUBS 0.007784f
C237 B.n56 VSUBS 0.017713f
C238 B.n57 VSUBS 0.007784f
C239 B.n58 VSUBS 0.007784f
C240 B.n59 VSUBS 0.007784f
C241 B.n60 VSUBS 0.007784f
C242 B.n61 VSUBS 0.007784f
C243 B.n62 VSUBS 0.007784f
C244 B.n63 VSUBS 0.007784f
C245 B.n64 VSUBS 0.007784f
C246 B.n65 VSUBS 0.007784f
C247 B.n66 VSUBS 0.007784f
C248 B.n67 VSUBS 0.007784f
C249 B.n68 VSUBS 0.007784f
C250 B.n69 VSUBS 0.007784f
C251 B.n70 VSUBS 0.007784f
C252 B.n71 VSUBS 0.007784f
C253 B.n72 VSUBS 0.007784f
C254 B.n73 VSUBS 0.007784f
C255 B.n74 VSUBS 0.007784f
C256 B.n75 VSUBS 0.007784f
C257 B.n76 VSUBS 0.007784f
C258 B.n77 VSUBS 0.007784f
C259 B.n78 VSUBS 0.007784f
C260 B.n79 VSUBS 0.007784f
C261 B.n80 VSUBS 0.007784f
C262 B.n81 VSUBS 0.007784f
C263 B.n82 VSUBS 0.007784f
C264 B.n83 VSUBS 0.007784f
C265 B.n84 VSUBS 0.007784f
C266 B.n85 VSUBS 0.007784f
C267 B.n86 VSUBS 0.007784f
C268 B.n87 VSUBS 0.007784f
C269 B.n88 VSUBS 0.007784f
C270 B.n89 VSUBS 0.007784f
C271 B.n90 VSUBS 0.007784f
C272 B.n91 VSUBS 0.007784f
C273 B.n92 VSUBS 0.017415f
C274 B.n93 VSUBS 0.007784f
C275 B.n94 VSUBS 0.007784f
C276 B.n95 VSUBS 0.007784f
C277 B.n96 VSUBS 0.007784f
C278 B.n97 VSUBS 0.007784f
C279 B.n98 VSUBS 0.007784f
C280 B.n99 VSUBS 0.007784f
C281 B.n100 VSUBS 0.007784f
C282 B.n101 VSUBS 0.007784f
C283 B.n102 VSUBS 0.007784f
C284 B.n103 VSUBS 0.007784f
C285 B.n104 VSUBS 0.007784f
C286 B.n105 VSUBS 0.007784f
C287 B.n106 VSUBS 0.00538f
C288 B.n107 VSUBS 0.007784f
C289 B.n108 VSUBS 0.007784f
C290 B.n109 VSUBS 0.007784f
C291 B.n110 VSUBS 0.007784f
C292 B.n111 VSUBS 0.007784f
C293 B.t5 VSUBS 0.123207f
C294 B.t4 VSUBS 0.140226f
C295 B.t3 VSUBS 0.4351f
C296 B.n112 VSUBS 0.238661f
C297 B.n113 VSUBS 0.191735f
C298 B.n114 VSUBS 0.007784f
C299 B.n115 VSUBS 0.007784f
C300 B.n116 VSUBS 0.007784f
C301 B.n117 VSUBS 0.007784f
C302 B.n118 VSUBS 0.007784f
C303 B.n119 VSUBS 0.007784f
C304 B.n120 VSUBS 0.007784f
C305 B.n121 VSUBS 0.007784f
C306 B.n122 VSUBS 0.007784f
C307 B.n123 VSUBS 0.007784f
C308 B.n124 VSUBS 0.007784f
C309 B.n125 VSUBS 0.007784f
C310 B.n126 VSUBS 0.007784f
C311 B.n127 VSUBS 0.016397f
C312 B.n128 VSUBS 0.007784f
C313 B.n129 VSUBS 0.007784f
C314 B.n130 VSUBS 0.007784f
C315 B.n131 VSUBS 0.007784f
C316 B.n132 VSUBS 0.007784f
C317 B.n133 VSUBS 0.007784f
C318 B.n134 VSUBS 0.007784f
C319 B.n135 VSUBS 0.007784f
C320 B.n136 VSUBS 0.007784f
C321 B.n137 VSUBS 0.007784f
C322 B.n138 VSUBS 0.007784f
C323 B.n139 VSUBS 0.007784f
C324 B.n140 VSUBS 0.007784f
C325 B.n141 VSUBS 0.007784f
C326 B.n142 VSUBS 0.007784f
C327 B.n143 VSUBS 0.007784f
C328 B.n144 VSUBS 0.007784f
C329 B.n145 VSUBS 0.007784f
C330 B.n146 VSUBS 0.007784f
C331 B.n147 VSUBS 0.007784f
C332 B.n148 VSUBS 0.007784f
C333 B.n149 VSUBS 0.007784f
C334 B.n150 VSUBS 0.007784f
C335 B.n151 VSUBS 0.007784f
C336 B.n152 VSUBS 0.007784f
C337 B.n153 VSUBS 0.007784f
C338 B.n154 VSUBS 0.007784f
C339 B.n155 VSUBS 0.007784f
C340 B.n156 VSUBS 0.007784f
C341 B.n157 VSUBS 0.007784f
C342 B.n158 VSUBS 0.007784f
C343 B.n159 VSUBS 0.007784f
C344 B.n160 VSUBS 0.007784f
C345 B.n161 VSUBS 0.007784f
C346 B.n162 VSUBS 0.007784f
C347 B.n163 VSUBS 0.007784f
C348 B.n164 VSUBS 0.007784f
C349 B.n165 VSUBS 0.007784f
C350 B.n166 VSUBS 0.007784f
C351 B.n167 VSUBS 0.007784f
C352 B.n168 VSUBS 0.007784f
C353 B.n169 VSUBS 0.007784f
C354 B.n170 VSUBS 0.007784f
C355 B.n171 VSUBS 0.007784f
C356 B.n172 VSUBS 0.007784f
C357 B.n173 VSUBS 0.007784f
C358 B.n174 VSUBS 0.007784f
C359 B.n175 VSUBS 0.007784f
C360 B.n176 VSUBS 0.007784f
C361 B.n177 VSUBS 0.007784f
C362 B.n178 VSUBS 0.007784f
C363 B.n179 VSUBS 0.007784f
C364 B.n180 VSUBS 0.007784f
C365 B.n181 VSUBS 0.007784f
C366 B.n182 VSUBS 0.007784f
C367 B.n183 VSUBS 0.007784f
C368 B.n184 VSUBS 0.007784f
C369 B.n185 VSUBS 0.007784f
C370 B.n186 VSUBS 0.007784f
C371 B.n187 VSUBS 0.007784f
C372 B.n188 VSUBS 0.007784f
C373 B.n189 VSUBS 0.007784f
C374 B.n190 VSUBS 0.007784f
C375 B.n191 VSUBS 0.007784f
C376 B.n192 VSUBS 0.007784f
C377 B.n193 VSUBS 0.007784f
C378 B.n194 VSUBS 0.016397f
C379 B.n195 VSUBS 0.017713f
C380 B.n196 VSUBS 0.017713f
C381 B.n197 VSUBS 0.007784f
C382 B.n198 VSUBS 0.007784f
C383 B.n199 VSUBS 0.007784f
C384 B.n200 VSUBS 0.007784f
C385 B.n201 VSUBS 0.007784f
C386 B.n202 VSUBS 0.007784f
C387 B.n203 VSUBS 0.007784f
C388 B.n204 VSUBS 0.007784f
C389 B.n205 VSUBS 0.007784f
C390 B.n206 VSUBS 0.007784f
C391 B.n207 VSUBS 0.007784f
C392 B.n208 VSUBS 0.007784f
C393 B.n209 VSUBS 0.007784f
C394 B.n210 VSUBS 0.007784f
C395 B.n211 VSUBS 0.007784f
C396 B.n212 VSUBS 0.007784f
C397 B.n213 VSUBS 0.007784f
C398 B.n214 VSUBS 0.007784f
C399 B.n215 VSUBS 0.007784f
C400 B.n216 VSUBS 0.007784f
C401 B.n217 VSUBS 0.007784f
C402 B.n218 VSUBS 0.007784f
C403 B.n219 VSUBS 0.007784f
C404 B.n220 VSUBS 0.007784f
C405 B.n221 VSUBS 0.007784f
C406 B.n222 VSUBS 0.007784f
C407 B.n223 VSUBS 0.007784f
C408 B.n224 VSUBS 0.007784f
C409 B.n225 VSUBS 0.007784f
C410 B.n226 VSUBS 0.007784f
C411 B.n227 VSUBS 0.007784f
C412 B.n228 VSUBS 0.007784f
C413 B.n229 VSUBS 0.007784f
C414 B.n230 VSUBS 0.007784f
C415 B.n231 VSUBS 0.007784f
C416 B.n232 VSUBS 0.007784f
C417 B.n233 VSUBS 0.007784f
C418 B.n234 VSUBS 0.007784f
C419 B.n235 VSUBS 0.007784f
C420 B.n236 VSUBS 0.00538f
C421 B.n237 VSUBS 0.018034f
C422 B.n238 VSUBS 0.006296f
C423 B.n239 VSUBS 0.007784f
C424 B.n240 VSUBS 0.007784f
C425 B.n241 VSUBS 0.007784f
C426 B.n242 VSUBS 0.007784f
C427 B.n243 VSUBS 0.007784f
C428 B.n244 VSUBS 0.007784f
C429 B.n245 VSUBS 0.007784f
C430 B.n246 VSUBS 0.007784f
C431 B.n247 VSUBS 0.007784f
C432 B.n248 VSUBS 0.007784f
C433 B.n249 VSUBS 0.007784f
C434 B.t11 VSUBS 0.12321f
C435 B.t10 VSUBS 0.140228f
C436 B.t9 VSUBS 0.4351f
C437 B.n250 VSUBS 0.238659f
C438 B.n251 VSUBS 0.191733f
C439 B.n252 VSUBS 0.018034f
C440 B.n253 VSUBS 0.006296f
C441 B.n254 VSUBS 0.007784f
C442 B.n255 VSUBS 0.007784f
C443 B.n256 VSUBS 0.007784f
C444 B.n257 VSUBS 0.007784f
C445 B.n258 VSUBS 0.007784f
C446 B.n259 VSUBS 0.007784f
C447 B.n260 VSUBS 0.007784f
C448 B.n261 VSUBS 0.007784f
C449 B.n262 VSUBS 0.007784f
C450 B.n263 VSUBS 0.007784f
C451 B.n264 VSUBS 0.007784f
C452 B.n265 VSUBS 0.007784f
C453 B.n266 VSUBS 0.007784f
C454 B.n267 VSUBS 0.007784f
C455 B.n268 VSUBS 0.007784f
C456 B.n269 VSUBS 0.007784f
C457 B.n270 VSUBS 0.007784f
C458 B.n271 VSUBS 0.007784f
C459 B.n272 VSUBS 0.007784f
C460 B.n273 VSUBS 0.007784f
C461 B.n274 VSUBS 0.007784f
C462 B.n275 VSUBS 0.007784f
C463 B.n276 VSUBS 0.007784f
C464 B.n277 VSUBS 0.007784f
C465 B.n278 VSUBS 0.007784f
C466 B.n279 VSUBS 0.007784f
C467 B.n280 VSUBS 0.007784f
C468 B.n281 VSUBS 0.007784f
C469 B.n282 VSUBS 0.007784f
C470 B.n283 VSUBS 0.007784f
C471 B.n284 VSUBS 0.007784f
C472 B.n285 VSUBS 0.007784f
C473 B.n286 VSUBS 0.007784f
C474 B.n287 VSUBS 0.007784f
C475 B.n288 VSUBS 0.007784f
C476 B.n289 VSUBS 0.007784f
C477 B.n290 VSUBS 0.007784f
C478 B.n291 VSUBS 0.007784f
C479 B.n292 VSUBS 0.007784f
C480 B.n293 VSUBS 0.007784f
C481 B.n294 VSUBS 0.007784f
C482 B.n295 VSUBS 0.016695f
C483 B.n296 VSUBS 0.017713f
C484 B.n297 VSUBS 0.016397f
C485 B.n298 VSUBS 0.007784f
C486 B.n299 VSUBS 0.007784f
C487 B.n300 VSUBS 0.007784f
C488 B.n301 VSUBS 0.007784f
C489 B.n302 VSUBS 0.007784f
C490 B.n303 VSUBS 0.007784f
C491 B.n304 VSUBS 0.007784f
C492 B.n305 VSUBS 0.007784f
C493 B.n306 VSUBS 0.007784f
C494 B.n307 VSUBS 0.007784f
C495 B.n308 VSUBS 0.007784f
C496 B.n309 VSUBS 0.007784f
C497 B.n310 VSUBS 0.007784f
C498 B.n311 VSUBS 0.007784f
C499 B.n312 VSUBS 0.007784f
C500 B.n313 VSUBS 0.007784f
C501 B.n314 VSUBS 0.007784f
C502 B.n315 VSUBS 0.007784f
C503 B.n316 VSUBS 0.007784f
C504 B.n317 VSUBS 0.007784f
C505 B.n318 VSUBS 0.007784f
C506 B.n319 VSUBS 0.007784f
C507 B.n320 VSUBS 0.007784f
C508 B.n321 VSUBS 0.007784f
C509 B.n322 VSUBS 0.007784f
C510 B.n323 VSUBS 0.007784f
C511 B.n324 VSUBS 0.007784f
C512 B.n325 VSUBS 0.007784f
C513 B.n326 VSUBS 0.007784f
C514 B.n327 VSUBS 0.007784f
C515 B.n328 VSUBS 0.007784f
C516 B.n329 VSUBS 0.007784f
C517 B.n330 VSUBS 0.007784f
C518 B.n331 VSUBS 0.007784f
C519 B.n332 VSUBS 0.007784f
C520 B.n333 VSUBS 0.007784f
C521 B.n334 VSUBS 0.007784f
C522 B.n335 VSUBS 0.007784f
C523 B.n336 VSUBS 0.007784f
C524 B.n337 VSUBS 0.007784f
C525 B.n338 VSUBS 0.007784f
C526 B.n339 VSUBS 0.007784f
C527 B.n340 VSUBS 0.007784f
C528 B.n341 VSUBS 0.007784f
C529 B.n342 VSUBS 0.007784f
C530 B.n343 VSUBS 0.007784f
C531 B.n344 VSUBS 0.007784f
C532 B.n345 VSUBS 0.007784f
C533 B.n346 VSUBS 0.007784f
C534 B.n347 VSUBS 0.007784f
C535 B.n348 VSUBS 0.007784f
C536 B.n349 VSUBS 0.007784f
C537 B.n350 VSUBS 0.007784f
C538 B.n351 VSUBS 0.007784f
C539 B.n352 VSUBS 0.007784f
C540 B.n353 VSUBS 0.007784f
C541 B.n354 VSUBS 0.007784f
C542 B.n355 VSUBS 0.007784f
C543 B.n356 VSUBS 0.007784f
C544 B.n357 VSUBS 0.007784f
C545 B.n358 VSUBS 0.007784f
C546 B.n359 VSUBS 0.007784f
C547 B.n360 VSUBS 0.007784f
C548 B.n361 VSUBS 0.007784f
C549 B.n362 VSUBS 0.007784f
C550 B.n363 VSUBS 0.007784f
C551 B.n364 VSUBS 0.007784f
C552 B.n365 VSUBS 0.007784f
C553 B.n366 VSUBS 0.007784f
C554 B.n367 VSUBS 0.007784f
C555 B.n368 VSUBS 0.007784f
C556 B.n369 VSUBS 0.007784f
C557 B.n370 VSUBS 0.007784f
C558 B.n371 VSUBS 0.007784f
C559 B.n372 VSUBS 0.007784f
C560 B.n373 VSUBS 0.007784f
C561 B.n374 VSUBS 0.007784f
C562 B.n375 VSUBS 0.007784f
C563 B.n376 VSUBS 0.007784f
C564 B.n377 VSUBS 0.007784f
C565 B.n378 VSUBS 0.007784f
C566 B.n379 VSUBS 0.007784f
C567 B.n380 VSUBS 0.007784f
C568 B.n381 VSUBS 0.007784f
C569 B.n382 VSUBS 0.007784f
C570 B.n383 VSUBS 0.007784f
C571 B.n384 VSUBS 0.007784f
C572 B.n385 VSUBS 0.007784f
C573 B.n386 VSUBS 0.007784f
C574 B.n387 VSUBS 0.007784f
C575 B.n388 VSUBS 0.007784f
C576 B.n389 VSUBS 0.007784f
C577 B.n390 VSUBS 0.007784f
C578 B.n391 VSUBS 0.007784f
C579 B.n392 VSUBS 0.007784f
C580 B.n393 VSUBS 0.007784f
C581 B.n394 VSUBS 0.007784f
C582 B.n395 VSUBS 0.007784f
C583 B.n396 VSUBS 0.007784f
C584 B.n397 VSUBS 0.007784f
C585 B.n398 VSUBS 0.007784f
C586 B.n399 VSUBS 0.007784f
C587 B.n400 VSUBS 0.007784f
C588 B.n401 VSUBS 0.007784f
C589 B.n402 VSUBS 0.007784f
C590 B.n403 VSUBS 0.016397f
C591 B.n404 VSUBS 0.016397f
C592 B.n405 VSUBS 0.017713f
C593 B.n406 VSUBS 0.007784f
C594 B.n407 VSUBS 0.007784f
C595 B.n408 VSUBS 0.007784f
C596 B.n409 VSUBS 0.007784f
C597 B.n410 VSUBS 0.007784f
C598 B.n411 VSUBS 0.007784f
C599 B.n412 VSUBS 0.007784f
C600 B.n413 VSUBS 0.007784f
C601 B.n414 VSUBS 0.007784f
C602 B.n415 VSUBS 0.007784f
C603 B.n416 VSUBS 0.007784f
C604 B.n417 VSUBS 0.007784f
C605 B.n418 VSUBS 0.007784f
C606 B.n419 VSUBS 0.007784f
C607 B.n420 VSUBS 0.007784f
C608 B.n421 VSUBS 0.007784f
C609 B.n422 VSUBS 0.007784f
C610 B.n423 VSUBS 0.007784f
C611 B.n424 VSUBS 0.007784f
C612 B.n425 VSUBS 0.007784f
C613 B.n426 VSUBS 0.007784f
C614 B.n427 VSUBS 0.007784f
C615 B.n428 VSUBS 0.007784f
C616 B.n429 VSUBS 0.007784f
C617 B.n430 VSUBS 0.007784f
C618 B.n431 VSUBS 0.007784f
C619 B.n432 VSUBS 0.007784f
C620 B.n433 VSUBS 0.007784f
C621 B.n434 VSUBS 0.007784f
C622 B.n435 VSUBS 0.007784f
C623 B.n436 VSUBS 0.007784f
C624 B.n437 VSUBS 0.007784f
C625 B.n438 VSUBS 0.007784f
C626 B.n439 VSUBS 0.007784f
C627 B.n440 VSUBS 0.007784f
C628 B.n441 VSUBS 0.007784f
C629 B.n442 VSUBS 0.007784f
C630 B.n443 VSUBS 0.007784f
C631 B.n444 VSUBS 0.007784f
C632 B.n445 VSUBS 0.00538f
C633 B.n446 VSUBS 0.007784f
C634 B.n447 VSUBS 0.007784f
C635 B.n448 VSUBS 0.006296f
C636 B.n449 VSUBS 0.007784f
C637 B.n450 VSUBS 0.007784f
C638 B.n451 VSUBS 0.007784f
C639 B.n452 VSUBS 0.007784f
C640 B.n453 VSUBS 0.007784f
C641 B.n454 VSUBS 0.007784f
C642 B.n455 VSUBS 0.007784f
C643 B.n456 VSUBS 0.007784f
C644 B.n457 VSUBS 0.007784f
C645 B.n458 VSUBS 0.007784f
C646 B.n459 VSUBS 0.007784f
C647 B.n460 VSUBS 0.006296f
C648 B.n461 VSUBS 0.018034f
C649 B.n462 VSUBS 0.00538f
C650 B.n463 VSUBS 0.007784f
C651 B.n464 VSUBS 0.007784f
C652 B.n465 VSUBS 0.007784f
C653 B.n466 VSUBS 0.007784f
C654 B.n467 VSUBS 0.007784f
C655 B.n468 VSUBS 0.007784f
C656 B.n469 VSUBS 0.007784f
C657 B.n470 VSUBS 0.007784f
C658 B.n471 VSUBS 0.007784f
C659 B.n472 VSUBS 0.007784f
C660 B.n473 VSUBS 0.007784f
C661 B.n474 VSUBS 0.007784f
C662 B.n475 VSUBS 0.007784f
C663 B.n476 VSUBS 0.007784f
C664 B.n477 VSUBS 0.007784f
C665 B.n478 VSUBS 0.007784f
C666 B.n479 VSUBS 0.007784f
C667 B.n480 VSUBS 0.007784f
C668 B.n481 VSUBS 0.007784f
C669 B.n482 VSUBS 0.007784f
C670 B.n483 VSUBS 0.007784f
C671 B.n484 VSUBS 0.007784f
C672 B.n485 VSUBS 0.007784f
C673 B.n486 VSUBS 0.007784f
C674 B.n487 VSUBS 0.007784f
C675 B.n488 VSUBS 0.007784f
C676 B.n489 VSUBS 0.007784f
C677 B.n490 VSUBS 0.007784f
C678 B.n491 VSUBS 0.007784f
C679 B.n492 VSUBS 0.007784f
C680 B.n493 VSUBS 0.007784f
C681 B.n494 VSUBS 0.007784f
C682 B.n495 VSUBS 0.007784f
C683 B.n496 VSUBS 0.007784f
C684 B.n497 VSUBS 0.007784f
C685 B.n498 VSUBS 0.007784f
C686 B.n499 VSUBS 0.007784f
C687 B.n500 VSUBS 0.007784f
C688 B.n501 VSUBS 0.007784f
C689 B.n502 VSUBS 0.017713f
C690 B.n503 VSUBS 0.017713f
C691 B.n504 VSUBS 0.016397f
C692 B.n505 VSUBS 0.007784f
C693 B.n506 VSUBS 0.007784f
C694 B.n507 VSUBS 0.007784f
C695 B.n508 VSUBS 0.007784f
C696 B.n509 VSUBS 0.007784f
C697 B.n510 VSUBS 0.007784f
C698 B.n511 VSUBS 0.007784f
C699 B.n512 VSUBS 0.007784f
C700 B.n513 VSUBS 0.007784f
C701 B.n514 VSUBS 0.007784f
C702 B.n515 VSUBS 0.007784f
C703 B.n516 VSUBS 0.007784f
C704 B.n517 VSUBS 0.007784f
C705 B.n518 VSUBS 0.007784f
C706 B.n519 VSUBS 0.007784f
C707 B.n520 VSUBS 0.007784f
C708 B.n521 VSUBS 0.007784f
C709 B.n522 VSUBS 0.007784f
C710 B.n523 VSUBS 0.007784f
C711 B.n524 VSUBS 0.007784f
C712 B.n525 VSUBS 0.007784f
C713 B.n526 VSUBS 0.007784f
C714 B.n527 VSUBS 0.007784f
C715 B.n528 VSUBS 0.007784f
C716 B.n529 VSUBS 0.007784f
C717 B.n530 VSUBS 0.007784f
C718 B.n531 VSUBS 0.007784f
C719 B.n532 VSUBS 0.007784f
C720 B.n533 VSUBS 0.007784f
C721 B.n534 VSUBS 0.007784f
C722 B.n535 VSUBS 0.007784f
C723 B.n536 VSUBS 0.007784f
C724 B.n537 VSUBS 0.007784f
C725 B.n538 VSUBS 0.007784f
C726 B.n539 VSUBS 0.007784f
C727 B.n540 VSUBS 0.007784f
C728 B.n541 VSUBS 0.007784f
C729 B.n542 VSUBS 0.007784f
C730 B.n543 VSUBS 0.007784f
C731 B.n544 VSUBS 0.007784f
C732 B.n545 VSUBS 0.007784f
C733 B.n546 VSUBS 0.007784f
C734 B.n547 VSUBS 0.007784f
C735 B.n548 VSUBS 0.007784f
C736 B.n549 VSUBS 0.007784f
C737 B.n550 VSUBS 0.007784f
C738 B.n551 VSUBS 0.007784f
C739 B.n552 VSUBS 0.007784f
C740 B.n553 VSUBS 0.007784f
C741 B.n554 VSUBS 0.007784f
C742 B.n555 VSUBS 0.010157f
C743 B.n556 VSUBS 0.01082f
C744 B.n557 VSUBS 0.021517f
C745 VTAIL.t12 VSUBS 0.172681f
C746 VTAIL.t8 VSUBS 0.172681f
C747 VTAIL.n0 VSUBS 1.10344f
C748 VTAIL.n1 VSUBS 0.790947f
C749 VTAIL.n2 VSUBS 0.032081f
C750 VTAIL.n3 VSUBS 0.030392f
C751 VTAIL.n4 VSUBS 0.016331f
C752 VTAIL.n5 VSUBS 0.038602f
C753 VTAIL.n6 VSUBS 0.017292f
C754 VTAIL.n7 VSUBS 0.030392f
C755 VTAIL.n8 VSUBS 0.016331f
C756 VTAIL.n9 VSUBS 0.038602f
C757 VTAIL.n10 VSUBS 0.017292f
C758 VTAIL.n11 VSUBS 0.852358f
C759 VTAIL.n12 VSUBS 0.016331f
C760 VTAIL.t2 VSUBS 0.082894f
C761 VTAIL.n13 VSUBS 0.173426f
C762 VTAIL.n14 VSUBS 0.029037f
C763 VTAIL.n15 VSUBS 0.028951f
C764 VTAIL.n16 VSUBS 0.038602f
C765 VTAIL.n17 VSUBS 0.017292f
C766 VTAIL.n18 VSUBS 0.016331f
C767 VTAIL.n19 VSUBS 0.030392f
C768 VTAIL.n20 VSUBS 0.030392f
C769 VTAIL.n21 VSUBS 0.016331f
C770 VTAIL.n22 VSUBS 0.017292f
C771 VTAIL.n23 VSUBS 0.038602f
C772 VTAIL.n24 VSUBS 0.038602f
C773 VTAIL.n25 VSUBS 0.017292f
C774 VTAIL.n26 VSUBS 0.016331f
C775 VTAIL.n27 VSUBS 0.030392f
C776 VTAIL.n28 VSUBS 0.030392f
C777 VTAIL.n29 VSUBS 0.016331f
C778 VTAIL.n30 VSUBS 0.017292f
C779 VTAIL.n31 VSUBS 0.038602f
C780 VTAIL.n32 VSUBS 0.094681f
C781 VTAIL.n33 VSUBS 0.017292f
C782 VTAIL.n34 VSUBS 0.032071f
C783 VTAIL.n35 VSUBS 0.074817f
C784 VTAIL.n36 VSUBS 0.071878f
C785 VTAIL.n37 VSUBS 0.270832f
C786 VTAIL.t7 VSUBS 0.172681f
C787 VTAIL.t4 VSUBS 0.172681f
C788 VTAIL.n38 VSUBS 1.10344f
C789 VTAIL.n39 VSUBS 0.83738f
C790 VTAIL.t3 VSUBS 0.172681f
C791 VTAIL.t1 VSUBS 0.172681f
C792 VTAIL.n40 VSUBS 1.10344f
C793 VTAIL.n41 VSUBS 1.98808f
C794 VTAIL.t9 VSUBS 0.172681f
C795 VTAIL.t17 VSUBS 0.172681f
C796 VTAIL.n42 VSUBS 1.10345f
C797 VTAIL.n43 VSUBS 1.98807f
C798 VTAIL.t16 VSUBS 0.172681f
C799 VTAIL.t14 VSUBS 0.172681f
C800 VTAIL.n44 VSUBS 1.10345f
C801 VTAIL.n45 VSUBS 0.837372f
C802 VTAIL.n46 VSUBS 0.032081f
C803 VTAIL.n47 VSUBS 0.030392f
C804 VTAIL.n48 VSUBS 0.016331f
C805 VTAIL.n49 VSUBS 0.038602f
C806 VTAIL.n50 VSUBS 0.017292f
C807 VTAIL.n51 VSUBS 0.030392f
C808 VTAIL.n52 VSUBS 0.016331f
C809 VTAIL.n53 VSUBS 0.038602f
C810 VTAIL.n54 VSUBS 0.017292f
C811 VTAIL.n55 VSUBS 0.852358f
C812 VTAIL.n56 VSUBS 0.016331f
C813 VTAIL.t13 VSUBS 0.082894f
C814 VTAIL.n57 VSUBS 0.173426f
C815 VTAIL.n58 VSUBS 0.029037f
C816 VTAIL.n59 VSUBS 0.028951f
C817 VTAIL.n60 VSUBS 0.038602f
C818 VTAIL.n61 VSUBS 0.017292f
C819 VTAIL.n62 VSUBS 0.016331f
C820 VTAIL.n63 VSUBS 0.030392f
C821 VTAIL.n64 VSUBS 0.030392f
C822 VTAIL.n65 VSUBS 0.016331f
C823 VTAIL.n66 VSUBS 0.017292f
C824 VTAIL.n67 VSUBS 0.038602f
C825 VTAIL.n68 VSUBS 0.038602f
C826 VTAIL.n69 VSUBS 0.017292f
C827 VTAIL.n70 VSUBS 0.016331f
C828 VTAIL.n71 VSUBS 0.030392f
C829 VTAIL.n72 VSUBS 0.030392f
C830 VTAIL.n73 VSUBS 0.016331f
C831 VTAIL.n74 VSUBS 0.017292f
C832 VTAIL.n75 VSUBS 0.038602f
C833 VTAIL.n76 VSUBS 0.094681f
C834 VTAIL.n77 VSUBS 0.017292f
C835 VTAIL.n78 VSUBS 0.032071f
C836 VTAIL.n79 VSUBS 0.074817f
C837 VTAIL.n80 VSUBS 0.071878f
C838 VTAIL.n81 VSUBS 0.270832f
C839 VTAIL.t6 VSUBS 0.172681f
C840 VTAIL.t5 VSUBS 0.172681f
C841 VTAIL.n82 VSUBS 1.10345f
C842 VTAIL.n83 VSUBS 0.817954f
C843 VTAIL.t18 VSUBS 0.172681f
C844 VTAIL.t0 VSUBS 0.172681f
C845 VTAIL.n84 VSUBS 1.10345f
C846 VTAIL.n85 VSUBS 0.837372f
C847 VTAIL.n86 VSUBS 0.032081f
C848 VTAIL.n87 VSUBS 0.030392f
C849 VTAIL.n88 VSUBS 0.016331f
C850 VTAIL.n89 VSUBS 0.038602f
C851 VTAIL.n90 VSUBS 0.017292f
C852 VTAIL.n91 VSUBS 0.030392f
C853 VTAIL.n92 VSUBS 0.016331f
C854 VTAIL.n93 VSUBS 0.038602f
C855 VTAIL.n94 VSUBS 0.017292f
C856 VTAIL.n95 VSUBS 0.852358f
C857 VTAIL.n96 VSUBS 0.016331f
C858 VTAIL.t19 VSUBS 0.082894f
C859 VTAIL.n97 VSUBS 0.173426f
C860 VTAIL.n98 VSUBS 0.029037f
C861 VTAIL.n99 VSUBS 0.028951f
C862 VTAIL.n100 VSUBS 0.038602f
C863 VTAIL.n101 VSUBS 0.017292f
C864 VTAIL.n102 VSUBS 0.016331f
C865 VTAIL.n103 VSUBS 0.030392f
C866 VTAIL.n104 VSUBS 0.030392f
C867 VTAIL.n105 VSUBS 0.016331f
C868 VTAIL.n106 VSUBS 0.017292f
C869 VTAIL.n107 VSUBS 0.038602f
C870 VTAIL.n108 VSUBS 0.038602f
C871 VTAIL.n109 VSUBS 0.017292f
C872 VTAIL.n110 VSUBS 0.016331f
C873 VTAIL.n111 VSUBS 0.030392f
C874 VTAIL.n112 VSUBS 0.030392f
C875 VTAIL.n113 VSUBS 0.016331f
C876 VTAIL.n114 VSUBS 0.017292f
C877 VTAIL.n115 VSUBS 0.038602f
C878 VTAIL.n116 VSUBS 0.094681f
C879 VTAIL.n117 VSUBS 0.017292f
C880 VTAIL.n118 VSUBS 0.032071f
C881 VTAIL.n119 VSUBS 0.074817f
C882 VTAIL.n120 VSUBS 0.071878f
C883 VTAIL.n121 VSUBS 1.31009f
C884 VTAIL.n122 VSUBS 0.032081f
C885 VTAIL.n123 VSUBS 0.030392f
C886 VTAIL.n124 VSUBS 0.016331f
C887 VTAIL.n125 VSUBS 0.038602f
C888 VTAIL.n126 VSUBS 0.017292f
C889 VTAIL.n127 VSUBS 0.030392f
C890 VTAIL.n128 VSUBS 0.016331f
C891 VTAIL.n129 VSUBS 0.038602f
C892 VTAIL.n130 VSUBS 0.017292f
C893 VTAIL.n131 VSUBS 0.852358f
C894 VTAIL.n132 VSUBS 0.016331f
C895 VTAIL.t11 VSUBS 0.082894f
C896 VTAIL.n133 VSUBS 0.173426f
C897 VTAIL.n134 VSUBS 0.029037f
C898 VTAIL.n135 VSUBS 0.028951f
C899 VTAIL.n136 VSUBS 0.038602f
C900 VTAIL.n137 VSUBS 0.017292f
C901 VTAIL.n138 VSUBS 0.016331f
C902 VTAIL.n139 VSUBS 0.030392f
C903 VTAIL.n140 VSUBS 0.030392f
C904 VTAIL.n141 VSUBS 0.016331f
C905 VTAIL.n142 VSUBS 0.017292f
C906 VTAIL.n143 VSUBS 0.038602f
C907 VTAIL.n144 VSUBS 0.038602f
C908 VTAIL.n145 VSUBS 0.017292f
C909 VTAIL.n146 VSUBS 0.016331f
C910 VTAIL.n147 VSUBS 0.030392f
C911 VTAIL.n148 VSUBS 0.030392f
C912 VTAIL.n149 VSUBS 0.016331f
C913 VTAIL.n150 VSUBS 0.017292f
C914 VTAIL.n151 VSUBS 0.038602f
C915 VTAIL.n152 VSUBS 0.094681f
C916 VTAIL.n153 VSUBS 0.017292f
C917 VTAIL.n154 VSUBS 0.032071f
C918 VTAIL.n155 VSUBS 0.074817f
C919 VTAIL.n156 VSUBS 0.071878f
C920 VTAIL.n157 VSUBS 1.31009f
C921 VTAIL.t10 VSUBS 0.172681f
C922 VTAIL.t15 VSUBS 0.172681f
C923 VTAIL.n158 VSUBS 1.10344f
C924 VTAIL.n159 VSUBS 0.73354f
C925 VDD2.n0 VSUBS 0.024199f
C926 VDD2.n1 VSUBS 0.022925f
C927 VDD2.n2 VSUBS 0.012319f
C928 VDD2.n3 VSUBS 0.029118f
C929 VDD2.n4 VSUBS 0.013044f
C930 VDD2.n5 VSUBS 0.022925f
C931 VDD2.n6 VSUBS 0.012319f
C932 VDD2.n7 VSUBS 0.029118f
C933 VDD2.n8 VSUBS 0.013044f
C934 VDD2.n9 VSUBS 0.642943f
C935 VDD2.n10 VSUBS 0.012319f
C936 VDD2.t1 VSUBS 0.062528f
C937 VDD2.n11 VSUBS 0.130817f
C938 VDD2.n12 VSUBS 0.021903f
C939 VDD2.n13 VSUBS 0.021838f
C940 VDD2.n14 VSUBS 0.029118f
C941 VDD2.n15 VSUBS 0.013044f
C942 VDD2.n16 VSUBS 0.012319f
C943 VDD2.n17 VSUBS 0.022925f
C944 VDD2.n18 VSUBS 0.022925f
C945 VDD2.n19 VSUBS 0.012319f
C946 VDD2.n20 VSUBS 0.013044f
C947 VDD2.n21 VSUBS 0.029118f
C948 VDD2.n22 VSUBS 0.029118f
C949 VDD2.n23 VSUBS 0.013044f
C950 VDD2.n24 VSUBS 0.012319f
C951 VDD2.n25 VSUBS 0.022925f
C952 VDD2.n26 VSUBS 0.022925f
C953 VDD2.n27 VSUBS 0.012319f
C954 VDD2.n28 VSUBS 0.013044f
C955 VDD2.n29 VSUBS 0.029118f
C956 VDD2.n30 VSUBS 0.071419f
C957 VDD2.n31 VSUBS 0.013044f
C958 VDD2.n32 VSUBS 0.024192f
C959 VDD2.n33 VSUBS 0.056436f
C960 VDD2.n34 VSUBS 0.07372f
C961 VDD2.t7 VSUBS 0.130255f
C962 VDD2.t2 VSUBS 0.130255f
C963 VDD2.n35 VSUBS 0.920753f
C964 VDD2.n36 VSUBS 0.639306f
C965 VDD2.t9 VSUBS 0.130255f
C966 VDD2.t4 VSUBS 0.130255f
C967 VDD2.n37 VSUBS 0.926735f
C968 VDD2.n38 VSUBS 1.92128f
C969 VDD2.n39 VSUBS 0.024199f
C970 VDD2.n40 VSUBS 0.022925f
C971 VDD2.n41 VSUBS 0.012319f
C972 VDD2.n42 VSUBS 0.029118f
C973 VDD2.n43 VSUBS 0.013044f
C974 VDD2.n44 VSUBS 0.022925f
C975 VDD2.n45 VSUBS 0.012319f
C976 VDD2.n46 VSUBS 0.029118f
C977 VDD2.n47 VSUBS 0.013044f
C978 VDD2.n48 VSUBS 0.642943f
C979 VDD2.n49 VSUBS 0.012319f
C980 VDD2.t8 VSUBS 0.062528f
C981 VDD2.n50 VSUBS 0.130817f
C982 VDD2.n51 VSUBS 0.021903f
C983 VDD2.n52 VSUBS 0.021838f
C984 VDD2.n53 VSUBS 0.029118f
C985 VDD2.n54 VSUBS 0.013044f
C986 VDD2.n55 VSUBS 0.012319f
C987 VDD2.n56 VSUBS 0.022925f
C988 VDD2.n57 VSUBS 0.022925f
C989 VDD2.n58 VSUBS 0.012319f
C990 VDD2.n59 VSUBS 0.013044f
C991 VDD2.n60 VSUBS 0.029118f
C992 VDD2.n61 VSUBS 0.029118f
C993 VDD2.n62 VSUBS 0.013044f
C994 VDD2.n63 VSUBS 0.012319f
C995 VDD2.n64 VSUBS 0.022925f
C996 VDD2.n65 VSUBS 0.022925f
C997 VDD2.n66 VSUBS 0.012319f
C998 VDD2.n67 VSUBS 0.013044f
C999 VDD2.n68 VSUBS 0.029118f
C1000 VDD2.n69 VSUBS 0.071419f
C1001 VDD2.n70 VSUBS 0.013044f
C1002 VDD2.n71 VSUBS 0.024192f
C1003 VDD2.n72 VSUBS 0.056436f
C1004 VDD2.n73 VSUBS 0.070023f
C1005 VDD2.n74 VSUBS 1.81447f
C1006 VDD2.t6 VSUBS 0.130255f
C1007 VDD2.t3 VSUBS 0.130255f
C1008 VDD2.n75 VSUBS 0.920758f
C1009 VDD2.n76 VSUBS 0.504656f
C1010 VDD2.t5 VSUBS 0.130255f
C1011 VDD2.t0 VSUBS 0.130255f
C1012 VDD2.n77 VSUBS 0.926709f
C1013 VN.n0 VSUBS 0.061632f
C1014 VN.t2 VSUBS 1.08279f
C1015 VN.n1 VSUBS 0.420976f
C1016 VN.n2 VSUBS 0.046188f
C1017 VN.t7 VSUBS 1.08279f
C1018 VN.n3 VSUBS 0.420976f
C1019 VN.n4 VSUBS 0.046188f
C1020 VN.t9 VSUBS 1.08279f
C1021 VN.n5 VSUBS 0.482925f
C1022 VN.t5 VSUBS 1.22225f
C1023 VN.n6 VSUBS 0.496473f
C1024 VN.n7 VSUBS 0.240719f
C1025 VN.n8 VSUBS 0.073469f
C1026 VN.n9 VSUBS 0.037713f
C1027 VN.n10 VSUBS 0.071513f
C1028 VN.n11 VSUBS 0.046188f
C1029 VN.n12 VSUBS 0.046188f
C1030 VN.n13 VSUBS 0.071513f
C1031 VN.n14 VSUBS 0.037713f
C1032 VN.n15 VSUBS 0.073469f
C1033 VN.n16 VSUBS 0.046188f
C1034 VN.n17 VSUBS 0.046188f
C1035 VN.n18 VSUBS 0.067743f
C1036 VN.n19 VSUBS 0.033084f
C1037 VN.t6 VSUBS 1.16912f
C1038 VN.n20 VSUBS 0.508548f
C1039 VN.n21 VSUBS 0.043257f
C1040 VN.n22 VSUBS 0.061632f
C1041 VN.t0 VSUBS 1.08279f
C1042 VN.n23 VSUBS 0.420976f
C1043 VN.n24 VSUBS 0.046188f
C1044 VN.t1 VSUBS 1.08279f
C1045 VN.n25 VSUBS 0.420976f
C1046 VN.n26 VSUBS 0.046188f
C1047 VN.t3 VSUBS 1.08279f
C1048 VN.n27 VSUBS 0.482925f
C1049 VN.t4 VSUBS 1.22225f
C1050 VN.n28 VSUBS 0.496473f
C1051 VN.n29 VSUBS 0.240719f
C1052 VN.n30 VSUBS 0.073469f
C1053 VN.n31 VSUBS 0.037713f
C1054 VN.n32 VSUBS 0.071513f
C1055 VN.n33 VSUBS 0.046188f
C1056 VN.n34 VSUBS 0.046188f
C1057 VN.n35 VSUBS 0.071513f
C1058 VN.n36 VSUBS 0.037713f
C1059 VN.n37 VSUBS 0.073469f
C1060 VN.n38 VSUBS 0.046188f
C1061 VN.n39 VSUBS 0.046188f
C1062 VN.n40 VSUBS 0.067743f
C1063 VN.n41 VSUBS 0.033084f
C1064 VN.t8 VSUBS 1.16912f
C1065 VN.n42 VSUBS 0.508548f
C1066 VN.n43 VSUBS 1.9584f
.ends

