* NGSPICE file created from diff_pair_sample_0668.ext - technology: sky130A

.subckt diff_pair_sample_0668 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3770_n1948# sky130_fd_pr__pfet_01v8 ad=1.911 pd=10.58 as=0 ps=0 w=4.9 l=2.47
X1 B.t8 B.t6 B.t7 w_n3770_n1948# sky130_fd_pr__pfet_01v8 ad=1.911 pd=10.58 as=0 ps=0 w=4.9 l=2.47
X2 VDD2.t7 VN.t0 VTAIL.t9 w_n3770_n1948# sky130_fd_pr__pfet_01v8 ad=0.8085 pd=5.23 as=1.911 ps=10.58 w=4.9 l=2.47
X3 VTAIL.t5 VP.t0 VDD1.t7 w_n3770_n1948# sky130_fd_pr__pfet_01v8 ad=1.911 pd=10.58 as=0.8085 ps=5.23 w=4.9 l=2.47
X4 VDD2.t6 VN.t1 VTAIL.t8 w_n3770_n1948# sky130_fd_pr__pfet_01v8 ad=0.8085 pd=5.23 as=1.911 ps=10.58 w=4.9 l=2.47
X5 VTAIL.t10 VN.t2 VDD2.t5 w_n3770_n1948# sky130_fd_pr__pfet_01v8 ad=1.911 pd=10.58 as=0.8085 ps=5.23 w=4.9 l=2.47
X6 B.t5 B.t3 B.t4 w_n3770_n1948# sky130_fd_pr__pfet_01v8 ad=1.911 pd=10.58 as=0 ps=0 w=4.9 l=2.47
X7 VDD2.t4 VN.t3 VTAIL.t12 w_n3770_n1948# sky130_fd_pr__pfet_01v8 ad=0.8085 pd=5.23 as=0.8085 ps=5.23 w=4.9 l=2.47
X8 VDD1.t6 VP.t1 VTAIL.t4 w_n3770_n1948# sky130_fd_pr__pfet_01v8 ad=0.8085 pd=5.23 as=1.911 ps=10.58 w=4.9 l=2.47
X9 B.t2 B.t0 B.t1 w_n3770_n1948# sky130_fd_pr__pfet_01v8 ad=1.911 pd=10.58 as=0 ps=0 w=4.9 l=2.47
X10 VTAIL.t15 VN.t4 VDD2.t3 w_n3770_n1948# sky130_fd_pr__pfet_01v8 ad=0.8085 pd=5.23 as=0.8085 ps=5.23 w=4.9 l=2.47
X11 VDD1.t5 VP.t2 VTAIL.t3 w_n3770_n1948# sky130_fd_pr__pfet_01v8 ad=0.8085 pd=5.23 as=0.8085 ps=5.23 w=4.9 l=2.47
X12 VDD2.t2 VN.t5 VTAIL.t11 w_n3770_n1948# sky130_fd_pr__pfet_01v8 ad=0.8085 pd=5.23 as=0.8085 ps=5.23 w=4.9 l=2.47
X13 VTAIL.t2 VP.t3 VDD1.t4 w_n3770_n1948# sky130_fd_pr__pfet_01v8 ad=1.911 pd=10.58 as=0.8085 ps=5.23 w=4.9 l=2.47
X14 VDD1.t3 VP.t4 VTAIL.t1 w_n3770_n1948# sky130_fd_pr__pfet_01v8 ad=0.8085 pd=5.23 as=1.911 ps=10.58 w=4.9 l=2.47
X15 VDD1.t2 VP.t5 VTAIL.t0 w_n3770_n1948# sky130_fd_pr__pfet_01v8 ad=0.8085 pd=5.23 as=0.8085 ps=5.23 w=4.9 l=2.47
X16 VTAIL.t6 VP.t6 VDD1.t1 w_n3770_n1948# sky130_fd_pr__pfet_01v8 ad=0.8085 pd=5.23 as=0.8085 ps=5.23 w=4.9 l=2.47
X17 VTAIL.t14 VN.t6 VDD2.t1 w_n3770_n1948# sky130_fd_pr__pfet_01v8 ad=0.8085 pd=5.23 as=0.8085 ps=5.23 w=4.9 l=2.47
X18 VTAIL.t13 VN.t7 VDD2.t0 w_n3770_n1948# sky130_fd_pr__pfet_01v8 ad=1.911 pd=10.58 as=0.8085 ps=5.23 w=4.9 l=2.47
X19 VTAIL.t7 VP.t7 VDD1.t0 w_n3770_n1948# sky130_fd_pr__pfet_01v8 ad=0.8085 pd=5.23 as=0.8085 ps=5.23 w=4.9 l=2.47
R0 B.n309 B.n106 585
R1 B.n308 B.n307 585
R2 B.n306 B.n107 585
R3 B.n305 B.n304 585
R4 B.n303 B.n108 585
R5 B.n302 B.n301 585
R6 B.n300 B.n109 585
R7 B.n299 B.n298 585
R8 B.n297 B.n110 585
R9 B.n296 B.n295 585
R10 B.n294 B.n111 585
R11 B.n293 B.n292 585
R12 B.n291 B.n112 585
R13 B.n290 B.n289 585
R14 B.n288 B.n113 585
R15 B.n287 B.n286 585
R16 B.n285 B.n114 585
R17 B.n284 B.n283 585
R18 B.n282 B.n115 585
R19 B.n281 B.n280 585
R20 B.n279 B.n116 585
R21 B.n278 B.n277 585
R22 B.n273 B.n117 585
R23 B.n272 B.n271 585
R24 B.n270 B.n118 585
R25 B.n269 B.n268 585
R26 B.n267 B.n119 585
R27 B.n266 B.n265 585
R28 B.n264 B.n120 585
R29 B.n263 B.n262 585
R30 B.n260 B.n121 585
R31 B.n259 B.n258 585
R32 B.n257 B.n124 585
R33 B.n256 B.n255 585
R34 B.n254 B.n125 585
R35 B.n253 B.n252 585
R36 B.n251 B.n126 585
R37 B.n250 B.n249 585
R38 B.n248 B.n127 585
R39 B.n247 B.n246 585
R40 B.n245 B.n128 585
R41 B.n244 B.n243 585
R42 B.n242 B.n129 585
R43 B.n241 B.n240 585
R44 B.n239 B.n130 585
R45 B.n238 B.n237 585
R46 B.n236 B.n131 585
R47 B.n235 B.n234 585
R48 B.n233 B.n132 585
R49 B.n232 B.n231 585
R50 B.n230 B.n133 585
R51 B.n311 B.n310 585
R52 B.n312 B.n105 585
R53 B.n314 B.n313 585
R54 B.n315 B.n104 585
R55 B.n317 B.n316 585
R56 B.n318 B.n103 585
R57 B.n320 B.n319 585
R58 B.n321 B.n102 585
R59 B.n323 B.n322 585
R60 B.n324 B.n101 585
R61 B.n326 B.n325 585
R62 B.n327 B.n100 585
R63 B.n329 B.n328 585
R64 B.n330 B.n99 585
R65 B.n332 B.n331 585
R66 B.n333 B.n98 585
R67 B.n335 B.n334 585
R68 B.n336 B.n97 585
R69 B.n338 B.n337 585
R70 B.n339 B.n96 585
R71 B.n341 B.n340 585
R72 B.n342 B.n95 585
R73 B.n344 B.n343 585
R74 B.n345 B.n94 585
R75 B.n347 B.n346 585
R76 B.n348 B.n93 585
R77 B.n350 B.n349 585
R78 B.n351 B.n92 585
R79 B.n353 B.n352 585
R80 B.n354 B.n91 585
R81 B.n356 B.n355 585
R82 B.n357 B.n90 585
R83 B.n359 B.n358 585
R84 B.n360 B.n89 585
R85 B.n362 B.n361 585
R86 B.n363 B.n88 585
R87 B.n365 B.n364 585
R88 B.n366 B.n87 585
R89 B.n368 B.n367 585
R90 B.n369 B.n86 585
R91 B.n371 B.n370 585
R92 B.n372 B.n85 585
R93 B.n374 B.n373 585
R94 B.n375 B.n84 585
R95 B.n377 B.n376 585
R96 B.n378 B.n83 585
R97 B.n380 B.n379 585
R98 B.n381 B.n82 585
R99 B.n383 B.n382 585
R100 B.n384 B.n81 585
R101 B.n386 B.n385 585
R102 B.n387 B.n80 585
R103 B.n389 B.n388 585
R104 B.n390 B.n79 585
R105 B.n392 B.n391 585
R106 B.n393 B.n78 585
R107 B.n395 B.n394 585
R108 B.n396 B.n77 585
R109 B.n398 B.n397 585
R110 B.n399 B.n76 585
R111 B.n401 B.n400 585
R112 B.n402 B.n75 585
R113 B.n404 B.n403 585
R114 B.n405 B.n74 585
R115 B.n407 B.n406 585
R116 B.n408 B.n73 585
R117 B.n410 B.n409 585
R118 B.n411 B.n72 585
R119 B.n413 B.n412 585
R120 B.n414 B.n71 585
R121 B.n416 B.n415 585
R122 B.n417 B.n70 585
R123 B.n419 B.n418 585
R124 B.n420 B.n69 585
R125 B.n422 B.n421 585
R126 B.n423 B.n68 585
R127 B.n425 B.n424 585
R128 B.n426 B.n67 585
R129 B.n428 B.n427 585
R130 B.n429 B.n66 585
R131 B.n431 B.n430 585
R132 B.n432 B.n65 585
R133 B.n434 B.n433 585
R134 B.n435 B.n64 585
R135 B.n437 B.n436 585
R136 B.n438 B.n63 585
R137 B.n440 B.n439 585
R138 B.n441 B.n62 585
R139 B.n443 B.n442 585
R140 B.n444 B.n61 585
R141 B.n446 B.n445 585
R142 B.n447 B.n60 585
R143 B.n449 B.n448 585
R144 B.n450 B.n59 585
R145 B.n452 B.n451 585
R146 B.n453 B.n58 585
R147 B.n455 B.n454 585
R148 B.n456 B.n57 585
R149 B.n458 B.n457 585
R150 B.n459 B.n56 585
R151 B.n538 B.n537 585
R152 B.n536 B.n27 585
R153 B.n535 B.n534 585
R154 B.n533 B.n28 585
R155 B.n532 B.n531 585
R156 B.n530 B.n29 585
R157 B.n529 B.n528 585
R158 B.n527 B.n30 585
R159 B.n526 B.n525 585
R160 B.n524 B.n31 585
R161 B.n523 B.n522 585
R162 B.n521 B.n32 585
R163 B.n520 B.n519 585
R164 B.n518 B.n33 585
R165 B.n517 B.n516 585
R166 B.n515 B.n34 585
R167 B.n514 B.n513 585
R168 B.n512 B.n35 585
R169 B.n511 B.n510 585
R170 B.n509 B.n36 585
R171 B.n508 B.n507 585
R172 B.n505 B.n37 585
R173 B.n504 B.n503 585
R174 B.n502 B.n40 585
R175 B.n501 B.n500 585
R176 B.n499 B.n41 585
R177 B.n498 B.n497 585
R178 B.n496 B.n42 585
R179 B.n495 B.n494 585
R180 B.n493 B.n43 585
R181 B.n491 B.n490 585
R182 B.n489 B.n46 585
R183 B.n488 B.n487 585
R184 B.n486 B.n47 585
R185 B.n485 B.n484 585
R186 B.n483 B.n48 585
R187 B.n482 B.n481 585
R188 B.n480 B.n49 585
R189 B.n479 B.n478 585
R190 B.n477 B.n50 585
R191 B.n476 B.n475 585
R192 B.n474 B.n51 585
R193 B.n473 B.n472 585
R194 B.n471 B.n52 585
R195 B.n470 B.n469 585
R196 B.n468 B.n53 585
R197 B.n467 B.n466 585
R198 B.n465 B.n54 585
R199 B.n464 B.n463 585
R200 B.n462 B.n55 585
R201 B.n461 B.n460 585
R202 B.n539 B.n26 585
R203 B.n541 B.n540 585
R204 B.n542 B.n25 585
R205 B.n544 B.n543 585
R206 B.n545 B.n24 585
R207 B.n547 B.n546 585
R208 B.n548 B.n23 585
R209 B.n550 B.n549 585
R210 B.n551 B.n22 585
R211 B.n553 B.n552 585
R212 B.n554 B.n21 585
R213 B.n556 B.n555 585
R214 B.n557 B.n20 585
R215 B.n559 B.n558 585
R216 B.n560 B.n19 585
R217 B.n562 B.n561 585
R218 B.n563 B.n18 585
R219 B.n565 B.n564 585
R220 B.n566 B.n17 585
R221 B.n568 B.n567 585
R222 B.n569 B.n16 585
R223 B.n571 B.n570 585
R224 B.n572 B.n15 585
R225 B.n574 B.n573 585
R226 B.n575 B.n14 585
R227 B.n577 B.n576 585
R228 B.n578 B.n13 585
R229 B.n580 B.n579 585
R230 B.n581 B.n12 585
R231 B.n583 B.n582 585
R232 B.n584 B.n11 585
R233 B.n586 B.n585 585
R234 B.n587 B.n10 585
R235 B.n589 B.n588 585
R236 B.n590 B.n9 585
R237 B.n592 B.n591 585
R238 B.n593 B.n8 585
R239 B.n595 B.n594 585
R240 B.n596 B.n7 585
R241 B.n598 B.n597 585
R242 B.n599 B.n6 585
R243 B.n601 B.n600 585
R244 B.n602 B.n5 585
R245 B.n604 B.n603 585
R246 B.n605 B.n4 585
R247 B.n607 B.n606 585
R248 B.n608 B.n3 585
R249 B.n610 B.n609 585
R250 B.n611 B.n0 585
R251 B.n2 B.n1 585
R252 B.n158 B.n157 585
R253 B.n160 B.n159 585
R254 B.n161 B.n156 585
R255 B.n163 B.n162 585
R256 B.n164 B.n155 585
R257 B.n166 B.n165 585
R258 B.n167 B.n154 585
R259 B.n169 B.n168 585
R260 B.n170 B.n153 585
R261 B.n172 B.n171 585
R262 B.n173 B.n152 585
R263 B.n175 B.n174 585
R264 B.n176 B.n151 585
R265 B.n178 B.n177 585
R266 B.n179 B.n150 585
R267 B.n181 B.n180 585
R268 B.n182 B.n149 585
R269 B.n184 B.n183 585
R270 B.n185 B.n148 585
R271 B.n187 B.n186 585
R272 B.n188 B.n147 585
R273 B.n190 B.n189 585
R274 B.n191 B.n146 585
R275 B.n193 B.n192 585
R276 B.n194 B.n145 585
R277 B.n196 B.n195 585
R278 B.n197 B.n144 585
R279 B.n199 B.n198 585
R280 B.n200 B.n143 585
R281 B.n202 B.n201 585
R282 B.n203 B.n142 585
R283 B.n205 B.n204 585
R284 B.n206 B.n141 585
R285 B.n208 B.n207 585
R286 B.n209 B.n140 585
R287 B.n211 B.n210 585
R288 B.n212 B.n139 585
R289 B.n214 B.n213 585
R290 B.n215 B.n138 585
R291 B.n217 B.n216 585
R292 B.n218 B.n137 585
R293 B.n220 B.n219 585
R294 B.n221 B.n136 585
R295 B.n223 B.n222 585
R296 B.n224 B.n135 585
R297 B.n226 B.n225 585
R298 B.n227 B.n134 585
R299 B.n229 B.n228 585
R300 B.n228 B.n133 468.476
R301 B.n310 B.n309 468.476
R302 B.n460 B.n459 468.476
R303 B.n539 B.n538 468.476
R304 B.n613 B.n612 256.663
R305 B.n122 B.t9 255.651
R306 B.n274 B.t6 255.651
R307 B.n44 B.t0 255.651
R308 B.n38 B.t3 255.651
R309 B.n612 B.n611 235.042
R310 B.n612 B.n2 235.042
R311 B.n274 B.t7 171.671
R312 B.n44 B.t2 171.671
R313 B.n122 B.t10 171.666
R314 B.n38 B.t5 171.666
R315 B.n232 B.n133 163.367
R316 B.n233 B.n232 163.367
R317 B.n234 B.n233 163.367
R318 B.n234 B.n131 163.367
R319 B.n238 B.n131 163.367
R320 B.n239 B.n238 163.367
R321 B.n240 B.n239 163.367
R322 B.n240 B.n129 163.367
R323 B.n244 B.n129 163.367
R324 B.n245 B.n244 163.367
R325 B.n246 B.n245 163.367
R326 B.n246 B.n127 163.367
R327 B.n250 B.n127 163.367
R328 B.n251 B.n250 163.367
R329 B.n252 B.n251 163.367
R330 B.n252 B.n125 163.367
R331 B.n256 B.n125 163.367
R332 B.n257 B.n256 163.367
R333 B.n258 B.n257 163.367
R334 B.n258 B.n121 163.367
R335 B.n263 B.n121 163.367
R336 B.n264 B.n263 163.367
R337 B.n265 B.n264 163.367
R338 B.n265 B.n119 163.367
R339 B.n269 B.n119 163.367
R340 B.n270 B.n269 163.367
R341 B.n271 B.n270 163.367
R342 B.n271 B.n117 163.367
R343 B.n278 B.n117 163.367
R344 B.n279 B.n278 163.367
R345 B.n280 B.n279 163.367
R346 B.n280 B.n115 163.367
R347 B.n284 B.n115 163.367
R348 B.n285 B.n284 163.367
R349 B.n286 B.n285 163.367
R350 B.n286 B.n113 163.367
R351 B.n290 B.n113 163.367
R352 B.n291 B.n290 163.367
R353 B.n292 B.n291 163.367
R354 B.n292 B.n111 163.367
R355 B.n296 B.n111 163.367
R356 B.n297 B.n296 163.367
R357 B.n298 B.n297 163.367
R358 B.n298 B.n109 163.367
R359 B.n302 B.n109 163.367
R360 B.n303 B.n302 163.367
R361 B.n304 B.n303 163.367
R362 B.n304 B.n107 163.367
R363 B.n308 B.n107 163.367
R364 B.n309 B.n308 163.367
R365 B.n459 B.n458 163.367
R366 B.n458 B.n57 163.367
R367 B.n454 B.n57 163.367
R368 B.n454 B.n453 163.367
R369 B.n453 B.n452 163.367
R370 B.n452 B.n59 163.367
R371 B.n448 B.n59 163.367
R372 B.n448 B.n447 163.367
R373 B.n447 B.n446 163.367
R374 B.n446 B.n61 163.367
R375 B.n442 B.n61 163.367
R376 B.n442 B.n441 163.367
R377 B.n441 B.n440 163.367
R378 B.n440 B.n63 163.367
R379 B.n436 B.n63 163.367
R380 B.n436 B.n435 163.367
R381 B.n435 B.n434 163.367
R382 B.n434 B.n65 163.367
R383 B.n430 B.n65 163.367
R384 B.n430 B.n429 163.367
R385 B.n429 B.n428 163.367
R386 B.n428 B.n67 163.367
R387 B.n424 B.n67 163.367
R388 B.n424 B.n423 163.367
R389 B.n423 B.n422 163.367
R390 B.n422 B.n69 163.367
R391 B.n418 B.n69 163.367
R392 B.n418 B.n417 163.367
R393 B.n417 B.n416 163.367
R394 B.n416 B.n71 163.367
R395 B.n412 B.n71 163.367
R396 B.n412 B.n411 163.367
R397 B.n411 B.n410 163.367
R398 B.n410 B.n73 163.367
R399 B.n406 B.n73 163.367
R400 B.n406 B.n405 163.367
R401 B.n405 B.n404 163.367
R402 B.n404 B.n75 163.367
R403 B.n400 B.n75 163.367
R404 B.n400 B.n399 163.367
R405 B.n399 B.n398 163.367
R406 B.n398 B.n77 163.367
R407 B.n394 B.n77 163.367
R408 B.n394 B.n393 163.367
R409 B.n393 B.n392 163.367
R410 B.n392 B.n79 163.367
R411 B.n388 B.n79 163.367
R412 B.n388 B.n387 163.367
R413 B.n387 B.n386 163.367
R414 B.n386 B.n81 163.367
R415 B.n382 B.n81 163.367
R416 B.n382 B.n381 163.367
R417 B.n381 B.n380 163.367
R418 B.n380 B.n83 163.367
R419 B.n376 B.n83 163.367
R420 B.n376 B.n375 163.367
R421 B.n375 B.n374 163.367
R422 B.n374 B.n85 163.367
R423 B.n370 B.n85 163.367
R424 B.n370 B.n369 163.367
R425 B.n369 B.n368 163.367
R426 B.n368 B.n87 163.367
R427 B.n364 B.n87 163.367
R428 B.n364 B.n363 163.367
R429 B.n363 B.n362 163.367
R430 B.n362 B.n89 163.367
R431 B.n358 B.n89 163.367
R432 B.n358 B.n357 163.367
R433 B.n357 B.n356 163.367
R434 B.n356 B.n91 163.367
R435 B.n352 B.n91 163.367
R436 B.n352 B.n351 163.367
R437 B.n351 B.n350 163.367
R438 B.n350 B.n93 163.367
R439 B.n346 B.n93 163.367
R440 B.n346 B.n345 163.367
R441 B.n345 B.n344 163.367
R442 B.n344 B.n95 163.367
R443 B.n340 B.n95 163.367
R444 B.n340 B.n339 163.367
R445 B.n339 B.n338 163.367
R446 B.n338 B.n97 163.367
R447 B.n334 B.n97 163.367
R448 B.n334 B.n333 163.367
R449 B.n333 B.n332 163.367
R450 B.n332 B.n99 163.367
R451 B.n328 B.n99 163.367
R452 B.n328 B.n327 163.367
R453 B.n327 B.n326 163.367
R454 B.n326 B.n101 163.367
R455 B.n322 B.n101 163.367
R456 B.n322 B.n321 163.367
R457 B.n321 B.n320 163.367
R458 B.n320 B.n103 163.367
R459 B.n316 B.n103 163.367
R460 B.n316 B.n315 163.367
R461 B.n315 B.n314 163.367
R462 B.n314 B.n105 163.367
R463 B.n310 B.n105 163.367
R464 B.n538 B.n27 163.367
R465 B.n534 B.n27 163.367
R466 B.n534 B.n533 163.367
R467 B.n533 B.n532 163.367
R468 B.n532 B.n29 163.367
R469 B.n528 B.n29 163.367
R470 B.n528 B.n527 163.367
R471 B.n527 B.n526 163.367
R472 B.n526 B.n31 163.367
R473 B.n522 B.n31 163.367
R474 B.n522 B.n521 163.367
R475 B.n521 B.n520 163.367
R476 B.n520 B.n33 163.367
R477 B.n516 B.n33 163.367
R478 B.n516 B.n515 163.367
R479 B.n515 B.n514 163.367
R480 B.n514 B.n35 163.367
R481 B.n510 B.n35 163.367
R482 B.n510 B.n509 163.367
R483 B.n509 B.n508 163.367
R484 B.n508 B.n37 163.367
R485 B.n503 B.n37 163.367
R486 B.n503 B.n502 163.367
R487 B.n502 B.n501 163.367
R488 B.n501 B.n41 163.367
R489 B.n497 B.n41 163.367
R490 B.n497 B.n496 163.367
R491 B.n496 B.n495 163.367
R492 B.n495 B.n43 163.367
R493 B.n490 B.n43 163.367
R494 B.n490 B.n489 163.367
R495 B.n489 B.n488 163.367
R496 B.n488 B.n47 163.367
R497 B.n484 B.n47 163.367
R498 B.n484 B.n483 163.367
R499 B.n483 B.n482 163.367
R500 B.n482 B.n49 163.367
R501 B.n478 B.n49 163.367
R502 B.n478 B.n477 163.367
R503 B.n477 B.n476 163.367
R504 B.n476 B.n51 163.367
R505 B.n472 B.n51 163.367
R506 B.n472 B.n471 163.367
R507 B.n471 B.n470 163.367
R508 B.n470 B.n53 163.367
R509 B.n466 B.n53 163.367
R510 B.n466 B.n465 163.367
R511 B.n465 B.n464 163.367
R512 B.n464 B.n55 163.367
R513 B.n460 B.n55 163.367
R514 B.n540 B.n539 163.367
R515 B.n540 B.n25 163.367
R516 B.n544 B.n25 163.367
R517 B.n545 B.n544 163.367
R518 B.n546 B.n545 163.367
R519 B.n546 B.n23 163.367
R520 B.n550 B.n23 163.367
R521 B.n551 B.n550 163.367
R522 B.n552 B.n551 163.367
R523 B.n552 B.n21 163.367
R524 B.n556 B.n21 163.367
R525 B.n557 B.n556 163.367
R526 B.n558 B.n557 163.367
R527 B.n558 B.n19 163.367
R528 B.n562 B.n19 163.367
R529 B.n563 B.n562 163.367
R530 B.n564 B.n563 163.367
R531 B.n564 B.n17 163.367
R532 B.n568 B.n17 163.367
R533 B.n569 B.n568 163.367
R534 B.n570 B.n569 163.367
R535 B.n570 B.n15 163.367
R536 B.n574 B.n15 163.367
R537 B.n575 B.n574 163.367
R538 B.n576 B.n575 163.367
R539 B.n576 B.n13 163.367
R540 B.n580 B.n13 163.367
R541 B.n581 B.n580 163.367
R542 B.n582 B.n581 163.367
R543 B.n582 B.n11 163.367
R544 B.n586 B.n11 163.367
R545 B.n587 B.n586 163.367
R546 B.n588 B.n587 163.367
R547 B.n588 B.n9 163.367
R548 B.n592 B.n9 163.367
R549 B.n593 B.n592 163.367
R550 B.n594 B.n593 163.367
R551 B.n594 B.n7 163.367
R552 B.n598 B.n7 163.367
R553 B.n599 B.n598 163.367
R554 B.n600 B.n599 163.367
R555 B.n600 B.n5 163.367
R556 B.n604 B.n5 163.367
R557 B.n605 B.n604 163.367
R558 B.n606 B.n605 163.367
R559 B.n606 B.n3 163.367
R560 B.n610 B.n3 163.367
R561 B.n611 B.n610 163.367
R562 B.n157 B.n2 163.367
R563 B.n160 B.n157 163.367
R564 B.n161 B.n160 163.367
R565 B.n162 B.n161 163.367
R566 B.n162 B.n155 163.367
R567 B.n166 B.n155 163.367
R568 B.n167 B.n166 163.367
R569 B.n168 B.n167 163.367
R570 B.n168 B.n153 163.367
R571 B.n172 B.n153 163.367
R572 B.n173 B.n172 163.367
R573 B.n174 B.n173 163.367
R574 B.n174 B.n151 163.367
R575 B.n178 B.n151 163.367
R576 B.n179 B.n178 163.367
R577 B.n180 B.n179 163.367
R578 B.n180 B.n149 163.367
R579 B.n184 B.n149 163.367
R580 B.n185 B.n184 163.367
R581 B.n186 B.n185 163.367
R582 B.n186 B.n147 163.367
R583 B.n190 B.n147 163.367
R584 B.n191 B.n190 163.367
R585 B.n192 B.n191 163.367
R586 B.n192 B.n145 163.367
R587 B.n196 B.n145 163.367
R588 B.n197 B.n196 163.367
R589 B.n198 B.n197 163.367
R590 B.n198 B.n143 163.367
R591 B.n202 B.n143 163.367
R592 B.n203 B.n202 163.367
R593 B.n204 B.n203 163.367
R594 B.n204 B.n141 163.367
R595 B.n208 B.n141 163.367
R596 B.n209 B.n208 163.367
R597 B.n210 B.n209 163.367
R598 B.n210 B.n139 163.367
R599 B.n214 B.n139 163.367
R600 B.n215 B.n214 163.367
R601 B.n216 B.n215 163.367
R602 B.n216 B.n137 163.367
R603 B.n220 B.n137 163.367
R604 B.n221 B.n220 163.367
R605 B.n222 B.n221 163.367
R606 B.n222 B.n135 163.367
R607 B.n226 B.n135 163.367
R608 B.n227 B.n226 163.367
R609 B.n228 B.n227 163.367
R610 B.n275 B.t8 117.368
R611 B.n45 B.t1 117.368
R612 B.n123 B.t11 117.362
R613 B.n39 B.t4 117.362
R614 B.n261 B.n123 59.5399
R615 B.n276 B.n275 59.5399
R616 B.n492 B.n45 59.5399
R617 B.n506 B.n39 59.5399
R618 B.n123 B.n122 54.3035
R619 B.n275 B.n274 54.3035
R620 B.n45 B.n44 54.3035
R621 B.n39 B.n38 54.3035
R622 B.n537 B.n26 30.4395
R623 B.n461 B.n56 30.4395
R624 B.n230 B.n229 30.4395
R625 B.n311 B.n106 30.4395
R626 B B.n613 18.0485
R627 B.n541 B.n26 10.6151
R628 B.n542 B.n541 10.6151
R629 B.n543 B.n542 10.6151
R630 B.n543 B.n24 10.6151
R631 B.n547 B.n24 10.6151
R632 B.n548 B.n547 10.6151
R633 B.n549 B.n548 10.6151
R634 B.n549 B.n22 10.6151
R635 B.n553 B.n22 10.6151
R636 B.n554 B.n553 10.6151
R637 B.n555 B.n554 10.6151
R638 B.n555 B.n20 10.6151
R639 B.n559 B.n20 10.6151
R640 B.n560 B.n559 10.6151
R641 B.n561 B.n560 10.6151
R642 B.n561 B.n18 10.6151
R643 B.n565 B.n18 10.6151
R644 B.n566 B.n565 10.6151
R645 B.n567 B.n566 10.6151
R646 B.n567 B.n16 10.6151
R647 B.n571 B.n16 10.6151
R648 B.n572 B.n571 10.6151
R649 B.n573 B.n572 10.6151
R650 B.n573 B.n14 10.6151
R651 B.n577 B.n14 10.6151
R652 B.n578 B.n577 10.6151
R653 B.n579 B.n578 10.6151
R654 B.n579 B.n12 10.6151
R655 B.n583 B.n12 10.6151
R656 B.n584 B.n583 10.6151
R657 B.n585 B.n584 10.6151
R658 B.n585 B.n10 10.6151
R659 B.n589 B.n10 10.6151
R660 B.n590 B.n589 10.6151
R661 B.n591 B.n590 10.6151
R662 B.n591 B.n8 10.6151
R663 B.n595 B.n8 10.6151
R664 B.n596 B.n595 10.6151
R665 B.n597 B.n596 10.6151
R666 B.n597 B.n6 10.6151
R667 B.n601 B.n6 10.6151
R668 B.n602 B.n601 10.6151
R669 B.n603 B.n602 10.6151
R670 B.n603 B.n4 10.6151
R671 B.n607 B.n4 10.6151
R672 B.n608 B.n607 10.6151
R673 B.n609 B.n608 10.6151
R674 B.n609 B.n0 10.6151
R675 B.n537 B.n536 10.6151
R676 B.n536 B.n535 10.6151
R677 B.n535 B.n28 10.6151
R678 B.n531 B.n28 10.6151
R679 B.n531 B.n530 10.6151
R680 B.n530 B.n529 10.6151
R681 B.n529 B.n30 10.6151
R682 B.n525 B.n30 10.6151
R683 B.n525 B.n524 10.6151
R684 B.n524 B.n523 10.6151
R685 B.n523 B.n32 10.6151
R686 B.n519 B.n32 10.6151
R687 B.n519 B.n518 10.6151
R688 B.n518 B.n517 10.6151
R689 B.n517 B.n34 10.6151
R690 B.n513 B.n34 10.6151
R691 B.n513 B.n512 10.6151
R692 B.n512 B.n511 10.6151
R693 B.n511 B.n36 10.6151
R694 B.n507 B.n36 10.6151
R695 B.n505 B.n504 10.6151
R696 B.n504 B.n40 10.6151
R697 B.n500 B.n40 10.6151
R698 B.n500 B.n499 10.6151
R699 B.n499 B.n498 10.6151
R700 B.n498 B.n42 10.6151
R701 B.n494 B.n42 10.6151
R702 B.n494 B.n493 10.6151
R703 B.n491 B.n46 10.6151
R704 B.n487 B.n46 10.6151
R705 B.n487 B.n486 10.6151
R706 B.n486 B.n485 10.6151
R707 B.n485 B.n48 10.6151
R708 B.n481 B.n48 10.6151
R709 B.n481 B.n480 10.6151
R710 B.n480 B.n479 10.6151
R711 B.n479 B.n50 10.6151
R712 B.n475 B.n50 10.6151
R713 B.n475 B.n474 10.6151
R714 B.n474 B.n473 10.6151
R715 B.n473 B.n52 10.6151
R716 B.n469 B.n52 10.6151
R717 B.n469 B.n468 10.6151
R718 B.n468 B.n467 10.6151
R719 B.n467 B.n54 10.6151
R720 B.n463 B.n54 10.6151
R721 B.n463 B.n462 10.6151
R722 B.n462 B.n461 10.6151
R723 B.n457 B.n56 10.6151
R724 B.n457 B.n456 10.6151
R725 B.n456 B.n455 10.6151
R726 B.n455 B.n58 10.6151
R727 B.n451 B.n58 10.6151
R728 B.n451 B.n450 10.6151
R729 B.n450 B.n449 10.6151
R730 B.n449 B.n60 10.6151
R731 B.n445 B.n60 10.6151
R732 B.n445 B.n444 10.6151
R733 B.n444 B.n443 10.6151
R734 B.n443 B.n62 10.6151
R735 B.n439 B.n62 10.6151
R736 B.n439 B.n438 10.6151
R737 B.n438 B.n437 10.6151
R738 B.n437 B.n64 10.6151
R739 B.n433 B.n64 10.6151
R740 B.n433 B.n432 10.6151
R741 B.n432 B.n431 10.6151
R742 B.n431 B.n66 10.6151
R743 B.n427 B.n66 10.6151
R744 B.n427 B.n426 10.6151
R745 B.n426 B.n425 10.6151
R746 B.n425 B.n68 10.6151
R747 B.n421 B.n68 10.6151
R748 B.n421 B.n420 10.6151
R749 B.n420 B.n419 10.6151
R750 B.n419 B.n70 10.6151
R751 B.n415 B.n70 10.6151
R752 B.n415 B.n414 10.6151
R753 B.n414 B.n413 10.6151
R754 B.n413 B.n72 10.6151
R755 B.n409 B.n72 10.6151
R756 B.n409 B.n408 10.6151
R757 B.n408 B.n407 10.6151
R758 B.n407 B.n74 10.6151
R759 B.n403 B.n74 10.6151
R760 B.n403 B.n402 10.6151
R761 B.n402 B.n401 10.6151
R762 B.n401 B.n76 10.6151
R763 B.n397 B.n76 10.6151
R764 B.n397 B.n396 10.6151
R765 B.n396 B.n395 10.6151
R766 B.n395 B.n78 10.6151
R767 B.n391 B.n78 10.6151
R768 B.n391 B.n390 10.6151
R769 B.n390 B.n389 10.6151
R770 B.n389 B.n80 10.6151
R771 B.n385 B.n80 10.6151
R772 B.n385 B.n384 10.6151
R773 B.n384 B.n383 10.6151
R774 B.n383 B.n82 10.6151
R775 B.n379 B.n82 10.6151
R776 B.n379 B.n378 10.6151
R777 B.n378 B.n377 10.6151
R778 B.n377 B.n84 10.6151
R779 B.n373 B.n84 10.6151
R780 B.n373 B.n372 10.6151
R781 B.n372 B.n371 10.6151
R782 B.n371 B.n86 10.6151
R783 B.n367 B.n86 10.6151
R784 B.n367 B.n366 10.6151
R785 B.n366 B.n365 10.6151
R786 B.n365 B.n88 10.6151
R787 B.n361 B.n88 10.6151
R788 B.n361 B.n360 10.6151
R789 B.n360 B.n359 10.6151
R790 B.n359 B.n90 10.6151
R791 B.n355 B.n90 10.6151
R792 B.n355 B.n354 10.6151
R793 B.n354 B.n353 10.6151
R794 B.n353 B.n92 10.6151
R795 B.n349 B.n92 10.6151
R796 B.n349 B.n348 10.6151
R797 B.n348 B.n347 10.6151
R798 B.n347 B.n94 10.6151
R799 B.n343 B.n94 10.6151
R800 B.n343 B.n342 10.6151
R801 B.n342 B.n341 10.6151
R802 B.n341 B.n96 10.6151
R803 B.n337 B.n96 10.6151
R804 B.n337 B.n336 10.6151
R805 B.n336 B.n335 10.6151
R806 B.n335 B.n98 10.6151
R807 B.n331 B.n98 10.6151
R808 B.n331 B.n330 10.6151
R809 B.n330 B.n329 10.6151
R810 B.n329 B.n100 10.6151
R811 B.n325 B.n100 10.6151
R812 B.n325 B.n324 10.6151
R813 B.n324 B.n323 10.6151
R814 B.n323 B.n102 10.6151
R815 B.n319 B.n102 10.6151
R816 B.n319 B.n318 10.6151
R817 B.n318 B.n317 10.6151
R818 B.n317 B.n104 10.6151
R819 B.n313 B.n104 10.6151
R820 B.n313 B.n312 10.6151
R821 B.n312 B.n311 10.6151
R822 B.n158 B.n1 10.6151
R823 B.n159 B.n158 10.6151
R824 B.n159 B.n156 10.6151
R825 B.n163 B.n156 10.6151
R826 B.n164 B.n163 10.6151
R827 B.n165 B.n164 10.6151
R828 B.n165 B.n154 10.6151
R829 B.n169 B.n154 10.6151
R830 B.n170 B.n169 10.6151
R831 B.n171 B.n170 10.6151
R832 B.n171 B.n152 10.6151
R833 B.n175 B.n152 10.6151
R834 B.n176 B.n175 10.6151
R835 B.n177 B.n176 10.6151
R836 B.n177 B.n150 10.6151
R837 B.n181 B.n150 10.6151
R838 B.n182 B.n181 10.6151
R839 B.n183 B.n182 10.6151
R840 B.n183 B.n148 10.6151
R841 B.n187 B.n148 10.6151
R842 B.n188 B.n187 10.6151
R843 B.n189 B.n188 10.6151
R844 B.n189 B.n146 10.6151
R845 B.n193 B.n146 10.6151
R846 B.n194 B.n193 10.6151
R847 B.n195 B.n194 10.6151
R848 B.n195 B.n144 10.6151
R849 B.n199 B.n144 10.6151
R850 B.n200 B.n199 10.6151
R851 B.n201 B.n200 10.6151
R852 B.n201 B.n142 10.6151
R853 B.n205 B.n142 10.6151
R854 B.n206 B.n205 10.6151
R855 B.n207 B.n206 10.6151
R856 B.n207 B.n140 10.6151
R857 B.n211 B.n140 10.6151
R858 B.n212 B.n211 10.6151
R859 B.n213 B.n212 10.6151
R860 B.n213 B.n138 10.6151
R861 B.n217 B.n138 10.6151
R862 B.n218 B.n217 10.6151
R863 B.n219 B.n218 10.6151
R864 B.n219 B.n136 10.6151
R865 B.n223 B.n136 10.6151
R866 B.n224 B.n223 10.6151
R867 B.n225 B.n224 10.6151
R868 B.n225 B.n134 10.6151
R869 B.n229 B.n134 10.6151
R870 B.n231 B.n230 10.6151
R871 B.n231 B.n132 10.6151
R872 B.n235 B.n132 10.6151
R873 B.n236 B.n235 10.6151
R874 B.n237 B.n236 10.6151
R875 B.n237 B.n130 10.6151
R876 B.n241 B.n130 10.6151
R877 B.n242 B.n241 10.6151
R878 B.n243 B.n242 10.6151
R879 B.n243 B.n128 10.6151
R880 B.n247 B.n128 10.6151
R881 B.n248 B.n247 10.6151
R882 B.n249 B.n248 10.6151
R883 B.n249 B.n126 10.6151
R884 B.n253 B.n126 10.6151
R885 B.n254 B.n253 10.6151
R886 B.n255 B.n254 10.6151
R887 B.n255 B.n124 10.6151
R888 B.n259 B.n124 10.6151
R889 B.n260 B.n259 10.6151
R890 B.n262 B.n120 10.6151
R891 B.n266 B.n120 10.6151
R892 B.n267 B.n266 10.6151
R893 B.n268 B.n267 10.6151
R894 B.n268 B.n118 10.6151
R895 B.n272 B.n118 10.6151
R896 B.n273 B.n272 10.6151
R897 B.n277 B.n273 10.6151
R898 B.n281 B.n116 10.6151
R899 B.n282 B.n281 10.6151
R900 B.n283 B.n282 10.6151
R901 B.n283 B.n114 10.6151
R902 B.n287 B.n114 10.6151
R903 B.n288 B.n287 10.6151
R904 B.n289 B.n288 10.6151
R905 B.n289 B.n112 10.6151
R906 B.n293 B.n112 10.6151
R907 B.n294 B.n293 10.6151
R908 B.n295 B.n294 10.6151
R909 B.n295 B.n110 10.6151
R910 B.n299 B.n110 10.6151
R911 B.n300 B.n299 10.6151
R912 B.n301 B.n300 10.6151
R913 B.n301 B.n108 10.6151
R914 B.n305 B.n108 10.6151
R915 B.n306 B.n305 10.6151
R916 B.n307 B.n306 10.6151
R917 B.n307 B.n106 10.6151
R918 B.n613 B.n0 8.11757
R919 B.n613 B.n1 8.11757
R920 B.n506 B.n505 6.5566
R921 B.n493 B.n492 6.5566
R922 B.n262 B.n261 6.5566
R923 B.n277 B.n276 6.5566
R924 B.n507 B.n506 4.05904
R925 B.n492 B.n491 4.05904
R926 B.n261 B.n260 4.05904
R927 B.n276 B.n116 4.05904
R928 VN.n51 VN.n27 161.3
R929 VN.n50 VN.n49 161.3
R930 VN.n48 VN.n28 161.3
R931 VN.n47 VN.n46 161.3
R932 VN.n45 VN.n29 161.3
R933 VN.n44 VN.n43 161.3
R934 VN.n42 VN.n41 161.3
R935 VN.n40 VN.n31 161.3
R936 VN.n39 VN.n38 161.3
R937 VN.n37 VN.n32 161.3
R938 VN.n36 VN.n35 161.3
R939 VN.n24 VN.n0 161.3
R940 VN.n23 VN.n22 161.3
R941 VN.n21 VN.n1 161.3
R942 VN.n20 VN.n19 161.3
R943 VN.n18 VN.n2 161.3
R944 VN.n17 VN.n16 161.3
R945 VN.n15 VN.n14 161.3
R946 VN.n13 VN.n4 161.3
R947 VN.n12 VN.n11 161.3
R948 VN.n10 VN.n5 161.3
R949 VN.n9 VN.n8 161.3
R950 VN.n26 VN.n25 101.072
R951 VN.n53 VN.n52 101.072
R952 VN.n6 VN.t2 81.4408
R953 VN.n33 VN.t1 81.4408
R954 VN.n19 VN.n1 56.5617
R955 VN.n46 VN.n28 56.5617
R956 VN.n7 VN.n6 52.9956
R957 VN.n34 VN.n33 52.9956
R958 VN.n7 VN.t3 47.8102
R959 VN.n3 VN.t6 47.8102
R960 VN.n25 VN.t0 47.8102
R961 VN.n34 VN.t4 47.8102
R962 VN.n30 VN.t5 47.8102
R963 VN.n52 VN.t7 47.8102
R964 VN VN.n53 45.1724
R965 VN.n12 VN.n5 40.577
R966 VN.n13 VN.n12 40.577
R967 VN.n39 VN.n32 40.577
R968 VN.n40 VN.n39 40.577
R969 VN.n8 VN.n5 24.5923
R970 VN.n14 VN.n13 24.5923
R971 VN.n18 VN.n17 24.5923
R972 VN.n19 VN.n18 24.5923
R973 VN.n23 VN.n1 24.5923
R974 VN.n24 VN.n23 24.5923
R975 VN.n35 VN.n32 24.5923
R976 VN.n46 VN.n45 24.5923
R977 VN.n45 VN.n44 24.5923
R978 VN.n41 VN.n40 24.5923
R979 VN.n51 VN.n50 24.5923
R980 VN.n50 VN.n28 24.5923
R981 VN.n8 VN.n7 19.674
R982 VN.n14 VN.n3 19.674
R983 VN.n35 VN.n34 19.674
R984 VN.n41 VN.n30 19.674
R985 VN.n25 VN.n24 9.83723
R986 VN.n52 VN.n51 9.83723
R987 VN.n36 VN.n33 6.84375
R988 VN.n9 VN.n6 6.84375
R989 VN.n17 VN.n3 4.91887
R990 VN.n44 VN.n30 4.91887
R991 VN.n53 VN.n27 0.278335
R992 VN.n26 VN.n0 0.278335
R993 VN.n49 VN.n27 0.189894
R994 VN.n49 VN.n48 0.189894
R995 VN.n48 VN.n47 0.189894
R996 VN.n47 VN.n29 0.189894
R997 VN.n43 VN.n29 0.189894
R998 VN.n43 VN.n42 0.189894
R999 VN.n42 VN.n31 0.189894
R1000 VN.n38 VN.n31 0.189894
R1001 VN.n38 VN.n37 0.189894
R1002 VN.n37 VN.n36 0.189894
R1003 VN.n10 VN.n9 0.189894
R1004 VN.n11 VN.n10 0.189894
R1005 VN.n11 VN.n4 0.189894
R1006 VN.n15 VN.n4 0.189894
R1007 VN.n16 VN.n15 0.189894
R1008 VN.n16 VN.n2 0.189894
R1009 VN.n20 VN.n2 0.189894
R1010 VN.n21 VN.n20 0.189894
R1011 VN.n22 VN.n21 0.189894
R1012 VN.n22 VN.n0 0.189894
R1013 VN VN.n26 0.153485
R1014 VTAIL.n11 VTAIL.t2 90.0077
R1015 VTAIL.n10 VTAIL.t8 90.0077
R1016 VTAIL.n7 VTAIL.t13 90.0077
R1017 VTAIL.n15 VTAIL.t9 90.0076
R1018 VTAIL.n2 VTAIL.t10 90.0076
R1019 VTAIL.n3 VTAIL.t4 90.0076
R1020 VTAIL.n6 VTAIL.t5 90.0076
R1021 VTAIL.n14 VTAIL.t1 90.0076
R1022 VTAIL.n13 VTAIL.n12 83.3741
R1023 VTAIL.n9 VTAIL.n8 83.3741
R1024 VTAIL.n1 VTAIL.n0 83.3739
R1025 VTAIL.n5 VTAIL.n4 83.3739
R1026 VTAIL.n15 VTAIL.n14 19.0048
R1027 VTAIL.n7 VTAIL.n6 19.0048
R1028 VTAIL.n0 VTAIL.t12 6.63417
R1029 VTAIL.n0 VTAIL.t14 6.63417
R1030 VTAIL.n4 VTAIL.t0 6.63417
R1031 VTAIL.n4 VTAIL.t7 6.63417
R1032 VTAIL.n12 VTAIL.t3 6.63417
R1033 VTAIL.n12 VTAIL.t6 6.63417
R1034 VTAIL.n8 VTAIL.t11 6.63417
R1035 VTAIL.n8 VTAIL.t15 6.63417
R1036 VTAIL.n9 VTAIL.n7 2.41429
R1037 VTAIL.n10 VTAIL.n9 2.41429
R1038 VTAIL.n13 VTAIL.n11 2.41429
R1039 VTAIL.n14 VTAIL.n13 2.41429
R1040 VTAIL.n6 VTAIL.n5 2.41429
R1041 VTAIL.n5 VTAIL.n3 2.41429
R1042 VTAIL.n2 VTAIL.n1 2.41429
R1043 VTAIL VTAIL.n15 2.3561
R1044 VTAIL.n11 VTAIL.n10 0.470328
R1045 VTAIL.n3 VTAIL.n2 0.470328
R1046 VTAIL VTAIL.n1 0.0586897
R1047 VDD2.n2 VDD2.n1 101.204
R1048 VDD2.n2 VDD2.n0 101.204
R1049 VDD2 VDD2.n5 101.201
R1050 VDD2.n4 VDD2.n3 100.052
R1051 VDD2.n4 VDD2.n2 38.8015
R1052 VDD2.n5 VDD2.t3 6.63417
R1053 VDD2.n5 VDD2.t6 6.63417
R1054 VDD2.n3 VDD2.t0 6.63417
R1055 VDD2.n3 VDD2.t2 6.63417
R1056 VDD2.n1 VDD2.t1 6.63417
R1057 VDD2.n1 VDD2.t7 6.63417
R1058 VDD2.n0 VDD2.t5 6.63417
R1059 VDD2.n0 VDD2.t4 6.63417
R1060 VDD2 VDD2.n4 1.26559
R1061 VP.n19 VP.n18 161.3
R1062 VP.n20 VP.n15 161.3
R1063 VP.n22 VP.n21 161.3
R1064 VP.n23 VP.n14 161.3
R1065 VP.n25 VP.n24 161.3
R1066 VP.n27 VP.n26 161.3
R1067 VP.n28 VP.n12 161.3
R1068 VP.n30 VP.n29 161.3
R1069 VP.n31 VP.n11 161.3
R1070 VP.n33 VP.n32 161.3
R1071 VP.n34 VP.n10 161.3
R1072 VP.n64 VP.n0 161.3
R1073 VP.n63 VP.n62 161.3
R1074 VP.n61 VP.n1 161.3
R1075 VP.n60 VP.n59 161.3
R1076 VP.n58 VP.n2 161.3
R1077 VP.n57 VP.n56 161.3
R1078 VP.n55 VP.n54 161.3
R1079 VP.n53 VP.n4 161.3
R1080 VP.n52 VP.n51 161.3
R1081 VP.n50 VP.n5 161.3
R1082 VP.n49 VP.n48 161.3
R1083 VP.n46 VP.n6 161.3
R1084 VP.n45 VP.n44 161.3
R1085 VP.n43 VP.n7 161.3
R1086 VP.n42 VP.n41 161.3
R1087 VP.n40 VP.n8 161.3
R1088 VP.n39 VP.n38 161.3
R1089 VP.n37 VP.n9 101.072
R1090 VP.n66 VP.n65 101.072
R1091 VP.n36 VP.n35 101.072
R1092 VP.n16 VP.t3 81.4408
R1093 VP.n41 VP.n7 56.5617
R1094 VP.n59 VP.n1 56.5617
R1095 VP.n29 VP.n11 56.5617
R1096 VP.n17 VP.n16 52.9956
R1097 VP.n9 VP.t0 47.8102
R1098 VP.n47 VP.t5 47.8102
R1099 VP.n3 VP.t7 47.8102
R1100 VP.n65 VP.t1 47.8102
R1101 VP.n35 VP.t4 47.8102
R1102 VP.n13 VP.t6 47.8102
R1103 VP.n17 VP.t2 47.8102
R1104 VP.n37 VP.n36 44.8936
R1105 VP.n52 VP.n5 40.577
R1106 VP.n53 VP.n52 40.577
R1107 VP.n23 VP.n22 40.577
R1108 VP.n22 VP.n15 40.577
R1109 VP.n40 VP.n39 24.5923
R1110 VP.n41 VP.n40 24.5923
R1111 VP.n45 VP.n7 24.5923
R1112 VP.n46 VP.n45 24.5923
R1113 VP.n48 VP.n5 24.5923
R1114 VP.n54 VP.n53 24.5923
R1115 VP.n58 VP.n57 24.5923
R1116 VP.n59 VP.n58 24.5923
R1117 VP.n63 VP.n1 24.5923
R1118 VP.n64 VP.n63 24.5923
R1119 VP.n33 VP.n11 24.5923
R1120 VP.n34 VP.n33 24.5923
R1121 VP.n24 VP.n23 24.5923
R1122 VP.n28 VP.n27 24.5923
R1123 VP.n29 VP.n28 24.5923
R1124 VP.n18 VP.n15 24.5923
R1125 VP.n48 VP.n47 19.674
R1126 VP.n54 VP.n3 19.674
R1127 VP.n24 VP.n13 19.674
R1128 VP.n18 VP.n17 19.674
R1129 VP.n39 VP.n9 9.83723
R1130 VP.n65 VP.n64 9.83723
R1131 VP.n35 VP.n34 9.83723
R1132 VP.n19 VP.n16 6.84375
R1133 VP.n47 VP.n46 4.91887
R1134 VP.n57 VP.n3 4.91887
R1135 VP.n27 VP.n13 4.91887
R1136 VP.n36 VP.n10 0.278335
R1137 VP.n38 VP.n37 0.278335
R1138 VP.n66 VP.n0 0.278335
R1139 VP.n20 VP.n19 0.189894
R1140 VP.n21 VP.n20 0.189894
R1141 VP.n21 VP.n14 0.189894
R1142 VP.n25 VP.n14 0.189894
R1143 VP.n26 VP.n25 0.189894
R1144 VP.n26 VP.n12 0.189894
R1145 VP.n30 VP.n12 0.189894
R1146 VP.n31 VP.n30 0.189894
R1147 VP.n32 VP.n31 0.189894
R1148 VP.n32 VP.n10 0.189894
R1149 VP.n38 VP.n8 0.189894
R1150 VP.n42 VP.n8 0.189894
R1151 VP.n43 VP.n42 0.189894
R1152 VP.n44 VP.n43 0.189894
R1153 VP.n44 VP.n6 0.189894
R1154 VP.n49 VP.n6 0.189894
R1155 VP.n50 VP.n49 0.189894
R1156 VP.n51 VP.n50 0.189894
R1157 VP.n51 VP.n4 0.189894
R1158 VP.n55 VP.n4 0.189894
R1159 VP.n56 VP.n55 0.189894
R1160 VP.n56 VP.n2 0.189894
R1161 VP.n60 VP.n2 0.189894
R1162 VP.n61 VP.n60 0.189894
R1163 VP.n62 VP.n61 0.189894
R1164 VP.n62 VP.n0 0.189894
R1165 VP VP.n66 0.153485
R1166 VDD1 VDD1.n0 101.319
R1167 VDD1.n3 VDD1.n2 101.204
R1168 VDD1.n3 VDD1.n1 101.204
R1169 VDD1.n5 VDD1.n4 100.052
R1170 VDD1.n5 VDD1.n3 39.3845
R1171 VDD1.n4 VDD1.t1 6.63417
R1172 VDD1.n4 VDD1.t3 6.63417
R1173 VDD1.n0 VDD1.t4 6.63417
R1174 VDD1.n0 VDD1.t5 6.63417
R1175 VDD1.n2 VDD1.t0 6.63417
R1176 VDD1.n2 VDD1.t6 6.63417
R1177 VDD1.n1 VDD1.t7 6.63417
R1178 VDD1.n1 VDD1.t2 6.63417
R1179 VDD1 VDD1.n5 1.14921
C0 VP B 1.96488f
C1 VP VDD1 4.12853f
C2 w_n3770_n1948# B 7.93817f
C3 w_n3770_n1948# VDD1 1.72395f
C4 VP w_n3770_n1948# 7.99435f
C5 VN VTAIL 4.63033f
C6 VDD2 B 1.50918f
C7 VDD1 VDD2 1.71044f
C8 VP VDD2 0.510575f
C9 w_n3770_n1948# VDD2 1.8329f
C10 B VTAIL 2.58932f
C11 VDD1 VTAIL 5.60297f
C12 VN B 1.14585f
C13 VP VTAIL 4.64443f
C14 VN VDD1 0.155725f
C15 VN VP 6.18408f
C16 w_n3770_n1948# VTAIL 2.58077f
C17 VN w_n3770_n1948# 7.50539f
C18 VDD2 VTAIL 5.65652f
C19 VDD1 B 1.41715f
C20 VN VDD2 3.77564f
C21 VDD2 VSUBS 1.499312f
C22 VDD1 VSUBS 2.125295f
C23 VTAIL VSUBS 0.656855f
C24 VN VSUBS 6.27464f
C25 VP VSUBS 2.953087f
C26 B VSUBS 4.019731f
C27 w_n3770_n1948# VSUBS 92.0634f
C28 VDD1.t4 VSUBS 0.095628f
C29 VDD1.t5 VSUBS 0.095628f
C30 VDD1.n0 VSUBS 0.605071f
C31 VDD1.t7 VSUBS 0.095628f
C32 VDD1.t2 VSUBS 0.095628f
C33 VDD1.n1 VSUBS 0.60422f
C34 VDD1.t0 VSUBS 0.095628f
C35 VDD1.t6 VSUBS 0.095628f
C36 VDD1.n2 VSUBS 0.60422f
C37 VDD1.n3 VSUBS 3.13361f
C38 VDD1.t1 VSUBS 0.095628f
C39 VDD1.t3 VSUBS 0.095628f
C40 VDD1.n4 VSUBS 0.596592f
C41 VDD1.n5 VSUBS 2.5288f
C42 VP.n0 VSUBS 0.054717f
C43 VP.t1 VSUBS 1.312f
C44 VP.n1 VSUBS 0.054592f
C45 VP.n2 VSUBS 0.041505f
C46 VP.t7 VSUBS 1.312f
C47 VP.n3 VSUBS 0.507253f
C48 VP.n4 VSUBS 0.041505f
C49 VP.n5 VSUBS 0.082056f
C50 VP.n6 VSUBS 0.041505f
C51 VP.t5 VSUBS 1.312f
C52 VP.n7 VSUBS 0.066075f
C53 VP.n8 VSUBS 0.041505f
C54 VP.t0 VSUBS 1.312f
C55 VP.n9 VSUBS 0.637874f
C56 VP.n10 VSUBS 0.054717f
C57 VP.t4 VSUBS 1.312f
C58 VP.n11 VSUBS 0.054592f
C59 VP.n12 VSUBS 0.041505f
C60 VP.t6 VSUBS 1.312f
C61 VP.n13 VSUBS 0.507253f
C62 VP.n14 VSUBS 0.041505f
C63 VP.n15 VSUBS 0.082056f
C64 VP.t3 VSUBS 1.62328f
C65 VP.n16 VSUBS 0.597502f
C66 VP.t2 VSUBS 1.312f
C67 VP.n17 VSUBS 0.635251f
C68 VP.n18 VSUBS 0.069367f
C69 VP.n19 VSUBS 0.395675f
C70 VP.n20 VSUBS 0.041505f
C71 VP.n21 VSUBS 0.041505f
C72 VP.n22 VSUBS 0.033522f
C73 VP.n23 VSUBS 0.082056f
C74 VP.n24 VSUBS 0.069367f
C75 VP.n25 VSUBS 0.041505f
C76 VP.n26 VSUBS 0.041505f
C77 VP.n27 VSUBS 0.04657f
C78 VP.n28 VSUBS 0.076967f
C79 VP.n29 VSUBS 0.066075f
C80 VP.n30 VSUBS 0.041505f
C81 VP.n31 VSUBS 0.041505f
C82 VP.n32 VSUBS 0.041505f
C83 VP.n33 VSUBS 0.076967f
C84 VP.n34 VSUBS 0.054169f
C85 VP.n35 VSUBS 0.637874f
C86 VP.n36 VSUBS 1.96053f
C87 VP.n37 VSUBS 1.99386f
C88 VP.n38 VSUBS 0.054717f
C89 VP.n39 VSUBS 0.054169f
C90 VP.n40 VSUBS 0.076967f
C91 VP.n41 VSUBS 0.054592f
C92 VP.n42 VSUBS 0.041505f
C93 VP.n43 VSUBS 0.041505f
C94 VP.n44 VSUBS 0.041505f
C95 VP.n45 VSUBS 0.076967f
C96 VP.n46 VSUBS 0.04657f
C97 VP.n47 VSUBS 0.507253f
C98 VP.n48 VSUBS 0.069367f
C99 VP.n49 VSUBS 0.041505f
C100 VP.n50 VSUBS 0.041505f
C101 VP.n51 VSUBS 0.041505f
C102 VP.n52 VSUBS 0.033522f
C103 VP.n53 VSUBS 0.082056f
C104 VP.n54 VSUBS 0.069367f
C105 VP.n55 VSUBS 0.041505f
C106 VP.n56 VSUBS 0.041505f
C107 VP.n57 VSUBS 0.04657f
C108 VP.n58 VSUBS 0.076967f
C109 VP.n59 VSUBS 0.066075f
C110 VP.n60 VSUBS 0.041505f
C111 VP.n61 VSUBS 0.041505f
C112 VP.n62 VSUBS 0.041505f
C113 VP.n63 VSUBS 0.076967f
C114 VP.n64 VSUBS 0.054169f
C115 VP.n65 VSUBS 0.637874f
C116 VP.n66 VSUBS 0.06602f
C117 VDD2.t5 VSUBS 0.094545f
C118 VDD2.t4 VSUBS 0.094545f
C119 VDD2.n0 VSUBS 0.597379f
C120 VDD2.t1 VSUBS 0.094545f
C121 VDD2.t7 VSUBS 0.094545f
C122 VDD2.n1 VSUBS 0.597379f
C123 VDD2.n2 VSUBS 3.04701f
C124 VDD2.t0 VSUBS 0.094545f
C125 VDD2.t2 VSUBS 0.094545f
C126 VDD2.n3 VSUBS 0.58984f
C127 VDD2.n4 VSUBS 2.47026f
C128 VDD2.t3 VSUBS 0.094545f
C129 VDD2.t6 VSUBS 0.094545f
C130 VDD2.n5 VSUBS 0.597352f
C131 VTAIL.t12 VSUBS 0.118159f
C132 VTAIL.t14 VSUBS 0.118159f
C133 VTAIL.n0 VSUBS 0.645341f
C134 VTAIL.n1 VSUBS 0.758193f
C135 VTAIL.t10 VSUBS 0.904988f
C136 VTAIL.n2 VSUBS 0.861274f
C137 VTAIL.t4 VSUBS 0.904988f
C138 VTAIL.n3 VSUBS 0.861274f
C139 VTAIL.t0 VSUBS 0.118159f
C140 VTAIL.t7 VSUBS 0.118159f
C141 VTAIL.n4 VSUBS 0.645341f
C142 VTAIL.n5 VSUBS 0.989813f
C143 VTAIL.t5 VSUBS 0.904988f
C144 VTAIL.n6 VSUBS 1.88228f
C145 VTAIL.t13 VSUBS 0.904993f
C146 VTAIL.n7 VSUBS 1.88227f
C147 VTAIL.t11 VSUBS 0.118159f
C148 VTAIL.t15 VSUBS 0.118159f
C149 VTAIL.n8 VSUBS 0.645345f
C150 VTAIL.n9 VSUBS 0.989809f
C151 VTAIL.t8 VSUBS 0.904993f
C152 VTAIL.n10 VSUBS 0.861269f
C153 VTAIL.t2 VSUBS 0.904993f
C154 VTAIL.n11 VSUBS 0.861269f
C155 VTAIL.t3 VSUBS 0.118159f
C156 VTAIL.t6 VSUBS 0.118159f
C157 VTAIL.n12 VSUBS 0.645345f
C158 VTAIL.n13 VSUBS 0.989809f
C159 VTAIL.t1 VSUBS 0.904988f
C160 VTAIL.n14 VSUBS 1.88228f
C161 VTAIL.t9 VSUBS 0.904988f
C162 VTAIL.n15 VSUBS 1.87656f
C163 VN.n0 VSUBS 0.052671f
C164 VN.t0 VSUBS 1.26295f
C165 VN.n1 VSUBS 0.052551f
C166 VN.n2 VSUBS 0.039953f
C167 VN.t6 VSUBS 1.26295f
C168 VN.n3 VSUBS 0.488288f
C169 VN.n4 VSUBS 0.039953f
C170 VN.n5 VSUBS 0.078988f
C171 VN.t2 VSUBS 1.56259f
C172 VN.n6 VSUBS 0.575163f
C173 VN.t3 VSUBS 1.26295f
C174 VN.n7 VSUBS 0.611501f
C175 VN.n8 VSUBS 0.066774f
C176 VN.n9 VSUBS 0.380881f
C177 VN.n10 VSUBS 0.039953f
C178 VN.n11 VSUBS 0.039953f
C179 VN.n12 VSUBS 0.032269f
C180 VN.n13 VSUBS 0.078988f
C181 VN.n14 VSUBS 0.066774f
C182 VN.n15 VSUBS 0.039953f
C183 VN.n16 VSUBS 0.039953f
C184 VN.n17 VSUBS 0.044828f
C185 VN.n18 VSUBS 0.074089f
C186 VN.n19 VSUBS 0.063605f
C187 VN.n20 VSUBS 0.039953f
C188 VN.n21 VSUBS 0.039953f
C189 VN.n22 VSUBS 0.039953f
C190 VN.n23 VSUBS 0.074089f
C191 VN.n24 VSUBS 0.052144f
C192 VN.n25 VSUBS 0.614026f
C193 VN.n26 VSUBS 0.063551f
C194 VN.n27 VSUBS 0.052671f
C195 VN.t7 VSUBS 1.26295f
C196 VN.n28 VSUBS 0.052551f
C197 VN.n29 VSUBS 0.039953f
C198 VN.t5 VSUBS 1.26295f
C199 VN.n30 VSUBS 0.488288f
C200 VN.n31 VSUBS 0.039953f
C201 VN.n32 VSUBS 0.078988f
C202 VN.t1 VSUBS 1.56259f
C203 VN.n33 VSUBS 0.575163f
C204 VN.t4 VSUBS 1.26295f
C205 VN.n34 VSUBS 0.611501f
C206 VN.n35 VSUBS 0.066774f
C207 VN.n36 VSUBS 0.380881f
C208 VN.n37 VSUBS 0.039953f
C209 VN.n38 VSUBS 0.039953f
C210 VN.n39 VSUBS 0.032269f
C211 VN.n40 VSUBS 0.078988f
C212 VN.n41 VSUBS 0.066774f
C213 VN.n42 VSUBS 0.039953f
C214 VN.n43 VSUBS 0.039953f
C215 VN.n44 VSUBS 0.044828f
C216 VN.n45 VSUBS 0.074089f
C217 VN.n46 VSUBS 0.063605f
C218 VN.n47 VSUBS 0.039953f
C219 VN.n48 VSUBS 0.039953f
C220 VN.n49 VSUBS 0.039953f
C221 VN.n50 VSUBS 0.074089f
C222 VN.n51 VSUBS 0.052144f
C223 VN.n52 VSUBS 0.614026f
C224 VN.n53 VSUBS 1.90908f
C225 B.n0 VSUBS 0.007558f
C226 B.n1 VSUBS 0.007558f
C227 B.n2 VSUBS 0.011178f
C228 B.n3 VSUBS 0.008566f
C229 B.n4 VSUBS 0.008566f
C230 B.n5 VSUBS 0.008566f
C231 B.n6 VSUBS 0.008566f
C232 B.n7 VSUBS 0.008566f
C233 B.n8 VSUBS 0.008566f
C234 B.n9 VSUBS 0.008566f
C235 B.n10 VSUBS 0.008566f
C236 B.n11 VSUBS 0.008566f
C237 B.n12 VSUBS 0.008566f
C238 B.n13 VSUBS 0.008566f
C239 B.n14 VSUBS 0.008566f
C240 B.n15 VSUBS 0.008566f
C241 B.n16 VSUBS 0.008566f
C242 B.n17 VSUBS 0.008566f
C243 B.n18 VSUBS 0.008566f
C244 B.n19 VSUBS 0.008566f
C245 B.n20 VSUBS 0.008566f
C246 B.n21 VSUBS 0.008566f
C247 B.n22 VSUBS 0.008566f
C248 B.n23 VSUBS 0.008566f
C249 B.n24 VSUBS 0.008566f
C250 B.n25 VSUBS 0.008566f
C251 B.n26 VSUBS 0.018843f
C252 B.n27 VSUBS 0.008566f
C253 B.n28 VSUBS 0.008566f
C254 B.n29 VSUBS 0.008566f
C255 B.n30 VSUBS 0.008566f
C256 B.n31 VSUBS 0.008566f
C257 B.n32 VSUBS 0.008566f
C258 B.n33 VSUBS 0.008566f
C259 B.n34 VSUBS 0.008566f
C260 B.n35 VSUBS 0.008566f
C261 B.n36 VSUBS 0.008566f
C262 B.n37 VSUBS 0.008566f
C263 B.t4 VSUBS 0.16663f
C264 B.t5 VSUBS 0.18965f
C265 B.t3 VSUBS 0.705258f
C266 B.n38 VSUBS 0.123287f
C267 B.n39 VSUBS 0.084988f
C268 B.n40 VSUBS 0.008566f
C269 B.n41 VSUBS 0.008566f
C270 B.n42 VSUBS 0.008566f
C271 B.n43 VSUBS 0.008566f
C272 B.t1 VSUBS 0.16663f
C273 B.t2 VSUBS 0.189649f
C274 B.t0 VSUBS 0.705258f
C275 B.n44 VSUBS 0.123288f
C276 B.n45 VSUBS 0.084988f
C277 B.n46 VSUBS 0.008566f
C278 B.n47 VSUBS 0.008566f
C279 B.n48 VSUBS 0.008566f
C280 B.n49 VSUBS 0.008566f
C281 B.n50 VSUBS 0.008566f
C282 B.n51 VSUBS 0.008566f
C283 B.n52 VSUBS 0.008566f
C284 B.n53 VSUBS 0.008566f
C285 B.n54 VSUBS 0.008566f
C286 B.n55 VSUBS 0.008566f
C287 B.n56 VSUBS 0.018843f
C288 B.n57 VSUBS 0.008566f
C289 B.n58 VSUBS 0.008566f
C290 B.n59 VSUBS 0.008566f
C291 B.n60 VSUBS 0.008566f
C292 B.n61 VSUBS 0.008566f
C293 B.n62 VSUBS 0.008566f
C294 B.n63 VSUBS 0.008566f
C295 B.n64 VSUBS 0.008566f
C296 B.n65 VSUBS 0.008566f
C297 B.n66 VSUBS 0.008566f
C298 B.n67 VSUBS 0.008566f
C299 B.n68 VSUBS 0.008566f
C300 B.n69 VSUBS 0.008566f
C301 B.n70 VSUBS 0.008566f
C302 B.n71 VSUBS 0.008566f
C303 B.n72 VSUBS 0.008566f
C304 B.n73 VSUBS 0.008566f
C305 B.n74 VSUBS 0.008566f
C306 B.n75 VSUBS 0.008566f
C307 B.n76 VSUBS 0.008566f
C308 B.n77 VSUBS 0.008566f
C309 B.n78 VSUBS 0.008566f
C310 B.n79 VSUBS 0.008566f
C311 B.n80 VSUBS 0.008566f
C312 B.n81 VSUBS 0.008566f
C313 B.n82 VSUBS 0.008566f
C314 B.n83 VSUBS 0.008566f
C315 B.n84 VSUBS 0.008566f
C316 B.n85 VSUBS 0.008566f
C317 B.n86 VSUBS 0.008566f
C318 B.n87 VSUBS 0.008566f
C319 B.n88 VSUBS 0.008566f
C320 B.n89 VSUBS 0.008566f
C321 B.n90 VSUBS 0.008566f
C322 B.n91 VSUBS 0.008566f
C323 B.n92 VSUBS 0.008566f
C324 B.n93 VSUBS 0.008566f
C325 B.n94 VSUBS 0.008566f
C326 B.n95 VSUBS 0.008566f
C327 B.n96 VSUBS 0.008566f
C328 B.n97 VSUBS 0.008566f
C329 B.n98 VSUBS 0.008566f
C330 B.n99 VSUBS 0.008566f
C331 B.n100 VSUBS 0.008566f
C332 B.n101 VSUBS 0.008566f
C333 B.n102 VSUBS 0.008566f
C334 B.n103 VSUBS 0.008566f
C335 B.n104 VSUBS 0.008566f
C336 B.n105 VSUBS 0.008566f
C337 B.n106 VSUBS 0.018366f
C338 B.n107 VSUBS 0.008566f
C339 B.n108 VSUBS 0.008566f
C340 B.n109 VSUBS 0.008566f
C341 B.n110 VSUBS 0.008566f
C342 B.n111 VSUBS 0.008566f
C343 B.n112 VSUBS 0.008566f
C344 B.n113 VSUBS 0.008566f
C345 B.n114 VSUBS 0.008566f
C346 B.n115 VSUBS 0.008566f
C347 B.n116 VSUBS 0.005921f
C348 B.n117 VSUBS 0.008566f
C349 B.n118 VSUBS 0.008566f
C350 B.n119 VSUBS 0.008566f
C351 B.n120 VSUBS 0.008566f
C352 B.n121 VSUBS 0.008566f
C353 B.t11 VSUBS 0.16663f
C354 B.t10 VSUBS 0.18965f
C355 B.t9 VSUBS 0.705258f
C356 B.n122 VSUBS 0.123287f
C357 B.n123 VSUBS 0.084988f
C358 B.n124 VSUBS 0.008566f
C359 B.n125 VSUBS 0.008566f
C360 B.n126 VSUBS 0.008566f
C361 B.n127 VSUBS 0.008566f
C362 B.n128 VSUBS 0.008566f
C363 B.n129 VSUBS 0.008566f
C364 B.n130 VSUBS 0.008566f
C365 B.n131 VSUBS 0.008566f
C366 B.n132 VSUBS 0.008566f
C367 B.n133 VSUBS 0.019452f
C368 B.n134 VSUBS 0.008566f
C369 B.n135 VSUBS 0.008566f
C370 B.n136 VSUBS 0.008566f
C371 B.n137 VSUBS 0.008566f
C372 B.n138 VSUBS 0.008566f
C373 B.n139 VSUBS 0.008566f
C374 B.n140 VSUBS 0.008566f
C375 B.n141 VSUBS 0.008566f
C376 B.n142 VSUBS 0.008566f
C377 B.n143 VSUBS 0.008566f
C378 B.n144 VSUBS 0.008566f
C379 B.n145 VSUBS 0.008566f
C380 B.n146 VSUBS 0.008566f
C381 B.n147 VSUBS 0.008566f
C382 B.n148 VSUBS 0.008566f
C383 B.n149 VSUBS 0.008566f
C384 B.n150 VSUBS 0.008566f
C385 B.n151 VSUBS 0.008566f
C386 B.n152 VSUBS 0.008566f
C387 B.n153 VSUBS 0.008566f
C388 B.n154 VSUBS 0.008566f
C389 B.n155 VSUBS 0.008566f
C390 B.n156 VSUBS 0.008566f
C391 B.n157 VSUBS 0.008566f
C392 B.n158 VSUBS 0.008566f
C393 B.n159 VSUBS 0.008566f
C394 B.n160 VSUBS 0.008566f
C395 B.n161 VSUBS 0.008566f
C396 B.n162 VSUBS 0.008566f
C397 B.n163 VSUBS 0.008566f
C398 B.n164 VSUBS 0.008566f
C399 B.n165 VSUBS 0.008566f
C400 B.n166 VSUBS 0.008566f
C401 B.n167 VSUBS 0.008566f
C402 B.n168 VSUBS 0.008566f
C403 B.n169 VSUBS 0.008566f
C404 B.n170 VSUBS 0.008566f
C405 B.n171 VSUBS 0.008566f
C406 B.n172 VSUBS 0.008566f
C407 B.n173 VSUBS 0.008566f
C408 B.n174 VSUBS 0.008566f
C409 B.n175 VSUBS 0.008566f
C410 B.n176 VSUBS 0.008566f
C411 B.n177 VSUBS 0.008566f
C412 B.n178 VSUBS 0.008566f
C413 B.n179 VSUBS 0.008566f
C414 B.n180 VSUBS 0.008566f
C415 B.n181 VSUBS 0.008566f
C416 B.n182 VSUBS 0.008566f
C417 B.n183 VSUBS 0.008566f
C418 B.n184 VSUBS 0.008566f
C419 B.n185 VSUBS 0.008566f
C420 B.n186 VSUBS 0.008566f
C421 B.n187 VSUBS 0.008566f
C422 B.n188 VSUBS 0.008566f
C423 B.n189 VSUBS 0.008566f
C424 B.n190 VSUBS 0.008566f
C425 B.n191 VSUBS 0.008566f
C426 B.n192 VSUBS 0.008566f
C427 B.n193 VSUBS 0.008566f
C428 B.n194 VSUBS 0.008566f
C429 B.n195 VSUBS 0.008566f
C430 B.n196 VSUBS 0.008566f
C431 B.n197 VSUBS 0.008566f
C432 B.n198 VSUBS 0.008566f
C433 B.n199 VSUBS 0.008566f
C434 B.n200 VSUBS 0.008566f
C435 B.n201 VSUBS 0.008566f
C436 B.n202 VSUBS 0.008566f
C437 B.n203 VSUBS 0.008566f
C438 B.n204 VSUBS 0.008566f
C439 B.n205 VSUBS 0.008566f
C440 B.n206 VSUBS 0.008566f
C441 B.n207 VSUBS 0.008566f
C442 B.n208 VSUBS 0.008566f
C443 B.n209 VSUBS 0.008566f
C444 B.n210 VSUBS 0.008566f
C445 B.n211 VSUBS 0.008566f
C446 B.n212 VSUBS 0.008566f
C447 B.n213 VSUBS 0.008566f
C448 B.n214 VSUBS 0.008566f
C449 B.n215 VSUBS 0.008566f
C450 B.n216 VSUBS 0.008566f
C451 B.n217 VSUBS 0.008566f
C452 B.n218 VSUBS 0.008566f
C453 B.n219 VSUBS 0.008566f
C454 B.n220 VSUBS 0.008566f
C455 B.n221 VSUBS 0.008566f
C456 B.n222 VSUBS 0.008566f
C457 B.n223 VSUBS 0.008566f
C458 B.n224 VSUBS 0.008566f
C459 B.n225 VSUBS 0.008566f
C460 B.n226 VSUBS 0.008566f
C461 B.n227 VSUBS 0.008566f
C462 B.n228 VSUBS 0.018843f
C463 B.n229 VSUBS 0.018843f
C464 B.n230 VSUBS 0.019452f
C465 B.n231 VSUBS 0.008566f
C466 B.n232 VSUBS 0.008566f
C467 B.n233 VSUBS 0.008566f
C468 B.n234 VSUBS 0.008566f
C469 B.n235 VSUBS 0.008566f
C470 B.n236 VSUBS 0.008566f
C471 B.n237 VSUBS 0.008566f
C472 B.n238 VSUBS 0.008566f
C473 B.n239 VSUBS 0.008566f
C474 B.n240 VSUBS 0.008566f
C475 B.n241 VSUBS 0.008566f
C476 B.n242 VSUBS 0.008566f
C477 B.n243 VSUBS 0.008566f
C478 B.n244 VSUBS 0.008566f
C479 B.n245 VSUBS 0.008566f
C480 B.n246 VSUBS 0.008566f
C481 B.n247 VSUBS 0.008566f
C482 B.n248 VSUBS 0.008566f
C483 B.n249 VSUBS 0.008566f
C484 B.n250 VSUBS 0.008566f
C485 B.n251 VSUBS 0.008566f
C486 B.n252 VSUBS 0.008566f
C487 B.n253 VSUBS 0.008566f
C488 B.n254 VSUBS 0.008566f
C489 B.n255 VSUBS 0.008566f
C490 B.n256 VSUBS 0.008566f
C491 B.n257 VSUBS 0.008566f
C492 B.n258 VSUBS 0.008566f
C493 B.n259 VSUBS 0.008566f
C494 B.n260 VSUBS 0.005921f
C495 B.n261 VSUBS 0.019846f
C496 B.n262 VSUBS 0.006928f
C497 B.n263 VSUBS 0.008566f
C498 B.n264 VSUBS 0.008566f
C499 B.n265 VSUBS 0.008566f
C500 B.n266 VSUBS 0.008566f
C501 B.n267 VSUBS 0.008566f
C502 B.n268 VSUBS 0.008566f
C503 B.n269 VSUBS 0.008566f
C504 B.n270 VSUBS 0.008566f
C505 B.n271 VSUBS 0.008566f
C506 B.n272 VSUBS 0.008566f
C507 B.n273 VSUBS 0.008566f
C508 B.t8 VSUBS 0.16663f
C509 B.t7 VSUBS 0.189649f
C510 B.t6 VSUBS 0.705258f
C511 B.n274 VSUBS 0.123288f
C512 B.n275 VSUBS 0.084988f
C513 B.n276 VSUBS 0.019846f
C514 B.n277 VSUBS 0.006928f
C515 B.n278 VSUBS 0.008566f
C516 B.n279 VSUBS 0.008566f
C517 B.n280 VSUBS 0.008566f
C518 B.n281 VSUBS 0.008566f
C519 B.n282 VSUBS 0.008566f
C520 B.n283 VSUBS 0.008566f
C521 B.n284 VSUBS 0.008566f
C522 B.n285 VSUBS 0.008566f
C523 B.n286 VSUBS 0.008566f
C524 B.n287 VSUBS 0.008566f
C525 B.n288 VSUBS 0.008566f
C526 B.n289 VSUBS 0.008566f
C527 B.n290 VSUBS 0.008566f
C528 B.n291 VSUBS 0.008566f
C529 B.n292 VSUBS 0.008566f
C530 B.n293 VSUBS 0.008566f
C531 B.n294 VSUBS 0.008566f
C532 B.n295 VSUBS 0.008566f
C533 B.n296 VSUBS 0.008566f
C534 B.n297 VSUBS 0.008566f
C535 B.n298 VSUBS 0.008566f
C536 B.n299 VSUBS 0.008566f
C537 B.n300 VSUBS 0.008566f
C538 B.n301 VSUBS 0.008566f
C539 B.n302 VSUBS 0.008566f
C540 B.n303 VSUBS 0.008566f
C541 B.n304 VSUBS 0.008566f
C542 B.n305 VSUBS 0.008566f
C543 B.n306 VSUBS 0.008566f
C544 B.n307 VSUBS 0.008566f
C545 B.n308 VSUBS 0.008566f
C546 B.n309 VSUBS 0.019452f
C547 B.n310 VSUBS 0.018843f
C548 B.n311 VSUBS 0.019929f
C549 B.n312 VSUBS 0.008566f
C550 B.n313 VSUBS 0.008566f
C551 B.n314 VSUBS 0.008566f
C552 B.n315 VSUBS 0.008566f
C553 B.n316 VSUBS 0.008566f
C554 B.n317 VSUBS 0.008566f
C555 B.n318 VSUBS 0.008566f
C556 B.n319 VSUBS 0.008566f
C557 B.n320 VSUBS 0.008566f
C558 B.n321 VSUBS 0.008566f
C559 B.n322 VSUBS 0.008566f
C560 B.n323 VSUBS 0.008566f
C561 B.n324 VSUBS 0.008566f
C562 B.n325 VSUBS 0.008566f
C563 B.n326 VSUBS 0.008566f
C564 B.n327 VSUBS 0.008566f
C565 B.n328 VSUBS 0.008566f
C566 B.n329 VSUBS 0.008566f
C567 B.n330 VSUBS 0.008566f
C568 B.n331 VSUBS 0.008566f
C569 B.n332 VSUBS 0.008566f
C570 B.n333 VSUBS 0.008566f
C571 B.n334 VSUBS 0.008566f
C572 B.n335 VSUBS 0.008566f
C573 B.n336 VSUBS 0.008566f
C574 B.n337 VSUBS 0.008566f
C575 B.n338 VSUBS 0.008566f
C576 B.n339 VSUBS 0.008566f
C577 B.n340 VSUBS 0.008566f
C578 B.n341 VSUBS 0.008566f
C579 B.n342 VSUBS 0.008566f
C580 B.n343 VSUBS 0.008566f
C581 B.n344 VSUBS 0.008566f
C582 B.n345 VSUBS 0.008566f
C583 B.n346 VSUBS 0.008566f
C584 B.n347 VSUBS 0.008566f
C585 B.n348 VSUBS 0.008566f
C586 B.n349 VSUBS 0.008566f
C587 B.n350 VSUBS 0.008566f
C588 B.n351 VSUBS 0.008566f
C589 B.n352 VSUBS 0.008566f
C590 B.n353 VSUBS 0.008566f
C591 B.n354 VSUBS 0.008566f
C592 B.n355 VSUBS 0.008566f
C593 B.n356 VSUBS 0.008566f
C594 B.n357 VSUBS 0.008566f
C595 B.n358 VSUBS 0.008566f
C596 B.n359 VSUBS 0.008566f
C597 B.n360 VSUBS 0.008566f
C598 B.n361 VSUBS 0.008566f
C599 B.n362 VSUBS 0.008566f
C600 B.n363 VSUBS 0.008566f
C601 B.n364 VSUBS 0.008566f
C602 B.n365 VSUBS 0.008566f
C603 B.n366 VSUBS 0.008566f
C604 B.n367 VSUBS 0.008566f
C605 B.n368 VSUBS 0.008566f
C606 B.n369 VSUBS 0.008566f
C607 B.n370 VSUBS 0.008566f
C608 B.n371 VSUBS 0.008566f
C609 B.n372 VSUBS 0.008566f
C610 B.n373 VSUBS 0.008566f
C611 B.n374 VSUBS 0.008566f
C612 B.n375 VSUBS 0.008566f
C613 B.n376 VSUBS 0.008566f
C614 B.n377 VSUBS 0.008566f
C615 B.n378 VSUBS 0.008566f
C616 B.n379 VSUBS 0.008566f
C617 B.n380 VSUBS 0.008566f
C618 B.n381 VSUBS 0.008566f
C619 B.n382 VSUBS 0.008566f
C620 B.n383 VSUBS 0.008566f
C621 B.n384 VSUBS 0.008566f
C622 B.n385 VSUBS 0.008566f
C623 B.n386 VSUBS 0.008566f
C624 B.n387 VSUBS 0.008566f
C625 B.n388 VSUBS 0.008566f
C626 B.n389 VSUBS 0.008566f
C627 B.n390 VSUBS 0.008566f
C628 B.n391 VSUBS 0.008566f
C629 B.n392 VSUBS 0.008566f
C630 B.n393 VSUBS 0.008566f
C631 B.n394 VSUBS 0.008566f
C632 B.n395 VSUBS 0.008566f
C633 B.n396 VSUBS 0.008566f
C634 B.n397 VSUBS 0.008566f
C635 B.n398 VSUBS 0.008566f
C636 B.n399 VSUBS 0.008566f
C637 B.n400 VSUBS 0.008566f
C638 B.n401 VSUBS 0.008566f
C639 B.n402 VSUBS 0.008566f
C640 B.n403 VSUBS 0.008566f
C641 B.n404 VSUBS 0.008566f
C642 B.n405 VSUBS 0.008566f
C643 B.n406 VSUBS 0.008566f
C644 B.n407 VSUBS 0.008566f
C645 B.n408 VSUBS 0.008566f
C646 B.n409 VSUBS 0.008566f
C647 B.n410 VSUBS 0.008566f
C648 B.n411 VSUBS 0.008566f
C649 B.n412 VSUBS 0.008566f
C650 B.n413 VSUBS 0.008566f
C651 B.n414 VSUBS 0.008566f
C652 B.n415 VSUBS 0.008566f
C653 B.n416 VSUBS 0.008566f
C654 B.n417 VSUBS 0.008566f
C655 B.n418 VSUBS 0.008566f
C656 B.n419 VSUBS 0.008566f
C657 B.n420 VSUBS 0.008566f
C658 B.n421 VSUBS 0.008566f
C659 B.n422 VSUBS 0.008566f
C660 B.n423 VSUBS 0.008566f
C661 B.n424 VSUBS 0.008566f
C662 B.n425 VSUBS 0.008566f
C663 B.n426 VSUBS 0.008566f
C664 B.n427 VSUBS 0.008566f
C665 B.n428 VSUBS 0.008566f
C666 B.n429 VSUBS 0.008566f
C667 B.n430 VSUBS 0.008566f
C668 B.n431 VSUBS 0.008566f
C669 B.n432 VSUBS 0.008566f
C670 B.n433 VSUBS 0.008566f
C671 B.n434 VSUBS 0.008566f
C672 B.n435 VSUBS 0.008566f
C673 B.n436 VSUBS 0.008566f
C674 B.n437 VSUBS 0.008566f
C675 B.n438 VSUBS 0.008566f
C676 B.n439 VSUBS 0.008566f
C677 B.n440 VSUBS 0.008566f
C678 B.n441 VSUBS 0.008566f
C679 B.n442 VSUBS 0.008566f
C680 B.n443 VSUBS 0.008566f
C681 B.n444 VSUBS 0.008566f
C682 B.n445 VSUBS 0.008566f
C683 B.n446 VSUBS 0.008566f
C684 B.n447 VSUBS 0.008566f
C685 B.n448 VSUBS 0.008566f
C686 B.n449 VSUBS 0.008566f
C687 B.n450 VSUBS 0.008566f
C688 B.n451 VSUBS 0.008566f
C689 B.n452 VSUBS 0.008566f
C690 B.n453 VSUBS 0.008566f
C691 B.n454 VSUBS 0.008566f
C692 B.n455 VSUBS 0.008566f
C693 B.n456 VSUBS 0.008566f
C694 B.n457 VSUBS 0.008566f
C695 B.n458 VSUBS 0.008566f
C696 B.n459 VSUBS 0.018843f
C697 B.n460 VSUBS 0.019452f
C698 B.n461 VSUBS 0.019452f
C699 B.n462 VSUBS 0.008566f
C700 B.n463 VSUBS 0.008566f
C701 B.n464 VSUBS 0.008566f
C702 B.n465 VSUBS 0.008566f
C703 B.n466 VSUBS 0.008566f
C704 B.n467 VSUBS 0.008566f
C705 B.n468 VSUBS 0.008566f
C706 B.n469 VSUBS 0.008566f
C707 B.n470 VSUBS 0.008566f
C708 B.n471 VSUBS 0.008566f
C709 B.n472 VSUBS 0.008566f
C710 B.n473 VSUBS 0.008566f
C711 B.n474 VSUBS 0.008566f
C712 B.n475 VSUBS 0.008566f
C713 B.n476 VSUBS 0.008566f
C714 B.n477 VSUBS 0.008566f
C715 B.n478 VSUBS 0.008566f
C716 B.n479 VSUBS 0.008566f
C717 B.n480 VSUBS 0.008566f
C718 B.n481 VSUBS 0.008566f
C719 B.n482 VSUBS 0.008566f
C720 B.n483 VSUBS 0.008566f
C721 B.n484 VSUBS 0.008566f
C722 B.n485 VSUBS 0.008566f
C723 B.n486 VSUBS 0.008566f
C724 B.n487 VSUBS 0.008566f
C725 B.n488 VSUBS 0.008566f
C726 B.n489 VSUBS 0.008566f
C727 B.n490 VSUBS 0.008566f
C728 B.n491 VSUBS 0.005921f
C729 B.n492 VSUBS 0.019846f
C730 B.n493 VSUBS 0.006928f
C731 B.n494 VSUBS 0.008566f
C732 B.n495 VSUBS 0.008566f
C733 B.n496 VSUBS 0.008566f
C734 B.n497 VSUBS 0.008566f
C735 B.n498 VSUBS 0.008566f
C736 B.n499 VSUBS 0.008566f
C737 B.n500 VSUBS 0.008566f
C738 B.n501 VSUBS 0.008566f
C739 B.n502 VSUBS 0.008566f
C740 B.n503 VSUBS 0.008566f
C741 B.n504 VSUBS 0.008566f
C742 B.n505 VSUBS 0.006928f
C743 B.n506 VSUBS 0.019846f
C744 B.n507 VSUBS 0.005921f
C745 B.n508 VSUBS 0.008566f
C746 B.n509 VSUBS 0.008566f
C747 B.n510 VSUBS 0.008566f
C748 B.n511 VSUBS 0.008566f
C749 B.n512 VSUBS 0.008566f
C750 B.n513 VSUBS 0.008566f
C751 B.n514 VSUBS 0.008566f
C752 B.n515 VSUBS 0.008566f
C753 B.n516 VSUBS 0.008566f
C754 B.n517 VSUBS 0.008566f
C755 B.n518 VSUBS 0.008566f
C756 B.n519 VSUBS 0.008566f
C757 B.n520 VSUBS 0.008566f
C758 B.n521 VSUBS 0.008566f
C759 B.n522 VSUBS 0.008566f
C760 B.n523 VSUBS 0.008566f
C761 B.n524 VSUBS 0.008566f
C762 B.n525 VSUBS 0.008566f
C763 B.n526 VSUBS 0.008566f
C764 B.n527 VSUBS 0.008566f
C765 B.n528 VSUBS 0.008566f
C766 B.n529 VSUBS 0.008566f
C767 B.n530 VSUBS 0.008566f
C768 B.n531 VSUBS 0.008566f
C769 B.n532 VSUBS 0.008566f
C770 B.n533 VSUBS 0.008566f
C771 B.n534 VSUBS 0.008566f
C772 B.n535 VSUBS 0.008566f
C773 B.n536 VSUBS 0.008566f
C774 B.n537 VSUBS 0.019452f
C775 B.n538 VSUBS 0.019452f
C776 B.n539 VSUBS 0.018843f
C777 B.n540 VSUBS 0.008566f
C778 B.n541 VSUBS 0.008566f
C779 B.n542 VSUBS 0.008566f
C780 B.n543 VSUBS 0.008566f
C781 B.n544 VSUBS 0.008566f
C782 B.n545 VSUBS 0.008566f
C783 B.n546 VSUBS 0.008566f
C784 B.n547 VSUBS 0.008566f
C785 B.n548 VSUBS 0.008566f
C786 B.n549 VSUBS 0.008566f
C787 B.n550 VSUBS 0.008566f
C788 B.n551 VSUBS 0.008566f
C789 B.n552 VSUBS 0.008566f
C790 B.n553 VSUBS 0.008566f
C791 B.n554 VSUBS 0.008566f
C792 B.n555 VSUBS 0.008566f
C793 B.n556 VSUBS 0.008566f
C794 B.n557 VSUBS 0.008566f
C795 B.n558 VSUBS 0.008566f
C796 B.n559 VSUBS 0.008566f
C797 B.n560 VSUBS 0.008566f
C798 B.n561 VSUBS 0.008566f
C799 B.n562 VSUBS 0.008566f
C800 B.n563 VSUBS 0.008566f
C801 B.n564 VSUBS 0.008566f
C802 B.n565 VSUBS 0.008566f
C803 B.n566 VSUBS 0.008566f
C804 B.n567 VSUBS 0.008566f
C805 B.n568 VSUBS 0.008566f
C806 B.n569 VSUBS 0.008566f
C807 B.n570 VSUBS 0.008566f
C808 B.n571 VSUBS 0.008566f
C809 B.n572 VSUBS 0.008566f
C810 B.n573 VSUBS 0.008566f
C811 B.n574 VSUBS 0.008566f
C812 B.n575 VSUBS 0.008566f
C813 B.n576 VSUBS 0.008566f
C814 B.n577 VSUBS 0.008566f
C815 B.n578 VSUBS 0.008566f
C816 B.n579 VSUBS 0.008566f
C817 B.n580 VSUBS 0.008566f
C818 B.n581 VSUBS 0.008566f
C819 B.n582 VSUBS 0.008566f
C820 B.n583 VSUBS 0.008566f
C821 B.n584 VSUBS 0.008566f
C822 B.n585 VSUBS 0.008566f
C823 B.n586 VSUBS 0.008566f
C824 B.n587 VSUBS 0.008566f
C825 B.n588 VSUBS 0.008566f
C826 B.n589 VSUBS 0.008566f
C827 B.n590 VSUBS 0.008566f
C828 B.n591 VSUBS 0.008566f
C829 B.n592 VSUBS 0.008566f
C830 B.n593 VSUBS 0.008566f
C831 B.n594 VSUBS 0.008566f
C832 B.n595 VSUBS 0.008566f
C833 B.n596 VSUBS 0.008566f
C834 B.n597 VSUBS 0.008566f
C835 B.n598 VSUBS 0.008566f
C836 B.n599 VSUBS 0.008566f
C837 B.n600 VSUBS 0.008566f
C838 B.n601 VSUBS 0.008566f
C839 B.n602 VSUBS 0.008566f
C840 B.n603 VSUBS 0.008566f
C841 B.n604 VSUBS 0.008566f
C842 B.n605 VSUBS 0.008566f
C843 B.n606 VSUBS 0.008566f
C844 B.n607 VSUBS 0.008566f
C845 B.n608 VSUBS 0.008566f
C846 B.n609 VSUBS 0.008566f
C847 B.n610 VSUBS 0.008566f
C848 B.n611 VSUBS 0.011178f
C849 B.n612 VSUBS 0.011908f
C850 B.n613 VSUBS 0.023679f
.ends

