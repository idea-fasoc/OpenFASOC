* NGSPICE file created from diff_pair_sample_0259.ext - technology: sky130A

.subckt diff_pair_sample_0259 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=0.12705 pd=1.1 as=0.12705 ps=1.1 w=0.77 l=1.87
X1 VDD1.t9 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.12705 pd=1.1 as=0.12705 ps=1.1 w=0.77 l=1.87
X2 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.32 as=0 ps=0 w=0.77 l=1.87
X3 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.32 as=0 ps=0 w=0.77 l=1.87
X4 VDD2.t5 VN.t1 VTAIL.t18 B.t5 sky130_fd_pr__nfet_01v8 ad=0.12705 pd=1.1 as=0.3003 ps=2.32 w=0.77 l=1.87
X5 VDD1.t8 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.12705 pd=1.1 as=0.12705 ps=1.1 w=0.77 l=1.87
X6 VTAIL.t9 VP.t2 VDD1.t7 B.t9 sky130_fd_pr__nfet_01v8 ad=0.12705 pd=1.1 as=0.12705 ps=1.1 w=0.77 l=1.87
X7 VTAIL.t17 VN.t2 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.12705 pd=1.1 as=0.12705 ps=1.1 w=0.77 l=1.87
X8 VDD2.t8 VN.t3 VTAIL.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.32 as=0.12705 ps=1.1 w=0.77 l=1.87
X9 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.32 as=0 ps=0 w=0.77 l=1.87
X10 VTAIL.t15 VN.t4 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.12705 pd=1.1 as=0.12705 ps=1.1 w=0.77 l=1.87
X11 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.32 as=0 ps=0 w=0.77 l=1.87
X12 VDD2.t9 VN.t5 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=0.12705 pd=1.1 as=0.12705 ps=1.1 w=0.77 l=1.87
X13 VDD1.t6 VP.t3 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.32 as=0.12705 ps=1.1 w=0.77 l=1.87
X14 VDD2.t1 VN.t6 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=0.12705 pd=1.1 as=0.12705 ps=1.1 w=0.77 l=1.87
X15 VTAIL.t3 VP.t4 VDD1.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=0.12705 pd=1.1 as=0.12705 ps=1.1 w=0.77 l=1.87
X16 VTAIL.t2 VP.t5 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.12705 pd=1.1 as=0.12705 ps=1.1 w=0.77 l=1.87
X17 VTAIL.t12 VN.t7 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.12705 pd=1.1 as=0.12705 ps=1.1 w=0.77 l=1.87
X18 VDD2.t7 VN.t8 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=0.12705 pd=1.1 as=0.3003 ps=2.32 w=0.77 l=1.87
X19 VDD1.t3 VP.t6 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.12705 pd=1.1 as=0.3003 ps=2.32 w=0.77 l=1.87
X20 VDD1.t2 VP.t7 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.32 as=0.12705 ps=1.1 w=0.77 l=1.87
X21 VDD2.t0 VN.t9 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=0.3003 pd=2.32 as=0.12705 ps=1.1 w=0.77 l=1.87
X22 VDD1.t1 VP.t8 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.12705 pd=1.1 as=0.3003 ps=2.32 w=0.77 l=1.87
X23 VTAIL.t4 VP.t9 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=0.12705 pd=1.1 as=0.12705 ps=1.1 w=0.77 l=1.87
R0 VN.n59 VN.n31 161.3
R1 VN.n58 VN.n57 161.3
R2 VN.n56 VN.n32 161.3
R3 VN.n55 VN.n54 161.3
R4 VN.n52 VN.n33 161.3
R5 VN.n51 VN.n50 161.3
R6 VN.n49 VN.n34 161.3
R7 VN.n48 VN.n47 161.3
R8 VN.n46 VN.n35 161.3
R9 VN.n45 VN.n44 161.3
R10 VN.n43 VN.n36 161.3
R11 VN.n42 VN.n41 161.3
R12 VN.n40 VN.n37 161.3
R13 VN.n28 VN.n0 161.3
R14 VN.n27 VN.n26 161.3
R15 VN.n25 VN.n1 161.3
R16 VN.n24 VN.n23 161.3
R17 VN.n21 VN.n2 161.3
R18 VN.n20 VN.n19 161.3
R19 VN.n18 VN.n3 161.3
R20 VN.n17 VN.n16 161.3
R21 VN.n15 VN.n4 161.3
R22 VN.n14 VN.n13 161.3
R23 VN.n12 VN.n5 161.3
R24 VN.n11 VN.n10 161.3
R25 VN.n9 VN.n6 161.3
R26 VN.n30 VN.n29 91.1828
R27 VN.n61 VN.n60 91.1828
R28 VN.n8 VN.n7 59.9592
R29 VN.n39 VN.n38 59.9592
R30 VN.n27 VN.n1 56.5193
R31 VN.n58 VN.n32 56.5193
R32 VN.n10 VN.n5 50.2061
R33 VN.n20 VN.n3 50.2061
R34 VN.n41 VN.n36 50.2061
R35 VN.n51 VN.n34 50.2061
R36 VN VN.n61 40.9072
R37 VN.n7 VN.t9 40.1933
R38 VN.n38 VN.t8 40.1933
R39 VN.n14 VN.n5 30.7807
R40 VN.n16 VN.n3 30.7807
R41 VN.n45 VN.n36 30.7807
R42 VN.n47 VN.n34 30.7807
R43 VN.n10 VN.n9 24.4675
R44 VN.n15 VN.n14 24.4675
R45 VN.n16 VN.n15 24.4675
R46 VN.n21 VN.n20 24.4675
R47 VN.n23 VN.n1 24.4675
R48 VN.n28 VN.n27 24.4675
R49 VN.n41 VN.n40 24.4675
R50 VN.n47 VN.n46 24.4675
R51 VN.n46 VN.n45 24.4675
R52 VN.n54 VN.n32 24.4675
R53 VN.n52 VN.n51 24.4675
R54 VN.n59 VN.n58 24.4675
R55 VN.n29 VN.n28 19.5741
R56 VN.n60 VN.n59 19.5741
R57 VN.n23 VN.n22 14.6807
R58 VN.n54 VN.n53 14.6807
R59 VN.n38 VN.n37 13.3649
R60 VN.n7 VN.n6 13.3649
R61 VN.n15 VN.t5 9.92403
R62 VN.n8 VN.t7 9.92403
R63 VN.n22 VN.t0 9.92403
R64 VN.n29 VN.t1 9.92403
R65 VN.n46 VN.t6 9.92403
R66 VN.n39 VN.t4 9.92403
R67 VN.n53 VN.t2 9.92403
R68 VN.n60 VN.t3 9.92403
R69 VN.n9 VN.n8 9.7873
R70 VN.n22 VN.n21 9.7873
R71 VN.n40 VN.n39 9.7873
R72 VN.n53 VN.n52 9.7873
R73 VN.n61 VN.n31 0.278367
R74 VN.n30 VN.n0 0.278367
R75 VN.n57 VN.n31 0.189894
R76 VN.n57 VN.n56 0.189894
R77 VN.n56 VN.n55 0.189894
R78 VN.n55 VN.n33 0.189894
R79 VN.n50 VN.n33 0.189894
R80 VN.n50 VN.n49 0.189894
R81 VN.n49 VN.n48 0.189894
R82 VN.n48 VN.n35 0.189894
R83 VN.n44 VN.n35 0.189894
R84 VN.n44 VN.n43 0.189894
R85 VN.n43 VN.n42 0.189894
R86 VN.n42 VN.n37 0.189894
R87 VN.n11 VN.n6 0.189894
R88 VN.n12 VN.n11 0.189894
R89 VN.n13 VN.n12 0.189894
R90 VN.n13 VN.n4 0.189894
R91 VN.n17 VN.n4 0.189894
R92 VN.n18 VN.n17 0.189894
R93 VN.n19 VN.n18 0.189894
R94 VN.n19 VN.n2 0.189894
R95 VN.n24 VN.n2 0.189894
R96 VN.n25 VN.n24 0.189894
R97 VN.n26 VN.n25 0.189894
R98 VN.n26 VN.n0 0.189894
R99 VN VN.n30 0.153454
R100 VDD2.n1 VDD2.t0 264.772
R101 VDD2.n4 VDD2.t8 262.875
R102 VDD2.n3 VDD2.n2 238.529
R103 VDD2 VDD2.n7 238.525
R104 VDD2.n6 VDD2.n5 237.161
R105 VDD2.n1 VDD2.n0 237.161
R106 VDD2.n4 VDD2.n3 33.3877
R107 VDD2.n7 VDD2.t3 25.7148
R108 VDD2.n7 VDD2.t7 25.7148
R109 VDD2.n5 VDD2.t4 25.7148
R110 VDD2.n5 VDD2.t1 25.7148
R111 VDD2.n2 VDD2.t6 25.7148
R112 VDD2.n2 VDD2.t5 25.7148
R113 VDD2.n0 VDD2.t2 25.7148
R114 VDD2.n0 VDD2.t9 25.7148
R115 VDD2.n6 VDD2.n4 1.89705
R116 VDD2 VDD2.n6 0.532828
R117 VDD2.n3 VDD2.n1 0.419292
R118 VTAIL.n17 VTAIL.t18 246.196
R119 VTAIL.n2 VTAIL.t7 246.196
R120 VTAIL.n16 VTAIL.t5 246.196
R121 VTAIL.n11 VTAIL.t11 246.196
R122 VTAIL.n19 VTAIL.n18 220.482
R123 VTAIL.n1 VTAIL.n0 220.482
R124 VTAIL.n4 VTAIL.n3 220.482
R125 VTAIL.n6 VTAIL.n5 220.482
R126 VTAIL.n15 VTAIL.n14 220.482
R127 VTAIL.n13 VTAIL.n12 220.482
R128 VTAIL.n10 VTAIL.n9 220.482
R129 VTAIL.n8 VTAIL.n7 220.482
R130 VTAIL.n18 VTAIL.t14 25.7148
R131 VTAIL.n18 VTAIL.t19 25.7148
R132 VTAIL.n0 VTAIL.t10 25.7148
R133 VTAIL.n0 VTAIL.t12 25.7148
R134 VTAIL.n3 VTAIL.t0 25.7148
R135 VTAIL.n3 VTAIL.t3 25.7148
R136 VTAIL.n5 VTAIL.t8 25.7148
R137 VTAIL.n5 VTAIL.t4 25.7148
R138 VTAIL.n14 VTAIL.t1 25.7148
R139 VTAIL.n14 VTAIL.t9 25.7148
R140 VTAIL.n12 VTAIL.t6 25.7148
R141 VTAIL.n12 VTAIL.t2 25.7148
R142 VTAIL.n9 VTAIL.t13 25.7148
R143 VTAIL.n9 VTAIL.t15 25.7148
R144 VTAIL.n7 VTAIL.t16 25.7148
R145 VTAIL.n7 VTAIL.t17 25.7148
R146 VTAIL.n8 VTAIL.n6 16.8238
R147 VTAIL.n17 VTAIL.n16 14.9272
R148 VTAIL.n10 VTAIL.n8 1.89705
R149 VTAIL.n11 VTAIL.n10 1.89705
R150 VTAIL.n15 VTAIL.n13 1.89705
R151 VTAIL.n16 VTAIL.n15 1.89705
R152 VTAIL.n6 VTAIL.n4 1.89705
R153 VTAIL.n4 VTAIL.n2 1.89705
R154 VTAIL.n19 VTAIL.n17 1.89705
R155 VTAIL VTAIL.n1 1.4811
R156 VTAIL.n13 VTAIL.n11 1.4186
R157 VTAIL.n2 VTAIL.n1 1.4186
R158 VTAIL VTAIL.n19 0.416448
R159 B.n522 B.n521 585
R160 B.n523 B.n522 585
R161 B.n155 B.n101 585
R162 B.n154 B.n153 585
R163 B.n152 B.n151 585
R164 B.n150 B.n149 585
R165 B.n148 B.n147 585
R166 B.n146 B.n145 585
R167 B.n144 B.n143 585
R168 B.n142 B.n141 585
R169 B.n140 B.n139 585
R170 B.n138 B.n137 585
R171 B.n136 B.n135 585
R172 B.n134 B.n133 585
R173 B.n132 B.n131 585
R174 B.n130 B.n129 585
R175 B.n128 B.n127 585
R176 B.n126 B.n125 585
R177 B.n124 B.n123 585
R178 B.n121 B.n120 585
R179 B.n119 B.n118 585
R180 B.n117 B.n116 585
R181 B.n115 B.n114 585
R182 B.n113 B.n112 585
R183 B.n111 B.n110 585
R184 B.n109 B.n108 585
R185 B.n88 B.n87 585
R186 B.n526 B.n525 585
R187 B.n520 B.n102 585
R188 B.n102 B.n85 585
R189 B.n519 B.n84 585
R190 B.n530 B.n84 585
R191 B.n518 B.n83 585
R192 B.n531 B.n83 585
R193 B.n517 B.n82 585
R194 B.n532 B.n82 585
R195 B.n516 B.n515 585
R196 B.n515 B.n78 585
R197 B.n514 B.n77 585
R198 B.n538 B.n77 585
R199 B.n513 B.n76 585
R200 B.n539 B.n76 585
R201 B.n512 B.n75 585
R202 B.n540 B.n75 585
R203 B.n511 B.n510 585
R204 B.n510 B.n71 585
R205 B.n509 B.n70 585
R206 B.n546 B.n70 585
R207 B.n508 B.n69 585
R208 B.n547 B.n69 585
R209 B.n507 B.n68 585
R210 B.n548 B.n68 585
R211 B.n506 B.n505 585
R212 B.n505 B.n64 585
R213 B.n504 B.n63 585
R214 B.n554 B.n63 585
R215 B.n503 B.n62 585
R216 B.n555 B.n62 585
R217 B.n502 B.n61 585
R218 B.n556 B.n61 585
R219 B.n501 B.n500 585
R220 B.n500 B.n60 585
R221 B.n499 B.n56 585
R222 B.n562 B.n56 585
R223 B.n498 B.n55 585
R224 B.n563 B.n55 585
R225 B.n497 B.n54 585
R226 B.n564 B.n54 585
R227 B.n496 B.n495 585
R228 B.n495 B.n50 585
R229 B.n494 B.n49 585
R230 B.n570 B.n49 585
R231 B.n493 B.n48 585
R232 B.n571 B.n48 585
R233 B.n492 B.n47 585
R234 B.n572 B.n47 585
R235 B.n491 B.n490 585
R236 B.n490 B.n43 585
R237 B.n489 B.n42 585
R238 B.n578 B.n42 585
R239 B.n488 B.n41 585
R240 B.n579 B.n41 585
R241 B.n487 B.n40 585
R242 B.n580 B.n40 585
R243 B.n486 B.n485 585
R244 B.n485 B.n36 585
R245 B.n484 B.n35 585
R246 B.n586 B.n35 585
R247 B.n483 B.n34 585
R248 B.n587 B.n34 585
R249 B.n482 B.n33 585
R250 B.n588 B.n33 585
R251 B.n481 B.n480 585
R252 B.n480 B.n29 585
R253 B.n479 B.n28 585
R254 B.n594 B.n28 585
R255 B.n478 B.n27 585
R256 B.n595 B.n27 585
R257 B.n477 B.n26 585
R258 B.n596 B.n26 585
R259 B.n476 B.n475 585
R260 B.n475 B.n22 585
R261 B.n474 B.n21 585
R262 B.n602 B.n21 585
R263 B.n473 B.n20 585
R264 B.n603 B.n20 585
R265 B.n472 B.n19 585
R266 B.n604 B.n19 585
R267 B.n471 B.n470 585
R268 B.n470 B.n15 585
R269 B.n469 B.n14 585
R270 B.n610 B.n14 585
R271 B.n468 B.n13 585
R272 B.n611 B.n13 585
R273 B.n467 B.n12 585
R274 B.n612 B.n12 585
R275 B.n466 B.n465 585
R276 B.n465 B.n8 585
R277 B.n464 B.n7 585
R278 B.n618 B.n7 585
R279 B.n463 B.n6 585
R280 B.n619 B.n6 585
R281 B.n462 B.n5 585
R282 B.n620 B.n5 585
R283 B.n461 B.n460 585
R284 B.n460 B.n4 585
R285 B.n459 B.n156 585
R286 B.n459 B.n458 585
R287 B.n449 B.n157 585
R288 B.n158 B.n157 585
R289 B.n451 B.n450 585
R290 B.n452 B.n451 585
R291 B.n448 B.n162 585
R292 B.n166 B.n162 585
R293 B.n447 B.n446 585
R294 B.n446 B.n445 585
R295 B.n164 B.n163 585
R296 B.n165 B.n164 585
R297 B.n438 B.n437 585
R298 B.n439 B.n438 585
R299 B.n436 B.n171 585
R300 B.n171 B.n170 585
R301 B.n435 B.n434 585
R302 B.n434 B.n433 585
R303 B.n173 B.n172 585
R304 B.n174 B.n173 585
R305 B.n426 B.n425 585
R306 B.n427 B.n426 585
R307 B.n424 B.n179 585
R308 B.n179 B.n178 585
R309 B.n423 B.n422 585
R310 B.n422 B.n421 585
R311 B.n181 B.n180 585
R312 B.n182 B.n181 585
R313 B.n414 B.n413 585
R314 B.n415 B.n414 585
R315 B.n412 B.n187 585
R316 B.n187 B.n186 585
R317 B.n411 B.n410 585
R318 B.n410 B.n409 585
R319 B.n189 B.n188 585
R320 B.n190 B.n189 585
R321 B.n402 B.n401 585
R322 B.n403 B.n402 585
R323 B.n400 B.n195 585
R324 B.n195 B.n194 585
R325 B.n399 B.n398 585
R326 B.n398 B.n397 585
R327 B.n197 B.n196 585
R328 B.n198 B.n197 585
R329 B.n390 B.n389 585
R330 B.n391 B.n390 585
R331 B.n388 B.n202 585
R332 B.n206 B.n202 585
R333 B.n387 B.n386 585
R334 B.n386 B.n385 585
R335 B.n204 B.n203 585
R336 B.n205 B.n204 585
R337 B.n378 B.n377 585
R338 B.n379 B.n378 585
R339 B.n376 B.n211 585
R340 B.n211 B.n210 585
R341 B.n375 B.n374 585
R342 B.n374 B.n373 585
R343 B.n213 B.n212 585
R344 B.n366 B.n213 585
R345 B.n365 B.n364 585
R346 B.n367 B.n365 585
R347 B.n363 B.n218 585
R348 B.n218 B.n217 585
R349 B.n362 B.n361 585
R350 B.n361 B.n360 585
R351 B.n220 B.n219 585
R352 B.n221 B.n220 585
R353 B.n353 B.n352 585
R354 B.n354 B.n353 585
R355 B.n351 B.n226 585
R356 B.n226 B.n225 585
R357 B.n350 B.n349 585
R358 B.n349 B.n348 585
R359 B.n228 B.n227 585
R360 B.n229 B.n228 585
R361 B.n341 B.n340 585
R362 B.n342 B.n341 585
R363 B.n339 B.n233 585
R364 B.n237 B.n233 585
R365 B.n338 B.n337 585
R366 B.n337 B.n336 585
R367 B.n235 B.n234 585
R368 B.n236 B.n235 585
R369 B.n329 B.n328 585
R370 B.n330 B.n329 585
R371 B.n327 B.n242 585
R372 B.n242 B.n241 585
R373 B.n326 B.n325 585
R374 B.n325 B.n324 585
R375 B.n244 B.n243 585
R376 B.n245 B.n244 585
R377 B.n320 B.n319 585
R378 B.n248 B.n247 585
R379 B.n316 B.n315 585
R380 B.n317 B.n316 585
R381 B.n314 B.n261 585
R382 B.n313 B.n312 585
R383 B.n311 B.n310 585
R384 B.n309 B.n308 585
R385 B.n307 B.n306 585
R386 B.n305 B.n304 585
R387 B.n303 B.n302 585
R388 B.n301 B.n300 585
R389 B.n299 B.n298 585
R390 B.n297 B.n296 585
R391 B.n295 B.n294 585
R392 B.n293 B.n292 585
R393 B.n291 B.n290 585
R394 B.n289 B.n288 585
R395 B.n287 B.n286 585
R396 B.n284 B.n283 585
R397 B.n282 B.n281 585
R398 B.n280 B.n279 585
R399 B.n278 B.n277 585
R400 B.n276 B.n275 585
R401 B.n274 B.n273 585
R402 B.n272 B.n271 585
R403 B.n270 B.n269 585
R404 B.n268 B.n267 585
R405 B.n321 B.n246 585
R406 B.n246 B.n245 585
R407 B.n323 B.n322 585
R408 B.n324 B.n323 585
R409 B.n240 B.n239 585
R410 B.n241 B.n240 585
R411 B.n332 B.n331 585
R412 B.n331 B.n330 585
R413 B.n333 B.n238 585
R414 B.n238 B.n236 585
R415 B.n335 B.n334 585
R416 B.n336 B.n335 585
R417 B.n232 B.n231 585
R418 B.n237 B.n232 585
R419 B.n344 B.n343 585
R420 B.n343 B.n342 585
R421 B.n345 B.n230 585
R422 B.n230 B.n229 585
R423 B.n347 B.n346 585
R424 B.n348 B.n347 585
R425 B.n224 B.n223 585
R426 B.n225 B.n224 585
R427 B.n356 B.n355 585
R428 B.n355 B.n354 585
R429 B.n357 B.n222 585
R430 B.n222 B.n221 585
R431 B.n359 B.n358 585
R432 B.n360 B.n359 585
R433 B.n216 B.n215 585
R434 B.n217 B.n216 585
R435 B.n369 B.n368 585
R436 B.n368 B.n367 585
R437 B.n370 B.n214 585
R438 B.n366 B.n214 585
R439 B.n372 B.n371 585
R440 B.n373 B.n372 585
R441 B.n209 B.n208 585
R442 B.n210 B.n209 585
R443 B.n381 B.n380 585
R444 B.n380 B.n379 585
R445 B.n382 B.n207 585
R446 B.n207 B.n205 585
R447 B.n384 B.n383 585
R448 B.n385 B.n384 585
R449 B.n201 B.n200 585
R450 B.n206 B.n201 585
R451 B.n393 B.n392 585
R452 B.n392 B.n391 585
R453 B.n394 B.n199 585
R454 B.n199 B.n198 585
R455 B.n396 B.n395 585
R456 B.n397 B.n396 585
R457 B.n193 B.n192 585
R458 B.n194 B.n193 585
R459 B.n405 B.n404 585
R460 B.n404 B.n403 585
R461 B.n406 B.n191 585
R462 B.n191 B.n190 585
R463 B.n408 B.n407 585
R464 B.n409 B.n408 585
R465 B.n185 B.n184 585
R466 B.n186 B.n185 585
R467 B.n417 B.n416 585
R468 B.n416 B.n415 585
R469 B.n418 B.n183 585
R470 B.n183 B.n182 585
R471 B.n420 B.n419 585
R472 B.n421 B.n420 585
R473 B.n177 B.n176 585
R474 B.n178 B.n177 585
R475 B.n429 B.n428 585
R476 B.n428 B.n427 585
R477 B.n430 B.n175 585
R478 B.n175 B.n174 585
R479 B.n432 B.n431 585
R480 B.n433 B.n432 585
R481 B.n169 B.n168 585
R482 B.n170 B.n169 585
R483 B.n441 B.n440 585
R484 B.n440 B.n439 585
R485 B.n442 B.n167 585
R486 B.n167 B.n165 585
R487 B.n444 B.n443 585
R488 B.n445 B.n444 585
R489 B.n161 B.n160 585
R490 B.n166 B.n161 585
R491 B.n454 B.n453 585
R492 B.n453 B.n452 585
R493 B.n455 B.n159 585
R494 B.n159 B.n158 585
R495 B.n457 B.n456 585
R496 B.n458 B.n457 585
R497 B.n2 B.n0 585
R498 B.n4 B.n2 585
R499 B.n3 B.n1 585
R500 B.n619 B.n3 585
R501 B.n617 B.n616 585
R502 B.n618 B.n617 585
R503 B.n615 B.n9 585
R504 B.n9 B.n8 585
R505 B.n614 B.n613 585
R506 B.n613 B.n612 585
R507 B.n11 B.n10 585
R508 B.n611 B.n11 585
R509 B.n609 B.n608 585
R510 B.n610 B.n609 585
R511 B.n607 B.n16 585
R512 B.n16 B.n15 585
R513 B.n606 B.n605 585
R514 B.n605 B.n604 585
R515 B.n18 B.n17 585
R516 B.n603 B.n18 585
R517 B.n601 B.n600 585
R518 B.n602 B.n601 585
R519 B.n599 B.n23 585
R520 B.n23 B.n22 585
R521 B.n598 B.n597 585
R522 B.n597 B.n596 585
R523 B.n25 B.n24 585
R524 B.n595 B.n25 585
R525 B.n593 B.n592 585
R526 B.n594 B.n593 585
R527 B.n591 B.n30 585
R528 B.n30 B.n29 585
R529 B.n590 B.n589 585
R530 B.n589 B.n588 585
R531 B.n32 B.n31 585
R532 B.n587 B.n32 585
R533 B.n585 B.n584 585
R534 B.n586 B.n585 585
R535 B.n583 B.n37 585
R536 B.n37 B.n36 585
R537 B.n582 B.n581 585
R538 B.n581 B.n580 585
R539 B.n39 B.n38 585
R540 B.n579 B.n39 585
R541 B.n577 B.n576 585
R542 B.n578 B.n577 585
R543 B.n575 B.n44 585
R544 B.n44 B.n43 585
R545 B.n574 B.n573 585
R546 B.n573 B.n572 585
R547 B.n46 B.n45 585
R548 B.n571 B.n46 585
R549 B.n569 B.n568 585
R550 B.n570 B.n569 585
R551 B.n567 B.n51 585
R552 B.n51 B.n50 585
R553 B.n566 B.n565 585
R554 B.n565 B.n564 585
R555 B.n53 B.n52 585
R556 B.n563 B.n53 585
R557 B.n561 B.n560 585
R558 B.n562 B.n561 585
R559 B.n559 B.n57 585
R560 B.n60 B.n57 585
R561 B.n558 B.n557 585
R562 B.n557 B.n556 585
R563 B.n59 B.n58 585
R564 B.n555 B.n59 585
R565 B.n553 B.n552 585
R566 B.n554 B.n553 585
R567 B.n551 B.n65 585
R568 B.n65 B.n64 585
R569 B.n550 B.n549 585
R570 B.n549 B.n548 585
R571 B.n67 B.n66 585
R572 B.n547 B.n67 585
R573 B.n545 B.n544 585
R574 B.n546 B.n545 585
R575 B.n543 B.n72 585
R576 B.n72 B.n71 585
R577 B.n542 B.n541 585
R578 B.n541 B.n540 585
R579 B.n74 B.n73 585
R580 B.n539 B.n74 585
R581 B.n537 B.n536 585
R582 B.n538 B.n537 585
R583 B.n535 B.n79 585
R584 B.n79 B.n78 585
R585 B.n534 B.n533 585
R586 B.n533 B.n532 585
R587 B.n81 B.n80 585
R588 B.n531 B.n81 585
R589 B.n529 B.n528 585
R590 B.n530 B.n529 585
R591 B.n527 B.n86 585
R592 B.n86 B.n85 585
R593 B.n622 B.n621 585
R594 B.n621 B.n620 585
R595 B.n319 B.n246 468.476
R596 B.n525 B.n86 468.476
R597 B.n267 B.n244 468.476
R598 B.n522 B.n102 468.476
R599 B.n265 B.t23 278.012
R600 B.n262 B.t13 278.012
R601 B.n106 B.t16 278.012
R602 B.n103 B.t19 278.012
R603 B.n523 B.n100 256.663
R604 B.n523 B.n99 256.663
R605 B.n523 B.n98 256.663
R606 B.n523 B.n97 256.663
R607 B.n523 B.n96 256.663
R608 B.n523 B.n95 256.663
R609 B.n523 B.n94 256.663
R610 B.n523 B.n93 256.663
R611 B.n523 B.n92 256.663
R612 B.n523 B.n91 256.663
R613 B.n523 B.n90 256.663
R614 B.n523 B.n89 256.663
R615 B.n524 B.n523 256.663
R616 B.n318 B.n317 256.663
R617 B.n317 B.n249 256.663
R618 B.n317 B.n250 256.663
R619 B.n317 B.n251 256.663
R620 B.n317 B.n252 256.663
R621 B.n317 B.n253 256.663
R622 B.n317 B.n254 256.663
R623 B.n317 B.n255 256.663
R624 B.n317 B.n256 256.663
R625 B.n317 B.n257 256.663
R626 B.n317 B.n258 256.663
R627 B.n317 B.n259 256.663
R628 B.n317 B.n260 256.663
R629 B.n266 B.t22 235.345
R630 B.n263 B.t12 235.345
R631 B.n107 B.t17 235.345
R632 B.n104 B.t20 235.345
R633 B.n317 B.n245 216.543
R634 B.n523 B.n85 216.543
R635 B.n265 B.t21 208.024
R636 B.n262 B.t10 208.024
R637 B.n106 B.t14 208.024
R638 B.n103 B.t18 208.024
R639 B.n323 B.n246 163.367
R640 B.n323 B.n240 163.367
R641 B.n331 B.n240 163.367
R642 B.n331 B.n238 163.367
R643 B.n335 B.n238 163.367
R644 B.n335 B.n232 163.367
R645 B.n343 B.n232 163.367
R646 B.n343 B.n230 163.367
R647 B.n347 B.n230 163.367
R648 B.n347 B.n224 163.367
R649 B.n355 B.n224 163.367
R650 B.n355 B.n222 163.367
R651 B.n359 B.n222 163.367
R652 B.n359 B.n216 163.367
R653 B.n368 B.n216 163.367
R654 B.n368 B.n214 163.367
R655 B.n372 B.n214 163.367
R656 B.n372 B.n209 163.367
R657 B.n380 B.n209 163.367
R658 B.n380 B.n207 163.367
R659 B.n384 B.n207 163.367
R660 B.n384 B.n201 163.367
R661 B.n392 B.n201 163.367
R662 B.n392 B.n199 163.367
R663 B.n396 B.n199 163.367
R664 B.n396 B.n193 163.367
R665 B.n404 B.n193 163.367
R666 B.n404 B.n191 163.367
R667 B.n408 B.n191 163.367
R668 B.n408 B.n185 163.367
R669 B.n416 B.n185 163.367
R670 B.n416 B.n183 163.367
R671 B.n420 B.n183 163.367
R672 B.n420 B.n177 163.367
R673 B.n428 B.n177 163.367
R674 B.n428 B.n175 163.367
R675 B.n432 B.n175 163.367
R676 B.n432 B.n169 163.367
R677 B.n440 B.n169 163.367
R678 B.n440 B.n167 163.367
R679 B.n444 B.n167 163.367
R680 B.n444 B.n161 163.367
R681 B.n453 B.n161 163.367
R682 B.n453 B.n159 163.367
R683 B.n457 B.n159 163.367
R684 B.n457 B.n2 163.367
R685 B.n621 B.n2 163.367
R686 B.n621 B.n3 163.367
R687 B.n617 B.n3 163.367
R688 B.n617 B.n9 163.367
R689 B.n613 B.n9 163.367
R690 B.n613 B.n11 163.367
R691 B.n609 B.n11 163.367
R692 B.n609 B.n16 163.367
R693 B.n605 B.n16 163.367
R694 B.n605 B.n18 163.367
R695 B.n601 B.n18 163.367
R696 B.n601 B.n23 163.367
R697 B.n597 B.n23 163.367
R698 B.n597 B.n25 163.367
R699 B.n593 B.n25 163.367
R700 B.n593 B.n30 163.367
R701 B.n589 B.n30 163.367
R702 B.n589 B.n32 163.367
R703 B.n585 B.n32 163.367
R704 B.n585 B.n37 163.367
R705 B.n581 B.n37 163.367
R706 B.n581 B.n39 163.367
R707 B.n577 B.n39 163.367
R708 B.n577 B.n44 163.367
R709 B.n573 B.n44 163.367
R710 B.n573 B.n46 163.367
R711 B.n569 B.n46 163.367
R712 B.n569 B.n51 163.367
R713 B.n565 B.n51 163.367
R714 B.n565 B.n53 163.367
R715 B.n561 B.n53 163.367
R716 B.n561 B.n57 163.367
R717 B.n557 B.n57 163.367
R718 B.n557 B.n59 163.367
R719 B.n553 B.n59 163.367
R720 B.n553 B.n65 163.367
R721 B.n549 B.n65 163.367
R722 B.n549 B.n67 163.367
R723 B.n545 B.n67 163.367
R724 B.n545 B.n72 163.367
R725 B.n541 B.n72 163.367
R726 B.n541 B.n74 163.367
R727 B.n537 B.n74 163.367
R728 B.n537 B.n79 163.367
R729 B.n533 B.n79 163.367
R730 B.n533 B.n81 163.367
R731 B.n529 B.n81 163.367
R732 B.n529 B.n86 163.367
R733 B.n316 B.n248 163.367
R734 B.n316 B.n261 163.367
R735 B.n312 B.n311 163.367
R736 B.n308 B.n307 163.367
R737 B.n304 B.n303 163.367
R738 B.n300 B.n299 163.367
R739 B.n296 B.n295 163.367
R740 B.n292 B.n291 163.367
R741 B.n288 B.n287 163.367
R742 B.n283 B.n282 163.367
R743 B.n279 B.n278 163.367
R744 B.n275 B.n274 163.367
R745 B.n271 B.n270 163.367
R746 B.n325 B.n244 163.367
R747 B.n325 B.n242 163.367
R748 B.n329 B.n242 163.367
R749 B.n329 B.n235 163.367
R750 B.n337 B.n235 163.367
R751 B.n337 B.n233 163.367
R752 B.n341 B.n233 163.367
R753 B.n341 B.n228 163.367
R754 B.n349 B.n228 163.367
R755 B.n349 B.n226 163.367
R756 B.n353 B.n226 163.367
R757 B.n353 B.n220 163.367
R758 B.n361 B.n220 163.367
R759 B.n361 B.n218 163.367
R760 B.n365 B.n218 163.367
R761 B.n365 B.n213 163.367
R762 B.n374 B.n213 163.367
R763 B.n374 B.n211 163.367
R764 B.n378 B.n211 163.367
R765 B.n378 B.n204 163.367
R766 B.n386 B.n204 163.367
R767 B.n386 B.n202 163.367
R768 B.n390 B.n202 163.367
R769 B.n390 B.n197 163.367
R770 B.n398 B.n197 163.367
R771 B.n398 B.n195 163.367
R772 B.n402 B.n195 163.367
R773 B.n402 B.n189 163.367
R774 B.n410 B.n189 163.367
R775 B.n410 B.n187 163.367
R776 B.n414 B.n187 163.367
R777 B.n414 B.n181 163.367
R778 B.n422 B.n181 163.367
R779 B.n422 B.n179 163.367
R780 B.n426 B.n179 163.367
R781 B.n426 B.n173 163.367
R782 B.n434 B.n173 163.367
R783 B.n434 B.n171 163.367
R784 B.n438 B.n171 163.367
R785 B.n438 B.n164 163.367
R786 B.n446 B.n164 163.367
R787 B.n446 B.n162 163.367
R788 B.n451 B.n162 163.367
R789 B.n451 B.n157 163.367
R790 B.n459 B.n157 163.367
R791 B.n460 B.n459 163.367
R792 B.n460 B.n5 163.367
R793 B.n6 B.n5 163.367
R794 B.n7 B.n6 163.367
R795 B.n465 B.n7 163.367
R796 B.n465 B.n12 163.367
R797 B.n13 B.n12 163.367
R798 B.n14 B.n13 163.367
R799 B.n470 B.n14 163.367
R800 B.n470 B.n19 163.367
R801 B.n20 B.n19 163.367
R802 B.n21 B.n20 163.367
R803 B.n475 B.n21 163.367
R804 B.n475 B.n26 163.367
R805 B.n27 B.n26 163.367
R806 B.n28 B.n27 163.367
R807 B.n480 B.n28 163.367
R808 B.n480 B.n33 163.367
R809 B.n34 B.n33 163.367
R810 B.n35 B.n34 163.367
R811 B.n485 B.n35 163.367
R812 B.n485 B.n40 163.367
R813 B.n41 B.n40 163.367
R814 B.n42 B.n41 163.367
R815 B.n490 B.n42 163.367
R816 B.n490 B.n47 163.367
R817 B.n48 B.n47 163.367
R818 B.n49 B.n48 163.367
R819 B.n495 B.n49 163.367
R820 B.n495 B.n54 163.367
R821 B.n55 B.n54 163.367
R822 B.n56 B.n55 163.367
R823 B.n500 B.n56 163.367
R824 B.n500 B.n61 163.367
R825 B.n62 B.n61 163.367
R826 B.n63 B.n62 163.367
R827 B.n505 B.n63 163.367
R828 B.n505 B.n68 163.367
R829 B.n69 B.n68 163.367
R830 B.n70 B.n69 163.367
R831 B.n510 B.n70 163.367
R832 B.n510 B.n75 163.367
R833 B.n76 B.n75 163.367
R834 B.n77 B.n76 163.367
R835 B.n515 B.n77 163.367
R836 B.n515 B.n82 163.367
R837 B.n83 B.n82 163.367
R838 B.n84 B.n83 163.367
R839 B.n102 B.n84 163.367
R840 B.n108 B.n88 163.367
R841 B.n112 B.n111 163.367
R842 B.n116 B.n115 163.367
R843 B.n120 B.n119 163.367
R844 B.n125 B.n124 163.367
R845 B.n129 B.n128 163.367
R846 B.n133 B.n132 163.367
R847 B.n137 B.n136 163.367
R848 B.n141 B.n140 163.367
R849 B.n145 B.n144 163.367
R850 B.n149 B.n148 163.367
R851 B.n153 B.n152 163.367
R852 B.n522 B.n101 163.367
R853 B.n324 B.n245 123.74
R854 B.n324 B.n241 123.74
R855 B.n330 B.n241 123.74
R856 B.n330 B.n236 123.74
R857 B.n336 B.n236 123.74
R858 B.n336 B.n237 123.74
R859 B.n342 B.n229 123.74
R860 B.n348 B.n229 123.74
R861 B.n348 B.n225 123.74
R862 B.n354 B.n225 123.74
R863 B.n354 B.n221 123.74
R864 B.n360 B.n221 123.74
R865 B.n360 B.n217 123.74
R866 B.n367 B.n217 123.74
R867 B.n367 B.n366 123.74
R868 B.n373 B.n210 123.74
R869 B.n379 B.n210 123.74
R870 B.n379 B.n205 123.74
R871 B.n385 B.n205 123.74
R872 B.n385 B.n206 123.74
R873 B.n391 B.n198 123.74
R874 B.n397 B.n198 123.74
R875 B.n397 B.n194 123.74
R876 B.n403 B.n194 123.74
R877 B.n403 B.n190 123.74
R878 B.n409 B.n190 123.74
R879 B.n415 B.n186 123.74
R880 B.n415 B.n182 123.74
R881 B.n421 B.n182 123.74
R882 B.n421 B.n178 123.74
R883 B.n427 B.n178 123.74
R884 B.n433 B.n174 123.74
R885 B.n433 B.n170 123.74
R886 B.n439 B.n170 123.74
R887 B.n439 B.n165 123.74
R888 B.n445 B.n165 123.74
R889 B.n445 B.n166 123.74
R890 B.n452 B.n158 123.74
R891 B.n458 B.n158 123.74
R892 B.n458 B.n4 123.74
R893 B.n620 B.n4 123.74
R894 B.n620 B.n619 123.74
R895 B.n619 B.n618 123.74
R896 B.n618 B.n8 123.74
R897 B.n612 B.n8 123.74
R898 B.n611 B.n610 123.74
R899 B.n610 B.n15 123.74
R900 B.n604 B.n15 123.74
R901 B.n604 B.n603 123.74
R902 B.n603 B.n602 123.74
R903 B.n602 B.n22 123.74
R904 B.n596 B.n595 123.74
R905 B.n595 B.n594 123.74
R906 B.n594 B.n29 123.74
R907 B.n588 B.n29 123.74
R908 B.n588 B.n587 123.74
R909 B.n586 B.n36 123.74
R910 B.n580 B.n36 123.74
R911 B.n580 B.n579 123.74
R912 B.n579 B.n578 123.74
R913 B.n578 B.n43 123.74
R914 B.n572 B.n43 123.74
R915 B.n571 B.n570 123.74
R916 B.n570 B.n50 123.74
R917 B.n564 B.n50 123.74
R918 B.n564 B.n563 123.74
R919 B.n563 B.n562 123.74
R920 B.n556 B.n60 123.74
R921 B.n556 B.n555 123.74
R922 B.n555 B.n554 123.74
R923 B.n554 B.n64 123.74
R924 B.n548 B.n64 123.74
R925 B.n548 B.n547 123.74
R926 B.n547 B.n546 123.74
R927 B.n546 B.n71 123.74
R928 B.n540 B.n71 123.74
R929 B.n539 B.n538 123.74
R930 B.n538 B.n78 123.74
R931 B.n532 B.n78 123.74
R932 B.n532 B.n531 123.74
R933 B.n531 B.n530 123.74
R934 B.n530 B.n85 123.74
R935 B.n452 B.t7 103.722
R936 B.n612 B.t6 103.722
R937 B.t0 B.n186 96.4438
R938 B.n587 B.t1 96.4438
R939 B.n206 B.t4 92.8045
R940 B.t9 B.n571 92.8045
R941 B.n373 B.t8 89.1651
R942 B.n562 B.t5 89.1651
R943 B.n427 B.t3 85.5257
R944 B.n596 B.t2 85.5257
R945 B.n237 B.t11 74.6076
R946 B.t15 B.n539 74.6076
R947 B.n319 B.n318 71.676
R948 B.n261 B.n249 71.676
R949 B.n311 B.n250 71.676
R950 B.n307 B.n251 71.676
R951 B.n303 B.n252 71.676
R952 B.n299 B.n253 71.676
R953 B.n295 B.n254 71.676
R954 B.n291 B.n255 71.676
R955 B.n287 B.n256 71.676
R956 B.n282 B.n257 71.676
R957 B.n278 B.n258 71.676
R958 B.n274 B.n259 71.676
R959 B.n270 B.n260 71.676
R960 B.n525 B.n524 71.676
R961 B.n108 B.n89 71.676
R962 B.n112 B.n90 71.676
R963 B.n116 B.n91 71.676
R964 B.n120 B.n92 71.676
R965 B.n125 B.n93 71.676
R966 B.n129 B.n94 71.676
R967 B.n133 B.n95 71.676
R968 B.n137 B.n96 71.676
R969 B.n141 B.n97 71.676
R970 B.n145 B.n98 71.676
R971 B.n149 B.n99 71.676
R972 B.n153 B.n100 71.676
R973 B.n101 B.n100 71.676
R974 B.n152 B.n99 71.676
R975 B.n148 B.n98 71.676
R976 B.n144 B.n97 71.676
R977 B.n140 B.n96 71.676
R978 B.n136 B.n95 71.676
R979 B.n132 B.n94 71.676
R980 B.n128 B.n93 71.676
R981 B.n124 B.n92 71.676
R982 B.n119 B.n91 71.676
R983 B.n115 B.n90 71.676
R984 B.n111 B.n89 71.676
R985 B.n524 B.n88 71.676
R986 B.n318 B.n248 71.676
R987 B.n312 B.n249 71.676
R988 B.n308 B.n250 71.676
R989 B.n304 B.n251 71.676
R990 B.n300 B.n252 71.676
R991 B.n296 B.n253 71.676
R992 B.n292 B.n254 71.676
R993 B.n288 B.n255 71.676
R994 B.n283 B.n256 71.676
R995 B.n279 B.n257 71.676
R996 B.n275 B.n258 71.676
R997 B.n271 B.n259 71.676
R998 B.n267 B.n260 71.676
R999 B.n285 B.n266 59.5399
R1000 B.n264 B.n263 59.5399
R1001 B.n122 B.n107 59.5399
R1002 B.n105 B.n104 59.5399
R1003 B.n342 B.t11 49.132
R1004 B.n540 B.t15 49.132
R1005 B.n266 B.n265 42.6672
R1006 B.n263 B.n262 42.6672
R1007 B.n107 B.n106 42.6672
R1008 B.n104 B.n103 42.6672
R1009 B.t3 B.n174 38.2139
R1010 B.t2 B.n22 38.2139
R1011 B.n366 B.t8 34.5745
R1012 B.n60 B.t5 34.5745
R1013 B.n391 B.t4 30.9352
R1014 B.n572 B.t9 30.9352
R1015 B.n527 B.n526 30.4395
R1016 B.n521 B.n520 30.4395
R1017 B.n268 B.n243 30.4395
R1018 B.n321 B.n320 30.4395
R1019 B.n409 B.t0 27.2958
R1020 B.t1 B.n586 27.2958
R1021 B.n166 B.t7 20.017
R1022 B.t6 B.n611 20.017
R1023 B B.n622 18.0485
R1024 B.n526 B.n87 10.6151
R1025 B.n109 B.n87 10.6151
R1026 B.n110 B.n109 10.6151
R1027 B.n113 B.n110 10.6151
R1028 B.n114 B.n113 10.6151
R1029 B.n117 B.n114 10.6151
R1030 B.n118 B.n117 10.6151
R1031 B.n121 B.n118 10.6151
R1032 B.n126 B.n123 10.6151
R1033 B.n127 B.n126 10.6151
R1034 B.n130 B.n127 10.6151
R1035 B.n131 B.n130 10.6151
R1036 B.n134 B.n131 10.6151
R1037 B.n135 B.n134 10.6151
R1038 B.n138 B.n135 10.6151
R1039 B.n139 B.n138 10.6151
R1040 B.n143 B.n142 10.6151
R1041 B.n146 B.n143 10.6151
R1042 B.n147 B.n146 10.6151
R1043 B.n150 B.n147 10.6151
R1044 B.n151 B.n150 10.6151
R1045 B.n154 B.n151 10.6151
R1046 B.n155 B.n154 10.6151
R1047 B.n521 B.n155 10.6151
R1048 B.n326 B.n243 10.6151
R1049 B.n327 B.n326 10.6151
R1050 B.n328 B.n327 10.6151
R1051 B.n328 B.n234 10.6151
R1052 B.n338 B.n234 10.6151
R1053 B.n339 B.n338 10.6151
R1054 B.n340 B.n339 10.6151
R1055 B.n340 B.n227 10.6151
R1056 B.n350 B.n227 10.6151
R1057 B.n351 B.n350 10.6151
R1058 B.n352 B.n351 10.6151
R1059 B.n352 B.n219 10.6151
R1060 B.n362 B.n219 10.6151
R1061 B.n363 B.n362 10.6151
R1062 B.n364 B.n363 10.6151
R1063 B.n364 B.n212 10.6151
R1064 B.n375 B.n212 10.6151
R1065 B.n376 B.n375 10.6151
R1066 B.n377 B.n376 10.6151
R1067 B.n377 B.n203 10.6151
R1068 B.n387 B.n203 10.6151
R1069 B.n388 B.n387 10.6151
R1070 B.n389 B.n388 10.6151
R1071 B.n389 B.n196 10.6151
R1072 B.n399 B.n196 10.6151
R1073 B.n400 B.n399 10.6151
R1074 B.n401 B.n400 10.6151
R1075 B.n401 B.n188 10.6151
R1076 B.n411 B.n188 10.6151
R1077 B.n412 B.n411 10.6151
R1078 B.n413 B.n412 10.6151
R1079 B.n413 B.n180 10.6151
R1080 B.n423 B.n180 10.6151
R1081 B.n424 B.n423 10.6151
R1082 B.n425 B.n424 10.6151
R1083 B.n425 B.n172 10.6151
R1084 B.n435 B.n172 10.6151
R1085 B.n436 B.n435 10.6151
R1086 B.n437 B.n436 10.6151
R1087 B.n437 B.n163 10.6151
R1088 B.n447 B.n163 10.6151
R1089 B.n448 B.n447 10.6151
R1090 B.n450 B.n448 10.6151
R1091 B.n450 B.n449 10.6151
R1092 B.n449 B.n156 10.6151
R1093 B.n461 B.n156 10.6151
R1094 B.n462 B.n461 10.6151
R1095 B.n463 B.n462 10.6151
R1096 B.n464 B.n463 10.6151
R1097 B.n466 B.n464 10.6151
R1098 B.n467 B.n466 10.6151
R1099 B.n468 B.n467 10.6151
R1100 B.n469 B.n468 10.6151
R1101 B.n471 B.n469 10.6151
R1102 B.n472 B.n471 10.6151
R1103 B.n473 B.n472 10.6151
R1104 B.n474 B.n473 10.6151
R1105 B.n476 B.n474 10.6151
R1106 B.n477 B.n476 10.6151
R1107 B.n478 B.n477 10.6151
R1108 B.n479 B.n478 10.6151
R1109 B.n481 B.n479 10.6151
R1110 B.n482 B.n481 10.6151
R1111 B.n483 B.n482 10.6151
R1112 B.n484 B.n483 10.6151
R1113 B.n486 B.n484 10.6151
R1114 B.n487 B.n486 10.6151
R1115 B.n488 B.n487 10.6151
R1116 B.n489 B.n488 10.6151
R1117 B.n491 B.n489 10.6151
R1118 B.n492 B.n491 10.6151
R1119 B.n493 B.n492 10.6151
R1120 B.n494 B.n493 10.6151
R1121 B.n496 B.n494 10.6151
R1122 B.n497 B.n496 10.6151
R1123 B.n498 B.n497 10.6151
R1124 B.n499 B.n498 10.6151
R1125 B.n501 B.n499 10.6151
R1126 B.n502 B.n501 10.6151
R1127 B.n503 B.n502 10.6151
R1128 B.n504 B.n503 10.6151
R1129 B.n506 B.n504 10.6151
R1130 B.n507 B.n506 10.6151
R1131 B.n508 B.n507 10.6151
R1132 B.n509 B.n508 10.6151
R1133 B.n511 B.n509 10.6151
R1134 B.n512 B.n511 10.6151
R1135 B.n513 B.n512 10.6151
R1136 B.n514 B.n513 10.6151
R1137 B.n516 B.n514 10.6151
R1138 B.n517 B.n516 10.6151
R1139 B.n518 B.n517 10.6151
R1140 B.n519 B.n518 10.6151
R1141 B.n520 B.n519 10.6151
R1142 B.n320 B.n247 10.6151
R1143 B.n315 B.n247 10.6151
R1144 B.n315 B.n314 10.6151
R1145 B.n314 B.n313 10.6151
R1146 B.n313 B.n310 10.6151
R1147 B.n310 B.n309 10.6151
R1148 B.n309 B.n306 10.6151
R1149 B.n306 B.n305 10.6151
R1150 B.n302 B.n301 10.6151
R1151 B.n301 B.n298 10.6151
R1152 B.n298 B.n297 10.6151
R1153 B.n297 B.n294 10.6151
R1154 B.n294 B.n293 10.6151
R1155 B.n293 B.n290 10.6151
R1156 B.n290 B.n289 10.6151
R1157 B.n289 B.n286 10.6151
R1158 B.n284 B.n281 10.6151
R1159 B.n281 B.n280 10.6151
R1160 B.n280 B.n277 10.6151
R1161 B.n277 B.n276 10.6151
R1162 B.n276 B.n273 10.6151
R1163 B.n273 B.n272 10.6151
R1164 B.n272 B.n269 10.6151
R1165 B.n269 B.n268 10.6151
R1166 B.n322 B.n321 10.6151
R1167 B.n322 B.n239 10.6151
R1168 B.n332 B.n239 10.6151
R1169 B.n333 B.n332 10.6151
R1170 B.n334 B.n333 10.6151
R1171 B.n334 B.n231 10.6151
R1172 B.n344 B.n231 10.6151
R1173 B.n345 B.n344 10.6151
R1174 B.n346 B.n345 10.6151
R1175 B.n346 B.n223 10.6151
R1176 B.n356 B.n223 10.6151
R1177 B.n357 B.n356 10.6151
R1178 B.n358 B.n357 10.6151
R1179 B.n358 B.n215 10.6151
R1180 B.n369 B.n215 10.6151
R1181 B.n370 B.n369 10.6151
R1182 B.n371 B.n370 10.6151
R1183 B.n371 B.n208 10.6151
R1184 B.n381 B.n208 10.6151
R1185 B.n382 B.n381 10.6151
R1186 B.n383 B.n382 10.6151
R1187 B.n383 B.n200 10.6151
R1188 B.n393 B.n200 10.6151
R1189 B.n394 B.n393 10.6151
R1190 B.n395 B.n394 10.6151
R1191 B.n395 B.n192 10.6151
R1192 B.n405 B.n192 10.6151
R1193 B.n406 B.n405 10.6151
R1194 B.n407 B.n406 10.6151
R1195 B.n407 B.n184 10.6151
R1196 B.n417 B.n184 10.6151
R1197 B.n418 B.n417 10.6151
R1198 B.n419 B.n418 10.6151
R1199 B.n419 B.n176 10.6151
R1200 B.n429 B.n176 10.6151
R1201 B.n430 B.n429 10.6151
R1202 B.n431 B.n430 10.6151
R1203 B.n431 B.n168 10.6151
R1204 B.n441 B.n168 10.6151
R1205 B.n442 B.n441 10.6151
R1206 B.n443 B.n442 10.6151
R1207 B.n443 B.n160 10.6151
R1208 B.n454 B.n160 10.6151
R1209 B.n455 B.n454 10.6151
R1210 B.n456 B.n455 10.6151
R1211 B.n456 B.n0 10.6151
R1212 B.n616 B.n1 10.6151
R1213 B.n616 B.n615 10.6151
R1214 B.n615 B.n614 10.6151
R1215 B.n614 B.n10 10.6151
R1216 B.n608 B.n10 10.6151
R1217 B.n608 B.n607 10.6151
R1218 B.n607 B.n606 10.6151
R1219 B.n606 B.n17 10.6151
R1220 B.n600 B.n17 10.6151
R1221 B.n600 B.n599 10.6151
R1222 B.n599 B.n598 10.6151
R1223 B.n598 B.n24 10.6151
R1224 B.n592 B.n24 10.6151
R1225 B.n592 B.n591 10.6151
R1226 B.n591 B.n590 10.6151
R1227 B.n590 B.n31 10.6151
R1228 B.n584 B.n31 10.6151
R1229 B.n584 B.n583 10.6151
R1230 B.n583 B.n582 10.6151
R1231 B.n582 B.n38 10.6151
R1232 B.n576 B.n38 10.6151
R1233 B.n576 B.n575 10.6151
R1234 B.n575 B.n574 10.6151
R1235 B.n574 B.n45 10.6151
R1236 B.n568 B.n45 10.6151
R1237 B.n568 B.n567 10.6151
R1238 B.n567 B.n566 10.6151
R1239 B.n566 B.n52 10.6151
R1240 B.n560 B.n52 10.6151
R1241 B.n560 B.n559 10.6151
R1242 B.n559 B.n558 10.6151
R1243 B.n558 B.n58 10.6151
R1244 B.n552 B.n58 10.6151
R1245 B.n552 B.n551 10.6151
R1246 B.n551 B.n550 10.6151
R1247 B.n550 B.n66 10.6151
R1248 B.n544 B.n66 10.6151
R1249 B.n544 B.n543 10.6151
R1250 B.n543 B.n542 10.6151
R1251 B.n542 B.n73 10.6151
R1252 B.n536 B.n73 10.6151
R1253 B.n536 B.n535 10.6151
R1254 B.n535 B.n534 10.6151
R1255 B.n534 B.n80 10.6151
R1256 B.n528 B.n80 10.6151
R1257 B.n528 B.n527 10.6151
R1258 B.n123 B.n122 6.5566
R1259 B.n139 B.n105 6.5566
R1260 B.n302 B.n264 6.5566
R1261 B.n286 B.n285 6.5566
R1262 B.n122 B.n121 4.05904
R1263 B.n142 B.n105 4.05904
R1264 B.n305 B.n264 4.05904
R1265 B.n285 B.n284 4.05904
R1266 B.n622 B.n0 2.81026
R1267 B.n622 B.n1 2.81026
R1268 VP.n18 VP.n15 161.3
R1269 VP.n20 VP.n19 161.3
R1270 VP.n21 VP.n14 161.3
R1271 VP.n23 VP.n22 161.3
R1272 VP.n24 VP.n13 161.3
R1273 VP.n26 VP.n25 161.3
R1274 VP.n27 VP.n12 161.3
R1275 VP.n29 VP.n28 161.3
R1276 VP.n30 VP.n11 161.3
R1277 VP.n33 VP.n32 161.3
R1278 VP.n34 VP.n10 161.3
R1279 VP.n36 VP.n35 161.3
R1280 VP.n37 VP.n9 161.3
R1281 VP.n68 VP.n0 161.3
R1282 VP.n67 VP.n66 161.3
R1283 VP.n65 VP.n1 161.3
R1284 VP.n64 VP.n63 161.3
R1285 VP.n61 VP.n2 161.3
R1286 VP.n60 VP.n59 161.3
R1287 VP.n58 VP.n3 161.3
R1288 VP.n57 VP.n56 161.3
R1289 VP.n55 VP.n4 161.3
R1290 VP.n54 VP.n53 161.3
R1291 VP.n52 VP.n5 161.3
R1292 VP.n51 VP.n50 161.3
R1293 VP.n49 VP.n6 161.3
R1294 VP.n47 VP.n46 161.3
R1295 VP.n45 VP.n7 161.3
R1296 VP.n44 VP.n43 161.3
R1297 VP.n42 VP.n8 161.3
R1298 VP.n41 VP.n40 91.1828
R1299 VP.n70 VP.n69 91.1828
R1300 VP.n39 VP.n38 91.1828
R1301 VP.n17 VP.n16 59.9592
R1302 VP.n43 VP.n7 56.5193
R1303 VP.n67 VP.n1 56.5193
R1304 VP.n36 VP.n10 56.5193
R1305 VP.n50 VP.n5 50.2061
R1306 VP.n60 VP.n3 50.2061
R1307 VP.n29 VP.n12 50.2061
R1308 VP.n19 VP.n14 50.2061
R1309 VP.n40 VP.n39 40.6284
R1310 VP.n16 VP.t7 40.1933
R1311 VP.n54 VP.n5 30.7807
R1312 VP.n56 VP.n3 30.7807
R1313 VP.n25 VP.n12 30.7807
R1314 VP.n23 VP.n14 30.7807
R1315 VP.n43 VP.n42 24.4675
R1316 VP.n47 VP.n7 24.4675
R1317 VP.n50 VP.n49 24.4675
R1318 VP.n55 VP.n54 24.4675
R1319 VP.n56 VP.n55 24.4675
R1320 VP.n61 VP.n60 24.4675
R1321 VP.n63 VP.n1 24.4675
R1322 VP.n68 VP.n67 24.4675
R1323 VP.n37 VP.n36 24.4675
R1324 VP.n30 VP.n29 24.4675
R1325 VP.n32 VP.n10 24.4675
R1326 VP.n24 VP.n23 24.4675
R1327 VP.n25 VP.n24 24.4675
R1328 VP.n19 VP.n18 24.4675
R1329 VP.n42 VP.n41 19.5741
R1330 VP.n69 VP.n68 19.5741
R1331 VP.n38 VP.n37 19.5741
R1332 VP.n48 VP.n47 14.6807
R1333 VP.n63 VP.n62 14.6807
R1334 VP.n32 VP.n31 14.6807
R1335 VP.n16 VP.n15 13.3649
R1336 VP.n55 VP.t0 9.92403
R1337 VP.n41 VP.t3 9.92403
R1338 VP.n48 VP.t9 9.92403
R1339 VP.n62 VP.t4 9.92403
R1340 VP.n69 VP.t6 9.92403
R1341 VP.n24 VP.t1 9.92403
R1342 VP.n38 VP.t8 9.92403
R1343 VP.n31 VP.t2 9.92403
R1344 VP.n17 VP.t5 9.92403
R1345 VP.n49 VP.n48 9.7873
R1346 VP.n62 VP.n61 9.7873
R1347 VP.n31 VP.n30 9.7873
R1348 VP.n18 VP.n17 9.7873
R1349 VP.n39 VP.n9 0.278367
R1350 VP.n40 VP.n8 0.278367
R1351 VP.n70 VP.n0 0.278367
R1352 VP.n20 VP.n15 0.189894
R1353 VP.n21 VP.n20 0.189894
R1354 VP.n22 VP.n21 0.189894
R1355 VP.n22 VP.n13 0.189894
R1356 VP.n26 VP.n13 0.189894
R1357 VP.n27 VP.n26 0.189894
R1358 VP.n28 VP.n27 0.189894
R1359 VP.n28 VP.n11 0.189894
R1360 VP.n33 VP.n11 0.189894
R1361 VP.n34 VP.n33 0.189894
R1362 VP.n35 VP.n34 0.189894
R1363 VP.n35 VP.n9 0.189894
R1364 VP.n44 VP.n8 0.189894
R1365 VP.n45 VP.n44 0.189894
R1366 VP.n46 VP.n45 0.189894
R1367 VP.n46 VP.n6 0.189894
R1368 VP.n51 VP.n6 0.189894
R1369 VP.n52 VP.n51 0.189894
R1370 VP.n53 VP.n52 0.189894
R1371 VP.n53 VP.n4 0.189894
R1372 VP.n57 VP.n4 0.189894
R1373 VP.n58 VP.n57 0.189894
R1374 VP.n59 VP.n58 0.189894
R1375 VP.n59 VP.n2 0.189894
R1376 VP.n64 VP.n2 0.189894
R1377 VP.n65 VP.n64 0.189894
R1378 VP.n66 VP.n65 0.189894
R1379 VP.n66 VP.n0 0.189894
R1380 VP VP.n70 0.153454
R1381 VDD1.n1 VDD1.t2 264.772
R1382 VDD1.n3 VDD1.t6 264.772
R1383 VDD1.n5 VDD1.n4 238.529
R1384 VDD1.n7 VDD1.n6 237.161
R1385 VDD1.n1 VDD1.n0 237.161
R1386 VDD1.n3 VDD1.n2 237.161
R1387 VDD1.n7 VDD1.n5 34.919
R1388 VDD1.n6 VDD1.t7 25.7148
R1389 VDD1.n6 VDD1.t1 25.7148
R1390 VDD1.n0 VDD1.t4 25.7148
R1391 VDD1.n0 VDD1.t8 25.7148
R1392 VDD1.n4 VDD1.t5 25.7148
R1393 VDD1.n4 VDD1.t3 25.7148
R1394 VDD1.n2 VDD1.t0 25.7148
R1395 VDD1.n2 VDD1.t9 25.7148
R1396 VDD1 VDD1.n7 1.36472
R1397 VDD1 VDD1.n1 0.532828
R1398 VDD1.n5 VDD1.n3 0.419292
C0 VTAIL VN 2.29196f
C1 VTAIL VP 2.30609f
C2 VN VP 5.25629f
C3 VTAIL VDD2 4.4122f
C4 VDD2 VN 1.10111f
C5 VDD2 VP 0.499796f
C6 VTAIL VDD1 4.36363f
C7 VDD1 VN 0.160027f
C8 VDD1 VP 1.43688f
C9 VDD1 VDD2 1.69803f
C10 VDD2 B 4.183246f
C11 VDD1 B 4.295817f
C12 VTAIL B 2.831999f
C13 VN B 13.64084f
C14 VP B 12.147769f
C15 VDD1.t2 B 0.062376f
C16 VDD1.t4 B 0.012838f
C17 VDD1.t8 B 0.012838f
C18 VDD1.n0 B 0.031169f
C19 VDD1.n1 B 0.415205f
C20 VDD1.t6 B 0.062376f
C21 VDD1.t0 B 0.012838f
C22 VDD1.t9 B 0.012838f
C23 VDD1.n2 B 0.031169f
C24 VDD1.n3 B 0.408654f
C25 VDD1.t5 B 0.012838f
C26 VDD1.t3 B 0.012838f
C27 VDD1.n4 B 0.032804f
C28 VDD1.n5 B 1.5373f
C29 VDD1.t7 B 0.012838f
C30 VDD1.t1 B 0.012838f
C31 VDD1.n6 B 0.031169f
C32 VDD1.n7 B 1.55614f
C33 VP.n0 B 0.043967f
C34 VP.t6 B 0.076316f
C35 VP.n1 B 0.05333f
C36 VP.n2 B 0.033349f
C37 VP.t4 B 0.076316f
C38 VP.n3 B 0.031504f
C39 VP.n4 B 0.033349f
C40 VP.t0 B 0.076316f
C41 VP.n5 B 0.031504f
C42 VP.n6 B 0.033349f
C43 VP.t9 B 0.076316f
C44 VP.n7 B 0.05333f
C45 VP.n8 B 0.043967f
C46 VP.t3 B 0.076316f
C47 VP.n9 B 0.043967f
C48 VP.t8 B 0.076316f
C49 VP.n10 B 0.05333f
C50 VP.n11 B 0.033349f
C51 VP.t2 B 0.076316f
C52 VP.n12 B 0.031504f
C53 VP.n13 B 0.033349f
C54 VP.t1 B 0.076316f
C55 VP.n14 B 0.031504f
C56 VP.n15 B 0.245707f
C57 VP.t5 B 0.076316f
C58 VP.t7 B 0.249292f
C59 VP.n16 B 0.134281f
C60 VP.n17 B 0.14852f
C61 VP.n18 B 0.043743f
C62 VP.n19 B 0.061208f
C63 VP.n20 B 0.033349f
C64 VP.n21 B 0.033349f
C65 VP.n22 B 0.033349f
C66 VP.n23 B 0.06681f
C67 VP.n24 B 0.107012f
C68 VP.n25 B 0.06681f
C69 VP.n26 B 0.033349f
C70 VP.n27 B 0.033349f
C71 VP.n28 B 0.033349f
C72 VP.n29 B 0.061208f
C73 VP.n30 B 0.043743f
C74 VP.n31 B 0.075544f
C75 VP.n32 B 0.04988f
C76 VP.n33 B 0.033349f
C77 VP.n34 B 0.033349f
C78 VP.n35 B 0.033349f
C79 VP.n36 B 0.044037f
C80 VP.n37 B 0.056017f
C81 VP.n38 B 0.170776f
C82 VP.n39 B 1.32825f
C83 VP.n40 B 1.35776f
C84 VP.n41 B 0.170776f
C85 VP.n42 B 0.056017f
C86 VP.n43 B 0.044037f
C87 VP.n44 B 0.033349f
C88 VP.n45 B 0.033349f
C89 VP.n46 B 0.033349f
C90 VP.n47 B 0.04988f
C91 VP.n48 B 0.075544f
C92 VP.n49 B 0.043743f
C93 VP.n50 B 0.061208f
C94 VP.n51 B 0.033349f
C95 VP.n52 B 0.033349f
C96 VP.n53 B 0.033349f
C97 VP.n54 B 0.06681f
C98 VP.n55 B 0.107012f
C99 VP.n56 B 0.06681f
C100 VP.n57 B 0.033349f
C101 VP.n58 B 0.033349f
C102 VP.n59 B 0.033349f
C103 VP.n60 B 0.061208f
C104 VP.n61 B 0.043743f
C105 VP.n62 B 0.075544f
C106 VP.n63 B 0.04988f
C107 VP.n64 B 0.033349f
C108 VP.n65 B 0.033349f
C109 VP.n66 B 0.033349f
C110 VP.n67 B 0.044037f
C111 VP.n68 B 0.056017f
C112 VP.n69 B 0.170776f
C113 VP.n70 B 0.039968f
C114 VTAIL.t10 B 0.030843f
C115 VTAIL.t12 B 0.030843f
C116 VTAIL.n0 B 0.065724f
C117 VTAIL.n1 B 0.544456f
C118 VTAIL.t7 B 0.137413f
C119 VTAIL.n2 B 0.624823f
C120 VTAIL.t0 B 0.030843f
C121 VTAIL.t3 B 0.030843f
C122 VTAIL.n3 B 0.065724f
C123 VTAIL.n4 B 0.69054f
C124 VTAIL.t8 B 0.030843f
C125 VTAIL.t4 B 0.030843f
C126 VTAIL.n5 B 0.065724f
C127 VTAIL.n6 B 1.79729f
C128 VTAIL.t16 B 0.030843f
C129 VTAIL.t17 B 0.030843f
C130 VTAIL.n7 B 0.065724f
C131 VTAIL.n8 B 1.79729f
C132 VTAIL.t13 B 0.030843f
C133 VTAIL.t15 B 0.030843f
C134 VTAIL.n9 B 0.065724f
C135 VTAIL.n10 B 0.69054f
C136 VTAIL.t11 B 0.137413f
C137 VTAIL.n11 B 0.624823f
C138 VTAIL.t6 B 0.030843f
C139 VTAIL.t2 B 0.030843f
C140 VTAIL.n12 B 0.065724f
C141 VTAIL.n13 B 0.612394f
C142 VTAIL.t1 B 0.030843f
C143 VTAIL.t9 B 0.030843f
C144 VTAIL.n14 B 0.065724f
C145 VTAIL.n15 B 0.69054f
C146 VTAIL.t5 B 0.137413f
C147 VTAIL.n16 B 1.49995f
C148 VTAIL.t18 B 0.137413f
C149 VTAIL.n17 B 1.49995f
C150 VTAIL.t14 B 0.030843f
C151 VTAIL.t19 B 0.030843f
C152 VTAIL.n18 B 0.065724f
C153 VTAIL.n19 B 0.448709f
C154 VDD2.t0 B 0.063501f
C155 VDD2.t2 B 0.01307f
C156 VDD2.t9 B 0.01307f
C157 VDD2.n0 B 0.031731f
C158 VDD2.n1 B 0.416022f
C159 VDD2.t6 B 0.01307f
C160 VDD2.t5 B 0.01307f
C161 VDD2.n2 B 0.033395f
C162 VDD2.n3 B 1.4822f
C163 VDD2.t8 B 0.062063f
C164 VDD2.n4 B 1.49857f
C165 VDD2.t4 B 0.01307f
C166 VDD2.t1 B 0.01307f
C167 VDD2.n5 B 0.031731f
C168 VDD2.n6 B 0.223504f
C169 VDD2.t3 B 0.01307f
C170 VDD2.t7 B 0.01307f
C171 VDD2.n7 B 0.033388f
C172 VN.n0 B 0.043698f
C173 VN.t1 B 0.075848f
C174 VN.n1 B 0.053003f
C175 VN.n2 B 0.033145f
C176 VN.t0 B 0.075848f
C177 VN.n3 B 0.031311f
C178 VN.n4 B 0.033145f
C179 VN.t5 B 0.075848f
C180 VN.n5 B 0.031311f
C181 VN.n6 B 0.2442f
C182 VN.t7 B 0.075848f
C183 VN.t9 B 0.247764f
C184 VN.n7 B 0.133458f
C185 VN.n8 B 0.14761f
C186 VN.n9 B 0.043475f
C187 VN.n10 B 0.060833f
C188 VN.n11 B 0.033145f
C189 VN.n12 B 0.033145f
C190 VN.n13 B 0.033145f
C191 VN.n14 B 0.0664f
C192 VN.n15 B 0.106356f
C193 VN.n16 B 0.0664f
C194 VN.n17 B 0.033145f
C195 VN.n18 B 0.033145f
C196 VN.n19 B 0.033145f
C197 VN.n20 B 0.060833f
C198 VN.n21 B 0.043475f
C199 VN.n22 B 0.07508f
C200 VN.n23 B 0.049574f
C201 VN.n24 B 0.033145f
C202 VN.n25 B 0.033145f
C203 VN.n26 B 0.033145f
C204 VN.n27 B 0.043767f
C205 VN.n28 B 0.055674f
C206 VN.n29 B 0.169729f
C207 VN.n30 B 0.039723f
C208 VN.n31 B 0.043698f
C209 VN.t3 B 0.075848f
C210 VN.n32 B 0.053003f
C211 VN.n33 B 0.033145f
C212 VN.t2 B 0.075848f
C213 VN.n34 B 0.031311f
C214 VN.n35 B 0.033145f
C215 VN.t6 B 0.075848f
C216 VN.n36 B 0.031311f
C217 VN.n37 B 0.2442f
C218 VN.t4 B 0.075848f
C219 VN.t8 B 0.247764f
C220 VN.n38 B 0.133458f
C221 VN.n39 B 0.14761f
C222 VN.n40 B 0.043475f
C223 VN.n41 B 0.060833f
C224 VN.n42 B 0.033145f
C225 VN.n43 B 0.033145f
C226 VN.n44 B 0.033145f
C227 VN.n45 B 0.0664f
C228 VN.n46 B 0.106356f
C229 VN.n47 B 0.0664f
C230 VN.n48 B 0.033145f
C231 VN.n49 B 0.033145f
C232 VN.n50 B 0.033145f
C233 VN.n51 B 0.060833f
C234 VN.n52 B 0.043475f
C235 VN.n53 B 0.07508f
C236 VN.n54 B 0.049574f
C237 VN.n55 B 0.033145f
C238 VN.n56 B 0.033145f
C239 VN.n57 B 0.033145f
C240 VN.n58 B 0.043767f
C241 VN.n59 B 0.055674f
C242 VN.n60 B 0.169729f
C243 VN.n61 B 1.33857f
.ends

