* NGSPICE file created from diff_pair_sample_0440.ext - technology: sky130A

.subckt diff_pair_sample_0440 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=4.9881 pd=26.36 as=0 ps=0 w=12.79 l=2.41
X1 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=4.9881 pd=26.36 as=0 ps=0 w=12.79 l=2.41
X2 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.9881 pd=26.36 as=0 ps=0 w=12.79 l=2.41
X3 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=4.9881 pd=26.36 as=4.9881 ps=26.36 w=12.79 l=2.41
X4 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.9881 pd=26.36 as=0 ps=0 w=12.79 l=2.41
X5 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=4.9881 pd=26.36 as=4.9881 ps=26.36 w=12.79 l=2.41
X6 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.9881 pd=26.36 as=4.9881 ps=26.36 w=12.79 l=2.41
X7 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.9881 pd=26.36 as=4.9881 ps=26.36 w=12.79 l=2.41
R0 B.n690 B.n689 585
R1 B.n691 B.n690 585
R2 B.n291 B.n96 585
R3 B.n290 B.n289 585
R4 B.n288 B.n287 585
R5 B.n286 B.n285 585
R6 B.n284 B.n283 585
R7 B.n282 B.n281 585
R8 B.n280 B.n279 585
R9 B.n278 B.n277 585
R10 B.n276 B.n275 585
R11 B.n274 B.n273 585
R12 B.n272 B.n271 585
R13 B.n270 B.n269 585
R14 B.n268 B.n267 585
R15 B.n266 B.n265 585
R16 B.n264 B.n263 585
R17 B.n262 B.n261 585
R18 B.n260 B.n259 585
R19 B.n258 B.n257 585
R20 B.n256 B.n255 585
R21 B.n254 B.n253 585
R22 B.n252 B.n251 585
R23 B.n250 B.n249 585
R24 B.n248 B.n247 585
R25 B.n246 B.n245 585
R26 B.n244 B.n243 585
R27 B.n242 B.n241 585
R28 B.n240 B.n239 585
R29 B.n238 B.n237 585
R30 B.n236 B.n235 585
R31 B.n234 B.n233 585
R32 B.n232 B.n231 585
R33 B.n230 B.n229 585
R34 B.n228 B.n227 585
R35 B.n226 B.n225 585
R36 B.n224 B.n223 585
R37 B.n222 B.n221 585
R38 B.n220 B.n219 585
R39 B.n218 B.n217 585
R40 B.n216 B.n215 585
R41 B.n214 B.n213 585
R42 B.n212 B.n211 585
R43 B.n210 B.n209 585
R44 B.n208 B.n207 585
R45 B.n205 B.n204 585
R46 B.n203 B.n202 585
R47 B.n201 B.n200 585
R48 B.n199 B.n198 585
R49 B.n197 B.n196 585
R50 B.n195 B.n194 585
R51 B.n193 B.n192 585
R52 B.n191 B.n190 585
R53 B.n189 B.n188 585
R54 B.n187 B.n186 585
R55 B.n185 B.n184 585
R56 B.n183 B.n182 585
R57 B.n181 B.n180 585
R58 B.n179 B.n178 585
R59 B.n177 B.n176 585
R60 B.n175 B.n174 585
R61 B.n173 B.n172 585
R62 B.n171 B.n170 585
R63 B.n169 B.n168 585
R64 B.n167 B.n166 585
R65 B.n165 B.n164 585
R66 B.n163 B.n162 585
R67 B.n161 B.n160 585
R68 B.n159 B.n158 585
R69 B.n157 B.n156 585
R70 B.n155 B.n154 585
R71 B.n153 B.n152 585
R72 B.n151 B.n150 585
R73 B.n149 B.n148 585
R74 B.n147 B.n146 585
R75 B.n145 B.n144 585
R76 B.n143 B.n142 585
R77 B.n141 B.n140 585
R78 B.n139 B.n138 585
R79 B.n137 B.n136 585
R80 B.n135 B.n134 585
R81 B.n133 B.n132 585
R82 B.n131 B.n130 585
R83 B.n129 B.n128 585
R84 B.n127 B.n126 585
R85 B.n125 B.n124 585
R86 B.n123 B.n122 585
R87 B.n121 B.n120 585
R88 B.n119 B.n118 585
R89 B.n117 B.n116 585
R90 B.n115 B.n114 585
R91 B.n113 B.n112 585
R92 B.n111 B.n110 585
R93 B.n109 B.n108 585
R94 B.n107 B.n106 585
R95 B.n105 B.n104 585
R96 B.n103 B.n102 585
R97 B.n46 B.n45 585
R98 B.n688 B.n47 585
R99 B.n692 B.n47 585
R100 B.n687 B.n686 585
R101 B.n686 B.n43 585
R102 B.n685 B.n42 585
R103 B.n698 B.n42 585
R104 B.n684 B.n41 585
R105 B.n699 B.n41 585
R106 B.n683 B.n40 585
R107 B.n700 B.n40 585
R108 B.n682 B.n681 585
R109 B.n681 B.n36 585
R110 B.n680 B.n35 585
R111 B.n706 B.n35 585
R112 B.n679 B.n34 585
R113 B.n707 B.n34 585
R114 B.n678 B.n33 585
R115 B.n708 B.n33 585
R116 B.n677 B.n676 585
R117 B.n676 B.n29 585
R118 B.n675 B.n28 585
R119 B.n714 B.n28 585
R120 B.n674 B.n27 585
R121 B.n715 B.n27 585
R122 B.n673 B.n26 585
R123 B.n716 B.n26 585
R124 B.n672 B.n671 585
R125 B.n671 B.n22 585
R126 B.n670 B.n21 585
R127 B.n722 B.n21 585
R128 B.n669 B.n20 585
R129 B.n723 B.n20 585
R130 B.n668 B.n19 585
R131 B.n724 B.n19 585
R132 B.n667 B.n666 585
R133 B.n666 B.n15 585
R134 B.n665 B.n14 585
R135 B.n730 B.n14 585
R136 B.n664 B.n13 585
R137 B.n731 B.n13 585
R138 B.n663 B.n12 585
R139 B.n732 B.n12 585
R140 B.n662 B.n661 585
R141 B.n661 B.n8 585
R142 B.n660 B.n7 585
R143 B.n738 B.n7 585
R144 B.n659 B.n6 585
R145 B.n739 B.n6 585
R146 B.n658 B.n5 585
R147 B.n740 B.n5 585
R148 B.n657 B.n656 585
R149 B.n656 B.n4 585
R150 B.n655 B.n292 585
R151 B.n655 B.n654 585
R152 B.n645 B.n293 585
R153 B.n294 B.n293 585
R154 B.n647 B.n646 585
R155 B.n648 B.n647 585
R156 B.n644 B.n299 585
R157 B.n299 B.n298 585
R158 B.n643 B.n642 585
R159 B.n642 B.n641 585
R160 B.n301 B.n300 585
R161 B.n302 B.n301 585
R162 B.n634 B.n633 585
R163 B.n635 B.n634 585
R164 B.n632 B.n307 585
R165 B.n307 B.n306 585
R166 B.n631 B.n630 585
R167 B.n630 B.n629 585
R168 B.n309 B.n308 585
R169 B.n310 B.n309 585
R170 B.n622 B.n621 585
R171 B.n623 B.n622 585
R172 B.n620 B.n315 585
R173 B.n315 B.n314 585
R174 B.n619 B.n618 585
R175 B.n618 B.n617 585
R176 B.n317 B.n316 585
R177 B.n318 B.n317 585
R178 B.n610 B.n609 585
R179 B.n611 B.n610 585
R180 B.n608 B.n322 585
R181 B.n326 B.n322 585
R182 B.n607 B.n606 585
R183 B.n606 B.n605 585
R184 B.n324 B.n323 585
R185 B.n325 B.n324 585
R186 B.n598 B.n597 585
R187 B.n599 B.n598 585
R188 B.n596 B.n331 585
R189 B.n331 B.n330 585
R190 B.n595 B.n594 585
R191 B.n594 B.n593 585
R192 B.n333 B.n332 585
R193 B.n334 B.n333 585
R194 B.n586 B.n585 585
R195 B.n587 B.n586 585
R196 B.n337 B.n336 585
R197 B.n393 B.n391 585
R198 B.n394 B.n390 585
R199 B.n394 B.n338 585
R200 B.n397 B.n396 585
R201 B.n398 B.n389 585
R202 B.n400 B.n399 585
R203 B.n402 B.n388 585
R204 B.n405 B.n404 585
R205 B.n406 B.n387 585
R206 B.n408 B.n407 585
R207 B.n410 B.n386 585
R208 B.n413 B.n412 585
R209 B.n414 B.n385 585
R210 B.n416 B.n415 585
R211 B.n418 B.n384 585
R212 B.n421 B.n420 585
R213 B.n422 B.n383 585
R214 B.n424 B.n423 585
R215 B.n426 B.n382 585
R216 B.n429 B.n428 585
R217 B.n430 B.n381 585
R218 B.n432 B.n431 585
R219 B.n434 B.n380 585
R220 B.n437 B.n436 585
R221 B.n438 B.n379 585
R222 B.n440 B.n439 585
R223 B.n442 B.n378 585
R224 B.n445 B.n444 585
R225 B.n446 B.n377 585
R226 B.n448 B.n447 585
R227 B.n450 B.n376 585
R228 B.n453 B.n452 585
R229 B.n454 B.n375 585
R230 B.n456 B.n455 585
R231 B.n458 B.n374 585
R232 B.n461 B.n460 585
R233 B.n462 B.n373 585
R234 B.n464 B.n463 585
R235 B.n466 B.n372 585
R236 B.n469 B.n468 585
R237 B.n470 B.n371 585
R238 B.n472 B.n471 585
R239 B.n474 B.n370 585
R240 B.n477 B.n476 585
R241 B.n479 B.n367 585
R242 B.n481 B.n480 585
R243 B.n483 B.n366 585
R244 B.n486 B.n485 585
R245 B.n487 B.n365 585
R246 B.n489 B.n488 585
R247 B.n491 B.n364 585
R248 B.n494 B.n493 585
R249 B.n495 B.n361 585
R250 B.n498 B.n497 585
R251 B.n500 B.n360 585
R252 B.n503 B.n502 585
R253 B.n504 B.n359 585
R254 B.n506 B.n505 585
R255 B.n508 B.n358 585
R256 B.n511 B.n510 585
R257 B.n512 B.n357 585
R258 B.n514 B.n513 585
R259 B.n516 B.n356 585
R260 B.n519 B.n518 585
R261 B.n520 B.n355 585
R262 B.n522 B.n521 585
R263 B.n524 B.n354 585
R264 B.n527 B.n526 585
R265 B.n528 B.n353 585
R266 B.n530 B.n529 585
R267 B.n532 B.n352 585
R268 B.n535 B.n534 585
R269 B.n536 B.n351 585
R270 B.n538 B.n537 585
R271 B.n540 B.n350 585
R272 B.n543 B.n542 585
R273 B.n544 B.n349 585
R274 B.n546 B.n545 585
R275 B.n548 B.n348 585
R276 B.n551 B.n550 585
R277 B.n552 B.n347 585
R278 B.n554 B.n553 585
R279 B.n556 B.n346 585
R280 B.n559 B.n558 585
R281 B.n560 B.n345 585
R282 B.n562 B.n561 585
R283 B.n564 B.n344 585
R284 B.n567 B.n566 585
R285 B.n568 B.n343 585
R286 B.n570 B.n569 585
R287 B.n572 B.n342 585
R288 B.n575 B.n574 585
R289 B.n576 B.n341 585
R290 B.n578 B.n577 585
R291 B.n580 B.n340 585
R292 B.n583 B.n582 585
R293 B.n584 B.n339 585
R294 B.n589 B.n588 585
R295 B.n588 B.n587 585
R296 B.n590 B.n335 585
R297 B.n335 B.n334 585
R298 B.n592 B.n591 585
R299 B.n593 B.n592 585
R300 B.n329 B.n328 585
R301 B.n330 B.n329 585
R302 B.n601 B.n600 585
R303 B.n600 B.n599 585
R304 B.n602 B.n327 585
R305 B.n327 B.n325 585
R306 B.n604 B.n603 585
R307 B.n605 B.n604 585
R308 B.n321 B.n320 585
R309 B.n326 B.n321 585
R310 B.n613 B.n612 585
R311 B.n612 B.n611 585
R312 B.n614 B.n319 585
R313 B.n319 B.n318 585
R314 B.n616 B.n615 585
R315 B.n617 B.n616 585
R316 B.n313 B.n312 585
R317 B.n314 B.n313 585
R318 B.n625 B.n624 585
R319 B.n624 B.n623 585
R320 B.n626 B.n311 585
R321 B.n311 B.n310 585
R322 B.n628 B.n627 585
R323 B.n629 B.n628 585
R324 B.n305 B.n304 585
R325 B.n306 B.n305 585
R326 B.n637 B.n636 585
R327 B.n636 B.n635 585
R328 B.n638 B.n303 585
R329 B.n303 B.n302 585
R330 B.n640 B.n639 585
R331 B.n641 B.n640 585
R332 B.n297 B.n296 585
R333 B.n298 B.n297 585
R334 B.n650 B.n649 585
R335 B.n649 B.n648 585
R336 B.n651 B.n295 585
R337 B.n295 B.n294 585
R338 B.n653 B.n652 585
R339 B.n654 B.n653 585
R340 B.n2 B.n0 585
R341 B.n4 B.n2 585
R342 B.n3 B.n1 585
R343 B.n739 B.n3 585
R344 B.n737 B.n736 585
R345 B.n738 B.n737 585
R346 B.n735 B.n9 585
R347 B.n9 B.n8 585
R348 B.n734 B.n733 585
R349 B.n733 B.n732 585
R350 B.n11 B.n10 585
R351 B.n731 B.n11 585
R352 B.n729 B.n728 585
R353 B.n730 B.n729 585
R354 B.n727 B.n16 585
R355 B.n16 B.n15 585
R356 B.n726 B.n725 585
R357 B.n725 B.n724 585
R358 B.n18 B.n17 585
R359 B.n723 B.n18 585
R360 B.n721 B.n720 585
R361 B.n722 B.n721 585
R362 B.n719 B.n23 585
R363 B.n23 B.n22 585
R364 B.n718 B.n717 585
R365 B.n717 B.n716 585
R366 B.n25 B.n24 585
R367 B.n715 B.n25 585
R368 B.n713 B.n712 585
R369 B.n714 B.n713 585
R370 B.n711 B.n30 585
R371 B.n30 B.n29 585
R372 B.n710 B.n709 585
R373 B.n709 B.n708 585
R374 B.n32 B.n31 585
R375 B.n707 B.n32 585
R376 B.n705 B.n704 585
R377 B.n706 B.n705 585
R378 B.n703 B.n37 585
R379 B.n37 B.n36 585
R380 B.n702 B.n701 585
R381 B.n701 B.n700 585
R382 B.n39 B.n38 585
R383 B.n699 B.n39 585
R384 B.n697 B.n696 585
R385 B.n698 B.n697 585
R386 B.n695 B.n44 585
R387 B.n44 B.n43 585
R388 B.n694 B.n693 585
R389 B.n693 B.n692 585
R390 B.n742 B.n741 585
R391 B.n741 B.n740 585
R392 B.n588 B.n337 574.183
R393 B.n693 B.n46 574.183
R394 B.n586 B.n339 574.183
R395 B.n690 B.n47 574.183
R396 B.n362 B.t15 348.993
R397 B.n97 B.t4 348.993
R398 B.n368 B.t9 348.993
R399 B.n99 B.t11 348.993
R400 B.n362 B.t13 335.642
R401 B.n368 B.t6 335.642
R402 B.n99 B.t10 335.642
R403 B.n97 B.t2 335.642
R404 B.n363 B.t14 295.853
R405 B.n98 B.t5 295.853
R406 B.n369 B.t8 295.853
R407 B.n100 B.t12 295.853
R408 B.n691 B.n95 256.663
R409 B.n691 B.n94 256.663
R410 B.n691 B.n93 256.663
R411 B.n691 B.n92 256.663
R412 B.n691 B.n91 256.663
R413 B.n691 B.n90 256.663
R414 B.n691 B.n89 256.663
R415 B.n691 B.n88 256.663
R416 B.n691 B.n87 256.663
R417 B.n691 B.n86 256.663
R418 B.n691 B.n85 256.663
R419 B.n691 B.n84 256.663
R420 B.n691 B.n83 256.663
R421 B.n691 B.n82 256.663
R422 B.n691 B.n81 256.663
R423 B.n691 B.n80 256.663
R424 B.n691 B.n79 256.663
R425 B.n691 B.n78 256.663
R426 B.n691 B.n77 256.663
R427 B.n691 B.n76 256.663
R428 B.n691 B.n75 256.663
R429 B.n691 B.n74 256.663
R430 B.n691 B.n73 256.663
R431 B.n691 B.n72 256.663
R432 B.n691 B.n71 256.663
R433 B.n691 B.n70 256.663
R434 B.n691 B.n69 256.663
R435 B.n691 B.n68 256.663
R436 B.n691 B.n67 256.663
R437 B.n691 B.n66 256.663
R438 B.n691 B.n65 256.663
R439 B.n691 B.n64 256.663
R440 B.n691 B.n63 256.663
R441 B.n691 B.n62 256.663
R442 B.n691 B.n61 256.663
R443 B.n691 B.n60 256.663
R444 B.n691 B.n59 256.663
R445 B.n691 B.n58 256.663
R446 B.n691 B.n57 256.663
R447 B.n691 B.n56 256.663
R448 B.n691 B.n55 256.663
R449 B.n691 B.n54 256.663
R450 B.n691 B.n53 256.663
R451 B.n691 B.n52 256.663
R452 B.n691 B.n51 256.663
R453 B.n691 B.n50 256.663
R454 B.n691 B.n49 256.663
R455 B.n691 B.n48 256.663
R456 B.n392 B.n338 256.663
R457 B.n395 B.n338 256.663
R458 B.n401 B.n338 256.663
R459 B.n403 B.n338 256.663
R460 B.n409 B.n338 256.663
R461 B.n411 B.n338 256.663
R462 B.n417 B.n338 256.663
R463 B.n419 B.n338 256.663
R464 B.n425 B.n338 256.663
R465 B.n427 B.n338 256.663
R466 B.n433 B.n338 256.663
R467 B.n435 B.n338 256.663
R468 B.n441 B.n338 256.663
R469 B.n443 B.n338 256.663
R470 B.n449 B.n338 256.663
R471 B.n451 B.n338 256.663
R472 B.n457 B.n338 256.663
R473 B.n459 B.n338 256.663
R474 B.n465 B.n338 256.663
R475 B.n467 B.n338 256.663
R476 B.n473 B.n338 256.663
R477 B.n475 B.n338 256.663
R478 B.n482 B.n338 256.663
R479 B.n484 B.n338 256.663
R480 B.n490 B.n338 256.663
R481 B.n492 B.n338 256.663
R482 B.n499 B.n338 256.663
R483 B.n501 B.n338 256.663
R484 B.n507 B.n338 256.663
R485 B.n509 B.n338 256.663
R486 B.n515 B.n338 256.663
R487 B.n517 B.n338 256.663
R488 B.n523 B.n338 256.663
R489 B.n525 B.n338 256.663
R490 B.n531 B.n338 256.663
R491 B.n533 B.n338 256.663
R492 B.n539 B.n338 256.663
R493 B.n541 B.n338 256.663
R494 B.n547 B.n338 256.663
R495 B.n549 B.n338 256.663
R496 B.n555 B.n338 256.663
R497 B.n557 B.n338 256.663
R498 B.n563 B.n338 256.663
R499 B.n565 B.n338 256.663
R500 B.n571 B.n338 256.663
R501 B.n573 B.n338 256.663
R502 B.n579 B.n338 256.663
R503 B.n581 B.n338 256.663
R504 B.n588 B.n335 163.367
R505 B.n592 B.n335 163.367
R506 B.n592 B.n329 163.367
R507 B.n600 B.n329 163.367
R508 B.n600 B.n327 163.367
R509 B.n604 B.n327 163.367
R510 B.n604 B.n321 163.367
R511 B.n612 B.n321 163.367
R512 B.n612 B.n319 163.367
R513 B.n616 B.n319 163.367
R514 B.n616 B.n313 163.367
R515 B.n624 B.n313 163.367
R516 B.n624 B.n311 163.367
R517 B.n628 B.n311 163.367
R518 B.n628 B.n305 163.367
R519 B.n636 B.n305 163.367
R520 B.n636 B.n303 163.367
R521 B.n640 B.n303 163.367
R522 B.n640 B.n297 163.367
R523 B.n649 B.n297 163.367
R524 B.n649 B.n295 163.367
R525 B.n653 B.n295 163.367
R526 B.n653 B.n2 163.367
R527 B.n741 B.n2 163.367
R528 B.n741 B.n3 163.367
R529 B.n737 B.n3 163.367
R530 B.n737 B.n9 163.367
R531 B.n733 B.n9 163.367
R532 B.n733 B.n11 163.367
R533 B.n729 B.n11 163.367
R534 B.n729 B.n16 163.367
R535 B.n725 B.n16 163.367
R536 B.n725 B.n18 163.367
R537 B.n721 B.n18 163.367
R538 B.n721 B.n23 163.367
R539 B.n717 B.n23 163.367
R540 B.n717 B.n25 163.367
R541 B.n713 B.n25 163.367
R542 B.n713 B.n30 163.367
R543 B.n709 B.n30 163.367
R544 B.n709 B.n32 163.367
R545 B.n705 B.n32 163.367
R546 B.n705 B.n37 163.367
R547 B.n701 B.n37 163.367
R548 B.n701 B.n39 163.367
R549 B.n697 B.n39 163.367
R550 B.n697 B.n44 163.367
R551 B.n693 B.n44 163.367
R552 B.n394 B.n393 163.367
R553 B.n396 B.n394 163.367
R554 B.n400 B.n389 163.367
R555 B.n404 B.n402 163.367
R556 B.n408 B.n387 163.367
R557 B.n412 B.n410 163.367
R558 B.n416 B.n385 163.367
R559 B.n420 B.n418 163.367
R560 B.n424 B.n383 163.367
R561 B.n428 B.n426 163.367
R562 B.n432 B.n381 163.367
R563 B.n436 B.n434 163.367
R564 B.n440 B.n379 163.367
R565 B.n444 B.n442 163.367
R566 B.n448 B.n377 163.367
R567 B.n452 B.n450 163.367
R568 B.n456 B.n375 163.367
R569 B.n460 B.n458 163.367
R570 B.n464 B.n373 163.367
R571 B.n468 B.n466 163.367
R572 B.n472 B.n371 163.367
R573 B.n476 B.n474 163.367
R574 B.n481 B.n367 163.367
R575 B.n485 B.n483 163.367
R576 B.n489 B.n365 163.367
R577 B.n493 B.n491 163.367
R578 B.n498 B.n361 163.367
R579 B.n502 B.n500 163.367
R580 B.n506 B.n359 163.367
R581 B.n510 B.n508 163.367
R582 B.n514 B.n357 163.367
R583 B.n518 B.n516 163.367
R584 B.n522 B.n355 163.367
R585 B.n526 B.n524 163.367
R586 B.n530 B.n353 163.367
R587 B.n534 B.n532 163.367
R588 B.n538 B.n351 163.367
R589 B.n542 B.n540 163.367
R590 B.n546 B.n349 163.367
R591 B.n550 B.n548 163.367
R592 B.n554 B.n347 163.367
R593 B.n558 B.n556 163.367
R594 B.n562 B.n345 163.367
R595 B.n566 B.n564 163.367
R596 B.n570 B.n343 163.367
R597 B.n574 B.n572 163.367
R598 B.n578 B.n341 163.367
R599 B.n582 B.n580 163.367
R600 B.n586 B.n333 163.367
R601 B.n594 B.n333 163.367
R602 B.n594 B.n331 163.367
R603 B.n598 B.n331 163.367
R604 B.n598 B.n324 163.367
R605 B.n606 B.n324 163.367
R606 B.n606 B.n322 163.367
R607 B.n610 B.n322 163.367
R608 B.n610 B.n317 163.367
R609 B.n618 B.n317 163.367
R610 B.n618 B.n315 163.367
R611 B.n622 B.n315 163.367
R612 B.n622 B.n309 163.367
R613 B.n630 B.n309 163.367
R614 B.n630 B.n307 163.367
R615 B.n634 B.n307 163.367
R616 B.n634 B.n301 163.367
R617 B.n642 B.n301 163.367
R618 B.n642 B.n299 163.367
R619 B.n647 B.n299 163.367
R620 B.n647 B.n293 163.367
R621 B.n655 B.n293 163.367
R622 B.n656 B.n655 163.367
R623 B.n656 B.n5 163.367
R624 B.n6 B.n5 163.367
R625 B.n7 B.n6 163.367
R626 B.n661 B.n7 163.367
R627 B.n661 B.n12 163.367
R628 B.n13 B.n12 163.367
R629 B.n14 B.n13 163.367
R630 B.n666 B.n14 163.367
R631 B.n666 B.n19 163.367
R632 B.n20 B.n19 163.367
R633 B.n21 B.n20 163.367
R634 B.n671 B.n21 163.367
R635 B.n671 B.n26 163.367
R636 B.n27 B.n26 163.367
R637 B.n28 B.n27 163.367
R638 B.n676 B.n28 163.367
R639 B.n676 B.n33 163.367
R640 B.n34 B.n33 163.367
R641 B.n35 B.n34 163.367
R642 B.n681 B.n35 163.367
R643 B.n681 B.n40 163.367
R644 B.n41 B.n40 163.367
R645 B.n42 B.n41 163.367
R646 B.n686 B.n42 163.367
R647 B.n686 B.n47 163.367
R648 B.n104 B.n103 163.367
R649 B.n108 B.n107 163.367
R650 B.n112 B.n111 163.367
R651 B.n116 B.n115 163.367
R652 B.n120 B.n119 163.367
R653 B.n124 B.n123 163.367
R654 B.n128 B.n127 163.367
R655 B.n132 B.n131 163.367
R656 B.n136 B.n135 163.367
R657 B.n140 B.n139 163.367
R658 B.n144 B.n143 163.367
R659 B.n148 B.n147 163.367
R660 B.n152 B.n151 163.367
R661 B.n156 B.n155 163.367
R662 B.n160 B.n159 163.367
R663 B.n164 B.n163 163.367
R664 B.n168 B.n167 163.367
R665 B.n172 B.n171 163.367
R666 B.n176 B.n175 163.367
R667 B.n180 B.n179 163.367
R668 B.n184 B.n183 163.367
R669 B.n188 B.n187 163.367
R670 B.n192 B.n191 163.367
R671 B.n196 B.n195 163.367
R672 B.n200 B.n199 163.367
R673 B.n204 B.n203 163.367
R674 B.n209 B.n208 163.367
R675 B.n213 B.n212 163.367
R676 B.n217 B.n216 163.367
R677 B.n221 B.n220 163.367
R678 B.n225 B.n224 163.367
R679 B.n229 B.n228 163.367
R680 B.n233 B.n232 163.367
R681 B.n237 B.n236 163.367
R682 B.n241 B.n240 163.367
R683 B.n245 B.n244 163.367
R684 B.n249 B.n248 163.367
R685 B.n253 B.n252 163.367
R686 B.n257 B.n256 163.367
R687 B.n261 B.n260 163.367
R688 B.n265 B.n264 163.367
R689 B.n269 B.n268 163.367
R690 B.n273 B.n272 163.367
R691 B.n277 B.n276 163.367
R692 B.n281 B.n280 163.367
R693 B.n285 B.n284 163.367
R694 B.n289 B.n288 163.367
R695 B.n690 B.n96 163.367
R696 B.n587 B.n338 84.6393
R697 B.n692 B.n691 84.6393
R698 B.n392 B.n337 71.676
R699 B.n396 B.n395 71.676
R700 B.n401 B.n400 71.676
R701 B.n404 B.n403 71.676
R702 B.n409 B.n408 71.676
R703 B.n412 B.n411 71.676
R704 B.n417 B.n416 71.676
R705 B.n420 B.n419 71.676
R706 B.n425 B.n424 71.676
R707 B.n428 B.n427 71.676
R708 B.n433 B.n432 71.676
R709 B.n436 B.n435 71.676
R710 B.n441 B.n440 71.676
R711 B.n444 B.n443 71.676
R712 B.n449 B.n448 71.676
R713 B.n452 B.n451 71.676
R714 B.n457 B.n456 71.676
R715 B.n460 B.n459 71.676
R716 B.n465 B.n464 71.676
R717 B.n468 B.n467 71.676
R718 B.n473 B.n472 71.676
R719 B.n476 B.n475 71.676
R720 B.n482 B.n481 71.676
R721 B.n485 B.n484 71.676
R722 B.n490 B.n489 71.676
R723 B.n493 B.n492 71.676
R724 B.n499 B.n498 71.676
R725 B.n502 B.n501 71.676
R726 B.n507 B.n506 71.676
R727 B.n510 B.n509 71.676
R728 B.n515 B.n514 71.676
R729 B.n518 B.n517 71.676
R730 B.n523 B.n522 71.676
R731 B.n526 B.n525 71.676
R732 B.n531 B.n530 71.676
R733 B.n534 B.n533 71.676
R734 B.n539 B.n538 71.676
R735 B.n542 B.n541 71.676
R736 B.n547 B.n546 71.676
R737 B.n550 B.n549 71.676
R738 B.n555 B.n554 71.676
R739 B.n558 B.n557 71.676
R740 B.n563 B.n562 71.676
R741 B.n566 B.n565 71.676
R742 B.n571 B.n570 71.676
R743 B.n574 B.n573 71.676
R744 B.n579 B.n578 71.676
R745 B.n582 B.n581 71.676
R746 B.n48 B.n46 71.676
R747 B.n104 B.n49 71.676
R748 B.n108 B.n50 71.676
R749 B.n112 B.n51 71.676
R750 B.n116 B.n52 71.676
R751 B.n120 B.n53 71.676
R752 B.n124 B.n54 71.676
R753 B.n128 B.n55 71.676
R754 B.n132 B.n56 71.676
R755 B.n136 B.n57 71.676
R756 B.n140 B.n58 71.676
R757 B.n144 B.n59 71.676
R758 B.n148 B.n60 71.676
R759 B.n152 B.n61 71.676
R760 B.n156 B.n62 71.676
R761 B.n160 B.n63 71.676
R762 B.n164 B.n64 71.676
R763 B.n168 B.n65 71.676
R764 B.n172 B.n66 71.676
R765 B.n176 B.n67 71.676
R766 B.n180 B.n68 71.676
R767 B.n184 B.n69 71.676
R768 B.n188 B.n70 71.676
R769 B.n192 B.n71 71.676
R770 B.n196 B.n72 71.676
R771 B.n200 B.n73 71.676
R772 B.n204 B.n74 71.676
R773 B.n209 B.n75 71.676
R774 B.n213 B.n76 71.676
R775 B.n217 B.n77 71.676
R776 B.n221 B.n78 71.676
R777 B.n225 B.n79 71.676
R778 B.n229 B.n80 71.676
R779 B.n233 B.n81 71.676
R780 B.n237 B.n82 71.676
R781 B.n241 B.n83 71.676
R782 B.n245 B.n84 71.676
R783 B.n249 B.n85 71.676
R784 B.n253 B.n86 71.676
R785 B.n257 B.n87 71.676
R786 B.n261 B.n88 71.676
R787 B.n265 B.n89 71.676
R788 B.n269 B.n90 71.676
R789 B.n273 B.n91 71.676
R790 B.n277 B.n92 71.676
R791 B.n281 B.n93 71.676
R792 B.n285 B.n94 71.676
R793 B.n289 B.n95 71.676
R794 B.n96 B.n95 71.676
R795 B.n288 B.n94 71.676
R796 B.n284 B.n93 71.676
R797 B.n280 B.n92 71.676
R798 B.n276 B.n91 71.676
R799 B.n272 B.n90 71.676
R800 B.n268 B.n89 71.676
R801 B.n264 B.n88 71.676
R802 B.n260 B.n87 71.676
R803 B.n256 B.n86 71.676
R804 B.n252 B.n85 71.676
R805 B.n248 B.n84 71.676
R806 B.n244 B.n83 71.676
R807 B.n240 B.n82 71.676
R808 B.n236 B.n81 71.676
R809 B.n232 B.n80 71.676
R810 B.n228 B.n79 71.676
R811 B.n224 B.n78 71.676
R812 B.n220 B.n77 71.676
R813 B.n216 B.n76 71.676
R814 B.n212 B.n75 71.676
R815 B.n208 B.n74 71.676
R816 B.n203 B.n73 71.676
R817 B.n199 B.n72 71.676
R818 B.n195 B.n71 71.676
R819 B.n191 B.n70 71.676
R820 B.n187 B.n69 71.676
R821 B.n183 B.n68 71.676
R822 B.n179 B.n67 71.676
R823 B.n175 B.n66 71.676
R824 B.n171 B.n65 71.676
R825 B.n167 B.n64 71.676
R826 B.n163 B.n63 71.676
R827 B.n159 B.n62 71.676
R828 B.n155 B.n61 71.676
R829 B.n151 B.n60 71.676
R830 B.n147 B.n59 71.676
R831 B.n143 B.n58 71.676
R832 B.n139 B.n57 71.676
R833 B.n135 B.n56 71.676
R834 B.n131 B.n55 71.676
R835 B.n127 B.n54 71.676
R836 B.n123 B.n53 71.676
R837 B.n119 B.n52 71.676
R838 B.n115 B.n51 71.676
R839 B.n111 B.n50 71.676
R840 B.n107 B.n49 71.676
R841 B.n103 B.n48 71.676
R842 B.n393 B.n392 71.676
R843 B.n395 B.n389 71.676
R844 B.n402 B.n401 71.676
R845 B.n403 B.n387 71.676
R846 B.n410 B.n409 71.676
R847 B.n411 B.n385 71.676
R848 B.n418 B.n417 71.676
R849 B.n419 B.n383 71.676
R850 B.n426 B.n425 71.676
R851 B.n427 B.n381 71.676
R852 B.n434 B.n433 71.676
R853 B.n435 B.n379 71.676
R854 B.n442 B.n441 71.676
R855 B.n443 B.n377 71.676
R856 B.n450 B.n449 71.676
R857 B.n451 B.n375 71.676
R858 B.n458 B.n457 71.676
R859 B.n459 B.n373 71.676
R860 B.n466 B.n465 71.676
R861 B.n467 B.n371 71.676
R862 B.n474 B.n473 71.676
R863 B.n475 B.n367 71.676
R864 B.n483 B.n482 71.676
R865 B.n484 B.n365 71.676
R866 B.n491 B.n490 71.676
R867 B.n492 B.n361 71.676
R868 B.n500 B.n499 71.676
R869 B.n501 B.n359 71.676
R870 B.n508 B.n507 71.676
R871 B.n509 B.n357 71.676
R872 B.n516 B.n515 71.676
R873 B.n517 B.n355 71.676
R874 B.n524 B.n523 71.676
R875 B.n525 B.n353 71.676
R876 B.n532 B.n531 71.676
R877 B.n533 B.n351 71.676
R878 B.n540 B.n539 71.676
R879 B.n541 B.n349 71.676
R880 B.n548 B.n547 71.676
R881 B.n549 B.n347 71.676
R882 B.n556 B.n555 71.676
R883 B.n557 B.n345 71.676
R884 B.n564 B.n563 71.676
R885 B.n565 B.n343 71.676
R886 B.n572 B.n571 71.676
R887 B.n573 B.n341 71.676
R888 B.n580 B.n579 71.676
R889 B.n581 B.n339 71.676
R890 B.n496 B.n363 59.5399
R891 B.n478 B.n369 59.5399
R892 B.n101 B.n100 59.5399
R893 B.n206 B.n98 59.5399
R894 B.n363 B.n362 53.1399
R895 B.n369 B.n368 53.1399
R896 B.n100 B.n99 53.1399
R897 B.n98 B.n97 53.1399
R898 B.n587 B.n334 41.4065
R899 B.n593 B.n334 41.4065
R900 B.n593 B.n330 41.4065
R901 B.n599 B.n330 41.4065
R902 B.n599 B.n325 41.4065
R903 B.n605 B.n325 41.4065
R904 B.n605 B.n326 41.4065
R905 B.n611 B.n318 41.4065
R906 B.n617 B.n318 41.4065
R907 B.n617 B.n314 41.4065
R908 B.n623 B.n314 41.4065
R909 B.n623 B.n310 41.4065
R910 B.n629 B.n310 41.4065
R911 B.n629 B.n306 41.4065
R912 B.n635 B.n306 41.4065
R913 B.n635 B.n302 41.4065
R914 B.n641 B.n302 41.4065
R915 B.n648 B.n298 41.4065
R916 B.n648 B.n294 41.4065
R917 B.n654 B.n294 41.4065
R918 B.n654 B.n4 41.4065
R919 B.n740 B.n4 41.4065
R920 B.n740 B.n739 41.4065
R921 B.n739 B.n738 41.4065
R922 B.n738 B.n8 41.4065
R923 B.n732 B.n8 41.4065
R924 B.n732 B.n731 41.4065
R925 B.n730 B.n15 41.4065
R926 B.n724 B.n15 41.4065
R927 B.n724 B.n723 41.4065
R928 B.n723 B.n722 41.4065
R929 B.n722 B.n22 41.4065
R930 B.n716 B.n22 41.4065
R931 B.n716 B.n715 41.4065
R932 B.n715 B.n714 41.4065
R933 B.n714 B.n29 41.4065
R934 B.n708 B.n29 41.4065
R935 B.n707 B.n706 41.4065
R936 B.n706 B.n36 41.4065
R937 B.n700 B.n36 41.4065
R938 B.n700 B.n699 41.4065
R939 B.n699 B.n698 41.4065
R940 B.n698 B.n43 41.4065
R941 B.n692 B.n43 41.4065
R942 B.n694 B.n45 37.3078
R943 B.n689 B.n688 37.3078
R944 B.n585 B.n584 37.3078
R945 B.n589 B.n336 37.3078
R946 B.n611 B.t7 37.1442
R947 B.n708 B.t3 37.1442
R948 B.t0 B.n298 26.1837
R949 B.n731 B.t1 26.1837
R950 B B.n742 18.0485
R951 B.n641 B.t0 15.2233
R952 B.t1 B.n730 15.2233
R953 B.n102 B.n45 10.6151
R954 B.n105 B.n102 10.6151
R955 B.n106 B.n105 10.6151
R956 B.n109 B.n106 10.6151
R957 B.n110 B.n109 10.6151
R958 B.n113 B.n110 10.6151
R959 B.n114 B.n113 10.6151
R960 B.n117 B.n114 10.6151
R961 B.n118 B.n117 10.6151
R962 B.n121 B.n118 10.6151
R963 B.n122 B.n121 10.6151
R964 B.n125 B.n122 10.6151
R965 B.n126 B.n125 10.6151
R966 B.n129 B.n126 10.6151
R967 B.n130 B.n129 10.6151
R968 B.n133 B.n130 10.6151
R969 B.n134 B.n133 10.6151
R970 B.n137 B.n134 10.6151
R971 B.n138 B.n137 10.6151
R972 B.n141 B.n138 10.6151
R973 B.n142 B.n141 10.6151
R974 B.n145 B.n142 10.6151
R975 B.n146 B.n145 10.6151
R976 B.n149 B.n146 10.6151
R977 B.n150 B.n149 10.6151
R978 B.n153 B.n150 10.6151
R979 B.n154 B.n153 10.6151
R980 B.n157 B.n154 10.6151
R981 B.n158 B.n157 10.6151
R982 B.n161 B.n158 10.6151
R983 B.n162 B.n161 10.6151
R984 B.n165 B.n162 10.6151
R985 B.n166 B.n165 10.6151
R986 B.n169 B.n166 10.6151
R987 B.n170 B.n169 10.6151
R988 B.n173 B.n170 10.6151
R989 B.n174 B.n173 10.6151
R990 B.n177 B.n174 10.6151
R991 B.n178 B.n177 10.6151
R992 B.n181 B.n178 10.6151
R993 B.n182 B.n181 10.6151
R994 B.n185 B.n182 10.6151
R995 B.n186 B.n185 10.6151
R996 B.n190 B.n189 10.6151
R997 B.n193 B.n190 10.6151
R998 B.n194 B.n193 10.6151
R999 B.n197 B.n194 10.6151
R1000 B.n198 B.n197 10.6151
R1001 B.n201 B.n198 10.6151
R1002 B.n202 B.n201 10.6151
R1003 B.n205 B.n202 10.6151
R1004 B.n210 B.n207 10.6151
R1005 B.n211 B.n210 10.6151
R1006 B.n214 B.n211 10.6151
R1007 B.n215 B.n214 10.6151
R1008 B.n218 B.n215 10.6151
R1009 B.n219 B.n218 10.6151
R1010 B.n222 B.n219 10.6151
R1011 B.n223 B.n222 10.6151
R1012 B.n226 B.n223 10.6151
R1013 B.n227 B.n226 10.6151
R1014 B.n230 B.n227 10.6151
R1015 B.n231 B.n230 10.6151
R1016 B.n234 B.n231 10.6151
R1017 B.n235 B.n234 10.6151
R1018 B.n238 B.n235 10.6151
R1019 B.n239 B.n238 10.6151
R1020 B.n242 B.n239 10.6151
R1021 B.n243 B.n242 10.6151
R1022 B.n246 B.n243 10.6151
R1023 B.n247 B.n246 10.6151
R1024 B.n250 B.n247 10.6151
R1025 B.n251 B.n250 10.6151
R1026 B.n254 B.n251 10.6151
R1027 B.n255 B.n254 10.6151
R1028 B.n258 B.n255 10.6151
R1029 B.n259 B.n258 10.6151
R1030 B.n262 B.n259 10.6151
R1031 B.n263 B.n262 10.6151
R1032 B.n266 B.n263 10.6151
R1033 B.n267 B.n266 10.6151
R1034 B.n270 B.n267 10.6151
R1035 B.n271 B.n270 10.6151
R1036 B.n274 B.n271 10.6151
R1037 B.n275 B.n274 10.6151
R1038 B.n278 B.n275 10.6151
R1039 B.n279 B.n278 10.6151
R1040 B.n282 B.n279 10.6151
R1041 B.n283 B.n282 10.6151
R1042 B.n286 B.n283 10.6151
R1043 B.n287 B.n286 10.6151
R1044 B.n290 B.n287 10.6151
R1045 B.n291 B.n290 10.6151
R1046 B.n689 B.n291 10.6151
R1047 B.n585 B.n332 10.6151
R1048 B.n595 B.n332 10.6151
R1049 B.n596 B.n595 10.6151
R1050 B.n597 B.n596 10.6151
R1051 B.n597 B.n323 10.6151
R1052 B.n607 B.n323 10.6151
R1053 B.n608 B.n607 10.6151
R1054 B.n609 B.n608 10.6151
R1055 B.n609 B.n316 10.6151
R1056 B.n619 B.n316 10.6151
R1057 B.n620 B.n619 10.6151
R1058 B.n621 B.n620 10.6151
R1059 B.n621 B.n308 10.6151
R1060 B.n631 B.n308 10.6151
R1061 B.n632 B.n631 10.6151
R1062 B.n633 B.n632 10.6151
R1063 B.n633 B.n300 10.6151
R1064 B.n643 B.n300 10.6151
R1065 B.n644 B.n643 10.6151
R1066 B.n646 B.n644 10.6151
R1067 B.n646 B.n645 10.6151
R1068 B.n645 B.n292 10.6151
R1069 B.n657 B.n292 10.6151
R1070 B.n658 B.n657 10.6151
R1071 B.n659 B.n658 10.6151
R1072 B.n660 B.n659 10.6151
R1073 B.n662 B.n660 10.6151
R1074 B.n663 B.n662 10.6151
R1075 B.n664 B.n663 10.6151
R1076 B.n665 B.n664 10.6151
R1077 B.n667 B.n665 10.6151
R1078 B.n668 B.n667 10.6151
R1079 B.n669 B.n668 10.6151
R1080 B.n670 B.n669 10.6151
R1081 B.n672 B.n670 10.6151
R1082 B.n673 B.n672 10.6151
R1083 B.n674 B.n673 10.6151
R1084 B.n675 B.n674 10.6151
R1085 B.n677 B.n675 10.6151
R1086 B.n678 B.n677 10.6151
R1087 B.n679 B.n678 10.6151
R1088 B.n680 B.n679 10.6151
R1089 B.n682 B.n680 10.6151
R1090 B.n683 B.n682 10.6151
R1091 B.n684 B.n683 10.6151
R1092 B.n685 B.n684 10.6151
R1093 B.n687 B.n685 10.6151
R1094 B.n688 B.n687 10.6151
R1095 B.n391 B.n336 10.6151
R1096 B.n391 B.n390 10.6151
R1097 B.n397 B.n390 10.6151
R1098 B.n398 B.n397 10.6151
R1099 B.n399 B.n398 10.6151
R1100 B.n399 B.n388 10.6151
R1101 B.n405 B.n388 10.6151
R1102 B.n406 B.n405 10.6151
R1103 B.n407 B.n406 10.6151
R1104 B.n407 B.n386 10.6151
R1105 B.n413 B.n386 10.6151
R1106 B.n414 B.n413 10.6151
R1107 B.n415 B.n414 10.6151
R1108 B.n415 B.n384 10.6151
R1109 B.n421 B.n384 10.6151
R1110 B.n422 B.n421 10.6151
R1111 B.n423 B.n422 10.6151
R1112 B.n423 B.n382 10.6151
R1113 B.n429 B.n382 10.6151
R1114 B.n430 B.n429 10.6151
R1115 B.n431 B.n430 10.6151
R1116 B.n431 B.n380 10.6151
R1117 B.n437 B.n380 10.6151
R1118 B.n438 B.n437 10.6151
R1119 B.n439 B.n438 10.6151
R1120 B.n439 B.n378 10.6151
R1121 B.n445 B.n378 10.6151
R1122 B.n446 B.n445 10.6151
R1123 B.n447 B.n446 10.6151
R1124 B.n447 B.n376 10.6151
R1125 B.n453 B.n376 10.6151
R1126 B.n454 B.n453 10.6151
R1127 B.n455 B.n454 10.6151
R1128 B.n455 B.n374 10.6151
R1129 B.n461 B.n374 10.6151
R1130 B.n462 B.n461 10.6151
R1131 B.n463 B.n462 10.6151
R1132 B.n463 B.n372 10.6151
R1133 B.n469 B.n372 10.6151
R1134 B.n470 B.n469 10.6151
R1135 B.n471 B.n470 10.6151
R1136 B.n471 B.n370 10.6151
R1137 B.n477 B.n370 10.6151
R1138 B.n480 B.n479 10.6151
R1139 B.n480 B.n366 10.6151
R1140 B.n486 B.n366 10.6151
R1141 B.n487 B.n486 10.6151
R1142 B.n488 B.n487 10.6151
R1143 B.n488 B.n364 10.6151
R1144 B.n494 B.n364 10.6151
R1145 B.n495 B.n494 10.6151
R1146 B.n497 B.n360 10.6151
R1147 B.n503 B.n360 10.6151
R1148 B.n504 B.n503 10.6151
R1149 B.n505 B.n504 10.6151
R1150 B.n505 B.n358 10.6151
R1151 B.n511 B.n358 10.6151
R1152 B.n512 B.n511 10.6151
R1153 B.n513 B.n512 10.6151
R1154 B.n513 B.n356 10.6151
R1155 B.n519 B.n356 10.6151
R1156 B.n520 B.n519 10.6151
R1157 B.n521 B.n520 10.6151
R1158 B.n521 B.n354 10.6151
R1159 B.n527 B.n354 10.6151
R1160 B.n528 B.n527 10.6151
R1161 B.n529 B.n528 10.6151
R1162 B.n529 B.n352 10.6151
R1163 B.n535 B.n352 10.6151
R1164 B.n536 B.n535 10.6151
R1165 B.n537 B.n536 10.6151
R1166 B.n537 B.n350 10.6151
R1167 B.n543 B.n350 10.6151
R1168 B.n544 B.n543 10.6151
R1169 B.n545 B.n544 10.6151
R1170 B.n545 B.n348 10.6151
R1171 B.n551 B.n348 10.6151
R1172 B.n552 B.n551 10.6151
R1173 B.n553 B.n552 10.6151
R1174 B.n553 B.n346 10.6151
R1175 B.n559 B.n346 10.6151
R1176 B.n560 B.n559 10.6151
R1177 B.n561 B.n560 10.6151
R1178 B.n561 B.n344 10.6151
R1179 B.n567 B.n344 10.6151
R1180 B.n568 B.n567 10.6151
R1181 B.n569 B.n568 10.6151
R1182 B.n569 B.n342 10.6151
R1183 B.n575 B.n342 10.6151
R1184 B.n576 B.n575 10.6151
R1185 B.n577 B.n576 10.6151
R1186 B.n577 B.n340 10.6151
R1187 B.n583 B.n340 10.6151
R1188 B.n584 B.n583 10.6151
R1189 B.n590 B.n589 10.6151
R1190 B.n591 B.n590 10.6151
R1191 B.n591 B.n328 10.6151
R1192 B.n601 B.n328 10.6151
R1193 B.n602 B.n601 10.6151
R1194 B.n603 B.n602 10.6151
R1195 B.n603 B.n320 10.6151
R1196 B.n613 B.n320 10.6151
R1197 B.n614 B.n613 10.6151
R1198 B.n615 B.n614 10.6151
R1199 B.n615 B.n312 10.6151
R1200 B.n625 B.n312 10.6151
R1201 B.n626 B.n625 10.6151
R1202 B.n627 B.n626 10.6151
R1203 B.n627 B.n304 10.6151
R1204 B.n637 B.n304 10.6151
R1205 B.n638 B.n637 10.6151
R1206 B.n639 B.n638 10.6151
R1207 B.n639 B.n296 10.6151
R1208 B.n650 B.n296 10.6151
R1209 B.n651 B.n650 10.6151
R1210 B.n652 B.n651 10.6151
R1211 B.n652 B.n0 10.6151
R1212 B.n736 B.n1 10.6151
R1213 B.n736 B.n735 10.6151
R1214 B.n735 B.n734 10.6151
R1215 B.n734 B.n10 10.6151
R1216 B.n728 B.n10 10.6151
R1217 B.n728 B.n727 10.6151
R1218 B.n727 B.n726 10.6151
R1219 B.n726 B.n17 10.6151
R1220 B.n720 B.n17 10.6151
R1221 B.n720 B.n719 10.6151
R1222 B.n719 B.n718 10.6151
R1223 B.n718 B.n24 10.6151
R1224 B.n712 B.n24 10.6151
R1225 B.n712 B.n711 10.6151
R1226 B.n711 B.n710 10.6151
R1227 B.n710 B.n31 10.6151
R1228 B.n704 B.n31 10.6151
R1229 B.n704 B.n703 10.6151
R1230 B.n703 B.n702 10.6151
R1231 B.n702 B.n38 10.6151
R1232 B.n696 B.n38 10.6151
R1233 B.n696 B.n695 10.6151
R1234 B.n695 B.n694 10.6151
R1235 B.n189 B.n101 6.5566
R1236 B.n206 B.n205 6.5566
R1237 B.n479 B.n478 6.5566
R1238 B.n496 B.n495 6.5566
R1239 B.n326 B.t7 4.26289
R1240 B.t3 B.n707 4.26289
R1241 B.n186 B.n101 4.05904
R1242 B.n207 B.n206 4.05904
R1243 B.n478 B.n477 4.05904
R1244 B.n497 B.n496 4.05904
R1245 B.n742 B.n0 2.81026
R1246 B.n742 B.n1 2.81026
R1247 VN VN.t1 221.918
R1248 VN VN.t0 177.407
R1249 VTAIL.n274 VTAIL.n210 289.615
R1250 VTAIL.n64 VTAIL.n0 289.615
R1251 VTAIL.n204 VTAIL.n140 289.615
R1252 VTAIL.n134 VTAIL.n70 289.615
R1253 VTAIL.n233 VTAIL.n232 185
R1254 VTAIL.n230 VTAIL.n229 185
R1255 VTAIL.n239 VTAIL.n238 185
R1256 VTAIL.n241 VTAIL.n240 185
R1257 VTAIL.n226 VTAIL.n225 185
R1258 VTAIL.n247 VTAIL.n246 185
R1259 VTAIL.n250 VTAIL.n249 185
R1260 VTAIL.n248 VTAIL.n222 185
R1261 VTAIL.n255 VTAIL.n221 185
R1262 VTAIL.n257 VTAIL.n256 185
R1263 VTAIL.n259 VTAIL.n258 185
R1264 VTAIL.n218 VTAIL.n217 185
R1265 VTAIL.n265 VTAIL.n264 185
R1266 VTAIL.n267 VTAIL.n266 185
R1267 VTAIL.n214 VTAIL.n213 185
R1268 VTAIL.n273 VTAIL.n272 185
R1269 VTAIL.n275 VTAIL.n274 185
R1270 VTAIL.n23 VTAIL.n22 185
R1271 VTAIL.n20 VTAIL.n19 185
R1272 VTAIL.n29 VTAIL.n28 185
R1273 VTAIL.n31 VTAIL.n30 185
R1274 VTAIL.n16 VTAIL.n15 185
R1275 VTAIL.n37 VTAIL.n36 185
R1276 VTAIL.n40 VTAIL.n39 185
R1277 VTAIL.n38 VTAIL.n12 185
R1278 VTAIL.n45 VTAIL.n11 185
R1279 VTAIL.n47 VTAIL.n46 185
R1280 VTAIL.n49 VTAIL.n48 185
R1281 VTAIL.n8 VTAIL.n7 185
R1282 VTAIL.n55 VTAIL.n54 185
R1283 VTAIL.n57 VTAIL.n56 185
R1284 VTAIL.n4 VTAIL.n3 185
R1285 VTAIL.n63 VTAIL.n62 185
R1286 VTAIL.n65 VTAIL.n64 185
R1287 VTAIL.n205 VTAIL.n204 185
R1288 VTAIL.n203 VTAIL.n202 185
R1289 VTAIL.n144 VTAIL.n143 185
R1290 VTAIL.n197 VTAIL.n196 185
R1291 VTAIL.n195 VTAIL.n194 185
R1292 VTAIL.n148 VTAIL.n147 185
R1293 VTAIL.n189 VTAIL.n188 185
R1294 VTAIL.n187 VTAIL.n186 185
R1295 VTAIL.n185 VTAIL.n151 185
R1296 VTAIL.n155 VTAIL.n152 185
R1297 VTAIL.n180 VTAIL.n179 185
R1298 VTAIL.n178 VTAIL.n177 185
R1299 VTAIL.n157 VTAIL.n156 185
R1300 VTAIL.n172 VTAIL.n171 185
R1301 VTAIL.n170 VTAIL.n169 185
R1302 VTAIL.n161 VTAIL.n160 185
R1303 VTAIL.n164 VTAIL.n163 185
R1304 VTAIL.n135 VTAIL.n134 185
R1305 VTAIL.n133 VTAIL.n132 185
R1306 VTAIL.n74 VTAIL.n73 185
R1307 VTAIL.n127 VTAIL.n126 185
R1308 VTAIL.n125 VTAIL.n124 185
R1309 VTAIL.n78 VTAIL.n77 185
R1310 VTAIL.n119 VTAIL.n118 185
R1311 VTAIL.n117 VTAIL.n116 185
R1312 VTAIL.n115 VTAIL.n81 185
R1313 VTAIL.n85 VTAIL.n82 185
R1314 VTAIL.n110 VTAIL.n109 185
R1315 VTAIL.n108 VTAIL.n107 185
R1316 VTAIL.n87 VTAIL.n86 185
R1317 VTAIL.n102 VTAIL.n101 185
R1318 VTAIL.n100 VTAIL.n99 185
R1319 VTAIL.n91 VTAIL.n90 185
R1320 VTAIL.n94 VTAIL.n93 185
R1321 VTAIL.t3 VTAIL.n231 149.524
R1322 VTAIL.t0 VTAIL.n21 149.524
R1323 VTAIL.t1 VTAIL.n162 149.524
R1324 VTAIL.t2 VTAIL.n92 149.524
R1325 VTAIL.n232 VTAIL.n229 104.615
R1326 VTAIL.n239 VTAIL.n229 104.615
R1327 VTAIL.n240 VTAIL.n239 104.615
R1328 VTAIL.n240 VTAIL.n225 104.615
R1329 VTAIL.n247 VTAIL.n225 104.615
R1330 VTAIL.n249 VTAIL.n247 104.615
R1331 VTAIL.n249 VTAIL.n248 104.615
R1332 VTAIL.n248 VTAIL.n221 104.615
R1333 VTAIL.n257 VTAIL.n221 104.615
R1334 VTAIL.n258 VTAIL.n257 104.615
R1335 VTAIL.n258 VTAIL.n217 104.615
R1336 VTAIL.n265 VTAIL.n217 104.615
R1337 VTAIL.n266 VTAIL.n265 104.615
R1338 VTAIL.n266 VTAIL.n213 104.615
R1339 VTAIL.n273 VTAIL.n213 104.615
R1340 VTAIL.n274 VTAIL.n273 104.615
R1341 VTAIL.n22 VTAIL.n19 104.615
R1342 VTAIL.n29 VTAIL.n19 104.615
R1343 VTAIL.n30 VTAIL.n29 104.615
R1344 VTAIL.n30 VTAIL.n15 104.615
R1345 VTAIL.n37 VTAIL.n15 104.615
R1346 VTAIL.n39 VTAIL.n37 104.615
R1347 VTAIL.n39 VTAIL.n38 104.615
R1348 VTAIL.n38 VTAIL.n11 104.615
R1349 VTAIL.n47 VTAIL.n11 104.615
R1350 VTAIL.n48 VTAIL.n47 104.615
R1351 VTAIL.n48 VTAIL.n7 104.615
R1352 VTAIL.n55 VTAIL.n7 104.615
R1353 VTAIL.n56 VTAIL.n55 104.615
R1354 VTAIL.n56 VTAIL.n3 104.615
R1355 VTAIL.n63 VTAIL.n3 104.615
R1356 VTAIL.n64 VTAIL.n63 104.615
R1357 VTAIL.n204 VTAIL.n203 104.615
R1358 VTAIL.n203 VTAIL.n143 104.615
R1359 VTAIL.n196 VTAIL.n143 104.615
R1360 VTAIL.n196 VTAIL.n195 104.615
R1361 VTAIL.n195 VTAIL.n147 104.615
R1362 VTAIL.n188 VTAIL.n147 104.615
R1363 VTAIL.n188 VTAIL.n187 104.615
R1364 VTAIL.n187 VTAIL.n151 104.615
R1365 VTAIL.n155 VTAIL.n151 104.615
R1366 VTAIL.n179 VTAIL.n155 104.615
R1367 VTAIL.n179 VTAIL.n178 104.615
R1368 VTAIL.n178 VTAIL.n156 104.615
R1369 VTAIL.n171 VTAIL.n156 104.615
R1370 VTAIL.n171 VTAIL.n170 104.615
R1371 VTAIL.n170 VTAIL.n160 104.615
R1372 VTAIL.n163 VTAIL.n160 104.615
R1373 VTAIL.n134 VTAIL.n133 104.615
R1374 VTAIL.n133 VTAIL.n73 104.615
R1375 VTAIL.n126 VTAIL.n73 104.615
R1376 VTAIL.n126 VTAIL.n125 104.615
R1377 VTAIL.n125 VTAIL.n77 104.615
R1378 VTAIL.n118 VTAIL.n77 104.615
R1379 VTAIL.n118 VTAIL.n117 104.615
R1380 VTAIL.n117 VTAIL.n81 104.615
R1381 VTAIL.n85 VTAIL.n81 104.615
R1382 VTAIL.n109 VTAIL.n85 104.615
R1383 VTAIL.n109 VTAIL.n108 104.615
R1384 VTAIL.n108 VTAIL.n86 104.615
R1385 VTAIL.n101 VTAIL.n86 104.615
R1386 VTAIL.n101 VTAIL.n100 104.615
R1387 VTAIL.n100 VTAIL.n90 104.615
R1388 VTAIL.n93 VTAIL.n90 104.615
R1389 VTAIL.n232 VTAIL.t3 52.3082
R1390 VTAIL.n22 VTAIL.t0 52.3082
R1391 VTAIL.n163 VTAIL.t1 52.3082
R1392 VTAIL.n93 VTAIL.t2 52.3082
R1393 VTAIL.n279 VTAIL.n278 31.2157
R1394 VTAIL.n69 VTAIL.n68 31.2157
R1395 VTAIL.n209 VTAIL.n208 31.2157
R1396 VTAIL.n139 VTAIL.n138 31.2157
R1397 VTAIL.n139 VTAIL.n69 28.1169
R1398 VTAIL.n279 VTAIL.n209 25.7548
R1399 VTAIL.n256 VTAIL.n255 13.1884
R1400 VTAIL.n46 VTAIL.n45 13.1884
R1401 VTAIL.n186 VTAIL.n185 13.1884
R1402 VTAIL.n116 VTAIL.n115 13.1884
R1403 VTAIL.n254 VTAIL.n222 12.8005
R1404 VTAIL.n259 VTAIL.n220 12.8005
R1405 VTAIL.n44 VTAIL.n12 12.8005
R1406 VTAIL.n49 VTAIL.n10 12.8005
R1407 VTAIL.n189 VTAIL.n150 12.8005
R1408 VTAIL.n184 VTAIL.n152 12.8005
R1409 VTAIL.n119 VTAIL.n80 12.8005
R1410 VTAIL.n114 VTAIL.n82 12.8005
R1411 VTAIL.n251 VTAIL.n250 12.0247
R1412 VTAIL.n260 VTAIL.n218 12.0247
R1413 VTAIL.n41 VTAIL.n40 12.0247
R1414 VTAIL.n50 VTAIL.n8 12.0247
R1415 VTAIL.n190 VTAIL.n148 12.0247
R1416 VTAIL.n181 VTAIL.n180 12.0247
R1417 VTAIL.n120 VTAIL.n78 12.0247
R1418 VTAIL.n111 VTAIL.n110 12.0247
R1419 VTAIL.n246 VTAIL.n224 11.249
R1420 VTAIL.n264 VTAIL.n263 11.249
R1421 VTAIL.n36 VTAIL.n14 11.249
R1422 VTAIL.n54 VTAIL.n53 11.249
R1423 VTAIL.n194 VTAIL.n193 11.249
R1424 VTAIL.n177 VTAIL.n154 11.249
R1425 VTAIL.n124 VTAIL.n123 11.249
R1426 VTAIL.n107 VTAIL.n84 11.249
R1427 VTAIL.n245 VTAIL.n226 10.4732
R1428 VTAIL.n267 VTAIL.n216 10.4732
R1429 VTAIL.n35 VTAIL.n16 10.4732
R1430 VTAIL.n57 VTAIL.n6 10.4732
R1431 VTAIL.n197 VTAIL.n146 10.4732
R1432 VTAIL.n176 VTAIL.n157 10.4732
R1433 VTAIL.n127 VTAIL.n76 10.4732
R1434 VTAIL.n106 VTAIL.n87 10.4732
R1435 VTAIL.n233 VTAIL.n231 10.2747
R1436 VTAIL.n23 VTAIL.n21 10.2747
R1437 VTAIL.n164 VTAIL.n162 10.2747
R1438 VTAIL.n94 VTAIL.n92 10.2747
R1439 VTAIL.n242 VTAIL.n241 9.69747
R1440 VTAIL.n268 VTAIL.n214 9.69747
R1441 VTAIL.n32 VTAIL.n31 9.69747
R1442 VTAIL.n58 VTAIL.n4 9.69747
R1443 VTAIL.n198 VTAIL.n144 9.69747
R1444 VTAIL.n173 VTAIL.n172 9.69747
R1445 VTAIL.n128 VTAIL.n74 9.69747
R1446 VTAIL.n103 VTAIL.n102 9.69747
R1447 VTAIL.n278 VTAIL.n277 9.45567
R1448 VTAIL.n68 VTAIL.n67 9.45567
R1449 VTAIL.n208 VTAIL.n207 9.45567
R1450 VTAIL.n138 VTAIL.n137 9.45567
R1451 VTAIL.n212 VTAIL.n211 9.3005
R1452 VTAIL.n271 VTAIL.n270 9.3005
R1453 VTAIL.n269 VTAIL.n268 9.3005
R1454 VTAIL.n216 VTAIL.n215 9.3005
R1455 VTAIL.n263 VTAIL.n262 9.3005
R1456 VTAIL.n261 VTAIL.n260 9.3005
R1457 VTAIL.n220 VTAIL.n219 9.3005
R1458 VTAIL.n235 VTAIL.n234 9.3005
R1459 VTAIL.n237 VTAIL.n236 9.3005
R1460 VTAIL.n228 VTAIL.n227 9.3005
R1461 VTAIL.n243 VTAIL.n242 9.3005
R1462 VTAIL.n245 VTAIL.n244 9.3005
R1463 VTAIL.n224 VTAIL.n223 9.3005
R1464 VTAIL.n252 VTAIL.n251 9.3005
R1465 VTAIL.n254 VTAIL.n253 9.3005
R1466 VTAIL.n277 VTAIL.n276 9.3005
R1467 VTAIL.n2 VTAIL.n1 9.3005
R1468 VTAIL.n61 VTAIL.n60 9.3005
R1469 VTAIL.n59 VTAIL.n58 9.3005
R1470 VTAIL.n6 VTAIL.n5 9.3005
R1471 VTAIL.n53 VTAIL.n52 9.3005
R1472 VTAIL.n51 VTAIL.n50 9.3005
R1473 VTAIL.n10 VTAIL.n9 9.3005
R1474 VTAIL.n25 VTAIL.n24 9.3005
R1475 VTAIL.n27 VTAIL.n26 9.3005
R1476 VTAIL.n18 VTAIL.n17 9.3005
R1477 VTAIL.n33 VTAIL.n32 9.3005
R1478 VTAIL.n35 VTAIL.n34 9.3005
R1479 VTAIL.n14 VTAIL.n13 9.3005
R1480 VTAIL.n42 VTAIL.n41 9.3005
R1481 VTAIL.n44 VTAIL.n43 9.3005
R1482 VTAIL.n67 VTAIL.n66 9.3005
R1483 VTAIL.n166 VTAIL.n165 9.3005
R1484 VTAIL.n168 VTAIL.n167 9.3005
R1485 VTAIL.n159 VTAIL.n158 9.3005
R1486 VTAIL.n174 VTAIL.n173 9.3005
R1487 VTAIL.n176 VTAIL.n175 9.3005
R1488 VTAIL.n154 VTAIL.n153 9.3005
R1489 VTAIL.n182 VTAIL.n181 9.3005
R1490 VTAIL.n184 VTAIL.n183 9.3005
R1491 VTAIL.n207 VTAIL.n206 9.3005
R1492 VTAIL.n142 VTAIL.n141 9.3005
R1493 VTAIL.n201 VTAIL.n200 9.3005
R1494 VTAIL.n199 VTAIL.n198 9.3005
R1495 VTAIL.n146 VTAIL.n145 9.3005
R1496 VTAIL.n193 VTAIL.n192 9.3005
R1497 VTAIL.n191 VTAIL.n190 9.3005
R1498 VTAIL.n150 VTAIL.n149 9.3005
R1499 VTAIL.n96 VTAIL.n95 9.3005
R1500 VTAIL.n98 VTAIL.n97 9.3005
R1501 VTAIL.n89 VTAIL.n88 9.3005
R1502 VTAIL.n104 VTAIL.n103 9.3005
R1503 VTAIL.n106 VTAIL.n105 9.3005
R1504 VTAIL.n84 VTAIL.n83 9.3005
R1505 VTAIL.n112 VTAIL.n111 9.3005
R1506 VTAIL.n114 VTAIL.n113 9.3005
R1507 VTAIL.n137 VTAIL.n136 9.3005
R1508 VTAIL.n72 VTAIL.n71 9.3005
R1509 VTAIL.n131 VTAIL.n130 9.3005
R1510 VTAIL.n129 VTAIL.n128 9.3005
R1511 VTAIL.n76 VTAIL.n75 9.3005
R1512 VTAIL.n123 VTAIL.n122 9.3005
R1513 VTAIL.n121 VTAIL.n120 9.3005
R1514 VTAIL.n80 VTAIL.n79 9.3005
R1515 VTAIL.n238 VTAIL.n228 8.92171
R1516 VTAIL.n272 VTAIL.n271 8.92171
R1517 VTAIL.n28 VTAIL.n18 8.92171
R1518 VTAIL.n62 VTAIL.n61 8.92171
R1519 VTAIL.n202 VTAIL.n201 8.92171
R1520 VTAIL.n169 VTAIL.n159 8.92171
R1521 VTAIL.n132 VTAIL.n131 8.92171
R1522 VTAIL.n99 VTAIL.n89 8.92171
R1523 VTAIL.n237 VTAIL.n230 8.14595
R1524 VTAIL.n275 VTAIL.n212 8.14595
R1525 VTAIL.n27 VTAIL.n20 8.14595
R1526 VTAIL.n65 VTAIL.n2 8.14595
R1527 VTAIL.n205 VTAIL.n142 8.14595
R1528 VTAIL.n168 VTAIL.n161 8.14595
R1529 VTAIL.n135 VTAIL.n72 8.14595
R1530 VTAIL.n98 VTAIL.n91 8.14595
R1531 VTAIL.n234 VTAIL.n233 7.3702
R1532 VTAIL.n276 VTAIL.n210 7.3702
R1533 VTAIL.n24 VTAIL.n23 7.3702
R1534 VTAIL.n66 VTAIL.n0 7.3702
R1535 VTAIL.n206 VTAIL.n140 7.3702
R1536 VTAIL.n165 VTAIL.n164 7.3702
R1537 VTAIL.n136 VTAIL.n70 7.3702
R1538 VTAIL.n95 VTAIL.n94 7.3702
R1539 VTAIL.n278 VTAIL.n210 6.59444
R1540 VTAIL.n68 VTAIL.n0 6.59444
R1541 VTAIL.n208 VTAIL.n140 6.59444
R1542 VTAIL.n138 VTAIL.n70 6.59444
R1543 VTAIL.n234 VTAIL.n230 5.81868
R1544 VTAIL.n276 VTAIL.n275 5.81868
R1545 VTAIL.n24 VTAIL.n20 5.81868
R1546 VTAIL.n66 VTAIL.n65 5.81868
R1547 VTAIL.n206 VTAIL.n205 5.81868
R1548 VTAIL.n165 VTAIL.n161 5.81868
R1549 VTAIL.n136 VTAIL.n135 5.81868
R1550 VTAIL.n95 VTAIL.n91 5.81868
R1551 VTAIL.n238 VTAIL.n237 5.04292
R1552 VTAIL.n272 VTAIL.n212 5.04292
R1553 VTAIL.n28 VTAIL.n27 5.04292
R1554 VTAIL.n62 VTAIL.n2 5.04292
R1555 VTAIL.n202 VTAIL.n142 5.04292
R1556 VTAIL.n169 VTAIL.n168 5.04292
R1557 VTAIL.n132 VTAIL.n72 5.04292
R1558 VTAIL.n99 VTAIL.n98 5.04292
R1559 VTAIL.n241 VTAIL.n228 4.26717
R1560 VTAIL.n271 VTAIL.n214 4.26717
R1561 VTAIL.n31 VTAIL.n18 4.26717
R1562 VTAIL.n61 VTAIL.n4 4.26717
R1563 VTAIL.n201 VTAIL.n144 4.26717
R1564 VTAIL.n172 VTAIL.n159 4.26717
R1565 VTAIL.n131 VTAIL.n74 4.26717
R1566 VTAIL.n102 VTAIL.n89 4.26717
R1567 VTAIL.n242 VTAIL.n226 3.49141
R1568 VTAIL.n268 VTAIL.n267 3.49141
R1569 VTAIL.n32 VTAIL.n16 3.49141
R1570 VTAIL.n58 VTAIL.n57 3.49141
R1571 VTAIL.n198 VTAIL.n197 3.49141
R1572 VTAIL.n173 VTAIL.n157 3.49141
R1573 VTAIL.n128 VTAIL.n127 3.49141
R1574 VTAIL.n103 VTAIL.n87 3.49141
R1575 VTAIL.n235 VTAIL.n231 2.84303
R1576 VTAIL.n25 VTAIL.n21 2.84303
R1577 VTAIL.n166 VTAIL.n162 2.84303
R1578 VTAIL.n96 VTAIL.n92 2.84303
R1579 VTAIL.n246 VTAIL.n245 2.71565
R1580 VTAIL.n264 VTAIL.n216 2.71565
R1581 VTAIL.n36 VTAIL.n35 2.71565
R1582 VTAIL.n54 VTAIL.n6 2.71565
R1583 VTAIL.n194 VTAIL.n146 2.71565
R1584 VTAIL.n177 VTAIL.n176 2.71565
R1585 VTAIL.n124 VTAIL.n76 2.71565
R1586 VTAIL.n107 VTAIL.n106 2.71565
R1587 VTAIL.n250 VTAIL.n224 1.93989
R1588 VTAIL.n263 VTAIL.n218 1.93989
R1589 VTAIL.n40 VTAIL.n14 1.93989
R1590 VTAIL.n53 VTAIL.n8 1.93989
R1591 VTAIL.n193 VTAIL.n148 1.93989
R1592 VTAIL.n180 VTAIL.n154 1.93989
R1593 VTAIL.n123 VTAIL.n78 1.93989
R1594 VTAIL.n110 VTAIL.n84 1.93989
R1595 VTAIL.n209 VTAIL.n139 1.65136
R1596 VTAIL.n251 VTAIL.n222 1.16414
R1597 VTAIL.n260 VTAIL.n259 1.16414
R1598 VTAIL.n41 VTAIL.n12 1.16414
R1599 VTAIL.n50 VTAIL.n49 1.16414
R1600 VTAIL.n190 VTAIL.n189 1.16414
R1601 VTAIL.n181 VTAIL.n152 1.16414
R1602 VTAIL.n120 VTAIL.n119 1.16414
R1603 VTAIL.n111 VTAIL.n82 1.16414
R1604 VTAIL VTAIL.n69 1.11903
R1605 VTAIL VTAIL.n279 0.532828
R1606 VTAIL.n255 VTAIL.n254 0.388379
R1607 VTAIL.n256 VTAIL.n220 0.388379
R1608 VTAIL.n45 VTAIL.n44 0.388379
R1609 VTAIL.n46 VTAIL.n10 0.388379
R1610 VTAIL.n186 VTAIL.n150 0.388379
R1611 VTAIL.n185 VTAIL.n184 0.388379
R1612 VTAIL.n116 VTAIL.n80 0.388379
R1613 VTAIL.n115 VTAIL.n114 0.388379
R1614 VTAIL.n236 VTAIL.n235 0.155672
R1615 VTAIL.n236 VTAIL.n227 0.155672
R1616 VTAIL.n243 VTAIL.n227 0.155672
R1617 VTAIL.n244 VTAIL.n243 0.155672
R1618 VTAIL.n244 VTAIL.n223 0.155672
R1619 VTAIL.n252 VTAIL.n223 0.155672
R1620 VTAIL.n253 VTAIL.n252 0.155672
R1621 VTAIL.n253 VTAIL.n219 0.155672
R1622 VTAIL.n261 VTAIL.n219 0.155672
R1623 VTAIL.n262 VTAIL.n261 0.155672
R1624 VTAIL.n262 VTAIL.n215 0.155672
R1625 VTAIL.n269 VTAIL.n215 0.155672
R1626 VTAIL.n270 VTAIL.n269 0.155672
R1627 VTAIL.n270 VTAIL.n211 0.155672
R1628 VTAIL.n277 VTAIL.n211 0.155672
R1629 VTAIL.n26 VTAIL.n25 0.155672
R1630 VTAIL.n26 VTAIL.n17 0.155672
R1631 VTAIL.n33 VTAIL.n17 0.155672
R1632 VTAIL.n34 VTAIL.n33 0.155672
R1633 VTAIL.n34 VTAIL.n13 0.155672
R1634 VTAIL.n42 VTAIL.n13 0.155672
R1635 VTAIL.n43 VTAIL.n42 0.155672
R1636 VTAIL.n43 VTAIL.n9 0.155672
R1637 VTAIL.n51 VTAIL.n9 0.155672
R1638 VTAIL.n52 VTAIL.n51 0.155672
R1639 VTAIL.n52 VTAIL.n5 0.155672
R1640 VTAIL.n59 VTAIL.n5 0.155672
R1641 VTAIL.n60 VTAIL.n59 0.155672
R1642 VTAIL.n60 VTAIL.n1 0.155672
R1643 VTAIL.n67 VTAIL.n1 0.155672
R1644 VTAIL.n207 VTAIL.n141 0.155672
R1645 VTAIL.n200 VTAIL.n141 0.155672
R1646 VTAIL.n200 VTAIL.n199 0.155672
R1647 VTAIL.n199 VTAIL.n145 0.155672
R1648 VTAIL.n192 VTAIL.n145 0.155672
R1649 VTAIL.n192 VTAIL.n191 0.155672
R1650 VTAIL.n191 VTAIL.n149 0.155672
R1651 VTAIL.n183 VTAIL.n149 0.155672
R1652 VTAIL.n183 VTAIL.n182 0.155672
R1653 VTAIL.n182 VTAIL.n153 0.155672
R1654 VTAIL.n175 VTAIL.n153 0.155672
R1655 VTAIL.n175 VTAIL.n174 0.155672
R1656 VTAIL.n174 VTAIL.n158 0.155672
R1657 VTAIL.n167 VTAIL.n158 0.155672
R1658 VTAIL.n167 VTAIL.n166 0.155672
R1659 VTAIL.n137 VTAIL.n71 0.155672
R1660 VTAIL.n130 VTAIL.n71 0.155672
R1661 VTAIL.n130 VTAIL.n129 0.155672
R1662 VTAIL.n129 VTAIL.n75 0.155672
R1663 VTAIL.n122 VTAIL.n75 0.155672
R1664 VTAIL.n122 VTAIL.n121 0.155672
R1665 VTAIL.n121 VTAIL.n79 0.155672
R1666 VTAIL.n113 VTAIL.n79 0.155672
R1667 VTAIL.n113 VTAIL.n112 0.155672
R1668 VTAIL.n112 VTAIL.n83 0.155672
R1669 VTAIL.n105 VTAIL.n83 0.155672
R1670 VTAIL.n105 VTAIL.n104 0.155672
R1671 VTAIL.n104 VTAIL.n88 0.155672
R1672 VTAIL.n97 VTAIL.n88 0.155672
R1673 VTAIL.n97 VTAIL.n96 0.155672
R1674 VDD2.n133 VDD2.n69 289.615
R1675 VDD2.n64 VDD2.n0 289.615
R1676 VDD2.n134 VDD2.n133 185
R1677 VDD2.n132 VDD2.n131 185
R1678 VDD2.n73 VDD2.n72 185
R1679 VDD2.n126 VDD2.n125 185
R1680 VDD2.n124 VDD2.n123 185
R1681 VDD2.n77 VDD2.n76 185
R1682 VDD2.n118 VDD2.n117 185
R1683 VDD2.n116 VDD2.n115 185
R1684 VDD2.n114 VDD2.n80 185
R1685 VDD2.n84 VDD2.n81 185
R1686 VDD2.n109 VDD2.n108 185
R1687 VDD2.n107 VDD2.n106 185
R1688 VDD2.n86 VDD2.n85 185
R1689 VDD2.n101 VDD2.n100 185
R1690 VDD2.n99 VDD2.n98 185
R1691 VDD2.n90 VDD2.n89 185
R1692 VDD2.n93 VDD2.n92 185
R1693 VDD2.n23 VDD2.n22 185
R1694 VDD2.n20 VDD2.n19 185
R1695 VDD2.n29 VDD2.n28 185
R1696 VDD2.n31 VDD2.n30 185
R1697 VDD2.n16 VDD2.n15 185
R1698 VDD2.n37 VDD2.n36 185
R1699 VDD2.n40 VDD2.n39 185
R1700 VDD2.n38 VDD2.n12 185
R1701 VDD2.n45 VDD2.n11 185
R1702 VDD2.n47 VDD2.n46 185
R1703 VDD2.n49 VDD2.n48 185
R1704 VDD2.n8 VDD2.n7 185
R1705 VDD2.n55 VDD2.n54 185
R1706 VDD2.n57 VDD2.n56 185
R1707 VDD2.n4 VDD2.n3 185
R1708 VDD2.n63 VDD2.n62 185
R1709 VDD2.n65 VDD2.n64 185
R1710 VDD2.t0 VDD2.n91 149.524
R1711 VDD2.t1 VDD2.n21 149.524
R1712 VDD2.n133 VDD2.n132 104.615
R1713 VDD2.n132 VDD2.n72 104.615
R1714 VDD2.n125 VDD2.n72 104.615
R1715 VDD2.n125 VDD2.n124 104.615
R1716 VDD2.n124 VDD2.n76 104.615
R1717 VDD2.n117 VDD2.n76 104.615
R1718 VDD2.n117 VDD2.n116 104.615
R1719 VDD2.n116 VDD2.n80 104.615
R1720 VDD2.n84 VDD2.n80 104.615
R1721 VDD2.n108 VDD2.n84 104.615
R1722 VDD2.n108 VDD2.n107 104.615
R1723 VDD2.n107 VDD2.n85 104.615
R1724 VDD2.n100 VDD2.n85 104.615
R1725 VDD2.n100 VDD2.n99 104.615
R1726 VDD2.n99 VDD2.n89 104.615
R1727 VDD2.n92 VDD2.n89 104.615
R1728 VDD2.n22 VDD2.n19 104.615
R1729 VDD2.n29 VDD2.n19 104.615
R1730 VDD2.n30 VDD2.n29 104.615
R1731 VDD2.n30 VDD2.n15 104.615
R1732 VDD2.n37 VDD2.n15 104.615
R1733 VDD2.n39 VDD2.n37 104.615
R1734 VDD2.n39 VDD2.n38 104.615
R1735 VDD2.n38 VDD2.n11 104.615
R1736 VDD2.n47 VDD2.n11 104.615
R1737 VDD2.n48 VDD2.n47 104.615
R1738 VDD2.n48 VDD2.n7 104.615
R1739 VDD2.n55 VDD2.n7 104.615
R1740 VDD2.n56 VDD2.n55 104.615
R1741 VDD2.n56 VDD2.n3 104.615
R1742 VDD2.n63 VDD2.n3 104.615
R1743 VDD2.n64 VDD2.n63 104.615
R1744 VDD2.n138 VDD2.n68 87.3039
R1745 VDD2.n92 VDD2.t0 52.3082
R1746 VDD2.n22 VDD2.t1 52.3082
R1747 VDD2.n138 VDD2.n137 47.8944
R1748 VDD2.n115 VDD2.n114 13.1884
R1749 VDD2.n46 VDD2.n45 13.1884
R1750 VDD2.n118 VDD2.n79 12.8005
R1751 VDD2.n113 VDD2.n81 12.8005
R1752 VDD2.n44 VDD2.n12 12.8005
R1753 VDD2.n49 VDD2.n10 12.8005
R1754 VDD2.n119 VDD2.n77 12.0247
R1755 VDD2.n110 VDD2.n109 12.0247
R1756 VDD2.n41 VDD2.n40 12.0247
R1757 VDD2.n50 VDD2.n8 12.0247
R1758 VDD2.n123 VDD2.n122 11.249
R1759 VDD2.n106 VDD2.n83 11.249
R1760 VDD2.n36 VDD2.n14 11.249
R1761 VDD2.n54 VDD2.n53 11.249
R1762 VDD2.n126 VDD2.n75 10.4732
R1763 VDD2.n105 VDD2.n86 10.4732
R1764 VDD2.n35 VDD2.n16 10.4732
R1765 VDD2.n57 VDD2.n6 10.4732
R1766 VDD2.n93 VDD2.n91 10.2747
R1767 VDD2.n23 VDD2.n21 10.2747
R1768 VDD2.n127 VDD2.n73 9.69747
R1769 VDD2.n102 VDD2.n101 9.69747
R1770 VDD2.n32 VDD2.n31 9.69747
R1771 VDD2.n58 VDD2.n4 9.69747
R1772 VDD2.n137 VDD2.n136 9.45567
R1773 VDD2.n68 VDD2.n67 9.45567
R1774 VDD2.n95 VDD2.n94 9.3005
R1775 VDD2.n97 VDD2.n96 9.3005
R1776 VDD2.n88 VDD2.n87 9.3005
R1777 VDD2.n103 VDD2.n102 9.3005
R1778 VDD2.n105 VDD2.n104 9.3005
R1779 VDD2.n83 VDD2.n82 9.3005
R1780 VDD2.n111 VDD2.n110 9.3005
R1781 VDD2.n113 VDD2.n112 9.3005
R1782 VDD2.n136 VDD2.n135 9.3005
R1783 VDD2.n71 VDD2.n70 9.3005
R1784 VDD2.n130 VDD2.n129 9.3005
R1785 VDD2.n128 VDD2.n127 9.3005
R1786 VDD2.n75 VDD2.n74 9.3005
R1787 VDD2.n122 VDD2.n121 9.3005
R1788 VDD2.n120 VDD2.n119 9.3005
R1789 VDD2.n79 VDD2.n78 9.3005
R1790 VDD2.n2 VDD2.n1 9.3005
R1791 VDD2.n61 VDD2.n60 9.3005
R1792 VDD2.n59 VDD2.n58 9.3005
R1793 VDD2.n6 VDD2.n5 9.3005
R1794 VDD2.n53 VDD2.n52 9.3005
R1795 VDD2.n51 VDD2.n50 9.3005
R1796 VDD2.n10 VDD2.n9 9.3005
R1797 VDD2.n25 VDD2.n24 9.3005
R1798 VDD2.n27 VDD2.n26 9.3005
R1799 VDD2.n18 VDD2.n17 9.3005
R1800 VDD2.n33 VDD2.n32 9.3005
R1801 VDD2.n35 VDD2.n34 9.3005
R1802 VDD2.n14 VDD2.n13 9.3005
R1803 VDD2.n42 VDD2.n41 9.3005
R1804 VDD2.n44 VDD2.n43 9.3005
R1805 VDD2.n67 VDD2.n66 9.3005
R1806 VDD2.n131 VDD2.n130 8.92171
R1807 VDD2.n98 VDD2.n88 8.92171
R1808 VDD2.n28 VDD2.n18 8.92171
R1809 VDD2.n62 VDD2.n61 8.92171
R1810 VDD2.n134 VDD2.n71 8.14595
R1811 VDD2.n97 VDD2.n90 8.14595
R1812 VDD2.n27 VDD2.n20 8.14595
R1813 VDD2.n65 VDD2.n2 8.14595
R1814 VDD2.n135 VDD2.n69 7.3702
R1815 VDD2.n94 VDD2.n93 7.3702
R1816 VDD2.n24 VDD2.n23 7.3702
R1817 VDD2.n66 VDD2.n0 7.3702
R1818 VDD2.n137 VDD2.n69 6.59444
R1819 VDD2.n68 VDD2.n0 6.59444
R1820 VDD2.n135 VDD2.n134 5.81868
R1821 VDD2.n94 VDD2.n90 5.81868
R1822 VDD2.n24 VDD2.n20 5.81868
R1823 VDD2.n66 VDD2.n65 5.81868
R1824 VDD2.n131 VDD2.n71 5.04292
R1825 VDD2.n98 VDD2.n97 5.04292
R1826 VDD2.n28 VDD2.n27 5.04292
R1827 VDD2.n62 VDD2.n2 5.04292
R1828 VDD2.n130 VDD2.n73 4.26717
R1829 VDD2.n101 VDD2.n88 4.26717
R1830 VDD2.n31 VDD2.n18 4.26717
R1831 VDD2.n61 VDD2.n4 4.26717
R1832 VDD2.n127 VDD2.n126 3.49141
R1833 VDD2.n102 VDD2.n86 3.49141
R1834 VDD2.n32 VDD2.n16 3.49141
R1835 VDD2.n58 VDD2.n57 3.49141
R1836 VDD2.n95 VDD2.n91 2.84303
R1837 VDD2.n25 VDD2.n21 2.84303
R1838 VDD2.n123 VDD2.n75 2.71565
R1839 VDD2.n106 VDD2.n105 2.71565
R1840 VDD2.n36 VDD2.n35 2.71565
R1841 VDD2.n54 VDD2.n6 2.71565
R1842 VDD2.n122 VDD2.n77 1.93989
R1843 VDD2.n109 VDD2.n83 1.93989
R1844 VDD2.n40 VDD2.n14 1.93989
R1845 VDD2.n53 VDD2.n8 1.93989
R1846 VDD2.n119 VDD2.n118 1.16414
R1847 VDD2.n110 VDD2.n81 1.16414
R1848 VDD2.n41 VDD2.n12 1.16414
R1849 VDD2.n50 VDD2.n49 1.16414
R1850 VDD2 VDD2.n138 0.649207
R1851 VDD2.n115 VDD2.n79 0.388379
R1852 VDD2.n114 VDD2.n113 0.388379
R1853 VDD2.n45 VDD2.n44 0.388379
R1854 VDD2.n46 VDD2.n10 0.388379
R1855 VDD2.n136 VDD2.n70 0.155672
R1856 VDD2.n129 VDD2.n70 0.155672
R1857 VDD2.n129 VDD2.n128 0.155672
R1858 VDD2.n128 VDD2.n74 0.155672
R1859 VDD2.n121 VDD2.n74 0.155672
R1860 VDD2.n121 VDD2.n120 0.155672
R1861 VDD2.n120 VDD2.n78 0.155672
R1862 VDD2.n112 VDD2.n78 0.155672
R1863 VDD2.n112 VDD2.n111 0.155672
R1864 VDD2.n111 VDD2.n82 0.155672
R1865 VDD2.n104 VDD2.n82 0.155672
R1866 VDD2.n104 VDD2.n103 0.155672
R1867 VDD2.n103 VDD2.n87 0.155672
R1868 VDD2.n96 VDD2.n87 0.155672
R1869 VDD2.n96 VDD2.n95 0.155672
R1870 VDD2.n26 VDD2.n25 0.155672
R1871 VDD2.n26 VDD2.n17 0.155672
R1872 VDD2.n33 VDD2.n17 0.155672
R1873 VDD2.n34 VDD2.n33 0.155672
R1874 VDD2.n34 VDD2.n13 0.155672
R1875 VDD2.n42 VDD2.n13 0.155672
R1876 VDD2.n43 VDD2.n42 0.155672
R1877 VDD2.n43 VDD2.n9 0.155672
R1878 VDD2.n51 VDD2.n9 0.155672
R1879 VDD2.n52 VDD2.n51 0.155672
R1880 VDD2.n52 VDD2.n5 0.155672
R1881 VDD2.n59 VDD2.n5 0.155672
R1882 VDD2.n60 VDD2.n59 0.155672
R1883 VDD2.n60 VDD2.n1 0.155672
R1884 VDD2.n67 VDD2.n1 0.155672
R1885 VP.n0 VP.t1 221.821
R1886 VP.n0 VP.t0 177.071
R1887 VP VP.n0 0.336784
R1888 VDD1.n64 VDD1.n0 289.615
R1889 VDD1.n133 VDD1.n69 289.615
R1890 VDD1.n65 VDD1.n64 185
R1891 VDD1.n63 VDD1.n62 185
R1892 VDD1.n4 VDD1.n3 185
R1893 VDD1.n57 VDD1.n56 185
R1894 VDD1.n55 VDD1.n54 185
R1895 VDD1.n8 VDD1.n7 185
R1896 VDD1.n49 VDD1.n48 185
R1897 VDD1.n47 VDD1.n46 185
R1898 VDD1.n45 VDD1.n11 185
R1899 VDD1.n15 VDD1.n12 185
R1900 VDD1.n40 VDD1.n39 185
R1901 VDD1.n38 VDD1.n37 185
R1902 VDD1.n17 VDD1.n16 185
R1903 VDD1.n32 VDD1.n31 185
R1904 VDD1.n30 VDD1.n29 185
R1905 VDD1.n21 VDD1.n20 185
R1906 VDD1.n24 VDD1.n23 185
R1907 VDD1.n92 VDD1.n91 185
R1908 VDD1.n89 VDD1.n88 185
R1909 VDD1.n98 VDD1.n97 185
R1910 VDD1.n100 VDD1.n99 185
R1911 VDD1.n85 VDD1.n84 185
R1912 VDD1.n106 VDD1.n105 185
R1913 VDD1.n109 VDD1.n108 185
R1914 VDD1.n107 VDD1.n81 185
R1915 VDD1.n114 VDD1.n80 185
R1916 VDD1.n116 VDD1.n115 185
R1917 VDD1.n118 VDD1.n117 185
R1918 VDD1.n77 VDD1.n76 185
R1919 VDD1.n124 VDD1.n123 185
R1920 VDD1.n126 VDD1.n125 185
R1921 VDD1.n73 VDD1.n72 185
R1922 VDD1.n132 VDD1.n131 185
R1923 VDD1.n134 VDD1.n133 185
R1924 VDD1.t0 VDD1.n22 149.524
R1925 VDD1.t1 VDD1.n90 149.524
R1926 VDD1.n64 VDD1.n63 104.615
R1927 VDD1.n63 VDD1.n3 104.615
R1928 VDD1.n56 VDD1.n3 104.615
R1929 VDD1.n56 VDD1.n55 104.615
R1930 VDD1.n55 VDD1.n7 104.615
R1931 VDD1.n48 VDD1.n7 104.615
R1932 VDD1.n48 VDD1.n47 104.615
R1933 VDD1.n47 VDD1.n11 104.615
R1934 VDD1.n15 VDD1.n11 104.615
R1935 VDD1.n39 VDD1.n15 104.615
R1936 VDD1.n39 VDD1.n38 104.615
R1937 VDD1.n38 VDD1.n16 104.615
R1938 VDD1.n31 VDD1.n16 104.615
R1939 VDD1.n31 VDD1.n30 104.615
R1940 VDD1.n30 VDD1.n20 104.615
R1941 VDD1.n23 VDD1.n20 104.615
R1942 VDD1.n91 VDD1.n88 104.615
R1943 VDD1.n98 VDD1.n88 104.615
R1944 VDD1.n99 VDD1.n98 104.615
R1945 VDD1.n99 VDD1.n84 104.615
R1946 VDD1.n106 VDD1.n84 104.615
R1947 VDD1.n108 VDD1.n106 104.615
R1948 VDD1.n108 VDD1.n107 104.615
R1949 VDD1.n107 VDD1.n80 104.615
R1950 VDD1.n116 VDD1.n80 104.615
R1951 VDD1.n117 VDD1.n116 104.615
R1952 VDD1.n117 VDD1.n76 104.615
R1953 VDD1.n124 VDD1.n76 104.615
R1954 VDD1.n125 VDD1.n124 104.615
R1955 VDD1.n125 VDD1.n72 104.615
R1956 VDD1.n132 VDD1.n72 104.615
R1957 VDD1.n133 VDD1.n132 104.615
R1958 VDD1 VDD1.n137 88.4192
R1959 VDD1.n23 VDD1.t0 52.3082
R1960 VDD1.n91 VDD1.t1 52.3082
R1961 VDD1 VDD1.n68 48.5431
R1962 VDD1.n46 VDD1.n45 13.1884
R1963 VDD1.n115 VDD1.n114 13.1884
R1964 VDD1.n49 VDD1.n10 12.8005
R1965 VDD1.n44 VDD1.n12 12.8005
R1966 VDD1.n113 VDD1.n81 12.8005
R1967 VDD1.n118 VDD1.n79 12.8005
R1968 VDD1.n50 VDD1.n8 12.0247
R1969 VDD1.n41 VDD1.n40 12.0247
R1970 VDD1.n110 VDD1.n109 12.0247
R1971 VDD1.n119 VDD1.n77 12.0247
R1972 VDD1.n54 VDD1.n53 11.249
R1973 VDD1.n37 VDD1.n14 11.249
R1974 VDD1.n105 VDD1.n83 11.249
R1975 VDD1.n123 VDD1.n122 11.249
R1976 VDD1.n57 VDD1.n6 10.4732
R1977 VDD1.n36 VDD1.n17 10.4732
R1978 VDD1.n104 VDD1.n85 10.4732
R1979 VDD1.n126 VDD1.n75 10.4732
R1980 VDD1.n24 VDD1.n22 10.2747
R1981 VDD1.n92 VDD1.n90 10.2747
R1982 VDD1.n58 VDD1.n4 9.69747
R1983 VDD1.n33 VDD1.n32 9.69747
R1984 VDD1.n101 VDD1.n100 9.69747
R1985 VDD1.n127 VDD1.n73 9.69747
R1986 VDD1.n68 VDD1.n67 9.45567
R1987 VDD1.n137 VDD1.n136 9.45567
R1988 VDD1.n26 VDD1.n25 9.3005
R1989 VDD1.n28 VDD1.n27 9.3005
R1990 VDD1.n19 VDD1.n18 9.3005
R1991 VDD1.n34 VDD1.n33 9.3005
R1992 VDD1.n36 VDD1.n35 9.3005
R1993 VDD1.n14 VDD1.n13 9.3005
R1994 VDD1.n42 VDD1.n41 9.3005
R1995 VDD1.n44 VDD1.n43 9.3005
R1996 VDD1.n67 VDD1.n66 9.3005
R1997 VDD1.n2 VDD1.n1 9.3005
R1998 VDD1.n61 VDD1.n60 9.3005
R1999 VDD1.n59 VDD1.n58 9.3005
R2000 VDD1.n6 VDD1.n5 9.3005
R2001 VDD1.n53 VDD1.n52 9.3005
R2002 VDD1.n51 VDD1.n50 9.3005
R2003 VDD1.n10 VDD1.n9 9.3005
R2004 VDD1.n71 VDD1.n70 9.3005
R2005 VDD1.n130 VDD1.n129 9.3005
R2006 VDD1.n128 VDD1.n127 9.3005
R2007 VDD1.n75 VDD1.n74 9.3005
R2008 VDD1.n122 VDD1.n121 9.3005
R2009 VDD1.n120 VDD1.n119 9.3005
R2010 VDD1.n79 VDD1.n78 9.3005
R2011 VDD1.n94 VDD1.n93 9.3005
R2012 VDD1.n96 VDD1.n95 9.3005
R2013 VDD1.n87 VDD1.n86 9.3005
R2014 VDD1.n102 VDD1.n101 9.3005
R2015 VDD1.n104 VDD1.n103 9.3005
R2016 VDD1.n83 VDD1.n82 9.3005
R2017 VDD1.n111 VDD1.n110 9.3005
R2018 VDD1.n113 VDD1.n112 9.3005
R2019 VDD1.n136 VDD1.n135 9.3005
R2020 VDD1.n62 VDD1.n61 8.92171
R2021 VDD1.n29 VDD1.n19 8.92171
R2022 VDD1.n97 VDD1.n87 8.92171
R2023 VDD1.n131 VDD1.n130 8.92171
R2024 VDD1.n65 VDD1.n2 8.14595
R2025 VDD1.n28 VDD1.n21 8.14595
R2026 VDD1.n96 VDD1.n89 8.14595
R2027 VDD1.n134 VDD1.n71 8.14595
R2028 VDD1.n66 VDD1.n0 7.3702
R2029 VDD1.n25 VDD1.n24 7.3702
R2030 VDD1.n93 VDD1.n92 7.3702
R2031 VDD1.n135 VDD1.n69 7.3702
R2032 VDD1.n68 VDD1.n0 6.59444
R2033 VDD1.n137 VDD1.n69 6.59444
R2034 VDD1.n66 VDD1.n65 5.81868
R2035 VDD1.n25 VDD1.n21 5.81868
R2036 VDD1.n93 VDD1.n89 5.81868
R2037 VDD1.n135 VDD1.n134 5.81868
R2038 VDD1.n62 VDD1.n2 5.04292
R2039 VDD1.n29 VDD1.n28 5.04292
R2040 VDD1.n97 VDD1.n96 5.04292
R2041 VDD1.n131 VDD1.n71 5.04292
R2042 VDD1.n61 VDD1.n4 4.26717
R2043 VDD1.n32 VDD1.n19 4.26717
R2044 VDD1.n100 VDD1.n87 4.26717
R2045 VDD1.n130 VDD1.n73 4.26717
R2046 VDD1.n58 VDD1.n57 3.49141
R2047 VDD1.n33 VDD1.n17 3.49141
R2048 VDD1.n101 VDD1.n85 3.49141
R2049 VDD1.n127 VDD1.n126 3.49141
R2050 VDD1.n26 VDD1.n22 2.84303
R2051 VDD1.n94 VDD1.n90 2.84303
R2052 VDD1.n54 VDD1.n6 2.71565
R2053 VDD1.n37 VDD1.n36 2.71565
R2054 VDD1.n105 VDD1.n104 2.71565
R2055 VDD1.n123 VDD1.n75 2.71565
R2056 VDD1.n53 VDD1.n8 1.93989
R2057 VDD1.n40 VDD1.n14 1.93989
R2058 VDD1.n109 VDD1.n83 1.93989
R2059 VDD1.n122 VDD1.n77 1.93989
R2060 VDD1.n50 VDD1.n49 1.16414
R2061 VDD1.n41 VDD1.n12 1.16414
R2062 VDD1.n110 VDD1.n81 1.16414
R2063 VDD1.n119 VDD1.n118 1.16414
R2064 VDD1.n46 VDD1.n10 0.388379
R2065 VDD1.n45 VDD1.n44 0.388379
R2066 VDD1.n114 VDD1.n113 0.388379
R2067 VDD1.n115 VDD1.n79 0.388379
R2068 VDD1.n67 VDD1.n1 0.155672
R2069 VDD1.n60 VDD1.n1 0.155672
R2070 VDD1.n60 VDD1.n59 0.155672
R2071 VDD1.n59 VDD1.n5 0.155672
R2072 VDD1.n52 VDD1.n5 0.155672
R2073 VDD1.n52 VDD1.n51 0.155672
R2074 VDD1.n51 VDD1.n9 0.155672
R2075 VDD1.n43 VDD1.n9 0.155672
R2076 VDD1.n43 VDD1.n42 0.155672
R2077 VDD1.n42 VDD1.n13 0.155672
R2078 VDD1.n35 VDD1.n13 0.155672
R2079 VDD1.n35 VDD1.n34 0.155672
R2080 VDD1.n34 VDD1.n18 0.155672
R2081 VDD1.n27 VDD1.n18 0.155672
R2082 VDD1.n27 VDD1.n26 0.155672
R2083 VDD1.n95 VDD1.n94 0.155672
R2084 VDD1.n95 VDD1.n86 0.155672
R2085 VDD1.n102 VDD1.n86 0.155672
R2086 VDD1.n103 VDD1.n102 0.155672
R2087 VDD1.n103 VDD1.n82 0.155672
R2088 VDD1.n111 VDD1.n82 0.155672
R2089 VDD1.n112 VDD1.n111 0.155672
R2090 VDD1.n112 VDD1.n78 0.155672
R2091 VDD1.n120 VDD1.n78 0.155672
R2092 VDD1.n121 VDD1.n120 0.155672
R2093 VDD1.n121 VDD1.n74 0.155672
R2094 VDD1.n128 VDD1.n74 0.155672
R2095 VDD1.n129 VDD1.n128 0.155672
R2096 VDD1.n129 VDD1.n70 0.155672
R2097 VDD1.n136 VDD1.n70 0.155672
C0 VDD2 VN 2.91129f
C1 VP VDD1 3.08563f
C2 VTAIL VDD1 5.25454f
C3 VP VTAIL 2.53864f
C4 VDD2 VDD1 0.651971f
C5 VP VDD2 0.325161f
C6 VDD2 VTAIL 5.30347f
C7 VDD1 VN 0.148035f
C8 VP VN 5.51238f
C9 VTAIL VN 2.52432f
C10 VDD2 B 4.505587f
C11 VDD1 B 7.26555f
C12 VTAIL B 7.605919f
C13 VN B 10.66937f
C14 VP B 6.214713f
C15 VDD1.n0 B 0.028602f
C16 VDD1.n1 B 0.020447f
C17 VDD1.n2 B 0.010987f
C18 VDD1.n3 B 0.02597f
C19 VDD1.n4 B 0.011633f
C20 VDD1.n5 B 0.020447f
C21 VDD1.n6 B 0.010987f
C22 VDD1.n7 B 0.02597f
C23 VDD1.n8 B 0.011633f
C24 VDD1.n9 B 0.020447f
C25 VDD1.n10 B 0.010987f
C26 VDD1.n11 B 0.02597f
C27 VDD1.n12 B 0.011633f
C28 VDD1.n13 B 0.020447f
C29 VDD1.n14 B 0.010987f
C30 VDD1.n15 B 0.02597f
C31 VDD1.n16 B 0.02597f
C32 VDD1.n17 B 0.011633f
C33 VDD1.n18 B 0.020447f
C34 VDD1.n19 B 0.010987f
C35 VDD1.n20 B 0.02597f
C36 VDD1.n21 B 0.011633f
C37 VDD1.n22 B 0.153619f
C38 VDD1.t0 B 0.043948f
C39 VDD1.n23 B 0.019477f
C40 VDD1.n24 B 0.018358f
C41 VDD1.n25 B 0.010987f
C42 VDD1.n26 B 1.10334f
C43 VDD1.n27 B 0.020447f
C44 VDD1.n28 B 0.010987f
C45 VDD1.n29 B 0.011633f
C46 VDD1.n30 B 0.02597f
C47 VDD1.n31 B 0.02597f
C48 VDD1.n32 B 0.011633f
C49 VDD1.n33 B 0.010987f
C50 VDD1.n34 B 0.020447f
C51 VDD1.n35 B 0.020447f
C52 VDD1.n36 B 0.010987f
C53 VDD1.n37 B 0.011633f
C54 VDD1.n38 B 0.02597f
C55 VDD1.n39 B 0.02597f
C56 VDD1.n40 B 0.011633f
C57 VDD1.n41 B 0.010987f
C58 VDD1.n42 B 0.020447f
C59 VDD1.n43 B 0.020447f
C60 VDD1.n44 B 0.010987f
C61 VDD1.n45 B 0.01131f
C62 VDD1.n46 B 0.01131f
C63 VDD1.n47 B 0.02597f
C64 VDD1.n48 B 0.02597f
C65 VDD1.n49 B 0.011633f
C66 VDD1.n50 B 0.010987f
C67 VDD1.n51 B 0.020447f
C68 VDD1.n52 B 0.020447f
C69 VDD1.n53 B 0.010987f
C70 VDD1.n54 B 0.011633f
C71 VDD1.n55 B 0.02597f
C72 VDD1.n56 B 0.02597f
C73 VDD1.n57 B 0.011633f
C74 VDD1.n58 B 0.010987f
C75 VDD1.n59 B 0.020447f
C76 VDD1.n60 B 0.020447f
C77 VDD1.n61 B 0.010987f
C78 VDD1.n62 B 0.011633f
C79 VDD1.n63 B 0.02597f
C80 VDD1.n64 B 0.055976f
C81 VDD1.n65 B 0.011633f
C82 VDD1.n66 B 0.010987f
C83 VDD1.n67 B 0.045865f
C84 VDD1.n68 B 0.046468f
C85 VDD1.n69 B 0.028602f
C86 VDD1.n70 B 0.020447f
C87 VDD1.n71 B 0.010987f
C88 VDD1.n72 B 0.02597f
C89 VDD1.n73 B 0.011633f
C90 VDD1.n74 B 0.020447f
C91 VDD1.n75 B 0.010987f
C92 VDD1.n76 B 0.02597f
C93 VDD1.n77 B 0.011633f
C94 VDD1.n78 B 0.020447f
C95 VDD1.n79 B 0.010987f
C96 VDD1.n80 B 0.02597f
C97 VDD1.n81 B 0.011633f
C98 VDD1.n82 B 0.020447f
C99 VDD1.n83 B 0.010987f
C100 VDD1.n84 B 0.02597f
C101 VDD1.n85 B 0.011633f
C102 VDD1.n86 B 0.020447f
C103 VDD1.n87 B 0.010987f
C104 VDD1.n88 B 0.02597f
C105 VDD1.n89 B 0.011633f
C106 VDD1.n90 B 0.153619f
C107 VDD1.t1 B 0.043948f
C108 VDD1.n91 B 0.019477f
C109 VDD1.n92 B 0.018358f
C110 VDD1.n93 B 0.010987f
C111 VDD1.n94 B 1.10334f
C112 VDD1.n95 B 0.020447f
C113 VDD1.n96 B 0.010987f
C114 VDD1.n97 B 0.011633f
C115 VDD1.n98 B 0.02597f
C116 VDD1.n99 B 0.02597f
C117 VDD1.n100 B 0.011633f
C118 VDD1.n101 B 0.010987f
C119 VDD1.n102 B 0.020447f
C120 VDD1.n103 B 0.020447f
C121 VDD1.n104 B 0.010987f
C122 VDD1.n105 B 0.011633f
C123 VDD1.n106 B 0.02597f
C124 VDD1.n107 B 0.02597f
C125 VDD1.n108 B 0.02597f
C126 VDD1.n109 B 0.011633f
C127 VDD1.n110 B 0.010987f
C128 VDD1.n111 B 0.020447f
C129 VDD1.n112 B 0.020447f
C130 VDD1.n113 B 0.010987f
C131 VDD1.n114 B 0.01131f
C132 VDD1.n115 B 0.01131f
C133 VDD1.n116 B 0.02597f
C134 VDD1.n117 B 0.02597f
C135 VDD1.n118 B 0.011633f
C136 VDD1.n119 B 0.010987f
C137 VDD1.n120 B 0.020447f
C138 VDD1.n121 B 0.020447f
C139 VDD1.n122 B 0.010987f
C140 VDD1.n123 B 0.011633f
C141 VDD1.n124 B 0.02597f
C142 VDD1.n125 B 0.02597f
C143 VDD1.n126 B 0.011633f
C144 VDD1.n127 B 0.010987f
C145 VDD1.n128 B 0.020447f
C146 VDD1.n129 B 0.020447f
C147 VDD1.n130 B 0.010987f
C148 VDD1.n131 B 0.011633f
C149 VDD1.n132 B 0.02597f
C150 VDD1.n133 B 0.055976f
C151 VDD1.n134 B 0.011633f
C152 VDD1.n135 B 0.010987f
C153 VDD1.n136 B 0.045865f
C154 VDD1.n137 B 0.659351f
C155 VP.t1 B 3.56547f
C156 VP.t0 B 3.06721f
C157 VP.n0 B 4.39496f
C158 VDD2.n0 B 0.028174f
C159 VDD2.n1 B 0.020141f
C160 VDD2.n2 B 0.010823f
C161 VDD2.n3 B 0.025581f
C162 VDD2.n4 B 0.01146f
C163 VDD2.n5 B 0.020141f
C164 VDD2.n6 B 0.010823f
C165 VDD2.n7 B 0.025581f
C166 VDD2.n8 B 0.01146f
C167 VDD2.n9 B 0.020141f
C168 VDD2.n10 B 0.010823f
C169 VDD2.n11 B 0.025581f
C170 VDD2.n12 B 0.01146f
C171 VDD2.n13 B 0.020141f
C172 VDD2.n14 B 0.010823f
C173 VDD2.n15 B 0.025581f
C174 VDD2.n16 B 0.01146f
C175 VDD2.n17 B 0.020141f
C176 VDD2.n18 B 0.010823f
C177 VDD2.n19 B 0.025581f
C178 VDD2.n20 B 0.01146f
C179 VDD2.n21 B 0.151322f
C180 VDD2.t1 B 0.043291f
C181 VDD2.n22 B 0.019186f
C182 VDD2.n23 B 0.018084f
C183 VDD2.n24 B 0.010823f
C184 VDD2.n25 B 1.08684f
C185 VDD2.n26 B 0.020141f
C186 VDD2.n27 B 0.010823f
C187 VDD2.n28 B 0.01146f
C188 VDD2.n29 B 0.025581f
C189 VDD2.n30 B 0.025581f
C190 VDD2.n31 B 0.01146f
C191 VDD2.n32 B 0.010823f
C192 VDD2.n33 B 0.020141f
C193 VDD2.n34 B 0.020141f
C194 VDD2.n35 B 0.010823f
C195 VDD2.n36 B 0.01146f
C196 VDD2.n37 B 0.025581f
C197 VDD2.n38 B 0.025581f
C198 VDD2.n39 B 0.025581f
C199 VDD2.n40 B 0.01146f
C200 VDD2.n41 B 0.010823f
C201 VDD2.n42 B 0.020141f
C202 VDD2.n43 B 0.020141f
C203 VDD2.n44 B 0.010823f
C204 VDD2.n45 B 0.011141f
C205 VDD2.n46 B 0.011141f
C206 VDD2.n47 B 0.025581f
C207 VDD2.n48 B 0.025581f
C208 VDD2.n49 B 0.01146f
C209 VDD2.n50 B 0.010823f
C210 VDD2.n51 B 0.020141f
C211 VDD2.n52 B 0.020141f
C212 VDD2.n53 B 0.010823f
C213 VDD2.n54 B 0.01146f
C214 VDD2.n55 B 0.025581f
C215 VDD2.n56 B 0.025581f
C216 VDD2.n57 B 0.01146f
C217 VDD2.n58 B 0.010823f
C218 VDD2.n59 B 0.020141f
C219 VDD2.n60 B 0.020141f
C220 VDD2.n61 B 0.010823f
C221 VDD2.n62 B 0.01146f
C222 VDD2.n63 B 0.025581f
C223 VDD2.n64 B 0.055139f
C224 VDD2.n65 B 0.01146f
C225 VDD2.n66 B 0.010823f
C226 VDD2.n67 B 0.045179f
C227 VDD2.n68 B 0.610448f
C228 VDD2.n69 B 0.028174f
C229 VDD2.n70 B 0.020141f
C230 VDD2.n71 B 0.010823f
C231 VDD2.n72 B 0.025581f
C232 VDD2.n73 B 0.01146f
C233 VDD2.n74 B 0.020141f
C234 VDD2.n75 B 0.010823f
C235 VDD2.n76 B 0.025581f
C236 VDD2.n77 B 0.01146f
C237 VDD2.n78 B 0.020141f
C238 VDD2.n79 B 0.010823f
C239 VDD2.n80 B 0.025581f
C240 VDD2.n81 B 0.01146f
C241 VDD2.n82 B 0.020141f
C242 VDD2.n83 B 0.010823f
C243 VDD2.n84 B 0.025581f
C244 VDD2.n85 B 0.025581f
C245 VDD2.n86 B 0.01146f
C246 VDD2.n87 B 0.020141f
C247 VDD2.n88 B 0.010823f
C248 VDD2.n89 B 0.025581f
C249 VDD2.n90 B 0.01146f
C250 VDD2.n91 B 0.151322f
C251 VDD2.t0 B 0.043291f
C252 VDD2.n92 B 0.019186f
C253 VDD2.n93 B 0.018084f
C254 VDD2.n94 B 0.010823f
C255 VDD2.n95 B 1.08684f
C256 VDD2.n96 B 0.020141f
C257 VDD2.n97 B 0.010823f
C258 VDD2.n98 B 0.01146f
C259 VDD2.n99 B 0.025581f
C260 VDD2.n100 B 0.025581f
C261 VDD2.n101 B 0.01146f
C262 VDD2.n102 B 0.010823f
C263 VDD2.n103 B 0.020141f
C264 VDD2.n104 B 0.020141f
C265 VDD2.n105 B 0.010823f
C266 VDD2.n106 B 0.01146f
C267 VDD2.n107 B 0.025581f
C268 VDD2.n108 B 0.025581f
C269 VDD2.n109 B 0.01146f
C270 VDD2.n110 B 0.010823f
C271 VDD2.n111 B 0.020141f
C272 VDD2.n112 B 0.020141f
C273 VDD2.n113 B 0.010823f
C274 VDD2.n114 B 0.011141f
C275 VDD2.n115 B 0.011141f
C276 VDD2.n116 B 0.025581f
C277 VDD2.n117 B 0.025581f
C278 VDD2.n118 B 0.01146f
C279 VDD2.n119 B 0.010823f
C280 VDD2.n120 B 0.020141f
C281 VDD2.n121 B 0.020141f
C282 VDD2.n122 B 0.010823f
C283 VDD2.n123 B 0.01146f
C284 VDD2.n124 B 0.025581f
C285 VDD2.n125 B 0.025581f
C286 VDD2.n126 B 0.01146f
C287 VDD2.n127 B 0.010823f
C288 VDD2.n128 B 0.020141f
C289 VDD2.n129 B 0.020141f
C290 VDD2.n130 B 0.010823f
C291 VDD2.n131 B 0.01146f
C292 VDD2.n132 B 0.025581f
C293 VDD2.n133 B 0.055139f
C294 VDD2.n134 B 0.01146f
C295 VDD2.n135 B 0.010823f
C296 VDD2.n136 B 0.045179f
C297 VDD2.n137 B 0.044703f
C298 VDD2.n138 B 2.48797f
C299 VTAIL.n0 B 0.028598f
C300 VTAIL.n1 B 0.020444f
C301 VTAIL.n2 B 0.010986f
C302 VTAIL.n3 B 0.025966f
C303 VTAIL.n4 B 0.011632f
C304 VTAIL.n5 B 0.020444f
C305 VTAIL.n6 B 0.010986f
C306 VTAIL.n7 B 0.025966f
C307 VTAIL.n8 B 0.011632f
C308 VTAIL.n9 B 0.020444f
C309 VTAIL.n10 B 0.010986f
C310 VTAIL.n11 B 0.025966f
C311 VTAIL.n12 B 0.011632f
C312 VTAIL.n13 B 0.020444f
C313 VTAIL.n14 B 0.010986f
C314 VTAIL.n15 B 0.025966f
C315 VTAIL.n16 B 0.011632f
C316 VTAIL.n17 B 0.020444f
C317 VTAIL.n18 B 0.010986f
C318 VTAIL.n19 B 0.025966f
C319 VTAIL.n20 B 0.011632f
C320 VTAIL.n21 B 0.153597f
C321 VTAIL.t0 B 0.043942f
C322 VTAIL.n22 B 0.019474f
C323 VTAIL.n23 B 0.018356f
C324 VTAIL.n24 B 0.010986f
C325 VTAIL.n25 B 1.10319f
C326 VTAIL.n26 B 0.020444f
C327 VTAIL.n27 B 0.010986f
C328 VTAIL.n28 B 0.011632f
C329 VTAIL.n29 B 0.025966f
C330 VTAIL.n30 B 0.025966f
C331 VTAIL.n31 B 0.011632f
C332 VTAIL.n32 B 0.010986f
C333 VTAIL.n33 B 0.020444f
C334 VTAIL.n34 B 0.020444f
C335 VTAIL.n35 B 0.010986f
C336 VTAIL.n36 B 0.011632f
C337 VTAIL.n37 B 0.025966f
C338 VTAIL.n38 B 0.025966f
C339 VTAIL.n39 B 0.025966f
C340 VTAIL.n40 B 0.011632f
C341 VTAIL.n41 B 0.010986f
C342 VTAIL.n42 B 0.020444f
C343 VTAIL.n43 B 0.020444f
C344 VTAIL.n44 B 0.010986f
C345 VTAIL.n45 B 0.011309f
C346 VTAIL.n46 B 0.011309f
C347 VTAIL.n47 B 0.025966f
C348 VTAIL.n48 B 0.025966f
C349 VTAIL.n49 B 0.011632f
C350 VTAIL.n50 B 0.010986f
C351 VTAIL.n51 B 0.020444f
C352 VTAIL.n52 B 0.020444f
C353 VTAIL.n53 B 0.010986f
C354 VTAIL.n54 B 0.011632f
C355 VTAIL.n55 B 0.025966f
C356 VTAIL.n56 B 0.025966f
C357 VTAIL.n57 B 0.011632f
C358 VTAIL.n58 B 0.010986f
C359 VTAIL.n59 B 0.020444f
C360 VTAIL.n60 B 0.020444f
C361 VTAIL.n61 B 0.010986f
C362 VTAIL.n62 B 0.011632f
C363 VTAIL.n63 B 0.025966f
C364 VTAIL.n64 B 0.055968f
C365 VTAIL.n65 B 0.011632f
C366 VTAIL.n66 B 0.010986f
C367 VTAIL.n67 B 0.045858f
C368 VTAIL.n68 B 0.031248f
C369 VTAIL.n69 B 1.40558f
C370 VTAIL.n70 B 0.028598f
C371 VTAIL.n71 B 0.020444f
C372 VTAIL.n72 B 0.010986f
C373 VTAIL.n73 B 0.025966f
C374 VTAIL.n74 B 0.011632f
C375 VTAIL.n75 B 0.020444f
C376 VTAIL.n76 B 0.010986f
C377 VTAIL.n77 B 0.025966f
C378 VTAIL.n78 B 0.011632f
C379 VTAIL.n79 B 0.020444f
C380 VTAIL.n80 B 0.010986f
C381 VTAIL.n81 B 0.025966f
C382 VTAIL.n82 B 0.011632f
C383 VTAIL.n83 B 0.020444f
C384 VTAIL.n84 B 0.010986f
C385 VTAIL.n85 B 0.025966f
C386 VTAIL.n86 B 0.025966f
C387 VTAIL.n87 B 0.011632f
C388 VTAIL.n88 B 0.020444f
C389 VTAIL.n89 B 0.010986f
C390 VTAIL.n90 B 0.025966f
C391 VTAIL.n91 B 0.011632f
C392 VTAIL.n92 B 0.153597f
C393 VTAIL.t2 B 0.043942f
C394 VTAIL.n93 B 0.019474f
C395 VTAIL.n94 B 0.018356f
C396 VTAIL.n95 B 0.010986f
C397 VTAIL.n96 B 1.10319f
C398 VTAIL.n97 B 0.020444f
C399 VTAIL.n98 B 0.010986f
C400 VTAIL.n99 B 0.011632f
C401 VTAIL.n100 B 0.025966f
C402 VTAIL.n101 B 0.025966f
C403 VTAIL.n102 B 0.011632f
C404 VTAIL.n103 B 0.010986f
C405 VTAIL.n104 B 0.020444f
C406 VTAIL.n105 B 0.020444f
C407 VTAIL.n106 B 0.010986f
C408 VTAIL.n107 B 0.011632f
C409 VTAIL.n108 B 0.025966f
C410 VTAIL.n109 B 0.025966f
C411 VTAIL.n110 B 0.011632f
C412 VTAIL.n111 B 0.010986f
C413 VTAIL.n112 B 0.020444f
C414 VTAIL.n113 B 0.020444f
C415 VTAIL.n114 B 0.010986f
C416 VTAIL.n115 B 0.011309f
C417 VTAIL.n116 B 0.011309f
C418 VTAIL.n117 B 0.025966f
C419 VTAIL.n118 B 0.025966f
C420 VTAIL.n119 B 0.011632f
C421 VTAIL.n120 B 0.010986f
C422 VTAIL.n121 B 0.020444f
C423 VTAIL.n122 B 0.020444f
C424 VTAIL.n123 B 0.010986f
C425 VTAIL.n124 B 0.011632f
C426 VTAIL.n125 B 0.025966f
C427 VTAIL.n126 B 0.025966f
C428 VTAIL.n127 B 0.011632f
C429 VTAIL.n128 B 0.010986f
C430 VTAIL.n129 B 0.020444f
C431 VTAIL.n130 B 0.020444f
C432 VTAIL.n131 B 0.010986f
C433 VTAIL.n132 B 0.011632f
C434 VTAIL.n133 B 0.025966f
C435 VTAIL.n134 B 0.055968f
C436 VTAIL.n135 B 0.011632f
C437 VTAIL.n136 B 0.010986f
C438 VTAIL.n137 B 0.045858f
C439 VTAIL.n138 B 0.031248f
C440 VTAIL.n139 B 1.44064f
C441 VTAIL.n140 B 0.028598f
C442 VTAIL.n141 B 0.020444f
C443 VTAIL.n142 B 0.010986f
C444 VTAIL.n143 B 0.025966f
C445 VTAIL.n144 B 0.011632f
C446 VTAIL.n145 B 0.020444f
C447 VTAIL.n146 B 0.010986f
C448 VTAIL.n147 B 0.025966f
C449 VTAIL.n148 B 0.011632f
C450 VTAIL.n149 B 0.020444f
C451 VTAIL.n150 B 0.010986f
C452 VTAIL.n151 B 0.025966f
C453 VTAIL.n152 B 0.011632f
C454 VTAIL.n153 B 0.020444f
C455 VTAIL.n154 B 0.010986f
C456 VTAIL.n155 B 0.025966f
C457 VTAIL.n156 B 0.025966f
C458 VTAIL.n157 B 0.011632f
C459 VTAIL.n158 B 0.020444f
C460 VTAIL.n159 B 0.010986f
C461 VTAIL.n160 B 0.025966f
C462 VTAIL.n161 B 0.011632f
C463 VTAIL.n162 B 0.153597f
C464 VTAIL.t1 B 0.043942f
C465 VTAIL.n163 B 0.019474f
C466 VTAIL.n164 B 0.018356f
C467 VTAIL.n165 B 0.010986f
C468 VTAIL.n166 B 1.10319f
C469 VTAIL.n167 B 0.020444f
C470 VTAIL.n168 B 0.010986f
C471 VTAIL.n169 B 0.011632f
C472 VTAIL.n170 B 0.025966f
C473 VTAIL.n171 B 0.025966f
C474 VTAIL.n172 B 0.011632f
C475 VTAIL.n173 B 0.010986f
C476 VTAIL.n174 B 0.020444f
C477 VTAIL.n175 B 0.020444f
C478 VTAIL.n176 B 0.010986f
C479 VTAIL.n177 B 0.011632f
C480 VTAIL.n178 B 0.025966f
C481 VTAIL.n179 B 0.025966f
C482 VTAIL.n180 B 0.011632f
C483 VTAIL.n181 B 0.010986f
C484 VTAIL.n182 B 0.020444f
C485 VTAIL.n183 B 0.020444f
C486 VTAIL.n184 B 0.010986f
C487 VTAIL.n185 B 0.011309f
C488 VTAIL.n186 B 0.011309f
C489 VTAIL.n187 B 0.025966f
C490 VTAIL.n188 B 0.025966f
C491 VTAIL.n189 B 0.011632f
C492 VTAIL.n190 B 0.010986f
C493 VTAIL.n191 B 0.020444f
C494 VTAIL.n192 B 0.020444f
C495 VTAIL.n193 B 0.010986f
C496 VTAIL.n194 B 0.011632f
C497 VTAIL.n195 B 0.025966f
C498 VTAIL.n196 B 0.025966f
C499 VTAIL.n197 B 0.011632f
C500 VTAIL.n198 B 0.010986f
C501 VTAIL.n199 B 0.020444f
C502 VTAIL.n200 B 0.020444f
C503 VTAIL.n201 B 0.010986f
C504 VTAIL.n202 B 0.011632f
C505 VTAIL.n203 B 0.025966f
C506 VTAIL.n204 B 0.055968f
C507 VTAIL.n205 B 0.011632f
C508 VTAIL.n206 B 0.010986f
C509 VTAIL.n207 B 0.045858f
C510 VTAIL.n208 B 0.031248f
C511 VTAIL.n209 B 1.28504f
C512 VTAIL.n210 B 0.028598f
C513 VTAIL.n211 B 0.020444f
C514 VTAIL.n212 B 0.010986f
C515 VTAIL.n213 B 0.025966f
C516 VTAIL.n214 B 0.011632f
C517 VTAIL.n215 B 0.020444f
C518 VTAIL.n216 B 0.010986f
C519 VTAIL.n217 B 0.025966f
C520 VTAIL.n218 B 0.011632f
C521 VTAIL.n219 B 0.020444f
C522 VTAIL.n220 B 0.010986f
C523 VTAIL.n221 B 0.025966f
C524 VTAIL.n222 B 0.011632f
C525 VTAIL.n223 B 0.020444f
C526 VTAIL.n224 B 0.010986f
C527 VTAIL.n225 B 0.025966f
C528 VTAIL.n226 B 0.011632f
C529 VTAIL.n227 B 0.020444f
C530 VTAIL.n228 B 0.010986f
C531 VTAIL.n229 B 0.025966f
C532 VTAIL.n230 B 0.011632f
C533 VTAIL.n231 B 0.153597f
C534 VTAIL.t3 B 0.043942f
C535 VTAIL.n232 B 0.019474f
C536 VTAIL.n233 B 0.018356f
C537 VTAIL.n234 B 0.010986f
C538 VTAIL.n235 B 1.10319f
C539 VTAIL.n236 B 0.020444f
C540 VTAIL.n237 B 0.010986f
C541 VTAIL.n238 B 0.011632f
C542 VTAIL.n239 B 0.025966f
C543 VTAIL.n240 B 0.025966f
C544 VTAIL.n241 B 0.011632f
C545 VTAIL.n242 B 0.010986f
C546 VTAIL.n243 B 0.020444f
C547 VTAIL.n244 B 0.020444f
C548 VTAIL.n245 B 0.010986f
C549 VTAIL.n246 B 0.011632f
C550 VTAIL.n247 B 0.025966f
C551 VTAIL.n248 B 0.025966f
C552 VTAIL.n249 B 0.025966f
C553 VTAIL.n250 B 0.011632f
C554 VTAIL.n251 B 0.010986f
C555 VTAIL.n252 B 0.020444f
C556 VTAIL.n253 B 0.020444f
C557 VTAIL.n254 B 0.010986f
C558 VTAIL.n255 B 0.011309f
C559 VTAIL.n256 B 0.011309f
C560 VTAIL.n257 B 0.025966f
C561 VTAIL.n258 B 0.025966f
C562 VTAIL.n259 B 0.011632f
C563 VTAIL.n260 B 0.010986f
C564 VTAIL.n261 B 0.020444f
C565 VTAIL.n262 B 0.020444f
C566 VTAIL.n263 B 0.010986f
C567 VTAIL.n264 B 0.011632f
C568 VTAIL.n265 B 0.025966f
C569 VTAIL.n266 B 0.025966f
C570 VTAIL.n267 B 0.011632f
C571 VTAIL.n268 B 0.010986f
C572 VTAIL.n269 B 0.020444f
C573 VTAIL.n270 B 0.020444f
C574 VTAIL.n271 B 0.010986f
C575 VTAIL.n272 B 0.011632f
C576 VTAIL.n273 B 0.025966f
C577 VTAIL.n274 B 0.055968f
C578 VTAIL.n275 B 0.011632f
C579 VTAIL.n276 B 0.010986f
C580 VTAIL.n277 B 0.045858f
C581 VTAIL.n278 B 0.031248f
C582 VTAIL.n279 B 1.21136f
C583 VN.t0 B 3.00139f
C584 VN.t1 B 3.48994f
.ends

