* NGSPICE file created from diff_pair_sample_0684.ext - technology: sky130A

.subckt diff_pair_sample_0684 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=4.0365 pd=21.48 as=4.0365 ps=21.48 w=10.35 l=3.25
X1 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.0365 pd=21.48 as=4.0365 ps=21.48 w=10.35 l=3.25
X2 VDD2.t0 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=4.0365 pd=21.48 as=4.0365 ps=21.48 w=10.35 l=3.25
X3 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.0365 pd=21.48 as=4.0365 ps=21.48 w=10.35 l=3.25
X4 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=4.0365 pd=21.48 as=0 ps=0 w=10.35 l=3.25
X5 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=4.0365 pd=21.48 as=0 ps=0 w=10.35 l=3.25
X6 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.0365 pd=21.48 as=0 ps=0 w=10.35 l=3.25
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.0365 pd=21.48 as=0 ps=0 w=10.35 l=3.25
R0 VN VN.t1 160.575
R1 VN VN.t0 116.064
R2 VTAIL.n1 VTAIL.t3 48.2991
R3 VTAIL.n3 VTAIL.t2 48.2988
R4 VTAIL.n0 VTAIL.t1 48.2988
R5 VTAIL.n2 VTAIL.t0 48.2988
R6 VTAIL.n1 VTAIL.n0 27.4617
R7 VTAIL.n3 VTAIL.n2 24.3755
R8 VTAIL.n2 VTAIL.n1 2.01343
R9 VTAIL VTAIL.n0 1.30007
R10 VTAIL VTAIL.n3 0.713862
R11 VDD2.n0 VDD2.t1 103.731
R12 VDD2.n0 VDD2.t0 64.9776
R13 VDD2 VDD2.n0 0.830241
R14 B.n661 B.n660 585
R15 B.n662 B.n661 585
R16 B.n266 B.n97 585
R17 B.n265 B.n264 585
R18 B.n263 B.n262 585
R19 B.n261 B.n260 585
R20 B.n259 B.n258 585
R21 B.n257 B.n256 585
R22 B.n255 B.n254 585
R23 B.n253 B.n252 585
R24 B.n251 B.n250 585
R25 B.n249 B.n248 585
R26 B.n247 B.n246 585
R27 B.n245 B.n244 585
R28 B.n243 B.n242 585
R29 B.n241 B.n240 585
R30 B.n239 B.n238 585
R31 B.n237 B.n236 585
R32 B.n235 B.n234 585
R33 B.n233 B.n232 585
R34 B.n231 B.n230 585
R35 B.n229 B.n228 585
R36 B.n227 B.n226 585
R37 B.n225 B.n224 585
R38 B.n223 B.n222 585
R39 B.n221 B.n220 585
R40 B.n219 B.n218 585
R41 B.n217 B.n216 585
R42 B.n215 B.n214 585
R43 B.n213 B.n212 585
R44 B.n211 B.n210 585
R45 B.n209 B.n208 585
R46 B.n207 B.n206 585
R47 B.n205 B.n204 585
R48 B.n203 B.n202 585
R49 B.n201 B.n200 585
R50 B.n199 B.n198 585
R51 B.n197 B.n196 585
R52 B.n195 B.n194 585
R53 B.n193 B.n192 585
R54 B.n191 B.n190 585
R55 B.n189 B.n188 585
R56 B.n187 B.n186 585
R57 B.n185 B.n184 585
R58 B.n183 B.n182 585
R59 B.n181 B.n180 585
R60 B.n179 B.n178 585
R61 B.n176 B.n175 585
R62 B.n174 B.n173 585
R63 B.n172 B.n171 585
R64 B.n170 B.n169 585
R65 B.n168 B.n167 585
R66 B.n166 B.n165 585
R67 B.n164 B.n163 585
R68 B.n162 B.n161 585
R69 B.n160 B.n159 585
R70 B.n158 B.n157 585
R71 B.n156 B.n155 585
R72 B.n154 B.n153 585
R73 B.n152 B.n151 585
R74 B.n150 B.n149 585
R75 B.n148 B.n147 585
R76 B.n146 B.n145 585
R77 B.n144 B.n143 585
R78 B.n142 B.n141 585
R79 B.n140 B.n139 585
R80 B.n138 B.n137 585
R81 B.n136 B.n135 585
R82 B.n134 B.n133 585
R83 B.n132 B.n131 585
R84 B.n130 B.n129 585
R85 B.n128 B.n127 585
R86 B.n126 B.n125 585
R87 B.n124 B.n123 585
R88 B.n122 B.n121 585
R89 B.n120 B.n119 585
R90 B.n118 B.n117 585
R91 B.n116 B.n115 585
R92 B.n114 B.n113 585
R93 B.n112 B.n111 585
R94 B.n110 B.n109 585
R95 B.n108 B.n107 585
R96 B.n106 B.n105 585
R97 B.n104 B.n103 585
R98 B.n659 B.n55 585
R99 B.n663 B.n55 585
R100 B.n658 B.n54 585
R101 B.n664 B.n54 585
R102 B.n657 B.n656 585
R103 B.n656 B.n50 585
R104 B.n655 B.n49 585
R105 B.n670 B.n49 585
R106 B.n654 B.n48 585
R107 B.n671 B.n48 585
R108 B.n653 B.n47 585
R109 B.n672 B.n47 585
R110 B.n652 B.n651 585
R111 B.n651 B.n43 585
R112 B.n650 B.n42 585
R113 B.n678 B.n42 585
R114 B.n649 B.n41 585
R115 B.n679 B.n41 585
R116 B.n648 B.n40 585
R117 B.n680 B.n40 585
R118 B.n647 B.n646 585
R119 B.n646 B.n36 585
R120 B.n645 B.n35 585
R121 B.n686 B.n35 585
R122 B.n644 B.n34 585
R123 B.n687 B.n34 585
R124 B.n643 B.n33 585
R125 B.n688 B.n33 585
R126 B.n642 B.n641 585
R127 B.n641 B.n29 585
R128 B.n640 B.n28 585
R129 B.n694 B.n28 585
R130 B.n639 B.n27 585
R131 B.n695 B.n27 585
R132 B.n638 B.n26 585
R133 B.n696 B.n26 585
R134 B.n637 B.n636 585
R135 B.n636 B.n22 585
R136 B.n635 B.n21 585
R137 B.n702 B.n21 585
R138 B.n634 B.n20 585
R139 B.n703 B.n20 585
R140 B.n633 B.n19 585
R141 B.n704 B.n19 585
R142 B.n632 B.n631 585
R143 B.n631 B.n18 585
R144 B.n630 B.n14 585
R145 B.n710 B.n14 585
R146 B.n629 B.n13 585
R147 B.n711 B.n13 585
R148 B.n628 B.n12 585
R149 B.n712 B.n12 585
R150 B.n627 B.n626 585
R151 B.n626 B.n8 585
R152 B.n625 B.n7 585
R153 B.n718 B.n7 585
R154 B.n624 B.n6 585
R155 B.n719 B.n6 585
R156 B.n623 B.n5 585
R157 B.n720 B.n5 585
R158 B.n622 B.n621 585
R159 B.n621 B.n4 585
R160 B.n620 B.n267 585
R161 B.n620 B.n619 585
R162 B.n610 B.n268 585
R163 B.n269 B.n268 585
R164 B.n612 B.n611 585
R165 B.n613 B.n612 585
R166 B.n609 B.n274 585
R167 B.n274 B.n273 585
R168 B.n608 B.n607 585
R169 B.n607 B.n606 585
R170 B.n276 B.n275 585
R171 B.n599 B.n276 585
R172 B.n598 B.n597 585
R173 B.n600 B.n598 585
R174 B.n596 B.n281 585
R175 B.n281 B.n280 585
R176 B.n595 B.n594 585
R177 B.n594 B.n593 585
R178 B.n283 B.n282 585
R179 B.n284 B.n283 585
R180 B.n586 B.n585 585
R181 B.n587 B.n586 585
R182 B.n584 B.n289 585
R183 B.n289 B.n288 585
R184 B.n583 B.n582 585
R185 B.n582 B.n581 585
R186 B.n291 B.n290 585
R187 B.n292 B.n291 585
R188 B.n574 B.n573 585
R189 B.n575 B.n574 585
R190 B.n572 B.n297 585
R191 B.n297 B.n296 585
R192 B.n571 B.n570 585
R193 B.n570 B.n569 585
R194 B.n299 B.n298 585
R195 B.n300 B.n299 585
R196 B.n562 B.n561 585
R197 B.n563 B.n562 585
R198 B.n560 B.n304 585
R199 B.n308 B.n304 585
R200 B.n559 B.n558 585
R201 B.n558 B.n557 585
R202 B.n306 B.n305 585
R203 B.n307 B.n306 585
R204 B.n550 B.n549 585
R205 B.n551 B.n550 585
R206 B.n548 B.n313 585
R207 B.n313 B.n312 585
R208 B.n547 B.n546 585
R209 B.n546 B.n545 585
R210 B.n315 B.n314 585
R211 B.n316 B.n315 585
R212 B.n538 B.n537 585
R213 B.n539 B.n538 585
R214 B.n536 B.n321 585
R215 B.n321 B.n320 585
R216 B.n530 B.n529 585
R217 B.n528 B.n364 585
R218 B.n527 B.n363 585
R219 B.n532 B.n363 585
R220 B.n526 B.n525 585
R221 B.n524 B.n523 585
R222 B.n522 B.n521 585
R223 B.n520 B.n519 585
R224 B.n518 B.n517 585
R225 B.n516 B.n515 585
R226 B.n514 B.n513 585
R227 B.n512 B.n511 585
R228 B.n510 B.n509 585
R229 B.n508 B.n507 585
R230 B.n506 B.n505 585
R231 B.n504 B.n503 585
R232 B.n502 B.n501 585
R233 B.n500 B.n499 585
R234 B.n498 B.n497 585
R235 B.n496 B.n495 585
R236 B.n494 B.n493 585
R237 B.n492 B.n491 585
R238 B.n490 B.n489 585
R239 B.n488 B.n487 585
R240 B.n486 B.n485 585
R241 B.n484 B.n483 585
R242 B.n482 B.n481 585
R243 B.n480 B.n479 585
R244 B.n478 B.n477 585
R245 B.n476 B.n475 585
R246 B.n474 B.n473 585
R247 B.n472 B.n471 585
R248 B.n470 B.n469 585
R249 B.n468 B.n467 585
R250 B.n466 B.n465 585
R251 B.n464 B.n463 585
R252 B.n462 B.n461 585
R253 B.n460 B.n459 585
R254 B.n458 B.n457 585
R255 B.n456 B.n455 585
R256 B.n454 B.n453 585
R257 B.n452 B.n451 585
R258 B.n450 B.n449 585
R259 B.n448 B.n447 585
R260 B.n446 B.n445 585
R261 B.n444 B.n443 585
R262 B.n442 B.n441 585
R263 B.n439 B.n438 585
R264 B.n437 B.n436 585
R265 B.n435 B.n434 585
R266 B.n433 B.n432 585
R267 B.n431 B.n430 585
R268 B.n429 B.n428 585
R269 B.n427 B.n426 585
R270 B.n425 B.n424 585
R271 B.n423 B.n422 585
R272 B.n421 B.n420 585
R273 B.n419 B.n418 585
R274 B.n417 B.n416 585
R275 B.n415 B.n414 585
R276 B.n413 B.n412 585
R277 B.n411 B.n410 585
R278 B.n409 B.n408 585
R279 B.n407 B.n406 585
R280 B.n405 B.n404 585
R281 B.n403 B.n402 585
R282 B.n401 B.n400 585
R283 B.n399 B.n398 585
R284 B.n397 B.n396 585
R285 B.n395 B.n394 585
R286 B.n393 B.n392 585
R287 B.n391 B.n390 585
R288 B.n389 B.n388 585
R289 B.n387 B.n386 585
R290 B.n385 B.n384 585
R291 B.n383 B.n382 585
R292 B.n381 B.n380 585
R293 B.n379 B.n378 585
R294 B.n377 B.n376 585
R295 B.n375 B.n374 585
R296 B.n373 B.n372 585
R297 B.n371 B.n370 585
R298 B.n323 B.n322 585
R299 B.n535 B.n534 585
R300 B.n319 B.n318 585
R301 B.n320 B.n319 585
R302 B.n541 B.n540 585
R303 B.n540 B.n539 585
R304 B.n542 B.n317 585
R305 B.n317 B.n316 585
R306 B.n544 B.n543 585
R307 B.n545 B.n544 585
R308 B.n311 B.n310 585
R309 B.n312 B.n311 585
R310 B.n553 B.n552 585
R311 B.n552 B.n551 585
R312 B.n554 B.n309 585
R313 B.n309 B.n307 585
R314 B.n556 B.n555 585
R315 B.n557 B.n556 585
R316 B.n303 B.n302 585
R317 B.n308 B.n303 585
R318 B.n565 B.n564 585
R319 B.n564 B.n563 585
R320 B.n566 B.n301 585
R321 B.n301 B.n300 585
R322 B.n568 B.n567 585
R323 B.n569 B.n568 585
R324 B.n295 B.n294 585
R325 B.n296 B.n295 585
R326 B.n577 B.n576 585
R327 B.n576 B.n575 585
R328 B.n578 B.n293 585
R329 B.n293 B.n292 585
R330 B.n580 B.n579 585
R331 B.n581 B.n580 585
R332 B.n287 B.n286 585
R333 B.n288 B.n287 585
R334 B.n589 B.n588 585
R335 B.n588 B.n587 585
R336 B.n590 B.n285 585
R337 B.n285 B.n284 585
R338 B.n592 B.n591 585
R339 B.n593 B.n592 585
R340 B.n279 B.n278 585
R341 B.n280 B.n279 585
R342 B.n602 B.n601 585
R343 B.n601 B.n600 585
R344 B.n603 B.n277 585
R345 B.n599 B.n277 585
R346 B.n605 B.n604 585
R347 B.n606 B.n605 585
R348 B.n272 B.n271 585
R349 B.n273 B.n272 585
R350 B.n615 B.n614 585
R351 B.n614 B.n613 585
R352 B.n616 B.n270 585
R353 B.n270 B.n269 585
R354 B.n618 B.n617 585
R355 B.n619 B.n618 585
R356 B.n2 B.n0 585
R357 B.n4 B.n2 585
R358 B.n3 B.n1 585
R359 B.n719 B.n3 585
R360 B.n717 B.n716 585
R361 B.n718 B.n717 585
R362 B.n715 B.n9 585
R363 B.n9 B.n8 585
R364 B.n714 B.n713 585
R365 B.n713 B.n712 585
R366 B.n11 B.n10 585
R367 B.n711 B.n11 585
R368 B.n709 B.n708 585
R369 B.n710 B.n709 585
R370 B.n707 B.n15 585
R371 B.n18 B.n15 585
R372 B.n706 B.n705 585
R373 B.n705 B.n704 585
R374 B.n17 B.n16 585
R375 B.n703 B.n17 585
R376 B.n701 B.n700 585
R377 B.n702 B.n701 585
R378 B.n699 B.n23 585
R379 B.n23 B.n22 585
R380 B.n698 B.n697 585
R381 B.n697 B.n696 585
R382 B.n25 B.n24 585
R383 B.n695 B.n25 585
R384 B.n693 B.n692 585
R385 B.n694 B.n693 585
R386 B.n691 B.n30 585
R387 B.n30 B.n29 585
R388 B.n690 B.n689 585
R389 B.n689 B.n688 585
R390 B.n32 B.n31 585
R391 B.n687 B.n32 585
R392 B.n685 B.n684 585
R393 B.n686 B.n685 585
R394 B.n683 B.n37 585
R395 B.n37 B.n36 585
R396 B.n682 B.n681 585
R397 B.n681 B.n680 585
R398 B.n39 B.n38 585
R399 B.n679 B.n39 585
R400 B.n677 B.n676 585
R401 B.n678 B.n677 585
R402 B.n675 B.n44 585
R403 B.n44 B.n43 585
R404 B.n674 B.n673 585
R405 B.n673 B.n672 585
R406 B.n46 B.n45 585
R407 B.n671 B.n46 585
R408 B.n669 B.n668 585
R409 B.n670 B.n669 585
R410 B.n667 B.n51 585
R411 B.n51 B.n50 585
R412 B.n666 B.n665 585
R413 B.n665 B.n664 585
R414 B.n53 B.n52 585
R415 B.n663 B.n53 585
R416 B.n722 B.n721 585
R417 B.n721 B.n720 585
R418 B.n530 B.n319 535.745
R419 B.n103 B.n53 535.745
R420 B.n534 B.n321 535.745
R421 B.n661 B.n55 535.745
R422 B.n368 B.t13 285.603
R423 B.n365 B.t2 285.603
R424 B.n101 B.t6 285.603
R425 B.n98 B.t10 285.603
R426 B.n662 B.n96 256.663
R427 B.n662 B.n95 256.663
R428 B.n662 B.n94 256.663
R429 B.n662 B.n93 256.663
R430 B.n662 B.n92 256.663
R431 B.n662 B.n91 256.663
R432 B.n662 B.n90 256.663
R433 B.n662 B.n89 256.663
R434 B.n662 B.n88 256.663
R435 B.n662 B.n87 256.663
R436 B.n662 B.n86 256.663
R437 B.n662 B.n85 256.663
R438 B.n662 B.n84 256.663
R439 B.n662 B.n83 256.663
R440 B.n662 B.n82 256.663
R441 B.n662 B.n81 256.663
R442 B.n662 B.n80 256.663
R443 B.n662 B.n79 256.663
R444 B.n662 B.n78 256.663
R445 B.n662 B.n77 256.663
R446 B.n662 B.n76 256.663
R447 B.n662 B.n75 256.663
R448 B.n662 B.n74 256.663
R449 B.n662 B.n73 256.663
R450 B.n662 B.n72 256.663
R451 B.n662 B.n71 256.663
R452 B.n662 B.n70 256.663
R453 B.n662 B.n69 256.663
R454 B.n662 B.n68 256.663
R455 B.n662 B.n67 256.663
R456 B.n662 B.n66 256.663
R457 B.n662 B.n65 256.663
R458 B.n662 B.n64 256.663
R459 B.n662 B.n63 256.663
R460 B.n662 B.n62 256.663
R461 B.n662 B.n61 256.663
R462 B.n662 B.n60 256.663
R463 B.n662 B.n59 256.663
R464 B.n662 B.n58 256.663
R465 B.n662 B.n57 256.663
R466 B.n662 B.n56 256.663
R467 B.n532 B.n531 256.663
R468 B.n532 B.n324 256.663
R469 B.n532 B.n325 256.663
R470 B.n532 B.n326 256.663
R471 B.n532 B.n327 256.663
R472 B.n532 B.n328 256.663
R473 B.n532 B.n329 256.663
R474 B.n532 B.n330 256.663
R475 B.n532 B.n331 256.663
R476 B.n532 B.n332 256.663
R477 B.n532 B.n333 256.663
R478 B.n532 B.n334 256.663
R479 B.n532 B.n335 256.663
R480 B.n532 B.n336 256.663
R481 B.n532 B.n337 256.663
R482 B.n532 B.n338 256.663
R483 B.n532 B.n339 256.663
R484 B.n532 B.n340 256.663
R485 B.n532 B.n341 256.663
R486 B.n532 B.n342 256.663
R487 B.n532 B.n343 256.663
R488 B.n532 B.n344 256.663
R489 B.n532 B.n345 256.663
R490 B.n532 B.n346 256.663
R491 B.n532 B.n347 256.663
R492 B.n532 B.n348 256.663
R493 B.n532 B.n349 256.663
R494 B.n532 B.n350 256.663
R495 B.n532 B.n351 256.663
R496 B.n532 B.n352 256.663
R497 B.n532 B.n353 256.663
R498 B.n532 B.n354 256.663
R499 B.n532 B.n355 256.663
R500 B.n532 B.n356 256.663
R501 B.n532 B.n357 256.663
R502 B.n532 B.n358 256.663
R503 B.n532 B.n359 256.663
R504 B.n532 B.n360 256.663
R505 B.n532 B.n361 256.663
R506 B.n532 B.n362 256.663
R507 B.n533 B.n532 256.663
R508 B.n540 B.n319 163.367
R509 B.n540 B.n317 163.367
R510 B.n544 B.n317 163.367
R511 B.n544 B.n311 163.367
R512 B.n552 B.n311 163.367
R513 B.n552 B.n309 163.367
R514 B.n556 B.n309 163.367
R515 B.n556 B.n303 163.367
R516 B.n564 B.n303 163.367
R517 B.n564 B.n301 163.367
R518 B.n568 B.n301 163.367
R519 B.n568 B.n295 163.367
R520 B.n576 B.n295 163.367
R521 B.n576 B.n293 163.367
R522 B.n580 B.n293 163.367
R523 B.n580 B.n287 163.367
R524 B.n588 B.n287 163.367
R525 B.n588 B.n285 163.367
R526 B.n592 B.n285 163.367
R527 B.n592 B.n279 163.367
R528 B.n601 B.n279 163.367
R529 B.n601 B.n277 163.367
R530 B.n605 B.n277 163.367
R531 B.n605 B.n272 163.367
R532 B.n614 B.n272 163.367
R533 B.n614 B.n270 163.367
R534 B.n618 B.n270 163.367
R535 B.n618 B.n2 163.367
R536 B.n721 B.n2 163.367
R537 B.n721 B.n3 163.367
R538 B.n717 B.n3 163.367
R539 B.n717 B.n9 163.367
R540 B.n713 B.n9 163.367
R541 B.n713 B.n11 163.367
R542 B.n709 B.n11 163.367
R543 B.n709 B.n15 163.367
R544 B.n705 B.n15 163.367
R545 B.n705 B.n17 163.367
R546 B.n701 B.n17 163.367
R547 B.n701 B.n23 163.367
R548 B.n697 B.n23 163.367
R549 B.n697 B.n25 163.367
R550 B.n693 B.n25 163.367
R551 B.n693 B.n30 163.367
R552 B.n689 B.n30 163.367
R553 B.n689 B.n32 163.367
R554 B.n685 B.n32 163.367
R555 B.n685 B.n37 163.367
R556 B.n681 B.n37 163.367
R557 B.n681 B.n39 163.367
R558 B.n677 B.n39 163.367
R559 B.n677 B.n44 163.367
R560 B.n673 B.n44 163.367
R561 B.n673 B.n46 163.367
R562 B.n669 B.n46 163.367
R563 B.n669 B.n51 163.367
R564 B.n665 B.n51 163.367
R565 B.n665 B.n53 163.367
R566 B.n364 B.n363 163.367
R567 B.n525 B.n363 163.367
R568 B.n523 B.n522 163.367
R569 B.n519 B.n518 163.367
R570 B.n515 B.n514 163.367
R571 B.n511 B.n510 163.367
R572 B.n507 B.n506 163.367
R573 B.n503 B.n502 163.367
R574 B.n499 B.n498 163.367
R575 B.n495 B.n494 163.367
R576 B.n491 B.n490 163.367
R577 B.n487 B.n486 163.367
R578 B.n483 B.n482 163.367
R579 B.n479 B.n478 163.367
R580 B.n475 B.n474 163.367
R581 B.n471 B.n470 163.367
R582 B.n467 B.n466 163.367
R583 B.n463 B.n462 163.367
R584 B.n459 B.n458 163.367
R585 B.n455 B.n454 163.367
R586 B.n451 B.n450 163.367
R587 B.n447 B.n446 163.367
R588 B.n443 B.n442 163.367
R589 B.n438 B.n437 163.367
R590 B.n434 B.n433 163.367
R591 B.n430 B.n429 163.367
R592 B.n426 B.n425 163.367
R593 B.n422 B.n421 163.367
R594 B.n418 B.n417 163.367
R595 B.n414 B.n413 163.367
R596 B.n410 B.n409 163.367
R597 B.n406 B.n405 163.367
R598 B.n402 B.n401 163.367
R599 B.n398 B.n397 163.367
R600 B.n394 B.n393 163.367
R601 B.n390 B.n389 163.367
R602 B.n386 B.n385 163.367
R603 B.n382 B.n381 163.367
R604 B.n378 B.n377 163.367
R605 B.n374 B.n373 163.367
R606 B.n370 B.n323 163.367
R607 B.n538 B.n321 163.367
R608 B.n538 B.n315 163.367
R609 B.n546 B.n315 163.367
R610 B.n546 B.n313 163.367
R611 B.n550 B.n313 163.367
R612 B.n550 B.n306 163.367
R613 B.n558 B.n306 163.367
R614 B.n558 B.n304 163.367
R615 B.n562 B.n304 163.367
R616 B.n562 B.n299 163.367
R617 B.n570 B.n299 163.367
R618 B.n570 B.n297 163.367
R619 B.n574 B.n297 163.367
R620 B.n574 B.n291 163.367
R621 B.n582 B.n291 163.367
R622 B.n582 B.n289 163.367
R623 B.n586 B.n289 163.367
R624 B.n586 B.n283 163.367
R625 B.n594 B.n283 163.367
R626 B.n594 B.n281 163.367
R627 B.n598 B.n281 163.367
R628 B.n598 B.n276 163.367
R629 B.n607 B.n276 163.367
R630 B.n607 B.n274 163.367
R631 B.n612 B.n274 163.367
R632 B.n612 B.n268 163.367
R633 B.n620 B.n268 163.367
R634 B.n621 B.n620 163.367
R635 B.n621 B.n5 163.367
R636 B.n6 B.n5 163.367
R637 B.n7 B.n6 163.367
R638 B.n626 B.n7 163.367
R639 B.n626 B.n12 163.367
R640 B.n13 B.n12 163.367
R641 B.n14 B.n13 163.367
R642 B.n631 B.n14 163.367
R643 B.n631 B.n19 163.367
R644 B.n20 B.n19 163.367
R645 B.n21 B.n20 163.367
R646 B.n636 B.n21 163.367
R647 B.n636 B.n26 163.367
R648 B.n27 B.n26 163.367
R649 B.n28 B.n27 163.367
R650 B.n641 B.n28 163.367
R651 B.n641 B.n33 163.367
R652 B.n34 B.n33 163.367
R653 B.n35 B.n34 163.367
R654 B.n646 B.n35 163.367
R655 B.n646 B.n40 163.367
R656 B.n41 B.n40 163.367
R657 B.n42 B.n41 163.367
R658 B.n651 B.n42 163.367
R659 B.n651 B.n47 163.367
R660 B.n48 B.n47 163.367
R661 B.n49 B.n48 163.367
R662 B.n656 B.n49 163.367
R663 B.n656 B.n54 163.367
R664 B.n55 B.n54 163.367
R665 B.n107 B.n106 163.367
R666 B.n111 B.n110 163.367
R667 B.n115 B.n114 163.367
R668 B.n119 B.n118 163.367
R669 B.n123 B.n122 163.367
R670 B.n127 B.n126 163.367
R671 B.n131 B.n130 163.367
R672 B.n135 B.n134 163.367
R673 B.n139 B.n138 163.367
R674 B.n143 B.n142 163.367
R675 B.n147 B.n146 163.367
R676 B.n151 B.n150 163.367
R677 B.n155 B.n154 163.367
R678 B.n159 B.n158 163.367
R679 B.n163 B.n162 163.367
R680 B.n167 B.n166 163.367
R681 B.n171 B.n170 163.367
R682 B.n175 B.n174 163.367
R683 B.n180 B.n179 163.367
R684 B.n184 B.n183 163.367
R685 B.n188 B.n187 163.367
R686 B.n192 B.n191 163.367
R687 B.n196 B.n195 163.367
R688 B.n200 B.n199 163.367
R689 B.n204 B.n203 163.367
R690 B.n208 B.n207 163.367
R691 B.n212 B.n211 163.367
R692 B.n216 B.n215 163.367
R693 B.n220 B.n219 163.367
R694 B.n224 B.n223 163.367
R695 B.n228 B.n227 163.367
R696 B.n232 B.n231 163.367
R697 B.n236 B.n235 163.367
R698 B.n240 B.n239 163.367
R699 B.n244 B.n243 163.367
R700 B.n248 B.n247 163.367
R701 B.n252 B.n251 163.367
R702 B.n256 B.n255 163.367
R703 B.n260 B.n259 163.367
R704 B.n264 B.n263 163.367
R705 B.n661 B.n97 163.367
R706 B.n368 B.t15 140.389
R707 B.n98 B.t11 140.389
R708 B.n365 B.t5 140.377
R709 B.n101 B.t8 140.377
R710 B.n532 B.n320 95.0405
R711 B.n663 B.n662 95.0405
R712 B.n531 B.n530 71.676
R713 B.n525 B.n324 71.676
R714 B.n522 B.n325 71.676
R715 B.n518 B.n326 71.676
R716 B.n514 B.n327 71.676
R717 B.n510 B.n328 71.676
R718 B.n506 B.n329 71.676
R719 B.n502 B.n330 71.676
R720 B.n498 B.n331 71.676
R721 B.n494 B.n332 71.676
R722 B.n490 B.n333 71.676
R723 B.n486 B.n334 71.676
R724 B.n482 B.n335 71.676
R725 B.n478 B.n336 71.676
R726 B.n474 B.n337 71.676
R727 B.n470 B.n338 71.676
R728 B.n466 B.n339 71.676
R729 B.n462 B.n340 71.676
R730 B.n458 B.n341 71.676
R731 B.n454 B.n342 71.676
R732 B.n450 B.n343 71.676
R733 B.n446 B.n344 71.676
R734 B.n442 B.n345 71.676
R735 B.n437 B.n346 71.676
R736 B.n433 B.n347 71.676
R737 B.n429 B.n348 71.676
R738 B.n425 B.n349 71.676
R739 B.n421 B.n350 71.676
R740 B.n417 B.n351 71.676
R741 B.n413 B.n352 71.676
R742 B.n409 B.n353 71.676
R743 B.n405 B.n354 71.676
R744 B.n401 B.n355 71.676
R745 B.n397 B.n356 71.676
R746 B.n393 B.n357 71.676
R747 B.n389 B.n358 71.676
R748 B.n385 B.n359 71.676
R749 B.n381 B.n360 71.676
R750 B.n377 B.n361 71.676
R751 B.n373 B.n362 71.676
R752 B.n533 B.n323 71.676
R753 B.n103 B.n56 71.676
R754 B.n107 B.n57 71.676
R755 B.n111 B.n58 71.676
R756 B.n115 B.n59 71.676
R757 B.n119 B.n60 71.676
R758 B.n123 B.n61 71.676
R759 B.n127 B.n62 71.676
R760 B.n131 B.n63 71.676
R761 B.n135 B.n64 71.676
R762 B.n139 B.n65 71.676
R763 B.n143 B.n66 71.676
R764 B.n147 B.n67 71.676
R765 B.n151 B.n68 71.676
R766 B.n155 B.n69 71.676
R767 B.n159 B.n70 71.676
R768 B.n163 B.n71 71.676
R769 B.n167 B.n72 71.676
R770 B.n171 B.n73 71.676
R771 B.n175 B.n74 71.676
R772 B.n180 B.n75 71.676
R773 B.n184 B.n76 71.676
R774 B.n188 B.n77 71.676
R775 B.n192 B.n78 71.676
R776 B.n196 B.n79 71.676
R777 B.n200 B.n80 71.676
R778 B.n204 B.n81 71.676
R779 B.n208 B.n82 71.676
R780 B.n212 B.n83 71.676
R781 B.n216 B.n84 71.676
R782 B.n220 B.n85 71.676
R783 B.n224 B.n86 71.676
R784 B.n228 B.n87 71.676
R785 B.n232 B.n88 71.676
R786 B.n236 B.n89 71.676
R787 B.n240 B.n90 71.676
R788 B.n244 B.n91 71.676
R789 B.n248 B.n92 71.676
R790 B.n252 B.n93 71.676
R791 B.n256 B.n94 71.676
R792 B.n260 B.n95 71.676
R793 B.n264 B.n96 71.676
R794 B.n97 B.n96 71.676
R795 B.n263 B.n95 71.676
R796 B.n259 B.n94 71.676
R797 B.n255 B.n93 71.676
R798 B.n251 B.n92 71.676
R799 B.n247 B.n91 71.676
R800 B.n243 B.n90 71.676
R801 B.n239 B.n89 71.676
R802 B.n235 B.n88 71.676
R803 B.n231 B.n87 71.676
R804 B.n227 B.n86 71.676
R805 B.n223 B.n85 71.676
R806 B.n219 B.n84 71.676
R807 B.n215 B.n83 71.676
R808 B.n211 B.n82 71.676
R809 B.n207 B.n81 71.676
R810 B.n203 B.n80 71.676
R811 B.n199 B.n79 71.676
R812 B.n195 B.n78 71.676
R813 B.n191 B.n77 71.676
R814 B.n187 B.n76 71.676
R815 B.n183 B.n75 71.676
R816 B.n179 B.n74 71.676
R817 B.n174 B.n73 71.676
R818 B.n170 B.n72 71.676
R819 B.n166 B.n71 71.676
R820 B.n162 B.n70 71.676
R821 B.n158 B.n69 71.676
R822 B.n154 B.n68 71.676
R823 B.n150 B.n67 71.676
R824 B.n146 B.n66 71.676
R825 B.n142 B.n65 71.676
R826 B.n138 B.n64 71.676
R827 B.n134 B.n63 71.676
R828 B.n130 B.n62 71.676
R829 B.n126 B.n61 71.676
R830 B.n122 B.n60 71.676
R831 B.n118 B.n59 71.676
R832 B.n114 B.n58 71.676
R833 B.n110 B.n57 71.676
R834 B.n106 B.n56 71.676
R835 B.n531 B.n364 71.676
R836 B.n523 B.n324 71.676
R837 B.n519 B.n325 71.676
R838 B.n515 B.n326 71.676
R839 B.n511 B.n327 71.676
R840 B.n507 B.n328 71.676
R841 B.n503 B.n329 71.676
R842 B.n499 B.n330 71.676
R843 B.n495 B.n331 71.676
R844 B.n491 B.n332 71.676
R845 B.n487 B.n333 71.676
R846 B.n483 B.n334 71.676
R847 B.n479 B.n335 71.676
R848 B.n475 B.n336 71.676
R849 B.n471 B.n337 71.676
R850 B.n467 B.n338 71.676
R851 B.n463 B.n339 71.676
R852 B.n459 B.n340 71.676
R853 B.n455 B.n341 71.676
R854 B.n451 B.n342 71.676
R855 B.n447 B.n343 71.676
R856 B.n443 B.n344 71.676
R857 B.n438 B.n345 71.676
R858 B.n434 B.n346 71.676
R859 B.n430 B.n347 71.676
R860 B.n426 B.n348 71.676
R861 B.n422 B.n349 71.676
R862 B.n418 B.n350 71.676
R863 B.n414 B.n351 71.676
R864 B.n410 B.n352 71.676
R865 B.n406 B.n353 71.676
R866 B.n402 B.n354 71.676
R867 B.n398 B.n355 71.676
R868 B.n394 B.n356 71.676
R869 B.n390 B.n357 71.676
R870 B.n386 B.n358 71.676
R871 B.n382 B.n359 71.676
R872 B.n378 B.n360 71.676
R873 B.n374 B.n361 71.676
R874 B.n370 B.n362 71.676
R875 B.n534 B.n533 71.676
R876 B.n369 B.t14 70.9595
R877 B.n99 B.t12 70.9595
R878 B.n366 B.t4 70.9468
R879 B.n102 B.t9 70.9468
R880 B.n369 B.n368 69.4308
R881 B.n366 B.n365 69.4308
R882 B.n102 B.n101 69.4308
R883 B.n99 B.n98 69.4308
R884 B.n440 B.n369 59.5399
R885 B.n367 B.n366 59.5399
R886 B.n177 B.n102 59.5399
R887 B.n100 B.n99 59.5399
R888 B.n539 B.n320 47.8725
R889 B.n539 B.n316 47.8725
R890 B.n545 B.n316 47.8725
R891 B.n545 B.n312 47.8725
R892 B.n551 B.n312 47.8725
R893 B.n551 B.n307 47.8725
R894 B.n557 B.n307 47.8725
R895 B.n557 B.n308 47.8725
R896 B.n563 B.n300 47.8725
R897 B.n569 B.n300 47.8725
R898 B.n569 B.n296 47.8725
R899 B.n575 B.n296 47.8725
R900 B.n575 B.n292 47.8725
R901 B.n581 B.n292 47.8725
R902 B.n581 B.n288 47.8725
R903 B.n587 B.n288 47.8725
R904 B.n587 B.n284 47.8725
R905 B.n593 B.n284 47.8725
R906 B.n593 B.n280 47.8725
R907 B.n600 B.n280 47.8725
R908 B.n600 B.n599 47.8725
R909 B.n606 B.n273 47.8725
R910 B.n613 B.n273 47.8725
R911 B.n613 B.n269 47.8725
R912 B.n619 B.n269 47.8725
R913 B.n619 B.n4 47.8725
R914 B.n720 B.n4 47.8725
R915 B.n720 B.n719 47.8725
R916 B.n719 B.n718 47.8725
R917 B.n718 B.n8 47.8725
R918 B.n712 B.n8 47.8725
R919 B.n712 B.n711 47.8725
R920 B.n711 B.n710 47.8725
R921 B.n704 B.n18 47.8725
R922 B.n704 B.n703 47.8725
R923 B.n703 B.n702 47.8725
R924 B.n702 B.n22 47.8725
R925 B.n696 B.n22 47.8725
R926 B.n696 B.n695 47.8725
R927 B.n695 B.n694 47.8725
R928 B.n694 B.n29 47.8725
R929 B.n688 B.n29 47.8725
R930 B.n688 B.n687 47.8725
R931 B.n687 B.n686 47.8725
R932 B.n686 B.n36 47.8725
R933 B.n680 B.n36 47.8725
R934 B.n679 B.n678 47.8725
R935 B.n678 B.n43 47.8725
R936 B.n672 B.n43 47.8725
R937 B.n672 B.n671 47.8725
R938 B.n671 B.n670 47.8725
R939 B.n670 B.n50 47.8725
R940 B.n664 B.n50 47.8725
R941 B.n664 B.n663 47.8725
R942 B.n606 B.t1 41.5365
R943 B.n710 B.t0 41.5365
R944 B.n660 B.n659 34.8103
R945 B.n104 B.n52 34.8103
R946 B.n536 B.n535 34.8103
R947 B.n529 B.n318 34.8103
R948 B.n563 B.t3 28.8645
R949 B.n680 B.t7 28.8645
R950 B.n308 B.t3 19.0085
R951 B.t7 B.n679 19.0085
R952 B B.n722 18.0485
R953 B.n105 B.n104 10.6151
R954 B.n108 B.n105 10.6151
R955 B.n109 B.n108 10.6151
R956 B.n112 B.n109 10.6151
R957 B.n113 B.n112 10.6151
R958 B.n116 B.n113 10.6151
R959 B.n117 B.n116 10.6151
R960 B.n120 B.n117 10.6151
R961 B.n121 B.n120 10.6151
R962 B.n124 B.n121 10.6151
R963 B.n125 B.n124 10.6151
R964 B.n128 B.n125 10.6151
R965 B.n129 B.n128 10.6151
R966 B.n132 B.n129 10.6151
R967 B.n133 B.n132 10.6151
R968 B.n136 B.n133 10.6151
R969 B.n137 B.n136 10.6151
R970 B.n140 B.n137 10.6151
R971 B.n141 B.n140 10.6151
R972 B.n144 B.n141 10.6151
R973 B.n145 B.n144 10.6151
R974 B.n148 B.n145 10.6151
R975 B.n149 B.n148 10.6151
R976 B.n152 B.n149 10.6151
R977 B.n153 B.n152 10.6151
R978 B.n156 B.n153 10.6151
R979 B.n157 B.n156 10.6151
R980 B.n160 B.n157 10.6151
R981 B.n161 B.n160 10.6151
R982 B.n164 B.n161 10.6151
R983 B.n165 B.n164 10.6151
R984 B.n168 B.n165 10.6151
R985 B.n169 B.n168 10.6151
R986 B.n172 B.n169 10.6151
R987 B.n173 B.n172 10.6151
R988 B.n176 B.n173 10.6151
R989 B.n181 B.n178 10.6151
R990 B.n182 B.n181 10.6151
R991 B.n185 B.n182 10.6151
R992 B.n186 B.n185 10.6151
R993 B.n189 B.n186 10.6151
R994 B.n190 B.n189 10.6151
R995 B.n193 B.n190 10.6151
R996 B.n194 B.n193 10.6151
R997 B.n198 B.n197 10.6151
R998 B.n201 B.n198 10.6151
R999 B.n202 B.n201 10.6151
R1000 B.n205 B.n202 10.6151
R1001 B.n206 B.n205 10.6151
R1002 B.n209 B.n206 10.6151
R1003 B.n210 B.n209 10.6151
R1004 B.n213 B.n210 10.6151
R1005 B.n214 B.n213 10.6151
R1006 B.n217 B.n214 10.6151
R1007 B.n218 B.n217 10.6151
R1008 B.n221 B.n218 10.6151
R1009 B.n222 B.n221 10.6151
R1010 B.n225 B.n222 10.6151
R1011 B.n226 B.n225 10.6151
R1012 B.n229 B.n226 10.6151
R1013 B.n230 B.n229 10.6151
R1014 B.n233 B.n230 10.6151
R1015 B.n234 B.n233 10.6151
R1016 B.n237 B.n234 10.6151
R1017 B.n238 B.n237 10.6151
R1018 B.n241 B.n238 10.6151
R1019 B.n242 B.n241 10.6151
R1020 B.n245 B.n242 10.6151
R1021 B.n246 B.n245 10.6151
R1022 B.n249 B.n246 10.6151
R1023 B.n250 B.n249 10.6151
R1024 B.n253 B.n250 10.6151
R1025 B.n254 B.n253 10.6151
R1026 B.n257 B.n254 10.6151
R1027 B.n258 B.n257 10.6151
R1028 B.n261 B.n258 10.6151
R1029 B.n262 B.n261 10.6151
R1030 B.n265 B.n262 10.6151
R1031 B.n266 B.n265 10.6151
R1032 B.n660 B.n266 10.6151
R1033 B.n537 B.n536 10.6151
R1034 B.n537 B.n314 10.6151
R1035 B.n547 B.n314 10.6151
R1036 B.n548 B.n547 10.6151
R1037 B.n549 B.n548 10.6151
R1038 B.n549 B.n305 10.6151
R1039 B.n559 B.n305 10.6151
R1040 B.n560 B.n559 10.6151
R1041 B.n561 B.n560 10.6151
R1042 B.n561 B.n298 10.6151
R1043 B.n571 B.n298 10.6151
R1044 B.n572 B.n571 10.6151
R1045 B.n573 B.n572 10.6151
R1046 B.n573 B.n290 10.6151
R1047 B.n583 B.n290 10.6151
R1048 B.n584 B.n583 10.6151
R1049 B.n585 B.n584 10.6151
R1050 B.n585 B.n282 10.6151
R1051 B.n595 B.n282 10.6151
R1052 B.n596 B.n595 10.6151
R1053 B.n597 B.n596 10.6151
R1054 B.n597 B.n275 10.6151
R1055 B.n608 B.n275 10.6151
R1056 B.n609 B.n608 10.6151
R1057 B.n611 B.n609 10.6151
R1058 B.n611 B.n610 10.6151
R1059 B.n610 B.n267 10.6151
R1060 B.n622 B.n267 10.6151
R1061 B.n623 B.n622 10.6151
R1062 B.n624 B.n623 10.6151
R1063 B.n625 B.n624 10.6151
R1064 B.n627 B.n625 10.6151
R1065 B.n628 B.n627 10.6151
R1066 B.n629 B.n628 10.6151
R1067 B.n630 B.n629 10.6151
R1068 B.n632 B.n630 10.6151
R1069 B.n633 B.n632 10.6151
R1070 B.n634 B.n633 10.6151
R1071 B.n635 B.n634 10.6151
R1072 B.n637 B.n635 10.6151
R1073 B.n638 B.n637 10.6151
R1074 B.n639 B.n638 10.6151
R1075 B.n640 B.n639 10.6151
R1076 B.n642 B.n640 10.6151
R1077 B.n643 B.n642 10.6151
R1078 B.n644 B.n643 10.6151
R1079 B.n645 B.n644 10.6151
R1080 B.n647 B.n645 10.6151
R1081 B.n648 B.n647 10.6151
R1082 B.n649 B.n648 10.6151
R1083 B.n650 B.n649 10.6151
R1084 B.n652 B.n650 10.6151
R1085 B.n653 B.n652 10.6151
R1086 B.n654 B.n653 10.6151
R1087 B.n655 B.n654 10.6151
R1088 B.n657 B.n655 10.6151
R1089 B.n658 B.n657 10.6151
R1090 B.n659 B.n658 10.6151
R1091 B.n529 B.n528 10.6151
R1092 B.n528 B.n527 10.6151
R1093 B.n527 B.n526 10.6151
R1094 B.n526 B.n524 10.6151
R1095 B.n524 B.n521 10.6151
R1096 B.n521 B.n520 10.6151
R1097 B.n520 B.n517 10.6151
R1098 B.n517 B.n516 10.6151
R1099 B.n516 B.n513 10.6151
R1100 B.n513 B.n512 10.6151
R1101 B.n512 B.n509 10.6151
R1102 B.n509 B.n508 10.6151
R1103 B.n508 B.n505 10.6151
R1104 B.n505 B.n504 10.6151
R1105 B.n504 B.n501 10.6151
R1106 B.n501 B.n500 10.6151
R1107 B.n500 B.n497 10.6151
R1108 B.n497 B.n496 10.6151
R1109 B.n496 B.n493 10.6151
R1110 B.n493 B.n492 10.6151
R1111 B.n492 B.n489 10.6151
R1112 B.n489 B.n488 10.6151
R1113 B.n488 B.n485 10.6151
R1114 B.n485 B.n484 10.6151
R1115 B.n484 B.n481 10.6151
R1116 B.n481 B.n480 10.6151
R1117 B.n480 B.n477 10.6151
R1118 B.n477 B.n476 10.6151
R1119 B.n476 B.n473 10.6151
R1120 B.n473 B.n472 10.6151
R1121 B.n472 B.n469 10.6151
R1122 B.n469 B.n468 10.6151
R1123 B.n468 B.n465 10.6151
R1124 B.n465 B.n464 10.6151
R1125 B.n464 B.n461 10.6151
R1126 B.n461 B.n460 10.6151
R1127 B.n457 B.n456 10.6151
R1128 B.n456 B.n453 10.6151
R1129 B.n453 B.n452 10.6151
R1130 B.n452 B.n449 10.6151
R1131 B.n449 B.n448 10.6151
R1132 B.n448 B.n445 10.6151
R1133 B.n445 B.n444 10.6151
R1134 B.n444 B.n441 10.6151
R1135 B.n439 B.n436 10.6151
R1136 B.n436 B.n435 10.6151
R1137 B.n435 B.n432 10.6151
R1138 B.n432 B.n431 10.6151
R1139 B.n431 B.n428 10.6151
R1140 B.n428 B.n427 10.6151
R1141 B.n427 B.n424 10.6151
R1142 B.n424 B.n423 10.6151
R1143 B.n423 B.n420 10.6151
R1144 B.n420 B.n419 10.6151
R1145 B.n419 B.n416 10.6151
R1146 B.n416 B.n415 10.6151
R1147 B.n415 B.n412 10.6151
R1148 B.n412 B.n411 10.6151
R1149 B.n411 B.n408 10.6151
R1150 B.n408 B.n407 10.6151
R1151 B.n407 B.n404 10.6151
R1152 B.n404 B.n403 10.6151
R1153 B.n403 B.n400 10.6151
R1154 B.n400 B.n399 10.6151
R1155 B.n399 B.n396 10.6151
R1156 B.n396 B.n395 10.6151
R1157 B.n395 B.n392 10.6151
R1158 B.n392 B.n391 10.6151
R1159 B.n391 B.n388 10.6151
R1160 B.n388 B.n387 10.6151
R1161 B.n387 B.n384 10.6151
R1162 B.n384 B.n383 10.6151
R1163 B.n383 B.n380 10.6151
R1164 B.n380 B.n379 10.6151
R1165 B.n379 B.n376 10.6151
R1166 B.n376 B.n375 10.6151
R1167 B.n375 B.n372 10.6151
R1168 B.n372 B.n371 10.6151
R1169 B.n371 B.n322 10.6151
R1170 B.n535 B.n322 10.6151
R1171 B.n541 B.n318 10.6151
R1172 B.n542 B.n541 10.6151
R1173 B.n543 B.n542 10.6151
R1174 B.n543 B.n310 10.6151
R1175 B.n553 B.n310 10.6151
R1176 B.n554 B.n553 10.6151
R1177 B.n555 B.n554 10.6151
R1178 B.n555 B.n302 10.6151
R1179 B.n565 B.n302 10.6151
R1180 B.n566 B.n565 10.6151
R1181 B.n567 B.n566 10.6151
R1182 B.n567 B.n294 10.6151
R1183 B.n577 B.n294 10.6151
R1184 B.n578 B.n577 10.6151
R1185 B.n579 B.n578 10.6151
R1186 B.n579 B.n286 10.6151
R1187 B.n589 B.n286 10.6151
R1188 B.n590 B.n589 10.6151
R1189 B.n591 B.n590 10.6151
R1190 B.n591 B.n278 10.6151
R1191 B.n602 B.n278 10.6151
R1192 B.n603 B.n602 10.6151
R1193 B.n604 B.n603 10.6151
R1194 B.n604 B.n271 10.6151
R1195 B.n615 B.n271 10.6151
R1196 B.n616 B.n615 10.6151
R1197 B.n617 B.n616 10.6151
R1198 B.n617 B.n0 10.6151
R1199 B.n716 B.n1 10.6151
R1200 B.n716 B.n715 10.6151
R1201 B.n715 B.n714 10.6151
R1202 B.n714 B.n10 10.6151
R1203 B.n708 B.n10 10.6151
R1204 B.n708 B.n707 10.6151
R1205 B.n707 B.n706 10.6151
R1206 B.n706 B.n16 10.6151
R1207 B.n700 B.n16 10.6151
R1208 B.n700 B.n699 10.6151
R1209 B.n699 B.n698 10.6151
R1210 B.n698 B.n24 10.6151
R1211 B.n692 B.n24 10.6151
R1212 B.n692 B.n691 10.6151
R1213 B.n691 B.n690 10.6151
R1214 B.n690 B.n31 10.6151
R1215 B.n684 B.n31 10.6151
R1216 B.n684 B.n683 10.6151
R1217 B.n683 B.n682 10.6151
R1218 B.n682 B.n38 10.6151
R1219 B.n676 B.n38 10.6151
R1220 B.n676 B.n675 10.6151
R1221 B.n675 B.n674 10.6151
R1222 B.n674 B.n45 10.6151
R1223 B.n668 B.n45 10.6151
R1224 B.n668 B.n667 10.6151
R1225 B.n667 B.n666 10.6151
R1226 B.n666 B.n52 10.6151
R1227 B.n178 B.n177 6.5566
R1228 B.n194 B.n100 6.5566
R1229 B.n457 B.n367 6.5566
R1230 B.n441 B.n440 6.5566
R1231 B.n599 B.t1 6.3365
R1232 B.n18 B.t0 6.3365
R1233 B.n177 B.n176 4.05904
R1234 B.n197 B.n100 4.05904
R1235 B.n460 B.n367 4.05904
R1236 B.n440 B.n439 4.05904
R1237 B.n722 B.n0 2.81026
R1238 B.n722 B.n1 2.81026
R1239 VP.n0 VP.t0 160.667
R1240 VP.n0 VP.t1 115.537
R1241 VP VP.n0 0.52637
R1242 VDD1 VDD1.t0 105.028
R1243 VDD1 VDD1.t1 65.8074
C0 VDD1 VDD2 0.753636f
C1 VDD1 VTAIL 4.76381f
C2 VDD1 VN 0.148421f
C3 VP VDD2 0.360261f
C4 VP VTAIL 2.30871f
C5 VN VP 5.45791f
C6 VDD1 VP 2.71771f
C7 VDD2 VTAIL 4.81968f
C8 VN VDD2 2.50788f
C9 VN VTAIL 2.29448f
C10 VDD2 B 4.36167f
C11 VDD1 B 7.51854f
C12 VTAIL B 7.001776f
C13 VN B 11.0137f
C14 VP B 7.106787f
C15 VDD1.t1 B 1.91673f
C16 VDD1.t0 B 2.4909f
C17 VP.t0 B 3.60408f
C18 VP.t1 B 2.96556f
C19 VP.n0 B 3.83283f
C20 VDD2.t1 B 2.41014f
C21 VDD2.t0 B 1.88138f
C22 VDD2.n0 B 2.85151f
C23 VTAIL.t1 B 1.90012f
C24 VTAIL.n0 B 1.70739f
C25 VTAIL.t3 B 1.90012f
C26 VTAIL.n1 B 1.75682f
C27 VTAIL.t0 B 1.90012f
C28 VTAIL.n2 B 1.54294f
C29 VTAIL.t2 B 1.90012f
C30 VTAIL.n3 B 1.45287f
C31 VN.t0 B 2.90222f
C32 VN.t1 B 3.5222f
.ends

