* NGSPICE file created from diff_pair_sample_0349.ext - technology: sky130A

.subckt diff_pair_sample_0349 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1802_n1278# sky130_fd_pr__pfet_01v8 ad=0.6045 pd=3.88 as=0 ps=0 w=1.55 l=1.75
X1 VDD1.t1 VP.t0 VTAIL.t3 w_n1802_n1278# sky130_fd_pr__pfet_01v8 ad=0.6045 pd=3.88 as=0.6045 ps=3.88 w=1.55 l=1.75
X2 VDD2.t1 VN.t0 VTAIL.t1 w_n1802_n1278# sky130_fd_pr__pfet_01v8 ad=0.6045 pd=3.88 as=0.6045 ps=3.88 w=1.55 l=1.75
X3 VDD2.t0 VN.t1 VTAIL.t0 w_n1802_n1278# sky130_fd_pr__pfet_01v8 ad=0.6045 pd=3.88 as=0.6045 ps=3.88 w=1.55 l=1.75
X4 B.t8 B.t6 B.t7 w_n1802_n1278# sky130_fd_pr__pfet_01v8 ad=0.6045 pd=3.88 as=0 ps=0 w=1.55 l=1.75
X5 VDD1.t0 VP.t1 VTAIL.t2 w_n1802_n1278# sky130_fd_pr__pfet_01v8 ad=0.6045 pd=3.88 as=0.6045 ps=3.88 w=1.55 l=1.75
X6 B.t5 B.t3 B.t4 w_n1802_n1278# sky130_fd_pr__pfet_01v8 ad=0.6045 pd=3.88 as=0 ps=0 w=1.55 l=1.75
X7 B.t2 B.t0 B.t1 w_n1802_n1278# sky130_fd_pr__pfet_01v8 ad=0.6045 pd=3.88 as=0 ps=0 w=1.55 l=1.75
R0 B.n158 B.n53 585
R1 B.n157 B.n156 585
R2 B.n155 B.n54 585
R3 B.n154 B.n153 585
R4 B.n152 B.n55 585
R5 B.n151 B.n150 585
R6 B.n149 B.n56 585
R7 B.n148 B.n147 585
R8 B.n146 B.n57 585
R9 B.n145 B.n144 585
R10 B.n143 B.n58 585
R11 B.n142 B.n141 585
R12 B.n137 B.n59 585
R13 B.n136 B.n135 585
R14 B.n134 B.n60 585
R15 B.n133 B.n132 585
R16 B.n131 B.n61 585
R17 B.n130 B.n129 585
R18 B.n128 B.n62 585
R19 B.n127 B.n126 585
R20 B.n124 B.n63 585
R21 B.n123 B.n122 585
R22 B.n121 B.n66 585
R23 B.n120 B.n119 585
R24 B.n118 B.n67 585
R25 B.n117 B.n116 585
R26 B.n115 B.n68 585
R27 B.n114 B.n113 585
R28 B.n112 B.n69 585
R29 B.n111 B.n110 585
R30 B.n109 B.n70 585
R31 B.n160 B.n159 585
R32 B.n161 B.n52 585
R33 B.n163 B.n162 585
R34 B.n164 B.n51 585
R35 B.n166 B.n165 585
R36 B.n167 B.n50 585
R37 B.n169 B.n168 585
R38 B.n170 B.n49 585
R39 B.n172 B.n171 585
R40 B.n173 B.n48 585
R41 B.n175 B.n174 585
R42 B.n176 B.n47 585
R43 B.n178 B.n177 585
R44 B.n179 B.n46 585
R45 B.n181 B.n180 585
R46 B.n182 B.n45 585
R47 B.n184 B.n183 585
R48 B.n185 B.n44 585
R49 B.n187 B.n186 585
R50 B.n188 B.n43 585
R51 B.n190 B.n189 585
R52 B.n191 B.n42 585
R53 B.n193 B.n192 585
R54 B.n194 B.n41 585
R55 B.n196 B.n195 585
R56 B.n197 B.n40 585
R57 B.n199 B.n198 585
R58 B.n200 B.n39 585
R59 B.n202 B.n201 585
R60 B.n203 B.n38 585
R61 B.n205 B.n204 585
R62 B.n206 B.n37 585
R63 B.n208 B.n207 585
R64 B.n209 B.n36 585
R65 B.n211 B.n210 585
R66 B.n212 B.n35 585
R67 B.n214 B.n213 585
R68 B.n215 B.n34 585
R69 B.n217 B.n216 585
R70 B.n218 B.n33 585
R71 B.n220 B.n219 585
R72 B.n221 B.n32 585
R73 B.n269 B.n12 585
R74 B.n268 B.n267 585
R75 B.n266 B.n13 585
R76 B.n265 B.n264 585
R77 B.n263 B.n14 585
R78 B.n262 B.n261 585
R79 B.n260 B.n15 585
R80 B.n259 B.n258 585
R81 B.n257 B.n16 585
R82 B.n256 B.n255 585
R83 B.n254 B.n17 585
R84 B.n252 B.n251 585
R85 B.n250 B.n20 585
R86 B.n249 B.n248 585
R87 B.n247 B.n21 585
R88 B.n246 B.n245 585
R89 B.n244 B.n22 585
R90 B.n243 B.n242 585
R91 B.n241 B.n23 585
R92 B.n240 B.n239 585
R93 B.n238 B.n237 585
R94 B.n236 B.n27 585
R95 B.n235 B.n234 585
R96 B.n233 B.n28 585
R97 B.n232 B.n231 585
R98 B.n230 B.n29 585
R99 B.n229 B.n228 585
R100 B.n227 B.n30 585
R101 B.n226 B.n225 585
R102 B.n224 B.n31 585
R103 B.n223 B.n222 585
R104 B.n271 B.n270 585
R105 B.n272 B.n11 585
R106 B.n274 B.n273 585
R107 B.n275 B.n10 585
R108 B.n277 B.n276 585
R109 B.n278 B.n9 585
R110 B.n280 B.n279 585
R111 B.n281 B.n8 585
R112 B.n283 B.n282 585
R113 B.n284 B.n7 585
R114 B.n286 B.n285 585
R115 B.n287 B.n6 585
R116 B.n289 B.n288 585
R117 B.n290 B.n5 585
R118 B.n292 B.n291 585
R119 B.n293 B.n4 585
R120 B.n295 B.n294 585
R121 B.n296 B.n3 585
R122 B.n298 B.n297 585
R123 B.n299 B.n0 585
R124 B.n2 B.n1 585
R125 B.n81 B.n80 585
R126 B.n82 B.n79 585
R127 B.n84 B.n83 585
R128 B.n85 B.n78 585
R129 B.n87 B.n86 585
R130 B.n88 B.n77 585
R131 B.n90 B.n89 585
R132 B.n91 B.n76 585
R133 B.n93 B.n92 585
R134 B.n94 B.n75 585
R135 B.n96 B.n95 585
R136 B.n97 B.n74 585
R137 B.n99 B.n98 585
R138 B.n100 B.n73 585
R139 B.n102 B.n101 585
R140 B.n103 B.n72 585
R141 B.n105 B.n104 585
R142 B.n106 B.n71 585
R143 B.n108 B.n107 585
R144 B.n109 B.n108 502.111
R145 B.n160 B.n53 502.111
R146 B.n222 B.n221 502.111
R147 B.n270 B.n269 502.111
R148 B.n138 B.t1 290.058
R149 B.n24 B.t11 290.058
R150 B.n64 B.t7 290.058
R151 B.n18 B.t5 290.058
R152 B.n301 B.n300 256.663
R153 B.n139 B.t2 249.719
R154 B.n25 B.t10 249.719
R155 B.n65 B.t8 249.718
R156 B.n19 B.t4 249.718
R157 B.n300 B.n299 235.042
R158 B.n300 B.n2 235.042
R159 B.n64 B.t6 227.609
R160 B.n138 B.t0 227.609
R161 B.n24 B.t9 227.609
R162 B.n18 B.t3 227.609
R163 B.n110 B.n109 163.367
R164 B.n110 B.n69 163.367
R165 B.n114 B.n69 163.367
R166 B.n115 B.n114 163.367
R167 B.n116 B.n115 163.367
R168 B.n116 B.n67 163.367
R169 B.n120 B.n67 163.367
R170 B.n121 B.n120 163.367
R171 B.n122 B.n121 163.367
R172 B.n122 B.n63 163.367
R173 B.n127 B.n63 163.367
R174 B.n128 B.n127 163.367
R175 B.n129 B.n128 163.367
R176 B.n129 B.n61 163.367
R177 B.n133 B.n61 163.367
R178 B.n134 B.n133 163.367
R179 B.n135 B.n134 163.367
R180 B.n135 B.n59 163.367
R181 B.n142 B.n59 163.367
R182 B.n143 B.n142 163.367
R183 B.n144 B.n143 163.367
R184 B.n144 B.n57 163.367
R185 B.n148 B.n57 163.367
R186 B.n149 B.n148 163.367
R187 B.n150 B.n149 163.367
R188 B.n150 B.n55 163.367
R189 B.n154 B.n55 163.367
R190 B.n155 B.n154 163.367
R191 B.n156 B.n155 163.367
R192 B.n156 B.n53 163.367
R193 B.n221 B.n220 163.367
R194 B.n220 B.n33 163.367
R195 B.n216 B.n33 163.367
R196 B.n216 B.n215 163.367
R197 B.n215 B.n214 163.367
R198 B.n214 B.n35 163.367
R199 B.n210 B.n35 163.367
R200 B.n210 B.n209 163.367
R201 B.n209 B.n208 163.367
R202 B.n208 B.n37 163.367
R203 B.n204 B.n37 163.367
R204 B.n204 B.n203 163.367
R205 B.n203 B.n202 163.367
R206 B.n202 B.n39 163.367
R207 B.n198 B.n39 163.367
R208 B.n198 B.n197 163.367
R209 B.n197 B.n196 163.367
R210 B.n196 B.n41 163.367
R211 B.n192 B.n41 163.367
R212 B.n192 B.n191 163.367
R213 B.n191 B.n190 163.367
R214 B.n190 B.n43 163.367
R215 B.n186 B.n43 163.367
R216 B.n186 B.n185 163.367
R217 B.n185 B.n184 163.367
R218 B.n184 B.n45 163.367
R219 B.n180 B.n45 163.367
R220 B.n180 B.n179 163.367
R221 B.n179 B.n178 163.367
R222 B.n178 B.n47 163.367
R223 B.n174 B.n47 163.367
R224 B.n174 B.n173 163.367
R225 B.n173 B.n172 163.367
R226 B.n172 B.n49 163.367
R227 B.n168 B.n49 163.367
R228 B.n168 B.n167 163.367
R229 B.n167 B.n166 163.367
R230 B.n166 B.n51 163.367
R231 B.n162 B.n51 163.367
R232 B.n162 B.n161 163.367
R233 B.n161 B.n160 163.367
R234 B.n269 B.n268 163.367
R235 B.n268 B.n13 163.367
R236 B.n264 B.n13 163.367
R237 B.n264 B.n263 163.367
R238 B.n263 B.n262 163.367
R239 B.n262 B.n15 163.367
R240 B.n258 B.n15 163.367
R241 B.n258 B.n257 163.367
R242 B.n257 B.n256 163.367
R243 B.n256 B.n17 163.367
R244 B.n251 B.n17 163.367
R245 B.n251 B.n250 163.367
R246 B.n250 B.n249 163.367
R247 B.n249 B.n21 163.367
R248 B.n245 B.n21 163.367
R249 B.n245 B.n244 163.367
R250 B.n244 B.n243 163.367
R251 B.n243 B.n23 163.367
R252 B.n239 B.n23 163.367
R253 B.n239 B.n238 163.367
R254 B.n238 B.n27 163.367
R255 B.n234 B.n27 163.367
R256 B.n234 B.n233 163.367
R257 B.n233 B.n232 163.367
R258 B.n232 B.n29 163.367
R259 B.n228 B.n29 163.367
R260 B.n228 B.n227 163.367
R261 B.n227 B.n226 163.367
R262 B.n226 B.n31 163.367
R263 B.n222 B.n31 163.367
R264 B.n270 B.n11 163.367
R265 B.n274 B.n11 163.367
R266 B.n275 B.n274 163.367
R267 B.n276 B.n275 163.367
R268 B.n276 B.n9 163.367
R269 B.n280 B.n9 163.367
R270 B.n281 B.n280 163.367
R271 B.n282 B.n281 163.367
R272 B.n282 B.n7 163.367
R273 B.n286 B.n7 163.367
R274 B.n287 B.n286 163.367
R275 B.n288 B.n287 163.367
R276 B.n288 B.n5 163.367
R277 B.n292 B.n5 163.367
R278 B.n293 B.n292 163.367
R279 B.n294 B.n293 163.367
R280 B.n294 B.n3 163.367
R281 B.n298 B.n3 163.367
R282 B.n299 B.n298 163.367
R283 B.n80 B.n2 163.367
R284 B.n80 B.n79 163.367
R285 B.n84 B.n79 163.367
R286 B.n85 B.n84 163.367
R287 B.n86 B.n85 163.367
R288 B.n86 B.n77 163.367
R289 B.n90 B.n77 163.367
R290 B.n91 B.n90 163.367
R291 B.n92 B.n91 163.367
R292 B.n92 B.n75 163.367
R293 B.n96 B.n75 163.367
R294 B.n97 B.n96 163.367
R295 B.n98 B.n97 163.367
R296 B.n98 B.n73 163.367
R297 B.n102 B.n73 163.367
R298 B.n103 B.n102 163.367
R299 B.n104 B.n103 163.367
R300 B.n104 B.n71 163.367
R301 B.n108 B.n71 163.367
R302 B.n125 B.n65 59.5399
R303 B.n140 B.n139 59.5399
R304 B.n26 B.n25 59.5399
R305 B.n253 B.n19 59.5399
R306 B.n65 B.n64 40.3399
R307 B.n139 B.n138 40.3399
R308 B.n25 B.n24 40.3399
R309 B.n19 B.n18 40.3399
R310 B.n271 B.n12 32.6249
R311 B.n223 B.n32 32.6249
R312 B.n159 B.n158 32.6249
R313 B.n107 B.n70 32.6249
R314 B B.n301 18.0485
R315 B.n272 B.n271 10.6151
R316 B.n273 B.n272 10.6151
R317 B.n273 B.n10 10.6151
R318 B.n277 B.n10 10.6151
R319 B.n278 B.n277 10.6151
R320 B.n279 B.n278 10.6151
R321 B.n279 B.n8 10.6151
R322 B.n283 B.n8 10.6151
R323 B.n284 B.n283 10.6151
R324 B.n285 B.n284 10.6151
R325 B.n285 B.n6 10.6151
R326 B.n289 B.n6 10.6151
R327 B.n290 B.n289 10.6151
R328 B.n291 B.n290 10.6151
R329 B.n291 B.n4 10.6151
R330 B.n295 B.n4 10.6151
R331 B.n296 B.n295 10.6151
R332 B.n297 B.n296 10.6151
R333 B.n297 B.n0 10.6151
R334 B.n267 B.n12 10.6151
R335 B.n267 B.n266 10.6151
R336 B.n266 B.n265 10.6151
R337 B.n265 B.n14 10.6151
R338 B.n261 B.n14 10.6151
R339 B.n261 B.n260 10.6151
R340 B.n260 B.n259 10.6151
R341 B.n259 B.n16 10.6151
R342 B.n255 B.n16 10.6151
R343 B.n255 B.n254 10.6151
R344 B.n252 B.n20 10.6151
R345 B.n248 B.n20 10.6151
R346 B.n248 B.n247 10.6151
R347 B.n247 B.n246 10.6151
R348 B.n246 B.n22 10.6151
R349 B.n242 B.n22 10.6151
R350 B.n242 B.n241 10.6151
R351 B.n241 B.n240 10.6151
R352 B.n237 B.n236 10.6151
R353 B.n236 B.n235 10.6151
R354 B.n235 B.n28 10.6151
R355 B.n231 B.n28 10.6151
R356 B.n231 B.n230 10.6151
R357 B.n230 B.n229 10.6151
R358 B.n229 B.n30 10.6151
R359 B.n225 B.n30 10.6151
R360 B.n225 B.n224 10.6151
R361 B.n224 B.n223 10.6151
R362 B.n219 B.n32 10.6151
R363 B.n219 B.n218 10.6151
R364 B.n218 B.n217 10.6151
R365 B.n217 B.n34 10.6151
R366 B.n213 B.n34 10.6151
R367 B.n213 B.n212 10.6151
R368 B.n212 B.n211 10.6151
R369 B.n211 B.n36 10.6151
R370 B.n207 B.n36 10.6151
R371 B.n207 B.n206 10.6151
R372 B.n206 B.n205 10.6151
R373 B.n205 B.n38 10.6151
R374 B.n201 B.n38 10.6151
R375 B.n201 B.n200 10.6151
R376 B.n200 B.n199 10.6151
R377 B.n199 B.n40 10.6151
R378 B.n195 B.n40 10.6151
R379 B.n195 B.n194 10.6151
R380 B.n194 B.n193 10.6151
R381 B.n193 B.n42 10.6151
R382 B.n189 B.n42 10.6151
R383 B.n189 B.n188 10.6151
R384 B.n188 B.n187 10.6151
R385 B.n187 B.n44 10.6151
R386 B.n183 B.n44 10.6151
R387 B.n183 B.n182 10.6151
R388 B.n182 B.n181 10.6151
R389 B.n181 B.n46 10.6151
R390 B.n177 B.n46 10.6151
R391 B.n177 B.n176 10.6151
R392 B.n176 B.n175 10.6151
R393 B.n175 B.n48 10.6151
R394 B.n171 B.n48 10.6151
R395 B.n171 B.n170 10.6151
R396 B.n170 B.n169 10.6151
R397 B.n169 B.n50 10.6151
R398 B.n165 B.n50 10.6151
R399 B.n165 B.n164 10.6151
R400 B.n164 B.n163 10.6151
R401 B.n163 B.n52 10.6151
R402 B.n159 B.n52 10.6151
R403 B.n81 B.n1 10.6151
R404 B.n82 B.n81 10.6151
R405 B.n83 B.n82 10.6151
R406 B.n83 B.n78 10.6151
R407 B.n87 B.n78 10.6151
R408 B.n88 B.n87 10.6151
R409 B.n89 B.n88 10.6151
R410 B.n89 B.n76 10.6151
R411 B.n93 B.n76 10.6151
R412 B.n94 B.n93 10.6151
R413 B.n95 B.n94 10.6151
R414 B.n95 B.n74 10.6151
R415 B.n99 B.n74 10.6151
R416 B.n100 B.n99 10.6151
R417 B.n101 B.n100 10.6151
R418 B.n101 B.n72 10.6151
R419 B.n105 B.n72 10.6151
R420 B.n106 B.n105 10.6151
R421 B.n107 B.n106 10.6151
R422 B.n111 B.n70 10.6151
R423 B.n112 B.n111 10.6151
R424 B.n113 B.n112 10.6151
R425 B.n113 B.n68 10.6151
R426 B.n117 B.n68 10.6151
R427 B.n118 B.n117 10.6151
R428 B.n119 B.n118 10.6151
R429 B.n119 B.n66 10.6151
R430 B.n123 B.n66 10.6151
R431 B.n124 B.n123 10.6151
R432 B.n126 B.n62 10.6151
R433 B.n130 B.n62 10.6151
R434 B.n131 B.n130 10.6151
R435 B.n132 B.n131 10.6151
R436 B.n132 B.n60 10.6151
R437 B.n136 B.n60 10.6151
R438 B.n137 B.n136 10.6151
R439 B.n141 B.n137 10.6151
R440 B.n145 B.n58 10.6151
R441 B.n146 B.n145 10.6151
R442 B.n147 B.n146 10.6151
R443 B.n147 B.n56 10.6151
R444 B.n151 B.n56 10.6151
R445 B.n152 B.n151 10.6151
R446 B.n153 B.n152 10.6151
R447 B.n153 B.n54 10.6151
R448 B.n157 B.n54 10.6151
R449 B.n158 B.n157 10.6151
R450 B.n301 B.n0 8.11757
R451 B.n301 B.n1 8.11757
R452 B.n253 B.n252 6.5566
R453 B.n240 B.n26 6.5566
R454 B.n126 B.n125 6.5566
R455 B.n141 B.n140 6.5566
R456 B.n254 B.n253 4.05904
R457 B.n237 B.n26 4.05904
R458 B.n125 B.n124 4.05904
R459 B.n140 B.n58 4.05904
R460 VP.n0 VP.t0 114.692
R461 VP.n0 VP.t1 80.207
R462 VP VP.n0 0.241678
R463 VTAIL.n1 VTAIL.t1 256.214
R464 VTAIL.n3 VTAIL.t0 256.214
R465 VTAIL.n0 VTAIL.t2 256.214
R466 VTAIL.n2 VTAIL.t3 256.214
R467 VTAIL.n1 VTAIL.n0 17.2893
R468 VTAIL.n3 VTAIL.n2 15.4962
R469 VTAIL.n2 VTAIL.n1 1.36688
R470 VTAIL VTAIL.n0 0.976793
R471 VTAIL VTAIL.n3 0.390586
R472 VDD1 VDD1.t0 302.447
R473 VDD1 VDD1.t1 273.399
R474 VN VN.t0 114.883
R475 VN VN.t1 80.4481
R476 VDD2.n0 VDD2.t0 301.474
R477 VDD2.n0 VDD2.t1 272.892
R478 VDD2 VDD2.n0 0.506965
C0 VDD2 w_n1802_n1278# 0.952832f
C1 VTAIL VP 0.782953f
C2 VTAIL VN 0.768811f
C3 VDD2 B 0.802576f
C4 w_n1802_n1278# VTAIL 1.17031f
C5 VDD1 VP 0.700015f
C6 VDD1 VN 0.154722f
C7 w_n1802_n1278# VDD1 0.938021f
C8 B VTAIL 1.01613f
C9 B VDD1 0.779673f
C10 VP VN 3.13135f
C11 VDD2 VTAIL 2.08291f
C12 w_n1802_n1278# VP 2.40742f
C13 w_n1802_n1278# VN 2.18574f
C14 VDD2 VDD1 0.572758f
C15 B VP 1.11735f
C16 B VN 0.747343f
C17 VTAIL VDD1 2.03575f
C18 w_n1802_n1278# B 4.97088f
C19 VDD2 VP 0.304208f
C20 VDD2 VN 0.552106f
C21 VDD2 VSUBS 0.465439f
C22 VDD1 VSUBS 2.286301f
C23 VTAIL VSUBS 0.312811f
C24 VN VSUBS 4.92818f
C25 VP VSUBS 0.95503f
C26 B VSUBS 2.258035f
C27 w_n1802_n1278# VSUBS 29.516802f
C28 VDD2.t0 VSUBS 0.202324f
C29 VDD2.t1 VSUBS 0.132647f
C30 VDD2.n0 VSUBS 1.68473f
C31 VN.t1 VSUBS 0.69019f
C32 VN.t0 VSUBS 1.26876f
C33 VDD1.t1 VSUBS 0.122891f
C34 VDD1.t0 VSUBS 0.193296f
C35 VTAIL.t2 VSUBS 0.149465f
C36 VTAIL.n0 VSUBS 0.91102f
C37 VTAIL.t1 VSUBS 0.149465f
C38 VTAIL.n1 VSUBS 0.938351f
C39 VTAIL.t3 VSUBS 0.149465f
C40 VTAIL.n2 VSUBS 0.812719f
C41 VTAIL.t0 VSUBS 0.149465f
C42 VTAIL.n3 VSUBS 0.744316f
C43 VP.t0 VSUBS 1.32546f
C44 VP.t1 VSUBS 0.726334f
C45 VP.n0 VSUBS 3.35966f
C46 B.n0 VSUBS 0.008811f
C47 B.n1 VSUBS 0.008811f
C48 B.n2 VSUBS 0.01303f
C49 B.n3 VSUBS 0.009985f
C50 B.n4 VSUBS 0.009985f
C51 B.n5 VSUBS 0.009985f
C52 B.n6 VSUBS 0.009985f
C53 B.n7 VSUBS 0.009985f
C54 B.n8 VSUBS 0.009985f
C55 B.n9 VSUBS 0.009985f
C56 B.n10 VSUBS 0.009985f
C57 B.n11 VSUBS 0.009985f
C58 B.n12 VSUBS 0.023593f
C59 B.n13 VSUBS 0.009985f
C60 B.n14 VSUBS 0.009985f
C61 B.n15 VSUBS 0.009985f
C62 B.n16 VSUBS 0.009985f
C63 B.n17 VSUBS 0.009985f
C64 B.t4 VSUBS 0.045116f
C65 B.t5 VSUBS 0.053032f
C66 B.t3 VSUBS 0.191536f
C67 B.n18 VSUBS 0.084154f
C68 B.n19 VSUBS 0.071167f
C69 B.n20 VSUBS 0.009985f
C70 B.n21 VSUBS 0.009985f
C71 B.n22 VSUBS 0.009985f
C72 B.n23 VSUBS 0.009985f
C73 B.t10 VSUBS 0.045116f
C74 B.t11 VSUBS 0.053032f
C75 B.t9 VSUBS 0.191536f
C76 B.n24 VSUBS 0.084154f
C77 B.n25 VSUBS 0.071167f
C78 B.n26 VSUBS 0.023135f
C79 B.n27 VSUBS 0.009985f
C80 B.n28 VSUBS 0.009985f
C81 B.n29 VSUBS 0.009985f
C82 B.n30 VSUBS 0.009985f
C83 B.n31 VSUBS 0.009985f
C84 B.n32 VSUBS 0.023103f
C85 B.n33 VSUBS 0.009985f
C86 B.n34 VSUBS 0.009985f
C87 B.n35 VSUBS 0.009985f
C88 B.n36 VSUBS 0.009985f
C89 B.n37 VSUBS 0.009985f
C90 B.n38 VSUBS 0.009985f
C91 B.n39 VSUBS 0.009985f
C92 B.n40 VSUBS 0.009985f
C93 B.n41 VSUBS 0.009985f
C94 B.n42 VSUBS 0.009985f
C95 B.n43 VSUBS 0.009985f
C96 B.n44 VSUBS 0.009985f
C97 B.n45 VSUBS 0.009985f
C98 B.n46 VSUBS 0.009985f
C99 B.n47 VSUBS 0.009985f
C100 B.n48 VSUBS 0.009985f
C101 B.n49 VSUBS 0.009985f
C102 B.n50 VSUBS 0.009985f
C103 B.n51 VSUBS 0.009985f
C104 B.n52 VSUBS 0.009985f
C105 B.n53 VSUBS 0.023593f
C106 B.n54 VSUBS 0.009985f
C107 B.n55 VSUBS 0.009985f
C108 B.n56 VSUBS 0.009985f
C109 B.n57 VSUBS 0.009985f
C110 B.n58 VSUBS 0.006902f
C111 B.n59 VSUBS 0.009985f
C112 B.n60 VSUBS 0.009985f
C113 B.n61 VSUBS 0.009985f
C114 B.n62 VSUBS 0.009985f
C115 B.n63 VSUBS 0.009985f
C116 B.t8 VSUBS 0.045116f
C117 B.t7 VSUBS 0.053032f
C118 B.t6 VSUBS 0.191536f
C119 B.n64 VSUBS 0.084154f
C120 B.n65 VSUBS 0.071167f
C121 B.n66 VSUBS 0.009985f
C122 B.n67 VSUBS 0.009985f
C123 B.n68 VSUBS 0.009985f
C124 B.n69 VSUBS 0.009985f
C125 B.n70 VSUBS 0.023593f
C126 B.n71 VSUBS 0.009985f
C127 B.n72 VSUBS 0.009985f
C128 B.n73 VSUBS 0.009985f
C129 B.n74 VSUBS 0.009985f
C130 B.n75 VSUBS 0.009985f
C131 B.n76 VSUBS 0.009985f
C132 B.n77 VSUBS 0.009985f
C133 B.n78 VSUBS 0.009985f
C134 B.n79 VSUBS 0.009985f
C135 B.n80 VSUBS 0.009985f
C136 B.n81 VSUBS 0.009985f
C137 B.n82 VSUBS 0.009985f
C138 B.n83 VSUBS 0.009985f
C139 B.n84 VSUBS 0.009985f
C140 B.n85 VSUBS 0.009985f
C141 B.n86 VSUBS 0.009985f
C142 B.n87 VSUBS 0.009985f
C143 B.n88 VSUBS 0.009985f
C144 B.n89 VSUBS 0.009985f
C145 B.n90 VSUBS 0.009985f
C146 B.n91 VSUBS 0.009985f
C147 B.n92 VSUBS 0.009985f
C148 B.n93 VSUBS 0.009985f
C149 B.n94 VSUBS 0.009985f
C150 B.n95 VSUBS 0.009985f
C151 B.n96 VSUBS 0.009985f
C152 B.n97 VSUBS 0.009985f
C153 B.n98 VSUBS 0.009985f
C154 B.n99 VSUBS 0.009985f
C155 B.n100 VSUBS 0.009985f
C156 B.n101 VSUBS 0.009985f
C157 B.n102 VSUBS 0.009985f
C158 B.n103 VSUBS 0.009985f
C159 B.n104 VSUBS 0.009985f
C160 B.n105 VSUBS 0.009985f
C161 B.n106 VSUBS 0.009985f
C162 B.n107 VSUBS 0.023103f
C163 B.n108 VSUBS 0.023103f
C164 B.n109 VSUBS 0.023593f
C165 B.n110 VSUBS 0.009985f
C166 B.n111 VSUBS 0.009985f
C167 B.n112 VSUBS 0.009985f
C168 B.n113 VSUBS 0.009985f
C169 B.n114 VSUBS 0.009985f
C170 B.n115 VSUBS 0.009985f
C171 B.n116 VSUBS 0.009985f
C172 B.n117 VSUBS 0.009985f
C173 B.n118 VSUBS 0.009985f
C174 B.n119 VSUBS 0.009985f
C175 B.n120 VSUBS 0.009985f
C176 B.n121 VSUBS 0.009985f
C177 B.n122 VSUBS 0.009985f
C178 B.n123 VSUBS 0.009985f
C179 B.n124 VSUBS 0.006902f
C180 B.n125 VSUBS 0.023135f
C181 B.n126 VSUBS 0.008076f
C182 B.n127 VSUBS 0.009985f
C183 B.n128 VSUBS 0.009985f
C184 B.n129 VSUBS 0.009985f
C185 B.n130 VSUBS 0.009985f
C186 B.n131 VSUBS 0.009985f
C187 B.n132 VSUBS 0.009985f
C188 B.n133 VSUBS 0.009985f
C189 B.n134 VSUBS 0.009985f
C190 B.n135 VSUBS 0.009985f
C191 B.n136 VSUBS 0.009985f
C192 B.n137 VSUBS 0.009985f
C193 B.t2 VSUBS 0.045116f
C194 B.t1 VSUBS 0.053032f
C195 B.t0 VSUBS 0.191536f
C196 B.n138 VSUBS 0.084154f
C197 B.n139 VSUBS 0.071167f
C198 B.n140 VSUBS 0.023135f
C199 B.n141 VSUBS 0.008076f
C200 B.n142 VSUBS 0.009985f
C201 B.n143 VSUBS 0.009985f
C202 B.n144 VSUBS 0.009985f
C203 B.n145 VSUBS 0.009985f
C204 B.n146 VSUBS 0.009985f
C205 B.n147 VSUBS 0.009985f
C206 B.n148 VSUBS 0.009985f
C207 B.n149 VSUBS 0.009985f
C208 B.n150 VSUBS 0.009985f
C209 B.n151 VSUBS 0.009985f
C210 B.n152 VSUBS 0.009985f
C211 B.n153 VSUBS 0.009985f
C212 B.n154 VSUBS 0.009985f
C213 B.n155 VSUBS 0.009985f
C214 B.n156 VSUBS 0.009985f
C215 B.n157 VSUBS 0.009985f
C216 B.n158 VSUBS 0.022412f
C217 B.n159 VSUBS 0.024284f
C218 B.n160 VSUBS 0.023103f
C219 B.n161 VSUBS 0.009985f
C220 B.n162 VSUBS 0.009985f
C221 B.n163 VSUBS 0.009985f
C222 B.n164 VSUBS 0.009985f
C223 B.n165 VSUBS 0.009985f
C224 B.n166 VSUBS 0.009985f
C225 B.n167 VSUBS 0.009985f
C226 B.n168 VSUBS 0.009985f
C227 B.n169 VSUBS 0.009985f
C228 B.n170 VSUBS 0.009985f
C229 B.n171 VSUBS 0.009985f
C230 B.n172 VSUBS 0.009985f
C231 B.n173 VSUBS 0.009985f
C232 B.n174 VSUBS 0.009985f
C233 B.n175 VSUBS 0.009985f
C234 B.n176 VSUBS 0.009985f
C235 B.n177 VSUBS 0.009985f
C236 B.n178 VSUBS 0.009985f
C237 B.n179 VSUBS 0.009985f
C238 B.n180 VSUBS 0.009985f
C239 B.n181 VSUBS 0.009985f
C240 B.n182 VSUBS 0.009985f
C241 B.n183 VSUBS 0.009985f
C242 B.n184 VSUBS 0.009985f
C243 B.n185 VSUBS 0.009985f
C244 B.n186 VSUBS 0.009985f
C245 B.n187 VSUBS 0.009985f
C246 B.n188 VSUBS 0.009985f
C247 B.n189 VSUBS 0.009985f
C248 B.n190 VSUBS 0.009985f
C249 B.n191 VSUBS 0.009985f
C250 B.n192 VSUBS 0.009985f
C251 B.n193 VSUBS 0.009985f
C252 B.n194 VSUBS 0.009985f
C253 B.n195 VSUBS 0.009985f
C254 B.n196 VSUBS 0.009985f
C255 B.n197 VSUBS 0.009985f
C256 B.n198 VSUBS 0.009985f
C257 B.n199 VSUBS 0.009985f
C258 B.n200 VSUBS 0.009985f
C259 B.n201 VSUBS 0.009985f
C260 B.n202 VSUBS 0.009985f
C261 B.n203 VSUBS 0.009985f
C262 B.n204 VSUBS 0.009985f
C263 B.n205 VSUBS 0.009985f
C264 B.n206 VSUBS 0.009985f
C265 B.n207 VSUBS 0.009985f
C266 B.n208 VSUBS 0.009985f
C267 B.n209 VSUBS 0.009985f
C268 B.n210 VSUBS 0.009985f
C269 B.n211 VSUBS 0.009985f
C270 B.n212 VSUBS 0.009985f
C271 B.n213 VSUBS 0.009985f
C272 B.n214 VSUBS 0.009985f
C273 B.n215 VSUBS 0.009985f
C274 B.n216 VSUBS 0.009985f
C275 B.n217 VSUBS 0.009985f
C276 B.n218 VSUBS 0.009985f
C277 B.n219 VSUBS 0.009985f
C278 B.n220 VSUBS 0.009985f
C279 B.n221 VSUBS 0.023103f
C280 B.n222 VSUBS 0.023593f
C281 B.n223 VSUBS 0.023593f
C282 B.n224 VSUBS 0.009985f
C283 B.n225 VSUBS 0.009985f
C284 B.n226 VSUBS 0.009985f
C285 B.n227 VSUBS 0.009985f
C286 B.n228 VSUBS 0.009985f
C287 B.n229 VSUBS 0.009985f
C288 B.n230 VSUBS 0.009985f
C289 B.n231 VSUBS 0.009985f
C290 B.n232 VSUBS 0.009985f
C291 B.n233 VSUBS 0.009985f
C292 B.n234 VSUBS 0.009985f
C293 B.n235 VSUBS 0.009985f
C294 B.n236 VSUBS 0.009985f
C295 B.n237 VSUBS 0.006902f
C296 B.n238 VSUBS 0.009985f
C297 B.n239 VSUBS 0.009985f
C298 B.n240 VSUBS 0.008076f
C299 B.n241 VSUBS 0.009985f
C300 B.n242 VSUBS 0.009985f
C301 B.n243 VSUBS 0.009985f
C302 B.n244 VSUBS 0.009985f
C303 B.n245 VSUBS 0.009985f
C304 B.n246 VSUBS 0.009985f
C305 B.n247 VSUBS 0.009985f
C306 B.n248 VSUBS 0.009985f
C307 B.n249 VSUBS 0.009985f
C308 B.n250 VSUBS 0.009985f
C309 B.n251 VSUBS 0.009985f
C310 B.n252 VSUBS 0.008076f
C311 B.n253 VSUBS 0.023135f
C312 B.n254 VSUBS 0.006902f
C313 B.n255 VSUBS 0.009985f
C314 B.n256 VSUBS 0.009985f
C315 B.n257 VSUBS 0.009985f
C316 B.n258 VSUBS 0.009985f
C317 B.n259 VSUBS 0.009985f
C318 B.n260 VSUBS 0.009985f
C319 B.n261 VSUBS 0.009985f
C320 B.n262 VSUBS 0.009985f
C321 B.n263 VSUBS 0.009985f
C322 B.n264 VSUBS 0.009985f
C323 B.n265 VSUBS 0.009985f
C324 B.n266 VSUBS 0.009985f
C325 B.n267 VSUBS 0.009985f
C326 B.n268 VSUBS 0.009985f
C327 B.n269 VSUBS 0.023593f
C328 B.n270 VSUBS 0.023103f
C329 B.n271 VSUBS 0.023103f
C330 B.n272 VSUBS 0.009985f
C331 B.n273 VSUBS 0.009985f
C332 B.n274 VSUBS 0.009985f
C333 B.n275 VSUBS 0.009985f
C334 B.n276 VSUBS 0.009985f
C335 B.n277 VSUBS 0.009985f
C336 B.n278 VSUBS 0.009985f
C337 B.n279 VSUBS 0.009985f
C338 B.n280 VSUBS 0.009985f
C339 B.n281 VSUBS 0.009985f
C340 B.n282 VSUBS 0.009985f
C341 B.n283 VSUBS 0.009985f
C342 B.n284 VSUBS 0.009985f
C343 B.n285 VSUBS 0.009985f
C344 B.n286 VSUBS 0.009985f
C345 B.n287 VSUBS 0.009985f
C346 B.n288 VSUBS 0.009985f
C347 B.n289 VSUBS 0.009985f
C348 B.n290 VSUBS 0.009985f
C349 B.n291 VSUBS 0.009985f
C350 B.n292 VSUBS 0.009985f
C351 B.n293 VSUBS 0.009985f
C352 B.n294 VSUBS 0.009985f
C353 B.n295 VSUBS 0.009985f
C354 B.n296 VSUBS 0.009985f
C355 B.n297 VSUBS 0.009985f
C356 B.n298 VSUBS 0.009985f
C357 B.n299 VSUBS 0.01303f
C358 B.n300 VSUBS 0.013881f
C359 B.n301 VSUBS 0.027603f
.ends

