* NGSPICE file created from diff_pair_sample_1717.ext - technology: sky130A

.subckt diff_pair_sample_1717 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.2884 pd=27.9 as=5.2884 ps=27.9 w=13.56 l=3.25
X1 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=5.2884 pd=27.9 as=0 ps=0 w=13.56 l=3.25
X2 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=5.2884 pd=27.9 as=0 ps=0 w=13.56 l=3.25
X3 VDD1.t0 VP.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=5.2884 pd=27.9 as=5.2884 ps=27.9 w=13.56 l=3.25
X4 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=5.2884 pd=27.9 as=5.2884 ps=27.9 w=13.56 l=3.25
X5 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.2884 pd=27.9 as=5.2884 ps=27.9 w=13.56 l=3.25
X6 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.2884 pd=27.9 as=0 ps=0 w=13.56 l=3.25
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=5.2884 pd=27.9 as=0 ps=0 w=13.56 l=3.25
R0 VP.n0 VP.t1 186.845
R1 VP.n0 VP.t0 139.284
R2 VP VP.n0 0.526368
R3 VTAIL.n290 VTAIL.n222 289.615
R4 VTAIL.n68 VTAIL.n0 289.615
R5 VTAIL.n216 VTAIL.n148 289.615
R6 VTAIL.n142 VTAIL.n74 289.615
R7 VTAIL.n247 VTAIL.n246 185
R8 VTAIL.n249 VTAIL.n248 185
R9 VTAIL.n242 VTAIL.n241 185
R10 VTAIL.n255 VTAIL.n254 185
R11 VTAIL.n257 VTAIL.n256 185
R12 VTAIL.n238 VTAIL.n237 185
R13 VTAIL.n264 VTAIL.n263 185
R14 VTAIL.n265 VTAIL.n236 185
R15 VTAIL.n267 VTAIL.n266 185
R16 VTAIL.n234 VTAIL.n233 185
R17 VTAIL.n273 VTAIL.n272 185
R18 VTAIL.n275 VTAIL.n274 185
R19 VTAIL.n230 VTAIL.n229 185
R20 VTAIL.n281 VTAIL.n280 185
R21 VTAIL.n283 VTAIL.n282 185
R22 VTAIL.n226 VTAIL.n225 185
R23 VTAIL.n289 VTAIL.n288 185
R24 VTAIL.n291 VTAIL.n290 185
R25 VTAIL.n25 VTAIL.n24 185
R26 VTAIL.n27 VTAIL.n26 185
R27 VTAIL.n20 VTAIL.n19 185
R28 VTAIL.n33 VTAIL.n32 185
R29 VTAIL.n35 VTAIL.n34 185
R30 VTAIL.n16 VTAIL.n15 185
R31 VTAIL.n42 VTAIL.n41 185
R32 VTAIL.n43 VTAIL.n14 185
R33 VTAIL.n45 VTAIL.n44 185
R34 VTAIL.n12 VTAIL.n11 185
R35 VTAIL.n51 VTAIL.n50 185
R36 VTAIL.n53 VTAIL.n52 185
R37 VTAIL.n8 VTAIL.n7 185
R38 VTAIL.n59 VTAIL.n58 185
R39 VTAIL.n61 VTAIL.n60 185
R40 VTAIL.n4 VTAIL.n3 185
R41 VTAIL.n67 VTAIL.n66 185
R42 VTAIL.n69 VTAIL.n68 185
R43 VTAIL.n217 VTAIL.n216 185
R44 VTAIL.n215 VTAIL.n214 185
R45 VTAIL.n152 VTAIL.n151 185
R46 VTAIL.n209 VTAIL.n208 185
R47 VTAIL.n207 VTAIL.n206 185
R48 VTAIL.n156 VTAIL.n155 185
R49 VTAIL.n201 VTAIL.n200 185
R50 VTAIL.n199 VTAIL.n198 185
R51 VTAIL.n160 VTAIL.n159 185
R52 VTAIL.n164 VTAIL.n162 185
R53 VTAIL.n193 VTAIL.n192 185
R54 VTAIL.n191 VTAIL.n190 185
R55 VTAIL.n166 VTAIL.n165 185
R56 VTAIL.n185 VTAIL.n184 185
R57 VTAIL.n183 VTAIL.n182 185
R58 VTAIL.n170 VTAIL.n169 185
R59 VTAIL.n177 VTAIL.n176 185
R60 VTAIL.n175 VTAIL.n174 185
R61 VTAIL.n143 VTAIL.n142 185
R62 VTAIL.n141 VTAIL.n140 185
R63 VTAIL.n78 VTAIL.n77 185
R64 VTAIL.n135 VTAIL.n134 185
R65 VTAIL.n133 VTAIL.n132 185
R66 VTAIL.n82 VTAIL.n81 185
R67 VTAIL.n127 VTAIL.n126 185
R68 VTAIL.n125 VTAIL.n124 185
R69 VTAIL.n86 VTAIL.n85 185
R70 VTAIL.n90 VTAIL.n88 185
R71 VTAIL.n119 VTAIL.n118 185
R72 VTAIL.n117 VTAIL.n116 185
R73 VTAIL.n92 VTAIL.n91 185
R74 VTAIL.n111 VTAIL.n110 185
R75 VTAIL.n109 VTAIL.n108 185
R76 VTAIL.n96 VTAIL.n95 185
R77 VTAIL.n103 VTAIL.n102 185
R78 VTAIL.n101 VTAIL.n100 185
R79 VTAIL.n245 VTAIL.t0 149.524
R80 VTAIL.n23 VTAIL.t1 149.524
R81 VTAIL.n173 VTAIL.t2 149.524
R82 VTAIL.n99 VTAIL.t3 149.524
R83 VTAIL.n248 VTAIL.n247 104.615
R84 VTAIL.n248 VTAIL.n241 104.615
R85 VTAIL.n255 VTAIL.n241 104.615
R86 VTAIL.n256 VTAIL.n255 104.615
R87 VTAIL.n256 VTAIL.n237 104.615
R88 VTAIL.n264 VTAIL.n237 104.615
R89 VTAIL.n265 VTAIL.n264 104.615
R90 VTAIL.n266 VTAIL.n265 104.615
R91 VTAIL.n266 VTAIL.n233 104.615
R92 VTAIL.n273 VTAIL.n233 104.615
R93 VTAIL.n274 VTAIL.n273 104.615
R94 VTAIL.n274 VTAIL.n229 104.615
R95 VTAIL.n281 VTAIL.n229 104.615
R96 VTAIL.n282 VTAIL.n281 104.615
R97 VTAIL.n282 VTAIL.n225 104.615
R98 VTAIL.n289 VTAIL.n225 104.615
R99 VTAIL.n290 VTAIL.n289 104.615
R100 VTAIL.n26 VTAIL.n25 104.615
R101 VTAIL.n26 VTAIL.n19 104.615
R102 VTAIL.n33 VTAIL.n19 104.615
R103 VTAIL.n34 VTAIL.n33 104.615
R104 VTAIL.n34 VTAIL.n15 104.615
R105 VTAIL.n42 VTAIL.n15 104.615
R106 VTAIL.n43 VTAIL.n42 104.615
R107 VTAIL.n44 VTAIL.n43 104.615
R108 VTAIL.n44 VTAIL.n11 104.615
R109 VTAIL.n51 VTAIL.n11 104.615
R110 VTAIL.n52 VTAIL.n51 104.615
R111 VTAIL.n52 VTAIL.n7 104.615
R112 VTAIL.n59 VTAIL.n7 104.615
R113 VTAIL.n60 VTAIL.n59 104.615
R114 VTAIL.n60 VTAIL.n3 104.615
R115 VTAIL.n67 VTAIL.n3 104.615
R116 VTAIL.n68 VTAIL.n67 104.615
R117 VTAIL.n216 VTAIL.n215 104.615
R118 VTAIL.n215 VTAIL.n151 104.615
R119 VTAIL.n208 VTAIL.n151 104.615
R120 VTAIL.n208 VTAIL.n207 104.615
R121 VTAIL.n207 VTAIL.n155 104.615
R122 VTAIL.n200 VTAIL.n155 104.615
R123 VTAIL.n200 VTAIL.n199 104.615
R124 VTAIL.n199 VTAIL.n159 104.615
R125 VTAIL.n164 VTAIL.n159 104.615
R126 VTAIL.n192 VTAIL.n164 104.615
R127 VTAIL.n192 VTAIL.n191 104.615
R128 VTAIL.n191 VTAIL.n165 104.615
R129 VTAIL.n184 VTAIL.n165 104.615
R130 VTAIL.n184 VTAIL.n183 104.615
R131 VTAIL.n183 VTAIL.n169 104.615
R132 VTAIL.n176 VTAIL.n169 104.615
R133 VTAIL.n176 VTAIL.n175 104.615
R134 VTAIL.n142 VTAIL.n141 104.615
R135 VTAIL.n141 VTAIL.n77 104.615
R136 VTAIL.n134 VTAIL.n77 104.615
R137 VTAIL.n134 VTAIL.n133 104.615
R138 VTAIL.n133 VTAIL.n81 104.615
R139 VTAIL.n126 VTAIL.n81 104.615
R140 VTAIL.n126 VTAIL.n125 104.615
R141 VTAIL.n125 VTAIL.n85 104.615
R142 VTAIL.n90 VTAIL.n85 104.615
R143 VTAIL.n118 VTAIL.n90 104.615
R144 VTAIL.n118 VTAIL.n117 104.615
R145 VTAIL.n117 VTAIL.n91 104.615
R146 VTAIL.n110 VTAIL.n91 104.615
R147 VTAIL.n110 VTAIL.n109 104.615
R148 VTAIL.n109 VTAIL.n95 104.615
R149 VTAIL.n102 VTAIL.n95 104.615
R150 VTAIL.n102 VTAIL.n101 104.615
R151 VTAIL.n247 VTAIL.t0 52.3082
R152 VTAIL.n25 VTAIL.t1 52.3082
R153 VTAIL.n175 VTAIL.t2 52.3082
R154 VTAIL.n101 VTAIL.t3 52.3082
R155 VTAIL.n295 VTAIL.n294 32.1853
R156 VTAIL.n73 VTAIL.n72 32.1853
R157 VTAIL.n221 VTAIL.n220 32.1853
R158 VTAIL.n147 VTAIL.n146 32.1853
R159 VTAIL.n147 VTAIL.n73 30.2289
R160 VTAIL.n295 VTAIL.n221 27.1427
R161 VTAIL.n267 VTAIL.n234 13.1884
R162 VTAIL.n45 VTAIL.n12 13.1884
R163 VTAIL.n162 VTAIL.n160 13.1884
R164 VTAIL.n88 VTAIL.n86 13.1884
R165 VTAIL.n268 VTAIL.n236 12.8005
R166 VTAIL.n272 VTAIL.n271 12.8005
R167 VTAIL.n46 VTAIL.n14 12.8005
R168 VTAIL.n50 VTAIL.n49 12.8005
R169 VTAIL.n198 VTAIL.n197 12.8005
R170 VTAIL.n194 VTAIL.n193 12.8005
R171 VTAIL.n124 VTAIL.n123 12.8005
R172 VTAIL.n120 VTAIL.n119 12.8005
R173 VTAIL.n263 VTAIL.n262 12.0247
R174 VTAIL.n275 VTAIL.n232 12.0247
R175 VTAIL.n41 VTAIL.n40 12.0247
R176 VTAIL.n53 VTAIL.n10 12.0247
R177 VTAIL.n201 VTAIL.n158 12.0247
R178 VTAIL.n190 VTAIL.n163 12.0247
R179 VTAIL.n127 VTAIL.n84 12.0247
R180 VTAIL.n116 VTAIL.n89 12.0247
R181 VTAIL.n261 VTAIL.n238 11.249
R182 VTAIL.n276 VTAIL.n230 11.249
R183 VTAIL.n39 VTAIL.n16 11.249
R184 VTAIL.n54 VTAIL.n8 11.249
R185 VTAIL.n202 VTAIL.n156 11.249
R186 VTAIL.n189 VTAIL.n166 11.249
R187 VTAIL.n128 VTAIL.n82 11.249
R188 VTAIL.n115 VTAIL.n92 11.249
R189 VTAIL.n258 VTAIL.n257 10.4732
R190 VTAIL.n280 VTAIL.n279 10.4732
R191 VTAIL.n36 VTAIL.n35 10.4732
R192 VTAIL.n58 VTAIL.n57 10.4732
R193 VTAIL.n206 VTAIL.n205 10.4732
R194 VTAIL.n186 VTAIL.n185 10.4732
R195 VTAIL.n132 VTAIL.n131 10.4732
R196 VTAIL.n112 VTAIL.n111 10.4732
R197 VTAIL.n246 VTAIL.n245 10.2747
R198 VTAIL.n24 VTAIL.n23 10.2747
R199 VTAIL.n174 VTAIL.n173 10.2747
R200 VTAIL.n100 VTAIL.n99 10.2747
R201 VTAIL.n254 VTAIL.n240 9.69747
R202 VTAIL.n283 VTAIL.n228 9.69747
R203 VTAIL.n32 VTAIL.n18 9.69747
R204 VTAIL.n61 VTAIL.n6 9.69747
R205 VTAIL.n209 VTAIL.n154 9.69747
R206 VTAIL.n182 VTAIL.n168 9.69747
R207 VTAIL.n135 VTAIL.n80 9.69747
R208 VTAIL.n108 VTAIL.n94 9.69747
R209 VTAIL.n294 VTAIL.n293 9.45567
R210 VTAIL.n72 VTAIL.n71 9.45567
R211 VTAIL.n220 VTAIL.n219 9.45567
R212 VTAIL.n146 VTAIL.n145 9.45567
R213 VTAIL.n293 VTAIL.n292 9.3005
R214 VTAIL.n287 VTAIL.n286 9.3005
R215 VTAIL.n285 VTAIL.n284 9.3005
R216 VTAIL.n228 VTAIL.n227 9.3005
R217 VTAIL.n279 VTAIL.n278 9.3005
R218 VTAIL.n277 VTAIL.n276 9.3005
R219 VTAIL.n232 VTAIL.n231 9.3005
R220 VTAIL.n271 VTAIL.n270 9.3005
R221 VTAIL.n244 VTAIL.n243 9.3005
R222 VTAIL.n251 VTAIL.n250 9.3005
R223 VTAIL.n253 VTAIL.n252 9.3005
R224 VTAIL.n240 VTAIL.n239 9.3005
R225 VTAIL.n259 VTAIL.n258 9.3005
R226 VTAIL.n261 VTAIL.n260 9.3005
R227 VTAIL.n262 VTAIL.n235 9.3005
R228 VTAIL.n269 VTAIL.n268 9.3005
R229 VTAIL.n224 VTAIL.n223 9.3005
R230 VTAIL.n71 VTAIL.n70 9.3005
R231 VTAIL.n65 VTAIL.n64 9.3005
R232 VTAIL.n63 VTAIL.n62 9.3005
R233 VTAIL.n6 VTAIL.n5 9.3005
R234 VTAIL.n57 VTAIL.n56 9.3005
R235 VTAIL.n55 VTAIL.n54 9.3005
R236 VTAIL.n10 VTAIL.n9 9.3005
R237 VTAIL.n49 VTAIL.n48 9.3005
R238 VTAIL.n22 VTAIL.n21 9.3005
R239 VTAIL.n29 VTAIL.n28 9.3005
R240 VTAIL.n31 VTAIL.n30 9.3005
R241 VTAIL.n18 VTAIL.n17 9.3005
R242 VTAIL.n37 VTAIL.n36 9.3005
R243 VTAIL.n39 VTAIL.n38 9.3005
R244 VTAIL.n40 VTAIL.n13 9.3005
R245 VTAIL.n47 VTAIL.n46 9.3005
R246 VTAIL.n2 VTAIL.n1 9.3005
R247 VTAIL.n172 VTAIL.n171 9.3005
R248 VTAIL.n179 VTAIL.n178 9.3005
R249 VTAIL.n181 VTAIL.n180 9.3005
R250 VTAIL.n168 VTAIL.n167 9.3005
R251 VTAIL.n187 VTAIL.n186 9.3005
R252 VTAIL.n189 VTAIL.n188 9.3005
R253 VTAIL.n163 VTAIL.n161 9.3005
R254 VTAIL.n195 VTAIL.n194 9.3005
R255 VTAIL.n219 VTAIL.n218 9.3005
R256 VTAIL.n150 VTAIL.n149 9.3005
R257 VTAIL.n213 VTAIL.n212 9.3005
R258 VTAIL.n211 VTAIL.n210 9.3005
R259 VTAIL.n154 VTAIL.n153 9.3005
R260 VTAIL.n205 VTAIL.n204 9.3005
R261 VTAIL.n203 VTAIL.n202 9.3005
R262 VTAIL.n158 VTAIL.n157 9.3005
R263 VTAIL.n197 VTAIL.n196 9.3005
R264 VTAIL.n98 VTAIL.n97 9.3005
R265 VTAIL.n105 VTAIL.n104 9.3005
R266 VTAIL.n107 VTAIL.n106 9.3005
R267 VTAIL.n94 VTAIL.n93 9.3005
R268 VTAIL.n113 VTAIL.n112 9.3005
R269 VTAIL.n115 VTAIL.n114 9.3005
R270 VTAIL.n89 VTAIL.n87 9.3005
R271 VTAIL.n121 VTAIL.n120 9.3005
R272 VTAIL.n145 VTAIL.n144 9.3005
R273 VTAIL.n76 VTAIL.n75 9.3005
R274 VTAIL.n139 VTAIL.n138 9.3005
R275 VTAIL.n137 VTAIL.n136 9.3005
R276 VTAIL.n80 VTAIL.n79 9.3005
R277 VTAIL.n131 VTAIL.n130 9.3005
R278 VTAIL.n129 VTAIL.n128 9.3005
R279 VTAIL.n84 VTAIL.n83 9.3005
R280 VTAIL.n123 VTAIL.n122 9.3005
R281 VTAIL.n253 VTAIL.n242 8.92171
R282 VTAIL.n284 VTAIL.n226 8.92171
R283 VTAIL.n31 VTAIL.n20 8.92171
R284 VTAIL.n62 VTAIL.n4 8.92171
R285 VTAIL.n210 VTAIL.n152 8.92171
R286 VTAIL.n181 VTAIL.n170 8.92171
R287 VTAIL.n136 VTAIL.n78 8.92171
R288 VTAIL.n107 VTAIL.n96 8.92171
R289 VTAIL.n250 VTAIL.n249 8.14595
R290 VTAIL.n288 VTAIL.n287 8.14595
R291 VTAIL.n28 VTAIL.n27 8.14595
R292 VTAIL.n66 VTAIL.n65 8.14595
R293 VTAIL.n214 VTAIL.n213 8.14595
R294 VTAIL.n178 VTAIL.n177 8.14595
R295 VTAIL.n140 VTAIL.n139 8.14595
R296 VTAIL.n104 VTAIL.n103 8.14595
R297 VTAIL.n246 VTAIL.n244 7.3702
R298 VTAIL.n291 VTAIL.n224 7.3702
R299 VTAIL.n294 VTAIL.n222 7.3702
R300 VTAIL.n24 VTAIL.n22 7.3702
R301 VTAIL.n69 VTAIL.n2 7.3702
R302 VTAIL.n72 VTAIL.n0 7.3702
R303 VTAIL.n220 VTAIL.n148 7.3702
R304 VTAIL.n217 VTAIL.n150 7.3702
R305 VTAIL.n174 VTAIL.n172 7.3702
R306 VTAIL.n146 VTAIL.n74 7.3702
R307 VTAIL.n143 VTAIL.n76 7.3702
R308 VTAIL.n100 VTAIL.n98 7.3702
R309 VTAIL.n292 VTAIL.n291 6.59444
R310 VTAIL.n292 VTAIL.n222 6.59444
R311 VTAIL.n70 VTAIL.n69 6.59444
R312 VTAIL.n70 VTAIL.n0 6.59444
R313 VTAIL.n218 VTAIL.n148 6.59444
R314 VTAIL.n218 VTAIL.n217 6.59444
R315 VTAIL.n144 VTAIL.n74 6.59444
R316 VTAIL.n144 VTAIL.n143 6.59444
R317 VTAIL.n249 VTAIL.n244 5.81868
R318 VTAIL.n288 VTAIL.n224 5.81868
R319 VTAIL.n27 VTAIL.n22 5.81868
R320 VTAIL.n66 VTAIL.n2 5.81868
R321 VTAIL.n214 VTAIL.n150 5.81868
R322 VTAIL.n177 VTAIL.n172 5.81868
R323 VTAIL.n140 VTAIL.n76 5.81868
R324 VTAIL.n103 VTAIL.n98 5.81868
R325 VTAIL.n250 VTAIL.n242 5.04292
R326 VTAIL.n287 VTAIL.n226 5.04292
R327 VTAIL.n28 VTAIL.n20 5.04292
R328 VTAIL.n65 VTAIL.n4 5.04292
R329 VTAIL.n213 VTAIL.n152 5.04292
R330 VTAIL.n178 VTAIL.n170 5.04292
R331 VTAIL.n139 VTAIL.n78 5.04292
R332 VTAIL.n104 VTAIL.n96 5.04292
R333 VTAIL.n254 VTAIL.n253 4.26717
R334 VTAIL.n284 VTAIL.n283 4.26717
R335 VTAIL.n32 VTAIL.n31 4.26717
R336 VTAIL.n62 VTAIL.n61 4.26717
R337 VTAIL.n210 VTAIL.n209 4.26717
R338 VTAIL.n182 VTAIL.n181 4.26717
R339 VTAIL.n136 VTAIL.n135 4.26717
R340 VTAIL.n108 VTAIL.n107 4.26717
R341 VTAIL.n257 VTAIL.n240 3.49141
R342 VTAIL.n280 VTAIL.n228 3.49141
R343 VTAIL.n35 VTAIL.n18 3.49141
R344 VTAIL.n58 VTAIL.n6 3.49141
R345 VTAIL.n206 VTAIL.n154 3.49141
R346 VTAIL.n185 VTAIL.n168 3.49141
R347 VTAIL.n132 VTAIL.n80 3.49141
R348 VTAIL.n111 VTAIL.n94 3.49141
R349 VTAIL.n245 VTAIL.n243 2.84303
R350 VTAIL.n23 VTAIL.n21 2.84303
R351 VTAIL.n173 VTAIL.n171 2.84303
R352 VTAIL.n99 VTAIL.n97 2.84303
R353 VTAIL.n258 VTAIL.n238 2.71565
R354 VTAIL.n279 VTAIL.n230 2.71565
R355 VTAIL.n36 VTAIL.n16 2.71565
R356 VTAIL.n57 VTAIL.n8 2.71565
R357 VTAIL.n205 VTAIL.n156 2.71565
R358 VTAIL.n186 VTAIL.n166 2.71565
R359 VTAIL.n131 VTAIL.n82 2.71565
R360 VTAIL.n112 VTAIL.n92 2.71565
R361 VTAIL.n221 VTAIL.n147 2.01343
R362 VTAIL.n263 VTAIL.n261 1.93989
R363 VTAIL.n276 VTAIL.n275 1.93989
R364 VTAIL.n41 VTAIL.n39 1.93989
R365 VTAIL.n54 VTAIL.n53 1.93989
R366 VTAIL.n202 VTAIL.n201 1.93989
R367 VTAIL.n190 VTAIL.n189 1.93989
R368 VTAIL.n128 VTAIL.n127 1.93989
R369 VTAIL.n116 VTAIL.n115 1.93989
R370 VTAIL VTAIL.n73 1.30007
R371 VTAIL.n262 VTAIL.n236 1.16414
R372 VTAIL.n272 VTAIL.n232 1.16414
R373 VTAIL.n40 VTAIL.n14 1.16414
R374 VTAIL.n50 VTAIL.n10 1.16414
R375 VTAIL.n198 VTAIL.n158 1.16414
R376 VTAIL.n193 VTAIL.n163 1.16414
R377 VTAIL.n124 VTAIL.n84 1.16414
R378 VTAIL.n119 VTAIL.n89 1.16414
R379 VTAIL VTAIL.n295 0.713862
R380 VTAIL.n268 VTAIL.n267 0.388379
R381 VTAIL.n271 VTAIL.n234 0.388379
R382 VTAIL.n46 VTAIL.n45 0.388379
R383 VTAIL.n49 VTAIL.n12 0.388379
R384 VTAIL.n197 VTAIL.n160 0.388379
R385 VTAIL.n194 VTAIL.n162 0.388379
R386 VTAIL.n123 VTAIL.n86 0.388379
R387 VTAIL.n120 VTAIL.n88 0.388379
R388 VTAIL.n251 VTAIL.n243 0.155672
R389 VTAIL.n252 VTAIL.n251 0.155672
R390 VTAIL.n252 VTAIL.n239 0.155672
R391 VTAIL.n259 VTAIL.n239 0.155672
R392 VTAIL.n260 VTAIL.n259 0.155672
R393 VTAIL.n260 VTAIL.n235 0.155672
R394 VTAIL.n269 VTAIL.n235 0.155672
R395 VTAIL.n270 VTAIL.n269 0.155672
R396 VTAIL.n270 VTAIL.n231 0.155672
R397 VTAIL.n277 VTAIL.n231 0.155672
R398 VTAIL.n278 VTAIL.n277 0.155672
R399 VTAIL.n278 VTAIL.n227 0.155672
R400 VTAIL.n285 VTAIL.n227 0.155672
R401 VTAIL.n286 VTAIL.n285 0.155672
R402 VTAIL.n286 VTAIL.n223 0.155672
R403 VTAIL.n293 VTAIL.n223 0.155672
R404 VTAIL.n29 VTAIL.n21 0.155672
R405 VTAIL.n30 VTAIL.n29 0.155672
R406 VTAIL.n30 VTAIL.n17 0.155672
R407 VTAIL.n37 VTAIL.n17 0.155672
R408 VTAIL.n38 VTAIL.n37 0.155672
R409 VTAIL.n38 VTAIL.n13 0.155672
R410 VTAIL.n47 VTAIL.n13 0.155672
R411 VTAIL.n48 VTAIL.n47 0.155672
R412 VTAIL.n48 VTAIL.n9 0.155672
R413 VTAIL.n55 VTAIL.n9 0.155672
R414 VTAIL.n56 VTAIL.n55 0.155672
R415 VTAIL.n56 VTAIL.n5 0.155672
R416 VTAIL.n63 VTAIL.n5 0.155672
R417 VTAIL.n64 VTAIL.n63 0.155672
R418 VTAIL.n64 VTAIL.n1 0.155672
R419 VTAIL.n71 VTAIL.n1 0.155672
R420 VTAIL.n219 VTAIL.n149 0.155672
R421 VTAIL.n212 VTAIL.n149 0.155672
R422 VTAIL.n212 VTAIL.n211 0.155672
R423 VTAIL.n211 VTAIL.n153 0.155672
R424 VTAIL.n204 VTAIL.n153 0.155672
R425 VTAIL.n204 VTAIL.n203 0.155672
R426 VTAIL.n203 VTAIL.n157 0.155672
R427 VTAIL.n196 VTAIL.n157 0.155672
R428 VTAIL.n196 VTAIL.n195 0.155672
R429 VTAIL.n195 VTAIL.n161 0.155672
R430 VTAIL.n188 VTAIL.n161 0.155672
R431 VTAIL.n188 VTAIL.n187 0.155672
R432 VTAIL.n187 VTAIL.n167 0.155672
R433 VTAIL.n180 VTAIL.n167 0.155672
R434 VTAIL.n180 VTAIL.n179 0.155672
R435 VTAIL.n179 VTAIL.n171 0.155672
R436 VTAIL.n145 VTAIL.n75 0.155672
R437 VTAIL.n138 VTAIL.n75 0.155672
R438 VTAIL.n138 VTAIL.n137 0.155672
R439 VTAIL.n137 VTAIL.n79 0.155672
R440 VTAIL.n130 VTAIL.n79 0.155672
R441 VTAIL.n130 VTAIL.n129 0.155672
R442 VTAIL.n129 VTAIL.n83 0.155672
R443 VTAIL.n122 VTAIL.n83 0.155672
R444 VTAIL.n122 VTAIL.n121 0.155672
R445 VTAIL.n121 VTAIL.n87 0.155672
R446 VTAIL.n114 VTAIL.n87 0.155672
R447 VTAIL.n114 VTAIL.n113 0.155672
R448 VTAIL.n113 VTAIL.n93 0.155672
R449 VTAIL.n106 VTAIL.n93 0.155672
R450 VTAIL.n106 VTAIL.n105 0.155672
R451 VTAIL.n105 VTAIL.n97 0.155672
R452 VDD1.n68 VDD1.n0 289.615
R453 VDD1.n141 VDD1.n73 289.615
R454 VDD1.n69 VDD1.n68 185
R455 VDD1.n67 VDD1.n66 185
R456 VDD1.n4 VDD1.n3 185
R457 VDD1.n61 VDD1.n60 185
R458 VDD1.n59 VDD1.n58 185
R459 VDD1.n8 VDD1.n7 185
R460 VDD1.n53 VDD1.n52 185
R461 VDD1.n51 VDD1.n50 185
R462 VDD1.n12 VDD1.n11 185
R463 VDD1.n16 VDD1.n14 185
R464 VDD1.n45 VDD1.n44 185
R465 VDD1.n43 VDD1.n42 185
R466 VDD1.n18 VDD1.n17 185
R467 VDD1.n37 VDD1.n36 185
R468 VDD1.n35 VDD1.n34 185
R469 VDD1.n22 VDD1.n21 185
R470 VDD1.n29 VDD1.n28 185
R471 VDD1.n27 VDD1.n26 185
R472 VDD1.n98 VDD1.n97 185
R473 VDD1.n100 VDD1.n99 185
R474 VDD1.n93 VDD1.n92 185
R475 VDD1.n106 VDD1.n105 185
R476 VDD1.n108 VDD1.n107 185
R477 VDD1.n89 VDD1.n88 185
R478 VDD1.n115 VDD1.n114 185
R479 VDD1.n116 VDD1.n87 185
R480 VDD1.n118 VDD1.n117 185
R481 VDD1.n85 VDD1.n84 185
R482 VDD1.n124 VDD1.n123 185
R483 VDD1.n126 VDD1.n125 185
R484 VDD1.n81 VDD1.n80 185
R485 VDD1.n132 VDD1.n131 185
R486 VDD1.n134 VDD1.n133 185
R487 VDD1.n77 VDD1.n76 185
R488 VDD1.n140 VDD1.n139 185
R489 VDD1.n142 VDD1.n141 185
R490 VDD1.n25 VDD1.t0 149.524
R491 VDD1.n96 VDD1.t1 149.524
R492 VDD1.n68 VDD1.n67 104.615
R493 VDD1.n67 VDD1.n3 104.615
R494 VDD1.n60 VDD1.n3 104.615
R495 VDD1.n60 VDD1.n59 104.615
R496 VDD1.n59 VDD1.n7 104.615
R497 VDD1.n52 VDD1.n7 104.615
R498 VDD1.n52 VDD1.n51 104.615
R499 VDD1.n51 VDD1.n11 104.615
R500 VDD1.n16 VDD1.n11 104.615
R501 VDD1.n44 VDD1.n16 104.615
R502 VDD1.n44 VDD1.n43 104.615
R503 VDD1.n43 VDD1.n17 104.615
R504 VDD1.n36 VDD1.n17 104.615
R505 VDD1.n36 VDD1.n35 104.615
R506 VDD1.n35 VDD1.n21 104.615
R507 VDD1.n28 VDD1.n21 104.615
R508 VDD1.n28 VDD1.n27 104.615
R509 VDD1.n99 VDD1.n98 104.615
R510 VDD1.n99 VDD1.n92 104.615
R511 VDD1.n106 VDD1.n92 104.615
R512 VDD1.n107 VDD1.n106 104.615
R513 VDD1.n107 VDD1.n88 104.615
R514 VDD1.n115 VDD1.n88 104.615
R515 VDD1.n116 VDD1.n115 104.615
R516 VDD1.n117 VDD1.n116 104.615
R517 VDD1.n117 VDD1.n84 104.615
R518 VDD1.n124 VDD1.n84 104.615
R519 VDD1.n125 VDD1.n124 104.615
R520 VDD1.n125 VDD1.n80 104.615
R521 VDD1.n132 VDD1.n80 104.615
R522 VDD1.n133 VDD1.n132 104.615
R523 VDD1.n133 VDD1.n76 104.615
R524 VDD1.n140 VDD1.n76 104.615
R525 VDD1.n141 VDD1.n140 104.615
R526 VDD1 VDD1.n145 91.682
R527 VDD1.n27 VDD1.t0 52.3082
R528 VDD1.n98 VDD1.t1 52.3082
R529 VDD1 VDD1.n72 49.6939
R530 VDD1.n14 VDD1.n12 13.1884
R531 VDD1.n118 VDD1.n85 13.1884
R532 VDD1.n50 VDD1.n49 12.8005
R533 VDD1.n46 VDD1.n45 12.8005
R534 VDD1.n119 VDD1.n87 12.8005
R535 VDD1.n123 VDD1.n122 12.8005
R536 VDD1.n53 VDD1.n10 12.0247
R537 VDD1.n42 VDD1.n15 12.0247
R538 VDD1.n114 VDD1.n113 12.0247
R539 VDD1.n126 VDD1.n83 12.0247
R540 VDD1.n54 VDD1.n8 11.249
R541 VDD1.n41 VDD1.n18 11.249
R542 VDD1.n112 VDD1.n89 11.249
R543 VDD1.n127 VDD1.n81 11.249
R544 VDD1.n58 VDD1.n57 10.4732
R545 VDD1.n38 VDD1.n37 10.4732
R546 VDD1.n109 VDD1.n108 10.4732
R547 VDD1.n131 VDD1.n130 10.4732
R548 VDD1.n26 VDD1.n25 10.2747
R549 VDD1.n97 VDD1.n96 10.2747
R550 VDD1.n61 VDD1.n6 9.69747
R551 VDD1.n34 VDD1.n20 9.69747
R552 VDD1.n105 VDD1.n91 9.69747
R553 VDD1.n134 VDD1.n79 9.69747
R554 VDD1.n72 VDD1.n71 9.45567
R555 VDD1.n145 VDD1.n144 9.45567
R556 VDD1.n24 VDD1.n23 9.3005
R557 VDD1.n31 VDD1.n30 9.3005
R558 VDD1.n33 VDD1.n32 9.3005
R559 VDD1.n20 VDD1.n19 9.3005
R560 VDD1.n39 VDD1.n38 9.3005
R561 VDD1.n41 VDD1.n40 9.3005
R562 VDD1.n15 VDD1.n13 9.3005
R563 VDD1.n47 VDD1.n46 9.3005
R564 VDD1.n71 VDD1.n70 9.3005
R565 VDD1.n2 VDD1.n1 9.3005
R566 VDD1.n65 VDD1.n64 9.3005
R567 VDD1.n63 VDD1.n62 9.3005
R568 VDD1.n6 VDD1.n5 9.3005
R569 VDD1.n57 VDD1.n56 9.3005
R570 VDD1.n55 VDD1.n54 9.3005
R571 VDD1.n10 VDD1.n9 9.3005
R572 VDD1.n49 VDD1.n48 9.3005
R573 VDD1.n144 VDD1.n143 9.3005
R574 VDD1.n138 VDD1.n137 9.3005
R575 VDD1.n136 VDD1.n135 9.3005
R576 VDD1.n79 VDD1.n78 9.3005
R577 VDD1.n130 VDD1.n129 9.3005
R578 VDD1.n128 VDD1.n127 9.3005
R579 VDD1.n83 VDD1.n82 9.3005
R580 VDD1.n122 VDD1.n121 9.3005
R581 VDD1.n95 VDD1.n94 9.3005
R582 VDD1.n102 VDD1.n101 9.3005
R583 VDD1.n104 VDD1.n103 9.3005
R584 VDD1.n91 VDD1.n90 9.3005
R585 VDD1.n110 VDD1.n109 9.3005
R586 VDD1.n112 VDD1.n111 9.3005
R587 VDD1.n113 VDD1.n86 9.3005
R588 VDD1.n120 VDD1.n119 9.3005
R589 VDD1.n75 VDD1.n74 9.3005
R590 VDD1.n62 VDD1.n4 8.92171
R591 VDD1.n33 VDD1.n22 8.92171
R592 VDD1.n104 VDD1.n93 8.92171
R593 VDD1.n135 VDD1.n77 8.92171
R594 VDD1.n66 VDD1.n65 8.14595
R595 VDD1.n30 VDD1.n29 8.14595
R596 VDD1.n101 VDD1.n100 8.14595
R597 VDD1.n139 VDD1.n138 8.14595
R598 VDD1.n72 VDD1.n0 7.3702
R599 VDD1.n69 VDD1.n2 7.3702
R600 VDD1.n26 VDD1.n24 7.3702
R601 VDD1.n97 VDD1.n95 7.3702
R602 VDD1.n142 VDD1.n75 7.3702
R603 VDD1.n145 VDD1.n73 7.3702
R604 VDD1.n70 VDD1.n0 6.59444
R605 VDD1.n70 VDD1.n69 6.59444
R606 VDD1.n143 VDD1.n142 6.59444
R607 VDD1.n143 VDD1.n73 6.59444
R608 VDD1.n66 VDD1.n2 5.81868
R609 VDD1.n29 VDD1.n24 5.81868
R610 VDD1.n100 VDD1.n95 5.81868
R611 VDD1.n139 VDD1.n75 5.81868
R612 VDD1.n65 VDD1.n4 5.04292
R613 VDD1.n30 VDD1.n22 5.04292
R614 VDD1.n101 VDD1.n93 5.04292
R615 VDD1.n138 VDD1.n77 5.04292
R616 VDD1.n62 VDD1.n61 4.26717
R617 VDD1.n34 VDD1.n33 4.26717
R618 VDD1.n105 VDD1.n104 4.26717
R619 VDD1.n135 VDD1.n134 4.26717
R620 VDD1.n58 VDD1.n6 3.49141
R621 VDD1.n37 VDD1.n20 3.49141
R622 VDD1.n108 VDD1.n91 3.49141
R623 VDD1.n131 VDD1.n79 3.49141
R624 VDD1.n25 VDD1.n23 2.84303
R625 VDD1.n96 VDD1.n94 2.84303
R626 VDD1.n57 VDD1.n8 2.71565
R627 VDD1.n38 VDD1.n18 2.71565
R628 VDD1.n109 VDD1.n89 2.71565
R629 VDD1.n130 VDD1.n81 2.71565
R630 VDD1.n54 VDD1.n53 1.93989
R631 VDD1.n42 VDD1.n41 1.93989
R632 VDD1.n114 VDD1.n112 1.93989
R633 VDD1.n127 VDD1.n126 1.93989
R634 VDD1.n50 VDD1.n10 1.16414
R635 VDD1.n45 VDD1.n15 1.16414
R636 VDD1.n113 VDD1.n87 1.16414
R637 VDD1.n123 VDD1.n83 1.16414
R638 VDD1.n49 VDD1.n12 0.388379
R639 VDD1.n46 VDD1.n14 0.388379
R640 VDD1.n119 VDD1.n118 0.388379
R641 VDD1.n122 VDD1.n85 0.388379
R642 VDD1.n71 VDD1.n1 0.155672
R643 VDD1.n64 VDD1.n1 0.155672
R644 VDD1.n64 VDD1.n63 0.155672
R645 VDD1.n63 VDD1.n5 0.155672
R646 VDD1.n56 VDD1.n5 0.155672
R647 VDD1.n56 VDD1.n55 0.155672
R648 VDD1.n55 VDD1.n9 0.155672
R649 VDD1.n48 VDD1.n9 0.155672
R650 VDD1.n48 VDD1.n47 0.155672
R651 VDD1.n47 VDD1.n13 0.155672
R652 VDD1.n40 VDD1.n13 0.155672
R653 VDD1.n40 VDD1.n39 0.155672
R654 VDD1.n39 VDD1.n19 0.155672
R655 VDD1.n32 VDD1.n19 0.155672
R656 VDD1.n32 VDD1.n31 0.155672
R657 VDD1.n31 VDD1.n23 0.155672
R658 VDD1.n102 VDD1.n94 0.155672
R659 VDD1.n103 VDD1.n102 0.155672
R660 VDD1.n103 VDD1.n90 0.155672
R661 VDD1.n110 VDD1.n90 0.155672
R662 VDD1.n111 VDD1.n110 0.155672
R663 VDD1.n111 VDD1.n86 0.155672
R664 VDD1.n120 VDD1.n86 0.155672
R665 VDD1.n121 VDD1.n120 0.155672
R666 VDD1.n121 VDD1.n82 0.155672
R667 VDD1.n128 VDD1.n82 0.155672
R668 VDD1.n129 VDD1.n128 0.155672
R669 VDD1.n129 VDD1.n78 0.155672
R670 VDD1.n136 VDD1.n78 0.155672
R671 VDD1.n137 VDD1.n136 0.155672
R672 VDD1.n137 VDD1.n74 0.155672
R673 VDD1.n144 VDD1.n74 0.155672
R674 B.n755 B.n754 585
R675 B.n313 B.n106 585
R676 B.n312 B.n311 585
R677 B.n310 B.n309 585
R678 B.n308 B.n307 585
R679 B.n306 B.n305 585
R680 B.n304 B.n303 585
R681 B.n302 B.n301 585
R682 B.n300 B.n299 585
R683 B.n298 B.n297 585
R684 B.n296 B.n295 585
R685 B.n294 B.n293 585
R686 B.n292 B.n291 585
R687 B.n290 B.n289 585
R688 B.n288 B.n287 585
R689 B.n286 B.n285 585
R690 B.n284 B.n283 585
R691 B.n282 B.n281 585
R692 B.n280 B.n279 585
R693 B.n278 B.n277 585
R694 B.n276 B.n275 585
R695 B.n274 B.n273 585
R696 B.n272 B.n271 585
R697 B.n270 B.n269 585
R698 B.n268 B.n267 585
R699 B.n266 B.n265 585
R700 B.n264 B.n263 585
R701 B.n262 B.n261 585
R702 B.n260 B.n259 585
R703 B.n258 B.n257 585
R704 B.n256 B.n255 585
R705 B.n254 B.n253 585
R706 B.n252 B.n251 585
R707 B.n250 B.n249 585
R708 B.n248 B.n247 585
R709 B.n246 B.n245 585
R710 B.n244 B.n243 585
R711 B.n242 B.n241 585
R712 B.n240 B.n239 585
R713 B.n238 B.n237 585
R714 B.n236 B.n235 585
R715 B.n234 B.n233 585
R716 B.n232 B.n231 585
R717 B.n230 B.n229 585
R718 B.n228 B.n227 585
R719 B.n226 B.n225 585
R720 B.n224 B.n223 585
R721 B.n222 B.n221 585
R722 B.n220 B.n219 585
R723 B.n218 B.n217 585
R724 B.n216 B.n215 585
R725 B.n214 B.n213 585
R726 B.n212 B.n211 585
R727 B.n210 B.n209 585
R728 B.n208 B.n207 585
R729 B.n206 B.n205 585
R730 B.n204 B.n203 585
R731 B.n202 B.n201 585
R732 B.n200 B.n199 585
R733 B.n198 B.n197 585
R734 B.n196 B.n195 585
R735 B.n194 B.n193 585
R736 B.n192 B.n191 585
R737 B.n190 B.n189 585
R738 B.n188 B.n187 585
R739 B.n186 B.n185 585
R740 B.n184 B.n183 585
R741 B.n182 B.n181 585
R742 B.n180 B.n179 585
R743 B.n178 B.n177 585
R744 B.n176 B.n175 585
R745 B.n174 B.n173 585
R746 B.n172 B.n171 585
R747 B.n170 B.n169 585
R748 B.n168 B.n167 585
R749 B.n166 B.n165 585
R750 B.n164 B.n163 585
R751 B.n162 B.n161 585
R752 B.n160 B.n159 585
R753 B.n158 B.n157 585
R754 B.n156 B.n155 585
R755 B.n154 B.n153 585
R756 B.n152 B.n151 585
R757 B.n150 B.n149 585
R758 B.n148 B.n147 585
R759 B.n146 B.n145 585
R760 B.n144 B.n143 585
R761 B.n142 B.n141 585
R762 B.n140 B.n139 585
R763 B.n138 B.n137 585
R764 B.n136 B.n135 585
R765 B.n134 B.n133 585
R766 B.n132 B.n131 585
R767 B.n130 B.n129 585
R768 B.n128 B.n127 585
R769 B.n126 B.n125 585
R770 B.n124 B.n123 585
R771 B.n122 B.n121 585
R772 B.n120 B.n119 585
R773 B.n118 B.n117 585
R774 B.n116 B.n115 585
R775 B.n114 B.n113 585
R776 B.n753 B.n55 585
R777 B.n758 B.n55 585
R778 B.n752 B.n54 585
R779 B.n759 B.n54 585
R780 B.n751 B.n750 585
R781 B.n750 B.n50 585
R782 B.n749 B.n49 585
R783 B.n765 B.n49 585
R784 B.n748 B.n48 585
R785 B.n766 B.n48 585
R786 B.n747 B.n47 585
R787 B.n767 B.n47 585
R788 B.n746 B.n745 585
R789 B.n745 B.n43 585
R790 B.n744 B.n42 585
R791 B.n773 B.n42 585
R792 B.n743 B.n41 585
R793 B.n774 B.n41 585
R794 B.n742 B.n40 585
R795 B.n775 B.n40 585
R796 B.n741 B.n740 585
R797 B.n740 B.n36 585
R798 B.n739 B.n35 585
R799 B.n781 B.n35 585
R800 B.n738 B.n34 585
R801 B.n782 B.n34 585
R802 B.n737 B.n33 585
R803 B.n783 B.n33 585
R804 B.n736 B.n735 585
R805 B.n735 B.n29 585
R806 B.n734 B.n28 585
R807 B.n789 B.n28 585
R808 B.n733 B.n27 585
R809 B.n790 B.n27 585
R810 B.n732 B.n26 585
R811 B.n791 B.n26 585
R812 B.n731 B.n730 585
R813 B.n730 B.n22 585
R814 B.n729 B.n21 585
R815 B.n797 B.n21 585
R816 B.n728 B.n20 585
R817 B.n798 B.n20 585
R818 B.n727 B.n19 585
R819 B.n799 B.n19 585
R820 B.n726 B.n725 585
R821 B.n725 B.n18 585
R822 B.n724 B.n14 585
R823 B.n805 B.n14 585
R824 B.n723 B.n13 585
R825 B.n806 B.n13 585
R826 B.n722 B.n12 585
R827 B.n807 B.n12 585
R828 B.n721 B.n720 585
R829 B.n720 B.n8 585
R830 B.n719 B.n7 585
R831 B.n813 B.n7 585
R832 B.n718 B.n6 585
R833 B.n814 B.n6 585
R834 B.n717 B.n5 585
R835 B.n815 B.n5 585
R836 B.n716 B.n715 585
R837 B.n715 B.n4 585
R838 B.n714 B.n314 585
R839 B.n714 B.n713 585
R840 B.n704 B.n315 585
R841 B.n316 B.n315 585
R842 B.n706 B.n705 585
R843 B.n707 B.n706 585
R844 B.n703 B.n321 585
R845 B.n321 B.n320 585
R846 B.n702 B.n701 585
R847 B.n701 B.n700 585
R848 B.n323 B.n322 585
R849 B.n693 B.n323 585
R850 B.n692 B.n691 585
R851 B.n694 B.n692 585
R852 B.n690 B.n328 585
R853 B.n328 B.n327 585
R854 B.n689 B.n688 585
R855 B.n688 B.n687 585
R856 B.n330 B.n329 585
R857 B.n331 B.n330 585
R858 B.n680 B.n679 585
R859 B.n681 B.n680 585
R860 B.n678 B.n336 585
R861 B.n336 B.n335 585
R862 B.n677 B.n676 585
R863 B.n676 B.n675 585
R864 B.n338 B.n337 585
R865 B.n339 B.n338 585
R866 B.n668 B.n667 585
R867 B.n669 B.n668 585
R868 B.n666 B.n344 585
R869 B.n344 B.n343 585
R870 B.n665 B.n664 585
R871 B.n664 B.n663 585
R872 B.n346 B.n345 585
R873 B.n347 B.n346 585
R874 B.n656 B.n655 585
R875 B.n657 B.n656 585
R876 B.n654 B.n351 585
R877 B.n355 B.n351 585
R878 B.n653 B.n652 585
R879 B.n652 B.n651 585
R880 B.n353 B.n352 585
R881 B.n354 B.n353 585
R882 B.n644 B.n643 585
R883 B.n645 B.n644 585
R884 B.n642 B.n360 585
R885 B.n360 B.n359 585
R886 B.n641 B.n640 585
R887 B.n640 B.n639 585
R888 B.n362 B.n361 585
R889 B.n363 B.n362 585
R890 B.n632 B.n631 585
R891 B.n633 B.n632 585
R892 B.n630 B.n368 585
R893 B.n368 B.n367 585
R894 B.n625 B.n624 585
R895 B.n623 B.n421 585
R896 B.n622 B.n420 585
R897 B.n627 B.n420 585
R898 B.n621 B.n620 585
R899 B.n619 B.n618 585
R900 B.n617 B.n616 585
R901 B.n615 B.n614 585
R902 B.n613 B.n612 585
R903 B.n611 B.n610 585
R904 B.n609 B.n608 585
R905 B.n607 B.n606 585
R906 B.n605 B.n604 585
R907 B.n603 B.n602 585
R908 B.n601 B.n600 585
R909 B.n599 B.n598 585
R910 B.n597 B.n596 585
R911 B.n595 B.n594 585
R912 B.n593 B.n592 585
R913 B.n591 B.n590 585
R914 B.n589 B.n588 585
R915 B.n587 B.n586 585
R916 B.n585 B.n584 585
R917 B.n583 B.n582 585
R918 B.n581 B.n580 585
R919 B.n579 B.n578 585
R920 B.n577 B.n576 585
R921 B.n575 B.n574 585
R922 B.n573 B.n572 585
R923 B.n571 B.n570 585
R924 B.n569 B.n568 585
R925 B.n567 B.n566 585
R926 B.n565 B.n564 585
R927 B.n563 B.n562 585
R928 B.n561 B.n560 585
R929 B.n559 B.n558 585
R930 B.n557 B.n556 585
R931 B.n555 B.n554 585
R932 B.n553 B.n552 585
R933 B.n551 B.n550 585
R934 B.n549 B.n548 585
R935 B.n547 B.n546 585
R936 B.n545 B.n544 585
R937 B.n543 B.n542 585
R938 B.n541 B.n540 585
R939 B.n539 B.n538 585
R940 B.n537 B.n536 585
R941 B.n534 B.n533 585
R942 B.n532 B.n531 585
R943 B.n530 B.n529 585
R944 B.n528 B.n527 585
R945 B.n526 B.n525 585
R946 B.n524 B.n523 585
R947 B.n522 B.n521 585
R948 B.n520 B.n519 585
R949 B.n518 B.n517 585
R950 B.n516 B.n515 585
R951 B.n513 B.n512 585
R952 B.n511 B.n510 585
R953 B.n509 B.n508 585
R954 B.n507 B.n506 585
R955 B.n505 B.n504 585
R956 B.n503 B.n502 585
R957 B.n501 B.n500 585
R958 B.n499 B.n498 585
R959 B.n497 B.n496 585
R960 B.n495 B.n494 585
R961 B.n493 B.n492 585
R962 B.n491 B.n490 585
R963 B.n489 B.n488 585
R964 B.n487 B.n486 585
R965 B.n485 B.n484 585
R966 B.n483 B.n482 585
R967 B.n481 B.n480 585
R968 B.n479 B.n478 585
R969 B.n477 B.n476 585
R970 B.n475 B.n474 585
R971 B.n473 B.n472 585
R972 B.n471 B.n470 585
R973 B.n469 B.n468 585
R974 B.n467 B.n466 585
R975 B.n465 B.n464 585
R976 B.n463 B.n462 585
R977 B.n461 B.n460 585
R978 B.n459 B.n458 585
R979 B.n457 B.n456 585
R980 B.n455 B.n454 585
R981 B.n453 B.n452 585
R982 B.n451 B.n450 585
R983 B.n449 B.n448 585
R984 B.n447 B.n446 585
R985 B.n445 B.n444 585
R986 B.n443 B.n442 585
R987 B.n441 B.n440 585
R988 B.n439 B.n438 585
R989 B.n437 B.n436 585
R990 B.n435 B.n434 585
R991 B.n433 B.n432 585
R992 B.n431 B.n430 585
R993 B.n429 B.n428 585
R994 B.n427 B.n426 585
R995 B.n370 B.n369 585
R996 B.n629 B.n628 585
R997 B.n628 B.n627 585
R998 B.n366 B.n365 585
R999 B.n367 B.n366 585
R1000 B.n635 B.n634 585
R1001 B.n634 B.n633 585
R1002 B.n636 B.n364 585
R1003 B.n364 B.n363 585
R1004 B.n638 B.n637 585
R1005 B.n639 B.n638 585
R1006 B.n358 B.n357 585
R1007 B.n359 B.n358 585
R1008 B.n647 B.n646 585
R1009 B.n646 B.n645 585
R1010 B.n648 B.n356 585
R1011 B.n356 B.n354 585
R1012 B.n650 B.n649 585
R1013 B.n651 B.n650 585
R1014 B.n350 B.n349 585
R1015 B.n355 B.n350 585
R1016 B.n659 B.n658 585
R1017 B.n658 B.n657 585
R1018 B.n660 B.n348 585
R1019 B.n348 B.n347 585
R1020 B.n662 B.n661 585
R1021 B.n663 B.n662 585
R1022 B.n342 B.n341 585
R1023 B.n343 B.n342 585
R1024 B.n671 B.n670 585
R1025 B.n670 B.n669 585
R1026 B.n672 B.n340 585
R1027 B.n340 B.n339 585
R1028 B.n674 B.n673 585
R1029 B.n675 B.n674 585
R1030 B.n334 B.n333 585
R1031 B.n335 B.n334 585
R1032 B.n683 B.n682 585
R1033 B.n682 B.n681 585
R1034 B.n684 B.n332 585
R1035 B.n332 B.n331 585
R1036 B.n686 B.n685 585
R1037 B.n687 B.n686 585
R1038 B.n326 B.n325 585
R1039 B.n327 B.n326 585
R1040 B.n696 B.n695 585
R1041 B.n695 B.n694 585
R1042 B.n697 B.n324 585
R1043 B.n693 B.n324 585
R1044 B.n699 B.n698 585
R1045 B.n700 B.n699 585
R1046 B.n319 B.n318 585
R1047 B.n320 B.n319 585
R1048 B.n709 B.n708 585
R1049 B.n708 B.n707 585
R1050 B.n710 B.n317 585
R1051 B.n317 B.n316 585
R1052 B.n712 B.n711 585
R1053 B.n713 B.n712 585
R1054 B.n2 B.n0 585
R1055 B.n4 B.n2 585
R1056 B.n3 B.n1 585
R1057 B.n814 B.n3 585
R1058 B.n812 B.n811 585
R1059 B.n813 B.n812 585
R1060 B.n810 B.n9 585
R1061 B.n9 B.n8 585
R1062 B.n809 B.n808 585
R1063 B.n808 B.n807 585
R1064 B.n11 B.n10 585
R1065 B.n806 B.n11 585
R1066 B.n804 B.n803 585
R1067 B.n805 B.n804 585
R1068 B.n802 B.n15 585
R1069 B.n18 B.n15 585
R1070 B.n801 B.n800 585
R1071 B.n800 B.n799 585
R1072 B.n17 B.n16 585
R1073 B.n798 B.n17 585
R1074 B.n796 B.n795 585
R1075 B.n797 B.n796 585
R1076 B.n794 B.n23 585
R1077 B.n23 B.n22 585
R1078 B.n793 B.n792 585
R1079 B.n792 B.n791 585
R1080 B.n25 B.n24 585
R1081 B.n790 B.n25 585
R1082 B.n788 B.n787 585
R1083 B.n789 B.n788 585
R1084 B.n786 B.n30 585
R1085 B.n30 B.n29 585
R1086 B.n785 B.n784 585
R1087 B.n784 B.n783 585
R1088 B.n32 B.n31 585
R1089 B.n782 B.n32 585
R1090 B.n780 B.n779 585
R1091 B.n781 B.n780 585
R1092 B.n778 B.n37 585
R1093 B.n37 B.n36 585
R1094 B.n777 B.n776 585
R1095 B.n776 B.n775 585
R1096 B.n39 B.n38 585
R1097 B.n774 B.n39 585
R1098 B.n772 B.n771 585
R1099 B.n773 B.n772 585
R1100 B.n770 B.n44 585
R1101 B.n44 B.n43 585
R1102 B.n769 B.n768 585
R1103 B.n768 B.n767 585
R1104 B.n46 B.n45 585
R1105 B.n766 B.n46 585
R1106 B.n764 B.n763 585
R1107 B.n765 B.n764 585
R1108 B.n762 B.n51 585
R1109 B.n51 B.n50 585
R1110 B.n761 B.n760 585
R1111 B.n760 B.n759 585
R1112 B.n53 B.n52 585
R1113 B.n758 B.n53 585
R1114 B.n817 B.n816 585
R1115 B.n816 B.n815 585
R1116 B.n625 B.n366 526.135
R1117 B.n113 B.n53 526.135
R1118 B.n628 B.n368 526.135
R1119 B.n755 B.n55 526.135
R1120 B.n424 B.t15 378.741
R1121 B.n107 B.t11 378.741
R1122 B.n422 B.t5 378.741
R1123 B.n110 B.t8 378.741
R1124 B.n424 B.t13 309.408
R1125 B.n422 B.t2 309.408
R1126 B.n110 B.t6 309.408
R1127 B.n107 B.t10 309.408
R1128 B.n425 B.t14 309.312
R1129 B.n108 B.t12 309.312
R1130 B.n423 B.t4 309.312
R1131 B.n111 B.t9 309.312
R1132 B.n757 B.n756 256.663
R1133 B.n757 B.n105 256.663
R1134 B.n757 B.n104 256.663
R1135 B.n757 B.n103 256.663
R1136 B.n757 B.n102 256.663
R1137 B.n757 B.n101 256.663
R1138 B.n757 B.n100 256.663
R1139 B.n757 B.n99 256.663
R1140 B.n757 B.n98 256.663
R1141 B.n757 B.n97 256.663
R1142 B.n757 B.n96 256.663
R1143 B.n757 B.n95 256.663
R1144 B.n757 B.n94 256.663
R1145 B.n757 B.n93 256.663
R1146 B.n757 B.n92 256.663
R1147 B.n757 B.n91 256.663
R1148 B.n757 B.n90 256.663
R1149 B.n757 B.n89 256.663
R1150 B.n757 B.n88 256.663
R1151 B.n757 B.n87 256.663
R1152 B.n757 B.n86 256.663
R1153 B.n757 B.n85 256.663
R1154 B.n757 B.n84 256.663
R1155 B.n757 B.n83 256.663
R1156 B.n757 B.n82 256.663
R1157 B.n757 B.n81 256.663
R1158 B.n757 B.n80 256.663
R1159 B.n757 B.n79 256.663
R1160 B.n757 B.n78 256.663
R1161 B.n757 B.n77 256.663
R1162 B.n757 B.n76 256.663
R1163 B.n757 B.n75 256.663
R1164 B.n757 B.n74 256.663
R1165 B.n757 B.n73 256.663
R1166 B.n757 B.n72 256.663
R1167 B.n757 B.n71 256.663
R1168 B.n757 B.n70 256.663
R1169 B.n757 B.n69 256.663
R1170 B.n757 B.n68 256.663
R1171 B.n757 B.n67 256.663
R1172 B.n757 B.n66 256.663
R1173 B.n757 B.n65 256.663
R1174 B.n757 B.n64 256.663
R1175 B.n757 B.n63 256.663
R1176 B.n757 B.n62 256.663
R1177 B.n757 B.n61 256.663
R1178 B.n757 B.n60 256.663
R1179 B.n757 B.n59 256.663
R1180 B.n757 B.n58 256.663
R1181 B.n757 B.n57 256.663
R1182 B.n757 B.n56 256.663
R1183 B.n627 B.n626 256.663
R1184 B.n627 B.n371 256.663
R1185 B.n627 B.n372 256.663
R1186 B.n627 B.n373 256.663
R1187 B.n627 B.n374 256.663
R1188 B.n627 B.n375 256.663
R1189 B.n627 B.n376 256.663
R1190 B.n627 B.n377 256.663
R1191 B.n627 B.n378 256.663
R1192 B.n627 B.n379 256.663
R1193 B.n627 B.n380 256.663
R1194 B.n627 B.n381 256.663
R1195 B.n627 B.n382 256.663
R1196 B.n627 B.n383 256.663
R1197 B.n627 B.n384 256.663
R1198 B.n627 B.n385 256.663
R1199 B.n627 B.n386 256.663
R1200 B.n627 B.n387 256.663
R1201 B.n627 B.n388 256.663
R1202 B.n627 B.n389 256.663
R1203 B.n627 B.n390 256.663
R1204 B.n627 B.n391 256.663
R1205 B.n627 B.n392 256.663
R1206 B.n627 B.n393 256.663
R1207 B.n627 B.n394 256.663
R1208 B.n627 B.n395 256.663
R1209 B.n627 B.n396 256.663
R1210 B.n627 B.n397 256.663
R1211 B.n627 B.n398 256.663
R1212 B.n627 B.n399 256.663
R1213 B.n627 B.n400 256.663
R1214 B.n627 B.n401 256.663
R1215 B.n627 B.n402 256.663
R1216 B.n627 B.n403 256.663
R1217 B.n627 B.n404 256.663
R1218 B.n627 B.n405 256.663
R1219 B.n627 B.n406 256.663
R1220 B.n627 B.n407 256.663
R1221 B.n627 B.n408 256.663
R1222 B.n627 B.n409 256.663
R1223 B.n627 B.n410 256.663
R1224 B.n627 B.n411 256.663
R1225 B.n627 B.n412 256.663
R1226 B.n627 B.n413 256.663
R1227 B.n627 B.n414 256.663
R1228 B.n627 B.n415 256.663
R1229 B.n627 B.n416 256.663
R1230 B.n627 B.n417 256.663
R1231 B.n627 B.n418 256.663
R1232 B.n627 B.n419 256.663
R1233 B.n634 B.n366 163.367
R1234 B.n634 B.n364 163.367
R1235 B.n638 B.n364 163.367
R1236 B.n638 B.n358 163.367
R1237 B.n646 B.n358 163.367
R1238 B.n646 B.n356 163.367
R1239 B.n650 B.n356 163.367
R1240 B.n650 B.n350 163.367
R1241 B.n658 B.n350 163.367
R1242 B.n658 B.n348 163.367
R1243 B.n662 B.n348 163.367
R1244 B.n662 B.n342 163.367
R1245 B.n670 B.n342 163.367
R1246 B.n670 B.n340 163.367
R1247 B.n674 B.n340 163.367
R1248 B.n674 B.n334 163.367
R1249 B.n682 B.n334 163.367
R1250 B.n682 B.n332 163.367
R1251 B.n686 B.n332 163.367
R1252 B.n686 B.n326 163.367
R1253 B.n695 B.n326 163.367
R1254 B.n695 B.n324 163.367
R1255 B.n699 B.n324 163.367
R1256 B.n699 B.n319 163.367
R1257 B.n708 B.n319 163.367
R1258 B.n708 B.n317 163.367
R1259 B.n712 B.n317 163.367
R1260 B.n712 B.n2 163.367
R1261 B.n816 B.n2 163.367
R1262 B.n816 B.n3 163.367
R1263 B.n812 B.n3 163.367
R1264 B.n812 B.n9 163.367
R1265 B.n808 B.n9 163.367
R1266 B.n808 B.n11 163.367
R1267 B.n804 B.n11 163.367
R1268 B.n804 B.n15 163.367
R1269 B.n800 B.n15 163.367
R1270 B.n800 B.n17 163.367
R1271 B.n796 B.n17 163.367
R1272 B.n796 B.n23 163.367
R1273 B.n792 B.n23 163.367
R1274 B.n792 B.n25 163.367
R1275 B.n788 B.n25 163.367
R1276 B.n788 B.n30 163.367
R1277 B.n784 B.n30 163.367
R1278 B.n784 B.n32 163.367
R1279 B.n780 B.n32 163.367
R1280 B.n780 B.n37 163.367
R1281 B.n776 B.n37 163.367
R1282 B.n776 B.n39 163.367
R1283 B.n772 B.n39 163.367
R1284 B.n772 B.n44 163.367
R1285 B.n768 B.n44 163.367
R1286 B.n768 B.n46 163.367
R1287 B.n764 B.n46 163.367
R1288 B.n764 B.n51 163.367
R1289 B.n760 B.n51 163.367
R1290 B.n760 B.n53 163.367
R1291 B.n421 B.n420 163.367
R1292 B.n620 B.n420 163.367
R1293 B.n618 B.n617 163.367
R1294 B.n614 B.n613 163.367
R1295 B.n610 B.n609 163.367
R1296 B.n606 B.n605 163.367
R1297 B.n602 B.n601 163.367
R1298 B.n598 B.n597 163.367
R1299 B.n594 B.n593 163.367
R1300 B.n590 B.n589 163.367
R1301 B.n586 B.n585 163.367
R1302 B.n582 B.n581 163.367
R1303 B.n578 B.n577 163.367
R1304 B.n574 B.n573 163.367
R1305 B.n570 B.n569 163.367
R1306 B.n566 B.n565 163.367
R1307 B.n562 B.n561 163.367
R1308 B.n558 B.n557 163.367
R1309 B.n554 B.n553 163.367
R1310 B.n550 B.n549 163.367
R1311 B.n546 B.n545 163.367
R1312 B.n542 B.n541 163.367
R1313 B.n538 B.n537 163.367
R1314 B.n533 B.n532 163.367
R1315 B.n529 B.n528 163.367
R1316 B.n525 B.n524 163.367
R1317 B.n521 B.n520 163.367
R1318 B.n517 B.n516 163.367
R1319 B.n512 B.n511 163.367
R1320 B.n508 B.n507 163.367
R1321 B.n504 B.n503 163.367
R1322 B.n500 B.n499 163.367
R1323 B.n496 B.n495 163.367
R1324 B.n492 B.n491 163.367
R1325 B.n488 B.n487 163.367
R1326 B.n484 B.n483 163.367
R1327 B.n480 B.n479 163.367
R1328 B.n476 B.n475 163.367
R1329 B.n472 B.n471 163.367
R1330 B.n468 B.n467 163.367
R1331 B.n464 B.n463 163.367
R1332 B.n460 B.n459 163.367
R1333 B.n456 B.n455 163.367
R1334 B.n452 B.n451 163.367
R1335 B.n448 B.n447 163.367
R1336 B.n444 B.n443 163.367
R1337 B.n440 B.n439 163.367
R1338 B.n436 B.n435 163.367
R1339 B.n432 B.n431 163.367
R1340 B.n428 B.n427 163.367
R1341 B.n628 B.n370 163.367
R1342 B.n632 B.n368 163.367
R1343 B.n632 B.n362 163.367
R1344 B.n640 B.n362 163.367
R1345 B.n640 B.n360 163.367
R1346 B.n644 B.n360 163.367
R1347 B.n644 B.n353 163.367
R1348 B.n652 B.n353 163.367
R1349 B.n652 B.n351 163.367
R1350 B.n656 B.n351 163.367
R1351 B.n656 B.n346 163.367
R1352 B.n664 B.n346 163.367
R1353 B.n664 B.n344 163.367
R1354 B.n668 B.n344 163.367
R1355 B.n668 B.n338 163.367
R1356 B.n676 B.n338 163.367
R1357 B.n676 B.n336 163.367
R1358 B.n680 B.n336 163.367
R1359 B.n680 B.n330 163.367
R1360 B.n688 B.n330 163.367
R1361 B.n688 B.n328 163.367
R1362 B.n692 B.n328 163.367
R1363 B.n692 B.n323 163.367
R1364 B.n701 B.n323 163.367
R1365 B.n701 B.n321 163.367
R1366 B.n706 B.n321 163.367
R1367 B.n706 B.n315 163.367
R1368 B.n714 B.n315 163.367
R1369 B.n715 B.n714 163.367
R1370 B.n715 B.n5 163.367
R1371 B.n6 B.n5 163.367
R1372 B.n7 B.n6 163.367
R1373 B.n720 B.n7 163.367
R1374 B.n720 B.n12 163.367
R1375 B.n13 B.n12 163.367
R1376 B.n14 B.n13 163.367
R1377 B.n725 B.n14 163.367
R1378 B.n725 B.n19 163.367
R1379 B.n20 B.n19 163.367
R1380 B.n21 B.n20 163.367
R1381 B.n730 B.n21 163.367
R1382 B.n730 B.n26 163.367
R1383 B.n27 B.n26 163.367
R1384 B.n28 B.n27 163.367
R1385 B.n735 B.n28 163.367
R1386 B.n735 B.n33 163.367
R1387 B.n34 B.n33 163.367
R1388 B.n35 B.n34 163.367
R1389 B.n740 B.n35 163.367
R1390 B.n740 B.n40 163.367
R1391 B.n41 B.n40 163.367
R1392 B.n42 B.n41 163.367
R1393 B.n745 B.n42 163.367
R1394 B.n745 B.n47 163.367
R1395 B.n48 B.n47 163.367
R1396 B.n49 B.n48 163.367
R1397 B.n750 B.n49 163.367
R1398 B.n750 B.n54 163.367
R1399 B.n55 B.n54 163.367
R1400 B.n117 B.n116 163.367
R1401 B.n121 B.n120 163.367
R1402 B.n125 B.n124 163.367
R1403 B.n129 B.n128 163.367
R1404 B.n133 B.n132 163.367
R1405 B.n137 B.n136 163.367
R1406 B.n141 B.n140 163.367
R1407 B.n145 B.n144 163.367
R1408 B.n149 B.n148 163.367
R1409 B.n153 B.n152 163.367
R1410 B.n157 B.n156 163.367
R1411 B.n161 B.n160 163.367
R1412 B.n165 B.n164 163.367
R1413 B.n169 B.n168 163.367
R1414 B.n173 B.n172 163.367
R1415 B.n177 B.n176 163.367
R1416 B.n181 B.n180 163.367
R1417 B.n185 B.n184 163.367
R1418 B.n189 B.n188 163.367
R1419 B.n193 B.n192 163.367
R1420 B.n197 B.n196 163.367
R1421 B.n201 B.n200 163.367
R1422 B.n205 B.n204 163.367
R1423 B.n209 B.n208 163.367
R1424 B.n213 B.n212 163.367
R1425 B.n217 B.n216 163.367
R1426 B.n221 B.n220 163.367
R1427 B.n225 B.n224 163.367
R1428 B.n229 B.n228 163.367
R1429 B.n233 B.n232 163.367
R1430 B.n237 B.n236 163.367
R1431 B.n241 B.n240 163.367
R1432 B.n245 B.n244 163.367
R1433 B.n249 B.n248 163.367
R1434 B.n253 B.n252 163.367
R1435 B.n257 B.n256 163.367
R1436 B.n261 B.n260 163.367
R1437 B.n265 B.n264 163.367
R1438 B.n269 B.n268 163.367
R1439 B.n273 B.n272 163.367
R1440 B.n277 B.n276 163.367
R1441 B.n281 B.n280 163.367
R1442 B.n285 B.n284 163.367
R1443 B.n289 B.n288 163.367
R1444 B.n293 B.n292 163.367
R1445 B.n297 B.n296 163.367
R1446 B.n301 B.n300 163.367
R1447 B.n305 B.n304 163.367
R1448 B.n309 B.n308 163.367
R1449 B.n311 B.n106 163.367
R1450 B.n627 B.n367 78.8431
R1451 B.n758 B.n757 78.8431
R1452 B.n626 B.n625 71.676
R1453 B.n620 B.n371 71.676
R1454 B.n617 B.n372 71.676
R1455 B.n613 B.n373 71.676
R1456 B.n609 B.n374 71.676
R1457 B.n605 B.n375 71.676
R1458 B.n601 B.n376 71.676
R1459 B.n597 B.n377 71.676
R1460 B.n593 B.n378 71.676
R1461 B.n589 B.n379 71.676
R1462 B.n585 B.n380 71.676
R1463 B.n581 B.n381 71.676
R1464 B.n577 B.n382 71.676
R1465 B.n573 B.n383 71.676
R1466 B.n569 B.n384 71.676
R1467 B.n565 B.n385 71.676
R1468 B.n561 B.n386 71.676
R1469 B.n557 B.n387 71.676
R1470 B.n553 B.n388 71.676
R1471 B.n549 B.n389 71.676
R1472 B.n545 B.n390 71.676
R1473 B.n541 B.n391 71.676
R1474 B.n537 B.n392 71.676
R1475 B.n532 B.n393 71.676
R1476 B.n528 B.n394 71.676
R1477 B.n524 B.n395 71.676
R1478 B.n520 B.n396 71.676
R1479 B.n516 B.n397 71.676
R1480 B.n511 B.n398 71.676
R1481 B.n507 B.n399 71.676
R1482 B.n503 B.n400 71.676
R1483 B.n499 B.n401 71.676
R1484 B.n495 B.n402 71.676
R1485 B.n491 B.n403 71.676
R1486 B.n487 B.n404 71.676
R1487 B.n483 B.n405 71.676
R1488 B.n479 B.n406 71.676
R1489 B.n475 B.n407 71.676
R1490 B.n471 B.n408 71.676
R1491 B.n467 B.n409 71.676
R1492 B.n463 B.n410 71.676
R1493 B.n459 B.n411 71.676
R1494 B.n455 B.n412 71.676
R1495 B.n451 B.n413 71.676
R1496 B.n447 B.n414 71.676
R1497 B.n443 B.n415 71.676
R1498 B.n439 B.n416 71.676
R1499 B.n435 B.n417 71.676
R1500 B.n431 B.n418 71.676
R1501 B.n427 B.n419 71.676
R1502 B.n113 B.n56 71.676
R1503 B.n117 B.n57 71.676
R1504 B.n121 B.n58 71.676
R1505 B.n125 B.n59 71.676
R1506 B.n129 B.n60 71.676
R1507 B.n133 B.n61 71.676
R1508 B.n137 B.n62 71.676
R1509 B.n141 B.n63 71.676
R1510 B.n145 B.n64 71.676
R1511 B.n149 B.n65 71.676
R1512 B.n153 B.n66 71.676
R1513 B.n157 B.n67 71.676
R1514 B.n161 B.n68 71.676
R1515 B.n165 B.n69 71.676
R1516 B.n169 B.n70 71.676
R1517 B.n173 B.n71 71.676
R1518 B.n177 B.n72 71.676
R1519 B.n181 B.n73 71.676
R1520 B.n185 B.n74 71.676
R1521 B.n189 B.n75 71.676
R1522 B.n193 B.n76 71.676
R1523 B.n197 B.n77 71.676
R1524 B.n201 B.n78 71.676
R1525 B.n205 B.n79 71.676
R1526 B.n209 B.n80 71.676
R1527 B.n213 B.n81 71.676
R1528 B.n217 B.n82 71.676
R1529 B.n221 B.n83 71.676
R1530 B.n225 B.n84 71.676
R1531 B.n229 B.n85 71.676
R1532 B.n233 B.n86 71.676
R1533 B.n237 B.n87 71.676
R1534 B.n241 B.n88 71.676
R1535 B.n245 B.n89 71.676
R1536 B.n249 B.n90 71.676
R1537 B.n253 B.n91 71.676
R1538 B.n257 B.n92 71.676
R1539 B.n261 B.n93 71.676
R1540 B.n265 B.n94 71.676
R1541 B.n269 B.n95 71.676
R1542 B.n273 B.n96 71.676
R1543 B.n277 B.n97 71.676
R1544 B.n281 B.n98 71.676
R1545 B.n285 B.n99 71.676
R1546 B.n289 B.n100 71.676
R1547 B.n293 B.n101 71.676
R1548 B.n297 B.n102 71.676
R1549 B.n301 B.n103 71.676
R1550 B.n305 B.n104 71.676
R1551 B.n309 B.n105 71.676
R1552 B.n756 B.n106 71.676
R1553 B.n756 B.n755 71.676
R1554 B.n311 B.n105 71.676
R1555 B.n308 B.n104 71.676
R1556 B.n304 B.n103 71.676
R1557 B.n300 B.n102 71.676
R1558 B.n296 B.n101 71.676
R1559 B.n292 B.n100 71.676
R1560 B.n288 B.n99 71.676
R1561 B.n284 B.n98 71.676
R1562 B.n280 B.n97 71.676
R1563 B.n276 B.n96 71.676
R1564 B.n272 B.n95 71.676
R1565 B.n268 B.n94 71.676
R1566 B.n264 B.n93 71.676
R1567 B.n260 B.n92 71.676
R1568 B.n256 B.n91 71.676
R1569 B.n252 B.n90 71.676
R1570 B.n248 B.n89 71.676
R1571 B.n244 B.n88 71.676
R1572 B.n240 B.n87 71.676
R1573 B.n236 B.n86 71.676
R1574 B.n232 B.n85 71.676
R1575 B.n228 B.n84 71.676
R1576 B.n224 B.n83 71.676
R1577 B.n220 B.n82 71.676
R1578 B.n216 B.n81 71.676
R1579 B.n212 B.n80 71.676
R1580 B.n208 B.n79 71.676
R1581 B.n204 B.n78 71.676
R1582 B.n200 B.n77 71.676
R1583 B.n196 B.n76 71.676
R1584 B.n192 B.n75 71.676
R1585 B.n188 B.n74 71.676
R1586 B.n184 B.n73 71.676
R1587 B.n180 B.n72 71.676
R1588 B.n176 B.n71 71.676
R1589 B.n172 B.n70 71.676
R1590 B.n168 B.n69 71.676
R1591 B.n164 B.n68 71.676
R1592 B.n160 B.n67 71.676
R1593 B.n156 B.n66 71.676
R1594 B.n152 B.n65 71.676
R1595 B.n148 B.n64 71.676
R1596 B.n144 B.n63 71.676
R1597 B.n140 B.n62 71.676
R1598 B.n136 B.n61 71.676
R1599 B.n132 B.n60 71.676
R1600 B.n128 B.n59 71.676
R1601 B.n124 B.n58 71.676
R1602 B.n120 B.n57 71.676
R1603 B.n116 B.n56 71.676
R1604 B.n626 B.n421 71.676
R1605 B.n618 B.n371 71.676
R1606 B.n614 B.n372 71.676
R1607 B.n610 B.n373 71.676
R1608 B.n606 B.n374 71.676
R1609 B.n602 B.n375 71.676
R1610 B.n598 B.n376 71.676
R1611 B.n594 B.n377 71.676
R1612 B.n590 B.n378 71.676
R1613 B.n586 B.n379 71.676
R1614 B.n582 B.n380 71.676
R1615 B.n578 B.n381 71.676
R1616 B.n574 B.n382 71.676
R1617 B.n570 B.n383 71.676
R1618 B.n566 B.n384 71.676
R1619 B.n562 B.n385 71.676
R1620 B.n558 B.n386 71.676
R1621 B.n554 B.n387 71.676
R1622 B.n550 B.n388 71.676
R1623 B.n546 B.n389 71.676
R1624 B.n542 B.n390 71.676
R1625 B.n538 B.n391 71.676
R1626 B.n533 B.n392 71.676
R1627 B.n529 B.n393 71.676
R1628 B.n525 B.n394 71.676
R1629 B.n521 B.n395 71.676
R1630 B.n517 B.n396 71.676
R1631 B.n512 B.n397 71.676
R1632 B.n508 B.n398 71.676
R1633 B.n504 B.n399 71.676
R1634 B.n500 B.n400 71.676
R1635 B.n496 B.n401 71.676
R1636 B.n492 B.n402 71.676
R1637 B.n488 B.n403 71.676
R1638 B.n484 B.n404 71.676
R1639 B.n480 B.n405 71.676
R1640 B.n476 B.n406 71.676
R1641 B.n472 B.n407 71.676
R1642 B.n468 B.n408 71.676
R1643 B.n464 B.n409 71.676
R1644 B.n460 B.n410 71.676
R1645 B.n456 B.n411 71.676
R1646 B.n452 B.n412 71.676
R1647 B.n448 B.n413 71.676
R1648 B.n444 B.n414 71.676
R1649 B.n440 B.n415 71.676
R1650 B.n436 B.n416 71.676
R1651 B.n432 B.n417 71.676
R1652 B.n428 B.n418 71.676
R1653 B.n419 B.n370 71.676
R1654 B.n425 B.n424 69.4308
R1655 B.n423 B.n422 69.4308
R1656 B.n111 B.n110 69.4308
R1657 B.n108 B.n107 69.4308
R1658 B.n514 B.n425 59.5399
R1659 B.n535 B.n423 59.5399
R1660 B.n112 B.n111 59.5399
R1661 B.n109 B.n108 59.5399
R1662 B.n633 B.n367 39.7138
R1663 B.n633 B.n363 39.7138
R1664 B.n639 B.n363 39.7138
R1665 B.n639 B.n359 39.7138
R1666 B.n645 B.n359 39.7138
R1667 B.n645 B.n354 39.7138
R1668 B.n651 B.n354 39.7138
R1669 B.n651 B.n355 39.7138
R1670 B.n657 B.n347 39.7138
R1671 B.n663 B.n347 39.7138
R1672 B.n663 B.n343 39.7138
R1673 B.n669 B.n343 39.7138
R1674 B.n669 B.n339 39.7138
R1675 B.n675 B.n339 39.7138
R1676 B.n675 B.n335 39.7138
R1677 B.n681 B.n335 39.7138
R1678 B.n681 B.n331 39.7138
R1679 B.n687 B.n331 39.7138
R1680 B.n687 B.n327 39.7138
R1681 B.n694 B.n327 39.7138
R1682 B.n694 B.n693 39.7138
R1683 B.n700 B.n320 39.7138
R1684 B.n707 B.n320 39.7138
R1685 B.n707 B.n316 39.7138
R1686 B.n713 B.n316 39.7138
R1687 B.n713 B.n4 39.7138
R1688 B.n815 B.n4 39.7138
R1689 B.n815 B.n814 39.7138
R1690 B.n814 B.n813 39.7138
R1691 B.n813 B.n8 39.7138
R1692 B.n807 B.n8 39.7138
R1693 B.n807 B.n806 39.7138
R1694 B.n806 B.n805 39.7138
R1695 B.n799 B.n18 39.7138
R1696 B.n799 B.n798 39.7138
R1697 B.n798 B.n797 39.7138
R1698 B.n797 B.n22 39.7138
R1699 B.n791 B.n22 39.7138
R1700 B.n791 B.n790 39.7138
R1701 B.n790 B.n789 39.7138
R1702 B.n789 B.n29 39.7138
R1703 B.n783 B.n29 39.7138
R1704 B.n783 B.n782 39.7138
R1705 B.n782 B.n781 39.7138
R1706 B.n781 B.n36 39.7138
R1707 B.n775 B.n36 39.7138
R1708 B.n774 B.n773 39.7138
R1709 B.n773 B.n43 39.7138
R1710 B.n767 B.n43 39.7138
R1711 B.n767 B.n766 39.7138
R1712 B.n766 B.n765 39.7138
R1713 B.n765 B.n50 39.7138
R1714 B.n759 B.n50 39.7138
R1715 B.n759 B.n758 39.7138
R1716 B.n700 B.t1 34.4576
R1717 B.n805 B.t0 34.4576
R1718 B.n114 B.n52 34.1859
R1719 B.n754 B.n753 34.1859
R1720 B.n630 B.n629 34.1859
R1721 B.n624 B.n365 34.1859
R1722 B.n657 B.t3 23.9453
R1723 B.n775 B.t7 23.9453
R1724 B B.n817 18.0485
R1725 B.n355 B.t3 15.769
R1726 B.t7 B.n774 15.769
R1727 B.n115 B.n114 10.6151
R1728 B.n118 B.n115 10.6151
R1729 B.n119 B.n118 10.6151
R1730 B.n122 B.n119 10.6151
R1731 B.n123 B.n122 10.6151
R1732 B.n126 B.n123 10.6151
R1733 B.n127 B.n126 10.6151
R1734 B.n130 B.n127 10.6151
R1735 B.n131 B.n130 10.6151
R1736 B.n134 B.n131 10.6151
R1737 B.n135 B.n134 10.6151
R1738 B.n138 B.n135 10.6151
R1739 B.n139 B.n138 10.6151
R1740 B.n142 B.n139 10.6151
R1741 B.n143 B.n142 10.6151
R1742 B.n146 B.n143 10.6151
R1743 B.n147 B.n146 10.6151
R1744 B.n150 B.n147 10.6151
R1745 B.n151 B.n150 10.6151
R1746 B.n154 B.n151 10.6151
R1747 B.n155 B.n154 10.6151
R1748 B.n158 B.n155 10.6151
R1749 B.n159 B.n158 10.6151
R1750 B.n162 B.n159 10.6151
R1751 B.n163 B.n162 10.6151
R1752 B.n166 B.n163 10.6151
R1753 B.n167 B.n166 10.6151
R1754 B.n170 B.n167 10.6151
R1755 B.n171 B.n170 10.6151
R1756 B.n174 B.n171 10.6151
R1757 B.n175 B.n174 10.6151
R1758 B.n178 B.n175 10.6151
R1759 B.n179 B.n178 10.6151
R1760 B.n182 B.n179 10.6151
R1761 B.n183 B.n182 10.6151
R1762 B.n186 B.n183 10.6151
R1763 B.n187 B.n186 10.6151
R1764 B.n190 B.n187 10.6151
R1765 B.n191 B.n190 10.6151
R1766 B.n194 B.n191 10.6151
R1767 B.n195 B.n194 10.6151
R1768 B.n198 B.n195 10.6151
R1769 B.n199 B.n198 10.6151
R1770 B.n202 B.n199 10.6151
R1771 B.n203 B.n202 10.6151
R1772 B.n207 B.n206 10.6151
R1773 B.n210 B.n207 10.6151
R1774 B.n211 B.n210 10.6151
R1775 B.n214 B.n211 10.6151
R1776 B.n215 B.n214 10.6151
R1777 B.n218 B.n215 10.6151
R1778 B.n219 B.n218 10.6151
R1779 B.n222 B.n219 10.6151
R1780 B.n223 B.n222 10.6151
R1781 B.n227 B.n226 10.6151
R1782 B.n230 B.n227 10.6151
R1783 B.n231 B.n230 10.6151
R1784 B.n234 B.n231 10.6151
R1785 B.n235 B.n234 10.6151
R1786 B.n238 B.n235 10.6151
R1787 B.n239 B.n238 10.6151
R1788 B.n242 B.n239 10.6151
R1789 B.n243 B.n242 10.6151
R1790 B.n246 B.n243 10.6151
R1791 B.n247 B.n246 10.6151
R1792 B.n250 B.n247 10.6151
R1793 B.n251 B.n250 10.6151
R1794 B.n254 B.n251 10.6151
R1795 B.n255 B.n254 10.6151
R1796 B.n258 B.n255 10.6151
R1797 B.n259 B.n258 10.6151
R1798 B.n262 B.n259 10.6151
R1799 B.n263 B.n262 10.6151
R1800 B.n266 B.n263 10.6151
R1801 B.n267 B.n266 10.6151
R1802 B.n270 B.n267 10.6151
R1803 B.n271 B.n270 10.6151
R1804 B.n274 B.n271 10.6151
R1805 B.n275 B.n274 10.6151
R1806 B.n278 B.n275 10.6151
R1807 B.n279 B.n278 10.6151
R1808 B.n282 B.n279 10.6151
R1809 B.n283 B.n282 10.6151
R1810 B.n286 B.n283 10.6151
R1811 B.n287 B.n286 10.6151
R1812 B.n290 B.n287 10.6151
R1813 B.n291 B.n290 10.6151
R1814 B.n294 B.n291 10.6151
R1815 B.n295 B.n294 10.6151
R1816 B.n298 B.n295 10.6151
R1817 B.n299 B.n298 10.6151
R1818 B.n302 B.n299 10.6151
R1819 B.n303 B.n302 10.6151
R1820 B.n306 B.n303 10.6151
R1821 B.n307 B.n306 10.6151
R1822 B.n310 B.n307 10.6151
R1823 B.n312 B.n310 10.6151
R1824 B.n313 B.n312 10.6151
R1825 B.n754 B.n313 10.6151
R1826 B.n631 B.n630 10.6151
R1827 B.n631 B.n361 10.6151
R1828 B.n641 B.n361 10.6151
R1829 B.n642 B.n641 10.6151
R1830 B.n643 B.n642 10.6151
R1831 B.n643 B.n352 10.6151
R1832 B.n653 B.n352 10.6151
R1833 B.n654 B.n653 10.6151
R1834 B.n655 B.n654 10.6151
R1835 B.n655 B.n345 10.6151
R1836 B.n665 B.n345 10.6151
R1837 B.n666 B.n665 10.6151
R1838 B.n667 B.n666 10.6151
R1839 B.n667 B.n337 10.6151
R1840 B.n677 B.n337 10.6151
R1841 B.n678 B.n677 10.6151
R1842 B.n679 B.n678 10.6151
R1843 B.n679 B.n329 10.6151
R1844 B.n689 B.n329 10.6151
R1845 B.n690 B.n689 10.6151
R1846 B.n691 B.n690 10.6151
R1847 B.n691 B.n322 10.6151
R1848 B.n702 B.n322 10.6151
R1849 B.n703 B.n702 10.6151
R1850 B.n705 B.n703 10.6151
R1851 B.n705 B.n704 10.6151
R1852 B.n704 B.n314 10.6151
R1853 B.n716 B.n314 10.6151
R1854 B.n717 B.n716 10.6151
R1855 B.n718 B.n717 10.6151
R1856 B.n719 B.n718 10.6151
R1857 B.n721 B.n719 10.6151
R1858 B.n722 B.n721 10.6151
R1859 B.n723 B.n722 10.6151
R1860 B.n724 B.n723 10.6151
R1861 B.n726 B.n724 10.6151
R1862 B.n727 B.n726 10.6151
R1863 B.n728 B.n727 10.6151
R1864 B.n729 B.n728 10.6151
R1865 B.n731 B.n729 10.6151
R1866 B.n732 B.n731 10.6151
R1867 B.n733 B.n732 10.6151
R1868 B.n734 B.n733 10.6151
R1869 B.n736 B.n734 10.6151
R1870 B.n737 B.n736 10.6151
R1871 B.n738 B.n737 10.6151
R1872 B.n739 B.n738 10.6151
R1873 B.n741 B.n739 10.6151
R1874 B.n742 B.n741 10.6151
R1875 B.n743 B.n742 10.6151
R1876 B.n744 B.n743 10.6151
R1877 B.n746 B.n744 10.6151
R1878 B.n747 B.n746 10.6151
R1879 B.n748 B.n747 10.6151
R1880 B.n749 B.n748 10.6151
R1881 B.n751 B.n749 10.6151
R1882 B.n752 B.n751 10.6151
R1883 B.n753 B.n752 10.6151
R1884 B.n624 B.n623 10.6151
R1885 B.n623 B.n622 10.6151
R1886 B.n622 B.n621 10.6151
R1887 B.n621 B.n619 10.6151
R1888 B.n619 B.n616 10.6151
R1889 B.n616 B.n615 10.6151
R1890 B.n615 B.n612 10.6151
R1891 B.n612 B.n611 10.6151
R1892 B.n611 B.n608 10.6151
R1893 B.n608 B.n607 10.6151
R1894 B.n607 B.n604 10.6151
R1895 B.n604 B.n603 10.6151
R1896 B.n603 B.n600 10.6151
R1897 B.n600 B.n599 10.6151
R1898 B.n599 B.n596 10.6151
R1899 B.n596 B.n595 10.6151
R1900 B.n595 B.n592 10.6151
R1901 B.n592 B.n591 10.6151
R1902 B.n591 B.n588 10.6151
R1903 B.n588 B.n587 10.6151
R1904 B.n587 B.n584 10.6151
R1905 B.n584 B.n583 10.6151
R1906 B.n583 B.n580 10.6151
R1907 B.n580 B.n579 10.6151
R1908 B.n579 B.n576 10.6151
R1909 B.n576 B.n575 10.6151
R1910 B.n575 B.n572 10.6151
R1911 B.n572 B.n571 10.6151
R1912 B.n571 B.n568 10.6151
R1913 B.n568 B.n567 10.6151
R1914 B.n567 B.n564 10.6151
R1915 B.n564 B.n563 10.6151
R1916 B.n563 B.n560 10.6151
R1917 B.n560 B.n559 10.6151
R1918 B.n559 B.n556 10.6151
R1919 B.n556 B.n555 10.6151
R1920 B.n555 B.n552 10.6151
R1921 B.n552 B.n551 10.6151
R1922 B.n551 B.n548 10.6151
R1923 B.n548 B.n547 10.6151
R1924 B.n547 B.n544 10.6151
R1925 B.n544 B.n543 10.6151
R1926 B.n543 B.n540 10.6151
R1927 B.n540 B.n539 10.6151
R1928 B.n539 B.n536 10.6151
R1929 B.n534 B.n531 10.6151
R1930 B.n531 B.n530 10.6151
R1931 B.n530 B.n527 10.6151
R1932 B.n527 B.n526 10.6151
R1933 B.n526 B.n523 10.6151
R1934 B.n523 B.n522 10.6151
R1935 B.n522 B.n519 10.6151
R1936 B.n519 B.n518 10.6151
R1937 B.n518 B.n515 10.6151
R1938 B.n513 B.n510 10.6151
R1939 B.n510 B.n509 10.6151
R1940 B.n509 B.n506 10.6151
R1941 B.n506 B.n505 10.6151
R1942 B.n505 B.n502 10.6151
R1943 B.n502 B.n501 10.6151
R1944 B.n501 B.n498 10.6151
R1945 B.n498 B.n497 10.6151
R1946 B.n497 B.n494 10.6151
R1947 B.n494 B.n493 10.6151
R1948 B.n493 B.n490 10.6151
R1949 B.n490 B.n489 10.6151
R1950 B.n489 B.n486 10.6151
R1951 B.n486 B.n485 10.6151
R1952 B.n485 B.n482 10.6151
R1953 B.n482 B.n481 10.6151
R1954 B.n481 B.n478 10.6151
R1955 B.n478 B.n477 10.6151
R1956 B.n477 B.n474 10.6151
R1957 B.n474 B.n473 10.6151
R1958 B.n473 B.n470 10.6151
R1959 B.n470 B.n469 10.6151
R1960 B.n469 B.n466 10.6151
R1961 B.n466 B.n465 10.6151
R1962 B.n465 B.n462 10.6151
R1963 B.n462 B.n461 10.6151
R1964 B.n461 B.n458 10.6151
R1965 B.n458 B.n457 10.6151
R1966 B.n457 B.n454 10.6151
R1967 B.n454 B.n453 10.6151
R1968 B.n453 B.n450 10.6151
R1969 B.n450 B.n449 10.6151
R1970 B.n449 B.n446 10.6151
R1971 B.n446 B.n445 10.6151
R1972 B.n445 B.n442 10.6151
R1973 B.n442 B.n441 10.6151
R1974 B.n441 B.n438 10.6151
R1975 B.n438 B.n437 10.6151
R1976 B.n437 B.n434 10.6151
R1977 B.n434 B.n433 10.6151
R1978 B.n433 B.n430 10.6151
R1979 B.n430 B.n429 10.6151
R1980 B.n429 B.n426 10.6151
R1981 B.n426 B.n369 10.6151
R1982 B.n629 B.n369 10.6151
R1983 B.n635 B.n365 10.6151
R1984 B.n636 B.n635 10.6151
R1985 B.n637 B.n636 10.6151
R1986 B.n637 B.n357 10.6151
R1987 B.n647 B.n357 10.6151
R1988 B.n648 B.n647 10.6151
R1989 B.n649 B.n648 10.6151
R1990 B.n649 B.n349 10.6151
R1991 B.n659 B.n349 10.6151
R1992 B.n660 B.n659 10.6151
R1993 B.n661 B.n660 10.6151
R1994 B.n661 B.n341 10.6151
R1995 B.n671 B.n341 10.6151
R1996 B.n672 B.n671 10.6151
R1997 B.n673 B.n672 10.6151
R1998 B.n673 B.n333 10.6151
R1999 B.n683 B.n333 10.6151
R2000 B.n684 B.n683 10.6151
R2001 B.n685 B.n684 10.6151
R2002 B.n685 B.n325 10.6151
R2003 B.n696 B.n325 10.6151
R2004 B.n697 B.n696 10.6151
R2005 B.n698 B.n697 10.6151
R2006 B.n698 B.n318 10.6151
R2007 B.n709 B.n318 10.6151
R2008 B.n710 B.n709 10.6151
R2009 B.n711 B.n710 10.6151
R2010 B.n711 B.n0 10.6151
R2011 B.n811 B.n1 10.6151
R2012 B.n811 B.n810 10.6151
R2013 B.n810 B.n809 10.6151
R2014 B.n809 B.n10 10.6151
R2015 B.n803 B.n10 10.6151
R2016 B.n803 B.n802 10.6151
R2017 B.n802 B.n801 10.6151
R2018 B.n801 B.n16 10.6151
R2019 B.n795 B.n16 10.6151
R2020 B.n795 B.n794 10.6151
R2021 B.n794 B.n793 10.6151
R2022 B.n793 B.n24 10.6151
R2023 B.n787 B.n24 10.6151
R2024 B.n787 B.n786 10.6151
R2025 B.n786 B.n785 10.6151
R2026 B.n785 B.n31 10.6151
R2027 B.n779 B.n31 10.6151
R2028 B.n779 B.n778 10.6151
R2029 B.n778 B.n777 10.6151
R2030 B.n777 B.n38 10.6151
R2031 B.n771 B.n38 10.6151
R2032 B.n771 B.n770 10.6151
R2033 B.n770 B.n769 10.6151
R2034 B.n769 B.n45 10.6151
R2035 B.n763 B.n45 10.6151
R2036 B.n763 B.n762 10.6151
R2037 B.n762 B.n761 10.6151
R2038 B.n761 B.n52 10.6151
R2039 B.n203 B.n112 9.36635
R2040 B.n226 B.n109 9.36635
R2041 B.n536 B.n535 9.36635
R2042 B.n514 B.n513 9.36635
R2043 B.n693 B.t1 5.25667
R2044 B.n18 B.t0 5.25667
R2045 B.n817 B.n0 2.81026
R2046 B.n817 B.n1 2.81026
R2047 B.n206 B.n112 1.24928
R2048 B.n223 B.n109 1.24928
R2049 B.n535 B.n534 1.24928
R2050 B.n515 B.n514 1.24928
R2051 VN VN.t0 186.752
R2052 VN VN.t1 139.81
R2053 VDD2.n141 VDD2.n73 289.615
R2054 VDD2.n68 VDD2.n0 289.615
R2055 VDD2.n142 VDD2.n141 185
R2056 VDD2.n140 VDD2.n139 185
R2057 VDD2.n77 VDD2.n76 185
R2058 VDD2.n134 VDD2.n133 185
R2059 VDD2.n132 VDD2.n131 185
R2060 VDD2.n81 VDD2.n80 185
R2061 VDD2.n126 VDD2.n125 185
R2062 VDD2.n124 VDD2.n123 185
R2063 VDD2.n85 VDD2.n84 185
R2064 VDD2.n89 VDD2.n87 185
R2065 VDD2.n118 VDD2.n117 185
R2066 VDD2.n116 VDD2.n115 185
R2067 VDD2.n91 VDD2.n90 185
R2068 VDD2.n110 VDD2.n109 185
R2069 VDD2.n108 VDD2.n107 185
R2070 VDD2.n95 VDD2.n94 185
R2071 VDD2.n102 VDD2.n101 185
R2072 VDD2.n100 VDD2.n99 185
R2073 VDD2.n25 VDD2.n24 185
R2074 VDD2.n27 VDD2.n26 185
R2075 VDD2.n20 VDD2.n19 185
R2076 VDD2.n33 VDD2.n32 185
R2077 VDD2.n35 VDD2.n34 185
R2078 VDD2.n16 VDD2.n15 185
R2079 VDD2.n42 VDD2.n41 185
R2080 VDD2.n43 VDD2.n14 185
R2081 VDD2.n45 VDD2.n44 185
R2082 VDD2.n12 VDD2.n11 185
R2083 VDD2.n51 VDD2.n50 185
R2084 VDD2.n53 VDD2.n52 185
R2085 VDD2.n8 VDD2.n7 185
R2086 VDD2.n59 VDD2.n58 185
R2087 VDD2.n61 VDD2.n60 185
R2088 VDD2.n4 VDD2.n3 185
R2089 VDD2.n67 VDD2.n66 185
R2090 VDD2.n69 VDD2.n68 185
R2091 VDD2.n98 VDD2.t1 149.524
R2092 VDD2.n23 VDD2.t0 149.524
R2093 VDD2.n141 VDD2.n140 104.615
R2094 VDD2.n140 VDD2.n76 104.615
R2095 VDD2.n133 VDD2.n76 104.615
R2096 VDD2.n133 VDD2.n132 104.615
R2097 VDD2.n132 VDD2.n80 104.615
R2098 VDD2.n125 VDD2.n80 104.615
R2099 VDD2.n125 VDD2.n124 104.615
R2100 VDD2.n124 VDD2.n84 104.615
R2101 VDD2.n89 VDD2.n84 104.615
R2102 VDD2.n117 VDD2.n89 104.615
R2103 VDD2.n117 VDD2.n116 104.615
R2104 VDD2.n116 VDD2.n90 104.615
R2105 VDD2.n109 VDD2.n90 104.615
R2106 VDD2.n109 VDD2.n108 104.615
R2107 VDD2.n108 VDD2.n94 104.615
R2108 VDD2.n101 VDD2.n94 104.615
R2109 VDD2.n101 VDD2.n100 104.615
R2110 VDD2.n26 VDD2.n25 104.615
R2111 VDD2.n26 VDD2.n19 104.615
R2112 VDD2.n33 VDD2.n19 104.615
R2113 VDD2.n34 VDD2.n33 104.615
R2114 VDD2.n34 VDD2.n15 104.615
R2115 VDD2.n42 VDD2.n15 104.615
R2116 VDD2.n43 VDD2.n42 104.615
R2117 VDD2.n44 VDD2.n43 104.615
R2118 VDD2.n44 VDD2.n11 104.615
R2119 VDD2.n51 VDD2.n11 104.615
R2120 VDD2.n52 VDD2.n51 104.615
R2121 VDD2.n52 VDD2.n7 104.615
R2122 VDD2.n59 VDD2.n7 104.615
R2123 VDD2.n60 VDD2.n59 104.615
R2124 VDD2.n60 VDD2.n3 104.615
R2125 VDD2.n67 VDD2.n3 104.615
R2126 VDD2.n68 VDD2.n67 104.615
R2127 VDD2.n146 VDD2.n72 90.3857
R2128 VDD2.n100 VDD2.t1 52.3082
R2129 VDD2.n25 VDD2.t0 52.3082
R2130 VDD2.n146 VDD2.n145 48.8641
R2131 VDD2.n87 VDD2.n85 13.1884
R2132 VDD2.n45 VDD2.n12 13.1884
R2133 VDD2.n123 VDD2.n122 12.8005
R2134 VDD2.n119 VDD2.n118 12.8005
R2135 VDD2.n46 VDD2.n14 12.8005
R2136 VDD2.n50 VDD2.n49 12.8005
R2137 VDD2.n126 VDD2.n83 12.0247
R2138 VDD2.n115 VDD2.n88 12.0247
R2139 VDD2.n41 VDD2.n40 12.0247
R2140 VDD2.n53 VDD2.n10 12.0247
R2141 VDD2.n127 VDD2.n81 11.249
R2142 VDD2.n114 VDD2.n91 11.249
R2143 VDD2.n39 VDD2.n16 11.249
R2144 VDD2.n54 VDD2.n8 11.249
R2145 VDD2.n131 VDD2.n130 10.4732
R2146 VDD2.n111 VDD2.n110 10.4732
R2147 VDD2.n36 VDD2.n35 10.4732
R2148 VDD2.n58 VDD2.n57 10.4732
R2149 VDD2.n99 VDD2.n98 10.2747
R2150 VDD2.n24 VDD2.n23 10.2747
R2151 VDD2.n134 VDD2.n79 9.69747
R2152 VDD2.n107 VDD2.n93 9.69747
R2153 VDD2.n32 VDD2.n18 9.69747
R2154 VDD2.n61 VDD2.n6 9.69747
R2155 VDD2.n145 VDD2.n144 9.45567
R2156 VDD2.n72 VDD2.n71 9.45567
R2157 VDD2.n97 VDD2.n96 9.3005
R2158 VDD2.n104 VDD2.n103 9.3005
R2159 VDD2.n106 VDD2.n105 9.3005
R2160 VDD2.n93 VDD2.n92 9.3005
R2161 VDD2.n112 VDD2.n111 9.3005
R2162 VDD2.n114 VDD2.n113 9.3005
R2163 VDD2.n88 VDD2.n86 9.3005
R2164 VDD2.n120 VDD2.n119 9.3005
R2165 VDD2.n144 VDD2.n143 9.3005
R2166 VDD2.n75 VDD2.n74 9.3005
R2167 VDD2.n138 VDD2.n137 9.3005
R2168 VDD2.n136 VDD2.n135 9.3005
R2169 VDD2.n79 VDD2.n78 9.3005
R2170 VDD2.n130 VDD2.n129 9.3005
R2171 VDD2.n128 VDD2.n127 9.3005
R2172 VDD2.n83 VDD2.n82 9.3005
R2173 VDD2.n122 VDD2.n121 9.3005
R2174 VDD2.n71 VDD2.n70 9.3005
R2175 VDD2.n65 VDD2.n64 9.3005
R2176 VDD2.n63 VDD2.n62 9.3005
R2177 VDD2.n6 VDD2.n5 9.3005
R2178 VDD2.n57 VDD2.n56 9.3005
R2179 VDD2.n55 VDD2.n54 9.3005
R2180 VDD2.n10 VDD2.n9 9.3005
R2181 VDD2.n49 VDD2.n48 9.3005
R2182 VDD2.n22 VDD2.n21 9.3005
R2183 VDD2.n29 VDD2.n28 9.3005
R2184 VDD2.n31 VDD2.n30 9.3005
R2185 VDD2.n18 VDD2.n17 9.3005
R2186 VDD2.n37 VDD2.n36 9.3005
R2187 VDD2.n39 VDD2.n38 9.3005
R2188 VDD2.n40 VDD2.n13 9.3005
R2189 VDD2.n47 VDD2.n46 9.3005
R2190 VDD2.n2 VDD2.n1 9.3005
R2191 VDD2.n135 VDD2.n77 8.92171
R2192 VDD2.n106 VDD2.n95 8.92171
R2193 VDD2.n31 VDD2.n20 8.92171
R2194 VDD2.n62 VDD2.n4 8.92171
R2195 VDD2.n139 VDD2.n138 8.14595
R2196 VDD2.n103 VDD2.n102 8.14595
R2197 VDD2.n28 VDD2.n27 8.14595
R2198 VDD2.n66 VDD2.n65 8.14595
R2199 VDD2.n145 VDD2.n73 7.3702
R2200 VDD2.n142 VDD2.n75 7.3702
R2201 VDD2.n99 VDD2.n97 7.3702
R2202 VDD2.n24 VDD2.n22 7.3702
R2203 VDD2.n69 VDD2.n2 7.3702
R2204 VDD2.n72 VDD2.n0 7.3702
R2205 VDD2.n143 VDD2.n73 6.59444
R2206 VDD2.n143 VDD2.n142 6.59444
R2207 VDD2.n70 VDD2.n69 6.59444
R2208 VDD2.n70 VDD2.n0 6.59444
R2209 VDD2.n139 VDD2.n75 5.81868
R2210 VDD2.n102 VDD2.n97 5.81868
R2211 VDD2.n27 VDD2.n22 5.81868
R2212 VDD2.n66 VDD2.n2 5.81868
R2213 VDD2.n138 VDD2.n77 5.04292
R2214 VDD2.n103 VDD2.n95 5.04292
R2215 VDD2.n28 VDD2.n20 5.04292
R2216 VDD2.n65 VDD2.n4 5.04292
R2217 VDD2.n135 VDD2.n134 4.26717
R2218 VDD2.n107 VDD2.n106 4.26717
R2219 VDD2.n32 VDD2.n31 4.26717
R2220 VDD2.n62 VDD2.n61 4.26717
R2221 VDD2.n131 VDD2.n79 3.49141
R2222 VDD2.n110 VDD2.n93 3.49141
R2223 VDD2.n35 VDD2.n18 3.49141
R2224 VDD2.n58 VDD2.n6 3.49141
R2225 VDD2.n98 VDD2.n96 2.84303
R2226 VDD2.n23 VDD2.n21 2.84303
R2227 VDD2.n130 VDD2.n81 2.71565
R2228 VDD2.n111 VDD2.n91 2.71565
R2229 VDD2.n36 VDD2.n16 2.71565
R2230 VDD2.n57 VDD2.n8 2.71565
R2231 VDD2.n127 VDD2.n126 1.93989
R2232 VDD2.n115 VDD2.n114 1.93989
R2233 VDD2.n41 VDD2.n39 1.93989
R2234 VDD2.n54 VDD2.n53 1.93989
R2235 VDD2.n123 VDD2.n83 1.16414
R2236 VDD2.n118 VDD2.n88 1.16414
R2237 VDD2.n40 VDD2.n14 1.16414
R2238 VDD2.n50 VDD2.n10 1.16414
R2239 VDD2 VDD2.n146 0.830241
R2240 VDD2.n122 VDD2.n85 0.388379
R2241 VDD2.n119 VDD2.n87 0.388379
R2242 VDD2.n46 VDD2.n45 0.388379
R2243 VDD2.n49 VDD2.n12 0.388379
R2244 VDD2.n144 VDD2.n74 0.155672
R2245 VDD2.n137 VDD2.n74 0.155672
R2246 VDD2.n137 VDD2.n136 0.155672
R2247 VDD2.n136 VDD2.n78 0.155672
R2248 VDD2.n129 VDD2.n78 0.155672
R2249 VDD2.n129 VDD2.n128 0.155672
R2250 VDD2.n128 VDD2.n82 0.155672
R2251 VDD2.n121 VDD2.n82 0.155672
R2252 VDD2.n121 VDD2.n120 0.155672
R2253 VDD2.n120 VDD2.n86 0.155672
R2254 VDD2.n113 VDD2.n86 0.155672
R2255 VDD2.n113 VDD2.n112 0.155672
R2256 VDD2.n112 VDD2.n92 0.155672
R2257 VDD2.n105 VDD2.n92 0.155672
R2258 VDD2.n105 VDD2.n104 0.155672
R2259 VDD2.n104 VDD2.n96 0.155672
R2260 VDD2.n29 VDD2.n21 0.155672
R2261 VDD2.n30 VDD2.n29 0.155672
R2262 VDD2.n30 VDD2.n17 0.155672
R2263 VDD2.n37 VDD2.n17 0.155672
R2264 VDD2.n38 VDD2.n37 0.155672
R2265 VDD2.n38 VDD2.n13 0.155672
R2266 VDD2.n47 VDD2.n13 0.155672
R2267 VDD2.n48 VDD2.n47 0.155672
R2268 VDD2.n48 VDD2.n9 0.155672
R2269 VDD2.n55 VDD2.n9 0.155672
R2270 VDD2.n56 VDD2.n55 0.155672
R2271 VDD2.n56 VDD2.n5 0.155672
R2272 VDD2.n63 VDD2.n5 0.155672
R2273 VDD2.n64 VDD2.n63 0.155672
R2274 VDD2.n64 VDD2.n1 0.155672
R2275 VDD2.n71 VDD2.n1 0.155672
C0 VDD1 VN 0.148086f
C1 VDD1 VDD2 0.753933f
C2 VN VP 6.05577f
C3 VP VDD2 0.36014f
C4 VDD1 VTAIL 5.58118f
C5 VP VTAIL 2.85952f
C6 VN VDD2 3.20774f
C7 VN VTAIL 2.84526f
C8 VDD2 VTAIL 5.63645f
C9 VDD1 VP 3.41731f
C10 VDD2 B 4.935604f
C11 VDD1 B 7.91566f
C12 VTAIL B 8.314223f
C13 VN B 11.72269f
C14 VP B 7.319036f
C15 VDD2.n0 B 0.029405f
C16 VDD2.n1 B 0.020146f
C17 VDD2.n2 B 0.010826f
C18 VDD2.n3 B 0.025588f
C19 VDD2.n4 B 0.011462f
C20 VDD2.n5 B 0.020146f
C21 VDD2.n6 B 0.010826f
C22 VDD2.n7 B 0.025588f
C23 VDD2.n8 B 0.011462f
C24 VDD2.n9 B 0.020146f
C25 VDD2.n10 B 0.010826f
C26 VDD2.n11 B 0.025588f
C27 VDD2.n12 B 0.011144f
C28 VDD2.n13 B 0.020146f
C29 VDD2.n14 B 0.011462f
C30 VDD2.n15 B 0.025588f
C31 VDD2.n16 B 0.011462f
C32 VDD2.n17 B 0.020146f
C33 VDD2.n18 B 0.010826f
C34 VDD2.n19 B 0.025588f
C35 VDD2.n20 B 0.011462f
C36 VDD2.n21 B 1.15612f
C37 VDD2.n22 B 0.010826f
C38 VDD2.t0 B 0.043385f
C39 VDD2.n23 B 0.157317f
C40 VDD2.n24 B 0.018089f
C41 VDD2.n25 B 0.019191f
C42 VDD2.n26 B 0.025588f
C43 VDD2.n27 B 0.011462f
C44 VDD2.n28 B 0.010826f
C45 VDD2.n29 B 0.020146f
C46 VDD2.n30 B 0.020146f
C47 VDD2.n31 B 0.010826f
C48 VDD2.n32 B 0.011462f
C49 VDD2.n33 B 0.025588f
C50 VDD2.n34 B 0.025588f
C51 VDD2.n35 B 0.011462f
C52 VDD2.n36 B 0.010826f
C53 VDD2.n37 B 0.020146f
C54 VDD2.n38 B 0.020146f
C55 VDD2.n39 B 0.010826f
C56 VDD2.n40 B 0.010826f
C57 VDD2.n41 B 0.011462f
C58 VDD2.n42 B 0.025588f
C59 VDD2.n43 B 0.025588f
C60 VDD2.n44 B 0.025588f
C61 VDD2.n45 B 0.011144f
C62 VDD2.n46 B 0.010826f
C63 VDD2.n47 B 0.020146f
C64 VDD2.n48 B 0.020146f
C65 VDD2.n49 B 0.010826f
C66 VDD2.n50 B 0.011462f
C67 VDD2.n51 B 0.025588f
C68 VDD2.n52 B 0.025588f
C69 VDD2.n53 B 0.011462f
C70 VDD2.n54 B 0.010826f
C71 VDD2.n55 B 0.020146f
C72 VDD2.n56 B 0.020146f
C73 VDD2.n57 B 0.010826f
C74 VDD2.n58 B 0.011462f
C75 VDD2.n59 B 0.025588f
C76 VDD2.n60 B 0.025588f
C77 VDD2.n61 B 0.011462f
C78 VDD2.n62 B 0.010826f
C79 VDD2.n63 B 0.020146f
C80 VDD2.n64 B 0.020146f
C81 VDD2.n65 B 0.010826f
C82 VDD2.n66 B 0.011462f
C83 VDD2.n67 B 0.025588f
C84 VDD2.n68 B 0.057316f
C85 VDD2.n69 B 0.011462f
C86 VDD2.n70 B 0.010826f
C87 VDD2.n71 B 0.046567f
C88 VDD2.n72 B 0.674258f
C89 VDD2.n73 B 0.029405f
C90 VDD2.n74 B 0.020146f
C91 VDD2.n75 B 0.010826f
C92 VDD2.n76 B 0.025588f
C93 VDD2.n77 B 0.011462f
C94 VDD2.n78 B 0.020146f
C95 VDD2.n79 B 0.010826f
C96 VDD2.n80 B 0.025588f
C97 VDD2.n81 B 0.011462f
C98 VDD2.n82 B 0.020146f
C99 VDD2.n83 B 0.010826f
C100 VDD2.n84 B 0.025588f
C101 VDD2.n85 B 0.011144f
C102 VDD2.n86 B 0.020146f
C103 VDD2.n87 B 0.011144f
C104 VDD2.n88 B 0.010826f
C105 VDD2.n89 B 0.025588f
C106 VDD2.n90 B 0.025588f
C107 VDD2.n91 B 0.011462f
C108 VDD2.n92 B 0.020146f
C109 VDD2.n93 B 0.010826f
C110 VDD2.n94 B 0.025588f
C111 VDD2.n95 B 0.011462f
C112 VDD2.n96 B 1.15612f
C113 VDD2.n97 B 0.010826f
C114 VDD2.t1 B 0.043385f
C115 VDD2.n98 B 0.157317f
C116 VDD2.n99 B 0.018089f
C117 VDD2.n100 B 0.019191f
C118 VDD2.n101 B 0.025588f
C119 VDD2.n102 B 0.011462f
C120 VDD2.n103 B 0.010826f
C121 VDD2.n104 B 0.020146f
C122 VDD2.n105 B 0.020146f
C123 VDD2.n106 B 0.010826f
C124 VDD2.n107 B 0.011462f
C125 VDD2.n108 B 0.025588f
C126 VDD2.n109 B 0.025588f
C127 VDD2.n110 B 0.011462f
C128 VDD2.n111 B 0.010826f
C129 VDD2.n112 B 0.020146f
C130 VDD2.n113 B 0.020146f
C131 VDD2.n114 B 0.010826f
C132 VDD2.n115 B 0.011462f
C133 VDD2.n116 B 0.025588f
C134 VDD2.n117 B 0.025588f
C135 VDD2.n118 B 0.011462f
C136 VDD2.n119 B 0.010826f
C137 VDD2.n120 B 0.020146f
C138 VDD2.n121 B 0.020146f
C139 VDD2.n122 B 0.010826f
C140 VDD2.n123 B 0.011462f
C141 VDD2.n124 B 0.025588f
C142 VDD2.n125 B 0.025588f
C143 VDD2.n126 B 0.011462f
C144 VDD2.n127 B 0.010826f
C145 VDD2.n128 B 0.020146f
C146 VDD2.n129 B 0.020146f
C147 VDD2.n130 B 0.010826f
C148 VDD2.n131 B 0.011462f
C149 VDD2.n132 B 0.025588f
C150 VDD2.n133 B 0.025588f
C151 VDD2.n134 B 0.011462f
C152 VDD2.n135 B 0.010826f
C153 VDD2.n136 B 0.020146f
C154 VDD2.n137 B 0.020146f
C155 VDD2.n138 B 0.010826f
C156 VDD2.n139 B 0.011462f
C157 VDD2.n140 B 0.025588f
C158 VDD2.n141 B 0.057316f
C159 VDD2.n142 B 0.011462f
C160 VDD2.n143 B 0.010826f
C161 VDD2.n144 B 0.046567f
C162 VDD2.n145 B 0.046179f
C163 VDD2.n146 B 2.69046f
C164 VN.t1 B 3.55331f
C165 VN.t0 B 4.17836f
C166 VDD1.n0 B 0.029821f
C167 VDD1.n1 B 0.020431f
C168 VDD1.n2 B 0.010979f
C169 VDD1.n3 B 0.02595f
C170 VDD1.n4 B 0.011625f
C171 VDD1.n5 B 0.020431f
C172 VDD1.n6 B 0.010979f
C173 VDD1.n7 B 0.02595f
C174 VDD1.n8 B 0.011625f
C175 VDD1.n9 B 0.020431f
C176 VDD1.n10 B 0.010979f
C177 VDD1.n11 B 0.02595f
C178 VDD1.n12 B 0.011302f
C179 VDD1.n13 B 0.020431f
C180 VDD1.n14 B 0.011302f
C181 VDD1.n15 B 0.010979f
C182 VDD1.n16 B 0.02595f
C183 VDD1.n17 B 0.02595f
C184 VDD1.n18 B 0.011625f
C185 VDD1.n19 B 0.020431f
C186 VDD1.n20 B 0.010979f
C187 VDD1.n21 B 0.02595f
C188 VDD1.n22 B 0.011625f
C189 VDD1.n23 B 1.17249f
C190 VDD1.n24 B 0.010979f
C191 VDD1.t0 B 0.043999f
C192 VDD1.n25 B 0.159543f
C193 VDD1.n26 B 0.018345f
C194 VDD1.n27 B 0.019462f
C195 VDD1.n28 B 0.02595f
C196 VDD1.n29 B 0.011625f
C197 VDD1.n30 B 0.010979f
C198 VDD1.n31 B 0.020431f
C199 VDD1.n32 B 0.020431f
C200 VDD1.n33 B 0.010979f
C201 VDD1.n34 B 0.011625f
C202 VDD1.n35 B 0.02595f
C203 VDD1.n36 B 0.02595f
C204 VDD1.n37 B 0.011625f
C205 VDD1.n38 B 0.010979f
C206 VDD1.n39 B 0.020431f
C207 VDD1.n40 B 0.020431f
C208 VDD1.n41 B 0.010979f
C209 VDD1.n42 B 0.011625f
C210 VDD1.n43 B 0.02595f
C211 VDD1.n44 B 0.02595f
C212 VDD1.n45 B 0.011625f
C213 VDD1.n46 B 0.010979f
C214 VDD1.n47 B 0.020431f
C215 VDD1.n48 B 0.020431f
C216 VDD1.n49 B 0.010979f
C217 VDD1.n50 B 0.011625f
C218 VDD1.n51 B 0.02595f
C219 VDD1.n52 B 0.02595f
C220 VDD1.n53 B 0.011625f
C221 VDD1.n54 B 0.010979f
C222 VDD1.n55 B 0.020431f
C223 VDD1.n56 B 0.020431f
C224 VDD1.n57 B 0.010979f
C225 VDD1.n58 B 0.011625f
C226 VDD1.n59 B 0.02595f
C227 VDD1.n60 B 0.02595f
C228 VDD1.n61 B 0.011625f
C229 VDD1.n62 B 0.010979f
C230 VDD1.n63 B 0.020431f
C231 VDD1.n64 B 0.020431f
C232 VDD1.n65 B 0.010979f
C233 VDD1.n66 B 0.011625f
C234 VDD1.n67 B 0.02595f
C235 VDD1.n68 B 0.058128f
C236 VDD1.n69 B 0.011625f
C237 VDD1.n70 B 0.010979f
C238 VDD1.n71 B 0.047226f
C239 VDD1.n72 B 0.048401f
C240 VDD1.n73 B 0.029821f
C241 VDD1.n74 B 0.020431f
C242 VDD1.n75 B 0.010979f
C243 VDD1.n76 B 0.02595f
C244 VDD1.n77 B 0.011625f
C245 VDD1.n78 B 0.020431f
C246 VDD1.n79 B 0.010979f
C247 VDD1.n80 B 0.02595f
C248 VDD1.n81 B 0.011625f
C249 VDD1.n82 B 0.020431f
C250 VDD1.n83 B 0.010979f
C251 VDD1.n84 B 0.02595f
C252 VDD1.n85 B 0.011302f
C253 VDD1.n86 B 0.020431f
C254 VDD1.n87 B 0.011625f
C255 VDD1.n88 B 0.02595f
C256 VDD1.n89 B 0.011625f
C257 VDD1.n90 B 0.020431f
C258 VDD1.n91 B 0.010979f
C259 VDD1.n92 B 0.02595f
C260 VDD1.n93 B 0.011625f
C261 VDD1.n94 B 1.17249f
C262 VDD1.n95 B 0.010979f
C263 VDD1.t1 B 0.043999f
C264 VDD1.n96 B 0.159543f
C265 VDD1.n97 B 0.018345f
C266 VDD1.n98 B 0.019462f
C267 VDD1.n99 B 0.02595f
C268 VDD1.n100 B 0.011625f
C269 VDD1.n101 B 0.010979f
C270 VDD1.n102 B 0.020431f
C271 VDD1.n103 B 0.020431f
C272 VDD1.n104 B 0.010979f
C273 VDD1.n105 B 0.011625f
C274 VDD1.n106 B 0.02595f
C275 VDD1.n107 B 0.02595f
C276 VDD1.n108 B 0.011625f
C277 VDD1.n109 B 0.010979f
C278 VDD1.n110 B 0.020431f
C279 VDD1.n111 B 0.020431f
C280 VDD1.n112 B 0.010979f
C281 VDD1.n113 B 0.010979f
C282 VDD1.n114 B 0.011625f
C283 VDD1.n115 B 0.02595f
C284 VDD1.n116 B 0.02595f
C285 VDD1.n117 B 0.02595f
C286 VDD1.n118 B 0.011302f
C287 VDD1.n119 B 0.010979f
C288 VDD1.n120 B 0.020431f
C289 VDD1.n121 B 0.020431f
C290 VDD1.n122 B 0.010979f
C291 VDD1.n123 B 0.011625f
C292 VDD1.n124 B 0.02595f
C293 VDD1.n125 B 0.02595f
C294 VDD1.n126 B 0.011625f
C295 VDD1.n127 B 0.010979f
C296 VDD1.n128 B 0.020431f
C297 VDD1.n129 B 0.020431f
C298 VDD1.n130 B 0.010979f
C299 VDD1.n131 B 0.011625f
C300 VDD1.n132 B 0.02595f
C301 VDD1.n133 B 0.02595f
C302 VDD1.n134 B 0.011625f
C303 VDD1.n135 B 0.010979f
C304 VDD1.n136 B 0.020431f
C305 VDD1.n137 B 0.020431f
C306 VDD1.n138 B 0.010979f
C307 VDD1.n139 B 0.011625f
C308 VDD1.n140 B 0.02595f
C309 VDD1.n141 B 0.058128f
C310 VDD1.n142 B 0.011625f
C311 VDD1.n143 B 0.010979f
C312 VDD1.n144 B 0.047226f
C313 VDD1.n145 B 0.729835f
C314 VTAIL.n0 B 0.030078f
C315 VTAIL.n1 B 0.020607f
C316 VTAIL.n2 B 0.011074f
C317 VTAIL.n3 B 0.026174f
C318 VTAIL.n4 B 0.011725f
C319 VTAIL.n5 B 0.020607f
C320 VTAIL.n6 B 0.011074f
C321 VTAIL.n7 B 0.026174f
C322 VTAIL.n8 B 0.011725f
C323 VTAIL.n9 B 0.020607f
C324 VTAIL.n10 B 0.011074f
C325 VTAIL.n11 B 0.026174f
C326 VTAIL.n12 B 0.011399f
C327 VTAIL.n13 B 0.020607f
C328 VTAIL.n14 B 0.011725f
C329 VTAIL.n15 B 0.026174f
C330 VTAIL.n16 B 0.011725f
C331 VTAIL.n17 B 0.020607f
C332 VTAIL.n18 B 0.011074f
C333 VTAIL.n19 B 0.026174f
C334 VTAIL.n20 B 0.011725f
C335 VTAIL.n21 B 1.1826f
C336 VTAIL.n22 B 0.011074f
C337 VTAIL.t1 B 0.044379f
C338 VTAIL.n23 B 0.16092f
C339 VTAIL.n24 B 0.018503f
C340 VTAIL.n25 B 0.01963f
C341 VTAIL.n26 B 0.026174f
C342 VTAIL.n27 B 0.011725f
C343 VTAIL.n28 B 0.011074f
C344 VTAIL.n29 B 0.020607f
C345 VTAIL.n30 B 0.020607f
C346 VTAIL.n31 B 0.011074f
C347 VTAIL.n32 B 0.011725f
C348 VTAIL.n33 B 0.026174f
C349 VTAIL.n34 B 0.026174f
C350 VTAIL.n35 B 0.011725f
C351 VTAIL.n36 B 0.011074f
C352 VTAIL.n37 B 0.020607f
C353 VTAIL.n38 B 0.020607f
C354 VTAIL.n39 B 0.011074f
C355 VTAIL.n40 B 0.011074f
C356 VTAIL.n41 B 0.011725f
C357 VTAIL.n42 B 0.026174f
C358 VTAIL.n43 B 0.026174f
C359 VTAIL.n44 B 0.026174f
C360 VTAIL.n45 B 0.011399f
C361 VTAIL.n46 B 0.011074f
C362 VTAIL.n47 B 0.020607f
C363 VTAIL.n48 B 0.020607f
C364 VTAIL.n49 B 0.011074f
C365 VTAIL.n50 B 0.011725f
C366 VTAIL.n51 B 0.026174f
C367 VTAIL.n52 B 0.026174f
C368 VTAIL.n53 B 0.011725f
C369 VTAIL.n54 B 0.011074f
C370 VTAIL.n55 B 0.020607f
C371 VTAIL.n56 B 0.020607f
C372 VTAIL.n57 B 0.011074f
C373 VTAIL.n58 B 0.011725f
C374 VTAIL.n59 B 0.026174f
C375 VTAIL.n60 B 0.026174f
C376 VTAIL.n61 B 0.011725f
C377 VTAIL.n62 B 0.011074f
C378 VTAIL.n63 B 0.020607f
C379 VTAIL.n64 B 0.020607f
C380 VTAIL.n65 B 0.011074f
C381 VTAIL.n66 B 0.011725f
C382 VTAIL.n67 B 0.026174f
C383 VTAIL.n68 B 0.058629f
C384 VTAIL.n69 B 0.011725f
C385 VTAIL.n70 B 0.011074f
C386 VTAIL.n71 B 0.047633f
C387 VTAIL.n72 B 0.033007f
C388 VTAIL.n73 B 1.5699f
C389 VTAIL.n74 B 0.030078f
C390 VTAIL.n75 B 0.020607f
C391 VTAIL.n76 B 0.011074f
C392 VTAIL.n77 B 0.026174f
C393 VTAIL.n78 B 0.011725f
C394 VTAIL.n79 B 0.020607f
C395 VTAIL.n80 B 0.011074f
C396 VTAIL.n81 B 0.026174f
C397 VTAIL.n82 B 0.011725f
C398 VTAIL.n83 B 0.020607f
C399 VTAIL.n84 B 0.011074f
C400 VTAIL.n85 B 0.026174f
C401 VTAIL.n86 B 0.011399f
C402 VTAIL.n87 B 0.020607f
C403 VTAIL.n88 B 0.011399f
C404 VTAIL.n89 B 0.011074f
C405 VTAIL.n90 B 0.026174f
C406 VTAIL.n91 B 0.026174f
C407 VTAIL.n92 B 0.011725f
C408 VTAIL.n93 B 0.020607f
C409 VTAIL.n94 B 0.011074f
C410 VTAIL.n95 B 0.026174f
C411 VTAIL.n96 B 0.011725f
C412 VTAIL.n97 B 1.1826f
C413 VTAIL.n98 B 0.011074f
C414 VTAIL.t3 B 0.044379f
C415 VTAIL.n99 B 0.16092f
C416 VTAIL.n100 B 0.018503f
C417 VTAIL.n101 B 0.01963f
C418 VTAIL.n102 B 0.026174f
C419 VTAIL.n103 B 0.011725f
C420 VTAIL.n104 B 0.011074f
C421 VTAIL.n105 B 0.020607f
C422 VTAIL.n106 B 0.020607f
C423 VTAIL.n107 B 0.011074f
C424 VTAIL.n108 B 0.011725f
C425 VTAIL.n109 B 0.026174f
C426 VTAIL.n110 B 0.026174f
C427 VTAIL.n111 B 0.011725f
C428 VTAIL.n112 B 0.011074f
C429 VTAIL.n113 B 0.020607f
C430 VTAIL.n114 B 0.020607f
C431 VTAIL.n115 B 0.011074f
C432 VTAIL.n116 B 0.011725f
C433 VTAIL.n117 B 0.026174f
C434 VTAIL.n118 B 0.026174f
C435 VTAIL.n119 B 0.011725f
C436 VTAIL.n120 B 0.011074f
C437 VTAIL.n121 B 0.020607f
C438 VTAIL.n122 B 0.020607f
C439 VTAIL.n123 B 0.011074f
C440 VTAIL.n124 B 0.011725f
C441 VTAIL.n125 B 0.026174f
C442 VTAIL.n126 B 0.026174f
C443 VTAIL.n127 B 0.011725f
C444 VTAIL.n128 B 0.011074f
C445 VTAIL.n129 B 0.020607f
C446 VTAIL.n130 B 0.020607f
C447 VTAIL.n131 B 0.011074f
C448 VTAIL.n132 B 0.011725f
C449 VTAIL.n133 B 0.026174f
C450 VTAIL.n134 B 0.026174f
C451 VTAIL.n135 B 0.011725f
C452 VTAIL.n136 B 0.011074f
C453 VTAIL.n137 B 0.020607f
C454 VTAIL.n138 B 0.020607f
C455 VTAIL.n139 B 0.011074f
C456 VTAIL.n140 B 0.011725f
C457 VTAIL.n141 B 0.026174f
C458 VTAIL.n142 B 0.058629f
C459 VTAIL.n143 B 0.011725f
C460 VTAIL.n144 B 0.011074f
C461 VTAIL.n145 B 0.047633f
C462 VTAIL.n146 B 0.033007f
C463 VTAIL.n147 B 1.61727f
C464 VTAIL.n148 B 0.030078f
C465 VTAIL.n149 B 0.020607f
C466 VTAIL.n150 B 0.011074f
C467 VTAIL.n151 B 0.026174f
C468 VTAIL.n152 B 0.011725f
C469 VTAIL.n153 B 0.020607f
C470 VTAIL.n154 B 0.011074f
C471 VTAIL.n155 B 0.026174f
C472 VTAIL.n156 B 0.011725f
C473 VTAIL.n157 B 0.020607f
C474 VTAIL.n158 B 0.011074f
C475 VTAIL.n159 B 0.026174f
C476 VTAIL.n160 B 0.011399f
C477 VTAIL.n161 B 0.020607f
C478 VTAIL.n162 B 0.011399f
C479 VTAIL.n163 B 0.011074f
C480 VTAIL.n164 B 0.026174f
C481 VTAIL.n165 B 0.026174f
C482 VTAIL.n166 B 0.011725f
C483 VTAIL.n167 B 0.020607f
C484 VTAIL.n168 B 0.011074f
C485 VTAIL.n169 B 0.026174f
C486 VTAIL.n170 B 0.011725f
C487 VTAIL.n171 B 1.1826f
C488 VTAIL.n172 B 0.011074f
C489 VTAIL.t2 B 0.044379f
C490 VTAIL.n173 B 0.16092f
C491 VTAIL.n174 B 0.018503f
C492 VTAIL.n175 B 0.01963f
C493 VTAIL.n176 B 0.026174f
C494 VTAIL.n177 B 0.011725f
C495 VTAIL.n178 B 0.011074f
C496 VTAIL.n179 B 0.020607f
C497 VTAIL.n180 B 0.020607f
C498 VTAIL.n181 B 0.011074f
C499 VTAIL.n182 B 0.011725f
C500 VTAIL.n183 B 0.026174f
C501 VTAIL.n184 B 0.026174f
C502 VTAIL.n185 B 0.011725f
C503 VTAIL.n186 B 0.011074f
C504 VTAIL.n187 B 0.020607f
C505 VTAIL.n188 B 0.020607f
C506 VTAIL.n189 B 0.011074f
C507 VTAIL.n190 B 0.011725f
C508 VTAIL.n191 B 0.026174f
C509 VTAIL.n192 B 0.026174f
C510 VTAIL.n193 B 0.011725f
C511 VTAIL.n194 B 0.011074f
C512 VTAIL.n195 B 0.020607f
C513 VTAIL.n196 B 0.020607f
C514 VTAIL.n197 B 0.011074f
C515 VTAIL.n198 B 0.011725f
C516 VTAIL.n199 B 0.026174f
C517 VTAIL.n200 B 0.026174f
C518 VTAIL.n201 B 0.011725f
C519 VTAIL.n202 B 0.011074f
C520 VTAIL.n203 B 0.020607f
C521 VTAIL.n204 B 0.020607f
C522 VTAIL.n205 B 0.011074f
C523 VTAIL.n206 B 0.011725f
C524 VTAIL.n207 B 0.026174f
C525 VTAIL.n208 B 0.026174f
C526 VTAIL.n209 B 0.011725f
C527 VTAIL.n210 B 0.011074f
C528 VTAIL.n211 B 0.020607f
C529 VTAIL.n212 B 0.020607f
C530 VTAIL.n213 B 0.011074f
C531 VTAIL.n214 B 0.011725f
C532 VTAIL.n215 B 0.026174f
C533 VTAIL.n216 B 0.058629f
C534 VTAIL.n217 B 0.011725f
C535 VTAIL.n218 B 0.011074f
C536 VTAIL.n219 B 0.047633f
C537 VTAIL.n220 B 0.033007f
C538 VTAIL.n221 B 1.41234f
C539 VTAIL.n222 B 0.030078f
C540 VTAIL.n223 B 0.020607f
C541 VTAIL.n224 B 0.011074f
C542 VTAIL.n225 B 0.026174f
C543 VTAIL.n226 B 0.011725f
C544 VTAIL.n227 B 0.020607f
C545 VTAIL.n228 B 0.011074f
C546 VTAIL.n229 B 0.026174f
C547 VTAIL.n230 B 0.011725f
C548 VTAIL.n231 B 0.020607f
C549 VTAIL.n232 B 0.011074f
C550 VTAIL.n233 B 0.026174f
C551 VTAIL.n234 B 0.011399f
C552 VTAIL.n235 B 0.020607f
C553 VTAIL.n236 B 0.011725f
C554 VTAIL.n237 B 0.026174f
C555 VTAIL.n238 B 0.011725f
C556 VTAIL.n239 B 0.020607f
C557 VTAIL.n240 B 0.011074f
C558 VTAIL.n241 B 0.026174f
C559 VTAIL.n242 B 0.011725f
C560 VTAIL.n243 B 1.1826f
C561 VTAIL.n244 B 0.011074f
C562 VTAIL.t0 B 0.044379f
C563 VTAIL.n245 B 0.16092f
C564 VTAIL.n246 B 0.018503f
C565 VTAIL.n247 B 0.01963f
C566 VTAIL.n248 B 0.026174f
C567 VTAIL.n249 B 0.011725f
C568 VTAIL.n250 B 0.011074f
C569 VTAIL.n251 B 0.020607f
C570 VTAIL.n252 B 0.020607f
C571 VTAIL.n253 B 0.011074f
C572 VTAIL.n254 B 0.011725f
C573 VTAIL.n255 B 0.026174f
C574 VTAIL.n256 B 0.026174f
C575 VTAIL.n257 B 0.011725f
C576 VTAIL.n258 B 0.011074f
C577 VTAIL.n259 B 0.020607f
C578 VTAIL.n260 B 0.020607f
C579 VTAIL.n261 B 0.011074f
C580 VTAIL.n262 B 0.011074f
C581 VTAIL.n263 B 0.011725f
C582 VTAIL.n264 B 0.026174f
C583 VTAIL.n265 B 0.026174f
C584 VTAIL.n266 B 0.026174f
C585 VTAIL.n267 B 0.011399f
C586 VTAIL.n268 B 0.011074f
C587 VTAIL.n269 B 0.020607f
C588 VTAIL.n270 B 0.020607f
C589 VTAIL.n271 B 0.011074f
C590 VTAIL.n272 B 0.011725f
C591 VTAIL.n273 B 0.026174f
C592 VTAIL.n274 B 0.026174f
C593 VTAIL.n275 B 0.011725f
C594 VTAIL.n276 B 0.011074f
C595 VTAIL.n277 B 0.020607f
C596 VTAIL.n278 B 0.020607f
C597 VTAIL.n279 B 0.011074f
C598 VTAIL.n280 B 0.011725f
C599 VTAIL.n281 B 0.026174f
C600 VTAIL.n282 B 0.026174f
C601 VTAIL.n283 B 0.011725f
C602 VTAIL.n284 B 0.011074f
C603 VTAIL.n285 B 0.020607f
C604 VTAIL.n286 B 0.020607f
C605 VTAIL.n287 B 0.011074f
C606 VTAIL.n288 B 0.011725f
C607 VTAIL.n289 B 0.026174f
C608 VTAIL.n290 B 0.058629f
C609 VTAIL.n291 B 0.011725f
C610 VTAIL.n292 B 0.011074f
C611 VTAIL.n293 B 0.047633f
C612 VTAIL.n294 B 0.033007f
C613 VTAIL.n295 B 1.32604f
C614 VP.t1 B 4.29524f
C615 VP.t0 B 3.64829f
C616 VP.n0 B 4.36293f
.ends

