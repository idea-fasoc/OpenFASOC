* NGSPICE file created from diff_pair_sample_0238.ext - technology: sky130A

.subckt diff_pair_sample_0238 VTAIL VN VP B VDD2 VDD1
X0 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=2.886 pd=15.58 as=0 ps=0 w=7.4 l=0.43
X1 VDD2.t5 VN.t0 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=2.886 pd=15.58 as=1.221 ps=7.73 w=7.4 l=0.43
X2 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=2.886 pd=15.58 as=0 ps=0 w=7.4 l=0.43
X3 B.t11 B.t9 B.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=2.886 pd=15.58 as=0 ps=0 w=7.4 l=0.43
X4 VTAIL.t8 VN.t1 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.221 pd=7.73 as=1.221 ps=7.73 w=7.4 l=0.43
X5 VDD1.t5 VP.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.221 pd=7.73 as=2.886 ps=15.58 w=7.4 l=0.43
X6 VTAIL.t5 VP.t1 VDD1.t4 B.t19 sky130_fd_pr__nfet_01v8 ad=1.221 pd=7.73 as=1.221 ps=7.73 w=7.4 l=0.43
X7 VDD2.t3 VN.t2 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.221 pd=7.73 as=2.886 ps=15.58 w=7.4 l=0.43
X8 VTAIL.t11 VN.t3 VDD2.t2 B.t19 sky130_fd_pr__nfet_01v8 ad=1.221 pd=7.73 as=1.221 ps=7.73 w=7.4 l=0.43
X9 VDD2.t1 VN.t4 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=2.886 pd=15.58 as=1.221 ps=7.73 w=7.4 l=0.43
X10 VDD1.t3 VP.t2 VTAIL.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.221 pd=7.73 as=2.886 ps=15.58 w=7.4 l=0.43
X11 VTAIL.t2 VP.t3 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=1.221 pd=7.73 as=1.221 ps=7.73 w=7.4 l=0.43
X12 VDD2.t0 VN.t5 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=1.221 pd=7.73 as=2.886 ps=15.58 w=7.4 l=0.43
X13 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=2.886 pd=15.58 as=0 ps=0 w=7.4 l=0.43
X14 VDD1.t1 VP.t4 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.886 pd=15.58 as=1.221 ps=7.73 w=7.4 l=0.43
X15 VDD1.t0 VP.t5 VTAIL.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.886 pd=15.58 as=1.221 ps=7.73 w=7.4 l=0.43
R0 B.n271 B.t12 623.114
R1 B.n269 B.t16 623.114
R2 B.n71 B.t9 623.114
R3 B.n68 B.t5 623.114
R4 B.n479 B.n478 585
R5 B.n202 B.n67 585
R6 B.n201 B.n200 585
R7 B.n199 B.n198 585
R8 B.n197 B.n196 585
R9 B.n195 B.n194 585
R10 B.n193 B.n192 585
R11 B.n191 B.n190 585
R12 B.n189 B.n188 585
R13 B.n187 B.n186 585
R14 B.n185 B.n184 585
R15 B.n183 B.n182 585
R16 B.n181 B.n180 585
R17 B.n179 B.n178 585
R18 B.n177 B.n176 585
R19 B.n175 B.n174 585
R20 B.n173 B.n172 585
R21 B.n171 B.n170 585
R22 B.n169 B.n168 585
R23 B.n167 B.n166 585
R24 B.n165 B.n164 585
R25 B.n163 B.n162 585
R26 B.n161 B.n160 585
R27 B.n159 B.n158 585
R28 B.n157 B.n156 585
R29 B.n155 B.n154 585
R30 B.n153 B.n152 585
R31 B.n151 B.n150 585
R32 B.n149 B.n148 585
R33 B.n147 B.n146 585
R34 B.n145 B.n144 585
R35 B.n143 B.n142 585
R36 B.n141 B.n140 585
R37 B.n139 B.n138 585
R38 B.n137 B.n136 585
R39 B.n135 B.n134 585
R40 B.n133 B.n132 585
R41 B.n131 B.n130 585
R42 B.n129 B.n128 585
R43 B.n127 B.n126 585
R44 B.n125 B.n124 585
R45 B.n123 B.n122 585
R46 B.n121 B.n120 585
R47 B.n119 B.n118 585
R48 B.n117 B.n116 585
R49 B.n115 B.n114 585
R50 B.n113 B.n112 585
R51 B.n111 B.n110 585
R52 B.n109 B.n108 585
R53 B.n107 B.n106 585
R54 B.n105 B.n104 585
R55 B.n103 B.n102 585
R56 B.n101 B.n100 585
R57 B.n99 B.n98 585
R58 B.n97 B.n96 585
R59 B.n95 B.n94 585
R60 B.n93 B.n92 585
R61 B.n91 B.n90 585
R62 B.n89 B.n88 585
R63 B.n87 B.n86 585
R64 B.n85 B.n84 585
R65 B.n83 B.n82 585
R66 B.n81 B.n80 585
R67 B.n79 B.n78 585
R68 B.n77 B.n76 585
R69 B.n75 B.n74 585
R70 B.n477 B.n34 585
R71 B.n482 B.n34 585
R72 B.n476 B.n33 585
R73 B.n483 B.n33 585
R74 B.n475 B.n474 585
R75 B.n474 B.n29 585
R76 B.n473 B.n28 585
R77 B.n489 B.n28 585
R78 B.n472 B.n27 585
R79 B.n490 B.n27 585
R80 B.n471 B.n26 585
R81 B.n491 B.n26 585
R82 B.n470 B.n469 585
R83 B.n469 B.n22 585
R84 B.n468 B.n21 585
R85 B.n497 B.n21 585
R86 B.n467 B.n20 585
R87 B.n498 B.n20 585
R88 B.n466 B.n19 585
R89 B.n499 B.n19 585
R90 B.n465 B.n464 585
R91 B.n464 B.n15 585
R92 B.n463 B.n14 585
R93 B.n505 B.n14 585
R94 B.n462 B.n13 585
R95 B.n506 B.n13 585
R96 B.n461 B.n12 585
R97 B.n507 B.n12 585
R98 B.n460 B.n459 585
R99 B.n459 B.n11 585
R100 B.n458 B.n7 585
R101 B.n513 B.n7 585
R102 B.n457 B.n6 585
R103 B.n514 B.n6 585
R104 B.n456 B.n5 585
R105 B.n515 B.n5 585
R106 B.n455 B.n454 585
R107 B.n454 B.n4 585
R108 B.n453 B.n203 585
R109 B.n453 B.n452 585
R110 B.n442 B.n204 585
R111 B.n445 B.n204 585
R112 B.n444 B.n443 585
R113 B.n446 B.n444 585
R114 B.n441 B.n208 585
R115 B.n212 B.n208 585
R116 B.n440 B.n439 585
R117 B.n439 B.n438 585
R118 B.n210 B.n209 585
R119 B.n211 B.n210 585
R120 B.n431 B.n430 585
R121 B.n432 B.n431 585
R122 B.n429 B.n217 585
R123 B.n217 B.n216 585
R124 B.n428 B.n427 585
R125 B.n427 B.n426 585
R126 B.n219 B.n218 585
R127 B.n220 B.n219 585
R128 B.n419 B.n418 585
R129 B.n420 B.n419 585
R130 B.n417 B.n224 585
R131 B.n228 B.n224 585
R132 B.n416 B.n415 585
R133 B.n415 B.n414 585
R134 B.n226 B.n225 585
R135 B.n227 B.n226 585
R136 B.n407 B.n406 585
R137 B.n408 B.n407 585
R138 B.n405 B.n233 585
R139 B.n233 B.n232 585
R140 B.n400 B.n399 585
R141 B.n398 B.n268 585
R142 B.n397 B.n267 585
R143 B.n402 B.n267 585
R144 B.n396 B.n395 585
R145 B.n394 B.n393 585
R146 B.n392 B.n391 585
R147 B.n390 B.n389 585
R148 B.n388 B.n387 585
R149 B.n386 B.n385 585
R150 B.n384 B.n383 585
R151 B.n382 B.n381 585
R152 B.n380 B.n379 585
R153 B.n378 B.n377 585
R154 B.n376 B.n375 585
R155 B.n374 B.n373 585
R156 B.n372 B.n371 585
R157 B.n370 B.n369 585
R158 B.n368 B.n367 585
R159 B.n366 B.n365 585
R160 B.n364 B.n363 585
R161 B.n362 B.n361 585
R162 B.n360 B.n359 585
R163 B.n358 B.n357 585
R164 B.n356 B.n355 585
R165 B.n354 B.n353 585
R166 B.n352 B.n351 585
R167 B.n350 B.n349 585
R168 B.n348 B.n347 585
R169 B.n345 B.n344 585
R170 B.n343 B.n342 585
R171 B.n341 B.n340 585
R172 B.n339 B.n338 585
R173 B.n337 B.n336 585
R174 B.n335 B.n334 585
R175 B.n333 B.n332 585
R176 B.n331 B.n330 585
R177 B.n329 B.n328 585
R178 B.n327 B.n326 585
R179 B.n324 B.n323 585
R180 B.n322 B.n321 585
R181 B.n320 B.n319 585
R182 B.n318 B.n317 585
R183 B.n316 B.n315 585
R184 B.n314 B.n313 585
R185 B.n312 B.n311 585
R186 B.n310 B.n309 585
R187 B.n308 B.n307 585
R188 B.n306 B.n305 585
R189 B.n304 B.n303 585
R190 B.n302 B.n301 585
R191 B.n300 B.n299 585
R192 B.n298 B.n297 585
R193 B.n296 B.n295 585
R194 B.n294 B.n293 585
R195 B.n292 B.n291 585
R196 B.n290 B.n289 585
R197 B.n288 B.n287 585
R198 B.n286 B.n285 585
R199 B.n284 B.n283 585
R200 B.n282 B.n281 585
R201 B.n280 B.n279 585
R202 B.n278 B.n277 585
R203 B.n276 B.n275 585
R204 B.n274 B.n273 585
R205 B.n235 B.n234 585
R206 B.n404 B.n403 585
R207 B.n403 B.n402 585
R208 B.n231 B.n230 585
R209 B.n232 B.n231 585
R210 B.n410 B.n409 585
R211 B.n409 B.n408 585
R212 B.n411 B.n229 585
R213 B.n229 B.n227 585
R214 B.n413 B.n412 585
R215 B.n414 B.n413 585
R216 B.n223 B.n222 585
R217 B.n228 B.n223 585
R218 B.n422 B.n421 585
R219 B.n421 B.n420 585
R220 B.n423 B.n221 585
R221 B.n221 B.n220 585
R222 B.n425 B.n424 585
R223 B.n426 B.n425 585
R224 B.n215 B.n214 585
R225 B.n216 B.n215 585
R226 B.n434 B.n433 585
R227 B.n433 B.n432 585
R228 B.n435 B.n213 585
R229 B.n213 B.n211 585
R230 B.n437 B.n436 585
R231 B.n438 B.n437 585
R232 B.n207 B.n206 585
R233 B.n212 B.n207 585
R234 B.n448 B.n447 585
R235 B.n447 B.n446 585
R236 B.n449 B.n205 585
R237 B.n445 B.n205 585
R238 B.n451 B.n450 585
R239 B.n452 B.n451 585
R240 B.n2 B.n0 585
R241 B.n4 B.n2 585
R242 B.n3 B.n1 585
R243 B.n514 B.n3 585
R244 B.n512 B.n511 585
R245 B.n513 B.n512 585
R246 B.n510 B.n8 585
R247 B.n11 B.n8 585
R248 B.n509 B.n508 585
R249 B.n508 B.n507 585
R250 B.n10 B.n9 585
R251 B.n506 B.n10 585
R252 B.n504 B.n503 585
R253 B.n505 B.n504 585
R254 B.n502 B.n16 585
R255 B.n16 B.n15 585
R256 B.n501 B.n500 585
R257 B.n500 B.n499 585
R258 B.n18 B.n17 585
R259 B.n498 B.n18 585
R260 B.n496 B.n495 585
R261 B.n497 B.n496 585
R262 B.n494 B.n23 585
R263 B.n23 B.n22 585
R264 B.n493 B.n492 585
R265 B.n492 B.n491 585
R266 B.n25 B.n24 585
R267 B.n490 B.n25 585
R268 B.n488 B.n487 585
R269 B.n489 B.n488 585
R270 B.n486 B.n30 585
R271 B.n30 B.n29 585
R272 B.n485 B.n484 585
R273 B.n484 B.n483 585
R274 B.n32 B.n31 585
R275 B.n482 B.n32 585
R276 B.n517 B.n516 585
R277 B.n516 B.n515 585
R278 B.n400 B.n231 487.695
R279 B.n74 B.n32 487.695
R280 B.n403 B.n233 487.695
R281 B.n479 B.n34 487.695
R282 B.n481 B.n480 256.663
R283 B.n481 B.n66 256.663
R284 B.n481 B.n65 256.663
R285 B.n481 B.n64 256.663
R286 B.n481 B.n63 256.663
R287 B.n481 B.n62 256.663
R288 B.n481 B.n61 256.663
R289 B.n481 B.n60 256.663
R290 B.n481 B.n59 256.663
R291 B.n481 B.n58 256.663
R292 B.n481 B.n57 256.663
R293 B.n481 B.n56 256.663
R294 B.n481 B.n55 256.663
R295 B.n481 B.n54 256.663
R296 B.n481 B.n53 256.663
R297 B.n481 B.n52 256.663
R298 B.n481 B.n51 256.663
R299 B.n481 B.n50 256.663
R300 B.n481 B.n49 256.663
R301 B.n481 B.n48 256.663
R302 B.n481 B.n47 256.663
R303 B.n481 B.n46 256.663
R304 B.n481 B.n45 256.663
R305 B.n481 B.n44 256.663
R306 B.n481 B.n43 256.663
R307 B.n481 B.n42 256.663
R308 B.n481 B.n41 256.663
R309 B.n481 B.n40 256.663
R310 B.n481 B.n39 256.663
R311 B.n481 B.n38 256.663
R312 B.n481 B.n37 256.663
R313 B.n481 B.n36 256.663
R314 B.n481 B.n35 256.663
R315 B.n402 B.n401 256.663
R316 B.n402 B.n236 256.663
R317 B.n402 B.n237 256.663
R318 B.n402 B.n238 256.663
R319 B.n402 B.n239 256.663
R320 B.n402 B.n240 256.663
R321 B.n402 B.n241 256.663
R322 B.n402 B.n242 256.663
R323 B.n402 B.n243 256.663
R324 B.n402 B.n244 256.663
R325 B.n402 B.n245 256.663
R326 B.n402 B.n246 256.663
R327 B.n402 B.n247 256.663
R328 B.n402 B.n248 256.663
R329 B.n402 B.n249 256.663
R330 B.n402 B.n250 256.663
R331 B.n402 B.n251 256.663
R332 B.n402 B.n252 256.663
R333 B.n402 B.n253 256.663
R334 B.n402 B.n254 256.663
R335 B.n402 B.n255 256.663
R336 B.n402 B.n256 256.663
R337 B.n402 B.n257 256.663
R338 B.n402 B.n258 256.663
R339 B.n402 B.n259 256.663
R340 B.n402 B.n260 256.663
R341 B.n402 B.n261 256.663
R342 B.n402 B.n262 256.663
R343 B.n402 B.n263 256.663
R344 B.n402 B.n264 256.663
R345 B.n402 B.n265 256.663
R346 B.n402 B.n266 256.663
R347 B.n271 B.t15 217.876
R348 B.n68 B.t7 217.876
R349 B.n269 B.t18 217.876
R350 B.n71 B.t10 217.876
R351 B.n272 B.t14 203.137
R352 B.n69 B.t8 203.137
R353 B.n270 B.t17 203.137
R354 B.n72 B.t11 203.137
R355 B.n409 B.n231 163.367
R356 B.n409 B.n229 163.367
R357 B.n413 B.n229 163.367
R358 B.n413 B.n223 163.367
R359 B.n421 B.n223 163.367
R360 B.n421 B.n221 163.367
R361 B.n425 B.n221 163.367
R362 B.n425 B.n215 163.367
R363 B.n433 B.n215 163.367
R364 B.n433 B.n213 163.367
R365 B.n437 B.n213 163.367
R366 B.n437 B.n207 163.367
R367 B.n447 B.n207 163.367
R368 B.n447 B.n205 163.367
R369 B.n451 B.n205 163.367
R370 B.n451 B.n2 163.367
R371 B.n516 B.n2 163.367
R372 B.n516 B.n3 163.367
R373 B.n512 B.n3 163.367
R374 B.n512 B.n8 163.367
R375 B.n508 B.n8 163.367
R376 B.n508 B.n10 163.367
R377 B.n504 B.n10 163.367
R378 B.n504 B.n16 163.367
R379 B.n500 B.n16 163.367
R380 B.n500 B.n18 163.367
R381 B.n496 B.n18 163.367
R382 B.n496 B.n23 163.367
R383 B.n492 B.n23 163.367
R384 B.n492 B.n25 163.367
R385 B.n488 B.n25 163.367
R386 B.n488 B.n30 163.367
R387 B.n484 B.n30 163.367
R388 B.n484 B.n32 163.367
R389 B.n268 B.n267 163.367
R390 B.n395 B.n267 163.367
R391 B.n393 B.n392 163.367
R392 B.n389 B.n388 163.367
R393 B.n385 B.n384 163.367
R394 B.n381 B.n380 163.367
R395 B.n377 B.n376 163.367
R396 B.n373 B.n372 163.367
R397 B.n369 B.n368 163.367
R398 B.n365 B.n364 163.367
R399 B.n361 B.n360 163.367
R400 B.n357 B.n356 163.367
R401 B.n353 B.n352 163.367
R402 B.n349 B.n348 163.367
R403 B.n344 B.n343 163.367
R404 B.n340 B.n339 163.367
R405 B.n336 B.n335 163.367
R406 B.n332 B.n331 163.367
R407 B.n328 B.n327 163.367
R408 B.n323 B.n322 163.367
R409 B.n319 B.n318 163.367
R410 B.n315 B.n314 163.367
R411 B.n311 B.n310 163.367
R412 B.n307 B.n306 163.367
R413 B.n303 B.n302 163.367
R414 B.n299 B.n298 163.367
R415 B.n295 B.n294 163.367
R416 B.n291 B.n290 163.367
R417 B.n287 B.n286 163.367
R418 B.n283 B.n282 163.367
R419 B.n279 B.n278 163.367
R420 B.n275 B.n274 163.367
R421 B.n403 B.n235 163.367
R422 B.n407 B.n233 163.367
R423 B.n407 B.n226 163.367
R424 B.n415 B.n226 163.367
R425 B.n415 B.n224 163.367
R426 B.n419 B.n224 163.367
R427 B.n419 B.n219 163.367
R428 B.n427 B.n219 163.367
R429 B.n427 B.n217 163.367
R430 B.n431 B.n217 163.367
R431 B.n431 B.n210 163.367
R432 B.n439 B.n210 163.367
R433 B.n439 B.n208 163.367
R434 B.n444 B.n208 163.367
R435 B.n444 B.n204 163.367
R436 B.n453 B.n204 163.367
R437 B.n454 B.n453 163.367
R438 B.n454 B.n5 163.367
R439 B.n6 B.n5 163.367
R440 B.n7 B.n6 163.367
R441 B.n459 B.n7 163.367
R442 B.n459 B.n12 163.367
R443 B.n13 B.n12 163.367
R444 B.n14 B.n13 163.367
R445 B.n464 B.n14 163.367
R446 B.n464 B.n19 163.367
R447 B.n20 B.n19 163.367
R448 B.n21 B.n20 163.367
R449 B.n469 B.n21 163.367
R450 B.n469 B.n26 163.367
R451 B.n27 B.n26 163.367
R452 B.n28 B.n27 163.367
R453 B.n474 B.n28 163.367
R454 B.n474 B.n33 163.367
R455 B.n34 B.n33 163.367
R456 B.n78 B.n77 163.367
R457 B.n82 B.n81 163.367
R458 B.n86 B.n85 163.367
R459 B.n90 B.n89 163.367
R460 B.n94 B.n93 163.367
R461 B.n98 B.n97 163.367
R462 B.n102 B.n101 163.367
R463 B.n106 B.n105 163.367
R464 B.n110 B.n109 163.367
R465 B.n114 B.n113 163.367
R466 B.n118 B.n117 163.367
R467 B.n122 B.n121 163.367
R468 B.n126 B.n125 163.367
R469 B.n130 B.n129 163.367
R470 B.n134 B.n133 163.367
R471 B.n138 B.n137 163.367
R472 B.n142 B.n141 163.367
R473 B.n146 B.n145 163.367
R474 B.n150 B.n149 163.367
R475 B.n154 B.n153 163.367
R476 B.n158 B.n157 163.367
R477 B.n162 B.n161 163.367
R478 B.n166 B.n165 163.367
R479 B.n170 B.n169 163.367
R480 B.n174 B.n173 163.367
R481 B.n178 B.n177 163.367
R482 B.n182 B.n181 163.367
R483 B.n186 B.n185 163.367
R484 B.n190 B.n189 163.367
R485 B.n194 B.n193 163.367
R486 B.n198 B.n197 163.367
R487 B.n200 B.n67 163.367
R488 B.n402 B.n232 110.218
R489 B.n482 B.n481 110.218
R490 B.n401 B.n400 71.676
R491 B.n395 B.n236 71.676
R492 B.n392 B.n237 71.676
R493 B.n388 B.n238 71.676
R494 B.n384 B.n239 71.676
R495 B.n380 B.n240 71.676
R496 B.n376 B.n241 71.676
R497 B.n372 B.n242 71.676
R498 B.n368 B.n243 71.676
R499 B.n364 B.n244 71.676
R500 B.n360 B.n245 71.676
R501 B.n356 B.n246 71.676
R502 B.n352 B.n247 71.676
R503 B.n348 B.n248 71.676
R504 B.n343 B.n249 71.676
R505 B.n339 B.n250 71.676
R506 B.n335 B.n251 71.676
R507 B.n331 B.n252 71.676
R508 B.n327 B.n253 71.676
R509 B.n322 B.n254 71.676
R510 B.n318 B.n255 71.676
R511 B.n314 B.n256 71.676
R512 B.n310 B.n257 71.676
R513 B.n306 B.n258 71.676
R514 B.n302 B.n259 71.676
R515 B.n298 B.n260 71.676
R516 B.n294 B.n261 71.676
R517 B.n290 B.n262 71.676
R518 B.n286 B.n263 71.676
R519 B.n282 B.n264 71.676
R520 B.n278 B.n265 71.676
R521 B.n274 B.n266 71.676
R522 B.n74 B.n35 71.676
R523 B.n78 B.n36 71.676
R524 B.n82 B.n37 71.676
R525 B.n86 B.n38 71.676
R526 B.n90 B.n39 71.676
R527 B.n94 B.n40 71.676
R528 B.n98 B.n41 71.676
R529 B.n102 B.n42 71.676
R530 B.n106 B.n43 71.676
R531 B.n110 B.n44 71.676
R532 B.n114 B.n45 71.676
R533 B.n118 B.n46 71.676
R534 B.n122 B.n47 71.676
R535 B.n126 B.n48 71.676
R536 B.n130 B.n49 71.676
R537 B.n134 B.n50 71.676
R538 B.n138 B.n51 71.676
R539 B.n142 B.n52 71.676
R540 B.n146 B.n53 71.676
R541 B.n150 B.n54 71.676
R542 B.n154 B.n55 71.676
R543 B.n158 B.n56 71.676
R544 B.n162 B.n57 71.676
R545 B.n166 B.n58 71.676
R546 B.n170 B.n59 71.676
R547 B.n174 B.n60 71.676
R548 B.n178 B.n61 71.676
R549 B.n182 B.n62 71.676
R550 B.n186 B.n63 71.676
R551 B.n190 B.n64 71.676
R552 B.n194 B.n65 71.676
R553 B.n198 B.n66 71.676
R554 B.n480 B.n67 71.676
R555 B.n480 B.n479 71.676
R556 B.n200 B.n66 71.676
R557 B.n197 B.n65 71.676
R558 B.n193 B.n64 71.676
R559 B.n189 B.n63 71.676
R560 B.n185 B.n62 71.676
R561 B.n181 B.n61 71.676
R562 B.n177 B.n60 71.676
R563 B.n173 B.n59 71.676
R564 B.n169 B.n58 71.676
R565 B.n165 B.n57 71.676
R566 B.n161 B.n56 71.676
R567 B.n157 B.n55 71.676
R568 B.n153 B.n54 71.676
R569 B.n149 B.n53 71.676
R570 B.n145 B.n52 71.676
R571 B.n141 B.n51 71.676
R572 B.n137 B.n50 71.676
R573 B.n133 B.n49 71.676
R574 B.n129 B.n48 71.676
R575 B.n125 B.n47 71.676
R576 B.n121 B.n46 71.676
R577 B.n117 B.n45 71.676
R578 B.n113 B.n44 71.676
R579 B.n109 B.n43 71.676
R580 B.n105 B.n42 71.676
R581 B.n101 B.n41 71.676
R582 B.n97 B.n40 71.676
R583 B.n93 B.n39 71.676
R584 B.n89 B.n38 71.676
R585 B.n85 B.n37 71.676
R586 B.n81 B.n36 71.676
R587 B.n77 B.n35 71.676
R588 B.n401 B.n268 71.676
R589 B.n393 B.n236 71.676
R590 B.n389 B.n237 71.676
R591 B.n385 B.n238 71.676
R592 B.n381 B.n239 71.676
R593 B.n377 B.n240 71.676
R594 B.n373 B.n241 71.676
R595 B.n369 B.n242 71.676
R596 B.n365 B.n243 71.676
R597 B.n361 B.n244 71.676
R598 B.n357 B.n245 71.676
R599 B.n353 B.n246 71.676
R600 B.n349 B.n247 71.676
R601 B.n344 B.n248 71.676
R602 B.n340 B.n249 71.676
R603 B.n336 B.n250 71.676
R604 B.n332 B.n251 71.676
R605 B.n328 B.n252 71.676
R606 B.n323 B.n253 71.676
R607 B.n319 B.n254 71.676
R608 B.n315 B.n255 71.676
R609 B.n311 B.n256 71.676
R610 B.n307 B.n257 71.676
R611 B.n303 B.n258 71.676
R612 B.n299 B.n259 71.676
R613 B.n295 B.n260 71.676
R614 B.n291 B.n261 71.676
R615 B.n287 B.n262 71.676
R616 B.n283 B.n263 71.676
R617 B.n279 B.n264 71.676
R618 B.n275 B.n265 71.676
R619 B.n266 B.n235 71.676
R620 B.n325 B.n272 59.5399
R621 B.n346 B.n270 59.5399
R622 B.n73 B.n72 59.5399
R623 B.n70 B.n69 59.5399
R624 B.n408 B.n232 59.0143
R625 B.n408 B.n227 59.0143
R626 B.n414 B.n227 59.0143
R627 B.n414 B.n228 59.0143
R628 B.n420 B.n220 59.0143
R629 B.n426 B.n220 59.0143
R630 B.n426 B.n216 59.0143
R631 B.n432 B.n216 59.0143
R632 B.n438 B.n211 59.0143
R633 B.n438 B.n212 59.0143
R634 B.n446 B.n445 59.0143
R635 B.n452 B.n4 59.0143
R636 B.n515 B.n4 59.0143
R637 B.n515 B.n514 59.0143
R638 B.n514 B.n513 59.0143
R639 B.n507 B.n11 59.0143
R640 B.n506 B.n505 59.0143
R641 B.n505 B.n15 59.0143
R642 B.n499 B.n498 59.0143
R643 B.n498 B.n497 59.0143
R644 B.n497 B.n22 59.0143
R645 B.n491 B.n22 59.0143
R646 B.n490 B.n489 59.0143
R647 B.n489 B.n29 59.0143
R648 B.n483 B.n29 59.0143
R649 B.n483 B.n482 59.0143
R650 B.n446 B.t19 56.4108
R651 B.n507 B.t4 56.4108
R652 B.n432 B.t0 47.7323
R653 B.n499 B.t3 47.7323
R654 B.n452 B.t1 42.5252
R655 B.n513 B.t2 42.5252
R656 B.n420 B.t13 37.3181
R657 B.n491 B.t6 37.3181
R658 B.n75 B.n31 31.6883
R659 B.n478 B.n477 31.6883
R660 B.n405 B.n404 31.6883
R661 B.n399 B.n230 31.6883
R662 B.n228 B.t13 21.6968
R663 B.t6 B.n490 21.6968
R664 B B.n517 18.0485
R665 B.n445 B.t1 16.4897
R666 B.n11 B.t2 16.4897
R667 B.n272 B.n271 14.7399
R668 B.n270 B.n269 14.7399
R669 B.n72 B.n71 14.7399
R670 B.n69 B.n68 14.7399
R671 B.t0 B.n211 11.2826
R672 B.t3 B.n15 11.2826
R673 B.n76 B.n75 10.6151
R674 B.n79 B.n76 10.6151
R675 B.n80 B.n79 10.6151
R676 B.n83 B.n80 10.6151
R677 B.n84 B.n83 10.6151
R678 B.n87 B.n84 10.6151
R679 B.n88 B.n87 10.6151
R680 B.n91 B.n88 10.6151
R681 B.n92 B.n91 10.6151
R682 B.n95 B.n92 10.6151
R683 B.n96 B.n95 10.6151
R684 B.n99 B.n96 10.6151
R685 B.n100 B.n99 10.6151
R686 B.n103 B.n100 10.6151
R687 B.n104 B.n103 10.6151
R688 B.n107 B.n104 10.6151
R689 B.n108 B.n107 10.6151
R690 B.n111 B.n108 10.6151
R691 B.n112 B.n111 10.6151
R692 B.n115 B.n112 10.6151
R693 B.n116 B.n115 10.6151
R694 B.n119 B.n116 10.6151
R695 B.n120 B.n119 10.6151
R696 B.n123 B.n120 10.6151
R697 B.n124 B.n123 10.6151
R698 B.n127 B.n124 10.6151
R699 B.n128 B.n127 10.6151
R700 B.n132 B.n131 10.6151
R701 B.n135 B.n132 10.6151
R702 B.n136 B.n135 10.6151
R703 B.n139 B.n136 10.6151
R704 B.n140 B.n139 10.6151
R705 B.n143 B.n140 10.6151
R706 B.n144 B.n143 10.6151
R707 B.n147 B.n144 10.6151
R708 B.n148 B.n147 10.6151
R709 B.n152 B.n151 10.6151
R710 B.n155 B.n152 10.6151
R711 B.n156 B.n155 10.6151
R712 B.n159 B.n156 10.6151
R713 B.n160 B.n159 10.6151
R714 B.n163 B.n160 10.6151
R715 B.n164 B.n163 10.6151
R716 B.n167 B.n164 10.6151
R717 B.n168 B.n167 10.6151
R718 B.n171 B.n168 10.6151
R719 B.n172 B.n171 10.6151
R720 B.n175 B.n172 10.6151
R721 B.n176 B.n175 10.6151
R722 B.n179 B.n176 10.6151
R723 B.n180 B.n179 10.6151
R724 B.n183 B.n180 10.6151
R725 B.n184 B.n183 10.6151
R726 B.n187 B.n184 10.6151
R727 B.n188 B.n187 10.6151
R728 B.n191 B.n188 10.6151
R729 B.n192 B.n191 10.6151
R730 B.n195 B.n192 10.6151
R731 B.n196 B.n195 10.6151
R732 B.n199 B.n196 10.6151
R733 B.n201 B.n199 10.6151
R734 B.n202 B.n201 10.6151
R735 B.n478 B.n202 10.6151
R736 B.n406 B.n405 10.6151
R737 B.n406 B.n225 10.6151
R738 B.n416 B.n225 10.6151
R739 B.n417 B.n416 10.6151
R740 B.n418 B.n417 10.6151
R741 B.n418 B.n218 10.6151
R742 B.n428 B.n218 10.6151
R743 B.n429 B.n428 10.6151
R744 B.n430 B.n429 10.6151
R745 B.n430 B.n209 10.6151
R746 B.n440 B.n209 10.6151
R747 B.n441 B.n440 10.6151
R748 B.n443 B.n441 10.6151
R749 B.n443 B.n442 10.6151
R750 B.n442 B.n203 10.6151
R751 B.n455 B.n203 10.6151
R752 B.n456 B.n455 10.6151
R753 B.n457 B.n456 10.6151
R754 B.n458 B.n457 10.6151
R755 B.n460 B.n458 10.6151
R756 B.n461 B.n460 10.6151
R757 B.n462 B.n461 10.6151
R758 B.n463 B.n462 10.6151
R759 B.n465 B.n463 10.6151
R760 B.n466 B.n465 10.6151
R761 B.n467 B.n466 10.6151
R762 B.n468 B.n467 10.6151
R763 B.n470 B.n468 10.6151
R764 B.n471 B.n470 10.6151
R765 B.n472 B.n471 10.6151
R766 B.n473 B.n472 10.6151
R767 B.n475 B.n473 10.6151
R768 B.n476 B.n475 10.6151
R769 B.n477 B.n476 10.6151
R770 B.n399 B.n398 10.6151
R771 B.n398 B.n397 10.6151
R772 B.n397 B.n396 10.6151
R773 B.n396 B.n394 10.6151
R774 B.n394 B.n391 10.6151
R775 B.n391 B.n390 10.6151
R776 B.n390 B.n387 10.6151
R777 B.n387 B.n386 10.6151
R778 B.n386 B.n383 10.6151
R779 B.n383 B.n382 10.6151
R780 B.n382 B.n379 10.6151
R781 B.n379 B.n378 10.6151
R782 B.n378 B.n375 10.6151
R783 B.n375 B.n374 10.6151
R784 B.n374 B.n371 10.6151
R785 B.n371 B.n370 10.6151
R786 B.n370 B.n367 10.6151
R787 B.n367 B.n366 10.6151
R788 B.n366 B.n363 10.6151
R789 B.n363 B.n362 10.6151
R790 B.n362 B.n359 10.6151
R791 B.n359 B.n358 10.6151
R792 B.n358 B.n355 10.6151
R793 B.n355 B.n354 10.6151
R794 B.n354 B.n351 10.6151
R795 B.n351 B.n350 10.6151
R796 B.n350 B.n347 10.6151
R797 B.n345 B.n342 10.6151
R798 B.n342 B.n341 10.6151
R799 B.n341 B.n338 10.6151
R800 B.n338 B.n337 10.6151
R801 B.n337 B.n334 10.6151
R802 B.n334 B.n333 10.6151
R803 B.n333 B.n330 10.6151
R804 B.n330 B.n329 10.6151
R805 B.n329 B.n326 10.6151
R806 B.n324 B.n321 10.6151
R807 B.n321 B.n320 10.6151
R808 B.n320 B.n317 10.6151
R809 B.n317 B.n316 10.6151
R810 B.n316 B.n313 10.6151
R811 B.n313 B.n312 10.6151
R812 B.n312 B.n309 10.6151
R813 B.n309 B.n308 10.6151
R814 B.n308 B.n305 10.6151
R815 B.n305 B.n304 10.6151
R816 B.n304 B.n301 10.6151
R817 B.n301 B.n300 10.6151
R818 B.n300 B.n297 10.6151
R819 B.n297 B.n296 10.6151
R820 B.n296 B.n293 10.6151
R821 B.n293 B.n292 10.6151
R822 B.n292 B.n289 10.6151
R823 B.n289 B.n288 10.6151
R824 B.n288 B.n285 10.6151
R825 B.n285 B.n284 10.6151
R826 B.n284 B.n281 10.6151
R827 B.n281 B.n280 10.6151
R828 B.n280 B.n277 10.6151
R829 B.n277 B.n276 10.6151
R830 B.n276 B.n273 10.6151
R831 B.n273 B.n234 10.6151
R832 B.n404 B.n234 10.6151
R833 B.n410 B.n230 10.6151
R834 B.n411 B.n410 10.6151
R835 B.n412 B.n411 10.6151
R836 B.n412 B.n222 10.6151
R837 B.n422 B.n222 10.6151
R838 B.n423 B.n422 10.6151
R839 B.n424 B.n423 10.6151
R840 B.n424 B.n214 10.6151
R841 B.n434 B.n214 10.6151
R842 B.n435 B.n434 10.6151
R843 B.n436 B.n435 10.6151
R844 B.n436 B.n206 10.6151
R845 B.n448 B.n206 10.6151
R846 B.n449 B.n448 10.6151
R847 B.n450 B.n449 10.6151
R848 B.n450 B.n0 10.6151
R849 B.n511 B.n1 10.6151
R850 B.n511 B.n510 10.6151
R851 B.n510 B.n509 10.6151
R852 B.n509 B.n9 10.6151
R853 B.n503 B.n9 10.6151
R854 B.n503 B.n502 10.6151
R855 B.n502 B.n501 10.6151
R856 B.n501 B.n17 10.6151
R857 B.n495 B.n17 10.6151
R858 B.n495 B.n494 10.6151
R859 B.n494 B.n493 10.6151
R860 B.n493 B.n24 10.6151
R861 B.n487 B.n24 10.6151
R862 B.n487 B.n486 10.6151
R863 B.n486 B.n485 10.6151
R864 B.n485 B.n31 10.6151
R865 B.n128 B.n73 9.36635
R866 B.n151 B.n70 9.36635
R867 B.n347 B.n346 9.36635
R868 B.n325 B.n324 9.36635
R869 B.n517 B.n0 2.81026
R870 B.n517 B.n1 2.81026
R871 B.n212 B.t19 2.60405
R872 B.t4 B.n506 2.60405
R873 B.n131 B.n73 1.24928
R874 B.n148 B.n70 1.24928
R875 B.n346 B.n345 1.24928
R876 B.n326 B.n325 1.24928
R877 VN.n0 VN.t0 532.241
R878 VN.n4 VN.t5 532.241
R879 VN.n2 VN.t2 513.794
R880 VN.n6 VN.t4 513.794
R881 VN.n1 VN.t1 507.221
R882 VN.n5 VN.t3 507.221
R883 VN.n3 VN.n2 161.3
R884 VN.n7 VN.n6 161.3
R885 VN.n7 VN.n4 71.6697
R886 VN.n3 VN.n0 71.6697
R887 VN.n2 VN.n1 41.6278
R888 VN.n6 VN.n5 41.6278
R889 VN VN.n7 37.1463
R890 VN.n5 VN.n4 18.4263
R891 VN.n1 VN.n0 18.4263
R892 VN VN.n3 0.0516364
R893 VTAIL.n162 VTAIL.n128 289.615
R894 VTAIL.n36 VTAIL.n2 289.615
R895 VTAIL.n122 VTAIL.n88 289.615
R896 VTAIL.n80 VTAIL.n46 289.615
R897 VTAIL.n140 VTAIL.n139 185
R898 VTAIL.n145 VTAIL.n144 185
R899 VTAIL.n147 VTAIL.n146 185
R900 VTAIL.n136 VTAIL.n135 185
R901 VTAIL.n153 VTAIL.n152 185
R902 VTAIL.n155 VTAIL.n154 185
R903 VTAIL.n132 VTAIL.n131 185
R904 VTAIL.n161 VTAIL.n160 185
R905 VTAIL.n163 VTAIL.n162 185
R906 VTAIL.n14 VTAIL.n13 185
R907 VTAIL.n19 VTAIL.n18 185
R908 VTAIL.n21 VTAIL.n20 185
R909 VTAIL.n10 VTAIL.n9 185
R910 VTAIL.n27 VTAIL.n26 185
R911 VTAIL.n29 VTAIL.n28 185
R912 VTAIL.n6 VTAIL.n5 185
R913 VTAIL.n35 VTAIL.n34 185
R914 VTAIL.n37 VTAIL.n36 185
R915 VTAIL.n123 VTAIL.n122 185
R916 VTAIL.n121 VTAIL.n120 185
R917 VTAIL.n92 VTAIL.n91 185
R918 VTAIL.n115 VTAIL.n114 185
R919 VTAIL.n113 VTAIL.n112 185
R920 VTAIL.n96 VTAIL.n95 185
R921 VTAIL.n107 VTAIL.n106 185
R922 VTAIL.n105 VTAIL.n104 185
R923 VTAIL.n100 VTAIL.n99 185
R924 VTAIL.n81 VTAIL.n80 185
R925 VTAIL.n79 VTAIL.n78 185
R926 VTAIL.n50 VTAIL.n49 185
R927 VTAIL.n73 VTAIL.n72 185
R928 VTAIL.n71 VTAIL.n70 185
R929 VTAIL.n54 VTAIL.n53 185
R930 VTAIL.n65 VTAIL.n64 185
R931 VTAIL.n63 VTAIL.n62 185
R932 VTAIL.n58 VTAIL.n57 185
R933 VTAIL.n141 VTAIL.t6 147.659
R934 VTAIL.n15 VTAIL.t3 147.659
R935 VTAIL.n101 VTAIL.t1 147.659
R936 VTAIL.n59 VTAIL.t7 147.659
R937 VTAIL.n145 VTAIL.n139 104.615
R938 VTAIL.n146 VTAIL.n145 104.615
R939 VTAIL.n146 VTAIL.n135 104.615
R940 VTAIL.n153 VTAIL.n135 104.615
R941 VTAIL.n154 VTAIL.n153 104.615
R942 VTAIL.n154 VTAIL.n131 104.615
R943 VTAIL.n161 VTAIL.n131 104.615
R944 VTAIL.n162 VTAIL.n161 104.615
R945 VTAIL.n19 VTAIL.n13 104.615
R946 VTAIL.n20 VTAIL.n19 104.615
R947 VTAIL.n20 VTAIL.n9 104.615
R948 VTAIL.n27 VTAIL.n9 104.615
R949 VTAIL.n28 VTAIL.n27 104.615
R950 VTAIL.n28 VTAIL.n5 104.615
R951 VTAIL.n35 VTAIL.n5 104.615
R952 VTAIL.n36 VTAIL.n35 104.615
R953 VTAIL.n122 VTAIL.n121 104.615
R954 VTAIL.n121 VTAIL.n91 104.615
R955 VTAIL.n114 VTAIL.n91 104.615
R956 VTAIL.n114 VTAIL.n113 104.615
R957 VTAIL.n113 VTAIL.n95 104.615
R958 VTAIL.n106 VTAIL.n95 104.615
R959 VTAIL.n106 VTAIL.n105 104.615
R960 VTAIL.n105 VTAIL.n99 104.615
R961 VTAIL.n80 VTAIL.n79 104.615
R962 VTAIL.n79 VTAIL.n49 104.615
R963 VTAIL.n72 VTAIL.n49 104.615
R964 VTAIL.n72 VTAIL.n71 104.615
R965 VTAIL.n71 VTAIL.n53 104.615
R966 VTAIL.n64 VTAIL.n53 104.615
R967 VTAIL.n64 VTAIL.n63 104.615
R968 VTAIL.n63 VTAIL.n57 104.615
R969 VTAIL.t6 VTAIL.n139 52.3082
R970 VTAIL.t3 VTAIL.n13 52.3082
R971 VTAIL.t1 VTAIL.n99 52.3082
R972 VTAIL.t7 VTAIL.n57 52.3082
R973 VTAIL.n87 VTAIL.n86 47.746
R974 VTAIL.n45 VTAIL.n44 47.746
R975 VTAIL.n1 VTAIL.n0 47.7458
R976 VTAIL.n43 VTAIL.n42 47.7458
R977 VTAIL.n167 VTAIL.n166 31.4096
R978 VTAIL.n41 VTAIL.n40 31.4096
R979 VTAIL.n127 VTAIL.n126 31.4096
R980 VTAIL.n85 VTAIL.n84 31.4096
R981 VTAIL.n45 VTAIL.n43 20.0565
R982 VTAIL.n167 VTAIL.n127 19.4014
R983 VTAIL.n141 VTAIL.n140 15.6677
R984 VTAIL.n15 VTAIL.n14 15.6677
R985 VTAIL.n101 VTAIL.n100 15.6677
R986 VTAIL.n59 VTAIL.n58 15.6677
R987 VTAIL.n144 VTAIL.n143 12.8005
R988 VTAIL.n18 VTAIL.n17 12.8005
R989 VTAIL.n104 VTAIL.n103 12.8005
R990 VTAIL.n62 VTAIL.n61 12.8005
R991 VTAIL.n147 VTAIL.n138 12.0247
R992 VTAIL.n21 VTAIL.n12 12.0247
R993 VTAIL.n107 VTAIL.n98 12.0247
R994 VTAIL.n65 VTAIL.n56 12.0247
R995 VTAIL.n148 VTAIL.n136 11.249
R996 VTAIL.n22 VTAIL.n10 11.249
R997 VTAIL.n108 VTAIL.n96 11.249
R998 VTAIL.n66 VTAIL.n54 11.249
R999 VTAIL.n152 VTAIL.n151 10.4732
R1000 VTAIL.n26 VTAIL.n25 10.4732
R1001 VTAIL.n112 VTAIL.n111 10.4732
R1002 VTAIL.n70 VTAIL.n69 10.4732
R1003 VTAIL.n155 VTAIL.n134 9.69747
R1004 VTAIL.n29 VTAIL.n8 9.69747
R1005 VTAIL.n115 VTAIL.n94 9.69747
R1006 VTAIL.n73 VTAIL.n52 9.69747
R1007 VTAIL.n166 VTAIL.n165 9.45567
R1008 VTAIL.n40 VTAIL.n39 9.45567
R1009 VTAIL.n126 VTAIL.n125 9.45567
R1010 VTAIL.n84 VTAIL.n83 9.45567
R1011 VTAIL.n165 VTAIL.n164 9.3005
R1012 VTAIL.n159 VTAIL.n158 9.3005
R1013 VTAIL.n157 VTAIL.n156 9.3005
R1014 VTAIL.n134 VTAIL.n133 9.3005
R1015 VTAIL.n151 VTAIL.n150 9.3005
R1016 VTAIL.n149 VTAIL.n148 9.3005
R1017 VTAIL.n138 VTAIL.n137 9.3005
R1018 VTAIL.n143 VTAIL.n142 9.3005
R1019 VTAIL.n130 VTAIL.n129 9.3005
R1020 VTAIL.n39 VTAIL.n38 9.3005
R1021 VTAIL.n33 VTAIL.n32 9.3005
R1022 VTAIL.n31 VTAIL.n30 9.3005
R1023 VTAIL.n8 VTAIL.n7 9.3005
R1024 VTAIL.n25 VTAIL.n24 9.3005
R1025 VTAIL.n23 VTAIL.n22 9.3005
R1026 VTAIL.n12 VTAIL.n11 9.3005
R1027 VTAIL.n17 VTAIL.n16 9.3005
R1028 VTAIL.n4 VTAIL.n3 9.3005
R1029 VTAIL.n125 VTAIL.n124 9.3005
R1030 VTAIL.n90 VTAIL.n89 9.3005
R1031 VTAIL.n119 VTAIL.n118 9.3005
R1032 VTAIL.n117 VTAIL.n116 9.3005
R1033 VTAIL.n94 VTAIL.n93 9.3005
R1034 VTAIL.n111 VTAIL.n110 9.3005
R1035 VTAIL.n109 VTAIL.n108 9.3005
R1036 VTAIL.n98 VTAIL.n97 9.3005
R1037 VTAIL.n103 VTAIL.n102 9.3005
R1038 VTAIL.n83 VTAIL.n82 9.3005
R1039 VTAIL.n48 VTAIL.n47 9.3005
R1040 VTAIL.n77 VTAIL.n76 9.3005
R1041 VTAIL.n75 VTAIL.n74 9.3005
R1042 VTAIL.n52 VTAIL.n51 9.3005
R1043 VTAIL.n69 VTAIL.n68 9.3005
R1044 VTAIL.n67 VTAIL.n66 9.3005
R1045 VTAIL.n56 VTAIL.n55 9.3005
R1046 VTAIL.n61 VTAIL.n60 9.3005
R1047 VTAIL.n156 VTAIL.n132 8.92171
R1048 VTAIL.n30 VTAIL.n6 8.92171
R1049 VTAIL.n116 VTAIL.n92 8.92171
R1050 VTAIL.n74 VTAIL.n50 8.92171
R1051 VTAIL.n160 VTAIL.n159 8.14595
R1052 VTAIL.n34 VTAIL.n33 8.14595
R1053 VTAIL.n120 VTAIL.n119 8.14595
R1054 VTAIL.n78 VTAIL.n77 8.14595
R1055 VTAIL.n163 VTAIL.n130 7.3702
R1056 VTAIL.n166 VTAIL.n128 7.3702
R1057 VTAIL.n37 VTAIL.n4 7.3702
R1058 VTAIL.n40 VTAIL.n2 7.3702
R1059 VTAIL.n126 VTAIL.n88 7.3702
R1060 VTAIL.n123 VTAIL.n90 7.3702
R1061 VTAIL.n84 VTAIL.n46 7.3702
R1062 VTAIL.n81 VTAIL.n48 7.3702
R1063 VTAIL.n164 VTAIL.n163 6.59444
R1064 VTAIL.n164 VTAIL.n128 6.59444
R1065 VTAIL.n38 VTAIL.n37 6.59444
R1066 VTAIL.n38 VTAIL.n2 6.59444
R1067 VTAIL.n124 VTAIL.n88 6.59444
R1068 VTAIL.n124 VTAIL.n123 6.59444
R1069 VTAIL.n82 VTAIL.n46 6.59444
R1070 VTAIL.n82 VTAIL.n81 6.59444
R1071 VTAIL.n160 VTAIL.n130 5.81868
R1072 VTAIL.n34 VTAIL.n4 5.81868
R1073 VTAIL.n120 VTAIL.n90 5.81868
R1074 VTAIL.n78 VTAIL.n48 5.81868
R1075 VTAIL.n159 VTAIL.n132 5.04292
R1076 VTAIL.n33 VTAIL.n6 5.04292
R1077 VTAIL.n119 VTAIL.n92 5.04292
R1078 VTAIL.n77 VTAIL.n50 5.04292
R1079 VTAIL.n102 VTAIL.n101 4.38565
R1080 VTAIL.n60 VTAIL.n59 4.38565
R1081 VTAIL.n142 VTAIL.n141 4.38565
R1082 VTAIL.n16 VTAIL.n15 4.38565
R1083 VTAIL.n156 VTAIL.n155 4.26717
R1084 VTAIL.n30 VTAIL.n29 4.26717
R1085 VTAIL.n116 VTAIL.n115 4.26717
R1086 VTAIL.n74 VTAIL.n73 4.26717
R1087 VTAIL.n152 VTAIL.n134 3.49141
R1088 VTAIL.n26 VTAIL.n8 3.49141
R1089 VTAIL.n112 VTAIL.n94 3.49141
R1090 VTAIL.n70 VTAIL.n52 3.49141
R1091 VTAIL.n151 VTAIL.n136 2.71565
R1092 VTAIL.n25 VTAIL.n10 2.71565
R1093 VTAIL.n111 VTAIL.n96 2.71565
R1094 VTAIL.n69 VTAIL.n54 2.71565
R1095 VTAIL.n0 VTAIL.t10 2.67618
R1096 VTAIL.n0 VTAIL.t8 2.67618
R1097 VTAIL.n42 VTAIL.t4 2.67618
R1098 VTAIL.n42 VTAIL.t5 2.67618
R1099 VTAIL.n86 VTAIL.t0 2.67618
R1100 VTAIL.n86 VTAIL.t2 2.67618
R1101 VTAIL.n44 VTAIL.t9 2.67618
R1102 VTAIL.n44 VTAIL.t11 2.67618
R1103 VTAIL.n148 VTAIL.n147 1.93989
R1104 VTAIL.n22 VTAIL.n21 1.93989
R1105 VTAIL.n108 VTAIL.n107 1.93989
R1106 VTAIL.n66 VTAIL.n65 1.93989
R1107 VTAIL.n144 VTAIL.n138 1.16414
R1108 VTAIL.n18 VTAIL.n12 1.16414
R1109 VTAIL.n104 VTAIL.n98 1.16414
R1110 VTAIL.n62 VTAIL.n56 1.16414
R1111 VTAIL.n87 VTAIL.n85 0.797914
R1112 VTAIL.n41 VTAIL.n1 0.797914
R1113 VTAIL.n85 VTAIL.n45 0.655672
R1114 VTAIL.n127 VTAIL.n87 0.655672
R1115 VTAIL.n43 VTAIL.n41 0.655672
R1116 VTAIL VTAIL.n167 0.43369
R1117 VTAIL.n143 VTAIL.n140 0.388379
R1118 VTAIL.n17 VTAIL.n14 0.388379
R1119 VTAIL.n103 VTAIL.n100 0.388379
R1120 VTAIL.n61 VTAIL.n58 0.388379
R1121 VTAIL VTAIL.n1 0.222483
R1122 VTAIL.n142 VTAIL.n137 0.155672
R1123 VTAIL.n149 VTAIL.n137 0.155672
R1124 VTAIL.n150 VTAIL.n149 0.155672
R1125 VTAIL.n150 VTAIL.n133 0.155672
R1126 VTAIL.n157 VTAIL.n133 0.155672
R1127 VTAIL.n158 VTAIL.n157 0.155672
R1128 VTAIL.n158 VTAIL.n129 0.155672
R1129 VTAIL.n165 VTAIL.n129 0.155672
R1130 VTAIL.n16 VTAIL.n11 0.155672
R1131 VTAIL.n23 VTAIL.n11 0.155672
R1132 VTAIL.n24 VTAIL.n23 0.155672
R1133 VTAIL.n24 VTAIL.n7 0.155672
R1134 VTAIL.n31 VTAIL.n7 0.155672
R1135 VTAIL.n32 VTAIL.n31 0.155672
R1136 VTAIL.n32 VTAIL.n3 0.155672
R1137 VTAIL.n39 VTAIL.n3 0.155672
R1138 VTAIL.n125 VTAIL.n89 0.155672
R1139 VTAIL.n118 VTAIL.n89 0.155672
R1140 VTAIL.n118 VTAIL.n117 0.155672
R1141 VTAIL.n117 VTAIL.n93 0.155672
R1142 VTAIL.n110 VTAIL.n93 0.155672
R1143 VTAIL.n110 VTAIL.n109 0.155672
R1144 VTAIL.n109 VTAIL.n97 0.155672
R1145 VTAIL.n102 VTAIL.n97 0.155672
R1146 VTAIL.n83 VTAIL.n47 0.155672
R1147 VTAIL.n76 VTAIL.n47 0.155672
R1148 VTAIL.n76 VTAIL.n75 0.155672
R1149 VTAIL.n75 VTAIL.n51 0.155672
R1150 VTAIL.n68 VTAIL.n51 0.155672
R1151 VTAIL.n68 VTAIL.n67 0.155672
R1152 VTAIL.n67 VTAIL.n55 0.155672
R1153 VTAIL.n60 VTAIL.n55 0.155672
R1154 VDD2.n75 VDD2.n41 289.615
R1155 VDD2.n34 VDD2.n0 289.615
R1156 VDD2.n76 VDD2.n75 185
R1157 VDD2.n74 VDD2.n73 185
R1158 VDD2.n45 VDD2.n44 185
R1159 VDD2.n68 VDD2.n67 185
R1160 VDD2.n66 VDD2.n65 185
R1161 VDD2.n49 VDD2.n48 185
R1162 VDD2.n60 VDD2.n59 185
R1163 VDD2.n58 VDD2.n57 185
R1164 VDD2.n53 VDD2.n52 185
R1165 VDD2.n12 VDD2.n11 185
R1166 VDD2.n17 VDD2.n16 185
R1167 VDD2.n19 VDD2.n18 185
R1168 VDD2.n8 VDD2.n7 185
R1169 VDD2.n25 VDD2.n24 185
R1170 VDD2.n27 VDD2.n26 185
R1171 VDD2.n4 VDD2.n3 185
R1172 VDD2.n33 VDD2.n32 185
R1173 VDD2.n35 VDD2.n34 185
R1174 VDD2.n54 VDD2.t1 147.659
R1175 VDD2.n13 VDD2.t5 147.659
R1176 VDD2.n75 VDD2.n74 104.615
R1177 VDD2.n74 VDD2.n44 104.615
R1178 VDD2.n67 VDD2.n44 104.615
R1179 VDD2.n67 VDD2.n66 104.615
R1180 VDD2.n66 VDD2.n48 104.615
R1181 VDD2.n59 VDD2.n48 104.615
R1182 VDD2.n59 VDD2.n58 104.615
R1183 VDD2.n58 VDD2.n52 104.615
R1184 VDD2.n17 VDD2.n11 104.615
R1185 VDD2.n18 VDD2.n17 104.615
R1186 VDD2.n18 VDD2.n7 104.615
R1187 VDD2.n25 VDD2.n7 104.615
R1188 VDD2.n26 VDD2.n25 104.615
R1189 VDD2.n26 VDD2.n3 104.615
R1190 VDD2.n33 VDD2.n3 104.615
R1191 VDD2.n34 VDD2.n33 104.615
R1192 VDD2.n40 VDD2.n39 64.533
R1193 VDD2 VDD2.n81 64.5302
R1194 VDD2.t1 VDD2.n52 52.3082
R1195 VDD2.t5 VDD2.n11 52.3082
R1196 VDD2.n40 VDD2.n38 48.5244
R1197 VDD2.n80 VDD2.n79 48.0884
R1198 VDD2.n80 VDD2.n40 32.2239
R1199 VDD2.n54 VDD2.n53 15.6677
R1200 VDD2.n13 VDD2.n12 15.6677
R1201 VDD2.n57 VDD2.n56 12.8005
R1202 VDD2.n16 VDD2.n15 12.8005
R1203 VDD2.n60 VDD2.n51 12.0247
R1204 VDD2.n19 VDD2.n10 12.0247
R1205 VDD2.n61 VDD2.n49 11.249
R1206 VDD2.n20 VDD2.n8 11.249
R1207 VDD2.n65 VDD2.n64 10.4732
R1208 VDD2.n24 VDD2.n23 10.4732
R1209 VDD2.n68 VDD2.n47 9.69747
R1210 VDD2.n27 VDD2.n6 9.69747
R1211 VDD2.n79 VDD2.n78 9.45567
R1212 VDD2.n38 VDD2.n37 9.45567
R1213 VDD2.n78 VDD2.n77 9.3005
R1214 VDD2.n43 VDD2.n42 9.3005
R1215 VDD2.n72 VDD2.n71 9.3005
R1216 VDD2.n70 VDD2.n69 9.3005
R1217 VDD2.n47 VDD2.n46 9.3005
R1218 VDD2.n64 VDD2.n63 9.3005
R1219 VDD2.n62 VDD2.n61 9.3005
R1220 VDD2.n51 VDD2.n50 9.3005
R1221 VDD2.n56 VDD2.n55 9.3005
R1222 VDD2.n37 VDD2.n36 9.3005
R1223 VDD2.n31 VDD2.n30 9.3005
R1224 VDD2.n29 VDD2.n28 9.3005
R1225 VDD2.n6 VDD2.n5 9.3005
R1226 VDD2.n23 VDD2.n22 9.3005
R1227 VDD2.n21 VDD2.n20 9.3005
R1228 VDD2.n10 VDD2.n9 9.3005
R1229 VDD2.n15 VDD2.n14 9.3005
R1230 VDD2.n2 VDD2.n1 9.3005
R1231 VDD2.n69 VDD2.n45 8.92171
R1232 VDD2.n28 VDD2.n4 8.92171
R1233 VDD2.n73 VDD2.n72 8.14595
R1234 VDD2.n32 VDD2.n31 8.14595
R1235 VDD2.n79 VDD2.n41 7.3702
R1236 VDD2.n76 VDD2.n43 7.3702
R1237 VDD2.n35 VDD2.n2 7.3702
R1238 VDD2.n38 VDD2.n0 7.3702
R1239 VDD2.n77 VDD2.n41 6.59444
R1240 VDD2.n77 VDD2.n76 6.59444
R1241 VDD2.n36 VDD2.n35 6.59444
R1242 VDD2.n36 VDD2.n0 6.59444
R1243 VDD2.n73 VDD2.n43 5.81868
R1244 VDD2.n32 VDD2.n2 5.81868
R1245 VDD2.n72 VDD2.n45 5.04292
R1246 VDD2.n31 VDD2.n4 5.04292
R1247 VDD2.n55 VDD2.n54 4.38565
R1248 VDD2.n14 VDD2.n13 4.38565
R1249 VDD2.n69 VDD2.n68 4.26717
R1250 VDD2.n28 VDD2.n27 4.26717
R1251 VDD2.n65 VDD2.n47 3.49141
R1252 VDD2.n24 VDD2.n6 3.49141
R1253 VDD2.n64 VDD2.n49 2.71565
R1254 VDD2.n23 VDD2.n8 2.71565
R1255 VDD2.n81 VDD2.t2 2.67618
R1256 VDD2.n81 VDD2.t0 2.67618
R1257 VDD2.n39 VDD2.t4 2.67618
R1258 VDD2.n39 VDD2.t3 2.67618
R1259 VDD2.n61 VDD2.n60 1.93989
R1260 VDD2.n20 VDD2.n19 1.93989
R1261 VDD2.n57 VDD2.n51 1.16414
R1262 VDD2.n16 VDD2.n10 1.16414
R1263 VDD2 VDD2.n80 0.550069
R1264 VDD2.n56 VDD2.n53 0.388379
R1265 VDD2.n15 VDD2.n12 0.388379
R1266 VDD2.n78 VDD2.n42 0.155672
R1267 VDD2.n71 VDD2.n42 0.155672
R1268 VDD2.n71 VDD2.n70 0.155672
R1269 VDD2.n70 VDD2.n46 0.155672
R1270 VDD2.n63 VDD2.n46 0.155672
R1271 VDD2.n63 VDD2.n62 0.155672
R1272 VDD2.n62 VDD2.n50 0.155672
R1273 VDD2.n55 VDD2.n50 0.155672
R1274 VDD2.n14 VDD2.n9 0.155672
R1275 VDD2.n21 VDD2.n9 0.155672
R1276 VDD2.n22 VDD2.n21 0.155672
R1277 VDD2.n22 VDD2.n5 0.155672
R1278 VDD2.n29 VDD2.n5 0.155672
R1279 VDD2.n30 VDD2.n29 0.155672
R1280 VDD2.n30 VDD2.n1 0.155672
R1281 VDD2.n37 VDD2.n1 0.155672
R1282 VP.n1 VP.t5 532.241
R1283 VP.n8 VP.t0 513.794
R1284 VP.n6 VP.t4 513.794
R1285 VP.n3 VP.t2 513.794
R1286 VP.n7 VP.t1 507.221
R1287 VP.n2 VP.t3 507.221
R1288 VP.n9 VP.n8 161.3
R1289 VP.n4 VP.n3 161.3
R1290 VP.n7 VP.n0 161.3
R1291 VP.n6 VP.n5 161.3
R1292 VP.n4 VP.n1 71.6697
R1293 VP.n7 VP.n6 41.6278
R1294 VP.n8 VP.n7 41.6278
R1295 VP.n3 VP.n2 41.6278
R1296 VP.n5 VP.n4 36.7657
R1297 VP.n2 VP.n1 18.4263
R1298 VP.n5 VP.n0 0.189894
R1299 VP.n9 VP.n0 0.189894
R1300 VP VP.n9 0.0516364
R1301 VDD1.n34 VDD1.n0 289.615
R1302 VDD1.n73 VDD1.n39 289.615
R1303 VDD1.n35 VDD1.n34 185
R1304 VDD1.n33 VDD1.n32 185
R1305 VDD1.n4 VDD1.n3 185
R1306 VDD1.n27 VDD1.n26 185
R1307 VDD1.n25 VDD1.n24 185
R1308 VDD1.n8 VDD1.n7 185
R1309 VDD1.n19 VDD1.n18 185
R1310 VDD1.n17 VDD1.n16 185
R1311 VDD1.n12 VDD1.n11 185
R1312 VDD1.n51 VDD1.n50 185
R1313 VDD1.n56 VDD1.n55 185
R1314 VDD1.n58 VDD1.n57 185
R1315 VDD1.n47 VDD1.n46 185
R1316 VDD1.n64 VDD1.n63 185
R1317 VDD1.n66 VDD1.n65 185
R1318 VDD1.n43 VDD1.n42 185
R1319 VDD1.n72 VDD1.n71 185
R1320 VDD1.n74 VDD1.n73 185
R1321 VDD1.n13 VDD1.t0 147.659
R1322 VDD1.n52 VDD1.t1 147.659
R1323 VDD1.n34 VDD1.n33 104.615
R1324 VDD1.n33 VDD1.n3 104.615
R1325 VDD1.n26 VDD1.n3 104.615
R1326 VDD1.n26 VDD1.n25 104.615
R1327 VDD1.n25 VDD1.n7 104.615
R1328 VDD1.n18 VDD1.n7 104.615
R1329 VDD1.n18 VDD1.n17 104.615
R1330 VDD1.n17 VDD1.n11 104.615
R1331 VDD1.n56 VDD1.n50 104.615
R1332 VDD1.n57 VDD1.n56 104.615
R1333 VDD1.n57 VDD1.n46 104.615
R1334 VDD1.n64 VDD1.n46 104.615
R1335 VDD1.n65 VDD1.n64 104.615
R1336 VDD1.n65 VDD1.n42 104.615
R1337 VDD1.n72 VDD1.n42 104.615
R1338 VDD1.n73 VDD1.n72 104.615
R1339 VDD1.n79 VDD1.n78 64.533
R1340 VDD1.n81 VDD1.n80 64.4246
R1341 VDD1.t0 VDD1.n11 52.3082
R1342 VDD1.t1 VDD1.n50 52.3082
R1343 VDD1 VDD1.n38 48.6379
R1344 VDD1.n79 VDD1.n77 48.5244
R1345 VDD1.n81 VDD1.n79 33.1345
R1346 VDD1.n13 VDD1.n12 15.6677
R1347 VDD1.n52 VDD1.n51 15.6677
R1348 VDD1.n16 VDD1.n15 12.8005
R1349 VDD1.n55 VDD1.n54 12.8005
R1350 VDD1.n19 VDD1.n10 12.0247
R1351 VDD1.n58 VDD1.n49 12.0247
R1352 VDD1.n20 VDD1.n8 11.249
R1353 VDD1.n59 VDD1.n47 11.249
R1354 VDD1.n24 VDD1.n23 10.4732
R1355 VDD1.n63 VDD1.n62 10.4732
R1356 VDD1.n27 VDD1.n6 9.69747
R1357 VDD1.n66 VDD1.n45 9.69747
R1358 VDD1.n38 VDD1.n37 9.45567
R1359 VDD1.n77 VDD1.n76 9.45567
R1360 VDD1.n37 VDD1.n36 9.3005
R1361 VDD1.n2 VDD1.n1 9.3005
R1362 VDD1.n31 VDD1.n30 9.3005
R1363 VDD1.n29 VDD1.n28 9.3005
R1364 VDD1.n6 VDD1.n5 9.3005
R1365 VDD1.n23 VDD1.n22 9.3005
R1366 VDD1.n21 VDD1.n20 9.3005
R1367 VDD1.n10 VDD1.n9 9.3005
R1368 VDD1.n15 VDD1.n14 9.3005
R1369 VDD1.n76 VDD1.n75 9.3005
R1370 VDD1.n70 VDD1.n69 9.3005
R1371 VDD1.n68 VDD1.n67 9.3005
R1372 VDD1.n45 VDD1.n44 9.3005
R1373 VDD1.n62 VDD1.n61 9.3005
R1374 VDD1.n60 VDD1.n59 9.3005
R1375 VDD1.n49 VDD1.n48 9.3005
R1376 VDD1.n54 VDD1.n53 9.3005
R1377 VDD1.n41 VDD1.n40 9.3005
R1378 VDD1.n28 VDD1.n4 8.92171
R1379 VDD1.n67 VDD1.n43 8.92171
R1380 VDD1.n32 VDD1.n31 8.14595
R1381 VDD1.n71 VDD1.n70 8.14595
R1382 VDD1.n38 VDD1.n0 7.3702
R1383 VDD1.n35 VDD1.n2 7.3702
R1384 VDD1.n74 VDD1.n41 7.3702
R1385 VDD1.n77 VDD1.n39 7.3702
R1386 VDD1.n36 VDD1.n0 6.59444
R1387 VDD1.n36 VDD1.n35 6.59444
R1388 VDD1.n75 VDD1.n74 6.59444
R1389 VDD1.n75 VDD1.n39 6.59444
R1390 VDD1.n32 VDD1.n2 5.81868
R1391 VDD1.n71 VDD1.n41 5.81868
R1392 VDD1.n31 VDD1.n4 5.04292
R1393 VDD1.n70 VDD1.n43 5.04292
R1394 VDD1.n14 VDD1.n13 4.38565
R1395 VDD1.n53 VDD1.n52 4.38565
R1396 VDD1.n28 VDD1.n27 4.26717
R1397 VDD1.n67 VDD1.n66 4.26717
R1398 VDD1.n24 VDD1.n6 3.49141
R1399 VDD1.n63 VDD1.n45 3.49141
R1400 VDD1.n23 VDD1.n8 2.71565
R1401 VDD1.n62 VDD1.n47 2.71565
R1402 VDD1.n80 VDD1.t2 2.67618
R1403 VDD1.n80 VDD1.t3 2.67618
R1404 VDD1.n78 VDD1.t4 2.67618
R1405 VDD1.n78 VDD1.t5 2.67618
R1406 VDD1.n20 VDD1.n19 1.93989
R1407 VDD1.n59 VDD1.n58 1.93989
R1408 VDD1.n16 VDD1.n10 1.16414
R1409 VDD1.n55 VDD1.n49 1.16414
R1410 VDD1.n15 VDD1.n12 0.388379
R1411 VDD1.n54 VDD1.n51 0.388379
R1412 VDD1.n37 VDD1.n1 0.155672
R1413 VDD1.n30 VDD1.n1 0.155672
R1414 VDD1.n30 VDD1.n29 0.155672
R1415 VDD1.n29 VDD1.n5 0.155672
R1416 VDD1.n22 VDD1.n5 0.155672
R1417 VDD1.n22 VDD1.n21 0.155672
R1418 VDD1.n21 VDD1.n9 0.155672
R1419 VDD1.n14 VDD1.n9 0.155672
R1420 VDD1.n53 VDD1.n48 0.155672
R1421 VDD1.n60 VDD1.n48 0.155672
R1422 VDD1.n61 VDD1.n60 0.155672
R1423 VDD1.n61 VDD1.n44 0.155672
R1424 VDD1.n68 VDD1.n44 0.155672
R1425 VDD1.n69 VDD1.n68 0.155672
R1426 VDD1.n69 VDD1.n40 0.155672
R1427 VDD1.n76 VDD1.n40 0.155672
R1428 VDD1 VDD1.n81 0.106103
C0 VDD1 VDD2 0.613385f
C1 VP VN 3.96696f
C2 VDD2 VN 2.18063f
C3 VDD2 VP 0.273734f
C4 VDD1 VTAIL 8.06937f
C5 VTAIL VN 1.96582f
C6 VTAIL VP 1.9803f
C7 VDD1 VN 0.147406f
C8 VDD1 VP 2.30381f
C9 VTAIL VDD2 8.103431f
C10 VDD2 B 3.469556f
C11 VDD1 B 3.441024f
C12 VTAIL B 4.471308f
C13 VN B 6.078691f
C14 VP B 4.629312f
C15 VDD1.n0 B 0.036507f
C16 VDD1.n1 B 0.025484f
C17 VDD1.n2 B 0.013694f
C18 VDD1.n3 B 0.032367f
C19 VDD1.n4 B 0.014499f
C20 VDD1.n5 B 0.025484f
C21 VDD1.n6 B 0.013694f
C22 VDD1.n7 B 0.032367f
C23 VDD1.n8 B 0.014499f
C24 VDD1.n9 B 0.025484f
C25 VDD1.n10 B 0.013694f
C26 VDD1.n11 B 0.024275f
C27 VDD1.n12 B 0.01912f
C28 VDD1.t0 B 0.05275f
C29 VDD1.n13 B 0.117745f
C30 VDD1.n14 B 0.770244f
C31 VDD1.n15 B 0.013694f
C32 VDD1.n16 B 0.014499f
C33 VDD1.n17 B 0.032367f
C34 VDD1.n18 B 0.032367f
C35 VDD1.n19 B 0.014499f
C36 VDD1.n20 B 0.013694f
C37 VDD1.n21 B 0.025484f
C38 VDD1.n22 B 0.025484f
C39 VDD1.n23 B 0.013694f
C40 VDD1.n24 B 0.014499f
C41 VDD1.n25 B 0.032367f
C42 VDD1.n26 B 0.032367f
C43 VDD1.n27 B 0.014499f
C44 VDD1.n28 B 0.013694f
C45 VDD1.n29 B 0.025484f
C46 VDD1.n30 B 0.025484f
C47 VDD1.n31 B 0.013694f
C48 VDD1.n32 B 0.014499f
C49 VDD1.n33 B 0.032367f
C50 VDD1.n34 B 0.071286f
C51 VDD1.n35 B 0.014499f
C52 VDD1.n36 B 0.013694f
C53 VDD1.n37 B 0.057512f
C54 VDD1.n38 B 0.058631f
C55 VDD1.n39 B 0.036507f
C56 VDD1.n40 B 0.025484f
C57 VDD1.n41 B 0.013694f
C58 VDD1.n42 B 0.032367f
C59 VDD1.n43 B 0.014499f
C60 VDD1.n44 B 0.025484f
C61 VDD1.n45 B 0.013694f
C62 VDD1.n46 B 0.032367f
C63 VDD1.n47 B 0.014499f
C64 VDD1.n48 B 0.025484f
C65 VDD1.n49 B 0.013694f
C66 VDD1.n50 B 0.024275f
C67 VDD1.n51 B 0.01912f
C68 VDD1.t1 B 0.05275f
C69 VDD1.n52 B 0.117745f
C70 VDD1.n53 B 0.770244f
C71 VDD1.n54 B 0.013694f
C72 VDD1.n55 B 0.014499f
C73 VDD1.n56 B 0.032367f
C74 VDD1.n57 B 0.032367f
C75 VDD1.n58 B 0.014499f
C76 VDD1.n59 B 0.013694f
C77 VDD1.n60 B 0.025484f
C78 VDD1.n61 B 0.025484f
C79 VDD1.n62 B 0.013694f
C80 VDD1.n63 B 0.014499f
C81 VDD1.n64 B 0.032367f
C82 VDD1.n65 B 0.032367f
C83 VDD1.n66 B 0.014499f
C84 VDD1.n67 B 0.013694f
C85 VDD1.n68 B 0.025484f
C86 VDD1.n69 B 0.025484f
C87 VDD1.n70 B 0.013694f
C88 VDD1.n71 B 0.014499f
C89 VDD1.n72 B 0.032367f
C90 VDD1.n73 B 0.071286f
C91 VDD1.n74 B 0.014499f
C92 VDD1.n75 B 0.013694f
C93 VDD1.n76 B 0.057512f
C94 VDD1.n77 B 0.058344f
C95 VDD1.t4 B 0.149021f
C96 VDD1.t5 B 0.149021f
C97 VDD1.n78 B 1.27201f
C98 VDD1.n79 B 1.56017f
C99 VDD1.t2 B 0.149021f
C100 VDD1.t3 B 0.149021f
C101 VDD1.n80 B 1.27153f
C102 VDD1.n81 B 1.84982f
C103 VP.n0 B 0.041676f
C104 VP.t4 B 0.384617f
C105 VP.t5 B 0.390549f
C106 VP.n1 B 0.165452f
C107 VP.t3 B 0.382523f
C108 VP.n2 B 0.178175f
C109 VP.t2 B 0.384617f
C110 VP.n3 B 0.171071f
C111 VP.n4 B 1.4573f
C112 VP.n5 B 1.40333f
C113 VP.n6 B 0.171071f
C114 VP.t1 B 0.382523f
C115 VP.n7 B 0.178175f
C116 VP.t0 B 0.384617f
C117 VP.n8 B 0.171071f
C118 VP.n9 B 0.032297f
C119 VDD2.n0 B 0.036486f
C120 VDD2.n1 B 0.025469f
C121 VDD2.n2 B 0.013686f
C122 VDD2.n3 B 0.032349f
C123 VDD2.n4 B 0.014491f
C124 VDD2.n5 B 0.025469f
C125 VDD2.n6 B 0.013686f
C126 VDD2.n7 B 0.032349f
C127 VDD2.n8 B 0.014491f
C128 VDD2.n9 B 0.025469f
C129 VDD2.n10 B 0.013686f
C130 VDD2.n11 B 0.024262f
C131 VDD2.n12 B 0.019109f
C132 VDD2.t5 B 0.05272f
C133 VDD2.n13 B 0.117677f
C134 VDD2.n14 B 0.769804f
C135 VDD2.n15 B 0.013686f
C136 VDD2.n16 B 0.014491f
C137 VDD2.n17 B 0.032349f
C138 VDD2.n18 B 0.032349f
C139 VDD2.n19 B 0.014491f
C140 VDD2.n20 B 0.013686f
C141 VDD2.n21 B 0.025469f
C142 VDD2.n22 B 0.025469f
C143 VDD2.n23 B 0.013686f
C144 VDD2.n24 B 0.014491f
C145 VDD2.n25 B 0.032349f
C146 VDD2.n26 B 0.032349f
C147 VDD2.n27 B 0.014491f
C148 VDD2.n28 B 0.013686f
C149 VDD2.n29 B 0.025469f
C150 VDD2.n30 B 0.025469f
C151 VDD2.n31 B 0.013686f
C152 VDD2.n32 B 0.014491f
C153 VDD2.n33 B 0.032349f
C154 VDD2.n34 B 0.071245f
C155 VDD2.n35 B 0.014491f
C156 VDD2.n36 B 0.013686f
C157 VDD2.n37 B 0.057479f
C158 VDD2.n38 B 0.05831f
C159 VDD2.t4 B 0.148936f
C160 VDD2.t3 B 0.148936f
C161 VDD2.n39 B 1.27129f
C162 VDD2.n40 B 1.48841f
C163 VDD2.n41 B 0.036486f
C164 VDD2.n42 B 0.025469f
C165 VDD2.n43 B 0.013686f
C166 VDD2.n44 B 0.032349f
C167 VDD2.n45 B 0.014491f
C168 VDD2.n46 B 0.025469f
C169 VDD2.n47 B 0.013686f
C170 VDD2.n48 B 0.032349f
C171 VDD2.n49 B 0.014491f
C172 VDD2.n50 B 0.025469f
C173 VDD2.n51 B 0.013686f
C174 VDD2.n52 B 0.024262f
C175 VDD2.n53 B 0.019109f
C176 VDD2.t1 B 0.05272f
C177 VDD2.n54 B 0.117677f
C178 VDD2.n55 B 0.769804f
C179 VDD2.n56 B 0.013686f
C180 VDD2.n57 B 0.014491f
C181 VDD2.n58 B 0.032349f
C182 VDD2.n59 B 0.032349f
C183 VDD2.n60 B 0.014491f
C184 VDD2.n61 B 0.013686f
C185 VDD2.n62 B 0.025469f
C186 VDD2.n63 B 0.025469f
C187 VDD2.n64 B 0.013686f
C188 VDD2.n65 B 0.014491f
C189 VDD2.n66 B 0.032349f
C190 VDD2.n67 B 0.032349f
C191 VDD2.n68 B 0.014491f
C192 VDD2.n69 B 0.013686f
C193 VDD2.n70 B 0.025469f
C194 VDD2.n71 B 0.025469f
C195 VDD2.n72 B 0.013686f
C196 VDD2.n73 B 0.014491f
C197 VDD2.n74 B 0.032349f
C198 VDD2.n75 B 0.071245f
C199 VDD2.n76 B 0.014491f
C200 VDD2.n77 B 0.013686f
C201 VDD2.n78 B 0.057479f
C202 VDD2.n79 B 0.057543f
C203 VDD2.n80 B 1.63507f
C204 VDD2.t2 B 0.148936f
C205 VDD2.t0 B 0.148936f
C206 VDD2.n81 B 1.27127f
C207 VTAIL.t10 B 0.127744f
C208 VTAIL.t8 B 0.127744f
C209 VTAIL.n0 B 1.02817f
C210 VTAIL.n1 B 0.284982f
C211 VTAIL.n2 B 0.031295f
C212 VTAIL.n3 B 0.021845f
C213 VTAIL.n4 B 0.011739f
C214 VTAIL.n5 B 0.027746f
C215 VTAIL.n6 B 0.012429f
C216 VTAIL.n7 B 0.021845f
C217 VTAIL.n8 B 0.011739f
C218 VTAIL.n9 B 0.027746f
C219 VTAIL.n10 B 0.012429f
C220 VTAIL.n11 B 0.021845f
C221 VTAIL.n12 B 0.011739f
C222 VTAIL.n13 B 0.020809f
C223 VTAIL.n14 B 0.01639f
C224 VTAIL.t3 B 0.045219f
C225 VTAIL.n15 B 0.100933f
C226 VTAIL.n16 B 0.660272f
C227 VTAIL.n17 B 0.011739f
C228 VTAIL.n18 B 0.012429f
C229 VTAIL.n19 B 0.027746f
C230 VTAIL.n20 B 0.027746f
C231 VTAIL.n21 B 0.012429f
C232 VTAIL.n22 B 0.011739f
C233 VTAIL.n23 B 0.021845f
C234 VTAIL.n24 B 0.021845f
C235 VTAIL.n25 B 0.011739f
C236 VTAIL.n26 B 0.012429f
C237 VTAIL.n27 B 0.027746f
C238 VTAIL.n28 B 0.027746f
C239 VTAIL.n29 B 0.012429f
C240 VTAIL.n30 B 0.011739f
C241 VTAIL.n31 B 0.021845f
C242 VTAIL.n32 B 0.021845f
C243 VTAIL.n33 B 0.011739f
C244 VTAIL.n34 B 0.012429f
C245 VTAIL.n35 B 0.027746f
C246 VTAIL.n36 B 0.061108f
C247 VTAIL.n37 B 0.012429f
C248 VTAIL.n38 B 0.011739f
C249 VTAIL.n39 B 0.0493f
C250 VTAIL.n40 B 0.034262f
C251 VTAIL.n41 B 0.120232f
C252 VTAIL.t4 B 0.127744f
C253 VTAIL.t5 B 0.127744f
C254 VTAIL.n42 B 1.02817f
C255 VTAIL.n43 B 1.09736f
C256 VTAIL.t9 B 0.127744f
C257 VTAIL.t11 B 0.127744f
C258 VTAIL.n44 B 1.02818f
C259 VTAIL.n45 B 1.09735f
C260 VTAIL.n46 B 0.031295f
C261 VTAIL.n47 B 0.021845f
C262 VTAIL.n48 B 0.011739f
C263 VTAIL.n49 B 0.027746f
C264 VTAIL.n50 B 0.012429f
C265 VTAIL.n51 B 0.021845f
C266 VTAIL.n52 B 0.011739f
C267 VTAIL.n53 B 0.027746f
C268 VTAIL.n54 B 0.012429f
C269 VTAIL.n55 B 0.021845f
C270 VTAIL.n56 B 0.011739f
C271 VTAIL.n57 B 0.020809f
C272 VTAIL.n58 B 0.01639f
C273 VTAIL.t7 B 0.045219f
C274 VTAIL.n59 B 0.100933f
C275 VTAIL.n60 B 0.660272f
C276 VTAIL.n61 B 0.011739f
C277 VTAIL.n62 B 0.012429f
C278 VTAIL.n63 B 0.027746f
C279 VTAIL.n64 B 0.027746f
C280 VTAIL.n65 B 0.012429f
C281 VTAIL.n66 B 0.011739f
C282 VTAIL.n67 B 0.021845f
C283 VTAIL.n68 B 0.021845f
C284 VTAIL.n69 B 0.011739f
C285 VTAIL.n70 B 0.012429f
C286 VTAIL.n71 B 0.027746f
C287 VTAIL.n72 B 0.027746f
C288 VTAIL.n73 B 0.012429f
C289 VTAIL.n74 B 0.011739f
C290 VTAIL.n75 B 0.021845f
C291 VTAIL.n76 B 0.021845f
C292 VTAIL.n77 B 0.011739f
C293 VTAIL.n78 B 0.012429f
C294 VTAIL.n79 B 0.027746f
C295 VTAIL.n80 B 0.061108f
C296 VTAIL.n81 B 0.012429f
C297 VTAIL.n82 B 0.011739f
C298 VTAIL.n83 B 0.0493f
C299 VTAIL.n84 B 0.034262f
C300 VTAIL.n85 B 0.120232f
C301 VTAIL.t0 B 0.127744f
C302 VTAIL.t2 B 0.127744f
C303 VTAIL.n86 B 1.02818f
C304 VTAIL.n87 B 0.315467f
C305 VTAIL.n88 B 0.031295f
C306 VTAIL.n89 B 0.021845f
C307 VTAIL.n90 B 0.011739f
C308 VTAIL.n91 B 0.027746f
C309 VTAIL.n92 B 0.012429f
C310 VTAIL.n93 B 0.021845f
C311 VTAIL.n94 B 0.011739f
C312 VTAIL.n95 B 0.027746f
C313 VTAIL.n96 B 0.012429f
C314 VTAIL.n97 B 0.021845f
C315 VTAIL.n98 B 0.011739f
C316 VTAIL.n99 B 0.020809f
C317 VTAIL.n100 B 0.01639f
C318 VTAIL.t1 B 0.045219f
C319 VTAIL.n101 B 0.100933f
C320 VTAIL.n102 B 0.660272f
C321 VTAIL.n103 B 0.011739f
C322 VTAIL.n104 B 0.012429f
C323 VTAIL.n105 B 0.027746f
C324 VTAIL.n106 B 0.027746f
C325 VTAIL.n107 B 0.012429f
C326 VTAIL.n108 B 0.011739f
C327 VTAIL.n109 B 0.021845f
C328 VTAIL.n110 B 0.021845f
C329 VTAIL.n111 B 0.011739f
C330 VTAIL.n112 B 0.012429f
C331 VTAIL.n113 B 0.027746f
C332 VTAIL.n114 B 0.027746f
C333 VTAIL.n115 B 0.012429f
C334 VTAIL.n116 B 0.011739f
C335 VTAIL.n117 B 0.021845f
C336 VTAIL.n118 B 0.021845f
C337 VTAIL.n119 B 0.011739f
C338 VTAIL.n120 B 0.012429f
C339 VTAIL.n121 B 0.027746f
C340 VTAIL.n122 B 0.061108f
C341 VTAIL.n123 B 0.012429f
C342 VTAIL.n124 B 0.011739f
C343 VTAIL.n125 B 0.0493f
C344 VTAIL.n126 B 0.034262f
C345 VTAIL.n127 B 0.856f
C346 VTAIL.n128 B 0.031295f
C347 VTAIL.n129 B 0.021845f
C348 VTAIL.n130 B 0.011739f
C349 VTAIL.n131 B 0.027746f
C350 VTAIL.n132 B 0.012429f
C351 VTAIL.n133 B 0.021845f
C352 VTAIL.n134 B 0.011739f
C353 VTAIL.n135 B 0.027746f
C354 VTAIL.n136 B 0.012429f
C355 VTAIL.n137 B 0.021845f
C356 VTAIL.n138 B 0.011739f
C357 VTAIL.n139 B 0.020809f
C358 VTAIL.n140 B 0.01639f
C359 VTAIL.t6 B 0.045219f
C360 VTAIL.n141 B 0.100933f
C361 VTAIL.n142 B 0.660272f
C362 VTAIL.n143 B 0.011739f
C363 VTAIL.n144 B 0.012429f
C364 VTAIL.n145 B 0.027746f
C365 VTAIL.n146 B 0.027746f
C366 VTAIL.n147 B 0.012429f
C367 VTAIL.n148 B 0.011739f
C368 VTAIL.n149 B 0.021845f
C369 VTAIL.n150 B 0.021845f
C370 VTAIL.n151 B 0.011739f
C371 VTAIL.n152 B 0.012429f
C372 VTAIL.n153 B 0.027746f
C373 VTAIL.n154 B 0.027746f
C374 VTAIL.n155 B 0.012429f
C375 VTAIL.n156 B 0.011739f
C376 VTAIL.n157 B 0.021845f
C377 VTAIL.n158 B 0.021845f
C378 VTAIL.n159 B 0.011739f
C379 VTAIL.n160 B 0.012429f
C380 VTAIL.n161 B 0.027746f
C381 VTAIL.n162 B 0.061108f
C382 VTAIL.n163 B 0.012429f
C383 VTAIL.n164 B 0.011739f
C384 VTAIL.n165 B 0.0493f
C385 VTAIL.n166 B 0.034262f
C386 VTAIL.n167 B 0.840374f
C387 VN.t0 B 0.380808f
C388 VN.n0 B 0.161326f
C389 VN.t1 B 0.372983f
C390 VN.n1 B 0.173732f
C391 VN.t2 B 0.375025f
C392 VN.n2 B 0.166804f
C393 VN.n3 B 0.123733f
C394 VN.t5 B 0.380808f
C395 VN.n4 B 0.161326f
C396 VN.t4 B 0.375025f
C397 VN.t3 B 0.372983f
C398 VN.n5 B 0.173732f
C399 VN.n6 B 0.166804f
C400 VN.n7 B 1.44786f
.ends

