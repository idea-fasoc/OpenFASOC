* NGSPICE file created from diff_pair_sample_0673.ext - technology: sky130A

.subckt diff_pair_sample_0673 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=3.17625 pd=19.58 as=3.17625 ps=19.58 w=19.25 l=2.57
X1 VDD2.t9 VN.t0 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=7.5075 pd=39.28 as=3.17625 ps=19.58 w=19.25 l=2.57
X2 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=7.5075 pd=39.28 as=0 ps=0 w=19.25 l=2.57
X3 VTAIL.t18 VP.t1 VDD1.t4 B.t9 sky130_fd_pr__nfet_01v8 ad=3.17625 pd=19.58 as=3.17625 ps=19.58 w=19.25 l=2.57
X4 VDD2.t8 VN.t1 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=3.17625 pd=19.58 as=3.17625 ps=19.58 w=19.25 l=2.57
X5 VDD2.t7 VN.t2 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=3.17625 pd=19.58 as=3.17625 ps=19.58 w=19.25 l=2.57
X6 VTAIL.t9 VN.t3 VDD2.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=3.17625 pd=19.58 as=3.17625 ps=19.58 w=19.25 l=2.57
X7 VTAIL.t17 VP.t2 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=3.17625 pd=19.58 as=3.17625 ps=19.58 w=19.25 l=2.57
X8 VDD2.t5 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=7.5075 pd=39.28 as=3.17625 ps=19.58 w=19.25 l=2.57
X9 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=7.5075 pd=39.28 as=0 ps=0 w=19.25 l=2.57
X10 VTAIL.t3 VN.t5 VDD2.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.17625 pd=19.58 as=3.17625 ps=19.58 w=19.25 l=2.57
X11 VDD1.t2 VP.t3 VTAIL.t16 B.t0 sky130_fd_pr__nfet_01v8 ad=7.5075 pd=39.28 as=3.17625 ps=19.58 w=19.25 l=2.57
X12 VDD2.t3 VN.t6 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.17625 pd=19.58 as=7.5075 ps=39.28 w=19.25 l=2.57
X13 VDD1.t1 VP.t4 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=3.17625 pd=19.58 as=3.17625 ps=19.58 w=19.25 l=2.57
X14 VTAIL.t5 VN.t7 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=3.17625 pd=19.58 as=3.17625 ps=19.58 w=19.25 l=2.57
X15 VTAIL.t1 VN.t8 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.17625 pd=19.58 as=3.17625 ps=19.58 w=19.25 l=2.57
X16 VDD2.t0 VN.t9 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.17625 pd=19.58 as=7.5075 ps=39.28 w=19.25 l=2.57
X17 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=7.5075 pd=39.28 as=0 ps=0 w=19.25 l=2.57
X18 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.5075 pd=39.28 as=0 ps=0 w=19.25 l=2.57
X19 VDD1.t0 VP.t5 VTAIL.t14 B.t2 sky130_fd_pr__nfet_01v8 ad=3.17625 pd=19.58 as=7.5075 ps=39.28 w=19.25 l=2.57
X20 VTAIL.t13 VP.t6 VDD1.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=3.17625 pd=19.58 as=3.17625 ps=19.58 w=19.25 l=2.57
X21 VDD1.t8 VP.t7 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=3.17625 pd=19.58 as=3.17625 ps=19.58 w=19.25 l=2.57
X22 VDD1.t7 VP.t8 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=3.17625 pd=19.58 as=7.5075 ps=39.28 w=19.25 l=2.57
X23 VDD1.t6 VP.t9 VTAIL.t10 B.t8 sky130_fd_pr__nfet_01v8 ad=7.5075 pd=39.28 as=3.17625 ps=19.58 w=19.25 l=2.57
R0 VP.n24 VP.t3 211.549
R1 VP.n56 VP.t9 180.517
R2 VP.n64 VP.t2 180.517
R3 VP.n76 VP.t4 180.517
R4 VP.n3 VP.t6 180.517
R5 VP.n95 VP.t8 180.517
R6 VP.n53 VP.t5 180.517
R7 VP.n16 VP.t0 180.517
R8 VP.n34 VP.t7 180.517
R9 VP.n23 VP.t1 180.517
R10 VP.n25 VP.n22 161.3
R11 VP.n27 VP.n26 161.3
R12 VP.n28 VP.n21 161.3
R13 VP.n30 VP.n29 161.3
R14 VP.n31 VP.n20 161.3
R15 VP.n33 VP.n32 161.3
R16 VP.n35 VP.n19 161.3
R17 VP.n37 VP.n36 161.3
R18 VP.n38 VP.n18 161.3
R19 VP.n40 VP.n39 161.3
R20 VP.n41 VP.n17 161.3
R21 VP.n43 VP.n42 161.3
R22 VP.n45 VP.n44 161.3
R23 VP.n46 VP.n15 161.3
R24 VP.n48 VP.n47 161.3
R25 VP.n49 VP.n14 161.3
R26 VP.n51 VP.n50 161.3
R27 VP.n52 VP.n13 161.3
R28 VP.n94 VP.n0 161.3
R29 VP.n93 VP.n92 161.3
R30 VP.n91 VP.n1 161.3
R31 VP.n90 VP.n89 161.3
R32 VP.n88 VP.n2 161.3
R33 VP.n87 VP.n86 161.3
R34 VP.n85 VP.n84 161.3
R35 VP.n83 VP.n4 161.3
R36 VP.n82 VP.n81 161.3
R37 VP.n80 VP.n5 161.3
R38 VP.n79 VP.n78 161.3
R39 VP.n77 VP.n6 161.3
R40 VP.n75 VP.n74 161.3
R41 VP.n73 VP.n7 161.3
R42 VP.n72 VP.n71 161.3
R43 VP.n70 VP.n8 161.3
R44 VP.n69 VP.n68 161.3
R45 VP.n67 VP.n9 161.3
R46 VP.n66 VP.n65 161.3
R47 VP.n63 VP.n10 161.3
R48 VP.n62 VP.n61 161.3
R49 VP.n60 VP.n11 161.3
R50 VP.n59 VP.n58 161.3
R51 VP.n57 VP.n12 161.3
R52 VP.n56 VP.n55 108.309
R53 VP.n96 VP.n95 108.309
R54 VP.n54 VP.n53 108.309
R55 VP.n24 VP.n23 65.3454
R56 VP.n55 VP.n54 58.3405
R57 VP.n71 VP.n70 56.5193
R58 VP.n82 VP.n5 56.5193
R59 VP.n40 VP.n18 56.5193
R60 VP.n29 VP.n28 56.5193
R61 VP.n62 VP.n11 50.2061
R62 VP.n89 VP.n1 50.2061
R63 VP.n47 VP.n14 50.2061
R64 VP.n63 VP.n62 30.7807
R65 VP.n89 VP.n88 30.7807
R66 VP.n47 VP.n46 30.7807
R67 VP.n58 VP.n57 24.4675
R68 VP.n58 VP.n11 24.4675
R69 VP.n65 VP.n63 24.4675
R70 VP.n69 VP.n9 24.4675
R71 VP.n70 VP.n69 24.4675
R72 VP.n71 VP.n7 24.4675
R73 VP.n75 VP.n7 24.4675
R74 VP.n78 VP.n77 24.4675
R75 VP.n78 VP.n5 24.4675
R76 VP.n83 VP.n82 24.4675
R77 VP.n84 VP.n83 24.4675
R78 VP.n88 VP.n87 24.4675
R79 VP.n93 VP.n1 24.4675
R80 VP.n94 VP.n93 24.4675
R81 VP.n51 VP.n14 24.4675
R82 VP.n52 VP.n51 24.4675
R83 VP.n41 VP.n40 24.4675
R84 VP.n42 VP.n41 24.4675
R85 VP.n46 VP.n45 24.4675
R86 VP.n29 VP.n20 24.4675
R87 VP.n33 VP.n20 24.4675
R88 VP.n36 VP.n35 24.4675
R89 VP.n36 VP.n18 24.4675
R90 VP.n27 VP.n22 24.4675
R91 VP.n28 VP.n27 24.4675
R92 VP.n65 VP.n64 17.1274
R93 VP.n87 VP.n3 17.1274
R94 VP.n45 VP.n16 17.1274
R95 VP.n76 VP.n75 12.234
R96 VP.n77 VP.n76 12.234
R97 VP.n34 VP.n33 12.234
R98 VP.n35 VP.n34 12.234
R99 VP.n64 VP.n9 7.3406
R100 VP.n84 VP.n3 7.3406
R101 VP.n42 VP.n16 7.3406
R102 VP.n23 VP.n22 7.3406
R103 VP.n25 VP.n24 7.32785
R104 VP.n57 VP.n56 2.4472
R105 VP.n95 VP.n94 2.4472
R106 VP.n53 VP.n52 2.4472
R107 VP.n54 VP.n13 0.278367
R108 VP.n55 VP.n12 0.278367
R109 VP.n96 VP.n0 0.278367
R110 VP.n26 VP.n25 0.189894
R111 VP.n26 VP.n21 0.189894
R112 VP.n30 VP.n21 0.189894
R113 VP.n31 VP.n30 0.189894
R114 VP.n32 VP.n31 0.189894
R115 VP.n32 VP.n19 0.189894
R116 VP.n37 VP.n19 0.189894
R117 VP.n38 VP.n37 0.189894
R118 VP.n39 VP.n38 0.189894
R119 VP.n39 VP.n17 0.189894
R120 VP.n43 VP.n17 0.189894
R121 VP.n44 VP.n43 0.189894
R122 VP.n44 VP.n15 0.189894
R123 VP.n48 VP.n15 0.189894
R124 VP.n49 VP.n48 0.189894
R125 VP.n50 VP.n49 0.189894
R126 VP.n50 VP.n13 0.189894
R127 VP.n59 VP.n12 0.189894
R128 VP.n60 VP.n59 0.189894
R129 VP.n61 VP.n60 0.189894
R130 VP.n61 VP.n10 0.189894
R131 VP.n66 VP.n10 0.189894
R132 VP.n67 VP.n66 0.189894
R133 VP.n68 VP.n67 0.189894
R134 VP.n68 VP.n8 0.189894
R135 VP.n72 VP.n8 0.189894
R136 VP.n73 VP.n72 0.189894
R137 VP.n74 VP.n73 0.189894
R138 VP.n74 VP.n6 0.189894
R139 VP.n79 VP.n6 0.189894
R140 VP.n80 VP.n79 0.189894
R141 VP.n81 VP.n80 0.189894
R142 VP.n81 VP.n4 0.189894
R143 VP.n85 VP.n4 0.189894
R144 VP.n86 VP.n85 0.189894
R145 VP.n86 VP.n2 0.189894
R146 VP.n90 VP.n2 0.189894
R147 VP.n91 VP.n90 0.189894
R148 VP.n92 VP.n91 0.189894
R149 VP.n92 VP.n0 0.189894
R150 VP VP.n96 0.153454
R151 VDD1.n1 VDD1.t2 62.7821
R152 VDD1.n3 VDD1.t6 62.7819
R153 VDD1.n5 VDD1.n4 61.0732
R154 VDD1.n1 VDD1.n0 59.2536
R155 VDD1.n3 VDD1.n2 59.2535
R156 VDD1.n7 VDD1.n6 59.2534
R157 VDD1.n7 VDD1.n5 54.0181
R158 VDD1 VDD1.n7 1.81731
R159 VDD1.n6 VDD1.t5 1.02907
R160 VDD1.n6 VDD1.t0 1.02907
R161 VDD1.n0 VDD1.t4 1.02907
R162 VDD1.n0 VDD1.t8 1.02907
R163 VDD1.n4 VDD1.t9 1.02907
R164 VDD1.n4 VDD1.t7 1.02907
R165 VDD1.n2 VDD1.t3 1.02907
R166 VDD1.n2 VDD1.t1 1.02907
R167 VDD1 VDD1.n1 0.68369
R168 VDD1.n5 VDD1.n3 0.570154
R169 VTAIL.n11 VTAIL.t4 43.6033
R170 VTAIL.n17 VTAIL.t2 43.6031
R171 VTAIL.n2 VTAIL.t11 43.6031
R172 VTAIL.n16 VTAIL.t14 43.6031
R173 VTAIL.n15 VTAIL.n14 42.5748
R174 VTAIL.n13 VTAIL.n12 42.5748
R175 VTAIL.n10 VTAIL.n9 42.5748
R176 VTAIL.n8 VTAIL.n7 42.5748
R177 VTAIL.n19 VTAIL.n18 42.5747
R178 VTAIL.n1 VTAIL.n0 42.5747
R179 VTAIL.n4 VTAIL.n3 42.5747
R180 VTAIL.n6 VTAIL.n5 42.5747
R181 VTAIL.n8 VTAIL.n6 33.9617
R182 VTAIL.n17 VTAIL.n16 31.4617
R183 VTAIL.n10 VTAIL.n8 2.5005
R184 VTAIL.n11 VTAIL.n10 2.5005
R185 VTAIL.n15 VTAIL.n13 2.5005
R186 VTAIL.n16 VTAIL.n15 2.5005
R187 VTAIL.n6 VTAIL.n4 2.5005
R188 VTAIL.n4 VTAIL.n2 2.5005
R189 VTAIL.n19 VTAIL.n17 2.5005
R190 VTAIL VTAIL.n1 1.93369
R191 VTAIL.n13 VTAIL.n11 1.72033
R192 VTAIL.n2 VTAIL.n1 1.72033
R193 VTAIL.n18 VTAIL.t6 1.02907
R194 VTAIL.n18 VTAIL.t1 1.02907
R195 VTAIL.n0 VTAIL.t0 1.02907
R196 VTAIL.n0 VTAIL.t9 1.02907
R197 VTAIL.n3 VTAIL.t15 1.02907
R198 VTAIL.n3 VTAIL.t13 1.02907
R199 VTAIL.n5 VTAIL.t10 1.02907
R200 VTAIL.n5 VTAIL.t17 1.02907
R201 VTAIL.n14 VTAIL.t12 1.02907
R202 VTAIL.n14 VTAIL.t19 1.02907
R203 VTAIL.n12 VTAIL.t16 1.02907
R204 VTAIL.n12 VTAIL.t18 1.02907
R205 VTAIL.n9 VTAIL.t7 1.02907
R206 VTAIL.n9 VTAIL.t3 1.02907
R207 VTAIL.n7 VTAIL.t8 1.02907
R208 VTAIL.n7 VTAIL.t5 1.02907
R209 VTAIL VTAIL.n19 0.56731
R210 B.n1161 B.n1160 585
R211 B.n1162 B.n1161 585
R212 B.n447 B.n177 585
R213 B.n446 B.n445 585
R214 B.n444 B.n443 585
R215 B.n442 B.n441 585
R216 B.n440 B.n439 585
R217 B.n438 B.n437 585
R218 B.n436 B.n435 585
R219 B.n434 B.n433 585
R220 B.n432 B.n431 585
R221 B.n430 B.n429 585
R222 B.n428 B.n427 585
R223 B.n426 B.n425 585
R224 B.n424 B.n423 585
R225 B.n422 B.n421 585
R226 B.n420 B.n419 585
R227 B.n418 B.n417 585
R228 B.n416 B.n415 585
R229 B.n414 B.n413 585
R230 B.n412 B.n411 585
R231 B.n410 B.n409 585
R232 B.n408 B.n407 585
R233 B.n406 B.n405 585
R234 B.n404 B.n403 585
R235 B.n402 B.n401 585
R236 B.n400 B.n399 585
R237 B.n398 B.n397 585
R238 B.n396 B.n395 585
R239 B.n394 B.n393 585
R240 B.n392 B.n391 585
R241 B.n390 B.n389 585
R242 B.n388 B.n387 585
R243 B.n386 B.n385 585
R244 B.n384 B.n383 585
R245 B.n382 B.n381 585
R246 B.n380 B.n379 585
R247 B.n378 B.n377 585
R248 B.n376 B.n375 585
R249 B.n374 B.n373 585
R250 B.n372 B.n371 585
R251 B.n370 B.n369 585
R252 B.n368 B.n367 585
R253 B.n366 B.n365 585
R254 B.n364 B.n363 585
R255 B.n362 B.n361 585
R256 B.n360 B.n359 585
R257 B.n358 B.n357 585
R258 B.n356 B.n355 585
R259 B.n354 B.n353 585
R260 B.n352 B.n351 585
R261 B.n350 B.n349 585
R262 B.n348 B.n347 585
R263 B.n346 B.n345 585
R264 B.n344 B.n343 585
R265 B.n342 B.n341 585
R266 B.n340 B.n339 585
R267 B.n338 B.n337 585
R268 B.n336 B.n335 585
R269 B.n334 B.n333 585
R270 B.n332 B.n331 585
R271 B.n330 B.n329 585
R272 B.n328 B.n327 585
R273 B.n326 B.n325 585
R274 B.n324 B.n323 585
R275 B.n322 B.n321 585
R276 B.n320 B.n319 585
R277 B.n318 B.n317 585
R278 B.n316 B.n315 585
R279 B.n314 B.n313 585
R280 B.n312 B.n311 585
R281 B.n310 B.n309 585
R282 B.n308 B.n307 585
R283 B.n305 B.n304 585
R284 B.n303 B.n302 585
R285 B.n301 B.n300 585
R286 B.n299 B.n298 585
R287 B.n297 B.n296 585
R288 B.n295 B.n294 585
R289 B.n293 B.n292 585
R290 B.n291 B.n290 585
R291 B.n289 B.n288 585
R292 B.n287 B.n286 585
R293 B.n285 B.n284 585
R294 B.n283 B.n282 585
R295 B.n281 B.n280 585
R296 B.n279 B.n278 585
R297 B.n277 B.n276 585
R298 B.n275 B.n274 585
R299 B.n273 B.n272 585
R300 B.n271 B.n270 585
R301 B.n269 B.n268 585
R302 B.n267 B.n266 585
R303 B.n265 B.n264 585
R304 B.n263 B.n262 585
R305 B.n261 B.n260 585
R306 B.n259 B.n258 585
R307 B.n257 B.n256 585
R308 B.n255 B.n254 585
R309 B.n253 B.n252 585
R310 B.n251 B.n250 585
R311 B.n249 B.n248 585
R312 B.n247 B.n246 585
R313 B.n245 B.n244 585
R314 B.n243 B.n242 585
R315 B.n241 B.n240 585
R316 B.n239 B.n238 585
R317 B.n237 B.n236 585
R318 B.n235 B.n234 585
R319 B.n233 B.n232 585
R320 B.n231 B.n230 585
R321 B.n229 B.n228 585
R322 B.n227 B.n226 585
R323 B.n225 B.n224 585
R324 B.n223 B.n222 585
R325 B.n221 B.n220 585
R326 B.n219 B.n218 585
R327 B.n217 B.n216 585
R328 B.n215 B.n214 585
R329 B.n213 B.n212 585
R330 B.n211 B.n210 585
R331 B.n209 B.n208 585
R332 B.n207 B.n206 585
R333 B.n205 B.n204 585
R334 B.n203 B.n202 585
R335 B.n201 B.n200 585
R336 B.n199 B.n198 585
R337 B.n197 B.n196 585
R338 B.n195 B.n194 585
R339 B.n193 B.n192 585
R340 B.n191 B.n190 585
R341 B.n189 B.n188 585
R342 B.n187 B.n186 585
R343 B.n185 B.n184 585
R344 B.n110 B.n109 585
R345 B.n1165 B.n1164 585
R346 B.n1159 B.n178 585
R347 B.n178 B.n107 585
R348 B.n1158 B.n106 585
R349 B.n1169 B.n106 585
R350 B.n1157 B.n105 585
R351 B.n1170 B.n105 585
R352 B.n1156 B.n104 585
R353 B.n1171 B.n104 585
R354 B.n1155 B.n1154 585
R355 B.n1154 B.n100 585
R356 B.n1153 B.n99 585
R357 B.n1177 B.n99 585
R358 B.n1152 B.n98 585
R359 B.n1178 B.n98 585
R360 B.n1151 B.n97 585
R361 B.n1179 B.n97 585
R362 B.n1150 B.n1149 585
R363 B.n1149 B.n93 585
R364 B.n1148 B.n92 585
R365 B.n1185 B.n92 585
R366 B.n1147 B.n91 585
R367 B.n1186 B.n91 585
R368 B.n1146 B.n90 585
R369 B.n1187 B.n90 585
R370 B.n1145 B.n1144 585
R371 B.n1144 B.n86 585
R372 B.n1143 B.n85 585
R373 B.n1193 B.n85 585
R374 B.n1142 B.n84 585
R375 B.n1194 B.n84 585
R376 B.n1141 B.n83 585
R377 B.n1195 B.n83 585
R378 B.n1140 B.n1139 585
R379 B.n1139 B.n79 585
R380 B.n1138 B.n78 585
R381 B.n1201 B.n78 585
R382 B.n1137 B.n77 585
R383 B.n1202 B.n77 585
R384 B.n1136 B.n76 585
R385 B.n1203 B.n76 585
R386 B.n1135 B.n1134 585
R387 B.n1134 B.n72 585
R388 B.n1133 B.n71 585
R389 B.n1209 B.n71 585
R390 B.n1132 B.n70 585
R391 B.n1210 B.n70 585
R392 B.n1131 B.n69 585
R393 B.n1211 B.n69 585
R394 B.n1130 B.n1129 585
R395 B.n1129 B.n65 585
R396 B.n1128 B.n64 585
R397 B.n1217 B.n64 585
R398 B.n1127 B.n63 585
R399 B.n1218 B.n63 585
R400 B.n1126 B.n62 585
R401 B.n1219 B.n62 585
R402 B.n1125 B.n1124 585
R403 B.n1124 B.n61 585
R404 B.n1123 B.n57 585
R405 B.n1225 B.n57 585
R406 B.n1122 B.n56 585
R407 B.n1226 B.n56 585
R408 B.n1121 B.n55 585
R409 B.n1227 B.n55 585
R410 B.n1120 B.n1119 585
R411 B.n1119 B.n51 585
R412 B.n1118 B.n50 585
R413 B.n1233 B.n50 585
R414 B.n1117 B.n49 585
R415 B.n1234 B.n49 585
R416 B.n1116 B.n48 585
R417 B.n1235 B.n48 585
R418 B.n1115 B.n1114 585
R419 B.n1114 B.n47 585
R420 B.n1113 B.n43 585
R421 B.n1241 B.n43 585
R422 B.n1112 B.n42 585
R423 B.n1242 B.n42 585
R424 B.n1111 B.n41 585
R425 B.n1243 B.n41 585
R426 B.n1110 B.n1109 585
R427 B.n1109 B.n37 585
R428 B.n1108 B.n36 585
R429 B.n1249 B.n36 585
R430 B.n1107 B.n35 585
R431 B.n1250 B.n35 585
R432 B.n1106 B.n34 585
R433 B.n1251 B.n34 585
R434 B.n1105 B.n1104 585
R435 B.n1104 B.n30 585
R436 B.n1103 B.n29 585
R437 B.n1257 B.n29 585
R438 B.n1102 B.n28 585
R439 B.n1258 B.n28 585
R440 B.n1101 B.n27 585
R441 B.n1259 B.n27 585
R442 B.n1100 B.n1099 585
R443 B.n1099 B.n23 585
R444 B.n1098 B.n22 585
R445 B.n1265 B.n22 585
R446 B.n1097 B.n21 585
R447 B.n1266 B.n21 585
R448 B.n1096 B.n20 585
R449 B.n1267 B.n20 585
R450 B.n1095 B.n1094 585
R451 B.n1094 B.n16 585
R452 B.n1093 B.n15 585
R453 B.n1273 B.n15 585
R454 B.n1092 B.n14 585
R455 B.n1274 B.n14 585
R456 B.n1091 B.n13 585
R457 B.n1275 B.n13 585
R458 B.n1090 B.n1089 585
R459 B.n1089 B.n12 585
R460 B.n1088 B.n1087 585
R461 B.n1088 B.n8 585
R462 B.n1086 B.n7 585
R463 B.n1282 B.n7 585
R464 B.n1085 B.n6 585
R465 B.n1283 B.n6 585
R466 B.n1084 B.n5 585
R467 B.n1284 B.n5 585
R468 B.n1083 B.n1082 585
R469 B.n1082 B.n4 585
R470 B.n1081 B.n448 585
R471 B.n1081 B.n1080 585
R472 B.n1071 B.n449 585
R473 B.n450 B.n449 585
R474 B.n1073 B.n1072 585
R475 B.n1074 B.n1073 585
R476 B.n1070 B.n455 585
R477 B.n455 B.n454 585
R478 B.n1069 B.n1068 585
R479 B.n1068 B.n1067 585
R480 B.n457 B.n456 585
R481 B.n458 B.n457 585
R482 B.n1060 B.n1059 585
R483 B.n1061 B.n1060 585
R484 B.n1058 B.n463 585
R485 B.n463 B.n462 585
R486 B.n1057 B.n1056 585
R487 B.n1056 B.n1055 585
R488 B.n465 B.n464 585
R489 B.n466 B.n465 585
R490 B.n1048 B.n1047 585
R491 B.n1049 B.n1048 585
R492 B.n1046 B.n471 585
R493 B.n471 B.n470 585
R494 B.n1045 B.n1044 585
R495 B.n1044 B.n1043 585
R496 B.n473 B.n472 585
R497 B.n474 B.n473 585
R498 B.n1036 B.n1035 585
R499 B.n1037 B.n1036 585
R500 B.n1034 B.n479 585
R501 B.n479 B.n478 585
R502 B.n1033 B.n1032 585
R503 B.n1032 B.n1031 585
R504 B.n481 B.n480 585
R505 B.n482 B.n481 585
R506 B.n1024 B.n1023 585
R507 B.n1025 B.n1024 585
R508 B.n1022 B.n487 585
R509 B.n487 B.n486 585
R510 B.n1021 B.n1020 585
R511 B.n1020 B.n1019 585
R512 B.n489 B.n488 585
R513 B.n1012 B.n489 585
R514 B.n1011 B.n1010 585
R515 B.n1013 B.n1011 585
R516 B.n1009 B.n494 585
R517 B.n494 B.n493 585
R518 B.n1008 B.n1007 585
R519 B.n1007 B.n1006 585
R520 B.n496 B.n495 585
R521 B.n497 B.n496 585
R522 B.n999 B.n998 585
R523 B.n1000 B.n999 585
R524 B.n997 B.n502 585
R525 B.n502 B.n501 585
R526 B.n996 B.n995 585
R527 B.n995 B.n994 585
R528 B.n504 B.n503 585
R529 B.n987 B.n504 585
R530 B.n986 B.n985 585
R531 B.n988 B.n986 585
R532 B.n984 B.n509 585
R533 B.n509 B.n508 585
R534 B.n983 B.n982 585
R535 B.n982 B.n981 585
R536 B.n511 B.n510 585
R537 B.n512 B.n511 585
R538 B.n974 B.n973 585
R539 B.n975 B.n974 585
R540 B.n972 B.n517 585
R541 B.n517 B.n516 585
R542 B.n971 B.n970 585
R543 B.n970 B.n969 585
R544 B.n519 B.n518 585
R545 B.n520 B.n519 585
R546 B.n962 B.n961 585
R547 B.n963 B.n962 585
R548 B.n960 B.n525 585
R549 B.n525 B.n524 585
R550 B.n959 B.n958 585
R551 B.n958 B.n957 585
R552 B.n527 B.n526 585
R553 B.n528 B.n527 585
R554 B.n950 B.n949 585
R555 B.n951 B.n950 585
R556 B.n948 B.n533 585
R557 B.n533 B.n532 585
R558 B.n947 B.n946 585
R559 B.n946 B.n945 585
R560 B.n535 B.n534 585
R561 B.n536 B.n535 585
R562 B.n938 B.n937 585
R563 B.n939 B.n938 585
R564 B.n936 B.n541 585
R565 B.n541 B.n540 585
R566 B.n935 B.n934 585
R567 B.n934 B.n933 585
R568 B.n543 B.n542 585
R569 B.n544 B.n543 585
R570 B.n926 B.n925 585
R571 B.n927 B.n926 585
R572 B.n924 B.n549 585
R573 B.n549 B.n548 585
R574 B.n923 B.n922 585
R575 B.n922 B.n921 585
R576 B.n551 B.n550 585
R577 B.n552 B.n551 585
R578 B.n914 B.n913 585
R579 B.n915 B.n914 585
R580 B.n912 B.n557 585
R581 B.n557 B.n556 585
R582 B.n911 B.n910 585
R583 B.n910 B.n909 585
R584 B.n559 B.n558 585
R585 B.n560 B.n559 585
R586 B.n905 B.n904 585
R587 B.n563 B.n562 585
R588 B.n901 B.n900 585
R589 B.n902 B.n901 585
R590 B.n899 B.n630 585
R591 B.n898 B.n897 585
R592 B.n896 B.n895 585
R593 B.n894 B.n893 585
R594 B.n892 B.n891 585
R595 B.n890 B.n889 585
R596 B.n888 B.n887 585
R597 B.n886 B.n885 585
R598 B.n884 B.n883 585
R599 B.n882 B.n881 585
R600 B.n880 B.n879 585
R601 B.n878 B.n877 585
R602 B.n876 B.n875 585
R603 B.n874 B.n873 585
R604 B.n872 B.n871 585
R605 B.n870 B.n869 585
R606 B.n868 B.n867 585
R607 B.n866 B.n865 585
R608 B.n864 B.n863 585
R609 B.n862 B.n861 585
R610 B.n860 B.n859 585
R611 B.n858 B.n857 585
R612 B.n856 B.n855 585
R613 B.n854 B.n853 585
R614 B.n852 B.n851 585
R615 B.n850 B.n849 585
R616 B.n848 B.n847 585
R617 B.n846 B.n845 585
R618 B.n844 B.n843 585
R619 B.n842 B.n841 585
R620 B.n840 B.n839 585
R621 B.n838 B.n837 585
R622 B.n836 B.n835 585
R623 B.n834 B.n833 585
R624 B.n832 B.n831 585
R625 B.n830 B.n829 585
R626 B.n828 B.n827 585
R627 B.n826 B.n825 585
R628 B.n824 B.n823 585
R629 B.n822 B.n821 585
R630 B.n820 B.n819 585
R631 B.n818 B.n817 585
R632 B.n816 B.n815 585
R633 B.n814 B.n813 585
R634 B.n812 B.n811 585
R635 B.n810 B.n809 585
R636 B.n808 B.n807 585
R637 B.n806 B.n805 585
R638 B.n804 B.n803 585
R639 B.n802 B.n801 585
R640 B.n800 B.n799 585
R641 B.n798 B.n797 585
R642 B.n796 B.n795 585
R643 B.n794 B.n793 585
R644 B.n792 B.n791 585
R645 B.n790 B.n789 585
R646 B.n788 B.n787 585
R647 B.n786 B.n785 585
R648 B.n784 B.n783 585
R649 B.n782 B.n781 585
R650 B.n780 B.n779 585
R651 B.n778 B.n777 585
R652 B.n776 B.n775 585
R653 B.n774 B.n773 585
R654 B.n772 B.n771 585
R655 B.n770 B.n769 585
R656 B.n768 B.n767 585
R657 B.n766 B.n765 585
R658 B.n764 B.n763 585
R659 B.n761 B.n760 585
R660 B.n759 B.n758 585
R661 B.n757 B.n756 585
R662 B.n755 B.n754 585
R663 B.n753 B.n752 585
R664 B.n751 B.n750 585
R665 B.n749 B.n748 585
R666 B.n747 B.n746 585
R667 B.n745 B.n744 585
R668 B.n743 B.n742 585
R669 B.n741 B.n740 585
R670 B.n739 B.n738 585
R671 B.n737 B.n736 585
R672 B.n735 B.n734 585
R673 B.n733 B.n732 585
R674 B.n731 B.n730 585
R675 B.n729 B.n728 585
R676 B.n727 B.n726 585
R677 B.n725 B.n724 585
R678 B.n723 B.n722 585
R679 B.n721 B.n720 585
R680 B.n719 B.n718 585
R681 B.n717 B.n716 585
R682 B.n715 B.n714 585
R683 B.n713 B.n712 585
R684 B.n711 B.n710 585
R685 B.n709 B.n708 585
R686 B.n707 B.n706 585
R687 B.n705 B.n704 585
R688 B.n703 B.n702 585
R689 B.n701 B.n700 585
R690 B.n699 B.n698 585
R691 B.n697 B.n696 585
R692 B.n695 B.n694 585
R693 B.n693 B.n692 585
R694 B.n691 B.n690 585
R695 B.n689 B.n688 585
R696 B.n687 B.n686 585
R697 B.n685 B.n684 585
R698 B.n683 B.n682 585
R699 B.n681 B.n680 585
R700 B.n679 B.n678 585
R701 B.n677 B.n676 585
R702 B.n675 B.n674 585
R703 B.n673 B.n672 585
R704 B.n671 B.n670 585
R705 B.n669 B.n668 585
R706 B.n667 B.n666 585
R707 B.n665 B.n664 585
R708 B.n663 B.n662 585
R709 B.n661 B.n660 585
R710 B.n659 B.n658 585
R711 B.n657 B.n656 585
R712 B.n655 B.n654 585
R713 B.n653 B.n652 585
R714 B.n651 B.n650 585
R715 B.n649 B.n648 585
R716 B.n647 B.n646 585
R717 B.n645 B.n644 585
R718 B.n643 B.n642 585
R719 B.n641 B.n640 585
R720 B.n639 B.n638 585
R721 B.n637 B.n636 585
R722 B.n906 B.n561 585
R723 B.n561 B.n560 585
R724 B.n908 B.n907 585
R725 B.n909 B.n908 585
R726 B.n555 B.n554 585
R727 B.n556 B.n555 585
R728 B.n917 B.n916 585
R729 B.n916 B.n915 585
R730 B.n918 B.n553 585
R731 B.n553 B.n552 585
R732 B.n920 B.n919 585
R733 B.n921 B.n920 585
R734 B.n547 B.n546 585
R735 B.n548 B.n547 585
R736 B.n929 B.n928 585
R737 B.n928 B.n927 585
R738 B.n930 B.n545 585
R739 B.n545 B.n544 585
R740 B.n932 B.n931 585
R741 B.n933 B.n932 585
R742 B.n539 B.n538 585
R743 B.n540 B.n539 585
R744 B.n941 B.n940 585
R745 B.n940 B.n939 585
R746 B.n942 B.n537 585
R747 B.n537 B.n536 585
R748 B.n944 B.n943 585
R749 B.n945 B.n944 585
R750 B.n531 B.n530 585
R751 B.n532 B.n531 585
R752 B.n953 B.n952 585
R753 B.n952 B.n951 585
R754 B.n954 B.n529 585
R755 B.n529 B.n528 585
R756 B.n956 B.n955 585
R757 B.n957 B.n956 585
R758 B.n523 B.n522 585
R759 B.n524 B.n523 585
R760 B.n965 B.n964 585
R761 B.n964 B.n963 585
R762 B.n966 B.n521 585
R763 B.n521 B.n520 585
R764 B.n968 B.n967 585
R765 B.n969 B.n968 585
R766 B.n515 B.n514 585
R767 B.n516 B.n515 585
R768 B.n977 B.n976 585
R769 B.n976 B.n975 585
R770 B.n978 B.n513 585
R771 B.n513 B.n512 585
R772 B.n980 B.n979 585
R773 B.n981 B.n980 585
R774 B.n507 B.n506 585
R775 B.n508 B.n507 585
R776 B.n990 B.n989 585
R777 B.n989 B.n988 585
R778 B.n991 B.n505 585
R779 B.n987 B.n505 585
R780 B.n993 B.n992 585
R781 B.n994 B.n993 585
R782 B.n500 B.n499 585
R783 B.n501 B.n500 585
R784 B.n1002 B.n1001 585
R785 B.n1001 B.n1000 585
R786 B.n1003 B.n498 585
R787 B.n498 B.n497 585
R788 B.n1005 B.n1004 585
R789 B.n1006 B.n1005 585
R790 B.n492 B.n491 585
R791 B.n493 B.n492 585
R792 B.n1015 B.n1014 585
R793 B.n1014 B.n1013 585
R794 B.n1016 B.n490 585
R795 B.n1012 B.n490 585
R796 B.n1018 B.n1017 585
R797 B.n1019 B.n1018 585
R798 B.n485 B.n484 585
R799 B.n486 B.n485 585
R800 B.n1027 B.n1026 585
R801 B.n1026 B.n1025 585
R802 B.n1028 B.n483 585
R803 B.n483 B.n482 585
R804 B.n1030 B.n1029 585
R805 B.n1031 B.n1030 585
R806 B.n477 B.n476 585
R807 B.n478 B.n477 585
R808 B.n1039 B.n1038 585
R809 B.n1038 B.n1037 585
R810 B.n1040 B.n475 585
R811 B.n475 B.n474 585
R812 B.n1042 B.n1041 585
R813 B.n1043 B.n1042 585
R814 B.n469 B.n468 585
R815 B.n470 B.n469 585
R816 B.n1051 B.n1050 585
R817 B.n1050 B.n1049 585
R818 B.n1052 B.n467 585
R819 B.n467 B.n466 585
R820 B.n1054 B.n1053 585
R821 B.n1055 B.n1054 585
R822 B.n461 B.n460 585
R823 B.n462 B.n461 585
R824 B.n1063 B.n1062 585
R825 B.n1062 B.n1061 585
R826 B.n1064 B.n459 585
R827 B.n459 B.n458 585
R828 B.n1066 B.n1065 585
R829 B.n1067 B.n1066 585
R830 B.n453 B.n452 585
R831 B.n454 B.n453 585
R832 B.n1076 B.n1075 585
R833 B.n1075 B.n1074 585
R834 B.n1077 B.n451 585
R835 B.n451 B.n450 585
R836 B.n1079 B.n1078 585
R837 B.n1080 B.n1079 585
R838 B.n3 B.n0 585
R839 B.n4 B.n3 585
R840 B.n1281 B.n1 585
R841 B.n1282 B.n1281 585
R842 B.n1280 B.n1279 585
R843 B.n1280 B.n8 585
R844 B.n1278 B.n9 585
R845 B.n12 B.n9 585
R846 B.n1277 B.n1276 585
R847 B.n1276 B.n1275 585
R848 B.n11 B.n10 585
R849 B.n1274 B.n11 585
R850 B.n1272 B.n1271 585
R851 B.n1273 B.n1272 585
R852 B.n1270 B.n17 585
R853 B.n17 B.n16 585
R854 B.n1269 B.n1268 585
R855 B.n1268 B.n1267 585
R856 B.n19 B.n18 585
R857 B.n1266 B.n19 585
R858 B.n1264 B.n1263 585
R859 B.n1265 B.n1264 585
R860 B.n1262 B.n24 585
R861 B.n24 B.n23 585
R862 B.n1261 B.n1260 585
R863 B.n1260 B.n1259 585
R864 B.n26 B.n25 585
R865 B.n1258 B.n26 585
R866 B.n1256 B.n1255 585
R867 B.n1257 B.n1256 585
R868 B.n1254 B.n31 585
R869 B.n31 B.n30 585
R870 B.n1253 B.n1252 585
R871 B.n1252 B.n1251 585
R872 B.n33 B.n32 585
R873 B.n1250 B.n33 585
R874 B.n1248 B.n1247 585
R875 B.n1249 B.n1248 585
R876 B.n1246 B.n38 585
R877 B.n38 B.n37 585
R878 B.n1245 B.n1244 585
R879 B.n1244 B.n1243 585
R880 B.n40 B.n39 585
R881 B.n1242 B.n40 585
R882 B.n1240 B.n1239 585
R883 B.n1241 B.n1240 585
R884 B.n1238 B.n44 585
R885 B.n47 B.n44 585
R886 B.n1237 B.n1236 585
R887 B.n1236 B.n1235 585
R888 B.n46 B.n45 585
R889 B.n1234 B.n46 585
R890 B.n1232 B.n1231 585
R891 B.n1233 B.n1232 585
R892 B.n1230 B.n52 585
R893 B.n52 B.n51 585
R894 B.n1229 B.n1228 585
R895 B.n1228 B.n1227 585
R896 B.n54 B.n53 585
R897 B.n1226 B.n54 585
R898 B.n1224 B.n1223 585
R899 B.n1225 B.n1224 585
R900 B.n1222 B.n58 585
R901 B.n61 B.n58 585
R902 B.n1221 B.n1220 585
R903 B.n1220 B.n1219 585
R904 B.n60 B.n59 585
R905 B.n1218 B.n60 585
R906 B.n1216 B.n1215 585
R907 B.n1217 B.n1216 585
R908 B.n1214 B.n66 585
R909 B.n66 B.n65 585
R910 B.n1213 B.n1212 585
R911 B.n1212 B.n1211 585
R912 B.n68 B.n67 585
R913 B.n1210 B.n68 585
R914 B.n1208 B.n1207 585
R915 B.n1209 B.n1208 585
R916 B.n1206 B.n73 585
R917 B.n73 B.n72 585
R918 B.n1205 B.n1204 585
R919 B.n1204 B.n1203 585
R920 B.n75 B.n74 585
R921 B.n1202 B.n75 585
R922 B.n1200 B.n1199 585
R923 B.n1201 B.n1200 585
R924 B.n1198 B.n80 585
R925 B.n80 B.n79 585
R926 B.n1197 B.n1196 585
R927 B.n1196 B.n1195 585
R928 B.n82 B.n81 585
R929 B.n1194 B.n82 585
R930 B.n1192 B.n1191 585
R931 B.n1193 B.n1192 585
R932 B.n1190 B.n87 585
R933 B.n87 B.n86 585
R934 B.n1189 B.n1188 585
R935 B.n1188 B.n1187 585
R936 B.n89 B.n88 585
R937 B.n1186 B.n89 585
R938 B.n1184 B.n1183 585
R939 B.n1185 B.n1184 585
R940 B.n1182 B.n94 585
R941 B.n94 B.n93 585
R942 B.n1181 B.n1180 585
R943 B.n1180 B.n1179 585
R944 B.n96 B.n95 585
R945 B.n1178 B.n96 585
R946 B.n1176 B.n1175 585
R947 B.n1177 B.n1176 585
R948 B.n1174 B.n101 585
R949 B.n101 B.n100 585
R950 B.n1173 B.n1172 585
R951 B.n1172 B.n1171 585
R952 B.n103 B.n102 585
R953 B.n1170 B.n103 585
R954 B.n1168 B.n1167 585
R955 B.n1169 B.n1168 585
R956 B.n1166 B.n108 585
R957 B.n108 B.n107 585
R958 B.n1285 B.n1284 585
R959 B.n1283 B.n2 585
R960 B.n1164 B.n108 502.111
R961 B.n1161 B.n178 502.111
R962 B.n636 B.n559 502.111
R963 B.n904 B.n561 502.111
R964 B.n182 B.t10 388.517
R965 B.n179 B.t18 388.517
R966 B.n634 B.t14 388.517
R967 B.n631 B.t21 388.517
R968 B.n1162 B.n176 256.663
R969 B.n1162 B.n175 256.663
R970 B.n1162 B.n174 256.663
R971 B.n1162 B.n173 256.663
R972 B.n1162 B.n172 256.663
R973 B.n1162 B.n171 256.663
R974 B.n1162 B.n170 256.663
R975 B.n1162 B.n169 256.663
R976 B.n1162 B.n168 256.663
R977 B.n1162 B.n167 256.663
R978 B.n1162 B.n166 256.663
R979 B.n1162 B.n165 256.663
R980 B.n1162 B.n164 256.663
R981 B.n1162 B.n163 256.663
R982 B.n1162 B.n162 256.663
R983 B.n1162 B.n161 256.663
R984 B.n1162 B.n160 256.663
R985 B.n1162 B.n159 256.663
R986 B.n1162 B.n158 256.663
R987 B.n1162 B.n157 256.663
R988 B.n1162 B.n156 256.663
R989 B.n1162 B.n155 256.663
R990 B.n1162 B.n154 256.663
R991 B.n1162 B.n153 256.663
R992 B.n1162 B.n152 256.663
R993 B.n1162 B.n151 256.663
R994 B.n1162 B.n150 256.663
R995 B.n1162 B.n149 256.663
R996 B.n1162 B.n148 256.663
R997 B.n1162 B.n147 256.663
R998 B.n1162 B.n146 256.663
R999 B.n1162 B.n145 256.663
R1000 B.n1162 B.n144 256.663
R1001 B.n1162 B.n143 256.663
R1002 B.n1162 B.n142 256.663
R1003 B.n1162 B.n141 256.663
R1004 B.n1162 B.n140 256.663
R1005 B.n1162 B.n139 256.663
R1006 B.n1162 B.n138 256.663
R1007 B.n1162 B.n137 256.663
R1008 B.n1162 B.n136 256.663
R1009 B.n1162 B.n135 256.663
R1010 B.n1162 B.n134 256.663
R1011 B.n1162 B.n133 256.663
R1012 B.n1162 B.n132 256.663
R1013 B.n1162 B.n131 256.663
R1014 B.n1162 B.n130 256.663
R1015 B.n1162 B.n129 256.663
R1016 B.n1162 B.n128 256.663
R1017 B.n1162 B.n127 256.663
R1018 B.n1162 B.n126 256.663
R1019 B.n1162 B.n125 256.663
R1020 B.n1162 B.n124 256.663
R1021 B.n1162 B.n123 256.663
R1022 B.n1162 B.n122 256.663
R1023 B.n1162 B.n121 256.663
R1024 B.n1162 B.n120 256.663
R1025 B.n1162 B.n119 256.663
R1026 B.n1162 B.n118 256.663
R1027 B.n1162 B.n117 256.663
R1028 B.n1162 B.n116 256.663
R1029 B.n1162 B.n115 256.663
R1030 B.n1162 B.n114 256.663
R1031 B.n1162 B.n113 256.663
R1032 B.n1162 B.n112 256.663
R1033 B.n1162 B.n111 256.663
R1034 B.n1163 B.n1162 256.663
R1035 B.n903 B.n902 256.663
R1036 B.n902 B.n564 256.663
R1037 B.n902 B.n565 256.663
R1038 B.n902 B.n566 256.663
R1039 B.n902 B.n567 256.663
R1040 B.n902 B.n568 256.663
R1041 B.n902 B.n569 256.663
R1042 B.n902 B.n570 256.663
R1043 B.n902 B.n571 256.663
R1044 B.n902 B.n572 256.663
R1045 B.n902 B.n573 256.663
R1046 B.n902 B.n574 256.663
R1047 B.n902 B.n575 256.663
R1048 B.n902 B.n576 256.663
R1049 B.n902 B.n577 256.663
R1050 B.n902 B.n578 256.663
R1051 B.n902 B.n579 256.663
R1052 B.n902 B.n580 256.663
R1053 B.n902 B.n581 256.663
R1054 B.n902 B.n582 256.663
R1055 B.n902 B.n583 256.663
R1056 B.n902 B.n584 256.663
R1057 B.n902 B.n585 256.663
R1058 B.n902 B.n586 256.663
R1059 B.n902 B.n587 256.663
R1060 B.n902 B.n588 256.663
R1061 B.n902 B.n589 256.663
R1062 B.n902 B.n590 256.663
R1063 B.n902 B.n591 256.663
R1064 B.n902 B.n592 256.663
R1065 B.n902 B.n593 256.663
R1066 B.n902 B.n594 256.663
R1067 B.n902 B.n595 256.663
R1068 B.n902 B.n596 256.663
R1069 B.n902 B.n597 256.663
R1070 B.n902 B.n598 256.663
R1071 B.n902 B.n599 256.663
R1072 B.n902 B.n600 256.663
R1073 B.n902 B.n601 256.663
R1074 B.n902 B.n602 256.663
R1075 B.n902 B.n603 256.663
R1076 B.n902 B.n604 256.663
R1077 B.n902 B.n605 256.663
R1078 B.n902 B.n606 256.663
R1079 B.n902 B.n607 256.663
R1080 B.n902 B.n608 256.663
R1081 B.n902 B.n609 256.663
R1082 B.n902 B.n610 256.663
R1083 B.n902 B.n611 256.663
R1084 B.n902 B.n612 256.663
R1085 B.n902 B.n613 256.663
R1086 B.n902 B.n614 256.663
R1087 B.n902 B.n615 256.663
R1088 B.n902 B.n616 256.663
R1089 B.n902 B.n617 256.663
R1090 B.n902 B.n618 256.663
R1091 B.n902 B.n619 256.663
R1092 B.n902 B.n620 256.663
R1093 B.n902 B.n621 256.663
R1094 B.n902 B.n622 256.663
R1095 B.n902 B.n623 256.663
R1096 B.n902 B.n624 256.663
R1097 B.n902 B.n625 256.663
R1098 B.n902 B.n626 256.663
R1099 B.n902 B.n627 256.663
R1100 B.n902 B.n628 256.663
R1101 B.n902 B.n629 256.663
R1102 B.n1287 B.n1286 256.663
R1103 B.n184 B.n110 163.367
R1104 B.n188 B.n187 163.367
R1105 B.n192 B.n191 163.367
R1106 B.n196 B.n195 163.367
R1107 B.n200 B.n199 163.367
R1108 B.n204 B.n203 163.367
R1109 B.n208 B.n207 163.367
R1110 B.n212 B.n211 163.367
R1111 B.n216 B.n215 163.367
R1112 B.n220 B.n219 163.367
R1113 B.n224 B.n223 163.367
R1114 B.n228 B.n227 163.367
R1115 B.n232 B.n231 163.367
R1116 B.n236 B.n235 163.367
R1117 B.n240 B.n239 163.367
R1118 B.n244 B.n243 163.367
R1119 B.n248 B.n247 163.367
R1120 B.n252 B.n251 163.367
R1121 B.n256 B.n255 163.367
R1122 B.n260 B.n259 163.367
R1123 B.n264 B.n263 163.367
R1124 B.n268 B.n267 163.367
R1125 B.n272 B.n271 163.367
R1126 B.n276 B.n275 163.367
R1127 B.n280 B.n279 163.367
R1128 B.n284 B.n283 163.367
R1129 B.n288 B.n287 163.367
R1130 B.n292 B.n291 163.367
R1131 B.n296 B.n295 163.367
R1132 B.n300 B.n299 163.367
R1133 B.n304 B.n303 163.367
R1134 B.n309 B.n308 163.367
R1135 B.n313 B.n312 163.367
R1136 B.n317 B.n316 163.367
R1137 B.n321 B.n320 163.367
R1138 B.n325 B.n324 163.367
R1139 B.n329 B.n328 163.367
R1140 B.n333 B.n332 163.367
R1141 B.n337 B.n336 163.367
R1142 B.n341 B.n340 163.367
R1143 B.n345 B.n344 163.367
R1144 B.n349 B.n348 163.367
R1145 B.n353 B.n352 163.367
R1146 B.n357 B.n356 163.367
R1147 B.n361 B.n360 163.367
R1148 B.n365 B.n364 163.367
R1149 B.n369 B.n368 163.367
R1150 B.n373 B.n372 163.367
R1151 B.n377 B.n376 163.367
R1152 B.n381 B.n380 163.367
R1153 B.n385 B.n384 163.367
R1154 B.n389 B.n388 163.367
R1155 B.n393 B.n392 163.367
R1156 B.n397 B.n396 163.367
R1157 B.n401 B.n400 163.367
R1158 B.n405 B.n404 163.367
R1159 B.n409 B.n408 163.367
R1160 B.n413 B.n412 163.367
R1161 B.n417 B.n416 163.367
R1162 B.n421 B.n420 163.367
R1163 B.n425 B.n424 163.367
R1164 B.n429 B.n428 163.367
R1165 B.n433 B.n432 163.367
R1166 B.n437 B.n436 163.367
R1167 B.n441 B.n440 163.367
R1168 B.n445 B.n444 163.367
R1169 B.n1161 B.n177 163.367
R1170 B.n910 B.n559 163.367
R1171 B.n910 B.n557 163.367
R1172 B.n914 B.n557 163.367
R1173 B.n914 B.n551 163.367
R1174 B.n922 B.n551 163.367
R1175 B.n922 B.n549 163.367
R1176 B.n926 B.n549 163.367
R1177 B.n926 B.n543 163.367
R1178 B.n934 B.n543 163.367
R1179 B.n934 B.n541 163.367
R1180 B.n938 B.n541 163.367
R1181 B.n938 B.n535 163.367
R1182 B.n946 B.n535 163.367
R1183 B.n946 B.n533 163.367
R1184 B.n950 B.n533 163.367
R1185 B.n950 B.n527 163.367
R1186 B.n958 B.n527 163.367
R1187 B.n958 B.n525 163.367
R1188 B.n962 B.n525 163.367
R1189 B.n962 B.n519 163.367
R1190 B.n970 B.n519 163.367
R1191 B.n970 B.n517 163.367
R1192 B.n974 B.n517 163.367
R1193 B.n974 B.n511 163.367
R1194 B.n982 B.n511 163.367
R1195 B.n982 B.n509 163.367
R1196 B.n986 B.n509 163.367
R1197 B.n986 B.n504 163.367
R1198 B.n995 B.n504 163.367
R1199 B.n995 B.n502 163.367
R1200 B.n999 B.n502 163.367
R1201 B.n999 B.n496 163.367
R1202 B.n1007 B.n496 163.367
R1203 B.n1007 B.n494 163.367
R1204 B.n1011 B.n494 163.367
R1205 B.n1011 B.n489 163.367
R1206 B.n1020 B.n489 163.367
R1207 B.n1020 B.n487 163.367
R1208 B.n1024 B.n487 163.367
R1209 B.n1024 B.n481 163.367
R1210 B.n1032 B.n481 163.367
R1211 B.n1032 B.n479 163.367
R1212 B.n1036 B.n479 163.367
R1213 B.n1036 B.n473 163.367
R1214 B.n1044 B.n473 163.367
R1215 B.n1044 B.n471 163.367
R1216 B.n1048 B.n471 163.367
R1217 B.n1048 B.n465 163.367
R1218 B.n1056 B.n465 163.367
R1219 B.n1056 B.n463 163.367
R1220 B.n1060 B.n463 163.367
R1221 B.n1060 B.n457 163.367
R1222 B.n1068 B.n457 163.367
R1223 B.n1068 B.n455 163.367
R1224 B.n1073 B.n455 163.367
R1225 B.n1073 B.n449 163.367
R1226 B.n1081 B.n449 163.367
R1227 B.n1082 B.n1081 163.367
R1228 B.n1082 B.n5 163.367
R1229 B.n6 B.n5 163.367
R1230 B.n7 B.n6 163.367
R1231 B.n1088 B.n7 163.367
R1232 B.n1089 B.n1088 163.367
R1233 B.n1089 B.n13 163.367
R1234 B.n14 B.n13 163.367
R1235 B.n15 B.n14 163.367
R1236 B.n1094 B.n15 163.367
R1237 B.n1094 B.n20 163.367
R1238 B.n21 B.n20 163.367
R1239 B.n22 B.n21 163.367
R1240 B.n1099 B.n22 163.367
R1241 B.n1099 B.n27 163.367
R1242 B.n28 B.n27 163.367
R1243 B.n29 B.n28 163.367
R1244 B.n1104 B.n29 163.367
R1245 B.n1104 B.n34 163.367
R1246 B.n35 B.n34 163.367
R1247 B.n36 B.n35 163.367
R1248 B.n1109 B.n36 163.367
R1249 B.n1109 B.n41 163.367
R1250 B.n42 B.n41 163.367
R1251 B.n43 B.n42 163.367
R1252 B.n1114 B.n43 163.367
R1253 B.n1114 B.n48 163.367
R1254 B.n49 B.n48 163.367
R1255 B.n50 B.n49 163.367
R1256 B.n1119 B.n50 163.367
R1257 B.n1119 B.n55 163.367
R1258 B.n56 B.n55 163.367
R1259 B.n57 B.n56 163.367
R1260 B.n1124 B.n57 163.367
R1261 B.n1124 B.n62 163.367
R1262 B.n63 B.n62 163.367
R1263 B.n64 B.n63 163.367
R1264 B.n1129 B.n64 163.367
R1265 B.n1129 B.n69 163.367
R1266 B.n70 B.n69 163.367
R1267 B.n71 B.n70 163.367
R1268 B.n1134 B.n71 163.367
R1269 B.n1134 B.n76 163.367
R1270 B.n77 B.n76 163.367
R1271 B.n78 B.n77 163.367
R1272 B.n1139 B.n78 163.367
R1273 B.n1139 B.n83 163.367
R1274 B.n84 B.n83 163.367
R1275 B.n85 B.n84 163.367
R1276 B.n1144 B.n85 163.367
R1277 B.n1144 B.n90 163.367
R1278 B.n91 B.n90 163.367
R1279 B.n92 B.n91 163.367
R1280 B.n1149 B.n92 163.367
R1281 B.n1149 B.n97 163.367
R1282 B.n98 B.n97 163.367
R1283 B.n99 B.n98 163.367
R1284 B.n1154 B.n99 163.367
R1285 B.n1154 B.n104 163.367
R1286 B.n105 B.n104 163.367
R1287 B.n106 B.n105 163.367
R1288 B.n178 B.n106 163.367
R1289 B.n901 B.n563 163.367
R1290 B.n901 B.n630 163.367
R1291 B.n897 B.n896 163.367
R1292 B.n893 B.n892 163.367
R1293 B.n889 B.n888 163.367
R1294 B.n885 B.n884 163.367
R1295 B.n881 B.n880 163.367
R1296 B.n877 B.n876 163.367
R1297 B.n873 B.n872 163.367
R1298 B.n869 B.n868 163.367
R1299 B.n865 B.n864 163.367
R1300 B.n861 B.n860 163.367
R1301 B.n857 B.n856 163.367
R1302 B.n853 B.n852 163.367
R1303 B.n849 B.n848 163.367
R1304 B.n845 B.n844 163.367
R1305 B.n841 B.n840 163.367
R1306 B.n837 B.n836 163.367
R1307 B.n833 B.n832 163.367
R1308 B.n829 B.n828 163.367
R1309 B.n825 B.n824 163.367
R1310 B.n821 B.n820 163.367
R1311 B.n817 B.n816 163.367
R1312 B.n813 B.n812 163.367
R1313 B.n809 B.n808 163.367
R1314 B.n805 B.n804 163.367
R1315 B.n801 B.n800 163.367
R1316 B.n797 B.n796 163.367
R1317 B.n793 B.n792 163.367
R1318 B.n789 B.n788 163.367
R1319 B.n785 B.n784 163.367
R1320 B.n781 B.n780 163.367
R1321 B.n777 B.n776 163.367
R1322 B.n773 B.n772 163.367
R1323 B.n769 B.n768 163.367
R1324 B.n765 B.n764 163.367
R1325 B.n760 B.n759 163.367
R1326 B.n756 B.n755 163.367
R1327 B.n752 B.n751 163.367
R1328 B.n748 B.n747 163.367
R1329 B.n744 B.n743 163.367
R1330 B.n740 B.n739 163.367
R1331 B.n736 B.n735 163.367
R1332 B.n732 B.n731 163.367
R1333 B.n728 B.n727 163.367
R1334 B.n724 B.n723 163.367
R1335 B.n720 B.n719 163.367
R1336 B.n716 B.n715 163.367
R1337 B.n712 B.n711 163.367
R1338 B.n708 B.n707 163.367
R1339 B.n704 B.n703 163.367
R1340 B.n700 B.n699 163.367
R1341 B.n696 B.n695 163.367
R1342 B.n692 B.n691 163.367
R1343 B.n688 B.n687 163.367
R1344 B.n684 B.n683 163.367
R1345 B.n680 B.n679 163.367
R1346 B.n676 B.n675 163.367
R1347 B.n672 B.n671 163.367
R1348 B.n668 B.n667 163.367
R1349 B.n664 B.n663 163.367
R1350 B.n660 B.n659 163.367
R1351 B.n656 B.n655 163.367
R1352 B.n652 B.n651 163.367
R1353 B.n648 B.n647 163.367
R1354 B.n644 B.n643 163.367
R1355 B.n640 B.n639 163.367
R1356 B.n908 B.n561 163.367
R1357 B.n908 B.n555 163.367
R1358 B.n916 B.n555 163.367
R1359 B.n916 B.n553 163.367
R1360 B.n920 B.n553 163.367
R1361 B.n920 B.n547 163.367
R1362 B.n928 B.n547 163.367
R1363 B.n928 B.n545 163.367
R1364 B.n932 B.n545 163.367
R1365 B.n932 B.n539 163.367
R1366 B.n940 B.n539 163.367
R1367 B.n940 B.n537 163.367
R1368 B.n944 B.n537 163.367
R1369 B.n944 B.n531 163.367
R1370 B.n952 B.n531 163.367
R1371 B.n952 B.n529 163.367
R1372 B.n956 B.n529 163.367
R1373 B.n956 B.n523 163.367
R1374 B.n964 B.n523 163.367
R1375 B.n964 B.n521 163.367
R1376 B.n968 B.n521 163.367
R1377 B.n968 B.n515 163.367
R1378 B.n976 B.n515 163.367
R1379 B.n976 B.n513 163.367
R1380 B.n980 B.n513 163.367
R1381 B.n980 B.n507 163.367
R1382 B.n989 B.n507 163.367
R1383 B.n989 B.n505 163.367
R1384 B.n993 B.n505 163.367
R1385 B.n993 B.n500 163.367
R1386 B.n1001 B.n500 163.367
R1387 B.n1001 B.n498 163.367
R1388 B.n1005 B.n498 163.367
R1389 B.n1005 B.n492 163.367
R1390 B.n1014 B.n492 163.367
R1391 B.n1014 B.n490 163.367
R1392 B.n1018 B.n490 163.367
R1393 B.n1018 B.n485 163.367
R1394 B.n1026 B.n485 163.367
R1395 B.n1026 B.n483 163.367
R1396 B.n1030 B.n483 163.367
R1397 B.n1030 B.n477 163.367
R1398 B.n1038 B.n477 163.367
R1399 B.n1038 B.n475 163.367
R1400 B.n1042 B.n475 163.367
R1401 B.n1042 B.n469 163.367
R1402 B.n1050 B.n469 163.367
R1403 B.n1050 B.n467 163.367
R1404 B.n1054 B.n467 163.367
R1405 B.n1054 B.n461 163.367
R1406 B.n1062 B.n461 163.367
R1407 B.n1062 B.n459 163.367
R1408 B.n1066 B.n459 163.367
R1409 B.n1066 B.n453 163.367
R1410 B.n1075 B.n453 163.367
R1411 B.n1075 B.n451 163.367
R1412 B.n1079 B.n451 163.367
R1413 B.n1079 B.n3 163.367
R1414 B.n1285 B.n3 163.367
R1415 B.n1281 B.n2 163.367
R1416 B.n1281 B.n1280 163.367
R1417 B.n1280 B.n9 163.367
R1418 B.n1276 B.n9 163.367
R1419 B.n1276 B.n11 163.367
R1420 B.n1272 B.n11 163.367
R1421 B.n1272 B.n17 163.367
R1422 B.n1268 B.n17 163.367
R1423 B.n1268 B.n19 163.367
R1424 B.n1264 B.n19 163.367
R1425 B.n1264 B.n24 163.367
R1426 B.n1260 B.n24 163.367
R1427 B.n1260 B.n26 163.367
R1428 B.n1256 B.n26 163.367
R1429 B.n1256 B.n31 163.367
R1430 B.n1252 B.n31 163.367
R1431 B.n1252 B.n33 163.367
R1432 B.n1248 B.n33 163.367
R1433 B.n1248 B.n38 163.367
R1434 B.n1244 B.n38 163.367
R1435 B.n1244 B.n40 163.367
R1436 B.n1240 B.n40 163.367
R1437 B.n1240 B.n44 163.367
R1438 B.n1236 B.n44 163.367
R1439 B.n1236 B.n46 163.367
R1440 B.n1232 B.n46 163.367
R1441 B.n1232 B.n52 163.367
R1442 B.n1228 B.n52 163.367
R1443 B.n1228 B.n54 163.367
R1444 B.n1224 B.n54 163.367
R1445 B.n1224 B.n58 163.367
R1446 B.n1220 B.n58 163.367
R1447 B.n1220 B.n60 163.367
R1448 B.n1216 B.n60 163.367
R1449 B.n1216 B.n66 163.367
R1450 B.n1212 B.n66 163.367
R1451 B.n1212 B.n68 163.367
R1452 B.n1208 B.n68 163.367
R1453 B.n1208 B.n73 163.367
R1454 B.n1204 B.n73 163.367
R1455 B.n1204 B.n75 163.367
R1456 B.n1200 B.n75 163.367
R1457 B.n1200 B.n80 163.367
R1458 B.n1196 B.n80 163.367
R1459 B.n1196 B.n82 163.367
R1460 B.n1192 B.n82 163.367
R1461 B.n1192 B.n87 163.367
R1462 B.n1188 B.n87 163.367
R1463 B.n1188 B.n89 163.367
R1464 B.n1184 B.n89 163.367
R1465 B.n1184 B.n94 163.367
R1466 B.n1180 B.n94 163.367
R1467 B.n1180 B.n96 163.367
R1468 B.n1176 B.n96 163.367
R1469 B.n1176 B.n101 163.367
R1470 B.n1172 B.n101 163.367
R1471 B.n1172 B.n103 163.367
R1472 B.n1168 B.n103 163.367
R1473 B.n1168 B.n108 163.367
R1474 B.n179 B.t19 127.495
R1475 B.n634 B.t17 127.495
R1476 B.n182 B.t12 127.469
R1477 B.n631 B.t23 127.469
R1478 B.n1164 B.n1163 71.676
R1479 B.n184 B.n111 71.676
R1480 B.n188 B.n112 71.676
R1481 B.n192 B.n113 71.676
R1482 B.n196 B.n114 71.676
R1483 B.n200 B.n115 71.676
R1484 B.n204 B.n116 71.676
R1485 B.n208 B.n117 71.676
R1486 B.n212 B.n118 71.676
R1487 B.n216 B.n119 71.676
R1488 B.n220 B.n120 71.676
R1489 B.n224 B.n121 71.676
R1490 B.n228 B.n122 71.676
R1491 B.n232 B.n123 71.676
R1492 B.n236 B.n124 71.676
R1493 B.n240 B.n125 71.676
R1494 B.n244 B.n126 71.676
R1495 B.n248 B.n127 71.676
R1496 B.n252 B.n128 71.676
R1497 B.n256 B.n129 71.676
R1498 B.n260 B.n130 71.676
R1499 B.n264 B.n131 71.676
R1500 B.n268 B.n132 71.676
R1501 B.n272 B.n133 71.676
R1502 B.n276 B.n134 71.676
R1503 B.n280 B.n135 71.676
R1504 B.n284 B.n136 71.676
R1505 B.n288 B.n137 71.676
R1506 B.n292 B.n138 71.676
R1507 B.n296 B.n139 71.676
R1508 B.n300 B.n140 71.676
R1509 B.n304 B.n141 71.676
R1510 B.n309 B.n142 71.676
R1511 B.n313 B.n143 71.676
R1512 B.n317 B.n144 71.676
R1513 B.n321 B.n145 71.676
R1514 B.n325 B.n146 71.676
R1515 B.n329 B.n147 71.676
R1516 B.n333 B.n148 71.676
R1517 B.n337 B.n149 71.676
R1518 B.n341 B.n150 71.676
R1519 B.n345 B.n151 71.676
R1520 B.n349 B.n152 71.676
R1521 B.n353 B.n153 71.676
R1522 B.n357 B.n154 71.676
R1523 B.n361 B.n155 71.676
R1524 B.n365 B.n156 71.676
R1525 B.n369 B.n157 71.676
R1526 B.n373 B.n158 71.676
R1527 B.n377 B.n159 71.676
R1528 B.n381 B.n160 71.676
R1529 B.n385 B.n161 71.676
R1530 B.n389 B.n162 71.676
R1531 B.n393 B.n163 71.676
R1532 B.n397 B.n164 71.676
R1533 B.n401 B.n165 71.676
R1534 B.n405 B.n166 71.676
R1535 B.n409 B.n167 71.676
R1536 B.n413 B.n168 71.676
R1537 B.n417 B.n169 71.676
R1538 B.n421 B.n170 71.676
R1539 B.n425 B.n171 71.676
R1540 B.n429 B.n172 71.676
R1541 B.n433 B.n173 71.676
R1542 B.n437 B.n174 71.676
R1543 B.n441 B.n175 71.676
R1544 B.n445 B.n176 71.676
R1545 B.n177 B.n176 71.676
R1546 B.n444 B.n175 71.676
R1547 B.n440 B.n174 71.676
R1548 B.n436 B.n173 71.676
R1549 B.n432 B.n172 71.676
R1550 B.n428 B.n171 71.676
R1551 B.n424 B.n170 71.676
R1552 B.n420 B.n169 71.676
R1553 B.n416 B.n168 71.676
R1554 B.n412 B.n167 71.676
R1555 B.n408 B.n166 71.676
R1556 B.n404 B.n165 71.676
R1557 B.n400 B.n164 71.676
R1558 B.n396 B.n163 71.676
R1559 B.n392 B.n162 71.676
R1560 B.n388 B.n161 71.676
R1561 B.n384 B.n160 71.676
R1562 B.n380 B.n159 71.676
R1563 B.n376 B.n158 71.676
R1564 B.n372 B.n157 71.676
R1565 B.n368 B.n156 71.676
R1566 B.n364 B.n155 71.676
R1567 B.n360 B.n154 71.676
R1568 B.n356 B.n153 71.676
R1569 B.n352 B.n152 71.676
R1570 B.n348 B.n151 71.676
R1571 B.n344 B.n150 71.676
R1572 B.n340 B.n149 71.676
R1573 B.n336 B.n148 71.676
R1574 B.n332 B.n147 71.676
R1575 B.n328 B.n146 71.676
R1576 B.n324 B.n145 71.676
R1577 B.n320 B.n144 71.676
R1578 B.n316 B.n143 71.676
R1579 B.n312 B.n142 71.676
R1580 B.n308 B.n141 71.676
R1581 B.n303 B.n140 71.676
R1582 B.n299 B.n139 71.676
R1583 B.n295 B.n138 71.676
R1584 B.n291 B.n137 71.676
R1585 B.n287 B.n136 71.676
R1586 B.n283 B.n135 71.676
R1587 B.n279 B.n134 71.676
R1588 B.n275 B.n133 71.676
R1589 B.n271 B.n132 71.676
R1590 B.n267 B.n131 71.676
R1591 B.n263 B.n130 71.676
R1592 B.n259 B.n129 71.676
R1593 B.n255 B.n128 71.676
R1594 B.n251 B.n127 71.676
R1595 B.n247 B.n126 71.676
R1596 B.n243 B.n125 71.676
R1597 B.n239 B.n124 71.676
R1598 B.n235 B.n123 71.676
R1599 B.n231 B.n122 71.676
R1600 B.n227 B.n121 71.676
R1601 B.n223 B.n120 71.676
R1602 B.n219 B.n119 71.676
R1603 B.n215 B.n118 71.676
R1604 B.n211 B.n117 71.676
R1605 B.n207 B.n116 71.676
R1606 B.n203 B.n115 71.676
R1607 B.n199 B.n114 71.676
R1608 B.n195 B.n113 71.676
R1609 B.n191 B.n112 71.676
R1610 B.n187 B.n111 71.676
R1611 B.n1163 B.n110 71.676
R1612 B.n904 B.n903 71.676
R1613 B.n630 B.n564 71.676
R1614 B.n896 B.n565 71.676
R1615 B.n892 B.n566 71.676
R1616 B.n888 B.n567 71.676
R1617 B.n884 B.n568 71.676
R1618 B.n880 B.n569 71.676
R1619 B.n876 B.n570 71.676
R1620 B.n872 B.n571 71.676
R1621 B.n868 B.n572 71.676
R1622 B.n864 B.n573 71.676
R1623 B.n860 B.n574 71.676
R1624 B.n856 B.n575 71.676
R1625 B.n852 B.n576 71.676
R1626 B.n848 B.n577 71.676
R1627 B.n844 B.n578 71.676
R1628 B.n840 B.n579 71.676
R1629 B.n836 B.n580 71.676
R1630 B.n832 B.n581 71.676
R1631 B.n828 B.n582 71.676
R1632 B.n824 B.n583 71.676
R1633 B.n820 B.n584 71.676
R1634 B.n816 B.n585 71.676
R1635 B.n812 B.n586 71.676
R1636 B.n808 B.n587 71.676
R1637 B.n804 B.n588 71.676
R1638 B.n800 B.n589 71.676
R1639 B.n796 B.n590 71.676
R1640 B.n792 B.n591 71.676
R1641 B.n788 B.n592 71.676
R1642 B.n784 B.n593 71.676
R1643 B.n780 B.n594 71.676
R1644 B.n776 B.n595 71.676
R1645 B.n772 B.n596 71.676
R1646 B.n768 B.n597 71.676
R1647 B.n764 B.n598 71.676
R1648 B.n759 B.n599 71.676
R1649 B.n755 B.n600 71.676
R1650 B.n751 B.n601 71.676
R1651 B.n747 B.n602 71.676
R1652 B.n743 B.n603 71.676
R1653 B.n739 B.n604 71.676
R1654 B.n735 B.n605 71.676
R1655 B.n731 B.n606 71.676
R1656 B.n727 B.n607 71.676
R1657 B.n723 B.n608 71.676
R1658 B.n719 B.n609 71.676
R1659 B.n715 B.n610 71.676
R1660 B.n711 B.n611 71.676
R1661 B.n707 B.n612 71.676
R1662 B.n703 B.n613 71.676
R1663 B.n699 B.n614 71.676
R1664 B.n695 B.n615 71.676
R1665 B.n691 B.n616 71.676
R1666 B.n687 B.n617 71.676
R1667 B.n683 B.n618 71.676
R1668 B.n679 B.n619 71.676
R1669 B.n675 B.n620 71.676
R1670 B.n671 B.n621 71.676
R1671 B.n667 B.n622 71.676
R1672 B.n663 B.n623 71.676
R1673 B.n659 B.n624 71.676
R1674 B.n655 B.n625 71.676
R1675 B.n651 B.n626 71.676
R1676 B.n647 B.n627 71.676
R1677 B.n643 B.n628 71.676
R1678 B.n639 B.n629 71.676
R1679 B.n903 B.n563 71.676
R1680 B.n897 B.n564 71.676
R1681 B.n893 B.n565 71.676
R1682 B.n889 B.n566 71.676
R1683 B.n885 B.n567 71.676
R1684 B.n881 B.n568 71.676
R1685 B.n877 B.n569 71.676
R1686 B.n873 B.n570 71.676
R1687 B.n869 B.n571 71.676
R1688 B.n865 B.n572 71.676
R1689 B.n861 B.n573 71.676
R1690 B.n857 B.n574 71.676
R1691 B.n853 B.n575 71.676
R1692 B.n849 B.n576 71.676
R1693 B.n845 B.n577 71.676
R1694 B.n841 B.n578 71.676
R1695 B.n837 B.n579 71.676
R1696 B.n833 B.n580 71.676
R1697 B.n829 B.n581 71.676
R1698 B.n825 B.n582 71.676
R1699 B.n821 B.n583 71.676
R1700 B.n817 B.n584 71.676
R1701 B.n813 B.n585 71.676
R1702 B.n809 B.n586 71.676
R1703 B.n805 B.n587 71.676
R1704 B.n801 B.n588 71.676
R1705 B.n797 B.n589 71.676
R1706 B.n793 B.n590 71.676
R1707 B.n789 B.n591 71.676
R1708 B.n785 B.n592 71.676
R1709 B.n781 B.n593 71.676
R1710 B.n777 B.n594 71.676
R1711 B.n773 B.n595 71.676
R1712 B.n769 B.n596 71.676
R1713 B.n765 B.n597 71.676
R1714 B.n760 B.n598 71.676
R1715 B.n756 B.n599 71.676
R1716 B.n752 B.n600 71.676
R1717 B.n748 B.n601 71.676
R1718 B.n744 B.n602 71.676
R1719 B.n740 B.n603 71.676
R1720 B.n736 B.n604 71.676
R1721 B.n732 B.n605 71.676
R1722 B.n728 B.n606 71.676
R1723 B.n724 B.n607 71.676
R1724 B.n720 B.n608 71.676
R1725 B.n716 B.n609 71.676
R1726 B.n712 B.n610 71.676
R1727 B.n708 B.n611 71.676
R1728 B.n704 B.n612 71.676
R1729 B.n700 B.n613 71.676
R1730 B.n696 B.n614 71.676
R1731 B.n692 B.n615 71.676
R1732 B.n688 B.n616 71.676
R1733 B.n684 B.n617 71.676
R1734 B.n680 B.n618 71.676
R1735 B.n676 B.n619 71.676
R1736 B.n672 B.n620 71.676
R1737 B.n668 B.n621 71.676
R1738 B.n664 B.n622 71.676
R1739 B.n660 B.n623 71.676
R1740 B.n656 B.n624 71.676
R1741 B.n652 B.n625 71.676
R1742 B.n648 B.n626 71.676
R1743 B.n644 B.n627 71.676
R1744 B.n640 B.n628 71.676
R1745 B.n636 B.n629 71.676
R1746 B.n1286 B.n1285 71.676
R1747 B.n1286 B.n2 71.676
R1748 B.n180 B.t20 71.2517
R1749 B.n635 B.t16 71.2517
R1750 B.n183 B.t13 71.226
R1751 B.n632 B.t22 71.226
R1752 B.n306 B.n183 59.5399
R1753 B.n181 B.n180 59.5399
R1754 B.n762 B.n635 59.5399
R1755 B.n633 B.n632 59.5399
R1756 B.n183 B.n182 56.2429
R1757 B.n180 B.n179 56.2429
R1758 B.n635 B.n634 56.2429
R1759 B.n632 B.n631 56.2429
R1760 B.n902 B.n560 48.8894
R1761 B.n1162 B.n107 48.8894
R1762 B.n906 B.n905 32.6249
R1763 B.n637 B.n558 32.6249
R1764 B.n1160 B.n1159 32.6249
R1765 B.n1166 B.n1165 32.6249
R1766 B.n909 B.n560 30.5
R1767 B.n909 B.n556 30.5
R1768 B.n915 B.n556 30.5
R1769 B.n915 B.n552 30.5
R1770 B.n921 B.n552 30.5
R1771 B.n921 B.n548 30.5
R1772 B.n927 B.n548 30.5
R1773 B.n933 B.n544 30.5
R1774 B.n933 B.n540 30.5
R1775 B.n939 B.n540 30.5
R1776 B.n939 B.n536 30.5
R1777 B.n945 B.n536 30.5
R1778 B.n945 B.n532 30.5
R1779 B.n951 B.n532 30.5
R1780 B.n951 B.n528 30.5
R1781 B.n957 B.n528 30.5
R1782 B.n957 B.n524 30.5
R1783 B.n963 B.n524 30.5
R1784 B.n969 B.n520 30.5
R1785 B.n969 B.n516 30.5
R1786 B.n975 B.n516 30.5
R1787 B.n975 B.n512 30.5
R1788 B.n981 B.n512 30.5
R1789 B.n981 B.n508 30.5
R1790 B.n988 B.n508 30.5
R1791 B.n988 B.n987 30.5
R1792 B.n994 B.n501 30.5
R1793 B.n1000 B.n501 30.5
R1794 B.n1000 B.n497 30.5
R1795 B.n1006 B.n497 30.5
R1796 B.n1006 B.n493 30.5
R1797 B.n1013 B.n493 30.5
R1798 B.n1013 B.n1012 30.5
R1799 B.n1019 B.n486 30.5
R1800 B.n1025 B.n486 30.5
R1801 B.n1025 B.n482 30.5
R1802 B.n1031 B.n482 30.5
R1803 B.n1031 B.n478 30.5
R1804 B.n1037 B.n478 30.5
R1805 B.n1037 B.n474 30.5
R1806 B.n1043 B.n474 30.5
R1807 B.n1049 B.n470 30.5
R1808 B.n1049 B.n466 30.5
R1809 B.n1055 B.n466 30.5
R1810 B.n1055 B.n462 30.5
R1811 B.n1061 B.n462 30.5
R1812 B.n1061 B.n458 30.5
R1813 B.n1067 B.n458 30.5
R1814 B.n1074 B.n454 30.5
R1815 B.n1074 B.n450 30.5
R1816 B.n1080 B.n450 30.5
R1817 B.n1080 B.n4 30.5
R1818 B.n1284 B.n4 30.5
R1819 B.n1284 B.n1283 30.5
R1820 B.n1283 B.n1282 30.5
R1821 B.n1282 B.n8 30.5
R1822 B.n12 B.n8 30.5
R1823 B.n1275 B.n12 30.5
R1824 B.n1275 B.n1274 30.5
R1825 B.n1273 B.n16 30.5
R1826 B.n1267 B.n16 30.5
R1827 B.n1267 B.n1266 30.5
R1828 B.n1266 B.n1265 30.5
R1829 B.n1265 B.n23 30.5
R1830 B.n1259 B.n23 30.5
R1831 B.n1259 B.n1258 30.5
R1832 B.n1257 B.n30 30.5
R1833 B.n1251 B.n30 30.5
R1834 B.n1251 B.n1250 30.5
R1835 B.n1250 B.n1249 30.5
R1836 B.n1249 B.n37 30.5
R1837 B.n1243 B.n37 30.5
R1838 B.n1243 B.n1242 30.5
R1839 B.n1242 B.n1241 30.5
R1840 B.n1235 B.n47 30.5
R1841 B.n1235 B.n1234 30.5
R1842 B.n1234 B.n1233 30.5
R1843 B.n1233 B.n51 30.5
R1844 B.n1227 B.n51 30.5
R1845 B.n1227 B.n1226 30.5
R1846 B.n1226 B.n1225 30.5
R1847 B.n1219 B.n61 30.5
R1848 B.n1219 B.n1218 30.5
R1849 B.n1218 B.n1217 30.5
R1850 B.n1217 B.n65 30.5
R1851 B.n1211 B.n65 30.5
R1852 B.n1211 B.n1210 30.5
R1853 B.n1210 B.n1209 30.5
R1854 B.n1209 B.n72 30.5
R1855 B.n1203 B.n1202 30.5
R1856 B.n1202 B.n1201 30.5
R1857 B.n1201 B.n79 30.5
R1858 B.n1195 B.n79 30.5
R1859 B.n1195 B.n1194 30.5
R1860 B.n1194 B.n1193 30.5
R1861 B.n1193 B.n86 30.5
R1862 B.n1187 B.n86 30.5
R1863 B.n1187 B.n1186 30.5
R1864 B.n1186 B.n1185 30.5
R1865 B.n1185 B.n93 30.5
R1866 B.n1179 B.n1178 30.5
R1867 B.n1178 B.n1177 30.5
R1868 B.n1177 B.n100 30.5
R1869 B.n1171 B.n100 30.5
R1870 B.n1171 B.n1170 30.5
R1871 B.n1170 B.n1169 30.5
R1872 B.n1169 B.n107 30.5
R1873 B.n994 B.t5 29.1544
R1874 B.n1225 B.t1 29.1544
R1875 B.t3 B.n470 27.3603
R1876 B.n1258 B.t9 27.3603
R1877 B.n927 B.t15 23.7722
R1878 B.n1179 B.t11 23.7722
R1879 B.n1067 B.t4 19.2869
R1880 B.t0 B.n1273 19.2869
R1881 B B.n1287 18.0485
R1882 B.n1012 B.t7 17.4929
R1883 B.n47 B.t6 17.4929
R1884 B.n963 B.t8 15.6988
R1885 B.n1203 B.t2 15.6988
R1886 B.t8 B.n520 14.8017
R1887 B.t2 B.n72 14.8017
R1888 B.n1019 B.t7 13.0076
R1889 B.n1241 B.t6 13.0076
R1890 B.t4 B.n454 11.2135
R1891 B.n1274 B.t0 11.2135
R1892 B.n907 B.n906 10.6151
R1893 B.n907 B.n554 10.6151
R1894 B.n917 B.n554 10.6151
R1895 B.n918 B.n917 10.6151
R1896 B.n919 B.n918 10.6151
R1897 B.n919 B.n546 10.6151
R1898 B.n929 B.n546 10.6151
R1899 B.n930 B.n929 10.6151
R1900 B.n931 B.n930 10.6151
R1901 B.n931 B.n538 10.6151
R1902 B.n941 B.n538 10.6151
R1903 B.n942 B.n941 10.6151
R1904 B.n943 B.n942 10.6151
R1905 B.n943 B.n530 10.6151
R1906 B.n953 B.n530 10.6151
R1907 B.n954 B.n953 10.6151
R1908 B.n955 B.n954 10.6151
R1909 B.n955 B.n522 10.6151
R1910 B.n965 B.n522 10.6151
R1911 B.n966 B.n965 10.6151
R1912 B.n967 B.n966 10.6151
R1913 B.n967 B.n514 10.6151
R1914 B.n977 B.n514 10.6151
R1915 B.n978 B.n977 10.6151
R1916 B.n979 B.n978 10.6151
R1917 B.n979 B.n506 10.6151
R1918 B.n990 B.n506 10.6151
R1919 B.n991 B.n990 10.6151
R1920 B.n992 B.n991 10.6151
R1921 B.n992 B.n499 10.6151
R1922 B.n1002 B.n499 10.6151
R1923 B.n1003 B.n1002 10.6151
R1924 B.n1004 B.n1003 10.6151
R1925 B.n1004 B.n491 10.6151
R1926 B.n1015 B.n491 10.6151
R1927 B.n1016 B.n1015 10.6151
R1928 B.n1017 B.n1016 10.6151
R1929 B.n1017 B.n484 10.6151
R1930 B.n1027 B.n484 10.6151
R1931 B.n1028 B.n1027 10.6151
R1932 B.n1029 B.n1028 10.6151
R1933 B.n1029 B.n476 10.6151
R1934 B.n1039 B.n476 10.6151
R1935 B.n1040 B.n1039 10.6151
R1936 B.n1041 B.n1040 10.6151
R1937 B.n1041 B.n468 10.6151
R1938 B.n1051 B.n468 10.6151
R1939 B.n1052 B.n1051 10.6151
R1940 B.n1053 B.n1052 10.6151
R1941 B.n1053 B.n460 10.6151
R1942 B.n1063 B.n460 10.6151
R1943 B.n1064 B.n1063 10.6151
R1944 B.n1065 B.n1064 10.6151
R1945 B.n1065 B.n452 10.6151
R1946 B.n1076 B.n452 10.6151
R1947 B.n1077 B.n1076 10.6151
R1948 B.n1078 B.n1077 10.6151
R1949 B.n1078 B.n0 10.6151
R1950 B.n905 B.n562 10.6151
R1951 B.n900 B.n562 10.6151
R1952 B.n900 B.n899 10.6151
R1953 B.n899 B.n898 10.6151
R1954 B.n898 B.n895 10.6151
R1955 B.n895 B.n894 10.6151
R1956 B.n894 B.n891 10.6151
R1957 B.n891 B.n890 10.6151
R1958 B.n890 B.n887 10.6151
R1959 B.n887 B.n886 10.6151
R1960 B.n886 B.n883 10.6151
R1961 B.n883 B.n882 10.6151
R1962 B.n882 B.n879 10.6151
R1963 B.n879 B.n878 10.6151
R1964 B.n878 B.n875 10.6151
R1965 B.n875 B.n874 10.6151
R1966 B.n874 B.n871 10.6151
R1967 B.n871 B.n870 10.6151
R1968 B.n870 B.n867 10.6151
R1969 B.n867 B.n866 10.6151
R1970 B.n866 B.n863 10.6151
R1971 B.n863 B.n862 10.6151
R1972 B.n862 B.n859 10.6151
R1973 B.n859 B.n858 10.6151
R1974 B.n858 B.n855 10.6151
R1975 B.n855 B.n854 10.6151
R1976 B.n854 B.n851 10.6151
R1977 B.n851 B.n850 10.6151
R1978 B.n850 B.n847 10.6151
R1979 B.n847 B.n846 10.6151
R1980 B.n846 B.n843 10.6151
R1981 B.n843 B.n842 10.6151
R1982 B.n842 B.n839 10.6151
R1983 B.n839 B.n838 10.6151
R1984 B.n838 B.n835 10.6151
R1985 B.n835 B.n834 10.6151
R1986 B.n834 B.n831 10.6151
R1987 B.n831 B.n830 10.6151
R1988 B.n830 B.n827 10.6151
R1989 B.n827 B.n826 10.6151
R1990 B.n826 B.n823 10.6151
R1991 B.n823 B.n822 10.6151
R1992 B.n822 B.n819 10.6151
R1993 B.n819 B.n818 10.6151
R1994 B.n818 B.n815 10.6151
R1995 B.n815 B.n814 10.6151
R1996 B.n814 B.n811 10.6151
R1997 B.n811 B.n810 10.6151
R1998 B.n810 B.n807 10.6151
R1999 B.n807 B.n806 10.6151
R2000 B.n806 B.n803 10.6151
R2001 B.n803 B.n802 10.6151
R2002 B.n802 B.n799 10.6151
R2003 B.n799 B.n798 10.6151
R2004 B.n798 B.n795 10.6151
R2005 B.n795 B.n794 10.6151
R2006 B.n794 B.n791 10.6151
R2007 B.n791 B.n790 10.6151
R2008 B.n790 B.n787 10.6151
R2009 B.n787 B.n786 10.6151
R2010 B.n786 B.n783 10.6151
R2011 B.n783 B.n782 10.6151
R2012 B.n779 B.n778 10.6151
R2013 B.n778 B.n775 10.6151
R2014 B.n775 B.n774 10.6151
R2015 B.n774 B.n771 10.6151
R2016 B.n771 B.n770 10.6151
R2017 B.n770 B.n767 10.6151
R2018 B.n767 B.n766 10.6151
R2019 B.n766 B.n763 10.6151
R2020 B.n761 B.n758 10.6151
R2021 B.n758 B.n757 10.6151
R2022 B.n757 B.n754 10.6151
R2023 B.n754 B.n753 10.6151
R2024 B.n753 B.n750 10.6151
R2025 B.n750 B.n749 10.6151
R2026 B.n749 B.n746 10.6151
R2027 B.n746 B.n745 10.6151
R2028 B.n745 B.n742 10.6151
R2029 B.n742 B.n741 10.6151
R2030 B.n741 B.n738 10.6151
R2031 B.n738 B.n737 10.6151
R2032 B.n737 B.n734 10.6151
R2033 B.n734 B.n733 10.6151
R2034 B.n733 B.n730 10.6151
R2035 B.n730 B.n729 10.6151
R2036 B.n729 B.n726 10.6151
R2037 B.n726 B.n725 10.6151
R2038 B.n725 B.n722 10.6151
R2039 B.n722 B.n721 10.6151
R2040 B.n721 B.n718 10.6151
R2041 B.n718 B.n717 10.6151
R2042 B.n717 B.n714 10.6151
R2043 B.n714 B.n713 10.6151
R2044 B.n713 B.n710 10.6151
R2045 B.n710 B.n709 10.6151
R2046 B.n709 B.n706 10.6151
R2047 B.n706 B.n705 10.6151
R2048 B.n705 B.n702 10.6151
R2049 B.n702 B.n701 10.6151
R2050 B.n701 B.n698 10.6151
R2051 B.n698 B.n697 10.6151
R2052 B.n697 B.n694 10.6151
R2053 B.n694 B.n693 10.6151
R2054 B.n693 B.n690 10.6151
R2055 B.n690 B.n689 10.6151
R2056 B.n689 B.n686 10.6151
R2057 B.n686 B.n685 10.6151
R2058 B.n685 B.n682 10.6151
R2059 B.n682 B.n681 10.6151
R2060 B.n681 B.n678 10.6151
R2061 B.n678 B.n677 10.6151
R2062 B.n677 B.n674 10.6151
R2063 B.n674 B.n673 10.6151
R2064 B.n673 B.n670 10.6151
R2065 B.n670 B.n669 10.6151
R2066 B.n669 B.n666 10.6151
R2067 B.n666 B.n665 10.6151
R2068 B.n665 B.n662 10.6151
R2069 B.n662 B.n661 10.6151
R2070 B.n661 B.n658 10.6151
R2071 B.n658 B.n657 10.6151
R2072 B.n657 B.n654 10.6151
R2073 B.n654 B.n653 10.6151
R2074 B.n653 B.n650 10.6151
R2075 B.n650 B.n649 10.6151
R2076 B.n649 B.n646 10.6151
R2077 B.n646 B.n645 10.6151
R2078 B.n645 B.n642 10.6151
R2079 B.n642 B.n641 10.6151
R2080 B.n641 B.n638 10.6151
R2081 B.n638 B.n637 10.6151
R2082 B.n911 B.n558 10.6151
R2083 B.n912 B.n911 10.6151
R2084 B.n913 B.n912 10.6151
R2085 B.n913 B.n550 10.6151
R2086 B.n923 B.n550 10.6151
R2087 B.n924 B.n923 10.6151
R2088 B.n925 B.n924 10.6151
R2089 B.n925 B.n542 10.6151
R2090 B.n935 B.n542 10.6151
R2091 B.n936 B.n935 10.6151
R2092 B.n937 B.n936 10.6151
R2093 B.n937 B.n534 10.6151
R2094 B.n947 B.n534 10.6151
R2095 B.n948 B.n947 10.6151
R2096 B.n949 B.n948 10.6151
R2097 B.n949 B.n526 10.6151
R2098 B.n959 B.n526 10.6151
R2099 B.n960 B.n959 10.6151
R2100 B.n961 B.n960 10.6151
R2101 B.n961 B.n518 10.6151
R2102 B.n971 B.n518 10.6151
R2103 B.n972 B.n971 10.6151
R2104 B.n973 B.n972 10.6151
R2105 B.n973 B.n510 10.6151
R2106 B.n983 B.n510 10.6151
R2107 B.n984 B.n983 10.6151
R2108 B.n985 B.n984 10.6151
R2109 B.n985 B.n503 10.6151
R2110 B.n996 B.n503 10.6151
R2111 B.n997 B.n996 10.6151
R2112 B.n998 B.n997 10.6151
R2113 B.n998 B.n495 10.6151
R2114 B.n1008 B.n495 10.6151
R2115 B.n1009 B.n1008 10.6151
R2116 B.n1010 B.n1009 10.6151
R2117 B.n1010 B.n488 10.6151
R2118 B.n1021 B.n488 10.6151
R2119 B.n1022 B.n1021 10.6151
R2120 B.n1023 B.n1022 10.6151
R2121 B.n1023 B.n480 10.6151
R2122 B.n1033 B.n480 10.6151
R2123 B.n1034 B.n1033 10.6151
R2124 B.n1035 B.n1034 10.6151
R2125 B.n1035 B.n472 10.6151
R2126 B.n1045 B.n472 10.6151
R2127 B.n1046 B.n1045 10.6151
R2128 B.n1047 B.n1046 10.6151
R2129 B.n1047 B.n464 10.6151
R2130 B.n1057 B.n464 10.6151
R2131 B.n1058 B.n1057 10.6151
R2132 B.n1059 B.n1058 10.6151
R2133 B.n1059 B.n456 10.6151
R2134 B.n1069 B.n456 10.6151
R2135 B.n1070 B.n1069 10.6151
R2136 B.n1072 B.n1070 10.6151
R2137 B.n1072 B.n1071 10.6151
R2138 B.n1071 B.n448 10.6151
R2139 B.n1083 B.n448 10.6151
R2140 B.n1084 B.n1083 10.6151
R2141 B.n1085 B.n1084 10.6151
R2142 B.n1086 B.n1085 10.6151
R2143 B.n1087 B.n1086 10.6151
R2144 B.n1090 B.n1087 10.6151
R2145 B.n1091 B.n1090 10.6151
R2146 B.n1092 B.n1091 10.6151
R2147 B.n1093 B.n1092 10.6151
R2148 B.n1095 B.n1093 10.6151
R2149 B.n1096 B.n1095 10.6151
R2150 B.n1097 B.n1096 10.6151
R2151 B.n1098 B.n1097 10.6151
R2152 B.n1100 B.n1098 10.6151
R2153 B.n1101 B.n1100 10.6151
R2154 B.n1102 B.n1101 10.6151
R2155 B.n1103 B.n1102 10.6151
R2156 B.n1105 B.n1103 10.6151
R2157 B.n1106 B.n1105 10.6151
R2158 B.n1107 B.n1106 10.6151
R2159 B.n1108 B.n1107 10.6151
R2160 B.n1110 B.n1108 10.6151
R2161 B.n1111 B.n1110 10.6151
R2162 B.n1112 B.n1111 10.6151
R2163 B.n1113 B.n1112 10.6151
R2164 B.n1115 B.n1113 10.6151
R2165 B.n1116 B.n1115 10.6151
R2166 B.n1117 B.n1116 10.6151
R2167 B.n1118 B.n1117 10.6151
R2168 B.n1120 B.n1118 10.6151
R2169 B.n1121 B.n1120 10.6151
R2170 B.n1122 B.n1121 10.6151
R2171 B.n1123 B.n1122 10.6151
R2172 B.n1125 B.n1123 10.6151
R2173 B.n1126 B.n1125 10.6151
R2174 B.n1127 B.n1126 10.6151
R2175 B.n1128 B.n1127 10.6151
R2176 B.n1130 B.n1128 10.6151
R2177 B.n1131 B.n1130 10.6151
R2178 B.n1132 B.n1131 10.6151
R2179 B.n1133 B.n1132 10.6151
R2180 B.n1135 B.n1133 10.6151
R2181 B.n1136 B.n1135 10.6151
R2182 B.n1137 B.n1136 10.6151
R2183 B.n1138 B.n1137 10.6151
R2184 B.n1140 B.n1138 10.6151
R2185 B.n1141 B.n1140 10.6151
R2186 B.n1142 B.n1141 10.6151
R2187 B.n1143 B.n1142 10.6151
R2188 B.n1145 B.n1143 10.6151
R2189 B.n1146 B.n1145 10.6151
R2190 B.n1147 B.n1146 10.6151
R2191 B.n1148 B.n1147 10.6151
R2192 B.n1150 B.n1148 10.6151
R2193 B.n1151 B.n1150 10.6151
R2194 B.n1152 B.n1151 10.6151
R2195 B.n1153 B.n1152 10.6151
R2196 B.n1155 B.n1153 10.6151
R2197 B.n1156 B.n1155 10.6151
R2198 B.n1157 B.n1156 10.6151
R2199 B.n1158 B.n1157 10.6151
R2200 B.n1159 B.n1158 10.6151
R2201 B.n1279 B.n1 10.6151
R2202 B.n1279 B.n1278 10.6151
R2203 B.n1278 B.n1277 10.6151
R2204 B.n1277 B.n10 10.6151
R2205 B.n1271 B.n10 10.6151
R2206 B.n1271 B.n1270 10.6151
R2207 B.n1270 B.n1269 10.6151
R2208 B.n1269 B.n18 10.6151
R2209 B.n1263 B.n18 10.6151
R2210 B.n1263 B.n1262 10.6151
R2211 B.n1262 B.n1261 10.6151
R2212 B.n1261 B.n25 10.6151
R2213 B.n1255 B.n25 10.6151
R2214 B.n1255 B.n1254 10.6151
R2215 B.n1254 B.n1253 10.6151
R2216 B.n1253 B.n32 10.6151
R2217 B.n1247 B.n32 10.6151
R2218 B.n1247 B.n1246 10.6151
R2219 B.n1246 B.n1245 10.6151
R2220 B.n1245 B.n39 10.6151
R2221 B.n1239 B.n39 10.6151
R2222 B.n1239 B.n1238 10.6151
R2223 B.n1238 B.n1237 10.6151
R2224 B.n1237 B.n45 10.6151
R2225 B.n1231 B.n45 10.6151
R2226 B.n1231 B.n1230 10.6151
R2227 B.n1230 B.n1229 10.6151
R2228 B.n1229 B.n53 10.6151
R2229 B.n1223 B.n53 10.6151
R2230 B.n1223 B.n1222 10.6151
R2231 B.n1222 B.n1221 10.6151
R2232 B.n1221 B.n59 10.6151
R2233 B.n1215 B.n59 10.6151
R2234 B.n1215 B.n1214 10.6151
R2235 B.n1214 B.n1213 10.6151
R2236 B.n1213 B.n67 10.6151
R2237 B.n1207 B.n67 10.6151
R2238 B.n1207 B.n1206 10.6151
R2239 B.n1206 B.n1205 10.6151
R2240 B.n1205 B.n74 10.6151
R2241 B.n1199 B.n74 10.6151
R2242 B.n1199 B.n1198 10.6151
R2243 B.n1198 B.n1197 10.6151
R2244 B.n1197 B.n81 10.6151
R2245 B.n1191 B.n81 10.6151
R2246 B.n1191 B.n1190 10.6151
R2247 B.n1190 B.n1189 10.6151
R2248 B.n1189 B.n88 10.6151
R2249 B.n1183 B.n88 10.6151
R2250 B.n1183 B.n1182 10.6151
R2251 B.n1182 B.n1181 10.6151
R2252 B.n1181 B.n95 10.6151
R2253 B.n1175 B.n95 10.6151
R2254 B.n1175 B.n1174 10.6151
R2255 B.n1174 B.n1173 10.6151
R2256 B.n1173 B.n102 10.6151
R2257 B.n1167 B.n102 10.6151
R2258 B.n1167 B.n1166 10.6151
R2259 B.n1165 B.n109 10.6151
R2260 B.n185 B.n109 10.6151
R2261 B.n186 B.n185 10.6151
R2262 B.n189 B.n186 10.6151
R2263 B.n190 B.n189 10.6151
R2264 B.n193 B.n190 10.6151
R2265 B.n194 B.n193 10.6151
R2266 B.n197 B.n194 10.6151
R2267 B.n198 B.n197 10.6151
R2268 B.n201 B.n198 10.6151
R2269 B.n202 B.n201 10.6151
R2270 B.n205 B.n202 10.6151
R2271 B.n206 B.n205 10.6151
R2272 B.n209 B.n206 10.6151
R2273 B.n210 B.n209 10.6151
R2274 B.n213 B.n210 10.6151
R2275 B.n214 B.n213 10.6151
R2276 B.n217 B.n214 10.6151
R2277 B.n218 B.n217 10.6151
R2278 B.n221 B.n218 10.6151
R2279 B.n222 B.n221 10.6151
R2280 B.n225 B.n222 10.6151
R2281 B.n226 B.n225 10.6151
R2282 B.n229 B.n226 10.6151
R2283 B.n230 B.n229 10.6151
R2284 B.n233 B.n230 10.6151
R2285 B.n234 B.n233 10.6151
R2286 B.n237 B.n234 10.6151
R2287 B.n238 B.n237 10.6151
R2288 B.n241 B.n238 10.6151
R2289 B.n242 B.n241 10.6151
R2290 B.n245 B.n242 10.6151
R2291 B.n246 B.n245 10.6151
R2292 B.n249 B.n246 10.6151
R2293 B.n250 B.n249 10.6151
R2294 B.n253 B.n250 10.6151
R2295 B.n254 B.n253 10.6151
R2296 B.n257 B.n254 10.6151
R2297 B.n258 B.n257 10.6151
R2298 B.n261 B.n258 10.6151
R2299 B.n262 B.n261 10.6151
R2300 B.n265 B.n262 10.6151
R2301 B.n266 B.n265 10.6151
R2302 B.n269 B.n266 10.6151
R2303 B.n270 B.n269 10.6151
R2304 B.n273 B.n270 10.6151
R2305 B.n274 B.n273 10.6151
R2306 B.n277 B.n274 10.6151
R2307 B.n278 B.n277 10.6151
R2308 B.n281 B.n278 10.6151
R2309 B.n282 B.n281 10.6151
R2310 B.n285 B.n282 10.6151
R2311 B.n286 B.n285 10.6151
R2312 B.n289 B.n286 10.6151
R2313 B.n290 B.n289 10.6151
R2314 B.n293 B.n290 10.6151
R2315 B.n294 B.n293 10.6151
R2316 B.n297 B.n294 10.6151
R2317 B.n298 B.n297 10.6151
R2318 B.n301 B.n298 10.6151
R2319 B.n302 B.n301 10.6151
R2320 B.n305 B.n302 10.6151
R2321 B.n310 B.n307 10.6151
R2322 B.n311 B.n310 10.6151
R2323 B.n314 B.n311 10.6151
R2324 B.n315 B.n314 10.6151
R2325 B.n318 B.n315 10.6151
R2326 B.n319 B.n318 10.6151
R2327 B.n322 B.n319 10.6151
R2328 B.n323 B.n322 10.6151
R2329 B.n327 B.n326 10.6151
R2330 B.n330 B.n327 10.6151
R2331 B.n331 B.n330 10.6151
R2332 B.n334 B.n331 10.6151
R2333 B.n335 B.n334 10.6151
R2334 B.n338 B.n335 10.6151
R2335 B.n339 B.n338 10.6151
R2336 B.n342 B.n339 10.6151
R2337 B.n343 B.n342 10.6151
R2338 B.n346 B.n343 10.6151
R2339 B.n347 B.n346 10.6151
R2340 B.n350 B.n347 10.6151
R2341 B.n351 B.n350 10.6151
R2342 B.n354 B.n351 10.6151
R2343 B.n355 B.n354 10.6151
R2344 B.n358 B.n355 10.6151
R2345 B.n359 B.n358 10.6151
R2346 B.n362 B.n359 10.6151
R2347 B.n363 B.n362 10.6151
R2348 B.n366 B.n363 10.6151
R2349 B.n367 B.n366 10.6151
R2350 B.n370 B.n367 10.6151
R2351 B.n371 B.n370 10.6151
R2352 B.n374 B.n371 10.6151
R2353 B.n375 B.n374 10.6151
R2354 B.n378 B.n375 10.6151
R2355 B.n379 B.n378 10.6151
R2356 B.n382 B.n379 10.6151
R2357 B.n383 B.n382 10.6151
R2358 B.n386 B.n383 10.6151
R2359 B.n387 B.n386 10.6151
R2360 B.n390 B.n387 10.6151
R2361 B.n391 B.n390 10.6151
R2362 B.n394 B.n391 10.6151
R2363 B.n395 B.n394 10.6151
R2364 B.n398 B.n395 10.6151
R2365 B.n399 B.n398 10.6151
R2366 B.n402 B.n399 10.6151
R2367 B.n403 B.n402 10.6151
R2368 B.n406 B.n403 10.6151
R2369 B.n407 B.n406 10.6151
R2370 B.n410 B.n407 10.6151
R2371 B.n411 B.n410 10.6151
R2372 B.n414 B.n411 10.6151
R2373 B.n415 B.n414 10.6151
R2374 B.n418 B.n415 10.6151
R2375 B.n419 B.n418 10.6151
R2376 B.n422 B.n419 10.6151
R2377 B.n423 B.n422 10.6151
R2378 B.n426 B.n423 10.6151
R2379 B.n427 B.n426 10.6151
R2380 B.n430 B.n427 10.6151
R2381 B.n431 B.n430 10.6151
R2382 B.n434 B.n431 10.6151
R2383 B.n435 B.n434 10.6151
R2384 B.n438 B.n435 10.6151
R2385 B.n439 B.n438 10.6151
R2386 B.n442 B.n439 10.6151
R2387 B.n443 B.n442 10.6151
R2388 B.n446 B.n443 10.6151
R2389 B.n447 B.n446 10.6151
R2390 B.n1160 B.n447 10.6151
R2391 B.n1287 B.n0 8.11757
R2392 B.n1287 B.n1 8.11757
R2393 B.t15 B.n544 6.72833
R2394 B.t11 B.n93 6.72833
R2395 B.n779 B.n633 6.5566
R2396 B.n763 B.n762 6.5566
R2397 B.n307 B.n306 6.5566
R2398 B.n323 B.n181 6.5566
R2399 B.n782 B.n633 4.05904
R2400 B.n762 B.n761 4.05904
R2401 B.n306 B.n305 4.05904
R2402 B.n326 B.n181 4.05904
R2403 B.n1043 B.t3 3.14015
R2404 B.t9 B.n1257 3.14015
R2405 B.n987 B.t5 1.34607
R2406 B.n61 B.t1 1.34607
R2407 VN.n11 VN.t4 211.549
R2408 VN.n53 VN.t9 211.549
R2409 VN.n10 VN.t3 180.517
R2410 VN.n21 VN.t2 180.517
R2411 VN.n3 VN.t8 180.517
R2412 VN.n40 VN.t6 180.517
R2413 VN.n52 VN.t5 180.517
R2414 VN.n63 VN.t1 180.517
R2415 VN.n45 VN.t7 180.517
R2416 VN.n82 VN.t0 180.517
R2417 VN.n81 VN.n42 161.3
R2418 VN.n80 VN.n79 161.3
R2419 VN.n78 VN.n43 161.3
R2420 VN.n77 VN.n76 161.3
R2421 VN.n75 VN.n44 161.3
R2422 VN.n74 VN.n73 161.3
R2423 VN.n72 VN.n71 161.3
R2424 VN.n70 VN.n46 161.3
R2425 VN.n69 VN.n68 161.3
R2426 VN.n67 VN.n47 161.3
R2427 VN.n66 VN.n65 161.3
R2428 VN.n64 VN.n48 161.3
R2429 VN.n62 VN.n61 161.3
R2430 VN.n60 VN.n49 161.3
R2431 VN.n59 VN.n58 161.3
R2432 VN.n57 VN.n50 161.3
R2433 VN.n56 VN.n55 161.3
R2434 VN.n54 VN.n51 161.3
R2435 VN.n39 VN.n0 161.3
R2436 VN.n38 VN.n37 161.3
R2437 VN.n36 VN.n1 161.3
R2438 VN.n35 VN.n34 161.3
R2439 VN.n33 VN.n2 161.3
R2440 VN.n32 VN.n31 161.3
R2441 VN.n30 VN.n29 161.3
R2442 VN.n28 VN.n4 161.3
R2443 VN.n27 VN.n26 161.3
R2444 VN.n25 VN.n5 161.3
R2445 VN.n24 VN.n23 161.3
R2446 VN.n22 VN.n6 161.3
R2447 VN.n20 VN.n19 161.3
R2448 VN.n18 VN.n7 161.3
R2449 VN.n17 VN.n16 161.3
R2450 VN.n15 VN.n8 161.3
R2451 VN.n14 VN.n13 161.3
R2452 VN.n12 VN.n9 161.3
R2453 VN.n41 VN.n40 108.309
R2454 VN.n83 VN.n82 108.309
R2455 VN.n11 VN.n10 65.3454
R2456 VN.n53 VN.n52 65.3454
R2457 VN VN.n83 58.6194
R2458 VN.n16 VN.n15 56.5193
R2459 VN.n27 VN.n5 56.5193
R2460 VN.n58 VN.n57 56.5193
R2461 VN.n69 VN.n47 56.5193
R2462 VN.n34 VN.n1 50.2061
R2463 VN.n76 VN.n43 50.2061
R2464 VN.n34 VN.n33 30.7807
R2465 VN.n76 VN.n75 30.7807
R2466 VN.n14 VN.n9 24.4675
R2467 VN.n15 VN.n14 24.4675
R2468 VN.n16 VN.n7 24.4675
R2469 VN.n20 VN.n7 24.4675
R2470 VN.n23 VN.n22 24.4675
R2471 VN.n23 VN.n5 24.4675
R2472 VN.n28 VN.n27 24.4675
R2473 VN.n29 VN.n28 24.4675
R2474 VN.n33 VN.n32 24.4675
R2475 VN.n38 VN.n1 24.4675
R2476 VN.n39 VN.n38 24.4675
R2477 VN.n57 VN.n56 24.4675
R2478 VN.n56 VN.n51 24.4675
R2479 VN.n65 VN.n47 24.4675
R2480 VN.n65 VN.n64 24.4675
R2481 VN.n62 VN.n49 24.4675
R2482 VN.n58 VN.n49 24.4675
R2483 VN.n75 VN.n74 24.4675
R2484 VN.n71 VN.n70 24.4675
R2485 VN.n70 VN.n69 24.4675
R2486 VN.n81 VN.n80 24.4675
R2487 VN.n80 VN.n43 24.4675
R2488 VN.n32 VN.n3 17.1274
R2489 VN.n74 VN.n45 17.1274
R2490 VN.n21 VN.n20 12.234
R2491 VN.n22 VN.n21 12.234
R2492 VN.n64 VN.n63 12.234
R2493 VN.n63 VN.n62 12.234
R2494 VN.n10 VN.n9 7.3406
R2495 VN.n29 VN.n3 7.3406
R2496 VN.n52 VN.n51 7.3406
R2497 VN.n71 VN.n45 7.3406
R2498 VN.n54 VN.n53 7.32785
R2499 VN.n12 VN.n11 7.32785
R2500 VN.n40 VN.n39 2.4472
R2501 VN.n82 VN.n81 2.4472
R2502 VN.n83 VN.n42 0.278367
R2503 VN.n41 VN.n0 0.278367
R2504 VN.n79 VN.n42 0.189894
R2505 VN.n79 VN.n78 0.189894
R2506 VN.n78 VN.n77 0.189894
R2507 VN.n77 VN.n44 0.189894
R2508 VN.n73 VN.n44 0.189894
R2509 VN.n73 VN.n72 0.189894
R2510 VN.n72 VN.n46 0.189894
R2511 VN.n68 VN.n46 0.189894
R2512 VN.n68 VN.n67 0.189894
R2513 VN.n67 VN.n66 0.189894
R2514 VN.n66 VN.n48 0.189894
R2515 VN.n61 VN.n48 0.189894
R2516 VN.n61 VN.n60 0.189894
R2517 VN.n60 VN.n59 0.189894
R2518 VN.n59 VN.n50 0.189894
R2519 VN.n55 VN.n50 0.189894
R2520 VN.n55 VN.n54 0.189894
R2521 VN.n13 VN.n12 0.189894
R2522 VN.n13 VN.n8 0.189894
R2523 VN.n17 VN.n8 0.189894
R2524 VN.n18 VN.n17 0.189894
R2525 VN.n19 VN.n18 0.189894
R2526 VN.n19 VN.n6 0.189894
R2527 VN.n24 VN.n6 0.189894
R2528 VN.n25 VN.n24 0.189894
R2529 VN.n26 VN.n25 0.189894
R2530 VN.n26 VN.n4 0.189894
R2531 VN.n30 VN.n4 0.189894
R2532 VN.n31 VN.n30 0.189894
R2533 VN.n31 VN.n2 0.189894
R2534 VN.n35 VN.n2 0.189894
R2535 VN.n36 VN.n35 0.189894
R2536 VN.n37 VN.n36 0.189894
R2537 VN.n37 VN.n0 0.189894
R2538 VN VN.n41 0.153454
R2539 VDD2.n1 VDD2.t5 62.7819
R2540 VDD2.n3 VDD2.n2 61.0732
R2541 VDD2 VDD2.n7 61.0702
R2542 VDD2.n4 VDD2.t9 60.2821
R2543 VDD2.n6 VDD2.n5 59.2536
R2544 VDD2.n1 VDD2.n0 59.2535
R2545 VDD2.n4 VDD2.n3 52.1851
R2546 VDD2.n6 VDD2.n4 2.5005
R2547 VDD2.n7 VDD2.t4 1.02907
R2548 VDD2.n7 VDD2.t0 1.02907
R2549 VDD2.n5 VDD2.t2 1.02907
R2550 VDD2.n5 VDD2.t8 1.02907
R2551 VDD2.n2 VDD2.t1 1.02907
R2552 VDD2.n2 VDD2.t3 1.02907
R2553 VDD2.n0 VDD2.t6 1.02907
R2554 VDD2.n0 VDD2.t7 1.02907
R2555 VDD2 VDD2.n6 0.68369
R2556 VDD2.n3 VDD2.n1 0.570154
C0 VP VTAIL 17.082f
C1 VTAIL VDD2 13.799f
C2 VN VTAIL 17.0676f
C3 VTAIL VDD1 13.75f
C4 VP VDD2 0.580372f
C5 VP VN 9.70121f
C6 VP VDD1 17.184f
C7 VN VDD2 16.7621f
C8 VDD1 VDD2 2.15596f
C9 VN VDD1 0.153326f
C10 VDD2 B 8.45626f
C11 VDD1 B 8.430911f
C12 VTAIL B 11.069127f
C13 VN B 18.617168f
C14 VP B 17.020077f
C15 VDD2.t5 B 4.1734f
C16 VDD2.t6 B 0.356061f
C17 VDD2.t7 B 0.356061f
C18 VDD2.n0 B 3.2499f
C19 VDD2.n1 B 0.873303f
C20 VDD2.t1 B 0.356061f
C21 VDD2.t3 B 0.356061f
C22 VDD2.n2 B 3.26578f
C23 VDD2.n3 B 3.13558f
C24 VDD2.t9 B 4.15502f
C25 VDD2.n4 B 3.4398f
C26 VDD2.t2 B 0.356061f
C27 VDD2.t8 B 0.356061f
C28 VDD2.n5 B 3.24989f
C29 VDD2.n6 B 0.437725f
C30 VDD2.t4 B 0.356061f
C31 VDD2.t0 B 0.356061f
C32 VDD2.n7 B 3.26573f
C33 VN.n0 B 0.027174f
C34 VN.t6 B 2.80822f
C35 VN.n1 B 0.03783f
C36 VN.n2 B 0.020612f
C37 VN.t8 B 2.80822f
C38 VN.n3 B 0.971534f
C39 VN.n4 B 0.020612f
C40 VN.n5 B 0.027218f
C41 VN.n6 B 0.020612f
C42 VN.t2 B 2.80822f
C43 VN.n7 B 0.038415f
C44 VN.n8 B 0.020612f
C45 VN.n9 B 0.025139f
C46 VN.t4 B 2.96897f
C47 VN.t3 B 2.80822f
C48 VN.n10 B 1.02739f
C49 VN.n11 B 1.01707f
C50 VN.n12 B 0.197983f
C51 VN.n13 B 0.020612f
C52 VN.n14 B 0.038415f
C53 VN.n15 B 0.032961f
C54 VN.n16 B 0.027218f
C55 VN.n17 B 0.020612f
C56 VN.n18 B 0.020612f
C57 VN.n19 B 0.020612f
C58 VN.n20 B 0.028932f
C59 VN.n21 B 0.971534f
C60 VN.n22 B 0.028932f
C61 VN.n23 B 0.038415f
C62 VN.n24 B 0.020612f
C63 VN.n25 B 0.020612f
C64 VN.n26 B 0.020612f
C65 VN.n27 B 0.032961f
C66 VN.n28 B 0.038415f
C67 VN.n29 B 0.025139f
C68 VN.n30 B 0.020612f
C69 VN.n31 B 0.020612f
C70 VN.n32 B 0.032725f
C71 VN.n33 B 0.041292f
C72 VN.n34 B 0.019471f
C73 VN.n35 B 0.020612f
C74 VN.n36 B 0.020612f
C75 VN.n37 B 0.020612f
C76 VN.n38 B 0.038415f
C77 VN.n39 B 0.021346f
C78 VN.n40 B 1.03166f
C79 VN.n41 B 0.036709f
C80 VN.n42 B 0.027174f
C81 VN.t0 B 2.80822f
C82 VN.n43 B 0.03783f
C83 VN.n44 B 0.020612f
C84 VN.t7 B 2.80822f
C85 VN.n45 B 0.971534f
C86 VN.n46 B 0.020612f
C87 VN.n47 B 0.027218f
C88 VN.n48 B 0.020612f
C89 VN.t1 B 2.80822f
C90 VN.n49 B 0.038415f
C91 VN.n50 B 0.020612f
C92 VN.n51 B 0.025139f
C93 VN.t9 B 2.96897f
C94 VN.t5 B 2.80822f
C95 VN.n52 B 1.02739f
C96 VN.n53 B 1.01707f
C97 VN.n54 B 0.197983f
C98 VN.n55 B 0.020612f
C99 VN.n56 B 0.038415f
C100 VN.n57 B 0.032961f
C101 VN.n58 B 0.027218f
C102 VN.n59 B 0.020612f
C103 VN.n60 B 0.020612f
C104 VN.n61 B 0.020612f
C105 VN.n62 B 0.028932f
C106 VN.n63 B 0.971534f
C107 VN.n64 B 0.028932f
C108 VN.n65 B 0.038415f
C109 VN.n66 B 0.020612f
C110 VN.n67 B 0.020612f
C111 VN.n68 B 0.020612f
C112 VN.n69 B 0.032961f
C113 VN.n70 B 0.038415f
C114 VN.n71 B 0.025139f
C115 VN.n72 B 0.020612f
C116 VN.n73 B 0.020612f
C117 VN.n74 B 0.032725f
C118 VN.n75 B 0.041292f
C119 VN.n76 B 0.019471f
C120 VN.n77 B 0.020612f
C121 VN.n78 B 0.020612f
C122 VN.n79 B 0.020612f
C123 VN.n80 B 0.038415f
C124 VN.n81 B 0.021346f
C125 VN.n82 B 1.03166f
C126 VN.n83 B 1.44076f
C127 VTAIL.t0 B 0.35771f
C128 VTAIL.t9 B 0.35771f
C129 VTAIL.n0 B 3.18891f
C130 VTAIL.n1 B 0.519414f
C131 VTAIL.t11 B 4.07467f
C132 VTAIL.n2 B 0.652174f
C133 VTAIL.t15 B 0.35771f
C134 VTAIL.t13 B 0.35771f
C135 VTAIL.n3 B 3.18891f
C136 VTAIL.n4 B 0.621476f
C137 VTAIL.t10 B 0.35771f
C138 VTAIL.t17 B 0.35771f
C139 VTAIL.n5 B 3.18891f
C140 VTAIL.n6 B 2.38773f
C141 VTAIL.t8 B 0.35771f
C142 VTAIL.t5 B 0.35771f
C143 VTAIL.n7 B 3.18891f
C144 VTAIL.n8 B 2.38774f
C145 VTAIL.t7 B 0.35771f
C146 VTAIL.t3 B 0.35771f
C147 VTAIL.n9 B 3.18891f
C148 VTAIL.n10 B 0.621483f
C149 VTAIL.t4 B 4.07468f
C150 VTAIL.n11 B 0.652169f
C151 VTAIL.t16 B 0.35771f
C152 VTAIL.t18 B 0.35771f
C153 VTAIL.n12 B 3.18891f
C154 VTAIL.n13 B 0.562369f
C155 VTAIL.t12 B 0.35771f
C156 VTAIL.t19 B 0.35771f
C157 VTAIL.n14 B 3.18891f
C158 VTAIL.n15 B 0.621483f
C159 VTAIL.t14 B 4.07467f
C160 VTAIL.n16 B 2.28812f
C161 VTAIL.t2 B 4.07467f
C162 VTAIL.n17 B 2.28812f
C163 VTAIL.t6 B 0.35771f
C164 VTAIL.t1 B 0.35771f
C165 VTAIL.n18 B 3.18891f
C166 VTAIL.n19 B 0.474996f
C167 VDD1.t2 B 4.2132f
C168 VDD1.t4 B 0.359456f
C169 VDD1.t8 B 0.359456f
C170 VDD1.n0 B 3.28088f
C171 VDD1.n1 B 0.889315f
C172 VDD1.t6 B 4.21319f
C173 VDD1.t3 B 0.359456f
C174 VDD1.t1 B 0.359456f
C175 VDD1.n2 B 3.28089f
C176 VDD1.n3 B 0.881629f
C177 VDD1.t9 B 0.359456f
C178 VDD1.t7 B 0.359456f
C179 VDD1.n4 B 3.29692f
C180 VDD1.n5 B 3.28686f
C181 VDD1.t5 B 0.359456f
C182 VDD1.t0 B 0.359456f
C183 VDD1.n6 B 3.28087f
C184 VDD1.n7 B 3.51025f
C185 VP.n0 B 0.027442f
C186 VP.t8 B 2.83587f
C187 VP.n1 B 0.038202f
C188 VP.n2 B 0.020815f
C189 VP.t6 B 2.83587f
C190 VP.n3 B 0.981099f
C191 VP.n4 B 0.020815f
C192 VP.n5 B 0.027485f
C193 VP.n6 B 0.020815f
C194 VP.t4 B 2.83587f
C195 VP.n7 B 0.038793f
C196 VP.n8 B 0.020815f
C197 VP.n9 B 0.025386f
C198 VP.n10 B 0.020815f
C199 VP.n11 B 0.038202f
C200 VP.n12 B 0.027442f
C201 VP.t9 B 2.83587f
C202 VP.n13 B 0.027442f
C203 VP.t5 B 2.83587f
C204 VP.n14 B 0.038202f
C205 VP.n15 B 0.020815f
C206 VP.t0 B 2.83587f
C207 VP.n16 B 0.981099f
C208 VP.n17 B 0.020815f
C209 VP.n18 B 0.027485f
C210 VP.n19 B 0.020815f
C211 VP.t7 B 2.83587f
C212 VP.n20 B 0.038793f
C213 VP.n21 B 0.020815f
C214 VP.n22 B 0.025386f
C215 VP.t3 B 2.9982f
C216 VP.t1 B 2.83587f
C217 VP.n23 B 1.03751f
C218 VP.n24 B 1.02709f
C219 VP.n25 B 0.199932f
C220 VP.n26 B 0.020815f
C221 VP.n27 B 0.038793f
C222 VP.n28 B 0.033286f
C223 VP.n29 B 0.027485f
C224 VP.n30 B 0.020815f
C225 VP.n31 B 0.020815f
C226 VP.n32 B 0.020815f
C227 VP.n33 B 0.029217f
C228 VP.n34 B 0.981099f
C229 VP.n35 B 0.029217f
C230 VP.n36 B 0.038793f
C231 VP.n37 B 0.020815f
C232 VP.n38 B 0.020815f
C233 VP.n39 B 0.020815f
C234 VP.n40 B 0.033286f
C235 VP.n41 B 0.038793f
C236 VP.n42 B 0.025386f
C237 VP.n43 B 0.020815f
C238 VP.n44 B 0.020815f
C239 VP.n45 B 0.033047f
C240 VP.n46 B 0.041699f
C241 VP.n47 B 0.019663f
C242 VP.n48 B 0.020815f
C243 VP.n49 B 0.020815f
C244 VP.n50 B 0.020815f
C245 VP.n51 B 0.038793f
C246 VP.n52 B 0.021556f
C247 VP.n53 B 1.04182f
C248 VP.n54 B 1.44401f
C249 VP.n55 B 1.45684f
C250 VP.n56 B 1.04182f
C251 VP.n57 B 0.021556f
C252 VP.n58 B 0.038793f
C253 VP.n59 B 0.020815f
C254 VP.n60 B 0.020815f
C255 VP.n61 B 0.020815f
C256 VP.n62 B 0.019663f
C257 VP.n63 B 0.041699f
C258 VP.t2 B 2.83587f
C259 VP.n64 B 0.981099f
C260 VP.n65 B 0.033047f
C261 VP.n66 B 0.020815f
C262 VP.n67 B 0.020815f
C263 VP.n68 B 0.020815f
C264 VP.n69 B 0.038793f
C265 VP.n70 B 0.033286f
C266 VP.n71 B 0.027485f
C267 VP.n72 B 0.020815f
C268 VP.n73 B 0.020815f
C269 VP.n74 B 0.020815f
C270 VP.n75 B 0.029217f
C271 VP.n76 B 0.981099f
C272 VP.n77 B 0.029217f
C273 VP.n78 B 0.038793f
C274 VP.n79 B 0.020815f
C275 VP.n80 B 0.020815f
C276 VP.n81 B 0.020815f
C277 VP.n82 B 0.033286f
C278 VP.n83 B 0.038793f
C279 VP.n84 B 0.025386f
C280 VP.n85 B 0.020815f
C281 VP.n86 B 0.020815f
C282 VP.n87 B 0.033047f
C283 VP.n88 B 0.041699f
C284 VP.n89 B 0.019663f
C285 VP.n90 B 0.020815f
C286 VP.n91 B 0.020815f
C287 VP.n92 B 0.020815f
C288 VP.n93 B 0.038793f
C289 VP.n94 B 0.021556f
C290 VP.n95 B 1.04182f
C291 VP.n96 B 0.03707f
.ends

