* NGSPICE file created from diff_pair_sample_1708.ext - technology: sky130A

.subckt diff_pair_sample_1708 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t9 w_n1634_n4096# sky130_fd_pr__pfet_01v8 ad=6.0996 pd=32.06 as=2.5806 ps=15.97 w=15.64 l=0.5
X1 B.t11 B.t9 B.t10 w_n1634_n4096# sky130_fd_pr__pfet_01v8 ad=6.0996 pd=32.06 as=0 ps=0 w=15.64 l=0.5
X2 VDD1.t4 VP.t1 VTAIL.t8 w_n1634_n4096# sky130_fd_pr__pfet_01v8 ad=6.0996 pd=32.06 as=2.5806 ps=15.97 w=15.64 l=0.5
X3 VDD2.t5 VN.t0 VTAIL.t5 w_n1634_n4096# sky130_fd_pr__pfet_01v8 ad=6.0996 pd=32.06 as=2.5806 ps=15.97 w=15.64 l=0.5
X4 B.t8 B.t6 B.t7 w_n1634_n4096# sky130_fd_pr__pfet_01v8 ad=6.0996 pd=32.06 as=0 ps=0 w=15.64 l=0.5
X5 B.t5 B.t3 B.t4 w_n1634_n4096# sky130_fd_pr__pfet_01v8 ad=6.0996 pd=32.06 as=0 ps=0 w=15.64 l=0.5
X6 VDD2.t4 VN.t1 VTAIL.t4 w_n1634_n4096# sky130_fd_pr__pfet_01v8 ad=2.5806 pd=15.97 as=6.0996 ps=32.06 w=15.64 l=0.5
X7 VDD2.t3 VN.t2 VTAIL.t0 w_n1634_n4096# sky130_fd_pr__pfet_01v8 ad=2.5806 pd=15.97 as=6.0996 ps=32.06 w=15.64 l=0.5
X8 VTAIL.t6 VP.t2 VDD1.t3 w_n1634_n4096# sky130_fd_pr__pfet_01v8 ad=2.5806 pd=15.97 as=2.5806 ps=15.97 w=15.64 l=0.5
X9 VDD1.t2 VP.t3 VTAIL.t11 w_n1634_n4096# sky130_fd_pr__pfet_01v8 ad=2.5806 pd=15.97 as=6.0996 ps=32.06 w=15.64 l=0.5
X10 VTAIL.t7 VP.t4 VDD1.t1 w_n1634_n4096# sky130_fd_pr__pfet_01v8 ad=2.5806 pd=15.97 as=2.5806 ps=15.97 w=15.64 l=0.5
X11 B.t2 B.t0 B.t1 w_n1634_n4096# sky130_fd_pr__pfet_01v8 ad=6.0996 pd=32.06 as=0 ps=0 w=15.64 l=0.5
X12 VDD1.t0 VP.t5 VTAIL.t10 w_n1634_n4096# sky130_fd_pr__pfet_01v8 ad=2.5806 pd=15.97 as=6.0996 ps=32.06 w=15.64 l=0.5
X13 VTAIL.t2 VN.t3 VDD2.t2 w_n1634_n4096# sky130_fd_pr__pfet_01v8 ad=2.5806 pd=15.97 as=2.5806 ps=15.97 w=15.64 l=0.5
X14 VTAIL.t3 VN.t4 VDD2.t1 w_n1634_n4096# sky130_fd_pr__pfet_01v8 ad=2.5806 pd=15.97 as=2.5806 ps=15.97 w=15.64 l=0.5
X15 VDD2.t0 VN.t5 VTAIL.t1 w_n1634_n4096# sky130_fd_pr__pfet_01v8 ad=6.0996 pd=32.06 as=2.5806 ps=15.97 w=15.64 l=0.5
R0 VP.n1 VP.t0 859.236
R1 VP.n6 VP.t1 832.414
R2 VP.n7 VP.t4 832.414
R3 VP.n8 VP.t5 832.414
R4 VP.n3 VP.t3 832.414
R5 VP.n2 VP.t2 832.414
R6 VP.n9 VP.n8 161.3
R7 VP.n4 VP.n3 161.3
R8 VP.n6 VP.n5 161.3
R9 VP.n7 VP.n0 80.6037
R10 VP.n7 VP.n6 48.2005
R11 VP.n8 VP.n7 48.2005
R12 VP.n3 VP.n2 48.2005
R13 VP.n4 VP.n1 45.1367
R14 VP.n5 VP.n4 43.1634
R15 VP.n2 VP.n1 13.3799
R16 VP.n5 VP.n0 0.285035
R17 VP.n9 VP.n0 0.285035
R18 VP VP.n9 0.0516364
R19 VTAIL.n7 VTAIL.t0 53.8717
R20 VTAIL.n11 VTAIL.t4 53.8716
R21 VTAIL.n2 VTAIL.t10 53.8716
R22 VTAIL.n10 VTAIL.t11 53.8716
R23 VTAIL.n9 VTAIL.n8 51.7935
R24 VTAIL.n6 VTAIL.n5 51.7935
R25 VTAIL.n1 VTAIL.n0 51.7932
R26 VTAIL.n4 VTAIL.n3 51.7932
R27 VTAIL.n6 VTAIL.n4 27.2807
R28 VTAIL.n11 VTAIL.n10 26.5652
R29 VTAIL.n0 VTAIL.t1 2.07882
R30 VTAIL.n0 VTAIL.t3 2.07882
R31 VTAIL.n3 VTAIL.t8 2.07882
R32 VTAIL.n3 VTAIL.t7 2.07882
R33 VTAIL.n8 VTAIL.t9 2.07882
R34 VTAIL.n8 VTAIL.t6 2.07882
R35 VTAIL.n5 VTAIL.t5 2.07882
R36 VTAIL.n5 VTAIL.t2 2.07882
R37 VTAIL.n9 VTAIL.n7 0.828086
R38 VTAIL.n2 VTAIL.n1 0.828086
R39 VTAIL.n7 VTAIL.n6 0.716017
R40 VTAIL.n10 VTAIL.n9 0.716017
R41 VTAIL.n4 VTAIL.n2 0.716017
R42 VTAIL VTAIL.n11 0.478948
R43 VTAIL VTAIL.n1 0.237569
R44 VDD1 VDD1.t5 71.1453
R45 VDD1.n1 VDD1.t4 71.0317
R46 VDD1.n1 VDD1.n0 68.5955
R47 VDD1.n3 VDD1.n2 68.4721
R48 VDD1.n3 VDD1.n1 40.4643
R49 VDD1.n2 VDD1.t3 2.07882
R50 VDD1.n2 VDD1.t2 2.07882
R51 VDD1.n0 VDD1.t1 2.07882
R52 VDD1.n0 VDD1.t0 2.07882
R53 VDD1 VDD1.n3 0.12119
R54 B.n118 B.t9 960.256
R55 B.n124 B.t6 960.256
R56 B.n38 B.t0 960.256
R57 B.n44 B.t3 960.256
R58 B.n415 B.n72 585
R59 B.n417 B.n416 585
R60 B.n418 B.n71 585
R61 B.n420 B.n419 585
R62 B.n421 B.n70 585
R63 B.n423 B.n422 585
R64 B.n424 B.n69 585
R65 B.n426 B.n425 585
R66 B.n427 B.n68 585
R67 B.n429 B.n428 585
R68 B.n430 B.n67 585
R69 B.n432 B.n431 585
R70 B.n433 B.n66 585
R71 B.n435 B.n434 585
R72 B.n436 B.n65 585
R73 B.n438 B.n437 585
R74 B.n439 B.n64 585
R75 B.n441 B.n440 585
R76 B.n442 B.n63 585
R77 B.n444 B.n443 585
R78 B.n445 B.n62 585
R79 B.n447 B.n446 585
R80 B.n448 B.n61 585
R81 B.n450 B.n449 585
R82 B.n451 B.n60 585
R83 B.n453 B.n452 585
R84 B.n454 B.n59 585
R85 B.n456 B.n455 585
R86 B.n457 B.n58 585
R87 B.n459 B.n458 585
R88 B.n460 B.n57 585
R89 B.n462 B.n461 585
R90 B.n463 B.n56 585
R91 B.n465 B.n464 585
R92 B.n466 B.n55 585
R93 B.n468 B.n467 585
R94 B.n469 B.n54 585
R95 B.n471 B.n470 585
R96 B.n472 B.n53 585
R97 B.n474 B.n473 585
R98 B.n475 B.n52 585
R99 B.n477 B.n476 585
R100 B.n478 B.n51 585
R101 B.n480 B.n479 585
R102 B.n481 B.n50 585
R103 B.n483 B.n482 585
R104 B.n484 B.n49 585
R105 B.n486 B.n485 585
R106 B.n487 B.n48 585
R107 B.n489 B.n488 585
R108 B.n490 B.n47 585
R109 B.n492 B.n491 585
R110 B.n494 B.n493 585
R111 B.n495 B.n43 585
R112 B.n497 B.n496 585
R113 B.n498 B.n42 585
R114 B.n500 B.n499 585
R115 B.n501 B.n41 585
R116 B.n503 B.n502 585
R117 B.n504 B.n40 585
R118 B.n506 B.n505 585
R119 B.n507 B.n37 585
R120 B.n510 B.n509 585
R121 B.n511 B.n36 585
R122 B.n513 B.n512 585
R123 B.n514 B.n35 585
R124 B.n516 B.n515 585
R125 B.n517 B.n34 585
R126 B.n519 B.n518 585
R127 B.n520 B.n33 585
R128 B.n522 B.n521 585
R129 B.n523 B.n32 585
R130 B.n525 B.n524 585
R131 B.n526 B.n31 585
R132 B.n528 B.n527 585
R133 B.n529 B.n30 585
R134 B.n531 B.n530 585
R135 B.n532 B.n29 585
R136 B.n534 B.n533 585
R137 B.n535 B.n28 585
R138 B.n537 B.n536 585
R139 B.n538 B.n27 585
R140 B.n540 B.n539 585
R141 B.n541 B.n26 585
R142 B.n543 B.n542 585
R143 B.n544 B.n25 585
R144 B.n546 B.n545 585
R145 B.n547 B.n24 585
R146 B.n549 B.n548 585
R147 B.n550 B.n23 585
R148 B.n552 B.n551 585
R149 B.n553 B.n22 585
R150 B.n555 B.n554 585
R151 B.n556 B.n21 585
R152 B.n558 B.n557 585
R153 B.n559 B.n20 585
R154 B.n561 B.n560 585
R155 B.n562 B.n19 585
R156 B.n564 B.n563 585
R157 B.n565 B.n18 585
R158 B.n567 B.n566 585
R159 B.n568 B.n17 585
R160 B.n570 B.n569 585
R161 B.n571 B.n16 585
R162 B.n573 B.n572 585
R163 B.n574 B.n15 585
R164 B.n576 B.n575 585
R165 B.n577 B.n14 585
R166 B.n579 B.n578 585
R167 B.n580 B.n13 585
R168 B.n582 B.n581 585
R169 B.n583 B.n12 585
R170 B.n585 B.n584 585
R171 B.n586 B.n11 585
R172 B.n414 B.n413 585
R173 B.n412 B.n73 585
R174 B.n411 B.n410 585
R175 B.n409 B.n74 585
R176 B.n408 B.n407 585
R177 B.n406 B.n75 585
R178 B.n405 B.n404 585
R179 B.n403 B.n76 585
R180 B.n402 B.n401 585
R181 B.n400 B.n77 585
R182 B.n399 B.n398 585
R183 B.n397 B.n78 585
R184 B.n396 B.n395 585
R185 B.n394 B.n79 585
R186 B.n393 B.n392 585
R187 B.n391 B.n80 585
R188 B.n390 B.n389 585
R189 B.n388 B.n81 585
R190 B.n387 B.n386 585
R191 B.n385 B.n82 585
R192 B.n384 B.n383 585
R193 B.n382 B.n83 585
R194 B.n381 B.n380 585
R195 B.n379 B.n84 585
R196 B.n378 B.n377 585
R197 B.n376 B.n85 585
R198 B.n375 B.n374 585
R199 B.n373 B.n86 585
R200 B.n372 B.n371 585
R201 B.n370 B.n87 585
R202 B.n369 B.n368 585
R203 B.n367 B.n88 585
R204 B.n366 B.n365 585
R205 B.n364 B.n89 585
R206 B.n363 B.n362 585
R207 B.n361 B.n90 585
R208 B.n360 B.n359 585
R209 B.n187 B.n152 585
R210 B.n189 B.n188 585
R211 B.n190 B.n151 585
R212 B.n192 B.n191 585
R213 B.n193 B.n150 585
R214 B.n195 B.n194 585
R215 B.n196 B.n149 585
R216 B.n198 B.n197 585
R217 B.n199 B.n148 585
R218 B.n201 B.n200 585
R219 B.n202 B.n147 585
R220 B.n204 B.n203 585
R221 B.n205 B.n146 585
R222 B.n207 B.n206 585
R223 B.n208 B.n145 585
R224 B.n210 B.n209 585
R225 B.n211 B.n144 585
R226 B.n213 B.n212 585
R227 B.n214 B.n143 585
R228 B.n216 B.n215 585
R229 B.n217 B.n142 585
R230 B.n219 B.n218 585
R231 B.n220 B.n141 585
R232 B.n222 B.n221 585
R233 B.n223 B.n140 585
R234 B.n225 B.n224 585
R235 B.n226 B.n139 585
R236 B.n228 B.n227 585
R237 B.n229 B.n138 585
R238 B.n231 B.n230 585
R239 B.n232 B.n137 585
R240 B.n234 B.n233 585
R241 B.n235 B.n136 585
R242 B.n237 B.n236 585
R243 B.n238 B.n135 585
R244 B.n240 B.n239 585
R245 B.n241 B.n134 585
R246 B.n243 B.n242 585
R247 B.n244 B.n133 585
R248 B.n246 B.n245 585
R249 B.n247 B.n132 585
R250 B.n249 B.n248 585
R251 B.n250 B.n131 585
R252 B.n252 B.n251 585
R253 B.n253 B.n130 585
R254 B.n255 B.n254 585
R255 B.n256 B.n129 585
R256 B.n258 B.n257 585
R257 B.n259 B.n128 585
R258 B.n261 B.n260 585
R259 B.n262 B.n127 585
R260 B.n264 B.n263 585
R261 B.n266 B.n265 585
R262 B.n267 B.n123 585
R263 B.n269 B.n268 585
R264 B.n270 B.n122 585
R265 B.n272 B.n271 585
R266 B.n273 B.n121 585
R267 B.n275 B.n274 585
R268 B.n276 B.n120 585
R269 B.n278 B.n277 585
R270 B.n279 B.n117 585
R271 B.n282 B.n281 585
R272 B.n283 B.n116 585
R273 B.n285 B.n284 585
R274 B.n286 B.n115 585
R275 B.n288 B.n287 585
R276 B.n289 B.n114 585
R277 B.n291 B.n290 585
R278 B.n292 B.n113 585
R279 B.n294 B.n293 585
R280 B.n295 B.n112 585
R281 B.n297 B.n296 585
R282 B.n298 B.n111 585
R283 B.n300 B.n299 585
R284 B.n301 B.n110 585
R285 B.n303 B.n302 585
R286 B.n304 B.n109 585
R287 B.n306 B.n305 585
R288 B.n307 B.n108 585
R289 B.n309 B.n308 585
R290 B.n310 B.n107 585
R291 B.n312 B.n311 585
R292 B.n313 B.n106 585
R293 B.n315 B.n314 585
R294 B.n316 B.n105 585
R295 B.n318 B.n317 585
R296 B.n319 B.n104 585
R297 B.n321 B.n320 585
R298 B.n322 B.n103 585
R299 B.n324 B.n323 585
R300 B.n325 B.n102 585
R301 B.n327 B.n326 585
R302 B.n328 B.n101 585
R303 B.n330 B.n329 585
R304 B.n331 B.n100 585
R305 B.n333 B.n332 585
R306 B.n334 B.n99 585
R307 B.n336 B.n335 585
R308 B.n337 B.n98 585
R309 B.n339 B.n338 585
R310 B.n340 B.n97 585
R311 B.n342 B.n341 585
R312 B.n343 B.n96 585
R313 B.n345 B.n344 585
R314 B.n346 B.n95 585
R315 B.n348 B.n347 585
R316 B.n349 B.n94 585
R317 B.n351 B.n350 585
R318 B.n352 B.n93 585
R319 B.n354 B.n353 585
R320 B.n355 B.n92 585
R321 B.n357 B.n356 585
R322 B.n358 B.n91 585
R323 B.n186 B.n185 585
R324 B.n184 B.n153 585
R325 B.n183 B.n182 585
R326 B.n181 B.n154 585
R327 B.n180 B.n179 585
R328 B.n178 B.n155 585
R329 B.n177 B.n176 585
R330 B.n175 B.n156 585
R331 B.n174 B.n173 585
R332 B.n172 B.n157 585
R333 B.n171 B.n170 585
R334 B.n169 B.n158 585
R335 B.n168 B.n167 585
R336 B.n166 B.n159 585
R337 B.n165 B.n164 585
R338 B.n163 B.n160 585
R339 B.n162 B.n161 585
R340 B.n2 B.n0 585
R341 B.n613 B.n1 585
R342 B.n612 B.n611 585
R343 B.n610 B.n3 585
R344 B.n609 B.n608 585
R345 B.n607 B.n4 585
R346 B.n606 B.n605 585
R347 B.n604 B.n5 585
R348 B.n603 B.n602 585
R349 B.n601 B.n6 585
R350 B.n600 B.n599 585
R351 B.n598 B.n7 585
R352 B.n597 B.n596 585
R353 B.n595 B.n8 585
R354 B.n594 B.n593 585
R355 B.n592 B.n9 585
R356 B.n591 B.n590 585
R357 B.n589 B.n10 585
R358 B.n588 B.n587 585
R359 B.n615 B.n614 585
R360 B.n187 B.n186 497.305
R361 B.n588 B.n11 497.305
R362 B.n360 B.n91 497.305
R363 B.n415 B.n414 497.305
R364 B.n186 B.n153 163.367
R365 B.n182 B.n153 163.367
R366 B.n182 B.n181 163.367
R367 B.n181 B.n180 163.367
R368 B.n180 B.n155 163.367
R369 B.n176 B.n155 163.367
R370 B.n176 B.n175 163.367
R371 B.n175 B.n174 163.367
R372 B.n174 B.n157 163.367
R373 B.n170 B.n157 163.367
R374 B.n170 B.n169 163.367
R375 B.n169 B.n168 163.367
R376 B.n168 B.n159 163.367
R377 B.n164 B.n159 163.367
R378 B.n164 B.n163 163.367
R379 B.n163 B.n162 163.367
R380 B.n162 B.n2 163.367
R381 B.n614 B.n2 163.367
R382 B.n614 B.n613 163.367
R383 B.n613 B.n612 163.367
R384 B.n612 B.n3 163.367
R385 B.n608 B.n3 163.367
R386 B.n608 B.n607 163.367
R387 B.n607 B.n606 163.367
R388 B.n606 B.n5 163.367
R389 B.n602 B.n5 163.367
R390 B.n602 B.n601 163.367
R391 B.n601 B.n600 163.367
R392 B.n600 B.n7 163.367
R393 B.n596 B.n7 163.367
R394 B.n596 B.n595 163.367
R395 B.n595 B.n594 163.367
R396 B.n594 B.n9 163.367
R397 B.n590 B.n9 163.367
R398 B.n590 B.n589 163.367
R399 B.n589 B.n588 163.367
R400 B.n188 B.n187 163.367
R401 B.n188 B.n151 163.367
R402 B.n192 B.n151 163.367
R403 B.n193 B.n192 163.367
R404 B.n194 B.n193 163.367
R405 B.n194 B.n149 163.367
R406 B.n198 B.n149 163.367
R407 B.n199 B.n198 163.367
R408 B.n200 B.n199 163.367
R409 B.n200 B.n147 163.367
R410 B.n204 B.n147 163.367
R411 B.n205 B.n204 163.367
R412 B.n206 B.n205 163.367
R413 B.n206 B.n145 163.367
R414 B.n210 B.n145 163.367
R415 B.n211 B.n210 163.367
R416 B.n212 B.n211 163.367
R417 B.n212 B.n143 163.367
R418 B.n216 B.n143 163.367
R419 B.n217 B.n216 163.367
R420 B.n218 B.n217 163.367
R421 B.n218 B.n141 163.367
R422 B.n222 B.n141 163.367
R423 B.n223 B.n222 163.367
R424 B.n224 B.n223 163.367
R425 B.n224 B.n139 163.367
R426 B.n228 B.n139 163.367
R427 B.n229 B.n228 163.367
R428 B.n230 B.n229 163.367
R429 B.n230 B.n137 163.367
R430 B.n234 B.n137 163.367
R431 B.n235 B.n234 163.367
R432 B.n236 B.n235 163.367
R433 B.n236 B.n135 163.367
R434 B.n240 B.n135 163.367
R435 B.n241 B.n240 163.367
R436 B.n242 B.n241 163.367
R437 B.n242 B.n133 163.367
R438 B.n246 B.n133 163.367
R439 B.n247 B.n246 163.367
R440 B.n248 B.n247 163.367
R441 B.n248 B.n131 163.367
R442 B.n252 B.n131 163.367
R443 B.n253 B.n252 163.367
R444 B.n254 B.n253 163.367
R445 B.n254 B.n129 163.367
R446 B.n258 B.n129 163.367
R447 B.n259 B.n258 163.367
R448 B.n260 B.n259 163.367
R449 B.n260 B.n127 163.367
R450 B.n264 B.n127 163.367
R451 B.n265 B.n264 163.367
R452 B.n265 B.n123 163.367
R453 B.n269 B.n123 163.367
R454 B.n270 B.n269 163.367
R455 B.n271 B.n270 163.367
R456 B.n271 B.n121 163.367
R457 B.n275 B.n121 163.367
R458 B.n276 B.n275 163.367
R459 B.n277 B.n276 163.367
R460 B.n277 B.n117 163.367
R461 B.n282 B.n117 163.367
R462 B.n283 B.n282 163.367
R463 B.n284 B.n283 163.367
R464 B.n284 B.n115 163.367
R465 B.n288 B.n115 163.367
R466 B.n289 B.n288 163.367
R467 B.n290 B.n289 163.367
R468 B.n290 B.n113 163.367
R469 B.n294 B.n113 163.367
R470 B.n295 B.n294 163.367
R471 B.n296 B.n295 163.367
R472 B.n296 B.n111 163.367
R473 B.n300 B.n111 163.367
R474 B.n301 B.n300 163.367
R475 B.n302 B.n301 163.367
R476 B.n302 B.n109 163.367
R477 B.n306 B.n109 163.367
R478 B.n307 B.n306 163.367
R479 B.n308 B.n307 163.367
R480 B.n308 B.n107 163.367
R481 B.n312 B.n107 163.367
R482 B.n313 B.n312 163.367
R483 B.n314 B.n313 163.367
R484 B.n314 B.n105 163.367
R485 B.n318 B.n105 163.367
R486 B.n319 B.n318 163.367
R487 B.n320 B.n319 163.367
R488 B.n320 B.n103 163.367
R489 B.n324 B.n103 163.367
R490 B.n325 B.n324 163.367
R491 B.n326 B.n325 163.367
R492 B.n326 B.n101 163.367
R493 B.n330 B.n101 163.367
R494 B.n331 B.n330 163.367
R495 B.n332 B.n331 163.367
R496 B.n332 B.n99 163.367
R497 B.n336 B.n99 163.367
R498 B.n337 B.n336 163.367
R499 B.n338 B.n337 163.367
R500 B.n338 B.n97 163.367
R501 B.n342 B.n97 163.367
R502 B.n343 B.n342 163.367
R503 B.n344 B.n343 163.367
R504 B.n344 B.n95 163.367
R505 B.n348 B.n95 163.367
R506 B.n349 B.n348 163.367
R507 B.n350 B.n349 163.367
R508 B.n350 B.n93 163.367
R509 B.n354 B.n93 163.367
R510 B.n355 B.n354 163.367
R511 B.n356 B.n355 163.367
R512 B.n356 B.n91 163.367
R513 B.n361 B.n360 163.367
R514 B.n362 B.n361 163.367
R515 B.n362 B.n89 163.367
R516 B.n366 B.n89 163.367
R517 B.n367 B.n366 163.367
R518 B.n368 B.n367 163.367
R519 B.n368 B.n87 163.367
R520 B.n372 B.n87 163.367
R521 B.n373 B.n372 163.367
R522 B.n374 B.n373 163.367
R523 B.n374 B.n85 163.367
R524 B.n378 B.n85 163.367
R525 B.n379 B.n378 163.367
R526 B.n380 B.n379 163.367
R527 B.n380 B.n83 163.367
R528 B.n384 B.n83 163.367
R529 B.n385 B.n384 163.367
R530 B.n386 B.n385 163.367
R531 B.n386 B.n81 163.367
R532 B.n390 B.n81 163.367
R533 B.n391 B.n390 163.367
R534 B.n392 B.n391 163.367
R535 B.n392 B.n79 163.367
R536 B.n396 B.n79 163.367
R537 B.n397 B.n396 163.367
R538 B.n398 B.n397 163.367
R539 B.n398 B.n77 163.367
R540 B.n402 B.n77 163.367
R541 B.n403 B.n402 163.367
R542 B.n404 B.n403 163.367
R543 B.n404 B.n75 163.367
R544 B.n408 B.n75 163.367
R545 B.n409 B.n408 163.367
R546 B.n410 B.n409 163.367
R547 B.n410 B.n73 163.367
R548 B.n414 B.n73 163.367
R549 B.n584 B.n11 163.367
R550 B.n584 B.n583 163.367
R551 B.n583 B.n582 163.367
R552 B.n582 B.n13 163.367
R553 B.n578 B.n13 163.367
R554 B.n578 B.n577 163.367
R555 B.n577 B.n576 163.367
R556 B.n576 B.n15 163.367
R557 B.n572 B.n15 163.367
R558 B.n572 B.n571 163.367
R559 B.n571 B.n570 163.367
R560 B.n570 B.n17 163.367
R561 B.n566 B.n17 163.367
R562 B.n566 B.n565 163.367
R563 B.n565 B.n564 163.367
R564 B.n564 B.n19 163.367
R565 B.n560 B.n19 163.367
R566 B.n560 B.n559 163.367
R567 B.n559 B.n558 163.367
R568 B.n558 B.n21 163.367
R569 B.n554 B.n21 163.367
R570 B.n554 B.n553 163.367
R571 B.n553 B.n552 163.367
R572 B.n552 B.n23 163.367
R573 B.n548 B.n23 163.367
R574 B.n548 B.n547 163.367
R575 B.n547 B.n546 163.367
R576 B.n546 B.n25 163.367
R577 B.n542 B.n25 163.367
R578 B.n542 B.n541 163.367
R579 B.n541 B.n540 163.367
R580 B.n540 B.n27 163.367
R581 B.n536 B.n27 163.367
R582 B.n536 B.n535 163.367
R583 B.n535 B.n534 163.367
R584 B.n534 B.n29 163.367
R585 B.n530 B.n29 163.367
R586 B.n530 B.n529 163.367
R587 B.n529 B.n528 163.367
R588 B.n528 B.n31 163.367
R589 B.n524 B.n31 163.367
R590 B.n524 B.n523 163.367
R591 B.n523 B.n522 163.367
R592 B.n522 B.n33 163.367
R593 B.n518 B.n33 163.367
R594 B.n518 B.n517 163.367
R595 B.n517 B.n516 163.367
R596 B.n516 B.n35 163.367
R597 B.n512 B.n35 163.367
R598 B.n512 B.n511 163.367
R599 B.n511 B.n510 163.367
R600 B.n510 B.n37 163.367
R601 B.n505 B.n37 163.367
R602 B.n505 B.n504 163.367
R603 B.n504 B.n503 163.367
R604 B.n503 B.n41 163.367
R605 B.n499 B.n41 163.367
R606 B.n499 B.n498 163.367
R607 B.n498 B.n497 163.367
R608 B.n497 B.n43 163.367
R609 B.n493 B.n43 163.367
R610 B.n493 B.n492 163.367
R611 B.n492 B.n47 163.367
R612 B.n488 B.n47 163.367
R613 B.n488 B.n487 163.367
R614 B.n487 B.n486 163.367
R615 B.n486 B.n49 163.367
R616 B.n482 B.n49 163.367
R617 B.n482 B.n481 163.367
R618 B.n481 B.n480 163.367
R619 B.n480 B.n51 163.367
R620 B.n476 B.n51 163.367
R621 B.n476 B.n475 163.367
R622 B.n475 B.n474 163.367
R623 B.n474 B.n53 163.367
R624 B.n470 B.n53 163.367
R625 B.n470 B.n469 163.367
R626 B.n469 B.n468 163.367
R627 B.n468 B.n55 163.367
R628 B.n464 B.n55 163.367
R629 B.n464 B.n463 163.367
R630 B.n463 B.n462 163.367
R631 B.n462 B.n57 163.367
R632 B.n458 B.n57 163.367
R633 B.n458 B.n457 163.367
R634 B.n457 B.n456 163.367
R635 B.n456 B.n59 163.367
R636 B.n452 B.n59 163.367
R637 B.n452 B.n451 163.367
R638 B.n451 B.n450 163.367
R639 B.n450 B.n61 163.367
R640 B.n446 B.n61 163.367
R641 B.n446 B.n445 163.367
R642 B.n445 B.n444 163.367
R643 B.n444 B.n63 163.367
R644 B.n440 B.n63 163.367
R645 B.n440 B.n439 163.367
R646 B.n439 B.n438 163.367
R647 B.n438 B.n65 163.367
R648 B.n434 B.n65 163.367
R649 B.n434 B.n433 163.367
R650 B.n433 B.n432 163.367
R651 B.n432 B.n67 163.367
R652 B.n428 B.n67 163.367
R653 B.n428 B.n427 163.367
R654 B.n427 B.n426 163.367
R655 B.n426 B.n69 163.367
R656 B.n422 B.n69 163.367
R657 B.n422 B.n421 163.367
R658 B.n421 B.n420 163.367
R659 B.n420 B.n71 163.367
R660 B.n416 B.n71 163.367
R661 B.n416 B.n415 163.367
R662 B.n118 B.t11 122.57
R663 B.n44 B.t4 122.57
R664 B.n124 B.t8 122.55
R665 B.n38 B.t1 122.55
R666 B.n119 B.t10 106.474
R667 B.n45 B.t5 106.474
R668 B.n125 B.t7 106.454
R669 B.n39 B.t2 106.454
R670 B.n280 B.n119 59.5399
R671 B.n126 B.n125 59.5399
R672 B.n508 B.n39 59.5399
R673 B.n46 B.n45 59.5399
R674 B.n587 B.n586 32.3127
R675 B.n413 B.n72 32.3127
R676 B.n359 B.n358 32.3127
R677 B.n185 B.n152 32.3127
R678 B B.n615 18.0485
R679 B.n119 B.n118 16.0975
R680 B.n125 B.n124 16.0975
R681 B.n39 B.n38 16.0975
R682 B.n45 B.n44 16.0975
R683 B.n586 B.n585 10.6151
R684 B.n585 B.n12 10.6151
R685 B.n581 B.n12 10.6151
R686 B.n581 B.n580 10.6151
R687 B.n580 B.n579 10.6151
R688 B.n579 B.n14 10.6151
R689 B.n575 B.n14 10.6151
R690 B.n575 B.n574 10.6151
R691 B.n574 B.n573 10.6151
R692 B.n573 B.n16 10.6151
R693 B.n569 B.n16 10.6151
R694 B.n569 B.n568 10.6151
R695 B.n568 B.n567 10.6151
R696 B.n567 B.n18 10.6151
R697 B.n563 B.n18 10.6151
R698 B.n563 B.n562 10.6151
R699 B.n562 B.n561 10.6151
R700 B.n561 B.n20 10.6151
R701 B.n557 B.n20 10.6151
R702 B.n557 B.n556 10.6151
R703 B.n556 B.n555 10.6151
R704 B.n555 B.n22 10.6151
R705 B.n551 B.n22 10.6151
R706 B.n551 B.n550 10.6151
R707 B.n550 B.n549 10.6151
R708 B.n549 B.n24 10.6151
R709 B.n545 B.n24 10.6151
R710 B.n545 B.n544 10.6151
R711 B.n544 B.n543 10.6151
R712 B.n543 B.n26 10.6151
R713 B.n539 B.n26 10.6151
R714 B.n539 B.n538 10.6151
R715 B.n538 B.n537 10.6151
R716 B.n537 B.n28 10.6151
R717 B.n533 B.n28 10.6151
R718 B.n533 B.n532 10.6151
R719 B.n532 B.n531 10.6151
R720 B.n531 B.n30 10.6151
R721 B.n527 B.n30 10.6151
R722 B.n527 B.n526 10.6151
R723 B.n526 B.n525 10.6151
R724 B.n525 B.n32 10.6151
R725 B.n521 B.n32 10.6151
R726 B.n521 B.n520 10.6151
R727 B.n520 B.n519 10.6151
R728 B.n519 B.n34 10.6151
R729 B.n515 B.n34 10.6151
R730 B.n515 B.n514 10.6151
R731 B.n514 B.n513 10.6151
R732 B.n513 B.n36 10.6151
R733 B.n509 B.n36 10.6151
R734 B.n507 B.n506 10.6151
R735 B.n506 B.n40 10.6151
R736 B.n502 B.n40 10.6151
R737 B.n502 B.n501 10.6151
R738 B.n501 B.n500 10.6151
R739 B.n500 B.n42 10.6151
R740 B.n496 B.n42 10.6151
R741 B.n496 B.n495 10.6151
R742 B.n495 B.n494 10.6151
R743 B.n491 B.n490 10.6151
R744 B.n490 B.n489 10.6151
R745 B.n489 B.n48 10.6151
R746 B.n485 B.n48 10.6151
R747 B.n485 B.n484 10.6151
R748 B.n484 B.n483 10.6151
R749 B.n483 B.n50 10.6151
R750 B.n479 B.n50 10.6151
R751 B.n479 B.n478 10.6151
R752 B.n478 B.n477 10.6151
R753 B.n477 B.n52 10.6151
R754 B.n473 B.n52 10.6151
R755 B.n473 B.n472 10.6151
R756 B.n472 B.n471 10.6151
R757 B.n471 B.n54 10.6151
R758 B.n467 B.n54 10.6151
R759 B.n467 B.n466 10.6151
R760 B.n466 B.n465 10.6151
R761 B.n465 B.n56 10.6151
R762 B.n461 B.n56 10.6151
R763 B.n461 B.n460 10.6151
R764 B.n460 B.n459 10.6151
R765 B.n459 B.n58 10.6151
R766 B.n455 B.n58 10.6151
R767 B.n455 B.n454 10.6151
R768 B.n454 B.n453 10.6151
R769 B.n453 B.n60 10.6151
R770 B.n449 B.n60 10.6151
R771 B.n449 B.n448 10.6151
R772 B.n448 B.n447 10.6151
R773 B.n447 B.n62 10.6151
R774 B.n443 B.n62 10.6151
R775 B.n443 B.n442 10.6151
R776 B.n442 B.n441 10.6151
R777 B.n441 B.n64 10.6151
R778 B.n437 B.n64 10.6151
R779 B.n437 B.n436 10.6151
R780 B.n436 B.n435 10.6151
R781 B.n435 B.n66 10.6151
R782 B.n431 B.n66 10.6151
R783 B.n431 B.n430 10.6151
R784 B.n430 B.n429 10.6151
R785 B.n429 B.n68 10.6151
R786 B.n425 B.n68 10.6151
R787 B.n425 B.n424 10.6151
R788 B.n424 B.n423 10.6151
R789 B.n423 B.n70 10.6151
R790 B.n419 B.n70 10.6151
R791 B.n419 B.n418 10.6151
R792 B.n418 B.n417 10.6151
R793 B.n417 B.n72 10.6151
R794 B.n359 B.n90 10.6151
R795 B.n363 B.n90 10.6151
R796 B.n364 B.n363 10.6151
R797 B.n365 B.n364 10.6151
R798 B.n365 B.n88 10.6151
R799 B.n369 B.n88 10.6151
R800 B.n370 B.n369 10.6151
R801 B.n371 B.n370 10.6151
R802 B.n371 B.n86 10.6151
R803 B.n375 B.n86 10.6151
R804 B.n376 B.n375 10.6151
R805 B.n377 B.n376 10.6151
R806 B.n377 B.n84 10.6151
R807 B.n381 B.n84 10.6151
R808 B.n382 B.n381 10.6151
R809 B.n383 B.n382 10.6151
R810 B.n383 B.n82 10.6151
R811 B.n387 B.n82 10.6151
R812 B.n388 B.n387 10.6151
R813 B.n389 B.n388 10.6151
R814 B.n389 B.n80 10.6151
R815 B.n393 B.n80 10.6151
R816 B.n394 B.n393 10.6151
R817 B.n395 B.n394 10.6151
R818 B.n395 B.n78 10.6151
R819 B.n399 B.n78 10.6151
R820 B.n400 B.n399 10.6151
R821 B.n401 B.n400 10.6151
R822 B.n401 B.n76 10.6151
R823 B.n405 B.n76 10.6151
R824 B.n406 B.n405 10.6151
R825 B.n407 B.n406 10.6151
R826 B.n407 B.n74 10.6151
R827 B.n411 B.n74 10.6151
R828 B.n412 B.n411 10.6151
R829 B.n413 B.n412 10.6151
R830 B.n189 B.n152 10.6151
R831 B.n190 B.n189 10.6151
R832 B.n191 B.n190 10.6151
R833 B.n191 B.n150 10.6151
R834 B.n195 B.n150 10.6151
R835 B.n196 B.n195 10.6151
R836 B.n197 B.n196 10.6151
R837 B.n197 B.n148 10.6151
R838 B.n201 B.n148 10.6151
R839 B.n202 B.n201 10.6151
R840 B.n203 B.n202 10.6151
R841 B.n203 B.n146 10.6151
R842 B.n207 B.n146 10.6151
R843 B.n208 B.n207 10.6151
R844 B.n209 B.n208 10.6151
R845 B.n209 B.n144 10.6151
R846 B.n213 B.n144 10.6151
R847 B.n214 B.n213 10.6151
R848 B.n215 B.n214 10.6151
R849 B.n215 B.n142 10.6151
R850 B.n219 B.n142 10.6151
R851 B.n220 B.n219 10.6151
R852 B.n221 B.n220 10.6151
R853 B.n221 B.n140 10.6151
R854 B.n225 B.n140 10.6151
R855 B.n226 B.n225 10.6151
R856 B.n227 B.n226 10.6151
R857 B.n227 B.n138 10.6151
R858 B.n231 B.n138 10.6151
R859 B.n232 B.n231 10.6151
R860 B.n233 B.n232 10.6151
R861 B.n233 B.n136 10.6151
R862 B.n237 B.n136 10.6151
R863 B.n238 B.n237 10.6151
R864 B.n239 B.n238 10.6151
R865 B.n239 B.n134 10.6151
R866 B.n243 B.n134 10.6151
R867 B.n244 B.n243 10.6151
R868 B.n245 B.n244 10.6151
R869 B.n245 B.n132 10.6151
R870 B.n249 B.n132 10.6151
R871 B.n250 B.n249 10.6151
R872 B.n251 B.n250 10.6151
R873 B.n251 B.n130 10.6151
R874 B.n255 B.n130 10.6151
R875 B.n256 B.n255 10.6151
R876 B.n257 B.n256 10.6151
R877 B.n257 B.n128 10.6151
R878 B.n261 B.n128 10.6151
R879 B.n262 B.n261 10.6151
R880 B.n263 B.n262 10.6151
R881 B.n267 B.n266 10.6151
R882 B.n268 B.n267 10.6151
R883 B.n268 B.n122 10.6151
R884 B.n272 B.n122 10.6151
R885 B.n273 B.n272 10.6151
R886 B.n274 B.n273 10.6151
R887 B.n274 B.n120 10.6151
R888 B.n278 B.n120 10.6151
R889 B.n279 B.n278 10.6151
R890 B.n281 B.n116 10.6151
R891 B.n285 B.n116 10.6151
R892 B.n286 B.n285 10.6151
R893 B.n287 B.n286 10.6151
R894 B.n287 B.n114 10.6151
R895 B.n291 B.n114 10.6151
R896 B.n292 B.n291 10.6151
R897 B.n293 B.n292 10.6151
R898 B.n293 B.n112 10.6151
R899 B.n297 B.n112 10.6151
R900 B.n298 B.n297 10.6151
R901 B.n299 B.n298 10.6151
R902 B.n299 B.n110 10.6151
R903 B.n303 B.n110 10.6151
R904 B.n304 B.n303 10.6151
R905 B.n305 B.n304 10.6151
R906 B.n305 B.n108 10.6151
R907 B.n309 B.n108 10.6151
R908 B.n310 B.n309 10.6151
R909 B.n311 B.n310 10.6151
R910 B.n311 B.n106 10.6151
R911 B.n315 B.n106 10.6151
R912 B.n316 B.n315 10.6151
R913 B.n317 B.n316 10.6151
R914 B.n317 B.n104 10.6151
R915 B.n321 B.n104 10.6151
R916 B.n322 B.n321 10.6151
R917 B.n323 B.n322 10.6151
R918 B.n323 B.n102 10.6151
R919 B.n327 B.n102 10.6151
R920 B.n328 B.n327 10.6151
R921 B.n329 B.n328 10.6151
R922 B.n329 B.n100 10.6151
R923 B.n333 B.n100 10.6151
R924 B.n334 B.n333 10.6151
R925 B.n335 B.n334 10.6151
R926 B.n335 B.n98 10.6151
R927 B.n339 B.n98 10.6151
R928 B.n340 B.n339 10.6151
R929 B.n341 B.n340 10.6151
R930 B.n341 B.n96 10.6151
R931 B.n345 B.n96 10.6151
R932 B.n346 B.n345 10.6151
R933 B.n347 B.n346 10.6151
R934 B.n347 B.n94 10.6151
R935 B.n351 B.n94 10.6151
R936 B.n352 B.n351 10.6151
R937 B.n353 B.n352 10.6151
R938 B.n353 B.n92 10.6151
R939 B.n357 B.n92 10.6151
R940 B.n358 B.n357 10.6151
R941 B.n185 B.n184 10.6151
R942 B.n184 B.n183 10.6151
R943 B.n183 B.n154 10.6151
R944 B.n179 B.n154 10.6151
R945 B.n179 B.n178 10.6151
R946 B.n178 B.n177 10.6151
R947 B.n177 B.n156 10.6151
R948 B.n173 B.n156 10.6151
R949 B.n173 B.n172 10.6151
R950 B.n172 B.n171 10.6151
R951 B.n171 B.n158 10.6151
R952 B.n167 B.n158 10.6151
R953 B.n167 B.n166 10.6151
R954 B.n166 B.n165 10.6151
R955 B.n165 B.n160 10.6151
R956 B.n161 B.n160 10.6151
R957 B.n161 B.n0 10.6151
R958 B.n611 B.n1 10.6151
R959 B.n611 B.n610 10.6151
R960 B.n610 B.n609 10.6151
R961 B.n609 B.n4 10.6151
R962 B.n605 B.n4 10.6151
R963 B.n605 B.n604 10.6151
R964 B.n604 B.n603 10.6151
R965 B.n603 B.n6 10.6151
R966 B.n599 B.n6 10.6151
R967 B.n599 B.n598 10.6151
R968 B.n598 B.n597 10.6151
R969 B.n597 B.n8 10.6151
R970 B.n593 B.n8 10.6151
R971 B.n593 B.n592 10.6151
R972 B.n592 B.n591 10.6151
R973 B.n591 B.n10 10.6151
R974 B.n587 B.n10 10.6151
R975 B.n509 B.n508 9.36635
R976 B.n491 B.n46 9.36635
R977 B.n263 B.n126 9.36635
R978 B.n281 B.n280 9.36635
R979 B.n615 B.n0 2.81026
R980 B.n615 B.n1 2.81026
R981 B.n508 B.n507 1.24928
R982 B.n494 B.n46 1.24928
R983 B.n266 B.n126 1.24928
R984 B.n280 B.n279 1.24928
R985 VN.n0 VN.t5 859.236
R986 VN.n4 VN.t2 859.236
R987 VN.n1 VN.t4 832.414
R988 VN.n2 VN.t1 832.414
R989 VN.n5 VN.t3 832.414
R990 VN.n6 VN.t0 832.414
R991 VN.n3 VN.n2 161.3
R992 VN.n7 VN.n6 161.3
R993 VN.n2 VN.n1 48.2005
R994 VN.n6 VN.n5 48.2005
R995 VN.n7 VN.n4 45.1367
R996 VN.n3 VN.n0 45.1367
R997 VN VN.n7 43.5441
R998 VN.n5 VN.n4 13.3799
R999 VN.n1 VN.n0 13.3799
R1000 VN VN.n3 0.0516364
R1001 VDD2.n1 VDD2.t0 71.0317
R1002 VDD2.n2 VDD2.t5 70.5505
R1003 VDD2.n1 VDD2.n0 68.5955
R1004 VDD2 VDD2.n3 68.5928
R1005 VDD2.n2 VDD2.n1 39.5235
R1006 VDD2.n3 VDD2.t2 2.07882
R1007 VDD2.n3 VDD2.t3 2.07882
R1008 VDD2.n0 VDD2.t1 2.07882
R1009 VDD2.n0 VDD2.t4 2.07882
R1010 VDD2 VDD2.n2 0.595328
C0 VP VDD2 0.281755f
C1 w_n1634_n4096# VDD1 2.02709f
C2 VTAIL VDD1 14.236402f
C3 VP VN 5.56067f
C4 B VP 1.09793f
C5 VN VDD2 4.64116f
C6 B VDD2 1.78181f
C7 w_n1634_n4096# VP 2.86332f
C8 VP VTAIL 4.12798f
C9 w_n1634_n4096# VDD2 2.04506f
C10 VDD2 VTAIL 14.266f
C11 B VN 0.765562f
C12 VP VDD1 4.76847f
C13 w_n1634_n4096# VN 2.65792f
C14 VN VTAIL 4.11313f
C15 B w_n1634_n4096# 7.79936f
C16 VDD2 VDD1 0.641079f
C17 B VTAIL 3.19158f
C18 w_n1634_n4096# VTAIL 3.54563f
C19 VN VDD1 0.148247f
C20 B VDD1 1.75748f
C21 VDD2 VSUBS 1.515858f
C22 VDD1 VSUBS 1.798659f
C23 VTAIL VSUBS 0.774262f
C24 VN VSUBS 4.74198f
C25 VP VSUBS 1.449627f
C26 B VSUBS 2.853954f
C27 w_n1634_n4096# VSUBS 82.020294f
C28 VDD2.t0 VSUBS 3.58857f
C29 VDD2.t1 VSUBS 0.338979f
C30 VDD2.t4 VSUBS 0.338979f
C31 VDD2.n0 VSUBS 2.75904f
C32 VDD2.n1 VSUBS 3.08258f
C33 VDD2.t5 VSUBS 3.58392f
C34 VDD2.n2 VSUBS 3.08657f
C35 VDD2.t2 VSUBS 0.338979f
C36 VDD2.t3 VSUBS 0.338979f
C37 VDD2.n3 VSUBS 2.75899f
C38 VN.t5 VSUBS 1.36416f
C39 VN.n0 VSUBS 0.506927f
C40 VN.t4 VSUBS 1.34786f
C41 VN.n1 VSUBS 0.535788f
C42 VN.t1 VSUBS 1.34786f
C43 VN.n2 VSUBS 0.522016f
C44 VN.n3 VSUBS 0.233872f
C45 VN.t2 VSUBS 1.36416f
C46 VN.n4 VSUBS 0.506927f
C47 VN.t3 VSUBS 1.34786f
C48 VN.n5 VSUBS 0.535788f
C49 VN.t0 VSUBS 1.34786f
C50 VN.n6 VSUBS 0.522016f
C51 VN.n7 VSUBS 2.84718f
C52 B.n0 VSUBS 0.004548f
C53 B.n1 VSUBS 0.004548f
C54 B.n2 VSUBS 0.007192f
C55 B.n3 VSUBS 0.007192f
C56 B.n4 VSUBS 0.007192f
C57 B.n5 VSUBS 0.007192f
C58 B.n6 VSUBS 0.007192f
C59 B.n7 VSUBS 0.007192f
C60 B.n8 VSUBS 0.007192f
C61 B.n9 VSUBS 0.007192f
C62 B.n10 VSUBS 0.007192f
C63 B.n11 VSUBS 0.016952f
C64 B.n12 VSUBS 0.007192f
C65 B.n13 VSUBS 0.007192f
C66 B.n14 VSUBS 0.007192f
C67 B.n15 VSUBS 0.007192f
C68 B.n16 VSUBS 0.007192f
C69 B.n17 VSUBS 0.007192f
C70 B.n18 VSUBS 0.007192f
C71 B.n19 VSUBS 0.007192f
C72 B.n20 VSUBS 0.007192f
C73 B.n21 VSUBS 0.007192f
C74 B.n22 VSUBS 0.007192f
C75 B.n23 VSUBS 0.007192f
C76 B.n24 VSUBS 0.007192f
C77 B.n25 VSUBS 0.007192f
C78 B.n26 VSUBS 0.007192f
C79 B.n27 VSUBS 0.007192f
C80 B.n28 VSUBS 0.007192f
C81 B.n29 VSUBS 0.007192f
C82 B.n30 VSUBS 0.007192f
C83 B.n31 VSUBS 0.007192f
C84 B.n32 VSUBS 0.007192f
C85 B.n33 VSUBS 0.007192f
C86 B.n34 VSUBS 0.007192f
C87 B.n35 VSUBS 0.007192f
C88 B.n36 VSUBS 0.007192f
C89 B.n37 VSUBS 0.007192f
C90 B.t2 VSUBS 0.536754f
C91 B.t1 VSUBS 0.543957f
C92 B.t0 VSUBS 0.320063f
C93 B.n38 VSUBS 0.143725f
C94 B.n39 VSUBS 0.065099f
C95 B.n40 VSUBS 0.007192f
C96 B.n41 VSUBS 0.007192f
C97 B.n42 VSUBS 0.007192f
C98 B.n43 VSUBS 0.007192f
C99 B.t5 VSUBS 0.536737f
C100 B.t4 VSUBS 0.543941f
C101 B.t3 VSUBS 0.320063f
C102 B.n44 VSUBS 0.14374f
C103 B.n45 VSUBS 0.065115f
C104 B.n46 VSUBS 0.016664f
C105 B.n47 VSUBS 0.007192f
C106 B.n48 VSUBS 0.007192f
C107 B.n49 VSUBS 0.007192f
C108 B.n50 VSUBS 0.007192f
C109 B.n51 VSUBS 0.007192f
C110 B.n52 VSUBS 0.007192f
C111 B.n53 VSUBS 0.007192f
C112 B.n54 VSUBS 0.007192f
C113 B.n55 VSUBS 0.007192f
C114 B.n56 VSUBS 0.007192f
C115 B.n57 VSUBS 0.007192f
C116 B.n58 VSUBS 0.007192f
C117 B.n59 VSUBS 0.007192f
C118 B.n60 VSUBS 0.007192f
C119 B.n61 VSUBS 0.007192f
C120 B.n62 VSUBS 0.007192f
C121 B.n63 VSUBS 0.007192f
C122 B.n64 VSUBS 0.007192f
C123 B.n65 VSUBS 0.007192f
C124 B.n66 VSUBS 0.007192f
C125 B.n67 VSUBS 0.007192f
C126 B.n68 VSUBS 0.007192f
C127 B.n69 VSUBS 0.007192f
C128 B.n70 VSUBS 0.007192f
C129 B.n71 VSUBS 0.007192f
C130 B.n72 VSUBS 0.016093f
C131 B.n73 VSUBS 0.007192f
C132 B.n74 VSUBS 0.007192f
C133 B.n75 VSUBS 0.007192f
C134 B.n76 VSUBS 0.007192f
C135 B.n77 VSUBS 0.007192f
C136 B.n78 VSUBS 0.007192f
C137 B.n79 VSUBS 0.007192f
C138 B.n80 VSUBS 0.007192f
C139 B.n81 VSUBS 0.007192f
C140 B.n82 VSUBS 0.007192f
C141 B.n83 VSUBS 0.007192f
C142 B.n84 VSUBS 0.007192f
C143 B.n85 VSUBS 0.007192f
C144 B.n86 VSUBS 0.007192f
C145 B.n87 VSUBS 0.007192f
C146 B.n88 VSUBS 0.007192f
C147 B.n89 VSUBS 0.007192f
C148 B.n90 VSUBS 0.007192f
C149 B.n91 VSUBS 0.016952f
C150 B.n92 VSUBS 0.007192f
C151 B.n93 VSUBS 0.007192f
C152 B.n94 VSUBS 0.007192f
C153 B.n95 VSUBS 0.007192f
C154 B.n96 VSUBS 0.007192f
C155 B.n97 VSUBS 0.007192f
C156 B.n98 VSUBS 0.007192f
C157 B.n99 VSUBS 0.007192f
C158 B.n100 VSUBS 0.007192f
C159 B.n101 VSUBS 0.007192f
C160 B.n102 VSUBS 0.007192f
C161 B.n103 VSUBS 0.007192f
C162 B.n104 VSUBS 0.007192f
C163 B.n105 VSUBS 0.007192f
C164 B.n106 VSUBS 0.007192f
C165 B.n107 VSUBS 0.007192f
C166 B.n108 VSUBS 0.007192f
C167 B.n109 VSUBS 0.007192f
C168 B.n110 VSUBS 0.007192f
C169 B.n111 VSUBS 0.007192f
C170 B.n112 VSUBS 0.007192f
C171 B.n113 VSUBS 0.007192f
C172 B.n114 VSUBS 0.007192f
C173 B.n115 VSUBS 0.007192f
C174 B.n116 VSUBS 0.007192f
C175 B.n117 VSUBS 0.007192f
C176 B.t10 VSUBS 0.536737f
C177 B.t11 VSUBS 0.543941f
C178 B.t9 VSUBS 0.320063f
C179 B.n118 VSUBS 0.14374f
C180 B.n119 VSUBS 0.065115f
C181 B.n120 VSUBS 0.007192f
C182 B.n121 VSUBS 0.007192f
C183 B.n122 VSUBS 0.007192f
C184 B.n123 VSUBS 0.007192f
C185 B.t7 VSUBS 0.536754f
C186 B.t8 VSUBS 0.543957f
C187 B.t6 VSUBS 0.320063f
C188 B.n124 VSUBS 0.143725f
C189 B.n125 VSUBS 0.065099f
C190 B.n126 VSUBS 0.016664f
C191 B.n127 VSUBS 0.007192f
C192 B.n128 VSUBS 0.007192f
C193 B.n129 VSUBS 0.007192f
C194 B.n130 VSUBS 0.007192f
C195 B.n131 VSUBS 0.007192f
C196 B.n132 VSUBS 0.007192f
C197 B.n133 VSUBS 0.007192f
C198 B.n134 VSUBS 0.007192f
C199 B.n135 VSUBS 0.007192f
C200 B.n136 VSUBS 0.007192f
C201 B.n137 VSUBS 0.007192f
C202 B.n138 VSUBS 0.007192f
C203 B.n139 VSUBS 0.007192f
C204 B.n140 VSUBS 0.007192f
C205 B.n141 VSUBS 0.007192f
C206 B.n142 VSUBS 0.007192f
C207 B.n143 VSUBS 0.007192f
C208 B.n144 VSUBS 0.007192f
C209 B.n145 VSUBS 0.007192f
C210 B.n146 VSUBS 0.007192f
C211 B.n147 VSUBS 0.007192f
C212 B.n148 VSUBS 0.007192f
C213 B.n149 VSUBS 0.007192f
C214 B.n150 VSUBS 0.007192f
C215 B.n151 VSUBS 0.007192f
C216 B.n152 VSUBS 0.016952f
C217 B.n153 VSUBS 0.007192f
C218 B.n154 VSUBS 0.007192f
C219 B.n155 VSUBS 0.007192f
C220 B.n156 VSUBS 0.007192f
C221 B.n157 VSUBS 0.007192f
C222 B.n158 VSUBS 0.007192f
C223 B.n159 VSUBS 0.007192f
C224 B.n160 VSUBS 0.007192f
C225 B.n161 VSUBS 0.007192f
C226 B.n162 VSUBS 0.007192f
C227 B.n163 VSUBS 0.007192f
C228 B.n164 VSUBS 0.007192f
C229 B.n165 VSUBS 0.007192f
C230 B.n166 VSUBS 0.007192f
C231 B.n167 VSUBS 0.007192f
C232 B.n168 VSUBS 0.007192f
C233 B.n169 VSUBS 0.007192f
C234 B.n170 VSUBS 0.007192f
C235 B.n171 VSUBS 0.007192f
C236 B.n172 VSUBS 0.007192f
C237 B.n173 VSUBS 0.007192f
C238 B.n174 VSUBS 0.007192f
C239 B.n175 VSUBS 0.007192f
C240 B.n176 VSUBS 0.007192f
C241 B.n177 VSUBS 0.007192f
C242 B.n178 VSUBS 0.007192f
C243 B.n179 VSUBS 0.007192f
C244 B.n180 VSUBS 0.007192f
C245 B.n181 VSUBS 0.007192f
C246 B.n182 VSUBS 0.007192f
C247 B.n183 VSUBS 0.007192f
C248 B.n184 VSUBS 0.007192f
C249 B.n185 VSUBS 0.016471f
C250 B.n186 VSUBS 0.016471f
C251 B.n187 VSUBS 0.016952f
C252 B.n188 VSUBS 0.007192f
C253 B.n189 VSUBS 0.007192f
C254 B.n190 VSUBS 0.007192f
C255 B.n191 VSUBS 0.007192f
C256 B.n192 VSUBS 0.007192f
C257 B.n193 VSUBS 0.007192f
C258 B.n194 VSUBS 0.007192f
C259 B.n195 VSUBS 0.007192f
C260 B.n196 VSUBS 0.007192f
C261 B.n197 VSUBS 0.007192f
C262 B.n198 VSUBS 0.007192f
C263 B.n199 VSUBS 0.007192f
C264 B.n200 VSUBS 0.007192f
C265 B.n201 VSUBS 0.007192f
C266 B.n202 VSUBS 0.007192f
C267 B.n203 VSUBS 0.007192f
C268 B.n204 VSUBS 0.007192f
C269 B.n205 VSUBS 0.007192f
C270 B.n206 VSUBS 0.007192f
C271 B.n207 VSUBS 0.007192f
C272 B.n208 VSUBS 0.007192f
C273 B.n209 VSUBS 0.007192f
C274 B.n210 VSUBS 0.007192f
C275 B.n211 VSUBS 0.007192f
C276 B.n212 VSUBS 0.007192f
C277 B.n213 VSUBS 0.007192f
C278 B.n214 VSUBS 0.007192f
C279 B.n215 VSUBS 0.007192f
C280 B.n216 VSUBS 0.007192f
C281 B.n217 VSUBS 0.007192f
C282 B.n218 VSUBS 0.007192f
C283 B.n219 VSUBS 0.007192f
C284 B.n220 VSUBS 0.007192f
C285 B.n221 VSUBS 0.007192f
C286 B.n222 VSUBS 0.007192f
C287 B.n223 VSUBS 0.007192f
C288 B.n224 VSUBS 0.007192f
C289 B.n225 VSUBS 0.007192f
C290 B.n226 VSUBS 0.007192f
C291 B.n227 VSUBS 0.007192f
C292 B.n228 VSUBS 0.007192f
C293 B.n229 VSUBS 0.007192f
C294 B.n230 VSUBS 0.007192f
C295 B.n231 VSUBS 0.007192f
C296 B.n232 VSUBS 0.007192f
C297 B.n233 VSUBS 0.007192f
C298 B.n234 VSUBS 0.007192f
C299 B.n235 VSUBS 0.007192f
C300 B.n236 VSUBS 0.007192f
C301 B.n237 VSUBS 0.007192f
C302 B.n238 VSUBS 0.007192f
C303 B.n239 VSUBS 0.007192f
C304 B.n240 VSUBS 0.007192f
C305 B.n241 VSUBS 0.007192f
C306 B.n242 VSUBS 0.007192f
C307 B.n243 VSUBS 0.007192f
C308 B.n244 VSUBS 0.007192f
C309 B.n245 VSUBS 0.007192f
C310 B.n246 VSUBS 0.007192f
C311 B.n247 VSUBS 0.007192f
C312 B.n248 VSUBS 0.007192f
C313 B.n249 VSUBS 0.007192f
C314 B.n250 VSUBS 0.007192f
C315 B.n251 VSUBS 0.007192f
C316 B.n252 VSUBS 0.007192f
C317 B.n253 VSUBS 0.007192f
C318 B.n254 VSUBS 0.007192f
C319 B.n255 VSUBS 0.007192f
C320 B.n256 VSUBS 0.007192f
C321 B.n257 VSUBS 0.007192f
C322 B.n258 VSUBS 0.007192f
C323 B.n259 VSUBS 0.007192f
C324 B.n260 VSUBS 0.007192f
C325 B.n261 VSUBS 0.007192f
C326 B.n262 VSUBS 0.007192f
C327 B.n263 VSUBS 0.006769f
C328 B.n264 VSUBS 0.007192f
C329 B.n265 VSUBS 0.007192f
C330 B.n266 VSUBS 0.004019f
C331 B.n267 VSUBS 0.007192f
C332 B.n268 VSUBS 0.007192f
C333 B.n269 VSUBS 0.007192f
C334 B.n270 VSUBS 0.007192f
C335 B.n271 VSUBS 0.007192f
C336 B.n272 VSUBS 0.007192f
C337 B.n273 VSUBS 0.007192f
C338 B.n274 VSUBS 0.007192f
C339 B.n275 VSUBS 0.007192f
C340 B.n276 VSUBS 0.007192f
C341 B.n277 VSUBS 0.007192f
C342 B.n278 VSUBS 0.007192f
C343 B.n279 VSUBS 0.004019f
C344 B.n280 VSUBS 0.016664f
C345 B.n281 VSUBS 0.006769f
C346 B.n282 VSUBS 0.007192f
C347 B.n283 VSUBS 0.007192f
C348 B.n284 VSUBS 0.007192f
C349 B.n285 VSUBS 0.007192f
C350 B.n286 VSUBS 0.007192f
C351 B.n287 VSUBS 0.007192f
C352 B.n288 VSUBS 0.007192f
C353 B.n289 VSUBS 0.007192f
C354 B.n290 VSUBS 0.007192f
C355 B.n291 VSUBS 0.007192f
C356 B.n292 VSUBS 0.007192f
C357 B.n293 VSUBS 0.007192f
C358 B.n294 VSUBS 0.007192f
C359 B.n295 VSUBS 0.007192f
C360 B.n296 VSUBS 0.007192f
C361 B.n297 VSUBS 0.007192f
C362 B.n298 VSUBS 0.007192f
C363 B.n299 VSUBS 0.007192f
C364 B.n300 VSUBS 0.007192f
C365 B.n301 VSUBS 0.007192f
C366 B.n302 VSUBS 0.007192f
C367 B.n303 VSUBS 0.007192f
C368 B.n304 VSUBS 0.007192f
C369 B.n305 VSUBS 0.007192f
C370 B.n306 VSUBS 0.007192f
C371 B.n307 VSUBS 0.007192f
C372 B.n308 VSUBS 0.007192f
C373 B.n309 VSUBS 0.007192f
C374 B.n310 VSUBS 0.007192f
C375 B.n311 VSUBS 0.007192f
C376 B.n312 VSUBS 0.007192f
C377 B.n313 VSUBS 0.007192f
C378 B.n314 VSUBS 0.007192f
C379 B.n315 VSUBS 0.007192f
C380 B.n316 VSUBS 0.007192f
C381 B.n317 VSUBS 0.007192f
C382 B.n318 VSUBS 0.007192f
C383 B.n319 VSUBS 0.007192f
C384 B.n320 VSUBS 0.007192f
C385 B.n321 VSUBS 0.007192f
C386 B.n322 VSUBS 0.007192f
C387 B.n323 VSUBS 0.007192f
C388 B.n324 VSUBS 0.007192f
C389 B.n325 VSUBS 0.007192f
C390 B.n326 VSUBS 0.007192f
C391 B.n327 VSUBS 0.007192f
C392 B.n328 VSUBS 0.007192f
C393 B.n329 VSUBS 0.007192f
C394 B.n330 VSUBS 0.007192f
C395 B.n331 VSUBS 0.007192f
C396 B.n332 VSUBS 0.007192f
C397 B.n333 VSUBS 0.007192f
C398 B.n334 VSUBS 0.007192f
C399 B.n335 VSUBS 0.007192f
C400 B.n336 VSUBS 0.007192f
C401 B.n337 VSUBS 0.007192f
C402 B.n338 VSUBS 0.007192f
C403 B.n339 VSUBS 0.007192f
C404 B.n340 VSUBS 0.007192f
C405 B.n341 VSUBS 0.007192f
C406 B.n342 VSUBS 0.007192f
C407 B.n343 VSUBS 0.007192f
C408 B.n344 VSUBS 0.007192f
C409 B.n345 VSUBS 0.007192f
C410 B.n346 VSUBS 0.007192f
C411 B.n347 VSUBS 0.007192f
C412 B.n348 VSUBS 0.007192f
C413 B.n349 VSUBS 0.007192f
C414 B.n350 VSUBS 0.007192f
C415 B.n351 VSUBS 0.007192f
C416 B.n352 VSUBS 0.007192f
C417 B.n353 VSUBS 0.007192f
C418 B.n354 VSUBS 0.007192f
C419 B.n355 VSUBS 0.007192f
C420 B.n356 VSUBS 0.007192f
C421 B.n357 VSUBS 0.007192f
C422 B.n358 VSUBS 0.016952f
C423 B.n359 VSUBS 0.016471f
C424 B.n360 VSUBS 0.016471f
C425 B.n361 VSUBS 0.007192f
C426 B.n362 VSUBS 0.007192f
C427 B.n363 VSUBS 0.007192f
C428 B.n364 VSUBS 0.007192f
C429 B.n365 VSUBS 0.007192f
C430 B.n366 VSUBS 0.007192f
C431 B.n367 VSUBS 0.007192f
C432 B.n368 VSUBS 0.007192f
C433 B.n369 VSUBS 0.007192f
C434 B.n370 VSUBS 0.007192f
C435 B.n371 VSUBS 0.007192f
C436 B.n372 VSUBS 0.007192f
C437 B.n373 VSUBS 0.007192f
C438 B.n374 VSUBS 0.007192f
C439 B.n375 VSUBS 0.007192f
C440 B.n376 VSUBS 0.007192f
C441 B.n377 VSUBS 0.007192f
C442 B.n378 VSUBS 0.007192f
C443 B.n379 VSUBS 0.007192f
C444 B.n380 VSUBS 0.007192f
C445 B.n381 VSUBS 0.007192f
C446 B.n382 VSUBS 0.007192f
C447 B.n383 VSUBS 0.007192f
C448 B.n384 VSUBS 0.007192f
C449 B.n385 VSUBS 0.007192f
C450 B.n386 VSUBS 0.007192f
C451 B.n387 VSUBS 0.007192f
C452 B.n388 VSUBS 0.007192f
C453 B.n389 VSUBS 0.007192f
C454 B.n390 VSUBS 0.007192f
C455 B.n391 VSUBS 0.007192f
C456 B.n392 VSUBS 0.007192f
C457 B.n393 VSUBS 0.007192f
C458 B.n394 VSUBS 0.007192f
C459 B.n395 VSUBS 0.007192f
C460 B.n396 VSUBS 0.007192f
C461 B.n397 VSUBS 0.007192f
C462 B.n398 VSUBS 0.007192f
C463 B.n399 VSUBS 0.007192f
C464 B.n400 VSUBS 0.007192f
C465 B.n401 VSUBS 0.007192f
C466 B.n402 VSUBS 0.007192f
C467 B.n403 VSUBS 0.007192f
C468 B.n404 VSUBS 0.007192f
C469 B.n405 VSUBS 0.007192f
C470 B.n406 VSUBS 0.007192f
C471 B.n407 VSUBS 0.007192f
C472 B.n408 VSUBS 0.007192f
C473 B.n409 VSUBS 0.007192f
C474 B.n410 VSUBS 0.007192f
C475 B.n411 VSUBS 0.007192f
C476 B.n412 VSUBS 0.007192f
C477 B.n413 VSUBS 0.017329f
C478 B.n414 VSUBS 0.016471f
C479 B.n415 VSUBS 0.016952f
C480 B.n416 VSUBS 0.007192f
C481 B.n417 VSUBS 0.007192f
C482 B.n418 VSUBS 0.007192f
C483 B.n419 VSUBS 0.007192f
C484 B.n420 VSUBS 0.007192f
C485 B.n421 VSUBS 0.007192f
C486 B.n422 VSUBS 0.007192f
C487 B.n423 VSUBS 0.007192f
C488 B.n424 VSUBS 0.007192f
C489 B.n425 VSUBS 0.007192f
C490 B.n426 VSUBS 0.007192f
C491 B.n427 VSUBS 0.007192f
C492 B.n428 VSUBS 0.007192f
C493 B.n429 VSUBS 0.007192f
C494 B.n430 VSUBS 0.007192f
C495 B.n431 VSUBS 0.007192f
C496 B.n432 VSUBS 0.007192f
C497 B.n433 VSUBS 0.007192f
C498 B.n434 VSUBS 0.007192f
C499 B.n435 VSUBS 0.007192f
C500 B.n436 VSUBS 0.007192f
C501 B.n437 VSUBS 0.007192f
C502 B.n438 VSUBS 0.007192f
C503 B.n439 VSUBS 0.007192f
C504 B.n440 VSUBS 0.007192f
C505 B.n441 VSUBS 0.007192f
C506 B.n442 VSUBS 0.007192f
C507 B.n443 VSUBS 0.007192f
C508 B.n444 VSUBS 0.007192f
C509 B.n445 VSUBS 0.007192f
C510 B.n446 VSUBS 0.007192f
C511 B.n447 VSUBS 0.007192f
C512 B.n448 VSUBS 0.007192f
C513 B.n449 VSUBS 0.007192f
C514 B.n450 VSUBS 0.007192f
C515 B.n451 VSUBS 0.007192f
C516 B.n452 VSUBS 0.007192f
C517 B.n453 VSUBS 0.007192f
C518 B.n454 VSUBS 0.007192f
C519 B.n455 VSUBS 0.007192f
C520 B.n456 VSUBS 0.007192f
C521 B.n457 VSUBS 0.007192f
C522 B.n458 VSUBS 0.007192f
C523 B.n459 VSUBS 0.007192f
C524 B.n460 VSUBS 0.007192f
C525 B.n461 VSUBS 0.007192f
C526 B.n462 VSUBS 0.007192f
C527 B.n463 VSUBS 0.007192f
C528 B.n464 VSUBS 0.007192f
C529 B.n465 VSUBS 0.007192f
C530 B.n466 VSUBS 0.007192f
C531 B.n467 VSUBS 0.007192f
C532 B.n468 VSUBS 0.007192f
C533 B.n469 VSUBS 0.007192f
C534 B.n470 VSUBS 0.007192f
C535 B.n471 VSUBS 0.007192f
C536 B.n472 VSUBS 0.007192f
C537 B.n473 VSUBS 0.007192f
C538 B.n474 VSUBS 0.007192f
C539 B.n475 VSUBS 0.007192f
C540 B.n476 VSUBS 0.007192f
C541 B.n477 VSUBS 0.007192f
C542 B.n478 VSUBS 0.007192f
C543 B.n479 VSUBS 0.007192f
C544 B.n480 VSUBS 0.007192f
C545 B.n481 VSUBS 0.007192f
C546 B.n482 VSUBS 0.007192f
C547 B.n483 VSUBS 0.007192f
C548 B.n484 VSUBS 0.007192f
C549 B.n485 VSUBS 0.007192f
C550 B.n486 VSUBS 0.007192f
C551 B.n487 VSUBS 0.007192f
C552 B.n488 VSUBS 0.007192f
C553 B.n489 VSUBS 0.007192f
C554 B.n490 VSUBS 0.007192f
C555 B.n491 VSUBS 0.006769f
C556 B.n492 VSUBS 0.007192f
C557 B.n493 VSUBS 0.007192f
C558 B.n494 VSUBS 0.004019f
C559 B.n495 VSUBS 0.007192f
C560 B.n496 VSUBS 0.007192f
C561 B.n497 VSUBS 0.007192f
C562 B.n498 VSUBS 0.007192f
C563 B.n499 VSUBS 0.007192f
C564 B.n500 VSUBS 0.007192f
C565 B.n501 VSUBS 0.007192f
C566 B.n502 VSUBS 0.007192f
C567 B.n503 VSUBS 0.007192f
C568 B.n504 VSUBS 0.007192f
C569 B.n505 VSUBS 0.007192f
C570 B.n506 VSUBS 0.007192f
C571 B.n507 VSUBS 0.004019f
C572 B.n508 VSUBS 0.016664f
C573 B.n509 VSUBS 0.006769f
C574 B.n510 VSUBS 0.007192f
C575 B.n511 VSUBS 0.007192f
C576 B.n512 VSUBS 0.007192f
C577 B.n513 VSUBS 0.007192f
C578 B.n514 VSUBS 0.007192f
C579 B.n515 VSUBS 0.007192f
C580 B.n516 VSUBS 0.007192f
C581 B.n517 VSUBS 0.007192f
C582 B.n518 VSUBS 0.007192f
C583 B.n519 VSUBS 0.007192f
C584 B.n520 VSUBS 0.007192f
C585 B.n521 VSUBS 0.007192f
C586 B.n522 VSUBS 0.007192f
C587 B.n523 VSUBS 0.007192f
C588 B.n524 VSUBS 0.007192f
C589 B.n525 VSUBS 0.007192f
C590 B.n526 VSUBS 0.007192f
C591 B.n527 VSUBS 0.007192f
C592 B.n528 VSUBS 0.007192f
C593 B.n529 VSUBS 0.007192f
C594 B.n530 VSUBS 0.007192f
C595 B.n531 VSUBS 0.007192f
C596 B.n532 VSUBS 0.007192f
C597 B.n533 VSUBS 0.007192f
C598 B.n534 VSUBS 0.007192f
C599 B.n535 VSUBS 0.007192f
C600 B.n536 VSUBS 0.007192f
C601 B.n537 VSUBS 0.007192f
C602 B.n538 VSUBS 0.007192f
C603 B.n539 VSUBS 0.007192f
C604 B.n540 VSUBS 0.007192f
C605 B.n541 VSUBS 0.007192f
C606 B.n542 VSUBS 0.007192f
C607 B.n543 VSUBS 0.007192f
C608 B.n544 VSUBS 0.007192f
C609 B.n545 VSUBS 0.007192f
C610 B.n546 VSUBS 0.007192f
C611 B.n547 VSUBS 0.007192f
C612 B.n548 VSUBS 0.007192f
C613 B.n549 VSUBS 0.007192f
C614 B.n550 VSUBS 0.007192f
C615 B.n551 VSUBS 0.007192f
C616 B.n552 VSUBS 0.007192f
C617 B.n553 VSUBS 0.007192f
C618 B.n554 VSUBS 0.007192f
C619 B.n555 VSUBS 0.007192f
C620 B.n556 VSUBS 0.007192f
C621 B.n557 VSUBS 0.007192f
C622 B.n558 VSUBS 0.007192f
C623 B.n559 VSUBS 0.007192f
C624 B.n560 VSUBS 0.007192f
C625 B.n561 VSUBS 0.007192f
C626 B.n562 VSUBS 0.007192f
C627 B.n563 VSUBS 0.007192f
C628 B.n564 VSUBS 0.007192f
C629 B.n565 VSUBS 0.007192f
C630 B.n566 VSUBS 0.007192f
C631 B.n567 VSUBS 0.007192f
C632 B.n568 VSUBS 0.007192f
C633 B.n569 VSUBS 0.007192f
C634 B.n570 VSUBS 0.007192f
C635 B.n571 VSUBS 0.007192f
C636 B.n572 VSUBS 0.007192f
C637 B.n573 VSUBS 0.007192f
C638 B.n574 VSUBS 0.007192f
C639 B.n575 VSUBS 0.007192f
C640 B.n576 VSUBS 0.007192f
C641 B.n577 VSUBS 0.007192f
C642 B.n578 VSUBS 0.007192f
C643 B.n579 VSUBS 0.007192f
C644 B.n580 VSUBS 0.007192f
C645 B.n581 VSUBS 0.007192f
C646 B.n582 VSUBS 0.007192f
C647 B.n583 VSUBS 0.007192f
C648 B.n584 VSUBS 0.007192f
C649 B.n585 VSUBS 0.007192f
C650 B.n586 VSUBS 0.016952f
C651 B.n587 VSUBS 0.016471f
C652 B.n588 VSUBS 0.016471f
C653 B.n589 VSUBS 0.007192f
C654 B.n590 VSUBS 0.007192f
C655 B.n591 VSUBS 0.007192f
C656 B.n592 VSUBS 0.007192f
C657 B.n593 VSUBS 0.007192f
C658 B.n594 VSUBS 0.007192f
C659 B.n595 VSUBS 0.007192f
C660 B.n596 VSUBS 0.007192f
C661 B.n597 VSUBS 0.007192f
C662 B.n598 VSUBS 0.007192f
C663 B.n599 VSUBS 0.007192f
C664 B.n600 VSUBS 0.007192f
C665 B.n601 VSUBS 0.007192f
C666 B.n602 VSUBS 0.007192f
C667 B.n603 VSUBS 0.007192f
C668 B.n604 VSUBS 0.007192f
C669 B.n605 VSUBS 0.007192f
C670 B.n606 VSUBS 0.007192f
C671 B.n607 VSUBS 0.007192f
C672 B.n608 VSUBS 0.007192f
C673 B.n609 VSUBS 0.007192f
C674 B.n610 VSUBS 0.007192f
C675 B.n611 VSUBS 0.007192f
C676 B.n612 VSUBS 0.007192f
C677 B.n613 VSUBS 0.007192f
C678 B.n614 VSUBS 0.007192f
C679 B.n615 VSUBS 0.016286f
C680 VDD1.t5 VSUBS 3.58954f
C681 VDD1.t4 VSUBS 3.58835f
C682 VDD1.t1 VSUBS 0.338958f
C683 VDD1.t0 VSUBS 0.338958f
C684 VDD1.n0 VSUBS 2.75887f
C685 VDD1.n1 VSUBS 3.16283f
C686 VDD1.t3 VSUBS 0.338958f
C687 VDD1.t2 VSUBS 0.338958f
C688 VDD1.n2 VSUBS 2.75773f
C689 VDD1.n3 VSUBS 3.0301f
C690 VTAIL.t1 VSUBS 0.368643f
C691 VTAIL.t3 VSUBS 0.368643f
C692 VTAIL.n0 VSUBS 2.8129f
C693 VTAIL.n1 VSUBS 0.832471f
C694 VTAIL.t10 VSUBS 3.68519f
C695 VTAIL.n2 VSUBS 1.01155f
C696 VTAIL.t8 VSUBS 0.368643f
C697 VTAIL.t7 VSUBS 0.368643f
C698 VTAIL.n3 VSUBS 2.8129f
C699 VTAIL.n4 VSUBS 2.63746f
C700 VTAIL.t5 VSUBS 0.368643f
C701 VTAIL.t2 VSUBS 0.368643f
C702 VTAIL.n5 VSUBS 2.81291f
C703 VTAIL.n6 VSUBS 2.63745f
C704 VTAIL.t0 VSUBS 3.68522f
C705 VTAIL.n7 VSUBS 1.01152f
C706 VTAIL.t9 VSUBS 0.368643f
C707 VTAIL.t6 VSUBS 0.368643f
C708 VTAIL.n8 VSUBS 2.81291f
C709 VTAIL.n9 VSUBS 0.878449f
C710 VTAIL.t11 VSUBS 3.68519f
C711 VTAIL.n10 VSUBS 2.70179f
C712 VTAIL.t4 VSUBS 3.68519f
C713 VTAIL.n11 VSUBS 2.679f
C714 VP.n0 VSUBS 0.083109f
C715 VP.t0 VSUBS 1.4033f
C716 VP.n1 VSUBS 0.521471f
C717 VP.t3 VSUBS 1.38653f
C718 VP.t2 VSUBS 1.38653f
C719 VP.n2 VSUBS 0.551161f
C720 VP.n3 VSUBS 0.536994f
C721 VP.n4 VSUBS 2.88795f
C722 VP.n5 VSUBS 2.76877f
C723 VP.t1 VSUBS 1.38653f
C724 VP.n6 VSUBS 0.536994f
C725 VP.t4 VSUBS 1.38653f
C726 VP.n7 VSUBS 0.55116f
C727 VP.t5 VSUBS 1.38653f
C728 VP.n8 VSUBS 0.536994f
C729 VP.n9 VSUBS 0.069255f
.ends

