* NGSPICE file created from diff_pair_sample_1658.ext - technology: sky130A

.subckt diff_pair_sample_1658 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1420_n4080# sky130_fd_pr__pfet_01v8 ad=6.0684 pd=31.9 as=0 ps=0 w=15.56 l=0.42
X1 VTAIL.t7 VN.t0 VDD2.t3 w_n1420_n4080# sky130_fd_pr__pfet_01v8 ad=6.0684 pd=31.9 as=2.5674 ps=15.89 w=15.56 l=0.42
X2 VTAIL.t1 VP.t0 VDD1.t3 w_n1420_n4080# sky130_fd_pr__pfet_01v8 ad=6.0684 pd=31.9 as=2.5674 ps=15.89 w=15.56 l=0.42
X3 B.t8 B.t6 B.t7 w_n1420_n4080# sky130_fd_pr__pfet_01v8 ad=6.0684 pd=31.9 as=0 ps=0 w=15.56 l=0.42
X4 VTAIL.t2 VP.t1 VDD1.t2 w_n1420_n4080# sky130_fd_pr__pfet_01v8 ad=6.0684 pd=31.9 as=2.5674 ps=15.89 w=15.56 l=0.42
X5 VDD2.t0 VN.t1 VTAIL.t6 w_n1420_n4080# sky130_fd_pr__pfet_01v8 ad=2.5674 pd=15.89 as=6.0684 ps=31.9 w=15.56 l=0.42
X6 VDD1.t1 VP.t2 VTAIL.t0 w_n1420_n4080# sky130_fd_pr__pfet_01v8 ad=2.5674 pd=15.89 as=6.0684 ps=31.9 w=15.56 l=0.42
X7 VDD1.t0 VP.t3 VTAIL.t3 w_n1420_n4080# sky130_fd_pr__pfet_01v8 ad=2.5674 pd=15.89 as=6.0684 ps=31.9 w=15.56 l=0.42
X8 B.t5 B.t3 B.t4 w_n1420_n4080# sky130_fd_pr__pfet_01v8 ad=6.0684 pd=31.9 as=0 ps=0 w=15.56 l=0.42
X9 VTAIL.t5 VN.t2 VDD2.t2 w_n1420_n4080# sky130_fd_pr__pfet_01v8 ad=6.0684 pd=31.9 as=2.5674 ps=15.89 w=15.56 l=0.42
X10 B.t2 B.t0 B.t1 w_n1420_n4080# sky130_fd_pr__pfet_01v8 ad=6.0684 pd=31.9 as=0 ps=0 w=15.56 l=0.42
X11 VDD2.t1 VN.t3 VTAIL.t4 w_n1420_n4080# sky130_fd_pr__pfet_01v8 ad=2.5674 pd=15.89 as=6.0684 ps=31.9 w=15.56 l=0.42
R0 B.n112 B.t3 1102.28
R1 B.n42 B.t6 1102.28
R2 B.n247 B.t0 1102.12
R3 B.n36 B.t9 1102.12
R4 B.n345 B.n344 585
R5 B.n343 B.n86 585
R6 B.n342 B.n341 585
R7 B.n340 B.n87 585
R8 B.n339 B.n338 585
R9 B.n337 B.n88 585
R10 B.n336 B.n335 585
R11 B.n334 B.n89 585
R12 B.n333 B.n332 585
R13 B.n331 B.n90 585
R14 B.n330 B.n329 585
R15 B.n328 B.n91 585
R16 B.n327 B.n326 585
R17 B.n325 B.n92 585
R18 B.n324 B.n323 585
R19 B.n322 B.n93 585
R20 B.n321 B.n320 585
R21 B.n319 B.n94 585
R22 B.n318 B.n317 585
R23 B.n316 B.n95 585
R24 B.n315 B.n314 585
R25 B.n313 B.n96 585
R26 B.n312 B.n311 585
R27 B.n310 B.n97 585
R28 B.n309 B.n308 585
R29 B.n307 B.n98 585
R30 B.n306 B.n305 585
R31 B.n304 B.n99 585
R32 B.n303 B.n302 585
R33 B.n301 B.n100 585
R34 B.n300 B.n299 585
R35 B.n298 B.n101 585
R36 B.n297 B.n296 585
R37 B.n295 B.n102 585
R38 B.n294 B.n293 585
R39 B.n292 B.n103 585
R40 B.n291 B.n290 585
R41 B.n289 B.n104 585
R42 B.n288 B.n287 585
R43 B.n286 B.n105 585
R44 B.n285 B.n284 585
R45 B.n283 B.n106 585
R46 B.n282 B.n281 585
R47 B.n280 B.n107 585
R48 B.n279 B.n278 585
R49 B.n277 B.n108 585
R50 B.n276 B.n275 585
R51 B.n274 B.n109 585
R52 B.n273 B.n272 585
R53 B.n271 B.n110 585
R54 B.n270 B.n269 585
R55 B.n268 B.n111 585
R56 B.n266 B.n265 585
R57 B.n264 B.n114 585
R58 B.n263 B.n262 585
R59 B.n261 B.n115 585
R60 B.n260 B.n259 585
R61 B.n258 B.n116 585
R62 B.n257 B.n256 585
R63 B.n255 B.n117 585
R64 B.n254 B.n253 585
R65 B.n252 B.n118 585
R66 B.n251 B.n250 585
R67 B.n246 B.n119 585
R68 B.n245 B.n244 585
R69 B.n243 B.n120 585
R70 B.n242 B.n241 585
R71 B.n240 B.n121 585
R72 B.n239 B.n238 585
R73 B.n237 B.n122 585
R74 B.n236 B.n235 585
R75 B.n234 B.n123 585
R76 B.n233 B.n232 585
R77 B.n231 B.n124 585
R78 B.n230 B.n229 585
R79 B.n228 B.n125 585
R80 B.n227 B.n226 585
R81 B.n225 B.n126 585
R82 B.n224 B.n223 585
R83 B.n222 B.n127 585
R84 B.n221 B.n220 585
R85 B.n219 B.n128 585
R86 B.n218 B.n217 585
R87 B.n216 B.n129 585
R88 B.n215 B.n214 585
R89 B.n213 B.n130 585
R90 B.n212 B.n211 585
R91 B.n210 B.n131 585
R92 B.n209 B.n208 585
R93 B.n207 B.n132 585
R94 B.n206 B.n205 585
R95 B.n204 B.n133 585
R96 B.n203 B.n202 585
R97 B.n201 B.n134 585
R98 B.n200 B.n199 585
R99 B.n198 B.n135 585
R100 B.n197 B.n196 585
R101 B.n195 B.n136 585
R102 B.n194 B.n193 585
R103 B.n192 B.n137 585
R104 B.n191 B.n190 585
R105 B.n189 B.n138 585
R106 B.n188 B.n187 585
R107 B.n186 B.n139 585
R108 B.n185 B.n184 585
R109 B.n183 B.n140 585
R110 B.n182 B.n181 585
R111 B.n180 B.n141 585
R112 B.n179 B.n178 585
R113 B.n177 B.n142 585
R114 B.n176 B.n175 585
R115 B.n174 B.n143 585
R116 B.n173 B.n172 585
R117 B.n171 B.n144 585
R118 B.n346 B.n85 585
R119 B.n348 B.n347 585
R120 B.n349 B.n84 585
R121 B.n351 B.n350 585
R122 B.n352 B.n83 585
R123 B.n354 B.n353 585
R124 B.n355 B.n82 585
R125 B.n357 B.n356 585
R126 B.n358 B.n81 585
R127 B.n360 B.n359 585
R128 B.n361 B.n80 585
R129 B.n363 B.n362 585
R130 B.n364 B.n79 585
R131 B.n366 B.n365 585
R132 B.n367 B.n78 585
R133 B.n369 B.n368 585
R134 B.n370 B.n77 585
R135 B.n372 B.n371 585
R136 B.n373 B.n76 585
R137 B.n375 B.n374 585
R138 B.n376 B.n75 585
R139 B.n378 B.n377 585
R140 B.n379 B.n74 585
R141 B.n381 B.n380 585
R142 B.n382 B.n73 585
R143 B.n384 B.n383 585
R144 B.n385 B.n72 585
R145 B.n387 B.n386 585
R146 B.n388 B.n71 585
R147 B.n390 B.n389 585
R148 B.n562 B.n9 585
R149 B.n561 B.n560 585
R150 B.n559 B.n10 585
R151 B.n558 B.n557 585
R152 B.n556 B.n11 585
R153 B.n555 B.n554 585
R154 B.n553 B.n12 585
R155 B.n552 B.n551 585
R156 B.n550 B.n13 585
R157 B.n549 B.n548 585
R158 B.n547 B.n14 585
R159 B.n546 B.n545 585
R160 B.n544 B.n15 585
R161 B.n543 B.n542 585
R162 B.n541 B.n16 585
R163 B.n540 B.n539 585
R164 B.n538 B.n17 585
R165 B.n537 B.n536 585
R166 B.n535 B.n18 585
R167 B.n534 B.n533 585
R168 B.n532 B.n19 585
R169 B.n531 B.n530 585
R170 B.n529 B.n20 585
R171 B.n528 B.n527 585
R172 B.n526 B.n21 585
R173 B.n525 B.n524 585
R174 B.n523 B.n22 585
R175 B.n522 B.n521 585
R176 B.n520 B.n23 585
R177 B.n519 B.n518 585
R178 B.n517 B.n24 585
R179 B.n516 B.n515 585
R180 B.n514 B.n25 585
R181 B.n513 B.n512 585
R182 B.n511 B.n26 585
R183 B.n510 B.n509 585
R184 B.n508 B.n27 585
R185 B.n507 B.n506 585
R186 B.n505 B.n28 585
R187 B.n504 B.n503 585
R188 B.n502 B.n29 585
R189 B.n501 B.n500 585
R190 B.n499 B.n30 585
R191 B.n498 B.n497 585
R192 B.n496 B.n31 585
R193 B.n495 B.n494 585
R194 B.n493 B.n32 585
R195 B.n492 B.n491 585
R196 B.n490 B.n33 585
R197 B.n489 B.n488 585
R198 B.n487 B.n34 585
R199 B.n486 B.n485 585
R200 B.n483 B.n35 585
R201 B.n482 B.n481 585
R202 B.n480 B.n38 585
R203 B.n479 B.n478 585
R204 B.n477 B.n39 585
R205 B.n476 B.n475 585
R206 B.n474 B.n40 585
R207 B.n473 B.n472 585
R208 B.n471 B.n41 585
R209 B.n470 B.n469 585
R210 B.n468 B.n467 585
R211 B.n466 B.n45 585
R212 B.n465 B.n464 585
R213 B.n463 B.n46 585
R214 B.n462 B.n461 585
R215 B.n460 B.n47 585
R216 B.n459 B.n458 585
R217 B.n457 B.n48 585
R218 B.n456 B.n455 585
R219 B.n454 B.n49 585
R220 B.n453 B.n452 585
R221 B.n451 B.n50 585
R222 B.n450 B.n449 585
R223 B.n448 B.n51 585
R224 B.n447 B.n446 585
R225 B.n445 B.n52 585
R226 B.n444 B.n443 585
R227 B.n442 B.n53 585
R228 B.n441 B.n440 585
R229 B.n439 B.n54 585
R230 B.n438 B.n437 585
R231 B.n436 B.n55 585
R232 B.n435 B.n434 585
R233 B.n433 B.n56 585
R234 B.n432 B.n431 585
R235 B.n430 B.n57 585
R236 B.n429 B.n428 585
R237 B.n427 B.n58 585
R238 B.n426 B.n425 585
R239 B.n424 B.n59 585
R240 B.n423 B.n422 585
R241 B.n421 B.n60 585
R242 B.n420 B.n419 585
R243 B.n418 B.n61 585
R244 B.n417 B.n416 585
R245 B.n415 B.n62 585
R246 B.n414 B.n413 585
R247 B.n412 B.n63 585
R248 B.n411 B.n410 585
R249 B.n409 B.n64 585
R250 B.n408 B.n407 585
R251 B.n406 B.n65 585
R252 B.n405 B.n404 585
R253 B.n403 B.n66 585
R254 B.n402 B.n401 585
R255 B.n400 B.n67 585
R256 B.n399 B.n398 585
R257 B.n397 B.n68 585
R258 B.n396 B.n395 585
R259 B.n394 B.n69 585
R260 B.n393 B.n392 585
R261 B.n391 B.n70 585
R262 B.n564 B.n563 585
R263 B.n565 B.n8 585
R264 B.n567 B.n566 585
R265 B.n568 B.n7 585
R266 B.n570 B.n569 585
R267 B.n571 B.n6 585
R268 B.n573 B.n572 585
R269 B.n574 B.n5 585
R270 B.n576 B.n575 585
R271 B.n577 B.n4 585
R272 B.n579 B.n578 585
R273 B.n580 B.n3 585
R274 B.n582 B.n581 585
R275 B.n583 B.n0 585
R276 B.n2 B.n1 585
R277 B.n152 B.n151 585
R278 B.n153 B.n150 585
R279 B.n155 B.n154 585
R280 B.n156 B.n149 585
R281 B.n158 B.n157 585
R282 B.n159 B.n148 585
R283 B.n161 B.n160 585
R284 B.n162 B.n147 585
R285 B.n164 B.n163 585
R286 B.n165 B.n146 585
R287 B.n167 B.n166 585
R288 B.n168 B.n145 585
R289 B.n170 B.n169 585
R290 B.n171 B.n170 516.524
R291 B.n344 B.n85 516.524
R292 B.n391 B.n390 516.524
R293 B.n564 B.n9 516.524
R294 B.n112 B.t4 454.611
R295 B.n42 B.t8 454.611
R296 B.n247 B.t1 454.611
R297 B.n36 B.t11 454.611
R298 B.n113 B.t5 440.065
R299 B.n43 B.t7 440.065
R300 B.n248 B.t2 440.065
R301 B.n37 B.t10 440.065
R302 B.n585 B.n584 256.663
R303 B.n584 B.n583 235.042
R304 B.n584 B.n2 235.042
R305 B.n172 B.n171 163.367
R306 B.n172 B.n143 163.367
R307 B.n176 B.n143 163.367
R308 B.n177 B.n176 163.367
R309 B.n178 B.n177 163.367
R310 B.n178 B.n141 163.367
R311 B.n182 B.n141 163.367
R312 B.n183 B.n182 163.367
R313 B.n184 B.n183 163.367
R314 B.n184 B.n139 163.367
R315 B.n188 B.n139 163.367
R316 B.n189 B.n188 163.367
R317 B.n190 B.n189 163.367
R318 B.n190 B.n137 163.367
R319 B.n194 B.n137 163.367
R320 B.n195 B.n194 163.367
R321 B.n196 B.n195 163.367
R322 B.n196 B.n135 163.367
R323 B.n200 B.n135 163.367
R324 B.n201 B.n200 163.367
R325 B.n202 B.n201 163.367
R326 B.n202 B.n133 163.367
R327 B.n206 B.n133 163.367
R328 B.n207 B.n206 163.367
R329 B.n208 B.n207 163.367
R330 B.n208 B.n131 163.367
R331 B.n212 B.n131 163.367
R332 B.n213 B.n212 163.367
R333 B.n214 B.n213 163.367
R334 B.n214 B.n129 163.367
R335 B.n218 B.n129 163.367
R336 B.n219 B.n218 163.367
R337 B.n220 B.n219 163.367
R338 B.n220 B.n127 163.367
R339 B.n224 B.n127 163.367
R340 B.n225 B.n224 163.367
R341 B.n226 B.n225 163.367
R342 B.n226 B.n125 163.367
R343 B.n230 B.n125 163.367
R344 B.n231 B.n230 163.367
R345 B.n232 B.n231 163.367
R346 B.n232 B.n123 163.367
R347 B.n236 B.n123 163.367
R348 B.n237 B.n236 163.367
R349 B.n238 B.n237 163.367
R350 B.n238 B.n121 163.367
R351 B.n242 B.n121 163.367
R352 B.n243 B.n242 163.367
R353 B.n244 B.n243 163.367
R354 B.n244 B.n119 163.367
R355 B.n251 B.n119 163.367
R356 B.n252 B.n251 163.367
R357 B.n253 B.n252 163.367
R358 B.n253 B.n117 163.367
R359 B.n257 B.n117 163.367
R360 B.n258 B.n257 163.367
R361 B.n259 B.n258 163.367
R362 B.n259 B.n115 163.367
R363 B.n263 B.n115 163.367
R364 B.n264 B.n263 163.367
R365 B.n265 B.n264 163.367
R366 B.n265 B.n111 163.367
R367 B.n270 B.n111 163.367
R368 B.n271 B.n270 163.367
R369 B.n272 B.n271 163.367
R370 B.n272 B.n109 163.367
R371 B.n276 B.n109 163.367
R372 B.n277 B.n276 163.367
R373 B.n278 B.n277 163.367
R374 B.n278 B.n107 163.367
R375 B.n282 B.n107 163.367
R376 B.n283 B.n282 163.367
R377 B.n284 B.n283 163.367
R378 B.n284 B.n105 163.367
R379 B.n288 B.n105 163.367
R380 B.n289 B.n288 163.367
R381 B.n290 B.n289 163.367
R382 B.n290 B.n103 163.367
R383 B.n294 B.n103 163.367
R384 B.n295 B.n294 163.367
R385 B.n296 B.n295 163.367
R386 B.n296 B.n101 163.367
R387 B.n300 B.n101 163.367
R388 B.n301 B.n300 163.367
R389 B.n302 B.n301 163.367
R390 B.n302 B.n99 163.367
R391 B.n306 B.n99 163.367
R392 B.n307 B.n306 163.367
R393 B.n308 B.n307 163.367
R394 B.n308 B.n97 163.367
R395 B.n312 B.n97 163.367
R396 B.n313 B.n312 163.367
R397 B.n314 B.n313 163.367
R398 B.n314 B.n95 163.367
R399 B.n318 B.n95 163.367
R400 B.n319 B.n318 163.367
R401 B.n320 B.n319 163.367
R402 B.n320 B.n93 163.367
R403 B.n324 B.n93 163.367
R404 B.n325 B.n324 163.367
R405 B.n326 B.n325 163.367
R406 B.n326 B.n91 163.367
R407 B.n330 B.n91 163.367
R408 B.n331 B.n330 163.367
R409 B.n332 B.n331 163.367
R410 B.n332 B.n89 163.367
R411 B.n336 B.n89 163.367
R412 B.n337 B.n336 163.367
R413 B.n338 B.n337 163.367
R414 B.n338 B.n87 163.367
R415 B.n342 B.n87 163.367
R416 B.n343 B.n342 163.367
R417 B.n344 B.n343 163.367
R418 B.n390 B.n71 163.367
R419 B.n386 B.n71 163.367
R420 B.n386 B.n385 163.367
R421 B.n385 B.n384 163.367
R422 B.n384 B.n73 163.367
R423 B.n380 B.n73 163.367
R424 B.n380 B.n379 163.367
R425 B.n379 B.n378 163.367
R426 B.n378 B.n75 163.367
R427 B.n374 B.n75 163.367
R428 B.n374 B.n373 163.367
R429 B.n373 B.n372 163.367
R430 B.n372 B.n77 163.367
R431 B.n368 B.n77 163.367
R432 B.n368 B.n367 163.367
R433 B.n367 B.n366 163.367
R434 B.n366 B.n79 163.367
R435 B.n362 B.n79 163.367
R436 B.n362 B.n361 163.367
R437 B.n361 B.n360 163.367
R438 B.n360 B.n81 163.367
R439 B.n356 B.n81 163.367
R440 B.n356 B.n355 163.367
R441 B.n355 B.n354 163.367
R442 B.n354 B.n83 163.367
R443 B.n350 B.n83 163.367
R444 B.n350 B.n349 163.367
R445 B.n349 B.n348 163.367
R446 B.n348 B.n85 163.367
R447 B.n560 B.n9 163.367
R448 B.n560 B.n559 163.367
R449 B.n559 B.n558 163.367
R450 B.n558 B.n11 163.367
R451 B.n554 B.n11 163.367
R452 B.n554 B.n553 163.367
R453 B.n553 B.n552 163.367
R454 B.n552 B.n13 163.367
R455 B.n548 B.n13 163.367
R456 B.n548 B.n547 163.367
R457 B.n547 B.n546 163.367
R458 B.n546 B.n15 163.367
R459 B.n542 B.n15 163.367
R460 B.n542 B.n541 163.367
R461 B.n541 B.n540 163.367
R462 B.n540 B.n17 163.367
R463 B.n536 B.n17 163.367
R464 B.n536 B.n535 163.367
R465 B.n535 B.n534 163.367
R466 B.n534 B.n19 163.367
R467 B.n530 B.n19 163.367
R468 B.n530 B.n529 163.367
R469 B.n529 B.n528 163.367
R470 B.n528 B.n21 163.367
R471 B.n524 B.n21 163.367
R472 B.n524 B.n523 163.367
R473 B.n523 B.n522 163.367
R474 B.n522 B.n23 163.367
R475 B.n518 B.n23 163.367
R476 B.n518 B.n517 163.367
R477 B.n517 B.n516 163.367
R478 B.n516 B.n25 163.367
R479 B.n512 B.n25 163.367
R480 B.n512 B.n511 163.367
R481 B.n511 B.n510 163.367
R482 B.n510 B.n27 163.367
R483 B.n506 B.n27 163.367
R484 B.n506 B.n505 163.367
R485 B.n505 B.n504 163.367
R486 B.n504 B.n29 163.367
R487 B.n500 B.n29 163.367
R488 B.n500 B.n499 163.367
R489 B.n499 B.n498 163.367
R490 B.n498 B.n31 163.367
R491 B.n494 B.n31 163.367
R492 B.n494 B.n493 163.367
R493 B.n493 B.n492 163.367
R494 B.n492 B.n33 163.367
R495 B.n488 B.n33 163.367
R496 B.n488 B.n487 163.367
R497 B.n487 B.n486 163.367
R498 B.n486 B.n35 163.367
R499 B.n481 B.n35 163.367
R500 B.n481 B.n480 163.367
R501 B.n480 B.n479 163.367
R502 B.n479 B.n39 163.367
R503 B.n475 B.n39 163.367
R504 B.n475 B.n474 163.367
R505 B.n474 B.n473 163.367
R506 B.n473 B.n41 163.367
R507 B.n469 B.n41 163.367
R508 B.n469 B.n468 163.367
R509 B.n468 B.n45 163.367
R510 B.n464 B.n45 163.367
R511 B.n464 B.n463 163.367
R512 B.n463 B.n462 163.367
R513 B.n462 B.n47 163.367
R514 B.n458 B.n47 163.367
R515 B.n458 B.n457 163.367
R516 B.n457 B.n456 163.367
R517 B.n456 B.n49 163.367
R518 B.n452 B.n49 163.367
R519 B.n452 B.n451 163.367
R520 B.n451 B.n450 163.367
R521 B.n450 B.n51 163.367
R522 B.n446 B.n51 163.367
R523 B.n446 B.n445 163.367
R524 B.n445 B.n444 163.367
R525 B.n444 B.n53 163.367
R526 B.n440 B.n53 163.367
R527 B.n440 B.n439 163.367
R528 B.n439 B.n438 163.367
R529 B.n438 B.n55 163.367
R530 B.n434 B.n55 163.367
R531 B.n434 B.n433 163.367
R532 B.n433 B.n432 163.367
R533 B.n432 B.n57 163.367
R534 B.n428 B.n57 163.367
R535 B.n428 B.n427 163.367
R536 B.n427 B.n426 163.367
R537 B.n426 B.n59 163.367
R538 B.n422 B.n59 163.367
R539 B.n422 B.n421 163.367
R540 B.n421 B.n420 163.367
R541 B.n420 B.n61 163.367
R542 B.n416 B.n61 163.367
R543 B.n416 B.n415 163.367
R544 B.n415 B.n414 163.367
R545 B.n414 B.n63 163.367
R546 B.n410 B.n63 163.367
R547 B.n410 B.n409 163.367
R548 B.n409 B.n408 163.367
R549 B.n408 B.n65 163.367
R550 B.n404 B.n65 163.367
R551 B.n404 B.n403 163.367
R552 B.n403 B.n402 163.367
R553 B.n402 B.n67 163.367
R554 B.n398 B.n67 163.367
R555 B.n398 B.n397 163.367
R556 B.n397 B.n396 163.367
R557 B.n396 B.n69 163.367
R558 B.n392 B.n69 163.367
R559 B.n392 B.n391 163.367
R560 B.n565 B.n564 163.367
R561 B.n566 B.n565 163.367
R562 B.n566 B.n7 163.367
R563 B.n570 B.n7 163.367
R564 B.n571 B.n570 163.367
R565 B.n572 B.n571 163.367
R566 B.n572 B.n5 163.367
R567 B.n576 B.n5 163.367
R568 B.n577 B.n576 163.367
R569 B.n578 B.n577 163.367
R570 B.n578 B.n3 163.367
R571 B.n582 B.n3 163.367
R572 B.n583 B.n582 163.367
R573 B.n152 B.n2 163.367
R574 B.n153 B.n152 163.367
R575 B.n154 B.n153 163.367
R576 B.n154 B.n149 163.367
R577 B.n158 B.n149 163.367
R578 B.n159 B.n158 163.367
R579 B.n160 B.n159 163.367
R580 B.n160 B.n147 163.367
R581 B.n164 B.n147 163.367
R582 B.n165 B.n164 163.367
R583 B.n166 B.n165 163.367
R584 B.n166 B.n145 163.367
R585 B.n170 B.n145 163.367
R586 B.n249 B.n248 59.5399
R587 B.n267 B.n113 59.5399
R588 B.n44 B.n43 59.5399
R589 B.n484 B.n37 59.5399
R590 B.n563 B.n562 33.5615
R591 B.n389 B.n70 33.5615
R592 B.n346 B.n345 33.5615
R593 B.n169 B.n144 33.5615
R594 B B.n585 18.0485
R595 B.n248 B.n247 14.546
R596 B.n113 B.n112 14.546
R597 B.n43 B.n42 14.546
R598 B.n37 B.n36 14.546
R599 B.n563 B.n8 10.6151
R600 B.n567 B.n8 10.6151
R601 B.n568 B.n567 10.6151
R602 B.n569 B.n568 10.6151
R603 B.n569 B.n6 10.6151
R604 B.n573 B.n6 10.6151
R605 B.n574 B.n573 10.6151
R606 B.n575 B.n574 10.6151
R607 B.n575 B.n4 10.6151
R608 B.n579 B.n4 10.6151
R609 B.n580 B.n579 10.6151
R610 B.n581 B.n580 10.6151
R611 B.n581 B.n0 10.6151
R612 B.n562 B.n561 10.6151
R613 B.n561 B.n10 10.6151
R614 B.n557 B.n10 10.6151
R615 B.n557 B.n556 10.6151
R616 B.n556 B.n555 10.6151
R617 B.n555 B.n12 10.6151
R618 B.n551 B.n12 10.6151
R619 B.n551 B.n550 10.6151
R620 B.n550 B.n549 10.6151
R621 B.n549 B.n14 10.6151
R622 B.n545 B.n14 10.6151
R623 B.n545 B.n544 10.6151
R624 B.n544 B.n543 10.6151
R625 B.n543 B.n16 10.6151
R626 B.n539 B.n16 10.6151
R627 B.n539 B.n538 10.6151
R628 B.n538 B.n537 10.6151
R629 B.n537 B.n18 10.6151
R630 B.n533 B.n18 10.6151
R631 B.n533 B.n532 10.6151
R632 B.n532 B.n531 10.6151
R633 B.n531 B.n20 10.6151
R634 B.n527 B.n20 10.6151
R635 B.n527 B.n526 10.6151
R636 B.n526 B.n525 10.6151
R637 B.n525 B.n22 10.6151
R638 B.n521 B.n22 10.6151
R639 B.n521 B.n520 10.6151
R640 B.n520 B.n519 10.6151
R641 B.n519 B.n24 10.6151
R642 B.n515 B.n24 10.6151
R643 B.n515 B.n514 10.6151
R644 B.n514 B.n513 10.6151
R645 B.n513 B.n26 10.6151
R646 B.n509 B.n26 10.6151
R647 B.n509 B.n508 10.6151
R648 B.n508 B.n507 10.6151
R649 B.n507 B.n28 10.6151
R650 B.n503 B.n28 10.6151
R651 B.n503 B.n502 10.6151
R652 B.n502 B.n501 10.6151
R653 B.n501 B.n30 10.6151
R654 B.n497 B.n30 10.6151
R655 B.n497 B.n496 10.6151
R656 B.n496 B.n495 10.6151
R657 B.n495 B.n32 10.6151
R658 B.n491 B.n32 10.6151
R659 B.n491 B.n490 10.6151
R660 B.n490 B.n489 10.6151
R661 B.n489 B.n34 10.6151
R662 B.n485 B.n34 10.6151
R663 B.n483 B.n482 10.6151
R664 B.n482 B.n38 10.6151
R665 B.n478 B.n38 10.6151
R666 B.n478 B.n477 10.6151
R667 B.n477 B.n476 10.6151
R668 B.n476 B.n40 10.6151
R669 B.n472 B.n40 10.6151
R670 B.n472 B.n471 10.6151
R671 B.n471 B.n470 10.6151
R672 B.n467 B.n466 10.6151
R673 B.n466 B.n465 10.6151
R674 B.n465 B.n46 10.6151
R675 B.n461 B.n46 10.6151
R676 B.n461 B.n460 10.6151
R677 B.n460 B.n459 10.6151
R678 B.n459 B.n48 10.6151
R679 B.n455 B.n48 10.6151
R680 B.n455 B.n454 10.6151
R681 B.n454 B.n453 10.6151
R682 B.n453 B.n50 10.6151
R683 B.n449 B.n50 10.6151
R684 B.n449 B.n448 10.6151
R685 B.n448 B.n447 10.6151
R686 B.n447 B.n52 10.6151
R687 B.n443 B.n52 10.6151
R688 B.n443 B.n442 10.6151
R689 B.n442 B.n441 10.6151
R690 B.n441 B.n54 10.6151
R691 B.n437 B.n54 10.6151
R692 B.n437 B.n436 10.6151
R693 B.n436 B.n435 10.6151
R694 B.n435 B.n56 10.6151
R695 B.n431 B.n56 10.6151
R696 B.n431 B.n430 10.6151
R697 B.n430 B.n429 10.6151
R698 B.n429 B.n58 10.6151
R699 B.n425 B.n58 10.6151
R700 B.n425 B.n424 10.6151
R701 B.n424 B.n423 10.6151
R702 B.n423 B.n60 10.6151
R703 B.n419 B.n60 10.6151
R704 B.n419 B.n418 10.6151
R705 B.n418 B.n417 10.6151
R706 B.n417 B.n62 10.6151
R707 B.n413 B.n62 10.6151
R708 B.n413 B.n412 10.6151
R709 B.n412 B.n411 10.6151
R710 B.n411 B.n64 10.6151
R711 B.n407 B.n64 10.6151
R712 B.n407 B.n406 10.6151
R713 B.n406 B.n405 10.6151
R714 B.n405 B.n66 10.6151
R715 B.n401 B.n66 10.6151
R716 B.n401 B.n400 10.6151
R717 B.n400 B.n399 10.6151
R718 B.n399 B.n68 10.6151
R719 B.n395 B.n68 10.6151
R720 B.n395 B.n394 10.6151
R721 B.n394 B.n393 10.6151
R722 B.n393 B.n70 10.6151
R723 B.n389 B.n388 10.6151
R724 B.n388 B.n387 10.6151
R725 B.n387 B.n72 10.6151
R726 B.n383 B.n72 10.6151
R727 B.n383 B.n382 10.6151
R728 B.n382 B.n381 10.6151
R729 B.n381 B.n74 10.6151
R730 B.n377 B.n74 10.6151
R731 B.n377 B.n376 10.6151
R732 B.n376 B.n375 10.6151
R733 B.n375 B.n76 10.6151
R734 B.n371 B.n76 10.6151
R735 B.n371 B.n370 10.6151
R736 B.n370 B.n369 10.6151
R737 B.n369 B.n78 10.6151
R738 B.n365 B.n78 10.6151
R739 B.n365 B.n364 10.6151
R740 B.n364 B.n363 10.6151
R741 B.n363 B.n80 10.6151
R742 B.n359 B.n80 10.6151
R743 B.n359 B.n358 10.6151
R744 B.n358 B.n357 10.6151
R745 B.n357 B.n82 10.6151
R746 B.n353 B.n82 10.6151
R747 B.n353 B.n352 10.6151
R748 B.n352 B.n351 10.6151
R749 B.n351 B.n84 10.6151
R750 B.n347 B.n84 10.6151
R751 B.n347 B.n346 10.6151
R752 B.n151 B.n1 10.6151
R753 B.n151 B.n150 10.6151
R754 B.n155 B.n150 10.6151
R755 B.n156 B.n155 10.6151
R756 B.n157 B.n156 10.6151
R757 B.n157 B.n148 10.6151
R758 B.n161 B.n148 10.6151
R759 B.n162 B.n161 10.6151
R760 B.n163 B.n162 10.6151
R761 B.n163 B.n146 10.6151
R762 B.n167 B.n146 10.6151
R763 B.n168 B.n167 10.6151
R764 B.n169 B.n168 10.6151
R765 B.n173 B.n144 10.6151
R766 B.n174 B.n173 10.6151
R767 B.n175 B.n174 10.6151
R768 B.n175 B.n142 10.6151
R769 B.n179 B.n142 10.6151
R770 B.n180 B.n179 10.6151
R771 B.n181 B.n180 10.6151
R772 B.n181 B.n140 10.6151
R773 B.n185 B.n140 10.6151
R774 B.n186 B.n185 10.6151
R775 B.n187 B.n186 10.6151
R776 B.n187 B.n138 10.6151
R777 B.n191 B.n138 10.6151
R778 B.n192 B.n191 10.6151
R779 B.n193 B.n192 10.6151
R780 B.n193 B.n136 10.6151
R781 B.n197 B.n136 10.6151
R782 B.n198 B.n197 10.6151
R783 B.n199 B.n198 10.6151
R784 B.n199 B.n134 10.6151
R785 B.n203 B.n134 10.6151
R786 B.n204 B.n203 10.6151
R787 B.n205 B.n204 10.6151
R788 B.n205 B.n132 10.6151
R789 B.n209 B.n132 10.6151
R790 B.n210 B.n209 10.6151
R791 B.n211 B.n210 10.6151
R792 B.n211 B.n130 10.6151
R793 B.n215 B.n130 10.6151
R794 B.n216 B.n215 10.6151
R795 B.n217 B.n216 10.6151
R796 B.n217 B.n128 10.6151
R797 B.n221 B.n128 10.6151
R798 B.n222 B.n221 10.6151
R799 B.n223 B.n222 10.6151
R800 B.n223 B.n126 10.6151
R801 B.n227 B.n126 10.6151
R802 B.n228 B.n227 10.6151
R803 B.n229 B.n228 10.6151
R804 B.n229 B.n124 10.6151
R805 B.n233 B.n124 10.6151
R806 B.n234 B.n233 10.6151
R807 B.n235 B.n234 10.6151
R808 B.n235 B.n122 10.6151
R809 B.n239 B.n122 10.6151
R810 B.n240 B.n239 10.6151
R811 B.n241 B.n240 10.6151
R812 B.n241 B.n120 10.6151
R813 B.n245 B.n120 10.6151
R814 B.n246 B.n245 10.6151
R815 B.n250 B.n246 10.6151
R816 B.n254 B.n118 10.6151
R817 B.n255 B.n254 10.6151
R818 B.n256 B.n255 10.6151
R819 B.n256 B.n116 10.6151
R820 B.n260 B.n116 10.6151
R821 B.n261 B.n260 10.6151
R822 B.n262 B.n261 10.6151
R823 B.n262 B.n114 10.6151
R824 B.n266 B.n114 10.6151
R825 B.n269 B.n268 10.6151
R826 B.n269 B.n110 10.6151
R827 B.n273 B.n110 10.6151
R828 B.n274 B.n273 10.6151
R829 B.n275 B.n274 10.6151
R830 B.n275 B.n108 10.6151
R831 B.n279 B.n108 10.6151
R832 B.n280 B.n279 10.6151
R833 B.n281 B.n280 10.6151
R834 B.n281 B.n106 10.6151
R835 B.n285 B.n106 10.6151
R836 B.n286 B.n285 10.6151
R837 B.n287 B.n286 10.6151
R838 B.n287 B.n104 10.6151
R839 B.n291 B.n104 10.6151
R840 B.n292 B.n291 10.6151
R841 B.n293 B.n292 10.6151
R842 B.n293 B.n102 10.6151
R843 B.n297 B.n102 10.6151
R844 B.n298 B.n297 10.6151
R845 B.n299 B.n298 10.6151
R846 B.n299 B.n100 10.6151
R847 B.n303 B.n100 10.6151
R848 B.n304 B.n303 10.6151
R849 B.n305 B.n304 10.6151
R850 B.n305 B.n98 10.6151
R851 B.n309 B.n98 10.6151
R852 B.n310 B.n309 10.6151
R853 B.n311 B.n310 10.6151
R854 B.n311 B.n96 10.6151
R855 B.n315 B.n96 10.6151
R856 B.n316 B.n315 10.6151
R857 B.n317 B.n316 10.6151
R858 B.n317 B.n94 10.6151
R859 B.n321 B.n94 10.6151
R860 B.n322 B.n321 10.6151
R861 B.n323 B.n322 10.6151
R862 B.n323 B.n92 10.6151
R863 B.n327 B.n92 10.6151
R864 B.n328 B.n327 10.6151
R865 B.n329 B.n328 10.6151
R866 B.n329 B.n90 10.6151
R867 B.n333 B.n90 10.6151
R868 B.n334 B.n333 10.6151
R869 B.n335 B.n334 10.6151
R870 B.n335 B.n88 10.6151
R871 B.n339 B.n88 10.6151
R872 B.n340 B.n339 10.6151
R873 B.n341 B.n340 10.6151
R874 B.n341 B.n86 10.6151
R875 B.n345 B.n86 10.6151
R876 B.n485 B.n484 9.52245
R877 B.n467 B.n44 9.52245
R878 B.n250 B.n249 9.52245
R879 B.n268 B.n267 9.52245
R880 B.n585 B.n0 8.11757
R881 B.n585 B.n1 8.11757
R882 B.n484 B.n483 1.09318
R883 B.n470 B.n44 1.09318
R884 B.n249 B.n118 1.09318
R885 B.n267 B.n266 1.09318
R886 VN.n0 VN.t0 1008.51
R887 VN.n1 VN.t1 1008.51
R888 VN.n0 VN.t3 1008.48
R889 VN.n1 VN.t2 1008.48
R890 VN VN.n1 112.829
R891 VN VN.n0 70.265
R892 VDD2.n2 VDD2.n0 113.204
R893 VDD2.n2 VDD2.n1 74.1368
R894 VDD2.n1 VDD2.t2 2.08951
R895 VDD2.n1 VDD2.t0 2.08951
R896 VDD2.n0 VDD2.t3 2.08951
R897 VDD2.n0 VDD2.t1 2.08951
R898 VDD2 VDD2.n2 0.0586897
R899 VTAIL.n682 VTAIL.n602 756.745
R900 VTAIL.n80 VTAIL.n0 756.745
R901 VTAIL.n166 VTAIL.n86 756.745
R902 VTAIL.n252 VTAIL.n172 756.745
R903 VTAIL.n596 VTAIL.n516 756.745
R904 VTAIL.n510 VTAIL.n430 756.745
R905 VTAIL.n424 VTAIL.n344 756.745
R906 VTAIL.n338 VTAIL.n258 756.745
R907 VTAIL.n631 VTAIL.n630 585
R908 VTAIL.n633 VTAIL.n632 585
R909 VTAIL.n626 VTAIL.n625 585
R910 VTAIL.n639 VTAIL.n638 585
R911 VTAIL.n641 VTAIL.n640 585
R912 VTAIL.n622 VTAIL.n621 585
R913 VTAIL.n647 VTAIL.n646 585
R914 VTAIL.n649 VTAIL.n648 585
R915 VTAIL.n618 VTAIL.n617 585
R916 VTAIL.n655 VTAIL.n654 585
R917 VTAIL.n657 VTAIL.n656 585
R918 VTAIL.n614 VTAIL.n613 585
R919 VTAIL.n663 VTAIL.n662 585
R920 VTAIL.n665 VTAIL.n664 585
R921 VTAIL.n610 VTAIL.n609 585
R922 VTAIL.n672 VTAIL.n671 585
R923 VTAIL.n673 VTAIL.n608 585
R924 VTAIL.n675 VTAIL.n674 585
R925 VTAIL.n606 VTAIL.n605 585
R926 VTAIL.n681 VTAIL.n680 585
R927 VTAIL.n683 VTAIL.n682 585
R928 VTAIL.n29 VTAIL.n28 585
R929 VTAIL.n31 VTAIL.n30 585
R930 VTAIL.n24 VTAIL.n23 585
R931 VTAIL.n37 VTAIL.n36 585
R932 VTAIL.n39 VTAIL.n38 585
R933 VTAIL.n20 VTAIL.n19 585
R934 VTAIL.n45 VTAIL.n44 585
R935 VTAIL.n47 VTAIL.n46 585
R936 VTAIL.n16 VTAIL.n15 585
R937 VTAIL.n53 VTAIL.n52 585
R938 VTAIL.n55 VTAIL.n54 585
R939 VTAIL.n12 VTAIL.n11 585
R940 VTAIL.n61 VTAIL.n60 585
R941 VTAIL.n63 VTAIL.n62 585
R942 VTAIL.n8 VTAIL.n7 585
R943 VTAIL.n70 VTAIL.n69 585
R944 VTAIL.n71 VTAIL.n6 585
R945 VTAIL.n73 VTAIL.n72 585
R946 VTAIL.n4 VTAIL.n3 585
R947 VTAIL.n79 VTAIL.n78 585
R948 VTAIL.n81 VTAIL.n80 585
R949 VTAIL.n115 VTAIL.n114 585
R950 VTAIL.n117 VTAIL.n116 585
R951 VTAIL.n110 VTAIL.n109 585
R952 VTAIL.n123 VTAIL.n122 585
R953 VTAIL.n125 VTAIL.n124 585
R954 VTAIL.n106 VTAIL.n105 585
R955 VTAIL.n131 VTAIL.n130 585
R956 VTAIL.n133 VTAIL.n132 585
R957 VTAIL.n102 VTAIL.n101 585
R958 VTAIL.n139 VTAIL.n138 585
R959 VTAIL.n141 VTAIL.n140 585
R960 VTAIL.n98 VTAIL.n97 585
R961 VTAIL.n147 VTAIL.n146 585
R962 VTAIL.n149 VTAIL.n148 585
R963 VTAIL.n94 VTAIL.n93 585
R964 VTAIL.n156 VTAIL.n155 585
R965 VTAIL.n157 VTAIL.n92 585
R966 VTAIL.n159 VTAIL.n158 585
R967 VTAIL.n90 VTAIL.n89 585
R968 VTAIL.n165 VTAIL.n164 585
R969 VTAIL.n167 VTAIL.n166 585
R970 VTAIL.n201 VTAIL.n200 585
R971 VTAIL.n203 VTAIL.n202 585
R972 VTAIL.n196 VTAIL.n195 585
R973 VTAIL.n209 VTAIL.n208 585
R974 VTAIL.n211 VTAIL.n210 585
R975 VTAIL.n192 VTAIL.n191 585
R976 VTAIL.n217 VTAIL.n216 585
R977 VTAIL.n219 VTAIL.n218 585
R978 VTAIL.n188 VTAIL.n187 585
R979 VTAIL.n225 VTAIL.n224 585
R980 VTAIL.n227 VTAIL.n226 585
R981 VTAIL.n184 VTAIL.n183 585
R982 VTAIL.n233 VTAIL.n232 585
R983 VTAIL.n235 VTAIL.n234 585
R984 VTAIL.n180 VTAIL.n179 585
R985 VTAIL.n242 VTAIL.n241 585
R986 VTAIL.n243 VTAIL.n178 585
R987 VTAIL.n245 VTAIL.n244 585
R988 VTAIL.n176 VTAIL.n175 585
R989 VTAIL.n251 VTAIL.n250 585
R990 VTAIL.n253 VTAIL.n252 585
R991 VTAIL.n597 VTAIL.n596 585
R992 VTAIL.n595 VTAIL.n594 585
R993 VTAIL.n520 VTAIL.n519 585
R994 VTAIL.n524 VTAIL.n522 585
R995 VTAIL.n589 VTAIL.n588 585
R996 VTAIL.n587 VTAIL.n586 585
R997 VTAIL.n526 VTAIL.n525 585
R998 VTAIL.n581 VTAIL.n580 585
R999 VTAIL.n579 VTAIL.n578 585
R1000 VTAIL.n530 VTAIL.n529 585
R1001 VTAIL.n573 VTAIL.n572 585
R1002 VTAIL.n571 VTAIL.n570 585
R1003 VTAIL.n534 VTAIL.n533 585
R1004 VTAIL.n565 VTAIL.n564 585
R1005 VTAIL.n563 VTAIL.n562 585
R1006 VTAIL.n538 VTAIL.n537 585
R1007 VTAIL.n557 VTAIL.n556 585
R1008 VTAIL.n555 VTAIL.n554 585
R1009 VTAIL.n542 VTAIL.n541 585
R1010 VTAIL.n549 VTAIL.n548 585
R1011 VTAIL.n547 VTAIL.n546 585
R1012 VTAIL.n511 VTAIL.n510 585
R1013 VTAIL.n509 VTAIL.n508 585
R1014 VTAIL.n434 VTAIL.n433 585
R1015 VTAIL.n438 VTAIL.n436 585
R1016 VTAIL.n503 VTAIL.n502 585
R1017 VTAIL.n501 VTAIL.n500 585
R1018 VTAIL.n440 VTAIL.n439 585
R1019 VTAIL.n495 VTAIL.n494 585
R1020 VTAIL.n493 VTAIL.n492 585
R1021 VTAIL.n444 VTAIL.n443 585
R1022 VTAIL.n487 VTAIL.n486 585
R1023 VTAIL.n485 VTAIL.n484 585
R1024 VTAIL.n448 VTAIL.n447 585
R1025 VTAIL.n479 VTAIL.n478 585
R1026 VTAIL.n477 VTAIL.n476 585
R1027 VTAIL.n452 VTAIL.n451 585
R1028 VTAIL.n471 VTAIL.n470 585
R1029 VTAIL.n469 VTAIL.n468 585
R1030 VTAIL.n456 VTAIL.n455 585
R1031 VTAIL.n463 VTAIL.n462 585
R1032 VTAIL.n461 VTAIL.n460 585
R1033 VTAIL.n425 VTAIL.n424 585
R1034 VTAIL.n423 VTAIL.n422 585
R1035 VTAIL.n348 VTAIL.n347 585
R1036 VTAIL.n352 VTAIL.n350 585
R1037 VTAIL.n417 VTAIL.n416 585
R1038 VTAIL.n415 VTAIL.n414 585
R1039 VTAIL.n354 VTAIL.n353 585
R1040 VTAIL.n409 VTAIL.n408 585
R1041 VTAIL.n407 VTAIL.n406 585
R1042 VTAIL.n358 VTAIL.n357 585
R1043 VTAIL.n401 VTAIL.n400 585
R1044 VTAIL.n399 VTAIL.n398 585
R1045 VTAIL.n362 VTAIL.n361 585
R1046 VTAIL.n393 VTAIL.n392 585
R1047 VTAIL.n391 VTAIL.n390 585
R1048 VTAIL.n366 VTAIL.n365 585
R1049 VTAIL.n385 VTAIL.n384 585
R1050 VTAIL.n383 VTAIL.n382 585
R1051 VTAIL.n370 VTAIL.n369 585
R1052 VTAIL.n377 VTAIL.n376 585
R1053 VTAIL.n375 VTAIL.n374 585
R1054 VTAIL.n339 VTAIL.n338 585
R1055 VTAIL.n337 VTAIL.n336 585
R1056 VTAIL.n262 VTAIL.n261 585
R1057 VTAIL.n266 VTAIL.n264 585
R1058 VTAIL.n331 VTAIL.n330 585
R1059 VTAIL.n329 VTAIL.n328 585
R1060 VTAIL.n268 VTAIL.n267 585
R1061 VTAIL.n323 VTAIL.n322 585
R1062 VTAIL.n321 VTAIL.n320 585
R1063 VTAIL.n272 VTAIL.n271 585
R1064 VTAIL.n315 VTAIL.n314 585
R1065 VTAIL.n313 VTAIL.n312 585
R1066 VTAIL.n276 VTAIL.n275 585
R1067 VTAIL.n307 VTAIL.n306 585
R1068 VTAIL.n305 VTAIL.n304 585
R1069 VTAIL.n280 VTAIL.n279 585
R1070 VTAIL.n299 VTAIL.n298 585
R1071 VTAIL.n297 VTAIL.n296 585
R1072 VTAIL.n284 VTAIL.n283 585
R1073 VTAIL.n291 VTAIL.n290 585
R1074 VTAIL.n289 VTAIL.n288 585
R1075 VTAIL.n629 VTAIL.t4 327.466
R1076 VTAIL.n27 VTAIL.t7 327.466
R1077 VTAIL.n113 VTAIL.t3 327.466
R1078 VTAIL.n199 VTAIL.t2 327.466
R1079 VTAIL.n545 VTAIL.t0 327.466
R1080 VTAIL.n459 VTAIL.t1 327.466
R1081 VTAIL.n373 VTAIL.t6 327.466
R1082 VTAIL.n287 VTAIL.t5 327.466
R1083 VTAIL.n632 VTAIL.n631 171.744
R1084 VTAIL.n632 VTAIL.n625 171.744
R1085 VTAIL.n639 VTAIL.n625 171.744
R1086 VTAIL.n640 VTAIL.n639 171.744
R1087 VTAIL.n640 VTAIL.n621 171.744
R1088 VTAIL.n647 VTAIL.n621 171.744
R1089 VTAIL.n648 VTAIL.n647 171.744
R1090 VTAIL.n648 VTAIL.n617 171.744
R1091 VTAIL.n655 VTAIL.n617 171.744
R1092 VTAIL.n656 VTAIL.n655 171.744
R1093 VTAIL.n656 VTAIL.n613 171.744
R1094 VTAIL.n663 VTAIL.n613 171.744
R1095 VTAIL.n664 VTAIL.n663 171.744
R1096 VTAIL.n664 VTAIL.n609 171.744
R1097 VTAIL.n672 VTAIL.n609 171.744
R1098 VTAIL.n673 VTAIL.n672 171.744
R1099 VTAIL.n674 VTAIL.n673 171.744
R1100 VTAIL.n674 VTAIL.n605 171.744
R1101 VTAIL.n681 VTAIL.n605 171.744
R1102 VTAIL.n682 VTAIL.n681 171.744
R1103 VTAIL.n30 VTAIL.n29 171.744
R1104 VTAIL.n30 VTAIL.n23 171.744
R1105 VTAIL.n37 VTAIL.n23 171.744
R1106 VTAIL.n38 VTAIL.n37 171.744
R1107 VTAIL.n38 VTAIL.n19 171.744
R1108 VTAIL.n45 VTAIL.n19 171.744
R1109 VTAIL.n46 VTAIL.n45 171.744
R1110 VTAIL.n46 VTAIL.n15 171.744
R1111 VTAIL.n53 VTAIL.n15 171.744
R1112 VTAIL.n54 VTAIL.n53 171.744
R1113 VTAIL.n54 VTAIL.n11 171.744
R1114 VTAIL.n61 VTAIL.n11 171.744
R1115 VTAIL.n62 VTAIL.n61 171.744
R1116 VTAIL.n62 VTAIL.n7 171.744
R1117 VTAIL.n70 VTAIL.n7 171.744
R1118 VTAIL.n71 VTAIL.n70 171.744
R1119 VTAIL.n72 VTAIL.n71 171.744
R1120 VTAIL.n72 VTAIL.n3 171.744
R1121 VTAIL.n79 VTAIL.n3 171.744
R1122 VTAIL.n80 VTAIL.n79 171.744
R1123 VTAIL.n116 VTAIL.n115 171.744
R1124 VTAIL.n116 VTAIL.n109 171.744
R1125 VTAIL.n123 VTAIL.n109 171.744
R1126 VTAIL.n124 VTAIL.n123 171.744
R1127 VTAIL.n124 VTAIL.n105 171.744
R1128 VTAIL.n131 VTAIL.n105 171.744
R1129 VTAIL.n132 VTAIL.n131 171.744
R1130 VTAIL.n132 VTAIL.n101 171.744
R1131 VTAIL.n139 VTAIL.n101 171.744
R1132 VTAIL.n140 VTAIL.n139 171.744
R1133 VTAIL.n140 VTAIL.n97 171.744
R1134 VTAIL.n147 VTAIL.n97 171.744
R1135 VTAIL.n148 VTAIL.n147 171.744
R1136 VTAIL.n148 VTAIL.n93 171.744
R1137 VTAIL.n156 VTAIL.n93 171.744
R1138 VTAIL.n157 VTAIL.n156 171.744
R1139 VTAIL.n158 VTAIL.n157 171.744
R1140 VTAIL.n158 VTAIL.n89 171.744
R1141 VTAIL.n165 VTAIL.n89 171.744
R1142 VTAIL.n166 VTAIL.n165 171.744
R1143 VTAIL.n202 VTAIL.n201 171.744
R1144 VTAIL.n202 VTAIL.n195 171.744
R1145 VTAIL.n209 VTAIL.n195 171.744
R1146 VTAIL.n210 VTAIL.n209 171.744
R1147 VTAIL.n210 VTAIL.n191 171.744
R1148 VTAIL.n217 VTAIL.n191 171.744
R1149 VTAIL.n218 VTAIL.n217 171.744
R1150 VTAIL.n218 VTAIL.n187 171.744
R1151 VTAIL.n225 VTAIL.n187 171.744
R1152 VTAIL.n226 VTAIL.n225 171.744
R1153 VTAIL.n226 VTAIL.n183 171.744
R1154 VTAIL.n233 VTAIL.n183 171.744
R1155 VTAIL.n234 VTAIL.n233 171.744
R1156 VTAIL.n234 VTAIL.n179 171.744
R1157 VTAIL.n242 VTAIL.n179 171.744
R1158 VTAIL.n243 VTAIL.n242 171.744
R1159 VTAIL.n244 VTAIL.n243 171.744
R1160 VTAIL.n244 VTAIL.n175 171.744
R1161 VTAIL.n251 VTAIL.n175 171.744
R1162 VTAIL.n252 VTAIL.n251 171.744
R1163 VTAIL.n596 VTAIL.n595 171.744
R1164 VTAIL.n595 VTAIL.n519 171.744
R1165 VTAIL.n524 VTAIL.n519 171.744
R1166 VTAIL.n588 VTAIL.n524 171.744
R1167 VTAIL.n588 VTAIL.n587 171.744
R1168 VTAIL.n587 VTAIL.n525 171.744
R1169 VTAIL.n580 VTAIL.n525 171.744
R1170 VTAIL.n580 VTAIL.n579 171.744
R1171 VTAIL.n579 VTAIL.n529 171.744
R1172 VTAIL.n572 VTAIL.n529 171.744
R1173 VTAIL.n572 VTAIL.n571 171.744
R1174 VTAIL.n571 VTAIL.n533 171.744
R1175 VTAIL.n564 VTAIL.n533 171.744
R1176 VTAIL.n564 VTAIL.n563 171.744
R1177 VTAIL.n563 VTAIL.n537 171.744
R1178 VTAIL.n556 VTAIL.n537 171.744
R1179 VTAIL.n556 VTAIL.n555 171.744
R1180 VTAIL.n555 VTAIL.n541 171.744
R1181 VTAIL.n548 VTAIL.n541 171.744
R1182 VTAIL.n548 VTAIL.n547 171.744
R1183 VTAIL.n510 VTAIL.n509 171.744
R1184 VTAIL.n509 VTAIL.n433 171.744
R1185 VTAIL.n438 VTAIL.n433 171.744
R1186 VTAIL.n502 VTAIL.n438 171.744
R1187 VTAIL.n502 VTAIL.n501 171.744
R1188 VTAIL.n501 VTAIL.n439 171.744
R1189 VTAIL.n494 VTAIL.n439 171.744
R1190 VTAIL.n494 VTAIL.n493 171.744
R1191 VTAIL.n493 VTAIL.n443 171.744
R1192 VTAIL.n486 VTAIL.n443 171.744
R1193 VTAIL.n486 VTAIL.n485 171.744
R1194 VTAIL.n485 VTAIL.n447 171.744
R1195 VTAIL.n478 VTAIL.n447 171.744
R1196 VTAIL.n478 VTAIL.n477 171.744
R1197 VTAIL.n477 VTAIL.n451 171.744
R1198 VTAIL.n470 VTAIL.n451 171.744
R1199 VTAIL.n470 VTAIL.n469 171.744
R1200 VTAIL.n469 VTAIL.n455 171.744
R1201 VTAIL.n462 VTAIL.n455 171.744
R1202 VTAIL.n462 VTAIL.n461 171.744
R1203 VTAIL.n424 VTAIL.n423 171.744
R1204 VTAIL.n423 VTAIL.n347 171.744
R1205 VTAIL.n352 VTAIL.n347 171.744
R1206 VTAIL.n416 VTAIL.n352 171.744
R1207 VTAIL.n416 VTAIL.n415 171.744
R1208 VTAIL.n415 VTAIL.n353 171.744
R1209 VTAIL.n408 VTAIL.n353 171.744
R1210 VTAIL.n408 VTAIL.n407 171.744
R1211 VTAIL.n407 VTAIL.n357 171.744
R1212 VTAIL.n400 VTAIL.n357 171.744
R1213 VTAIL.n400 VTAIL.n399 171.744
R1214 VTAIL.n399 VTAIL.n361 171.744
R1215 VTAIL.n392 VTAIL.n361 171.744
R1216 VTAIL.n392 VTAIL.n391 171.744
R1217 VTAIL.n391 VTAIL.n365 171.744
R1218 VTAIL.n384 VTAIL.n365 171.744
R1219 VTAIL.n384 VTAIL.n383 171.744
R1220 VTAIL.n383 VTAIL.n369 171.744
R1221 VTAIL.n376 VTAIL.n369 171.744
R1222 VTAIL.n376 VTAIL.n375 171.744
R1223 VTAIL.n338 VTAIL.n337 171.744
R1224 VTAIL.n337 VTAIL.n261 171.744
R1225 VTAIL.n266 VTAIL.n261 171.744
R1226 VTAIL.n330 VTAIL.n266 171.744
R1227 VTAIL.n330 VTAIL.n329 171.744
R1228 VTAIL.n329 VTAIL.n267 171.744
R1229 VTAIL.n322 VTAIL.n267 171.744
R1230 VTAIL.n322 VTAIL.n321 171.744
R1231 VTAIL.n321 VTAIL.n271 171.744
R1232 VTAIL.n314 VTAIL.n271 171.744
R1233 VTAIL.n314 VTAIL.n313 171.744
R1234 VTAIL.n313 VTAIL.n275 171.744
R1235 VTAIL.n306 VTAIL.n275 171.744
R1236 VTAIL.n306 VTAIL.n305 171.744
R1237 VTAIL.n305 VTAIL.n279 171.744
R1238 VTAIL.n298 VTAIL.n279 171.744
R1239 VTAIL.n298 VTAIL.n297 171.744
R1240 VTAIL.n297 VTAIL.n283 171.744
R1241 VTAIL.n290 VTAIL.n283 171.744
R1242 VTAIL.n290 VTAIL.n289 171.744
R1243 VTAIL.n631 VTAIL.t4 85.8723
R1244 VTAIL.n29 VTAIL.t7 85.8723
R1245 VTAIL.n115 VTAIL.t3 85.8723
R1246 VTAIL.n201 VTAIL.t2 85.8723
R1247 VTAIL.n547 VTAIL.t0 85.8723
R1248 VTAIL.n461 VTAIL.t1 85.8723
R1249 VTAIL.n375 VTAIL.t6 85.8723
R1250 VTAIL.n289 VTAIL.t5 85.8723
R1251 VTAIL.n687 VTAIL.n686 36.0641
R1252 VTAIL.n85 VTAIL.n84 36.0641
R1253 VTAIL.n171 VTAIL.n170 36.0641
R1254 VTAIL.n257 VTAIL.n256 36.0641
R1255 VTAIL.n601 VTAIL.n600 36.0641
R1256 VTAIL.n515 VTAIL.n514 36.0641
R1257 VTAIL.n429 VTAIL.n428 36.0641
R1258 VTAIL.n343 VTAIL.n342 36.0641
R1259 VTAIL.n687 VTAIL.n601 26.4272
R1260 VTAIL.n343 VTAIL.n257 26.4272
R1261 VTAIL.n630 VTAIL.n629 16.3895
R1262 VTAIL.n28 VTAIL.n27 16.3895
R1263 VTAIL.n114 VTAIL.n113 16.3895
R1264 VTAIL.n200 VTAIL.n199 16.3895
R1265 VTAIL.n546 VTAIL.n545 16.3895
R1266 VTAIL.n460 VTAIL.n459 16.3895
R1267 VTAIL.n374 VTAIL.n373 16.3895
R1268 VTAIL.n288 VTAIL.n287 16.3895
R1269 VTAIL.n675 VTAIL.n606 13.1884
R1270 VTAIL.n73 VTAIL.n4 13.1884
R1271 VTAIL.n159 VTAIL.n90 13.1884
R1272 VTAIL.n245 VTAIL.n176 13.1884
R1273 VTAIL.n522 VTAIL.n520 13.1884
R1274 VTAIL.n436 VTAIL.n434 13.1884
R1275 VTAIL.n350 VTAIL.n348 13.1884
R1276 VTAIL.n264 VTAIL.n262 13.1884
R1277 VTAIL.n633 VTAIL.n628 12.8005
R1278 VTAIL.n676 VTAIL.n608 12.8005
R1279 VTAIL.n680 VTAIL.n679 12.8005
R1280 VTAIL.n31 VTAIL.n26 12.8005
R1281 VTAIL.n74 VTAIL.n6 12.8005
R1282 VTAIL.n78 VTAIL.n77 12.8005
R1283 VTAIL.n117 VTAIL.n112 12.8005
R1284 VTAIL.n160 VTAIL.n92 12.8005
R1285 VTAIL.n164 VTAIL.n163 12.8005
R1286 VTAIL.n203 VTAIL.n198 12.8005
R1287 VTAIL.n246 VTAIL.n178 12.8005
R1288 VTAIL.n250 VTAIL.n249 12.8005
R1289 VTAIL.n594 VTAIL.n593 12.8005
R1290 VTAIL.n590 VTAIL.n589 12.8005
R1291 VTAIL.n549 VTAIL.n544 12.8005
R1292 VTAIL.n508 VTAIL.n507 12.8005
R1293 VTAIL.n504 VTAIL.n503 12.8005
R1294 VTAIL.n463 VTAIL.n458 12.8005
R1295 VTAIL.n422 VTAIL.n421 12.8005
R1296 VTAIL.n418 VTAIL.n417 12.8005
R1297 VTAIL.n377 VTAIL.n372 12.8005
R1298 VTAIL.n336 VTAIL.n335 12.8005
R1299 VTAIL.n332 VTAIL.n331 12.8005
R1300 VTAIL.n291 VTAIL.n286 12.8005
R1301 VTAIL.n634 VTAIL.n626 12.0247
R1302 VTAIL.n671 VTAIL.n670 12.0247
R1303 VTAIL.n683 VTAIL.n604 12.0247
R1304 VTAIL.n32 VTAIL.n24 12.0247
R1305 VTAIL.n69 VTAIL.n68 12.0247
R1306 VTAIL.n81 VTAIL.n2 12.0247
R1307 VTAIL.n118 VTAIL.n110 12.0247
R1308 VTAIL.n155 VTAIL.n154 12.0247
R1309 VTAIL.n167 VTAIL.n88 12.0247
R1310 VTAIL.n204 VTAIL.n196 12.0247
R1311 VTAIL.n241 VTAIL.n240 12.0247
R1312 VTAIL.n253 VTAIL.n174 12.0247
R1313 VTAIL.n597 VTAIL.n518 12.0247
R1314 VTAIL.n586 VTAIL.n523 12.0247
R1315 VTAIL.n550 VTAIL.n542 12.0247
R1316 VTAIL.n511 VTAIL.n432 12.0247
R1317 VTAIL.n500 VTAIL.n437 12.0247
R1318 VTAIL.n464 VTAIL.n456 12.0247
R1319 VTAIL.n425 VTAIL.n346 12.0247
R1320 VTAIL.n414 VTAIL.n351 12.0247
R1321 VTAIL.n378 VTAIL.n370 12.0247
R1322 VTAIL.n339 VTAIL.n260 12.0247
R1323 VTAIL.n328 VTAIL.n265 12.0247
R1324 VTAIL.n292 VTAIL.n284 12.0247
R1325 VTAIL.n638 VTAIL.n637 11.249
R1326 VTAIL.n669 VTAIL.n610 11.249
R1327 VTAIL.n684 VTAIL.n602 11.249
R1328 VTAIL.n36 VTAIL.n35 11.249
R1329 VTAIL.n67 VTAIL.n8 11.249
R1330 VTAIL.n82 VTAIL.n0 11.249
R1331 VTAIL.n122 VTAIL.n121 11.249
R1332 VTAIL.n153 VTAIL.n94 11.249
R1333 VTAIL.n168 VTAIL.n86 11.249
R1334 VTAIL.n208 VTAIL.n207 11.249
R1335 VTAIL.n239 VTAIL.n180 11.249
R1336 VTAIL.n254 VTAIL.n172 11.249
R1337 VTAIL.n598 VTAIL.n516 11.249
R1338 VTAIL.n585 VTAIL.n526 11.249
R1339 VTAIL.n554 VTAIL.n553 11.249
R1340 VTAIL.n512 VTAIL.n430 11.249
R1341 VTAIL.n499 VTAIL.n440 11.249
R1342 VTAIL.n468 VTAIL.n467 11.249
R1343 VTAIL.n426 VTAIL.n344 11.249
R1344 VTAIL.n413 VTAIL.n354 11.249
R1345 VTAIL.n382 VTAIL.n381 11.249
R1346 VTAIL.n340 VTAIL.n258 11.249
R1347 VTAIL.n327 VTAIL.n268 11.249
R1348 VTAIL.n296 VTAIL.n295 11.249
R1349 VTAIL.n641 VTAIL.n624 10.4732
R1350 VTAIL.n666 VTAIL.n665 10.4732
R1351 VTAIL.n39 VTAIL.n22 10.4732
R1352 VTAIL.n64 VTAIL.n63 10.4732
R1353 VTAIL.n125 VTAIL.n108 10.4732
R1354 VTAIL.n150 VTAIL.n149 10.4732
R1355 VTAIL.n211 VTAIL.n194 10.4732
R1356 VTAIL.n236 VTAIL.n235 10.4732
R1357 VTAIL.n582 VTAIL.n581 10.4732
R1358 VTAIL.n557 VTAIL.n540 10.4732
R1359 VTAIL.n496 VTAIL.n495 10.4732
R1360 VTAIL.n471 VTAIL.n454 10.4732
R1361 VTAIL.n410 VTAIL.n409 10.4732
R1362 VTAIL.n385 VTAIL.n368 10.4732
R1363 VTAIL.n324 VTAIL.n323 10.4732
R1364 VTAIL.n299 VTAIL.n282 10.4732
R1365 VTAIL.n642 VTAIL.n622 9.69747
R1366 VTAIL.n662 VTAIL.n612 9.69747
R1367 VTAIL.n40 VTAIL.n20 9.69747
R1368 VTAIL.n60 VTAIL.n10 9.69747
R1369 VTAIL.n126 VTAIL.n106 9.69747
R1370 VTAIL.n146 VTAIL.n96 9.69747
R1371 VTAIL.n212 VTAIL.n192 9.69747
R1372 VTAIL.n232 VTAIL.n182 9.69747
R1373 VTAIL.n578 VTAIL.n528 9.69747
R1374 VTAIL.n558 VTAIL.n538 9.69747
R1375 VTAIL.n492 VTAIL.n442 9.69747
R1376 VTAIL.n472 VTAIL.n452 9.69747
R1377 VTAIL.n406 VTAIL.n356 9.69747
R1378 VTAIL.n386 VTAIL.n366 9.69747
R1379 VTAIL.n320 VTAIL.n270 9.69747
R1380 VTAIL.n300 VTAIL.n280 9.69747
R1381 VTAIL.n686 VTAIL.n685 9.45567
R1382 VTAIL.n84 VTAIL.n83 9.45567
R1383 VTAIL.n170 VTAIL.n169 9.45567
R1384 VTAIL.n256 VTAIL.n255 9.45567
R1385 VTAIL.n600 VTAIL.n599 9.45567
R1386 VTAIL.n514 VTAIL.n513 9.45567
R1387 VTAIL.n428 VTAIL.n427 9.45567
R1388 VTAIL.n342 VTAIL.n341 9.45567
R1389 VTAIL.n685 VTAIL.n684 9.3005
R1390 VTAIL.n604 VTAIL.n603 9.3005
R1391 VTAIL.n679 VTAIL.n678 9.3005
R1392 VTAIL.n651 VTAIL.n650 9.3005
R1393 VTAIL.n620 VTAIL.n619 9.3005
R1394 VTAIL.n645 VTAIL.n644 9.3005
R1395 VTAIL.n643 VTAIL.n642 9.3005
R1396 VTAIL.n624 VTAIL.n623 9.3005
R1397 VTAIL.n637 VTAIL.n636 9.3005
R1398 VTAIL.n635 VTAIL.n634 9.3005
R1399 VTAIL.n628 VTAIL.n627 9.3005
R1400 VTAIL.n653 VTAIL.n652 9.3005
R1401 VTAIL.n616 VTAIL.n615 9.3005
R1402 VTAIL.n659 VTAIL.n658 9.3005
R1403 VTAIL.n661 VTAIL.n660 9.3005
R1404 VTAIL.n612 VTAIL.n611 9.3005
R1405 VTAIL.n667 VTAIL.n666 9.3005
R1406 VTAIL.n669 VTAIL.n668 9.3005
R1407 VTAIL.n670 VTAIL.n607 9.3005
R1408 VTAIL.n677 VTAIL.n676 9.3005
R1409 VTAIL.n83 VTAIL.n82 9.3005
R1410 VTAIL.n2 VTAIL.n1 9.3005
R1411 VTAIL.n77 VTAIL.n76 9.3005
R1412 VTAIL.n49 VTAIL.n48 9.3005
R1413 VTAIL.n18 VTAIL.n17 9.3005
R1414 VTAIL.n43 VTAIL.n42 9.3005
R1415 VTAIL.n41 VTAIL.n40 9.3005
R1416 VTAIL.n22 VTAIL.n21 9.3005
R1417 VTAIL.n35 VTAIL.n34 9.3005
R1418 VTAIL.n33 VTAIL.n32 9.3005
R1419 VTAIL.n26 VTAIL.n25 9.3005
R1420 VTAIL.n51 VTAIL.n50 9.3005
R1421 VTAIL.n14 VTAIL.n13 9.3005
R1422 VTAIL.n57 VTAIL.n56 9.3005
R1423 VTAIL.n59 VTAIL.n58 9.3005
R1424 VTAIL.n10 VTAIL.n9 9.3005
R1425 VTAIL.n65 VTAIL.n64 9.3005
R1426 VTAIL.n67 VTAIL.n66 9.3005
R1427 VTAIL.n68 VTAIL.n5 9.3005
R1428 VTAIL.n75 VTAIL.n74 9.3005
R1429 VTAIL.n169 VTAIL.n168 9.3005
R1430 VTAIL.n88 VTAIL.n87 9.3005
R1431 VTAIL.n163 VTAIL.n162 9.3005
R1432 VTAIL.n135 VTAIL.n134 9.3005
R1433 VTAIL.n104 VTAIL.n103 9.3005
R1434 VTAIL.n129 VTAIL.n128 9.3005
R1435 VTAIL.n127 VTAIL.n126 9.3005
R1436 VTAIL.n108 VTAIL.n107 9.3005
R1437 VTAIL.n121 VTAIL.n120 9.3005
R1438 VTAIL.n119 VTAIL.n118 9.3005
R1439 VTAIL.n112 VTAIL.n111 9.3005
R1440 VTAIL.n137 VTAIL.n136 9.3005
R1441 VTAIL.n100 VTAIL.n99 9.3005
R1442 VTAIL.n143 VTAIL.n142 9.3005
R1443 VTAIL.n145 VTAIL.n144 9.3005
R1444 VTAIL.n96 VTAIL.n95 9.3005
R1445 VTAIL.n151 VTAIL.n150 9.3005
R1446 VTAIL.n153 VTAIL.n152 9.3005
R1447 VTAIL.n154 VTAIL.n91 9.3005
R1448 VTAIL.n161 VTAIL.n160 9.3005
R1449 VTAIL.n255 VTAIL.n254 9.3005
R1450 VTAIL.n174 VTAIL.n173 9.3005
R1451 VTAIL.n249 VTAIL.n248 9.3005
R1452 VTAIL.n221 VTAIL.n220 9.3005
R1453 VTAIL.n190 VTAIL.n189 9.3005
R1454 VTAIL.n215 VTAIL.n214 9.3005
R1455 VTAIL.n213 VTAIL.n212 9.3005
R1456 VTAIL.n194 VTAIL.n193 9.3005
R1457 VTAIL.n207 VTAIL.n206 9.3005
R1458 VTAIL.n205 VTAIL.n204 9.3005
R1459 VTAIL.n198 VTAIL.n197 9.3005
R1460 VTAIL.n223 VTAIL.n222 9.3005
R1461 VTAIL.n186 VTAIL.n185 9.3005
R1462 VTAIL.n229 VTAIL.n228 9.3005
R1463 VTAIL.n231 VTAIL.n230 9.3005
R1464 VTAIL.n182 VTAIL.n181 9.3005
R1465 VTAIL.n237 VTAIL.n236 9.3005
R1466 VTAIL.n239 VTAIL.n238 9.3005
R1467 VTAIL.n240 VTAIL.n177 9.3005
R1468 VTAIL.n247 VTAIL.n246 9.3005
R1469 VTAIL.n532 VTAIL.n531 9.3005
R1470 VTAIL.n575 VTAIL.n574 9.3005
R1471 VTAIL.n577 VTAIL.n576 9.3005
R1472 VTAIL.n528 VTAIL.n527 9.3005
R1473 VTAIL.n583 VTAIL.n582 9.3005
R1474 VTAIL.n585 VTAIL.n584 9.3005
R1475 VTAIL.n523 VTAIL.n521 9.3005
R1476 VTAIL.n591 VTAIL.n590 9.3005
R1477 VTAIL.n599 VTAIL.n598 9.3005
R1478 VTAIL.n518 VTAIL.n517 9.3005
R1479 VTAIL.n593 VTAIL.n592 9.3005
R1480 VTAIL.n569 VTAIL.n568 9.3005
R1481 VTAIL.n567 VTAIL.n566 9.3005
R1482 VTAIL.n536 VTAIL.n535 9.3005
R1483 VTAIL.n561 VTAIL.n560 9.3005
R1484 VTAIL.n559 VTAIL.n558 9.3005
R1485 VTAIL.n540 VTAIL.n539 9.3005
R1486 VTAIL.n553 VTAIL.n552 9.3005
R1487 VTAIL.n551 VTAIL.n550 9.3005
R1488 VTAIL.n544 VTAIL.n543 9.3005
R1489 VTAIL.n446 VTAIL.n445 9.3005
R1490 VTAIL.n489 VTAIL.n488 9.3005
R1491 VTAIL.n491 VTAIL.n490 9.3005
R1492 VTAIL.n442 VTAIL.n441 9.3005
R1493 VTAIL.n497 VTAIL.n496 9.3005
R1494 VTAIL.n499 VTAIL.n498 9.3005
R1495 VTAIL.n437 VTAIL.n435 9.3005
R1496 VTAIL.n505 VTAIL.n504 9.3005
R1497 VTAIL.n513 VTAIL.n512 9.3005
R1498 VTAIL.n432 VTAIL.n431 9.3005
R1499 VTAIL.n507 VTAIL.n506 9.3005
R1500 VTAIL.n483 VTAIL.n482 9.3005
R1501 VTAIL.n481 VTAIL.n480 9.3005
R1502 VTAIL.n450 VTAIL.n449 9.3005
R1503 VTAIL.n475 VTAIL.n474 9.3005
R1504 VTAIL.n473 VTAIL.n472 9.3005
R1505 VTAIL.n454 VTAIL.n453 9.3005
R1506 VTAIL.n467 VTAIL.n466 9.3005
R1507 VTAIL.n465 VTAIL.n464 9.3005
R1508 VTAIL.n458 VTAIL.n457 9.3005
R1509 VTAIL.n360 VTAIL.n359 9.3005
R1510 VTAIL.n403 VTAIL.n402 9.3005
R1511 VTAIL.n405 VTAIL.n404 9.3005
R1512 VTAIL.n356 VTAIL.n355 9.3005
R1513 VTAIL.n411 VTAIL.n410 9.3005
R1514 VTAIL.n413 VTAIL.n412 9.3005
R1515 VTAIL.n351 VTAIL.n349 9.3005
R1516 VTAIL.n419 VTAIL.n418 9.3005
R1517 VTAIL.n427 VTAIL.n426 9.3005
R1518 VTAIL.n346 VTAIL.n345 9.3005
R1519 VTAIL.n421 VTAIL.n420 9.3005
R1520 VTAIL.n397 VTAIL.n396 9.3005
R1521 VTAIL.n395 VTAIL.n394 9.3005
R1522 VTAIL.n364 VTAIL.n363 9.3005
R1523 VTAIL.n389 VTAIL.n388 9.3005
R1524 VTAIL.n387 VTAIL.n386 9.3005
R1525 VTAIL.n368 VTAIL.n367 9.3005
R1526 VTAIL.n381 VTAIL.n380 9.3005
R1527 VTAIL.n379 VTAIL.n378 9.3005
R1528 VTAIL.n372 VTAIL.n371 9.3005
R1529 VTAIL.n274 VTAIL.n273 9.3005
R1530 VTAIL.n317 VTAIL.n316 9.3005
R1531 VTAIL.n319 VTAIL.n318 9.3005
R1532 VTAIL.n270 VTAIL.n269 9.3005
R1533 VTAIL.n325 VTAIL.n324 9.3005
R1534 VTAIL.n327 VTAIL.n326 9.3005
R1535 VTAIL.n265 VTAIL.n263 9.3005
R1536 VTAIL.n333 VTAIL.n332 9.3005
R1537 VTAIL.n341 VTAIL.n340 9.3005
R1538 VTAIL.n260 VTAIL.n259 9.3005
R1539 VTAIL.n335 VTAIL.n334 9.3005
R1540 VTAIL.n311 VTAIL.n310 9.3005
R1541 VTAIL.n309 VTAIL.n308 9.3005
R1542 VTAIL.n278 VTAIL.n277 9.3005
R1543 VTAIL.n303 VTAIL.n302 9.3005
R1544 VTAIL.n301 VTAIL.n300 9.3005
R1545 VTAIL.n282 VTAIL.n281 9.3005
R1546 VTAIL.n295 VTAIL.n294 9.3005
R1547 VTAIL.n293 VTAIL.n292 9.3005
R1548 VTAIL.n286 VTAIL.n285 9.3005
R1549 VTAIL.n646 VTAIL.n645 8.92171
R1550 VTAIL.n661 VTAIL.n614 8.92171
R1551 VTAIL.n44 VTAIL.n43 8.92171
R1552 VTAIL.n59 VTAIL.n12 8.92171
R1553 VTAIL.n130 VTAIL.n129 8.92171
R1554 VTAIL.n145 VTAIL.n98 8.92171
R1555 VTAIL.n216 VTAIL.n215 8.92171
R1556 VTAIL.n231 VTAIL.n184 8.92171
R1557 VTAIL.n577 VTAIL.n530 8.92171
R1558 VTAIL.n562 VTAIL.n561 8.92171
R1559 VTAIL.n491 VTAIL.n444 8.92171
R1560 VTAIL.n476 VTAIL.n475 8.92171
R1561 VTAIL.n405 VTAIL.n358 8.92171
R1562 VTAIL.n390 VTAIL.n389 8.92171
R1563 VTAIL.n319 VTAIL.n272 8.92171
R1564 VTAIL.n304 VTAIL.n303 8.92171
R1565 VTAIL.n649 VTAIL.n620 8.14595
R1566 VTAIL.n658 VTAIL.n657 8.14595
R1567 VTAIL.n47 VTAIL.n18 8.14595
R1568 VTAIL.n56 VTAIL.n55 8.14595
R1569 VTAIL.n133 VTAIL.n104 8.14595
R1570 VTAIL.n142 VTAIL.n141 8.14595
R1571 VTAIL.n219 VTAIL.n190 8.14595
R1572 VTAIL.n228 VTAIL.n227 8.14595
R1573 VTAIL.n574 VTAIL.n573 8.14595
R1574 VTAIL.n565 VTAIL.n536 8.14595
R1575 VTAIL.n488 VTAIL.n487 8.14595
R1576 VTAIL.n479 VTAIL.n450 8.14595
R1577 VTAIL.n402 VTAIL.n401 8.14595
R1578 VTAIL.n393 VTAIL.n364 8.14595
R1579 VTAIL.n316 VTAIL.n315 8.14595
R1580 VTAIL.n307 VTAIL.n278 8.14595
R1581 VTAIL.n650 VTAIL.n618 7.3702
R1582 VTAIL.n654 VTAIL.n616 7.3702
R1583 VTAIL.n48 VTAIL.n16 7.3702
R1584 VTAIL.n52 VTAIL.n14 7.3702
R1585 VTAIL.n134 VTAIL.n102 7.3702
R1586 VTAIL.n138 VTAIL.n100 7.3702
R1587 VTAIL.n220 VTAIL.n188 7.3702
R1588 VTAIL.n224 VTAIL.n186 7.3702
R1589 VTAIL.n570 VTAIL.n532 7.3702
R1590 VTAIL.n566 VTAIL.n534 7.3702
R1591 VTAIL.n484 VTAIL.n446 7.3702
R1592 VTAIL.n480 VTAIL.n448 7.3702
R1593 VTAIL.n398 VTAIL.n360 7.3702
R1594 VTAIL.n394 VTAIL.n362 7.3702
R1595 VTAIL.n312 VTAIL.n274 7.3702
R1596 VTAIL.n308 VTAIL.n276 7.3702
R1597 VTAIL.n653 VTAIL.n618 6.59444
R1598 VTAIL.n654 VTAIL.n653 6.59444
R1599 VTAIL.n51 VTAIL.n16 6.59444
R1600 VTAIL.n52 VTAIL.n51 6.59444
R1601 VTAIL.n137 VTAIL.n102 6.59444
R1602 VTAIL.n138 VTAIL.n137 6.59444
R1603 VTAIL.n223 VTAIL.n188 6.59444
R1604 VTAIL.n224 VTAIL.n223 6.59444
R1605 VTAIL.n570 VTAIL.n569 6.59444
R1606 VTAIL.n569 VTAIL.n534 6.59444
R1607 VTAIL.n484 VTAIL.n483 6.59444
R1608 VTAIL.n483 VTAIL.n448 6.59444
R1609 VTAIL.n398 VTAIL.n397 6.59444
R1610 VTAIL.n397 VTAIL.n362 6.59444
R1611 VTAIL.n312 VTAIL.n311 6.59444
R1612 VTAIL.n311 VTAIL.n276 6.59444
R1613 VTAIL.n650 VTAIL.n649 5.81868
R1614 VTAIL.n657 VTAIL.n616 5.81868
R1615 VTAIL.n48 VTAIL.n47 5.81868
R1616 VTAIL.n55 VTAIL.n14 5.81868
R1617 VTAIL.n134 VTAIL.n133 5.81868
R1618 VTAIL.n141 VTAIL.n100 5.81868
R1619 VTAIL.n220 VTAIL.n219 5.81868
R1620 VTAIL.n227 VTAIL.n186 5.81868
R1621 VTAIL.n573 VTAIL.n532 5.81868
R1622 VTAIL.n566 VTAIL.n565 5.81868
R1623 VTAIL.n487 VTAIL.n446 5.81868
R1624 VTAIL.n480 VTAIL.n479 5.81868
R1625 VTAIL.n401 VTAIL.n360 5.81868
R1626 VTAIL.n394 VTAIL.n393 5.81868
R1627 VTAIL.n315 VTAIL.n274 5.81868
R1628 VTAIL.n308 VTAIL.n307 5.81868
R1629 VTAIL.n646 VTAIL.n620 5.04292
R1630 VTAIL.n658 VTAIL.n614 5.04292
R1631 VTAIL.n44 VTAIL.n18 5.04292
R1632 VTAIL.n56 VTAIL.n12 5.04292
R1633 VTAIL.n130 VTAIL.n104 5.04292
R1634 VTAIL.n142 VTAIL.n98 5.04292
R1635 VTAIL.n216 VTAIL.n190 5.04292
R1636 VTAIL.n228 VTAIL.n184 5.04292
R1637 VTAIL.n574 VTAIL.n530 5.04292
R1638 VTAIL.n562 VTAIL.n536 5.04292
R1639 VTAIL.n488 VTAIL.n444 5.04292
R1640 VTAIL.n476 VTAIL.n450 5.04292
R1641 VTAIL.n402 VTAIL.n358 5.04292
R1642 VTAIL.n390 VTAIL.n364 5.04292
R1643 VTAIL.n316 VTAIL.n272 5.04292
R1644 VTAIL.n304 VTAIL.n278 5.04292
R1645 VTAIL.n645 VTAIL.n622 4.26717
R1646 VTAIL.n662 VTAIL.n661 4.26717
R1647 VTAIL.n43 VTAIL.n20 4.26717
R1648 VTAIL.n60 VTAIL.n59 4.26717
R1649 VTAIL.n129 VTAIL.n106 4.26717
R1650 VTAIL.n146 VTAIL.n145 4.26717
R1651 VTAIL.n215 VTAIL.n192 4.26717
R1652 VTAIL.n232 VTAIL.n231 4.26717
R1653 VTAIL.n578 VTAIL.n577 4.26717
R1654 VTAIL.n561 VTAIL.n538 4.26717
R1655 VTAIL.n492 VTAIL.n491 4.26717
R1656 VTAIL.n475 VTAIL.n452 4.26717
R1657 VTAIL.n406 VTAIL.n405 4.26717
R1658 VTAIL.n389 VTAIL.n366 4.26717
R1659 VTAIL.n320 VTAIL.n319 4.26717
R1660 VTAIL.n303 VTAIL.n280 4.26717
R1661 VTAIL.n629 VTAIL.n627 3.70982
R1662 VTAIL.n27 VTAIL.n25 3.70982
R1663 VTAIL.n113 VTAIL.n111 3.70982
R1664 VTAIL.n199 VTAIL.n197 3.70982
R1665 VTAIL.n545 VTAIL.n543 3.70982
R1666 VTAIL.n459 VTAIL.n457 3.70982
R1667 VTAIL.n373 VTAIL.n371 3.70982
R1668 VTAIL.n287 VTAIL.n285 3.70982
R1669 VTAIL.n642 VTAIL.n641 3.49141
R1670 VTAIL.n665 VTAIL.n612 3.49141
R1671 VTAIL.n40 VTAIL.n39 3.49141
R1672 VTAIL.n63 VTAIL.n10 3.49141
R1673 VTAIL.n126 VTAIL.n125 3.49141
R1674 VTAIL.n149 VTAIL.n96 3.49141
R1675 VTAIL.n212 VTAIL.n211 3.49141
R1676 VTAIL.n235 VTAIL.n182 3.49141
R1677 VTAIL.n581 VTAIL.n528 3.49141
R1678 VTAIL.n558 VTAIL.n557 3.49141
R1679 VTAIL.n495 VTAIL.n442 3.49141
R1680 VTAIL.n472 VTAIL.n471 3.49141
R1681 VTAIL.n409 VTAIL.n356 3.49141
R1682 VTAIL.n386 VTAIL.n385 3.49141
R1683 VTAIL.n323 VTAIL.n270 3.49141
R1684 VTAIL.n300 VTAIL.n299 3.49141
R1685 VTAIL.n638 VTAIL.n624 2.71565
R1686 VTAIL.n666 VTAIL.n610 2.71565
R1687 VTAIL.n686 VTAIL.n602 2.71565
R1688 VTAIL.n36 VTAIL.n22 2.71565
R1689 VTAIL.n64 VTAIL.n8 2.71565
R1690 VTAIL.n84 VTAIL.n0 2.71565
R1691 VTAIL.n122 VTAIL.n108 2.71565
R1692 VTAIL.n150 VTAIL.n94 2.71565
R1693 VTAIL.n170 VTAIL.n86 2.71565
R1694 VTAIL.n208 VTAIL.n194 2.71565
R1695 VTAIL.n236 VTAIL.n180 2.71565
R1696 VTAIL.n256 VTAIL.n172 2.71565
R1697 VTAIL.n600 VTAIL.n516 2.71565
R1698 VTAIL.n582 VTAIL.n526 2.71565
R1699 VTAIL.n554 VTAIL.n540 2.71565
R1700 VTAIL.n514 VTAIL.n430 2.71565
R1701 VTAIL.n496 VTAIL.n440 2.71565
R1702 VTAIL.n468 VTAIL.n454 2.71565
R1703 VTAIL.n428 VTAIL.n344 2.71565
R1704 VTAIL.n410 VTAIL.n354 2.71565
R1705 VTAIL.n382 VTAIL.n368 2.71565
R1706 VTAIL.n342 VTAIL.n258 2.71565
R1707 VTAIL.n324 VTAIL.n268 2.71565
R1708 VTAIL.n296 VTAIL.n282 2.71565
R1709 VTAIL.n637 VTAIL.n626 1.93989
R1710 VTAIL.n671 VTAIL.n669 1.93989
R1711 VTAIL.n684 VTAIL.n683 1.93989
R1712 VTAIL.n35 VTAIL.n24 1.93989
R1713 VTAIL.n69 VTAIL.n67 1.93989
R1714 VTAIL.n82 VTAIL.n81 1.93989
R1715 VTAIL.n121 VTAIL.n110 1.93989
R1716 VTAIL.n155 VTAIL.n153 1.93989
R1717 VTAIL.n168 VTAIL.n167 1.93989
R1718 VTAIL.n207 VTAIL.n196 1.93989
R1719 VTAIL.n241 VTAIL.n239 1.93989
R1720 VTAIL.n254 VTAIL.n253 1.93989
R1721 VTAIL.n598 VTAIL.n597 1.93989
R1722 VTAIL.n586 VTAIL.n585 1.93989
R1723 VTAIL.n553 VTAIL.n542 1.93989
R1724 VTAIL.n512 VTAIL.n511 1.93989
R1725 VTAIL.n500 VTAIL.n499 1.93989
R1726 VTAIL.n467 VTAIL.n456 1.93989
R1727 VTAIL.n426 VTAIL.n425 1.93989
R1728 VTAIL.n414 VTAIL.n413 1.93989
R1729 VTAIL.n381 VTAIL.n370 1.93989
R1730 VTAIL.n340 VTAIL.n339 1.93989
R1731 VTAIL.n328 VTAIL.n327 1.93989
R1732 VTAIL.n295 VTAIL.n284 1.93989
R1733 VTAIL.n634 VTAIL.n633 1.16414
R1734 VTAIL.n670 VTAIL.n608 1.16414
R1735 VTAIL.n680 VTAIL.n604 1.16414
R1736 VTAIL.n32 VTAIL.n31 1.16414
R1737 VTAIL.n68 VTAIL.n6 1.16414
R1738 VTAIL.n78 VTAIL.n2 1.16414
R1739 VTAIL.n118 VTAIL.n117 1.16414
R1740 VTAIL.n154 VTAIL.n92 1.16414
R1741 VTAIL.n164 VTAIL.n88 1.16414
R1742 VTAIL.n204 VTAIL.n203 1.16414
R1743 VTAIL.n240 VTAIL.n178 1.16414
R1744 VTAIL.n250 VTAIL.n174 1.16414
R1745 VTAIL.n594 VTAIL.n518 1.16414
R1746 VTAIL.n589 VTAIL.n523 1.16414
R1747 VTAIL.n550 VTAIL.n549 1.16414
R1748 VTAIL.n508 VTAIL.n432 1.16414
R1749 VTAIL.n503 VTAIL.n437 1.16414
R1750 VTAIL.n464 VTAIL.n463 1.16414
R1751 VTAIL.n422 VTAIL.n346 1.16414
R1752 VTAIL.n417 VTAIL.n351 1.16414
R1753 VTAIL.n378 VTAIL.n377 1.16414
R1754 VTAIL.n336 VTAIL.n260 1.16414
R1755 VTAIL.n331 VTAIL.n265 1.16414
R1756 VTAIL.n292 VTAIL.n291 1.16414
R1757 VTAIL.n429 VTAIL.n343 0.647052
R1758 VTAIL.n601 VTAIL.n515 0.647052
R1759 VTAIL.n257 VTAIL.n171 0.647052
R1760 VTAIL.n515 VTAIL.n429 0.470328
R1761 VTAIL.n171 VTAIL.n85 0.470328
R1762 VTAIL.n630 VTAIL.n628 0.388379
R1763 VTAIL.n676 VTAIL.n675 0.388379
R1764 VTAIL.n679 VTAIL.n606 0.388379
R1765 VTAIL.n28 VTAIL.n26 0.388379
R1766 VTAIL.n74 VTAIL.n73 0.388379
R1767 VTAIL.n77 VTAIL.n4 0.388379
R1768 VTAIL.n114 VTAIL.n112 0.388379
R1769 VTAIL.n160 VTAIL.n159 0.388379
R1770 VTAIL.n163 VTAIL.n90 0.388379
R1771 VTAIL.n200 VTAIL.n198 0.388379
R1772 VTAIL.n246 VTAIL.n245 0.388379
R1773 VTAIL.n249 VTAIL.n176 0.388379
R1774 VTAIL.n593 VTAIL.n520 0.388379
R1775 VTAIL.n590 VTAIL.n522 0.388379
R1776 VTAIL.n546 VTAIL.n544 0.388379
R1777 VTAIL.n507 VTAIL.n434 0.388379
R1778 VTAIL.n504 VTAIL.n436 0.388379
R1779 VTAIL.n460 VTAIL.n458 0.388379
R1780 VTAIL.n421 VTAIL.n348 0.388379
R1781 VTAIL.n418 VTAIL.n350 0.388379
R1782 VTAIL.n374 VTAIL.n372 0.388379
R1783 VTAIL.n335 VTAIL.n262 0.388379
R1784 VTAIL.n332 VTAIL.n264 0.388379
R1785 VTAIL.n288 VTAIL.n286 0.388379
R1786 VTAIL VTAIL.n85 0.381966
R1787 VTAIL VTAIL.n687 0.265586
R1788 VTAIL.n635 VTAIL.n627 0.155672
R1789 VTAIL.n636 VTAIL.n635 0.155672
R1790 VTAIL.n636 VTAIL.n623 0.155672
R1791 VTAIL.n643 VTAIL.n623 0.155672
R1792 VTAIL.n644 VTAIL.n643 0.155672
R1793 VTAIL.n644 VTAIL.n619 0.155672
R1794 VTAIL.n651 VTAIL.n619 0.155672
R1795 VTAIL.n652 VTAIL.n651 0.155672
R1796 VTAIL.n652 VTAIL.n615 0.155672
R1797 VTAIL.n659 VTAIL.n615 0.155672
R1798 VTAIL.n660 VTAIL.n659 0.155672
R1799 VTAIL.n660 VTAIL.n611 0.155672
R1800 VTAIL.n667 VTAIL.n611 0.155672
R1801 VTAIL.n668 VTAIL.n667 0.155672
R1802 VTAIL.n668 VTAIL.n607 0.155672
R1803 VTAIL.n677 VTAIL.n607 0.155672
R1804 VTAIL.n678 VTAIL.n677 0.155672
R1805 VTAIL.n678 VTAIL.n603 0.155672
R1806 VTAIL.n685 VTAIL.n603 0.155672
R1807 VTAIL.n33 VTAIL.n25 0.155672
R1808 VTAIL.n34 VTAIL.n33 0.155672
R1809 VTAIL.n34 VTAIL.n21 0.155672
R1810 VTAIL.n41 VTAIL.n21 0.155672
R1811 VTAIL.n42 VTAIL.n41 0.155672
R1812 VTAIL.n42 VTAIL.n17 0.155672
R1813 VTAIL.n49 VTAIL.n17 0.155672
R1814 VTAIL.n50 VTAIL.n49 0.155672
R1815 VTAIL.n50 VTAIL.n13 0.155672
R1816 VTAIL.n57 VTAIL.n13 0.155672
R1817 VTAIL.n58 VTAIL.n57 0.155672
R1818 VTAIL.n58 VTAIL.n9 0.155672
R1819 VTAIL.n65 VTAIL.n9 0.155672
R1820 VTAIL.n66 VTAIL.n65 0.155672
R1821 VTAIL.n66 VTAIL.n5 0.155672
R1822 VTAIL.n75 VTAIL.n5 0.155672
R1823 VTAIL.n76 VTAIL.n75 0.155672
R1824 VTAIL.n76 VTAIL.n1 0.155672
R1825 VTAIL.n83 VTAIL.n1 0.155672
R1826 VTAIL.n119 VTAIL.n111 0.155672
R1827 VTAIL.n120 VTAIL.n119 0.155672
R1828 VTAIL.n120 VTAIL.n107 0.155672
R1829 VTAIL.n127 VTAIL.n107 0.155672
R1830 VTAIL.n128 VTAIL.n127 0.155672
R1831 VTAIL.n128 VTAIL.n103 0.155672
R1832 VTAIL.n135 VTAIL.n103 0.155672
R1833 VTAIL.n136 VTAIL.n135 0.155672
R1834 VTAIL.n136 VTAIL.n99 0.155672
R1835 VTAIL.n143 VTAIL.n99 0.155672
R1836 VTAIL.n144 VTAIL.n143 0.155672
R1837 VTAIL.n144 VTAIL.n95 0.155672
R1838 VTAIL.n151 VTAIL.n95 0.155672
R1839 VTAIL.n152 VTAIL.n151 0.155672
R1840 VTAIL.n152 VTAIL.n91 0.155672
R1841 VTAIL.n161 VTAIL.n91 0.155672
R1842 VTAIL.n162 VTAIL.n161 0.155672
R1843 VTAIL.n162 VTAIL.n87 0.155672
R1844 VTAIL.n169 VTAIL.n87 0.155672
R1845 VTAIL.n205 VTAIL.n197 0.155672
R1846 VTAIL.n206 VTAIL.n205 0.155672
R1847 VTAIL.n206 VTAIL.n193 0.155672
R1848 VTAIL.n213 VTAIL.n193 0.155672
R1849 VTAIL.n214 VTAIL.n213 0.155672
R1850 VTAIL.n214 VTAIL.n189 0.155672
R1851 VTAIL.n221 VTAIL.n189 0.155672
R1852 VTAIL.n222 VTAIL.n221 0.155672
R1853 VTAIL.n222 VTAIL.n185 0.155672
R1854 VTAIL.n229 VTAIL.n185 0.155672
R1855 VTAIL.n230 VTAIL.n229 0.155672
R1856 VTAIL.n230 VTAIL.n181 0.155672
R1857 VTAIL.n237 VTAIL.n181 0.155672
R1858 VTAIL.n238 VTAIL.n237 0.155672
R1859 VTAIL.n238 VTAIL.n177 0.155672
R1860 VTAIL.n247 VTAIL.n177 0.155672
R1861 VTAIL.n248 VTAIL.n247 0.155672
R1862 VTAIL.n248 VTAIL.n173 0.155672
R1863 VTAIL.n255 VTAIL.n173 0.155672
R1864 VTAIL.n599 VTAIL.n517 0.155672
R1865 VTAIL.n592 VTAIL.n517 0.155672
R1866 VTAIL.n592 VTAIL.n591 0.155672
R1867 VTAIL.n591 VTAIL.n521 0.155672
R1868 VTAIL.n584 VTAIL.n521 0.155672
R1869 VTAIL.n584 VTAIL.n583 0.155672
R1870 VTAIL.n583 VTAIL.n527 0.155672
R1871 VTAIL.n576 VTAIL.n527 0.155672
R1872 VTAIL.n576 VTAIL.n575 0.155672
R1873 VTAIL.n575 VTAIL.n531 0.155672
R1874 VTAIL.n568 VTAIL.n531 0.155672
R1875 VTAIL.n568 VTAIL.n567 0.155672
R1876 VTAIL.n567 VTAIL.n535 0.155672
R1877 VTAIL.n560 VTAIL.n535 0.155672
R1878 VTAIL.n560 VTAIL.n559 0.155672
R1879 VTAIL.n559 VTAIL.n539 0.155672
R1880 VTAIL.n552 VTAIL.n539 0.155672
R1881 VTAIL.n552 VTAIL.n551 0.155672
R1882 VTAIL.n551 VTAIL.n543 0.155672
R1883 VTAIL.n513 VTAIL.n431 0.155672
R1884 VTAIL.n506 VTAIL.n431 0.155672
R1885 VTAIL.n506 VTAIL.n505 0.155672
R1886 VTAIL.n505 VTAIL.n435 0.155672
R1887 VTAIL.n498 VTAIL.n435 0.155672
R1888 VTAIL.n498 VTAIL.n497 0.155672
R1889 VTAIL.n497 VTAIL.n441 0.155672
R1890 VTAIL.n490 VTAIL.n441 0.155672
R1891 VTAIL.n490 VTAIL.n489 0.155672
R1892 VTAIL.n489 VTAIL.n445 0.155672
R1893 VTAIL.n482 VTAIL.n445 0.155672
R1894 VTAIL.n482 VTAIL.n481 0.155672
R1895 VTAIL.n481 VTAIL.n449 0.155672
R1896 VTAIL.n474 VTAIL.n449 0.155672
R1897 VTAIL.n474 VTAIL.n473 0.155672
R1898 VTAIL.n473 VTAIL.n453 0.155672
R1899 VTAIL.n466 VTAIL.n453 0.155672
R1900 VTAIL.n466 VTAIL.n465 0.155672
R1901 VTAIL.n465 VTAIL.n457 0.155672
R1902 VTAIL.n427 VTAIL.n345 0.155672
R1903 VTAIL.n420 VTAIL.n345 0.155672
R1904 VTAIL.n420 VTAIL.n419 0.155672
R1905 VTAIL.n419 VTAIL.n349 0.155672
R1906 VTAIL.n412 VTAIL.n349 0.155672
R1907 VTAIL.n412 VTAIL.n411 0.155672
R1908 VTAIL.n411 VTAIL.n355 0.155672
R1909 VTAIL.n404 VTAIL.n355 0.155672
R1910 VTAIL.n404 VTAIL.n403 0.155672
R1911 VTAIL.n403 VTAIL.n359 0.155672
R1912 VTAIL.n396 VTAIL.n359 0.155672
R1913 VTAIL.n396 VTAIL.n395 0.155672
R1914 VTAIL.n395 VTAIL.n363 0.155672
R1915 VTAIL.n388 VTAIL.n363 0.155672
R1916 VTAIL.n388 VTAIL.n387 0.155672
R1917 VTAIL.n387 VTAIL.n367 0.155672
R1918 VTAIL.n380 VTAIL.n367 0.155672
R1919 VTAIL.n380 VTAIL.n379 0.155672
R1920 VTAIL.n379 VTAIL.n371 0.155672
R1921 VTAIL.n341 VTAIL.n259 0.155672
R1922 VTAIL.n334 VTAIL.n259 0.155672
R1923 VTAIL.n334 VTAIL.n333 0.155672
R1924 VTAIL.n333 VTAIL.n263 0.155672
R1925 VTAIL.n326 VTAIL.n263 0.155672
R1926 VTAIL.n326 VTAIL.n325 0.155672
R1927 VTAIL.n325 VTAIL.n269 0.155672
R1928 VTAIL.n318 VTAIL.n269 0.155672
R1929 VTAIL.n318 VTAIL.n317 0.155672
R1930 VTAIL.n317 VTAIL.n273 0.155672
R1931 VTAIL.n310 VTAIL.n273 0.155672
R1932 VTAIL.n310 VTAIL.n309 0.155672
R1933 VTAIL.n309 VTAIL.n277 0.155672
R1934 VTAIL.n302 VTAIL.n277 0.155672
R1935 VTAIL.n302 VTAIL.n301 0.155672
R1936 VTAIL.n301 VTAIL.n281 0.155672
R1937 VTAIL.n294 VTAIL.n281 0.155672
R1938 VTAIL.n294 VTAIL.n293 0.155672
R1939 VTAIL.n293 VTAIL.n285 0.155672
R1940 VP.n0 VP.t0 1008.51
R1941 VP.n0 VP.t2 1008.48
R1942 VP.n2 VP.t1 987.527
R1943 VP.n3 VP.t3 987.527
R1944 VP.n4 VP.n3 161.3
R1945 VP.n2 VP.n1 161.3
R1946 VP.n1 VP.n0 112.448
R1947 VP.n3 VP.n2 48.2005
R1948 VP.n4 VP.n1 0.189894
R1949 VP VP.n4 0.0516364
R1950 VDD1 VDD1.n1 113.73
R1951 VDD1 VDD1.n0 74.1949
R1952 VDD1.n0 VDD1.t3 2.08951
R1953 VDD1.n0 VDD1.t1 2.08951
R1954 VDD1.n1 VDD1.t2 2.08951
R1955 VDD1.n1 VDD1.t0 2.08951
C0 w_n1420_n4080# VDD2 1.10573f
C1 VP VTAIL 2.50054f
C2 VDD1 VTAIL 10.3134f
C3 B VTAIL 4.52058f
C4 VN VTAIL 2.48644f
C5 VP VDD2 0.25536f
C6 VP w_n1420_n4080# 2.25459f
C7 VDD1 VDD2 0.506056f
C8 VDD1 w_n1420_n4080# 1.09661f
C9 B VDD2 0.989594f
C10 B w_n1420_n4080# 7.56769f
C11 VN VDD2 3.11346f
C12 VN w_n1420_n4080# 2.07756f
C13 VDD1 VP 3.22183f
C14 B VP 1.01712f
C15 VP VN 5.2847f
C16 VDD1 B 0.971971f
C17 VDD1 VN 0.146801f
C18 B VN 0.733489f
C19 VTAIL VDD2 10.353f
C20 VTAIL w_n1420_n4080# 5.1569f
C21 VDD2 VSUBS 0.730785f
C22 VDD1 VSUBS 5.763757f
C23 VTAIL VSUBS 0.918489f
C24 VN VSUBS 6.67555f
C25 VP VSUBS 1.28088f
C26 B VSUBS 2.680968f
C27 w_n1420_n4080# VSUBS 71.0057f
C28 VDD1.t3 VSUBS 0.37857f
C29 VDD1.t1 VSUBS 0.37857f
C30 VDD1.n0 VSUBS 3.10556f
C31 VDD1.t2 VSUBS 0.37857f
C32 VDD1.t0 VSUBS 0.37857f
C33 VDD1.n1 VSUBS 3.94406f
C34 VP.t2 VSUBS 1.31272f
C35 VP.t0 VSUBS 1.31274f
C36 VP.n0 VSUBS 2.1214f
C37 VP.n1 VSUBS 4.85574f
C38 VP.t1 VSUBS 1.30217f
C39 VP.n2 VSUBS 0.507777f
C40 VP.t3 VSUBS 1.30217f
C41 VP.n3 VSUBS 0.507777f
C42 VP.n4 VSUBS 0.054366f
C43 VTAIL.n0 VSUBS 0.026731f
C44 VTAIL.n1 VSUBS 0.024048f
C45 VTAIL.n2 VSUBS 0.012923f
C46 VTAIL.n3 VSUBS 0.030544f
C47 VTAIL.n4 VSUBS 0.013303f
C48 VTAIL.n5 VSUBS 0.024048f
C49 VTAIL.n6 VSUBS 0.013683f
C50 VTAIL.n7 VSUBS 0.030544f
C51 VTAIL.n8 VSUBS 0.013683f
C52 VTAIL.n9 VSUBS 0.024048f
C53 VTAIL.n10 VSUBS 0.012923f
C54 VTAIL.n11 VSUBS 0.030544f
C55 VTAIL.n12 VSUBS 0.013683f
C56 VTAIL.n13 VSUBS 0.024048f
C57 VTAIL.n14 VSUBS 0.012923f
C58 VTAIL.n15 VSUBS 0.030544f
C59 VTAIL.n16 VSUBS 0.013683f
C60 VTAIL.n17 VSUBS 0.024048f
C61 VTAIL.n18 VSUBS 0.012923f
C62 VTAIL.n19 VSUBS 0.030544f
C63 VTAIL.n20 VSUBS 0.013683f
C64 VTAIL.n21 VSUBS 0.024048f
C65 VTAIL.n22 VSUBS 0.012923f
C66 VTAIL.n23 VSUBS 0.030544f
C67 VTAIL.n24 VSUBS 0.013683f
C68 VTAIL.n25 VSUBS 1.59668f
C69 VTAIL.n26 VSUBS 0.012923f
C70 VTAIL.t7 VSUBS 0.065423f
C71 VTAIL.n27 VSUBS 0.173494f
C72 VTAIL.n28 VSUBS 0.019431f
C73 VTAIL.n29 VSUBS 0.022908f
C74 VTAIL.n30 VSUBS 0.030544f
C75 VTAIL.n31 VSUBS 0.013683f
C76 VTAIL.n32 VSUBS 0.012923f
C77 VTAIL.n33 VSUBS 0.024048f
C78 VTAIL.n34 VSUBS 0.024048f
C79 VTAIL.n35 VSUBS 0.012923f
C80 VTAIL.n36 VSUBS 0.013683f
C81 VTAIL.n37 VSUBS 0.030544f
C82 VTAIL.n38 VSUBS 0.030544f
C83 VTAIL.n39 VSUBS 0.013683f
C84 VTAIL.n40 VSUBS 0.012923f
C85 VTAIL.n41 VSUBS 0.024048f
C86 VTAIL.n42 VSUBS 0.024048f
C87 VTAIL.n43 VSUBS 0.012923f
C88 VTAIL.n44 VSUBS 0.013683f
C89 VTAIL.n45 VSUBS 0.030544f
C90 VTAIL.n46 VSUBS 0.030544f
C91 VTAIL.n47 VSUBS 0.013683f
C92 VTAIL.n48 VSUBS 0.012923f
C93 VTAIL.n49 VSUBS 0.024048f
C94 VTAIL.n50 VSUBS 0.024048f
C95 VTAIL.n51 VSUBS 0.012923f
C96 VTAIL.n52 VSUBS 0.013683f
C97 VTAIL.n53 VSUBS 0.030544f
C98 VTAIL.n54 VSUBS 0.030544f
C99 VTAIL.n55 VSUBS 0.013683f
C100 VTAIL.n56 VSUBS 0.012923f
C101 VTAIL.n57 VSUBS 0.024048f
C102 VTAIL.n58 VSUBS 0.024048f
C103 VTAIL.n59 VSUBS 0.012923f
C104 VTAIL.n60 VSUBS 0.013683f
C105 VTAIL.n61 VSUBS 0.030544f
C106 VTAIL.n62 VSUBS 0.030544f
C107 VTAIL.n63 VSUBS 0.013683f
C108 VTAIL.n64 VSUBS 0.012923f
C109 VTAIL.n65 VSUBS 0.024048f
C110 VTAIL.n66 VSUBS 0.024048f
C111 VTAIL.n67 VSUBS 0.012923f
C112 VTAIL.n68 VSUBS 0.012923f
C113 VTAIL.n69 VSUBS 0.013683f
C114 VTAIL.n70 VSUBS 0.030544f
C115 VTAIL.n71 VSUBS 0.030544f
C116 VTAIL.n72 VSUBS 0.030544f
C117 VTAIL.n73 VSUBS 0.013303f
C118 VTAIL.n74 VSUBS 0.012923f
C119 VTAIL.n75 VSUBS 0.024048f
C120 VTAIL.n76 VSUBS 0.024048f
C121 VTAIL.n77 VSUBS 0.012923f
C122 VTAIL.n78 VSUBS 0.013683f
C123 VTAIL.n79 VSUBS 0.030544f
C124 VTAIL.n80 VSUBS 0.074991f
C125 VTAIL.n81 VSUBS 0.013683f
C126 VTAIL.n82 VSUBS 0.012923f
C127 VTAIL.n83 VSUBS 0.062158f
C128 VTAIL.n84 VSUBS 0.037951f
C129 VTAIL.n85 VSUBS 0.090224f
C130 VTAIL.n86 VSUBS 0.026731f
C131 VTAIL.n87 VSUBS 0.024048f
C132 VTAIL.n88 VSUBS 0.012923f
C133 VTAIL.n89 VSUBS 0.030544f
C134 VTAIL.n90 VSUBS 0.013303f
C135 VTAIL.n91 VSUBS 0.024048f
C136 VTAIL.n92 VSUBS 0.013683f
C137 VTAIL.n93 VSUBS 0.030544f
C138 VTAIL.n94 VSUBS 0.013683f
C139 VTAIL.n95 VSUBS 0.024048f
C140 VTAIL.n96 VSUBS 0.012923f
C141 VTAIL.n97 VSUBS 0.030544f
C142 VTAIL.n98 VSUBS 0.013683f
C143 VTAIL.n99 VSUBS 0.024048f
C144 VTAIL.n100 VSUBS 0.012923f
C145 VTAIL.n101 VSUBS 0.030544f
C146 VTAIL.n102 VSUBS 0.013683f
C147 VTAIL.n103 VSUBS 0.024048f
C148 VTAIL.n104 VSUBS 0.012923f
C149 VTAIL.n105 VSUBS 0.030544f
C150 VTAIL.n106 VSUBS 0.013683f
C151 VTAIL.n107 VSUBS 0.024048f
C152 VTAIL.n108 VSUBS 0.012923f
C153 VTAIL.n109 VSUBS 0.030544f
C154 VTAIL.n110 VSUBS 0.013683f
C155 VTAIL.n111 VSUBS 1.59668f
C156 VTAIL.n112 VSUBS 0.012923f
C157 VTAIL.t3 VSUBS 0.065423f
C158 VTAIL.n113 VSUBS 0.173494f
C159 VTAIL.n114 VSUBS 0.019431f
C160 VTAIL.n115 VSUBS 0.022908f
C161 VTAIL.n116 VSUBS 0.030544f
C162 VTAIL.n117 VSUBS 0.013683f
C163 VTAIL.n118 VSUBS 0.012923f
C164 VTAIL.n119 VSUBS 0.024048f
C165 VTAIL.n120 VSUBS 0.024048f
C166 VTAIL.n121 VSUBS 0.012923f
C167 VTAIL.n122 VSUBS 0.013683f
C168 VTAIL.n123 VSUBS 0.030544f
C169 VTAIL.n124 VSUBS 0.030544f
C170 VTAIL.n125 VSUBS 0.013683f
C171 VTAIL.n126 VSUBS 0.012923f
C172 VTAIL.n127 VSUBS 0.024048f
C173 VTAIL.n128 VSUBS 0.024048f
C174 VTAIL.n129 VSUBS 0.012923f
C175 VTAIL.n130 VSUBS 0.013683f
C176 VTAIL.n131 VSUBS 0.030544f
C177 VTAIL.n132 VSUBS 0.030544f
C178 VTAIL.n133 VSUBS 0.013683f
C179 VTAIL.n134 VSUBS 0.012923f
C180 VTAIL.n135 VSUBS 0.024048f
C181 VTAIL.n136 VSUBS 0.024048f
C182 VTAIL.n137 VSUBS 0.012923f
C183 VTAIL.n138 VSUBS 0.013683f
C184 VTAIL.n139 VSUBS 0.030544f
C185 VTAIL.n140 VSUBS 0.030544f
C186 VTAIL.n141 VSUBS 0.013683f
C187 VTAIL.n142 VSUBS 0.012923f
C188 VTAIL.n143 VSUBS 0.024048f
C189 VTAIL.n144 VSUBS 0.024048f
C190 VTAIL.n145 VSUBS 0.012923f
C191 VTAIL.n146 VSUBS 0.013683f
C192 VTAIL.n147 VSUBS 0.030544f
C193 VTAIL.n148 VSUBS 0.030544f
C194 VTAIL.n149 VSUBS 0.013683f
C195 VTAIL.n150 VSUBS 0.012923f
C196 VTAIL.n151 VSUBS 0.024048f
C197 VTAIL.n152 VSUBS 0.024048f
C198 VTAIL.n153 VSUBS 0.012923f
C199 VTAIL.n154 VSUBS 0.012923f
C200 VTAIL.n155 VSUBS 0.013683f
C201 VTAIL.n156 VSUBS 0.030544f
C202 VTAIL.n157 VSUBS 0.030544f
C203 VTAIL.n158 VSUBS 0.030544f
C204 VTAIL.n159 VSUBS 0.013303f
C205 VTAIL.n160 VSUBS 0.012923f
C206 VTAIL.n161 VSUBS 0.024048f
C207 VTAIL.n162 VSUBS 0.024048f
C208 VTAIL.n163 VSUBS 0.012923f
C209 VTAIL.n164 VSUBS 0.013683f
C210 VTAIL.n165 VSUBS 0.030544f
C211 VTAIL.n166 VSUBS 0.074991f
C212 VTAIL.n167 VSUBS 0.013683f
C213 VTAIL.n168 VSUBS 0.012923f
C214 VTAIL.n169 VSUBS 0.062158f
C215 VTAIL.n170 VSUBS 0.037951f
C216 VTAIL.n171 VSUBS 0.110765f
C217 VTAIL.n172 VSUBS 0.026731f
C218 VTAIL.n173 VSUBS 0.024048f
C219 VTAIL.n174 VSUBS 0.012923f
C220 VTAIL.n175 VSUBS 0.030544f
C221 VTAIL.n176 VSUBS 0.013303f
C222 VTAIL.n177 VSUBS 0.024048f
C223 VTAIL.n178 VSUBS 0.013683f
C224 VTAIL.n179 VSUBS 0.030544f
C225 VTAIL.n180 VSUBS 0.013683f
C226 VTAIL.n181 VSUBS 0.024048f
C227 VTAIL.n182 VSUBS 0.012923f
C228 VTAIL.n183 VSUBS 0.030544f
C229 VTAIL.n184 VSUBS 0.013683f
C230 VTAIL.n185 VSUBS 0.024048f
C231 VTAIL.n186 VSUBS 0.012923f
C232 VTAIL.n187 VSUBS 0.030544f
C233 VTAIL.n188 VSUBS 0.013683f
C234 VTAIL.n189 VSUBS 0.024048f
C235 VTAIL.n190 VSUBS 0.012923f
C236 VTAIL.n191 VSUBS 0.030544f
C237 VTAIL.n192 VSUBS 0.013683f
C238 VTAIL.n193 VSUBS 0.024048f
C239 VTAIL.n194 VSUBS 0.012923f
C240 VTAIL.n195 VSUBS 0.030544f
C241 VTAIL.n196 VSUBS 0.013683f
C242 VTAIL.n197 VSUBS 1.59668f
C243 VTAIL.n198 VSUBS 0.012923f
C244 VTAIL.t2 VSUBS 0.065423f
C245 VTAIL.n199 VSUBS 0.173494f
C246 VTAIL.n200 VSUBS 0.019431f
C247 VTAIL.n201 VSUBS 0.022908f
C248 VTAIL.n202 VSUBS 0.030544f
C249 VTAIL.n203 VSUBS 0.013683f
C250 VTAIL.n204 VSUBS 0.012923f
C251 VTAIL.n205 VSUBS 0.024048f
C252 VTAIL.n206 VSUBS 0.024048f
C253 VTAIL.n207 VSUBS 0.012923f
C254 VTAIL.n208 VSUBS 0.013683f
C255 VTAIL.n209 VSUBS 0.030544f
C256 VTAIL.n210 VSUBS 0.030544f
C257 VTAIL.n211 VSUBS 0.013683f
C258 VTAIL.n212 VSUBS 0.012923f
C259 VTAIL.n213 VSUBS 0.024048f
C260 VTAIL.n214 VSUBS 0.024048f
C261 VTAIL.n215 VSUBS 0.012923f
C262 VTAIL.n216 VSUBS 0.013683f
C263 VTAIL.n217 VSUBS 0.030544f
C264 VTAIL.n218 VSUBS 0.030544f
C265 VTAIL.n219 VSUBS 0.013683f
C266 VTAIL.n220 VSUBS 0.012923f
C267 VTAIL.n221 VSUBS 0.024048f
C268 VTAIL.n222 VSUBS 0.024048f
C269 VTAIL.n223 VSUBS 0.012923f
C270 VTAIL.n224 VSUBS 0.013683f
C271 VTAIL.n225 VSUBS 0.030544f
C272 VTAIL.n226 VSUBS 0.030544f
C273 VTAIL.n227 VSUBS 0.013683f
C274 VTAIL.n228 VSUBS 0.012923f
C275 VTAIL.n229 VSUBS 0.024048f
C276 VTAIL.n230 VSUBS 0.024048f
C277 VTAIL.n231 VSUBS 0.012923f
C278 VTAIL.n232 VSUBS 0.013683f
C279 VTAIL.n233 VSUBS 0.030544f
C280 VTAIL.n234 VSUBS 0.030544f
C281 VTAIL.n235 VSUBS 0.013683f
C282 VTAIL.n236 VSUBS 0.012923f
C283 VTAIL.n237 VSUBS 0.024048f
C284 VTAIL.n238 VSUBS 0.024048f
C285 VTAIL.n239 VSUBS 0.012923f
C286 VTAIL.n240 VSUBS 0.012923f
C287 VTAIL.n241 VSUBS 0.013683f
C288 VTAIL.n242 VSUBS 0.030544f
C289 VTAIL.n243 VSUBS 0.030544f
C290 VTAIL.n244 VSUBS 0.030544f
C291 VTAIL.n245 VSUBS 0.013303f
C292 VTAIL.n246 VSUBS 0.012923f
C293 VTAIL.n247 VSUBS 0.024048f
C294 VTAIL.n248 VSUBS 0.024048f
C295 VTAIL.n249 VSUBS 0.012923f
C296 VTAIL.n250 VSUBS 0.013683f
C297 VTAIL.n251 VSUBS 0.030544f
C298 VTAIL.n252 VSUBS 0.074991f
C299 VTAIL.n253 VSUBS 0.013683f
C300 VTAIL.n254 VSUBS 0.012923f
C301 VTAIL.n255 VSUBS 0.062158f
C302 VTAIL.n256 VSUBS 0.037951f
C303 VTAIL.n257 VSUBS 1.49056f
C304 VTAIL.n258 VSUBS 0.026731f
C305 VTAIL.n259 VSUBS 0.024048f
C306 VTAIL.n260 VSUBS 0.012923f
C307 VTAIL.n261 VSUBS 0.030544f
C308 VTAIL.n262 VSUBS 0.013303f
C309 VTAIL.n263 VSUBS 0.024048f
C310 VTAIL.n264 VSUBS 0.013303f
C311 VTAIL.n265 VSUBS 0.012923f
C312 VTAIL.n266 VSUBS 0.030544f
C313 VTAIL.n267 VSUBS 0.030544f
C314 VTAIL.n268 VSUBS 0.013683f
C315 VTAIL.n269 VSUBS 0.024048f
C316 VTAIL.n270 VSUBS 0.012923f
C317 VTAIL.n271 VSUBS 0.030544f
C318 VTAIL.n272 VSUBS 0.013683f
C319 VTAIL.n273 VSUBS 0.024048f
C320 VTAIL.n274 VSUBS 0.012923f
C321 VTAIL.n275 VSUBS 0.030544f
C322 VTAIL.n276 VSUBS 0.013683f
C323 VTAIL.n277 VSUBS 0.024048f
C324 VTAIL.n278 VSUBS 0.012923f
C325 VTAIL.n279 VSUBS 0.030544f
C326 VTAIL.n280 VSUBS 0.013683f
C327 VTAIL.n281 VSUBS 0.024048f
C328 VTAIL.n282 VSUBS 0.012923f
C329 VTAIL.n283 VSUBS 0.030544f
C330 VTAIL.n284 VSUBS 0.013683f
C331 VTAIL.n285 VSUBS 1.59668f
C332 VTAIL.n286 VSUBS 0.012923f
C333 VTAIL.t5 VSUBS 0.065423f
C334 VTAIL.n287 VSUBS 0.173494f
C335 VTAIL.n288 VSUBS 0.019431f
C336 VTAIL.n289 VSUBS 0.022908f
C337 VTAIL.n290 VSUBS 0.030544f
C338 VTAIL.n291 VSUBS 0.013683f
C339 VTAIL.n292 VSUBS 0.012923f
C340 VTAIL.n293 VSUBS 0.024048f
C341 VTAIL.n294 VSUBS 0.024048f
C342 VTAIL.n295 VSUBS 0.012923f
C343 VTAIL.n296 VSUBS 0.013683f
C344 VTAIL.n297 VSUBS 0.030544f
C345 VTAIL.n298 VSUBS 0.030544f
C346 VTAIL.n299 VSUBS 0.013683f
C347 VTAIL.n300 VSUBS 0.012923f
C348 VTAIL.n301 VSUBS 0.024048f
C349 VTAIL.n302 VSUBS 0.024048f
C350 VTAIL.n303 VSUBS 0.012923f
C351 VTAIL.n304 VSUBS 0.013683f
C352 VTAIL.n305 VSUBS 0.030544f
C353 VTAIL.n306 VSUBS 0.030544f
C354 VTAIL.n307 VSUBS 0.013683f
C355 VTAIL.n308 VSUBS 0.012923f
C356 VTAIL.n309 VSUBS 0.024048f
C357 VTAIL.n310 VSUBS 0.024048f
C358 VTAIL.n311 VSUBS 0.012923f
C359 VTAIL.n312 VSUBS 0.013683f
C360 VTAIL.n313 VSUBS 0.030544f
C361 VTAIL.n314 VSUBS 0.030544f
C362 VTAIL.n315 VSUBS 0.013683f
C363 VTAIL.n316 VSUBS 0.012923f
C364 VTAIL.n317 VSUBS 0.024048f
C365 VTAIL.n318 VSUBS 0.024048f
C366 VTAIL.n319 VSUBS 0.012923f
C367 VTAIL.n320 VSUBS 0.013683f
C368 VTAIL.n321 VSUBS 0.030544f
C369 VTAIL.n322 VSUBS 0.030544f
C370 VTAIL.n323 VSUBS 0.013683f
C371 VTAIL.n324 VSUBS 0.012923f
C372 VTAIL.n325 VSUBS 0.024048f
C373 VTAIL.n326 VSUBS 0.024048f
C374 VTAIL.n327 VSUBS 0.012923f
C375 VTAIL.n328 VSUBS 0.013683f
C376 VTAIL.n329 VSUBS 0.030544f
C377 VTAIL.n330 VSUBS 0.030544f
C378 VTAIL.n331 VSUBS 0.013683f
C379 VTAIL.n332 VSUBS 0.012923f
C380 VTAIL.n333 VSUBS 0.024048f
C381 VTAIL.n334 VSUBS 0.024048f
C382 VTAIL.n335 VSUBS 0.012923f
C383 VTAIL.n336 VSUBS 0.013683f
C384 VTAIL.n337 VSUBS 0.030544f
C385 VTAIL.n338 VSUBS 0.074991f
C386 VTAIL.n339 VSUBS 0.013683f
C387 VTAIL.n340 VSUBS 0.012923f
C388 VTAIL.n341 VSUBS 0.062158f
C389 VTAIL.n342 VSUBS 0.037951f
C390 VTAIL.n343 VSUBS 1.49056f
C391 VTAIL.n344 VSUBS 0.026731f
C392 VTAIL.n345 VSUBS 0.024048f
C393 VTAIL.n346 VSUBS 0.012923f
C394 VTAIL.n347 VSUBS 0.030544f
C395 VTAIL.n348 VSUBS 0.013303f
C396 VTAIL.n349 VSUBS 0.024048f
C397 VTAIL.n350 VSUBS 0.013303f
C398 VTAIL.n351 VSUBS 0.012923f
C399 VTAIL.n352 VSUBS 0.030544f
C400 VTAIL.n353 VSUBS 0.030544f
C401 VTAIL.n354 VSUBS 0.013683f
C402 VTAIL.n355 VSUBS 0.024048f
C403 VTAIL.n356 VSUBS 0.012923f
C404 VTAIL.n357 VSUBS 0.030544f
C405 VTAIL.n358 VSUBS 0.013683f
C406 VTAIL.n359 VSUBS 0.024048f
C407 VTAIL.n360 VSUBS 0.012923f
C408 VTAIL.n361 VSUBS 0.030544f
C409 VTAIL.n362 VSUBS 0.013683f
C410 VTAIL.n363 VSUBS 0.024048f
C411 VTAIL.n364 VSUBS 0.012923f
C412 VTAIL.n365 VSUBS 0.030544f
C413 VTAIL.n366 VSUBS 0.013683f
C414 VTAIL.n367 VSUBS 0.024048f
C415 VTAIL.n368 VSUBS 0.012923f
C416 VTAIL.n369 VSUBS 0.030544f
C417 VTAIL.n370 VSUBS 0.013683f
C418 VTAIL.n371 VSUBS 1.59668f
C419 VTAIL.n372 VSUBS 0.012923f
C420 VTAIL.t6 VSUBS 0.065423f
C421 VTAIL.n373 VSUBS 0.173494f
C422 VTAIL.n374 VSUBS 0.019431f
C423 VTAIL.n375 VSUBS 0.022908f
C424 VTAIL.n376 VSUBS 0.030544f
C425 VTAIL.n377 VSUBS 0.013683f
C426 VTAIL.n378 VSUBS 0.012923f
C427 VTAIL.n379 VSUBS 0.024048f
C428 VTAIL.n380 VSUBS 0.024048f
C429 VTAIL.n381 VSUBS 0.012923f
C430 VTAIL.n382 VSUBS 0.013683f
C431 VTAIL.n383 VSUBS 0.030544f
C432 VTAIL.n384 VSUBS 0.030544f
C433 VTAIL.n385 VSUBS 0.013683f
C434 VTAIL.n386 VSUBS 0.012923f
C435 VTAIL.n387 VSUBS 0.024048f
C436 VTAIL.n388 VSUBS 0.024048f
C437 VTAIL.n389 VSUBS 0.012923f
C438 VTAIL.n390 VSUBS 0.013683f
C439 VTAIL.n391 VSUBS 0.030544f
C440 VTAIL.n392 VSUBS 0.030544f
C441 VTAIL.n393 VSUBS 0.013683f
C442 VTAIL.n394 VSUBS 0.012923f
C443 VTAIL.n395 VSUBS 0.024048f
C444 VTAIL.n396 VSUBS 0.024048f
C445 VTAIL.n397 VSUBS 0.012923f
C446 VTAIL.n398 VSUBS 0.013683f
C447 VTAIL.n399 VSUBS 0.030544f
C448 VTAIL.n400 VSUBS 0.030544f
C449 VTAIL.n401 VSUBS 0.013683f
C450 VTAIL.n402 VSUBS 0.012923f
C451 VTAIL.n403 VSUBS 0.024048f
C452 VTAIL.n404 VSUBS 0.024048f
C453 VTAIL.n405 VSUBS 0.012923f
C454 VTAIL.n406 VSUBS 0.013683f
C455 VTAIL.n407 VSUBS 0.030544f
C456 VTAIL.n408 VSUBS 0.030544f
C457 VTAIL.n409 VSUBS 0.013683f
C458 VTAIL.n410 VSUBS 0.012923f
C459 VTAIL.n411 VSUBS 0.024048f
C460 VTAIL.n412 VSUBS 0.024048f
C461 VTAIL.n413 VSUBS 0.012923f
C462 VTAIL.n414 VSUBS 0.013683f
C463 VTAIL.n415 VSUBS 0.030544f
C464 VTAIL.n416 VSUBS 0.030544f
C465 VTAIL.n417 VSUBS 0.013683f
C466 VTAIL.n418 VSUBS 0.012923f
C467 VTAIL.n419 VSUBS 0.024048f
C468 VTAIL.n420 VSUBS 0.024048f
C469 VTAIL.n421 VSUBS 0.012923f
C470 VTAIL.n422 VSUBS 0.013683f
C471 VTAIL.n423 VSUBS 0.030544f
C472 VTAIL.n424 VSUBS 0.074991f
C473 VTAIL.n425 VSUBS 0.013683f
C474 VTAIL.n426 VSUBS 0.012923f
C475 VTAIL.n427 VSUBS 0.062158f
C476 VTAIL.n428 VSUBS 0.037951f
C477 VTAIL.n429 VSUBS 0.110765f
C478 VTAIL.n430 VSUBS 0.026731f
C479 VTAIL.n431 VSUBS 0.024048f
C480 VTAIL.n432 VSUBS 0.012923f
C481 VTAIL.n433 VSUBS 0.030544f
C482 VTAIL.n434 VSUBS 0.013303f
C483 VTAIL.n435 VSUBS 0.024048f
C484 VTAIL.n436 VSUBS 0.013303f
C485 VTAIL.n437 VSUBS 0.012923f
C486 VTAIL.n438 VSUBS 0.030544f
C487 VTAIL.n439 VSUBS 0.030544f
C488 VTAIL.n440 VSUBS 0.013683f
C489 VTAIL.n441 VSUBS 0.024048f
C490 VTAIL.n442 VSUBS 0.012923f
C491 VTAIL.n443 VSUBS 0.030544f
C492 VTAIL.n444 VSUBS 0.013683f
C493 VTAIL.n445 VSUBS 0.024048f
C494 VTAIL.n446 VSUBS 0.012923f
C495 VTAIL.n447 VSUBS 0.030544f
C496 VTAIL.n448 VSUBS 0.013683f
C497 VTAIL.n449 VSUBS 0.024048f
C498 VTAIL.n450 VSUBS 0.012923f
C499 VTAIL.n451 VSUBS 0.030544f
C500 VTAIL.n452 VSUBS 0.013683f
C501 VTAIL.n453 VSUBS 0.024048f
C502 VTAIL.n454 VSUBS 0.012923f
C503 VTAIL.n455 VSUBS 0.030544f
C504 VTAIL.n456 VSUBS 0.013683f
C505 VTAIL.n457 VSUBS 1.59668f
C506 VTAIL.n458 VSUBS 0.012923f
C507 VTAIL.t1 VSUBS 0.065423f
C508 VTAIL.n459 VSUBS 0.173494f
C509 VTAIL.n460 VSUBS 0.019431f
C510 VTAIL.n461 VSUBS 0.022908f
C511 VTAIL.n462 VSUBS 0.030544f
C512 VTAIL.n463 VSUBS 0.013683f
C513 VTAIL.n464 VSUBS 0.012923f
C514 VTAIL.n465 VSUBS 0.024048f
C515 VTAIL.n466 VSUBS 0.024048f
C516 VTAIL.n467 VSUBS 0.012923f
C517 VTAIL.n468 VSUBS 0.013683f
C518 VTAIL.n469 VSUBS 0.030544f
C519 VTAIL.n470 VSUBS 0.030544f
C520 VTAIL.n471 VSUBS 0.013683f
C521 VTAIL.n472 VSUBS 0.012923f
C522 VTAIL.n473 VSUBS 0.024048f
C523 VTAIL.n474 VSUBS 0.024048f
C524 VTAIL.n475 VSUBS 0.012923f
C525 VTAIL.n476 VSUBS 0.013683f
C526 VTAIL.n477 VSUBS 0.030544f
C527 VTAIL.n478 VSUBS 0.030544f
C528 VTAIL.n479 VSUBS 0.013683f
C529 VTAIL.n480 VSUBS 0.012923f
C530 VTAIL.n481 VSUBS 0.024048f
C531 VTAIL.n482 VSUBS 0.024048f
C532 VTAIL.n483 VSUBS 0.012923f
C533 VTAIL.n484 VSUBS 0.013683f
C534 VTAIL.n485 VSUBS 0.030544f
C535 VTAIL.n486 VSUBS 0.030544f
C536 VTAIL.n487 VSUBS 0.013683f
C537 VTAIL.n488 VSUBS 0.012923f
C538 VTAIL.n489 VSUBS 0.024048f
C539 VTAIL.n490 VSUBS 0.024048f
C540 VTAIL.n491 VSUBS 0.012923f
C541 VTAIL.n492 VSUBS 0.013683f
C542 VTAIL.n493 VSUBS 0.030544f
C543 VTAIL.n494 VSUBS 0.030544f
C544 VTAIL.n495 VSUBS 0.013683f
C545 VTAIL.n496 VSUBS 0.012923f
C546 VTAIL.n497 VSUBS 0.024048f
C547 VTAIL.n498 VSUBS 0.024048f
C548 VTAIL.n499 VSUBS 0.012923f
C549 VTAIL.n500 VSUBS 0.013683f
C550 VTAIL.n501 VSUBS 0.030544f
C551 VTAIL.n502 VSUBS 0.030544f
C552 VTAIL.n503 VSUBS 0.013683f
C553 VTAIL.n504 VSUBS 0.012923f
C554 VTAIL.n505 VSUBS 0.024048f
C555 VTAIL.n506 VSUBS 0.024048f
C556 VTAIL.n507 VSUBS 0.012923f
C557 VTAIL.n508 VSUBS 0.013683f
C558 VTAIL.n509 VSUBS 0.030544f
C559 VTAIL.n510 VSUBS 0.074991f
C560 VTAIL.n511 VSUBS 0.013683f
C561 VTAIL.n512 VSUBS 0.012923f
C562 VTAIL.n513 VSUBS 0.062158f
C563 VTAIL.n514 VSUBS 0.037951f
C564 VTAIL.n515 VSUBS 0.110765f
C565 VTAIL.n516 VSUBS 0.026731f
C566 VTAIL.n517 VSUBS 0.024048f
C567 VTAIL.n518 VSUBS 0.012923f
C568 VTAIL.n519 VSUBS 0.030544f
C569 VTAIL.n520 VSUBS 0.013303f
C570 VTAIL.n521 VSUBS 0.024048f
C571 VTAIL.n522 VSUBS 0.013303f
C572 VTAIL.n523 VSUBS 0.012923f
C573 VTAIL.n524 VSUBS 0.030544f
C574 VTAIL.n525 VSUBS 0.030544f
C575 VTAIL.n526 VSUBS 0.013683f
C576 VTAIL.n527 VSUBS 0.024048f
C577 VTAIL.n528 VSUBS 0.012923f
C578 VTAIL.n529 VSUBS 0.030544f
C579 VTAIL.n530 VSUBS 0.013683f
C580 VTAIL.n531 VSUBS 0.024048f
C581 VTAIL.n532 VSUBS 0.012923f
C582 VTAIL.n533 VSUBS 0.030544f
C583 VTAIL.n534 VSUBS 0.013683f
C584 VTAIL.n535 VSUBS 0.024048f
C585 VTAIL.n536 VSUBS 0.012923f
C586 VTAIL.n537 VSUBS 0.030544f
C587 VTAIL.n538 VSUBS 0.013683f
C588 VTAIL.n539 VSUBS 0.024048f
C589 VTAIL.n540 VSUBS 0.012923f
C590 VTAIL.n541 VSUBS 0.030544f
C591 VTAIL.n542 VSUBS 0.013683f
C592 VTAIL.n543 VSUBS 1.59668f
C593 VTAIL.n544 VSUBS 0.012923f
C594 VTAIL.t0 VSUBS 0.065423f
C595 VTAIL.n545 VSUBS 0.173494f
C596 VTAIL.n546 VSUBS 0.019431f
C597 VTAIL.n547 VSUBS 0.022908f
C598 VTAIL.n548 VSUBS 0.030544f
C599 VTAIL.n549 VSUBS 0.013683f
C600 VTAIL.n550 VSUBS 0.012923f
C601 VTAIL.n551 VSUBS 0.024048f
C602 VTAIL.n552 VSUBS 0.024048f
C603 VTAIL.n553 VSUBS 0.012923f
C604 VTAIL.n554 VSUBS 0.013683f
C605 VTAIL.n555 VSUBS 0.030544f
C606 VTAIL.n556 VSUBS 0.030544f
C607 VTAIL.n557 VSUBS 0.013683f
C608 VTAIL.n558 VSUBS 0.012923f
C609 VTAIL.n559 VSUBS 0.024048f
C610 VTAIL.n560 VSUBS 0.024048f
C611 VTAIL.n561 VSUBS 0.012923f
C612 VTAIL.n562 VSUBS 0.013683f
C613 VTAIL.n563 VSUBS 0.030544f
C614 VTAIL.n564 VSUBS 0.030544f
C615 VTAIL.n565 VSUBS 0.013683f
C616 VTAIL.n566 VSUBS 0.012923f
C617 VTAIL.n567 VSUBS 0.024048f
C618 VTAIL.n568 VSUBS 0.024048f
C619 VTAIL.n569 VSUBS 0.012923f
C620 VTAIL.n570 VSUBS 0.013683f
C621 VTAIL.n571 VSUBS 0.030544f
C622 VTAIL.n572 VSUBS 0.030544f
C623 VTAIL.n573 VSUBS 0.013683f
C624 VTAIL.n574 VSUBS 0.012923f
C625 VTAIL.n575 VSUBS 0.024048f
C626 VTAIL.n576 VSUBS 0.024048f
C627 VTAIL.n577 VSUBS 0.012923f
C628 VTAIL.n578 VSUBS 0.013683f
C629 VTAIL.n579 VSUBS 0.030544f
C630 VTAIL.n580 VSUBS 0.030544f
C631 VTAIL.n581 VSUBS 0.013683f
C632 VTAIL.n582 VSUBS 0.012923f
C633 VTAIL.n583 VSUBS 0.024048f
C634 VTAIL.n584 VSUBS 0.024048f
C635 VTAIL.n585 VSUBS 0.012923f
C636 VTAIL.n586 VSUBS 0.013683f
C637 VTAIL.n587 VSUBS 0.030544f
C638 VTAIL.n588 VSUBS 0.030544f
C639 VTAIL.n589 VSUBS 0.013683f
C640 VTAIL.n590 VSUBS 0.012923f
C641 VTAIL.n591 VSUBS 0.024048f
C642 VTAIL.n592 VSUBS 0.024048f
C643 VTAIL.n593 VSUBS 0.012923f
C644 VTAIL.n594 VSUBS 0.013683f
C645 VTAIL.n595 VSUBS 0.030544f
C646 VTAIL.n596 VSUBS 0.074991f
C647 VTAIL.n597 VSUBS 0.013683f
C648 VTAIL.n598 VSUBS 0.012923f
C649 VTAIL.n599 VSUBS 0.062158f
C650 VTAIL.n600 VSUBS 0.037951f
C651 VTAIL.n601 VSUBS 1.49056f
C652 VTAIL.n602 VSUBS 0.026731f
C653 VTAIL.n603 VSUBS 0.024048f
C654 VTAIL.n604 VSUBS 0.012923f
C655 VTAIL.n605 VSUBS 0.030544f
C656 VTAIL.n606 VSUBS 0.013303f
C657 VTAIL.n607 VSUBS 0.024048f
C658 VTAIL.n608 VSUBS 0.013683f
C659 VTAIL.n609 VSUBS 0.030544f
C660 VTAIL.n610 VSUBS 0.013683f
C661 VTAIL.n611 VSUBS 0.024048f
C662 VTAIL.n612 VSUBS 0.012923f
C663 VTAIL.n613 VSUBS 0.030544f
C664 VTAIL.n614 VSUBS 0.013683f
C665 VTAIL.n615 VSUBS 0.024048f
C666 VTAIL.n616 VSUBS 0.012923f
C667 VTAIL.n617 VSUBS 0.030544f
C668 VTAIL.n618 VSUBS 0.013683f
C669 VTAIL.n619 VSUBS 0.024048f
C670 VTAIL.n620 VSUBS 0.012923f
C671 VTAIL.n621 VSUBS 0.030544f
C672 VTAIL.n622 VSUBS 0.013683f
C673 VTAIL.n623 VSUBS 0.024048f
C674 VTAIL.n624 VSUBS 0.012923f
C675 VTAIL.n625 VSUBS 0.030544f
C676 VTAIL.n626 VSUBS 0.013683f
C677 VTAIL.n627 VSUBS 1.59668f
C678 VTAIL.n628 VSUBS 0.012923f
C679 VTAIL.t4 VSUBS 0.065423f
C680 VTAIL.n629 VSUBS 0.173494f
C681 VTAIL.n630 VSUBS 0.019431f
C682 VTAIL.n631 VSUBS 0.022908f
C683 VTAIL.n632 VSUBS 0.030544f
C684 VTAIL.n633 VSUBS 0.013683f
C685 VTAIL.n634 VSUBS 0.012923f
C686 VTAIL.n635 VSUBS 0.024048f
C687 VTAIL.n636 VSUBS 0.024048f
C688 VTAIL.n637 VSUBS 0.012923f
C689 VTAIL.n638 VSUBS 0.013683f
C690 VTAIL.n639 VSUBS 0.030544f
C691 VTAIL.n640 VSUBS 0.030544f
C692 VTAIL.n641 VSUBS 0.013683f
C693 VTAIL.n642 VSUBS 0.012923f
C694 VTAIL.n643 VSUBS 0.024048f
C695 VTAIL.n644 VSUBS 0.024048f
C696 VTAIL.n645 VSUBS 0.012923f
C697 VTAIL.n646 VSUBS 0.013683f
C698 VTAIL.n647 VSUBS 0.030544f
C699 VTAIL.n648 VSUBS 0.030544f
C700 VTAIL.n649 VSUBS 0.013683f
C701 VTAIL.n650 VSUBS 0.012923f
C702 VTAIL.n651 VSUBS 0.024048f
C703 VTAIL.n652 VSUBS 0.024048f
C704 VTAIL.n653 VSUBS 0.012923f
C705 VTAIL.n654 VSUBS 0.013683f
C706 VTAIL.n655 VSUBS 0.030544f
C707 VTAIL.n656 VSUBS 0.030544f
C708 VTAIL.n657 VSUBS 0.013683f
C709 VTAIL.n658 VSUBS 0.012923f
C710 VTAIL.n659 VSUBS 0.024048f
C711 VTAIL.n660 VSUBS 0.024048f
C712 VTAIL.n661 VSUBS 0.012923f
C713 VTAIL.n662 VSUBS 0.013683f
C714 VTAIL.n663 VSUBS 0.030544f
C715 VTAIL.n664 VSUBS 0.030544f
C716 VTAIL.n665 VSUBS 0.013683f
C717 VTAIL.n666 VSUBS 0.012923f
C718 VTAIL.n667 VSUBS 0.024048f
C719 VTAIL.n668 VSUBS 0.024048f
C720 VTAIL.n669 VSUBS 0.012923f
C721 VTAIL.n670 VSUBS 0.012923f
C722 VTAIL.n671 VSUBS 0.013683f
C723 VTAIL.n672 VSUBS 0.030544f
C724 VTAIL.n673 VSUBS 0.030544f
C725 VTAIL.n674 VSUBS 0.030544f
C726 VTAIL.n675 VSUBS 0.013303f
C727 VTAIL.n676 VSUBS 0.012923f
C728 VTAIL.n677 VSUBS 0.024048f
C729 VTAIL.n678 VSUBS 0.024048f
C730 VTAIL.n679 VSUBS 0.012923f
C731 VTAIL.n680 VSUBS 0.013683f
C732 VTAIL.n681 VSUBS 0.030544f
C733 VTAIL.n682 VSUBS 0.074991f
C734 VTAIL.n683 VSUBS 0.013683f
C735 VTAIL.n684 VSUBS 0.012923f
C736 VTAIL.n685 VSUBS 0.062158f
C737 VTAIL.n686 VSUBS 0.037951f
C738 VTAIL.n687 VSUBS 1.461f
C739 VDD2.t3 VSUBS 0.381786f
C740 VDD2.t1 VSUBS 0.381786f
C741 VDD2.n0 VSUBS 3.9486f
C742 VDD2.t2 VSUBS 0.381786f
C743 VDD2.t0 VSUBS 0.381786f
C744 VDD2.n1 VSUBS 3.13142f
C745 VDD2.n2 VSUBS 4.82146f
C746 VN.t0 VSUBS 1.27368f
C747 VN.t3 VSUBS 1.27367f
C748 VN.n0 VSUBS 0.965033f
C749 VN.t1 VSUBS 1.27368f
C750 VN.t2 VSUBS 1.27367f
C751 VN.n1 VSUBS 2.08129f
C752 B.n0 VSUBS 0.007305f
C753 B.n1 VSUBS 0.007305f
C754 B.n2 VSUBS 0.010804f
C755 B.n3 VSUBS 0.008279f
C756 B.n4 VSUBS 0.008279f
C757 B.n5 VSUBS 0.008279f
C758 B.n6 VSUBS 0.008279f
C759 B.n7 VSUBS 0.008279f
C760 B.n8 VSUBS 0.008279f
C761 B.n9 VSUBS 0.020455f
C762 B.n10 VSUBS 0.008279f
C763 B.n11 VSUBS 0.008279f
C764 B.n12 VSUBS 0.008279f
C765 B.n13 VSUBS 0.008279f
C766 B.n14 VSUBS 0.008279f
C767 B.n15 VSUBS 0.008279f
C768 B.n16 VSUBS 0.008279f
C769 B.n17 VSUBS 0.008279f
C770 B.n18 VSUBS 0.008279f
C771 B.n19 VSUBS 0.008279f
C772 B.n20 VSUBS 0.008279f
C773 B.n21 VSUBS 0.008279f
C774 B.n22 VSUBS 0.008279f
C775 B.n23 VSUBS 0.008279f
C776 B.n24 VSUBS 0.008279f
C777 B.n25 VSUBS 0.008279f
C778 B.n26 VSUBS 0.008279f
C779 B.n27 VSUBS 0.008279f
C780 B.n28 VSUBS 0.008279f
C781 B.n29 VSUBS 0.008279f
C782 B.n30 VSUBS 0.008279f
C783 B.n31 VSUBS 0.008279f
C784 B.n32 VSUBS 0.008279f
C785 B.n33 VSUBS 0.008279f
C786 B.n34 VSUBS 0.008279f
C787 B.n35 VSUBS 0.008279f
C788 B.t10 VSUBS 0.346571f
C789 B.t11 VSUBS 0.357152f
C790 B.t9 VSUBS 0.305211f
C791 B.n36 VSUBS 0.416851f
C792 B.n37 VSUBS 0.342506f
C793 B.n38 VSUBS 0.008279f
C794 B.n39 VSUBS 0.008279f
C795 B.n40 VSUBS 0.008279f
C796 B.n41 VSUBS 0.008279f
C797 B.t7 VSUBS 0.346575f
C798 B.t8 VSUBS 0.357156f
C799 B.t6 VSUBS 0.305222f
C800 B.n42 VSUBS 0.416833f
C801 B.n43 VSUBS 0.342502f
C802 B.n44 VSUBS 0.019182f
C803 B.n45 VSUBS 0.008279f
C804 B.n46 VSUBS 0.008279f
C805 B.n47 VSUBS 0.008279f
C806 B.n48 VSUBS 0.008279f
C807 B.n49 VSUBS 0.008279f
C808 B.n50 VSUBS 0.008279f
C809 B.n51 VSUBS 0.008279f
C810 B.n52 VSUBS 0.008279f
C811 B.n53 VSUBS 0.008279f
C812 B.n54 VSUBS 0.008279f
C813 B.n55 VSUBS 0.008279f
C814 B.n56 VSUBS 0.008279f
C815 B.n57 VSUBS 0.008279f
C816 B.n58 VSUBS 0.008279f
C817 B.n59 VSUBS 0.008279f
C818 B.n60 VSUBS 0.008279f
C819 B.n61 VSUBS 0.008279f
C820 B.n62 VSUBS 0.008279f
C821 B.n63 VSUBS 0.008279f
C822 B.n64 VSUBS 0.008279f
C823 B.n65 VSUBS 0.008279f
C824 B.n66 VSUBS 0.008279f
C825 B.n67 VSUBS 0.008279f
C826 B.n68 VSUBS 0.008279f
C827 B.n69 VSUBS 0.008279f
C828 B.n70 VSUBS 0.020455f
C829 B.n71 VSUBS 0.008279f
C830 B.n72 VSUBS 0.008279f
C831 B.n73 VSUBS 0.008279f
C832 B.n74 VSUBS 0.008279f
C833 B.n75 VSUBS 0.008279f
C834 B.n76 VSUBS 0.008279f
C835 B.n77 VSUBS 0.008279f
C836 B.n78 VSUBS 0.008279f
C837 B.n79 VSUBS 0.008279f
C838 B.n80 VSUBS 0.008279f
C839 B.n81 VSUBS 0.008279f
C840 B.n82 VSUBS 0.008279f
C841 B.n83 VSUBS 0.008279f
C842 B.n84 VSUBS 0.008279f
C843 B.n85 VSUBS 0.018992f
C844 B.n86 VSUBS 0.008279f
C845 B.n87 VSUBS 0.008279f
C846 B.n88 VSUBS 0.008279f
C847 B.n89 VSUBS 0.008279f
C848 B.n90 VSUBS 0.008279f
C849 B.n91 VSUBS 0.008279f
C850 B.n92 VSUBS 0.008279f
C851 B.n93 VSUBS 0.008279f
C852 B.n94 VSUBS 0.008279f
C853 B.n95 VSUBS 0.008279f
C854 B.n96 VSUBS 0.008279f
C855 B.n97 VSUBS 0.008279f
C856 B.n98 VSUBS 0.008279f
C857 B.n99 VSUBS 0.008279f
C858 B.n100 VSUBS 0.008279f
C859 B.n101 VSUBS 0.008279f
C860 B.n102 VSUBS 0.008279f
C861 B.n103 VSUBS 0.008279f
C862 B.n104 VSUBS 0.008279f
C863 B.n105 VSUBS 0.008279f
C864 B.n106 VSUBS 0.008279f
C865 B.n107 VSUBS 0.008279f
C866 B.n108 VSUBS 0.008279f
C867 B.n109 VSUBS 0.008279f
C868 B.n110 VSUBS 0.008279f
C869 B.n111 VSUBS 0.008279f
C870 B.t5 VSUBS 0.346575f
C871 B.t4 VSUBS 0.357156f
C872 B.t3 VSUBS 0.305222f
C873 B.n112 VSUBS 0.416833f
C874 B.n113 VSUBS 0.342502f
C875 B.n114 VSUBS 0.008279f
C876 B.n115 VSUBS 0.008279f
C877 B.n116 VSUBS 0.008279f
C878 B.n117 VSUBS 0.008279f
C879 B.n118 VSUBS 0.004566f
C880 B.n119 VSUBS 0.008279f
C881 B.n120 VSUBS 0.008279f
C882 B.n121 VSUBS 0.008279f
C883 B.n122 VSUBS 0.008279f
C884 B.n123 VSUBS 0.008279f
C885 B.n124 VSUBS 0.008279f
C886 B.n125 VSUBS 0.008279f
C887 B.n126 VSUBS 0.008279f
C888 B.n127 VSUBS 0.008279f
C889 B.n128 VSUBS 0.008279f
C890 B.n129 VSUBS 0.008279f
C891 B.n130 VSUBS 0.008279f
C892 B.n131 VSUBS 0.008279f
C893 B.n132 VSUBS 0.008279f
C894 B.n133 VSUBS 0.008279f
C895 B.n134 VSUBS 0.008279f
C896 B.n135 VSUBS 0.008279f
C897 B.n136 VSUBS 0.008279f
C898 B.n137 VSUBS 0.008279f
C899 B.n138 VSUBS 0.008279f
C900 B.n139 VSUBS 0.008279f
C901 B.n140 VSUBS 0.008279f
C902 B.n141 VSUBS 0.008279f
C903 B.n142 VSUBS 0.008279f
C904 B.n143 VSUBS 0.008279f
C905 B.n144 VSUBS 0.020455f
C906 B.n145 VSUBS 0.008279f
C907 B.n146 VSUBS 0.008279f
C908 B.n147 VSUBS 0.008279f
C909 B.n148 VSUBS 0.008279f
C910 B.n149 VSUBS 0.008279f
C911 B.n150 VSUBS 0.008279f
C912 B.n151 VSUBS 0.008279f
C913 B.n152 VSUBS 0.008279f
C914 B.n153 VSUBS 0.008279f
C915 B.n154 VSUBS 0.008279f
C916 B.n155 VSUBS 0.008279f
C917 B.n156 VSUBS 0.008279f
C918 B.n157 VSUBS 0.008279f
C919 B.n158 VSUBS 0.008279f
C920 B.n159 VSUBS 0.008279f
C921 B.n160 VSUBS 0.008279f
C922 B.n161 VSUBS 0.008279f
C923 B.n162 VSUBS 0.008279f
C924 B.n163 VSUBS 0.008279f
C925 B.n164 VSUBS 0.008279f
C926 B.n165 VSUBS 0.008279f
C927 B.n166 VSUBS 0.008279f
C928 B.n167 VSUBS 0.008279f
C929 B.n168 VSUBS 0.008279f
C930 B.n169 VSUBS 0.018992f
C931 B.n170 VSUBS 0.018992f
C932 B.n171 VSUBS 0.020455f
C933 B.n172 VSUBS 0.008279f
C934 B.n173 VSUBS 0.008279f
C935 B.n174 VSUBS 0.008279f
C936 B.n175 VSUBS 0.008279f
C937 B.n176 VSUBS 0.008279f
C938 B.n177 VSUBS 0.008279f
C939 B.n178 VSUBS 0.008279f
C940 B.n179 VSUBS 0.008279f
C941 B.n180 VSUBS 0.008279f
C942 B.n181 VSUBS 0.008279f
C943 B.n182 VSUBS 0.008279f
C944 B.n183 VSUBS 0.008279f
C945 B.n184 VSUBS 0.008279f
C946 B.n185 VSUBS 0.008279f
C947 B.n186 VSUBS 0.008279f
C948 B.n187 VSUBS 0.008279f
C949 B.n188 VSUBS 0.008279f
C950 B.n189 VSUBS 0.008279f
C951 B.n190 VSUBS 0.008279f
C952 B.n191 VSUBS 0.008279f
C953 B.n192 VSUBS 0.008279f
C954 B.n193 VSUBS 0.008279f
C955 B.n194 VSUBS 0.008279f
C956 B.n195 VSUBS 0.008279f
C957 B.n196 VSUBS 0.008279f
C958 B.n197 VSUBS 0.008279f
C959 B.n198 VSUBS 0.008279f
C960 B.n199 VSUBS 0.008279f
C961 B.n200 VSUBS 0.008279f
C962 B.n201 VSUBS 0.008279f
C963 B.n202 VSUBS 0.008279f
C964 B.n203 VSUBS 0.008279f
C965 B.n204 VSUBS 0.008279f
C966 B.n205 VSUBS 0.008279f
C967 B.n206 VSUBS 0.008279f
C968 B.n207 VSUBS 0.008279f
C969 B.n208 VSUBS 0.008279f
C970 B.n209 VSUBS 0.008279f
C971 B.n210 VSUBS 0.008279f
C972 B.n211 VSUBS 0.008279f
C973 B.n212 VSUBS 0.008279f
C974 B.n213 VSUBS 0.008279f
C975 B.n214 VSUBS 0.008279f
C976 B.n215 VSUBS 0.008279f
C977 B.n216 VSUBS 0.008279f
C978 B.n217 VSUBS 0.008279f
C979 B.n218 VSUBS 0.008279f
C980 B.n219 VSUBS 0.008279f
C981 B.n220 VSUBS 0.008279f
C982 B.n221 VSUBS 0.008279f
C983 B.n222 VSUBS 0.008279f
C984 B.n223 VSUBS 0.008279f
C985 B.n224 VSUBS 0.008279f
C986 B.n225 VSUBS 0.008279f
C987 B.n226 VSUBS 0.008279f
C988 B.n227 VSUBS 0.008279f
C989 B.n228 VSUBS 0.008279f
C990 B.n229 VSUBS 0.008279f
C991 B.n230 VSUBS 0.008279f
C992 B.n231 VSUBS 0.008279f
C993 B.n232 VSUBS 0.008279f
C994 B.n233 VSUBS 0.008279f
C995 B.n234 VSUBS 0.008279f
C996 B.n235 VSUBS 0.008279f
C997 B.n236 VSUBS 0.008279f
C998 B.n237 VSUBS 0.008279f
C999 B.n238 VSUBS 0.008279f
C1000 B.n239 VSUBS 0.008279f
C1001 B.n240 VSUBS 0.008279f
C1002 B.n241 VSUBS 0.008279f
C1003 B.n242 VSUBS 0.008279f
C1004 B.n243 VSUBS 0.008279f
C1005 B.n244 VSUBS 0.008279f
C1006 B.n245 VSUBS 0.008279f
C1007 B.n246 VSUBS 0.008279f
C1008 B.t2 VSUBS 0.346571f
C1009 B.t1 VSUBS 0.357152f
C1010 B.t0 VSUBS 0.305211f
C1011 B.n247 VSUBS 0.416851f
C1012 B.n248 VSUBS 0.342506f
C1013 B.n249 VSUBS 0.019182f
C1014 B.n250 VSUBS 0.007853f
C1015 B.n251 VSUBS 0.008279f
C1016 B.n252 VSUBS 0.008279f
C1017 B.n253 VSUBS 0.008279f
C1018 B.n254 VSUBS 0.008279f
C1019 B.n255 VSUBS 0.008279f
C1020 B.n256 VSUBS 0.008279f
C1021 B.n257 VSUBS 0.008279f
C1022 B.n258 VSUBS 0.008279f
C1023 B.n259 VSUBS 0.008279f
C1024 B.n260 VSUBS 0.008279f
C1025 B.n261 VSUBS 0.008279f
C1026 B.n262 VSUBS 0.008279f
C1027 B.n263 VSUBS 0.008279f
C1028 B.n264 VSUBS 0.008279f
C1029 B.n265 VSUBS 0.008279f
C1030 B.n266 VSUBS 0.004566f
C1031 B.n267 VSUBS 0.019182f
C1032 B.n268 VSUBS 0.007853f
C1033 B.n269 VSUBS 0.008279f
C1034 B.n270 VSUBS 0.008279f
C1035 B.n271 VSUBS 0.008279f
C1036 B.n272 VSUBS 0.008279f
C1037 B.n273 VSUBS 0.008279f
C1038 B.n274 VSUBS 0.008279f
C1039 B.n275 VSUBS 0.008279f
C1040 B.n276 VSUBS 0.008279f
C1041 B.n277 VSUBS 0.008279f
C1042 B.n278 VSUBS 0.008279f
C1043 B.n279 VSUBS 0.008279f
C1044 B.n280 VSUBS 0.008279f
C1045 B.n281 VSUBS 0.008279f
C1046 B.n282 VSUBS 0.008279f
C1047 B.n283 VSUBS 0.008279f
C1048 B.n284 VSUBS 0.008279f
C1049 B.n285 VSUBS 0.008279f
C1050 B.n286 VSUBS 0.008279f
C1051 B.n287 VSUBS 0.008279f
C1052 B.n288 VSUBS 0.008279f
C1053 B.n289 VSUBS 0.008279f
C1054 B.n290 VSUBS 0.008279f
C1055 B.n291 VSUBS 0.008279f
C1056 B.n292 VSUBS 0.008279f
C1057 B.n293 VSUBS 0.008279f
C1058 B.n294 VSUBS 0.008279f
C1059 B.n295 VSUBS 0.008279f
C1060 B.n296 VSUBS 0.008279f
C1061 B.n297 VSUBS 0.008279f
C1062 B.n298 VSUBS 0.008279f
C1063 B.n299 VSUBS 0.008279f
C1064 B.n300 VSUBS 0.008279f
C1065 B.n301 VSUBS 0.008279f
C1066 B.n302 VSUBS 0.008279f
C1067 B.n303 VSUBS 0.008279f
C1068 B.n304 VSUBS 0.008279f
C1069 B.n305 VSUBS 0.008279f
C1070 B.n306 VSUBS 0.008279f
C1071 B.n307 VSUBS 0.008279f
C1072 B.n308 VSUBS 0.008279f
C1073 B.n309 VSUBS 0.008279f
C1074 B.n310 VSUBS 0.008279f
C1075 B.n311 VSUBS 0.008279f
C1076 B.n312 VSUBS 0.008279f
C1077 B.n313 VSUBS 0.008279f
C1078 B.n314 VSUBS 0.008279f
C1079 B.n315 VSUBS 0.008279f
C1080 B.n316 VSUBS 0.008279f
C1081 B.n317 VSUBS 0.008279f
C1082 B.n318 VSUBS 0.008279f
C1083 B.n319 VSUBS 0.008279f
C1084 B.n320 VSUBS 0.008279f
C1085 B.n321 VSUBS 0.008279f
C1086 B.n322 VSUBS 0.008279f
C1087 B.n323 VSUBS 0.008279f
C1088 B.n324 VSUBS 0.008279f
C1089 B.n325 VSUBS 0.008279f
C1090 B.n326 VSUBS 0.008279f
C1091 B.n327 VSUBS 0.008279f
C1092 B.n328 VSUBS 0.008279f
C1093 B.n329 VSUBS 0.008279f
C1094 B.n330 VSUBS 0.008279f
C1095 B.n331 VSUBS 0.008279f
C1096 B.n332 VSUBS 0.008279f
C1097 B.n333 VSUBS 0.008279f
C1098 B.n334 VSUBS 0.008279f
C1099 B.n335 VSUBS 0.008279f
C1100 B.n336 VSUBS 0.008279f
C1101 B.n337 VSUBS 0.008279f
C1102 B.n338 VSUBS 0.008279f
C1103 B.n339 VSUBS 0.008279f
C1104 B.n340 VSUBS 0.008279f
C1105 B.n341 VSUBS 0.008279f
C1106 B.n342 VSUBS 0.008279f
C1107 B.n343 VSUBS 0.008279f
C1108 B.n344 VSUBS 0.020455f
C1109 B.n345 VSUBS 0.019503f
C1110 B.n346 VSUBS 0.019944f
C1111 B.n347 VSUBS 0.008279f
C1112 B.n348 VSUBS 0.008279f
C1113 B.n349 VSUBS 0.008279f
C1114 B.n350 VSUBS 0.008279f
C1115 B.n351 VSUBS 0.008279f
C1116 B.n352 VSUBS 0.008279f
C1117 B.n353 VSUBS 0.008279f
C1118 B.n354 VSUBS 0.008279f
C1119 B.n355 VSUBS 0.008279f
C1120 B.n356 VSUBS 0.008279f
C1121 B.n357 VSUBS 0.008279f
C1122 B.n358 VSUBS 0.008279f
C1123 B.n359 VSUBS 0.008279f
C1124 B.n360 VSUBS 0.008279f
C1125 B.n361 VSUBS 0.008279f
C1126 B.n362 VSUBS 0.008279f
C1127 B.n363 VSUBS 0.008279f
C1128 B.n364 VSUBS 0.008279f
C1129 B.n365 VSUBS 0.008279f
C1130 B.n366 VSUBS 0.008279f
C1131 B.n367 VSUBS 0.008279f
C1132 B.n368 VSUBS 0.008279f
C1133 B.n369 VSUBS 0.008279f
C1134 B.n370 VSUBS 0.008279f
C1135 B.n371 VSUBS 0.008279f
C1136 B.n372 VSUBS 0.008279f
C1137 B.n373 VSUBS 0.008279f
C1138 B.n374 VSUBS 0.008279f
C1139 B.n375 VSUBS 0.008279f
C1140 B.n376 VSUBS 0.008279f
C1141 B.n377 VSUBS 0.008279f
C1142 B.n378 VSUBS 0.008279f
C1143 B.n379 VSUBS 0.008279f
C1144 B.n380 VSUBS 0.008279f
C1145 B.n381 VSUBS 0.008279f
C1146 B.n382 VSUBS 0.008279f
C1147 B.n383 VSUBS 0.008279f
C1148 B.n384 VSUBS 0.008279f
C1149 B.n385 VSUBS 0.008279f
C1150 B.n386 VSUBS 0.008279f
C1151 B.n387 VSUBS 0.008279f
C1152 B.n388 VSUBS 0.008279f
C1153 B.n389 VSUBS 0.018992f
C1154 B.n390 VSUBS 0.018992f
C1155 B.n391 VSUBS 0.020455f
C1156 B.n392 VSUBS 0.008279f
C1157 B.n393 VSUBS 0.008279f
C1158 B.n394 VSUBS 0.008279f
C1159 B.n395 VSUBS 0.008279f
C1160 B.n396 VSUBS 0.008279f
C1161 B.n397 VSUBS 0.008279f
C1162 B.n398 VSUBS 0.008279f
C1163 B.n399 VSUBS 0.008279f
C1164 B.n400 VSUBS 0.008279f
C1165 B.n401 VSUBS 0.008279f
C1166 B.n402 VSUBS 0.008279f
C1167 B.n403 VSUBS 0.008279f
C1168 B.n404 VSUBS 0.008279f
C1169 B.n405 VSUBS 0.008279f
C1170 B.n406 VSUBS 0.008279f
C1171 B.n407 VSUBS 0.008279f
C1172 B.n408 VSUBS 0.008279f
C1173 B.n409 VSUBS 0.008279f
C1174 B.n410 VSUBS 0.008279f
C1175 B.n411 VSUBS 0.008279f
C1176 B.n412 VSUBS 0.008279f
C1177 B.n413 VSUBS 0.008279f
C1178 B.n414 VSUBS 0.008279f
C1179 B.n415 VSUBS 0.008279f
C1180 B.n416 VSUBS 0.008279f
C1181 B.n417 VSUBS 0.008279f
C1182 B.n418 VSUBS 0.008279f
C1183 B.n419 VSUBS 0.008279f
C1184 B.n420 VSUBS 0.008279f
C1185 B.n421 VSUBS 0.008279f
C1186 B.n422 VSUBS 0.008279f
C1187 B.n423 VSUBS 0.008279f
C1188 B.n424 VSUBS 0.008279f
C1189 B.n425 VSUBS 0.008279f
C1190 B.n426 VSUBS 0.008279f
C1191 B.n427 VSUBS 0.008279f
C1192 B.n428 VSUBS 0.008279f
C1193 B.n429 VSUBS 0.008279f
C1194 B.n430 VSUBS 0.008279f
C1195 B.n431 VSUBS 0.008279f
C1196 B.n432 VSUBS 0.008279f
C1197 B.n433 VSUBS 0.008279f
C1198 B.n434 VSUBS 0.008279f
C1199 B.n435 VSUBS 0.008279f
C1200 B.n436 VSUBS 0.008279f
C1201 B.n437 VSUBS 0.008279f
C1202 B.n438 VSUBS 0.008279f
C1203 B.n439 VSUBS 0.008279f
C1204 B.n440 VSUBS 0.008279f
C1205 B.n441 VSUBS 0.008279f
C1206 B.n442 VSUBS 0.008279f
C1207 B.n443 VSUBS 0.008279f
C1208 B.n444 VSUBS 0.008279f
C1209 B.n445 VSUBS 0.008279f
C1210 B.n446 VSUBS 0.008279f
C1211 B.n447 VSUBS 0.008279f
C1212 B.n448 VSUBS 0.008279f
C1213 B.n449 VSUBS 0.008279f
C1214 B.n450 VSUBS 0.008279f
C1215 B.n451 VSUBS 0.008279f
C1216 B.n452 VSUBS 0.008279f
C1217 B.n453 VSUBS 0.008279f
C1218 B.n454 VSUBS 0.008279f
C1219 B.n455 VSUBS 0.008279f
C1220 B.n456 VSUBS 0.008279f
C1221 B.n457 VSUBS 0.008279f
C1222 B.n458 VSUBS 0.008279f
C1223 B.n459 VSUBS 0.008279f
C1224 B.n460 VSUBS 0.008279f
C1225 B.n461 VSUBS 0.008279f
C1226 B.n462 VSUBS 0.008279f
C1227 B.n463 VSUBS 0.008279f
C1228 B.n464 VSUBS 0.008279f
C1229 B.n465 VSUBS 0.008279f
C1230 B.n466 VSUBS 0.008279f
C1231 B.n467 VSUBS 0.007853f
C1232 B.n468 VSUBS 0.008279f
C1233 B.n469 VSUBS 0.008279f
C1234 B.n470 VSUBS 0.004566f
C1235 B.n471 VSUBS 0.008279f
C1236 B.n472 VSUBS 0.008279f
C1237 B.n473 VSUBS 0.008279f
C1238 B.n474 VSUBS 0.008279f
C1239 B.n475 VSUBS 0.008279f
C1240 B.n476 VSUBS 0.008279f
C1241 B.n477 VSUBS 0.008279f
C1242 B.n478 VSUBS 0.008279f
C1243 B.n479 VSUBS 0.008279f
C1244 B.n480 VSUBS 0.008279f
C1245 B.n481 VSUBS 0.008279f
C1246 B.n482 VSUBS 0.008279f
C1247 B.n483 VSUBS 0.004566f
C1248 B.n484 VSUBS 0.019182f
C1249 B.n485 VSUBS 0.007853f
C1250 B.n486 VSUBS 0.008279f
C1251 B.n487 VSUBS 0.008279f
C1252 B.n488 VSUBS 0.008279f
C1253 B.n489 VSUBS 0.008279f
C1254 B.n490 VSUBS 0.008279f
C1255 B.n491 VSUBS 0.008279f
C1256 B.n492 VSUBS 0.008279f
C1257 B.n493 VSUBS 0.008279f
C1258 B.n494 VSUBS 0.008279f
C1259 B.n495 VSUBS 0.008279f
C1260 B.n496 VSUBS 0.008279f
C1261 B.n497 VSUBS 0.008279f
C1262 B.n498 VSUBS 0.008279f
C1263 B.n499 VSUBS 0.008279f
C1264 B.n500 VSUBS 0.008279f
C1265 B.n501 VSUBS 0.008279f
C1266 B.n502 VSUBS 0.008279f
C1267 B.n503 VSUBS 0.008279f
C1268 B.n504 VSUBS 0.008279f
C1269 B.n505 VSUBS 0.008279f
C1270 B.n506 VSUBS 0.008279f
C1271 B.n507 VSUBS 0.008279f
C1272 B.n508 VSUBS 0.008279f
C1273 B.n509 VSUBS 0.008279f
C1274 B.n510 VSUBS 0.008279f
C1275 B.n511 VSUBS 0.008279f
C1276 B.n512 VSUBS 0.008279f
C1277 B.n513 VSUBS 0.008279f
C1278 B.n514 VSUBS 0.008279f
C1279 B.n515 VSUBS 0.008279f
C1280 B.n516 VSUBS 0.008279f
C1281 B.n517 VSUBS 0.008279f
C1282 B.n518 VSUBS 0.008279f
C1283 B.n519 VSUBS 0.008279f
C1284 B.n520 VSUBS 0.008279f
C1285 B.n521 VSUBS 0.008279f
C1286 B.n522 VSUBS 0.008279f
C1287 B.n523 VSUBS 0.008279f
C1288 B.n524 VSUBS 0.008279f
C1289 B.n525 VSUBS 0.008279f
C1290 B.n526 VSUBS 0.008279f
C1291 B.n527 VSUBS 0.008279f
C1292 B.n528 VSUBS 0.008279f
C1293 B.n529 VSUBS 0.008279f
C1294 B.n530 VSUBS 0.008279f
C1295 B.n531 VSUBS 0.008279f
C1296 B.n532 VSUBS 0.008279f
C1297 B.n533 VSUBS 0.008279f
C1298 B.n534 VSUBS 0.008279f
C1299 B.n535 VSUBS 0.008279f
C1300 B.n536 VSUBS 0.008279f
C1301 B.n537 VSUBS 0.008279f
C1302 B.n538 VSUBS 0.008279f
C1303 B.n539 VSUBS 0.008279f
C1304 B.n540 VSUBS 0.008279f
C1305 B.n541 VSUBS 0.008279f
C1306 B.n542 VSUBS 0.008279f
C1307 B.n543 VSUBS 0.008279f
C1308 B.n544 VSUBS 0.008279f
C1309 B.n545 VSUBS 0.008279f
C1310 B.n546 VSUBS 0.008279f
C1311 B.n547 VSUBS 0.008279f
C1312 B.n548 VSUBS 0.008279f
C1313 B.n549 VSUBS 0.008279f
C1314 B.n550 VSUBS 0.008279f
C1315 B.n551 VSUBS 0.008279f
C1316 B.n552 VSUBS 0.008279f
C1317 B.n553 VSUBS 0.008279f
C1318 B.n554 VSUBS 0.008279f
C1319 B.n555 VSUBS 0.008279f
C1320 B.n556 VSUBS 0.008279f
C1321 B.n557 VSUBS 0.008279f
C1322 B.n558 VSUBS 0.008279f
C1323 B.n559 VSUBS 0.008279f
C1324 B.n560 VSUBS 0.008279f
C1325 B.n561 VSUBS 0.008279f
C1326 B.n562 VSUBS 0.020455f
C1327 B.n563 VSUBS 0.018992f
C1328 B.n564 VSUBS 0.018992f
C1329 B.n565 VSUBS 0.008279f
C1330 B.n566 VSUBS 0.008279f
C1331 B.n567 VSUBS 0.008279f
C1332 B.n568 VSUBS 0.008279f
C1333 B.n569 VSUBS 0.008279f
C1334 B.n570 VSUBS 0.008279f
C1335 B.n571 VSUBS 0.008279f
C1336 B.n572 VSUBS 0.008279f
C1337 B.n573 VSUBS 0.008279f
C1338 B.n574 VSUBS 0.008279f
C1339 B.n575 VSUBS 0.008279f
C1340 B.n576 VSUBS 0.008279f
C1341 B.n577 VSUBS 0.008279f
C1342 B.n578 VSUBS 0.008279f
C1343 B.n579 VSUBS 0.008279f
C1344 B.n580 VSUBS 0.008279f
C1345 B.n581 VSUBS 0.008279f
C1346 B.n582 VSUBS 0.008279f
C1347 B.n583 VSUBS 0.010804f
C1348 B.n584 VSUBS 0.011509f
C1349 B.n585 VSUBS 0.022886f
.ends

