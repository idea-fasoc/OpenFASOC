* NGSPICE file created from diff_pair_sample_0873.ext - technology: sky130A

.subckt diff_pair_sample_0873 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t11 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=6.6456 pd=34.86 as=2.8116 ps=17.37 w=17.04 l=3.83
X1 VDD2.t9 VN.t0 VTAIL.t7 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=6.6456 pd=34.86 as=2.8116 ps=17.37 w=17.04 l=3.83
X2 VDD1.t8 VP.t1 VTAIL.t14 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=2.8116 pd=17.37 as=2.8116 ps=17.37 w=17.04 l=3.83
X3 VTAIL.t5 VN.t1 VDD2.t8 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=2.8116 pd=17.37 as=2.8116 ps=17.37 w=17.04 l=3.83
X4 VTAIL.t2 VN.t2 VDD2.t7 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=2.8116 pd=17.37 as=2.8116 ps=17.37 w=17.04 l=3.83
X5 VTAIL.t13 VP.t2 VDD1.t7 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=2.8116 pd=17.37 as=2.8116 ps=17.37 w=17.04 l=3.83
X6 VDD2.t6 VN.t3 VTAIL.t8 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=6.6456 pd=34.86 as=2.8116 ps=17.37 w=17.04 l=3.83
X7 VDD2.t5 VN.t4 VTAIL.t1 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=2.8116 pd=17.37 as=2.8116 ps=17.37 w=17.04 l=3.83
X8 VDD1.t6 VP.t3 VTAIL.t15 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=2.8116 pd=17.37 as=6.6456 ps=34.86 w=17.04 l=3.83
X9 VTAIL.t16 VP.t4 VDD1.t5 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=2.8116 pd=17.37 as=2.8116 ps=17.37 w=17.04 l=3.83
X10 VTAIL.t12 VP.t5 VDD1.t4 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=2.8116 pd=17.37 as=2.8116 ps=17.37 w=17.04 l=3.83
X11 VTAIL.t18 VP.t6 VDD1.t3 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=2.8116 pd=17.37 as=2.8116 ps=17.37 w=17.04 l=3.83
X12 VDD2.t4 VN.t5 VTAIL.t6 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=2.8116 pd=17.37 as=6.6456 ps=34.86 w=17.04 l=3.83
X13 B.t11 B.t9 B.t10 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=6.6456 pd=34.86 as=0 ps=0 w=17.04 l=3.83
X14 VDD1.t2 VP.t7 VTAIL.t10 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=2.8116 pd=17.37 as=6.6456 ps=34.86 w=17.04 l=3.83
X15 VDD1.t1 VP.t8 VTAIL.t17 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=2.8116 pd=17.37 as=2.8116 ps=17.37 w=17.04 l=3.83
X16 VTAIL.t19 VN.t6 VDD2.t3 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=2.8116 pd=17.37 as=2.8116 ps=17.37 w=17.04 l=3.83
X17 VDD2.t2 VN.t7 VTAIL.t4 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=2.8116 pd=17.37 as=2.8116 ps=17.37 w=17.04 l=3.83
X18 B.t8 B.t6 B.t7 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=6.6456 pd=34.86 as=0 ps=0 w=17.04 l=3.83
X19 VDD2.t1 VN.t8 VTAIL.t3 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=2.8116 pd=17.37 as=6.6456 ps=34.86 w=17.04 l=3.83
X20 B.t5 B.t3 B.t4 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=6.6456 pd=34.86 as=0 ps=0 w=17.04 l=3.83
X21 VTAIL.t0 VN.t9 VDD2.t0 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=2.8116 pd=17.37 as=2.8116 ps=17.37 w=17.04 l=3.83
X22 VDD1.t0 VP.t9 VTAIL.t9 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=6.6456 pd=34.86 as=2.8116 ps=17.37 w=17.04 l=3.83
X23 B.t2 B.t0 B.t1 w_n5962_n4376# sky130_fd_pr__pfet_01v8 ad=6.6456 pd=34.86 as=0 ps=0 w=17.04 l=3.83
R0 VP.n34 VP.n33 161.3
R1 VP.n35 VP.n30 161.3
R2 VP.n37 VP.n36 161.3
R3 VP.n38 VP.n29 161.3
R4 VP.n40 VP.n39 161.3
R5 VP.n41 VP.n28 161.3
R6 VP.n43 VP.n42 161.3
R7 VP.n44 VP.n27 161.3
R8 VP.n47 VP.n46 161.3
R9 VP.n48 VP.n26 161.3
R10 VP.n50 VP.n49 161.3
R11 VP.n51 VP.n25 161.3
R12 VP.n53 VP.n52 161.3
R13 VP.n54 VP.n24 161.3
R14 VP.n56 VP.n55 161.3
R15 VP.n57 VP.n23 161.3
R16 VP.n60 VP.n59 161.3
R17 VP.n61 VP.n22 161.3
R18 VP.n63 VP.n62 161.3
R19 VP.n64 VP.n21 161.3
R20 VP.n66 VP.n65 161.3
R21 VP.n67 VP.n20 161.3
R22 VP.n69 VP.n68 161.3
R23 VP.n70 VP.n19 161.3
R24 VP.n72 VP.n71 161.3
R25 VP.n129 VP.n128 161.3
R26 VP.n127 VP.n1 161.3
R27 VP.n126 VP.n125 161.3
R28 VP.n124 VP.n2 161.3
R29 VP.n123 VP.n122 161.3
R30 VP.n121 VP.n3 161.3
R31 VP.n120 VP.n119 161.3
R32 VP.n118 VP.n4 161.3
R33 VP.n117 VP.n116 161.3
R34 VP.n114 VP.n5 161.3
R35 VP.n113 VP.n112 161.3
R36 VP.n111 VP.n6 161.3
R37 VP.n110 VP.n109 161.3
R38 VP.n108 VP.n7 161.3
R39 VP.n107 VP.n106 161.3
R40 VP.n105 VP.n8 161.3
R41 VP.n104 VP.n103 161.3
R42 VP.n101 VP.n9 161.3
R43 VP.n100 VP.n99 161.3
R44 VP.n98 VP.n10 161.3
R45 VP.n97 VP.n96 161.3
R46 VP.n95 VP.n11 161.3
R47 VP.n94 VP.n93 161.3
R48 VP.n92 VP.n12 161.3
R49 VP.n91 VP.n90 161.3
R50 VP.n88 VP.n13 161.3
R51 VP.n87 VP.n86 161.3
R52 VP.n85 VP.n14 161.3
R53 VP.n84 VP.n83 161.3
R54 VP.n82 VP.n15 161.3
R55 VP.n81 VP.n80 161.3
R56 VP.n79 VP.n16 161.3
R57 VP.n78 VP.n77 161.3
R58 VP.n76 VP.n17 161.3
R59 VP.n31 VP.t0 140.311
R60 VP.n75 VP.t9 107.224
R61 VP.n89 VP.t5 107.224
R62 VP.n102 VP.t8 107.224
R63 VP.n115 VP.t6 107.224
R64 VP.n0 VP.t7 107.224
R65 VP.n18 VP.t3 107.224
R66 VP.n58 VP.t4 107.224
R67 VP.n45 VP.t1 107.224
R68 VP.n32 VP.t2 107.224
R69 VP.n75 VP.n74 86.8027
R70 VP.n130 VP.n0 86.8027
R71 VP.n73 VP.n18 86.8027
R72 VP.n74 VP.n73 63.6889
R73 VP.n96 VP.n95 56.5617
R74 VP.n109 VP.n108 56.5617
R75 VP.n52 VP.n51 56.5617
R76 VP.n39 VP.n38 56.5617
R77 VP.n32 VP.n31 55.106
R78 VP.n83 VP.n82 41.5458
R79 VP.n122 VP.n121 41.5458
R80 VP.n65 VP.n64 41.5458
R81 VP.n82 VP.n81 39.6083
R82 VP.n122 VP.n2 39.6083
R83 VP.n65 VP.n20 39.6083
R84 VP.n77 VP.n76 24.5923
R85 VP.n77 VP.n16 24.5923
R86 VP.n81 VP.n16 24.5923
R87 VP.n83 VP.n14 24.5923
R88 VP.n87 VP.n14 24.5923
R89 VP.n88 VP.n87 24.5923
R90 VP.n90 VP.n12 24.5923
R91 VP.n94 VP.n12 24.5923
R92 VP.n95 VP.n94 24.5923
R93 VP.n96 VP.n10 24.5923
R94 VP.n100 VP.n10 24.5923
R95 VP.n101 VP.n100 24.5923
R96 VP.n103 VP.n8 24.5923
R97 VP.n107 VP.n8 24.5923
R98 VP.n108 VP.n107 24.5923
R99 VP.n109 VP.n6 24.5923
R100 VP.n113 VP.n6 24.5923
R101 VP.n114 VP.n113 24.5923
R102 VP.n116 VP.n4 24.5923
R103 VP.n120 VP.n4 24.5923
R104 VP.n121 VP.n120 24.5923
R105 VP.n126 VP.n2 24.5923
R106 VP.n127 VP.n126 24.5923
R107 VP.n128 VP.n127 24.5923
R108 VP.n69 VP.n20 24.5923
R109 VP.n70 VP.n69 24.5923
R110 VP.n71 VP.n70 24.5923
R111 VP.n52 VP.n24 24.5923
R112 VP.n56 VP.n24 24.5923
R113 VP.n57 VP.n56 24.5923
R114 VP.n59 VP.n22 24.5923
R115 VP.n63 VP.n22 24.5923
R116 VP.n64 VP.n63 24.5923
R117 VP.n39 VP.n28 24.5923
R118 VP.n43 VP.n28 24.5923
R119 VP.n44 VP.n43 24.5923
R120 VP.n46 VP.n26 24.5923
R121 VP.n50 VP.n26 24.5923
R122 VP.n51 VP.n50 24.5923
R123 VP.n33 VP.n30 24.5923
R124 VP.n37 VP.n30 24.5923
R125 VP.n38 VP.n37 24.5923
R126 VP.n90 VP.n89 20.1658
R127 VP.n115 VP.n114 20.1658
R128 VP.n58 VP.n57 20.1658
R129 VP.n33 VP.n32 20.1658
R130 VP.n102 VP.n101 12.2964
R131 VP.n103 VP.n102 12.2964
R132 VP.n45 VP.n44 12.2964
R133 VP.n46 VP.n45 12.2964
R134 VP.n89 VP.n88 4.42703
R135 VP.n116 VP.n115 4.42703
R136 VP.n59 VP.n58 4.42703
R137 VP.n76 VP.n75 3.44336
R138 VP.n128 VP.n0 3.44336
R139 VP.n71 VP.n18 3.44336
R140 VP.n34 VP.n31 2.44068
R141 VP.n73 VP.n72 0.354861
R142 VP.n74 VP.n17 0.354861
R143 VP.n130 VP.n129 0.354861
R144 VP VP.n130 0.267071
R145 VP.n35 VP.n34 0.189894
R146 VP.n36 VP.n35 0.189894
R147 VP.n36 VP.n29 0.189894
R148 VP.n40 VP.n29 0.189894
R149 VP.n41 VP.n40 0.189894
R150 VP.n42 VP.n41 0.189894
R151 VP.n42 VP.n27 0.189894
R152 VP.n47 VP.n27 0.189894
R153 VP.n48 VP.n47 0.189894
R154 VP.n49 VP.n48 0.189894
R155 VP.n49 VP.n25 0.189894
R156 VP.n53 VP.n25 0.189894
R157 VP.n54 VP.n53 0.189894
R158 VP.n55 VP.n54 0.189894
R159 VP.n55 VP.n23 0.189894
R160 VP.n60 VP.n23 0.189894
R161 VP.n61 VP.n60 0.189894
R162 VP.n62 VP.n61 0.189894
R163 VP.n62 VP.n21 0.189894
R164 VP.n66 VP.n21 0.189894
R165 VP.n67 VP.n66 0.189894
R166 VP.n68 VP.n67 0.189894
R167 VP.n68 VP.n19 0.189894
R168 VP.n72 VP.n19 0.189894
R169 VP.n78 VP.n17 0.189894
R170 VP.n79 VP.n78 0.189894
R171 VP.n80 VP.n79 0.189894
R172 VP.n80 VP.n15 0.189894
R173 VP.n84 VP.n15 0.189894
R174 VP.n85 VP.n84 0.189894
R175 VP.n86 VP.n85 0.189894
R176 VP.n86 VP.n13 0.189894
R177 VP.n91 VP.n13 0.189894
R178 VP.n92 VP.n91 0.189894
R179 VP.n93 VP.n92 0.189894
R180 VP.n93 VP.n11 0.189894
R181 VP.n97 VP.n11 0.189894
R182 VP.n98 VP.n97 0.189894
R183 VP.n99 VP.n98 0.189894
R184 VP.n99 VP.n9 0.189894
R185 VP.n104 VP.n9 0.189894
R186 VP.n105 VP.n104 0.189894
R187 VP.n106 VP.n105 0.189894
R188 VP.n106 VP.n7 0.189894
R189 VP.n110 VP.n7 0.189894
R190 VP.n111 VP.n110 0.189894
R191 VP.n112 VP.n111 0.189894
R192 VP.n112 VP.n5 0.189894
R193 VP.n117 VP.n5 0.189894
R194 VP.n118 VP.n117 0.189894
R195 VP.n119 VP.n118 0.189894
R196 VP.n119 VP.n3 0.189894
R197 VP.n123 VP.n3 0.189894
R198 VP.n124 VP.n123 0.189894
R199 VP.n125 VP.n124 0.189894
R200 VP.n125 VP.n1 0.189894
R201 VP.n129 VP.n1 0.189894
R202 VTAIL.n11 VTAIL.t6 52.1036
R203 VTAIL.n17 VTAIL.t3 52.1035
R204 VTAIL.n2 VTAIL.t10 52.1035
R205 VTAIL.n16 VTAIL.t15 52.1035
R206 VTAIL.n15 VTAIL.n14 50.1961
R207 VTAIL.n13 VTAIL.n12 50.1961
R208 VTAIL.n10 VTAIL.n9 50.1961
R209 VTAIL.n8 VTAIL.n7 50.1961
R210 VTAIL.n19 VTAIL.n18 50.1959
R211 VTAIL.n1 VTAIL.n0 50.1959
R212 VTAIL.n4 VTAIL.n3 50.1959
R213 VTAIL.n6 VTAIL.n5 50.1959
R214 VTAIL.n8 VTAIL.n6 34.2289
R215 VTAIL.n17 VTAIL.n16 30.6427
R216 VTAIL.n10 VTAIL.n8 3.58671
R217 VTAIL.n11 VTAIL.n10 3.58671
R218 VTAIL.n15 VTAIL.n13 3.58671
R219 VTAIL.n16 VTAIL.n15 3.58671
R220 VTAIL.n6 VTAIL.n4 3.58671
R221 VTAIL.n4 VTAIL.n2 3.58671
R222 VTAIL.n19 VTAIL.n17 3.58671
R223 VTAIL VTAIL.n1 2.74834
R224 VTAIL.n13 VTAIL.n11 2.26343
R225 VTAIL.n2 VTAIL.n1 2.26343
R226 VTAIL.n18 VTAIL.t4 1.90807
R227 VTAIL.n18 VTAIL.t0 1.90807
R228 VTAIL.n0 VTAIL.t8 1.90807
R229 VTAIL.n0 VTAIL.t5 1.90807
R230 VTAIL.n3 VTAIL.t17 1.90807
R231 VTAIL.n3 VTAIL.t18 1.90807
R232 VTAIL.n5 VTAIL.t9 1.90807
R233 VTAIL.n5 VTAIL.t12 1.90807
R234 VTAIL.n14 VTAIL.t14 1.90807
R235 VTAIL.n14 VTAIL.t16 1.90807
R236 VTAIL.n12 VTAIL.t11 1.90807
R237 VTAIL.n12 VTAIL.t13 1.90807
R238 VTAIL.n9 VTAIL.t1 1.90807
R239 VTAIL.n9 VTAIL.t19 1.90807
R240 VTAIL.n7 VTAIL.t7 1.90807
R241 VTAIL.n7 VTAIL.t2 1.90807
R242 VTAIL VTAIL.n19 0.838862
R243 VDD1.n1 VDD1.t9 72.3686
R244 VDD1.n3 VDD1.t0 72.3685
R245 VDD1.n5 VDD1.n4 69.509
R246 VDD1.n1 VDD1.n0 66.8749
R247 VDD1.n7 VDD1.n6 66.8747
R248 VDD1.n3 VDD1.n2 66.8747
R249 VDD1.n7 VDD1.n5 57.8155
R250 VDD1 VDD1.n7 2.63197
R251 VDD1.n6 VDD1.t5 1.90807
R252 VDD1.n6 VDD1.t6 1.90807
R253 VDD1.n0 VDD1.t7 1.90807
R254 VDD1.n0 VDD1.t8 1.90807
R255 VDD1.n4 VDD1.t3 1.90807
R256 VDD1.n4 VDD1.t2 1.90807
R257 VDD1.n2 VDD1.t4 1.90807
R258 VDD1.n2 VDD1.t1 1.90807
R259 VDD1 VDD1.n1 0.955241
R260 VDD1.n5 VDD1.n3 0.841706
R261 VN.n110 VN.n109 161.3
R262 VN.n108 VN.n57 161.3
R263 VN.n107 VN.n106 161.3
R264 VN.n105 VN.n58 161.3
R265 VN.n104 VN.n103 161.3
R266 VN.n102 VN.n59 161.3
R267 VN.n101 VN.n100 161.3
R268 VN.n99 VN.n60 161.3
R269 VN.n98 VN.n97 161.3
R270 VN.n95 VN.n61 161.3
R271 VN.n94 VN.n93 161.3
R272 VN.n92 VN.n62 161.3
R273 VN.n91 VN.n90 161.3
R274 VN.n89 VN.n63 161.3
R275 VN.n88 VN.n87 161.3
R276 VN.n86 VN.n64 161.3
R277 VN.n85 VN.n84 161.3
R278 VN.n82 VN.n65 161.3
R279 VN.n81 VN.n80 161.3
R280 VN.n79 VN.n66 161.3
R281 VN.n78 VN.n77 161.3
R282 VN.n76 VN.n67 161.3
R283 VN.n75 VN.n74 161.3
R284 VN.n73 VN.n68 161.3
R285 VN.n72 VN.n71 161.3
R286 VN.n54 VN.n53 161.3
R287 VN.n52 VN.n1 161.3
R288 VN.n51 VN.n50 161.3
R289 VN.n49 VN.n2 161.3
R290 VN.n48 VN.n47 161.3
R291 VN.n46 VN.n3 161.3
R292 VN.n45 VN.n44 161.3
R293 VN.n43 VN.n4 161.3
R294 VN.n42 VN.n41 161.3
R295 VN.n39 VN.n5 161.3
R296 VN.n38 VN.n37 161.3
R297 VN.n36 VN.n6 161.3
R298 VN.n35 VN.n34 161.3
R299 VN.n33 VN.n7 161.3
R300 VN.n32 VN.n31 161.3
R301 VN.n30 VN.n8 161.3
R302 VN.n29 VN.n28 161.3
R303 VN.n26 VN.n9 161.3
R304 VN.n25 VN.n24 161.3
R305 VN.n23 VN.n10 161.3
R306 VN.n22 VN.n21 161.3
R307 VN.n20 VN.n11 161.3
R308 VN.n19 VN.n18 161.3
R309 VN.n17 VN.n12 161.3
R310 VN.n16 VN.n15 161.3
R311 VN.n69 VN.t5 140.311
R312 VN.n13 VN.t3 140.311
R313 VN.n14 VN.t1 107.224
R314 VN.n27 VN.t7 107.224
R315 VN.n40 VN.t9 107.224
R316 VN.n0 VN.t8 107.224
R317 VN.n70 VN.t6 107.224
R318 VN.n83 VN.t4 107.224
R319 VN.n96 VN.t2 107.224
R320 VN.n56 VN.t0 107.224
R321 VN.n55 VN.n0 86.8027
R322 VN.n111 VN.n56 86.8027
R323 VN VN.n111 63.8542
R324 VN.n21 VN.n20 56.5617
R325 VN.n34 VN.n33 56.5617
R326 VN.n77 VN.n76 56.5617
R327 VN.n90 VN.n89 56.5617
R328 VN.n14 VN.n13 55.106
R329 VN.n70 VN.n69 55.106
R330 VN.n47 VN.n46 41.5458
R331 VN.n103 VN.n102 41.5458
R332 VN.n47 VN.n2 39.6083
R333 VN.n103 VN.n58 39.6083
R334 VN.n15 VN.n12 24.5923
R335 VN.n19 VN.n12 24.5923
R336 VN.n20 VN.n19 24.5923
R337 VN.n21 VN.n10 24.5923
R338 VN.n25 VN.n10 24.5923
R339 VN.n26 VN.n25 24.5923
R340 VN.n28 VN.n8 24.5923
R341 VN.n32 VN.n8 24.5923
R342 VN.n33 VN.n32 24.5923
R343 VN.n34 VN.n6 24.5923
R344 VN.n38 VN.n6 24.5923
R345 VN.n39 VN.n38 24.5923
R346 VN.n41 VN.n4 24.5923
R347 VN.n45 VN.n4 24.5923
R348 VN.n46 VN.n45 24.5923
R349 VN.n51 VN.n2 24.5923
R350 VN.n52 VN.n51 24.5923
R351 VN.n53 VN.n52 24.5923
R352 VN.n76 VN.n75 24.5923
R353 VN.n75 VN.n68 24.5923
R354 VN.n71 VN.n68 24.5923
R355 VN.n89 VN.n88 24.5923
R356 VN.n88 VN.n64 24.5923
R357 VN.n84 VN.n64 24.5923
R358 VN.n82 VN.n81 24.5923
R359 VN.n81 VN.n66 24.5923
R360 VN.n77 VN.n66 24.5923
R361 VN.n102 VN.n101 24.5923
R362 VN.n101 VN.n60 24.5923
R363 VN.n97 VN.n60 24.5923
R364 VN.n95 VN.n94 24.5923
R365 VN.n94 VN.n62 24.5923
R366 VN.n90 VN.n62 24.5923
R367 VN.n109 VN.n108 24.5923
R368 VN.n108 VN.n107 24.5923
R369 VN.n107 VN.n58 24.5923
R370 VN.n15 VN.n14 20.1658
R371 VN.n40 VN.n39 20.1658
R372 VN.n71 VN.n70 20.1658
R373 VN.n96 VN.n95 20.1658
R374 VN.n27 VN.n26 12.2964
R375 VN.n28 VN.n27 12.2964
R376 VN.n84 VN.n83 12.2964
R377 VN.n83 VN.n82 12.2964
R378 VN.n41 VN.n40 4.42703
R379 VN.n97 VN.n96 4.42703
R380 VN.n53 VN.n0 3.44336
R381 VN.n109 VN.n56 3.44336
R382 VN.n16 VN.n13 2.44069
R383 VN.n72 VN.n69 2.44069
R384 VN.n111 VN.n110 0.354861
R385 VN.n55 VN.n54 0.354861
R386 VN VN.n55 0.267071
R387 VN.n110 VN.n57 0.189894
R388 VN.n106 VN.n57 0.189894
R389 VN.n106 VN.n105 0.189894
R390 VN.n105 VN.n104 0.189894
R391 VN.n104 VN.n59 0.189894
R392 VN.n100 VN.n59 0.189894
R393 VN.n100 VN.n99 0.189894
R394 VN.n99 VN.n98 0.189894
R395 VN.n98 VN.n61 0.189894
R396 VN.n93 VN.n61 0.189894
R397 VN.n93 VN.n92 0.189894
R398 VN.n92 VN.n91 0.189894
R399 VN.n91 VN.n63 0.189894
R400 VN.n87 VN.n63 0.189894
R401 VN.n87 VN.n86 0.189894
R402 VN.n86 VN.n85 0.189894
R403 VN.n85 VN.n65 0.189894
R404 VN.n80 VN.n65 0.189894
R405 VN.n80 VN.n79 0.189894
R406 VN.n79 VN.n78 0.189894
R407 VN.n78 VN.n67 0.189894
R408 VN.n74 VN.n67 0.189894
R409 VN.n74 VN.n73 0.189894
R410 VN.n73 VN.n72 0.189894
R411 VN.n17 VN.n16 0.189894
R412 VN.n18 VN.n17 0.189894
R413 VN.n18 VN.n11 0.189894
R414 VN.n22 VN.n11 0.189894
R415 VN.n23 VN.n22 0.189894
R416 VN.n24 VN.n23 0.189894
R417 VN.n24 VN.n9 0.189894
R418 VN.n29 VN.n9 0.189894
R419 VN.n30 VN.n29 0.189894
R420 VN.n31 VN.n30 0.189894
R421 VN.n31 VN.n7 0.189894
R422 VN.n35 VN.n7 0.189894
R423 VN.n36 VN.n35 0.189894
R424 VN.n37 VN.n36 0.189894
R425 VN.n37 VN.n5 0.189894
R426 VN.n42 VN.n5 0.189894
R427 VN.n43 VN.n42 0.189894
R428 VN.n44 VN.n43 0.189894
R429 VN.n44 VN.n3 0.189894
R430 VN.n48 VN.n3 0.189894
R431 VN.n49 VN.n48 0.189894
R432 VN.n50 VN.n49 0.189894
R433 VN.n50 VN.n1 0.189894
R434 VN.n54 VN.n1 0.189894
R435 VDD2.n1 VDD2.t6 72.3685
R436 VDD2.n3 VDD2.n2 69.509
R437 VDD2 VDD2.n7 69.5062
R438 VDD2.n4 VDD2.t9 68.7824
R439 VDD2.n6 VDD2.n5 66.8749
R440 VDD2.n1 VDD2.n0 66.8747
R441 VDD2.n4 VDD2.n3 55.4394
R442 VDD2.n6 VDD2.n4 3.58671
R443 VDD2.n7 VDD2.t3 1.90807
R444 VDD2.n7 VDD2.t4 1.90807
R445 VDD2.n5 VDD2.t7 1.90807
R446 VDD2.n5 VDD2.t5 1.90807
R447 VDD2.n2 VDD2.t0 1.90807
R448 VDD2.n2 VDD2.t1 1.90807
R449 VDD2.n0 VDD2.t8 1.90807
R450 VDD2.n0 VDD2.t2 1.90807
R451 VDD2 VDD2.n6 0.955241
R452 VDD2.n3 VDD2.n1 0.841706
R453 B.n600 B.n599 585
R454 B.n598 B.n191 585
R455 B.n597 B.n596 585
R456 B.n595 B.n192 585
R457 B.n594 B.n593 585
R458 B.n592 B.n193 585
R459 B.n591 B.n590 585
R460 B.n589 B.n194 585
R461 B.n588 B.n587 585
R462 B.n586 B.n195 585
R463 B.n585 B.n584 585
R464 B.n583 B.n196 585
R465 B.n582 B.n581 585
R466 B.n580 B.n197 585
R467 B.n579 B.n578 585
R468 B.n577 B.n198 585
R469 B.n576 B.n575 585
R470 B.n574 B.n199 585
R471 B.n573 B.n572 585
R472 B.n571 B.n200 585
R473 B.n570 B.n569 585
R474 B.n568 B.n201 585
R475 B.n567 B.n566 585
R476 B.n565 B.n202 585
R477 B.n564 B.n563 585
R478 B.n562 B.n203 585
R479 B.n561 B.n560 585
R480 B.n559 B.n204 585
R481 B.n558 B.n557 585
R482 B.n556 B.n205 585
R483 B.n555 B.n554 585
R484 B.n553 B.n206 585
R485 B.n552 B.n551 585
R486 B.n550 B.n207 585
R487 B.n549 B.n548 585
R488 B.n547 B.n208 585
R489 B.n546 B.n545 585
R490 B.n544 B.n209 585
R491 B.n543 B.n542 585
R492 B.n541 B.n210 585
R493 B.n540 B.n539 585
R494 B.n538 B.n211 585
R495 B.n537 B.n536 585
R496 B.n535 B.n212 585
R497 B.n534 B.n533 585
R498 B.n532 B.n213 585
R499 B.n531 B.n530 585
R500 B.n529 B.n214 585
R501 B.n528 B.n527 585
R502 B.n526 B.n215 585
R503 B.n525 B.n524 585
R504 B.n523 B.n216 585
R505 B.n522 B.n521 585
R506 B.n520 B.n217 585
R507 B.n519 B.n518 585
R508 B.n517 B.n218 585
R509 B.n515 B.n514 585
R510 B.n513 B.n221 585
R511 B.n512 B.n511 585
R512 B.n510 B.n222 585
R513 B.n509 B.n508 585
R514 B.n507 B.n223 585
R515 B.n506 B.n505 585
R516 B.n504 B.n224 585
R517 B.n503 B.n502 585
R518 B.n501 B.n225 585
R519 B.n500 B.n499 585
R520 B.n495 B.n226 585
R521 B.n494 B.n493 585
R522 B.n492 B.n227 585
R523 B.n491 B.n490 585
R524 B.n489 B.n228 585
R525 B.n488 B.n487 585
R526 B.n486 B.n229 585
R527 B.n485 B.n484 585
R528 B.n483 B.n230 585
R529 B.n482 B.n481 585
R530 B.n480 B.n231 585
R531 B.n479 B.n478 585
R532 B.n477 B.n232 585
R533 B.n476 B.n475 585
R534 B.n474 B.n233 585
R535 B.n473 B.n472 585
R536 B.n471 B.n234 585
R537 B.n470 B.n469 585
R538 B.n468 B.n235 585
R539 B.n467 B.n466 585
R540 B.n465 B.n236 585
R541 B.n464 B.n463 585
R542 B.n462 B.n237 585
R543 B.n461 B.n460 585
R544 B.n459 B.n238 585
R545 B.n458 B.n457 585
R546 B.n456 B.n239 585
R547 B.n455 B.n454 585
R548 B.n453 B.n240 585
R549 B.n452 B.n451 585
R550 B.n450 B.n241 585
R551 B.n449 B.n448 585
R552 B.n447 B.n242 585
R553 B.n446 B.n445 585
R554 B.n444 B.n243 585
R555 B.n443 B.n442 585
R556 B.n441 B.n244 585
R557 B.n440 B.n439 585
R558 B.n438 B.n245 585
R559 B.n437 B.n436 585
R560 B.n435 B.n246 585
R561 B.n434 B.n433 585
R562 B.n432 B.n247 585
R563 B.n431 B.n430 585
R564 B.n429 B.n248 585
R565 B.n428 B.n427 585
R566 B.n426 B.n249 585
R567 B.n425 B.n424 585
R568 B.n423 B.n250 585
R569 B.n422 B.n421 585
R570 B.n420 B.n251 585
R571 B.n419 B.n418 585
R572 B.n417 B.n252 585
R573 B.n416 B.n415 585
R574 B.n414 B.n253 585
R575 B.n601 B.n190 585
R576 B.n603 B.n602 585
R577 B.n604 B.n189 585
R578 B.n606 B.n605 585
R579 B.n607 B.n188 585
R580 B.n609 B.n608 585
R581 B.n610 B.n187 585
R582 B.n612 B.n611 585
R583 B.n613 B.n186 585
R584 B.n615 B.n614 585
R585 B.n616 B.n185 585
R586 B.n618 B.n617 585
R587 B.n619 B.n184 585
R588 B.n621 B.n620 585
R589 B.n622 B.n183 585
R590 B.n624 B.n623 585
R591 B.n625 B.n182 585
R592 B.n627 B.n626 585
R593 B.n628 B.n181 585
R594 B.n630 B.n629 585
R595 B.n631 B.n180 585
R596 B.n633 B.n632 585
R597 B.n634 B.n179 585
R598 B.n636 B.n635 585
R599 B.n637 B.n178 585
R600 B.n639 B.n638 585
R601 B.n640 B.n177 585
R602 B.n642 B.n641 585
R603 B.n643 B.n176 585
R604 B.n645 B.n644 585
R605 B.n646 B.n175 585
R606 B.n648 B.n647 585
R607 B.n649 B.n174 585
R608 B.n651 B.n650 585
R609 B.n652 B.n173 585
R610 B.n654 B.n653 585
R611 B.n655 B.n172 585
R612 B.n657 B.n656 585
R613 B.n658 B.n171 585
R614 B.n660 B.n659 585
R615 B.n661 B.n170 585
R616 B.n663 B.n662 585
R617 B.n664 B.n169 585
R618 B.n666 B.n665 585
R619 B.n667 B.n168 585
R620 B.n669 B.n668 585
R621 B.n670 B.n167 585
R622 B.n672 B.n671 585
R623 B.n673 B.n166 585
R624 B.n675 B.n674 585
R625 B.n676 B.n165 585
R626 B.n678 B.n677 585
R627 B.n679 B.n164 585
R628 B.n681 B.n680 585
R629 B.n682 B.n163 585
R630 B.n684 B.n683 585
R631 B.n685 B.n162 585
R632 B.n687 B.n686 585
R633 B.n688 B.n161 585
R634 B.n690 B.n689 585
R635 B.n691 B.n160 585
R636 B.n693 B.n692 585
R637 B.n694 B.n159 585
R638 B.n696 B.n695 585
R639 B.n697 B.n158 585
R640 B.n699 B.n698 585
R641 B.n700 B.n157 585
R642 B.n702 B.n701 585
R643 B.n703 B.n156 585
R644 B.n705 B.n704 585
R645 B.n706 B.n155 585
R646 B.n708 B.n707 585
R647 B.n709 B.n154 585
R648 B.n711 B.n710 585
R649 B.n712 B.n153 585
R650 B.n714 B.n713 585
R651 B.n715 B.n152 585
R652 B.n717 B.n716 585
R653 B.n718 B.n151 585
R654 B.n720 B.n719 585
R655 B.n721 B.n150 585
R656 B.n723 B.n722 585
R657 B.n724 B.n149 585
R658 B.n726 B.n725 585
R659 B.n727 B.n148 585
R660 B.n729 B.n728 585
R661 B.n730 B.n147 585
R662 B.n732 B.n731 585
R663 B.n733 B.n146 585
R664 B.n735 B.n734 585
R665 B.n736 B.n145 585
R666 B.n738 B.n737 585
R667 B.n739 B.n144 585
R668 B.n741 B.n740 585
R669 B.n742 B.n143 585
R670 B.n744 B.n743 585
R671 B.n745 B.n142 585
R672 B.n747 B.n746 585
R673 B.n748 B.n141 585
R674 B.n750 B.n749 585
R675 B.n751 B.n140 585
R676 B.n753 B.n752 585
R677 B.n754 B.n139 585
R678 B.n756 B.n755 585
R679 B.n757 B.n138 585
R680 B.n759 B.n758 585
R681 B.n760 B.n137 585
R682 B.n762 B.n761 585
R683 B.n763 B.n136 585
R684 B.n765 B.n764 585
R685 B.n766 B.n135 585
R686 B.n768 B.n767 585
R687 B.n769 B.n134 585
R688 B.n771 B.n770 585
R689 B.n772 B.n133 585
R690 B.n774 B.n773 585
R691 B.n775 B.n132 585
R692 B.n777 B.n776 585
R693 B.n778 B.n131 585
R694 B.n780 B.n779 585
R695 B.n781 B.n130 585
R696 B.n783 B.n782 585
R697 B.n784 B.n129 585
R698 B.n786 B.n785 585
R699 B.n787 B.n128 585
R700 B.n789 B.n788 585
R701 B.n790 B.n127 585
R702 B.n792 B.n791 585
R703 B.n793 B.n126 585
R704 B.n795 B.n794 585
R705 B.n796 B.n125 585
R706 B.n798 B.n797 585
R707 B.n799 B.n124 585
R708 B.n801 B.n800 585
R709 B.n802 B.n123 585
R710 B.n804 B.n803 585
R711 B.n805 B.n122 585
R712 B.n807 B.n806 585
R713 B.n808 B.n121 585
R714 B.n810 B.n809 585
R715 B.n811 B.n120 585
R716 B.n813 B.n812 585
R717 B.n814 B.n119 585
R718 B.n816 B.n815 585
R719 B.n817 B.n118 585
R720 B.n819 B.n818 585
R721 B.n820 B.n117 585
R722 B.n822 B.n821 585
R723 B.n823 B.n116 585
R724 B.n825 B.n824 585
R725 B.n826 B.n115 585
R726 B.n828 B.n827 585
R727 B.n829 B.n114 585
R728 B.n831 B.n830 585
R729 B.n832 B.n113 585
R730 B.n834 B.n833 585
R731 B.n835 B.n112 585
R732 B.n837 B.n836 585
R733 B.n838 B.n111 585
R734 B.n840 B.n839 585
R735 B.n841 B.n110 585
R736 B.n843 B.n842 585
R737 B.n844 B.n109 585
R738 B.n846 B.n845 585
R739 B.n1030 B.n1029 585
R740 B.n1028 B.n43 585
R741 B.n1027 B.n1026 585
R742 B.n1025 B.n44 585
R743 B.n1024 B.n1023 585
R744 B.n1022 B.n45 585
R745 B.n1021 B.n1020 585
R746 B.n1019 B.n46 585
R747 B.n1018 B.n1017 585
R748 B.n1016 B.n47 585
R749 B.n1015 B.n1014 585
R750 B.n1013 B.n48 585
R751 B.n1012 B.n1011 585
R752 B.n1010 B.n49 585
R753 B.n1009 B.n1008 585
R754 B.n1007 B.n50 585
R755 B.n1006 B.n1005 585
R756 B.n1004 B.n51 585
R757 B.n1003 B.n1002 585
R758 B.n1001 B.n52 585
R759 B.n1000 B.n999 585
R760 B.n998 B.n53 585
R761 B.n997 B.n996 585
R762 B.n995 B.n54 585
R763 B.n994 B.n993 585
R764 B.n992 B.n55 585
R765 B.n991 B.n990 585
R766 B.n989 B.n56 585
R767 B.n988 B.n987 585
R768 B.n986 B.n57 585
R769 B.n985 B.n984 585
R770 B.n983 B.n58 585
R771 B.n982 B.n981 585
R772 B.n980 B.n59 585
R773 B.n979 B.n978 585
R774 B.n977 B.n60 585
R775 B.n976 B.n975 585
R776 B.n974 B.n61 585
R777 B.n973 B.n972 585
R778 B.n971 B.n62 585
R779 B.n970 B.n969 585
R780 B.n968 B.n63 585
R781 B.n967 B.n966 585
R782 B.n965 B.n64 585
R783 B.n964 B.n963 585
R784 B.n962 B.n65 585
R785 B.n961 B.n960 585
R786 B.n959 B.n66 585
R787 B.n958 B.n957 585
R788 B.n956 B.n67 585
R789 B.n955 B.n954 585
R790 B.n953 B.n68 585
R791 B.n952 B.n951 585
R792 B.n950 B.n69 585
R793 B.n949 B.n948 585
R794 B.n947 B.n70 585
R795 B.n946 B.n945 585
R796 B.n944 B.n71 585
R797 B.n943 B.n942 585
R798 B.n941 B.n75 585
R799 B.n940 B.n939 585
R800 B.n938 B.n76 585
R801 B.n937 B.n936 585
R802 B.n935 B.n77 585
R803 B.n934 B.n933 585
R804 B.n932 B.n78 585
R805 B.n930 B.n929 585
R806 B.n928 B.n81 585
R807 B.n927 B.n926 585
R808 B.n925 B.n82 585
R809 B.n924 B.n923 585
R810 B.n922 B.n83 585
R811 B.n921 B.n920 585
R812 B.n919 B.n84 585
R813 B.n918 B.n917 585
R814 B.n916 B.n85 585
R815 B.n915 B.n914 585
R816 B.n913 B.n86 585
R817 B.n912 B.n911 585
R818 B.n910 B.n87 585
R819 B.n909 B.n908 585
R820 B.n907 B.n88 585
R821 B.n906 B.n905 585
R822 B.n904 B.n89 585
R823 B.n903 B.n902 585
R824 B.n901 B.n90 585
R825 B.n900 B.n899 585
R826 B.n898 B.n91 585
R827 B.n897 B.n896 585
R828 B.n895 B.n92 585
R829 B.n894 B.n893 585
R830 B.n892 B.n93 585
R831 B.n891 B.n890 585
R832 B.n889 B.n94 585
R833 B.n888 B.n887 585
R834 B.n886 B.n95 585
R835 B.n885 B.n884 585
R836 B.n883 B.n96 585
R837 B.n882 B.n881 585
R838 B.n880 B.n97 585
R839 B.n879 B.n878 585
R840 B.n877 B.n98 585
R841 B.n876 B.n875 585
R842 B.n874 B.n99 585
R843 B.n873 B.n872 585
R844 B.n871 B.n100 585
R845 B.n870 B.n869 585
R846 B.n868 B.n101 585
R847 B.n867 B.n866 585
R848 B.n865 B.n102 585
R849 B.n864 B.n863 585
R850 B.n862 B.n103 585
R851 B.n861 B.n860 585
R852 B.n859 B.n104 585
R853 B.n858 B.n857 585
R854 B.n856 B.n105 585
R855 B.n855 B.n854 585
R856 B.n853 B.n106 585
R857 B.n852 B.n851 585
R858 B.n850 B.n107 585
R859 B.n849 B.n848 585
R860 B.n847 B.n108 585
R861 B.n1031 B.n42 585
R862 B.n1033 B.n1032 585
R863 B.n1034 B.n41 585
R864 B.n1036 B.n1035 585
R865 B.n1037 B.n40 585
R866 B.n1039 B.n1038 585
R867 B.n1040 B.n39 585
R868 B.n1042 B.n1041 585
R869 B.n1043 B.n38 585
R870 B.n1045 B.n1044 585
R871 B.n1046 B.n37 585
R872 B.n1048 B.n1047 585
R873 B.n1049 B.n36 585
R874 B.n1051 B.n1050 585
R875 B.n1052 B.n35 585
R876 B.n1054 B.n1053 585
R877 B.n1055 B.n34 585
R878 B.n1057 B.n1056 585
R879 B.n1058 B.n33 585
R880 B.n1060 B.n1059 585
R881 B.n1061 B.n32 585
R882 B.n1063 B.n1062 585
R883 B.n1064 B.n31 585
R884 B.n1066 B.n1065 585
R885 B.n1067 B.n30 585
R886 B.n1069 B.n1068 585
R887 B.n1070 B.n29 585
R888 B.n1072 B.n1071 585
R889 B.n1073 B.n28 585
R890 B.n1075 B.n1074 585
R891 B.n1076 B.n27 585
R892 B.n1078 B.n1077 585
R893 B.n1079 B.n26 585
R894 B.n1081 B.n1080 585
R895 B.n1082 B.n25 585
R896 B.n1084 B.n1083 585
R897 B.n1085 B.n24 585
R898 B.n1087 B.n1086 585
R899 B.n1088 B.n23 585
R900 B.n1090 B.n1089 585
R901 B.n1091 B.n22 585
R902 B.n1093 B.n1092 585
R903 B.n1094 B.n21 585
R904 B.n1096 B.n1095 585
R905 B.n1097 B.n20 585
R906 B.n1099 B.n1098 585
R907 B.n1100 B.n19 585
R908 B.n1102 B.n1101 585
R909 B.n1103 B.n18 585
R910 B.n1105 B.n1104 585
R911 B.n1106 B.n17 585
R912 B.n1108 B.n1107 585
R913 B.n1109 B.n16 585
R914 B.n1111 B.n1110 585
R915 B.n1112 B.n15 585
R916 B.n1114 B.n1113 585
R917 B.n1115 B.n14 585
R918 B.n1117 B.n1116 585
R919 B.n1118 B.n13 585
R920 B.n1120 B.n1119 585
R921 B.n1121 B.n12 585
R922 B.n1123 B.n1122 585
R923 B.n1124 B.n11 585
R924 B.n1126 B.n1125 585
R925 B.n1127 B.n10 585
R926 B.n1129 B.n1128 585
R927 B.n1130 B.n9 585
R928 B.n1132 B.n1131 585
R929 B.n1133 B.n8 585
R930 B.n1135 B.n1134 585
R931 B.n1136 B.n7 585
R932 B.n1138 B.n1137 585
R933 B.n1139 B.n6 585
R934 B.n1141 B.n1140 585
R935 B.n1142 B.n5 585
R936 B.n1144 B.n1143 585
R937 B.n1145 B.n4 585
R938 B.n1147 B.n1146 585
R939 B.n1148 B.n3 585
R940 B.n1150 B.n1149 585
R941 B.n1151 B.n0 585
R942 B.n2 B.n1 585
R943 B.n294 B.n293 585
R944 B.n296 B.n295 585
R945 B.n297 B.n292 585
R946 B.n299 B.n298 585
R947 B.n300 B.n291 585
R948 B.n302 B.n301 585
R949 B.n303 B.n290 585
R950 B.n305 B.n304 585
R951 B.n306 B.n289 585
R952 B.n308 B.n307 585
R953 B.n309 B.n288 585
R954 B.n311 B.n310 585
R955 B.n312 B.n287 585
R956 B.n314 B.n313 585
R957 B.n315 B.n286 585
R958 B.n317 B.n316 585
R959 B.n318 B.n285 585
R960 B.n320 B.n319 585
R961 B.n321 B.n284 585
R962 B.n323 B.n322 585
R963 B.n324 B.n283 585
R964 B.n326 B.n325 585
R965 B.n327 B.n282 585
R966 B.n329 B.n328 585
R967 B.n330 B.n281 585
R968 B.n332 B.n331 585
R969 B.n333 B.n280 585
R970 B.n335 B.n334 585
R971 B.n336 B.n279 585
R972 B.n338 B.n337 585
R973 B.n339 B.n278 585
R974 B.n341 B.n340 585
R975 B.n342 B.n277 585
R976 B.n344 B.n343 585
R977 B.n345 B.n276 585
R978 B.n347 B.n346 585
R979 B.n348 B.n275 585
R980 B.n350 B.n349 585
R981 B.n351 B.n274 585
R982 B.n353 B.n352 585
R983 B.n354 B.n273 585
R984 B.n356 B.n355 585
R985 B.n357 B.n272 585
R986 B.n359 B.n358 585
R987 B.n360 B.n271 585
R988 B.n362 B.n361 585
R989 B.n363 B.n270 585
R990 B.n365 B.n364 585
R991 B.n366 B.n269 585
R992 B.n368 B.n367 585
R993 B.n369 B.n268 585
R994 B.n371 B.n370 585
R995 B.n372 B.n267 585
R996 B.n374 B.n373 585
R997 B.n375 B.n266 585
R998 B.n377 B.n376 585
R999 B.n378 B.n265 585
R1000 B.n380 B.n379 585
R1001 B.n381 B.n264 585
R1002 B.n383 B.n382 585
R1003 B.n384 B.n263 585
R1004 B.n386 B.n385 585
R1005 B.n387 B.n262 585
R1006 B.n389 B.n388 585
R1007 B.n390 B.n261 585
R1008 B.n392 B.n391 585
R1009 B.n393 B.n260 585
R1010 B.n395 B.n394 585
R1011 B.n396 B.n259 585
R1012 B.n398 B.n397 585
R1013 B.n399 B.n258 585
R1014 B.n401 B.n400 585
R1015 B.n402 B.n257 585
R1016 B.n404 B.n403 585
R1017 B.n405 B.n256 585
R1018 B.n407 B.n406 585
R1019 B.n408 B.n255 585
R1020 B.n410 B.n409 585
R1021 B.n411 B.n254 585
R1022 B.n413 B.n412 585
R1023 B.n414 B.n413 540.549
R1024 B.n599 B.n190 540.549
R1025 B.n845 B.n108 540.549
R1026 B.n1031 B.n1030 540.549
R1027 B.n496 B.t6 316.589
R1028 B.n219 B.t9 316.589
R1029 B.n79 B.t0 316.589
R1030 B.n72 B.t3 316.589
R1031 B.n1153 B.n1152 256.663
R1032 B.n1152 B.n1151 235.042
R1033 B.n1152 B.n2 235.042
R1034 B.n219 B.t10 187.76
R1035 B.n79 B.t2 187.76
R1036 B.n496 B.t7 187.738
R1037 B.n72 B.t5 187.738
R1038 B.n415 B.n414 163.367
R1039 B.n415 B.n252 163.367
R1040 B.n419 B.n252 163.367
R1041 B.n420 B.n419 163.367
R1042 B.n421 B.n420 163.367
R1043 B.n421 B.n250 163.367
R1044 B.n425 B.n250 163.367
R1045 B.n426 B.n425 163.367
R1046 B.n427 B.n426 163.367
R1047 B.n427 B.n248 163.367
R1048 B.n431 B.n248 163.367
R1049 B.n432 B.n431 163.367
R1050 B.n433 B.n432 163.367
R1051 B.n433 B.n246 163.367
R1052 B.n437 B.n246 163.367
R1053 B.n438 B.n437 163.367
R1054 B.n439 B.n438 163.367
R1055 B.n439 B.n244 163.367
R1056 B.n443 B.n244 163.367
R1057 B.n444 B.n443 163.367
R1058 B.n445 B.n444 163.367
R1059 B.n445 B.n242 163.367
R1060 B.n449 B.n242 163.367
R1061 B.n450 B.n449 163.367
R1062 B.n451 B.n450 163.367
R1063 B.n451 B.n240 163.367
R1064 B.n455 B.n240 163.367
R1065 B.n456 B.n455 163.367
R1066 B.n457 B.n456 163.367
R1067 B.n457 B.n238 163.367
R1068 B.n461 B.n238 163.367
R1069 B.n462 B.n461 163.367
R1070 B.n463 B.n462 163.367
R1071 B.n463 B.n236 163.367
R1072 B.n467 B.n236 163.367
R1073 B.n468 B.n467 163.367
R1074 B.n469 B.n468 163.367
R1075 B.n469 B.n234 163.367
R1076 B.n473 B.n234 163.367
R1077 B.n474 B.n473 163.367
R1078 B.n475 B.n474 163.367
R1079 B.n475 B.n232 163.367
R1080 B.n479 B.n232 163.367
R1081 B.n480 B.n479 163.367
R1082 B.n481 B.n480 163.367
R1083 B.n481 B.n230 163.367
R1084 B.n485 B.n230 163.367
R1085 B.n486 B.n485 163.367
R1086 B.n487 B.n486 163.367
R1087 B.n487 B.n228 163.367
R1088 B.n491 B.n228 163.367
R1089 B.n492 B.n491 163.367
R1090 B.n493 B.n492 163.367
R1091 B.n493 B.n226 163.367
R1092 B.n500 B.n226 163.367
R1093 B.n501 B.n500 163.367
R1094 B.n502 B.n501 163.367
R1095 B.n502 B.n224 163.367
R1096 B.n506 B.n224 163.367
R1097 B.n507 B.n506 163.367
R1098 B.n508 B.n507 163.367
R1099 B.n508 B.n222 163.367
R1100 B.n512 B.n222 163.367
R1101 B.n513 B.n512 163.367
R1102 B.n514 B.n513 163.367
R1103 B.n514 B.n218 163.367
R1104 B.n519 B.n218 163.367
R1105 B.n520 B.n519 163.367
R1106 B.n521 B.n520 163.367
R1107 B.n521 B.n216 163.367
R1108 B.n525 B.n216 163.367
R1109 B.n526 B.n525 163.367
R1110 B.n527 B.n526 163.367
R1111 B.n527 B.n214 163.367
R1112 B.n531 B.n214 163.367
R1113 B.n532 B.n531 163.367
R1114 B.n533 B.n532 163.367
R1115 B.n533 B.n212 163.367
R1116 B.n537 B.n212 163.367
R1117 B.n538 B.n537 163.367
R1118 B.n539 B.n538 163.367
R1119 B.n539 B.n210 163.367
R1120 B.n543 B.n210 163.367
R1121 B.n544 B.n543 163.367
R1122 B.n545 B.n544 163.367
R1123 B.n545 B.n208 163.367
R1124 B.n549 B.n208 163.367
R1125 B.n550 B.n549 163.367
R1126 B.n551 B.n550 163.367
R1127 B.n551 B.n206 163.367
R1128 B.n555 B.n206 163.367
R1129 B.n556 B.n555 163.367
R1130 B.n557 B.n556 163.367
R1131 B.n557 B.n204 163.367
R1132 B.n561 B.n204 163.367
R1133 B.n562 B.n561 163.367
R1134 B.n563 B.n562 163.367
R1135 B.n563 B.n202 163.367
R1136 B.n567 B.n202 163.367
R1137 B.n568 B.n567 163.367
R1138 B.n569 B.n568 163.367
R1139 B.n569 B.n200 163.367
R1140 B.n573 B.n200 163.367
R1141 B.n574 B.n573 163.367
R1142 B.n575 B.n574 163.367
R1143 B.n575 B.n198 163.367
R1144 B.n579 B.n198 163.367
R1145 B.n580 B.n579 163.367
R1146 B.n581 B.n580 163.367
R1147 B.n581 B.n196 163.367
R1148 B.n585 B.n196 163.367
R1149 B.n586 B.n585 163.367
R1150 B.n587 B.n586 163.367
R1151 B.n587 B.n194 163.367
R1152 B.n591 B.n194 163.367
R1153 B.n592 B.n591 163.367
R1154 B.n593 B.n592 163.367
R1155 B.n593 B.n192 163.367
R1156 B.n597 B.n192 163.367
R1157 B.n598 B.n597 163.367
R1158 B.n599 B.n598 163.367
R1159 B.n845 B.n844 163.367
R1160 B.n844 B.n843 163.367
R1161 B.n843 B.n110 163.367
R1162 B.n839 B.n110 163.367
R1163 B.n839 B.n838 163.367
R1164 B.n838 B.n837 163.367
R1165 B.n837 B.n112 163.367
R1166 B.n833 B.n112 163.367
R1167 B.n833 B.n832 163.367
R1168 B.n832 B.n831 163.367
R1169 B.n831 B.n114 163.367
R1170 B.n827 B.n114 163.367
R1171 B.n827 B.n826 163.367
R1172 B.n826 B.n825 163.367
R1173 B.n825 B.n116 163.367
R1174 B.n821 B.n116 163.367
R1175 B.n821 B.n820 163.367
R1176 B.n820 B.n819 163.367
R1177 B.n819 B.n118 163.367
R1178 B.n815 B.n118 163.367
R1179 B.n815 B.n814 163.367
R1180 B.n814 B.n813 163.367
R1181 B.n813 B.n120 163.367
R1182 B.n809 B.n120 163.367
R1183 B.n809 B.n808 163.367
R1184 B.n808 B.n807 163.367
R1185 B.n807 B.n122 163.367
R1186 B.n803 B.n122 163.367
R1187 B.n803 B.n802 163.367
R1188 B.n802 B.n801 163.367
R1189 B.n801 B.n124 163.367
R1190 B.n797 B.n124 163.367
R1191 B.n797 B.n796 163.367
R1192 B.n796 B.n795 163.367
R1193 B.n795 B.n126 163.367
R1194 B.n791 B.n126 163.367
R1195 B.n791 B.n790 163.367
R1196 B.n790 B.n789 163.367
R1197 B.n789 B.n128 163.367
R1198 B.n785 B.n128 163.367
R1199 B.n785 B.n784 163.367
R1200 B.n784 B.n783 163.367
R1201 B.n783 B.n130 163.367
R1202 B.n779 B.n130 163.367
R1203 B.n779 B.n778 163.367
R1204 B.n778 B.n777 163.367
R1205 B.n777 B.n132 163.367
R1206 B.n773 B.n132 163.367
R1207 B.n773 B.n772 163.367
R1208 B.n772 B.n771 163.367
R1209 B.n771 B.n134 163.367
R1210 B.n767 B.n134 163.367
R1211 B.n767 B.n766 163.367
R1212 B.n766 B.n765 163.367
R1213 B.n765 B.n136 163.367
R1214 B.n761 B.n136 163.367
R1215 B.n761 B.n760 163.367
R1216 B.n760 B.n759 163.367
R1217 B.n759 B.n138 163.367
R1218 B.n755 B.n138 163.367
R1219 B.n755 B.n754 163.367
R1220 B.n754 B.n753 163.367
R1221 B.n753 B.n140 163.367
R1222 B.n749 B.n140 163.367
R1223 B.n749 B.n748 163.367
R1224 B.n748 B.n747 163.367
R1225 B.n747 B.n142 163.367
R1226 B.n743 B.n142 163.367
R1227 B.n743 B.n742 163.367
R1228 B.n742 B.n741 163.367
R1229 B.n741 B.n144 163.367
R1230 B.n737 B.n144 163.367
R1231 B.n737 B.n736 163.367
R1232 B.n736 B.n735 163.367
R1233 B.n735 B.n146 163.367
R1234 B.n731 B.n146 163.367
R1235 B.n731 B.n730 163.367
R1236 B.n730 B.n729 163.367
R1237 B.n729 B.n148 163.367
R1238 B.n725 B.n148 163.367
R1239 B.n725 B.n724 163.367
R1240 B.n724 B.n723 163.367
R1241 B.n723 B.n150 163.367
R1242 B.n719 B.n150 163.367
R1243 B.n719 B.n718 163.367
R1244 B.n718 B.n717 163.367
R1245 B.n717 B.n152 163.367
R1246 B.n713 B.n152 163.367
R1247 B.n713 B.n712 163.367
R1248 B.n712 B.n711 163.367
R1249 B.n711 B.n154 163.367
R1250 B.n707 B.n154 163.367
R1251 B.n707 B.n706 163.367
R1252 B.n706 B.n705 163.367
R1253 B.n705 B.n156 163.367
R1254 B.n701 B.n156 163.367
R1255 B.n701 B.n700 163.367
R1256 B.n700 B.n699 163.367
R1257 B.n699 B.n158 163.367
R1258 B.n695 B.n158 163.367
R1259 B.n695 B.n694 163.367
R1260 B.n694 B.n693 163.367
R1261 B.n693 B.n160 163.367
R1262 B.n689 B.n160 163.367
R1263 B.n689 B.n688 163.367
R1264 B.n688 B.n687 163.367
R1265 B.n687 B.n162 163.367
R1266 B.n683 B.n162 163.367
R1267 B.n683 B.n682 163.367
R1268 B.n682 B.n681 163.367
R1269 B.n681 B.n164 163.367
R1270 B.n677 B.n164 163.367
R1271 B.n677 B.n676 163.367
R1272 B.n676 B.n675 163.367
R1273 B.n675 B.n166 163.367
R1274 B.n671 B.n166 163.367
R1275 B.n671 B.n670 163.367
R1276 B.n670 B.n669 163.367
R1277 B.n669 B.n168 163.367
R1278 B.n665 B.n168 163.367
R1279 B.n665 B.n664 163.367
R1280 B.n664 B.n663 163.367
R1281 B.n663 B.n170 163.367
R1282 B.n659 B.n170 163.367
R1283 B.n659 B.n658 163.367
R1284 B.n658 B.n657 163.367
R1285 B.n657 B.n172 163.367
R1286 B.n653 B.n172 163.367
R1287 B.n653 B.n652 163.367
R1288 B.n652 B.n651 163.367
R1289 B.n651 B.n174 163.367
R1290 B.n647 B.n174 163.367
R1291 B.n647 B.n646 163.367
R1292 B.n646 B.n645 163.367
R1293 B.n645 B.n176 163.367
R1294 B.n641 B.n176 163.367
R1295 B.n641 B.n640 163.367
R1296 B.n640 B.n639 163.367
R1297 B.n639 B.n178 163.367
R1298 B.n635 B.n178 163.367
R1299 B.n635 B.n634 163.367
R1300 B.n634 B.n633 163.367
R1301 B.n633 B.n180 163.367
R1302 B.n629 B.n180 163.367
R1303 B.n629 B.n628 163.367
R1304 B.n628 B.n627 163.367
R1305 B.n627 B.n182 163.367
R1306 B.n623 B.n182 163.367
R1307 B.n623 B.n622 163.367
R1308 B.n622 B.n621 163.367
R1309 B.n621 B.n184 163.367
R1310 B.n617 B.n184 163.367
R1311 B.n617 B.n616 163.367
R1312 B.n616 B.n615 163.367
R1313 B.n615 B.n186 163.367
R1314 B.n611 B.n186 163.367
R1315 B.n611 B.n610 163.367
R1316 B.n610 B.n609 163.367
R1317 B.n609 B.n188 163.367
R1318 B.n605 B.n188 163.367
R1319 B.n605 B.n604 163.367
R1320 B.n604 B.n603 163.367
R1321 B.n603 B.n190 163.367
R1322 B.n1030 B.n43 163.367
R1323 B.n1026 B.n43 163.367
R1324 B.n1026 B.n1025 163.367
R1325 B.n1025 B.n1024 163.367
R1326 B.n1024 B.n45 163.367
R1327 B.n1020 B.n45 163.367
R1328 B.n1020 B.n1019 163.367
R1329 B.n1019 B.n1018 163.367
R1330 B.n1018 B.n47 163.367
R1331 B.n1014 B.n47 163.367
R1332 B.n1014 B.n1013 163.367
R1333 B.n1013 B.n1012 163.367
R1334 B.n1012 B.n49 163.367
R1335 B.n1008 B.n49 163.367
R1336 B.n1008 B.n1007 163.367
R1337 B.n1007 B.n1006 163.367
R1338 B.n1006 B.n51 163.367
R1339 B.n1002 B.n51 163.367
R1340 B.n1002 B.n1001 163.367
R1341 B.n1001 B.n1000 163.367
R1342 B.n1000 B.n53 163.367
R1343 B.n996 B.n53 163.367
R1344 B.n996 B.n995 163.367
R1345 B.n995 B.n994 163.367
R1346 B.n994 B.n55 163.367
R1347 B.n990 B.n55 163.367
R1348 B.n990 B.n989 163.367
R1349 B.n989 B.n988 163.367
R1350 B.n988 B.n57 163.367
R1351 B.n984 B.n57 163.367
R1352 B.n984 B.n983 163.367
R1353 B.n983 B.n982 163.367
R1354 B.n982 B.n59 163.367
R1355 B.n978 B.n59 163.367
R1356 B.n978 B.n977 163.367
R1357 B.n977 B.n976 163.367
R1358 B.n976 B.n61 163.367
R1359 B.n972 B.n61 163.367
R1360 B.n972 B.n971 163.367
R1361 B.n971 B.n970 163.367
R1362 B.n970 B.n63 163.367
R1363 B.n966 B.n63 163.367
R1364 B.n966 B.n965 163.367
R1365 B.n965 B.n964 163.367
R1366 B.n964 B.n65 163.367
R1367 B.n960 B.n65 163.367
R1368 B.n960 B.n959 163.367
R1369 B.n959 B.n958 163.367
R1370 B.n958 B.n67 163.367
R1371 B.n954 B.n67 163.367
R1372 B.n954 B.n953 163.367
R1373 B.n953 B.n952 163.367
R1374 B.n952 B.n69 163.367
R1375 B.n948 B.n69 163.367
R1376 B.n948 B.n947 163.367
R1377 B.n947 B.n946 163.367
R1378 B.n946 B.n71 163.367
R1379 B.n942 B.n71 163.367
R1380 B.n942 B.n941 163.367
R1381 B.n941 B.n940 163.367
R1382 B.n940 B.n76 163.367
R1383 B.n936 B.n76 163.367
R1384 B.n936 B.n935 163.367
R1385 B.n935 B.n934 163.367
R1386 B.n934 B.n78 163.367
R1387 B.n929 B.n78 163.367
R1388 B.n929 B.n928 163.367
R1389 B.n928 B.n927 163.367
R1390 B.n927 B.n82 163.367
R1391 B.n923 B.n82 163.367
R1392 B.n923 B.n922 163.367
R1393 B.n922 B.n921 163.367
R1394 B.n921 B.n84 163.367
R1395 B.n917 B.n84 163.367
R1396 B.n917 B.n916 163.367
R1397 B.n916 B.n915 163.367
R1398 B.n915 B.n86 163.367
R1399 B.n911 B.n86 163.367
R1400 B.n911 B.n910 163.367
R1401 B.n910 B.n909 163.367
R1402 B.n909 B.n88 163.367
R1403 B.n905 B.n88 163.367
R1404 B.n905 B.n904 163.367
R1405 B.n904 B.n903 163.367
R1406 B.n903 B.n90 163.367
R1407 B.n899 B.n90 163.367
R1408 B.n899 B.n898 163.367
R1409 B.n898 B.n897 163.367
R1410 B.n897 B.n92 163.367
R1411 B.n893 B.n92 163.367
R1412 B.n893 B.n892 163.367
R1413 B.n892 B.n891 163.367
R1414 B.n891 B.n94 163.367
R1415 B.n887 B.n94 163.367
R1416 B.n887 B.n886 163.367
R1417 B.n886 B.n885 163.367
R1418 B.n885 B.n96 163.367
R1419 B.n881 B.n96 163.367
R1420 B.n881 B.n880 163.367
R1421 B.n880 B.n879 163.367
R1422 B.n879 B.n98 163.367
R1423 B.n875 B.n98 163.367
R1424 B.n875 B.n874 163.367
R1425 B.n874 B.n873 163.367
R1426 B.n873 B.n100 163.367
R1427 B.n869 B.n100 163.367
R1428 B.n869 B.n868 163.367
R1429 B.n868 B.n867 163.367
R1430 B.n867 B.n102 163.367
R1431 B.n863 B.n102 163.367
R1432 B.n863 B.n862 163.367
R1433 B.n862 B.n861 163.367
R1434 B.n861 B.n104 163.367
R1435 B.n857 B.n104 163.367
R1436 B.n857 B.n856 163.367
R1437 B.n856 B.n855 163.367
R1438 B.n855 B.n106 163.367
R1439 B.n851 B.n106 163.367
R1440 B.n851 B.n850 163.367
R1441 B.n850 B.n849 163.367
R1442 B.n849 B.n108 163.367
R1443 B.n1032 B.n1031 163.367
R1444 B.n1032 B.n41 163.367
R1445 B.n1036 B.n41 163.367
R1446 B.n1037 B.n1036 163.367
R1447 B.n1038 B.n1037 163.367
R1448 B.n1038 B.n39 163.367
R1449 B.n1042 B.n39 163.367
R1450 B.n1043 B.n1042 163.367
R1451 B.n1044 B.n1043 163.367
R1452 B.n1044 B.n37 163.367
R1453 B.n1048 B.n37 163.367
R1454 B.n1049 B.n1048 163.367
R1455 B.n1050 B.n1049 163.367
R1456 B.n1050 B.n35 163.367
R1457 B.n1054 B.n35 163.367
R1458 B.n1055 B.n1054 163.367
R1459 B.n1056 B.n1055 163.367
R1460 B.n1056 B.n33 163.367
R1461 B.n1060 B.n33 163.367
R1462 B.n1061 B.n1060 163.367
R1463 B.n1062 B.n1061 163.367
R1464 B.n1062 B.n31 163.367
R1465 B.n1066 B.n31 163.367
R1466 B.n1067 B.n1066 163.367
R1467 B.n1068 B.n1067 163.367
R1468 B.n1068 B.n29 163.367
R1469 B.n1072 B.n29 163.367
R1470 B.n1073 B.n1072 163.367
R1471 B.n1074 B.n1073 163.367
R1472 B.n1074 B.n27 163.367
R1473 B.n1078 B.n27 163.367
R1474 B.n1079 B.n1078 163.367
R1475 B.n1080 B.n1079 163.367
R1476 B.n1080 B.n25 163.367
R1477 B.n1084 B.n25 163.367
R1478 B.n1085 B.n1084 163.367
R1479 B.n1086 B.n1085 163.367
R1480 B.n1086 B.n23 163.367
R1481 B.n1090 B.n23 163.367
R1482 B.n1091 B.n1090 163.367
R1483 B.n1092 B.n1091 163.367
R1484 B.n1092 B.n21 163.367
R1485 B.n1096 B.n21 163.367
R1486 B.n1097 B.n1096 163.367
R1487 B.n1098 B.n1097 163.367
R1488 B.n1098 B.n19 163.367
R1489 B.n1102 B.n19 163.367
R1490 B.n1103 B.n1102 163.367
R1491 B.n1104 B.n1103 163.367
R1492 B.n1104 B.n17 163.367
R1493 B.n1108 B.n17 163.367
R1494 B.n1109 B.n1108 163.367
R1495 B.n1110 B.n1109 163.367
R1496 B.n1110 B.n15 163.367
R1497 B.n1114 B.n15 163.367
R1498 B.n1115 B.n1114 163.367
R1499 B.n1116 B.n1115 163.367
R1500 B.n1116 B.n13 163.367
R1501 B.n1120 B.n13 163.367
R1502 B.n1121 B.n1120 163.367
R1503 B.n1122 B.n1121 163.367
R1504 B.n1122 B.n11 163.367
R1505 B.n1126 B.n11 163.367
R1506 B.n1127 B.n1126 163.367
R1507 B.n1128 B.n1127 163.367
R1508 B.n1128 B.n9 163.367
R1509 B.n1132 B.n9 163.367
R1510 B.n1133 B.n1132 163.367
R1511 B.n1134 B.n1133 163.367
R1512 B.n1134 B.n7 163.367
R1513 B.n1138 B.n7 163.367
R1514 B.n1139 B.n1138 163.367
R1515 B.n1140 B.n1139 163.367
R1516 B.n1140 B.n5 163.367
R1517 B.n1144 B.n5 163.367
R1518 B.n1145 B.n1144 163.367
R1519 B.n1146 B.n1145 163.367
R1520 B.n1146 B.n3 163.367
R1521 B.n1150 B.n3 163.367
R1522 B.n1151 B.n1150 163.367
R1523 B.n294 B.n2 163.367
R1524 B.n295 B.n294 163.367
R1525 B.n295 B.n292 163.367
R1526 B.n299 B.n292 163.367
R1527 B.n300 B.n299 163.367
R1528 B.n301 B.n300 163.367
R1529 B.n301 B.n290 163.367
R1530 B.n305 B.n290 163.367
R1531 B.n306 B.n305 163.367
R1532 B.n307 B.n306 163.367
R1533 B.n307 B.n288 163.367
R1534 B.n311 B.n288 163.367
R1535 B.n312 B.n311 163.367
R1536 B.n313 B.n312 163.367
R1537 B.n313 B.n286 163.367
R1538 B.n317 B.n286 163.367
R1539 B.n318 B.n317 163.367
R1540 B.n319 B.n318 163.367
R1541 B.n319 B.n284 163.367
R1542 B.n323 B.n284 163.367
R1543 B.n324 B.n323 163.367
R1544 B.n325 B.n324 163.367
R1545 B.n325 B.n282 163.367
R1546 B.n329 B.n282 163.367
R1547 B.n330 B.n329 163.367
R1548 B.n331 B.n330 163.367
R1549 B.n331 B.n280 163.367
R1550 B.n335 B.n280 163.367
R1551 B.n336 B.n335 163.367
R1552 B.n337 B.n336 163.367
R1553 B.n337 B.n278 163.367
R1554 B.n341 B.n278 163.367
R1555 B.n342 B.n341 163.367
R1556 B.n343 B.n342 163.367
R1557 B.n343 B.n276 163.367
R1558 B.n347 B.n276 163.367
R1559 B.n348 B.n347 163.367
R1560 B.n349 B.n348 163.367
R1561 B.n349 B.n274 163.367
R1562 B.n353 B.n274 163.367
R1563 B.n354 B.n353 163.367
R1564 B.n355 B.n354 163.367
R1565 B.n355 B.n272 163.367
R1566 B.n359 B.n272 163.367
R1567 B.n360 B.n359 163.367
R1568 B.n361 B.n360 163.367
R1569 B.n361 B.n270 163.367
R1570 B.n365 B.n270 163.367
R1571 B.n366 B.n365 163.367
R1572 B.n367 B.n366 163.367
R1573 B.n367 B.n268 163.367
R1574 B.n371 B.n268 163.367
R1575 B.n372 B.n371 163.367
R1576 B.n373 B.n372 163.367
R1577 B.n373 B.n266 163.367
R1578 B.n377 B.n266 163.367
R1579 B.n378 B.n377 163.367
R1580 B.n379 B.n378 163.367
R1581 B.n379 B.n264 163.367
R1582 B.n383 B.n264 163.367
R1583 B.n384 B.n383 163.367
R1584 B.n385 B.n384 163.367
R1585 B.n385 B.n262 163.367
R1586 B.n389 B.n262 163.367
R1587 B.n390 B.n389 163.367
R1588 B.n391 B.n390 163.367
R1589 B.n391 B.n260 163.367
R1590 B.n395 B.n260 163.367
R1591 B.n396 B.n395 163.367
R1592 B.n397 B.n396 163.367
R1593 B.n397 B.n258 163.367
R1594 B.n401 B.n258 163.367
R1595 B.n402 B.n401 163.367
R1596 B.n403 B.n402 163.367
R1597 B.n403 B.n256 163.367
R1598 B.n407 B.n256 163.367
R1599 B.n408 B.n407 163.367
R1600 B.n409 B.n408 163.367
R1601 B.n409 B.n254 163.367
R1602 B.n413 B.n254 163.367
R1603 B.n220 B.t11 107.081
R1604 B.n80 B.t1 107.081
R1605 B.n497 B.t8 107.058
R1606 B.n73 B.t4 107.058
R1607 B.n497 B.n496 80.6793
R1608 B.n220 B.n219 80.6793
R1609 B.n80 B.n79 80.6793
R1610 B.n73 B.n72 80.6793
R1611 B.n498 B.n497 59.5399
R1612 B.n516 B.n220 59.5399
R1613 B.n931 B.n80 59.5399
R1614 B.n74 B.n73 59.5399
R1615 B.n1029 B.n42 35.1225
R1616 B.n847 B.n846 35.1225
R1617 B.n601 B.n600 35.1225
R1618 B.n412 B.n253 35.1225
R1619 B B.n1153 18.0485
R1620 B.n1033 B.n42 10.6151
R1621 B.n1034 B.n1033 10.6151
R1622 B.n1035 B.n1034 10.6151
R1623 B.n1035 B.n40 10.6151
R1624 B.n1039 B.n40 10.6151
R1625 B.n1040 B.n1039 10.6151
R1626 B.n1041 B.n1040 10.6151
R1627 B.n1041 B.n38 10.6151
R1628 B.n1045 B.n38 10.6151
R1629 B.n1046 B.n1045 10.6151
R1630 B.n1047 B.n1046 10.6151
R1631 B.n1047 B.n36 10.6151
R1632 B.n1051 B.n36 10.6151
R1633 B.n1052 B.n1051 10.6151
R1634 B.n1053 B.n1052 10.6151
R1635 B.n1053 B.n34 10.6151
R1636 B.n1057 B.n34 10.6151
R1637 B.n1058 B.n1057 10.6151
R1638 B.n1059 B.n1058 10.6151
R1639 B.n1059 B.n32 10.6151
R1640 B.n1063 B.n32 10.6151
R1641 B.n1064 B.n1063 10.6151
R1642 B.n1065 B.n1064 10.6151
R1643 B.n1065 B.n30 10.6151
R1644 B.n1069 B.n30 10.6151
R1645 B.n1070 B.n1069 10.6151
R1646 B.n1071 B.n1070 10.6151
R1647 B.n1071 B.n28 10.6151
R1648 B.n1075 B.n28 10.6151
R1649 B.n1076 B.n1075 10.6151
R1650 B.n1077 B.n1076 10.6151
R1651 B.n1077 B.n26 10.6151
R1652 B.n1081 B.n26 10.6151
R1653 B.n1082 B.n1081 10.6151
R1654 B.n1083 B.n1082 10.6151
R1655 B.n1083 B.n24 10.6151
R1656 B.n1087 B.n24 10.6151
R1657 B.n1088 B.n1087 10.6151
R1658 B.n1089 B.n1088 10.6151
R1659 B.n1089 B.n22 10.6151
R1660 B.n1093 B.n22 10.6151
R1661 B.n1094 B.n1093 10.6151
R1662 B.n1095 B.n1094 10.6151
R1663 B.n1095 B.n20 10.6151
R1664 B.n1099 B.n20 10.6151
R1665 B.n1100 B.n1099 10.6151
R1666 B.n1101 B.n1100 10.6151
R1667 B.n1101 B.n18 10.6151
R1668 B.n1105 B.n18 10.6151
R1669 B.n1106 B.n1105 10.6151
R1670 B.n1107 B.n1106 10.6151
R1671 B.n1107 B.n16 10.6151
R1672 B.n1111 B.n16 10.6151
R1673 B.n1112 B.n1111 10.6151
R1674 B.n1113 B.n1112 10.6151
R1675 B.n1113 B.n14 10.6151
R1676 B.n1117 B.n14 10.6151
R1677 B.n1118 B.n1117 10.6151
R1678 B.n1119 B.n1118 10.6151
R1679 B.n1119 B.n12 10.6151
R1680 B.n1123 B.n12 10.6151
R1681 B.n1124 B.n1123 10.6151
R1682 B.n1125 B.n1124 10.6151
R1683 B.n1125 B.n10 10.6151
R1684 B.n1129 B.n10 10.6151
R1685 B.n1130 B.n1129 10.6151
R1686 B.n1131 B.n1130 10.6151
R1687 B.n1131 B.n8 10.6151
R1688 B.n1135 B.n8 10.6151
R1689 B.n1136 B.n1135 10.6151
R1690 B.n1137 B.n1136 10.6151
R1691 B.n1137 B.n6 10.6151
R1692 B.n1141 B.n6 10.6151
R1693 B.n1142 B.n1141 10.6151
R1694 B.n1143 B.n1142 10.6151
R1695 B.n1143 B.n4 10.6151
R1696 B.n1147 B.n4 10.6151
R1697 B.n1148 B.n1147 10.6151
R1698 B.n1149 B.n1148 10.6151
R1699 B.n1149 B.n0 10.6151
R1700 B.n1029 B.n1028 10.6151
R1701 B.n1028 B.n1027 10.6151
R1702 B.n1027 B.n44 10.6151
R1703 B.n1023 B.n44 10.6151
R1704 B.n1023 B.n1022 10.6151
R1705 B.n1022 B.n1021 10.6151
R1706 B.n1021 B.n46 10.6151
R1707 B.n1017 B.n46 10.6151
R1708 B.n1017 B.n1016 10.6151
R1709 B.n1016 B.n1015 10.6151
R1710 B.n1015 B.n48 10.6151
R1711 B.n1011 B.n48 10.6151
R1712 B.n1011 B.n1010 10.6151
R1713 B.n1010 B.n1009 10.6151
R1714 B.n1009 B.n50 10.6151
R1715 B.n1005 B.n50 10.6151
R1716 B.n1005 B.n1004 10.6151
R1717 B.n1004 B.n1003 10.6151
R1718 B.n1003 B.n52 10.6151
R1719 B.n999 B.n52 10.6151
R1720 B.n999 B.n998 10.6151
R1721 B.n998 B.n997 10.6151
R1722 B.n997 B.n54 10.6151
R1723 B.n993 B.n54 10.6151
R1724 B.n993 B.n992 10.6151
R1725 B.n992 B.n991 10.6151
R1726 B.n991 B.n56 10.6151
R1727 B.n987 B.n56 10.6151
R1728 B.n987 B.n986 10.6151
R1729 B.n986 B.n985 10.6151
R1730 B.n985 B.n58 10.6151
R1731 B.n981 B.n58 10.6151
R1732 B.n981 B.n980 10.6151
R1733 B.n980 B.n979 10.6151
R1734 B.n979 B.n60 10.6151
R1735 B.n975 B.n60 10.6151
R1736 B.n975 B.n974 10.6151
R1737 B.n974 B.n973 10.6151
R1738 B.n973 B.n62 10.6151
R1739 B.n969 B.n62 10.6151
R1740 B.n969 B.n968 10.6151
R1741 B.n968 B.n967 10.6151
R1742 B.n967 B.n64 10.6151
R1743 B.n963 B.n64 10.6151
R1744 B.n963 B.n962 10.6151
R1745 B.n962 B.n961 10.6151
R1746 B.n961 B.n66 10.6151
R1747 B.n957 B.n66 10.6151
R1748 B.n957 B.n956 10.6151
R1749 B.n956 B.n955 10.6151
R1750 B.n955 B.n68 10.6151
R1751 B.n951 B.n68 10.6151
R1752 B.n951 B.n950 10.6151
R1753 B.n950 B.n949 10.6151
R1754 B.n949 B.n70 10.6151
R1755 B.n945 B.n944 10.6151
R1756 B.n944 B.n943 10.6151
R1757 B.n943 B.n75 10.6151
R1758 B.n939 B.n75 10.6151
R1759 B.n939 B.n938 10.6151
R1760 B.n938 B.n937 10.6151
R1761 B.n937 B.n77 10.6151
R1762 B.n933 B.n77 10.6151
R1763 B.n933 B.n932 10.6151
R1764 B.n930 B.n81 10.6151
R1765 B.n926 B.n81 10.6151
R1766 B.n926 B.n925 10.6151
R1767 B.n925 B.n924 10.6151
R1768 B.n924 B.n83 10.6151
R1769 B.n920 B.n83 10.6151
R1770 B.n920 B.n919 10.6151
R1771 B.n919 B.n918 10.6151
R1772 B.n918 B.n85 10.6151
R1773 B.n914 B.n85 10.6151
R1774 B.n914 B.n913 10.6151
R1775 B.n913 B.n912 10.6151
R1776 B.n912 B.n87 10.6151
R1777 B.n908 B.n87 10.6151
R1778 B.n908 B.n907 10.6151
R1779 B.n907 B.n906 10.6151
R1780 B.n906 B.n89 10.6151
R1781 B.n902 B.n89 10.6151
R1782 B.n902 B.n901 10.6151
R1783 B.n901 B.n900 10.6151
R1784 B.n900 B.n91 10.6151
R1785 B.n896 B.n91 10.6151
R1786 B.n896 B.n895 10.6151
R1787 B.n895 B.n894 10.6151
R1788 B.n894 B.n93 10.6151
R1789 B.n890 B.n93 10.6151
R1790 B.n890 B.n889 10.6151
R1791 B.n889 B.n888 10.6151
R1792 B.n888 B.n95 10.6151
R1793 B.n884 B.n95 10.6151
R1794 B.n884 B.n883 10.6151
R1795 B.n883 B.n882 10.6151
R1796 B.n882 B.n97 10.6151
R1797 B.n878 B.n97 10.6151
R1798 B.n878 B.n877 10.6151
R1799 B.n877 B.n876 10.6151
R1800 B.n876 B.n99 10.6151
R1801 B.n872 B.n99 10.6151
R1802 B.n872 B.n871 10.6151
R1803 B.n871 B.n870 10.6151
R1804 B.n870 B.n101 10.6151
R1805 B.n866 B.n101 10.6151
R1806 B.n866 B.n865 10.6151
R1807 B.n865 B.n864 10.6151
R1808 B.n864 B.n103 10.6151
R1809 B.n860 B.n103 10.6151
R1810 B.n860 B.n859 10.6151
R1811 B.n859 B.n858 10.6151
R1812 B.n858 B.n105 10.6151
R1813 B.n854 B.n105 10.6151
R1814 B.n854 B.n853 10.6151
R1815 B.n853 B.n852 10.6151
R1816 B.n852 B.n107 10.6151
R1817 B.n848 B.n107 10.6151
R1818 B.n848 B.n847 10.6151
R1819 B.n846 B.n109 10.6151
R1820 B.n842 B.n109 10.6151
R1821 B.n842 B.n841 10.6151
R1822 B.n841 B.n840 10.6151
R1823 B.n840 B.n111 10.6151
R1824 B.n836 B.n111 10.6151
R1825 B.n836 B.n835 10.6151
R1826 B.n835 B.n834 10.6151
R1827 B.n834 B.n113 10.6151
R1828 B.n830 B.n113 10.6151
R1829 B.n830 B.n829 10.6151
R1830 B.n829 B.n828 10.6151
R1831 B.n828 B.n115 10.6151
R1832 B.n824 B.n115 10.6151
R1833 B.n824 B.n823 10.6151
R1834 B.n823 B.n822 10.6151
R1835 B.n822 B.n117 10.6151
R1836 B.n818 B.n117 10.6151
R1837 B.n818 B.n817 10.6151
R1838 B.n817 B.n816 10.6151
R1839 B.n816 B.n119 10.6151
R1840 B.n812 B.n119 10.6151
R1841 B.n812 B.n811 10.6151
R1842 B.n811 B.n810 10.6151
R1843 B.n810 B.n121 10.6151
R1844 B.n806 B.n121 10.6151
R1845 B.n806 B.n805 10.6151
R1846 B.n805 B.n804 10.6151
R1847 B.n804 B.n123 10.6151
R1848 B.n800 B.n123 10.6151
R1849 B.n800 B.n799 10.6151
R1850 B.n799 B.n798 10.6151
R1851 B.n798 B.n125 10.6151
R1852 B.n794 B.n125 10.6151
R1853 B.n794 B.n793 10.6151
R1854 B.n793 B.n792 10.6151
R1855 B.n792 B.n127 10.6151
R1856 B.n788 B.n127 10.6151
R1857 B.n788 B.n787 10.6151
R1858 B.n787 B.n786 10.6151
R1859 B.n786 B.n129 10.6151
R1860 B.n782 B.n129 10.6151
R1861 B.n782 B.n781 10.6151
R1862 B.n781 B.n780 10.6151
R1863 B.n780 B.n131 10.6151
R1864 B.n776 B.n131 10.6151
R1865 B.n776 B.n775 10.6151
R1866 B.n775 B.n774 10.6151
R1867 B.n774 B.n133 10.6151
R1868 B.n770 B.n133 10.6151
R1869 B.n770 B.n769 10.6151
R1870 B.n769 B.n768 10.6151
R1871 B.n768 B.n135 10.6151
R1872 B.n764 B.n135 10.6151
R1873 B.n764 B.n763 10.6151
R1874 B.n763 B.n762 10.6151
R1875 B.n762 B.n137 10.6151
R1876 B.n758 B.n137 10.6151
R1877 B.n758 B.n757 10.6151
R1878 B.n757 B.n756 10.6151
R1879 B.n756 B.n139 10.6151
R1880 B.n752 B.n139 10.6151
R1881 B.n752 B.n751 10.6151
R1882 B.n751 B.n750 10.6151
R1883 B.n750 B.n141 10.6151
R1884 B.n746 B.n141 10.6151
R1885 B.n746 B.n745 10.6151
R1886 B.n745 B.n744 10.6151
R1887 B.n744 B.n143 10.6151
R1888 B.n740 B.n143 10.6151
R1889 B.n740 B.n739 10.6151
R1890 B.n739 B.n738 10.6151
R1891 B.n738 B.n145 10.6151
R1892 B.n734 B.n145 10.6151
R1893 B.n734 B.n733 10.6151
R1894 B.n733 B.n732 10.6151
R1895 B.n732 B.n147 10.6151
R1896 B.n728 B.n147 10.6151
R1897 B.n728 B.n727 10.6151
R1898 B.n727 B.n726 10.6151
R1899 B.n726 B.n149 10.6151
R1900 B.n722 B.n149 10.6151
R1901 B.n722 B.n721 10.6151
R1902 B.n721 B.n720 10.6151
R1903 B.n720 B.n151 10.6151
R1904 B.n716 B.n151 10.6151
R1905 B.n716 B.n715 10.6151
R1906 B.n715 B.n714 10.6151
R1907 B.n714 B.n153 10.6151
R1908 B.n710 B.n153 10.6151
R1909 B.n710 B.n709 10.6151
R1910 B.n709 B.n708 10.6151
R1911 B.n708 B.n155 10.6151
R1912 B.n704 B.n155 10.6151
R1913 B.n704 B.n703 10.6151
R1914 B.n703 B.n702 10.6151
R1915 B.n702 B.n157 10.6151
R1916 B.n698 B.n157 10.6151
R1917 B.n698 B.n697 10.6151
R1918 B.n697 B.n696 10.6151
R1919 B.n696 B.n159 10.6151
R1920 B.n692 B.n159 10.6151
R1921 B.n692 B.n691 10.6151
R1922 B.n691 B.n690 10.6151
R1923 B.n690 B.n161 10.6151
R1924 B.n686 B.n161 10.6151
R1925 B.n686 B.n685 10.6151
R1926 B.n685 B.n684 10.6151
R1927 B.n684 B.n163 10.6151
R1928 B.n680 B.n163 10.6151
R1929 B.n680 B.n679 10.6151
R1930 B.n679 B.n678 10.6151
R1931 B.n678 B.n165 10.6151
R1932 B.n674 B.n165 10.6151
R1933 B.n674 B.n673 10.6151
R1934 B.n673 B.n672 10.6151
R1935 B.n672 B.n167 10.6151
R1936 B.n668 B.n167 10.6151
R1937 B.n668 B.n667 10.6151
R1938 B.n667 B.n666 10.6151
R1939 B.n666 B.n169 10.6151
R1940 B.n662 B.n169 10.6151
R1941 B.n662 B.n661 10.6151
R1942 B.n661 B.n660 10.6151
R1943 B.n660 B.n171 10.6151
R1944 B.n656 B.n171 10.6151
R1945 B.n656 B.n655 10.6151
R1946 B.n655 B.n654 10.6151
R1947 B.n654 B.n173 10.6151
R1948 B.n650 B.n173 10.6151
R1949 B.n650 B.n649 10.6151
R1950 B.n649 B.n648 10.6151
R1951 B.n648 B.n175 10.6151
R1952 B.n644 B.n175 10.6151
R1953 B.n644 B.n643 10.6151
R1954 B.n643 B.n642 10.6151
R1955 B.n642 B.n177 10.6151
R1956 B.n638 B.n177 10.6151
R1957 B.n638 B.n637 10.6151
R1958 B.n637 B.n636 10.6151
R1959 B.n636 B.n179 10.6151
R1960 B.n632 B.n179 10.6151
R1961 B.n632 B.n631 10.6151
R1962 B.n631 B.n630 10.6151
R1963 B.n630 B.n181 10.6151
R1964 B.n626 B.n181 10.6151
R1965 B.n626 B.n625 10.6151
R1966 B.n625 B.n624 10.6151
R1967 B.n624 B.n183 10.6151
R1968 B.n620 B.n183 10.6151
R1969 B.n620 B.n619 10.6151
R1970 B.n619 B.n618 10.6151
R1971 B.n618 B.n185 10.6151
R1972 B.n614 B.n185 10.6151
R1973 B.n614 B.n613 10.6151
R1974 B.n613 B.n612 10.6151
R1975 B.n612 B.n187 10.6151
R1976 B.n608 B.n187 10.6151
R1977 B.n608 B.n607 10.6151
R1978 B.n607 B.n606 10.6151
R1979 B.n606 B.n189 10.6151
R1980 B.n602 B.n189 10.6151
R1981 B.n602 B.n601 10.6151
R1982 B.n293 B.n1 10.6151
R1983 B.n296 B.n293 10.6151
R1984 B.n297 B.n296 10.6151
R1985 B.n298 B.n297 10.6151
R1986 B.n298 B.n291 10.6151
R1987 B.n302 B.n291 10.6151
R1988 B.n303 B.n302 10.6151
R1989 B.n304 B.n303 10.6151
R1990 B.n304 B.n289 10.6151
R1991 B.n308 B.n289 10.6151
R1992 B.n309 B.n308 10.6151
R1993 B.n310 B.n309 10.6151
R1994 B.n310 B.n287 10.6151
R1995 B.n314 B.n287 10.6151
R1996 B.n315 B.n314 10.6151
R1997 B.n316 B.n315 10.6151
R1998 B.n316 B.n285 10.6151
R1999 B.n320 B.n285 10.6151
R2000 B.n321 B.n320 10.6151
R2001 B.n322 B.n321 10.6151
R2002 B.n322 B.n283 10.6151
R2003 B.n326 B.n283 10.6151
R2004 B.n327 B.n326 10.6151
R2005 B.n328 B.n327 10.6151
R2006 B.n328 B.n281 10.6151
R2007 B.n332 B.n281 10.6151
R2008 B.n333 B.n332 10.6151
R2009 B.n334 B.n333 10.6151
R2010 B.n334 B.n279 10.6151
R2011 B.n338 B.n279 10.6151
R2012 B.n339 B.n338 10.6151
R2013 B.n340 B.n339 10.6151
R2014 B.n340 B.n277 10.6151
R2015 B.n344 B.n277 10.6151
R2016 B.n345 B.n344 10.6151
R2017 B.n346 B.n345 10.6151
R2018 B.n346 B.n275 10.6151
R2019 B.n350 B.n275 10.6151
R2020 B.n351 B.n350 10.6151
R2021 B.n352 B.n351 10.6151
R2022 B.n352 B.n273 10.6151
R2023 B.n356 B.n273 10.6151
R2024 B.n357 B.n356 10.6151
R2025 B.n358 B.n357 10.6151
R2026 B.n358 B.n271 10.6151
R2027 B.n362 B.n271 10.6151
R2028 B.n363 B.n362 10.6151
R2029 B.n364 B.n363 10.6151
R2030 B.n364 B.n269 10.6151
R2031 B.n368 B.n269 10.6151
R2032 B.n369 B.n368 10.6151
R2033 B.n370 B.n369 10.6151
R2034 B.n370 B.n267 10.6151
R2035 B.n374 B.n267 10.6151
R2036 B.n375 B.n374 10.6151
R2037 B.n376 B.n375 10.6151
R2038 B.n376 B.n265 10.6151
R2039 B.n380 B.n265 10.6151
R2040 B.n381 B.n380 10.6151
R2041 B.n382 B.n381 10.6151
R2042 B.n382 B.n263 10.6151
R2043 B.n386 B.n263 10.6151
R2044 B.n387 B.n386 10.6151
R2045 B.n388 B.n387 10.6151
R2046 B.n388 B.n261 10.6151
R2047 B.n392 B.n261 10.6151
R2048 B.n393 B.n392 10.6151
R2049 B.n394 B.n393 10.6151
R2050 B.n394 B.n259 10.6151
R2051 B.n398 B.n259 10.6151
R2052 B.n399 B.n398 10.6151
R2053 B.n400 B.n399 10.6151
R2054 B.n400 B.n257 10.6151
R2055 B.n404 B.n257 10.6151
R2056 B.n405 B.n404 10.6151
R2057 B.n406 B.n405 10.6151
R2058 B.n406 B.n255 10.6151
R2059 B.n410 B.n255 10.6151
R2060 B.n411 B.n410 10.6151
R2061 B.n412 B.n411 10.6151
R2062 B.n416 B.n253 10.6151
R2063 B.n417 B.n416 10.6151
R2064 B.n418 B.n417 10.6151
R2065 B.n418 B.n251 10.6151
R2066 B.n422 B.n251 10.6151
R2067 B.n423 B.n422 10.6151
R2068 B.n424 B.n423 10.6151
R2069 B.n424 B.n249 10.6151
R2070 B.n428 B.n249 10.6151
R2071 B.n429 B.n428 10.6151
R2072 B.n430 B.n429 10.6151
R2073 B.n430 B.n247 10.6151
R2074 B.n434 B.n247 10.6151
R2075 B.n435 B.n434 10.6151
R2076 B.n436 B.n435 10.6151
R2077 B.n436 B.n245 10.6151
R2078 B.n440 B.n245 10.6151
R2079 B.n441 B.n440 10.6151
R2080 B.n442 B.n441 10.6151
R2081 B.n442 B.n243 10.6151
R2082 B.n446 B.n243 10.6151
R2083 B.n447 B.n446 10.6151
R2084 B.n448 B.n447 10.6151
R2085 B.n448 B.n241 10.6151
R2086 B.n452 B.n241 10.6151
R2087 B.n453 B.n452 10.6151
R2088 B.n454 B.n453 10.6151
R2089 B.n454 B.n239 10.6151
R2090 B.n458 B.n239 10.6151
R2091 B.n459 B.n458 10.6151
R2092 B.n460 B.n459 10.6151
R2093 B.n460 B.n237 10.6151
R2094 B.n464 B.n237 10.6151
R2095 B.n465 B.n464 10.6151
R2096 B.n466 B.n465 10.6151
R2097 B.n466 B.n235 10.6151
R2098 B.n470 B.n235 10.6151
R2099 B.n471 B.n470 10.6151
R2100 B.n472 B.n471 10.6151
R2101 B.n472 B.n233 10.6151
R2102 B.n476 B.n233 10.6151
R2103 B.n477 B.n476 10.6151
R2104 B.n478 B.n477 10.6151
R2105 B.n478 B.n231 10.6151
R2106 B.n482 B.n231 10.6151
R2107 B.n483 B.n482 10.6151
R2108 B.n484 B.n483 10.6151
R2109 B.n484 B.n229 10.6151
R2110 B.n488 B.n229 10.6151
R2111 B.n489 B.n488 10.6151
R2112 B.n490 B.n489 10.6151
R2113 B.n490 B.n227 10.6151
R2114 B.n494 B.n227 10.6151
R2115 B.n495 B.n494 10.6151
R2116 B.n499 B.n495 10.6151
R2117 B.n503 B.n225 10.6151
R2118 B.n504 B.n503 10.6151
R2119 B.n505 B.n504 10.6151
R2120 B.n505 B.n223 10.6151
R2121 B.n509 B.n223 10.6151
R2122 B.n510 B.n509 10.6151
R2123 B.n511 B.n510 10.6151
R2124 B.n511 B.n221 10.6151
R2125 B.n515 B.n221 10.6151
R2126 B.n518 B.n517 10.6151
R2127 B.n518 B.n217 10.6151
R2128 B.n522 B.n217 10.6151
R2129 B.n523 B.n522 10.6151
R2130 B.n524 B.n523 10.6151
R2131 B.n524 B.n215 10.6151
R2132 B.n528 B.n215 10.6151
R2133 B.n529 B.n528 10.6151
R2134 B.n530 B.n529 10.6151
R2135 B.n530 B.n213 10.6151
R2136 B.n534 B.n213 10.6151
R2137 B.n535 B.n534 10.6151
R2138 B.n536 B.n535 10.6151
R2139 B.n536 B.n211 10.6151
R2140 B.n540 B.n211 10.6151
R2141 B.n541 B.n540 10.6151
R2142 B.n542 B.n541 10.6151
R2143 B.n542 B.n209 10.6151
R2144 B.n546 B.n209 10.6151
R2145 B.n547 B.n546 10.6151
R2146 B.n548 B.n547 10.6151
R2147 B.n548 B.n207 10.6151
R2148 B.n552 B.n207 10.6151
R2149 B.n553 B.n552 10.6151
R2150 B.n554 B.n553 10.6151
R2151 B.n554 B.n205 10.6151
R2152 B.n558 B.n205 10.6151
R2153 B.n559 B.n558 10.6151
R2154 B.n560 B.n559 10.6151
R2155 B.n560 B.n203 10.6151
R2156 B.n564 B.n203 10.6151
R2157 B.n565 B.n564 10.6151
R2158 B.n566 B.n565 10.6151
R2159 B.n566 B.n201 10.6151
R2160 B.n570 B.n201 10.6151
R2161 B.n571 B.n570 10.6151
R2162 B.n572 B.n571 10.6151
R2163 B.n572 B.n199 10.6151
R2164 B.n576 B.n199 10.6151
R2165 B.n577 B.n576 10.6151
R2166 B.n578 B.n577 10.6151
R2167 B.n578 B.n197 10.6151
R2168 B.n582 B.n197 10.6151
R2169 B.n583 B.n582 10.6151
R2170 B.n584 B.n583 10.6151
R2171 B.n584 B.n195 10.6151
R2172 B.n588 B.n195 10.6151
R2173 B.n589 B.n588 10.6151
R2174 B.n590 B.n589 10.6151
R2175 B.n590 B.n193 10.6151
R2176 B.n594 B.n193 10.6151
R2177 B.n595 B.n594 10.6151
R2178 B.n596 B.n595 10.6151
R2179 B.n596 B.n191 10.6151
R2180 B.n600 B.n191 10.6151
R2181 B.n74 B.n70 9.36635
R2182 B.n931 B.n930 9.36635
R2183 B.n499 B.n498 9.36635
R2184 B.n517 B.n516 9.36635
R2185 B.n1153 B.n0 8.11757
R2186 B.n1153 B.n1 8.11757
R2187 B.n945 B.n74 1.24928
R2188 B.n932 B.n931 1.24928
R2189 B.n498 B.n225 1.24928
R2190 B.n516 B.n515 1.24928
C0 VN VTAIL 16.866901f
C1 w_n5962_n4376# VN 13.2036f
C2 B VTAIL 5.39766f
C3 w_n5962_n4376# B 14.0276f
C4 VP VTAIL 16.882f
C5 VDD1 VDD2 2.97547f
C6 w_n5962_n4376# VP 13.9837f
C7 B VN 1.66025f
C8 VP VN 11.136299f
C9 B VP 2.97868f
C10 VTAIL VDD1 12.979f
C11 w_n5962_n4376# VDD1 3.59353f
C12 VTAIL VDD2 13.038401f
C13 w_n5962_n4376# VDD2 3.80101f
C14 VN VDD1 0.156403f
C15 VN VDD2 15.94f
C16 B VDD1 3.36494f
C17 VP VDD1 16.52f
C18 B VDD2 3.53075f
C19 w_n5962_n4376# VTAIL 4.05972f
C20 VP VDD2 0.740263f
C21 VDD2 VSUBS 2.71339f
C22 VDD1 VSUBS 2.595108f
C23 VTAIL VSUBS 1.765073f
C24 VN VSUBS 9.88876f
C25 VP VSUBS 5.9838f
C26 B VSUBS 7.315865f
C27 w_n5962_n4376# VSUBS 0.319301p
C28 B.n0 VSUBS 0.006787f
C29 B.n1 VSUBS 0.006787f
C30 B.n2 VSUBS 0.010038f
C31 B.n3 VSUBS 0.007692f
C32 B.n4 VSUBS 0.007692f
C33 B.n5 VSUBS 0.007692f
C34 B.n6 VSUBS 0.007692f
C35 B.n7 VSUBS 0.007692f
C36 B.n8 VSUBS 0.007692f
C37 B.n9 VSUBS 0.007692f
C38 B.n10 VSUBS 0.007692f
C39 B.n11 VSUBS 0.007692f
C40 B.n12 VSUBS 0.007692f
C41 B.n13 VSUBS 0.007692f
C42 B.n14 VSUBS 0.007692f
C43 B.n15 VSUBS 0.007692f
C44 B.n16 VSUBS 0.007692f
C45 B.n17 VSUBS 0.007692f
C46 B.n18 VSUBS 0.007692f
C47 B.n19 VSUBS 0.007692f
C48 B.n20 VSUBS 0.007692f
C49 B.n21 VSUBS 0.007692f
C50 B.n22 VSUBS 0.007692f
C51 B.n23 VSUBS 0.007692f
C52 B.n24 VSUBS 0.007692f
C53 B.n25 VSUBS 0.007692f
C54 B.n26 VSUBS 0.007692f
C55 B.n27 VSUBS 0.007692f
C56 B.n28 VSUBS 0.007692f
C57 B.n29 VSUBS 0.007692f
C58 B.n30 VSUBS 0.007692f
C59 B.n31 VSUBS 0.007692f
C60 B.n32 VSUBS 0.007692f
C61 B.n33 VSUBS 0.007692f
C62 B.n34 VSUBS 0.007692f
C63 B.n35 VSUBS 0.007692f
C64 B.n36 VSUBS 0.007692f
C65 B.n37 VSUBS 0.007692f
C66 B.n38 VSUBS 0.007692f
C67 B.n39 VSUBS 0.007692f
C68 B.n40 VSUBS 0.007692f
C69 B.n41 VSUBS 0.007692f
C70 B.n42 VSUBS 0.018633f
C71 B.n43 VSUBS 0.007692f
C72 B.n44 VSUBS 0.007692f
C73 B.n45 VSUBS 0.007692f
C74 B.n46 VSUBS 0.007692f
C75 B.n47 VSUBS 0.007692f
C76 B.n48 VSUBS 0.007692f
C77 B.n49 VSUBS 0.007692f
C78 B.n50 VSUBS 0.007692f
C79 B.n51 VSUBS 0.007692f
C80 B.n52 VSUBS 0.007692f
C81 B.n53 VSUBS 0.007692f
C82 B.n54 VSUBS 0.007692f
C83 B.n55 VSUBS 0.007692f
C84 B.n56 VSUBS 0.007692f
C85 B.n57 VSUBS 0.007692f
C86 B.n58 VSUBS 0.007692f
C87 B.n59 VSUBS 0.007692f
C88 B.n60 VSUBS 0.007692f
C89 B.n61 VSUBS 0.007692f
C90 B.n62 VSUBS 0.007692f
C91 B.n63 VSUBS 0.007692f
C92 B.n64 VSUBS 0.007692f
C93 B.n65 VSUBS 0.007692f
C94 B.n66 VSUBS 0.007692f
C95 B.n67 VSUBS 0.007692f
C96 B.n68 VSUBS 0.007692f
C97 B.n69 VSUBS 0.007692f
C98 B.n70 VSUBS 0.007239f
C99 B.n71 VSUBS 0.007692f
C100 B.t4 VSUBS 0.629604f
C101 B.t5 VSUBS 0.661346f
C102 B.t3 VSUBS 3.28052f
C103 B.n72 VSUBS 0.406606f
C104 B.n73 VSUBS 0.084833f
C105 B.n74 VSUBS 0.017821f
C106 B.n75 VSUBS 0.007692f
C107 B.n76 VSUBS 0.007692f
C108 B.n77 VSUBS 0.007692f
C109 B.n78 VSUBS 0.007692f
C110 B.t1 VSUBS 0.629582f
C111 B.t2 VSUBS 0.66133f
C112 B.t0 VSUBS 3.28052f
C113 B.n79 VSUBS 0.406622f
C114 B.n80 VSUBS 0.084855f
C115 B.n81 VSUBS 0.007692f
C116 B.n82 VSUBS 0.007692f
C117 B.n83 VSUBS 0.007692f
C118 B.n84 VSUBS 0.007692f
C119 B.n85 VSUBS 0.007692f
C120 B.n86 VSUBS 0.007692f
C121 B.n87 VSUBS 0.007692f
C122 B.n88 VSUBS 0.007692f
C123 B.n89 VSUBS 0.007692f
C124 B.n90 VSUBS 0.007692f
C125 B.n91 VSUBS 0.007692f
C126 B.n92 VSUBS 0.007692f
C127 B.n93 VSUBS 0.007692f
C128 B.n94 VSUBS 0.007692f
C129 B.n95 VSUBS 0.007692f
C130 B.n96 VSUBS 0.007692f
C131 B.n97 VSUBS 0.007692f
C132 B.n98 VSUBS 0.007692f
C133 B.n99 VSUBS 0.007692f
C134 B.n100 VSUBS 0.007692f
C135 B.n101 VSUBS 0.007692f
C136 B.n102 VSUBS 0.007692f
C137 B.n103 VSUBS 0.007692f
C138 B.n104 VSUBS 0.007692f
C139 B.n105 VSUBS 0.007692f
C140 B.n106 VSUBS 0.007692f
C141 B.n107 VSUBS 0.007692f
C142 B.n108 VSUBS 0.019148f
C143 B.n109 VSUBS 0.007692f
C144 B.n110 VSUBS 0.007692f
C145 B.n111 VSUBS 0.007692f
C146 B.n112 VSUBS 0.007692f
C147 B.n113 VSUBS 0.007692f
C148 B.n114 VSUBS 0.007692f
C149 B.n115 VSUBS 0.007692f
C150 B.n116 VSUBS 0.007692f
C151 B.n117 VSUBS 0.007692f
C152 B.n118 VSUBS 0.007692f
C153 B.n119 VSUBS 0.007692f
C154 B.n120 VSUBS 0.007692f
C155 B.n121 VSUBS 0.007692f
C156 B.n122 VSUBS 0.007692f
C157 B.n123 VSUBS 0.007692f
C158 B.n124 VSUBS 0.007692f
C159 B.n125 VSUBS 0.007692f
C160 B.n126 VSUBS 0.007692f
C161 B.n127 VSUBS 0.007692f
C162 B.n128 VSUBS 0.007692f
C163 B.n129 VSUBS 0.007692f
C164 B.n130 VSUBS 0.007692f
C165 B.n131 VSUBS 0.007692f
C166 B.n132 VSUBS 0.007692f
C167 B.n133 VSUBS 0.007692f
C168 B.n134 VSUBS 0.007692f
C169 B.n135 VSUBS 0.007692f
C170 B.n136 VSUBS 0.007692f
C171 B.n137 VSUBS 0.007692f
C172 B.n138 VSUBS 0.007692f
C173 B.n139 VSUBS 0.007692f
C174 B.n140 VSUBS 0.007692f
C175 B.n141 VSUBS 0.007692f
C176 B.n142 VSUBS 0.007692f
C177 B.n143 VSUBS 0.007692f
C178 B.n144 VSUBS 0.007692f
C179 B.n145 VSUBS 0.007692f
C180 B.n146 VSUBS 0.007692f
C181 B.n147 VSUBS 0.007692f
C182 B.n148 VSUBS 0.007692f
C183 B.n149 VSUBS 0.007692f
C184 B.n150 VSUBS 0.007692f
C185 B.n151 VSUBS 0.007692f
C186 B.n152 VSUBS 0.007692f
C187 B.n153 VSUBS 0.007692f
C188 B.n154 VSUBS 0.007692f
C189 B.n155 VSUBS 0.007692f
C190 B.n156 VSUBS 0.007692f
C191 B.n157 VSUBS 0.007692f
C192 B.n158 VSUBS 0.007692f
C193 B.n159 VSUBS 0.007692f
C194 B.n160 VSUBS 0.007692f
C195 B.n161 VSUBS 0.007692f
C196 B.n162 VSUBS 0.007692f
C197 B.n163 VSUBS 0.007692f
C198 B.n164 VSUBS 0.007692f
C199 B.n165 VSUBS 0.007692f
C200 B.n166 VSUBS 0.007692f
C201 B.n167 VSUBS 0.007692f
C202 B.n168 VSUBS 0.007692f
C203 B.n169 VSUBS 0.007692f
C204 B.n170 VSUBS 0.007692f
C205 B.n171 VSUBS 0.007692f
C206 B.n172 VSUBS 0.007692f
C207 B.n173 VSUBS 0.007692f
C208 B.n174 VSUBS 0.007692f
C209 B.n175 VSUBS 0.007692f
C210 B.n176 VSUBS 0.007692f
C211 B.n177 VSUBS 0.007692f
C212 B.n178 VSUBS 0.007692f
C213 B.n179 VSUBS 0.007692f
C214 B.n180 VSUBS 0.007692f
C215 B.n181 VSUBS 0.007692f
C216 B.n182 VSUBS 0.007692f
C217 B.n183 VSUBS 0.007692f
C218 B.n184 VSUBS 0.007692f
C219 B.n185 VSUBS 0.007692f
C220 B.n186 VSUBS 0.007692f
C221 B.n187 VSUBS 0.007692f
C222 B.n188 VSUBS 0.007692f
C223 B.n189 VSUBS 0.007692f
C224 B.n190 VSUBS 0.018633f
C225 B.n191 VSUBS 0.007692f
C226 B.n192 VSUBS 0.007692f
C227 B.n193 VSUBS 0.007692f
C228 B.n194 VSUBS 0.007692f
C229 B.n195 VSUBS 0.007692f
C230 B.n196 VSUBS 0.007692f
C231 B.n197 VSUBS 0.007692f
C232 B.n198 VSUBS 0.007692f
C233 B.n199 VSUBS 0.007692f
C234 B.n200 VSUBS 0.007692f
C235 B.n201 VSUBS 0.007692f
C236 B.n202 VSUBS 0.007692f
C237 B.n203 VSUBS 0.007692f
C238 B.n204 VSUBS 0.007692f
C239 B.n205 VSUBS 0.007692f
C240 B.n206 VSUBS 0.007692f
C241 B.n207 VSUBS 0.007692f
C242 B.n208 VSUBS 0.007692f
C243 B.n209 VSUBS 0.007692f
C244 B.n210 VSUBS 0.007692f
C245 B.n211 VSUBS 0.007692f
C246 B.n212 VSUBS 0.007692f
C247 B.n213 VSUBS 0.007692f
C248 B.n214 VSUBS 0.007692f
C249 B.n215 VSUBS 0.007692f
C250 B.n216 VSUBS 0.007692f
C251 B.n217 VSUBS 0.007692f
C252 B.n218 VSUBS 0.007692f
C253 B.t11 VSUBS 0.629582f
C254 B.t10 VSUBS 0.66133f
C255 B.t9 VSUBS 3.28052f
C256 B.n219 VSUBS 0.406622f
C257 B.n220 VSUBS 0.084855f
C258 B.n221 VSUBS 0.007692f
C259 B.n222 VSUBS 0.007692f
C260 B.n223 VSUBS 0.007692f
C261 B.n224 VSUBS 0.007692f
C262 B.n225 VSUBS 0.004298f
C263 B.n226 VSUBS 0.007692f
C264 B.n227 VSUBS 0.007692f
C265 B.n228 VSUBS 0.007692f
C266 B.n229 VSUBS 0.007692f
C267 B.n230 VSUBS 0.007692f
C268 B.n231 VSUBS 0.007692f
C269 B.n232 VSUBS 0.007692f
C270 B.n233 VSUBS 0.007692f
C271 B.n234 VSUBS 0.007692f
C272 B.n235 VSUBS 0.007692f
C273 B.n236 VSUBS 0.007692f
C274 B.n237 VSUBS 0.007692f
C275 B.n238 VSUBS 0.007692f
C276 B.n239 VSUBS 0.007692f
C277 B.n240 VSUBS 0.007692f
C278 B.n241 VSUBS 0.007692f
C279 B.n242 VSUBS 0.007692f
C280 B.n243 VSUBS 0.007692f
C281 B.n244 VSUBS 0.007692f
C282 B.n245 VSUBS 0.007692f
C283 B.n246 VSUBS 0.007692f
C284 B.n247 VSUBS 0.007692f
C285 B.n248 VSUBS 0.007692f
C286 B.n249 VSUBS 0.007692f
C287 B.n250 VSUBS 0.007692f
C288 B.n251 VSUBS 0.007692f
C289 B.n252 VSUBS 0.007692f
C290 B.n253 VSUBS 0.019148f
C291 B.n254 VSUBS 0.007692f
C292 B.n255 VSUBS 0.007692f
C293 B.n256 VSUBS 0.007692f
C294 B.n257 VSUBS 0.007692f
C295 B.n258 VSUBS 0.007692f
C296 B.n259 VSUBS 0.007692f
C297 B.n260 VSUBS 0.007692f
C298 B.n261 VSUBS 0.007692f
C299 B.n262 VSUBS 0.007692f
C300 B.n263 VSUBS 0.007692f
C301 B.n264 VSUBS 0.007692f
C302 B.n265 VSUBS 0.007692f
C303 B.n266 VSUBS 0.007692f
C304 B.n267 VSUBS 0.007692f
C305 B.n268 VSUBS 0.007692f
C306 B.n269 VSUBS 0.007692f
C307 B.n270 VSUBS 0.007692f
C308 B.n271 VSUBS 0.007692f
C309 B.n272 VSUBS 0.007692f
C310 B.n273 VSUBS 0.007692f
C311 B.n274 VSUBS 0.007692f
C312 B.n275 VSUBS 0.007692f
C313 B.n276 VSUBS 0.007692f
C314 B.n277 VSUBS 0.007692f
C315 B.n278 VSUBS 0.007692f
C316 B.n279 VSUBS 0.007692f
C317 B.n280 VSUBS 0.007692f
C318 B.n281 VSUBS 0.007692f
C319 B.n282 VSUBS 0.007692f
C320 B.n283 VSUBS 0.007692f
C321 B.n284 VSUBS 0.007692f
C322 B.n285 VSUBS 0.007692f
C323 B.n286 VSUBS 0.007692f
C324 B.n287 VSUBS 0.007692f
C325 B.n288 VSUBS 0.007692f
C326 B.n289 VSUBS 0.007692f
C327 B.n290 VSUBS 0.007692f
C328 B.n291 VSUBS 0.007692f
C329 B.n292 VSUBS 0.007692f
C330 B.n293 VSUBS 0.007692f
C331 B.n294 VSUBS 0.007692f
C332 B.n295 VSUBS 0.007692f
C333 B.n296 VSUBS 0.007692f
C334 B.n297 VSUBS 0.007692f
C335 B.n298 VSUBS 0.007692f
C336 B.n299 VSUBS 0.007692f
C337 B.n300 VSUBS 0.007692f
C338 B.n301 VSUBS 0.007692f
C339 B.n302 VSUBS 0.007692f
C340 B.n303 VSUBS 0.007692f
C341 B.n304 VSUBS 0.007692f
C342 B.n305 VSUBS 0.007692f
C343 B.n306 VSUBS 0.007692f
C344 B.n307 VSUBS 0.007692f
C345 B.n308 VSUBS 0.007692f
C346 B.n309 VSUBS 0.007692f
C347 B.n310 VSUBS 0.007692f
C348 B.n311 VSUBS 0.007692f
C349 B.n312 VSUBS 0.007692f
C350 B.n313 VSUBS 0.007692f
C351 B.n314 VSUBS 0.007692f
C352 B.n315 VSUBS 0.007692f
C353 B.n316 VSUBS 0.007692f
C354 B.n317 VSUBS 0.007692f
C355 B.n318 VSUBS 0.007692f
C356 B.n319 VSUBS 0.007692f
C357 B.n320 VSUBS 0.007692f
C358 B.n321 VSUBS 0.007692f
C359 B.n322 VSUBS 0.007692f
C360 B.n323 VSUBS 0.007692f
C361 B.n324 VSUBS 0.007692f
C362 B.n325 VSUBS 0.007692f
C363 B.n326 VSUBS 0.007692f
C364 B.n327 VSUBS 0.007692f
C365 B.n328 VSUBS 0.007692f
C366 B.n329 VSUBS 0.007692f
C367 B.n330 VSUBS 0.007692f
C368 B.n331 VSUBS 0.007692f
C369 B.n332 VSUBS 0.007692f
C370 B.n333 VSUBS 0.007692f
C371 B.n334 VSUBS 0.007692f
C372 B.n335 VSUBS 0.007692f
C373 B.n336 VSUBS 0.007692f
C374 B.n337 VSUBS 0.007692f
C375 B.n338 VSUBS 0.007692f
C376 B.n339 VSUBS 0.007692f
C377 B.n340 VSUBS 0.007692f
C378 B.n341 VSUBS 0.007692f
C379 B.n342 VSUBS 0.007692f
C380 B.n343 VSUBS 0.007692f
C381 B.n344 VSUBS 0.007692f
C382 B.n345 VSUBS 0.007692f
C383 B.n346 VSUBS 0.007692f
C384 B.n347 VSUBS 0.007692f
C385 B.n348 VSUBS 0.007692f
C386 B.n349 VSUBS 0.007692f
C387 B.n350 VSUBS 0.007692f
C388 B.n351 VSUBS 0.007692f
C389 B.n352 VSUBS 0.007692f
C390 B.n353 VSUBS 0.007692f
C391 B.n354 VSUBS 0.007692f
C392 B.n355 VSUBS 0.007692f
C393 B.n356 VSUBS 0.007692f
C394 B.n357 VSUBS 0.007692f
C395 B.n358 VSUBS 0.007692f
C396 B.n359 VSUBS 0.007692f
C397 B.n360 VSUBS 0.007692f
C398 B.n361 VSUBS 0.007692f
C399 B.n362 VSUBS 0.007692f
C400 B.n363 VSUBS 0.007692f
C401 B.n364 VSUBS 0.007692f
C402 B.n365 VSUBS 0.007692f
C403 B.n366 VSUBS 0.007692f
C404 B.n367 VSUBS 0.007692f
C405 B.n368 VSUBS 0.007692f
C406 B.n369 VSUBS 0.007692f
C407 B.n370 VSUBS 0.007692f
C408 B.n371 VSUBS 0.007692f
C409 B.n372 VSUBS 0.007692f
C410 B.n373 VSUBS 0.007692f
C411 B.n374 VSUBS 0.007692f
C412 B.n375 VSUBS 0.007692f
C413 B.n376 VSUBS 0.007692f
C414 B.n377 VSUBS 0.007692f
C415 B.n378 VSUBS 0.007692f
C416 B.n379 VSUBS 0.007692f
C417 B.n380 VSUBS 0.007692f
C418 B.n381 VSUBS 0.007692f
C419 B.n382 VSUBS 0.007692f
C420 B.n383 VSUBS 0.007692f
C421 B.n384 VSUBS 0.007692f
C422 B.n385 VSUBS 0.007692f
C423 B.n386 VSUBS 0.007692f
C424 B.n387 VSUBS 0.007692f
C425 B.n388 VSUBS 0.007692f
C426 B.n389 VSUBS 0.007692f
C427 B.n390 VSUBS 0.007692f
C428 B.n391 VSUBS 0.007692f
C429 B.n392 VSUBS 0.007692f
C430 B.n393 VSUBS 0.007692f
C431 B.n394 VSUBS 0.007692f
C432 B.n395 VSUBS 0.007692f
C433 B.n396 VSUBS 0.007692f
C434 B.n397 VSUBS 0.007692f
C435 B.n398 VSUBS 0.007692f
C436 B.n399 VSUBS 0.007692f
C437 B.n400 VSUBS 0.007692f
C438 B.n401 VSUBS 0.007692f
C439 B.n402 VSUBS 0.007692f
C440 B.n403 VSUBS 0.007692f
C441 B.n404 VSUBS 0.007692f
C442 B.n405 VSUBS 0.007692f
C443 B.n406 VSUBS 0.007692f
C444 B.n407 VSUBS 0.007692f
C445 B.n408 VSUBS 0.007692f
C446 B.n409 VSUBS 0.007692f
C447 B.n410 VSUBS 0.007692f
C448 B.n411 VSUBS 0.007692f
C449 B.n412 VSUBS 0.018633f
C450 B.n413 VSUBS 0.018633f
C451 B.n414 VSUBS 0.019148f
C452 B.n415 VSUBS 0.007692f
C453 B.n416 VSUBS 0.007692f
C454 B.n417 VSUBS 0.007692f
C455 B.n418 VSUBS 0.007692f
C456 B.n419 VSUBS 0.007692f
C457 B.n420 VSUBS 0.007692f
C458 B.n421 VSUBS 0.007692f
C459 B.n422 VSUBS 0.007692f
C460 B.n423 VSUBS 0.007692f
C461 B.n424 VSUBS 0.007692f
C462 B.n425 VSUBS 0.007692f
C463 B.n426 VSUBS 0.007692f
C464 B.n427 VSUBS 0.007692f
C465 B.n428 VSUBS 0.007692f
C466 B.n429 VSUBS 0.007692f
C467 B.n430 VSUBS 0.007692f
C468 B.n431 VSUBS 0.007692f
C469 B.n432 VSUBS 0.007692f
C470 B.n433 VSUBS 0.007692f
C471 B.n434 VSUBS 0.007692f
C472 B.n435 VSUBS 0.007692f
C473 B.n436 VSUBS 0.007692f
C474 B.n437 VSUBS 0.007692f
C475 B.n438 VSUBS 0.007692f
C476 B.n439 VSUBS 0.007692f
C477 B.n440 VSUBS 0.007692f
C478 B.n441 VSUBS 0.007692f
C479 B.n442 VSUBS 0.007692f
C480 B.n443 VSUBS 0.007692f
C481 B.n444 VSUBS 0.007692f
C482 B.n445 VSUBS 0.007692f
C483 B.n446 VSUBS 0.007692f
C484 B.n447 VSUBS 0.007692f
C485 B.n448 VSUBS 0.007692f
C486 B.n449 VSUBS 0.007692f
C487 B.n450 VSUBS 0.007692f
C488 B.n451 VSUBS 0.007692f
C489 B.n452 VSUBS 0.007692f
C490 B.n453 VSUBS 0.007692f
C491 B.n454 VSUBS 0.007692f
C492 B.n455 VSUBS 0.007692f
C493 B.n456 VSUBS 0.007692f
C494 B.n457 VSUBS 0.007692f
C495 B.n458 VSUBS 0.007692f
C496 B.n459 VSUBS 0.007692f
C497 B.n460 VSUBS 0.007692f
C498 B.n461 VSUBS 0.007692f
C499 B.n462 VSUBS 0.007692f
C500 B.n463 VSUBS 0.007692f
C501 B.n464 VSUBS 0.007692f
C502 B.n465 VSUBS 0.007692f
C503 B.n466 VSUBS 0.007692f
C504 B.n467 VSUBS 0.007692f
C505 B.n468 VSUBS 0.007692f
C506 B.n469 VSUBS 0.007692f
C507 B.n470 VSUBS 0.007692f
C508 B.n471 VSUBS 0.007692f
C509 B.n472 VSUBS 0.007692f
C510 B.n473 VSUBS 0.007692f
C511 B.n474 VSUBS 0.007692f
C512 B.n475 VSUBS 0.007692f
C513 B.n476 VSUBS 0.007692f
C514 B.n477 VSUBS 0.007692f
C515 B.n478 VSUBS 0.007692f
C516 B.n479 VSUBS 0.007692f
C517 B.n480 VSUBS 0.007692f
C518 B.n481 VSUBS 0.007692f
C519 B.n482 VSUBS 0.007692f
C520 B.n483 VSUBS 0.007692f
C521 B.n484 VSUBS 0.007692f
C522 B.n485 VSUBS 0.007692f
C523 B.n486 VSUBS 0.007692f
C524 B.n487 VSUBS 0.007692f
C525 B.n488 VSUBS 0.007692f
C526 B.n489 VSUBS 0.007692f
C527 B.n490 VSUBS 0.007692f
C528 B.n491 VSUBS 0.007692f
C529 B.n492 VSUBS 0.007692f
C530 B.n493 VSUBS 0.007692f
C531 B.n494 VSUBS 0.007692f
C532 B.n495 VSUBS 0.007692f
C533 B.t8 VSUBS 0.629604f
C534 B.t7 VSUBS 0.661346f
C535 B.t6 VSUBS 3.28052f
C536 B.n496 VSUBS 0.406606f
C537 B.n497 VSUBS 0.084833f
C538 B.n498 VSUBS 0.017821f
C539 B.n499 VSUBS 0.007239f
C540 B.n500 VSUBS 0.007692f
C541 B.n501 VSUBS 0.007692f
C542 B.n502 VSUBS 0.007692f
C543 B.n503 VSUBS 0.007692f
C544 B.n504 VSUBS 0.007692f
C545 B.n505 VSUBS 0.007692f
C546 B.n506 VSUBS 0.007692f
C547 B.n507 VSUBS 0.007692f
C548 B.n508 VSUBS 0.007692f
C549 B.n509 VSUBS 0.007692f
C550 B.n510 VSUBS 0.007692f
C551 B.n511 VSUBS 0.007692f
C552 B.n512 VSUBS 0.007692f
C553 B.n513 VSUBS 0.007692f
C554 B.n514 VSUBS 0.007692f
C555 B.n515 VSUBS 0.004298f
C556 B.n516 VSUBS 0.017821f
C557 B.n517 VSUBS 0.007239f
C558 B.n518 VSUBS 0.007692f
C559 B.n519 VSUBS 0.007692f
C560 B.n520 VSUBS 0.007692f
C561 B.n521 VSUBS 0.007692f
C562 B.n522 VSUBS 0.007692f
C563 B.n523 VSUBS 0.007692f
C564 B.n524 VSUBS 0.007692f
C565 B.n525 VSUBS 0.007692f
C566 B.n526 VSUBS 0.007692f
C567 B.n527 VSUBS 0.007692f
C568 B.n528 VSUBS 0.007692f
C569 B.n529 VSUBS 0.007692f
C570 B.n530 VSUBS 0.007692f
C571 B.n531 VSUBS 0.007692f
C572 B.n532 VSUBS 0.007692f
C573 B.n533 VSUBS 0.007692f
C574 B.n534 VSUBS 0.007692f
C575 B.n535 VSUBS 0.007692f
C576 B.n536 VSUBS 0.007692f
C577 B.n537 VSUBS 0.007692f
C578 B.n538 VSUBS 0.007692f
C579 B.n539 VSUBS 0.007692f
C580 B.n540 VSUBS 0.007692f
C581 B.n541 VSUBS 0.007692f
C582 B.n542 VSUBS 0.007692f
C583 B.n543 VSUBS 0.007692f
C584 B.n544 VSUBS 0.007692f
C585 B.n545 VSUBS 0.007692f
C586 B.n546 VSUBS 0.007692f
C587 B.n547 VSUBS 0.007692f
C588 B.n548 VSUBS 0.007692f
C589 B.n549 VSUBS 0.007692f
C590 B.n550 VSUBS 0.007692f
C591 B.n551 VSUBS 0.007692f
C592 B.n552 VSUBS 0.007692f
C593 B.n553 VSUBS 0.007692f
C594 B.n554 VSUBS 0.007692f
C595 B.n555 VSUBS 0.007692f
C596 B.n556 VSUBS 0.007692f
C597 B.n557 VSUBS 0.007692f
C598 B.n558 VSUBS 0.007692f
C599 B.n559 VSUBS 0.007692f
C600 B.n560 VSUBS 0.007692f
C601 B.n561 VSUBS 0.007692f
C602 B.n562 VSUBS 0.007692f
C603 B.n563 VSUBS 0.007692f
C604 B.n564 VSUBS 0.007692f
C605 B.n565 VSUBS 0.007692f
C606 B.n566 VSUBS 0.007692f
C607 B.n567 VSUBS 0.007692f
C608 B.n568 VSUBS 0.007692f
C609 B.n569 VSUBS 0.007692f
C610 B.n570 VSUBS 0.007692f
C611 B.n571 VSUBS 0.007692f
C612 B.n572 VSUBS 0.007692f
C613 B.n573 VSUBS 0.007692f
C614 B.n574 VSUBS 0.007692f
C615 B.n575 VSUBS 0.007692f
C616 B.n576 VSUBS 0.007692f
C617 B.n577 VSUBS 0.007692f
C618 B.n578 VSUBS 0.007692f
C619 B.n579 VSUBS 0.007692f
C620 B.n580 VSUBS 0.007692f
C621 B.n581 VSUBS 0.007692f
C622 B.n582 VSUBS 0.007692f
C623 B.n583 VSUBS 0.007692f
C624 B.n584 VSUBS 0.007692f
C625 B.n585 VSUBS 0.007692f
C626 B.n586 VSUBS 0.007692f
C627 B.n587 VSUBS 0.007692f
C628 B.n588 VSUBS 0.007692f
C629 B.n589 VSUBS 0.007692f
C630 B.n590 VSUBS 0.007692f
C631 B.n591 VSUBS 0.007692f
C632 B.n592 VSUBS 0.007692f
C633 B.n593 VSUBS 0.007692f
C634 B.n594 VSUBS 0.007692f
C635 B.n595 VSUBS 0.007692f
C636 B.n596 VSUBS 0.007692f
C637 B.n597 VSUBS 0.007692f
C638 B.n598 VSUBS 0.007692f
C639 B.n599 VSUBS 0.019148f
C640 B.n600 VSUBS 0.018303f
C641 B.n601 VSUBS 0.019478f
C642 B.n602 VSUBS 0.007692f
C643 B.n603 VSUBS 0.007692f
C644 B.n604 VSUBS 0.007692f
C645 B.n605 VSUBS 0.007692f
C646 B.n606 VSUBS 0.007692f
C647 B.n607 VSUBS 0.007692f
C648 B.n608 VSUBS 0.007692f
C649 B.n609 VSUBS 0.007692f
C650 B.n610 VSUBS 0.007692f
C651 B.n611 VSUBS 0.007692f
C652 B.n612 VSUBS 0.007692f
C653 B.n613 VSUBS 0.007692f
C654 B.n614 VSUBS 0.007692f
C655 B.n615 VSUBS 0.007692f
C656 B.n616 VSUBS 0.007692f
C657 B.n617 VSUBS 0.007692f
C658 B.n618 VSUBS 0.007692f
C659 B.n619 VSUBS 0.007692f
C660 B.n620 VSUBS 0.007692f
C661 B.n621 VSUBS 0.007692f
C662 B.n622 VSUBS 0.007692f
C663 B.n623 VSUBS 0.007692f
C664 B.n624 VSUBS 0.007692f
C665 B.n625 VSUBS 0.007692f
C666 B.n626 VSUBS 0.007692f
C667 B.n627 VSUBS 0.007692f
C668 B.n628 VSUBS 0.007692f
C669 B.n629 VSUBS 0.007692f
C670 B.n630 VSUBS 0.007692f
C671 B.n631 VSUBS 0.007692f
C672 B.n632 VSUBS 0.007692f
C673 B.n633 VSUBS 0.007692f
C674 B.n634 VSUBS 0.007692f
C675 B.n635 VSUBS 0.007692f
C676 B.n636 VSUBS 0.007692f
C677 B.n637 VSUBS 0.007692f
C678 B.n638 VSUBS 0.007692f
C679 B.n639 VSUBS 0.007692f
C680 B.n640 VSUBS 0.007692f
C681 B.n641 VSUBS 0.007692f
C682 B.n642 VSUBS 0.007692f
C683 B.n643 VSUBS 0.007692f
C684 B.n644 VSUBS 0.007692f
C685 B.n645 VSUBS 0.007692f
C686 B.n646 VSUBS 0.007692f
C687 B.n647 VSUBS 0.007692f
C688 B.n648 VSUBS 0.007692f
C689 B.n649 VSUBS 0.007692f
C690 B.n650 VSUBS 0.007692f
C691 B.n651 VSUBS 0.007692f
C692 B.n652 VSUBS 0.007692f
C693 B.n653 VSUBS 0.007692f
C694 B.n654 VSUBS 0.007692f
C695 B.n655 VSUBS 0.007692f
C696 B.n656 VSUBS 0.007692f
C697 B.n657 VSUBS 0.007692f
C698 B.n658 VSUBS 0.007692f
C699 B.n659 VSUBS 0.007692f
C700 B.n660 VSUBS 0.007692f
C701 B.n661 VSUBS 0.007692f
C702 B.n662 VSUBS 0.007692f
C703 B.n663 VSUBS 0.007692f
C704 B.n664 VSUBS 0.007692f
C705 B.n665 VSUBS 0.007692f
C706 B.n666 VSUBS 0.007692f
C707 B.n667 VSUBS 0.007692f
C708 B.n668 VSUBS 0.007692f
C709 B.n669 VSUBS 0.007692f
C710 B.n670 VSUBS 0.007692f
C711 B.n671 VSUBS 0.007692f
C712 B.n672 VSUBS 0.007692f
C713 B.n673 VSUBS 0.007692f
C714 B.n674 VSUBS 0.007692f
C715 B.n675 VSUBS 0.007692f
C716 B.n676 VSUBS 0.007692f
C717 B.n677 VSUBS 0.007692f
C718 B.n678 VSUBS 0.007692f
C719 B.n679 VSUBS 0.007692f
C720 B.n680 VSUBS 0.007692f
C721 B.n681 VSUBS 0.007692f
C722 B.n682 VSUBS 0.007692f
C723 B.n683 VSUBS 0.007692f
C724 B.n684 VSUBS 0.007692f
C725 B.n685 VSUBS 0.007692f
C726 B.n686 VSUBS 0.007692f
C727 B.n687 VSUBS 0.007692f
C728 B.n688 VSUBS 0.007692f
C729 B.n689 VSUBS 0.007692f
C730 B.n690 VSUBS 0.007692f
C731 B.n691 VSUBS 0.007692f
C732 B.n692 VSUBS 0.007692f
C733 B.n693 VSUBS 0.007692f
C734 B.n694 VSUBS 0.007692f
C735 B.n695 VSUBS 0.007692f
C736 B.n696 VSUBS 0.007692f
C737 B.n697 VSUBS 0.007692f
C738 B.n698 VSUBS 0.007692f
C739 B.n699 VSUBS 0.007692f
C740 B.n700 VSUBS 0.007692f
C741 B.n701 VSUBS 0.007692f
C742 B.n702 VSUBS 0.007692f
C743 B.n703 VSUBS 0.007692f
C744 B.n704 VSUBS 0.007692f
C745 B.n705 VSUBS 0.007692f
C746 B.n706 VSUBS 0.007692f
C747 B.n707 VSUBS 0.007692f
C748 B.n708 VSUBS 0.007692f
C749 B.n709 VSUBS 0.007692f
C750 B.n710 VSUBS 0.007692f
C751 B.n711 VSUBS 0.007692f
C752 B.n712 VSUBS 0.007692f
C753 B.n713 VSUBS 0.007692f
C754 B.n714 VSUBS 0.007692f
C755 B.n715 VSUBS 0.007692f
C756 B.n716 VSUBS 0.007692f
C757 B.n717 VSUBS 0.007692f
C758 B.n718 VSUBS 0.007692f
C759 B.n719 VSUBS 0.007692f
C760 B.n720 VSUBS 0.007692f
C761 B.n721 VSUBS 0.007692f
C762 B.n722 VSUBS 0.007692f
C763 B.n723 VSUBS 0.007692f
C764 B.n724 VSUBS 0.007692f
C765 B.n725 VSUBS 0.007692f
C766 B.n726 VSUBS 0.007692f
C767 B.n727 VSUBS 0.007692f
C768 B.n728 VSUBS 0.007692f
C769 B.n729 VSUBS 0.007692f
C770 B.n730 VSUBS 0.007692f
C771 B.n731 VSUBS 0.007692f
C772 B.n732 VSUBS 0.007692f
C773 B.n733 VSUBS 0.007692f
C774 B.n734 VSUBS 0.007692f
C775 B.n735 VSUBS 0.007692f
C776 B.n736 VSUBS 0.007692f
C777 B.n737 VSUBS 0.007692f
C778 B.n738 VSUBS 0.007692f
C779 B.n739 VSUBS 0.007692f
C780 B.n740 VSUBS 0.007692f
C781 B.n741 VSUBS 0.007692f
C782 B.n742 VSUBS 0.007692f
C783 B.n743 VSUBS 0.007692f
C784 B.n744 VSUBS 0.007692f
C785 B.n745 VSUBS 0.007692f
C786 B.n746 VSUBS 0.007692f
C787 B.n747 VSUBS 0.007692f
C788 B.n748 VSUBS 0.007692f
C789 B.n749 VSUBS 0.007692f
C790 B.n750 VSUBS 0.007692f
C791 B.n751 VSUBS 0.007692f
C792 B.n752 VSUBS 0.007692f
C793 B.n753 VSUBS 0.007692f
C794 B.n754 VSUBS 0.007692f
C795 B.n755 VSUBS 0.007692f
C796 B.n756 VSUBS 0.007692f
C797 B.n757 VSUBS 0.007692f
C798 B.n758 VSUBS 0.007692f
C799 B.n759 VSUBS 0.007692f
C800 B.n760 VSUBS 0.007692f
C801 B.n761 VSUBS 0.007692f
C802 B.n762 VSUBS 0.007692f
C803 B.n763 VSUBS 0.007692f
C804 B.n764 VSUBS 0.007692f
C805 B.n765 VSUBS 0.007692f
C806 B.n766 VSUBS 0.007692f
C807 B.n767 VSUBS 0.007692f
C808 B.n768 VSUBS 0.007692f
C809 B.n769 VSUBS 0.007692f
C810 B.n770 VSUBS 0.007692f
C811 B.n771 VSUBS 0.007692f
C812 B.n772 VSUBS 0.007692f
C813 B.n773 VSUBS 0.007692f
C814 B.n774 VSUBS 0.007692f
C815 B.n775 VSUBS 0.007692f
C816 B.n776 VSUBS 0.007692f
C817 B.n777 VSUBS 0.007692f
C818 B.n778 VSUBS 0.007692f
C819 B.n779 VSUBS 0.007692f
C820 B.n780 VSUBS 0.007692f
C821 B.n781 VSUBS 0.007692f
C822 B.n782 VSUBS 0.007692f
C823 B.n783 VSUBS 0.007692f
C824 B.n784 VSUBS 0.007692f
C825 B.n785 VSUBS 0.007692f
C826 B.n786 VSUBS 0.007692f
C827 B.n787 VSUBS 0.007692f
C828 B.n788 VSUBS 0.007692f
C829 B.n789 VSUBS 0.007692f
C830 B.n790 VSUBS 0.007692f
C831 B.n791 VSUBS 0.007692f
C832 B.n792 VSUBS 0.007692f
C833 B.n793 VSUBS 0.007692f
C834 B.n794 VSUBS 0.007692f
C835 B.n795 VSUBS 0.007692f
C836 B.n796 VSUBS 0.007692f
C837 B.n797 VSUBS 0.007692f
C838 B.n798 VSUBS 0.007692f
C839 B.n799 VSUBS 0.007692f
C840 B.n800 VSUBS 0.007692f
C841 B.n801 VSUBS 0.007692f
C842 B.n802 VSUBS 0.007692f
C843 B.n803 VSUBS 0.007692f
C844 B.n804 VSUBS 0.007692f
C845 B.n805 VSUBS 0.007692f
C846 B.n806 VSUBS 0.007692f
C847 B.n807 VSUBS 0.007692f
C848 B.n808 VSUBS 0.007692f
C849 B.n809 VSUBS 0.007692f
C850 B.n810 VSUBS 0.007692f
C851 B.n811 VSUBS 0.007692f
C852 B.n812 VSUBS 0.007692f
C853 B.n813 VSUBS 0.007692f
C854 B.n814 VSUBS 0.007692f
C855 B.n815 VSUBS 0.007692f
C856 B.n816 VSUBS 0.007692f
C857 B.n817 VSUBS 0.007692f
C858 B.n818 VSUBS 0.007692f
C859 B.n819 VSUBS 0.007692f
C860 B.n820 VSUBS 0.007692f
C861 B.n821 VSUBS 0.007692f
C862 B.n822 VSUBS 0.007692f
C863 B.n823 VSUBS 0.007692f
C864 B.n824 VSUBS 0.007692f
C865 B.n825 VSUBS 0.007692f
C866 B.n826 VSUBS 0.007692f
C867 B.n827 VSUBS 0.007692f
C868 B.n828 VSUBS 0.007692f
C869 B.n829 VSUBS 0.007692f
C870 B.n830 VSUBS 0.007692f
C871 B.n831 VSUBS 0.007692f
C872 B.n832 VSUBS 0.007692f
C873 B.n833 VSUBS 0.007692f
C874 B.n834 VSUBS 0.007692f
C875 B.n835 VSUBS 0.007692f
C876 B.n836 VSUBS 0.007692f
C877 B.n837 VSUBS 0.007692f
C878 B.n838 VSUBS 0.007692f
C879 B.n839 VSUBS 0.007692f
C880 B.n840 VSUBS 0.007692f
C881 B.n841 VSUBS 0.007692f
C882 B.n842 VSUBS 0.007692f
C883 B.n843 VSUBS 0.007692f
C884 B.n844 VSUBS 0.007692f
C885 B.n845 VSUBS 0.018633f
C886 B.n846 VSUBS 0.018633f
C887 B.n847 VSUBS 0.019148f
C888 B.n848 VSUBS 0.007692f
C889 B.n849 VSUBS 0.007692f
C890 B.n850 VSUBS 0.007692f
C891 B.n851 VSUBS 0.007692f
C892 B.n852 VSUBS 0.007692f
C893 B.n853 VSUBS 0.007692f
C894 B.n854 VSUBS 0.007692f
C895 B.n855 VSUBS 0.007692f
C896 B.n856 VSUBS 0.007692f
C897 B.n857 VSUBS 0.007692f
C898 B.n858 VSUBS 0.007692f
C899 B.n859 VSUBS 0.007692f
C900 B.n860 VSUBS 0.007692f
C901 B.n861 VSUBS 0.007692f
C902 B.n862 VSUBS 0.007692f
C903 B.n863 VSUBS 0.007692f
C904 B.n864 VSUBS 0.007692f
C905 B.n865 VSUBS 0.007692f
C906 B.n866 VSUBS 0.007692f
C907 B.n867 VSUBS 0.007692f
C908 B.n868 VSUBS 0.007692f
C909 B.n869 VSUBS 0.007692f
C910 B.n870 VSUBS 0.007692f
C911 B.n871 VSUBS 0.007692f
C912 B.n872 VSUBS 0.007692f
C913 B.n873 VSUBS 0.007692f
C914 B.n874 VSUBS 0.007692f
C915 B.n875 VSUBS 0.007692f
C916 B.n876 VSUBS 0.007692f
C917 B.n877 VSUBS 0.007692f
C918 B.n878 VSUBS 0.007692f
C919 B.n879 VSUBS 0.007692f
C920 B.n880 VSUBS 0.007692f
C921 B.n881 VSUBS 0.007692f
C922 B.n882 VSUBS 0.007692f
C923 B.n883 VSUBS 0.007692f
C924 B.n884 VSUBS 0.007692f
C925 B.n885 VSUBS 0.007692f
C926 B.n886 VSUBS 0.007692f
C927 B.n887 VSUBS 0.007692f
C928 B.n888 VSUBS 0.007692f
C929 B.n889 VSUBS 0.007692f
C930 B.n890 VSUBS 0.007692f
C931 B.n891 VSUBS 0.007692f
C932 B.n892 VSUBS 0.007692f
C933 B.n893 VSUBS 0.007692f
C934 B.n894 VSUBS 0.007692f
C935 B.n895 VSUBS 0.007692f
C936 B.n896 VSUBS 0.007692f
C937 B.n897 VSUBS 0.007692f
C938 B.n898 VSUBS 0.007692f
C939 B.n899 VSUBS 0.007692f
C940 B.n900 VSUBS 0.007692f
C941 B.n901 VSUBS 0.007692f
C942 B.n902 VSUBS 0.007692f
C943 B.n903 VSUBS 0.007692f
C944 B.n904 VSUBS 0.007692f
C945 B.n905 VSUBS 0.007692f
C946 B.n906 VSUBS 0.007692f
C947 B.n907 VSUBS 0.007692f
C948 B.n908 VSUBS 0.007692f
C949 B.n909 VSUBS 0.007692f
C950 B.n910 VSUBS 0.007692f
C951 B.n911 VSUBS 0.007692f
C952 B.n912 VSUBS 0.007692f
C953 B.n913 VSUBS 0.007692f
C954 B.n914 VSUBS 0.007692f
C955 B.n915 VSUBS 0.007692f
C956 B.n916 VSUBS 0.007692f
C957 B.n917 VSUBS 0.007692f
C958 B.n918 VSUBS 0.007692f
C959 B.n919 VSUBS 0.007692f
C960 B.n920 VSUBS 0.007692f
C961 B.n921 VSUBS 0.007692f
C962 B.n922 VSUBS 0.007692f
C963 B.n923 VSUBS 0.007692f
C964 B.n924 VSUBS 0.007692f
C965 B.n925 VSUBS 0.007692f
C966 B.n926 VSUBS 0.007692f
C967 B.n927 VSUBS 0.007692f
C968 B.n928 VSUBS 0.007692f
C969 B.n929 VSUBS 0.007692f
C970 B.n930 VSUBS 0.007239f
C971 B.n931 VSUBS 0.017821f
C972 B.n932 VSUBS 0.004298f
C973 B.n933 VSUBS 0.007692f
C974 B.n934 VSUBS 0.007692f
C975 B.n935 VSUBS 0.007692f
C976 B.n936 VSUBS 0.007692f
C977 B.n937 VSUBS 0.007692f
C978 B.n938 VSUBS 0.007692f
C979 B.n939 VSUBS 0.007692f
C980 B.n940 VSUBS 0.007692f
C981 B.n941 VSUBS 0.007692f
C982 B.n942 VSUBS 0.007692f
C983 B.n943 VSUBS 0.007692f
C984 B.n944 VSUBS 0.007692f
C985 B.n945 VSUBS 0.004298f
C986 B.n946 VSUBS 0.007692f
C987 B.n947 VSUBS 0.007692f
C988 B.n948 VSUBS 0.007692f
C989 B.n949 VSUBS 0.007692f
C990 B.n950 VSUBS 0.007692f
C991 B.n951 VSUBS 0.007692f
C992 B.n952 VSUBS 0.007692f
C993 B.n953 VSUBS 0.007692f
C994 B.n954 VSUBS 0.007692f
C995 B.n955 VSUBS 0.007692f
C996 B.n956 VSUBS 0.007692f
C997 B.n957 VSUBS 0.007692f
C998 B.n958 VSUBS 0.007692f
C999 B.n959 VSUBS 0.007692f
C1000 B.n960 VSUBS 0.007692f
C1001 B.n961 VSUBS 0.007692f
C1002 B.n962 VSUBS 0.007692f
C1003 B.n963 VSUBS 0.007692f
C1004 B.n964 VSUBS 0.007692f
C1005 B.n965 VSUBS 0.007692f
C1006 B.n966 VSUBS 0.007692f
C1007 B.n967 VSUBS 0.007692f
C1008 B.n968 VSUBS 0.007692f
C1009 B.n969 VSUBS 0.007692f
C1010 B.n970 VSUBS 0.007692f
C1011 B.n971 VSUBS 0.007692f
C1012 B.n972 VSUBS 0.007692f
C1013 B.n973 VSUBS 0.007692f
C1014 B.n974 VSUBS 0.007692f
C1015 B.n975 VSUBS 0.007692f
C1016 B.n976 VSUBS 0.007692f
C1017 B.n977 VSUBS 0.007692f
C1018 B.n978 VSUBS 0.007692f
C1019 B.n979 VSUBS 0.007692f
C1020 B.n980 VSUBS 0.007692f
C1021 B.n981 VSUBS 0.007692f
C1022 B.n982 VSUBS 0.007692f
C1023 B.n983 VSUBS 0.007692f
C1024 B.n984 VSUBS 0.007692f
C1025 B.n985 VSUBS 0.007692f
C1026 B.n986 VSUBS 0.007692f
C1027 B.n987 VSUBS 0.007692f
C1028 B.n988 VSUBS 0.007692f
C1029 B.n989 VSUBS 0.007692f
C1030 B.n990 VSUBS 0.007692f
C1031 B.n991 VSUBS 0.007692f
C1032 B.n992 VSUBS 0.007692f
C1033 B.n993 VSUBS 0.007692f
C1034 B.n994 VSUBS 0.007692f
C1035 B.n995 VSUBS 0.007692f
C1036 B.n996 VSUBS 0.007692f
C1037 B.n997 VSUBS 0.007692f
C1038 B.n998 VSUBS 0.007692f
C1039 B.n999 VSUBS 0.007692f
C1040 B.n1000 VSUBS 0.007692f
C1041 B.n1001 VSUBS 0.007692f
C1042 B.n1002 VSUBS 0.007692f
C1043 B.n1003 VSUBS 0.007692f
C1044 B.n1004 VSUBS 0.007692f
C1045 B.n1005 VSUBS 0.007692f
C1046 B.n1006 VSUBS 0.007692f
C1047 B.n1007 VSUBS 0.007692f
C1048 B.n1008 VSUBS 0.007692f
C1049 B.n1009 VSUBS 0.007692f
C1050 B.n1010 VSUBS 0.007692f
C1051 B.n1011 VSUBS 0.007692f
C1052 B.n1012 VSUBS 0.007692f
C1053 B.n1013 VSUBS 0.007692f
C1054 B.n1014 VSUBS 0.007692f
C1055 B.n1015 VSUBS 0.007692f
C1056 B.n1016 VSUBS 0.007692f
C1057 B.n1017 VSUBS 0.007692f
C1058 B.n1018 VSUBS 0.007692f
C1059 B.n1019 VSUBS 0.007692f
C1060 B.n1020 VSUBS 0.007692f
C1061 B.n1021 VSUBS 0.007692f
C1062 B.n1022 VSUBS 0.007692f
C1063 B.n1023 VSUBS 0.007692f
C1064 B.n1024 VSUBS 0.007692f
C1065 B.n1025 VSUBS 0.007692f
C1066 B.n1026 VSUBS 0.007692f
C1067 B.n1027 VSUBS 0.007692f
C1068 B.n1028 VSUBS 0.007692f
C1069 B.n1029 VSUBS 0.019148f
C1070 B.n1030 VSUBS 0.019148f
C1071 B.n1031 VSUBS 0.018633f
C1072 B.n1032 VSUBS 0.007692f
C1073 B.n1033 VSUBS 0.007692f
C1074 B.n1034 VSUBS 0.007692f
C1075 B.n1035 VSUBS 0.007692f
C1076 B.n1036 VSUBS 0.007692f
C1077 B.n1037 VSUBS 0.007692f
C1078 B.n1038 VSUBS 0.007692f
C1079 B.n1039 VSUBS 0.007692f
C1080 B.n1040 VSUBS 0.007692f
C1081 B.n1041 VSUBS 0.007692f
C1082 B.n1042 VSUBS 0.007692f
C1083 B.n1043 VSUBS 0.007692f
C1084 B.n1044 VSUBS 0.007692f
C1085 B.n1045 VSUBS 0.007692f
C1086 B.n1046 VSUBS 0.007692f
C1087 B.n1047 VSUBS 0.007692f
C1088 B.n1048 VSUBS 0.007692f
C1089 B.n1049 VSUBS 0.007692f
C1090 B.n1050 VSUBS 0.007692f
C1091 B.n1051 VSUBS 0.007692f
C1092 B.n1052 VSUBS 0.007692f
C1093 B.n1053 VSUBS 0.007692f
C1094 B.n1054 VSUBS 0.007692f
C1095 B.n1055 VSUBS 0.007692f
C1096 B.n1056 VSUBS 0.007692f
C1097 B.n1057 VSUBS 0.007692f
C1098 B.n1058 VSUBS 0.007692f
C1099 B.n1059 VSUBS 0.007692f
C1100 B.n1060 VSUBS 0.007692f
C1101 B.n1061 VSUBS 0.007692f
C1102 B.n1062 VSUBS 0.007692f
C1103 B.n1063 VSUBS 0.007692f
C1104 B.n1064 VSUBS 0.007692f
C1105 B.n1065 VSUBS 0.007692f
C1106 B.n1066 VSUBS 0.007692f
C1107 B.n1067 VSUBS 0.007692f
C1108 B.n1068 VSUBS 0.007692f
C1109 B.n1069 VSUBS 0.007692f
C1110 B.n1070 VSUBS 0.007692f
C1111 B.n1071 VSUBS 0.007692f
C1112 B.n1072 VSUBS 0.007692f
C1113 B.n1073 VSUBS 0.007692f
C1114 B.n1074 VSUBS 0.007692f
C1115 B.n1075 VSUBS 0.007692f
C1116 B.n1076 VSUBS 0.007692f
C1117 B.n1077 VSUBS 0.007692f
C1118 B.n1078 VSUBS 0.007692f
C1119 B.n1079 VSUBS 0.007692f
C1120 B.n1080 VSUBS 0.007692f
C1121 B.n1081 VSUBS 0.007692f
C1122 B.n1082 VSUBS 0.007692f
C1123 B.n1083 VSUBS 0.007692f
C1124 B.n1084 VSUBS 0.007692f
C1125 B.n1085 VSUBS 0.007692f
C1126 B.n1086 VSUBS 0.007692f
C1127 B.n1087 VSUBS 0.007692f
C1128 B.n1088 VSUBS 0.007692f
C1129 B.n1089 VSUBS 0.007692f
C1130 B.n1090 VSUBS 0.007692f
C1131 B.n1091 VSUBS 0.007692f
C1132 B.n1092 VSUBS 0.007692f
C1133 B.n1093 VSUBS 0.007692f
C1134 B.n1094 VSUBS 0.007692f
C1135 B.n1095 VSUBS 0.007692f
C1136 B.n1096 VSUBS 0.007692f
C1137 B.n1097 VSUBS 0.007692f
C1138 B.n1098 VSUBS 0.007692f
C1139 B.n1099 VSUBS 0.007692f
C1140 B.n1100 VSUBS 0.007692f
C1141 B.n1101 VSUBS 0.007692f
C1142 B.n1102 VSUBS 0.007692f
C1143 B.n1103 VSUBS 0.007692f
C1144 B.n1104 VSUBS 0.007692f
C1145 B.n1105 VSUBS 0.007692f
C1146 B.n1106 VSUBS 0.007692f
C1147 B.n1107 VSUBS 0.007692f
C1148 B.n1108 VSUBS 0.007692f
C1149 B.n1109 VSUBS 0.007692f
C1150 B.n1110 VSUBS 0.007692f
C1151 B.n1111 VSUBS 0.007692f
C1152 B.n1112 VSUBS 0.007692f
C1153 B.n1113 VSUBS 0.007692f
C1154 B.n1114 VSUBS 0.007692f
C1155 B.n1115 VSUBS 0.007692f
C1156 B.n1116 VSUBS 0.007692f
C1157 B.n1117 VSUBS 0.007692f
C1158 B.n1118 VSUBS 0.007692f
C1159 B.n1119 VSUBS 0.007692f
C1160 B.n1120 VSUBS 0.007692f
C1161 B.n1121 VSUBS 0.007692f
C1162 B.n1122 VSUBS 0.007692f
C1163 B.n1123 VSUBS 0.007692f
C1164 B.n1124 VSUBS 0.007692f
C1165 B.n1125 VSUBS 0.007692f
C1166 B.n1126 VSUBS 0.007692f
C1167 B.n1127 VSUBS 0.007692f
C1168 B.n1128 VSUBS 0.007692f
C1169 B.n1129 VSUBS 0.007692f
C1170 B.n1130 VSUBS 0.007692f
C1171 B.n1131 VSUBS 0.007692f
C1172 B.n1132 VSUBS 0.007692f
C1173 B.n1133 VSUBS 0.007692f
C1174 B.n1134 VSUBS 0.007692f
C1175 B.n1135 VSUBS 0.007692f
C1176 B.n1136 VSUBS 0.007692f
C1177 B.n1137 VSUBS 0.007692f
C1178 B.n1138 VSUBS 0.007692f
C1179 B.n1139 VSUBS 0.007692f
C1180 B.n1140 VSUBS 0.007692f
C1181 B.n1141 VSUBS 0.007692f
C1182 B.n1142 VSUBS 0.007692f
C1183 B.n1143 VSUBS 0.007692f
C1184 B.n1144 VSUBS 0.007692f
C1185 B.n1145 VSUBS 0.007692f
C1186 B.n1146 VSUBS 0.007692f
C1187 B.n1147 VSUBS 0.007692f
C1188 B.n1148 VSUBS 0.007692f
C1189 B.n1149 VSUBS 0.007692f
C1190 B.n1150 VSUBS 0.007692f
C1191 B.n1151 VSUBS 0.010038f
C1192 B.n1152 VSUBS 0.010692f
C1193 B.n1153 VSUBS 0.021263f
C1194 VDD2.t6 VSUBS 4.27311f
C1195 VDD2.t8 VSUBS 0.395665f
C1196 VDD2.t2 VSUBS 0.395665f
C1197 VDD2.n0 VSUBS 3.25117f
C1198 VDD2.n1 VSUBS 2.00535f
C1199 VDD2.t0 VSUBS 0.395665f
C1200 VDD2.t1 VSUBS 0.395665f
C1201 VDD2.n2 VSUBS 3.29625f
C1202 VDD2.n3 VSUBS 4.87486f
C1203 VDD2.t9 VSUBS 4.22115f
C1204 VDD2.n4 VSUBS 5.0636f
C1205 VDD2.t7 VSUBS 0.395665f
C1206 VDD2.t5 VSUBS 0.395665f
C1207 VDD2.n5 VSUBS 3.25118f
C1208 VDD2.n6 VSUBS 1.01835f
C1209 VDD2.t3 VSUBS 0.395665f
C1210 VDD2.t4 VSUBS 0.395665f
C1211 VDD2.n7 VSUBS 3.29617f
C1212 VN.t8 VSUBS 3.68204f
C1213 VN.n0 VSUBS 1.34833f
C1214 VN.n1 VSUBS 0.020533f
C1215 VN.n2 VSUBS 0.040785f
C1216 VN.n3 VSUBS 0.020533f
C1217 VN.n4 VSUBS 0.038077f
C1218 VN.n5 VSUBS 0.020533f
C1219 VN.t9 VSUBS 3.68204f
C1220 VN.n6 VSUBS 0.038077f
C1221 VN.n7 VSUBS 0.020533f
C1222 VN.n8 VSUBS 0.038077f
C1223 VN.n9 VSUBS 0.020533f
C1224 VN.t7 VSUBS 3.68204f
C1225 VN.n10 VSUBS 0.038077f
C1226 VN.n11 VSUBS 0.020533f
C1227 VN.n12 VSUBS 0.038077f
C1228 VN.t3 VSUBS 4.02025f
C1229 VN.n13 VSUBS 1.28509f
C1230 VN.t1 VSUBS 3.68204f
C1231 VN.n14 VSUBS 1.35057f
C1232 VN.n15 VSUBS 0.034694f
C1233 VN.n16 VSUBS 0.264206f
C1234 VN.n17 VSUBS 0.020533f
C1235 VN.n18 VSUBS 0.020533f
C1236 VN.n19 VSUBS 0.038077f
C1237 VN.n20 VSUBS 0.025304f
C1238 VN.n21 VSUBS 0.034393f
C1239 VN.n22 VSUBS 0.020533f
C1240 VN.n23 VSUBS 0.020533f
C1241 VN.n24 VSUBS 0.020533f
C1242 VN.n25 VSUBS 0.038077f
C1243 VN.n26 VSUBS 0.028678f
C1244 VN.n27 VSUBS 1.27063f
C1245 VN.n28 VSUBS 0.028678f
C1246 VN.n29 VSUBS 0.020533f
C1247 VN.n30 VSUBS 0.020533f
C1248 VN.n31 VSUBS 0.020533f
C1249 VN.n32 VSUBS 0.038077f
C1250 VN.n33 VSUBS 0.034393f
C1251 VN.n34 VSUBS 0.025304f
C1252 VN.n35 VSUBS 0.020533f
C1253 VN.n36 VSUBS 0.020533f
C1254 VN.n37 VSUBS 0.020533f
C1255 VN.n38 VSUBS 0.038077f
C1256 VN.n39 VSUBS 0.034694f
C1257 VN.n40 VSUBS 1.27063f
C1258 VN.n41 VSUBS 0.022663f
C1259 VN.n42 VSUBS 0.020533f
C1260 VN.n43 VSUBS 0.020533f
C1261 VN.n44 VSUBS 0.020533f
C1262 VN.n45 VSUBS 0.038077f
C1263 VN.n46 VSUBS 0.040378f
C1264 VN.n47 VSUBS 0.01661f
C1265 VN.n48 VSUBS 0.020533f
C1266 VN.n49 VSUBS 0.020533f
C1267 VN.n50 VSUBS 0.020533f
C1268 VN.n51 VSUBS 0.038077f
C1269 VN.n52 VSUBS 0.038077f
C1270 VN.n53 VSUBS 0.021911f
C1271 VN.n54 VSUBS 0.033135f
C1272 VN.n55 VSUBS 0.062998f
C1273 VN.t0 VSUBS 3.68204f
C1274 VN.n56 VSUBS 1.34833f
C1275 VN.n57 VSUBS 0.020533f
C1276 VN.n58 VSUBS 0.040785f
C1277 VN.n59 VSUBS 0.020533f
C1278 VN.n60 VSUBS 0.038077f
C1279 VN.n61 VSUBS 0.020533f
C1280 VN.t2 VSUBS 3.68204f
C1281 VN.n62 VSUBS 0.038077f
C1282 VN.n63 VSUBS 0.020533f
C1283 VN.n64 VSUBS 0.038077f
C1284 VN.n65 VSUBS 0.020533f
C1285 VN.t4 VSUBS 3.68204f
C1286 VN.n66 VSUBS 0.038077f
C1287 VN.n67 VSUBS 0.020533f
C1288 VN.n68 VSUBS 0.038077f
C1289 VN.t5 VSUBS 4.02025f
C1290 VN.n69 VSUBS 1.28509f
C1291 VN.t6 VSUBS 3.68204f
C1292 VN.n70 VSUBS 1.35057f
C1293 VN.n71 VSUBS 0.034694f
C1294 VN.n72 VSUBS 0.264206f
C1295 VN.n73 VSUBS 0.020533f
C1296 VN.n74 VSUBS 0.020533f
C1297 VN.n75 VSUBS 0.038077f
C1298 VN.n76 VSUBS 0.025304f
C1299 VN.n77 VSUBS 0.034393f
C1300 VN.n78 VSUBS 0.020533f
C1301 VN.n79 VSUBS 0.020533f
C1302 VN.n80 VSUBS 0.020533f
C1303 VN.n81 VSUBS 0.038077f
C1304 VN.n82 VSUBS 0.028678f
C1305 VN.n83 VSUBS 1.27063f
C1306 VN.n84 VSUBS 0.028678f
C1307 VN.n85 VSUBS 0.020533f
C1308 VN.n86 VSUBS 0.020533f
C1309 VN.n87 VSUBS 0.020533f
C1310 VN.n88 VSUBS 0.038077f
C1311 VN.n89 VSUBS 0.034393f
C1312 VN.n90 VSUBS 0.025304f
C1313 VN.n91 VSUBS 0.020533f
C1314 VN.n92 VSUBS 0.020533f
C1315 VN.n93 VSUBS 0.020533f
C1316 VN.n94 VSUBS 0.038077f
C1317 VN.n95 VSUBS 0.034694f
C1318 VN.n96 VSUBS 1.27063f
C1319 VN.n97 VSUBS 0.022663f
C1320 VN.n98 VSUBS 0.020533f
C1321 VN.n99 VSUBS 0.020533f
C1322 VN.n100 VSUBS 0.020533f
C1323 VN.n101 VSUBS 0.038077f
C1324 VN.n102 VSUBS 0.040378f
C1325 VN.n103 VSUBS 0.01661f
C1326 VN.n104 VSUBS 0.020533f
C1327 VN.n105 VSUBS 0.020533f
C1328 VN.n106 VSUBS 0.020533f
C1329 VN.n107 VSUBS 0.038077f
C1330 VN.n108 VSUBS 0.038077f
C1331 VN.n109 VSUBS 0.021911f
C1332 VN.n110 VSUBS 0.033135f
C1333 VN.n111 VSUBS 1.64882f
C1334 VDD1.t9 VSUBS 4.29394f
C1335 VDD1.t7 VSUBS 0.397593f
C1336 VDD1.t8 VSUBS 0.397593f
C1337 VDD1.n0 VSUBS 3.26701f
C1338 VDD1.n1 VSUBS 2.02508f
C1339 VDD1.t0 VSUBS 4.29392f
C1340 VDD1.t4 VSUBS 0.397593f
C1341 VDD1.t1 VSUBS 0.397593f
C1342 VDD1.n2 VSUBS 3.26701f
C1343 VDD1.n3 VSUBS 2.01512f
C1344 VDD1.t3 VSUBS 0.397593f
C1345 VDD1.t2 VSUBS 0.397593f
C1346 VDD1.n4 VSUBS 3.31231f
C1347 VDD1.n5 VSUBS 5.09077f
C1348 VDD1.t5 VSUBS 0.397593f
C1349 VDD1.t6 VSUBS 0.397593f
C1350 VDD1.n6 VSUBS 3.267f
C1351 VDD1.n7 VSUBS 5.1459f
C1352 VTAIL.t8 VSUBS 0.382264f
C1353 VTAIL.t5 VSUBS 0.382264f
C1354 VTAIL.n0 VSUBS 2.95395f
C1355 VTAIL.n1 VSUBS 1.17535f
C1356 VTAIL.t10 VSUBS 3.86415f
C1357 VTAIL.n2 VSUBS 1.38437f
C1358 VTAIL.t17 VSUBS 0.382264f
C1359 VTAIL.t18 VSUBS 0.382264f
C1360 VTAIL.n3 VSUBS 2.95395f
C1361 VTAIL.n4 VSUBS 1.37308f
C1362 VTAIL.t9 VSUBS 0.382264f
C1363 VTAIL.t12 VSUBS 0.382264f
C1364 VTAIL.n5 VSUBS 2.95395f
C1365 VTAIL.n6 VSUBS 3.43046f
C1366 VTAIL.t7 VSUBS 0.382264f
C1367 VTAIL.t2 VSUBS 0.382264f
C1368 VTAIL.n7 VSUBS 2.95396f
C1369 VTAIL.n8 VSUBS 3.43045f
C1370 VTAIL.t1 VSUBS 0.382264f
C1371 VTAIL.t19 VSUBS 0.382264f
C1372 VTAIL.n9 VSUBS 2.95396f
C1373 VTAIL.n10 VSUBS 1.37307f
C1374 VTAIL.t6 VSUBS 3.86419f
C1375 VTAIL.n11 VSUBS 1.38434f
C1376 VTAIL.t11 VSUBS 0.382264f
C1377 VTAIL.t13 VSUBS 0.382264f
C1378 VTAIL.n12 VSUBS 2.95396f
C1379 VTAIL.n13 VSUBS 1.25203f
C1380 VTAIL.t14 VSUBS 0.382264f
C1381 VTAIL.t16 VSUBS 0.382264f
C1382 VTAIL.n14 VSUBS 2.95396f
C1383 VTAIL.n15 VSUBS 1.37307f
C1384 VTAIL.t15 VSUBS 3.86415f
C1385 VTAIL.n16 VSUBS 3.23475f
C1386 VTAIL.t3 VSUBS 3.86415f
C1387 VTAIL.n17 VSUBS 3.23475f
C1388 VTAIL.t4 VSUBS 0.382264f
C1389 VTAIL.t0 VSUBS 0.382264f
C1390 VTAIL.n18 VSUBS 2.95395f
C1391 VTAIL.n19 VSUBS 1.12173f
C1392 VP.t7 VSUBS 3.96778f
C1393 VP.n0 VSUBS 1.45296f
C1394 VP.n1 VSUBS 0.022127f
C1395 VP.n2 VSUBS 0.04395f
C1396 VP.n3 VSUBS 0.022127f
C1397 VP.n4 VSUBS 0.041032f
C1398 VP.n5 VSUBS 0.022127f
C1399 VP.t6 VSUBS 3.96778f
C1400 VP.n6 VSUBS 0.041032f
C1401 VP.n7 VSUBS 0.022127f
C1402 VP.n8 VSUBS 0.041032f
C1403 VP.n9 VSUBS 0.022127f
C1404 VP.t8 VSUBS 3.96778f
C1405 VP.n10 VSUBS 0.041032f
C1406 VP.n11 VSUBS 0.022127f
C1407 VP.n12 VSUBS 0.041032f
C1408 VP.n13 VSUBS 0.022127f
C1409 VP.t5 VSUBS 3.96778f
C1410 VP.n14 VSUBS 0.041032f
C1411 VP.n15 VSUBS 0.022127f
C1412 VP.n16 VSUBS 0.041032f
C1413 VP.n17 VSUBS 0.035707f
C1414 VP.t9 VSUBS 3.96778f
C1415 VP.t3 VSUBS 3.96778f
C1416 VP.n18 VSUBS 1.45296f
C1417 VP.n19 VSUBS 0.022127f
C1418 VP.n20 VSUBS 0.04395f
C1419 VP.n21 VSUBS 0.022127f
C1420 VP.n22 VSUBS 0.041032f
C1421 VP.n23 VSUBS 0.022127f
C1422 VP.t4 VSUBS 3.96778f
C1423 VP.n24 VSUBS 0.041032f
C1424 VP.n25 VSUBS 0.022127f
C1425 VP.n26 VSUBS 0.041032f
C1426 VP.n27 VSUBS 0.022127f
C1427 VP.t1 VSUBS 3.96778f
C1428 VP.n28 VSUBS 0.041032f
C1429 VP.n29 VSUBS 0.022127f
C1430 VP.n30 VSUBS 0.041032f
C1431 VP.t0 VSUBS 4.33223f
C1432 VP.n31 VSUBS 1.38482f
C1433 VP.t2 VSUBS 3.96778f
C1434 VP.n32 VSUBS 1.45538f
C1435 VP.n33 VSUBS 0.037386f
C1436 VP.n34 VSUBS 0.28471f
C1437 VP.n35 VSUBS 0.022127f
C1438 VP.n36 VSUBS 0.022127f
C1439 VP.n37 VSUBS 0.041032f
C1440 VP.n38 VSUBS 0.027267f
C1441 VP.n39 VSUBS 0.037062f
C1442 VP.n40 VSUBS 0.022127f
C1443 VP.n41 VSUBS 0.022127f
C1444 VP.n42 VSUBS 0.022127f
C1445 VP.n43 VSUBS 0.041032f
C1446 VP.n44 VSUBS 0.030904f
C1447 VP.n45 VSUBS 1.36924f
C1448 VP.n46 VSUBS 0.030904f
C1449 VP.n47 VSUBS 0.022127f
C1450 VP.n48 VSUBS 0.022127f
C1451 VP.n49 VSUBS 0.022127f
C1452 VP.n50 VSUBS 0.041032f
C1453 VP.n51 VSUBS 0.037062f
C1454 VP.n52 VSUBS 0.027267f
C1455 VP.n53 VSUBS 0.022127f
C1456 VP.n54 VSUBS 0.022127f
C1457 VP.n55 VSUBS 0.022127f
C1458 VP.n56 VSUBS 0.041032f
C1459 VP.n57 VSUBS 0.037386f
C1460 VP.n58 VSUBS 1.36924f
C1461 VP.n59 VSUBS 0.024422f
C1462 VP.n60 VSUBS 0.022127f
C1463 VP.n61 VSUBS 0.022127f
C1464 VP.n62 VSUBS 0.022127f
C1465 VP.n63 VSUBS 0.041032f
C1466 VP.n64 VSUBS 0.043512f
C1467 VP.n65 VSUBS 0.017899f
C1468 VP.n66 VSUBS 0.022127f
C1469 VP.n67 VSUBS 0.022127f
C1470 VP.n68 VSUBS 0.022127f
C1471 VP.n69 VSUBS 0.041032f
C1472 VP.n70 VSUBS 0.041032f
C1473 VP.n71 VSUBS 0.023612f
C1474 VP.n72 VSUBS 0.035707f
C1475 VP.n73 VSUBS 1.76839f
C1476 VP.n74 VSUBS 1.78092f
C1477 VP.n75 VSUBS 1.45296f
C1478 VP.n76 VSUBS 0.023612f
C1479 VP.n77 VSUBS 0.041032f
C1480 VP.n78 VSUBS 0.022127f
C1481 VP.n79 VSUBS 0.022127f
C1482 VP.n80 VSUBS 0.022127f
C1483 VP.n81 VSUBS 0.04395f
C1484 VP.n82 VSUBS 0.017899f
C1485 VP.n83 VSUBS 0.043512f
C1486 VP.n84 VSUBS 0.022127f
C1487 VP.n85 VSUBS 0.022127f
C1488 VP.n86 VSUBS 0.022127f
C1489 VP.n87 VSUBS 0.041032f
C1490 VP.n88 VSUBS 0.024422f
C1491 VP.n89 VSUBS 1.36924f
C1492 VP.n90 VSUBS 0.037386f
C1493 VP.n91 VSUBS 0.022127f
C1494 VP.n92 VSUBS 0.022127f
C1495 VP.n93 VSUBS 0.022127f
C1496 VP.n94 VSUBS 0.041032f
C1497 VP.n95 VSUBS 0.027267f
C1498 VP.n96 VSUBS 0.037062f
C1499 VP.n97 VSUBS 0.022127f
C1500 VP.n98 VSUBS 0.022127f
C1501 VP.n99 VSUBS 0.022127f
C1502 VP.n100 VSUBS 0.041032f
C1503 VP.n101 VSUBS 0.030904f
C1504 VP.n102 VSUBS 1.36924f
C1505 VP.n103 VSUBS 0.030904f
C1506 VP.n104 VSUBS 0.022127f
C1507 VP.n105 VSUBS 0.022127f
C1508 VP.n106 VSUBS 0.022127f
C1509 VP.n107 VSUBS 0.041032f
C1510 VP.n108 VSUBS 0.037062f
C1511 VP.n109 VSUBS 0.027267f
C1512 VP.n110 VSUBS 0.022127f
C1513 VP.n111 VSUBS 0.022127f
C1514 VP.n112 VSUBS 0.022127f
C1515 VP.n113 VSUBS 0.041032f
C1516 VP.n114 VSUBS 0.037386f
C1517 VP.n115 VSUBS 1.36924f
C1518 VP.n116 VSUBS 0.024422f
C1519 VP.n117 VSUBS 0.022127f
C1520 VP.n118 VSUBS 0.022127f
C1521 VP.n119 VSUBS 0.022127f
C1522 VP.n120 VSUBS 0.041032f
C1523 VP.n121 VSUBS 0.043512f
C1524 VP.n122 VSUBS 0.017899f
C1525 VP.n123 VSUBS 0.022127f
C1526 VP.n124 VSUBS 0.022127f
C1527 VP.n125 VSUBS 0.022127f
C1528 VP.n126 VSUBS 0.041032f
C1529 VP.n127 VSUBS 0.041032f
C1530 VP.n128 VSUBS 0.023612f
C1531 VP.n129 VSUBS 0.035707f
C1532 VP.n130 VSUBS 0.067886f
.ends

