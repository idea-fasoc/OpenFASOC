* NGSPICE file created from diff_pair_sample_1091.ext - technology: sky130A

.subckt diff_pair_sample_1091 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t11 w_n4394_n2506# sky130_fd_pr__pfet_01v8 ad=2.9991 pd=16.16 as=1.26885 ps=8.02 w=7.69 l=3.95
X1 B.t11 B.t9 B.t10 w_n4394_n2506# sky130_fd_pr__pfet_01v8 ad=2.9991 pd=16.16 as=0 ps=0 w=7.69 l=3.95
X2 VDD1.t5 VP.t0 VTAIL.t2 w_n4394_n2506# sky130_fd_pr__pfet_01v8 ad=2.9991 pd=16.16 as=1.26885 ps=8.02 w=7.69 l=3.95
X3 VDD1.t4 VP.t1 VTAIL.t3 w_n4394_n2506# sky130_fd_pr__pfet_01v8 ad=1.26885 pd=8.02 as=2.9991 ps=16.16 w=7.69 l=3.95
X4 VTAIL.t7 VN.t1 VDD2.t4 w_n4394_n2506# sky130_fd_pr__pfet_01v8 ad=1.26885 pd=8.02 as=1.26885 ps=8.02 w=7.69 l=3.95
X5 VDD2.t3 VN.t2 VTAIL.t6 w_n4394_n2506# sky130_fd_pr__pfet_01v8 ad=1.26885 pd=8.02 as=2.9991 ps=16.16 w=7.69 l=3.95
X6 B.t8 B.t6 B.t7 w_n4394_n2506# sky130_fd_pr__pfet_01v8 ad=2.9991 pd=16.16 as=0 ps=0 w=7.69 l=3.95
X7 VTAIL.t0 VP.t2 VDD1.t3 w_n4394_n2506# sky130_fd_pr__pfet_01v8 ad=1.26885 pd=8.02 as=1.26885 ps=8.02 w=7.69 l=3.95
X8 VTAIL.t5 VP.t3 VDD1.t2 w_n4394_n2506# sky130_fd_pr__pfet_01v8 ad=1.26885 pd=8.02 as=1.26885 ps=8.02 w=7.69 l=3.95
X9 VDD2.t2 VN.t3 VTAIL.t8 w_n4394_n2506# sky130_fd_pr__pfet_01v8 ad=2.9991 pd=16.16 as=1.26885 ps=8.02 w=7.69 l=3.95
X10 VDD2.t1 VN.t4 VTAIL.t9 w_n4394_n2506# sky130_fd_pr__pfet_01v8 ad=1.26885 pd=8.02 as=2.9991 ps=16.16 w=7.69 l=3.95
X11 VDD1.t1 VP.t4 VTAIL.t4 w_n4394_n2506# sky130_fd_pr__pfet_01v8 ad=2.9991 pd=16.16 as=1.26885 ps=8.02 w=7.69 l=3.95
X12 B.t5 B.t3 B.t4 w_n4394_n2506# sky130_fd_pr__pfet_01v8 ad=2.9991 pd=16.16 as=0 ps=0 w=7.69 l=3.95
X13 VTAIL.t10 VN.t5 VDD2.t0 w_n4394_n2506# sky130_fd_pr__pfet_01v8 ad=1.26885 pd=8.02 as=1.26885 ps=8.02 w=7.69 l=3.95
X14 VDD1.t0 VP.t5 VTAIL.t1 w_n4394_n2506# sky130_fd_pr__pfet_01v8 ad=1.26885 pd=8.02 as=2.9991 ps=16.16 w=7.69 l=3.95
X15 B.t2 B.t0 B.t1 w_n4394_n2506# sky130_fd_pr__pfet_01v8 ad=2.9991 pd=16.16 as=0 ps=0 w=7.69 l=3.95
R0 VN.n42 VN.n41 161.3
R1 VN.n40 VN.n23 161.3
R2 VN.n39 VN.n38 161.3
R3 VN.n37 VN.n24 161.3
R4 VN.n36 VN.n35 161.3
R5 VN.n34 VN.n25 161.3
R6 VN.n33 VN.n32 161.3
R7 VN.n31 VN.n26 161.3
R8 VN.n30 VN.n29 161.3
R9 VN.n20 VN.n19 161.3
R10 VN.n18 VN.n1 161.3
R11 VN.n17 VN.n16 161.3
R12 VN.n15 VN.n2 161.3
R13 VN.n14 VN.n13 161.3
R14 VN.n12 VN.n3 161.3
R15 VN.n11 VN.n10 161.3
R16 VN.n9 VN.n4 161.3
R17 VN.n8 VN.n7 161.3
R18 VN.n21 VN.n0 88.5994
R19 VN.n43 VN.n22 88.5994
R20 VN.n27 VN.t2 79.3417
R21 VN.n5 VN.t0 79.3417
R22 VN.n6 VN.n5 62.9319
R23 VN.n28 VN.n27 62.9319
R24 VN.n13 VN.n12 51.1773
R25 VN.n35 VN.n34 51.1773
R26 VN VN.n43 50.9374
R27 VN.n6 VN.t1 46.9192
R28 VN.n0 VN.t4 46.9192
R29 VN.n28 VN.t5 46.9192
R30 VN.n22 VN.t3 46.9192
R31 VN.n13 VN.n2 29.8095
R32 VN.n35 VN.n24 29.8095
R33 VN.n7 VN.n4 24.4675
R34 VN.n11 VN.n4 24.4675
R35 VN.n12 VN.n11 24.4675
R36 VN.n17 VN.n2 24.4675
R37 VN.n18 VN.n17 24.4675
R38 VN.n19 VN.n18 24.4675
R39 VN.n34 VN.n33 24.4675
R40 VN.n33 VN.n26 24.4675
R41 VN.n29 VN.n26 24.4675
R42 VN.n41 VN.n40 24.4675
R43 VN.n40 VN.n39 24.4675
R44 VN.n39 VN.n24 24.4675
R45 VN.n7 VN.n6 12.234
R46 VN.n29 VN.n28 12.234
R47 VN.n30 VN.n27 2.50011
R48 VN.n8 VN.n5 2.50011
R49 VN.n19 VN.n0 1.46852
R50 VN.n41 VN.n22 1.46852
R51 VN.n43 VN.n42 0.354971
R52 VN.n21 VN.n20 0.354971
R53 VN VN.n21 0.26696
R54 VN.n42 VN.n23 0.189894
R55 VN.n38 VN.n23 0.189894
R56 VN.n38 VN.n37 0.189894
R57 VN.n37 VN.n36 0.189894
R58 VN.n36 VN.n25 0.189894
R59 VN.n32 VN.n25 0.189894
R60 VN.n32 VN.n31 0.189894
R61 VN.n31 VN.n30 0.189894
R62 VN.n9 VN.n8 0.189894
R63 VN.n10 VN.n9 0.189894
R64 VN.n10 VN.n3 0.189894
R65 VN.n14 VN.n3 0.189894
R66 VN.n15 VN.n14 0.189894
R67 VN.n16 VN.n15 0.189894
R68 VN.n16 VN.n1 0.189894
R69 VN.n20 VN.n1 0.189894
R70 VTAIL.n10 VTAIL.t1 69.3969
R71 VTAIL.n7 VTAIL.t6 69.3968
R72 VTAIL.n11 VTAIL.t9 69.3967
R73 VTAIL.n2 VTAIL.t3 69.3967
R74 VTAIL.n9 VTAIL.n8 65.17
R75 VTAIL.n6 VTAIL.n5 65.17
R76 VTAIL.n1 VTAIL.n0 65.1699
R77 VTAIL.n4 VTAIL.n3 65.1699
R78 VTAIL.n6 VTAIL.n4 26.3755
R79 VTAIL.n11 VTAIL.n10 22.6858
R80 VTAIL.n0 VTAIL.t11 4.22742
R81 VTAIL.n0 VTAIL.t7 4.22742
R82 VTAIL.n3 VTAIL.t4 4.22742
R83 VTAIL.n3 VTAIL.t5 4.22742
R84 VTAIL.n8 VTAIL.t2 4.22742
R85 VTAIL.n8 VTAIL.t0 4.22742
R86 VTAIL.n5 VTAIL.t8 4.22742
R87 VTAIL.n5 VTAIL.t10 4.22742
R88 VTAIL.n7 VTAIL.n6 3.69016
R89 VTAIL.n10 VTAIL.n9 3.69016
R90 VTAIL.n4 VTAIL.n2 3.69016
R91 VTAIL VTAIL.n11 2.70955
R92 VTAIL.n9 VTAIL.n7 2.31516
R93 VTAIL.n2 VTAIL.n1 2.31516
R94 VTAIL VTAIL.n1 0.981103
R95 VDD2.n1 VDD2.t5 88.7874
R96 VDD2.n2 VDD2.t2 86.0756
R97 VDD2.n1 VDD2.n0 82.7158
R98 VDD2 VDD2.n3 82.713
R99 VDD2.n2 VDD2.n1 42.336
R100 VDD2.n3 VDD2.t0 4.22742
R101 VDD2.n3 VDD2.t3 4.22742
R102 VDD2.n0 VDD2.t4 4.22742
R103 VDD2.n0 VDD2.t1 4.22742
R104 VDD2 VDD2.n2 2.82593
R105 B.n381 B.n128 585
R106 B.n380 B.n379 585
R107 B.n378 B.n129 585
R108 B.n377 B.n376 585
R109 B.n375 B.n130 585
R110 B.n374 B.n373 585
R111 B.n372 B.n131 585
R112 B.n371 B.n370 585
R113 B.n369 B.n132 585
R114 B.n368 B.n367 585
R115 B.n366 B.n133 585
R116 B.n365 B.n364 585
R117 B.n363 B.n134 585
R118 B.n362 B.n361 585
R119 B.n360 B.n135 585
R120 B.n359 B.n358 585
R121 B.n357 B.n136 585
R122 B.n356 B.n355 585
R123 B.n354 B.n137 585
R124 B.n353 B.n352 585
R125 B.n351 B.n138 585
R126 B.n350 B.n349 585
R127 B.n348 B.n139 585
R128 B.n347 B.n346 585
R129 B.n345 B.n140 585
R130 B.n344 B.n343 585
R131 B.n342 B.n141 585
R132 B.n341 B.n340 585
R133 B.n339 B.n142 585
R134 B.n338 B.n337 585
R135 B.n333 B.n143 585
R136 B.n332 B.n331 585
R137 B.n330 B.n144 585
R138 B.n329 B.n328 585
R139 B.n327 B.n145 585
R140 B.n326 B.n325 585
R141 B.n324 B.n146 585
R142 B.n323 B.n322 585
R143 B.n320 B.n147 585
R144 B.n319 B.n318 585
R145 B.n317 B.n150 585
R146 B.n316 B.n315 585
R147 B.n314 B.n151 585
R148 B.n313 B.n312 585
R149 B.n311 B.n152 585
R150 B.n310 B.n309 585
R151 B.n308 B.n153 585
R152 B.n307 B.n306 585
R153 B.n305 B.n154 585
R154 B.n304 B.n303 585
R155 B.n302 B.n155 585
R156 B.n301 B.n300 585
R157 B.n299 B.n156 585
R158 B.n298 B.n297 585
R159 B.n296 B.n157 585
R160 B.n295 B.n294 585
R161 B.n293 B.n158 585
R162 B.n292 B.n291 585
R163 B.n290 B.n159 585
R164 B.n289 B.n288 585
R165 B.n287 B.n160 585
R166 B.n286 B.n285 585
R167 B.n284 B.n161 585
R168 B.n283 B.n282 585
R169 B.n281 B.n162 585
R170 B.n280 B.n279 585
R171 B.n278 B.n163 585
R172 B.n383 B.n382 585
R173 B.n384 B.n127 585
R174 B.n386 B.n385 585
R175 B.n387 B.n126 585
R176 B.n389 B.n388 585
R177 B.n390 B.n125 585
R178 B.n392 B.n391 585
R179 B.n393 B.n124 585
R180 B.n395 B.n394 585
R181 B.n396 B.n123 585
R182 B.n398 B.n397 585
R183 B.n399 B.n122 585
R184 B.n401 B.n400 585
R185 B.n402 B.n121 585
R186 B.n404 B.n403 585
R187 B.n405 B.n120 585
R188 B.n407 B.n406 585
R189 B.n408 B.n119 585
R190 B.n410 B.n409 585
R191 B.n411 B.n118 585
R192 B.n413 B.n412 585
R193 B.n414 B.n117 585
R194 B.n416 B.n415 585
R195 B.n417 B.n116 585
R196 B.n419 B.n418 585
R197 B.n420 B.n115 585
R198 B.n422 B.n421 585
R199 B.n423 B.n114 585
R200 B.n425 B.n424 585
R201 B.n426 B.n113 585
R202 B.n428 B.n427 585
R203 B.n429 B.n112 585
R204 B.n431 B.n430 585
R205 B.n432 B.n111 585
R206 B.n434 B.n433 585
R207 B.n435 B.n110 585
R208 B.n437 B.n436 585
R209 B.n438 B.n109 585
R210 B.n440 B.n439 585
R211 B.n441 B.n108 585
R212 B.n443 B.n442 585
R213 B.n444 B.n107 585
R214 B.n446 B.n445 585
R215 B.n447 B.n106 585
R216 B.n449 B.n448 585
R217 B.n450 B.n105 585
R218 B.n452 B.n451 585
R219 B.n453 B.n104 585
R220 B.n455 B.n454 585
R221 B.n456 B.n103 585
R222 B.n458 B.n457 585
R223 B.n459 B.n102 585
R224 B.n461 B.n460 585
R225 B.n462 B.n101 585
R226 B.n464 B.n463 585
R227 B.n465 B.n100 585
R228 B.n467 B.n466 585
R229 B.n468 B.n99 585
R230 B.n470 B.n469 585
R231 B.n471 B.n98 585
R232 B.n473 B.n472 585
R233 B.n474 B.n97 585
R234 B.n476 B.n475 585
R235 B.n477 B.n96 585
R236 B.n479 B.n478 585
R237 B.n480 B.n95 585
R238 B.n482 B.n481 585
R239 B.n483 B.n94 585
R240 B.n485 B.n484 585
R241 B.n486 B.n93 585
R242 B.n488 B.n487 585
R243 B.n489 B.n92 585
R244 B.n491 B.n490 585
R245 B.n492 B.n91 585
R246 B.n494 B.n493 585
R247 B.n495 B.n90 585
R248 B.n497 B.n496 585
R249 B.n498 B.n89 585
R250 B.n500 B.n499 585
R251 B.n501 B.n88 585
R252 B.n503 B.n502 585
R253 B.n504 B.n87 585
R254 B.n506 B.n505 585
R255 B.n507 B.n86 585
R256 B.n509 B.n508 585
R257 B.n510 B.n85 585
R258 B.n512 B.n511 585
R259 B.n513 B.n84 585
R260 B.n515 B.n514 585
R261 B.n516 B.n83 585
R262 B.n518 B.n517 585
R263 B.n519 B.n82 585
R264 B.n521 B.n520 585
R265 B.n522 B.n81 585
R266 B.n524 B.n523 585
R267 B.n525 B.n80 585
R268 B.n527 B.n526 585
R269 B.n528 B.n79 585
R270 B.n530 B.n529 585
R271 B.n531 B.n78 585
R272 B.n533 B.n532 585
R273 B.n534 B.n77 585
R274 B.n536 B.n535 585
R275 B.n537 B.n76 585
R276 B.n539 B.n538 585
R277 B.n540 B.n75 585
R278 B.n542 B.n541 585
R279 B.n543 B.n74 585
R280 B.n545 B.n544 585
R281 B.n546 B.n73 585
R282 B.n548 B.n547 585
R283 B.n549 B.n72 585
R284 B.n551 B.n550 585
R285 B.n552 B.n71 585
R286 B.n554 B.n553 585
R287 B.n555 B.n70 585
R288 B.n557 B.n556 585
R289 B.n558 B.n69 585
R290 B.n660 B.n31 585
R291 B.n659 B.n658 585
R292 B.n657 B.n32 585
R293 B.n656 B.n655 585
R294 B.n654 B.n33 585
R295 B.n653 B.n652 585
R296 B.n651 B.n34 585
R297 B.n650 B.n649 585
R298 B.n648 B.n35 585
R299 B.n647 B.n646 585
R300 B.n645 B.n36 585
R301 B.n644 B.n643 585
R302 B.n642 B.n37 585
R303 B.n641 B.n640 585
R304 B.n639 B.n38 585
R305 B.n638 B.n637 585
R306 B.n636 B.n39 585
R307 B.n635 B.n634 585
R308 B.n633 B.n40 585
R309 B.n632 B.n631 585
R310 B.n630 B.n41 585
R311 B.n629 B.n628 585
R312 B.n627 B.n42 585
R313 B.n626 B.n625 585
R314 B.n624 B.n43 585
R315 B.n623 B.n622 585
R316 B.n621 B.n44 585
R317 B.n620 B.n619 585
R318 B.n618 B.n45 585
R319 B.n616 B.n615 585
R320 B.n614 B.n48 585
R321 B.n613 B.n612 585
R322 B.n611 B.n49 585
R323 B.n610 B.n609 585
R324 B.n608 B.n50 585
R325 B.n607 B.n606 585
R326 B.n605 B.n51 585
R327 B.n604 B.n603 585
R328 B.n602 B.n601 585
R329 B.n600 B.n55 585
R330 B.n599 B.n598 585
R331 B.n597 B.n56 585
R332 B.n596 B.n595 585
R333 B.n594 B.n57 585
R334 B.n593 B.n592 585
R335 B.n591 B.n58 585
R336 B.n590 B.n589 585
R337 B.n588 B.n59 585
R338 B.n587 B.n586 585
R339 B.n585 B.n60 585
R340 B.n584 B.n583 585
R341 B.n582 B.n61 585
R342 B.n581 B.n580 585
R343 B.n579 B.n62 585
R344 B.n578 B.n577 585
R345 B.n576 B.n63 585
R346 B.n575 B.n574 585
R347 B.n573 B.n64 585
R348 B.n572 B.n571 585
R349 B.n570 B.n65 585
R350 B.n569 B.n568 585
R351 B.n567 B.n66 585
R352 B.n566 B.n565 585
R353 B.n564 B.n67 585
R354 B.n563 B.n562 585
R355 B.n561 B.n68 585
R356 B.n560 B.n559 585
R357 B.n662 B.n661 585
R358 B.n663 B.n30 585
R359 B.n665 B.n664 585
R360 B.n666 B.n29 585
R361 B.n668 B.n667 585
R362 B.n669 B.n28 585
R363 B.n671 B.n670 585
R364 B.n672 B.n27 585
R365 B.n674 B.n673 585
R366 B.n675 B.n26 585
R367 B.n677 B.n676 585
R368 B.n678 B.n25 585
R369 B.n680 B.n679 585
R370 B.n681 B.n24 585
R371 B.n683 B.n682 585
R372 B.n684 B.n23 585
R373 B.n686 B.n685 585
R374 B.n687 B.n22 585
R375 B.n689 B.n688 585
R376 B.n690 B.n21 585
R377 B.n692 B.n691 585
R378 B.n693 B.n20 585
R379 B.n695 B.n694 585
R380 B.n696 B.n19 585
R381 B.n698 B.n697 585
R382 B.n699 B.n18 585
R383 B.n701 B.n700 585
R384 B.n702 B.n17 585
R385 B.n704 B.n703 585
R386 B.n705 B.n16 585
R387 B.n707 B.n706 585
R388 B.n708 B.n15 585
R389 B.n710 B.n709 585
R390 B.n711 B.n14 585
R391 B.n713 B.n712 585
R392 B.n714 B.n13 585
R393 B.n716 B.n715 585
R394 B.n717 B.n12 585
R395 B.n719 B.n718 585
R396 B.n720 B.n11 585
R397 B.n722 B.n721 585
R398 B.n723 B.n10 585
R399 B.n725 B.n724 585
R400 B.n726 B.n9 585
R401 B.n728 B.n727 585
R402 B.n729 B.n8 585
R403 B.n731 B.n730 585
R404 B.n732 B.n7 585
R405 B.n734 B.n733 585
R406 B.n735 B.n6 585
R407 B.n737 B.n736 585
R408 B.n738 B.n5 585
R409 B.n740 B.n739 585
R410 B.n741 B.n4 585
R411 B.n743 B.n742 585
R412 B.n744 B.n3 585
R413 B.n746 B.n745 585
R414 B.n747 B.n0 585
R415 B.n2 B.n1 585
R416 B.n193 B.n192 585
R417 B.n194 B.n191 585
R418 B.n196 B.n195 585
R419 B.n197 B.n190 585
R420 B.n199 B.n198 585
R421 B.n200 B.n189 585
R422 B.n202 B.n201 585
R423 B.n203 B.n188 585
R424 B.n205 B.n204 585
R425 B.n206 B.n187 585
R426 B.n208 B.n207 585
R427 B.n209 B.n186 585
R428 B.n211 B.n210 585
R429 B.n212 B.n185 585
R430 B.n214 B.n213 585
R431 B.n215 B.n184 585
R432 B.n217 B.n216 585
R433 B.n218 B.n183 585
R434 B.n220 B.n219 585
R435 B.n221 B.n182 585
R436 B.n223 B.n222 585
R437 B.n224 B.n181 585
R438 B.n226 B.n225 585
R439 B.n227 B.n180 585
R440 B.n229 B.n228 585
R441 B.n230 B.n179 585
R442 B.n232 B.n231 585
R443 B.n233 B.n178 585
R444 B.n235 B.n234 585
R445 B.n236 B.n177 585
R446 B.n238 B.n237 585
R447 B.n239 B.n176 585
R448 B.n241 B.n240 585
R449 B.n242 B.n175 585
R450 B.n244 B.n243 585
R451 B.n245 B.n174 585
R452 B.n247 B.n246 585
R453 B.n248 B.n173 585
R454 B.n250 B.n249 585
R455 B.n251 B.n172 585
R456 B.n253 B.n252 585
R457 B.n254 B.n171 585
R458 B.n256 B.n255 585
R459 B.n257 B.n170 585
R460 B.n259 B.n258 585
R461 B.n260 B.n169 585
R462 B.n262 B.n261 585
R463 B.n263 B.n168 585
R464 B.n265 B.n264 585
R465 B.n266 B.n167 585
R466 B.n268 B.n267 585
R467 B.n269 B.n166 585
R468 B.n271 B.n270 585
R469 B.n272 B.n165 585
R470 B.n274 B.n273 585
R471 B.n275 B.n164 585
R472 B.n277 B.n276 585
R473 B.n276 B.n163 530.939
R474 B.n382 B.n381 530.939
R475 B.n560 B.n69 530.939
R476 B.n662 B.n31 530.939
R477 B.n334 B.t0 257.053
R478 B.n52 B.t9 257.053
R479 B.n148 B.t3 256.815
R480 B.n46 B.t6 256.815
R481 B.n749 B.n748 256.663
R482 B.n748 B.n747 235.042
R483 B.n748 B.n2 235.042
R484 B.n334 B.t1 196.207
R485 B.n52 B.t11 196.207
R486 B.n148 B.t4 196.198
R487 B.n46 B.t8 196.198
R488 B.n280 B.n163 163.367
R489 B.n281 B.n280 163.367
R490 B.n282 B.n281 163.367
R491 B.n282 B.n161 163.367
R492 B.n286 B.n161 163.367
R493 B.n287 B.n286 163.367
R494 B.n288 B.n287 163.367
R495 B.n288 B.n159 163.367
R496 B.n292 B.n159 163.367
R497 B.n293 B.n292 163.367
R498 B.n294 B.n293 163.367
R499 B.n294 B.n157 163.367
R500 B.n298 B.n157 163.367
R501 B.n299 B.n298 163.367
R502 B.n300 B.n299 163.367
R503 B.n300 B.n155 163.367
R504 B.n304 B.n155 163.367
R505 B.n305 B.n304 163.367
R506 B.n306 B.n305 163.367
R507 B.n306 B.n153 163.367
R508 B.n310 B.n153 163.367
R509 B.n311 B.n310 163.367
R510 B.n312 B.n311 163.367
R511 B.n312 B.n151 163.367
R512 B.n316 B.n151 163.367
R513 B.n317 B.n316 163.367
R514 B.n318 B.n317 163.367
R515 B.n318 B.n147 163.367
R516 B.n323 B.n147 163.367
R517 B.n324 B.n323 163.367
R518 B.n325 B.n324 163.367
R519 B.n325 B.n145 163.367
R520 B.n329 B.n145 163.367
R521 B.n330 B.n329 163.367
R522 B.n331 B.n330 163.367
R523 B.n331 B.n143 163.367
R524 B.n338 B.n143 163.367
R525 B.n339 B.n338 163.367
R526 B.n340 B.n339 163.367
R527 B.n340 B.n141 163.367
R528 B.n344 B.n141 163.367
R529 B.n345 B.n344 163.367
R530 B.n346 B.n345 163.367
R531 B.n346 B.n139 163.367
R532 B.n350 B.n139 163.367
R533 B.n351 B.n350 163.367
R534 B.n352 B.n351 163.367
R535 B.n352 B.n137 163.367
R536 B.n356 B.n137 163.367
R537 B.n357 B.n356 163.367
R538 B.n358 B.n357 163.367
R539 B.n358 B.n135 163.367
R540 B.n362 B.n135 163.367
R541 B.n363 B.n362 163.367
R542 B.n364 B.n363 163.367
R543 B.n364 B.n133 163.367
R544 B.n368 B.n133 163.367
R545 B.n369 B.n368 163.367
R546 B.n370 B.n369 163.367
R547 B.n370 B.n131 163.367
R548 B.n374 B.n131 163.367
R549 B.n375 B.n374 163.367
R550 B.n376 B.n375 163.367
R551 B.n376 B.n129 163.367
R552 B.n380 B.n129 163.367
R553 B.n381 B.n380 163.367
R554 B.n556 B.n69 163.367
R555 B.n556 B.n555 163.367
R556 B.n555 B.n554 163.367
R557 B.n554 B.n71 163.367
R558 B.n550 B.n71 163.367
R559 B.n550 B.n549 163.367
R560 B.n549 B.n548 163.367
R561 B.n548 B.n73 163.367
R562 B.n544 B.n73 163.367
R563 B.n544 B.n543 163.367
R564 B.n543 B.n542 163.367
R565 B.n542 B.n75 163.367
R566 B.n538 B.n75 163.367
R567 B.n538 B.n537 163.367
R568 B.n537 B.n536 163.367
R569 B.n536 B.n77 163.367
R570 B.n532 B.n77 163.367
R571 B.n532 B.n531 163.367
R572 B.n531 B.n530 163.367
R573 B.n530 B.n79 163.367
R574 B.n526 B.n79 163.367
R575 B.n526 B.n525 163.367
R576 B.n525 B.n524 163.367
R577 B.n524 B.n81 163.367
R578 B.n520 B.n81 163.367
R579 B.n520 B.n519 163.367
R580 B.n519 B.n518 163.367
R581 B.n518 B.n83 163.367
R582 B.n514 B.n83 163.367
R583 B.n514 B.n513 163.367
R584 B.n513 B.n512 163.367
R585 B.n512 B.n85 163.367
R586 B.n508 B.n85 163.367
R587 B.n508 B.n507 163.367
R588 B.n507 B.n506 163.367
R589 B.n506 B.n87 163.367
R590 B.n502 B.n87 163.367
R591 B.n502 B.n501 163.367
R592 B.n501 B.n500 163.367
R593 B.n500 B.n89 163.367
R594 B.n496 B.n89 163.367
R595 B.n496 B.n495 163.367
R596 B.n495 B.n494 163.367
R597 B.n494 B.n91 163.367
R598 B.n490 B.n91 163.367
R599 B.n490 B.n489 163.367
R600 B.n489 B.n488 163.367
R601 B.n488 B.n93 163.367
R602 B.n484 B.n93 163.367
R603 B.n484 B.n483 163.367
R604 B.n483 B.n482 163.367
R605 B.n482 B.n95 163.367
R606 B.n478 B.n95 163.367
R607 B.n478 B.n477 163.367
R608 B.n477 B.n476 163.367
R609 B.n476 B.n97 163.367
R610 B.n472 B.n97 163.367
R611 B.n472 B.n471 163.367
R612 B.n471 B.n470 163.367
R613 B.n470 B.n99 163.367
R614 B.n466 B.n99 163.367
R615 B.n466 B.n465 163.367
R616 B.n465 B.n464 163.367
R617 B.n464 B.n101 163.367
R618 B.n460 B.n101 163.367
R619 B.n460 B.n459 163.367
R620 B.n459 B.n458 163.367
R621 B.n458 B.n103 163.367
R622 B.n454 B.n103 163.367
R623 B.n454 B.n453 163.367
R624 B.n453 B.n452 163.367
R625 B.n452 B.n105 163.367
R626 B.n448 B.n105 163.367
R627 B.n448 B.n447 163.367
R628 B.n447 B.n446 163.367
R629 B.n446 B.n107 163.367
R630 B.n442 B.n107 163.367
R631 B.n442 B.n441 163.367
R632 B.n441 B.n440 163.367
R633 B.n440 B.n109 163.367
R634 B.n436 B.n109 163.367
R635 B.n436 B.n435 163.367
R636 B.n435 B.n434 163.367
R637 B.n434 B.n111 163.367
R638 B.n430 B.n111 163.367
R639 B.n430 B.n429 163.367
R640 B.n429 B.n428 163.367
R641 B.n428 B.n113 163.367
R642 B.n424 B.n113 163.367
R643 B.n424 B.n423 163.367
R644 B.n423 B.n422 163.367
R645 B.n422 B.n115 163.367
R646 B.n418 B.n115 163.367
R647 B.n418 B.n417 163.367
R648 B.n417 B.n416 163.367
R649 B.n416 B.n117 163.367
R650 B.n412 B.n117 163.367
R651 B.n412 B.n411 163.367
R652 B.n411 B.n410 163.367
R653 B.n410 B.n119 163.367
R654 B.n406 B.n119 163.367
R655 B.n406 B.n405 163.367
R656 B.n405 B.n404 163.367
R657 B.n404 B.n121 163.367
R658 B.n400 B.n121 163.367
R659 B.n400 B.n399 163.367
R660 B.n399 B.n398 163.367
R661 B.n398 B.n123 163.367
R662 B.n394 B.n123 163.367
R663 B.n394 B.n393 163.367
R664 B.n393 B.n392 163.367
R665 B.n392 B.n125 163.367
R666 B.n388 B.n125 163.367
R667 B.n388 B.n387 163.367
R668 B.n387 B.n386 163.367
R669 B.n386 B.n127 163.367
R670 B.n382 B.n127 163.367
R671 B.n658 B.n31 163.367
R672 B.n658 B.n657 163.367
R673 B.n657 B.n656 163.367
R674 B.n656 B.n33 163.367
R675 B.n652 B.n33 163.367
R676 B.n652 B.n651 163.367
R677 B.n651 B.n650 163.367
R678 B.n650 B.n35 163.367
R679 B.n646 B.n35 163.367
R680 B.n646 B.n645 163.367
R681 B.n645 B.n644 163.367
R682 B.n644 B.n37 163.367
R683 B.n640 B.n37 163.367
R684 B.n640 B.n639 163.367
R685 B.n639 B.n638 163.367
R686 B.n638 B.n39 163.367
R687 B.n634 B.n39 163.367
R688 B.n634 B.n633 163.367
R689 B.n633 B.n632 163.367
R690 B.n632 B.n41 163.367
R691 B.n628 B.n41 163.367
R692 B.n628 B.n627 163.367
R693 B.n627 B.n626 163.367
R694 B.n626 B.n43 163.367
R695 B.n622 B.n43 163.367
R696 B.n622 B.n621 163.367
R697 B.n621 B.n620 163.367
R698 B.n620 B.n45 163.367
R699 B.n615 B.n45 163.367
R700 B.n615 B.n614 163.367
R701 B.n614 B.n613 163.367
R702 B.n613 B.n49 163.367
R703 B.n609 B.n49 163.367
R704 B.n609 B.n608 163.367
R705 B.n608 B.n607 163.367
R706 B.n607 B.n51 163.367
R707 B.n603 B.n51 163.367
R708 B.n603 B.n602 163.367
R709 B.n602 B.n55 163.367
R710 B.n598 B.n55 163.367
R711 B.n598 B.n597 163.367
R712 B.n597 B.n596 163.367
R713 B.n596 B.n57 163.367
R714 B.n592 B.n57 163.367
R715 B.n592 B.n591 163.367
R716 B.n591 B.n590 163.367
R717 B.n590 B.n59 163.367
R718 B.n586 B.n59 163.367
R719 B.n586 B.n585 163.367
R720 B.n585 B.n584 163.367
R721 B.n584 B.n61 163.367
R722 B.n580 B.n61 163.367
R723 B.n580 B.n579 163.367
R724 B.n579 B.n578 163.367
R725 B.n578 B.n63 163.367
R726 B.n574 B.n63 163.367
R727 B.n574 B.n573 163.367
R728 B.n573 B.n572 163.367
R729 B.n572 B.n65 163.367
R730 B.n568 B.n65 163.367
R731 B.n568 B.n567 163.367
R732 B.n567 B.n566 163.367
R733 B.n566 B.n67 163.367
R734 B.n562 B.n67 163.367
R735 B.n562 B.n561 163.367
R736 B.n561 B.n560 163.367
R737 B.n663 B.n662 163.367
R738 B.n664 B.n663 163.367
R739 B.n664 B.n29 163.367
R740 B.n668 B.n29 163.367
R741 B.n669 B.n668 163.367
R742 B.n670 B.n669 163.367
R743 B.n670 B.n27 163.367
R744 B.n674 B.n27 163.367
R745 B.n675 B.n674 163.367
R746 B.n676 B.n675 163.367
R747 B.n676 B.n25 163.367
R748 B.n680 B.n25 163.367
R749 B.n681 B.n680 163.367
R750 B.n682 B.n681 163.367
R751 B.n682 B.n23 163.367
R752 B.n686 B.n23 163.367
R753 B.n687 B.n686 163.367
R754 B.n688 B.n687 163.367
R755 B.n688 B.n21 163.367
R756 B.n692 B.n21 163.367
R757 B.n693 B.n692 163.367
R758 B.n694 B.n693 163.367
R759 B.n694 B.n19 163.367
R760 B.n698 B.n19 163.367
R761 B.n699 B.n698 163.367
R762 B.n700 B.n699 163.367
R763 B.n700 B.n17 163.367
R764 B.n704 B.n17 163.367
R765 B.n705 B.n704 163.367
R766 B.n706 B.n705 163.367
R767 B.n706 B.n15 163.367
R768 B.n710 B.n15 163.367
R769 B.n711 B.n710 163.367
R770 B.n712 B.n711 163.367
R771 B.n712 B.n13 163.367
R772 B.n716 B.n13 163.367
R773 B.n717 B.n716 163.367
R774 B.n718 B.n717 163.367
R775 B.n718 B.n11 163.367
R776 B.n722 B.n11 163.367
R777 B.n723 B.n722 163.367
R778 B.n724 B.n723 163.367
R779 B.n724 B.n9 163.367
R780 B.n728 B.n9 163.367
R781 B.n729 B.n728 163.367
R782 B.n730 B.n729 163.367
R783 B.n730 B.n7 163.367
R784 B.n734 B.n7 163.367
R785 B.n735 B.n734 163.367
R786 B.n736 B.n735 163.367
R787 B.n736 B.n5 163.367
R788 B.n740 B.n5 163.367
R789 B.n741 B.n740 163.367
R790 B.n742 B.n741 163.367
R791 B.n742 B.n3 163.367
R792 B.n746 B.n3 163.367
R793 B.n747 B.n746 163.367
R794 B.n192 B.n2 163.367
R795 B.n192 B.n191 163.367
R796 B.n196 B.n191 163.367
R797 B.n197 B.n196 163.367
R798 B.n198 B.n197 163.367
R799 B.n198 B.n189 163.367
R800 B.n202 B.n189 163.367
R801 B.n203 B.n202 163.367
R802 B.n204 B.n203 163.367
R803 B.n204 B.n187 163.367
R804 B.n208 B.n187 163.367
R805 B.n209 B.n208 163.367
R806 B.n210 B.n209 163.367
R807 B.n210 B.n185 163.367
R808 B.n214 B.n185 163.367
R809 B.n215 B.n214 163.367
R810 B.n216 B.n215 163.367
R811 B.n216 B.n183 163.367
R812 B.n220 B.n183 163.367
R813 B.n221 B.n220 163.367
R814 B.n222 B.n221 163.367
R815 B.n222 B.n181 163.367
R816 B.n226 B.n181 163.367
R817 B.n227 B.n226 163.367
R818 B.n228 B.n227 163.367
R819 B.n228 B.n179 163.367
R820 B.n232 B.n179 163.367
R821 B.n233 B.n232 163.367
R822 B.n234 B.n233 163.367
R823 B.n234 B.n177 163.367
R824 B.n238 B.n177 163.367
R825 B.n239 B.n238 163.367
R826 B.n240 B.n239 163.367
R827 B.n240 B.n175 163.367
R828 B.n244 B.n175 163.367
R829 B.n245 B.n244 163.367
R830 B.n246 B.n245 163.367
R831 B.n246 B.n173 163.367
R832 B.n250 B.n173 163.367
R833 B.n251 B.n250 163.367
R834 B.n252 B.n251 163.367
R835 B.n252 B.n171 163.367
R836 B.n256 B.n171 163.367
R837 B.n257 B.n256 163.367
R838 B.n258 B.n257 163.367
R839 B.n258 B.n169 163.367
R840 B.n262 B.n169 163.367
R841 B.n263 B.n262 163.367
R842 B.n264 B.n263 163.367
R843 B.n264 B.n167 163.367
R844 B.n268 B.n167 163.367
R845 B.n269 B.n268 163.367
R846 B.n270 B.n269 163.367
R847 B.n270 B.n165 163.367
R848 B.n274 B.n165 163.367
R849 B.n275 B.n274 163.367
R850 B.n276 B.n275 163.367
R851 B.n335 B.t2 113.201
R852 B.n53 B.t10 113.201
R853 B.n149 B.t5 113.192
R854 B.n47 B.t7 113.192
R855 B.n149 B.n148 83.0066
R856 B.n335 B.n334 83.0066
R857 B.n53 B.n52 83.0066
R858 B.n47 B.n46 83.0066
R859 B.n321 B.n149 59.5399
R860 B.n336 B.n335 59.5399
R861 B.n54 B.n53 59.5399
R862 B.n617 B.n47 59.5399
R863 B.n661 B.n660 34.4981
R864 B.n559 B.n558 34.4981
R865 B.n383 B.n128 34.4981
R866 B.n278 B.n277 34.4981
R867 B B.n749 18.0485
R868 B.n661 B.n30 10.6151
R869 B.n665 B.n30 10.6151
R870 B.n666 B.n665 10.6151
R871 B.n667 B.n666 10.6151
R872 B.n667 B.n28 10.6151
R873 B.n671 B.n28 10.6151
R874 B.n672 B.n671 10.6151
R875 B.n673 B.n672 10.6151
R876 B.n673 B.n26 10.6151
R877 B.n677 B.n26 10.6151
R878 B.n678 B.n677 10.6151
R879 B.n679 B.n678 10.6151
R880 B.n679 B.n24 10.6151
R881 B.n683 B.n24 10.6151
R882 B.n684 B.n683 10.6151
R883 B.n685 B.n684 10.6151
R884 B.n685 B.n22 10.6151
R885 B.n689 B.n22 10.6151
R886 B.n690 B.n689 10.6151
R887 B.n691 B.n690 10.6151
R888 B.n691 B.n20 10.6151
R889 B.n695 B.n20 10.6151
R890 B.n696 B.n695 10.6151
R891 B.n697 B.n696 10.6151
R892 B.n697 B.n18 10.6151
R893 B.n701 B.n18 10.6151
R894 B.n702 B.n701 10.6151
R895 B.n703 B.n702 10.6151
R896 B.n703 B.n16 10.6151
R897 B.n707 B.n16 10.6151
R898 B.n708 B.n707 10.6151
R899 B.n709 B.n708 10.6151
R900 B.n709 B.n14 10.6151
R901 B.n713 B.n14 10.6151
R902 B.n714 B.n713 10.6151
R903 B.n715 B.n714 10.6151
R904 B.n715 B.n12 10.6151
R905 B.n719 B.n12 10.6151
R906 B.n720 B.n719 10.6151
R907 B.n721 B.n720 10.6151
R908 B.n721 B.n10 10.6151
R909 B.n725 B.n10 10.6151
R910 B.n726 B.n725 10.6151
R911 B.n727 B.n726 10.6151
R912 B.n727 B.n8 10.6151
R913 B.n731 B.n8 10.6151
R914 B.n732 B.n731 10.6151
R915 B.n733 B.n732 10.6151
R916 B.n733 B.n6 10.6151
R917 B.n737 B.n6 10.6151
R918 B.n738 B.n737 10.6151
R919 B.n739 B.n738 10.6151
R920 B.n739 B.n4 10.6151
R921 B.n743 B.n4 10.6151
R922 B.n744 B.n743 10.6151
R923 B.n745 B.n744 10.6151
R924 B.n745 B.n0 10.6151
R925 B.n660 B.n659 10.6151
R926 B.n659 B.n32 10.6151
R927 B.n655 B.n32 10.6151
R928 B.n655 B.n654 10.6151
R929 B.n654 B.n653 10.6151
R930 B.n653 B.n34 10.6151
R931 B.n649 B.n34 10.6151
R932 B.n649 B.n648 10.6151
R933 B.n648 B.n647 10.6151
R934 B.n647 B.n36 10.6151
R935 B.n643 B.n36 10.6151
R936 B.n643 B.n642 10.6151
R937 B.n642 B.n641 10.6151
R938 B.n641 B.n38 10.6151
R939 B.n637 B.n38 10.6151
R940 B.n637 B.n636 10.6151
R941 B.n636 B.n635 10.6151
R942 B.n635 B.n40 10.6151
R943 B.n631 B.n40 10.6151
R944 B.n631 B.n630 10.6151
R945 B.n630 B.n629 10.6151
R946 B.n629 B.n42 10.6151
R947 B.n625 B.n42 10.6151
R948 B.n625 B.n624 10.6151
R949 B.n624 B.n623 10.6151
R950 B.n623 B.n44 10.6151
R951 B.n619 B.n44 10.6151
R952 B.n619 B.n618 10.6151
R953 B.n616 B.n48 10.6151
R954 B.n612 B.n48 10.6151
R955 B.n612 B.n611 10.6151
R956 B.n611 B.n610 10.6151
R957 B.n610 B.n50 10.6151
R958 B.n606 B.n50 10.6151
R959 B.n606 B.n605 10.6151
R960 B.n605 B.n604 10.6151
R961 B.n601 B.n600 10.6151
R962 B.n600 B.n599 10.6151
R963 B.n599 B.n56 10.6151
R964 B.n595 B.n56 10.6151
R965 B.n595 B.n594 10.6151
R966 B.n594 B.n593 10.6151
R967 B.n593 B.n58 10.6151
R968 B.n589 B.n58 10.6151
R969 B.n589 B.n588 10.6151
R970 B.n588 B.n587 10.6151
R971 B.n587 B.n60 10.6151
R972 B.n583 B.n60 10.6151
R973 B.n583 B.n582 10.6151
R974 B.n582 B.n581 10.6151
R975 B.n581 B.n62 10.6151
R976 B.n577 B.n62 10.6151
R977 B.n577 B.n576 10.6151
R978 B.n576 B.n575 10.6151
R979 B.n575 B.n64 10.6151
R980 B.n571 B.n64 10.6151
R981 B.n571 B.n570 10.6151
R982 B.n570 B.n569 10.6151
R983 B.n569 B.n66 10.6151
R984 B.n565 B.n66 10.6151
R985 B.n565 B.n564 10.6151
R986 B.n564 B.n563 10.6151
R987 B.n563 B.n68 10.6151
R988 B.n559 B.n68 10.6151
R989 B.n558 B.n557 10.6151
R990 B.n557 B.n70 10.6151
R991 B.n553 B.n70 10.6151
R992 B.n553 B.n552 10.6151
R993 B.n552 B.n551 10.6151
R994 B.n551 B.n72 10.6151
R995 B.n547 B.n72 10.6151
R996 B.n547 B.n546 10.6151
R997 B.n546 B.n545 10.6151
R998 B.n545 B.n74 10.6151
R999 B.n541 B.n74 10.6151
R1000 B.n541 B.n540 10.6151
R1001 B.n540 B.n539 10.6151
R1002 B.n539 B.n76 10.6151
R1003 B.n535 B.n76 10.6151
R1004 B.n535 B.n534 10.6151
R1005 B.n534 B.n533 10.6151
R1006 B.n533 B.n78 10.6151
R1007 B.n529 B.n78 10.6151
R1008 B.n529 B.n528 10.6151
R1009 B.n528 B.n527 10.6151
R1010 B.n527 B.n80 10.6151
R1011 B.n523 B.n80 10.6151
R1012 B.n523 B.n522 10.6151
R1013 B.n522 B.n521 10.6151
R1014 B.n521 B.n82 10.6151
R1015 B.n517 B.n82 10.6151
R1016 B.n517 B.n516 10.6151
R1017 B.n516 B.n515 10.6151
R1018 B.n515 B.n84 10.6151
R1019 B.n511 B.n84 10.6151
R1020 B.n511 B.n510 10.6151
R1021 B.n510 B.n509 10.6151
R1022 B.n509 B.n86 10.6151
R1023 B.n505 B.n86 10.6151
R1024 B.n505 B.n504 10.6151
R1025 B.n504 B.n503 10.6151
R1026 B.n503 B.n88 10.6151
R1027 B.n499 B.n88 10.6151
R1028 B.n499 B.n498 10.6151
R1029 B.n498 B.n497 10.6151
R1030 B.n497 B.n90 10.6151
R1031 B.n493 B.n90 10.6151
R1032 B.n493 B.n492 10.6151
R1033 B.n492 B.n491 10.6151
R1034 B.n491 B.n92 10.6151
R1035 B.n487 B.n92 10.6151
R1036 B.n487 B.n486 10.6151
R1037 B.n486 B.n485 10.6151
R1038 B.n485 B.n94 10.6151
R1039 B.n481 B.n94 10.6151
R1040 B.n481 B.n480 10.6151
R1041 B.n480 B.n479 10.6151
R1042 B.n479 B.n96 10.6151
R1043 B.n475 B.n96 10.6151
R1044 B.n475 B.n474 10.6151
R1045 B.n474 B.n473 10.6151
R1046 B.n473 B.n98 10.6151
R1047 B.n469 B.n98 10.6151
R1048 B.n469 B.n468 10.6151
R1049 B.n468 B.n467 10.6151
R1050 B.n467 B.n100 10.6151
R1051 B.n463 B.n100 10.6151
R1052 B.n463 B.n462 10.6151
R1053 B.n462 B.n461 10.6151
R1054 B.n461 B.n102 10.6151
R1055 B.n457 B.n102 10.6151
R1056 B.n457 B.n456 10.6151
R1057 B.n456 B.n455 10.6151
R1058 B.n455 B.n104 10.6151
R1059 B.n451 B.n104 10.6151
R1060 B.n451 B.n450 10.6151
R1061 B.n450 B.n449 10.6151
R1062 B.n449 B.n106 10.6151
R1063 B.n445 B.n106 10.6151
R1064 B.n445 B.n444 10.6151
R1065 B.n444 B.n443 10.6151
R1066 B.n443 B.n108 10.6151
R1067 B.n439 B.n108 10.6151
R1068 B.n439 B.n438 10.6151
R1069 B.n438 B.n437 10.6151
R1070 B.n437 B.n110 10.6151
R1071 B.n433 B.n110 10.6151
R1072 B.n433 B.n432 10.6151
R1073 B.n432 B.n431 10.6151
R1074 B.n431 B.n112 10.6151
R1075 B.n427 B.n112 10.6151
R1076 B.n427 B.n426 10.6151
R1077 B.n426 B.n425 10.6151
R1078 B.n425 B.n114 10.6151
R1079 B.n421 B.n114 10.6151
R1080 B.n421 B.n420 10.6151
R1081 B.n420 B.n419 10.6151
R1082 B.n419 B.n116 10.6151
R1083 B.n415 B.n116 10.6151
R1084 B.n415 B.n414 10.6151
R1085 B.n414 B.n413 10.6151
R1086 B.n413 B.n118 10.6151
R1087 B.n409 B.n118 10.6151
R1088 B.n409 B.n408 10.6151
R1089 B.n408 B.n407 10.6151
R1090 B.n407 B.n120 10.6151
R1091 B.n403 B.n120 10.6151
R1092 B.n403 B.n402 10.6151
R1093 B.n402 B.n401 10.6151
R1094 B.n401 B.n122 10.6151
R1095 B.n397 B.n122 10.6151
R1096 B.n397 B.n396 10.6151
R1097 B.n396 B.n395 10.6151
R1098 B.n395 B.n124 10.6151
R1099 B.n391 B.n124 10.6151
R1100 B.n391 B.n390 10.6151
R1101 B.n390 B.n389 10.6151
R1102 B.n389 B.n126 10.6151
R1103 B.n385 B.n126 10.6151
R1104 B.n385 B.n384 10.6151
R1105 B.n384 B.n383 10.6151
R1106 B.n193 B.n1 10.6151
R1107 B.n194 B.n193 10.6151
R1108 B.n195 B.n194 10.6151
R1109 B.n195 B.n190 10.6151
R1110 B.n199 B.n190 10.6151
R1111 B.n200 B.n199 10.6151
R1112 B.n201 B.n200 10.6151
R1113 B.n201 B.n188 10.6151
R1114 B.n205 B.n188 10.6151
R1115 B.n206 B.n205 10.6151
R1116 B.n207 B.n206 10.6151
R1117 B.n207 B.n186 10.6151
R1118 B.n211 B.n186 10.6151
R1119 B.n212 B.n211 10.6151
R1120 B.n213 B.n212 10.6151
R1121 B.n213 B.n184 10.6151
R1122 B.n217 B.n184 10.6151
R1123 B.n218 B.n217 10.6151
R1124 B.n219 B.n218 10.6151
R1125 B.n219 B.n182 10.6151
R1126 B.n223 B.n182 10.6151
R1127 B.n224 B.n223 10.6151
R1128 B.n225 B.n224 10.6151
R1129 B.n225 B.n180 10.6151
R1130 B.n229 B.n180 10.6151
R1131 B.n230 B.n229 10.6151
R1132 B.n231 B.n230 10.6151
R1133 B.n231 B.n178 10.6151
R1134 B.n235 B.n178 10.6151
R1135 B.n236 B.n235 10.6151
R1136 B.n237 B.n236 10.6151
R1137 B.n237 B.n176 10.6151
R1138 B.n241 B.n176 10.6151
R1139 B.n242 B.n241 10.6151
R1140 B.n243 B.n242 10.6151
R1141 B.n243 B.n174 10.6151
R1142 B.n247 B.n174 10.6151
R1143 B.n248 B.n247 10.6151
R1144 B.n249 B.n248 10.6151
R1145 B.n249 B.n172 10.6151
R1146 B.n253 B.n172 10.6151
R1147 B.n254 B.n253 10.6151
R1148 B.n255 B.n254 10.6151
R1149 B.n255 B.n170 10.6151
R1150 B.n259 B.n170 10.6151
R1151 B.n260 B.n259 10.6151
R1152 B.n261 B.n260 10.6151
R1153 B.n261 B.n168 10.6151
R1154 B.n265 B.n168 10.6151
R1155 B.n266 B.n265 10.6151
R1156 B.n267 B.n266 10.6151
R1157 B.n267 B.n166 10.6151
R1158 B.n271 B.n166 10.6151
R1159 B.n272 B.n271 10.6151
R1160 B.n273 B.n272 10.6151
R1161 B.n273 B.n164 10.6151
R1162 B.n277 B.n164 10.6151
R1163 B.n279 B.n278 10.6151
R1164 B.n279 B.n162 10.6151
R1165 B.n283 B.n162 10.6151
R1166 B.n284 B.n283 10.6151
R1167 B.n285 B.n284 10.6151
R1168 B.n285 B.n160 10.6151
R1169 B.n289 B.n160 10.6151
R1170 B.n290 B.n289 10.6151
R1171 B.n291 B.n290 10.6151
R1172 B.n291 B.n158 10.6151
R1173 B.n295 B.n158 10.6151
R1174 B.n296 B.n295 10.6151
R1175 B.n297 B.n296 10.6151
R1176 B.n297 B.n156 10.6151
R1177 B.n301 B.n156 10.6151
R1178 B.n302 B.n301 10.6151
R1179 B.n303 B.n302 10.6151
R1180 B.n303 B.n154 10.6151
R1181 B.n307 B.n154 10.6151
R1182 B.n308 B.n307 10.6151
R1183 B.n309 B.n308 10.6151
R1184 B.n309 B.n152 10.6151
R1185 B.n313 B.n152 10.6151
R1186 B.n314 B.n313 10.6151
R1187 B.n315 B.n314 10.6151
R1188 B.n315 B.n150 10.6151
R1189 B.n319 B.n150 10.6151
R1190 B.n320 B.n319 10.6151
R1191 B.n322 B.n146 10.6151
R1192 B.n326 B.n146 10.6151
R1193 B.n327 B.n326 10.6151
R1194 B.n328 B.n327 10.6151
R1195 B.n328 B.n144 10.6151
R1196 B.n332 B.n144 10.6151
R1197 B.n333 B.n332 10.6151
R1198 B.n337 B.n333 10.6151
R1199 B.n341 B.n142 10.6151
R1200 B.n342 B.n341 10.6151
R1201 B.n343 B.n342 10.6151
R1202 B.n343 B.n140 10.6151
R1203 B.n347 B.n140 10.6151
R1204 B.n348 B.n347 10.6151
R1205 B.n349 B.n348 10.6151
R1206 B.n349 B.n138 10.6151
R1207 B.n353 B.n138 10.6151
R1208 B.n354 B.n353 10.6151
R1209 B.n355 B.n354 10.6151
R1210 B.n355 B.n136 10.6151
R1211 B.n359 B.n136 10.6151
R1212 B.n360 B.n359 10.6151
R1213 B.n361 B.n360 10.6151
R1214 B.n361 B.n134 10.6151
R1215 B.n365 B.n134 10.6151
R1216 B.n366 B.n365 10.6151
R1217 B.n367 B.n366 10.6151
R1218 B.n367 B.n132 10.6151
R1219 B.n371 B.n132 10.6151
R1220 B.n372 B.n371 10.6151
R1221 B.n373 B.n372 10.6151
R1222 B.n373 B.n130 10.6151
R1223 B.n377 B.n130 10.6151
R1224 B.n378 B.n377 10.6151
R1225 B.n379 B.n378 10.6151
R1226 B.n379 B.n128 10.6151
R1227 B.n749 B.n0 8.11757
R1228 B.n749 B.n1 8.11757
R1229 B.n617 B.n616 6.4005
R1230 B.n604 B.n54 6.4005
R1231 B.n322 B.n321 6.4005
R1232 B.n337 B.n336 6.4005
R1233 B.n618 B.n617 4.21513
R1234 B.n601 B.n54 4.21513
R1235 B.n321 B.n320 4.21513
R1236 B.n336 B.n142 4.21513
R1237 VP.n18 VP.n17 161.3
R1238 VP.n19 VP.n14 161.3
R1239 VP.n21 VP.n20 161.3
R1240 VP.n22 VP.n13 161.3
R1241 VP.n24 VP.n23 161.3
R1242 VP.n25 VP.n12 161.3
R1243 VP.n27 VP.n26 161.3
R1244 VP.n28 VP.n11 161.3
R1245 VP.n30 VP.n29 161.3
R1246 VP.n61 VP.n60 161.3
R1247 VP.n59 VP.n1 161.3
R1248 VP.n58 VP.n57 161.3
R1249 VP.n56 VP.n2 161.3
R1250 VP.n55 VP.n54 161.3
R1251 VP.n53 VP.n3 161.3
R1252 VP.n52 VP.n51 161.3
R1253 VP.n50 VP.n4 161.3
R1254 VP.n49 VP.n48 161.3
R1255 VP.n46 VP.n5 161.3
R1256 VP.n45 VP.n44 161.3
R1257 VP.n43 VP.n6 161.3
R1258 VP.n42 VP.n41 161.3
R1259 VP.n40 VP.n7 161.3
R1260 VP.n39 VP.n38 161.3
R1261 VP.n37 VP.n8 161.3
R1262 VP.n36 VP.n35 161.3
R1263 VP.n34 VP.n9 161.3
R1264 VP.n33 VP.n32 88.5994
R1265 VP.n62 VP.n0 88.5994
R1266 VP.n31 VP.n10 88.5994
R1267 VP.n15 VP.t0 79.3416
R1268 VP.n16 VP.n15 62.9319
R1269 VP.n41 VP.n40 51.1773
R1270 VP.n54 VP.n53 51.1773
R1271 VP.n23 VP.n22 51.1773
R1272 VP.n32 VP.n31 50.7721
R1273 VP.n33 VP.t4 46.9192
R1274 VP.n47 VP.t3 46.9192
R1275 VP.n0 VP.t1 46.9192
R1276 VP.n10 VP.t5 46.9192
R1277 VP.n16 VP.t2 46.9192
R1278 VP.n40 VP.n39 29.8095
R1279 VP.n54 VP.n2 29.8095
R1280 VP.n23 VP.n12 29.8095
R1281 VP.n35 VP.n34 24.4675
R1282 VP.n35 VP.n8 24.4675
R1283 VP.n39 VP.n8 24.4675
R1284 VP.n41 VP.n6 24.4675
R1285 VP.n45 VP.n6 24.4675
R1286 VP.n46 VP.n45 24.4675
R1287 VP.n48 VP.n4 24.4675
R1288 VP.n52 VP.n4 24.4675
R1289 VP.n53 VP.n52 24.4675
R1290 VP.n58 VP.n2 24.4675
R1291 VP.n59 VP.n58 24.4675
R1292 VP.n60 VP.n59 24.4675
R1293 VP.n27 VP.n12 24.4675
R1294 VP.n28 VP.n27 24.4675
R1295 VP.n29 VP.n28 24.4675
R1296 VP.n17 VP.n14 24.4675
R1297 VP.n21 VP.n14 24.4675
R1298 VP.n22 VP.n21 24.4675
R1299 VP.n47 VP.n46 12.234
R1300 VP.n48 VP.n47 12.234
R1301 VP.n17 VP.n16 12.234
R1302 VP.n18 VP.n15 2.5001
R1303 VP.n34 VP.n33 1.46852
R1304 VP.n60 VP.n0 1.46852
R1305 VP.n29 VP.n10 1.46852
R1306 VP.n31 VP.n30 0.354971
R1307 VP.n32 VP.n9 0.354971
R1308 VP.n62 VP.n61 0.354971
R1309 VP VP.n62 0.26696
R1310 VP.n19 VP.n18 0.189894
R1311 VP.n20 VP.n19 0.189894
R1312 VP.n20 VP.n13 0.189894
R1313 VP.n24 VP.n13 0.189894
R1314 VP.n25 VP.n24 0.189894
R1315 VP.n26 VP.n25 0.189894
R1316 VP.n26 VP.n11 0.189894
R1317 VP.n30 VP.n11 0.189894
R1318 VP.n36 VP.n9 0.189894
R1319 VP.n37 VP.n36 0.189894
R1320 VP.n38 VP.n37 0.189894
R1321 VP.n38 VP.n7 0.189894
R1322 VP.n42 VP.n7 0.189894
R1323 VP.n43 VP.n42 0.189894
R1324 VP.n44 VP.n43 0.189894
R1325 VP.n44 VP.n5 0.189894
R1326 VP.n49 VP.n5 0.189894
R1327 VP.n50 VP.n49 0.189894
R1328 VP.n51 VP.n50 0.189894
R1329 VP.n51 VP.n3 0.189894
R1330 VP.n55 VP.n3 0.189894
R1331 VP.n56 VP.n55 0.189894
R1332 VP.n57 VP.n56 0.189894
R1333 VP.n57 VP.n1 0.189894
R1334 VP.n61 VP.n1 0.189894
R1335 VDD1 VDD1.t5 88.901
R1336 VDD1.n1 VDD1.t1 88.7874
R1337 VDD1.n1 VDD1.n0 82.7158
R1338 VDD1.n3 VDD1.n2 81.8488
R1339 VDD1.n3 VDD1.n1 44.7638
R1340 VDD1.n2 VDD1.t3 4.22742
R1341 VDD1.n2 VDD1.t0 4.22742
R1342 VDD1.n0 VDD1.t2 4.22742
R1343 VDD1.n0 VDD1.t4 4.22742
R1344 VDD1 VDD1.n3 0.864724
C0 B VDD1 2.094f
C1 VDD2 w_n4394_n2506# 2.45054f
C2 B VTAIL 3.15454f
C3 VN VDD2 4.75051f
C4 VP w_n4394_n2506# 9.15217f
C5 VDD2 VDD1 1.93352f
C6 VP VN 7.44021f
C7 VDD2 VTAIL 6.94493f
C8 VP VDD1 5.16798f
C9 B VDD2 2.20047f
C10 VN w_n4394_n2506# 8.58033f
C11 VP VTAIL 5.46285f
C12 VDD1 w_n4394_n2506# 2.3223f
C13 B VP 2.36901f
C14 VN VDD1 0.152606f
C15 VTAIL w_n4394_n2506# 2.50526f
C16 B w_n4394_n2506# 10.3501f
C17 VN VTAIL 5.44825f
C18 VP VDD2 0.572186f
C19 B VN 1.40745f
C20 VDD1 VTAIL 6.88336f
C21 VDD2 VSUBS 2.199848f
C22 VDD1 VSUBS 2.77874f
C23 VTAIL VSUBS 1.31493f
C24 VN VSUBS 7.14626f
C25 VP VSUBS 3.830885f
C26 B VSUBS 5.607995f
C27 w_n4394_n2506# VSUBS 0.136724p
C28 VDD1.t5 VSUBS 1.75215f
C29 VDD1.t1 VSUBS 1.75069f
C30 VDD1.t2 VSUBS 0.184715f
C31 VDD1.t4 VSUBS 0.184715f
C32 VDD1.n0 VSUBS 1.30953f
C33 VDD1.n1 VSUBS 4.67323f
C34 VDD1.t3 VSUBS 0.184715f
C35 VDD1.t0 VSUBS 0.184715f
C36 VDD1.n2 VSUBS 1.2991f
C37 VDD1.n3 VSUBS 3.73953f
C38 VP.t1 VSUBS 2.66835f
C39 VP.n0 VSUBS 1.08598f
C40 VP.n1 VSUBS 0.032796f
C41 VP.n2 VSUBS 0.065339f
C42 VP.n3 VSUBS 0.032796f
C43 VP.n4 VSUBS 0.061123f
C44 VP.n5 VSUBS 0.032796f
C45 VP.t3 VSUBS 2.66835f
C46 VP.n6 VSUBS 0.061123f
C47 VP.n7 VSUBS 0.032796f
C48 VP.n8 VSUBS 0.061123f
C49 VP.n9 VSUBS 0.052932f
C50 VP.t4 VSUBS 2.66835f
C51 VP.t5 VSUBS 2.66835f
C52 VP.n10 VSUBS 1.08598f
C53 VP.n11 VSUBS 0.032796f
C54 VP.n12 VSUBS 0.065339f
C55 VP.n13 VSUBS 0.032796f
C56 VP.n14 VSUBS 0.061123f
C57 VP.t0 VSUBS 3.16976f
C58 VP.n15 VSUBS 1.04018f
C59 VP.t2 VSUBS 2.66835f
C60 VP.n16 VSUBS 1.08024f
C61 VP.n17 VSUBS 0.046035f
C62 VP.n18 VSUBS 0.428878f
C63 VP.n19 VSUBS 0.032796f
C64 VP.n20 VSUBS 0.032796f
C65 VP.n21 VSUBS 0.061123f
C66 VP.n22 VSUBS 0.059545f
C67 VP.n23 VSUBS 0.03199f
C68 VP.n24 VSUBS 0.032796f
C69 VP.n25 VSUBS 0.032796f
C70 VP.n26 VSUBS 0.032796f
C71 VP.n27 VSUBS 0.061123f
C72 VP.n28 VSUBS 0.061123f
C73 VP.n29 VSUBS 0.032757f
C74 VP.n30 VSUBS 0.052932f
C75 VP.n31 VSUBS 1.93399f
C76 VP.n32 VSUBS 1.95721f
C77 VP.n33 VSUBS 1.08598f
C78 VP.n34 VSUBS 0.032757f
C79 VP.n35 VSUBS 0.061123f
C80 VP.n36 VSUBS 0.032796f
C81 VP.n37 VSUBS 0.032796f
C82 VP.n38 VSUBS 0.032796f
C83 VP.n39 VSUBS 0.065339f
C84 VP.n40 VSUBS 0.03199f
C85 VP.n41 VSUBS 0.059545f
C86 VP.n42 VSUBS 0.032796f
C87 VP.n43 VSUBS 0.032796f
C88 VP.n44 VSUBS 0.032796f
C89 VP.n45 VSUBS 0.061123f
C90 VP.n46 VSUBS 0.046035f
C91 VP.n47 VSUBS 0.960772f
C92 VP.n48 VSUBS 0.046035f
C93 VP.n49 VSUBS 0.032796f
C94 VP.n50 VSUBS 0.032796f
C95 VP.n51 VSUBS 0.032796f
C96 VP.n52 VSUBS 0.061123f
C97 VP.n53 VSUBS 0.059545f
C98 VP.n54 VSUBS 0.03199f
C99 VP.n55 VSUBS 0.032796f
C100 VP.n56 VSUBS 0.032796f
C101 VP.n57 VSUBS 0.032796f
C102 VP.n58 VSUBS 0.061123f
C103 VP.n59 VSUBS 0.061123f
C104 VP.n60 VSUBS 0.032757f
C105 VP.n61 VSUBS 0.052932f
C106 VP.n62 VSUBS 0.104901f
C107 B.n0 VSUBS 0.008874f
C108 B.n1 VSUBS 0.008874f
C109 B.n2 VSUBS 0.013124f
C110 B.n3 VSUBS 0.010057f
C111 B.n4 VSUBS 0.010057f
C112 B.n5 VSUBS 0.010057f
C113 B.n6 VSUBS 0.010057f
C114 B.n7 VSUBS 0.010057f
C115 B.n8 VSUBS 0.010057f
C116 B.n9 VSUBS 0.010057f
C117 B.n10 VSUBS 0.010057f
C118 B.n11 VSUBS 0.010057f
C119 B.n12 VSUBS 0.010057f
C120 B.n13 VSUBS 0.010057f
C121 B.n14 VSUBS 0.010057f
C122 B.n15 VSUBS 0.010057f
C123 B.n16 VSUBS 0.010057f
C124 B.n17 VSUBS 0.010057f
C125 B.n18 VSUBS 0.010057f
C126 B.n19 VSUBS 0.010057f
C127 B.n20 VSUBS 0.010057f
C128 B.n21 VSUBS 0.010057f
C129 B.n22 VSUBS 0.010057f
C130 B.n23 VSUBS 0.010057f
C131 B.n24 VSUBS 0.010057f
C132 B.n25 VSUBS 0.010057f
C133 B.n26 VSUBS 0.010057f
C134 B.n27 VSUBS 0.010057f
C135 B.n28 VSUBS 0.010057f
C136 B.n29 VSUBS 0.010057f
C137 B.n30 VSUBS 0.010057f
C138 B.n31 VSUBS 0.02469f
C139 B.n32 VSUBS 0.010057f
C140 B.n33 VSUBS 0.010057f
C141 B.n34 VSUBS 0.010057f
C142 B.n35 VSUBS 0.010057f
C143 B.n36 VSUBS 0.010057f
C144 B.n37 VSUBS 0.010057f
C145 B.n38 VSUBS 0.010057f
C146 B.n39 VSUBS 0.010057f
C147 B.n40 VSUBS 0.010057f
C148 B.n41 VSUBS 0.010057f
C149 B.n42 VSUBS 0.010057f
C150 B.n43 VSUBS 0.010057f
C151 B.n44 VSUBS 0.010057f
C152 B.n45 VSUBS 0.010057f
C153 B.t7 VSUBS 0.338688f
C154 B.t8 VSUBS 0.379398f
C155 B.t6 VSUBS 2.08146f
C156 B.n46 VSUBS 0.224234f
C157 B.n47 VSUBS 0.110569f
C158 B.n48 VSUBS 0.010057f
C159 B.n49 VSUBS 0.010057f
C160 B.n50 VSUBS 0.010057f
C161 B.n51 VSUBS 0.010057f
C162 B.t10 VSUBS 0.338685f
C163 B.t11 VSUBS 0.379395f
C164 B.t9 VSUBS 2.08159f
C165 B.n52 VSUBS 0.224107f
C166 B.n53 VSUBS 0.110572f
C167 B.n54 VSUBS 0.0233f
C168 B.n55 VSUBS 0.010057f
C169 B.n56 VSUBS 0.010057f
C170 B.n57 VSUBS 0.010057f
C171 B.n58 VSUBS 0.010057f
C172 B.n59 VSUBS 0.010057f
C173 B.n60 VSUBS 0.010057f
C174 B.n61 VSUBS 0.010057f
C175 B.n62 VSUBS 0.010057f
C176 B.n63 VSUBS 0.010057f
C177 B.n64 VSUBS 0.010057f
C178 B.n65 VSUBS 0.010057f
C179 B.n66 VSUBS 0.010057f
C180 B.n67 VSUBS 0.010057f
C181 B.n68 VSUBS 0.010057f
C182 B.n69 VSUBS 0.024114f
C183 B.n70 VSUBS 0.010057f
C184 B.n71 VSUBS 0.010057f
C185 B.n72 VSUBS 0.010057f
C186 B.n73 VSUBS 0.010057f
C187 B.n74 VSUBS 0.010057f
C188 B.n75 VSUBS 0.010057f
C189 B.n76 VSUBS 0.010057f
C190 B.n77 VSUBS 0.010057f
C191 B.n78 VSUBS 0.010057f
C192 B.n79 VSUBS 0.010057f
C193 B.n80 VSUBS 0.010057f
C194 B.n81 VSUBS 0.010057f
C195 B.n82 VSUBS 0.010057f
C196 B.n83 VSUBS 0.010057f
C197 B.n84 VSUBS 0.010057f
C198 B.n85 VSUBS 0.010057f
C199 B.n86 VSUBS 0.010057f
C200 B.n87 VSUBS 0.010057f
C201 B.n88 VSUBS 0.010057f
C202 B.n89 VSUBS 0.010057f
C203 B.n90 VSUBS 0.010057f
C204 B.n91 VSUBS 0.010057f
C205 B.n92 VSUBS 0.010057f
C206 B.n93 VSUBS 0.010057f
C207 B.n94 VSUBS 0.010057f
C208 B.n95 VSUBS 0.010057f
C209 B.n96 VSUBS 0.010057f
C210 B.n97 VSUBS 0.010057f
C211 B.n98 VSUBS 0.010057f
C212 B.n99 VSUBS 0.010057f
C213 B.n100 VSUBS 0.010057f
C214 B.n101 VSUBS 0.010057f
C215 B.n102 VSUBS 0.010057f
C216 B.n103 VSUBS 0.010057f
C217 B.n104 VSUBS 0.010057f
C218 B.n105 VSUBS 0.010057f
C219 B.n106 VSUBS 0.010057f
C220 B.n107 VSUBS 0.010057f
C221 B.n108 VSUBS 0.010057f
C222 B.n109 VSUBS 0.010057f
C223 B.n110 VSUBS 0.010057f
C224 B.n111 VSUBS 0.010057f
C225 B.n112 VSUBS 0.010057f
C226 B.n113 VSUBS 0.010057f
C227 B.n114 VSUBS 0.010057f
C228 B.n115 VSUBS 0.010057f
C229 B.n116 VSUBS 0.010057f
C230 B.n117 VSUBS 0.010057f
C231 B.n118 VSUBS 0.010057f
C232 B.n119 VSUBS 0.010057f
C233 B.n120 VSUBS 0.010057f
C234 B.n121 VSUBS 0.010057f
C235 B.n122 VSUBS 0.010057f
C236 B.n123 VSUBS 0.010057f
C237 B.n124 VSUBS 0.010057f
C238 B.n125 VSUBS 0.010057f
C239 B.n126 VSUBS 0.010057f
C240 B.n127 VSUBS 0.010057f
C241 B.n128 VSUBS 0.023566f
C242 B.n129 VSUBS 0.010057f
C243 B.n130 VSUBS 0.010057f
C244 B.n131 VSUBS 0.010057f
C245 B.n132 VSUBS 0.010057f
C246 B.n133 VSUBS 0.010057f
C247 B.n134 VSUBS 0.010057f
C248 B.n135 VSUBS 0.010057f
C249 B.n136 VSUBS 0.010057f
C250 B.n137 VSUBS 0.010057f
C251 B.n138 VSUBS 0.010057f
C252 B.n139 VSUBS 0.010057f
C253 B.n140 VSUBS 0.010057f
C254 B.n141 VSUBS 0.010057f
C255 B.n142 VSUBS 0.007025f
C256 B.n143 VSUBS 0.010057f
C257 B.n144 VSUBS 0.010057f
C258 B.n145 VSUBS 0.010057f
C259 B.n146 VSUBS 0.010057f
C260 B.n147 VSUBS 0.010057f
C261 B.t5 VSUBS 0.338688f
C262 B.t4 VSUBS 0.379398f
C263 B.t3 VSUBS 2.08146f
C264 B.n148 VSUBS 0.224234f
C265 B.n149 VSUBS 0.110569f
C266 B.n150 VSUBS 0.010057f
C267 B.n151 VSUBS 0.010057f
C268 B.n152 VSUBS 0.010057f
C269 B.n153 VSUBS 0.010057f
C270 B.n154 VSUBS 0.010057f
C271 B.n155 VSUBS 0.010057f
C272 B.n156 VSUBS 0.010057f
C273 B.n157 VSUBS 0.010057f
C274 B.n158 VSUBS 0.010057f
C275 B.n159 VSUBS 0.010057f
C276 B.n160 VSUBS 0.010057f
C277 B.n161 VSUBS 0.010057f
C278 B.n162 VSUBS 0.010057f
C279 B.n163 VSUBS 0.02469f
C280 B.n164 VSUBS 0.010057f
C281 B.n165 VSUBS 0.010057f
C282 B.n166 VSUBS 0.010057f
C283 B.n167 VSUBS 0.010057f
C284 B.n168 VSUBS 0.010057f
C285 B.n169 VSUBS 0.010057f
C286 B.n170 VSUBS 0.010057f
C287 B.n171 VSUBS 0.010057f
C288 B.n172 VSUBS 0.010057f
C289 B.n173 VSUBS 0.010057f
C290 B.n174 VSUBS 0.010057f
C291 B.n175 VSUBS 0.010057f
C292 B.n176 VSUBS 0.010057f
C293 B.n177 VSUBS 0.010057f
C294 B.n178 VSUBS 0.010057f
C295 B.n179 VSUBS 0.010057f
C296 B.n180 VSUBS 0.010057f
C297 B.n181 VSUBS 0.010057f
C298 B.n182 VSUBS 0.010057f
C299 B.n183 VSUBS 0.010057f
C300 B.n184 VSUBS 0.010057f
C301 B.n185 VSUBS 0.010057f
C302 B.n186 VSUBS 0.010057f
C303 B.n187 VSUBS 0.010057f
C304 B.n188 VSUBS 0.010057f
C305 B.n189 VSUBS 0.010057f
C306 B.n190 VSUBS 0.010057f
C307 B.n191 VSUBS 0.010057f
C308 B.n192 VSUBS 0.010057f
C309 B.n193 VSUBS 0.010057f
C310 B.n194 VSUBS 0.010057f
C311 B.n195 VSUBS 0.010057f
C312 B.n196 VSUBS 0.010057f
C313 B.n197 VSUBS 0.010057f
C314 B.n198 VSUBS 0.010057f
C315 B.n199 VSUBS 0.010057f
C316 B.n200 VSUBS 0.010057f
C317 B.n201 VSUBS 0.010057f
C318 B.n202 VSUBS 0.010057f
C319 B.n203 VSUBS 0.010057f
C320 B.n204 VSUBS 0.010057f
C321 B.n205 VSUBS 0.010057f
C322 B.n206 VSUBS 0.010057f
C323 B.n207 VSUBS 0.010057f
C324 B.n208 VSUBS 0.010057f
C325 B.n209 VSUBS 0.010057f
C326 B.n210 VSUBS 0.010057f
C327 B.n211 VSUBS 0.010057f
C328 B.n212 VSUBS 0.010057f
C329 B.n213 VSUBS 0.010057f
C330 B.n214 VSUBS 0.010057f
C331 B.n215 VSUBS 0.010057f
C332 B.n216 VSUBS 0.010057f
C333 B.n217 VSUBS 0.010057f
C334 B.n218 VSUBS 0.010057f
C335 B.n219 VSUBS 0.010057f
C336 B.n220 VSUBS 0.010057f
C337 B.n221 VSUBS 0.010057f
C338 B.n222 VSUBS 0.010057f
C339 B.n223 VSUBS 0.010057f
C340 B.n224 VSUBS 0.010057f
C341 B.n225 VSUBS 0.010057f
C342 B.n226 VSUBS 0.010057f
C343 B.n227 VSUBS 0.010057f
C344 B.n228 VSUBS 0.010057f
C345 B.n229 VSUBS 0.010057f
C346 B.n230 VSUBS 0.010057f
C347 B.n231 VSUBS 0.010057f
C348 B.n232 VSUBS 0.010057f
C349 B.n233 VSUBS 0.010057f
C350 B.n234 VSUBS 0.010057f
C351 B.n235 VSUBS 0.010057f
C352 B.n236 VSUBS 0.010057f
C353 B.n237 VSUBS 0.010057f
C354 B.n238 VSUBS 0.010057f
C355 B.n239 VSUBS 0.010057f
C356 B.n240 VSUBS 0.010057f
C357 B.n241 VSUBS 0.010057f
C358 B.n242 VSUBS 0.010057f
C359 B.n243 VSUBS 0.010057f
C360 B.n244 VSUBS 0.010057f
C361 B.n245 VSUBS 0.010057f
C362 B.n246 VSUBS 0.010057f
C363 B.n247 VSUBS 0.010057f
C364 B.n248 VSUBS 0.010057f
C365 B.n249 VSUBS 0.010057f
C366 B.n250 VSUBS 0.010057f
C367 B.n251 VSUBS 0.010057f
C368 B.n252 VSUBS 0.010057f
C369 B.n253 VSUBS 0.010057f
C370 B.n254 VSUBS 0.010057f
C371 B.n255 VSUBS 0.010057f
C372 B.n256 VSUBS 0.010057f
C373 B.n257 VSUBS 0.010057f
C374 B.n258 VSUBS 0.010057f
C375 B.n259 VSUBS 0.010057f
C376 B.n260 VSUBS 0.010057f
C377 B.n261 VSUBS 0.010057f
C378 B.n262 VSUBS 0.010057f
C379 B.n263 VSUBS 0.010057f
C380 B.n264 VSUBS 0.010057f
C381 B.n265 VSUBS 0.010057f
C382 B.n266 VSUBS 0.010057f
C383 B.n267 VSUBS 0.010057f
C384 B.n268 VSUBS 0.010057f
C385 B.n269 VSUBS 0.010057f
C386 B.n270 VSUBS 0.010057f
C387 B.n271 VSUBS 0.010057f
C388 B.n272 VSUBS 0.010057f
C389 B.n273 VSUBS 0.010057f
C390 B.n274 VSUBS 0.010057f
C391 B.n275 VSUBS 0.010057f
C392 B.n276 VSUBS 0.024114f
C393 B.n277 VSUBS 0.024114f
C394 B.n278 VSUBS 0.02469f
C395 B.n279 VSUBS 0.010057f
C396 B.n280 VSUBS 0.010057f
C397 B.n281 VSUBS 0.010057f
C398 B.n282 VSUBS 0.010057f
C399 B.n283 VSUBS 0.010057f
C400 B.n284 VSUBS 0.010057f
C401 B.n285 VSUBS 0.010057f
C402 B.n286 VSUBS 0.010057f
C403 B.n287 VSUBS 0.010057f
C404 B.n288 VSUBS 0.010057f
C405 B.n289 VSUBS 0.010057f
C406 B.n290 VSUBS 0.010057f
C407 B.n291 VSUBS 0.010057f
C408 B.n292 VSUBS 0.010057f
C409 B.n293 VSUBS 0.010057f
C410 B.n294 VSUBS 0.010057f
C411 B.n295 VSUBS 0.010057f
C412 B.n296 VSUBS 0.010057f
C413 B.n297 VSUBS 0.010057f
C414 B.n298 VSUBS 0.010057f
C415 B.n299 VSUBS 0.010057f
C416 B.n300 VSUBS 0.010057f
C417 B.n301 VSUBS 0.010057f
C418 B.n302 VSUBS 0.010057f
C419 B.n303 VSUBS 0.010057f
C420 B.n304 VSUBS 0.010057f
C421 B.n305 VSUBS 0.010057f
C422 B.n306 VSUBS 0.010057f
C423 B.n307 VSUBS 0.010057f
C424 B.n308 VSUBS 0.010057f
C425 B.n309 VSUBS 0.010057f
C426 B.n310 VSUBS 0.010057f
C427 B.n311 VSUBS 0.010057f
C428 B.n312 VSUBS 0.010057f
C429 B.n313 VSUBS 0.010057f
C430 B.n314 VSUBS 0.010057f
C431 B.n315 VSUBS 0.010057f
C432 B.n316 VSUBS 0.010057f
C433 B.n317 VSUBS 0.010057f
C434 B.n318 VSUBS 0.010057f
C435 B.n319 VSUBS 0.010057f
C436 B.n320 VSUBS 0.007025f
C437 B.n321 VSUBS 0.0233f
C438 B.n322 VSUBS 0.00806f
C439 B.n323 VSUBS 0.010057f
C440 B.n324 VSUBS 0.010057f
C441 B.n325 VSUBS 0.010057f
C442 B.n326 VSUBS 0.010057f
C443 B.n327 VSUBS 0.010057f
C444 B.n328 VSUBS 0.010057f
C445 B.n329 VSUBS 0.010057f
C446 B.n330 VSUBS 0.010057f
C447 B.n331 VSUBS 0.010057f
C448 B.n332 VSUBS 0.010057f
C449 B.n333 VSUBS 0.010057f
C450 B.t2 VSUBS 0.338685f
C451 B.t1 VSUBS 0.379395f
C452 B.t0 VSUBS 2.08159f
C453 B.n334 VSUBS 0.224107f
C454 B.n335 VSUBS 0.110572f
C455 B.n336 VSUBS 0.0233f
C456 B.n337 VSUBS 0.00806f
C457 B.n338 VSUBS 0.010057f
C458 B.n339 VSUBS 0.010057f
C459 B.n340 VSUBS 0.010057f
C460 B.n341 VSUBS 0.010057f
C461 B.n342 VSUBS 0.010057f
C462 B.n343 VSUBS 0.010057f
C463 B.n344 VSUBS 0.010057f
C464 B.n345 VSUBS 0.010057f
C465 B.n346 VSUBS 0.010057f
C466 B.n347 VSUBS 0.010057f
C467 B.n348 VSUBS 0.010057f
C468 B.n349 VSUBS 0.010057f
C469 B.n350 VSUBS 0.010057f
C470 B.n351 VSUBS 0.010057f
C471 B.n352 VSUBS 0.010057f
C472 B.n353 VSUBS 0.010057f
C473 B.n354 VSUBS 0.010057f
C474 B.n355 VSUBS 0.010057f
C475 B.n356 VSUBS 0.010057f
C476 B.n357 VSUBS 0.010057f
C477 B.n358 VSUBS 0.010057f
C478 B.n359 VSUBS 0.010057f
C479 B.n360 VSUBS 0.010057f
C480 B.n361 VSUBS 0.010057f
C481 B.n362 VSUBS 0.010057f
C482 B.n363 VSUBS 0.010057f
C483 B.n364 VSUBS 0.010057f
C484 B.n365 VSUBS 0.010057f
C485 B.n366 VSUBS 0.010057f
C486 B.n367 VSUBS 0.010057f
C487 B.n368 VSUBS 0.010057f
C488 B.n369 VSUBS 0.010057f
C489 B.n370 VSUBS 0.010057f
C490 B.n371 VSUBS 0.010057f
C491 B.n372 VSUBS 0.010057f
C492 B.n373 VSUBS 0.010057f
C493 B.n374 VSUBS 0.010057f
C494 B.n375 VSUBS 0.010057f
C495 B.n376 VSUBS 0.010057f
C496 B.n377 VSUBS 0.010057f
C497 B.n378 VSUBS 0.010057f
C498 B.n379 VSUBS 0.010057f
C499 B.n380 VSUBS 0.010057f
C500 B.n381 VSUBS 0.02469f
C501 B.n382 VSUBS 0.024114f
C502 B.n383 VSUBS 0.025239f
C503 B.n384 VSUBS 0.010057f
C504 B.n385 VSUBS 0.010057f
C505 B.n386 VSUBS 0.010057f
C506 B.n387 VSUBS 0.010057f
C507 B.n388 VSUBS 0.010057f
C508 B.n389 VSUBS 0.010057f
C509 B.n390 VSUBS 0.010057f
C510 B.n391 VSUBS 0.010057f
C511 B.n392 VSUBS 0.010057f
C512 B.n393 VSUBS 0.010057f
C513 B.n394 VSUBS 0.010057f
C514 B.n395 VSUBS 0.010057f
C515 B.n396 VSUBS 0.010057f
C516 B.n397 VSUBS 0.010057f
C517 B.n398 VSUBS 0.010057f
C518 B.n399 VSUBS 0.010057f
C519 B.n400 VSUBS 0.010057f
C520 B.n401 VSUBS 0.010057f
C521 B.n402 VSUBS 0.010057f
C522 B.n403 VSUBS 0.010057f
C523 B.n404 VSUBS 0.010057f
C524 B.n405 VSUBS 0.010057f
C525 B.n406 VSUBS 0.010057f
C526 B.n407 VSUBS 0.010057f
C527 B.n408 VSUBS 0.010057f
C528 B.n409 VSUBS 0.010057f
C529 B.n410 VSUBS 0.010057f
C530 B.n411 VSUBS 0.010057f
C531 B.n412 VSUBS 0.010057f
C532 B.n413 VSUBS 0.010057f
C533 B.n414 VSUBS 0.010057f
C534 B.n415 VSUBS 0.010057f
C535 B.n416 VSUBS 0.010057f
C536 B.n417 VSUBS 0.010057f
C537 B.n418 VSUBS 0.010057f
C538 B.n419 VSUBS 0.010057f
C539 B.n420 VSUBS 0.010057f
C540 B.n421 VSUBS 0.010057f
C541 B.n422 VSUBS 0.010057f
C542 B.n423 VSUBS 0.010057f
C543 B.n424 VSUBS 0.010057f
C544 B.n425 VSUBS 0.010057f
C545 B.n426 VSUBS 0.010057f
C546 B.n427 VSUBS 0.010057f
C547 B.n428 VSUBS 0.010057f
C548 B.n429 VSUBS 0.010057f
C549 B.n430 VSUBS 0.010057f
C550 B.n431 VSUBS 0.010057f
C551 B.n432 VSUBS 0.010057f
C552 B.n433 VSUBS 0.010057f
C553 B.n434 VSUBS 0.010057f
C554 B.n435 VSUBS 0.010057f
C555 B.n436 VSUBS 0.010057f
C556 B.n437 VSUBS 0.010057f
C557 B.n438 VSUBS 0.010057f
C558 B.n439 VSUBS 0.010057f
C559 B.n440 VSUBS 0.010057f
C560 B.n441 VSUBS 0.010057f
C561 B.n442 VSUBS 0.010057f
C562 B.n443 VSUBS 0.010057f
C563 B.n444 VSUBS 0.010057f
C564 B.n445 VSUBS 0.010057f
C565 B.n446 VSUBS 0.010057f
C566 B.n447 VSUBS 0.010057f
C567 B.n448 VSUBS 0.010057f
C568 B.n449 VSUBS 0.010057f
C569 B.n450 VSUBS 0.010057f
C570 B.n451 VSUBS 0.010057f
C571 B.n452 VSUBS 0.010057f
C572 B.n453 VSUBS 0.010057f
C573 B.n454 VSUBS 0.010057f
C574 B.n455 VSUBS 0.010057f
C575 B.n456 VSUBS 0.010057f
C576 B.n457 VSUBS 0.010057f
C577 B.n458 VSUBS 0.010057f
C578 B.n459 VSUBS 0.010057f
C579 B.n460 VSUBS 0.010057f
C580 B.n461 VSUBS 0.010057f
C581 B.n462 VSUBS 0.010057f
C582 B.n463 VSUBS 0.010057f
C583 B.n464 VSUBS 0.010057f
C584 B.n465 VSUBS 0.010057f
C585 B.n466 VSUBS 0.010057f
C586 B.n467 VSUBS 0.010057f
C587 B.n468 VSUBS 0.010057f
C588 B.n469 VSUBS 0.010057f
C589 B.n470 VSUBS 0.010057f
C590 B.n471 VSUBS 0.010057f
C591 B.n472 VSUBS 0.010057f
C592 B.n473 VSUBS 0.010057f
C593 B.n474 VSUBS 0.010057f
C594 B.n475 VSUBS 0.010057f
C595 B.n476 VSUBS 0.010057f
C596 B.n477 VSUBS 0.010057f
C597 B.n478 VSUBS 0.010057f
C598 B.n479 VSUBS 0.010057f
C599 B.n480 VSUBS 0.010057f
C600 B.n481 VSUBS 0.010057f
C601 B.n482 VSUBS 0.010057f
C602 B.n483 VSUBS 0.010057f
C603 B.n484 VSUBS 0.010057f
C604 B.n485 VSUBS 0.010057f
C605 B.n486 VSUBS 0.010057f
C606 B.n487 VSUBS 0.010057f
C607 B.n488 VSUBS 0.010057f
C608 B.n489 VSUBS 0.010057f
C609 B.n490 VSUBS 0.010057f
C610 B.n491 VSUBS 0.010057f
C611 B.n492 VSUBS 0.010057f
C612 B.n493 VSUBS 0.010057f
C613 B.n494 VSUBS 0.010057f
C614 B.n495 VSUBS 0.010057f
C615 B.n496 VSUBS 0.010057f
C616 B.n497 VSUBS 0.010057f
C617 B.n498 VSUBS 0.010057f
C618 B.n499 VSUBS 0.010057f
C619 B.n500 VSUBS 0.010057f
C620 B.n501 VSUBS 0.010057f
C621 B.n502 VSUBS 0.010057f
C622 B.n503 VSUBS 0.010057f
C623 B.n504 VSUBS 0.010057f
C624 B.n505 VSUBS 0.010057f
C625 B.n506 VSUBS 0.010057f
C626 B.n507 VSUBS 0.010057f
C627 B.n508 VSUBS 0.010057f
C628 B.n509 VSUBS 0.010057f
C629 B.n510 VSUBS 0.010057f
C630 B.n511 VSUBS 0.010057f
C631 B.n512 VSUBS 0.010057f
C632 B.n513 VSUBS 0.010057f
C633 B.n514 VSUBS 0.010057f
C634 B.n515 VSUBS 0.010057f
C635 B.n516 VSUBS 0.010057f
C636 B.n517 VSUBS 0.010057f
C637 B.n518 VSUBS 0.010057f
C638 B.n519 VSUBS 0.010057f
C639 B.n520 VSUBS 0.010057f
C640 B.n521 VSUBS 0.010057f
C641 B.n522 VSUBS 0.010057f
C642 B.n523 VSUBS 0.010057f
C643 B.n524 VSUBS 0.010057f
C644 B.n525 VSUBS 0.010057f
C645 B.n526 VSUBS 0.010057f
C646 B.n527 VSUBS 0.010057f
C647 B.n528 VSUBS 0.010057f
C648 B.n529 VSUBS 0.010057f
C649 B.n530 VSUBS 0.010057f
C650 B.n531 VSUBS 0.010057f
C651 B.n532 VSUBS 0.010057f
C652 B.n533 VSUBS 0.010057f
C653 B.n534 VSUBS 0.010057f
C654 B.n535 VSUBS 0.010057f
C655 B.n536 VSUBS 0.010057f
C656 B.n537 VSUBS 0.010057f
C657 B.n538 VSUBS 0.010057f
C658 B.n539 VSUBS 0.010057f
C659 B.n540 VSUBS 0.010057f
C660 B.n541 VSUBS 0.010057f
C661 B.n542 VSUBS 0.010057f
C662 B.n543 VSUBS 0.010057f
C663 B.n544 VSUBS 0.010057f
C664 B.n545 VSUBS 0.010057f
C665 B.n546 VSUBS 0.010057f
C666 B.n547 VSUBS 0.010057f
C667 B.n548 VSUBS 0.010057f
C668 B.n549 VSUBS 0.010057f
C669 B.n550 VSUBS 0.010057f
C670 B.n551 VSUBS 0.010057f
C671 B.n552 VSUBS 0.010057f
C672 B.n553 VSUBS 0.010057f
C673 B.n554 VSUBS 0.010057f
C674 B.n555 VSUBS 0.010057f
C675 B.n556 VSUBS 0.010057f
C676 B.n557 VSUBS 0.010057f
C677 B.n558 VSUBS 0.024114f
C678 B.n559 VSUBS 0.02469f
C679 B.n560 VSUBS 0.02469f
C680 B.n561 VSUBS 0.010057f
C681 B.n562 VSUBS 0.010057f
C682 B.n563 VSUBS 0.010057f
C683 B.n564 VSUBS 0.010057f
C684 B.n565 VSUBS 0.010057f
C685 B.n566 VSUBS 0.010057f
C686 B.n567 VSUBS 0.010057f
C687 B.n568 VSUBS 0.010057f
C688 B.n569 VSUBS 0.010057f
C689 B.n570 VSUBS 0.010057f
C690 B.n571 VSUBS 0.010057f
C691 B.n572 VSUBS 0.010057f
C692 B.n573 VSUBS 0.010057f
C693 B.n574 VSUBS 0.010057f
C694 B.n575 VSUBS 0.010057f
C695 B.n576 VSUBS 0.010057f
C696 B.n577 VSUBS 0.010057f
C697 B.n578 VSUBS 0.010057f
C698 B.n579 VSUBS 0.010057f
C699 B.n580 VSUBS 0.010057f
C700 B.n581 VSUBS 0.010057f
C701 B.n582 VSUBS 0.010057f
C702 B.n583 VSUBS 0.010057f
C703 B.n584 VSUBS 0.010057f
C704 B.n585 VSUBS 0.010057f
C705 B.n586 VSUBS 0.010057f
C706 B.n587 VSUBS 0.010057f
C707 B.n588 VSUBS 0.010057f
C708 B.n589 VSUBS 0.010057f
C709 B.n590 VSUBS 0.010057f
C710 B.n591 VSUBS 0.010057f
C711 B.n592 VSUBS 0.010057f
C712 B.n593 VSUBS 0.010057f
C713 B.n594 VSUBS 0.010057f
C714 B.n595 VSUBS 0.010057f
C715 B.n596 VSUBS 0.010057f
C716 B.n597 VSUBS 0.010057f
C717 B.n598 VSUBS 0.010057f
C718 B.n599 VSUBS 0.010057f
C719 B.n600 VSUBS 0.010057f
C720 B.n601 VSUBS 0.007025f
C721 B.n602 VSUBS 0.010057f
C722 B.n603 VSUBS 0.010057f
C723 B.n604 VSUBS 0.00806f
C724 B.n605 VSUBS 0.010057f
C725 B.n606 VSUBS 0.010057f
C726 B.n607 VSUBS 0.010057f
C727 B.n608 VSUBS 0.010057f
C728 B.n609 VSUBS 0.010057f
C729 B.n610 VSUBS 0.010057f
C730 B.n611 VSUBS 0.010057f
C731 B.n612 VSUBS 0.010057f
C732 B.n613 VSUBS 0.010057f
C733 B.n614 VSUBS 0.010057f
C734 B.n615 VSUBS 0.010057f
C735 B.n616 VSUBS 0.00806f
C736 B.n617 VSUBS 0.0233f
C737 B.n618 VSUBS 0.007025f
C738 B.n619 VSUBS 0.010057f
C739 B.n620 VSUBS 0.010057f
C740 B.n621 VSUBS 0.010057f
C741 B.n622 VSUBS 0.010057f
C742 B.n623 VSUBS 0.010057f
C743 B.n624 VSUBS 0.010057f
C744 B.n625 VSUBS 0.010057f
C745 B.n626 VSUBS 0.010057f
C746 B.n627 VSUBS 0.010057f
C747 B.n628 VSUBS 0.010057f
C748 B.n629 VSUBS 0.010057f
C749 B.n630 VSUBS 0.010057f
C750 B.n631 VSUBS 0.010057f
C751 B.n632 VSUBS 0.010057f
C752 B.n633 VSUBS 0.010057f
C753 B.n634 VSUBS 0.010057f
C754 B.n635 VSUBS 0.010057f
C755 B.n636 VSUBS 0.010057f
C756 B.n637 VSUBS 0.010057f
C757 B.n638 VSUBS 0.010057f
C758 B.n639 VSUBS 0.010057f
C759 B.n640 VSUBS 0.010057f
C760 B.n641 VSUBS 0.010057f
C761 B.n642 VSUBS 0.010057f
C762 B.n643 VSUBS 0.010057f
C763 B.n644 VSUBS 0.010057f
C764 B.n645 VSUBS 0.010057f
C765 B.n646 VSUBS 0.010057f
C766 B.n647 VSUBS 0.010057f
C767 B.n648 VSUBS 0.010057f
C768 B.n649 VSUBS 0.010057f
C769 B.n650 VSUBS 0.010057f
C770 B.n651 VSUBS 0.010057f
C771 B.n652 VSUBS 0.010057f
C772 B.n653 VSUBS 0.010057f
C773 B.n654 VSUBS 0.010057f
C774 B.n655 VSUBS 0.010057f
C775 B.n656 VSUBS 0.010057f
C776 B.n657 VSUBS 0.010057f
C777 B.n658 VSUBS 0.010057f
C778 B.n659 VSUBS 0.010057f
C779 B.n660 VSUBS 0.02469f
C780 B.n661 VSUBS 0.024114f
C781 B.n662 VSUBS 0.024114f
C782 B.n663 VSUBS 0.010057f
C783 B.n664 VSUBS 0.010057f
C784 B.n665 VSUBS 0.010057f
C785 B.n666 VSUBS 0.010057f
C786 B.n667 VSUBS 0.010057f
C787 B.n668 VSUBS 0.010057f
C788 B.n669 VSUBS 0.010057f
C789 B.n670 VSUBS 0.010057f
C790 B.n671 VSUBS 0.010057f
C791 B.n672 VSUBS 0.010057f
C792 B.n673 VSUBS 0.010057f
C793 B.n674 VSUBS 0.010057f
C794 B.n675 VSUBS 0.010057f
C795 B.n676 VSUBS 0.010057f
C796 B.n677 VSUBS 0.010057f
C797 B.n678 VSUBS 0.010057f
C798 B.n679 VSUBS 0.010057f
C799 B.n680 VSUBS 0.010057f
C800 B.n681 VSUBS 0.010057f
C801 B.n682 VSUBS 0.010057f
C802 B.n683 VSUBS 0.010057f
C803 B.n684 VSUBS 0.010057f
C804 B.n685 VSUBS 0.010057f
C805 B.n686 VSUBS 0.010057f
C806 B.n687 VSUBS 0.010057f
C807 B.n688 VSUBS 0.010057f
C808 B.n689 VSUBS 0.010057f
C809 B.n690 VSUBS 0.010057f
C810 B.n691 VSUBS 0.010057f
C811 B.n692 VSUBS 0.010057f
C812 B.n693 VSUBS 0.010057f
C813 B.n694 VSUBS 0.010057f
C814 B.n695 VSUBS 0.010057f
C815 B.n696 VSUBS 0.010057f
C816 B.n697 VSUBS 0.010057f
C817 B.n698 VSUBS 0.010057f
C818 B.n699 VSUBS 0.010057f
C819 B.n700 VSUBS 0.010057f
C820 B.n701 VSUBS 0.010057f
C821 B.n702 VSUBS 0.010057f
C822 B.n703 VSUBS 0.010057f
C823 B.n704 VSUBS 0.010057f
C824 B.n705 VSUBS 0.010057f
C825 B.n706 VSUBS 0.010057f
C826 B.n707 VSUBS 0.010057f
C827 B.n708 VSUBS 0.010057f
C828 B.n709 VSUBS 0.010057f
C829 B.n710 VSUBS 0.010057f
C830 B.n711 VSUBS 0.010057f
C831 B.n712 VSUBS 0.010057f
C832 B.n713 VSUBS 0.010057f
C833 B.n714 VSUBS 0.010057f
C834 B.n715 VSUBS 0.010057f
C835 B.n716 VSUBS 0.010057f
C836 B.n717 VSUBS 0.010057f
C837 B.n718 VSUBS 0.010057f
C838 B.n719 VSUBS 0.010057f
C839 B.n720 VSUBS 0.010057f
C840 B.n721 VSUBS 0.010057f
C841 B.n722 VSUBS 0.010057f
C842 B.n723 VSUBS 0.010057f
C843 B.n724 VSUBS 0.010057f
C844 B.n725 VSUBS 0.010057f
C845 B.n726 VSUBS 0.010057f
C846 B.n727 VSUBS 0.010057f
C847 B.n728 VSUBS 0.010057f
C848 B.n729 VSUBS 0.010057f
C849 B.n730 VSUBS 0.010057f
C850 B.n731 VSUBS 0.010057f
C851 B.n732 VSUBS 0.010057f
C852 B.n733 VSUBS 0.010057f
C853 B.n734 VSUBS 0.010057f
C854 B.n735 VSUBS 0.010057f
C855 B.n736 VSUBS 0.010057f
C856 B.n737 VSUBS 0.010057f
C857 B.n738 VSUBS 0.010057f
C858 B.n739 VSUBS 0.010057f
C859 B.n740 VSUBS 0.010057f
C860 B.n741 VSUBS 0.010057f
C861 B.n742 VSUBS 0.010057f
C862 B.n743 VSUBS 0.010057f
C863 B.n744 VSUBS 0.010057f
C864 B.n745 VSUBS 0.010057f
C865 B.n746 VSUBS 0.010057f
C866 B.n747 VSUBS 0.013124f
C867 B.n748 VSUBS 0.01398f
C868 B.n749 VSUBS 0.0278f
C869 VDD2.t5 VSUBS 1.752f
C870 VDD2.t4 VSUBS 0.184853f
C871 VDD2.t1 VSUBS 0.184853f
C872 VDD2.n0 VSUBS 1.31051f
C873 VDD2.n1 VSUBS 4.48733f
C874 VDD2.t2 VSUBS 1.7247f
C875 VDD2.n2 VSUBS 3.72947f
C876 VDD2.t0 VSUBS 0.184853f
C877 VDD2.t3 VSUBS 0.184853f
C878 VDD2.n3 VSUBS 1.31047f
C879 VTAIL.t11 VSUBS 0.200142f
C880 VTAIL.t7 VSUBS 0.200142f
C881 VTAIL.n0 VSUBS 1.26062f
C882 VTAIL.n1 VSUBS 1.03251f
C883 VTAIL.t3 VSUBS 1.70862f
C884 VTAIL.n2 VSUBS 1.41785f
C885 VTAIL.t4 VSUBS 0.200142f
C886 VTAIL.t5 VSUBS 0.200142f
C887 VTAIL.n3 VSUBS 1.26062f
C888 VTAIL.n4 VSUBS 3.00841f
C889 VTAIL.t8 VSUBS 0.200142f
C890 VTAIL.t10 VSUBS 0.200142f
C891 VTAIL.n5 VSUBS 1.26062f
C892 VTAIL.n6 VSUBS 3.0084f
C893 VTAIL.t6 VSUBS 1.70863f
C894 VTAIL.n7 VSUBS 1.41784f
C895 VTAIL.t2 VSUBS 0.200142f
C896 VTAIL.t0 VSUBS 0.200142f
C897 VTAIL.n8 VSUBS 1.26062f
C898 VTAIL.n9 VSUBS 1.32f
C899 VTAIL.t1 VSUBS 1.70862f
C900 VTAIL.n10 VSUBS 2.71468f
C901 VTAIL.t9 VSUBS 1.70862f
C902 VTAIL.n11 VSUBS 2.61063f
C903 VN.t4 VSUBS 2.35025f
C904 VN.n0 VSUBS 0.956517f
C905 VN.n1 VSUBS 0.028886f
C906 VN.n2 VSUBS 0.05755f
C907 VN.n3 VSUBS 0.028886f
C908 VN.n4 VSUBS 0.053836f
C909 VN.t0 VSUBS 2.79188f
C910 VN.n5 VSUBS 0.916177f
C911 VN.t1 VSUBS 2.35025f
C912 VN.n6 VSUBS 0.95146f
C913 VN.n7 VSUBS 0.040547f
C914 VN.n8 VSUBS 0.37775f
C915 VN.n9 VSUBS 0.028886f
C916 VN.n10 VSUBS 0.028886f
C917 VN.n11 VSUBS 0.053836f
C918 VN.n12 VSUBS 0.052447f
C919 VN.n13 VSUBS 0.028177f
C920 VN.n14 VSUBS 0.028886f
C921 VN.n15 VSUBS 0.028886f
C922 VN.n16 VSUBS 0.028886f
C923 VN.n17 VSUBS 0.053836f
C924 VN.n18 VSUBS 0.053836f
C925 VN.n19 VSUBS 0.028852f
C926 VN.n20 VSUBS 0.046622f
C927 VN.n21 VSUBS 0.092395f
C928 VN.t3 VSUBS 2.35025f
C929 VN.n22 VSUBS 0.956517f
C930 VN.n23 VSUBS 0.028886f
C931 VN.n24 VSUBS 0.05755f
C932 VN.n25 VSUBS 0.028886f
C933 VN.n26 VSUBS 0.053836f
C934 VN.t2 VSUBS 2.79188f
C935 VN.n27 VSUBS 0.916177f
C936 VN.t5 VSUBS 2.35025f
C937 VN.n28 VSUBS 0.95146f
C938 VN.n29 VSUBS 0.040547f
C939 VN.n30 VSUBS 0.37775f
C940 VN.n31 VSUBS 0.028886f
C941 VN.n32 VSUBS 0.028886f
C942 VN.n33 VSUBS 0.053836f
C943 VN.n34 VSUBS 0.052447f
C944 VN.n35 VSUBS 0.028177f
C945 VN.n36 VSUBS 0.028886f
C946 VN.n37 VSUBS 0.028886f
C947 VN.n38 VSUBS 0.028886f
C948 VN.n39 VSUBS 0.053836f
C949 VN.n40 VSUBS 0.053836f
C950 VN.n41 VSUBS 0.028852f
C951 VN.n42 VSUBS 0.046622f
C952 VN.n43 VSUBS 1.71519f
.ends

