* NGSPICE file created from diff_pair_sample_0862.ext - technology: sky130A

.subckt diff_pair_sample_0862 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1630_n2606# sky130_fd_pr__pfet_01v8 ad=3.89025 pd=17.33 as=0 ps=0 w=8.19 l=0.16
X1 VDD2.t7 VN.t0 VTAIL.t14 w_n1630_n2606# sky130_fd_pr__pfet_01v8 ad=2.0475 pd=8.69 as=2.0475 ps=8.69 w=8.19 l=0.16
X2 B.t8 B.t6 B.t7 w_n1630_n2606# sky130_fd_pr__pfet_01v8 ad=3.89025 pd=17.33 as=0 ps=0 w=8.19 l=0.16
X3 VDD2.t6 VN.t1 VTAIL.t13 w_n1630_n2606# sky130_fd_pr__pfet_01v8 ad=2.0475 pd=8.69 as=2.0475 ps=8.69 w=8.19 l=0.16
X4 B.t5 B.t3 B.t4 w_n1630_n2606# sky130_fd_pr__pfet_01v8 ad=3.89025 pd=17.33 as=0 ps=0 w=8.19 l=0.16
X5 VTAIL.t9 VN.t2 VDD2.t5 w_n1630_n2606# sky130_fd_pr__pfet_01v8 ad=3.89025 pd=17.33 as=2.0475 ps=8.69 w=8.19 l=0.16
X6 VDD1.t7 VP.t0 VTAIL.t15 w_n1630_n2606# sky130_fd_pr__pfet_01v8 ad=2.0475 pd=8.69 as=2.0475 ps=8.69 w=8.19 l=0.16
X7 VDD2.t4 VN.t3 VTAIL.t7 w_n1630_n2606# sky130_fd_pr__pfet_01v8 ad=2.0475 pd=8.69 as=3.89025 ps=17.33 w=8.19 l=0.16
X8 VDD2.t3 VN.t4 VTAIL.t8 w_n1630_n2606# sky130_fd_pr__pfet_01v8 ad=2.0475 pd=8.69 as=3.89025 ps=17.33 w=8.19 l=0.16
X9 VTAIL.t2 VP.t1 VDD1.t6 w_n1630_n2606# sky130_fd_pr__pfet_01v8 ad=3.89025 pd=17.33 as=2.0475 ps=8.69 w=8.19 l=0.16
X10 VTAIL.t11 VN.t5 VDD2.t2 w_n1630_n2606# sky130_fd_pr__pfet_01v8 ad=3.89025 pd=17.33 as=2.0475 ps=8.69 w=8.19 l=0.16
X11 B.t2 B.t0 B.t1 w_n1630_n2606# sky130_fd_pr__pfet_01v8 ad=3.89025 pd=17.33 as=0 ps=0 w=8.19 l=0.16
X12 VTAIL.t10 VN.t6 VDD2.t1 w_n1630_n2606# sky130_fd_pr__pfet_01v8 ad=2.0475 pd=8.69 as=2.0475 ps=8.69 w=8.19 l=0.16
X13 VDD1.t5 VP.t2 VTAIL.t1 w_n1630_n2606# sky130_fd_pr__pfet_01v8 ad=2.0475 pd=8.69 as=3.89025 ps=17.33 w=8.19 l=0.16
X14 VTAIL.t6 VP.t3 VDD1.t4 w_n1630_n2606# sky130_fd_pr__pfet_01v8 ad=2.0475 pd=8.69 as=2.0475 ps=8.69 w=8.19 l=0.16
X15 VTAIL.t5 VP.t4 VDD1.t3 w_n1630_n2606# sky130_fd_pr__pfet_01v8 ad=3.89025 pd=17.33 as=2.0475 ps=8.69 w=8.19 l=0.16
X16 VTAIL.t12 VN.t7 VDD2.t0 w_n1630_n2606# sky130_fd_pr__pfet_01v8 ad=2.0475 pd=8.69 as=2.0475 ps=8.69 w=8.19 l=0.16
X17 VDD1.t2 VP.t5 VTAIL.t0 w_n1630_n2606# sky130_fd_pr__pfet_01v8 ad=2.0475 pd=8.69 as=2.0475 ps=8.69 w=8.19 l=0.16
X18 VDD1.t1 VP.t6 VTAIL.t4 w_n1630_n2606# sky130_fd_pr__pfet_01v8 ad=2.0475 pd=8.69 as=3.89025 ps=17.33 w=8.19 l=0.16
X19 VTAIL.t3 VP.t7 VDD1.t0 w_n1630_n2606# sky130_fd_pr__pfet_01v8 ad=2.0475 pd=8.69 as=2.0475 ps=8.69 w=8.19 l=0.16
R0 B.n84 B.t3 1485.03
R1 B.n92 B.t0 1485.03
R2 B.n26 B.t9 1485.03
R3 B.n34 B.t6 1485.03
R4 B.n305 B.n50 585
R5 B.n307 B.n306 585
R6 B.n308 B.n49 585
R7 B.n310 B.n309 585
R8 B.n311 B.n48 585
R9 B.n313 B.n312 585
R10 B.n314 B.n47 585
R11 B.n316 B.n315 585
R12 B.n317 B.n46 585
R13 B.n319 B.n318 585
R14 B.n320 B.n45 585
R15 B.n322 B.n321 585
R16 B.n323 B.n44 585
R17 B.n325 B.n324 585
R18 B.n326 B.n43 585
R19 B.n328 B.n327 585
R20 B.n329 B.n42 585
R21 B.n331 B.n330 585
R22 B.n332 B.n41 585
R23 B.n334 B.n333 585
R24 B.n335 B.n40 585
R25 B.n337 B.n336 585
R26 B.n338 B.n39 585
R27 B.n340 B.n339 585
R28 B.n341 B.n38 585
R29 B.n343 B.n342 585
R30 B.n344 B.n37 585
R31 B.n346 B.n345 585
R32 B.n347 B.n36 585
R33 B.n349 B.n348 585
R34 B.n351 B.n33 585
R35 B.n353 B.n352 585
R36 B.n354 B.n32 585
R37 B.n356 B.n355 585
R38 B.n357 B.n31 585
R39 B.n359 B.n358 585
R40 B.n360 B.n30 585
R41 B.n362 B.n361 585
R42 B.n363 B.n29 585
R43 B.n365 B.n364 585
R44 B.n367 B.n366 585
R45 B.n368 B.n25 585
R46 B.n370 B.n369 585
R47 B.n371 B.n24 585
R48 B.n373 B.n372 585
R49 B.n374 B.n23 585
R50 B.n376 B.n375 585
R51 B.n377 B.n22 585
R52 B.n379 B.n378 585
R53 B.n380 B.n21 585
R54 B.n382 B.n381 585
R55 B.n383 B.n20 585
R56 B.n385 B.n384 585
R57 B.n386 B.n19 585
R58 B.n388 B.n387 585
R59 B.n389 B.n18 585
R60 B.n391 B.n390 585
R61 B.n392 B.n17 585
R62 B.n394 B.n393 585
R63 B.n395 B.n16 585
R64 B.n397 B.n396 585
R65 B.n398 B.n15 585
R66 B.n400 B.n399 585
R67 B.n401 B.n14 585
R68 B.n403 B.n402 585
R69 B.n404 B.n13 585
R70 B.n406 B.n405 585
R71 B.n407 B.n12 585
R72 B.n409 B.n408 585
R73 B.n410 B.n11 585
R74 B.n304 B.n303 585
R75 B.n302 B.n51 585
R76 B.n301 B.n300 585
R77 B.n299 B.n52 585
R78 B.n298 B.n297 585
R79 B.n296 B.n53 585
R80 B.n295 B.n294 585
R81 B.n293 B.n54 585
R82 B.n292 B.n291 585
R83 B.n290 B.n55 585
R84 B.n289 B.n288 585
R85 B.n287 B.n56 585
R86 B.n286 B.n285 585
R87 B.n284 B.n57 585
R88 B.n283 B.n282 585
R89 B.n281 B.n58 585
R90 B.n280 B.n279 585
R91 B.n278 B.n59 585
R92 B.n277 B.n276 585
R93 B.n275 B.n60 585
R94 B.n274 B.n273 585
R95 B.n272 B.n61 585
R96 B.n271 B.n270 585
R97 B.n269 B.n62 585
R98 B.n268 B.n267 585
R99 B.n266 B.n63 585
R100 B.n265 B.n264 585
R101 B.n263 B.n64 585
R102 B.n262 B.n261 585
R103 B.n260 B.n65 585
R104 B.n259 B.n258 585
R105 B.n257 B.n66 585
R106 B.n256 B.n255 585
R107 B.n254 B.n67 585
R108 B.n253 B.n252 585
R109 B.n251 B.n68 585
R110 B.n250 B.n249 585
R111 B.n143 B.n108 585
R112 B.n145 B.n144 585
R113 B.n146 B.n107 585
R114 B.n148 B.n147 585
R115 B.n149 B.n106 585
R116 B.n151 B.n150 585
R117 B.n152 B.n105 585
R118 B.n154 B.n153 585
R119 B.n155 B.n104 585
R120 B.n157 B.n156 585
R121 B.n158 B.n103 585
R122 B.n160 B.n159 585
R123 B.n161 B.n102 585
R124 B.n163 B.n162 585
R125 B.n164 B.n101 585
R126 B.n166 B.n165 585
R127 B.n167 B.n100 585
R128 B.n169 B.n168 585
R129 B.n170 B.n99 585
R130 B.n172 B.n171 585
R131 B.n173 B.n98 585
R132 B.n175 B.n174 585
R133 B.n176 B.n97 585
R134 B.n178 B.n177 585
R135 B.n179 B.n96 585
R136 B.n181 B.n180 585
R137 B.n182 B.n95 585
R138 B.n184 B.n183 585
R139 B.n185 B.n94 585
R140 B.n187 B.n186 585
R141 B.n189 B.n91 585
R142 B.n191 B.n190 585
R143 B.n192 B.n90 585
R144 B.n194 B.n193 585
R145 B.n195 B.n89 585
R146 B.n197 B.n196 585
R147 B.n198 B.n88 585
R148 B.n200 B.n199 585
R149 B.n201 B.n87 585
R150 B.n203 B.n202 585
R151 B.n205 B.n204 585
R152 B.n206 B.n83 585
R153 B.n208 B.n207 585
R154 B.n209 B.n82 585
R155 B.n211 B.n210 585
R156 B.n212 B.n81 585
R157 B.n214 B.n213 585
R158 B.n215 B.n80 585
R159 B.n217 B.n216 585
R160 B.n218 B.n79 585
R161 B.n220 B.n219 585
R162 B.n221 B.n78 585
R163 B.n223 B.n222 585
R164 B.n224 B.n77 585
R165 B.n226 B.n225 585
R166 B.n227 B.n76 585
R167 B.n229 B.n228 585
R168 B.n230 B.n75 585
R169 B.n232 B.n231 585
R170 B.n233 B.n74 585
R171 B.n235 B.n234 585
R172 B.n236 B.n73 585
R173 B.n238 B.n237 585
R174 B.n239 B.n72 585
R175 B.n241 B.n240 585
R176 B.n242 B.n71 585
R177 B.n244 B.n243 585
R178 B.n245 B.n70 585
R179 B.n247 B.n246 585
R180 B.n248 B.n69 585
R181 B.n142 B.n141 585
R182 B.n140 B.n109 585
R183 B.n139 B.n138 585
R184 B.n137 B.n110 585
R185 B.n136 B.n135 585
R186 B.n134 B.n111 585
R187 B.n133 B.n132 585
R188 B.n131 B.n112 585
R189 B.n130 B.n129 585
R190 B.n128 B.n113 585
R191 B.n127 B.n126 585
R192 B.n125 B.n114 585
R193 B.n124 B.n123 585
R194 B.n122 B.n115 585
R195 B.n121 B.n120 585
R196 B.n119 B.n116 585
R197 B.n118 B.n117 585
R198 B.n2 B.n0 585
R199 B.n437 B.n1 585
R200 B.n436 B.n435 585
R201 B.n434 B.n3 585
R202 B.n433 B.n432 585
R203 B.n431 B.n4 585
R204 B.n430 B.n429 585
R205 B.n428 B.n5 585
R206 B.n427 B.n426 585
R207 B.n425 B.n6 585
R208 B.n424 B.n423 585
R209 B.n422 B.n7 585
R210 B.n421 B.n420 585
R211 B.n419 B.n8 585
R212 B.n418 B.n417 585
R213 B.n416 B.n9 585
R214 B.n415 B.n414 585
R215 B.n413 B.n10 585
R216 B.n412 B.n411 585
R217 B.n439 B.n438 585
R218 B.n143 B.n142 502.111
R219 B.n412 B.n11 502.111
R220 B.n250 B.n69 502.111
R221 B.n305 B.n304 502.111
R222 B.n142 B.n109 163.367
R223 B.n138 B.n109 163.367
R224 B.n138 B.n137 163.367
R225 B.n137 B.n136 163.367
R226 B.n136 B.n111 163.367
R227 B.n132 B.n111 163.367
R228 B.n132 B.n131 163.367
R229 B.n131 B.n130 163.367
R230 B.n130 B.n113 163.367
R231 B.n126 B.n113 163.367
R232 B.n126 B.n125 163.367
R233 B.n125 B.n124 163.367
R234 B.n124 B.n115 163.367
R235 B.n120 B.n115 163.367
R236 B.n120 B.n119 163.367
R237 B.n119 B.n118 163.367
R238 B.n118 B.n2 163.367
R239 B.n438 B.n2 163.367
R240 B.n438 B.n437 163.367
R241 B.n437 B.n436 163.367
R242 B.n436 B.n3 163.367
R243 B.n432 B.n3 163.367
R244 B.n432 B.n431 163.367
R245 B.n431 B.n430 163.367
R246 B.n430 B.n5 163.367
R247 B.n426 B.n5 163.367
R248 B.n426 B.n425 163.367
R249 B.n425 B.n424 163.367
R250 B.n424 B.n7 163.367
R251 B.n420 B.n7 163.367
R252 B.n420 B.n419 163.367
R253 B.n419 B.n418 163.367
R254 B.n418 B.n9 163.367
R255 B.n414 B.n9 163.367
R256 B.n414 B.n413 163.367
R257 B.n413 B.n412 163.367
R258 B.n144 B.n143 163.367
R259 B.n144 B.n107 163.367
R260 B.n148 B.n107 163.367
R261 B.n149 B.n148 163.367
R262 B.n150 B.n149 163.367
R263 B.n150 B.n105 163.367
R264 B.n154 B.n105 163.367
R265 B.n155 B.n154 163.367
R266 B.n156 B.n155 163.367
R267 B.n156 B.n103 163.367
R268 B.n160 B.n103 163.367
R269 B.n161 B.n160 163.367
R270 B.n162 B.n161 163.367
R271 B.n162 B.n101 163.367
R272 B.n166 B.n101 163.367
R273 B.n167 B.n166 163.367
R274 B.n168 B.n167 163.367
R275 B.n168 B.n99 163.367
R276 B.n172 B.n99 163.367
R277 B.n173 B.n172 163.367
R278 B.n174 B.n173 163.367
R279 B.n174 B.n97 163.367
R280 B.n178 B.n97 163.367
R281 B.n179 B.n178 163.367
R282 B.n180 B.n179 163.367
R283 B.n180 B.n95 163.367
R284 B.n184 B.n95 163.367
R285 B.n185 B.n184 163.367
R286 B.n186 B.n185 163.367
R287 B.n186 B.n91 163.367
R288 B.n191 B.n91 163.367
R289 B.n192 B.n191 163.367
R290 B.n193 B.n192 163.367
R291 B.n193 B.n89 163.367
R292 B.n197 B.n89 163.367
R293 B.n198 B.n197 163.367
R294 B.n199 B.n198 163.367
R295 B.n199 B.n87 163.367
R296 B.n203 B.n87 163.367
R297 B.n204 B.n203 163.367
R298 B.n204 B.n83 163.367
R299 B.n208 B.n83 163.367
R300 B.n209 B.n208 163.367
R301 B.n210 B.n209 163.367
R302 B.n210 B.n81 163.367
R303 B.n214 B.n81 163.367
R304 B.n215 B.n214 163.367
R305 B.n216 B.n215 163.367
R306 B.n216 B.n79 163.367
R307 B.n220 B.n79 163.367
R308 B.n221 B.n220 163.367
R309 B.n222 B.n221 163.367
R310 B.n222 B.n77 163.367
R311 B.n226 B.n77 163.367
R312 B.n227 B.n226 163.367
R313 B.n228 B.n227 163.367
R314 B.n228 B.n75 163.367
R315 B.n232 B.n75 163.367
R316 B.n233 B.n232 163.367
R317 B.n234 B.n233 163.367
R318 B.n234 B.n73 163.367
R319 B.n238 B.n73 163.367
R320 B.n239 B.n238 163.367
R321 B.n240 B.n239 163.367
R322 B.n240 B.n71 163.367
R323 B.n244 B.n71 163.367
R324 B.n245 B.n244 163.367
R325 B.n246 B.n245 163.367
R326 B.n246 B.n69 163.367
R327 B.n251 B.n250 163.367
R328 B.n252 B.n251 163.367
R329 B.n252 B.n67 163.367
R330 B.n256 B.n67 163.367
R331 B.n257 B.n256 163.367
R332 B.n258 B.n257 163.367
R333 B.n258 B.n65 163.367
R334 B.n262 B.n65 163.367
R335 B.n263 B.n262 163.367
R336 B.n264 B.n263 163.367
R337 B.n264 B.n63 163.367
R338 B.n268 B.n63 163.367
R339 B.n269 B.n268 163.367
R340 B.n270 B.n269 163.367
R341 B.n270 B.n61 163.367
R342 B.n274 B.n61 163.367
R343 B.n275 B.n274 163.367
R344 B.n276 B.n275 163.367
R345 B.n276 B.n59 163.367
R346 B.n280 B.n59 163.367
R347 B.n281 B.n280 163.367
R348 B.n282 B.n281 163.367
R349 B.n282 B.n57 163.367
R350 B.n286 B.n57 163.367
R351 B.n287 B.n286 163.367
R352 B.n288 B.n287 163.367
R353 B.n288 B.n55 163.367
R354 B.n292 B.n55 163.367
R355 B.n293 B.n292 163.367
R356 B.n294 B.n293 163.367
R357 B.n294 B.n53 163.367
R358 B.n298 B.n53 163.367
R359 B.n299 B.n298 163.367
R360 B.n300 B.n299 163.367
R361 B.n300 B.n51 163.367
R362 B.n304 B.n51 163.367
R363 B.n408 B.n11 163.367
R364 B.n408 B.n407 163.367
R365 B.n407 B.n406 163.367
R366 B.n406 B.n13 163.367
R367 B.n402 B.n13 163.367
R368 B.n402 B.n401 163.367
R369 B.n401 B.n400 163.367
R370 B.n400 B.n15 163.367
R371 B.n396 B.n15 163.367
R372 B.n396 B.n395 163.367
R373 B.n395 B.n394 163.367
R374 B.n394 B.n17 163.367
R375 B.n390 B.n17 163.367
R376 B.n390 B.n389 163.367
R377 B.n389 B.n388 163.367
R378 B.n388 B.n19 163.367
R379 B.n384 B.n19 163.367
R380 B.n384 B.n383 163.367
R381 B.n383 B.n382 163.367
R382 B.n382 B.n21 163.367
R383 B.n378 B.n21 163.367
R384 B.n378 B.n377 163.367
R385 B.n377 B.n376 163.367
R386 B.n376 B.n23 163.367
R387 B.n372 B.n23 163.367
R388 B.n372 B.n371 163.367
R389 B.n371 B.n370 163.367
R390 B.n370 B.n25 163.367
R391 B.n366 B.n25 163.367
R392 B.n366 B.n365 163.367
R393 B.n365 B.n29 163.367
R394 B.n361 B.n29 163.367
R395 B.n361 B.n360 163.367
R396 B.n360 B.n359 163.367
R397 B.n359 B.n31 163.367
R398 B.n355 B.n31 163.367
R399 B.n355 B.n354 163.367
R400 B.n354 B.n353 163.367
R401 B.n353 B.n33 163.367
R402 B.n348 B.n33 163.367
R403 B.n348 B.n347 163.367
R404 B.n347 B.n346 163.367
R405 B.n346 B.n37 163.367
R406 B.n342 B.n37 163.367
R407 B.n342 B.n341 163.367
R408 B.n341 B.n340 163.367
R409 B.n340 B.n39 163.367
R410 B.n336 B.n39 163.367
R411 B.n336 B.n335 163.367
R412 B.n335 B.n334 163.367
R413 B.n334 B.n41 163.367
R414 B.n330 B.n41 163.367
R415 B.n330 B.n329 163.367
R416 B.n329 B.n328 163.367
R417 B.n328 B.n43 163.367
R418 B.n324 B.n43 163.367
R419 B.n324 B.n323 163.367
R420 B.n323 B.n322 163.367
R421 B.n322 B.n45 163.367
R422 B.n318 B.n45 163.367
R423 B.n318 B.n317 163.367
R424 B.n317 B.n316 163.367
R425 B.n316 B.n47 163.367
R426 B.n312 B.n47 163.367
R427 B.n312 B.n311 163.367
R428 B.n311 B.n310 163.367
R429 B.n310 B.n49 163.367
R430 B.n306 B.n49 163.367
R431 B.n306 B.n305 163.367
R432 B.n84 B.t5 123.957
R433 B.n34 B.t7 123.957
R434 B.n92 B.t2 123.948
R435 B.n26 B.t10 123.948
R436 B.n85 B.t4 111.156
R437 B.n35 B.t8 111.156
R438 B.n93 B.t1 111.147
R439 B.n27 B.t11 111.147
R440 B.n86 B.n85 59.5399
R441 B.n188 B.n93 59.5399
R442 B.n28 B.n27 59.5399
R443 B.n350 B.n35 59.5399
R444 B.n411 B.n410 32.6249
R445 B.n303 B.n50 32.6249
R446 B.n249 B.n248 32.6249
R447 B.n141 B.n108 32.6249
R448 B B.n439 18.0485
R449 B.n85 B.n84 12.8005
R450 B.n93 B.n92 12.8005
R451 B.n27 B.n26 12.8005
R452 B.n35 B.n34 12.8005
R453 B.n410 B.n409 10.6151
R454 B.n409 B.n12 10.6151
R455 B.n405 B.n12 10.6151
R456 B.n405 B.n404 10.6151
R457 B.n404 B.n403 10.6151
R458 B.n403 B.n14 10.6151
R459 B.n399 B.n14 10.6151
R460 B.n399 B.n398 10.6151
R461 B.n398 B.n397 10.6151
R462 B.n397 B.n16 10.6151
R463 B.n393 B.n16 10.6151
R464 B.n393 B.n392 10.6151
R465 B.n392 B.n391 10.6151
R466 B.n391 B.n18 10.6151
R467 B.n387 B.n18 10.6151
R468 B.n387 B.n386 10.6151
R469 B.n386 B.n385 10.6151
R470 B.n385 B.n20 10.6151
R471 B.n381 B.n20 10.6151
R472 B.n381 B.n380 10.6151
R473 B.n380 B.n379 10.6151
R474 B.n379 B.n22 10.6151
R475 B.n375 B.n22 10.6151
R476 B.n375 B.n374 10.6151
R477 B.n374 B.n373 10.6151
R478 B.n373 B.n24 10.6151
R479 B.n369 B.n24 10.6151
R480 B.n369 B.n368 10.6151
R481 B.n368 B.n367 10.6151
R482 B.n364 B.n363 10.6151
R483 B.n363 B.n362 10.6151
R484 B.n362 B.n30 10.6151
R485 B.n358 B.n30 10.6151
R486 B.n358 B.n357 10.6151
R487 B.n357 B.n356 10.6151
R488 B.n356 B.n32 10.6151
R489 B.n352 B.n32 10.6151
R490 B.n352 B.n351 10.6151
R491 B.n349 B.n36 10.6151
R492 B.n345 B.n36 10.6151
R493 B.n345 B.n344 10.6151
R494 B.n344 B.n343 10.6151
R495 B.n343 B.n38 10.6151
R496 B.n339 B.n38 10.6151
R497 B.n339 B.n338 10.6151
R498 B.n338 B.n337 10.6151
R499 B.n337 B.n40 10.6151
R500 B.n333 B.n40 10.6151
R501 B.n333 B.n332 10.6151
R502 B.n332 B.n331 10.6151
R503 B.n331 B.n42 10.6151
R504 B.n327 B.n42 10.6151
R505 B.n327 B.n326 10.6151
R506 B.n326 B.n325 10.6151
R507 B.n325 B.n44 10.6151
R508 B.n321 B.n44 10.6151
R509 B.n321 B.n320 10.6151
R510 B.n320 B.n319 10.6151
R511 B.n319 B.n46 10.6151
R512 B.n315 B.n46 10.6151
R513 B.n315 B.n314 10.6151
R514 B.n314 B.n313 10.6151
R515 B.n313 B.n48 10.6151
R516 B.n309 B.n48 10.6151
R517 B.n309 B.n308 10.6151
R518 B.n308 B.n307 10.6151
R519 B.n307 B.n50 10.6151
R520 B.n249 B.n68 10.6151
R521 B.n253 B.n68 10.6151
R522 B.n254 B.n253 10.6151
R523 B.n255 B.n254 10.6151
R524 B.n255 B.n66 10.6151
R525 B.n259 B.n66 10.6151
R526 B.n260 B.n259 10.6151
R527 B.n261 B.n260 10.6151
R528 B.n261 B.n64 10.6151
R529 B.n265 B.n64 10.6151
R530 B.n266 B.n265 10.6151
R531 B.n267 B.n266 10.6151
R532 B.n267 B.n62 10.6151
R533 B.n271 B.n62 10.6151
R534 B.n272 B.n271 10.6151
R535 B.n273 B.n272 10.6151
R536 B.n273 B.n60 10.6151
R537 B.n277 B.n60 10.6151
R538 B.n278 B.n277 10.6151
R539 B.n279 B.n278 10.6151
R540 B.n279 B.n58 10.6151
R541 B.n283 B.n58 10.6151
R542 B.n284 B.n283 10.6151
R543 B.n285 B.n284 10.6151
R544 B.n285 B.n56 10.6151
R545 B.n289 B.n56 10.6151
R546 B.n290 B.n289 10.6151
R547 B.n291 B.n290 10.6151
R548 B.n291 B.n54 10.6151
R549 B.n295 B.n54 10.6151
R550 B.n296 B.n295 10.6151
R551 B.n297 B.n296 10.6151
R552 B.n297 B.n52 10.6151
R553 B.n301 B.n52 10.6151
R554 B.n302 B.n301 10.6151
R555 B.n303 B.n302 10.6151
R556 B.n145 B.n108 10.6151
R557 B.n146 B.n145 10.6151
R558 B.n147 B.n146 10.6151
R559 B.n147 B.n106 10.6151
R560 B.n151 B.n106 10.6151
R561 B.n152 B.n151 10.6151
R562 B.n153 B.n152 10.6151
R563 B.n153 B.n104 10.6151
R564 B.n157 B.n104 10.6151
R565 B.n158 B.n157 10.6151
R566 B.n159 B.n158 10.6151
R567 B.n159 B.n102 10.6151
R568 B.n163 B.n102 10.6151
R569 B.n164 B.n163 10.6151
R570 B.n165 B.n164 10.6151
R571 B.n165 B.n100 10.6151
R572 B.n169 B.n100 10.6151
R573 B.n170 B.n169 10.6151
R574 B.n171 B.n170 10.6151
R575 B.n171 B.n98 10.6151
R576 B.n175 B.n98 10.6151
R577 B.n176 B.n175 10.6151
R578 B.n177 B.n176 10.6151
R579 B.n177 B.n96 10.6151
R580 B.n181 B.n96 10.6151
R581 B.n182 B.n181 10.6151
R582 B.n183 B.n182 10.6151
R583 B.n183 B.n94 10.6151
R584 B.n187 B.n94 10.6151
R585 B.n190 B.n189 10.6151
R586 B.n190 B.n90 10.6151
R587 B.n194 B.n90 10.6151
R588 B.n195 B.n194 10.6151
R589 B.n196 B.n195 10.6151
R590 B.n196 B.n88 10.6151
R591 B.n200 B.n88 10.6151
R592 B.n201 B.n200 10.6151
R593 B.n202 B.n201 10.6151
R594 B.n206 B.n205 10.6151
R595 B.n207 B.n206 10.6151
R596 B.n207 B.n82 10.6151
R597 B.n211 B.n82 10.6151
R598 B.n212 B.n211 10.6151
R599 B.n213 B.n212 10.6151
R600 B.n213 B.n80 10.6151
R601 B.n217 B.n80 10.6151
R602 B.n218 B.n217 10.6151
R603 B.n219 B.n218 10.6151
R604 B.n219 B.n78 10.6151
R605 B.n223 B.n78 10.6151
R606 B.n224 B.n223 10.6151
R607 B.n225 B.n224 10.6151
R608 B.n225 B.n76 10.6151
R609 B.n229 B.n76 10.6151
R610 B.n230 B.n229 10.6151
R611 B.n231 B.n230 10.6151
R612 B.n231 B.n74 10.6151
R613 B.n235 B.n74 10.6151
R614 B.n236 B.n235 10.6151
R615 B.n237 B.n236 10.6151
R616 B.n237 B.n72 10.6151
R617 B.n241 B.n72 10.6151
R618 B.n242 B.n241 10.6151
R619 B.n243 B.n242 10.6151
R620 B.n243 B.n70 10.6151
R621 B.n247 B.n70 10.6151
R622 B.n248 B.n247 10.6151
R623 B.n141 B.n140 10.6151
R624 B.n140 B.n139 10.6151
R625 B.n139 B.n110 10.6151
R626 B.n135 B.n110 10.6151
R627 B.n135 B.n134 10.6151
R628 B.n134 B.n133 10.6151
R629 B.n133 B.n112 10.6151
R630 B.n129 B.n112 10.6151
R631 B.n129 B.n128 10.6151
R632 B.n128 B.n127 10.6151
R633 B.n127 B.n114 10.6151
R634 B.n123 B.n114 10.6151
R635 B.n123 B.n122 10.6151
R636 B.n122 B.n121 10.6151
R637 B.n121 B.n116 10.6151
R638 B.n117 B.n116 10.6151
R639 B.n117 B.n0 10.6151
R640 B.n435 B.n1 10.6151
R641 B.n435 B.n434 10.6151
R642 B.n434 B.n433 10.6151
R643 B.n433 B.n4 10.6151
R644 B.n429 B.n4 10.6151
R645 B.n429 B.n428 10.6151
R646 B.n428 B.n427 10.6151
R647 B.n427 B.n6 10.6151
R648 B.n423 B.n6 10.6151
R649 B.n423 B.n422 10.6151
R650 B.n422 B.n421 10.6151
R651 B.n421 B.n8 10.6151
R652 B.n417 B.n8 10.6151
R653 B.n417 B.n416 10.6151
R654 B.n416 B.n415 10.6151
R655 B.n415 B.n10 10.6151
R656 B.n411 B.n10 10.6151
R657 B.n367 B.n28 9.36635
R658 B.n350 B.n349 9.36635
R659 B.n188 B.n187 9.36635
R660 B.n205 B.n86 9.36635
R661 B.n439 B.n0 2.81026
R662 B.n439 B.n1 2.81026
R663 B.n364 B.n28 1.24928
R664 B.n351 B.n350 1.24928
R665 B.n189 B.n188 1.24928
R666 B.n202 B.n86 1.24928
R667 VN.n7 VN.t4 1465.99
R668 VN.n2 VN.t2 1465.99
R669 VN.n16 VN.t5 1465.99
R670 VN.n11 VN.t3 1465.99
R671 VN.n6 VN.t7 1430.94
R672 VN.n1 VN.t1 1430.94
R673 VN.n15 VN.t0 1430.94
R674 VN.n10 VN.t6 1430.94
R675 VN.n12 VN.n11 161.489
R676 VN.n3 VN.n2 161.489
R677 VN.n8 VN.n7 161.3
R678 VN.n17 VN.n16 161.3
R679 VN.n14 VN.n9 161.3
R680 VN.n13 VN.n12 161.3
R681 VN.n5 VN.n0 161.3
R682 VN.n4 VN.n3 161.3
R683 VN.n5 VN.n4 73.0308
R684 VN.n14 VN.n13 73.0308
R685 VN.n2 VN.n1 61.346
R686 VN.n7 VN.n6 61.346
R687 VN.n16 VN.n15 61.346
R688 VN.n11 VN.n10 61.346
R689 VN VN.n17 37.813
R690 VN.n4 VN.n1 11.6853
R691 VN.n6 VN.n5 11.6853
R692 VN.n15 VN.n14 11.6853
R693 VN.n13 VN.n10 11.6853
R694 VN.n17 VN.n9 0.189894
R695 VN.n12 VN.n9 0.189894
R696 VN.n3 VN.n0 0.189894
R697 VN.n8 VN.n0 0.189894
R698 VN VN.n8 0.0516364
R699 VTAIL.n11 VTAIL.t5 71.2012
R700 VTAIL.n10 VTAIL.t7 71.2012
R701 VTAIL.n7 VTAIL.t11 71.2012
R702 VTAIL.n15 VTAIL.t8 71.2011
R703 VTAIL.n2 VTAIL.t9 71.2011
R704 VTAIL.n3 VTAIL.t1 71.2011
R705 VTAIL.n6 VTAIL.t2 71.2011
R706 VTAIL.n14 VTAIL.t4 71.2011
R707 VTAIL.n13 VTAIL.n12 65.1879
R708 VTAIL.n9 VTAIL.n8 65.1879
R709 VTAIL.n1 VTAIL.n0 65.1876
R710 VTAIL.n5 VTAIL.n4 65.1876
R711 VTAIL.n15 VTAIL.n14 19.9962
R712 VTAIL.n7 VTAIL.n6 19.9962
R713 VTAIL.n0 VTAIL.t13 6.01393
R714 VTAIL.n0 VTAIL.t12 6.01393
R715 VTAIL.n4 VTAIL.t0 6.01393
R716 VTAIL.n4 VTAIL.t3 6.01393
R717 VTAIL.n12 VTAIL.t15 6.01393
R718 VTAIL.n12 VTAIL.t6 6.01393
R719 VTAIL.n8 VTAIL.t14 6.01393
R720 VTAIL.n8 VTAIL.t10 6.01393
R721 VTAIL.n9 VTAIL.n7 0.569465
R722 VTAIL.n10 VTAIL.n9 0.569465
R723 VTAIL.n13 VTAIL.n11 0.569465
R724 VTAIL.n14 VTAIL.n13 0.569465
R725 VTAIL.n6 VTAIL.n5 0.569465
R726 VTAIL.n5 VTAIL.n3 0.569465
R727 VTAIL.n2 VTAIL.n1 0.569465
R728 VTAIL VTAIL.n15 0.511276
R729 VTAIL.n11 VTAIL.n10 0.470328
R730 VTAIL.n3 VTAIL.n2 0.470328
R731 VTAIL VTAIL.n1 0.0586897
R732 VDD2.n2 VDD2.n1 82.0955
R733 VDD2.n2 VDD2.n0 82.0955
R734 VDD2 VDD2.n5 82.0928
R735 VDD2.n4 VDD2.n3 81.8667
R736 VDD2.n4 VDD2.n2 33.336
R737 VDD2.n5 VDD2.t1 6.01393
R738 VDD2.n5 VDD2.t4 6.01393
R739 VDD2.n3 VDD2.t2 6.01393
R740 VDD2.n3 VDD2.t7 6.01393
R741 VDD2.n1 VDD2.t0 6.01393
R742 VDD2.n1 VDD2.t3 6.01393
R743 VDD2.n0 VDD2.t5 6.01393
R744 VDD2.n0 VDD2.t6 6.01393
R745 VDD2 VDD2.n4 0.343172
R746 VP.n17 VP.t2 1465.99
R747 VP.n11 VP.t1 1465.99
R748 VP.n4 VP.t4 1465.99
R749 VP.n9 VP.t6 1465.99
R750 VP.n16 VP.t7 1430.94
R751 VP.n1 VP.t5 1430.94
R752 VP.n3 VP.t0 1430.94
R753 VP.n8 VP.t3 1430.94
R754 VP.n5 VP.n4 161.489
R755 VP.n18 VP.n17 161.3
R756 VP.n6 VP.n5 161.3
R757 VP.n7 VP.n2 161.3
R758 VP.n10 VP.n9 161.3
R759 VP.n15 VP.n0 161.3
R760 VP.n14 VP.n13 161.3
R761 VP.n12 VP.n11 161.3
R762 VP.n15 VP.n14 73.0308
R763 VP.n7 VP.n6 73.0308
R764 VP.n11 VP.n1 61.346
R765 VP.n17 VP.n16 61.346
R766 VP.n4 VP.n3 61.346
R767 VP.n9 VP.n8 61.346
R768 VP.n12 VP.n10 37.4323
R769 VP.n14 VP.n1 11.6853
R770 VP.n16 VP.n15 11.6853
R771 VP.n6 VP.n3 11.6853
R772 VP.n8 VP.n7 11.6853
R773 VP.n5 VP.n2 0.189894
R774 VP.n10 VP.n2 0.189894
R775 VP.n13 VP.n12 0.189894
R776 VP.n13 VP.n0 0.189894
R777 VP.n18 VP.n0 0.189894
R778 VP VP.n18 0.0516364
R779 VDD1 VDD1.n0 82.2093
R780 VDD1.n3 VDD1.n2 82.0955
R781 VDD1.n3 VDD1.n1 82.0955
R782 VDD1.n5 VDD1.n4 81.8665
R783 VDD1.n5 VDD1.n3 33.919
R784 VDD1.n4 VDD1.t4 6.01393
R785 VDD1.n4 VDD1.t1 6.01393
R786 VDD1.n0 VDD1.t3 6.01393
R787 VDD1.n0 VDD1.t7 6.01393
R788 VDD1.n2 VDD1.t0 6.01393
R789 VDD1.n2 VDD1.t5 6.01393
R790 VDD1.n1 VDD1.t6 6.01393
R791 VDD1.n1 VDD1.t2 6.01393
R792 VDD1 VDD1.n5 0.226793
C0 VTAIL VDD1 11.856f
C1 w_n1630_n2606# VN 2.54377f
C2 VTAIL VN 1.26818f
C3 B VDD2 0.885003f
C4 B VP 0.960312f
C5 VDD2 VP 0.277496f
C6 B w_n1630_n2606# 5.57439f
C7 w_n1630_n2606# VDD2 1.06955f
C8 B VTAIL 2.54648f
C9 VN VDD1 0.147059f
C10 w_n1630_n2606# VP 2.74868f
C11 VTAIL VDD2 11.895201f
C12 VTAIL VP 1.28229f
C13 VTAIL w_n1630_n2606# 3.32141f
C14 B VDD1 0.859737f
C15 VDD2 VDD1 0.644877f
C16 B VN 0.628951f
C17 VDD1 VP 1.77107f
C18 VDD2 VN 1.64072f
C19 w_n1630_n2606# VDD1 1.04998f
C20 VN VP 4.16925f
C21 VDD2 VSUBS 1.042468f
C22 VDD1 VSUBS 1.262319f
C23 VTAIL VSUBS 0.596113f
C24 VN VSUBS 3.48465f
C25 VP VSUBS 0.965152f
C26 B VSUBS 2.068122f
C27 w_n1630_n2606# VSUBS 52.675102f
C28 VDD1.t3 VSUBS 0.238618f
C29 VDD1.t7 VSUBS 0.238618f
C30 VDD1.n0 VSUBS 1.30732f
C31 VDD1.t6 VSUBS 0.238618f
C32 VDD1.t2 VSUBS 0.238618f
C33 VDD1.n1 VSUBS 1.30661f
C34 VDD1.t0 VSUBS 0.238618f
C35 VDD1.t5 VSUBS 0.238618f
C36 VDD1.n2 VSUBS 1.30661f
C37 VDD1.n3 VSUBS 2.16684f
C38 VDD1.t4 VSUBS 0.238618f
C39 VDD1.t1 VSUBS 0.238618f
C40 VDD1.n4 VSUBS 1.30524f
C41 VDD1.n5 VSUBS 2.05717f
C42 VP.n0 VSUBS 0.05689f
C43 VP.t7 VSUBS 0.211555f
C44 VP.t5 VSUBS 0.211555f
C45 VP.n1 VSUBS 0.098316f
C46 VP.n2 VSUBS 0.05689f
C47 VP.t3 VSUBS 0.211555f
C48 VP.t0 VSUBS 0.211555f
C49 VP.n3 VSUBS 0.098316f
C50 VP.t4 VSUBS 0.213823f
C51 VP.n4 VSUBS 0.117098f
C52 VP.n5 VSUBS 0.118618f
C53 VP.n6 VSUBS 0.021678f
C54 VP.n7 VSUBS 0.021678f
C55 VP.n8 VSUBS 0.098316f
C56 VP.t6 VSUBS 0.213823f
C57 VP.n9 VSUBS 0.117026f
C58 VP.n10 VSUBS 1.92231f
C59 VP.t1 VSUBS 0.213823f
C60 VP.n11 VSUBS 0.117026f
C61 VP.n12 VSUBS 1.97694f
C62 VP.n13 VSUBS 0.05689f
C63 VP.n14 VSUBS 0.021678f
C64 VP.n15 VSUBS 0.021678f
C65 VP.n16 VSUBS 0.098316f
C66 VP.t2 VSUBS 0.213823f
C67 VP.n17 VSUBS 0.117026f
C68 VP.n18 VSUBS 0.044087f
C69 VDD2.t5 VSUBS 0.240434f
C70 VDD2.t6 VSUBS 0.240434f
C71 VDD2.n0 VSUBS 1.31656f
C72 VDD2.t0 VSUBS 0.240434f
C73 VDD2.t3 VSUBS 0.240434f
C74 VDD2.n1 VSUBS 1.31656f
C75 VDD2.n2 VSUBS 2.13052f
C76 VDD2.t2 VSUBS 0.240434f
C77 VDD2.t7 VSUBS 0.240434f
C78 VDD2.n3 VSUBS 1.31518f
C79 VDD2.n4 VSUBS 2.04425f
C80 VDD2.t1 VSUBS 0.240434f
C81 VDD2.t4 VSUBS 0.240434f
C82 VDD2.n5 VSUBS 1.31653f
C83 VTAIL.t13 VSUBS 0.233903f
C84 VTAIL.t12 VSUBS 0.233903f
C85 VTAIL.n0 VSUBS 1.17591f
C86 VTAIL.n1 VSUBS 0.528528f
C87 VTAIL.t9 VSUBS 1.48182f
C88 VTAIL.n2 VSUBS 0.675288f
C89 VTAIL.t1 VSUBS 1.48182f
C90 VTAIL.n3 VSUBS 0.675288f
C91 VTAIL.t0 VSUBS 0.233903f
C92 VTAIL.t3 VSUBS 0.233903f
C93 VTAIL.n4 VSUBS 1.17591f
C94 VTAIL.n5 VSUBS 0.567786f
C95 VTAIL.t2 VSUBS 1.48182f
C96 VTAIL.n6 VSUBS 1.54958f
C97 VTAIL.t11 VSUBS 1.48183f
C98 VTAIL.n7 VSUBS 1.54957f
C99 VTAIL.t14 VSUBS 0.233903f
C100 VTAIL.t10 VSUBS 0.233903f
C101 VTAIL.n8 VSUBS 1.17592f
C102 VTAIL.n9 VSUBS 0.567782f
C103 VTAIL.t7 VSUBS 1.48183f
C104 VTAIL.n10 VSUBS 0.675278f
C105 VTAIL.t5 VSUBS 1.48183f
C106 VTAIL.n11 VSUBS 0.675278f
C107 VTAIL.t15 VSUBS 0.233903f
C108 VTAIL.t6 VSUBS 0.233903f
C109 VTAIL.n12 VSUBS 1.17592f
C110 VTAIL.n13 VSUBS 0.567782f
C111 VTAIL.t4 VSUBS 1.48182f
C112 VTAIL.n14 VSUBS 1.54958f
C113 VTAIL.t8 VSUBS 1.48182f
C114 VTAIL.n15 VSUBS 1.5451f
C115 VN.n0 VSUBS 0.054608f
C116 VN.t7 VSUBS 0.20307f
C117 VN.t1 VSUBS 0.20307f
C118 VN.n1 VSUBS 0.094373f
C119 VN.t2 VSUBS 0.205246f
C120 VN.n2 VSUBS 0.112402f
C121 VN.n3 VSUBS 0.11386f
C122 VN.n4 VSUBS 0.020809f
C123 VN.n5 VSUBS 0.020809f
C124 VN.n6 VSUBS 0.094373f
C125 VN.t4 VSUBS 0.205246f
C126 VN.n7 VSUBS 0.112332f
C127 VN.n8 VSUBS 0.042319f
C128 VN.n9 VSUBS 0.054608f
C129 VN.t5 VSUBS 0.205246f
C130 VN.t0 VSUBS 0.20307f
C131 VN.t6 VSUBS 0.20307f
C132 VN.n10 VSUBS 0.094373f
C133 VN.t3 VSUBS 0.205246f
C134 VN.n11 VSUBS 0.112402f
C135 VN.n12 VSUBS 0.11386f
C136 VN.n13 VSUBS 0.020809f
C137 VN.n14 VSUBS 0.020809f
C138 VN.n15 VSUBS 0.094373f
C139 VN.n16 VSUBS 0.112332f
C140 VN.n17 VSUBS 1.88132f
C141 B.n0 VSUBS 0.005708f
C142 B.n1 VSUBS 0.005708f
C143 B.n2 VSUBS 0.009026f
C144 B.n3 VSUBS 0.009026f
C145 B.n4 VSUBS 0.009026f
C146 B.n5 VSUBS 0.009026f
C147 B.n6 VSUBS 0.009026f
C148 B.n7 VSUBS 0.009026f
C149 B.n8 VSUBS 0.009026f
C150 B.n9 VSUBS 0.009026f
C151 B.n10 VSUBS 0.009026f
C152 B.n11 VSUBS 0.021275f
C153 B.n12 VSUBS 0.009026f
C154 B.n13 VSUBS 0.009026f
C155 B.n14 VSUBS 0.009026f
C156 B.n15 VSUBS 0.009026f
C157 B.n16 VSUBS 0.009026f
C158 B.n17 VSUBS 0.009026f
C159 B.n18 VSUBS 0.009026f
C160 B.n19 VSUBS 0.009026f
C161 B.n20 VSUBS 0.009026f
C162 B.n21 VSUBS 0.009026f
C163 B.n22 VSUBS 0.009026f
C164 B.n23 VSUBS 0.009026f
C165 B.n24 VSUBS 0.009026f
C166 B.n25 VSUBS 0.009026f
C167 B.t11 VSUBS 0.365813f
C168 B.t10 VSUBS 0.373401f
C169 B.t9 VSUBS 0.065762f
C170 B.n26 VSUBS 0.099085f
C171 B.n27 VSUBS 0.086357f
C172 B.n28 VSUBS 0.020913f
C173 B.n29 VSUBS 0.009026f
C174 B.n30 VSUBS 0.009026f
C175 B.n31 VSUBS 0.009026f
C176 B.n32 VSUBS 0.009026f
C177 B.n33 VSUBS 0.009026f
C178 B.t8 VSUBS 0.365811f
C179 B.t7 VSUBS 0.373399f
C180 B.t6 VSUBS 0.065762f
C181 B.n34 VSUBS 0.099088f
C182 B.n35 VSUBS 0.086359f
C183 B.n36 VSUBS 0.009026f
C184 B.n37 VSUBS 0.009026f
C185 B.n38 VSUBS 0.009026f
C186 B.n39 VSUBS 0.009026f
C187 B.n40 VSUBS 0.009026f
C188 B.n41 VSUBS 0.009026f
C189 B.n42 VSUBS 0.009026f
C190 B.n43 VSUBS 0.009026f
C191 B.n44 VSUBS 0.009026f
C192 B.n45 VSUBS 0.009026f
C193 B.n46 VSUBS 0.009026f
C194 B.n47 VSUBS 0.009026f
C195 B.n48 VSUBS 0.009026f
C196 B.n49 VSUBS 0.009026f
C197 B.n50 VSUBS 0.020207f
C198 B.n51 VSUBS 0.009026f
C199 B.n52 VSUBS 0.009026f
C200 B.n53 VSUBS 0.009026f
C201 B.n54 VSUBS 0.009026f
C202 B.n55 VSUBS 0.009026f
C203 B.n56 VSUBS 0.009026f
C204 B.n57 VSUBS 0.009026f
C205 B.n58 VSUBS 0.009026f
C206 B.n59 VSUBS 0.009026f
C207 B.n60 VSUBS 0.009026f
C208 B.n61 VSUBS 0.009026f
C209 B.n62 VSUBS 0.009026f
C210 B.n63 VSUBS 0.009026f
C211 B.n64 VSUBS 0.009026f
C212 B.n65 VSUBS 0.009026f
C213 B.n66 VSUBS 0.009026f
C214 B.n67 VSUBS 0.009026f
C215 B.n68 VSUBS 0.009026f
C216 B.n69 VSUBS 0.021275f
C217 B.n70 VSUBS 0.009026f
C218 B.n71 VSUBS 0.009026f
C219 B.n72 VSUBS 0.009026f
C220 B.n73 VSUBS 0.009026f
C221 B.n74 VSUBS 0.009026f
C222 B.n75 VSUBS 0.009026f
C223 B.n76 VSUBS 0.009026f
C224 B.n77 VSUBS 0.009026f
C225 B.n78 VSUBS 0.009026f
C226 B.n79 VSUBS 0.009026f
C227 B.n80 VSUBS 0.009026f
C228 B.n81 VSUBS 0.009026f
C229 B.n82 VSUBS 0.009026f
C230 B.n83 VSUBS 0.009026f
C231 B.t4 VSUBS 0.365811f
C232 B.t5 VSUBS 0.373399f
C233 B.t3 VSUBS 0.065762f
C234 B.n84 VSUBS 0.099088f
C235 B.n85 VSUBS 0.086359f
C236 B.n86 VSUBS 0.020913f
C237 B.n87 VSUBS 0.009026f
C238 B.n88 VSUBS 0.009026f
C239 B.n89 VSUBS 0.009026f
C240 B.n90 VSUBS 0.009026f
C241 B.n91 VSUBS 0.009026f
C242 B.t1 VSUBS 0.365813f
C243 B.t2 VSUBS 0.373401f
C244 B.t0 VSUBS 0.065762f
C245 B.n92 VSUBS 0.099085f
C246 B.n93 VSUBS 0.086357f
C247 B.n94 VSUBS 0.009026f
C248 B.n95 VSUBS 0.009026f
C249 B.n96 VSUBS 0.009026f
C250 B.n97 VSUBS 0.009026f
C251 B.n98 VSUBS 0.009026f
C252 B.n99 VSUBS 0.009026f
C253 B.n100 VSUBS 0.009026f
C254 B.n101 VSUBS 0.009026f
C255 B.n102 VSUBS 0.009026f
C256 B.n103 VSUBS 0.009026f
C257 B.n104 VSUBS 0.009026f
C258 B.n105 VSUBS 0.009026f
C259 B.n106 VSUBS 0.009026f
C260 B.n107 VSUBS 0.009026f
C261 B.n108 VSUBS 0.021275f
C262 B.n109 VSUBS 0.009026f
C263 B.n110 VSUBS 0.009026f
C264 B.n111 VSUBS 0.009026f
C265 B.n112 VSUBS 0.009026f
C266 B.n113 VSUBS 0.009026f
C267 B.n114 VSUBS 0.009026f
C268 B.n115 VSUBS 0.009026f
C269 B.n116 VSUBS 0.009026f
C270 B.n117 VSUBS 0.009026f
C271 B.n118 VSUBS 0.009026f
C272 B.n119 VSUBS 0.009026f
C273 B.n120 VSUBS 0.009026f
C274 B.n121 VSUBS 0.009026f
C275 B.n122 VSUBS 0.009026f
C276 B.n123 VSUBS 0.009026f
C277 B.n124 VSUBS 0.009026f
C278 B.n125 VSUBS 0.009026f
C279 B.n126 VSUBS 0.009026f
C280 B.n127 VSUBS 0.009026f
C281 B.n128 VSUBS 0.009026f
C282 B.n129 VSUBS 0.009026f
C283 B.n130 VSUBS 0.009026f
C284 B.n131 VSUBS 0.009026f
C285 B.n132 VSUBS 0.009026f
C286 B.n133 VSUBS 0.009026f
C287 B.n134 VSUBS 0.009026f
C288 B.n135 VSUBS 0.009026f
C289 B.n136 VSUBS 0.009026f
C290 B.n137 VSUBS 0.009026f
C291 B.n138 VSUBS 0.009026f
C292 B.n139 VSUBS 0.009026f
C293 B.n140 VSUBS 0.009026f
C294 B.n141 VSUBS 0.020936f
C295 B.n142 VSUBS 0.020936f
C296 B.n143 VSUBS 0.021275f
C297 B.n144 VSUBS 0.009026f
C298 B.n145 VSUBS 0.009026f
C299 B.n146 VSUBS 0.009026f
C300 B.n147 VSUBS 0.009026f
C301 B.n148 VSUBS 0.009026f
C302 B.n149 VSUBS 0.009026f
C303 B.n150 VSUBS 0.009026f
C304 B.n151 VSUBS 0.009026f
C305 B.n152 VSUBS 0.009026f
C306 B.n153 VSUBS 0.009026f
C307 B.n154 VSUBS 0.009026f
C308 B.n155 VSUBS 0.009026f
C309 B.n156 VSUBS 0.009026f
C310 B.n157 VSUBS 0.009026f
C311 B.n158 VSUBS 0.009026f
C312 B.n159 VSUBS 0.009026f
C313 B.n160 VSUBS 0.009026f
C314 B.n161 VSUBS 0.009026f
C315 B.n162 VSUBS 0.009026f
C316 B.n163 VSUBS 0.009026f
C317 B.n164 VSUBS 0.009026f
C318 B.n165 VSUBS 0.009026f
C319 B.n166 VSUBS 0.009026f
C320 B.n167 VSUBS 0.009026f
C321 B.n168 VSUBS 0.009026f
C322 B.n169 VSUBS 0.009026f
C323 B.n170 VSUBS 0.009026f
C324 B.n171 VSUBS 0.009026f
C325 B.n172 VSUBS 0.009026f
C326 B.n173 VSUBS 0.009026f
C327 B.n174 VSUBS 0.009026f
C328 B.n175 VSUBS 0.009026f
C329 B.n176 VSUBS 0.009026f
C330 B.n177 VSUBS 0.009026f
C331 B.n178 VSUBS 0.009026f
C332 B.n179 VSUBS 0.009026f
C333 B.n180 VSUBS 0.009026f
C334 B.n181 VSUBS 0.009026f
C335 B.n182 VSUBS 0.009026f
C336 B.n183 VSUBS 0.009026f
C337 B.n184 VSUBS 0.009026f
C338 B.n185 VSUBS 0.009026f
C339 B.n186 VSUBS 0.009026f
C340 B.n187 VSUBS 0.008495f
C341 B.n188 VSUBS 0.020913f
C342 B.n189 VSUBS 0.005044f
C343 B.n190 VSUBS 0.009026f
C344 B.n191 VSUBS 0.009026f
C345 B.n192 VSUBS 0.009026f
C346 B.n193 VSUBS 0.009026f
C347 B.n194 VSUBS 0.009026f
C348 B.n195 VSUBS 0.009026f
C349 B.n196 VSUBS 0.009026f
C350 B.n197 VSUBS 0.009026f
C351 B.n198 VSUBS 0.009026f
C352 B.n199 VSUBS 0.009026f
C353 B.n200 VSUBS 0.009026f
C354 B.n201 VSUBS 0.009026f
C355 B.n202 VSUBS 0.005044f
C356 B.n203 VSUBS 0.009026f
C357 B.n204 VSUBS 0.009026f
C358 B.n205 VSUBS 0.008495f
C359 B.n206 VSUBS 0.009026f
C360 B.n207 VSUBS 0.009026f
C361 B.n208 VSUBS 0.009026f
C362 B.n209 VSUBS 0.009026f
C363 B.n210 VSUBS 0.009026f
C364 B.n211 VSUBS 0.009026f
C365 B.n212 VSUBS 0.009026f
C366 B.n213 VSUBS 0.009026f
C367 B.n214 VSUBS 0.009026f
C368 B.n215 VSUBS 0.009026f
C369 B.n216 VSUBS 0.009026f
C370 B.n217 VSUBS 0.009026f
C371 B.n218 VSUBS 0.009026f
C372 B.n219 VSUBS 0.009026f
C373 B.n220 VSUBS 0.009026f
C374 B.n221 VSUBS 0.009026f
C375 B.n222 VSUBS 0.009026f
C376 B.n223 VSUBS 0.009026f
C377 B.n224 VSUBS 0.009026f
C378 B.n225 VSUBS 0.009026f
C379 B.n226 VSUBS 0.009026f
C380 B.n227 VSUBS 0.009026f
C381 B.n228 VSUBS 0.009026f
C382 B.n229 VSUBS 0.009026f
C383 B.n230 VSUBS 0.009026f
C384 B.n231 VSUBS 0.009026f
C385 B.n232 VSUBS 0.009026f
C386 B.n233 VSUBS 0.009026f
C387 B.n234 VSUBS 0.009026f
C388 B.n235 VSUBS 0.009026f
C389 B.n236 VSUBS 0.009026f
C390 B.n237 VSUBS 0.009026f
C391 B.n238 VSUBS 0.009026f
C392 B.n239 VSUBS 0.009026f
C393 B.n240 VSUBS 0.009026f
C394 B.n241 VSUBS 0.009026f
C395 B.n242 VSUBS 0.009026f
C396 B.n243 VSUBS 0.009026f
C397 B.n244 VSUBS 0.009026f
C398 B.n245 VSUBS 0.009026f
C399 B.n246 VSUBS 0.009026f
C400 B.n247 VSUBS 0.009026f
C401 B.n248 VSUBS 0.021275f
C402 B.n249 VSUBS 0.020936f
C403 B.n250 VSUBS 0.020936f
C404 B.n251 VSUBS 0.009026f
C405 B.n252 VSUBS 0.009026f
C406 B.n253 VSUBS 0.009026f
C407 B.n254 VSUBS 0.009026f
C408 B.n255 VSUBS 0.009026f
C409 B.n256 VSUBS 0.009026f
C410 B.n257 VSUBS 0.009026f
C411 B.n258 VSUBS 0.009026f
C412 B.n259 VSUBS 0.009026f
C413 B.n260 VSUBS 0.009026f
C414 B.n261 VSUBS 0.009026f
C415 B.n262 VSUBS 0.009026f
C416 B.n263 VSUBS 0.009026f
C417 B.n264 VSUBS 0.009026f
C418 B.n265 VSUBS 0.009026f
C419 B.n266 VSUBS 0.009026f
C420 B.n267 VSUBS 0.009026f
C421 B.n268 VSUBS 0.009026f
C422 B.n269 VSUBS 0.009026f
C423 B.n270 VSUBS 0.009026f
C424 B.n271 VSUBS 0.009026f
C425 B.n272 VSUBS 0.009026f
C426 B.n273 VSUBS 0.009026f
C427 B.n274 VSUBS 0.009026f
C428 B.n275 VSUBS 0.009026f
C429 B.n276 VSUBS 0.009026f
C430 B.n277 VSUBS 0.009026f
C431 B.n278 VSUBS 0.009026f
C432 B.n279 VSUBS 0.009026f
C433 B.n280 VSUBS 0.009026f
C434 B.n281 VSUBS 0.009026f
C435 B.n282 VSUBS 0.009026f
C436 B.n283 VSUBS 0.009026f
C437 B.n284 VSUBS 0.009026f
C438 B.n285 VSUBS 0.009026f
C439 B.n286 VSUBS 0.009026f
C440 B.n287 VSUBS 0.009026f
C441 B.n288 VSUBS 0.009026f
C442 B.n289 VSUBS 0.009026f
C443 B.n290 VSUBS 0.009026f
C444 B.n291 VSUBS 0.009026f
C445 B.n292 VSUBS 0.009026f
C446 B.n293 VSUBS 0.009026f
C447 B.n294 VSUBS 0.009026f
C448 B.n295 VSUBS 0.009026f
C449 B.n296 VSUBS 0.009026f
C450 B.n297 VSUBS 0.009026f
C451 B.n298 VSUBS 0.009026f
C452 B.n299 VSUBS 0.009026f
C453 B.n300 VSUBS 0.009026f
C454 B.n301 VSUBS 0.009026f
C455 B.n302 VSUBS 0.009026f
C456 B.n303 VSUBS 0.022004f
C457 B.n304 VSUBS 0.020936f
C458 B.n305 VSUBS 0.021275f
C459 B.n306 VSUBS 0.009026f
C460 B.n307 VSUBS 0.009026f
C461 B.n308 VSUBS 0.009026f
C462 B.n309 VSUBS 0.009026f
C463 B.n310 VSUBS 0.009026f
C464 B.n311 VSUBS 0.009026f
C465 B.n312 VSUBS 0.009026f
C466 B.n313 VSUBS 0.009026f
C467 B.n314 VSUBS 0.009026f
C468 B.n315 VSUBS 0.009026f
C469 B.n316 VSUBS 0.009026f
C470 B.n317 VSUBS 0.009026f
C471 B.n318 VSUBS 0.009026f
C472 B.n319 VSUBS 0.009026f
C473 B.n320 VSUBS 0.009026f
C474 B.n321 VSUBS 0.009026f
C475 B.n322 VSUBS 0.009026f
C476 B.n323 VSUBS 0.009026f
C477 B.n324 VSUBS 0.009026f
C478 B.n325 VSUBS 0.009026f
C479 B.n326 VSUBS 0.009026f
C480 B.n327 VSUBS 0.009026f
C481 B.n328 VSUBS 0.009026f
C482 B.n329 VSUBS 0.009026f
C483 B.n330 VSUBS 0.009026f
C484 B.n331 VSUBS 0.009026f
C485 B.n332 VSUBS 0.009026f
C486 B.n333 VSUBS 0.009026f
C487 B.n334 VSUBS 0.009026f
C488 B.n335 VSUBS 0.009026f
C489 B.n336 VSUBS 0.009026f
C490 B.n337 VSUBS 0.009026f
C491 B.n338 VSUBS 0.009026f
C492 B.n339 VSUBS 0.009026f
C493 B.n340 VSUBS 0.009026f
C494 B.n341 VSUBS 0.009026f
C495 B.n342 VSUBS 0.009026f
C496 B.n343 VSUBS 0.009026f
C497 B.n344 VSUBS 0.009026f
C498 B.n345 VSUBS 0.009026f
C499 B.n346 VSUBS 0.009026f
C500 B.n347 VSUBS 0.009026f
C501 B.n348 VSUBS 0.009026f
C502 B.n349 VSUBS 0.008495f
C503 B.n350 VSUBS 0.020913f
C504 B.n351 VSUBS 0.005044f
C505 B.n352 VSUBS 0.009026f
C506 B.n353 VSUBS 0.009026f
C507 B.n354 VSUBS 0.009026f
C508 B.n355 VSUBS 0.009026f
C509 B.n356 VSUBS 0.009026f
C510 B.n357 VSUBS 0.009026f
C511 B.n358 VSUBS 0.009026f
C512 B.n359 VSUBS 0.009026f
C513 B.n360 VSUBS 0.009026f
C514 B.n361 VSUBS 0.009026f
C515 B.n362 VSUBS 0.009026f
C516 B.n363 VSUBS 0.009026f
C517 B.n364 VSUBS 0.005044f
C518 B.n365 VSUBS 0.009026f
C519 B.n366 VSUBS 0.009026f
C520 B.n367 VSUBS 0.008495f
C521 B.n368 VSUBS 0.009026f
C522 B.n369 VSUBS 0.009026f
C523 B.n370 VSUBS 0.009026f
C524 B.n371 VSUBS 0.009026f
C525 B.n372 VSUBS 0.009026f
C526 B.n373 VSUBS 0.009026f
C527 B.n374 VSUBS 0.009026f
C528 B.n375 VSUBS 0.009026f
C529 B.n376 VSUBS 0.009026f
C530 B.n377 VSUBS 0.009026f
C531 B.n378 VSUBS 0.009026f
C532 B.n379 VSUBS 0.009026f
C533 B.n380 VSUBS 0.009026f
C534 B.n381 VSUBS 0.009026f
C535 B.n382 VSUBS 0.009026f
C536 B.n383 VSUBS 0.009026f
C537 B.n384 VSUBS 0.009026f
C538 B.n385 VSUBS 0.009026f
C539 B.n386 VSUBS 0.009026f
C540 B.n387 VSUBS 0.009026f
C541 B.n388 VSUBS 0.009026f
C542 B.n389 VSUBS 0.009026f
C543 B.n390 VSUBS 0.009026f
C544 B.n391 VSUBS 0.009026f
C545 B.n392 VSUBS 0.009026f
C546 B.n393 VSUBS 0.009026f
C547 B.n394 VSUBS 0.009026f
C548 B.n395 VSUBS 0.009026f
C549 B.n396 VSUBS 0.009026f
C550 B.n397 VSUBS 0.009026f
C551 B.n398 VSUBS 0.009026f
C552 B.n399 VSUBS 0.009026f
C553 B.n400 VSUBS 0.009026f
C554 B.n401 VSUBS 0.009026f
C555 B.n402 VSUBS 0.009026f
C556 B.n403 VSUBS 0.009026f
C557 B.n404 VSUBS 0.009026f
C558 B.n405 VSUBS 0.009026f
C559 B.n406 VSUBS 0.009026f
C560 B.n407 VSUBS 0.009026f
C561 B.n408 VSUBS 0.009026f
C562 B.n409 VSUBS 0.009026f
C563 B.n410 VSUBS 0.021275f
C564 B.n411 VSUBS 0.020936f
C565 B.n412 VSUBS 0.020936f
C566 B.n413 VSUBS 0.009026f
C567 B.n414 VSUBS 0.009026f
C568 B.n415 VSUBS 0.009026f
C569 B.n416 VSUBS 0.009026f
C570 B.n417 VSUBS 0.009026f
C571 B.n418 VSUBS 0.009026f
C572 B.n419 VSUBS 0.009026f
C573 B.n420 VSUBS 0.009026f
C574 B.n421 VSUBS 0.009026f
C575 B.n422 VSUBS 0.009026f
C576 B.n423 VSUBS 0.009026f
C577 B.n424 VSUBS 0.009026f
C578 B.n425 VSUBS 0.009026f
C579 B.n426 VSUBS 0.009026f
C580 B.n427 VSUBS 0.009026f
C581 B.n428 VSUBS 0.009026f
C582 B.n429 VSUBS 0.009026f
C583 B.n430 VSUBS 0.009026f
C584 B.n431 VSUBS 0.009026f
C585 B.n432 VSUBS 0.009026f
C586 B.n433 VSUBS 0.009026f
C587 B.n434 VSUBS 0.009026f
C588 B.n435 VSUBS 0.009026f
C589 B.n436 VSUBS 0.009026f
C590 B.n437 VSUBS 0.009026f
C591 B.n438 VSUBS 0.009026f
C592 B.n439 VSUBS 0.020439f
.ends

