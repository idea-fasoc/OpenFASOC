* NGSPICE file created from diff_pair_sample_0511.ext - technology: sky130A

.subckt diff_pair_sample_0511 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=4.017 ps=21.38 w=10.3 l=2.9
X1 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=4.017 pd=21.38 as=0 ps=0 w=10.3 l=2.9
X2 VDD1.t4 VP.t1 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=4.017 pd=21.38 as=1.6995 ps=10.63 w=10.3 l=2.9
X3 VDD2.t5 VN.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=4.017 pd=21.38 as=1.6995 ps=10.63 w=10.3 l=2.9
X4 VDD1.t3 VP.t2 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=4.017 pd=21.38 as=1.6995 ps=10.63 w=10.3 l=2.9
X5 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=4.017 pd=21.38 as=0 ps=0 w=10.3 l=2.9
X6 VTAIL.t9 VP.t3 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=1.6995 ps=10.63 w=10.3 l=2.9
X7 VDD2.t4 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=4.017 pd=21.38 as=1.6995 ps=10.63 w=10.3 l=2.9
X8 VDD2.t3 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=4.017 ps=21.38 w=10.3 l=2.9
X9 VDD1.t1 VP.t4 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=4.017 ps=21.38 w=10.3 l=2.9
X10 VDD2.t2 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=4.017 ps=21.38 w=10.3 l=2.9
X11 VTAIL.t7 VP.t5 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=1.6995 ps=10.63 w=10.3 l=2.9
X12 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=4.017 pd=21.38 as=0 ps=0 w=10.3 l=2.9
X13 VTAIL.t5 VN.t4 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=1.6995 ps=10.63 w=10.3 l=2.9
X14 VTAIL.t1 VN.t5 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6995 pd=10.63 as=1.6995 ps=10.63 w=10.3 l=2.9
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.017 pd=21.38 as=0 ps=0 w=10.3 l=2.9
R0 VP.n13 VP.n10 161.3
R1 VP.n15 VP.n14 161.3
R2 VP.n16 VP.n9 161.3
R3 VP.n18 VP.n17 161.3
R4 VP.n19 VP.n8 161.3
R5 VP.n21 VP.n20 161.3
R6 VP.n43 VP.n42 161.3
R7 VP.n41 VP.n1 161.3
R8 VP.n40 VP.n39 161.3
R9 VP.n38 VP.n2 161.3
R10 VP.n37 VP.n36 161.3
R11 VP.n35 VP.n3 161.3
R12 VP.n33 VP.n32 161.3
R13 VP.n31 VP.n4 161.3
R14 VP.n30 VP.n29 161.3
R15 VP.n28 VP.n5 161.3
R16 VP.n27 VP.n26 161.3
R17 VP.n25 VP.n6 161.3
R18 VP.n11 VP.t1 117.368
R19 VP.n23 VP.t2 85.5971
R20 VP.n34 VP.t5 85.5971
R21 VP.n0 VP.t0 85.5971
R22 VP.n7 VP.t4 85.5971
R23 VP.n12 VP.t3 85.5971
R24 VP.n24 VP.n23 66.5213
R25 VP.n44 VP.n0 66.5213
R26 VP.n22 VP.n7 66.5213
R27 VP.n12 VP.n11 61.4167
R28 VP.n29 VP.n28 53.5561
R29 VP.n40 VP.n2 53.5561
R30 VP.n18 VP.n9 53.5561
R31 VP.n24 VP.n22 48.715
R32 VP.n28 VP.n27 27.2651
R33 VP.n41 VP.n40 27.2651
R34 VP.n19 VP.n18 27.2651
R35 VP.n27 VP.n6 24.3439
R36 VP.n29 VP.n4 24.3439
R37 VP.n33 VP.n4 24.3439
R38 VP.n36 VP.n35 24.3439
R39 VP.n36 VP.n2 24.3439
R40 VP.n42 VP.n41 24.3439
R41 VP.n20 VP.n19 24.3439
R42 VP.n14 VP.n13 24.3439
R43 VP.n14 VP.n9 24.3439
R44 VP.n23 VP.n6 23.3702
R45 VP.n42 VP.n0 23.3702
R46 VP.n20 VP.n7 23.3702
R47 VP.n34 VP.n33 12.1722
R48 VP.n35 VP.n34 12.1722
R49 VP.n13 VP.n12 12.1722
R50 VP.n11 VP.n10 5.30778
R51 VP.n22 VP.n21 0.355081
R52 VP.n25 VP.n24 0.355081
R53 VP.n44 VP.n43 0.355081
R54 VP VP.n44 0.26685
R55 VP.n15 VP.n10 0.189894
R56 VP.n16 VP.n15 0.189894
R57 VP.n17 VP.n16 0.189894
R58 VP.n17 VP.n8 0.189894
R59 VP.n21 VP.n8 0.189894
R60 VP.n26 VP.n25 0.189894
R61 VP.n26 VP.n5 0.189894
R62 VP.n30 VP.n5 0.189894
R63 VP.n31 VP.n30 0.189894
R64 VP.n32 VP.n31 0.189894
R65 VP.n32 VP.n3 0.189894
R66 VP.n37 VP.n3 0.189894
R67 VP.n38 VP.n37 0.189894
R68 VP.n39 VP.n38 0.189894
R69 VP.n39 VP.n1 0.189894
R70 VP.n43 VP.n1 0.189894
R71 VTAIL.n7 VTAIL.t0 47.3387
R72 VTAIL.n11 VTAIL.t3 47.3384
R73 VTAIL.n2 VTAIL.t10 47.3384
R74 VTAIL.n10 VTAIL.t8 47.3384
R75 VTAIL.n9 VTAIL.n8 45.4163
R76 VTAIL.n6 VTAIL.n5 45.4163
R77 VTAIL.n1 VTAIL.n0 45.4161
R78 VTAIL.n4 VTAIL.n3 45.4161
R79 VTAIL.n6 VTAIL.n4 26.8152
R80 VTAIL.n11 VTAIL.n10 24.0307
R81 VTAIL.n7 VTAIL.n6 2.78498
R82 VTAIL.n10 VTAIL.n9 2.78498
R83 VTAIL.n4 VTAIL.n2 2.78498
R84 VTAIL VTAIL.n11 2.03067
R85 VTAIL.n0 VTAIL.t4 1.92283
R86 VTAIL.n0 VTAIL.t1 1.92283
R87 VTAIL.n3 VTAIL.t11 1.92283
R88 VTAIL.n3 VTAIL.t7 1.92283
R89 VTAIL.n8 VTAIL.t6 1.92283
R90 VTAIL.n8 VTAIL.t9 1.92283
R91 VTAIL.n5 VTAIL.t2 1.92283
R92 VTAIL.n5 VTAIL.t5 1.92283
R93 VTAIL.n9 VTAIL.n7 1.86257
R94 VTAIL.n2 VTAIL.n1 1.86257
R95 VTAIL VTAIL.n1 0.75481
R96 VDD1 VDD1.t4 66.164
R97 VDD1.n1 VDD1.t3 66.0502
R98 VDD1.n1 VDD1.n0 62.7357
R99 VDD1.n3 VDD1.n2 62.0949
R100 VDD1.n3 VDD1.n1 43.6194
R101 VDD1.n2 VDD1.t2 1.92283
R102 VDD1.n2 VDD1.t1 1.92283
R103 VDD1.n0 VDD1.t0 1.92283
R104 VDD1.n0 VDD1.t5 1.92283
R105 VDD1 VDD1.n3 0.638431
R106 B.n632 B.n132 585
R107 B.n132 B.n85 585
R108 B.n634 B.n633 585
R109 B.n636 B.n131 585
R110 B.n639 B.n638 585
R111 B.n640 B.n130 585
R112 B.n642 B.n641 585
R113 B.n644 B.n129 585
R114 B.n647 B.n646 585
R115 B.n648 B.n128 585
R116 B.n650 B.n649 585
R117 B.n652 B.n127 585
R118 B.n655 B.n654 585
R119 B.n656 B.n126 585
R120 B.n658 B.n657 585
R121 B.n660 B.n125 585
R122 B.n663 B.n662 585
R123 B.n664 B.n124 585
R124 B.n666 B.n665 585
R125 B.n668 B.n123 585
R126 B.n671 B.n670 585
R127 B.n672 B.n122 585
R128 B.n674 B.n673 585
R129 B.n676 B.n121 585
R130 B.n679 B.n678 585
R131 B.n680 B.n120 585
R132 B.n682 B.n681 585
R133 B.n684 B.n119 585
R134 B.n687 B.n686 585
R135 B.n688 B.n118 585
R136 B.n690 B.n689 585
R137 B.n692 B.n117 585
R138 B.n695 B.n694 585
R139 B.n696 B.n116 585
R140 B.n698 B.n697 585
R141 B.n700 B.n115 585
R142 B.n702 B.n701 585
R143 B.n704 B.n703 585
R144 B.n707 B.n706 585
R145 B.n708 B.n110 585
R146 B.n710 B.n709 585
R147 B.n712 B.n109 585
R148 B.n715 B.n714 585
R149 B.n716 B.n108 585
R150 B.n718 B.n717 585
R151 B.n720 B.n107 585
R152 B.n723 B.n722 585
R153 B.n725 B.n104 585
R154 B.n727 B.n726 585
R155 B.n729 B.n103 585
R156 B.n732 B.n731 585
R157 B.n733 B.n102 585
R158 B.n735 B.n734 585
R159 B.n737 B.n101 585
R160 B.n740 B.n739 585
R161 B.n741 B.n100 585
R162 B.n743 B.n742 585
R163 B.n745 B.n99 585
R164 B.n748 B.n747 585
R165 B.n749 B.n98 585
R166 B.n751 B.n750 585
R167 B.n753 B.n97 585
R168 B.n756 B.n755 585
R169 B.n757 B.n96 585
R170 B.n759 B.n758 585
R171 B.n761 B.n95 585
R172 B.n764 B.n763 585
R173 B.n765 B.n94 585
R174 B.n767 B.n766 585
R175 B.n769 B.n93 585
R176 B.n772 B.n771 585
R177 B.n773 B.n92 585
R178 B.n775 B.n774 585
R179 B.n777 B.n91 585
R180 B.n780 B.n779 585
R181 B.n781 B.n90 585
R182 B.n783 B.n782 585
R183 B.n785 B.n89 585
R184 B.n788 B.n787 585
R185 B.n789 B.n88 585
R186 B.n791 B.n790 585
R187 B.n793 B.n87 585
R188 B.n796 B.n795 585
R189 B.n797 B.n86 585
R190 B.n631 B.n84 585
R191 B.n800 B.n84 585
R192 B.n630 B.n83 585
R193 B.n801 B.n83 585
R194 B.n629 B.n82 585
R195 B.n802 B.n82 585
R196 B.n628 B.n627 585
R197 B.n627 B.n78 585
R198 B.n626 B.n77 585
R199 B.n808 B.n77 585
R200 B.n625 B.n76 585
R201 B.n809 B.n76 585
R202 B.n624 B.n75 585
R203 B.n810 B.n75 585
R204 B.n623 B.n622 585
R205 B.n622 B.n74 585
R206 B.n621 B.n70 585
R207 B.n816 B.n70 585
R208 B.n620 B.n69 585
R209 B.n817 B.n69 585
R210 B.n619 B.n68 585
R211 B.n818 B.n68 585
R212 B.n618 B.n617 585
R213 B.n617 B.n64 585
R214 B.n616 B.n63 585
R215 B.n824 B.n63 585
R216 B.n615 B.n62 585
R217 B.n825 B.n62 585
R218 B.n614 B.n61 585
R219 B.n826 B.n61 585
R220 B.n613 B.n612 585
R221 B.n612 B.n57 585
R222 B.n611 B.n56 585
R223 B.n832 B.n56 585
R224 B.n610 B.n55 585
R225 B.n833 B.n55 585
R226 B.n609 B.n54 585
R227 B.n834 B.n54 585
R228 B.n608 B.n607 585
R229 B.n607 B.n50 585
R230 B.n606 B.n49 585
R231 B.n840 B.n49 585
R232 B.n605 B.n48 585
R233 B.n841 B.n48 585
R234 B.n604 B.n47 585
R235 B.n842 B.n47 585
R236 B.n603 B.n602 585
R237 B.n602 B.n43 585
R238 B.n601 B.n42 585
R239 B.n848 B.n42 585
R240 B.n600 B.n41 585
R241 B.n849 B.n41 585
R242 B.n599 B.n40 585
R243 B.n850 B.n40 585
R244 B.n598 B.n597 585
R245 B.n597 B.n36 585
R246 B.n596 B.n35 585
R247 B.n856 B.n35 585
R248 B.n595 B.n34 585
R249 B.n857 B.n34 585
R250 B.n594 B.n33 585
R251 B.n858 B.n33 585
R252 B.n593 B.n592 585
R253 B.n592 B.n29 585
R254 B.n591 B.n28 585
R255 B.n864 B.n28 585
R256 B.n590 B.n27 585
R257 B.n865 B.n27 585
R258 B.n589 B.n26 585
R259 B.n866 B.n26 585
R260 B.n588 B.n587 585
R261 B.n587 B.n22 585
R262 B.n586 B.n21 585
R263 B.n872 B.n21 585
R264 B.n585 B.n20 585
R265 B.n873 B.n20 585
R266 B.n584 B.n19 585
R267 B.n874 B.n19 585
R268 B.n583 B.n582 585
R269 B.n582 B.n18 585
R270 B.n581 B.n14 585
R271 B.n880 B.n14 585
R272 B.n580 B.n13 585
R273 B.n881 B.n13 585
R274 B.n579 B.n12 585
R275 B.n882 B.n12 585
R276 B.n578 B.n577 585
R277 B.n577 B.n8 585
R278 B.n576 B.n7 585
R279 B.n888 B.n7 585
R280 B.n575 B.n6 585
R281 B.n889 B.n6 585
R282 B.n574 B.n5 585
R283 B.n890 B.n5 585
R284 B.n573 B.n572 585
R285 B.n572 B.n4 585
R286 B.n571 B.n133 585
R287 B.n571 B.n570 585
R288 B.n561 B.n134 585
R289 B.n135 B.n134 585
R290 B.n563 B.n562 585
R291 B.n564 B.n563 585
R292 B.n560 B.n140 585
R293 B.n140 B.n139 585
R294 B.n559 B.n558 585
R295 B.n558 B.n557 585
R296 B.n142 B.n141 585
R297 B.n550 B.n142 585
R298 B.n549 B.n548 585
R299 B.n551 B.n549 585
R300 B.n547 B.n147 585
R301 B.n147 B.n146 585
R302 B.n546 B.n545 585
R303 B.n545 B.n544 585
R304 B.n149 B.n148 585
R305 B.n150 B.n149 585
R306 B.n537 B.n536 585
R307 B.n538 B.n537 585
R308 B.n535 B.n155 585
R309 B.n155 B.n154 585
R310 B.n534 B.n533 585
R311 B.n533 B.n532 585
R312 B.n157 B.n156 585
R313 B.n158 B.n157 585
R314 B.n525 B.n524 585
R315 B.n526 B.n525 585
R316 B.n523 B.n163 585
R317 B.n163 B.n162 585
R318 B.n522 B.n521 585
R319 B.n521 B.n520 585
R320 B.n165 B.n164 585
R321 B.n166 B.n165 585
R322 B.n513 B.n512 585
R323 B.n514 B.n513 585
R324 B.n511 B.n171 585
R325 B.n171 B.n170 585
R326 B.n510 B.n509 585
R327 B.n509 B.n508 585
R328 B.n173 B.n172 585
R329 B.n174 B.n173 585
R330 B.n501 B.n500 585
R331 B.n502 B.n501 585
R332 B.n499 B.n179 585
R333 B.n179 B.n178 585
R334 B.n498 B.n497 585
R335 B.n497 B.n496 585
R336 B.n181 B.n180 585
R337 B.n182 B.n181 585
R338 B.n489 B.n488 585
R339 B.n490 B.n489 585
R340 B.n487 B.n187 585
R341 B.n187 B.n186 585
R342 B.n486 B.n485 585
R343 B.n485 B.n484 585
R344 B.n189 B.n188 585
R345 B.n190 B.n189 585
R346 B.n477 B.n476 585
R347 B.n478 B.n477 585
R348 B.n475 B.n195 585
R349 B.n195 B.n194 585
R350 B.n474 B.n473 585
R351 B.n473 B.n472 585
R352 B.n197 B.n196 585
R353 B.n198 B.n197 585
R354 B.n465 B.n464 585
R355 B.n466 B.n465 585
R356 B.n463 B.n203 585
R357 B.n203 B.n202 585
R358 B.n462 B.n461 585
R359 B.n461 B.n460 585
R360 B.n205 B.n204 585
R361 B.n453 B.n205 585
R362 B.n452 B.n451 585
R363 B.n454 B.n452 585
R364 B.n450 B.n210 585
R365 B.n210 B.n209 585
R366 B.n449 B.n448 585
R367 B.n448 B.n447 585
R368 B.n212 B.n211 585
R369 B.n213 B.n212 585
R370 B.n440 B.n439 585
R371 B.n441 B.n440 585
R372 B.n438 B.n218 585
R373 B.n218 B.n217 585
R374 B.n437 B.n436 585
R375 B.n436 B.n435 585
R376 B.n432 B.n222 585
R377 B.n431 B.n430 585
R378 B.n428 B.n223 585
R379 B.n428 B.n221 585
R380 B.n427 B.n426 585
R381 B.n425 B.n424 585
R382 B.n423 B.n225 585
R383 B.n421 B.n420 585
R384 B.n419 B.n226 585
R385 B.n418 B.n417 585
R386 B.n415 B.n227 585
R387 B.n413 B.n412 585
R388 B.n411 B.n228 585
R389 B.n410 B.n409 585
R390 B.n407 B.n229 585
R391 B.n405 B.n404 585
R392 B.n403 B.n230 585
R393 B.n402 B.n401 585
R394 B.n399 B.n231 585
R395 B.n397 B.n396 585
R396 B.n395 B.n232 585
R397 B.n394 B.n393 585
R398 B.n391 B.n233 585
R399 B.n389 B.n388 585
R400 B.n387 B.n234 585
R401 B.n386 B.n385 585
R402 B.n383 B.n235 585
R403 B.n381 B.n380 585
R404 B.n379 B.n236 585
R405 B.n378 B.n377 585
R406 B.n375 B.n237 585
R407 B.n373 B.n372 585
R408 B.n371 B.n238 585
R409 B.n370 B.n369 585
R410 B.n367 B.n239 585
R411 B.n365 B.n364 585
R412 B.n363 B.n240 585
R413 B.n362 B.n361 585
R414 B.n359 B.n358 585
R415 B.n357 B.n356 585
R416 B.n355 B.n245 585
R417 B.n353 B.n352 585
R418 B.n351 B.n246 585
R419 B.n350 B.n349 585
R420 B.n347 B.n247 585
R421 B.n345 B.n344 585
R422 B.n343 B.n248 585
R423 B.n341 B.n340 585
R424 B.n338 B.n251 585
R425 B.n336 B.n335 585
R426 B.n334 B.n252 585
R427 B.n333 B.n332 585
R428 B.n330 B.n253 585
R429 B.n328 B.n327 585
R430 B.n326 B.n254 585
R431 B.n325 B.n324 585
R432 B.n322 B.n255 585
R433 B.n320 B.n319 585
R434 B.n318 B.n256 585
R435 B.n317 B.n316 585
R436 B.n314 B.n257 585
R437 B.n312 B.n311 585
R438 B.n310 B.n258 585
R439 B.n309 B.n308 585
R440 B.n306 B.n259 585
R441 B.n304 B.n303 585
R442 B.n302 B.n260 585
R443 B.n301 B.n300 585
R444 B.n298 B.n261 585
R445 B.n296 B.n295 585
R446 B.n294 B.n262 585
R447 B.n293 B.n292 585
R448 B.n290 B.n263 585
R449 B.n288 B.n287 585
R450 B.n286 B.n264 585
R451 B.n285 B.n284 585
R452 B.n282 B.n265 585
R453 B.n280 B.n279 585
R454 B.n278 B.n266 585
R455 B.n277 B.n276 585
R456 B.n274 B.n267 585
R457 B.n272 B.n271 585
R458 B.n270 B.n269 585
R459 B.n220 B.n219 585
R460 B.n434 B.n433 585
R461 B.n435 B.n434 585
R462 B.n216 B.n215 585
R463 B.n217 B.n216 585
R464 B.n443 B.n442 585
R465 B.n442 B.n441 585
R466 B.n444 B.n214 585
R467 B.n214 B.n213 585
R468 B.n446 B.n445 585
R469 B.n447 B.n446 585
R470 B.n208 B.n207 585
R471 B.n209 B.n208 585
R472 B.n456 B.n455 585
R473 B.n455 B.n454 585
R474 B.n457 B.n206 585
R475 B.n453 B.n206 585
R476 B.n459 B.n458 585
R477 B.n460 B.n459 585
R478 B.n201 B.n200 585
R479 B.n202 B.n201 585
R480 B.n468 B.n467 585
R481 B.n467 B.n466 585
R482 B.n469 B.n199 585
R483 B.n199 B.n198 585
R484 B.n471 B.n470 585
R485 B.n472 B.n471 585
R486 B.n193 B.n192 585
R487 B.n194 B.n193 585
R488 B.n480 B.n479 585
R489 B.n479 B.n478 585
R490 B.n481 B.n191 585
R491 B.n191 B.n190 585
R492 B.n483 B.n482 585
R493 B.n484 B.n483 585
R494 B.n185 B.n184 585
R495 B.n186 B.n185 585
R496 B.n492 B.n491 585
R497 B.n491 B.n490 585
R498 B.n493 B.n183 585
R499 B.n183 B.n182 585
R500 B.n495 B.n494 585
R501 B.n496 B.n495 585
R502 B.n177 B.n176 585
R503 B.n178 B.n177 585
R504 B.n504 B.n503 585
R505 B.n503 B.n502 585
R506 B.n505 B.n175 585
R507 B.n175 B.n174 585
R508 B.n507 B.n506 585
R509 B.n508 B.n507 585
R510 B.n169 B.n168 585
R511 B.n170 B.n169 585
R512 B.n516 B.n515 585
R513 B.n515 B.n514 585
R514 B.n517 B.n167 585
R515 B.n167 B.n166 585
R516 B.n519 B.n518 585
R517 B.n520 B.n519 585
R518 B.n161 B.n160 585
R519 B.n162 B.n161 585
R520 B.n528 B.n527 585
R521 B.n527 B.n526 585
R522 B.n529 B.n159 585
R523 B.n159 B.n158 585
R524 B.n531 B.n530 585
R525 B.n532 B.n531 585
R526 B.n153 B.n152 585
R527 B.n154 B.n153 585
R528 B.n540 B.n539 585
R529 B.n539 B.n538 585
R530 B.n541 B.n151 585
R531 B.n151 B.n150 585
R532 B.n543 B.n542 585
R533 B.n544 B.n543 585
R534 B.n145 B.n144 585
R535 B.n146 B.n145 585
R536 B.n553 B.n552 585
R537 B.n552 B.n551 585
R538 B.n554 B.n143 585
R539 B.n550 B.n143 585
R540 B.n556 B.n555 585
R541 B.n557 B.n556 585
R542 B.n138 B.n137 585
R543 B.n139 B.n138 585
R544 B.n566 B.n565 585
R545 B.n565 B.n564 585
R546 B.n567 B.n136 585
R547 B.n136 B.n135 585
R548 B.n569 B.n568 585
R549 B.n570 B.n569 585
R550 B.n2 B.n0 585
R551 B.n4 B.n2 585
R552 B.n3 B.n1 585
R553 B.n889 B.n3 585
R554 B.n887 B.n886 585
R555 B.n888 B.n887 585
R556 B.n885 B.n9 585
R557 B.n9 B.n8 585
R558 B.n884 B.n883 585
R559 B.n883 B.n882 585
R560 B.n11 B.n10 585
R561 B.n881 B.n11 585
R562 B.n879 B.n878 585
R563 B.n880 B.n879 585
R564 B.n877 B.n15 585
R565 B.n18 B.n15 585
R566 B.n876 B.n875 585
R567 B.n875 B.n874 585
R568 B.n17 B.n16 585
R569 B.n873 B.n17 585
R570 B.n871 B.n870 585
R571 B.n872 B.n871 585
R572 B.n869 B.n23 585
R573 B.n23 B.n22 585
R574 B.n868 B.n867 585
R575 B.n867 B.n866 585
R576 B.n25 B.n24 585
R577 B.n865 B.n25 585
R578 B.n863 B.n862 585
R579 B.n864 B.n863 585
R580 B.n861 B.n30 585
R581 B.n30 B.n29 585
R582 B.n860 B.n859 585
R583 B.n859 B.n858 585
R584 B.n32 B.n31 585
R585 B.n857 B.n32 585
R586 B.n855 B.n854 585
R587 B.n856 B.n855 585
R588 B.n853 B.n37 585
R589 B.n37 B.n36 585
R590 B.n852 B.n851 585
R591 B.n851 B.n850 585
R592 B.n39 B.n38 585
R593 B.n849 B.n39 585
R594 B.n847 B.n846 585
R595 B.n848 B.n847 585
R596 B.n845 B.n44 585
R597 B.n44 B.n43 585
R598 B.n844 B.n843 585
R599 B.n843 B.n842 585
R600 B.n46 B.n45 585
R601 B.n841 B.n46 585
R602 B.n839 B.n838 585
R603 B.n840 B.n839 585
R604 B.n837 B.n51 585
R605 B.n51 B.n50 585
R606 B.n836 B.n835 585
R607 B.n835 B.n834 585
R608 B.n53 B.n52 585
R609 B.n833 B.n53 585
R610 B.n831 B.n830 585
R611 B.n832 B.n831 585
R612 B.n829 B.n58 585
R613 B.n58 B.n57 585
R614 B.n828 B.n827 585
R615 B.n827 B.n826 585
R616 B.n60 B.n59 585
R617 B.n825 B.n60 585
R618 B.n823 B.n822 585
R619 B.n824 B.n823 585
R620 B.n821 B.n65 585
R621 B.n65 B.n64 585
R622 B.n820 B.n819 585
R623 B.n819 B.n818 585
R624 B.n67 B.n66 585
R625 B.n817 B.n67 585
R626 B.n815 B.n814 585
R627 B.n816 B.n815 585
R628 B.n813 B.n71 585
R629 B.n74 B.n71 585
R630 B.n812 B.n811 585
R631 B.n811 B.n810 585
R632 B.n73 B.n72 585
R633 B.n809 B.n73 585
R634 B.n807 B.n806 585
R635 B.n808 B.n807 585
R636 B.n805 B.n79 585
R637 B.n79 B.n78 585
R638 B.n804 B.n803 585
R639 B.n803 B.n802 585
R640 B.n81 B.n80 585
R641 B.n801 B.n81 585
R642 B.n799 B.n798 585
R643 B.n800 B.n799 585
R644 B.n892 B.n891 585
R645 B.n891 B.n890 585
R646 B.n434 B.n222 502.111
R647 B.n799 B.n86 502.111
R648 B.n436 B.n220 502.111
R649 B.n132 B.n84 502.111
R650 B.n249 B.t10 294.055
R651 B.n241 B.t6 294.055
R652 B.n105 B.t13 294.055
R653 B.n111 B.t17 294.055
R654 B.n635 B.n85 256.663
R655 B.n637 B.n85 256.663
R656 B.n643 B.n85 256.663
R657 B.n645 B.n85 256.663
R658 B.n651 B.n85 256.663
R659 B.n653 B.n85 256.663
R660 B.n659 B.n85 256.663
R661 B.n661 B.n85 256.663
R662 B.n667 B.n85 256.663
R663 B.n669 B.n85 256.663
R664 B.n675 B.n85 256.663
R665 B.n677 B.n85 256.663
R666 B.n683 B.n85 256.663
R667 B.n685 B.n85 256.663
R668 B.n691 B.n85 256.663
R669 B.n693 B.n85 256.663
R670 B.n699 B.n85 256.663
R671 B.n114 B.n85 256.663
R672 B.n705 B.n85 256.663
R673 B.n711 B.n85 256.663
R674 B.n713 B.n85 256.663
R675 B.n719 B.n85 256.663
R676 B.n721 B.n85 256.663
R677 B.n728 B.n85 256.663
R678 B.n730 B.n85 256.663
R679 B.n736 B.n85 256.663
R680 B.n738 B.n85 256.663
R681 B.n744 B.n85 256.663
R682 B.n746 B.n85 256.663
R683 B.n752 B.n85 256.663
R684 B.n754 B.n85 256.663
R685 B.n760 B.n85 256.663
R686 B.n762 B.n85 256.663
R687 B.n768 B.n85 256.663
R688 B.n770 B.n85 256.663
R689 B.n776 B.n85 256.663
R690 B.n778 B.n85 256.663
R691 B.n784 B.n85 256.663
R692 B.n786 B.n85 256.663
R693 B.n792 B.n85 256.663
R694 B.n794 B.n85 256.663
R695 B.n429 B.n221 256.663
R696 B.n224 B.n221 256.663
R697 B.n422 B.n221 256.663
R698 B.n416 B.n221 256.663
R699 B.n414 B.n221 256.663
R700 B.n408 B.n221 256.663
R701 B.n406 B.n221 256.663
R702 B.n400 B.n221 256.663
R703 B.n398 B.n221 256.663
R704 B.n392 B.n221 256.663
R705 B.n390 B.n221 256.663
R706 B.n384 B.n221 256.663
R707 B.n382 B.n221 256.663
R708 B.n376 B.n221 256.663
R709 B.n374 B.n221 256.663
R710 B.n368 B.n221 256.663
R711 B.n366 B.n221 256.663
R712 B.n360 B.n221 256.663
R713 B.n244 B.n221 256.663
R714 B.n354 B.n221 256.663
R715 B.n348 B.n221 256.663
R716 B.n346 B.n221 256.663
R717 B.n339 B.n221 256.663
R718 B.n337 B.n221 256.663
R719 B.n331 B.n221 256.663
R720 B.n329 B.n221 256.663
R721 B.n323 B.n221 256.663
R722 B.n321 B.n221 256.663
R723 B.n315 B.n221 256.663
R724 B.n313 B.n221 256.663
R725 B.n307 B.n221 256.663
R726 B.n305 B.n221 256.663
R727 B.n299 B.n221 256.663
R728 B.n297 B.n221 256.663
R729 B.n291 B.n221 256.663
R730 B.n289 B.n221 256.663
R731 B.n283 B.n221 256.663
R732 B.n281 B.n221 256.663
R733 B.n275 B.n221 256.663
R734 B.n273 B.n221 256.663
R735 B.n268 B.n221 256.663
R736 B.n434 B.n216 163.367
R737 B.n442 B.n216 163.367
R738 B.n442 B.n214 163.367
R739 B.n446 B.n214 163.367
R740 B.n446 B.n208 163.367
R741 B.n455 B.n208 163.367
R742 B.n455 B.n206 163.367
R743 B.n459 B.n206 163.367
R744 B.n459 B.n201 163.367
R745 B.n467 B.n201 163.367
R746 B.n467 B.n199 163.367
R747 B.n471 B.n199 163.367
R748 B.n471 B.n193 163.367
R749 B.n479 B.n193 163.367
R750 B.n479 B.n191 163.367
R751 B.n483 B.n191 163.367
R752 B.n483 B.n185 163.367
R753 B.n491 B.n185 163.367
R754 B.n491 B.n183 163.367
R755 B.n495 B.n183 163.367
R756 B.n495 B.n177 163.367
R757 B.n503 B.n177 163.367
R758 B.n503 B.n175 163.367
R759 B.n507 B.n175 163.367
R760 B.n507 B.n169 163.367
R761 B.n515 B.n169 163.367
R762 B.n515 B.n167 163.367
R763 B.n519 B.n167 163.367
R764 B.n519 B.n161 163.367
R765 B.n527 B.n161 163.367
R766 B.n527 B.n159 163.367
R767 B.n531 B.n159 163.367
R768 B.n531 B.n153 163.367
R769 B.n539 B.n153 163.367
R770 B.n539 B.n151 163.367
R771 B.n543 B.n151 163.367
R772 B.n543 B.n145 163.367
R773 B.n552 B.n145 163.367
R774 B.n552 B.n143 163.367
R775 B.n556 B.n143 163.367
R776 B.n556 B.n138 163.367
R777 B.n565 B.n138 163.367
R778 B.n565 B.n136 163.367
R779 B.n569 B.n136 163.367
R780 B.n569 B.n2 163.367
R781 B.n891 B.n2 163.367
R782 B.n891 B.n3 163.367
R783 B.n887 B.n3 163.367
R784 B.n887 B.n9 163.367
R785 B.n883 B.n9 163.367
R786 B.n883 B.n11 163.367
R787 B.n879 B.n11 163.367
R788 B.n879 B.n15 163.367
R789 B.n875 B.n15 163.367
R790 B.n875 B.n17 163.367
R791 B.n871 B.n17 163.367
R792 B.n871 B.n23 163.367
R793 B.n867 B.n23 163.367
R794 B.n867 B.n25 163.367
R795 B.n863 B.n25 163.367
R796 B.n863 B.n30 163.367
R797 B.n859 B.n30 163.367
R798 B.n859 B.n32 163.367
R799 B.n855 B.n32 163.367
R800 B.n855 B.n37 163.367
R801 B.n851 B.n37 163.367
R802 B.n851 B.n39 163.367
R803 B.n847 B.n39 163.367
R804 B.n847 B.n44 163.367
R805 B.n843 B.n44 163.367
R806 B.n843 B.n46 163.367
R807 B.n839 B.n46 163.367
R808 B.n839 B.n51 163.367
R809 B.n835 B.n51 163.367
R810 B.n835 B.n53 163.367
R811 B.n831 B.n53 163.367
R812 B.n831 B.n58 163.367
R813 B.n827 B.n58 163.367
R814 B.n827 B.n60 163.367
R815 B.n823 B.n60 163.367
R816 B.n823 B.n65 163.367
R817 B.n819 B.n65 163.367
R818 B.n819 B.n67 163.367
R819 B.n815 B.n67 163.367
R820 B.n815 B.n71 163.367
R821 B.n811 B.n71 163.367
R822 B.n811 B.n73 163.367
R823 B.n807 B.n73 163.367
R824 B.n807 B.n79 163.367
R825 B.n803 B.n79 163.367
R826 B.n803 B.n81 163.367
R827 B.n799 B.n81 163.367
R828 B.n430 B.n428 163.367
R829 B.n428 B.n427 163.367
R830 B.n424 B.n423 163.367
R831 B.n421 B.n226 163.367
R832 B.n417 B.n415 163.367
R833 B.n413 B.n228 163.367
R834 B.n409 B.n407 163.367
R835 B.n405 B.n230 163.367
R836 B.n401 B.n399 163.367
R837 B.n397 B.n232 163.367
R838 B.n393 B.n391 163.367
R839 B.n389 B.n234 163.367
R840 B.n385 B.n383 163.367
R841 B.n381 B.n236 163.367
R842 B.n377 B.n375 163.367
R843 B.n373 B.n238 163.367
R844 B.n369 B.n367 163.367
R845 B.n365 B.n240 163.367
R846 B.n361 B.n359 163.367
R847 B.n356 B.n355 163.367
R848 B.n353 B.n246 163.367
R849 B.n349 B.n347 163.367
R850 B.n345 B.n248 163.367
R851 B.n340 B.n338 163.367
R852 B.n336 B.n252 163.367
R853 B.n332 B.n330 163.367
R854 B.n328 B.n254 163.367
R855 B.n324 B.n322 163.367
R856 B.n320 B.n256 163.367
R857 B.n316 B.n314 163.367
R858 B.n312 B.n258 163.367
R859 B.n308 B.n306 163.367
R860 B.n304 B.n260 163.367
R861 B.n300 B.n298 163.367
R862 B.n296 B.n262 163.367
R863 B.n292 B.n290 163.367
R864 B.n288 B.n264 163.367
R865 B.n284 B.n282 163.367
R866 B.n280 B.n266 163.367
R867 B.n276 B.n274 163.367
R868 B.n272 B.n269 163.367
R869 B.n436 B.n218 163.367
R870 B.n440 B.n218 163.367
R871 B.n440 B.n212 163.367
R872 B.n448 B.n212 163.367
R873 B.n448 B.n210 163.367
R874 B.n452 B.n210 163.367
R875 B.n452 B.n205 163.367
R876 B.n461 B.n205 163.367
R877 B.n461 B.n203 163.367
R878 B.n465 B.n203 163.367
R879 B.n465 B.n197 163.367
R880 B.n473 B.n197 163.367
R881 B.n473 B.n195 163.367
R882 B.n477 B.n195 163.367
R883 B.n477 B.n189 163.367
R884 B.n485 B.n189 163.367
R885 B.n485 B.n187 163.367
R886 B.n489 B.n187 163.367
R887 B.n489 B.n181 163.367
R888 B.n497 B.n181 163.367
R889 B.n497 B.n179 163.367
R890 B.n501 B.n179 163.367
R891 B.n501 B.n173 163.367
R892 B.n509 B.n173 163.367
R893 B.n509 B.n171 163.367
R894 B.n513 B.n171 163.367
R895 B.n513 B.n165 163.367
R896 B.n521 B.n165 163.367
R897 B.n521 B.n163 163.367
R898 B.n525 B.n163 163.367
R899 B.n525 B.n157 163.367
R900 B.n533 B.n157 163.367
R901 B.n533 B.n155 163.367
R902 B.n537 B.n155 163.367
R903 B.n537 B.n149 163.367
R904 B.n545 B.n149 163.367
R905 B.n545 B.n147 163.367
R906 B.n549 B.n147 163.367
R907 B.n549 B.n142 163.367
R908 B.n558 B.n142 163.367
R909 B.n558 B.n140 163.367
R910 B.n563 B.n140 163.367
R911 B.n563 B.n134 163.367
R912 B.n571 B.n134 163.367
R913 B.n572 B.n571 163.367
R914 B.n572 B.n5 163.367
R915 B.n6 B.n5 163.367
R916 B.n7 B.n6 163.367
R917 B.n577 B.n7 163.367
R918 B.n577 B.n12 163.367
R919 B.n13 B.n12 163.367
R920 B.n14 B.n13 163.367
R921 B.n582 B.n14 163.367
R922 B.n582 B.n19 163.367
R923 B.n20 B.n19 163.367
R924 B.n21 B.n20 163.367
R925 B.n587 B.n21 163.367
R926 B.n587 B.n26 163.367
R927 B.n27 B.n26 163.367
R928 B.n28 B.n27 163.367
R929 B.n592 B.n28 163.367
R930 B.n592 B.n33 163.367
R931 B.n34 B.n33 163.367
R932 B.n35 B.n34 163.367
R933 B.n597 B.n35 163.367
R934 B.n597 B.n40 163.367
R935 B.n41 B.n40 163.367
R936 B.n42 B.n41 163.367
R937 B.n602 B.n42 163.367
R938 B.n602 B.n47 163.367
R939 B.n48 B.n47 163.367
R940 B.n49 B.n48 163.367
R941 B.n607 B.n49 163.367
R942 B.n607 B.n54 163.367
R943 B.n55 B.n54 163.367
R944 B.n56 B.n55 163.367
R945 B.n612 B.n56 163.367
R946 B.n612 B.n61 163.367
R947 B.n62 B.n61 163.367
R948 B.n63 B.n62 163.367
R949 B.n617 B.n63 163.367
R950 B.n617 B.n68 163.367
R951 B.n69 B.n68 163.367
R952 B.n70 B.n69 163.367
R953 B.n622 B.n70 163.367
R954 B.n622 B.n75 163.367
R955 B.n76 B.n75 163.367
R956 B.n77 B.n76 163.367
R957 B.n627 B.n77 163.367
R958 B.n627 B.n82 163.367
R959 B.n83 B.n82 163.367
R960 B.n84 B.n83 163.367
R961 B.n795 B.n793 163.367
R962 B.n791 B.n88 163.367
R963 B.n787 B.n785 163.367
R964 B.n783 B.n90 163.367
R965 B.n779 B.n777 163.367
R966 B.n775 B.n92 163.367
R967 B.n771 B.n769 163.367
R968 B.n767 B.n94 163.367
R969 B.n763 B.n761 163.367
R970 B.n759 B.n96 163.367
R971 B.n755 B.n753 163.367
R972 B.n751 B.n98 163.367
R973 B.n747 B.n745 163.367
R974 B.n743 B.n100 163.367
R975 B.n739 B.n737 163.367
R976 B.n735 B.n102 163.367
R977 B.n731 B.n729 163.367
R978 B.n727 B.n104 163.367
R979 B.n722 B.n720 163.367
R980 B.n718 B.n108 163.367
R981 B.n714 B.n712 163.367
R982 B.n710 B.n110 163.367
R983 B.n706 B.n704 163.367
R984 B.n701 B.n700 163.367
R985 B.n698 B.n116 163.367
R986 B.n694 B.n692 163.367
R987 B.n690 B.n118 163.367
R988 B.n686 B.n684 163.367
R989 B.n682 B.n120 163.367
R990 B.n678 B.n676 163.367
R991 B.n674 B.n122 163.367
R992 B.n670 B.n668 163.367
R993 B.n666 B.n124 163.367
R994 B.n662 B.n660 163.367
R995 B.n658 B.n126 163.367
R996 B.n654 B.n652 163.367
R997 B.n650 B.n128 163.367
R998 B.n646 B.n644 163.367
R999 B.n642 B.n130 163.367
R1000 B.n638 B.n636 163.367
R1001 B.n634 B.n132 163.367
R1002 B.n249 B.t12 132.642
R1003 B.n111 B.t18 132.642
R1004 B.n241 B.t9 132.629
R1005 B.n105 B.t15 132.629
R1006 B.n435 B.n221 92.5206
R1007 B.n800 B.n85 92.5206
R1008 B.n429 B.n222 71.676
R1009 B.n427 B.n224 71.676
R1010 B.n423 B.n422 71.676
R1011 B.n416 B.n226 71.676
R1012 B.n415 B.n414 71.676
R1013 B.n408 B.n228 71.676
R1014 B.n407 B.n406 71.676
R1015 B.n400 B.n230 71.676
R1016 B.n399 B.n398 71.676
R1017 B.n392 B.n232 71.676
R1018 B.n391 B.n390 71.676
R1019 B.n384 B.n234 71.676
R1020 B.n383 B.n382 71.676
R1021 B.n376 B.n236 71.676
R1022 B.n375 B.n374 71.676
R1023 B.n368 B.n238 71.676
R1024 B.n367 B.n366 71.676
R1025 B.n360 B.n240 71.676
R1026 B.n359 B.n244 71.676
R1027 B.n355 B.n354 71.676
R1028 B.n348 B.n246 71.676
R1029 B.n347 B.n346 71.676
R1030 B.n339 B.n248 71.676
R1031 B.n338 B.n337 71.676
R1032 B.n331 B.n252 71.676
R1033 B.n330 B.n329 71.676
R1034 B.n323 B.n254 71.676
R1035 B.n322 B.n321 71.676
R1036 B.n315 B.n256 71.676
R1037 B.n314 B.n313 71.676
R1038 B.n307 B.n258 71.676
R1039 B.n306 B.n305 71.676
R1040 B.n299 B.n260 71.676
R1041 B.n298 B.n297 71.676
R1042 B.n291 B.n262 71.676
R1043 B.n290 B.n289 71.676
R1044 B.n283 B.n264 71.676
R1045 B.n282 B.n281 71.676
R1046 B.n275 B.n266 71.676
R1047 B.n274 B.n273 71.676
R1048 B.n269 B.n268 71.676
R1049 B.n794 B.n86 71.676
R1050 B.n793 B.n792 71.676
R1051 B.n786 B.n88 71.676
R1052 B.n785 B.n784 71.676
R1053 B.n778 B.n90 71.676
R1054 B.n777 B.n776 71.676
R1055 B.n770 B.n92 71.676
R1056 B.n769 B.n768 71.676
R1057 B.n762 B.n94 71.676
R1058 B.n761 B.n760 71.676
R1059 B.n754 B.n96 71.676
R1060 B.n753 B.n752 71.676
R1061 B.n746 B.n98 71.676
R1062 B.n745 B.n744 71.676
R1063 B.n738 B.n100 71.676
R1064 B.n737 B.n736 71.676
R1065 B.n730 B.n102 71.676
R1066 B.n729 B.n728 71.676
R1067 B.n721 B.n104 71.676
R1068 B.n720 B.n719 71.676
R1069 B.n713 B.n108 71.676
R1070 B.n712 B.n711 71.676
R1071 B.n705 B.n110 71.676
R1072 B.n704 B.n114 71.676
R1073 B.n700 B.n699 71.676
R1074 B.n693 B.n116 71.676
R1075 B.n692 B.n691 71.676
R1076 B.n685 B.n118 71.676
R1077 B.n684 B.n683 71.676
R1078 B.n677 B.n120 71.676
R1079 B.n676 B.n675 71.676
R1080 B.n669 B.n122 71.676
R1081 B.n668 B.n667 71.676
R1082 B.n661 B.n124 71.676
R1083 B.n660 B.n659 71.676
R1084 B.n653 B.n126 71.676
R1085 B.n652 B.n651 71.676
R1086 B.n645 B.n128 71.676
R1087 B.n644 B.n643 71.676
R1088 B.n637 B.n130 71.676
R1089 B.n636 B.n635 71.676
R1090 B.n635 B.n634 71.676
R1091 B.n638 B.n637 71.676
R1092 B.n643 B.n642 71.676
R1093 B.n646 B.n645 71.676
R1094 B.n651 B.n650 71.676
R1095 B.n654 B.n653 71.676
R1096 B.n659 B.n658 71.676
R1097 B.n662 B.n661 71.676
R1098 B.n667 B.n666 71.676
R1099 B.n670 B.n669 71.676
R1100 B.n675 B.n674 71.676
R1101 B.n678 B.n677 71.676
R1102 B.n683 B.n682 71.676
R1103 B.n686 B.n685 71.676
R1104 B.n691 B.n690 71.676
R1105 B.n694 B.n693 71.676
R1106 B.n699 B.n698 71.676
R1107 B.n701 B.n114 71.676
R1108 B.n706 B.n705 71.676
R1109 B.n711 B.n710 71.676
R1110 B.n714 B.n713 71.676
R1111 B.n719 B.n718 71.676
R1112 B.n722 B.n721 71.676
R1113 B.n728 B.n727 71.676
R1114 B.n731 B.n730 71.676
R1115 B.n736 B.n735 71.676
R1116 B.n739 B.n738 71.676
R1117 B.n744 B.n743 71.676
R1118 B.n747 B.n746 71.676
R1119 B.n752 B.n751 71.676
R1120 B.n755 B.n754 71.676
R1121 B.n760 B.n759 71.676
R1122 B.n763 B.n762 71.676
R1123 B.n768 B.n767 71.676
R1124 B.n771 B.n770 71.676
R1125 B.n776 B.n775 71.676
R1126 B.n779 B.n778 71.676
R1127 B.n784 B.n783 71.676
R1128 B.n787 B.n786 71.676
R1129 B.n792 B.n791 71.676
R1130 B.n795 B.n794 71.676
R1131 B.n430 B.n429 71.676
R1132 B.n424 B.n224 71.676
R1133 B.n422 B.n421 71.676
R1134 B.n417 B.n416 71.676
R1135 B.n414 B.n413 71.676
R1136 B.n409 B.n408 71.676
R1137 B.n406 B.n405 71.676
R1138 B.n401 B.n400 71.676
R1139 B.n398 B.n397 71.676
R1140 B.n393 B.n392 71.676
R1141 B.n390 B.n389 71.676
R1142 B.n385 B.n384 71.676
R1143 B.n382 B.n381 71.676
R1144 B.n377 B.n376 71.676
R1145 B.n374 B.n373 71.676
R1146 B.n369 B.n368 71.676
R1147 B.n366 B.n365 71.676
R1148 B.n361 B.n360 71.676
R1149 B.n356 B.n244 71.676
R1150 B.n354 B.n353 71.676
R1151 B.n349 B.n348 71.676
R1152 B.n346 B.n345 71.676
R1153 B.n340 B.n339 71.676
R1154 B.n337 B.n336 71.676
R1155 B.n332 B.n331 71.676
R1156 B.n329 B.n328 71.676
R1157 B.n324 B.n323 71.676
R1158 B.n321 B.n320 71.676
R1159 B.n316 B.n315 71.676
R1160 B.n313 B.n312 71.676
R1161 B.n308 B.n307 71.676
R1162 B.n305 B.n304 71.676
R1163 B.n300 B.n299 71.676
R1164 B.n297 B.n296 71.676
R1165 B.n292 B.n291 71.676
R1166 B.n289 B.n288 71.676
R1167 B.n284 B.n283 71.676
R1168 B.n281 B.n280 71.676
R1169 B.n276 B.n275 71.676
R1170 B.n273 B.n272 71.676
R1171 B.n268 B.n220 71.676
R1172 B.n250 B.t11 69.9991
R1173 B.n112 B.t19 69.9991
R1174 B.n242 B.t8 69.9864
R1175 B.n106 B.t16 69.9864
R1176 B.n250 B.n249 62.6429
R1177 B.n242 B.n241 62.6429
R1178 B.n106 B.n105 62.6429
R1179 B.n112 B.n111 62.6429
R1180 B.n342 B.n250 59.5399
R1181 B.n243 B.n242 59.5399
R1182 B.n724 B.n106 59.5399
R1183 B.n113 B.n112 59.5399
R1184 B.n435 B.n217 48.0262
R1185 B.n441 B.n217 48.0262
R1186 B.n441 B.n213 48.0262
R1187 B.n447 B.n213 48.0262
R1188 B.n447 B.n209 48.0262
R1189 B.n454 B.n209 48.0262
R1190 B.n454 B.n453 48.0262
R1191 B.n460 B.n202 48.0262
R1192 B.n466 B.n202 48.0262
R1193 B.n466 B.n198 48.0262
R1194 B.n472 B.n198 48.0262
R1195 B.n472 B.n194 48.0262
R1196 B.n478 B.n194 48.0262
R1197 B.n478 B.n190 48.0262
R1198 B.n484 B.n190 48.0262
R1199 B.n484 B.n186 48.0262
R1200 B.n490 B.n186 48.0262
R1201 B.n490 B.n182 48.0262
R1202 B.n496 B.n182 48.0262
R1203 B.n502 B.n178 48.0262
R1204 B.n502 B.n174 48.0262
R1205 B.n508 B.n174 48.0262
R1206 B.n508 B.n170 48.0262
R1207 B.n514 B.n170 48.0262
R1208 B.n514 B.n166 48.0262
R1209 B.n520 B.n166 48.0262
R1210 B.n520 B.n162 48.0262
R1211 B.n526 B.n162 48.0262
R1212 B.n532 B.n158 48.0262
R1213 B.n532 B.n154 48.0262
R1214 B.n538 B.n154 48.0262
R1215 B.n538 B.n150 48.0262
R1216 B.n544 B.n150 48.0262
R1217 B.n544 B.n146 48.0262
R1218 B.n551 B.n146 48.0262
R1219 B.n551 B.n550 48.0262
R1220 B.n557 B.n139 48.0262
R1221 B.n564 B.n139 48.0262
R1222 B.n564 B.n135 48.0262
R1223 B.n570 B.n135 48.0262
R1224 B.n570 B.n4 48.0262
R1225 B.n890 B.n4 48.0262
R1226 B.n890 B.n889 48.0262
R1227 B.n889 B.n888 48.0262
R1228 B.n888 B.n8 48.0262
R1229 B.n882 B.n8 48.0262
R1230 B.n882 B.n881 48.0262
R1231 B.n881 B.n880 48.0262
R1232 B.n874 B.n18 48.0262
R1233 B.n874 B.n873 48.0262
R1234 B.n873 B.n872 48.0262
R1235 B.n872 B.n22 48.0262
R1236 B.n866 B.n22 48.0262
R1237 B.n866 B.n865 48.0262
R1238 B.n865 B.n864 48.0262
R1239 B.n864 B.n29 48.0262
R1240 B.n858 B.n857 48.0262
R1241 B.n857 B.n856 48.0262
R1242 B.n856 B.n36 48.0262
R1243 B.n850 B.n36 48.0262
R1244 B.n850 B.n849 48.0262
R1245 B.n849 B.n848 48.0262
R1246 B.n848 B.n43 48.0262
R1247 B.n842 B.n43 48.0262
R1248 B.n842 B.n841 48.0262
R1249 B.n840 B.n50 48.0262
R1250 B.n834 B.n50 48.0262
R1251 B.n834 B.n833 48.0262
R1252 B.n833 B.n832 48.0262
R1253 B.n832 B.n57 48.0262
R1254 B.n826 B.n57 48.0262
R1255 B.n826 B.n825 48.0262
R1256 B.n825 B.n824 48.0262
R1257 B.n824 B.n64 48.0262
R1258 B.n818 B.n64 48.0262
R1259 B.n818 B.n817 48.0262
R1260 B.n817 B.n816 48.0262
R1261 B.n810 B.n74 48.0262
R1262 B.n810 B.n809 48.0262
R1263 B.n809 B.n808 48.0262
R1264 B.n808 B.n78 48.0262
R1265 B.n802 B.n78 48.0262
R1266 B.n802 B.n801 48.0262
R1267 B.n801 B.n800 48.0262
R1268 B.n453 B.t7 45.2011
R1269 B.n74 B.t14 45.2011
R1270 B.t5 B.n158 40.9636
R1271 B.t1 B.n29 40.9636
R1272 B.n798 B.n797 32.6249
R1273 B.n632 B.n631 32.6249
R1274 B.n437 B.n219 32.6249
R1275 B.n433 B.n432 32.6249
R1276 B.n496 B.t2 31.0759
R1277 B.n550 B.t0 31.0759
R1278 B.n18 B.t4 31.0759
R1279 B.t3 B.n840 31.0759
R1280 B B.n892 18.0485
R1281 B.t2 B.n178 16.9507
R1282 B.n557 B.t0 16.9507
R1283 B.n880 B.t4 16.9507
R1284 B.n841 B.t3 16.9507
R1285 B.n797 B.n796 10.6151
R1286 B.n796 B.n87 10.6151
R1287 B.n790 B.n87 10.6151
R1288 B.n790 B.n789 10.6151
R1289 B.n789 B.n788 10.6151
R1290 B.n788 B.n89 10.6151
R1291 B.n782 B.n89 10.6151
R1292 B.n782 B.n781 10.6151
R1293 B.n781 B.n780 10.6151
R1294 B.n780 B.n91 10.6151
R1295 B.n774 B.n91 10.6151
R1296 B.n774 B.n773 10.6151
R1297 B.n773 B.n772 10.6151
R1298 B.n772 B.n93 10.6151
R1299 B.n766 B.n93 10.6151
R1300 B.n766 B.n765 10.6151
R1301 B.n765 B.n764 10.6151
R1302 B.n764 B.n95 10.6151
R1303 B.n758 B.n95 10.6151
R1304 B.n758 B.n757 10.6151
R1305 B.n757 B.n756 10.6151
R1306 B.n756 B.n97 10.6151
R1307 B.n750 B.n97 10.6151
R1308 B.n750 B.n749 10.6151
R1309 B.n749 B.n748 10.6151
R1310 B.n748 B.n99 10.6151
R1311 B.n742 B.n99 10.6151
R1312 B.n742 B.n741 10.6151
R1313 B.n741 B.n740 10.6151
R1314 B.n740 B.n101 10.6151
R1315 B.n734 B.n101 10.6151
R1316 B.n734 B.n733 10.6151
R1317 B.n733 B.n732 10.6151
R1318 B.n732 B.n103 10.6151
R1319 B.n726 B.n103 10.6151
R1320 B.n726 B.n725 10.6151
R1321 B.n723 B.n107 10.6151
R1322 B.n717 B.n107 10.6151
R1323 B.n717 B.n716 10.6151
R1324 B.n716 B.n715 10.6151
R1325 B.n715 B.n109 10.6151
R1326 B.n709 B.n109 10.6151
R1327 B.n709 B.n708 10.6151
R1328 B.n708 B.n707 10.6151
R1329 B.n703 B.n702 10.6151
R1330 B.n702 B.n115 10.6151
R1331 B.n697 B.n115 10.6151
R1332 B.n697 B.n696 10.6151
R1333 B.n696 B.n695 10.6151
R1334 B.n695 B.n117 10.6151
R1335 B.n689 B.n117 10.6151
R1336 B.n689 B.n688 10.6151
R1337 B.n688 B.n687 10.6151
R1338 B.n687 B.n119 10.6151
R1339 B.n681 B.n119 10.6151
R1340 B.n681 B.n680 10.6151
R1341 B.n680 B.n679 10.6151
R1342 B.n679 B.n121 10.6151
R1343 B.n673 B.n121 10.6151
R1344 B.n673 B.n672 10.6151
R1345 B.n672 B.n671 10.6151
R1346 B.n671 B.n123 10.6151
R1347 B.n665 B.n123 10.6151
R1348 B.n665 B.n664 10.6151
R1349 B.n664 B.n663 10.6151
R1350 B.n663 B.n125 10.6151
R1351 B.n657 B.n125 10.6151
R1352 B.n657 B.n656 10.6151
R1353 B.n656 B.n655 10.6151
R1354 B.n655 B.n127 10.6151
R1355 B.n649 B.n127 10.6151
R1356 B.n649 B.n648 10.6151
R1357 B.n648 B.n647 10.6151
R1358 B.n647 B.n129 10.6151
R1359 B.n641 B.n129 10.6151
R1360 B.n641 B.n640 10.6151
R1361 B.n640 B.n639 10.6151
R1362 B.n639 B.n131 10.6151
R1363 B.n633 B.n131 10.6151
R1364 B.n633 B.n632 10.6151
R1365 B.n438 B.n437 10.6151
R1366 B.n439 B.n438 10.6151
R1367 B.n439 B.n211 10.6151
R1368 B.n449 B.n211 10.6151
R1369 B.n450 B.n449 10.6151
R1370 B.n451 B.n450 10.6151
R1371 B.n451 B.n204 10.6151
R1372 B.n462 B.n204 10.6151
R1373 B.n463 B.n462 10.6151
R1374 B.n464 B.n463 10.6151
R1375 B.n464 B.n196 10.6151
R1376 B.n474 B.n196 10.6151
R1377 B.n475 B.n474 10.6151
R1378 B.n476 B.n475 10.6151
R1379 B.n476 B.n188 10.6151
R1380 B.n486 B.n188 10.6151
R1381 B.n487 B.n486 10.6151
R1382 B.n488 B.n487 10.6151
R1383 B.n488 B.n180 10.6151
R1384 B.n498 B.n180 10.6151
R1385 B.n499 B.n498 10.6151
R1386 B.n500 B.n499 10.6151
R1387 B.n500 B.n172 10.6151
R1388 B.n510 B.n172 10.6151
R1389 B.n511 B.n510 10.6151
R1390 B.n512 B.n511 10.6151
R1391 B.n512 B.n164 10.6151
R1392 B.n522 B.n164 10.6151
R1393 B.n523 B.n522 10.6151
R1394 B.n524 B.n523 10.6151
R1395 B.n524 B.n156 10.6151
R1396 B.n534 B.n156 10.6151
R1397 B.n535 B.n534 10.6151
R1398 B.n536 B.n535 10.6151
R1399 B.n536 B.n148 10.6151
R1400 B.n546 B.n148 10.6151
R1401 B.n547 B.n546 10.6151
R1402 B.n548 B.n547 10.6151
R1403 B.n548 B.n141 10.6151
R1404 B.n559 B.n141 10.6151
R1405 B.n560 B.n559 10.6151
R1406 B.n562 B.n560 10.6151
R1407 B.n562 B.n561 10.6151
R1408 B.n561 B.n133 10.6151
R1409 B.n573 B.n133 10.6151
R1410 B.n574 B.n573 10.6151
R1411 B.n575 B.n574 10.6151
R1412 B.n576 B.n575 10.6151
R1413 B.n578 B.n576 10.6151
R1414 B.n579 B.n578 10.6151
R1415 B.n580 B.n579 10.6151
R1416 B.n581 B.n580 10.6151
R1417 B.n583 B.n581 10.6151
R1418 B.n584 B.n583 10.6151
R1419 B.n585 B.n584 10.6151
R1420 B.n586 B.n585 10.6151
R1421 B.n588 B.n586 10.6151
R1422 B.n589 B.n588 10.6151
R1423 B.n590 B.n589 10.6151
R1424 B.n591 B.n590 10.6151
R1425 B.n593 B.n591 10.6151
R1426 B.n594 B.n593 10.6151
R1427 B.n595 B.n594 10.6151
R1428 B.n596 B.n595 10.6151
R1429 B.n598 B.n596 10.6151
R1430 B.n599 B.n598 10.6151
R1431 B.n600 B.n599 10.6151
R1432 B.n601 B.n600 10.6151
R1433 B.n603 B.n601 10.6151
R1434 B.n604 B.n603 10.6151
R1435 B.n605 B.n604 10.6151
R1436 B.n606 B.n605 10.6151
R1437 B.n608 B.n606 10.6151
R1438 B.n609 B.n608 10.6151
R1439 B.n610 B.n609 10.6151
R1440 B.n611 B.n610 10.6151
R1441 B.n613 B.n611 10.6151
R1442 B.n614 B.n613 10.6151
R1443 B.n615 B.n614 10.6151
R1444 B.n616 B.n615 10.6151
R1445 B.n618 B.n616 10.6151
R1446 B.n619 B.n618 10.6151
R1447 B.n620 B.n619 10.6151
R1448 B.n621 B.n620 10.6151
R1449 B.n623 B.n621 10.6151
R1450 B.n624 B.n623 10.6151
R1451 B.n625 B.n624 10.6151
R1452 B.n626 B.n625 10.6151
R1453 B.n628 B.n626 10.6151
R1454 B.n629 B.n628 10.6151
R1455 B.n630 B.n629 10.6151
R1456 B.n631 B.n630 10.6151
R1457 B.n432 B.n431 10.6151
R1458 B.n431 B.n223 10.6151
R1459 B.n426 B.n223 10.6151
R1460 B.n426 B.n425 10.6151
R1461 B.n425 B.n225 10.6151
R1462 B.n420 B.n225 10.6151
R1463 B.n420 B.n419 10.6151
R1464 B.n419 B.n418 10.6151
R1465 B.n418 B.n227 10.6151
R1466 B.n412 B.n227 10.6151
R1467 B.n412 B.n411 10.6151
R1468 B.n411 B.n410 10.6151
R1469 B.n410 B.n229 10.6151
R1470 B.n404 B.n229 10.6151
R1471 B.n404 B.n403 10.6151
R1472 B.n403 B.n402 10.6151
R1473 B.n402 B.n231 10.6151
R1474 B.n396 B.n231 10.6151
R1475 B.n396 B.n395 10.6151
R1476 B.n395 B.n394 10.6151
R1477 B.n394 B.n233 10.6151
R1478 B.n388 B.n233 10.6151
R1479 B.n388 B.n387 10.6151
R1480 B.n387 B.n386 10.6151
R1481 B.n386 B.n235 10.6151
R1482 B.n380 B.n235 10.6151
R1483 B.n380 B.n379 10.6151
R1484 B.n379 B.n378 10.6151
R1485 B.n378 B.n237 10.6151
R1486 B.n372 B.n237 10.6151
R1487 B.n372 B.n371 10.6151
R1488 B.n371 B.n370 10.6151
R1489 B.n370 B.n239 10.6151
R1490 B.n364 B.n239 10.6151
R1491 B.n364 B.n363 10.6151
R1492 B.n363 B.n362 10.6151
R1493 B.n358 B.n357 10.6151
R1494 B.n357 B.n245 10.6151
R1495 B.n352 B.n245 10.6151
R1496 B.n352 B.n351 10.6151
R1497 B.n351 B.n350 10.6151
R1498 B.n350 B.n247 10.6151
R1499 B.n344 B.n247 10.6151
R1500 B.n344 B.n343 10.6151
R1501 B.n341 B.n251 10.6151
R1502 B.n335 B.n251 10.6151
R1503 B.n335 B.n334 10.6151
R1504 B.n334 B.n333 10.6151
R1505 B.n333 B.n253 10.6151
R1506 B.n327 B.n253 10.6151
R1507 B.n327 B.n326 10.6151
R1508 B.n326 B.n325 10.6151
R1509 B.n325 B.n255 10.6151
R1510 B.n319 B.n255 10.6151
R1511 B.n319 B.n318 10.6151
R1512 B.n318 B.n317 10.6151
R1513 B.n317 B.n257 10.6151
R1514 B.n311 B.n257 10.6151
R1515 B.n311 B.n310 10.6151
R1516 B.n310 B.n309 10.6151
R1517 B.n309 B.n259 10.6151
R1518 B.n303 B.n259 10.6151
R1519 B.n303 B.n302 10.6151
R1520 B.n302 B.n301 10.6151
R1521 B.n301 B.n261 10.6151
R1522 B.n295 B.n261 10.6151
R1523 B.n295 B.n294 10.6151
R1524 B.n294 B.n293 10.6151
R1525 B.n293 B.n263 10.6151
R1526 B.n287 B.n263 10.6151
R1527 B.n287 B.n286 10.6151
R1528 B.n286 B.n285 10.6151
R1529 B.n285 B.n265 10.6151
R1530 B.n279 B.n265 10.6151
R1531 B.n279 B.n278 10.6151
R1532 B.n278 B.n277 10.6151
R1533 B.n277 B.n267 10.6151
R1534 B.n271 B.n267 10.6151
R1535 B.n271 B.n270 10.6151
R1536 B.n270 B.n219 10.6151
R1537 B.n433 B.n215 10.6151
R1538 B.n443 B.n215 10.6151
R1539 B.n444 B.n443 10.6151
R1540 B.n445 B.n444 10.6151
R1541 B.n445 B.n207 10.6151
R1542 B.n456 B.n207 10.6151
R1543 B.n457 B.n456 10.6151
R1544 B.n458 B.n457 10.6151
R1545 B.n458 B.n200 10.6151
R1546 B.n468 B.n200 10.6151
R1547 B.n469 B.n468 10.6151
R1548 B.n470 B.n469 10.6151
R1549 B.n470 B.n192 10.6151
R1550 B.n480 B.n192 10.6151
R1551 B.n481 B.n480 10.6151
R1552 B.n482 B.n481 10.6151
R1553 B.n482 B.n184 10.6151
R1554 B.n492 B.n184 10.6151
R1555 B.n493 B.n492 10.6151
R1556 B.n494 B.n493 10.6151
R1557 B.n494 B.n176 10.6151
R1558 B.n504 B.n176 10.6151
R1559 B.n505 B.n504 10.6151
R1560 B.n506 B.n505 10.6151
R1561 B.n506 B.n168 10.6151
R1562 B.n516 B.n168 10.6151
R1563 B.n517 B.n516 10.6151
R1564 B.n518 B.n517 10.6151
R1565 B.n518 B.n160 10.6151
R1566 B.n528 B.n160 10.6151
R1567 B.n529 B.n528 10.6151
R1568 B.n530 B.n529 10.6151
R1569 B.n530 B.n152 10.6151
R1570 B.n540 B.n152 10.6151
R1571 B.n541 B.n540 10.6151
R1572 B.n542 B.n541 10.6151
R1573 B.n542 B.n144 10.6151
R1574 B.n553 B.n144 10.6151
R1575 B.n554 B.n553 10.6151
R1576 B.n555 B.n554 10.6151
R1577 B.n555 B.n137 10.6151
R1578 B.n566 B.n137 10.6151
R1579 B.n567 B.n566 10.6151
R1580 B.n568 B.n567 10.6151
R1581 B.n568 B.n0 10.6151
R1582 B.n886 B.n1 10.6151
R1583 B.n886 B.n885 10.6151
R1584 B.n885 B.n884 10.6151
R1585 B.n884 B.n10 10.6151
R1586 B.n878 B.n10 10.6151
R1587 B.n878 B.n877 10.6151
R1588 B.n877 B.n876 10.6151
R1589 B.n876 B.n16 10.6151
R1590 B.n870 B.n16 10.6151
R1591 B.n870 B.n869 10.6151
R1592 B.n869 B.n868 10.6151
R1593 B.n868 B.n24 10.6151
R1594 B.n862 B.n24 10.6151
R1595 B.n862 B.n861 10.6151
R1596 B.n861 B.n860 10.6151
R1597 B.n860 B.n31 10.6151
R1598 B.n854 B.n31 10.6151
R1599 B.n854 B.n853 10.6151
R1600 B.n853 B.n852 10.6151
R1601 B.n852 B.n38 10.6151
R1602 B.n846 B.n38 10.6151
R1603 B.n846 B.n845 10.6151
R1604 B.n845 B.n844 10.6151
R1605 B.n844 B.n45 10.6151
R1606 B.n838 B.n45 10.6151
R1607 B.n838 B.n837 10.6151
R1608 B.n837 B.n836 10.6151
R1609 B.n836 B.n52 10.6151
R1610 B.n830 B.n52 10.6151
R1611 B.n830 B.n829 10.6151
R1612 B.n829 B.n828 10.6151
R1613 B.n828 B.n59 10.6151
R1614 B.n822 B.n59 10.6151
R1615 B.n822 B.n821 10.6151
R1616 B.n821 B.n820 10.6151
R1617 B.n820 B.n66 10.6151
R1618 B.n814 B.n66 10.6151
R1619 B.n814 B.n813 10.6151
R1620 B.n813 B.n812 10.6151
R1621 B.n812 B.n72 10.6151
R1622 B.n806 B.n72 10.6151
R1623 B.n806 B.n805 10.6151
R1624 B.n805 B.n804 10.6151
R1625 B.n804 B.n80 10.6151
R1626 B.n798 B.n80 10.6151
R1627 B.n526 B.t5 7.0631
R1628 B.n858 B.t1 7.0631
R1629 B.n724 B.n723 6.5566
R1630 B.n707 B.n113 6.5566
R1631 B.n358 B.n243 6.5566
R1632 B.n343 B.n342 6.5566
R1633 B.n725 B.n724 4.05904
R1634 B.n703 B.n113 4.05904
R1635 B.n362 B.n243 4.05904
R1636 B.n342 B.n341 4.05904
R1637 B.n460 B.t7 2.82554
R1638 B.n816 B.t14 2.82554
R1639 B.n892 B.n0 2.81026
R1640 B.n892 B.n1 2.81026
R1641 VN.n30 VN.n29 161.3
R1642 VN.n28 VN.n17 161.3
R1643 VN.n27 VN.n26 161.3
R1644 VN.n25 VN.n18 161.3
R1645 VN.n24 VN.n23 161.3
R1646 VN.n22 VN.n19 161.3
R1647 VN.n14 VN.n13 161.3
R1648 VN.n12 VN.n1 161.3
R1649 VN.n11 VN.n10 161.3
R1650 VN.n9 VN.n2 161.3
R1651 VN.n8 VN.n7 161.3
R1652 VN.n6 VN.n3 161.3
R1653 VN.n20 VN.t3 117.368
R1654 VN.n4 VN.t0 117.368
R1655 VN.n5 VN.t5 85.5971
R1656 VN.n0 VN.t2 85.5971
R1657 VN.n21 VN.t4 85.5971
R1658 VN.n16 VN.t1 85.5971
R1659 VN.n15 VN.n0 66.5213
R1660 VN.n31 VN.n16 66.5213
R1661 VN.n5 VN.n4 61.4167
R1662 VN.n21 VN.n20 61.4167
R1663 VN.n11 VN.n2 53.5561
R1664 VN.n27 VN.n18 53.5561
R1665 VN VN.n31 48.8805
R1666 VN.n12 VN.n11 27.2651
R1667 VN.n28 VN.n27 27.2651
R1668 VN.n7 VN.n6 24.3439
R1669 VN.n7 VN.n2 24.3439
R1670 VN.n13 VN.n12 24.3439
R1671 VN.n23 VN.n18 24.3439
R1672 VN.n23 VN.n22 24.3439
R1673 VN.n29 VN.n28 24.3439
R1674 VN.n13 VN.n0 23.3702
R1675 VN.n29 VN.n16 23.3702
R1676 VN.n6 VN.n5 12.1722
R1677 VN.n22 VN.n21 12.1722
R1678 VN.n20 VN.n19 5.30782
R1679 VN.n4 VN.n3 5.30782
R1680 VN.n31 VN.n30 0.355081
R1681 VN.n15 VN.n14 0.355081
R1682 VN VN.n15 0.26685
R1683 VN.n30 VN.n17 0.189894
R1684 VN.n26 VN.n17 0.189894
R1685 VN.n26 VN.n25 0.189894
R1686 VN.n25 VN.n24 0.189894
R1687 VN.n24 VN.n19 0.189894
R1688 VN.n8 VN.n3 0.189894
R1689 VN.n9 VN.n8 0.189894
R1690 VN.n10 VN.n9 0.189894
R1691 VN.n10 VN.n1 0.189894
R1692 VN.n14 VN.n1 0.189894
R1693 VDD2.n1 VDD2.t5 66.0502
R1694 VDD2.n2 VDD2.t4 64.0174
R1695 VDD2.n1 VDD2.n0 62.7357
R1696 VDD2 VDD2.n3 62.7329
R1697 VDD2.n2 VDD2.n1 41.6442
R1698 VDD2 VDD2.n2 2.14705
R1699 VDD2.n3 VDD2.t1 1.92283
R1700 VDD2.n3 VDD2.t2 1.92283
R1701 VDD2.n0 VDD2.t0 1.92283
R1702 VDD2.n0 VDD2.t3 1.92283
C0 VTAIL VDD1 7.20618f
C1 VDD1 VP 6.26977f
C2 VN VDD1 0.15084f
C3 VDD2 VTAIL 7.259681f
C4 VDD2 VP 0.483318f
C5 VTAIL VP 6.26389f
C6 VDD2 VN 5.94015f
C7 VN VTAIL 6.24965f
C8 VN VP 6.91024f
C9 VDD2 VDD1 1.52394f
C10 VDD2 B 5.914577f
C11 VDD1 B 6.254151f
C12 VTAIL B 7.335035f
C13 VN B 13.63908f
C14 VP B 12.324059f
C15 VDD2.t5 B 1.97333f
C16 VDD2.t0 B 0.174649f
C17 VDD2.t3 B 0.174649f
C18 VDD2.n0 B 1.54493f
C19 VDD2.n1 B 2.51308f
C20 VDD2.t4 B 1.96162f
C21 VDD2.n2 B 2.35425f
C22 VDD2.t1 B 0.174649f
C23 VDD2.t2 B 0.174649f
C24 VDD2.n3 B 1.5449f
C25 VN.t2 B 1.78959f
C26 VN.n0 B 0.727621f
C27 VN.n1 B 0.022093f
C28 VN.n2 B 0.039154f
C29 VN.n3 B 0.234964f
C30 VN.t5 B 1.78959f
C31 VN.t0 B 2.00242f
C32 VN.n4 B 0.684007f
C33 VN.n5 B 0.706397f
C34 VN.n6 B 0.031167f
C35 VN.n7 B 0.041383f
C36 VN.n8 B 0.022093f
C37 VN.n9 B 0.022093f
C38 VN.n10 B 0.022093f
C39 VN.n11 B 0.023705f
C40 VN.n12 B 0.04331f
C41 VN.n13 B 0.040566f
C42 VN.n14 B 0.035664f
C43 VN.n15 B 0.041639f
C44 VN.t1 B 1.78959f
C45 VN.n16 B 0.727621f
C46 VN.n17 B 0.022093f
C47 VN.n18 B 0.039154f
C48 VN.n19 B 0.234964f
C49 VN.t4 B 1.78959f
C50 VN.t3 B 2.00242f
C51 VN.n20 B 0.684007f
C52 VN.n21 B 0.706397f
C53 VN.n22 B 0.031167f
C54 VN.n23 B 0.041383f
C55 VN.n24 B 0.022093f
C56 VN.n25 B 0.022093f
C57 VN.n26 B 0.022093f
C58 VN.n27 B 0.023705f
C59 VN.n28 B 0.04331f
C60 VN.n29 B 0.040566f
C61 VN.n30 B 0.035664f
C62 VN.n31 B 1.20756f
C63 VDD1.t4 B 2.00703f
C64 VDD1.t3 B 2.00613f
C65 VDD1.t0 B 0.177552f
C66 VDD1.t5 B 0.177552f
C67 VDD1.n0 B 1.57061f
C68 VDD1.n1 B 2.66875f
C69 VDD1.t2 B 0.177552f
C70 VDD1.t1 B 0.177552f
C71 VDD1.n2 B 1.56623f
C72 VDD1.n3 B 2.39352f
C73 VTAIL.t4 B 0.199538f
C74 VTAIL.t1 B 0.199538f
C75 VTAIL.n0 B 1.68813f
C76 VTAIL.n1 B 0.446238f
C77 VTAIL.t10 B 2.14977f
C78 VTAIL.n2 B 0.689156f
C79 VTAIL.t11 B 0.199538f
C80 VTAIL.t7 B 0.199538f
C81 VTAIL.n3 B 1.68813f
C82 VTAIL.n4 B 1.93384f
C83 VTAIL.t2 B 0.199538f
C84 VTAIL.t5 B 0.199538f
C85 VTAIL.n5 B 1.68814f
C86 VTAIL.n6 B 1.93384f
C87 VTAIL.t0 B 2.14978f
C88 VTAIL.n7 B 0.689151f
C89 VTAIL.t6 B 0.199538f
C90 VTAIL.t9 B 0.199538f
C91 VTAIL.n8 B 1.68814f
C92 VTAIL.n9 B 0.606602f
C93 VTAIL.t8 B 2.14977f
C94 VTAIL.n10 B 1.79644f
C95 VTAIL.t3 B 2.14977f
C96 VTAIL.n11 B 1.73685f
C97 VP.t0 B 1.83969f
C98 VP.n0 B 0.747991f
C99 VP.n1 B 0.022712f
C100 VP.n2 B 0.04025f
C101 VP.n3 B 0.022712f
C102 VP.t5 B 1.83969f
C103 VP.n4 B 0.042542f
C104 VP.n5 B 0.022712f
C105 VP.n6 B 0.041702f
C106 VP.t4 B 1.83969f
C107 VP.n7 B 0.747991f
C108 VP.n8 B 0.022712f
C109 VP.n9 B 0.04025f
C110 VP.n10 B 0.241542f
C111 VP.t3 B 1.83969f
C112 VP.t1 B 2.05848f
C113 VP.n11 B 0.703158f
C114 VP.n12 B 0.726173f
C115 VP.n13 B 0.03204f
C116 VP.n14 B 0.042542f
C117 VP.n15 B 0.022712f
C118 VP.n16 B 0.022712f
C119 VP.n17 B 0.022712f
C120 VP.n18 B 0.024369f
C121 VP.n19 B 0.044522f
C122 VP.n20 B 0.041702f
C123 VP.n21 B 0.036662f
C124 VP.n22 B 1.23199f
C125 VP.t2 B 1.83969f
C126 VP.n23 B 0.747991f
C127 VP.n24 B 1.2487f
C128 VP.n25 B 0.036662f
C129 VP.n26 B 0.022712f
C130 VP.n27 B 0.044522f
C131 VP.n28 B 0.024369f
C132 VP.n29 B 0.04025f
C133 VP.n30 B 0.022712f
C134 VP.n31 B 0.022712f
C135 VP.n32 B 0.022712f
C136 VP.n33 B 0.03204f
C137 VP.n34 B 0.654744f
C138 VP.n35 B 0.03204f
C139 VP.n36 B 0.042542f
C140 VP.n37 B 0.022712f
C141 VP.n38 B 0.022712f
C142 VP.n39 B 0.022712f
C143 VP.n40 B 0.024369f
C144 VP.n41 B 0.044522f
C145 VP.n42 B 0.041702f
C146 VP.n43 B 0.036662f
C147 VP.n44 B 0.042805f
.ends

