* NGSPICE file created from diff_pair_sample_0767.ext - technology: sky130A

.subckt diff_pair_sample_0767 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t2 w_n2146_n4910# sky130_fd_pr__pfet_01v8 ad=3.25215 pd=20.04 as=3.25215 ps=20.04 w=19.71 l=1.14
X1 VTAIL.t2 VP.t0 VDD1.t5 w_n2146_n4910# sky130_fd_pr__pfet_01v8 ad=3.25215 pd=20.04 as=3.25215 ps=20.04 w=19.71 l=1.14
X2 B.t11 B.t9 B.t10 w_n2146_n4910# sky130_fd_pr__pfet_01v8 ad=7.6869 pd=40.2 as=0 ps=0 w=19.71 l=1.14
X3 B.t8 B.t6 B.t7 w_n2146_n4910# sky130_fd_pr__pfet_01v8 ad=7.6869 pd=40.2 as=0 ps=0 w=19.71 l=1.14
X4 B.t5 B.t3 B.t4 w_n2146_n4910# sky130_fd_pr__pfet_01v8 ad=7.6869 pd=40.2 as=0 ps=0 w=19.71 l=1.14
X5 VDD1.t4 VP.t1 VTAIL.t3 w_n2146_n4910# sky130_fd_pr__pfet_01v8 ad=3.25215 pd=20.04 as=7.6869 ps=40.2 w=19.71 l=1.14
X6 VDD2.t1 VN.t1 VTAIL.t10 w_n2146_n4910# sky130_fd_pr__pfet_01v8 ad=3.25215 pd=20.04 as=7.6869 ps=40.2 w=19.71 l=1.14
X7 VTAIL.t9 VN.t2 VDD2.t3 w_n2146_n4910# sky130_fd_pr__pfet_01v8 ad=3.25215 pd=20.04 as=3.25215 ps=20.04 w=19.71 l=1.14
X8 VDD2.t4 VN.t3 VTAIL.t8 w_n2146_n4910# sky130_fd_pr__pfet_01v8 ad=7.6869 pd=40.2 as=3.25215 ps=20.04 w=19.71 l=1.14
X9 B.t2 B.t0 B.t1 w_n2146_n4910# sky130_fd_pr__pfet_01v8 ad=7.6869 pd=40.2 as=0 ps=0 w=19.71 l=1.14
X10 VDD2.t0 VN.t4 VTAIL.t7 w_n2146_n4910# sky130_fd_pr__pfet_01v8 ad=7.6869 pd=40.2 as=3.25215 ps=20.04 w=19.71 l=1.14
X11 VDD1.t3 VP.t2 VTAIL.t0 w_n2146_n4910# sky130_fd_pr__pfet_01v8 ad=7.6869 pd=40.2 as=3.25215 ps=20.04 w=19.71 l=1.14
X12 VDD1.t2 VP.t3 VTAIL.t4 w_n2146_n4910# sky130_fd_pr__pfet_01v8 ad=7.6869 pd=40.2 as=3.25215 ps=20.04 w=19.71 l=1.14
X13 VTAIL.t1 VP.t4 VDD1.t1 w_n2146_n4910# sky130_fd_pr__pfet_01v8 ad=3.25215 pd=20.04 as=3.25215 ps=20.04 w=19.71 l=1.14
X14 VDD1.t0 VP.t5 VTAIL.t5 w_n2146_n4910# sky130_fd_pr__pfet_01v8 ad=3.25215 pd=20.04 as=7.6869 ps=40.2 w=19.71 l=1.14
X15 VDD2.t5 VN.t5 VTAIL.t6 w_n2146_n4910# sky130_fd_pr__pfet_01v8 ad=3.25215 pd=20.04 as=7.6869 ps=40.2 w=19.71 l=1.14
R0 VN.n1 VN.t4 474.664
R1 VN.n7 VN.t1 474.664
R2 VN.n4 VN.t5 451.346
R3 VN.n10 VN.t3 451.346
R4 VN.n2 VN.t0 416.676
R5 VN.n8 VN.t2 416.676
R6 VN.n9 VN.n6 161.3
R7 VN.n3 VN.n0 161.3
R8 VN.n11 VN.n10 80.6037
R9 VN.n5 VN.n4 80.6037
R10 VN.n4 VN.n3 51.6259
R11 VN.n10 VN.n9 51.6259
R12 VN VN.n11 49.3059
R13 VN.n2 VN.n1 32.927
R14 VN.n8 VN.n7 32.927
R15 VN.n7 VN.n6 27.9957
R16 VN.n1 VN.n0 27.9957
R17 VN.n3 VN.n2 24.4675
R18 VN.n9 VN.n8 24.4675
R19 VN.n11 VN.n6 0.285035
R20 VN.n5 VN.n0 0.285035
R21 VN VN.n5 0.146778
R22 VDD2.n215 VDD2.n111 756.745
R23 VDD2.n104 VDD2.n0 756.745
R24 VDD2.n216 VDD2.n215 585
R25 VDD2.n214 VDD2.n213 585
R26 VDD2.n115 VDD2.n114 585
R27 VDD2.n208 VDD2.n207 585
R28 VDD2.n206 VDD2.n205 585
R29 VDD2.n119 VDD2.n118 585
R30 VDD2.n200 VDD2.n199 585
R31 VDD2.n198 VDD2.n197 585
R32 VDD2.n123 VDD2.n122 585
R33 VDD2.n127 VDD2.n125 585
R34 VDD2.n192 VDD2.n191 585
R35 VDD2.n190 VDD2.n189 585
R36 VDD2.n129 VDD2.n128 585
R37 VDD2.n184 VDD2.n183 585
R38 VDD2.n182 VDD2.n181 585
R39 VDD2.n133 VDD2.n132 585
R40 VDD2.n176 VDD2.n175 585
R41 VDD2.n174 VDD2.n173 585
R42 VDD2.n137 VDD2.n136 585
R43 VDD2.n168 VDD2.n167 585
R44 VDD2.n166 VDD2.n165 585
R45 VDD2.n141 VDD2.n140 585
R46 VDD2.n160 VDD2.n159 585
R47 VDD2.n158 VDD2.n157 585
R48 VDD2.n145 VDD2.n144 585
R49 VDD2.n152 VDD2.n151 585
R50 VDD2.n150 VDD2.n149 585
R51 VDD2.n37 VDD2.n36 585
R52 VDD2.n39 VDD2.n38 585
R53 VDD2.n32 VDD2.n31 585
R54 VDD2.n45 VDD2.n44 585
R55 VDD2.n47 VDD2.n46 585
R56 VDD2.n28 VDD2.n27 585
R57 VDD2.n53 VDD2.n52 585
R58 VDD2.n55 VDD2.n54 585
R59 VDD2.n24 VDD2.n23 585
R60 VDD2.n61 VDD2.n60 585
R61 VDD2.n63 VDD2.n62 585
R62 VDD2.n20 VDD2.n19 585
R63 VDD2.n69 VDD2.n68 585
R64 VDD2.n71 VDD2.n70 585
R65 VDD2.n16 VDD2.n15 585
R66 VDD2.n78 VDD2.n77 585
R67 VDD2.n79 VDD2.n14 585
R68 VDD2.n81 VDD2.n80 585
R69 VDD2.n12 VDD2.n11 585
R70 VDD2.n87 VDD2.n86 585
R71 VDD2.n89 VDD2.n88 585
R72 VDD2.n8 VDD2.n7 585
R73 VDD2.n95 VDD2.n94 585
R74 VDD2.n97 VDD2.n96 585
R75 VDD2.n4 VDD2.n3 585
R76 VDD2.n103 VDD2.n102 585
R77 VDD2.n105 VDD2.n104 585
R78 VDD2.n148 VDD2.t4 327.466
R79 VDD2.n35 VDD2.t0 327.466
R80 VDD2.n215 VDD2.n214 171.744
R81 VDD2.n214 VDD2.n114 171.744
R82 VDD2.n207 VDD2.n114 171.744
R83 VDD2.n207 VDD2.n206 171.744
R84 VDD2.n206 VDD2.n118 171.744
R85 VDD2.n199 VDD2.n118 171.744
R86 VDD2.n199 VDD2.n198 171.744
R87 VDD2.n198 VDD2.n122 171.744
R88 VDD2.n127 VDD2.n122 171.744
R89 VDD2.n191 VDD2.n127 171.744
R90 VDD2.n191 VDD2.n190 171.744
R91 VDD2.n190 VDD2.n128 171.744
R92 VDD2.n183 VDD2.n128 171.744
R93 VDD2.n183 VDD2.n182 171.744
R94 VDD2.n182 VDD2.n132 171.744
R95 VDD2.n175 VDD2.n132 171.744
R96 VDD2.n175 VDD2.n174 171.744
R97 VDD2.n174 VDD2.n136 171.744
R98 VDD2.n167 VDD2.n136 171.744
R99 VDD2.n167 VDD2.n166 171.744
R100 VDD2.n166 VDD2.n140 171.744
R101 VDD2.n159 VDD2.n140 171.744
R102 VDD2.n159 VDD2.n158 171.744
R103 VDD2.n158 VDD2.n144 171.744
R104 VDD2.n151 VDD2.n144 171.744
R105 VDD2.n151 VDD2.n150 171.744
R106 VDD2.n38 VDD2.n37 171.744
R107 VDD2.n38 VDD2.n31 171.744
R108 VDD2.n45 VDD2.n31 171.744
R109 VDD2.n46 VDD2.n45 171.744
R110 VDD2.n46 VDD2.n27 171.744
R111 VDD2.n53 VDD2.n27 171.744
R112 VDD2.n54 VDD2.n53 171.744
R113 VDD2.n54 VDD2.n23 171.744
R114 VDD2.n61 VDD2.n23 171.744
R115 VDD2.n62 VDD2.n61 171.744
R116 VDD2.n62 VDD2.n19 171.744
R117 VDD2.n69 VDD2.n19 171.744
R118 VDD2.n70 VDD2.n69 171.744
R119 VDD2.n70 VDD2.n15 171.744
R120 VDD2.n78 VDD2.n15 171.744
R121 VDD2.n79 VDD2.n78 171.744
R122 VDD2.n80 VDD2.n79 171.744
R123 VDD2.n80 VDD2.n11 171.744
R124 VDD2.n87 VDD2.n11 171.744
R125 VDD2.n88 VDD2.n87 171.744
R126 VDD2.n88 VDD2.n7 171.744
R127 VDD2.n95 VDD2.n7 171.744
R128 VDD2.n96 VDD2.n95 171.744
R129 VDD2.n96 VDD2.n3 171.744
R130 VDD2.n103 VDD2.n3 171.744
R131 VDD2.n104 VDD2.n103 171.744
R132 VDD2.n150 VDD2.t4 85.8723
R133 VDD2.n37 VDD2.t0 85.8723
R134 VDD2.n110 VDD2.n109 68.9529
R135 VDD2 VDD2.n221 68.95
R136 VDD2.n110 VDD2.n108 50.341
R137 VDD2.n220 VDD2.n219 49.446
R138 VDD2.n220 VDD2.n110 44.8252
R139 VDD2.n149 VDD2.n148 16.3895
R140 VDD2.n36 VDD2.n35 16.3895
R141 VDD2.n125 VDD2.n123 13.1884
R142 VDD2.n81 VDD2.n12 13.1884
R143 VDD2.n197 VDD2.n196 12.8005
R144 VDD2.n193 VDD2.n192 12.8005
R145 VDD2.n152 VDD2.n147 12.8005
R146 VDD2.n39 VDD2.n34 12.8005
R147 VDD2.n82 VDD2.n14 12.8005
R148 VDD2.n86 VDD2.n85 12.8005
R149 VDD2.n200 VDD2.n121 12.0247
R150 VDD2.n189 VDD2.n126 12.0247
R151 VDD2.n153 VDD2.n145 12.0247
R152 VDD2.n40 VDD2.n32 12.0247
R153 VDD2.n77 VDD2.n76 12.0247
R154 VDD2.n89 VDD2.n10 12.0247
R155 VDD2.n201 VDD2.n119 11.249
R156 VDD2.n188 VDD2.n129 11.249
R157 VDD2.n157 VDD2.n156 11.249
R158 VDD2.n44 VDD2.n43 11.249
R159 VDD2.n75 VDD2.n16 11.249
R160 VDD2.n90 VDD2.n8 11.249
R161 VDD2.n205 VDD2.n204 10.4732
R162 VDD2.n185 VDD2.n184 10.4732
R163 VDD2.n160 VDD2.n143 10.4732
R164 VDD2.n47 VDD2.n30 10.4732
R165 VDD2.n72 VDD2.n71 10.4732
R166 VDD2.n94 VDD2.n93 10.4732
R167 VDD2.n208 VDD2.n117 9.69747
R168 VDD2.n181 VDD2.n131 9.69747
R169 VDD2.n161 VDD2.n141 9.69747
R170 VDD2.n48 VDD2.n28 9.69747
R171 VDD2.n68 VDD2.n18 9.69747
R172 VDD2.n97 VDD2.n6 9.69747
R173 VDD2.n219 VDD2.n218 9.45567
R174 VDD2.n108 VDD2.n107 9.45567
R175 VDD2.n135 VDD2.n134 9.3005
R176 VDD2.n178 VDD2.n177 9.3005
R177 VDD2.n180 VDD2.n179 9.3005
R178 VDD2.n131 VDD2.n130 9.3005
R179 VDD2.n186 VDD2.n185 9.3005
R180 VDD2.n188 VDD2.n187 9.3005
R181 VDD2.n126 VDD2.n124 9.3005
R182 VDD2.n194 VDD2.n193 9.3005
R183 VDD2.n218 VDD2.n217 9.3005
R184 VDD2.n113 VDD2.n112 9.3005
R185 VDD2.n212 VDD2.n211 9.3005
R186 VDD2.n210 VDD2.n209 9.3005
R187 VDD2.n117 VDD2.n116 9.3005
R188 VDD2.n204 VDD2.n203 9.3005
R189 VDD2.n202 VDD2.n201 9.3005
R190 VDD2.n121 VDD2.n120 9.3005
R191 VDD2.n196 VDD2.n195 9.3005
R192 VDD2.n172 VDD2.n171 9.3005
R193 VDD2.n170 VDD2.n169 9.3005
R194 VDD2.n139 VDD2.n138 9.3005
R195 VDD2.n164 VDD2.n163 9.3005
R196 VDD2.n162 VDD2.n161 9.3005
R197 VDD2.n143 VDD2.n142 9.3005
R198 VDD2.n156 VDD2.n155 9.3005
R199 VDD2.n154 VDD2.n153 9.3005
R200 VDD2.n147 VDD2.n146 9.3005
R201 VDD2.n107 VDD2.n106 9.3005
R202 VDD2.n101 VDD2.n100 9.3005
R203 VDD2.n99 VDD2.n98 9.3005
R204 VDD2.n6 VDD2.n5 9.3005
R205 VDD2.n93 VDD2.n92 9.3005
R206 VDD2.n91 VDD2.n90 9.3005
R207 VDD2.n10 VDD2.n9 9.3005
R208 VDD2.n85 VDD2.n84 9.3005
R209 VDD2.n57 VDD2.n56 9.3005
R210 VDD2.n26 VDD2.n25 9.3005
R211 VDD2.n51 VDD2.n50 9.3005
R212 VDD2.n49 VDD2.n48 9.3005
R213 VDD2.n30 VDD2.n29 9.3005
R214 VDD2.n43 VDD2.n42 9.3005
R215 VDD2.n41 VDD2.n40 9.3005
R216 VDD2.n34 VDD2.n33 9.3005
R217 VDD2.n59 VDD2.n58 9.3005
R218 VDD2.n22 VDD2.n21 9.3005
R219 VDD2.n65 VDD2.n64 9.3005
R220 VDD2.n67 VDD2.n66 9.3005
R221 VDD2.n18 VDD2.n17 9.3005
R222 VDD2.n73 VDD2.n72 9.3005
R223 VDD2.n75 VDD2.n74 9.3005
R224 VDD2.n76 VDD2.n13 9.3005
R225 VDD2.n83 VDD2.n82 9.3005
R226 VDD2.n2 VDD2.n1 9.3005
R227 VDD2.n209 VDD2.n115 8.92171
R228 VDD2.n180 VDD2.n133 8.92171
R229 VDD2.n165 VDD2.n164 8.92171
R230 VDD2.n52 VDD2.n51 8.92171
R231 VDD2.n67 VDD2.n20 8.92171
R232 VDD2.n98 VDD2.n4 8.92171
R233 VDD2.n213 VDD2.n212 8.14595
R234 VDD2.n177 VDD2.n176 8.14595
R235 VDD2.n168 VDD2.n139 8.14595
R236 VDD2.n55 VDD2.n26 8.14595
R237 VDD2.n64 VDD2.n63 8.14595
R238 VDD2.n102 VDD2.n101 8.14595
R239 VDD2.n219 VDD2.n111 7.3702
R240 VDD2.n216 VDD2.n113 7.3702
R241 VDD2.n173 VDD2.n135 7.3702
R242 VDD2.n169 VDD2.n137 7.3702
R243 VDD2.n56 VDD2.n24 7.3702
R244 VDD2.n60 VDD2.n22 7.3702
R245 VDD2.n105 VDD2.n2 7.3702
R246 VDD2.n108 VDD2.n0 7.3702
R247 VDD2.n217 VDD2.n111 6.59444
R248 VDD2.n217 VDD2.n216 6.59444
R249 VDD2.n173 VDD2.n172 6.59444
R250 VDD2.n172 VDD2.n137 6.59444
R251 VDD2.n59 VDD2.n24 6.59444
R252 VDD2.n60 VDD2.n59 6.59444
R253 VDD2.n106 VDD2.n105 6.59444
R254 VDD2.n106 VDD2.n0 6.59444
R255 VDD2.n213 VDD2.n113 5.81868
R256 VDD2.n176 VDD2.n135 5.81868
R257 VDD2.n169 VDD2.n168 5.81868
R258 VDD2.n56 VDD2.n55 5.81868
R259 VDD2.n63 VDD2.n22 5.81868
R260 VDD2.n102 VDD2.n2 5.81868
R261 VDD2.n212 VDD2.n115 5.04292
R262 VDD2.n177 VDD2.n133 5.04292
R263 VDD2.n165 VDD2.n139 5.04292
R264 VDD2.n52 VDD2.n26 5.04292
R265 VDD2.n64 VDD2.n20 5.04292
R266 VDD2.n101 VDD2.n4 5.04292
R267 VDD2.n209 VDD2.n208 4.26717
R268 VDD2.n181 VDD2.n180 4.26717
R269 VDD2.n164 VDD2.n141 4.26717
R270 VDD2.n51 VDD2.n28 4.26717
R271 VDD2.n68 VDD2.n67 4.26717
R272 VDD2.n98 VDD2.n97 4.26717
R273 VDD2.n148 VDD2.n146 3.70982
R274 VDD2.n35 VDD2.n33 3.70982
R275 VDD2.n205 VDD2.n117 3.49141
R276 VDD2.n184 VDD2.n131 3.49141
R277 VDD2.n161 VDD2.n160 3.49141
R278 VDD2.n48 VDD2.n47 3.49141
R279 VDD2.n71 VDD2.n18 3.49141
R280 VDD2.n94 VDD2.n6 3.49141
R281 VDD2.n204 VDD2.n119 2.71565
R282 VDD2.n185 VDD2.n129 2.71565
R283 VDD2.n157 VDD2.n143 2.71565
R284 VDD2.n44 VDD2.n30 2.71565
R285 VDD2.n72 VDD2.n16 2.71565
R286 VDD2.n93 VDD2.n8 2.71565
R287 VDD2.n201 VDD2.n200 1.93989
R288 VDD2.n189 VDD2.n188 1.93989
R289 VDD2.n156 VDD2.n145 1.93989
R290 VDD2.n43 VDD2.n32 1.93989
R291 VDD2.n77 VDD2.n75 1.93989
R292 VDD2.n90 VDD2.n89 1.93989
R293 VDD2.n221 VDD2.t3 1.64966
R294 VDD2.n221 VDD2.t1 1.64966
R295 VDD2.n109 VDD2.t2 1.64966
R296 VDD2.n109 VDD2.t5 1.64966
R297 VDD2.n197 VDD2.n121 1.16414
R298 VDD2.n192 VDD2.n126 1.16414
R299 VDD2.n153 VDD2.n152 1.16414
R300 VDD2.n40 VDD2.n39 1.16414
R301 VDD2.n76 VDD2.n14 1.16414
R302 VDD2.n86 VDD2.n10 1.16414
R303 VDD2 VDD2.n220 1.00912
R304 VDD2.n196 VDD2.n123 0.388379
R305 VDD2.n193 VDD2.n125 0.388379
R306 VDD2.n149 VDD2.n147 0.388379
R307 VDD2.n36 VDD2.n34 0.388379
R308 VDD2.n82 VDD2.n81 0.388379
R309 VDD2.n85 VDD2.n12 0.388379
R310 VDD2.n218 VDD2.n112 0.155672
R311 VDD2.n211 VDD2.n112 0.155672
R312 VDD2.n211 VDD2.n210 0.155672
R313 VDD2.n210 VDD2.n116 0.155672
R314 VDD2.n203 VDD2.n116 0.155672
R315 VDD2.n203 VDD2.n202 0.155672
R316 VDD2.n202 VDD2.n120 0.155672
R317 VDD2.n195 VDD2.n120 0.155672
R318 VDD2.n195 VDD2.n194 0.155672
R319 VDD2.n194 VDD2.n124 0.155672
R320 VDD2.n187 VDD2.n124 0.155672
R321 VDD2.n187 VDD2.n186 0.155672
R322 VDD2.n186 VDD2.n130 0.155672
R323 VDD2.n179 VDD2.n130 0.155672
R324 VDD2.n179 VDD2.n178 0.155672
R325 VDD2.n178 VDD2.n134 0.155672
R326 VDD2.n171 VDD2.n134 0.155672
R327 VDD2.n171 VDD2.n170 0.155672
R328 VDD2.n170 VDD2.n138 0.155672
R329 VDD2.n163 VDD2.n138 0.155672
R330 VDD2.n163 VDD2.n162 0.155672
R331 VDD2.n162 VDD2.n142 0.155672
R332 VDD2.n155 VDD2.n142 0.155672
R333 VDD2.n155 VDD2.n154 0.155672
R334 VDD2.n154 VDD2.n146 0.155672
R335 VDD2.n41 VDD2.n33 0.155672
R336 VDD2.n42 VDD2.n41 0.155672
R337 VDD2.n42 VDD2.n29 0.155672
R338 VDD2.n49 VDD2.n29 0.155672
R339 VDD2.n50 VDD2.n49 0.155672
R340 VDD2.n50 VDD2.n25 0.155672
R341 VDD2.n57 VDD2.n25 0.155672
R342 VDD2.n58 VDD2.n57 0.155672
R343 VDD2.n58 VDD2.n21 0.155672
R344 VDD2.n65 VDD2.n21 0.155672
R345 VDD2.n66 VDD2.n65 0.155672
R346 VDD2.n66 VDD2.n17 0.155672
R347 VDD2.n73 VDD2.n17 0.155672
R348 VDD2.n74 VDD2.n73 0.155672
R349 VDD2.n74 VDD2.n13 0.155672
R350 VDD2.n83 VDD2.n13 0.155672
R351 VDD2.n84 VDD2.n83 0.155672
R352 VDD2.n84 VDD2.n9 0.155672
R353 VDD2.n91 VDD2.n9 0.155672
R354 VDD2.n92 VDD2.n91 0.155672
R355 VDD2.n92 VDD2.n5 0.155672
R356 VDD2.n99 VDD2.n5 0.155672
R357 VDD2.n100 VDD2.n99 0.155672
R358 VDD2.n100 VDD2.n1 0.155672
R359 VDD2.n107 VDD2.n1 0.155672
R360 VTAIL.n442 VTAIL.n338 756.745
R361 VTAIL.n106 VTAIL.n2 756.745
R362 VTAIL.n332 VTAIL.n228 756.745
R363 VTAIL.n220 VTAIL.n116 756.745
R364 VTAIL.n375 VTAIL.n374 585
R365 VTAIL.n377 VTAIL.n376 585
R366 VTAIL.n370 VTAIL.n369 585
R367 VTAIL.n383 VTAIL.n382 585
R368 VTAIL.n385 VTAIL.n384 585
R369 VTAIL.n366 VTAIL.n365 585
R370 VTAIL.n391 VTAIL.n390 585
R371 VTAIL.n393 VTAIL.n392 585
R372 VTAIL.n362 VTAIL.n361 585
R373 VTAIL.n399 VTAIL.n398 585
R374 VTAIL.n401 VTAIL.n400 585
R375 VTAIL.n358 VTAIL.n357 585
R376 VTAIL.n407 VTAIL.n406 585
R377 VTAIL.n409 VTAIL.n408 585
R378 VTAIL.n354 VTAIL.n353 585
R379 VTAIL.n416 VTAIL.n415 585
R380 VTAIL.n417 VTAIL.n352 585
R381 VTAIL.n419 VTAIL.n418 585
R382 VTAIL.n350 VTAIL.n349 585
R383 VTAIL.n425 VTAIL.n424 585
R384 VTAIL.n427 VTAIL.n426 585
R385 VTAIL.n346 VTAIL.n345 585
R386 VTAIL.n433 VTAIL.n432 585
R387 VTAIL.n435 VTAIL.n434 585
R388 VTAIL.n342 VTAIL.n341 585
R389 VTAIL.n441 VTAIL.n440 585
R390 VTAIL.n443 VTAIL.n442 585
R391 VTAIL.n39 VTAIL.n38 585
R392 VTAIL.n41 VTAIL.n40 585
R393 VTAIL.n34 VTAIL.n33 585
R394 VTAIL.n47 VTAIL.n46 585
R395 VTAIL.n49 VTAIL.n48 585
R396 VTAIL.n30 VTAIL.n29 585
R397 VTAIL.n55 VTAIL.n54 585
R398 VTAIL.n57 VTAIL.n56 585
R399 VTAIL.n26 VTAIL.n25 585
R400 VTAIL.n63 VTAIL.n62 585
R401 VTAIL.n65 VTAIL.n64 585
R402 VTAIL.n22 VTAIL.n21 585
R403 VTAIL.n71 VTAIL.n70 585
R404 VTAIL.n73 VTAIL.n72 585
R405 VTAIL.n18 VTAIL.n17 585
R406 VTAIL.n80 VTAIL.n79 585
R407 VTAIL.n81 VTAIL.n16 585
R408 VTAIL.n83 VTAIL.n82 585
R409 VTAIL.n14 VTAIL.n13 585
R410 VTAIL.n89 VTAIL.n88 585
R411 VTAIL.n91 VTAIL.n90 585
R412 VTAIL.n10 VTAIL.n9 585
R413 VTAIL.n97 VTAIL.n96 585
R414 VTAIL.n99 VTAIL.n98 585
R415 VTAIL.n6 VTAIL.n5 585
R416 VTAIL.n105 VTAIL.n104 585
R417 VTAIL.n107 VTAIL.n106 585
R418 VTAIL.n333 VTAIL.n332 585
R419 VTAIL.n331 VTAIL.n330 585
R420 VTAIL.n232 VTAIL.n231 585
R421 VTAIL.n325 VTAIL.n324 585
R422 VTAIL.n323 VTAIL.n322 585
R423 VTAIL.n236 VTAIL.n235 585
R424 VTAIL.n317 VTAIL.n316 585
R425 VTAIL.n315 VTAIL.n314 585
R426 VTAIL.n240 VTAIL.n239 585
R427 VTAIL.n244 VTAIL.n242 585
R428 VTAIL.n309 VTAIL.n308 585
R429 VTAIL.n307 VTAIL.n306 585
R430 VTAIL.n246 VTAIL.n245 585
R431 VTAIL.n301 VTAIL.n300 585
R432 VTAIL.n299 VTAIL.n298 585
R433 VTAIL.n250 VTAIL.n249 585
R434 VTAIL.n293 VTAIL.n292 585
R435 VTAIL.n291 VTAIL.n290 585
R436 VTAIL.n254 VTAIL.n253 585
R437 VTAIL.n285 VTAIL.n284 585
R438 VTAIL.n283 VTAIL.n282 585
R439 VTAIL.n258 VTAIL.n257 585
R440 VTAIL.n277 VTAIL.n276 585
R441 VTAIL.n275 VTAIL.n274 585
R442 VTAIL.n262 VTAIL.n261 585
R443 VTAIL.n269 VTAIL.n268 585
R444 VTAIL.n267 VTAIL.n266 585
R445 VTAIL.n221 VTAIL.n220 585
R446 VTAIL.n219 VTAIL.n218 585
R447 VTAIL.n120 VTAIL.n119 585
R448 VTAIL.n213 VTAIL.n212 585
R449 VTAIL.n211 VTAIL.n210 585
R450 VTAIL.n124 VTAIL.n123 585
R451 VTAIL.n205 VTAIL.n204 585
R452 VTAIL.n203 VTAIL.n202 585
R453 VTAIL.n128 VTAIL.n127 585
R454 VTAIL.n132 VTAIL.n130 585
R455 VTAIL.n197 VTAIL.n196 585
R456 VTAIL.n195 VTAIL.n194 585
R457 VTAIL.n134 VTAIL.n133 585
R458 VTAIL.n189 VTAIL.n188 585
R459 VTAIL.n187 VTAIL.n186 585
R460 VTAIL.n138 VTAIL.n137 585
R461 VTAIL.n181 VTAIL.n180 585
R462 VTAIL.n179 VTAIL.n178 585
R463 VTAIL.n142 VTAIL.n141 585
R464 VTAIL.n173 VTAIL.n172 585
R465 VTAIL.n171 VTAIL.n170 585
R466 VTAIL.n146 VTAIL.n145 585
R467 VTAIL.n165 VTAIL.n164 585
R468 VTAIL.n163 VTAIL.n162 585
R469 VTAIL.n150 VTAIL.n149 585
R470 VTAIL.n157 VTAIL.n156 585
R471 VTAIL.n155 VTAIL.n154 585
R472 VTAIL.n373 VTAIL.t6 327.466
R473 VTAIL.n37 VTAIL.t3 327.466
R474 VTAIL.n265 VTAIL.t5 327.466
R475 VTAIL.n153 VTAIL.t10 327.466
R476 VTAIL.n376 VTAIL.n375 171.744
R477 VTAIL.n376 VTAIL.n369 171.744
R478 VTAIL.n383 VTAIL.n369 171.744
R479 VTAIL.n384 VTAIL.n383 171.744
R480 VTAIL.n384 VTAIL.n365 171.744
R481 VTAIL.n391 VTAIL.n365 171.744
R482 VTAIL.n392 VTAIL.n391 171.744
R483 VTAIL.n392 VTAIL.n361 171.744
R484 VTAIL.n399 VTAIL.n361 171.744
R485 VTAIL.n400 VTAIL.n399 171.744
R486 VTAIL.n400 VTAIL.n357 171.744
R487 VTAIL.n407 VTAIL.n357 171.744
R488 VTAIL.n408 VTAIL.n407 171.744
R489 VTAIL.n408 VTAIL.n353 171.744
R490 VTAIL.n416 VTAIL.n353 171.744
R491 VTAIL.n417 VTAIL.n416 171.744
R492 VTAIL.n418 VTAIL.n417 171.744
R493 VTAIL.n418 VTAIL.n349 171.744
R494 VTAIL.n425 VTAIL.n349 171.744
R495 VTAIL.n426 VTAIL.n425 171.744
R496 VTAIL.n426 VTAIL.n345 171.744
R497 VTAIL.n433 VTAIL.n345 171.744
R498 VTAIL.n434 VTAIL.n433 171.744
R499 VTAIL.n434 VTAIL.n341 171.744
R500 VTAIL.n441 VTAIL.n341 171.744
R501 VTAIL.n442 VTAIL.n441 171.744
R502 VTAIL.n40 VTAIL.n39 171.744
R503 VTAIL.n40 VTAIL.n33 171.744
R504 VTAIL.n47 VTAIL.n33 171.744
R505 VTAIL.n48 VTAIL.n47 171.744
R506 VTAIL.n48 VTAIL.n29 171.744
R507 VTAIL.n55 VTAIL.n29 171.744
R508 VTAIL.n56 VTAIL.n55 171.744
R509 VTAIL.n56 VTAIL.n25 171.744
R510 VTAIL.n63 VTAIL.n25 171.744
R511 VTAIL.n64 VTAIL.n63 171.744
R512 VTAIL.n64 VTAIL.n21 171.744
R513 VTAIL.n71 VTAIL.n21 171.744
R514 VTAIL.n72 VTAIL.n71 171.744
R515 VTAIL.n72 VTAIL.n17 171.744
R516 VTAIL.n80 VTAIL.n17 171.744
R517 VTAIL.n81 VTAIL.n80 171.744
R518 VTAIL.n82 VTAIL.n81 171.744
R519 VTAIL.n82 VTAIL.n13 171.744
R520 VTAIL.n89 VTAIL.n13 171.744
R521 VTAIL.n90 VTAIL.n89 171.744
R522 VTAIL.n90 VTAIL.n9 171.744
R523 VTAIL.n97 VTAIL.n9 171.744
R524 VTAIL.n98 VTAIL.n97 171.744
R525 VTAIL.n98 VTAIL.n5 171.744
R526 VTAIL.n105 VTAIL.n5 171.744
R527 VTAIL.n106 VTAIL.n105 171.744
R528 VTAIL.n332 VTAIL.n331 171.744
R529 VTAIL.n331 VTAIL.n231 171.744
R530 VTAIL.n324 VTAIL.n231 171.744
R531 VTAIL.n324 VTAIL.n323 171.744
R532 VTAIL.n323 VTAIL.n235 171.744
R533 VTAIL.n316 VTAIL.n235 171.744
R534 VTAIL.n316 VTAIL.n315 171.744
R535 VTAIL.n315 VTAIL.n239 171.744
R536 VTAIL.n244 VTAIL.n239 171.744
R537 VTAIL.n308 VTAIL.n244 171.744
R538 VTAIL.n308 VTAIL.n307 171.744
R539 VTAIL.n307 VTAIL.n245 171.744
R540 VTAIL.n300 VTAIL.n245 171.744
R541 VTAIL.n300 VTAIL.n299 171.744
R542 VTAIL.n299 VTAIL.n249 171.744
R543 VTAIL.n292 VTAIL.n249 171.744
R544 VTAIL.n292 VTAIL.n291 171.744
R545 VTAIL.n291 VTAIL.n253 171.744
R546 VTAIL.n284 VTAIL.n253 171.744
R547 VTAIL.n284 VTAIL.n283 171.744
R548 VTAIL.n283 VTAIL.n257 171.744
R549 VTAIL.n276 VTAIL.n257 171.744
R550 VTAIL.n276 VTAIL.n275 171.744
R551 VTAIL.n275 VTAIL.n261 171.744
R552 VTAIL.n268 VTAIL.n261 171.744
R553 VTAIL.n268 VTAIL.n267 171.744
R554 VTAIL.n220 VTAIL.n219 171.744
R555 VTAIL.n219 VTAIL.n119 171.744
R556 VTAIL.n212 VTAIL.n119 171.744
R557 VTAIL.n212 VTAIL.n211 171.744
R558 VTAIL.n211 VTAIL.n123 171.744
R559 VTAIL.n204 VTAIL.n123 171.744
R560 VTAIL.n204 VTAIL.n203 171.744
R561 VTAIL.n203 VTAIL.n127 171.744
R562 VTAIL.n132 VTAIL.n127 171.744
R563 VTAIL.n196 VTAIL.n132 171.744
R564 VTAIL.n196 VTAIL.n195 171.744
R565 VTAIL.n195 VTAIL.n133 171.744
R566 VTAIL.n188 VTAIL.n133 171.744
R567 VTAIL.n188 VTAIL.n187 171.744
R568 VTAIL.n187 VTAIL.n137 171.744
R569 VTAIL.n180 VTAIL.n137 171.744
R570 VTAIL.n180 VTAIL.n179 171.744
R571 VTAIL.n179 VTAIL.n141 171.744
R572 VTAIL.n172 VTAIL.n141 171.744
R573 VTAIL.n172 VTAIL.n171 171.744
R574 VTAIL.n171 VTAIL.n145 171.744
R575 VTAIL.n164 VTAIL.n145 171.744
R576 VTAIL.n164 VTAIL.n163 171.744
R577 VTAIL.n163 VTAIL.n149 171.744
R578 VTAIL.n156 VTAIL.n149 171.744
R579 VTAIL.n156 VTAIL.n155 171.744
R580 VTAIL.n375 VTAIL.t6 85.8723
R581 VTAIL.n39 VTAIL.t3 85.8723
R582 VTAIL.n267 VTAIL.t5 85.8723
R583 VTAIL.n155 VTAIL.t10 85.8723
R584 VTAIL.n227 VTAIL.n226 52.0128
R585 VTAIL.n115 VTAIL.n114 52.0128
R586 VTAIL.n1 VTAIL.n0 52.0126
R587 VTAIL.n113 VTAIL.n112 52.0126
R588 VTAIL.n447 VTAIL.n446 32.7672
R589 VTAIL.n111 VTAIL.n110 32.7672
R590 VTAIL.n337 VTAIL.n336 32.7672
R591 VTAIL.n225 VTAIL.n224 32.7672
R592 VTAIL.n115 VTAIL.n113 31.8927
R593 VTAIL.n447 VTAIL.n337 30.6255
R594 VTAIL.n374 VTAIL.n373 16.3895
R595 VTAIL.n38 VTAIL.n37 16.3895
R596 VTAIL.n266 VTAIL.n265 16.3895
R597 VTAIL.n154 VTAIL.n153 16.3895
R598 VTAIL.n419 VTAIL.n350 13.1884
R599 VTAIL.n83 VTAIL.n14 13.1884
R600 VTAIL.n242 VTAIL.n240 13.1884
R601 VTAIL.n130 VTAIL.n128 13.1884
R602 VTAIL.n377 VTAIL.n372 12.8005
R603 VTAIL.n420 VTAIL.n352 12.8005
R604 VTAIL.n424 VTAIL.n423 12.8005
R605 VTAIL.n41 VTAIL.n36 12.8005
R606 VTAIL.n84 VTAIL.n16 12.8005
R607 VTAIL.n88 VTAIL.n87 12.8005
R608 VTAIL.n314 VTAIL.n313 12.8005
R609 VTAIL.n310 VTAIL.n309 12.8005
R610 VTAIL.n269 VTAIL.n264 12.8005
R611 VTAIL.n202 VTAIL.n201 12.8005
R612 VTAIL.n198 VTAIL.n197 12.8005
R613 VTAIL.n157 VTAIL.n152 12.8005
R614 VTAIL.n378 VTAIL.n370 12.0247
R615 VTAIL.n415 VTAIL.n414 12.0247
R616 VTAIL.n427 VTAIL.n348 12.0247
R617 VTAIL.n42 VTAIL.n34 12.0247
R618 VTAIL.n79 VTAIL.n78 12.0247
R619 VTAIL.n91 VTAIL.n12 12.0247
R620 VTAIL.n317 VTAIL.n238 12.0247
R621 VTAIL.n306 VTAIL.n243 12.0247
R622 VTAIL.n270 VTAIL.n262 12.0247
R623 VTAIL.n205 VTAIL.n126 12.0247
R624 VTAIL.n194 VTAIL.n131 12.0247
R625 VTAIL.n158 VTAIL.n150 12.0247
R626 VTAIL.n382 VTAIL.n381 11.249
R627 VTAIL.n413 VTAIL.n354 11.249
R628 VTAIL.n428 VTAIL.n346 11.249
R629 VTAIL.n46 VTAIL.n45 11.249
R630 VTAIL.n77 VTAIL.n18 11.249
R631 VTAIL.n92 VTAIL.n10 11.249
R632 VTAIL.n318 VTAIL.n236 11.249
R633 VTAIL.n305 VTAIL.n246 11.249
R634 VTAIL.n274 VTAIL.n273 11.249
R635 VTAIL.n206 VTAIL.n124 11.249
R636 VTAIL.n193 VTAIL.n134 11.249
R637 VTAIL.n162 VTAIL.n161 11.249
R638 VTAIL.n385 VTAIL.n368 10.4732
R639 VTAIL.n410 VTAIL.n409 10.4732
R640 VTAIL.n432 VTAIL.n431 10.4732
R641 VTAIL.n49 VTAIL.n32 10.4732
R642 VTAIL.n74 VTAIL.n73 10.4732
R643 VTAIL.n96 VTAIL.n95 10.4732
R644 VTAIL.n322 VTAIL.n321 10.4732
R645 VTAIL.n302 VTAIL.n301 10.4732
R646 VTAIL.n277 VTAIL.n260 10.4732
R647 VTAIL.n210 VTAIL.n209 10.4732
R648 VTAIL.n190 VTAIL.n189 10.4732
R649 VTAIL.n165 VTAIL.n148 10.4732
R650 VTAIL.n386 VTAIL.n366 9.69747
R651 VTAIL.n406 VTAIL.n356 9.69747
R652 VTAIL.n435 VTAIL.n344 9.69747
R653 VTAIL.n50 VTAIL.n30 9.69747
R654 VTAIL.n70 VTAIL.n20 9.69747
R655 VTAIL.n99 VTAIL.n8 9.69747
R656 VTAIL.n325 VTAIL.n234 9.69747
R657 VTAIL.n298 VTAIL.n248 9.69747
R658 VTAIL.n278 VTAIL.n258 9.69747
R659 VTAIL.n213 VTAIL.n122 9.69747
R660 VTAIL.n186 VTAIL.n136 9.69747
R661 VTAIL.n166 VTAIL.n146 9.69747
R662 VTAIL.n446 VTAIL.n445 9.45567
R663 VTAIL.n110 VTAIL.n109 9.45567
R664 VTAIL.n336 VTAIL.n335 9.45567
R665 VTAIL.n224 VTAIL.n223 9.45567
R666 VTAIL.n445 VTAIL.n444 9.3005
R667 VTAIL.n439 VTAIL.n438 9.3005
R668 VTAIL.n437 VTAIL.n436 9.3005
R669 VTAIL.n344 VTAIL.n343 9.3005
R670 VTAIL.n431 VTAIL.n430 9.3005
R671 VTAIL.n429 VTAIL.n428 9.3005
R672 VTAIL.n348 VTAIL.n347 9.3005
R673 VTAIL.n423 VTAIL.n422 9.3005
R674 VTAIL.n395 VTAIL.n394 9.3005
R675 VTAIL.n364 VTAIL.n363 9.3005
R676 VTAIL.n389 VTAIL.n388 9.3005
R677 VTAIL.n387 VTAIL.n386 9.3005
R678 VTAIL.n368 VTAIL.n367 9.3005
R679 VTAIL.n381 VTAIL.n380 9.3005
R680 VTAIL.n379 VTAIL.n378 9.3005
R681 VTAIL.n372 VTAIL.n371 9.3005
R682 VTAIL.n397 VTAIL.n396 9.3005
R683 VTAIL.n360 VTAIL.n359 9.3005
R684 VTAIL.n403 VTAIL.n402 9.3005
R685 VTAIL.n405 VTAIL.n404 9.3005
R686 VTAIL.n356 VTAIL.n355 9.3005
R687 VTAIL.n411 VTAIL.n410 9.3005
R688 VTAIL.n413 VTAIL.n412 9.3005
R689 VTAIL.n414 VTAIL.n351 9.3005
R690 VTAIL.n421 VTAIL.n420 9.3005
R691 VTAIL.n340 VTAIL.n339 9.3005
R692 VTAIL.n109 VTAIL.n108 9.3005
R693 VTAIL.n103 VTAIL.n102 9.3005
R694 VTAIL.n101 VTAIL.n100 9.3005
R695 VTAIL.n8 VTAIL.n7 9.3005
R696 VTAIL.n95 VTAIL.n94 9.3005
R697 VTAIL.n93 VTAIL.n92 9.3005
R698 VTAIL.n12 VTAIL.n11 9.3005
R699 VTAIL.n87 VTAIL.n86 9.3005
R700 VTAIL.n59 VTAIL.n58 9.3005
R701 VTAIL.n28 VTAIL.n27 9.3005
R702 VTAIL.n53 VTAIL.n52 9.3005
R703 VTAIL.n51 VTAIL.n50 9.3005
R704 VTAIL.n32 VTAIL.n31 9.3005
R705 VTAIL.n45 VTAIL.n44 9.3005
R706 VTAIL.n43 VTAIL.n42 9.3005
R707 VTAIL.n36 VTAIL.n35 9.3005
R708 VTAIL.n61 VTAIL.n60 9.3005
R709 VTAIL.n24 VTAIL.n23 9.3005
R710 VTAIL.n67 VTAIL.n66 9.3005
R711 VTAIL.n69 VTAIL.n68 9.3005
R712 VTAIL.n20 VTAIL.n19 9.3005
R713 VTAIL.n75 VTAIL.n74 9.3005
R714 VTAIL.n77 VTAIL.n76 9.3005
R715 VTAIL.n78 VTAIL.n15 9.3005
R716 VTAIL.n85 VTAIL.n84 9.3005
R717 VTAIL.n4 VTAIL.n3 9.3005
R718 VTAIL.n252 VTAIL.n251 9.3005
R719 VTAIL.n295 VTAIL.n294 9.3005
R720 VTAIL.n297 VTAIL.n296 9.3005
R721 VTAIL.n248 VTAIL.n247 9.3005
R722 VTAIL.n303 VTAIL.n302 9.3005
R723 VTAIL.n305 VTAIL.n304 9.3005
R724 VTAIL.n243 VTAIL.n241 9.3005
R725 VTAIL.n311 VTAIL.n310 9.3005
R726 VTAIL.n335 VTAIL.n334 9.3005
R727 VTAIL.n230 VTAIL.n229 9.3005
R728 VTAIL.n329 VTAIL.n328 9.3005
R729 VTAIL.n327 VTAIL.n326 9.3005
R730 VTAIL.n234 VTAIL.n233 9.3005
R731 VTAIL.n321 VTAIL.n320 9.3005
R732 VTAIL.n319 VTAIL.n318 9.3005
R733 VTAIL.n238 VTAIL.n237 9.3005
R734 VTAIL.n313 VTAIL.n312 9.3005
R735 VTAIL.n289 VTAIL.n288 9.3005
R736 VTAIL.n287 VTAIL.n286 9.3005
R737 VTAIL.n256 VTAIL.n255 9.3005
R738 VTAIL.n281 VTAIL.n280 9.3005
R739 VTAIL.n279 VTAIL.n278 9.3005
R740 VTAIL.n260 VTAIL.n259 9.3005
R741 VTAIL.n273 VTAIL.n272 9.3005
R742 VTAIL.n271 VTAIL.n270 9.3005
R743 VTAIL.n264 VTAIL.n263 9.3005
R744 VTAIL.n140 VTAIL.n139 9.3005
R745 VTAIL.n183 VTAIL.n182 9.3005
R746 VTAIL.n185 VTAIL.n184 9.3005
R747 VTAIL.n136 VTAIL.n135 9.3005
R748 VTAIL.n191 VTAIL.n190 9.3005
R749 VTAIL.n193 VTAIL.n192 9.3005
R750 VTAIL.n131 VTAIL.n129 9.3005
R751 VTAIL.n199 VTAIL.n198 9.3005
R752 VTAIL.n223 VTAIL.n222 9.3005
R753 VTAIL.n118 VTAIL.n117 9.3005
R754 VTAIL.n217 VTAIL.n216 9.3005
R755 VTAIL.n215 VTAIL.n214 9.3005
R756 VTAIL.n122 VTAIL.n121 9.3005
R757 VTAIL.n209 VTAIL.n208 9.3005
R758 VTAIL.n207 VTAIL.n206 9.3005
R759 VTAIL.n126 VTAIL.n125 9.3005
R760 VTAIL.n201 VTAIL.n200 9.3005
R761 VTAIL.n177 VTAIL.n176 9.3005
R762 VTAIL.n175 VTAIL.n174 9.3005
R763 VTAIL.n144 VTAIL.n143 9.3005
R764 VTAIL.n169 VTAIL.n168 9.3005
R765 VTAIL.n167 VTAIL.n166 9.3005
R766 VTAIL.n148 VTAIL.n147 9.3005
R767 VTAIL.n161 VTAIL.n160 9.3005
R768 VTAIL.n159 VTAIL.n158 9.3005
R769 VTAIL.n152 VTAIL.n151 9.3005
R770 VTAIL.n390 VTAIL.n389 8.92171
R771 VTAIL.n405 VTAIL.n358 8.92171
R772 VTAIL.n436 VTAIL.n342 8.92171
R773 VTAIL.n54 VTAIL.n53 8.92171
R774 VTAIL.n69 VTAIL.n22 8.92171
R775 VTAIL.n100 VTAIL.n6 8.92171
R776 VTAIL.n326 VTAIL.n232 8.92171
R777 VTAIL.n297 VTAIL.n250 8.92171
R778 VTAIL.n282 VTAIL.n281 8.92171
R779 VTAIL.n214 VTAIL.n120 8.92171
R780 VTAIL.n185 VTAIL.n138 8.92171
R781 VTAIL.n170 VTAIL.n169 8.92171
R782 VTAIL.n393 VTAIL.n364 8.14595
R783 VTAIL.n402 VTAIL.n401 8.14595
R784 VTAIL.n440 VTAIL.n439 8.14595
R785 VTAIL.n57 VTAIL.n28 8.14595
R786 VTAIL.n66 VTAIL.n65 8.14595
R787 VTAIL.n104 VTAIL.n103 8.14595
R788 VTAIL.n330 VTAIL.n329 8.14595
R789 VTAIL.n294 VTAIL.n293 8.14595
R790 VTAIL.n285 VTAIL.n256 8.14595
R791 VTAIL.n218 VTAIL.n217 8.14595
R792 VTAIL.n182 VTAIL.n181 8.14595
R793 VTAIL.n173 VTAIL.n144 8.14595
R794 VTAIL.n394 VTAIL.n362 7.3702
R795 VTAIL.n398 VTAIL.n360 7.3702
R796 VTAIL.n443 VTAIL.n340 7.3702
R797 VTAIL.n446 VTAIL.n338 7.3702
R798 VTAIL.n58 VTAIL.n26 7.3702
R799 VTAIL.n62 VTAIL.n24 7.3702
R800 VTAIL.n107 VTAIL.n4 7.3702
R801 VTAIL.n110 VTAIL.n2 7.3702
R802 VTAIL.n336 VTAIL.n228 7.3702
R803 VTAIL.n333 VTAIL.n230 7.3702
R804 VTAIL.n290 VTAIL.n252 7.3702
R805 VTAIL.n286 VTAIL.n254 7.3702
R806 VTAIL.n224 VTAIL.n116 7.3702
R807 VTAIL.n221 VTAIL.n118 7.3702
R808 VTAIL.n178 VTAIL.n140 7.3702
R809 VTAIL.n174 VTAIL.n142 7.3702
R810 VTAIL.n397 VTAIL.n362 6.59444
R811 VTAIL.n398 VTAIL.n397 6.59444
R812 VTAIL.n444 VTAIL.n443 6.59444
R813 VTAIL.n444 VTAIL.n338 6.59444
R814 VTAIL.n61 VTAIL.n26 6.59444
R815 VTAIL.n62 VTAIL.n61 6.59444
R816 VTAIL.n108 VTAIL.n107 6.59444
R817 VTAIL.n108 VTAIL.n2 6.59444
R818 VTAIL.n334 VTAIL.n228 6.59444
R819 VTAIL.n334 VTAIL.n333 6.59444
R820 VTAIL.n290 VTAIL.n289 6.59444
R821 VTAIL.n289 VTAIL.n254 6.59444
R822 VTAIL.n222 VTAIL.n116 6.59444
R823 VTAIL.n222 VTAIL.n221 6.59444
R824 VTAIL.n178 VTAIL.n177 6.59444
R825 VTAIL.n177 VTAIL.n142 6.59444
R826 VTAIL.n394 VTAIL.n393 5.81868
R827 VTAIL.n401 VTAIL.n360 5.81868
R828 VTAIL.n440 VTAIL.n340 5.81868
R829 VTAIL.n58 VTAIL.n57 5.81868
R830 VTAIL.n65 VTAIL.n24 5.81868
R831 VTAIL.n104 VTAIL.n4 5.81868
R832 VTAIL.n330 VTAIL.n230 5.81868
R833 VTAIL.n293 VTAIL.n252 5.81868
R834 VTAIL.n286 VTAIL.n285 5.81868
R835 VTAIL.n218 VTAIL.n118 5.81868
R836 VTAIL.n181 VTAIL.n140 5.81868
R837 VTAIL.n174 VTAIL.n173 5.81868
R838 VTAIL.n390 VTAIL.n364 5.04292
R839 VTAIL.n402 VTAIL.n358 5.04292
R840 VTAIL.n439 VTAIL.n342 5.04292
R841 VTAIL.n54 VTAIL.n28 5.04292
R842 VTAIL.n66 VTAIL.n22 5.04292
R843 VTAIL.n103 VTAIL.n6 5.04292
R844 VTAIL.n329 VTAIL.n232 5.04292
R845 VTAIL.n294 VTAIL.n250 5.04292
R846 VTAIL.n282 VTAIL.n256 5.04292
R847 VTAIL.n217 VTAIL.n120 5.04292
R848 VTAIL.n182 VTAIL.n138 5.04292
R849 VTAIL.n170 VTAIL.n144 5.04292
R850 VTAIL.n389 VTAIL.n366 4.26717
R851 VTAIL.n406 VTAIL.n405 4.26717
R852 VTAIL.n436 VTAIL.n435 4.26717
R853 VTAIL.n53 VTAIL.n30 4.26717
R854 VTAIL.n70 VTAIL.n69 4.26717
R855 VTAIL.n100 VTAIL.n99 4.26717
R856 VTAIL.n326 VTAIL.n325 4.26717
R857 VTAIL.n298 VTAIL.n297 4.26717
R858 VTAIL.n281 VTAIL.n258 4.26717
R859 VTAIL.n214 VTAIL.n213 4.26717
R860 VTAIL.n186 VTAIL.n185 4.26717
R861 VTAIL.n169 VTAIL.n146 4.26717
R862 VTAIL.n373 VTAIL.n371 3.70982
R863 VTAIL.n37 VTAIL.n35 3.70982
R864 VTAIL.n265 VTAIL.n263 3.70982
R865 VTAIL.n153 VTAIL.n151 3.70982
R866 VTAIL.n386 VTAIL.n385 3.49141
R867 VTAIL.n409 VTAIL.n356 3.49141
R868 VTAIL.n432 VTAIL.n344 3.49141
R869 VTAIL.n50 VTAIL.n49 3.49141
R870 VTAIL.n73 VTAIL.n20 3.49141
R871 VTAIL.n96 VTAIL.n8 3.49141
R872 VTAIL.n322 VTAIL.n234 3.49141
R873 VTAIL.n301 VTAIL.n248 3.49141
R874 VTAIL.n278 VTAIL.n277 3.49141
R875 VTAIL.n210 VTAIL.n122 3.49141
R876 VTAIL.n189 VTAIL.n136 3.49141
R877 VTAIL.n166 VTAIL.n165 3.49141
R878 VTAIL.n382 VTAIL.n368 2.71565
R879 VTAIL.n410 VTAIL.n354 2.71565
R880 VTAIL.n431 VTAIL.n346 2.71565
R881 VTAIL.n46 VTAIL.n32 2.71565
R882 VTAIL.n74 VTAIL.n18 2.71565
R883 VTAIL.n95 VTAIL.n10 2.71565
R884 VTAIL.n321 VTAIL.n236 2.71565
R885 VTAIL.n302 VTAIL.n246 2.71565
R886 VTAIL.n274 VTAIL.n260 2.71565
R887 VTAIL.n209 VTAIL.n124 2.71565
R888 VTAIL.n190 VTAIL.n134 2.71565
R889 VTAIL.n162 VTAIL.n148 2.71565
R890 VTAIL.n381 VTAIL.n370 1.93989
R891 VTAIL.n415 VTAIL.n413 1.93989
R892 VTAIL.n428 VTAIL.n427 1.93989
R893 VTAIL.n45 VTAIL.n34 1.93989
R894 VTAIL.n79 VTAIL.n77 1.93989
R895 VTAIL.n92 VTAIL.n91 1.93989
R896 VTAIL.n318 VTAIL.n317 1.93989
R897 VTAIL.n306 VTAIL.n305 1.93989
R898 VTAIL.n273 VTAIL.n262 1.93989
R899 VTAIL.n206 VTAIL.n205 1.93989
R900 VTAIL.n194 VTAIL.n193 1.93989
R901 VTAIL.n161 VTAIL.n150 1.93989
R902 VTAIL.n0 VTAIL.t7 1.64966
R903 VTAIL.n0 VTAIL.t11 1.64966
R904 VTAIL.n112 VTAIL.t4 1.64966
R905 VTAIL.n112 VTAIL.t2 1.64966
R906 VTAIL.n226 VTAIL.t0 1.64966
R907 VTAIL.n226 VTAIL.t1 1.64966
R908 VTAIL.n114 VTAIL.t8 1.64966
R909 VTAIL.n114 VTAIL.t9 1.64966
R910 VTAIL.n225 VTAIL.n115 1.26774
R911 VTAIL.n337 VTAIL.n227 1.26774
R912 VTAIL.n113 VTAIL.n111 1.26774
R913 VTAIL.n378 VTAIL.n377 1.16414
R914 VTAIL.n414 VTAIL.n352 1.16414
R915 VTAIL.n424 VTAIL.n348 1.16414
R916 VTAIL.n42 VTAIL.n41 1.16414
R917 VTAIL.n78 VTAIL.n16 1.16414
R918 VTAIL.n88 VTAIL.n12 1.16414
R919 VTAIL.n314 VTAIL.n238 1.16414
R920 VTAIL.n309 VTAIL.n243 1.16414
R921 VTAIL.n270 VTAIL.n269 1.16414
R922 VTAIL.n202 VTAIL.n126 1.16414
R923 VTAIL.n197 VTAIL.n131 1.16414
R924 VTAIL.n158 VTAIL.n157 1.16414
R925 VTAIL.n227 VTAIL.n225 1.10395
R926 VTAIL.n111 VTAIL.n1 1.10395
R927 VTAIL VTAIL.n447 0.892741
R928 VTAIL.n374 VTAIL.n372 0.388379
R929 VTAIL.n420 VTAIL.n419 0.388379
R930 VTAIL.n423 VTAIL.n350 0.388379
R931 VTAIL.n38 VTAIL.n36 0.388379
R932 VTAIL.n84 VTAIL.n83 0.388379
R933 VTAIL.n87 VTAIL.n14 0.388379
R934 VTAIL.n313 VTAIL.n240 0.388379
R935 VTAIL.n310 VTAIL.n242 0.388379
R936 VTAIL.n266 VTAIL.n264 0.388379
R937 VTAIL.n201 VTAIL.n128 0.388379
R938 VTAIL.n198 VTAIL.n130 0.388379
R939 VTAIL.n154 VTAIL.n152 0.388379
R940 VTAIL VTAIL.n1 0.3755
R941 VTAIL.n379 VTAIL.n371 0.155672
R942 VTAIL.n380 VTAIL.n379 0.155672
R943 VTAIL.n380 VTAIL.n367 0.155672
R944 VTAIL.n387 VTAIL.n367 0.155672
R945 VTAIL.n388 VTAIL.n387 0.155672
R946 VTAIL.n388 VTAIL.n363 0.155672
R947 VTAIL.n395 VTAIL.n363 0.155672
R948 VTAIL.n396 VTAIL.n395 0.155672
R949 VTAIL.n396 VTAIL.n359 0.155672
R950 VTAIL.n403 VTAIL.n359 0.155672
R951 VTAIL.n404 VTAIL.n403 0.155672
R952 VTAIL.n404 VTAIL.n355 0.155672
R953 VTAIL.n411 VTAIL.n355 0.155672
R954 VTAIL.n412 VTAIL.n411 0.155672
R955 VTAIL.n412 VTAIL.n351 0.155672
R956 VTAIL.n421 VTAIL.n351 0.155672
R957 VTAIL.n422 VTAIL.n421 0.155672
R958 VTAIL.n422 VTAIL.n347 0.155672
R959 VTAIL.n429 VTAIL.n347 0.155672
R960 VTAIL.n430 VTAIL.n429 0.155672
R961 VTAIL.n430 VTAIL.n343 0.155672
R962 VTAIL.n437 VTAIL.n343 0.155672
R963 VTAIL.n438 VTAIL.n437 0.155672
R964 VTAIL.n438 VTAIL.n339 0.155672
R965 VTAIL.n445 VTAIL.n339 0.155672
R966 VTAIL.n43 VTAIL.n35 0.155672
R967 VTAIL.n44 VTAIL.n43 0.155672
R968 VTAIL.n44 VTAIL.n31 0.155672
R969 VTAIL.n51 VTAIL.n31 0.155672
R970 VTAIL.n52 VTAIL.n51 0.155672
R971 VTAIL.n52 VTAIL.n27 0.155672
R972 VTAIL.n59 VTAIL.n27 0.155672
R973 VTAIL.n60 VTAIL.n59 0.155672
R974 VTAIL.n60 VTAIL.n23 0.155672
R975 VTAIL.n67 VTAIL.n23 0.155672
R976 VTAIL.n68 VTAIL.n67 0.155672
R977 VTAIL.n68 VTAIL.n19 0.155672
R978 VTAIL.n75 VTAIL.n19 0.155672
R979 VTAIL.n76 VTAIL.n75 0.155672
R980 VTAIL.n76 VTAIL.n15 0.155672
R981 VTAIL.n85 VTAIL.n15 0.155672
R982 VTAIL.n86 VTAIL.n85 0.155672
R983 VTAIL.n86 VTAIL.n11 0.155672
R984 VTAIL.n93 VTAIL.n11 0.155672
R985 VTAIL.n94 VTAIL.n93 0.155672
R986 VTAIL.n94 VTAIL.n7 0.155672
R987 VTAIL.n101 VTAIL.n7 0.155672
R988 VTAIL.n102 VTAIL.n101 0.155672
R989 VTAIL.n102 VTAIL.n3 0.155672
R990 VTAIL.n109 VTAIL.n3 0.155672
R991 VTAIL.n335 VTAIL.n229 0.155672
R992 VTAIL.n328 VTAIL.n229 0.155672
R993 VTAIL.n328 VTAIL.n327 0.155672
R994 VTAIL.n327 VTAIL.n233 0.155672
R995 VTAIL.n320 VTAIL.n233 0.155672
R996 VTAIL.n320 VTAIL.n319 0.155672
R997 VTAIL.n319 VTAIL.n237 0.155672
R998 VTAIL.n312 VTAIL.n237 0.155672
R999 VTAIL.n312 VTAIL.n311 0.155672
R1000 VTAIL.n311 VTAIL.n241 0.155672
R1001 VTAIL.n304 VTAIL.n241 0.155672
R1002 VTAIL.n304 VTAIL.n303 0.155672
R1003 VTAIL.n303 VTAIL.n247 0.155672
R1004 VTAIL.n296 VTAIL.n247 0.155672
R1005 VTAIL.n296 VTAIL.n295 0.155672
R1006 VTAIL.n295 VTAIL.n251 0.155672
R1007 VTAIL.n288 VTAIL.n251 0.155672
R1008 VTAIL.n288 VTAIL.n287 0.155672
R1009 VTAIL.n287 VTAIL.n255 0.155672
R1010 VTAIL.n280 VTAIL.n255 0.155672
R1011 VTAIL.n280 VTAIL.n279 0.155672
R1012 VTAIL.n279 VTAIL.n259 0.155672
R1013 VTAIL.n272 VTAIL.n259 0.155672
R1014 VTAIL.n272 VTAIL.n271 0.155672
R1015 VTAIL.n271 VTAIL.n263 0.155672
R1016 VTAIL.n223 VTAIL.n117 0.155672
R1017 VTAIL.n216 VTAIL.n117 0.155672
R1018 VTAIL.n216 VTAIL.n215 0.155672
R1019 VTAIL.n215 VTAIL.n121 0.155672
R1020 VTAIL.n208 VTAIL.n121 0.155672
R1021 VTAIL.n208 VTAIL.n207 0.155672
R1022 VTAIL.n207 VTAIL.n125 0.155672
R1023 VTAIL.n200 VTAIL.n125 0.155672
R1024 VTAIL.n200 VTAIL.n199 0.155672
R1025 VTAIL.n199 VTAIL.n129 0.155672
R1026 VTAIL.n192 VTAIL.n129 0.155672
R1027 VTAIL.n192 VTAIL.n191 0.155672
R1028 VTAIL.n191 VTAIL.n135 0.155672
R1029 VTAIL.n184 VTAIL.n135 0.155672
R1030 VTAIL.n184 VTAIL.n183 0.155672
R1031 VTAIL.n183 VTAIL.n139 0.155672
R1032 VTAIL.n176 VTAIL.n139 0.155672
R1033 VTAIL.n176 VTAIL.n175 0.155672
R1034 VTAIL.n175 VTAIL.n143 0.155672
R1035 VTAIL.n168 VTAIL.n143 0.155672
R1036 VTAIL.n168 VTAIL.n167 0.155672
R1037 VTAIL.n167 VTAIL.n147 0.155672
R1038 VTAIL.n160 VTAIL.n147 0.155672
R1039 VTAIL.n160 VTAIL.n159 0.155672
R1040 VTAIL.n159 VTAIL.n151 0.155672
R1041 VP.n3 VP.t2 474.664
R1042 VP.n8 VP.t3 451.346
R1043 VP.n14 VP.t1 451.346
R1044 VP.n6 VP.t5 451.346
R1045 VP.n12 VP.t0 416.676
R1046 VP.n4 VP.t4 416.676
R1047 VP.n5 VP.n2 161.3
R1048 VP.n13 VP.n0 161.3
R1049 VP.n12 VP.n11 161.3
R1050 VP.n10 VP.n1 161.3
R1051 VP.n7 VP.n6 80.6037
R1052 VP.n15 VP.n14 80.6037
R1053 VP.n9 VP.n8 80.6037
R1054 VP.n8 VP.n1 51.6259
R1055 VP.n14 VP.n13 51.6259
R1056 VP.n6 VP.n5 51.6259
R1057 VP.n9 VP.n7 49.0203
R1058 VP.n4 VP.n3 32.927
R1059 VP.n3 VP.n2 27.9957
R1060 VP.n12 VP.n1 24.4675
R1061 VP.n13 VP.n12 24.4675
R1062 VP.n5 VP.n4 24.4675
R1063 VP.n7 VP.n2 0.285035
R1064 VP.n10 VP.n9 0.285035
R1065 VP.n15 VP.n0 0.285035
R1066 VP.n11 VP.n10 0.189894
R1067 VP.n11 VP.n0 0.189894
R1068 VP VP.n15 0.146778
R1069 VDD1.n104 VDD1.n0 756.745
R1070 VDD1.n213 VDD1.n109 756.745
R1071 VDD1.n105 VDD1.n104 585
R1072 VDD1.n103 VDD1.n102 585
R1073 VDD1.n4 VDD1.n3 585
R1074 VDD1.n97 VDD1.n96 585
R1075 VDD1.n95 VDD1.n94 585
R1076 VDD1.n8 VDD1.n7 585
R1077 VDD1.n89 VDD1.n88 585
R1078 VDD1.n87 VDD1.n86 585
R1079 VDD1.n12 VDD1.n11 585
R1080 VDD1.n16 VDD1.n14 585
R1081 VDD1.n81 VDD1.n80 585
R1082 VDD1.n79 VDD1.n78 585
R1083 VDD1.n18 VDD1.n17 585
R1084 VDD1.n73 VDD1.n72 585
R1085 VDD1.n71 VDD1.n70 585
R1086 VDD1.n22 VDD1.n21 585
R1087 VDD1.n65 VDD1.n64 585
R1088 VDD1.n63 VDD1.n62 585
R1089 VDD1.n26 VDD1.n25 585
R1090 VDD1.n57 VDD1.n56 585
R1091 VDD1.n55 VDD1.n54 585
R1092 VDD1.n30 VDD1.n29 585
R1093 VDD1.n49 VDD1.n48 585
R1094 VDD1.n47 VDD1.n46 585
R1095 VDD1.n34 VDD1.n33 585
R1096 VDD1.n41 VDD1.n40 585
R1097 VDD1.n39 VDD1.n38 585
R1098 VDD1.n146 VDD1.n145 585
R1099 VDD1.n148 VDD1.n147 585
R1100 VDD1.n141 VDD1.n140 585
R1101 VDD1.n154 VDD1.n153 585
R1102 VDD1.n156 VDD1.n155 585
R1103 VDD1.n137 VDD1.n136 585
R1104 VDD1.n162 VDD1.n161 585
R1105 VDD1.n164 VDD1.n163 585
R1106 VDD1.n133 VDD1.n132 585
R1107 VDD1.n170 VDD1.n169 585
R1108 VDD1.n172 VDD1.n171 585
R1109 VDD1.n129 VDD1.n128 585
R1110 VDD1.n178 VDD1.n177 585
R1111 VDD1.n180 VDD1.n179 585
R1112 VDD1.n125 VDD1.n124 585
R1113 VDD1.n187 VDD1.n186 585
R1114 VDD1.n188 VDD1.n123 585
R1115 VDD1.n190 VDD1.n189 585
R1116 VDD1.n121 VDD1.n120 585
R1117 VDD1.n196 VDD1.n195 585
R1118 VDD1.n198 VDD1.n197 585
R1119 VDD1.n117 VDD1.n116 585
R1120 VDD1.n204 VDD1.n203 585
R1121 VDD1.n206 VDD1.n205 585
R1122 VDD1.n113 VDD1.n112 585
R1123 VDD1.n212 VDD1.n211 585
R1124 VDD1.n214 VDD1.n213 585
R1125 VDD1.n37 VDD1.t3 327.466
R1126 VDD1.n144 VDD1.t2 327.466
R1127 VDD1.n104 VDD1.n103 171.744
R1128 VDD1.n103 VDD1.n3 171.744
R1129 VDD1.n96 VDD1.n3 171.744
R1130 VDD1.n96 VDD1.n95 171.744
R1131 VDD1.n95 VDD1.n7 171.744
R1132 VDD1.n88 VDD1.n7 171.744
R1133 VDD1.n88 VDD1.n87 171.744
R1134 VDD1.n87 VDD1.n11 171.744
R1135 VDD1.n16 VDD1.n11 171.744
R1136 VDD1.n80 VDD1.n16 171.744
R1137 VDD1.n80 VDD1.n79 171.744
R1138 VDD1.n79 VDD1.n17 171.744
R1139 VDD1.n72 VDD1.n17 171.744
R1140 VDD1.n72 VDD1.n71 171.744
R1141 VDD1.n71 VDD1.n21 171.744
R1142 VDD1.n64 VDD1.n21 171.744
R1143 VDD1.n64 VDD1.n63 171.744
R1144 VDD1.n63 VDD1.n25 171.744
R1145 VDD1.n56 VDD1.n25 171.744
R1146 VDD1.n56 VDD1.n55 171.744
R1147 VDD1.n55 VDD1.n29 171.744
R1148 VDD1.n48 VDD1.n29 171.744
R1149 VDD1.n48 VDD1.n47 171.744
R1150 VDD1.n47 VDD1.n33 171.744
R1151 VDD1.n40 VDD1.n33 171.744
R1152 VDD1.n40 VDD1.n39 171.744
R1153 VDD1.n147 VDD1.n146 171.744
R1154 VDD1.n147 VDD1.n140 171.744
R1155 VDD1.n154 VDD1.n140 171.744
R1156 VDD1.n155 VDD1.n154 171.744
R1157 VDD1.n155 VDD1.n136 171.744
R1158 VDD1.n162 VDD1.n136 171.744
R1159 VDD1.n163 VDD1.n162 171.744
R1160 VDD1.n163 VDD1.n132 171.744
R1161 VDD1.n170 VDD1.n132 171.744
R1162 VDD1.n171 VDD1.n170 171.744
R1163 VDD1.n171 VDD1.n128 171.744
R1164 VDD1.n178 VDD1.n128 171.744
R1165 VDD1.n179 VDD1.n178 171.744
R1166 VDD1.n179 VDD1.n124 171.744
R1167 VDD1.n187 VDD1.n124 171.744
R1168 VDD1.n188 VDD1.n187 171.744
R1169 VDD1.n189 VDD1.n188 171.744
R1170 VDD1.n189 VDD1.n120 171.744
R1171 VDD1.n196 VDD1.n120 171.744
R1172 VDD1.n197 VDD1.n196 171.744
R1173 VDD1.n197 VDD1.n116 171.744
R1174 VDD1.n204 VDD1.n116 171.744
R1175 VDD1.n205 VDD1.n204 171.744
R1176 VDD1.n205 VDD1.n112 171.744
R1177 VDD1.n212 VDD1.n112 171.744
R1178 VDD1.n213 VDD1.n212 171.744
R1179 VDD1.n39 VDD1.t3 85.8723
R1180 VDD1.n146 VDD1.t2 85.8723
R1181 VDD1.n219 VDD1.n218 68.9529
R1182 VDD1.n221 VDD1.n220 68.6914
R1183 VDD1 VDD1.n108 50.4546
R1184 VDD1.n219 VDD1.n217 50.341
R1185 VDD1.n221 VDD1.n219 46.0418
R1186 VDD1.n38 VDD1.n37 16.3895
R1187 VDD1.n145 VDD1.n144 16.3895
R1188 VDD1.n14 VDD1.n12 13.1884
R1189 VDD1.n190 VDD1.n121 13.1884
R1190 VDD1.n86 VDD1.n85 12.8005
R1191 VDD1.n82 VDD1.n81 12.8005
R1192 VDD1.n41 VDD1.n36 12.8005
R1193 VDD1.n148 VDD1.n143 12.8005
R1194 VDD1.n191 VDD1.n123 12.8005
R1195 VDD1.n195 VDD1.n194 12.8005
R1196 VDD1.n89 VDD1.n10 12.0247
R1197 VDD1.n78 VDD1.n15 12.0247
R1198 VDD1.n42 VDD1.n34 12.0247
R1199 VDD1.n149 VDD1.n141 12.0247
R1200 VDD1.n186 VDD1.n185 12.0247
R1201 VDD1.n198 VDD1.n119 12.0247
R1202 VDD1.n90 VDD1.n8 11.249
R1203 VDD1.n77 VDD1.n18 11.249
R1204 VDD1.n46 VDD1.n45 11.249
R1205 VDD1.n153 VDD1.n152 11.249
R1206 VDD1.n184 VDD1.n125 11.249
R1207 VDD1.n199 VDD1.n117 11.249
R1208 VDD1.n94 VDD1.n93 10.4732
R1209 VDD1.n74 VDD1.n73 10.4732
R1210 VDD1.n49 VDD1.n32 10.4732
R1211 VDD1.n156 VDD1.n139 10.4732
R1212 VDD1.n181 VDD1.n180 10.4732
R1213 VDD1.n203 VDD1.n202 10.4732
R1214 VDD1.n97 VDD1.n6 9.69747
R1215 VDD1.n70 VDD1.n20 9.69747
R1216 VDD1.n50 VDD1.n30 9.69747
R1217 VDD1.n157 VDD1.n137 9.69747
R1218 VDD1.n177 VDD1.n127 9.69747
R1219 VDD1.n206 VDD1.n115 9.69747
R1220 VDD1.n108 VDD1.n107 9.45567
R1221 VDD1.n217 VDD1.n216 9.45567
R1222 VDD1.n24 VDD1.n23 9.3005
R1223 VDD1.n67 VDD1.n66 9.3005
R1224 VDD1.n69 VDD1.n68 9.3005
R1225 VDD1.n20 VDD1.n19 9.3005
R1226 VDD1.n75 VDD1.n74 9.3005
R1227 VDD1.n77 VDD1.n76 9.3005
R1228 VDD1.n15 VDD1.n13 9.3005
R1229 VDD1.n83 VDD1.n82 9.3005
R1230 VDD1.n107 VDD1.n106 9.3005
R1231 VDD1.n2 VDD1.n1 9.3005
R1232 VDD1.n101 VDD1.n100 9.3005
R1233 VDD1.n99 VDD1.n98 9.3005
R1234 VDD1.n6 VDD1.n5 9.3005
R1235 VDD1.n93 VDD1.n92 9.3005
R1236 VDD1.n91 VDD1.n90 9.3005
R1237 VDD1.n10 VDD1.n9 9.3005
R1238 VDD1.n85 VDD1.n84 9.3005
R1239 VDD1.n61 VDD1.n60 9.3005
R1240 VDD1.n59 VDD1.n58 9.3005
R1241 VDD1.n28 VDD1.n27 9.3005
R1242 VDD1.n53 VDD1.n52 9.3005
R1243 VDD1.n51 VDD1.n50 9.3005
R1244 VDD1.n32 VDD1.n31 9.3005
R1245 VDD1.n45 VDD1.n44 9.3005
R1246 VDD1.n43 VDD1.n42 9.3005
R1247 VDD1.n36 VDD1.n35 9.3005
R1248 VDD1.n216 VDD1.n215 9.3005
R1249 VDD1.n210 VDD1.n209 9.3005
R1250 VDD1.n208 VDD1.n207 9.3005
R1251 VDD1.n115 VDD1.n114 9.3005
R1252 VDD1.n202 VDD1.n201 9.3005
R1253 VDD1.n200 VDD1.n199 9.3005
R1254 VDD1.n119 VDD1.n118 9.3005
R1255 VDD1.n194 VDD1.n193 9.3005
R1256 VDD1.n166 VDD1.n165 9.3005
R1257 VDD1.n135 VDD1.n134 9.3005
R1258 VDD1.n160 VDD1.n159 9.3005
R1259 VDD1.n158 VDD1.n157 9.3005
R1260 VDD1.n139 VDD1.n138 9.3005
R1261 VDD1.n152 VDD1.n151 9.3005
R1262 VDD1.n150 VDD1.n149 9.3005
R1263 VDD1.n143 VDD1.n142 9.3005
R1264 VDD1.n168 VDD1.n167 9.3005
R1265 VDD1.n131 VDD1.n130 9.3005
R1266 VDD1.n174 VDD1.n173 9.3005
R1267 VDD1.n176 VDD1.n175 9.3005
R1268 VDD1.n127 VDD1.n126 9.3005
R1269 VDD1.n182 VDD1.n181 9.3005
R1270 VDD1.n184 VDD1.n183 9.3005
R1271 VDD1.n185 VDD1.n122 9.3005
R1272 VDD1.n192 VDD1.n191 9.3005
R1273 VDD1.n111 VDD1.n110 9.3005
R1274 VDD1.n98 VDD1.n4 8.92171
R1275 VDD1.n69 VDD1.n22 8.92171
R1276 VDD1.n54 VDD1.n53 8.92171
R1277 VDD1.n161 VDD1.n160 8.92171
R1278 VDD1.n176 VDD1.n129 8.92171
R1279 VDD1.n207 VDD1.n113 8.92171
R1280 VDD1.n102 VDD1.n101 8.14595
R1281 VDD1.n66 VDD1.n65 8.14595
R1282 VDD1.n57 VDD1.n28 8.14595
R1283 VDD1.n164 VDD1.n135 8.14595
R1284 VDD1.n173 VDD1.n172 8.14595
R1285 VDD1.n211 VDD1.n210 8.14595
R1286 VDD1.n108 VDD1.n0 7.3702
R1287 VDD1.n105 VDD1.n2 7.3702
R1288 VDD1.n62 VDD1.n24 7.3702
R1289 VDD1.n58 VDD1.n26 7.3702
R1290 VDD1.n165 VDD1.n133 7.3702
R1291 VDD1.n169 VDD1.n131 7.3702
R1292 VDD1.n214 VDD1.n111 7.3702
R1293 VDD1.n217 VDD1.n109 7.3702
R1294 VDD1.n106 VDD1.n0 6.59444
R1295 VDD1.n106 VDD1.n105 6.59444
R1296 VDD1.n62 VDD1.n61 6.59444
R1297 VDD1.n61 VDD1.n26 6.59444
R1298 VDD1.n168 VDD1.n133 6.59444
R1299 VDD1.n169 VDD1.n168 6.59444
R1300 VDD1.n215 VDD1.n214 6.59444
R1301 VDD1.n215 VDD1.n109 6.59444
R1302 VDD1.n102 VDD1.n2 5.81868
R1303 VDD1.n65 VDD1.n24 5.81868
R1304 VDD1.n58 VDD1.n57 5.81868
R1305 VDD1.n165 VDD1.n164 5.81868
R1306 VDD1.n172 VDD1.n131 5.81868
R1307 VDD1.n211 VDD1.n111 5.81868
R1308 VDD1.n101 VDD1.n4 5.04292
R1309 VDD1.n66 VDD1.n22 5.04292
R1310 VDD1.n54 VDD1.n28 5.04292
R1311 VDD1.n161 VDD1.n135 5.04292
R1312 VDD1.n173 VDD1.n129 5.04292
R1313 VDD1.n210 VDD1.n113 5.04292
R1314 VDD1.n98 VDD1.n97 4.26717
R1315 VDD1.n70 VDD1.n69 4.26717
R1316 VDD1.n53 VDD1.n30 4.26717
R1317 VDD1.n160 VDD1.n137 4.26717
R1318 VDD1.n177 VDD1.n176 4.26717
R1319 VDD1.n207 VDD1.n206 4.26717
R1320 VDD1.n37 VDD1.n35 3.70982
R1321 VDD1.n144 VDD1.n142 3.70982
R1322 VDD1.n94 VDD1.n6 3.49141
R1323 VDD1.n73 VDD1.n20 3.49141
R1324 VDD1.n50 VDD1.n49 3.49141
R1325 VDD1.n157 VDD1.n156 3.49141
R1326 VDD1.n180 VDD1.n127 3.49141
R1327 VDD1.n203 VDD1.n115 3.49141
R1328 VDD1.n93 VDD1.n8 2.71565
R1329 VDD1.n74 VDD1.n18 2.71565
R1330 VDD1.n46 VDD1.n32 2.71565
R1331 VDD1.n153 VDD1.n139 2.71565
R1332 VDD1.n181 VDD1.n125 2.71565
R1333 VDD1.n202 VDD1.n117 2.71565
R1334 VDD1.n90 VDD1.n89 1.93989
R1335 VDD1.n78 VDD1.n77 1.93989
R1336 VDD1.n45 VDD1.n34 1.93989
R1337 VDD1.n152 VDD1.n141 1.93989
R1338 VDD1.n186 VDD1.n184 1.93989
R1339 VDD1.n199 VDD1.n198 1.93989
R1340 VDD1.n220 VDD1.t1 1.64966
R1341 VDD1.n220 VDD1.t0 1.64966
R1342 VDD1.n218 VDD1.t5 1.64966
R1343 VDD1.n218 VDD1.t4 1.64966
R1344 VDD1.n86 VDD1.n10 1.16414
R1345 VDD1.n81 VDD1.n15 1.16414
R1346 VDD1.n42 VDD1.n41 1.16414
R1347 VDD1.n149 VDD1.n148 1.16414
R1348 VDD1.n185 VDD1.n123 1.16414
R1349 VDD1.n195 VDD1.n119 1.16414
R1350 VDD1.n85 VDD1.n12 0.388379
R1351 VDD1.n82 VDD1.n14 0.388379
R1352 VDD1.n38 VDD1.n36 0.388379
R1353 VDD1.n145 VDD1.n143 0.388379
R1354 VDD1.n191 VDD1.n190 0.388379
R1355 VDD1.n194 VDD1.n121 0.388379
R1356 VDD1 VDD1.n221 0.259121
R1357 VDD1.n107 VDD1.n1 0.155672
R1358 VDD1.n100 VDD1.n1 0.155672
R1359 VDD1.n100 VDD1.n99 0.155672
R1360 VDD1.n99 VDD1.n5 0.155672
R1361 VDD1.n92 VDD1.n5 0.155672
R1362 VDD1.n92 VDD1.n91 0.155672
R1363 VDD1.n91 VDD1.n9 0.155672
R1364 VDD1.n84 VDD1.n9 0.155672
R1365 VDD1.n84 VDD1.n83 0.155672
R1366 VDD1.n83 VDD1.n13 0.155672
R1367 VDD1.n76 VDD1.n13 0.155672
R1368 VDD1.n76 VDD1.n75 0.155672
R1369 VDD1.n75 VDD1.n19 0.155672
R1370 VDD1.n68 VDD1.n19 0.155672
R1371 VDD1.n68 VDD1.n67 0.155672
R1372 VDD1.n67 VDD1.n23 0.155672
R1373 VDD1.n60 VDD1.n23 0.155672
R1374 VDD1.n60 VDD1.n59 0.155672
R1375 VDD1.n59 VDD1.n27 0.155672
R1376 VDD1.n52 VDD1.n27 0.155672
R1377 VDD1.n52 VDD1.n51 0.155672
R1378 VDD1.n51 VDD1.n31 0.155672
R1379 VDD1.n44 VDD1.n31 0.155672
R1380 VDD1.n44 VDD1.n43 0.155672
R1381 VDD1.n43 VDD1.n35 0.155672
R1382 VDD1.n150 VDD1.n142 0.155672
R1383 VDD1.n151 VDD1.n150 0.155672
R1384 VDD1.n151 VDD1.n138 0.155672
R1385 VDD1.n158 VDD1.n138 0.155672
R1386 VDD1.n159 VDD1.n158 0.155672
R1387 VDD1.n159 VDD1.n134 0.155672
R1388 VDD1.n166 VDD1.n134 0.155672
R1389 VDD1.n167 VDD1.n166 0.155672
R1390 VDD1.n167 VDD1.n130 0.155672
R1391 VDD1.n174 VDD1.n130 0.155672
R1392 VDD1.n175 VDD1.n174 0.155672
R1393 VDD1.n175 VDD1.n126 0.155672
R1394 VDD1.n182 VDD1.n126 0.155672
R1395 VDD1.n183 VDD1.n182 0.155672
R1396 VDD1.n183 VDD1.n122 0.155672
R1397 VDD1.n192 VDD1.n122 0.155672
R1398 VDD1.n193 VDD1.n192 0.155672
R1399 VDD1.n193 VDD1.n118 0.155672
R1400 VDD1.n200 VDD1.n118 0.155672
R1401 VDD1.n201 VDD1.n200 0.155672
R1402 VDD1.n201 VDD1.n114 0.155672
R1403 VDD1.n208 VDD1.n114 0.155672
R1404 VDD1.n209 VDD1.n208 0.155672
R1405 VDD1.n209 VDD1.n110 0.155672
R1406 VDD1.n216 VDD1.n110 0.155672
R1407 B.n328 B.t3 620.467
R1408 B.n147 B.t0 620.467
R1409 B.n55 B.t9 620.467
R1410 B.n48 B.t6 620.467
R1411 B.n444 B.n443 585
R1412 B.n442 B.n115 585
R1413 B.n441 B.n440 585
R1414 B.n439 B.n116 585
R1415 B.n438 B.n437 585
R1416 B.n436 B.n117 585
R1417 B.n435 B.n434 585
R1418 B.n433 B.n118 585
R1419 B.n432 B.n431 585
R1420 B.n430 B.n119 585
R1421 B.n429 B.n428 585
R1422 B.n427 B.n120 585
R1423 B.n426 B.n425 585
R1424 B.n424 B.n121 585
R1425 B.n423 B.n422 585
R1426 B.n421 B.n122 585
R1427 B.n420 B.n419 585
R1428 B.n418 B.n123 585
R1429 B.n417 B.n416 585
R1430 B.n415 B.n124 585
R1431 B.n414 B.n413 585
R1432 B.n412 B.n125 585
R1433 B.n411 B.n410 585
R1434 B.n409 B.n126 585
R1435 B.n408 B.n407 585
R1436 B.n406 B.n127 585
R1437 B.n405 B.n404 585
R1438 B.n403 B.n128 585
R1439 B.n402 B.n401 585
R1440 B.n400 B.n129 585
R1441 B.n399 B.n398 585
R1442 B.n397 B.n130 585
R1443 B.n396 B.n395 585
R1444 B.n394 B.n131 585
R1445 B.n393 B.n392 585
R1446 B.n391 B.n132 585
R1447 B.n390 B.n389 585
R1448 B.n388 B.n133 585
R1449 B.n387 B.n386 585
R1450 B.n385 B.n134 585
R1451 B.n384 B.n383 585
R1452 B.n382 B.n135 585
R1453 B.n381 B.n380 585
R1454 B.n379 B.n136 585
R1455 B.n378 B.n377 585
R1456 B.n376 B.n137 585
R1457 B.n375 B.n374 585
R1458 B.n373 B.n138 585
R1459 B.n372 B.n371 585
R1460 B.n370 B.n139 585
R1461 B.n369 B.n368 585
R1462 B.n367 B.n140 585
R1463 B.n366 B.n365 585
R1464 B.n364 B.n141 585
R1465 B.n363 B.n362 585
R1466 B.n361 B.n142 585
R1467 B.n360 B.n359 585
R1468 B.n358 B.n143 585
R1469 B.n357 B.n356 585
R1470 B.n355 B.n144 585
R1471 B.n354 B.n353 585
R1472 B.n352 B.n145 585
R1473 B.n351 B.n350 585
R1474 B.n349 B.n146 585
R1475 B.n347 B.n346 585
R1476 B.n345 B.n149 585
R1477 B.n344 B.n343 585
R1478 B.n342 B.n150 585
R1479 B.n341 B.n340 585
R1480 B.n339 B.n151 585
R1481 B.n338 B.n337 585
R1482 B.n336 B.n152 585
R1483 B.n335 B.n334 585
R1484 B.n333 B.n153 585
R1485 B.n332 B.n331 585
R1486 B.n327 B.n154 585
R1487 B.n326 B.n325 585
R1488 B.n324 B.n155 585
R1489 B.n323 B.n322 585
R1490 B.n321 B.n156 585
R1491 B.n320 B.n319 585
R1492 B.n318 B.n157 585
R1493 B.n317 B.n316 585
R1494 B.n315 B.n158 585
R1495 B.n314 B.n313 585
R1496 B.n312 B.n159 585
R1497 B.n311 B.n310 585
R1498 B.n309 B.n160 585
R1499 B.n308 B.n307 585
R1500 B.n306 B.n161 585
R1501 B.n305 B.n304 585
R1502 B.n303 B.n162 585
R1503 B.n302 B.n301 585
R1504 B.n300 B.n163 585
R1505 B.n299 B.n298 585
R1506 B.n297 B.n164 585
R1507 B.n296 B.n295 585
R1508 B.n294 B.n165 585
R1509 B.n293 B.n292 585
R1510 B.n291 B.n166 585
R1511 B.n290 B.n289 585
R1512 B.n288 B.n167 585
R1513 B.n287 B.n286 585
R1514 B.n285 B.n168 585
R1515 B.n284 B.n283 585
R1516 B.n282 B.n169 585
R1517 B.n281 B.n280 585
R1518 B.n279 B.n170 585
R1519 B.n278 B.n277 585
R1520 B.n276 B.n171 585
R1521 B.n275 B.n274 585
R1522 B.n273 B.n172 585
R1523 B.n272 B.n271 585
R1524 B.n270 B.n173 585
R1525 B.n269 B.n268 585
R1526 B.n267 B.n174 585
R1527 B.n266 B.n265 585
R1528 B.n264 B.n175 585
R1529 B.n263 B.n262 585
R1530 B.n261 B.n176 585
R1531 B.n260 B.n259 585
R1532 B.n258 B.n177 585
R1533 B.n257 B.n256 585
R1534 B.n255 B.n178 585
R1535 B.n254 B.n253 585
R1536 B.n252 B.n179 585
R1537 B.n251 B.n250 585
R1538 B.n249 B.n180 585
R1539 B.n248 B.n247 585
R1540 B.n246 B.n181 585
R1541 B.n245 B.n244 585
R1542 B.n243 B.n182 585
R1543 B.n242 B.n241 585
R1544 B.n240 B.n183 585
R1545 B.n239 B.n238 585
R1546 B.n237 B.n184 585
R1547 B.n236 B.n235 585
R1548 B.n234 B.n185 585
R1549 B.n445 B.n114 585
R1550 B.n447 B.n446 585
R1551 B.n448 B.n113 585
R1552 B.n450 B.n449 585
R1553 B.n451 B.n112 585
R1554 B.n453 B.n452 585
R1555 B.n454 B.n111 585
R1556 B.n456 B.n455 585
R1557 B.n457 B.n110 585
R1558 B.n459 B.n458 585
R1559 B.n460 B.n109 585
R1560 B.n462 B.n461 585
R1561 B.n463 B.n108 585
R1562 B.n465 B.n464 585
R1563 B.n466 B.n107 585
R1564 B.n468 B.n467 585
R1565 B.n469 B.n106 585
R1566 B.n471 B.n470 585
R1567 B.n472 B.n105 585
R1568 B.n474 B.n473 585
R1569 B.n475 B.n104 585
R1570 B.n477 B.n476 585
R1571 B.n478 B.n103 585
R1572 B.n480 B.n479 585
R1573 B.n481 B.n102 585
R1574 B.n483 B.n482 585
R1575 B.n484 B.n101 585
R1576 B.n486 B.n485 585
R1577 B.n487 B.n100 585
R1578 B.n489 B.n488 585
R1579 B.n490 B.n99 585
R1580 B.n492 B.n491 585
R1581 B.n493 B.n98 585
R1582 B.n495 B.n494 585
R1583 B.n496 B.n97 585
R1584 B.n498 B.n497 585
R1585 B.n499 B.n96 585
R1586 B.n501 B.n500 585
R1587 B.n502 B.n95 585
R1588 B.n504 B.n503 585
R1589 B.n505 B.n94 585
R1590 B.n507 B.n506 585
R1591 B.n508 B.n93 585
R1592 B.n510 B.n509 585
R1593 B.n511 B.n92 585
R1594 B.n513 B.n512 585
R1595 B.n514 B.n91 585
R1596 B.n516 B.n515 585
R1597 B.n517 B.n90 585
R1598 B.n519 B.n518 585
R1599 B.n520 B.n89 585
R1600 B.n522 B.n521 585
R1601 B.n730 B.n729 585
R1602 B.n728 B.n15 585
R1603 B.n727 B.n726 585
R1604 B.n725 B.n16 585
R1605 B.n724 B.n723 585
R1606 B.n722 B.n17 585
R1607 B.n721 B.n720 585
R1608 B.n719 B.n18 585
R1609 B.n718 B.n717 585
R1610 B.n716 B.n19 585
R1611 B.n715 B.n714 585
R1612 B.n713 B.n20 585
R1613 B.n712 B.n711 585
R1614 B.n710 B.n21 585
R1615 B.n709 B.n708 585
R1616 B.n707 B.n22 585
R1617 B.n706 B.n705 585
R1618 B.n704 B.n23 585
R1619 B.n703 B.n702 585
R1620 B.n701 B.n24 585
R1621 B.n700 B.n699 585
R1622 B.n698 B.n25 585
R1623 B.n697 B.n696 585
R1624 B.n695 B.n26 585
R1625 B.n694 B.n693 585
R1626 B.n692 B.n27 585
R1627 B.n691 B.n690 585
R1628 B.n689 B.n28 585
R1629 B.n688 B.n687 585
R1630 B.n686 B.n29 585
R1631 B.n685 B.n684 585
R1632 B.n683 B.n30 585
R1633 B.n682 B.n681 585
R1634 B.n680 B.n31 585
R1635 B.n679 B.n678 585
R1636 B.n677 B.n32 585
R1637 B.n676 B.n675 585
R1638 B.n674 B.n33 585
R1639 B.n673 B.n672 585
R1640 B.n671 B.n34 585
R1641 B.n670 B.n669 585
R1642 B.n668 B.n35 585
R1643 B.n667 B.n666 585
R1644 B.n665 B.n36 585
R1645 B.n664 B.n663 585
R1646 B.n662 B.n37 585
R1647 B.n661 B.n660 585
R1648 B.n659 B.n38 585
R1649 B.n658 B.n657 585
R1650 B.n656 B.n39 585
R1651 B.n655 B.n654 585
R1652 B.n653 B.n40 585
R1653 B.n652 B.n651 585
R1654 B.n650 B.n41 585
R1655 B.n649 B.n648 585
R1656 B.n647 B.n42 585
R1657 B.n646 B.n645 585
R1658 B.n644 B.n43 585
R1659 B.n643 B.n642 585
R1660 B.n641 B.n44 585
R1661 B.n640 B.n639 585
R1662 B.n638 B.n45 585
R1663 B.n637 B.n636 585
R1664 B.n635 B.n46 585
R1665 B.n634 B.n633 585
R1666 B.n632 B.n47 585
R1667 B.n631 B.n630 585
R1668 B.n629 B.n51 585
R1669 B.n628 B.n627 585
R1670 B.n626 B.n52 585
R1671 B.n625 B.n624 585
R1672 B.n623 B.n53 585
R1673 B.n622 B.n621 585
R1674 B.n620 B.n54 585
R1675 B.n618 B.n617 585
R1676 B.n616 B.n57 585
R1677 B.n615 B.n614 585
R1678 B.n613 B.n58 585
R1679 B.n612 B.n611 585
R1680 B.n610 B.n59 585
R1681 B.n609 B.n608 585
R1682 B.n607 B.n60 585
R1683 B.n606 B.n605 585
R1684 B.n604 B.n61 585
R1685 B.n603 B.n602 585
R1686 B.n601 B.n62 585
R1687 B.n600 B.n599 585
R1688 B.n598 B.n63 585
R1689 B.n597 B.n596 585
R1690 B.n595 B.n64 585
R1691 B.n594 B.n593 585
R1692 B.n592 B.n65 585
R1693 B.n591 B.n590 585
R1694 B.n589 B.n66 585
R1695 B.n588 B.n587 585
R1696 B.n586 B.n67 585
R1697 B.n585 B.n584 585
R1698 B.n583 B.n68 585
R1699 B.n582 B.n581 585
R1700 B.n580 B.n69 585
R1701 B.n579 B.n578 585
R1702 B.n577 B.n70 585
R1703 B.n576 B.n575 585
R1704 B.n574 B.n71 585
R1705 B.n573 B.n572 585
R1706 B.n571 B.n72 585
R1707 B.n570 B.n569 585
R1708 B.n568 B.n73 585
R1709 B.n567 B.n566 585
R1710 B.n565 B.n74 585
R1711 B.n564 B.n563 585
R1712 B.n562 B.n75 585
R1713 B.n561 B.n560 585
R1714 B.n559 B.n76 585
R1715 B.n558 B.n557 585
R1716 B.n556 B.n77 585
R1717 B.n555 B.n554 585
R1718 B.n553 B.n78 585
R1719 B.n552 B.n551 585
R1720 B.n550 B.n79 585
R1721 B.n549 B.n548 585
R1722 B.n547 B.n80 585
R1723 B.n546 B.n545 585
R1724 B.n544 B.n81 585
R1725 B.n543 B.n542 585
R1726 B.n541 B.n82 585
R1727 B.n540 B.n539 585
R1728 B.n538 B.n83 585
R1729 B.n537 B.n536 585
R1730 B.n535 B.n84 585
R1731 B.n534 B.n533 585
R1732 B.n532 B.n85 585
R1733 B.n531 B.n530 585
R1734 B.n529 B.n86 585
R1735 B.n528 B.n527 585
R1736 B.n526 B.n87 585
R1737 B.n525 B.n524 585
R1738 B.n523 B.n88 585
R1739 B.n731 B.n14 585
R1740 B.n733 B.n732 585
R1741 B.n734 B.n13 585
R1742 B.n736 B.n735 585
R1743 B.n737 B.n12 585
R1744 B.n739 B.n738 585
R1745 B.n740 B.n11 585
R1746 B.n742 B.n741 585
R1747 B.n743 B.n10 585
R1748 B.n745 B.n744 585
R1749 B.n746 B.n9 585
R1750 B.n748 B.n747 585
R1751 B.n749 B.n8 585
R1752 B.n751 B.n750 585
R1753 B.n752 B.n7 585
R1754 B.n754 B.n753 585
R1755 B.n755 B.n6 585
R1756 B.n757 B.n756 585
R1757 B.n758 B.n5 585
R1758 B.n760 B.n759 585
R1759 B.n761 B.n4 585
R1760 B.n763 B.n762 585
R1761 B.n764 B.n3 585
R1762 B.n766 B.n765 585
R1763 B.n767 B.n0 585
R1764 B.n2 B.n1 585
R1765 B.n198 B.n197 585
R1766 B.n200 B.n199 585
R1767 B.n201 B.n196 585
R1768 B.n203 B.n202 585
R1769 B.n204 B.n195 585
R1770 B.n206 B.n205 585
R1771 B.n207 B.n194 585
R1772 B.n209 B.n208 585
R1773 B.n210 B.n193 585
R1774 B.n212 B.n211 585
R1775 B.n213 B.n192 585
R1776 B.n215 B.n214 585
R1777 B.n216 B.n191 585
R1778 B.n218 B.n217 585
R1779 B.n219 B.n190 585
R1780 B.n221 B.n220 585
R1781 B.n222 B.n189 585
R1782 B.n224 B.n223 585
R1783 B.n225 B.n188 585
R1784 B.n227 B.n226 585
R1785 B.n228 B.n187 585
R1786 B.n230 B.n229 585
R1787 B.n231 B.n186 585
R1788 B.n233 B.n232 585
R1789 B.n147 B.t1 543.227
R1790 B.n55 B.t11 543.227
R1791 B.n328 B.t4 543.227
R1792 B.n48 B.t8 543.227
R1793 B.n148 B.t2 514.718
R1794 B.n56 B.t10 514.718
R1795 B.n329 B.t5 514.718
R1796 B.n49 B.t7 514.718
R1797 B.n234 B.n233 497.305
R1798 B.n443 B.n114 497.305
R1799 B.n521 B.n88 497.305
R1800 B.n731 B.n730 497.305
R1801 B.n769 B.n768 256.663
R1802 B.n768 B.n767 235.042
R1803 B.n768 B.n2 235.042
R1804 B.n235 B.n234 163.367
R1805 B.n235 B.n184 163.367
R1806 B.n239 B.n184 163.367
R1807 B.n240 B.n239 163.367
R1808 B.n241 B.n240 163.367
R1809 B.n241 B.n182 163.367
R1810 B.n245 B.n182 163.367
R1811 B.n246 B.n245 163.367
R1812 B.n247 B.n246 163.367
R1813 B.n247 B.n180 163.367
R1814 B.n251 B.n180 163.367
R1815 B.n252 B.n251 163.367
R1816 B.n253 B.n252 163.367
R1817 B.n253 B.n178 163.367
R1818 B.n257 B.n178 163.367
R1819 B.n258 B.n257 163.367
R1820 B.n259 B.n258 163.367
R1821 B.n259 B.n176 163.367
R1822 B.n263 B.n176 163.367
R1823 B.n264 B.n263 163.367
R1824 B.n265 B.n264 163.367
R1825 B.n265 B.n174 163.367
R1826 B.n269 B.n174 163.367
R1827 B.n270 B.n269 163.367
R1828 B.n271 B.n270 163.367
R1829 B.n271 B.n172 163.367
R1830 B.n275 B.n172 163.367
R1831 B.n276 B.n275 163.367
R1832 B.n277 B.n276 163.367
R1833 B.n277 B.n170 163.367
R1834 B.n281 B.n170 163.367
R1835 B.n282 B.n281 163.367
R1836 B.n283 B.n282 163.367
R1837 B.n283 B.n168 163.367
R1838 B.n287 B.n168 163.367
R1839 B.n288 B.n287 163.367
R1840 B.n289 B.n288 163.367
R1841 B.n289 B.n166 163.367
R1842 B.n293 B.n166 163.367
R1843 B.n294 B.n293 163.367
R1844 B.n295 B.n294 163.367
R1845 B.n295 B.n164 163.367
R1846 B.n299 B.n164 163.367
R1847 B.n300 B.n299 163.367
R1848 B.n301 B.n300 163.367
R1849 B.n301 B.n162 163.367
R1850 B.n305 B.n162 163.367
R1851 B.n306 B.n305 163.367
R1852 B.n307 B.n306 163.367
R1853 B.n307 B.n160 163.367
R1854 B.n311 B.n160 163.367
R1855 B.n312 B.n311 163.367
R1856 B.n313 B.n312 163.367
R1857 B.n313 B.n158 163.367
R1858 B.n317 B.n158 163.367
R1859 B.n318 B.n317 163.367
R1860 B.n319 B.n318 163.367
R1861 B.n319 B.n156 163.367
R1862 B.n323 B.n156 163.367
R1863 B.n324 B.n323 163.367
R1864 B.n325 B.n324 163.367
R1865 B.n325 B.n154 163.367
R1866 B.n332 B.n154 163.367
R1867 B.n333 B.n332 163.367
R1868 B.n334 B.n333 163.367
R1869 B.n334 B.n152 163.367
R1870 B.n338 B.n152 163.367
R1871 B.n339 B.n338 163.367
R1872 B.n340 B.n339 163.367
R1873 B.n340 B.n150 163.367
R1874 B.n344 B.n150 163.367
R1875 B.n345 B.n344 163.367
R1876 B.n346 B.n345 163.367
R1877 B.n346 B.n146 163.367
R1878 B.n351 B.n146 163.367
R1879 B.n352 B.n351 163.367
R1880 B.n353 B.n352 163.367
R1881 B.n353 B.n144 163.367
R1882 B.n357 B.n144 163.367
R1883 B.n358 B.n357 163.367
R1884 B.n359 B.n358 163.367
R1885 B.n359 B.n142 163.367
R1886 B.n363 B.n142 163.367
R1887 B.n364 B.n363 163.367
R1888 B.n365 B.n364 163.367
R1889 B.n365 B.n140 163.367
R1890 B.n369 B.n140 163.367
R1891 B.n370 B.n369 163.367
R1892 B.n371 B.n370 163.367
R1893 B.n371 B.n138 163.367
R1894 B.n375 B.n138 163.367
R1895 B.n376 B.n375 163.367
R1896 B.n377 B.n376 163.367
R1897 B.n377 B.n136 163.367
R1898 B.n381 B.n136 163.367
R1899 B.n382 B.n381 163.367
R1900 B.n383 B.n382 163.367
R1901 B.n383 B.n134 163.367
R1902 B.n387 B.n134 163.367
R1903 B.n388 B.n387 163.367
R1904 B.n389 B.n388 163.367
R1905 B.n389 B.n132 163.367
R1906 B.n393 B.n132 163.367
R1907 B.n394 B.n393 163.367
R1908 B.n395 B.n394 163.367
R1909 B.n395 B.n130 163.367
R1910 B.n399 B.n130 163.367
R1911 B.n400 B.n399 163.367
R1912 B.n401 B.n400 163.367
R1913 B.n401 B.n128 163.367
R1914 B.n405 B.n128 163.367
R1915 B.n406 B.n405 163.367
R1916 B.n407 B.n406 163.367
R1917 B.n407 B.n126 163.367
R1918 B.n411 B.n126 163.367
R1919 B.n412 B.n411 163.367
R1920 B.n413 B.n412 163.367
R1921 B.n413 B.n124 163.367
R1922 B.n417 B.n124 163.367
R1923 B.n418 B.n417 163.367
R1924 B.n419 B.n418 163.367
R1925 B.n419 B.n122 163.367
R1926 B.n423 B.n122 163.367
R1927 B.n424 B.n423 163.367
R1928 B.n425 B.n424 163.367
R1929 B.n425 B.n120 163.367
R1930 B.n429 B.n120 163.367
R1931 B.n430 B.n429 163.367
R1932 B.n431 B.n430 163.367
R1933 B.n431 B.n118 163.367
R1934 B.n435 B.n118 163.367
R1935 B.n436 B.n435 163.367
R1936 B.n437 B.n436 163.367
R1937 B.n437 B.n116 163.367
R1938 B.n441 B.n116 163.367
R1939 B.n442 B.n441 163.367
R1940 B.n443 B.n442 163.367
R1941 B.n521 B.n520 163.367
R1942 B.n520 B.n519 163.367
R1943 B.n519 B.n90 163.367
R1944 B.n515 B.n90 163.367
R1945 B.n515 B.n514 163.367
R1946 B.n514 B.n513 163.367
R1947 B.n513 B.n92 163.367
R1948 B.n509 B.n92 163.367
R1949 B.n509 B.n508 163.367
R1950 B.n508 B.n507 163.367
R1951 B.n507 B.n94 163.367
R1952 B.n503 B.n94 163.367
R1953 B.n503 B.n502 163.367
R1954 B.n502 B.n501 163.367
R1955 B.n501 B.n96 163.367
R1956 B.n497 B.n96 163.367
R1957 B.n497 B.n496 163.367
R1958 B.n496 B.n495 163.367
R1959 B.n495 B.n98 163.367
R1960 B.n491 B.n98 163.367
R1961 B.n491 B.n490 163.367
R1962 B.n490 B.n489 163.367
R1963 B.n489 B.n100 163.367
R1964 B.n485 B.n100 163.367
R1965 B.n485 B.n484 163.367
R1966 B.n484 B.n483 163.367
R1967 B.n483 B.n102 163.367
R1968 B.n479 B.n102 163.367
R1969 B.n479 B.n478 163.367
R1970 B.n478 B.n477 163.367
R1971 B.n477 B.n104 163.367
R1972 B.n473 B.n104 163.367
R1973 B.n473 B.n472 163.367
R1974 B.n472 B.n471 163.367
R1975 B.n471 B.n106 163.367
R1976 B.n467 B.n106 163.367
R1977 B.n467 B.n466 163.367
R1978 B.n466 B.n465 163.367
R1979 B.n465 B.n108 163.367
R1980 B.n461 B.n108 163.367
R1981 B.n461 B.n460 163.367
R1982 B.n460 B.n459 163.367
R1983 B.n459 B.n110 163.367
R1984 B.n455 B.n110 163.367
R1985 B.n455 B.n454 163.367
R1986 B.n454 B.n453 163.367
R1987 B.n453 B.n112 163.367
R1988 B.n449 B.n112 163.367
R1989 B.n449 B.n448 163.367
R1990 B.n448 B.n447 163.367
R1991 B.n447 B.n114 163.367
R1992 B.n730 B.n15 163.367
R1993 B.n726 B.n15 163.367
R1994 B.n726 B.n725 163.367
R1995 B.n725 B.n724 163.367
R1996 B.n724 B.n17 163.367
R1997 B.n720 B.n17 163.367
R1998 B.n720 B.n719 163.367
R1999 B.n719 B.n718 163.367
R2000 B.n718 B.n19 163.367
R2001 B.n714 B.n19 163.367
R2002 B.n714 B.n713 163.367
R2003 B.n713 B.n712 163.367
R2004 B.n712 B.n21 163.367
R2005 B.n708 B.n21 163.367
R2006 B.n708 B.n707 163.367
R2007 B.n707 B.n706 163.367
R2008 B.n706 B.n23 163.367
R2009 B.n702 B.n23 163.367
R2010 B.n702 B.n701 163.367
R2011 B.n701 B.n700 163.367
R2012 B.n700 B.n25 163.367
R2013 B.n696 B.n25 163.367
R2014 B.n696 B.n695 163.367
R2015 B.n695 B.n694 163.367
R2016 B.n694 B.n27 163.367
R2017 B.n690 B.n27 163.367
R2018 B.n690 B.n689 163.367
R2019 B.n689 B.n688 163.367
R2020 B.n688 B.n29 163.367
R2021 B.n684 B.n29 163.367
R2022 B.n684 B.n683 163.367
R2023 B.n683 B.n682 163.367
R2024 B.n682 B.n31 163.367
R2025 B.n678 B.n31 163.367
R2026 B.n678 B.n677 163.367
R2027 B.n677 B.n676 163.367
R2028 B.n676 B.n33 163.367
R2029 B.n672 B.n33 163.367
R2030 B.n672 B.n671 163.367
R2031 B.n671 B.n670 163.367
R2032 B.n670 B.n35 163.367
R2033 B.n666 B.n35 163.367
R2034 B.n666 B.n665 163.367
R2035 B.n665 B.n664 163.367
R2036 B.n664 B.n37 163.367
R2037 B.n660 B.n37 163.367
R2038 B.n660 B.n659 163.367
R2039 B.n659 B.n658 163.367
R2040 B.n658 B.n39 163.367
R2041 B.n654 B.n39 163.367
R2042 B.n654 B.n653 163.367
R2043 B.n653 B.n652 163.367
R2044 B.n652 B.n41 163.367
R2045 B.n648 B.n41 163.367
R2046 B.n648 B.n647 163.367
R2047 B.n647 B.n646 163.367
R2048 B.n646 B.n43 163.367
R2049 B.n642 B.n43 163.367
R2050 B.n642 B.n641 163.367
R2051 B.n641 B.n640 163.367
R2052 B.n640 B.n45 163.367
R2053 B.n636 B.n45 163.367
R2054 B.n636 B.n635 163.367
R2055 B.n635 B.n634 163.367
R2056 B.n634 B.n47 163.367
R2057 B.n630 B.n47 163.367
R2058 B.n630 B.n629 163.367
R2059 B.n629 B.n628 163.367
R2060 B.n628 B.n52 163.367
R2061 B.n624 B.n52 163.367
R2062 B.n624 B.n623 163.367
R2063 B.n623 B.n622 163.367
R2064 B.n622 B.n54 163.367
R2065 B.n617 B.n54 163.367
R2066 B.n617 B.n616 163.367
R2067 B.n616 B.n615 163.367
R2068 B.n615 B.n58 163.367
R2069 B.n611 B.n58 163.367
R2070 B.n611 B.n610 163.367
R2071 B.n610 B.n609 163.367
R2072 B.n609 B.n60 163.367
R2073 B.n605 B.n60 163.367
R2074 B.n605 B.n604 163.367
R2075 B.n604 B.n603 163.367
R2076 B.n603 B.n62 163.367
R2077 B.n599 B.n62 163.367
R2078 B.n599 B.n598 163.367
R2079 B.n598 B.n597 163.367
R2080 B.n597 B.n64 163.367
R2081 B.n593 B.n64 163.367
R2082 B.n593 B.n592 163.367
R2083 B.n592 B.n591 163.367
R2084 B.n591 B.n66 163.367
R2085 B.n587 B.n66 163.367
R2086 B.n587 B.n586 163.367
R2087 B.n586 B.n585 163.367
R2088 B.n585 B.n68 163.367
R2089 B.n581 B.n68 163.367
R2090 B.n581 B.n580 163.367
R2091 B.n580 B.n579 163.367
R2092 B.n579 B.n70 163.367
R2093 B.n575 B.n70 163.367
R2094 B.n575 B.n574 163.367
R2095 B.n574 B.n573 163.367
R2096 B.n573 B.n72 163.367
R2097 B.n569 B.n72 163.367
R2098 B.n569 B.n568 163.367
R2099 B.n568 B.n567 163.367
R2100 B.n567 B.n74 163.367
R2101 B.n563 B.n74 163.367
R2102 B.n563 B.n562 163.367
R2103 B.n562 B.n561 163.367
R2104 B.n561 B.n76 163.367
R2105 B.n557 B.n76 163.367
R2106 B.n557 B.n556 163.367
R2107 B.n556 B.n555 163.367
R2108 B.n555 B.n78 163.367
R2109 B.n551 B.n78 163.367
R2110 B.n551 B.n550 163.367
R2111 B.n550 B.n549 163.367
R2112 B.n549 B.n80 163.367
R2113 B.n545 B.n80 163.367
R2114 B.n545 B.n544 163.367
R2115 B.n544 B.n543 163.367
R2116 B.n543 B.n82 163.367
R2117 B.n539 B.n82 163.367
R2118 B.n539 B.n538 163.367
R2119 B.n538 B.n537 163.367
R2120 B.n537 B.n84 163.367
R2121 B.n533 B.n84 163.367
R2122 B.n533 B.n532 163.367
R2123 B.n532 B.n531 163.367
R2124 B.n531 B.n86 163.367
R2125 B.n527 B.n86 163.367
R2126 B.n527 B.n526 163.367
R2127 B.n526 B.n525 163.367
R2128 B.n525 B.n88 163.367
R2129 B.n732 B.n731 163.367
R2130 B.n732 B.n13 163.367
R2131 B.n736 B.n13 163.367
R2132 B.n737 B.n736 163.367
R2133 B.n738 B.n737 163.367
R2134 B.n738 B.n11 163.367
R2135 B.n742 B.n11 163.367
R2136 B.n743 B.n742 163.367
R2137 B.n744 B.n743 163.367
R2138 B.n744 B.n9 163.367
R2139 B.n748 B.n9 163.367
R2140 B.n749 B.n748 163.367
R2141 B.n750 B.n749 163.367
R2142 B.n750 B.n7 163.367
R2143 B.n754 B.n7 163.367
R2144 B.n755 B.n754 163.367
R2145 B.n756 B.n755 163.367
R2146 B.n756 B.n5 163.367
R2147 B.n760 B.n5 163.367
R2148 B.n761 B.n760 163.367
R2149 B.n762 B.n761 163.367
R2150 B.n762 B.n3 163.367
R2151 B.n766 B.n3 163.367
R2152 B.n767 B.n766 163.367
R2153 B.n198 B.n2 163.367
R2154 B.n199 B.n198 163.367
R2155 B.n199 B.n196 163.367
R2156 B.n203 B.n196 163.367
R2157 B.n204 B.n203 163.367
R2158 B.n205 B.n204 163.367
R2159 B.n205 B.n194 163.367
R2160 B.n209 B.n194 163.367
R2161 B.n210 B.n209 163.367
R2162 B.n211 B.n210 163.367
R2163 B.n211 B.n192 163.367
R2164 B.n215 B.n192 163.367
R2165 B.n216 B.n215 163.367
R2166 B.n217 B.n216 163.367
R2167 B.n217 B.n190 163.367
R2168 B.n221 B.n190 163.367
R2169 B.n222 B.n221 163.367
R2170 B.n223 B.n222 163.367
R2171 B.n223 B.n188 163.367
R2172 B.n227 B.n188 163.367
R2173 B.n228 B.n227 163.367
R2174 B.n229 B.n228 163.367
R2175 B.n229 B.n186 163.367
R2176 B.n233 B.n186 163.367
R2177 B.n330 B.n329 59.5399
R2178 B.n348 B.n148 59.5399
R2179 B.n619 B.n56 59.5399
R2180 B.n50 B.n49 59.5399
R2181 B.n729 B.n14 32.3127
R2182 B.n523 B.n522 32.3127
R2183 B.n445 B.n444 32.3127
R2184 B.n232 B.n185 32.3127
R2185 B.n329 B.n328 28.5096
R2186 B.n148 B.n147 28.5096
R2187 B.n56 B.n55 28.5096
R2188 B.n49 B.n48 28.5096
R2189 B B.n769 18.0485
R2190 B.n733 B.n14 10.6151
R2191 B.n734 B.n733 10.6151
R2192 B.n735 B.n734 10.6151
R2193 B.n735 B.n12 10.6151
R2194 B.n739 B.n12 10.6151
R2195 B.n740 B.n739 10.6151
R2196 B.n741 B.n740 10.6151
R2197 B.n741 B.n10 10.6151
R2198 B.n745 B.n10 10.6151
R2199 B.n746 B.n745 10.6151
R2200 B.n747 B.n746 10.6151
R2201 B.n747 B.n8 10.6151
R2202 B.n751 B.n8 10.6151
R2203 B.n752 B.n751 10.6151
R2204 B.n753 B.n752 10.6151
R2205 B.n753 B.n6 10.6151
R2206 B.n757 B.n6 10.6151
R2207 B.n758 B.n757 10.6151
R2208 B.n759 B.n758 10.6151
R2209 B.n759 B.n4 10.6151
R2210 B.n763 B.n4 10.6151
R2211 B.n764 B.n763 10.6151
R2212 B.n765 B.n764 10.6151
R2213 B.n765 B.n0 10.6151
R2214 B.n729 B.n728 10.6151
R2215 B.n728 B.n727 10.6151
R2216 B.n727 B.n16 10.6151
R2217 B.n723 B.n16 10.6151
R2218 B.n723 B.n722 10.6151
R2219 B.n722 B.n721 10.6151
R2220 B.n721 B.n18 10.6151
R2221 B.n717 B.n18 10.6151
R2222 B.n717 B.n716 10.6151
R2223 B.n716 B.n715 10.6151
R2224 B.n715 B.n20 10.6151
R2225 B.n711 B.n20 10.6151
R2226 B.n711 B.n710 10.6151
R2227 B.n710 B.n709 10.6151
R2228 B.n709 B.n22 10.6151
R2229 B.n705 B.n22 10.6151
R2230 B.n705 B.n704 10.6151
R2231 B.n704 B.n703 10.6151
R2232 B.n703 B.n24 10.6151
R2233 B.n699 B.n24 10.6151
R2234 B.n699 B.n698 10.6151
R2235 B.n698 B.n697 10.6151
R2236 B.n697 B.n26 10.6151
R2237 B.n693 B.n26 10.6151
R2238 B.n693 B.n692 10.6151
R2239 B.n692 B.n691 10.6151
R2240 B.n691 B.n28 10.6151
R2241 B.n687 B.n28 10.6151
R2242 B.n687 B.n686 10.6151
R2243 B.n686 B.n685 10.6151
R2244 B.n685 B.n30 10.6151
R2245 B.n681 B.n30 10.6151
R2246 B.n681 B.n680 10.6151
R2247 B.n680 B.n679 10.6151
R2248 B.n679 B.n32 10.6151
R2249 B.n675 B.n32 10.6151
R2250 B.n675 B.n674 10.6151
R2251 B.n674 B.n673 10.6151
R2252 B.n673 B.n34 10.6151
R2253 B.n669 B.n34 10.6151
R2254 B.n669 B.n668 10.6151
R2255 B.n668 B.n667 10.6151
R2256 B.n667 B.n36 10.6151
R2257 B.n663 B.n36 10.6151
R2258 B.n663 B.n662 10.6151
R2259 B.n662 B.n661 10.6151
R2260 B.n661 B.n38 10.6151
R2261 B.n657 B.n38 10.6151
R2262 B.n657 B.n656 10.6151
R2263 B.n656 B.n655 10.6151
R2264 B.n655 B.n40 10.6151
R2265 B.n651 B.n40 10.6151
R2266 B.n651 B.n650 10.6151
R2267 B.n650 B.n649 10.6151
R2268 B.n649 B.n42 10.6151
R2269 B.n645 B.n42 10.6151
R2270 B.n645 B.n644 10.6151
R2271 B.n644 B.n643 10.6151
R2272 B.n643 B.n44 10.6151
R2273 B.n639 B.n44 10.6151
R2274 B.n639 B.n638 10.6151
R2275 B.n638 B.n637 10.6151
R2276 B.n637 B.n46 10.6151
R2277 B.n633 B.n632 10.6151
R2278 B.n632 B.n631 10.6151
R2279 B.n631 B.n51 10.6151
R2280 B.n627 B.n51 10.6151
R2281 B.n627 B.n626 10.6151
R2282 B.n626 B.n625 10.6151
R2283 B.n625 B.n53 10.6151
R2284 B.n621 B.n53 10.6151
R2285 B.n621 B.n620 10.6151
R2286 B.n618 B.n57 10.6151
R2287 B.n614 B.n57 10.6151
R2288 B.n614 B.n613 10.6151
R2289 B.n613 B.n612 10.6151
R2290 B.n612 B.n59 10.6151
R2291 B.n608 B.n59 10.6151
R2292 B.n608 B.n607 10.6151
R2293 B.n607 B.n606 10.6151
R2294 B.n606 B.n61 10.6151
R2295 B.n602 B.n61 10.6151
R2296 B.n602 B.n601 10.6151
R2297 B.n601 B.n600 10.6151
R2298 B.n600 B.n63 10.6151
R2299 B.n596 B.n63 10.6151
R2300 B.n596 B.n595 10.6151
R2301 B.n595 B.n594 10.6151
R2302 B.n594 B.n65 10.6151
R2303 B.n590 B.n65 10.6151
R2304 B.n590 B.n589 10.6151
R2305 B.n589 B.n588 10.6151
R2306 B.n588 B.n67 10.6151
R2307 B.n584 B.n67 10.6151
R2308 B.n584 B.n583 10.6151
R2309 B.n583 B.n582 10.6151
R2310 B.n582 B.n69 10.6151
R2311 B.n578 B.n69 10.6151
R2312 B.n578 B.n577 10.6151
R2313 B.n577 B.n576 10.6151
R2314 B.n576 B.n71 10.6151
R2315 B.n572 B.n71 10.6151
R2316 B.n572 B.n571 10.6151
R2317 B.n571 B.n570 10.6151
R2318 B.n570 B.n73 10.6151
R2319 B.n566 B.n73 10.6151
R2320 B.n566 B.n565 10.6151
R2321 B.n565 B.n564 10.6151
R2322 B.n564 B.n75 10.6151
R2323 B.n560 B.n75 10.6151
R2324 B.n560 B.n559 10.6151
R2325 B.n559 B.n558 10.6151
R2326 B.n558 B.n77 10.6151
R2327 B.n554 B.n77 10.6151
R2328 B.n554 B.n553 10.6151
R2329 B.n553 B.n552 10.6151
R2330 B.n552 B.n79 10.6151
R2331 B.n548 B.n79 10.6151
R2332 B.n548 B.n547 10.6151
R2333 B.n547 B.n546 10.6151
R2334 B.n546 B.n81 10.6151
R2335 B.n542 B.n81 10.6151
R2336 B.n542 B.n541 10.6151
R2337 B.n541 B.n540 10.6151
R2338 B.n540 B.n83 10.6151
R2339 B.n536 B.n83 10.6151
R2340 B.n536 B.n535 10.6151
R2341 B.n535 B.n534 10.6151
R2342 B.n534 B.n85 10.6151
R2343 B.n530 B.n85 10.6151
R2344 B.n530 B.n529 10.6151
R2345 B.n529 B.n528 10.6151
R2346 B.n528 B.n87 10.6151
R2347 B.n524 B.n87 10.6151
R2348 B.n524 B.n523 10.6151
R2349 B.n522 B.n89 10.6151
R2350 B.n518 B.n89 10.6151
R2351 B.n518 B.n517 10.6151
R2352 B.n517 B.n516 10.6151
R2353 B.n516 B.n91 10.6151
R2354 B.n512 B.n91 10.6151
R2355 B.n512 B.n511 10.6151
R2356 B.n511 B.n510 10.6151
R2357 B.n510 B.n93 10.6151
R2358 B.n506 B.n93 10.6151
R2359 B.n506 B.n505 10.6151
R2360 B.n505 B.n504 10.6151
R2361 B.n504 B.n95 10.6151
R2362 B.n500 B.n95 10.6151
R2363 B.n500 B.n499 10.6151
R2364 B.n499 B.n498 10.6151
R2365 B.n498 B.n97 10.6151
R2366 B.n494 B.n97 10.6151
R2367 B.n494 B.n493 10.6151
R2368 B.n493 B.n492 10.6151
R2369 B.n492 B.n99 10.6151
R2370 B.n488 B.n99 10.6151
R2371 B.n488 B.n487 10.6151
R2372 B.n487 B.n486 10.6151
R2373 B.n486 B.n101 10.6151
R2374 B.n482 B.n101 10.6151
R2375 B.n482 B.n481 10.6151
R2376 B.n481 B.n480 10.6151
R2377 B.n480 B.n103 10.6151
R2378 B.n476 B.n103 10.6151
R2379 B.n476 B.n475 10.6151
R2380 B.n475 B.n474 10.6151
R2381 B.n474 B.n105 10.6151
R2382 B.n470 B.n105 10.6151
R2383 B.n470 B.n469 10.6151
R2384 B.n469 B.n468 10.6151
R2385 B.n468 B.n107 10.6151
R2386 B.n464 B.n107 10.6151
R2387 B.n464 B.n463 10.6151
R2388 B.n463 B.n462 10.6151
R2389 B.n462 B.n109 10.6151
R2390 B.n458 B.n109 10.6151
R2391 B.n458 B.n457 10.6151
R2392 B.n457 B.n456 10.6151
R2393 B.n456 B.n111 10.6151
R2394 B.n452 B.n111 10.6151
R2395 B.n452 B.n451 10.6151
R2396 B.n451 B.n450 10.6151
R2397 B.n450 B.n113 10.6151
R2398 B.n446 B.n113 10.6151
R2399 B.n446 B.n445 10.6151
R2400 B.n197 B.n1 10.6151
R2401 B.n200 B.n197 10.6151
R2402 B.n201 B.n200 10.6151
R2403 B.n202 B.n201 10.6151
R2404 B.n202 B.n195 10.6151
R2405 B.n206 B.n195 10.6151
R2406 B.n207 B.n206 10.6151
R2407 B.n208 B.n207 10.6151
R2408 B.n208 B.n193 10.6151
R2409 B.n212 B.n193 10.6151
R2410 B.n213 B.n212 10.6151
R2411 B.n214 B.n213 10.6151
R2412 B.n214 B.n191 10.6151
R2413 B.n218 B.n191 10.6151
R2414 B.n219 B.n218 10.6151
R2415 B.n220 B.n219 10.6151
R2416 B.n220 B.n189 10.6151
R2417 B.n224 B.n189 10.6151
R2418 B.n225 B.n224 10.6151
R2419 B.n226 B.n225 10.6151
R2420 B.n226 B.n187 10.6151
R2421 B.n230 B.n187 10.6151
R2422 B.n231 B.n230 10.6151
R2423 B.n232 B.n231 10.6151
R2424 B.n236 B.n185 10.6151
R2425 B.n237 B.n236 10.6151
R2426 B.n238 B.n237 10.6151
R2427 B.n238 B.n183 10.6151
R2428 B.n242 B.n183 10.6151
R2429 B.n243 B.n242 10.6151
R2430 B.n244 B.n243 10.6151
R2431 B.n244 B.n181 10.6151
R2432 B.n248 B.n181 10.6151
R2433 B.n249 B.n248 10.6151
R2434 B.n250 B.n249 10.6151
R2435 B.n250 B.n179 10.6151
R2436 B.n254 B.n179 10.6151
R2437 B.n255 B.n254 10.6151
R2438 B.n256 B.n255 10.6151
R2439 B.n256 B.n177 10.6151
R2440 B.n260 B.n177 10.6151
R2441 B.n261 B.n260 10.6151
R2442 B.n262 B.n261 10.6151
R2443 B.n262 B.n175 10.6151
R2444 B.n266 B.n175 10.6151
R2445 B.n267 B.n266 10.6151
R2446 B.n268 B.n267 10.6151
R2447 B.n268 B.n173 10.6151
R2448 B.n272 B.n173 10.6151
R2449 B.n273 B.n272 10.6151
R2450 B.n274 B.n273 10.6151
R2451 B.n274 B.n171 10.6151
R2452 B.n278 B.n171 10.6151
R2453 B.n279 B.n278 10.6151
R2454 B.n280 B.n279 10.6151
R2455 B.n280 B.n169 10.6151
R2456 B.n284 B.n169 10.6151
R2457 B.n285 B.n284 10.6151
R2458 B.n286 B.n285 10.6151
R2459 B.n286 B.n167 10.6151
R2460 B.n290 B.n167 10.6151
R2461 B.n291 B.n290 10.6151
R2462 B.n292 B.n291 10.6151
R2463 B.n292 B.n165 10.6151
R2464 B.n296 B.n165 10.6151
R2465 B.n297 B.n296 10.6151
R2466 B.n298 B.n297 10.6151
R2467 B.n298 B.n163 10.6151
R2468 B.n302 B.n163 10.6151
R2469 B.n303 B.n302 10.6151
R2470 B.n304 B.n303 10.6151
R2471 B.n304 B.n161 10.6151
R2472 B.n308 B.n161 10.6151
R2473 B.n309 B.n308 10.6151
R2474 B.n310 B.n309 10.6151
R2475 B.n310 B.n159 10.6151
R2476 B.n314 B.n159 10.6151
R2477 B.n315 B.n314 10.6151
R2478 B.n316 B.n315 10.6151
R2479 B.n316 B.n157 10.6151
R2480 B.n320 B.n157 10.6151
R2481 B.n321 B.n320 10.6151
R2482 B.n322 B.n321 10.6151
R2483 B.n322 B.n155 10.6151
R2484 B.n326 B.n155 10.6151
R2485 B.n327 B.n326 10.6151
R2486 B.n331 B.n327 10.6151
R2487 B.n335 B.n153 10.6151
R2488 B.n336 B.n335 10.6151
R2489 B.n337 B.n336 10.6151
R2490 B.n337 B.n151 10.6151
R2491 B.n341 B.n151 10.6151
R2492 B.n342 B.n341 10.6151
R2493 B.n343 B.n342 10.6151
R2494 B.n343 B.n149 10.6151
R2495 B.n347 B.n149 10.6151
R2496 B.n350 B.n349 10.6151
R2497 B.n350 B.n145 10.6151
R2498 B.n354 B.n145 10.6151
R2499 B.n355 B.n354 10.6151
R2500 B.n356 B.n355 10.6151
R2501 B.n356 B.n143 10.6151
R2502 B.n360 B.n143 10.6151
R2503 B.n361 B.n360 10.6151
R2504 B.n362 B.n361 10.6151
R2505 B.n362 B.n141 10.6151
R2506 B.n366 B.n141 10.6151
R2507 B.n367 B.n366 10.6151
R2508 B.n368 B.n367 10.6151
R2509 B.n368 B.n139 10.6151
R2510 B.n372 B.n139 10.6151
R2511 B.n373 B.n372 10.6151
R2512 B.n374 B.n373 10.6151
R2513 B.n374 B.n137 10.6151
R2514 B.n378 B.n137 10.6151
R2515 B.n379 B.n378 10.6151
R2516 B.n380 B.n379 10.6151
R2517 B.n380 B.n135 10.6151
R2518 B.n384 B.n135 10.6151
R2519 B.n385 B.n384 10.6151
R2520 B.n386 B.n385 10.6151
R2521 B.n386 B.n133 10.6151
R2522 B.n390 B.n133 10.6151
R2523 B.n391 B.n390 10.6151
R2524 B.n392 B.n391 10.6151
R2525 B.n392 B.n131 10.6151
R2526 B.n396 B.n131 10.6151
R2527 B.n397 B.n396 10.6151
R2528 B.n398 B.n397 10.6151
R2529 B.n398 B.n129 10.6151
R2530 B.n402 B.n129 10.6151
R2531 B.n403 B.n402 10.6151
R2532 B.n404 B.n403 10.6151
R2533 B.n404 B.n127 10.6151
R2534 B.n408 B.n127 10.6151
R2535 B.n409 B.n408 10.6151
R2536 B.n410 B.n409 10.6151
R2537 B.n410 B.n125 10.6151
R2538 B.n414 B.n125 10.6151
R2539 B.n415 B.n414 10.6151
R2540 B.n416 B.n415 10.6151
R2541 B.n416 B.n123 10.6151
R2542 B.n420 B.n123 10.6151
R2543 B.n421 B.n420 10.6151
R2544 B.n422 B.n421 10.6151
R2545 B.n422 B.n121 10.6151
R2546 B.n426 B.n121 10.6151
R2547 B.n427 B.n426 10.6151
R2548 B.n428 B.n427 10.6151
R2549 B.n428 B.n119 10.6151
R2550 B.n432 B.n119 10.6151
R2551 B.n433 B.n432 10.6151
R2552 B.n434 B.n433 10.6151
R2553 B.n434 B.n117 10.6151
R2554 B.n438 B.n117 10.6151
R2555 B.n439 B.n438 10.6151
R2556 B.n440 B.n439 10.6151
R2557 B.n440 B.n115 10.6151
R2558 B.n444 B.n115 10.6151
R2559 B.n50 B.n46 9.36635
R2560 B.n619 B.n618 9.36635
R2561 B.n331 B.n330 9.36635
R2562 B.n349 B.n348 9.36635
R2563 B.n769 B.n0 8.11757
R2564 B.n769 B.n1 8.11757
R2565 B.n633 B.n50 1.24928
R2566 B.n620 B.n619 1.24928
R2567 B.n330 B.n153 1.24928
R2568 B.n348 B.n347 1.24928
C0 VTAIL B 4.46861f
C1 VDD2 w_n2146_n4910# 2.52508f
C2 VTAIL VP 8.094879f
C3 VN B 0.948647f
C4 VN VP 6.93234f
C5 VDD1 B 2.2689f
C6 VN VTAIL 8.08015f
C7 VDD2 B 2.30822f
C8 VDD1 VP 8.75266f
C9 VTAIL VDD1 12.5195f
C10 VDD2 VP 0.33581f
C11 VTAIL VDD2 12.5546f
C12 VN VDD1 0.148805f
C13 w_n2146_n4910# B 9.82179f
C14 VN VDD2 8.57189f
C15 w_n2146_n4910# VP 4.11846f
C16 VDD1 VDD2 0.874416f
C17 VTAIL w_n2146_n4910# 4.07002f
C18 VN w_n2146_n4910# 3.84508f
C19 B VP 1.39773f
C20 VDD1 w_n2146_n4910# 2.48709f
C21 VDD2 VSUBS 1.785766f
C22 VDD1 VSUBS 1.554288f
C23 VTAIL VSUBS 1.149f
C24 VN VSUBS 5.19754f
C25 VP VSUBS 2.113932f
C26 B VSUBS 3.849201f
C27 w_n2146_n4910# VSUBS 0.128683p
C28 B.n0 VSUBS 0.007314f
C29 B.n1 VSUBS 0.007314f
C30 B.n2 VSUBS 0.010817f
C31 B.n3 VSUBS 0.008289f
C32 B.n4 VSUBS 0.008289f
C33 B.n5 VSUBS 0.008289f
C34 B.n6 VSUBS 0.008289f
C35 B.n7 VSUBS 0.008289f
C36 B.n8 VSUBS 0.008289f
C37 B.n9 VSUBS 0.008289f
C38 B.n10 VSUBS 0.008289f
C39 B.n11 VSUBS 0.008289f
C40 B.n12 VSUBS 0.008289f
C41 B.n13 VSUBS 0.008289f
C42 B.n14 VSUBS 0.018935f
C43 B.n15 VSUBS 0.008289f
C44 B.n16 VSUBS 0.008289f
C45 B.n17 VSUBS 0.008289f
C46 B.n18 VSUBS 0.008289f
C47 B.n19 VSUBS 0.008289f
C48 B.n20 VSUBS 0.008289f
C49 B.n21 VSUBS 0.008289f
C50 B.n22 VSUBS 0.008289f
C51 B.n23 VSUBS 0.008289f
C52 B.n24 VSUBS 0.008289f
C53 B.n25 VSUBS 0.008289f
C54 B.n26 VSUBS 0.008289f
C55 B.n27 VSUBS 0.008289f
C56 B.n28 VSUBS 0.008289f
C57 B.n29 VSUBS 0.008289f
C58 B.n30 VSUBS 0.008289f
C59 B.n31 VSUBS 0.008289f
C60 B.n32 VSUBS 0.008289f
C61 B.n33 VSUBS 0.008289f
C62 B.n34 VSUBS 0.008289f
C63 B.n35 VSUBS 0.008289f
C64 B.n36 VSUBS 0.008289f
C65 B.n37 VSUBS 0.008289f
C66 B.n38 VSUBS 0.008289f
C67 B.n39 VSUBS 0.008289f
C68 B.n40 VSUBS 0.008289f
C69 B.n41 VSUBS 0.008289f
C70 B.n42 VSUBS 0.008289f
C71 B.n43 VSUBS 0.008289f
C72 B.n44 VSUBS 0.008289f
C73 B.n45 VSUBS 0.008289f
C74 B.n46 VSUBS 0.007802f
C75 B.n47 VSUBS 0.008289f
C76 B.t7 VSUBS 0.465345f
C77 B.t8 VSUBS 0.486017f
C78 B.t6 VSUBS 1.10195f
C79 B.n48 VSUBS 0.628312f
C80 B.n49 VSUBS 0.405716f
C81 B.n50 VSUBS 0.019206f
C82 B.n51 VSUBS 0.008289f
C83 B.n52 VSUBS 0.008289f
C84 B.n53 VSUBS 0.008289f
C85 B.n54 VSUBS 0.008289f
C86 B.t10 VSUBS 0.465349f
C87 B.t11 VSUBS 0.486021f
C88 B.t9 VSUBS 1.10195f
C89 B.n55 VSUBS 0.628308f
C90 B.n56 VSUBS 0.405711f
C91 B.n57 VSUBS 0.008289f
C92 B.n58 VSUBS 0.008289f
C93 B.n59 VSUBS 0.008289f
C94 B.n60 VSUBS 0.008289f
C95 B.n61 VSUBS 0.008289f
C96 B.n62 VSUBS 0.008289f
C97 B.n63 VSUBS 0.008289f
C98 B.n64 VSUBS 0.008289f
C99 B.n65 VSUBS 0.008289f
C100 B.n66 VSUBS 0.008289f
C101 B.n67 VSUBS 0.008289f
C102 B.n68 VSUBS 0.008289f
C103 B.n69 VSUBS 0.008289f
C104 B.n70 VSUBS 0.008289f
C105 B.n71 VSUBS 0.008289f
C106 B.n72 VSUBS 0.008289f
C107 B.n73 VSUBS 0.008289f
C108 B.n74 VSUBS 0.008289f
C109 B.n75 VSUBS 0.008289f
C110 B.n76 VSUBS 0.008289f
C111 B.n77 VSUBS 0.008289f
C112 B.n78 VSUBS 0.008289f
C113 B.n79 VSUBS 0.008289f
C114 B.n80 VSUBS 0.008289f
C115 B.n81 VSUBS 0.008289f
C116 B.n82 VSUBS 0.008289f
C117 B.n83 VSUBS 0.008289f
C118 B.n84 VSUBS 0.008289f
C119 B.n85 VSUBS 0.008289f
C120 B.n86 VSUBS 0.008289f
C121 B.n87 VSUBS 0.008289f
C122 B.n88 VSUBS 0.019587f
C123 B.n89 VSUBS 0.008289f
C124 B.n90 VSUBS 0.008289f
C125 B.n91 VSUBS 0.008289f
C126 B.n92 VSUBS 0.008289f
C127 B.n93 VSUBS 0.008289f
C128 B.n94 VSUBS 0.008289f
C129 B.n95 VSUBS 0.008289f
C130 B.n96 VSUBS 0.008289f
C131 B.n97 VSUBS 0.008289f
C132 B.n98 VSUBS 0.008289f
C133 B.n99 VSUBS 0.008289f
C134 B.n100 VSUBS 0.008289f
C135 B.n101 VSUBS 0.008289f
C136 B.n102 VSUBS 0.008289f
C137 B.n103 VSUBS 0.008289f
C138 B.n104 VSUBS 0.008289f
C139 B.n105 VSUBS 0.008289f
C140 B.n106 VSUBS 0.008289f
C141 B.n107 VSUBS 0.008289f
C142 B.n108 VSUBS 0.008289f
C143 B.n109 VSUBS 0.008289f
C144 B.n110 VSUBS 0.008289f
C145 B.n111 VSUBS 0.008289f
C146 B.n112 VSUBS 0.008289f
C147 B.n113 VSUBS 0.008289f
C148 B.n114 VSUBS 0.018935f
C149 B.n115 VSUBS 0.008289f
C150 B.n116 VSUBS 0.008289f
C151 B.n117 VSUBS 0.008289f
C152 B.n118 VSUBS 0.008289f
C153 B.n119 VSUBS 0.008289f
C154 B.n120 VSUBS 0.008289f
C155 B.n121 VSUBS 0.008289f
C156 B.n122 VSUBS 0.008289f
C157 B.n123 VSUBS 0.008289f
C158 B.n124 VSUBS 0.008289f
C159 B.n125 VSUBS 0.008289f
C160 B.n126 VSUBS 0.008289f
C161 B.n127 VSUBS 0.008289f
C162 B.n128 VSUBS 0.008289f
C163 B.n129 VSUBS 0.008289f
C164 B.n130 VSUBS 0.008289f
C165 B.n131 VSUBS 0.008289f
C166 B.n132 VSUBS 0.008289f
C167 B.n133 VSUBS 0.008289f
C168 B.n134 VSUBS 0.008289f
C169 B.n135 VSUBS 0.008289f
C170 B.n136 VSUBS 0.008289f
C171 B.n137 VSUBS 0.008289f
C172 B.n138 VSUBS 0.008289f
C173 B.n139 VSUBS 0.008289f
C174 B.n140 VSUBS 0.008289f
C175 B.n141 VSUBS 0.008289f
C176 B.n142 VSUBS 0.008289f
C177 B.n143 VSUBS 0.008289f
C178 B.n144 VSUBS 0.008289f
C179 B.n145 VSUBS 0.008289f
C180 B.n146 VSUBS 0.008289f
C181 B.t2 VSUBS 0.465349f
C182 B.t1 VSUBS 0.486021f
C183 B.t0 VSUBS 1.10195f
C184 B.n147 VSUBS 0.628308f
C185 B.n148 VSUBS 0.405711f
C186 B.n149 VSUBS 0.008289f
C187 B.n150 VSUBS 0.008289f
C188 B.n151 VSUBS 0.008289f
C189 B.n152 VSUBS 0.008289f
C190 B.n153 VSUBS 0.004632f
C191 B.n154 VSUBS 0.008289f
C192 B.n155 VSUBS 0.008289f
C193 B.n156 VSUBS 0.008289f
C194 B.n157 VSUBS 0.008289f
C195 B.n158 VSUBS 0.008289f
C196 B.n159 VSUBS 0.008289f
C197 B.n160 VSUBS 0.008289f
C198 B.n161 VSUBS 0.008289f
C199 B.n162 VSUBS 0.008289f
C200 B.n163 VSUBS 0.008289f
C201 B.n164 VSUBS 0.008289f
C202 B.n165 VSUBS 0.008289f
C203 B.n166 VSUBS 0.008289f
C204 B.n167 VSUBS 0.008289f
C205 B.n168 VSUBS 0.008289f
C206 B.n169 VSUBS 0.008289f
C207 B.n170 VSUBS 0.008289f
C208 B.n171 VSUBS 0.008289f
C209 B.n172 VSUBS 0.008289f
C210 B.n173 VSUBS 0.008289f
C211 B.n174 VSUBS 0.008289f
C212 B.n175 VSUBS 0.008289f
C213 B.n176 VSUBS 0.008289f
C214 B.n177 VSUBS 0.008289f
C215 B.n178 VSUBS 0.008289f
C216 B.n179 VSUBS 0.008289f
C217 B.n180 VSUBS 0.008289f
C218 B.n181 VSUBS 0.008289f
C219 B.n182 VSUBS 0.008289f
C220 B.n183 VSUBS 0.008289f
C221 B.n184 VSUBS 0.008289f
C222 B.n185 VSUBS 0.019587f
C223 B.n186 VSUBS 0.008289f
C224 B.n187 VSUBS 0.008289f
C225 B.n188 VSUBS 0.008289f
C226 B.n189 VSUBS 0.008289f
C227 B.n190 VSUBS 0.008289f
C228 B.n191 VSUBS 0.008289f
C229 B.n192 VSUBS 0.008289f
C230 B.n193 VSUBS 0.008289f
C231 B.n194 VSUBS 0.008289f
C232 B.n195 VSUBS 0.008289f
C233 B.n196 VSUBS 0.008289f
C234 B.n197 VSUBS 0.008289f
C235 B.n198 VSUBS 0.008289f
C236 B.n199 VSUBS 0.008289f
C237 B.n200 VSUBS 0.008289f
C238 B.n201 VSUBS 0.008289f
C239 B.n202 VSUBS 0.008289f
C240 B.n203 VSUBS 0.008289f
C241 B.n204 VSUBS 0.008289f
C242 B.n205 VSUBS 0.008289f
C243 B.n206 VSUBS 0.008289f
C244 B.n207 VSUBS 0.008289f
C245 B.n208 VSUBS 0.008289f
C246 B.n209 VSUBS 0.008289f
C247 B.n210 VSUBS 0.008289f
C248 B.n211 VSUBS 0.008289f
C249 B.n212 VSUBS 0.008289f
C250 B.n213 VSUBS 0.008289f
C251 B.n214 VSUBS 0.008289f
C252 B.n215 VSUBS 0.008289f
C253 B.n216 VSUBS 0.008289f
C254 B.n217 VSUBS 0.008289f
C255 B.n218 VSUBS 0.008289f
C256 B.n219 VSUBS 0.008289f
C257 B.n220 VSUBS 0.008289f
C258 B.n221 VSUBS 0.008289f
C259 B.n222 VSUBS 0.008289f
C260 B.n223 VSUBS 0.008289f
C261 B.n224 VSUBS 0.008289f
C262 B.n225 VSUBS 0.008289f
C263 B.n226 VSUBS 0.008289f
C264 B.n227 VSUBS 0.008289f
C265 B.n228 VSUBS 0.008289f
C266 B.n229 VSUBS 0.008289f
C267 B.n230 VSUBS 0.008289f
C268 B.n231 VSUBS 0.008289f
C269 B.n232 VSUBS 0.018935f
C270 B.n233 VSUBS 0.018935f
C271 B.n234 VSUBS 0.019587f
C272 B.n235 VSUBS 0.008289f
C273 B.n236 VSUBS 0.008289f
C274 B.n237 VSUBS 0.008289f
C275 B.n238 VSUBS 0.008289f
C276 B.n239 VSUBS 0.008289f
C277 B.n240 VSUBS 0.008289f
C278 B.n241 VSUBS 0.008289f
C279 B.n242 VSUBS 0.008289f
C280 B.n243 VSUBS 0.008289f
C281 B.n244 VSUBS 0.008289f
C282 B.n245 VSUBS 0.008289f
C283 B.n246 VSUBS 0.008289f
C284 B.n247 VSUBS 0.008289f
C285 B.n248 VSUBS 0.008289f
C286 B.n249 VSUBS 0.008289f
C287 B.n250 VSUBS 0.008289f
C288 B.n251 VSUBS 0.008289f
C289 B.n252 VSUBS 0.008289f
C290 B.n253 VSUBS 0.008289f
C291 B.n254 VSUBS 0.008289f
C292 B.n255 VSUBS 0.008289f
C293 B.n256 VSUBS 0.008289f
C294 B.n257 VSUBS 0.008289f
C295 B.n258 VSUBS 0.008289f
C296 B.n259 VSUBS 0.008289f
C297 B.n260 VSUBS 0.008289f
C298 B.n261 VSUBS 0.008289f
C299 B.n262 VSUBS 0.008289f
C300 B.n263 VSUBS 0.008289f
C301 B.n264 VSUBS 0.008289f
C302 B.n265 VSUBS 0.008289f
C303 B.n266 VSUBS 0.008289f
C304 B.n267 VSUBS 0.008289f
C305 B.n268 VSUBS 0.008289f
C306 B.n269 VSUBS 0.008289f
C307 B.n270 VSUBS 0.008289f
C308 B.n271 VSUBS 0.008289f
C309 B.n272 VSUBS 0.008289f
C310 B.n273 VSUBS 0.008289f
C311 B.n274 VSUBS 0.008289f
C312 B.n275 VSUBS 0.008289f
C313 B.n276 VSUBS 0.008289f
C314 B.n277 VSUBS 0.008289f
C315 B.n278 VSUBS 0.008289f
C316 B.n279 VSUBS 0.008289f
C317 B.n280 VSUBS 0.008289f
C318 B.n281 VSUBS 0.008289f
C319 B.n282 VSUBS 0.008289f
C320 B.n283 VSUBS 0.008289f
C321 B.n284 VSUBS 0.008289f
C322 B.n285 VSUBS 0.008289f
C323 B.n286 VSUBS 0.008289f
C324 B.n287 VSUBS 0.008289f
C325 B.n288 VSUBS 0.008289f
C326 B.n289 VSUBS 0.008289f
C327 B.n290 VSUBS 0.008289f
C328 B.n291 VSUBS 0.008289f
C329 B.n292 VSUBS 0.008289f
C330 B.n293 VSUBS 0.008289f
C331 B.n294 VSUBS 0.008289f
C332 B.n295 VSUBS 0.008289f
C333 B.n296 VSUBS 0.008289f
C334 B.n297 VSUBS 0.008289f
C335 B.n298 VSUBS 0.008289f
C336 B.n299 VSUBS 0.008289f
C337 B.n300 VSUBS 0.008289f
C338 B.n301 VSUBS 0.008289f
C339 B.n302 VSUBS 0.008289f
C340 B.n303 VSUBS 0.008289f
C341 B.n304 VSUBS 0.008289f
C342 B.n305 VSUBS 0.008289f
C343 B.n306 VSUBS 0.008289f
C344 B.n307 VSUBS 0.008289f
C345 B.n308 VSUBS 0.008289f
C346 B.n309 VSUBS 0.008289f
C347 B.n310 VSUBS 0.008289f
C348 B.n311 VSUBS 0.008289f
C349 B.n312 VSUBS 0.008289f
C350 B.n313 VSUBS 0.008289f
C351 B.n314 VSUBS 0.008289f
C352 B.n315 VSUBS 0.008289f
C353 B.n316 VSUBS 0.008289f
C354 B.n317 VSUBS 0.008289f
C355 B.n318 VSUBS 0.008289f
C356 B.n319 VSUBS 0.008289f
C357 B.n320 VSUBS 0.008289f
C358 B.n321 VSUBS 0.008289f
C359 B.n322 VSUBS 0.008289f
C360 B.n323 VSUBS 0.008289f
C361 B.n324 VSUBS 0.008289f
C362 B.n325 VSUBS 0.008289f
C363 B.n326 VSUBS 0.008289f
C364 B.n327 VSUBS 0.008289f
C365 B.t5 VSUBS 0.465345f
C366 B.t4 VSUBS 0.486017f
C367 B.t3 VSUBS 1.10195f
C368 B.n328 VSUBS 0.628312f
C369 B.n329 VSUBS 0.405716f
C370 B.n330 VSUBS 0.019206f
C371 B.n331 VSUBS 0.007802f
C372 B.n332 VSUBS 0.008289f
C373 B.n333 VSUBS 0.008289f
C374 B.n334 VSUBS 0.008289f
C375 B.n335 VSUBS 0.008289f
C376 B.n336 VSUBS 0.008289f
C377 B.n337 VSUBS 0.008289f
C378 B.n338 VSUBS 0.008289f
C379 B.n339 VSUBS 0.008289f
C380 B.n340 VSUBS 0.008289f
C381 B.n341 VSUBS 0.008289f
C382 B.n342 VSUBS 0.008289f
C383 B.n343 VSUBS 0.008289f
C384 B.n344 VSUBS 0.008289f
C385 B.n345 VSUBS 0.008289f
C386 B.n346 VSUBS 0.008289f
C387 B.n347 VSUBS 0.004632f
C388 B.n348 VSUBS 0.019206f
C389 B.n349 VSUBS 0.007802f
C390 B.n350 VSUBS 0.008289f
C391 B.n351 VSUBS 0.008289f
C392 B.n352 VSUBS 0.008289f
C393 B.n353 VSUBS 0.008289f
C394 B.n354 VSUBS 0.008289f
C395 B.n355 VSUBS 0.008289f
C396 B.n356 VSUBS 0.008289f
C397 B.n357 VSUBS 0.008289f
C398 B.n358 VSUBS 0.008289f
C399 B.n359 VSUBS 0.008289f
C400 B.n360 VSUBS 0.008289f
C401 B.n361 VSUBS 0.008289f
C402 B.n362 VSUBS 0.008289f
C403 B.n363 VSUBS 0.008289f
C404 B.n364 VSUBS 0.008289f
C405 B.n365 VSUBS 0.008289f
C406 B.n366 VSUBS 0.008289f
C407 B.n367 VSUBS 0.008289f
C408 B.n368 VSUBS 0.008289f
C409 B.n369 VSUBS 0.008289f
C410 B.n370 VSUBS 0.008289f
C411 B.n371 VSUBS 0.008289f
C412 B.n372 VSUBS 0.008289f
C413 B.n373 VSUBS 0.008289f
C414 B.n374 VSUBS 0.008289f
C415 B.n375 VSUBS 0.008289f
C416 B.n376 VSUBS 0.008289f
C417 B.n377 VSUBS 0.008289f
C418 B.n378 VSUBS 0.008289f
C419 B.n379 VSUBS 0.008289f
C420 B.n380 VSUBS 0.008289f
C421 B.n381 VSUBS 0.008289f
C422 B.n382 VSUBS 0.008289f
C423 B.n383 VSUBS 0.008289f
C424 B.n384 VSUBS 0.008289f
C425 B.n385 VSUBS 0.008289f
C426 B.n386 VSUBS 0.008289f
C427 B.n387 VSUBS 0.008289f
C428 B.n388 VSUBS 0.008289f
C429 B.n389 VSUBS 0.008289f
C430 B.n390 VSUBS 0.008289f
C431 B.n391 VSUBS 0.008289f
C432 B.n392 VSUBS 0.008289f
C433 B.n393 VSUBS 0.008289f
C434 B.n394 VSUBS 0.008289f
C435 B.n395 VSUBS 0.008289f
C436 B.n396 VSUBS 0.008289f
C437 B.n397 VSUBS 0.008289f
C438 B.n398 VSUBS 0.008289f
C439 B.n399 VSUBS 0.008289f
C440 B.n400 VSUBS 0.008289f
C441 B.n401 VSUBS 0.008289f
C442 B.n402 VSUBS 0.008289f
C443 B.n403 VSUBS 0.008289f
C444 B.n404 VSUBS 0.008289f
C445 B.n405 VSUBS 0.008289f
C446 B.n406 VSUBS 0.008289f
C447 B.n407 VSUBS 0.008289f
C448 B.n408 VSUBS 0.008289f
C449 B.n409 VSUBS 0.008289f
C450 B.n410 VSUBS 0.008289f
C451 B.n411 VSUBS 0.008289f
C452 B.n412 VSUBS 0.008289f
C453 B.n413 VSUBS 0.008289f
C454 B.n414 VSUBS 0.008289f
C455 B.n415 VSUBS 0.008289f
C456 B.n416 VSUBS 0.008289f
C457 B.n417 VSUBS 0.008289f
C458 B.n418 VSUBS 0.008289f
C459 B.n419 VSUBS 0.008289f
C460 B.n420 VSUBS 0.008289f
C461 B.n421 VSUBS 0.008289f
C462 B.n422 VSUBS 0.008289f
C463 B.n423 VSUBS 0.008289f
C464 B.n424 VSUBS 0.008289f
C465 B.n425 VSUBS 0.008289f
C466 B.n426 VSUBS 0.008289f
C467 B.n427 VSUBS 0.008289f
C468 B.n428 VSUBS 0.008289f
C469 B.n429 VSUBS 0.008289f
C470 B.n430 VSUBS 0.008289f
C471 B.n431 VSUBS 0.008289f
C472 B.n432 VSUBS 0.008289f
C473 B.n433 VSUBS 0.008289f
C474 B.n434 VSUBS 0.008289f
C475 B.n435 VSUBS 0.008289f
C476 B.n436 VSUBS 0.008289f
C477 B.n437 VSUBS 0.008289f
C478 B.n438 VSUBS 0.008289f
C479 B.n439 VSUBS 0.008289f
C480 B.n440 VSUBS 0.008289f
C481 B.n441 VSUBS 0.008289f
C482 B.n442 VSUBS 0.008289f
C483 B.n443 VSUBS 0.019587f
C484 B.n444 VSUBS 0.018597f
C485 B.n445 VSUBS 0.019925f
C486 B.n446 VSUBS 0.008289f
C487 B.n447 VSUBS 0.008289f
C488 B.n448 VSUBS 0.008289f
C489 B.n449 VSUBS 0.008289f
C490 B.n450 VSUBS 0.008289f
C491 B.n451 VSUBS 0.008289f
C492 B.n452 VSUBS 0.008289f
C493 B.n453 VSUBS 0.008289f
C494 B.n454 VSUBS 0.008289f
C495 B.n455 VSUBS 0.008289f
C496 B.n456 VSUBS 0.008289f
C497 B.n457 VSUBS 0.008289f
C498 B.n458 VSUBS 0.008289f
C499 B.n459 VSUBS 0.008289f
C500 B.n460 VSUBS 0.008289f
C501 B.n461 VSUBS 0.008289f
C502 B.n462 VSUBS 0.008289f
C503 B.n463 VSUBS 0.008289f
C504 B.n464 VSUBS 0.008289f
C505 B.n465 VSUBS 0.008289f
C506 B.n466 VSUBS 0.008289f
C507 B.n467 VSUBS 0.008289f
C508 B.n468 VSUBS 0.008289f
C509 B.n469 VSUBS 0.008289f
C510 B.n470 VSUBS 0.008289f
C511 B.n471 VSUBS 0.008289f
C512 B.n472 VSUBS 0.008289f
C513 B.n473 VSUBS 0.008289f
C514 B.n474 VSUBS 0.008289f
C515 B.n475 VSUBS 0.008289f
C516 B.n476 VSUBS 0.008289f
C517 B.n477 VSUBS 0.008289f
C518 B.n478 VSUBS 0.008289f
C519 B.n479 VSUBS 0.008289f
C520 B.n480 VSUBS 0.008289f
C521 B.n481 VSUBS 0.008289f
C522 B.n482 VSUBS 0.008289f
C523 B.n483 VSUBS 0.008289f
C524 B.n484 VSUBS 0.008289f
C525 B.n485 VSUBS 0.008289f
C526 B.n486 VSUBS 0.008289f
C527 B.n487 VSUBS 0.008289f
C528 B.n488 VSUBS 0.008289f
C529 B.n489 VSUBS 0.008289f
C530 B.n490 VSUBS 0.008289f
C531 B.n491 VSUBS 0.008289f
C532 B.n492 VSUBS 0.008289f
C533 B.n493 VSUBS 0.008289f
C534 B.n494 VSUBS 0.008289f
C535 B.n495 VSUBS 0.008289f
C536 B.n496 VSUBS 0.008289f
C537 B.n497 VSUBS 0.008289f
C538 B.n498 VSUBS 0.008289f
C539 B.n499 VSUBS 0.008289f
C540 B.n500 VSUBS 0.008289f
C541 B.n501 VSUBS 0.008289f
C542 B.n502 VSUBS 0.008289f
C543 B.n503 VSUBS 0.008289f
C544 B.n504 VSUBS 0.008289f
C545 B.n505 VSUBS 0.008289f
C546 B.n506 VSUBS 0.008289f
C547 B.n507 VSUBS 0.008289f
C548 B.n508 VSUBS 0.008289f
C549 B.n509 VSUBS 0.008289f
C550 B.n510 VSUBS 0.008289f
C551 B.n511 VSUBS 0.008289f
C552 B.n512 VSUBS 0.008289f
C553 B.n513 VSUBS 0.008289f
C554 B.n514 VSUBS 0.008289f
C555 B.n515 VSUBS 0.008289f
C556 B.n516 VSUBS 0.008289f
C557 B.n517 VSUBS 0.008289f
C558 B.n518 VSUBS 0.008289f
C559 B.n519 VSUBS 0.008289f
C560 B.n520 VSUBS 0.008289f
C561 B.n521 VSUBS 0.018935f
C562 B.n522 VSUBS 0.018935f
C563 B.n523 VSUBS 0.019587f
C564 B.n524 VSUBS 0.008289f
C565 B.n525 VSUBS 0.008289f
C566 B.n526 VSUBS 0.008289f
C567 B.n527 VSUBS 0.008289f
C568 B.n528 VSUBS 0.008289f
C569 B.n529 VSUBS 0.008289f
C570 B.n530 VSUBS 0.008289f
C571 B.n531 VSUBS 0.008289f
C572 B.n532 VSUBS 0.008289f
C573 B.n533 VSUBS 0.008289f
C574 B.n534 VSUBS 0.008289f
C575 B.n535 VSUBS 0.008289f
C576 B.n536 VSUBS 0.008289f
C577 B.n537 VSUBS 0.008289f
C578 B.n538 VSUBS 0.008289f
C579 B.n539 VSUBS 0.008289f
C580 B.n540 VSUBS 0.008289f
C581 B.n541 VSUBS 0.008289f
C582 B.n542 VSUBS 0.008289f
C583 B.n543 VSUBS 0.008289f
C584 B.n544 VSUBS 0.008289f
C585 B.n545 VSUBS 0.008289f
C586 B.n546 VSUBS 0.008289f
C587 B.n547 VSUBS 0.008289f
C588 B.n548 VSUBS 0.008289f
C589 B.n549 VSUBS 0.008289f
C590 B.n550 VSUBS 0.008289f
C591 B.n551 VSUBS 0.008289f
C592 B.n552 VSUBS 0.008289f
C593 B.n553 VSUBS 0.008289f
C594 B.n554 VSUBS 0.008289f
C595 B.n555 VSUBS 0.008289f
C596 B.n556 VSUBS 0.008289f
C597 B.n557 VSUBS 0.008289f
C598 B.n558 VSUBS 0.008289f
C599 B.n559 VSUBS 0.008289f
C600 B.n560 VSUBS 0.008289f
C601 B.n561 VSUBS 0.008289f
C602 B.n562 VSUBS 0.008289f
C603 B.n563 VSUBS 0.008289f
C604 B.n564 VSUBS 0.008289f
C605 B.n565 VSUBS 0.008289f
C606 B.n566 VSUBS 0.008289f
C607 B.n567 VSUBS 0.008289f
C608 B.n568 VSUBS 0.008289f
C609 B.n569 VSUBS 0.008289f
C610 B.n570 VSUBS 0.008289f
C611 B.n571 VSUBS 0.008289f
C612 B.n572 VSUBS 0.008289f
C613 B.n573 VSUBS 0.008289f
C614 B.n574 VSUBS 0.008289f
C615 B.n575 VSUBS 0.008289f
C616 B.n576 VSUBS 0.008289f
C617 B.n577 VSUBS 0.008289f
C618 B.n578 VSUBS 0.008289f
C619 B.n579 VSUBS 0.008289f
C620 B.n580 VSUBS 0.008289f
C621 B.n581 VSUBS 0.008289f
C622 B.n582 VSUBS 0.008289f
C623 B.n583 VSUBS 0.008289f
C624 B.n584 VSUBS 0.008289f
C625 B.n585 VSUBS 0.008289f
C626 B.n586 VSUBS 0.008289f
C627 B.n587 VSUBS 0.008289f
C628 B.n588 VSUBS 0.008289f
C629 B.n589 VSUBS 0.008289f
C630 B.n590 VSUBS 0.008289f
C631 B.n591 VSUBS 0.008289f
C632 B.n592 VSUBS 0.008289f
C633 B.n593 VSUBS 0.008289f
C634 B.n594 VSUBS 0.008289f
C635 B.n595 VSUBS 0.008289f
C636 B.n596 VSUBS 0.008289f
C637 B.n597 VSUBS 0.008289f
C638 B.n598 VSUBS 0.008289f
C639 B.n599 VSUBS 0.008289f
C640 B.n600 VSUBS 0.008289f
C641 B.n601 VSUBS 0.008289f
C642 B.n602 VSUBS 0.008289f
C643 B.n603 VSUBS 0.008289f
C644 B.n604 VSUBS 0.008289f
C645 B.n605 VSUBS 0.008289f
C646 B.n606 VSUBS 0.008289f
C647 B.n607 VSUBS 0.008289f
C648 B.n608 VSUBS 0.008289f
C649 B.n609 VSUBS 0.008289f
C650 B.n610 VSUBS 0.008289f
C651 B.n611 VSUBS 0.008289f
C652 B.n612 VSUBS 0.008289f
C653 B.n613 VSUBS 0.008289f
C654 B.n614 VSUBS 0.008289f
C655 B.n615 VSUBS 0.008289f
C656 B.n616 VSUBS 0.008289f
C657 B.n617 VSUBS 0.008289f
C658 B.n618 VSUBS 0.007802f
C659 B.n619 VSUBS 0.019206f
C660 B.n620 VSUBS 0.004632f
C661 B.n621 VSUBS 0.008289f
C662 B.n622 VSUBS 0.008289f
C663 B.n623 VSUBS 0.008289f
C664 B.n624 VSUBS 0.008289f
C665 B.n625 VSUBS 0.008289f
C666 B.n626 VSUBS 0.008289f
C667 B.n627 VSUBS 0.008289f
C668 B.n628 VSUBS 0.008289f
C669 B.n629 VSUBS 0.008289f
C670 B.n630 VSUBS 0.008289f
C671 B.n631 VSUBS 0.008289f
C672 B.n632 VSUBS 0.008289f
C673 B.n633 VSUBS 0.004632f
C674 B.n634 VSUBS 0.008289f
C675 B.n635 VSUBS 0.008289f
C676 B.n636 VSUBS 0.008289f
C677 B.n637 VSUBS 0.008289f
C678 B.n638 VSUBS 0.008289f
C679 B.n639 VSUBS 0.008289f
C680 B.n640 VSUBS 0.008289f
C681 B.n641 VSUBS 0.008289f
C682 B.n642 VSUBS 0.008289f
C683 B.n643 VSUBS 0.008289f
C684 B.n644 VSUBS 0.008289f
C685 B.n645 VSUBS 0.008289f
C686 B.n646 VSUBS 0.008289f
C687 B.n647 VSUBS 0.008289f
C688 B.n648 VSUBS 0.008289f
C689 B.n649 VSUBS 0.008289f
C690 B.n650 VSUBS 0.008289f
C691 B.n651 VSUBS 0.008289f
C692 B.n652 VSUBS 0.008289f
C693 B.n653 VSUBS 0.008289f
C694 B.n654 VSUBS 0.008289f
C695 B.n655 VSUBS 0.008289f
C696 B.n656 VSUBS 0.008289f
C697 B.n657 VSUBS 0.008289f
C698 B.n658 VSUBS 0.008289f
C699 B.n659 VSUBS 0.008289f
C700 B.n660 VSUBS 0.008289f
C701 B.n661 VSUBS 0.008289f
C702 B.n662 VSUBS 0.008289f
C703 B.n663 VSUBS 0.008289f
C704 B.n664 VSUBS 0.008289f
C705 B.n665 VSUBS 0.008289f
C706 B.n666 VSUBS 0.008289f
C707 B.n667 VSUBS 0.008289f
C708 B.n668 VSUBS 0.008289f
C709 B.n669 VSUBS 0.008289f
C710 B.n670 VSUBS 0.008289f
C711 B.n671 VSUBS 0.008289f
C712 B.n672 VSUBS 0.008289f
C713 B.n673 VSUBS 0.008289f
C714 B.n674 VSUBS 0.008289f
C715 B.n675 VSUBS 0.008289f
C716 B.n676 VSUBS 0.008289f
C717 B.n677 VSUBS 0.008289f
C718 B.n678 VSUBS 0.008289f
C719 B.n679 VSUBS 0.008289f
C720 B.n680 VSUBS 0.008289f
C721 B.n681 VSUBS 0.008289f
C722 B.n682 VSUBS 0.008289f
C723 B.n683 VSUBS 0.008289f
C724 B.n684 VSUBS 0.008289f
C725 B.n685 VSUBS 0.008289f
C726 B.n686 VSUBS 0.008289f
C727 B.n687 VSUBS 0.008289f
C728 B.n688 VSUBS 0.008289f
C729 B.n689 VSUBS 0.008289f
C730 B.n690 VSUBS 0.008289f
C731 B.n691 VSUBS 0.008289f
C732 B.n692 VSUBS 0.008289f
C733 B.n693 VSUBS 0.008289f
C734 B.n694 VSUBS 0.008289f
C735 B.n695 VSUBS 0.008289f
C736 B.n696 VSUBS 0.008289f
C737 B.n697 VSUBS 0.008289f
C738 B.n698 VSUBS 0.008289f
C739 B.n699 VSUBS 0.008289f
C740 B.n700 VSUBS 0.008289f
C741 B.n701 VSUBS 0.008289f
C742 B.n702 VSUBS 0.008289f
C743 B.n703 VSUBS 0.008289f
C744 B.n704 VSUBS 0.008289f
C745 B.n705 VSUBS 0.008289f
C746 B.n706 VSUBS 0.008289f
C747 B.n707 VSUBS 0.008289f
C748 B.n708 VSUBS 0.008289f
C749 B.n709 VSUBS 0.008289f
C750 B.n710 VSUBS 0.008289f
C751 B.n711 VSUBS 0.008289f
C752 B.n712 VSUBS 0.008289f
C753 B.n713 VSUBS 0.008289f
C754 B.n714 VSUBS 0.008289f
C755 B.n715 VSUBS 0.008289f
C756 B.n716 VSUBS 0.008289f
C757 B.n717 VSUBS 0.008289f
C758 B.n718 VSUBS 0.008289f
C759 B.n719 VSUBS 0.008289f
C760 B.n720 VSUBS 0.008289f
C761 B.n721 VSUBS 0.008289f
C762 B.n722 VSUBS 0.008289f
C763 B.n723 VSUBS 0.008289f
C764 B.n724 VSUBS 0.008289f
C765 B.n725 VSUBS 0.008289f
C766 B.n726 VSUBS 0.008289f
C767 B.n727 VSUBS 0.008289f
C768 B.n728 VSUBS 0.008289f
C769 B.n729 VSUBS 0.019587f
C770 B.n730 VSUBS 0.019587f
C771 B.n731 VSUBS 0.018935f
C772 B.n732 VSUBS 0.008289f
C773 B.n733 VSUBS 0.008289f
C774 B.n734 VSUBS 0.008289f
C775 B.n735 VSUBS 0.008289f
C776 B.n736 VSUBS 0.008289f
C777 B.n737 VSUBS 0.008289f
C778 B.n738 VSUBS 0.008289f
C779 B.n739 VSUBS 0.008289f
C780 B.n740 VSUBS 0.008289f
C781 B.n741 VSUBS 0.008289f
C782 B.n742 VSUBS 0.008289f
C783 B.n743 VSUBS 0.008289f
C784 B.n744 VSUBS 0.008289f
C785 B.n745 VSUBS 0.008289f
C786 B.n746 VSUBS 0.008289f
C787 B.n747 VSUBS 0.008289f
C788 B.n748 VSUBS 0.008289f
C789 B.n749 VSUBS 0.008289f
C790 B.n750 VSUBS 0.008289f
C791 B.n751 VSUBS 0.008289f
C792 B.n752 VSUBS 0.008289f
C793 B.n753 VSUBS 0.008289f
C794 B.n754 VSUBS 0.008289f
C795 B.n755 VSUBS 0.008289f
C796 B.n756 VSUBS 0.008289f
C797 B.n757 VSUBS 0.008289f
C798 B.n758 VSUBS 0.008289f
C799 B.n759 VSUBS 0.008289f
C800 B.n760 VSUBS 0.008289f
C801 B.n761 VSUBS 0.008289f
C802 B.n762 VSUBS 0.008289f
C803 B.n763 VSUBS 0.008289f
C804 B.n764 VSUBS 0.008289f
C805 B.n765 VSUBS 0.008289f
C806 B.n766 VSUBS 0.008289f
C807 B.n767 VSUBS 0.010817f
C808 B.n768 VSUBS 0.011523f
C809 B.n769 VSUBS 0.022915f
C810 VDD1.n0 VSUBS 0.030919f
C811 VDD1.n1 VSUBS 0.027093f
C812 VDD1.n2 VSUBS 0.014558f
C813 VDD1.n3 VSUBS 0.034411f
C814 VDD1.n4 VSUBS 0.015415f
C815 VDD1.n5 VSUBS 0.027093f
C816 VDD1.n6 VSUBS 0.014558f
C817 VDD1.n7 VSUBS 0.034411f
C818 VDD1.n8 VSUBS 0.015415f
C819 VDD1.n9 VSUBS 0.027093f
C820 VDD1.n10 VSUBS 0.014558f
C821 VDD1.n11 VSUBS 0.034411f
C822 VDD1.n12 VSUBS 0.014987f
C823 VDD1.n13 VSUBS 0.027093f
C824 VDD1.n14 VSUBS 0.014987f
C825 VDD1.n15 VSUBS 0.014558f
C826 VDD1.n16 VSUBS 0.034411f
C827 VDD1.n17 VSUBS 0.034411f
C828 VDD1.n18 VSUBS 0.015415f
C829 VDD1.n19 VSUBS 0.027093f
C830 VDD1.n20 VSUBS 0.014558f
C831 VDD1.n21 VSUBS 0.034411f
C832 VDD1.n22 VSUBS 0.015415f
C833 VDD1.n23 VSUBS 0.027093f
C834 VDD1.n24 VSUBS 0.014558f
C835 VDD1.n25 VSUBS 0.034411f
C836 VDD1.n26 VSUBS 0.015415f
C837 VDD1.n27 VSUBS 0.027093f
C838 VDD1.n28 VSUBS 0.014558f
C839 VDD1.n29 VSUBS 0.034411f
C840 VDD1.n30 VSUBS 0.015415f
C841 VDD1.n31 VSUBS 0.027093f
C842 VDD1.n32 VSUBS 0.014558f
C843 VDD1.n33 VSUBS 0.034411f
C844 VDD1.n34 VSUBS 0.015415f
C845 VDD1.n35 VSUBS 2.30922f
C846 VDD1.n36 VSUBS 0.014558f
C847 VDD1.t3 VSUBS 0.073984f
C848 VDD1.n37 VSUBS 0.228618f
C849 VDD1.n38 VSUBS 0.02189f
C850 VDD1.n39 VSUBS 0.025808f
C851 VDD1.n40 VSUBS 0.034411f
C852 VDD1.n41 VSUBS 0.015415f
C853 VDD1.n42 VSUBS 0.014558f
C854 VDD1.n43 VSUBS 0.027093f
C855 VDD1.n44 VSUBS 0.027093f
C856 VDD1.n45 VSUBS 0.014558f
C857 VDD1.n46 VSUBS 0.015415f
C858 VDD1.n47 VSUBS 0.034411f
C859 VDD1.n48 VSUBS 0.034411f
C860 VDD1.n49 VSUBS 0.015415f
C861 VDD1.n50 VSUBS 0.014558f
C862 VDD1.n51 VSUBS 0.027093f
C863 VDD1.n52 VSUBS 0.027093f
C864 VDD1.n53 VSUBS 0.014558f
C865 VDD1.n54 VSUBS 0.015415f
C866 VDD1.n55 VSUBS 0.034411f
C867 VDD1.n56 VSUBS 0.034411f
C868 VDD1.n57 VSUBS 0.015415f
C869 VDD1.n58 VSUBS 0.014558f
C870 VDD1.n59 VSUBS 0.027093f
C871 VDD1.n60 VSUBS 0.027093f
C872 VDD1.n61 VSUBS 0.014558f
C873 VDD1.n62 VSUBS 0.015415f
C874 VDD1.n63 VSUBS 0.034411f
C875 VDD1.n64 VSUBS 0.034411f
C876 VDD1.n65 VSUBS 0.015415f
C877 VDD1.n66 VSUBS 0.014558f
C878 VDD1.n67 VSUBS 0.027093f
C879 VDD1.n68 VSUBS 0.027093f
C880 VDD1.n69 VSUBS 0.014558f
C881 VDD1.n70 VSUBS 0.015415f
C882 VDD1.n71 VSUBS 0.034411f
C883 VDD1.n72 VSUBS 0.034411f
C884 VDD1.n73 VSUBS 0.015415f
C885 VDD1.n74 VSUBS 0.014558f
C886 VDD1.n75 VSUBS 0.027093f
C887 VDD1.n76 VSUBS 0.027093f
C888 VDD1.n77 VSUBS 0.014558f
C889 VDD1.n78 VSUBS 0.015415f
C890 VDD1.n79 VSUBS 0.034411f
C891 VDD1.n80 VSUBS 0.034411f
C892 VDD1.n81 VSUBS 0.015415f
C893 VDD1.n82 VSUBS 0.014558f
C894 VDD1.n83 VSUBS 0.027093f
C895 VDD1.n84 VSUBS 0.027093f
C896 VDD1.n85 VSUBS 0.014558f
C897 VDD1.n86 VSUBS 0.015415f
C898 VDD1.n87 VSUBS 0.034411f
C899 VDD1.n88 VSUBS 0.034411f
C900 VDD1.n89 VSUBS 0.015415f
C901 VDD1.n90 VSUBS 0.014558f
C902 VDD1.n91 VSUBS 0.027093f
C903 VDD1.n92 VSUBS 0.027093f
C904 VDD1.n93 VSUBS 0.014558f
C905 VDD1.n94 VSUBS 0.015415f
C906 VDD1.n95 VSUBS 0.034411f
C907 VDD1.n96 VSUBS 0.034411f
C908 VDD1.n97 VSUBS 0.015415f
C909 VDD1.n98 VSUBS 0.014558f
C910 VDD1.n99 VSUBS 0.027093f
C911 VDD1.n100 VSUBS 0.027093f
C912 VDD1.n101 VSUBS 0.014558f
C913 VDD1.n102 VSUBS 0.015415f
C914 VDD1.n103 VSUBS 0.034411f
C915 VDD1.n104 VSUBS 0.087222f
C916 VDD1.n105 VSUBS 0.015415f
C917 VDD1.n106 VSUBS 0.014558f
C918 VDD1.n107 VSUBS 0.063734f
C919 VDD1.n108 VSUBS 0.065585f
C920 VDD1.n109 VSUBS 0.030919f
C921 VDD1.n110 VSUBS 0.027093f
C922 VDD1.n111 VSUBS 0.014558f
C923 VDD1.n112 VSUBS 0.034411f
C924 VDD1.n113 VSUBS 0.015415f
C925 VDD1.n114 VSUBS 0.027093f
C926 VDD1.n115 VSUBS 0.014558f
C927 VDD1.n116 VSUBS 0.034411f
C928 VDD1.n117 VSUBS 0.015415f
C929 VDD1.n118 VSUBS 0.027093f
C930 VDD1.n119 VSUBS 0.014558f
C931 VDD1.n120 VSUBS 0.034411f
C932 VDD1.n121 VSUBS 0.014987f
C933 VDD1.n122 VSUBS 0.027093f
C934 VDD1.n123 VSUBS 0.015415f
C935 VDD1.n124 VSUBS 0.034411f
C936 VDD1.n125 VSUBS 0.015415f
C937 VDD1.n126 VSUBS 0.027093f
C938 VDD1.n127 VSUBS 0.014558f
C939 VDD1.n128 VSUBS 0.034411f
C940 VDD1.n129 VSUBS 0.015415f
C941 VDD1.n130 VSUBS 0.027093f
C942 VDD1.n131 VSUBS 0.014558f
C943 VDD1.n132 VSUBS 0.034411f
C944 VDD1.n133 VSUBS 0.015415f
C945 VDD1.n134 VSUBS 0.027093f
C946 VDD1.n135 VSUBS 0.014558f
C947 VDD1.n136 VSUBS 0.034411f
C948 VDD1.n137 VSUBS 0.015415f
C949 VDD1.n138 VSUBS 0.027093f
C950 VDD1.n139 VSUBS 0.014558f
C951 VDD1.n140 VSUBS 0.034411f
C952 VDD1.n141 VSUBS 0.015415f
C953 VDD1.n142 VSUBS 2.30922f
C954 VDD1.n143 VSUBS 0.014558f
C955 VDD1.t2 VSUBS 0.073984f
C956 VDD1.n144 VSUBS 0.228618f
C957 VDD1.n145 VSUBS 0.02189f
C958 VDD1.n146 VSUBS 0.025808f
C959 VDD1.n147 VSUBS 0.034411f
C960 VDD1.n148 VSUBS 0.015415f
C961 VDD1.n149 VSUBS 0.014558f
C962 VDD1.n150 VSUBS 0.027093f
C963 VDD1.n151 VSUBS 0.027093f
C964 VDD1.n152 VSUBS 0.014558f
C965 VDD1.n153 VSUBS 0.015415f
C966 VDD1.n154 VSUBS 0.034411f
C967 VDD1.n155 VSUBS 0.034411f
C968 VDD1.n156 VSUBS 0.015415f
C969 VDD1.n157 VSUBS 0.014558f
C970 VDD1.n158 VSUBS 0.027093f
C971 VDD1.n159 VSUBS 0.027093f
C972 VDD1.n160 VSUBS 0.014558f
C973 VDD1.n161 VSUBS 0.015415f
C974 VDD1.n162 VSUBS 0.034411f
C975 VDD1.n163 VSUBS 0.034411f
C976 VDD1.n164 VSUBS 0.015415f
C977 VDD1.n165 VSUBS 0.014558f
C978 VDD1.n166 VSUBS 0.027093f
C979 VDD1.n167 VSUBS 0.027093f
C980 VDD1.n168 VSUBS 0.014558f
C981 VDD1.n169 VSUBS 0.015415f
C982 VDD1.n170 VSUBS 0.034411f
C983 VDD1.n171 VSUBS 0.034411f
C984 VDD1.n172 VSUBS 0.015415f
C985 VDD1.n173 VSUBS 0.014558f
C986 VDD1.n174 VSUBS 0.027093f
C987 VDD1.n175 VSUBS 0.027093f
C988 VDD1.n176 VSUBS 0.014558f
C989 VDD1.n177 VSUBS 0.015415f
C990 VDD1.n178 VSUBS 0.034411f
C991 VDD1.n179 VSUBS 0.034411f
C992 VDD1.n180 VSUBS 0.015415f
C993 VDD1.n181 VSUBS 0.014558f
C994 VDD1.n182 VSUBS 0.027093f
C995 VDD1.n183 VSUBS 0.027093f
C996 VDD1.n184 VSUBS 0.014558f
C997 VDD1.n185 VSUBS 0.014558f
C998 VDD1.n186 VSUBS 0.015415f
C999 VDD1.n187 VSUBS 0.034411f
C1000 VDD1.n188 VSUBS 0.034411f
C1001 VDD1.n189 VSUBS 0.034411f
C1002 VDD1.n190 VSUBS 0.014987f
C1003 VDD1.n191 VSUBS 0.014558f
C1004 VDD1.n192 VSUBS 0.027093f
C1005 VDD1.n193 VSUBS 0.027093f
C1006 VDD1.n194 VSUBS 0.014558f
C1007 VDD1.n195 VSUBS 0.015415f
C1008 VDD1.n196 VSUBS 0.034411f
C1009 VDD1.n197 VSUBS 0.034411f
C1010 VDD1.n198 VSUBS 0.015415f
C1011 VDD1.n199 VSUBS 0.014558f
C1012 VDD1.n200 VSUBS 0.027093f
C1013 VDD1.n201 VSUBS 0.027093f
C1014 VDD1.n202 VSUBS 0.014558f
C1015 VDD1.n203 VSUBS 0.015415f
C1016 VDD1.n204 VSUBS 0.034411f
C1017 VDD1.n205 VSUBS 0.034411f
C1018 VDD1.n206 VSUBS 0.015415f
C1019 VDD1.n207 VSUBS 0.014558f
C1020 VDD1.n208 VSUBS 0.027093f
C1021 VDD1.n209 VSUBS 0.027093f
C1022 VDD1.n210 VSUBS 0.014558f
C1023 VDD1.n211 VSUBS 0.015415f
C1024 VDD1.n212 VSUBS 0.034411f
C1025 VDD1.n213 VSUBS 0.087222f
C1026 VDD1.n214 VSUBS 0.015415f
C1027 VDD1.n215 VSUBS 0.014558f
C1028 VDD1.n216 VSUBS 0.063734f
C1029 VDD1.n217 VSUBS 0.06511f
C1030 VDD1.t5 VSUBS 0.421979f
C1031 VDD1.t4 VSUBS 0.421979f
C1032 VDD1.n218 VSUBS 3.54746f
C1033 VDD1.n219 VSUBS 3.14921f
C1034 VDD1.t1 VSUBS 0.421979f
C1035 VDD1.t0 VSUBS 0.421979f
C1036 VDD1.n220 VSUBS 3.54486f
C1037 VDD1.n221 VSUBS 3.53053f
C1038 VP.n0 VSUBS 0.057912f
C1039 VP.t0 VSUBS 2.68666f
C1040 VP.n1 VSUBS 0.060007f
C1041 VP.n2 VSUBS 0.244831f
C1042 VP.t5 VSUBS 2.76246f
C1043 VP.t4 VSUBS 2.68666f
C1044 VP.t2 VSUBS 2.81357f
C1045 VP.n3 VSUBS 1.00797f
C1046 VP.n4 VSUBS 1.02405f
C1047 VP.n5 VSUBS 0.060007f
C1048 VP.n6 VSUBS 1.02909f
C1049 VP.n7 VSUBS 2.30544f
C1050 VP.t3 VSUBS 2.76246f
C1051 VP.n8 VSUBS 1.02909f
C1052 VP.n9 VSUBS 2.33727f
C1053 VP.n10 VSUBS 0.057912f
C1054 VP.n11 VSUBS 0.0434f
C1055 VP.n12 VSUBS 0.991847f
C1056 VP.n13 VSUBS 0.060007f
C1057 VP.t1 VSUBS 2.76246f
C1058 VP.n14 VSUBS 1.02909f
C1059 VP.n15 VSUBS 0.040646f
C1060 VTAIL.t7 VSUBS 0.423701f
C1061 VTAIL.t11 VSUBS 0.423701f
C1062 VTAIL.n0 VSUBS 3.38735f
C1063 VTAIL.n1 VSUBS 0.806071f
C1064 VTAIL.n2 VSUBS 0.031045f
C1065 VTAIL.n3 VSUBS 0.027203f
C1066 VTAIL.n4 VSUBS 0.014618f
C1067 VTAIL.n5 VSUBS 0.034551f
C1068 VTAIL.n6 VSUBS 0.015478f
C1069 VTAIL.n7 VSUBS 0.027203f
C1070 VTAIL.n8 VSUBS 0.014618f
C1071 VTAIL.n9 VSUBS 0.034551f
C1072 VTAIL.n10 VSUBS 0.015478f
C1073 VTAIL.n11 VSUBS 0.027203f
C1074 VTAIL.n12 VSUBS 0.014618f
C1075 VTAIL.n13 VSUBS 0.034551f
C1076 VTAIL.n14 VSUBS 0.015048f
C1077 VTAIL.n15 VSUBS 0.027203f
C1078 VTAIL.n16 VSUBS 0.015478f
C1079 VTAIL.n17 VSUBS 0.034551f
C1080 VTAIL.n18 VSUBS 0.015478f
C1081 VTAIL.n19 VSUBS 0.027203f
C1082 VTAIL.n20 VSUBS 0.014618f
C1083 VTAIL.n21 VSUBS 0.034551f
C1084 VTAIL.n22 VSUBS 0.015478f
C1085 VTAIL.n23 VSUBS 0.027203f
C1086 VTAIL.n24 VSUBS 0.014618f
C1087 VTAIL.n25 VSUBS 0.034551f
C1088 VTAIL.n26 VSUBS 0.015478f
C1089 VTAIL.n27 VSUBS 0.027203f
C1090 VTAIL.n28 VSUBS 0.014618f
C1091 VTAIL.n29 VSUBS 0.034551f
C1092 VTAIL.n30 VSUBS 0.015478f
C1093 VTAIL.n31 VSUBS 0.027203f
C1094 VTAIL.n32 VSUBS 0.014618f
C1095 VTAIL.n33 VSUBS 0.034551f
C1096 VTAIL.n34 VSUBS 0.015478f
C1097 VTAIL.n35 VSUBS 2.31864f
C1098 VTAIL.n36 VSUBS 0.014618f
C1099 VTAIL.t3 VSUBS 0.074286f
C1100 VTAIL.n37 VSUBS 0.229551f
C1101 VTAIL.n38 VSUBS 0.02198f
C1102 VTAIL.n39 VSUBS 0.025913f
C1103 VTAIL.n40 VSUBS 0.034551f
C1104 VTAIL.n41 VSUBS 0.015478f
C1105 VTAIL.n42 VSUBS 0.014618f
C1106 VTAIL.n43 VSUBS 0.027203f
C1107 VTAIL.n44 VSUBS 0.027203f
C1108 VTAIL.n45 VSUBS 0.014618f
C1109 VTAIL.n46 VSUBS 0.015478f
C1110 VTAIL.n47 VSUBS 0.034551f
C1111 VTAIL.n48 VSUBS 0.034551f
C1112 VTAIL.n49 VSUBS 0.015478f
C1113 VTAIL.n50 VSUBS 0.014618f
C1114 VTAIL.n51 VSUBS 0.027203f
C1115 VTAIL.n52 VSUBS 0.027203f
C1116 VTAIL.n53 VSUBS 0.014618f
C1117 VTAIL.n54 VSUBS 0.015478f
C1118 VTAIL.n55 VSUBS 0.034551f
C1119 VTAIL.n56 VSUBS 0.034551f
C1120 VTAIL.n57 VSUBS 0.015478f
C1121 VTAIL.n58 VSUBS 0.014618f
C1122 VTAIL.n59 VSUBS 0.027203f
C1123 VTAIL.n60 VSUBS 0.027203f
C1124 VTAIL.n61 VSUBS 0.014618f
C1125 VTAIL.n62 VSUBS 0.015478f
C1126 VTAIL.n63 VSUBS 0.034551f
C1127 VTAIL.n64 VSUBS 0.034551f
C1128 VTAIL.n65 VSUBS 0.015478f
C1129 VTAIL.n66 VSUBS 0.014618f
C1130 VTAIL.n67 VSUBS 0.027203f
C1131 VTAIL.n68 VSUBS 0.027203f
C1132 VTAIL.n69 VSUBS 0.014618f
C1133 VTAIL.n70 VSUBS 0.015478f
C1134 VTAIL.n71 VSUBS 0.034551f
C1135 VTAIL.n72 VSUBS 0.034551f
C1136 VTAIL.n73 VSUBS 0.015478f
C1137 VTAIL.n74 VSUBS 0.014618f
C1138 VTAIL.n75 VSUBS 0.027203f
C1139 VTAIL.n76 VSUBS 0.027203f
C1140 VTAIL.n77 VSUBS 0.014618f
C1141 VTAIL.n78 VSUBS 0.014618f
C1142 VTAIL.n79 VSUBS 0.015478f
C1143 VTAIL.n80 VSUBS 0.034551f
C1144 VTAIL.n81 VSUBS 0.034551f
C1145 VTAIL.n82 VSUBS 0.034551f
C1146 VTAIL.n83 VSUBS 0.015048f
C1147 VTAIL.n84 VSUBS 0.014618f
C1148 VTAIL.n85 VSUBS 0.027203f
C1149 VTAIL.n86 VSUBS 0.027203f
C1150 VTAIL.n87 VSUBS 0.014618f
C1151 VTAIL.n88 VSUBS 0.015478f
C1152 VTAIL.n89 VSUBS 0.034551f
C1153 VTAIL.n90 VSUBS 0.034551f
C1154 VTAIL.n91 VSUBS 0.015478f
C1155 VTAIL.n92 VSUBS 0.014618f
C1156 VTAIL.n93 VSUBS 0.027203f
C1157 VTAIL.n94 VSUBS 0.027203f
C1158 VTAIL.n95 VSUBS 0.014618f
C1159 VTAIL.n96 VSUBS 0.015478f
C1160 VTAIL.n97 VSUBS 0.034551f
C1161 VTAIL.n98 VSUBS 0.034551f
C1162 VTAIL.n99 VSUBS 0.015478f
C1163 VTAIL.n100 VSUBS 0.014618f
C1164 VTAIL.n101 VSUBS 0.027203f
C1165 VTAIL.n102 VSUBS 0.027203f
C1166 VTAIL.n103 VSUBS 0.014618f
C1167 VTAIL.n104 VSUBS 0.015478f
C1168 VTAIL.n105 VSUBS 0.034551f
C1169 VTAIL.n106 VSUBS 0.087578f
C1170 VTAIL.n107 VSUBS 0.015478f
C1171 VTAIL.n108 VSUBS 0.014618f
C1172 VTAIL.n109 VSUBS 0.063994f
C1173 VTAIL.n110 VSUBS 0.044251f
C1174 VTAIL.n111 VSUBS 0.231665f
C1175 VTAIL.t4 VSUBS 0.423701f
C1176 VTAIL.t2 VSUBS 0.423701f
C1177 VTAIL.n112 VSUBS 3.38735f
C1178 VTAIL.n113 VSUBS 2.86861f
C1179 VTAIL.t8 VSUBS 0.423701f
C1180 VTAIL.t9 VSUBS 0.423701f
C1181 VTAIL.n114 VSUBS 3.38737f
C1182 VTAIL.n115 VSUBS 2.86859f
C1183 VTAIL.n116 VSUBS 0.031045f
C1184 VTAIL.n117 VSUBS 0.027203f
C1185 VTAIL.n118 VSUBS 0.014618f
C1186 VTAIL.n119 VSUBS 0.034551f
C1187 VTAIL.n120 VSUBS 0.015478f
C1188 VTAIL.n121 VSUBS 0.027203f
C1189 VTAIL.n122 VSUBS 0.014618f
C1190 VTAIL.n123 VSUBS 0.034551f
C1191 VTAIL.n124 VSUBS 0.015478f
C1192 VTAIL.n125 VSUBS 0.027203f
C1193 VTAIL.n126 VSUBS 0.014618f
C1194 VTAIL.n127 VSUBS 0.034551f
C1195 VTAIL.n128 VSUBS 0.015048f
C1196 VTAIL.n129 VSUBS 0.027203f
C1197 VTAIL.n130 VSUBS 0.015048f
C1198 VTAIL.n131 VSUBS 0.014618f
C1199 VTAIL.n132 VSUBS 0.034551f
C1200 VTAIL.n133 VSUBS 0.034551f
C1201 VTAIL.n134 VSUBS 0.015478f
C1202 VTAIL.n135 VSUBS 0.027203f
C1203 VTAIL.n136 VSUBS 0.014618f
C1204 VTAIL.n137 VSUBS 0.034551f
C1205 VTAIL.n138 VSUBS 0.015478f
C1206 VTAIL.n139 VSUBS 0.027203f
C1207 VTAIL.n140 VSUBS 0.014618f
C1208 VTAIL.n141 VSUBS 0.034551f
C1209 VTAIL.n142 VSUBS 0.015478f
C1210 VTAIL.n143 VSUBS 0.027203f
C1211 VTAIL.n144 VSUBS 0.014618f
C1212 VTAIL.n145 VSUBS 0.034551f
C1213 VTAIL.n146 VSUBS 0.015478f
C1214 VTAIL.n147 VSUBS 0.027203f
C1215 VTAIL.n148 VSUBS 0.014618f
C1216 VTAIL.n149 VSUBS 0.034551f
C1217 VTAIL.n150 VSUBS 0.015478f
C1218 VTAIL.n151 VSUBS 2.31864f
C1219 VTAIL.n152 VSUBS 0.014618f
C1220 VTAIL.t10 VSUBS 0.074286f
C1221 VTAIL.n153 VSUBS 0.229551f
C1222 VTAIL.n154 VSUBS 0.02198f
C1223 VTAIL.n155 VSUBS 0.025913f
C1224 VTAIL.n156 VSUBS 0.034551f
C1225 VTAIL.n157 VSUBS 0.015478f
C1226 VTAIL.n158 VSUBS 0.014618f
C1227 VTAIL.n159 VSUBS 0.027203f
C1228 VTAIL.n160 VSUBS 0.027203f
C1229 VTAIL.n161 VSUBS 0.014618f
C1230 VTAIL.n162 VSUBS 0.015478f
C1231 VTAIL.n163 VSUBS 0.034551f
C1232 VTAIL.n164 VSUBS 0.034551f
C1233 VTAIL.n165 VSUBS 0.015478f
C1234 VTAIL.n166 VSUBS 0.014618f
C1235 VTAIL.n167 VSUBS 0.027203f
C1236 VTAIL.n168 VSUBS 0.027203f
C1237 VTAIL.n169 VSUBS 0.014618f
C1238 VTAIL.n170 VSUBS 0.015478f
C1239 VTAIL.n171 VSUBS 0.034551f
C1240 VTAIL.n172 VSUBS 0.034551f
C1241 VTAIL.n173 VSUBS 0.015478f
C1242 VTAIL.n174 VSUBS 0.014618f
C1243 VTAIL.n175 VSUBS 0.027203f
C1244 VTAIL.n176 VSUBS 0.027203f
C1245 VTAIL.n177 VSUBS 0.014618f
C1246 VTAIL.n178 VSUBS 0.015478f
C1247 VTAIL.n179 VSUBS 0.034551f
C1248 VTAIL.n180 VSUBS 0.034551f
C1249 VTAIL.n181 VSUBS 0.015478f
C1250 VTAIL.n182 VSUBS 0.014618f
C1251 VTAIL.n183 VSUBS 0.027203f
C1252 VTAIL.n184 VSUBS 0.027203f
C1253 VTAIL.n185 VSUBS 0.014618f
C1254 VTAIL.n186 VSUBS 0.015478f
C1255 VTAIL.n187 VSUBS 0.034551f
C1256 VTAIL.n188 VSUBS 0.034551f
C1257 VTAIL.n189 VSUBS 0.015478f
C1258 VTAIL.n190 VSUBS 0.014618f
C1259 VTAIL.n191 VSUBS 0.027203f
C1260 VTAIL.n192 VSUBS 0.027203f
C1261 VTAIL.n193 VSUBS 0.014618f
C1262 VTAIL.n194 VSUBS 0.015478f
C1263 VTAIL.n195 VSUBS 0.034551f
C1264 VTAIL.n196 VSUBS 0.034551f
C1265 VTAIL.n197 VSUBS 0.015478f
C1266 VTAIL.n198 VSUBS 0.014618f
C1267 VTAIL.n199 VSUBS 0.027203f
C1268 VTAIL.n200 VSUBS 0.027203f
C1269 VTAIL.n201 VSUBS 0.014618f
C1270 VTAIL.n202 VSUBS 0.015478f
C1271 VTAIL.n203 VSUBS 0.034551f
C1272 VTAIL.n204 VSUBS 0.034551f
C1273 VTAIL.n205 VSUBS 0.015478f
C1274 VTAIL.n206 VSUBS 0.014618f
C1275 VTAIL.n207 VSUBS 0.027203f
C1276 VTAIL.n208 VSUBS 0.027203f
C1277 VTAIL.n209 VSUBS 0.014618f
C1278 VTAIL.n210 VSUBS 0.015478f
C1279 VTAIL.n211 VSUBS 0.034551f
C1280 VTAIL.n212 VSUBS 0.034551f
C1281 VTAIL.n213 VSUBS 0.015478f
C1282 VTAIL.n214 VSUBS 0.014618f
C1283 VTAIL.n215 VSUBS 0.027203f
C1284 VTAIL.n216 VSUBS 0.027203f
C1285 VTAIL.n217 VSUBS 0.014618f
C1286 VTAIL.n218 VSUBS 0.015478f
C1287 VTAIL.n219 VSUBS 0.034551f
C1288 VTAIL.n220 VSUBS 0.087578f
C1289 VTAIL.n221 VSUBS 0.015478f
C1290 VTAIL.n222 VSUBS 0.014618f
C1291 VTAIL.n223 VSUBS 0.063994f
C1292 VTAIL.n224 VSUBS 0.044251f
C1293 VTAIL.n225 VSUBS 0.231665f
C1294 VTAIL.t0 VSUBS 0.423701f
C1295 VTAIL.t1 VSUBS 0.423701f
C1296 VTAIL.n226 VSUBS 3.38737f
C1297 VTAIL.n227 VSUBS 0.884261f
C1298 VTAIL.n228 VSUBS 0.031045f
C1299 VTAIL.n229 VSUBS 0.027203f
C1300 VTAIL.n230 VSUBS 0.014618f
C1301 VTAIL.n231 VSUBS 0.034551f
C1302 VTAIL.n232 VSUBS 0.015478f
C1303 VTAIL.n233 VSUBS 0.027203f
C1304 VTAIL.n234 VSUBS 0.014618f
C1305 VTAIL.n235 VSUBS 0.034551f
C1306 VTAIL.n236 VSUBS 0.015478f
C1307 VTAIL.n237 VSUBS 0.027203f
C1308 VTAIL.n238 VSUBS 0.014618f
C1309 VTAIL.n239 VSUBS 0.034551f
C1310 VTAIL.n240 VSUBS 0.015048f
C1311 VTAIL.n241 VSUBS 0.027203f
C1312 VTAIL.n242 VSUBS 0.015048f
C1313 VTAIL.n243 VSUBS 0.014618f
C1314 VTAIL.n244 VSUBS 0.034551f
C1315 VTAIL.n245 VSUBS 0.034551f
C1316 VTAIL.n246 VSUBS 0.015478f
C1317 VTAIL.n247 VSUBS 0.027203f
C1318 VTAIL.n248 VSUBS 0.014618f
C1319 VTAIL.n249 VSUBS 0.034551f
C1320 VTAIL.n250 VSUBS 0.015478f
C1321 VTAIL.n251 VSUBS 0.027203f
C1322 VTAIL.n252 VSUBS 0.014618f
C1323 VTAIL.n253 VSUBS 0.034551f
C1324 VTAIL.n254 VSUBS 0.015478f
C1325 VTAIL.n255 VSUBS 0.027203f
C1326 VTAIL.n256 VSUBS 0.014618f
C1327 VTAIL.n257 VSUBS 0.034551f
C1328 VTAIL.n258 VSUBS 0.015478f
C1329 VTAIL.n259 VSUBS 0.027203f
C1330 VTAIL.n260 VSUBS 0.014618f
C1331 VTAIL.n261 VSUBS 0.034551f
C1332 VTAIL.n262 VSUBS 0.015478f
C1333 VTAIL.n263 VSUBS 2.31864f
C1334 VTAIL.n264 VSUBS 0.014618f
C1335 VTAIL.t5 VSUBS 0.074286f
C1336 VTAIL.n265 VSUBS 0.229551f
C1337 VTAIL.n266 VSUBS 0.02198f
C1338 VTAIL.n267 VSUBS 0.025913f
C1339 VTAIL.n268 VSUBS 0.034551f
C1340 VTAIL.n269 VSUBS 0.015478f
C1341 VTAIL.n270 VSUBS 0.014618f
C1342 VTAIL.n271 VSUBS 0.027203f
C1343 VTAIL.n272 VSUBS 0.027203f
C1344 VTAIL.n273 VSUBS 0.014618f
C1345 VTAIL.n274 VSUBS 0.015478f
C1346 VTAIL.n275 VSUBS 0.034551f
C1347 VTAIL.n276 VSUBS 0.034551f
C1348 VTAIL.n277 VSUBS 0.015478f
C1349 VTAIL.n278 VSUBS 0.014618f
C1350 VTAIL.n279 VSUBS 0.027203f
C1351 VTAIL.n280 VSUBS 0.027203f
C1352 VTAIL.n281 VSUBS 0.014618f
C1353 VTAIL.n282 VSUBS 0.015478f
C1354 VTAIL.n283 VSUBS 0.034551f
C1355 VTAIL.n284 VSUBS 0.034551f
C1356 VTAIL.n285 VSUBS 0.015478f
C1357 VTAIL.n286 VSUBS 0.014618f
C1358 VTAIL.n287 VSUBS 0.027203f
C1359 VTAIL.n288 VSUBS 0.027203f
C1360 VTAIL.n289 VSUBS 0.014618f
C1361 VTAIL.n290 VSUBS 0.015478f
C1362 VTAIL.n291 VSUBS 0.034551f
C1363 VTAIL.n292 VSUBS 0.034551f
C1364 VTAIL.n293 VSUBS 0.015478f
C1365 VTAIL.n294 VSUBS 0.014618f
C1366 VTAIL.n295 VSUBS 0.027203f
C1367 VTAIL.n296 VSUBS 0.027203f
C1368 VTAIL.n297 VSUBS 0.014618f
C1369 VTAIL.n298 VSUBS 0.015478f
C1370 VTAIL.n299 VSUBS 0.034551f
C1371 VTAIL.n300 VSUBS 0.034551f
C1372 VTAIL.n301 VSUBS 0.015478f
C1373 VTAIL.n302 VSUBS 0.014618f
C1374 VTAIL.n303 VSUBS 0.027203f
C1375 VTAIL.n304 VSUBS 0.027203f
C1376 VTAIL.n305 VSUBS 0.014618f
C1377 VTAIL.n306 VSUBS 0.015478f
C1378 VTAIL.n307 VSUBS 0.034551f
C1379 VTAIL.n308 VSUBS 0.034551f
C1380 VTAIL.n309 VSUBS 0.015478f
C1381 VTAIL.n310 VSUBS 0.014618f
C1382 VTAIL.n311 VSUBS 0.027203f
C1383 VTAIL.n312 VSUBS 0.027203f
C1384 VTAIL.n313 VSUBS 0.014618f
C1385 VTAIL.n314 VSUBS 0.015478f
C1386 VTAIL.n315 VSUBS 0.034551f
C1387 VTAIL.n316 VSUBS 0.034551f
C1388 VTAIL.n317 VSUBS 0.015478f
C1389 VTAIL.n318 VSUBS 0.014618f
C1390 VTAIL.n319 VSUBS 0.027203f
C1391 VTAIL.n320 VSUBS 0.027203f
C1392 VTAIL.n321 VSUBS 0.014618f
C1393 VTAIL.n322 VSUBS 0.015478f
C1394 VTAIL.n323 VSUBS 0.034551f
C1395 VTAIL.n324 VSUBS 0.034551f
C1396 VTAIL.n325 VSUBS 0.015478f
C1397 VTAIL.n326 VSUBS 0.014618f
C1398 VTAIL.n327 VSUBS 0.027203f
C1399 VTAIL.n328 VSUBS 0.027203f
C1400 VTAIL.n329 VSUBS 0.014618f
C1401 VTAIL.n330 VSUBS 0.015478f
C1402 VTAIL.n331 VSUBS 0.034551f
C1403 VTAIL.n332 VSUBS 0.087578f
C1404 VTAIL.n333 VSUBS 0.015478f
C1405 VTAIL.n334 VSUBS 0.014618f
C1406 VTAIL.n335 VSUBS 0.063994f
C1407 VTAIL.n336 VSUBS 0.044251f
C1408 VTAIL.n337 VSUBS 2.10492f
C1409 VTAIL.n338 VSUBS 0.031045f
C1410 VTAIL.n339 VSUBS 0.027203f
C1411 VTAIL.n340 VSUBS 0.014618f
C1412 VTAIL.n341 VSUBS 0.034551f
C1413 VTAIL.n342 VSUBS 0.015478f
C1414 VTAIL.n343 VSUBS 0.027203f
C1415 VTAIL.n344 VSUBS 0.014618f
C1416 VTAIL.n345 VSUBS 0.034551f
C1417 VTAIL.n346 VSUBS 0.015478f
C1418 VTAIL.n347 VSUBS 0.027203f
C1419 VTAIL.n348 VSUBS 0.014618f
C1420 VTAIL.n349 VSUBS 0.034551f
C1421 VTAIL.n350 VSUBS 0.015048f
C1422 VTAIL.n351 VSUBS 0.027203f
C1423 VTAIL.n352 VSUBS 0.015478f
C1424 VTAIL.n353 VSUBS 0.034551f
C1425 VTAIL.n354 VSUBS 0.015478f
C1426 VTAIL.n355 VSUBS 0.027203f
C1427 VTAIL.n356 VSUBS 0.014618f
C1428 VTAIL.n357 VSUBS 0.034551f
C1429 VTAIL.n358 VSUBS 0.015478f
C1430 VTAIL.n359 VSUBS 0.027203f
C1431 VTAIL.n360 VSUBS 0.014618f
C1432 VTAIL.n361 VSUBS 0.034551f
C1433 VTAIL.n362 VSUBS 0.015478f
C1434 VTAIL.n363 VSUBS 0.027203f
C1435 VTAIL.n364 VSUBS 0.014618f
C1436 VTAIL.n365 VSUBS 0.034551f
C1437 VTAIL.n366 VSUBS 0.015478f
C1438 VTAIL.n367 VSUBS 0.027203f
C1439 VTAIL.n368 VSUBS 0.014618f
C1440 VTAIL.n369 VSUBS 0.034551f
C1441 VTAIL.n370 VSUBS 0.015478f
C1442 VTAIL.n371 VSUBS 2.31864f
C1443 VTAIL.n372 VSUBS 0.014618f
C1444 VTAIL.t6 VSUBS 0.074286f
C1445 VTAIL.n373 VSUBS 0.229551f
C1446 VTAIL.n374 VSUBS 0.02198f
C1447 VTAIL.n375 VSUBS 0.025913f
C1448 VTAIL.n376 VSUBS 0.034551f
C1449 VTAIL.n377 VSUBS 0.015478f
C1450 VTAIL.n378 VSUBS 0.014618f
C1451 VTAIL.n379 VSUBS 0.027203f
C1452 VTAIL.n380 VSUBS 0.027203f
C1453 VTAIL.n381 VSUBS 0.014618f
C1454 VTAIL.n382 VSUBS 0.015478f
C1455 VTAIL.n383 VSUBS 0.034551f
C1456 VTAIL.n384 VSUBS 0.034551f
C1457 VTAIL.n385 VSUBS 0.015478f
C1458 VTAIL.n386 VSUBS 0.014618f
C1459 VTAIL.n387 VSUBS 0.027203f
C1460 VTAIL.n388 VSUBS 0.027203f
C1461 VTAIL.n389 VSUBS 0.014618f
C1462 VTAIL.n390 VSUBS 0.015478f
C1463 VTAIL.n391 VSUBS 0.034551f
C1464 VTAIL.n392 VSUBS 0.034551f
C1465 VTAIL.n393 VSUBS 0.015478f
C1466 VTAIL.n394 VSUBS 0.014618f
C1467 VTAIL.n395 VSUBS 0.027203f
C1468 VTAIL.n396 VSUBS 0.027203f
C1469 VTAIL.n397 VSUBS 0.014618f
C1470 VTAIL.n398 VSUBS 0.015478f
C1471 VTAIL.n399 VSUBS 0.034551f
C1472 VTAIL.n400 VSUBS 0.034551f
C1473 VTAIL.n401 VSUBS 0.015478f
C1474 VTAIL.n402 VSUBS 0.014618f
C1475 VTAIL.n403 VSUBS 0.027203f
C1476 VTAIL.n404 VSUBS 0.027203f
C1477 VTAIL.n405 VSUBS 0.014618f
C1478 VTAIL.n406 VSUBS 0.015478f
C1479 VTAIL.n407 VSUBS 0.034551f
C1480 VTAIL.n408 VSUBS 0.034551f
C1481 VTAIL.n409 VSUBS 0.015478f
C1482 VTAIL.n410 VSUBS 0.014618f
C1483 VTAIL.n411 VSUBS 0.027203f
C1484 VTAIL.n412 VSUBS 0.027203f
C1485 VTAIL.n413 VSUBS 0.014618f
C1486 VTAIL.n414 VSUBS 0.014618f
C1487 VTAIL.n415 VSUBS 0.015478f
C1488 VTAIL.n416 VSUBS 0.034551f
C1489 VTAIL.n417 VSUBS 0.034551f
C1490 VTAIL.n418 VSUBS 0.034551f
C1491 VTAIL.n419 VSUBS 0.015048f
C1492 VTAIL.n420 VSUBS 0.014618f
C1493 VTAIL.n421 VSUBS 0.027203f
C1494 VTAIL.n422 VSUBS 0.027203f
C1495 VTAIL.n423 VSUBS 0.014618f
C1496 VTAIL.n424 VSUBS 0.015478f
C1497 VTAIL.n425 VSUBS 0.034551f
C1498 VTAIL.n426 VSUBS 0.034551f
C1499 VTAIL.n427 VSUBS 0.015478f
C1500 VTAIL.n428 VSUBS 0.014618f
C1501 VTAIL.n429 VSUBS 0.027203f
C1502 VTAIL.n430 VSUBS 0.027203f
C1503 VTAIL.n431 VSUBS 0.014618f
C1504 VTAIL.n432 VSUBS 0.015478f
C1505 VTAIL.n433 VSUBS 0.034551f
C1506 VTAIL.n434 VSUBS 0.034551f
C1507 VTAIL.n435 VSUBS 0.015478f
C1508 VTAIL.n436 VSUBS 0.014618f
C1509 VTAIL.n437 VSUBS 0.027203f
C1510 VTAIL.n438 VSUBS 0.027203f
C1511 VTAIL.n439 VSUBS 0.014618f
C1512 VTAIL.n440 VSUBS 0.015478f
C1513 VTAIL.n441 VSUBS 0.034551f
C1514 VTAIL.n442 VSUBS 0.087578f
C1515 VTAIL.n443 VSUBS 0.015478f
C1516 VTAIL.n444 VSUBS 0.014618f
C1517 VTAIL.n445 VSUBS 0.063994f
C1518 VTAIL.n446 VSUBS 0.044251f
C1519 VTAIL.n447 VSUBS 2.07205f
C1520 VDD2.n0 VSUBS 0.030919f
C1521 VDD2.n1 VSUBS 0.027093f
C1522 VDD2.n2 VSUBS 0.014558f
C1523 VDD2.n3 VSUBS 0.034411f
C1524 VDD2.n4 VSUBS 0.015415f
C1525 VDD2.n5 VSUBS 0.027093f
C1526 VDD2.n6 VSUBS 0.014558f
C1527 VDD2.n7 VSUBS 0.034411f
C1528 VDD2.n8 VSUBS 0.015415f
C1529 VDD2.n9 VSUBS 0.027093f
C1530 VDD2.n10 VSUBS 0.014558f
C1531 VDD2.n11 VSUBS 0.034411f
C1532 VDD2.n12 VSUBS 0.014987f
C1533 VDD2.n13 VSUBS 0.027093f
C1534 VDD2.n14 VSUBS 0.015415f
C1535 VDD2.n15 VSUBS 0.034411f
C1536 VDD2.n16 VSUBS 0.015415f
C1537 VDD2.n17 VSUBS 0.027093f
C1538 VDD2.n18 VSUBS 0.014558f
C1539 VDD2.n19 VSUBS 0.034411f
C1540 VDD2.n20 VSUBS 0.015415f
C1541 VDD2.n21 VSUBS 0.027093f
C1542 VDD2.n22 VSUBS 0.014558f
C1543 VDD2.n23 VSUBS 0.034411f
C1544 VDD2.n24 VSUBS 0.015415f
C1545 VDD2.n25 VSUBS 0.027093f
C1546 VDD2.n26 VSUBS 0.014558f
C1547 VDD2.n27 VSUBS 0.034411f
C1548 VDD2.n28 VSUBS 0.015415f
C1549 VDD2.n29 VSUBS 0.027093f
C1550 VDD2.n30 VSUBS 0.014558f
C1551 VDD2.n31 VSUBS 0.034411f
C1552 VDD2.n32 VSUBS 0.015415f
C1553 VDD2.n33 VSUBS 2.30922f
C1554 VDD2.n34 VSUBS 0.014558f
C1555 VDD2.t0 VSUBS 0.073984f
C1556 VDD2.n35 VSUBS 0.228619f
C1557 VDD2.n36 VSUBS 0.021891f
C1558 VDD2.n37 VSUBS 0.025808f
C1559 VDD2.n38 VSUBS 0.034411f
C1560 VDD2.n39 VSUBS 0.015415f
C1561 VDD2.n40 VSUBS 0.014558f
C1562 VDD2.n41 VSUBS 0.027093f
C1563 VDD2.n42 VSUBS 0.027093f
C1564 VDD2.n43 VSUBS 0.014558f
C1565 VDD2.n44 VSUBS 0.015415f
C1566 VDD2.n45 VSUBS 0.034411f
C1567 VDD2.n46 VSUBS 0.034411f
C1568 VDD2.n47 VSUBS 0.015415f
C1569 VDD2.n48 VSUBS 0.014558f
C1570 VDD2.n49 VSUBS 0.027093f
C1571 VDD2.n50 VSUBS 0.027093f
C1572 VDD2.n51 VSUBS 0.014558f
C1573 VDD2.n52 VSUBS 0.015415f
C1574 VDD2.n53 VSUBS 0.034411f
C1575 VDD2.n54 VSUBS 0.034411f
C1576 VDD2.n55 VSUBS 0.015415f
C1577 VDD2.n56 VSUBS 0.014558f
C1578 VDD2.n57 VSUBS 0.027093f
C1579 VDD2.n58 VSUBS 0.027093f
C1580 VDD2.n59 VSUBS 0.014558f
C1581 VDD2.n60 VSUBS 0.015415f
C1582 VDD2.n61 VSUBS 0.034411f
C1583 VDD2.n62 VSUBS 0.034411f
C1584 VDD2.n63 VSUBS 0.015415f
C1585 VDD2.n64 VSUBS 0.014558f
C1586 VDD2.n65 VSUBS 0.027093f
C1587 VDD2.n66 VSUBS 0.027093f
C1588 VDD2.n67 VSUBS 0.014558f
C1589 VDD2.n68 VSUBS 0.015415f
C1590 VDD2.n69 VSUBS 0.034411f
C1591 VDD2.n70 VSUBS 0.034411f
C1592 VDD2.n71 VSUBS 0.015415f
C1593 VDD2.n72 VSUBS 0.014558f
C1594 VDD2.n73 VSUBS 0.027093f
C1595 VDD2.n74 VSUBS 0.027093f
C1596 VDD2.n75 VSUBS 0.014558f
C1597 VDD2.n76 VSUBS 0.014558f
C1598 VDD2.n77 VSUBS 0.015415f
C1599 VDD2.n78 VSUBS 0.034411f
C1600 VDD2.n79 VSUBS 0.034411f
C1601 VDD2.n80 VSUBS 0.034411f
C1602 VDD2.n81 VSUBS 0.014987f
C1603 VDD2.n82 VSUBS 0.014558f
C1604 VDD2.n83 VSUBS 0.027093f
C1605 VDD2.n84 VSUBS 0.027093f
C1606 VDD2.n85 VSUBS 0.014558f
C1607 VDD2.n86 VSUBS 0.015415f
C1608 VDD2.n87 VSUBS 0.034411f
C1609 VDD2.n88 VSUBS 0.034411f
C1610 VDD2.n89 VSUBS 0.015415f
C1611 VDD2.n90 VSUBS 0.014558f
C1612 VDD2.n91 VSUBS 0.027093f
C1613 VDD2.n92 VSUBS 0.027093f
C1614 VDD2.n93 VSUBS 0.014558f
C1615 VDD2.n94 VSUBS 0.015415f
C1616 VDD2.n95 VSUBS 0.034411f
C1617 VDD2.n96 VSUBS 0.034411f
C1618 VDD2.n97 VSUBS 0.015415f
C1619 VDD2.n98 VSUBS 0.014558f
C1620 VDD2.n99 VSUBS 0.027093f
C1621 VDD2.n100 VSUBS 0.027093f
C1622 VDD2.n101 VSUBS 0.014558f
C1623 VDD2.n102 VSUBS 0.015415f
C1624 VDD2.n103 VSUBS 0.034411f
C1625 VDD2.n104 VSUBS 0.087222f
C1626 VDD2.n105 VSUBS 0.015415f
C1627 VDD2.n106 VSUBS 0.014558f
C1628 VDD2.n107 VSUBS 0.063734f
C1629 VDD2.n108 VSUBS 0.06511f
C1630 VDD2.t2 VSUBS 0.42198f
C1631 VDD2.t5 VSUBS 0.42198f
C1632 VDD2.n109 VSUBS 3.54747f
C1633 VDD2.n110 VSUBS 3.0514f
C1634 VDD2.n111 VSUBS 0.030919f
C1635 VDD2.n112 VSUBS 0.027093f
C1636 VDD2.n113 VSUBS 0.014558f
C1637 VDD2.n114 VSUBS 0.034411f
C1638 VDD2.n115 VSUBS 0.015415f
C1639 VDD2.n116 VSUBS 0.027093f
C1640 VDD2.n117 VSUBS 0.014558f
C1641 VDD2.n118 VSUBS 0.034411f
C1642 VDD2.n119 VSUBS 0.015415f
C1643 VDD2.n120 VSUBS 0.027093f
C1644 VDD2.n121 VSUBS 0.014558f
C1645 VDD2.n122 VSUBS 0.034411f
C1646 VDD2.n123 VSUBS 0.014987f
C1647 VDD2.n124 VSUBS 0.027093f
C1648 VDD2.n125 VSUBS 0.014987f
C1649 VDD2.n126 VSUBS 0.014558f
C1650 VDD2.n127 VSUBS 0.034411f
C1651 VDD2.n128 VSUBS 0.034411f
C1652 VDD2.n129 VSUBS 0.015415f
C1653 VDD2.n130 VSUBS 0.027093f
C1654 VDD2.n131 VSUBS 0.014558f
C1655 VDD2.n132 VSUBS 0.034411f
C1656 VDD2.n133 VSUBS 0.015415f
C1657 VDD2.n134 VSUBS 0.027093f
C1658 VDD2.n135 VSUBS 0.014558f
C1659 VDD2.n136 VSUBS 0.034411f
C1660 VDD2.n137 VSUBS 0.015415f
C1661 VDD2.n138 VSUBS 0.027093f
C1662 VDD2.n139 VSUBS 0.014558f
C1663 VDD2.n140 VSUBS 0.034411f
C1664 VDD2.n141 VSUBS 0.015415f
C1665 VDD2.n142 VSUBS 0.027093f
C1666 VDD2.n143 VSUBS 0.014558f
C1667 VDD2.n144 VSUBS 0.034411f
C1668 VDD2.n145 VSUBS 0.015415f
C1669 VDD2.n146 VSUBS 2.30922f
C1670 VDD2.n147 VSUBS 0.014558f
C1671 VDD2.t4 VSUBS 0.073984f
C1672 VDD2.n148 VSUBS 0.228619f
C1673 VDD2.n149 VSUBS 0.021891f
C1674 VDD2.n150 VSUBS 0.025808f
C1675 VDD2.n151 VSUBS 0.034411f
C1676 VDD2.n152 VSUBS 0.015415f
C1677 VDD2.n153 VSUBS 0.014558f
C1678 VDD2.n154 VSUBS 0.027093f
C1679 VDD2.n155 VSUBS 0.027093f
C1680 VDD2.n156 VSUBS 0.014558f
C1681 VDD2.n157 VSUBS 0.015415f
C1682 VDD2.n158 VSUBS 0.034411f
C1683 VDD2.n159 VSUBS 0.034411f
C1684 VDD2.n160 VSUBS 0.015415f
C1685 VDD2.n161 VSUBS 0.014558f
C1686 VDD2.n162 VSUBS 0.027093f
C1687 VDD2.n163 VSUBS 0.027093f
C1688 VDD2.n164 VSUBS 0.014558f
C1689 VDD2.n165 VSUBS 0.015415f
C1690 VDD2.n166 VSUBS 0.034411f
C1691 VDD2.n167 VSUBS 0.034411f
C1692 VDD2.n168 VSUBS 0.015415f
C1693 VDD2.n169 VSUBS 0.014558f
C1694 VDD2.n170 VSUBS 0.027093f
C1695 VDD2.n171 VSUBS 0.027093f
C1696 VDD2.n172 VSUBS 0.014558f
C1697 VDD2.n173 VSUBS 0.015415f
C1698 VDD2.n174 VSUBS 0.034411f
C1699 VDD2.n175 VSUBS 0.034411f
C1700 VDD2.n176 VSUBS 0.015415f
C1701 VDD2.n177 VSUBS 0.014558f
C1702 VDD2.n178 VSUBS 0.027093f
C1703 VDD2.n179 VSUBS 0.027093f
C1704 VDD2.n180 VSUBS 0.014558f
C1705 VDD2.n181 VSUBS 0.015415f
C1706 VDD2.n182 VSUBS 0.034411f
C1707 VDD2.n183 VSUBS 0.034411f
C1708 VDD2.n184 VSUBS 0.015415f
C1709 VDD2.n185 VSUBS 0.014558f
C1710 VDD2.n186 VSUBS 0.027093f
C1711 VDD2.n187 VSUBS 0.027093f
C1712 VDD2.n188 VSUBS 0.014558f
C1713 VDD2.n189 VSUBS 0.015415f
C1714 VDD2.n190 VSUBS 0.034411f
C1715 VDD2.n191 VSUBS 0.034411f
C1716 VDD2.n192 VSUBS 0.015415f
C1717 VDD2.n193 VSUBS 0.014558f
C1718 VDD2.n194 VSUBS 0.027093f
C1719 VDD2.n195 VSUBS 0.027093f
C1720 VDD2.n196 VSUBS 0.014558f
C1721 VDD2.n197 VSUBS 0.015415f
C1722 VDD2.n198 VSUBS 0.034411f
C1723 VDD2.n199 VSUBS 0.034411f
C1724 VDD2.n200 VSUBS 0.015415f
C1725 VDD2.n201 VSUBS 0.014558f
C1726 VDD2.n202 VSUBS 0.027093f
C1727 VDD2.n203 VSUBS 0.027093f
C1728 VDD2.n204 VSUBS 0.014558f
C1729 VDD2.n205 VSUBS 0.015415f
C1730 VDD2.n206 VSUBS 0.034411f
C1731 VDD2.n207 VSUBS 0.034411f
C1732 VDD2.n208 VSUBS 0.015415f
C1733 VDD2.n209 VSUBS 0.014558f
C1734 VDD2.n210 VSUBS 0.027093f
C1735 VDD2.n211 VSUBS 0.027093f
C1736 VDD2.n212 VSUBS 0.014558f
C1737 VDD2.n213 VSUBS 0.015415f
C1738 VDD2.n214 VSUBS 0.034411f
C1739 VDD2.n215 VSUBS 0.087222f
C1740 VDD2.n216 VSUBS 0.015415f
C1741 VDD2.n217 VSUBS 0.014558f
C1742 VDD2.n218 VSUBS 0.063734f
C1743 VDD2.n219 VSUBS 0.062769f
C1744 VDD2.n220 VSUBS 2.98575f
C1745 VDD2.t3 VSUBS 0.42198f
C1746 VDD2.t1 VSUBS 0.42198f
C1747 VDD2.n221 VSUBS 3.54743f
C1748 VN.n0 VSUBS 0.239919f
C1749 VN.t0 VSUBS 2.63276f
C1750 VN.t4 VSUBS 2.75712f
C1751 VN.n1 VSUBS 0.987751f
C1752 VN.n2 VSUBS 1.00351f
C1753 VN.n3 VSUBS 0.058803f
C1754 VN.t5 VSUBS 2.70703f
C1755 VN.n4 VSUBS 1.00844f
C1756 VN.n5 VSUBS 0.03983f
C1757 VN.n6 VSUBS 0.239919f
C1758 VN.t2 VSUBS 2.63276f
C1759 VN.t1 VSUBS 2.75712f
C1760 VN.n7 VSUBS 0.987751f
C1761 VN.n8 VSUBS 1.00351f
C1762 VN.n9 VSUBS 0.058803f
C1763 VN.t3 VSUBS 2.70703f
C1764 VN.n10 VSUBS 1.00844f
C1765 VN.n11 VSUBS 2.28245f
.ends

