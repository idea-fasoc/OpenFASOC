* NGSPICE file created from diff_pair_sample_1754.ext - technology: sky130A

.subckt diff_pair_sample_1754 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t15 B.t1 sky130_fd_pr__nfet_01v8 ad=0.91245 pd=5.86 as=0.91245 ps=5.86 w=5.53 l=1.16
X1 VTAIL.t6 VP.t0 VDD1.t7 B.t20 sky130_fd_pr__nfet_01v8 ad=0.91245 pd=5.86 as=0.91245 ps=5.86 w=5.53 l=1.16
X2 VDD2.t6 VN.t1 VTAIL.t10 B.t21 sky130_fd_pr__nfet_01v8 ad=0.91245 pd=5.86 as=0.91245 ps=5.86 w=5.53 l=1.16
X3 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=2.1567 pd=11.84 as=0 ps=0 w=5.53 l=1.16
X4 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=2.1567 pd=11.84 as=0 ps=0 w=5.53 l=1.16
X5 VTAIL.t4 VP.t1 VDD1.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=0.91245 pd=5.86 as=0.91245 ps=5.86 w=5.53 l=1.16
X6 VDD1.t5 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.91245 pd=5.86 as=0.91245 ps=5.86 w=5.53 l=1.16
X7 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.1567 pd=11.84 as=0 ps=0 w=5.53 l=1.16
X8 VTAIL.t13 VN.t2 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=0.91245 pd=5.86 as=0.91245 ps=5.86 w=5.53 l=1.16
X9 VTAIL.t2 VP.t3 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1567 pd=11.84 as=0.91245 ps=5.86 w=5.53 l=1.16
X10 VTAIL.t8 VN.t3 VDD2.t4 B.t20 sky130_fd_pr__nfet_01v8 ad=0.91245 pd=5.86 as=0.91245 ps=5.86 w=5.53 l=1.16
X11 VDD2.t3 VN.t4 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=0.91245 pd=5.86 as=2.1567 ps=11.84 w=5.53 l=1.16
X12 VDD1.t3 VP.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.91245 pd=5.86 as=2.1567 ps=11.84 w=5.53 l=1.16
X13 VTAIL.t11 VN.t5 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1567 pd=11.84 as=0.91245 ps=5.86 w=5.53 l=1.16
X14 VDD1.t2 VP.t5 VTAIL.t7 B.t21 sky130_fd_pr__nfet_01v8 ad=0.91245 pd=5.86 as=0.91245 ps=5.86 w=5.53 l=1.16
X15 VDD2.t1 VN.t6 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=0.91245 pd=5.86 as=2.1567 ps=11.84 w=5.53 l=1.16
X16 VDD1.t1 VP.t6 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.91245 pd=5.86 as=2.1567 ps=11.84 w=5.53 l=1.16
X17 VTAIL.t0 VP.t7 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1567 pd=11.84 as=0.91245 ps=5.86 w=5.53 l=1.16
X18 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.1567 pd=11.84 as=0 ps=0 w=5.53 l=1.16
X19 VTAIL.t14 VN.t7 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1567 pd=11.84 as=0.91245 ps=5.86 w=5.53 l=1.16
R0 VN.n16 VN.n15 174.268
R1 VN.n33 VN.n32 174.268
R2 VN.n31 VN.n17 161.3
R3 VN.n30 VN.n29 161.3
R4 VN.n28 VN.n18 161.3
R5 VN.n27 VN.n26 161.3
R6 VN.n25 VN.n19 161.3
R7 VN.n24 VN.n23 161.3
R8 VN.n14 VN.n0 161.3
R9 VN.n13 VN.n12 161.3
R10 VN.n11 VN.n1 161.3
R11 VN.n10 VN.n9 161.3
R12 VN.n7 VN.n2 161.3
R13 VN.n6 VN.n5 161.3
R14 VN.n4 VN.t5 144.495
R15 VN.n22 VN.t4 144.495
R16 VN.n3 VN.t0 114.891
R17 VN.n8 VN.t3 114.891
R18 VN.n15 VN.t6 114.891
R19 VN.n21 VN.t2 114.891
R20 VN.n20 VN.t1 114.891
R21 VN.n32 VN.t7 114.891
R22 VN.n4 VN.n3 51.7518
R23 VN.n22 VN.n21 51.7518
R24 VN.n13 VN.n1 41.4647
R25 VN.n30 VN.n18 41.4647
R26 VN.n7 VN.n6 40.4934
R27 VN.n9 VN.n7 40.4934
R28 VN.n25 VN.n24 40.4934
R29 VN.n26 VN.n25 40.4934
R30 VN.n14 VN.n13 39.5221
R31 VN.n31 VN.n30 39.5221
R32 VN VN.n33 39.5024
R33 VN.n23 VN.n22 27.1667
R34 VN.n5 VN.n4 27.1667
R35 VN.n8 VN.n1 12.4787
R36 VN.n20 VN.n18 12.4787
R37 VN.n6 VN.n3 11.9893
R38 VN.n9 VN.n8 11.9893
R39 VN.n24 VN.n21 11.9893
R40 VN.n26 VN.n20 11.9893
R41 VN.n15 VN.n14 11.5
R42 VN.n32 VN.n31 11.5
R43 VN.n33 VN.n17 0.189894
R44 VN.n29 VN.n17 0.189894
R45 VN.n29 VN.n28 0.189894
R46 VN.n28 VN.n27 0.189894
R47 VN.n27 VN.n19 0.189894
R48 VN.n23 VN.n19 0.189894
R49 VN.n5 VN.n2 0.189894
R50 VN.n10 VN.n2 0.189894
R51 VN.n11 VN.n10 0.189894
R52 VN.n12 VN.n11 0.189894
R53 VN.n12 VN.n0 0.189894
R54 VN.n16 VN.n0 0.189894
R55 VN VN.n16 0.0516364
R56 VTAIL.n11 VTAIL.t2 52.6384
R57 VTAIL.n10 VTAIL.t12 52.6384
R58 VTAIL.n7 VTAIL.t14 52.6384
R59 VTAIL.n15 VTAIL.t9 52.6382
R60 VTAIL.n2 VTAIL.t11 52.6382
R61 VTAIL.n3 VTAIL.t5 52.6382
R62 VTAIL.n6 VTAIL.t0 52.6382
R63 VTAIL.n14 VTAIL.t3 52.6382
R64 VTAIL.n13 VTAIL.n12 49.0579
R65 VTAIL.n9 VTAIL.n8 49.0579
R66 VTAIL.n1 VTAIL.n0 49.0577
R67 VTAIL.n5 VTAIL.n4 49.0577
R68 VTAIL.n15 VTAIL.n14 18.4186
R69 VTAIL.n7 VTAIL.n6 18.4186
R70 VTAIL.n0 VTAIL.t15 3.58097
R71 VTAIL.n0 VTAIL.t8 3.58097
R72 VTAIL.n4 VTAIL.t7 3.58097
R73 VTAIL.n4 VTAIL.t4 3.58097
R74 VTAIL.n12 VTAIL.t1 3.58097
R75 VTAIL.n12 VTAIL.t6 3.58097
R76 VTAIL.n8 VTAIL.t10 3.58097
R77 VTAIL.n8 VTAIL.t13 3.58097
R78 VTAIL.n9 VTAIL.n7 1.28498
R79 VTAIL.n10 VTAIL.n9 1.28498
R80 VTAIL.n13 VTAIL.n11 1.28498
R81 VTAIL.n14 VTAIL.n13 1.28498
R82 VTAIL.n6 VTAIL.n5 1.28498
R83 VTAIL.n5 VTAIL.n3 1.28498
R84 VTAIL.n2 VTAIL.n1 1.28498
R85 VTAIL VTAIL.n15 1.22679
R86 VTAIL.n11 VTAIL.n10 0.470328
R87 VTAIL.n3 VTAIL.n2 0.470328
R88 VTAIL VTAIL.n1 0.0586897
R89 VDD2.n2 VDD2.n1 66.3234
R90 VDD2.n2 VDD2.n0 66.3234
R91 VDD2 VDD2.n5 66.3206
R92 VDD2.n4 VDD2.n3 65.7367
R93 VDD2.n4 VDD2.n2 34.2627
R94 VDD2.n5 VDD2.t5 3.58097
R95 VDD2.n5 VDD2.t3 3.58097
R96 VDD2.n3 VDD2.t0 3.58097
R97 VDD2.n3 VDD2.t6 3.58097
R98 VDD2.n1 VDD2.t4 3.58097
R99 VDD2.n1 VDD2.t1 3.58097
R100 VDD2.n0 VDD2.t2 3.58097
R101 VDD2.n0 VDD2.t7 3.58097
R102 VDD2 VDD2.n4 0.700931
R103 B.n420 B.n419 585
R104 B.n420 B.n57 585
R105 B.n423 B.n422 585
R106 B.n424 B.n89 585
R107 B.n426 B.n425 585
R108 B.n428 B.n88 585
R109 B.n431 B.n430 585
R110 B.n432 B.n87 585
R111 B.n434 B.n433 585
R112 B.n436 B.n86 585
R113 B.n439 B.n438 585
R114 B.n440 B.n85 585
R115 B.n442 B.n441 585
R116 B.n444 B.n84 585
R117 B.n447 B.n446 585
R118 B.n448 B.n83 585
R119 B.n450 B.n449 585
R120 B.n452 B.n82 585
R121 B.n455 B.n454 585
R122 B.n456 B.n81 585
R123 B.n458 B.n457 585
R124 B.n460 B.n80 585
R125 B.n463 B.n462 585
R126 B.n464 B.n77 585
R127 B.n467 B.n466 585
R128 B.n469 B.n76 585
R129 B.n472 B.n471 585
R130 B.n473 B.n75 585
R131 B.n475 B.n474 585
R132 B.n477 B.n74 585
R133 B.n480 B.n479 585
R134 B.n481 B.n70 585
R135 B.n483 B.n482 585
R136 B.n485 B.n69 585
R137 B.n488 B.n487 585
R138 B.n489 B.n68 585
R139 B.n491 B.n490 585
R140 B.n493 B.n67 585
R141 B.n496 B.n495 585
R142 B.n497 B.n66 585
R143 B.n499 B.n498 585
R144 B.n501 B.n65 585
R145 B.n504 B.n503 585
R146 B.n505 B.n64 585
R147 B.n507 B.n506 585
R148 B.n509 B.n63 585
R149 B.n512 B.n511 585
R150 B.n513 B.n62 585
R151 B.n515 B.n514 585
R152 B.n517 B.n61 585
R153 B.n520 B.n519 585
R154 B.n521 B.n60 585
R155 B.n523 B.n522 585
R156 B.n525 B.n59 585
R157 B.n528 B.n527 585
R158 B.n529 B.n58 585
R159 B.n418 B.n56 585
R160 B.n532 B.n56 585
R161 B.n417 B.n55 585
R162 B.n533 B.n55 585
R163 B.n416 B.n54 585
R164 B.n534 B.n54 585
R165 B.n415 B.n414 585
R166 B.n414 B.n50 585
R167 B.n413 B.n49 585
R168 B.n540 B.n49 585
R169 B.n412 B.n48 585
R170 B.n541 B.n48 585
R171 B.n411 B.n47 585
R172 B.n542 B.n47 585
R173 B.n410 B.n409 585
R174 B.n409 B.n43 585
R175 B.n408 B.n42 585
R176 B.n548 B.n42 585
R177 B.n407 B.n41 585
R178 B.n549 B.n41 585
R179 B.n406 B.n40 585
R180 B.n550 B.n40 585
R181 B.n405 B.n404 585
R182 B.n404 B.n36 585
R183 B.n403 B.n35 585
R184 B.n556 B.n35 585
R185 B.n402 B.n34 585
R186 B.n557 B.n34 585
R187 B.n401 B.n33 585
R188 B.n558 B.n33 585
R189 B.n400 B.n399 585
R190 B.n399 B.n29 585
R191 B.n398 B.n28 585
R192 B.n564 B.n28 585
R193 B.n397 B.n27 585
R194 B.n565 B.n27 585
R195 B.n396 B.n26 585
R196 B.n566 B.n26 585
R197 B.n395 B.n394 585
R198 B.n394 B.n22 585
R199 B.n393 B.n21 585
R200 B.n572 B.n21 585
R201 B.n392 B.n20 585
R202 B.n573 B.n20 585
R203 B.n391 B.n19 585
R204 B.n574 B.n19 585
R205 B.n390 B.n389 585
R206 B.n389 B.n15 585
R207 B.n388 B.n14 585
R208 B.n580 B.n14 585
R209 B.n387 B.n13 585
R210 B.n581 B.n13 585
R211 B.n386 B.n12 585
R212 B.n582 B.n12 585
R213 B.n385 B.n384 585
R214 B.n384 B.n8 585
R215 B.n383 B.n7 585
R216 B.n588 B.n7 585
R217 B.n382 B.n6 585
R218 B.n589 B.n6 585
R219 B.n381 B.n5 585
R220 B.n590 B.n5 585
R221 B.n380 B.n379 585
R222 B.n379 B.n4 585
R223 B.n378 B.n90 585
R224 B.n378 B.n377 585
R225 B.n368 B.n91 585
R226 B.n92 B.n91 585
R227 B.n370 B.n369 585
R228 B.n371 B.n370 585
R229 B.n367 B.n97 585
R230 B.n97 B.n96 585
R231 B.n366 B.n365 585
R232 B.n365 B.n364 585
R233 B.n99 B.n98 585
R234 B.n100 B.n99 585
R235 B.n357 B.n356 585
R236 B.n358 B.n357 585
R237 B.n355 B.n104 585
R238 B.n108 B.n104 585
R239 B.n354 B.n353 585
R240 B.n353 B.n352 585
R241 B.n106 B.n105 585
R242 B.n107 B.n106 585
R243 B.n345 B.n344 585
R244 B.n346 B.n345 585
R245 B.n343 B.n112 585
R246 B.n116 B.n112 585
R247 B.n342 B.n341 585
R248 B.n341 B.n340 585
R249 B.n114 B.n113 585
R250 B.n115 B.n114 585
R251 B.n333 B.n332 585
R252 B.n334 B.n333 585
R253 B.n331 B.n120 585
R254 B.n124 B.n120 585
R255 B.n330 B.n329 585
R256 B.n329 B.n328 585
R257 B.n122 B.n121 585
R258 B.n123 B.n122 585
R259 B.n321 B.n320 585
R260 B.n322 B.n321 585
R261 B.n319 B.n129 585
R262 B.n129 B.n128 585
R263 B.n318 B.n317 585
R264 B.n317 B.n316 585
R265 B.n131 B.n130 585
R266 B.n132 B.n131 585
R267 B.n309 B.n308 585
R268 B.n310 B.n309 585
R269 B.n307 B.n136 585
R270 B.n140 B.n136 585
R271 B.n306 B.n305 585
R272 B.n305 B.n304 585
R273 B.n138 B.n137 585
R274 B.n139 B.n138 585
R275 B.n297 B.n296 585
R276 B.n298 B.n297 585
R277 B.n295 B.n145 585
R278 B.n145 B.n144 585
R279 B.n294 B.n293 585
R280 B.n293 B.n292 585
R281 B.n289 B.n149 585
R282 B.n288 B.n287 585
R283 B.n285 B.n150 585
R284 B.n285 B.n148 585
R285 B.n284 B.n283 585
R286 B.n282 B.n281 585
R287 B.n280 B.n152 585
R288 B.n278 B.n277 585
R289 B.n276 B.n153 585
R290 B.n275 B.n274 585
R291 B.n272 B.n154 585
R292 B.n270 B.n269 585
R293 B.n268 B.n155 585
R294 B.n267 B.n266 585
R295 B.n264 B.n156 585
R296 B.n262 B.n261 585
R297 B.n260 B.n157 585
R298 B.n259 B.n258 585
R299 B.n256 B.n158 585
R300 B.n254 B.n253 585
R301 B.n252 B.n159 585
R302 B.n251 B.n250 585
R303 B.n248 B.n160 585
R304 B.n246 B.n245 585
R305 B.n243 B.n161 585
R306 B.n242 B.n241 585
R307 B.n239 B.n164 585
R308 B.n237 B.n236 585
R309 B.n235 B.n165 585
R310 B.n234 B.n233 585
R311 B.n231 B.n166 585
R312 B.n229 B.n228 585
R313 B.n227 B.n167 585
R314 B.n225 B.n224 585
R315 B.n222 B.n170 585
R316 B.n220 B.n219 585
R317 B.n218 B.n171 585
R318 B.n217 B.n216 585
R319 B.n214 B.n172 585
R320 B.n212 B.n211 585
R321 B.n210 B.n173 585
R322 B.n209 B.n208 585
R323 B.n206 B.n174 585
R324 B.n204 B.n203 585
R325 B.n202 B.n175 585
R326 B.n201 B.n200 585
R327 B.n198 B.n176 585
R328 B.n196 B.n195 585
R329 B.n194 B.n177 585
R330 B.n193 B.n192 585
R331 B.n190 B.n178 585
R332 B.n188 B.n187 585
R333 B.n186 B.n179 585
R334 B.n185 B.n184 585
R335 B.n182 B.n180 585
R336 B.n147 B.n146 585
R337 B.n291 B.n290 585
R338 B.n292 B.n291 585
R339 B.n143 B.n142 585
R340 B.n144 B.n143 585
R341 B.n300 B.n299 585
R342 B.n299 B.n298 585
R343 B.n301 B.n141 585
R344 B.n141 B.n139 585
R345 B.n303 B.n302 585
R346 B.n304 B.n303 585
R347 B.n135 B.n134 585
R348 B.n140 B.n135 585
R349 B.n312 B.n311 585
R350 B.n311 B.n310 585
R351 B.n313 B.n133 585
R352 B.n133 B.n132 585
R353 B.n315 B.n314 585
R354 B.n316 B.n315 585
R355 B.n127 B.n126 585
R356 B.n128 B.n127 585
R357 B.n324 B.n323 585
R358 B.n323 B.n322 585
R359 B.n325 B.n125 585
R360 B.n125 B.n123 585
R361 B.n327 B.n326 585
R362 B.n328 B.n327 585
R363 B.n119 B.n118 585
R364 B.n124 B.n119 585
R365 B.n336 B.n335 585
R366 B.n335 B.n334 585
R367 B.n337 B.n117 585
R368 B.n117 B.n115 585
R369 B.n339 B.n338 585
R370 B.n340 B.n339 585
R371 B.n111 B.n110 585
R372 B.n116 B.n111 585
R373 B.n348 B.n347 585
R374 B.n347 B.n346 585
R375 B.n349 B.n109 585
R376 B.n109 B.n107 585
R377 B.n351 B.n350 585
R378 B.n352 B.n351 585
R379 B.n103 B.n102 585
R380 B.n108 B.n103 585
R381 B.n360 B.n359 585
R382 B.n359 B.n358 585
R383 B.n361 B.n101 585
R384 B.n101 B.n100 585
R385 B.n363 B.n362 585
R386 B.n364 B.n363 585
R387 B.n95 B.n94 585
R388 B.n96 B.n95 585
R389 B.n373 B.n372 585
R390 B.n372 B.n371 585
R391 B.n374 B.n93 585
R392 B.n93 B.n92 585
R393 B.n376 B.n375 585
R394 B.n377 B.n376 585
R395 B.n2 B.n0 585
R396 B.n4 B.n2 585
R397 B.n3 B.n1 585
R398 B.n589 B.n3 585
R399 B.n587 B.n586 585
R400 B.n588 B.n587 585
R401 B.n585 B.n9 585
R402 B.n9 B.n8 585
R403 B.n584 B.n583 585
R404 B.n583 B.n582 585
R405 B.n11 B.n10 585
R406 B.n581 B.n11 585
R407 B.n579 B.n578 585
R408 B.n580 B.n579 585
R409 B.n577 B.n16 585
R410 B.n16 B.n15 585
R411 B.n576 B.n575 585
R412 B.n575 B.n574 585
R413 B.n18 B.n17 585
R414 B.n573 B.n18 585
R415 B.n571 B.n570 585
R416 B.n572 B.n571 585
R417 B.n569 B.n23 585
R418 B.n23 B.n22 585
R419 B.n568 B.n567 585
R420 B.n567 B.n566 585
R421 B.n25 B.n24 585
R422 B.n565 B.n25 585
R423 B.n563 B.n562 585
R424 B.n564 B.n563 585
R425 B.n561 B.n30 585
R426 B.n30 B.n29 585
R427 B.n560 B.n559 585
R428 B.n559 B.n558 585
R429 B.n32 B.n31 585
R430 B.n557 B.n32 585
R431 B.n555 B.n554 585
R432 B.n556 B.n555 585
R433 B.n553 B.n37 585
R434 B.n37 B.n36 585
R435 B.n552 B.n551 585
R436 B.n551 B.n550 585
R437 B.n39 B.n38 585
R438 B.n549 B.n39 585
R439 B.n547 B.n546 585
R440 B.n548 B.n547 585
R441 B.n545 B.n44 585
R442 B.n44 B.n43 585
R443 B.n544 B.n543 585
R444 B.n543 B.n542 585
R445 B.n46 B.n45 585
R446 B.n541 B.n46 585
R447 B.n539 B.n538 585
R448 B.n540 B.n539 585
R449 B.n537 B.n51 585
R450 B.n51 B.n50 585
R451 B.n536 B.n535 585
R452 B.n535 B.n534 585
R453 B.n53 B.n52 585
R454 B.n533 B.n53 585
R455 B.n531 B.n530 585
R456 B.n532 B.n531 585
R457 B.n592 B.n591 585
R458 B.n591 B.n590 585
R459 B.n291 B.n149 482.89
R460 B.n531 B.n58 482.89
R461 B.n293 B.n147 482.89
R462 B.n420 B.n56 482.89
R463 B.n168 B.t14 318.793
R464 B.n162 B.t10 318.793
R465 B.n71 B.t6 318.793
R466 B.n78 B.t17 318.793
R467 B.n421 B.n57 256.663
R468 B.n427 B.n57 256.663
R469 B.n429 B.n57 256.663
R470 B.n435 B.n57 256.663
R471 B.n437 B.n57 256.663
R472 B.n443 B.n57 256.663
R473 B.n445 B.n57 256.663
R474 B.n451 B.n57 256.663
R475 B.n453 B.n57 256.663
R476 B.n459 B.n57 256.663
R477 B.n461 B.n57 256.663
R478 B.n468 B.n57 256.663
R479 B.n470 B.n57 256.663
R480 B.n476 B.n57 256.663
R481 B.n478 B.n57 256.663
R482 B.n484 B.n57 256.663
R483 B.n486 B.n57 256.663
R484 B.n492 B.n57 256.663
R485 B.n494 B.n57 256.663
R486 B.n500 B.n57 256.663
R487 B.n502 B.n57 256.663
R488 B.n508 B.n57 256.663
R489 B.n510 B.n57 256.663
R490 B.n516 B.n57 256.663
R491 B.n518 B.n57 256.663
R492 B.n524 B.n57 256.663
R493 B.n526 B.n57 256.663
R494 B.n286 B.n148 256.663
R495 B.n151 B.n148 256.663
R496 B.n279 B.n148 256.663
R497 B.n273 B.n148 256.663
R498 B.n271 B.n148 256.663
R499 B.n265 B.n148 256.663
R500 B.n263 B.n148 256.663
R501 B.n257 B.n148 256.663
R502 B.n255 B.n148 256.663
R503 B.n249 B.n148 256.663
R504 B.n247 B.n148 256.663
R505 B.n240 B.n148 256.663
R506 B.n238 B.n148 256.663
R507 B.n232 B.n148 256.663
R508 B.n230 B.n148 256.663
R509 B.n223 B.n148 256.663
R510 B.n221 B.n148 256.663
R511 B.n215 B.n148 256.663
R512 B.n213 B.n148 256.663
R513 B.n207 B.n148 256.663
R514 B.n205 B.n148 256.663
R515 B.n199 B.n148 256.663
R516 B.n197 B.n148 256.663
R517 B.n191 B.n148 256.663
R518 B.n189 B.n148 256.663
R519 B.n183 B.n148 256.663
R520 B.n181 B.n148 256.663
R521 B.n291 B.n143 163.367
R522 B.n299 B.n143 163.367
R523 B.n299 B.n141 163.367
R524 B.n303 B.n141 163.367
R525 B.n303 B.n135 163.367
R526 B.n311 B.n135 163.367
R527 B.n311 B.n133 163.367
R528 B.n315 B.n133 163.367
R529 B.n315 B.n127 163.367
R530 B.n323 B.n127 163.367
R531 B.n323 B.n125 163.367
R532 B.n327 B.n125 163.367
R533 B.n327 B.n119 163.367
R534 B.n335 B.n119 163.367
R535 B.n335 B.n117 163.367
R536 B.n339 B.n117 163.367
R537 B.n339 B.n111 163.367
R538 B.n347 B.n111 163.367
R539 B.n347 B.n109 163.367
R540 B.n351 B.n109 163.367
R541 B.n351 B.n103 163.367
R542 B.n359 B.n103 163.367
R543 B.n359 B.n101 163.367
R544 B.n363 B.n101 163.367
R545 B.n363 B.n95 163.367
R546 B.n372 B.n95 163.367
R547 B.n372 B.n93 163.367
R548 B.n376 B.n93 163.367
R549 B.n376 B.n2 163.367
R550 B.n591 B.n2 163.367
R551 B.n591 B.n3 163.367
R552 B.n587 B.n3 163.367
R553 B.n587 B.n9 163.367
R554 B.n583 B.n9 163.367
R555 B.n583 B.n11 163.367
R556 B.n579 B.n11 163.367
R557 B.n579 B.n16 163.367
R558 B.n575 B.n16 163.367
R559 B.n575 B.n18 163.367
R560 B.n571 B.n18 163.367
R561 B.n571 B.n23 163.367
R562 B.n567 B.n23 163.367
R563 B.n567 B.n25 163.367
R564 B.n563 B.n25 163.367
R565 B.n563 B.n30 163.367
R566 B.n559 B.n30 163.367
R567 B.n559 B.n32 163.367
R568 B.n555 B.n32 163.367
R569 B.n555 B.n37 163.367
R570 B.n551 B.n37 163.367
R571 B.n551 B.n39 163.367
R572 B.n547 B.n39 163.367
R573 B.n547 B.n44 163.367
R574 B.n543 B.n44 163.367
R575 B.n543 B.n46 163.367
R576 B.n539 B.n46 163.367
R577 B.n539 B.n51 163.367
R578 B.n535 B.n51 163.367
R579 B.n535 B.n53 163.367
R580 B.n531 B.n53 163.367
R581 B.n287 B.n285 163.367
R582 B.n285 B.n284 163.367
R583 B.n281 B.n280 163.367
R584 B.n278 B.n153 163.367
R585 B.n274 B.n272 163.367
R586 B.n270 B.n155 163.367
R587 B.n266 B.n264 163.367
R588 B.n262 B.n157 163.367
R589 B.n258 B.n256 163.367
R590 B.n254 B.n159 163.367
R591 B.n250 B.n248 163.367
R592 B.n246 B.n161 163.367
R593 B.n241 B.n239 163.367
R594 B.n237 B.n165 163.367
R595 B.n233 B.n231 163.367
R596 B.n229 B.n167 163.367
R597 B.n224 B.n222 163.367
R598 B.n220 B.n171 163.367
R599 B.n216 B.n214 163.367
R600 B.n212 B.n173 163.367
R601 B.n208 B.n206 163.367
R602 B.n204 B.n175 163.367
R603 B.n200 B.n198 163.367
R604 B.n196 B.n177 163.367
R605 B.n192 B.n190 163.367
R606 B.n188 B.n179 163.367
R607 B.n184 B.n182 163.367
R608 B.n293 B.n145 163.367
R609 B.n297 B.n145 163.367
R610 B.n297 B.n138 163.367
R611 B.n305 B.n138 163.367
R612 B.n305 B.n136 163.367
R613 B.n309 B.n136 163.367
R614 B.n309 B.n131 163.367
R615 B.n317 B.n131 163.367
R616 B.n317 B.n129 163.367
R617 B.n321 B.n129 163.367
R618 B.n321 B.n122 163.367
R619 B.n329 B.n122 163.367
R620 B.n329 B.n120 163.367
R621 B.n333 B.n120 163.367
R622 B.n333 B.n114 163.367
R623 B.n341 B.n114 163.367
R624 B.n341 B.n112 163.367
R625 B.n345 B.n112 163.367
R626 B.n345 B.n106 163.367
R627 B.n353 B.n106 163.367
R628 B.n353 B.n104 163.367
R629 B.n357 B.n104 163.367
R630 B.n357 B.n99 163.367
R631 B.n365 B.n99 163.367
R632 B.n365 B.n97 163.367
R633 B.n370 B.n97 163.367
R634 B.n370 B.n91 163.367
R635 B.n378 B.n91 163.367
R636 B.n379 B.n378 163.367
R637 B.n379 B.n5 163.367
R638 B.n6 B.n5 163.367
R639 B.n7 B.n6 163.367
R640 B.n384 B.n7 163.367
R641 B.n384 B.n12 163.367
R642 B.n13 B.n12 163.367
R643 B.n14 B.n13 163.367
R644 B.n389 B.n14 163.367
R645 B.n389 B.n19 163.367
R646 B.n20 B.n19 163.367
R647 B.n21 B.n20 163.367
R648 B.n394 B.n21 163.367
R649 B.n394 B.n26 163.367
R650 B.n27 B.n26 163.367
R651 B.n28 B.n27 163.367
R652 B.n399 B.n28 163.367
R653 B.n399 B.n33 163.367
R654 B.n34 B.n33 163.367
R655 B.n35 B.n34 163.367
R656 B.n404 B.n35 163.367
R657 B.n404 B.n40 163.367
R658 B.n41 B.n40 163.367
R659 B.n42 B.n41 163.367
R660 B.n409 B.n42 163.367
R661 B.n409 B.n47 163.367
R662 B.n48 B.n47 163.367
R663 B.n49 B.n48 163.367
R664 B.n414 B.n49 163.367
R665 B.n414 B.n54 163.367
R666 B.n55 B.n54 163.367
R667 B.n56 B.n55 163.367
R668 B.n527 B.n525 163.367
R669 B.n523 B.n60 163.367
R670 B.n519 B.n517 163.367
R671 B.n515 B.n62 163.367
R672 B.n511 B.n509 163.367
R673 B.n507 B.n64 163.367
R674 B.n503 B.n501 163.367
R675 B.n499 B.n66 163.367
R676 B.n495 B.n493 163.367
R677 B.n491 B.n68 163.367
R678 B.n487 B.n485 163.367
R679 B.n483 B.n70 163.367
R680 B.n479 B.n477 163.367
R681 B.n475 B.n75 163.367
R682 B.n471 B.n469 163.367
R683 B.n467 B.n77 163.367
R684 B.n462 B.n460 163.367
R685 B.n458 B.n81 163.367
R686 B.n454 B.n452 163.367
R687 B.n450 B.n83 163.367
R688 B.n446 B.n444 163.367
R689 B.n442 B.n85 163.367
R690 B.n438 B.n436 163.367
R691 B.n434 B.n87 163.367
R692 B.n430 B.n428 163.367
R693 B.n426 B.n89 163.367
R694 B.n422 B.n420 163.367
R695 B.n292 B.n148 127.257
R696 B.n532 B.n57 127.257
R697 B.n168 B.t16 100.388
R698 B.n78 B.t18 100.388
R699 B.n162 B.t13 100.382
R700 B.n71 B.t8 100.382
R701 B.n286 B.n149 71.676
R702 B.n284 B.n151 71.676
R703 B.n280 B.n279 71.676
R704 B.n273 B.n153 71.676
R705 B.n272 B.n271 71.676
R706 B.n265 B.n155 71.676
R707 B.n264 B.n263 71.676
R708 B.n257 B.n157 71.676
R709 B.n256 B.n255 71.676
R710 B.n249 B.n159 71.676
R711 B.n248 B.n247 71.676
R712 B.n240 B.n161 71.676
R713 B.n239 B.n238 71.676
R714 B.n232 B.n165 71.676
R715 B.n231 B.n230 71.676
R716 B.n223 B.n167 71.676
R717 B.n222 B.n221 71.676
R718 B.n215 B.n171 71.676
R719 B.n214 B.n213 71.676
R720 B.n207 B.n173 71.676
R721 B.n206 B.n205 71.676
R722 B.n199 B.n175 71.676
R723 B.n198 B.n197 71.676
R724 B.n191 B.n177 71.676
R725 B.n190 B.n189 71.676
R726 B.n183 B.n179 71.676
R727 B.n182 B.n181 71.676
R728 B.n526 B.n58 71.676
R729 B.n525 B.n524 71.676
R730 B.n518 B.n60 71.676
R731 B.n517 B.n516 71.676
R732 B.n510 B.n62 71.676
R733 B.n509 B.n508 71.676
R734 B.n502 B.n64 71.676
R735 B.n501 B.n500 71.676
R736 B.n494 B.n66 71.676
R737 B.n493 B.n492 71.676
R738 B.n486 B.n68 71.676
R739 B.n485 B.n484 71.676
R740 B.n478 B.n70 71.676
R741 B.n477 B.n476 71.676
R742 B.n470 B.n75 71.676
R743 B.n469 B.n468 71.676
R744 B.n461 B.n77 71.676
R745 B.n460 B.n459 71.676
R746 B.n453 B.n81 71.676
R747 B.n452 B.n451 71.676
R748 B.n445 B.n83 71.676
R749 B.n444 B.n443 71.676
R750 B.n437 B.n85 71.676
R751 B.n436 B.n435 71.676
R752 B.n429 B.n87 71.676
R753 B.n428 B.n427 71.676
R754 B.n421 B.n89 71.676
R755 B.n422 B.n421 71.676
R756 B.n427 B.n426 71.676
R757 B.n430 B.n429 71.676
R758 B.n435 B.n434 71.676
R759 B.n438 B.n437 71.676
R760 B.n443 B.n442 71.676
R761 B.n446 B.n445 71.676
R762 B.n451 B.n450 71.676
R763 B.n454 B.n453 71.676
R764 B.n459 B.n458 71.676
R765 B.n462 B.n461 71.676
R766 B.n468 B.n467 71.676
R767 B.n471 B.n470 71.676
R768 B.n476 B.n475 71.676
R769 B.n479 B.n478 71.676
R770 B.n484 B.n483 71.676
R771 B.n487 B.n486 71.676
R772 B.n492 B.n491 71.676
R773 B.n495 B.n494 71.676
R774 B.n500 B.n499 71.676
R775 B.n503 B.n502 71.676
R776 B.n508 B.n507 71.676
R777 B.n511 B.n510 71.676
R778 B.n516 B.n515 71.676
R779 B.n519 B.n518 71.676
R780 B.n524 B.n523 71.676
R781 B.n527 B.n526 71.676
R782 B.n287 B.n286 71.676
R783 B.n281 B.n151 71.676
R784 B.n279 B.n278 71.676
R785 B.n274 B.n273 71.676
R786 B.n271 B.n270 71.676
R787 B.n266 B.n265 71.676
R788 B.n263 B.n262 71.676
R789 B.n258 B.n257 71.676
R790 B.n255 B.n254 71.676
R791 B.n250 B.n249 71.676
R792 B.n247 B.n246 71.676
R793 B.n241 B.n240 71.676
R794 B.n238 B.n237 71.676
R795 B.n233 B.n232 71.676
R796 B.n230 B.n229 71.676
R797 B.n224 B.n223 71.676
R798 B.n221 B.n220 71.676
R799 B.n216 B.n215 71.676
R800 B.n213 B.n212 71.676
R801 B.n208 B.n207 71.676
R802 B.n205 B.n204 71.676
R803 B.n200 B.n199 71.676
R804 B.n197 B.n196 71.676
R805 B.n192 B.n191 71.676
R806 B.n189 B.n188 71.676
R807 B.n184 B.n183 71.676
R808 B.n181 B.n147 71.676
R809 B.n169 B.t15 71.4903
R810 B.n79 B.t19 71.4903
R811 B.n163 B.t12 71.4845
R812 B.n72 B.t9 71.4845
R813 B.n292 B.n144 69.2277
R814 B.n298 B.n144 69.2277
R815 B.n298 B.n139 69.2277
R816 B.n304 B.n139 69.2277
R817 B.n304 B.n140 69.2277
R818 B.n310 B.n132 69.2277
R819 B.n316 B.n132 69.2277
R820 B.n316 B.n128 69.2277
R821 B.n322 B.n128 69.2277
R822 B.n322 B.n123 69.2277
R823 B.n328 B.n123 69.2277
R824 B.n328 B.n124 69.2277
R825 B.n334 B.n115 69.2277
R826 B.n340 B.n115 69.2277
R827 B.n340 B.n116 69.2277
R828 B.n346 B.n107 69.2277
R829 B.n352 B.n107 69.2277
R830 B.n352 B.n108 69.2277
R831 B.n358 B.n100 69.2277
R832 B.n364 B.n100 69.2277
R833 B.n364 B.n96 69.2277
R834 B.n371 B.n96 69.2277
R835 B.n377 B.n92 69.2277
R836 B.n377 B.n4 69.2277
R837 B.n590 B.n4 69.2277
R838 B.n590 B.n589 69.2277
R839 B.n589 B.n588 69.2277
R840 B.n588 B.n8 69.2277
R841 B.n582 B.n581 69.2277
R842 B.n581 B.n580 69.2277
R843 B.n580 B.n15 69.2277
R844 B.n574 B.n15 69.2277
R845 B.n573 B.n572 69.2277
R846 B.n572 B.n22 69.2277
R847 B.n566 B.n22 69.2277
R848 B.n565 B.n564 69.2277
R849 B.n564 B.n29 69.2277
R850 B.n558 B.n29 69.2277
R851 B.n557 B.n556 69.2277
R852 B.n556 B.n36 69.2277
R853 B.n550 B.n36 69.2277
R854 B.n550 B.n549 69.2277
R855 B.n549 B.n548 69.2277
R856 B.n548 B.n43 69.2277
R857 B.n542 B.n43 69.2277
R858 B.n541 B.n540 69.2277
R859 B.n540 B.n50 69.2277
R860 B.n534 B.n50 69.2277
R861 B.n534 B.n533 69.2277
R862 B.n533 B.n532 69.2277
R863 B.n334 B.t0 65.1555
R864 B.n558 B.t3 65.1555
R865 B.n226 B.n169 59.5399
R866 B.n244 B.n163 59.5399
R867 B.n73 B.n72 59.5399
R868 B.n465 B.n79 59.5399
R869 B.n108 B.t4 57.0111
R870 B.t1 B.n573 57.0111
R871 B.t5 B.n92 54.975
R872 B.t2 B.n8 54.975
R873 B.n346 B.t21 38.6863
R874 B.n566 B.t20 38.6863
R875 B.n310 B.t11 36.6502
R876 B.n542 B.t7 36.6502
R877 B.n140 B.t11 32.578
R878 B.t7 B.n541 32.578
R879 B.n530 B.n529 31.3761
R880 B.n419 B.n418 31.3761
R881 B.n294 B.n146 31.3761
R882 B.n290 B.n289 31.3761
R883 B.n116 B.t21 30.5419
R884 B.t20 B.n565 30.5419
R885 B.n169 B.n168 28.8975
R886 B.n163 B.n162 28.8975
R887 B.n72 B.n71 28.8975
R888 B.n79 B.n78 28.8975
R889 B B.n592 18.0485
R890 B.n371 B.t5 14.2532
R891 B.n582 B.t2 14.2532
R892 B.n358 B.t4 12.2171
R893 B.n574 B.t1 12.2171
R894 B.n529 B.n528 10.6151
R895 B.n528 B.n59 10.6151
R896 B.n522 B.n59 10.6151
R897 B.n522 B.n521 10.6151
R898 B.n521 B.n520 10.6151
R899 B.n520 B.n61 10.6151
R900 B.n514 B.n61 10.6151
R901 B.n514 B.n513 10.6151
R902 B.n513 B.n512 10.6151
R903 B.n512 B.n63 10.6151
R904 B.n506 B.n63 10.6151
R905 B.n506 B.n505 10.6151
R906 B.n505 B.n504 10.6151
R907 B.n504 B.n65 10.6151
R908 B.n498 B.n65 10.6151
R909 B.n498 B.n497 10.6151
R910 B.n497 B.n496 10.6151
R911 B.n496 B.n67 10.6151
R912 B.n490 B.n67 10.6151
R913 B.n490 B.n489 10.6151
R914 B.n489 B.n488 10.6151
R915 B.n488 B.n69 10.6151
R916 B.n482 B.n481 10.6151
R917 B.n481 B.n480 10.6151
R918 B.n480 B.n74 10.6151
R919 B.n474 B.n74 10.6151
R920 B.n474 B.n473 10.6151
R921 B.n473 B.n472 10.6151
R922 B.n472 B.n76 10.6151
R923 B.n466 B.n76 10.6151
R924 B.n464 B.n463 10.6151
R925 B.n463 B.n80 10.6151
R926 B.n457 B.n80 10.6151
R927 B.n457 B.n456 10.6151
R928 B.n456 B.n455 10.6151
R929 B.n455 B.n82 10.6151
R930 B.n449 B.n82 10.6151
R931 B.n449 B.n448 10.6151
R932 B.n448 B.n447 10.6151
R933 B.n447 B.n84 10.6151
R934 B.n441 B.n84 10.6151
R935 B.n441 B.n440 10.6151
R936 B.n440 B.n439 10.6151
R937 B.n439 B.n86 10.6151
R938 B.n433 B.n86 10.6151
R939 B.n433 B.n432 10.6151
R940 B.n432 B.n431 10.6151
R941 B.n431 B.n88 10.6151
R942 B.n425 B.n88 10.6151
R943 B.n425 B.n424 10.6151
R944 B.n424 B.n423 10.6151
R945 B.n423 B.n419 10.6151
R946 B.n295 B.n294 10.6151
R947 B.n296 B.n295 10.6151
R948 B.n296 B.n137 10.6151
R949 B.n306 B.n137 10.6151
R950 B.n307 B.n306 10.6151
R951 B.n308 B.n307 10.6151
R952 B.n308 B.n130 10.6151
R953 B.n318 B.n130 10.6151
R954 B.n319 B.n318 10.6151
R955 B.n320 B.n319 10.6151
R956 B.n320 B.n121 10.6151
R957 B.n330 B.n121 10.6151
R958 B.n331 B.n330 10.6151
R959 B.n332 B.n331 10.6151
R960 B.n332 B.n113 10.6151
R961 B.n342 B.n113 10.6151
R962 B.n343 B.n342 10.6151
R963 B.n344 B.n343 10.6151
R964 B.n344 B.n105 10.6151
R965 B.n354 B.n105 10.6151
R966 B.n355 B.n354 10.6151
R967 B.n356 B.n355 10.6151
R968 B.n356 B.n98 10.6151
R969 B.n366 B.n98 10.6151
R970 B.n367 B.n366 10.6151
R971 B.n369 B.n367 10.6151
R972 B.n369 B.n368 10.6151
R973 B.n368 B.n90 10.6151
R974 B.n380 B.n90 10.6151
R975 B.n381 B.n380 10.6151
R976 B.n382 B.n381 10.6151
R977 B.n383 B.n382 10.6151
R978 B.n385 B.n383 10.6151
R979 B.n386 B.n385 10.6151
R980 B.n387 B.n386 10.6151
R981 B.n388 B.n387 10.6151
R982 B.n390 B.n388 10.6151
R983 B.n391 B.n390 10.6151
R984 B.n392 B.n391 10.6151
R985 B.n393 B.n392 10.6151
R986 B.n395 B.n393 10.6151
R987 B.n396 B.n395 10.6151
R988 B.n397 B.n396 10.6151
R989 B.n398 B.n397 10.6151
R990 B.n400 B.n398 10.6151
R991 B.n401 B.n400 10.6151
R992 B.n402 B.n401 10.6151
R993 B.n403 B.n402 10.6151
R994 B.n405 B.n403 10.6151
R995 B.n406 B.n405 10.6151
R996 B.n407 B.n406 10.6151
R997 B.n408 B.n407 10.6151
R998 B.n410 B.n408 10.6151
R999 B.n411 B.n410 10.6151
R1000 B.n412 B.n411 10.6151
R1001 B.n413 B.n412 10.6151
R1002 B.n415 B.n413 10.6151
R1003 B.n416 B.n415 10.6151
R1004 B.n417 B.n416 10.6151
R1005 B.n418 B.n417 10.6151
R1006 B.n289 B.n288 10.6151
R1007 B.n288 B.n150 10.6151
R1008 B.n283 B.n150 10.6151
R1009 B.n283 B.n282 10.6151
R1010 B.n282 B.n152 10.6151
R1011 B.n277 B.n152 10.6151
R1012 B.n277 B.n276 10.6151
R1013 B.n276 B.n275 10.6151
R1014 B.n275 B.n154 10.6151
R1015 B.n269 B.n154 10.6151
R1016 B.n269 B.n268 10.6151
R1017 B.n268 B.n267 10.6151
R1018 B.n267 B.n156 10.6151
R1019 B.n261 B.n156 10.6151
R1020 B.n261 B.n260 10.6151
R1021 B.n260 B.n259 10.6151
R1022 B.n259 B.n158 10.6151
R1023 B.n253 B.n158 10.6151
R1024 B.n253 B.n252 10.6151
R1025 B.n252 B.n251 10.6151
R1026 B.n251 B.n160 10.6151
R1027 B.n245 B.n160 10.6151
R1028 B.n243 B.n242 10.6151
R1029 B.n242 B.n164 10.6151
R1030 B.n236 B.n164 10.6151
R1031 B.n236 B.n235 10.6151
R1032 B.n235 B.n234 10.6151
R1033 B.n234 B.n166 10.6151
R1034 B.n228 B.n166 10.6151
R1035 B.n228 B.n227 10.6151
R1036 B.n225 B.n170 10.6151
R1037 B.n219 B.n170 10.6151
R1038 B.n219 B.n218 10.6151
R1039 B.n218 B.n217 10.6151
R1040 B.n217 B.n172 10.6151
R1041 B.n211 B.n172 10.6151
R1042 B.n211 B.n210 10.6151
R1043 B.n210 B.n209 10.6151
R1044 B.n209 B.n174 10.6151
R1045 B.n203 B.n174 10.6151
R1046 B.n203 B.n202 10.6151
R1047 B.n202 B.n201 10.6151
R1048 B.n201 B.n176 10.6151
R1049 B.n195 B.n176 10.6151
R1050 B.n195 B.n194 10.6151
R1051 B.n194 B.n193 10.6151
R1052 B.n193 B.n178 10.6151
R1053 B.n187 B.n178 10.6151
R1054 B.n187 B.n186 10.6151
R1055 B.n186 B.n185 10.6151
R1056 B.n185 B.n180 10.6151
R1057 B.n180 B.n146 10.6151
R1058 B.n290 B.n142 10.6151
R1059 B.n300 B.n142 10.6151
R1060 B.n301 B.n300 10.6151
R1061 B.n302 B.n301 10.6151
R1062 B.n302 B.n134 10.6151
R1063 B.n312 B.n134 10.6151
R1064 B.n313 B.n312 10.6151
R1065 B.n314 B.n313 10.6151
R1066 B.n314 B.n126 10.6151
R1067 B.n324 B.n126 10.6151
R1068 B.n325 B.n324 10.6151
R1069 B.n326 B.n325 10.6151
R1070 B.n326 B.n118 10.6151
R1071 B.n336 B.n118 10.6151
R1072 B.n337 B.n336 10.6151
R1073 B.n338 B.n337 10.6151
R1074 B.n338 B.n110 10.6151
R1075 B.n348 B.n110 10.6151
R1076 B.n349 B.n348 10.6151
R1077 B.n350 B.n349 10.6151
R1078 B.n350 B.n102 10.6151
R1079 B.n360 B.n102 10.6151
R1080 B.n361 B.n360 10.6151
R1081 B.n362 B.n361 10.6151
R1082 B.n362 B.n94 10.6151
R1083 B.n373 B.n94 10.6151
R1084 B.n374 B.n373 10.6151
R1085 B.n375 B.n374 10.6151
R1086 B.n375 B.n0 10.6151
R1087 B.n586 B.n1 10.6151
R1088 B.n586 B.n585 10.6151
R1089 B.n585 B.n584 10.6151
R1090 B.n584 B.n10 10.6151
R1091 B.n578 B.n10 10.6151
R1092 B.n578 B.n577 10.6151
R1093 B.n577 B.n576 10.6151
R1094 B.n576 B.n17 10.6151
R1095 B.n570 B.n17 10.6151
R1096 B.n570 B.n569 10.6151
R1097 B.n569 B.n568 10.6151
R1098 B.n568 B.n24 10.6151
R1099 B.n562 B.n24 10.6151
R1100 B.n562 B.n561 10.6151
R1101 B.n561 B.n560 10.6151
R1102 B.n560 B.n31 10.6151
R1103 B.n554 B.n31 10.6151
R1104 B.n554 B.n553 10.6151
R1105 B.n553 B.n552 10.6151
R1106 B.n552 B.n38 10.6151
R1107 B.n546 B.n38 10.6151
R1108 B.n546 B.n545 10.6151
R1109 B.n545 B.n544 10.6151
R1110 B.n544 B.n45 10.6151
R1111 B.n538 B.n45 10.6151
R1112 B.n538 B.n537 10.6151
R1113 B.n537 B.n536 10.6151
R1114 B.n536 B.n52 10.6151
R1115 B.n530 B.n52 10.6151
R1116 B.n482 B.n73 6.5566
R1117 B.n466 B.n465 6.5566
R1118 B.n244 B.n243 6.5566
R1119 B.n227 B.n226 6.5566
R1120 B.n124 B.t0 4.07269
R1121 B.t3 B.n557 4.07269
R1122 B.n73 B.n69 4.05904
R1123 B.n465 B.n464 4.05904
R1124 B.n245 B.n244 4.05904
R1125 B.n226 B.n225 4.05904
R1126 B.n592 B.n0 2.81026
R1127 B.n592 B.n1 2.81026
R1128 VP.n23 VP.n5 174.268
R1129 VP.n40 VP.n39 174.268
R1130 VP.n22 VP.n21 174.268
R1131 VP.n12 VP.n11 161.3
R1132 VP.n13 VP.n8 161.3
R1133 VP.n16 VP.n15 161.3
R1134 VP.n17 VP.n7 161.3
R1135 VP.n19 VP.n18 161.3
R1136 VP.n20 VP.n6 161.3
R1137 VP.n38 VP.n0 161.3
R1138 VP.n37 VP.n36 161.3
R1139 VP.n35 VP.n1 161.3
R1140 VP.n34 VP.n33 161.3
R1141 VP.n31 VP.n2 161.3
R1142 VP.n30 VP.n29 161.3
R1143 VP.n28 VP.n27 161.3
R1144 VP.n26 VP.n4 161.3
R1145 VP.n25 VP.n24 161.3
R1146 VP.n10 VP.t3 144.495
R1147 VP.n5 VP.t7 114.891
R1148 VP.n3 VP.t5 114.891
R1149 VP.n32 VP.t1 114.891
R1150 VP.n39 VP.t6 114.891
R1151 VP.n21 VP.t4 114.891
R1152 VP.n14 VP.t0 114.891
R1153 VP.n9 VP.t2 114.891
R1154 VP.n10 VP.n9 51.7518
R1155 VP.n27 VP.n26 41.4647
R1156 VP.n37 VP.n1 41.4647
R1157 VP.n19 VP.n7 41.4647
R1158 VP.n31 VP.n30 40.4934
R1159 VP.n33 VP.n31 40.4934
R1160 VP.n15 VP.n13 40.4934
R1161 VP.n13 VP.n12 40.4934
R1162 VP.n26 VP.n25 39.5221
R1163 VP.n38 VP.n37 39.5221
R1164 VP.n20 VP.n19 39.5221
R1165 VP.n23 VP.n22 39.1217
R1166 VP.n11 VP.n10 27.1667
R1167 VP.n27 VP.n3 12.4787
R1168 VP.n32 VP.n1 12.4787
R1169 VP.n14 VP.n7 12.4787
R1170 VP.n30 VP.n3 11.9893
R1171 VP.n33 VP.n32 11.9893
R1172 VP.n15 VP.n14 11.9893
R1173 VP.n12 VP.n9 11.9893
R1174 VP.n25 VP.n5 11.5
R1175 VP.n39 VP.n38 11.5
R1176 VP.n21 VP.n20 11.5
R1177 VP.n11 VP.n8 0.189894
R1178 VP.n16 VP.n8 0.189894
R1179 VP.n17 VP.n16 0.189894
R1180 VP.n18 VP.n17 0.189894
R1181 VP.n18 VP.n6 0.189894
R1182 VP.n22 VP.n6 0.189894
R1183 VP.n24 VP.n23 0.189894
R1184 VP.n24 VP.n4 0.189894
R1185 VP.n28 VP.n4 0.189894
R1186 VP.n29 VP.n28 0.189894
R1187 VP.n29 VP.n2 0.189894
R1188 VP.n34 VP.n2 0.189894
R1189 VP.n35 VP.n34 0.189894
R1190 VP.n36 VP.n35 0.189894
R1191 VP.n36 VP.n0 0.189894
R1192 VP.n40 VP.n0 0.189894
R1193 VP VP.n40 0.0516364
R1194 VDD1 VDD1.n0 66.4371
R1195 VDD1.n3 VDD1.n2 66.3234
R1196 VDD1.n3 VDD1.n1 66.3234
R1197 VDD1.n5 VDD1.n4 65.7365
R1198 VDD1.n5 VDD1.n3 34.8457
R1199 VDD1.n4 VDD1.t7 3.58097
R1200 VDD1.n4 VDD1.t3 3.58097
R1201 VDD1.n0 VDD1.t4 3.58097
R1202 VDD1.n0 VDD1.t5 3.58097
R1203 VDD1.n2 VDD1.t6 3.58097
R1204 VDD1.n2 VDD1.t1 3.58097
R1205 VDD1.n1 VDD1.t0 3.58097
R1206 VDD1.n1 VDD1.t2 3.58097
R1207 VDD1 VDD1.n5 0.584552
C0 VP VDD1 3.6334f
C1 VN VDD2 3.41675f
C2 VN VP 4.70738f
C3 VP VDD2 0.365931f
C4 VTAIL VDD1 5.57725f
C5 VN VTAIL 3.68784f
C6 VN VDD1 0.148616f
C7 VTAIL VDD2 5.62201f
C8 VDD1 VDD2 1.05283f
C9 VP VTAIL 3.70194f
C10 VDD2 B 3.413425f
C11 VDD1 B 3.6995f
C12 VTAIL B 5.4244f
C13 VN B 9.41679f
C14 VP B 7.897849f
C15 VDD1.t4 B 0.111374f
C16 VDD1.t5 B 0.111374f
C17 VDD1.n0 B 0.922739f
C18 VDD1.t0 B 0.111374f
C19 VDD1.t2 B 0.111374f
C20 VDD1.n1 B 0.922019f
C21 VDD1.t6 B 0.111374f
C22 VDD1.t1 B 0.111374f
C23 VDD1.n2 B 0.922019f
C24 VDD1.n3 B 2.13744f
C25 VDD1.t7 B 0.111374f
C26 VDD1.t3 B 0.111374f
C27 VDD1.n4 B 0.918737f
C28 VDD1.n5 B 2.00544f
C29 VP.n0 B 0.038168f
C30 VP.t6 B 0.644797f
C31 VP.n1 B 0.058241f
C32 VP.n2 B 0.038168f
C33 VP.t5 B 0.644797f
C34 VP.n3 B 0.263835f
C35 VP.n4 B 0.038168f
C36 VP.t7 B 0.644797f
C37 VP.n5 B 0.322849f
C38 VP.n6 B 0.038168f
C39 VP.t4 B 0.644797f
C40 VP.n7 B 0.058241f
C41 VP.n8 B 0.038168f
C42 VP.t2 B 0.644797f
C43 VP.n9 B 0.318861f
C44 VP.t3 B 0.721204f
C45 VP.n10 B 0.340027f
C46 VP.n11 B 0.196779f
C47 VP.n12 B 0.057945f
C48 VP.n13 B 0.030855f
C49 VP.t0 B 0.644797f
C50 VP.n14 B 0.263835f
C51 VP.n15 B 0.057945f
C52 VP.n16 B 0.038168f
C53 VP.n17 B 0.038168f
C54 VP.n18 B 0.038168f
C55 VP.n19 B 0.030904f
C56 VP.n20 B 0.057601f
C57 VP.n21 B 0.322849f
C58 VP.n22 B 1.40019f
C59 VP.n23 B 1.43526f
C60 VP.n24 B 0.038168f
C61 VP.n25 B 0.057601f
C62 VP.n26 B 0.030904f
C63 VP.n27 B 0.058241f
C64 VP.n28 B 0.038168f
C65 VP.n29 B 0.038168f
C66 VP.n30 B 0.057945f
C67 VP.n31 B 0.030855f
C68 VP.t1 B 0.644797f
C69 VP.n32 B 0.263835f
C70 VP.n33 B 0.057945f
C71 VP.n34 B 0.038168f
C72 VP.n35 B 0.038168f
C73 VP.n36 B 0.038168f
C74 VP.n37 B 0.030904f
C75 VP.n38 B 0.057601f
C76 VP.n39 B 0.322849f
C77 VP.n40 B 0.034323f
C78 VDD2.t2 B 0.110079f
C79 VDD2.t7 B 0.110079f
C80 VDD2.n0 B 0.9113f
C81 VDD2.t4 B 0.110079f
C82 VDD2.t1 B 0.110079f
C83 VDD2.n1 B 0.9113f
C84 VDD2.n2 B 2.05896f
C85 VDD2.t0 B 0.110079f
C86 VDD2.t6 B 0.110079f
C87 VDD2.n3 B 0.90806f
C88 VDD2.n4 B 1.95216f
C89 VDD2.t5 B 0.110079f
C90 VDD2.t3 B 0.110079f
C91 VDD2.n5 B 0.911273f
C92 VTAIL.t15 B 0.095838f
C93 VTAIL.t8 B 0.095838f
C94 VTAIL.n0 B 0.731773f
C95 VTAIL.n1 B 0.301018f
C96 VTAIL.t11 B 0.932113f
C97 VTAIL.n2 B 0.391143f
C98 VTAIL.t5 B 0.932113f
C99 VTAIL.n3 B 0.391143f
C100 VTAIL.t7 B 0.095838f
C101 VTAIL.t4 B 0.095838f
C102 VTAIL.n4 B 0.731773f
C103 VTAIL.n5 B 0.387676f
C104 VTAIL.t0 B 0.932113f
C105 VTAIL.n6 B 1.0835f
C106 VTAIL.t14 B 0.932118f
C107 VTAIL.n7 B 1.0835f
C108 VTAIL.t10 B 0.095838f
C109 VTAIL.t13 B 0.095838f
C110 VTAIL.n8 B 0.731777f
C111 VTAIL.n9 B 0.387672f
C112 VTAIL.t12 B 0.932118f
C113 VTAIL.n10 B 0.391139f
C114 VTAIL.t2 B 0.932118f
C115 VTAIL.n11 B 0.391139f
C116 VTAIL.t1 B 0.095838f
C117 VTAIL.t6 B 0.095838f
C118 VTAIL.n12 B 0.731777f
C119 VTAIL.n13 B 0.387672f
C120 VTAIL.t3 B 0.932113f
C121 VTAIL.n14 B 1.0835f
C122 VTAIL.t9 B 0.932113f
C123 VTAIL.n15 B 1.07939f
C124 VN.n0 B 0.037365f
C125 VN.t6 B 0.631228f
C126 VN.n1 B 0.057015f
C127 VN.n2 B 0.037365f
C128 VN.t0 B 0.631228f
C129 VN.n3 B 0.312151f
C130 VN.t5 B 0.706027f
C131 VN.n4 B 0.332872f
C132 VN.n5 B 0.192638f
C133 VN.n6 B 0.056726f
C134 VN.n7 B 0.030206f
C135 VN.t3 B 0.631228f
C136 VN.n8 B 0.258283f
C137 VN.n9 B 0.056726f
C138 VN.n10 B 0.037365f
C139 VN.n11 B 0.037365f
C140 VN.n12 B 0.037365f
C141 VN.n13 B 0.030254f
C142 VN.n14 B 0.056389f
C143 VN.n15 B 0.316056f
C144 VN.n16 B 0.033601f
C145 VN.n17 B 0.037365f
C146 VN.t7 B 0.631228f
C147 VN.n18 B 0.057015f
C148 VN.n19 B 0.037365f
C149 VN.t1 B 0.631228f
C150 VN.n20 B 0.258283f
C151 VN.t2 B 0.631228f
C152 VN.n21 B 0.312151f
C153 VN.t4 B 0.706027f
C154 VN.n22 B 0.332872f
C155 VN.n23 B 0.192638f
C156 VN.n24 B 0.056726f
C157 VN.n25 B 0.030206f
C158 VN.n26 B 0.056726f
C159 VN.n27 B 0.037365f
C160 VN.n28 B 0.037365f
C161 VN.n29 B 0.037365f
C162 VN.n30 B 0.030254f
C163 VN.n31 B 0.056389f
C164 VN.n32 B 0.316056f
C165 VN.n33 B 1.39536f
.ends

