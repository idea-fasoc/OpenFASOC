* NGSPICE file created from diff_pair_sample_0300.ext - technology: sky130A

.subckt diff_pair_sample_0300 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t7 B.t9 sky130_fd_pr__nfet_01v8 ad=2.65815 pd=16.44 as=2.65815 ps=16.44 w=16.11 l=2.34
X1 VTAIL.t0 VN.t0 VDD2.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=2.65815 pd=16.44 as=2.65815 ps=16.44 w=16.11 l=2.34
X2 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=6.2829 pd=33 as=0 ps=0 w=16.11 l=2.34
X3 VTAIL.t4 VN.t1 VDD2.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=2.65815 pd=16.44 as=2.65815 ps=16.44 w=16.11 l=2.34
X4 VDD1.t6 VP.t1 VTAIL.t18 B.t8 sky130_fd_pr__nfet_01v8 ad=2.65815 pd=16.44 as=6.2829 ps=33 w=16.11 l=2.34
X5 VTAIL.t5 VN.t2 VDD2.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=2.65815 pd=16.44 as=2.65815 ps=16.44 w=16.11 l=2.34
X6 VDD1.t3 VP.t2 VTAIL.t17 B.t7 sky130_fd_pr__nfet_01v8 ad=2.65815 pd=16.44 as=2.65815 ps=16.44 w=16.11 l=2.34
X7 VDD1.t2 VP.t3 VTAIL.t16 B.t6 sky130_fd_pr__nfet_01v8 ad=2.65815 pd=16.44 as=6.2829 ps=33 w=16.11 l=2.34
X8 VTAIL.t9 VN.t3 VDD2.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=2.65815 pd=16.44 as=2.65815 ps=16.44 w=16.11 l=2.34
X9 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=6.2829 pd=33 as=0 ps=0 w=16.11 l=2.34
X10 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=6.2829 pd=33 as=0 ps=0 w=16.11 l=2.34
X11 VDD1.t5 VP.t4 VTAIL.t15 B.t3 sky130_fd_pr__nfet_01v8 ad=2.65815 pd=16.44 as=2.65815 ps=16.44 w=16.11 l=2.34
X12 VDD1.t4 VP.t5 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=6.2829 pd=33 as=2.65815 ps=16.44 w=16.11 l=2.34
X13 VDD2.t5 VN.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.2829 pd=33 as=2.65815 ps=16.44 w=16.11 l=2.34
X14 VDD1.t9 VP.t6 VTAIL.t13 B.t2 sky130_fd_pr__nfet_01v8 ad=6.2829 pd=33 as=2.65815 ps=16.44 w=16.11 l=2.34
X15 VDD2.t4 VN.t5 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.65815 pd=16.44 as=6.2829 ps=33 w=16.11 l=2.34
X16 VDD2.t3 VN.t6 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.65815 pd=16.44 as=2.65815 ps=16.44 w=16.11 l=2.34
X17 VTAIL.t12 VP.t7 VDD1.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=2.65815 pd=16.44 as=2.65815 ps=16.44 w=16.11 l=2.34
X18 VDD2.t2 VN.t7 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.2829 pd=33 as=2.65815 ps=16.44 w=16.11 l=2.34
X19 VTAIL.t11 VP.t8 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.65815 pd=16.44 as=2.65815 ps=16.44 w=16.11 l=2.34
X20 VDD2.t1 VN.t8 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.65815 pd=16.44 as=2.65815 ps=16.44 w=16.11 l=2.34
X21 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.2829 pd=33 as=0 ps=0 w=16.11 l=2.34
X22 VDD2.t0 VN.t9 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=2.65815 pd=16.44 as=6.2829 ps=33 w=16.11 l=2.34
X23 VTAIL.t10 VP.t9 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=2.65815 pd=16.44 as=2.65815 ps=16.44 w=16.11 l=2.34
R0 VP.n19 VP.t5 198.988
R1 VP.n5 VP.t4 165.919
R2 VP.n49 VP.t6 165.919
R3 VP.n57 VP.t0 165.919
R4 VP.n75 VP.t9 165.919
R5 VP.n83 VP.t3 165.919
R6 VP.n16 VP.t2 165.919
R7 VP.n46 VP.t1 165.919
R8 VP.n38 VP.t7 165.919
R9 VP.n20 VP.t8 165.919
R10 VP.n22 VP.n21 161.3
R11 VP.n23 VP.n18 161.3
R12 VP.n25 VP.n24 161.3
R13 VP.n26 VP.n17 161.3
R14 VP.n28 VP.n27 161.3
R15 VP.n29 VP.n16 161.3
R16 VP.n31 VP.n30 161.3
R17 VP.n32 VP.n15 161.3
R18 VP.n34 VP.n33 161.3
R19 VP.n35 VP.n14 161.3
R20 VP.n37 VP.n36 161.3
R21 VP.n39 VP.n13 161.3
R22 VP.n41 VP.n40 161.3
R23 VP.n42 VP.n12 161.3
R24 VP.n44 VP.n43 161.3
R25 VP.n45 VP.n11 161.3
R26 VP.n82 VP.n0 161.3
R27 VP.n81 VP.n80 161.3
R28 VP.n79 VP.n1 161.3
R29 VP.n78 VP.n77 161.3
R30 VP.n76 VP.n2 161.3
R31 VP.n74 VP.n73 161.3
R32 VP.n72 VP.n3 161.3
R33 VP.n71 VP.n70 161.3
R34 VP.n69 VP.n4 161.3
R35 VP.n68 VP.n67 161.3
R36 VP.n66 VP.n5 161.3
R37 VP.n65 VP.n64 161.3
R38 VP.n63 VP.n6 161.3
R39 VP.n62 VP.n61 161.3
R40 VP.n60 VP.n7 161.3
R41 VP.n59 VP.n58 161.3
R42 VP.n56 VP.n8 161.3
R43 VP.n55 VP.n54 161.3
R44 VP.n53 VP.n9 161.3
R45 VP.n52 VP.n51 161.3
R46 VP.n50 VP.n10 161.3
R47 VP.n49 VP.n48 94.1189
R48 VP.n84 VP.n83 94.1189
R49 VP.n47 VP.n46 94.1189
R50 VP.n20 VP.n19 63.5395
R51 VP.n63 VP.n62 56.5193
R52 VP.n70 VP.n69 56.5193
R53 VP.n33 VP.n32 56.5193
R54 VP.n26 VP.n25 56.5193
R55 VP.n48 VP.n47 54.8746
R56 VP.n51 VP.n9 40.979
R57 VP.n81 VP.n1 40.979
R58 VP.n44 VP.n12 40.979
R59 VP.n55 VP.n9 40.0078
R60 VP.n77 VP.n1 40.0078
R61 VP.n40 VP.n12 40.0078
R62 VP.n51 VP.n50 24.4675
R63 VP.n56 VP.n55 24.4675
R64 VP.n58 VP.n7 24.4675
R65 VP.n62 VP.n7 24.4675
R66 VP.n64 VP.n63 24.4675
R67 VP.n64 VP.n5 24.4675
R68 VP.n68 VP.n5 24.4675
R69 VP.n69 VP.n68 24.4675
R70 VP.n70 VP.n3 24.4675
R71 VP.n74 VP.n3 24.4675
R72 VP.n77 VP.n76 24.4675
R73 VP.n82 VP.n81 24.4675
R74 VP.n45 VP.n44 24.4675
R75 VP.n33 VP.n14 24.4675
R76 VP.n37 VP.n14 24.4675
R77 VP.n40 VP.n39 24.4675
R78 VP.n27 VP.n26 24.4675
R79 VP.n27 VP.n16 24.4675
R80 VP.n31 VP.n16 24.4675
R81 VP.n32 VP.n31 24.4675
R82 VP.n21 VP.n18 24.4675
R83 VP.n25 VP.n18 24.4675
R84 VP.n50 VP.n49 16.6381
R85 VP.n83 VP.n82 16.6381
R86 VP.n46 VP.n45 16.6381
R87 VP.n57 VP.n56 16.1487
R88 VP.n76 VP.n75 16.1487
R89 VP.n39 VP.n38 16.1487
R90 VP.n22 VP.n19 9.31187
R91 VP.n58 VP.n57 8.31928
R92 VP.n75 VP.n74 8.31928
R93 VP.n38 VP.n37 8.31928
R94 VP.n21 VP.n20 8.31928
R95 VP.n47 VP.n11 0.278367
R96 VP.n48 VP.n10 0.278367
R97 VP.n84 VP.n0 0.278367
R98 VP.n23 VP.n22 0.189894
R99 VP.n24 VP.n23 0.189894
R100 VP.n24 VP.n17 0.189894
R101 VP.n28 VP.n17 0.189894
R102 VP.n29 VP.n28 0.189894
R103 VP.n30 VP.n29 0.189894
R104 VP.n30 VP.n15 0.189894
R105 VP.n34 VP.n15 0.189894
R106 VP.n35 VP.n34 0.189894
R107 VP.n36 VP.n35 0.189894
R108 VP.n36 VP.n13 0.189894
R109 VP.n41 VP.n13 0.189894
R110 VP.n42 VP.n41 0.189894
R111 VP.n43 VP.n42 0.189894
R112 VP.n43 VP.n11 0.189894
R113 VP.n52 VP.n10 0.189894
R114 VP.n53 VP.n52 0.189894
R115 VP.n54 VP.n53 0.189894
R116 VP.n54 VP.n8 0.189894
R117 VP.n59 VP.n8 0.189894
R118 VP.n60 VP.n59 0.189894
R119 VP.n61 VP.n60 0.189894
R120 VP.n61 VP.n6 0.189894
R121 VP.n65 VP.n6 0.189894
R122 VP.n66 VP.n65 0.189894
R123 VP.n67 VP.n66 0.189894
R124 VP.n67 VP.n4 0.189894
R125 VP.n71 VP.n4 0.189894
R126 VP.n72 VP.n71 0.189894
R127 VP.n73 VP.n72 0.189894
R128 VP.n73 VP.n2 0.189894
R129 VP.n78 VP.n2 0.189894
R130 VP.n79 VP.n78 0.189894
R131 VP.n80 VP.n79 0.189894
R132 VP.n80 VP.n0 0.189894
R133 VP VP.n84 0.153454
R134 VDD1.n84 VDD1.n0 289.615
R135 VDD1.n175 VDD1.n91 289.615
R136 VDD1.n85 VDD1.n84 185
R137 VDD1.n83 VDD1.n82 185
R138 VDD1.n4 VDD1.n3 185
R139 VDD1.n77 VDD1.n76 185
R140 VDD1.n75 VDD1.n6 185
R141 VDD1.n74 VDD1.n73 185
R142 VDD1.n9 VDD1.n7 185
R143 VDD1.n68 VDD1.n67 185
R144 VDD1.n66 VDD1.n65 185
R145 VDD1.n13 VDD1.n12 185
R146 VDD1.n60 VDD1.n59 185
R147 VDD1.n58 VDD1.n57 185
R148 VDD1.n17 VDD1.n16 185
R149 VDD1.n52 VDD1.n51 185
R150 VDD1.n50 VDD1.n49 185
R151 VDD1.n21 VDD1.n20 185
R152 VDD1.n44 VDD1.n43 185
R153 VDD1.n42 VDD1.n41 185
R154 VDD1.n25 VDD1.n24 185
R155 VDD1.n36 VDD1.n35 185
R156 VDD1.n34 VDD1.n33 185
R157 VDD1.n29 VDD1.n28 185
R158 VDD1.n119 VDD1.n118 185
R159 VDD1.n124 VDD1.n123 185
R160 VDD1.n126 VDD1.n125 185
R161 VDD1.n115 VDD1.n114 185
R162 VDD1.n132 VDD1.n131 185
R163 VDD1.n134 VDD1.n133 185
R164 VDD1.n111 VDD1.n110 185
R165 VDD1.n140 VDD1.n139 185
R166 VDD1.n142 VDD1.n141 185
R167 VDD1.n107 VDD1.n106 185
R168 VDD1.n148 VDD1.n147 185
R169 VDD1.n150 VDD1.n149 185
R170 VDD1.n103 VDD1.n102 185
R171 VDD1.n156 VDD1.n155 185
R172 VDD1.n158 VDD1.n157 185
R173 VDD1.n99 VDD1.n98 185
R174 VDD1.n165 VDD1.n164 185
R175 VDD1.n166 VDD1.n97 185
R176 VDD1.n168 VDD1.n167 185
R177 VDD1.n95 VDD1.n94 185
R178 VDD1.n174 VDD1.n173 185
R179 VDD1.n176 VDD1.n175 185
R180 VDD1.n30 VDD1.t4 147.659
R181 VDD1.n120 VDD1.t9 147.659
R182 VDD1.n84 VDD1.n83 104.615
R183 VDD1.n83 VDD1.n3 104.615
R184 VDD1.n76 VDD1.n3 104.615
R185 VDD1.n76 VDD1.n75 104.615
R186 VDD1.n75 VDD1.n74 104.615
R187 VDD1.n74 VDD1.n7 104.615
R188 VDD1.n67 VDD1.n7 104.615
R189 VDD1.n67 VDD1.n66 104.615
R190 VDD1.n66 VDD1.n12 104.615
R191 VDD1.n59 VDD1.n12 104.615
R192 VDD1.n59 VDD1.n58 104.615
R193 VDD1.n58 VDD1.n16 104.615
R194 VDD1.n51 VDD1.n16 104.615
R195 VDD1.n51 VDD1.n50 104.615
R196 VDD1.n50 VDD1.n20 104.615
R197 VDD1.n43 VDD1.n20 104.615
R198 VDD1.n43 VDD1.n42 104.615
R199 VDD1.n42 VDD1.n24 104.615
R200 VDD1.n35 VDD1.n24 104.615
R201 VDD1.n35 VDD1.n34 104.615
R202 VDD1.n34 VDD1.n28 104.615
R203 VDD1.n124 VDD1.n118 104.615
R204 VDD1.n125 VDD1.n124 104.615
R205 VDD1.n125 VDD1.n114 104.615
R206 VDD1.n132 VDD1.n114 104.615
R207 VDD1.n133 VDD1.n132 104.615
R208 VDD1.n133 VDD1.n110 104.615
R209 VDD1.n140 VDD1.n110 104.615
R210 VDD1.n141 VDD1.n140 104.615
R211 VDD1.n141 VDD1.n106 104.615
R212 VDD1.n148 VDD1.n106 104.615
R213 VDD1.n149 VDD1.n148 104.615
R214 VDD1.n149 VDD1.n102 104.615
R215 VDD1.n156 VDD1.n102 104.615
R216 VDD1.n157 VDD1.n156 104.615
R217 VDD1.n157 VDD1.n98 104.615
R218 VDD1.n165 VDD1.n98 104.615
R219 VDD1.n166 VDD1.n165 104.615
R220 VDD1.n167 VDD1.n166 104.615
R221 VDD1.n167 VDD1.n94 104.615
R222 VDD1.n174 VDD1.n94 104.615
R223 VDD1.n175 VDD1.n174 104.615
R224 VDD1.n183 VDD1.n182 63.0303
R225 VDD1.n90 VDD1.n89 61.3595
R226 VDD1.n185 VDD1.n184 61.3594
R227 VDD1.n181 VDD1.n180 61.3594
R228 VDD1.t4 VDD1.n28 52.3082
R229 VDD1.t9 VDD1.n118 52.3082
R230 VDD1.n90 VDD1.n88 51.7477
R231 VDD1.n181 VDD1.n179 51.7477
R232 VDD1.n185 VDD1.n183 50.2703
R233 VDD1.n30 VDD1.n29 15.6677
R234 VDD1.n120 VDD1.n119 15.6677
R235 VDD1.n77 VDD1.n6 13.1884
R236 VDD1.n168 VDD1.n97 13.1884
R237 VDD1.n78 VDD1.n4 12.8005
R238 VDD1.n73 VDD1.n8 12.8005
R239 VDD1.n33 VDD1.n32 12.8005
R240 VDD1.n123 VDD1.n122 12.8005
R241 VDD1.n164 VDD1.n163 12.8005
R242 VDD1.n169 VDD1.n95 12.8005
R243 VDD1.n82 VDD1.n81 12.0247
R244 VDD1.n72 VDD1.n9 12.0247
R245 VDD1.n36 VDD1.n27 12.0247
R246 VDD1.n126 VDD1.n117 12.0247
R247 VDD1.n162 VDD1.n99 12.0247
R248 VDD1.n173 VDD1.n172 12.0247
R249 VDD1.n85 VDD1.n2 11.249
R250 VDD1.n69 VDD1.n68 11.249
R251 VDD1.n37 VDD1.n25 11.249
R252 VDD1.n127 VDD1.n115 11.249
R253 VDD1.n159 VDD1.n158 11.249
R254 VDD1.n176 VDD1.n93 11.249
R255 VDD1.n86 VDD1.n0 10.4732
R256 VDD1.n65 VDD1.n11 10.4732
R257 VDD1.n41 VDD1.n40 10.4732
R258 VDD1.n131 VDD1.n130 10.4732
R259 VDD1.n155 VDD1.n101 10.4732
R260 VDD1.n177 VDD1.n91 10.4732
R261 VDD1.n64 VDD1.n13 9.69747
R262 VDD1.n44 VDD1.n23 9.69747
R263 VDD1.n134 VDD1.n113 9.69747
R264 VDD1.n154 VDD1.n103 9.69747
R265 VDD1.n88 VDD1.n87 9.45567
R266 VDD1.n179 VDD1.n178 9.45567
R267 VDD1.n56 VDD1.n55 9.3005
R268 VDD1.n15 VDD1.n14 9.3005
R269 VDD1.n62 VDD1.n61 9.3005
R270 VDD1.n64 VDD1.n63 9.3005
R271 VDD1.n11 VDD1.n10 9.3005
R272 VDD1.n70 VDD1.n69 9.3005
R273 VDD1.n72 VDD1.n71 9.3005
R274 VDD1.n8 VDD1.n5 9.3005
R275 VDD1.n87 VDD1.n86 9.3005
R276 VDD1.n2 VDD1.n1 9.3005
R277 VDD1.n81 VDD1.n80 9.3005
R278 VDD1.n79 VDD1.n78 9.3005
R279 VDD1.n54 VDD1.n53 9.3005
R280 VDD1.n19 VDD1.n18 9.3005
R281 VDD1.n48 VDD1.n47 9.3005
R282 VDD1.n46 VDD1.n45 9.3005
R283 VDD1.n23 VDD1.n22 9.3005
R284 VDD1.n40 VDD1.n39 9.3005
R285 VDD1.n38 VDD1.n37 9.3005
R286 VDD1.n27 VDD1.n26 9.3005
R287 VDD1.n32 VDD1.n31 9.3005
R288 VDD1.n178 VDD1.n177 9.3005
R289 VDD1.n93 VDD1.n92 9.3005
R290 VDD1.n172 VDD1.n171 9.3005
R291 VDD1.n170 VDD1.n169 9.3005
R292 VDD1.n109 VDD1.n108 9.3005
R293 VDD1.n138 VDD1.n137 9.3005
R294 VDD1.n136 VDD1.n135 9.3005
R295 VDD1.n113 VDD1.n112 9.3005
R296 VDD1.n130 VDD1.n129 9.3005
R297 VDD1.n128 VDD1.n127 9.3005
R298 VDD1.n117 VDD1.n116 9.3005
R299 VDD1.n122 VDD1.n121 9.3005
R300 VDD1.n144 VDD1.n143 9.3005
R301 VDD1.n146 VDD1.n145 9.3005
R302 VDD1.n105 VDD1.n104 9.3005
R303 VDD1.n152 VDD1.n151 9.3005
R304 VDD1.n154 VDD1.n153 9.3005
R305 VDD1.n101 VDD1.n100 9.3005
R306 VDD1.n160 VDD1.n159 9.3005
R307 VDD1.n162 VDD1.n161 9.3005
R308 VDD1.n163 VDD1.n96 9.3005
R309 VDD1.n61 VDD1.n60 8.92171
R310 VDD1.n45 VDD1.n21 8.92171
R311 VDD1.n135 VDD1.n111 8.92171
R312 VDD1.n151 VDD1.n150 8.92171
R313 VDD1.n57 VDD1.n15 8.14595
R314 VDD1.n49 VDD1.n48 8.14595
R315 VDD1.n139 VDD1.n138 8.14595
R316 VDD1.n147 VDD1.n105 8.14595
R317 VDD1.n56 VDD1.n17 7.3702
R318 VDD1.n52 VDD1.n19 7.3702
R319 VDD1.n142 VDD1.n109 7.3702
R320 VDD1.n146 VDD1.n107 7.3702
R321 VDD1.n53 VDD1.n17 6.59444
R322 VDD1.n53 VDD1.n52 6.59444
R323 VDD1.n143 VDD1.n142 6.59444
R324 VDD1.n143 VDD1.n107 6.59444
R325 VDD1.n57 VDD1.n56 5.81868
R326 VDD1.n49 VDD1.n19 5.81868
R327 VDD1.n139 VDD1.n109 5.81868
R328 VDD1.n147 VDD1.n146 5.81868
R329 VDD1.n60 VDD1.n15 5.04292
R330 VDD1.n48 VDD1.n21 5.04292
R331 VDD1.n138 VDD1.n111 5.04292
R332 VDD1.n150 VDD1.n105 5.04292
R333 VDD1.n31 VDD1.n30 4.38563
R334 VDD1.n121 VDD1.n120 4.38563
R335 VDD1.n61 VDD1.n13 4.26717
R336 VDD1.n45 VDD1.n44 4.26717
R337 VDD1.n135 VDD1.n134 4.26717
R338 VDD1.n151 VDD1.n103 4.26717
R339 VDD1.n88 VDD1.n0 3.49141
R340 VDD1.n65 VDD1.n64 3.49141
R341 VDD1.n41 VDD1.n23 3.49141
R342 VDD1.n131 VDD1.n113 3.49141
R343 VDD1.n155 VDD1.n154 3.49141
R344 VDD1.n179 VDD1.n91 3.49141
R345 VDD1.n86 VDD1.n85 2.71565
R346 VDD1.n68 VDD1.n11 2.71565
R347 VDD1.n40 VDD1.n25 2.71565
R348 VDD1.n130 VDD1.n115 2.71565
R349 VDD1.n158 VDD1.n101 2.71565
R350 VDD1.n177 VDD1.n176 2.71565
R351 VDD1.n82 VDD1.n2 1.93989
R352 VDD1.n69 VDD1.n9 1.93989
R353 VDD1.n37 VDD1.n36 1.93989
R354 VDD1.n127 VDD1.n126 1.93989
R355 VDD1.n159 VDD1.n99 1.93989
R356 VDD1.n173 VDD1.n93 1.93989
R357 VDD1 VDD1.n185 1.6686
R358 VDD1.n184 VDD1.t8 1.22955
R359 VDD1.n184 VDD1.t6 1.22955
R360 VDD1.n89 VDD1.t1 1.22955
R361 VDD1.n89 VDD1.t3 1.22955
R362 VDD1.n182 VDD1.t0 1.22955
R363 VDD1.n182 VDD1.t2 1.22955
R364 VDD1.n180 VDD1.t7 1.22955
R365 VDD1.n180 VDD1.t5 1.22955
R366 VDD1.n81 VDD1.n4 1.16414
R367 VDD1.n73 VDD1.n72 1.16414
R368 VDD1.n33 VDD1.n27 1.16414
R369 VDD1.n123 VDD1.n117 1.16414
R370 VDD1.n164 VDD1.n162 1.16414
R371 VDD1.n172 VDD1.n95 1.16414
R372 VDD1 VDD1.n90 0.634121
R373 VDD1.n183 VDD1.n181 0.520585
R374 VDD1.n78 VDD1.n77 0.388379
R375 VDD1.n8 VDD1.n6 0.388379
R376 VDD1.n32 VDD1.n29 0.388379
R377 VDD1.n122 VDD1.n119 0.388379
R378 VDD1.n163 VDD1.n97 0.388379
R379 VDD1.n169 VDD1.n168 0.388379
R380 VDD1.n87 VDD1.n1 0.155672
R381 VDD1.n80 VDD1.n1 0.155672
R382 VDD1.n80 VDD1.n79 0.155672
R383 VDD1.n79 VDD1.n5 0.155672
R384 VDD1.n71 VDD1.n5 0.155672
R385 VDD1.n71 VDD1.n70 0.155672
R386 VDD1.n70 VDD1.n10 0.155672
R387 VDD1.n63 VDD1.n10 0.155672
R388 VDD1.n63 VDD1.n62 0.155672
R389 VDD1.n62 VDD1.n14 0.155672
R390 VDD1.n55 VDD1.n14 0.155672
R391 VDD1.n55 VDD1.n54 0.155672
R392 VDD1.n54 VDD1.n18 0.155672
R393 VDD1.n47 VDD1.n18 0.155672
R394 VDD1.n47 VDD1.n46 0.155672
R395 VDD1.n46 VDD1.n22 0.155672
R396 VDD1.n39 VDD1.n22 0.155672
R397 VDD1.n39 VDD1.n38 0.155672
R398 VDD1.n38 VDD1.n26 0.155672
R399 VDD1.n31 VDD1.n26 0.155672
R400 VDD1.n121 VDD1.n116 0.155672
R401 VDD1.n128 VDD1.n116 0.155672
R402 VDD1.n129 VDD1.n128 0.155672
R403 VDD1.n129 VDD1.n112 0.155672
R404 VDD1.n136 VDD1.n112 0.155672
R405 VDD1.n137 VDD1.n136 0.155672
R406 VDD1.n137 VDD1.n108 0.155672
R407 VDD1.n144 VDD1.n108 0.155672
R408 VDD1.n145 VDD1.n144 0.155672
R409 VDD1.n145 VDD1.n104 0.155672
R410 VDD1.n152 VDD1.n104 0.155672
R411 VDD1.n153 VDD1.n152 0.155672
R412 VDD1.n153 VDD1.n100 0.155672
R413 VDD1.n160 VDD1.n100 0.155672
R414 VDD1.n161 VDD1.n160 0.155672
R415 VDD1.n161 VDD1.n96 0.155672
R416 VDD1.n170 VDD1.n96 0.155672
R417 VDD1.n171 VDD1.n170 0.155672
R418 VDD1.n171 VDD1.n92 0.155672
R419 VDD1.n178 VDD1.n92 0.155672
R420 VTAIL.n368 VTAIL.n284 289.615
R421 VTAIL.n86 VTAIL.n2 289.615
R422 VTAIL.n278 VTAIL.n194 289.615
R423 VTAIL.n184 VTAIL.n100 289.615
R424 VTAIL.n312 VTAIL.n311 185
R425 VTAIL.n317 VTAIL.n316 185
R426 VTAIL.n319 VTAIL.n318 185
R427 VTAIL.n308 VTAIL.n307 185
R428 VTAIL.n325 VTAIL.n324 185
R429 VTAIL.n327 VTAIL.n326 185
R430 VTAIL.n304 VTAIL.n303 185
R431 VTAIL.n333 VTAIL.n332 185
R432 VTAIL.n335 VTAIL.n334 185
R433 VTAIL.n300 VTAIL.n299 185
R434 VTAIL.n341 VTAIL.n340 185
R435 VTAIL.n343 VTAIL.n342 185
R436 VTAIL.n296 VTAIL.n295 185
R437 VTAIL.n349 VTAIL.n348 185
R438 VTAIL.n351 VTAIL.n350 185
R439 VTAIL.n292 VTAIL.n291 185
R440 VTAIL.n358 VTAIL.n357 185
R441 VTAIL.n359 VTAIL.n290 185
R442 VTAIL.n361 VTAIL.n360 185
R443 VTAIL.n288 VTAIL.n287 185
R444 VTAIL.n367 VTAIL.n366 185
R445 VTAIL.n369 VTAIL.n368 185
R446 VTAIL.n30 VTAIL.n29 185
R447 VTAIL.n35 VTAIL.n34 185
R448 VTAIL.n37 VTAIL.n36 185
R449 VTAIL.n26 VTAIL.n25 185
R450 VTAIL.n43 VTAIL.n42 185
R451 VTAIL.n45 VTAIL.n44 185
R452 VTAIL.n22 VTAIL.n21 185
R453 VTAIL.n51 VTAIL.n50 185
R454 VTAIL.n53 VTAIL.n52 185
R455 VTAIL.n18 VTAIL.n17 185
R456 VTAIL.n59 VTAIL.n58 185
R457 VTAIL.n61 VTAIL.n60 185
R458 VTAIL.n14 VTAIL.n13 185
R459 VTAIL.n67 VTAIL.n66 185
R460 VTAIL.n69 VTAIL.n68 185
R461 VTAIL.n10 VTAIL.n9 185
R462 VTAIL.n76 VTAIL.n75 185
R463 VTAIL.n77 VTAIL.n8 185
R464 VTAIL.n79 VTAIL.n78 185
R465 VTAIL.n6 VTAIL.n5 185
R466 VTAIL.n85 VTAIL.n84 185
R467 VTAIL.n87 VTAIL.n86 185
R468 VTAIL.n279 VTAIL.n278 185
R469 VTAIL.n277 VTAIL.n276 185
R470 VTAIL.n198 VTAIL.n197 185
R471 VTAIL.n271 VTAIL.n270 185
R472 VTAIL.n269 VTAIL.n200 185
R473 VTAIL.n268 VTAIL.n267 185
R474 VTAIL.n203 VTAIL.n201 185
R475 VTAIL.n262 VTAIL.n261 185
R476 VTAIL.n260 VTAIL.n259 185
R477 VTAIL.n207 VTAIL.n206 185
R478 VTAIL.n254 VTAIL.n253 185
R479 VTAIL.n252 VTAIL.n251 185
R480 VTAIL.n211 VTAIL.n210 185
R481 VTAIL.n246 VTAIL.n245 185
R482 VTAIL.n244 VTAIL.n243 185
R483 VTAIL.n215 VTAIL.n214 185
R484 VTAIL.n238 VTAIL.n237 185
R485 VTAIL.n236 VTAIL.n235 185
R486 VTAIL.n219 VTAIL.n218 185
R487 VTAIL.n230 VTAIL.n229 185
R488 VTAIL.n228 VTAIL.n227 185
R489 VTAIL.n223 VTAIL.n222 185
R490 VTAIL.n185 VTAIL.n184 185
R491 VTAIL.n183 VTAIL.n182 185
R492 VTAIL.n104 VTAIL.n103 185
R493 VTAIL.n177 VTAIL.n176 185
R494 VTAIL.n175 VTAIL.n106 185
R495 VTAIL.n174 VTAIL.n173 185
R496 VTAIL.n109 VTAIL.n107 185
R497 VTAIL.n168 VTAIL.n167 185
R498 VTAIL.n166 VTAIL.n165 185
R499 VTAIL.n113 VTAIL.n112 185
R500 VTAIL.n160 VTAIL.n159 185
R501 VTAIL.n158 VTAIL.n157 185
R502 VTAIL.n117 VTAIL.n116 185
R503 VTAIL.n152 VTAIL.n151 185
R504 VTAIL.n150 VTAIL.n149 185
R505 VTAIL.n121 VTAIL.n120 185
R506 VTAIL.n144 VTAIL.n143 185
R507 VTAIL.n142 VTAIL.n141 185
R508 VTAIL.n125 VTAIL.n124 185
R509 VTAIL.n136 VTAIL.n135 185
R510 VTAIL.n134 VTAIL.n133 185
R511 VTAIL.n129 VTAIL.n128 185
R512 VTAIL.n313 VTAIL.t8 147.659
R513 VTAIL.n31 VTAIL.t16 147.659
R514 VTAIL.n224 VTAIL.t18 147.659
R515 VTAIL.n130 VTAIL.t6 147.659
R516 VTAIL.n317 VTAIL.n311 104.615
R517 VTAIL.n318 VTAIL.n317 104.615
R518 VTAIL.n318 VTAIL.n307 104.615
R519 VTAIL.n325 VTAIL.n307 104.615
R520 VTAIL.n326 VTAIL.n325 104.615
R521 VTAIL.n326 VTAIL.n303 104.615
R522 VTAIL.n333 VTAIL.n303 104.615
R523 VTAIL.n334 VTAIL.n333 104.615
R524 VTAIL.n334 VTAIL.n299 104.615
R525 VTAIL.n341 VTAIL.n299 104.615
R526 VTAIL.n342 VTAIL.n341 104.615
R527 VTAIL.n342 VTAIL.n295 104.615
R528 VTAIL.n349 VTAIL.n295 104.615
R529 VTAIL.n350 VTAIL.n349 104.615
R530 VTAIL.n350 VTAIL.n291 104.615
R531 VTAIL.n358 VTAIL.n291 104.615
R532 VTAIL.n359 VTAIL.n358 104.615
R533 VTAIL.n360 VTAIL.n359 104.615
R534 VTAIL.n360 VTAIL.n287 104.615
R535 VTAIL.n367 VTAIL.n287 104.615
R536 VTAIL.n368 VTAIL.n367 104.615
R537 VTAIL.n35 VTAIL.n29 104.615
R538 VTAIL.n36 VTAIL.n35 104.615
R539 VTAIL.n36 VTAIL.n25 104.615
R540 VTAIL.n43 VTAIL.n25 104.615
R541 VTAIL.n44 VTAIL.n43 104.615
R542 VTAIL.n44 VTAIL.n21 104.615
R543 VTAIL.n51 VTAIL.n21 104.615
R544 VTAIL.n52 VTAIL.n51 104.615
R545 VTAIL.n52 VTAIL.n17 104.615
R546 VTAIL.n59 VTAIL.n17 104.615
R547 VTAIL.n60 VTAIL.n59 104.615
R548 VTAIL.n60 VTAIL.n13 104.615
R549 VTAIL.n67 VTAIL.n13 104.615
R550 VTAIL.n68 VTAIL.n67 104.615
R551 VTAIL.n68 VTAIL.n9 104.615
R552 VTAIL.n76 VTAIL.n9 104.615
R553 VTAIL.n77 VTAIL.n76 104.615
R554 VTAIL.n78 VTAIL.n77 104.615
R555 VTAIL.n78 VTAIL.n5 104.615
R556 VTAIL.n85 VTAIL.n5 104.615
R557 VTAIL.n86 VTAIL.n85 104.615
R558 VTAIL.n278 VTAIL.n277 104.615
R559 VTAIL.n277 VTAIL.n197 104.615
R560 VTAIL.n270 VTAIL.n197 104.615
R561 VTAIL.n270 VTAIL.n269 104.615
R562 VTAIL.n269 VTAIL.n268 104.615
R563 VTAIL.n268 VTAIL.n201 104.615
R564 VTAIL.n261 VTAIL.n201 104.615
R565 VTAIL.n261 VTAIL.n260 104.615
R566 VTAIL.n260 VTAIL.n206 104.615
R567 VTAIL.n253 VTAIL.n206 104.615
R568 VTAIL.n253 VTAIL.n252 104.615
R569 VTAIL.n252 VTAIL.n210 104.615
R570 VTAIL.n245 VTAIL.n210 104.615
R571 VTAIL.n245 VTAIL.n244 104.615
R572 VTAIL.n244 VTAIL.n214 104.615
R573 VTAIL.n237 VTAIL.n214 104.615
R574 VTAIL.n237 VTAIL.n236 104.615
R575 VTAIL.n236 VTAIL.n218 104.615
R576 VTAIL.n229 VTAIL.n218 104.615
R577 VTAIL.n229 VTAIL.n228 104.615
R578 VTAIL.n228 VTAIL.n222 104.615
R579 VTAIL.n184 VTAIL.n183 104.615
R580 VTAIL.n183 VTAIL.n103 104.615
R581 VTAIL.n176 VTAIL.n103 104.615
R582 VTAIL.n176 VTAIL.n175 104.615
R583 VTAIL.n175 VTAIL.n174 104.615
R584 VTAIL.n174 VTAIL.n107 104.615
R585 VTAIL.n167 VTAIL.n107 104.615
R586 VTAIL.n167 VTAIL.n166 104.615
R587 VTAIL.n166 VTAIL.n112 104.615
R588 VTAIL.n159 VTAIL.n112 104.615
R589 VTAIL.n159 VTAIL.n158 104.615
R590 VTAIL.n158 VTAIL.n116 104.615
R591 VTAIL.n151 VTAIL.n116 104.615
R592 VTAIL.n151 VTAIL.n150 104.615
R593 VTAIL.n150 VTAIL.n120 104.615
R594 VTAIL.n143 VTAIL.n120 104.615
R595 VTAIL.n143 VTAIL.n142 104.615
R596 VTAIL.n142 VTAIL.n124 104.615
R597 VTAIL.n135 VTAIL.n124 104.615
R598 VTAIL.n135 VTAIL.n134 104.615
R599 VTAIL.n134 VTAIL.n128 104.615
R600 VTAIL.t8 VTAIL.n311 52.3082
R601 VTAIL.t16 VTAIL.n29 52.3082
R602 VTAIL.t18 VTAIL.n222 52.3082
R603 VTAIL.t6 VTAIL.n128 52.3082
R604 VTAIL.n193 VTAIL.n192 44.6808
R605 VTAIL.n191 VTAIL.n190 44.6808
R606 VTAIL.n99 VTAIL.n98 44.6808
R607 VTAIL.n97 VTAIL.n96 44.6808
R608 VTAIL.n375 VTAIL.n374 44.6806
R609 VTAIL.n1 VTAIL.n0 44.6806
R610 VTAIL.n93 VTAIL.n92 44.6806
R611 VTAIL.n95 VTAIL.n94 44.6806
R612 VTAIL.n373 VTAIL.n372 32.7672
R613 VTAIL.n91 VTAIL.n90 32.7672
R614 VTAIL.n283 VTAIL.n282 32.7672
R615 VTAIL.n189 VTAIL.n188 32.7672
R616 VTAIL.n97 VTAIL.n95 30.8583
R617 VTAIL.n373 VTAIL.n283 28.5565
R618 VTAIL.n313 VTAIL.n312 15.6677
R619 VTAIL.n31 VTAIL.n30 15.6677
R620 VTAIL.n224 VTAIL.n223 15.6677
R621 VTAIL.n130 VTAIL.n129 15.6677
R622 VTAIL.n361 VTAIL.n290 13.1884
R623 VTAIL.n79 VTAIL.n8 13.1884
R624 VTAIL.n271 VTAIL.n200 13.1884
R625 VTAIL.n177 VTAIL.n106 13.1884
R626 VTAIL.n316 VTAIL.n315 12.8005
R627 VTAIL.n357 VTAIL.n356 12.8005
R628 VTAIL.n362 VTAIL.n288 12.8005
R629 VTAIL.n34 VTAIL.n33 12.8005
R630 VTAIL.n75 VTAIL.n74 12.8005
R631 VTAIL.n80 VTAIL.n6 12.8005
R632 VTAIL.n272 VTAIL.n198 12.8005
R633 VTAIL.n267 VTAIL.n202 12.8005
R634 VTAIL.n227 VTAIL.n226 12.8005
R635 VTAIL.n178 VTAIL.n104 12.8005
R636 VTAIL.n173 VTAIL.n108 12.8005
R637 VTAIL.n133 VTAIL.n132 12.8005
R638 VTAIL.n319 VTAIL.n310 12.0247
R639 VTAIL.n355 VTAIL.n292 12.0247
R640 VTAIL.n366 VTAIL.n365 12.0247
R641 VTAIL.n37 VTAIL.n28 12.0247
R642 VTAIL.n73 VTAIL.n10 12.0247
R643 VTAIL.n84 VTAIL.n83 12.0247
R644 VTAIL.n276 VTAIL.n275 12.0247
R645 VTAIL.n266 VTAIL.n203 12.0247
R646 VTAIL.n230 VTAIL.n221 12.0247
R647 VTAIL.n182 VTAIL.n181 12.0247
R648 VTAIL.n172 VTAIL.n109 12.0247
R649 VTAIL.n136 VTAIL.n127 12.0247
R650 VTAIL.n320 VTAIL.n308 11.249
R651 VTAIL.n352 VTAIL.n351 11.249
R652 VTAIL.n369 VTAIL.n286 11.249
R653 VTAIL.n38 VTAIL.n26 11.249
R654 VTAIL.n70 VTAIL.n69 11.249
R655 VTAIL.n87 VTAIL.n4 11.249
R656 VTAIL.n279 VTAIL.n196 11.249
R657 VTAIL.n263 VTAIL.n262 11.249
R658 VTAIL.n231 VTAIL.n219 11.249
R659 VTAIL.n185 VTAIL.n102 11.249
R660 VTAIL.n169 VTAIL.n168 11.249
R661 VTAIL.n137 VTAIL.n125 11.249
R662 VTAIL.n324 VTAIL.n323 10.4732
R663 VTAIL.n348 VTAIL.n294 10.4732
R664 VTAIL.n370 VTAIL.n284 10.4732
R665 VTAIL.n42 VTAIL.n41 10.4732
R666 VTAIL.n66 VTAIL.n12 10.4732
R667 VTAIL.n88 VTAIL.n2 10.4732
R668 VTAIL.n280 VTAIL.n194 10.4732
R669 VTAIL.n259 VTAIL.n205 10.4732
R670 VTAIL.n235 VTAIL.n234 10.4732
R671 VTAIL.n186 VTAIL.n100 10.4732
R672 VTAIL.n165 VTAIL.n111 10.4732
R673 VTAIL.n141 VTAIL.n140 10.4732
R674 VTAIL.n327 VTAIL.n306 9.69747
R675 VTAIL.n347 VTAIL.n296 9.69747
R676 VTAIL.n45 VTAIL.n24 9.69747
R677 VTAIL.n65 VTAIL.n14 9.69747
R678 VTAIL.n258 VTAIL.n207 9.69747
R679 VTAIL.n238 VTAIL.n217 9.69747
R680 VTAIL.n164 VTAIL.n113 9.69747
R681 VTAIL.n144 VTAIL.n123 9.69747
R682 VTAIL.n372 VTAIL.n371 9.45567
R683 VTAIL.n90 VTAIL.n89 9.45567
R684 VTAIL.n282 VTAIL.n281 9.45567
R685 VTAIL.n188 VTAIL.n187 9.45567
R686 VTAIL.n371 VTAIL.n370 9.3005
R687 VTAIL.n286 VTAIL.n285 9.3005
R688 VTAIL.n365 VTAIL.n364 9.3005
R689 VTAIL.n363 VTAIL.n362 9.3005
R690 VTAIL.n302 VTAIL.n301 9.3005
R691 VTAIL.n331 VTAIL.n330 9.3005
R692 VTAIL.n329 VTAIL.n328 9.3005
R693 VTAIL.n306 VTAIL.n305 9.3005
R694 VTAIL.n323 VTAIL.n322 9.3005
R695 VTAIL.n321 VTAIL.n320 9.3005
R696 VTAIL.n310 VTAIL.n309 9.3005
R697 VTAIL.n315 VTAIL.n314 9.3005
R698 VTAIL.n337 VTAIL.n336 9.3005
R699 VTAIL.n339 VTAIL.n338 9.3005
R700 VTAIL.n298 VTAIL.n297 9.3005
R701 VTAIL.n345 VTAIL.n344 9.3005
R702 VTAIL.n347 VTAIL.n346 9.3005
R703 VTAIL.n294 VTAIL.n293 9.3005
R704 VTAIL.n353 VTAIL.n352 9.3005
R705 VTAIL.n355 VTAIL.n354 9.3005
R706 VTAIL.n356 VTAIL.n289 9.3005
R707 VTAIL.n89 VTAIL.n88 9.3005
R708 VTAIL.n4 VTAIL.n3 9.3005
R709 VTAIL.n83 VTAIL.n82 9.3005
R710 VTAIL.n81 VTAIL.n80 9.3005
R711 VTAIL.n20 VTAIL.n19 9.3005
R712 VTAIL.n49 VTAIL.n48 9.3005
R713 VTAIL.n47 VTAIL.n46 9.3005
R714 VTAIL.n24 VTAIL.n23 9.3005
R715 VTAIL.n41 VTAIL.n40 9.3005
R716 VTAIL.n39 VTAIL.n38 9.3005
R717 VTAIL.n28 VTAIL.n27 9.3005
R718 VTAIL.n33 VTAIL.n32 9.3005
R719 VTAIL.n55 VTAIL.n54 9.3005
R720 VTAIL.n57 VTAIL.n56 9.3005
R721 VTAIL.n16 VTAIL.n15 9.3005
R722 VTAIL.n63 VTAIL.n62 9.3005
R723 VTAIL.n65 VTAIL.n64 9.3005
R724 VTAIL.n12 VTAIL.n11 9.3005
R725 VTAIL.n71 VTAIL.n70 9.3005
R726 VTAIL.n73 VTAIL.n72 9.3005
R727 VTAIL.n74 VTAIL.n7 9.3005
R728 VTAIL.n250 VTAIL.n249 9.3005
R729 VTAIL.n209 VTAIL.n208 9.3005
R730 VTAIL.n256 VTAIL.n255 9.3005
R731 VTAIL.n258 VTAIL.n257 9.3005
R732 VTAIL.n205 VTAIL.n204 9.3005
R733 VTAIL.n264 VTAIL.n263 9.3005
R734 VTAIL.n266 VTAIL.n265 9.3005
R735 VTAIL.n202 VTAIL.n199 9.3005
R736 VTAIL.n281 VTAIL.n280 9.3005
R737 VTAIL.n196 VTAIL.n195 9.3005
R738 VTAIL.n275 VTAIL.n274 9.3005
R739 VTAIL.n273 VTAIL.n272 9.3005
R740 VTAIL.n248 VTAIL.n247 9.3005
R741 VTAIL.n213 VTAIL.n212 9.3005
R742 VTAIL.n242 VTAIL.n241 9.3005
R743 VTAIL.n240 VTAIL.n239 9.3005
R744 VTAIL.n217 VTAIL.n216 9.3005
R745 VTAIL.n234 VTAIL.n233 9.3005
R746 VTAIL.n232 VTAIL.n231 9.3005
R747 VTAIL.n221 VTAIL.n220 9.3005
R748 VTAIL.n226 VTAIL.n225 9.3005
R749 VTAIL.n156 VTAIL.n155 9.3005
R750 VTAIL.n115 VTAIL.n114 9.3005
R751 VTAIL.n162 VTAIL.n161 9.3005
R752 VTAIL.n164 VTAIL.n163 9.3005
R753 VTAIL.n111 VTAIL.n110 9.3005
R754 VTAIL.n170 VTAIL.n169 9.3005
R755 VTAIL.n172 VTAIL.n171 9.3005
R756 VTAIL.n108 VTAIL.n105 9.3005
R757 VTAIL.n187 VTAIL.n186 9.3005
R758 VTAIL.n102 VTAIL.n101 9.3005
R759 VTAIL.n181 VTAIL.n180 9.3005
R760 VTAIL.n179 VTAIL.n178 9.3005
R761 VTAIL.n154 VTAIL.n153 9.3005
R762 VTAIL.n119 VTAIL.n118 9.3005
R763 VTAIL.n148 VTAIL.n147 9.3005
R764 VTAIL.n146 VTAIL.n145 9.3005
R765 VTAIL.n123 VTAIL.n122 9.3005
R766 VTAIL.n140 VTAIL.n139 9.3005
R767 VTAIL.n138 VTAIL.n137 9.3005
R768 VTAIL.n127 VTAIL.n126 9.3005
R769 VTAIL.n132 VTAIL.n131 9.3005
R770 VTAIL.n328 VTAIL.n304 8.92171
R771 VTAIL.n344 VTAIL.n343 8.92171
R772 VTAIL.n46 VTAIL.n22 8.92171
R773 VTAIL.n62 VTAIL.n61 8.92171
R774 VTAIL.n255 VTAIL.n254 8.92171
R775 VTAIL.n239 VTAIL.n215 8.92171
R776 VTAIL.n161 VTAIL.n160 8.92171
R777 VTAIL.n145 VTAIL.n121 8.92171
R778 VTAIL.n332 VTAIL.n331 8.14595
R779 VTAIL.n340 VTAIL.n298 8.14595
R780 VTAIL.n50 VTAIL.n49 8.14595
R781 VTAIL.n58 VTAIL.n16 8.14595
R782 VTAIL.n251 VTAIL.n209 8.14595
R783 VTAIL.n243 VTAIL.n242 8.14595
R784 VTAIL.n157 VTAIL.n115 8.14595
R785 VTAIL.n149 VTAIL.n148 8.14595
R786 VTAIL.n335 VTAIL.n302 7.3702
R787 VTAIL.n339 VTAIL.n300 7.3702
R788 VTAIL.n53 VTAIL.n20 7.3702
R789 VTAIL.n57 VTAIL.n18 7.3702
R790 VTAIL.n250 VTAIL.n211 7.3702
R791 VTAIL.n246 VTAIL.n213 7.3702
R792 VTAIL.n156 VTAIL.n117 7.3702
R793 VTAIL.n152 VTAIL.n119 7.3702
R794 VTAIL.n336 VTAIL.n335 6.59444
R795 VTAIL.n336 VTAIL.n300 6.59444
R796 VTAIL.n54 VTAIL.n53 6.59444
R797 VTAIL.n54 VTAIL.n18 6.59444
R798 VTAIL.n247 VTAIL.n211 6.59444
R799 VTAIL.n247 VTAIL.n246 6.59444
R800 VTAIL.n153 VTAIL.n117 6.59444
R801 VTAIL.n153 VTAIL.n152 6.59444
R802 VTAIL.n332 VTAIL.n302 5.81868
R803 VTAIL.n340 VTAIL.n339 5.81868
R804 VTAIL.n50 VTAIL.n20 5.81868
R805 VTAIL.n58 VTAIL.n57 5.81868
R806 VTAIL.n251 VTAIL.n250 5.81868
R807 VTAIL.n243 VTAIL.n213 5.81868
R808 VTAIL.n157 VTAIL.n156 5.81868
R809 VTAIL.n149 VTAIL.n119 5.81868
R810 VTAIL.n331 VTAIL.n304 5.04292
R811 VTAIL.n343 VTAIL.n298 5.04292
R812 VTAIL.n49 VTAIL.n22 5.04292
R813 VTAIL.n61 VTAIL.n16 5.04292
R814 VTAIL.n254 VTAIL.n209 5.04292
R815 VTAIL.n242 VTAIL.n215 5.04292
R816 VTAIL.n160 VTAIL.n115 5.04292
R817 VTAIL.n148 VTAIL.n121 5.04292
R818 VTAIL.n314 VTAIL.n313 4.38563
R819 VTAIL.n32 VTAIL.n31 4.38563
R820 VTAIL.n225 VTAIL.n224 4.38563
R821 VTAIL.n131 VTAIL.n130 4.38563
R822 VTAIL.n328 VTAIL.n327 4.26717
R823 VTAIL.n344 VTAIL.n296 4.26717
R824 VTAIL.n46 VTAIL.n45 4.26717
R825 VTAIL.n62 VTAIL.n14 4.26717
R826 VTAIL.n255 VTAIL.n207 4.26717
R827 VTAIL.n239 VTAIL.n238 4.26717
R828 VTAIL.n161 VTAIL.n113 4.26717
R829 VTAIL.n145 VTAIL.n144 4.26717
R830 VTAIL.n324 VTAIL.n306 3.49141
R831 VTAIL.n348 VTAIL.n347 3.49141
R832 VTAIL.n372 VTAIL.n284 3.49141
R833 VTAIL.n42 VTAIL.n24 3.49141
R834 VTAIL.n66 VTAIL.n65 3.49141
R835 VTAIL.n90 VTAIL.n2 3.49141
R836 VTAIL.n282 VTAIL.n194 3.49141
R837 VTAIL.n259 VTAIL.n258 3.49141
R838 VTAIL.n235 VTAIL.n217 3.49141
R839 VTAIL.n188 VTAIL.n100 3.49141
R840 VTAIL.n165 VTAIL.n164 3.49141
R841 VTAIL.n141 VTAIL.n123 3.49141
R842 VTAIL.n323 VTAIL.n308 2.71565
R843 VTAIL.n351 VTAIL.n294 2.71565
R844 VTAIL.n370 VTAIL.n369 2.71565
R845 VTAIL.n41 VTAIL.n26 2.71565
R846 VTAIL.n69 VTAIL.n12 2.71565
R847 VTAIL.n88 VTAIL.n87 2.71565
R848 VTAIL.n280 VTAIL.n279 2.71565
R849 VTAIL.n262 VTAIL.n205 2.71565
R850 VTAIL.n234 VTAIL.n219 2.71565
R851 VTAIL.n186 VTAIL.n185 2.71565
R852 VTAIL.n168 VTAIL.n111 2.71565
R853 VTAIL.n140 VTAIL.n125 2.71565
R854 VTAIL.n99 VTAIL.n97 2.30222
R855 VTAIL.n189 VTAIL.n99 2.30222
R856 VTAIL.n193 VTAIL.n191 2.30222
R857 VTAIL.n283 VTAIL.n193 2.30222
R858 VTAIL.n95 VTAIL.n93 2.30222
R859 VTAIL.n93 VTAIL.n91 2.30222
R860 VTAIL.n375 VTAIL.n373 2.30222
R861 VTAIL.n320 VTAIL.n319 1.93989
R862 VTAIL.n352 VTAIL.n292 1.93989
R863 VTAIL.n366 VTAIL.n286 1.93989
R864 VTAIL.n38 VTAIL.n37 1.93989
R865 VTAIL.n70 VTAIL.n10 1.93989
R866 VTAIL.n84 VTAIL.n4 1.93989
R867 VTAIL.n276 VTAIL.n196 1.93989
R868 VTAIL.n263 VTAIL.n203 1.93989
R869 VTAIL.n231 VTAIL.n230 1.93989
R870 VTAIL.n182 VTAIL.n102 1.93989
R871 VTAIL.n169 VTAIL.n109 1.93989
R872 VTAIL.n137 VTAIL.n136 1.93989
R873 VTAIL VTAIL.n1 1.78498
R874 VTAIL.n191 VTAIL.n189 1.62119
R875 VTAIL.n91 VTAIL.n1 1.62119
R876 VTAIL.n374 VTAIL.t7 1.22955
R877 VTAIL.n374 VTAIL.t5 1.22955
R878 VTAIL.n0 VTAIL.t1 1.22955
R879 VTAIL.n0 VTAIL.t0 1.22955
R880 VTAIL.n92 VTAIL.t15 1.22955
R881 VTAIL.n92 VTAIL.t10 1.22955
R882 VTAIL.n94 VTAIL.t13 1.22955
R883 VTAIL.n94 VTAIL.t19 1.22955
R884 VTAIL.n192 VTAIL.t17 1.22955
R885 VTAIL.n192 VTAIL.t12 1.22955
R886 VTAIL.n190 VTAIL.t14 1.22955
R887 VTAIL.n190 VTAIL.t11 1.22955
R888 VTAIL.n98 VTAIL.t3 1.22955
R889 VTAIL.n98 VTAIL.t4 1.22955
R890 VTAIL.n96 VTAIL.t2 1.22955
R891 VTAIL.n96 VTAIL.t9 1.22955
R892 VTAIL.n316 VTAIL.n310 1.16414
R893 VTAIL.n357 VTAIL.n355 1.16414
R894 VTAIL.n365 VTAIL.n288 1.16414
R895 VTAIL.n34 VTAIL.n28 1.16414
R896 VTAIL.n75 VTAIL.n73 1.16414
R897 VTAIL.n83 VTAIL.n6 1.16414
R898 VTAIL.n275 VTAIL.n198 1.16414
R899 VTAIL.n267 VTAIL.n266 1.16414
R900 VTAIL.n227 VTAIL.n221 1.16414
R901 VTAIL.n181 VTAIL.n104 1.16414
R902 VTAIL.n173 VTAIL.n172 1.16414
R903 VTAIL.n133 VTAIL.n127 1.16414
R904 VTAIL VTAIL.n375 0.517741
R905 VTAIL.n315 VTAIL.n312 0.388379
R906 VTAIL.n356 VTAIL.n290 0.388379
R907 VTAIL.n362 VTAIL.n361 0.388379
R908 VTAIL.n33 VTAIL.n30 0.388379
R909 VTAIL.n74 VTAIL.n8 0.388379
R910 VTAIL.n80 VTAIL.n79 0.388379
R911 VTAIL.n272 VTAIL.n271 0.388379
R912 VTAIL.n202 VTAIL.n200 0.388379
R913 VTAIL.n226 VTAIL.n223 0.388379
R914 VTAIL.n178 VTAIL.n177 0.388379
R915 VTAIL.n108 VTAIL.n106 0.388379
R916 VTAIL.n132 VTAIL.n129 0.388379
R917 VTAIL.n314 VTAIL.n309 0.155672
R918 VTAIL.n321 VTAIL.n309 0.155672
R919 VTAIL.n322 VTAIL.n321 0.155672
R920 VTAIL.n322 VTAIL.n305 0.155672
R921 VTAIL.n329 VTAIL.n305 0.155672
R922 VTAIL.n330 VTAIL.n329 0.155672
R923 VTAIL.n330 VTAIL.n301 0.155672
R924 VTAIL.n337 VTAIL.n301 0.155672
R925 VTAIL.n338 VTAIL.n337 0.155672
R926 VTAIL.n338 VTAIL.n297 0.155672
R927 VTAIL.n345 VTAIL.n297 0.155672
R928 VTAIL.n346 VTAIL.n345 0.155672
R929 VTAIL.n346 VTAIL.n293 0.155672
R930 VTAIL.n353 VTAIL.n293 0.155672
R931 VTAIL.n354 VTAIL.n353 0.155672
R932 VTAIL.n354 VTAIL.n289 0.155672
R933 VTAIL.n363 VTAIL.n289 0.155672
R934 VTAIL.n364 VTAIL.n363 0.155672
R935 VTAIL.n364 VTAIL.n285 0.155672
R936 VTAIL.n371 VTAIL.n285 0.155672
R937 VTAIL.n32 VTAIL.n27 0.155672
R938 VTAIL.n39 VTAIL.n27 0.155672
R939 VTAIL.n40 VTAIL.n39 0.155672
R940 VTAIL.n40 VTAIL.n23 0.155672
R941 VTAIL.n47 VTAIL.n23 0.155672
R942 VTAIL.n48 VTAIL.n47 0.155672
R943 VTAIL.n48 VTAIL.n19 0.155672
R944 VTAIL.n55 VTAIL.n19 0.155672
R945 VTAIL.n56 VTAIL.n55 0.155672
R946 VTAIL.n56 VTAIL.n15 0.155672
R947 VTAIL.n63 VTAIL.n15 0.155672
R948 VTAIL.n64 VTAIL.n63 0.155672
R949 VTAIL.n64 VTAIL.n11 0.155672
R950 VTAIL.n71 VTAIL.n11 0.155672
R951 VTAIL.n72 VTAIL.n71 0.155672
R952 VTAIL.n72 VTAIL.n7 0.155672
R953 VTAIL.n81 VTAIL.n7 0.155672
R954 VTAIL.n82 VTAIL.n81 0.155672
R955 VTAIL.n82 VTAIL.n3 0.155672
R956 VTAIL.n89 VTAIL.n3 0.155672
R957 VTAIL.n281 VTAIL.n195 0.155672
R958 VTAIL.n274 VTAIL.n195 0.155672
R959 VTAIL.n274 VTAIL.n273 0.155672
R960 VTAIL.n273 VTAIL.n199 0.155672
R961 VTAIL.n265 VTAIL.n199 0.155672
R962 VTAIL.n265 VTAIL.n264 0.155672
R963 VTAIL.n264 VTAIL.n204 0.155672
R964 VTAIL.n257 VTAIL.n204 0.155672
R965 VTAIL.n257 VTAIL.n256 0.155672
R966 VTAIL.n256 VTAIL.n208 0.155672
R967 VTAIL.n249 VTAIL.n208 0.155672
R968 VTAIL.n249 VTAIL.n248 0.155672
R969 VTAIL.n248 VTAIL.n212 0.155672
R970 VTAIL.n241 VTAIL.n212 0.155672
R971 VTAIL.n241 VTAIL.n240 0.155672
R972 VTAIL.n240 VTAIL.n216 0.155672
R973 VTAIL.n233 VTAIL.n216 0.155672
R974 VTAIL.n233 VTAIL.n232 0.155672
R975 VTAIL.n232 VTAIL.n220 0.155672
R976 VTAIL.n225 VTAIL.n220 0.155672
R977 VTAIL.n187 VTAIL.n101 0.155672
R978 VTAIL.n180 VTAIL.n101 0.155672
R979 VTAIL.n180 VTAIL.n179 0.155672
R980 VTAIL.n179 VTAIL.n105 0.155672
R981 VTAIL.n171 VTAIL.n105 0.155672
R982 VTAIL.n171 VTAIL.n170 0.155672
R983 VTAIL.n170 VTAIL.n110 0.155672
R984 VTAIL.n163 VTAIL.n110 0.155672
R985 VTAIL.n163 VTAIL.n162 0.155672
R986 VTAIL.n162 VTAIL.n114 0.155672
R987 VTAIL.n155 VTAIL.n114 0.155672
R988 VTAIL.n155 VTAIL.n154 0.155672
R989 VTAIL.n154 VTAIL.n118 0.155672
R990 VTAIL.n147 VTAIL.n118 0.155672
R991 VTAIL.n147 VTAIL.n146 0.155672
R992 VTAIL.n146 VTAIL.n122 0.155672
R993 VTAIL.n139 VTAIL.n122 0.155672
R994 VTAIL.n139 VTAIL.n138 0.155672
R995 VTAIL.n138 VTAIL.n126 0.155672
R996 VTAIL.n131 VTAIL.n126 0.155672
R997 B.n1035 B.n1034 585
R998 B.n1036 B.n1035 585
R999 B.n394 B.n160 585
R1000 B.n393 B.n392 585
R1001 B.n391 B.n390 585
R1002 B.n389 B.n388 585
R1003 B.n387 B.n386 585
R1004 B.n385 B.n384 585
R1005 B.n383 B.n382 585
R1006 B.n381 B.n380 585
R1007 B.n379 B.n378 585
R1008 B.n377 B.n376 585
R1009 B.n375 B.n374 585
R1010 B.n373 B.n372 585
R1011 B.n371 B.n370 585
R1012 B.n369 B.n368 585
R1013 B.n367 B.n366 585
R1014 B.n365 B.n364 585
R1015 B.n363 B.n362 585
R1016 B.n361 B.n360 585
R1017 B.n359 B.n358 585
R1018 B.n357 B.n356 585
R1019 B.n355 B.n354 585
R1020 B.n353 B.n352 585
R1021 B.n351 B.n350 585
R1022 B.n349 B.n348 585
R1023 B.n347 B.n346 585
R1024 B.n345 B.n344 585
R1025 B.n343 B.n342 585
R1026 B.n341 B.n340 585
R1027 B.n339 B.n338 585
R1028 B.n337 B.n336 585
R1029 B.n335 B.n334 585
R1030 B.n333 B.n332 585
R1031 B.n331 B.n330 585
R1032 B.n329 B.n328 585
R1033 B.n327 B.n326 585
R1034 B.n325 B.n324 585
R1035 B.n323 B.n322 585
R1036 B.n321 B.n320 585
R1037 B.n319 B.n318 585
R1038 B.n317 B.n316 585
R1039 B.n315 B.n314 585
R1040 B.n313 B.n312 585
R1041 B.n311 B.n310 585
R1042 B.n309 B.n308 585
R1043 B.n307 B.n306 585
R1044 B.n305 B.n304 585
R1045 B.n303 B.n302 585
R1046 B.n301 B.n300 585
R1047 B.n299 B.n298 585
R1048 B.n297 B.n296 585
R1049 B.n295 B.n294 585
R1050 B.n293 B.n292 585
R1051 B.n291 B.n290 585
R1052 B.n288 B.n287 585
R1053 B.n286 B.n285 585
R1054 B.n284 B.n283 585
R1055 B.n282 B.n281 585
R1056 B.n280 B.n279 585
R1057 B.n278 B.n277 585
R1058 B.n276 B.n275 585
R1059 B.n274 B.n273 585
R1060 B.n272 B.n271 585
R1061 B.n270 B.n269 585
R1062 B.n268 B.n267 585
R1063 B.n266 B.n265 585
R1064 B.n264 B.n263 585
R1065 B.n262 B.n261 585
R1066 B.n260 B.n259 585
R1067 B.n258 B.n257 585
R1068 B.n256 B.n255 585
R1069 B.n254 B.n253 585
R1070 B.n252 B.n251 585
R1071 B.n250 B.n249 585
R1072 B.n248 B.n247 585
R1073 B.n246 B.n245 585
R1074 B.n244 B.n243 585
R1075 B.n242 B.n241 585
R1076 B.n240 B.n239 585
R1077 B.n238 B.n237 585
R1078 B.n236 B.n235 585
R1079 B.n234 B.n233 585
R1080 B.n232 B.n231 585
R1081 B.n230 B.n229 585
R1082 B.n228 B.n227 585
R1083 B.n226 B.n225 585
R1084 B.n224 B.n223 585
R1085 B.n222 B.n221 585
R1086 B.n220 B.n219 585
R1087 B.n218 B.n217 585
R1088 B.n216 B.n215 585
R1089 B.n214 B.n213 585
R1090 B.n212 B.n211 585
R1091 B.n210 B.n209 585
R1092 B.n208 B.n207 585
R1093 B.n206 B.n205 585
R1094 B.n204 B.n203 585
R1095 B.n202 B.n201 585
R1096 B.n200 B.n199 585
R1097 B.n198 B.n197 585
R1098 B.n196 B.n195 585
R1099 B.n194 B.n193 585
R1100 B.n192 B.n191 585
R1101 B.n190 B.n189 585
R1102 B.n188 B.n187 585
R1103 B.n186 B.n185 585
R1104 B.n184 B.n183 585
R1105 B.n182 B.n181 585
R1106 B.n180 B.n179 585
R1107 B.n178 B.n177 585
R1108 B.n176 B.n175 585
R1109 B.n174 B.n173 585
R1110 B.n172 B.n171 585
R1111 B.n170 B.n169 585
R1112 B.n168 B.n167 585
R1113 B.n102 B.n101 585
R1114 B.n1039 B.n1038 585
R1115 B.n1033 B.n161 585
R1116 B.n161 B.n99 585
R1117 B.n1032 B.n98 585
R1118 B.n1043 B.n98 585
R1119 B.n1031 B.n97 585
R1120 B.n1044 B.n97 585
R1121 B.n1030 B.n96 585
R1122 B.n1045 B.n96 585
R1123 B.n1029 B.n1028 585
R1124 B.n1028 B.n92 585
R1125 B.n1027 B.n91 585
R1126 B.n1051 B.n91 585
R1127 B.n1026 B.n90 585
R1128 B.n1052 B.n90 585
R1129 B.n1025 B.n89 585
R1130 B.t11 B.n89 585
R1131 B.n1024 B.n1023 585
R1132 B.n1023 B.n85 585
R1133 B.n1022 B.n84 585
R1134 B.n1058 B.n84 585
R1135 B.n1021 B.n83 585
R1136 B.n1059 B.n83 585
R1137 B.n1020 B.n82 585
R1138 B.n1060 B.n82 585
R1139 B.n1019 B.n1018 585
R1140 B.n1018 B.n78 585
R1141 B.n1017 B.n77 585
R1142 B.n1066 B.n77 585
R1143 B.n1016 B.n76 585
R1144 B.n1067 B.n76 585
R1145 B.n1015 B.n75 585
R1146 B.n1068 B.n75 585
R1147 B.n1014 B.n1013 585
R1148 B.n1013 B.n71 585
R1149 B.n1012 B.n70 585
R1150 B.n1074 B.n70 585
R1151 B.n1011 B.n69 585
R1152 B.n1075 B.n69 585
R1153 B.n1010 B.n68 585
R1154 B.n1076 B.n68 585
R1155 B.n1009 B.n1008 585
R1156 B.n1008 B.n64 585
R1157 B.n1007 B.n63 585
R1158 B.n1082 B.n63 585
R1159 B.n1006 B.n62 585
R1160 B.n1083 B.n62 585
R1161 B.n1005 B.n61 585
R1162 B.n1084 B.n61 585
R1163 B.n1004 B.n1003 585
R1164 B.n1003 B.n57 585
R1165 B.n1002 B.n56 585
R1166 B.n1090 B.n56 585
R1167 B.n1001 B.n55 585
R1168 B.n1091 B.n55 585
R1169 B.n1000 B.n54 585
R1170 B.n1092 B.n54 585
R1171 B.n999 B.n998 585
R1172 B.n998 B.n50 585
R1173 B.n997 B.n49 585
R1174 B.n1098 B.n49 585
R1175 B.n996 B.n48 585
R1176 B.n1099 B.n48 585
R1177 B.n995 B.n47 585
R1178 B.n1100 B.n47 585
R1179 B.n994 B.n993 585
R1180 B.n993 B.n43 585
R1181 B.n992 B.n42 585
R1182 B.n1106 B.n42 585
R1183 B.n991 B.n41 585
R1184 B.n1107 B.n41 585
R1185 B.n990 B.n40 585
R1186 B.n1108 B.n40 585
R1187 B.n989 B.n988 585
R1188 B.n988 B.n36 585
R1189 B.n987 B.n35 585
R1190 B.n1114 B.n35 585
R1191 B.n986 B.n34 585
R1192 B.n1115 B.n34 585
R1193 B.n985 B.n33 585
R1194 B.n1116 B.n33 585
R1195 B.n984 B.n983 585
R1196 B.n983 B.n29 585
R1197 B.n982 B.n28 585
R1198 B.n1122 B.n28 585
R1199 B.n981 B.n27 585
R1200 B.n1123 B.n27 585
R1201 B.n980 B.n26 585
R1202 B.n1124 B.n26 585
R1203 B.n979 B.n978 585
R1204 B.n978 B.n22 585
R1205 B.n977 B.n21 585
R1206 B.n1130 B.n21 585
R1207 B.n976 B.n20 585
R1208 B.n1131 B.n20 585
R1209 B.n975 B.n19 585
R1210 B.n1132 B.n19 585
R1211 B.n974 B.n973 585
R1212 B.n973 B.n15 585
R1213 B.n972 B.n14 585
R1214 B.n1138 B.n14 585
R1215 B.n971 B.n13 585
R1216 B.n1139 B.n13 585
R1217 B.n970 B.n12 585
R1218 B.n1140 B.n12 585
R1219 B.n969 B.n968 585
R1220 B.n968 B.n8 585
R1221 B.n967 B.n7 585
R1222 B.n1146 B.n7 585
R1223 B.n966 B.n6 585
R1224 B.n1147 B.n6 585
R1225 B.n965 B.n5 585
R1226 B.n1148 B.n5 585
R1227 B.n964 B.n963 585
R1228 B.n963 B.n4 585
R1229 B.n962 B.n395 585
R1230 B.n962 B.n961 585
R1231 B.n952 B.n396 585
R1232 B.n397 B.n396 585
R1233 B.n954 B.n953 585
R1234 B.n955 B.n954 585
R1235 B.n951 B.n402 585
R1236 B.n402 B.n401 585
R1237 B.n950 B.n949 585
R1238 B.n949 B.n948 585
R1239 B.n404 B.n403 585
R1240 B.n405 B.n404 585
R1241 B.n941 B.n940 585
R1242 B.n942 B.n941 585
R1243 B.n939 B.n410 585
R1244 B.n410 B.n409 585
R1245 B.n938 B.n937 585
R1246 B.n937 B.n936 585
R1247 B.n412 B.n411 585
R1248 B.n413 B.n412 585
R1249 B.n929 B.n928 585
R1250 B.n930 B.n929 585
R1251 B.n927 B.n418 585
R1252 B.n418 B.n417 585
R1253 B.n926 B.n925 585
R1254 B.n925 B.n924 585
R1255 B.n420 B.n419 585
R1256 B.n421 B.n420 585
R1257 B.n917 B.n916 585
R1258 B.n918 B.n917 585
R1259 B.n915 B.n426 585
R1260 B.n426 B.n425 585
R1261 B.n914 B.n913 585
R1262 B.n913 B.n912 585
R1263 B.n428 B.n427 585
R1264 B.n429 B.n428 585
R1265 B.n905 B.n904 585
R1266 B.n906 B.n905 585
R1267 B.n903 B.n434 585
R1268 B.n434 B.n433 585
R1269 B.n902 B.n901 585
R1270 B.n901 B.n900 585
R1271 B.n436 B.n435 585
R1272 B.n437 B.n436 585
R1273 B.n893 B.n892 585
R1274 B.n894 B.n893 585
R1275 B.n891 B.n442 585
R1276 B.n442 B.n441 585
R1277 B.n890 B.n889 585
R1278 B.n889 B.n888 585
R1279 B.n444 B.n443 585
R1280 B.n445 B.n444 585
R1281 B.n881 B.n880 585
R1282 B.n882 B.n881 585
R1283 B.n879 B.n450 585
R1284 B.n450 B.n449 585
R1285 B.n878 B.n877 585
R1286 B.n877 B.n876 585
R1287 B.n452 B.n451 585
R1288 B.n453 B.n452 585
R1289 B.n869 B.n868 585
R1290 B.n870 B.n869 585
R1291 B.n867 B.n458 585
R1292 B.n458 B.n457 585
R1293 B.n866 B.n865 585
R1294 B.n865 B.n864 585
R1295 B.n460 B.n459 585
R1296 B.n461 B.n460 585
R1297 B.n857 B.n856 585
R1298 B.n858 B.n857 585
R1299 B.n855 B.n465 585
R1300 B.n469 B.n465 585
R1301 B.n854 B.n853 585
R1302 B.n853 B.n852 585
R1303 B.n467 B.n466 585
R1304 B.n468 B.n467 585
R1305 B.n845 B.n844 585
R1306 B.n846 B.n845 585
R1307 B.n843 B.n474 585
R1308 B.n474 B.n473 585
R1309 B.n842 B.n841 585
R1310 B.n841 B.n840 585
R1311 B.n476 B.n475 585
R1312 B.n477 B.n476 585
R1313 B.n833 B.n832 585
R1314 B.n834 B.n833 585
R1315 B.n831 B.n482 585
R1316 B.n482 B.n481 585
R1317 B.n830 B.n829 585
R1318 B.n829 B.n828 585
R1319 B.n484 B.n483 585
R1320 B.n485 B.n484 585
R1321 B.n822 B.n821 585
R1322 B.t15 B.n822 585
R1323 B.n820 B.n490 585
R1324 B.n490 B.n489 585
R1325 B.n819 B.n818 585
R1326 B.n818 B.n817 585
R1327 B.n492 B.n491 585
R1328 B.n493 B.n492 585
R1329 B.n810 B.n809 585
R1330 B.n811 B.n810 585
R1331 B.n808 B.n498 585
R1332 B.n498 B.n497 585
R1333 B.n807 B.n806 585
R1334 B.n806 B.n805 585
R1335 B.n500 B.n499 585
R1336 B.n501 B.n500 585
R1337 B.n801 B.n800 585
R1338 B.n504 B.n503 585
R1339 B.n797 B.n796 585
R1340 B.n798 B.n797 585
R1341 B.n795 B.n562 585
R1342 B.n794 B.n793 585
R1343 B.n792 B.n791 585
R1344 B.n790 B.n789 585
R1345 B.n788 B.n787 585
R1346 B.n786 B.n785 585
R1347 B.n784 B.n783 585
R1348 B.n782 B.n781 585
R1349 B.n780 B.n779 585
R1350 B.n778 B.n777 585
R1351 B.n776 B.n775 585
R1352 B.n774 B.n773 585
R1353 B.n772 B.n771 585
R1354 B.n770 B.n769 585
R1355 B.n768 B.n767 585
R1356 B.n766 B.n765 585
R1357 B.n764 B.n763 585
R1358 B.n762 B.n761 585
R1359 B.n760 B.n759 585
R1360 B.n758 B.n757 585
R1361 B.n756 B.n755 585
R1362 B.n754 B.n753 585
R1363 B.n752 B.n751 585
R1364 B.n750 B.n749 585
R1365 B.n748 B.n747 585
R1366 B.n746 B.n745 585
R1367 B.n744 B.n743 585
R1368 B.n742 B.n741 585
R1369 B.n740 B.n739 585
R1370 B.n738 B.n737 585
R1371 B.n736 B.n735 585
R1372 B.n734 B.n733 585
R1373 B.n732 B.n731 585
R1374 B.n730 B.n729 585
R1375 B.n728 B.n727 585
R1376 B.n726 B.n725 585
R1377 B.n724 B.n723 585
R1378 B.n722 B.n721 585
R1379 B.n720 B.n719 585
R1380 B.n718 B.n717 585
R1381 B.n716 B.n715 585
R1382 B.n714 B.n713 585
R1383 B.n712 B.n711 585
R1384 B.n710 B.n709 585
R1385 B.n708 B.n707 585
R1386 B.n706 B.n705 585
R1387 B.n704 B.n703 585
R1388 B.n702 B.n701 585
R1389 B.n700 B.n699 585
R1390 B.n698 B.n697 585
R1391 B.n696 B.n695 585
R1392 B.n693 B.n692 585
R1393 B.n691 B.n690 585
R1394 B.n689 B.n688 585
R1395 B.n687 B.n686 585
R1396 B.n685 B.n684 585
R1397 B.n683 B.n682 585
R1398 B.n681 B.n680 585
R1399 B.n679 B.n678 585
R1400 B.n677 B.n676 585
R1401 B.n675 B.n674 585
R1402 B.n673 B.n672 585
R1403 B.n671 B.n670 585
R1404 B.n669 B.n668 585
R1405 B.n667 B.n666 585
R1406 B.n665 B.n664 585
R1407 B.n663 B.n662 585
R1408 B.n661 B.n660 585
R1409 B.n659 B.n658 585
R1410 B.n657 B.n656 585
R1411 B.n655 B.n654 585
R1412 B.n653 B.n652 585
R1413 B.n651 B.n650 585
R1414 B.n649 B.n648 585
R1415 B.n647 B.n646 585
R1416 B.n645 B.n644 585
R1417 B.n643 B.n642 585
R1418 B.n641 B.n640 585
R1419 B.n639 B.n638 585
R1420 B.n637 B.n636 585
R1421 B.n635 B.n634 585
R1422 B.n633 B.n632 585
R1423 B.n631 B.n630 585
R1424 B.n629 B.n628 585
R1425 B.n627 B.n626 585
R1426 B.n625 B.n624 585
R1427 B.n623 B.n622 585
R1428 B.n621 B.n620 585
R1429 B.n619 B.n618 585
R1430 B.n617 B.n616 585
R1431 B.n615 B.n614 585
R1432 B.n613 B.n612 585
R1433 B.n611 B.n610 585
R1434 B.n609 B.n608 585
R1435 B.n607 B.n606 585
R1436 B.n605 B.n604 585
R1437 B.n603 B.n602 585
R1438 B.n601 B.n600 585
R1439 B.n599 B.n598 585
R1440 B.n597 B.n596 585
R1441 B.n595 B.n594 585
R1442 B.n593 B.n592 585
R1443 B.n591 B.n590 585
R1444 B.n589 B.n588 585
R1445 B.n587 B.n586 585
R1446 B.n585 B.n584 585
R1447 B.n583 B.n582 585
R1448 B.n581 B.n580 585
R1449 B.n579 B.n578 585
R1450 B.n577 B.n576 585
R1451 B.n575 B.n574 585
R1452 B.n573 B.n572 585
R1453 B.n571 B.n570 585
R1454 B.n569 B.n568 585
R1455 B.n802 B.n502 585
R1456 B.n502 B.n501 585
R1457 B.n804 B.n803 585
R1458 B.n805 B.n804 585
R1459 B.n496 B.n495 585
R1460 B.n497 B.n496 585
R1461 B.n813 B.n812 585
R1462 B.n812 B.n811 585
R1463 B.n814 B.n494 585
R1464 B.n494 B.n493 585
R1465 B.n816 B.n815 585
R1466 B.n817 B.n816 585
R1467 B.n488 B.n487 585
R1468 B.n489 B.n488 585
R1469 B.n824 B.n823 585
R1470 B.n823 B.t15 585
R1471 B.n825 B.n486 585
R1472 B.n486 B.n485 585
R1473 B.n827 B.n826 585
R1474 B.n828 B.n827 585
R1475 B.n480 B.n479 585
R1476 B.n481 B.n480 585
R1477 B.n836 B.n835 585
R1478 B.n835 B.n834 585
R1479 B.n837 B.n478 585
R1480 B.n478 B.n477 585
R1481 B.n839 B.n838 585
R1482 B.n840 B.n839 585
R1483 B.n472 B.n471 585
R1484 B.n473 B.n472 585
R1485 B.n848 B.n847 585
R1486 B.n847 B.n846 585
R1487 B.n849 B.n470 585
R1488 B.n470 B.n468 585
R1489 B.n851 B.n850 585
R1490 B.n852 B.n851 585
R1491 B.n464 B.n463 585
R1492 B.n469 B.n464 585
R1493 B.n860 B.n859 585
R1494 B.n859 B.n858 585
R1495 B.n861 B.n462 585
R1496 B.n462 B.n461 585
R1497 B.n863 B.n862 585
R1498 B.n864 B.n863 585
R1499 B.n456 B.n455 585
R1500 B.n457 B.n456 585
R1501 B.n872 B.n871 585
R1502 B.n871 B.n870 585
R1503 B.n873 B.n454 585
R1504 B.n454 B.n453 585
R1505 B.n875 B.n874 585
R1506 B.n876 B.n875 585
R1507 B.n448 B.n447 585
R1508 B.n449 B.n448 585
R1509 B.n884 B.n883 585
R1510 B.n883 B.n882 585
R1511 B.n885 B.n446 585
R1512 B.n446 B.n445 585
R1513 B.n887 B.n886 585
R1514 B.n888 B.n887 585
R1515 B.n440 B.n439 585
R1516 B.n441 B.n440 585
R1517 B.n896 B.n895 585
R1518 B.n895 B.n894 585
R1519 B.n897 B.n438 585
R1520 B.n438 B.n437 585
R1521 B.n899 B.n898 585
R1522 B.n900 B.n899 585
R1523 B.n432 B.n431 585
R1524 B.n433 B.n432 585
R1525 B.n908 B.n907 585
R1526 B.n907 B.n906 585
R1527 B.n909 B.n430 585
R1528 B.n430 B.n429 585
R1529 B.n911 B.n910 585
R1530 B.n912 B.n911 585
R1531 B.n424 B.n423 585
R1532 B.n425 B.n424 585
R1533 B.n920 B.n919 585
R1534 B.n919 B.n918 585
R1535 B.n921 B.n422 585
R1536 B.n422 B.n421 585
R1537 B.n923 B.n922 585
R1538 B.n924 B.n923 585
R1539 B.n416 B.n415 585
R1540 B.n417 B.n416 585
R1541 B.n932 B.n931 585
R1542 B.n931 B.n930 585
R1543 B.n933 B.n414 585
R1544 B.n414 B.n413 585
R1545 B.n935 B.n934 585
R1546 B.n936 B.n935 585
R1547 B.n408 B.n407 585
R1548 B.n409 B.n408 585
R1549 B.n944 B.n943 585
R1550 B.n943 B.n942 585
R1551 B.n945 B.n406 585
R1552 B.n406 B.n405 585
R1553 B.n947 B.n946 585
R1554 B.n948 B.n947 585
R1555 B.n400 B.n399 585
R1556 B.n401 B.n400 585
R1557 B.n957 B.n956 585
R1558 B.n956 B.n955 585
R1559 B.n958 B.n398 585
R1560 B.n398 B.n397 585
R1561 B.n960 B.n959 585
R1562 B.n961 B.n960 585
R1563 B.n2 B.n0 585
R1564 B.n4 B.n2 585
R1565 B.n3 B.n1 585
R1566 B.n1147 B.n3 585
R1567 B.n1145 B.n1144 585
R1568 B.n1146 B.n1145 585
R1569 B.n1143 B.n9 585
R1570 B.n9 B.n8 585
R1571 B.n1142 B.n1141 585
R1572 B.n1141 B.n1140 585
R1573 B.n11 B.n10 585
R1574 B.n1139 B.n11 585
R1575 B.n1137 B.n1136 585
R1576 B.n1138 B.n1137 585
R1577 B.n1135 B.n16 585
R1578 B.n16 B.n15 585
R1579 B.n1134 B.n1133 585
R1580 B.n1133 B.n1132 585
R1581 B.n18 B.n17 585
R1582 B.n1131 B.n18 585
R1583 B.n1129 B.n1128 585
R1584 B.n1130 B.n1129 585
R1585 B.n1127 B.n23 585
R1586 B.n23 B.n22 585
R1587 B.n1126 B.n1125 585
R1588 B.n1125 B.n1124 585
R1589 B.n25 B.n24 585
R1590 B.n1123 B.n25 585
R1591 B.n1121 B.n1120 585
R1592 B.n1122 B.n1121 585
R1593 B.n1119 B.n30 585
R1594 B.n30 B.n29 585
R1595 B.n1118 B.n1117 585
R1596 B.n1117 B.n1116 585
R1597 B.n32 B.n31 585
R1598 B.n1115 B.n32 585
R1599 B.n1113 B.n1112 585
R1600 B.n1114 B.n1113 585
R1601 B.n1111 B.n37 585
R1602 B.n37 B.n36 585
R1603 B.n1110 B.n1109 585
R1604 B.n1109 B.n1108 585
R1605 B.n39 B.n38 585
R1606 B.n1107 B.n39 585
R1607 B.n1105 B.n1104 585
R1608 B.n1106 B.n1105 585
R1609 B.n1103 B.n44 585
R1610 B.n44 B.n43 585
R1611 B.n1102 B.n1101 585
R1612 B.n1101 B.n1100 585
R1613 B.n46 B.n45 585
R1614 B.n1099 B.n46 585
R1615 B.n1097 B.n1096 585
R1616 B.n1098 B.n1097 585
R1617 B.n1095 B.n51 585
R1618 B.n51 B.n50 585
R1619 B.n1094 B.n1093 585
R1620 B.n1093 B.n1092 585
R1621 B.n53 B.n52 585
R1622 B.n1091 B.n53 585
R1623 B.n1089 B.n1088 585
R1624 B.n1090 B.n1089 585
R1625 B.n1087 B.n58 585
R1626 B.n58 B.n57 585
R1627 B.n1086 B.n1085 585
R1628 B.n1085 B.n1084 585
R1629 B.n60 B.n59 585
R1630 B.n1083 B.n60 585
R1631 B.n1081 B.n1080 585
R1632 B.n1082 B.n1081 585
R1633 B.n1079 B.n65 585
R1634 B.n65 B.n64 585
R1635 B.n1078 B.n1077 585
R1636 B.n1077 B.n1076 585
R1637 B.n67 B.n66 585
R1638 B.n1075 B.n67 585
R1639 B.n1073 B.n1072 585
R1640 B.n1074 B.n1073 585
R1641 B.n1071 B.n72 585
R1642 B.n72 B.n71 585
R1643 B.n1070 B.n1069 585
R1644 B.n1069 B.n1068 585
R1645 B.n74 B.n73 585
R1646 B.n1067 B.n74 585
R1647 B.n1065 B.n1064 585
R1648 B.n1066 B.n1065 585
R1649 B.n1063 B.n79 585
R1650 B.n79 B.n78 585
R1651 B.n1062 B.n1061 585
R1652 B.n1061 B.n1060 585
R1653 B.n81 B.n80 585
R1654 B.n1059 B.n81 585
R1655 B.n1057 B.n1056 585
R1656 B.n1058 B.n1057 585
R1657 B.n1055 B.n86 585
R1658 B.n86 B.n85 585
R1659 B.n1054 B.n1053 585
R1660 B.n1053 B.t11 585
R1661 B.n88 B.n87 585
R1662 B.n1052 B.n88 585
R1663 B.n1050 B.n1049 585
R1664 B.n1051 B.n1050 585
R1665 B.n1048 B.n93 585
R1666 B.n93 B.n92 585
R1667 B.n1047 B.n1046 585
R1668 B.n1046 B.n1045 585
R1669 B.n95 B.n94 585
R1670 B.n1044 B.n95 585
R1671 B.n1042 B.n1041 585
R1672 B.n1043 B.n1042 585
R1673 B.n1040 B.n100 585
R1674 B.n100 B.n99 585
R1675 B.n1150 B.n1149 585
R1676 B.n1149 B.n1148 585
R1677 B.n800 B.n502 535.745
R1678 B.n1038 B.n100 535.745
R1679 B.n568 B.n500 535.745
R1680 B.n1035 B.n161 535.745
R1681 B.n565 B.t23 404.647
R1682 B.n162 B.t19 404.647
R1683 B.n563 B.t17 404.647
R1684 B.n164 B.t12 404.647
R1685 B.n565 B.t21 373.538
R1686 B.n563 B.t14 373.538
R1687 B.n164 B.t10 373.538
R1688 B.n162 B.t18 373.538
R1689 B.n566 B.t22 352.865
R1690 B.n163 B.t20 352.865
R1691 B.n564 B.t16 352.865
R1692 B.n165 B.t13 352.865
R1693 B.n1036 B.n159 256.663
R1694 B.n1036 B.n158 256.663
R1695 B.n1036 B.n157 256.663
R1696 B.n1036 B.n156 256.663
R1697 B.n1036 B.n155 256.663
R1698 B.n1036 B.n154 256.663
R1699 B.n1036 B.n153 256.663
R1700 B.n1036 B.n152 256.663
R1701 B.n1036 B.n151 256.663
R1702 B.n1036 B.n150 256.663
R1703 B.n1036 B.n149 256.663
R1704 B.n1036 B.n148 256.663
R1705 B.n1036 B.n147 256.663
R1706 B.n1036 B.n146 256.663
R1707 B.n1036 B.n145 256.663
R1708 B.n1036 B.n144 256.663
R1709 B.n1036 B.n143 256.663
R1710 B.n1036 B.n142 256.663
R1711 B.n1036 B.n141 256.663
R1712 B.n1036 B.n140 256.663
R1713 B.n1036 B.n139 256.663
R1714 B.n1036 B.n138 256.663
R1715 B.n1036 B.n137 256.663
R1716 B.n1036 B.n136 256.663
R1717 B.n1036 B.n135 256.663
R1718 B.n1036 B.n134 256.663
R1719 B.n1036 B.n133 256.663
R1720 B.n1036 B.n132 256.663
R1721 B.n1036 B.n131 256.663
R1722 B.n1036 B.n130 256.663
R1723 B.n1036 B.n129 256.663
R1724 B.n1036 B.n128 256.663
R1725 B.n1036 B.n127 256.663
R1726 B.n1036 B.n126 256.663
R1727 B.n1036 B.n125 256.663
R1728 B.n1036 B.n124 256.663
R1729 B.n1036 B.n123 256.663
R1730 B.n1036 B.n122 256.663
R1731 B.n1036 B.n121 256.663
R1732 B.n1036 B.n120 256.663
R1733 B.n1036 B.n119 256.663
R1734 B.n1036 B.n118 256.663
R1735 B.n1036 B.n117 256.663
R1736 B.n1036 B.n116 256.663
R1737 B.n1036 B.n115 256.663
R1738 B.n1036 B.n114 256.663
R1739 B.n1036 B.n113 256.663
R1740 B.n1036 B.n112 256.663
R1741 B.n1036 B.n111 256.663
R1742 B.n1036 B.n110 256.663
R1743 B.n1036 B.n109 256.663
R1744 B.n1036 B.n108 256.663
R1745 B.n1036 B.n107 256.663
R1746 B.n1036 B.n106 256.663
R1747 B.n1036 B.n105 256.663
R1748 B.n1036 B.n104 256.663
R1749 B.n1036 B.n103 256.663
R1750 B.n1037 B.n1036 256.663
R1751 B.n799 B.n798 256.663
R1752 B.n798 B.n505 256.663
R1753 B.n798 B.n506 256.663
R1754 B.n798 B.n507 256.663
R1755 B.n798 B.n508 256.663
R1756 B.n798 B.n509 256.663
R1757 B.n798 B.n510 256.663
R1758 B.n798 B.n511 256.663
R1759 B.n798 B.n512 256.663
R1760 B.n798 B.n513 256.663
R1761 B.n798 B.n514 256.663
R1762 B.n798 B.n515 256.663
R1763 B.n798 B.n516 256.663
R1764 B.n798 B.n517 256.663
R1765 B.n798 B.n518 256.663
R1766 B.n798 B.n519 256.663
R1767 B.n798 B.n520 256.663
R1768 B.n798 B.n521 256.663
R1769 B.n798 B.n522 256.663
R1770 B.n798 B.n523 256.663
R1771 B.n798 B.n524 256.663
R1772 B.n798 B.n525 256.663
R1773 B.n798 B.n526 256.663
R1774 B.n798 B.n527 256.663
R1775 B.n798 B.n528 256.663
R1776 B.n798 B.n529 256.663
R1777 B.n798 B.n530 256.663
R1778 B.n798 B.n531 256.663
R1779 B.n798 B.n532 256.663
R1780 B.n798 B.n533 256.663
R1781 B.n798 B.n534 256.663
R1782 B.n798 B.n535 256.663
R1783 B.n798 B.n536 256.663
R1784 B.n798 B.n537 256.663
R1785 B.n798 B.n538 256.663
R1786 B.n798 B.n539 256.663
R1787 B.n798 B.n540 256.663
R1788 B.n798 B.n541 256.663
R1789 B.n798 B.n542 256.663
R1790 B.n798 B.n543 256.663
R1791 B.n798 B.n544 256.663
R1792 B.n798 B.n545 256.663
R1793 B.n798 B.n546 256.663
R1794 B.n798 B.n547 256.663
R1795 B.n798 B.n548 256.663
R1796 B.n798 B.n549 256.663
R1797 B.n798 B.n550 256.663
R1798 B.n798 B.n551 256.663
R1799 B.n798 B.n552 256.663
R1800 B.n798 B.n553 256.663
R1801 B.n798 B.n554 256.663
R1802 B.n798 B.n555 256.663
R1803 B.n798 B.n556 256.663
R1804 B.n798 B.n557 256.663
R1805 B.n798 B.n558 256.663
R1806 B.n798 B.n559 256.663
R1807 B.n798 B.n560 256.663
R1808 B.n798 B.n561 256.663
R1809 B.n804 B.n502 163.367
R1810 B.n804 B.n496 163.367
R1811 B.n812 B.n496 163.367
R1812 B.n812 B.n494 163.367
R1813 B.n816 B.n494 163.367
R1814 B.n816 B.n488 163.367
R1815 B.n823 B.n488 163.367
R1816 B.n823 B.n486 163.367
R1817 B.n827 B.n486 163.367
R1818 B.n827 B.n480 163.367
R1819 B.n835 B.n480 163.367
R1820 B.n835 B.n478 163.367
R1821 B.n839 B.n478 163.367
R1822 B.n839 B.n472 163.367
R1823 B.n847 B.n472 163.367
R1824 B.n847 B.n470 163.367
R1825 B.n851 B.n470 163.367
R1826 B.n851 B.n464 163.367
R1827 B.n859 B.n464 163.367
R1828 B.n859 B.n462 163.367
R1829 B.n863 B.n462 163.367
R1830 B.n863 B.n456 163.367
R1831 B.n871 B.n456 163.367
R1832 B.n871 B.n454 163.367
R1833 B.n875 B.n454 163.367
R1834 B.n875 B.n448 163.367
R1835 B.n883 B.n448 163.367
R1836 B.n883 B.n446 163.367
R1837 B.n887 B.n446 163.367
R1838 B.n887 B.n440 163.367
R1839 B.n895 B.n440 163.367
R1840 B.n895 B.n438 163.367
R1841 B.n899 B.n438 163.367
R1842 B.n899 B.n432 163.367
R1843 B.n907 B.n432 163.367
R1844 B.n907 B.n430 163.367
R1845 B.n911 B.n430 163.367
R1846 B.n911 B.n424 163.367
R1847 B.n919 B.n424 163.367
R1848 B.n919 B.n422 163.367
R1849 B.n923 B.n422 163.367
R1850 B.n923 B.n416 163.367
R1851 B.n931 B.n416 163.367
R1852 B.n931 B.n414 163.367
R1853 B.n935 B.n414 163.367
R1854 B.n935 B.n408 163.367
R1855 B.n943 B.n408 163.367
R1856 B.n943 B.n406 163.367
R1857 B.n947 B.n406 163.367
R1858 B.n947 B.n400 163.367
R1859 B.n956 B.n400 163.367
R1860 B.n956 B.n398 163.367
R1861 B.n960 B.n398 163.367
R1862 B.n960 B.n2 163.367
R1863 B.n1149 B.n2 163.367
R1864 B.n1149 B.n3 163.367
R1865 B.n1145 B.n3 163.367
R1866 B.n1145 B.n9 163.367
R1867 B.n1141 B.n9 163.367
R1868 B.n1141 B.n11 163.367
R1869 B.n1137 B.n11 163.367
R1870 B.n1137 B.n16 163.367
R1871 B.n1133 B.n16 163.367
R1872 B.n1133 B.n18 163.367
R1873 B.n1129 B.n18 163.367
R1874 B.n1129 B.n23 163.367
R1875 B.n1125 B.n23 163.367
R1876 B.n1125 B.n25 163.367
R1877 B.n1121 B.n25 163.367
R1878 B.n1121 B.n30 163.367
R1879 B.n1117 B.n30 163.367
R1880 B.n1117 B.n32 163.367
R1881 B.n1113 B.n32 163.367
R1882 B.n1113 B.n37 163.367
R1883 B.n1109 B.n37 163.367
R1884 B.n1109 B.n39 163.367
R1885 B.n1105 B.n39 163.367
R1886 B.n1105 B.n44 163.367
R1887 B.n1101 B.n44 163.367
R1888 B.n1101 B.n46 163.367
R1889 B.n1097 B.n46 163.367
R1890 B.n1097 B.n51 163.367
R1891 B.n1093 B.n51 163.367
R1892 B.n1093 B.n53 163.367
R1893 B.n1089 B.n53 163.367
R1894 B.n1089 B.n58 163.367
R1895 B.n1085 B.n58 163.367
R1896 B.n1085 B.n60 163.367
R1897 B.n1081 B.n60 163.367
R1898 B.n1081 B.n65 163.367
R1899 B.n1077 B.n65 163.367
R1900 B.n1077 B.n67 163.367
R1901 B.n1073 B.n67 163.367
R1902 B.n1073 B.n72 163.367
R1903 B.n1069 B.n72 163.367
R1904 B.n1069 B.n74 163.367
R1905 B.n1065 B.n74 163.367
R1906 B.n1065 B.n79 163.367
R1907 B.n1061 B.n79 163.367
R1908 B.n1061 B.n81 163.367
R1909 B.n1057 B.n81 163.367
R1910 B.n1057 B.n86 163.367
R1911 B.n1053 B.n86 163.367
R1912 B.n1053 B.n88 163.367
R1913 B.n1050 B.n88 163.367
R1914 B.n1050 B.n93 163.367
R1915 B.n1046 B.n93 163.367
R1916 B.n1046 B.n95 163.367
R1917 B.n1042 B.n95 163.367
R1918 B.n1042 B.n100 163.367
R1919 B.n797 B.n504 163.367
R1920 B.n797 B.n562 163.367
R1921 B.n793 B.n792 163.367
R1922 B.n789 B.n788 163.367
R1923 B.n785 B.n784 163.367
R1924 B.n781 B.n780 163.367
R1925 B.n777 B.n776 163.367
R1926 B.n773 B.n772 163.367
R1927 B.n769 B.n768 163.367
R1928 B.n765 B.n764 163.367
R1929 B.n761 B.n760 163.367
R1930 B.n757 B.n756 163.367
R1931 B.n753 B.n752 163.367
R1932 B.n749 B.n748 163.367
R1933 B.n745 B.n744 163.367
R1934 B.n741 B.n740 163.367
R1935 B.n737 B.n736 163.367
R1936 B.n733 B.n732 163.367
R1937 B.n729 B.n728 163.367
R1938 B.n725 B.n724 163.367
R1939 B.n721 B.n720 163.367
R1940 B.n717 B.n716 163.367
R1941 B.n713 B.n712 163.367
R1942 B.n709 B.n708 163.367
R1943 B.n705 B.n704 163.367
R1944 B.n701 B.n700 163.367
R1945 B.n697 B.n696 163.367
R1946 B.n692 B.n691 163.367
R1947 B.n688 B.n687 163.367
R1948 B.n684 B.n683 163.367
R1949 B.n680 B.n679 163.367
R1950 B.n676 B.n675 163.367
R1951 B.n672 B.n671 163.367
R1952 B.n668 B.n667 163.367
R1953 B.n664 B.n663 163.367
R1954 B.n660 B.n659 163.367
R1955 B.n656 B.n655 163.367
R1956 B.n652 B.n651 163.367
R1957 B.n648 B.n647 163.367
R1958 B.n644 B.n643 163.367
R1959 B.n640 B.n639 163.367
R1960 B.n636 B.n635 163.367
R1961 B.n632 B.n631 163.367
R1962 B.n628 B.n627 163.367
R1963 B.n624 B.n623 163.367
R1964 B.n620 B.n619 163.367
R1965 B.n616 B.n615 163.367
R1966 B.n612 B.n611 163.367
R1967 B.n608 B.n607 163.367
R1968 B.n604 B.n603 163.367
R1969 B.n600 B.n599 163.367
R1970 B.n596 B.n595 163.367
R1971 B.n592 B.n591 163.367
R1972 B.n588 B.n587 163.367
R1973 B.n584 B.n583 163.367
R1974 B.n580 B.n579 163.367
R1975 B.n576 B.n575 163.367
R1976 B.n572 B.n571 163.367
R1977 B.n806 B.n500 163.367
R1978 B.n806 B.n498 163.367
R1979 B.n810 B.n498 163.367
R1980 B.n810 B.n492 163.367
R1981 B.n818 B.n492 163.367
R1982 B.n818 B.n490 163.367
R1983 B.n822 B.n490 163.367
R1984 B.n822 B.n484 163.367
R1985 B.n829 B.n484 163.367
R1986 B.n829 B.n482 163.367
R1987 B.n833 B.n482 163.367
R1988 B.n833 B.n476 163.367
R1989 B.n841 B.n476 163.367
R1990 B.n841 B.n474 163.367
R1991 B.n845 B.n474 163.367
R1992 B.n845 B.n467 163.367
R1993 B.n853 B.n467 163.367
R1994 B.n853 B.n465 163.367
R1995 B.n857 B.n465 163.367
R1996 B.n857 B.n460 163.367
R1997 B.n865 B.n460 163.367
R1998 B.n865 B.n458 163.367
R1999 B.n869 B.n458 163.367
R2000 B.n869 B.n452 163.367
R2001 B.n877 B.n452 163.367
R2002 B.n877 B.n450 163.367
R2003 B.n881 B.n450 163.367
R2004 B.n881 B.n444 163.367
R2005 B.n889 B.n444 163.367
R2006 B.n889 B.n442 163.367
R2007 B.n893 B.n442 163.367
R2008 B.n893 B.n436 163.367
R2009 B.n901 B.n436 163.367
R2010 B.n901 B.n434 163.367
R2011 B.n905 B.n434 163.367
R2012 B.n905 B.n428 163.367
R2013 B.n913 B.n428 163.367
R2014 B.n913 B.n426 163.367
R2015 B.n917 B.n426 163.367
R2016 B.n917 B.n420 163.367
R2017 B.n925 B.n420 163.367
R2018 B.n925 B.n418 163.367
R2019 B.n929 B.n418 163.367
R2020 B.n929 B.n412 163.367
R2021 B.n937 B.n412 163.367
R2022 B.n937 B.n410 163.367
R2023 B.n941 B.n410 163.367
R2024 B.n941 B.n404 163.367
R2025 B.n949 B.n404 163.367
R2026 B.n949 B.n402 163.367
R2027 B.n954 B.n402 163.367
R2028 B.n954 B.n396 163.367
R2029 B.n962 B.n396 163.367
R2030 B.n963 B.n962 163.367
R2031 B.n963 B.n5 163.367
R2032 B.n6 B.n5 163.367
R2033 B.n7 B.n6 163.367
R2034 B.n968 B.n7 163.367
R2035 B.n968 B.n12 163.367
R2036 B.n13 B.n12 163.367
R2037 B.n14 B.n13 163.367
R2038 B.n973 B.n14 163.367
R2039 B.n973 B.n19 163.367
R2040 B.n20 B.n19 163.367
R2041 B.n21 B.n20 163.367
R2042 B.n978 B.n21 163.367
R2043 B.n978 B.n26 163.367
R2044 B.n27 B.n26 163.367
R2045 B.n28 B.n27 163.367
R2046 B.n983 B.n28 163.367
R2047 B.n983 B.n33 163.367
R2048 B.n34 B.n33 163.367
R2049 B.n35 B.n34 163.367
R2050 B.n988 B.n35 163.367
R2051 B.n988 B.n40 163.367
R2052 B.n41 B.n40 163.367
R2053 B.n42 B.n41 163.367
R2054 B.n993 B.n42 163.367
R2055 B.n993 B.n47 163.367
R2056 B.n48 B.n47 163.367
R2057 B.n49 B.n48 163.367
R2058 B.n998 B.n49 163.367
R2059 B.n998 B.n54 163.367
R2060 B.n55 B.n54 163.367
R2061 B.n56 B.n55 163.367
R2062 B.n1003 B.n56 163.367
R2063 B.n1003 B.n61 163.367
R2064 B.n62 B.n61 163.367
R2065 B.n63 B.n62 163.367
R2066 B.n1008 B.n63 163.367
R2067 B.n1008 B.n68 163.367
R2068 B.n69 B.n68 163.367
R2069 B.n70 B.n69 163.367
R2070 B.n1013 B.n70 163.367
R2071 B.n1013 B.n75 163.367
R2072 B.n76 B.n75 163.367
R2073 B.n77 B.n76 163.367
R2074 B.n1018 B.n77 163.367
R2075 B.n1018 B.n82 163.367
R2076 B.n83 B.n82 163.367
R2077 B.n84 B.n83 163.367
R2078 B.n1023 B.n84 163.367
R2079 B.n1023 B.n89 163.367
R2080 B.n90 B.n89 163.367
R2081 B.n91 B.n90 163.367
R2082 B.n1028 B.n91 163.367
R2083 B.n1028 B.n96 163.367
R2084 B.n97 B.n96 163.367
R2085 B.n98 B.n97 163.367
R2086 B.n161 B.n98 163.367
R2087 B.n167 B.n102 163.367
R2088 B.n171 B.n170 163.367
R2089 B.n175 B.n174 163.367
R2090 B.n179 B.n178 163.367
R2091 B.n183 B.n182 163.367
R2092 B.n187 B.n186 163.367
R2093 B.n191 B.n190 163.367
R2094 B.n195 B.n194 163.367
R2095 B.n199 B.n198 163.367
R2096 B.n203 B.n202 163.367
R2097 B.n207 B.n206 163.367
R2098 B.n211 B.n210 163.367
R2099 B.n215 B.n214 163.367
R2100 B.n219 B.n218 163.367
R2101 B.n223 B.n222 163.367
R2102 B.n227 B.n226 163.367
R2103 B.n231 B.n230 163.367
R2104 B.n235 B.n234 163.367
R2105 B.n239 B.n238 163.367
R2106 B.n243 B.n242 163.367
R2107 B.n247 B.n246 163.367
R2108 B.n251 B.n250 163.367
R2109 B.n255 B.n254 163.367
R2110 B.n259 B.n258 163.367
R2111 B.n263 B.n262 163.367
R2112 B.n267 B.n266 163.367
R2113 B.n271 B.n270 163.367
R2114 B.n275 B.n274 163.367
R2115 B.n279 B.n278 163.367
R2116 B.n283 B.n282 163.367
R2117 B.n287 B.n286 163.367
R2118 B.n292 B.n291 163.367
R2119 B.n296 B.n295 163.367
R2120 B.n300 B.n299 163.367
R2121 B.n304 B.n303 163.367
R2122 B.n308 B.n307 163.367
R2123 B.n312 B.n311 163.367
R2124 B.n316 B.n315 163.367
R2125 B.n320 B.n319 163.367
R2126 B.n324 B.n323 163.367
R2127 B.n328 B.n327 163.367
R2128 B.n332 B.n331 163.367
R2129 B.n336 B.n335 163.367
R2130 B.n340 B.n339 163.367
R2131 B.n344 B.n343 163.367
R2132 B.n348 B.n347 163.367
R2133 B.n352 B.n351 163.367
R2134 B.n356 B.n355 163.367
R2135 B.n360 B.n359 163.367
R2136 B.n364 B.n363 163.367
R2137 B.n368 B.n367 163.367
R2138 B.n372 B.n371 163.367
R2139 B.n376 B.n375 163.367
R2140 B.n380 B.n379 163.367
R2141 B.n384 B.n383 163.367
R2142 B.n388 B.n387 163.367
R2143 B.n392 B.n391 163.367
R2144 B.n1035 B.n160 163.367
R2145 B.n800 B.n799 71.676
R2146 B.n562 B.n505 71.676
R2147 B.n792 B.n506 71.676
R2148 B.n788 B.n507 71.676
R2149 B.n784 B.n508 71.676
R2150 B.n780 B.n509 71.676
R2151 B.n776 B.n510 71.676
R2152 B.n772 B.n511 71.676
R2153 B.n768 B.n512 71.676
R2154 B.n764 B.n513 71.676
R2155 B.n760 B.n514 71.676
R2156 B.n756 B.n515 71.676
R2157 B.n752 B.n516 71.676
R2158 B.n748 B.n517 71.676
R2159 B.n744 B.n518 71.676
R2160 B.n740 B.n519 71.676
R2161 B.n736 B.n520 71.676
R2162 B.n732 B.n521 71.676
R2163 B.n728 B.n522 71.676
R2164 B.n724 B.n523 71.676
R2165 B.n720 B.n524 71.676
R2166 B.n716 B.n525 71.676
R2167 B.n712 B.n526 71.676
R2168 B.n708 B.n527 71.676
R2169 B.n704 B.n528 71.676
R2170 B.n700 B.n529 71.676
R2171 B.n696 B.n530 71.676
R2172 B.n691 B.n531 71.676
R2173 B.n687 B.n532 71.676
R2174 B.n683 B.n533 71.676
R2175 B.n679 B.n534 71.676
R2176 B.n675 B.n535 71.676
R2177 B.n671 B.n536 71.676
R2178 B.n667 B.n537 71.676
R2179 B.n663 B.n538 71.676
R2180 B.n659 B.n539 71.676
R2181 B.n655 B.n540 71.676
R2182 B.n651 B.n541 71.676
R2183 B.n647 B.n542 71.676
R2184 B.n643 B.n543 71.676
R2185 B.n639 B.n544 71.676
R2186 B.n635 B.n545 71.676
R2187 B.n631 B.n546 71.676
R2188 B.n627 B.n547 71.676
R2189 B.n623 B.n548 71.676
R2190 B.n619 B.n549 71.676
R2191 B.n615 B.n550 71.676
R2192 B.n611 B.n551 71.676
R2193 B.n607 B.n552 71.676
R2194 B.n603 B.n553 71.676
R2195 B.n599 B.n554 71.676
R2196 B.n595 B.n555 71.676
R2197 B.n591 B.n556 71.676
R2198 B.n587 B.n557 71.676
R2199 B.n583 B.n558 71.676
R2200 B.n579 B.n559 71.676
R2201 B.n575 B.n560 71.676
R2202 B.n571 B.n561 71.676
R2203 B.n1038 B.n1037 71.676
R2204 B.n167 B.n103 71.676
R2205 B.n171 B.n104 71.676
R2206 B.n175 B.n105 71.676
R2207 B.n179 B.n106 71.676
R2208 B.n183 B.n107 71.676
R2209 B.n187 B.n108 71.676
R2210 B.n191 B.n109 71.676
R2211 B.n195 B.n110 71.676
R2212 B.n199 B.n111 71.676
R2213 B.n203 B.n112 71.676
R2214 B.n207 B.n113 71.676
R2215 B.n211 B.n114 71.676
R2216 B.n215 B.n115 71.676
R2217 B.n219 B.n116 71.676
R2218 B.n223 B.n117 71.676
R2219 B.n227 B.n118 71.676
R2220 B.n231 B.n119 71.676
R2221 B.n235 B.n120 71.676
R2222 B.n239 B.n121 71.676
R2223 B.n243 B.n122 71.676
R2224 B.n247 B.n123 71.676
R2225 B.n251 B.n124 71.676
R2226 B.n255 B.n125 71.676
R2227 B.n259 B.n126 71.676
R2228 B.n263 B.n127 71.676
R2229 B.n267 B.n128 71.676
R2230 B.n271 B.n129 71.676
R2231 B.n275 B.n130 71.676
R2232 B.n279 B.n131 71.676
R2233 B.n283 B.n132 71.676
R2234 B.n287 B.n133 71.676
R2235 B.n292 B.n134 71.676
R2236 B.n296 B.n135 71.676
R2237 B.n300 B.n136 71.676
R2238 B.n304 B.n137 71.676
R2239 B.n308 B.n138 71.676
R2240 B.n312 B.n139 71.676
R2241 B.n316 B.n140 71.676
R2242 B.n320 B.n141 71.676
R2243 B.n324 B.n142 71.676
R2244 B.n328 B.n143 71.676
R2245 B.n332 B.n144 71.676
R2246 B.n336 B.n145 71.676
R2247 B.n340 B.n146 71.676
R2248 B.n344 B.n147 71.676
R2249 B.n348 B.n148 71.676
R2250 B.n352 B.n149 71.676
R2251 B.n356 B.n150 71.676
R2252 B.n360 B.n151 71.676
R2253 B.n364 B.n152 71.676
R2254 B.n368 B.n153 71.676
R2255 B.n372 B.n154 71.676
R2256 B.n376 B.n155 71.676
R2257 B.n380 B.n156 71.676
R2258 B.n384 B.n157 71.676
R2259 B.n388 B.n158 71.676
R2260 B.n392 B.n159 71.676
R2261 B.n160 B.n159 71.676
R2262 B.n391 B.n158 71.676
R2263 B.n387 B.n157 71.676
R2264 B.n383 B.n156 71.676
R2265 B.n379 B.n155 71.676
R2266 B.n375 B.n154 71.676
R2267 B.n371 B.n153 71.676
R2268 B.n367 B.n152 71.676
R2269 B.n363 B.n151 71.676
R2270 B.n359 B.n150 71.676
R2271 B.n355 B.n149 71.676
R2272 B.n351 B.n148 71.676
R2273 B.n347 B.n147 71.676
R2274 B.n343 B.n146 71.676
R2275 B.n339 B.n145 71.676
R2276 B.n335 B.n144 71.676
R2277 B.n331 B.n143 71.676
R2278 B.n327 B.n142 71.676
R2279 B.n323 B.n141 71.676
R2280 B.n319 B.n140 71.676
R2281 B.n315 B.n139 71.676
R2282 B.n311 B.n138 71.676
R2283 B.n307 B.n137 71.676
R2284 B.n303 B.n136 71.676
R2285 B.n299 B.n135 71.676
R2286 B.n295 B.n134 71.676
R2287 B.n291 B.n133 71.676
R2288 B.n286 B.n132 71.676
R2289 B.n282 B.n131 71.676
R2290 B.n278 B.n130 71.676
R2291 B.n274 B.n129 71.676
R2292 B.n270 B.n128 71.676
R2293 B.n266 B.n127 71.676
R2294 B.n262 B.n126 71.676
R2295 B.n258 B.n125 71.676
R2296 B.n254 B.n124 71.676
R2297 B.n250 B.n123 71.676
R2298 B.n246 B.n122 71.676
R2299 B.n242 B.n121 71.676
R2300 B.n238 B.n120 71.676
R2301 B.n234 B.n119 71.676
R2302 B.n230 B.n118 71.676
R2303 B.n226 B.n117 71.676
R2304 B.n222 B.n116 71.676
R2305 B.n218 B.n115 71.676
R2306 B.n214 B.n114 71.676
R2307 B.n210 B.n113 71.676
R2308 B.n206 B.n112 71.676
R2309 B.n202 B.n111 71.676
R2310 B.n198 B.n110 71.676
R2311 B.n194 B.n109 71.676
R2312 B.n190 B.n108 71.676
R2313 B.n186 B.n107 71.676
R2314 B.n182 B.n106 71.676
R2315 B.n178 B.n105 71.676
R2316 B.n174 B.n104 71.676
R2317 B.n170 B.n103 71.676
R2318 B.n1037 B.n102 71.676
R2319 B.n799 B.n504 71.676
R2320 B.n793 B.n505 71.676
R2321 B.n789 B.n506 71.676
R2322 B.n785 B.n507 71.676
R2323 B.n781 B.n508 71.676
R2324 B.n777 B.n509 71.676
R2325 B.n773 B.n510 71.676
R2326 B.n769 B.n511 71.676
R2327 B.n765 B.n512 71.676
R2328 B.n761 B.n513 71.676
R2329 B.n757 B.n514 71.676
R2330 B.n753 B.n515 71.676
R2331 B.n749 B.n516 71.676
R2332 B.n745 B.n517 71.676
R2333 B.n741 B.n518 71.676
R2334 B.n737 B.n519 71.676
R2335 B.n733 B.n520 71.676
R2336 B.n729 B.n521 71.676
R2337 B.n725 B.n522 71.676
R2338 B.n721 B.n523 71.676
R2339 B.n717 B.n524 71.676
R2340 B.n713 B.n525 71.676
R2341 B.n709 B.n526 71.676
R2342 B.n705 B.n527 71.676
R2343 B.n701 B.n528 71.676
R2344 B.n697 B.n529 71.676
R2345 B.n692 B.n530 71.676
R2346 B.n688 B.n531 71.676
R2347 B.n684 B.n532 71.676
R2348 B.n680 B.n533 71.676
R2349 B.n676 B.n534 71.676
R2350 B.n672 B.n535 71.676
R2351 B.n668 B.n536 71.676
R2352 B.n664 B.n537 71.676
R2353 B.n660 B.n538 71.676
R2354 B.n656 B.n539 71.676
R2355 B.n652 B.n540 71.676
R2356 B.n648 B.n541 71.676
R2357 B.n644 B.n542 71.676
R2358 B.n640 B.n543 71.676
R2359 B.n636 B.n544 71.676
R2360 B.n632 B.n545 71.676
R2361 B.n628 B.n546 71.676
R2362 B.n624 B.n547 71.676
R2363 B.n620 B.n548 71.676
R2364 B.n616 B.n549 71.676
R2365 B.n612 B.n550 71.676
R2366 B.n608 B.n551 71.676
R2367 B.n604 B.n552 71.676
R2368 B.n600 B.n553 71.676
R2369 B.n596 B.n554 71.676
R2370 B.n592 B.n555 71.676
R2371 B.n588 B.n556 71.676
R2372 B.n584 B.n557 71.676
R2373 B.n580 B.n558 71.676
R2374 B.n576 B.n559 71.676
R2375 B.n572 B.n560 71.676
R2376 B.n568 B.n561 71.676
R2377 B.n798 B.n501 71.4992
R2378 B.n1036 B.n99 71.4992
R2379 B.n567 B.n566 59.5399
R2380 B.n694 B.n564 59.5399
R2381 B.n166 B.n165 59.5399
R2382 B.n289 B.n163 59.5399
R2383 B.n566 B.n565 51.7823
R2384 B.n564 B.n563 51.7823
R2385 B.n165 B.n164 51.7823
R2386 B.n163 B.n162 51.7823
R2387 B.n805 B.n501 34.9783
R2388 B.n805 B.n497 34.9783
R2389 B.n811 B.n497 34.9783
R2390 B.n811 B.n493 34.9783
R2391 B.n817 B.n493 34.9783
R2392 B.n817 B.n489 34.9783
R2393 B.t15 B.n489 34.9783
R2394 B.t15 B.n485 34.9783
R2395 B.n828 B.n485 34.9783
R2396 B.n828 B.n481 34.9783
R2397 B.n834 B.n481 34.9783
R2398 B.n834 B.n477 34.9783
R2399 B.n840 B.n477 34.9783
R2400 B.n840 B.n473 34.9783
R2401 B.n846 B.n473 34.9783
R2402 B.n846 B.n468 34.9783
R2403 B.n852 B.n468 34.9783
R2404 B.n852 B.n469 34.9783
R2405 B.n858 B.n461 34.9783
R2406 B.n864 B.n461 34.9783
R2407 B.n864 B.n457 34.9783
R2408 B.n870 B.n457 34.9783
R2409 B.n870 B.n453 34.9783
R2410 B.n876 B.n453 34.9783
R2411 B.n882 B.n449 34.9783
R2412 B.n882 B.n445 34.9783
R2413 B.n888 B.n445 34.9783
R2414 B.n888 B.n441 34.9783
R2415 B.n894 B.n441 34.9783
R2416 B.n894 B.n437 34.9783
R2417 B.n900 B.n437 34.9783
R2418 B.n906 B.n433 34.9783
R2419 B.n906 B.n429 34.9783
R2420 B.n912 B.n429 34.9783
R2421 B.n912 B.n425 34.9783
R2422 B.n918 B.n425 34.9783
R2423 B.n918 B.n421 34.9783
R2424 B.n924 B.n421 34.9783
R2425 B.n930 B.n417 34.9783
R2426 B.n930 B.n413 34.9783
R2427 B.n936 B.n413 34.9783
R2428 B.n936 B.n409 34.9783
R2429 B.n942 B.n409 34.9783
R2430 B.n942 B.n405 34.9783
R2431 B.n948 B.n405 34.9783
R2432 B.n955 B.n401 34.9783
R2433 B.n955 B.n397 34.9783
R2434 B.n961 B.n397 34.9783
R2435 B.n961 B.n4 34.9783
R2436 B.n1148 B.n4 34.9783
R2437 B.n1148 B.n1147 34.9783
R2438 B.n1147 B.n1146 34.9783
R2439 B.n1146 B.n8 34.9783
R2440 B.n1140 B.n8 34.9783
R2441 B.n1140 B.n1139 34.9783
R2442 B.n1138 B.n15 34.9783
R2443 B.n1132 B.n15 34.9783
R2444 B.n1132 B.n1131 34.9783
R2445 B.n1131 B.n1130 34.9783
R2446 B.n1130 B.n22 34.9783
R2447 B.n1124 B.n22 34.9783
R2448 B.n1124 B.n1123 34.9783
R2449 B.n1122 B.n29 34.9783
R2450 B.n1116 B.n29 34.9783
R2451 B.n1116 B.n1115 34.9783
R2452 B.n1115 B.n1114 34.9783
R2453 B.n1114 B.n36 34.9783
R2454 B.n1108 B.n36 34.9783
R2455 B.n1108 B.n1107 34.9783
R2456 B.n1106 B.n43 34.9783
R2457 B.n1100 B.n43 34.9783
R2458 B.n1100 B.n1099 34.9783
R2459 B.n1099 B.n1098 34.9783
R2460 B.n1098 B.n50 34.9783
R2461 B.n1092 B.n50 34.9783
R2462 B.n1092 B.n1091 34.9783
R2463 B.n1090 B.n57 34.9783
R2464 B.n1084 B.n57 34.9783
R2465 B.n1084 B.n1083 34.9783
R2466 B.n1083 B.n1082 34.9783
R2467 B.n1082 B.n64 34.9783
R2468 B.n1076 B.n64 34.9783
R2469 B.n1075 B.n1074 34.9783
R2470 B.n1074 B.n71 34.9783
R2471 B.n1068 B.n71 34.9783
R2472 B.n1068 B.n1067 34.9783
R2473 B.n1067 B.n1066 34.9783
R2474 B.n1066 B.n78 34.9783
R2475 B.n1060 B.n78 34.9783
R2476 B.n1060 B.n1059 34.9783
R2477 B.n1059 B.n1058 34.9783
R2478 B.n1058 B.n85 34.9783
R2479 B.t11 B.n85 34.9783
R2480 B.t11 B.n1052 34.9783
R2481 B.n1052 B.n1051 34.9783
R2482 B.n1051 B.n92 34.9783
R2483 B.n1045 B.n92 34.9783
R2484 B.n1045 B.n1044 34.9783
R2485 B.n1044 B.n1043 34.9783
R2486 B.n1043 B.n99 34.9783
R2487 B.n1040 B.n1039 34.8103
R2488 B.n1034 B.n1033 34.8103
R2489 B.n569 B.n499 34.8103
R2490 B.n802 B.n801 34.8103
R2491 B.n858 B.t2 32.9208
R2492 B.n1076 B.t8 32.9208
R2493 B.n876 B.t9 31.892
R2494 B.t5 B.n1090 31.892
R2495 B.n900 B.t3 26.7482
R2496 B.t7 B.n1106 26.7482
R2497 B.n924 B.t4 21.6044
R2498 B.t0 B.n1122 21.6044
R2499 B.t6 B.n401 18.5182
R2500 B.n1139 B.t1 18.5182
R2501 B B.n1150 18.0485
R2502 B.n948 B.t6 16.4606
R2503 B.t1 B.n1138 16.4606
R2504 B.t4 B.n417 13.3744
R2505 B.n1123 B.t0 13.3744
R2506 B.n1039 B.n101 10.6151
R2507 B.n168 B.n101 10.6151
R2508 B.n169 B.n168 10.6151
R2509 B.n172 B.n169 10.6151
R2510 B.n173 B.n172 10.6151
R2511 B.n176 B.n173 10.6151
R2512 B.n177 B.n176 10.6151
R2513 B.n180 B.n177 10.6151
R2514 B.n181 B.n180 10.6151
R2515 B.n184 B.n181 10.6151
R2516 B.n185 B.n184 10.6151
R2517 B.n188 B.n185 10.6151
R2518 B.n189 B.n188 10.6151
R2519 B.n192 B.n189 10.6151
R2520 B.n193 B.n192 10.6151
R2521 B.n196 B.n193 10.6151
R2522 B.n197 B.n196 10.6151
R2523 B.n200 B.n197 10.6151
R2524 B.n201 B.n200 10.6151
R2525 B.n204 B.n201 10.6151
R2526 B.n205 B.n204 10.6151
R2527 B.n208 B.n205 10.6151
R2528 B.n209 B.n208 10.6151
R2529 B.n212 B.n209 10.6151
R2530 B.n213 B.n212 10.6151
R2531 B.n216 B.n213 10.6151
R2532 B.n217 B.n216 10.6151
R2533 B.n220 B.n217 10.6151
R2534 B.n221 B.n220 10.6151
R2535 B.n224 B.n221 10.6151
R2536 B.n225 B.n224 10.6151
R2537 B.n228 B.n225 10.6151
R2538 B.n229 B.n228 10.6151
R2539 B.n232 B.n229 10.6151
R2540 B.n233 B.n232 10.6151
R2541 B.n236 B.n233 10.6151
R2542 B.n237 B.n236 10.6151
R2543 B.n240 B.n237 10.6151
R2544 B.n241 B.n240 10.6151
R2545 B.n244 B.n241 10.6151
R2546 B.n245 B.n244 10.6151
R2547 B.n248 B.n245 10.6151
R2548 B.n249 B.n248 10.6151
R2549 B.n252 B.n249 10.6151
R2550 B.n253 B.n252 10.6151
R2551 B.n256 B.n253 10.6151
R2552 B.n257 B.n256 10.6151
R2553 B.n260 B.n257 10.6151
R2554 B.n261 B.n260 10.6151
R2555 B.n264 B.n261 10.6151
R2556 B.n265 B.n264 10.6151
R2557 B.n268 B.n265 10.6151
R2558 B.n269 B.n268 10.6151
R2559 B.n273 B.n272 10.6151
R2560 B.n276 B.n273 10.6151
R2561 B.n277 B.n276 10.6151
R2562 B.n280 B.n277 10.6151
R2563 B.n281 B.n280 10.6151
R2564 B.n284 B.n281 10.6151
R2565 B.n285 B.n284 10.6151
R2566 B.n288 B.n285 10.6151
R2567 B.n293 B.n290 10.6151
R2568 B.n294 B.n293 10.6151
R2569 B.n297 B.n294 10.6151
R2570 B.n298 B.n297 10.6151
R2571 B.n301 B.n298 10.6151
R2572 B.n302 B.n301 10.6151
R2573 B.n305 B.n302 10.6151
R2574 B.n306 B.n305 10.6151
R2575 B.n309 B.n306 10.6151
R2576 B.n310 B.n309 10.6151
R2577 B.n313 B.n310 10.6151
R2578 B.n314 B.n313 10.6151
R2579 B.n317 B.n314 10.6151
R2580 B.n318 B.n317 10.6151
R2581 B.n321 B.n318 10.6151
R2582 B.n322 B.n321 10.6151
R2583 B.n325 B.n322 10.6151
R2584 B.n326 B.n325 10.6151
R2585 B.n329 B.n326 10.6151
R2586 B.n330 B.n329 10.6151
R2587 B.n333 B.n330 10.6151
R2588 B.n334 B.n333 10.6151
R2589 B.n337 B.n334 10.6151
R2590 B.n338 B.n337 10.6151
R2591 B.n341 B.n338 10.6151
R2592 B.n342 B.n341 10.6151
R2593 B.n345 B.n342 10.6151
R2594 B.n346 B.n345 10.6151
R2595 B.n349 B.n346 10.6151
R2596 B.n350 B.n349 10.6151
R2597 B.n353 B.n350 10.6151
R2598 B.n354 B.n353 10.6151
R2599 B.n357 B.n354 10.6151
R2600 B.n358 B.n357 10.6151
R2601 B.n361 B.n358 10.6151
R2602 B.n362 B.n361 10.6151
R2603 B.n365 B.n362 10.6151
R2604 B.n366 B.n365 10.6151
R2605 B.n369 B.n366 10.6151
R2606 B.n370 B.n369 10.6151
R2607 B.n373 B.n370 10.6151
R2608 B.n374 B.n373 10.6151
R2609 B.n377 B.n374 10.6151
R2610 B.n378 B.n377 10.6151
R2611 B.n381 B.n378 10.6151
R2612 B.n382 B.n381 10.6151
R2613 B.n385 B.n382 10.6151
R2614 B.n386 B.n385 10.6151
R2615 B.n389 B.n386 10.6151
R2616 B.n390 B.n389 10.6151
R2617 B.n393 B.n390 10.6151
R2618 B.n394 B.n393 10.6151
R2619 B.n1034 B.n394 10.6151
R2620 B.n807 B.n499 10.6151
R2621 B.n808 B.n807 10.6151
R2622 B.n809 B.n808 10.6151
R2623 B.n809 B.n491 10.6151
R2624 B.n819 B.n491 10.6151
R2625 B.n820 B.n819 10.6151
R2626 B.n821 B.n820 10.6151
R2627 B.n821 B.n483 10.6151
R2628 B.n830 B.n483 10.6151
R2629 B.n831 B.n830 10.6151
R2630 B.n832 B.n831 10.6151
R2631 B.n832 B.n475 10.6151
R2632 B.n842 B.n475 10.6151
R2633 B.n843 B.n842 10.6151
R2634 B.n844 B.n843 10.6151
R2635 B.n844 B.n466 10.6151
R2636 B.n854 B.n466 10.6151
R2637 B.n855 B.n854 10.6151
R2638 B.n856 B.n855 10.6151
R2639 B.n856 B.n459 10.6151
R2640 B.n866 B.n459 10.6151
R2641 B.n867 B.n866 10.6151
R2642 B.n868 B.n867 10.6151
R2643 B.n868 B.n451 10.6151
R2644 B.n878 B.n451 10.6151
R2645 B.n879 B.n878 10.6151
R2646 B.n880 B.n879 10.6151
R2647 B.n880 B.n443 10.6151
R2648 B.n890 B.n443 10.6151
R2649 B.n891 B.n890 10.6151
R2650 B.n892 B.n891 10.6151
R2651 B.n892 B.n435 10.6151
R2652 B.n902 B.n435 10.6151
R2653 B.n903 B.n902 10.6151
R2654 B.n904 B.n903 10.6151
R2655 B.n904 B.n427 10.6151
R2656 B.n914 B.n427 10.6151
R2657 B.n915 B.n914 10.6151
R2658 B.n916 B.n915 10.6151
R2659 B.n916 B.n419 10.6151
R2660 B.n926 B.n419 10.6151
R2661 B.n927 B.n926 10.6151
R2662 B.n928 B.n927 10.6151
R2663 B.n928 B.n411 10.6151
R2664 B.n938 B.n411 10.6151
R2665 B.n939 B.n938 10.6151
R2666 B.n940 B.n939 10.6151
R2667 B.n940 B.n403 10.6151
R2668 B.n950 B.n403 10.6151
R2669 B.n951 B.n950 10.6151
R2670 B.n953 B.n951 10.6151
R2671 B.n953 B.n952 10.6151
R2672 B.n952 B.n395 10.6151
R2673 B.n964 B.n395 10.6151
R2674 B.n965 B.n964 10.6151
R2675 B.n966 B.n965 10.6151
R2676 B.n967 B.n966 10.6151
R2677 B.n969 B.n967 10.6151
R2678 B.n970 B.n969 10.6151
R2679 B.n971 B.n970 10.6151
R2680 B.n972 B.n971 10.6151
R2681 B.n974 B.n972 10.6151
R2682 B.n975 B.n974 10.6151
R2683 B.n976 B.n975 10.6151
R2684 B.n977 B.n976 10.6151
R2685 B.n979 B.n977 10.6151
R2686 B.n980 B.n979 10.6151
R2687 B.n981 B.n980 10.6151
R2688 B.n982 B.n981 10.6151
R2689 B.n984 B.n982 10.6151
R2690 B.n985 B.n984 10.6151
R2691 B.n986 B.n985 10.6151
R2692 B.n987 B.n986 10.6151
R2693 B.n989 B.n987 10.6151
R2694 B.n990 B.n989 10.6151
R2695 B.n991 B.n990 10.6151
R2696 B.n992 B.n991 10.6151
R2697 B.n994 B.n992 10.6151
R2698 B.n995 B.n994 10.6151
R2699 B.n996 B.n995 10.6151
R2700 B.n997 B.n996 10.6151
R2701 B.n999 B.n997 10.6151
R2702 B.n1000 B.n999 10.6151
R2703 B.n1001 B.n1000 10.6151
R2704 B.n1002 B.n1001 10.6151
R2705 B.n1004 B.n1002 10.6151
R2706 B.n1005 B.n1004 10.6151
R2707 B.n1006 B.n1005 10.6151
R2708 B.n1007 B.n1006 10.6151
R2709 B.n1009 B.n1007 10.6151
R2710 B.n1010 B.n1009 10.6151
R2711 B.n1011 B.n1010 10.6151
R2712 B.n1012 B.n1011 10.6151
R2713 B.n1014 B.n1012 10.6151
R2714 B.n1015 B.n1014 10.6151
R2715 B.n1016 B.n1015 10.6151
R2716 B.n1017 B.n1016 10.6151
R2717 B.n1019 B.n1017 10.6151
R2718 B.n1020 B.n1019 10.6151
R2719 B.n1021 B.n1020 10.6151
R2720 B.n1022 B.n1021 10.6151
R2721 B.n1024 B.n1022 10.6151
R2722 B.n1025 B.n1024 10.6151
R2723 B.n1026 B.n1025 10.6151
R2724 B.n1027 B.n1026 10.6151
R2725 B.n1029 B.n1027 10.6151
R2726 B.n1030 B.n1029 10.6151
R2727 B.n1031 B.n1030 10.6151
R2728 B.n1032 B.n1031 10.6151
R2729 B.n1033 B.n1032 10.6151
R2730 B.n801 B.n503 10.6151
R2731 B.n796 B.n503 10.6151
R2732 B.n796 B.n795 10.6151
R2733 B.n795 B.n794 10.6151
R2734 B.n794 B.n791 10.6151
R2735 B.n791 B.n790 10.6151
R2736 B.n790 B.n787 10.6151
R2737 B.n787 B.n786 10.6151
R2738 B.n786 B.n783 10.6151
R2739 B.n783 B.n782 10.6151
R2740 B.n782 B.n779 10.6151
R2741 B.n779 B.n778 10.6151
R2742 B.n778 B.n775 10.6151
R2743 B.n775 B.n774 10.6151
R2744 B.n774 B.n771 10.6151
R2745 B.n771 B.n770 10.6151
R2746 B.n770 B.n767 10.6151
R2747 B.n767 B.n766 10.6151
R2748 B.n766 B.n763 10.6151
R2749 B.n763 B.n762 10.6151
R2750 B.n762 B.n759 10.6151
R2751 B.n759 B.n758 10.6151
R2752 B.n758 B.n755 10.6151
R2753 B.n755 B.n754 10.6151
R2754 B.n754 B.n751 10.6151
R2755 B.n751 B.n750 10.6151
R2756 B.n750 B.n747 10.6151
R2757 B.n747 B.n746 10.6151
R2758 B.n746 B.n743 10.6151
R2759 B.n743 B.n742 10.6151
R2760 B.n742 B.n739 10.6151
R2761 B.n739 B.n738 10.6151
R2762 B.n738 B.n735 10.6151
R2763 B.n735 B.n734 10.6151
R2764 B.n734 B.n731 10.6151
R2765 B.n731 B.n730 10.6151
R2766 B.n730 B.n727 10.6151
R2767 B.n727 B.n726 10.6151
R2768 B.n726 B.n723 10.6151
R2769 B.n723 B.n722 10.6151
R2770 B.n722 B.n719 10.6151
R2771 B.n719 B.n718 10.6151
R2772 B.n718 B.n715 10.6151
R2773 B.n715 B.n714 10.6151
R2774 B.n714 B.n711 10.6151
R2775 B.n711 B.n710 10.6151
R2776 B.n710 B.n707 10.6151
R2777 B.n707 B.n706 10.6151
R2778 B.n706 B.n703 10.6151
R2779 B.n703 B.n702 10.6151
R2780 B.n702 B.n699 10.6151
R2781 B.n699 B.n698 10.6151
R2782 B.n698 B.n695 10.6151
R2783 B.n693 B.n690 10.6151
R2784 B.n690 B.n689 10.6151
R2785 B.n689 B.n686 10.6151
R2786 B.n686 B.n685 10.6151
R2787 B.n685 B.n682 10.6151
R2788 B.n682 B.n681 10.6151
R2789 B.n681 B.n678 10.6151
R2790 B.n678 B.n677 10.6151
R2791 B.n674 B.n673 10.6151
R2792 B.n673 B.n670 10.6151
R2793 B.n670 B.n669 10.6151
R2794 B.n669 B.n666 10.6151
R2795 B.n666 B.n665 10.6151
R2796 B.n665 B.n662 10.6151
R2797 B.n662 B.n661 10.6151
R2798 B.n661 B.n658 10.6151
R2799 B.n658 B.n657 10.6151
R2800 B.n657 B.n654 10.6151
R2801 B.n654 B.n653 10.6151
R2802 B.n653 B.n650 10.6151
R2803 B.n650 B.n649 10.6151
R2804 B.n649 B.n646 10.6151
R2805 B.n646 B.n645 10.6151
R2806 B.n645 B.n642 10.6151
R2807 B.n642 B.n641 10.6151
R2808 B.n641 B.n638 10.6151
R2809 B.n638 B.n637 10.6151
R2810 B.n637 B.n634 10.6151
R2811 B.n634 B.n633 10.6151
R2812 B.n633 B.n630 10.6151
R2813 B.n630 B.n629 10.6151
R2814 B.n629 B.n626 10.6151
R2815 B.n626 B.n625 10.6151
R2816 B.n625 B.n622 10.6151
R2817 B.n622 B.n621 10.6151
R2818 B.n621 B.n618 10.6151
R2819 B.n618 B.n617 10.6151
R2820 B.n617 B.n614 10.6151
R2821 B.n614 B.n613 10.6151
R2822 B.n613 B.n610 10.6151
R2823 B.n610 B.n609 10.6151
R2824 B.n609 B.n606 10.6151
R2825 B.n606 B.n605 10.6151
R2826 B.n605 B.n602 10.6151
R2827 B.n602 B.n601 10.6151
R2828 B.n601 B.n598 10.6151
R2829 B.n598 B.n597 10.6151
R2830 B.n597 B.n594 10.6151
R2831 B.n594 B.n593 10.6151
R2832 B.n593 B.n590 10.6151
R2833 B.n590 B.n589 10.6151
R2834 B.n589 B.n586 10.6151
R2835 B.n586 B.n585 10.6151
R2836 B.n585 B.n582 10.6151
R2837 B.n582 B.n581 10.6151
R2838 B.n581 B.n578 10.6151
R2839 B.n578 B.n577 10.6151
R2840 B.n577 B.n574 10.6151
R2841 B.n574 B.n573 10.6151
R2842 B.n573 B.n570 10.6151
R2843 B.n570 B.n569 10.6151
R2844 B.n803 B.n802 10.6151
R2845 B.n803 B.n495 10.6151
R2846 B.n813 B.n495 10.6151
R2847 B.n814 B.n813 10.6151
R2848 B.n815 B.n814 10.6151
R2849 B.n815 B.n487 10.6151
R2850 B.n824 B.n487 10.6151
R2851 B.n825 B.n824 10.6151
R2852 B.n826 B.n825 10.6151
R2853 B.n826 B.n479 10.6151
R2854 B.n836 B.n479 10.6151
R2855 B.n837 B.n836 10.6151
R2856 B.n838 B.n837 10.6151
R2857 B.n838 B.n471 10.6151
R2858 B.n848 B.n471 10.6151
R2859 B.n849 B.n848 10.6151
R2860 B.n850 B.n849 10.6151
R2861 B.n850 B.n463 10.6151
R2862 B.n860 B.n463 10.6151
R2863 B.n861 B.n860 10.6151
R2864 B.n862 B.n861 10.6151
R2865 B.n862 B.n455 10.6151
R2866 B.n872 B.n455 10.6151
R2867 B.n873 B.n872 10.6151
R2868 B.n874 B.n873 10.6151
R2869 B.n874 B.n447 10.6151
R2870 B.n884 B.n447 10.6151
R2871 B.n885 B.n884 10.6151
R2872 B.n886 B.n885 10.6151
R2873 B.n886 B.n439 10.6151
R2874 B.n896 B.n439 10.6151
R2875 B.n897 B.n896 10.6151
R2876 B.n898 B.n897 10.6151
R2877 B.n898 B.n431 10.6151
R2878 B.n908 B.n431 10.6151
R2879 B.n909 B.n908 10.6151
R2880 B.n910 B.n909 10.6151
R2881 B.n910 B.n423 10.6151
R2882 B.n920 B.n423 10.6151
R2883 B.n921 B.n920 10.6151
R2884 B.n922 B.n921 10.6151
R2885 B.n922 B.n415 10.6151
R2886 B.n932 B.n415 10.6151
R2887 B.n933 B.n932 10.6151
R2888 B.n934 B.n933 10.6151
R2889 B.n934 B.n407 10.6151
R2890 B.n944 B.n407 10.6151
R2891 B.n945 B.n944 10.6151
R2892 B.n946 B.n945 10.6151
R2893 B.n946 B.n399 10.6151
R2894 B.n957 B.n399 10.6151
R2895 B.n958 B.n957 10.6151
R2896 B.n959 B.n958 10.6151
R2897 B.n959 B.n0 10.6151
R2898 B.n1144 B.n1 10.6151
R2899 B.n1144 B.n1143 10.6151
R2900 B.n1143 B.n1142 10.6151
R2901 B.n1142 B.n10 10.6151
R2902 B.n1136 B.n10 10.6151
R2903 B.n1136 B.n1135 10.6151
R2904 B.n1135 B.n1134 10.6151
R2905 B.n1134 B.n17 10.6151
R2906 B.n1128 B.n17 10.6151
R2907 B.n1128 B.n1127 10.6151
R2908 B.n1127 B.n1126 10.6151
R2909 B.n1126 B.n24 10.6151
R2910 B.n1120 B.n24 10.6151
R2911 B.n1120 B.n1119 10.6151
R2912 B.n1119 B.n1118 10.6151
R2913 B.n1118 B.n31 10.6151
R2914 B.n1112 B.n31 10.6151
R2915 B.n1112 B.n1111 10.6151
R2916 B.n1111 B.n1110 10.6151
R2917 B.n1110 B.n38 10.6151
R2918 B.n1104 B.n38 10.6151
R2919 B.n1104 B.n1103 10.6151
R2920 B.n1103 B.n1102 10.6151
R2921 B.n1102 B.n45 10.6151
R2922 B.n1096 B.n45 10.6151
R2923 B.n1096 B.n1095 10.6151
R2924 B.n1095 B.n1094 10.6151
R2925 B.n1094 B.n52 10.6151
R2926 B.n1088 B.n52 10.6151
R2927 B.n1088 B.n1087 10.6151
R2928 B.n1087 B.n1086 10.6151
R2929 B.n1086 B.n59 10.6151
R2930 B.n1080 B.n59 10.6151
R2931 B.n1080 B.n1079 10.6151
R2932 B.n1079 B.n1078 10.6151
R2933 B.n1078 B.n66 10.6151
R2934 B.n1072 B.n66 10.6151
R2935 B.n1072 B.n1071 10.6151
R2936 B.n1071 B.n1070 10.6151
R2937 B.n1070 B.n73 10.6151
R2938 B.n1064 B.n73 10.6151
R2939 B.n1064 B.n1063 10.6151
R2940 B.n1063 B.n1062 10.6151
R2941 B.n1062 B.n80 10.6151
R2942 B.n1056 B.n80 10.6151
R2943 B.n1056 B.n1055 10.6151
R2944 B.n1055 B.n1054 10.6151
R2945 B.n1054 B.n87 10.6151
R2946 B.n1049 B.n87 10.6151
R2947 B.n1049 B.n1048 10.6151
R2948 B.n1048 B.n1047 10.6151
R2949 B.n1047 B.n94 10.6151
R2950 B.n1041 B.n94 10.6151
R2951 B.n1041 B.n1040 10.6151
R2952 B.t3 B.n433 8.23057
R2953 B.n1107 B.t7 8.23057
R2954 B.n272 B.n166 6.5566
R2955 B.n289 B.n288 6.5566
R2956 B.n694 B.n693 6.5566
R2957 B.n677 B.n567 6.5566
R2958 B.n269 B.n166 4.05904
R2959 B.n290 B.n289 4.05904
R2960 B.n695 B.n694 4.05904
R2961 B.n674 B.n567 4.05904
R2962 B.t9 B.n449 3.08678
R2963 B.n1091 B.t5 3.08678
R2964 B.n1150 B.n0 2.81026
R2965 B.n1150 B.n1 2.81026
R2966 B.n469 B.t2 2.05802
R2967 B.t8 B.n1075 2.05802
R2968 VN.n8 VN.t7 198.988
R2969 VN.n45 VN.t5 198.988
R2970 VN.n5 VN.t6 165.919
R2971 VN.n9 VN.t0 165.919
R2972 VN.n27 VN.t2 165.919
R2973 VN.n35 VN.t9 165.919
R2974 VN.n42 VN.t8 165.919
R2975 VN.n46 VN.t1 165.919
R2976 VN.n64 VN.t3 165.919
R2977 VN.n72 VN.t4 165.919
R2978 VN.n71 VN.n37 161.3
R2979 VN.n70 VN.n69 161.3
R2980 VN.n68 VN.n38 161.3
R2981 VN.n67 VN.n66 161.3
R2982 VN.n65 VN.n39 161.3
R2983 VN.n63 VN.n62 161.3
R2984 VN.n61 VN.n40 161.3
R2985 VN.n60 VN.n59 161.3
R2986 VN.n58 VN.n41 161.3
R2987 VN.n57 VN.n56 161.3
R2988 VN.n55 VN.n42 161.3
R2989 VN.n54 VN.n53 161.3
R2990 VN.n52 VN.n43 161.3
R2991 VN.n51 VN.n50 161.3
R2992 VN.n49 VN.n44 161.3
R2993 VN.n48 VN.n47 161.3
R2994 VN.n34 VN.n0 161.3
R2995 VN.n33 VN.n32 161.3
R2996 VN.n31 VN.n1 161.3
R2997 VN.n30 VN.n29 161.3
R2998 VN.n28 VN.n2 161.3
R2999 VN.n26 VN.n25 161.3
R3000 VN.n24 VN.n3 161.3
R3001 VN.n23 VN.n22 161.3
R3002 VN.n21 VN.n4 161.3
R3003 VN.n20 VN.n19 161.3
R3004 VN.n18 VN.n5 161.3
R3005 VN.n17 VN.n16 161.3
R3006 VN.n15 VN.n6 161.3
R3007 VN.n14 VN.n13 161.3
R3008 VN.n12 VN.n7 161.3
R3009 VN.n11 VN.n10 161.3
R3010 VN.n36 VN.n35 94.1189
R3011 VN.n73 VN.n72 94.1189
R3012 VN.n9 VN.n8 63.5395
R3013 VN.n46 VN.n45 63.5395
R3014 VN.n15 VN.n14 56.5193
R3015 VN.n22 VN.n21 56.5193
R3016 VN.n52 VN.n51 56.5193
R3017 VN.n59 VN.n58 56.5193
R3018 VN VN.n73 55.1535
R3019 VN.n33 VN.n1 40.979
R3020 VN.n70 VN.n38 40.979
R3021 VN.n29 VN.n1 40.0078
R3022 VN.n66 VN.n38 40.0078
R3023 VN.n10 VN.n7 24.4675
R3024 VN.n14 VN.n7 24.4675
R3025 VN.n16 VN.n15 24.4675
R3026 VN.n16 VN.n5 24.4675
R3027 VN.n20 VN.n5 24.4675
R3028 VN.n21 VN.n20 24.4675
R3029 VN.n22 VN.n3 24.4675
R3030 VN.n26 VN.n3 24.4675
R3031 VN.n29 VN.n28 24.4675
R3032 VN.n34 VN.n33 24.4675
R3033 VN.n51 VN.n44 24.4675
R3034 VN.n47 VN.n44 24.4675
R3035 VN.n58 VN.n57 24.4675
R3036 VN.n57 VN.n42 24.4675
R3037 VN.n53 VN.n42 24.4675
R3038 VN.n53 VN.n52 24.4675
R3039 VN.n66 VN.n65 24.4675
R3040 VN.n63 VN.n40 24.4675
R3041 VN.n59 VN.n40 24.4675
R3042 VN.n71 VN.n70 24.4675
R3043 VN.n35 VN.n34 16.6381
R3044 VN.n72 VN.n71 16.6381
R3045 VN.n28 VN.n27 16.1487
R3046 VN.n65 VN.n64 16.1487
R3047 VN.n48 VN.n45 9.31187
R3048 VN.n11 VN.n8 9.31187
R3049 VN.n10 VN.n9 8.31928
R3050 VN.n27 VN.n26 8.31928
R3051 VN.n47 VN.n46 8.31928
R3052 VN.n64 VN.n63 8.31928
R3053 VN.n73 VN.n37 0.278367
R3054 VN.n36 VN.n0 0.278367
R3055 VN.n69 VN.n37 0.189894
R3056 VN.n69 VN.n68 0.189894
R3057 VN.n68 VN.n67 0.189894
R3058 VN.n67 VN.n39 0.189894
R3059 VN.n62 VN.n39 0.189894
R3060 VN.n62 VN.n61 0.189894
R3061 VN.n61 VN.n60 0.189894
R3062 VN.n60 VN.n41 0.189894
R3063 VN.n56 VN.n41 0.189894
R3064 VN.n56 VN.n55 0.189894
R3065 VN.n55 VN.n54 0.189894
R3066 VN.n54 VN.n43 0.189894
R3067 VN.n50 VN.n43 0.189894
R3068 VN.n50 VN.n49 0.189894
R3069 VN.n49 VN.n48 0.189894
R3070 VN.n12 VN.n11 0.189894
R3071 VN.n13 VN.n12 0.189894
R3072 VN.n13 VN.n6 0.189894
R3073 VN.n17 VN.n6 0.189894
R3074 VN.n18 VN.n17 0.189894
R3075 VN.n19 VN.n18 0.189894
R3076 VN.n19 VN.n4 0.189894
R3077 VN.n23 VN.n4 0.189894
R3078 VN.n24 VN.n23 0.189894
R3079 VN.n25 VN.n24 0.189894
R3080 VN.n25 VN.n2 0.189894
R3081 VN.n30 VN.n2 0.189894
R3082 VN.n31 VN.n30 0.189894
R3083 VN.n32 VN.n31 0.189894
R3084 VN.n32 VN.n0 0.189894
R3085 VN VN.n36 0.153454
R3086 VDD2.n177 VDD2.n93 289.615
R3087 VDD2.n84 VDD2.n0 289.615
R3088 VDD2.n178 VDD2.n177 185
R3089 VDD2.n176 VDD2.n175 185
R3090 VDD2.n97 VDD2.n96 185
R3091 VDD2.n170 VDD2.n169 185
R3092 VDD2.n168 VDD2.n99 185
R3093 VDD2.n167 VDD2.n166 185
R3094 VDD2.n102 VDD2.n100 185
R3095 VDD2.n161 VDD2.n160 185
R3096 VDD2.n159 VDD2.n158 185
R3097 VDD2.n106 VDD2.n105 185
R3098 VDD2.n153 VDD2.n152 185
R3099 VDD2.n151 VDD2.n150 185
R3100 VDD2.n110 VDD2.n109 185
R3101 VDD2.n145 VDD2.n144 185
R3102 VDD2.n143 VDD2.n142 185
R3103 VDD2.n114 VDD2.n113 185
R3104 VDD2.n137 VDD2.n136 185
R3105 VDD2.n135 VDD2.n134 185
R3106 VDD2.n118 VDD2.n117 185
R3107 VDD2.n129 VDD2.n128 185
R3108 VDD2.n127 VDD2.n126 185
R3109 VDD2.n122 VDD2.n121 185
R3110 VDD2.n28 VDD2.n27 185
R3111 VDD2.n33 VDD2.n32 185
R3112 VDD2.n35 VDD2.n34 185
R3113 VDD2.n24 VDD2.n23 185
R3114 VDD2.n41 VDD2.n40 185
R3115 VDD2.n43 VDD2.n42 185
R3116 VDD2.n20 VDD2.n19 185
R3117 VDD2.n49 VDD2.n48 185
R3118 VDD2.n51 VDD2.n50 185
R3119 VDD2.n16 VDD2.n15 185
R3120 VDD2.n57 VDD2.n56 185
R3121 VDD2.n59 VDD2.n58 185
R3122 VDD2.n12 VDD2.n11 185
R3123 VDD2.n65 VDD2.n64 185
R3124 VDD2.n67 VDD2.n66 185
R3125 VDD2.n8 VDD2.n7 185
R3126 VDD2.n74 VDD2.n73 185
R3127 VDD2.n75 VDD2.n6 185
R3128 VDD2.n77 VDD2.n76 185
R3129 VDD2.n4 VDD2.n3 185
R3130 VDD2.n83 VDD2.n82 185
R3131 VDD2.n85 VDD2.n84 185
R3132 VDD2.n123 VDD2.t5 147.659
R3133 VDD2.n29 VDD2.t2 147.659
R3134 VDD2.n177 VDD2.n176 104.615
R3135 VDD2.n176 VDD2.n96 104.615
R3136 VDD2.n169 VDD2.n96 104.615
R3137 VDD2.n169 VDD2.n168 104.615
R3138 VDD2.n168 VDD2.n167 104.615
R3139 VDD2.n167 VDD2.n100 104.615
R3140 VDD2.n160 VDD2.n100 104.615
R3141 VDD2.n160 VDD2.n159 104.615
R3142 VDD2.n159 VDD2.n105 104.615
R3143 VDD2.n152 VDD2.n105 104.615
R3144 VDD2.n152 VDD2.n151 104.615
R3145 VDD2.n151 VDD2.n109 104.615
R3146 VDD2.n144 VDD2.n109 104.615
R3147 VDD2.n144 VDD2.n143 104.615
R3148 VDD2.n143 VDD2.n113 104.615
R3149 VDD2.n136 VDD2.n113 104.615
R3150 VDD2.n136 VDD2.n135 104.615
R3151 VDD2.n135 VDD2.n117 104.615
R3152 VDD2.n128 VDD2.n117 104.615
R3153 VDD2.n128 VDD2.n127 104.615
R3154 VDD2.n127 VDD2.n121 104.615
R3155 VDD2.n33 VDD2.n27 104.615
R3156 VDD2.n34 VDD2.n33 104.615
R3157 VDD2.n34 VDD2.n23 104.615
R3158 VDD2.n41 VDD2.n23 104.615
R3159 VDD2.n42 VDD2.n41 104.615
R3160 VDD2.n42 VDD2.n19 104.615
R3161 VDD2.n49 VDD2.n19 104.615
R3162 VDD2.n50 VDD2.n49 104.615
R3163 VDD2.n50 VDD2.n15 104.615
R3164 VDD2.n57 VDD2.n15 104.615
R3165 VDD2.n58 VDD2.n57 104.615
R3166 VDD2.n58 VDD2.n11 104.615
R3167 VDD2.n65 VDD2.n11 104.615
R3168 VDD2.n66 VDD2.n65 104.615
R3169 VDD2.n66 VDD2.n7 104.615
R3170 VDD2.n74 VDD2.n7 104.615
R3171 VDD2.n75 VDD2.n74 104.615
R3172 VDD2.n76 VDD2.n75 104.615
R3173 VDD2.n76 VDD2.n3 104.615
R3174 VDD2.n83 VDD2.n3 104.615
R3175 VDD2.n84 VDD2.n83 104.615
R3176 VDD2.n92 VDD2.n91 63.0303
R3177 VDD2 VDD2.n185 63.0275
R3178 VDD2.n184 VDD2.n183 61.3595
R3179 VDD2.n90 VDD2.n89 61.3594
R3180 VDD2.t5 VDD2.n121 52.3082
R3181 VDD2.t2 VDD2.n27 52.3082
R3182 VDD2.n90 VDD2.n88 51.7477
R3183 VDD2.n182 VDD2.n181 49.446
R3184 VDD2.n182 VDD2.n92 48.5364
R3185 VDD2.n123 VDD2.n122 15.6677
R3186 VDD2.n29 VDD2.n28 15.6677
R3187 VDD2.n170 VDD2.n99 13.1884
R3188 VDD2.n77 VDD2.n6 13.1884
R3189 VDD2.n171 VDD2.n97 12.8005
R3190 VDD2.n166 VDD2.n101 12.8005
R3191 VDD2.n126 VDD2.n125 12.8005
R3192 VDD2.n32 VDD2.n31 12.8005
R3193 VDD2.n73 VDD2.n72 12.8005
R3194 VDD2.n78 VDD2.n4 12.8005
R3195 VDD2.n175 VDD2.n174 12.0247
R3196 VDD2.n165 VDD2.n102 12.0247
R3197 VDD2.n129 VDD2.n120 12.0247
R3198 VDD2.n35 VDD2.n26 12.0247
R3199 VDD2.n71 VDD2.n8 12.0247
R3200 VDD2.n82 VDD2.n81 12.0247
R3201 VDD2.n178 VDD2.n95 11.249
R3202 VDD2.n162 VDD2.n161 11.249
R3203 VDD2.n130 VDD2.n118 11.249
R3204 VDD2.n36 VDD2.n24 11.249
R3205 VDD2.n68 VDD2.n67 11.249
R3206 VDD2.n85 VDD2.n2 11.249
R3207 VDD2.n179 VDD2.n93 10.4732
R3208 VDD2.n158 VDD2.n104 10.4732
R3209 VDD2.n134 VDD2.n133 10.4732
R3210 VDD2.n40 VDD2.n39 10.4732
R3211 VDD2.n64 VDD2.n10 10.4732
R3212 VDD2.n86 VDD2.n0 10.4732
R3213 VDD2.n157 VDD2.n106 9.69747
R3214 VDD2.n137 VDD2.n116 9.69747
R3215 VDD2.n43 VDD2.n22 9.69747
R3216 VDD2.n63 VDD2.n12 9.69747
R3217 VDD2.n181 VDD2.n180 9.45567
R3218 VDD2.n88 VDD2.n87 9.45567
R3219 VDD2.n149 VDD2.n148 9.3005
R3220 VDD2.n108 VDD2.n107 9.3005
R3221 VDD2.n155 VDD2.n154 9.3005
R3222 VDD2.n157 VDD2.n156 9.3005
R3223 VDD2.n104 VDD2.n103 9.3005
R3224 VDD2.n163 VDD2.n162 9.3005
R3225 VDD2.n165 VDD2.n164 9.3005
R3226 VDD2.n101 VDD2.n98 9.3005
R3227 VDD2.n180 VDD2.n179 9.3005
R3228 VDD2.n95 VDD2.n94 9.3005
R3229 VDD2.n174 VDD2.n173 9.3005
R3230 VDD2.n172 VDD2.n171 9.3005
R3231 VDD2.n147 VDD2.n146 9.3005
R3232 VDD2.n112 VDD2.n111 9.3005
R3233 VDD2.n141 VDD2.n140 9.3005
R3234 VDD2.n139 VDD2.n138 9.3005
R3235 VDD2.n116 VDD2.n115 9.3005
R3236 VDD2.n133 VDD2.n132 9.3005
R3237 VDD2.n131 VDD2.n130 9.3005
R3238 VDD2.n120 VDD2.n119 9.3005
R3239 VDD2.n125 VDD2.n124 9.3005
R3240 VDD2.n87 VDD2.n86 9.3005
R3241 VDD2.n2 VDD2.n1 9.3005
R3242 VDD2.n81 VDD2.n80 9.3005
R3243 VDD2.n79 VDD2.n78 9.3005
R3244 VDD2.n18 VDD2.n17 9.3005
R3245 VDD2.n47 VDD2.n46 9.3005
R3246 VDD2.n45 VDD2.n44 9.3005
R3247 VDD2.n22 VDD2.n21 9.3005
R3248 VDD2.n39 VDD2.n38 9.3005
R3249 VDD2.n37 VDD2.n36 9.3005
R3250 VDD2.n26 VDD2.n25 9.3005
R3251 VDD2.n31 VDD2.n30 9.3005
R3252 VDD2.n53 VDD2.n52 9.3005
R3253 VDD2.n55 VDD2.n54 9.3005
R3254 VDD2.n14 VDD2.n13 9.3005
R3255 VDD2.n61 VDD2.n60 9.3005
R3256 VDD2.n63 VDD2.n62 9.3005
R3257 VDD2.n10 VDD2.n9 9.3005
R3258 VDD2.n69 VDD2.n68 9.3005
R3259 VDD2.n71 VDD2.n70 9.3005
R3260 VDD2.n72 VDD2.n5 9.3005
R3261 VDD2.n154 VDD2.n153 8.92171
R3262 VDD2.n138 VDD2.n114 8.92171
R3263 VDD2.n44 VDD2.n20 8.92171
R3264 VDD2.n60 VDD2.n59 8.92171
R3265 VDD2.n150 VDD2.n108 8.14595
R3266 VDD2.n142 VDD2.n141 8.14595
R3267 VDD2.n48 VDD2.n47 8.14595
R3268 VDD2.n56 VDD2.n14 8.14595
R3269 VDD2.n149 VDD2.n110 7.3702
R3270 VDD2.n145 VDD2.n112 7.3702
R3271 VDD2.n51 VDD2.n18 7.3702
R3272 VDD2.n55 VDD2.n16 7.3702
R3273 VDD2.n146 VDD2.n110 6.59444
R3274 VDD2.n146 VDD2.n145 6.59444
R3275 VDD2.n52 VDD2.n51 6.59444
R3276 VDD2.n52 VDD2.n16 6.59444
R3277 VDD2.n150 VDD2.n149 5.81868
R3278 VDD2.n142 VDD2.n112 5.81868
R3279 VDD2.n48 VDD2.n18 5.81868
R3280 VDD2.n56 VDD2.n55 5.81868
R3281 VDD2.n153 VDD2.n108 5.04292
R3282 VDD2.n141 VDD2.n114 5.04292
R3283 VDD2.n47 VDD2.n20 5.04292
R3284 VDD2.n59 VDD2.n14 5.04292
R3285 VDD2.n124 VDD2.n123 4.38563
R3286 VDD2.n30 VDD2.n29 4.38563
R3287 VDD2.n154 VDD2.n106 4.26717
R3288 VDD2.n138 VDD2.n137 4.26717
R3289 VDD2.n44 VDD2.n43 4.26717
R3290 VDD2.n60 VDD2.n12 4.26717
R3291 VDD2.n181 VDD2.n93 3.49141
R3292 VDD2.n158 VDD2.n157 3.49141
R3293 VDD2.n134 VDD2.n116 3.49141
R3294 VDD2.n40 VDD2.n22 3.49141
R3295 VDD2.n64 VDD2.n63 3.49141
R3296 VDD2.n88 VDD2.n0 3.49141
R3297 VDD2.n179 VDD2.n178 2.71565
R3298 VDD2.n161 VDD2.n104 2.71565
R3299 VDD2.n133 VDD2.n118 2.71565
R3300 VDD2.n39 VDD2.n24 2.71565
R3301 VDD2.n67 VDD2.n10 2.71565
R3302 VDD2.n86 VDD2.n85 2.71565
R3303 VDD2.n184 VDD2.n182 2.30222
R3304 VDD2.n175 VDD2.n95 1.93989
R3305 VDD2.n162 VDD2.n102 1.93989
R3306 VDD2.n130 VDD2.n129 1.93989
R3307 VDD2.n36 VDD2.n35 1.93989
R3308 VDD2.n68 VDD2.n8 1.93989
R3309 VDD2.n82 VDD2.n2 1.93989
R3310 VDD2.n185 VDD2.t8 1.22955
R3311 VDD2.n185 VDD2.t4 1.22955
R3312 VDD2.n183 VDD2.t6 1.22955
R3313 VDD2.n183 VDD2.t1 1.22955
R3314 VDD2.n91 VDD2.t7 1.22955
R3315 VDD2.n91 VDD2.t0 1.22955
R3316 VDD2.n89 VDD2.t9 1.22955
R3317 VDD2.n89 VDD2.t3 1.22955
R3318 VDD2.n174 VDD2.n97 1.16414
R3319 VDD2.n166 VDD2.n165 1.16414
R3320 VDD2.n126 VDD2.n120 1.16414
R3321 VDD2.n32 VDD2.n26 1.16414
R3322 VDD2.n73 VDD2.n71 1.16414
R3323 VDD2.n81 VDD2.n4 1.16414
R3324 VDD2 VDD2.n184 0.634121
R3325 VDD2.n92 VDD2.n90 0.520585
R3326 VDD2.n171 VDD2.n170 0.388379
R3327 VDD2.n101 VDD2.n99 0.388379
R3328 VDD2.n125 VDD2.n122 0.388379
R3329 VDD2.n31 VDD2.n28 0.388379
R3330 VDD2.n72 VDD2.n6 0.388379
R3331 VDD2.n78 VDD2.n77 0.388379
R3332 VDD2.n180 VDD2.n94 0.155672
R3333 VDD2.n173 VDD2.n94 0.155672
R3334 VDD2.n173 VDD2.n172 0.155672
R3335 VDD2.n172 VDD2.n98 0.155672
R3336 VDD2.n164 VDD2.n98 0.155672
R3337 VDD2.n164 VDD2.n163 0.155672
R3338 VDD2.n163 VDD2.n103 0.155672
R3339 VDD2.n156 VDD2.n103 0.155672
R3340 VDD2.n156 VDD2.n155 0.155672
R3341 VDD2.n155 VDD2.n107 0.155672
R3342 VDD2.n148 VDD2.n107 0.155672
R3343 VDD2.n148 VDD2.n147 0.155672
R3344 VDD2.n147 VDD2.n111 0.155672
R3345 VDD2.n140 VDD2.n111 0.155672
R3346 VDD2.n140 VDD2.n139 0.155672
R3347 VDD2.n139 VDD2.n115 0.155672
R3348 VDD2.n132 VDD2.n115 0.155672
R3349 VDD2.n132 VDD2.n131 0.155672
R3350 VDD2.n131 VDD2.n119 0.155672
R3351 VDD2.n124 VDD2.n119 0.155672
R3352 VDD2.n30 VDD2.n25 0.155672
R3353 VDD2.n37 VDD2.n25 0.155672
R3354 VDD2.n38 VDD2.n37 0.155672
R3355 VDD2.n38 VDD2.n21 0.155672
R3356 VDD2.n45 VDD2.n21 0.155672
R3357 VDD2.n46 VDD2.n45 0.155672
R3358 VDD2.n46 VDD2.n17 0.155672
R3359 VDD2.n53 VDD2.n17 0.155672
R3360 VDD2.n54 VDD2.n53 0.155672
R3361 VDD2.n54 VDD2.n13 0.155672
R3362 VDD2.n61 VDD2.n13 0.155672
R3363 VDD2.n62 VDD2.n61 0.155672
R3364 VDD2.n62 VDD2.n9 0.155672
R3365 VDD2.n69 VDD2.n9 0.155672
R3366 VDD2.n70 VDD2.n69 0.155672
R3367 VDD2.n70 VDD2.n5 0.155672
R3368 VDD2.n79 VDD2.n5 0.155672
R3369 VDD2.n80 VDD2.n79 0.155672
R3370 VDD2.n80 VDD2.n1 0.155672
R3371 VDD2.n87 VDD2.n1 0.155672
C0 VDD1 VDD2 2.00473f
C1 VDD1 VN 0.15262f
C2 VDD2 VN 13.838099f
C3 VDD1 VTAIL 12.367901f
C4 VDD2 VTAIL 12.4158f
C5 VN VTAIL 14.1912f
C6 VDD1 VP 14.231501f
C7 VDD2 VP 0.550629f
C8 VN VP 8.77472f
C9 VTAIL VP 14.2055f
C10 VDD2 B 7.634338f
C11 VDD1 B 7.605136f
C12 VTAIL B 9.624571f
C13 VN B 17.26358f
C14 VP B 15.692297f
C15 VDD2.n0 B 0.031701f
C16 VDD2.n1 B 0.023572f
C17 VDD2.n2 B 0.012666f
C18 VDD2.n3 B 0.029939f
C19 VDD2.n4 B 0.013411f
C20 VDD2.n5 B 0.023572f
C21 VDD2.n6 B 0.013039f
C22 VDD2.n7 B 0.029939f
C23 VDD2.n8 B 0.013411f
C24 VDD2.n9 B 0.023572f
C25 VDD2.n10 B 0.012666f
C26 VDD2.n11 B 0.029939f
C27 VDD2.n12 B 0.013411f
C28 VDD2.n13 B 0.023572f
C29 VDD2.n14 B 0.012666f
C30 VDD2.n15 B 0.029939f
C31 VDD2.n16 B 0.013411f
C32 VDD2.n17 B 0.023572f
C33 VDD2.n18 B 0.012666f
C34 VDD2.n19 B 0.029939f
C35 VDD2.n20 B 0.013411f
C36 VDD2.n21 B 0.023572f
C37 VDD2.n22 B 0.012666f
C38 VDD2.n23 B 0.029939f
C39 VDD2.n24 B 0.013411f
C40 VDD2.n25 B 0.023572f
C41 VDD2.n26 B 0.012666f
C42 VDD2.n27 B 0.022454f
C43 VDD2.n28 B 0.017686f
C44 VDD2.t2 B 0.049455f
C45 VDD2.n29 B 0.160299f
C46 VDD2.n30 B 1.65351f
C47 VDD2.n31 B 0.012666f
C48 VDD2.n32 B 0.013411f
C49 VDD2.n33 B 0.029939f
C50 VDD2.n34 B 0.029939f
C51 VDD2.n35 B 0.013411f
C52 VDD2.n36 B 0.012666f
C53 VDD2.n37 B 0.023572f
C54 VDD2.n38 B 0.023572f
C55 VDD2.n39 B 0.012666f
C56 VDD2.n40 B 0.013411f
C57 VDD2.n41 B 0.029939f
C58 VDD2.n42 B 0.029939f
C59 VDD2.n43 B 0.013411f
C60 VDD2.n44 B 0.012666f
C61 VDD2.n45 B 0.023572f
C62 VDD2.n46 B 0.023572f
C63 VDD2.n47 B 0.012666f
C64 VDD2.n48 B 0.013411f
C65 VDD2.n49 B 0.029939f
C66 VDD2.n50 B 0.029939f
C67 VDD2.n51 B 0.013411f
C68 VDD2.n52 B 0.012666f
C69 VDD2.n53 B 0.023572f
C70 VDD2.n54 B 0.023572f
C71 VDD2.n55 B 0.012666f
C72 VDD2.n56 B 0.013411f
C73 VDD2.n57 B 0.029939f
C74 VDD2.n58 B 0.029939f
C75 VDD2.n59 B 0.013411f
C76 VDD2.n60 B 0.012666f
C77 VDD2.n61 B 0.023572f
C78 VDD2.n62 B 0.023572f
C79 VDD2.n63 B 0.012666f
C80 VDD2.n64 B 0.013411f
C81 VDD2.n65 B 0.029939f
C82 VDD2.n66 B 0.029939f
C83 VDD2.n67 B 0.013411f
C84 VDD2.n68 B 0.012666f
C85 VDD2.n69 B 0.023572f
C86 VDD2.n70 B 0.023572f
C87 VDD2.n71 B 0.012666f
C88 VDD2.n72 B 0.012666f
C89 VDD2.n73 B 0.013411f
C90 VDD2.n74 B 0.029939f
C91 VDD2.n75 B 0.029939f
C92 VDD2.n76 B 0.029939f
C93 VDD2.n77 B 0.013039f
C94 VDD2.n78 B 0.012666f
C95 VDD2.n79 B 0.023572f
C96 VDD2.n80 B 0.023572f
C97 VDD2.n81 B 0.012666f
C98 VDD2.n82 B 0.013411f
C99 VDD2.n83 B 0.029939f
C100 VDD2.n84 B 0.062281f
C101 VDD2.n85 B 0.013411f
C102 VDD2.n86 B 0.012666f
C103 VDD2.n87 B 0.05545f
C104 VDD2.n88 B 0.060706f
C105 VDD2.t9 B 0.30008f
C106 VDD2.t3 B 0.30008f
C107 VDD2.n89 B 2.72169f
C108 VDD2.n90 B 0.619918f
C109 VDD2.t7 B 0.30008f
C110 VDD2.t0 B 0.30008f
C111 VDD2.n91 B 2.73508f
C112 VDD2.n92 B 2.85196f
C113 VDD2.n93 B 0.031701f
C114 VDD2.n94 B 0.023572f
C115 VDD2.n95 B 0.012666f
C116 VDD2.n96 B 0.029939f
C117 VDD2.n97 B 0.013411f
C118 VDD2.n98 B 0.023572f
C119 VDD2.n99 B 0.013039f
C120 VDD2.n100 B 0.029939f
C121 VDD2.n101 B 0.012666f
C122 VDD2.n102 B 0.013411f
C123 VDD2.n103 B 0.023572f
C124 VDD2.n104 B 0.012666f
C125 VDD2.n105 B 0.029939f
C126 VDD2.n106 B 0.013411f
C127 VDD2.n107 B 0.023572f
C128 VDD2.n108 B 0.012666f
C129 VDD2.n109 B 0.029939f
C130 VDD2.n110 B 0.013411f
C131 VDD2.n111 B 0.023572f
C132 VDD2.n112 B 0.012666f
C133 VDD2.n113 B 0.029939f
C134 VDD2.n114 B 0.013411f
C135 VDD2.n115 B 0.023572f
C136 VDD2.n116 B 0.012666f
C137 VDD2.n117 B 0.029939f
C138 VDD2.n118 B 0.013411f
C139 VDD2.n119 B 0.023572f
C140 VDD2.n120 B 0.012666f
C141 VDD2.n121 B 0.022454f
C142 VDD2.n122 B 0.017686f
C143 VDD2.t5 B 0.049455f
C144 VDD2.n123 B 0.160299f
C145 VDD2.n124 B 1.65351f
C146 VDD2.n125 B 0.012666f
C147 VDD2.n126 B 0.013411f
C148 VDD2.n127 B 0.029939f
C149 VDD2.n128 B 0.029939f
C150 VDD2.n129 B 0.013411f
C151 VDD2.n130 B 0.012666f
C152 VDD2.n131 B 0.023572f
C153 VDD2.n132 B 0.023572f
C154 VDD2.n133 B 0.012666f
C155 VDD2.n134 B 0.013411f
C156 VDD2.n135 B 0.029939f
C157 VDD2.n136 B 0.029939f
C158 VDD2.n137 B 0.013411f
C159 VDD2.n138 B 0.012666f
C160 VDD2.n139 B 0.023572f
C161 VDD2.n140 B 0.023572f
C162 VDD2.n141 B 0.012666f
C163 VDD2.n142 B 0.013411f
C164 VDD2.n143 B 0.029939f
C165 VDD2.n144 B 0.029939f
C166 VDD2.n145 B 0.013411f
C167 VDD2.n146 B 0.012666f
C168 VDD2.n147 B 0.023572f
C169 VDD2.n148 B 0.023572f
C170 VDD2.n149 B 0.012666f
C171 VDD2.n150 B 0.013411f
C172 VDD2.n151 B 0.029939f
C173 VDD2.n152 B 0.029939f
C174 VDD2.n153 B 0.013411f
C175 VDD2.n154 B 0.012666f
C176 VDD2.n155 B 0.023572f
C177 VDD2.n156 B 0.023572f
C178 VDD2.n157 B 0.012666f
C179 VDD2.n158 B 0.013411f
C180 VDD2.n159 B 0.029939f
C181 VDD2.n160 B 0.029939f
C182 VDD2.n161 B 0.013411f
C183 VDD2.n162 B 0.012666f
C184 VDD2.n163 B 0.023572f
C185 VDD2.n164 B 0.023572f
C186 VDD2.n165 B 0.012666f
C187 VDD2.n166 B 0.013411f
C188 VDD2.n167 B 0.029939f
C189 VDD2.n168 B 0.029939f
C190 VDD2.n169 B 0.029939f
C191 VDD2.n170 B 0.013039f
C192 VDD2.n171 B 0.012666f
C193 VDD2.n172 B 0.023572f
C194 VDD2.n173 B 0.023572f
C195 VDD2.n174 B 0.012666f
C196 VDD2.n175 B 0.013411f
C197 VDD2.n176 B 0.029939f
C198 VDD2.n177 B 0.062281f
C199 VDD2.n178 B 0.013411f
C200 VDD2.n179 B 0.012666f
C201 VDD2.n180 B 0.05545f
C202 VDD2.n181 B 0.050886f
C203 VDD2.n182 B 2.92707f
C204 VDD2.t6 B 0.30008f
C205 VDD2.t1 B 0.30008f
C206 VDD2.n183 B 2.72169f
C207 VDD2.n184 B 0.416537f
C208 VDD2.t8 B 0.30008f
C209 VDD2.t4 B 0.30008f
C210 VDD2.n185 B 2.73504f
C211 VN.n0 B 0.029369f
C212 VN.t9 B 2.30466f
C213 VN.n1 B 0.018016f
C214 VN.n2 B 0.022276f
C215 VN.t2 B 2.30466f
C216 VN.n3 B 0.041517f
C217 VN.n4 B 0.022276f
C218 VN.t6 B 2.30466f
C219 VN.n5 B 0.825968f
C220 VN.n6 B 0.022276f
C221 VN.n7 B 0.041517f
C222 VN.t7 B 2.45953f
C223 VN.n8 B 0.852415f
C224 VN.t0 B 2.30466f
C225 VN.n9 B 0.861756f
C226 VN.n10 B 0.027989f
C227 VN.n11 B 0.192676f
C228 VN.n12 B 0.022276f
C229 VN.n13 B 0.022276f
C230 VN.n14 B 0.027245f
C231 VN.n15 B 0.037797f
C232 VN.n16 B 0.041517f
C233 VN.n17 B 0.022276f
C234 VN.n18 B 0.022276f
C235 VN.n19 B 0.022276f
C236 VN.n20 B 0.041517f
C237 VN.n21 B 0.037797f
C238 VN.n22 B 0.027245f
C239 VN.n23 B 0.022276f
C240 VN.n24 B 0.022276f
C241 VN.n25 B 0.022276f
C242 VN.n26 B 0.027989f
C243 VN.n27 B 0.804948f
C244 VN.n28 B 0.034548f
C245 VN.n29 B 0.044383f
C246 VN.n30 B 0.022276f
C247 VN.n31 B 0.022276f
C248 VN.n32 B 0.022276f
C249 VN.n33 B 0.04416f
C250 VN.n34 B 0.034958f
C251 VN.n35 B 0.880252f
C252 VN.n36 B 0.030554f
C253 VN.n37 B 0.029369f
C254 VN.t4 B 2.30466f
C255 VN.n38 B 0.018016f
C256 VN.n39 B 0.022276f
C257 VN.t3 B 2.30466f
C258 VN.n40 B 0.041517f
C259 VN.n41 B 0.022276f
C260 VN.t8 B 2.30466f
C261 VN.n42 B 0.825968f
C262 VN.n43 B 0.022276f
C263 VN.n44 B 0.041517f
C264 VN.t5 B 2.45953f
C265 VN.n45 B 0.852415f
C266 VN.t1 B 2.30466f
C267 VN.n46 B 0.861756f
C268 VN.n47 B 0.027989f
C269 VN.n48 B 0.192676f
C270 VN.n49 B 0.022276f
C271 VN.n50 B 0.022276f
C272 VN.n51 B 0.027245f
C273 VN.n52 B 0.037797f
C274 VN.n53 B 0.041517f
C275 VN.n54 B 0.022276f
C276 VN.n55 B 0.022276f
C277 VN.n56 B 0.022276f
C278 VN.n57 B 0.041517f
C279 VN.n58 B 0.037797f
C280 VN.n59 B 0.027245f
C281 VN.n60 B 0.022276f
C282 VN.n61 B 0.022276f
C283 VN.n62 B 0.022276f
C284 VN.n63 B 0.027989f
C285 VN.n64 B 0.804948f
C286 VN.n65 B 0.034548f
C287 VN.n66 B 0.044383f
C288 VN.n67 B 0.022276f
C289 VN.n68 B 0.022276f
C290 VN.n69 B 0.022276f
C291 VN.n70 B 0.04416f
C292 VN.n71 B 0.034958f
C293 VN.n72 B 0.880252f
C294 VN.n73 B 1.42323f
C295 VTAIL.t1 B 0.304009f
C296 VTAIL.t0 B 0.304009f
C297 VTAIL.n0 B 2.68581f
C298 VTAIL.n1 B 0.497214f
C299 VTAIL.n2 B 0.032116f
C300 VTAIL.n3 B 0.02388f
C301 VTAIL.n4 B 0.012832f
C302 VTAIL.n5 B 0.030331f
C303 VTAIL.n6 B 0.013587f
C304 VTAIL.n7 B 0.02388f
C305 VTAIL.n8 B 0.01321f
C306 VTAIL.n9 B 0.030331f
C307 VTAIL.n10 B 0.013587f
C308 VTAIL.n11 B 0.02388f
C309 VTAIL.n12 B 0.012832f
C310 VTAIL.n13 B 0.030331f
C311 VTAIL.n14 B 0.013587f
C312 VTAIL.n15 B 0.02388f
C313 VTAIL.n16 B 0.012832f
C314 VTAIL.n17 B 0.030331f
C315 VTAIL.n18 B 0.013587f
C316 VTAIL.n19 B 0.02388f
C317 VTAIL.n20 B 0.012832f
C318 VTAIL.n21 B 0.030331f
C319 VTAIL.n22 B 0.013587f
C320 VTAIL.n23 B 0.02388f
C321 VTAIL.n24 B 0.012832f
C322 VTAIL.n25 B 0.030331f
C323 VTAIL.n26 B 0.013587f
C324 VTAIL.n27 B 0.02388f
C325 VTAIL.n28 B 0.012832f
C326 VTAIL.n29 B 0.022748f
C327 VTAIL.n30 B 0.017917f
C328 VTAIL.t16 B 0.050102f
C329 VTAIL.n31 B 0.162398f
C330 VTAIL.n32 B 1.67516f
C331 VTAIL.n33 B 0.012832f
C332 VTAIL.n34 B 0.013587f
C333 VTAIL.n35 B 0.030331f
C334 VTAIL.n36 B 0.030331f
C335 VTAIL.n37 B 0.013587f
C336 VTAIL.n38 B 0.012832f
C337 VTAIL.n39 B 0.02388f
C338 VTAIL.n40 B 0.02388f
C339 VTAIL.n41 B 0.012832f
C340 VTAIL.n42 B 0.013587f
C341 VTAIL.n43 B 0.030331f
C342 VTAIL.n44 B 0.030331f
C343 VTAIL.n45 B 0.013587f
C344 VTAIL.n46 B 0.012832f
C345 VTAIL.n47 B 0.02388f
C346 VTAIL.n48 B 0.02388f
C347 VTAIL.n49 B 0.012832f
C348 VTAIL.n50 B 0.013587f
C349 VTAIL.n51 B 0.030331f
C350 VTAIL.n52 B 0.030331f
C351 VTAIL.n53 B 0.013587f
C352 VTAIL.n54 B 0.012832f
C353 VTAIL.n55 B 0.02388f
C354 VTAIL.n56 B 0.02388f
C355 VTAIL.n57 B 0.012832f
C356 VTAIL.n58 B 0.013587f
C357 VTAIL.n59 B 0.030331f
C358 VTAIL.n60 B 0.030331f
C359 VTAIL.n61 B 0.013587f
C360 VTAIL.n62 B 0.012832f
C361 VTAIL.n63 B 0.02388f
C362 VTAIL.n64 B 0.02388f
C363 VTAIL.n65 B 0.012832f
C364 VTAIL.n66 B 0.013587f
C365 VTAIL.n67 B 0.030331f
C366 VTAIL.n68 B 0.030331f
C367 VTAIL.n69 B 0.013587f
C368 VTAIL.n70 B 0.012832f
C369 VTAIL.n71 B 0.02388f
C370 VTAIL.n72 B 0.02388f
C371 VTAIL.n73 B 0.012832f
C372 VTAIL.n74 B 0.012832f
C373 VTAIL.n75 B 0.013587f
C374 VTAIL.n76 B 0.030331f
C375 VTAIL.n77 B 0.030331f
C376 VTAIL.n78 B 0.030331f
C377 VTAIL.n79 B 0.01321f
C378 VTAIL.n80 B 0.012832f
C379 VTAIL.n81 B 0.02388f
C380 VTAIL.n82 B 0.02388f
C381 VTAIL.n83 B 0.012832f
C382 VTAIL.n84 B 0.013587f
C383 VTAIL.n85 B 0.030331f
C384 VTAIL.n86 B 0.063096f
C385 VTAIL.n87 B 0.013587f
C386 VTAIL.n88 B 0.012832f
C387 VTAIL.n89 B 0.056177f
C388 VTAIL.n90 B 0.035071f
C389 VTAIL.n91 B 0.322767f
C390 VTAIL.t15 B 0.304009f
C391 VTAIL.t10 B 0.304009f
C392 VTAIL.n92 B 2.68581f
C393 VTAIL.n93 B 0.589418f
C394 VTAIL.t13 B 0.304009f
C395 VTAIL.t19 B 0.304009f
C396 VTAIL.n94 B 2.68581f
C397 VTAIL.n95 B 2.15955f
C398 VTAIL.t2 B 0.304009f
C399 VTAIL.t9 B 0.304009f
C400 VTAIL.n96 B 2.68582f
C401 VTAIL.n97 B 2.15954f
C402 VTAIL.t3 B 0.304009f
C403 VTAIL.t4 B 0.304009f
C404 VTAIL.n98 B 2.68582f
C405 VTAIL.n99 B 0.589405f
C406 VTAIL.n100 B 0.032116f
C407 VTAIL.n101 B 0.02388f
C408 VTAIL.n102 B 0.012832f
C409 VTAIL.n103 B 0.030331f
C410 VTAIL.n104 B 0.013587f
C411 VTAIL.n105 B 0.02388f
C412 VTAIL.n106 B 0.01321f
C413 VTAIL.n107 B 0.030331f
C414 VTAIL.n108 B 0.012832f
C415 VTAIL.n109 B 0.013587f
C416 VTAIL.n110 B 0.02388f
C417 VTAIL.n111 B 0.012832f
C418 VTAIL.n112 B 0.030331f
C419 VTAIL.n113 B 0.013587f
C420 VTAIL.n114 B 0.02388f
C421 VTAIL.n115 B 0.012832f
C422 VTAIL.n116 B 0.030331f
C423 VTAIL.n117 B 0.013587f
C424 VTAIL.n118 B 0.02388f
C425 VTAIL.n119 B 0.012832f
C426 VTAIL.n120 B 0.030331f
C427 VTAIL.n121 B 0.013587f
C428 VTAIL.n122 B 0.02388f
C429 VTAIL.n123 B 0.012832f
C430 VTAIL.n124 B 0.030331f
C431 VTAIL.n125 B 0.013587f
C432 VTAIL.n126 B 0.02388f
C433 VTAIL.n127 B 0.012832f
C434 VTAIL.n128 B 0.022748f
C435 VTAIL.n129 B 0.017917f
C436 VTAIL.t6 B 0.050102f
C437 VTAIL.n130 B 0.162398f
C438 VTAIL.n131 B 1.67516f
C439 VTAIL.n132 B 0.012832f
C440 VTAIL.n133 B 0.013587f
C441 VTAIL.n134 B 0.030331f
C442 VTAIL.n135 B 0.030331f
C443 VTAIL.n136 B 0.013587f
C444 VTAIL.n137 B 0.012832f
C445 VTAIL.n138 B 0.02388f
C446 VTAIL.n139 B 0.02388f
C447 VTAIL.n140 B 0.012832f
C448 VTAIL.n141 B 0.013587f
C449 VTAIL.n142 B 0.030331f
C450 VTAIL.n143 B 0.030331f
C451 VTAIL.n144 B 0.013587f
C452 VTAIL.n145 B 0.012832f
C453 VTAIL.n146 B 0.02388f
C454 VTAIL.n147 B 0.02388f
C455 VTAIL.n148 B 0.012832f
C456 VTAIL.n149 B 0.013587f
C457 VTAIL.n150 B 0.030331f
C458 VTAIL.n151 B 0.030331f
C459 VTAIL.n152 B 0.013587f
C460 VTAIL.n153 B 0.012832f
C461 VTAIL.n154 B 0.02388f
C462 VTAIL.n155 B 0.02388f
C463 VTAIL.n156 B 0.012832f
C464 VTAIL.n157 B 0.013587f
C465 VTAIL.n158 B 0.030331f
C466 VTAIL.n159 B 0.030331f
C467 VTAIL.n160 B 0.013587f
C468 VTAIL.n161 B 0.012832f
C469 VTAIL.n162 B 0.02388f
C470 VTAIL.n163 B 0.02388f
C471 VTAIL.n164 B 0.012832f
C472 VTAIL.n165 B 0.013587f
C473 VTAIL.n166 B 0.030331f
C474 VTAIL.n167 B 0.030331f
C475 VTAIL.n168 B 0.013587f
C476 VTAIL.n169 B 0.012832f
C477 VTAIL.n170 B 0.02388f
C478 VTAIL.n171 B 0.02388f
C479 VTAIL.n172 B 0.012832f
C480 VTAIL.n173 B 0.013587f
C481 VTAIL.n174 B 0.030331f
C482 VTAIL.n175 B 0.030331f
C483 VTAIL.n176 B 0.030331f
C484 VTAIL.n177 B 0.01321f
C485 VTAIL.n178 B 0.012832f
C486 VTAIL.n179 B 0.02388f
C487 VTAIL.n180 B 0.02388f
C488 VTAIL.n181 B 0.012832f
C489 VTAIL.n182 B 0.013587f
C490 VTAIL.n183 B 0.030331f
C491 VTAIL.n184 B 0.063096f
C492 VTAIL.n185 B 0.013587f
C493 VTAIL.n186 B 0.012832f
C494 VTAIL.n187 B 0.056177f
C495 VTAIL.n188 B 0.035071f
C496 VTAIL.n189 B 0.322767f
C497 VTAIL.t14 B 0.304009f
C498 VTAIL.t11 B 0.304009f
C499 VTAIL.n190 B 2.68582f
C500 VTAIL.n191 B 0.537001f
C501 VTAIL.t17 B 0.304009f
C502 VTAIL.t12 B 0.304009f
C503 VTAIL.n192 B 2.68582f
C504 VTAIL.n193 B 0.589405f
C505 VTAIL.n194 B 0.032116f
C506 VTAIL.n195 B 0.02388f
C507 VTAIL.n196 B 0.012832f
C508 VTAIL.n197 B 0.030331f
C509 VTAIL.n198 B 0.013587f
C510 VTAIL.n199 B 0.02388f
C511 VTAIL.n200 B 0.01321f
C512 VTAIL.n201 B 0.030331f
C513 VTAIL.n202 B 0.012832f
C514 VTAIL.n203 B 0.013587f
C515 VTAIL.n204 B 0.02388f
C516 VTAIL.n205 B 0.012832f
C517 VTAIL.n206 B 0.030331f
C518 VTAIL.n207 B 0.013587f
C519 VTAIL.n208 B 0.02388f
C520 VTAIL.n209 B 0.012832f
C521 VTAIL.n210 B 0.030331f
C522 VTAIL.n211 B 0.013587f
C523 VTAIL.n212 B 0.02388f
C524 VTAIL.n213 B 0.012832f
C525 VTAIL.n214 B 0.030331f
C526 VTAIL.n215 B 0.013587f
C527 VTAIL.n216 B 0.02388f
C528 VTAIL.n217 B 0.012832f
C529 VTAIL.n218 B 0.030331f
C530 VTAIL.n219 B 0.013587f
C531 VTAIL.n220 B 0.02388f
C532 VTAIL.n221 B 0.012832f
C533 VTAIL.n222 B 0.022748f
C534 VTAIL.n223 B 0.017917f
C535 VTAIL.t18 B 0.050102f
C536 VTAIL.n224 B 0.162398f
C537 VTAIL.n225 B 1.67516f
C538 VTAIL.n226 B 0.012832f
C539 VTAIL.n227 B 0.013587f
C540 VTAIL.n228 B 0.030331f
C541 VTAIL.n229 B 0.030331f
C542 VTAIL.n230 B 0.013587f
C543 VTAIL.n231 B 0.012832f
C544 VTAIL.n232 B 0.02388f
C545 VTAIL.n233 B 0.02388f
C546 VTAIL.n234 B 0.012832f
C547 VTAIL.n235 B 0.013587f
C548 VTAIL.n236 B 0.030331f
C549 VTAIL.n237 B 0.030331f
C550 VTAIL.n238 B 0.013587f
C551 VTAIL.n239 B 0.012832f
C552 VTAIL.n240 B 0.02388f
C553 VTAIL.n241 B 0.02388f
C554 VTAIL.n242 B 0.012832f
C555 VTAIL.n243 B 0.013587f
C556 VTAIL.n244 B 0.030331f
C557 VTAIL.n245 B 0.030331f
C558 VTAIL.n246 B 0.013587f
C559 VTAIL.n247 B 0.012832f
C560 VTAIL.n248 B 0.02388f
C561 VTAIL.n249 B 0.02388f
C562 VTAIL.n250 B 0.012832f
C563 VTAIL.n251 B 0.013587f
C564 VTAIL.n252 B 0.030331f
C565 VTAIL.n253 B 0.030331f
C566 VTAIL.n254 B 0.013587f
C567 VTAIL.n255 B 0.012832f
C568 VTAIL.n256 B 0.02388f
C569 VTAIL.n257 B 0.02388f
C570 VTAIL.n258 B 0.012832f
C571 VTAIL.n259 B 0.013587f
C572 VTAIL.n260 B 0.030331f
C573 VTAIL.n261 B 0.030331f
C574 VTAIL.n262 B 0.013587f
C575 VTAIL.n263 B 0.012832f
C576 VTAIL.n264 B 0.02388f
C577 VTAIL.n265 B 0.02388f
C578 VTAIL.n266 B 0.012832f
C579 VTAIL.n267 B 0.013587f
C580 VTAIL.n268 B 0.030331f
C581 VTAIL.n269 B 0.030331f
C582 VTAIL.n270 B 0.030331f
C583 VTAIL.n271 B 0.01321f
C584 VTAIL.n272 B 0.012832f
C585 VTAIL.n273 B 0.02388f
C586 VTAIL.n274 B 0.02388f
C587 VTAIL.n275 B 0.012832f
C588 VTAIL.n276 B 0.013587f
C589 VTAIL.n277 B 0.030331f
C590 VTAIL.n278 B 0.063096f
C591 VTAIL.n279 B 0.013587f
C592 VTAIL.n280 B 0.012832f
C593 VTAIL.n281 B 0.056177f
C594 VTAIL.n282 B 0.035071f
C595 VTAIL.n283 B 1.76819f
C596 VTAIL.n284 B 0.032116f
C597 VTAIL.n285 B 0.02388f
C598 VTAIL.n286 B 0.012832f
C599 VTAIL.n287 B 0.030331f
C600 VTAIL.n288 B 0.013587f
C601 VTAIL.n289 B 0.02388f
C602 VTAIL.n290 B 0.01321f
C603 VTAIL.n291 B 0.030331f
C604 VTAIL.n292 B 0.013587f
C605 VTAIL.n293 B 0.02388f
C606 VTAIL.n294 B 0.012832f
C607 VTAIL.n295 B 0.030331f
C608 VTAIL.n296 B 0.013587f
C609 VTAIL.n297 B 0.02388f
C610 VTAIL.n298 B 0.012832f
C611 VTAIL.n299 B 0.030331f
C612 VTAIL.n300 B 0.013587f
C613 VTAIL.n301 B 0.02388f
C614 VTAIL.n302 B 0.012832f
C615 VTAIL.n303 B 0.030331f
C616 VTAIL.n304 B 0.013587f
C617 VTAIL.n305 B 0.02388f
C618 VTAIL.n306 B 0.012832f
C619 VTAIL.n307 B 0.030331f
C620 VTAIL.n308 B 0.013587f
C621 VTAIL.n309 B 0.02388f
C622 VTAIL.n310 B 0.012832f
C623 VTAIL.n311 B 0.022748f
C624 VTAIL.n312 B 0.017917f
C625 VTAIL.t8 B 0.050102f
C626 VTAIL.n313 B 0.162398f
C627 VTAIL.n314 B 1.67516f
C628 VTAIL.n315 B 0.012832f
C629 VTAIL.n316 B 0.013587f
C630 VTAIL.n317 B 0.030331f
C631 VTAIL.n318 B 0.030331f
C632 VTAIL.n319 B 0.013587f
C633 VTAIL.n320 B 0.012832f
C634 VTAIL.n321 B 0.02388f
C635 VTAIL.n322 B 0.02388f
C636 VTAIL.n323 B 0.012832f
C637 VTAIL.n324 B 0.013587f
C638 VTAIL.n325 B 0.030331f
C639 VTAIL.n326 B 0.030331f
C640 VTAIL.n327 B 0.013587f
C641 VTAIL.n328 B 0.012832f
C642 VTAIL.n329 B 0.02388f
C643 VTAIL.n330 B 0.02388f
C644 VTAIL.n331 B 0.012832f
C645 VTAIL.n332 B 0.013587f
C646 VTAIL.n333 B 0.030331f
C647 VTAIL.n334 B 0.030331f
C648 VTAIL.n335 B 0.013587f
C649 VTAIL.n336 B 0.012832f
C650 VTAIL.n337 B 0.02388f
C651 VTAIL.n338 B 0.02388f
C652 VTAIL.n339 B 0.012832f
C653 VTAIL.n340 B 0.013587f
C654 VTAIL.n341 B 0.030331f
C655 VTAIL.n342 B 0.030331f
C656 VTAIL.n343 B 0.013587f
C657 VTAIL.n344 B 0.012832f
C658 VTAIL.n345 B 0.02388f
C659 VTAIL.n346 B 0.02388f
C660 VTAIL.n347 B 0.012832f
C661 VTAIL.n348 B 0.013587f
C662 VTAIL.n349 B 0.030331f
C663 VTAIL.n350 B 0.030331f
C664 VTAIL.n351 B 0.013587f
C665 VTAIL.n352 B 0.012832f
C666 VTAIL.n353 B 0.02388f
C667 VTAIL.n354 B 0.02388f
C668 VTAIL.n355 B 0.012832f
C669 VTAIL.n356 B 0.012832f
C670 VTAIL.n357 B 0.013587f
C671 VTAIL.n358 B 0.030331f
C672 VTAIL.n359 B 0.030331f
C673 VTAIL.n360 B 0.030331f
C674 VTAIL.n361 B 0.01321f
C675 VTAIL.n362 B 0.012832f
C676 VTAIL.n363 B 0.02388f
C677 VTAIL.n364 B 0.02388f
C678 VTAIL.n365 B 0.012832f
C679 VTAIL.n366 B 0.013587f
C680 VTAIL.n367 B 0.030331f
C681 VTAIL.n368 B 0.063096f
C682 VTAIL.n369 B 0.013587f
C683 VTAIL.n370 B 0.012832f
C684 VTAIL.n371 B 0.056177f
C685 VTAIL.n372 B 0.035071f
C686 VTAIL.n373 B 1.76819f
C687 VTAIL.t7 B 0.304009f
C688 VTAIL.t5 B 0.304009f
C689 VTAIL.n374 B 2.68581f
C690 VTAIL.n375 B 0.452106f
C691 VDD1.n0 B 0.032051f
C692 VDD1.n1 B 0.023832f
C693 VDD1.n2 B 0.012806f
C694 VDD1.n3 B 0.03027f
C695 VDD1.n4 B 0.01356f
C696 VDD1.n5 B 0.023832f
C697 VDD1.n6 B 0.013183f
C698 VDD1.n7 B 0.03027f
C699 VDD1.n8 B 0.012806f
C700 VDD1.n9 B 0.01356f
C701 VDD1.n10 B 0.023832f
C702 VDD1.n11 B 0.012806f
C703 VDD1.n12 B 0.03027f
C704 VDD1.n13 B 0.01356f
C705 VDD1.n14 B 0.023832f
C706 VDD1.n15 B 0.012806f
C707 VDD1.n16 B 0.03027f
C708 VDD1.n17 B 0.01356f
C709 VDD1.n18 B 0.023832f
C710 VDD1.n19 B 0.012806f
C711 VDD1.n20 B 0.03027f
C712 VDD1.n21 B 0.01356f
C713 VDD1.n22 B 0.023832f
C714 VDD1.n23 B 0.012806f
C715 VDD1.n24 B 0.03027f
C716 VDD1.n25 B 0.01356f
C717 VDD1.n26 B 0.023832f
C718 VDD1.n27 B 0.012806f
C719 VDD1.n28 B 0.022702f
C720 VDD1.n29 B 0.017881f
C721 VDD1.t4 B 0.050002f
C722 VDD1.n30 B 0.162072f
C723 VDD1.n31 B 1.6718f
C724 VDD1.n32 B 0.012806f
C725 VDD1.n33 B 0.01356f
C726 VDD1.n34 B 0.03027f
C727 VDD1.n35 B 0.03027f
C728 VDD1.n36 B 0.01356f
C729 VDD1.n37 B 0.012806f
C730 VDD1.n38 B 0.023832f
C731 VDD1.n39 B 0.023832f
C732 VDD1.n40 B 0.012806f
C733 VDD1.n41 B 0.01356f
C734 VDD1.n42 B 0.03027f
C735 VDD1.n43 B 0.03027f
C736 VDD1.n44 B 0.01356f
C737 VDD1.n45 B 0.012806f
C738 VDD1.n46 B 0.023832f
C739 VDD1.n47 B 0.023832f
C740 VDD1.n48 B 0.012806f
C741 VDD1.n49 B 0.01356f
C742 VDD1.n50 B 0.03027f
C743 VDD1.n51 B 0.03027f
C744 VDD1.n52 B 0.01356f
C745 VDD1.n53 B 0.012806f
C746 VDD1.n54 B 0.023832f
C747 VDD1.n55 B 0.023832f
C748 VDD1.n56 B 0.012806f
C749 VDD1.n57 B 0.01356f
C750 VDD1.n58 B 0.03027f
C751 VDD1.n59 B 0.03027f
C752 VDD1.n60 B 0.01356f
C753 VDD1.n61 B 0.012806f
C754 VDD1.n62 B 0.023832f
C755 VDD1.n63 B 0.023832f
C756 VDD1.n64 B 0.012806f
C757 VDD1.n65 B 0.01356f
C758 VDD1.n66 B 0.03027f
C759 VDD1.n67 B 0.03027f
C760 VDD1.n68 B 0.01356f
C761 VDD1.n69 B 0.012806f
C762 VDD1.n70 B 0.023832f
C763 VDD1.n71 B 0.023832f
C764 VDD1.n72 B 0.012806f
C765 VDD1.n73 B 0.01356f
C766 VDD1.n74 B 0.03027f
C767 VDD1.n75 B 0.03027f
C768 VDD1.n76 B 0.03027f
C769 VDD1.n77 B 0.013183f
C770 VDD1.n78 B 0.012806f
C771 VDD1.n79 B 0.023832f
C772 VDD1.n80 B 0.023832f
C773 VDD1.n81 B 0.012806f
C774 VDD1.n82 B 0.01356f
C775 VDD1.n83 B 0.03027f
C776 VDD1.n84 B 0.06297f
C777 VDD1.n85 B 0.01356f
C778 VDD1.n86 B 0.012806f
C779 VDD1.n87 B 0.056064f
C780 VDD1.n88 B 0.061377f
C781 VDD1.t1 B 0.3034f
C782 VDD1.t3 B 0.3034f
C783 VDD1.n89 B 2.7518f
C784 VDD1.n90 B 0.634424f
C785 VDD1.n91 B 0.032051f
C786 VDD1.n92 B 0.023832f
C787 VDD1.n93 B 0.012806f
C788 VDD1.n94 B 0.03027f
C789 VDD1.n95 B 0.01356f
C790 VDD1.n96 B 0.023832f
C791 VDD1.n97 B 0.013183f
C792 VDD1.n98 B 0.03027f
C793 VDD1.n99 B 0.01356f
C794 VDD1.n100 B 0.023832f
C795 VDD1.n101 B 0.012806f
C796 VDD1.n102 B 0.03027f
C797 VDD1.n103 B 0.01356f
C798 VDD1.n104 B 0.023832f
C799 VDD1.n105 B 0.012806f
C800 VDD1.n106 B 0.03027f
C801 VDD1.n107 B 0.01356f
C802 VDD1.n108 B 0.023832f
C803 VDD1.n109 B 0.012806f
C804 VDD1.n110 B 0.03027f
C805 VDD1.n111 B 0.01356f
C806 VDD1.n112 B 0.023832f
C807 VDD1.n113 B 0.012806f
C808 VDD1.n114 B 0.03027f
C809 VDD1.n115 B 0.01356f
C810 VDD1.n116 B 0.023832f
C811 VDD1.n117 B 0.012806f
C812 VDD1.n118 B 0.022702f
C813 VDD1.n119 B 0.017881f
C814 VDD1.t9 B 0.050002f
C815 VDD1.n120 B 0.162072f
C816 VDD1.n121 B 1.6718f
C817 VDD1.n122 B 0.012806f
C818 VDD1.n123 B 0.01356f
C819 VDD1.n124 B 0.03027f
C820 VDD1.n125 B 0.03027f
C821 VDD1.n126 B 0.01356f
C822 VDD1.n127 B 0.012806f
C823 VDD1.n128 B 0.023832f
C824 VDD1.n129 B 0.023832f
C825 VDD1.n130 B 0.012806f
C826 VDD1.n131 B 0.01356f
C827 VDD1.n132 B 0.03027f
C828 VDD1.n133 B 0.03027f
C829 VDD1.n134 B 0.01356f
C830 VDD1.n135 B 0.012806f
C831 VDD1.n136 B 0.023832f
C832 VDD1.n137 B 0.023832f
C833 VDD1.n138 B 0.012806f
C834 VDD1.n139 B 0.01356f
C835 VDD1.n140 B 0.03027f
C836 VDD1.n141 B 0.03027f
C837 VDD1.n142 B 0.01356f
C838 VDD1.n143 B 0.012806f
C839 VDD1.n144 B 0.023832f
C840 VDD1.n145 B 0.023832f
C841 VDD1.n146 B 0.012806f
C842 VDD1.n147 B 0.01356f
C843 VDD1.n148 B 0.03027f
C844 VDD1.n149 B 0.03027f
C845 VDD1.n150 B 0.01356f
C846 VDD1.n151 B 0.012806f
C847 VDD1.n152 B 0.023832f
C848 VDD1.n153 B 0.023832f
C849 VDD1.n154 B 0.012806f
C850 VDD1.n155 B 0.01356f
C851 VDD1.n156 B 0.03027f
C852 VDD1.n157 B 0.03027f
C853 VDD1.n158 B 0.01356f
C854 VDD1.n159 B 0.012806f
C855 VDD1.n160 B 0.023832f
C856 VDD1.n161 B 0.023832f
C857 VDD1.n162 B 0.012806f
C858 VDD1.n163 B 0.012806f
C859 VDD1.n164 B 0.01356f
C860 VDD1.n165 B 0.03027f
C861 VDD1.n166 B 0.03027f
C862 VDD1.n167 B 0.03027f
C863 VDD1.n168 B 0.013183f
C864 VDD1.n169 B 0.012806f
C865 VDD1.n170 B 0.023832f
C866 VDD1.n171 B 0.023832f
C867 VDD1.n172 B 0.012806f
C868 VDD1.n173 B 0.01356f
C869 VDD1.n174 B 0.03027f
C870 VDD1.n175 B 0.06297f
C871 VDD1.n176 B 0.01356f
C872 VDD1.n177 B 0.012806f
C873 VDD1.n178 B 0.056064f
C874 VDD1.n179 B 0.061377f
C875 VDD1.t7 B 0.3034f
C876 VDD1.t5 B 0.3034f
C877 VDD1.n180 B 2.7518f
C878 VDD1.n181 B 0.626776f
C879 VDD1.t0 B 0.3034f
C880 VDD1.t2 B 0.3034f
C881 VDD1.n182 B 2.76534f
C882 VDD1.n183 B 2.99843f
C883 VDD1.t8 B 0.3034f
C884 VDD1.t6 B 0.3034f
C885 VDD1.n184 B 2.7518f
C886 VDD1.n185 B 3.21955f
C887 VP.n0 B 0.029713f
C888 VP.t3 B 2.3317f
C889 VP.n1 B 0.018227f
C890 VP.n2 B 0.022537f
C891 VP.t9 B 2.3317f
C892 VP.n3 B 0.042004f
C893 VP.n4 B 0.022537f
C894 VP.t4 B 2.3317f
C895 VP.n5 B 0.835657f
C896 VP.n6 B 0.022537f
C897 VP.n7 B 0.042004f
C898 VP.n8 B 0.022537f
C899 VP.t0 B 2.3317f
C900 VP.n9 B 0.018227f
C901 VP.n10 B 0.029713f
C902 VP.t6 B 2.3317f
C903 VP.n11 B 0.029713f
C904 VP.t1 B 2.3317f
C905 VP.n12 B 0.018227f
C906 VP.n13 B 0.022537f
C907 VP.t7 B 2.3317f
C908 VP.n14 B 0.042004f
C909 VP.n15 B 0.022537f
C910 VP.t2 B 2.3317f
C911 VP.n16 B 0.835657f
C912 VP.n17 B 0.022537f
C913 VP.n18 B 0.042004f
C914 VP.t5 B 2.48839f
C915 VP.n19 B 0.862414f
C916 VP.t8 B 2.3317f
C917 VP.n20 B 0.871865f
C918 VP.n21 B 0.028317f
C919 VP.n22 B 0.194937f
C920 VP.n23 B 0.022537f
C921 VP.n24 B 0.022537f
C922 VP.n25 B 0.027564f
C923 VP.n26 B 0.03824f
C924 VP.n27 B 0.042004f
C925 VP.n28 B 0.022537f
C926 VP.n29 B 0.022537f
C927 VP.n30 B 0.022537f
C928 VP.n31 B 0.042004f
C929 VP.n32 B 0.03824f
C930 VP.n33 B 0.027564f
C931 VP.n34 B 0.022537f
C932 VP.n35 B 0.022537f
C933 VP.n36 B 0.022537f
C934 VP.n37 B 0.028317f
C935 VP.n38 B 0.814391f
C936 VP.n39 B 0.034953f
C937 VP.n40 B 0.044904f
C938 VP.n41 B 0.022537f
C939 VP.n42 B 0.022537f
C940 VP.n43 B 0.022537f
C941 VP.n44 B 0.044677f
C942 VP.n45 B 0.035368f
C943 VP.n46 B 0.890578f
C944 VP.n47 B 1.42799f
C945 VP.n48 B 1.44275f
C946 VP.n49 B 0.890578f
C947 VP.n50 B 0.035368f
C948 VP.n51 B 0.044677f
C949 VP.n52 B 0.022537f
C950 VP.n53 B 0.022537f
C951 VP.n54 B 0.022537f
C952 VP.n55 B 0.044904f
C953 VP.n56 B 0.034953f
C954 VP.n57 B 0.814391f
C955 VP.n58 B 0.028317f
C956 VP.n59 B 0.022537f
C957 VP.n60 B 0.022537f
C958 VP.n61 B 0.022537f
C959 VP.n62 B 0.027564f
C960 VP.n63 B 0.03824f
C961 VP.n64 B 0.042004f
C962 VP.n65 B 0.022537f
C963 VP.n66 B 0.022537f
C964 VP.n67 B 0.022537f
C965 VP.n68 B 0.042004f
C966 VP.n69 B 0.03824f
C967 VP.n70 B 0.027564f
C968 VP.n71 B 0.022537f
C969 VP.n72 B 0.022537f
C970 VP.n73 B 0.022537f
C971 VP.n74 B 0.028317f
C972 VP.n75 B 0.814391f
C973 VP.n76 B 0.034953f
C974 VP.n77 B 0.044904f
C975 VP.n78 B 0.022537f
C976 VP.n79 B 0.022537f
C977 VP.n80 B 0.022537f
C978 VP.n81 B 0.044677f
C979 VP.n82 B 0.035368f
C980 VP.n83 B 0.890578f
C981 VP.n84 B 0.030913f
.ends

