* NGSPICE file created from diff_pair_sample_1426.ext - technology: sky130A

.subckt diff_pair_sample_1426 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1534_n1608# sky130_fd_pr__pfet_01v8 ad=1.248 pd=7.18 as=0 ps=0 w=3.2 l=0.61
X1 VDD1.t3 VP.t0 VTAIL.t7 w_n1534_n1608# sky130_fd_pr__pfet_01v8 ad=0.528 pd=3.53 as=1.248 ps=7.18 w=3.2 l=0.61
X2 B.t8 B.t6 B.t7 w_n1534_n1608# sky130_fd_pr__pfet_01v8 ad=1.248 pd=7.18 as=0 ps=0 w=3.2 l=0.61
X3 B.t5 B.t3 B.t4 w_n1534_n1608# sky130_fd_pr__pfet_01v8 ad=1.248 pd=7.18 as=0 ps=0 w=3.2 l=0.61
X4 VTAIL.t6 VP.t1 VDD1.t2 w_n1534_n1608# sky130_fd_pr__pfet_01v8 ad=1.248 pd=7.18 as=0.528 ps=3.53 w=3.2 l=0.61
X5 VDD2.t3 VN.t0 VTAIL.t1 w_n1534_n1608# sky130_fd_pr__pfet_01v8 ad=0.528 pd=3.53 as=1.248 ps=7.18 w=3.2 l=0.61
X6 VDD2.t2 VN.t1 VTAIL.t2 w_n1534_n1608# sky130_fd_pr__pfet_01v8 ad=0.528 pd=3.53 as=1.248 ps=7.18 w=3.2 l=0.61
X7 B.t2 B.t0 B.t1 w_n1534_n1608# sky130_fd_pr__pfet_01v8 ad=1.248 pd=7.18 as=0 ps=0 w=3.2 l=0.61
X8 VDD1.t1 VP.t2 VTAIL.t4 w_n1534_n1608# sky130_fd_pr__pfet_01v8 ad=0.528 pd=3.53 as=1.248 ps=7.18 w=3.2 l=0.61
X9 VTAIL.t0 VN.t2 VDD2.t1 w_n1534_n1608# sky130_fd_pr__pfet_01v8 ad=1.248 pd=7.18 as=0.528 ps=3.53 w=3.2 l=0.61
X10 VTAIL.t3 VN.t3 VDD2.t0 w_n1534_n1608# sky130_fd_pr__pfet_01v8 ad=1.248 pd=7.18 as=0.528 ps=3.53 w=3.2 l=0.61
X11 VTAIL.t5 VP.t3 VDD1.t0 w_n1534_n1608# sky130_fd_pr__pfet_01v8 ad=1.248 pd=7.18 as=0.528 ps=3.53 w=3.2 l=0.61
R0 B.n169 B.n52 585
R1 B.n168 B.n167 585
R2 B.n166 B.n53 585
R3 B.n165 B.n164 585
R4 B.n163 B.n54 585
R5 B.n162 B.n161 585
R6 B.n160 B.n55 585
R7 B.n159 B.n158 585
R8 B.n157 B.n56 585
R9 B.n156 B.n155 585
R10 B.n154 B.n57 585
R11 B.n153 B.n152 585
R12 B.n151 B.n58 585
R13 B.n150 B.n149 585
R14 B.n148 B.n59 585
R15 B.n147 B.n146 585
R16 B.n145 B.n144 585
R17 B.n143 B.n63 585
R18 B.n142 B.n141 585
R19 B.n140 B.n64 585
R20 B.n139 B.n138 585
R21 B.n137 B.n65 585
R22 B.n136 B.n135 585
R23 B.n134 B.n66 585
R24 B.n133 B.n132 585
R25 B.n130 B.n67 585
R26 B.n129 B.n128 585
R27 B.n127 B.n70 585
R28 B.n126 B.n125 585
R29 B.n124 B.n71 585
R30 B.n123 B.n122 585
R31 B.n121 B.n72 585
R32 B.n120 B.n119 585
R33 B.n118 B.n73 585
R34 B.n117 B.n116 585
R35 B.n115 B.n74 585
R36 B.n114 B.n113 585
R37 B.n112 B.n75 585
R38 B.n111 B.n110 585
R39 B.n109 B.n76 585
R40 B.n108 B.n107 585
R41 B.n171 B.n170 585
R42 B.n172 B.n51 585
R43 B.n174 B.n173 585
R44 B.n175 B.n50 585
R45 B.n177 B.n176 585
R46 B.n178 B.n49 585
R47 B.n180 B.n179 585
R48 B.n181 B.n48 585
R49 B.n183 B.n182 585
R50 B.n184 B.n47 585
R51 B.n186 B.n185 585
R52 B.n187 B.n46 585
R53 B.n189 B.n188 585
R54 B.n190 B.n45 585
R55 B.n192 B.n191 585
R56 B.n193 B.n44 585
R57 B.n195 B.n194 585
R58 B.n196 B.n43 585
R59 B.n198 B.n197 585
R60 B.n199 B.n42 585
R61 B.n201 B.n200 585
R62 B.n202 B.n41 585
R63 B.n204 B.n203 585
R64 B.n205 B.n40 585
R65 B.n207 B.n206 585
R66 B.n208 B.n39 585
R67 B.n210 B.n209 585
R68 B.n211 B.n38 585
R69 B.n213 B.n212 585
R70 B.n214 B.n37 585
R71 B.n216 B.n215 585
R72 B.n217 B.n36 585
R73 B.n219 B.n218 585
R74 B.n220 B.n35 585
R75 B.n283 B.n10 585
R76 B.n282 B.n281 585
R77 B.n280 B.n11 585
R78 B.n279 B.n278 585
R79 B.n277 B.n12 585
R80 B.n276 B.n275 585
R81 B.n274 B.n13 585
R82 B.n273 B.n272 585
R83 B.n271 B.n14 585
R84 B.n270 B.n269 585
R85 B.n268 B.n15 585
R86 B.n267 B.n266 585
R87 B.n265 B.n16 585
R88 B.n264 B.n263 585
R89 B.n262 B.n17 585
R90 B.n261 B.n260 585
R91 B.n259 B.n258 585
R92 B.n257 B.n21 585
R93 B.n256 B.n255 585
R94 B.n254 B.n22 585
R95 B.n253 B.n252 585
R96 B.n251 B.n23 585
R97 B.n250 B.n249 585
R98 B.n248 B.n24 585
R99 B.n247 B.n246 585
R100 B.n244 B.n25 585
R101 B.n243 B.n242 585
R102 B.n241 B.n28 585
R103 B.n240 B.n239 585
R104 B.n238 B.n29 585
R105 B.n237 B.n236 585
R106 B.n235 B.n30 585
R107 B.n234 B.n233 585
R108 B.n232 B.n31 585
R109 B.n231 B.n230 585
R110 B.n229 B.n32 585
R111 B.n228 B.n227 585
R112 B.n226 B.n33 585
R113 B.n225 B.n224 585
R114 B.n223 B.n34 585
R115 B.n222 B.n221 585
R116 B.n285 B.n284 585
R117 B.n286 B.n9 585
R118 B.n288 B.n287 585
R119 B.n289 B.n8 585
R120 B.n291 B.n290 585
R121 B.n292 B.n7 585
R122 B.n294 B.n293 585
R123 B.n295 B.n6 585
R124 B.n297 B.n296 585
R125 B.n298 B.n5 585
R126 B.n300 B.n299 585
R127 B.n301 B.n4 585
R128 B.n303 B.n302 585
R129 B.n304 B.n3 585
R130 B.n306 B.n305 585
R131 B.n307 B.n0 585
R132 B.n2 B.n1 585
R133 B.n85 B.n84 585
R134 B.n87 B.n86 585
R135 B.n88 B.n83 585
R136 B.n90 B.n89 585
R137 B.n91 B.n82 585
R138 B.n93 B.n92 585
R139 B.n94 B.n81 585
R140 B.n96 B.n95 585
R141 B.n97 B.n80 585
R142 B.n99 B.n98 585
R143 B.n100 B.n79 585
R144 B.n102 B.n101 585
R145 B.n103 B.n78 585
R146 B.n105 B.n104 585
R147 B.n106 B.n77 585
R148 B.n108 B.n77 487.695
R149 B.n170 B.n169 487.695
R150 B.n222 B.n35 487.695
R151 B.n284 B.n283 487.695
R152 B.n68 B.t9 330.661
R153 B.n60 B.t3 330.661
R154 B.n26 B.t6 330.661
R155 B.n18 B.t0 330.661
R156 B.n309 B.n308 256.663
R157 B.n60 B.t4 243.792
R158 B.n26 B.t8 243.792
R159 B.n68 B.t10 243.791
R160 B.n18 B.t2 243.791
R161 B.n308 B.n307 235.042
R162 B.n308 B.n2 235.042
R163 B.n61 B.t5 225.56
R164 B.n27 B.t7 225.56
R165 B.n69 B.t11 225.56
R166 B.n19 B.t1 225.56
R167 B.n109 B.n108 163.367
R168 B.n110 B.n109 163.367
R169 B.n110 B.n75 163.367
R170 B.n114 B.n75 163.367
R171 B.n115 B.n114 163.367
R172 B.n116 B.n115 163.367
R173 B.n116 B.n73 163.367
R174 B.n120 B.n73 163.367
R175 B.n121 B.n120 163.367
R176 B.n122 B.n121 163.367
R177 B.n122 B.n71 163.367
R178 B.n126 B.n71 163.367
R179 B.n127 B.n126 163.367
R180 B.n128 B.n127 163.367
R181 B.n128 B.n67 163.367
R182 B.n133 B.n67 163.367
R183 B.n134 B.n133 163.367
R184 B.n135 B.n134 163.367
R185 B.n135 B.n65 163.367
R186 B.n139 B.n65 163.367
R187 B.n140 B.n139 163.367
R188 B.n141 B.n140 163.367
R189 B.n141 B.n63 163.367
R190 B.n145 B.n63 163.367
R191 B.n146 B.n145 163.367
R192 B.n146 B.n59 163.367
R193 B.n150 B.n59 163.367
R194 B.n151 B.n150 163.367
R195 B.n152 B.n151 163.367
R196 B.n152 B.n57 163.367
R197 B.n156 B.n57 163.367
R198 B.n157 B.n156 163.367
R199 B.n158 B.n157 163.367
R200 B.n158 B.n55 163.367
R201 B.n162 B.n55 163.367
R202 B.n163 B.n162 163.367
R203 B.n164 B.n163 163.367
R204 B.n164 B.n53 163.367
R205 B.n168 B.n53 163.367
R206 B.n169 B.n168 163.367
R207 B.n218 B.n35 163.367
R208 B.n218 B.n217 163.367
R209 B.n217 B.n216 163.367
R210 B.n216 B.n37 163.367
R211 B.n212 B.n37 163.367
R212 B.n212 B.n211 163.367
R213 B.n211 B.n210 163.367
R214 B.n210 B.n39 163.367
R215 B.n206 B.n39 163.367
R216 B.n206 B.n205 163.367
R217 B.n205 B.n204 163.367
R218 B.n204 B.n41 163.367
R219 B.n200 B.n41 163.367
R220 B.n200 B.n199 163.367
R221 B.n199 B.n198 163.367
R222 B.n198 B.n43 163.367
R223 B.n194 B.n43 163.367
R224 B.n194 B.n193 163.367
R225 B.n193 B.n192 163.367
R226 B.n192 B.n45 163.367
R227 B.n188 B.n45 163.367
R228 B.n188 B.n187 163.367
R229 B.n187 B.n186 163.367
R230 B.n186 B.n47 163.367
R231 B.n182 B.n47 163.367
R232 B.n182 B.n181 163.367
R233 B.n181 B.n180 163.367
R234 B.n180 B.n49 163.367
R235 B.n176 B.n49 163.367
R236 B.n176 B.n175 163.367
R237 B.n175 B.n174 163.367
R238 B.n174 B.n51 163.367
R239 B.n170 B.n51 163.367
R240 B.n283 B.n282 163.367
R241 B.n282 B.n11 163.367
R242 B.n278 B.n11 163.367
R243 B.n278 B.n277 163.367
R244 B.n277 B.n276 163.367
R245 B.n276 B.n13 163.367
R246 B.n272 B.n13 163.367
R247 B.n272 B.n271 163.367
R248 B.n271 B.n270 163.367
R249 B.n270 B.n15 163.367
R250 B.n266 B.n15 163.367
R251 B.n266 B.n265 163.367
R252 B.n265 B.n264 163.367
R253 B.n264 B.n17 163.367
R254 B.n260 B.n17 163.367
R255 B.n260 B.n259 163.367
R256 B.n259 B.n21 163.367
R257 B.n255 B.n21 163.367
R258 B.n255 B.n254 163.367
R259 B.n254 B.n253 163.367
R260 B.n253 B.n23 163.367
R261 B.n249 B.n23 163.367
R262 B.n249 B.n248 163.367
R263 B.n248 B.n247 163.367
R264 B.n247 B.n25 163.367
R265 B.n242 B.n25 163.367
R266 B.n242 B.n241 163.367
R267 B.n241 B.n240 163.367
R268 B.n240 B.n29 163.367
R269 B.n236 B.n29 163.367
R270 B.n236 B.n235 163.367
R271 B.n235 B.n234 163.367
R272 B.n234 B.n31 163.367
R273 B.n230 B.n31 163.367
R274 B.n230 B.n229 163.367
R275 B.n229 B.n228 163.367
R276 B.n228 B.n33 163.367
R277 B.n224 B.n33 163.367
R278 B.n224 B.n223 163.367
R279 B.n223 B.n222 163.367
R280 B.n284 B.n9 163.367
R281 B.n288 B.n9 163.367
R282 B.n289 B.n288 163.367
R283 B.n290 B.n289 163.367
R284 B.n290 B.n7 163.367
R285 B.n294 B.n7 163.367
R286 B.n295 B.n294 163.367
R287 B.n296 B.n295 163.367
R288 B.n296 B.n5 163.367
R289 B.n300 B.n5 163.367
R290 B.n301 B.n300 163.367
R291 B.n302 B.n301 163.367
R292 B.n302 B.n3 163.367
R293 B.n306 B.n3 163.367
R294 B.n307 B.n306 163.367
R295 B.n85 B.n2 163.367
R296 B.n86 B.n85 163.367
R297 B.n86 B.n83 163.367
R298 B.n90 B.n83 163.367
R299 B.n91 B.n90 163.367
R300 B.n92 B.n91 163.367
R301 B.n92 B.n81 163.367
R302 B.n96 B.n81 163.367
R303 B.n97 B.n96 163.367
R304 B.n98 B.n97 163.367
R305 B.n98 B.n79 163.367
R306 B.n102 B.n79 163.367
R307 B.n103 B.n102 163.367
R308 B.n104 B.n103 163.367
R309 B.n104 B.n77 163.367
R310 B.n131 B.n69 59.5399
R311 B.n62 B.n61 59.5399
R312 B.n245 B.n27 59.5399
R313 B.n20 B.n19 59.5399
R314 B.n285 B.n10 31.6883
R315 B.n221 B.n220 31.6883
R316 B.n171 B.n52 31.6883
R317 B.n107 B.n106 31.6883
R318 B.n69 B.n68 18.2308
R319 B.n61 B.n60 18.2308
R320 B.n27 B.n26 18.2308
R321 B.n19 B.n18 18.2308
R322 B B.n309 18.0485
R323 B.n286 B.n285 10.6151
R324 B.n287 B.n286 10.6151
R325 B.n287 B.n8 10.6151
R326 B.n291 B.n8 10.6151
R327 B.n292 B.n291 10.6151
R328 B.n293 B.n292 10.6151
R329 B.n293 B.n6 10.6151
R330 B.n297 B.n6 10.6151
R331 B.n298 B.n297 10.6151
R332 B.n299 B.n298 10.6151
R333 B.n299 B.n4 10.6151
R334 B.n303 B.n4 10.6151
R335 B.n304 B.n303 10.6151
R336 B.n305 B.n304 10.6151
R337 B.n305 B.n0 10.6151
R338 B.n281 B.n10 10.6151
R339 B.n281 B.n280 10.6151
R340 B.n280 B.n279 10.6151
R341 B.n279 B.n12 10.6151
R342 B.n275 B.n12 10.6151
R343 B.n275 B.n274 10.6151
R344 B.n274 B.n273 10.6151
R345 B.n273 B.n14 10.6151
R346 B.n269 B.n14 10.6151
R347 B.n269 B.n268 10.6151
R348 B.n268 B.n267 10.6151
R349 B.n267 B.n16 10.6151
R350 B.n263 B.n16 10.6151
R351 B.n263 B.n262 10.6151
R352 B.n262 B.n261 10.6151
R353 B.n258 B.n257 10.6151
R354 B.n257 B.n256 10.6151
R355 B.n256 B.n22 10.6151
R356 B.n252 B.n22 10.6151
R357 B.n252 B.n251 10.6151
R358 B.n251 B.n250 10.6151
R359 B.n250 B.n24 10.6151
R360 B.n246 B.n24 10.6151
R361 B.n244 B.n243 10.6151
R362 B.n243 B.n28 10.6151
R363 B.n239 B.n28 10.6151
R364 B.n239 B.n238 10.6151
R365 B.n238 B.n237 10.6151
R366 B.n237 B.n30 10.6151
R367 B.n233 B.n30 10.6151
R368 B.n233 B.n232 10.6151
R369 B.n232 B.n231 10.6151
R370 B.n231 B.n32 10.6151
R371 B.n227 B.n32 10.6151
R372 B.n227 B.n226 10.6151
R373 B.n226 B.n225 10.6151
R374 B.n225 B.n34 10.6151
R375 B.n221 B.n34 10.6151
R376 B.n220 B.n219 10.6151
R377 B.n219 B.n36 10.6151
R378 B.n215 B.n36 10.6151
R379 B.n215 B.n214 10.6151
R380 B.n214 B.n213 10.6151
R381 B.n213 B.n38 10.6151
R382 B.n209 B.n38 10.6151
R383 B.n209 B.n208 10.6151
R384 B.n208 B.n207 10.6151
R385 B.n207 B.n40 10.6151
R386 B.n203 B.n40 10.6151
R387 B.n203 B.n202 10.6151
R388 B.n202 B.n201 10.6151
R389 B.n201 B.n42 10.6151
R390 B.n197 B.n42 10.6151
R391 B.n197 B.n196 10.6151
R392 B.n196 B.n195 10.6151
R393 B.n195 B.n44 10.6151
R394 B.n191 B.n44 10.6151
R395 B.n191 B.n190 10.6151
R396 B.n190 B.n189 10.6151
R397 B.n189 B.n46 10.6151
R398 B.n185 B.n46 10.6151
R399 B.n185 B.n184 10.6151
R400 B.n184 B.n183 10.6151
R401 B.n183 B.n48 10.6151
R402 B.n179 B.n48 10.6151
R403 B.n179 B.n178 10.6151
R404 B.n178 B.n177 10.6151
R405 B.n177 B.n50 10.6151
R406 B.n173 B.n50 10.6151
R407 B.n173 B.n172 10.6151
R408 B.n172 B.n171 10.6151
R409 B.n84 B.n1 10.6151
R410 B.n87 B.n84 10.6151
R411 B.n88 B.n87 10.6151
R412 B.n89 B.n88 10.6151
R413 B.n89 B.n82 10.6151
R414 B.n93 B.n82 10.6151
R415 B.n94 B.n93 10.6151
R416 B.n95 B.n94 10.6151
R417 B.n95 B.n80 10.6151
R418 B.n99 B.n80 10.6151
R419 B.n100 B.n99 10.6151
R420 B.n101 B.n100 10.6151
R421 B.n101 B.n78 10.6151
R422 B.n105 B.n78 10.6151
R423 B.n106 B.n105 10.6151
R424 B.n107 B.n76 10.6151
R425 B.n111 B.n76 10.6151
R426 B.n112 B.n111 10.6151
R427 B.n113 B.n112 10.6151
R428 B.n113 B.n74 10.6151
R429 B.n117 B.n74 10.6151
R430 B.n118 B.n117 10.6151
R431 B.n119 B.n118 10.6151
R432 B.n119 B.n72 10.6151
R433 B.n123 B.n72 10.6151
R434 B.n124 B.n123 10.6151
R435 B.n125 B.n124 10.6151
R436 B.n125 B.n70 10.6151
R437 B.n129 B.n70 10.6151
R438 B.n130 B.n129 10.6151
R439 B.n132 B.n66 10.6151
R440 B.n136 B.n66 10.6151
R441 B.n137 B.n136 10.6151
R442 B.n138 B.n137 10.6151
R443 B.n138 B.n64 10.6151
R444 B.n142 B.n64 10.6151
R445 B.n143 B.n142 10.6151
R446 B.n144 B.n143 10.6151
R447 B.n148 B.n147 10.6151
R448 B.n149 B.n148 10.6151
R449 B.n149 B.n58 10.6151
R450 B.n153 B.n58 10.6151
R451 B.n154 B.n153 10.6151
R452 B.n155 B.n154 10.6151
R453 B.n155 B.n56 10.6151
R454 B.n159 B.n56 10.6151
R455 B.n160 B.n159 10.6151
R456 B.n161 B.n160 10.6151
R457 B.n161 B.n54 10.6151
R458 B.n165 B.n54 10.6151
R459 B.n166 B.n165 10.6151
R460 B.n167 B.n166 10.6151
R461 B.n167 B.n52 10.6151
R462 B.n309 B.n0 8.11757
R463 B.n309 B.n1 8.11757
R464 B.n258 B.n20 6.5566
R465 B.n246 B.n245 6.5566
R466 B.n132 B.n131 6.5566
R467 B.n144 B.n62 6.5566
R468 B.n261 B.n20 4.05904
R469 B.n245 B.n244 4.05904
R470 B.n131 B.n130 4.05904
R471 B.n147 B.n62 4.05904
R472 VP.n0 VP.t3 211.806
R473 VP.n0 VP.t0 211.782
R474 VP.n2 VP.t1 190.826
R475 VP.n3 VP.t2 190.826
R476 VP.n4 VP.n3 161.3
R477 VP.n2 VP.n1 161.3
R478 VP.n1 VP.n0 103.805
R479 VP.n3 VP.n2 48.2005
R480 VP.n4 VP.n1 0.189894
R481 VP VP.n4 0.0516364
R482 VTAIL.n122 VTAIL.n112 756.745
R483 VTAIL.n10 VTAIL.n0 756.745
R484 VTAIL.n26 VTAIL.n16 756.745
R485 VTAIL.n42 VTAIL.n32 756.745
R486 VTAIL.n106 VTAIL.n96 756.745
R487 VTAIL.n90 VTAIL.n80 756.745
R488 VTAIL.n74 VTAIL.n64 756.745
R489 VTAIL.n58 VTAIL.n48 756.745
R490 VTAIL.n116 VTAIL.n115 585
R491 VTAIL.n121 VTAIL.n120 585
R492 VTAIL.n123 VTAIL.n122 585
R493 VTAIL.n4 VTAIL.n3 585
R494 VTAIL.n9 VTAIL.n8 585
R495 VTAIL.n11 VTAIL.n10 585
R496 VTAIL.n20 VTAIL.n19 585
R497 VTAIL.n25 VTAIL.n24 585
R498 VTAIL.n27 VTAIL.n26 585
R499 VTAIL.n36 VTAIL.n35 585
R500 VTAIL.n41 VTAIL.n40 585
R501 VTAIL.n43 VTAIL.n42 585
R502 VTAIL.n107 VTAIL.n106 585
R503 VTAIL.n105 VTAIL.n104 585
R504 VTAIL.n100 VTAIL.n99 585
R505 VTAIL.n91 VTAIL.n90 585
R506 VTAIL.n89 VTAIL.n88 585
R507 VTAIL.n84 VTAIL.n83 585
R508 VTAIL.n75 VTAIL.n74 585
R509 VTAIL.n73 VTAIL.n72 585
R510 VTAIL.n68 VTAIL.n67 585
R511 VTAIL.n59 VTAIL.n58 585
R512 VTAIL.n57 VTAIL.n56 585
R513 VTAIL.n52 VTAIL.n51 585
R514 VTAIL.n117 VTAIL.t2 336.901
R515 VTAIL.n5 VTAIL.t3 336.901
R516 VTAIL.n21 VTAIL.t4 336.901
R517 VTAIL.n37 VTAIL.t6 336.901
R518 VTAIL.n101 VTAIL.t7 336.901
R519 VTAIL.n85 VTAIL.t5 336.901
R520 VTAIL.n69 VTAIL.t1 336.901
R521 VTAIL.n53 VTAIL.t0 336.901
R522 VTAIL.n121 VTAIL.n115 171.744
R523 VTAIL.n122 VTAIL.n121 171.744
R524 VTAIL.n9 VTAIL.n3 171.744
R525 VTAIL.n10 VTAIL.n9 171.744
R526 VTAIL.n25 VTAIL.n19 171.744
R527 VTAIL.n26 VTAIL.n25 171.744
R528 VTAIL.n41 VTAIL.n35 171.744
R529 VTAIL.n42 VTAIL.n41 171.744
R530 VTAIL.n106 VTAIL.n105 171.744
R531 VTAIL.n105 VTAIL.n99 171.744
R532 VTAIL.n90 VTAIL.n89 171.744
R533 VTAIL.n89 VTAIL.n83 171.744
R534 VTAIL.n74 VTAIL.n73 171.744
R535 VTAIL.n73 VTAIL.n67 171.744
R536 VTAIL.n58 VTAIL.n57 171.744
R537 VTAIL.n57 VTAIL.n51 171.744
R538 VTAIL.t2 VTAIL.n115 85.8723
R539 VTAIL.t3 VTAIL.n3 85.8723
R540 VTAIL.t4 VTAIL.n19 85.8723
R541 VTAIL.t6 VTAIL.n35 85.8723
R542 VTAIL.t7 VTAIL.n99 85.8723
R543 VTAIL.t5 VTAIL.n83 85.8723
R544 VTAIL.t1 VTAIL.n67 85.8723
R545 VTAIL.t0 VTAIL.n51 85.8723
R546 VTAIL.n127 VTAIL.n126 33.7369
R547 VTAIL.n15 VTAIL.n14 33.7369
R548 VTAIL.n31 VTAIL.n30 33.7369
R549 VTAIL.n47 VTAIL.n46 33.7369
R550 VTAIL.n111 VTAIL.n110 33.7369
R551 VTAIL.n95 VTAIL.n94 33.7369
R552 VTAIL.n79 VTAIL.n78 33.7369
R553 VTAIL.n63 VTAIL.n62 33.7369
R554 VTAIL.n117 VTAIL.n116 16.193
R555 VTAIL.n5 VTAIL.n4 16.193
R556 VTAIL.n21 VTAIL.n20 16.193
R557 VTAIL.n37 VTAIL.n36 16.193
R558 VTAIL.n101 VTAIL.n100 16.193
R559 VTAIL.n85 VTAIL.n84 16.193
R560 VTAIL.n69 VTAIL.n68 16.193
R561 VTAIL.n53 VTAIL.n52 16.193
R562 VTAIL.n127 VTAIL.n111 15.9358
R563 VTAIL.n63 VTAIL.n47 15.9358
R564 VTAIL.n120 VTAIL.n119 12.8005
R565 VTAIL.n8 VTAIL.n7 12.8005
R566 VTAIL.n24 VTAIL.n23 12.8005
R567 VTAIL.n40 VTAIL.n39 12.8005
R568 VTAIL.n104 VTAIL.n103 12.8005
R569 VTAIL.n88 VTAIL.n87 12.8005
R570 VTAIL.n72 VTAIL.n71 12.8005
R571 VTAIL.n56 VTAIL.n55 12.8005
R572 VTAIL.n123 VTAIL.n114 12.0247
R573 VTAIL.n11 VTAIL.n2 12.0247
R574 VTAIL.n27 VTAIL.n18 12.0247
R575 VTAIL.n43 VTAIL.n34 12.0247
R576 VTAIL.n107 VTAIL.n98 12.0247
R577 VTAIL.n91 VTAIL.n82 12.0247
R578 VTAIL.n75 VTAIL.n66 12.0247
R579 VTAIL.n59 VTAIL.n50 12.0247
R580 VTAIL.n124 VTAIL.n112 11.249
R581 VTAIL.n12 VTAIL.n0 11.249
R582 VTAIL.n28 VTAIL.n16 11.249
R583 VTAIL.n44 VTAIL.n32 11.249
R584 VTAIL.n108 VTAIL.n96 11.249
R585 VTAIL.n92 VTAIL.n80 11.249
R586 VTAIL.n76 VTAIL.n64 11.249
R587 VTAIL.n60 VTAIL.n48 11.249
R588 VTAIL.n126 VTAIL.n125 9.45567
R589 VTAIL.n14 VTAIL.n13 9.45567
R590 VTAIL.n30 VTAIL.n29 9.45567
R591 VTAIL.n46 VTAIL.n45 9.45567
R592 VTAIL.n110 VTAIL.n109 9.45567
R593 VTAIL.n94 VTAIL.n93 9.45567
R594 VTAIL.n78 VTAIL.n77 9.45567
R595 VTAIL.n62 VTAIL.n61 9.45567
R596 VTAIL.n125 VTAIL.n124 9.3005
R597 VTAIL.n114 VTAIL.n113 9.3005
R598 VTAIL.n119 VTAIL.n118 9.3005
R599 VTAIL.n13 VTAIL.n12 9.3005
R600 VTAIL.n2 VTAIL.n1 9.3005
R601 VTAIL.n7 VTAIL.n6 9.3005
R602 VTAIL.n29 VTAIL.n28 9.3005
R603 VTAIL.n18 VTAIL.n17 9.3005
R604 VTAIL.n23 VTAIL.n22 9.3005
R605 VTAIL.n45 VTAIL.n44 9.3005
R606 VTAIL.n34 VTAIL.n33 9.3005
R607 VTAIL.n39 VTAIL.n38 9.3005
R608 VTAIL.n109 VTAIL.n108 9.3005
R609 VTAIL.n98 VTAIL.n97 9.3005
R610 VTAIL.n103 VTAIL.n102 9.3005
R611 VTAIL.n93 VTAIL.n92 9.3005
R612 VTAIL.n82 VTAIL.n81 9.3005
R613 VTAIL.n87 VTAIL.n86 9.3005
R614 VTAIL.n77 VTAIL.n76 9.3005
R615 VTAIL.n66 VTAIL.n65 9.3005
R616 VTAIL.n71 VTAIL.n70 9.3005
R617 VTAIL.n61 VTAIL.n60 9.3005
R618 VTAIL.n50 VTAIL.n49 9.3005
R619 VTAIL.n55 VTAIL.n54 9.3005
R620 VTAIL.n102 VTAIL.n101 3.91276
R621 VTAIL.n86 VTAIL.n85 3.91276
R622 VTAIL.n70 VTAIL.n69 3.91276
R623 VTAIL.n54 VTAIL.n53 3.91276
R624 VTAIL.n118 VTAIL.n117 3.91276
R625 VTAIL.n6 VTAIL.n5 3.91276
R626 VTAIL.n22 VTAIL.n21 3.91276
R627 VTAIL.n38 VTAIL.n37 3.91276
R628 VTAIL.n126 VTAIL.n112 2.71565
R629 VTAIL.n14 VTAIL.n0 2.71565
R630 VTAIL.n30 VTAIL.n16 2.71565
R631 VTAIL.n46 VTAIL.n32 2.71565
R632 VTAIL.n110 VTAIL.n96 2.71565
R633 VTAIL.n94 VTAIL.n80 2.71565
R634 VTAIL.n78 VTAIL.n64 2.71565
R635 VTAIL.n62 VTAIL.n48 2.71565
R636 VTAIL.n124 VTAIL.n123 1.93989
R637 VTAIL.n12 VTAIL.n11 1.93989
R638 VTAIL.n28 VTAIL.n27 1.93989
R639 VTAIL.n44 VTAIL.n43 1.93989
R640 VTAIL.n108 VTAIL.n107 1.93989
R641 VTAIL.n92 VTAIL.n91 1.93989
R642 VTAIL.n76 VTAIL.n75 1.93989
R643 VTAIL.n60 VTAIL.n59 1.93989
R644 VTAIL.n120 VTAIL.n114 1.16414
R645 VTAIL.n8 VTAIL.n2 1.16414
R646 VTAIL.n24 VTAIL.n18 1.16414
R647 VTAIL.n40 VTAIL.n34 1.16414
R648 VTAIL.n104 VTAIL.n98 1.16414
R649 VTAIL.n88 VTAIL.n82 1.16414
R650 VTAIL.n72 VTAIL.n66 1.16414
R651 VTAIL.n56 VTAIL.n50 1.16414
R652 VTAIL.n79 VTAIL.n63 0.810845
R653 VTAIL.n111 VTAIL.n95 0.810845
R654 VTAIL.n47 VTAIL.n31 0.810845
R655 VTAIL.n95 VTAIL.n79 0.470328
R656 VTAIL.n31 VTAIL.n15 0.470328
R657 VTAIL VTAIL.n15 0.463862
R658 VTAIL.n119 VTAIL.n116 0.388379
R659 VTAIL.n7 VTAIL.n4 0.388379
R660 VTAIL.n23 VTAIL.n20 0.388379
R661 VTAIL.n39 VTAIL.n36 0.388379
R662 VTAIL.n103 VTAIL.n100 0.388379
R663 VTAIL.n87 VTAIL.n84 0.388379
R664 VTAIL.n71 VTAIL.n68 0.388379
R665 VTAIL.n55 VTAIL.n52 0.388379
R666 VTAIL VTAIL.n127 0.347483
R667 VTAIL.n118 VTAIL.n113 0.155672
R668 VTAIL.n125 VTAIL.n113 0.155672
R669 VTAIL.n6 VTAIL.n1 0.155672
R670 VTAIL.n13 VTAIL.n1 0.155672
R671 VTAIL.n22 VTAIL.n17 0.155672
R672 VTAIL.n29 VTAIL.n17 0.155672
R673 VTAIL.n38 VTAIL.n33 0.155672
R674 VTAIL.n45 VTAIL.n33 0.155672
R675 VTAIL.n109 VTAIL.n97 0.155672
R676 VTAIL.n102 VTAIL.n97 0.155672
R677 VTAIL.n93 VTAIL.n81 0.155672
R678 VTAIL.n86 VTAIL.n81 0.155672
R679 VTAIL.n77 VTAIL.n65 0.155672
R680 VTAIL.n70 VTAIL.n65 0.155672
R681 VTAIL.n61 VTAIL.n49 0.155672
R682 VTAIL.n54 VTAIL.n49 0.155672
R683 VDD1 VDD1.n1 158.832
R684 VDD1 VDD1.n0 129.46
R685 VDD1.n0 VDD1.t0 10.1583
R686 VDD1.n0 VDD1.t3 10.1583
R687 VDD1.n1 VDD1.t2 10.1583
R688 VDD1.n1 VDD1.t1 10.1583
R689 VN.n0 VN.t3 211.806
R690 VN.n1 VN.t0 211.806
R691 VN.n0 VN.t1 211.782
R692 VN.n1 VN.t2 211.782
R693 VN VN.n1 104.186
R694 VN VN.n0 70.265
R695 VDD2.n2 VDD2.n0 158.306
R696 VDD2.n2 VDD2.n1 129.403
R697 VDD2.n1 VDD2.t1 10.1583
R698 VDD2.n1 VDD2.t3 10.1583
R699 VDD2.n0 VDD2.t0 10.1583
R700 VDD2.n0 VDD2.t2 10.1583
R701 VDD2 VDD2.n2 0.0586897
C0 B VDD1 0.672076f
C1 VP w_n1534_n1608# 2.22431f
C2 B w_n1534_n1608# 4.32251f
C3 VDD2 VN 0.996284f
C4 VDD2 VP 0.273314f
C5 B VDD2 0.692418f
C6 VP VN 3.12802f
C7 B VN 0.620933f
C8 B VP 0.930192f
C9 VDD1 VTAIL 2.94467f
C10 VTAIL w_n1534_n1608# 1.86501f
C11 VDD2 VTAIL 2.98553f
C12 VDD1 w_n1534_n1608# 0.806795f
C13 VTAIL VN 1.01139f
C14 VTAIL VP 1.0255f
C15 VDD1 VDD2 0.548062f
C16 B VTAIL 1.38464f
C17 VDD2 w_n1534_n1608# 0.819078f
C18 VDD1 VN 0.152404f
C19 VN w_n1534_n1608# 2.03415f
C20 VDD1 VP 1.11652f
C21 VDD2 VSUBS 0.42365f
C22 VDD1 VSUBS 2.55616f
C23 VTAIL VSUBS 0.348305f
C24 VN VSUBS 4.08553f
C25 VP VSUBS 0.842283f
C26 B VSUBS 1.720181f
C27 w_n1534_n1608# VSUBS 31.201601f
C28 VDD2.t0 VSUBS 0.052749f
C29 VDD2.t2 VSUBS 0.052749f
C30 VDD2.n0 VSUBS 0.442585f
C31 VDD2.t1 VSUBS 0.052749f
C32 VDD2.t3 VSUBS 0.052749f
C33 VDD2.n1 VSUBS 0.284488f
C34 VDD2.n2 VSUBS 2.00297f
C35 VN.t3 VSUBS 0.324448f
C36 VN.t1 VSUBS 0.324422f
C37 VN.n0 VSUBS 0.31851f
C38 VN.t0 VSUBS 0.324448f
C39 VN.t2 VSUBS 0.324422f
C40 VN.n1 VSUBS 0.824669f
C41 VDD1.t0 VSUBS 0.049714f
C42 VDD1.t3 VSUBS 0.049714f
C43 VDD1.n0 VSUBS 0.268262f
C44 VDD1.t2 VSUBS 0.049714f
C45 VDD1.t1 VSUBS 0.049714f
C46 VDD1.n1 VSUBS 0.426855f
C47 VTAIL.n0 VSUBS 0.016279f
C48 VTAIL.n1 VSUBS 0.015348f
C49 VTAIL.n2 VSUBS 0.008247f
C50 VTAIL.n3 VSUBS 0.01462f
C51 VTAIL.n4 VSUBS 0.012035f
C52 VTAIL.t3 VSUBS 0.043456f
C53 VTAIL.n5 VSUBS 0.055774f
C54 VTAIL.n6 VSUBS 0.15501f
C55 VTAIL.n7 VSUBS 0.008247f
C56 VTAIL.n8 VSUBS 0.008732f
C57 VTAIL.n9 VSUBS 0.019493f
C58 VTAIL.n10 VSUBS 0.0452f
C59 VTAIL.n11 VSUBS 0.008732f
C60 VTAIL.n12 VSUBS 0.008247f
C61 VTAIL.n13 VSUBS 0.037152f
C62 VTAIL.n14 VSUBS 0.022692f
C63 VTAIL.n15 VSUBS 0.060205f
C64 VTAIL.n16 VSUBS 0.016279f
C65 VTAIL.n17 VSUBS 0.015348f
C66 VTAIL.n18 VSUBS 0.008247f
C67 VTAIL.n19 VSUBS 0.01462f
C68 VTAIL.n20 VSUBS 0.012035f
C69 VTAIL.t4 VSUBS 0.043456f
C70 VTAIL.n21 VSUBS 0.055774f
C71 VTAIL.n22 VSUBS 0.15501f
C72 VTAIL.n23 VSUBS 0.008247f
C73 VTAIL.n24 VSUBS 0.008732f
C74 VTAIL.n25 VSUBS 0.019493f
C75 VTAIL.n26 VSUBS 0.0452f
C76 VTAIL.n27 VSUBS 0.008732f
C77 VTAIL.n28 VSUBS 0.008247f
C78 VTAIL.n29 VSUBS 0.037152f
C79 VTAIL.n30 VSUBS 0.022692f
C80 VTAIL.n31 VSUBS 0.077365f
C81 VTAIL.n32 VSUBS 0.016279f
C82 VTAIL.n33 VSUBS 0.015348f
C83 VTAIL.n34 VSUBS 0.008247f
C84 VTAIL.n35 VSUBS 0.01462f
C85 VTAIL.n36 VSUBS 0.012035f
C86 VTAIL.t6 VSUBS 0.043456f
C87 VTAIL.n37 VSUBS 0.055774f
C88 VTAIL.n38 VSUBS 0.15501f
C89 VTAIL.n39 VSUBS 0.008247f
C90 VTAIL.n40 VSUBS 0.008732f
C91 VTAIL.n41 VSUBS 0.019493f
C92 VTAIL.n42 VSUBS 0.0452f
C93 VTAIL.n43 VSUBS 0.008732f
C94 VTAIL.n44 VSUBS 0.008247f
C95 VTAIL.n45 VSUBS 0.037152f
C96 VTAIL.n46 VSUBS 0.022692f
C97 VTAIL.n47 VSUBS 0.439106f
C98 VTAIL.n48 VSUBS 0.016279f
C99 VTAIL.n49 VSUBS 0.015348f
C100 VTAIL.n50 VSUBS 0.008247f
C101 VTAIL.n51 VSUBS 0.01462f
C102 VTAIL.n52 VSUBS 0.012035f
C103 VTAIL.t0 VSUBS 0.043456f
C104 VTAIL.n53 VSUBS 0.055774f
C105 VTAIL.n54 VSUBS 0.15501f
C106 VTAIL.n55 VSUBS 0.008247f
C107 VTAIL.n56 VSUBS 0.008732f
C108 VTAIL.n57 VSUBS 0.019493f
C109 VTAIL.n58 VSUBS 0.0452f
C110 VTAIL.n59 VSUBS 0.008732f
C111 VTAIL.n60 VSUBS 0.008247f
C112 VTAIL.n61 VSUBS 0.037152f
C113 VTAIL.n62 VSUBS 0.022692f
C114 VTAIL.n63 VSUBS 0.439106f
C115 VTAIL.n64 VSUBS 0.016279f
C116 VTAIL.n65 VSUBS 0.015348f
C117 VTAIL.n66 VSUBS 0.008247f
C118 VTAIL.n67 VSUBS 0.01462f
C119 VTAIL.n68 VSUBS 0.012035f
C120 VTAIL.t1 VSUBS 0.043456f
C121 VTAIL.n69 VSUBS 0.055774f
C122 VTAIL.n70 VSUBS 0.15501f
C123 VTAIL.n71 VSUBS 0.008247f
C124 VTAIL.n72 VSUBS 0.008732f
C125 VTAIL.n73 VSUBS 0.019493f
C126 VTAIL.n74 VSUBS 0.0452f
C127 VTAIL.n75 VSUBS 0.008732f
C128 VTAIL.n76 VSUBS 0.008247f
C129 VTAIL.n77 VSUBS 0.037152f
C130 VTAIL.n78 VSUBS 0.022692f
C131 VTAIL.n79 VSUBS 0.077365f
C132 VTAIL.n80 VSUBS 0.016279f
C133 VTAIL.n81 VSUBS 0.015348f
C134 VTAIL.n82 VSUBS 0.008247f
C135 VTAIL.n83 VSUBS 0.01462f
C136 VTAIL.n84 VSUBS 0.012035f
C137 VTAIL.t5 VSUBS 0.043456f
C138 VTAIL.n85 VSUBS 0.055774f
C139 VTAIL.n86 VSUBS 0.15501f
C140 VTAIL.n87 VSUBS 0.008247f
C141 VTAIL.n88 VSUBS 0.008732f
C142 VTAIL.n89 VSUBS 0.019493f
C143 VTAIL.n90 VSUBS 0.0452f
C144 VTAIL.n91 VSUBS 0.008732f
C145 VTAIL.n92 VSUBS 0.008247f
C146 VTAIL.n93 VSUBS 0.037152f
C147 VTAIL.n94 VSUBS 0.022692f
C148 VTAIL.n95 VSUBS 0.077365f
C149 VTAIL.n96 VSUBS 0.016279f
C150 VTAIL.n97 VSUBS 0.015348f
C151 VTAIL.n98 VSUBS 0.008247f
C152 VTAIL.n99 VSUBS 0.01462f
C153 VTAIL.n100 VSUBS 0.012035f
C154 VTAIL.t7 VSUBS 0.043456f
C155 VTAIL.n101 VSUBS 0.055774f
C156 VTAIL.n102 VSUBS 0.15501f
C157 VTAIL.n103 VSUBS 0.008247f
C158 VTAIL.n104 VSUBS 0.008732f
C159 VTAIL.n105 VSUBS 0.019493f
C160 VTAIL.n106 VSUBS 0.0452f
C161 VTAIL.n107 VSUBS 0.008732f
C162 VTAIL.n108 VSUBS 0.008247f
C163 VTAIL.n109 VSUBS 0.037152f
C164 VTAIL.n110 VSUBS 0.022692f
C165 VTAIL.n111 VSUBS 0.439106f
C166 VTAIL.n112 VSUBS 0.016279f
C167 VTAIL.n113 VSUBS 0.015348f
C168 VTAIL.n114 VSUBS 0.008247f
C169 VTAIL.n115 VSUBS 0.01462f
C170 VTAIL.n116 VSUBS 0.012035f
C171 VTAIL.t2 VSUBS 0.043456f
C172 VTAIL.n117 VSUBS 0.055774f
C173 VTAIL.n118 VSUBS 0.15501f
C174 VTAIL.n119 VSUBS 0.008247f
C175 VTAIL.n120 VSUBS 0.008732f
C176 VTAIL.n121 VSUBS 0.019493f
C177 VTAIL.n122 VSUBS 0.0452f
C178 VTAIL.n123 VSUBS 0.008732f
C179 VTAIL.n124 VSUBS 0.008247f
C180 VTAIL.n125 VSUBS 0.037152f
C181 VTAIL.n126 VSUBS 0.022692f
C182 VTAIL.n127 VSUBS 0.416191f
C183 VP.t0 VSUBS 0.342109f
C184 VP.t3 VSUBS 0.342137f
C185 VP.n0 VSUBS 0.853602f
C186 VP.n1 VSUBS 2.66785f
C187 VP.t1 VSUBS 0.323673f
C188 VP.n2 VSUBS 0.186301f
C189 VP.t2 VSUBS 0.323673f
C190 VP.n3 VSUBS 0.186301f
C191 VP.n4 VSUBS 0.043029f
C192 B.n0 VSUBS 0.00698f
C193 B.n1 VSUBS 0.00698f
C194 B.n2 VSUBS 0.010323f
C195 B.n3 VSUBS 0.00791f
C196 B.n4 VSUBS 0.00791f
C197 B.n5 VSUBS 0.00791f
C198 B.n6 VSUBS 0.00791f
C199 B.n7 VSUBS 0.00791f
C200 B.n8 VSUBS 0.00791f
C201 B.n9 VSUBS 0.00791f
C202 B.n10 VSUBS 0.018511f
C203 B.n11 VSUBS 0.00791f
C204 B.n12 VSUBS 0.00791f
C205 B.n13 VSUBS 0.00791f
C206 B.n14 VSUBS 0.00791f
C207 B.n15 VSUBS 0.00791f
C208 B.n16 VSUBS 0.00791f
C209 B.n17 VSUBS 0.00791f
C210 B.t1 VSUBS 0.053257f
C211 B.t2 VSUBS 0.059961f
C212 B.t0 VSUBS 0.099566f
C213 B.n18 VSUBS 0.109135f
C214 B.n19 VSUBS 0.10094f
C215 B.n20 VSUBS 0.018327f
C216 B.n21 VSUBS 0.00791f
C217 B.n22 VSUBS 0.00791f
C218 B.n23 VSUBS 0.00791f
C219 B.n24 VSUBS 0.00791f
C220 B.n25 VSUBS 0.00791f
C221 B.t7 VSUBS 0.053257f
C222 B.t8 VSUBS 0.059962f
C223 B.t6 VSUBS 0.099566f
C224 B.n26 VSUBS 0.109135f
C225 B.n27 VSUBS 0.100939f
C226 B.n28 VSUBS 0.00791f
C227 B.n29 VSUBS 0.00791f
C228 B.n30 VSUBS 0.00791f
C229 B.n31 VSUBS 0.00791f
C230 B.n32 VSUBS 0.00791f
C231 B.n33 VSUBS 0.00791f
C232 B.n34 VSUBS 0.00791f
C233 B.n35 VSUBS 0.017783f
C234 B.n36 VSUBS 0.00791f
C235 B.n37 VSUBS 0.00791f
C236 B.n38 VSUBS 0.00791f
C237 B.n39 VSUBS 0.00791f
C238 B.n40 VSUBS 0.00791f
C239 B.n41 VSUBS 0.00791f
C240 B.n42 VSUBS 0.00791f
C241 B.n43 VSUBS 0.00791f
C242 B.n44 VSUBS 0.00791f
C243 B.n45 VSUBS 0.00791f
C244 B.n46 VSUBS 0.00791f
C245 B.n47 VSUBS 0.00791f
C246 B.n48 VSUBS 0.00791f
C247 B.n49 VSUBS 0.00791f
C248 B.n50 VSUBS 0.00791f
C249 B.n51 VSUBS 0.00791f
C250 B.n52 VSUBS 0.017548f
C251 B.n53 VSUBS 0.00791f
C252 B.n54 VSUBS 0.00791f
C253 B.n55 VSUBS 0.00791f
C254 B.n56 VSUBS 0.00791f
C255 B.n57 VSUBS 0.00791f
C256 B.n58 VSUBS 0.00791f
C257 B.n59 VSUBS 0.00791f
C258 B.t5 VSUBS 0.053257f
C259 B.t4 VSUBS 0.059962f
C260 B.t3 VSUBS 0.099566f
C261 B.n60 VSUBS 0.109135f
C262 B.n61 VSUBS 0.100939f
C263 B.n62 VSUBS 0.018327f
C264 B.n63 VSUBS 0.00791f
C265 B.n64 VSUBS 0.00791f
C266 B.n65 VSUBS 0.00791f
C267 B.n66 VSUBS 0.00791f
C268 B.n67 VSUBS 0.00791f
C269 B.t11 VSUBS 0.053257f
C270 B.t10 VSUBS 0.059961f
C271 B.t9 VSUBS 0.099566f
C272 B.n68 VSUBS 0.109135f
C273 B.n69 VSUBS 0.10094f
C274 B.n70 VSUBS 0.00791f
C275 B.n71 VSUBS 0.00791f
C276 B.n72 VSUBS 0.00791f
C277 B.n73 VSUBS 0.00791f
C278 B.n74 VSUBS 0.00791f
C279 B.n75 VSUBS 0.00791f
C280 B.n76 VSUBS 0.00791f
C281 B.n77 VSUBS 0.017783f
C282 B.n78 VSUBS 0.00791f
C283 B.n79 VSUBS 0.00791f
C284 B.n80 VSUBS 0.00791f
C285 B.n81 VSUBS 0.00791f
C286 B.n82 VSUBS 0.00791f
C287 B.n83 VSUBS 0.00791f
C288 B.n84 VSUBS 0.00791f
C289 B.n85 VSUBS 0.00791f
C290 B.n86 VSUBS 0.00791f
C291 B.n87 VSUBS 0.00791f
C292 B.n88 VSUBS 0.00791f
C293 B.n89 VSUBS 0.00791f
C294 B.n90 VSUBS 0.00791f
C295 B.n91 VSUBS 0.00791f
C296 B.n92 VSUBS 0.00791f
C297 B.n93 VSUBS 0.00791f
C298 B.n94 VSUBS 0.00791f
C299 B.n95 VSUBS 0.00791f
C300 B.n96 VSUBS 0.00791f
C301 B.n97 VSUBS 0.00791f
C302 B.n98 VSUBS 0.00791f
C303 B.n99 VSUBS 0.00791f
C304 B.n100 VSUBS 0.00791f
C305 B.n101 VSUBS 0.00791f
C306 B.n102 VSUBS 0.00791f
C307 B.n103 VSUBS 0.00791f
C308 B.n104 VSUBS 0.00791f
C309 B.n105 VSUBS 0.00791f
C310 B.n106 VSUBS 0.017783f
C311 B.n107 VSUBS 0.018511f
C312 B.n108 VSUBS 0.018511f
C313 B.n109 VSUBS 0.00791f
C314 B.n110 VSUBS 0.00791f
C315 B.n111 VSUBS 0.00791f
C316 B.n112 VSUBS 0.00791f
C317 B.n113 VSUBS 0.00791f
C318 B.n114 VSUBS 0.00791f
C319 B.n115 VSUBS 0.00791f
C320 B.n116 VSUBS 0.00791f
C321 B.n117 VSUBS 0.00791f
C322 B.n118 VSUBS 0.00791f
C323 B.n119 VSUBS 0.00791f
C324 B.n120 VSUBS 0.00791f
C325 B.n121 VSUBS 0.00791f
C326 B.n122 VSUBS 0.00791f
C327 B.n123 VSUBS 0.00791f
C328 B.n124 VSUBS 0.00791f
C329 B.n125 VSUBS 0.00791f
C330 B.n126 VSUBS 0.00791f
C331 B.n127 VSUBS 0.00791f
C332 B.n128 VSUBS 0.00791f
C333 B.n129 VSUBS 0.00791f
C334 B.n130 VSUBS 0.005467f
C335 B.n131 VSUBS 0.018327f
C336 B.n132 VSUBS 0.006398f
C337 B.n133 VSUBS 0.00791f
C338 B.n134 VSUBS 0.00791f
C339 B.n135 VSUBS 0.00791f
C340 B.n136 VSUBS 0.00791f
C341 B.n137 VSUBS 0.00791f
C342 B.n138 VSUBS 0.00791f
C343 B.n139 VSUBS 0.00791f
C344 B.n140 VSUBS 0.00791f
C345 B.n141 VSUBS 0.00791f
C346 B.n142 VSUBS 0.00791f
C347 B.n143 VSUBS 0.00791f
C348 B.n144 VSUBS 0.006398f
C349 B.n145 VSUBS 0.00791f
C350 B.n146 VSUBS 0.00791f
C351 B.n147 VSUBS 0.005467f
C352 B.n148 VSUBS 0.00791f
C353 B.n149 VSUBS 0.00791f
C354 B.n150 VSUBS 0.00791f
C355 B.n151 VSUBS 0.00791f
C356 B.n152 VSUBS 0.00791f
C357 B.n153 VSUBS 0.00791f
C358 B.n154 VSUBS 0.00791f
C359 B.n155 VSUBS 0.00791f
C360 B.n156 VSUBS 0.00791f
C361 B.n157 VSUBS 0.00791f
C362 B.n158 VSUBS 0.00791f
C363 B.n159 VSUBS 0.00791f
C364 B.n160 VSUBS 0.00791f
C365 B.n161 VSUBS 0.00791f
C366 B.n162 VSUBS 0.00791f
C367 B.n163 VSUBS 0.00791f
C368 B.n164 VSUBS 0.00791f
C369 B.n165 VSUBS 0.00791f
C370 B.n166 VSUBS 0.00791f
C371 B.n167 VSUBS 0.00791f
C372 B.n168 VSUBS 0.00791f
C373 B.n169 VSUBS 0.018511f
C374 B.n170 VSUBS 0.017783f
C375 B.n171 VSUBS 0.018746f
C376 B.n172 VSUBS 0.00791f
C377 B.n173 VSUBS 0.00791f
C378 B.n174 VSUBS 0.00791f
C379 B.n175 VSUBS 0.00791f
C380 B.n176 VSUBS 0.00791f
C381 B.n177 VSUBS 0.00791f
C382 B.n178 VSUBS 0.00791f
C383 B.n179 VSUBS 0.00791f
C384 B.n180 VSUBS 0.00791f
C385 B.n181 VSUBS 0.00791f
C386 B.n182 VSUBS 0.00791f
C387 B.n183 VSUBS 0.00791f
C388 B.n184 VSUBS 0.00791f
C389 B.n185 VSUBS 0.00791f
C390 B.n186 VSUBS 0.00791f
C391 B.n187 VSUBS 0.00791f
C392 B.n188 VSUBS 0.00791f
C393 B.n189 VSUBS 0.00791f
C394 B.n190 VSUBS 0.00791f
C395 B.n191 VSUBS 0.00791f
C396 B.n192 VSUBS 0.00791f
C397 B.n193 VSUBS 0.00791f
C398 B.n194 VSUBS 0.00791f
C399 B.n195 VSUBS 0.00791f
C400 B.n196 VSUBS 0.00791f
C401 B.n197 VSUBS 0.00791f
C402 B.n198 VSUBS 0.00791f
C403 B.n199 VSUBS 0.00791f
C404 B.n200 VSUBS 0.00791f
C405 B.n201 VSUBS 0.00791f
C406 B.n202 VSUBS 0.00791f
C407 B.n203 VSUBS 0.00791f
C408 B.n204 VSUBS 0.00791f
C409 B.n205 VSUBS 0.00791f
C410 B.n206 VSUBS 0.00791f
C411 B.n207 VSUBS 0.00791f
C412 B.n208 VSUBS 0.00791f
C413 B.n209 VSUBS 0.00791f
C414 B.n210 VSUBS 0.00791f
C415 B.n211 VSUBS 0.00791f
C416 B.n212 VSUBS 0.00791f
C417 B.n213 VSUBS 0.00791f
C418 B.n214 VSUBS 0.00791f
C419 B.n215 VSUBS 0.00791f
C420 B.n216 VSUBS 0.00791f
C421 B.n217 VSUBS 0.00791f
C422 B.n218 VSUBS 0.00791f
C423 B.n219 VSUBS 0.00791f
C424 B.n220 VSUBS 0.017783f
C425 B.n221 VSUBS 0.018511f
C426 B.n222 VSUBS 0.018511f
C427 B.n223 VSUBS 0.00791f
C428 B.n224 VSUBS 0.00791f
C429 B.n225 VSUBS 0.00791f
C430 B.n226 VSUBS 0.00791f
C431 B.n227 VSUBS 0.00791f
C432 B.n228 VSUBS 0.00791f
C433 B.n229 VSUBS 0.00791f
C434 B.n230 VSUBS 0.00791f
C435 B.n231 VSUBS 0.00791f
C436 B.n232 VSUBS 0.00791f
C437 B.n233 VSUBS 0.00791f
C438 B.n234 VSUBS 0.00791f
C439 B.n235 VSUBS 0.00791f
C440 B.n236 VSUBS 0.00791f
C441 B.n237 VSUBS 0.00791f
C442 B.n238 VSUBS 0.00791f
C443 B.n239 VSUBS 0.00791f
C444 B.n240 VSUBS 0.00791f
C445 B.n241 VSUBS 0.00791f
C446 B.n242 VSUBS 0.00791f
C447 B.n243 VSUBS 0.00791f
C448 B.n244 VSUBS 0.005467f
C449 B.n245 VSUBS 0.018327f
C450 B.n246 VSUBS 0.006398f
C451 B.n247 VSUBS 0.00791f
C452 B.n248 VSUBS 0.00791f
C453 B.n249 VSUBS 0.00791f
C454 B.n250 VSUBS 0.00791f
C455 B.n251 VSUBS 0.00791f
C456 B.n252 VSUBS 0.00791f
C457 B.n253 VSUBS 0.00791f
C458 B.n254 VSUBS 0.00791f
C459 B.n255 VSUBS 0.00791f
C460 B.n256 VSUBS 0.00791f
C461 B.n257 VSUBS 0.00791f
C462 B.n258 VSUBS 0.006398f
C463 B.n259 VSUBS 0.00791f
C464 B.n260 VSUBS 0.00791f
C465 B.n261 VSUBS 0.005467f
C466 B.n262 VSUBS 0.00791f
C467 B.n263 VSUBS 0.00791f
C468 B.n264 VSUBS 0.00791f
C469 B.n265 VSUBS 0.00791f
C470 B.n266 VSUBS 0.00791f
C471 B.n267 VSUBS 0.00791f
C472 B.n268 VSUBS 0.00791f
C473 B.n269 VSUBS 0.00791f
C474 B.n270 VSUBS 0.00791f
C475 B.n271 VSUBS 0.00791f
C476 B.n272 VSUBS 0.00791f
C477 B.n273 VSUBS 0.00791f
C478 B.n274 VSUBS 0.00791f
C479 B.n275 VSUBS 0.00791f
C480 B.n276 VSUBS 0.00791f
C481 B.n277 VSUBS 0.00791f
C482 B.n278 VSUBS 0.00791f
C483 B.n279 VSUBS 0.00791f
C484 B.n280 VSUBS 0.00791f
C485 B.n281 VSUBS 0.00791f
C486 B.n282 VSUBS 0.00791f
C487 B.n283 VSUBS 0.018511f
C488 B.n284 VSUBS 0.017783f
C489 B.n285 VSUBS 0.017783f
C490 B.n286 VSUBS 0.00791f
C491 B.n287 VSUBS 0.00791f
C492 B.n288 VSUBS 0.00791f
C493 B.n289 VSUBS 0.00791f
C494 B.n290 VSUBS 0.00791f
C495 B.n291 VSUBS 0.00791f
C496 B.n292 VSUBS 0.00791f
C497 B.n293 VSUBS 0.00791f
C498 B.n294 VSUBS 0.00791f
C499 B.n295 VSUBS 0.00791f
C500 B.n296 VSUBS 0.00791f
C501 B.n297 VSUBS 0.00791f
C502 B.n298 VSUBS 0.00791f
C503 B.n299 VSUBS 0.00791f
C504 B.n300 VSUBS 0.00791f
C505 B.n301 VSUBS 0.00791f
C506 B.n302 VSUBS 0.00791f
C507 B.n303 VSUBS 0.00791f
C508 B.n304 VSUBS 0.00791f
C509 B.n305 VSUBS 0.00791f
C510 B.n306 VSUBS 0.00791f
C511 B.n307 VSUBS 0.010323f
C512 B.n308 VSUBS 0.010996f
C513 B.n309 VSUBS 0.021867f
.ends

