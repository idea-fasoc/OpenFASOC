* NGSPICE file created from diff_pair_sample_0791.ext - technology: sky130A

.subckt diff_pair_sample_0791 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t7 w_n3234_n2520# sky130_fd_pr__pfet_01v8 ad=1.2804 pd=8.09 as=3.0264 ps=16.3 w=7.76 l=2.5
X1 VTAIL.t9 VP.t1 VDD1.t4 w_n3234_n2520# sky130_fd_pr__pfet_01v8 ad=1.2804 pd=8.09 as=1.2804 ps=8.09 w=7.76 l=2.5
X2 VDD2.t5 VN.t0 VTAIL.t0 w_n3234_n2520# sky130_fd_pr__pfet_01v8 ad=3.0264 pd=16.3 as=1.2804 ps=8.09 w=7.76 l=2.5
X3 B.t11 B.t9 B.t10 w_n3234_n2520# sky130_fd_pr__pfet_01v8 ad=3.0264 pd=16.3 as=0 ps=0 w=7.76 l=2.5
X4 B.t8 B.t6 B.t7 w_n3234_n2520# sky130_fd_pr__pfet_01v8 ad=3.0264 pd=16.3 as=0 ps=0 w=7.76 l=2.5
X5 VDD1.t3 VP.t2 VTAIL.t11 w_n3234_n2520# sky130_fd_pr__pfet_01v8 ad=1.2804 pd=8.09 as=3.0264 ps=16.3 w=7.76 l=2.5
X6 B.t5 B.t3 B.t4 w_n3234_n2520# sky130_fd_pr__pfet_01v8 ad=3.0264 pd=16.3 as=0 ps=0 w=7.76 l=2.5
X7 VDD2.t4 VN.t1 VTAIL.t5 w_n3234_n2520# sky130_fd_pr__pfet_01v8 ad=1.2804 pd=8.09 as=3.0264 ps=16.3 w=7.76 l=2.5
X8 B.t2 B.t0 B.t1 w_n3234_n2520# sky130_fd_pr__pfet_01v8 ad=3.0264 pd=16.3 as=0 ps=0 w=7.76 l=2.5
X9 VTAIL.t4 VN.t2 VDD2.t3 w_n3234_n2520# sky130_fd_pr__pfet_01v8 ad=1.2804 pd=8.09 as=1.2804 ps=8.09 w=7.76 l=2.5
X10 VTAIL.t2 VN.t3 VDD2.t2 w_n3234_n2520# sky130_fd_pr__pfet_01v8 ad=1.2804 pd=8.09 as=1.2804 ps=8.09 w=7.76 l=2.5
X11 VDD2.t1 VN.t4 VTAIL.t1 w_n3234_n2520# sky130_fd_pr__pfet_01v8 ad=1.2804 pd=8.09 as=3.0264 ps=16.3 w=7.76 l=2.5
X12 VDD1.t2 VP.t3 VTAIL.t6 w_n3234_n2520# sky130_fd_pr__pfet_01v8 ad=3.0264 pd=16.3 as=1.2804 ps=8.09 w=7.76 l=2.5
X13 VDD1.t1 VP.t4 VTAIL.t8 w_n3234_n2520# sky130_fd_pr__pfet_01v8 ad=3.0264 pd=16.3 as=1.2804 ps=8.09 w=7.76 l=2.5
X14 VDD2.t0 VN.t5 VTAIL.t3 w_n3234_n2520# sky130_fd_pr__pfet_01v8 ad=3.0264 pd=16.3 as=1.2804 ps=8.09 w=7.76 l=2.5
X15 VTAIL.t10 VP.t5 VDD1.t0 w_n3234_n2520# sky130_fd_pr__pfet_01v8 ad=1.2804 pd=8.09 as=1.2804 ps=8.09 w=7.76 l=2.5
R0 VP.n13 VP.n12 161.3
R1 VP.n14 VP.n9 161.3
R2 VP.n16 VP.n15 161.3
R3 VP.n17 VP.n8 161.3
R4 VP.n19 VP.n18 161.3
R5 VP.n20 VP.n7 161.3
R6 VP.n42 VP.n0 161.3
R7 VP.n41 VP.n40 161.3
R8 VP.n39 VP.n1 161.3
R9 VP.n38 VP.n37 161.3
R10 VP.n36 VP.n2 161.3
R11 VP.n35 VP.n34 161.3
R12 VP.n33 VP.n32 161.3
R13 VP.n31 VP.n4 161.3
R14 VP.n30 VP.n29 161.3
R15 VP.n28 VP.n5 161.3
R16 VP.n27 VP.n26 161.3
R17 VP.n25 VP.n6 161.3
R18 VP.n24 VP.n23 106.974
R19 VP.n44 VP.n43 106.974
R20 VP.n22 VP.n21 106.974
R21 VP.n11 VP.t4 106.558
R22 VP.n24 VP.t3 74.8069
R23 VP.n3 VP.t5 74.8069
R24 VP.n43 VP.t2 74.8069
R25 VP.n21 VP.t0 74.8069
R26 VP.n10 VP.t1 74.8069
R27 VP.n11 VP.n10 60.0034
R28 VP.n30 VP.n5 56.5617
R29 VP.n37 VP.n1 56.5617
R30 VP.n15 VP.n8 56.5617
R31 VP.n23 VP.n22 44.9731
R32 VP.n26 VP.n25 24.5923
R33 VP.n26 VP.n5 24.5923
R34 VP.n31 VP.n30 24.5923
R35 VP.n32 VP.n31 24.5923
R36 VP.n36 VP.n35 24.5923
R37 VP.n37 VP.n36 24.5923
R38 VP.n41 VP.n1 24.5923
R39 VP.n42 VP.n41 24.5923
R40 VP.n19 VP.n8 24.5923
R41 VP.n20 VP.n19 24.5923
R42 VP.n14 VP.n13 24.5923
R43 VP.n15 VP.n14 24.5923
R44 VP.n32 VP.n3 12.2964
R45 VP.n35 VP.n3 12.2964
R46 VP.n13 VP.n10 12.2964
R47 VP.n12 VP.n11 7.21347
R48 VP.n25 VP.n24 3.93519
R49 VP.n43 VP.n42 3.93519
R50 VP.n21 VP.n20 3.93519
R51 VP.n22 VP.n7 0.278335
R52 VP.n23 VP.n6 0.278335
R53 VP.n44 VP.n0 0.278335
R54 VP.n12 VP.n9 0.189894
R55 VP.n16 VP.n9 0.189894
R56 VP.n17 VP.n16 0.189894
R57 VP.n18 VP.n17 0.189894
R58 VP.n18 VP.n7 0.189894
R59 VP.n27 VP.n6 0.189894
R60 VP.n28 VP.n27 0.189894
R61 VP.n29 VP.n28 0.189894
R62 VP.n29 VP.n4 0.189894
R63 VP.n33 VP.n4 0.189894
R64 VP.n34 VP.n33 0.189894
R65 VP.n34 VP.n2 0.189894
R66 VP.n38 VP.n2 0.189894
R67 VP.n39 VP.n38 0.189894
R68 VP.n40 VP.n39 0.189894
R69 VP.n40 VP.n0 0.189894
R70 VP VP.n44 0.153485
R71 VTAIL.n10 VTAIL.t7 70.7163
R72 VTAIL.n7 VTAIL.t5 70.7163
R73 VTAIL.n11 VTAIL.t1 70.7161
R74 VTAIL.n2 VTAIL.t11 70.7161
R75 VTAIL.n9 VTAIL.n8 66.5275
R76 VTAIL.n6 VTAIL.n5 66.5275
R77 VTAIL.n1 VTAIL.n0 66.5275
R78 VTAIL.n4 VTAIL.n3 66.5275
R79 VTAIL.n6 VTAIL.n4 23.9358
R80 VTAIL.n11 VTAIL.n10 21.4962
R81 VTAIL.n0 VTAIL.t0 4.18929
R82 VTAIL.n0 VTAIL.t2 4.18929
R83 VTAIL.n3 VTAIL.t6 4.18929
R84 VTAIL.n3 VTAIL.t10 4.18929
R85 VTAIL.n8 VTAIL.t8 4.18929
R86 VTAIL.n8 VTAIL.t9 4.18929
R87 VTAIL.n5 VTAIL.t3 4.18929
R88 VTAIL.n5 VTAIL.t4 4.18929
R89 VTAIL.n7 VTAIL.n6 2.44016
R90 VTAIL.n10 VTAIL.n9 2.44016
R91 VTAIL.n4 VTAIL.n2 2.44016
R92 VTAIL VTAIL.n11 1.77205
R93 VTAIL.n9 VTAIL.n7 1.69016
R94 VTAIL.n2 VTAIL.n1 1.69016
R95 VTAIL VTAIL.n1 0.668603
R96 VDD1 VDD1.t1 89.283
R97 VDD1.n1 VDD1.t2 89.1693
R98 VDD1.n1 VDD1.n0 83.7608
R99 VDD1.n3 VDD1.n2 83.2063
R100 VDD1.n3 VDD1.n1 40.1367
R101 VDD1.n2 VDD1.t4 4.18929
R102 VDD1.n2 VDD1.t5 4.18929
R103 VDD1.n0 VDD1.t0 4.18929
R104 VDD1.n0 VDD1.t3 4.18929
R105 VDD1 VDD1.n3 0.552224
R106 VN.n29 VN.n16 161.3
R107 VN.n28 VN.n27 161.3
R108 VN.n26 VN.n17 161.3
R109 VN.n25 VN.n24 161.3
R110 VN.n23 VN.n18 161.3
R111 VN.n22 VN.n21 161.3
R112 VN.n13 VN.n0 161.3
R113 VN.n12 VN.n11 161.3
R114 VN.n10 VN.n1 161.3
R115 VN.n9 VN.n8 161.3
R116 VN.n7 VN.n2 161.3
R117 VN.n6 VN.n5 161.3
R118 VN.n15 VN.n14 106.974
R119 VN.n31 VN.n30 106.974
R120 VN.n4 VN.t0 106.558
R121 VN.n20 VN.t1 106.558
R122 VN.n3 VN.t3 74.8069
R123 VN.n14 VN.t4 74.8069
R124 VN.n19 VN.t2 74.8069
R125 VN.n30 VN.t5 74.8069
R126 VN.n4 VN.n3 60.0034
R127 VN.n20 VN.n19 60.0034
R128 VN.n8 VN.n1 56.5617
R129 VN.n24 VN.n17 56.5617
R130 VN VN.n31 45.252
R131 VN.n7 VN.n6 24.5923
R132 VN.n8 VN.n7 24.5923
R133 VN.n12 VN.n1 24.5923
R134 VN.n13 VN.n12 24.5923
R135 VN.n24 VN.n23 24.5923
R136 VN.n23 VN.n22 24.5923
R137 VN.n29 VN.n28 24.5923
R138 VN.n28 VN.n17 24.5923
R139 VN.n6 VN.n3 12.2964
R140 VN.n22 VN.n19 12.2964
R141 VN.n21 VN.n20 7.21347
R142 VN.n5 VN.n4 7.21347
R143 VN.n14 VN.n13 3.93519
R144 VN.n30 VN.n29 3.93519
R145 VN.n31 VN.n16 0.278335
R146 VN.n15 VN.n0 0.278335
R147 VN.n27 VN.n16 0.189894
R148 VN.n27 VN.n26 0.189894
R149 VN.n26 VN.n25 0.189894
R150 VN.n25 VN.n18 0.189894
R151 VN.n21 VN.n18 0.189894
R152 VN.n5 VN.n2 0.189894
R153 VN.n9 VN.n2 0.189894
R154 VN.n10 VN.n9 0.189894
R155 VN.n11 VN.n10 0.189894
R156 VN.n11 VN.n0 0.189894
R157 VN VN.n15 0.153485
R158 VDD2.n1 VDD2.t5 89.1693
R159 VDD2.n2 VDD2.t0 87.3951
R160 VDD2.n1 VDD2.n0 83.7608
R161 VDD2 VDD2.n3 83.758
R162 VDD2.n2 VDD2.n1 38.3338
R163 VDD2.n3 VDD2.t3 4.18929
R164 VDD2.n3 VDD2.t4 4.18929
R165 VDD2.n0 VDD2.t2 4.18929
R166 VDD2.n0 VDD2.t1 4.18929
R167 VDD2 VDD2.n2 1.88843
R168 B.n324 B.n103 585
R169 B.n323 B.n322 585
R170 B.n321 B.n104 585
R171 B.n320 B.n319 585
R172 B.n318 B.n105 585
R173 B.n317 B.n316 585
R174 B.n315 B.n106 585
R175 B.n314 B.n313 585
R176 B.n312 B.n107 585
R177 B.n311 B.n310 585
R178 B.n309 B.n108 585
R179 B.n308 B.n307 585
R180 B.n306 B.n109 585
R181 B.n305 B.n304 585
R182 B.n303 B.n110 585
R183 B.n302 B.n301 585
R184 B.n300 B.n111 585
R185 B.n299 B.n298 585
R186 B.n297 B.n112 585
R187 B.n296 B.n295 585
R188 B.n294 B.n113 585
R189 B.n293 B.n292 585
R190 B.n291 B.n114 585
R191 B.n290 B.n289 585
R192 B.n288 B.n115 585
R193 B.n287 B.n286 585
R194 B.n285 B.n116 585
R195 B.n284 B.n283 585
R196 B.n282 B.n117 585
R197 B.n280 B.n279 585
R198 B.n278 B.n120 585
R199 B.n277 B.n276 585
R200 B.n275 B.n121 585
R201 B.n274 B.n273 585
R202 B.n272 B.n122 585
R203 B.n271 B.n270 585
R204 B.n269 B.n123 585
R205 B.n268 B.n267 585
R206 B.n266 B.n124 585
R207 B.n265 B.n264 585
R208 B.n260 B.n125 585
R209 B.n259 B.n258 585
R210 B.n257 B.n126 585
R211 B.n256 B.n255 585
R212 B.n254 B.n127 585
R213 B.n253 B.n252 585
R214 B.n251 B.n128 585
R215 B.n250 B.n249 585
R216 B.n248 B.n129 585
R217 B.n247 B.n246 585
R218 B.n245 B.n130 585
R219 B.n244 B.n243 585
R220 B.n242 B.n131 585
R221 B.n241 B.n240 585
R222 B.n239 B.n132 585
R223 B.n238 B.n237 585
R224 B.n236 B.n133 585
R225 B.n235 B.n234 585
R226 B.n233 B.n134 585
R227 B.n232 B.n231 585
R228 B.n230 B.n135 585
R229 B.n229 B.n228 585
R230 B.n227 B.n136 585
R231 B.n226 B.n225 585
R232 B.n224 B.n137 585
R233 B.n223 B.n222 585
R234 B.n221 B.n138 585
R235 B.n220 B.n219 585
R236 B.n326 B.n325 585
R237 B.n327 B.n102 585
R238 B.n329 B.n328 585
R239 B.n330 B.n101 585
R240 B.n332 B.n331 585
R241 B.n333 B.n100 585
R242 B.n335 B.n334 585
R243 B.n336 B.n99 585
R244 B.n338 B.n337 585
R245 B.n339 B.n98 585
R246 B.n341 B.n340 585
R247 B.n342 B.n97 585
R248 B.n344 B.n343 585
R249 B.n345 B.n96 585
R250 B.n347 B.n346 585
R251 B.n348 B.n95 585
R252 B.n350 B.n349 585
R253 B.n351 B.n94 585
R254 B.n353 B.n352 585
R255 B.n354 B.n93 585
R256 B.n356 B.n355 585
R257 B.n357 B.n92 585
R258 B.n359 B.n358 585
R259 B.n360 B.n91 585
R260 B.n362 B.n361 585
R261 B.n363 B.n90 585
R262 B.n365 B.n364 585
R263 B.n366 B.n89 585
R264 B.n368 B.n367 585
R265 B.n369 B.n88 585
R266 B.n371 B.n370 585
R267 B.n372 B.n87 585
R268 B.n374 B.n373 585
R269 B.n375 B.n86 585
R270 B.n377 B.n376 585
R271 B.n378 B.n85 585
R272 B.n380 B.n379 585
R273 B.n381 B.n84 585
R274 B.n383 B.n382 585
R275 B.n384 B.n83 585
R276 B.n386 B.n385 585
R277 B.n387 B.n82 585
R278 B.n389 B.n388 585
R279 B.n390 B.n81 585
R280 B.n392 B.n391 585
R281 B.n393 B.n80 585
R282 B.n395 B.n394 585
R283 B.n396 B.n79 585
R284 B.n398 B.n397 585
R285 B.n399 B.n78 585
R286 B.n401 B.n400 585
R287 B.n402 B.n77 585
R288 B.n404 B.n403 585
R289 B.n405 B.n76 585
R290 B.n407 B.n406 585
R291 B.n408 B.n75 585
R292 B.n410 B.n409 585
R293 B.n411 B.n74 585
R294 B.n413 B.n412 585
R295 B.n414 B.n73 585
R296 B.n416 B.n415 585
R297 B.n417 B.n72 585
R298 B.n419 B.n418 585
R299 B.n420 B.n71 585
R300 B.n422 B.n421 585
R301 B.n423 B.n70 585
R302 B.n425 B.n424 585
R303 B.n426 B.n69 585
R304 B.n428 B.n427 585
R305 B.n429 B.n68 585
R306 B.n431 B.n430 585
R307 B.n432 B.n67 585
R308 B.n434 B.n433 585
R309 B.n435 B.n66 585
R310 B.n437 B.n436 585
R311 B.n438 B.n65 585
R312 B.n440 B.n439 585
R313 B.n441 B.n64 585
R314 B.n443 B.n442 585
R315 B.n444 B.n63 585
R316 B.n446 B.n445 585
R317 B.n447 B.n62 585
R318 B.n449 B.n448 585
R319 B.n450 B.n61 585
R320 B.n554 B.n553 585
R321 B.n552 B.n23 585
R322 B.n551 B.n550 585
R323 B.n549 B.n24 585
R324 B.n548 B.n547 585
R325 B.n546 B.n25 585
R326 B.n545 B.n544 585
R327 B.n543 B.n26 585
R328 B.n542 B.n541 585
R329 B.n540 B.n27 585
R330 B.n539 B.n538 585
R331 B.n537 B.n28 585
R332 B.n536 B.n535 585
R333 B.n534 B.n29 585
R334 B.n533 B.n532 585
R335 B.n531 B.n30 585
R336 B.n530 B.n529 585
R337 B.n528 B.n31 585
R338 B.n527 B.n526 585
R339 B.n525 B.n32 585
R340 B.n524 B.n523 585
R341 B.n522 B.n33 585
R342 B.n521 B.n520 585
R343 B.n519 B.n34 585
R344 B.n518 B.n517 585
R345 B.n516 B.n35 585
R346 B.n515 B.n514 585
R347 B.n513 B.n36 585
R348 B.n512 B.n511 585
R349 B.n509 B.n37 585
R350 B.n508 B.n507 585
R351 B.n506 B.n40 585
R352 B.n505 B.n504 585
R353 B.n503 B.n41 585
R354 B.n502 B.n501 585
R355 B.n500 B.n42 585
R356 B.n499 B.n498 585
R357 B.n497 B.n43 585
R358 B.n496 B.n495 585
R359 B.n494 B.n493 585
R360 B.n492 B.n47 585
R361 B.n491 B.n490 585
R362 B.n489 B.n48 585
R363 B.n488 B.n487 585
R364 B.n486 B.n49 585
R365 B.n485 B.n484 585
R366 B.n483 B.n50 585
R367 B.n482 B.n481 585
R368 B.n480 B.n51 585
R369 B.n479 B.n478 585
R370 B.n477 B.n52 585
R371 B.n476 B.n475 585
R372 B.n474 B.n53 585
R373 B.n473 B.n472 585
R374 B.n471 B.n54 585
R375 B.n470 B.n469 585
R376 B.n468 B.n55 585
R377 B.n467 B.n466 585
R378 B.n465 B.n56 585
R379 B.n464 B.n463 585
R380 B.n462 B.n57 585
R381 B.n461 B.n460 585
R382 B.n459 B.n58 585
R383 B.n458 B.n457 585
R384 B.n456 B.n59 585
R385 B.n455 B.n454 585
R386 B.n453 B.n60 585
R387 B.n452 B.n451 585
R388 B.n555 B.n22 585
R389 B.n557 B.n556 585
R390 B.n558 B.n21 585
R391 B.n560 B.n559 585
R392 B.n561 B.n20 585
R393 B.n563 B.n562 585
R394 B.n564 B.n19 585
R395 B.n566 B.n565 585
R396 B.n567 B.n18 585
R397 B.n569 B.n568 585
R398 B.n570 B.n17 585
R399 B.n572 B.n571 585
R400 B.n573 B.n16 585
R401 B.n575 B.n574 585
R402 B.n576 B.n15 585
R403 B.n578 B.n577 585
R404 B.n579 B.n14 585
R405 B.n581 B.n580 585
R406 B.n582 B.n13 585
R407 B.n584 B.n583 585
R408 B.n585 B.n12 585
R409 B.n587 B.n586 585
R410 B.n588 B.n11 585
R411 B.n590 B.n589 585
R412 B.n591 B.n10 585
R413 B.n593 B.n592 585
R414 B.n594 B.n9 585
R415 B.n596 B.n595 585
R416 B.n597 B.n8 585
R417 B.n599 B.n598 585
R418 B.n600 B.n7 585
R419 B.n602 B.n601 585
R420 B.n603 B.n6 585
R421 B.n605 B.n604 585
R422 B.n606 B.n5 585
R423 B.n608 B.n607 585
R424 B.n609 B.n4 585
R425 B.n611 B.n610 585
R426 B.n612 B.n3 585
R427 B.n614 B.n613 585
R428 B.n615 B.n0 585
R429 B.n2 B.n1 585
R430 B.n160 B.n159 585
R431 B.n161 B.n158 585
R432 B.n163 B.n162 585
R433 B.n164 B.n157 585
R434 B.n166 B.n165 585
R435 B.n167 B.n156 585
R436 B.n169 B.n168 585
R437 B.n170 B.n155 585
R438 B.n172 B.n171 585
R439 B.n173 B.n154 585
R440 B.n175 B.n174 585
R441 B.n176 B.n153 585
R442 B.n178 B.n177 585
R443 B.n179 B.n152 585
R444 B.n181 B.n180 585
R445 B.n182 B.n151 585
R446 B.n184 B.n183 585
R447 B.n185 B.n150 585
R448 B.n187 B.n186 585
R449 B.n188 B.n149 585
R450 B.n190 B.n189 585
R451 B.n191 B.n148 585
R452 B.n193 B.n192 585
R453 B.n194 B.n147 585
R454 B.n196 B.n195 585
R455 B.n197 B.n146 585
R456 B.n199 B.n198 585
R457 B.n200 B.n145 585
R458 B.n202 B.n201 585
R459 B.n203 B.n144 585
R460 B.n205 B.n204 585
R461 B.n206 B.n143 585
R462 B.n208 B.n207 585
R463 B.n209 B.n142 585
R464 B.n211 B.n210 585
R465 B.n212 B.n141 585
R466 B.n214 B.n213 585
R467 B.n215 B.n140 585
R468 B.n217 B.n216 585
R469 B.n218 B.n139 585
R470 B.n220 B.n139 473.281
R471 B.n326 B.n103 473.281
R472 B.n452 B.n61 473.281
R473 B.n555 B.n554 473.281
R474 B.n261 B.t0 282.697
R475 B.n118 B.t9 282.697
R476 B.n44 B.t6 282.697
R477 B.n38 B.t3 282.697
R478 B.n617 B.n616 256.663
R479 B.n616 B.n615 235.042
R480 B.n616 B.n2 235.042
R481 B.n118 B.t10 169.212
R482 B.n44 B.t8 169.212
R483 B.n261 B.t1 169.202
R484 B.n38 B.t5 169.202
R485 B.n221 B.n220 163.367
R486 B.n222 B.n221 163.367
R487 B.n222 B.n137 163.367
R488 B.n226 B.n137 163.367
R489 B.n227 B.n226 163.367
R490 B.n228 B.n227 163.367
R491 B.n228 B.n135 163.367
R492 B.n232 B.n135 163.367
R493 B.n233 B.n232 163.367
R494 B.n234 B.n233 163.367
R495 B.n234 B.n133 163.367
R496 B.n238 B.n133 163.367
R497 B.n239 B.n238 163.367
R498 B.n240 B.n239 163.367
R499 B.n240 B.n131 163.367
R500 B.n244 B.n131 163.367
R501 B.n245 B.n244 163.367
R502 B.n246 B.n245 163.367
R503 B.n246 B.n129 163.367
R504 B.n250 B.n129 163.367
R505 B.n251 B.n250 163.367
R506 B.n252 B.n251 163.367
R507 B.n252 B.n127 163.367
R508 B.n256 B.n127 163.367
R509 B.n257 B.n256 163.367
R510 B.n258 B.n257 163.367
R511 B.n258 B.n125 163.367
R512 B.n265 B.n125 163.367
R513 B.n266 B.n265 163.367
R514 B.n267 B.n266 163.367
R515 B.n267 B.n123 163.367
R516 B.n271 B.n123 163.367
R517 B.n272 B.n271 163.367
R518 B.n273 B.n272 163.367
R519 B.n273 B.n121 163.367
R520 B.n277 B.n121 163.367
R521 B.n278 B.n277 163.367
R522 B.n279 B.n278 163.367
R523 B.n279 B.n117 163.367
R524 B.n284 B.n117 163.367
R525 B.n285 B.n284 163.367
R526 B.n286 B.n285 163.367
R527 B.n286 B.n115 163.367
R528 B.n290 B.n115 163.367
R529 B.n291 B.n290 163.367
R530 B.n292 B.n291 163.367
R531 B.n292 B.n113 163.367
R532 B.n296 B.n113 163.367
R533 B.n297 B.n296 163.367
R534 B.n298 B.n297 163.367
R535 B.n298 B.n111 163.367
R536 B.n302 B.n111 163.367
R537 B.n303 B.n302 163.367
R538 B.n304 B.n303 163.367
R539 B.n304 B.n109 163.367
R540 B.n308 B.n109 163.367
R541 B.n309 B.n308 163.367
R542 B.n310 B.n309 163.367
R543 B.n310 B.n107 163.367
R544 B.n314 B.n107 163.367
R545 B.n315 B.n314 163.367
R546 B.n316 B.n315 163.367
R547 B.n316 B.n105 163.367
R548 B.n320 B.n105 163.367
R549 B.n321 B.n320 163.367
R550 B.n322 B.n321 163.367
R551 B.n322 B.n103 163.367
R552 B.n448 B.n61 163.367
R553 B.n448 B.n447 163.367
R554 B.n447 B.n446 163.367
R555 B.n446 B.n63 163.367
R556 B.n442 B.n63 163.367
R557 B.n442 B.n441 163.367
R558 B.n441 B.n440 163.367
R559 B.n440 B.n65 163.367
R560 B.n436 B.n65 163.367
R561 B.n436 B.n435 163.367
R562 B.n435 B.n434 163.367
R563 B.n434 B.n67 163.367
R564 B.n430 B.n67 163.367
R565 B.n430 B.n429 163.367
R566 B.n429 B.n428 163.367
R567 B.n428 B.n69 163.367
R568 B.n424 B.n69 163.367
R569 B.n424 B.n423 163.367
R570 B.n423 B.n422 163.367
R571 B.n422 B.n71 163.367
R572 B.n418 B.n71 163.367
R573 B.n418 B.n417 163.367
R574 B.n417 B.n416 163.367
R575 B.n416 B.n73 163.367
R576 B.n412 B.n73 163.367
R577 B.n412 B.n411 163.367
R578 B.n411 B.n410 163.367
R579 B.n410 B.n75 163.367
R580 B.n406 B.n75 163.367
R581 B.n406 B.n405 163.367
R582 B.n405 B.n404 163.367
R583 B.n404 B.n77 163.367
R584 B.n400 B.n77 163.367
R585 B.n400 B.n399 163.367
R586 B.n399 B.n398 163.367
R587 B.n398 B.n79 163.367
R588 B.n394 B.n79 163.367
R589 B.n394 B.n393 163.367
R590 B.n393 B.n392 163.367
R591 B.n392 B.n81 163.367
R592 B.n388 B.n81 163.367
R593 B.n388 B.n387 163.367
R594 B.n387 B.n386 163.367
R595 B.n386 B.n83 163.367
R596 B.n382 B.n83 163.367
R597 B.n382 B.n381 163.367
R598 B.n381 B.n380 163.367
R599 B.n380 B.n85 163.367
R600 B.n376 B.n85 163.367
R601 B.n376 B.n375 163.367
R602 B.n375 B.n374 163.367
R603 B.n374 B.n87 163.367
R604 B.n370 B.n87 163.367
R605 B.n370 B.n369 163.367
R606 B.n369 B.n368 163.367
R607 B.n368 B.n89 163.367
R608 B.n364 B.n89 163.367
R609 B.n364 B.n363 163.367
R610 B.n363 B.n362 163.367
R611 B.n362 B.n91 163.367
R612 B.n358 B.n91 163.367
R613 B.n358 B.n357 163.367
R614 B.n357 B.n356 163.367
R615 B.n356 B.n93 163.367
R616 B.n352 B.n93 163.367
R617 B.n352 B.n351 163.367
R618 B.n351 B.n350 163.367
R619 B.n350 B.n95 163.367
R620 B.n346 B.n95 163.367
R621 B.n346 B.n345 163.367
R622 B.n345 B.n344 163.367
R623 B.n344 B.n97 163.367
R624 B.n340 B.n97 163.367
R625 B.n340 B.n339 163.367
R626 B.n339 B.n338 163.367
R627 B.n338 B.n99 163.367
R628 B.n334 B.n99 163.367
R629 B.n334 B.n333 163.367
R630 B.n333 B.n332 163.367
R631 B.n332 B.n101 163.367
R632 B.n328 B.n101 163.367
R633 B.n328 B.n327 163.367
R634 B.n327 B.n326 163.367
R635 B.n554 B.n23 163.367
R636 B.n550 B.n23 163.367
R637 B.n550 B.n549 163.367
R638 B.n549 B.n548 163.367
R639 B.n548 B.n25 163.367
R640 B.n544 B.n25 163.367
R641 B.n544 B.n543 163.367
R642 B.n543 B.n542 163.367
R643 B.n542 B.n27 163.367
R644 B.n538 B.n27 163.367
R645 B.n538 B.n537 163.367
R646 B.n537 B.n536 163.367
R647 B.n536 B.n29 163.367
R648 B.n532 B.n29 163.367
R649 B.n532 B.n531 163.367
R650 B.n531 B.n530 163.367
R651 B.n530 B.n31 163.367
R652 B.n526 B.n31 163.367
R653 B.n526 B.n525 163.367
R654 B.n525 B.n524 163.367
R655 B.n524 B.n33 163.367
R656 B.n520 B.n33 163.367
R657 B.n520 B.n519 163.367
R658 B.n519 B.n518 163.367
R659 B.n518 B.n35 163.367
R660 B.n514 B.n35 163.367
R661 B.n514 B.n513 163.367
R662 B.n513 B.n512 163.367
R663 B.n512 B.n37 163.367
R664 B.n507 B.n37 163.367
R665 B.n507 B.n506 163.367
R666 B.n506 B.n505 163.367
R667 B.n505 B.n41 163.367
R668 B.n501 B.n41 163.367
R669 B.n501 B.n500 163.367
R670 B.n500 B.n499 163.367
R671 B.n499 B.n43 163.367
R672 B.n495 B.n43 163.367
R673 B.n495 B.n494 163.367
R674 B.n494 B.n47 163.367
R675 B.n490 B.n47 163.367
R676 B.n490 B.n489 163.367
R677 B.n489 B.n488 163.367
R678 B.n488 B.n49 163.367
R679 B.n484 B.n49 163.367
R680 B.n484 B.n483 163.367
R681 B.n483 B.n482 163.367
R682 B.n482 B.n51 163.367
R683 B.n478 B.n51 163.367
R684 B.n478 B.n477 163.367
R685 B.n477 B.n476 163.367
R686 B.n476 B.n53 163.367
R687 B.n472 B.n53 163.367
R688 B.n472 B.n471 163.367
R689 B.n471 B.n470 163.367
R690 B.n470 B.n55 163.367
R691 B.n466 B.n55 163.367
R692 B.n466 B.n465 163.367
R693 B.n465 B.n464 163.367
R694 B.n464 B.n57 163.367
R695 B.n460 B.n57 163.367
R696 B.n460 B.n459 163.367
R697 B.n459 B.n458 163.367
R698 B.n458 B.n59 163.367
R699 B.n454 B.n59 163.367
R700 B.n454 B.n453 163.367
R701 B.n453 B.n452 163.367
R702 B.n556 B.n555 163.367
R703 B.n556 B.n21 163.367
R704 B.n560 B.n21 163.367
R705 B.n561 B.n560 163.367
R706 B.n562 B.n561 163.367
R707 B.n562 B.n19 163.367
R708 B.n566 B.n19 163.367
R709 B.n567 B.n566 163.367
R710 B.n568 B.n567 163.367
R711 B.n568 B.n17 163.367
R712 B.n572 B.n17 163.367
R713 B.n573 B.n572 163.367
R714 B.n574 B.n573 163.367
R715 B.n574 B.n15 163.367
R716 B.n578 B.n15 163.367
R717 B.n579 B.n578 163.367
R718 B.n580 B.n579 163.367
R719 B.n580 B.n13 163.367
R720 B.n584 B.n13 163.367
R721 B.n585 B.n584 163.367
R722 B.n586 B.n585 163.367
R723 B.n586 B.n11 163.367
R724 B.n590 B.n11 163.367
R725 B.n591 B.n590 163.367
R726 B.n592 B.n591 163.367
R727 B.n592 B.n9 163.367
R728 B.n596 B.n9 163.367
R729 B.n597 B.n596 163.367
R730 B.n598 B.n597 163.367
R731 B.n598 B.n7 163.367
R732 B.n602 B.n7 163.367
R733 B.n603 B.n602 163.367
R734 B.n604 B.n603 163.367
R735 B.n604 B.n5 163.367
R736 B.n608 B.n5 163.367
R737 B.n609 B.n608 163.367
R738 B.n610 B.n609 163.367
R739 B.n610 B.n3 163.367
R740 B.n614 B.n3 163.367
R741 B.n615 B.n614 163.367
R742 B.n160 B.n2 163.367
R743 B.n161 B.n160 163.367
R744 B.n162 B.n161 163.367
R745 B.n162 B.n157 163.367
R746 B.n166 B.n157 163.367
R747 B.n167 B.n166 163.367
R748 B.n168 B.n167 163.367
R749 B.n168 B.n155 163.367
R750 B.n172 B.n155 163.367
R751 B.n173 B.n172 163.367
R752 B.n174 B.n173 163.367
R753 B.n174 B.n153 163.367
R754 B.n178 B.n153 163.367
R755 B.n179 B.n178 163.367
R756 B.n180 B.n179 163.367
R757 B.n180 B.n151 163.367
R758 B.n184 B.n151 163.367
R759 B.n185 B.n184 163.367
R760 B.n186 B.n185 163.367
R761 B.n186 B.n149 163.367
R762 B.n190 B.n149 163.367
R763 B.n191 B.n190 163.367
R764 B.n192 B.n191 163.367
R765 B.n192 B.n147 163.367
R766 B.n196 B.n147 163.367
R767 B.n197 B.n196 163.367
R768 B.n198 B.n197 163.367
R769 B.n198 B.n145 163.367
R770 B.n202 B.n145 163.367
R771 B.n203 B.n202 163.367
R772 B.n204 B.n203 163.367
R773 B.n204 B.n143 163.367
R774 B.n208 B.n143 163.367
R775 B.n209 B.n208 163.367
R776 B.n210 B.n209 163.367
R777 B.n210 B.n141 163.367
R778 B.n214 B.n141 163.367
R779 B.n215 B.n214 163.367
R780 B.n216 B.n215 163.367
R781 B.n216 B.n139 163.367
R782 B.n119 B.t11 114.326
R783 B.n45 B.t7 114.326
R784 B.n262 B.t2 114.319
R785 B.n39 B.t4 114.319
R786 B.n263 B.n262 59.5399
R787 B.n281 B.n119 59.5399
R788 B.n46 B.n45 59.5399
R789 B.n510 B.n39 59.5399
R790 B.n262 B.n261 54.8853
R791 B.n119 B.n118 54.8853
R792 B.n45 B.n44 54.8853
R793 B.n39 B.n38 54.8853
R794 B.n553 B.n22 30.7517
R795 B.n451 B.n450 30.7517
R796 B.n325 B.n324 30.7517
R797 B.n219 B.n218 30.7517
R798 B B.n617 18.0485
R799 B.n557 B.n22 10.6151
R800 B.n558 B.n557 10.6151
R801 B.n559 B.n558 10.6151
R802 B.n559 B.n20 10.6151
R803 B.n563 B.n20 10.6151
R804 B.n564 B.n563 10.6151
R805 B.n565 B.n564 10.6151
R806 B.n565 B.n18 10.6151
R807 B.n569 B.n18 10.6151
R808 B.n570 B.n569 10.6151
R809 B.n571 B.n570 10.6151
R810 B.n571 B.n16 10.6151
R811 B.n575 B.n16 10.6151
R812 B.n576 B.n575 10.6151
R813 B.n577 B.n576 10.6151
R814 B.n577 B.n14 10.6151
R815 B.n581 B.n14 10.6151
R816 B.n582 B.n581 10.6151
R817 B.n583 B.n582 10.6151
R818 B.n583 B.n12 10.6151
R819 B.n587 B.n12 10.6151
R820 B.n588 B.n587 10.6151
R821 B.n589 B.n588 10.6151
R822 B.n589 B.n10 10.6151
R823 B.n593 B.n10 10.6151
R824 B.n594 B.n593 10.6151
R825 B.n595 B.n594 10.6151
R826 B.n595 B.n8 10.6151
R827 B.n599 B.n8 10.6151
R828 B.n600 B.n599 10.6151
R829 B.n601 B.n600 10.6151
R830 B.n601 B.n6 10.6151
R831 B.n605 B.n6 10.6151
R832 B.n606 B.n605 10.6151
R833 B.n607 B.n606 10.6151
R834 B.n607 B.n4 10.6151
R835 B.n611 B.n4 10.6151
R836 B.n612 B.n611 10.6151
R837 B.n613 B.n612 10.6151
R838 B.n613 B.n0 10.6151
R839 B.n553 B.n552 10.6151
R840 B.n552 B.n551 10.6151
R841 B.n551 B.n24 10.6151
R842 B.n547 B.n24 10.6151
R843 B.n547 B.n546 10.6151
R844 B.n546 B.n545 10.6151
R845 B.n545 B.n26 10.6151
R846 B.n541 B.n26 10.6151
R847 B.n541 B.n540 10.6151
R848 B.n540 B.n539 10.6151
R849 B.n539 B.n28 10.6151
R850 B.n535 B.n28 10.6151
R851 B.n535 B.n534 10.6151
R852 B.n534 B.n533 10.6151
R853 B.n533 B.n30 10.6151
R854 B.n529 B.n30 10.6151
R855 B.n529 B.n528 10.6151
R856 B.n528 B.n527 10.6151
R857 B.n527 B.n32 10.6151
R858 B.n523 B.n32 10.6151
R859 B.n523 B.n522 10.6151
R860 B.n522 B.n521 10.6151
R861 B.n521 B.n34 10.6151
R862 B.n517 B.n34 10.6151
R863 B.n517 B.n516 10.6151
R864 B.n516 B.n515 10.6151
R865 B.n515 B.n36 10.6151
R866 B.n511 B.n36 10.6151
R867 B.n509 B.n508 10.6151
R868 B.n508 B.n40 10.6151
R869 B.n504 B.n40 10.6151
R870 B.n504 B.n503 10.6151
R871 B.n503 B.n502 10.6151
R872 B.n502 B.n42 10.6151
R873 B.n498 B.n42 10.6151
R874 B.n498 B.n497 10.6151
R875 B.n497 B.n496 10.6151
R876 B.n493 B.n492 10.6151
R877 B.n492 B.n491 10.6151
R878 B.n491 B.n48 10.6151
R879 B.n487 B.n48 10.6151
R880 B.n487 B.n486 10.6151
R881 B.n486 B.n485 10.6151
R882 B.n485 B.n50 10.6151
R883 B.n481 B.n50 10.6151
R884 B.n481 B.n480 10.6151
R885 B.n480 B.n479 10.6151
R886 B.n479 B.n52 10.6151
R887 B.n475 B.n52 10.6151
R888 B.n475 B.n474 10.6151
R889 B.n474 B.n473 10.6151
R890 B.n473 B.n54 10.6151
R891 B.n469 B.n54 10.6151
R892 B.n469 B.n468 10.6151
R893 B.n468 B.n467 10.6151
R894 B.n467 B.n56 10.6151
R895 B.n463 B.n56 10.6151
R896 B.n463 B.n462 10.6151
R897 B.n462 B.n461 10.6151
R898 B.n461 B.n58 10.6151
R899 B.n457 B.n58 10.6151
R900 B.n457 B.n456 10.6151
R901 B.n456 B.n455 10.6151
R902 B.n455 B.n60 10.6151
R903 B.n451 B.n60 10.6151
R904 B.n450 B.n449 10.6151
R905 B.n449 B.n62 10.6151
R906 B.n445 B.n62 10.6151
R907 B.n445 B.n444 10.6151
R908 B.n444 B.n443 10.6151
R909 B.n443 B.n64 10.6151
R910 B.n439 B.n64 10.6151
R911 B.n439 B.n438 10.6151
R912 B.n438 B.n437 10.6151
R913 B.n437 B.n66 10.6151
R914 B.n433 B.n66 10.6151
R915 B.n433 B.n432 10.6151
R916 B.n432 B.n431 10.6151
R917 B.n431 B.n68 10.6151
R918 B.n427 B.n68 10.6151
R919 B.n427 B.n426 10.6151
R920 B.n426 B.n425 10.6151
R921 B.n425 B.n70 10.6151
R922 B.n421 B.n70 10.6151
R923 B.n421 B.n420 10.6151
R924 B.n420 B.n419 10.6151
R925 B.n419 B.n72 10.6151
R926 B.n415 B.n72 10.6151
R927 B.n415 B.n414 10.6151
R928 B.n414 B.n413 10.6151
R929 B.n413 B.n74 10.6151
R930 B.n409 B.n74 10.6151
R931 B.n409 B.n408 10.6151
R932 B.n408 B.n407 10.6151
R933 B.n407 B.n76 10.6151
R934 B.n403 B.n76 10.6151
R935 B.n403 B.n402 10.6151
R936 B.n402 B.n401 10.6151
R937 B.n401 B.n78 10.6151
R938 B.n397 B.n78 10.6151
R939 B.n397 B.n396 10.6151
R940 B.n396 B.n395 10.6151
R941 B.n395 B.n80 10.6151
R942 B.n391 B.n80 10.6151
R943 B.n391 B.n390 10.6151
R944 B.n390 B.n389 10.6151
R945 B.n389 B.n82 10.6151
R946 B.n385 B.n82 10.6151
R947 B.n385 B.n384 10.6151
R948 B.n384 B.n383 10.6151
R949 B.n383 B.n84 10.6151
R950 B.n379 B.n84 10.6151
R951 B.n379 B.n378 10.6151
R952 B.n378 B.n377 10.6151
R953 B.n377 B.n86 10.6151
R954 B.n373 B.n86 10.6151
R955 B.n373 B.n372 10.6151
R956 B.n372 B.n371 10.6151
R957 B.n371 B.n88 10.6151
R958 B.n367 B.n88 10.6151
R959 B.n367 B.n366 10.6151
R960 B.n366 B.n365 10.6151
R961 B.n365 B.n90 10.6151
R962 B.n361 B.n90 10.6151
R963 B.n361 B.n360 10.6151
R964 B.n360 B.n359 10.6151
R965 B.n359 B.n92 10.6151
R966 B.n355 B.n92 10.6151
R967 B.n355 B.n354 10.6151
R968 B.n354 B.n353 10.6151
R969 B.n353 B.n94 10.6151
R970 B.n349 B.n94 10.6151
R971 B.n349 B.n348 10.6151
R972 B.n348 B.n347 10.6151
R973 B.n347 B.n96 10.6151
R974 B.n343 B.n96 10.6151
R975 B.n343 B.n342 10.6151
R976 B.n342 B.n341 10.6151
R977 B.n341 B.n98 10.6151
R978 B.n337 B.n98 10.6151
R979 B.n337 B.n336 10.6151
R980 B.n336 B.n335 10.6151
R981 B.n335 B.n100 10.6151
R982 B.n331 B.n100 10.6151
R983 B.n331 B.n330 10.6151
R984 B.n330 B.n329 10.6151
R985 B.n329 B.n102 10.6151
R986 B.n325 B.n102 10.6151
R987 B.n159 B.n1 10.6151
R988 B.n159 B.n158 10.6151
R989 B.n163 B.n158 10.6151
R990 B.n164 B.n163 10.6151
R991 B.n165 B.n164 10.6151
R992 B.n165 B.n156 10.6151
R993 B.n169 B.n156 10.6151
R994 B.n170 B.n169 10.6151
R995 B.n171 B.n170 10.6151
R996 B.n171 B.n154 10.6151
R997 B.n175 B.n154 10.6151
R998 B.n176 B.n175 10.6151
R999 B.n177 B.n176 10.6151
R1000 B.n177 B.n152 10.6151
R1001 B.n181 B.n152 10.6151
R1002 B.n182 B.n181 10.6151
R1003 B.n183 B.n182 10.6151
R1004 B.n183 B.n150 10.6151
R1005 B.n187 B.n150 10.6151
R1006 B.n188 B.n187 10.6151
R1007 B.n189 B.n188 10.6151
R1008 B.n189 B.n148 10.6151
R1009 B.n193 B.n148 10.6151
R1010 B.n194 B.n193 10.6151
R1011 B.n195 B.n194 10.6151
R1012 B.n195 B.n146 10.6151
R1013 B.n199 B.n146 10.6151
R1014 B.n200 B.n199 10.6151
R1015 B.n201 B.n200 10.6151
R1016 B.n201 B.n144 10.6151
R1017 B.n205 B.n144 10.6151
R1018 B.n206 B.n205 10.6151
R1019 B.n207 B.n206 10.6151
R1020 B.n207 B.n142 10.6151
R1021 B.n211 B.n142 10.6151
R1022 B.n212 B.n211 10.6151
R1023 B.n213 B.n212 10.6151
R1024 B.n213 B.n140 10.6151
R1025 B.n217 B.n140 10.6151
R1026 B.n218 B.n217 10.6151
R1027 B.n219 B.n138 10.6151
R1028 B.n223 B.n138 10.6151
R1029 B.n224 B.n223 10.6151
R1030 B.n225 B.n224 10.6151
R1031 B.n225 B.n136 10.6151
R1032 B.n229 B.n136 10.6151
R1033 B.n230 B.n229 10.6151
R1034 B.n231 B.n230 10.6151
R1035 B.n231 B.n134 10.6151
R1036 B.n235 B.n134 10.6151
R1037 B.n236 B.n235 10.6151
R1038 B.n237 B.n236 10.6151
R1039 B.n237 B.n132 10.6151
R1040 B.n241 B.n132 10.6151
R1041 B.n242 B.n241 10.6151
R1042 B.n243 B.n242 10.6151
R1043 B.n243 B.n130 10.6151
R1044 B.n247 B.n130 10.6151
R1045 B.n248 B.n247 10.6151
R1046 B.n249 B.n248 10.6151
R1047 B.n249 B.n128 10.6151
R1048 B.n253 B.n128 10.6151
R1049 B.n254 B.n253 10.6151
R1050 B.n255 B.n254 10.6151
R1051 B.n255 B.n126 10.6151
R1052 B.n259 B.n126 10.6151
R1053 B.n260 B.n259 10.6151
R1054 B.n264 B.n260 10.6151
R1055 B.n268 B.n124 10.6151
R1056 B.n269 B.n268 10.6151
R1057 B.n270 B.n269 10.6151
R1058 B.n270 B.n122 10.6151
R1059 B.n274 B.n122 10.6151
R1060 B.n275 B.n274 10.6151
R1061 B.n276 B.n275 10.6151
R1062 B.n276 B.n120 10.6151
R1063 B.n280 B.n120 10.6151
R1064 B.n283 B.n282 10.6151
R1065 B.n283 B.n116 10.6151
R1066 B.n287 B.n116 10.6151
R1067 B.n288 B.n287 10.6151
R1068 B.n289 B.n288 10.6151
R1069 B.n289 B.n114 10.6151
R1070 B.n293 B.n114 10.6151
R1071 B.n294 B.n293 10.6151
R1072 B.n295 B.n294 10.6151
R1073 B.n295 B.n112 10.6151
R1074 B.n299 B.n112 10.6151
R1075 B.n300 B.n299 10.6151
R1076 B.n301 B.n300 10.6151
R1077 B.n301 B.n110 10.6151
R1078 B.n305 B.n110 10.6151
R1079 B.n306 B.n305 10.6151
R1080 B.n307 B.n306 10.6151
R1081 B.n307 B.n108 10.6151
R1082 B.n311 B.n108 10.6151
R1083 B.n312 B.n311 10.6151
R1084 B.n313 B.n312 10.6151
R1085 B.n313 B.n106 10.6151
R1086 B.n317 B.n106 10.6151
R1087 B.n318 B.n317 10.6151
R1088 B.n319 B.n318 10.6151
R1089 B.n319 B.n104 10.6151
R1090 B.n323 B.n104 10.6151
R1091 B.n324 B.n323 10.6151
R1092 B.n511 B.n510 9.36635
R1093 B.n493 B.n46 9.36635
R1094 B.n264 B.n263 9.36635
R1095 B.n282 B.n281 9.36635
R1096 B.n617 B.n0 8.11757
R1097 B.n617 B.n1 8.11757
R1098 B.n510 B.n509 1.24928
R1099 B.n496 B.n46 1.24928
R1100 B.n263 B.n124 1.24928
R1101 B.n281 B.n280 1.24928
C0 VDD1 B 1.73199f
C1 VDD2 w_n3234_n2520# 2.05533f
C2 VP VN 6.04395f
C3 w_n3234_n2520# VN 6.02464f
C4 VDD2 VTAIL 6.20524f
C5 VP w_n3234_n2520# 6.442471f
C6 VDD2 VDD1 1.36802f
C7 VDD2 B 1.80368f
C8 VTAIL VN 4.76797f
C9 VTAIL VP 4.7822f
C10 VDD1 VN 0.151007f
C11 VN B 1.09994f
C12 VDD1 VP 4.74321f
C13 VP B 1.79705f
C14 VTAIL w_n3234_n2520# 2.37655f
C15 VDD1 w_n3234_n2520# 1.97347f
C16 w_n3234_n2520# B 8.34928f
C17 VDD2 VN 4.44677f
C18 VDD2 VP 0.449902f
C19 VDD1 VTAIL 6.15416f
C20 VTAIL B 2.70981f
C21 VDD2 VSUBS 1.651466f
C22 VDD1 VSUBS 1.980438f
C23 VTAIL VSUBS 1.024154f
C24 VN VSUBS 5.59911f
C25 VP VSUBS 2.697385f
C26 B VSUBS 4.180428f
C27 w_n3234_n2520# VSUBS 0.101172p
C28 B.n0 VSUBS 0.00623f
C29 B.n1 VSUBS 0.00623f
C30 B.n2 VSUBS 0.009214f
C31 B.n3 VSUBS 0.007061f
C32 B.n4 VSUBS 0.007061f
C33 B.n5 VSUBS 0.007061f
C34 B.n6 VSUBS 0.007061f
C35 B.n7 VSUBS 0.007061f
C36 B.n8 VSUBS 0.007061f
C37 B.n9 VSUBS 0.007061f
C38 B.n10 VSUBS 0.007061f
C39 B.n11 VSUBS 0.007061f
C40 B.n12 VSUBS 0.007061f
C41 B.n13 VSUBS 0.007061f
C42 B.n14 VSUBS 0.007061f
C43 B.n15 VSUBS 0.007061f
C44 B.n16 VSUBS 0.007061f
C45 B.n17 VSUBS 0.007061f
C46 B.n18 VSUBS 0.007061f
C47 B.n19 VSUBS 0.007061f
C48 B.n20 VSUBS 0.007061f
C49 B.n21 VSUBS 0.007061f
C50 B.n22 VSUBS 0.015487f
C51 B.n23 VSUBS 0.007061f
C52 B.n24 VSUBS 0.007061f
C53 B.n25 VSUBS 0.007061f
C54 B.n26 VSUBS 0.007061f
C55 B.n27 VSUBS 0.007061f
C56 B.n28 VSUBS 0.007061f
C57 B.n29 VSUBS 0.007061f
C58 B.n30 VSUBS 0.007061f
C59 B.n31 VSUBS 0.007061f
C60 B.n32 VSUBS 0.007061f
C61 B.n33 VSUBS 0.007061f
C62 B.n34 VSUBS 0.007061f
C63 B.n35 VSUBS 0.007061f
C64 B.n36 VSUBS 0.007061f
C65 B.n37 VSUBS 0.007061f
C66 B.t4 VSUBS 0.240214f
C67 B.t5 VSUBS 0.260181f
C68 B.t3 VSUBS 0.911811f
C69 B.n38 VSUBS 0.141603f
C70 B.n39 VSUBS 0.071626f
C71 B.n40 VSUBS 0.007061f
C72 B.n41 VSUBS 0.007061f
C73 B.n42 VSUBS 0.007061f
C74 B.n43 VSUBS 0.007061f
C75 B.t7 VSUBS 0.240212f
C76 B.t8 VSUBS 0.260178f
C77 B.t6 VSUBS 0.911811f
C78 B.n44 VSUBS 0.141606f
C79 B.n45 VSUBS 0.071628f
C80 B.n46 VSUBS 0.01636f
C81 B.n47 VSUBS 0.007061f
C82 B.n48 VSUBS 0.007061f
C83 B.n49 VSUBS 0.007061f
C84 B.n50 VSUBS 0.007061f
C85 B.n51 VSUBS 0.007061f
C86 B.n52 VSUBS 0.007061f
C87 B.n53 VSUBS 0.007061f
C88 B.n54 VSUBS 0.007061f
C89 B.n55 VSUBS 0.007061f
C90 B.n56 VSUBS 0.007061f
C91 B.n57 VSUBS 0.007061f
C92 B.n58 VSUBS 0.007061f
C93 B.n59 VSUBS 0.007061f
C94 B.n60 VSUBS 0.007061f
C95 B.n61 VSUBS 0.015487f
C96 B.n62 VSUBS 0.007061f
C97 B.n63 VSUBS 0.007061f
C98 B.n64 VSUBS 0.007061f
C99 B.n65 VSUBS 0.007061f
C100 B.n66 VSUBS 0.007061f
C101 B.n67 VSUBS 0.007061f
C102 B.n68 VSUBS 0.007061f
C103 B.n69 VSUBS 0.007061f
C104 B.n70 VSUBS 0.007061f
C105 B.n71 VSUBS 0.007061f
C106 B.n72 VSUBS 0.007061f
C107 B.n73 VSUBS 0.007061f
C108 B.n74 VSUBS 0.007061f
C109 B.n75 VSUBS 0.007061f
C110 B.n76 VSUBS 0.007061f
C111 B.n77 VSUBS 0.007061f
C112 B.n78 VSUBS 0.007061f
C113 B.n79 VSUBS 0.007061f
C114 B.n80 VSUBS 0.007061f
C115 B.n81 VSUBS 0.007061f
C116 B.n82 VSUBS 0.007061f
C117 B.n83 VSUBS 0.007061f
C118 B.n84 VSUBS 0.007061f
C119 B.n85 VSUBS 0.007061f
C120 B.n86 VSUBS 0.007061f
C121 B.n87 VSUBS 0.007061f
C122 B.n88 VSUBS 0.007061f
C123 B.n89 VSUBS 0.007061f
C124 B.n90 VSUBS 0.007061f
C125 B.n91 VSUBS 0.007061f
C126 B.n92 VSUBS 0.007061f
C127 B.n93 VSUBS 0.007061f
C128 B.n94 VSUBS 0.007061f
C129 B.n95 VSUBS 0.007061f
C130 B.n96 VSUBS 0.007061f
C131 B.n97 VSUBS 0.007061f
C132 B.n98 VSUBS 0.007061f
C133 B.n99 VSUBS 0.007061f
C134 B.n100 VSUBS 0.007061f
C135 B.n101 VSUBS 0.007061f
C136 B.n102 VSUBS 0.007061f
C137 B.n103 VSUBS 0.016287f
C138 B.n104 VSUBS 0.007061f
C139 B.n105 VSUBS 0.007061f
C140 B.n106 VSUBS 0.007061f
C141 B.n107 VSUBS 0.007061f
C142 B.n108 VSUBS 0.007061f
C143 B.n109 VSUBS 0.007061f
C144 B.n110 VSUBS 0.007061f
C145 B.n111 VSUBS 0.007061f
C146 B.n112 VSUBS 0.007061f
C147 B.n113 VSUBS 0.007061f
C148 B.n114 VSUBS 0.007061f
C149 B.n115 VSUBS 0.007061f
C150 B.n116 VSUBS 0.007061f
C151 B.n117 VSUBS 0.007061f
C152 B.t11 VSUBS 0.240212f
C153 B.t10 VSUBS 0.260178f
C154 B.t9 VSUBS 0.911811f
C155 B.n118 VSUBS 0.141606f
C156 B.n119 VSUBS 0.071628f
C157 B.n120 VSUBS 0.007061f
C158 B.n121 VSUBS 0.007061f
C159 B.n122 VSUBS 0.007061f
C160 B.n123 VSUBS 0.007061f
C161 B.n124 VSUBS 0.003946f
C162 B.n125 VSUBS 0.007061f
C163 B.n126 VSUBS 0.007061f
C164 B.n127 VSUBS 0.007061f
C165 B.n128 VSUBS 0.007061f
C166 B.n129 VSUBS 0.007061f
C167 B.n130 VSUBS 0.007061f
C168 B.n131 VSUBS 0.007061f
C169 B.n132 VSUBS 0.007061f
C170 B.n133 VSUBS 0.007061f
C171 B.n134 VSUBS 0.007061f
C172 B.n135 VSUBS 0.007061f
C173 B.n136 VSUBS 0.007061f
C174 B.n137 VSUBS 0.007061f
C175 B.n138 VSUBS 0.007061f
C176 B.n139 VSUBS 0.015487f
C177 B.n140 VSUBS 0.007061f
C178 B.n141 VSUBS 0.007061f
C179 B.n142 VSUBS 0.007061f
C180 B.n143 VSUBS 0.007061f
C181 B.n144 VSUBS 0.007061f
C182 B.n145 VSUBS 0.007061f
C183 B.n146 VSUBS 0.007061f
C184 B.n147 VSUBS 0.007061f
C185 B.n148 VSUBS 0.007061f
C186 B.n149 VSUBS 0.007061f
C187 B.n150 VSUBS 0.007061f
C188 B.n151 VSUBS 0.007061f
C189 B.n152 VSUBS 0.007061f
C190 B.n153 VSUBS 0.007061f
C191 B.n154 VSUBS 0.007061f
C192 B.n155 VSUBS 0.007061f
C193 B.n156 VSUBS 0.007061f
C194 B.n157 VSUBS 0.007061f
C195 B.n158 VSUBS 0.007061f
C196 B.n159 VSUBS 0.007061f
C197 B.n160 VSUBS 0.007061f
C198 B.n161 VSUBS 0.007061f
C199 B.n162 VSUBS 0.007061f
C200 B.n163 VSUBS 0.007061f
C201 B.n164 VSUBS 0.007061f
C202 B.n165 VSUBS 0.007061f
C203 B.n166 VSUBS 0.007061f
C204 B.n167 VSUBS 0.007061f
C205 B.n168 VSUBS 0.007061f
C206 B.n169 VSUBS 0.007061f
C207 B.n170 VSUBS 0.007061f
C208 B.n171 VSUBS 0.007061f
C209 B.n172 VSUBS 0.007061f
C210 B.n173 VSUBS 0.007061f
C211 B.n174 VSUBS 0.007061f
C212 B.n175 VSUBS 0.007061f
C213 B.n176 VSUBS 0.007061f
C214 B.n177 VSUBS 0.007061f
C215 B.n178 VSUBS 0.007061f
C216 B.n179 VSUBS 0.007061f
C217 B.n180 VSUBS 0.007061f
C218 B.n181 VSUBS 0.007061f
C219 B.n182 VSUBS 0.007061f
C220 B.n183 VSUBS 0.007061f
C221 B.n184 VSUBS 0.007061f
C222 B.n185 VSUBS 0.007061f
C223 B.n186 VSUBS 0.007061f
C224 B.n187 VSUBS 0.007061f
C225 B.n188 VSUBS 0.007061f
C226 B.n189 VSUBS 0.007061f
C227 B.n190 VSUBS 0.007061f
C228 B.n191 VSUBS 0.007061f
C229 B.n192 VSUBS 0.007061f
C230 B.n193 VSUBS 0.007061f
C231 B.n194 VSUBS 0.007061f
C232 B.n195 VSUBS 0.007061f
C233 B.n196 VSUBS 0.007061f
C234 B.n197 VSUBS 0.007061f
C235 B.n198 VSUBS 0.007061f
C236 B.n199 VSUBS 0.007061f
C237 B.n200 VSUBS 0.007061f
C238 B.n201 VSUBS 0.007061f
C239 B.n202 VSUBS 0.007061f
C240 B.n203 VSUBS 0.007061f
C241 B.n204 VSUBS 0.007061f
C242 B.n205 VSUBS 0.007061f
C243 B.n206 VSUBS 0.007061f
C244 B.n207 VSUBS 0.007061f
C245 B.n208 VSUBS 0.007061f
C246 B.n209 VSUBS 0.007061f
C247 B.n210 VSUBS 0.007061f
C248 B.n211 VSUBS 0.007061f
C249 B.n212 VSUBS 0.007061f
C250 B.n213 VSUBS 0.007061f
C251 B.n214 VSUBS 0.007061f
C252 B.n215 VSUBS 0.007061f
C253 B.n216 VSUBS 0.007061f
C254 B.n217 VSUBS 0.007061f
C255 B.n218 VSUBS 0.015487f
C256 B.n219 VSUBS 0.016287f
C257 B.n220 VSUBS 0.016287f
C258 B.n221 VSUBS 0.007061f
C259 B.n222 VSUBS 0.007061f
C260 B.n223 VSUBS 0.007061f
C261 B.n224 VSUBS 0.007061f
C262 B.n225 VSUBS 0.007061f
C263 B.n226 VSUBS 0.007061f
C264 B.n227 VSUBS 0.007061f
C265 B.n228 VSUBS 0.007061f
C266 B.n229 VSUBS 0.007061f
C267 B.n230 VSUBS 0.007061f
C268 B.n231 VSUBS 0.007061f
C269 B.n232 VSUBS 0.007061f
C270 B.n233 VSUBS 0.007061f
C271 B.n234 VSUBS 0.007061f
C272 B.n235 VSUBS 0.007061f
C273 B.n236 VSUBS 0.007061f
C274 B.n237 VSUBS 0.007061f
C275 B.n238 VSUBS 0.007061f
C276 B.n239 VSUBS 0.007061f
C277 B.n240 VSUBS 0.007061f
C278 B.n241 VSUBS 0.007061f
C279 B.n242 VSUBS 0.007061f
C280 B.n243 VSUBS 0.007061f
C281 B.n244 VSUBS 0.007061f
C282 B.n245 VSUBS 0.007061f
C283 B.n246 VSUBS 0.007061f
C284 B.n247 VSUBS 0.007061f
C285 B.n248 VSUBS 0.007061f
C286 B.n249 VSUBS 0.007061f
C287 B.n250 VSUBS 0.007061f
C288 B.n251 VSUBS 0.007061f
C289 B.n252 VSUBS 0.007061f
C290 B.n253 VSUBS 0.007061f
C291 B.n254 VSUBS 0.007061f
C292 B.n255 VSUBS 0.007061f
C293 B.n256 VSUBS 0.007061f
C294 B.n257 VSUBS 0.007061f
C295 B.n258 VSUBS 0.007061f
C296 B.n259 VSUBS 0.007061f
C297 B.n260 VSUBS 0.007061f
C298 B.t2 VSUBS 0.240214f
C299 B.t1 VSUBS 0.260181f
C300 B.t0 VSUBS 0.911811f
C301 B.n261 VSUBS 0.141603f
C302 B.n262 VSUBS 0.071626f
C303 B.n263 VSUBS 0.01636f
C304 B.n264 VSUBS 0.006646f
C305 B.n265 VSUBS 0.007061f
C306 B.n266 VSUBS 0.007061f
C307 B.n267 VSUBS 0.007061f
C308 B.n268 VSUBS 0.007061f
C309 B.n269 VSUBS 0.007061f
C310 B.n270 VSUBS 0.007061f
C311 B.n271 VSUBS 0.007061f
C312 B.n272 VSUBS 0.007061f
C313 B.n273 VSUBS 0.007061f
C314 B.n274 VSUBS 0.007061f
C315 B.n275 VSUBS 0.007061f
C316 B.n276 VSUBS 0.007061f
C317 B.n277 VSUBS 0.007061f
C318 B.n278 VSUBS 0.007061f
C319 B.n279 VSUBS 0.007061f
C320 B.n280 VSUBS 0.003946f
C321 B.n281 VSUBS 0.01636f
C322 B.n282 VSUBS 0.006646f
C323 B.n283 VSUBS 0.007061f
C324 B.n284 VSUBS 0.007061f
C325 B.n285 VSUBS 0.007061f
C326 B.n286 VSUBS 0.007061f
C327 B.n287 VSUBS 0.007061f
C328 B.n288 VSUBS 0.007061f
C329 B.n289 VSUBS 0.007061f
C330 B.n290 VSUBS 0.007061f
C331 B.n291 VSUBS 0.007061f
C332 B.n292 VSUBS 0.007061f
C333 B.n293 VSUBS 0.007061f
C334 B.n294 VSUBS 0.007061f
C335 B.n295 VSUBS 0.007061f
C336 B.n296 VSUBS 0.007061f
C337 B.n297 VSUBS 0.007061f
C338 B.n298 VSUBS 0.007061f
C339 B.n299 VSUBS 0.007061f
C340 B.n300 VSUBS 0.007061f
C341 B.n301 VSUBS 0.007061f
C342 B.n302 VSUBS 0.007061f
C343 B.n303 VSUBS 0.007061f
C344 B.n304 VSUBS 0.007061f
C345 B.n305 VSUBS 0.007061f
C346 B.n306 VSUBS 0.007061f
C347 B.n307 VSUBS 0.007061f
C348 B.n308 VSUBS 0.007061f
C349 B.n309 VSUBS 0.007061f
C350 B.n310 VSUBS 0.007061f
C351 B.n311 VSUBS 0.007061f
C352 B.n312 VSUBS 0.007061f
C353 B.n313 VSUBS 0.007061f
C354 B.n314 VSUBS 0.007061f
C355 B.n315 VSUBS 0.007061f
C356 B.n316 VSUBS 0.007061f
C357 B.n317 VSUBS 0.007061f
C358 B.n318 VSUBS 0.007061f
C359 B.n319 VSUBS 0.007061f
C360 B.n320 VSUBS 0.007061f
C361 B.n321 VSUBS 0.007061f
C362 B.n322 VSUBS 0.007061f
C363 B.n323 VSUBS 0.007061f
C364 B.n324 VSUBS 0.015401f
C365 B.n325 VSUBS 0.016373f
C366 B.n326 VSUBS 0.015487f
C367 B.n327 VSUBS 0.007061f
C368 B.n328 VSUBS 0.007061f
C369 B.n329 VSUBS 0.007061f
C370 B.n330 VSUBS 0.007061f
C371 B.n331 VSUBS 0.007061f
C372 B.n332 VSUBS 0.007061f
C373 B.n333 VSUBS 0.007061f
C374 B.n334 VSUBS 0.007061f
C375 B.n335 VSUBS 0.007061f
C376 B.n336 VSUBS 0.007061f
C377 B.n337 VSUBS 0.007061f
C378 B.n338 VSUBS 0.007061f
C379 B.n339 VSUBS 0.007061f
C380 B.n340 VSUBS 0.007061f
C381 B.n341 VSUBS 0.007061f
C382 B.n342 VSUBS 0.007061f
C383 B.n343 VSUBS 0.007061f
C384 B.n344 VSUBS 0.007061f
C385 B.n345 VSUBS 0.007061f
C386 B.n346 VSUBS 0.007061f
C387 B.n347 VSUBS 0.007061f
C388 B.n348 VSUBS 0.007061f
C389 B.n349 VSUBS 0.007061f
C390 B.n350 VSUBS 0.007061f
C391 B.n351 VSUBS 0.007061f
C392 B.n352 VSUBS 0.007061f
C393 B.n353 VSUBS 0.007061f
C394 B.n354 VSUBS 0.007061f
C395 B.n355 VSUBS 0.007061f
C396 B.n356 VSUBS 0.007061f
C397 B.n357 VSUBS 0.007061f
C398 B.n358 VSUBS 0.007061f
C399 B.n359 VSUBS 0.007061f
C400 B.n360 VSUBS 0.007061f
C401 B.n361 VSUBS 0.007061f
C402 B.n362 VSUBS 0.007061f
C403 B.n363 VSUBS 0.007061f
C404 B.n364 VSUBS 0.007061f
C405 B.n365 VSUBS 0.007061f
C406 B.n366 VSUBS 0.007061f
C407 B.n367 VSUBS 0.007061f
C408 B.n368 VSUBS 0.007061f
C409 B.n369 VSUBS 0.007061f
C410 B.n370 VSUBS 0.007061f
C411 B.n371 VSUBS 0.007061f
C412 B.n372 VSUBS 0.007061f
C413 B.n373 VSUBS 0.007061f
C414 B.n374 VSUBS 0.007061f
C415 B.n375 VSUBS 0.007061f
C416 B.n376 VSUBS 0.007061f
C417 B.n377 VSUBS 0.007061f
C418 B.n378 VSUBS 0.007061f
C419 B.n379 VSUBS 0.007061f
C420 B.n380 VSUBS 0.007061f
C421 B.n381 VSUBS 0.007061f
C422 B.n382 VSUBS 0.007061f
C423 B.n383 VSUBS 0.007061f
C424 B.n384 VSUBS 0.007061f
C425 B.n385 VSUBS 0.007061f
C426 B.n386 VSUBS 0.007061f
C427 B.n387 VSUBS 0.007061f
C428 B.n388 VSUBS 0.007061f
C429 B.n389 VSUBS 0.007061f
C430 B.n390 VSUBS 0.007061f
C431 B.n391 VSUBS 0.007061f
C432 B.n392 VSUBS 0.007061f
C433 B.n393 VSUBS 0.007061f
C434 B.n394 VSUBS 0.007061f
C435 B.n395 VSUBS 0.007061f
C436 B.n396 VSUBS 0.007061f
C437 B.n397 VSUBS 0.007061f
C438 B.n398 VSUBS 0.007061f
C439 B.n399 VSUBS 0.007061f
C440 B.n400 VSUBS 0.007061f
C441 B.n401 VSUBS 0.007061f
C442 B.n402 VSUBS 0.007061f
C443 B.n403 VSUBS 0.007061f
C444 B.n404 VSUBS 0.007061f
C445 B.n405 VSUBS 0.007061f
C446 B.n406 VSUBS 0.007061f
C447 B.n407 VSUBS 0.007061f
C448 B.n408 VSUBS 0.007061f
C449 B.n409 VSUBS 0.007061f
C450 B.n410 VSUBS 0.007061f
C451 B.n411 VSUBS 0.007061f
C452 B.n412 VSUBS 0.007061f
C453 B.n413 VSUBS 0.007061f
C454 B.n414 VSUBS 0.007061f
C455 B.n415 VSUBS 0.007061f
C456 B.n416 VSUBS 0.007061f
C457 B.n417 VSUBS 0.007061f
C458 B.n418 VSUBS 0.007061f
C459 B.n419 VSUBS 0.007061f
C460 B.n420 VSUBS 0.007061f
C461 B.n421 VSUBS 0.007061f
C462 B.n422 VSUBS 0.007061f
C463 B.n423 VSUBS 0.007061f
C464 B.n424 VSUBS 0.007061f
C465 B.n425 VSUBS 0.007061f
C466 B.n426 VSUBS 0.007061f
C467 B.n427 VSUBS 0.007061f
C468 B.n428 VSUBS 0.007061f
C469 B.n429 VSUBS 0.007061f
C470 B.n430 VSUBS 0.007061f
C471 B.n431 VSUBS 0.007061f
C472 B.n432 VSUBS 0.007061f
C473 B.n433 VSUBS 0.007061f
C474 B.n434 VSUBS 0.007061f
C475 B.n435 VSUBS 0.007061f
C476 B.n436 VSUBS 0.007061f
C477 B.n437 VSUBS 0.007061f
C478 B.n438 VSUBS 0.007061f
C479 B.n439 VSUBS 0.007061f
C480 B.n440 VSUBS 0.007061f
C481 B.n441 VSUBS 0.007061f
C482 B.n442 VSUBS 0.007061f
C483 B.n443 VSUBS 0.007061f
C484 B.n444 VSUBS 0.007061f
C485 B.n445 VSUBS 0.007061f
C486 B.n446 VSUBS 0.007061f
C487 B.n447 VSUBS 0.007061f
C488 B.n448 VSUBS 0.007061f
C489 B.n449 VSUBS 0.007061f
C490 B.n450 VSUBS 0.015487f
C491 B.n451 VSUBS 0.016287f
C492 B.n452 VSUBS 0.016287f
C493 B.n453 VSUBS 0.007061f
C494 B.n454 VSUBS 0.007061f
C495 B.n455 VSUBS 0.007061f
C496 B.n456 VSUBS 0.007061f
C497 B.n457 VSUBS 0.007061f
C498 B.n458 VSUBS 0.007061f
C499 B.n459 VSUBS 0.007061f
C500 B.n460 VSUBS 0.007061f
C501 B.n461 VSUBS 0.007061f
C502 B.n462 VSUBS 0.007061f
C503 B.n463 VSUBS 0.007061f
C504 B.n464 VSUBS 0.007061f
C505 B.n465 VSUBS 0.007061f
C506 B.n466 VSUBS 0.007061f
C507 B.n467 VSUBS 0.007061f
C508 B.n468 VSUBS 0.007061f
C509 B.n469 VSUBS 0.007061f
C510 B.n470 VSUBS 0.007061f
C511 B.n471 VSUBS 0.007061f
C512 B.n472 VSUBS 0.007061f
C513 B.n473 VSUBS 0.007061f
C514 B.n474 VSUBS 0.007061f
C515 B.n475 VSUBS 0.007061f
C516 B.n476 VSUBS 0.007061f
C517 B.n477 VSUBS 0.007061f
C518 B.n478 VSUBS 0.007061f
C519 B.n479 VSUBS 0.007061f
C520 B.n480 VSUBS 0.007061f
C521 B.n481 VSUBS 0.007061f
C522 B.n482 VSUBS 0.007061f
C523 B.n483 VSUBS 0.007061f
C524 B.n484 VSUBS 0.007061f
C525 B.n485 VSUBS 0.007061f
C526 B.n486 VSUBS 0.007061f
C527 B.n487 VSUBS 0.007061f
C528 B.n488 VSUBS 0.007061f
C529 B.n489 VSUBS 0.007061f
C530 B.n490 VSUBS 0.007061f
C531 B.n491 VSUBS 0.007061f
C532 B.n492 VSUBS 0.007061f
C533 B.n493 VSUBS 0.006646f
C534 B.n494 VSUBS 0.007061f
C535 B.n495 VSUBS 0.007061f
C536 B.n496 VSUBS 0.003946f
C537 B.n497 VSUBS 0.007061f
C538 B.n498 VSUBS 0.007061f
C539 B.n499 VSUBS 0.007061f
C540 B.n500 VSUBS 0.007061f
C541 B.n501 VSUBS 0.007061f
C542 B.n502 VSUBS 0.007061f
C543 B.n503 VSUBS 0.007061f
C544 B.n504 VSUBS 0.007061f
C545 B.n505 VSUBS 0.007061f
C546 B.n506 VSUBS 0.007061f
C547 B.n507 VSUBS 0.007061f
C548 B.n508 VSUBS 0.007061f
C549 B.n509 VSUBS 0.003946f
C550 B.n510 VSUBS 0.01636f
C551 B.n511 VSUBS 0.006646f
C552 B.n512 VSUBS 0.007061f
C553 B.n513 VSUBS 0.007061f
C554 B.n514 VSUBS 0.007061f
C555 B.n515 VSUBS 0.007061f
C556 B.n516 VSUBS 0.007061f
C557 B.n517 VSUBS 0.007061f
C558 B.n518 VSUBS 0.007061f
C559 B.n519 VSUBS 0.007061f
C560 B.n520 VSUBS 0.007061f
C561 B.n521 VSUBS 0.007061f
C562 B.n522 VSUBS 0.007061f
C563 B.n523 VSUBS 0.007061f
C564 B.n524 VSUBS 0.007061f
C565 B.n525 VSUBS 0.007061f
C566 B.n526 VSUBS 0.007061f
C567 B.n527 VSUBS 0.007061f
C568 B.n528 VSUBS 0.007061f
C569 B.n529 VSUBS 0.007061f
C570 B.n530 VSUBS 0.007061f
C571 B.n531 VSUBS 0.007061f
C572 B.n532 VSUBS 0.007061f
C573 B.n533 VSUBS 0.007061f
C574 B.n534 VSUBS 0.007061f
C575 B.n535 VSUBS 0.007061f
C576 B.n536 VSUBS 0.007061f
C577 B.n537 VSUBS 0.007061f
C578 B.n538 VSUBS 0.007061f
C579 B.n539 VSUBS 0.007061f
C580 B.n540 VSUBS 0.007061f
C581 B.n541 VSUBS 0.007061f
C582 B.n542 VSUBS 0.007061f
C583 B.n543 VSUBS 0.007061f
C584 B.n544 VSUBS 0.007061f
C585 B.n545 VSUBS 0.007061f
C586 B.n546 VSUBS 0.007061f
C587 B.n547 VSUBS 0.007061f
C588 B.n548 VSUBS 0.007061f
C589 B.n549 VSUBS 0.007061f
C590 B.n550 VSUBS 0.007061f
C591 B.n551 VSUBS 0.007061f
C592 B.n552 VSUBS 0.007061f
C593 B.n553 VSUBS 0.016287f
C594 B.n554 VSUBS 0.016287f
C595 B.n555 VSUBS 0.015487f
C596 B.n556 VSUBS 0.007061f
C597 B.n557 VSUBS 0.007061f
C598 B.n558 VSUBS 0.007061f
C599 B.n559 VSUBS 0.007061f
C600 B.n560 VSUBS 0.007061f
C601 B.n561 VSUBS 0.007061f
C602 B.n562 VSUBS 0.007061f
C603 B.n563 VSUBS 0.007061f
C604 B.n564 VSUBS 0.007061f
C605 B.n565 VSUBS 0.007061f
C606 B.n566 VSUBS 0.007061f
C607 B.n567 VSUBS 0.007061f
C608 B.n568 VSUBS 0.007061f
C609 B.n569 VSUBS 0.007061f
C610 B.n570 VSUBS 0.007061f
C611 B.n571 VSUBS 0.007061f
C612 B.n572 VSUBS 0.007061f
C613 B.n573 VSUBS 0.007061f
C614 B.n574 VSUBS 0.007061f
C615 B.n575 VSUBS 0.007061f
C616 B.n576 VSUBS 0.007061f
C617 B.n577 VSUBS 0.007061f
C618 B.n578 VSUBS 0.007061f
C619 B.n579 VSUBS 0.007061f
C620 B.n580 VSUBS 0.007061f
C621 B.n581 VSUBS 0.007061f
C622 B.n582 VSUBS 0.007061f
C623 B.n583 VSUBS 0.007061f
C624 B.n584 VSUBS 0.007061f
C625 B.n585 VSUBS 0.007061f
C626 B.n586 VSUBS 0.007061f
C627 B.n587 VSUBS 0.007061f
C628 B.n588 VSUBS 0.007061f
C629 B.n589 VSUBS 0.007061f
C630 B.n590 VSUBS 0.007061f
C631 B.n591 VSUBS 0.007061f
C632 B.n592 VSUBS 0.007061f
C633 B.n593 VSUBS 0.007061f
C634 B.n594 VSUBS 0.007061f
C635 B.n595 VSUBS 0.007061f
C636 B.n596 VSUBS 0.007061f
C637 B.n597 VSUBS 0.007061f
C638 B.n598 VSUBS 0.007061f
C639 B.n599 VSUBS 0.007061f
C640 B.n600 VSUBS 0.007061f
C641 B.n601 VSUBS 0.007061f
C642 B.n602 VSUBS 0.007061f
C643 B.n603 VSUBS 0.007061f
C644 B.n604 VSUBS 0.007061f
C645 B.n605 VSUBS 0.007061f
C646 B.n606 VSUBS 0.007061f
C647 B.n607 VSUBS 0.007061f
C648 B.n608 VSUBS 0.007061f
C649 B.n609 VSUBS 0.007061f
C650 B.n610 VSUBS 0.007061f
C651 B.n611 VSUBS 0.007061f
C652 B.n612 VSUBS 0.007061f
C653 B.n613 VSUBS 0.007061f
C654 B.n614 VSUBS 0.007061f
C655 B.n615 VSUBS 0.009214f
C656 B.n616 VSUBS 0.009815f
C657 B.n617 VSUBS 0.019519f
C658 VDD2.t5 VSUBS 1.498f
C659 VDD2.t2 VSUBS 0.158353f
C660 VDD2.t1 VSUBS 0.158353f
C661 VDD2.n0 VSUBS 1.12412f
C662 VDD2.n1 VSUBS 3.1689f
C663 VDD2.t0 VSUBS 1.48451f
C664 VDD2.n2 VSUBS 2.75631f
C665 VDD2.t3 VSUBS 0.158353f
C666 VDD2.t4 VSUBS 0.158353f
C667 VDD2.n3 VSUBS 1.12409f
C668 VN.n0 VSUBS 0.046405f
C669 VN.t4 VSUBS 1.83156f
C670 VN.n1 VSUBS 0.059447f
C671 VN.n2 VSUBS 0.0352f
C672 VN.t3 VSUBS 1.83156f
C673 VN.n3 VSUBS 0.76862f
C674 VN.t0 VSUBS 2.09314f
C675 VN.n4 VSUBS 0.750683f
C676 VN.n5 VSUBS 0.33566f
C677 VN.n6 VSUBS 0.049163f
C678 VN.n7 VSUBS 0.065276f
C679 VN.n8 VSUBS 0.042891f
C680 VN.n9 VSUBS 0.0352f
C681 VN.n10 VSUBS 0.0352f
C682 VN.n11 VSUBS 0.0352f
C683 VN.n12 VSUBS 0.065276f
C684 VN.n13 VSUBS 0.038207f
C685 VN.n14 VSUBS 0.771582f
C686 VN.n15 VSUBS 0.060731f
C687 VN.n16 VSUBS 0.046405f
C688 VN.t5 VSUBS 1.83156f
C689 VN.n17 VSUBS 0.059447f
C690 VN.n18 VSUBS 0.0352f
C691 VN.t2 VSUBS 1.83156f
C692 VN.n19 VSUBS 0.76862f
C693 VN.t1 VSUBS 2.09314f
C694 VN.n20 VSUBS 0.750683f
C695 VN.n21 VSUBS 0.33566f
C696 VN.n22 VSUBS 0.049163f
C697 VN.n23 VSUBS 0.065276f
C698 VN.n24 VSUBS 0.042891f
C699 VN.n25 VSUBS 0.0352f
C700 VN.n26 VSUBS 0.0352f
C701 VN.n27 VSUBS 0.0352f
C702 VN.n28 VSUBS 0.065276f
C703 VN.n29 VSUBS 0.038207f
C704 VN.n30 VSUBS 0.771582f
C705 VN.n31 VSUBS 1.69012f
C706 VDD1.t1 VSUBS 1.27699f
C707 VDD1.t2 VSUBS 1.2761f
C708 VDD1.t0 VSUBS 0.134896f
C709 VDD1.t3 VSUBS 0.134896f
C710 VDD1.n0 VSUBS 0.957601f
C711 VDD1.n1 VSUBS 2.80321f
C712 VDD1.t4 VSUBS 0.134896f
C713 VDD1.t5 VSUBS 0.134896f
C714 VDD1.n2 VSUBS 0.953578f
C715 VDD1.n3 VSUBS 2.34689f
C716 VTAIL.t0 VSUBS 0.192203f
C717 VTAIL.t2 VSUBS 0.192203f
C718 VTAIL.n0 VSUBS 1.2223f
C719 VTAIL.n1 VSUBS 0.881817f
C720 VTAIL.t11 VSUBS 1.65442f
C721 VTAIL.n2 VSUBS 1.15281f
C722 VTAIL.t6 VSUBS 0.192203f
C723 VTAIL.t10 VSUBS 0.192203f
C724 VTAIL.n3 VSUBS 1.2223f
C725 VTAIL.n4 VSUBS 2.48426f
C726 VTAIL.t3 VSUBS 0.192203f
C727 VTAIL.t4 VSUBS 0.192203f
C728 VTAIL.n5 VSUBS 1.22231f
C729 VTAIL.n6 VSUBS 2.48426f
C730 VTAIL.t5 VSUBS 1.65443f
C731 VTAIL.n7 VSUBS 1.1528f
C732 VTAIL.t8 VSUBS 0.192203f
C733 VTAIL.t9 VSUBS 0.192203f
C734 VTAIL.n8 VSUBS 1.22231f
C735 VTAIL.n9 VSUBS 1.06073f
C736 VTAIL.t7 VSUBS 1.65443f
C737 VTAIL.n10 VSUBS 2.32993f
C738 VTAIL.t1 VSUBS 1.65442f
C739 VTAIL.n11 VSUBS 2.26246f
C740 VP.n0 VSUBS 0.04805f
C741 VP.t2 VSUBS 1.89647f
C742 VP.n1 VSUBS 0.061554f
C743 VP.n2 VSUBS 0.036448f
C744 VP.t5 VSUBS 1.89647f
C745 VP.n3 VSUBS 0.693896f
C746 VP.n4 VSUBS 0.036448f
C747 VP.n5 VSUBS 0.061554f
C748 VP.n6 VSUBS 0.04805f
C749 VP.t3 VSUBS 1.89647f
C750 VP.n7 VSUBS 0.04805f
C751 VP.t0 VSUBS 1.89647f
C752 VP.n8 VSUBS 0.061554f
C753 VP.n9 VSUBS 0.036448f
C754 VP.t1 VSUBS 1.89647f
C755 VP.n10 VSUBS 0.795857f
C756 VP.t4 VSUBS 2.16732f
C757 VP.n11 VSUBS 0.777284f
C758 VP.n12 VSUBS 0.347554f
C759 VP.n13 VSUBS 0.050905f
C760 VP.n14 VSUBS 0.067589f
C761 VP.n15 VSUBS 0.044411f
C762 VP.n16 VSUBS 0.036448f
C763 VP.n17 VSUBS 0.036448f
C764 VP.n18 VSUBS 0.036448f
C765 VP.n19 VSUBS 0.067589f
C766 VP.n20 VSUBS 0.039561f
C767 VP.n21 VSUBS 0.798924f
C768 VP.n22 VSUBS 1.73007f
C769 VP.n23 VSUBS 1.75929f
C770 VP.n24 VSUBS 0.798924f
C771 VP.n25 VSUBS 0.039561f
C772 VP.n26 VSUBS 0.067589f
C773 VP.n27 VSUBS 0.036448f
C774 VP.n28 VSUBS 0.036448f
C775 VP.n29 VSUBS 0.036448f
C776 VP.n30 VSUBS 0.044411f
C777 VP.n31 VSUBS 0.067589f
C778 VP.n32 VSUBS 0.050905f
C779 VP.n33 VSUBS 0.036448f
C780 VP.n34 VSUBS 0.036448f
C781 VP.n35 VSUBS 0.050905f
C782 VP.n36 VSUBS 0.067589f
C783 VP.n37 VSUBS 0.044411f
C784 VP.n38 VSUBS 0.036448f
C785 VP.n39 VSUBS 0.036448f
C786 VP.n40 VSUBS 0.036448f
C787 VP.n41 VSUBS 0.067589f
C788 VP.n42 VSUBS 0.039561f
C789 VP.n43 VSUBS 0.798924f
C790 VP.n44 VSUBS 0.062883f
.ends

