* NGSPICE file created from diff_pair_sample_1571.ext - technology: sky130A

.subckt diff_pair_sample_1571 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=0.7878 pd=4.82 as=0 ps=0 w=2.02 l=1.28
X1 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=0.7878 pd=4.82 as=0 ps=0 w=2.02 l=1.28
X2 VDD1.t7 VP.t0 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3333 pd=2.35 as=0.7878 ps=4.82 w=2.02 l=1.28
X3 VTAIL.t5 VN.t0 VDD2.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=0.3333 pd=2.35 as=0.3333 ps=2.35 w=2.02 l=1.28
X4 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=0.7878 pd=4.82 as=0 ps=0 w=2.02 l=1.28
X5 VTAIL.t13 VP.t1 VDD1.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=0.3333 pd=2.35 as=0.3333 ps=2.35 w=2.02 l=1.28
X6 VDD2.t6 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3333 pd=2.35 as=0.3333 ps=2.35 w=2.02 l=1.28
X7 VDD2.t5 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.3333 pd=2.35 as=0.7878 ps=4.82 w=2.02 l=1.28
X8 VTAIL.t12 VP.t2 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.7878 pd=4.82 as=0.3333 ps=2.35 w=2.02 l=1.28
X9 VTAIL.t4 VN.t3 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.3333 pd=2.35 as=0.3333 ps=2.35 w=2.02 l=1.28
X10 VDD2.t3 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3333 pd=2.35 as=0.7878 ps=4.82 w=2.02 l=1.28
X11 VDD1.t4 VP.t3 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3333 pd=2.35 as=0.3333 ps=2.35 w=2.02 l=1.28
X12 VDD1.t3 VP.t4 VTAIL.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=0.3333 pd=2.35 as=0.7878 ps=4.82 w=2.02 l=1.28
X13 VTAIL.t9 VP.t5 VDD1.t2 B.t6 sky130_fd_pr__nfet_01v8 ad=0.7878 pd=4.82 as=0.3333 ps=2.35 w=2.02 l=1.28
X14 VTAIL.t10 VP.t6 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=0.3333 pd=2.35 as=0.3333 ps=2.35 w=2.02 l=1.28
X15 VTAIL.t2 VN.t5 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.7878 pd=4.82 as=0.3333 ps=2.35 w=2.02 l=1.28
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.7878 pd=4.82 as=0 ps=0 w=2.02 l=1.28
X17 VDD2.t1 VN.t6 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.3333 pd=2.35 as=0.3333 ps=2.35 w=2.02 l=1.28
X18 VDD1.t0 VP.t7 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=0.3333 pd=2.35 as=0.3333 ps=2.35 w=2.02 l=1.28
X19 VTAIL.t6 VN.t7 VDD2.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=0.7878 pd=4.82 as=0.3333 ps=2.35 w=2.02 l=1.28
R0 B.n438 B.n437 585
R1 B.n147 B.n78 585
R2 B.n146 B.n145 585
R3 B.n144 B.n143 585
R4 B.n142 B.n141 585
R5 B.n140 B.n139 585
R6 B.n138 B.n137 585
R7 B.n136 B.n135 585
R8 B.n134 B.n133 585
R9 B.n132 B.n131 585
R10 B.n130 B.n129 585
R11 B.n128 B.n127 585
R12 B.n126 B.n125 585
R13 B.n124 B.n123 585
R14 B.n122 B.n121 585
R15 B.n120 B.n119 585
R16 B.n118 B.n117 585
R17 B.n116 B.n115 585
R18 B.n114 B.n113 585
R19 B.n112 B.n111 585
R20 B.n110 B.n109 585
R21 B.n108 B.n107 585
R22 B.n106 B.n105 585
R23 B.n104 B.n103 585
R24 B.n102 B.n101 585
R25 B.n100 B.n99 585
R26 B.n98 B.n97 585
R27 B.n96 B.n95 585
R28 B.n94 B.n93 585
R29 B.n92 B.n91 585
R30 B.n90 B.n89 585
R31 B.n88 B.n87 585
R32 B.n86 B.n85 585
R33 B.n60 B.n59 585
R34 B.n436 B.n61 585
R35 B.n441 B.n61 585
R36 B.n435 B.n434 585
R37 B.n434 B.n57 585
R38 B.n433 B.n56 585
R39 B.n447 B.n56 585
R40 B.n432 B.n55 585
R41 B.n448 B.n55 585
R42 B.n431 B.n54 585
R43 B.n449 B.n54 585
R44 B.n430 B.n429 585
R45 B.n429 B.n53 585
R46 B.n428 B.n49 585
R47 B.n455 B.n49 585
R48 B.n427 B.n48 585
R49 B.n456 B.n48 585
R50 B.n426 B.n47 585
R51 B.n457 B.n47 585
R52 B.n425 B.n424 585
R53 B.n424 B.n43 585
R54 B.n423 B.n42 585
R55 B.n463 B.n42 585
R56 B.n422 B.n41 585
R57 B.n464 B.n41 585
R58 B.n421 B.n40 585
R59 B.n465 B.n40 585
R60 B.n420 B.n419 585
R61 B.n419 B.n39 585
R62 B.n418 B.n35 585
R63 B.n471 B.n35 585
R64 B.n417 B.n34 585
R65 B.n472 B.n34 585
R66 B.n416 B.n33 585
R67 B.n473 B.n33 585
R68 B.n415 B.n414 585
R69 B.n414 B.n29 585
R70 B.n413 B.n28 585
R71 B.n479 B.n28 585
R72 B.n412 B.n27 585
R73 B.n480 B.n27 585
R74 B.n411 B.n26 585
R75 B.n481 B.n26 585
R76 B.n410 B.n409 585
R77 B.n409 B.n22 585
R78 B.n408 B.n21 585
R79 B.n487 B.n21 585
R80 B.n407 B.n20 585
R81 B.n488 B.n20 585
R82 B.n406 B.n19 585
R83 B.n489 B.n19 585
R84 B.n405 B.n404 585
R85 B.n404 B.n15 585
R86 B.n403 B.n14 585
R87 B.n495 B.n14 585
R88 B.n402 B.n13 585
R89 B.n496 B.n13 585
R90 B.n401 B.n12 585
R91 B.n497 B.n12 585
R92 B.n400 B.n399 585
R93 B.n399 B.n8 585
R94 B.n398 B.n7 585
R95 B.n503 B.n7 585
R96 B.n397 B.n6 585
R97 B.n504 B.n6 585
R98 B.n396 B.n5 585
R99 B.n505 B.n5 585
R100 B.n395 B.n394 585
R101 B.n394 B.n4 585
R102 B.n393 B.n148 585
R103 B.n393 B.n392 585
R104 B.n383 B.n149 585
R105 B.n150 B.n149 585
R106 B.n385 B.n384 585
R107 B.n386 B.n385 585
R108 B.n382 B.n155 585
R109 B.n155 B.n154 585
R110 B.n381 B.n380 585
R111 B.n380 B.n379 585
R112 B.n157 B.n156 585
R113 B.n158 B.n157 585
R114 B.n372 B.n371 585
R115 B.n373 B.n372 585
R116 B.n370 B.n162 585
R117 B.n166 B.n162 585
R118 B.n369 B.n368 585
R119 B.n368 B.n367 585
R120 B.n164 B.n163 585
R121 B.n165 B.n164 585
R122 B.n360 B.n359 585
R123 B.n361 B.n360 585
R124 B.n358 B.n171 585
R125 B.n171 B.n170 585
R126 B.n357 B.n356 585
R127 B.n356 B.n355 585
R128 B.n173 B.n172 585
R129 B.n174 B.n173 585
R130 B.n348 B.n347 585
R131 B.n349 B.n348 585
R132 B.n346 B.n179 585
R133 B.n179 B.n178 585
R134 B.n345 B.n344 585
R135 B.n344 B.n343 585
R136 B.n181 B.n180 585
R137 B.n336 B.n181 585
R138 B.n335 B.n334 585
R139 B.n337 B.n335 585
R140 B.n333 B.n186 585
R141 B.n186 B.n185 585
R142 B.n332 B.n331 585
R143 B.n331 B.n330 585
R144 B.n188 B.n187 585
R145 B.n189 B.n188 585
R146 B.n323 B.n322 585
R147 B.n324 B.n323 585
R148 B.n321 B.n194 585
R149 B.n194 B.n193 585
R150 B.n320 B.n319 585
R151 B.n319 B.n318 585
R152 B.n196 B.n195 585
R153 B.n311 B.n196 585
R154 B.n310 B.n309 585
R155 B.n312 B.n310 585
R156 B.n308 B.n201 585
R157 B.n201 B.n200 585
R158 B.n307 B.n306 585
R159 B.n306 B.n305 585
R160 B.n203 B.n202 585
R161 B.n204 B.n203 585
R162 B.n298 B.n297 585
R163 B.n299 B.n298 585
R164 B.n207 B.n206 585
R165 B.n230 B.n228 585
R166 B.n231 B.n227 585
R167 B.n231 B.n208 585
R168 B.n234 B.n233 585
R169 B.n235 B.n226 585
R170 B.n237 B.n236 585
R171 B.n239 B.n225 585
R172 B.n242 B.n241 585
R173 B.n243 B.n224 585
R174 B.n245 B.n244 585
R175 B.n247 B.n223 585
R176 B.n250 B.n249 585
R177 B.n252 B.n220 585
R178 B.n254 B.n253 585
R179 B.n256 B.n219 585
R180 B.n259 B.n258 585
R181 B.n260 B.n218 585
R182 B.n262 B.n261 585
R183 B.n264 B.n217 585
R184 B.n267 B.n266 585
R185 B.n268 B.n216 585
R186 B.n273 B.n272 585
R187 B.n275 B.n215 585
R188 B.n278 B.n277 585
R189 B.n279 B.n214 585
R190 B.n281 B.n280 585
R191 B.n283 B.n213 585
R192 B.n286 B.n285 585
R193 B.n287 B.n212 585
R194 B.n289 B.n288 585
R195 B.n291 B.n211 585
R196 B.n292 B.n210 585
R197 B.n295 B.n294 585
R198 B.n296 B.n209 585
R199 B.n209 B.n208 585
R200 B.n301 B.n300 585
R201 B.n300 B.n299 585
R202 B.n302 B.n205 585
R203 B.n205 B.n204 585
R204 B.n304 B.n303 585
R205 B.n305 B.n304 585
R206 B.n199 B.n198 585
R207 B.n200 B.n199 585
R208 B.n314 B.n313 585
R209 B.n313 B.n312 585
R210 B.n315 B.n197 585
R211 B.n311 B.n197 585
R212 B.n317 B.n316 585
R213 B.n318 B.n317 585
R214 B.n192 B.n191 585
R215 B.n193 B.n192 585
R216 B.n326 B.n325 585
R217 B.n325 B.n324 585
R218 B.n327 B.n190 585
R219 B.n190 B.n189 585
R220 B.n329 B.n328 585
R221 B.n330 B.n329 585
R222 B.n184 B.n183 585
R223 B.n185 B.n184 585
R224 B.n339 B.n338 585
R225 B.n338 B.n337 585
R226 B.n340 B.n182 585
R227 B.n336 B.n182 585
R228 B.n342 B.n341 585
R229 B.n343 B.n342 585
R230 B.n177 B.n176 585
R231 B.n178 B.n177 585
R232 B.n351 B.n350 585
R233 B.n350 B.n349 585
R234 B.n352 B.n175 585
R235 B.n175 B.n174 585
R236 B.n354 B.n353 585
R237 B.n355 B.n354 585
R238 B.n169 B.n168 585
R239 B.n170 B.n169 585
R240 B.n363 B.n362 585
R241 B.n362 B.n361 585
R242 B.n364 B.n167 585
R243 B.n167 B.n165 585
R244 B.n366 B.n365 585
R245 B.n367 B.n366 585
R246 B.n161 B.n160 585
R247 B.n166 B.n161 585
R248 B.n375 B.n374 585
R249 B.n374 B.n373 585
R250 B.n376 B.n159 585
R251 B.n159 B.n158 585
R252 B.n378 B.n377 585
R253 B.n379 B.n378 585
R254 B.n153 B.n152 585
R255 B.n154 B.n153 585
R256 B.n388 B.n387 585
R257 B.n387 B.n386 585
R258 B.n389 B.n151 585
R259 B.n151 B.n150 585
R260 B.n391 B.n390 585
R261 B.n392 B.n391 585
R262 B.n2 B.n0 585
R263 B.n4 B.n2 585
R264 B.n3 B.n1 585
R265 B.n504 B.n3 585
R266 B.n502 B.n501 585
R267 B.n503 B.n502 585
R268 B.n500 B.n9 585
R269 B.n9 B.n8 585
R270 B.n499 B.n498 585
R271 B.n498 B.n497 585
R272 B.n11 B.n10 585
R273 B.n496 B.n11 585
R274 B.n494 B.n493 585
R275 B.n495 B.n494 585
R276 B.n492 B.n16 585
R277 B.n16 B.n15 585
R278 B.n491 B.n490 585
R279 B.n490 B.n489 585
R280 B.n18 B.n17 585
R281 B.n488 B.n18 585
R282 B.n486 B.n485 585
R283 B.n487 B.n486 585
R284 B.n484 B.n23 585
R285 B.n23 B.n22 585
R286 B.n483 B.n482 585
R287 B.n482 B.n481 585
R288 B.n25 B.n24 585
R289 B.n480 B.n25 585
R290 B.n478 B.n477 585
R291 B.n479 B.n478 585
R292 B.n476 B.n30 585
R293 B.n30 B.n29 585
R294 B.n475 B.n474 585
R295 B.n474 B.n473 585
R296 B.n32 B.n31 585
R297 B.n472 B.n32 585
R298 B.n470 B.n469 585
R299 B.n471 B.n470 585
R300 B.n468 B.n36 585
R301 B.n39 B.n36 585
R302 B.n467 B.n466 585
R303 B.n466 B.n465 585
R304 B.n38 B.n37 585
R305 B.n464 B.n38 585
R306 B.n462 B.n461 585
R307 B.n463 B.n462 585
R308 B.n460 B.n44 585
R309 B.n44 B.n43 585
R310 B.n459 B.n458 585
R311 B.n458 B.n457 585
R312 B.n46 B.n45 585
R313 B.n456 B.n46 585
R314 B.n454 B.n453 585
R315 B.n455 B.n454 585
R316 B.n452 B.n50 585
R317 B.n53 B.n50 585
R318 B.n451 B.n450 585
R319 B.n450 B.n449 585
R320 B.n52 B.n51 585
R321 B.n448 B.n52 585
R322 B.n446 B.n445 585
R323 B.n447 B.n446 585
R324 B.n444 B.n58 585
R325 B.n58 B.n57 585
R326 B.n443 B.n442 585
R327 B.n442 B.n441 585
R328 B.n507 B.n506 585
R329 B.n506 B.n505 585
R330 B.n300 B.n207 473.281
R331 B.n442 B.n60 473.281
R332 B.n298 B.n209 473.281
R333 B.n438 B.n61 473.281
R334 B.n440 B.n439 256.663
R335 B.n440 B.n77 256.663
R336 B.n440 B.n76 256.663
R337 B.n440 B.n75 256.663
R338 B.n440 B.n74 256.663
R339 B.n440 B.n73 256.663
R340 B.n440 B.n72 256.663
R341 B.n440 B.n71 256.663
R342 B.n440 B.n70 256.663
R343 B.n440 B.n69 256.663
R344 B.n440 B.n68 256.663
R345 B.n440 B.n67 256.663
R346 B.n440 B.n66 256.663
R347 B.n440 B.n65 256.663
R348 B.n440 B.n64 256.663
R349 B.n440 B.n63 256.663
R350 B.n440 B.n62 256.663
R351 B.n229 B.n208 256.663
R352 B.n232 B.n208 256.663
R353 B.n238 B.n208 256.663
R354 B.n240 B.n208 256.663
R355 B.n246 B.n208 256.663
R356 B.n248 B.n208 256.663
R357 B.n255 B.n208 256.663
R358 B.n257 B.n208 256.663
R359 B.n263 B.n208 256.663
R360 B.n265 B.n208 256.663
R361 B.n274 B.n208 256.663
R362 B.n276 B.n208 256.663
R363 B.n282 B.n208 256.663
R364 B.n284 B.n208 256.663
R365 B.n290 B.n208 256.663
R366 B.n293 B.n208 256.663
R367 B.n269 B.t19 242.548
R368 B.n221 B.t15 242.548
R369 B.n82 B.t12 242.548
R370 B.n79 B.t8 242.548
R371 B.n299 B.n208 164.359
R372 B.n441 B.n440 164.359
R373 B.n300 B.n205 163.367
R374 B.n304 B.n205 163.367
R375 B.n304 B.n199 163.367
R376 B.n313 B.n199 163.367
R377 B.n313 B.n197 163.367
R378 B.n317 B.n197 163.367
R379 B.n317 B.n192 163.367
R380 B.n325 B.n192 163.367
R381 B.n325 B.n190 163.367
R382 B.n329 B.n190 163.367
R383 B.n329 B.n184 163.367
R384 B.n338 B.n184 163.367
R385 B.n338 B.n182 163.367
R386 B.n342 B.n182 163.367
R387 B.n342 B.n177 163.367
R388 B.n350 B.n177 163.367
R389 B.n350 B.n175 163.367
R390 B.n354 B.n175 163.367
R391 B.n354 B.n169 163.367
R392 B.n362 B.n169 163.367
R393 B.n362 B.n167 163.367
R394 B.n366 B.n167 163.367
R395 B.n366 B.n161 163.367
R396 B.n374 B.n161 163.367
R397 B.n374 B.n159 163.367
R398 B.n378 B.n159 163.367
R399 B.n378 B.n153 163.367
R400 B.n387 B.n153 163.367
R401 B.n387 B.n151 163.367
R402 B.n391 B.n151 163.367
R403 B.n391 B.n2 163.367
R404 B.n506 B.n2 163.367
R405 B.n506 B.n3 163.367
R406 B.n502 B.n3 163.367
R407 B.n502 B.n9 163.367
R408 B.n498 B.n9 163.367
R409 B.n498 B.n11 163.367
R410 B.n494 B.n11 163.367
R411 B.n494 B.n16 163.367
R412 B.n490 B.n16 163.367
R413 B.n490 B.n18 163.367
R414 B.n486 B.n18 163.367
R415 B.n486 B.n23 163.367
R416 B.n482 B.n23 163.367
R417 B.n482 B.n25 163.367
R418 B.n478 B.n25 163.367
R419 B.n478 B.n30 163.367
R420 B.n474 B.n30 163.367
R421 B.n474 B.n32 163.367
R422 B.n470 B.n32 163.367
R423 B.n470 B.n36 163.367
R424 B.n466 B.n36 163.367
R425 B.n466 B.n38 163.367
R426 B.n462 B.n38 163.367
R427 B.n462 B.n44 163.367
R428 B.n458 B.n44 163.367
R429 B.n458 B.n46 163.367
R430 B.n454 B.n46 163.367
R431 B.n454 B.n50 163.367
R432 B.n450 B.n50 163.367
R433 B.n450 B.n52 163.367
R434 B.n446 B.n52 163.367
R435 B.n446 B.n58 163.367
R436 B.n442 B.n58 163.367
R437 B.n231 B.n230 163.367
R438 B.n233 B.n231 163.367
R439 B.n237 B.n226 163.367
R440 B.n241 B.n239 163.367
R441 B.n245 B.n224 163.367
R442 B.n249 B.n247 163.367
R443 B.n254 B.n220 163.367
R444 B.n258 B.n256 163.367
R445 B.n262 B.n218 163.367
R446 B.n266 B.n264 163.367
R447 B.n273 B.n216 163.367
R448 B.n277 B.n275 163.367
R449 B.n281 B.n214 163.367
R450 B.n285 B.n283 163.367
R451 B.n289 B.n212 163.367
R452 B.n292 B.n291 163.367
R453 B.n294 B.n209 163.367
R454 B.n298 B.n203 163.367
R455 B.n306 B.n203 163.367
R456 B.n306 B.n201 163.367
R457 B.n310 B.n201 163.367
R458 B.n310 B.n196 163.367
R459 B.n319 B.n196 163.367
R460 B.n319 B.n194 163.367
R461 B.n323 B.n194 163.367
R462 B.n323 B.n188 163.367
R463 B.n331 B.n188 163.367
R464 B.n331 B.n186 163.367
R465 B.n335 B.n186 163.367
R466 B.n335 B.n181 163.367
R467 B.n344 B.n181 163.367
R468 B.n344 B.n179 163.367
R469 B.n348 B.n179 163.367
R470 B.n348 B.n173 163.367
R471 B.n356 B.n173 163.367
R472 B.n356 B.n171 163.367
R473 B.n360 B.n171 163.367
R474 B.n360 B.n164 163.367
R475 B.n368 B.n164 163.367
R476 B.n368 B.n162 163.367
R477 B.n372 B.n162 163.367
R478 B.n372 B.n157 163.367
R479 B.n380 B.n157 163.367
R480 B.n380 B.n155 163.367
R481 B.n385 B.n155 163.367
R482 B.n385 B.n149 163.367
R483 B.n393 B.n149 163.367
R484 B.n394 B.n393 163.367
R485 B.n394 B.n5 163.367
R486 B.n6 B.n5 163.367
R487 B.n7 B.n6 163.367
R488 B.n399 B.n7 163.367
R489 B.n399 B.n12 163.367
R490 B.n13 B.n12 163.367
R491 B.n14 B.n13 163.367
R492 B.n404 B.n14 163.367
R493 B.n404 B.n19 163.367
R494 B.n20 B.n19 163.367
R495 B.n21 B.n20 163.367
R496 B.n409 B.n21 163.367
R497 B.n409 B.n26 163.367
R498 B.n27 B.n26 163.367
R499 B.n28 B.n27 163.367
R500 B.n414 B.n28 163.367
R501 B.n414 B.n33 163.367
R502 B.n34 B.n33 163.367
R503 B.n35 B.n34 163.367
R504 B.n419 B.n35 163.367
R505 B.n419 B.n40 163.367
R506 B.n41 B.n40 163.367
R507 B.n42 B.n41 163.367
R508 B.n424 B.n42 163.367
R509 B.n424 B.n47 163.367
R510 B.n48 B.n47 163.367
R511 B.n49 B.n48 163.367
R512 B.n429 B.n49 163.367
R513 B.n429 B.n54 163.367
R514 B.n55 B.n54 163.367
R515 B.n56 B.n55 163.367
R516 B.n434 B.n56 163.367
R517 B.n434 B.n61 163.367
R518 B.n87 B.n86 163.367
R519 B.n91 B.n90 163.367
R520 B.n95 B.n94 163.367
R521 B.n99 B.n98 163.367
R522 B.n103 B.n102 163.367
R523 B.n107 B.n106 163.367
R524 B.n111 B.n110 163.367
R525 B.n115 B.n114 163.367
R526 B.n119 B.n118 163.367
R527 B.n123 B.n122 163.367
R528 B.n127 B.n126 163.367
R529 B.n131 B.n130 163.367
R530 B.n135 B.n134 163.367
R531 B.n139 B.n138 163.367
R532 B.n143 B.n142 163.367
R533 B.n145 B.n78 163.367
R534 B.n269 B.t21 154.631
R535 B.n79 B.t10 154.631
R536 B.n221 B.t18 154.631
R537 B.n82 B.t13 154.631
R538 B.n270 B.t20 123.406
R539 B.n80 B.t11 123.406
R540 B.n222 B.t17 123.406
R541 B.n83 B.t14 123.406
R542 B.n299 B.n204 102.537
R543 B.n305 B.n204 102.537
R544 B.n305 B.n200 102.537
R545 B.n312 B.n200 102.537
R546 B.n312 B.n311 102.537
R547 B.n318 B.n193 102.537
R548 B.n324 B.n193 102.537
R549 B.n324 B.n189 102.537
R550 B.n330 B.n189 102.537
R551 B.n330 B.n185 102.537
R552 B.n337 B.n185 102.537
R553 B.n337 B.n336 102.537
R554 B.n343 B.n178 102.537
R555 B.n349 B.n178 102.537
R556 B.n349 B.n174 102.537
R557 B.n355 B.n174 102.537
R558 B.n361 B.n170 102.537
R559 B.n361 B.n165 102.537
R560 B.n367 B.n165 102.537
R561 B.n367 B.n166 102.537
R562 B.n373 B.n158 102.537
R563 B.n379 B.n158 102.537
R564 B.n379 B.n154 102.537
R565 B.n386 B.n154 102.537
R566 B.n392 B.n150 102.537
R567 B.n392 B.n4 102.537
R568 B.n505 B.n4 102.537
R569 B.n505 B.n504 102.537
R570 B.n504 B.n503 102.537
R571 B.n503 B.n8 102.537
R572 B.n497 B.n496 102.537
R573 B.n496 B.n495 102.537
R574 B.n495 B.n15 102.537
R575 B.n489 B.n15 102.537
R576 B.n488 B.n487 102.537
R577 B.n487 B.n22 102.537
R578 B.n481 B.n22 102.537
R579 B.n481 B.n480 102.537
R580 B.n479 B.n29 102.537
R581 B.n473 B.n29 102.537
R582 B.n473 B.n472 102.537
R583 B.n472 B.n471 102.537
R584 B.n465 B.n39 102.537
R585 B.n465 B.n464 102.537
R586 B.n464 B.n463 102.537
R587 B.n463 B.n43 102.537
R588 B.n457 B.n43 102.537
R589 B.n457 B.n456 102.537
R590 B.n456 B.n455 102.537
R591 B.n449 B.n53 102.537
R592 B.n449 B.n448 102.537
R593 B.n448 B.n447 102.537
R594 B.n447 B.n57 102.537
R595 B.n441 B.n57 102.537
R596 B.t0 B.n150 99.5207
R597 B.t6 B.n8 99.5207
R598 B.n311 B.t16 90.4734
R599 B.n53 B.t9 90.4734
R600 B.n336 B.t2 84.4419
R601 B.n39 B.t3 84.4419
R602 B.n373 B.t4 72.3788
R603 B.n489 B.t7 72.3788
R604 B.n229 B.n207 71.676
R605 B.n233 B.n232 71.676
R606 B.n238 B.n237 71.676
R607 B.n241 B.n240 71.676
R608 B.n246 B.n245 71.676
R609 B.n249 B.n248 71.676
R610 B.n255 B.n254 71.676
R611 B.n258 B.n257 71.676
R612 B.n263 B.n262 71.676
R613 B.n266 B.n265 71.676
R614 B.n274 B.n273 71.676
R615 B.n277 B.n276 71.676
R616 B.n282 B.n281 71.676
R617 B.n285 B.n284 71.676
R618 B.n290 B.n289 71.676
R619 B.n293 B.n292 71.676
R620 B.n62 B.n60 71.676
R621 B.n87 B.n63 71.676
R622 B.n91 B.n64 71.676
R623 B.n95 B.n65 71.676
R624 B.n99 B.n66 71.676
R625 B.n103 B.n67 71.676
R626 B.n107 B.n68 71.676
R627 B.n111 B.n69 71.676
R628 B.n115 B.n70 71.676
R629 B.n119 B.n71 71.676
R630 B.n123 B.n72 71.676
R631 B.n127 B.n73 71.676
R632 B.n131 B.n74 71.676
R633 B.n135 B.n75 71.676
R634 B.n139 B.n76 71.676
R635 B.n143 B.n77 71.676
R636 B.n439 B.n78 71.676
R637 B.n439 B.n438 71.676
R638 B.n145 B.n77 71.676
R639 B.n142 B.n76 71.676
R640 B.n138 B.n75 71.676
R641 B.n134 B.n74 71.676
R642 B.n130 B.n73 71.676
R643 B.n126 B.n72 71.676
R644 B.n122 B.n71 71.676
R645 B.n118 B.n70 71.676
R646 B.n114 B.n69 71.676
R647 B.n110 B.n68 71.676
R648 B.n106 B.n67 71.676
R649 B.n102 B.n66 71.676
R650 B.n98 B.n65 71.676
R651 B.n94 B.n64 71.676
R652 B.n90 B.n63 71.676
R653 B.n86 B.n62 71.676
R654 B.n230 B.n229 71.676
R655 B.n232 B.n226 71.676
R656 B.n239 B.n238 71.676
R657 B.n240 B.n224 71.676
R658 B.n247 B.n246 71.676
R659 B.n248 B.n220 71.676
R660 B.n256 B.n255 71.676
R661 B.n257 B.n218 71.676
R662 B.n264 B.n263 71.676
R663 B.n265 B.n216 71.676
R664 B.n275 B.n274 71.676
R665 B.n276 B.n214 71.676
R666 B.n283 B.n282 71.676
R667 B.n284 B.n212 71.676
R668 B.n291 B.n290 71.676
R669 B.n294 B.n293 71.676
R670 B.n271 B.n270 59.5399
R671 B.n251 B.n222 59.5399
R672 B.n84 B.n83 59.5399
R673 B.n81 B.n80 59.5399
R674 B.n355 B.t1 57.3
R675 B.t5 B.n479 57.3
R676 B.t1 B.n170 45.237
R677 B.n480 B.t5 45.237
R678 B.n270 B.n269 31.2247
R679 B.n222 B.n221 31.2247
R680 B.n83 B.n82 31.2247
R681 B.n80 B.n79 31.2247
R682 B.n443 B.n59 30.7517
R683 B.n437 B.n436 30.7517
R684 B.n297 B.n296 30.7517
R685 B.n301 B.n206 30.7517
R686 B.n166 B.t4 30.1581
R687 B.t7 B.n488 30.1581
R688 B.n343 B.t2 18.0951
R689 B.n471 B.t3 18.0951
R690 B B.n507 18.0485
R691 B.n318 B.t16 12.0636
R692 B.n455 B.t9 12.0636
R693 B.n85 B.n59 10.6151
R694 B.n88 B.n85 10.6151
R695 B.n89 B.n88 10.6151
R696 B.n92 B.n89 10.6151
R697 B.n93 B.n92 10.6151
R698 B.n96 B.n93 10.6151
R699 B.n97 B.n96 10.6151
R700 B.n100 B.n97 10.6151
R701 B.n101 B.n100 10.6151
R702 B.n104 B.n101 10.6151
R703 B.n105 B.n104 10.6151
R704 B.n109 B.n108 10.6151
R705 B.n112 B.n109 10.6151
R706 B.n113 B.n112 10.6151
R707 B.n116 B.n113 10.6151
R708 B.n117 B.n116 10.6151
R709 B.n120 B.n117 10.6151
R710 B.n121 B.n120 10.6151
R711 B.n124 B.n121 10.6151
R712 B.n125 B.n124 10.6151
R713 B.n129 B.n128 10.6151
R714 B.n132 B.n129 10.6151
R715 B.n133 B.n132 10.6151
R716 B.n136 B.n133 10.6151
R717 B.n137 B.n136 10.6151
R718 B.n140 B.n137 10.6151
R719 B.n141 B.n140 10.6151
R720 B.n144 B.n141 10.6151
R721 B.n146 B.n144 10.6151
R722 B.n147 B.n146 10.6151
R723 B.n437 B.n147 10.6151
R724 B.n297 B.n202 10.6151
R725 B.n307 B.n202 10.6151
R726 B.n308 B.n307 10.6151
R727 B.n309 B.n308 10.6151
R728 B.n309 B.n195 10.6151
R729 B.n320 B.n195 10.6151
R730 B.n321 B.n320 10.6151
R731 B.n322 B.n321 10.6151
R732 B.n322 B.n187 10.6151
R733 B.n332 B.n187 10.6151
R734 B.n333 B.n332 10.6151
R735 B.n334 B.n333 10.6151
R736 B.n334 B.n180 10.6151
R737 B.n345 B.n180 10.6151
R738 B.n346 B.n345 10.6151
R739 B.n347 B.n346 10.6151
R740 B.n347 B.n172 10.6151
R741 B.n357 B.n172 10.6151
R742 B.n358 B.n357 10.6151
R743 B.n359 B.n358 10.6151
R744 B.n359 B.n163 10.6151
R745 B.n369 B.n163 10.6151
R746 B.n370 B.n369 10.6151
R747 B.n371 B.n370 10.6151
R748 B.n371 B.n156 10.6151
R749 B.n381 B.n156 10.6151
R750 B.n382 B.n381 10.6151
R751 B.n384 B.n382 10.6151
R752 B.n384 B.n383 10.6151
R753 B.n383 B.n148 10.6151
R754 B.n395 B.n148 10.6151
R755 B.n396 B.n395 10.6151
R756 B.n397 B.n396 10.6151
R757 B.n398 B.n397 10.6151
R758 B.n400 B.n398 10.6151
R759 B.n401 B.n400 10.6151
R760 B.n402 B.n401 10.6151
R761 B.n403 B.n402 10.6151
R762 B.n405 B.n403 10.6151
R763 B.n406 B.n405 10.6151
R764 B.n407 B.n406 10.6151
R765 B.n408 B.n407 10.6151
R766 B.n410 B.n408 10.6151
R767 B.n411 B.n410 10.6151
R768 B.n412 B.n411 10.6151
R769 B.n413 B.n412 10.6151
R770 B.n415 B.n413 10.6151
R771 B.n416 B.n415 10.6151
R772 B.n417 B.n416 10.6151
R773 B.n418 B.n417 10.6151
R774 B.n420 B.n418 10.6151
R775 B.n421 B.n420 10.6151
R776 B.n422 B.n421 10.6151
R777 B.n423 B.n422 10.6151
R778 B.n425 B.n423 10.6151
R779 B.n426 B.n425 10.6151
R780 B.n427 B.n426 10.6151
R781 B.n428 B.n427 10.6151
R782 B.n430 B.n428 10.6151
R783 B.n431 B.n430 10.6151
R784 B.n432 B.n431 10.6151
R785 B.n433 B.n432 10.6151
R786 B.n435 B.n433 10.6151
R787 B.n436 B.n435 10.6151
R788 B.n228 B.n206 10.6151
R789 B.n228 B.n227 10.6151
R790 B.n234 B.n227 10.6151
R791 B.n235 B.n234 10.6151
R792 B.n236 B.n235 10.6151
R793 B.n236 B.n225 10.6151
R794 B.n242 B.n225 10.6151
R795 B.n243 B.n242 10.6151
R796 B.n244 B.n243 10.6151
R797 B.n244 B.n223 10.6151
R798 B.n250 B.n223 10.6151
R799 B.n253 B.n252 10.6151
R800 B.n253 B.n219 10.6151
R801 B.n259 B.n219 10.6151
R802 B.n260 B.n259 10.6151
R803 B.n261 B.n260 10.6151
R804 B.n261 B.n217 10.6151
R805 B.n267 B.n217 10.6151
R806 B.n268 B.n267 10.6151
R807 B.n272 B.n268 10.6151
R808 B.n278 B.n215 10.6151
R809 B.n279 B.n278 10.6151
R810 B.n280 B.n279 10.6151
R811 B.n280 B.n213 10.6151
R812 B.n286 B.n213 10.6151
R813 B.n287 B.n286 10.6151
R814 B.n288 B.n287 10.6151
R815 B.n288 B.n211 10.6151
R816 B.n211 B.n210 10.6151
R817 B.n295 B.n210 10.6151
R818 B.n296 B.n295 10.6151
R819 B.n302 B.n301 10.6151
R820 B.n303 B.n302 10.6151
R821 B.n303 B.n198 10.6151
R822 B.n314 B.n198 10.6151
R823 B.n315 B.n314 10.6151
R824 B.n316 B.n315 10.6151
R825 B.n316 B.n191 10.6151
R826 B.n326 B.n191 10.6151
R827 B.n327 B.n326 10.6151
R828 B.n328 B.n327 10.6151
R829 B.n328 B.n183 10.6151
R830 B.n339 B.n183 10.6151
R831 B.n340 B.n339 10.6151
R832 B.n341 B.n340 10.6151
R833 B.n341 B.n176 10.6151
R834 B.n351 B.n176 10.6151
R835 B.n352 B.n351 10.6151
R836 B.n353 B.n352 10.6151
R837 B.n353 B.n168 10.6151
R838 B.n363 B.n168 10.6151
R839 B.n364 B.n363 10.6151
R840 B.n365 B.n364 10.6151
R841 B.n365 B.n160 10.6151
R842 B.n375 B.n160 10.6151
R843 B.n376 B.n375 10.6151
R844 B.n377 B.n376 10.6151
R845 B.n377 B.n152 10.6151
R846 B.n388 B.n152 10.6151
R847 B.n389 B.n388 10.6151
R848 B.n390 B.n389 10.6151
R849 B.n390 B.n0 10.6151
R850 B.n501 B.n1 10.6151
R851 B.n501 B.n500 10.6151
R852 B.n500 B.n499 10.6151
R853 B.n499 B.n10 10.6151
R854 B.n493 B.n10 10.6151
R855 B.n493 B.n492 10.6151
R856 B.n492 B.n491 10.6151
R857 B.n491 B.n17 10.6151
R858 B.n485 B.n17 10.6151
R859 B.n485 B.n484 10.6151
R860 B.n484 B.n483 10.6151
R861 B.n483 B.n24 10.6151
R862 B.n477 B.n24 10.6151
R863 B.n477 B.n476 10.6151
R864 B.n476 B.n475 10.6151
R865 B.n475 B.n31 10.6151
R866 B.n469 B.n31 10.6151
R867 B.n469 B.n468 10.6151
R868 B.n468 B.n467 10.6151
R869 B.n467 B.n37 10.6151
R870 B.n461 B.n37 10.6151
R871 B.n461 B.n460 10.6151
R872 B.n460 B.n459 10.6151
R873 B.n459 B.n45 10.6151
R874 B.n453 B.n45 10.6151
R875 B.n453 B.n452 10.6151
R876 B.n452 B.n451 10.6151
R877 B.n451 B.n51 10.6151
R878 B.n445 B.n51 10.6151
R879 B.n445 B.n444 10.6151
R880 B.n444 B.n443 10.6151
R881 B.n105 B.n84 9.36635
R882 B.n128 B.n81 9.36635
R883 B.n251 B.n250 9.36635
R884 B.n271 B.n215 9.36635
R885 B.n386 B.t0 3.01626
R886 B.n497 B.t6 3.01626
R887 B.n507 B.n0 2.81026
R888 B.n507 B.n1 2.81026
R889 B.n108 B.n84 1.24928
R890 B.n125 B.n81 1.24928
R891 B.n252 B.n251 1.24928
R892 B.n272 B.n271 1.24928
R893 VP.n11 VP.n10 161.3
R894 VP.n12 VP.n7 161.3
R895 VP.n14 VP.n13 161.3
R896 VP.n16 VP.n15 161.3
R897 VP.n17 VP.n5 161.3
R898 VP.n32 VP.n0 161.3
R899 VP.n31 VP.n30 161.3
R900 VP.n29 VP.n28 161.3
R901 VP.n27 VP.n2 161.3
R902 VP.n26 VP.n25 161.3
R903 VP.n24 VP.n23 161.3
R904 VP.n22 VP.n4 161.3
R905 VP.n9 VP.t5 89.99
R906 VP.n19 VP.n18 80.6037
R907 VP.n34 VP.n33 80.6037
R908 VP.n21 VP.n20 80.6037
R909 VP.n21 VP.t2 69.0997
R910 VP.n33 VP.t0 69.0997
R911 VP.n18 VP.t4 69.0997
R912 VP.n9 VP.n8 42.1122
R913 VP.n27 VP.n26 40.4106
R914 VP.n28 VP.n27 40.4106
R915 VP.n13 VP.n12 40.4106
R916 VP.n12 VP.n11 40.4106
R917 VP.n22 VP.n21 40.1672
R918 VP.n33 VP.n32 40.1672
R919 VP.n18 VP.n17 40.1672
R920 VP.n3 VP.t3 38.0333
R921 VP.n1 VP.t1 38.0333
R922 VP.n6 VP.t6 38.0333
R923 VP.n8 VP.t7 38.0333
R924 VP.n20 VP.n19 37.3802
R925 VP.n23 VP.n22 29.6995
R926 VP.n32 VP.n31 29.6995
R927 VP.n17 VP.n16 29.6995
R928 VP.n10 VP.n9 28.9373
R929 VP.n26 VP.n3 14.85
R930 VP.n28 VP.n1 14.85
R931 VP.n13 VP.n6 14.85
R932 VP.n11 VP.n8 14.85
R933 VP.n23 VP.n3 9.49444
R934 VP.n31 VP.n1 9.49444
R935 VP.n16 VP.n6 9.49444
R936 VP.n19 VP.n5 0.285035
R937 VP.n20 VP.n4 0.285035
R938 VP.n34 VP.n0 0.285035
R939 VP.n10 VP.n7 0.189894
R940 VP.n14 VP.n7 0.189894
R941 VP.n15 VP.n14 0.189894
R942 VP.n15 VP.n5 0.189894
R943 VP.n24 VP.n4 0.189894
R944 VP.n25 VP.n24 0.189894
R945 VP.n25 VP.n2 0.189894
R946 VP.n29 VP.n2 0.189894
R947 VP.n30 VP.n29 0.189894
R948 VP.n30 VP.n0 0.189894
R949 VP VP.n34 0.146778
R950 VTAIL.n66 VTAIL.n64 289.615
R951 VTAIL.n4 VTAIL.n2 289.615
R952 VTAIL.n12 VTAIL.n10 289.615
R953 VTAIL.n22 VTAIL.n20 289.615
R954 VTAIL.n58 VTAIL.n56 289.615
R955 VTAIL.n48 VTAIL.n46 289.615
R956 VTAIL.n40 VTAIL.n38 289.615
R957 VTAIL.n30 VTAIL.n28 289.615
R958 VTAIL.n67 VTAIL.n66 185
R959 VTAIL.n5 VTAIL.n4 185
R960 VTAIL.n13 VTAIL.n12 185
R961 VTAIL.n23 VTAIL.n22 185
R962 VTAIL.n59 VTAIL.n58 185
R963 VTAIL.n49 VTAIL.n48 185
R964 VTAIL.n41 VTAIL.n40 185
R965 VTAIL.n31 VTAIL.n30 185
R966 VTAIL.t3 VTAIL.n65 167.117
R967 VTAIL.t6 VTAIL.n3 167.117
R968 VTAIL.t8 VTAIL.n11 167.117
R969 VTAIL.t12 VTAIL.n21 167.117
R970 VTAIL.t14 VTAIL.n57 167.117
R971 VTAIL.t9 VTAIL.n47 167.117
R972 VTAIL.t0 VTAIL.n39 167.117
R973 VTAIL.t2 VTAIL.n29 167.117
R974 VTAIL.n55 VTAIL.n54 84.5047
R975 VTAIL.n37 VTAIL.n36 84.5047
R976 VTAIL.n1 VTAIL.n0 84.5047
R977 VTAIL.n19 VTAIL.n18 84.5047
R978 VTAIL.n66 VTAIL.t3 52.3082
R979 VTAIL.n4 VTAIL.t6 52.3082
R980 VTAIL.n12 VTAIL.t8 52.3082
R981 VTAIL.n22 VTAIL.t12 52.3082
R982 VTAIL.n58 VTAIL.t14 52.3082
R983 VTAIL.n48 VTAIL.t9 52.3082
R984 VTAIL.n40 VTAIL.t0 52.3082
R985 VTAIL.n30 VTAIL.t2 52.3082
R986 VTAIL.n71 VTAIL.n70 31.7975
R987 VTAIL.n9 VTAIL.n8 31.7975
R988 VTAIL.n17 VTAIL.n16 31.7975
R989 VTAIL.n27 VTAIL.n26 31.7975
R990 VTAIL.n63 VTAIL.n62 31.7975
R991 VTAIL.n53 VTAIL.n52 31.7975
R992 VTAIL.n45 VTAIL.n44 31.7975
R993 VTAIL.n35 VTAIL.n34 31.7975
R994 VTAIL.n71 VTAIL.n63 15.4962
R995 VTAIL.n35 VTAIL.n27 15.4962
R996 VTAIL.n0 VTAIL.t7 9.80248
R997 VTAIL.n0 VTAIL.t5 9.80248
R998 VTAIL.n18 VTAIL.t11 9.80248
R999 VTAIL.n18 VTAIL.t13 9.80248
R1000 VTAIL.n54 VTAIL.t15 9.80248
R1001 VTAIL.n54 VTAIL.t10 9.80248
R1002 VTAIL.n36 VTAIL.t1 9.80248
R1003 VTAIL.n36 VTAIL.t4 9.80248
R1004 VTAIL.n67 VTAIL.n65 9.71174
R1005 VTAIL.n5 VTAIL.n3 9.71174
R1006 VTAIL.n13 VTAIL.n11 9.71174
R1007 VTAIL.n23 VTAIL.n21 9.71174
R1008 VTAIL.n59 VTAIL.n57 9.71174
R1009 VTAIL.n49 VTAIL.n47 9.71174
R1010 VTAIL.n41 VTAIL.n39 9.71174
R1011 VTAIL.n31 VTAIL.n29 9.71174
R1012 VTAIL.n70 VTAIL.n69 9.45567
R1013 VTAIL.n8 VTAIL.n7 9.45567
R1014 VTAIL.n16 VTAIL.n15 9.45567
R1015 VTAIL.n26 VTAIL.n25 9.45567
R1016 VTAIL.n62 VTAIL.n61 9.45567
R1017 VTAIL.n52 VTAIL.n51 9.45567
R1018 VTAIL.n44 VTAIL.n43 9.45567
R1019 VTAIL.n34 VTAIL.n33 9.45567
R1020 VTAIL.n69 VTAIL.n68 9.3005
R1021 VTAIL.n7 VTAIL.n6 9.3005
R1022 VTAIL.n15 VTAIL.n14 9.3005
R1023 VTAIL.n25 VTAIL.n24 9.3005
R1024 VTAIL.n61 VTAIL.n60 9.3005
R1025 VTAIL.n51 VTAIL.n50 9.3005
R1026 VTAIL.n43 VTAIL.n42 9.3005
R1027 VTAIL.n33 VTAIL.n32 9.3005
R1028 VTAIL.n70 VTAIL.n64 8.14595
R1029 VTAIL.n8 VTAIL.n2 8.14595
R1030 VTAIL.n16 VTAIL.n10 8.14595
R1031 VTAIL.n26 VTAIL.n20 8.14595
R1032 VTAIL.n62 VTAIL.n56 8.14595
R1033 VTAIL.n52 VTAIL.n46 8.14595
R1034 VTAIL.n44 VTAIL.n38 8.14595
R1035 VTAIL.n34 VTAIL.n28 8.14595
R1036 VTAIL.n68 VTAIL.n67 7.3702
R1037 VTAIL.n6 VTAIL.n5 7.3702
R1038 VTAIL.n14 VTAIL.n13 7.3702
R1039 VTAIL.n24 VTAIL.n23 7.3702
R1040 VTAIL.n60 VTAIL.n59 7.3702
R1041 VTAIL.n50 VTAIL.n49 7.3702
R1042 VTAIL.n42 VTAIL.n41 7.3702
R1043 VTAIL.n32 VTAIL.n31 7.3702
R1044 VTAIL.n68 VTAIL.n64 5.81868
R1045 VTAIL.n6 VTAIL.n2 5.81868
R1046 VTAIL.n14 VTAIL.n10 5.81868
R1047 VTAIL.n24 VTAIL.n20 5.81868
R1048 VTAIL.n60 VTAIL.n56 5.81868
R1049 VTAIL.n50 VTAIL.n46 5.81868
R1050 VTAIL.n42 VTAIL.n38 5.81868
R1051 VTAIL.n32 VTAIL.n28 5.81868
R1052 VTAIL.n69 VTAIL.n65 3.44771
R1053 VTAIL.n7 VTAIL.n3 3.44771
R1054 VTAIL.n15 VTAIL.n11 3.44771
R1055 VTAIL.n25 VTAIL.n21 3.44771
R1056 VTAIL.n61 VTAIL.n57 3.44771
R1057 VTAIL.n51 VTAIL.n47 3.44771
R1058 VTAIL.n43 VTAIL.n39 3.44771
R1059 VTAIL.n33 VTAIL.n29 3.44771
R1060 VTAIL.n37 VTAIL.n35 1.38843
R1061 VTAIL.n45 VTAIL.n37 1.38843
R1062 VTAIL.n55 VTAIL.n53 1.38843
R1063 VTAIL.n63 VTAIL.n55 1.38843
R1064 VTAIL.n27 VTAIL.n19 1.38843
R1065 VTAIL.n19 VTAIL.n17 1.38843
R1066 VTAIL.n9 VTAIL.n1 1.38843
R1067 VTAIL VTAIL.n71 1.33024
R1068 VTAIL.n53 VTAIL.n45 0.470328
R1069 VTAIL.n17 VTAIL.n9 0.470328
R1070 VTAIL VTAIL.n1 0.0586897
R1071 VDD1 VDD1.n0 101.936
R1072 VDD1.n3 VDD1.n2 101.823
R1073 VDD1.n3 VDD1.n1 101.823
R1074 VDD1.n5 VDD1.n4 101.183
R1075 VDD1.n5 VDD1.n3 32.2854
R1076 VDD1.n4 VDD1.t1 9.80248
R1077 VDD1.n4 VDD1.t3 9.80248
R1078 VDD1.n0 VDD1.t2 9.80248
R1079 VDD1.n0 VDD1.t0 9.80248
R1080 VDD1.n2 VDD1.t6 9.80248
R1081 VDD1.n2 VDD1.t7 9.80248
R1082 VDD1.n1 VDD1.t5 9.80248
R1083 VDD1.n1 VDD1.t4 9.80248
R1084 VDD1 VDD1.n5 0.636276
R1085 VN.n27 VN.n15 161.3
R1086 VN.n26 VN.n25 161.3
R1087 VN.n24 VN.n23 161.3
R1088 VN.n22 VN.n17 161.3
R1089 VN.n21 VN.n20 161.3
R1090 VN.n12 VN.n0 161.3
R1091 VN.n11 VN.n10 161.3
R1092 VN.n9 VN.n8 161.3
R1093 VN.n7 VN.n2 161.3
R1094 VN.n6 VN.n5 161.3
R1095 VN.n4 VN.t7 89.99
R1096 VN.n19 VN.t4 89.99
R1097 VN.n29 VN.n28 80.6037
R1098 VN.n14 VN.n13 80.6037
R1099 VN.n13 VN.t2 69.0997
R1100 VN.n28 VN.t5 69.0997
R1101 VN.n4 VN.n3 42.1122
R1102 VN.n19 VN.n18 42.1122
R1103 VN.n7 VN.n6 40.4106
R1104 VN.n8 VN.n7 40.4106
R1105 VN.n22 VN.n21 40.4106
R1106 VN.n23 VN.n22 40.4106
R1107 VN.n13 VN.n12 40.1672
R1108 VN.n28 VN.n27 40.1672
R1109 VN.n3 VN.t6 38.0333
R1110 VN.n1 VN.t0 38.0333
R1111 VN.n18 VN.t3 38.0333
R1112 VN.n16 VN.t1 38.0333
R1113 VN VN.n29 37.6657
R1114 VN.n12 VN.n11 29.6995
R1115 VN.n27 VN.n26 29.6995
R1116 VN.n20 VN.n19 28.9373
R1117 VN.n5 VN.n4 28.9373
R1118 VN.n6 VN.n3 14.85
R1119 VN.n8 VN.n1 14.85
R1120 VN.n21 VN.n18 14.85
R1121 VN.n23 VN.n16 14.85
R1122 VN.n11 VN.n1 9.49444
R1123 VN.n26 VN.n16 9.49444
R1124 VN.n29 VN.n15 0.285035
R1125 VN.n14 VN.n0 0.285035
R1126 VN.n25 VN.n15 0.189894
R1127 VN.n25 VN.n24 0.189894
R1128 VN.n24 VN.n17 0.189894
R1129 VN.n20 VN.n17 0.189894
R1130 VN.n5 VN.n2 0.189894
R1131 VN.n9 VN.n2 0.189894
R1132 VN.n10 VN.n9 0.189894
R1133 VN.n10 VN.n0 0.189894
R1134 VN VN.n14 0.146778
R1135 VDD2.n2 VDD2.n1 101.823
R1136 VDD2.n2 VDD2.n0 101.823
R1137 VDD2 VDD2.n5 101.82
R1138 VDD2.n4 VDD2.n3 101.183
R1139 VDD2.n4 VDD2.n2 31.7024
R1140 VDD2.n5 VDD2.t4 9.80248
R1141 VDD2.n5 VDD2.t3 9.80248
R1142 VDD2.n3 VDD2.t2 9.80248
R1143 VDD2.n3 VDD2.t6 9.80248
R1144 VDD2.n1 VDD2.t7 9.80248
R1145 VDD2.n1 VDD2.t5 9.80248
R1146 VDD2.n0 VDD2.t0 9.80248
R1147 VDD2.n0 VDD2.t1 9.80248
R1148 VDD2 VDD2.n4 0.752655
C0 VDD1 VDD2 1.11609f
C1 VN VP 4.20783f
C2 VTAIL VP 2.1023f
C3 VN VDD2 1.55309f
C4 VTAIL VDD2 3.76958f
C5 VDD1 VN 0.154658f
C6 VDD1 VTAIL 3.72401f
C7 VTAIL VN 2.08819f
C8 VDD2 VP 0.385382f
C9 VDD1 VP 1.78213f
C10 VDD2 B 3.106872f
C11 VDD1 B 3.383143f
C12 VTAIL B 3.403431f
C13 VN B 9.27939f
C14 VP B 8.045511f
C15 VDD2.t0 B 0.028166f
C16 VDD2.t1 B 0.028166f
C17 VDD2.n0 B 0.178748f
C18 VDD2.t7 B 0.028166f
C19 VDD2.t5 B 0.028166f
C20 VDD2.n1 B 0.178748f
C21 VDD2.n2 B 1.33598f
C22 VDD2.t2 B 0.028166f
C23 VDD2.t6 B 0.028166f
C24 VDD2.n3 B 0.177126f
C25 VDD2.n4 B 1.19009f
C26 VDD2.t4 B 0.028166f
C27 VDD2.t3 B 0.028166f
C28 VDD2.n5 B 0.178736f
C29 VN.n0 B 0.042356f
C30 VN.t0 B 0.192052f
C31 VN.n1 B 0.106025f
C32 VN.n2 B 0.031742f
C33 VN.t6 B 0.192052f
C34 VN.n3 B 0.150537f
C35 VN.t7 B 0.296114f
C36 VN.n4 B 0.159565f
C37 VN.n5 B 0.169081f
C38 VN.n6 B 0.051976f
C39 VN.n7 B 0.025687f
C40 VN.n8 B 0.051976f
C41 VN.n9 B 0.031742f
C42 VN.n10 B 0.031742f
C43 VN.n11 B 0.045678f
C44 VN.n12 B 0.027048f
C45 VN.t2 B 0.254678f
C46 VN.n13 B 0.171217f
C47 VN.n14 B 0.029728f
C48 VN.n15 B 0.042356f
C49 VN.t1 B 0.192052f
C50 VN.n16 B 0.106025f
C51 VN.n17 B 0.031742f
C52 VN.t3 B 0.192052f
C53 VN.n18 B 0.150537f
C54 VN.t4 B 0.296114f
C55 VN.n19 B 0.159565f
C56 VN.n20 B 0.169081f
C57 VN.n21 B 0.051976f
C58 VN.n22 B 0.025687f
C59 VN.n23 B 0.051976f
C60 VN.n24 B 0.031742f
C61 VN.n25 B 0.031742f
C62 VN.n26 B 0.045678f
C63 VN.n27 B 0.027048f
C64 VN.t5 B 0.254678f
C65 VN.n28 B 0.171217f
C66 VN.n29 B 1.0994f
C67 VDD1.t2 B 0.026962f
C68 VDD1.t0 B 0.026962f
C69 VDD1.n0 B 0.171425f
C70 VDD1.t5 B 0.026962f
C71 VDD1.t4 B 0.026962f
C72 VDD1.n1 B 0.171109f
C73 VDD1.t6 B 0.026962f
C74 VDD1.t7 B 0.026962f
C75 VDD1.n2 B 0.171109f
C76 VDD1.n3 B 1.31479f
C77 VDD1.t1 B 0.026962f
C78 VDD1.t3 B 0.026962f
C79 VDD1.n4 B 0.169557f
C80 VDD1.n5 B 1.15939f
C81 VTAIL.t7 B 0.044856f
C82 VTAIL.t5 B 0.044856f
C83 VTAIL.n0 B 0.240458f
C84 VTAIL.n1 B 0.350596f
C85 VTAIL.n2 B 0.041393f
C86 VTAIL.n3 B 0.091458f
C87 VTAIL.t6 B 0.068579f
C88 VTAIL.n4 B 0.071694f
C89 VTAIL.n5 B 0.022895f
C90 VTAIL.n6 B 0.0151f
C91 VTAIL.n7 B 0.202333f
C92 VTAIL.n8 B 0.045429f
C93 VTAIL.n9 B 0.191778f
C94 VTAIL.n10 B 0.041393f
C95 VTAIL.n11 B 0.091458f
C96 VTAIL.t8 B 0.068579f
C97 VTAIL.n12 B 0.071694f
C98 VTAIL.n13 B 0.022895f
C99 VTAIL.n14 B 0.0151f
C100 VTAIL.n15 B 0.202333f
C101 VTAIL.n16 B 0.045429f
C102 VTAIL.n17 B 0.191778f
C103 VTAIL.t11 B 0.044856f
C104 VTAIL.t13 B 0.044856f
C105 VTAIL.n18 B 0.240458f
C106 VTAIL.n19 B 0.470998f
C107 VTAIL.n20 B 0.041393f
C108 VTAIL.n21 B 0.091458f
C109 VTAIL.t12 B 0.068579f
C110 VTAIL.n22 B 0.071694f
C111 VTAIL.n23 B 0.022895f
C112 VTAIL.n24 B 0.0151f
C113 VTAIL.n25 B 0.202333f
C114 VTAIL.n26 B 0.045429f
C115 VTAIL.n27 B 0.814291f
C116 VTAIL.n28 B 0.041393f
C117 VTAIL.n29 B 0.091458f
C118 VTAIL.t2 B 0.068579f
C119 VTAIL.n30 B 0.071694f
C120 VTAIL.n31 B 0.022895f
C121 VTAIL.n32 B 0.0151f
C122 VTAIL.n33 B 0.202333f
C123 VTAIL.n34 B 0.045429f
C124 VTAIL.n35 B 0.814291f
C125 VTAIL.t1 B 0.044856f
C126 VTAIL.t4 B 0.044856f
C127 VTAIL.n36 B 0.24046f
C128 VTAIL.n37 B 0.470997f
C129 VTAIL.n38 B 0.041393f
C130 VTAIL.n39 B 0.091458f
C131 VTAIL.t0 B 0.068579f
C132 VTAIL.n40 B 0.071694f
C133 VTAIL.n41 B 0.022895f
C134 VTAIL.n42 B 0.0151f
C135 VTAIL.n43 B 0.202333f
C136 VTAIL.n44 B 0.045429f
C137 VTAIL.n45 B 0.191778f
C138 VTAIL.n46 B 0.041393f
C139 VTAIL.n47 B 0.091458f
C140 VTAIL.t9 B 0.068579f
C141 VTAIL.n48 B 0.071694f
C142 VTAIL.n49 B 0.022895f
C143 VTAIL.n50 B 0.0151f
C144 VTAIL.n51 B 0.202333f
C145 VTAIL.n52 B 0.045429f
C146 VTAIL.n53 B 0.191778f
C147 VTAIL.t15 B 0.044856f
C148 VTAIL.t10 B 0.044856f
C149 VTAIL.n54 B 0.24046f
C150 VTAIL.n55 B 0.470997f
C151 VTAIL.n56 B 0.041393f
C152 VTAIL.n57 B 0.091458f
C153 VTAIL.t14 B 0.068579f
C154 VTAIL.n58 B 0.071694f
C155 VTAIL.n59 B 0.022895f
C156 VTAIL.n60 B 0.0151f
C157 VTAIL.n61 B 0.202333f
C158 VTAIL.n62 B 0.045429f
C159 VTAIL.n63 B 0.814291f
C160 VTAIL.n64 B 0.041393f
C161 VTAIL.n65 B 0.091458f
C162 VTAIL.t3 B 0.068579f
C163 VTAIL.n66 B 0.071694f
C164 VTAIL.n67 B 0.022895f
C165 VTAIL.n68 B 0.0151f
C166 VTAIL.n69 B 0.202333f
C167 VTAIL.n70 B 0.045429f
C168 VTAIL.n71 B 0.809022f
C169 VP.n0 B 0.042658f
C170 VP.t1 B 0.193422f
C171 VP.n1 B 0.106781f
C172 VP.n2 B 0.031969f
C173 VP.t3 B 0.193422f
C174 VP.n3 B 0.106781f
C175 VP.n4 B 0.042658f
C176 VP.n5 B 0.042658f
C177 VP.t4 B 0.256495f
C178 VP.t6 B 0.193422f
C179 VP.n6 B 0.106781f
C180 VP.n7 B 0.031969f
C181 VP.t7 B 0.193422f
C182 VP.n8 B 0.151611f
C183 VP.t5 B 0.298226f
C184 VP.n9 B 0.160703f
C185 VP.n10 B 0.170287f
C186 VP.n11 B 0.052347f
C187 VP.n12 B 0.02587f
C188 VP.n13 B 0.052347f
C189 VP.n14 B 0.031969f
C190 VP.n15 B 0.031969f
C191 VP.n16 B 0.046004f
C192 VP.n17 B 0.027241f
C193 VP.n18 B 0.172438f
C194 VP.n19 B 1.08891f
C195 VP.n20 B 1.11957f
C196 VP.t2 B 0.256495f
C197 VP.n21 B 0.172438f
C198 VP.n22 B 0.027241f
C199 VP.n23 B 0.046004f
C200 VP.n24 B 0.031969f
C201 VP.n25 B 0.031969f
C202 VP.n26 B 0.052347f
C203 VP.n27 B 0.02587f
C204 VP.n28 B 0.052347f
C205 VP.n29 B 0.031969f
C206 VP.n30 B 0.031969f
C207 VP.n31 B 0.046004f
C208 VP.n32 B 0.027241f
C209 VP.t0 B 0.256495f
C210 VP.n33 B 0.172438f
C211 VP.n34 B 0.02994f
.ends

