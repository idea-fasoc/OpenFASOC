* NGSPICE file created from diff_pair_sample_1596.ext - technology: sky130A

.subckt diff_pair_sample_1596 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=5.7135 pd=30.08 as=0 ps=0 w=14.65 l=0.91
X1 VDD2.t5 VN.t0 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=2.41725 pd=14.98 as=5.7135 ps=30.08 w=14.65 l=0.91
X2 VDD2.t4 VN.t1 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=5.7135 pd=30.08 as=2.41725 ps=14.98 w=14.65 l=0.91
X3 VDD1.t5 VP.t0 VTAIL.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=2.41725 pd=14.98 as=5.7135 ps=30.08 w=14.65 l=0.91
X4 VDD1.t4 VP.t1 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=5.7135 pd=30.08 as=2.41725 ps=14.98 w=14.65 l=0.91
X5 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=5.7135 pd=30.08 as=0 ps=0 w=14.65 l=0.91
X6 VTAIL.t7 VN.t2 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=2.41725 pd=14.98 as=2.41725 ps=14.98 w=14.65 l=0.91
X7 VTAIL.t8 VN.t3 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.41725 pd=14.98 as=2.41725 ps=14.98 w=14.65 l=0.91
X8 VTAIL.t1 VP.t2 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=2.41725 pd=14.98 as=2.41725 ps=14.98 w=14.65 l=0.91
X9 VDD2.t1 VN.t4 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=5.7135 pd=30.08 as=2.41725 ps=14.98 w=14.65 l=0.91
X10 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.7135 pd=30.08 as=0 ps=0 w=14.65 l=0.91
X11 VTAIL.t0 VP.t3 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.41725 pd=14.98 as=2.41725 ps=14.98 w=14.65 l=0.91
X12 VDD1.t1 VP.t4 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.41725 pd=14.98 as=5.7135 ps=30.08 w=14.65 l=0.91
X13 VDD2.t0 VN.t5 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=2.41725 pd=14.98 as=5.7135 ps=30.08 w=14.65 l=0.91
X14 VDD1.t0 VP.t5 VTAIL.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=5.7135 pd=30.08 as=2.41725 ps=14.98 w=14.65 l=0.91
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.7135 pd=30.08 as=0 ps=0 w=14.65 l=0.91
R0 B.n70 B.t6 590.259
R1 B.n78 B.t14 590.259
R2 B.n177 B.t10 590.259
R3 B.n169 B.t17 590.259
R4 B.n518 B.n517 585
R5 B.n520 B.n103 585
R6 B.n523 B.n522 585
R7 B.n524 B.n102 585
R8 B.n526 B.n525 585
R9 B.n528 B.n101 585
R10 B.n531 B.n530 585
R11 B.n532 B.n100 585
R12 B.n534 B.n533 585
R13 B.n536 B.n99 585
R14 B.n539 B.n538 585
R15 B.n540 B.n98 585
R16 B.n542 B.n541 585
R17 B.n544 B.n97 585
R18 B.n547 B.n546 585
R19 B.n548 B.n96 585
R20 B.n550 B.n549 585
R21 B.n552 B.n95 585
R22 B.n555 B.n554 585
R23 B.n556 B.n94 585
R24 B.n558 B.n557 585
R25 B.n560 B.n93 585
R26 B.n563 B.n562 585
R27 B.n564 B.n92 585
R28 B.n566 B.n565 585
R29 B.n568 B.n91 585
R30 B.n571 B.n570 585
R31 B.n572 B.n90 585
R32 B.n574 B.n573 585
R33 B.n576 B.n89 585
R34 B.n579 B.n578 585
R35 B.n580 B.n88 585
R36 B.n582 B.n581 585
R37 B.n584 B.n87 585
R38 B.n587 B.n586 585
R39 B.n588 B.n86 585
R40 B.n590 B.n589 585
R41 B.n592 B.n85 585
R42 B.n595 B.n594 585
R43 B.n596 B.n84 585
R44 B.n598 B.n597 585
R45 B.n600 B.n83 585
R46 B.n603 B.n602 585
R47 B.n604 B.n82 585
R48 B.n606 B.n605 585
R49 B.n608 B.n81 585
R50 B.n611 B.n610 585
R51 B.n612 B.n77 585
R52 B.n614 B.n613 585
R53 B.n616 B.n76 585
R54 B.n619 B.n618 585
R55 B.n620 B.n75 585
R56 B.n622 B.n621 585
R57 B.n624 B.n74 585
R58 B.n627 B.n626 585
R59 B.n628 B.n73 585
R60 B.n630 B.n629 585
R61 B.n632 B.n72 585
R62 B.n635 B.n634 585
R63 B.n637 B.n69 585
R64 B.n639 B.n638 585
R65 B.n641 B.n68 585
R66 B.n644 B.n643 585
R67 B.n645 B.n67 585
R68 B.n647 B.n646 585
R69 B.n649 B.n66 585
R70 B.n652 B.n651 585
R71 B.n653 B.n65 585
R72 B.n655 B.n654 585
R73 B.n657 B.n64 585
R74 B.n660 B.n659 585
R75 B.n661 B.n63 585
R76 B.n663 B.n662 585
R77 B.n665 B.n62 585
R78 B.n668 B.n667 585
R79 B.n669 B.n61 585
R80 B.n671 B.n670 585
R81 B.n673 B.n60 585
R82 B.n676 B.n675 585
R83 B.n677 B.n59 585
R84 B.n679 B.n678 585
R85 B.n681 B.n58 585
R86 B.n684 B.n683 585
R87 B.n685 B.n57 585
R88 B.n687 B.n686 585
R89 B.n689 B.n56 585
R90 B.n692 B.n691 585
R91 B.n693 B.n55 585
R92 B.n695 B.n694 585
R93 B.n697 B.n54 585
R94 B.n700 B.n699 585
R95 B.n701 B.n53 585
R96 B.n703 B.n702 585
R97 B.n705 B.n52 585
R98 B.n708 B.n707 585
R99 B.n709 B.n51 585
R100 B.n711 B.n710 585
R101 B.n713 B.n50 585
R102 B.n716 B.n715 585
R103 B.n717 B.n49 585
R104 B.n719 B.n718 585
R105 B.n721 B.n48 585
R106 B.n724 B.n723 585
R107 B.n725 B.n47 585
R108 B.n727 B.n726 585
R109 B.n729 B.n46 585
R110 B.n732 B.n731 585
R111 B.n733 B.n45 585
R112 B.n516 B.n43 585
R113 B.n736 B.n43 585
R114 B.n515 B.n42 585
R115 B.n737 B.n42 585
R116 B.n514 B.n41 585
R117 B.n738 B.n41 585
R118 B.n513 B.n512 585
R119 B.n512 B.n37 585
R120 B.n511 B.n36 585
R121 B.n744 B.n36 585
R122 B.n510 B.n35 585
R123 B.n745 B.n35 585
R124 B.n509 B.n34 585
R125 B.n746 B.n34 585
R126 B.n508 B.n507 585
R127 B.n507 B.n30 585
R128 B.n506 B.n29 585
R129 B.n752 B.n29 585
R130 B.n505 B.n28 585
R131 B.n753 B.n28 585
R132 B.n504 B.n27 585
R133 B.n754 B.n27 585
R134 B.n503 B.n502 585
R135 B.n502 B.n26 585
R136 B.n501 B.n22 585
R137 B.n760 B.n22 585
R138 B.n500 B.n21 585
R139 B.n761 B.n21 585
R140 B.n499 B.n20 585
R141 B.n762 B.n20 585
R142 B.n498 B.n497 585
R143 B.n497 B.n19 585
R144 B.n496 B.n15 585
R145 B.n768 B.n15 585
R146 B.n495 B.n14 585
R147 B.n769 B.n14 585
R148 B.n494 B.n13 585
R149 B.n770 B.n13 585
R150 B.n493 B.n492 585
R151 B.n492 B.n12 585
R152 B.n491 B.n490 585
R153 B.n491 B.n8 585
R154 B.n489 B.n7 585
R155 B.n777 B.n7 585
R156 B.n488 B.n6 585
R157 B.n778 B.n6 585
R158 B.n487 B.n5 585
R159 B.n779 B.n5 585
R160 B.n486 B.n485 585
R161 B.n485 B.n4 585
R162 B.n484 B.n104 585
R163 B.n484 B.n483 585
R164 B.n473 B.n105 585
R165 B.n476 B.n105 585
R166 B.n475 B.n474 585
R167 B.n477 B.n475 585
R168 B.n472 B.n110 585
R169 B.n110 B.n109 585
R170 B.n471 B.n470 585
R171 B.n470 B.n469 585
R172 B.n112 B.n111 585
R173 B.n462 B.n112 585
R174 B.n461 B.n460 585
R175 B.n463 B.n461 585
R176 B.n459 B.n117 585
R177 B.n117 B.n116 585
R178 B.n458 B.n457 585
R179 B.n457 B.n456 585
R180 B.n119 B.n118 585
R181 B.n449 B.n119 585
R182 B.n448 B.n447 585
R183 B.n450 B.n448 585
R184 B.n446 B.n124 585
R185 B.n124 B.n123 585
R186 B.n445 B.n444 585
R187 B.n444 B.n443 585
R188 B.n126 B.n125 585
R189 B.n127 B.n126 585
R190 B.n436 B.n435 585
R191 B.n437 B.n436 585
R192 B.n434 B.n132 585
R193 B.n132 B.n131 585
R194 B.n433 B.n432 585
R195 B.n432 B.n431 585
R196 B.n134 B.n133 585
R197 B.n135 B.n134 585
R198 B.n424 B.n423 585
R199 B.n425 B.n424 585
R200 B.n422 B.n140 585
R201 B.n140 B.n139 585
R202 B.n421 B.n420 585
R203 B.n420 B.n419 585
R204 B.n416 B.n144 585
R205 B.n415 B.n414 585
R206 B.n412 B.n145 585
R207 B.n412 B.n143 585
R208 B.n411 B.n410 585
R209 B.n409 B.n408 585
R210 B.n407 B.n147 585
R211 B.n405 B.n404 585
R212 B.n403 B.n148 585
R213 B.n402 B.n401 585
R214 B.n399 B.n149 585
R215 B.n397 B.n396 585
R216 B.n395 B.n150 585
R217 B.n394 B.n393 585
R218 B.n391 B.n151 585
R219 B.n389 B.n388 585
R220 B.n387 B.n152 585
R221 B.n386 B.n385 585
R222 B.n383 B.n153 585
R223 B.n381 B.n380 585
R224 B.n379 B.n154 585
R225 B.n378 B.n377 585
R226 B.n375 B.n155 585
R227 B.n373 B.n372 585
R228 B.n371 B.n156 585
R229 B.n370 B.n369 585
R230 B.n367 B.n157 585
R231 B.n365 B.n364 585
R232 B.n363 B.n158 585
R233 B.n362 B.n361 585
R234 B.n359 B.n159 585
R235 B.n357 B.n356 585
R236 B.n355 B.n160 585
R237 B.n354 B.n353 585
R238 B.n351 B.n161 585
R239 B.n349 B.n348 585
R240 B.n347 B.n162 585
R241 B.n346 B.n345 585
R242 B.n343 B.n163 585
R243 B.n341 B.n340 585
R244 B.n339 B.n164 585
R245 B.n338 B.n337 585
R246 B.n335 B.n165 585
R247 B.n333 B.n332 585
R248 B.n331 B.n166 585
R249 B.n330 B.n329 585
R250 B.n327 B.n167 585
R251 B.n325 B.n324 585
R252 B.n323 B.n168 585
R253 B.n322 B.n321 585
R254 B.n319 B.n318 585
R255 B.n317 B.n316 585
R256 B.n315 B.n173 585
R257 B.n313 B.n312 585
R258 B.n311 B.n174 585
R259 B.n310 B.n309 585
R260 B.n307 B.n175 585
R261 B.n305 B.n304 585
R262 B.n303 B.n176 585
R263 B.n302 B.n301 585
R264 B.n299 B.n298 585
R265 B.n297 B.n296 585
R266 B.n295 B.n181 585
R267 B.n293 B.n292 585
R268 B.n291 B.n182 585
R269 B.n290 B.n289 585
R270 B.n287 B.n183 585
R271 B.n285 B.n284 585
R272 B.n283 B.n184 585
R273 B.n282 B.n281 585
R274 B.n279 B.n185 585
R275 B.n277 B.n276 585
R276 B.n275 B.n186 585
R277 B.n274 B.n273 585
R278 B.n271 B.n187 585
R279 B.n269 B.n268 585
R280 B.n267 B.n188 585
R281 B.n266 B.n265 585
R282 B.n263 B.n189 585
R283 B.n261 B.n260 585
R284 B.n259 B.n190 585
R285 B.n258 B.n257 585
R286 B.n255 B.n191 585
R287 B.n253 B.n252 585
R288 B.n251 B.n192 585
R289 B.n250 B.n249 585
R290 B.n247 B.n193 585
R291 B.n245 B.n244 585
R292 B.n243 B.n194 585
R293 B.n242 B.n241 585
R294 B.n239 B.n195 585
R295 B.n237 B.n236 585
R296 B.n235 B.n196 585
R297 B.n234 B.n233 585
R298 B.n231 B.n197 585
R299 B.n229 B.n228 585
R300 B.n227 B.n198 585
R301 B.n226 B.n225 585
R302 B.n223 B.n199 585
R303 B.n221 B.n220 585
R304 B.n219 B.n200 585
R305 B.n218 B.n217 585
R306 B.n215 B.n201 585
R307 B.n213 B.n212 585
R308 B.n211 B.n202 585
R309 B.n210 B.n209 585
R310 B.n207 B.n203 585
R311 B.n205 B.n204 585
R312 B.n142 B.n141 585
R313 B.n143 B.n142 585
R314 B.n418 B.n417 585
R315 B.n419 B.n418 585
R316 B.n138 B.n137 585
R317 B.n139 B.n138 585
R318 B.n427 B.n426 585
R319 B.n426 B.n425 585
R320 B.n428 B.n136 585
R321 B.n136 B.n135 585
R322 B.n430 B.n429 585
R323 B.n431 B.n430 585
R324 B.n130 B.n129 585
R325 B.n131 B.n130 585
R326 B.n439 B.n438 585
R327 B.n438 B.n437 585
R328 B.n440 B.n128 585
R329 B.n128 B.n127 585
R330 B.n442 B.n441 585
R331 B.n443 B.n442 585
R332 B.n122 B.n121 585
R333 B.n123 B.n122 585
R334 B.n452 B.n451 585
R335 B.n451 B.n450 585
R336 B.n453 B.n120 585
R337 B.n449 B.n120 585
R338 B.n455 B.n454 585
R339 B.n456 B.n455 585
R340 B.n115 B.n114 585
R341 B.n116 B.n115 585
R342 B.n465 B.n464 585
R343 B.n464 B.n463 585
R344 B.n466 B.n113 585
R345 B.n462 B.n113 585
R346 B.n468 B.n467 585
R347 B.n469 B.n468 585
R348 B.n108 B.n107 585
R349 B.n109 B.n108 585
R350 B.n479 B.n478 585
R351 B.n478 B.n477 585
R352 B.n480 B.n106 585
R353 B.n476 B.n106 585
R354 B.n482 B.n481 585
R355 B.n483 B.n482 585
R356 B.n3 B.n0 585
R357 B.n4 B.n3 585
R358 B.n776 B.n1 585
R359 B.n777 B.n776 585
R360 B.n775 B.n774 585
R361 B.n775 B.n8 585
R362 B.n773 B.n9 585
R363 B.n12 B.n9 585
R364 B.n772 B.n771 585
R365 B.n771 B.n770 585
R366 B.n11 B.n10 585
R367 B.n769 B.n11 585
R368 B.n767 B.n766 585
R369 B.n768 B.n767 585
R370 B.n765 B.n16 585
R371 B.n19 B.n16 585
R372 B.n764 B.n763 585
R373 B.n763 B.n762 585
R374 B.n18 B.n17 585
R375 B.n761 B.n18 585
R376 B.n759 B.n758 585
R377 B.n760 B.n759 585
R378 B.n757 B.n23 585
R379 B.n26 B.n23 585
R380 B.n756 B.n755 585
R381 B.n755 B.n754 585
R382 B.n25 B.n24 585
R383 B.n753 B.n25 585
R384 B.n751 B.n750 585
R385 B.n752 B.n751 585
R386 B.n749 B.n31 585
R387 B.n31 B.n30 585
R388 B.n748 B.n747 585
R389 B.n747 B.n746 585
R390 B.n33 B.n32 585
R391 B.n745 B.n33 585
R392 B.n743 B.n742 585
R393 B.n744 B.n743 585
R394 B.n741 B.n38 585
R395 B.n38 B.n37 585
R396 B.n740 B.n739 585
R397 B.n739 B.n738 585
R398 B.n40 B.n39 585
R399 B.n737 B.n40 585
R400 B.n735 B.n734 585
R401 B.n736 B.n735 585
R402 B.n780 B.n779 585
R403 B.n778 B.n2 585
R404 B.n735 B.n45 564.573
R405 B.n518 B.n43 564.573
R406 B.n420 B.n142 564.573
R407 B.n418 B.n144 564.573
R408 B.n78 B.t15 351.548
R409 B.n177 B.t13 351.548
R410 B.n70 B.t8 351.548
R411 B.n169 B.t19 351.548
R412 B.n79 B.t16 327.5
R413 B.n178 B.t12 327.5
R414 B.n71 B.t9 327.5
R415 B.n170 B.t18 327.5
R416 B.n519 B.n44 256.663
R417 B.n521 B.n44 256.663
R418 B.n527 B.n44 256.663
R419 B.n529 B.n44 256.663
R420 B.n535 B.n44 256.663
R421 B.n537 B.n44 256.663
R422 B.n543 B.n44 256.663
R423 B.n545 B.n44 256.663
R424 B.n551 B.n44 256.663
R425 B.n553 B.n44 256.663
R426 B.n559 B.n44 256.663
R427 B.n561 B.n44 256.663
R428 B.n567 B.n44 256.663
R429 B.n569 B.n44 256.663
R430 B.n575 B.n44 256.663
R431 B.n577 B.n44 256.663
R432 B.n583 B.n44 256.663
R433 B.n585 B.n44 256.663
R434 B.n591 B.n44 256.663
R435 B.n593 B.n44 256.663
R436 B.n599 B.n44 256.663
R437 B.n601 B.n44 256.663
R438 B.n607 B.n44 256.663
R439 B.n609 B.n44 256.663
R440 B.n615 B.n44 256.663
R441 B.n617 B.n44 256.663
R442 B.n623 B.n44 256.663
R443 B.n625 B.n44 256.663
R444 B.n631 B.n44 256.663
R445 B.n633 B.n44 256.663
R446 B.n640 B.n44 256.663
R447 B.n642 B.n44 256.663
R448 B.n648 B.n44 256.663
R449 B.n650 B.n44 256.663
R450 B.n656 B.n44 256.663
R451 B.n658 B.n44 256.663
R452 B.n664 B.n44 256.663
R453 B.n666 B.n44 256.663
R454 B.n672 B.n44 256.663
R455 B.n674 B.n44 256.663
R456 B.n680 B.n44 256.663
R457 B.n682 B.n44 256.663
R458 B.n688 B.n44 256.663
R459 B.n690 B.n44 256.663
R460 B.n696 B.n44 256.663
R461 B.n698 B.n44 256.663
R462 B.n704 B.n44 256.663
R463 B.n706 B.n44 256.663
R464 B.n712 B.n44 256.663
R465 B.n714 B.n44 256.663
R466 B.n720 B.n44 256.663
R467 B.n722 B.n44 256.663
R468 B.n728 B.n44 256.663
R469 B.n730 B.n44 256.663
R470 B.n413 B.n143 256.663
R471 B.n146 B.n143 256.663
R472 B.n406 B.n143 256.663
R473 B.n400 B.n143 256.663
R474 B.n398 B.n143 256.663
R475 B.n392 B.n143 256.663
R476 B.n390 B.n143 256.663
R477 B.n384 B.n143 256.663
R478 B.n382 B.n143 256.663
R479 B.n376 B.n143 256.663
R480 B.n374 B.n143 256.663
R481 B.n368 B.n143 256.663
R482 B.n366 B.n143 256.663
R483 B.n360 B.n143 256.663
R484 B.n358 B.n143 256.663
R485 B.n352 B.n143 256.663
R486 B.n350 B.n143 256.663
R487 B.n344 B.n143 256.663
R488 B.n342 B.n143 256.663
R489 B.n336 B.n143 256.663
R490 B.n334 B.n143 256.663
R491 B.n328 B.n143 256.663
R492 B.n326 B.n143 256.663
R493 B.n320 B.n143 256.663
R494 B.n172 B.n143 256.663
R495 B.n314 B.n143 256.663
R496 B.n308 B.n143 256.663
R497 B.n306 B.n143 256.663
R498 B.n300 B.n143 256.663
R499 B.n180 B.n143 256.663
R500 B.n294 B.n143 256.663
R501 B.n288 B.n143 256.663
R502 B.n286 B.n143 256.663
R503 B.n280 B.n143 256.663
R504 B.n278 B.n143 256.663
R505 B.n272 B.n143 256.663
R506 B.n270 B.n143 256.663
R507 B.n264 B.n143 256.663
R508 B.n262 B.n143 256.663
R509 B.n256 B.n143 256.663
R510 B.n254 B.n143 256.663
R511 B.n248 B.n143 256.663
R512 B.n246 B.n143 256.663
R513 B.n240 B.n143 256.663
R514 B.n238 B.n143 256.663
R515 B.n232 B.n143 256.663
R516 B.n230 B.n143 256.663
R517 B.n224 B.n143 256.663
R518 B.n222 B.n143 256.663
R519 B.n216 B.n143 256.663
R520 B.n214 B.n143 256.663
R521 B.n208 B.n143 256.663
R522 B.n206 B.n143 256.663
R523 B.n782 B.n781 256.663
R524 B.n731 B.n729 163.367
R525 B.n727 B.n47 163.367
R526 B.n723 B.n721 163.367
R527 B.n719 B.n49 163.367
R528 B.n715 B.n713 163.367
R529 B.n711 B.n51 163.367
R530 B.n707 B.n705 163.367
R531 B.n703 B.n53 163.367
R532 B.n699 B.n697 163.367
R533 B.n695 B.n55 163.367
R534 B.n691 B.n689 163.367
R535 B.n687 B.n57 163.367
R536 B.n683 B.n681 163.367
R537 B.n679 B.n59 163.367
R538 B.n675 B.n673 163.367
R539 B.n671 B.n61 163.367
R540 B.n667 B.n665 163.367
R541 B.n663 B.n63 163.367
R542 B.n659 B.n657 163.367
R543 B.n655 B.n65 163.367
R544 B.n651 B.n649 163.367
R545 B.n647 B.n67 163.367
R546 B.n643 B.n641 163.367
R547 B.n639 B.n69 163.367
R548 B.n634 B.n632 163.367
R549 B.n630 B.n73 163.367
R550 B.n626 B.n624 163.367
R551 B.n622 B.n75 163.367
R552 B.n618 B.n616 163.367
R553 B.n614 B.n77 163.367
R554 B.n610 B.n608 163.367
R555 B.n606 B.n82 163.367
R556 B.n602 B.n600 163.367
R557 B.n598 B.n84 163.367
R558 B.n594 B.n592 163.367
R559 B.n590 B.n86 163.367
R560 B.n586 B.n584 163.367
R561 B.n582 B.n88 163.367
R562 B.n578 B.n576 163.367
R563 B.n574 B.n90 163.367
R564 B.n570 B.n568 163.367
R565 B.n566 B.n92 163.367
R566 B.n562 B.n560 163.367
R567 B.n558 B.n94 163.367
R568 B.n554 B.n552 163.367
R569 B.n550 B.n96 163.367
R570 B.n546 B.n544 163.367
R571 B.n542 B.n98 163.367
R572 B.n538 B.n536 163.367
R573 B.n534 B.n100 163.367
R574 B.n530 B.n528 163.367
R575 B.n526 B.n102 163.367
R576 B.n522 B.n520 163.367
R577 B.n420 B.n140 163.367
R578 B.n424 B.n140 163.367
R579 B.n424 B.n134 163.367
R580 B.n432 B.n134 163.367
R581 B.n432 B.n132 163.367
R582 B.n436 B.n132 163.367
R583 B.n436 B.n126 163.367
R584 B.n444 B.n126 163.367
R585 B.n444 B.n124 163.367
R586 B.n448 B.n124 163.367
R587 B.n448 B.n119 163.367
R588 B.n457 B.n119 163.367
R589 B.n457 B.n117 163.367
R590 B.n461 B.n117 163.367
R591 B.n461 B.n112 163.367
R592 B.n470 B.n112 163.367
R593 B.n470 B.n110 163.367
R594 B.n475 B.n110 163.367
R595 B.n475 B.n105 163.367
R596 B.n484 B.n105 163.367
R597 B.n485 B.n484 163.367
R598 B.n485 B.n5 163.367
R599 B.n6 B.n5 163.367
R600 B.n7 B.n6 163.367
R601 B.n491 B.n7 163.367
R602 B.n492 B.n491 163.367
R603 B.n492 B.n13 163.367
R604 B.n14 B.n13 163.367
R605 B.n15 B.n14 163.367
R606 B.n497 B.n15 163.367
R607 B.n497 B.n20 163.367
R608 B.n21 B.n20 163.367
R609 B.n22 B.n21 163.367
R610 B.n502 B.n22 163.367
R611 B.n502 B.n27 163.367
R612 B.n28 B.n27 163.367
R613 B.n29 B.n28 163.367
R614 B.n507 B.n29 163.367
R615 B.n507 B.n34 163.367
R616 B.n35 B.n34 163.367
R617 B.n36 B.n35 163.367
R618 B.n512 B.n36 163.367
R619 B.n512 B.n41 163.367
R620 B.n42 B.n41 163.367
R621 B.n43 B.n42 163.367
R622 B.n414 B.n412 163.367
R623 B.n412 B.n411 163.367
R624 B.n408 B.n407 163.367
R625 B.n405 B.n148 163.367
R626 B.n401 B.n399 163.367
R627 B.n397 B.n150 163.367
R628 B.n393 B.n391 163.367
R629 B.n389 B.n152 163.367
R630 B.n385 B.n383 163.367
R631 B.n381 B.n154 163.367
R632 B.n377 B.n375 163.367
R633 B.n373 B.n156 163.367
R634 B.n369 B.n367 163.367
R635 B.n365 B.n158 163.367
R636 B.n361 B.n359 163.367
R637 B.n357 B.n160 163.367
R638 B.n353 B.n351 163.367
R639 B.n349 B.n162 163.367
R640 B.n345 B.n343 163.367
R641 B.n341 B.n164 163.367
R642 B.n337 B.n335 163.367
R643 B.n333 B.n166 163.367
R644 B.n329 B.n327 163.367
R645 B.n325 B.n168 163.367
R646 B.n321 B.n319 163.367
R647 B.n316 B.n315 163.367
R648 B.n313 B.n174 163.367
R649 B.n309 B.n307 163.367
R650 B.n305 B.n176 163.367
R651 B.n301 B.n299 163.367
R652 B.n296 B.n295 163.367
R653 B.n293 B.n182 163.367
R654 B.n289 B.n287 163.367
R655 B.n285 B.n184 163.367
R656 B.n281 B.n279 163.367
R657 B.n277 B.n186 163.367
R658 B.n273 B.n271 163.367
R659 B.n269 B.n188 163.367
R660 B.n265 B.n263 163.367
R661 B.n261 B.n190 163.367
R662 B.n257 B.n255 163.367
R663 B.n253 B.n192 163.367
R664 B.n249 B.n247 163.367
R665 B.n245 B.n194 163.367
R666 B.n241 B.n239 163.367
R667 B.n237 B.n196 163.367
R668 B.n233 B.n231 163.367
R669 B.n229 B.n198 163.367
R670 B.n225 B.n223 163.367
R671 B.n221 B.n200 163.367
R672 B.n217 B.n215 163.367
R673 B.n213 B.n202 163.367
R674 B.n209 B.n207 163.367
R675 B.n205 B.n142 163.367
R676 B.n418 B.n138 163.367
R677 B.n426 B.n138 163.367
R678 B.n426 B.n136 163.367
R679 B.n430 B.n136 163.367
R680 B.n430 B.n130 163.367
R681 B.n438 B.n130 163.367
R682 B.n438 B.n128 163.367
R683 B.n442 B.n128 163.367
R684 B.n442 B.n122 163.367
R685 B.n451 B.n122 163.367
R686 B.n451 B.n120 163.367
R687 B.n455 B.n120 163.367
R688 B.n455 B.n115 163.367
R689 B.n464 B.n115 163.367
R690 B.n464 B.n113 163.367
R691 B.n468 B.n113 163.367
R692 B.n468 B.n108 163.367
R693 B.n478 B.n108 163.367
R694 B.n478 B.n106 163.367
R695 B.n482 B.n106 163.367
R696 B.n482 B.n3 163.367
R697 B.n780 B.n3 163.367
R698 B.n776 B.n2 163.367
R699 B.n776 B.n775 163.367
R700 B.n775 B.n9 163.367
R701 B.n771 B.n9 163.367
R702 B.n771 B.n11 163.367
R703 B.n767 B.n11 163.367
R704 B.n767 B.n16 163.367
R705 B.n763 B.n16 163.367
R706 B.n763 B.n18 163.367
R707 B.n759 B.n18 163.367
R708 B.n759 B.n23 163.367
R709 B.n755 B.n23 163.367
R710 B.n755 B.n25 163.367
R711 B.n751 B.n25 163.367
R712 B.n751 B.n31 163.367
R713 B.n747 B.n31 163.367
R714 B.n747 B.n33 163.367
R715 B.n743 B.n33 163.367
R716 B.n743 B.n38 163.367
R717 B.n739 B.n38 163.367
R718 B.n739 B.n40 163.367
R719 B.n735 B.n40 163.367
R720 B.n419 B.n143 75.6341
R721 B.n736 B.n44 75.6341
R722 B.n730 B.n45 71.676
R723 B.n729 B.n728 71.676
R724 B.n722 B.n47 71.676
R725 B.n721 B.n720 71.676
R726 B.n714 B.n49 71.676
R727 B.n713 B.n712 71.676
R728 B.n706 B.n51 71.676
R729 B.n705 B.n704 71.676
R730 B.n698 B.n53 71.676
R731 B.n697 B.n696 71.676
R732 B.n690 B.n55 71.676
R733 B.n689 B.n688 71.676
R734 B.n682 B.n57 71.676
R735 B.n681 B.n680 71.676
R736 B.n674 B.n59 71.676
R737 B.n673 B.n672 71.676
R738 B.n666 B.n61 71.676
R739 B.n665 B.n664 71.676
R740 B.n658 B.n63 71.676
R741 B.n657 B.n656 71.676
R742 B.n650 B.n65 71.676
R743 B.n649 B.n648 71.676
R744 B.n642 B.n67 71.676
R745 B.n641 B.n640 71.676
R746 B.n633 B.n69 71.676
R747 B.n632 B.n631 71.676
R748 B.n625 B.n73 71.676
R749 B.n624 B.n623 71.676
R750 B.n617 B.n75 71.676
R751 B.n616 B.n615 71.676
R752 B.n609 B.n77 71.676
R753 B.n608 B.n607 71.676
R754 B.n601 B.n82 71.676
R755 B.n600 B.n599 71.676
R756 B.n593 B.n84 71.676
R757 B.n592 B.n591 71.676
R758 B.n585 B.n86 71.676
R759 B.n584 B.n583 71.676
R760 B.n577 B.n88 71.676
R761 B.n576 B.n575 71.676
R762 B.n569 B.n90 71.676
R763 B.n568 B.n567 71.676
R764 B.n561 B.n92 71.676
R765 B.n560 B.n559 71.676
R766 B.n553 B.n94 71.676
R767 B.n552 B.n551 71.676
R768 B.n545 B.n96 71.676
R769 B.n544 B.n543 71.676
R770 B.n537 B.n98 71.676
R771 B.n536 B.n535 71.676
R772 B.n529 B.n100 71.676
R773 B.n528 B.n527 71.676
R774 B.n521 B.n102 71.676
R775 B.n520 B.n519 71.676
R776 B.n519 B.n518 71.676
R777 B.n522 B.n521 71.676
R778 B.n527 B.n526 71.676
R779 B.n530 B.n529 71.676
R780 B.n535 B.n534 71.676
R781 B.n538 B.n537 71.676
R782 B.n543 B.n542 71.676
R783 B.n546 B.n545 71.676
R784 B.n551 B.n550 71.676
R785 B.n554 B.n553 71.676
R786 B.n559 B.n558 71.676
R787 B.n562 B.n561 71.676
R788 B.n567 B.n566 71.676
R789 B.n570 B.n569 71.676
R790 B.n575 B.n574 71.676
R791 B.n578 B.n577 71.676
R792 B.n583 B.n582 71.676
R793 B.n586 B.n585 71.676
R794 B.n591 B.n590 71.676
R795 B.n594 B.n593 71.676
R796 B.n599 B.n598 71.676
R797 B.n602 B.n601 71.676
R798 B.n607 B.n606 71.676
R799 B.n610 B.n609 71.676
R800 B.n615 B.n614 71.676
R801 B.n618 B.n617 71.676
R802 B.n623 B.n622 71.676
R803 B.n626 B.n625 71.676
R804 B.n631 B.n630 71.676
R805 B.n634 B.n633 71.676
R806 B.n640 B.n639 71.676
R807 B.n643 B.n642 71.676
R808 B.n648 B.n647 71.676
R809 B.n651 B.n650 71.676
R810 B.n656 B.n655 71.676
R811 B.n659 B.n658 71.676
R812 B.n664 B.n663 71.676
R813 B.n667 B.n666 71.676
R814 B.n672 B.n671 71.676
R815 B.n675 B.n674 71.676
R816 B.n680 B.n679 71.676
R817 B.n683 B.n682 71.676
R818 B.n688 B.n687 71.676
R819 B.n691 B.n690 71.676
R820 B.n696 B.n695 71.676
R821 B.n699 B.n698 71.676
R822 B.n704 B.n703 71.676
R823 B.n707 B.n706 71.676
R824 B.n712 B.n711 71.676
R825 B.n715 B.n714 71.676
R826 B.n720 B.n719 71.676
R827 B.n723 B.n722 71.676
R828 B.n728 B.n727 71.676
R829 B.n731 B.n730 71.676
R830 B.n413 B.n144 71.676
R831 B.n411 B.n146 71.676
R832 B.n407 B.n406 71.676
R833 B.n400 B.n148 71.676
R834 B.n399 B.n398 71.676
R835 B.n392 B.n150 71.676
R836 B.n391 B.n390 71.676
R837 B.n384 B.n152 71.676
R838 B.n383 B.n382 71.676
R839 B.n376 B.n154 71.676
R840 B.n375 B.n374 71.676
R841 B.n368 B.n156 71.676
R842 B.n367 B.n366 71.676
R843 B.n360 B.n158 71.676
R844 B.n359 B.n358 71.676
R845 B.n352 B.n160 71.676
R846 B.n351 B.n350 71.676
R847 B.n344 B.n162 71.676
R848 B.n343 B.n342 71.676
R849 B.n336 B.n164 71.676
R850 B.n335 B.n334 71.676
R851 B.n328 B.n166 71.676
R852 B.n327 B.n326 71.676
R853 B.n320 B.n168 71.676
R854 B.n319 B.n172 71.676
R855 B.n315 B.n314 71.676
R856 B.n308 B.n174 71.676
R857 B.n307 B.n306 71.676
R858 B.n300 B.n176 71.676
R859 B.n299 B.n180 71.676
R860 B.n295 B.n294 71.676
R861 B.n288 B.n182 71.676
R862 B.n287 B.n286 71.676
R863 B.n280 B.n184 71.676
R864 B.n279 B.n278 71.676
R865 B.n272 B.n186 71.676
R866 B.n271 B.n270 71.676
R867 B.n264 B.n188 71.676
R868 B.n263 B.n262 71.676
R869 B.n256 B.n190 71.676
R870 B.n255 B.n254 71.676
R871 B.n248 B.n192 71.676
R872 B.n247 B.n246 71.676
R873 B.n240 B.n194 71.676
R874 B.n239 B.n238 71.676
R875 B.n232 B.n196 71.676
R876 B.n231 B.n230 71.676
R877 B.n224 B.n198 71.676
R878 B.n223 B.n222 71.676
R879 B.n216 B.n200 71.676
R880 B.n215 B.n214 71.676
R881 B.n208 B.n202 71.676
R882 B.n207 B.n206 71.676
R883 B.n414 B.n413 71.676
R884 B.n408 B.n146 71.676
R885 B.n406 B.n405 71.676
R886 B.n401 B.n400 71.676
R887 B.n398 B.n397 71.676
R888 B.n393 B.n392 71.676
R889 B.n390 B.n389 71.676
R890 B.n385 B.n384 71.676
R891 B.n382 B.n381 71.676
R892 B.n377 B.n376 71.676
R893 B.n374 B.n373 71.676
R894 B.n369 B.n368 71.676
R895 B.n366 B.n365 71.676
R896 B.n361 B.n360 71.676
R897 B.n358 B.n357 71.676
R898 B.n353 B.n352 71.676
R899 B.n350 B.n349 71.676
R900 B.n345 B.n344 71.676
R901 B.n342 B.n341 71.676
R902 B.n337 B.n336 71.676
R903 B.n334 B.n333 71.676
R904 B.n329 B.n328 71.676
R905 B.n326 B.n325 71.676
R906 B.n321 B.n320 71.676
R907 B.n316 B.n172 71.676
R908 B.n314 B.n313 71.676
R909 B.n309 B.n308 71.676
R910 B.n306 B.n305 71.676
R911 B.n301 B.n300 71.676
R912 B.n296 B.n180 71.676
R913 B.n294 B.n293 71.676
R914 B.n289 B.n288 71.676
R915 B.n286 B.n285 71.676
R916 B.n281 B.n280 71.676
R917 B.n278 B.n277 71.676
R918 B.n273 B.n272 71.676
R919 B.n270 B.n269 71.676
R920 B.n265 B.n264 71.676
R921 B.n262 B.n261 71.676
R922 B.n257 B.n256 71.676
R923 B.n254 B.n253 71.676
R924 B.n249 B.n248 71.676
R925 B.n246 B.n245 71.676
R926 B.n241 B.n240 71.676
R927 B.n238 B.n237 71.676
R928 B.n233 B.n232 71.676
R929 B.n230 B.n229 71.676
R930 B.n225 B.n224 71.676
R931 B.n222 B.n221 71.676
R932 B.n217 B.n216 71.676
R933 B.n214 B.n213 71.676
R934 B.n209 B.n208 71.676
R935 B.n206 B.n205 71.676
R936 B.n781 B.n780 71.676
R937 B.n781 B.n2 71.676
R938 B.n636 B.n71 59.5399
R939 B.n80 B.n79 59.5399
R940 B.n179 B.n178 59.5399
R941 B.n171 B.n170 59.5399
R942 B.n419 B.n139 37.5413
R943 B.n425 B.n139 37.5413
R944 B.n425 B.n135 37.5413
R945 B.n431 B.n135 37.5413
R946 B.n437 B.n131 37.5413
R947 B.n437 B.n127 37.5413
R948 B.n443 B.n127 37.5413
R949 B.n443 B.n123 37.5413
R950 B.n450 B.n123 37.5413
R951 B.n450 B.n449 37.5413
R952 B.n456 B.n116 37.5413
R953 B.n463 B.n116 37.5413
R954 B.n463 B.n462 37.5413
R955 B.n469 B.n109 37.5413
R956 B.n477 B.n109 37.5413
R957 B.n477 B.n476 37.5413
R958 B.n483 B.n4 37.5413
R959 B.n779 B.n4 37.5413
R960 B.n779 B.n778 37.5413
R961 B.n778 B.n777 37.5413
R962 B.n777 B.n8 37.5413
R963 B.n770 B.n12 37.5413
R964 B.n770 B.n769 37.5413
R965 B.n769 B.n768 37.5413
R966 B.n762 B.n19 37.5413
R967 B.n762 B.n761 37.5413
R968 B.n761 B.n760 37.5413
R969 B.n754 B.n26 37.5413
R970 B.n754 B.n753 37.5413
R971 B.n753 B.n752 37.5413
R972 B.n752 B.n30 37.5413
R973 B.n746 B.n30 37.5413
R974 B.n746 B.n745 37.5413
R975 B.n744 B.n37 37.5413
R976 B.n738 B.n37 37.5413
R977 B.n738 B.n737 37.5413
R978 B.n737 B.n736 37.5413
R979 B.n417 B.n416 36.6834
R980 B.n421 B.n141 36.6834
R981 B.n517 B.n516 36.6834
R982 B.n734 B.n733 36.6834
R983 B.n431 B.t11 34.7809
R984 B.n483 B.t5 34.7809
R985 B.t4 B.n8 34.7809
R986 B.t7 B.n744 34.7809
R987 B.n449 B.t1 29.2602
R988 B.n26 B.t0 29.2602
R989 B.n71 B.n70 24.049
R990 B.n79 B.n78 24.049
R991 B.n178 B.n177 24.049
R992 B.n170 B.n169 24.049
R993 B.n469 B.t2 21.5312
R994 B.n768 B.t3 21.5312
R995 B B.n782 18.0485
R996 B.n462 B.t2 16.0105
R997 B.n19 B.t3 16.0105
R998 B.n417 B.n137 10.6151
R999 B.n427 B.n137 10.6151
R1000 B.n428 B.n427 10.6151
R1001 B.n429 B.n428 10.6151
R1002 B.n429 B.n129 10.6151
R1003 B.n439 B.n129 10.6151
R1004 B.n440 B.n439 10.6151
R1005 B.n441 B.n440 10.6151
R1006 B.n441 B.n121 10.6151
R1007 B.n452 B.n121 10.6151
R1008 B.n453 B.n452 10.6151
R1009 B.n454 B.n453 10.6151
R1010 B.n454 B.n114 10.6151
R1011 B.n465 B.n114 10.6151
R1012 B.n466 B.n465 10.6151
R1013 B.n467 B.n466 10.6151
R1014 B.n467 B.n107 10.6151
R1015 B.n479 B.n107 10.6151
R1016 B.n480 B.n479 10.6151
R1017 B.n481 B.n480 10.6151
R1018 B.n481 B.n0 10.6151
R1019 B.n416 B.n415 10.6151
R1020 B.n415 B.n145 10.6151
R1021 B.n410 B.n145 10.6151
R1022 B.n410 B.n409 10.6151
R1023 B.n409 B.n147 10.6151
R1024 B.n404 B.n147 10.6151
R1025 B.n404 B.n403 10.6151
R1026 B.n403 B.n402 10.6151
R1027 B.n402 B.n149 10.6151
R1028 B.n396 B.n149 10.6151
R1029 B.n396 B.n395 10.6151
R1030 B.n395 B.n394 10.6151
R1031 B.n394 B.n151 10.6151
R1032 B.n388 B.n151 10.6151
R1033 B.n388 B.n387 10.6151
R1034 B.n387 B.n386 10.6151
R1035 B.n386 B.n153 10.6151
R1036 B.n380 B.n153 10.6151
R1037 B.n380 B.n379 10.6151
R1038 B.n379 B.n378 10.6151
R1039 B.n378 B.n155 10.6151
R1040 B.n372 B.n155 10.6151
R1041 B.n372 B.n371 10.6151
R1042 B.n371 B.n370 10.6151
R1043 B.n370 B.n157 10.6151
R1044 B.n364 B.n157 10.6151
R1045 B.n364 B.n363 10.6151
R1046 B.n363 B.n362 10.6151
R1047 B.n362 B.n159 10.6151
R1048 B.n356 B.n159 10.6151
R1049 B.n356 B.n355 10.6151
R1050 B.n355 B.n354 10.6151
R1051 B.n354 B.n161 10.6151
R1052 B.n348 B.n161 10.6151
R1053 B.n348 B.n347 10.6151
R1054 B.n347 B.n346 10.6151
R1055 B.n346 B.n163 10.6151
R1056 B.n340 B.n163 10.6151
R1057 B.n340 B.n339 10.6151
R1058 B.n339 B.n338 10.6151
R1059 B.n338 B.n165 10.6151
R1060 B.n332 B.n165 10.6151
R1061 B.n332 B.n331 10.6151
R1062 B.n331 B.n330 10.6151
R1063 B.n330 B.n167 10.6151
R1064 B.n324 B.n167 10.6151
R1065 B.n324 B.n323 10.6151
R1066 B.n323 B.n322 10.6151
R1067 B.n318 B.n317 10.6151
R1068 B.n317 B.n173 10.6151
R1069 B.n312 B.n173 10.6151
R1070 B.n312 B.n311 10.6151
R1071 B.n311 B.n310 10.6151
R1072 B.n310 B.n175 10.6151
R1073 B.n304 B.n175 10.6151
R1074 B.n304 B.n303 10.6151
R1075 B.n303 B.n302 10.6151
R1076 B.n298 B.n297 10.6151
R1077 B.n297 B.n181 10.6151
R1078 B.n292 B.n181 10.6151
R1079 B.n292 B.n291 10.6151
R1080 B.n291 B.n290 10.6151
R1081 B.n290 B.n183 10.6151
R1082 B.n284 B.n183 10.6151
R1083 B.n284 B.n283 10.6151
R1084 B.n283 B.n282 10.6151
R1085 B.n282 B.n185 10.6151
R1086 B.n276 B.n185 10.6151
R1087 B.n276 B.n275 10.6151
R1088 B.n275 B.n274 10.6151
R1089 B.n274 B.n187 10.6151
R1090 B.n268 B.n187 10.6151
R1091 B.n268 B.n267 10.6151
R1092 B.n267 B.n266 10.6151
R1093 B.n266 B.n189 10.6151
R1094 B.n260 B.n189 10.6151
R1095 B.n260 B.n259 10.6151
R1096 B.n259 B.n258 10.6151
R1097 B.n258 B.n191 10.6151
R1098 B.n252 B.n191 10.6151
R1099 B.n252 B.n251 10.6151
R1100 B.n251 B.n250 10.6151
R1101 B.n250 B.n193 10.6151
R1102 B.n244 B.n193 10.6151
R1103 B.n244 B.n243 10.6151
R1104 B.n243 B.n242 10.6151
R1105 B.n242 B.n195 10.6151
R1106 B.n236 B.n195 10.6151
R1107 B.n236 B.n235 10.6151
R1108 B.n235 B.n234 10.6151
R1109 B.n234 B.n197 10.6151
R1110 B.n228 B.n197 10.6151
R1111 B.n228 B.n227 10.6151
R1112 B.n227 B.n226 10.6151
R1113 B.n226 B.n199 10.6151
R1114 B.n220 B.n199 10.6151
R1115 B.n220 B.n219 10.6151
R1116 B.n219 B.n218 10.6151
R1117 B.n218 B.n201 10.6151
R1118 B.n212 B.n201 10.6151
R1119 B.n212 B.n211 10.6151
R1120 B.n211 B.n210 10.6151
R1121 B.n210 B.n203 10.6151
R1122 B.n204 B.n203 10.6151
R1123 B.n204 B.n141 10.6151
R1124 B.n422 B.n421 10.6151
R1125 B.n423 B.n422 10.6151
R1126 B.n423 B.n133 10.6151
R1127 B.n433 B.n133 10.6151
R1128 B.n434 B.n433 10.6151
R1129 B.n435 B.n434 10.6151
R1130 B.n435 B.n125 10.6151
R1131 B.n445 B.n125 10.6151
R1132 B.n446 B.n445 10.6151
R1133 B.n447 B.n446 10.6151
R1134 B.n447 B.n118 10.6151
R1135 B.n458 B.n118 10.6151
R1136 B.n459 B.n458 10.6151
R1137 B.n460 B.n459 10.6151
R1138 B.n460 B.n111 10.6151
R1139 B.n471 B.n111 10.6151
R1140 B.n472 B.n471 10.6151
R1141 B.n474 B.n472 10.6151
R1142 B.n474 B.n473 10.6151
R1143 B.n473 B.n104 10.6151
R1144 B.n486 B.n104 10.6151
R1145 B.n487 B.n486 10.6151
R1146 B.n488 B.n487 10.6151
R1147 B.n489 B.n488 10.6151
R1148 B.n490 B.n489 10.6151
R1149 B.n493 B.n490 10.6151
R1150 B.n494 B.n493 10.6151
R1151 B.n495 B.n494 10.6151
R1152 B.n496 B.n495 10.6151
R1153 B.n498 B.n496 10.6151
R1154 B.n499 B.n498 10.6151
R1155 B.n500 B.n499 10.6151
R1156 B.n501 B.n500 10.6151
R1157 B.n503 B.n501 10.6151
R1158 B.n504 B.n503 10.6151
R1159 B.n505 B.n504 10.6151
R1160 B.n506 B.n505 10.6151
R1161 B.n508 B.n506 10.6151
R1162 B.n509 B.n508 10.6151
R1163 B.n510 B.n509 10.6151
R1164 B.n511 B.n510 10.6151
R1165 B.n513 B.n511 10.6151
R1166 B.n514 B.n513 10.6151
R1167 B.n515 B.n514 10.6151
R1168 B.n516 B.n515 10.6151
R1169 B.n774 B.n1 10.6151
R1170 B.n774 B.n773 10.6151
R1171 B.n773 B.n772 10.6151
R1172 B.n772 B.n10 10.6151
R1173 B.n766 B.n10 10.6151
R1174 B.n766 B.n765 10.6151
R1175 B.n765 B.n764 10.6151
R1176 B.n764 B.n17 10.6151
R1177 B.n758 B.n17 10.6151
R1178 B.n758 B.n757 10.6151
R1179 B.n757 B.n756 10.6151
R1180 B.n756 B.n24 10.6151
R1181 B.n750 B.n24 10.6151
R1182 B.n750 B.n749 10.6151
R1183 B.n749 B.n748 10.6151
R1184 B.n748 B.n32 10.6151
R1185 B.n742 B.n32 10.6151
R1186 B.n742 B.n741 10.6151
R1187 B.n741 B.n740 10.6151
R1188 B.n740 B.n39 10.6151
R1189 B.n734 B.n39 10.6151
R1190 B.n733 B.n732 10.6151
R1191 B.n732 B.n46 10.6151
R1192 B.n726 B.n46 10.6151
R1193 B.n726 B.n725 10.6151
R1194 B.n725 B.n724 10.6151
R1195 B.n724 B.n48 10.6151
R1196 B.n718 B.n48 10.6151
R1197 B.n718 B.n717 10.6151
R1198 B.n717 B.n716 10.6151
R1199 B.n716 B.n50 10.6151
R1200 B.n710 B.n50 10.6151
R1201 B.n710 B.n709 10.6151
R1202 B.n709 B.n708 10.6151
R1203 B.n708 B.n52 10.6151
R1204 B.n702 B.n52 10.6151
R1205 B.n702 B.n701 10.6151
R1206 B.n701 B.n700 10.6151
R1207 B.n700 B.n54 10.6151
R1208 B.n694 B.n54 10.6151
R1209 B.n694 B.n693 10.6151
R1210 B.n693 B.n692 10.6151
R1211 B.n692 B.n56 10.6151
R1212 B.n686 B.n56 10.6151
R1213 B.n686 B.n685 10.6151
R1214 B.n685 B.n684 10.6151
R1215 B.n684 B.n58 10.6151
R1216 B.n678 B.n58 10.6151
R1217 B.n678 B.n677 10.6151
R1218 B.n677 B.n676 10.6151
R1219 B.n676 B.n60 10.6151
R1220 B.n670 B.n60 10.6151
R1221 B.n670 B.n669 10.6151
R1222 B.n669 B.n668 10.6151
R1223 B.n668 B.n62 10.6151
R1224 B.n662 B.n62 10.6151
R1225 B.n662 B.n661 10.6151
R1226 B.n661 B.n660 10.6151
R1227 B.n660 B.n64 10.6151
R1228 B.n654 B.n64 10.6151
R1229 B.n654 B.n653 10.6151
R1230 B.n653 B.n652 10.6151
R1231 B.n652 B.n66 10.6151
R1232 B.n646 B.n66 10.6151
R1233 B.n646 B.n645 10.6151
R1234 B.n645 B.n644 10.6151
R1235 B.n644 B.n68 10.6151
R1236 B.n638 B.n68 10.6151
R1237 B.n638 B.n637 10.6151
R1238 B.n635 B.n72 10.6151
R1239 B.n629 B.n72 10.6151
R1240 B.n629 B.n628 10.6151
R1241 B.n628 B.n627 10.6151
R1242 B.n627 B.n74 10.6151
R1243 B.n621 B.n74 10.6151
R1244 B.n621 B.n620 10.6151
R1245 B.n620 B.n619 10.6151
R1246 B.n619 B.n76 10.6151
R1247 B.n613 B.n612 10.6151
R1248 B.n612 B.n611 10.6151
R1249 B.n611 B.n81 10.6151
R1250 B.n605 B.n81 10.6151
R1251 B.n605 B.n604 10.6151
R1252 B.n604 B.n603 10.6151
R1253 B.n603 B.n83 10.6151
R1254 B.n597 B.n83 10.6151
R1255 B.n597 B.n596 10.6151
R1256 B.n596 B.n595 10.6151
R1257 B.n595 B.n85 10.6151
R1258 B.n589 B.n85 10.6151
R1259 B.n589 B.n588 10.6151
R1260 B.n588 B.n587 10.6151
R1261 B.n587 B.n87 10.6151
R1262 B.n581 B.n87 10.6151
R1263 B.n581 B.n580 10.6151
R1264 B.n580 B.n579 10.6151
R1265 B.n579 B.n89 10.6151
R1266 B.n573 B.n89 10.6151
R1267 B.n573 B.n572 10.6151
R1268 B.n572 B.n571 10.6151
R1269 B.n571 B.n91 10.6151
R1270 B.n565 B.n91 10.6151
R1271 B.n565 B.n564 10.6151
R1272 B.n564 B.n563 10.6151
R1273 B.n563 B.n93 10.6151
R1274 B.n557 B.n93 10.6151
R1275 B.n557 B.n556 10.6151
R1276 B.n556 B.n555 10.6151
R1277 B.n555 B.n95 10.6151
R1278 B.n549 B.n95 10.6151
R1279 B.n549 B.n548 10.6151
R1280 B.n548 B.n547 10.6151
R1281 B.n547 B.n97 10.6151
R1282 B.n541 B.n97 10.6151
R1283 B.n541 B.n540 10.6151
R1284 B.n540 B.n539 10.6151
R1285 B.n539 B.n99 10.6151
R1286 B.n533 B.n99 10.6151
R1287 B.n533 B.n532 10.6151
R1288 B.n532 B.n531 10.6151
R1289 B.n531 B.n101 10.6151
R1290 B.n525 B.n101 10.6151
R1291 B.n525 B.n524 10.6151
R1292 B.n524 B.n523 10.6151
R1293 B.n523 B.n103 10.6151
R1294 B.n517 B.n103 10.6151
R1295 B.n322 B.n171 9.36635
R1296 B.n298 B.n179 9.36635
R1297 B.n637 B.n636 9.36635
R1298 B.n613 B.n80 9.36635
R1299 B.n456 B.t1 8.28155
R1300 B.n760 B.t0 8.28155
R1301 B.n782 B.n0 8.11757
R1302 B.n782 B.n1 8.11757
R1303 B.t11 B.n131 2.76085
R1304 B.n476 B.t5 2.76085
R1305 B.n12 B.t4 2.76085
R1306 B.n745 B.t7 2.76085
R1307 B.n318 B.n171 1.24928
R1308 B.n302 B.n179 1.24928
R1309 B.n636 B.n635 1.24928
R1310 B.n80 B.n76 1.24928
R1311 VN.n2 VN.t1 448.873
R1312 VN.n10 VN.t5 448.873
R1313 VN.n6 VN.t0 431.418
R1314 VN.n14 VN.t4 431.418
R1315 VN.n1 VN.t3 387.985
R1316 VN.n9 VN.t2 387.985
R1317 VN.n7 VN.n6 161.3
R1318 VN.n15 VN.n14 161.3
R1319 VN.n13 VN.n8 161.3
R1320 VN.n12 VN.n11 161.3
R1321 VN.n5 VN.n0 161.3
R1322 VN.n4 VN.n3 161.3
R1323 VN.n5 VN.n4 53.1199
R1324 VN.n13 VN.n12 53.1199
R1325 VN VN.n15 44.4342
R1326 VN.n11 VN.n10 43.5004
R1327 VN.n3 VN.n2 43.5004
R1328 VN.n2 VN.n1 42.494
R1329 VN.n10 VN.n9 42.494
R1330 VN.n4 VN.n1 12.234
R1331 VN.n12 VN.n9 12.234
R1332 VN.n6 VN.n5 5.11262
R1333 VN.n14 VN.n13 5.11262
R1334 VN.n15 VN.n8 0.189894
R1335 VN.n11 VN.n8 0.189894
R1336 VN.n3 VN.n0 0.189894
R1337 VN.n7 VN.n0 0.189894
R1338 VN VN.n7 0.0516364
R1339 VTAIL.n330 VTAIL.n254 289.615
R1340 VTAIL.n78 VTAIL.n2 289.615
R1341 VTAIL.n248 VTAIL.n172 289.615
R1342 VTAIL.n164 VTAIL.n88 289.615
R1343 VTAIL.n281 VTAIL.n280 185
R1344 VTAIL.n278 VTAIL.n277 185
R1345 VTAIL.n287 VTAIL.n286 185
R1346 VTAIL.n289 VTAIL.n288 185
R1347 VTAIL.n274 VTAIL.n273 185
R1348 VTAIL.n295 VTAIL.n294 185
R1349 VTAIL.n297 VTAIL.n296 185
R1350 VTAIL.n270 VTAIL.n269 185
R1351 VTAIL.n303 VTAIL.n302 185
R1352 VTAIL.n305 VTAIL.n304 185
R1353 VTAIL.n266 VTAIL.n265 185
R1354 VTAIL.n311 VTAIL.n310 185
R1355 VTAIL.n313 VTAIL.n312 185
R1356 VTAIL.n262 VTAIL.n261 185
R1357 VTAIL.n319 VTAIL.n318 185
R1358 VTAIL.n322 VTAIL.n321 185
R1359 VTAIL.n320 VTAIL.n258 185
R1360 VTAIL.n327 VTAIL.n257 185
R1361 VTAIL.n329 VTAIL.n328 185
R1362 VTAIL.n331 VTAIL.n330 185
R1363 VTAIL.n29 VTAIL.n28 185
R1364 VTAIL.n26 VTAIL.n25 185
R1365 VTAIL.n35 VTAIL.n34 185
R1366 VTAIL.n37 VTAIL.n36 185
R1367 VTAIL.n22 VTAIL.n21 185
R1368 VTAIL.n43 VTAIL.n42 185
R1369 VTAIL.n45 VTAIL.n44 185
R1370 VTAIL.n18 VTAIL.n17 185
R1371 VTAIL.n51 VTAIL.n50 185
R1372 VTAIL.n53 VTAIL.n52 185
R1373 VTAIL.n14 VTAIL.n13 185
R1374 VTAIL.n59 VTAIL.n58 185
R1375 VTAIL.n61 VTAIL.n60 185
R1376 VTAIL.n10 VTAIL.n9 185
R1377 VTAIL.n67 VTAIL.n66 185
R1378 VTAIL.n70 VTAIL.n69 185
R1379 VTAIL.n68 VTAIL.n6 185
R1380 VTAIL.n75 VTAIL.n5 185
R1381 VTAIL.n77 VTAIL.n76 185
R1382 VTAIL.n79 VTAIL.n78 185
R1383 VTAIL.n249 VTAIL.n248 185
R1384 VTAIL.n247 VTAIL.n246 185
R1385 VTAIL.n245 VTAIL.n175 185
R1386 VTAIL.n179 VTAIL.n176 185
R1387 VTAIL.n240 VTAIL.n239 185
R1388 VTAIL.n238 VTAIL.n237 185
R1389 VTAIL.n181 VTAIL.n180 185
R1390 VTAIL.n232 VTAIL.n231 185
R1391 VTAIL.n230 VTAIL.n229 185
R1392 VTAIL.n185 VTAIL.n184 185
R1393 VTAIL.n224 VTAIL.n223 185
R1394 VTAIL.n222 VTAIL.n221 185
R1395 VTAIL.n189 VTAIL.n188 185
R1396 VTAIL.n216 VTAIL.n215 185
R1397 VTAIL.n214 VTAIL.n213 185
R1398 VTAIL.n193 VTAIL.n192 185
R1399 VTAIL.n208 VTAIL.n207 185
R1400 VTAIL.n206 VTAIL.n205 185
R1401 VTAIL.n197 VTAIL.n196 185
R1402 VTAIL.n200 VTAIL.n199 185
R1403 VTAIL.n165 VTAIL.n164 185
R1404 VTAIL.n163 VTAIL.n162 185
R1405 VTAIL.n161 VTAIL.n91 185
R1406 VTAIL.n95 VTAIL.n92 185
R1407 VTAIL.n156 VTAIL.n155 185
R1408 VTAIL.n154 VTAIL.n153 185
R1409 VTAIL.n97 VTAIL.n96 185
R1410 VTAIL.n148 VTAIL.n147 185
R1411 VTAIL.n146 VTAIL.n145 185
R1412 VTAIL.n101 VTAIL.n100 185
R1413 VTAIL.n140 VTAIL.n139 185
R1414 VTAIL.n138 VTAIL.n137 185
R1415 VTAIL.n105 VTAIL.n104 185
R1416 VTAIL.n132 VTAIL.n131 185
R1417 VTAIL.n130 VTAIL.n129 185
R1418 VTAIL.n109 VTAIL.n108 185
R1419 VTAIL.n124 VTAIL.n123 185
R1420 VTAIL.n122 VTAIL.n121 185
R1421 VTAIL.n113 VTAIL.n112 185
R1422 VTAIL.n116 VTAIL.n115 185
R1423 VTAIL.t2 VTAIL.n198 147.659
R1424 VTAIL.t10 VTAIL.n114 147.659
R1425 VTAIL.t5 VTAIL.n279 147.659
R1426 VTAIL.t4 VTAIL.n27 147.659
R1427 VTAIL.n280 VTAIL.n277 104.615
R1428 VTAIL.n287 VTAIL.n277 104.615
R1429 VTAIL.n288 VTAIL.n287 104.615
R1430 VTAIL.n288 VTAIL.n273 104.615
R1431 VTAIL.n295 VTAIL.n273 104.615
R1432 VTAIL.n296 VTAIL.n295 104.615
R1433 VTAIL.n296 VTAIL.n269 104.615
R1434 VTAIL.n303 VTAIL.n269 104.615
R1435 VTAIL.n304 VTAIL.n303 104.615
R1436 VTAIL.n304 VTAIL.n265 104.615
R1437 VTAIL.n311 VTAIL.n265 104.615
R1438 VTAIL.n312 VTAIL.n311 104.615
R1439 VTAIL.n312 VTAIL.n261 104.615
R1440 VTAIL.n319 VTAIL.n261 104.615
R1441 VTAIL.n321 VTAIL.n319 104.615
R1442 VTAIL.n321 VTAIL.n320 104.615
R1443 VTAIL.n320 VTAIL.n257 104.615
R1444 VTAIL.n329 VTAIL.n257 104.615
R1445 VTAIL.n330 VTAIL.n329 104.615
R1446 VTAIL.n28 VTAIL.n25 104.615
R1447 VTAIL.n35 VTAIL.n25 104.615
R1448 VTAIL.n36 VTAIL.n35 104.615
R1449 VTAIL.n36 VTAIL.n21 104.615
R1450 VTAIL.n43 VTAIL.n21 104.615
R1451 VTAIL.n44 VTAIL.n43 104.615
R1452 VTAIL.n44 VTAIL.n17 104.615
R1453 VTAIL.n51 VTAIL.n17 104.615
R1454 VTAIL.n52 VTAIL.n51 104.615
R1455 VTAIL.n52 VTAIL.n13 104.615
R1456 VTAIL.n59 VTAIL.n13 104.615
R1457 VTAIL.n60 VTAIL.n59 104.615
R1458 VTAIL.n60 VTAIL.n9 104.615
R1459 VTAIL.n67 VTAIL.n9 104.615
R1460 VTAIL.n69 VTAIL.n67 104.615
R1461 VTAIL.n69 VTAIL.n68 104.615
R1462 VTAIL.n68 VTAIL.n5 104.615
R1463 VTAIL.n77 VTAIL.n5 104.615
R1464 VTAIL.n78 VTAIL.n77 104.615
R1465 VTAIL.n248 VTAIL.n247 104.615
R1466 VTAIL.n247 VTAIL.n175 104.615
R1467 VTAIL.n179 VTAIL.n175 104.615
R1468 VTAIL.n239 VTAIL.n179 104.615
R1469 VTAIL.n239 VTAIL.n238 104.615
R1470 VTAIL.n238 VTAIL.n180 104.615
R1471 VTAIL.n231 VTAIL.n180 104.615
R1472 VTAIL.n231 VTAIL.n230 104.615
R1473 VTAIL.n230 VTAIL.n184 104.615
R1474 VTAIL.n223 VTAIL.n184 104.615
R1475 VTAIL.n223 VTAIL.n222 104.615
R1476 VTAIL.n222 VTAIL.n188 104.615
R1477 VTAIL.n215 VTAIL.n188 104.615
R1478 VTAIL.n215 VTAIL.n214 104.615
R1479 VTAIL.n214 VTAIL.n192 104.615
R1480 VTAIL.n207 VTAIL.n192 104.615
R1481 VTAIL.n207 VTAIL.n206 104.615
R1482 VTAIL.n206 VTAIL.n196 104.615
R1483 VTAIL.n199 VTAIL.n196 104.615
R1484 VTAIL.n164 VTAIL.n163 104.615
R1485 VTAIL.n163 VTAIL.n91 104.615
R1486 VTAIL.n95 VTAIL.n91 104.615
R1487 VTAIL.n155 VTAIL.n95 104.615
R1488 VTAIL.n155 VTAIL.n154 104.615
R1489 VTAIL.n154 VTAIL.n96 104.615
R1490 VTAIL.n147 VTAIL.n96 104.615
R1491 VTAIL.n147 VTAIL.n146 104.615
R1492 VTAIL.n146 VTAIL.n100 104.615
R1493 VTAIL.n139 VTAIL.n100 104.615
R1494 VTAIL.n139 VTAIL.n138 104.615
R1495 VTAIL.n138 VTAIL.n104 104.615
R1496 VTAIL.n131 VTAIL.n104 104.615
R1497 VTAIL.n131 VTAIL.n130 104.615
R1498 VTAIL.n130 VTAIL.n108 104.615
R1499 VTAIL.n123 VTAIL.n108 104.615
R1500 VTAIL.n123 VTAIL.n122 104.615
R1501 VTAIL.n122 VTAIL.n112 104.615
R1502 VTAIL.n115 VTAIL.n112 104.615
R1503 VTAIL.n280 VTAIL.t5 52.3082
R1504 VTAIL.n28 VTAIL.t4 52.3082
R1505 VTAIL.n199 VTAIL.t2 52.3082
R1506 VTAIL.n115 VTAIL.t10 52.3082
R1507 VTAIL.n171 VTAIL.n170 44.4362
R1508 VTAIL.n87 VTAIL.n86 44.4362
R1509 VTAIL.n1 VTAIL.n0 44.4361
R1510 VTAIL.n85 VTAIL.n84 44.4361
R1511 VTAIL.n335 VTAIL.n334 32.3793
R1512 VTAIL.n83 VTAIL.n82 32.3793
R1513 VTAIL.n253 VTAIL.n252 32.3793
R1514 VTAIL.n169 VTAIL.n168 32.3793
R1515 VTAIL.n87 VTAIL.n85 27.1341
R1516 VTAIL.n335 VTAIL.n253 26.0652
R1517 VTAIL.n281 VTAIL.n279 15.6677
R1518 VTAIL.n29 VTAIL.n27 15.6677
R1519 VTAIL.n200 VTAIL.n198 15.6677
R1520 VTAIL.n116 VTAIL.n114 15.6677
R1521 VTAIL.n328 VTAIL.n327 13.1884
R1522 VTAIL.n76 VTAIL.n75 13.1884
R1523 VTAIL.n246 VTAIL.n245 13.1884
R1524 VTAIL.n162 VTAIL.n161 13.1884
R1525 VTAIL.n282 VTAIL.n278 12.8005
R1526 VTAIL.n326 VTAIL.n258 12.8005
R1527 VTAIL.n331 VTAIL.n256 12.8005
R1528 VTAIL.n30 VTAIL.n26 12.8005
R1529 VTAIL.n74 VTAIL.n6 12.8005
R1530 VTAIL.n79 VTAIL.n4 12.8005
R1531 VTAIL.n249 VTAIL.n174 12.8005
R1532 VTAIL.n244 VTAIL.n176 12.8005
R1533 VTAIL.n201 VTAIL.n197 12.8005
R1534 VTAIL.n165 VTAIL.n90 12.8005
R1535 VTAIL.n160 VTAIL.n92 12.8005
R1536 VTAIL.n117 VTAIL.n113 12.8005
R1537 VTAIL.n286 VTAIL.n285 12.0247
R1538 VTAIL.n323 VTAIL.n322 12.0247
R1539 VTAIL.n332 VTAIL.n254 12.0247
R1540 VTAIL.n34 VTAIL.n33 12.0247
R1541 VTAIL.n71 VTAIL.n70 12.0247
R1542 VTAIL.n80 VTAIL.n2 12.0247
R1543 VTAIL.n250 VTAIL.n172 12.0247
R1544 VTAIL.n241 VTAIL.n240 12.0247
R1545 VTAIL.n205 VTAIL.n204 12.0247
R1546 VTAIL.n166 VTAIL.n88 12.0247
R1547 VTAIL.n157 VTAIL.n156 12.0247
R1548 VTAIL.n121 VTAIL.n120 12.0247
R1549 VTAIL.n289 VTAIL.n276 11.249
R1550 VTAIL.n318 VTAIL.n260 11.249
R1551 VTAIL.n37 VTAIL.n24 11.249
R1552 VTAIL.n66 VTAIL.n8 11.249
R1553 VTAIL.n237 VTAIL.n178 11.249
R1554 VTAIL.n208 VTAIL.n195 11.249
R1555 VTAIL.n153 VTAIL.n94 11.249
R1556 VTAIL.n124 VTAIL.n111 11.249
R1557 VTAIL.n290 VTAIL.n274 10.4732
R1558 VTAIL.n317 VTAIL.n262 10.4732
R1559 VTAIL.n38 VTAIL.n22 10.4732
R1560 VTAIL.n65 VTAIL.n10 10.4732
R1561 VTAIL.n236 VTAIL.n181 10.4732
R1562 VTAIL.n209 VTAIL.n193 10.4732
R1563 VTAIL.n152 VTAIL.n97 10.4732
R1564 VTAIL.n125 VTAIL.n109 10.4732
R1565 VTAIL.n294 VTAIL.n293 9.69747
R1566 VTAIL.n314 VTAIL.n313 9.69747
R1567 VTAIL.n42 VTAIL.n41 9.69747
R1568 VTAIL.n62 VTAIL.n61 9.69747
R1569 VTAIL.n233 VTAIL.n232 9.69747
R1570 VTAIL.n213 VTAIL.n212 9.69747
R1571 VTAIL.n149 VTAIL.n148 9.69747
R1572 VTAIL.n129 VTAIL.n128 9.69747
R1573 VTAIL.n334 VTAIL.n333 9.45567
R1574 VTAIL.n82 VTAIL.n81 9.45567
R1575 VTAIL.n252 VTAIL.n251 9.45567
R1576 VTAIL.n168 VTAIL.n167 9.45567
R1577 VTAIL.n333 VTAIL.n332 9.3005
R1578 VTAIL.n256 VTAIL.n255 9.3005
R1579 VTAIL.n301 VTAIL.n300 9.3005
R1580 VTAIL.n299 VTAIL.n298 9.3005
R1581 VTAIL.n272 VTAIL.n271 9.3005
R1582 VTAIL.n293 VTAIL.n292 9.3005
R1583 VTAIL.n291 VTAIL.n290 9.3005
R1584 VTAIL.n276 VTAIL.n275 9.3005
R1585 VTAIL.n285 VTAIL.n284 9.3005
R1586 VTAIL.n283 VTAIL.n282 9.3005
R1587 VTAIL.n268 VTAIL.n267 9.3005
R1588 VTAIL.n307 VTAIL.n306 9.3005
R1589 VTAIL.n309 VTAIL.n308 9.3005
R1590 VTAIL.n264 VTAIL.n263 9.3005
R1591 VTAIL.n315 VTAIL.n314 9.3005
R1592 VTAIL.n317 VTAIL.n316 9.3005
R1593 VTAIL.n260 VTAIL.n259 9.3005
R1594 VTAIL.n324 VTAIL.n323 9.3005
R1595 VTAIL.n326 VTAIL.n325 9.3005
R1596 VTAIL.n81 VTAIL.n80 9.3005
R1597 VTAIL.n4 VTAIL.n3 9.3005
R1598 VTAIL.n49 VTAIL.n48 9.3005
R1599 VTAIL.n47 VTAIL.n46 9.3005
R1600 VTAIL.n20 VTAIL.n19 9.3005
R1601 VTAIL.n41 VTAIL.n40 9.3005
R1602 VTAIL.n39 VTAIL.n38 9.3005
R1603 VTAIL.n24 VTAIL.n23 9.3005
R1604 VTAIL.n33 VTAIL.n32 9.3005
R1605 VTAIL.n31 VTAIL.n30 9.3005
R1606 VTAIL.n16 VTAIL.n15 9.3005
R1607 VTAIL.n55 VTAIL.n54 9.3005
R1608 VTAIL.n57 VTAIL.n56 9.3005
R1609 VTAIL.n12 VTAIL.n11 9.3005
R1610 VTAIL.n63 VTAIL.n62 9.3005
R1611 VTAIL.n65 VTAIL.n64 9.3005
R1612 VTAIL.n8 VTAIL.n7 9.3005
R1613 VTAIL.n72 VTAIL.n71 9.3005
R1614 VTAIL.n74 VTAIL.n73 9.3005
R1615 VTAIL.n226 VTAIL.n225 9.3005
R1616 VTAIL.n228 VTAIL.n227 9.3005
R1617 VTAIL.n183 VTAIL.n182 9.3005
R1618 VTAIL.n234 VTAIL.n233 9.3005
R1619 VTAIL.n236 VTAIL.n235 9.3005
R1620 VTAIL.n178 VTAIL.n177 9.3005
R1621 VTAIL.n242 VTAIL.n241 9.3005
R1622 VTAIL.n244 VTAIL.n243 9.3005
R1623 VTAIL.n251 VTAIL.n250 9.3005
R1624 VTAIL.n174 VTAIL.n173 9.3005
R1625 VTAIL.n187 VTAIL.n186 9.3005
R1626 VTAIL.n220 VTAIL.n219 9.3005
R1627 VTAIL.n218 VTAIL.n217 9.3005
R1628 VTAIL.n191 VTAIL.n190 9.3005
R1629 VTAIL.n212 VTAIL.n211 9.3005
R1630 VTAIL.n210 VTAIL.n209 9.3005
R1631 VTAIL.n195 VTAIL.n194 9.3005
R1632 VTAIL.n204 VTAIL.n203 9.3005
R1633 VTAIL.n202 VTAIL.n201 9.3005
R1634 VTAIL.n142 VTAIL.n141 9.3005
R1635 VTAIL.n144 VTAIL.n143 9.3005
R1636 VTAIL.n99 VTAIL.n98 9.3005
R1637 VTAIL.n150 VTAIL.n149 9.3005
R1638 VTAIL.n152 VTAIL.n151 9.3005
R1639 VTAIL.n94 VTAIL.n93 9.3005
R1640 VTAIL.n158 VTAIL.n157 9.3005
R1641 VTAIL.n160 VTAIL.n159 9.3005
R1642 VTAIL.n167 VTAIL.n166 9.3005
R1643 VTAIL.n90 VTAIL.n89 9.3005
R1644 VTAIL.n103 VTAIL.n102 9.3005
R1645 VTAIL.n136 VTAIL.n135 9.3005
R1646 VTAIL.n134 VTAIL.n133 9.3005
R1647 VTAIL.n107 VTAIL.n106 9.3005
R1648 VTAIL.n128 VTAIL.n127 9.3005
R1649 VTAIL.n126 VTAIL.n125 9.3005
R1650 VTAIL.n111 VTAIL.n110 9.3005
R1651 VTAIL.n120 VTAIL.n119 9.3005
R1652 VTAIL.n118 VTAIL.n117 9.3005
R1653 VTAIL.n297 VTAIL.n272 8.92171
R1654 VTAIL.n310 VTAIL.n264 8.92171
R1655 VTAIL.n45 VTAIL.n20 8.92171
R1656 VTAIL.n58 VTAIL.n12 8.92171
R1657 VTAIL.n229 VTAIL.n183 8.92171
R1658 VTAIL.n216 VTAIL.n191 8.92171
R1659 VTAIL.n145 VTAIL.n99 8.92171
R1660 VTAIL.n132 VTAIL.n107 8.92171
R1661 VTAIL.n298 VTAIL.n270 8.14595
R1662 VTAIL.n309 VTAIL.n266 8.14595
R1663 VTAIL.n46 VTAIL.n18 8.14595
R1664 VTAIL.n57 VTAIL.n14 8.14595
R1665 VTAIL.n228 VTAIL.n185 8.14595
R1666 VTAIL.n217 VTAIL.n189 8.14595
R1667 VTAIL.n144 VTAIL.n101 8.14595
R1668 VTAIL.n133 VTAIL.n105 8.14595
R1669 VTAIL.n302 VTAIL.n301 7.3702
R1670 VTAIL.n306 VTAIL.n305 7.3702
R1671 VTAIL.n50 VTAIL.n49 7.3702
R1672 VTAIL.n54 VTAIL.n53 7.3702
R1673 VTAIL.n225 VTAIL.n224 7.3702
R1674 VTAIL.n221 VTAIL.n220 7.3702
R1675 VTAIL.n141 VTAIL.n140 7.3702
R1676 VTAIL.n137 VTAIL.n136 7.3702
R1677 VTAIL.n302 VTAIL.n268 6.59444
R1678 VTAIL.n305 VTAIL.n268 6.59444
R1679 VTAIL.n50 VTAIL.n16 6.59444
R1680 VTAIL.n53 VTAIL.n16 6.59444
R1681 VTAIL.n224 VTAIL.n187 6.59444
R1682 VTAIL.n221 VTAIL.n187 6.59444
R1683 VTAIL.n140 VTAIL.n103 6.59444
R1684 VTAIL.n137 VTAIL.n103 6.59444
R1685 VTAIL.n301 VTAIL.n270 5.81868
R1686 VTAIL.n306 VTAIL.n266 5.81868
R1687 VTAIL.n49 VTAIL.n18 5.81868
R1688 VTAIL.n54 VTAIL.n14 5.81868
R1689 VTAIL.n225 VTAIL.n185 5.81868
R1690 VTAIL.n220 VTAIL.n189 5.81868
R1691 VTAIL.n141 VTAIL.n101 5.81868
R1692 VTAIL.n136 VTAIL.n105 5.81868
R1693 VTAIL.n298 VTAIL.n297 5.04292
R1694 VTAIL.n310 VTAIL.n309 5.04292
R1695 VTAIL.n46 VTAIL.n45 5.04292
R1696 VTAIL.n58 VTAIL.n57 5.04292
R1697 VTAIL.n229 VTAIL.n228 5.04292
R1698 VTAIL.n217 VTAIL.n216 5.04292
R1699 VTAIL.n145 VTAIL.n144 5.04292
R1700 VTAIL.n133 VTAIL.n132 5.04292
R1701 VTAIL.n202 VTAIL.n198 4.38563
R1702 VTAIL.n118 VTAIL.n114 4.38563
R1703 VTAIL.n283 VTAIL.n279 4.38563
R1704 VTAIL.n31 VTAIL.n27 4.38563
R1705 VTAIL.n294 VTAIL.n272 4.26717
R1706 VTAIL.n313 VTAIL.n264 4.26717
R1707 VTAIL.n42 VTAIL.n20 4.26717
R1708 VTAIL.n61 VTAIL.n12 4.26717
R1709 VTAIL.n232 VTAIL.n183 4.26717
R1710 VTAIL.n213 VTAIL.n191 4.26717
R1711 VTAIL.n148 VTAIL.n99 4.26717
R1712 VTAIL.n129 VTAIL.n107 4.26717
R1713 VTAIL.n293 VTAIL.n274 3.49141
R1714 VTAIL.n314 VTAIL.n262 3.49141
R1715 VTAIL.n41 VTAIL.n22 3.49141
R1716 VTAIL.n62 VTAIL.n10 3.49141
R1717 VTAIL.n233 VTAIL.n181 3.49141
R1718 VTAIL.n212 VTAIL.n193 3.49141
R1719 VTAIL.n149 VTAIL.n97 3.49141
R1720 VTAIL.n128 VTAIL.n109 3.49141
R1721 VTAIL.n290 VTAIL.n289 2.71565
R1722 VTAIL.n318 VTAIL.n317 2.71565
R1723 VTAIL.n38 VTAIL.n37 2.71565
R1724 VTAIL.n66 VTAIL.n65 2.71565
R1725 VTAIL.n237 VTAIL.n236 2.71565
R1726 VTAIL.n209 VTAIL.n208 2.71565
R1727 VTAIL.n153 VTAIL.n152 2.71565
R1728 VTAIL.n125 VTAIL.n124 2.71565
R1729 VTAIL.n286 VTAIL.n276 1.93989
R1730 VTAIL.n322 VTAIL.n260 1.93989
R1731 VTAIL.n334 VTAIL.n254 1.93989
R1732 VTAIL.n34 VTAIL.n24 1.93989
R1733 VTAIL.n70 VTAIL.n8 1.93989
R1734 VTAIL.n82 VTAIL.n2 1.93989
R1735 VTAIL.n252 VTAIL.n172 1.93989
R1736 VTAIL.n240 VTAIL.n178 1.93989
R1737 VTAIL.n205 VTAIL.n195 1.93989
R1738 VTAIL.n168 VTAIL.n88 1.93989
R1739 VTAIL.n156 VTAIL.n94 1.93989
R1740 VTAIL.n121 VTAIL.n111 1.93989
R1741 VTAIL.n0 VTAIL.t6 1.35204
R1742 VTAIL.n0 VTAIL.t8 1.35204
R1743 VTAIL.n84 VTAIL.t11 1.35204
R1744 VTAIL.n84 VTAIL.t1 1.35204
R1745 VTAIL.n170 VTAIL.t3 1.35204
R1746 VTAIL.n170 VTAIL.t0 1.35204
R1747 VTAIL.n86 VTAIL.t9 1.35204
R1748 VTAIL.n86 VTAIL.t7 1.35204
R1749 VTAIL.n285 VTAIL.n278 1.16414
R1750 VTAIL.n323 VTAIL.n258 1.16414
R1751 VTAIL.n332 VTAIL.n331 1.16414
R1752 VTAIL.n33 VTAIL.n26 1.16414
R1753 VTAIL.n71 VTAIL.n6 1.16414
R1754 VTAIL.n80 VTAIL.n79 1.16414
R1755 VTAIL.n250 VTAIL.n249 1.16414
R1756 VTAIL.n241 VTAIL.n176 1.16414
R1757 VTAIL.n204 VTAIL.n197 1.16414
R1758 VTAIL.n166 VTAIL.n165 1.16414
R1759 VTAIL.n157 VTAIL.n92 1.16414
R1760 VTAIL.n120 VTAIL.n113 1.16414
R1761 VTAIL.n169 VTAIL.n87 1.06947
R1762 VTAIL.n253 VTAIL.n171 1.06947
R1763 VTAIL.n85 VTAIL.n83 1.06947
R1764 VTAIL.n171 VTAIL.n169 1.00481
R1765 VTAIL.n83 VTAIL.n1 1.00481
R1766 VTAIL VTAIL.n335 0.744035
R1767 VTAIL.n282 VTAIL.n281 0.388379
R1768 VTAIL.n327 VTAIL.n326 0.388379
R1769 VTAIL.n328 VTAIL.n256 0.388379
R1770 VTAIL.n30 VTAIL.n29 0.388379
R1771 VTAIL.n75 VTAIL.n74 0.388379
R1772 VTAIL.n76 VTAIL.n4 0.388379
R1773 VTAIL.n246 VTAIL.n174 0.388379
R1774 VTAIL.n245 VTAIL.n244 0.388379
R1775 VTAIL.n201 VTAIL.n200 0.388379
R1776 VTAIL.n162 VTAIL.n90 0.388379
R1777 VTAIL.n161 VTAIL.n160 0.388379
R1778 VTAIL.n117 VTAIL.n116 0.388379
R1779 VTAIL VTAIL.n1 0.325931
R1780 VTAIL.n284 VTAIL.n283 0.155672
R1781 VTAIL.n284 VTAIL.n275 0.155672
R1782 VTAIL.n291 VTAIL.n275 0.155672
R1783 VTAIL.n292 VTAIL.n291 0.155672
R1784 VTAIL.n292 VTAIL.n271 0.155672
R1785 VTAIL.n299 VTAIL.n271 0.155672
R1786 VTAIL.n300 VTAIL.n299 0.155672
R1787 VTAIL.n300 VTAIL.n267 0.155672
R1788 VTAIL.n307 VTAIL.n267 0.155672
R1789 VTAIL.n308 VTAIL.n307 0.155672
R1790 VTAIL.n308 VTAIL.n263 0.155672
R1791 VTAIL.n315 VTAIL.n263 0.155672
R1792 VTAIL.n316 VTAIL.n315 0.155672
R1793 VTAIL.n316 VTAIL.n259 0.155672
R1794 VTAIL.n324 VTAIL.n259 0.155672
R1795 VTAIL.n325 VTAIL.n324 0.155672
R1796 VTAIL.n325 VTAIL.n255 0.155672
R1797 VTAIL.n333 VTAIL.n255 0.155672
R1798 VTAIL.n32 VTAIL.n31 0.155672
R1799 VTAIL.n32 VTAIL.n23 0.155672
R1800 VTAIL.n39 VTAIL.n23 0.155672
R1801 VTAIL.n40 VTAIL.n39 0.155672
R1802 VTAIL.n40 VTAIL.n19 0.155672
R1803 VTAIL.n47 VTAIL.n19 0.155672
R1804 VTAIL.n48 VTAIL.n47 0.155672
R1805 VTAIL.n48 VTAIL.n15 0.155672
R1806 VTAIL.n55 VTAIL.n15 0.155672
R1807 VTAIL.n56 VTAIL.n55 0.155672
R1808 VTAIL.n56 VTAIL.n11 0.155672
R1809 VTAIL.n63 VTAIL.n11 0.155672
R1810 VTAIL.n64 VTAIL.n63 0.155672
R1811 VTAIL.n64 VTAIL.n7 0.155672
R1812 VTAIL.n72 VTAIL.n7 0.155672
R1813 VTAIL.n73 VTAIL.n72 0.155672
R1814 VTAIL.n73 VTAIL.n3 0.155672
R1815 VTAIL.n81 VTAIL.n3 0.155672
R1816 VTAIL.n251 VTAIL.n173 0.155672
R1817 VTAIL.n243 VTAIL.n173 0.155672
R1818 VTAIL.n243 VTAIL.n242 0.155672
R1819 VTAIL.n242 VTAIL.n177 0.155672
R1820 VTAIL.n235 VTAIL.n177 0.155672
R1821 VTAIL.n235 VTAIL.n234 0.155672
R1822 VTAIL.n234 VTAIL.n182 0.155672
R1823 VTAIL.n227 VTAIL.n182 0.155672
R1824 VTAIL.n227 VTAIL.n226 0.155672
R1825 VTAIL.n226 VTAIL.n186 0.155672
R1826 VTAIL.n219 VTAIL.n186 0.155672
R1827 VTAIL.n219 VTAIL.n218 0.155672
R1828 VTAIL.n218 VTAIL.n190 0.155672
R1829 VTAIL.n211 VTAIL.n190 0.155672
R1830 VTAIL.n211 VTAIL.n210 0.155672
R1831 VTAIL.n210 VTAIL.n194 0.155672
R1832 VTAIL.n203 VTAIL.n194 0.155672
R1833 VTAIL.n203 VTAIL.n202 0.155672
R1834 VTAIL.n167 VTAIL.n89 0.155672
R1835 VTAIL.n159 VTAIL.n89 0.155672
R1836 VTAIL.n159 VTAIL.n158 0.155672
R1837 VTAIL.n158 VTAIL.n93 0.155672
R1838 VTAIL.n151 VTAIL.n93 0.155672
R1839 VTAIL.n151 VTAIL.n150 0.155672
R1840 VTAIL.n150 VTAIL.n98 0.155672
R1841 VTAIL.n143 VTAIL.n98 0.155672
R1842 VTAIL.n143 VTAIL.n142 0.155672
R1843 VTAIL.n142 VTAIL.n102 0.155672
R1844 VTAIL.n135 VTAIL.n102 0.155672
R1845 VTAIL.n135 VTAIL.n134 0.155672
R1846 VTAIL.n134 VTAIL.n106 0.155672
R1847 VTAIL.n127 VTAIL.n106 0.155672
R1848 VTAIL.n127 VTAIL.n126 0.155672
R1849 VTAIL.n126 VTAIL.n110 0.155672
R1850 VTAIL.n119 VTAIL.n110 0.155672
R1851 VTAIL.n119 VTAIL.n118 0.155672
R1852 VDD2.n159 VDD2.n83 289.615
R1853 VDD2.n76 VDD2.n0 289.615
R1854 VDD2.n160 VDD2.n159 185
R1855 VDD2.n158 VDD2.n157 185
R1856 VDD2.n156 VDD2.n86 185
R1857 VDD2.n90 VDD2.n87 185
R1858 VDD2.n151 VDD2.n150 185
R1859 VDD2.n149 VDD2.n148 185
R1860 VDD2.n92 VDD2.n91 185
R1861 VDD2.n143 VDD2.n142 185
R1862 VDD2.n141 VDD2.n140 185
R1863 VDD2.n96 VDD2.n95 185
R1864 VDD2.n135 VDD2.n134 185
R1865 VDD2.n133 VDD2.n132 185
R1866 VDD2.n100 VDD2.n99 185
R1867 VDD2.n127 VDD2.n126 185
R1868 VDD2.n125 VDD2.n124 185
R1869 VDD2.n104 VDD2.n103 185
R1870 VDD2.n119 VDD2.n118 185
R1871 VDD2.n117 VDD2.n116 185
R1872 VDD2.n108 VDD2.n107 185
R1873 VDD2.n111 VDD2.n110 185
R1874 VDD2.n27 VDD2.n26 185
R1875 VDD2.n24 VDD2.n23 185
R1876 VDD2.n33 VDD2.n32 185
R1877 VDD2.n35 VDD2.n34 185
R1878 VDD2.n20 VDD2.n19 185
R1879 VDD2.n41 VDD2.n40 185
R1880 VDD2.n43 VDD2.n42 185
R1881 VDD2.n16 VDD2.n15 185
R1882 VDD2.n49 VDD2.n48 185
R1883 VDD2.n51 VDD2.n50 185
R1884 VDD2.n12 VDD2.n11 185
R1885 VDD2.n57 VDD2.n56 185
R1886 VDD2.n59 VDD2.n58 185
R1887 VDD2.n8 VDD2.n7 185
R1888 VDD2.n65 VDD2.n64 185
R1889 VDD2.n68 VDD2.n67 185
R1890 VDD2.n66 VDD2.n4 185
R1891 VDD2.n73 VDD2.n3 185
R1892 VDD2.n75 VDD2.n74 185
R1893 VDD2.n77 VDD2.n76 185
R1894 VDD2.t1 VDD2.n109 147.659
R1895 VDD2.t4 VDD2.n25 147.659
R1896 VDD2.n159 VDD2.n158 104.615
R1897 VDD2.n158 VDD2.n86 104.615
R1898 VDD2.n90 VDD2.n86 104.615
R1899 VDD2.n150 VDD2.n90 104.615
R1900 VDD2.n150 VDD2.n149 104.615
R1901 VDD2.n149 VDD2.n91 104.615
R1902 VDD2.n142 VDD2.n91 104.615
R1903 VDD2.n142 VDD2.n141 104.615
R1904 VDD2.n141 VDD2.n95 104.615
R1905 VDD2.n134 VDD2.n95 104.615
R1906 VDD2.n134 VDD2.n133 104.615
R1907 VDD2.n133 VDD2.n99 104.615
R1908 VDD2.n126 VDD2.n99 104.615
R1909 VDD2.n126 VDD2.n125 104.615
R1910 VDD2.n125 VDD2.n103 104.615
R1911 VDD2.n118 VDD2.n103 104.615
R1912 VDD2.n118 VDD2.n117 104.615
R1913 VDD2.n117 VDD2.n107 104.615
R1914 VDD2.n110 VDD2.n107 104.615
R1915 VDD2.n26 VDD2.n23 104.615
R1916 VDD2.n33 VDD2.n23 104.615
R1917 VDD2.n34 VDD2.n33 104.615
R1918 VDD2.n34 VDD2.n19 104.615
R1919 VDD2.n41 VDD2.n19 104.615
R1920 VDD2.n42 VDD2.n41 104.615
R1921 VDD2.n42 VDD2.n15 104.615
R1922 VDD2.n49 VDD2.n15 104.615
R1923 VDD2.n50 VDD2.n49 104.615
R1924 VDD2.n50 VDD2.n11 104.615
R1925 VDD2.n57 VDD2.n11 104.615
R1926 VDD2.n58 VDD2.n57 104.615
R1927 VDD2.n58 VDD2.n7 104.615
R1928 VDD2.n65 VDD2.n7 104.615
R1929 VDD2.n67 VDD2.n65 104.615
R1930 VDD2.n67 VDD2.n66 104.615
R1931 VDD2.n66 VDD2.n3 104.615
R1932 VDD2.n75 VDD2.n3 104.615
R1933 VDD2.n76 VDD2.n75 104.615
R1934 VDD2.n82 VDD2.n81 61.3267
R1935 VDD2 VDD2.n165 61.3239
R1936 VDD2.n110 VDD2.t1 52.3082
R1937 VDD2.n26 VDD2.t4 52.3082
R1938 VDD2.n82 VDD2.n80 49.8045
R1939 VDD2.n164 VDD2.n163 49.0581
R1940 VDD2.n164 VDD2.n82 39.8187
R1941 VDD2.n111 VDD2.n109 15.6677
R1942 VDD2.n27 VDD2.n25 15.6677
R1943 VDD2.n157 VDD2.n156 13.1884
R1944 VDD2.n74 VDD2.n73 13.1884
R1945 VDD2.n160 VDD2.n85 12.8005
R1946 VDD2.n155 VDD2.n87 12.8005
R1947 VDD2.n112 VDD2.n108 12.8005
R1948 VDD2.n28 VDD2.n24 12.8005
R1949 VDD2.n72 VDD2.n4 12.8005
R1950 VDD2.n77 VDD2.n2 12.8005
R1951 VDD2.n161 VDD2.n83 12.0247
R1952 VDD2.n152 VDD2.n151 12.0247
R1953 VDD2.n116 VDD2.n115 12.0247
R1954 VDD2.n32 VDD2.n31 12.0247
R1955 VDD2.n69 VDD2.n68 12.0247
R1956 VDD2.n78 VDD2.n0 12.0247
R1957 VDD2.n148 VDD2.n89 11.249
R1958 VDD2.n119 VDD2.n106 11.249
R1959 VDD2.n35 VDD2.n22 11.249
R1960 VDD2.n64 VDD2.n6 11.249
R1961 VDD2.n147 VDD2.n92 10.4732
R1962 VDD2.n120 VDD2.n104 10.4732
R1963 VDD2.n36 VDD2.n20 10.4732
R1964 VDD2.n63 VDD2.n8 10.4732
R1965 VDD2.n144 VDD2.n143 9.69747
R1966 VDD2.n124 VDD2.n123 9.69747
R1967 VDD2.n40 VDD2.n39 9.69747
R1968 VDD2.n60 VDD2.n59 9.69747
R1969 VDD2.n163 VDD2.n162 9.45567
R1970 VDD2.n80 VDD2.n79 9.45567
R1971 VDD2.n137 VDD2.n136 9.3005
R1972 VDD2.n139 VDD2.n138 9.3005
R1973 VDD2.n94 VDD2.n93 9.3005
R1974 VDD2.n145 VDD2.n144 9.3005
R1975 VDD2.n147 VDD2.n146 9.3005
R1976 VDD2.n89 VDD2.n88 9.3005
R1977 VDD2.n153 VDD2.n152 9.3005
R1978 VDD2.n155 VDD2.n154 9.3005
R1979 VDD2.n162 VDD2.n161 9.3005
R1980 VDD2.n85 VDD2.n84 9.3005
R1981 VDD2.n98 VDD2.n97 9.3005
R1982 VDD2.n131 VDD2.n130 9.3005
R1983 VDD2.n129 VDD2.n128 9.3005
R1984 VDD2.n102 VDD2.n101 9.3005
R1985 VDD2.n123 VDD2.n122 9.3005
R1986 VDD2.n121 VDD2.n120 9.3005
R1987 VDD2.n106 VDD2.n105 9.3005
R1988 VDD2.n115 VDD2.n114 9.3005
R1989 VDD2.n113 VDD2.n112 9.3005
R1990 VDD2.n79 VDD2.n78 9.3005
R1991 VDD2.n2 VDD2.n1 9.3005
R1992 VDD2.n47 VDD2.n46 9.3005
R1993 VDD2.n45 VDD2.n44 9.3005
R1994 VDD2.n18 VDD2.n17 9.3005
R1995 VDD2.n39 VDD2.n38 9.3005
R1996 VDD2.n37 VDD2.n36 9.3005
R1997 VDD2.n22 VDD2.n21 9.3005
R1998 VDD2.n31 VDD2.n30 9.3005
R1999 VDD2.n29 VDD2.n28 9.3005
R2000 VDD2.n14 VDD2.n13 9.3005
R2001 VDD2.n53 VDD2.n52 9.3005
R2002 VDD2.n55 VDD2.n54 9.3005
R2003 VDD2.n10 VDD2.n9 9.3005
R2004 VDD2.n61 VDD2.n60 9.3005
R2005 VDD2.n63 VDD2.n62 9.3005
R2006 VDD2.n6 VDD2.n5 9.3005
R2007 VDD2.n70 VDD2.n69 9.3005
R2008 VDD2.n72 VDD2.n71 9.3005
R2009 VDD2.n140 VDD2.n94 8.92171
R2010 VDD2.n127 VDD2.n102 8.92171
R2011 VDD2.n43 VDD2.n18 8.92171
R2012 VDD2.n56 VDD2.n10 8.92171
R2013 VDD2.n139 VDD2.n96 8.14595
R2014 VDD2.n128 VDD2.n100 8.14595
R2015 VDD2.n44 VDD2.n16 8.14595
R2016 VDD2.n55 VDD2.n12 8.14595
R2017 VDD2.n136 VDD2.n135 7.3702
R2018 VDD2.n132 VDD2.n131 7.3702
R2019 VDD2.n48 VDD2.n47 7.3702
R2020 VDD2.n52 VDD2.n51 7.3702
R2021 VDD2.n135 VDD2.n98 6.59444
R2022 VDD2.n132 VDD2.n98 6.59444
R2023 VDD2.n48 VDD2.n14 6.59444
R2024 VDD2.n51 VDD2.n14 6.59444
R2025 VDD2.n136 VDD2.n96 5.81868
R2026 VDD2.n131 VDD2.n100 5.81868
R2027 VDD2.n47 VDD2.n16 5.81868
R2028 VDD2.n52 VDD2.n12 5.81868
R2029 VDD2.n140 VDD2.n139 5.04292
R2030 VDD2.n128 VDD2.n127 5.04292
R2031 VDD2.n44 VDD2.n43 5.04292
R2032 VDD2.n56 VDD2.n55 5.04292
R2033 VDD2.n113 VDD2.n109 4.38563
R2034 VDD2.n29 VDD2.n25 4.38563
R2035 VDD2.n143 VDD2.n94 4.26717
R2036 VDD2.n124 VDD2.n102 4.26717
R2037 VDD2.n40 VDD2.n18 4.26717
R2038 VDD2.n59 VDD2.n10 4.26717
R2039 VDD2.n144 VDD2.n92 3.49141
R2040 VDD2.n123 VDD2.n104 3.49141
R2041 VDD2.n39 VDD2.n20 3.49141
R2042 VDD2.n60 VDD2.n8 3.49141
R2043 VDD2.n148 VDD2.n147 2.71565
R2044 VDD2.n120 VDD2.n119 2.71565
R2045 VDD2.n36 VDD2.n35 2.71565
R2046 VDD2.n64 VDD2.n63 2.71565
R2047 VDD2.n163 VDD2.n83 1.93989
R2048 VDD2.n151 VDD2.n89 1.93989
R2049 VDD2.n116 VDD2.n106 1.93989
R2050 VDD2.n32 VDD2.n22 1.93989
R2051 VDD2.n68 VDD2.n6 1.93989
R2052 VDD2.n80 VDD2.n0 1.93989
R2053 VDD2.n165 VDD2.t3 1.35204
R2054 VDD2.n165 VDD2.t0 1.35204
R2055 VDD2.n81 VDD2.t2 1.35204
R2056 VDD2.n81 VDD2.t5 1.35204
R2057 VDD2.n161 VDD2.n160 1.16414
R2058 VDD2.n152 VDD2.n87 1.16414
R2059 VDD2.n115 VDD2.n108 1.16414
R2060 VDD2.n31 VDD2.n24 1.16414
R2061 VDD2.n69 VDD2.n4 1.16414
R2062 VDD2.n78 VDD2.n77 1.16414
R2063 VDD2 VDD2.n164 0.860414
R2064 VDD2.n157 VDD2.n85 0.388379
R2065 VDD2.n156 VDD2.n155 0.388379
R2066 VDD2.n112 VDD2.n111 0.388379
R2067 VDD2.n28 VDD2.n27 0.388379
R2068 VDD2.n73 VDD2.n72 0.388379
R2069 VDD2.n74 VDD2.n2 0.388379
R2070 VDD2.n162 VDD2.n84 0.155672
R2071 VDD2.n154 VDD2.n84 0.155672
R2072 VDD2.n154 VDD2.n153 0.155672
R2073 VDD2.n153 VDD2.n88 0.155672
R2074 VDD2.n146 VDD2.n88 0.155672
R2075 VDD2.n146 VDD2.n145 0.155672
R2076 VDD2.n145 VDD2.n93 0.155672
R2077 VDD2.n138 VDD2.n93 0.155672
R2078 VDD2.n138 VDD2.n137 0.155672
R2079 VDD2.n137 VDD2.n97 0.155672
R2080 VDD2.n130 VDD2.n97 0.155672
R2081 VDD2.n130 VDD2.n129 0.155672
R2082 VDD2.n129 VDD2.n101 0.155672
R2083 VDD2.n122 VDD2.n101 0.155672
R2084 VDD2.n122 VDD2.n121 0.155672
R2085 VDD2.n121 VDD2.n105 0.155672
R2086 VDD2.n114 VDD2.n105 0.155672
R2087 VDD2.n114 VDD2.n113 0.155672
R2088 VDD2.n30 VDD2.n29 0.155672
R2089 VDD2.n30 VDD2.n21 0.155672
R2090 VDD2.n37 VDD2.n21 0.155672
R2091 VDD2.n38 VDD2.n37 0.155672
R2092 VDD2.n38 VDD2.n17 0.155672
R2093 VDD2.n45 VDD2.n17 0.155672
R2094 VDD2.n46 VDD2.n45 0.155672
R2095 VDD2.n46 VDD2.n13 0.155672
R2096 VDD2.n53 VDD2.n13 0.155672
R2097 VDD2.n54 VDD2.n53 0.155672
R2098 VDD2.n54 VDD2.n9 0.155672
R2099 VDD2.n61 VDD2.n9 0.155672
R2100 VDD2.n62 VDD2.n61 0.155672
R2101 VDD2.n62 VDD2.n5 0.155672
R2102 VDD2.n70 VDD2.n5 0.155672
R2103 VDD2.n71 VDD2.n70 0.155672
R2104 VDD2.n71 VDD2.n1 0.155672
R2105 VDD2.n79 VDD2.n1 0.155672
R2106 VP.n5 VP.t5 448.873
R2107 VP.n12 VP.t1 431.418
R2108 VP.n19 VP.t0 431.418
R2109 VP.n9 VP.t4 431.418
R2110 VP.n1 VP.t2 387.985
R2111 VP.n4 VP.t3 387.985
R2112 VP.n20 VP.n19 161.3
R2113 VP.n7 VP.n6 161.3
R2114 VP.n8 VP.n3 161.3
R2115 VP.n10 VP.n9 161.3
R2116 VP.n18 VP.n0 161.3
R2117 VP.n17 VP.n16 161.3
R2118 VP.n15 VP.n14 161.3
R2119 VP.n13 VP.n2 161.3
R2120 VP.n12 VP.n11 161.3
R2121 VP.n14 VP.n13 53.1199
R2122 VP.n18 VP.n17 53.1199
R2123 VP.n8 VP.n7 53.1199
R2124 VP.n11 VP.n10 44.0535
R2125 VP.n6 VP.n5 43.5004
R2126 VP.n5 VP.n4 42.494
R2127 VP.n14 VP.n1 12.234
R2128 VP.n17 VP.n1 12.234
R2129 VP.n7 VP.n4 12.234
R2130 VP.n13 VP.n12 5.11262
R2131 VP.n19 VP.n18 5.11262
R2132 VP.n9 VP.n8 5.11262
R2133 VP.n6 VP.n3 0.189894
R2134 VP.n10 VP.n3 0.189894
R2135 VP.n11 VP.n2 0.189894
R2136 VP.n15 VP.n2 0.189894
R2137 VP.n16 VP.n15 0.189894
R2138 VP.n16 VP.n0 0.189894
R2139 VP.n20 VP.n0 0.189894
R2140 VP VP.n20 0.0516364
R2141 VDD1.n76 VDD1.n0 289.615
R2142 VDD1.n157 VDD1.n81 289.615
R2143 VDD1.n77 VDD1.n76 185
R2144 VDD1.n75 VDD1.n74 185
R2145 VDD1.n73 VDD1.n3 185
R2146 VDD1.n7 VDD1.n4 185
R2147 VDD1.n68 VDD1.n67 185
R2148 VDD1.n66 VDD1.n65 185
R2149 VDD1.n9 VDD1.n8 185
R2150 VDD1.n60 VDD1.n59 185
R2151 VDD1.n58 VDD1.n57 185
R2152 VDD1.n13 VDD1.n12 185
R2153 VDD1.n52 VDD1.n51 185
R2154 VDD1.n50 VDD1.n49 185
R2155 VDD1.n17 VDD1.n16 185
R2156 VDD1.n44 VDD1.n43 185
R2157 VDD1.n42 VDD1.n41 185
R2158 VDD1.n21 VDD1.n20 185
R2159 VDD1.n36 VDD1.n35 185
R2160 VDD1.n34 VDD1.n33 185
R2161 VDD1.n25 VDD1.n24 185
R2162 VDD1.n28 VDD1.n27 185
R2163 VDD1.n108 VDD1.n107 185
R2164 VDD1.n105 VDD1.n104 185
R2165 VDD1.n114 VDD1.n113 185
R2166 VDD1.n116 VDD1.n115 185
R2167 VDD1.n101 VDD1.n100 185
R2168 VDD1.n122 VDD1.n121 185
R2169 VDD1.n124 VDD1.n123 185
R2170 VDD1.n97 VDD1.n96 185
R2171 VDD1.n130 VDD1.n129 185
R2172 VDD1.n132 VDD1.n131 185
R2173 VDD1.n93 VDD1.n92 185
R2174 VDD1.n138 VDD1.n137 185
R2175 VDD1.n140 VDD1.n139 185
R2176 VDD1.n89 VDD1.n88 185
R2177 VDD1.n146 VDD1.n145 185
R2178 VDD1.n149 VDD1.n148 185
R2179 VDD1.n147 VDD1.n85 185
R2180 VDD1.n154 VDD1.n84 185
R2181 VDD1.n156 VDD1.n155 185
R2182 VDD1.n158 VDD1.n157 185
R2183 VDD1.t0 VDD1.n26 147.659
R2184 VDD1.t4 VDD1.n106 147.659
R2185 VDD1.n76 VDD1.n75 104.615
R2186 VDD1.n75 VDD1.n3 104.615
R2187 VDD1.n7 VDD1.n3 104.615
R2188 VDD1.n67 VDD1.n7 104.615
R2189 VDD1.n67 VDD1.n66 104.615
R2190 VDD1.n66 VDD1.n8 104.615
R2191 VDD1.n59 VDD1.n8 104.615
R2192 VDD1.n59 VDD1.n58 104.615
R2193 VDD1.n58 VDD1.n12 104.615
R2194 VDD1.n51 VDD1.n12 104.615
R2195 VDD1.n51 VDD1.n50 104.615
R2196 VDD1.n50 VDD1.n16 104.615
R2197 VDD1.n43 VDD1.n16 104.615
R2198 VDD1.n43 VDD1.n42 104.615
R2199 VDD1.n42 VDD1.n20 104.615
R2200 VDD1.n35 VDD1.n20 104.615
R2201 VDD1.n35 VDD1.n34 104.615
R2202 VDD1.n34 VDD1.n24 104.615
R2203 VDD1.n27 VDD1.n24 104.615
R2204 VDD1.n107 VDD1.n104 104.615
R2205 VDD1.n114 VDD1.n104 104.615
R2206 VDD1.n115 VDD1.n114 104.615
R2207 VDD1.n115 VDD1.n100 104.615
R2208 VDD1.n122 VDD1.n100 104.615
R2209 VDD1.n123 VDD1.n122 104.615
R2210 VDD1.n123 VDD1.n96 104.615
R2211 VDD1.n130 VDD1.n96 104.615
R2212 VDD1.n131 VDD1.n130 104.615
R2213 VDD1.n131 VDD1.n92 104.615
R2214 VDD1.n138 VDD1.n92 104.615
R2215 VDD1.n139 VDD1.n138 104.615
R2216 VDD1.n139 VDD1.n88 104.615
R2217 VDD1.n146 VDD1.n88 104.615
R2218 VDD1.n148 VDD1.n146 104.615
R2219 VDD1.n148 VDD1.n147 104.615
R2220 VDD1.n147 VDD1.n84 104.615
R2221 VDD1.n156 VDD1.n84 104.615
R2222 VDD1.n157 VDD1.n156 104.615
R2223 VDD1.n163 VDD1.n162 61.3267
R2224 VDD1.n165 VDD1.n164 61.1149
R2225 VDD1.n27 VDD1.t0 52.3082
R2226 VDD1.n107 VDD1.t4 52.3082
R2227 VDD1 VDD1.n80 49.918
R2228 VDD1.n163 VDD1.n161 49.8045
R2229 VDD1.n165 VDD1.n163 40.9362
R2230 VDD1.n28 VDD1.n26 15.6677
R2231 VDD1.n108 VDD1.n106 15.6677
R2232 VDD1.n74 VDD1.n73 13.1884
R2233 VDD1.n155 VDD1.n154 13.1884
R2234 VDD1.n77 VDD1.n2 12.8005
R2235 VDD1.n72 VDD1.n4 12.8005
R2236 VDD1.n29 VDD1.n25 12.8005
R2237 VDD1.n109 VDD1.n105 12.8005
R2238 VDD1.n153 VDD1.n85 12.8005
R2239 VDD1.n158 VDD1.n83 12.8005
R2240 VDD1.n78 VDD1.n0 12.0247
R2241 VDD1.n69 VDD1.n68 12.0247
R2242 VDD1.n33 VDD1.n32 12.0247
R2243 VDD1.n113 VDD1.n112 12.0247
R2244 VDD1.n150 VDD1.n149 12.0247
R2245 VDD1.n159 VDD1.n81 12.0247
R2246 VDD1.n65 VDD1.n6 11.249
R2247 VDD1.n36 VDD1.n23 11.249
R2248 VDD1.n116 VDD1.n103 11.249
R2249 VDD1.n145 VDD1.n87 11.249
R2250 VDD1.n64 VDD1.n9 10.4732
R2251 VDD1.n37 VDD1.n21 10.4732
R2252 VDD1.n117 VDD1.n101 10.4732
R2253 VDD1.n144 VDD1.n89 10.4732
R2254 VDD1.n61 VDD1.n60 9.69747
R2255 VDD1.n41 VDD1.n40 9.69747
R2256 VDD1.n121 VDD1.n120 9.69747
R2257 VDD1.n141 VDD1.n140 9.69747
R2258 VDD1.n80 VDD1.n79 9.45567
R2259 VDD1.n161 VDD1.n160 9.45567
R2260 VDD1.n54 VDD1.n53 9.3005
R2261 VDD1.n56 VDD1.n55 9.3005
R2262 VDD1.n11 VDD1.n10 9.3005
R2263 VDD1.n62 VDD1.n61 9.3005
R2264 VDD1.n64 VDD1.n63 9.3005
R2265 VDD1.n6 VDD1.n5 9.3005
R2266 VDD1.n70 VDD1.n69 9.3005
R2267 VDD1.n72 VDD1.n71 9.3005
R2268 VDD1.n79 VDD1.n78 9.3005
R2269 VDD1.n2 VDD1.n1 9.3005
R2270 VDD1.n15 VDD1.n14 9.3005
R2271 VDD1.n48 VDD1.n47 9.3005
R2272 VDD1.n46 VDD1.n45 9.3005
R2273 VDD1.n19 VDD1.n18 9.3005
R2274 VDD1.n40 VDD1.n39 9.3005
R2275 VDD1.n38 VDD1.n37 9.3005
R2276 VDD1.n23 VDD1.n22 9.3005
R2277 VDD1.n32 VDD1.n31 9.3005
R2278 VDD1.n30 VDD1.n29 9.3005
R2279 VDD1.n160 VDD1.n159 9.3005
R2280 VDD1.n83 VDD1.n82 9.3005
R2281 VDD1.n128 VDD1.n127 9.3005
R2282 VDD1.n126 VDD1.n125 9.3005
R2283 VDD1.n99 VDD1.n98 9.3005
R2284 VDD1.n120 VDD1.n119 9.3005
R2285 VDD1.n118 VDD1.n117 9.3005
R2286 VDD1.n103 VDD1.n102 9.3005
R2287 VDD1.n112 VDD1.n111 9.3005
R2288 VDD1.n110 VDD1.n109 9.3005
R2289 VDD1.n95 VDD1.n94 9.3005
R2290 VDD1.n134 VDD1.n133 9.3005
R2291 VDD1.n136 VDD1.n135 9.3005
R2292 VDD1.n91 VDD1.n90 9.3005
R2293 VDD1.n142 VDD1.n141 9.3005
R2294 VDD1.n144 VDD1.n143 9.3005
R2295 VDD1.n87 VDD1.n86 9.3005
R2296 VDD1.n151 VDD1.n150 9.3005
R2297 VDD1.n153 VDD1.n152 9.3005
R2298 VDD1.n57 VDD1.n11 8.92171
R2299 VDD1.n44 VDD1.n19 8.92171
R2300 VDD1.n124 VDD1.n99 8.92171
R2301 VDD1.n137 VDD1.n91 8.92171
R2302 VDD1.n56 VDD1.n13 8.14595
R2303 VDD1.n45 VDD1.n17 8.14595
R2304 VDD1.n125 VDD1.n97 8.14595
R2305 VDD1.n136 VDD1.n93 8.14595
R2306 VDD1.n53 VDD1.n52 7.3702
R2307 VDD1.n49 VDD1.n48 7.3702
R2308 VDD1.n129 VDD1.n128 7.3702
R2309 VDD1.n133 VDD1.n132 7.3702
R2310 VDD1.n52 VDD1.n15 6.59444
R2311 VDD1.n49 VDD1.n15 6.59444
R2312 VDD1.n129 VDD1.n95 6.59444
R2313 VDD1.n132 VDD1.n95 6.59444
R2314 VDD1.n53 VDD1.n13 5.81868
R2315 VDD1.n48 VDD1.n17 5.81868
R2316 VDD1.n128 VDD1.n97 5.81868
R2317 VDD1.n133 VDD1.n93 5.81868
R2318 VDD1.n57 VDD1.n56 5.04292
R2319 VDD1.n45 VDD1.n44 5.04292
R2320 VDD1.n125 VDD1.n124 5.04292
R2321 VDD1.n137 VDD1.n136 5.04292
R2322 VDD1.n30 VDD1.n26 4.38563
R2323 VDD1.n110 VDD1.n106 4.38563
R2324 VDD1.n60 VDD1.n11 4.26717
R2325 VDD1.n41 VDD1.n19 4.26717
R2326 VDD1.n121 VDD1.n99 4.26717
R2327 VDD1.n140 VDD1.n91 4.26717
R2328 VDD1.n61 VDD1.n9 3.49141
R2329 VDD1.n40 VDD1.n21 3.49141
R2330 VDD1.n120 VDD1.n101 3.49141
R2331 VDD1.n141 VDD1.n89 3.49141
R2332 VDD1.n65 VDD1.n64 2.71565
R2333 VDD1.n37 VDD1.n36 2.71565
R2334 VDD1.n117 VDD1.n116 2.71565
R2335 VDD1.n145 VDD1.n144 2.71565
R2336 VDD1.n80 VDD1.n0 1.93989
R2337 VDD1.n68 VDD1.n6 1.93989
R2338 VDD1.n33 VDD1.n23 1.93989
R2339 VDD1.n113 VDD1.n103 1.93989
R2340 VDD1.n149 VDD1.n87 1.93989
R2341 VDD1.n161 VDD1.n81 1.93989
R2342 VDD1.n164 VDD1.t2 1.35204
R2343 VDD1.n164 VDD1.t1 1.35204
R2344 VDD1.n162 VDD1.t3 1.35204
R2345 VDD1.n162 VDD1.t5 1.35204
R2346 VDD1.n78 VDD1.n77 1.16414
R2347 VDD1.n69 VDD1.n4 1.16414
R2348 VDD1.n32 VDD1.n25 1.16414
R2349 VDD1.n112 VDD1.n105 1.16414
R2350 VDD1.n150 VDD1.n85 1.16414
R2351 VDD1.n159 VDD1.n158 1.16414
R2352 VDD1.n74 VDD1.n2 0.388379
R2353 VDD1.n73 VDD1.n72 0.388379
R2354 VDD1.n29 VDD1.n28 0.388379
R2355 VDD1.n109 VDD1.n108 0.388379
R2356 VDD1.n154 VDD1.n153 0.388379
R2357 VDD1.n155 VDD1.n83 0.388379
R2358 VDD1 VDD1.n165 0.209552
R2359 VDD1.n79 VDD1.n1 0.155672
R2360 VDD1.n71 VDD1.n1 0.155672
R2361 VDD1.n71 VDD1.n70 0.155672
R2362 VDD1.n70 VDD1.n5 0.155672
R2363 VDD1.n63 VDD1.n5 0.155672
R2364 VDD1.n63 VDD1.n62 0.155672
R2365 VDD1.n62 VDD1.n10 0.155672
R2366 VDD1.n55 VDD1.n10 0.155672
R2367 VDD1.n55 VDD1.n54 0.155672
R2368 VDD1.n54 VDD1.n14 0.155672
R2369 VDD1.n47 VDD1.n14 0.155672
R2370 VDD1.n47 VDD1.n46 0.155672
R2371 VDD1.n46 VDD1.n18 0.155672
R2372 VDD1.n39 VDD1.n18 0.155672
R2373 VDD1.n39 VDD1.n38 0.155672
R2374 VDD1.n38 VDD1.n22 0.155672
R2375 VDD1.n31 VDD1.n22 0.155672
R2376 VDD1.n31 VDD1.n30 0.155672
R2377 VDD1.n111 VDD1.n110 0.155672
R2378 VDD1.n111 VDD1.n102 0.155672
R2379 VDD1.n118 VDD1.n102 0.155672
R2380 VDD1.n119 VDD1.n118 0.155672
R2381 VDD1.n119 VDD1.n98 0.155672
R2382 VDD1.n126 VDD1.n98 0.155672
R2383 VDD1.n127 VDD1.n126 0.155672
R2384 VDD1.n127 VDD1.n94 0.155672
R2385 VDD1.n134 VDD1.n94 0.155672
R2386 VDD1.n135 VDD1.n134 0.155672
R2387 VDD1.n135 VDD1.n90 0.155672
R2388 VDD1.n142 VDD1.n90 0.155672
R2389 VDD1.n143 VDD1.n142 0.155672
R2390 VDD1.n143 VDD1.n86 0.155672
R2391 VDD1.n151 VDD1.n86 0.155672
R2392 VDD1.n152 VDD1.n151 0.155672
R2393 VDD1.n152 VDD1.n82 0.155672
R2394 VDD1.n160 VDD1.n82 0.155672
C0 VP VTAIL 5.54927f
C1 VP VDD1 6.06057f
C2 VP VN 5.77482f
C3 VTAIL VDD2 10.656401f
C4 VDD1 VDD2 0.787847f
C5 VN VDD2 5.89838f
C6 VP VDD2 0.315699f
C7 VTAIL VDD1 10.6215f
C8 VN VTAIL 5.53463f
C9 VN VDD1 0.148417f
C10 VDD2 B 5.129645f
C11 VDD1 B 5.16428f
C12 VTAIL B 7.56524f
C13 VN B 8.54093f
C14 VP B 6.574522f
C15 VDD1.n0 B 0.028934f
C16 VDD1.n1 B 0.022651f
C17 VDD1.n2 B 0.012172f
C18 VDD1.n3 B 0.02877f
C19 VDD1.n4 B 0.012888f
C20 VDD1.n5 B 0.022651f
C21 VDD1.n6 B 0.012172f
C22 VDD1.n7 B 0.02877f
C23 VDD1.n8 B 0.02877f
C24 VDD1.n9 B 0.012888f
C25 VDD1.n10 B 0.022651f
C26 VDD1.n11 B 0.012172f
C27 VDD1.n12 B 0.02877f
C28 VDD1.n13 B 0.012888f
C29 VDD1.n14 B 0.022651f
C30 VDD1.n15 B 0.012172f
C31 VDD1.n16 B 0.02877f
C32 VDD1.n17 B 0.012888f
C33 VDD1.n18 B 0.022651f
C34 VDD1.n19 B 0.012172f
C35 VDD1.n20 B 0.02877f
C36 VDD1.n21 B 0.012888f
C37 VDD1.n22 B 0.022651f
C38 VDD1.n23 B 0.012172f
C39 VDD1.n24 B 0.02877f
C40 VDD1.n25 B 0.012888f
C41 VDD1.n26 B 0.145747f
C42 VDD1.t0 B 0.04741f
C43 VDD1.n27 B 0.021577f
C44 VDD1.n28 B 0.016995f
C45 VDD1.n29 B 0.012172f
C46 VDD1.n30 B 1.43738f
C47 VDD1.n31 B 0.022651f
C48 VDD1.n32 B 0.012172f
C49 VDD1.n33 B 0.012888f
C50 VDD1.n34 B 0.02877f
C51 VDD1.n35 B 0.02877f
C52 VDD1.n36 B 0.012888f
C53 VDD1.n37 B 0.012172f
C54 VDD1.n38 B 0.022651f
C55 VDD1.n39 B 0.022651f
C56 VDD1.n40 B 0.012172f
C57 VDD1.n41 B 0.012888f
C58 VDD1.n42 B 0.02877f
C59 VDD1.n43 B 0.02877f
C60 VDD1.n44 B 0.012888f
C61 VDD1.n45 B 0.012172f
C62 VDD1.n46 B 0.022651f
C63 VDD1.n47 B 0.022651f
C64 VDD1.n48 B 0.012172f
C65 VDD1.n49 B 0.012888f
C66 VDD1.n50 B 0.02877f
C67 VDD1.n51 B 0.02877f
C68 VDD1.n52 B 0.012888f
C69 VDD1.n53 B 0.012172f
C70 VDD1.n54 B 0.022651f
C71 VDD1.n55 B 0.022651f
C72 VDD1.n56 B 0.012172f
C73 VDD1.n57 B 0.012888f
C74 VDD1.n58 B 0.02877f
C75 VDD1.n59 B 0.02877f
C76 VDD1.n60 B 0.012888f
C77 VDD1.n61 B 0.012172f
C78 VDD1.n62 B 0.022651f
C79 VDD1.n63 B 0.022651f
C80 VDD1.n64 B 0.012172f
C81 VDD1.n65 B 0.012888f
C82 VDD1.n66 B 0.02877f
C83 VDD1.n67 B 0.02877f
C84 VDD1.n68 B 0.012888f
C85 VDD1.n69 B 0.012172f
C86 VDD1.n70 B 0.022651f
C87 VDD1.n71 B 0.022651f
C88 VDD1.n72 B 0.012172f
C89 VDD1.n73 B 0.01253f
C90 VDD1.n74 B 0.01253f
C91 VDD1.n75 B 0.02877f
C92 VDD1.n76 B 0.057146f
C93 VDD1.n77 B 0.012888f
C94 VDD1.n78 B 0.012172f
C95 VDD1.n79 B 0.052666f
C96 VDD1.n80 B 0.04893f
C97 VDD1.n81 B 0.028934f
C98 VDD1.n82 B 0.022651f
C99 VDD1.n83 B 0.012172f
C100 VDD1.n84 B 0.02877f
C101 VDD1.n85 B 0.012888f
C102 VDD1.n86 B 0.022651f
C103 VDD1.n87 B 0.012172f
C104 VDD1.n88 B 0.02877f
C105 VDD1.n89 B 0.012888f
C106 VDD1.n90 B 0.022651f
C107 VDD1.n91 B 0.012172f
C108 VDD1.n92 B 0.02877f
C109 VDD1.n93 B 0.012888f
C110 VDD1.n94 B 0.022651f
C111 VDD1.n95 B 0.012172f
C112 VDD1.n96 B 0.02877f
C113 VDD1.n97 B 0.012888f
C114 VDD1.n98 B 0.022651f
C115 VDD1.n99 B 0.012172f
C116 VDD1.n100 B 0.02877f
C117 VDD1.n101 B 0.012888f
C118 VDD1.n102 B 0.022651f
C119 VDD1.n103 B 0.012172f
C120 VDD1.n104 B 0.02877f
C121 VDD1.n105 B 0.012888f
C122 VDD1.n106 B 0.145747f
C123 VDD1.t4 B 0.04741f
C124 VDD1.n107 B 0.021577f
C125 VDD1.n108 B 0.016995f
C126 VDD1.n109 B 0.012172f
C127 VDD1.n110 B 1.43738f
C128 VDD1.n111 B 0.022651f
C129 VDD1.n112 B 0.012172f
C130 VDD1.n113 B 0.012888f
C131 VDD1.n114 B 0.02877f
C132 VDD1.n115 B 0.02877f
C133 VDD1.n116 B 0.012888f
C134 VDD1.n117 B 0.012172f
C135 VDD1.n118 B 0.022651f
C136 VDD1.n119 B 0.022651f
C137 VDD1.n120 B 0.012172f
C138 VDD1.n121 B 0.012888f
C139 VDD1.n122 B 0.02877f
C140 VDD1.n123 B 0.02877f
C141 VDD1.n124 B 0.012888f
C142 VDD1.n125 B 0.012172f
C143 VDD1.n126 B 0.022651f
C144 VDD1.n127 B 0.022651f
C145 VDD1.n128 B 0.012172f
C146 VDD1.n129 B 0.012888f
C147 VDD1.n130 B 0.02877f
C148 VDD1.n131 B 0.02877f
C149 VDD1.n132 B 0.012888f
C150 VDD1.n133 B 0.012172f
C151 VDD1.n134 B 0.022651f
C152 VDD1.n135 B 0.022651f
C153 VDD1.n136 B 0.012172f
C154 VDD1.n137 B 0.012888f
C155 VDD1.n138 B 0.02877f
C156 VDD1.n139 B 0.02877f
C157 VDD1.n140 B 0.012888f
C158 VDD1.n141 B 0.012172f
C159 VDD1.n142 B 0.022651f
C160 VDD1.n143 B 0.022651f
C161 VDD1.n144 B 0.012172f
C162 VDD1.n145 B 0.012888f
C163 VDD1.n146 B 0.02877f
C164 VDD1.n147 B 0.02877f
C165 VDD1.n148 B 0.02877f
C166 VDD1.n149 B 0.012888f
C167 VDD1.n150 B 0.012172f
C168 VDD1.n151 B 0.022651f
C169 VDD1.n152 B 0.022651f
C170 VDD1.n153 B 0.012172f
C171 VDD1.n154 B 0.01253f
C172 VDD1.n155 B 0.01253f
C173 VDD1.n156 B 0.02877f
C174 VDD1.n157 B 0.057146f
C175 VDD1.n158 B 0.012888f
C176 VDD1.n159 B 0.012172f
C177 VDD1.n160 B 0.052666f
C178 VDD1.n161 B 0.048578f
C179 VDD1.t3 B 0.262228f
C180 VDD1.t5 B 0.262228f
C181 VDD1.n162 B 2.36883f
C182 VDD1.n163 B 1.98257f
C183 VDD1.t2 B 0.262228f
C184 VDD1.t1 B 0.262228f
C185 VDD1.n164 B 2.36783f
C186 VDD1.n165 B 2.27924f
C187 VP.n0 B 0.04179f
C188 VP.t2 B 1.52579f
C189 VP.n1 B 0.558891f
C190 VP.n2 B 0.04179f
C191 VP.n3 B 0.04179f
C192 VP.t4 B 1.58405f
C193 VP.t3 B 1.52579f
C194 VP.n4 B 0.59845f
C195 VP.t5 B 1.60799f
C196 VP.n5 B 0.610217f
C197 VP.n6 B 0.176336f
C198 VP.n7 B 0.054923f
C199 VP.n8 B 0.013895f
C200 VP.n9 B 0.604028f
C201 VP.n10 B 1.86547f
C202 VP.n11 B 1.89957f
C203 VP.t1 B 1.58405f
C204 VP.n12 B 0.604028f
C205 VP.n13 B 0.013895f
C206 VP.n14 B 0.054923f
C207 VP.n15 B 0.04179f
C208 VP.n16 B 0.04179f
C209 VP.n17 B 0.054923f
C210 VP.n18 B 0.013895f
C211 VP.t0 B 1.58405f
C212 VP.n19 B 0.604028f
C213 VP.n20 B 0.032386f
C214 VDD2.n0 B 0.028906f
C215 VDD2.n1 B 0.022629f
C216 VDD2.n2 B 0.01216f
C217 VDD2.n3 B 0.028741f
C218 VDD2.n4 B 0.012875f
C219 VDD2.n5 B 0.022629f
C220 VDD2.n6 B 0.01216f
C221 VDD2.n7 B 0.028741f
C222 VDD2.n8 B 0.012875f
C223 VDD2.n9 B 0.022629f
C224 VDD2.n10 B 0.01216f
C225 VDD2.n11 B 0.028741f
C226 VDD2.n12 B 0.012875f
C227 VDD2.n13 B 0.022629f
C228 VDD2.n14 B 0.01216f
C229 VDD2.n15 B 0.028741f
C230 VDD2.n16 B 0.012875f
C231 VDD2.n17 B 0.022629f
C232 VDD2.n18 B 0.01216f
C233 VDD2.n19 B 0.028741f
C234 VDD2.n20 B 0.012875f
C235 VDD2.n21 B 0.022629f
C236 VDD2.n22 B 0.01216f
C237 VDD2.n23 B 0.028741f
C238 VDD2.n24 B 0.012875f
C239 VDD2.n25 B 0.145604f
C240 VDD2.t4 B 0.047363f
C241 VDD2.n26 B 0.021556f
C242 VDD2.n27 B 0.016978f
C243 VDD2.n28 B 0.01216f
C244 VDD2.n29 B 1.43596f
C245 VDD2.n30 B 0.022629f
C246 VDD2.n31 B 0.01216f
C247 VDD2.n32 B 0.012875f
C248 VDD2.n33 B 0.028741f
C249 VDD2.n34 B 0.028741f
C250 VDD2.n35 B 0.012875f
C251 VDD2.n36 B 0.01216f
C252 VDD2.n37 B 0.022629f
C253 VDD2.n38 B 0.022629f
C254 VDD2.n39 B 0.01216f
C255 VDD2.n40 B 0.012875f
C256 VDD2.n41 B 0.028741f
C257 VDD2.n42 B 0.028741f
C258 VDD2.n43 B 0.012875f
C259 VDD2.n44 B 0.01216f
C260 VDD2.n45 B 0.022629f
C261 VDD2.n46 B 0.022629f
C262 VDD2.n47 B 0.01216f
C263 VDD2.n48 B 0.012875f
C264 VDD2.n49 B 0.028741f
C265 VDD2.n50 B 0.028741f
C266 VDD2.n51 B 0.012875f
C267 VDD2.n52 B 0.01216f
C268 VDD2.n53 B 0.022629f
C269 VDD2.n54 B 0.022629f
C270 VDD2.n55 B 0.01216f
C271 VDD2.n56 B 0.012875f
C272 VDD2.n57 B 0.028741f
C273 VDD2.n58 B 0.028741f
C274 VDD2.n59 B 0.012875f
C275 VDD2.n60 B 0.01216f
C276 VDD2.n61 B 0.022629f
C277 VDD2.n62 B 0.022629f
C278 VDD2.n63 B 0.01216f
C279 VDD2.n64 B 0.012875f
C280 VDD2.n65 B 0.028741f
C281 VDD2.n66 B 0.028741f
C282 VDD2.n67 B 0.028741f
C283 VDD2.n68 B 0.012875f
C284 VDD2.n69 B 0.01216f
C285 VDD2.n70 B 0.022629f
C286 VDD2.n71 B 0.022629f
C287 VDD2.n72 B 0.01216f
C288 VDD2.n73 B 0.012517f
C289 VDD2.n74 B 0.012517f
C290 VDD2.n75 B 0.028741f
C291 VDD2.n76 B 0.05709f
C292 VDD2.n77 B 0.012875f
C293 VDD2.n78 B 0.01216f
C294 VDD2.n79 B 0.052614f
C295 VDD2.n80 B 0.04853f
C296 VDD2.t2 B 0.261971f
C297 VDD2.t5 B 0.261971f
C298 VDD2.n81 B 2.3665f
C299 VDD2.n82 B 1.90551f
C300 VDD2.n83 B 0.028906f
C301 VDD2.n84 B 0.022629f
C302 VDD2.n85 B 0.01216f
C303 VDD2.n86 B 0.028741f
C304 VDD2.n87 B 0.012875f
C305 VDD2.n88 B 0.022629f
C306 VDD2.n89 B 0.01216f
C307 VDD2.n90 B 0.028741f
C308 VDD2.n91 B 0.028741f
C309 VDD2.n92 B 0.012875f
C310 VDD2.n93 B 0.022629f
C311 VDD2.n94 B 0.01216f
C312 VDD2.n95 B 0.028741f
C313 VDD2.n96 B 0.012875f
C314 VDD2.n97 B 0.022629f
C315 VDD2.n98 B 0.01216f
C316 VDD2.n99 B 0.028741f
C317 VDD2.n100 B 0.012875f
C318 VDD2.n101 B 0.022629f
C319 VDD2.n102 B 0.01216f
C320 VDD2.n103 B 0.028741f
C321 VDD2.n104 B 0.012875f
C322 VDD2.n105 B 0.022629f
C323 VDD2.n106 B 0.01216f
C324 VDD2.n107 B 0.028741f
C325 VDD2.n108 B 0.012875f
C326 VDD2.n109 B 0.145604f
C327 VDD2.t1 B 0.047363f
C328 VDD2.n110 B 0.021556f
C329 VDD2.n111 B 0.016978f
C330 VDD2.n112 B 0.01216f
C331 VDD2.n113 B 1.43596f
C332 VDD2.n114 B 0.022629f
C333 VDD2.n115 B 0.01216f
C334 VDD2.n116 B 0.012875f
C335 VDD2.n117 B 0.028741f
C336 VDD2.n118 B 0.028741f
C337 VDD2.n119 B 0.012875f
C338 VDD2.n120 B 0.01216f
C339 VDD2.n121 B 0.022629f
C340 VDD2.n122 B 0.022629f
C341 VDD2.n123 B 0.01216f
C342 VDD2.n124 B 0.012875f
C343 VDD2.n125 B 0.028741f
C344 VDD2.n126 B 0.028741f
C345 VDD2.n127 B 0.012875f
C346 VDD2.n128 B 0.01216f
C347 VDD2.n129 B 0.022629f
C348 VDD2.n130 B 0.022629f
C349 VDD2.n131 B 0.01216f
C350 VDD2.n132 B 0.012875f
C351 VDD2.n133 B 0.028741f
C352 VDD2.n134 B 0.028741f
C353 VDD2.n135 B 0.012875f
C354 VDD2.n136 B 0.01216f
C355 VDD2.n137 B 0.022629f
C356 VDD2.n138 B 0.022629f
C357 VDD2.n139 B 0.01216f
C358 VDD2.n140 B 0.012875f
C359 VDD2.n141 B 0.028741f
C360 VDD2.n142 B 0.028741f
C361 VDD2.n143 B 0.012875f
C362 VDD2.n144 B 0.01216f
C363 VDD2.n145 B 0.022629f
C364 VDD2.n146 B 0.022629f
C365 VDD2.n147 B 0.01216f
C366 VDD2.n148 B 0.012875f
C367 VDD2.n149 B 0.028741f
C368 VDD2.n150 B 0.028741f
C369 VDD2.n151 B 0.012875f
C370 VDD2.n152 B 0.01216f
C371 VDD2.n153 B 0.022629f
C372 VDD2.n154 B 0.022629f
C373 VDD2.n155 B 0.01216f
C374 VDD2.n156 B 0.012517f
C375 VDD2.n157 B 0.012517f
C376 VDD2.n158 B 0.028741f
C377 VDD2.n159 B 0.05709f
C378 VDD2.n160 B 0.012875f
C379 VDD2.n161 B 0.01216f
C380 VDD2.n162 B 0.052614f
C381 VDD2.n163 B 0.047049f
C382 VDD2.n164 B 2.08791f
C383 VDD2.t3 B 0.261971f
C384 VDD2.t0 B 0.261971f
C385 VDD2.n165 B 2.36648f
C386 VTAIL.t6 B 0.26942f
C387 VTAIL.t8 B 0.26942f
C388 VTAIL.n0 B 2.36311f
C389 VTAIL.n1 B 0.327769f
C390 VTAIL.n2 B 0.029728f
C391 VTAIL.n3 B 0.023272f
C392 VTAIL.n4 B 0.012506f
C393 VTAIL.n5 B 0.029559f
C394 VTAIL.n6 B 0.013241f
C395 VTAIL.n7 B 0.023272f
C396 VTAIL.n8 B 0.012506f
C397 VTAIL.n9 B 0.029559f
C398 VTAIL.n10 B 0.013241f
C399 VTAIL.n11 B 0.023272f
C400 VTAIL.n12 B 0.012506f
C401 VTAIL.n13 B 0.029559f
C402 VTAIL.n14 B 0.013241f
C403 VTAIL.n15 B 0.023272f
C404 VTAIL.n16 B 0.012506f
C405 VTAIL.n17 B 0.029559f
C406 VTAIL.n18 B 0.013241f
C407 VTAIL.n19 B 0.023272f
C408 VTAIL.n20 B 0.012506f
C409 VTAIL.n21 B 0.029559f
C410 VTAIL.n22 B 0.013241f
C411 VTAIL.n23 B 0.023272f
C412 VTAIL.n24 B 0.012506f
C413 VTAIL.n25 B 0.029559f
C414 VTAIL.n26 B 0.013241f
C415 VTAIL.n27 B 0.149745f
C416 VTAIL.t4 B 0.04871f
C417 VTAIL.n28 B 0.022169f
C418 VTAIL.n29 B 0.017461f
C419 VTAIL.n30 B 0.012506f
C420 VTAIL.n31 B 1.4768f
C421 VTAIL.n32 B 0.023272f
C422 VTAIL.n33 B 0.012506f
C423 VTAIL.n34 B 0.013241f
C424 VTAIL.n35 B 0.029559f
C425 VTAIL.n36 B 0.029559f
C426 VTAIL.n37 B 0.013241f
C427 VTAIL.n38 B 0.012506f
C428 VTAIL.n39 B 0.023272f
C429 VTAIL.n40 B 0.023272f
C430 VTAIL.n41 B 0.012506f
C431 VTAIL.n42 B 0.013241f
C432 VTAIL.n43 B 0.029559f
C433 VTAIL.n44 B 0.029559f
C434 VTAIL.n45 B 0.013241f
C435 VTAIL.n46 B 0.012506f
C436 VTAIL.n47 B 0.023272f
C437 VTAIL.n48 B 0.023272f
C438 VTAIL.n49 B 0.012506f
C439 VTAIL.n50 B 0.013241f
C440 VTAIL.n51 B 0.029559f
C441 VTAIL.n52 B 0.029559f
C442 VTAIL.n53 B 0.013241f
C443 VTAIL.n54 B 0.012506f
C444 VTAIL.n55 B 0.023272f
C445 VTAIL.n56 B 0.023272f
C446 VTAIL.n57 B 0.012506f
C447 VTAIL.n58 B 0.013241f
C448 VTAIL.n59 B 0.029559f
C449 VTAIL.n60 B 0.029559f
C450 VTAIL.n61 B 0.013241f
C451 VTAIL.n62 B 0.012506f
C452 VTAIL.n63 B 0.023272f
C453 VTAIL.n64 B 0.023272f
C454 VTAIL.n65 B 0.012506f
C455 VTAIL.n66 B 0.013241f
C456 VTAIL.n67 B 0.029559f
C457 VTAIL.n68 B 0.029559f
C458 VTAIL.n69 B 0.029559f
C459 VTAIL.n70 B 0.013241f
C460 VTAIL.n71 B 0.012506f
C461 VTAIL.n72 B 0.023272f
C462 VTAIL.n73 B 0.023272f
C463 VTAIL.n74 B 0.012506f
C464 VTAIL.n75 B 0.012873f
C465 VTAIL.n76 B 0.012873f
C466 VTAIL.n77 B 0.029559f
C467 VTAIL.n78 B 0.058713f
C468 VTAIL.n79 B 0.013241f
C469 VTAIL.n80 B 0.012506f
C470 VTAIL.n81 B 0.054111f
C471 VTAIL.n82 B 0.03232f
C472 VTAIL.n83 B 0.175528f
C473 VTAIL.t11 B 0.26942f
C474 VTAIL.t1 B 0.26942f
C475 VTAIL.n84 B 2.36311f
C476 VTAIL.n85 B 1.73171f
C477 VTAIL.t9 B 0.26942f
C478 VTAIL.t7 B 0.26942f
C479 VTAIL.n86 B 2.36312f
C480 VTAIL.n87 B 1.7317f
C481 VTAIL.n88 B 0.029728f
C482 VTAIL.n89 B 0.023272f
C483 VTAIL.n90 B 0.012506f
C484 VTAIL.n91 B 0.029559f
C485 VTAIL.n92 B 0.013241f
C486 VTAIL.n93 B 0.023272f
C487 VTAIL.n94 B 0.012506f
C488 VTAIL.n95 B 0.029559f
C489 VTAIL.n96 B 0.029559f
C490 VTAIL.n97 B 0.013241f
C491 VTAIL.n98 B 0.023272f
C492 VTAIL.n99 B 0.012506f
C493 VTAIL.n100 B 0.029559f
C494 VTAIL.n101 B 0.013241f
C495 VTAIL.n102 B 0.023272f
C496 VTAIL.n103 B 0.012506f
C497 VTAIL.n104 B 0.029559f
C498 VTAIL.n105 B 0.013241f
C499 VTAIL.n106 B 0.023272f
C500 VTAIL.n107 B 0.012506f
C501 VTAIL.n108 B 0.029559f
C502 VTAIL.n109 B 0.013241f
C503 VTAIL.n110 B 0.023272f
C504 VTAIL.n111 B 0.012506f
C505 VTAIL.n112 B 0.029559f
C506 VTAIL.n113 B 0.013241f
C507 VTAIL.n114 B 0.149745f
C508 VTAIL.t10 B 0.04871f
C509 VTAIL.n115 B 0.022169f
C510 VTAIL.n116 B 0.017461f
C511 VTAIL.n117 B 0.012506f
C512 VTAIL.n118 B 1.4768f
C513 VTAIL.n119 B 0.023272f
C514 VTAIL.n120 B 0.012506f
C515 VTAIL.n121 B 0.013241f
C516 VTAIL.n122 B 0.029559f
C517 VTAIL.n123 B 0.029559f
C518 VTAIL.n124 B 0.013241f
C519 VTAIL.n125 B 0.012506f
C520 VTAIL.n126 B 0.023272f
C521 VTAIL.n127 B 0.023272f
C522 VTAIL.n128 B 0.012506f
C523 VTAIL.n129 B 0.013241f
C524 VTAIL.n130 B 0.029559f
C525 VTAIL.n131 B 0.029559f
C526 VTAIL.n132 B 0.013241f
C527 VTAIL.n133 B 0.012506f
C528 VTAIL.n134 B 0.023272f
C529 VTAIL.n135 B 0.023272f
C530 VTAIL.n136 B 0.012506f
C531 VTAIL.n137 B 0.013241f
C532 VTAIL.n138 B 0.029559f
C533 VTAIL.n139 B 0.029559f
C534 VTAIL.n140 B 0.013241f
C535 VTAIL.n141 B 0.012506f
C536 VTAIL.n142 B 0.023272f
C537 VTAIL.n143 B 0.023272f
C538 VTAIL.n144 B 0.012506f
C539 VTAIL.n145 B 0.013241f
C540 VTAIL.n146 B 0.029559f
C541 VTAIL.n147 B 0.029559f
C542 VTAIL.n148 B 0.013241f
C543 VTAIL.n149 B 0.012506f
C544 VTAIL.n150 B 0.023272f
C545 VTAIL.n151 B 0.023272f
C546 VTAIL.n152 B 0.012506f
C547 VTAIL.n153 B 0.013241f
C548 VTAIL.n154 B 0.029559f
C549 VTAIL.n155 B 0.029559f
C550 VTAIL.n156 B 0.013241f
C551 VTAIL.n157 B 0.012506f
C552 VTAIL.n158 B 0.023272f
C553 VTAIL.n159 B 0.023272f
C554 VTAIL.n160 B 0.012506f
C555 VTAIL.n161 B 0.012873f
C556 VTAIL.n162 B 0.012873f
C557 VTAIL.n163 B 0.029559f
C558 VTAIL.n164 B 0.058713f
C559 VTAIL.n165 B 0.013241f
C560 VTAIL.n166 B 0.012506f
C561 VTAIL.n167 B 0.054111f
C562 VTAIL.n168 B 0.03232f
C563 VTAIL.n169 B 0.175528f
C564 VTAIL.t3 B 0.26942f
C565 VTAIL.t0 B 0.26942f
C566 VTAIL.n170 B 2.36312f
C567 VTAIL.n171 B 0.383513f
C568 VTAIL.n172 B 0.029728f
C569 VTAIL.n173 B 0.023272f
C570 VTAIL.n174 B 0.012506f
C571 VTAIL.n175 B 0.029559f
C572 VTAIL.n176 B 0.013241f
C573 VTAIL.n177 B 0.023272f
C574 VTAIL.n178 B 0.012506f
C575 VTAIL.n179 B 0.029559f
C576 VTAIL.n180 B 0.029559f
C577 VTAIL.n181 B 0.013241f
C578 VTAIL.n182 B 0.023272f
C579 VTAIL.n183 B 0.012506f
C580 VTAIL.n184 B 0.029559f
C581 VTAIL.n185 B 0.013241f
C582 VTAIL.n186 B 0.023272f
C583 VTAIL.n187 B 0.012506f
C584 VTAIL.n188 B 0.029559f
C585 VTAIL.n189 B 0.013241f
C586 VTAIL.n190 B 0.023272f
C587 VTAIL.n191 B 0.012506f
C588 VTAIL.n192 B 0.029559f
C589 VTAIL.n193 B 0.013241f
C590 VTAIL.n194 B 0.023272f
C591 VTAIL.n195 B 0.012506f
C592 VTAIL.n196 B 0.029559f
C593 VTAIL.n197 B 0.013241f
C594 VTAIL.n198 B 0.149745f
C595 VTAIL.t2 B 0.04871f
C596 VTAIL.n199 B 0.022169f
C597 VTAIL.n200 B 0.017461f
C598 VTAIL.n201 B 0.012506f
C599 VTAIL.n202 B 1.4768f
C600 VTAIL.n203 B 0.023272f
C601 VTAIL.n204 B 0.012506f
C602 VTAIL.n205 B 0.013241f
C603 VTAIL.n206 B 0.029559f
C604 VTAIL.n207 B 0.029559f
C605 VTAIL.n208 B 0.013241f
C606 VTAIL.n209 B 0.012506f
C607 VTAIL.n210 B 0.023272f
C608 VTAIL.n211 B 0.023272f
C609 VTAIL.n212 B 0.012506f
C610 VTAIL.n213 B 0.013241f
C611 VTAIL.n214 B 0.029559f
C612 VTAIL.n215 B 0.029559f
C613 VTAIL.n216 B 0.013241f
C614 VTAIL.n217 B 0.012506f
C615 VTAIL.n218 B 0.023272f
C616 VTAIL.n219 B 0.023272f
C617 VTAIL.n220 B 0.012506f
C618 VTAIL.n221 B 0.013241f
C619 VTAIL.n222 B 0.029559f
C620 VTAIL.n223 B 0.029559f
C621 VTAIL.n224 B 0.013241f
C622 VTAIL.n225 B 0.012506f
C623 VTAIL.n226 B 0.023272f
C624 VTAIL.n227 B 0.023272f
C625 VTAIL.n228 B 0.012506f
C626 VTAIL.n229 B 0.013241f
C627 VTAIL.n230 B 0.029559f
C628 VTAIL.n231 B 0.029559f
C629 VTAIL.n232 B 0.013241f
C630 VTAIL.n233 B 0.012506f
C631 VTAIL.n234 B 0.023272f
C632 VTAIL.n235 B 0.023272f
C633 VTAIL.n236 B 0.012506f
C634 VTAIL.n237 B 0.013241f
C635 VTAIL.n238 B 0.029559f
C636 VTAIL.n239 B 0.029559f
C637 VTAIL.n240 B 0.013241f
C638 VTAIL.n241 B 0.012506f
C639 VTAIL.n242 B 0.023272f
C640 VTAIL.n243 B 0.023272f
C641 VTAIL.n244 B 0.012506f
C642 VTAIL.n245 B 0.012873f
C643 VTAIL.n246 B 0.012873f
C644 VTAIL.n247 B 0.029559f
C645 VTAIL.n248 B 0.058713f
C646 VTAIL.n249 B 0.013241f
C647 VTAIL.n250 B 0.012506f
C648 VTAIL.n251 B 0.054111f
C649 VTAIL.n252 B 0.03232f
C650 VTAIL.n253 B 1.44356f
C651 VTAIL.n254 B 0.029728f
C652 VTAIL.n255 B 0.023272f
C653 VTAIL.n256 B 0.012506f
C654 VTAIL.n257 B 0.029559f
C655 VTAIL.n258 B 0.013241f
C656 VTAIL.n259 B 0.023272f
C657 VTAIL.n260 B 0.012506f
C658 VTAIL.n261 B 0.029559f
C659 VTAIL.n262 B 0.013241f
C660 VTAIL.n263 B 0.023272f
C661 VTAIL.n264 B 0.012506f
C662 VTAIL.n265 B 0.029559f
C663 VTAIL.n266 B 0.013241f
C664 VTAIL.n267 B 0.023272f
C665 VTAIL.n268 B 0.012506f
C666 VTAIL.n269 B 0.029559f
C667 VTAIL.n270 B 0.013241f
C668 VTAIL.n271 B 0.023272f
C669 VTAIL.n272 B 0.012506f
C670 VTAIL.n273 B 0.029559f
C671 VTAIL.n274 B 0.013241f
C672 VTAIL.n275 B 0.023272f
C673 VTAIL.n276 B 0.012506f
C674 VTAIL.n277 B 0.029559f
C675 VTAIL.n278 B 0.013241f
C676 VTAIL.n279 B 0.149745f
C677 VTAIL.t5 B 0.04871f
C678 VTAIL.n280 B 0.022169f
C679 VTAIL.n281 B 0.017461f
C680 VTAIL.n282 B 0.012506f
C681 VTAIL.n283 B 1.4768f
C682 VTAIL.n284 B 0.023272f
C683 VTAIL.n285 B 0.012506f
C684 VTAIL.n286 B 0.013241f
C685 VTAIL.n287 B 0.029559f
C686 VTAIL.n288 B 0.029559f
C687 VTAIL.n289 B 0.013241f
C688 VTAIL.n290 B 0.012506f
C689 VTAIL.n291 B 0.023272f
C690 VTAIL.n292 B 0.023272f
C691 VTAIL.n293 B 0.012506f
C692 VTAIL.n294 B 0.013241f
C693 VTAIL.n295 B 0.029559f
C694 VTAIL.n296 B 0.029559f
C695 VTAIL.n297 B 0.013241f
C696 VTAIL.n298 B 0.012506f
C697 VTAIL.n299 B 0.023272f
C698 VTAIL.n300 B 0.023272f
C699 VTAIL.n301 B 0.012506f
C700 VTAIL.n302 B 0.013241f
C701 VTAIL.n303 B 0.029559f
C702 VTAIL.n304 B 0.029559f
C703 VTAIL.n305 B 0.013241f
C704 VTAIL.n306 B 0.012506f
C705 VTAIL.n307 B 0.023272f
C706 VTAIL.n308 B 0.023272f
C707 VTAIL.n309 B 0.012506f
C708 VTAIL.n310 B 0.013241f
C709 VTAIL.n311 B 0.029559f
C710 VTAIL.n312 B 0.029559f
C711 VTAIL.n313 B 0.013241f
C712 VTAIL.n314 B 0.012506f
C713 VTAIL.n315 B 0.023272f
C714 VTAIL.n316 B 0.023272f
C715 VTAIL.n317 B 0.012506f
C716 VTAIL.n318 B 0.013241f
C717 VTAIL.n319 B 0.029559f
C718 VTAIL.n320 B 0.029559f
C719 VTAIL.n321 B 0.029559f
C720 VTAIL.n322 B 0.013241f
C721 VTAIL.n323 B 0.012506f
C722 VTAIL.n324 B 0.023272f
C723 VTAIL.n325 B 0.023272f
C724 VTAIL.n326 B 0.012506f
C725 VTAIL.n327 B 0.012873f
C726 VTAIL.n328 B 0.012873f
C727 VTAIL.n329 B 0.029559f
C728 VTAIL.n330 B 0.058713f
C729 VTAIL.n331 B 0.013241f
C730 VTAIL.n332 B 0.012506f
C731 VTAIL.n333 B 0.054111f
C732 VTAIL.n334 B 0.03232f
C733 VTAIL.n335 B 1.41915f
C734 VN.n0 B 0.041171f
C735 VN.t3 B 1.50318f
C736 VN.n1 B 0.589581f
C737 VN.t1 B 1.58416f
C738 VN.n2 B 0.601174f
C739 VN.n3 B 0.173723f
C740 VN.n4 B 0.054109f
C741 VN.n5 B 0.013689f
C742 VN.t0 B 1.56058f
C743 VN.n6 B 0.595076f
C744 VN.n7 B 0.031906f
C745 VN.n8 B 0.041171f
C746 VN.t2 B 1.50318f
C747 VN.n9 B 0.589581f
C748 VN.t5 B 1.58416f
C749 VN.n10 B 0.601174f
C750 VN.n11 B 0.173723f
C751 VN.n12 B 0.054109f
C752 VN.n13 B 0.013689f
C753 VN.t4 B 1.56058f
C754 VN.n14 B 0.595076f
C755 VN.n15 B 1.86478f
.ends

